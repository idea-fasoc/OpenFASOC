* NGSPICE file created from diff_pair_sample_0816.ext - technology: sky130A

.subckt diff_pair_sample_0816 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=0 ps=0 w=18.88 l=3.91
X2 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=0 ps=0 w=18.88 l=3.91
X3 VTAIL.t13 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=3.1152 ps=19.21 w=18.88 l=3.91
X4 VTAIL.t9 VN.t1 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=3.1152 ps=19.21 w=18.88 l=3.91
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=0 ps=0 w=18.88 l=3.91
X6 VTAIL.t15 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X7 VTAIL.t8 VN.t2 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X8 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X9 VDD1.t4 VP.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=7.3632 ps=38.54 w=18.88 l=3.91
X10 VDD2.t6 VN.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=7.3632 ps=38.54 w=18.88 l=3.91
X11 VTAIL.t6 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=3.1152 ps=19.21 w=18.88 l=3.91
X12 VDD2.t2 VN.t5 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=7.3632 ps=38.54 w=18.88 l=3.91
X13 VDD1.t3 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X14 VDD1.t2 VP.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=7.3632 ps=38.54 w=18.88 l=3.91
X15 VTAIL.t0 VP.t6 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X16 VDD2.t1 VN.t6 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X17 VTAIL.t14 VP.t7 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=3.1152 ps=19.21 w=18.88 l=3.91
X18 VDD2.t0 VN.t7 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1152 pd=19.21 as=3.1152 ps=19.21 w=18.88 l=3.91
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.3632 pd=38.54 as=0 ps=0 w=18.88 l=3.91
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n42 161.3
R7 VN.n65 VN.n64 161.3
R8 VN.n62 VN.n43 161.3
R9 VN.n61 VN.n60 161.3
R10 VN.n59 VN.n44 161.3
R11 VN.n58 VN.n57 161.3
R12 VN.n56 VN.n45 161.3
R13 VN.n55 VN.n54 161.3
R14 VN.n53 VN.n46 161.3
R15 VN.n52 VN.n51 161.3
R16 VN.n50 VN.n47 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n3 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n23 VN.n4 161.3
R26 VN.n22 VN.n21 161.3
R27 VN.n20 VN.n5 161.3
R28 VN.n19 VN.n18 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n9 VN.t1 148.778
R35 VN.n48 VN.t3 148.778
R36 VN.n10 VN.t7 116.371
R37 VN.n24 VN.t0 116.371
R38 VN.n37 VN.t5 116.371
R39 VN.n49 VN.t2 116.371
R40 VN.n63 VN.t6 116.371
R41 VN.n76 VN.t4 116.371
R42 VN.n10 VN.n9 69.3059
R43 VN.n49 VN.n48 69.3059
R44 VN.n38 VN.n37 64.6738
R45 VN.n77 VN.n76 64.6738
R46 VN VN.n77 62.4589
R47 VN.n31 VN.n30 56.5617
R48 VN.n70 VN.n69 56.5617
R49 VN.n17 VN.n16 40.577
R50 VN.n18 VN.n17 40.577
R51 VN.n56 VN.n55 40.577
R52 VN.n57 VN.n56 40.577
R53 VN.n12 VN.n11 24.5923
R54 VN.n12 VN.n7 24.5923
R55 VN.n16 VN.n7 24.5923
R56 VN.n18 VN.n5 24.5923
R57 VN.n22 VN.n5 24.5923
R58 VN.n23 VN.n22 24.5923
R59 VN.n25 VN.n3 24.5923
R60 VN.n29 VN.n3 24.5923
R61 VN.n30 VN.n29 24.5923
R62 VN.n31 VN.n1 24.5923
R63 VN.n35 VN.n1 24.5923
R64 VN.n36 VN.n35 24.5923
R65 VN.n55 VN.n46 24.5923
R66 VN.n51 VN.n46 24.5923
R67 VN.n51 VN.n50 24.5923
R68 VN.n69 VN.n68 24.5923
R69 VN.n68 VN.n42 24.5923
R70 VN.n64 VN.n42 24.5923
R71 VN.n62 VN.n61 24.5923
R72 VN.n61 VN.n44 24.5923
R73 VN.n57 VN.n44 24.5923
R74 VN.n75 VN.n74 24.5923
R75 VN.n74 VN.n40 24.5923
R76 VN.n70 VN.n40 24.5923
R77 VN.n25 VN.n24 18.6903
R78 VN.n64 VN.n63 18.6903
R79 VN.n37 VN.n36 17.7066
R80 VN.n76 VN.n75 17.7066
R81 VN.n11 VN.n10 5.90254
R82 VN.n24 VN.n23 5.90254
R83 VN.n50 VN.n49 5.90254
R84 VN.n63 VN.n62 5.90254
R85 VN.n48 VN.n47 2.76475
R86 VN.n9 VN.n8 2.76475
R87 VN.n77 VN.n39 0.417304
R88 VN.n38 VN.n0 0.417304
R89 VN VN.n38 0.394524
R90 VN.n73 VN.n39 0.189894
R91 VN.n73 VN.n72 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n41 0.189894
R94 VN.n67 VN.n41 0.189894
R95 VN.n67 VN.n66 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n43 0.189894
R98 VN.n60 VN.n43 0.189894
R99 VN.n60 VN.n59 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n45 0.189894
R102 VN.n54 VN.n45 0.189894
R103 VN.n54 VN.n53 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n47 0.189894
R106 VN.n13 VN.n8 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n15 VN.n14 0.189894
R109 VN.n15 VN.n6 0.189894
R110 VN.n19 VN.n6 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n21 VN.n20 0.189894
R113 VN.n21 VN.n4 0.189894
R114 VN.n26 VN.n4 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n28 VN.n27 0.189894
R117 VN.n28 VN.n2 0.189894
R118 VN.n32 VN.n2 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n34 VN.n33 0.189894
R121 VN.n34 VN.n0 0.189894
R122 VDD2.n2 VDD2.n1 60.8427
R123 VDD2.n2 VDD2.n0 60.8427
R124 VDD2 VDD2.n5 60.8397
R125 VDD2.n4 VDD2.n3 59.0705
R126 VDD2.n4 VDD2.n2 56.4394
R127 VDD2 VDD2.n4 1.88628
R128 VDD2.n5 VDD2.t3 1.04923
R129 VDD2.n5 VDD2.t6 1.04923
R130 VDD2.n3 VDD2.t5 1.04923
R131 VDD2.n3 VDD2.t1 1.04923
R132 VDD2.n1 VDD2.t7 1.04923
R133 VDD2.n1 VDD2.t2 1.04923
R134 VDD2.n0 VDD2.t4 1.04923
R135 VDD2.n0 VDD2.t0 1.04923
R136 VTAIL.n850 VTAIL.n750 289.615
R137 VTAIL.n102 VTAIL.n2 289.615
R138 VTAIL.n208 VTAIL.n108 289.615
R139 VTAIL.n316 VTAIL.n216 289.615
R140 VTAIL.n744 VTAIL.n644 289.615
R141 VTAIL.n636 VTAIL.n536 289.615
R142 VTAIL.n530 VTAIL.n430 289.615
R143 VTAIL.n422 VTAIL.n322 289.615
R144 VTAIL.n785 VTAIL.n784 185
R145 VTAIL.n782 VTAIL.n781 185
R146 VTAIL.n791 VTAIL.n790 185
R147 VTAIL.n793 VTAIL.n792 185
R148 VTAIL.n778 VTAIL.n777 185
R149 VTAIL.n799 VTAIL.n798 185
R150 VTAIL.n801 VTAIL.n800 185
R151 VTAIL.n774 VTAIL.n773 185
R152 VTAIL.n807 VTAIL.n806 185
R153 VTAIL.n809 VTAIL.n808 185
R154 VTAIL.n770 VTAIL.n769 185
R155 VTAIL.n815 VTAIL.n814 185
R156 VTAIL.n817 VTAIL.n816 185
R157 VTAIL.n766 VTAIL.n765 185
R158 VTAIL.n823 VTAIL.n822 185
R159 VTAIL.n826 VTAIL.n825 185
R160 VTAIL.n824 VTAIL.n762 185
R161 VTAIL.n831 VTAIL.n761 185
R162 VTAIL.n833 VTAIL.n832 185
R163 VTAIL.n835 VTAIL.n834 185
R164 VTAIL.n758 VTAIL.n757 185
R165 VTAIL.n841 VTAIL.n840 185
R166 VTAIL.n843 VTAIL.n842 185
R167 VTAIL.n754 VTAIL.n753 185
R168 VTAIL.n849 VTAIL.n848 185
R169 VTAIL.n851 VTAIL.n850 185
R170 VTAIL.n37 VTAIL.n36 185
R171 VTAIL.n34 VTAIL.n33 185
R172 VTAIL.n43 VTAIL.n42 185
R173 VTAIL.n45 VTAIL.n44 185
R174 VTAIL.n30 VTAIL.n29 185
R175 VTAIL.n51 VTAIL.n50 185
R176 VTAIL.n53 VTAIL.n52 185
R177 VTAIL.n26 VTAIL.n25 185
R178 VTAIL.n59 VTAIL.n58 185
R179 VTAIL.n61 VTAIL.n60 185
R180 VTAIL.n22 VTAIL.n21 185
R181 VTAIL.n67 VTAIL.n66 185
R182 VTAIL.n69 VTAIL.n68 185
R183 VTAIL.n18 VTAIL.n17 185
R184 VTAIL.n75 VTAIL.n74 185
R185 VTAIL.n78 VTAIL.n77 185
R186 VTAIL.n76 VTAIL.n14 185
R187 VTAIL.n83 VTAIL.n13 185
R188 VTAIL.n85 VTAIL.n84 185
R189 VTAIL.n87 VTAIL.n86 185
R190 VTAIL.n10 VTAIL.n9 185
R191 VTAIL.n93 VTAIL.n92 185
R192 VTAIL.n95 VTAIL.n94 185
R193 VTAIL.n6 VTAIL.n5 185
R194 VTAIL.n101 VTAIL.n100 185
R195 VTAIL.n103 VTAIL.n102 185
R196 VTAIL.n143 VTAIL.n142 185
R197 VTAIL.n140 VTAIL.n139 185
R198 VTAIL.n149 VTAIL.n148 185
R199 VTAIL.n151 VTAIL.n150 185
R200 VTAIL.n136 VTAIL.n135 185
R201 VTAIL.n157 VTAIL.n156 185
R202 VTAIL.n159 VTAIL.n158 185
R203 VTAIL.n132 VTAIL.n131 185
R204 VTAIL.n165 VTAIL.n164 185
R205 VTAIL.n167 VTAIL.n166 185
R206 VTAIL.n128 VTAIL.n127 185
R207 VTAIL.n173 VTAIL.n172 185
R208 VTAIL.n175 VTAIL.n174 185
R209 VTAIL.n124 VTAIL.n123 185
R210 VTAIL.n181 VTAIL.n180 185
R211 VTAIL.n184 VTAIL.n183 185
R212 VTAIL.n182 VTAIL.n120 185
R213 VTAIL.n189 VTAIL.n119 185
R214 VTAIL.n191 VTAIL.n190 185
R215 VTAIL.n193 VTAIL.n192 185
R216 VTAIL.n116 VTAIL.n115 185
R217 VTAIL.n199 VTAIL.n198 185
R218 VTAIL.n201 VTAIL.n200 185
R219 VTAIL.n112 VTAIL.n111 185
R220 VTAIL.n207 VTAIL.n206 185
R221 VTAIL.n209 VTAIL.n208 185
R222 VTAIL.n251 VTAIL.n250 185
R223 VTAIL.n248 VTAIL.n247 185
R224 VTAIL.n257 VTAIL.n256 185
R225 VTAIL.n259 VTAIL.n258 185
R226 VTAIL.n244 VTAIL.n243 185
R227 VTAIL.n265 VTAIL.n264 185
R228 VTAIL.n267 VTAIL.n266 185
R229 VTAIL.n240 VTAIL.n239 185
R230 VTAIL.n273 VTAIL.n272 185
R231 VTAIL.n275 VTAIL.n274 185
R232 VTAIL.n236 VTAIL.n235 185
R233 VTAIL.n281 VTAIL.n280 185
R234 VTAIL.n283 VTAIL.n282 185
R235 VTAIL.n232 VTAIL.n231 185
R236 VTAIL.n289 VTAIL.n288 185
R237 VTAIL.n292 VTAIL.n291 185
R238 VTAIL.n290 VTAIL.n228 185
R239 VTAIL.n297 VTAIL.n227 185
R240 VTAIL.n299 VTAIL.n298 185
R241 VTAIL.n301 VTAIL.n300 185
R242 VTAIL.n224 VTAIL.n223 185
R243 VTAIL.n307 VTAIL.n306 185
R244 VTAIL.n309 VTAIL.n308 185
R245 VTAIL.n220 VTAIL.n219 185
R246 VTAIL.n315 VTAIL.n314 185
R247 VTAIL.n317 VTAIL.n316 185
R248 VTAIL.n745 VTAIL.n744 185
R249 VTAIL.n743 VTAIL.n742 185
R250 VTAIL.n648 VTAIL.n647 185
R251 VTAIL.n737 VTAIL.n736 185
R252 VTAIL.n735 VTAIL.n734 185
R253 VTAIL.n652 VTAIL.n651 185
R254 VTAIL.n729 VTAIL.n728 185
R255 VTAIL.n727 VTAIL.n726 185
R256 VTAIL.n725 VTAIL.n655 185
R257 VTAIL.n659 VTAIL.n656 185
R258 VTAIL.n720 VTAIL.n719 185
R259 VTAIL.n718 VTAIL.n717 185
R260 VTAIL.n661 VTAIL.n660 185
R261 VTAIL.n712 VTAIL.n711 185
R262 VTAIL.n710 VTAIL.n709 185
R263 VTAIL.n665 VTAIL.n664 185
R264 VTAIL.n704 VTAIL.n703 185
R265 VTAIL.n702 VTAIL.n701 185
R266 VTAIL.n669 VTAIL.n668 185
R267 VTAIL.n696 VTAIL.n695 185
R268 VTAIL.n694 VTAIL.n693 185
R269 VTAIL.n673 VTAIL.n672 185
R270 VTAIL.n688 VTAIL.n687 185
R271 VTAIL.n686 VTAIL.n685 185
R272 VTAIL.n677 VTAIL.n676 185
R273 VTAIL.n680 VTAIL.n679 185
R274 VTAIL.n637 VTAIL.n636 185
R275 VTAIL.n635 VTAIL.n634 185
R276 VTAIL.n540 VTAIL.n539 185
R277 VTAIL.n629 VTAIL.n628 185
R278 VTAIL.n627 VTAIL.n626 185
R279 VTAIL.n544 VTAIL.n543 185
R280 VTAIL.n621 VTAIL.n620 185
R281 VTAIL.n619 VTAIL.n618 185
R282 VTAIL.n617 VTAIL.n547 185
R283 VTAIL.n551 VTAIL.n548 185
R284 VTAIL.n612 VTAIL.n611 185
R285 VTAIL.n610 VTAIL.n609 185
R286 VTAIL.n553 VTAIL.n552 185
R287 VTAIL.n604 VTAIL.n603 185
R288 VTAIL.n602 VTAIL.n601 185
R289 VTAIL.n557 VTAIL.n556 185
R290 VTAIL.n596 VTAIL.n595 185
R291 VTAIL.n594 VTAIL.n593 185
R292 VTAIL.n561 VTAIL.n560 185
R293 VTAIL.n588 VTAIL.n587 185
R294 VTAIL.n586 VTAIL.n585 185
R295 VTAIL.n565 VTAIL.n564 185
R296 VTAIL.n580 VTAIL.n579 185
R297 VTAIL.n578 VTAIL.n577 185
R298 VTAIL.n569 VTAIL.n568 185
R299 VTAIL.n572 VTAIL.n571 185
R300 VTAIL.n531 VTAIL.n530 185
R301 VTAIL.n529 VTAIL.n528 185
R302 VTAIL.n434 VTAIL.n433 185
R303 VTAIL.n523 VTAIL.n522 185
R304 VTAIL.n521 VTAIL.n520 185
R305 VTAIL.n438 VTAIL.n437 185
R306 VTAIL.n515 VTAIL.n514 185
R307 VTAIL.n513 VTAIL.n512 185
R308 VTAIL.n511 VTAIL.n441 185
R309 VTAIL.n445 VTAIL.n442 185
R310 VTAIL.n506 VTAIL.n505 185
R311 VTAIL.n504 VTAIL.n503 185
R312 VTAIL.n447 VTAIL.n446 185
R313 VTAIL.n498 VTAIL.n497 185
R314 VTAIL.n496 VTAIL.n495 185
R315 VTAIL.n451 VTAIL.n450 185
R316 VTAIL.n490 VTAIL.n489 185
R317 VTAIL.n488 VTAIL.n487 185
R318 VTAIL.n455 VTAIL.n454 185
R319 VTAIL.n482 VTAIL.n481 185
R320 VTAIL.n480 VTAIL.n479 185
R321 VTAIL.n459 VTAIL.n458 185
R322 VTAIL.n474 VTAIL.n473 185
R323 VTAIL.n472 VTAIL.n471 185
R324 VTAIL.n463 VTAIL.n462 185
R325 VTAIL.n466 VTAIL.n465 185
R326 VTAIL.n423 VTAIL.n422 185
R327 VTAIL.n421 VTAIL.n420 185
R328 VTAIL.n326 VTAIL.n325 185
R329 VTAIL.n415 VTAIL.n414 185
R330 VTAIL.n413 VTAIL.n412 185
R331 VTAIL.n330 VTAIL.n329 185
R332 VTAIL.n407 VTAIL.n406 185
R333 VTAIL.n405 VTAIL.n404 185
R334 VTAIL.n403 VTAIL.n333 185
R335 VTAIL.n337 VTAIL.n334 185
R336 VTAIL.n398 VTAIL.n397 185
R337 VTAIL.n396 VTAIL.n395 185
R338 VTAIL.n339 VTAIL.n338 185
R339 VTAIL.n390 VTAIL.n389 185
R340 VTAIL.n388 VTAIL.n387 185
R341 VTAIL.n343 VTAIL.n342 185
R342 VTAIL.n382 VTAIL.n381 185
R343 VTAIL.n380 VTAIL.n379 185
R344 VTAIL.n347 VTAIL.n346 185
R345 VTAIL.n374 VTAIL.n373 185
R346 VTAIL.n372 VTAIL.n371 185
R347 VTAIL.n351 VTAIL.n350 185
R348 VTAIL.n366 VTAIL.n365 185
R349 VTAIL.n364 VTAIL.n363 185
R350 VTAIL.n355 VTAIL.n354 185
R351 VTAIL.n358 VTAIL.n357 185
R352 VTAIL.t12 VTAIL.n678 147.659
R353 VTAIL.t14 VTAIL.n570 147.659
R354 VTAIL.t7 VTAIL.n464 147.659
R355 VTAIL.t6 VTAIL.n356 147.659
R356 VTAIL.t5 VTAIL.n783 147.659
R357 VTAIL.t9 VTAIL.n35 147.659
R358 VTAIL.t11 VTAIL.n141 147.659
R359 VTAIL.t13 VTAIL.n249 147.659
R360 VTAIL.n784 VTAIL.n781 104.615
R361 VTAIL.n791 VTAIL.n781 104.615
R362 VTAIL.n792 VTAIL.n791 104.615
R363 VTAIL.n792 VTAIL.n777 104.615
R364 VTAIL.n799 VTAIL.n777 104.615
R365 VTAIL.n800 VTAIL.n799 104.615
R366 VTAIL.n800 VTAIL.n773 104.615
R367 VTAIL.n807 VTAIL.n773 104.615
R368 VTAIL.n808 VTAIL.n807 104.615
R369 VTAIL.n808 VTAIL.n769 104.615
R370 VTAIL.n815 VTAIL.n769 104.615
R371 VTAIL.n816 VTAIL.n815 104.615
R372 VTAIL.n816 VTAIL.n765 104.615
R373 VTAIL.n823 VTAIL.n765 104.615
R374 VTAIL.n825 VTAIL.n823 104.615
R375 VTAIL.n825 VTAIL.n824 104.615
R376 VTAIL.n824 VTAIL.n761 104.615
R377 VTAIL.n833 VTAIL.n761 104.615
R378 VTAIL.n834 VTAIL.n833 104.615
R379 VTAIL.n834 VTAIL.n757 104.615
R380 VTAIL.n841 VTAIL.n757 104.615
R381 VTAIL.n842 VTAIL.n841 104.615
R382 VTAIL.n842 VTAIL.n753 104.615
R383 VTAIL.n849 VTAIL.n753 104.615
R384 VTAIL.n850 VTAIL.n849 104.615
R385 VTAIL.n36 VTAIL.n33 104.615
R386 VTAIL.n43 VTAIL.n33 104.615
R387 VTAIL.n44 VTAIL.n43 104.615
R388 VTAIL.n44 VTAIL.n29 104.615
R389 VTAIL.n51 VTAIL.n29 104.615
R390 VTAIL.n52 VTAIL.n51 104.615
R391 VTAIL.n52 VTAIL.n25 104.615
R392 VTAIL.n59 VTAIL.n25 104.615
R393 VTAIL.n60 VTAIL.n59 104.615
R394 VTAIL.n60 VTAIL.n21 104.615
R395 VTAIL.n67 VTAIL.n21 104.615
R396 VTAIL.n68 VTAIL.n67 104.615
R397 VTAIL.n68 VTAIL.n17 104.615
R398 VTAIL.n75 VTAIL.n17 104.615
R399 VTAIL.n77 VTAIL.n75 104.615
R400 VTAIL.n77 VTAIL.n76 104.615
R401 VTAIL.n76 VTAIL.n13 104.615
R402 VTAIL.n85 VTAIL.n13 104.615
R403 VTAIL.n86 VTAIL.n85 104.615
R404 VTAIL.n86 VTAIL.n9 104.615
R405 VTAIL.n93 VTAIL.n9 104.615
R406 VTAIL.n94 VTAIL.n93 104.615
R407 VTAIL.n94 VTAIL.n5 104.615
R408 VTAIL.n101 VTAIL.n5 104.615
R409 VTAIL.n102 VTAIL.n101 104.615
R410 VTAIL.n142 VTAIL.n139 104.615
R411 VTAIL.n149 VTAIL.n139 104.615
R412 VTAIL.n150 VTAIL.n149 104.615
R413 VTAIL.n150 VTAIL.n135 104.615
R414 VTAIL.n157 VTAIL.n135 104.615
R415 VTAIL.n158 VTAIL.n157 104.615
R416 VTAIL.n158 VTAIL.n131 104.615
R417 VTAIL.n165 VTAIL.n131 104.615
R418 VTAIL.n166 VTAIL.n165 104.615
R419 VTAIL.n166 VTAIL.n127 104.615
R420 VTAIL.n173 VTAIL.n127 104.615
R421 VTAIL.n174 VTAIL.n173 104.615
R422 VTAIL.n174 VTAIL.n123 104.615
R423 VTAIL.n181 VTAIL.n123 104.615
R424 VTAIL.n183 VTAIL.n181 104.615
R425 VTAIL.n183 VTAIL.n182 104.615
R426 VTAIL.n182 VTAIL.n119 104.615
R427 VTAIL.n191 VTAIL.n119 104.615
R428 VTAIL.n192 VTAIL.n191 104.615
R429 VTAIL.n192 VTAIL.n115 104.615
R430 VTAIL.n199 VTAIL.n115 104.615
R431 VTAIL.n200 VTAIL.n199 104.615
R432 VTAIL.n200 VTAIL.n111 104.615
R433 VTAIL.n207 VTAIL.n111 104.615
R434 VTAIL.n208 VTAIL.n207 104.615
R435 VTAIL.n250 VTAIL.n247 104.615
R436 VTAIL.n257 VTAIL.n247 104.615
R437 VTAIL.n258 VTAIL.n257 104.615
R438 VTAIL.n258 VTAIL.n243 104.615
R439 VTAIL.n265 VTAIL.n243 104.615
R440 VTAIL.n266 VTAIL.n265 104.615
R441 VTAIL.n266 VTAIL.n239 104.615
R442 VTAIL.n273 VTAIL.n239 104.615
R443 VTAIL.n274 VTAIL.n273 104.615
R444 VTAIL.n274 VTAIL.n235 104.615
R445 VTAIL.n281 VTAIL.n235 104.615
R446 VTAIL.n282 VTAIL.n281 104.615
R447 VTAIL.n282 VTAIL.n231 104.615
R448 VTAIL.n289 VTAIL.n231 104.615
R449 VTAIL.n291 VTAIL.n289 104.615
R450 VTAIL.n291 VTAIL.n290 104.615
R451 VTAIL.n290 VTAIL.n227 104.615
R452 VTAIL.n299 VTAIL.n227 104.615
R453 VTAIL.n300 VTAIL.n299 104.615
R454 VTAIL.n300 VTAIL.n223 104.615
R455 VTAIL.n307 VTAIL.n223 104.615
R456 VTAIL.n308 VTAIL.n307 104.615
R457 VTAIL.n308 VTAIL.n219 104.615
R458 VTAIL.n315 VTAIL.n219 104.615
R459 VTAIL.n316 VTAIL.n315 104.615
R460 VTAIL.n744 VTAIL.n743 104.615
R461 VTAIL.n743 VTAIL.n647 104.615
R462 VTAIL.n736 VTAIL.n647 104.615
R463 VTAIL.n736 VTAIL.n735 104.615
R464 VTAIL.n735 VTAIL.n651 104.615
R465 VTAIL.n728 VTAIL.n651 104.615
R466 VTAIL.n728 VTAIL.n727 104.615
R467 VTAIL.n727 VTAIL.n655 104.615
R468 VTAIL.n659 VTAIL.n655 104.615
R469 VTAIL.n719 VTAIL.n659 104.615
R470 VTAIL.n719 VTAIL.n718 104.615
R471 VTAIL.n718 VTAIL.n660 104.615
R472 VTAIL.n711 VTAIL.n660 104.615
R473 VTAIL.n711 VTAIL.n710 104.615
R474 VTAIL.n710 VTAIL.n664 104.615
R475 VTAIL.n703 VTAIL.n664 104.615
R476 VTAIL.n703 VTAIL.n702 104.615
R477 VTAIL.n702 VTAIL.n668 104.615
R478 VTAIL.n695 VTAIL.n668 104.615
R479 VTAIL.n695 VTAIL.n694 104.615
R480 VTAIL.n694 VTAIL.n672 104.615
R481 VTAIL.n687 VTAIL.n672 104.615
R482 VTAIL.n687 VTAIL.n686 104.615
R483 VTAIL.n686 VTAIL.n676 104.615
R484 VTAIL.n679 VTAIL.n676 104.615
R485 VTAIL.n636 VTAIL.n635 104.615
R486 VTAIL.n635 VTAIL.n539 104.615
R487 VTAIL.n628 VTAIL.n539 104.615
R488 VTAIL.n628 VTAIL.n627 104.615
R489 VTAIL.n627 VTAIL.n543 104.615
R490 VTAIL.n620 VTAIL.n543 104.615
R491 VTAIL.n620 VTAIL.n619 104.615
R492 VTAIL.n619 VTAIL.n547 104.615
R493 VTAIL.n551 VTAIL.n547 104.615
R494 VTAIL.n611 VTAIL.n551 104.615
R495 VTAIL.n611 VTAIL.n610 104.615
R496 VTAIL.n610 VTAIL.n552 104.615
R497 VTAIL.n603 VTAIL.n552 104.615
R498 VTAIL.n603 VTAIL.n602 104.615
R499 VTAIL.n602 VTAIL.n556 104.615
R500 VTAIL.n595 VTAIL.n556 104.615
R501 VTAIL.n595 VTAIL.n594 104.615
R502 VTAIL.n594 VTAIL.n560 104.615
R503 VTAIL.n587 VTAIL.n560 104.615
R504 VTAIL.n587 VTAIL.n586 104.615
R505 VTAIL.n586 VTAIL.n564 104.615
R506 VTAIL.n579 VTAIL.n564 104.615
R507 VTAIL.n579 VTAIL.n578 104.615
R508 VTAIL.n578 VTAIL.n568 104.615
R509 VTAIL.n571 VTAIL.n568 104.615
R510 VTAIL.n530 VTAIL.n529 104.615
R511 VTAIL.n529 VTAIL.n433 104.615
R512 VTAIL.n522 VTAIL.n433 104.615
R513 VTAIL.n522 VTAIL.n521 104.615
R514 VTAIL.n521 VTAIL.n437 104.615
R515 VTAIL.n514 VTAIL.n437 104.615
R516 VTAIL.n514 VTAIL.n513 104.615
R517 VTAIL.n513 VTAIL.n441 104.615
R518 VTAIL.n445 VTAIL.n441 104.615
R519 VTAIL.n505 VTAIL.n445 104.615
R520 VTAIL.n505 VTAIL.n504 104.615
R521 VTAIL.n504 VTAIL.n446 104.615
R522 VTAIL.n497 VTAIL.n446 104.615
R523 VTAIL.n497 VTAIL.n496 104.615
R524 VTAIL.n496 VTAIL.n450 104.615
R525 VTAIL.n489 VTAIL.n450 104.615
R526 VTAIL.n489 VTAIL.n488 104.615
R527 VTAIL.n488 VTAIL.n454 104.615
R528 VTAIL.n481 VTAIL.n454 104.615
R529 VTAIL.n481 VTAIL.n480 104.615
R530 VTAIL.n480 VTAIL.n458 104.615
R531 VTAIL.n473 VTAIL.n458 104.615
R532 VTAIL.n473 VTAIL.n472 104.615
R533 VTAIL.n472 VTAIL.n462 104.615
R534 VTAIL.n465 VTAIL.n462 104.615
R535 VTAIL.n422 VTAIL.n421 104.615
R536 VTAIL.n421 VTAIL.n325 104.615
R537 VTAIL.n414 VTAIL.n325 104.615
R538 VTAIL.n414 VTAIL.n413 104.615
R539 VTAIL.n413 VTAIL.n329 104.615
R540 VTAIL.n406 VTAIL.n329 104.615
R541 VTAIL.n406 VTAIL.n405 104.615
R542 VTAIL.n405 VTAIL.n333 104.615
R543 VTAIL.n337 VTAIL.n333 104.615
R544 VTAIL.n397 VTAIL.n337 104.615
R545 VTAIL.n397 VTAIL.n396 104.615
R546 VTAIL.n396 VTAIL.n338 104.615
R547 VTAIL.n389 VTAIL.n338 104.615
R548 VTAIL.n389 VTAIL.n388 104.615
R549 VTAIL.n388 VTAIL.n342 104.615
R550 VTAIL.n381 VTAIL.n342 104.615
R551 VTAIL.n381 VTAIL.n380 104.615
R552 VTAIL.n380 VTAIL.n346 104.615
R553 VTAIL.n373 VTAIL.n346 104.615
R554 VTAIL.n373 VTAIL.n372 104.615
R555 VTAIL.n372 VTAIL.n350 104.615
R556 VTAIL.n365 VTAIL.n350 104.615
R557 VTAIL.n365 VTAIL.n364 104.615
R558 VTAIL.n364 VTAIL.n354 104.615
R559 VTAIL.n357 VTAIL.n354 104.615
R560 VTAIL.n784 VTAIL.t5 52.3082
R561 VTAIL.n36 VTAIL.t9 52.3082
R562 VTAIL.n142 VTAIL.t11 52.3082
R563 VTAIL.n250 VTAIL.t13 52.3082
R564 VTAIL.n679 VTAIL.t12 52.3082
R565 VTAIL.n571 VTAIL.t14 52.3082
R566 VTAIL.n465 VTAIL.t7 52.3082
R567 VTAIL.n357 VTAIL.t6 52.3082
R568 VTAIL.n1 VTAIL.n0 42.3917
R569 VTAIL.n215 VTAIL.n214 42.3917
R570 VTAIL.n643 VTAIL.n642 42.3917
R571 VTAIL.n429 VTAIL.n428 42.3917
R572 VTAIL.n855 VTAIL.n749 32.2979
R573 VTAIL.n427 VTAIL.n321 32.2979
R574 VTAIL.n855 VTAIL.n854 30.6338
R575 VTAIL.n107 VTAIL.n106 30.6338
R576 VTAIL.n213 VTAIL.n212 30.6338
R577 VTAIL.n321 VTAIL.n320 30.6338
R578 VTAIL.n749 VTAIL.n748 30.6338
R579 VTAIL.n641 VTAIL.n640 30.6338
R580 VTAIL.n535 VTAIL.n534 30.6338
R581 VTAIL.n427 VTAIL.n426 30.6338
R582 VTAIL.n785 VTAIL.n783 15.6677
R583 VTAIL.n37 VTAIL.n35 15.6677
R584 VTAIL.n143 VTAIL.n141 15.6677
R585 VTAIL.n251 VTAIL.n249 15.6677
R586 VTAIL.n680 VTAIL.n678 15.6677
R587 VTAIL.n572 VTAIL.n570 15.6677
R588 VTAIL.n466 VTAIL.n464 15.6677
R589 VTAIL.n358 VTAIL.n356 15.6677
R590 VTAIL.n832 VTAIL.n831 13.1884
R591 VTAIL.n84 VTAIL.n83 13.1884
R592 VTAIL.n190 VTAIL.n189 13.1884
R593 VTAIL.n298 VTAIL.n297 13.1884
R594 VTAIL.n726 VTAIL.n725 13.1884
R595 VTAIL.n618 VTAIL.n617 13.1884
R596 VTAIL.n512 VTAIL.n511 13.1884
R597 VTAIL.n404 VTAIL.n403 13.1884
R598 VTAIL.n786 VTAIL.n782 12.8005
R599 VTAIL.n830 VTAIL.n762 12.8005
R600 VTAIL.n835 VTAIL.n760 12.8005
R601 VTAIL.n38 VTAIL.n34 12.8005
R602 VTAIL.n82 VTAIL.n14 12.8005
R603 VTAIL.n87 VTAIL.n12 12.8005
R604 VTAIL.n144 VTAIL.n140 12.8005
R605 VTAIL.n188 VTAIL.n120 12.8005
R606 VTAIL.n193 VTAIL.n118 12.8005
R607 VTAIL.n252 VTAIL.n248 12.8005
R608 VTAIL.n296 VTAIL.n228 12.8005
R609 VTAIL.n301 VTAIL.n226 12.8005
R610 VTAIL.n729 VTAIL.n654 12.8005
R611 VTAIL.n724 VTAIL.n656 12.8005
R612 VTAIL.n681 VTAIL.n677 12.8005
R613 VTAIL.n621 VTAIL.n546 12.8005
R614 VTAIL.n616 VTAIL.n548 12.8005
R615 VTAIL.n573 VTAIL.n569 12.8005
R616 VTAIL.n515 VTAIL.n440 12.8005
R617 VTAIL.n510 VTAIL.n442 12.8005
R618 VTAIL.n467 VTAIL.n463 12.8005
R619 VTAIL.n407 VTAIL.n332 12.8005
R620 VTAIL.n402 VTAIL.n334 12.8005
R621 VTAIL.n359 VTAIL.n355 12.8005
R622 VTAIL.n790 VTAIL.n789 12.0247
R623 VTAIL.n827 VTAIL.n826 12.0247
R624 VTAIL.n836 VTAIL.n758 12.0247
R625 VTAIL.n42 VTAIL.n41 12.0247
R626 VTAIL.n79 VTAIL.n78 12.0247
R627 VTAIL.n88 VTAIL.n10 12.0247
R628 VTAIL.n148 VTAIL.n147 12.0247
R629 VTAIL.n185 VTAIL.n184 12.0247
R630 VTAIL.n194 VTAIL.n116 12.0247
R631 VTAIL.n256 VTAIL.n255 12.0247
R632 VTAIL.n293 VTAIL.n292 12.0247
R633 VTAIL.n302 VTAIL.n224 12.0247
R634 VTAIL.n730 VTAIL.n652 12.0247
R635 VTAIL.n721 VTAIL.n720 12.0247
R636 VTAIL.n685 VTAIL.n684 12.0247
R637 VTAIL.n622 VTAIL.n544 12.0247
R638 VTAIL.n613 VTAIL.n612 12.0247
R639 VTAIL.n577 VTAIL.n576 12.0247
R640 VTAIL.n516 VTAIL.n438 12.0247
R641 VTAIL.n507 VTAIL.n506 12.0247
R642 VTAIL.n471 VTAIL.n470 12.0247
R643 VTAIL.n408 VTAIL.n330 12.0247
R644 VTAIL.n399 VTAIL.n398 12.0247
R645 VTAIL.n363 VTAIL.n362 12.0247
R646 VTAIL.n793 VTAIL.n780 11.249
R647 VTAIL.n822 VTAIL.n764 11.249
R648 VTAIL.n840 VTAIL.n839 11.249
R649 VTAIL.n45 VTAIL.n32 11.249
R650 VTAIL.n74 VTAIL.n16 11.249
R651 VTAIL.n92 VTAIL.n91 11.249
R652 VTAIL.n151 VTAIL.n138 11.249
R653 VTAIL.n180 VTAIL.n122 11.249
R654 VTAIL.n198 VTAIL.n197 11.249
R655 VTAIL.n259 VTAIL.n246 11.249
R656 VTAIL.n288 VTAIL.n230 11.249
R657 VTAIL.n306 VTAIL.n305 11.249
R658 VTAIL.n734 VTAIL.n733 11.249
R659 VTAIL.n717 VTAIL.n658 11.249
R660 VTAIL.n688 VTAIL.n675 11.249
R661 VTAIL.n626 VTAIL.n625 11.249
R662 VTAIL.n609 VTAIL.n550 11.249
R663 VTAIL.n580 VTAIL.n567 11.249
R664 VTAIL.n520 VTAIL.n519 11.249
R665 VTAIL.n503 VTAIL.n444 11.249
R666 VTAIL.n474 VTAIL.n461 11.249
R667 VTAIL.n412 VTAIL.n411 11.249
R668 VTAIL.n395 VTAIL.n336 11.249
R669 VTAIL.n366 VTAIL.n353 11.249
R670 VTAIL.n794 VTAIL.n778 10.4732
R671 VTAIL.n821 VTAIL.n766 10.4732
R672 VTAIL.n843 VTAIL.n756 10.4732
R673 VTAIL.n46 VTAIL.n30 10.4732
R674 VTAIL.n73 VTAIL.n18 10.4732
R675 VTAIL.n95 VTAIL.n8 10.4732
R676 VTAIL.n152 VTAIL.n136 10.4732
R677 VTAIL.n179 VTAIL.n124 10.4732
R678 VTAIL.n201 VTAIL.n114 10.4732
R679 VTAIL.n260 VTAIL.n244 10.4732
R680 VTAIL.n287 VTAIL.n232 10.4732
R681 VTAIL.n309 VTAIL.n222 10.4732
R682 VTAIL.n737 VTAIL.n650 10.4732
R683 VTAIL.n716 VTAIL.n661 10.4732
R684 VTAIL.n689 VTAIL.n673 10.4732
R685 VTAIL.n629 VTAIL.n542 10.4732
R686 VTAIL.n608 VTAIL.n553 10.4732
R687 VTAIL.n581 VTAIL.n565 10.4732
R688 VTAIL.n523 VTAIL.n436 10.4732
R689 VTAIL.n502 VTAIL.n447 10.4732
R690 VTAIL.n475 VTAIL.n459 10.4732
R691 VTAIL.n415 VTAIL.n328 10.4732
R692 VTAIL.n394 VTAIL.n339 10.4732
R693 VTAIL.n367 VTAIL.n351 10.4732
R694 VTAIL.n798 VTAIL.n797 9.69747
R695 VTAIL.n818 VTAIL.n817 9.69747
R696 VTAIL.n844 VTAIL.n754 9.69747
R697 VTAIL.n50 VTAIL.n49 9.69747
R698 VTAIL.n70 VTAIL.n69 9.69747
R699 VTAIL.n96 VTAIL.n6 9.69747
R700 VTAIL.n156 VTAIL.n155 9.69747
R701 VTAIL.n176 VTAIL.n175 9.69747
R702 VTAIL.n202 VTAIL.n112 9.69747
R703 VTAIL.n264 VTAIL.n263 9.69747
R704 VTAIL.n284 VTAIL.n283 9.69747
R705 VTAIL.n310 VTAIL.n220 9.69747
R706 VTAIL.n738 VTAIL.n648 9.69747
R707 VTAIL.n713 VTAIL.n712 9.69747
R708 VTAIL.n693 VTAIL.n692 9.69747
R709 VTAIL.n630 VTAIL.n540 9.69747
R710 VTAIL.n605 VTAIL.n604 9.69747
R711 VTAIL.n585 VTAIL.n584 9.69747
R712 VTAIL.n524 VTAIL.n434 9.69747
R713 VTAIL.n499 VTAIL.n498 9.69747
R714 VTAIL.n479 VTAIL.n478 9.69747
R715 VTAIL.n416 VTAIL.n326 9.69747
R716 VTAIL.n391 VTAIL.n390 9.69747
R717 VTAIL.n371 VTAIL.n370 9.69747
R718 VTAIL.n854 VTAIL.n853 9.45567
R719 VTAIL.n106 VTAIL.n105 9.45567
R720 VTAIL.n212 VTAIL.n211 9.45567
R721 VTAIL.n320 VTAIL.n319 9.45567
R722 VTAIL.n748 VTAIL.n747 9.45567
R723 VTAIL.n640 VTAIL.n639 9.45567
R724 VTAIL.n534 VTAIL.n533 9.45567
R725 VTAIL.n426 VTAIL.n425 9.45567
R726 VTAIL.n752 VTAIL.n751 9.3005
R727 VTAIL.n847 VTAIL.n846 9.3005
R728 VTAIL.n845 VTAIL.n844 9.3005
R729 VTAIL.n756 VTAIL.n755 9.3005
R730 VTAIL.n839 VTAIL.n838 9.3005
R731 VTAIL.n837 VTAIL.n836 9.3005
R732 VTAIL.n760 VTAIL.n759 9.3005
R733 VTAIL.n805 VTAIL.n804 9.3005
R734 VTAIL.n803 VTAIL.n802 9.3005
R735 VTAIL.n776 VTAIL.n775 9.3005
R736 VTAIL.n797 VTAIL.n796 9.3005
R737 VTAIL.n795 VTAIL.n794 9.3005
R738 VTAIL.n780 VTAIL.n779 9.3005
R739 VTAIL.n789 VTAIL.n788 9.3005
R740 VTAIL.n787 VTAIL.n786 9.3005
R741 VTAIL.n772 VTAIL.n771 9.3005
R742 VTAIL.n811 VTAIL.n810 9.3005
R743 VTAIL.n813 VTAIL.n812 9.3005
R744 VTAIL.n768 VTAIL.n767 9.3005
R745 VTAIL.n819 VTAIL.n818 9.3005
R746 VTAIL.n821 VTAIL.n820 9.3005
R747 VTAIL.n764 VTAIL.n763 9.3005
R748 VTAIL.n828 VTAIL.n827 9.3005
R749 VTAIL.n830 VTAIL.n829 9.3005
R750 VTAIL.n853 VTAIL.n852 9.3005
R751 VTAIL.n4 VTAIL.n3 9.3005
R752 VTAIL.n99 VTAIL.n98 9.3005
R753 VTAIL.n97 VTAIL.n96 9.3005
R754 VTAIL.n8 VTAIL.n7 9.3005
R755 VTAIL.n91 VTAIL.n90 9.3005
R756 VTAIL.n89 VTAIL.n88 9.3005
R757 VTAIL.n12 VTAIL.n11 9.3005
R758 VTAIL.n57 VTAIL.n56 9.3005
R759 VTAIL.n55 VTAIL.n54 9.3005
R760 VTAIL.n28 VTAIL.n27 9.3005
R761 VTAIL.n49 VTAIL.n48 9.3005
R762 VTAIL.n47 VTAIL.n46 9.3005
R763 VTAIL.n32 VTAIL.n31 9.3005
R764 VTAIL.n41 VTAIL.n40 9.3005
R765 VTAIL.n39 VTAIL.n38 9.3005
R766 VTAIL.n24 VTAIL.n23 9.3005
R767 VTAIL.n63 VTAIL.n62 9.3005
R768 VTAIL.n65 VTAIL.n64 9.3005
R769 VTAIL.n20 VTAIL.n19 9.3005
R770 VTAIL.n71 VTAIL.n70 9.3005
R771 VTAIL.n73 VTAIL.n72 9.3005
R772 VTAIL.n16 VTAIL.n15 9.3005
R773 VTAIL.n80 VTAIL.n79 9.3005
R774 VTAIL.n82 VTAIL.n81 9.3005
R775 VTAIL.n105 VTAIL.n104 9.3005
R776 VTAIL.n110 VTAIL.n109 9.3005
R777 VTAIL.n205 VTAIL.n204 9.3005
R778 VTAIL.n203 VTAIL.n202 9.3005
R779 VTAIL.n114 VTAIL.n113 9.3005
R780 VTAIL.n197 VTAIL.n196 9.3005
R781 VTAIL.n195 VTAIL.n194 9.3005
R782 VTAIL.n118 VTAIL.n117 9.3005
R783 VTAIL.n163 VTAIL.n162 9.3005
R784 VTAIL.n161 VTAIL.n160 9.3005
R785 VTAIL.n134 VTAIL.n133 9.3005
R786 VTAIL.n155 VTAIL.n154 9.3005
R787 VTAIL.n153 VTAIL.n152 9.3005
R788 VTAIL.n138 VTAIL.n137 9.3005
R789 VTAIL.n147 VTAIL.n146 9.3005
R790 VTAIL.n145 VTAIL.n144 9.3005
R791 VTAIL.n130 VTAIL.n129 9.3005
R792 VTAIL.n169 VTAIL.n168 9.3005
R793 VTAIL.n171 VTAIL.n170 9.3005
R794 VTAIL.n126 VTAIL.n125 9.3005
R795 VTAIL.n177 VTAIL.n176 9.3005
R796 VTAIL.n179 VTAIL.n178 9.3005
R797 VTAIL.n122 VTAIL.n121 9.3005
R798 VTAIL.n186 VTAIL.n185 9.3005
R799 VTAIL.n188 VTAIL.n187 9.3005
R800 VTAIL.n211 VTAIL.n210 9.3005
R801 VTAIL.n218 VTAIL.n217 9.3005
R802 VTAIL.n313 VTAIL.n312 9.3005
R803 VTAIL.n311 VTAIL.n310 9.3005
R804 VTAIL.n222 VTAIL.n221 9.3005
R805 VTAIL.n305 VTAIL.n304 9.3005
R806 VTAIL.n303 VTAIL.n302 9.3005
R807 VTAIL.n226 VTAIL.n225 9.3005
R808 VTAIL.n271 VTAIL.n270 9.3005
R809 VTAIL.n269 VTAIL.n268 9.3005
R810 VTAIL.n242 VTAIL.n241 9.3005
R811 VTAIL.n263 VTAIL.n262 9.3005
R812 VTAIL.n261 VTAIL.n260 9.3005
R813 VTAIL.n246 VTAIL.n245 9.3005
R814 VTAIL.n255 VTAIL.n254 9.3005
R815 VTAIL.n253 VTAIL.n252 9.3005
R816 VTAIL.n238 VTAIL.n237 9.3005
R817 VTAIL.n277 VTAIL.n276 9.3005
R818 VTAIL.n279 VTAIL.n278 9.3005
R819 VTAIL.n234 VTAIL.n233 9.3005
R820 VTAIL.n285 VTAIL.n284 9.3005
R821 VTAIL.n287 VTAIL.n286 9.3005
R822 VTAIL.n230 VTAIL.n229 9.3005
R823 VTAIL.n294 VTAIL.n293 9.3005
R824 VTAIL.n296 VTAIL.n295 9.3005
R825 VTAIL.n319 VTAIL.n318 9.3005
R826 VTAIL.n706 VTAIL.n705 9.3005
R827 VTAIL.n708 VTAIL.n707 9.3005
R828 VTAIL.n663 VTAIL.n662 9.3005
R829 VTAIL.n714 VTAIL.n713 9.3005
R830 VTAIL.n716 VTAIL.n715 9.3005
R831 VTAIL.n658 VTAIL.n657 9.3005
R832 VTAIL.n722 VTAIL.n721 9.3005
R833 VTAIL.n724 VTAIL.n723 9.3005
R834 VTAIL.n747 VTAIL.n746 9.3005
R835 VTAIL.n646 VTAIL.n645 9.3005
R836 VTAIL.n741 VTAIL.n740 9.3005
R837 VTAIL.n739 VTAIL.n738 9.3005
R838 VTAIL.n650 VTAIL.n649 9.3005
R839 VTAIL.n733 VTAIL.n732 9.3005
R840 VTAIL.n731 VTAIL.n730 9.3005
R841 VTAIL.n654 VTAIL.n653 9.3005
R842 VTAIL.n667 VTAIL.n666 9.3005
R843 VTAIL.n700 VTAIL.n699 9.3005
R844 VTAIL.n698 VTAIL.n697 9.3005
R845 VTAIL.n671 VTAIL.n670 9.3005
R846 VTAIL.n692 VTAIL.n691 9.3005
R847 VTAIL.n690 VTAIL.n689 9.3005
R848 VTAIL.n675 VTAIL.n674 9.3005
R849 VTAIL.n684 VTAIL.n683 9.3005
R850 VTAIL.n682 VTAIL.n681 9.3005
R851 VTAIL.n598 VTAIL.n597 9.3005
R852 VTAIL.n600 VTAIL.n599 9.3005
R853 VTAIL.n555 VTAIL.n554 9.3005
R854 VTAIL.n606 VTAIL.n605 9.3005
R855 VTAIL.n608 VTAIL.n607 9.3005
R856 VTAIL.n550 VTAIL.n549 9.3005
R857 VTAIL.n614 VTAIL.n613 9.3005
R858 VTAIL.n616 VTAIL.n615 9.3005
R859 VTAIL.n639 VTAIL.n638 9.3005
R860 VTAIL.n538 VTAIL.n537 9.3005
R861 VTAIL.n633 VTAIL.n632 9.3005
R862 VTAIL.n631 VTAIL.n630 9.3005
R863 VTAIL.n542 VTAIL.n541 9.3005
R864 VTAIL.n625 VTAIL.n624 9.3005
R865 VTAIL.n623 VTAIL.n622 9.3005
R866 VTAIL.n546 VTAIL.n545 9.3005
R867 VTAIL.n559 VTAIL.n558 9.3005
R868 VTAIL.n592 VTAIL.n591 9.3005
R869 VTAIL.n590 VTAIL.n589 9.3005
R870 VTAIL.n563 VTAIL.n562 9.3005
R871 VTAIL.n584 VTAIL.n583 9.3005
R872 VTAIL.n582 VTAIL.n581 9.3005
R873 VTAIL.n567 VTAIL.n566 9.3005
R874 VTAIL.n576 VTAIL.n575 9.3005
R875 VTAIL.n574 VTAIL.n573 9.3005
R876 VTAIL.n492 VTAIL.n491 9.3005
R877 VTAIL.n494 VTAIL.n493 9.3005
R878 VTAIL.n449 VTAIL.n448 9.3005
R879 VTAIL.n500 VTAIL.n499 9.3005
R880 VTAIL.n502 VTAIL.n501 9.3005
R881 VTAIL.n444 VTAIL.n443 9.3005
R882 VTAIL.n508 VTAIL.n507 9.3005
R883 VTAIL.n510 VTAIL.n509 9.3005
R884 VTAIL.n533 VTAIL.n532 9.3005
R885 VTAIL.n432 VTAIL.n431 9.3005
R886 VTAIL.n527 VTAIL.n526 9.3005
R887 VTAIL.n525 VTAIL.n524 9.3005
R888 VTAIL.n436 VTAIL.n435 9.3005
R889 VTAIL.n519 VTAIL.n518 9.3005
R890 VTAIL.n517 VTAIL.n516 9.3005
R891 VTAIL.n440 VTAIL.n439 9.3005
R892 VTAIL.n453 VTAIL.n452 9.3005
R893 VTAIL.n486 VTAIL.n485 9.3005
R894 VTAIL.n484 VTAIL.n483 9.3005
R895 VTAIL.n457 VTAIL.n456 9.3005
R896 VTAIL.n478 VTAIL.n477 9.3005
R897 VTAIL.n476 VTAIL.n475 9.3005
R898 VTAIL.n461 VTAIL.n460 9.3005
R899 VTAIL.n470 VTAIL.n469 9.3005
R900 VTAIL.n468 VTAIL.n467 9.3005
R901 VTAIL.n384 VTAIL.n383 9.3005
R902 VTAIL.n386 VTAIL.n385 9.3005
R903 VTAIL.n341 VTAIL.n340 9.3005
R904 VTAIL.n392 VTAIL.n391 9.3005
R905 VTAIL.n394 VTAIL.n393 9.3005
R906 VTAIL.n336 VTAIL.n335 9.3005
R907 VTAIL.n400 VTAIL.n399 9.3005
R908 VTAIL.n402 VTAIL.n401 9.3005
R909 VTAIL.n425 VTAIL.n424 9.3005
R910 VTAIL.n324 VTAIL.n323 9.3005
R911 VTAIL.n419 VTAIL.n418 9.3005
R912 VTAIL.n417 VTAIL.n416 9.3005
R913 VTAIL.n328 VTAIL.n327 9.3005
R914 VTAIL.n411 VTAIL.n410 9.3005
R915 VTAIL.n409 VTAIL.n408 9.3005
R916 VTAIL.n332 VTAIL.n331 9.3005
R917 VTAIL.n345 VTAIL.n344 9.3005
R918 VTAIL.n378 VTAIL.n377 9.3005
R919 VTAIL.n376 VTAIL.n375 9.3005
R920 VTAIL.n349 VTAIL.n348 9.3005
R921 VTAIL.n370 VTAIL.n369 9.3005
R922 VTAIL.n368 VTAIL.n367 9.3005
R923 VTAIL.n353 VTAIL.n352 9.3005
R924 VTAIL.n362 VTAIL.n361 9.3005
R925 VTAIL.n360 VTAIL.n359 9.3005
R926 VTAIL.n801 VTAIL.n776 8.92171
R927 VTAIL.n814 VTAIL.n768 8.92171
R928 VTAIL.n848 VTAIL.n847 8.92171
R929 VTAIL.n53 VTAIL.n28 8.92171
R930 VTAIL.n66 VTAIL.n20 8.92171
R931 VTAIL.n100 VTAIL.n99 8.92171
R932 VTAIL.n159 VTAIL.n134 8.92171
R933 VTAIL.n172 VTAIL.n126 8.92171
R934 VTAIL.n206 VTAIL.n205 8.92171
R935 VTAIL.n267 VTAIL.n242 8.92171
R936 VTAIL.n280 VTAIL.n234 8.92171
R937 VTAIL.n314 VTAIL.n313 8.92171
R938 VTAIL.n742 VTAIL.n741 8.92171
R939 VTAIL.n709 VTAIL.n663 8.92171
R940 VTAIL.n696 VTAIL.n671 8.92171
R941 VTAIL.n634 VTAIL.n633 8.92171
R942 VTAIL.n601 VTAIL.n555 8.92171
R943 VTAIL.n588 VTAIL.n563 8.92171
R944 VTAIL.n528 VTAIL.n527 8.92171
R945 VTAIL.n495 VTAIL.n449 8.92171
R946 VTAIL.n482 VTAIL.n457 8.92171
R947 VTAIL.n420 VTAIL.n419 8.92171
R948 VTAIL.n387 VTAIL.n341 8.92171
R949 VTAIL.n374 VTAIL.n349 8.92171
R950 VTAIL.n802 VTAIL.n774 8.14595
R951 VTAIL.n813 VTAIL.n770 8.14595
R952 VTAIL.n851 VTAIL.n752 8.14595
R953 VTAIL.n54 VTAIL.n26 8.14595
R954 VTAIL.n65 VTAIL.n22 8.14595
R955 VTAIL.n103 VTAIL.n4 8.14595
R956 VTAIL.n160 VTAIL.n132 8.14595
R957 VTAIL.n171 VTAIL.n128 8.14595
R958 VTAIL.n209 VTAIL.n110 8.14595
R959 VTAIL.n268 VTAIL.n240 8.14595
R960 VTAIL.n279 VTAIL.n236 8.14595
R961 VTAIL.n317 VTAIL.n218 8.14595
R962 VTAIL.n745 VTAIL.n646 8.14595
R963 VTAIL.n708 VTAIL.n665 8.14595
R964 VTAIL.n697 VTAIL.n669 8.14595
R965 VTAIL.n637 VTAIL.n538 8.14595
R966 VTAIL.n600 VTAIL.n557 8.14595
R967 VTAIL.n589 VTAIL.n561 8.14595
R968 VTAIL.n531 VTAIL.n432 8.14595
R969 VTAIL.n494 VTAIL.n451 8.14595
R970 VTAIL.n483 VTAIL.n455 8.14595
R971 VTAIL.n423 VTAIL.n324 8.14595
R972 VTAIL.n386 VTAIL.n343 8.14595
R973 VTAIL.n375 VTAIL.n347 8.14595
R974 VTAIL.n806 VTAIL.n805 7.3702
R975 VTAIL.n810 VTAIL.n809 7.3702
R976 VTAIL.n852 VTAIL.n750 7.3702
R977 VTAIL.n58 VTAIL.n57 7.3702
R978 VTAIL.n62 VTAIL.n61 7.3702
R979 VTAIL.n104 VTAIL.n2 7.3702
R980 VTAIL.n164 VTAIL.n163 7.3702
R981 VTAIL.n168 VTAIL.n167 7.3702
R982 VTAIL.n210 VTAIL.n108 7.3702
R983 VTAIL.n272 VTAIL.n271 7.3702
R984 VTAIL.n276 VTAIL.n275 7.3702
R985 VTAIL.n318 VTAIL.n216 7.3702
R986 VTAIL.n746 VTAIL.n644 7.3702
R987 VTAIL.n705 VTAIL.n704 7.3702
R988 VTAIL.n701 VTAIL.n700 7.3702
R989 VTAIL.n638 VTAIL.n536 7.3702
R990 VTAIL.n597 VTAIL.n596 7.3702
R991 VTAIL.n593 VTAIL.n592 7.3702
R992 VTAIL.n532 VTAIL.n430 7.3702
R993 VTAIL.n491 VTAIL.n490 7.3702
R994 VTAIL.n487 VTAIL.n486 7.3702
R995 VTAIL.n424 VTAIL.n322 7.3702
R996 VTAIL.n383 VTAIL.n382 7.3702
R997 VTAIL.n379 VTAIL.n378 7.3702
R998 VTAIL.n806 VTAIL.n772 6.59444
R999 VTAIL.n809 VTAIL.n772 6.59444
R1000 VTAIL.n854 VTAIL.n750 6.59444
R1001 VTAIL.n58 VTAIL.n24 6.59444
R1002 VTAIL.n61 VTAIL.n24 6.59444
R1003 VTAIL.n106 VTAIL.n2 6.59444
R1004 VTAIL.n164 VTAIL.n130 6.59444
R1005 VTAIL.n167 VTAIL.n130 6.59444
R1006 VTAIL.n212 VTAIL.n108 6.59444
R1007 VTAIL.n272 VTAIL.n238 6.59444
R1008 VTAIL.n275 VTAIL.n238 6.59444
R1009 VTAIL.n320 VTAIL.n216 6.59444
R1010 VTAIL.n748 VTAIL.n644 6.59444
R1011 VTAIL.n704 VTAIL.n667 6.59444
R1012 VTAIL.n701 VTAIL.n667 6.59444
R1013 VTAIL.n640 VTAIL.n536 6.59444
R1014 VTAIL.n596 VTAIL.n559 6.59444
R1015 VTAIL.n593 VTAIL.n559 6.59444
R1016 VTAIL.n534 VTAIL.n430 6.59444
R1017 VTAIL.n490 VTAIL.n453 6.59444
R1018 VTAIL.n487 VTAIL.n453 6.59444
R1019 VTAIL.n426 VTAIL.n322 6.59444
R1020 VTAIL.n382 VTAIL.n345 6.59444
R1021 VTAIL.n379 VTAIL.n345 6.59444
R1022 VTAIL.n805 VTAIL.n774 5.81868
R1023 VTAIL.n810 VTAIL.n770 5.81868
R1024 VTAIL.n852 VTAIL.n851 5.81868
R1025 VTAIL.n57 VTAIL.n26 5.81868
R1026 VTAIL.n62 VTAIL.n22 5.81868
R1027 VTAIL.n104 VTAIL.n103 5.81868
R1028 VTAIL.n163 VTAIL.n132 5.81868
R1029 VTAIL.n168 VTAIL.n128 5.81868
R1030 VTAIL.n210 VTAIL.n209 5.81868
R1031 VTAIL.n271 VTAIL.n240 5.81868
R1032 VTAIL.n276 VTAIL.n236 5.81868
R1033 VTAIL.n318 VTAIL.n317 5.81868
R1034 VTAIL.n746 VTAIL.n745 5.81868
R1035 VTAIL.n705 VTAIL.n665 5.81868
R1036 VTAIL.n700 VTAIL.n669 5.81868
R1037 VTAIL.n638 VTAIL.n637 5.81868
R1038 VTAIL.n597 VTAIL.n557 5.81868
R1039 VTAIL.n592 VTAIL.n561 5.81868
R1040 VTAIL.n532 VTAIL.n531 5.81868
R1041 VTAIL.n491 VTAIL.n451 5.81868
R1042 VTAIL.n486 VTAIL.n455 5.81868
R1043 VTAIL.n424 VTAIL.n423 5.81868
R1044 VTAIL.n383 VTAIL.n343 5.81868
R1045 VTAIL.n378 VTAIL.n347 5.81868
R1046 VTAIL.n802 VTAIL.n801 5.04292
R1047 VTAIL.n814 VTAIL.n813 5.04292
R1048 VTAIL.n848 VTAIL.n752 5.04292
R1049 VTAIL.n54 VTAIL.n53 5.04292
R1050 VTAIL.n66 VTAIL.n65 5.04292
R1051 VTAIL.n100 VTAIL.n4 5.04292
R1052 VTAIL.n160 VTAIL.n159 5.04292
R1053 VTAIL.n172 VTAIL.n171 5.04292
R1054 VTAIL.n206 VTAIL.n110 5.04292
R1055 VTAIL.n268 VTAIL.n267 5.04292
R1056 VTAIL.n280 VTAIL.n279 5.04292
R1057 VTAIL.n314 VTAIL.n218 5.04292
R1058 VTAIL.n742 VTAIL.n646 5.04292
R1059 VTAIL.n709 VTAIL.n708 5.04292
R1060 VTAIL.n697 VTAIL.n696 5.04292
R1061 VTAIL.n634 VTAIL.n538 5.04292
R1062 VTAIL.n601 VTAIL.n600 5.04292
R1063 VTAIL.n589 VTAIL.n588 5.04292
R1064 VTAIL.n528 VTAIL.n432 5.04292
R1065 VTAIL.n495 VTAIL.n494 5.04292
R1066 VTAIL.n483 VTAIL.n482 5.04292
R1067 VTAIL.n420 VTAIL.n324 5.04292
R1068 VTAIL.n387 VTAIL.n386 5.04292
R1069 VTAIL.n375 VTAIL.n374 5.04292
R1070 VTAIL.n682 VTAIL.n678 4.38563
R1071 VTAIL.n574 VTAIL.n570 4.38563
R1072 VTAIL.n468 VTAIL.n464 4.38563
R1073 VTAIL.n360 VTAIL.n356 4.38563
R1074 VTAIL.n787 VTAIL.n783 4.38563
R1075 VTAIL.n39 VTAIL.n35 4.38563
R1076 VTAIL.n145 VTAIL.n141 4.38563
R1077 VTAIL.n253 VTAIL.n249 4.38563
R1078 VTAIL.n798 VTAIL.n776 4.26717
R1079 VTAIL.n817 VTAIL.n768 4.26717
R1080 VTAIL.n847 VTAIL.n754 4.26717
R1081 VTAIL.n50 VTAIL.n28 4.26717
R1082 VTAIL.n69 VTAIL.n20 4.26717
R1083 VTAIL.n99 VTAIL.n6 4.26717
R1084 VTAIL.n156 VTAIL.n134 4.26717
R1085 VTAIL.n175 VTAIL.n126 4.26717
R1086 VTAIL.n205 VTAIL.n112 4.26717
R1087 VTAIL.n264 VTAIL.n242 4.26717
R1088 VTAIL.n283 VTAIL.n234 4.26717
R1089 VTAIL.n313 VTAIL.n220 4.26717
R1090 VTAIL.n741 VTAIL.n648 4.26717
R1091 VTAIL.n712 VTAIL.n663 4.26717
R1092 VTAIL.n693 VTAIL.n671 4.26717
R1093 VTAIL.n633 VTAIL.n540 4.26717
R1094 VTAIL.n604 VTAIL.n555 4.26717
R1095 VTAIL.n585 VTAIL.n563 4.26717
R1096 VTAIL.n527 VTAIL.n434 4.26717
R1097 VTAIL.n498 VTAIL.n449 4.26717
R1098 VTAIL.n479 VTAIL.n457 4.26717
R1099 VTAIL.n419 VTAIL.n326 4.26717
R1100 VTAIL.n390 VTAIL.n341 4.26717
R1101 VTAIL.n371 VTAIL.n349 4.26717
R1102 VTAIL.n429 VTAIL.n427 3.65567
R1103 VTAIL.n535 VTAIL.n429 3.65567
R1104 VTAIL.n643 VTAIL.n641 3.65567
R1105 VTAIL.n749 VTAIL.n643 3.65567
R1106 VTAIL.n321 VTAIL.n215 3.65567
R1107 VTAIL.n215 VTAIL.n213 3.65567
R1108 VTAIL.n107 VTAIL.n1 3.65567
R1109 VTAIL VTAIL.n855 3.59748
R1110 VTAIL.n797 VTAIL.n778 3.49141
R1111 VTAIL.n818 VTAIL.n766 3.49141
R1112 VTAIL.n844 VTAIL.n843 3.49141
R1113 VTAIL.n49 VTAIL.n30 3.49141
R1114 VTAIL.n70 VTAIL.n18 3.49141
R1115 VTAIL.n96 VTAIL.n95 3.49141
R1116 VTAIL.n155 VTAIL.n136 3.49141
R1117 VTAIL.n176 VTAIL.n124 3.49141
R1118 VTAIL.n202 VTAIL.n201 3.49141
R1119 VTAIL.n263 VTAIL.n244 3.49141
R1120 VTAIL.n284 VTAIL.n232 3.49141
R1121 VTAIL.n310 VTAIL.n309 3.49141
R1122 VTAIL.n738 VTAIL.n737 3.49141
R1123 VTAIL.n713 VTAIL.n661 3.49141
R1124 VTAIL.n692 VTAIL.n673 3.49141
R1125 VTAIL.n630 VTAIL.n629 3.49141
R1126 VTAIL.n605 VTAIL.n553 3.49141
R1127 VTAIL.n584 VTAIL.n565 3.49141
R1128 VTAIL.n524 VTAIL.n523 3.49141
R1129 VTAIL.n499 VTAIL.n447 3.49141
R1130 VTAIL.n478 VTAIL.n459 3.49141
R1131 VTAIL.n416 VTAIL.n415 3.49141
R1132 VTAIL.n391 VTAIL.n339 3.49141
R1133 VTAIL.n370 VTAIL.n351 3.49141
R1134 VTAIL.n794 VTAIL.n793 2.71565
R1135 VTAIL.n822 VTAIL.n821 2.71565
R1136 VTAIL.n840 VTAIL.n756 2.71565
R1137 VTAIL.n46 VTAIL.n45 2.71565
R1138 VTAIL.n74 VTAIL.n73 2.71565
R1139 VTAIL.n92 VTAIL.n8 2.71565
R1140 VTAIL.n152 VTAIL.n151 2.71565
R1141 VTAIL.n180 VTAIL.n179 2.71565
R1142 VTAIL.n198 VTAIL.n114 2.71565
R1143 VTAIL.n260 VTAIL.n259 2.71565
R1144 VTAIL.n288 VTAIL.n287 2.71565
R1145 VTAIL.n306 VTAIL.n222 2.71565
R1146 VTAIL.n734 VTAIL.n650 2.71565
R1147 VTAIL.n717 VTAIL.n716 2.71565
R1148 VTAIL.n689 VTAIL.n688 2.71565
R1149 VTAIL.n626 VTAIL.n542 2.71565
R1150 VTAIL.n609 VTAIL.n608 2.71565
R1151 VTAIL.n581 VTAIL.n580 2.71565
R1152 VTAIL.n520 VTAIL.n436 2.71565
R1153 VTAIL.n503 VTAIL.n502 2.71565
R1154 VTAIL.n475 VTAIL.n474 2.71565
R1155 VTAIL.n412 VTAIL.n328 2.71565
R1156 VTAIL.n395 VTAIL.n394 2.71565
R1157 VTAIL.n367 VTAIL.n366 2.71565
R1158 VTAIL.n790 VTAIL.n780 1.93989
R1159 VTAIL.n826 VTAIL.n764 1.93989
R1160 VTAIL.n839 VTAIL.n758 1.93989
R1161 VTAIL.n42 VTAIL.n32 1.93989
R1162 VTAIL.n78 VTAIL.n16 1.93989
R1163 VTAIL.n91 VTAIL.n10 1.93989
R1164 VTAIL.n148 VTAIL.n138 1.93989
R1165 VTAIL.n184 VTAIL.n122 1.93989
R1166 VTAIL.n197 VTAIL.n116 1.93989
R1167 VTAIL.n256 VTAIL.n246 1.93989
R1168 VTAIL.n292 VTAIL.n230 1.93989
R1169 VTAIL.n305 VTAIL.n224 1.93989
R1170 VTAIL.n733 VTAIL.n652 1.93989
R1171 VTAIL.n720 VTAIL.n658 1.93989
R1172 VTAIL.n685 VTAIL.n675 1.93989
R1173 VTAIL.n625 VTAIL.n544 1.93989
R1174 VTAIL.n612 VTAIL.n550 1.93989
R1175 VTAIL.n577 VTAIL.n567 1.93989
R1176 VTAIL.n519 VTAIL.n438 1.93989
R1177 VTAIL.n506 VTAIL.n444 1.93989
R1178 VTAIL.n471 VTAIL.n461 1.93989
R1179 VTAIL.n411 VTAIL.n330 1.93989
R1180 VTAIL.n398 VTAIL.n336 1.93989
R1181 VTAIL.n363 VTAIL.n353 1.93989
R1182 VTAIL.n789 VTAIL.n782 1.16414
R1183 VTAIL.n827 VTAIL.n762 1.16414
R1184 VTAIL.n836 VTAIL.n835 1.16414
R1185 VTAIL.n41 VTAIL.n34 1.16414
R1186 VTAIL.n79 VTAIL.n14 1.16414
R1187 VTAIL.n88 VTAIL.n87 1.16414
R1188 VTAIL.n147 VTAIL.n140 1.16414
R1189 VTAIL.n185 VTAIL.n120 1.16414
R1190 VTAIL.n194 VTAIL.n193 1.16414
R1191 VTAIL.n255 VTAIL.n248 1.16414
R1192 VTAIL.n293 VTAIL.n228 1.16414
R1193 VTAIL.n302 VTAIL.n301 1.16414
R1194 VTAIL.n730 VTAIL.n729 1.16414
R1195 VTAIL.n721 VTAIL.n656 1.16414
R1196 VTAIL.n684 VTAIL.n677 1.16414
R1197 VTAIL.n622 VTAIL.n621 1.16414
R1198 VTAIL.n613 VTAIL.n548 1.16414
R1199 VTAIL.n576 VTAIL.n569 1.16414
R1200 VTAIL.n516 VTAIL.n515 1.16414
R1201 VTAIL.n507 VTAIL.n442 1.16414
R1202 VTAIL.n470 VTAIL.n463 1.16414
R1203 VTAIL.n408 VTAIL.n407 1.16414
R1204 VTAIL.n399 VTAIL.n334 1.16414
R1205 VTAIL.n362 VTAIL.n355 1.16414
R1206 VTAIL.n0 VTAIL.t3 1.04923
R1207 VTAIL.n0 VTAIL.t10 1.04923
R1208 VTAIL.n214 VTAIL.t2 1.04923
R1209 VTAIL.n214 VTAIL.t15 1.04923
R1210 VTAIL.n642 VTAIL.t1 1.04923
R1211 VTAIL.n642 VTAIL.t0 1.04923
R1212 VTAIL.n428 VTAIL.t4 1.04923
R1213 VTAIL.n428 VTAIL.t8 1.04923
R1214 VTAIL.n641 VTAIL.n535 0.470328
R1215 VTAIL.n213 VTAIL.n107 0.470328
R1216 VTAIL.n786 VTAIL.n785 0.388379
R1217 VTAIL.n831 VTAIL.n830 0.388379
R1218 VTAIL.n832 VTAIL.n760 0.388379
R1219 VTAIL.n38 VTAIL.n37 0.388379
R1220 VTAIL.n83 VTAIL.n82 0.388379
R1221 VTAIL.n84 VTAIL.n12 0.388379
R1222 VTAIL.n144 VTAIL.n143 0.388379
R1223 VTAIL.n189 VTAIL.n188 0.388379
R1224 VTAIL.n190 VTAIL.n118 0.388379
R1225 VTAIL.n252 VTAIL.n251 0.388379
R1226 VTAIL.n297 VTAIL.n296 0.388379
R1227 VTAIL.n298 VTAIL.n226 0.388379
R1228 VTAIL.n726 VTAIL.n654 0.388379
R1229 VTAIL.n725 VTAIL.n724 0.388379
R1230 VTAIL.n681 VTAIL.n680 0.388379
R1231 VTAIL.n618 VTAIL.n546 0.388379
R1232 VTAIL.n617 VTAIL.n616 0.388379
R1233 VTAIL.n573 VTAIL.n572 0.388379
R1234 VTAIL.n512 VTAIL.n440 0.388379
R1235 VTAIL.n511 VTAIL.n510 0.388379
R1236 VTAIL.n467 VTAIL.n466 0.388379
R1237 VTAIL.n404 VTAIL.n332 0.388379
R1238 VTAIL.n403 VTAIL.n402 0.388379
R1239 VTAIL.n359 VTAIL.n358 0.388379
R1240 VTAIL.n788 VTAIL.n787 0.155672
R1241 VTAIL.n788 VTAIL.n779 0.155672
R1242 VTAIL.n795 VTAIL.n779 0.155672
R1243 VTAIL.n796 VTAIL.n795 0.155672
R1244 VTAIL.n796 VTAIL.n775 0.155672
R1245 VTAIL.n803 VTAIL.n775 0.155672
R1246 VTAIL.n804 VTAIL.n803 0.155672
R1247 VTAIL.n804 VTAIL.n771 0.155672
R1248 VTAIL.n811 VTAIL.n771 0.155672
R1249 VTAIL.n812 VTAIL.n811 0.155672
R1250 VTAIL.n812 VTAIL.n767 0.155672
R1251 VTAIL.n819 VTAIL.n767 0.155672
R1252 VTAIL.n820 VTAIL.n819 0.155672
R1253 VTAIL.n820 VTAIL.n763 0.155672
R1254 VTAIL.n828 VTAIL.n763 0.155672
R1255 VTAIL.n829 VTAIL.n828 0.155672
R1256 VTAIL.n829 VTAIL.n759 0.155672
R1257 VTAIL.n837 VTAIL.n759 0.155672
R1258 VTAIL.n838 VTAIL.n837 0.155672
R1259 VTAIL.n838 VTAIL.n755 0.155672
R1260 VTAIL.n845 VTAIL.n755 0.155672
R1261 VTAIL.n846 VTAIL.n845 0.155672
R1262 VTAIL.n846 VTAIL.n751 0.155672
R1263 VTAIL.n853 VTAIL.n751 0.155672
R1264 VTAIL.n40 VTAIL.n39 0.155672
R1265 VTAIL.n40 VTAIL.n31 0.155672
R1266 VTAIL.n47 VTAIL.n31 0.155672
R1267 VTAIL.n48 VTAIL.n47 0.155672
R1268 VTAIL.n48 VTAIL.n27 0.155672
R1269 VTAIL.n55 VTAIL.n27 0.155672
R1270 VTAIL.n56 VTAIL.n55 0.155672
R1271 VTAIL.n56 VTAIL.n23 0.155672
R1272 VTAIL.n63 VTAIL.n23 0.155672
R1273 VTAIL.n64 VTAIL.n63 0.155672
R1274 VTAIL.n64 VTAIL.n19 0.155672
R1275 VTAIL.n71 VTAIL.n19 0.155672
R1276 VTAIL.n72 VTAIL.n71 0.155672
R1277 VTAIL.n72 VTAIL.n15 0.155672
R1278 VTAIL.n80 VTAIL.n15 0.155672
R1279 VTAIL.n81 VTAIL.n80 0.155672
R1280 VTAIL.n81 VTAIL.n11 0.155672
R1281 VTAIL.n89 VTAIL.n11 0.155672
R1282 VTAIL.n90 VTAIL.n89 0.155672
R1283 VTAIL.n90 VTAIL.n7 0.155672
R1284 VTAIL.n97 VTAIL.n7 0.155672
R1285 VTAIL.n98 VTAIL.n97 0.155672
R1286 VTAIL.n98 VTAIL.n3 0.155672
R1287 VTAIL.n105 VTAIL.n3 0.155672
R1288 VTAIL.n146 VTAIL.n145 0.155672
R1289 VTAIL.n146 VTAIL.n137 0.155672
R1290 VTAIL.n153 VTAIL.n137 0.155672
R1291 VTAIL.n154 VTAIL.n153 0.155672
R1292 VTAIL.n154 VTAIL.n133 0.155672
R1293 VTAIL.n161 VTAIL.n133 0.155672
R1294 VTAIL.n162 VTAIL.n161 0.155672
R1295 VTAIL.n162 VTAIL.n129 0.155672
R1296 VTAIL.n169 VTAIL.n129 0.155672
R1297 VTAIL.n170 VTAIL.n169 0.155672
R1298 VTAIL.n170 VTAIL.n125 0.155672
R1299 VTAIL.n177 VTAIL.n125 0.155672
R1300 VTAIL.n178 VTAIL.n177 0.155672
R1301 VTAIL.n178 VTAIL.n121 0.155672
R1302 VTAIL.n186 VTAIL.n121 0.155672
R1303 VTAIL.n187 VTAIL.n186 0.155672
R1304 VTAIL.n187 VTAIL.n117 0.155672
R1305 VTAIL.n195 VTAIL.n117 0.155672
R1306 VTAIL.n196 VTAIL.n195 0.155672
R1307 VTAIL.n196 VTAIL.n113 0.155672
R1308 VTAIL.n203 VTAIL.n113 0.155672
R1309 VTAIL.n204 VTAIL.n203 0.155672
R1310 VTAIL.n204 VTAIL.n109 0.155672
R1311 VTAIL.n211 VTAIL.n109 0.155672
R1312 VTAIL.n254 VTAIL.n253 0.155672
R1313 VTAIL.n254 VTAIL.n245 0.155672
R1314 VTAIL.n261 VTAIL.n245 0.155672
R1315 VTAIL.n262 VTAIL.n261 0.155672
R1316 VTAIL.n262 VTAIL.n241 0.155672
R1317 VTAIL.n269 VTAIL.n241 0.155672
R1318 VTAIL.n270 VTAIL.n269 0.155672
R1319 VTAIL.n270 VTAIL.n237 0.155672
R1320 VTAIL.n277 VTAIL.n237 0.155672
R1321 VTAIL.n278 VTAIL.n277 0.155672
R1322 VTAIL.n278 VTAIL.n233 0.155672
R1323 VTAIL.n285 VTAIL.n233 0.155672
R1324 VTAIL.n286 VTAIL.n285 0.155672
R1325 VTAIL.n286 VTAIL.n229 0.155672
R1326 VTAIL.n294 VTAIL.n229 0.155672
R1327 VTAIL.n295 VTAIL.n294 0.155672
R1328 VTAIL.n295 VTAIL.n225 0.155672
R1329 VTAIL.n303 VTAIL.n225 0.155672
R1330 VTAIL.n304 VTAIL.n303 0.155672
R1331 VTAIL.n304 VTAIL.n221 0.155672
R1332 VTAIL.n311 VTAIL.n221 0.155672
R1333 VTAIL.n312 VTAIL.n311 0.155672
R1334 VTAIL.n312 VTAIL.n217 0.155672
R1335 VTAIL.n319 VTAIL.n217 0.155672
R1336 VTAIL.n747 VTAIL.n645 0.155672
R1337 VTAIL.n740 VTAIL.n645 0.155672
R1338 VTAIL.n740 VTAIL.n739 0.155672
R1339 VTAIL.n739 VTAIL.n649 0.155672
R1340 VTAIL.n732 VTAIL.n649 0.155672
R1341 VTAIL.n732 VTAIL.n731 0.155672
R1342 VTAIL.n731 VTAIL.n653 0.155672
R1343 VTAIL.n723 VTAIL.n653 0.155672
R1344 VTAIL.n723 VTAIL.n722 0.155672
R1345 VTAIL.n722 VTAIL.n657 0.155672
R1346 VTAIL.n715 VTAIL.n657 0.155672
R1347 VTAIL.n715 VTAIL.n714 0.155672
R1348 VTAIL.n714 VTAIL.n662 0.155672
R1349 VTAIL.n707 VTAIL.n662 0.155672
R1350 VTAIL.n707 VTAIL.n706 0.155672
R1351 VTAIL.n706 VTAIL.n666 0.155672
R1352 VTAIL.n699 VTAIL.n666 0.155672
R1353 VTAIL.n699 VTAIL.n698 0.155672
R1354 VTAIL.n698 VTAIL.n670 0.155672
R1355 VTAIL.n691 VTAIL.n670 0.155672
R1356 VTAIL.n691 VTAIL.n690 0.155672
R1357 VTAIL.n690 VTAIL.n674 0.155672
R1358 VTAIL.n683 VTAIL.n674 0.155672
R1359 VTAIL.n683 VTAIL.n682 0.155672
R1360 VTAIL.n639 VTAIL.n537 0.155672
R1361 VTAIL.n632 VTAIL.n537 0.155672
R1362 VTAIL.n632 VTAIL.n631 0.155672
R1363 VTAIL.n631 VTAIL.n541 0.155672
R1364 VTAIL.n624 VTAIL.n541 0.155672
R1365 VTAIL.n624 VTAIL.n623 0.155672
R1366 VTAIL.n623 VTAIL.n545 0.155672
R1367 VTAIL.n615 VTAIL.n545 0.155672
R1368 VTAIL.n615 VTAIL.n614 0.155672
R1369 VTAIL.n614 VTAIL.n549 0.155672
R1370 VTAIL.n607 VTAIL.n549 0.155672
R1371 VTAIL.n607 VTAIL.n606 0.155672
R1372 VTAIL.n606 VTAIL.n554 0.155672
R1373 VTAIL.n599 VTAIL.n554 0.155672
R1374 VTAIL.n599 VTAIL.n598 0.155672
R1375 VTAIL.n598 VTAIL.n558 0.155672
R1376 VTAIL.n591 VTAIL.n558 0.155672
R1377 VTAIL.n591 VTAIL.n590 0.155672
R1378 VTAIL.n590 VTAIL.n562 0.155672
R1379 VTAIL.n583 VTAIL.n562 0.155672
R1380 VTAIL.n583 VTAIL.n582 0.155672
R1381 VTAIL.n582 VTAIL.n566 0.155672
R1382 VTAIL.n575 VTAIL.n566 0.155672
R1383 VTAIL.n575 VTAIL.n574 0.155672
R1384 VTAIL.n533 VTAIL.n431 0.155672
R1385 VTAIL.n526 VTAIL.n431 0.155672
R1386 VTAIL.n526 VTAIL.n525 0.155672
R1387 VTAIL.n525 VTAIL.n435 0.155672
R1388 VTAIL.n518 VTAIL.n435 0.155672
R1389 VTAIL.n518 VTAIL.n517 0.155672
R1390 VTAIL.n517 VTAIL.n439 0.155672
R1391 VTAIL.n509 VTAIL.n439 0.155672
R1392 VTAIL.n509 VTAIL.n508 0.155672
R1393 VTAIL.n508 VTAIL.n443 0.155672
R1394 VTAIL.n501 VTAIL.n443 0.155672
R1395 VTAIL.n501 VTAIL.n500 0.155672
R1396 VTAIL.n500 VTAIL.n448 0.155672
R1397 VTAIL.n493 VTAIL.n448 0.155672
R1398 VTAIL.n493 VTAIL.n492 0.155672
R1399 VTAIL.n492 VTAIL.n452 0.155672
R1400 VTAIL.n485 VTAIL.n452 0.155672
R1401 VTAIL.n485 VTAIL.n484 0.155672
R1402 VTAIL.n484 VTAIL.n456 0.155672
R1403 VTAIL.n477 VTAIL.n456 0.155672
R1404 VTAIL.n477 VTAIL.n476 0.155672
R1405 VTAIL.n476 VTAIL.n460 0.155672
R1406 VTAIL.n469 VTAIL.n460 0.155672
R1407 VTAIL.n469 VTAIL.n468 0.155672
R1408 VTAIL.n425 VTAIL.n323 0.155672
R1409 VTAIL.n418 VTAIL.n323 0.155672
R1410 VTAIL.n418 VTAIL.n417 0.155672
R1411 VTAIL.n417 VTAIL.n327 0.155672
R1412 VTAIL.n410 VTAIL.n327 0.155672
R1413 VTAIL.n410 VTAIL.n409 0.155672
R1414 VTAIL.n409 VTAIL.n331 0.155672
R1415 VTAIL.n401 VTAIL.n331 0.155672
R1416 VTAIL.n401 VTAIL.n400 0.155672
R1417 VTAIL.n400 VTAIL.n335 0.155672
R1418 VTAIL.n393 VTAIL.n335 0.155672
R1419 VTAIL.n393 VTAIL.n392 0.155672
R1420 VTAIL.n392 VTAIL.n340 0.155672
R1421 VTAIL.n385 VTAIL.n340 0.155672
R1422 VTAIL.n385 VTAIL.n384 0.155672
R1423 VTAIL.n384 VTAIL.n344 0.155672
R1424 VTAIL.n377 VTAIL.n344 0.155672
R1425 VTAIL.n377 VTAIL.n376 0.155672
R1426 VTAIL.n376 VTAIL.n348 0.155672
R1427 VTAIL.n369 VTAIL.n348 0.155672
R1428 VTAIL.n369 VTAIL.n368 0.155672
R1429 VTAIL.n368 VTAIL.n352 0.155672
R1430 VTAIL.n361 VTAIL.n352 0.155672
R1431 VTAIL.n361 VTAIL.n360 0.155672
R1432 VTAIL VTAIL.n1 0.0586897
R1433 B.n977 B.n976 585
R1434 B.n977 B.n128 585
R1435 B.n980 B.n979 585
R1436 B.n981 B.n199 585
R1437 B.n983 B.n982 585
R1438 B.n985 B.n198 585
R1439 B.n988 B.n987 585
R1440 B.n989 B.n197 585
R1441 B.n991 B.n990 585
R1442 B.n993 B.n196 585
R1443 B.n996 B.n995 585
R1444 B.n997 B.n195 585
R1445 B.n999 B.n998 585
R1446 B.n1001 B.n194 585
R1447 B.n1004 B.n1003 585
R1448 B.n1005 B.n193 585
R1449 B.n1007 B.n1006 585
R1450 B.n1009 B.n192 585
R1451 B.n1012 B.n1011 585
R1452 B.n1013 B.n191 585
R1453 B.n1015 B.n1014 585
R1454 B.n1017 B.n190 585
R1455 B.n1020 B.n1019 585
R1456 B.n1021 B.n189 585
R1457 B.n1023 B.n1022 585
R1458 B.n1025 B.n188 585
R1459 B.n1028 B.n1027 585
R1460 B.n1029 B.n187 585
R1461 B.n1031 B.n1030 585
R1462 B.n1033 B.n186 585
R1463 B.n1036 B.n1035 585
R1464 B.n1037 B.n185 585
R1465 B.n1039 B.n1038 585
R1466 B.n1041 B.n184 585
R1467 B.n1044 B.n1043 585
R1468 B.n1045 B.n183 585
R1469 B.n1047 B.n1046 585
R1470 B.n1049 B.n182 585
R1471 B.n1052 B.n1051 585
R1472 B.n1053 B.n181 585
R1473 B.n1055 B.n1054 585
R1474 B.n1057 B.n180 585
R1475 B.n1060 B.n1059 585
R1476 B.n1061 B.n179 585
R1477 B.n1063 B.n1062 585
R1478 B.n1065 B.n178 585
R1479 B.n1068 B.n1067 585
R1480 B.n1069 B.n177 585
R1481 B.n1071 B.n1070 585
R1482 B.n1073 B.n176 585
R1483 B.n1076 B.n1075 585
R1484 B.n1077 B.n175 585
R1485 B.n1079 B.n1078 585
R1486 B.n1081 B.n174 585
R1487 B.n1084 B.n1083 585
R1488 B.n1085 B.n173 585
R1489 B.n1087 B.n1086 585
R1490 B.n1089 B.n172 585
R1491 B.n1092 B.n1091 585
R1492 B.n1093 B.n171 585
R1493 B.n1095 B.n1094 585
R1494 B.n1097 B.n170 585
R1495 B.n1100 B.n1099 585
R1496 B.n1102 B.n167 585
R1497 B.n1104 B.n1103 585
R1498 B.n1106 B.n166 585
R1499 B.n1109 B.n1108 585
R1500 B.n1110 B.n165 585
R1501 B.n1112 B.n1111 585
R1502 B.n1114 B.n164 585
R1503 B.n1116 B.n1115 585
R1504 B.n1118 B.n1117 585
R1505 B.n1121 B.n1120 585
R1506 B.n1122 B.n159 585
R1507 B.n1124 B.n1123 585
R1508 B.n1126 B.n158 585
R1509 B.n1129 B.n1128 585
R1510 B.n1130 B.n157 585
R1511 B.n1132 B.n1131 585
R1512 B.n1134 B.n156 585
R1513 B.n1137 B.n1136 585
R1514 B.n1138 B.n155 585
R1515 B.n1140 B.n1139 585
R1516 B.n1142 B.n154 585
R1517 B.n1145 B.n1144 585
R1518 B.n1146 B.n153 585
R1519 B.n1148 B.n1147 585
R1520 B.n1150 B.n152 585
R1521 B.n1153 B.n1152 585
R1522 B.n1154 B.n151 585
R1523 B.n1156 B.n1155 585
R1524 B.n1158 B.n150 585
R1525 B.n1161 B.n1160 585
R1526 B.n1162 B.n149 585
R1527 B.n1164 B.n1163 585
R1528 B.n1166 B.n148 585
R1529 B.n1169 B.n1168 585
R1530 B.n1170 B.n147 585
R1531 B.n1172 B.n1171 585
R1532 B.n1174 B.n146 585
R1533 B.n1177 B.n1176 585
R1534 B.n1178 B.n145 585
R1535 B.n1180 B.n1179 585
R1536 B.n1182 B.n144 585
R1537 B.n1185 B.n1184 585
R1538 B.n1186 B.n143 585
R1539 B.n1188 B.n1187 585
R1540 B.n1190 B.n142 585
R1541 B.n1193 B.n1192 585
R1542 B.n1194 B.n141 585
R1543 B.n1196 B.n1195 585
R1544 B.n1198 B.n140 585
R1545 B.n1201 B.n1200 585
R1546 B.n1202 B.n139 585
R1547 B.n1204 B.n1203 585
R1548 B.n1206 B.n138 585
R1549 B.n1209 B.n1208 585
R1550 B.n1210 B.n137 585
R1551 B.n1212 B.n1211 585
R1552 B.n1214 B.n136 585
R1553 B.n1217 B.n1216 585
R1554 B.n1218 B.n135 585
R1555 B.n1220 B.n1219 585
R1556 B.n1222 B.n134 585
R1557 B.n1225 B.n1224 585
R1558 B.n1226 B.n133 585
R1559 B.n1228 B.n1227 585
R1560 B.n1230 B.n132 585
R1561 B.n1233 B.n1232 585
R1562 B.n1234 B.n131 585
R1563 B.n1236 B.n1235 585
R1564 B.n1238 B.n130 585
R1565 B.n1241 B.n1240 585
R1566 B.n1242 B.n129 585
R1567 B.n975 B.n127 585
R1568 B.n1245 B.n127 585
R1569 B.n974 B.n126 585
R1570 B.n1246 B.n126 585
R1571 B.n973 B.n125 585
R1572 B.n1247 B.n125 585
R1573 B.n972 B.n971 585
R1574 B.n971 B.n121 585
R1575 B.n970 B.n120 585
R1576 B.n1253 B.n120 585
R1577 B.n969 B.n119 585
R1578 B.n1254 B.n119 585
R1579 B.n968 B.n118 585
R1580 B.n1255 B.n118 585
R1581 B.n967 B.n966 585
R1582 B.n966 B.n114 585
R1583 B.n965 B.n113 585
R1584 B.n1261 B.n113 585
R1585 B.n964 B.n112 585
R1586 B.n1262 B.n112 585
R1587 B.n963 B.n111 585
R1588 B.n1263 B.n111 585
R1589 B.n962 B.n961 585
R1590 B.n961 B.n107 585
R1591 B.n960 B.n106 585
R1592 B.n1269 B.n106 585
R1593 B.n959 B.n105 585
R1594 B.n1270 B.n105 585
R1595 B.n958 B.n104 585
R1596 B.n1271 B.n104 585
R1597 B.n957 B.n956 585
R1598 B.n956 B.n100 585
R1599 B.n955 B.n99 585
R1600 B.n1277 B.n99 585
R1601 B.n954 B.n98 585
R1602 B.n1278 B.n98 585
R1603 B.n953 B.n97 585
R1604 B.n1279 B.n97 585
R1605 B.n952 B.n951 585
R1606 B.n951 B.n93 585
R1607 B.n950 B.n92 585
R1608 B.n1285 B.n92 585
R1609 B.n949 B.n91 585
R1610 B.n1286 B.n91 585
R1611 B.n948 B.n90 585
R1612 B.n1287 B.n90 585
R1613 B.n947 B.n946 585
R1614 B.n946 B.n86 585
R1615 B.n945 B.n85 585
R1616 B.n1293 B.n85 585
R1617 B.n944 B.n84 585
R1618 B.n1294 B.n84 585
R1619 B.n943 B.n83 585
R1620 B.n1295 B.n83 585
R1621 B.n942 B.n941 585
R1622 B.n941 B.n79 585
R1623 B.n940 B.n78 585
R1624 B.n1301 B.n78 585
R1625 B.n939 B.n77 585
R1626 B.n1302 B.n77 585
R1627 B.n938 B.n76 585
R1628 B.n1303 B.n76 585
R1629 B.n937 B.n936 585
R1630 B.n936 B.n72 585
R1631 B.n935 B.n71 585
R1632 B.n1309 B.n71 585
R1633 B.n934 B.n70 585
R1634 B.n1310 B.n70 585
R1635 B.n933 B.n69 585
R1636 B.n1311 B.n69 585
R1637 B.n932 B.n931 585
R1638 B.n931 B.n65 585
R1639 B.n930 B.n64 585
R1640 B.n1317 B.n64 585
R1641 B.n929 B.n63 585
R1642 B.n1318 B.n63 585
R1643 B.n928 B.n62 585
R1644 B.n1319 B.n62 585
R1645 B.n927 B.n926 585
R1646 B.n926 B.n58 585
R1647 B.n925 B.n57 585
R1648 B.n1325 B.n57 585
R1649 B.n924 B.n56 585
R1650 B.n1326 B.n56 585
R1651 B.n923 B.n55 585
R1652 B.n1327 B.n55 585
R1653 B.n922 B.n921 585
R1654 B.n921 B.n51 585
R1655 B.n920 B.n50 585
R1656 B.n1333 B.n50 585
R1657 B.n919 B.n49 585
R1658 B.n1334 B.n49 585
R1659 B.n918 B.n48 585
R1660 B.n1335 B.n48 585
R1661 B.n917 B.n916 585
R1662 B.n916 B.n44 585
R1663 B.n915 B.n43 585
R1664 B.n1341 B.n43 585
R1665 B.n914 B.n42 585
R1666 B.n1342 B.n42 585
R1667 B.n913 B.n41 585
R1668 B.n1343 B.n41 585
R1669 B.n912 B.n911 585
R1670 B.n911 B.n37 585
R1671 B.n910 B.n36 585
R1672 B.n1349 B.n36 585
R1673 B.n909 B.n35 585
R1674 B.n1350 B.n35 585
R1675 B.n908 B.n34 585
R1676 B.n1351 B.n34 585
R1677 B.n907 B.n906 585
R1678 B.n906 B.n30 585
R1679 B.n905 B.n29 585
R1680 B.n1357 B.n29 585
R1681 B.n904 B.n28 585
R1682 B.n1358 B.n28 585
R1683 B.n903 B.n27 585
R1684 B.n1359 B.n27 585
R1685 B.n902 B.n901 585
R1686 B.n901 B.n23 585
R1687 B.n900 B.n22 585
R1688 B.n1365 B.n22 585
R1689 B.n899 B.n21 585
R1690 B.n1366 B.n21 585
R1691 B.n898 B.n20 585
R1692 B.n1367 B.n20 585
R1693 B.n897 B.n896 585
R1694 B.n896 B.n16 585
R1695 B.n895 B.n15 585
R1696 B.n1373 B.n15 585
R1697 B.n894 B.n14 585
R1698 B.n1374 B.n14 585
R1699 B.n893 B.n13 585
R1700 B.n1375 B.n13 585
R1701 B.n892 B.n891 585
R1702 B.n891 B.n12 585
R1703 B.n890 B.n889 585
R1704 B.n890 B.n8 585
R1705 B.n888 B.n7 585
R1706 B.n1382 B.n7 585
R1707 B.n887 B.n6 585
R1708 B.n1383 B.n6 585
R1709 B.n886 B.n5 585
R1710 B.n1384 B.n5 585
R1711 B.n885 B.n884 585
R1712 B.n884 B.n4 585
R1713 B.n883 B.n200 585
R1714 B.n883 B.n882 585
R1715 B.n873 B.n201 585
R1716 B.n202 B.n201 585
R1717 B.n875 B.n874 585
R1718 B.n876 B.n875 585
R1719 B.n872 B.n207 585
R1720 B.n207 B.n206 585
R1721 B.n871 B.n870 585
R1722 B.n870 B.n869 585
R1723 B.n209 B.n208 585
R1724 B.n210 B.n209 585
R1725 B.n862 B.n861 585
R1726 B.n863 B.n862 585
R1727 B.n860 B.n215 585
R1728 B.n215 B.n214 585
R1729 B.n859 B.n858 585
R1730 B.n858 B.n857 585
R1731 B.n217 B.n216 585
R1732 B.n218 B.n217 585
R1733 B.n850 B.n849 585
R1734 B.n851 B.n850 585
R1735 B.n848 B.n223 585
R1736 B.n223 B.n222 585
R1737 B.n847 B.n846 585
R1738 B.n846 B.n845 585
R1739 B.n225 B.n224 585
R1740 B.n226 B.n225 585
R1741 B.n838 B.n837 585
R1742 B.n839 B.n838 585
R1743 B.n836 B.n231 585
R1744 B.n231 B.n230 585
R1745 B.n835 B.n834 585
R1746 B.n834 B.n833 585
R1747 B.n233 B.n232 585
R1748 B.n234 B.n233 585
R1749 B.n826 B.n825 585
R1750 B.n827 B.n826 585
R1751 B.n824 B.n239 585
R1752 B.n239 B.n238 585
R1753 B.n823 B.n822 585
R1754 B.n822 B.n821 585
R1755 B.n241 B.n240 585
R1756 B.n242 B.n241 585
R1757 B.n814 B.n813 585
R1758 B.n815 B.n814 585
R1759 B.n812 B.n247 585
R1760 B.n247 B.n246 585
R1761 B.n811 B.n810 585
R1762 B.n810 B.n809 585
R1763 B.n249 B.n248 585
R1764 B.n250 B.n249 585
R1765 B.n802 B.n801 585
R1766 B.n803 B.n802 585
R1767 B.n800 B.n255 585
R1768 B.n255 B.n254 585
R1769 B.n799 B.n798 585
R1770 B.n798 B.n797 585
R1771 B.n257 B.n256 585
R1772 B.n258 B.n257 585
R1773 B.n790 B.n789 585
R1774 B.n791 B.n790 585
R1775 B.n788 B.n262 585
R1776 B.n266 B.n262 585
R1777 B.n787 B.n786 585
R1778 B.n786 B.n785 585
R1779 B.n264 B.n263 585
R1780 B.n265 B.n264 585
R1781 B.n778 B.n777 585
R1782 B.n779 B.n778 585
R1783 B.n776 B.n271 585
R1784 B.n271 B.n270 585
R1785 B.n775 B.n774 585
R1786 B.n774 B.n773 585
R1787 B.n273 B.n272 585
R1788 B.n274 B.n273 585
R1789 B.n766 B.n765 585
R1790 B.n767 B.n766 585
R1791 B.n764 B.n279 585
R1792 B.n279 B.n278 585
R1793 B.n763 B.n762 585
R1794 B.n762 B.n761 585
R1795 B.n281 B.n280 585
R1796 B.n282 B.n281 585
R1797 B.n754 B.n753 585
R1798 B.n755 B.n754 585
R1799 B.n752 B.n286 585
R1800 B.n290 B.n286 585
R1801 B.n751 B.n750 585
R1802 B.n750 B.n749 585
R1803 B.n288 B.n287 585
R1804 B.n289 B.n288 585
R1805 B.n742 B.n741 585
R1806 B.n743 B.n742 585
R1807 B.n740 B.n295 585
R1808 B.n295 B.n294 585
R1809 B.n739 B.n738 585
R1810 B.n738 B.n737 585
R1811 B.n297 B.n296 585
R1812 B.n298 B.n297 585
R1813 B.n730 B.n729 585
R1814 B.n731 B.n730 585
R1815 B.n728 B.n303 585
R1816 B.n303 B.n302 585
R1817 B.n727 B.n726 585
R1818 B.n726 B.n725 585
R1819 B.n305 B.n304 585
R1820 B.n306 B.n305 585
R1821 B.n718 B.n717 585
R1822 B.n719 B.n718 585
R1823 B.n716 B.n311 585
R1824 B.n311 B.n310 585
R1825 B.n715 B.n714 585
R1826 B.n714 B.n713 585
R1827 B.n313 B.n312 585
R1828 B.n314 B.n313 585
R1829 B.n706 B.n705 585
R1830 B.n707 B.n706 585
R1831 B.n704 B.n318 585
R1832 B.n322 B.n318 585
R1833 B.n703 B.n702 585
R1834 B.n702 B.n701 585
R1835 B.n320 B.n319 585
R1836 B.n321 B.n320 585
R1837 B.n694 B.n693 585
R1838 B.n695 B.n694 585
R1839 B.n692 B.n327 585
R1840 B.n327 B.n326 585
R1841 B.n691 B.n690 585
R1842 B.n690 B.n689 585
R1843 B.n329 B.n328 585
R1844 B.n330 B.n329 585
R1845 B.n682 B.n681 585
R1846 B.n683 B.n682 585
R1847 B.n680 B.n335 585
R1848 B.n335 B.n334 585
R1849 B.n679 B.n678 585
R1850 B.n678 B.n677 585
R1851 B.n674 B.n339 585
R1852 B.n673 B.n672 585
R1853 B.n670 B.n340 585
R1854 B.n670 B.n338 585
R1855 B.n669 B.n668 585
R1856 B.n667 B.n666 585
R1857 B.n665 B.n342 585
R1858 B.n663 B.n662 585
R1859 B.n661 B.n343 585
R1860 B.n660 B.n659 585
R1861 B.n657 B.n344 585
R1862 B.n655 B.n654 585
R1863 B.n653 B.n345 585
R1864 B.n652 B.n651 585
R1865 B.n649 B.n346 585
R1866 B.n647 B.n646 585
R1867 B.n645 B.n347 585
R1868 B.n644 B.n643 585
R1869 B.n641 B.n348 585
R1870 B.n639 B.n638 585
R1871 B.n637 B.n349 585
R1872 B.n636 B.n635 585
R1873 B.n633 B.n350 585
R1874 B.n631 B.n630 585
R1875 B.n629 B.n351 585
R1876 B.n628 B.n627 585
R1877 B.n625 B.n352 585
R1878 B.n623 B.n622 585
R1879 B.n621 B.n353 585
R1880 B.n620 B.n619 585
R1881 B.n617 B.n354 585
R1882 B.n615 B.n614 585
R1883 B.n613 B.n355 585
R1884 B.n612 B.n611 585
R1885 B.n609 B.n356 585
R1886 B.n607 B.n606 585
R1887 B.n605 B.n357 585
R1888 B.n604 B.n603 585
R1889 B.n601 B.n358 585
R1890 B.n599 B.n598 585
R1891 B.n597 B.n359 585
R1892 B.n596 B.n595 585
R1893 B.n593 B.n360 585
R1894 B.n591 B.n590 585
R1895 B.n589 B.n361 585
R1896 B.n588 B.n587 585
R1897 B.n585 B.n362 585
R1898 B.n583 B.n582 585
R1899 B.n581 B.n363 585
R1900 B.n580 B.n579 585
R1901 B.n577 B.n364 585
R1902 B.n575 B.n574 585
R1903 B.n573 B.n365 585
R1904 B.n572 B.n571 585
R1905 B.n569 B.n366 585
R1906 B.n567 B.n566 585
R1907 B.n565 B.n367 585
R1908 B.n564 B.n563 585
R1909 B.n561 B.n368 585
R1910 B.n559 B.n558 585
R1911 B.n557 B.n369 585
R1912 B.n556 B.n555 585
R1913 B.n553 B.n370 585
R1914 B.n551 B.n550 585
R1915 B.n549 B.n371 585
R1916 B.n548 B.n547 585
R1917 B.n545 B.n375 585
R1918 B.n543 B.n542 585
R1919 B.n541 B.n376 585
R1920 B.n540 B.n539 585
R1921 B.n537 B.n377 585
R1922 B.n535 B.n534 585
R1923 B.n532 B.n378 585
R1924 B.n531 B.n530 585
R1925 B.n528 B.n381 585
R1926 B.n526 B.n525 585
R1927 B.n524 B.n382 585
R1928 B.n523 B.n522 585
R1929 B.n520 B.n383 585
R1930 B.n518 B.n517 585
R1931 B.n516 B.n384 585
R1932 B.n515 B.n514 585
R1933 B.n512 B.n385 585
R1934 B.n510 B.n509 585
R1935 B.n508 B.n386 585
R1936 B.n507 B.n506 585
R1937 B.n504 B.n387 585
R1938 B.n502 B.n501 585
R1939 B.n500 B.n388 585
R1940 B.n499 B.n498 585
R1941 B.n496 B.n389 585
R1942 B.n494 B.n493 585
R1943 B.n492 B.n390 585
R1944 B.n491 B.n490 585
R1945 B.n488 B.n391 585
R1946 B.n486 B.n485 585
R1947 B.n484 B.n392 585
R1948 B.n483 B.n482 585
R1949 B.n480 B.n393 585
R1950 B.n478 B.n477 585
R1951 B.n476 B.n394 585
R1952 B.n475 B.n474 585
R1953 B.n472 B.n395 585
R1954 B.n470 B.n469 585
R1955 B.n468 B.n396 585
R1956 B.n467 B.n466 585
R1957 B.n464 B.n397 585
R1958 B.n462 B.n461 585
R1959 B.n460 B.n398 585
R1960 B.n459 B.n458 585
R1961 B.n456 B.n399 585
R1962 B.n454 B.n453 585
R1963 B.n452 B.n400 585
R1964 B.n451 B.n450 585
R1965 B.n448 B.n401 585
R1966 B.n446 B.n445 585
R1967 B.n444 B.n402 585
R1968 B.n443 B.n442 585
R1969 B.n440 B.n403 585
R1970 B.n438 B.n437 585
R1971 B.n436 B.n404 585
R1972 B.n435 B.n434 585
R1973 B.n432 B.n405 585
R1974 B.n430 B.n429 585
R1975 B.n428 B.n406 585
R1976 B.n427 B.n426 585
R1977 B.n424 B.n407 585
R1978 B.n422 B.n421 585
R1979 B.n420 B.n408 585
R1980 B.n419 B.n418 585
R1981 B.n416 B.n409 585
R1982 B.n414 B.n413 585
R1983 B.n412 B.n411 585
R1984 B.n337 B.n336 585
R1985 B.n676 B.n675 585
R1986 B.n677 B.n676 585
R1987 B.n333 B.n332 585
R1988 B.n334 B.n333 585
R1989 B.n685 B.n684 585
R1990 B.n684 B.n683 585
R1991 B.n686 B.n331 585
R1992 B.n331 B.n330 585
R1993 B.n688 B.n687 585
R1994 B.n689 B.n688 585
R1995 B.n325 B.n324 585
R1996 B.n326 B.n325 585
R1997 B.n697 B.n696 585
R1998 B.n696 B.n695 585
R1999 B.n698 B.n323 585
R2000 B.n323 B.n321 585
R2001 B.n700 B.n699 585
R2002 B.n701 B.n700 585
R2003 B.n317 B.n316 585
R2004 B.n322 B.n317 585
R2005 B.n709 B.n708 585
R2006 B.n708 B.n707 585
R2007 B.n710 B.n315 585
R2008 B.n315 B.n314 585
R2009 B.n712 B.n711 585
R2010 B.n713 B.n712 585
R2011 B.n309 B.n308 585
R2012 B.n310 B.n309 585
R2013 B.n721 B.n720 585
R2014 B.n720 B.n719 585
R2015 B.n722 B.n307 585
R2016 B.n307 B.n306 585
R2017 B.n724 B.n723 585
R2018 B.n725 B.n724 585
R2019 B.n301 B.n300 585
R2020 B.n302 B.n301 585
R2021 B.n733 B.n732 585
R2022 B.n732 B.n731 585
R2023 B.n734 B.n299 585
R2024 B.n299 B.n298 585
R2025 B.n736 B.n735 585
R2026 B.n737 B.n736 585
R2027 B.n293 B.n292 585
R2028 B.n294 B.n293 585
R2029 B.n745 B.n744 585
R2030 B.n744 B.n743 585
R2031 B.n746 B.n291 585
R2032 B.n291 B.n289 585
R2033 B.n748 B.n747 585
R2034 B.n749 B.n748 585
R2035 B.n285 B.n284 585
R2036 B.n290 B.n285 585
R2037 B.n757 B.n756 585
R2038 B.n756 B.n755 585
R2039 B.n758 B.n283 585
R2040 B.n283 B.n282 585
R2041 B.n760 B.n759 585
R2042 B.n761 B.n760 585
R2043 B.n277 B.n276 585
R2044 B.n278 B.n277 585
R2045 B.n769 B.n768 585
R2046 B.n768 B.n767 585
R2047 B.n770 B.n275 585
R2048 B.n275 B.n274 585
R2049 B.n772 B.n771 585
R2050 B.n773 B.n772 585
R2051 B.n269 B.n268 585
R2052 B.n270 B.n269 585
R2053 B.n781 B.n780 585
R2054 B.n780 B.n779 585
R2055 B.n782 B.n267 585
R2056 B.n267 B.n265 585
R2057 B.n784 B.n783 585
R2058 B.n785 B.n784 585
R2059 B.n261 B.n260 585
R2060 B.n266 B.n261 585
R2061 B.n793 B.n792 585
R2062 B.n792 B.n791 585
R2063 B.n794 B.n259 585
R2064 B.n259 B.n258 585
R2065 B.n796 B.n795 585
R2066 B.n797 B.n796 585
R2067 B.n253 B.n252 585
R2068 B.n254 B.n253 585
R2069 B.n805 B.n804 585
R2070 B.n804 B.n803 585
R2071 B.n806 B.n251 585
R2072 B.n251 B.n250 585
R2073 B.n808 B.n807 585
R2074 B.n809 B.n808 585
R2075 B.n245 B.n244 585
R2076 B.n246 B.n245 585
R2077 B.n817 B.n816 585
R2078 B.n816 B.n815 585
R2079 B.n818 B.n243 585
R2080 B.n243 B.n242 585
R2081 B.n820 B.n819 585
R2082 B.n821 B.n820 585
R2083 B.n237 B.n236 585
R2084 B.n238 B.n237 585
R2085 B.n829 B.n828 585
R2086 B.n828 B.n827 585
R2087 B.n830 B.n235 585
R2088 B.n235 B.n234 585
R2089 B.n832 B.n831 585
R2090 B.n833 B.n832 585
R2091 B.n229 B.n228 585
R2092 B.n230 B.n229 585
R2093 B.n841 B.n840 585
R2094 B.n840 B.n839 585
R2095 B.n842 B.n227 585
R2096 B.n227 B.n226 585
R2097 B.n844 B.n843 585
R2098 B.n845 B.n844 585
R2099 B.n221 B.n220 585
R2100 B.n222 B.n221 585
R2101 B.n853 B.n852 585
R2102 B.n852 B.n851 585
R2103 B.n854 B.n219 585
R2104 B.n219 B.n218 585
R2105 B.n856 B.n855 585
R2106 B.n857 B.n856 585
R2107 B.n213 B.n212 585
R2108 B.n214 B.n213 585
R2109 B.n865 B.n864 585
R2110 B.n864 B.n863 585
R2111 B.n866 B.n211 585
R2112 B.n211 B.n210 585
R2113 B.n868 B.n867 585
R2114 B.n869 B.n868 585
R2115 B.n205 B.n204 585
R2116 B.n206 B.n205 585
R2117 B.n878 B.n877 585
R2118 B.n877 B.n876 585
R2119 B.n879 B.n203 585
R2120 B.n203 B.n202 585
R2121 B.n881 B.n880 585
R2122 B.n882 B.n881 585
R2123 B.n3 B.n0 585
R2124 B.n4 B.n3 585
R2125 B.n1381 B.n1 585
R2126 B.n1382 B.n1381 585
R2127 B.n1380 B.n1379 585
R2128 B.n1380 B.n8 585
R2129 B.n1378 B.n9 585
R2130 B.n12 B.n9 585
R2131 B.n1377 B.n1376 585
R2132 B.n1376 B.n1375 585
R2133 B.n11 B.n10 585
R2134 B.n1374 B.n11 585
R2135 B.n1372 B.n1371 585
R2136 B.n1373 B.n1372 585
R2137 B.n1370 B.n17 585
R2138 B.n17 B.n16 585
R2139 B.n1369 B.n1368 585
R2140 B.n1368 B.n1367 585
R2141 B.n19 B.n18 585
R2142 B.n1366 B.n19 585
R2143 B.n1364 B.n1363 585
R2144 B.n1365 B.n1364 585
R2145 B.n1362 B.n24 585
R2146 B.n24 B.n23 585
R2147 B.n1361 B.n1360 585
R2148 B.n1360 B.n1359 585
R2149 B.n26 B.n25 585
R2150 B.n1358 B.n26 585
R2151 B.n1356 B.n1355 585
R2152 B.n1357 B.n1356 585
R2153 B.n1354 B.n31 585
R2154 B.n31 B.n30 585
R2155 B.n1353 B.n1352 585
R2156 B.n1352 B.n1351 585
R2157 B.n33 B.n32 585
R2158 B.n1350 B.n33 585
R2159 B.n1348 B.n1347 585
R2160 B.n1349 B.n1348 585
R2161 B.n1346 B.n38 585
R2162 B.n38 B.n37 585
R2163 B.n1345 B.n1344 585
R2164 B.n1344 B.n1343 585
R2165 B.n40 B.n39 585
R2166 B.n1342 B.n40 585
R2167 B.n1340 B.n1339 585
R2168 B.n1341 B.n1340 585
R2169 B.n1338 B.n45 585
R2170 B.n45 B.n44 585
R2171 B.n1337 B.n1336 585
R2172 B.n1336 B.n1335 585
R2173 B.n47 B.n46 585
R2174 B.n1334 B.n47 585
R2175 B.n1332 B.n1331 585
R2176 B.n1333 B.n1332 585
R2177 B.n1330 B.n52 585
R2178 B.n52 B.n51 585
R2179 B.n1329 B.n1328 585
R2180 B.n1328 B.n1327 585
R2181 B.n54 B.n53 585
R2182 B.n1326 B.n54 585
R2183 B.n1324 B.n1323 585
R2184 B.n1325 B.n1324 585
R2185 B.n1322 B.n59 585
R2186 B.n59 B.n58 585
R2187 B.n1321 B.n1320 585
R2188 B.n1320 B.n1319 585
R2189 B.n61 B.n60 585
R2190 B.n1318 B.n61 585
R2191 B.n1316 B.n1315 585
R2192 B.n1317 B.n1316 585
R2193 B.n1314 B.n66 585
R2194 B.n66 B.n65 585
R2195 B.n1313 B.n1312 585
R2196 B.n1312 B.n1311 585
R2197 B.n68 B.n67 585
R2198 B.n1310 B.n68 585
R2199 B.n1308 B.n1307 585
R2200 B.n1309 B.n1308 585
R2201 B.n1306 B.n73 585
R2202 B.n73 B.n72 585
R2203 B.n1305 B.n1304 585
R2204 B.n1304 B.n1303 585
R2205 B.n75 B.n74 585
R2206 B.n1302 B.n75 585
R2207 B.n1300 B.n1299 585
R2208 B.n1301 B.n1300 585
R2209 B.n1298 B.n80 585
R2210 B.n80 B.n79 585
R2211 B.n1297 B.n1296 585
R2212 B.n1296 B.n1295 585
R2213 B.n82 B.n81 585
R2214 B.n1294 B.n82 585
R2215 B.n1292 B.n1291 585
R2216 B.n1293 B.n1292 585
R2217 B.n1290 B.n87 585
R2218 B.n87 B.n86 585
R2219 B.n1289 B.n1288 585
R2220 B.n1288 B.n1287 585
R2221 B.n89 B.n88 585
R2222 B.n1286 B.n89 585
R2223 B.n1284 B.n1283 585
R2224 B.n1285 B.n1284 585
R2225 B.n1282 B.n94 585
R2226 B.n94 B.n93 585
R2227 B.n1281 B.n1280 585
R2228 B.n1280 B.n1279 585
R2229 B.n96 B.n95 585
R2230 B.n1278 B.n96 585
R2231 B.n1276 B.n1275 585
R2232 B.n1277 B.n1276 585
R2233 B.n1274 B.n101 585
R2234 B.n101 B.n100 585
R2235 B.n1273 B.n1272 585
R2236 B.n1272 B.n1271 585
R2237 B.n103 B.n102 585
R2238 B.n1270 B.n103 585
R2239 B.n1268 B.n1267 585
R2240 B.n1269 B.n1268 585
R2241 B.n1266 B.n108 585
R2242 B.n108 B.n107 585
R2243 B.n1265 B.n1264 585
R2244 B.n1264 B.n1263 585
R2245 B.n110 B.n109 585
R2246 B.n1262 B.n110 585
R2247 B.n1260 B.n1259 585
R2248 B.n1261 B.n1260 585
R2249 B.n1258 B.n115 585
R2250 B.n115 B.n114 585
R2251 B.n1257 B.n1256 585
R2252 B.n1256 B.n1255 585
R2253 B.n117 B.n116 585
R2254 B.n1254 B.n117 585
R2255 B.n1252 B.n1251 585
R2256 B.n1253 B.n1252 585
R2257 B.n1250 B.n122 585
R2258 B.n122 B.n121 585
R2259 B.n1249 B.n1248 585
R2260 B.n1248 B.n1247 585
R2261 B.n124 B.n123 585
R2262 B.n1246 B.n124 585
R2263 B.n1244 B.n1243 585
R2264 B.n1245 B.n1244 585
R2265 B.n1385 B.n1384 585
R2266 B.n1383 B.n2 585
R2267 B.n1244 B.n129 516.524
R2268 B.n977 B.n127 516.524
R2269 B.n678 B.n337 516.524
R2270 B.n676 B.n339 516.524
R2271 B.n168 B.t14 482.914
R2272 B.n379 B.t11 482.914
R2273 B.n160 B.t20 482.914
R2274 B.n372 B.t18 482.914
R2275 B.n169 B.t15 400.683
R2276 B.n380 B.t10 400.683
R2277 B.n161 B.t21 400.683
R2278 B.n373 B.t17 400.683
R2279 B.n160 B.t19 325.798
R2280 B.n168 B.t12 325.798
R2281 B.n379 B.t8 325.798
R2282 B.n372 B.t16 325.798
R2283 B.n978 B.n128 256.663
R2284 B.n984 B.n128 256.663
R2285 B.n986 B.n128 256.663
R2286 B.n992 B.n128 256.663
R2287 B.n994 B.n128 256.663
R2288 B.n1000 B.n128 256.663
R2289 B.n1002 B.n128 256.663
R2290 B.n1008 B.n128 256.663
R2291 B.n1010 B.n128 256.663
R2292 B.n1016 B.n128 256.663
R2293 B.n1018 B.n128 256.663
R2294 B.n1024 B.n128 256.663
R2295 B.n1026 B.n128 256.663
R2296 B.n1032 B.n128 256.663
R2297 B.n1034 B.n128 256.663
R2298 B.n1040 B.n128 256.663
R2299 B.n1042 B.n128 256.663
R2300 B.n1048 B.n128 256.663
R2301 B.n1050 B.n128 256.663
R2302 B.n1056 B.n128 256.663
R2303 B.n1058 B.n128 256.663
R2304 B.n1064 B.n128 256.663
R2305 B.n1066 B.n128 256.663
R2306 B.n1072 B.n128 256.663
R2307 B.n1074 B.n128 256.663
R2308 B.n1080 B.n128 256.663
R2309 B.n1082 B.n128 256.663
R2310 B.n1088 B.n128 256.663
R2311 B.n1090 B.n128 256.663
R2312 B.n1096 B.n128 256.663
R2313 B.n1098 B.n128 256.663
R2314 B.n1105 B.n128 256.663
R2315 B.n1107 B.n128 256.663
R2316 B.n1113 B.n128 256.663
R2317 B.n163 B.n128 256.663
R2318 B.n1119 B.n128 256.663
R2319 B.n1125 B.n128 256.663
R2320 B.n1127 B.n128 256.663
R2321 B.n1133 B.n128 256.663
R2322 B.n1135 B.n128 256.663
R2323 B.n1141 B.n128 256.663
R2324 B.n1143 B.n128 256.663
R2325 B.n1149 B.n128 256.663
R2326 B.n1151 B.n128 256.663
R2327 B.n1157 B.n128 256.663
R2328 B.n1159 B.n128 256.663
R2329 B.n1165 B.n128 256.663
R2330 B.n1167 B.n128 256.663
R2331 B.n1173 B.n128 256.663
R2332 B.n1175 B.n128 256.663
R2333 B.n1181 B.n128 256.663
R2334 B.n1183 B.n128 256.663
R2335 B.n1189 B.n128 256.663
R2336 B.n1191 B.n128 256.663
R2337 B.n1197 B.n128 256.663
R2338 B.n1199 B.n128 256.663
R2339 B.n1205 B.n128 256.663
R2340 B.n1207 B.n128 256.663
R2341 B.n1213 B.n128 256.663
R2342 B.n1215 B.n128 256.663
R2343 B.n1221 B.n128 256.663
R2344 B.n1223 B.n128 256.663
R2345 B.n1229 B.n128 256.663
R2346 B.n1231 B.n128 256.663
R2347 B.n1237 B.n128 256.663
R2348 B.n1239 B.n128 256.663
R2349 B.n671 B.n338 256.663
R2350 B.n341 B.n338 256.663
R2351 B.n664 B.n338 256.663
R2352 B.n658 B.n338 256.663
R2353 B.n656 B.n338 256.663
R2354 B.n650 B.n338 256.663
R2355 B.n648 B.n338 256.663
R2356 B.n642 B.n338 256.663
R2357 B.n640 B.n338 256.663
R2358 B.n634 B.n338 256.663
R2359 B.n632 B.n338 256.663
R2360 B.n626 B.n338 256.663
R2361 B.n624 B.n338 256.663
R2362 B.n618 B.n338 256.663
R2363 B.n616 B.n338 256.663
R2364 B.n610 B.n338 256.663
R2365 B.n608 B.n338 256.663
R2366 B.n602 B.n338 256.663
R2367 B.n600 B.n338 256.663
R2368 B.n594 B.n338 256.663
R2369 B.n592 B.n338 256.663
R2370 B.n586 B.n338 256.663
R2371 B.n584 B.n338 256.663
R2372 B.n578 B.n338 256.663
R2373 B.n576 B.n338 256.663
R2374 B.n570 B.n338 256.663
R2375 B.n568 B.n338 256.663
R2376 B.n562 B.n338 256.663
R2377 B.n560 B.n338 256.663
R2378 B.n554 B.n338 256.663
R2379 B.n552 B.n338 256.663
R2380 B.n546 B.n338 256.663
R2381 B.n544 B.n338 256.663
R2382 B.n538 B.n338 256.663
R2383 B.n536 B.n338 256.663
R2384 B.n529 B.n338 256.663
R2385 B.n527 B.n338 256.663
R2386 B.n521 B.n338 256.663
R2387 B.n519 B.n338 256.663
R2388 B.n513 B.n338 256.663
R2389 B.n511 B.n338 256.663
R2390 B.n505 B.n338 256.663
R2391 B.n503 B.n338 256.663
R2392 B.n497 B.n338 256.663
R2393 B.n495 B.n338 256.663
R2394 B.n489 B.n338 256.663
R2395 B.n487 B.n338 256.663
R2396 B.n481 B.n338 256.663
R2397 B.n479 B.n338 256.663
R2398 B.n473 B.n338 256.663
R2399 B.n471 B.n338 256.663
R2400 B.n465 B.n338 256.663
R2401 B.n463 B.n338 256.663
R2402 B.n457 B.n338 256.663
R2403 B.n455 B.n338 256.663
R2404 B.n449 B.n338 256.663
R2405 B.n447 B.n338 256.663
R2406 B.n441 B.n338 256.663
R2407 B.n439 B.n338 256.663
R2408 B.n433 B.n338 256.663
R2409 B.n431 B.n338 256.663
R2410 B.n425 B.n338 256.663
R2411 B.n423 B.n338 256.663
R2412 B.n417 B.n338 256.663
R2413 B.n415 B.n338 256.663
R2414 B.n410 B.n338 256.663
R2415 B.n1387 B.n1386 256.663
R2416 B.n1240 B.n1238 163.367
R2417 B.n1236 B.n131 163.367
R2418 B.n1232 B.n1230 163.367
R2419 B.n1228 B.n133 163.367
R2420 B.n1224 B.n1222 163.367
R2421 B.n1220 B.n135 163.367
R2422 B.n1216 B.n1214 163.367
R2423 B.n1212 B.n137 163.367
R2424 B.n1208 B.n1206 163.367
R2425 B.n1204 B.n139 163.367
R2426 B.n1200 B.n1198 163.367
R2427 B.n1196 B.n141 163.367
R2428 B.n1192 B.n1190 163.367
R2429 B.n1188 B.n143 163.367
R2430 B.n1184 B.n1182 163.367
R2431 B.n1180 B.n145 163.367
R2432 B.n1176 B.n1174 163.367
R2433 B.n1172 B.n147 163.367
R2434 B.n1168 B.n1166 163.367
R2435 B.n1164 B.n149 163.367
R2436 B.n1160 B.n1158 163.367
R2437 B.n1156 B.n151 163.367
R2438 B.n1152 B.n1150 163.367
R2439 B.n1148 B.n153 163.367
R2440 B.n1144 B.n1142 163.367
R2441 B.n1140 B.n155 163.367
R2442 B.n1136 B.n1134 163.367
R2443 B.n1132 B.n157 163.367
R2444 B.n1128 B.n1126 163.367
R2445 B.n1124 B.n159 163.367
R2446 B.n1120 B.n1118 163.367
R2447 B.n1115 B.n1114 163.367
R2448 B.n1112 B.n165 163.367
R2449 B.n1108 B.n1106 163.367
R2450 B.n1104 B.n167 163.367
R2451 B.n1099 B.n1097 163.367
R2452 B.n1095 B.n171 163.367
R2453 B.n1091 B.n1089 163.367
R2454 B.n1087 B.n173 163.367
R2455 B.n1083 B.n1081 163.367
R2456 B.n1079 B.n175 163.367
R2457 B.n1075 B.n1073 163.367
R2458 B.n1071 B.n177 163.367
R2459 B.n1067 B.n1065 163.367
R2460 B.n1063 B.n179 163.367
R2461 B.n1059 B.n1057 163.367
R2462 B.n1055 B.n181 163.367
R2463 B.n1051 B.n1049 163.367
R2464 B.n1047 B.n183 163.367
R2465 B.n1043 B.n1041 163.367
R2466 B.n1039 B.n185 163.367
R2467 B.n1035 B.n1033 163.367
R2468 B.n1031 B.n187 163.367
R2469 B.n1027 B.n1025 163.367
R2470 B.n1023 B.n189 163.367
R2471 B.n1019 B.n1017 163.367
R2472 B.n1015 B.n191 163.367
R2473 B.n1011 B.n1009 163.367
R2474 B.n1007 B.n193 163.367
R2475 B.n1003 B.n1001 163.367
R2476 B.n999 B.n195 163.367
R2477 B.n995 B.n993 163.367
R2478 B.n991 B.n197 163.367
R2479 B.n987 B.n985 163.367
R2480 B.n983 B.n199 163.367
R2481 B.n979 B.n977 163.367
R2482 B.n678 B.n335 163.367
R2483 B.n682 B.n335 163.367
R2484 B.n682 B.n329 163.367
R2485 B.n690 B.n329 163.367
R2486 B.n690 B.n327 163.367
R2487 B.n694 B.n327 163.367
R2488 B.n694 B.n320 163.367
R2489 B.n702 B.n320 163.367
R2490 B.n702 B.n318 163.367
R2491 B.n706 B.n318 163.367
R2492 B.n706 B.n313 163.367
R2493 B.n714 B.n313 163.367
R2494 B.n714 B.n311 163.367
R2495 B.n718 B.n311 163.367
R2496 B.n718 B.n305 163.367
R2497 B.n726 B.n305 163.367
R2498 B.n726 B.n303 163.367
R2499 B.n730 B.n303 163.367
R2500 B.n730 B.n297 163.367
R2501 B.n738 B.n297 163.367
R2502 B.n738 B.n295 163.367
R2503 B.n742 B.n295 163.367
R2504 B.n742 B.n288 163.367
R2505 B.n750 B.n288 163.367
R2506 B.n750 B.n286 163.367
R2507 B.n754 B.n286 163.367
R2508 B.n754 B.n281 163.367
R2509 B.n762 B.n281 163.367
R2510 B.n762 B.n279 163.367
R2511 B.n766 B.n279 163.367
R2512 B.n766 B.n273 163.367
R2513 B.n774 B.n273 163.367
R2514 B.n774 B.n271 163.367
R2515 B.n778 B.n271 163.367
R2516 B.n778 B.n264 163.367
R2517 B.n786 B.n264 163.367
R2518 B.n786 B.n262 163.367
R2519 B.n790 B.n262 163.367
R2520 B.n790 B.n257 163.367
R2521 B.n798 B.n257 163.367
R2522 B.n798 B.n255 163.367
R2523 B.n802 B.n255 163.367
R2524 B.n802 B.n249 163.367
R2525 B.n810 B.n249 163.367
R2526 B.n810 B.n247 163.367
R2527 B.n814 B.n247 163.367
R2528 B.n814 B.n241 163.367
R2529 B.n822 B.n241 163.367
R2530 B.n822 B.n239 163.367
R2531 B.n826 B.n239 163.367
R2532 B.n826 B.n233 163.367
R2533 B.n834 B.n233 163.367
R2534 B.n834 B.n231 163.367
R2535 B.n838 B.n231 163.367
R2536 B.n838 B.n225 163.367
R2537 B.n846 B.n225 163.367
R2538 B.n846 B.n223 163.367
R2539 B.n850 B.n223 163.367
R2540 B.n850 B.n217 163.367
R2541 B.n858 B.n217 163.367
R2542 B.n858 B.n215 163.367
R2543 B.n862 B.n215 163.367
R2544 B.n862 B.n209 163.367
R2545 B.n870 B.n209 163.367
R2546 B.n870 B.n207 163.367
R2547 B.n875 B.n207 163.367
R2548 B.n875 B.n201 163.367
R2549 B.n883 B.n201 163.367
R2550 B.n884 B.n883 163.367
R2551 B.n884 B.n5 163.367
R2552 B.n6 B.n5 163.367
R2553 B.n7 B.n6 163.367
R2554 B.n890 B.n7 163.367
R2555 B.n891 B.n890 163.367
R2556 B.n891 B.n13 163.367
R2557 B.n14 B.n13 163.367
R2558 B.n15 B.n14 163.367
R2559 B.n896 B.n15 163.367
R2560 B.n896 B.n20 163.367
R2561 B.n21 B.n20 163.367
R2562 B.n22 B.n21 163.367
R2563 B.n901 B.n22 163.367
R2564 B.n901 B.n27 163.367
R2565 B.n28 B.n27 163.367
R2566 B.n29 B.n28 163.367
R2567 B.n906 B.n29 163.367
R2568 B.n906 B.n34 163.367
R2569 B.n35 B.n34 163.367
R2570 B.n36 B.n35 163.367
R2571 B.n911 B.n36 163.367
R2572 B.n911 B.n41 163.367
R2573 B.n42 B.n41 163.367
R2574 B.n43 B.n42 163.367
R2575 B.n916 B.n43 163.367
R2576 B.n916 B.n48 163.367
R2577 B.n49 B.n48 163.367
R2578 B.n50 B.n49 163.367
R2579 B.n921 B.n50 163.367
R2580 B.n921 B.n55 163.367
R2581 B.n56 B.n55 163.367
R2582 B.n57 B.n56 163.367
R2583 B.n926 B.n57 163.367
R2584 B.n926 B.n62 163.367
R2585 B.n63 B.n62 163.367
R2586 B.n64 B.n63 163.367
R2587 B.n931 B.n64 163.367
R2588 B.n931 B.n69 163.367
R2589 B.n70 B.n69 163.367
R2590 B.n71 B.n70 163.367
R2591 B.n936 B.n71 163.367
R2592 B.n936 B.n76 163.367
R2593 B.n77 B.n76 163.367
R2594 B.n78 B.n77 163.367
R2595 B.n941 B.n78 163.367
R2596 B.n941 B.n83 163.367
R2597 B.n84 B.n83 163.367
R2598 B.n85 B.n84 163.367
R2599 B.n946 B.n85 163.367
R2600 B.n946 B.n90 163.367
R2601 B.n91 B.n90 163.367
R2602 B.n92 B.n91 163.367
R2603 B.n951 B.n92 163.367
R2604 B.n951 B.n97 163.367
R2605 B.n98 B.n97 163.367
R2606 B.n99 B.n98 163.367
R2607 B.n956 B.n99 163.367
R2608 B.n956 B.n104 163.367
R2609 B.n105 B.n104 163.367
R2610 B.n106 B.n105 163.367
R2611 B.n961 B.n106 163.367
R2612 B.n961 B.n111 163.367
R2613 B.n112 B.n111 163.367
R2614 B.n113 B.n112 163.367
R2615 B.n966 B.n113 163.367
R2616 B.n966 B.n118 163.367
R2617 B.n119 B.n118 163.367
R2618 B.n120 B.n119 163.367
R2619 B.n971 B.n120 163.367
R2620 B.n971 B.n125 163.367
R2621 B.n126 B.n125 163.367
R2622 B.n127 B.n126 163.367
R2623 B.n672 B.n670 163.367
R2624 B.n670 B.n669 163.367
R2625 B.n666 B.n665 163.367
R2626 B.n663 B.n343 163.367
R2627 B.n659 B.n657 163.367
R2628 B.n655 B.n345 163.367
R2629 B.n651 B.n649 163.367
R2630 B.n647 B.n347 163.367
R2631 B.n643 B.n641 163.367
R2632 B.n639 B.n349 163.367
R2633 B.n635 B.n633 163.367
R2634 B.n631 B.n351 163.367
R2635 B.n627 B.n625 163.367
R2636 B.n623 B.n353 163.367
R2637 B.n619 B.n617 163.367
R2638 B.n615 B.n355 163.367
R2639 B.n611 B.n609 163.367
R2640 B.n607 B.n357 163.367
R2641 B.n603 B.n601 163.367
R2642 B.n599 B.n359 163.367
R2643 B.n595 B.n593 163.367
R2644 B.n591 B.n361 163.367
R2645 B.n587 B.n585 163.367
R2646 B.n583 B.n363 163.367
R2647 B.n579 B.n577 163.367
R2648 B.n575 B.n365 163.367
R2649 B.n571 B.n569 163.367
R2650 B.n567 B.n367 163.367
R2651 B.n563 B.n561 163.367
R2652 B.n559 B.n369 163.367
R2653 B.n555 B.n553 163.367
R2654 B.n551 B.n371 163.367
R2655 B.n547 B.n545 163.367
R2656 B.n543 B.n376 163.367
R2657 B.n539 B.n537 163.367
R2658 B.n535 B.n378 163.367
R2659 B.n530 B.n528 163.367
R2660 B.n526 B.n382 163.367
R2661 B.n522 B.n520 163.367
R2662 B.n518 B.n384 163.367
R2663 B.n514 B.n512 163.367
R2664 B.n510 B.n386 163.367
R2665 B.n506 B.n504 163.367
R2666 B.n502 B.n388 163.367
R2667 B.n498 B.n496 163.367
R2668 B.n494 B.n390 163.367
R2669 B.n490 B.n488 163.367
R2670 B.n486 B.n392 163.367
R2671 B.n482 B.n480 163.367
R2672 B.n478 B.n394 163.367
R2673 B.n474 B.n472 163.367
R2674 B.n470 B.n396 163.367
R2675 B.n466 B.n464 163.367
R2676 B.n462 B.n398 163.367
R2677 B.n458 B.n456 163.367
R2678 B.n454 B.n400 163.367
R2679 B.n450 B.n448 163.367
R2680 B.n446 B.n402 163.367
R2681 B.n442 B.n440 163.367
R2682 B.n438 B.n404 163.367
R2683 B.n434 B.n432 163.367
R2684 B.n430 B.n406 163.367
R2685 B.n426 B.n424 163.367
R2686 B.n422 B.n408 163.367
R2687 B.n418 B.n416 163.367
R2688 B.n414 B.n411 163.367
R2689 B.n676 B.n333 163.367
R2690 B.n684 B.n333 163.367
R2691 B.n684 B.n331 163.367
R2692 B.n688 B.n331 163.367
R2693 B.n688 B.n325 163.367
R2694 B.n696 B.n325 163.367
R2695 B.n696 B.n323 163.367
R2696 B.n700 B.n323 163.367
R2697 B.n700 B.n317 163.367
R2698 B.n708 B.n317 163.367
R2699 B.n708 B.n315 163.367
R2700 B.n712 B.n315 163.367
R2701 B.n712 B.n309 163.367
R2702 B.n720 B.n309 163.367
R2703 B.n720 B.n307 163.367
R2704 B.n724 B.n307 163.367
R2705 B.n724 B.n301 163.367
R2706 B.n732 B.n301 163.367
R2707 B.n732 B.n299 163.367
R2708 B.n736 B.n299 163.367
R2709 B.n736 B.n293 163.367
R2710 B.n744 B.n293 163.367
R2711 B.n744 B.n291 163.367
R2712 B.n748 B.n291 163.367
R2713 B.n748 B.n285 163.367
R2714 B.n756 B.n285 163.367
R2715 B.n756 B.n283 163.367
R2716 B.n760 B.n283 163.367
R2717 B.n760 B.n277 163.367
R2718 B.n768 B.n277 163.367
R2719 B.n768 B.n275 163.367
R2720 B.n772 B.n275 163.367
R2721 B.n772 B.n269 163.367
R2722 B.n780 B.n269 163.367
R2723 B.n780 B.n267 163.367
R2724 B.n784 B.n267 163.367
R2725 B.n784 B.n261 163.367
R2726 B.n792 B.n261 163.367
R2727 B.n792 B.n259 163.367
R2728 B.n796 B.n259 163.367
R2729 B.n796 B.n253 163.367
R2730 B.n804 B.n253 163.367
R2731 B.n804 B.n251 163.367
R2732 B.n808 B.n251 163.367
R2733 B.n808 B.n245 163.367
R2734 B.n816 B.n245 163.367
R2735 B.n816 B.n243 163.367
R2736 B.n820 B.n243 163.367
R2737 B.n820 B.n237 163.367
R2738 B.n828 B.n237 163.367
R2739 B.n828 B.n235 163.367
R2740 B.n832 B.n235 163.367
R2741 B.n832 B.n229 163.367
R2742 B.n840 B.n229 163.367
R2743 B.n840 B.n227 163.367
R2744 B.n844 B.n227 163.367
R2745 B.n844 B.n221 163.367
R2746 B.n852 B.n221 163.367
R2747 B.n852 B.n219 163.367
R2748 B.n856 B.n219 163.367
R2749 B.n856 B.n213 163.367
R2750 B.n864 B.n213 163.367
R2751 B.n864 B.n211 163.367
R2752 B.n868 B.n211 163.367
R2753 B.n868 B.n205 163.367
R2754 B.n877 B.n205 163.367
R2755 B.n877 B.n203 163.367
R2756 B.n881 B.n203 163.367
R2757 B.n881 B.n3 163.367
R2758 B.n1385 B.n3 163.367
R2759 B.n1381 B.n2 163.367
R2760 B.n1381 B.n1380 163.367
R2761 B.n1380 B.n9 163.367
R2762 B.n1376 B.n9 163.367
R2763 B.n1376 B.n11 163.367
R2764 B.n1372 B.n11 163.367
R2765 B.n1372 B.n17 163.367
R2766 B.n1368 B.n17 163.367
R2767 B.n1368 B.n19 163.367
R2768 B.n1364 B.n19 163.367
R2769 B.n1364 B.n24 163.367
R2770 B.n1360 B.n24 163.367
R2771 B.n1360 B.n26 163.367
R2772 B.n1356 B.n26 163.367
R2773 B.n1356 B.n31 163.367
R2774 B.n1352 B.n31 163.367
R2775 B.n1352 B.n33 163.367
R2776 B.n1348 B.n33 163.367
R2777 B.n1348 B.n38 163.367
R2778 B.n1344 B.n38 163.367
R2779 B.n1344 B.n40 163.367
R2780 B.n1340 B.n40 163.367
R2781 B.n1340 B.n45 163.367
R2782 B.n1336 B.n45 163.367
R2783 B.n1336 B.n47 163.367
R2784 B.n1332 B.n47 163.367
R2785 B.n1332 B.n52 163.367
R2786 B.n1328 B.n52 163.367
R2787 B.n1328 B.n54 163.367
R2788 B.n1324 B.n54 163.367
R2789 B.n1324 B.n59 163.367
R2790 B.n1320 B.n59 163.367
R2791 B.n1320 B.n61 163.367
R2792 B.n1316 B.n61 163.367
R2793 B.n1316 B.n66 163.367
R2794 B.n1312 B.n66 163.367
R2795 B.n1312 B.n68 163.367
R2796 B.n1308 B.n68 163.367
R2797 B.n1308 B.n73 163.367
R2798 B.n1304 B.n73 163.367
R2799 B.n1304 B.n75 163.367
R2800 B.n1300 B.n75 163.367
R2801 B.n1300 B.n80 163.367
R2802 B.n1296 B.n80 163.367
R2803 B.n1296 B.n82 163.367
R2804 B.n1292 B.n82 163.367
R2805 B.n1292 B.n87 163.367
R2806 B.n1288 B.n87 163.367
R2807 B.n1288 B.n89 163.367
R2808 B.n1284 B.n89 163.367
R2809 B.n1284 B.n94 163.367
R2810 B.n1280 B.n94 163.367
R2811 B.n1280 B.n96 163.367
R2812 B.n1276 B.n96 163.367
R2813 B.n1276 B.n101 163.367
R2814 B.n1272 B.n101 163.367
R2815 B.n1272 B.n103 163.367
R2816 B.n1268 B.n103 163.367
R2817 B.n1268 B.n108 163.367
R2818 B.n1264 B.n108 163.367
R2819 B.n1264 B.n110 163.367
R2820 B.n1260 B.n110 163.367
R2821 B.n1260 B.n115 163.367
R2822 B.n1256 B.n115 163.367
R2823 B.n1256 B.n117 163.367
R2824 B.n1252 B.n117 163.367
R2825 B.n1252 B.n122 163.367
R2826 B.n1248 B.n122 163.367
R2827 B.n1248 B.n124 163.367
R2828 B.n1244 B.n124 163.367
R2829 B.n161 B.n160 82.2308
R2830 B.n169 B.n168 82.2308
R2831 B.n380 B.n379 82.2308
R2832 B.n373 B.n372 82.2308
R2833 B.n1239 B.n129 71.676
R2834 B.n1238 B.n1237 71.676
R2835 B.n1231 B.n131 71.676
R2836 B.n1230 B.n1229 71.676
R2837 B.n1223 B.n133 71.676
R2838 B.n1222 B.n1221 71.676
R2839 B.n1215 B.n135 71.676
R2840 B.n1214 B.n1213 71.676
R2841 B.n1207 B.n137 71.676
R2842 B.n1206 B.n1205 71.676
R2843 B.n1199 B.n139 71.676
R2844 B.n1198 B.n1197 71.676
R2845 B.n1191 B.n141 71.676
R2846 B.n1190 B.n1189 71.676
R2847 B.n1183 B.n143 71.676
R2848 B.n1182 B.n1181 71.676
R2849 B.n1175 B.n145 71.676
R2850 B.n1174 B.n1173 71.676
R2851 B.n1167 B.n147 71.676
R2852 B.n1166 B.n1165 71.676
R2853 B.n1159 B.n149 71.676
R2854 B.n1158 B.n1157 71.676
R2855 B.n1151 B.n151 71.676
R2856 B.n1150 B.n1149 71.676
R2857 B.n1143 B.n153 71.676
R2858 B.n1142 B.n1141 71.676
R2859 B.n1135 B.n155 71.676
R2860 B.n1134 B.n1133 71.676
R2861 B.n1127 B.n157 71.676
R2862 B.n1126 B.n1125 71.676
R2863 B.n1119 B.n159 71.676
R2864 B.n1118 B.n163 71.676
R2865 B.n1114 B.n1113 71.676
R2866 B.n1107 B.n165 71.676
R2867 B.n1106 B.n1105 71.676
R2868 B.n1098 B.n167 71.676
R2869 B.n1097 B.n1096 71.676
R2870 B.n1090 B.n171 71.676
R2871 B.n1089 B.n1088 71.676
R2872 B.n1082 B.n173 71.676
R2873 B.n1081 B.n1080 71.676
R2874 B.n1074 B.n175 71.676
R2875 B.n1073 B.n1072 71.676
R2876 B.n1066 B.n177 71.676
R2877 B.n1065 B.n1064 71.676
R2878 B.n1058 B.n179 71.676
R2879 B.n1057 B.n1056 71.676
R2880 B.n1050 B.n181 71.676
R2881 B.n1049 B.n1048 71.676
R2882 B.n1042 B.n183 71.676
R2883 B.n1041 B.n1040 71.676
R2884 B.n1034 B.n185 71.676
R2885 B.n1033 B.n1032 71.676
R2886 B.n1026 B.n187 71.676
R2887 B.n1025 B.n1024 71.676
R2888 B.n1018 B.n189 71.676
R2889 B.n1017 B.n1016 71.676
R2890 B.n1010 B.n191 71.676
R2891 B.n1009 B.n1008 71.676
R2892 B.n1002 B.n193 71.676
R2893 B.n1001 B.n1000 71.676
R2894 B.n994 B.n195 71.676
R2895 B.n993 B.n992 71.676
R2896 B.n986 B.n197 71.676
R2897 B.n985 B.n984 71.676
R2898 B.n978 B.n199 71.676
R2899 B.n979 B.n978 71.676
R2900 B.n984 B.n983 71.676
R2901 B.n987 B.n986 71.676
R2902 B.n992 B.n991 71.676
R2903 B.n995 B.n994 71.676
R2904 B.n1000 B.n999 71.676
R2905 B.n1003 B.n1002 71.676
R2906 B.n1008 B.n1007 71.676
R2907 B.n1011 B.n1010 71.676
R2908 B.n1016 B.n1015 71.676
R2909 B.n1019 B.n1018 71.676
R2910 B.n1024 B.n1023 71.676
R2911 B.n1027 B.n1026 71.676
R2912 B.n1032 B.n1031 71.676
R2913 B.n1035 B.n1034 71.676
R2914 B.n1040 B.n1039 71.676
R2915 B.n1043 B.n1042 71.676
R2916 B.n1048 B.n1047 71.676
R2917 B.n1051 B.n1050 71.676
R2918 B.n1056 B.n1055 71.676
R2919 B.n1059 B.n1058 71.676
R2920 B.n1064 B.n1063 71.676
R2921 B.n1067 B.n1066 71.676
R2922 B.n1072 B.n1071 71.676
R2923 B.n1075 B.n1074 71.676
R2924 B.n1080 B.n1079 71.676
R2925 B.n1083 B.n1082 71.676
R2926 B.n1088 B.n1087 71.676
R2927 B.n1091 B.n1090 71.676
R2928 B.n1096 B.n1095 71.676
R2929 B.n1099 B.n1098 71.676
R2930 B.n1105 B.n1104 71.676
R2931 B.n1108 B.n1107 71.676
R2932 B.n1113 B.n1112 71.676
R2933 B.n1115 B.n163 71.676
R2934 B.n1120 B.n1119 71.676
R2935 B.n1125 B.n1124 71.676
R2936 B.n1128 B.n1127 71.676
R2937 B.n1133 B.n1132 71.676
R2938 B.n1136 B.n1135 71.676
R2939 B.n1141 B.n1140 71.676
R2940 B.n1144 B.n1143 71.676
R2941 B.n1149 B.n1148 71.676
R2942 B.n1152 B.n1151 71.676
R2943 B.n1157 B.n1156 71.676
R2944 B.n1160 B.n1159 71.676
R2945 B.n1165 B.n1164 71.676
R2946 B.n1168 B.n1167 71.676
R2947 B.n1173 B.n1172 71.676
R2948 B.n1176 B.n1175 71.676
R2949 B.n1181 B.n1180 71.676
R2950 B.n1184 B.n1183 71.676
R2951 B.n1189 B.n1188 71.676
R2952 B.n1192 B.n1191 71.676
R2953 B.n1197 B.n1196 71.676
R2954 B.n1200 B.n1199 71.676
R2955 B.n1205 B.n1204 71.676
R2956 B.n1208 B.n1207 71.676
R2957 B.n1213 B.n1212 71.676
R2958 B.n1216 B.n1215 71.676
R2959 B.n1221 B.n1220 71.676
R2960 B.n1224 B.n1223 71.676
R2961 B.n1229 B.n1228 71.676
R2962 B.n1232 B.n1231 71.676
R2963 B.n1237 B.n1236 71.676
R2964 B.n1240 B.n1239 71.676
R2965 B.n671 B.n339 71.676
R2966 B.n669 B.n341 71.676
R2967 B.n665 B.n664 71.676
R2968 B.n658 B.n343 71.676
R2969 B.n657 B.n656 71.676
R2970 B.n650 B.n345 71.676
R2971 B.n649 B.n648 71.676
R2972 B.n642 B.n347 71.676
R2973 B.n641 B.n640 71.676
R2974 B.n634 B.n349 71.676
R2975 B.n633 B.n632 71.676
R2976 B.n626 B.n351 71.676
R2977 B.n625 B.n624 71.676
R2978 B.n618 B.n353 71.676
R2979 B.n617 B.n616 71.676
R2980 B.n610 B.n355 71.676
R2981 B.n609 B.n608 71.676
R2982 B.n602 B.n357 71.676
R2983 B.n601 B.n600 71.676
R2984 B.n594 B.n359 71.676
R2985 B.n593 B.n592 71.676
R2986 B.n586 B.n361 71.676
R2987 B.n585 B.n584 71.676
R2988 B.n578 B.n363 71.676
R2989 B.n577 B.n576 71.676
R2990 B.n570 B.n365 71.676
R2991 B.n569 B.n568 71.676
R2992 B.n562 B.n367 71.676
R2993 B.n561 B.n560 71.676
R2994 B.n554 B.n369 71.676
R2995 B.n553 B.n552 71.676
R2996 B.n546 B.n371 71.676
R2997 B.n545 B.n544 71.676
R2998 B.n538 B.n376 71.676
R2999 B.n537 B.n536 71.676
R3000 B.n529 B.n378 71.676
R3001 B.n528 B.n527 71.676
R3002 B.n521 B.n382 71.676
R3003 B.n520 B.n519 71.676
R3004 B.n513 B.n384 71.676
R3005 B.n512 B.n511 71.676
R3006 B.n505 B.n386 71.676
R3007 B.n504 B.n503 71.676
R3008 B.n497 B.n388 71.676
R3009 B.n496 B.n495 71.676
R3010 B.n489 B.n390 71.676
R3011 B.n488 B.n487 71.676
R3012 B.n481 B.n392 71.676
R3013 B.n480 B.n479 71.676
R3014 B.n473 B.n394 71.676
R3015 B.n472 B.n471 71.676
R3016 B.n465 B.n396 71.676
R3017 B.n464 B.n463 71.676
R3018 B.n457 B.n398 71.676
R3019 B.n456 B.n455 71.676
R3020 B.n449 B.n400 71.676
R3021 B.n448 B.n447 71.676
R3022 B.n441 B.n402 71.676
R3023 B.n440 B.n439 71.676
R3024 B.n433 B.n404 71.676
R3025 B.n432 B.n431 71.676
R3026 B.n425 B.n406 71.676
R3027 B.n424 B.n423 71.676
R3028 B.n417 B.n408 71.676
R3029 B.n416 B.n415 71.676
R3030 B.n411 B.n410 71.676
R3031 B.n672 B.n671 71.676
R3032 B.n666 B.n341 71.676
R3033 B.n664 B.n663 71.676
R3034 B.n659 B.n658 71.676
R3035 B.n656 B.n655 71.676
R3036 B.n651 B.n650 71.676
R3037 B.n648 B.n647 71.676
R3038 B.n643 B.n642 71.676
R3039 B.n640 B.n639 71.676
R3040 B.n635 B.n634 71.676
R3041 B.n632 B.n631 71.676
R3042 B.n627 B.n626 71.676
R3043 B.n624 B.n623 71.676
R3044 B.n619 B.n618 71.676
R3045 B.n616 B.n615 71.676
R3046 B.n611 B.n610 71.676
R3047 B.n608 B.n607 71.676
R3048 B.n603 B.n602 71.676
R3049 B.n600 B.n599 71.676
R3050 B.n595 B.n594 71.676
R3051 B.n592 B.n591 71.676
R3052 B.n587 B.n586 71.676
R3053 B.n584 B.n583 71.676
R3054 B.n579 B.n578 71.676
R3055 B.n576 B.n575 71.676
R3056 B.n571 B.n570 71.676
R3057 B.n568 B.n567 71.676
R3058 B.n563 B.n562 71.676
R3059 B.n560 B.n559 71.676
R3060 B.n555 B.n554 71.676
R3061 B.n552 B.n551 71.676
R3062 B.n547 B.n546 71.676
R3063 B.n544 B.n543 71.676
R3064 B.n539 B.n538 71.676
R3065 B.n536 B.n535 71.676
R3066 B.n530 B.n529 71.676
R3067 B.n527 B.n526 71.676
R3068 B.n522 B.n521 71.676
R3069 B.n519 B.n518 71.676
R3070 B.n514 B.n513 71.676
R3071 B.n511 B.n510 71.676
R3072 B.n506 B.n505 71.676
R3073 B.n503 B.n502 71.676
R3074 B.n498 B.n497 71.676
R3075 B.n495 B.n494 71.676
R3076 B.n490 B.n489 71.676
R3077 B.n487 B.n486 71.676
R3078 B.n482 B.n481 71.676
R3079 B.n479 B.n478 71.676
R3080 B.n474 B.n473 71.676
R3081 B.n471 B.n470 71.676
R3082 B.n466 B.n465 71.676
R3083 B.n463 B.n462 71.676
R3084 B.n458 B.n457 71.676
R3085 B.n455 B.n454 71.676
R3086 B.n450 B.n449 71.676
R3087 B.n447 B.n446 71.676
R3088 B.n442 B.n441 71.676
R3089 B.n439 B.n438 71.676
R3090 B.n434 B.n433 71.676
R3091 B.n431 B.n430 71.676
R3092 B.n426 B.n425 71.676
R3093 B.n423 B.n422 71.676
R3094 B.n418 B.n417 71.676
R3095 B.n415 B.n414 71.676
R3096 B.n410 B.n337 71.676
R3097 B.n1386 B.n1385 71.676
R3098 B.n1386 B.n2 71.676
R3099 B.n162 B.n161 59.5399
R3100 B.n1101 B.n169 59.5399
R3101 B.n533 B.n380 59.5399
R3102 B.n374 B.n373 59.5399
R3103 B.n677 B.n338 55.103
R3104 B.n1245 B.n128 55.103
R3105 B.n675 B.n674 33.5615
R3106 B.n679 B.n336 33.5615
R3107 B.n976 B.n975 33.5615
R3108 B.n1243 B.n1242 33.5615
R3109 B.n677 B.n334 30.9672
R3110 B.n683 B.n334 30.9672
R3111 B.n683 B.n330 30.9672
R3112 B.n689 B.n330 30.9672
R3113 B.n689 B.n326 30.9672
R3114 B.n695 B.n326 30.9672
R3115 B.n695 B.n321 30.9672
R3116 B.n701 B.n321 30.9672
R3117 B.n701 B.n322 30.9672
R3118 B.n707 B.n314 30.9672
R3119 B.n713 B.n314 30.9672
R3120 B.n713 B.n310 30.9672
R3121 B.n719 B.n310 30.9672
R3122 B.n719 B.n306 30.9672
R3123 B.n725 B.n306 30.9672
R3124 B.n725 B.n302 30.9672
R3125 B.n731 B.n302 30.9672
R3126 B.n731 B.n298 30.9672
R3127 B.n737 B.n298 30.9672
R3128 B.n737 B.n294 30.9672
R3129 B.n743 B.n294 30.9672
R3130 B.n743 B.n289 30.9672
R3131 B.n749 B.n289 30.9672
R3132 B.n749 B.n290 30.9672
R3133 B.n755 B.n282 30.9672
R3134 B.n761 B.n282 30.9672
R3135 B.n761 B.n278 30.9672
R3136 B.n767 B.n278 30.9672
R3137 B.n767 B.n274 30.9672
R3138 B.n773 B.n274 30.9672
R3139 B.n773 B.n270 30.9672
R3140 B.n779 B.n270 30.9672
R3141 B.n779 B.n265 30.9672
R3142 B.n785 B.n265 30.9672
R3143 B.n785 B.n266 30.9672
R3144 B.n791 B.n258 30.9672
R3145 B.n797 B.n258 30.9672
R3146 B.n797 B.n254 30.9672
R3147 B.n803 B.n254 30.9672
R3148 B.n803 B.n250 30.9672
R3149 B.n809 B.n250 30.9672
R3150 B.n809 B.n246 30.9672
R3151 B.n815 B.n246 30.9672
R3152 B.n815 B.n242 30.9672
R3153 B.n821 B.n242 30.9672
R3154 B.n821 B.n238 30.9672
R3155 B.n827 B.n238 30.9672
R3156 B.n833 B.n234 30.9672
R3157 B.n833 B.n230 30.9672
R3158 B.n839 B.n230 30.9672
R3159 B.n839 B.n226 30.9672
R3160 B.n845 B.n226 30.9672
R3161 B.n845 B.n222 30.9672
R3162 B.n851 B.n222 30.9672
R3163 B.n851 B.n218 30.9672
R3164 B.n857 B.n218 30.9672
R3165 B.n857 B.n214 30.9672
R3166 B.n863 B.n214 30.9672
R3167 B.n869 B.n210 30.9672
R3168 B.n869 B.n206 30.9672
R3169 B.n876 B.n206 30.9672
R3170 B.n876 B.n202 30.9672
R3171 B.n882 B.n202 30.9672
R3172 B.n882 B.n4 30.9672
R3173 B.n1384 B.n4 30.9672
R3174 B.n1384 B.n1383 30.9672
R3175 B.n1383 B.n1382 30.9672
R3176 B.n1382 B.n8 30.9672
R3177 B.n12 B.n8 30.9672
R3178 B.n1375 B.n12 30.9672
R3179 B.n1375 B.n1374 30.9672
R3180 B.n1374 B.n1373 30.9672
R3181 B.n1373 B.n16 30.9672
R3182 B.n1367 B.n1366 30.9672
R3183 B.n1366 B.n1365 30.9672
R3184 B.n1365 B.n23 30.9672
R3185 B.n1359 B.n23 30.9672
R3186 B.n1359 B.n1358 30.9672
R3187 B.n1358 B.n1357 30.9672
R3188 B.n1357 B.n30 30.9672
R3189 B.n1351 B.n30 30.9672
R3190 B.n1351 B.n1350 30.9672
R3191 B.n1350 B.n1349 30.9672
R3192 B.n1349 B.n37 30.9672
R3193 B.n1343 B.n1342 30.9672
R3194 B.n1342 B.n1341 30.9672
R3195 B.n1341 B.n44 30.9672
R3196 B.n1335 B.n44 30.9672
R3197 B.n1335 B.n1334 30.9672
R3198 B.n1334 B.n1333 30.9672
R3199 B.n1333 B.n51 30.9672
R3200 B.n1327 B.n51 30.9672
R3201 B.n1327 B.n1326 30.9672
R3202 B.n1326 B.n1325 30.9672
R3203 B.n1325 B.n58 30.9672
R3204 B.n1319 B.n58 30.9672
R3205 B.n1318 B.n1317 30.9672
R3206 B.n1317 B.n65 30.9672
R3207 B.n1311 B.n65 30.9672
R3208 B.n1311 B.n1310 30.9672
R3209 B.n1310 B.n1309 30.9672
R3210 B.n1309 B.n72 30.9672
R3211 B.n1303 B.n72 30.9672
R3212 B.n1303 B.n1302 30.9672
R3213 B.n1302 B.n1301 30.9672
R3214 B.n1301 B.n79 30.9672
R3215 B.n1295 B.n79 30.9672
R3216 B.n1294 B.n1293 30.9672
R3217 B.n1293 B.n86 30.9672
R3218 B.n1287 B.n86 30.9672
R3219 B.n1287 B.n1286 30.9672
R3220 B.n1286 B.n1285 30.9672
R3221 B.n1285 B.n93 30.9672
R3222 B.n1279 B.n93 30.9672
R3223 B.n1279 B.n1278 30.9672
R3224 B.n1278 B.n1277 30.9672
R3225 B.n1277 B.n100 30.9672
R3226 B.n1271 B.n100 30.9672
R3227 B.n1271 B.n1270 30.9672
R3228 B.n1270 B.n1269 30.9672
R3229 B.n1269 B.n107 30.9672
R3230 B.n1263 B.n107 30.9672
R3231 B.n1262 B.n1261 30.9672
R3232 B.n1261 B.n114 30.9672
R3233 B.n1255 B.n114 30.9672
R3234 B.n1255 B.n1254 30.9672
R3235 B.n1254 B.n1253 30.9672
R3236 B.n1253 B.n121 30.9672
R3237 B.n1247 B.n121 30.9672
R3238 B.n1247 B.n1246 30.9672
R3239 B.n1246 B.n1245 30.9672
R3240 B.t6 B.n234 25.0471
R3241 B.t1 B.n37 25.0471
R3242 B.n755 B.t4 23.2255
R3243 B.n1295 B.t3 23.2255
R3244 B.n266 B.t2 22.3147
R3245 B.t0 B.n1318 22.3147
R3246 B.n863 B.t5 20.4932
R3247 B.n1367 B.t7 20.4932
R3248 B B.n1387 18.0485
R3249 B.n322 B.t9 17.7608
R3250 B.t13 B.n1262 17.7608
R3251 B.n707 B.t9 13.2069
R3252 B.n1263 B.t13 13.2069
R3253 B.n675 B.n332 10.6151
R3254 B.n685 B.n332 10.6151
R3255 B.n686 B.n685 10.6151
R3256 B.n687 B.n686 10.6151
R3257 B.n687 B.n324 10.6151
R3258 B.n697 B.n324 10.6151
R3259 B.n698 B.n697 10.6151
R3260 B.n699 B.n698 10.6151
R3261 B.n699 B.n316 10.6151
R3262 B.n709 B.n316 10.6151
R3263 B.n710 B.n709 10.6151
R3264 B.n711 B.n710 10.6151
R3265 B.n711 B.n308 10.6151
R3266 B.n721 B.n308 10.6151
R3267 B.n722 B.n721 10.6151
R3268 B.n723 B.n722 10.6151
R3269 B.n723 B.n300 10.6151
R3270 B.n733 B.n300 10.6151
R3271 B.n734 B.n733 10.6151
R3272 B.n735 B.n734 10.6151
R3273 B.n735 B.n292 10.6151
R3274 B.n745 B.n292 10.6151
R3275 B.n746 B.n745 10.6151
R3276 B.n747 B.n746 10.6151
R3277 B.n747 B.n284 10.6151
R3278 B.n757 B.n284 10.6151
R3279 B.n758 B.n757 10.6151
R3280 B.n759 B.n758 10.6151
R3281 B.n759 B.n276 10.6151
R3282 B.n769 B.n276 10.6151
R3283 B.n770 B.n769 10.6151
R3284 B.n771 B.n770 10.6151
R3285 B.n771 B.n268 10.6151
R3286 B.n781 B.n268 10.6151
R3287 B.n782 B.n781 10.6151
R3288 B.n783 B.n782 10.6151
R3289 B.n783 B.n260 10.6151
R3290 B.n793 B.n260 10.6151
R3291 B.n794 B.n793 10.6151
R3292 B.n795 B.n794 10.6151
R3293 B.n795 B.n252 10.6151
R3294 B.n805 B.n252 10.6151
R3295 B.n806 B.n805 10.6151
R3296 B.n807 B.n806 10.6151
R3297 B.n807 B.n244 10.6151
R3298 B.n817 B.n244 10.6151
R3299 B.n818 B.n817 10.6151
R3300 B.n819 B.n818 10.6151
R3301 B.n819 B.n236 10.6151
R3302 B.n829 B.n236 10.6151
R3303 B.n830 B.n829 10.6151
R3304 B.n831 B.n830 10.6151
R3305 B.n831 B.n228 10.6151
R3306 B.n841 B.n228 10.6151
R3307 B.n842 B.n841 10.6151
R3308 B.n843 B.n842 10.6151
R3309 B.n843 B.n220 10.6151
R3310 B.n853 B.n220 10.6151
R3311 B.n854 B.n853 10.6151
R3312 B.n855 B.n854 10.6151
R3313 B.n855 B.n212 10.6151
R3314 B.n865 B.n212 10.6151
R3315 B.n866 B.n865 10.6151
R3316 B.n867 B.n866 10.6151
R3317 B.n867 B.n204 10.6151
R3318 B.n878 B.n204 10.6151
R3319 B.n879 B.n878 10.6151
R3320 B.n880 B.n879 10.6151
R3321 B.n880 B.n0 10.6151
R3322 B.n674 B.n673 10.6151
R3323 B.n673 B.n340 10.6151
R3324 B.n668 B.n340 10.6151
R3325 B.n668 B.n667 10.6151
R3326 B.n667 B.n342 10.6151
R3327 B.n662 B.n342 10.6151
R3328 B.n662 B.n661 10.6151
R3329 B.n661 B.n660 10.6151
R3330 B.n660 B.n344 10.6151
R3331 B.n654 B.n344 10.6151
R3332 B.n654 B.n653 10.6151
R3333 B.n653 B.n652 10.6151
R3334 B.n652 B.n346 10.6151
R3335 B.n646 B.n346 10.6151
R3336 B.n646 B.n645 10.6151
R3337 B.n645 B.n644 10.6151
R3338 B.n644 B.n348 10.6151
R3339 B.n638 B.n348 10.6151
R3340 B.n638 B.n637 10.6151
R3341 B.n637 B.n636 10.6151
R3342 B.n636 B.n350 10.6151
R3343 B.n630 B.n350 10.6151
R3344 B.n630 B.n629 10.6151
R3345 B.n629 B.n628 10.6151
R3346 B.n628 B.n352 10.6151
R3347 B.n622 B.n352 10.6151
R3348 B.n622 B.n621 10.6151
R3349 B.n621 B.n620 10.6151
R3350 B.n620 B.n354 10.6151
R3351 B.n614 B.n354 10.6151
R3352 B.n614 B.n613 10.6151
R3353 B.n613 B.n612 10.6151
R3354 B.n612 B.n356 10.6151
R3355 B.n606 B.n356 10.6151
R3356 B.n606 B.n605 10.6151
R3357 B.n605 B.n604 10.6151
R3358 B.n604 B.n358 10.6151
R3359 B.n598 B.n358 10.6151
R3360 B.n598 B.n597 10.6151
R3361 B.n597 B.n596 10.6151
R3362 B.n596 B.n360 10.6151
R3363 B.n590 B.n360 10.6151
R3364 B.n590 B.n589 10.6151
R3365 B.n589 B.n588 10.6151
R3366 B.n588 B.n362 10.6151
R3367 B.n582 B.n362 10.6151
R3368 B.n582 B.n581 10.6151
R3369 B.n581 B.n580 10.6151
R3370 B.n580 B.n364 10.6151
R3371 B.n574 B.n364 10.6151
R3372 B.n574 B.n573 10.6151
R3373 B.n573 B.n572 10.6151
R3374 B.n572 B.n366 10.6151
R3375 B.n566 B.n366 10.6151
R3376 B.n566 B.n565 10.6151
R3377 B.n565 B.n564 10.6151
R3378 B.n564 B.n368 10.6151
R3379 B.n558 B.n368 10.6151
R3380 B.n558 B.n557 10.6151
R3381 B.n557 B.n556 10.6151
R3382 B.n556 B.n370 10.6151
R3383 B.n550 B.n549 10.6151
R3384 B.n549 B.n548 10.6151
R3385 B.n548 B.n375 10.6151
R3386 B.n542 B.n375 10.6151
R3387 B.n542 B.n541 10.6151
R3388 B.n541 B.n540 10.6151
R3389 B.n540 B.n377 10.6151
R3390 B.n534 B.n377 10.6151
R3391 B.n532 B.n531 10.6151
R3392 B.n531 B.n381 10.6151
R3393 B.n525 B.n381 10.6151
R3394 B.n525 B.n524 10.6151
R3395 B.n524 B.n523 10.6151
R3396 B.n523 B.n383 10.6151
R3397 B.n517 B.n383 10.6151
R3398 B.n517 B.n516 10.6151
R3399 B.n516 B.n515 10.6151
R3400 B.n515 B.n385 10.6151
R3401 B.n509 B.n385 10.6151
R3402 B.n509 B.n508 10.6151
R3403 B.n508 B.n507 10.6151
R3404 B.n507 B.n387 10.6151
R3405 B.n501 B.n387 10.6151
R3406 B.n501 B.n500 10.6151
R3407 B.n500 B.n499 10.6151
R3408 B.n499 B.n389 10.6151
R3409 B.n493 B.n389 10.6151
R3410 B.n493 B.n492 10.6151
R3411 B.n492 B.n491 10.6151
R3412 B.n491 B.n391 10.6151
R3413 B.n485 B.n391 10.6151
R3414 B.n485 B.n484 10.6151
R3415 B.n484 B.n483 10.6151
R3416 B.n483 B.n393 10.6151
R3417 B.n477 B.n393 10.6151
R3418 B.n477 B.n476 10.6151
R3419 B.n476 B.n475 10.6151
R3420 B.n475 B.n395 10.6151
R3421 B.n469 B.n395 10.6151
R3422 B.n469 B.n468 10.6151
R3423 B.n468 B.n467 10.6151
R3424 B.n467 B.n397 10.6151
R3425 B.n461 B.n397 10.6151
R3426 B.n461 B.n460 10.6151
R3427 B.n460 B.n459 10.6151
R3428 B.n459 B.n399 10.6151
R3429 B.n453 B.n399 10.6151
R3430 B.n453 B.n452 10.6151
R3431 B.n452 B.n451 10.6151
R3432 B.n451 B.n401 10.6151
R3433 B.n445 B.n401 10.6151
R3434 B.n445 B.n444 10.6151
R3435 B.n444 B.n443 10.6151
R3436 B.n443 B.n403 10.6151
R3437 B.n437 B.n403 10.6151
R3438 B.n437 B.n436 10.6151
R3439 B.n436 B.n435 10.6151
R3440 B.n435 B.n405 10.6151
R3441 B.n429 B.n405 10.6151
R3442 B.n429 B.n428 10.6151
R3443 B.n428 B.n427 10.6151
R3444 B.n427 B.n407 10.6151
R3445 B.n421 B.n407 10.6151
R3446 B.n421 B.n420 10.6151
R3447 B.n420 B.n419 10.6151
R3448 B.n419 B.n409 10.6151
R3449 B.n413 B.n409 10.6151
R3450 B.n413 B.n412 10.6151
R3451 B.n412 B.n336 10.6151
R3452 B.n680 B.n679 10.6151
R3453 B.n681 B.n680 10.6151
R3454 B.n681 B.n328 10.6151
R3455 B.n691 B.n328 10.6151
R3456 B.n692 B.n691 10.6151
R3457 B.n693 B.n692 10.6151
R3458 B.n693 B.n319 10.6151
R3459 B.n703 B.n319 10.6151
R3460 B.n704 B.n703 10.6151
R3461 B.n705 B.n704 10.6151
R3462 B.n705 B.n312 10.6151
R3463 B.n715 B.n312 10.6151
R3464 B.n716 B.n715 10.6151
R3465 B.n717 B.n716 10.6151
R3466 B.n717 B.n304 10.6151
R3467 B.n727 B.n304 10.6151
R3468 B.n728 B.n727 10.6151
R3469 B.n729 B.n728 10.6151
R3470 B.n729 B.n296 10.6151
R3471 B.n739 B.n296 10.6151
R3472 B.n740 B.n739 10.6151
R3473 B.n741 B.n740 10.6151
R3474 B.n741 B.n287 10.6151
R3475 B.n751 B.n287 10.6151
R3476 B.n752 B.n751 10.6151
R3477 B.n753 B.n752 10.6151
R3478 B.n753 B.n280 10.6151
R3479 B.n763 B.n280 10.6151
R3480 B.n764 B.n763 10.6151
R3481 B.n765 B.n764 10.6151
R3482 B.n765 B.n272 10.6151
R3483 B.n775 B.n272 10.6151
R3484 B.n776 B.n775 10.6151
R3485 B.n777 B.n776 10.6151
R3486 B.n777 B.n263 10.6151
R3487 B.n787 B.n263 10.6151
R3488 B.n788 B.n787 10.6151
R3489 B.n789 B.n788 10.6151
R3490 B.n789 B.n256 10.6151
R3491 B.n799 B.n256 10.6151
R3492 B.n800 B.n799 10.6151
R3493 B.n801 B.n800 10.6151
R3494 B.n801 B.n248 10.6151
R3495 B.n811 B.n248 10.6151
R3496 B.n812 B.n811 10.6151
R3497 B.n813 B.n812 10.6151
R3498 B.n813 B.n240 10.6151
R3499 B.n823 B.n240 10.6151
R3500 B.n824 B.n823 10.6151
R3501 B.n825 B.n824 10.6151
R3502 B.n825 B.n232 10.6151
R3503 B.n835 B.n232 10.6151
R3504 B.n836 B.n835 10.6151
R3505 B.n837 B.n836 10.6151
R3506 B.n837 B.n224 10.6151
R3507 B.n847 B.n224 10.6151
R3508 B.n848 B.n847 10.6151
R3509 B.n849 B.n848 10.6151
R3510 B.n849 B.n216 10.6151
R3511 B.n859 B.n216 10.6151
R3512 B.n860 B.n859 10.6151
R3513 B.n861 B.n860 10.6151
R3514 B.n861 B.n208 10.6151
R3515 B.n871 B.n208 10.6151
R3516 B.n872 B.n871 10.6151
R3517 B.n874 B.n872 10.6151
R3518 B.n874 B.n873 10.6151
R3519 B.n873 B.n200 10.6151
R3520 B.n885 B.n200 10.6151
R3521 B.n886 B.n885 10.6151
R3522 B.n887 B.n886 10.6151
R3523 B.n888 B.n887 10.6151
R3524 B.n889 B.n888 10.6151
R3525 B.n892 B.n889 10.6151
R3526 B.n893 B.n892 10.6151
R3527 B.n894 B.n893 10.6151
R3528 B.n895 B.n894 10.6151
R3529 B.n897 B.n895 10.6151
R3530 B.n898 B.n897 10.6151
R3531 B.n899 B.n898 10.6151
R3532 B.n900 B.n899 10.6151
R3533 B.n902 B.n900 10.6151
R3534 B.n903 B.n902 10.6151
R3535 B.n904 B.n903 10.6151
R3536 B.n905 B.n904 10.6151
R3537 B.n907 B.n905 10.6151
R3538 B.n908 B.n907 10.6151
R3539 B.n909 B.n908 10.6151
R3540 B.n910 B.n909 10.6151
R3541 B.n912 B.n910 10.6151
R3542 B.n913 B.n912 10.6151
R3543 B.n914 B.n913 10.6151
R3544 B.n915 B.n914 10.6151
R3545 B.n917 B.n915 10.6151
R3546 B.n918 B.n917 10.6151
R3547 B.n919 B.n918 10.6151
R3548 B.n920 B.n919 10.6151
R3549 B.n922 B.n920 10.6151
R3550 B.n923 B.n922 10.6151
R3551 B.n924 B.n923 10.6151
R3552 B.n925 B.n924 10.6151
R3553 B.n927 B.n925 10.6151
R3554 B.n928 B.n927 10.6151
R3555 B.n929 B.n928 10.6151
R3556 B.n930 B.n929 10.6151
R3557 B.n932 B.n930 10.6151
R3558 B.n933 B.n932 10.6151
R3559 B.n934 B.n933 10.6151
R3560 B.n935 B.n934 10.6151
R3561 B.n937 B.n935 10.6151
R3562 B.n938 B.n937 10.6151
R3563 B.n939 B.n938 10.6151
R3564 B.n940 B.n939 10.6151
R3565 B.n942 B.n940 10.6151
R3566 B.n943 B.n942 10.6151
R3567 B.n944 B.n943 10.6151
R3568 B.n945 B.n944 10.6151
R3569 B.n947 B.n945 10.6151
R3570 B.n948 B.n947 10.6151
R3571 B.n949 B.n948 10.6151
R3572 B.n950 B.n949 10.6151
R3573 B.n952 B.n950 10.6151
R3574 B.n953 B.n952 10.6151
R3575 B.n954 B.n953 10.6151
R3576 B.n955 B.n954 10.6151
R3577 B.n957 B.n955 10.6151
R3578 B.n958 B.n957 10.6151
R3579 B.n959 B.n958 10.6151
R3580 B.n960 B.n959 10.6151
R3581 B.n962 B.n960 10.6151
R3582 B.n963 B.n962 10.6151
R3583 B.n964 B.n963 10.6151
R3584 B.n965 B.n964 10.6151
R3585 B.n967 B.n965 10.6151
R3586 B.n968 B.n967 10.6151
R3587 B.n969 B.n968 10.6151
R3588 B.n970 B.n969 10.6151
R3589 B.n972 B.n970 10.6151
R3590 B.n973 B.n972 10.6151
R3591 B.n974 B.n973 10.6151
R3592 B.n975 B.n974 10.6151
R3593 B.n1379 B.n1 10.6151
R3594 B.n1379 B.n1378 10.6151
R3595 B.n1378 B.n1377 10.6151
R3596 B.n1377 B.n10 10.6151
R3597 B.n1371 B.n10 10.6151
R3598 B.n1371 B.n1370 10.6151
R3599 B.n1370 B.n1369 10.6151
R3600 B.n1369 B.n18 10.6151
R3601 B.n1363 B.n18 10.6151
R3602 B.n1363 B.n1362 10.6151
R3603 B.n1362 B.n1361 10.6151
R3604 B.n1361 B.n25 10.6151
R3605 B.n1355 B.n25 10.6151
R3606 B.n1355 B.n1354 10.6151
R3607 B.n1354 B.n1353 10.6151
R3608 B.n1353 B.n32 10.6151
R3609 B.n1347 B.n32 10.6151
R3610 B.n1347 B.n1346 10.6151
R3611 B.n1346 B.n1345 10.6151
R3612 B.n1345 B.n39 10.6151
R3613 B.n1339 B.n39 10.6151
R3614 B.n1339 B.n1338 10.6151
R3615 B.n1338 B.n1337 10.6151
R3616 B.n1337 B.n46 10.6151
R3617 B.n1331 B.n46 10.6151
R3618 B.n1331 B.n1330 10.6151
R3619 B.n1330 B.n1329 10.6151
R3620 B.n1329 B.n53 10.6151
R3621 B.n1323 B.n53 10.6151
R3622 B.n1323 B.n1322 10.6151
R3623 B.n1322 B.n1321 10.6151
R3624 B.n1321 B.n60 10.6151
R3625 B.n1315 B.n60 10.6151
R3626 B.n1315 B.n1314 10.6151
R3627 B.n1314 B.n1313 10.6151
R3628 B.n1313 B.n67 10.6151
R3629 B.n1307 B.n67 10.6151
R3630 B.n1307 B.n1306 10.6151
R3631 B.n1306 B.n1305 10.6151
R3632 B.n1305 B.n74 10.6151
R3633 B.n1299 B.n74 10.6151
R3634 B.n1299 B.n1298 10.6151
R3635 B.n1298 B.n1297 10.6151
R3636 B.n1297 B.n81 10.6151
R3637 B.n1291 B.n81 10.6151
R3638 B.n1291 B.n1290 10.6151
R3639 B.n1290 B.n1289 10.6151
R3640 B.n1289 B.n88 10.6151
R3641 B.n1283 B.n88 10.6151
R3642 B.n1283 B.n1282 10.6151
R3643 B.n1282 B.n1281 10.6151
R3644 B.n1281 B.n95 10.6151
R3645 B.n1275 B.n95 10.6151
R3646 B.n1275 B.n1274 10.6151
R3647 B.n1274 B.n1273 10.6151
R3648 B.n1273 B.n102 10.6151
R3649 B.n1267 B.n102 10.6151
R3650 B.n1267 B.n1266 10.6151
R3651 B.n1266 B.n1265 10.6151
R3652 B.n1265 B.n109 10.6151
R3653 B.n1259 B.n109 10.6151
R3654 B.n1259 B.n1258 10.6151
R3655 B.n1258 B.n1257 10.6151
R3656 B.n1257 B.n116 10.6151
R3657 B.n1251 B.n116 10.6151
R3658 B.n1251 B.n1250 10.6151
R3659 B.n1250 B.n1249 10.6151
R3660 B.n1249 B.n123 10.6151
R3661 B.n1243 B.n123 10.6151
R3662 B.n1242 B.n1241 10.6151
R3663 B.n1241 B.n130 10.6151
R3664 B.n1235 B.n130 10.6151
R3665 B.n1235 B.n1234 10.6151
R3666 B.n1234 B.n1233 10.6151
R3667 B.n1233 B.n132 10.6151
R3668 B.n1227 B.n132 10.6151
R3669 B.n1227 B.n1226 10.6151
R3670 B.n1226 B.n1225 10.6151
R3671 B.n1225 B.n134 10.6151
R3672 B.n1219 B.n134 10.6151
R3673 B.n1219 B.n1218 10.6151
R3674 B.n1218 B.n1217 10.6151
R3675 B.n1217 B.n136 10.6151
R3676 B.n1211 B.n136 10.6151
R3677 B.n1211 B.n1210 10.6151
R3678 B.n1210 B.n1209 10.6151
R3679 B.n1209 B.n138 10.6151
R3680 B.n1203 B.n138 10.6151
R3681 B.n1203 B.n1202 10.6151
R3682 B.n1202 B.n1201 10.6151
R3683 B.n1201 B.n140 10.6151
R3684 B.n1195 B.n140 10.6151
R3685 B.n1195 B.n1194 10.6151
R3686 B.n1194 B.n1193 10.6151
R3687 B.n1193 B.n142 10.6151
R3688 B.n1187 B.n142 10.6151
R3689 B.n1187 B.n1186 10.6151
R3690 B.n1186 B.n1185 10.6151
R3691 B.n1185 B.n144 10.6151
R3692 B.n1179 B.n144 10.6151
R3693 B.n1179 B.n1178 10.6151
R3694 B.n1178 B.n1177 10.6151
R3695 B.n1177 B.n146 10.6151
R3696 B.n1171 B.n146 10.6151
R3697 B.n1171 B.n1170 10.6151
R3698 B.n1170 B.n1169 10.6151
R3699 B.n1169 B.n148 10.6151
R3700 B.n1163 B.n148 10.6151
R3701 B.n1163 B.n1162 10.6151
R3702 B.n1162 B.n1161 10.6151
R3703 B.n1161 B.n150 10.6151
R3704 B.n1155 B.n150 10.6151
R3705 B.n1155 B.n1154 10.6151
R3706 B.n1154 B.n1153 10.6151
R3707 B.n1153 B.n152 10.6151
R3708 B.n1147 B.n152 10.6151
R3709 B.n1147 B.n1146 10.6151
R3710 B.n1146 B.n1145 10.6151
R3711 B.n1145 B.n154 10.6151
R3712 B.n1139 B.n154 10.6151
R3713 B.n1139 B.n1138 10.6151
R3714 B.n1138 B.n1137 10.6151
R3715 B.n1137 B.n156 10.6151
R3716 B.n1131 B.n156 10.6151
R3717 B.n1131 B.n1130 10.6151
R3718 B.n1130 B.n1129 10.6151
R3719 B.n1129 B.n158 10.6151
R3720 B.n1123 B.n158 10.6151
R3721 B.n1123 B.n1122 10.6151
R3722 B.n1122 B.n1121 10.6151
R3723 B.n1117 B.n1116 10.6151
R3724 B.n1116 B.n164 10.6151
R3725 B.n1111 B.n164 10.6151
R3726 B.n1111 B.n1110 10.6151
R3727 B.n1110 B.n1109 10.6151
R3728 B.n1109 B.n166 10.6151
R3729 B.n1103 B.n166 10.6151
R3730 B.n1103 B.n1102 10.6151
R3731 B.n1100 B.n170 10.6151
R3732 B.n1094 B.n170 10.6151
R3733 B.n1094 B.n1093 10.6151
R3734 B.n1093 B.n1092 10.6151
R3735 B.n1092 B.n172 10.6151
R3736 B.n1086 B.n172 10.6151
R3737 B.n1086 B.n1085 10.6151
R3738 B.n1085 B.n1084 10.6151
R3739 B.n1084 B.n174 10.6151
R3740 B.n1078 B.n174 10.6151
R3741 B.n1078 B.n1077 10.6151
R3742 B.n1077 B.n1076 10.6151
R3743 B.n1076 B.n176 10.6151
R3744 B.n1070 B.n176 10.6151
R3745 B.n1070 B.n1069 10.6151
R3746 B.n1069 B.n1068 10.6151
R3747 B.n1068 B.n178 10.6151
R3748 B.n1062 B.n178 10.6151
R3749 B.n1062 B.n1061 10.6151
R3750 B.n1061 B.n1060 10.6151
R3751 B.n1060 B.n180 10.6151
R3752 B.n1054 B.n180 10.6151
R3753 B.n1054 B.n1053 10.6151
R3754 B.n1053 B.n1052 10.6151
R3755 B.n1052 B.n182 10.6151
R3756 B.n1046 B.n182 10.6151
R3757 B.n1046 B.n1045 10.6151
R3758 B.n1045 B.n1044 10.6151
R3759 B.n1044 B.n184 10.6151
R3760 B.n1038 B.n184 10.6151
R3761 B.n1038 B.n1037 10.6151
R3762 B.n1037 B.n1036 10.6151
R3763 B.n1036 B.n186 10.6151
R3764 B.n1030 B.n186 10.6151
R3765 B.n1030 B.n1029 10.6151
R3766 B.n1029 B.n1028 10.6151
R3767 B.n1028 B.n188 10.6151
R3768 B.n1022 B.n188 10.6151
R3769 B.n1022 B.n1021 10.6151
R3770 B.n1021 B.n1020 10.6151
R3771 B.n1020 B.n190 10.6151
R3772 B.n1014 B.n190 10.6151
R3773 B.n1014 B.n1013 10.6151
R3774 B.n1013 B.n1012 10.6151
R3775 B.n1012 B.n192 10.6151
R3776 B.n1006 B.n192 10.6151
R3777 B.n1006 B.n1005 10.6151
R3778 B.n1005 B.n1004 10.6151
R3779 B.n1004 B.n194 10.6151
R3780 B.n998 B.n194 10.6151
R3781 B.n998 B.n997 10.6151
R3782 B.n997 B.n996 10.6151
R3783 B.n996 B.n196 10.6151
R3784 B.n990 B.n196 10.6151
R3785 B.n990 B.n989 10.6151
R3786 B.n989 B.n988 10.6151
R3787 B.n988 B.n198 10.6151
R3788 B.n982 B.n198 10.6151
R3789 B.n982 B.n981 10.6151
R3790 B.n981 B.n980 10.6151
R3791 B.n980 B.n976 10.6151
R3792 B.t5 B.n210 10.4745
R3793 B.t7 B.n16 10.4745
R3794 B.n791 B.t2 8.65295
R3795 B.n1319 B.t0 8.65295
R3796 B.n1387 B.n0 8.11757
R3797 B.n1387 B.n1 8.11757
R3798 B.n290 B.t4 7.74217
R3799 B.t3 B.n1294 7.74217
R3800 B.n550 B.n374 6.5566
R3801 B.n534 B.n533 6.5566
R3802 B.n1117 B.n162 6.5566
R3803 B.n1102 B.n1101 6.5566
R3804 B.n827 B.t6 5.9206
R3805 B.n1343 B.t1 5.9206
R3806 B.n374 B.n370 4.05904
R3807 B.n533 B.n532 4.05904
R3808 B.n1121 B.n162 4.05904
R3809 B.n1101 B.n1100 4.05904
R3810 VP.n24 VP.n21 161.3
R3811 VP.n26 VP.n25 161.3
R3812 VP.n27 VP.n20 161.3
R3813 VP.n29 VP.n28 161.3
R3814 VP.n30 VP.n19 161.3
R3815 VP.n32 VP.n31 161.3
R3816 VP.n33 VP.n18 161.3
R3817 VP.n35 VP.n34 161.3
R3818 VP.n36 VP.n17 161.3
R3819 VP.n39 VP.n38 161.3
R3820 VP.n40 VP.n16 161.3
R3821 VP.n42 VP.n41 161.3
R3822 VP.n43 VP.n15 161.3
R3823 VP.n45 VP.n44 161.3
R3824 VP.n46 VP.n14 161.3
R3825 VP.n48 VP.n47 161.3
R3826 VP.n49 VP.n13 161.3
R3827 VP.n92 VP.n0 161.3
R3828 VP.n91 VP.n90 161.3
R3829 VP.n89 VP.n1 161.3
R3830 VP.n88 VP.n87 161.3
R3831 VP.n86 VP.n2 161.3
R3832 VP.n85 VP.n84 161.3
R3833 VP.n83 VP.n3 161.3
R3834 VP.n82 VP.n81 161.3
R3835 VP.n79 VP.n4 161.3
R3836 VP.n78 VP.n77 161.3
R3837 VP.n76 VP.n5 161.3
R3838 VP.n75 VP.n74 161.3
R3839 VP.n73 VP.n6 161.3
R3840 VP.n72 VP.n71 161.3
R3841 VP.n70 VP.n7 161.3
R3842 VP.n69 VP.n68 161.3
R3843 VP.n67 VP.n8 161.3
R3844 VP.n65 VP.n64 161.3
R3845 VP.n63 VP.n9 161.3
R3846 VP.n62 VP.n61 161.3
R3847 VP.n60 VP.n10 161.3
R3848 VP.n59 VP.n58 161.3
R3849 VP.n57 VP.n11 161.3
R3850 VP.n56 VP.n55 161.3
R3851 VP.n54 VP.n12 161.3
R3852 VP.n22 VP.t7 148.778
R3853 VP.n53 VP.t0 116.371
R3854 VP.n66 VP.t2 116.371
R3855 VP.n80 VP.t1 116.371
R3856 VP.n93 VP.t5 116.371
R3857 VP.n50 VP.t3 116.371
R3858 VP.n37 VP.t6 116.371
R3859 VP.n23 VP.t4 116.371
R3860 VP.n23 VP.n22 69.3059
R3861 VP.n53 VP.n52 64.6738
R3862 VP.n94 VP.n93 64.6738
R3863 VP.n51 VP.n50 64.6738
R3864 VP.n52 VP.n51 62.4211
R3865 VP.n87 VP.n86 56.5617
R3866 VP.n60 VP.n59 56.5617
R3867 VP.n44 VP.n43 56.5617
R3868 VP.n73 VP.n72 40.577
R3869 VP.n74 VP.n73 40.577
R3870 VP.n31 VP.n30 40.577
R3871 VP.n30 VP.n29 40.577
R3872 VP.n55 VP.n54 24.5923
R3873 VP.n55 VP.n11 24.5923
R3874 VP.n59 VP.n11 24.5923
R3875 VP.n61 VP.n60 24.5923
R3876 VP.n61 VP.n9 24.5923
R3877 VP.n65 VP.n9 24.5923
R3878 VP.n68 VP.n67 24.5923
R3879 VP.n68 VP.n7 24.5923
R3880 VP.n72 VP.n7 24.5923
R3881 VP.n74 VP.n5 24.5923
R3882 VP.n78 VP.n5 24.5923
R3883 VP.n79 VP.n78 24.5923
R3884 VP.n81 VP.n3 24.5923
R3885 VP.n85 VP.n3 24.5923
R3886 VP.n86 VP.n85 24.5923
R3887 VP.n87 VP.n1 24.5923
R3888 VP.n91 VP.n1 24.5923
R3889 VP.n92 VP.n91 24.5923
R3890 VP.n44 VP.n14 24.5923
R3891 VP.n48 VP.n14 24.5923
R3892 VP.n49 VP.n48 24.5923
R3893 VP.n31 VP.n18 24.5923
R3894 VP.n35 VP.n18 24.5923
R3895 VP.n36 VP.n35 24.5923
R3896 VP.n38 VP.n16 24.5923
R3897 VP.n42 VP.n16 24.5923
R3898 VP.n43 VP.n42 24.5923
R3899 VP.n25 VP.n24 24.5923
R3900 VP.n25 VP.n20 24.5923
R3901 VP.n29 VP.n20 24.5923
R3902 VP.n66 VP.n65 18.6903
R3903 VP.n81 VP.n80 18.6903
R3904 VP.n38 VP.n37 18.6903
R3905 VP.n54 VP.n53 17.7066
R3906 VP.n93 VP.n92 17.7066
R3907 VP.n50 VP.n49 17.7066
R3908 VP.n67 VP.n66 5.90254
R3909 VP.n80 VP.n79 5.90254
R3910 VP.n37 VP.n36 5.90254
R3911 VP.n24 VP.n23 5.90254
R3912 VP.n22 VP.n21 2.76473
R3913 VP.n51 VP.n13 0.417304
R3914 VP.n52 VP.n12 0.417304
R3915 VP.n94 VP.n0 0.417304
R3916 VP VP.n94 0.394524
R3917 VP.n26 VP.n21 0.189894
R3918 VP.n27 VP.n26 0.189894
R3919 VP.n28 VP.n27 0.189894
R3920 VP.n28 VP.n19 0.189894
R3921 VP.n32 VP.n19 0.189894
R3922 VP.n33 VP.n32 0.189894
R3923 VP.n34 VP.n33 0.189894
R3924 VP.n34 VP.n17 0.189894
R3925 VP.n39 VP.n17 0.189894
R3926 VP.n40 VP.n39 0.189894
R3927 VP.n41 VP.n40 0.189894
R3928 VP.n41 VP.n15 0.189894
R3929 VP.n45 VP.n15 0.189894
R3930 VP.n46 VP.n45 0.189894
R3931 VP.n47 VP.n46 0.189894
R3932 VP.n47 VP.n13 0.189894
R3933 VP.n56 VP.n12 0.189894
R3934 VP.n57 VP.n56 0.189894
R3935 VP.n58 VP.n57 0.189894
R3936 VP.n58 VP.n10 0.189894
R3937 VP.n62 VP.n10 0.189894
R3938 VP.n63 VP.n62 0.189894
R3939 VP.n64 VP.n63 0.189894
R3940 VP.n64 VP.n8 0.189894
R3941 VP.n69 VP.n8 0.189894
R3942 VP.n70 VP.n69 0.189894
R3943 VP.n71 VP.n70 0.189894
R3944 VP.n71 VP.n6 0.189894
R3945 VP.n75 VP.n6 0.189894
R3946 VP.n76 VP.n75 0.189894
R3947 VP.n77 VP.n76 0.189894
R3948 VP.n77 VP.n4 0.189894
R3949 VP.n82 VP.n4 0.189894
R3950 VP.n83 VP.n82 0.189894
R3951 VP.n84 VP.n83 0.189894
R3952 VP.n84 VP.n2 0.189894
R3953 VP.n88 VP.n2 0.189894
R3954 VP.n89 VP.n88 0.189894
R3955 VP.n90 VP.n89 0.189894
R3956 VP.n90 VP.n0 0.189894
R3957 VDD1 VDD1.n0 60.9562
R3958 VDD1.n3 VDD1.n2 60.8427
R3959 VDD1.n3 VDD1.n1 60.8427
R3960 VDD1.n5 VDD1.n4 59.0703
R3961 VDD1.n5 VDD1.n3 57.0224
R3962 VDD1 VDD1.n5 1.7699
R3963 VDD1.n4 VDD1.t1 1.04923
R3964 VDD1.n4 VDD1.t4 1.04923
R3965 VDD1.n0 VDD1.t0 1.04923
R3966 VDD1.n0 VDD1.t3 1.04923
R3967 VDD1.n2 VDD1.t6 1.04923
R3968 VDD1.n2 VDD1.t2 1.04923
R3969 VDD1.n1 VDD1.t7 1.04923
R3970 VDD1.n1 VDD1.t5 1.04923
C0 VTAIL VDD2 10.619201f
C1 VDD1 VDD2 2.45874f
C2 VTAIL VDD1 10.556f
C3 VDD2 VP 0.659553f
C4 VTAIL VP 14.872299f
C5 VDD2 VN 14.345401f
C6 VTAIL VN 14.8581f
C7 VDD1 VP 14.8483f
C8 VDD1 VN 0.154581f
C9 VP VN 10.5368f
C10 VDD2 B 7.224166f
C11 VDD1 B 7.80208f
C12 VTAIL B 15.532107f
C13 VN B 21.105122f
C14 VP B 19.712936f
C15 VDD1.t0 B 0.398984f
C16 VDD1.t3 B 0.398984f
C17 VDD1.n0 B 3.6608f
C18 VDD1.t7 B 0.398984f
C19 VDD1.t5 B 0.398984f
C20 VDD1.n1 B 3.65924f
C21 VDD1.t6 B 0.398984f
C22 VDD1.t2 B 0.398984f
C23 VDD1.n2 B 3.65924f
C24 VDD1.n3 B 4.84938f
C25 VDD1.t1 B 0.398984f
C26 VDD1.t4 B 0.398984f
C27 VDD1.n4 B 3.63871f
C28 VDD1.n5 B 4.23393f
C29 VP.n0 B 0.030143f
C30 VP.t5 B 3.25767f
C31 VP.n1 B 0.029725f
C32 VP.n2 B 0.01603f
C33 VP.n3 B 0.029725f
C34 VP.n4 B 0.01603f
C35 VP.t1 B 3.25767f
C36 VP.n5 B 0.029725f
C37 VP.n6 B 0.01603f
C38 VP.n7 B 0.029725f
C39 VP.n8 B 0.01603f
C40 VP.t2 B 3.25767f
C41 VP.n9 B 0.029725f
C42 VP.n10 B 0.01603f
C43 VP.n11 B 0.029725f
C44 VP.n12 B 0.030143f
C45 VP.t0 B 3.25767f
C46 VP.n13 B 0.030143f
C47 VP.t3 B 3.25767f
C48 VP.n14 B 0.029725f
C49 VP.n15 B 0.01603f
C50 VP.n16 B 0.029725f
C51 VP.n17 B 0.01603f
C52 VP.t6 B 3.25767f
C53 VP.n18 B 0.029725f
C54 VP.n19 B 0.01603f
C55 VP.n20 B 0.029725f
C56 VP.n21 B 0.213872f
C57 VP.t4 B 3.25767f
C58 VP.t7 B 3.52842f
C59 VP.n22 B 1.12059f
C60 VP.n23 B 1.17409f
C61 VP.n24 B 0.018573f
C62 VP.n25 B 0.029725f
C63 VP.n26 B 0.01603f
C64 VP.n27 B 0.01603f
C65 VP.n28 B 0.01603f
C66 VP.n29 B 0.031691f
C67 VP.n30 B 0.012947f
C68 VP.n31 B 0.031691f
C69 VP.n32 B 0.01603f
C70 VP.n33 B 0.01603f
C71 VP.n34 B 0.01603f
C72 VP.n35 B 0.029725f
C73 VP.n36 B 0.018573f
C74 VP.n37 B 1.12008f
C75 VP.n38 B 0.026204f
C76 VP.n39 B 0.01603f
C77 VP.n40 B 0.01603f
C78 VP.n41 B 0.01603f
C79 VP.n42 B 0.029725f
C80 VP.n43 B 0.022858f
C81 VP.n44 B 0.023745f
C82 VP.n45 B 0.01603f
C83 VP.n46 B 0.01603f
C84 VP.n47 B 0.01603f
C85 VP.n48 B 0.029725f
C86 VP.n49 B 0.025617f
C87 VP.n50 B 1.18629f
C88 VP.n51 B 1.25872f
C89 VP.n52 B 1.26798f
C90 VP.n53 B 1.18629f
C91 VP.n54 B 0.025617f
C92 VP.n55 B 0.029725f
C93 VP.n56 B 0.01603f
C94 VP.n57 B 0.01603f
C95 VP.n58 B 0.01603f
C96 VP.n59 B 0.023745f
C97 VP.n60 B 0.022858f
C98 VP.n61 B 0.029725f
C99 VP.n62 B 0.01603f
C100 VP.n63 B 0.01603f
C101 VP.n64 B 0.01603f
C102 VP.n65 B 0.026204f
C103 VP.n66 B 1.12008f
C104 VP.n67 B 0.018573f
C105 VP.n68 B 0.029725f
C106 VP.n69 B 0.01603f
C107 VP.n70 B 0.01603f
C108 VP.n71 B 0.01603f
C109 VP.n72 B 0.031691f
C110 VP.n73 B 0.012947f
C111 VP.n74 B 0.031691f
C112 VP.n75 B 0.01603f
C113 VP.n76 B 0.01603f
C114 VP.n77 B 0.01603f
C115 VP.n78 B 0.029725f
C116 VP.n79 B 0.018573f
C117 VP.n80 B 1.12008f
C118 VP.n81 B 0.026204f
C119 VP.n82 B 0.01603f
C120 VP.n83 B 0.01603f
C121 VP.n84 B 0.01603f
C122 VP.n85 B 0.029725f
C123 VP.n86 B 0.022858f
C124 VP.n87 B 0.023745f
C125 VP.n88 B 0.01603f
C126 VP.n89 B 0.01603f
C127 VP.n90 B 0.01603f
C128 VP.n91 B 0.029725f
C129 VP.n92 B 0.025617f
C130 VP.n93 B 1.18629f
C131 VP.n94 B 0.0527f
C132 VTAIL.t3 B 0.285155f
C133 VTAIL.t10 B 0.285155f
C134 VTAIL.n0 B 2.53856f
C135 VTAIL.n1 B 0.426082f
C136 VTAIL.n2 B 0.026349f
C137 VTAIL.n3 B 0.019113f
C138 VTAIL.n4 B 0.01027f
C139 VTAIL.n5 B 0.024275f
C140 VTAIL.n6 B 0.010875f
C141 VTAIL.n7 B 0.019113f
C142 VTAIL.n8 B 0.01027f
C143 VTAIL.n9 B 0.024275f
C144 VTAIL.n10 B 0.010875f
C145 VTAIL.n11 B 0.019113f
C146 VTAIL.n12 B 0.01027f
C147 VTAIL.n13 B 0.024275f
C148 VTAIL.n14 B 0.010875f
C149 VTAIL.n15 B 0.019113f
C150 VTAIL.n16 B 0.01027f
C151 VTAIL.n17 B 0.024275f
C152 VTAIL.n18 B 0.010875f
C153 VTAIL.n19 B 0.019113f
C154 VTAIL.n20 B 0.01027f
C155 VTAIL.n21 B 0.024275f
C156 VTAIL.n22 B 0.010875f
C157 VTAIL.n23 B 0.019113f
C158 VTAIL.n24 B 0.01027f
C159 VTAIL.n25 B 0.024275f
C160 VTAIL.n26 B 0.010875f
C161 VTAIL.n27 B 0.019113f
C162 VTAIL.n28 B 0.01027f
C163 VTAIL.n29 B 0.024275f
C164 VTAIL.n30 B 0.010875f
C165 VTAIL.n31 B 0.019113f
C166 VTAIL.n32 B 0.01027f
C167 VTAIL.n33 B 0.024275f
C168 VTAIL.n34 B 0.010875f
C169 VTAIL.n35 B 0.143251f
C170 VTAIL.t9 B 0.040282f
C171 VTAIL.n36 B 0.018207f
C172 VTAIL.n37 B 0.01434f
C173 VTAIL.n38 B 0.01027f
C174 VTAIL.n39 B 1.58338f
C175 VTAIL.n40 B 0.019113f
C176 VTAIL.n41 B 0.01027f
C177 VTAIL.n42 B 0.010875f
C178 VTAIL.n43 B 0.024275f
C179 VTAIL.n44 B 0.024275f
C180 VTAIL.n45 B 0.010875f
C181 VTAIL.n46 B 0.01027f
C182 VTAIL.n47 B 0.019113f
C183 VTAIL.n48 B 0.019113f
C184 VTAIL.n49 B 0.01027f
C185 VTAIL.n50 B 0.010875f
C186 VTAIL.n51 B 0.024275f
C187 VTAIL.n52 B 0.024275f
C188 VTAIL.n53 B 0.010875f
C189 VTAIL.n54 B 0.01027f
C190 VTAIL.n55 B 0.019113f
C191 VTAIL.n56 B 0.019113f
C192 VTAIL.n57 B 0.01027f
C193 VTAIL.n58 B 0.010875f
C194 VTAIL.n59 B 0.024275f
C195 VTAIL.n60 B 0.024275f
C196 VTAIL.n61 B 0.010875f
C197 VTAIL.n62 B 0.01027f
C198 VTAIL.n63 B 0.019113f
C199 VTAIL.n64 B 0.019113f
C200 VTAIL.n65 B 0.01027f
C201 VTAIL.n66 B 0.010875f
C202 VTAIL.n67 B 0.024275f
C203 VTAIL.n68 B 0.024275f
C204 VTAIL.n69 B 0.010875f
C205 VTAIL.n70 B 0.01027f
C206 VTAIL.n71 B 0.019113f
C207 VTAIL.n72 B 0.019113f
C208 VTAIL.n73 B 0.01027f
C209 VTAIL.n74 B 0.010875f
C210 VTAIL.n75 B 0.024275f
C211 VTAIL.n76 B 0.024275f
C212 VTAIL.n77 B 0.024275f
C213 VTAIL.n78 B 0.010875f
C214 VTAIL.n79 B 0.01027f
C215 VTAIL.n80 B 0.019113f
C216 VTAIL.n81 B 0.019113f
C217 VTAIL.n82 B 0.01027f
C218 VTAIL.n83 B 0.010573f
C219 VTAIL.n84 B 0.010573f
C220 VTAIL.n85 B 0.024275f
C221 VTAIL.n86 B 0.024275f
C222 VTAIL.n87 B 0.010875f
C223 VTAIL.n88 B 0.01027f
C224 VTAIL.n89 B 0.019113f
C225 VTAIL.n90 B 0.019113f
C226 VTAIL.n91 B 0.01027f
C227 VTAIL.n92 B 0.010875f
C228 VTAIL.n93 B 0.024275f
C229 VTAIL.n94 B 0.024275f
C230 VTAIL.n95 B 0.010875f
C231 VTAIL.n96 B 0.01027f
C232 VTAIL.n97 B 0.019113f
C233 VTAIL.n98 B 0.019113f
C234 VTAIL.n99 B 0.01027f
C235 VTAIL.n100 B 0.010875f
C236 VTAIL.n101 B 0.024275f
C237 VTAIL.n102 B 0.05164f
C238 VTAIL.n103 B 0.010875f
C239 VTAIL.n104 B 0.01027f
C240 VTAIL.n105 B 0.04209f
C241 VTAIL.n106 B 0.028735f
C242 VTAIL.n107 B 0.269188f
C243 VTAIL.n108 B 0.026349f
C244 VTAIL.n109 B 0.019113f
C245 VTAIL.n110 B 0.01027f
C246 VTAIL.n111 B 0.024275f
C247 VTAIL.n112 B 0.010875f
C248 VTAIL.n113 B 0.019113f
C249 VTAIL.n114 B 0.01027f
C250 VTAIL.n115 B 0.024275f
C251 VTAIL.n116 B 0.010875f
C252 VTAIL.n117 B 0.019113f
C253 VTAIL.n118 B 0.01027f
C254 VTAIL.n119 B 0.024275f
C255 VTAIL.n120 B 0.010875f
C256 VTAIL.n121 B 0.019113f
C257 VTAIL.n122 B 0.01027f
C258 VTAIL.n123 B 0.024275f
C259 VTAIL.n124 B 0.010875f
C260 VTAIL.n125 B 0.019113f
C261 VTAIL.n126 B 0.01027f
C262 VTAIL.n127 B 0.024275f
C263 VTAIL.n128 B 0.010875f
C264 VTAIL.n129 B 0.019113f
C265 VTAIL.n130 B 0.01027f
C266 VTAIL.n131 B 0.024275f
C267 VTAIL.n132 B 0.010875f
C268 VTAIL.n133 B 0.019113f
C269 VTAIL.n134 B 0.01027f
C270 VTAIL.n135 B 0.024275f
C271 VTAIL.n136 B 0.010875f
C272 VTAIL.n137 B 0.019113f
C273 VTAIL.n138 B 0.01027f
C274 VTAIL.n139 B 0.024275f
C275 VTAIL.n140 B 0.010875f
C276 VTAIL.n141 B 0.143251f
C277 VTAIL.t11 B 0.040282f
C278 VTAIL.n142 B 0.018207f
C279 VTAIL.n143 B 0.01434f
C280 VTAIL.n144 B 0.01027f
C281 VTAIL.n145 B 1.58338f
C282 VTAIL.n146 B 0.019113f
C283 VTAIL.n147 B 0.01027f
C284 VTAIL.n148 B 0.010875f
C285 VTAIL.n149 B 0.024275f
C286 VTAIL.n150 B 0.024275f
C287 VTAIL.n151 B 0.010875f
C288 VTAIL.n152 B 0.01027f
C289 VTAIL.n153 B 0.019113f
C290 VTAIL.n154 B 0.019113f
C291 VTAIL.n155 B 0.01027f
C292 VTAIL.n156 B 0.010875f
C293 VTAIL.n157 B 0.024275f
C294 VTAIL.n158 B 0.024275f
C295 VTAIL.n159 B 0.010875f
C296 VTAIL.n160 B 0.01027f
C297 VTAIL.n161 B 0.019113f
C298 VTAIL.n162 B 0.019113f
C299 VTAIL.n163 B 0.01027f
C300 VTAIL.n164 B 0.010875f
C301 VTAIL.n165 B 0.024275f
C302 VTAIL.n166 B 0.024275f
C303 VTAIL.n167 B 0.010875f
C304 VTAIL.n168 B 0.01027f
C305 VTAIL.n169 B 0.019113f
C306 VTAIL.n170 B 0.019113f
C307 VTAIL.n171 B 0.01027f
C308 VTAIL.n172 B 0.010875f
C309 VTAIL.n173 B 0.024275f
C310 VTAIL.n174 B 0.024275f
C311 VTAIL.n175 B 0.010875f
C312 VTAIL.n176 B 0.01027f
C313 VTAIL.n177 B 0.019113f
C314 VTAIL.n178 B 0.019113f
C315 VTAIL.n179 B 0.01027f
C316 VTAIL.n180 B 0.010875f
C317 VTAIL.n181 B 0.024275f
C318 VTAIL.n182 B 0.024275f
C319 VTAIL.n183 B 0.024275f
C320 VTAIL.n184 B 0.010875f
C321 VTAIL.n185 B 0.01027f
C322 VTAIL.n186 B 0.019113f
C323 VTAIL.n187 B 0.019113f
C324 VTAIL.n188 B 0.01027f
C325 VTAIL.n189 B 0.010573f
C326 VTAIL.n190 B 0.010573f
C327 VTAIL.n191 B 0.024275f
C328 VTAIL.n192 B 0.024275f
C329 VTAIL.n193 B 0.010875f
C330 VTAIL.n194 B 0.01027f
C331 VTAIL.n195 B 0.019113f
C332 VTAIL.n196 B 0.019113f
C333 VTAIL.n197 B 0.01027f
C334 VTAIL.n198 B 0.010875f
C335 VTAIL.n199 B 0.024275f
C336 VTAIL.n200 B 0.024275f
C337 VTAIL.n201 B 0.010875f
C338 VTAIL.n202 B 0.01027f
C339 VTAIL.n203 B 0.019113f
C340 VTAIL.n204 B 0.019113f
C341 VTAIL.n205 B 0.01027f
C342 VTAIL.n206 B 0.010875f
C343 VTAIL.n207 B 0.024275f
C344 VTAIL.n208 B 0.05164f
C345 VTAIL.n209 B 0.010875f
C346 VTAIL.n210 B 0.01027f
C347 VTAIL.n211 B 0.04209f
C348 VTAIL.n212 B 0.028735f
C349 VTAIL.n213 B 0.269188f
C350 VTAIL.t2 B 0.285155f
C351 VTAIL.t15 B 0.285155f
C352 VTAIL.n214 B 2.53856f
C353 VTAIL.n215 B 0.647605f
C354 VTAIL.n216 B 0.026349f
C355 VTAIL.n217 B 0.019113f
C356 VTAIL.n218 B 0.01027f
C357 VTAIL.n219 B 0.024275f
C358 VTAIL.n220 B 0.010875f
C359 VTAIL.n221 B 0.019113f
C360 VTAIL.n222 B 0.01027f
C361 VTAIL.n223 B 0.024275f
C362 VTAIL.n224 B 0.010875f
C363 VTAIL.n225 B 0.019113f
C364 VTAIL.n226 B 0.01027f
C365 VTAIL.n227 B 0.024275f
C366 VTAIL.n228 B 0.010875f
C367 VTAIL.n229 B 0.019113f
C368 VTAIL.n230 B 0.01027f
C369 VTAIL.n231 B 0.024275f
C370 VTAIL.n232 B 0.010875f
C371 VTAIL.n233 B 0.019113f
C372 VTAIL.n234 B 0.01027f
C373 VTAIL.n235 B 0.024275f
C374 VTAIL.n236 B 0.010875f
C375 VTAIL.n237 B 0.019113f
C376 VTAIL.n238 B 0.01027f
C377 VTAIL.n239 B 0.024275f
C378 VTAIL.n240 B 0.010875f
C379 VTAIL.n241 B 0.019113f
C380 VTAIL.n242 B 0.01027f
C381 VTAIL.n243 B 0.024275f
C382 VTAIL.n244 B 0.010875f
C383 VTAIL.n245 B 0.019113f
C384 VTAIL.n246 B 0.01027f
C385 VTAIL.n247 B 0.024275f
C386 VTAIL.n248 B 0.010875f
C387 VTAIL.n249 B 0.143251f
C388 VTAIL.t13 B 0.040282f
C389 VTAIL.n250 B 0.018207f
C390 VTAIL.n251 B 0.01434f
C391 VTAIL.n252 B 0.01027f
C392 VTAIL.n253 B 1.58338f
C393 VTAIL.n254 B 0.019113f
C394 VTAIL.n255 B 0.01027f
C395 VTAIL.n256 B 0.010875f
C396 VTAIL.n257 B 0.024275f
C397 VTAIL.n258 B 0.024275f
C398 VTAIL.n259 B 0.010875f
C399 VTAIL.n260 B 0.01027f
C400 VTAIL.n261 B 0.019113f
C401 VTAIL.n262 B 0.019113f
C402 VTAIL.n263 B 0.01027f
C403 VTAIL.n264 B 0.010875f
C404 VTAIL.n265 B 0.024275f
C405 VTAIL.n266 B 0.024275f
C406 VTAIL.n267 B 0.010875f
C407 VTAIL.n268 B 0.01027f
C408 VTAIL.n269 B 0.019113f
C409 VTAIL.n270 B 0.019113f
C410 VTAIL.n271 B 0.01027f
C411 VTAIL.n272 B 0.010875f
C412 VTAIL.n273 B 0.024275f
C413 VTAIL.n274 B 0.024275f
C414 VTAIL.n275 B 0.010875f
C415 VTAIL.n276 B 0.01027f
C416 VTAIL.n277 B 0.019113f
C417 VTAIL.n278 B 0.019113f
C418 VTAIL.n279 B 0.01027f
C419 VTAIL.n280 B 0.010875f
C420 VTAIL.n281 B 0.024275f
C421 VTAIL.n282 B 0.024275f
C422 VTAIL.n283 B 0.010875f
C423 VTAIL.n284 B 0.01027f
C424 VTAIL.n285 B 0.019113f
C425 VTAIL.n286 B 0.019113f
C426 VTAIL.n287 B 0.01027f
C427 VTAIL.n288 B 0.010875f
C428 VTAIL.n289 B 0.024275f
C429 VTAIL.n290 B 0.024275f
C430 VTAIL.n291 B 0.024275f
C431 VTAIL.n292 B 0.010875f
C432 VTAIL.n293 B 0.01027f
C433 VTAIL.n294 B 0.019113f
C434 VTAIL.n295 B 0.019113f
C435 VTAIL.n296 B 0.01027f
C436 VTAIL.n297 B 0.010573f
C437 VTAIL.n298 B 0.010573f
C438 VTAIL.n299 B 0.024275f
C439 VTAIL.n300 B 0.024275f
C440 VTAIL.n301 B 0.010875f
C441 VTAIL.n302 B 0.01027f
C442 VTAIL.n303 B 0.019113f
C443 VTAIL.n304 B 0.019113f
C444 VTAIL.n305 B 0.01027f
C445 VTAIL.n306 B 0.010875f
C446 VTAIL.n307 B 0.024275f
C447 VTAIL.n308 B 0.024275f
C448 VTAIL.n309 B 0.010875f
C449 VTAIL.n310 B 0.01027f
C450 VTAIL.n311 B 0.019113f
C451 VTAIL.n312 B 0.019113f
C452 VTAIL.n313 B 0.01027f
C453 VTAIL.n314 B 0.010875f
C454 VTAIL.n315 B 0.024275f
C455 VTAIL.n316 B 0.05164f
C456 VTAIL.n317 B 0.010875f
C457 VTAIL.n318 B 0.01027f
C458 VTAIL.n319 B 0.04209f
C459 VTAIL.n320 B 0.028735f
C460 VTAIL.n321 B 1.72735f
C461 VTAIL.n322 B 0.026349f
C462 VTAIL.n323 B 0.019113f
C463 VTAIL.n324 B 0.01027f
C464 VTAIL.n325 B 0.024275f
C465 VTAIL.n326 B 0.010875f
C466 VTAIL.n327 B 0.019113f
C467 VTAIL.n328 B 0.01027f
C468 VTAIL.n329 B 0.024275f
C469 VTAIL.n330 B 0.010875f
C470 VTAIL.n331 B 0.019113f
C471 VTAIL.n332 B 0.01027f
C472 VTAIL.n333 B 0.024275f
C473 VTAIL.n334 B 0.010875f
C474 VTAIL.n335 B 0.019113f
C475 VTAIL.n336 B 0.01027f
C476 VTAIL.n337 B 0.024275f
C477 VTAIL.n338 B 0.024275f
C478 VTAIL.n339 B 0.010875f
C479 VTAIL.n340 B 0.019113f
C480 VTAIL.n341 B 0.01027f
C481 VTAIL.n342 B 0.024275f
C482 VTAIL.n343 B 0.010875f
C483 VTAIL.n344 B 0.019113f
C484 VTAIL.n345 B 0.01027f
C485 VTAIL.n346 B 0.024275f
C486 VTAIL.n347 B 0.010875f
C487 VTAIL.n348 B 0.019113f
C488 VTAIL.n349 B 0.01027f
C489 VTAIL.n350 B 0.024275f
C490 VTAIL.n351 B 0.010875f
C491 VTAIL.n352 B 0.019113f
C492 VTAIL.n353 B 0.01027f
C493 VTAIL.n354 B 0.024275f
C494 VTAIL.n355 B 0.010875f
C495 VTAIL.n356 B 0.143251f
C496 VTAIL.t6 B 0.040282f
C497 VTAIL.n357 B 0.018207f
C498 VTAIL.n358 B 0.01434f
C499 VTAIL.n359 B 0.01027f
C500 VTAIL.n360 B 1.58338f
C501 VTAIL.n361 B 0.019113f
C502 VTAIL.n362 B 0.01027f
C503 VTAIL.n363 B 0.010875f
C504 VTAIL.n364 B 0.024275f
C505 VTAIL.n365 B 0.024275f
C506 VTAIL.n366 B 0.010875f
C507 VTAIL.n367 B 0.01027f
C508 VTAIL.n368 B 0.019113f
C509 VTAIL.n369 B 0.019113f
C510 VTAIL.n370 B 0.01027f
C511 VTAIL.n371 B 0.010875f
C512 VTAIL.n372 B 0.024275f
C513 VTAIL.n373 B 0.024275f
C514 VTAIL.n374 B 0.010875f
C515 VTAIL.n375 B 0.01027f
C516 VTAIL.n376 B 0.019113f
C517 VTAIL.n377 B 0.019113f
C518 VTAIL.n378 B 0.01027f
C519 VTAIL.n379 B 0.010875f
C520 VTAIL.n380 B 0.024275f
C521 VTAIL.n381 B 0.024275f
C522 VTAIL.n382 B 0.010875f
C523 VTAIL.n383 B 0.01027f
C524 VTAIL.n384 B 0.019113f
C525 VTAIL.n385 B 0.019113f
C526 VTAIL.n386 B 0.01027f
C527 VTAIL.n387 B 0.010875f
C528 VTAIL.n388 B 0.024275f
C529 VTAIL.n389 B 0.024275f
C530 VTAIL.n390 B 0.010875f
C531 VTAIL.n391 B 0.01027f
C532 VTAIL.n392 B 0.019113f
C533 VTAIL.n393 B 0.019113f
C534 VTAIL.n394 B 0.01027f
C535 VTAIL.n395 B 0.010875f
C536 VTAIL.n396 B 0.024275f
C537 VTAIL.n397 B 0.024275f
C538 VTAIL.n398 B 0.010875f
C539 VTAIL.n399 B 0.01027f
C540 VTAIL.n400 B 0.019113f
C541 VTAIL.n401 B 0.019113f
C542 VTAIL.n402 B 0.01027f
C543 VTAIL.n403 B 0.010573f
C544 VTAIL.n404 B 0.010573f
C545 VTAIL.n405 B 0.024275f
C546 VTAIL.n406 B 0.024275f
C547 VTAIL.n407 B 0.010875f
C548 VTAIL.n408 B 0.01027f
C549 VTAIL.n409 B 0.019113f
C550 VTAIL.n410 B 0.019113f
C551 VTAIL.n411 B 0.01027f
C552 VTAIL.n412 B 0.010875f
C553 VTAIL.n413 B 0.024275f
C554 VTAIL.n414 B 0.024275f
C555 VTAIL.n415 B 0.010875f
C556 VTAIL.n416 B 0.01027f
C557 VTAIL.n417 B 0.019113f
C558 VTAIL.n418 B 0.019113f
C559 VTAIL.n419 B 0.01027f
C560 VTAIL.n420 B 0.010875f
C561 VTAIL.n421 B 0.024275f
C562 VTAIL.n422 B 0.05164f
C563 VTAIL.n423 B 0.010875f
C564 VTAIL.n424 B 0.01027f
C565 VTAIL.n425 B 0.04209f
C566 VTAIL.n426 B 0.028735f
C567 VTAIL.n427 B 1.72735f
C568 VTAIL.t4 B 0.285155f
C569 VTAIL.t8 B 0.285155f
C570 VTAIL.n428 B 2.53856f
C571 VTAIL.n429 B 0.647604f
C572 VTAIL.n430 B 0.026349f
C573 VTAIL.n431 B 0.019113f
C574 VTAIL.n432 B 0.01027f
C575 VTAIL.n433 B 0.024275f
C576 VTAIL.n434 B 0.010875f
C577 VTAIL.n435 B 0.019113f
C578 VTAIL.n436 B 0.01027f
C579 VTAIL.n437 B 0.024275f
C580 VTAIL.n438 B 0.010875f
C581 VTAIL.n439 B 0.019113f
C582 VTAIL.n440 B 0.01027f
C583 VTAIL.n441 B 0.024275f
C584 VTAIL.n442 B 0.010875f
C585 VTAIL.n443 B 0.019113f
C586 VTAIL.n444 B 0.01027f
C587 VTAIL.n445 B 0.024275f
C588 VTAIL.n446 B 0.024275f
C589 VTAIL.n447 B 0.010875f
C590 VTAIL.n448 B 0.019113f
C591 VTAIL.n449 B 0.01027f
C592 VTAIL.n450 B 0.024275f
C593 VTAIL.n451 B 0.010875f
C594 VTAIL.n452 B 0.019113f
C595 VTAIL.n453 B 0.01027f
C596 VTAIL.n454 B 0.024275f
C597 VTAIL.n455 B 0.010875f
C598 VTAIL.n456 B 0.019113f
C599 VTAIL.n457 B 0.01027f
C600 VTAIL.n458 B 0.024275f
C601 VTAIL.n459 B 0.010875f
C602 VTAIL.n460 B 0.019113f
C603 VTAIL.n461 B 0.01027f
C604 VTAIL.n462 B 0.024275f
C605 VTAIL.n463 B 0.010875f
C606 VTAIL.n464 B 0.143251f
C607 VTAIL.t7 B 0.040282f
C608 VTAIL.n465 B 0.018207f
C609 VTAIL.n466 B 0.01434f
C610 VTAIL.n467 B 0.01027f
C611 VTAIL.n468 B 1.58338f
C612 VTAIL.n469 B 0.019113f
C613 VTAIL.n470 B 0.01027f
C614 VTAIL.n471 B 0.010875f
C615 VTAIL.n472 B 0.024275f
C616 VTAIL.n473 B 0.024275f
C617 VTAIL.n474 B 0.010875f
C618 VTAIL.n475 B 0.01027f
C619 VTAIL.n476 B 0.019113f
C620 VTAIL.n477 B 0.019113f
C621 VTAIL.n478 B 0.01027f
C622 VTAIL.n479 B 0.010875f
C623 VTAIL.n480 B 0.024275f
C624 VTAIL.n481 B 0.024275f
C625 VTAIL.n482 B 0.010875f
C626 VTAIL.n483 B 0.01027f
C627 VTAIL.n484 B 0.019113f
C628 VTAIL.n485 B 0.019113f
C629 VTAIL.n486 B 0.01027f
C630 VTAIL.n487 B 0.010875f
C631 VTAIL.n488 B 0.024275f
C632 VTAIL.n489 B 0.024275f
C633 VTAIL.n490 B 0.010875f
C634 VTAIL.n491 B 0.01027f
C635 VTAIL.n492 B 0.019113f
C636 VTAIL.n493 B 0.019113f
C637 VTAIL.n494 B 0.01027f
C638 VTAIL.n495 B 0.010875f
C639 VTAIL.n496 B 0.024275f
C640 VTAIL.n497 B 0.024275f
C641 VTAIL.n498 B 0.010875f
C642 VTAIL.n499 B 0.01027f
C643 VTAIL.n500 B 0.019113f
C644 VTAIL.n501 B 0.019113f
C645 VTAIL.n502 B 0.01027f
C646 VTAIL.n503 B 0.010875f
C647 VTAIL.n504 B 0.024275f
C648 VTAIL.n505 B 0.024275f
C649 VTAIL.n506 B 0.010875f
C650 VTAIL.n507 B 0.01027f
C651 VTAIL.n508 B 0.019113f
C652 VTAIL.n509 B 0.019113f
C653 VTAIL.n510 B 0.01027f
C654 VTAIL.n511 B 0.010573f
C655 VTAIL.n512 B 0.010573f
C656 VTAIL.n513 B 0.024275f
C657 VTAIL.n514 B 0.024275f
C658 VTAIL.n515 B 0.010875f
C659 VTAIL.n516 B 0.01027f
C660 VTAIL.n517 B 0.019113f
C661 VTAIL.n518 B 0.019113f
C662 VTAIL.n519 B 0.01027f
C663 VTAIL.n520 B 0.010875f
C664 VTAIL.n521 B 0.024275f
C665 VTAIL.n522 B 0.024275f
C666 VTAIL.n523 B 0.010875f
C667 VTAIL.n524 B 0.01027f
C668 VTAIL.n525 B 0.019113f
C669 VTAIL.n526 B 0.019113f
C670 VTAIL.n527 B 0.01027f
C671 VTAIL.n528 B 0.010875f
C672 VTAIL.n529 B 0.024275f
C673 VTAIL.n530 B 0.05164f
C674 VTAIL.n531 B 0.010875f
C675 VTAIL.n532 B 0.01027f
C676 VTAIL.n533 B 0.04209f
C677 VTAIL.n534 B 0.028735f
C678 VTAIL.n535 B 0.269188f
C679 VTAIL.n536 B 0.026349f
C680 VTAIL.n537 B 0.019113f
C681 VTAIL.n538 B 0.01027f
C682 VTAIL.n539 B 0.024275f
C683 VTAIL.n540 B 0.010875f
C684 VTAIL.n541 B 0.019113f
C685 VTAIL.n542 B 0.01027f
C686 VTAIL.n543 B 0.024275f
C687 VTAIL.n544 B 0.010875f
C688 VTAIL.n545 B 0.019113f
C689 VTAIL.n546 B 0.01027f
C690 VTAIL.n547 B 0.024275f
C691 VTAIL.n548 B 0.010875f
C692 VTAIL.n549 B 0.019113f
C693 VTAIL.n550 B 0.01027f
C694 VTAIL.n551 B 0.024275f
C695 VTAIL.n552 B 0.024275f
C696 VTAIL.n553 B 0.010875f
C697 VTAIL.n554 B 0.019113f
C698 VTAIL.n555 B 0.01027f
C699 VTAIL.n556 B 0.024275f
C700 VTAIL.n557 B 0.010875f
C701 VTAIL.n558 B 0.019113f
C702 VTAIL.n559 B 0.01027f
C703 VTAIL.n560 B 0.024275f
C704 VTAIL.n561 B 0.010875f
C705 VTAIL.n562 B 0.019113f
C706 VTAIL.n563 B 0.01027f
C707 VTAIL.n564 B 0.024275f
C708 VTAIL.n565 B 0.010875f
C709 VTAIL.n566 B 0.019113f
C710 VTAIL.n567 B 0.01027f
C711 VTAIL.n568 B 0.024275f
C712 VTAIL.n569 B 0.010875f
C713 VTAIL.n570 B 0.143251f
C714 VTAIL.t14 B 0.040282f
C715 VTAIL.n571 B 0.018207f
C716 VTAIL.n572 B 0.01434f
C717 VTAIL.n573 B 0.01027f
C718 VTAIL.n574 B 1.58338f
C719 VTAIL.n575 B 0.019113f
C720 VTAIL.n576 B 0.01027f
C721 VTAIL.n577 B 0.010875f
C722 VTAIL.n578 B 0.024275f
C723 VTAIL.n579 B 0.024275f
C724 VTAIL.n580 B 0.010875f
C725 VTAIL.n581 B 0.01027f
C726 VTAIL.n582 B 0.019113f
C727 VTAIL.n583 B 0.019113f
C728 VTAIL.n584 B 0.01027f
C729 VTAIL.n585 B 0.010875f
C730 VTAIL.n586 B 0.024275f
C731 VTAIL.n587 B 0.024275f
C732 VTAIL.n588 B 0.010875f
C733 VTAIL.n589 B 0.01027f
C734 VTAIL.n590 B 0.019113f
C735 VTAIL.n591 B 0.019113f
C736 VTAIL.n592 B 0.01027f
C737 VTAIL.n593 B 0.010875f
C738 VTAIL.n594 B 0.024275f
C739 VTAIL.n595 B 0.024275f
C740 VTAIL.n596 B 0.010875f
C741 VTAIL.n597 B 0.01027f
C742 VTAIL.n598 B 0.019113f
C743 VTAIL.n599 B 0.019113f
C744 VTAIL.n600 B 0.01027f
C745 VTAIL.n601 B 0.010875f
C746 VTAIL.n602 B 0.024275f
C747 VTAIL.n603 B 0.024275f
C748 VTAIL.n604 B 0.010875f
C749 VTAIL.n605 B 0.01027f
C750 VTAIL.n606 B 0.019113f
C751 VTAIL.n607 B 0.019113f
C752 VTAIL.n608 B 0.01027f
C753 VTAIL.n609 B 0.010875f
C754 VTAIL.n610 B 0.024275f
C755 VTAIL.n611 B 0.024275f
C756 VTAIL.n612 B 0.010875f
C757 VTAIL.n613 B 0.01027f
C758 VTAIL.n614 B 0.019113f
C759 VTAIL.n615 B 0.019113f
C760 VTAIL.n616 B 0.01027f
C761 VTAIL.n617 B 0.010573f
C762 VTAIL.n618 B 0.010573f
C763 VTAIL.n619 B 0.024275f
C764 VTAIL.n620 B 0.024275f
C765 VTAIL.n621 B 0.010875f
C766 VTAIL.n622 B 0.01027f
C767 VTAIL.n623 B 0.019113f
C768 VTAIL.n624 B 0.019113f
C769 VTAIL.n625 B 0.01027f
C770 VTAIL.n626 B 0.010875f
C771 VTAIL.n627 B 0.024275f
C772 VTAIL.n628 B 0.024275f
C773 VTAIL.n629 B 0.010875f
C774 VTAIL.n630 B 0.01027f
C775 VTAIL.n631 B 0.019113f
C776 VTAIL.n632 B 0.019113f
C777 VTAIL.n633 B 0.01027f
C778 VTAIL.n634 B 0.010875f
C779 VTAIL.n635 B 0.024275f
C780 VTAIL.n636 B 0.05164f
C781 VTAIL.n637 B 0.010875f
C782 VTAIL.n638 B 0.01027f
C783 VTAIL.n639 B 0.04209f
C784 VTAIL.n640 B 0.028735f
C785 VTAIL.n641 B 0.269188f
C786 VTAIL.t1 B 0.285155f
C787 VTAIL.t0 B 0.285155f
C788 VTAIL.n642 B 2.53856f
C789 VTAIL.n643 B 0.647604f
C790 VTAIL.n644 B 0.026349f
C791 VTAIL.n645 B 0.019113f
C792 VTAIL.n646 B 0.01027f
C793 VTAIL.n647 B 0.024275f
C794 VTAIL.n648 B 0.010875f
C795 VTAIL.n649 B 0.019113f
C796 VTAIL.n650 B 0.01027f
C797 VTAIL.n651 B 0.024275f
C798 VTAIL.n652 B 0.010875f
C799 VTAIL.n653 B 0.019113f
C800 VTAIL.n654 B 0.01027f
C801 VTAIL.n655 B 0.024275f
C802 VTAIL.n656 B 0.010875f
C803 VTAIL.n657 B 0.019113f
C804 VTAIL.n658 B 0.01027f
C805 VTAIL.n659 B 0.024275f
C806 VTAIL.n660 B 0.024275f
C807 VTAIL.n661 B 0.010875f
C808 VTAIL.n662 B 0.019113f
C809 VTAIL.n663 B 0.01027f
C810 VTAIL.n664 B 0.024275f
C811 VTAIL.n665 B 0.010875f
C812 VTAIL.n666 B 0.019113f
C813 VTAIL.n667 B 0.01027f
C814 VTAIL.n668 B 0.024275f
C815 VTAIL.n669 B 0.010875f
C816 VTAIL.n670 B 0.019113f
C817 VTAIL.n671 B 0.01027f
C818 VTAIL.n672 B 0.024275f
C819 VTAIL.n673 B 0.010875f
C820 VTAIL.n674 B 0.019113f
C821 VTAIL.n675 B 0.01027f
C822 VTAIL.n676 B 0.024275f
C823 VTAIL.n677 B 0.010875f
C824 VTAIL.n678 B 0.143251f
C825 VTAIL.t12 B 0.040282f
C826 VTAIL.n679 B 0.018207f
C827 VTAIL.n680 B 0.01434f
C828 VTAIL.n681 B 0.01027f
C829 VTAIL.n682 B 1.58338f
C830 VTAIL.n683 B 0.019113f
C831 VTAIL.n684 B 0.01027f
C832 VTAIL.n685 B 0.010875f
C833 VTAIL.n686 B 0.024275f
C834 VTAIL.n687 B 0.024275f
C835 VTAIL.n688 B 0.010875f
C836 VTAIL.n689 B 0.01027f
C837 VTAIL.n690 B 0.019113f
C838 VTAIL.n691 B 0.019113f
C839 VTAIL.n692 B 0.01027f
C840 VTAIL.n693 B 0.010875f
C841 VTAIL.n694 B 0.024275f
C842 VTAIL.n695 B 0.024275f
C843 VTAIL.n696 B 0.010875f
C844 VTAIL.n697 B 0.01027f
C845 VTAIL.n698 B 0.019113f
C846 VTAIL.n699 B 0.019113f
C847 VTAIL.n700 B 0.01027f
C848 VTAIL.n701 B 0.010875f
C849 VTAIL.n702 B 0.024275f
C850 VTAIL.n703 B 0.024275f
C851 VTAIL.n704 B 0.010875f
C852 VTAIL.n705 B 0.01027f
C853 VTAIL.n706 B 0.019113f
C854 VTAIL.n707 B 0.019113f
C855 VTAIL.n708 B 0.01027f
C856 VTAIL.n709 B 0.010875f
C857 VTAIL.n710 B 0.024275f
C858 VTAIL.n711 B 0.024275f
C859 VTAIL.n712 B 0.010875f
C860 VTAIL.n713 B 0.01027f
C861 VTAIL.n714 B 0.019113f
C862 VTAIL.n715 B 0.019113f
C863 VTAIL.n716 B 0.01027f
C864 VTAIL.n717 B 0.010875f
C865 VTAIL.n718 B 0.024275f
C866 VTAIL.n719 B 0.024275f
C867 VTAIL.n720 B 0.010875f
C868 VTAIL.n721 B 0.01027f
C869 VTAIL.n722 B 0.019113f
C870 VTAIL.n723 B 0.019113f
C871 VTAIL.n724 B 0.01027f
C872 VTAIL.n725 B 0.010573f
C873 VTAIL.n726 B 0.010573f
C874 VTAIL.n727 B 0.024275f
C875 VTAIL.n728 B 0.024275f
C876 VTAIL.n729 B 0.010875f
C877 VTAIL.n730 B 0.01027f
C878 VTAIL.n731 B 0.019113f
C879 VTAIL.n732 B 0.019113f
C880 VTAIL.n733 B 0.01027f
C881 VTAIL.n734 B 0.010875f
C882 VTAIL.n735 B 0.024275f
C883 VTAIL.n736 B 0.024275f
C884 VTAIL.n737 B 0.010875f
C885 VTAIL.n738 B 0.01027f
C886 VTAIL.n739 B 0.019113f
C887 VTAIL.n740 B 0.019113f
C888 VTAIL.n741 B 0.01027f
C889 VTAIL.n742 B 0.010875f
C890 VTAIL.n743 B 0.024275f
C891 VTAIL.n744 B 0.05164f
C892 VTAIL.n745 B 0.010875f
C893 VTAIL.n746 B 0.01027f
C894 VTAIL.n747 B 0.04209f
C895 VTAIL.n748 B 0.028735f
C896 VTAIL.n749 B 1.72735f
C897 VTAIL.n750 B 0.026349f
C898 VTAIL.n751 B 0.019113f
C899 VTAIL.n752 B 0.01027f
C900 VTAIL.n753 B 0.024275f
C901 VTAIL.n754 B 0.010875f
C902 VTAIL.n755 B 0.019113f
C903 VTAIL.n756 B 0.01027f
C904 VTAIL.n757 B 0.024275f
C905 VTAIL.n758 B 0.010875f
C906 VTAIL.n759 B 0.019113f
C907 VTAIL.n760 B 0.01027f
C908 VTAIL.n761 B 0.024275f
C909 VTAIL.n762 B 0.010875f
C910 VTAIL.n763 B 0.019113f
C911 VTAIL.n764 B 0.01027f
C912 VTAIL.n765 B 0.024275f
C913 VTAIL.n766 B 0.010875f
C914 VTAIL.n767 B 0.019113f
C915 VTAIL.n768 B 0.01027f
C916 VTAIL.n769 B 0.024275f
C917 VTAIL.n770 B 0.010875f
C918 VTAIL.n771 B 0.019113f
C919 VTAIL.n772 B 0.01027f
C920 VTAIL.n773 B 0.024275f
C921 VTAIL.n774 B 0.010875f
C922 VTAIL.n775 B 0.019113f
C923 VTAIL.n776 B 0.01027f
C924 VTAIL.n777 B 0.024275f
C925 VTAIL.n778 B 0.010875f
C926 VTAIL.n779 B 0.019113f
C927 VTAIL.n780 B 0.01027f
C928 VTAIL.n781 B 0.024275f
C929 VTAIL.n782 B 0.010875f
C930 VTAIL.n783 B 0.143251f
C931 VTAIL.t5 B 0.040282f
C932 VTAIL.n784 B 0.018207f
C933 VTAIL.n785 B 0.01434f
C934 VTAIL.n786 B 0.01027f
C935 VTAIL.n787 B 1.58338f
C936 VTAIL.n788 B 0.019113f
C937 VTAIL.n789 B 0.01027f
C938 VTAIL.n790 B 0.010875f
C939 VTAIL.n791 B 0.024275f
C940 VTAIL.n792 B 0.024275f
C941 VTAIL.n793 B 0.010875f
C942 VTAIL.n794 B 0.01027f
C943 VTAIL.n795 B 0.019113f
C944 VTAIL.n796 B 0.019113f
C945 VTAIL.n797 B 0.01027f
C946 VTAIL.n798 B 0.010875f
C947 VTAIL.n799 B 0.024275f
C948 VTAIL.n800 B 0.024275f
C949 VTAIL.n801 B 0.010875f
C950 VTAIL.n802 B 0.01027f
C951 VTAIL.n803 B 0.019113f
C952 VTAIL.n804 B 0.019113f
C953 VTAIL.n805 B 0.01027f
C954 VTAIL.n806 B 0.010875f
C955 VTAIL.n807 B 0.024275f
C956 VTAIL.n808 B 0.024275f
C957 VTAIL.n809 B 0.010875f
C958 VTAIL.n810 B 0.01027f
C959 VTAIL.n811 B 0.019113f
C960 VTAIL.n812 B 0.019113f
C961 VTAIL.n813 B 0.01027f
C962 VTAIL.n814 B 0.010875f
C963 VTAIL.n815 B 0.024275f
C964 VTAIL.n816 B 0.024275f
C965 VTAIL.n817 B 0.010875f
C966 VTAIL.n818 B 0.01027f
C967 VTAIL.n819 B 0.019113f
C968 VTAIL.n820 B 0.019113f
C969 VTAIL.n821 B 0.01027f
C970 VTAIL.n822 B 0.010875f
C971 VTAIL.n823 B 0.024275f
C972 VTAIL.n824 B 0.024275f
C973 VTAIL.n825 B 0.024275f
C974 VTAIL.n826 B 0.010875f
C975 VTAIL.n827 B 0.01027f
C976 VTAIL.n828 B 0.019113f
C977 VTAIL.n829 B 0.019113f
C978 VTAIL.n830 B 0.01027f
C979 VTAIL.n831 B 0.010573f
C980 VTAIL.n832 B 0.010573f
C981 VTAIL.n833 B 0.024275f
C982 VTAIL.n834 B 0.024275f
C983 VTAIL.n835 B 0.010875f
C984 VTAIL.n836 B 0.01027f
C985 VTAIL.n837 B 0.019113f
C986 VTAIL.n838 B 0.019113f
C987 VTAIL.n839 B 0.01027f
C988 VTAIL.n840 B 0.010875f
C989 VTAIL.n841 B 0.024275f
C990 VTAIL.n842 B 0.024275f
C991 VTAIL.n843 B 0.010875f
C992 VTAIL.n844 B 0.01027f
C993 VTAIL.n845 B 0.019113f
C994 VTAIL.n846 B 0.019113f
C995 VTAIL.n847 B 0.01027f
C996 VTAIL.n848 B 0.010875f
C997 VTAIL.n849 B 0.024275f
C998 VTAIL.n850 B 0.05164f
C999 VTAIL.n851 B 0.010875f
C1000 VTAIL.n852 B 0.01027f
C1001 VTAIL.n853 B 0.04209f
C1002 VTAIL.n854 B 0.028735f
C1003 VTAIL.n855 B 1.72376f
C1004 VDD2.t4 B 0.393226f
C1005 VDD2.t0 B 0.393226f
C1006 VDD2.n0 B 3.60643f
C1007 VDD2.t7 B 0.393226f
C1008 VDD2.t2 B 0.393226f
C1009 VDD2.n1 B 3.60643f
C1010 VDD2.n2 B 4.72544f
C1011 VDD2.t5 B 0.393226f
C1012 VDD2.t1 B 0.393226f
C1013 VDD2.n3 B 3.5862f
C1014 VDD2.n4 B 4.13929f
C1015 VDD2.t3 B 0.393226f
C1016 VDD2.t6 B 0.393226f
C1017 VDD2.n5 B 3.60637f
C1018 VN.n0 B 0.029751f
C1019 VN.t5 B 3.21535f
C1020 VN.n1 B 0.029339f
C1021 VN.n2 B 0.015821f
C1022 VN.n3 B 0.029339f
C1023 VN.n4 B 0.015821f
C1024 VN.t0 B 3.21535f
C1025 VN.n5 B 0.029339f
C1026 VN.n6 B 0.015821f
C1027 VN.n7 B 0.029339f
C1028 VN.n8 B 0.211093f
C1029 VN.t7 B 3.21535f
C1030 VN.t1 B 3.48259f
C1031 VN.n9 B 1.10603f
C1032 VN.n10 B 1.15884f
C1033 VN.n11 B 0.018331f
C1034 VN.n12 B 0.029339f
C1035 VN.n13 B 0.015821f
C1036 VN.n14 B 0.015821f
C1037 VN.n15 B 0.015821f
C1038 VN.n16 B 0.031279f
C1039 VN.n17 B 0.012778f
C1040 VN.n18 B 0.031279f
C1041 VN.n19 B 0.015821f
C1042 VN.n20 B 0.015821f
C1043 VN.n21 B 0.015821f
C1044 VN.n22 B 0.029339f
C1045 VN.n23 B 0.018331f
C1046 VN.n24 B 1.10553f
C1047 VN.n25 B 0.025863f
C1048 VN.n26 B 0.015821f
C1049 VN.n27 B 0.015821f
C1050 VN.n28 B 0.015821f
C1051 VN.n29 B 0.029339f
C1052 VN.n30 B 0.022561f
C1053 VN.n31 B 0.023437f
C1054 VN.n32 B 0.015821f
C1055 VN.n33 B 0.015821f
C1056 VN.n34 B 0.015821f
C1057 VN.n35 B 0.029339f
C1058 VN.n36 B 0.025284f
C1059 VN.n37 B 1.17088f
C1060 VN.n38 B 0.052015f
C1061 VN.n39 B 0.029751f
C1062 VN.t4 B 3.21535f
C1063 VN.n40 B 0.029339f
C1064 VN.n41 B 0.015821f
C1065 VN.n42 B 0.029339f
C1066 VN.n43 B 0.015821f
C1067 VN.t6 B 3.21535f
C1068 VN.n44 B 0.029339f
C1069 VN.n45 B 0.015821f
C1070 VN.n46 B 0.029339f
C1071 VN.n47 B 0.211093f
C1072 VN.t2 B 3.21535f
C1073 VN.t3 B 3.48259f
C1074 VN.n48 B 1.10603f
C1075 VN.n49 B 1.15884f
C1076 VN.n50 B 0.018331f
C1077 VN.n51 B 0.029339f
C1078 VN.n52 B 0.015821f
C1079 VN.n53 B 0.015821f
C1080 VN.n54 B 0.015821f
C1081 VN.n55 B 0.031279f
C1082 VN.n56 B 0.012778f
C1083 VN.n57 B 0.031279f
C1084 VN.n58 B 0.015821f
C1085 VN.n59 B 0.015821f
C1086 VN.n60 B 0.015821f
C1087 VN.n61 B 0.029339f
C1088 VN.n62 B 0.018331f
C1089 VN.n63 B 1.10553f
C1090 VN.n64 B 0.025863f
C1091 VN.n65 B 0.015821f
C1092 VN.n66 B 0.015821f
C1093 VN.n67 B 0.015821f
C1094 VN.n68 B 0.029339f
C1095 VN.n69 B 0.022561f
C1096 VN.n70 B 0.023437f
C1097 VN.n71 B 0.015821f
C1098 VN.n72 B 0.015821f
C1099 VN.n73 B 0.015821f
C1100 VN.n74 B 0.029339f
C1101 VN.n75 B 0.025284f
C1102 VN.n76 B 1.17088f
C1103 VN.n77 B 1.24589f
.ends

