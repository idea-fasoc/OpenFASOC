* NGSPICE file created from diff_pair_sample_0354.ext - technology: sky130A

.subckt diff_pair_sample_0354 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=7.6011 ps=39.76 w=19.49 l=2.9
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=0 ps=0 w=19.49 l=2.9
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=0 ps=0 w=19.49 l=2.9
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=7.6011 ps=39.76 w=19.49 l=2.9
X4 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=7.6011 ps=39.76 w=19.49 l=2.9
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=0 ps=0 w=19.49 l=2.9
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=7.6011 ps=39.76 w=19.49 l=2.9
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6011 pd=39.76 as=0 ps=0 w=19.49 l=2.9
R0 VP.n0 VP.t0 254.191
R1 VP.n0 VP.t1 203.065
R2 VP VP.n0 0.431811
R3 VTAIL.n418 VTAIL.n318 214.453
R4 VTAIL.n100 VTAIL.n0 214.453
R5 VTAIL.n312 VTAIL.n212 214.453
R6 VTAIL.n206 VTAIL.n106 214.453
R7 VTAIL.n353 VTAIL.n352 185
R8 VTAIL.n350 VTAIL.n349 185
R9 VTAIL.n359 VTAIL.n358 185
R10 VTAIL.n361 VTAIL.n360 185
R11 VTAIL.n346 VTAIL.n345 185
R12 VTAIL.n367 VTAIL.n366 185
R13 VTAIL.n370 VTAIL.n369 185
R14 VTAIL.n368 VTAIL.n342 185
R15 VTAIL.n375 VTAIL.n341 185
R16 VTAIL.n377 VTAIL.n376 185
R17 VTAIL.n379 VTAIL.n378 185
R18 VTAIL.n338 VTAIL.n337 185
R19 VTAIL.n385 VTAIL.n384 185
R20 VTAIL.n387 VTAIL.n386 185
R21 VTAIL.n334 VTAIL.n333 185
R22 VTAIL.n393 VTAIL.n392 185
R23 VTAIL.n395 VTAIL.n394 185
R24 VTAIL.n330 VTAIL.n329 185
R25 VTAIL.n401 VTAIL.n400 185
R26 VTAIL.n403 VTAIL.n402 185
R27 VTAIL.n326 VTAIL.n325 185
R28 VTAIL.n409 VTAIL.n408 185
R29 VTAIL.n411 VTAIL.n410 185
R30 VTAIL.n322 VTAIL.n321 185
R31 VTAIL.n417 VTAIL.n416 185
R32 VTAIL.n419 VTAIL.n418 185
R33 VTAIL.n35 VTAIL.n34 185
R34 VTAIL.n32 VTAIL.n31 185
R35 VTAIL.n41 VTAIL.n40 185
R36 VTAIL.n43 VTAIL.n42 185
R37 VTAIL.n28 VTAIL.n27 185
R38 VTAIL.n49 VTAIL.n48 185
R39 VTAIL.n52 VTAIL.n51 185
R40 VTAIL.n50 VTAIL.n24 185
R41 VTAIL.n57 VTAIL.n23 185
R42 VTAIL.n59 VTAIL.n58 185
R43 VTAIL.n61 VTAIL.n60 185
R44 VTAIL.n20 VTAIL.n19 185
R45 VTAIL.n67 VTAIL.n66 185
R46 VTAIL.n69 VTAIL.n68 185
R47 VTAIL.n16 VTAIL.n15 185
R48 VTAIL.n75 VTAIL.n74 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n12 VTAIL.n11 185
R51 VTAIL.n83 VTAIL.n82 185
R52 VTAIL.n85 VTAIL.n84 185
R53 VTAIL.n8 VTAIL.n7 185
R54 VTAIL.n91 VTAIL.n90 185
R55 VTAIL.n93 VTAIL.n92 185
R56 VTAIL.n4 VTAIL.n3 185
R57 VTAIL.n99 VTAIL.n98 185
R58 VTAIL.n101 VTAIL.n100 185
R59 VTAIL.n313 VTAIL.n312 185
R60 VTAIL.n311 VTAIL.n310 185
R61 VTAIL.n216 VTAIL.n215 185
R62 VTAIL.n305 VTAIL.n304 185
R63 VTAIL.n303 VTAIL.n302 185
R64 VTAIL.n220 VTAIL.n219 185
R65 VTAIL.n297 VTAIL.n296 185
R66 VTAIL.n295 VTAIL.n294 185
R67 VTAIL.n224 VTAIL.n223 185
R68 VTAIL.n289 VTAIL.n288 185
R69 VTAIL.n287 VTAIL.n286 185
R70 VTAIL.n228 VTAIL.n227 185
R71 VTAIL.n281 VTAIL.n280 185
R72 VTAIL.n279 VTAIL.n278 185
R73 VTAIL.n232 VTAIL.n231 185
R74 VTAIL.n273 VTAIL.n272 185
R75 VTAIL.n271 VTAIL.n270 185
R76 VTAIL.n269 VTAIL.n235 185
R77 VTAIL.n239 VTAIL.n236 185
R78 VTAIL.n264 VTAIL.n263 185
R79 VTAIL.n262 VTAIL.n261 185
R80 VTAIL.n241 VTAIL.n240 185
R81 VTAIL.n256 VTAIL.n255 185
R82 VTAIL.n254 VTAIL.n253 185
R83 VTAIL.n245 VTAIL.n244 185
R84 VTAIL.n248 VTAIL.n247 185
R85 VTAIL.n207 VTAIL.n206 185
R86 VTAIL.n205 VTAIL.n204 185
R87 VTAIL.n110 VTAIL.n109 185
R88 VTAIL.n199 VTAIL.n198 185
R89 VTAIL.n197 VTAIL.n196 185
R90 VTAIL.n114 VTAIL.n113 185
R91 VTAIL.n191 VTAIL.n190 185
R92 VTAIL.n189 VTAIL.n188 185
R93 VTAIL.n118 VTAIL.n117 185
R94 VTAIL.n183 VTAIL.n182 185
R95 VTAIL.n181 VTAIL.n180 185
R96 VTAIL.n122 VTAIL.n121 185
R97 VTAIL.n175 VTAIL.n174 185
R98 VTAIL.n173 VTAIL.n172 185
R99 VTAIL.n126 VTAIL.n125 185
R100 VTAIL.n167 VTAIL.n166 185
R101 VTAIL.n165 VTAIL.n164 185
R102 VTAIL.n163 VTAIL.n129 185
R103 VTAIL.n133 VTAIL.n130 185
R104 VTAIL.n158 VTAIL.n157 185
R105 VTAIL.n156 VTAIL.n155 185
R106 VTAIL.n135 VTAIL.n134 185
R107 VTAIL.n150 VTAIL.n149 185
R108 VTAIL.n148 VTAIL.n147 185
R109 VTAIL.n139 VTAIL.n138 185
R110 VTAIL.n142 VTAIL.n141 185
R111 VTAIL.t0 VTAIL.n351 149.524
R112 VTAIL.t3 VTAIL.n33 149.524
R113 VTAIL.t2 VTAIL.n246 149.524
R114 VTAIL.t1 VTAIL.n140 149.524
R115 VTAIL.n352 VTAIL.n349 104.615
R116 VTAIL.n359 VTAIL.n349 104.615
R117 VTAIL.n360 VTAIL.n359 104.615
R118 VTAIL.n360 VTAIL.n345 104.615
R119 VTAIL.n367 VTAIL.n345 104.615
R120 VTAIL.n369 VTAIL.n367 104.615
R121 VTAIL.n369 VTAIL.n368 104.615
R122 VTAIL.n368 VTAIL.n341 104.615
R123 VTAIL.n377 VTAIL.n341 104.615
R124 VTAIL.n378 VTAIL.n377 104.615
R125 VTAIL.n378 VTAIL.n337 104.615
R126 VTAIL.n385 VTAIL.n337 104.615
R127 VTAIL.n386 VTAIL.n385 104.615
R128 VTAIL.n386 VTAIL.n333 104.615
R129 VTAIL.n393 VTAIL.n333 104.615
R130 VTAIL.n394 VTAIL.n393 104.615
R131 VTAIL.n394 VTAIL.n329 104.615
R132 VTAIL.n401 VTAIL.n329 104.615
R133 VTAIL.n402 VTAIL.n401 104.615
R134 VTAIL.n402 VTAIL.n325 104.615
R135 VTAIL.n409 VTAIL.n325 104.615
R136 VTAIL.n410 VTAIL.n409 104.615
R137 VTAIL.n410 VTAIL.n321 104.615
R138 VTAIL.n417 VTAIL.n321 104.615
R139 VTAIL.n418 VTAIL.n417 104.615
R140 VTAIL.n34 VTAIL.n31 104.615
R141 VTAIL.n41 VTAIL.n31 104.615
R142 VTAIL.n42 VTAIL.n41 104.615
R143 VTAIL.n42 VTAIL.n27 104.615
R144 VTAIL.n49 VTAIL.n27 104.615
R145 VTAIL.n51 VTAIL.n49 104.615
R146 VTAIL.n51 VTAIL.n50 104.615
R147 VTAIL.n50 VTAIL.n23 104.615
R148 VTAIL.n59 VTAIL.n23 104.615
R149 VTAIL.n60 VTAIL.n59 104.615
R150 VTAIL.n60 VTAIL.n19 104.615
R151 VTAIL.n67 VTAIL.n19 104.615
R152 VTAIL.n68 VTAIL.n67 104.615
R153 VTAIL.n68 VTAIL.n15 104.615
R154 VTAIL.n75 VTAIL.n15 104.615
R155 VTAIL.n76 VTAIL.n75 104.615
R156 VTAIL.n76 VTAIL.n11 104.615
R157 VTAIL.n83 VTAIL.n11 104.615
R158 VTAIL.n84 VTAIL.n83 104.615
R159 VTAIL.n84 VTAIL.n7 104.615
R160 VTAIL.n91 VTAIL.n7 104.615
R161 VTAIL.n92 VTAIL.n91 104.615
R162 VTAIL.n92 VTAIL.n3 104.615
R163 VTAIL.n99 VTAIL.n3 104.615
R164 VTAIL.n100 VTAIL.n99 104.615
R165 VTAIL.n312 VTAIL.n311 104.615
R166 VTAIL.n311 VTAIL.n215 104.615
R167 VTAIL.n304 VTAIL.n215 104.615
R168 VTAIL.n304 VTAIL.n303 104.615
R169 VTAIL.n303 VTAIL.n219 104.615
R170 VTAIL.n296 VTAIL.n219 104.615
R171 VTAIL.n296 VTAIL.n295 104.615
R172 VTAIL.n295 VTAIL.n223 104.615
R173 VTAIL.n288 VTAIL.n223 104.615
R174 VTAIL.n288 VTAIL.n287 104.615
R175 VTAIL.n287 VTAIL.n227 104.615
R176 VTAIL.n280 VTAIL.n227 104.615
R177 VTAIL.n280 VTAIL.n279 104.615
R178 VTAIL.n279 VTAIL.n231 104.615
R179 VTAIL.n272 VTAIL.n231 104.615
R180 VTAIL.n272 VTAIL.n271 104.615
R181 VTAIL.n271 VTAIL.n235 104.615
R182 VTAIL.n239 VTAIL.n235 104.615
R183 VTAIL.n263 VTAIL.n239 104.615
R184 VTAIL.n263 VTAIL.n262 104.615
R185 VTAIL.n262 VTAIL.n240 104.615
R186 VTAIL.n255 VTAIL.n240 104.615
R187 VTAIL.n255 VTAIL.n254 104.615
R188 VTAIL.n254 VTAIL.n244 104.615
R189 VTAIL.n247 VTAIL.n244 104.615
R190 VTAIL.n206 VTAIL.n205 104.615
R191 VTAIL.n205 VTAIL.n109 104.615
R192 VTAIL.n198 VTAIL.n109 104.615
R193 VTAIL.n198 VTAIL.n197 104.615
R194 VTAIL.n197 VTAIL.n113 104.615
R195 VTAIL.n190 VTAIL.n113 104.615
R196 VTAIL.n190 VTAIL.n189 104.615
R197 VTAIL.n189 VTAIL.n117 104.615
R198 VTAIL.n182 VTAIL.n117 104.615
R199 VTAIL.n182 VTAIL.n181 104.615
R200 VTAIL.n181 VTAIL.n121 104.615
R201 VTAIL.n174 VTAIL.n121 104.615
R202 VTAIL.n174 VTAIL.n173 104.615
R203 VTAIL.n173 VTAIL.n125 104.615
R204 VTAIL.n166 VTAIL.n125 104.615
R205 VTAIL.n166 VTAIL.n165 104.615
R206 VTAIL.n165 VTAIL.n129 104.615
R207 VTAIL.n133 VTAIL.n129 104.615
R208 VTAIL.n157 VTAIL.n133 104.615
R209 VTAIL.n157 VTAIL.n156 104.615
R210 VTAIL.n156 VTAIL.n134 104.615
R211 VTAIL.n149 VTAIL.n134 104.615
R212 VTAIL.n149 VTAIL.n148 104.615
R213 VTAIL.n148 VTAIL.n138 104.615
R214 VTAIL.n141 VTAIL.n138 104.615
R215 VTAIL.n352 VTAIL.t0 52.3082
R216 VTAIL.n34 VTAIL.t3 52.3082
R217 VTAIL.n247 VTAIL.t2 52.3082
R218 VTAIL.n141 VTAIL.t1 52.3082
R219 VTAIL.n423 VTAIL.n422 35.4823
R220 VTAIL.n105 VTAIL.n104 35.4823
R221 VTAIL.n317 VTAIL.n316 35.4823
R222 VTAIL.n211 VTAIL.n210 35.4823
R223 VTAIL.n211 VTAIL.n105 34.7376
R224 VTAIL.n423 VTAIL.n317 31.9531
R225 VTAIL.n376 VTAIL.n375 13.1884
R226 VTAIL.n58 VTAIL.n57 13.1884
R227 VTAIL.n270 VTAIL.n269 13.1884
R228 VTAIL.n164 VTAIL.n163 13.1884
R229 VTAIL.n374 VTAIL.n342 12.8005
R230 VTAIL.n379 VTAIL.n340 12.8005
R231 VTAIL.n420 VTAIL.n419 12.8005
R232 VTAIL.n56 VTAIL.n24 12.8005
R233 VTAIL.n61 VTAIL.n22 12.8005
R234 VTAIL.n102 VTAIL.n101 12.8005
R235 VTAIL.n314 VTAIL.n313 12.8005
R236 VTAIL.n273 VTAIL.n234 12.8005
R237 VTAIL.n268 VTAIL.n236 12.8005
R238 VTAIL.n208 VTAIL.n207 12.8005
R239 VTAIL.n167 VTAIL.n128 12.8005
R240 VTAIL.n162 VTAIL.n130 12.8005
R241 VTAIL.n371 VTAIL.n370 12.0247
R242 VTAIL.n380 VTAIL.n338 12.0247
R243 VTAIL.n416 VTAIL.n320 12.0247
R244 VTAIL.n53 VTAIL.n52 12.0247
R245 VTAIL.n62 VTAIL.n20 12.0247
R246 VTAIL.n98 VTAIL.n2 12.0247
R247 VTAIL.n310 VTAIL.n214 12.0247
R248 VTAIL.n274 VTAIL.n232 12.0247
R249 VTAIL.n265 VTAIL.n264 12.0247
R250 VTAIL.n204 VTAIL.n108 12.0247
R251 VTAIL.n168 VTAIL.n126 12.0247
R252 VTAIL.n159 VTAIL.n158 12.0247
R253 VTAIL.n366 VTAIL.n344 11.249
R254 VTAIL.n384 VTAIL.n383 11.249
R255 VTAIL.n415 VTAIL.n322 11.249
R256 VTAIL.n48 VTAIL.n26 11.249
R257 VTAIL.n66 VTAIL.n65 11.249
R258 VTAIL.n97 VTAIL.n4 11.249
R259 VTAIL.n309 VTAIL.n216 11.249
R260 VTAIL.n278 VTAIL.n277 11.249
R261 VTAIL.n261 VTAIL.n238 11.249
R262 VTAIL.n203 VTAIL.n110 11.249
R263 VTAIL.n172 VTAIL.n171 11.249
R264 VTAIL.n155 VTAIL.n132 11.249
R265 VTAIL.n365 VTAIL.n346 10.4732
R266 VTAIL.n387 VTAIL.n336 10.4732
R267 VTAIL.n412 VTAIL.n411 10.4732
R268 VTAIL.n47 VTAIL.n28 10.4732
R269 VTAIL.n69 VTAIL.n18 10.4732
R270 VTAIL.n94 VTAIL.n93 10.4732
R271 VTAIL.n306 VTAIL.n305 10.4732
R272 VTAIL.n281 VTAIL.n230 10.4732
R273 VTAIL.n260 VTAIL.n241 10.4732
R274 VTAIL.n200 VTAIL.n199 10.4732
R275 VTAIL.n175 VTAIL.n124 10.4732
R276 VTAIL.n154 VTAIL.n135 10.4732
R277 VTAIL.n353 VTAIL.n351 10.2747
R278 VTAIL.n35 VTAIL.n33 10.2747
R279 VTAIL.n248 VTAIL.n246 10.2747
R280 VTAIL.n142 VTAIL.n140 10.2747
R281 VTAIL.n362 VTAIL.n361 9.69747
R282 VTAIL.n388 VTAIL.n334 9.69747
R283 VTAIL.n408 VTAIL.n324 9.69747
R284 VTAIL.n44 VTAIL.n43 9.69747
R285 VTAIL.n70 VTAIL.n16 9.69747
R286 VTAIL.n90 VTAIL.n6 9.69747
R287 VTAIL.n302 VTAIL.n218 9.69747
R288 VTAIL.n282 VTAIL.n228 9.69747
R289 VTAIL.n257 VTAIL.n256 9.69747
R290 VTAIL.n196 VTAIL.n112 9.69747
R291 VTAIL.n176 VTAIL.n122 9.69747
R292 VTAIL.n151 VTAIL.n150 9.69747
R293 VTAIL.n422 VTAIL.n421 9.45567
R294 VTAIL.n104 VTAIL.n103 9.45567
R295 VTAIL.n316 VTAIL.n315 9.45567
R296 VTAIL.n210 VTAIL.n209 9.45567
R297 VTAIL.n397 VTAIL.n396 9.3005
R298 VTAIL.n332 VTAIL.n331 9.3005
R299 VTAIL.n391 VTAIL.n390 9.3005
R300 VTAIL.n389 VTAIL.n388 9.3005
R301 VTAIL.n336 VTAIL.n335 9.3005
R302 VTAIL.n383 VTAIL.n382 9.3005
R303 VTAIL.n381 VTAIL.n380 9.3005
R304 VTAIL.n340 VTAIL.n339 9.3005
R305 VTAIL.n355 VTAIL.n354 9.3005
R306 VTAIL.n357 VTAIL.n356 9.3005
R307 VTAIL.n348 VTAIL.n347 9.3005
R308 VTAIL.n363 VTAIL.n362 9.3005
R309 VTAIL.n365 VTAIL.n364 9.3005
R310 VTAIL.n344 VTAIL.n343 9.3005
R311 VTAIL.n372 VTAIL.n371 9.3005
R312 VTAIL.n374 VTAIL.n373 9.3005
R313 VTAIL.n399 VTAIL.n398 9.3005
R314 VTAIL.n328 VTAIL.n327 9.3005
R315 VTAIL.n405 VTAIL.n404 9.3005
R316 VTAIL.n407 VTAIL.n406 9.3005
R317 VTAIL.n324 VTAIL.n323 9.3005
R318 VTAIL.n413 VTAIL.n412 9.3005
R319 VTAIL.n415 VTAIL.n414 9.3005
R320 VTAIL.n320 VTAIL.n319 9.3005
R321 VTAIL.n421 VTAIL.n420 9.3005
R322 VTAIL.n79 VTAIL.n78 9.3005
R323 VTAIL.n14 VTAIL.n13 9.3005
R324 VTAIL.n73 VTAIL.n72 9.3005
R325 VTAIL.n71 VTAIL.n70 9.3005
R326 VTAIL.n18 VTAIL.n17 9.3005
R327 VTAIL.n65 VTAIL.n64 9.3005
R328 VTAIL.n63 VTAIL.n62 9.3005
R329 VTAIL.n22 VTAIL.n21 9.3005
R330 VTAIL.n37 VTAIL.n36 9.3005
R331 VTAIL.n39 VTAIL.n38 9.3005
R332 VTAIL.n30 VTAIL.n29 9.3005
R333 VTAIL.n45 VTAIL.n44 9.3005
R334 VTAIL.n47 VTAIL.n46 9.3005
R335 VTAIL.n26 VTAIL.n25 9.3005
R336 VTAIL.n54 VTAIL.n53 9.3005
R337 VTAIL.n56 VTAIL.n55 9.3005
R338 VTAIL.n81 VTAIL.n80 9.3005
R339 VTAIL.n10 VTAIL.n9 9.3005
R340 VTAIL.n87 VTAIL.n86 9.3005
R341 VTAIL.n89 VTAIL.n88 9.3005
R342 VTAIL.n6 VTAIL.n5 9.3005
R343 VTAIL.n95 VTAIL.n94 9.3005
R344 VTAIL.n97 VTAIL.n96 9.3005
R345 VTAIL.n2 VTAIL.n1 9.3005
R346 VTAIL.n103 VTAIL.n102 9.3005
R347 VTAIL.n250 VTAIL.n249 9.3005
R348 VTAIL.n252 VTAIL.n251 9.3005
R349 VTAIL.n243 VTAIL.n242 9.3005
R350 VTAIL.n258 VTAIL.n257 9.3005
R351 VTAIL.n260 VTAIL.n259 9.3005
R352 VTAIL.n238 VTAIL.n237 9.3005
R353 VTAIL.n266 VTAIL.n265 9.3005
R354 VTAIL.n268 VTAIL.n267 9.3005
R355 VTAIL.n222 VTAIL.n221 9.3005
R356 VTAIL.n299 VTAIL.n298 9.3005
R357 VTAIL.n301 VTAIL.n300 9.3005
R358 VTAIL.n218 VTAIL.n217 9.3005
R359 VTAIL.n307 VTAIL.n306 9.3005
R360 VTAIL.n309 VTAIL.n308 9.3005
R361 VTAIL.n214 VTAIL.n213 9.3005
R362 VTAIL.n315 VTAIL.n314 9.3005
R363 VTAIL.n293 VTAIL.n292 9.3005
R364 VTAIL.n291 VTAIL.n290 9.3005
R365 VTAIL.n226 VTAIL.n225 9.3005
R366 VTAIL.n285 VTAIL.n284 9.3005
R367 VTAIL.n283 VTAIL.n282 9.3005
R368 VTAIL.n230 VTAIL.n229 9.3005
R369 VTAIL.n277 VTAIL.n276 9.3005
R370 VTAIL.n275 VTAIL.n274 9.3005
R371 VTAIL.n234 VTAIL.n233 9.3005
R372 VTAIL.n144 VTAIL.n143 9.3005
R373 VTAIL.n146 VTAIL.n145 9.3005
R374 VTAIL.n137 VTAIL.n136 9.3005
R375 VTAIL.n152 VTAIL.n151 9.3005
R376 VTAIL.n154 VTAIL.n153 9.3005
R377 VTAIL.n132 VTAIL.n131 9.3005
R378 VTAIL.n160 VTAIL.n159 9.3005
R379 VTAIL.n162 VTAIL.n161 9.3005
R380 VTAIL.n116 VTAIL.n115 9.3005
R381 VTAIL.n193 VTAIL.n192 9.3005
R382 VTAIL.n195 VTAIL.n194 9.3005
R383 VTAIL.n112 VTAIL.n111 9.3005
R384 VTAIL.n201 VTAIL.n200 9.3005
R385 VTAIL.n203 VTAIL.n202 9.3005
R386 VTAIL.n108 VTAIL.n107 9.3005
R387 VTAIL.n209 VTAIL.n208 9.3005
R388 VTAIL.n187 VTAIL.n186 9.3005
R389 VTAIL.n185 VTAIL.n184 9.3005
R390 VTAIL.n120 VTAIL.n119 9.3005
R391 VTAIL.n179 VTAIL.n178 9.3005
R392 VTAIL.n177 VTAIL.n176 9.3005
R393 VTAIL.n124 VTAIL.n123 9.3005
R394 VTAIL.n171 VTAIL.n170 9.3005
R395 VTAIL.n169 VTAIL.n168 9.3005
R396 VTAIL.n128 VTAIL.n127 9.3005
R397 VTAIL.n358 VTAIL.n348 8.92171
R398 VTAIL.n392 VTAIL.n391 8.92171
R399 VTAIL.n407 VTAIL.n326 8.92171
R400 VTAIL.n40 VTAIL.n30 8.92171
R401 VTAIL.n74 VTAIL.n73 8.92171
R402 VTAIL.n89 VTAIL.n8 8.92171
R403 VTAIL.n301 VTAIL.n220 8.92171
R404 VTAIL.n286 VTAIL.n285 8.92171
R405 VTAIL.n253 VTAIL.n243 8.92171
R406 VTAIL.n195 VTAIL.n114 8.92171
R407 VTAIL.n180 VTAIL.n179 8.92171
R408 VTAIL.n147 VTAIL.n137 8.92171
R409 VTAIL.n422 VTAIL.n318 8.2187
R410 VTAIL.n104 VTAIL.n0 8.2187
R411 VTAIL.n316 VTAIL.n212 8.2187
R412 VTAIL.n210 VTAIL.n106 8.2187
R413 VTAIL.n357 VTAIL.n350 8.14595
R414 VTAIL.n395 VTAIL.n332 8.14595
R415 VTAIL.n404 VTAIL.n403 8.14595
R416 VTAIL.n39 VTAIL.n32 8.14595
R417 VTAIL.n77 VTAIL.n14 8.14595
R418 VTAIL.n86 VTAIL.n85 8.14595
R419 VTAIL.n298 VTAIL.n297 8.14595
R420 VTAIL.n289 VTAIL.n226 8.14595
R421 VTAIL.n252 VTAIL.n245 8.14595
R422 VTAIL.n192 VTAIL.n191 8.14595
R423 VTAIL.n183 VTAIL.n120 8.14595
R424 VTAIL.n146 VTAIL.n139 8.14595
R425 VTAIL.n354 VTAIL.n353 7.3702
R426 VTAIL.n396 VTAIL.n330 7.3702
R427 VTAIL.n400 VTAIL.n328 7.3702
R428 VTAIL.n36 VTAIL.n35 7.3702
R429 VTAIL.n78 VTAIL.n12 7.3702
R430 VTAIL.n82 VTAIL.n10 7.3702
R431 VTAIL.n294 VTAIL.n222 7.3702
R432 VTAIL.n290 VTAIL.n224 7.3702
R433 VTAIL.n249 VTAIL.n248 7.3702
R434 VTAIL.n188 VTAIL.n116 7.3702
R435 VTAIL.n184 VTAIL.n118 7.3702
R436 VTAIL.n143 VTAIL.n142 7.3702
R437 VTAIL.n399 VTAIL.n330 6.59444
R438 VTAIL.n400 VTAIL.n399 6.59444
R439 VTAIL.n81 VTAIL.n12 6.59444
R440 VTAIL.n82 VTAIL.n81 6.59444
R441 VTAIL.n294 VTAIL.n293 6.59444
R442 VTAIL.n293 VTAIL.n224 6.59444
R443 VTAIL.n188 VTAIL.n187 6.59444
R444 VTAIL.n187 VTAIL.n118 6.59444
R445 VTAIL.n354 VTAIL.n350 5.81868
R446 VTAIL.n396 VTAIL.n395 5.81868
R447 VTAIL.n403 VTAIL.n328 5.81868
R448 VTAIL.n36 VTAIL.n32 5.81868
R449 VTAIL.n78 VTAIL.n77 5.81868
R450 VTAIL.n85 VTAIL.n10 5.81868
R451 VTAIL.n297 VTAIL.n222 5.81868
R452 VTAIL.n290 VTAIL.n289 5.81868
R453 VTAIL.n249 VTAIL.n245 5.81868
R454 VTAIL.n191 VTAIL.n116 5.81868
R455 VTAIL.n184 VTAIL.n183 5.81868
R456 VTAIL.n143 VTAIL.n139 5.81868
R457 VTAIL.n420 VTAIL.n318 5.3904
R458 VTAIL.n102 VTAIL.n0 5.3904
R459 VTAIL.n314 VTAIL.n212 5.3904
R460 VTAIL.n208 VTAIL.n106 5.3904
R461 VTAIL.n358 VTAIL.n357 5.04292
R462 VTAIL.n392 VTAIL.n332 5.04292
R463 VTAIL.n404 VTAIL.n326 5.04292
R464 VTAIL.n40 VTAIL.n39 5.04292
R465 VTAIL.n74 VTAIL.n14 5.04292
R466 VTAIL.n86 VTAIL.n8 5.04292
R467 VTAIL.n298 VTAIL.n220 5.04292
R468 VTAIL.n286 VTAIL.n226 5.04292
R469 VTAIL.n253 VTAIL.n252 5.04292
R470 VTAIL.n192 VTAIL.n114 5.04292
R471 VTAIL.n180 VTAIL.n120 5.04292
R472 VTAIL.n147 VTAIL.n146 5.04292
R473 VTAIL.n361 VTAIL.n348 4.26717
R474 VTAIL.n391 VTAIL.n334 4.26717
R475 VTAIL.n408 VTAIL.n407 4.26717
R476 VTAIL.n43 VTAIL.n30 4.26717
R477 VTAIL.n73 VTAIL.n16 4.26717
R478 VTAIL.n90 VTAIL.n89 4.26717
R479 VTAIL.n302 VTAIL.n301 4.26717
R480 VTAIL.n285 VTAIL.n228 4.26717
R481 VTAIL.n256 VTAIL.n243 4.26717
R482 VTAIL.n196 VTAIL.n195 4.26717
R483 VTAIL.n179 VTAIL.n122 4.26717
R484 VTAIL.n150 VTAIL.n137 4.26717
R485 VTAIL.n362 VTAIL.n346 3.49141
R486 VTAIL.n388 VTAIL.n387 3.49141
R487 VTAIL.n411 VTAIL.n324 3.49141
R488 VTAIL.n44 VTAIL.n28 3.49141
R489 VTAIL.n70 VTAIL.n69 3.49141
R490 VTAIL.n93 VTAIL.n6 3.49141
R491 VTAIL.n305 VTAIL.n218 3.49141
R492 VTAIL.n282 VTAIL.n281 3.49141
R493 VTAIL.n257 VTAIL.n241 3.49141
R494 VTAIL.n199 VTAIL.n112 3.49141
R495 VTAIL.n176 VTAIL.n175 3.49141
R496 VTAIL.n151 VTAIL.n135 3.49141
R497 VTAIL.n355 VTAIL.n351 2.84303
R498 VTAIL.n37 VTAIL.n33 2.84303
R499 VTAIL.n250 VTAIL.n246 2.84303
R500 VTAIL.n144 VTAIL.n140 2.84303
R501 VTAIL.n366 VTAIL.n365 2.71565
R502 VTAIL.n384 VTAIL.n336 2.71565
R503 VTAIL.n412 VTAIL.n322 2.71565
R504 VTAIL.n48 VTAIL.n47 2.71565
R505 VTAIL.n66 VTAIL.n18 2.71565
R506 VTAIL.n94 VTAIL.n4 2.71565
R507 VTAIL.n306 VTAIL.n216 2.71565
R508 VTAIL.n278 VTAIL.n230 2.71565
R509 VTAIL.n261 VTAIL.n260 2.71565
R510 VTAIL.n200 VTAIL.n110 2.71565
R511 VTAIL.n172 VTAIL.n124 2.71565
R512 VTAIL.n155 VTAIL.n154 2.71565
R513 VTAIL.n370 VTAIL.n344 1.93989
R514 VTAIL.n383 VTAIL.n338 1.93989
R515 VTAIL.n416 VTAIL.n415 1.93989
R516 VTAIL.n52 VTAIL.n26 1.93989
R517 VTAIL.n65 VTAIL.n20 1.93989
R518 VTAIL.n98 VTAIL.n97 1.93989
R519 VTAIL.n310 VTAIL.n309 1.93989
R520 VTAIL.n277 VTAIL.n232 1.93989
R521 VTAIL.n264 VTAIL.n238 1.93989
R522 VTAIL.n204 VTAIL.n203 1.93989
R523 VTAIL.n171 VTAIL.n126 1.93989
R524 VTAIL.n158 VTAIL.n132 1.93989
R525 VTAIL.n317 VTAIL.n211 1.86257
R526 VTAIL VTAIL.n105 1.22464
R527 VTAIL.n371 VTAIL.n342 1.16414
R528 VTAIL.n380 VTAIL.n379 1.16414
R529 VTAIL.n419 VTAIL.n320 1.16414
R530 VTAIL.n53 VTAIL.n24 1.16414
R531 VTAIL.n62 VTAIL.n61 1.16414
R532 VTAIL.n101 VTAIL.n2 1.16414
R533 VTAIL.n313 VTAIL.n214 1.16414
R534 VTAIL.n274 VTAIL.n273 1.16414
R535 VTAIL.n265 VTAIL.n236 1.16414
R536 VTAIL.n207 VTAIL.n108 1.16414
R537 VTAIL.n168 VTAIL.n167 1.16414
R538 VTAIL.n159 VTAIL.n130 1.16414
R539 VTAIL VTAIL.n423 0.638431
R540 VTAIL.n375 VTAIL.n374 0.388379
R541 VTAIL.n376 VTAIL.n340 0.388379
R542 VTAIL.n57 VTAIL.n56 0.388379
R543 VTAIL.n58 VTAIL.n22 0.388379
R544 VTAIL.n270 VTAIL.n234 0.388379
R545 VTAIL.n269 VTAIL.n268 0.388379
R546 VTAIL.n164 VTAIL.n128 0.388379
R547 VTAIL.n163 VTAIL.n162 0.388379
R548 VTAIL.n356 VTAIL.n355 0.155672
R549 VTAIL.n356 VTAIL.n347 0.155672
R550 VTAIL.n363 VTAIL.n347 0.155672
R551 VTAIL.n364 VTAIL.n363 0.155672
R552 VTAIL.n364 VTAIL.n343 0.155672
R553 VTAIL.n372 VTAIL.n343 0.155672
R554 VTAIL.n373 VTAIL.n372 0.155672
R555 VTAIL.n373 VTAIL.n339 0.155672
R556 VTAIL.n381 VTAIL.n339 0.155672
R557 VTAIL.n382 VTAIL.n381 0.155672
R558 VTAIL.n382 VTAIL.n335 0.155672
R559 VTAIL.n389 VTAIL.n335 0.155672
R560 VTAIL.n390 VTAIL.n389 0.155672
R561 VTAIL.n390 VTAIL.n331 0.155672
R562 VTAIL.n397 VTAIL.n331 0.155672
R563 VTAIL.n398 VTAIL.n397 0.155672
R564 VTAIL.n398 VTAIL.n327 0.155672
R565 VTAIL.n405 VTAIL.n327 0.155672
R566 VTAIL.n406 VTAIL.n405 0.155672
R567 VTAIL.n406 VTAIL.n323 0.155672
R568 VTAIL.n413 VTAIL.n323 0.155672
R569 VTAIL.n414 VTAIL.n413 0.155672
R570 VTAIL.n414 VTAIL.n319 0.155672
R571 VTAIL.n421 VTAIL.n319 0.155672
R572 VTAIL.n38 VTAIL.n37 0.155672
R573 VTAIL.n38 VTAIL.n29 0.155672
R574 VTAIL.n45 VTAIL.n29 0.155672
R575 VTAIL.n46 VTAIL.n45 0.155672
R576 VTAIL.n46 VTAIL.n25 0.155672
R577 VTAIL.n54 VTAIL.n25 0.155672
R578 VTAIL.n55 VTAIL.n54 0.155672
R579 VTAIL.n55 VTAIL.n21 0.155672
R580 VTAIL.n63 VTAIL.n21 0.155672
R581 VTAIL.n64 VTAIL.n63 0.155672
R582 VTAIL.n64 VTAIL.n17 0.155672
R583 VTAIL.n71 VTAIL.n17 0.155672
R584 VTAIL.n72 VTAIL.n71 0.155672
R585 VTAIL.n72 VTAIL.n13 0.155672
R586 VTAIL.n79 VTAIL.n13 0.155672
R587 VTAIL.n80 VTAIL.n79 0.155672
R588 VTAIL.n80 VTAIL.n9 0.155672
R589 VTAIL.n87 VTAIL.n9 0.155672
R590 VTAIL.n88 VTAIL.n87 0.155672
R591 VTAIL.n88 VTAIL.n5 0.155672
R592 VTAIL.n95 VTAIL.n5 0.155672
R593 VTAIL.n96 VTAIL.n95 0.155672
R594 VTAIL.n96 VTAIL.n1 0.155672
R595 VTAIL.n103 VTAIL.n1 0.155672
R596 VTAIL.n315 VTAIL.n213 0.155672
R597 VTAIL.n308 VTAIL.n213 0.155672
R598 VTAIL.n308 VTAIL.n307 0.155672
R599 VTAIL.n307 VTAIL.n217 0.155672
R600 VTAIL.n300 VTAIL.n217 0.155672
R601 VTAIL.n300 VTAIL.n299 0.155672
R602 VTAIL.n299 VTAIL.n221 0.155672
R603 VTAIL.n292 VTAIL.n221 0.155672
R604 VTAIL.n292 VTAIL.n291 0.155672
R605 VTAIL.n291 VTAIL.n225 0.155672
R606 VTAIL.n284 VTAIL.n225 0.155672
R607 VTAIL.n284 VTAIL.n283 0.155672
R608 VTAIL.n283 VTAIL.n229 0.155672
R609 VTAIL.n276 VTAIL.n229 0.155672
R610 VTAIL.n276 VTAIL.n275 0.155672
R611 VTAIL.n275 VTAIL.n233 0.155672
R612 VTAIL.n267 VTAIL.n233 0.155672
R613 VTAIL.n267 VTAIL.n266 0.155672
R614 VTAIL.n266 VTAIL.n237 0.155672
R615 VTAIL.n259 VTAIL.n237 0.155672
R616 VTAIL.n259 VTAIL.n258 0.155672
R617 VTAIL.n258 VTAIL.n242 0.155672
R618 VTAIL.n251 VTAIL.n242 0.155672
R619 VTAIL.n251 VTAIL.n250 0.155672
R620 VTAIL.n209 VTAIL.n107 0.155672
R621 VTAIL.n202 VTAIL.n107 0.155672
R622 VTAIL.n202 VTAIL.n201 0.155672
R623 VTAIL.n201 VTAIL.n111 0.155672
R624 VTAIL.n194 VTAIL.n111 0.155672
R625 VTAIL.n194 VTAIL.n193 0.155672
R626 VTAIL.n193 VTAIL.n115 0.155672
R627 VTAIL.n186 VTAIL.n115 0.155672
R628 VTAIL.n186 VTAIL.n185 0.155672
R629 VTAIL.n185 VTAIL.n119 0.155672
R630 VTAIL.n178 VTAIL.n119 0.155672
R631 VTAIL.n178 VTAIL.n177 0.155672
R632 VTAIL.n177 VTAIL.n123 0.155672
R633 VTAIL.n170 VTAIL.n123 0.155672
R634 VTAIL.n170 VTAIL.n169 0.155672
R635 VTAIL.n169 VTAIL.n127 0.155672
R636 VTAIL.n161 VTAIL.n127 0.155672
R637 VTAIL.n161 VTAIL.n160 0.155672
R638 VTAIL.n160 VTAIL.n131 0.155672
R639 VTAIL.n153 VTAIL.n131 0.155672
R640 VTAIL.n153 VTAIL.n152 0.155672
R641 VTAIL.n152 VTAIL.n136 0.155672
R642 VTAIL.n145 VTAIL.n136 0.155672
R643 VTAIL.n145 VTAIL.n144 0.155672
R644 VDD1.n100 VDD1.n0 214.453
R645 VDD1.n205 VDD1.n105 214.453
R646 VDD1.n101 VDD1.n100 185
R647 VDD1.n99 VDD1.n98 185
R648 VDD1.n4 VDD1.n3 185
R649 VDD1.n93 VDD1.n92 185
R650 VDD1.n91 VDD1.n90 185
R651 VDD1.n8 VDD1.n7 185
R652 VDD1.n85 VDD1.n84 185
R653 VDD1.n83 VDD1.n82 185
R654 VDD1.n12 VDD1.n11 185
R655 VDD1.n77 VDD1.n76 185
R656 VDD1.n75 VDD1.n74 185
R657 VDD1.n16 VDD1.n15 185
R658 VDD1.n69 VDD1.n68 185
R659 VDD1.n67 VDD1.n66 185
R660 VDD1.n20 VDD1.n19 185
R661 VDD1.n61 VDD1.n60 185
R662 VDD1.n59 VDD1.n58 185
R663 VDD1.n57 VDD1.n23 185
R664 VDD1.n27 VDD1.n24 185
R665 VDD1.n52 VDD1.n51 185
R666 VDD1.n50 VDD1.n49 185
R667 VDD1.n29 VDD1.n28 185
R668 VDD1.n44 VDD1.n43 185
R669 VDD1.n42 VDD1.n41 185
R670 VDD1.n33 VDD1.n32 185
R671 VDD1.n36 VDD1.n35 185
R672 VDD1.n140 VDD1.n139 185
R673 VDD1.n137 VDD1.n136 185
R674 VDD1.n146 VDD1.n145 185
R675 VDD1.n148 VDD1.n147 185
R676 VDD1.n133 VDD1.n132 185
R677 VDD1.n154 VDD1.n153 185
R678 VDD1.n157 VDD1.n156 185
R679 VDD1.n155 VDD1.n129 185
R680 VDD1.n162 VDD1.n128 185
R681 VDD1.n164 VDD1.n163 185
R682 VDD1.n166 VDD1.n165 185
R683 VDD1.n125 VDD1.n124 185
R684 VDD1.n172 VDD1.n171 185
R685 VDD1.n174 VDD1.n173 185
R686 VDD1.n121 VDD1.n120 185
R687 VDD1.n180 VDD1.n179 185
R688 VDD1.n182 VDD1.n181 185
R689 VDD1.n117 VDD1.n116 185
R690 VDD1.n188 VDD1.n187 185
R691 VDD1.n190 VDD1.n189 185
R692 VDD1.n113 VDD1.n112 185
R693 VDD1.n196 VDD1.n195 185
R694 VDD1.n198 VDD1.n197 185
R695 VDD1.n109 VDD1.n108 185
R696 VDD1.n204 VDD1.n203 185
R697 VDD1.n206 VDD1.n205 185
R698 VDD1.t1 VDD1.n34 149.524
R699 VDD1.t0 VDD1.n138 149.524
R700 VDD1.n100 VDD1.n99 104.615
R701 VDD1.n99 VDD1.n3 104.615
R702 VDD1.n92 VDD1.n3 104.615
R703 VDD1.n92 VDD1.n91 104.615
R704 VDD1.n91 VDD1.n7 104.615
R705 VDD1.n84 VDD1.n7 104.615
R706 VDD1.n84 VDD1.n83 104.615
R707 VDD1.n83 VDD1.n11 104.615
R708 VDD1.n76 VDD1.n11 104.615
R709 VDD1.n76 VDD1.n75 104.615
R710 VDD1.n75 VDD1.n15 104.615
R711 VDD1.n68 VDD1.n15 104.615
R712 VDD1.n68 VDD1.n67 104.615
R713 VDD1.n67 VDD1.n19 104.615
R714 VDD1.n60 VDD1.n19 104.615
R715 VDD1.n60 VDD1.n59 104.615
R716 VDD1.n59 VDD1.n23 104.615
R717 VDD1.n27 VDD1.n23 104.615
R718 VDD1.n51 VDD1.n27 104.615
R719 VDD1.n51 VDD1.n50 104.615
R720 VDD1.n50 VDD1.n28 104.615
R721 VDD1.n43 VDD1.n28 104.615
R722 VDD1.n43 VDD1.n42 104.615
R723 VDD1.n42 VDD1.n32 104.615
R724 VDD1.n35 VDD1.n32 104.615
R725 VDD1.n139 VDD1.n136 104.615
R726 VDD1.n146 VDD1.n136 104.615
R727 VDD1.n147 VDD1.n146 104.615
R728 VDD1.n147 VDD1.n132 104.615
R729 VDD1.n154 VDD1.n132 104.615
R730 VDD1.n156 VDD1.n154 104.615
R731 VDD1.n156 VDD1.n155 104.615
R732 VDD1.n155 VDD1.n128 104.615
R733 VDD1.n164 VDD1.n128 104.615
R734 VDD1.n165 VDD1.n164 104.615
R735 VDD1.n165 VDD1.n124 104.615
R736 VDD1.n172 VDD1.n124 104.615
R737 VDD1.n173 VDD1.n172 104.615
R738 VDD1.n173 VDD1.n120 104.615
R739 VDD1.n180 VDD1.n120 104.615
R740 VDD1.n181 VDD1.n180 104.615
R741 VDD1.n181 VDD1.n116 104.615
R742 VDD1.n188 VDD1.n116 104.615
R743 VDD1.n189 VDD1.n188 104.615
R744 VDD1.n189 VDD1.n112 104.615
R745 VDD1.n196 VDD1.n112 104.615
R746 VDD1.n197 VDD1.n196 104.615
R747 VDD1.n197 VDD1.n108 104.615
R748 VDD1.n204 VDD1.n108 104.615
R749 VDD1.n205 VDD1.n204 104.615
R750 VDD1 VDD1.n209 99.4122
R751 VDD1 VDD1.n104 52.9154
R752 VDD1.n35 VDD1.t1 52.3082
R753 VDD1.n139 VDD1.t0 52.3082
R754 VDD1.n58 VDD1.n57 13.1884
R755 VDD1.n163 VDD1.n162 13.1884
R756 VDD1.n102 VDD1.n101 12.8005
R757 VDD1.n61 VDD1.n22 12.8005
R758 VDD1.n56 VDD1.n24 12.8005
R759 VDD1.n161 VDD1.n129 12.8005
R760 VDD1.n166 VDD1.n127 12.8005
R761 VDD1.n207 VDD1.n206 12.8005
R762 VDD1.n98 VDD1.n2 12.0247
R763 VDD1.n62 VDD1.n20 12.0247
R764 VDD1.n53 VDD1.n52 12.0247
R765 VDD1.n158 VDD1.n157 12.0247
R766 VDD1.n167 VDD1.n125 12.0247
R767 VDD1.n203 VDD1.n107 12.0247
R768 VDD1.n97 VDD1.n4 11.249
R769 VDD1.n66 VDD1.n65 11.249
R770 VDD1.n49 VDD1.n26 11.249
R771 VDD1.n153 VDD1.n131 11.249
R772 VDD1.n171 VDD1.n170 11.249
R773 VDD1.n202 VDD1.n109 11.249
R774 VDD1.n94 VDD1.n93 10.4732
R775 VDD1.n69 VDD1.n18 10.4732
R776 VDD1.n48 VDD1.n29 10.4732
R777 VDD1.n152 VDD1.n133 10.4732
R778 VDD1.n174 VDD1.n123 10.4732
R779 VDD1.n199 VDD1.n198 10.4732
R780 VDD1.n36 VDD1.n34 10.2747
R781 VDD1.n140 VDD1.n138 10.2747
R782 VDD1.n90 VDD1.n6 9.69747
R783 VDD1.n70 VDD1.n16 9.69747
R784 VDD1.n45 VDD1.n44 9.69747
R785 VDD1.n149 VDD1.n148 9.69747
R786 VDD1.n175 VDD1.n121 9.69747
R787 VDD1.n195 VDD1.n111 9.69747
R788 VDD1.n104 VDD1.n103 9.45567
R789 VDD1.n209 VDD1.n208 9.45567
R790 VDD1.n38 VDD1.n37 9.3005
R791 VDD1.n40 VDD1.n39 9.3005
R792 VDD1.n31 VDD1.n30 9.3005
R793 VDD1.n46 VDD1.n45 9.3005
R794 VDD1.n48 VDD1.n47 9.3005
R795 VDD1.n26 VDD1.n25 9.3005
R796 VDD1.n54 VDD1.n53 9.3005
R797 VDD1.n56 VDD1.n55 9.3005
R798 VDD1.n10 VDD1.n9 9.3005
R799 VDD1.n87 VDD1.n86 9.3005
R800 VDD1.n89 VDD1.n88 9.3005
R801 VDD1.n6 VDD1.n5 9.3005
R802 VDD1.n95 VDD1.n94 9.3005
R803 VDD1.n97 VDD1.n96 9.3005
R804 VDD1.n2 VDD1.n1 9.3005
R805 VDD1.n103 VDD1.n102 9.3005
R806 VDD1.n81 VDD1.n80 9.3005
R807 VDD1.n79 VDD1.n78 9.3005
R808 VDD1.n14 VDD1.n13 9.3005
R809 VDD1.n73 VDD1.n72 9.3005
R810 VDD1.n71 VDD1.n70 9.3005
R811 VDD1.n18 VDD1.n17 9.3005
R812 VDD1.n65 VDD1.n64 9.3005
R813 VDD1.n63 VDD1.n62 9.3005
R814 VDD1.n22 VDD1.n21 9.3005
R815 VDD1.n184 VDD1.n183 9.3005
R816 VDD1.n119 VDD1.n118 9.3005
R817 VDD1.n178 VDD1.n177 9.3005
R818 VDD1.n176 VDD1.n175 9.3005
R819 VDD1.n123 VDD1.n122 9.3005
R820 VDD1.n170 VDD1.n169 9.3005
R821 VDD1.n168 VDD1.n167 9.3005
R822 VDD1.n127 VDD1.n126 9.3005
R823 VDD1.n142 VDD1.n141 9.3005
R824 VDD1.n144 VDD1.n143 9.3005
R825 VDD1.n135 VDD1.n134 9.3005
R826 VDD1.n150 VDD1.n149 9.3005
R827 VDD1.n152 VDD1.n151 9.3005
R828 VDD1.n131 VDD1.n130 9.3005
R829 VDD1.n159 VDD1.n158 9.3005
R830 VDD1.n161 VDD1.n160 9.3005
R831 VDD1.n186 VDD1.n185 9.3005
R832 VDD1.n115 VDD1.n114 9.3005
R833 VDD1.n192 VDD1.n191 9.3005
R834 VDD1.n194 VDD1.n193 9.3005
R835 VDD1.n111 VDD1.n110 9.3005
R836 VDD1.n200 VDD1.n199 9.3005
R837 VDD1.n202 VDD1.n201 9.3005
R838 VDD1.n107 VDD1.n106 9.3005
R839 VDD1.n208 VDD1.n207 9.3005
R840 VDD1.n89 VDD1.n8 8.92171
R841 VDD1.n74 VDD1.n73 8.92171
R842 VDD1.n41 VDD1.n31 8.92171
R843 VDD1.n145 VDD1.n135 8.92171
R844 VDD1.n179 VDD1.n178 8.92171
R845 VDD1.n194 VDD1.n113 8.92171
R846 VDD1.n104 VDD1.n0 8.2187
R847 VDD1.n209 VDD1.n105 8.2187
R848 VDD1.n86 VDD1.n85 8.14595
R849 VDD1.n77 VDD1.n14 8.14595
R850 VDD1.n40 VDD1.n33 8.14595
R851 VDD1.n144 VDD1.n137 8.14595
R852 VDD1.n182 VDD1.n119 8.14595
R853 VDD1.n191 VDD1.n190 8.14595
R854 VDD1.n82 VDD1.n10 7.3702
R855 VDD1.n78 VDD1.n12 7.3702
R856 VDD1.n37 VDD1.n36 7.3702
R857 VDD1.n141 VDD1.n140 7.3702
R858 VDD1.n183 VDD1.n117 7.3702
R859 VDD1.n187 VDD1.n115 7.3702
R860 VDD1.n82 VDD1.n81 6.59444
R861 VDD1.n81 VDD1.n12 6.59444
R862 VDD1.n186 VDD1.n117 6.59444
R863 VDD1.n187 VDD1.n186 6.59444
R864 VDD1.n85 VDD1.n10 5.81868
R865 VDD1.n78 VDD1.n77 5.81868
R866 VDD1.n37 VDD1.n33 5.81868
R867 VDD1.n141 VDD1.n137 5.81868
R868 VDD1.n183 VDD1.n182 5.81868
R869 VDD1.n190 VDD1.n115 5.81868
R870 VDD1.n102 VDD1.n0 5.3904
R871 VDD1.n207 VDD1.n105 5.3904
R872 VDD1.n86 VDD1.n8 5.04292
R873 VDD1.n74 VDD1.n14 5.04292
R874 VDD1.n41 VDD1.n40 5.04292
R875 VDD1.n145 VDD1.n144 5.04292
R876 VDD1.n179 VDD1.n119 5.04292
R877 VDD1.n191 VDD1.n113 5.04292
R878 VDD1.n90 VDD1.n89 4.26717
R879 VDD1.n73 VDD1.n16 4.26717
R880 VDD1.n44 VDD1.n31 4.26717
R881 VDD1.n148 VDD1.n135 4.26717
R882 VDD1.n178 VDD1.n121 4.26717
R883 VDD1.n195 VDD1.n194 4.26717
R884 VDD1.n93 VDD1.n6 3.49141
R885 VDD1.n70 VDD1.n69 3.49141
R886 VDD1.n45 VDD1.n29 3.49141
R887 VDD1.n149 VDD1.n133 3.49141
R888 VDD1.n175 VDD1.n174 3.49141
R889 VDD1.n198 VDD1.n111 3.49141
R890 VDD1.n142 VDD1.n138 2.84303
R891 VDD1.n38 VDD1.n34 2.84303
R892 VDD1.n94 VDD1.n4 2.71565
R893 VDD1.n66 VDD1.n18 2.71565
R894 VDD1.n49 VDD1.n48 2.71565
R895 VDD1.n153 VDD1.n152 2.71565
R896 VDD1.n171 VDD1.n123 2.71565
R897 VDD1.n199 VDD1.n109 2.71565
R898 VDD1.n98 VDD1.n97 1.93989
R899 VDD1.n65 VDD1.n20 1.93989
R900 VDD1.n52 VDD1.n26 1.93989
R901 VDD1.n157 VDD1.n131 1.93989
R902 VDD1.n170 VDD1.n125 1.93989
R903 VDD1.n203 VDD1.n202 1.93989
R904 VDD1.n101 VDD1.n2 1.16414
R905 VDD1.n62 VDD1.n61 1.16414
R906 VDD1.n53 VDD1.n24 1.16414
R907 VDD1.n158 VDD1.n129 1.16414
R908 VDD1.n167 VDD1.n166 1.16414
R909 VDD1.n206 VDD1.n107 1.16414
R910 VDD1.n58 VDD1.n22 0.388379
R911 VDD1.n57 VDD1.n56 0.388379
R912 VDD1.n162 VDD1.n161 0.388379
R913 VDD1.n163 VDD1.n127 0.388379
R914 VDD1.n103 VDD1.n1 0.155672
R915 VDD1.n96 VDD1.n1 0.155672
R916 VDD1.n96 VDD1.n95 0.155672
R917 VDD1.n95 VDD1.n5 0.155672
R918 VDD1.n88 VDD1.n5 0.155672
R919 VDD1.n88 VDD1.n87 0.155672
R920 VDD1.n87 VDD1.n9 0.155672
R921 VDD1.n80 VDD1.n9 0.155672
R922 VDD1.n80 VDD1.n79 0.155672
R923 VDD1.n79 VDD1.n13 0.155672
R924 VDD1.n72 VDD1.n13 0.155672
R925 VDD1.n72 VDD1.n71 0.155672
R926 VDD1.n71 VDD1.n17 0.155672
R927 VDD1.n64 VDD1.n17 0.155672
R928 VDD1.n64 VDD1.n63 0.155672
R929 VDD1.n63 VDD1.n21 0.155672
R930 VDD1.n55 VDD1.n21 0.155672
R931 VDD1.n55 VDD1.n54 0.155672
R932 VDD1.n54 VDD1.n25 0.155672
R933 VDD1.n47 VDD1.n25 0.155672
R934 VDD1.n47 VDD1.n46 0.155672
R935 VDD1.n46 VDD1.n30 0.155672
R936 VDD1.n39 VDD1.n30 0.155672
R937 VDD1.n39 VDD1.n38 0.155672
R938 VDD1.n143 VDD1.n142 0.155672
R939 VDD1.n143 VDD1.n134 0.155672
R940 VDD1.n150 VDD1.n134 0.155672
R941 VDD1.n151 VDD1.n150 0.155672
R942 VDD1.n151 VDD1.n130 0.155672
R943 VDD1.n159 VDD1.n130 0.155672
R944 VDD1.n160 VDD1.n159 0.155672
R945 VDD1.n160 VDD1.n126 0.155672
R946 VDD1.n168 VDD1.n126 0.155672
R947 VDD1.n169 VDD1.n168 0.155672
R948 VDD1.n169 VDD1.n122 0.155672
R949 VDD1.n176 VDD1.n122 0.155672
R950 VDD1.n177 VDD1.n176 0.155672
R951 VDD1.n177 VDD1.n118 0.155672
R952 VDD1.n184 VDD1.n118 0.155672
R953 VDD1.n185 VDD1.n184 0.155672
R954 VDD1.n185 VDD1.n114 0.155672
R955 VDD1.n192 VDD1.n114 0.155672
R956 VDD1.n193 VDD1.n192 0.155672
R957 VDD1.n193 VDD1.n110 0.155672
R958 VDD1.n200 VDD1.n110 0.155672
R959 VDD1.n201 VDD1.n200 0.155672
R960 VDD1.n201 VDD1.n106 0.155672
R961 VDD1.n208 VDD1.n106 0.155672
R962 B.n912 B.n911 585
R963 B.n913 B.n912 585
R964 B.n395 B.n121 585
R965 B.n394 B.n393 585
R966 B.n392 B.n391 585
R967 B.n390 B.n389 585
R968 B.n388 B.n387 585
R969 B.n386 B.n385 585
R970 B.n384 B.n383 585
R971 B.n382 B.n381 585
R972 B.n380 B.n379 585
R973 B.n378 B.n377 585
R974 B.n376 B.n375 585
R975 B.n374 B.n373 585
R976 B.n372 B.n371 585
R977 B.n370 B.n369 585
R978 B.n368 B.n367 585
R979 B.n366 B.n365 585
R980 B.n364 B.n363 585
R981 B.n362 B.n361 585
R982 B.n360 B.n359 585
R983 B.n358 B.n357 585
R984 B.n356 B.n355 585
R985 B.n354 B.n353 585
R986 B.n352 B.n351 585
R987 B.n350 B.n349 585
R988 B.n348 B.n347 585
R989 B.n346 B.n345 585
R990 B.n344 B.n343 585
R991 B.n342 B.n341 585
R992 B.n340 B.n339 585
R993 B.n338 B.n337 585
R994 B.n336 B.n335 585
R995 B.n334 B.n333 585
R996 B.n332 B.n331 585
R997 B.n330 B.n329 585
R998 B.n328 B.n327 585
R999 B.n326 B.n325 585
R1000 B.n324 B.n323 585
R1001 B.n322 B.n321 585
R1002 B.n320 B.n319 585
R1003 B.n318 B.n317 585
R1004 B.n316 B.n315 585
R1005 B.n314 B.n313 585
R1006 B.n312 B.n311 585
R1007 B.n310 B.n309 585
R1008 B.n308 B.n307 585
R1009 B.n306 B.n305 585
R1010 B.n304 B.n303 585
R1011 B.n302 B.n301 585
R1012 B.n300 B.n299 585
R1013 B.n298 B.n297 585
R1014 B.n296 B.n295 585
R1015 B.n294 B.n293 585
R1016 B.n292 B.n291 585
R1017 B.n290 B.n289 585
R1018 B.n288 B.n287 585
R1019 B.n286 B.n285 585
R1020 B.n284 B.n283 585
R1021 B.n282 B.n281 585
R1022 B.n280 B.n279 585
R1023 B.n278 B.n277 585
R1024 B.n276 B.n275 585
R1025 B.n274 B.n273 585
R1026 B.n272 B.n271 585
R1027 B.n269 B.n268 585
R1028 B.n267 B.n266 585
R1029 B.n265 B.n264 585
R1030 B.n263 B.n262 585
R1031 B.n261 B.n260 585
R1032 B.n259 B.n258 585
R1033 B.n257 B.n256 585
R1034 B.n255 B.n254 585
R1035 B.n253 B.n252 585
R1036 B.n251 B.n250 585
R1037 B.n249 B.n248 585
R1038 B.n247 B.n246 585
R1039 B.n245 B.n244 585
R1040 B.n243 B.n242 585
R1041 B.n241 B.n240 585
R1042 B.n239 B.n238 585
R1043 B.n237 B.n236 585
R1044 B.n235 B.n234 585
R1045 B.n233 B.n232 585
R1046 B.n231 B.n230 585
R1047 B.n229 B.n228 585
R1048 B.n227 B.n226 585
R1049 B.n225 B.n224 585
R1050 B.n223 B.n222 585
R1051 B.n221 B.n220 585
R1052 B.n219 B.n218 585
R1053 B.n217 B.n216 585
R1054 B.n215 B.n214 585
R1055 B.n213 B.n212 585
R1056 B.n211 B.n210 585
R1057 B.n209 B.n208 585
R1058 B.n207 B.n206 585
R1059 B.n205 B.n204 585
R1060 B.n203 B.n202 585
R1061 B.n201 B.n200 585
R1062 B.n199 B.n198 585
R1063 B.n197 B.n196 585
R1064 B.n195 B.n194 585
R1065 B.n193 B.n192 585
R1066 B.n191 B.n190 585
R1067 B.n189 B.n188 585
R1068 B.n187 B.n186 585
R1069 B.n185 B.n184 585
R1070 B.n183 B.n182 585
R1071 B.n181 B.n180 585
R1072 B.n179 B.n178 585
R1073 B.n177 B.n176 585
R1074 B.n175 B.n174 585
R1075 B.n173 B.n172 585
R1076 B.n171 B.n170 585
R1077 B.n169 B.n168 585
R1078 B.n167 B.n166 585
R1079 B.n165 B.n164 585
R1080 B.n163 B.n162 585
R1081 B.n161 B.n160 585
R1082 B.n159 B.n158 585
R1083 B.n157 B.n156 585
R1084 B.n155 B.n154 585
R1085 B.n153 B.n152 585
R1086 B.n151 B.n150 585
R1087 B.n149 B.n148 585
R1088 B.n147 B.n146 585
R1089 B.n145 B.n144 585
R1090 B.n143 B.n142 585
R1091 B.n141 B.n140 585
R1092 B.n139 B.n138 585
R1093 B.n137 B.n136 585
R1094 B.n135 B.n134 585
R1095 B.n133 B.n132 585
R1096 B.n131 B.n130 585
R1097 B.n129 B.n128 585
R1098 B.n53 B.n52 585
R1099 B.n916 B.n915 585
R1100 B.n910 B.n122 585
R1101 B.n122 B.n50 585
R1102 B.n909 B.n49 585
R1103 B.n920 B.n49 585
R1104 B.n908 B.n48 585
R1105 B.n921 B.n48 585
R1106 B.n907 B.n47 585
R1107 B.n922 B.n47 585
R1108 B.n906 B.n905 585
R1109 B.n905 B.n43 585
R1110 B.n904 B.n42 585
R1111 B.n928 B.n42 585
R1112 B.n903 B.n41 585
R1113 B.n929 B.n41 585
R1114 B.n902 B.n40 585
R1115 B.n930 B.n40 585
R1116 B.n901 B.n900 585
R1117 B.n900 B.n36 585
R1118 B.n899 B.n35 585
R1119 B.n936 B.n35 585
R1120 B.n898 B.n34 585
R1121 B.n937 B.n34 585
R1122 B.n897 B.n33 585
R1123 B.n938 B.n33 585
R1124 B.n896 B.n895 585
R1125 B.n895 B.n29 585
R1126 B.n894 B.n28 585
R1127 B.n944 B.n28 585
R1128 B.n893 B.n27 585
R1129 B.n945 B.n27 585
R1130 B.n892 B.n26 585
R1131 B.n946 B.n26 585
R1132 B.n891 B.n890 585
R1133 B.n890 B.n22 585
R1134 B.n889 B.n21 585
R1135 B.n952 B.n21 585
R1136 B.n888 B.n20 585
R1137 B.n953 B.n20 585
R1138 B.n887 B.n19 585
R1139 B.n954 B.n19 585
R1140 B.n886 B.n885 585
R1141 B.n885 B.n18 585
R1142 B.n884 B.n14 585
R1143 B.n960 B.n14 585
R1144 B.n883 B.n13 585
R1145 B.n961 B.n13 585
R1146 B.n882 B.n12 585
R1147 B.n962 B.n12 585
R1148 B.n881 B.n880 585
R1149 B.n880 B.n8 585
R1150 B.n879 B.n7 585
R1151 B.n968 B.n7 585
R1152 B.n878 B.n6 585
R1153 B.n969 B.n6 585
R1154 B.n877 B.n5 585
R1155 B.n970 B.n5 585
R1156 B.n876 B.n875 585
R1157 B.n875 B.n4 585
R1158 B.n874 B.n396 585
R1159 B.n874 B.n873 585
R1160 B.n864 B.n397 585
R1161 B.n398 B.n397 585
R1162 B.n866 B.n865 585
R1163 B.n867 B.n866 585
R1164 B.n863 B.n403 585
R1165 B.n403 B.n402 585
R1166 B.n862 B.n861 585
R1167 B.n861 B.n860 585
R1168 B.n405 B.n404 585
R1169 B.n853 B.n405 585
R1170 B.n852 B.n851 585
R1171 B.n854 B.n852 585
R1172 B.n850 B.n410 585
R1173 B.n410 B.n409 585
R1174 B.n849 B.n848 585
R1175 B.n848 B.n847 585
R1176 B.n412 B.n411 585
R1177 B.n413 B.n412 585
R1178 B.n840 B.n839 585
R1179 B.n841 B.n840 585
R1180 B.n838 B.n418 585
R1181 B.n418 B.n417 585
R1182 B.n837 B.n836 585
R1183 B.n836 B.n835 585
R1184 B.n420 B.n419 585
R1185 B.n421 B.n420 585
R1186 B.n828 B.n827 585
R1187 B.n829 B.n828 585
R1188 B.n826 B.n426 585
R1189 B.n426 B.n425 585
R1190 B.n825 B.n824 585
R1191 B.n824 B.n823 585
R1192 B.n428 B.n427 585
R1193 B.n429 B.n428 585
R1194 B.n816 B.n815 585
R1195 B.n817 B.n816 585
R1196 B.n814 B.n434 585
R1197 B.n434 B.n433 585
R1198 B.n813 B.n812 585
R1199 B.n812 B.n811 585
R1200 B.n436 B.n435 585
R1201 B.n437 B.n436 585
R1202 B.n804 B.n803 585
R1203 B.n805 B.n804 585
R1204 B.n802 B.n442 585
R1205 B.n442 B.n441 585
R1206 B.n801 B.n800 585
R1207 B.n800 B.n799 585
R1208 B.n444 B.n443 585
R1209 B.n445 B.n444 585
R1210 B.n795 B.n794 585
R1211 B.n448 B.n447 585
R1212 B.n791 B.n790 585
R1213 B.n792 B.n791 585
R1214 B.n789 B.n516 585
R1215 B.n788 B.n787 585
R1216 B.n786 B.n785 585
R1217 B.n784 B.n783 585
R1218 B.n782 B.n781 585
R1219 B.n780 B.n779 585
R1220 B.n778 B.n777 585
R1221 B.n776 B.n775 585
R1222 B.n774 B.n773 585
R1223 B.n772 B.n771 585
R1224 B.n770 B.n769 585
R1225 B.n768 B.n767 585
R1226 B.n766 B.n765 585
R1227 B.n764 B.n763 585
R1228 B.n762 B.n761 585
R1229 B.n760 B.n759 585
R1230 B.n758 B.n757 585
R1231 B.n756 B.n755 585
R1232 B.n754 B.n753 585
R1233 B.n752 B.n751 585
R1234 B.n750 B.n749 585
R1235 B.n748 B.n747 585
R1236 B.n746 B.n745 585
R1237 B.n744 B.n743 585
R1238 B.n742 B.n741 585
R1239 B.n740 B.n739 585
R1240 B.n738 B.n737 585
R1241 B.n736 B.n735 585
R1242 B.n734 B.n733 585
R1243 B.n732 B.n731 585
R1244 B.n730 B.n729 585
R1245 B.n728 B.n727 585
R1246 B.n726 B.n725 585
R1247 B.n724 B.n723 585
R1248 B.n722 B.n721 585
R1249 B.n720 B.n719 585
R1250 B.n718 B.n717 585
R1251 B.n716 B.n715 585
R1252 B.n714 B.n713 585
R1253 B.n712 B.n711 585
R1254 B.n710 B.n709 585
R1255 B.n708 B.n707 585
R1256 B.n706 B.n705 585
R1257 B.n704 B.n703 585
R1258 B.n702 B.n701 585
R1259 B.n700 B.n699 585
R1260 B.n698 B.n697 585
R1261 B.n696 B.n695 585
R1262 B.n694 B.n693 585
R1263 B.n692 B.n691 585
R1264 B.n690 B.n689 585
R1265 B.n688 B.n687 585
R1266 B.n686 B.n685 585
R1267 B.n684 B.n683 585
R1268 B.n682 B.n681 585
R1269 B.n680 B.n679 585
R1270 B.n678 B.n677 585
R1271 B.n676 B.n675 585
R1272 B.n674 B.n673 585
R1273 B.n672 B.n671 585
R1274 B.n670 B.n669 585
R1275 B.n667 B.n666 585
R1276 B.n665 B.n664 585
R1277 B.n663 B.n662 585
R1278 B.n661 B.n660 585
R1279 B.n659 B.n658 585
R1280 B.n657 B.n656 585
R1281 B.n655 B.n654 585
R1282 B.n653 B.n652 585
R1283 B.n651 B.n650 585
R1284 B.n649 B.n648 585
R1285 B.n647 B.n646 585
R1286 B.n645 B.n644 585
R1287 B.n643 B.n642 585
R1288 B.n641 B.n640 585
R1289 B.n639 B.n638 585
R1290 B.n637 B.n636 585
R1291 B.n635 B.n634 585
R1292 B.n633 B.n632 585
R1293 B.n631 B.n630 585
R1294 B.n629 B.n628 585
R1295 B.n627 B.n626 585
R1296 B.n625 B.n624 585
R1297 B.n623 B.n622 585
R1298 B.n621 B.n620 585
R1299 B.n619 B.n618 585
R1300 B.n617 B.n616 585
R1301 B.n615 B.n614 585
R1302 B.n613 B.n612 585
R1303 B.n611 B.n610 585
R1304 B.n609 B.n608 585
R1305 B.n607 B.n606 585
R1306 B.n605 B.n604 585
R1307 B.n603 B.n602 585
R1308 B.n601 B.n600 585
R1309 B.n599 B.n598 585
R1310 B.n597 B.n596 585
R1311 B.n595 B.n594 585
R1312 B.n593 B.n592 585
R1313 B.n591 B.n590 585
R1314 B.n589 B.n588 585
R1315 B.n587 B.n586 585
R1316 B.n585 B.n584 585
R1317 B.n583 B.n582 585
R1318 B.n581 B.n580 585
R1319 B.n579 B.n578 585
R1320 B.n577 B.n576 585
R1321 B.n575 B.n574 585
R1322 B.n573 B.n572 585
R1323 B.n571 B.n570 585
R1324 B.n569 B.n568 585
R1325 B.n567 B.n566 585
R1326 B.n565 B.n564 585
R1327 B.n563 B.n562 585
R1328 B.n561 B.n560 585
R1329 B.n559 B.n558 585
R1330 B.n557 B.n556 585
R1331 B.n555 B.n554 585
R1332 B.n553 B.n552 585
R1333 B.n551 B.n550 585
R1334 B.n549 B.n548 585
R1335 B.n547 B.n546 585
R1336 B.n545 B.n544 585
R1337 B.n543 B.n542 585
R1338 B.n541 B.n540 585
R1339 B.n539 B.n538 585
R1340 B.n537 B.n536 585
R1341 B.n535 B.n534 585
R1342 B.n533 B.n532 585
R1343 B.n531 B.n530 585
R1344 B.n529 B.n528 585
R1345 B.n527 B.n526 585
R1346 B.n525 B.n524 585
R1347 B.n523 B.n522 585
R1348 B.n796 B.n446 585
R1349 B.n446 B.n445 585
R1350 B.n798 B.n797 585
R1351 B.n799 B.n798 585
R1352 B.n440 B.n439 585
R1353 B.n441 B.n440 585
R1354 B.n807 B.n806 585
R1355 B.n806 B.n805 585
R1356 B.n808 B.n438 585
R1357 B.n438 B.n437 585
R1358 B.n810 B.n809 585
R1359 B.n811 B.n810 585
R1360 B.n432 B.n431 585
R1361 B.n433 B.n432 585
R1362 B.n819 B.n818 585
R1363 B.n818 B.n817 585
R1364 B.n820 B.n430 585
R1365 B.n430 B.n429 585
R1366 B.n822 B.n821 585
R1367 B.n823 B.n822 585
R1368 B.n424 B.n423 585
R1369 B.n425 B.n424 585
R1370 B.n831 B.n830 585
R1371 B.n830 B.n829 585
R1372 B.n832 B.n422 585
R1373 B.n422 B.n421 585
R1374 B.n834 B.n833 585
R1375 B.n835 B.n834 585
R1376 B.n416 B.n415 585
R1377 B.n417 B.n416 585
R1378 B.n843 B.n842 585
R1379 B.n842 B.n841 585
R1380 B.n844 B.n414 585
R1381 B.n414 B.n413 585
R1382 B.n846 B.n845 585
R1383 B.n847 B.n846 585
R1384 B.n408 B.n407 585
R1385 B.n409 B.n408 585
R1386 B.n856 B.n855 585
R1387 B.n855 B.n854 585
R1388 B.n857 B.n406 585
R1389 B.n853 B.n406 585
R1390 B.n859 B.n858 585
R1391 B.n860 B.n859 585
R1392 B.n401 B.n400 585
R1393 B.n402 B.n401 585
R1394 B.n869 B.n868 585
R1395 B.n868 B.n867 585
R1396 B.n870 B.n399 585
R1397 B.n399 B.n398 585
R1398 B.n872 B.n871 585
R1399 B.n873 B.n872 585
R1400 B.n2 B.n0 585
R1401 B.n4 B.n2 585
R1402 B.n3 B.n1 585
R1403 B.n969 B.n3 585
R1404 B.n967 B.n966 585
R1405 B.n968 B.n967 585
R1406 B.n965 B.n9 585
R1407 B.n9 B.n8 585
R1408 B.n964 B.n963 585
R1409 B.n963 B.n962 585
R1410 B.n11 B.n10 585
R1411 B.n961 B.n11 585
R1412 B.n959 B.n958 585
R1413 B.n960 B.n959 585
R1414 B.n957 B.n15 585
R1415 B.n18 B.n15 585
R1416 B.n956 B.n955 585
R1417 B.n955 B.n954 585
R1418 B.n17 B.n16 585
R1419 B.n953 B.n17 585
R1420 B.n951 B.n950 585
R1421 B.n952 B.n951 585
R1422 B.n949 B.n23 585
R1423 B.n23 B.n22 585
R1424 B.n948 B.n947 585
R1425 B.n947 B.n946 585
R1426 B.n25 B.n24 585
R1427 B.n945 B.n25 585
R1428 B.n943 B.n942 585
R1429 B.n944 B.n943 585
R1430 B.n941 B.n30 585
R1431 B.n30 B.n29 585
R1432 B.n940 B.n939 585
R1433 B.n939 B.n938 585
R1434 B.n32 B.n31 585
R1435 B.n937 B.n32 585
R1436 B.n935 B.n934 585
R1437 B.n936 B.n935 585
R1438 B.n933 B.n37 585
R1439 B.n37 B.n36 585
R1440 B.n932 B.n931 585
R1441 B.n931 B.n930 585
R1442 B.n39 B.n38 585
R1443 B.n929 B.n39 585
R1444 B.n927 B.n926 585
R1445 B.n928 B.n927 585
R1446 B.n925 B.n44 585
R1447 B.n44 B.n43 585
R1448 B.n924 B.n923 585
R1449 B.n923 B.n922 585
R1450 B.n46 B.n45 585
R1451 B.n921 B.n46 585
R1452 B.n919 B.n918 585
R1453 B.n920 B.n919 585
R1454 B.n917 B.n51 585
R1455 B.n51 B.n50 585
R1456 B.n972 B.n971 585
R1457 B.n971 B.n970 585
R1458 B.n794 B.n446 506.916
R1459 B.n915 B.n51 506.916
R1460 B.n522 B.n444 506.916
R1461 B.n912 B.n122 506.916
R1462 B.n519 B.t15 473.68
R1463 B.n123 B.t11 473.68
R1464 B.n517 B.t9 473.68
R1465 B.n125 B.t4 473.68
R1466 B.n520 B.t14 411.038
R1467 B.n124 B.t12 411.038
R1468 B.n518 B.t8 411.038
R1469 B.n126 B.t5 411.038
R1470 B.n519 B.t13 370.428
R1471 B.n517 B.t6 370.428
R1472 B.n125 B.t2 370.428
R1473 B.n123 B.t10 370.428
R1474 B.n913 B.n120 256.663
R1475 B.n913 B.n119 256.663
R1476 B.n913 B.n118 256.663
R1477 B.n913 B.n117 256.663
R1478 B.n913 B.n116 256.663
R1479 B.n913 B.n115 256.663
R1480 B.n913 B.n114 256.663
R1481 B.n913 B.n113 256.663
R1482 B.n913 B.n112 256.663
R1483 B.n913 B.n111 256.663
R1484 B.n913 B.n110 256.663
R1485 B.n913 B.n109 256.663
R1486 B.n913 B.n108 256.663
R1487 B.n913 B.n107 256.663
R1488 B.n913 B.n106 256.663
R1489 B.n913 B.n105 256.663
R1490 B.n913 B.n104 256.663
R1491 B.n913 B.n103 256.663
R1492 B.n913 B.n102 256.663
R1493 B.n913 B.n101 256.663
R1494 B.n913 B.n100 256.663
R1495 B.n913 B.n99 256.663
R1496 B.n913 B.n98 256.663
R1497 B.n913 B.n97 256.663
R1498 B.n913 B.n96 256.663
R1499 B.n913 B.n95 256.663
R1500 B.n913 B.n94 256.663
R1501 B.n913 B.n93 256.663
R1502 B.n913 B.n92 256.663
R1503 B.n913 B.n91 256.663
R1504 B.n913 B.n90 256.663
R1505 B.n913 B.n89 256.663
R1506 B.n913 B.n88 256.663
R1507 B.n913 B.n87 256.663
R1508 B.n913 B.n86 256.663
R1509 B.n913 B.n85 256.663
R1510 B.n913 B.n84 256.663
R1511 B.n913 B.n83 256.663
R1512 B.n913 B.n82 256.663
R1513 B.n913 B.n81 256.663
R1514 B.n913 B.n80 256.663
R1515 B.n913 B.n79 256.663
R1516 B.n913 B.n78 256.663
R1517 B.n913 B.n77 256.663
R1518 B.n913 B.n76 256.663
R1519 B.n913 B.n75 256.663
R1520 B.n913 B.n74 256.663
R1521 B.n913 B.n73 256.663
R1522 B.n913 B.n72 256.663
R1523 B.n913 B.n71 256.663
R1524 B.n913 B.n70 256.663
R1525 B.n913 B.n69 256.663
R1526 B.n913 B.n68 256.663
R1527 B.n913 B.n67 256.663
R1528 B.n913 B.n66 256.663
R1529 B.n913 B.n65 256.663
R1530 B.n913 B.n64 256.663
R1531 B.n913 B.n63 256.663
R1532 B.n913 B.n62 256.663
R1533 B.n913 B.n61 256.663
R1534 B.n913 B.n60 256.663
R1535 B.n913 B.n59 256.663
R1536 B.n913 B.n58 256.663
R1537 B.n913 B.n57 256.663
R1538 B.n913 B.n56 256.663
R1539 B.n913 B.n55 256.663
R1540 B.n913 B.n54 256.663
R1541 B.n914 B.n913 256.663
R1542 B.n793 B.n792 256.663
R1543 B.n792 B.n449 256.663
R1544 B.n792 B.n450 256.663
R1545 B.n792 B.n451 256.663
R1546 B.n792 B.n452 256.663
R1547 B.n792 B.n453 256.663
R1548 B.n792 B.n454 256.663
R1549 B.n792 B.n455 256.663
R1550 B.n792 B.n456 256.663
R1551 B.n792 B.n457 256.663
R1552 B.n792 B.n458 256.663
R1553 B.n792 B.n459 256.663
R1554 B.n792 B.n460 256.663
R1555 B.n792 B.n461 256.663
R1556 B.n792 B.n462 256.663
R1557 B.n792 B.n463 256.663
R1558 B.n792 B.n464 256.663
R1559 B.n792 B.n465 256.663
R1560 B.n792 B.n466 256.663
R1561 B.n792 B.n467 256.663
R1562 B.n792 B.n468 256.663
R1563 B.n792 B.n469 256.663
R1564 B.n792 B.n470 256.663
R1565 B.n792 B.n471 256.663
R1566 B.n792 B.n472 256.663
R1567 B.n792 B.n473 256.663
R1568 B.n792 B.n474 256.663
R1569 B.n792 B.n475 256.663
R1570 B.n792 B.n476 256.663
R1571 B.n792 B.n477 256.663
R1572 B.n792 B.n478 256.663
R1573 B.n792 B.n479 256.663
R1574 B.n792 B.n480 256.663
R1575 B.n792 B.n481 256.663
R1576 B.n792 B.n482 256.663
R1577 B.n792 B.n483 256.663
R1578 B.n792 B.n484 256.663
R1579 B.n792 B.n485 256.663
R1580 B.n792 B.n486 256.663
R1581 B.n792 B.n487 256.663
R1582 B.n792 B.n488 256.663
R1583 B.n792 B.n489 256.663
R1584 B.n792 B.n490 256.663
R1585 B.n792 B.n491 256.663
R1586 B.n792 B.n492 256.663
R1587 B.n792 B.n493 256.663
R1588 B.n792 B.n494 256.663
R1589 B.n792 B.n495 256.663
R1590 B.n792 B.n496 256.663
R1591 B.n792 B.n497 256.663
R1592 B.n792 B.n498 256.663
R1593 B.n792 B.n499 256.663
R1594 B.n792 B.n500 256.663
R1595 B.n792 B.n501 256.663
R1596 B.n792 B.n502 256.663
R1597 B.n792 B.n503 256.663
R1598 B.n792 B.n504 256.663
R1599 B.n792 B.n505 256.663
R1600 B.n792 B.n506 256.663
R1601 B.n792 B.n507 256.663
R1602 B.n792 B.n508 256.663
R1603 B.n792 B.n509 256.663
R1604 B.n792 B.n510 256.663
R1605 B.n792 B.n511 256.663
R1606 B.n792 B.n512 256.663
R1607 B.n792 B.n513 256.663
R1608 B.n792 B.n514 256.663
R1609 B.n792 B.n515 256.663
R1610 B.n798 B.n446 163.367
R1611 B.n798 B.n440 163.367
R1612 B.n806 B.n440 163.367
R1613 B.n806 B.n438 163.367
R1614 B.n810 B.n438 163.367
R1615 B.n810 B.n432 163.367
R1616 B.n818 B.n432 163.367
R1617 B.n818 B.n430 163.367
R1618 B.n822 B.n430 163.367
R1619 B.n822 B.n424 163.367
R1620 B.n830 B.n424 163.367
R1621 B.n830 B.n422 163.367
R1622 B.n834 B.n422 163.367
R1623 B.n834 B.n416 163.367
R1624 B.n842 B.n416 163.367
R1625 B.n842 B.n414 163.367
R1626 B.n846 B.n414 163.367
R1627 B.n846 B.n408 163.367
R1628 B.n855 B.n408 163.367
R1629 B.n855 B.n406 163.367
R1630 B.n859 B.n406 163.367
R1631 B.n859 B.n401 163.367
R1632 B.n868 B.n401 163.367
R1633 B.n868 B.n399 163.367
R1634 B.n872 B.n399 163.367
R1635 B.n872 B.n2 163.367
R1636 B.n971 B.n2 163.367
R1637 B.n971 B.n3 163.367
R1638 B.n967 B.n3 163.367
R1639 B.n967 B.n9 163.367
R1640 B.n963 B.n9 163.367
R1641 B.n963 B.n11 163.367
R1642 B.n959 B.n11 163.367
R1643 B.n959 B.n15 163.367
R1644 B.n955 B.n15 163.367
R1645 B.n955 B.n17 163.367
R1646 B.n951 B.n17 163.367
R1647 B.n951 B.n23 163.367
R1648 B.n947 B.n23 163.367
R1649 B.n947 B.n25 163.367
R1650 B.n943 B.n25 163.367
R1651 B.n943 B.n30 163.367
R1652 B.n939 B.n30 163.367
R1653 B.n939 B.n32 163.367
R1654 B.n935 B.n32 163.367
R1655 B.n935 B.n37 163.367
R1656 B.n931 B.n37 163.367
R1657 B.n931 B.n39 163.367
R1658 B.n927 B.n39 163.367
R1659 B.n927 B.n44 163.367
R1660 B.n923 B.n44 163.367
R1661 B.n923 B.n46 163.367
R1662 B.n919 B.n46 163.367
R1663 B.n919 B.n51 163.367
R1664 B.n791 B.n448 163.367
R1665 B.n791 B.n516 163.367
R1666 B.n787 B.n786 163.367
R1667 B.n783 B.n782 163.367
R1668 B.n779 B.n778 163.367
R1669 B.n775 B.n774 163.367
R1670 B.n771 B.n770 163.367
R1671 B.n767 B.n766 163.367
R1672 B.n763 B.n762 163.367
R1673 B.n759 B.n758 163.367
R1674 B.n755 B.n754 163.367
R1675 B.n751 B.n750 163.367
R1676 B.n747 B.n746 163.367
R1677 B.n743 B.n742 163.367
R1678 B.n739 B.n738 163.367
R1679 B.n735 B.n734 163.367
R1680 B.n731 B.n730 163.367
R1681 B.n727 B.n726 163.367
R1682 B.n723 B.n722 163.367
R1683 B.n719 B.n718 163.367
R1684 B.n715 B.n714 163.367
R1685 B.n711 B.n710 163.367
R1686 B.n707 B.n706 163.367
R1687 B.n703 B.n702 163.367
R1688 B.n699 B.n698 163.367
R1689 B.n695 B.n694 163.367
R1690 B.n691 B.n690 163.367
R1691 B.n687 B.n686 163.367
R1692 B.n683 B.n682 163.367
R1693 B.n679 B.n678 163.367
R1694 B.n675 B.n674 163.367
R1695 B.n671 B.n670 163.367
R1696 B.n666 B.n665 163.367
R1697 B.n662 B.n661 163.367
R1698 B.n658 B.n657 163.367
R1699 B.n654 B.n653 163.367
R1700 B.n650 B.n649 163.367
R1701 B.n646 B.n645 163.367
R1702 B.n642 B.n641 163.367
R1703 B.n638 B.n637 163.367
R1704 B.n634 B.n633 163.367
R1705 B.n630 B.n629 163.367
R1706 B.n626 B.n625 163.367
R1707 B.n622 B.n621 163.367
R1708 B.n618 B.n617 163.367
R1709 B.n614 B.n613 163.367
R1710 B.n610 B.n609 163.367
R1711 B.n606 B.n605 163.367
R1712 B.n602 B.n601 163.367
R1713 B.n598 B.n597 163.367
R1714 B.n594 B.n593 163.367
R1715 B.n590 B.n589 163.367
R1716 B.n586 B.n585 163.367
R1717 B.n582 B.n581 163.367
R1718 B.n578 B.n577 163.367
R1719 B.n574 B.n573 163.367
R1720 B.n570 B.n569 163.367
R1721 B.n566 B.n565 163.367
R1722 B.n562 B.n561 163.367
R1723 B.n558 B.n557 163.367
R1724 B.n554 B.n553 163.367
R1725 B.n550 B.n549 163.367
R1726 B.n546 B.n545 163.367
R1727 B.n542 B.n541 163.367
R1728 B.n538 B.n537 163.367
R1729 B.n534 B.n533 163.367
R1730 B.n530 B.n529 163.367
R1731 B.n526 B.n525 163.367
R1732 B.n800 B.n444 163.367
R1733 B.n800 B.n442 163.367
R1734 B.n804 B.n442 163.367
R1735 B.n804 B.n436 163.367
R1736 B.n812 B.n436 163.367
R1737 B.n812 B.n434 163.367
R1738 B.n816 B.n434 163.367
R1739 B.n816 B.n428 163.367
R1740 B.n824 B.n428 163.367
R1741 B.n824 B.n426 163.367
R1742 B.n828 B.n426 163.367
R1743 B.n828 B.n420 163.367
R1744 B.n836 B.n420 163.367
R1745 B.n836 B.n418 163.367
R1746 B.n840 B.n418 163.367
R1747 B.n840 B.n412 163.367
R1748 B.n848 B.n412 163.367
R1749 B.n848 B.n410 163.367
R1750 B.n852 B.n410 163.367
R1751 B.n852 B.n405 163.367
R1752 B.n861 B.n405 163.367
R1753 B.n861 B.n403 163.367
R1754 B.n866 B.n403 163.367
R1755 B.n866 B.n397 163.367
R1756 B.n874 B.n397 163.367
R1757 B.n875 B.n874 163.367
R1758 B.n875 B.n5 163.367
R1759 B.n6 B.n5 163.367
R1760 B.n7 B.n6 163.367
R1761 B.n880 B.n7 163.367
R1762 B.n880 B.n12 163.367
R1763 B.n13 B.n12 163.367
R1764 B.n14 B.n13 163.367
R1765 B.n885 B.n14 163.367
R1766 B.n885 B.n19 163.367
R1767 B.n20 B.n19 163.367
R1768 B.n21 B.n20 163.367
R1769 B.n890 B.n21 163.367
R1770 B.n890 B.n26 163.367
R1771 B.n27 B.n26 163.367
R1772 B.n28 B.n27 163.367
R1773 B.n895 B.n28 163.367
R1774 B.n895 B.n33 163.367
R1775 B.n34 B.n33 163.367
R1776 B.n35 B.n34 163.367
R1777 B.n900 B.n35 163.367
R1778 B.n900 B.n40 163.367
R1779 B.n41 B.n40 163.367
R1780 B.n42 B.n41 163.367
R1781 B.n905 B.n42 163.367
R1782 B.n905 B.n47 163.367
R1783 B.n48 B.n47 163.367
R1784 B.n49 B.n48 163.367
R1785 B.n122 B.n49 163.367
R1786 B.n128 B.n53 163.367
R1787 B.n132 B.n131 163.367
R1788 B.n136 B.n135 163.367
R1789 B.n140 B.n139 163.367
R1790 B.n144 B.n143 163.367
R1791 B.n148 B.n147 163.367
R1792 B.n152 B.n151 163.367
R1793 B.n156 B.n155 163.367
R1794 B.n160 B.n159 163.367
R1795 B.n164 B.n163 163.367
R1796 B.n168 B.n167 163.367
R1797 B.n172 B.n171 163.367
R1798 B.n176 B.n175 163.367
R1799 B.n180 B.n179 163.367
R1800 B.n184 B.n183 163.367
R1801 B.n188 B.n187 163.367
R1802 B.n192 B.n191 163.367
R1803 B.n196 B.n195 163.367
R1804 B.n200 B.n199 163.367
R1805 B.n204 B.n203 163.367
R1806 B.n208 B.n207 163.367
R1807 B.n212 B.n211 163.367
R1808 B.n216 B.n215 163.367
R1809 B.n220 B.n219 163.367
R1810 B.n224 B.n223 163.367
R1811 B.n228 B.n227 163.367
R1812 B.n232 B.n231 163.367
R1813 B.n236 B.n235 163.367
R1814 B.n240 B.n239 163.367
R1815 B.n244 B.n243 163.367
R1816 B.n248 B.n247 163.367
R1817 B.n252 B.n251 163.367
R1818 B.n256 B.n255 163.367
R1819 B.n260 B.n259 163.367
R1820 B.n264 B.n263 163.367
R1821 B.n268 B.n267 163.367
R1822 B.n273 B.n272 163.367
R1823 B.n277 B.n276 163.367
R1824 B.n281 B.n280 163.367
R1825 B.n285 B.n284 163.367
R1826 B.n289 B.n288 163.367
R1827 B.n293 B.n292 163.367
R1828 B.n297 B.n296 163.367
R1829 B.n301 B.n300 163.367
R1830 B.n305 B.n304 163.367
R1831 B.n309 B.n308 163.367
R1832 B.n313 B.n312 163.367
R1833 B.n317 B.n316 163.367
R1834 B.n321 B.n320 163.367
R1835 B.n325 B.n324 163.367
R1836 B.n329 B.n328 163.367
R1837 B.n333 B.n332 163.367
R1838 B.n337 B.n336 163.367
R1839 B.n341 B.n340 163.367
R1840 B.n345 B.n344 163.367
R1841 B.n349 B.n348 163.367
R1842 B.n353 B.n352 163.367
R1843 B.n357 B.n356 163.367
R1844 B.n361 B.n360 163.367
R1845 B.n365 B.n364 163.367
R1846 B.n369 B.n368 163.367
R1847 B.n373 B.n372 163.367
R1848 B.n377 B.n376 163.367
R1849 B.n381 B.n380 163.367
R1850 B.n385 B.n384 163.367
R1851 B.n389 B.n388 163.367
R1852 B.n393 B.n392 163.367
R1853 B.n912 B.n121 163.367
R1854 B.n794 B.n793 71.676
R1855 B.n516 B.n449 71.676
R1856 B.n786 B.n450 71.676
R1857 B.n782 B.n451 71.676
R1858 B.n778 B.n452 71.676
R1859 B.n774 B.n453 71.676
R1860 B.n770 B.n454 71.676
R1861 B.n766 B.n455 71.676
R1862 B.n762 B.n456 71.676
R1863 B.n758 B.n457 71.676
R1864 B.n754 B.n458 71.676
R1865 B.n750 B.n459 71.676
R1866 B.n746 B.n460 71.676
R1867 B.n742 B.n461 71.676
R1868 B.n738 B.n462 71.676
R1869 B.n734 B.n463 71.676
R1870 B.n730 B.n464 71.676
R1871 B.n726 B.n465 71.676
R1872 B.n722 B.n466 71.676
R1873 B.n718 B.n467 71.676
R1874 B.n714 B.n468 71.676
R1875 B.n710 B.n469 71.676
R1876 B.n706 B.n470 71.676
R1877 B.n702 B.n471 71.676
R1878 B.n698 B.n472 71.676
R1879 B.n694 B.n473 71.676
R1880 B.n690 B.n474 71.676
R1881 B.n686 B.n475 71.676
R1882 B.n682 B.n476 71.676
R1883 B.n678 B.n477 71.676
R1884 B.n674 B.n478 71.676
R1885 B.n670 B.n479 71.676
R1886 B.n665 B.n480 71.676
R1887 B.n661 B.n481 71.676
R1888 B.n657 B.n482 71.676
R1889 B.n653 B.n483 71.676
R1890 B.n649 B.n484 71.676
R1891 B.n645 B.n485 71.676
R1892 B.n641 B.n486 71.676
R1893 B.n637 B.n487 71.676
R1894 B.n633 B.n488 71.676
R1895 B.n629 B.n489 71.676
R1896 B.n625 B.n490 71.676
R1897 B.n621 B.n491 71.676
R1898 B.n617 B.n492 71.676
R1899 B.n613 B.n493 71.676
R1900 B.n609 B.n494 71.676
R1901 B.n605 B.n495 71.676
R1902 B.n601 B.n496 71.676
R1903 B.n597 B.n497 71.676
R1904 B.n593 B.n498 71.676
R1905 B.n589 B.n499 71.676
R1906 B.n585 B.n500 71.676
R1907 B.n581 B.n501 71.676
R1908 B.n577 B.n502 71.676
R1909 B.n573 B.n503 71.676
R1910 B.n569 B.n504 71.676
R1911 B.n565 B.n505 71.676
R1912 B.n561 B.n506 71.676
R1913 B.n557 B.n507 71.676
R1914 B.n553 B.n508 71.676
R1915 B.n549 B.n509 71.676
R1916 B.n545 B.n510 71.676
R1917 B.n541 B.n511 71.676
R1918 B.n537 B.n512 71.676
R1919 B.n533 B.n513 71.676
R1920 B.n529 B.n514 71.676
R1921 B.n525 B.n515 71.676
R1922 B.n915 B.n914 71.676
R1923 B.n128 B.n54 71.676
R1924 B.n132 B.n55 71.676
R1925 B.n136 B.n56 71.676
R1926 B.n140 B.n57 71.676
R1927 B.n144 B.n58 71.676
R1928 B.n148 B.n59 71.676
R1929 B.n152 B.n60 71.676
R1930 B.n156 B.n61 71.676
R1931 B.n160 B.n62 71.676
R1932 B.n164 B.n63 71.676
R1933 B.n168 B.n64 71.676
R1934 B.n172 B.n65 71.676
R1935 B.n176 B.n66 71.676
R1936 B.n180 B.n67 71.676
R1937 B.n184 B.n68 71.676
R1938 B.n188 B.n69 71.676
R1939 B.n192 B.n70 71.676
R1940 B.n196 B.n71 71.676
R1941 B.n200 B.n72 71.676
R1942 B.n204 B.n73 71.676
R1943 B.n208 B.n74 71.676
R1944 B.n212 B.n75 71.676
R1945 B.n216 B.n76 71.676
R1946 B.n220 B.n77 71.676
R1947 B.n224 B.n78 71.676
R1948 B.n228 B.n79 71.676
R1949 B.n232 B.n80 71.676
R1950 B.n236 B.n81 71.676
R1951 B.n240 B.n82 71.676
R1952 B.n244 B.n83 71.676
R1953 B.n248 B.n84 71.676
R1954 B.n252 B.n85 71.676
R1955 B.n256 B.n86 71.676
R1956 B.n260 B.n87 71.676
R1957 B.n264 B.n88 71.676
R1958 B.n268 B.n89 71.676
R1959 B.n273 B.n90 71.676
R1960 B.n277 B.n91 71.676
R1961 B.n281 B.n92 71.676
R1962 B.n285 B.n93 71.676
R1963 B.n289 B.n94 71.676
R1964 B.n293 B.n95 71.676
R1965 B.n297 B.n96 71.676
R1966 B.n301 B.n97 71.676
R1967 B.n305 B.n98 71.676
R1968 B.n309 B.n99 71.676
R1969 B.n313 B.n100 71.676
R1970 B.n317 B.n101 71.676
R1971 B.n321 B.n102 71.676
R1972 B.n325 B.n103 71.676
R1973 B.n329 B.n104 71.676
R1974 B.n333 B.n105 71.676
R1975 B.n337 B.n106 71.676
R1976 B.n341 B.n107 71.676
R1977 B.n345 B.n108 71.676
R1978 B.n349 B.n109 71.676
R1979 B.n353 B.n110 71.676
R1980 B.n357 B.n111 71.676
R1981 B.n361 B.n112 71.676
R1982 B.n365 B.n113 71.676
R1983 B.n369 B.n114 71.676
R1984 B.n373 B.n115 71.676
R1985 B.n377 B.n116 71.676
R1986 B.n381 B.n117 71.676
R1987 B.n385 B.n118 71.676
R1988 B.n389 B.n119 71.676
R1989 B.n393 B.n120 71.676
R1990 B.n121 B.n120 71.676
R1991 B.n392 B.n119 71.676
R1992 B.n388 B.n118 71.676
R1993 B.n384 B.n117 71.676
R1994 B.n380 B.n116 71.676
R1995 B.n376 B.n115 71.676
R1996 B.n372 B.n114 71.676
R1997 B.n368 B.n113 71.676
R1998 B.n364 B.n112 71.676
R1999 B.n360 B.n111 71.676
R2000 B.n356 B.n110 71.676
R2001 B.n352 B.n109 71.676
R2002 B.n348 B.n108 71.676
R2003 B.n344 B.n107 71.676
R2004 B.n340 B.n106 71.676
R2005 B.n336 B.n105 71.676
R2006 B.n332 B.n104 71.676
R2007 B.n328 B.n103 71.676
R2008 B.n324 B.n102 71.676
R2009 B.n320 B.n101 71.676
R2010 B.n316 B.n100 71.676
R2011 B.n312 B.n99 71.676
R2012 B.n308 B.n98 71.676
R2013 B.n304 B.n97 71.676
R2014 B.n300 B.n96 71.676
R2015 B.n296 B.n95 71.676
R2016 B.n292 B.n94 71.676
R2017 B.n288 B.n93 71.676
R2018 B.n284 B.n92 71.676
R2019 B.n280 B.n91 71.676
R2020 B.n276 B.n90 71.676
R2021 B.n272 B.n89 71.676
R2022 B.n267 B.n88 71.676
R2023 B.n263 B.n87 71.676
R2024 B.n259 B.n86 71.676
R2025 B.n255 B.n85 71.676
R2026 B.n251 B.n84 71.676
R2027 B.n247 B.n83 71.676
R2028 B.n243 B.n82 71.676
R2029 B.n239 B.n81 71.676
R2030 B.n235 B.n80 71.676
R2031 B.n231 B.n79 71.676
R2032 B.n227 B.n78 71.676
R2033 B.n223 B.n77 71.676
R2034 B.n219 B.n76 71.676
R2035 B.n215 B.n75 71.676
R2036 B.n211 B.n74 71.676
R2037 B.n207 B.n73 71.676
R2038 B.n203 B.n72 71.676
R2039 B.n199 B.n71 71.676
R2040 B.n195 B.n70 71.676
R2041 B.n191 B.n69 71.676
R2042 B.n187 B.n68 71.676
R2043 B.n183 B.n67 71.676
R2044 B.n179 B.n66 71.676
R2045 B.n175 B.n65 71.676
R2046 B.n171 B.n64 71.676
R2047 B.n167 B.n63 71.676
R2048 B.n163 B.n62 71.676
R2049 B.n159 B.n61 71.676
R2050 B.n155 B.n60 71.676
R2051 B.n151 B.n59 71.676
R2052 B.n147 B.n58 71.676
R2053 B.n143 B.n57 71.676
R2054 B.n139 B.n56 71.676
R2055 B.n135 B.n55 71.676
R2056 B.n131 B.n54 71.676
R2057 B.n914 B.n53 71.676
R2058 B.n793 B.n448 71.676
R2059 B.n787 B.n449 71.676
R2060 B.n783 B.n450 71.676
R2061 B.n779 B.n451 71.676
R2062 B.n775 B.n452 71.676
R2063 B.n771 B.n453 71.676
R2064 B.n767 B.n454 71.676
R2065 B.n763 B.n455 71.676
R2066 B.n759 B.n456 71.676
R2067 B.n755 B.n457 71.676
R2068 B.n751 B.n458 71.676
R2069 B.n747 B.n459 71.676
R2070 B.n743 B.n460 71.676
R2071 B.n739 B.n461 71.676
R2072 B.n735 B.n462 71.676
R2073 B.n731 B.n463 71.676
R2074 B.n727 B.n464 71.676
R2075 B.n723 B.n465 71.676
R2076 B.n719 B.n466 71.676
R2077 B.n715 B.n467 71.676
R2078 B.n711 B.n468 71.676
R2079 B.n707 B.n469 71.676
R2080 B.n703 B.n470 71.676
R2081 B.n699 B.n471 71.676
R2082 B.n695 B.n472 71.676
R2083 B.n691 B.n473 71.676
R2084 B.n687 B.n474 71.676
R2085 B.n683 B.n475 71.676
R2086 B.n679 B.n476 71.676
R2087 B.n675 B.n477 71.676
R2088 B.n671 B.n478 71.676
R2089 B.n666 B.n479 71.676
R2090 B.n662 B.n480 71.676
R2091 B.n658 B.n481 71.676
R2092 B.n654 B.n482 71.676
R2093 B.n650 B.n483 71.676
R2094 B.n646 B.n484 71.676
R2095 B.n642 B.n485 71.676
R2096 B.n638 B.n486 71.676
R2097 B.n634 B.n487 71.676
R2098 B.n630 B.n488 71.676
R2099 B.n626 B.n489 71.676
R2100 B.n622 B.n490 71.676
R2101 B.n618 B.n491 71.676
R2102 B.n614 B.n492 71.676
R2103 B.n610 B.n493 71.676
R2104 B.n606 B.n494 71.676
R2105 B.n602 B.n495 71.676
R2106 B.n598 B.n496 71.676
R2107 B.n594 B.n497 71.676
R2108 B.n590 B.n498 71.676
R2109 B.n586 B.n499 71.676
R2110 B.n582 B.n500 71.676
R2111 B.n578 B.n501 71.676
R2112 B.n574 B.n502 71.676
R2113 B.n570 B.n503 71.676
R2114 B.n566 B.n504 71.676
R2115 B.n562 B.n505 71.676
R2116 B.n558 B.n506 71.676
R2117 B.n554 B.n507 71.676
R2118 B.n550 B.n508 71.676
R2119 B.n546 B.n509 71.676
R2120 B.n542 B.n510 71.676
R2121 B.n538 B.n511 71.676
R2122 B.n534 B.n512 71.676
R2123 B.n530 B.n513 71.676
R2124 B.n526 B.n514 71.676
R2125 B.n522 B.n515 71.676
R2126 B.n520 B.n519 62.6429
R2127 B.n518 B.n517 62.6429
R2128 B.n126 B.n125 62.6429
R2129 B.n124 B.n123 62.6429
R2130 B.n521 B.n520 59.5399
R2131 B.n668 B.n518 59.5399
R2132 B.n127 B.n126 59.5399
R2133 B.n270 B.n124 59.5399
R2134 B.n792 B.n445 58.1875
R2135 B.n913 B.n50 58.1875
R2136 B.n917 B.n916 32.9371
R2137 B.n911 B.n910 32.9371
R2138 B.n523 B.n443 32.9371
R2139 B.n796 B.n795 32.9371
R2140 B.n799 B.n445 30.2044
R2141 B.n799 B.n441 30.2044
R2142 B.n805 B.n441 30.2044
R2143 B.n805 B.n437 30.2044
R2144 B.n811 B.n437 30.2044
R2145 B.n811 B.n433 30.2044
R2146 B.n817 B.n433 30.2044
R2147 B.n823 B.n429 30.2044
R2148 B.n823 B.n425 30.2044
R2149 B.n829 B.n425 30.2044
R2150 B.n829 B.n421 30.2044
R2151 B.n835 B.n421 30.2044
R2152 B.n835 B.n417 30.2044
R2153 B.n841 B.n417 30.2044
R2154 B.n841 B.n413 30.2044
R2155 B.n847 B.n413 30.2044
R2156 B.n847 B.n409 30.2044
R2157 B.n854 B.n409 30.2044
R2158 B.n854 B.n853 30.2044
R2159 B.n860 B.n402 30.2044
R2160 B.n867 B.n402 30.2044
R2161 B.n867 B.n398 30.2044
R2162 B.n873 B.n398 30.2044
R2163 B.n873 B.n4 30.2044
R2164 B.n970 B.n4 30.2044
R2165 B.n970 B.n969 30.2044
R2166 B.n969 B.n968 30.2044
R2167 B.n968 B.n8 30.2044
R2168 B.n962 B.n8 30.2044
R2169 B.n962 B.n961 30.2044
R2170 B.n961 B.n960 30.2044
R2171 B.n954 B.n18 30.2044
R2172 B.n954 B.n953 30.2044
R2173 B.n953 B.n952 30.2044
R2174 B.n952 B.n22 30.2044
R2175 B.n946 B.n22 30.2044
R2176 B.n946 B.n945 30.2044
R2177 B.n945 B.n944 30.2044
R2178 B.n944 B.n29 30.2044
R2179 B.n938 B.n29 30.2044
R2180 B.n938 B.n937 30.2044
R2181 B.n937 B.n936 30.2044
R2182 B.n936 B.n36 30.2044
R2183 B.n930 B.n929 30.2044
R2184 B.n929 B.n928 30.2044
R2185 B.n928 B.n43 30.2044
R2186 B.n922 B.n43 30.2044
R2187 B.n922 B.n921 30.2044
R2188 B.n921 B.n920 30.2044
R2189 B.n920 B.n50 30.2044
R2190 B.n817 B.t7 28.4277
R2191 B.n930 B.t3 28.4277
R2192 B.n853 B.t1 19.5442
R2193 B.n18 B.t0 19.5442
R2194 B B.n972 18.0485
R2195 B.n860 B.t1 10.6607
R2196 B.n960 B.t0 10.6607
R2197 B.n916 B.n52 10.6151
R2198 B.n129 B.n52 10.6151
R2199 B.n130 B.n129 10.6151
R2200 B.n133 B.n130 10.6151
R2201 B.n134 B.n133 10.6151
R2202 B.n137 B.n134 10.6151
R2203 B.n138 B.n137 10.6151
R2204 B.n141 B.n138 10.6151
R2205 B.n142 B.n141 10.6151
R2206 B.n145 B.n142 10.6151
R2207 B.n146 B.n145 10.6151
R2208 B.n149 B.n146 10.6151
R2209 B.n150 B.n149 10.6151
R2210 B.n153 B.n150 10.6151
R2211 B.n154 B.n153 10.6151
R2212 B.n157 B.n154 10.6151
R2213 B.n158 B.n157 10.6151
R2214 B.n161 B.n158 10.6151
R2215 B.n162 B.n161 10.6151
R2216 B.n165 B.n162 10.6151
R2217 B.n166 B.n165 10.6151
R2218 B.n169 B.n166 10.6151
R2219 B.n170 B.n169 10.6151
R2220 B.n173 B.n170 10.6151
R2221 B.n174 B.n173 10.6151
R2222 B.n177 B.n174 10.6151
R2223 B.n178 B.n177 10.6151
R2224 B.n181 B.n178 10.6151
R2225 B.n182 B.n181 10.6151
R2226 B.n185 B.n182 10.6151
R2227 B.n186 B.n185 10.6151
R2228 B.n189 B.n186 10.6151
R2229 B.n190 B.n189 10.6151
R2230 B.n193 B.n190 10.6151
R2231 B.n194 B.n193 10.6151
R2232 B.n197 B.n194 10.6151
R2233 B.n198 B.n197 10.6151
R2234 B.n201 B.n198 10.6151
R2235 B.n202 B.n201 10.6151
R2236 B.n205 B.n202 10.6151
R2237 B.n206 B.n205 10.6151
R2238 B.n209 B.n206 10.6151
R2239 B.n210 B.n209 10.6151
R2240 B.n213 B.n210 10.6151
R2241 B.n214 B.n213 10.6151
R2242 B.n217 B.n214 10.6151
R2243 B.n218 B.n217 10.6151
R2244 B.n221 B.n218 10.6151
R2245 B.n222 B.n221 10.6151
R2246 B.n225 B.n222 10.6151
R2247 B.n226 B.n225 10.6151
R2248 B.n229 B.n226 10.6151
R2249 B.n230 B.n229 10.6151
R2250 B.n233 B.n230 10.6151
R2251 B.n234 B.n233 10.6151
R2252 B.n237 B.n234 10.6151
R2253 B.n238 B.n237 10.6151
R2254 B.n241 B.n238 10.6151
R2255 B.n242 B.n241 10.6151
R2256 B.n245 B.n242 10.6151
R2257 B.n246 B.n245 10.6151
R2258 B.n249 B.n246 10.6151
R2259 B.n250 B.n249 10.6151
R2260 B.n254 B.n253 10.6151
R2261 B.n257 B.n254 10.6151
R2262 B.n258 B.n257 10.6151
R2263 B.n261 B.n258 10.6151
R2264 B.n262 B.n261 10.6151
R2265 B.n265 B.n262 10.6151
R2266 B.n266 B.n265 10.6151
R2267 B.n269 B.n266 10.6151
R2268 B.n274 B.n271 10.6151
R2269 B.n275 B.n274 10.6151
R2270 B.n278 B.n275 10.6151
R2271 B.n279 B.n278 10.6151
R2272 B.n282 B.n279 10.6151
R2273 B.n283 B.n282 10.6151
R2274 B.n286 B.n283 10.6151
R2275 B.n287 B.n286 10.6151
R2276 B.n290 B.n287 10.6151
R2277 B.n291 B.n290 10.6151
R2278 B.n294 B.n291 10.6151
R2279 B.n295 B.n294 10.6151
R2280 B.n298 B.n295 10.6151
R2281 B.n299 B.n298 10.6151
R2282 B.n302 B.n299 10.6151
R2283 B.n303 B.n302 10.6151
R2284 B.n306 B.n303 10.6151
R2285 B.n307 B.n306 10.6151
R2286 B.n310 B.n307 10.6151
R2287 B.n311 B.n310 10.6151
R2288 B.n314 B.n311 10.6151
R2289 B.n315 B.n314 10.6151
R2290 B.n318 B.n315 10.6151
R2291 B.n319 B.n318 10.6151
R2292 B.n322 B.n319 10.6151
R2293 B.n323 B.n322 10.6151
R2294 B.n326 B.n323 10.6151
R2295 B.n327 B.n326 10.6151
R2296 B.n330 B.n327 10.6151
R2297 B.n331 B.n330 10.6151
R2298 B.n334 B.n331 10.6151
R2299 B.n335 B.n334 10.6151
R2300 B.n338 B.n335 10.6151
R2301 B.n339 B.n338 10.6151
R2302 B.n342 B.n339 10.6151
R2303 B.n343 B.n342 10.6151
R2304 B.n346 B.n343 10.6151
R2305 B.n347 B.n346 10.6151
R2306 B.n350 B.n347 10.6151
R2307 B.n351 B.n350 10.6151
R2308 B.n354 B.n351 10.6151
R2309 B.n355 B.n354 10.6151
R2310 B.n358 B.n355 10.6151
R2311 B.n359 B.n358 10.6151
R2312 B.n362 B.n359 10.6151
R2313 B.n363 B.n362 10.6151
R2314 B.n366 B.n363 10.6151
R2315 B.n367 B.n366 10.6151
R2316 B.n370 B.n367 10.6151
R2317 B.n371 B.n370 10.6151
R2318 B.n374 B.n371 10.6151
R2319 B.n375 B.n374 10.6151
R2320 B.n378 B.n375 10.6151
R2321 B.n379 B.n378 10.6151
R2322 B.n382 B.n379 10.6151
R2323 B.n383 B.n382 10.6151
R2324 B.n386 B.n383 10.6151
R2325 B.n387 B.n386 10.6151
R2326 B.n390 B.n387 10.6151
R2327 B.n391 B.n390 10.6151
R2328 B.n394 B.n391 10.6151
R2329 B.n395 B.n394 10.6151
R2330 B.n911 B.n395 10.6151
R2331 B.n801 B.n443 10.6151
R2332 B.n802 B.n801 10.6151
R2333 B.n803 B.n802 10.6151
R2334 B.n803 B.n435 10.6151
R2335 B.n813 B.n435 10.6151
R2336 B.n814 B.n813 10.6151
R2337 B.n815 B.n814 10.6151
R2338 B.n815 B.n427 10.6151
R2339 B.n825 B.n427 10.6151
R2340 B.n826 B.n825 10.6151
R2341 B.n827 B.n826 10.6151
R2342 B.n827 B.n419 10.6151
R2343 B.n837 B.n419 10.6151
R2344 B.n838 B.n837 10.6151
R2345 B.n839 B.n838 10.6151
R2346 B.n839 B.n411 10.6151
R2347 B.n849 B.n411 10.6151
R2348 B.n850 B.n849 10.6151
R2349 B.n851 B.n850 10.6151
R2350 B.n851 B.n404 10.6151
R2351 B.n862 B.n404 10.6151
R2352 B.n863 B.n862 10.6151
R2353 B.n865 B.n863 10.6151
R2354 B.n865 B.n864 10.6151
R2355 B.n864 B.n396 10.6151
R2356 B.n876 B.n396 10.6151
R2357 B.n877 B.n876 10.6151
R2358 B.n878 B.n877 10.6151
R2359 B.n879 B.n878 10.6151
R2360 B.n881 B.n879 10.6151
R2361 B.n882 B.n881 10.6151
R2362 B.n883 B.n882 10.6151
R2363 B.n884 B.n883 10.6151
R2364 B.n886 B.n884 10.6151
R2365 B.n887 B.n886 10.6151
R2366 B.n888 B.n887 10.6151
R2367 B.n889 B.n888 10.6151
R2368 B.n891 B.n889 10.6151
R2369 B.n892 B.n891 10.6151
R2370 B.n893 B.n892 10.6151
R2371 B.n894 B.n893 10.6151
R2372 B.n896 B.n894 10.6151
R2373 B.n897 B.n896 10.6151
R2374 B.n898 B.n897 10.6151
R2375 B.n899 B.n898 10.6151
R2376 B.n901 B.n899 10.6151
R2377 B.n902 B.n901 10.6151
R2378 B.n903 B.n902 10.6151
R2379 B.n904 B.n903 10.6151
R2380 B.n906 B.n904 10.6151
R2381 B.n907 B.n906 10.6151
R2382 B.n908 B.n907 10.6151
R2383 B.n909 B.n908 10.6151
R2384 B.n910 B.n909 10.6151
R2385 B.n795 B.n447 10.6151
R2386 B.n790 B.n447 10.6151
R2387 B.n790 B.n789 10.6151
R2388 B.n789 B.n788 10.6151
R2389 B.n788 B.n785 10.6151
R2390 B.n785 B.n784 10.6151
R2391 B.n784 B.n781 10.6151
R2392 B.n781 B.n780 10.6151
R2393 B.n780 B.n777 10.6151
R2394 B.n777 B.n776 10.6151
R2395 B.n776 B.n773 10.6151
R2396 B.n773 B.n772 10.6151
R2397 B.n772 B.n769 10.6151
R2398 B.n769 B.n768 10.6151
R2399 B.n768 B.n765 10.6151
R2400 B.n765 B.n764 10.6151
R2401 B.n764 B.n761 10.6151
R2402 B.n761 B.n760 10.6151
R2403 B.n760 B.n757 10.6151
R2404 B.n757 B.n756 10.6151
R2405 B.n756 B.n753 10.6151
R2406 B.n753 B.n752 10.6151
R2407 B.n752 B.n749 10.6151
R2408 B.n749 B.n748 10.6151
R2409 B.n748 B.n745 10.6151
R2410 B.n745 B.n744 10.6151
R2411 B.n744 B.n741 10.6151
R2412 B.n741 B.n740 10.6151
R2413 B.n740 B.n737 10.6151
R2414 B.n737 B.n736 10.6151
R2415 B.n736 B.n733 10.6151
R2416 B.n733 B.n732 10.6151
R2417 B.n732 B.n729 10.6151
R2418 B.n729 B.n728 10.6151
R2419 B.n728 B.n725 10.6151
R2420 B.n725 B.n724 10.6151
R2421 B.n724 B.n721 10.6151
R2422 B.n721 B.n720 10.6151
R2423 B.n720 B.n717 10.6151
R2424 B.n717 B.n716 10.6151
R2425 B.n716 B.n713 10.6151
R2426 B.n713 B.n712 10.6151
R2427 B.n712 B.n709 10.6151
R2428 B.n709 B.n708 10.6151
R2429 B.n708 B.n705 10.6151
R2430 B.n705 B.n704 10.6151
R2431 B.n704 B.n701 10.6151
R2432 B.n701 B.n700 10.6151
R2433 B.n700 B.n697 10.6151
R2434 B.n697 B.n696 10.6151
R2435 B.n696 B.n693 10.6151
R2436 B.n693 B.n692 10.6151
R2437 B.n692 B.n689 10.6151
R2438 B.n689 B.n688 10.6151
R2439 B.n688 B.n685 10.6151
R2440 B.n685 B.n684 10.6151
R2441 B.n684 B.n681 10.6151
R2442 B.n681 B.n680 10.6151
R2443 B.n680 B.n677 10.6151
R2444 B.n677 B.n676 10.6151
R2445 B.n676 B.n673 10.6151
R2446 B.n673 B.n672 10.6151
R2447 B.n672 B.n669 10.6151
R2448 B.n667 B.n664 10.6151
R2449 B.n664 B.n663 10.6151
R2450 B.n663 B.n660 10.6151
R2451 B.n660 B.n659 10.6151
R2452 B.n659 B.n656 10.6151
R2453 B.n656 B.n655 10.6151
R2454 B.n655 B.n652 10.6151
R2455 B.n652 B.n651 10.6151
R2456 B.n648 B.n647 10.6151
R2457 B.n647 B.n644 10.6151
R2458 B.n644 B.n643 10.6151
R2459 B.n643 B.n640 10.6151
R2460 B.n640 B.n639 10.6151
R2461 B.n639 B.n636 10.6151
R2462 B.n636 B.n635 10.6151
R2463 B.n635 B.n632 10.6151
R2464 B.n632 B.n631 10.6151
R2465 B.n631 B.n628 10.6151
R2466 B.n628 B.n627 10.6151
R2467 B.n627 B.n624 10.6151
R2468 B.n624 B.n623 10.6151
R2469 B.n623 B.n620 10.6151
R2470 B.n620 B.n619 10.6151
R2471 B.n619 B.n616 10.6151
R2472 B.n616 B.n615 10.6151
R2473 B.n615 B.n612 10.6151
R2474 B.n612 B.n611 10.6151
R2475 B.n611 B.n608 10.6151
R2476 B.n608 B.n607 10.6151
R2477 B.n607 B.n604 10.6151
R2478 B.n604 B.n603 10.6151
R2479 B.n603 B.n600 10.6151
R2480 B.n600 B.n599 10.6151
R2481 B.n599 B.n596 10.6151
R2482 B.n596 B.n595 10.6151
R2483 B.n595 B.n592 10.6151
R2484 B.n592 B.n591 10.6151
R2485 B.n591 B.n588 10.6151
R2486 B.n588 B.n587 10.6151
R2487 B.n587 B.n584 10.6151
R2488 B.n584 B.n583 10.6151
R2489 B.n583 B.n580 10.6151
R2490 B.n580 B.n579 10.6151
R2491 B.n579 B.n576 10.6151
R2492 B.n576 B.n575 10.6151
R2493 B.n575 B.n572 10.6151
R2494 B.n572 B.n571 10.6151
R2495 B.n571 B.n568 10.6151
R2496 B.n568 B.n567 10.6151
R2497 B.n567 B.n564 10.6151
R2498 B.n564 B.n563 10.6151
R2499 B.n563 B.n560 10.6151
R2500 B.n560 B.n559 10.6151
R2501 B.n559 B.n556 10.6151
R2502 B.n556 B.n555 10.6151
R2503 B.n555 B.n552 10.6151
R2504 B.n552 B.n551 10.6151
R2505 B.n551 B.n548 10.6151
R2506 B.n548 B.n547 10.6151
R2507 B.n547 B.n544 10.6151
R2508 B.n544 B.n543 10.6151
R2509 B.n543 B.n540 10.6151
R2510 B.n540 B.n539 10.6151
R2511 B.n539 B.n536 10.6151
R2512 B.n536 B.n535 10.6151
R2513 B.n535 B.n532 10.6151
R2514 B.n532 B.n531 10.6151
R2515 B.n531 B.n528 10.6151
R2516 B.n528 B.n527 10.6151
R2517 B.n527 B.n524 10.6151
R2518 B.n524 B.n523 10.6151
R2519 B.n797 B.n796 10.6151
R2520 B.n797 B.n439 10.6151
R2521 B.n807 B.n439 10.6151
R2522 B.n808 B.n807 10.6151
R2523 B.n809 B.n808 10.6151
R2524 B.n809 B.n431 10.6151
R2525 B.n819 B.n431 10.6151
R2526 B.n820 B.n819 10.6151
R2527 B.n821 B.n820 10.6151
R2528 B.n821 B.n423 10.6151
R2529 B.n831 B.n423 10.6151
R2530 B.n832 B.n831 10.6151
R2531 B.n833 B.n832 10.6151
R2532 B.n833 B.n415 10.6151
R2533 B.n843 B.n415 10.6151
R2534 B.n844 B.n843 10.6151
R2535 B.n845 B.n844 10.6151
R2536 B.n845 B.n407 10.6151
R2537 B.n856 B.n407 10.6151
R2538 B.n857 B.n856 10.6151
R2539 B.n858 B.n857 10.6151
R2540 B.n858 B.n400 10.6151
R2541 B.n869 B.n400 10.6151
R2542 B.n870 B.n869 10.6151
R2543 B.n871 B.n870 10.6151
R2544 B.n871 B.n0 10.6151
R2545 B.n966 B.n1 10.6151
R2546 B.n966 B.n965 10.6151
R2547 B.n965 B.n964 10.6151
R2548 B.n964 B.n10 10.6151
R2549 B.n958 B.n10 10.6151
R2550 B.n958 B.n957 10.6151
R2551 B.n957 B.n956 10.6151
R2552 B.n956 B.n16 10.6151
R2553 B.n950 B.n16 10.6151
R2554 B.n950 B.n949 10.6151
R2555 B.n949 B.n948 10.6151
R2556 B.n948 B.n24 10.6151
R2557 B.n942 B.n24 10.6151
R2558 B.n942 B.n941 10.6151
R2559 B.n941 B.n940 10.6151
R2560 B.n940 B.n31 10.6151
R2561 B.n934 B.n31 10.6151
R2562 B.n934 B.n933 10.6151
R2563 B.n933 B.n932 10.6151
R2564 B.n932 B.n38 10.6151
R2565 B.n926 B.n38 10.6151
R2566 B.n926 B.n925 10.6151
R2567 B.n925 B.n924 10.6151
R2568 B.n924 B.n45 10.6151
R2569 B.n918 B.n45 10.6151
R2570 B.n918 B.n917 10.6151
R2571 B.n253 B.n127 6.5566
R2572 B.n270 B.n269 6.5566
R2573 B.n668 B.n667 6.5566
R2574 B.n651 B.n521 6.5566
R2575 B.n250 B.n127 4.05904
R2576 B.n271 B.n270 4.05904
R2577 B.n669 B.n668 4.05904
R2578 B.n648 B.n521 4.05904
R2579 B.n972 B.n0 2.81026
R2580 B.n972 B.n1 2.81026
R2581 B.t7 B.n429 1.7772
R2582 B.t3 B.n36 1.7772
R2583 VN VN.t0 254.194
R2584 VN VN.t1 203.496
R2585 VDD2.n205 VDD2.n105 214.453
R2586 VDD2.n100 VDD2.n0 214.453
R2587 VDD2.n206 VDD2.n205 185
R2588 VDD2.n204 VDD2.n203 185
R2589 VDD2.n109 VDD2.n108 185
R2590 VDD2.n198 VDD2.n197 185
R2591 VDD2.n196 VDD2.n195 185
R2592 VDD2.n113 VDD2.n112 185
R2593 VDD2.n190 VDD2.n189 185
R2594 VDD2.n188 VDD2.n187 185
R2595 VDD2.n117 VDD2.n116 185
R2596 VDD2.n182 VDD2.n181 185
R2597 VDD2.n180 VDD2.n179 185
R2598 VDD2.n121 VDD2.n120 185
R2599 VDD2.n174 VDD2.n173 185
R2600 VDD2.n172 VDD2.n171 185
R2601 VDD2.n125 VDD2.n124 185
R2602 VDD2.n166 VDD2.n165 185
R2603 VDD2.n164 VDD2.n163 185
R2604 VDD2.n162 VDD2.n128 185
R2605 VDD2.n132 VDD2.n129 185
R2606 VDD2.n157 VDD2.n156 185
R2607 VDD2.n155 VDD2.n154 185
R2608 VDD2.n134 VDD2.n133 185
R2609 VDD2.n149 VDD2.n148 185
R2610 VDD2.n147 VDD2.n146 185
R2611 VDD2.n138 VDD2.n137 185
R2612 VDD2.n141 VDD2.n140 185
R2613 VDD2.n35 VDD2.n34 185
R2614 VDD2.n32 VDD2.n31 185
R2615 VDD2.n41 VDD2.n40 185
R2616 VDD2.n43 VDD2.n42 185
R2617 VDD2.n28 VDD2.n27 185
R2618 VDD2.n49 VDD2.n48 185
R2619 VDD2.n52 VDD2.n51 185
R2620 VDD2.n50 VDD2.n24 185
R2621 VDD2.n57 VDD2.n23 185
R2622 VDD2.n59 VDD2.n58 185
R2623 VDD2.n61 VDD2.n60 185
R2624 VDD2.n20 VDD2.n19 185
R2625 VDD2.n67 VDD2.n66 185
R2626 VDD2.n69 VDD2.n68 185
R2627 VDD2.n16 VDD2.n15 185
R2628 VDD2.n75 VDD2.n74 185
R2629 VDD2.n77 VDD2.n76 185
R2630 VDD2.n12 VDD2.n11 185
R2631 VDD2.n83 VDD2.n82 185
R2632 VDD2.n85 VDD2.n84 185
R2633 VDD2.n8 VDD2.n7 185
R2634 VDD2.n91 VDD2.n90 185
R2635 VDD2.n93 VDD2.n92 185
R2636 VDD2.n4 VDD2.n3 185
R2637 VDD2.n99 VDD2.n98 185
R2638 VDD2.n101 VDD2.n100 185
R2639 VDD2.t1 VDD2.n139 149.524
R2640 VDD2.t0 VDD2.n33 149.524
R2641 VDD2.n205 VDD2.n204 104.615
R2642 VDD2.n204 VDD2.n108 104.615
R2643 VDD2.n197 VDD2.n108 104.615
R2644 VDD2.n197 VDD2.n196 104.615
R2645 VDD2.n196 VDD2.n112 104.615
R2646 VDD2.n189 VDD2.n112 104.615
R2647 VDD2.n189 VDD2.n188 104.615
R2648 VDD2.n188 VDD2.n116 104.615
R2649 VDD2.n181 VDD2.n116 104.615
R2650 VDD2.n181 VDD2.n180 104.615
R2651 VDD2.n180 VDD2.n120 104.615
R2652 VDD2.n173 VDD2.n120 104.615
R2653 VDD2.n173 VDD2.n172 104.615
R2654 VDD2.n172 VDD2.n124 104.615
R2655 VDD2.n165 VDD2.n124 104.615
R2656 VDD2.n165 VDD2.n164 104.615
R2657 VDD2.n164 VDD2.n128 104.615
R2658 VDD2.n132 VDD2.n128 104.615
R2659 VDD2.n156 VDD2.n132 104.615
R2660 VDD2.n156 VDD2.n155 104.615
R2661 VDD2.n155 VDD2.n133 104.615
R2662 VDD2.n148 VDD2.n133 104.615
R2663 VDD2.n148 VDD2.n147 104.615
R2664 VDD2.n147 VDD2.n137 104.615
R2665 VDD2.n140 VDD2.n137 104.615
R2666 VDD2.n34 VDD2.n31 104.615
R2667 VDD2.n41 VDD2.n31 104.615
R2668 VDD2.n42 VDD2.n41 104.615
R2669 VDD2.n42 VDD2.n27 104.615
R2670 VDD2.n49 VDD2.n27 104.615
R2671 VDD2.n51 VDD2.n49 104.615
R2672 VDD2.n51 VDD2.n50 104.615
R2673 VDD2.n50 VDD2.n23 104.615
R2674 VDD2.n59 VDD2.n23 104.615
R2675 VDD2.n60 VDD2.n59 104.615
R2676 VDD2.n60 VDD2.n19 104.615
R2677 VDD2.n67 VDD2.n19 104.615
R2678 VDD2.n68 VDD2.n67 104.615
R2679 VDD2.n68 VDD2.n15 104.615
R2680 VDD2.n75 VDD2.n15 104.615
R2681 VDD2.n76 VDD2.n75 104.615
R2682 VDD2.n76 VDD2.n11 104.615
R2683 VDD2.n83 VDD2.n11 104.615
R2684 VDD2.n84 VDD2.n83 104.615
R2685 VDD2.n84 VDD2.n7 104.615
R2686 VDD2.n91 VDD2.n7 104.615
R2687 VDD2.n92 VDD2.n91 104.615
R2688 VDD2.n92 VDD2.n3 104.615
R2689 VDD2.n99 VDD2.n3 104.615
R2690 VDD2.n100 VDD2.n99 104.615
R2691 VDD2.n210 VDD2.n104 98.1912
R2692 VDD2.n140 VDD2.t1 52.3082
R2693 VDD2.n34 VDD2.t0 52.3082
R2694 VDD2.n210 VDD2.n209 52.1611
R2695 VDD2.n163 VDD2.n162 13.1884
R2696 VDD2.n58 VDD2.n57 13.1884
R2697 VDD2.n207 VDD2.n206 12.8005
R2698 VDD2.n166 VDD2.n127 12.8005
R2699 VDD2.n161 VDD2.n129 12.8005
R2700 VDD2.n56 VDD2.n24 12.8005
R2701 VDD2.n61 VDD2.n22 12.8005
R2702 VDD2.n102 VDD2.n101 12.8005
R2703 VDD2.n203 VDD2.n107 12.0247
R2704 VDD2.n167 VDD2.n125 12.0247
R2705 VDD2.n158 VDD2.n157 12.0247
R2706 VDD2.n53 VDD2.n52 12.0247
R2707 VDD2.n62 VDD2.n20 12.0247
R2708 VDD2.n98 VDD2.n2 12.0247
R2709 VDD2.n202 VDD2.n109 11.249
R2710 VDD2.n171 VDD2.n170 11.249
R2711 VDD2.n154 VDD2.n131 11.249
R2712 VDD2.n48 VDD2.n26 11.249
R2713 VDD2.n66 VDD2.n65 11.249
R2714 VDD2.n97 VDD2.n4 11.249
R2715 VDD2.n199 VDD2.n198 10.4732
R2716 VDD2.n174 VDD2.n123 10.4732
R2717 VDD2.n153 VDD2.n134 10.4732
R2718 VDD2.n47 VDD2.n28 10.4732
R2719 VDD2.n69 VDD2.n18 10.4732
R2720 VDD2.n94 VDD2.n93 10.4732
R2721 VDD2.n141 VDD2.n139 10.2747
R2722 VDD2.n35 VDD2.n33 10.2747
R2723 VDD2.n195 VDD2.n111 9.69747
R2724 VDD2.n175 VDD2.n121 9.69747
R2725 VDD2.n150 VDD2.n149 9.69747
R2726 VDD2.n44 VDD2.n43 9.69747
R2727 VDD2.n70 VDD2.n16 9.69747
R2728 VDD2.n90 VDD2.n6 9.69747
R2729 VDD2.n209 VDD2.n208 9.45567
R2730 VDD2.n104 VDD2.n103 9.45567
R2731 VDD2.n143 VDD2.n142 9.3005
R2732 VDD2.n145 VDD2.n144 9.3005
R2733 VDD2.n136 VDD2.n135 9.3005
R2734 VDD2.n151 VDD2.n150 9.3005
R2735 VDD2.n153 VDD2.n152 9.3005
R2736 VDD2.n131 VDD2.n130 9.3005
R2737 VDD2.n159 VDD2.n158 9.3005
R2738 VDD2.n161 VDD2.n160 9.3005
R2739 VDD2.n115 VDD2.n114 9.3005
R2740 VDD2.n192 VDD2.n191 9.3005
R2741 VDD2.n194 VDD2.n193 9.3005
R2742 VDD2.n111 VDD2.n110 9.3005
R2743 VDD2.n200 VDD2.n199 9.3005
R2744 VDD2.n202 VDD2.n201 9.3005
R2745 VDD2.n107 VDD2.n106 9.3005
R2746 VDD2.n208 VDD2.n207 9.3005
R2747 VDD2.n186 VDD2.n185 9.3005
R2748 VDD2.n184 VDD2.n183 9.3005
R2749 VDD2.n119 VDD2.n118 9.3005
R2750 VDD2.n178 VDD2.n177 9.3005
R2751 VDD2.n176 VDD2.n175 9.3005
R2752 VDD2.n123 VDD2.n122 9.3005
R2753 VDD2.n170 VDD2.n169 9.3005
R2754 VDD2.n168 VDD2.n167 9.3005
R2755 VDD2.n127 VDD2.n126 9.3005
R2756 VDD2.n79 VDD2.n78 9.3005
R2757 VDD2.n14 VDD2.n13 9.3005
R2758 VDD2.n73 VDD2.n72 9.3005
R2759 VDD2.n71 VDD2.n70 9.3005
R2760 VDD2.n18 VDD2.n17 9.3005
R2761 VDD2.n65 VDD2.n64 9.3005
R2762 VDD2.n63 VDD2.n62 9.3005
R2763 VDD2.n22 VDD2.n21 9.3005
R2764 VDD2.n37 VDD2.n36 9.3005
R2765 VDD2.n39 VDD2.n38 9.3005
R2766 VDD2.n30 VDD2.n29 9.3005
R2767 VDD2.n45 VDD2.n44 9.3005
R2768 VDD2.n47 VDD2.n46 9.3005
R2769 VDD2.n26 VDD2.n25 9.3005
R2770 VDD2.n54 VDD2.n53 9.3005
R2771 VDD2.n56 VDD2.n55 9.3005
R2772 VDD2.n81 VDD2.n80 9.3005
R2773 VDD2.n10 VDD2.n9 9.3005
R2774 VDD2.n87 VDD2.n86 9.3005
R2775 VDD2.n89 VDD2.n88 9.3005
R2776 VDD2.n6 VDD2.n5 9.3005
R2777 VDD2.n95 VDD2.n94 9.3005
R2778 VDD2.n97 VDD2.n96 9.3005
R2779 VDD2.n2 VDD2.n1 9.3005
R2780 VDD2.n103 VDD2.n102 9.3005
R2781 VDD2.n194 VDD2.n113 8.92171
R2782 VDD2.n179 VDD2.n178 8.92171
R2783 VDD2.n146 VDD2.n136 8.92171
R2784 VDD2.n40 VDD2.n30 8.92171
R2785 VDD2.n74 VDD2.n73 8.92171
R2786 VDD2.n89 VDD2.n8 8.92171
R2787 VDD2.n209 VDD2.n105 8.2187
R2788 VDD2.n104 VDD2.n0 8.2187
R2789 VDD2.n191 VDD2.n190 8.14595
R2790 VDD2.n182 VDD2.n119 8.14595
R2791 VDD2.n145 VDD2.n138 8.14595
R2792 VDD2.n39 VDD2.n32 8.14595
R2793 VDD2.n77 VDD2.n14 8.14595
R2794 VDD2.n86 VDD2.n85 8.14595
R2795 VDD2.n187 VDD2.n115 7.3702
R2796 VDD2.n183 VDD2.n117 7.3702
R2797 VDD2.n142 VDD2.n141 7.3702
R2798 VDD2.n36 VDD2.n35 7.3702
R2799 VDD2.n78 VDD2.n12 7.3702
R2800 VDD2.n82 VDD2.n10 7.3702
R2801 VDD2.n187 VDD2.n186 6.59444
R2802 VDD2.n186 VDD2.n117 6.59444
R2803 VDD2.n81 VDD2.n12 6.59444
R2804 VDD2.n82 VDD2.n81 6.59444
R2805 VDD2.n190 VDD2.n115 5.81868
R2806 VDD2.n183 VDD2.n182 5.81868
R2807 VDD2.n142 VDD2.n138 5.81868
R2808 VDD2.n36 VDD2.n32 5.81868
R2809 VDD2.n78 VDD2.n77 5.81868
R2810 VDD2.n85 VDD2.n10 5.81868
R2811 VDD2.n207 VDD2.n105 5.3904
R2812 VDD2.n102 VDD2.n0 5.3904
R2813 VDD2.n191 VDD2.n113 5.04292
R2814 VDD2.n179 VDD2.n119 5.04292
R2815 VDD2.n146 VDD2.n145 5.04292
R2816 VDD2.n40 VDD2.n39 5.04292
R2817 VDD2.n74 VDD2.n14 5.04292
R2818 VDD2.n86 VDD2.n8 5.04292
R2819 VDD2.n195 VDD2.n194 4.26717
R2820 VDD2.n178 VDD2.n121 4.26717
R2821 VDD2.n149 VDD2.n136 4.26717
R2822 VDD2.n43 VDD2.n30 4.26717
R2823 VDD2.n73 VDD2.n16 4.26717
R2824 VDD2.n90 VDD2.n89 4.26717
R2825 VDD2.n198 VDD2.n111 3.49141
R2826 VDD2.n175 VDD2.n174 3.49141
R2827 VDD2.n150 VDD2.n134 3.49141
R2828 VDD2.n44 VDD2.n28 3.49141
R2829 VDD2.n70 VDD2.n69 3.49141
R2830 VDD2.n93 VDD2.n6 3.49141
R2831 VDD2.n37 VDD2.n33 2.84303
R2832 VDD2.n143 VDD2.n139 2.84303
R2833 VDD2.n199 VDD2.n109 2.71565
R2834 VDD2.n171 VDD2.n123 2.71565
R2835 VDD2.n154 VDD2.n153 2.71565
R2836 VDD2.n48 VDD2.n47 2.71565
R2837 VDD2.n66 VDD2.n18 2.71565
R2838 VDD2.n94 VDD2.n4 2.71565
R2839 VDD2.n203 VDD2.n202 1.93989
R2840 VDD2.n170 VDD2.n125 1.93989
R2841 VDD2.n157 VDD2.n131 1.93989
R2842 VDD2.n52 VDD2.n26 1.93989
R2843 VDD2.n65 VDD2.n20 1.93989
R2844 VDD2.n98 VDD2.n97 1.93989
R2845 VDD2.n206 VDD2.n107 1.16414
R2846 VDD2.n167 VDD2.n166 1.16414
R2847 VDD2.n158 VDD2.n129 1.16414
R2848 VDD2.n53 VDD2.n24 1.16414
R2849 VDD2.n62 VDD2.n61 1.16414
R2850 VDD2.n101 VDD2.n2 1.16414
R2851 VDD2 VDD2.n210 0.75481
R2852 VDD2.n163 VDD2.n127 0.388379
R2853 VDD2.n162 VDD2.n161 0.388379
R2854 VDD2.n57 VDD2.n56 0.388379
R2855 VDD2.n58 VDD2.n22 0.388379
R2856 VDD2.n208 VDD2.n106 0.155672
R2857 VDD2.n201 VDD2.n106 0.155672
R2858 VDD2.n201 VDD2.n200 0.155672
R2859 VDD2.n200 VDD2.n110 0.155672
R2860 VDD2.n193 VDD2.n110 0.155672
R2861 VDD2.n193 VDD2.n192 0.155672
R2862 VDD2.n192 VDD2.n114 0.155672
R2863 VDD2.n185 VDD2.n114 0.155672
R2864 VDD2.n185 VDD2.n184 0.155672
R2865 VDD2.n184 VDD2.n118 0.155672
R2866 VDD2.n177 VDD2.n118 0.155672
R2867 VDD2.n177 VDD2.n176 0.155672
R2868 VDD2.n176 VDD2.n122 0.155672
R2869 VDD2.n169 VDD2.n122 0.155672
R2870 VDD2.n169 VDD2.n168 0.155672
R2871 VDD2.n168 VDD2.n126 0.155672
R2872 VDD2.n160 VDD2.n126 0.155672
R2873 VDD2.n160 VDD2.n159 0.155672
R2874 VDD2.n159 VDD2.n130 0.155672
R2875 VDD2.n152 VDD2.n130 0.155672
R2876 VDD2.n152 VDD2.n151 0.155672
R2877 VDD2.n151 VDD2.n135 0.155672
R2878 VDD2.n144 VDD2.n135 0.155672
R2879 VDD2.n144 VDD2.n143 0.155672
R2880 VDD2.n38 VDD2.n37 0.155672
R2881 VDD2.n38 VDD2.n29 0.155672
R2882 VDD2.n45 VDD2.n29 0.155672
R2883 VDD2.n46 VDD2.n45 0.155672
R2884 VDD2.n46 VDD2.n25 0.155672
R2885 VDD2.n54 VDD2.n25 0.155672
R2886 VDD2.n55 VDD2.n54 0.155672
R2887 VDD2.n55 VDD2.n21 0.155672
R2888 VDD2.n63 VDD2.n21 0.155672
R2889 VDD2.n64 VDD2.n63 0.155672
R2890 VDD2.n64 VDD2.n17 0.155672
R2891 VDD2.n71 VDD2.n17 0.155672
R2892 VDD2.n72 VDD2.n71 0.155672
R2893 VDD2.n72 VDD2.n13 0.155672
R2894 VDD2.n79 VDD2.n13 0.155672
R2895 VDD2.n80 VDD2.n79 0.155672
R2896 VDD2.n80 VDD2.n9 0.155672
R2897 VDD2.n87 VDD2.n9 0.155672
R2898 VDD2.n88 VDD2.n87 0.155672
R2899 VDD2.n88 VDD2.n5 0.155672
R2900 VDD2.n95 VDD2.n5 0.155672
R2901 VDD2.n96 VDD2.n95 0.155672
R2902 VDD2.n96 VDD2.n1 0.155672
R2903 VDD2.n103 VDD2.n1 0.155672
C0 VDD2 VN 4.43174f
C1 VDD2 VTAIL 7.10693f
C2 VDD1 VN 0.14826f
C3 VDD1 VTAIL 7.05557f
C4 VP VN 6.98355f
C5 VDD1 VDD2 0.711725f
C6 VP VTAIL 3.79992f
C7 VDD2 VP 0.346212f
C8 VDD1 VP 4.62611f
C9 VN VTAIL 3.78556f
C10 VDD2 B 5.877414f
C11 VDD1 B 9.24822f
C12 VTAIL B 10.558885f
C13 VN B 12.773499f
C14 VP B 7.274028f
C15 VDD2.n0 B 0.027341f
C16 VDD2.n1 B 0.019824f
C17 VDD2.n2 B 0.010652f
C18 VDD2.n3 B 0.025178f
C19 VDD2.n4 B 0.011279f
C20 VDD2.n5 B 0.019824f
C21 VDD2.n6 B 0.010652f
C22 VDD2.n7 B 0.025178f
C23 VDD2.n8 B 0.011279f
C24 VDD2.n9 B 0.019824f
C25 VDD2.n10 B 0.010652f
C26 VDD2.n11 B 0.025178f
C27 VDD2.n12 B 0.011279f
C28 VDD2.n13 B 0.019824f
C29 VDD2.n14 B 0.010652f
C30 VDD2.n15 B 0.025178f
C31 VDD2.n16 B 0.011279f
C32 VDD2.n17 B 0.019824f
C33 VDD2.n18 B 0.010652f
C34 VDD2.n19 B 0.025178f
C35 VDD2.n20 B 0.011279f
C36 VDD2.n21 B 0.019824f
C37 VDD2.n22 B 0.010652f
C38 VDD2.n23 B 0.025178f
C39 VDD2.n24 B 0.011279f
C40 VDD2.n25 B 0.019824f
C41 VDD2.n26 B 0.010652f
C42 VDD2.n27 B 0.025178f
C43 VDD2.n28 B 0.011279f
C44 VDD2.n29 B 0.019824f
C45 VDD2.n30 B 0.010652f
C46 VDD2.n31 B 0.025178f
C47 VDD2.n32 B 0.011279f
C48 VDD2.n33 B 0.19993f
C49 VDD2.t0 B 0.043324f
C50 VDD2.n34 B 0.018884f
C51 VDD2.n35 B 0.017799f
C52 VDD2.n36 B 0.010652f
C53 VDD2.n37 B 1.66048f
C54 VDD2.n38 B 0.019824f
C55 VDD2.n39 B 0.010652f
C56 VDD2.n40 B 0.011279f
C57 VDD2.n41 B 0.025178f
C58 VDD2.n42 B 0.025178f
C59 VDD2.n43 B 0.011279f
C60 VDD2.n44 B 0.010652f
C61 VDD2.n45 B 0.019824f
C62 VDD2.n46 B 0.019824f
C63 VDD2.n47 B 0.010652f
C64 VDD2.n48 B 0.011279f
C65 VDD2.n49 B 0.025178f
C66 VDD2.n50 B 0.025178f
C67 VDD2.n51 B 0.025178f
C68 VDD2.n52 B 0.011279f
C69 VDD2.n53 B 0.010652f
C70 VDD2.n54 B 0.019824f
C71 VDD2.n55 B 0.019824f
C72 VDD2.n56 B 0.010652f
C73 VDD2.n57 B 0.010966f
C74 VDD2.n58 B 0.010966f
C75 VDD2.n59 B 0.025178f
C76 VDD2.n60 B 0.025178f
C77 VDD2.n61 B 0.011279f
C78 VDD2.n62 B 0.010652f
C79 VDD2.n63 B 0.019824f
C80 VDD2.n64 B 0.019824f
C81 VDD2.n65 B 0.010652f
C82 VDD2.n66 B 0.011279f
C83 VDD2.n67 B 0.025178f
C84 VDD2.n68 B 0.025178f
C85 VDD2.n69 B 0.011279f
C86 VDD2.n70 B 0.010652f
C87 VDD2.n71 B 0.019824f
C88 VDD2.n72 B 0.019824f
C89 VDD2.n73 B 0.010652f
C90 VDD2.n74 B 0.011279f
C91 VDD2.n75 B 0.025178f
C92 VDD2.n76 B 0.025178f
C93 VDD2.n77 B 0.011279f
C94 VDD2.n78 B 0.010652f
C95 VDD2.n79 B 0.019824f
C96 VDD2.n80 B 0.019824f
C97 VDD2.n81 B 0.010652f
C98 VDD2.n82 B 0.011279f
C99 VDD2.n83 B 0.025178f
C100 VDD2.n84 B 0.025178f
C101 VDD2.n85 B 0.011279f
C102 VDD2.n86 B 0.010652f
C103 VDD2.n87 B 0.019824f
C104 VDD2.n88 B 0.019824f
C105 VDD2.n89 B 0.010652f
C106 VDD2.n90 B 0.011279f
C107 VDD2.n91 B 0.025178f
C108 VDD2.n92 B 0.025178f
C109 VDD2.n93 B 0.011279f
C110 VDD2.n94 B 0.010652f
C111 VDD2.n95 B 0.019824f
C112 VDD2.n96 B 0.019824f
C113 VDD2.n97 B 0.010652f
C114 VDD2.n98 B 0.011279f
C115 VDD2.n99 B 0.025178f
C116 VDD2.n100 B 0.051763f
C117 VDD2.n101 B 0.011279f
C118 VDD2.n102 B 0.020829f
C119 VDD2.n103 B 0.050425f
C120 VDD2.n104 B 0.82279f
C121 VDD2.n105 B 0.027341f
C122 VDD2.n106 B 0.019824f
C123 VDD2.n107 B 0.010652f
C124 VDD2.n108 B 0.025178f
C125 VDD2.n109 B 0.011279f
C126 VDD2.n110 B 0.019824f
C127 VDD2.n111 B 0.010652f
C128 VDD2.n112 B 0.025178f
C129 VDD2.n113 B 0.011279f
C130 VDD2.n114 B 0.019824f
C131 VDD2.n115 B 0.010652f
C132 VDD2.n116 B 0.025178f
C133 VDD2.n117 B 0.011279f
C134 VDD2.n118 B 0.019824f
C135 VDD2.n119 B 0.010652f
C136 VDD2.n120 B 0.025178f
C137 VDD2.n121 B 0.011279f
C138 VDD2.n122 B 0.019824f
C139 VDD2.n123 B 0.010652f
C140 VDD2.n124 B 0.025178f
C141 VDD2.n125 B 0.011279f
C142 VDD2.n126 B 0.019824f
C143 VDD2.n127 B 0.010652f
C144 VDD2.n128 B 0.025178f
C145 VDD2.n129 B 0.011279f
C146 VDD2.n130 B 0.019824f
C147 VDD2.n131 B 0.010652f
C148 VDD2.n132 B 0.025178f
C149 VDD2.n133 B 0.025178f
C150 VDD2.n134 B 0.011279f
C151 VDD2.n135 B 0.019824f
C152 VDD2.n136 B 0.010652f
C153 VDD2.n137 B 0.025178f
C154 VDD2.n138 B 0.011279f
C155 VDD2.n139 B 0.19993f
C156 VDD2.t1 B 0.043324f
C157 VDD2.n140 B 0.018884f
C158 VDD2.n141 B 0.017799f
C159 VDD2.n142 B 0.010652f
C160 VDD2.n143 B 1.66048f
C161 VDD2.n144 B 0.019824f
C162 VDD2.n145 B 0.010652f
C163 VDD2.n146 B 0.011279f
C164 VDD2.n147 B 0.025178f
C165 VDD2.n148 B 0.025178f
C166 VDD2.n149 B 0.011279f
C167 VDD2.n150 B 0.010652f
C168 VDD2.n151 B 0.019824f
C169 VDD2.n152 B 0.019824f
C170 VDD2.n153 B 0.010652f
C171 VDD2.n154 B 0.011279f
C172 VDD2.n155 B 0.025178f
C173 VDD2.n156 B 0.025178f
C174 VDD2.n157 B 0.011279f
C175 VDD2.n158 B 0.010652f
C176 VDD2.n159 B 0.019824f
C177 VDD2.n160 B 0.019824f
C178 VDD2.n161 B 0.010652f
C179 VDD2.n162 B 0.010966f
C180 VDD2.n163 B 0.010966f
C181 VDD2.n164 B 0.025178f
C182 VDD2.n165 B 0.025178f
C183 VDD2.n166 B 0.011279f
C184 VDD2.n167 B 0.010652f
C185 VDD2.n168 B 0.019824f
C186 VDD2.n169 B 0.019824f
C187 VDD2.n170 B 0.010652f
C188 VDD2.n171 B 0.011279f
C189 VDD2.n172 B 0.025178f
C190 VDD2.n173 B 0.025178f
C191 VDD2.n174 B 0.011279f
C192 VDD2.n175 B 0.010652f
C193 VDD2.n176 B 0.019824f
C194 VDD2.n177 B 0.019824f
C195 VDD2.n178 B 0.010652f
C196 VDD2.n179 B 0.011279f
C197 VDD2.n180 B 0.025178f
C198 VDD2.n181 B 0.025178f
C199 VDD2.n182 B 0.011279f
C200 VDD2.n183 B 0.010652f
C201 VDD2.n184 B 0.019824f
C202 VDD2.n185 B 0.019824f
C203 VDD2.n186 B 0.010652f
C204 VDD2.n187 B 0.011279f
C205 VDD2.n188 B 0.025178f
C206 VDD2.n189 B 0.025178f
C207 VDD2.n190 B 0.011279f
C208 VDD2.n191 B 0.010652f
C209 VDD2.n192 B 0.019824f
C210 VDD2.n193 B 0.019824f
C211 VDD2.n194 B 0.010652f
C212 VDD2.n195 B 0.011279f
C213 VDD2.n196 B 0.025178f
C214 VDD2.n197 B 0.025178f
C215 VDD2.n198 B 0.011279f
C216 VDD2.n199 B 0.010652f
C217 VDD2.n200 B 0.019824f
C218 VDD2.n201 B 0.019824f
C219 VDD2.n202 B 0.010652f
C220 VDD2.n203 B 0.011279f
C221 VDD2.n204 B 0.025178f
C222 VDD2.n205 B 0.051763f
C223 VDD2.n206 B 0.011279f
C224 VDD2.n207 B 0.020829f
C225 VDD2.n208 B 0.050425f
C226 VDD2.n209 B 0.067415f
C227 VDD2.n210 B 3.09612f
C228 VN.t1 B 4.57177f
C229 VN.t0 B 5.17381f
C230 VDD1.n0 B 0.02764f
C231 VDD1.n1 B 0.020041f
C232 VDD1.n2 B 0.010769f
C233 VDD1.n3 B 0.025454f
C234 VDD1.n4 B 0.011402f
C235 VDD1.n5 B 0.020041f
C236 VDD1.n6 B 0.010769f
C237 VDD1.n7 B 0.025454f
C238 VDD1.n8 B 0.011402f
C239 VDD1.n9 B 0.020041f
C240 VDD1.n10 B 0.010769f
C241 VDD1.n11 B 0.025454f
C242 VDD1.n12 B 0.011402f
C243 VDD1.n13 B 0.020041f
C244 VDD1.n14 B 0.010769f
C245 VDD1.n15 B 0.025454f
C246 VDD1.n16 B 0.011402f
C247 VDD1.n17 B 0.020041f
C248 VDD1.n18 B 0.010769f
C249 VDD1.n19 B 0.025454f
C250 VDD1.n20 B 0.011402f
C251 VDD1.n21 B 0.020041f
C252 VDD1.n22 B 0.010769f
C253 VDD1.n23 B 0.025454f
C254 VDD1.n24 B 0.011402f
C255 VDD1.n25 B 0.020041f
C256 VDD1.n26 B 0.010769f
C257 VDD1.n27 B 0.025454f
C258 VDD1.n28 B 0.025454f
C259 VDD1.n29 B 0.011402f
C260 VDD1.n30 B 0.020041f
C261 VDD1.n31 B 0.010769f
C262 VDD1.n32 B 0.025454f
C263 VDD1.n33 B 0.011402f
C264 VDD1.n34 B 0.20212f
C265 VDD1.t1 B 0.043799f
C266 VDD1.n35 B 0.019091f
C267 VDD1.n36 B 0.017994f
C268 VDD1.n37 B 0.010769f
C269 VDD1.n38 B 1.67867f
C270 VDD1.n39 B 0.020041f
C271 VDD1.n40 B 0.010769f
C272 VDD1.n41 B 0.011402f
C273 VDD1.n42 B 0.025454f
C274 VDD1.n43 B 0.025454f
C275 VDD1.n44 B 0.011402f
C276 VDD1.n45 B 0.010769f
C277 VDD1.n46 B 0.020041f
C278 VDD1.n47 B 0.020041f
C279 VDD1.n48 B 0.010769f
C280 VDD1.n49 B 0.011402f
C281 VDD1.n50 B 0.025454f
C282 VDD1.n51 B 0.025454f
C283 VDD1.n52 B 0.011402f
C284 VDD1.n53 B 0.010769f
C285 VDD1.n54 B 0.020041f
C286 VDD1.n55 B 0.020041f
C287 VDD1.n56 B 0.010769f
C288 VDD1.n57 B 0.011086f
C289 VDD1.n58 B 0.011086f
C290 VDD1.n59 B 0.025454f
C291 VDD1.n60 B 0.025454f
C292 VDD1.n61 B 0.011402f
C293 VDD1.n62 B 0.010769f
C294 VDD1.n63 B 0.020041f
C295 VDD1.n64 B 0.020041f
C296 VDD1.n65 B 0.010769f
C297 VDD1.n66 B 0.011402f
C298 VDD1.n67 B 0.025454f
C299 VDD1.n68 B 0.025454f
C300 VDD1.n69 B 0.011402f
C301 VDD1.n70 B 0.010769f
C302 VDD1.n71 B 0.020041f
C303 VDD1.n72 B 0.020041f
C304 VDD1.n73 B 0.010769f
C305 VDD1.n74 B 0.011402f
C306 VDD1.n75 B 0.025454f
C307 VDD1.n76 B 0.025454f
C308 VDD1.n77 B 0.011402f
C309 VDD1.n78 B 0.010769f
C310 VDD1.n79 B 0.020041f
C311 VDD1.n80 B 0.020041f
C312 VDD1.n81 B 0.010769f
C313 VDD1.n82 B 0.011402f
C314 VDD1.n83 B 0.025454f
C315 VDD1.n84 B 0.025454f
C316 VDD1.n85 B 0.011402f
C317 VDD1.n86 B 0.010769f
C318 VDD1.n87 B 0.020041f
C319 VDD1.n88 B 0.020041f
C320 VDD1.n89 B 0.010769f
C321 VDD1.n90 B 0.011402f
C322 VDD1.n91 B 0.025454f
C323 VDD1.n92 B 0.025454f
C324 VDD1.n93 B 0.011402f
C325 VDD1.n94 B 0.010769f
C326 VDD1.n95 B 0.020041f
C327 VDD1.n96 B 0.020041f
C328 VDD1.n97 B 0.010769f
C329 VDD1.n98 B 0.011402f
C330 VDD1.n99 B 0.025454f
C331 VDD1.n100 B 0.05233f
C332 VDD1.n101 B 0.011402f
C333 VDD1.n102 B 0.021057f
C334 VDD1.n103 B 0.050977f
C335 VDD1.n104 B 0.069436f
C336 VDD1.n105 B 0.02764f
C337 VDD1.n106 B 0.020041f
C338 VDD1.n107 B 0.010769f
C339 VDD1.n108 B 0.025454f
C340 VDD1.n109 B 0.011402f
C341 VDD1.n110 B 0.020041f
C342 VDD1.n111 B 0.010769f
C343 VDD1.n112 B 0.025454f
C344 VDD1.n113 B 0.011402f
C345 VDD1.n114 B 0.020041f
C346 VDD1.n115 B 0.010769f
C347 VDD1.n116 B 0.025454f
C348 VDD1.n117 B 0.011402f
C349 VDD1.n118 B 0.020041f
C350 VDD1.n119 B 0.010769f
C351 VDD1.n120 B 0.025454f
C352 VDD1.n121 B 0.011402f
C353 VDD1.n122 B 0.020041f
C354 VDD1.n123 B 0.010769f
C355 VDD1.n124 B 0.025454f
C356 VDD1.n125 B 0.011402f
C357 VDD1.n126 B 0.020041f
C358 VDD1.n127 B 0.010769f
C359 VDD1.n128 B 0.025454f
C360 VDD1.n129 B 0.011402f
C361 VDD1.n130 B 0.020041f
C362 VDD1.n131 B 0.010769f
C363 VDD1.n132 B 0.025454f
C364 VDD1.n133 B 0.011402f
C365 VDD1.n134 B 0.020041f
C366 VDD1.n135 B 0.010769f
C367 VDD1.n136 B 0.025454f
C368 VDD1.n137 B 0.011402f
C369 VDD1.n138 B 0.20212f
C370 VDD1.t0 B 0.043799f
C371 VDD1.n139 B 0.019091f
C372 VDD1.n140 B 0.017994f
C373 VDD1.n141 B 0.010769f
C374 VDD1.n142 B 1.67867f
C375 VDD1.n143 B 0.020041f
C376 VDD1.n144 B 0.010769f
C377 VDD1.n145 B 0.011402f
C378 VDD1.n146 B 0.025454f
C379 VDD1.n147 B 0.025454f
C380 VDD1.n148 B 0.011402f
C381 VDD1.n149 B 0.010769f
C382 VDD1.n150 B 0.020041f
C383 VDD1.n151 B 0.020041f
C384 VDD1.n152 B 0.010769f
C385 VDD1.n153 B 0.011402f
C386 VDD1.n154 B 0.025454f
C387 VDD1.n155 B 0.025454f
C388 VDD1.n156 B 0.025454f
C389 VDD1.n157 B 0.011402f
C390 VDD1.n158 B 0.010769f
C391 VDD1.n159 B 0.020041f
C392 VDD1.n160 B 0.020041f
C393 VDD1.n161 B 0.010769f
C394 VDD1.n162 B 0.011086f
C395 VDD1.n163 B 0.011086f
C396 VDD1.n164 B 0.025454f
C397 VDD1.n165 B 0.025454f
C398 VDD1.n166 B 0.011402f
C399 VDD1.n167 B 0.010769f
C400 VDD1.n168 B 0.020041f
C401 VDD1.n169 B 0.020041f
C402 VDD1.n170 B 0.010769f
C403 VDD1.n171 B 0.011402f
C404 VDD1.n172 B 0.025454f
C405 VDD1.n173 B 0.025454f
C406 VDD1.n174 B 0.011402f
C407 VDD1.n175 B 0.010769f
C408 VDD1.n176 B 0.020041f
C409 VDD1.n177 B 0.020041f
C410 VDD1.n178 B 0.010769f
C411 VDD1.n179 B 0.011402f
C412 VDD1.n180 B 0.025454f
C413 VDD1.n181 B 0.025454f
C414 VDD1.n182 B 0.011402f
C415 VDD1.n183 B 0.010769f
C416 VDD1.n184 B 0.020041f
C417 VDD1.n185 B 0.020041f
C418 VDD1.n186 B 0.010769f
C419 VDD1.n187 B 0.011402f
C420 VDD1.n188 B 0.025454f
C421 VDD1.n189 B 0.025454f
C422 VDD1.n190 B 0.011402f
C423 VDD1.n191 B 0.010769f
C424 VDD1.n192 B 0.020041f
C425 VDD1.n193 B 0.020041f
C426 VDD1.n194 B 0.010769f
C427 VDD1.n195 B 0.011402f
C428 VDD1.n196 B 0.025454f
C429 VDD1.n197 B 0.025454f
C430 VDD1.n198 B 0.011402f
C431 VDD1.n199 B 0.010769f
C432 VDD1.n200 B 0.020041f
C433 VDD1.n201 B 0.020041f
C434 VDD1.n202 B 0.010769f
C435 VDD1.n203 B 0.011402f
C436 VDD1.n204 B 0.025454f
C437 VDD1.n205 B 0.05233f
C438 VDD1.n206 B 0.011402f
C439 VDD1.n207 B 0.021057f
C440 VDD1.n208 B 0.050977f
C441 VDD1.n209 B 0.876897f
C442 VTAIL.n0 B 0.027144f
C443 VTAIL.n1 B 0.019681f
C444 VTAIL.n2 B 0.010576f
C445 VTAIL.n3 B 0.024997f
C446 VTAIL.n4 B 0.011198f
C447 VTAIL.n5 B 0.019681f
C448 VTAIL.n6 B 0.010576f
C449 VTAIL.n7 B 0.024997f
C450 VTAIL.n8 B 0.011198f
C451 VTAIL.n9 B 0.019681f
C452 VTAIL.n10 B 0.010576f
C453 VTAIL.n11 B 0.024997f
C454 VTAIL.n12 B 0.011198f
C455 VTAIL.n13 B 0.019681f
C456 VTAIL.n14 B 0.010576f
C457 VTAIL.n15 B 0.024997f
C458 VTAIL.n16 B 0.011198f
C459 VTAIL.n17 B 0.019681f
C460 VTAIL.n18 B 0.010576f
C461 VTAIL.n19 B 0.024997f
C462 VTAIL.n20 B 0.011198f
C463 VTAIL.n21 B 0.019681f
C464 VTAIL.n22 B 0.010576f
C465 VTAIL.n23 B 0.024997f
C466 VTAIL.n24 B 0.011198f
C467 VTAIL.n25 B 0.019681f
C468 VTAIL.n26 B 0.010576f
C469 VTAIL.n27 B 0.024997f
C470 VTAIL.n28 B 0.011198f
C471 VTAIL.n29 B 0.019681f
C472 VTAIL.n30 B 0.010576f
C473 VTAIL.n31 B 0.024997f
C474 VTAIL.n32 B 0.011198f
C475 VTAIL.n33 B 0.19849f
C476 VTAIL.t3 B 0.043012f
C477 VTAIL.n34 B 0.018748f
C478 VTAIL.n35 B 0.017671f
C479 VTAIL.n36 B 0.010576f
C480 VTAIL.n37 B 1.64852f
C481 VTAIL.n38 B 0.019681f
C482 VTAIL.n39 B 0.010576f
C483 VTAIL.n40 B 0.011198f
C484 VTAIL.n41 B 0.024997f
C485 VTAIL.n42 B 0.024997f
C486 VTAIL.n43 B 0.011198f
C487 VTAIL.n44 B 0.010576f
C488 VTAIL.n45 B 0.019681f
C489 VTAIL.n46 B 0.019681f
C490 VTAIL.n47 B 0.010576f
C491 VTAIL.n48 B 0.011198f
C492 VTAIL.n49 B 0.024997f
C493 VTAIL.n50 B 0.024997f
C494 VTAIL.n51 B 0.024997f
C495 VTAIL.n52 B 0.011198f
C496 VTAIL.n53 B 0.010576f
C497 VTAIL.n54 B 0.019681f
C498 VTAIL.n55 B 0.019681f
C499 VTAIL.n56 B 0.010576f
C500 VTAIL.n57 B 0.010887f
C501 VTAIL.n58 B 0.010887f
C502 VTAIL.n59 B 0.024997f
C503 VTAIL.n60 B 0.024997f
C504 VTAIL.n61 B 0.011198f
C505 VTAIL.n62 B 0.010576f
C506 VTAIL.n63 B 0.019681f
C507 VTAIL.n64 B 0.019681f
C508 VTAIL.n65 B 0.010576f
C509 VTAIL.n66 B 0.011198f
C510 VTAIL.n67 B 0.024997f
C511 VTAIL.n68 B 0.024997f
C512 VTAIL.n69 B 0.011198f
C513 VTAIL.n70 B 0.010576f
C514 VTAIL.n71 B 0.019681f
C515 VTAIL.n72 B 0.019681f
C516 VTAIL.n73 B 0.010576f
C517 VTAIL.n74 B 0.011198f
C518 VTAIL.n75 B 0.024997f
C519 VTAIL.n76 B 0.024997f
C520 VTAIL.n77 B 0.011198f
C521 VTAIL.n78 B 0.010576f
C522 VTAIL.n79 B 0.019681f
C523 VTAIL.n80 B 0.019681f
C524 VTAIL.n81 B 0.010576f
C525 VTAIL.n82 B 0.011198f
C526 VTAIL.n83 B 0.024997f
C527 VTAIL.n84 B 0.024997f
C528 VTAIL.n85 B 0.011198f
C529 VTAIL.n86 B 0.010576f
C530 VTAIL.n87 B 0.019681f
C531 VTAIL.n88 B 0.019681f
C532 VTAIL.n89 B 0.010576f
C533 VTAIL.n90 B 0.011198f
C534 VTAIL.n91 B 0.024997f
C535 VTAIL.n92 B 0.024997f
C536 VTAIL.n93 B 0.011198f
C537 VTAIL.n94 B 0.010576f
C538 VTAIL.n95 B 0.019681f
C539 VTAIL.n96 B 0.019681f
C540 VTAIL.n97 B 0.010576f
C541 VTAIL.n98 B 0.011198f
C542 VTAIL.n99 B 0.024997f
C543 VTAIL.n100 B 0.05139f
C544 VTAIL.n101 B 0.011198f
C545 VTAIL.n102 B 0.020679f
C546 VTAIL.n103 B 0.050062f
C547 VTAIL.n104 B 0.053372f
C548 VTAIL.n105 B 1.78303f
C549 VTAIL.n106 B 0.027144f
C550 VTAIL.n107 B 0.019681f
C551 VTAIL.n108 B 0.010576f
C552 VTAIL.n109 B 0.024997f
C553 VTAIL.n110 B 0.011198f
C554 VTAIL.n111 B 0.019681f
C555 VTAIL.n112 B 0.010576f
C556 VTAIL.n113 B 0.024997f
C557 VTAIL.n114 B 0.011198f
C558 VTAIL.n115 B 0.019681f
C559 VTAIL.n116 B 0.010576f
C560 VTAIL.n117 B 0.024997f
C561 VTAIL.n118 B 0.011198f
C562 VTAIL.n119 B 0.019681f
C563 VTAIL.n120 B 0.010576f
C564 VTAIL.n121 B 0.024997f
C565 VTAIL.n122 B 0.011198f
C566 VTAIL.n123 B 0.019681f
C567 VTAIL.n124 B 0.010576f
C568 VTAIL.n125 B 0.024997f
C569 VTAIL.n126 B 0.011198f
C570 VTAIL.n127 B 0.019681f
C571 VTAIL.n128 B 0.010576f
C572 VTAIL.n129 B 0.024997f
C573 VTAIL.n130 B 0.011198f
C574 VTAIL.n131 B 0.019681f
C575 VTAIL.n132 B 0.010576f
C576 VTAIL.n133 B 0.024997f
C577 VTAIL.n134 B 0.024997f
C578 VTAIL.n135 B 0.011198f
C579 VTAIL.n136 B 0.019681f
C580 VTAIL.n137 B 0.010576f
C581 VTAIL.n138 B 0.024997f
C582 VTAIL.n139 B 0.011198f
C583 VTAIL.n140 B 0.19849f
C584 VTAIL.t1 B 0.043012f
C585 VTAIL.n141 B 0.018748f
C586 VTAIL.n142 B 0.017671f
C587 VTAIL.n143 B 0.010576f
C588 VTAIL.n144 B 1.64852f
C589 VTAIL.n145 B 0.019681f
C590 VTAIL.n146 B 0.010576f
C591 VTAIL.n147 B 0.011198f
C592 VTAIL.n148 B 0.024997f
C593 VTAIL.n149 B 0.024997f
C594 VTAIL.n150 B 0.011198f
C595 VTAIL.n151 B 0.010576f
C596 VTAIL.n152 B 0.019681f
C597 VTAIL.n153 B 0.019681f
C598 VTAIL.n154 B 0.010576f
C599 VTAIL.n155 B 0.011198f
C600 VTAIL.n156 B 0.024997f
C601 VTAIL.n157 B 0.024997f
C602 VTAIL.n158 B 0.011198f
C603 VTAIL.n159 B 0.010576f
C604 VTAIL.n160 B 0.019681f
C605 VTAIL.n161 B 0.019681f
C606 VTAIL.n162 B 0.010576f
C607 VTAIL.n163 B 0.010887f
C608 VTAIL.n164 B 0.010887f
C609 VTAIL.n165 B 0.024997f
C610 VTAIL.n166 B 0.024997f
C611 VTAIL.n167 B 0.011198f
C612 VTAIL.n168 B 0.010576f
C613 VTAIL.n169 B 0.019681f
C614 VTAIL.n170 B 0.019681f
C615 VTAIL.n171 B 0.010576f
C616 VTAIL.n172 B 0.011198f
C617 VTAIL.n173 B 0.024997f
C618 VTAIL.n174 B 0.024997f
C619 VTAIL.n175 B 0.011198f
C620 VTAIL.n176 B 0.010576f
C621 VTAIL.n177 B 0.019681f
C622 VTAIL.n178 B 0.019681f
C623 VTAIL.n179 B 0.010576f
C624 VTAIL.n180 B 0.011198f
C625 VTAIL.n181 B 0.024997f
C626 VTAIL.n182 B 0.024997f
C627 VTAIL.n183 B 0.011198f
C628 VTAIL.n184 B 0.010576f
C629 VTAIL.n185 B 0.019681f
C630 VTAIL.n186 B 0.019681f
C631 VTAIL.n187 B 0.010576f
C632 VTAIL.n188 B 0.011198f
C633 VTAIL.n189 B 0.024997f
C634 VTAIL.n190 B 0.024997f
C635 VTAIL.n191 B 0.011198f
C636 VTAIL.n192 B 0.010576f
C637 VTAIL.n193 B 0.019681f
C638 VTAIL.n194 B 0.019681f
C639 VTAIL.n195 B 0.010576f
C640 VTAIL.n196 B 0.011198f
C641 VTAIL.n197 B 0.024997f
C642 VTAIL.n198 B 0.024997f
C643 VTAIL.n199 B 0.011198f
C644 VTAIL.n200 B 0.010576f
C645 VTAIL.n201 B 0.019681f
C646 VTAIL.n202 B 0.019681f
C647 VTAIL.n203 B 0.010576f
C648 VTAIL.n204 B 0.011198f
C649 VTAIL.n205 B 0.024997f
C650 VTAIL.n206 B 0.05139f
C651 VTAIL.n207 B 0.011198f
C652 VTAIL.n208 B 0.020679f
C653 VTAIL.n209 B 0.050062f
C654 VTAIL.n210 B 0.053372f
C655 VTAIL.n211 B 1.82348f
C656 VTAIL.n212 B 0.027144f
C657 VTAIL.n213 B 0.019681f
C658 VTAIL.n214 B 0.010576f
C659 VTAIL.n215 B 0.024997f
C660 VTAIL.n216 B 0.011198f
C661 VTAIL.n217 B 0.019681f
C662 VTAIL.n218 B 0.010576f
C663 VTAIL.n219 B 0.024997f
C664 VTAIL.n220 B 0.011198f
C665 VTAIL.n221 B 0.019681f
C666 VTAIL.n222 B 0.010576f
C667 VTAIL.n223 B 0.024997f
C668 VTAIL.n224 B 0.011198f
C669 VTAIL.n225 B 0.019681f
C670 VTAIL.n226 B 0.010576f
C671 VTAIL.n227 B 0.024997f
C672 VTAIL.n228 B 0.011198f
C673 VTAIL.n229 B 0.019681f
C674 VTAIL.n230 B 0.010576f
C675 VTAIL.n231 B 0.024997f
C676 VTAIL.n232 B 0.011198f
C677 VTAIL.n233 B 0.019681f
C678 VTAIL.n234 B 0.010576f
C679 VTAIL.n235 B 0.024997f
C680 VTAIL.n236 B 0.011198f
C681 VTAIL.n237 B 0.019681f
C682 VTAIL.n238 B 0.010576f
C683 VTAIL.n239 B 0.024997f
C684 VTAIL.n240 B 0.024997f
C685 VTAIL.n241 B 0.011198f
C686 VTAIL.n242 B 0.019681f
C687 VTAIL.n243 B 0.010576f
C688 VTAIL.n244 B 0.024997f
C689 VTAIL.n245 B 0.011198f
C690 VTAIL.n246 B 0.19849f
C691 VTAIL.t2 B 0.043012f
C692 VTAIL.n247 B 0.018748f
C693 VTAIL.n248 B 0.017671f
C694 VTAIL.n249 B 0.010576f
C695 VTAIL.n250 B 1.64852f
C696 VTAIL.n251 B 0.019681f
C697 VTAIL.n252 B 0.010576f
C698 VTAIL.n253 B 0.011198f
C699 VTAIL.n254 B 0.024997f
C700 VTAIL.n255 B 0.024997f
C701 VTAIL.n256 B 0.011198f
C702 VTAIL.n257 B 0.010576f
C703 VTAIL.n258 B 0.019681f
C704 VTAIL.n259 B 0.019681f
C705 VTAIL.n260 B 0.010576f
C706 VTAIL.n261 B 0.011198f
C707 VTAIL.n262 B 0.024997f
C708 VTAIL.n263 B 0.024997f
C709 VTAIL.n264 B 0.011198f
C710 VTAIL.n265 B 0.010576f
C711 VTAIL.n266 B 0.019681f
C712 VTAIL.n267 B 0.019681f
C713 VTAIL.n268 B 0.010576f
C714 VTAIL.n269 B 0.010887f
C715 VTAIL.n270 B 0.010887f
C716 VTAIL.n271 B 0.024997f
C717 VTAIL.n272 B 0.024997f
C718 VTAIL.n273 B 0.011198f
C719 VTAIL.n274 B 0.010576f
C720 VTAIL.n275 B 0.019681f
C721 VTAIL.n276 B 0.019681f
C722 VTAIL.n277 B 0.010576f
C723 VTAIL.n278 B 0.011198f
C724 VTAIL.n279 B 0.024997f
C725 VTAIL.n280 B 0.024997f
C726 VTAIL.n281 B 0.011198f
C727 VTAIL.n282 B 0.010576f
C728 VTAIL.n283 B 0.019681f
C729 VTAIL.n284 B 0.019681f
C730 VTAIL.n285 B 0.010576f
C731 VTAIL.n286 B 0.011198f
C732 VTAIL.n287 B 0.024997f
C733 VTAIL.n288 B 0.024997f
C734 VTAIL.n289 B 0.011198f
C735 VTAIL.n290 B 0.010576f
C736 VTAIL.n291 B 0.019681f
C737 VTAIL.n292 B 0.019681f
C738 VTAIL.n293 B 0.010576f
C739 VTAIL.n294 B 0.011198f
C740 VTAIL.n295 B 0.024997f
C741 VTAIL.n296 B 0.024997f
C742 VTAIL.n297 B 0.011198f
C743 VTAIL.n298 B 0.010576f
C744 VTAIL.n299 B 0.019681f
C745 VTAIL.n300 B 0.019681f
C746 VTAIL.n301 B 0.010576f
C747 VTAIL.n302 B 0.011198f
C748 VTAIL.n303 B 0.024997f
C749 VTAIL.n304 B 0.024997f
C750 VTAIL.n305 B 0.011198f
C751 VTAIL.n306 B 0.010576f
C752 VTAIL.n307 B 0.019681f
C753 VTAIL.n308 B 0.019681f
C754 VTAIL.n309 B 0.010576f
C755 VTAIL.n310 B 0.011198f
C756 VTAIL.n311 B 0.024997f
C757 VTAIL.n312 B 0.05139f
C758 VTAIL.n313 B 0.011198f
C759 VTAIL.n314 B 0.020679f
C760 VTAIL.n315 B 0.050062f
C761 VTAIL.n316 B 0.053372f
C762 VTAIL.n317 B 1.6469f
C763 VTAIL.n318 B 0.027144f
C764 VTAIL.n319 B 0.019681f
C765 VTAIL.n320 B 0.010576f
C766 VTAIL.n321 B 0.024997f
C767 VTAIL.n322 B 0.011198f
C768 VTAIL.n323 B 0.019681f
C769 VTAIL.n324 B 0.010576f
C770 VTAIL.n325 B 0.024997f
C771 VTAIL.n326 B 0.011198f
C772 VTAIL.n327 B 0.019681f
C773 VTAIL.n328 B 0.010576f
C774 VTAIL.n329 B 0.024997f
C775 VTAIL.n330 B 0.011198f
C776 VTAIL.n331 B 0.019681f
C777 VTAIL.n332 B 0.010576f
C778 VTAIL.n333 B 0.024997f
C779 VTAIL.n334 B 0.011198f
C780 VTAIL.n335 B 0.019681f
C781 VTAIL.n336 B 0.010576f
C782 VTAIL.n337 B 0.024997f
C783 VTAIL.n338 B 0.011198f
C784 VTAIL.n339 B 0.019681f
C785 VTAIL.n340 B 0.010576f
C786 VTAIL.n341 B 0.024997f
C787 VTAIL.n342 B 0.011198f
C788 VTAIL.n343 B 0.019681f
C789 VTAIL.n344 B 0.010576f
C790 VTAIL.n345 B 0.024997f
C791 VTAIL.n346 B 0.011198f
C792 VTAIL.n347 B 0.019681f
C793 VTAIL.n348 B 0.010576f
C794 VTAIL.n349 B 0.024997f
C795 VTAIL.n350 B 0.011198f
C796 VTAIL.n351 B 0.19849f
C797 VTAIL.t0 B 0.043012f
C798 VTAIL.n352 B 0.018748f
C799 VTAIL.n353 B 0.017671f
C800 VTAIL.n354 B 0.010576f
C801 VTAIL.n355 B 1.64852f
C802 VTAIL.n356 B 0.019681f
C803 VTAIL.n357 B 0.010576f
C804 VTAIL.n358 B 0.011198f
C805 VTAIL.n359 B 0.024997f
C806 VTAIL.n360 B 0.024997f
C807 VTAIL.n361 B 0.011198f
C808 VTAIL.n362 B 0.010576f
C809 VTAIL.n363 B 0.019681f
C810 VTAIL.n364 B 0.019681f
C811 VTAIL.n365 B 0.010576f
C812 VTAIL.n366 B 0.011198f
C813 VTAIL.n367 B 0.024997f
C814 VTAIL.n368 B 0.024997f
C815 VTAIL.n369 B 0.024997f
C816 VTAIL.n370 B 0.011198f
C817 VTAIL.n371 B 0.010576f
C818 VTAIL.n372 B 0.019681f
C819 VTAIL.n373 B 0.019681f
C820 VTAIL.n374 B 0.010576f
C821 VTAIL.n375 B 0.010887f
C822 VTAIL.n376 B 0.010887f
C823 VTAIL.n377 B 0.024997f
C824 VTAIL.n378 B 0.024997f
C825 VTAIL.n379 B 0.011198f
C826 VTAIL.n380 B 0.010576f
C827 VTAIL.n381 B 0.019681f
C828 VTAIL.n382 B 0.019681f
C829 VTAIL.n383 B 0.010576f
C830 VTAIL.n384 B 0.011198f
C831 VTAIL.n385 B 0.024997f
C832 VTAIL.n386 B 0.024997f
C833 VTAIL.n387 B 0.011198f
C834 VTAIL.n388 B 0.010576f
C835 VTAIL.n389 B 0.019681f
C836 VTAIL.n390 B 0.019681f
C837 VTAIL.n391 B 0.010576f
C838 VTAIL.n392 B 0.011198f
C839 VTAIL.n393 B 0.024997f
C840 VTAIL.n394 B 0.024997f
C841 VTAIL.n395 B 0.011198f
C842 VTAIL.n396 B 0.010576f
C843 VTAIL.n397 B 0.019681f
C844 VTAIL.n398 B 0.019681f
C845 VTAIL.n399 B 0.010576f
C846 VTAIL.n400 B 0.011198f
C847 VTAIL.n401 B 0.024997f
C848 VTAIL.n402 B 0.024997f
C849 VTAIL.n403 B 0.011198f
C850 VTAIL.n404 B 0.010576f
C851 VTAIL.n405 B 0.019681f
C852 VTAIL.n406 B 0.019681f
C853 VTAIL.n407 B 0.010576f
C854 VTAIL.n408 B 0.011198f
C855 VTAIL.n409 B 0.024997f
C856 VTAIL.n410 B 0.024997f
C857 VTAIL.n411 B 0.011198f
C858 VTAIL.n412 B 0.010576f
C859 VTAIL.n413 B 0.019681f
C860 VTAIL.n414 B 0.019681f
C861 VTAIL.n415 B 0.010576f
C862 VTAIL.n416 B 0.011198f
C863 VTAIL.n417 B 0.024997f
C864 VTAIL.n418 B 0.05139f
C865 VTAIL.n419 B 0.011198f
C866 VTAIL.n420 B 0.020679f
C867 VTAIL.n421 B 0.050062f
C868 VTAIL.n422 B 0.053372f
C869 VTAIL.n423 B 1.56927f
C870 VP.t1 B 4.64045f
C871 VP.t0 B 5.25388f
C872 VP.n0 B 5.42624f
.ends

