* NGSPICE file created from diff_pair_sample_1116.ext - technology: sky130A

.subckt diff_pair_sample_1116 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=5.9631 ps=31.36 w=15.29 l=2.07
X1 VDD2.t9 VN.t0 VTAIL.t5 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=2.52285 ps=15.62 w=15.29 l=2.07
X2 B.t11 B.t9 B.t10 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=0 ps=0 w=15.29 l=2.07
X3 VDD1.t8 VP.t1 VTAIL.t11 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=5.9631 ps=31.36 w=15.29 l=2.07
X4 VTAIL.t12 VP.t2 VDD1.t7 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X5 VDD2.t8 VN.t1 VTAIL.t8 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=5.9631 ps=31.36 w=15.29 l=2.07
X6 VTAIL.t16 VP.t3 VDD1.t6 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X7 VTAIL.t1 VN.t2 VDD2.t7 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X8 VTAIL.t2 VN.t3 VDD2.t6 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X9 B.t8 B.t6 B.t7 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=0 ps=0 w=15.29 l=2.07
X10 VDD2.t5 VN.t4 VTAIL.t4 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=5.9631 ps=31.36 w=15.29 l=2.07
X11 VTAIL.t9 VN.t5 VDD2.t4 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X12 VTAIL.t13 VP.t4 VDD1.t5 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X13 VDD1.t4 VP.t5 VTAIL.t17 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X14 VDD2.t3 VN.t6 VTAIL.t7 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X15 B.t5 B.t3 B.t4 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=0 ps=0 w=15.29 l=2.07
X16 VDD1.t3 VP.t6 VTAIL.t18 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=2.52285 ps=15.62 w=15.29 l=2.07
X17 B.t2 B.t0 B.t1 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=0 ps=0 w=15.29 l=2.07
X18 VTAIL.t0 VN.t7 VDD2.t2 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X19 VDD2.t1 VN.t8 VTAIL.t3 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=2.52285 ps=15.62 w=15.29 l=2.07
X20 VDD1.t2 VP.t7 VTAIL.t19 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=5.9631 pd=31.36 as=2.52285 ps=15.62 w=15.29 l=2.07
X21 VDD2.t0 VN.t9 VTAIL.t6 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X22 VTAIL.t15 VP.t8 VDD1.t1 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
X23 VDD1.t0 VP.t9 VTAIL.t14 w_n3850_n4026# sky130_fd_pr__pfet_01v8 ad=2.52285 pd=15.62 as=2.52285 ps=15.62 w=15.29 l=2.07
R0 VP.n18 VP.t6 210.953
R1 VP.n60 VP.t9 178.014
R2 VP.n44 VP.t7 178.014
R3 VP.n7 VP.t8 178.014
R4 VP.n67 VP.t2 178.014
R5 VP.n75 VP.t1 178.014
R6 VP.n26 VP.t5 178.014
R7 VP.n41 VP.t0 178.014
R8 VP.n33 VP.t3 178.014
R9 VP.n17 VP.t4 178.014
R10 VP.n20 VP.n19 161.3
R11 VP.n21 VP.n16 161.3
R12 VP.n23 VP.n22 161.3
R13 VP.n24 VP.n15 161.3
R14 VP.n26 VP.n25 161.3
R15 VP.n27 VP.n14 161.3
R16 VP.n29 VP.n28 161.3
R17 VP.n30 VP.n13 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n34 VP.n12 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n37 VP.n11 161.3
R22 VP.n39 VP.n38 161.3
R23 VP.n40 VP.n10 161.3
R24 VP.n74 VP.n0 161.3
R25 VP.n73 VP.n72 161.3
R26 VP.n71 VP.n1 161.3
R27 VP.n70 VP.n69 161.3
R28 VP.n68 VP.n2 161.3
R29 VP.n66 VP.n65 161.3
R30 VP.n64 VP.n3 161.3
R31 VP.n63 VP.n62 161.3
R32 VP.n61 VP.n4 161.3
R33 VP.n60 VP.n59 161.3
R34 VP.n58 VP.n5 161.3
R35 VP.n57 VP.n56 161.3
R36 VP.n55 VP.n6 161.3
R37 VP.n54 VP.n53 161.3
R38 VP.n52 VP.n51 161.3
R39 VP.n50 VP.n8 161.3
R40 VP.n49 VP.n48 161.3
R41 VP.n47 VP.n9 161.3
R42 VP.n46 VP.n45 161.3
R43 VP.n44 VP.n43 96.0763
R44 VP.n76 VP.n75 96.0763
R45 VP.n42 VP.n41 96.0763
R46 VP.n56 VP.n55 56.5193
R47 VP.n62 VP.n3 56.5193
R48 VP.n28 VP.n13 56.5193
R49 VP.n22 VP.n21 56.5193
R50 VP.n43 VP.n42 52.689
R51 VP.n18 VP.n17 51.1767
R52 VP.n49 VP.n9 50.2061
R53 VP.n73 VP.n1 50.2061
R54 VP.n39 VP.n11 50.2061
R55 VP.n50 VP.n49 30.7807
R56 VP.n69 VP.n1 30.7807
R57 VP.n35 VP.n11 30.7807
R58 VP.n45 VP.n9 24.4675
R59 VP.n51 VP.n50 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n5 24.4675
R62 VP.n60 VP.n5 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n62 VP.n61 24.4675
R65 VP.n66 VP.n3 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n74 VP.n73 24.4675
R68 VP.n40 VP.n39 24.4675
R69 VP.n32 VP.n13 24.4675
R70 VP.n35 VP.n34 24.4675
R71 VP.n22 VP.n15 24.4675
R72 VP.n26 VP.n15 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 19.5741
R77 VP.n67 VP.n66 19.5741
R78 VP.n33 VP.n32 19.5741
R79 VP.n20 VP.n17 19.5741
R80 VP.n45 VP.n44 14.6807
R81 VP.n75 VP.n74 14.6807
R82 VP.n41 VP.n40 14.6807
R83 VP.n19 VP.n18 9.46762
R84 VP.n51 VP.n7 4.8939
R85 VP.n68 VP.n67 4.8939
R86 VP.n34 VP.n33 4.8939
R87 VP.n42 VP.n10 0.278367
R88 VP.n46 VP.n43 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153454
R122 VTAIL.n16 VTAIL.t10 54.8796
R123 VTAIL.n11 VTAIL.t4 54.8796
R124 VTAIL.n17 VTAIL.t8 54.8794
R125 VTAIL.n2 VTAIL.t11 54.8794
R126 VTAIL.n15 VTAIL.n14 52.7538
R127 VTAIL.n13 VTAIL.n12 52.7538
R128 VTAIL.n10 VTAIL.n9 52.7538
R129 VTAIL.n8 VTAIL.n7 52.7538
R130 VTAIL.n19 VTAIL.n18 52.7535
R131 VTAIL.n1 VTAIL.n0 52.7535
R132 VTAIL.n4 VTAIL.n3 52.7535
R133 VTAIL.n6 VTAIL.n5 52.7535
R134 VTAIL.n8 VTAIL.n6 29.6858
R135 VTAIL.n17 VTAIL.n16 27.6169
R136 VTAIL.n18 VTAIL.t6 2.1264
R137 VTAIL.n18 VTAIL.t2 2.1264
R138 VTAIL.n0 VTAIL.t3 2.1264
R139 VTAIL.n0 VTAIL.t0 2.1264
R140 VTAIL.n3 VTAIL.t14 2.1264
R141 VTAIL.n3 VTAIL.t12 2.1264
R142 VTAIL.n5 VTAIL.t19 2.1264
R143 VTAIL.n5 VTAIL.t15 2.1264
R144 VTAIL.n14 VTAIL.t17 2.1264
R145 VTAIL.n14 VTAIL.t16 2.1264
R146 VTAIL.n12 VTAIL.t18 2.1264
R147 VTAIL.n12 VTAIL.t13 2.1264
R148 VTAIL.n9 VTAIL.t7 2.1264
R149 VTAIL.n9 VTAIL.t9 2.1264
R150 VTAIL.n7 VTAIL.t5 2.1264
R151 VTAIL.n7 VTAIL.t1 2.1264
R152 VTAIL.n10 VTAIL.n8 2.06947
R153 VTAIL.n11 VTAIL.n10 2.06947
R154 VTAIL.n15 VTAIL.n13 2.06947
R155 VTAIL.n16 VTAIL.n15 2.06947
R156 VTAIL.n6 VTAIL.n4 2.06947
R157 VTAIL.n4 VTAIL.n2 2.06947
R158 VTAIL.n19 VTAIL.n17 2.06947
R159 VTAIL VTAIL.n1 1.61041
R160 VTAIL.n13 VTAIL.n11 1.50481
R161 VTAIL.n2 VTAIL.n1 1.50481
R162 VTAIL VTAIL.n19 0.459552
R163 VDD1.n1 VDD1.t3 73.6274
R164 VDD1.n3 VDD1.t2 73.6272
R165 VDD1.n5 VDD1.n4 70.9287
R166 VDD1.n7 VDD1.n6 69.4325
R167 VDD1.n1 VDD1.n0 69.4325
R168 VDD1.n3 VDD1.n2 69.4323
R169 VDD1.n7 VDD1.n5 48.3414
R170 VDD1.n6 VDD1.t6 2.1264
R171 VDD1.n6 VDD1.t9 2.1264
R172 VDD1.n0 VDD1.t5 2.1264
R173 VDD1.n0 VDD1.t4 2.1264
R174 VDD1.n4 VDD1.t7 2.1264
R175 VDD1.n4 VDD1.t8 2.1264
R176 VDD1.n2 VDD1.t1 2.1264
R177 VDD1.n2 VDD1.t0 2.1264
R178 VDD1 VDD1.n7 1.49403
R179 VDD1 VDD1.n1 0.575931
R180 VDD1.n5 VDD1.n3 0.462395
R181 VN.n8 VN.t8 210.953
R182 VN.n41 VN.t4 210.953
R183 VN.n16 VN.t9 178.014
R184 VN.n7 VN.t7 178.014
R185 VN.n23 VN.t3 178.014
R186 VN.n31 VN.t1 178.014
R187 VN.n49 VN.t6 178.014
R188 VN.n40 VN.t5 178.014
R189 VN.n56 VN.t2 178.014
R190 VN.n64 VN.t0 178.014
R191 VN.n63 VN.n33 161.3
R192 VN.n62 VN.n61 161.3
R193 VN.n60 VN.n34 161.3
R194 VN.n59 VN.n58 161.3
R195 VN.n57 VN.n35 161.3
R196 VN.n55 VN.n54 161.3
R197 VN.n53 VN.n36 161.3
R198 VN.n52 VN.n51 161.3
R199 VN.n50 VN.n37 161.3
R200 VN.n49 VN.n48 161.3
R201 VN.n47 VN.n38 161.3
R202 VN.n46 VN.n45 161.3
R203 VN.n44 VN.n39 161.3
R204 VN.n43 VN.n42 161.3
R205 VN.n30 VN.n0 161.3
R206 VN.n29 VN.n28 161.3
R207 VN.n27 VN.n1 161.3
R208 VN.n26 VN.n25 161.3
R209 VN.n24 VN.n2 161.3
R210 VN.n22 VN.n21 161.3
R211 VN.n20 VN.n3 161.3
R212 VN.n19 VN.n18 161.3
R213 VN.n17 VN.n4 161.3
R214 VN.n16 VN.n15 161.3
R215 VN.n14 VN.n5 161.3
R216 VN.n13 VN.n12 161.3
R217 VN.n11 VN.n6 161.3
R218 VN.n10 VN.n9 161.3
R219 VN.n32 VN.n31 96.0763
R220 VN.n65 VN.n64 96.0763
R221 VN.n12 VN.n11 56.5193
R222 VN.n18 VN.n3 56.5193
R223 VN.n45 VN.n44 56.5193
R224 VN.n51 VN.n36 56.5193
R225 VN VN.n65 52.9678
R226 VN.n8 VN.n7 51.1767
R227 VN.n41 VN.n40 51.1767
R228 VN.n29 VN.n1 50.2061
R229 VN.n62 VN.n34 50.2061
R230 VN.n25 VN.n1 30.7807
R231 VN.n58 VN.n34 30.7807
R232 VN.n11 VN.n10 24.4675
R233 VN.n12 VN.n5 24.4675
R234 VN.n16 VN.n5 24.4675
R235 VN.n17 VN.n16 24.4675
R236 VN.n18 VN.n17 24.4675
R237 VN.n22 VN.n3 24.4675
R238 VN.n25 VN.n24 24.4675
R239 VN.n30 VN.n29 24.4675
R240 VN.n44 VN.n43 24.4675
R241 VN.n51 VN.n50 24.4675
R242 VN.n50 VN.n49 24.4675
R243 VN.n49 VN.n38 24.4675
R244 VN.n45 VN.n38 24.4675
R245 VN.n58 VN.n57 24.4675
R246 VN.n55 VN.n36 24.4675
R247 VN.n63 VN.n62 24.4675
R248 VN.n10 VN.n7 19.5741
R249 VN.n23 VN.n22 19.5741
R250 VN.n43 VN.n40 19.5741
R251 VN.n56 VN.n55 19.5741
R252 VN.n31 VN.n30 14.6807
R253 VN.n64 VN.n63 14.6807
R254 VN.n42 VN.n41 9.46762
R255 VN.n9 VN.n8 9.46762
R256 VN.n24 VN.n23 4.8939
R257 VN.n57 VN.n56 4.8939
R258 VN.n65 VN.n33 0.278367
R259 VN.n32 VN.n0 0.278367
R260 VN.n61 VN.n33 0.189894
R261 VN.n61 VN.n60 0.189894
R262 VN.n60 VN.n59 0.189894
R263 VN.n59 VN.n35 0.189894
R264 VN.n54 VN.n35 0.189894
R265 VN.n54 VN.n53 0.189894
R266 VN.n53 VN.n52 0.189894
R267 VN.n52 VN.n37 0.189894
R268 VN.n48 VN.n37 0.189894
R269 VN.n48 VN.n47 0.189894
R270 VN.n47 VN.n46 0.189894
R271 VN.n46 VN.n39 0.189894
R272 VN.n42 VN.n39 0.189894
R273 VN.n9 VN.n6 0.189894
R274 VN.n13 VN.n6 0.189894
R275 VN.n14 VN.n13 0.189894
R276 VN.n15 VN.n14 0.189894
R277 VN.n15 VN.n4 0.189894
R278 VN.n19 VN.n4 0.189894
R279 VN.n20 VN.n19 0.189894
R280 VN.n21 VN.n20 0.189894
R281 VN.n21 VN.n2 0.189894
R282 VN.n26 VN.n2 0.189894
R283 VN.n27 VN.n26 0.189894
R284 VN.n28 VN.n27 0.189894
R285 VN.n28 VN.n0 0.189894
R286 VN VN.n32 0.153454
R287 VDD2.n1 VDD2.t1 73.6272
R288 VDD2.n4 VDD2.t9 71.5584
R289 VDD2.n3 VDD2.n2 70.9287
R290 VDD2 VDD2.n7 70.9261
R291 VDD2.n6 VDD2.n5 69.4325
R292 VDD2.n1 VDD2.n0 69.4323
R293 VDD2.n4 VDD2.n3 46.7239
R294 VDD2.n7 VDD2.t4 2.1264
R295 VDD2.n7 VDD2.t5 2.1264
R296 VDD2.n5 VDD2.t7 2.1264
R297 VDD2.n5 VDD2.t3 2.1264
R298 VDD2.n2 VDD2.t6 2.1264
R299 VDD2.n2 VDD2.t8 2.1264
R300 VDD2.n0 VDD2.t2 2.1264
R301 VDD2.n0 VDD2.t0 2.1264
R302 VDD2.n6 VDD2.n4 2.06947
R303 VDD2 VDD2.n6 0.575931
R304 VDD2.n3 VDD2.n1 0.462395
R305 B.n466 B.n139 585
R306 B.n465 B.n464 585
R307 B.n463 B.n140 585
R308 B.n462 B.n461 585
R309 B.n460 B.n141 585
R310 B.n459 B.n458 585
R311 B.n457 B.n142 585
R312 B.n456 B.n455 585
R313 B.n454 B.n143 585
R314 B.n453 B.n452 585
R315 B.n451 B.n144 585
R316 B.n450 B.n449 585
R317 B.n448 B.n145 585
R318 B.n447 B.n446 585
R319 B.n445 B.n146 585
R320 B.n444 B.n443 585
R321 B.n442 B.n147 585
R322 B.n441 B.n440 585
R323 B.n439 B.n148 585
R324 B.n438 B.n437 585
R325 B.n436 B.n149 585
R326 B.n435 B.n434 585
R327 B.n433 B.n150 585
R328 B.n432 B.n431 585
R329 B.n430 B.n151 585
R330 B.n429 B.n428 585
R331 B.n427 B.n152 585
R332 B.n426 B.n425 585
R333 B.n424 B.n153 585
R334 B.n423 B.n422 585
R335 B.n421 B.n154 585
R336 B.n420 B.n419 585
R337 B.n418 B.n155 585
R338 B.n417 B.n416 585
R339 B.n415 B.n156 585
R340 B.n414 B.n413 585
R341 B.n412 B.n157 585
R342 B.n411 B.n410 585
R343 B.n409 B.n158 585
R344 B.n408 B.n407 585
R345 B.n406 B.n159 585
R346 B.n405 B.n404 585
R347 B.n403 B.n160 585
R348 B.n402 B.n401 585
R349 B.n400 B.n161 585
R350 B.n399 B.n398 585
R351 B.n397 B.n162 585
R352 B.n396 B.n395 585
R353 B.n394 B.n163 585
R354 B.n393 B.n392 585
R355 B.n391 B.n164 585
R356 B.n389 B.n388 585
R357 B.n387 B.n167 585
R358 B.n386 B.n385 585
R359 B.n384 B.n168 585
R360 B.n383 B.n382 585
R361 B.n381 B.n169 585
R362 B.n380 B.n379 585
R363 B.n378 B.n170 585
R364 B.n377 B.n376 585
R365 B.n375 B.n171 585
R366 B.n374 B.n373 585
R367 B.n369 B.n172 585
R368 B.n368 B.n367 585
R369 B.n366 B.n173 585
R370 B.n365 B.n364 585
R371 B.n363 B.n174 585
R372 B.n362 B.n361 585
R373 B.n360 B.n175 585
R374 B.n359 B.n358 585
R375 B.n357 B.n176 585
R376 B.n356 B.n355 585
R377 B.n354 B.n177 585
R378 B.n353 B.n352 585
R379 B.n351 B.n178 585
R380 B.n350 B.n349 585
R381 B.n348 B.n179 585
R382 B.n347 B.n346 585
R383 B.n345 B.n180 585
R384 B.n344 B.n343 585
R385 B.n342 B.n181 585
R386 B.n341 B.n340 585
R387 B.n339 B.n182 585
R388 B.n338 B.n337 585
R389 B.n336 B.n183 585
R390 B.n335 B.n334 585
R391 B.n333 B.n184 585
R392 B.n332 B.n331 585
R393 B.n330 B.n185 585
R394 B.n329 B.n328 585
R395 B.n327 B.n186 585
R396 B.n326 B.n325 585
R397 B.n324 B.n187 585
R398 B.n323 B.n322 585
R399 B.n321 B.n188 585
R400 B.n320 B.n319 585
R401 B.n318 B.n189 585
R402 B.n317 B.n316 585
R403 B.n315 B.n190 585
R404 B.n314 B.n313 585
R405 B.n312 B.n191 585
R406 B.n311 B.n310 585
R407 B.n309 B.n192 585
R408 B.n308 B.n307 585
R409 B.n306 B.n193 585
R410 B.n305 B.n304 585
R411 B.n303 B.n194 585
R412 B.n302 B.n301 585
R413 B.n300 B.n195 585
R414 B.n299 B.n298 585
R415 B.n297 B.n196 585
R416 B.n296 B.n295 585
R417 B.n468 B.n467 585
R418 B.n469 B.n138 585
R419 B.n471 B.n470 585
R420 B.n472 B.n137 585
R421 B.n474 B.n473 585
R422 B.n475 B.n136 585
R423 B.n477 B.n476 585
R424 B.n478 B.n135 585
R425 B.n480 B.n479 585
R426 B.n481 B.n134 585
R427 B.n483 B.n482 585
R428 B.n484 B.n133 585
R429 B.n486 B.n485 585
R430 B.n487 B.n132 585
R431 B.n489 B.n488 585
R432 B.n490 B.n131 585
R433 B.n492 B.n491 585
R434 B.n493 B.n130 585
R435 B.n495 B.n494 585
R436 B.n496 B.n129 585
R437 B.n498 B.n497 585
R438 B.n499 B.n128 585
R439 B.n501 B.n500 585
R440 B.n502 B.n127 585
R441 B.n504 B.n503 585
R442 B.n505 B.n126 585
R443 B.n507 B.n506 585
R444 B.n508 B.n125 585
R445 B.n510 B.n509 585
R446 B.n511 B.n124 585
R447 B.n513 B.n512 585
R448 B.n514 B.n123 585
R449 B.n516 B.n515 585
R450 B.n517 B.n122 585
R451 B.n519 B.n518 585
R452 B.n520 B.n121 585
R453 B.n522 B.n521 585
R454 B.n523 B.n120 585
R455 B.n525 B.n524 585
R456 B.n526 B.n119 585
R457 B.n528 B.n527 585
R458 B.n529 B.n118 585
R459 B.n531 B.n530 585
R460 B.n532 B.n117 585
R461 B.n534 B.n533 585
R462 B.n535 B.n116 585
R463 B.n537 B.n536 585
R464 B.n538 B.n115 585
R465 B.n540 B.n539 585
R466 B.n541 B.n114 585
R467 B.n543 B.n542 585
R468 B.n544 B.n113 585
R469 B.n546 B.n545 585
R470 B.n547 B.n112 585
R471 B.n549 B.n548 585
R472 B.n550 B.n111 585
R473 B.n552 B.n551 585
R474 B.n553 B.n110 585
R475 B.n555 B.n554 585
R476 B.n556 B.n109 585
R477 B.n558 B.n557 585
R478 B.n559 B.n108 585
R479 B.n561 B.n560 585
R480 B.n562 B.n107 585
R481 B.n564 B.n563 585
R482 B.n565 B.n106 585
R483 B.n567 B.n566 585
R484 B.n568 B.n105 585
R485 B.n570 B.n569 585
R486 B.n571 B.n104 585
R487 B.n573 B.n572 585
R488 B.n574 B.n103 585
R489 B.n576 B.n575 585
R490 B.n577 B.n102 585
R491 B.n579 B.n578 585
R492 B.n580 B.n101 585
R493 B.n582 B.n581 585
R494 B.n583 B.n100 585
R495 B.n585 B.n584 585
R496 B.n586 B.n99 585
R497 B.n588 B.n587 585
R498 B.n589 B.n98 585
R499 B.n591 B.n590 585
R500 B.n592 B.n97 585
R501 B.n594 B.n593 585
R502 B.n595 B.n96 585
R503 B.n597 B.n596 585
R504 B.n598 B.n95 585
R505 B.n600 B.n599 585
R506 B.n601 B.n94 585
R507 B.n603 B.n602 585
R508 B.n604 B.n93 585
R509 B.n606 B.n605 585
R510 B.n607 B.n92 585
R511 B.n609 B.n608 585
R512 B.n610 B.n91 585
R513 B.n612 B.n611 585
R514 B.n613 B.n90 585
R515 B.n615 B.n614 585
R516 B.n616 B.n89 585
R517 B.n618 B.n617 585
R518 B.n619 B.n88 585
R519 B.n788 B.n27 585
R520 B.n787 B.n786 585
R521 B.n785 B.n28 585
R522 B.n784 B.n783 585
R523 B.n782 B.n29 585
R524 B.n781 B.n780 585
R525 B.n779 B.n30 585
R526 B.n778 B.n777 585
R527 B.n776 B.n31 585
R528 B.n775 B.n774 585
R529 B.n773 B.n32 585
R530 B.n772 B.n771 585
R531 B.n770 B.n33 585
R532 B.n769 B.n768 585
R533 B.n767 B.n34 585
R534 B.n766 B.n765 585
R535 B.n764 B.n35 585
R536 B.n763 B.n762 585
R537 B.n761 B.n36 585
R538 B.n760 B.n759 585
R539 B.n758 B.n37 585
R540 B.n757 B.n756 585
R541 B.n755 B.n38 585
R542 B.n754 B.n753 585
R543 B.n752 B.n39 585
R544 B.n751 B.n750 585
R545 B.n749 B.n40 585
R546 B.n748 B.n747 585
R547 B.n746 B.n41 585
R548 B.n745 B.n744 585
R549 B.n743 B.n42 585
R550 B.n742 B.n741 585
R551 B.n740 B.n43 585
R552 B.n739 B.n738 585
R553 B.n737 B.n44 585
R554 B.n736 B.n735 585
R555 B.n734 B.n45 585
R556 B.n733 B.n732 585
R557 B.n731 B.n46 585
R558 B.n730 B.n729 585
R559 B.n728 B.n47 585
R560 B.n727 B.n726 585
R561 B.n725 B.n48 585
R562 B.n724 B.n723 585
R563 B.n722 B.n49 585
R564 B.n721 B.n720 585
R565 B.n719 B.n50 585
R566 B.n718 B.n717 585
R567 B.n716 B.n51 585
R568 B.n715 B.n714 585
R569 B.n713 B.n52 585
R570 B.n712 B.n711 585
R571 B.n710 B.n53 585
R572 B.n709 B.n708 585
R573 B.n707 B.n57 585
R574 B.n706 B.n705 585
R575 B.n704 B.n58 585
R576 B.n703 B.n702 585
R577 B.n701 B.n59 585
R578 B.n700 B.n699 585
R579 B.n698 B.n60 585
R580 B.n696 B.n695 585
R581 B.n694 B.n63 585
R582 B.n693 B.n692 585
R583 B.n691 B.n64 585
R584 B.n690 B.n689 585
R585 B.n688 B.n65 585
R586 B.n687 B.n686 585
R587 B.n685 B.n66 585
R588 B.n684 B.n683 585
R589 B.n682 B.n67 585
R590 B.n681 B.n680 585
R591 B.n679 B.n68 585
R592 B.n678 B.n677 585
R593 B.n676 B.n69 585
R594 B.n675 B.n674 585
R595 B.n673 B.n70 585
R596 B.n672 B.n671 585
R597 B.n670 B.n71 585
R598 B.n669 B.n668 585
R599 B.n667 B.n72 585
R600 B.n666 B.n665 585
R601 B.n664 B.n73 585
R602 B.n663 B.n662 585
R603 B.n661 B.n74 585
R604 B.n660 B.n659 585
R605 B.n658 B.n75 585
R606 B.n657 B.n656 585
R607 B.n655 B.n76 585
R608 B.n654 B.n653 585
R609 B.n652 B.n77 585
R610 B.n651 B.n650 585
R611 B.n649 B.n78 585
R612 B.n648 B.n647 585
R613 B.n646 B.n79 585
R614 B.n645 B.n644 585
R615 B.n643 B.n80 585
R616 B.n642 B.n641 585
R617 B.n640 B.n81 585
R618 B.n639 B.n638 585
R619 B.n637 B.n82 585
R620 B.n636 B.n635 585
R621 B.n634 B.n83 585
R622 B.n633 B.n632 585
R623 B.n631 B.n84 585
R624 B.n630 B.n629 585
R625 B.n628 B.n85 585
R626 B.n627 B.n626 585
R627 B.n625 B.n86 585
R628 B.n624 B.n623 585
R629 B.n622 B.n87 585
R630 B.n621 B.n620 585
R631 B.n790 B.n789 585
R632 B.n791 B.n26 585
R633 B.n793 B.n792 585
R634 B.n794 B.n25 585
R635 B.n796 B.n795 585
R636 B.n797 B.n24 585
R637 B.n799 B.n798 585
R638 B.n800 B.n23 585
R639 B.n802 B.n801 585
R640 B.n803 B.n22 585
R641 B.n805 B.n804 585
R642 B.n806 B.n21 585
R643 B.n808 B.n807 585
R644 B.n809 B.n20 585
R645 B.n811 B.n810 585
R646 B.n812 B.n19 585
R647 B.n814 B.n813 585
R648 B.n815 B.n18 585
R649 B.n817 B.n816 585
R650 B.n818 B.n17 585
R651 B.n820 B.n819 585
R652 B.n821 B.n16 585
R653 B.n823 B.n822 585
R654 B.n824 B.n15 585
R655 B.n826 B.n825 585
R656 B.n827 B.n14 585
R657 B.n829 B.n828 585
R658 B.n830 B.n13 585
R659 B.n832 B.n831 585
R660 B.n833 B.n12 585
R661 B.n835 B.n834 585
R662 B.n836 B.n11 585
R663 B.n838 B.n837 585
R664 B.n839 B.n10 585
R665 B.n841 B.n840 585
R666 B.n842 B.n9 585
R667 B.n844 B.n843 585
R668 B.n845 B.n8 585
R669 B.n847 B.n846 585
R670 B.n848 B.n7 585
R671 B.n850 B.n849 585
R672 B.n851 B.n6 585
R673 B.n853 B.n852 585
R674 B.n854 B.n5 585
R675 B.n856 B.n855 585
R676 B.n857 B.n4 585
R677 B.n859 B.n858 585
R678 B.n860 B.n3 585
R679 B.n862 B.n861 585
R680 B.n863 B.n0 585
R681 B.n2 B.n1 585
R682 B.n222 B.n221 585
R683 B.n224 B.n223 585
R684 B.n225 B.n220 585
R685 B.n227 B.n226 585
R686 B.n228 B.n219 585
R687 B.n230 B.n229 585
R688 B.n231 B.n218 585
R689 B.n233 B.n232 585
R690 B.n234 B.n217 585
R691 B.n236 B.n235 585
R692 B.n237 B.n216 585
R693 B.n239 B.n238 585
R694 B.n240 B.n215 585
R695 B.n242 B.n241 585
R696 B.n243 B.n214 585
R697 B.n245 B.n244 585
R698 B.n246 B.n213 585
R699 B.n248 B.n247 585
R700 B.n249 B.n212 585
R701 B.n251 B.n250 585
R702 B.n252 B.n211 585
R703 B.n254 B.n253 585
R704 B.n255 B.n210 585
R705 B.n257 B.n256 585
R706 B.n258 B.n209 585
R707 B.n260 B.n259 585
R708 B.n261 B.n208 585
R709 B.n263 B.n262 585
R710 B.n264 B.n207 585
R711 B.n266 B.n265 585
R712 B.n267 B.n206 585
R713 B.n269 B.n268 585
R714 B.n270 B.n205 585
R715 B.n272 B.n271 585
R716 B.n273 B.n204 585
R717 B.n275 B.n274 585
R718 B.n276 B.n203 585
R719 B.n278 B.n277 585
R720 B.n279 B.n202 585
R721 B.n281 B.n280 585
R722 B.n282 B.n201 585
R723 B.n284 B.n283 585
R724 B.n285 B.n200 585
R725 B.n287 B.n286 585
R726 B.n288 B.n199 585
R727 B.n290 B.n289 585
R728 B.n291 B.n198 585
R729 B.n293 B.n292 585
R730 B.n294 B.n197 585
R731 B.n295 B.n294 506.916
R732 B.n467 B.n466 506.916
R733 B.n621 B.n88 506.916
R734 B.n790 B.n27 506.916
R735 B.n370 B.t6 385.091
R736 B.n165 B.t9 385.091
R737 B.n61 B.t3 385.091
R738 B.n54 B.t0 385.091
R739 B.n865 B.n864 256.663
R740 B.n864 B.n863 235.042
R741 B.n864 B.n2 235.042
R742 B.n295 B.n196 163.367
R743 B.n299 B.n196 163.367
R744 B.n300 B.n299 163.367
R745 B.n301 B.n300 163.367
R746 B.n301 B.n194 163.367
R747 B.n305 B.n194 163.367
R748 B.n306 B.n305 163.367
R749 B.n307 B.n306 163.367
R750 B.n307 B.n192 163.367
R751 B.n311 B.n192 163.367
R752 B.n312 B.n311 163.367
R753 B.n313 B.n312 163.367
R754 B.n313 B.n190 163.367
R755 B.n317 B.n190 163.367
R756 B.n318 B.n317 163.367
R757 B.n319 B.n318 163.367
R758 B.n319 B.n188 163.367
R759 B.n323 B.n188 163.367
R760 B.n324 B.n323 163.367
R761 B.n325 B.n324 163.367
R762 B.n325 B.n186 163.367
R763 B.n329 B.n186 163.367
R764 B.n330 B.n329 163.367
R765 B.n331 B.n330 163.367
R766 B.n331 B.n184 163.367
R767 B.n335 B.n184 163.367
R768 B.n336 B.n335 163.367
R769 B.n337 B.n336 163.367
R770 B.n337 B.n182 163.367
R771 B.n341 B.n182 163.367
R772 B.n342 B.n341 163.367
R773 B.n343 B.n342 163.367
R774 B.n343 B.n180 163.367
R775 B.n347 B.n180 163.367
R776 B.n348 B.n347 163.367
R777 B.n349 B.n348 163.367
R778 B.n349 B.n178 163.367
R779 B.n353 B.n178 163.367
R780 B.n354 B.n353 163.367
R781 B.n355 B.n354 163.367
R782 B.n355 B.n176 163.367
R783 B.n359 B.n176 163.367
R784 B.n360 B.n359 163.367
R785 B.n361 B.n360 163.367
R786 B.n361 B.n174 163.367
R787 B.n365 B.n174 163.367
R788 B.n366 B.n365 163.367
R789 B.n367 B.n366 163.367
R790 B.n367 B.n172 163.367
R791 B.n374 B.n172 163.367
R792 B.n375 B.n374 163.367
R793 B.n376 B.n375 163.367
R794 B.n376 B.n170 163.367
R795 B.n380 B.n170 163.367
R796 B.n381 B.n380 163.367
R797 B.n382 B.n381 163.367
R798 B.n382 B.n168 163.367
R799 B.n386 B.n168 163.367
R800 B.n387 B.n386 163.367
R801 B.n388 B.n387 163.367
R802 B.n388 B.n164 163.367
R803 B.n393 B.n164 163.367
R804 B.n394 B.n393 163.367
R805 B.n395 B.n394 163.367
R806 B.n395 B.n162 163.367
R807 B.n399 B.n162 163.367
R808 B.n400 B.n399 163.367
R809 B.n401 B.n400 163.367
R810 B.n401 B.n160 163.367
R811 B.n405 B.n160 163.367
R812 B.n406 B.n405 163.367
R813 B.n407 B.n406 163.367
R814 B.n407 B.n158 163.367
R815 B.n411 B.n158 163.367
R816 B.n412 B.n411 163.367
R817 B.n413 B.n412 163.367
R818 B.n413 B.n156 163.367
R819 B.n417 B.n156 163.367
R820 B.n418 B.n417 163.367
R821 B.n419 B.n418 163.367
R822 B.n419 B.n154 163.367
R823 B.n423 B.n154 163.367
R824 B.n424 B.n423 163.367
R825 B.n425 B.n424 163.367
R826 B.n425 B.n152 163.367
R827 B.n429 B.n152 163.367
R828 B.n430 B.n429 163.367
R829 B.n431 B.n430 163.367
R830 B.n431 B.n150 163.367
R831 B.n435 B.n150 163.367
R832 B.n436 B.n435 163.367
R833 B.n437 B.n436 163.367
R834 B.n437 B.n148 163.367
R835 B.n441 B.n148 163.367
R836 B.n442 B.n441 163.367
R837 B.n443 B.n442 163.367
R838 B.n443 B.n146 163.367
R839 B.n447 B.n146 163.367
R840 B.n448 B.n447 163.367
R841 B.n449 B.n448 163.367
R842 B.n449 B.n144 163.367
R843 B.n453 B.n144 163.367
R844 B.n454 B.n453 163.367
R845 B.n455 B.n454 163.367
R846 B.n455 B.n142 163.367
R847 B.n459 B.n142 163.367
R848 B.n460 B.n459 163.367
R849 B.n461 B.n460 163.367
R850 B.n461 B.n140 163.367
R851 B.n465 B.n140 163.367
R852 B.n466 B.n465 163.367
R853 B.n617 B.n88 163.367
R854 B.n617 B.n616 163.367
R855 B.n616 B.n615 163.367
R856 B.n615 B.n90 163.367
R857 B.n611 B.n90 163.367
R858 B.n611 B.n610 163.367
R859 B.n610 B.n609 163.367
R860 B.n609 B.n92 163.367
R861 B.n605 B.n92 163.367
R862 B.n605 B.n604 163.367
R863 B.n604 B.n603 163.367
R864 B.n603 B.n94 163.367
R865 B.n599 B.n94 163.367
R866 B.n599 B.n598 163.367
R867 B.n598 B.n597 163.367
R868 B.n597 B.n96 163.367
R869 B.n593 B.n96 163.367
R870 B.n593 B.n592 163.367
R871 B.n592 B.n591 163.367
R872 B.n591 B.n98 163.367
R873 B.n587 B.n98 163.367
R874 B.n587 B.n586 163.367
R875 B.n586 B.n585 163.367
R876 B.n585 B.n100 163.367
R877 B.n581 B.n100 163.367
R878 B.n581 B.n580 163.367
R879 B.n580 B.n579 163.367
R880 B.n579 B.n102 163.367
R881 B.n575 B.n102 163.367
R882 B.n575 B.n574 163.367
R883 B.n574 B.n573 163.367
R884 B.n573 B.n104 163.367
R885 B.n569 B.n104 163.367
R886 B.n569 B.n568 163.367
R887 B.n568 B.n567 163.367
R888 B.n567 B.n106 163.367
R889 B.n563 B.n106 163.367
R890 B.n563 B.n562 163.367
R891 B.n562 B.n561 163.367
R892 B.n561 B.n108 163.367
R893 B.n557 B.n108 163.367
R894 B.n557 B.n556 163.367
R895 B.n556 B.n555 163.367
R896 B.n555 B.n110 163.367
R897 B.n551 B.n110 163.367
R898 B.n551 B.n550 163.367
R899 B.n550 B.n549 163.367
R900 B.n549 B.n112 163.367
R901 B.n545 B.n112 163.367
R902 B.n545 B.n544 163.367
R903 B.n544 B.n543 163.367
R904 B.n543 B.n114 163.367
R905 B.n539 B.n114 163.367
R906 B.n539 B.n538 163.367
R907 B.n538 B.n537 163.367
R908 B.n537 B.n116 163.367
R909 B.n533 B.n116 163.367
R910 B.n533 B.n532 163.367
R911 B.n532 B.n531 163.367
R912 B.n531 B.n118 163.367
R913 B.n527 B.n118 163.367
R914 B.n527 B.n526 163.367
R915 B.n526 B.n525 163.367
R916 B.n525 B.n120 163.367
R917 B.n521 B.n120 163.367
R918 B.n521 B.n520 163.367
R919 B.n520 B.n519 163.367
R920 B.n519 B.n122 163.367
R921 B.n515 B.n122 163.367
R922 B.n515 B.n514 163.367
R923 B.n514 B.n513 163.367
R924 B.n513 B.n124 163.367
R925 B.n509 B.n124 163.367
R926 B.n509 B.n508 163.367
R927 B.n508 B.n507 163.367
R928 B.n507 B.n126 163.367
R929 B.n503 B.n126 163.367
R930 B.n503 B.n502 163.367
R931 B.n502 B.n501 163.367
R932 B.n501 B.n128 163.367
R933 B.n497 B.n128 163.367
R934 B.n497 B.n496 163.367
R935 B.n496 B.n495 163.367
R936 B.n495 B.n130 163.367
R937 B.n491 B.n130 163.367
R938 B.n491 B.n490 163.367
R939 B.n490 B.n489 163.367
R940 B.n489 B.n132 163.367
R941 B.n485 B.n132 163.367
R942 B.n485 B.n484 163.367
R943 B.n484 B.n483 163.367
R944 B.n483 B.n134 163.367
R945 B.n479 B.n134 163.367
R946 B.n479 B.n478 163.367
R947 B.n478 B.n477 163.367
R948 B.n477 B.n136 163.367
R949 B.n473 B.n136 163.367
R950 B.n473 B.n472 163.367
R951 B.n472 B.n471 163.367
R952 B.n471 B.n138 163.367
R953 B.n467 B.n138 163.367
R954 B.n786 B.n27 163.367
R955 B.n786 B.n785 163.367
R956 B.n785 B.n784 163.367
R957 B.n784 B.n29 163.367
R958 B.n780 B.n29 163.367
R959 B.n780 B.n779 163.367
R960 B.n779 B.n778 163.367
R961 B.n778 B.n31 163.367
R962 B.n774 B.n31 163.367
R963 B.n774 B.n773 163.367
R964 B.n773 B.n772 163.367
R965 B.n772 B.n33 163.367
R966 B.n768 B.n33 163.367
R967 B.n768 B.n767 163.367
R968 B.n767 B.n766 163.367
R969 B.n766 B.n35 163.367
R970 B.n762 B.n35 163.367
R971 B.n762 B.n761 163.367
R972 B.n761 B.n760 163.367
R973 B.n760 B.n37 163.367
R974 B.n756 B.n37 163.367
R975 B.n756 B.n755 163.367
R976 B.n755 B.n754 163.367
R977 B.n754 B.n39 163.367
R978 B.n750 B.n39 163.367
R979 B.n750 B.n749 163.367
R980 B.n749 B.n748 163.367
R981 B.n748 B.n41 163.367
R982 B.n744 B.n41 163.367
R983 B.n744 B.n743 163.367
R984 B.n743 B.n742 163.367
R985 B.n742 B.n43 163.367
R986 B.n738 B.n43 163.367
R987 B.n738 B.n737 163.367
R988 B.n737 B.n736 163.367
R989 B.n736 B.n45 163.367
R990 B.n732 B.n45 163.367
R991 B.n732 B.n731 163.367
R992 B.n731 B.n730 163.367
R993 B.n730 B.n47 163.367
R994 B.n726 B.n47 163.367
R995 B.n726 B.n725 163.367
R996 B.n725 B.n724 163.367
R997 B.n724 B.n49 163.367
R998 B.n720 B.n49 163.367
R999 B.n720 B.n719 163.367
R1000 B.n719 B.n718 163.367
R1001 B.n718 B.n51 163.367
R1002 B.n714 B.n51 163.367
R1003 B.n714 B.n713 163.367
R1004 B.n713 B.n712 163.367
R1005 B.n712 B.n53 163.367
R1006 B.n708 B.n53 163.367
R1007 B.n708 B.n707 163.367
R1008 B.n707 B.n706 163.367
R1009 B.n706 B.n58 163.367
R1010 B.n702 B.n58 163.367
R1011 B.n702 B.n701 163.367
R1012 B.n701 B.n700 163.367
R1013 B.n700 B.n60 163.367
R1014 B.n695 B.n60 163.367
R1015 B.n695 B.n694 163.367
R1016 B.n694 B.n693 163.367
R1017 B.n693 B.n64 163.367
R1018 B.n689 B.n64 163.367
R1019 B.n689 B.n688 163.367
R1020 B.n688 B.n687 163.367
R1021 B.n687 B.n66 163.367
R1022 B.n683 B.n66 163.367
R1023 B.n683 B.n682 163.367
R1024 B.n682 B.n681 163.367
R1025 B.n681 B.n68 163.367
R1026 B.n677 B.n68 163.367
R1027 B.n677 B.n676 163.367
R1028 B.n676 B.n675 163.367
R1029 B.n675 B.n70 163.367
R1030 B.n671 B.n70 163.367
R1031 B.n671 B.n670 163.367
R1032 B.n670 B.n669 163.367
R1033 B.n669 B.n72 163.367
R1034 B.n665 B.n72 163.367
R1035 B.n665 B.n664 163.367
R1036 B.n664 B.n663 163.367
R1037 B.n663 B.n74 163.367
R1038 B.n659 B.n74 163.367
R1039 B.n659 B.n658 163.367
R1040 B.n658 B.n657 163.367
R1041 B.n657 B.n76 163.367
R1042 B.n653 B.n76 163.367
R1043 B.n653 B.n652 163.367
R1044 B.n652 B.n651 163.367
R1045 B.n651 B.n78 163.367
R1046 B.n647 B.n78 163.367
R1047 B.n647 B.n646 163.367
R1048 B.n646 B.n645 163.367
R1049 B.n645 B.n80 163.367
R1050 B.n641 B.n80 163.367
R1051 B.n641 B.n640 163.367
R1052 B.n640 B.n639 163.367
R1053 B.n639 B.n82 163.367
R1054 B.n635 B.n82 163.367
R1055 B.n635 B.n634 163.367
R1056 B.n634 B.n633 163.367
R1057 B.n633 B.n84 163.367
R1058 B.n629 B.n84 163.367
R1059 B.n629 B.n628 163.367
R1060 B.n628 B.n627 163.367
R1061 B.n627 B.n86 163.367
R1062 B.n623 B.n86 163.367
R1063 B.n623 B.n622 163.367
R1064 B.n622 B.n621 163.367
R1065 B.n791 B.n790 163.367
R1066 B.n792 B.n791 163.367
R1067 B.n792 B.n25 163.367
R1068 B.n796 B.n25 163.367
R1069 B.n797 B.n796 163.367
R1070 B.n798 B.n797 163.367
R1071 B.n798 B.n23 163.367
R1072 B.n802 B.n23 163.367
R1073 B.n803 B.n802 163.367
R1074 B.n804 B.n803 163.367
R1075 B.n804 B.n21 163.367
R1076 B.n808 B.n21 163.367
R1077 B.n809 B.n808 163.367
R1078 B.n810 B.n809 163.367
R1079 B.n810 B.n19 163.367
R1080 B.n814 B.n19 163.367
R1081 B.n815 B.n814 163.367
R1082 B.n816 B.n815 163.367
R1083 B.n816 B.n17 163.367
R1084 B.n820 B.n17 163.367
R1085 B.n821 B.n820 163.367
R1086 B.n822 B.n821 163.367
R1087 B.n822 B.n15 163.367
R1088 B.n826 B.n15 163.367
R1089 B.n827 B.n826 163.367
R1090 B.n828 B.n827 163.367
R1091 B.n828 B.n13 163.367
R1092 B.n832 B.n13 163.367
R1093 B.n833 B.n832 163.367
R1094 B.n834 B.n833 163.367
R1095 B.n834 B.n11 163.367
R1096 B.n838 B.n11 163.367
R1097 B.n839 B.n838 163.367
R1098 B.n840 B.n839 163.367
R1099 B.n840 B.n9 163.367
R1100 B.n844 B.n9 163.367
R1101 B.n845 B.n844 163.367
R1102 B.n846 B.n845 163.367
R1103 B.n846 B.n7 163.367
R1104 B.n850 B.n7 163.367
R1105 B.n851 B.n850 163.367
R1106 B.n852 B.n851 163.367
R1107 B.n852 B.n5 163.367
R1108 B.n856 B.n5 163.367
R1109 B.n857 B.n856 163.367
R1110 B.n858 B.n857 163.367
R1111 B.n858 B.n3 163.367
R1112 B.n862 B.n3 163.367
R1113 B.n863 B.n862 163.367
R1114 B.n222 B.n2 163.367
R1115 B.n223 B.n222 163.367
R1116 B.n223 B.n220 163.367
R1117 B.n227 B.n220 163.367
R1118 B.n228 B.n227 163.367
R1119 B.n229 B.n228 163.367
R1120 B.n229 B.n218 163.367
R1121 B.n233 B.n218 163.367
R1122 B.n234 B.n233 163.367
R1123 B.n235 B.n234 163.367
R1124 B.n235 B.n216 163.367
R1125 B.n239 B.n216 163.367
R1126 B.n240 B.n239 163.367
R1127 B.n241 B.n240 163.367
R1128 B.n241 B.n214 163.367
R1129 B.n245 B.n214 163.367
R1130 B.n246 B.n245 163.367
R1131 B.n247 B.n246 163.367
R1132 B.n247 B.n212 163.367
R1133 B.n251 B.n212 163.367
R1134 B.n252 B.n251 163.367
R1135 B.n253 B.n252 163.367
R1136 B.n253 B.n210 163.367
R1137 B.n257 B.n210 163.367
R1138 B.n258 B.n257 163.367
R1139 B.n259 B.n258 163.367
R1140 B.n259 B.n208 163.367
R1141 B.n263 B.n208 163.367
R1142 B.n264 B.n263 163.367
R1143 B.n265 B.n264 163.367
R1144 B.n265 B.n206 163.367
R1145 B.n269 B.n206 163.367
R1146 B.n270 B.n269 163.367
R1147 B.n271 B.n270 163.367
R1148 B.n271 B.n204 163.367
R1149 B.n275 B.n204 163.367
R1150 B.n276 B.n275 163.367
R1151 B.n277 B.n276 163.367
R1152 B.n277 B.n202 163.367
R1153 B.n281 B.n202 163.367
R1154 B.n282 B.n281 163.367
R1155 B.n283 B.n282 163.367
R1156 B.n283 B.n200 163.367
R1157 B.n287 B.n200 163.367
R1158 B.n288 B.n287 163.367
R1159 B.n289 B.n288 163.367
R1160 B.n289 B.n198 163.367
R1161 B.n293 B.n198 163.367
R1162 B.n294 B.n293 163.367
R1163 B.n165 B.t10 159.465
R1164 B.n61 B.t5 159.465
R1165 B.n370 B.t7 159.446
R1166 B.n54 B.t2 159.446
R1167 B.n166 B.t11 112.921
R1168 B.n62 B.t4 112.921
R1169 B.n371 B.t8 112.901
R1170 B.n55 B.t1 112.901
R1171 B.n372 B.n371 59.5399
R1172 B.n390 B.n166 59.5399
R1173 B.n697 B.n62 59.5399
R1174 B.n56 B.n55 59.5399
R1175 B.n371 B.n370 46.546
R1176 B.n166 B.n165 46.546
R1177 B.n62 B.n61 46.546
R1178 B.n55 B.n54 46.546
R1179 B.n789 B.n788 32.9371
R1180 B.n620 B.n619 32.9371
R1181 B.n468 B.n139 32.9371
R1182 B.n296 B.n197 32.9371
R1183 B B.n865 18.0485
R1184 B.n789 B.n26 10.6151
R1185 B.n793 B.n26 10.6151
R1186 B.n794 B.n793 10.6151
R1187 B.n795 B.n794 10.6151
R1188 B.n795 B.n24 10.6151
R1189 B.n799 B.n24 10.6151
R1190 B.n800 B.n799 10.6151
R1191 B.n801 B.n800 10.6151
R1192 B.n801 B.n22 10.6151
R1193 B.n805 B.n22 10.6151
R1194 B.n806 B.n805 10.6151
R1195 B.n807 B.n806 10.6151
R1196 B.n807 B.n20 10.6151
R1197 B.n811 B.n20 10.6151
R1198 B.n812 B.n811 10.6151
R1199 B.n813 B.n812 10.6151
R1200 B.n813 B.n18 10.6151
R1201 B.n817 B.n18 10.6151
R1202 B.n818 B.n817 10.6151
R1203 B.n819 B.n818 10.6151
R1204 B.n819 B.n16 10.6151
R1205 B.n823 B.n16 10.6151
R1206 B.n824 B.n823 10.6151
R1207 B.n825 B.n824 10.6151
R1208 B.n825 B.n14 10.6151
R1209 B.n829 B.n14 10.6151
R1210 B.n830 B.n829 10.6151
R1211 B.n831 B.n830 10.6151
R1212 B.n831 B.n12 10.6151
R1213 B.n835 B.n12 10.6151
R1214 B.n836 B.n835 10.6151
R1215 B.n837 B.n836 10.6151
R1216 B.n837 B.n10 10.6151
R1217 B.n841 B.n10 10.6151
R1218 B.n842 B.n841 10.6151
R1219 B.n843 B.n842 10.6151
R1220 B.n843 B.n8 10.6151
R1221 B.n847 B.n8 10.6151
R1222 B.n848 B.n847 10.6151
R1223 B.n849 B.n848 10.6151
R1224 B.n849 B.n6 10.6151
R1225 B.n853 B.n6 10.6151
R1226 B.n854 B.n853 10.6151
R1227 B.n855 B.n854 10.6151
R1228 B.n855 B.n4 10.6151
R1229 B.n859 B.n4 10.6151
R1230 B.n860 B.n859 10.6151
R1231 B.n861 B.n860 10.6151
R1232 B.n861 B.n0 10.6151
R1233 B.n788 B.n787 10.6151
R1234 B.n787 B.n28 10.6151
R1235 B.n783 B.n28 10.6151
R1236 B.n783 B.n782 10.6151
R1237 B.n782 B.n781 10.6151
R1238 B.n781 B.n30 10.6151
R1239 B.n777 B.n30 10.6151
R1240 B.n777 B.n776 10.6151
R1241 B.n776 B.n775 10.6151
R1242 B.n775 B.n32 10.6151
R1243 B.n771 B.n32 10.6151
R1244 B.n771 B.n770 10.6151
R1245 B.n770 B.n769 10.6151
R1246 B.n769 B.n34 10.6151
R1247 B.n765 B.n34 10.6151
R1248 B.n765 B.n764 10.6151
R1249 B.n764 B.n763 10.6151
R1250 B.n763 B.n36 10.6151
R1251 B.n759 B.n36 10.6151
R1252 B.n759 B.n758 10.6151
R1253 B.n758 B.n757 10.6151
R1254 B.n757 B.n38 10.6151
R1255 B.n753 B.n38 10.6151
R1256 B.n753 B.n752 10.6151
R1257 B.n752 B.n751 10.6151
R1258 B.n751 B.n40 10.6151
R1259 B.n747 B.n40 10.6151
R1260 B.n747 B.n746 10.6151
R1261 B.n746 B.n745 10.6151
R1262 B.n745 B.n42 10.6151
R1263 B.n741 B.n42 10.6151
R1264 B.n741 B.n740 10.6151
R1265 B.n740 B.n739 10.6151
R1266 B.n739 B.n44 10.6151
R1267 B.n735 B.n44 10.6151
R1268 B.n735 B.n734 10.6151
R1269 B.n734 B.n733 10.6151
R1270 B.n733 B.n46 10.6151
R1271 B.n729 B.n46 10.6151
R1272 B.n729 B.n728 10.6151
R1273 B.n728 B.n727 10.6151
R1274 B.n727 B.n48 10.6151
R1275 B.n723 B.n48 10.6151
R1276 B.n723 B.n722 10.6151
R1277 B.n722 B.n721 10.6151
R1278 B.n721 B.n50 10.6151
R1279 B.n717 B.n50 10.6151
R1280 B.n717 B.n716 10.6151
R1281 B.n716 B.n715 10.6151
R1282 B.n715 B.n52 10.6151
R1283 B.n711 B.n710 10.6151
R1284 B.n710 B.n709 10.6151
R1285 B.n709 B.n57 10.6151
R1286 B.n705 B.n57 10.6151
R1287 B.n705 B.n704 10.6151
R1288 B.n704 B.n703 10.6151
R1289 B.n703 B.n59 10.6151
R1290 B.n699 B.n59 10.6151
R1291 B.n699 B.n698 10.6151
R1292 B.n696 B.n63 10.6151
R1293 B.n692 B.n63 10.6151
R1294 B.n692 B.n691 10.6151
R1295 B.n691 B.n690 10.6151
R1296 B.n690 B.n65 10.6151
R1297 B.n686 B.n65 10.6151
R1298 B.n686 B.n685 10.6151
R1299 B.n685 B.n684 10.6151
R1300 B.n684 B.n67 10.6151
R1301 B.n680 B.n67 10.6151
R1302 B.n680 B.n679 10.6151
R1303 B.n679 B.n678 10.6151
R1304 B.n678 B.n69 10.6151
R1305 B.n674 B.n69 10.6151
R1306 B.n674 B.n673 10.6151
R1307 B.n673 B.n672 10.6151
R1308 B.n672 B.n71 10.6151
R1309 B.n668 B.n71 10.6151
R1310 B.n668 B.n667 10.6151
R1311 B.n667 B.n666 10.6151
R1312 B.n666 B.n73 10.6151
R1313 B.n662 B.n73 10.6151
R1314 B.n662 B.n661 10.6151
R1315 B.n661 B.n660 10.6151
R1316 B.n660 B.n75 10.6151
R1317 B.n656 B.n75 10.6151
R1318 B.n656 B.n655 10.6151
R1319 B.n655 B.n654 10.6151
R1320 B.n654 B.n77 10.6151
R1321 B.n650 B.n77 10.6151
R1322 B.n650 B.n649 10.6151
R1323 B.n649 B.n648 10.6151
R1324 B.n648 B.n79 10.6151
R1325 B.n644 B.n79 10.6151
R1326 B.n644 B.n643 10.6151
R1327 B.n643 B.n642 10.6151
R1328 B.n642 B.n81 10.6151
R1329 B.n638 B.n81 10.6151
R1330 B.n638 B.n637 10.6151
R1331 B.n637 B.n636 10.6151
R1332 B.n636 B.n83 10.6151
R1333 B.n632 B.n83 10.6151
R1334 B.n632 B.n631 10.6151
R1335 B.n631 B.n630 10.6151
R1336 B.n630 B.n85 10.6151
R1337 B.n626 B.n85 10.6151
R1338 B.n626 B.n625 10.6151
R1339 B.n625 B.n624 10.6151
R1340 B.n624 B.n87 10.6151
R1341 B.n620 B.n87 10.6151
R1342 B.n619 B.n618 10.6151
R1343 B.n618 B.n89 10.6151
R1344 B.n614 B.n89 10.6151
R1345 B.n614 B.n613 10.6151
R1346 B.n613 B.n612 10.6151
R1347 B.n612 B.n91 10.6151
R1348 B.n608 B.n91 10.6151
R1349 B.n608 B.n607 10.6151
R1350 B.n607 B.n606 10.6151
R1351 B.n606 B.n93 10.6151
R1352 B.n602 B.n93 10.6151
R1353 B.n602 B.n601 10.6151
R1354 B.n601 B.n600 10.6151
R1355 B.n600 B.n95 10.6151
R1356 B.n596 B.n95 10.6151
R1357 B.n596 B.n595 10.6151
R1358 B.n595 B.n594 10.6151
R1359 B.n594 B.n97 10.6151
R1360 B.n590 B.n97 10.6151
R1361 B.n590 B.n589 10.6151
R1362 B.n589 B.n588 10.6151
R1363 B.n588 B.n99 10.6151
R1364 B.n584 B.n99 10.6151
R1365 B.n584 B.n583 10.6151
R1366 B.n583 B.n582 10.6151
R1367 B.n582 B.n101 10.6151
R1368 B.n578 B.n101 10.6151
R1369 B.n578 B.n577 10.6151
R1370 B.n577 B.n576 10.6151
R1371 B.n576 B.n103 10.6151
R1372 B.n572 B.n103 10.6151
R1373 B.n572 B.n571 10.6151
R1374 B.n571 B.n570 10.6151
R1375 B.n570 B.n105 10.6151
R1376 B.n566 B.n105 10.6151
R1377 B.n566 B.n565 10.6151
R1378 B.n565 B.n564 10.6151
R1379 B.n564 B.n107 10.6151
R1380 B.n560 B.n107 10.6151
R1381 B.n560 B.n559 10.6151
R1382 B.n559 B.n558 10.6151
R1383 B.n558 B.n109 10.6151
R1384 B.n554 B.n109 10.6151
R1385 B.n554 B.n553 10.6151
R1386 B.n553 B.n552 10.6151
R1387 B.n552 B.n111 10.6151
R1388 B.n548 B.n111 10.6151
R1389 B.n548 B.n547 10.6151
R1390 B.n547 B.n546 10.6151
R1391 B.n546 B.n113 10.6151
R1392 B.n542 B.n113 10.6151
R1393 B.n542 B.n541 10.6151
R1394 B.n541 B.n540 10.6151
R1395 B.n540 B.n115 10.6151
R1396 B.n536 B.n115 10.6151
R1397 B.n536 B.n535 10.6151
R1398 B.n535 B.n534 10.6151
R1399 B.n534 B.n117 10.6151
R1400 B.n530 B.n117 10.6151
R1401 B.n530 B.n529 10.6151
R1402 B.n529 B.n528 10.6151
R1403 B.n528 B.n119 10.6151
R1404 B.n524 B.n119 10.6151
R1405 B.n524 B.n523 10.6151
R1406 B.n523 B.n522 10.6151
R1407 B.n522 B.n121 10.6151
R1408 B.n518 B.n121 10.6151
R1409 B.n518 B.n517 10.6151
R1410 B.n517 B.n516 10.6151
R1411 B.n516 B.n123 10.6151
R1412 B.n512 B.n123 10.6151
R1413 B.n512 B.n511 10.6151
R1414 B.n511 B.n510 10.6151
R1415 B.n510 B.n125 10.6151
R1416 B.n506 B.n125 10.6151
R1417 B.n506 B.n505 10.6151
R1418 B.n505 B.n504 10.6151
R1419 B.n504 B.n127 10.6151
R1420 B.n500 B.n127 10.6151
R1421 B.n500 B.n499 10.6151
R1422 B.n499 B.n498 10.6151
R1423 B.n498 B.n129 10.6151
R1424 B.n494 B.n129 10.6151
R1425 B.n494 B.n493 10.6151
R1426 B.n493 B.n492 10.6151
R1427 B.n492 B.n131 10.6151
R1428 B.n488 B.n131 10.6151
R1429 B.n488 B.n487 10.6151
R1430 B.n487 B.n486 10.6151
R1431 B.n486 B.n133 10.6151
R1432 B.n482 B.n133 10.6151
R1433 B.n482 B.n481 10.6151
R1434 B.n481 B.n480 10.6151
R1435 B.n480 B.n135 10.6151
R1436 B.n476 B.n135 10.6151
R1437 B.n476 B.n475 10.6151
R1438 B.n475 B.n474 10.6151
R1439 B.n474 B.n137 10.6151
R1440 B.n470 B.n137 10.6151
R1441 B.n470 B.n469 10.6151
R1442 B.n469 B.n468 10.6151
R1443 B.n221 B.n1 10.6151
R1444 B.n224 B.n221 10.6151
R1445 B.n225 B.n224 10.6151
R1446 B.n226 B.n225 10.6151
R1447 B.n226 B.n219 10.6151
R1448 B.n230 B.n219 10.6151
R1449 B.n231 B.n230 10.6151
R1450 B.n232 B.n231 10.6151
R1451 B.n232 B.n217 10.6151
R1452 B.n236 B.n217 10.6151
R1453 B.n237 B.n236 10.6151
R1454 B.n238 B.n237 10.6151
R1455 B.n238 B.n215 10.6151
R1456 B.n242 B.n215 10.6151
R1457 B.n243 B.n242 10.6151
R1458 B.n244 B.n243 10.6151
R1459 B.n244 B.n213 10.6151
R1460 B.n248 B.n213 10.6151
R1461 B.n249 B.n248 10.6151
R1462 B.n250 B.n249 10.6151
R1463 B.n250 B.n211 10.6151
R1464 B.n254 B.n211 10.6151
R1465 B.n255 B.n254 10.6151
R1466 B.n256 B.n255 10.6151
R1467 B.n256 B.n209 10.6151
R1468 B.n260 B.n209 10.6151
R1469 B.n261 B.n260 10.6151
R1470 B.n262 B.n261 10.6151
R1471 B.n262 B.n207 10.6151
R1472 B.n266 B.n207 10.6151
R1473 B.n267 B.n266 10.6151
R1474 B.n268 B.n267 10.6151
R1475 B.n268 B.n205 10.6151
R1476 B.n272 B.n205 10.6151
R1477 B.n273 B.n272 10.6151
R1478 B.n274 B.n273 10.6151
R1479 B.n274 B.n203 10.6151
R1480 B.n278 B.n203 10.6151
R1481 B.n279 B.n278 10.6151
R1482 B.n280 B.n279 10.6151
R1483 B.n280 B.n201 10.6151
R1484 B.n284 B.n201 10.6151
R1485 B.n285 B.n284 10.6151
R1486 B.n286 B.n285 10.6151
R1487 B.n286 B.n199 10.6151
R1488 B.n290 B.n199 10.6151
R1489 B.n291 B.n290 10.6151
R1490 B.n292 B.n291 10.6151
R1491 B.n292 B.n197 10.6151
R1492 B.n297 B.n296 10.6151
R1493 B.n298 B.n297 10.6151
R1494 B.n298 B.n195 10.6151
R1495 B.n302 B.n195 10.6151
R1496 B.n303 B.n302 10.6151
R1497 B.n304 B.n303 10.6151
R1498 B.n304 B.n193 10.6151
R1499 B.n308 B.n193 10.6151
R1500 B.n309 B.n308 10.6151
R1501 B.n310 B.n309 10.6151
R1502 B.n310 B.n191 10.6151
R1503 B.n314 B.n191 10.6151
R1504 B.n315 B.n314 10.6151
R1505 B.n316 B.n315 10.6151
R1506 B.n316 B.n189 10.6151
R1507 B.n320 B.n189 10.6151
R1508 B.n321 B.n320 10.6151
R1509 B.n322 B.n321 10.6151
R1510 B.n322 B.n187 10.6151
R1511 B.n326 B.n187 10.6151
R1512 B.n327 B.n326 10.6151
R1513 B.n328 B.n327 10.6151
R1514 B.n328 B.n185 10.6151
R1515 B.n332 B.n185 10.6151
R1516 B.n333 B.n332 10.6151
R1517 B.n334 B.n333 10.6151
R1518 B.n334 B.n183 10.6151
R1519 B.n338 B.n183 10.6151
R1520 B.n339 B.n338 10.6151
R1521 B.n340 B.n339 10.6151
R1522 B.n340 B.n181 10.6151
R1523 B.n344 B.n181 10.6151
R1524 B.n345 B.n344 10.6151
R1525 B.n346 B.n345 10.6151
R1526 B.n346 B.n179 10.6151
R1527 B.n350 B.n179 10.6151
R1528 B.n351 B.n350 10.6151
R1529 B.n352 B.n351 10.6151
R1530 B.n352 B.n177 10.6151
R1531 B.n356 B.n177 10.6151
R1532 B.n357 B.n356 10.6151
R1533 B.n358 B.n357 10.6151
R1534 B.n358 B.n175 10.6151
R1535 B.n362 B.n175 10.6151
R1536 B.n363 B.n362 10.6151
R1537 B.n364 B.n363 10.6151
R1538 B.n364 B.n173 10.6151
R1539 B.n368 B.n173 10.6151
R1540 B.n369 B.n368 10.6151
R1541 B.n373 B.n369 10.6151
R1542 B.n377 B.n171 10.6151
R1543 B.n378 B.n377 10.6151
R1544 B.n379 B.n378 10.6151
R1545 B.n379 B.n169 10.6151
R1546 B.n383 B.n169 10.6151
R1547 B.n384 B.n383 10.6151
R1548 B.n385 B.n384 10.6151
R1549 B.n385 B.n167 10.6151
R1550 B.n389 B.n167 10.6151
R1551 B.n392 B.n391 10.6151
R1552 B.n392 B.n163 10.6151
R1553 B.n396 B.n163 10.6151
R1554 B.n397 B.n396 10.6151
R1555 B.n398 B.n397 10.6151
R1556 B.n398 B.n161 10.6151
R1557 B.n402 B.n161 10.6151
R1558 B.n403 B.n402 10.6151
R1559 B.n404 B.n403 10.6151
R1560 B.n404 B.n159 10.6151
R1561 B.n408 B.n159 10.6151
R1562 B.n409 B.n408 10.6151
R1563 B.n410 B.n409 10.6151
R1564 B.n410 B.n157 10.6151
R1565 B.n414 B.n157 10.6151
R1566 B.n415 B.n414 10.6151
R1567 B.n416 B.n415 10.6151
R1568 B.n416 B.n155 10.6151
R1569 B.n420 B.n155 10.6151
R1570 B.n421 B.n420 10.6151
R1571 B.n422 B.n421 10.6151
R1572 B.n422 B.n153 10.6151
R1573 B.n426 B.n153 10.6151
R1574 B.n427 B.n426 10.6151
R1575 B.n428 B.n427 10.6151
R1576 B.n428 B.n151 10.6151
R1577 B.n432 B.n151 10.6151
R1578 B.n433 B.n432 10.6151
R1579 B.n434 B.n433 10.6151
R1580 B.n434 B.n149 10.6151
R1581 B.n438 B.n149 10.6151
R1582 B.n439 B.n438 10.6151
R1583 B.n440 B.n439 10.6151
R1584 B.n440 B.n147 10.6151
R1585 B.n444 B.n147 10.6151
R1586 B.n445 B.n444 10.6151
R1587 B.n446 B.n445 10.6151
R1588 B.n446 B.n145 10.6151
R1589 B.n450 B.n145 10.6151
R1590 B.n451 B.n450 10.6151
R1591 B.n452 B.n451 10.6151
R1592 B.n452 B.n143 10.6151
R1593 B.n456 B.n143 10.6151
R1594 B.n457 B.n456 10.6151
R1595 B.n458 B.n457 10.6151
R1596 B.n458 B.n141 10.6151
R1597 B.n462 B.n141 10.6151
R1598 B.n463 B.n462 10.6151
R1599 B.n464 B.n463 10.6151
R1600 B.n464 B.n139 10.6151
R1601 B.n56 B.n52 9.36635
R1602 B.n697 B.n696 9.36635
R1603 B.n373 B.n372 9.36635
R1604 B.n391 B.n390 9.36635
R1605 B.n865 B.n0 8.11757
R1606 B.n865 B.n1 8.11757
R1607 B.n711 B.n56 1.24928
R1608 B.n698 B.n697 1.24928
R1609 B.n372 B.n171 1.24928
R1610 B.n390 B.n389 1.24928
C0 VDD2 B 2.6252f
C1 VP VTAIL 13.0795f
C2 B VTAIL 4.20541f
C3 VDD1 w_n3850_n4026# 2.81896f
C4 VDD2 VTAIL 12.169299f
C5 VN w_n3850_n4026# 8.143229f
C6 VP VDD1 13.1431f
C7 VP VN 8.23041f
C8 B VDD1 2.52792f
C9 B VN 1.18718f
C10 VDD2 VDD1 1.83024f
C11 VDD2 VN 12.7835f
C12 VDD1 VTAIL 12.123501f
C13 VN VTAIL 13.0651f
C14 VP w_n3850_n4026# 8.642839f
C15 VDD1 VN 0.152175f
C16 B w_n3850_n4026# 10.577901f
C17 VDD2 w_n3850_n4026# 2.93506f
C18 w_n3850_n4026# VTAIL 3.61233f
C19 VP B 2.02439f
C20 VDD2 VP 0.516332f
C21 VDD2 VSUBS 2.02188f
C22 VDD1 VSUBS 1.822433f
C23 VTAIL VSUBS 1.288598f
C24 VN VSUBS 6.96158f
C25 VP VSUBS 3.685325f
C26 B VSUBS 4.986558f
C27 w_n3850_n4026# VSUBS 0.190021p
C28 B.n0 VSUBS 0.007836f
C29 B.n1 VSUBS 0.007836f
C30 B.n2 VSUBS 0.011588f
C31 B.n3 VSUBS 0.00888f
C32 B.n4 VSUBS 0.00888f
C33 B.n5 VSUBS 0.00888f
C34 B.n6 VSUBS 0.00888f
C35 B.n7 VSUBS 0.00888f
C36 B.n8 VSUBS 0.00888f
C37 B.n9 VSUBS 0.00888f
C38 B.n10 VSUBS 0.00888f
C39 B.n11 VSUBS 0.00888f
C40 B.n12 VSUBS 0.00888f
C41 B.n13 VSUBS 0.00888f
C42 B.n14 VSUBS 0.00888f
C43 B.n15 VSUBS 0.00888f
C44 B.n16 VSUBS 0.00888f
C45 B.n17 VSUBS 0.00888f
C46 B.n18 VSUBS 0.00888f
C47 B.n19 VSUBS 0.00888f
C48 B.n20 VSUBS 0.00888f
C49 B.n21 VSUBS 0.00888f
C50 B.n22 VSUBS 0.00888f
C51 B.n23 VSUBS 0.00888f
C52 B.n24 VSUBS 0.00888f
C53 B.n25 VSUBS 0.00888f
C54 B.n26 VSUBS 0.00888f
C55 B.n27 VSUBS 0.021289f
C56 B.n28 VSUBS 0.00888f
C57 B.n29 VSUBS 0.00888f
C58 B.n30 VSUBS 0.00888f
C59 B.n31 VSUBS 0.00888f
C60 B.n32 VSUBS 0.00888f
C61 B.n33 VSUBS 0.00888f
C62 B.n34 VSUBS 0.00888f
C63 B.n35 VSUBS 0.00888f
C64 B.n36 VSUBS 0.00888f
C65 B.n37 VSUBS 0.00888f
C66 B.n38 VSUBS 0.00888f
C67 B.n39 VSUBS 0.00888f
C68 B.n40 VSUBS 0.00888f
C69 B.n41 VSUBS 0.00888f
C70 B.n42 VSUBS 0.00888f
C71 B.n43 VSUBS 0.00888f
C72 B.n44 VSUBS 0.00888f
C73 B.n45 VSUBS 0.00888f
C74 B.n46 VSUBS 0.00888f
C75 B.n47 VSUBS 0.00888f
C76 B.n48 VSUBS 0.00888f
C77 B.n49 VSUBS 0.00888f
C78 B.n50 VSUBS 0.00888f
C79 B.n51 VSUBS 0.00888f
C80 B.n52 VSUBS 0.008358f
C81 B.n53 VSUBS 0.00888f
C82 B.t1 VSUBS 0.646789f
C83 B.t2 VSUBS 0.668935f
C84 B.t0 VSUBS 1.77045f
C85 B.n54 VSUBS 0.331708f
C86 B.n55 VSUBS 0.088528f
C87 B.n56 VSUBS 0.020575f
C88 B.n57 VSUBS 0.00888f
C89 B.n58 VSUBS 0.00888f
C90 B.n59 VSUBS 0.00888f
C91 B.n60 VSUBS 0.00888f
C92 B.t4 VSUBS 0.646771f
C93 B.t5 VSUBS 0.668919f
C94 B.t3 VSUBS 1.77045f
C95 B.n61 VSUBS 0.331724f
C96 B.n62 VSUBS 0.088546f
C97 B.n63 VSUBS 0.00888f
C98 B.n64 VSUBS 0.00888f
C99 B.n65 VSUBS 0.00888f
C100 B.n66 VSUBS 0.00888f
C101 B.n67 VSUBS 0.00888f
C102 B.n68 VSUBS 0.00888f
C103 B.n69 VSUBS 0.00888f
C104 B.n70 VSUBS 0.00888f
C105 B.n71 VSUBS 0.00888f
C106 B.n72 VSUBS 0.00888f
C107 B.n73 VSUBS 0.00888f
C108 B.n74 VSUBS 0.00888f
C109 B.n75 VSUBS 0.00888f
C110 B.n76 VSUBS 0.00888f
C111 B.n77 VSUBS 0.00888f
C112 B.n78 VSUBS 0.00888f
C113 B.n79 VSUBS 0.00888f
C114 B.n80 VSUBS 0.00888f
C115 B.n81 VSUBS 0.00888f
C116 B.n82 VSUBS 0.00888f
C117 B.n83 VSUBS 0.00888f
C118 B.n84 VSUBS 0.00888f
C119 B.n85 VSUBS 0.00888f
C120 B.n86 VSUBS 0.00888f
C121 B.n87 VSUBS 0.00888f
C122 B.n88 VSUBS 0.020502f
C123 B.n89 VSUBS 0.00888f
C124 B.n90 VSUBS 0.00888f
C125 B.n91 VSUBS 0.00888f
C126 B.n92 VSUBS 0.00888f
C127 B.n93 VSUBS 0.00888f
C128 B.n94 VSUBS 0.00888f
C129 B.n95 VSUBS 0.00888f
C130 B.n96 VSUBS 0.00888f
C131 B.n97 VSUBS 0.00888f
C132 B.n98 VSUBS 0.00888f
C133 B.n99 VSUBS 0.00888f
C134 B.n100 VSUBS 0.00888f
C135 B.n101 VSUBS 0.00888f
C136 B.n102 VSUBS 0.00888f
C137 B.n103 VSUBS 0.00888f
C138 B.n104 VSUBS 0.00888f
C139 B.n105 VSUBS 0.00888f
C140 B.n106 VSUBS 0.00888f
C141 B.n107 VSUBS 0.00888f
C142 B.n108 VSUBS 0.00888f
C143 B.n109 VSUBS 0.00888f
C144 B.n110 VSUBS 0.00888f
C145 B.n111 VSUBS 0.00888f
C146 B.n112 VSUBS 0.00888f
C147 B.n113 VSUBS 0.00888f
C148 B.n114 VSUBS 0.00888f
C149 B.n115 VSUBS 0.00888f
C150 B.n116 VSUBS 0.00888f
C151 B.n117 VSUBS 0.00888f
C152 B.n118 VSUBS 0.00888f
C153 B.n119 VSUBS 0.00888f
C154 B.n120 VSUBS 0.00888f
C155 B.n121 VSUBS 0.00888f
C156 B.n122 VSUBS 0.00888f
C157 B.n123 VSUBS 0.00888f
C158 B.n124 VSUBS 0.00888f
C159 B.n125 VSUBS 0.00888f
C160 B.n126 VSUBS 0.00888f
C161 B.n127 VSUBS 0.00888f
C162 B.n128 VSUBS 0.00888f
C163 B.n129 VSUBS 0.00888f
C164 B.n130 VSUBS 0.00888f
C165 B.n131 VSUBS 0.00888f
C166 B.n132 VSUBS 0.00888f
C167 B.n133 VSUBS 0.00888f
C168 B.n134 VSUBS 0.00888f
C169 B.n135 VSUBS 0.00888f
C170 B.n136 VSUBS 0.00888f
C171 B.n137 VSUBS 0.00888f
C172 B.n138 VSUBS 0.00888f
C173 B.n139 VSUBS 0.020248f
C174 B.n140 VSUBS 0.00888f
C175 B.n141 VSUBS 0.00888f
C176 B.n142 VSUBS 0.00888f
C177 B.n143 VSUBS 0.00888f
C178 B.n144 VSUBS 0.00888f
C179 B.n145 VSUBS 0.00888f
C180 B.n146 VSUBS 0.00888f
C181 B.n147 VSUBS 0.00888f
C182 B.n148 VSUBS 0.00888f
C183 B.n149 VSUBS 0.00888f
C184 B.n150 VSUBS 0.00888f
C185 B.n151 VSUBS 0.00888f
C186 B.n152 VSUBS 0.00888f
C187 B.n153 VSUBS 0.00888f
C188 B.n154 VSUBS 0.00888f
C189 B.n155 VSUBS 0.00888f
C190 B.n156 VSUBS 0.00888f
C191 B.n157 VSUBS 0.00888f
C192 B.n158 VSUBS 0.00888f
C193 B.n159 VSUBS 0.00888f
C194 B.n160 VSUBS 0.00888f
C195 B.n161 VSUBS 0.00888f
C196 B.n162 VSUBS 0.00888f
C197 B.n163 VSUBS 0.00888f
C198 B.n164 VSUBS 0.00888f
C199 B.t11 VSUBS 0.646771f
C200 B.t10 VSUBS 0.668919f
C201 B.t9 VSUBS 1.77045f
C202 B.n165 VSUBS 0.331724f
C203 B.n166 VSUBS 0.088546f
C204 B.n167 VSUBS 0.00888f
C205 B.n168 VSUBS 0.00888f
C206 B.n169 VSUBS 0.00888f
C207 B.n170 VSUBS 0.00888f
C208 B.n171 VSUBS 0.004963f
C209 B.n172 VSUBS 0.00888f
C210 B.n173 VSUBS 0.00888f
C211 B.n174 VSUBS 0.00888f
C212 B.n175 VSUBS 0.00888f
C213 B.n176 VSUBS 0.00888f
C214 B.n177 VSUBS 0.00888f
C215 B.n178 VSUBS 0.00888f
C216 B.n179 VSUBS 0.00888f
C217 B.n180 VSUBS 0.00888f
C218 B.n181 VSUBS 0.00888f
C219 B.n182 VSUBS 0.00888f
C220 B.n183 VSUBS 0.00888f
C221 B.n184 VSUBS 0.00888f
C222 B.n185 VSUBS 0.00888f
C223 B.n186 VSUBS 0.00888f
C224 B.n187 VSUBS 0.00888f
C225 B.n188 VSUBS 0.00888f
C226 B.n189 VSUBS 0.00888f
C227 B.n190 VSUBS 0.00888f
C228 B.n191 VSUBS 0.00888f
C229 B.n192 VSUBS 0.00888f
C230 B.n193 VSUBS 0.00888f
C231 B.n194 VSUBS 0.00888f
C232 B.n195 VSUBS 0.00888f
C233 B.n196 VSUBS 0.00888f
C234 B.n197 VSUBS 0.020502f
C235 B.n198 VSUBS 0.00888f
C236 B.n199 VSUBS 0.00888f
C237 B.n200 VSUBS 0.00888f
C238 B.n201 VSUBS 0.00888f
C239 B.n202 VSUBS 0.00888f
C240 B.n203 VSUBS 0.00888f
C241 B.n204 VSUBS 0.00888f
C242 B.n205 VSUBS 0.00888f
C243 B.n206 VSUBS 0.00888f
C244 B.n207 VSUBS 0.00888f
C245 B.n208 VSUBS 0.00888f
C246 B.n209 VSUBS 0.00888f
C247 B.n210 VSUBS 0.00888f
C248 B.n211 VSUBS 0.00888f
C249 B.n212 VSUBS 0.00888f
C250 B.n213 VSUBS 0.00888f
C251 B.n214 VSUBS 0.00888f
C252 B.n215 VSUBS 0.00888f
C253 B.n216 VSUBS 0.00888f
C254 B.n217 VSUBS 0.00888f
C255 B.n218 VSUBS 0.00888f
C256 B.n219 VSUBS 0.00888f
C257 B.n220 VSUBS 0.00888f
C258 B.n221 VSUBS 0.00888f
C259 B.n222 VSUBS 0.00888f
C260 B.n223 VSUBS 0.00888f
C261 B.n224 VSUBS 0.00888f
C262 B.n225 VSUBS 0.00888f
C263 B.n226 VSUBS 0.00888f
C264 B.n227 VSUBS 0.00888f
C265 B.n228 VSUBS 0.00888f
C266 B.n229 VSUBS 0.00888f
C267 B.n230 VSUBS 0.00888f
C268 B.n231 VSUBS 0.00888f
C269 B.n232 VSUBS 0.00888f
C270 B.n233 VSUBS 0.00888f
C271 B.n234 VSUBS 0.00888f
C272 B.n235 VSUBS 0.00888f
C273 B.n236 VSUBS 0.00888f
C274 B.n237 VSUBS 0.00888f
C275 B.n238 VSUBS 0.00888f
C276 B.n239 VSUBS 0.00888f
C277 B.n240 VSUBS 0.00888f
C278 B.n241 VSUBS 0.00888f
C279 B.n242 VSUBS 0.00888f
C280 B.n243 VSUBS 0.00888f
C281 B.n244 VSUBS 0.00888f
C282 B.n245 VSUBS 0.00888f
C283 B.n246 VSUBS 0.00888f
C284 B.n247 VSUBS 0.00888f
C285 B.n248 VSUBS 0.00888f
C286 B.n249 VSUBS 0.00888f
C287 B.n250 VSUBS 0.00888f
C288 B.n251 VSUBS 0.00888f
C289 B.n252 VSUBS 0.00888f
C290 B.n253 VSUBS 0.00888f
C291 B.n254 VSUBS 0.00888f
C292 B.n255 VSUBS 0.00888f
C293 B.n256 VSUBS 0.00888f
C294 B.n257 VSUBS 0.00888f
C295 B.n258 VSUBS 0.00888f
C296 B.n259 VSUBS 0.00888f
C297 B.n260 VSUBS 0.00888f
C298 B.n261 VSUBS 0.00888f
C299 B.n262 VSUBS 0.00888f
C300 B.n263 VSUBS 0.00888f
C301 B.n264 VSUBS 0.00888f
C302 B.n265 VSUBS 0.00888f
C303 B.n266 VSUBS 0.00888f
C304 B.n267 VSUBS 0.00888f
C305 B.n268 VSUBS 0.00888f
C306 B.n269 VSUBS 0.00888f
C307 B.n270 VSUBS 0.00888f
C308 B.n271 VSUBS 0.00888f
C309 B.n272 VSUBS 0.00888f
C310 B.n273 VSUBS 0.00888f
C311 B.n274 VSUBS 0.00888f
C312 B.n275 VSUBS 0.00888f
C313 B.n276 VSUBS 0.00888f
C314 B.n277 VSUBS 0.00888f
C315 B.n278 VSUBS 0.00888f
C316 B.n279 VSUBS 0.00888f
C317 B.n280 VSUBS 0.00888f
C318 B.n281 VSUBS 0.00888f
C319 B.n282 VSUBS 0.00888f
C320 B.n283 VSUBS 0.00888f
C321 B.n284 VSUBS 0.00888f
C322 B.n285 VSUBS 0.00888f
C323 B.n286 VSUBS 0.00888f
C324 B.n287 VSUBS 0.00888f
C325 B.n288 VSUBS 0.00888f
C326 B.n289 VSUBS 0.00888f
C327 B.n290 VSUBS 0.00888f
C328 B.n291 VSUBS 0.00888f
C329 B.n292 VSUBS 0.00888f
C330 B.n293 VSUBS 0.00888f
C331 B.n294 VSUBS 0.020502f
C332 B.n295 VSUBS 0.021289f
C333 B.n296 VSUBS 0.021289f
C334 B.n297 VSUBS 0.00888f
C335 B.n298 VSUBS 0.00888f
C336 B.n299 VSUBS 0.00888f
C337 B.n300 VSUBS 0.00888f
C338 B.n301 VSUBS 0.00888f
C339 B.n302 VSUBS 0.00888f
C340 B.n303 VSUBS 0.00888f
C341 B.n304 VSUBS 0.00888f
C342 B.n305 VSUBS 0.00888f
C343 B.n306 VSUBS 0.00888f
C344 B.n307 VSUBS 0.00888f
C345 B.n308 VSUBS 0.00888f
C346 B.n309 VSUBS 0.00888f
C347 B.n310 VSUBS 0.00888f
C348 B.n311 VSUBS 0.00888f
C349 B.n312 VSUBS 0.00888f
C350 B.n313 VSUBS 0.00888f
C351 B.n314 VSUBS 0.00888f
C352 B.n315 VSUBS 0.00888f
C353 B.n316 VSUBS 0.00888f
C354 B.n317 VSUBS 0.00888f
C355 B.n318 VSUBS 0.00888f
C356 B.n319 VSUBS 0.00888f
C357 B.n320 VSUBS 0.00888f
C358 B.n321 VSUBS 0.00888f
C359 B.n322 VSUBS 0.00888f
C360 B.n323 VSUBS 0.00888f
C361 B.n324 VSUBS 0.00888f
C362 B.n325 VSUBS 0.00888f
C363 B.n326 VSUBS 0.00888f
C364 B.n327 VSUBS 0.00888f
C365 B.n328 VSUBS 0.00888f
C366 B.n329 VSUBS 0.00888f
C367 B.n330 VSUBS 0.00888f
C368 B.n331 VSUBS 0.00888f
C369 B.n332 VSUBS 0.00888f
C370 B.n333 VSUBS 0.00888f
C371 B.n334 VSUBS 0.00888f
C372 B.n335 VSUBS 0.00888f
C373 B.n336 VSUBS 0.00888f
C374 B.n337 VSUBS 0.00888f
C375 B.n338 VSUBS 0.00888f
C376 B.n339 VSUBS 0.00888f
C377 B.n340 VSUBS 0.00888f
C378 B.n341 VSUBS 0.00888f
C379 B.n342 VSUBS 0.00888f
C380 B.n343 VSUBS 0.00888f
C381 B.n344 VSUBS 0.00888f
C382 B.n345 VSUBS 0.00888f
C383 B.n346 VSUBS 0.00888f
C384 B.n347 VSUBS 0.00888f
C385 B.n348 VSUBS 0.00888f
C386 B.n349 VSUBS 0.00888f
C387 B.n350 VSUBS 0.00888f
C388 B.n351 VSUBS 0.00888f
C389 B.n352 VSUBS 0.00888f
C390 B.n353 VSUBS 0.00888f
C391 B.n354 VSUBS 0.00888f
C392 B.n355 VSUBS 0.00888f
C393 B.n356 VSUBS 0.00888f
C394 B.n357 VSUBS 0.00888f
C395 B.n358 VSUBS 0.00888f
C396 B.n359 VSUBS 0.00888f
C397 B.n360 VSUBS 0.00888f
C398 B.n361 VSUBS 0.00888f
C399 B.n362 VSUBS 0.00888f
C400 B.n363 VSUBS 0.00888f
C401 B.n364 VSUBS 0.00888f
C402 B.n365 VSUBS 0.00888f
C403 B.n366 VSUBS 0.00888f
C404 B.n367 VSUBS 0.00888f
C405 B.n368 VSUBS 0.00888f
C406 B.n369 VSUBS 0.00888f
C407 B.t8 VSUBS 0.646789f
C408 B.t7 VSUBS 0.668935f
C409 B.t6 VSUBS 1.77045f
C410 B.n370 VSUBS 0.331708f
C411 B.n371 VSUBS 0.088528f
C412 B.n372 VSUBS 0.020575f
C413 B.n373 VSUBS 0.008358f
C414 B.n374 VSUBS 0.00888f
C415 B.n375 VSUBS 0.00888f
C416 B.n376 VSUBS 0.00888f
C417 B.n377 VSUBS 0.00888f
C418 B.n378 VSUBS 0.00888f
C419 B.n379 VSUBS 0.00888f
C420 B.n380 VSUBS 0.00888f
C421 B.n381 VSUBS 0.00888f
C422 B.n382 VSUBS 0.00888f
C423 B.n383 VSUBS 0.00888f
C424 B.n384 VSUBS 0.00888f
C425 B.n385 VSUBS 0.00888f
C426 B.n386 VSUBS 0.00888f
C427 B.n387 VSUBS 0.00888f
C428 B.n388 VSUBS 0.00888f
C429 B.n389 VSUBS 0.004963f
C430 B.n390 VSUBS 0.020575f
C431 B.n391 VSUBS 0.008358f
C432 B.n392 VSUBS 0.00888f
C433 B.n393 VSUBS 0.00888f
C434 B.n394 VSUBS 0.00888f
C435 B.n395 VSUBS 0.00888f
C436 B.n396 VSUBS 0.00888f
C437 B.n397 VSUBS 0.00888f
C438 B.n398 VSUBS 0.00888f
C439 B.n399 VSUBS 0.00888f
C440 B.n400 VSUBS 0.00888f
C441 B.n401 VSUBS 0.00888f
C442 B.n402 VSUBS 0.00888f
C443 B.n403 VSUBS 0.00888f
C444 B.n404 VSUBS 0.00888f
C445 B.n405 VSUBS 0.00888f
C446 B.n406 VSUBS 0.00888f
C447 B.n407 VSUBS 0.00888f
C448 B.n408 VSUBS 0.00888f
C449 B.n409 VSUBS 0.00888f
C450 B.n410 VSUBS 0.00888f
C451 B.n411 VSUBS 0.00888f
C452 B.n412 VSUBS 0.00888f
C453 B.n413 VSUBS 0.00888f
C454 B.n414 VSUBS 0.00888f
C455 B.n415 VSUBS 0.00888f
C456 B.n416 VSUBS 0.00888f
C457 B.n417 VSUBS 0.00888f
C458 B.n418 VSUBS 0.00888f
C459 B.n419 VSUBS 0.00888f
C460 B.n420 VSUBS 0.00888f
C461 B.n421 VSUBS 0.00888f
C462 B.n422 VSUBS 0.00888f
C463 B.n423 VSUBS 0.00888f
C464 B.n424 VSUBS 0.00888f
C465 B.n425 VSUBS 0.00888f
C466 B.n426 VSUBS 0.00888f
C467 B.n427 VSUBS 0.00888f
C468 B.n428 VSUBS 0.00888f
C469 B.n429 VSUBS 0.00888f
C470 B.n430 VSUBS 0.00888f
C471 B.n431 VSUBS 0.00888f
C472 B.n432 VSUBS 0.00888f
C473 B.n433 VSUBS 0.00888f
C474 B.n434 VSUBS 0.00888f
C475 B.n435 VSUBS 0.00888f
C476 B.n436 VSUBS 0.00888f
C477 B.n437 VSUBS 0.00888f
C478 B.n438 VSUBS 0.00888f
C479 B.n439 VSUBS 0.00888f
C480 B.n440 VSUBS 0.00888f
C481 B.n441 VSUBS 0.00888f
C482 B.n442 VSUBS 0.00888f
C483 B.n443 VSUBS 0.00888f
C484 B.n444 VSUBS 0.00888f
C485 B.n445 VSUBS 0.00888f
C486 B.n446 VSUBS 0.00888f
C487 B.n447 VSUBS 0.00888f
C488 B.n448 VSUBS 0.00888f
C489 B.n449 VSUBS 0.00888f
C490 B.n450 VSUBS 0.00888f
C491 B.n451 VSUBS 0.00888f
C492 B.n452 VSUBS 0.00888f
C493 B.n453 VSUBS 0.00888f
C494 B.n454 VSUBS 0.00888f
C495 B.n455 VSUBS 0.00888f
C496 B.n456 VSUBS 0.00888f
C497 B.n457 VSUBS 0.00888f
C498 B.n458 VSUBS 0.00888f
C499 B.n459 VSUBS 0.00888f
C500 B.n460 VSUBS 0.00888f
C501 B.n461 VSUBS 0.00888f
C502 B.n462 VSUBS 0.00888f
C503 B.n463 VSUBS 0.00888f
C504 B.n464 VSUBS 0.00888f
C505 B.n465 VSUBS 0.00888f
C506 B.n466 VSUBS 0.021289f
C507 B.n467 VSUBS 0.020502f
C508 B.n468 VSUBS 0.021542f
C509 B.n469 VSUBS 0.00888f
C510 B.n470 VSUBS 0.00888f
C511 B.n471 VSUBS 0.00888f
C512 B.n472 VSUBS 0.00888f
C513 B.n473 VSUBS 0.00888f
C514 B.n474 VSUBS 0.00888f
C515 B.n475 VSUBS 0.00888f
C516 B.n476 VSUBS 0.00888f
C517 B.n477 VSUBS 0.00888f
C518 B.n478 VSUBS 0.00888f
C519 B.n479 VSUBS 0.00888f
C520 B.n480 VSUBS 0.00888f
C521 B.n481 VSUBS 0.00888f
C522 B.n482 VSUBS 0.00888f
C523 B.n483 VSUBS 0.00888f
C524 B.n484 VSUBS 0.00888f
C525 B.n485 VSUBS 0.00888f
C526 B.n486 VSUBS 0.00888f
C527 B.n487 VSUBS 0.00888f
C528 B.n488 VSUBS 0.00888f
C529 B.n489 VSUBS 0.00888f
C530 B.n490 VSUBS 0.00888f
C531 B.n491 VSUBS 0.00888f
C532 B.n492 VSUBS 0.00888f
C533 B.n493 VSUBS 0.00888f
C534 B.n494 VSUBS 0.00888f
C535 B.n495 VSUBS 0.00888f
C536 B.n496 VSUBS 0.00888f
C537 B.n497 VSUBS 0.00888f
C538 B.n498 VSUBS 0.00888f
C539 B.n499 VSUBS 0.00888f
C540 B.n500 VSUBS 0.00888f
C541 B.n501 VSUBS 0.00888f
C542 B.n502 VSUBS 0.00888f
C543 B.n503 VSUBS 0.00888f
C544 B.n504 VSUBS 0.00888f
C545 B.n505 VSUBS 0.00888f
C546 B.n506 VSUBS 0.00888f
C547 B.n507 VSUBS 0.00888f
C548 B.n508 VSUBS 0.00888f
C549 B.n509 VSUBS 0.00888f
C550 B.n510 VSUBS 0.00888f
C551 B.n511 VSUBS 0.00888f
C552 B.n512 VSUBS 0.00888f
C553 B.n513 VSUBS 0.00888f
C554 B.n514 VSUBS 0.00888f
C555 B.n515 VSUBS 0.00888f
C556 B.n516 VSUBS 0.00888f
C557 B.n517 VSUBS 0.00888f
C558 B.n518 VSUBS 0.00888f
C559 B.n519 VSUBS 0.00888f
C560 B.n520 VSUBS 0.00888f
C561 B.n521 VSUBS 0.00888f
C562 B.n522 VSUBS 0.00888f
C563 B.n523 VSUBS 0.00888f
C564 B.n524 VSUBS 0.00888f
C565 B.n525 VSUBS 0.00888f
C566 B.n526 VSUBS 0.00888f
C567 B.n527 VSUBS 0.00888f
C568 B.n528 VSUBS 0.00888f
C569 B.n529 VSUBS 0.00888f
C570 B.n530 VSUBS 0.00888f
C571 B.n531 VSUBS 0.00888f
C572 B.n532 VSUBS 0.00888f
C573 B.n533 VSUBS 0.00888f
C574 B.n534 VSUBS 0.00888f
C575 B.n535 VSUBS 0.00888f
C576 B.n536 VSUBS 0.00888f
C577 B.n537 VSUBS 0.00888f
C578 B.n538 VSUBS 0.00888f
C579 B.n539 VSUBS 0.00888f
C580 B.n540 VSUBS 0.00888f
C581 B.n541 VSUBS 0.00888f
C582 B.n542 VSUBS 0.00888f
C583 B.n543 VSUBS 0.00888f
C584 B.n544 VSUBS 0.00888f
C585 B.n545 VSUBS 0.00888f
C586 B.n546 VSUBS 0.00888f
C587 B.n547 VSUBS 0.00888f
C588 B.n548 VSUBS 0.00888f
C589 B.n549 VSUBS 0.00888f
C590 B.n550 VSUBS 0.00888f
C591 B.n551 VSUBS 0.00888f
C592 B.n552 VSUBS 0.00888f
C593 B.n553 VSUBS 0.00888f
C594 B.n554 VSUBS 0.00888f
C595 B.n555 VSUBS 0.00888f
C596 B.n556 VSUBS 0.00888f
C597 B.n557 VSUBS 0.00888f
C598 B.n558 VSUBS 0.00888f
C599 B.n559 VSUBS 0.00888f
C600 B.n560 VSUBS 0.00888f
C601 B.n561 VSUBS 0.00888f
C602 B.n562 VSUBS 0.00888f
C603 B.n563 VSUBS 0.00888f
C604 B.n564 VSUBS 0.00888f
C605 B.n565 VSUBS 0.00888f
C606 B.n566 VSUBS 0.00888f
C607 B.n567 VSUBS 0.00888f
C608 B.n568 VSUBS 0.00888f
C609 B.n569 VSUBS 0.00888f
C610 B.n570 VSUBS 0.00888f
C611 B.n571 VSUBS 0.00888f
C612 B.n572 VSUBS 0.00888f
C613 B.n573 VSUBS 0.00888f
C614 B.n574 VSUBS 0.00888f
C615 B.n575 VSUBS 0.00888f
C616 B.n576 VSUBS 0.00888f
C617 B.n577 VSUBS 0.00888f
C618 B.n578 VSUBS 0.00888f
C619 B.n579 VSUBS 0.00888f
C620 B.n580 VSUBS 0.00888f
C621 B.n581 VSUBS 0.00888f
C622 B.n582 VSUBS 0.00888f
C623 B.n583 VSUBS 0.00888f
C624 B.n584 VSUBS 0.00888f
C625 B.n585 VSUBS 0.00888f
C626 B.n586 VSUBS 0.00888f
C627 B.n587 VSUBS 0.00888f
C628 B.n588 VSUBS 0.00888f
C629 B.n589 VSUBS 0.00888f
C630 B.n590 VSUBS 0.00888f
C631 B.n591 VSUBS 0.00888f
C632 B.n592 VSUBS 0.00888f
C633 B.n593 VSUBS 0.00888f
C634 B.n594 VSUBS 0.00888f
C635 B.n595 VSUBS 0.00888f
C636 B.n596 VSUBS 0.00888f
C637 B.n597 VSUBS 0.00888f
C638 B.n598 VSUBS 0.00888f
C639 B.n599 VSUBS 0.00888f
C640 B.n600 VSUBS 0.00888f
C641 B.n601 VSUBS 0.00888f
C642 B.n602 VSUBS 0.00888f
C643 B.n603 VSUBS 0.00888f
C644 B.n604 VSUBS 0.00888f
C645 B.n605 VSUBS 0.00888f
C646 B.n606 VSUBS 0.00888f
C647 B.n607 VSUBS 0.00888f
C648 B.n608 VSUBS 0.00888f
C649 B.n609 VSUBS 0.00888f
C650 B.n610 VSUBS 0.00888f
C651 B.n611 VSUBS 0.00888f
C652 B.n612 VSUBS 0.00888f
C653 B.n613 VSUBS 0.00888f
C654 B.n614 VSUBS 0.00888f
C655 B.n615 VSUBS 0.00888f
C656 B.n616 VSUBS 0.00888f
C657 B.n617 VSUBS 0.00888f
C658 B.n618 VSUBS 0.00888f
C659 B.n619 VSUBS 0.020502f
C660 B.n620 VSUBS 0.021289f
C661 B.n621 VSUBS 0.021289f
C662 B.n622 VSUBS 0.00888f
C663 B.n623 VSUBS 0.00888f
C664 B.n624 VSUBS 0.00888f
C665 B.n625 VSUBS 0.00888f
C666 B.n626 VSUBS 0.00888f
C667 B.n627 VSUBS 0.00888f
C668 B.n628 VSUBS 0.00888f
C669 B.n629 VSUBS 0.00888f
C670 B.n630 VSUBS 0.00888f
C671 B.n631 VSUBS 0.00888f
C672 B.n632 VSUBS 0.00888f
C673 B.n633 VSUBS 0.00888f
C674 B.n634 VSUBS 0.00888f
C675 B.n635 VSUBS 0.00888f
C676 B.n636 VSUBS 0.00888f
C677 B.n637 VSUBS 0.00888f
C678 B.n638 VSUBS 0.00888f
C679 B.n639 VSUBS 0.00888f
C680 B.n640 VSUBS 0.00888f
C681 B.n641 VSUBS 0.00888f
C682 B.n642 VSUBS 0.00888f
C683 B.n643 VSUBS 0.00888f
C684 B.n644 VSUBS 0.00888f
C685 B.n645 VSUBS 0.00888f
C686 B.n646 VSUBS 0.00888f
C687 B.n647 VSUBS 0.00888f
C688 B.n648 VSUBS 0.00888f
C689 B.n649 VSUBS 0.00888f
C690 B.n650 VSUBS 0.00888f
C691 B.n651 VSUBS 0.00888f
C692 B.n652 VSUBS 0.00888f
C693 B.n653 VSUBS 0.00888f
C694 B.n654 VSUBS 0.00888f
C695 B.n655 VSUBS 0.00888f
C696 B.n656 VSUBS 0.00888f
C697 B.n657 VSUBS 0.00888f
C698 B.n658 VSUBS 0.00888f
C699 B.n659 VSUBS 0.00888f
C700 B.n660 VSUBS 0.00888f
C701 B.n661 VSUBS 0.00888f
C702 B.n662 VSUBS 0.00888f
C703 B.n663 VSUBS 0.00888f
C704 B.n664 VSUBS 0.00888f
C705 B.n665 VSUBS 0.00888f
C706 B.n666 VSUBS 0.00888f
C707 B.n667 VSUBS 0.00888f
C708 B.n668 VSUBS 0.00888f
C709 B.n669 VSUBS 0.00888f
C710 B.n670 VSUBS 0.00888f
C711 B.n671 VSUBS 0.00888f
C712 B.n672 VSUBS 0.00888f
C713 B.n673 VSUBS 0.00888f
C714 B.n674 VSUBS 0.00888f
C715 B.n675 VSUBS 0.00888f
C716 B.n676 VSUBS 0.00888f
C717 B.n677 VSUBS 0.00888f
C718 B.n678 VSUBS 0.00888f
C719 B.n679 VSUBS 0.00888f
C720 B.n680 VSUBS 0.00888f
C721 B.n681 VSUBS 0.00888f
C722 B.n682 VSUBS 0.00888f
C723 B.n683 VSUBS 0.00888f
C724 B.n684 VSUBS 0.00888f
C725 B.n685 VSUBS 0.00888f
C726 B.n686 VSUBS 0.00888f
C727 B.n687 VSUBS 0.00888f
C728 B.n688 VSUBS 0.00888f
C729 B.n689 VSUBS 0.00888f
C730 B.n690 VSUBS 0.00888f
C731 B.n691 VSUBS 0.00888f
C732 B.n692 VSUBS 0.00888f
C733 B.n693 VSUBS 0.00888f
C734 B.n694 VSUBS 0.00888f
C735 B.n695 VSUBS 0.00888f
C736 B.n696 VSUBS 0.008358f
C737 B.n697 VSUBS 0.020575f
C738 B.n698 VSUBS 0.004963f
C739 B.n699 VSUBS 0.00888f
C740 B.n700 VSUBS 0.00888f
C741 B.n701 VSUBS 0.00888f
C742 B.n702 VSUBS 0.00888f
C743 B.n703 VSUBS 0.00888f
C744 B.n704 VSUBS 0.00888f
C745 B.n705 VSUBS 0.00888f
C746 B.n706 VSUBS 0.00888f
C747 B.n707 VSUBS 0.00888f
C748 B.n708 VSUBS 0.00888f
C749 B.n709 VSUBS 0.00888f
C750 B.n710 VSUBS 0.00888f
C751 B.n711 VSUBS 0.004963f
C752 B.n712 VSUBS 0.00888f
C753 B.n713 VSUBS 0.00888f
C754 B.n714 VSUBS 0.00888f
C755 B.n715 VSUBS 0.00888f
C756 B.n716 VSUBS 0.00888f
C757 B.n717 VSUBS 0.00888f
C758 B.n718 VSUBS 0.00888f
C759 B.n719 VSUBS 0.00888f
C760 B.n720 VSUBS 0.00888f
C761 B.n721 VSUBS 0.00888f
C762 B.n722 VSUBS 0.00888f
C763 B.n723 VSUBS 0.00888f
C764 B.n724 VSUBS 0.00888f
C765 B.n725 VSUBS 0.00888f
C766 B.n726 VSUBS 0.00888f
C767 B.n727 VSUBS 0.00888f
C768 B.n728 VSUBS 0.00888f
C769 B.n729 VSUBS 0.00888f
C770 B.n730 VSUBS 0.00888f
C771 B.n731 VSUBS 0.00888f
C772 B.n732 VSUBS 0.00888f
C773 B.n733 VSUBS 0.00888f
C774 B.n734 VSUBS 0.00888f
C775 B.n735 VSUBS 0.00888f
C776 B.n736 VSUBS 0.00888f
C777 B.n737 VSUBS 0.00888f
C778 B.n738 VSUBS 0.00888f
C779 B.n739 VSUBS 0.00888f
C780 B.n740 VSUBS 0.00888f
C781 B.n741 VSUBS 0.00888f
C782 B.n742 VSUBS 0.00888f
C783 B.n743 VSUBS 0.00888f
C784 B.n744 VSUBS 0.00888f
C785 B.n745 VSUBS 0.00888f
C786 B.n746 VSUBS 0.00888f
C787 B.n747 VSUBS 0.00888f
C788 B.n748 VSUBS 0.00888f
C789 B.n749 VSUBS 0.00888f
C790 B.n750 VSUBS 0.00888f
C791 B.n751 VSUBS 0.00888f
C792 B.n752 VSUBS 0.00888f
C793 B.n753 VSUBS 0.00888f
C794 B.n754 VSUBS 0.00888f
C795 B.n755 VSUBS 0.00888f
C796 B.n756 VSUBS 0.00888f
C797 B.n757 VSUBS 0.00888f
C798 B.n758 VSUBS 0.00888f
C799 B.n759 VSUBS 0.00888f
C800 B.n760 VSUBS 0.00888f
C801 B.n761 VSUBS 0.00888f
C802 B.n762 VSUBS 0.00888f
C803 B.n763 VSUBS 0.00888f
C804 B.n764 VSUBS 0.00888f
C805 B.n765 VSUBS 0.00888f
C806 B.n766 VSUBS 0.00888f
C807 B.n767 VSUBS 0.00888f
C808 B.n768 VSUBS 0.00888f
C809 B.n769 VSUBS 0.00888f
C810 B.n770 VSUBS 0.00888f
C811 B.n771 VSUBS 0.00888f
C812 B.n772 VSUBS 0.00888f
C813 B.n773 VSUBS 0.00888f
C814 B.n774 VSUBS 0.00888f
C815 B.n775 VSUBS 0.00888f
C816 B.n776 VSUBS 0.00888f
C817 B.n777 VSUBS 0.00888f
C818 B.n778 VSUBS 0.00888f
C819 B.n779 VSUBS 0.00888f
C820 B.n780 VSUBS 0.00888f
C821 B.n781 VSUBS 0.00888f
C822 B.n782 VSUBS 0.00888f
C823 B.n783 VSUBS 0.00888f
C824 B.n784 VSUBS 0.00888f
C825 B.n785 VSUBS 0.00888f
C826 B.n786 VSUBS 0.00888f
C827 B.n787 VSUBS 0.00888f
C828 B.n788 VSUBS 0.021289f
C829 B.n789 VSUBS 0.020502f
C830 B.n790 VSUBS 0.020502f
C831 B.n791 VSUBS 0.00888f
C832 B.n792 VSUBS 0.00888f
C833 B.n793 VSUBS 0.00888f
C834 B.n794 VSUBS 0.00888f
C835 B.n795 VSUBS 0.00888f
C836 B.n796 VSUBS 0.00888f
C837 B.n797 VSUBS 0.00888f
C838 B.n798 VSUBS 0.00888f
C839 B.n799 VSUBS 0.00888f
C840 B.n800 VSUBS 0.00888f
C841 B.n801 VSUBS 0.00888f
C842 B.n802 VSUBS 0.00888f
C843 B.n803 VSUBS 0.00888f
C844 B.n804 VSUBS 0.00888f
C845 B.n805 VSUBS 0.00888f
C846 B.n806 VSUBS 0.00888f
C847 B.n807 VSUBS 0.00888f
C848 B.n808 VSUBS 0.00888f
C849 B.n809 VSUBS 0.00888f
C850 B.n810 VSUBS 0.00888f
C851 B.n811 VSUBS 0.00888f
C852 B.n812 VSUBS 0.00888f
C853 B.n813 VSUBS 0.00888f
C854 B.n814 VSUBS 0.00888f
C855 B.n815 VSUBS 0.00888f
C856 B.n816 VSUBS 0.00888f
C857 B.n817 VSUBS 0.00888f
C858 B.n818 VSUBS 0.00888f
C859 B.n819 VSUBS 0.00888f
C860 B.n820 VSUBS 0.00888f
C861 B.n821 VSUBS 0.00888f
C862 B.n822 VSUBS 0.00888f
C863 B.n823 VSUBS 0.00888f
C864 B.n824 VSUBS 0.00888f
C865 B.n825 VSUBS 0.00888f
C866 B.n826 VSUBS 0.00888f
C867 B.n827 VSUBS 0.00888f
C868 B.n828 VSUBS 0.00888f
C869 B.n829 VSUBS 0.00888f
C870 B.n830 VSUBS 0.00888f
C871 B.n831 VSUBS 0.00888f
C872 B.n832 VSUBS 0.00888f
C873 B.n833 VSUBS 0.00888f
C874 B.n834 VSUBS 0.00888f
C875 B.n835 VSUBS 0.00888f
C876 B.n836 VSUBS 0.00888f
C877 B.n837 VSUBS 0.00888f
C878 B.n838 VSUBS 0.00888f
C879 B.n839 VSUBS 0.00888f
C880 B.n840 VSUBS 0.00888f
C881 B.n841 VSUBS 0.00888f
C882 B.n842 VSUBS 0.00888f
C883 B.n843 VSUBS 0.00888f
C884 B.n844 VSUBS 0.00888f
C885 B.n845 VSUBS 0.00888f
C886 B.n846 VSUBS 0.00888f
C887 B.n847 VSUBS 0.00888f
C888 B.n848 VSUBS 0.00888f
C889 B.n849 VSUBS 0.00888f
C890 B.n850 VSUBS 0.00888f
C891 B.n851 VSUBS 0.00888f
C892 B.n852 VSUBS 0.00888f
C893 B.n853 VSUBS 0.00888f
C894 B.n854 VSUBS 0.00888f
C895 B.n855 VSUBS 0.00888f
C896 B.n856 VSUBS 0.00888f
C897 B.n857 VSUBS 0.00888f
C898 B.n858 VSUBS 0.00888f
C899 B.n859 VSUBS 0.00888f
C900 B.n860 VSUBS 0.00888f
C901 B.n861 VSUBS 0.00888f
C902 B.n862 VSUBS 0.00888f
C903 B.n863 VSUBS 0.011588f
C904 B.n864 VSUBS 0.012345f
C905 B.n865 VSUBS 0.024549f
C906 VDD2.t1 VSUBS 3.44855f
C907 VDD2.t2 VSUBS 0.325702f
C908 VDD2.t0 VSUBS 0.325702f
C909 VDD2.n0 VSUBS 2.63212f
C910 VDD2.n1 VSUBS 1.55474f
C911 VDD2.t6 VSUBS 0.325702f
C912 VDD2.t8 VSUBS 0.325702f
C913 VDD2.n2 VSUBS 2.65019f
C914 VDD2.n3 VSUBS 3.36208f
C915 VDD2.t9 VSUBS 3.42549f
C916 VDD2.n4 VSUBS 3.75615f
C917 VDD2.t7 VSUBS 0.325702f
C918 VDD2.t3 VSUBS 0.325702f
C919 VDD2.n5 VSUBS 2.63212f
C920 VDD2.n6 VSUBS 0.765257f
C921 VDD2.t4 VSUBS 0.325702f
C922 VDD2.t5 VSUBS 0.325702f
C923 VDD2.n7 VSUBS 2.65015f
C924 VN.n0 VSUBS 0.039543f
C925 VN.t1 VSUBS 2.60235f
C926 VN.n1 VSUBS 0.028334f
C927 VN.n2 VSUBS 0.029993f
C928 VN.t3 VSUBS 2.60235f
C929 VN.n3 VSUBS 0.047963f
C930 VN.n4 VSUBS 0.029993f
C931 VN.t9 VSUBS 2.60235f
C932 VN.n5 VSUBS 0.055899f
C933 VN.n6 VSUBS 0.029993f
C934 VN.t7 VSUBS 2.60235f
C935 VN.n7 VSUBS 0.997037f
C936 VN.t8 VSUBS 2.76929f
C937 VN.n8 VSUBS 0.983101f
C938 VN.n9 VSUBS 0.251537f
C939 VN.n10 VSUBS 0.05038f
C940 VN.n11 VSUBS 0.047963f
C941 VN.n12 VSUBS 0.039605f
C942 VN.n13 VSUBS 0.029993f
C943 VN.n14 VSUBS 0.029993f
C944 VN.n15 VSUBS 0.029993f
C945 VN.n16 VSUBS 0.942682f
C946 VN.n17 VSUBS 0.055899f
C947 VN.n18 VSUBS 0.039605f
C948 VN.n19 VSUBS 0.029993f
C949 VN.n20 VSUBS 0.029993f
C950 VN.n21 VSUBS 0.029993f
C951 VN.n22 VSUBS 0.05038f
C952 VN.n23 VSUBS 0.91438f
C953 VN.n24 VSUBS 0.033821f
C954 VN.n25 VSUBS 0.060086f
C955 VN.n26 VSUBS 0.029993f
C956 VN.n27 VSUBS 0.029993f
C957 VN.n28 VSUBS 0.029993f
C958 VN.n29 VSUBS 0.055048f
C959 VN.n30 VSUBS 0.04486f
C960 VN.n31 VSUBS 1.00062f
C961 VN.n32 VSUBS 0.04087f
C962 VN.n33 VSUBS 0.039543f
C963 VN.t0 VSUBS 2.60235f
C964 VN.n34 VSUBS 0.028334f
C965 VN.n35 VSUBS 0.029993f
C966 VN.t2 VSUBS 2.60235f
C967 VN.n36 VSUBS 0.047963f
C968 VN.n37 VSUBS 0.029993f
C969 VN.t6 VSUBS 2.60235f
C970 VN.n38 VSUBS 0.055899f
C971 VN.n39 VSUBS 0.029993f
C972 VN.t5 VSUBS 2.60235f
C973 VN.n40 VSUBS 0.997037f
C974 VN.t4 VSUBS 2.76929f
C975 VN.n41 VSUBS 0.983101f
C976 VN.n42 VSUBS 0.251537f
C977 VN.n43 VSUBS 0.05038f
C978 VN.n44 VSUBS 0.047963f
C979 VN.n45 VSUBS 0.039605f
C980 VN.n46 VSUBS 0.029993f
C981 VN.n47 VSUBS 0.029993f
C982 VN.n48 VSUBS 0.029993f
C983 VN.n49 VSUBS 0.942682f
C984 VN.n50 VSUBS 0.055899f
C985 VN.n51 VSUBS 0.039605f
C986 VN.n52 VSUBS 0.029993f
C987 VN.n53 VSUBS 0.029993f
C988 VN.n54 VSUBS 0.029993f
C989 VN.n55 VSUBS 0.05038f
C990 VN.n56 VSUBS 0.91438f
C991 VN.n57 VSUBS 0.033821f
C992 VN.n58 VSUBS 0.060086f
C993 VN.n59 VSUBS 0.029993f
C994 VN.n60 VSUBS 0.029993f
C995 VN.n61 VSUBS 0.029993f
C996 VN.n62 VSUBS 0.055048f
C997 VN.n63 VSUBS 0.04486f
C998 VN.n64 VSUBS 1.00062f
C999 VN.n65 VSUBS 1.80732f
C1000 VDD1.t3 VSUBS 3.43735f
C1001 VDD1.t5 VSUBS 0.324642f
C1002 VDD1.t4 VSUBS 0.324642f
C1003 VDD1.n0 VSUBS 2.62356f
C1004 VDD1.n1 VSUBS 1.55814f
C1005 VDD1.t2 VSUBS 3.43733f
C1006 VDD1.t1 VSUBS 0.324642f
C1007 VDD1.t0 VSUBS 0.324642f
C1008 VDD1.n2 VSUBS 2.62355f
C1009 VDD1.n3 VSUBS 1.54968f
C1010 VDD1.t7 VSUBS 0.324642f
C1011 VDD1.t8 VSUBS 0.324642f
C1012 VDD1.n4 VSUBS 2.64156f
C1013 VDD1.n5 VSUBS 3.47246f
C1014 VDD1.t6 VSUBS 0.324642f
C1015 VDD1.t9 VSUBS 0.324642f
C1016 VDD1.n6 VSUBS 2.62356f
C1017 VDD1.n7 VSUBS 3.75655f
C1018 VTAIL.t3 VSUBS 0.333965f
C1019 VTAIL.t0 VSUBS 0.333965f
C1020 VTAIL.n0 VSUBS 2.52693f
C1021 VTAIL.n1 VSUBS 0.96092f
C1022 VTAIL.t11 VSUBS 3.31751f
C1023 VTAIL.n2 VSUBS 1.12204f
C1024 VTAIL.t14 VSUBS 0.333965f
C1025 VTAIL.t12 VSUBS 0.333965f
C1026 VTAIL.n3 VSUBS 2.52693f
C1027 VTAIL.n4 VSUBS 1.05209f
C1028 VTAIL.t19 VSUBS 0.333965f
C1029 VTAIL.t15 VSUBS 0.333965f
C1030 VTAIL.n5 VSUBS 2.52693f
C1031 VTAIL.n6 VSUBS 2.78576f
C1032 VTAIL.t5 VSUBS 0.333965f
C1033 VTAIL.t1 VSUBS 0.333965f
C1034 VTAIL.n7 VSUBS 2.52694f
C1035 VTAIL.n8 VSUBS 2.78575f
C1036 VTAIL.t7 VSUBS 0.333965f
C1037 VTAIL.t9 VSUBS 0.333965f
C1038 VTAIL.n9 VSUBS 2.52694f
C1039 VTAIL.n10 VSUBS 1.05208f
C1040 VTAIL.t4 VSUBS 3.31753f
C1041 VTAIL.n11 VSUBS 1.12202f
C1042 VTAIL.t18 VSUBS 0.333965f
C1043 VTAIL.t13 VSUBS 0.333965f
C1044 VTAIL.n12 VSUBS 2.52694f
C1045 VTAIL.n13 VSUBS 1.00179f
C1046 VTAIL.t17 VSUBS 0.333965f
C1047 VTAIL.t16 VSUBS 0.333965f
C1048 VTAIL.n14 VSUBS 2.52694f
C1049 VTAIL.n15 VSUBS 1.05208f
C1050 VTAIL.t10 VSUBS 3.31752f
C1051 VTAIL.n16 VSUBS 2.72171f
C1052 VTAIL.t8 VSUBS 3.31751f
C1053 VTAIL.n17 VSUBS 2.72173f
C1054 VTAIL.t6 VSUBS 0.333965f
C1055 VTAIL.t2 VSUBS 0.333965f
C1056 VTAIL.n18 VSUBS 2.52693f
C1057 VTAIL.n19 VSUBS 0.908711f
C1058 VP.n0 VSUBS 0.042209f
C1059 VP.t1 VSUBS 2.77779f
C1060 VP.n1 VSUBS 0.030244f
C1061 VP.n2 VSUBS 0.032015f
C1062 VP.t2 VSUBS 2.77779f
C1063 VP.n3 VSUBS 0.051197f
C1064 VP.n4 VSUBS 0.032015f
C1065 VP.t9 VSUBS 2.77779f
C1066 VP.n5 VSUBS 0.059668f
C1067 VP.n6 VSUBS 0.032015f
C1068 VP.t8 VSUBS 2.77779f
C1069 VP.n7 VSUBS 0.976025f
C1070 VP.n8 VSUBS 0.032015f
C1071 VP.n9 VSUBS 0.058759f
C1072 VP.n10 VSUBS 0.042209f
C1073 VP.t0 VSUBS 2.77779f
C1074 VP.n11 VSUBS 0.030244f
C1075 VP.n12 VSUBS 0.032015f
C1076 VP.t3 VSUBS 2.77779f
C1077 VP.n13 VSUBS 0.051197f
C1078 VP.n14 VSUBS 0.032015f
C1079 VP.t5 VSUBS 2.77779f
C1080 VP.n15 VSUBS 0.059668f
C1081 VP.n16 VSUBS 0.032015f
C1082 VP.t4 VSUBS 2.77779f
C1083 VP.n17 VSUBS 1.06425f
C1084 VP.t6 VSUBS 2.95599f
C1085 VP.n18 VSUBS 1.04938f
C1086 VP.n19 VSUBS 0.268495f
C1087 VP.n20 VSUBS 0.053776f
C1088 VP.n21 VSUBS 0.051197f
C1089 VP.n22 VSUBS 0.042275f
C1090 VP.n23 VSUBS 0.032015f
C1091 VP.n24 VSUBS 0.032015f
C1092 VP.n25 VSUBS 0.032015f
C1093 VP.n26 VSUBS 1.00623f
C1094 VP.n27 VSUBS 0.059668f
C1095 VP.n28 VSUBS 0.042275f
C1096 VP.n29 VSUBS 0.032015f
C1097 VP.n30 VSUBS 0.032015f
C1098 VP.n31 VSUBS 0.032015f
C1099 VP.n32 VSUBS 0.053776f
C1100 VP.n33 VSUBS 0.976025f
C1101 VP.n34 VSUBS 0.036101f
C1102 VP.n35 VSUBS 0.064137f
C1103 VP.n36 VSUBS 0.032015f
C1104 VP.n37 VSUBS 0.032015f
C1105 VP.n38 VSUBS 0.032015f
C1106 VP.n39 VSUBS 0.058759f
C1107 VP.n40 VSUBS 0.047885f
C1108 VP.n41 VSUBS 1.06808f
C1109 VP.n42 VSUBS 1.91209f
C1110 VP.n43 VSUBS 1.93394f
C1111 VP.t7 VSUBS 2.77779f
C1112 VP.n44 VSUBS 1.06808f
C1113 VP.n45 VSUBS 0.047885f
C1114 VP.n46 VSUBS 0.042209f
C1115 VP.n47 VSUBS 0.032015f
C1116 VP.n48 VSUBS 0.032015f
C1117 VP.n49 VSUBS 0.030244f
C1118 VP.n50 VSUBS 0.064137f
C1119 VP.n51 VSUBS 0.036101f
C1120 VP.n52 VSUBS 0.032015f
C1121 VP.n53 VSUBS 0.032015f
C1122 VP.n54 VSUBS 0.053776f
C1123 VP.n55 VSUBS 0.051197f
C1124 VP.n56 VSUBS 0.042275f
C1125 VP.n57 VSUBS 0.032015f
C1126 VP.n58 VSUBS 0.032015f
C1127 VP.n59 VSUBS 0.032015f
C1128 VP.n60 VSUBS 1.00623f
C1129 VP.n61 VSUBS 0.059668f
C1130 VP.n62 VSUBS 0.042275f
C1131 VP.n63 VSUBS 0.032015f
C1132 VP.n64 VSUBS 0.032015f
C1133 VP.n65 VSUBS 0.032015f
C1134 VP.n66 VSUBS 0.053776f
C1135 VP.n67 VSUBS 0.976025f
C1136 VP.n68 VSUBS 0.036101f
C1137 VP.n69 VSUBS 0.064137f
C1138 VP.n70 VSUBS 0.032015f
C1139 VP.n71 VSUBS 0.032015f
C1140 VP.n72 VSUBS 0.032015f
C1141 VP.n73 VSUBS 0.058759f
C1142 VP.n74 VSUBS 0.047885f
C1143 VP.n75 VSUBS 1.06808f
C1144 VP.n76 VSUBS 0.043626f
.ends

