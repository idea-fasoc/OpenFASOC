* NGSPICE file created from diff_pair_sample_1773.ext - technology: sky130A

.subckt diff_pair_sample_1773 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=0 ps=0 w=13.53 l=2.4
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=5.2767 ps=27.84 w=13.53 l=2.4
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=0 ps=0 w=13.53 l=2.4
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=5.2767 ps=27.84 w=13.53 l=2.4
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=0 ps=0 w=13.53 l=2.4
X5 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=5.2767 ps=27.84 w=13.53 l=2.4
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=5.2767 ps=27.84 w=13.53 l=2.4
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2767 pd=27.84 as=0 ps=0 w=13.53 l=2.4
R0 B.n714 B.n713 585
R1 B.n303 B.n98 585
R2 B.n302 B.n301 585
R3 B.n300 B.n299 585
R4 B.n298 B.n297 585
R5 B.n296 B.n295 585
R6 B.n294 B.n293 585
R7 B.n292 B.n291 585
R8 B.n290 B.n289 585
R9 B.n288 B.n287 585
R10 B.n286 B.n285 585
R11 B.n284 B.n283 585
R12 B.n282 B.n281 585
R13 B.n280 B.n279 585
R14 B.n278 B.n277 585
R15 B.n276 B.n275 585
R16 B.n274 B.n273 585
R17 B.n272 B.n271 585
R18 B.n270 B.n269 585
R19 B.n268 B.n267 585
R20 B.n266 B.n265 585
R21 B.n264 B.n263 585
R22 B.n262 B.n261 585
R23 B.n260 B.n259 585
R24 B.n258 B.n257 585
R25 B.n256 B.n255 585
R26 B.n254 B.n253 585
R27 B.n252 B.n251 585
R28 B.n250 B.n249 585
R29 B.n248 B.n247 585
R30 B.n246 B.n245 585
R31 B.n244 B.n243 585
R32 B.n242 B.n241 585
R33 B.n240 B.n239 585
R34 B.n238 B.n237 585
R35 B.n236 B.n235 585
R36 B.n234 B.n233 585
R37 B.n232 B.n231 585
R38 B.n230 B.n229 585
R39 B.n228 B.n227 585
R40 B.n226 B.n225 585
R41 B.n224 B.n223 585
R42 B.n222 B.n221 585
R43 B.n220 B.n219 585
R44 B.n218 B.n217 585
R45 B.n216 B.n215 585
R46 B.n214 B.n213 585
R47 B.n212 B.n211 585
R48 B.n210 B.n209 585
R49 B.n208 B.n207 585
R50 B.n206 B.n205 585
R51 B.n204 B.n203 585
R52 B.n202 B.n201 585
R53 B.n200 B.n199 585
R54 B.n198 B.n197 585
R55 B.n196 B.n195 585
R56 B.n194 B.n193 585
R57 B.n192 B.n191 585
R58 B.n190 B.n189 585
R59 B.n188 B.n187 585
R60 B.n186 B.n185 585
R61 B.n184 B.n183 585
R62 B.n182 B.n181 585
R63 B.n180 B.n179 585
R64 B.n178 B.n177 585
R65 B.n176 B.n175 585
R66 B.n174 B.n173 585
R67 B.n172 B.n171 585
R68 B.n170 B.n169 585
R69 B.n168 B.n167 585
R70 B.n166 B.n165 585
R71 B.n164 B.n163 585
R72 B.n162 B.n161 585
R73 B.n160 B.n159 585
R74 B.n158 B.n157 585
R75 B.n156 B.n155 585
R76 B.n154 B.n153 585
R77 B.n152 B.n151 585
R78 B.n150 B.n149 585
R79 B.n148 B.n147 585
R80 B.n146 B.n145 585
R81 B.n144 B.n143 585
R82 B.n142 B.n141 585
R83 B.n140 B.n139 585
R84 B.n138 B.n137 585
R85 B.n136 B.n135 585
R86 B.n134 B.n133 585
R87 B.n132 B.n131 585
R88 B.n130 B.n129 585
R89 B.n128 B.n127 585
R90 B.n126 B.n125 585
R91 B.n124 B.n123 585
R92 B.n122 B.n121 585
R93 B.n120 B.n119 585
R94 B.n118 B.n117 585
R95 B.n116 B.n115 585
R96 B.n114 B.n113 585
R97 B.n112 B.n111 585
R98 B.n110 B.n109 585
R99 B.n108 B.n107 585
R100 B.n106 B.n105 585
R101 B.n46 B.n45 585
R102 B.n712 B.n47 585
R103 B.n717 B.n47 585
R104 B.n711 B.n710 585
R105 B.n710 B.n43 585
R106 B.n709 B.n42 585
R107 B.n723 B.n42 585
R108 B.n708 B.n41 585
R109 B.n724 B.n41 585
R110 B.n707 B.n40 585
R111 B.n725 B.n40 585
R112 B.n706 B.n705 585
R113 B.n705 B.n36 585
R114 B.n704 B.n35 585
R115 B.n731 B.n35 585
R116 B.n703 B.n34 585
R117 B.n732 B.n34 585
R118 B.n702 B.n33 585
R119 B.n733 B.n33 585
R120 B.n701 B.n700 585
R121 B.n700 B.n29 585
R122 B.n699 B.n28 585
R123 B.n739 B.n28 585
R124 B.n698 B.n27 585
R125 B.n740 B.n27 585
R126 B.n697 B.n26 585
R127 B.n741 B.n26 585
R128 B.n696 B.n695 585
R129 B.n695 B.n22 585
R130 B.n694 B.n21 585
R131 B.n747 B.n21 585
R132 B.n693 B.n20 585
R133 B.n748 B.n20 585
R134 B.n692 B.n19 585
R135 B.n749 B.n19 585
R136 B.n691 B.n690 585
R137 B.n690 B.n15 585
R138 B.n689 B.n14 585
R139 B.n755 B.n14 585
R140 B.n688 B.n13 585
R141 B.n756 B.n13 585
R142 B.n687 B.n12 585
R143 B.n757 B.n12 585
R144 B.n686 B.n685 585
R145 B.n685 B.n8 585
R146 B.n684 B.n7 585
R147 B.n763 B.n7 585
R148 B.n683 B.n6 585
R149 B.n764 B.n6 585
R150 B.n682 B.n5 585
R151 B.n765 B.n5 585
R152 B.n681 B.n680 585
R153 B.n680 B.n4 585
R154 B.n679 B.n304 585
R155 B.n679 B.n678 585
R156 B.n669 B.n305 585
R157 B.n306 B.n305 585
R158 B.n671 B.n670 585
R159 B.n672 B.n671 585
R160 B.n668 B.n311 585
R161 B.n311 B.n310 585
R162 B.n667 B.n666 585
R163 B.n666 B.n665 585
R164 B.n313 B.n312 585
R165 B.n314 B.n313 585
R166 B.n658 B.n657 585
R167 B.n659 B.n658 585
R168 B.n656 B.n319 585
R169 B.n319 B.n318 585
R170 B.n655 B.n654 585
R171 B.n654 B.n653 585
R172 B.n321 B.n320 585
R173 B.n322 B.n321 585
R174 B.n646 B.n645 585
R175 B.n647 B.n646 585
R176 B.n644 B.n327 585
R177 B.n327 B.n326 585
R178 B.n643 B.n642 585
R179 B.n642 B.n641 585
R180 B.n329 B.n328 585
R181 B.n330 B.n329 585
R182 B.n634 B.n633 585
R183 B.n635 B.n634 585
R184 B.n632 B.n334 585
R185 B.n338 B.n334 585
R186 B.n631 B.n630 585
R187 B.n630 B.n629 585
R188 B.n336 B.n335 585
R189 B.n337 B.n336 585
R190 B.n622 B.n621 585
R191 B.n623 B.n622 585
R192 B.n620 B.n343 585
R193 B.n343 B.n342 585
R194 B.n619 B.n618 585
R195 B.n618 B.n617 585
R196 B.n345 B.n344 585
R197 B.n346 B.n345 585
R198 B.n610 B.n609 585
R199 B.n611 B.n610 585
R200 B.n349 B.n348 585
R201 B.n406 B.n404 585
R202 B.n407 B.n403 585
R203 B.n407 B.n350 585
R204 B.n410 B.n409 585
R205 B.n411 B.n402 585
R206 B.n413 B.n412 585
R207 B.n415 B.n401 585
R208 B.n418 B.n417 585
R209 B.n419 B.n400 585
R210 B.n421 B.n420 585
R211 B.n423 B.n399 585
R212 B.n426 B.n425 585
R213 B.n427 B.n398 585
R214 B.n429 B.n428 585
R215 B.n431 B.n397 585
R216 B.n434 B.n433 585
R217 B.n435 B.n396 585
R218 B.n437 B.n436 585
R219 B.n439 B.n395 585
R220 B.n442 B.n441 585
R221 B.n443 B.n394 585
R222 B.n445 B.n444 585
R223 B.n447 B.n393 585
R224 B.n450 B.n449 585
R225 B.n451 B.n392 585
R226 B.n453 B.n452 585
R227 B.n455 B.n391 585
R228 B.n458 B.n457 585
R229 B.n459 B.n390 585
R230 B.n461 B.n460 585
R231 B.n463 B.n389 585
R232 B.n466 B.n465 585
R233 B.n467 B.n388 585
R234 B.n469 B.n468 585
R235 B.n471 B.n387 585
R236 B.n474 B.n473 585
R237 B.n475 B.n386 585
R238 B.n477 B.n476 585
R239 B.n479 B.n385 585
R240 B.n482 B.n481 585
R241 B.n483 B.n384 585
R242 B.n485 B.n484 585
R243 B.n487 B.n383 585
R244 B.n490 B.n489 585
R245 B.n491 B.n382 585
R246 B.n496 B.n495 585
R247 B.n498 B.n381 585
R248 B.n501 B.n500 585
R249 B.n502 B.n380 585
R250 B.n504 B.n503 585
R251 B.n506 B.n379 585
R252 B.n509 B.n508 585
R253 B.n510 B.n378 585
R254 B.n512 B.n511 585
R255 B.n514 B.n377 585
R256 B.n517 B.n516 585
R257 B.n519 B.n374 585
R258 B.n521 B.n520 585
R259 B.n523 B.n373 585
R260 B.n526 B.n525 585
R261 B.n527 B.n372 585
R262 B.n529 B.n528 585
R263 B.n531 B.n371 585
R264 B.n534 B.n533 585
R265 B.n535 B.n370 585
R266 B.n537 B.n536 585
R267 B.n539 B.n369 585
R268 B.n542 B.n541 585
R269 B.n543 B.n368 585
R270 B.n545 B.n544 585
R271 B.n547 B.n367 585
R272 B.n550 B.n549 585
R273 B.n551 B.n366 585
R274 B.n553 B.n552 585
R275 B.n555 B.n365 585
R276 B.n558 B.n557 585
R277 B.n559 B.n364 585
R278 B.n561 B.n560 585
R279 B.n563 B.n363 585
R280 B.n566 B.n565 585
R281 B.n567 B.n362 585
R282 B.n569 B.n568 585
R283 B.n571 B.n361 585
R284 B.n574 B.n573 585
R285 B.n575 B.n360 585
R286 B.n577 B.n576 585
R287 B.n579 B.n359 585
R288 B.n582 B.n581 585
R289 B.n583 B.n358 585
R290 B.n585 B.n584 585
R291 B.n587 B.n357 585
R292 B.n590 B.n589 585
R293 B.n591 B.n356 585
R294 B.n593 B.n592 585
R295 B.n595 B.n355 585
R296 B.n598 B.n597 585
R297 B.n599 B.n354 585
R298 B.n601 B.n600 585
R299 B.n603 B.n353 585
R300 B.n604 B.n352 585
R301 B.n607 B.n606 585
R302 B.n608 B.n351 585
R303 B.n351 B.n350 585
R304 B.n613 B.n612 585
R305 B.n612 B.n611 585
R306 B.n614 B.n347 585
R307 B.n347 B.n346 585
R308 B.n616 B.n615 585
R309 B.n617 B.n616 585
R310 B.n341 B.n340 585
R311 B.n342 B.n341 585
R312 B.n625 B.n624 585
R313 B.n624 B.n623 585
R314 B.n626 B.n339 585
R315 B.n339 B.n337 585
R316 B.n628 B.n627 585
R317 B.n629 B.n628 585
R318 B.n333 B.n332 585
R319 B.n338 B.n333 585
R320 B.n637 B.n636 585
R321 B.n636 B.n635 585
R322 B.n638 B.n331 585
R323 B.n331 B.n330 585
R324 B.n640 B.n639 585
R325 B.n641 B.n640 585
R326 B.n325 B.n324 585
R327 B.n326 B.n325 585
R328 B.n649 B.n648 585
R329 B.n648 B.n647 585
R330 B.n650 B.n323 585
R331 B.n323 B.n322 585
R332 B.n652 B.n651 585
R333 B.n653 B.n652 585
R334 B.n317 B.n316 585
R335 B.n318 B.n317 585
R336 B.n661 B.n660 585
R337 B.n660 B.n659 585
R338 B.n662 B.n315 585
R339 B.n315 B.n314 585
R340 B.n664 B.n663 585
R341 B.n665 B.n664 585
R342 B.n309 B.n308 585
R343 B.n310 B.n309 585
R344 B.n674 B.n673 585
R345 B.n673 B.n672 585
R346 B.n675 B.n307 585
R347 B.n307 B.n306 585
R348 B.n677 B.n676 585
R349 B.n678 B.n677 585
R350 B.n2 B.n0 585
R351 B.n4 B.n2 585
R352 B.n3 B.n1 585
R353 B.n764 B.n3 585
R354 B.n762 B.n761 585
R355 B.n763 B.n762 585
R356 B.n760 B.n9 585
R357 B.n9 B.n8 585
R358 B.n759 B.n758 585
R359 B.n758 B.n757 585
R360 B.n11 B.n10 585
R361 B.n756 B.n11 585
R362 B.n754 B.n753 585
R363 B.n755 B.n754 585
R364 B.n752 B.n16 585
R365 B.n16 B.n15 585
R366 B.n751 B.n750 585
R367 B.n750 B.n749 585
R368 B.n18 B.n17 585
R369 B.n748 B.n18 585
R370 B.n746 B.n745 585
R371 B.n747 B.n746 585
R372 B.n744 B.n23 585
R373 B.n23 B.n22 585
R374 B.n743 B.n742 585
R375 B.n742 B.n741 585
R376 B.n25 B.n24 585
R377 B.n740 B.n25 585
R378 B.n738 B.n737 585
R379 B.n739 B.n738 585
R380 B.n736 B.n30 585
R381 B.n30 B.n29 585
R382 B.n735 B.n734 585
R383 B.n734 B.n733 585
R384 B.n32 B.n31 585
R385 B.n732 B.n32 585
R386 B.n730 B.n729 585
R387 B.n731 B.n730 585
R388 B.n728 B.n37 585
R389 B.n37 B.n36 585
R390 B.n727 B.n726 585
R391 B.n726 B.n725 585
R392 B.n39 B.n38 585
R393 B.n724 B.n39 585
R394 B.n722 B.n721 585
R395 B.n723 B.n722 585
R396 B.n720 B.n44 585
R397 B.n44 B.n43 585
R398 B.n719 B.n718 585
R399 B.n718 B.n717 585
R400 B.n767 B.n766 585
R401 B.n766 B.n765 585
R402 B.n612 B.n349 511.721
R403 B.n718 B.n46 511.721
R404 B.n610 B.n351 511.721
R405 B.n714 B.n47 511.721
R406 B.n375 B.t12 361.675
R407 B.n99 B.t14 361.675
R408 B.n492 B.t5 361.675
R409 B.n102 B.t8 361.675
R410 B.n375 B.t10 343.587
R411 B.n492 B.t2 343.587
R412 B.n102 B.t6 343.587
R413 B.n99 B.t13 343.587
R414 B.n376 B.t11 308.729
R415 B.n100 B.t15 308.729
R416 B.n493 B.t4 308.729
R417 B.n103 B.t9 308.729
R418 B.n716 B.n715 256.663
R419 B.n716 B.n97 256.663
R420 B.n716 B.n96 256.663
R421 B.n716 B.n95 256.663
R422 B.n716 B.n94 256.663
R423 B.n716 B.n93 256.663
R424 B.n716 B.n92 256.663
R425 B.n716 B.n91 256.663
R426 B.n716 B.n90 256.663
R427 B.n716 B.n89 256.663
R428 B.n716 B.n88 256.663
R429 B.n716 B.n87 256.663
R430 B.n716 B.n86 256.663
R431 B.n716 B.n85 256.663
R432 B.n716 B.n84 256.663
R433 B.n716 B.n83 256.663
R434 B.n716 B.n82 256.663
R435 B.n716 B.n81 256.663
R436 B.n716 B.n80 256.663
R437 B.n716 B.n79 256.663
R438 B.n716 B.n78 256.663
R439 B.n716 B.n77 256.663
R440 B.n716 B.n76 256.663
R441 B.n716 B.n75 256.663
R442 B.n716 B.n74 256.663
R443 B.n716 B.n73 256.663
R444 B.n716 B.n72 256.663
R445 B.n716 B.n71 256.663
R446 B.n716 B.n70 256.663
R447 B.n716 B.n69 256.663
R448 B.n716 B.n68 256.663
R449 B.n716 B.n67 256.663
R450 B.n716 B.n66 256.663
R451 B.n716 B.n65 256.663
R452 B.n716 B.n64 256.663
R453 B.n716 B.n63 256.663
R454 B.n716 B.n62 256.663
R455 B.n716 B.n61 256.663
R456 B.n716 B.n60 256.663
R457 B.n716 B.n59 256.663
R458 B.n716 B.n58 256.663
R459 B.n716 B.n57 256.663
R460 B.n716 B.n56 256.663
R461 B.n716 B.n55 256.663
R462 B.n716 B.n54 256.663
R463 B.n716 B.n53 256.663
R464 B.n716 B.n52 256.663
R465 B.n716 B.n51 256.663
R466 B.n716 B.n50 256.663
R467 B.n716 B.n49 256.663
R468 B.n716 B.n48 256.663
R469 B.n405 B.n350 256.663
R470 B.n408 B.n350 256.663
R471 B.n414 B.n350 256.663
R472 B.n416 B.n350 256.663
R473 B.n422 B.n350 256.663
R474 B.n424 B.n350 256.663
R475 B.n430 B.n350 256.663
R476 B.n432 B.n350 256.663
R477 B.n438 B.n350 256.663
R478 B.n440 B.n350 256.663
R479 B.n446 B.n350 256.663
R480 B.n448 B.n350 256.663
R481 B.n454 B.n350 256.663
R482 B.n456 B.n350 256.663
R483 B.n462 B.n350 256.663
R484 B.n464 B.n350 256.663
R485 B.n470 B.n350 256.663
R486 B.n472 B.n350 256.663
R487 B.n478 B.n350 256.663
R488 B.n480 B.n350 256.663
R489 B.n486 B.n350 256.663
R490 B.n488 B.n350 256.663
R491 B.n497 B.n350 256.663
R492 B.n499 B.n350 256.663
R493 B.n505 B.n350 256.663
R494 B.n507 B.n350 256.663
R495 B.n513 B.n350 256.663
R496 B.n515 B.n350 256.663
R497 B.n522 B.n350 256.663
R498 B.n524 B.n350 256.663
R499 B.n530 B.n350 256.663
R500 B.n532 B.n350 256.663
R501 B.n538 B.n350 256.663
R502 B.n540 B.n350 256.663
R503 B.n546 B.n350 256.663
R504 B.n548 B.n350 256.663
R505 B.n554 B.n350 256.663
R506 B.n556 B.n350 256.663
R507 B.n562 B.n350 256.663
R508 B.n564 B.n350 256.663
R509 B.n570 B.n350 256.663
R510 B.n572 B.n350 256.663
R511 B.n578 B.n350 256.663
R512 B.n580 B.n350 256.663
R513 B.n586 B.n350 256.663
R514 B.n588 B.n350 256.663
R515 B.n594 B.n350 256.663
R516 B.n596 B.n350 256.663
R517 B.n602 B.n350 256.663
R518 B.n605 B.n350 256.663
R519 B.n612 B.n347 163.367
R520 B.n616 B.n347 163.367
R521 B.n616 B.n341 163.367
R522 B.n624 B.n341 163.367
R523 B.n624 B.n339 163.367
R524 B.n628 B.n339 163.367
R525 B.n628 B.n333 163.367
R526 B.n636 B.n333 163.367
R527 B.n636 B.n331 163.367
R528 B.n640 B.n331 163.367
R529 B.n640 B.n325 163.367
R530 B.n648 B.n325 163.367
R531 B.n648 B.n323 163.367
R532 B.n652 B.n323 163.367
R533 B.n652 B.n317 163.367
R534 B.n660 B.n317 163.367
R535 B.n660 B.n315 163.367
R536 B.n664 B.n315 163.367
R537 B.n664 B.n309 163.367
R538 B.n673 B.n309 163.367
R539 B.n673 B.n307 163.367
R540 B.n677 B.n307 163.367
R541 B.n677 B.n2 163.367
R542 B.n766 B.n2 163.367
R543 B.n766 B.n3 163.367
R544 B.n762 B.n3 163.367
R545 B.n762 B.n9 163.367
R546 B.n758 B.n9 163.367
R547 B.n758 B.n11 163.367
R548 B.n754 B.n11 163.367
R549 B.n754 B.n16 163.367
R550 B.n750 B.n16 163.367
R551 B.n750 B.n18 163.367
R552 B.n746 B.n18 163.367
R553 B.n746 B.n23 163.367
R554 B.n742 B.n23 163.367
R555 B.n742 B.n25 163.367
R556 B.n738 B.n25 163.367
R557 B.n738 B.n30 163.367
R558 B.n734 B.n30 163.367
R559 B.n734 B.n32 163.367
R560 B.n730 B.n32 163.367
R561 B.n730 B.n37 163.367
R562 B.n726 B.n37 163.367
R563 B.n726 B.n39 163.367
R564 B.n722 B.n39 163.367
R565 B.n722 B.n44 163.367
R566 B.n718 B.n44 163.367
R567 B.n407 B.n406 163.367
R568 B.n409 B.n407 163.367
R569 B.n413 B.n402 163.367
R570 B.n417 B.n415 163.367
R571 B.n421 B.n400 163.367
R572 B.n425 B.n423 163.367
R573 B.n429 B.n398 163.367
R574 B.n433 B.n431 163.367
R575 B.n437 B.n396 163.367
R576 B.n441 B.n439 163.367
R577 B.n445 B.n394 163.367
R578 B.n449 B.n447 163.367
R579 B.n453 B.n392 163.367
R580 B.n457 B.n455 163.367
R581 B.n461 B.n390 163.367
R582 B.n465 B.n463 163.367
R583 B.n469 B.n388 163.367
R584 B.n473 B.n471 163.367
R585 B.n477 B.n386 163.367
R586 B.n481 B.n479 163.367
R587 B.n485 B.n384 163.367
R588 B.n489 B.n487 163.367
R589 B.n496 B.n382 163.367
R590 B.n500 B.n498 163.367
R591 B.n504 B.n380 163.367
R592 B.n508 B.n506 163.367
R593 B.n512 B.n378 163.367
R594 B.n516 B.n514 163.367
R595 B.n521 B.n374 163.367
R596 B.n525 B.n523 163.367
R597 B.n529 B.n372 163.367
R598 B.n533 B.n531 163.367
R599 B.n537 B.n370 163.367
R600 B.n541 B.n539 163.367
R601 B.n545 B.n368 163.367
R602 B.n549 B.n547 163.367
R603 B.n553 B.n366 163.367
R604 B.n557 B.n555 163.367
R605 B.n561 B.n364 163.367
R606 B.n565 B.n563 163.367
R607 B.n569 B.n362 163.367
R608 B.n573 B.n571 163.367
R609 B.n577 B.n360 163.367
R610 B.n581 B.n579 163.367
R611 B.n585 B.n358 163.367
R612 B.n589 B.n587 163.367
R613 B.n593 B.n356 163.367
R614 B.n597 B.n595 163.367
R615 B.n601 B.n354 163.367
R616 B.n604 B.n603 163.367
R617 B.n606 B.n351 163.367
R618 B.n610 B.n345 163.367
R619 B.n618 B.n345 163.367
R620 B.n618 B.n343 163.367
R621 B.n622 B.n343 163.367
R622 B.n622 B.n336 163.367
R623 B.n630 B.n336 163.367
R624 B.n630 B.n334 163.367
R625 B.n634 B.n334 163.367
R626 B.n634 B.n329 163.367
R627 B.n642 B.n329 163.367
R628 B.n642 B.n327 163.367
R629 B.n646 B.n327 163.367
R630 B.n646 B.n321 163.367
R631 B.n654 B.n321 163.367
R632 B.n654 B.n319 163.367
R633 B.n658 B.n319 163.367
R634 B.n658 B.n313 163.367
R635 B.n666 B.n313 163.367
R636 B.n666 B.n311 163.367
R637 B.n671 B.n311 163.367
R638 B.n671 B.n305 163.367
R639 B.n679 B.n305 163.367
R640 B.n680 B.n679 163.367
R641 B.n680 B.n5 163.367
R642 B.n6 B.n5 163.367
R643 B.n7 B.n6 163.367
R644 B.n685 B.n7 163.367
R645 B.n685 B.n12 163.367
R646 B.n13 B.n12 163.367
R647 B.n14 B.n13 163.367
R648 B.n690 B.n14 163.367
R649 B.n690 B.n19 163.367
R650 B.n20 B.n19 163.367
R651 B.n21 B.n20 163.367
R652 B.n695 B.n21 163.367
R653 B.n695 B.n26 163.367
R654 B.n27 B.n26 163.367
R655 B.n28 B.n27 163.367
R656 B.n700 B.n28 163.367
R657 B.n700 B.n33 163.367
R658 B.n34 B.n33 163.367
R659 B.n35 B.n34 163.367
R660 B.n705 B.n35 163.367
R661 B.n705 B.n40 163.367
R662 B.n41 B.n40 163.367
R663 B.n42 B.n41 163.367
R664 B.n710 B.n42 163.367
R665 B.n710 B.n47 163.367
R666 B.n107 B.n106 163.367
R667 B.n111 B.n110 163.367
R668 B.n115 B.n114 163.367
R669 B.n119 B.n118 163.367
R670 B.n123 B.n122 163.367
R671 B.n127 B.n126 163.367
R672 B.n131 B.n130 163.367
R673 B.n135 B.n134 163.367
R674 B.n139 B.n138 163.367
R675 B.n143 B.n142 163.367
R676 B.n147 B.n146 163.367
R677 B.n151 B.n150 163.367
R678 B.n155 B.n154 163.367
R679 B.n159 B.n158 163.367
R680 B.n163 B.n162 163.367
R681 B.n167 B.n166 163.367
R682 B.n171 B.n170 163.367
R683 B.n175 B.n174 163.367
R684 B.n179 B.n178 163.367
R685 B.n183 B.n182 163.367
R686 B.n187 B.n186 163.367
R687 B.n191 B.n190 163.367
R688 B.n195 B.n194 163.367
R689 B.n199 B.n198 163.367
R690 B.n203 B.n202 163.367
R691 B.n207 B.n206 163.367
R692 B.n211 B.n210 163.367
R693 B.n215 B.n214 163.367
R694 B.n219 B.n218 163.367
R695 B.n223 B.n222 163.367
R696 B.n227 B.n226 163.367
R697 B.n231 B.n230 163.367
R698 B.n235 B.n234 163.367
R699 B.n239 B.n238 163.367
R700 B.n243 B.n242 163.367
R701 B.n247 B.n246 163.367
R702 B.n251 B.n250 163.367
R703 B.n255 B.n254 163.367
R704 B.n259 B.n258 163.367
R705 B.n263 B.n262 163.367
R706 B.n267 B.n266 163.367
R707 B.n271 B.n270 163.367
R708 B.n275 B.n274 163.367
R709 B.n279 B.n278 163.367
R710 B.n283 B.n282 163.367
R711 B.n287 B.n286 163.367
R712 B.n291 B.n290 163.367
R713 B.n295 B.n294 163.367
R714 B.n299 B.n298 163.367
R715 B.n301 B.n98 163.367
R716 B.n611 B.n350 78.9689
R717 B.n717 B.n716 78.9689
R718 B.n405 B.n349 71.676
R719 B.n409 B.n408 71.676
R720 B.n414 B.n413 71.676
R721 B.n417 B.n416 71.676
R722 B.n422 B.n421 71.676
R723 B.n425 B.n424 71.676
R724 B.n430 B.n429 71.676
R725 B.n433 B.n432 71.676
R726 B.n438 B.n437 71.676
R727 B.n441 B.n440 71.676
R728 B.n446 B.n445 71.676
R729 B.n449 B.n448 71.676
R730 B.n454 B.n453 71.676
R731 B.n457 B.n456 71.676
R732 B.n462 B.n461 71.676
R733 B.n465 B.n464 71.676
R734 B.n470 B.n469 71.676
R735 B.n473 B.n472 71.676
R736 B.n478 B.n477 71.676
R737 B.n481 B.n480 71.676
R738 B.n486 B.n485 71.676
R739 B.n489 B.n488 71.676
R740 B.n497 B.n496 71.676
R741 B.n500 B.n499 71.676
R742 B.n505 B.n504 71.676
R743 B.n508 B.n507 71.676
R744 B.n513 B.n512 71.676
R745 B.n516 B.n515 71.676
R746 B.n522 B.n521 71.676
R747 B.n525 B.n524 71.676
R748 B.n530 B.n529 71.676
R749 B.n533 B.n532 71.676
R750 B.n538 B.n537 71.676
R751 B.n541 B.n540 71.676
R752 B.n546 B.n545 71.676
R753 B.n549 B.n548 71.676
R754 B.n554 B.n553 71.676
R755 B.n557 B.n556 71.676
R756 B.n562 B.n561 71.676
R757 B.n565 B.n564 71.676
R758 B.n570 B.n569 71.676
R759 B.n573 B.n572 71.676
R760 B.n578 B.n577 71.676
R761 B.n581 B.n580 71.676
R762 B.n586 B.n585 71.676
R763 B.n589 B.n588 71.676
R764 B.n594 B.n593 71.676
R765 B.n597 B.n596 71.676
R766 B.n602 B.n601 71.676
R767 B.n605 B.n604 71.676
R768 B.n48 B.n46 71.676
R769 B.n107 B.n49 71.676
R770 B.n111 B.n50 71.676
R771 B.n115 B.n51 71.676
R772 B.n119 B.n52 71.676
R773 B.n123 B.n53 71.676
R774 B.n127 B.n54 71.676
R775 B.n131 B.n55 71.676
R776 B.n135 B.n56 71.676
R777 B.n139 B.n57 71.676
R778 B.n143 B.n58 71.676
R779 B.n147 B.n59 71.676
R780 B.n151 B.n60 71.676
R781 B.n155 B.n61 71.676
R782 B.n159 B.n62 71.676
R783 B.n163 B.n63 71.676
R784 B.n167 B.n64 71.676
R785 B.n171 B.n65 71.676
R786 B.n175 B.n66 71.676
R787 B.n179 B.n67 71.676
R788 B.n183 B.n68 71.676
R789 B.n187 B.n69 71.676
R790 B.n191 B.n70 71.676
R791 B.n195 B.n71 71.676
R792 B.n199 B.n72 71.676
R793 B.n203 B.n73 71.676
R794 B.n207 B.n74 71.676
R795 B.n211 B.n75 71.676
R796 B.n215 B.n76 71.676
R797 B.n219 B.n77 71.676
R798 B.n223 B.n78 71.676
R799 B.n227 B.n79 71.676
R800 B.n231 B.n80 71.676
R801 B.n235 B.n81 71.676
R802 B.n239 B.n82 71.676
R803 B.n243 B.n83 71.676
R804 B.n247 B.n84 71.676
R805 B.n251 B.n85 71.676
R806 B.n255 B.n86 71.676
R807 B.n259 B.n87 71.676
R808 B.n263 B.n88 71.676
R809 B.n267 B.n89 71.676
R810 B.n271 B.n90 71.676
R811 B.n275 B.n91 71.676
R812 B.n279 B.n92 71.676
R813 B.n283 B.n93 71.676
R814 B.n287 B.n94 71.676
R815 B.n291 B.n95 71.676
R816 B.n295 B.n96 71.676
R817 B.n299 B.n97 71.676
R818 B.n715 B.n98 71.676
R819 B.n715 B.n714 71.676
R820 B.n301 B.n97 71.676
R821 B.n298 B.n96 71.676
R822 B.n294 B.n95 71.676
R823 B.n290 B.n94 71.676
R824 B.n286 B.n93 71.676
R825 B.n282 B.n92 71.676
R826 B.n278 B.n91 71.676
R827 B.n274 B.n90 71.676
R828 B.n270 B.n89 71.676
R829 B.n266 B.n88 71.676
R830 B.n262 B.n87 71.676
R831 B.n258 B.n86 71.676
R832 B.n254 B.n85 71.676
R833 B.n250 B.n84 71.676
R834 B.n246 B.n83 71.676
R835 B.n242 B.n82 71.676
R836 B.n238 B.n81 71.676
R837 B.n234 B.n80 71.676
R838 B.n230 B.n79 71.676
R839 B.n226 B.n78 71.676
R840 B.n222 B.n77 71.676
R841 B.n218 B.n76 71.676
R842 B.n214 B.n75 71.676
R843 B.n210 B.n74 71.676
R844 B.n206 B.n73 71.676
R845 B.n202 B.n72 71.676
R846 B.n198 B.n71 71.676
R847 B.n194 B.n70 71.676
R848 B.n190 B.n69 71.676
R849 B.n186 B.n68 71.676
R850 B.n182 B.n67 71.676
R851 B.n178 B.n66 71.676
R852 B.n174 B.n65 71.676
R853 B.n170 B.n64 71.676
R854 B.n166 B.n63 71.676
R855 B.n162 B.n62 71.676
R856 B.n158 B.n61 71.676
R857 B.n154 B.n60 71.676
R858 B.n150 B.n59 71.676
R859 B.n146 B.n58 71.676
R860 B.n142 B.n57 71.676
R861 B.n138 B.n56 71.676
R862 B.n134 B.n55 71.676
R863 B.n130 B.n54 71.676
R864 B.n126 B.n53 71.676
R865 B.n122 B.n52 71.676
R866 B.n118 B.n51 71.676
R867 B.n114 B.n50 71.676
R868 B.n110 B.n49 71.676
R869 B.n106 B.n48 71.676
R870 B.n406 B.n405 71.676
R871 B.n408 B.n402 71.676
R872 B.n415 B.n414 71.676
R873 B.n416 B.n400 71.676
R874 B.n423 B.n422 71.676
R875 B.n424 B.n398 71.676
R876 B.n431 B.n430 71.676
R877 B.n432 B.n396 71.676
R878 B.n439 B.n438 71.676
R879 B.n440 B.n394 71.676
R880 B.n447 B.n446 71.676
R881 B.n448 B.n392 71.676
R882 B.n455 B.n454 71.676
R883 B.n456 B.n390 71.676
R884 B.n463 B.n462 71.676
R885 B.n464 B.n388 71.676
R886 B.n471 B.n470 71.676
R887 B.n472 B.n386 71.676
R888 B.n479 B.n478 71.676
R889 B.n480 B.n384 71.676
R890 B.n487 B.n486 71.676
R891 B.n488 B.n382 71.676
R892 B.n498 B.n497 71.676
R893 B.n499 B.n380 71.676
R894 B.n506 B.n505 71.676
R895 B.n507 B.n378 71.676
R896 B.n514 B.n513 71.676
R897 B.n515 B.n374 71.676
R898 B.n523 B.n522 71.676
R899 B.n524 B.n372 71.676
R900 B.n531 B.n530 71.676
R901 B.n532 B.n370 71.676
R902 B.n539 B.n538 71.676
R903 B.n540 B.n368 71.676
R904 B.n547 B.n546 71.676
R905 B.n548 B.n366 71.676
R906 B.n555 B.n554 71.676
R907 B.n556 B.n364 71.676
R908 B.n563 B.n562 71.676
R909 B.n564 B.n362 71.676
R910 B.n571 B.n570 71.676
R911 B.n572 B.n360 71.676
R912 B.n579 B.n578 71.676
R913 B.n580 B.n358 71.676
R914 B.n587 B.n586 71.676
R915 B.n588 B.n356 71.676
R916 B.n595 B.n594 71.676
R917 B.n596 B.n354 71.676
R918 B.n603 B.n602 71.676
R919 B.n606 B.n605 71.676
R920 B.n518 B.n376 59.5399
R921 B.n494 B.n493 59.5399
R922 B.n104 B.n103 59.5399
R923 B.n101 B.n100 59.5399
R924 B.n376 B.n375 52.946
R925 B.n493 B.n492 52.946
R926 B.n103 B.n102 52.946
R927 B.n100 B.n99 52.946
R928 B.n611 B.n346 39.7772
R929 B.n617 B.n346 39.7772
R930 B.n617 B.n342 39.7772
R931 B.n623 B.n342 39.7772
R932 B.n623 B.n337 39.7772
R933 B.n629 B.n337 39.7772
R934 B.n629 B.n338 39.7772
R935 B.n635 B.n330 39.7772
R936 B.n641 B.n330 39.7772
R937 B.n641 B.n326 39.7772
R938 B.n647 B.n326 39.7772
R939 B.n647 B.n322 39.7772
R940 B.n653 B.n322 39.7772
R941 B.n653 B.n318 39.7772
R942 B.n659 B.n318 39.7772
R943 B.n659 B.n314 39.7772
R944 B.n665 B.n314 39.7772
R945 B.n672 B.n310 39.7772
R946 B.n672 B.n306 39.7772
R947 B.n678 B.n306 39.7772
R948 B.n678 B.n4 39.7772
R949 B.n765 B.n4 39.7772
R950 B.n765 B.n764 39.7772
R951 B.n764 B.n763 39.7772
R952 B.n763 B.n8 39.7772
R953 B.n757 B.n8 39.7772
R954 B.n757 B.n756 39.7772
R955 B.n755 B.n15 39.7772
R956 B.n749 B.n15 39.7772
R957 B.n749 B.n748 39.7772
R958 B.n748 B.n747 39.7772
R959 B.n747 B.n22 39.7772
R960 B.n741 B.n22 39.7772
R961 B.n741 B.n740 39.7772
R962 B.n740 B.n739 39.7772
R963 B.n739 B.n29 39.7772
R964 B.n733 B.n29 39.7772
R965 B.n732 B.n731 39.7772
R966 B.n731 B.n36 39.7772
R967 B.n725 B.n36 39.7772
R968 B.n725 B.n724 39.7772
R969 B.n724 B.n723 39.7772
R970 B.n723 B.n43 39.7772
R971 B.n717 B.n43 39.7772
R972 B.n635 B.t3 33.9276
R973 B.n733 B.t7 33.9276
R974 B.n719 B.n45 33.2493
R975 B.n713 B.n712 33.2493
R976 B.n609 B.n608 33.2493
R977 B.n613 B.n348 33.2493
R978 B.t0 B.n310 24.5684
R979 B.n756 B.t1 24.5684
R980 B B.n767 18.0485
R981 B.n665 B.t0 15.2092
R982 B.t1 B.n755 15.2092
R983 B.n105 B.n45 10.6151
R984 B.n108 B.n105 10.6151
R985 B.n109 B.n108 10.6151
R986 B.n112 B.n109 10.6151
R987 B.n113 B.n112 10.6151
R988 B.n116 B.n113 10.6151
R989 B.n117 B.n116 10.6151
R990 B.n120 B.n117 10.6151
R991 B.n121 B.n120 10.6151
R992 B.n124 B.n121 10.6151
R993 B.n125 B.n124 10.6151
R994 B.n128 B.n125 10.6151
R995 B.n129 B.n128 10.6151
R996 B.n132 B.n129 10.6151
R997 B.n133 B.n132 10.6151
R998 B.n136 B.n133 10.6151
R999 B.n137 B.n136 10.6151
R1000 B.n140 B.n137 10.6151
R1001 B.n141 B.n140 10.6151
R1002 B.n144 B.n141 10.6151
R1003 B.n145 B.n144 10.6151
R1004 B.n148 B.n145 10.6151
R1005 B.n149 B.n148 10.6151
R1006 B.n152 B.n149 10.6151
R1007 B.n153 B.n152 10.6151
R1008 B.n156 B.n153 10.6151
R1009 B.n157 B.n156 10.6151
R1010 B.n160 B.n157 10.6151
R1011 B.n161 B.n160 10.6151
R1012 B.n164 B.n161 10.6151
R1013 B.n165 B.n164 10.6151
R1014 B.n168 B.n165 10.6151
R1015 B.n169 B.n168 10.6151
R1016 B.n172 B.n169 10.6151
R1017 B.n173 B.n172 10.6151
R1018 B.n176 B.n173 10.6151
R1019 B.n177 B.n176 10.6151
R1020 B.n180 B.n177 10.6151
R1021 B.n181 B.n180 10.6151
R1022 B.n184 B.n181 10.6151
R1023 B.n185 B.n184 10.6151
R1024 B.n188 B.n185 10.6151
R1025 B.n189 B.n188 10.6151
R1026 B.n192 B.n189 10.6151
R1027 B.n193 B.n192 10.6151
R1028 B.n197 B.n196 10.6151
R1029 B.n200 B.n197 10.6151
R1030 B.n201 B.n200 10.6151
R1031 B.n204 B.n201 10.6151
R1032 B.n205 B.n204 10.6151
R1033 B.n208 B.n205 10.6151
R1034 B.n209 B.n208 10.6151
R1035 B.n212 B.n209 10.6151
R1036 B.n213 B.n212 10.6151
R1037 B.n217 B.n216 10.6151
R1038 B.n220 B.n217 10.6151
R1039 B.n221 B.n220 10.6151
R1040 B.n224 B.n221 10.6151
R1041 B.n225 B.n224 10.6151
R1042 B.n228 B.n225 10.6151
R1043 B.n229 B.n228 10.6151
R1044 B.n232 B.n229 10.6151
R1045 B.n233 B.n232 10.6151
R1046 B.n236 B.n233 10.6151
R1047 B.n237 B.n236 10.6151
R1048 B.n240 B.n237 10.6151
R1049 B.n241 B.n240 10.6151
R1050 B.n244 B.n241 10.6151
R1051 B.n245 B.n244 10.6151
R1052 B.n248 B.n245 10.6151
R1053 B.n249 B.n248 10.6151
R1054 B.n252 B.n249 10.6151
R1055 B.n253 B.n252 10.6151
R1056 B.n256 B.n253 10.6151
R1057 B.n257 B.n256 10.6151
R1058 B.n260 B.n257 10.6151
R1059 B.n261 B.n260 10.6151
R1060 B.n264 B.n261 10.6151
R1061 B.n265 B.n264 10.6151
R1062 B.n268 B.n265 10.6151
R1063 B.n269 B.n268 10.6151
R1064 B.n272 B.n269 10.6151
R1065 B.n273 B.n272 10.6151
R1066 B.n276 B.n273 10.6151
R1067 B.n277 B.n276 10.6151
R1068 B.n280 B.n277 10.6151
R1069 B.n281 B.n280 10.6151
R1070 B.n284 B.n281 10.6151
R1071 B.n285 B.n284 10.6151
R1072 B.n288 B.n285 10.6151
R1073 B.n289 B.n288 10.6151
R1074 B.n292 B.n289 10.6151
R1075 B.n293 B.n292 10.6151
R1076 B.n296 B.n293 10.6151
R1077 B.n297 B.n296 10.6151
R1078 B.n300 B.n297 10.6151
R1079 B.n302 B.n300 10.6151
R1080 B.n303 B.n302 10.6151
R1081 B.n713 B.n303 10.6151
R1082 B.n609 B.n344 10.6151
R1083 B.n619 B.n344 10.6151
R1084 B.n620 B.n619 10.6151
R1085 B.n621 B.n620 10.6151
R1086 B.n621 B.n335 10.6151
R1087 B.n631 B.n335 10.6151
R1088 B.n632 B.n631 10.6151
R1089 B.n633 B.n632 10.6151
R1090 B.n633 B.n328 10.6151
R1091 B.n643 B.n328 10.6151
R1092 B.n644 B.n643 10.6151
R1093 B.n645 B.n644 10.6151
R1094 B.n645 B.n320 10.6151
R1095 B.n655 B.n320 10.6151
R1096 B.n656 B.n655 10.6151
R1097 B.n657 B.n656 10.6151
R1098 B.n657 B.n312 10.6151
R1099 B.n667 B.n312 10.6151
R1100 B.n668 B.n667 10.6151
R1101 B.n670 B.n668 10.6151
R1102 B.n670 B.n669 10.6151
R1103 B.n669 B.n304 10.6151
R1104 B.n681 B.n304 10.6151
R1105 B.n682 B.n681 10.6151
R1106 B.n683 B.n682 10.6151
R1107 B.n684 B.n683 10.6151
R1108 B.n686 B.n684 10.6151
R1109 B.n687 B.n686 10.6151
R1110 B.n688 B.n687 10.6151
R1111 B.n689 B.n688 10.6151
R1112 B.n691 B.n689 10.6151
R1113 B.n692 B.n691 10.6151
R1114 B.n693 B.n692 10.6151
R1115 B.n694 B.n693 10.6151
R1116 B.n696 B.n694 10.6151
R1117 B.n697 B.n696 10.6151
R1118 B.n698 B.n697 10.6151
R1119 B.n699 B.n698 10.6151
R1120 B.n701 B.n699 10.6151
R1121 B.n702 B.n701 10.6151
R1122 B.n703 B.n702 10.6151
R1123 B.n704 B.n703 10.6151
R1124 B.n706 B.n704 10.6151
R1125 B.n707 B.n706 10.6151
R1126 B.n708 B.n707 10.6151
R1127 B.n709 B.n708 10.6151
R1128 B.n711 B.n709 10.6151
R1129 B.n712 B.n711 10.6151
R1130 B.n404 B.n348 10.6151
R1131 B.n404 B.n403 10.6151
R1132 B.n410 B.n403 10.6151
R1133 B.n411 B.n410 10.6151
R1134 B.n412 B.n411 10.6151
R1135 B.n412 B.n401 10.6151
R1136 B.n418 B.n401 10.6151
R1137 B.n419 B.n418 10.6151
R1138 B.n420 B.n419 10.6151
R1139 B.n420 B.n399 10.6151
R1140 B.n426 B.n399 10.6151
R1141 B.n427 B.n426 10.6151
R1142 B.n428 B.n427 10.6151
R1143 B.n428 B.n397 10.6151
R1144 B.n434 B.n397 10.6151
R1145 B.n435 B.n434 10.6151
R1146 B.n436 B.n435 10.6151
R1147 B.n436 B.n395 10.6151
R1148 B.n442 B.n395 10.6151
R1149 B.n443 B.n442 10.6151
R1150 B.n444 B.n443 10.6151
R1151 B.n444 B.n393 10.6151
R1152 B.n450 B.n393 10.6151
R1153 B.n451 B.n450 10.6151
R1154 B.n452 B.n451 10.6151
R1155 B.n452 B.n391 10.6151
R1156 B.n458 B.n391 10.6151
R1157 B.n459 B.n458 10.6151
R1158 B.n460 B.n459 10.6151
R1159 B.n460 B.n389 10.6151
R1160 B.n466 B.n389 10.6151
R1161 B.n467 B.n466 10.6151
R1162 B.n468 B.n467 10.6151
R1163 B.n468 B.n387 10.6151
R1164 B.n474 B.n387 10.6151
R1165 B.n475 B.n474 10.6151
R1166 B.n476 B.n475 10.6151
R1167 B.n476 B.n385 10.6151
R1168 B.n482 B.n385 10.6151
R1169 B.n483 B.n482 10.6151
R1170 B.n484 B.n483 10.6151
R1171 B.n484 B.n383 10.6151
R1172 B.n490 B.n383 10.6151
R1173 B.n491 B.n490 10.6151
R1174 B.n495 B.n491 10.6151
R1175 B.n501 B.n381 10.6151
R1176 B.n502 B.n501 10.6151
R1177 B.n503 B.n502 10.6151
R1178 B.n503 B.n379 10.6151
R1179 B.n509 B.n379 10.6151
R1180 B.n510 B.n509 10.6151
R1181 B.n511 B.n510 10.6151
R1182 B.n511 B.n377 10.6151
R1183 B.n517 B.n377 10.6151
R1184 B.n520 B.n519 10.6151
R1185 B.n520 B.n373 10.6151
R1186 B.n526 B.n373 10.6151
R1187 B.n527 B.n526 10.6151
R1188 B.n528 B.n527 10.6151
R1189 B.n528 B.n371 10.6151
R1190 B.n534 B.n371 10.6151
R1191 B.n535 B.n534 10.6151
R1192 B.n536 B.n535 10.6151
R1193 B.n536 B.n369 10.6151
R1194 B.n542 B.n369 10.6151
R1195 B.n543 B.n542 10.6151
R1196 B.n544 B.n543 10.6151
R1197 B.n544 B.n367 10.6151
R1198 B.n550 B.n367 10.6151
R1199 B.n551 B.n550 10.6151
R1200 B.n552 B.n551 10.6151
R1201 B.n552 B.n365 10.6151
R1202 B.n558 B.n365 10.6151
R1203 B.n559 B.n558 10.6151
R1204 B.n560 B.n559 10.6151
R1205 B.n560 B.n363 10.6151
R1206 B.n566 B.n363 10.6151
R1207 B.n567 B.n566 10.6151
R1208 B.n568 B.n567 10.6151
R1209 B.n568 B.n361 10.6151
R1210 B.n574 B.n361 10.6151
R1211 B.n575 B.n574 10.6151
R1212 B.n576 B.n575 10.6151
R1213 B.n576 B.n359 10.6151
R1214 B.n582 B.n359 10.6151
R1215 B.n583 B.n582 10.6151
R1216 B.n584 B.n583 10.6151
R1217 B.n584 B.n357 10.6151
R1218 B.n590 B.n357 10.6151
R1219 B.n591 B.n590 10.6151
R1220 B.n592 B.n591 10.6151
R1221 B.n592 B.n355 10.6151
R1222 B.n598 B.n355 10.6151
R1223 B.n599 B.n598 10.6151
R1224 B.n600 B.n599 10.6151
R1225 B.n600 B.n353 10.6151
R1226 B.n353 B.n352 10.6151
R1227 B.n607 B.n352 10.6151
R1228 B.n608 B.n607 10.6151
R1229 B.n614 B.n613 10.6151
R1230 B.n615 B.n614 10.6151
R1231 B.n615 B.n340 10.6151
R1232 B.n625 B.n340 10.6151
R1233 B.n626 B.n625 10.6151
R1234 B.n627 B.n626 10.6151
R1235 B.n627 B.n332 10.6151
R1236 B.n637 B.n332 10.6151
R1237 B.n638 B.n637 10.6151
R1238 B.n639 B.n638 10.6151
R1239 B.n639 B.n324 10.6151
R1240 B.n649 B.n324 10.6151
R1241 B.n650 B.n649 10.6151
R1242 B.n651 B.n650 10.6151
R1243 B.n651 B.n316 10.6151
R1244 B.n661 B.n316 10.6151
R1245 B.n662 B.n661 10.6151
R1246 B.n663 B.n662 10.6151
R1247 B.n663 B.n308 10.6151
R1248 B.n674 B.n308 10.6151
R1249 B.n675 B.n674 10.6151
R1250 B.n676 B.n675 10.6151
R1251 B.n676 B.n0 10.6151
R1252 B.n761 B.n1 10.6151
R1253 B.n761 B.n760 10.6151
R1254 B.n760 B.n759 10.6151
R1255 B.n759 B.n10 10.6151
R1256 B.n753 B.n10 10.6151
R1257 B.n753 B.n752 10.6151
R1258 B.n752 B.n751 10.6151
R1259 B.n751 B.n17 10.6151
R1260 B.n745 B.n17 10.6151
R1261 B.n745 B.n744 10.6151
R1262 B.n744 B.n743 10.6151
R1263 B.n743 B.n24 10.6151
R1264 B.n737 B.n24 10.6151
R1265 B.n737 B.n736 10.6151
R1266 B.n736 B.n735 10.6151
R1267 B.n735 B.n31 10.6151
R1268 B.n729 B.n31 10.6151
R1269 B.n729 B.n728 10.6151
R1270 B.n728 B.n727 10.6151
R1271 B.n727 B.n38 10.6151
R1272 B.n721 B.n38 10.6151
R1273 B.n721 B.n720 10.6151
R1274 B.n720 B.n719 10.6151
R1275 B.n193 B.n104 9.36635
R1276 B.n216 B.n101 9.36635
R1277 B.n495 B.n494 9.36635
R1278 B.n519 B.n518 9.36635
R1279 B.n338 B.t3 5.85001
R1280 B.t7 B.n732 5.85001
R1281 B.n767 B.n0 2.81026
R1282 B.n767 B.n1 2.81026
R1283 B.n196 B.n104 1.24928
R1284 B.n213 B.n101 1.24928
R1285 B.n494 B.n381 1.24928
R1286 B.n518 B.n517 1.24928
R1287 VP.n0 VP.t1 230.32
R1288 VP.n0 VP.t0 185.035
R1289 VP VP.n0 0.336784
R1290 VTAIL.n290 VTAIL.n222 289.615
R1291 VTAIL.n68 VTAIL.n0 289.615
R1292 VTAIL.n216 VTAIL.n148 289.615
R1293 VTAIL.n142 VTAIL.n74 289.615
R1294 VTAIL.n247 VTAIL.n246 185
R1295 VTAIL.n249 VTAIL.n248 185
R1296 VTAIL.n242 VTAIL.n241 185
R1297 VTAIL.n255 VTAIL.n254 185
R1298 VTAIL.n257 VTAIL.n256 185
R1299 VTAIL.n238 VTAIL.n237 185
R1300 VTAIL.n264 VTAIL.n263 185
R1301 VTAIL.n265 VTAIL.n236 185
R1302 VTAIL.n267 VTAIL.n266 185
R1303 VTAIL.n234 VTAIL.n233 185
R1304 VTAIL.n273 VTAIL.n272 185
R1305 VTAIL.n275 VTAIL.n274 185
R1306 VTAIL.n230 VTAIL.n229 185
R1307 VTAIL.n281 VTAIL.n280 185
R1308 VTAIL.n283 VTAIL.n282 185
R1309 VTAIL.n226 VTAIL.n225 185
R1310 VTAIL.n289 VTAIL.n288 185
R1311 VTAIL.n291 VTAIL.n290 185
R1312 VTAIL.n25 VTAIL.n24 185
R1313 VTAIL.n27 VTAIL.n26 185
R1314 VTAIL.n20 VTAIL.n19 185
R1315 VTAIL.n33 VTAIL.n32 185
R1316 VTAIL.n35 VTAIL.n34 185
R1317 VTAIL.n16 VTAIL.n15 185
R1318 VTAIL.n42 VTAIL.n41 185
R1319 VTAIL.n43 VTAIL.n14 185
R1320 VTAIL.n45 VTAIL.n44 185
R1321 VTAIL.n12 VTAIL.n11 185
R1322 VTAIL.n51 VTAIL.n50 185
R1323 VTAIL.n53 VTAIL.n52 185
R1324 VTAIL.n8 VTAIL.n7 185
R1325 VTAIL.n59 VTAIL.n58 185
R1326 VTAIL.n61 VTAIL.n60 185
R1327 VTAIL.n4 VTAIL.n3 185
R1328 VTAIL.n67 VTAIL.n66 185
R1329 VTAIL.n69 VTAIL.n68 185
R1330 VTAIL.n217 VTAIL.n216 185
R1331 VTAIL.n215 VTAIL.n214 185
R1332 VTAIL.n152 VTAIL.n151 185
R1333 VTAIL.n209 VTAIL.n208 185
R1334 VTAIL.n207 VTAIL.n206 185
R1335 VTAIL.n156 VTAIL.n155 185
R1336 VTAIL.n201 VTAIL.n200 185
R1337 VTAIL.n199 VTAIL.n198 185
R1338 VTAIL.n160 VTAIL.n159 185
R1339 VTAIL.n164 VTAIL.n162 185
R1340 VTAIL.n193 VTAIL.n192 185
R1341 VTAIL.n191 VTAIL.n190 185
R1342 VTAIL.n166 VTAIL.n165 185
R1343 VTAIL.n185 VTAIL.n184 185
R1344 VTAIL.n183 VTAIL.n182 185
R1345 VTAIL.n170 VTAIL.n169 185
R1346 VTAIL.n177 VTAIL.n176 185
R1347 VTAIL.n175 VTAIL.n174 185
R1348 VTAIL.n143 VTAIL.n142 185
R1349 VTAIL.n141 VTAIL.n140 185
R1350 VTAIL.n78 VTAIL.n77 185
R1351 VTAIL.n135 VTAIL.n134 185
R1352 VTAIL.n133 VTAIL.n132 185
R1353 VTAIL.n82 VTAIL.n81 185
R1354 VTAIL.n127 VTAIL.n126 185
R1355 VTAIL.n125 VTAIL.n124 185
R1356 VTAIL.n86 VTAIL.n85 185
R1357 VTAIL.n90 VTAIL.n88 185
R1358 VTAIL.n119 VTAIL.n118 185
R1359 VTAIL.n117 VTAIL.n116 185
R1360 VTAIL.n92 VTAIL.n91 185
R1361 VTAIL.n111 VTAIL.n110 185
R1362 VTAIL.n109 VTAIL.n108 185
R1363 VTAIL.n96 VTAIL.n95 185
R1364 VTAIL.n103 VTAIL.n102 185
R1365 VTAIL.n101 VTAIL.n100 185
R1366 VTAIL.n245 VTAIL.t1 149.524
R1367 VTAIL.n23 VTAIL.t2 149.524
R1368 VTAIL.n173 VTAIL.t3 149.524
R1369 VTAIL.n99 VTAIL.t0 149.524
R1370 VTAIL.n248 VTAIL.n247 104.615
R1371 VTAIL.n248 VTAIL.n241 104.615
R1372 VTAIL.n255 VTAIL.n241 104.615
R1373 VTAIL.n256 VTAIL.n255 104.615
R1374 VTAIL.n256 VTAIL.n237 104.615
R1375 VTAIL.n264 VTAIL.n237 104.615
R1376 VTAIL.n265 VTAIL.n264 104.615
R1377 VTAIL.n266 VTAIL.n265 104.615
R1378 VTAIL.n266 VTAIL.n233 104.615
R1379 VTAIL.n273 VTAIL.n233 104.615
R1380 VTAIL.n274 VTAIL.n273 104.615
R1381 VTAIL.n274 VTAIL.n229 104.615
R1382 VTAIL.n281 VTAIL.n229 104.615
R1383 VTAIL.n282 VTAIL.n281 104.615
R1384 VTAIL.n282 VTAIL.n225 104.615
R1385 VTAIL.n289 VTAIL.n225 104.615
R1386 VTAIL.n290 VTAIL.n289 104.615
R1387 VTAIL.n26 VTAIL.n25 104.615
R1388 VTAIL.n26 VTAIL.n19 104.615
R1389 VTAIL.n33 VTAIL.n19 104.615
R1390 VTAIL.n34 VTAIL.n33 104.615
R1391 VTAIL.n34 VTAIL.n15 104.615
R1392 VTAIL.n42 VTAIL.n15 104.615
R1393 VTAIL.n43 VTAIL.n42 104.615
R1394 VTAIL.n44 VTAIL.n43 104.615
R1395 VTAIL.n44 VTAIL.n11 104.615
R1396 VTAIL.n51 VTAIL.n11 104.615
R1397 VTAIL.n52 VTAIL.n51 104.615
R1398 VTAIL.n52 VTAIL.n7 104.615
R1399 VTAIL.n59 VTAIL.n7 104.615
R1400 VTAIL.n60 VTAIL.n59 104.615
R1401 VTAIL.n60 VTAIL.n3 104.615
R1402 VTAIL.n67 VTAIL.n3 104.615
R1403 VTAIL.n68 VTAIL.n67 104.615
R1404 VTAIL.n216 VTAIL.n215 104.615
R1405 VTAIL.n215 VTAIL.n151 104.615
R1406 VTAIL.n208 VTAIL.n151 104.615
R1407 VTAIL.n208 VTAIL.n207 104.615
R1408 VTAIL.n207 VTAIL.n155 104.615
R1409 VTAIL.n200 VTAIL.n155 104.615
R1410 VTAIL.n200 VTAIL.n199 104.615
R1411 VTAIL.n199 VTAIL.n159 104.615
R1412 VTAIL.n164 VTAIL.n159 104.615
R1413 VTAIL.n192 VTAIL.n164 104.615
R1414 VTAIL.n192 VTAIL.n191 104.615
R1415 VTAIL.n191 VTAIL.n165 104.615
R1416 VTAIL.n184 VTAIL.n165 104.615
R1417 VTAIL.n184 VTAIL.n183 104.615
R1418 VTAIL.n183 VTAIL.n169 104.615
R1419 VTAIL.n176 VTAIL.n169 104.615
R1420 VTAIL.n176 VTAIL.n175 104.615
R1421 VTAIL.n142 VTAIL.n141 104.615
R1422 VTAIL.n141 VTAIL.n77 104.615
R1423 VTAIL.n134 VTAIL.n77 104.615
R1424 VTAIL.n134 VTAIL.n133 104.615
R1425 VTAIL.n133 VTAIL.n81 104.615
R1426 VTAIL.n126 VTAIL.n81 104.615
R1427 VTAIL.n126 VTAIL.n125 104.615
R1428 VTAIL.n125 VTAIL.n85 104.615
R1429 VTAIL.n90 VTAIL.n85 104.615
R1430 VTAIL.n118 VTAIL.n90 104.615
R1431 VTAIL.n118 VTAIL.n117 104.615
R1432 VTAIL.n117 VTAIL.n91 104.615
R1433 VTAIL.n110 VTAIL.n91 104.615
R1434 VTAIL.n110 VTAIL.n109 104.615
R1435 VTAIL.n109 VTAIL.n95 104.615
R1436 VTAIL.n102 VTAIL.n95 104.615
R1437 VTAIL.n102 VTAIL.n101 104.615
R1438 VTAIL.n247 VTAIL.t1 52.3082
R1439 VTAIL.n25 VTAIL.t2 52.3082
R1440 VTAIL.n175 VTAIL.t3 52.3082
R1441 VTAIL.n101 VTAIL.t0 52.3082
R1442 VTAIL.n295 VTAIL.n294 31.6035
R1443 VTAIL.n73 VTAIL.n72 31.6035
R1444 VTAIL.n221 VTAIL.n220 31.6035
R1445 VTAIL.n147 VTAIL.n146 31.6035
R1446 VTAIL.n147 VTAIL.n73 28.7376
R1447 VTAIL.n295 VTAIL.n221 26.3841
R1448 VTAIL.n267 VTAIL.n234 13.1884
R1449 VTAIL.n45 VTAIL.n12 13.1884
R1450 VTAIL.n162 VTAIL.n160 13.1884
R1451 VTAIL.n88 VTAIL.n86 13.1884
R1452 VTAIL.n268 VTAIL.n236 12.8005
R1453 VTAIL.n272 VTAIL.n271 12.8005
R1454 VTAIL.n46 VTAIL.n14 12.8005
R1455 VTAIL.n50 VTAIL.n49 12.8005
R1456 VTAIL.n198 VTAIL.n197 12.8005
R1457 VTAIL.n194 VTAIL.n193 12.8005
R1458 VTAIL.n124 VTAIL.n123 12.8005
R1459 VTAIL.n120 VTAIL.n119 12.8005
R1460 VTAIL.n263 VTAIL.n262 12.0247
R1461 VTAIL.n275 VTAIL.n232 12.0247
R1462 VTAIL.n41 VTAIL.n40 12.0247
R1463 VTAIL.n53 VTAIL.n10 12.0247
R1464 VTAIL.n201 VTAIL.n158 12.0247
R1465 VTAIL.n190 VTAIL.n163 12.0247
R1466 VTAIL.n127 VTAIL.n84 12.0247
R1467 VTAIL.n116 VTAIL.n89 12.0247
R1468 VTAIL.n261 VTAIL.n238 11.249
R1469 VTAIL.n276 VTAIL.n230 11.249
R1470 VTAIL.n39 VTAIL.n16 11.249
R1471 VTAIL.n54 VTAIL.n8 11.249
R1472 VTAIL.n202 VTAIL.n156 11.249
R1473 VTAIL.n189 VTAIL.n166 11.249
R1474 VTAIL.n128 VTAIL.n82 11.249
R1475 VTAIL.n115 VTAIL.n92 11.249
R1476 VTAIL.n258 VTAIL.n257 10.4732
R1477 VTAIL.n280 VTAIL.n279 10.4732
R1478 VTAIL.n36 VTAIL.n35 10.4732
R1479 VTAIL.n58 VTAIL.n57 10.4732
R1480 VTAIL.n206 VTAIL.n205 10.4732
R1481 VTAIL.n186 VTAIL.n185 10.4732
R1482 VTAIL.n132 VTAIL.n131 10.4732
R1483 VTAIL.n112 VTAIL.n111 10.4732
R1484 VTAIL.n246 VTAIL.n245 10.2747
R1485 VTAIL.n24 VTAIL.n23 10.2747
R1486 VTAIL.n174 VTAIL.n173 10.2747
R1487 VTAIL.n100 VTAIL.n99 10.2747
R1488 VTAIL.n254 VTAIL.n240 9.69747
R1489 VTAIL.n283 VTAIL.n228 9.69747
R1490 VTAIL.n32 VTAIL.n18 9.69747
R1491 VTAIL.n61 VTAIL.n6 9.69747
R1492 VTAIL.n209 VTAIL.n154 9.69747
R1493 VTAIL.n182 VTAIL.n168 9.69747
R1494 VTAIL.n135 VTAIL.n80 9.69747
R1495 VTAIL.n108 VTAIL.n94 9.69747
R1496 VTAIL.n294 VTAIL.n293 9.45567
R1497 VTAIL.n72 VTAIL.n71 9.45567
R1498 VTAIL.n220 VTAIL.n219 9.45567
R1499 VTAIL.n146 VTAIL.n145 9.45567
R1500 VTAIL.n293 VTAIL.n292 9.3005
R1501 VTAIL.n287 VTAIL.n286 9.3005
R1502 VTAIL.n285 VTAIL.n284 9.3005
R1503 VTAIL.n228 VTAIL.n227 9.3005
R1504 VTAIL.n279 VTAIL.n278 9.3005
R1505 VTAIL.n277 VTAIL.n276 9.3005
R1506 VTAIL.n232 VTAIL.n231 9.3005
R1507 VTAIL.n271 VTAIL.n270 9.3005
R1508 VTAIL.n244 VTAIL.n243 9.3005
R1509 VTAIL.n251 VTAIL.n250 9.3005
R1510 VTAIL.n253 VTAIL.n252 9.3005
R1511 VTAIL.n240 VTAIL.n239 9.3005
R1512 VTAIL.n259 VTAIL.n258 9.3005
R1513 VTAIL.n261 VTAIL.n260 9.3005
R1514 VTAIL.n262 VTAIL.n235 9.3005
R1515 VTAIL.n269 VTAIL.n268 9.3005
R1516 VTAIL.n224 VTAIL.n223 9.3005
R1517 VTAIL.n71 VTAIL.n70 9.3005
R1518 VTAIL.n65 VTAIL.n64 9.3005
R1519 VTAIL.n63 VTAIL.n62 9.3005
R1520 VTAIL.n6 VTAIL.n5 9.3005
R1521 VTAIL.n57 VTAIL.n56 9.3005
R1522 VTAIL.n55 VTAIL.n54 9.3005
R1523 VTAIL.n10 VTAIL.n9 9.3005
R1524 VTAIL.n49 VTAIL.n48 9.3005
R1525 VTAIL.n22 VTAIL.n21 9.3005
R1526 VTAIL.n29 VTAIL.n28 9.3005
R1527 VTAIL.n31 VTAIL.n30 9.3005
R1528 VTAIL.n18 VTAIL.n17 9.3005
R1529 VTAIL.n37 VTAIL.n36 9.3005
R1530 VTAIL.n39 VTAIL.n38 9.3005
R1531 VTAIL.n40 VTAIL.n13 9.3005
R1532 VTAIL.n47 VTAIL.n46 9.3005
R1533 VTAIL.n2 VTAIL.n1 9.3005
R1534 VTAIL.n172 VTAIL.n171 9.3005
R1535 VTAIL.n179 VTAIL.n178 9.3005
R1536 VTAIL.n181 VTAIL.n180 9.3005
R1537 VTAIL.n168 VTAIL.n167 9.3005
R1538 VTAIL.n187 VTAIL.n186 9.3005
R1539 VTAIL.n189 VTAIL.n188 9.3005
R1540 VTAIL.n163 VTAIL.n161 9.3005
R1541 VTAIL.n195 VTAIL.n194 9.3005
R1542 VTAIL.n219 VTAIL.n218 9.3005
R1543 VTAIL.n150 VTAIL.n149 9.3005
R1544 VTAIL.n213 VTAIL.n212 9.3005
R1545 VTAIL.n211 VTAIL.n210 9.3005
R1546 VTAIL.n154 VTAIL.n153 9.3005
R1547 VTAIL.n205 VTAIL.n204 9.3005
R1548 VTAIL.n203 VTAIL.n202 9.3005
R1549 VTAIL.n158 VTAIL.n157 9.3005
R1550 VTAIL.n197 VTAIL.n196 9.3005
R1551 VTAIL.n98 VTAIL.n97 9.3005
R1552 VTAIL.n105 VTAIL.n104 9.3005
R1553 VTAIL.n107 VTAIL.n106 9.3005
R1554 VTAIL.n94 VTAIL.n93 9.3005
R1555 VTAIL.n113 VTAIL.n112 9.3005
R1556 VTAIL.n115 VTAIL.n114 9.3005
R1557 VTAIL.n89 VTAIL.n87 9.3005
R1558 VTAIL.n121 VTAIL.n120 9.3005
R1559 VTAIL.n145 VTAIL.n144 9.3005
R1560 VTAIL.n76 VTAIL.n75 9.3005
R1561 VTAIL.n139 VTAIL.n138 9.3005
R1562 VTAIL.n137 VTAIL.n136 9.3005
R1563 VTAIL.n80 VTAIL.n79 9.3005
R1564 VTAIL.n131 VTAIL.n130 9.3005
R1565 VTAIL.n129 VTAIL.n128 9.3005
R1566 VTAIL.n84 VTAIL.n83 9.3005
R1567 VTAIL.n123 VTAIL.n122 9.3005
R1568 VTAIL.n253 VTAIL.n242 8.92171
R1569 VTAIL.n284 VTAIL.n226 8.92171
R1570 VTAIL.n31 VTAIL.n20 8.92171
R1571 VTAIL.n62 VTAIL.n4 8.92171
R1572 VTAIL.n210 VTAIL.n152 8.92171
R1573 VTAIL.n181 VTAIL.n170 8.92171
R1574 VTAIL.n136 VTAIL.n78 8.92171
R1575 VTAIL.n107 VTAIL.n96 8.92171
R1576 VTAIL.n250 VTAIL.n249 8.14595
R1577 VTAIL.n288 VTAIL.n287 8.14595
R1578 VTAIL.n28 VTAIL.n27 8.14595
R1579 VTAIL.n66 VTAIL.n65 8.14595
R1580 VTAIL.n214 VTAIL.n213 8.14595
R1581 VTAIL.n178 VTAIL.n177 8.14595
R1582 VTAIL.n140 VTAIL.n139 8.14595
R1583 VTAIL.n104 VTAIL.n103 8.14595
R1584 VTAIL.n246 VTAIL.n244 7.3702
R1585 VTAIL.n291 VTAIL.n224 7.3702
R1586 VTAIL.n294 VTAIL.n222 7.3702
R1587 VTAIL.n24 VTAIL.n22 7.3702
R1588 VTAIL.n69 VTAIL.n2 7.3702
R1589 VTAIL.n72 VTAIL.n0 7.3702
R1590 VTAIL.n220 VTAIL.n148 7.3702
R1591 VTAIL.n217 VTAIL.n150 7.3702
R1592 VTAIL.n174 VTAIL.n172 7.3702
R1593 VTAIL.n146 VTAIL.n74 7.3702
R1594 VTAIL.n143 VTAIL.n76 7.3702
R1595 VTAIL.n100 VTAIL.n98 7.3702
R1596 VTAIL.n292 VTAIL.n291 6.59444
R1597 VTAIL.n292 VTAIL.n222 6.59444
R1598 VTAIL.n70 VTAIL.n69 6.59444
R1599 VTAIL.n70 VTAIL.n0 6.59444
R1600 VTAIL.n218 VTAIL.n148 6.59444
R1601 VTAIL.n218 VTAIL.n217 6.59444
R1602 VTAIL.n144 VTAIL.n74 6.59444
R1603 VTAIL.n144 VTAIL.n143 6.59444
R1604 VTAIL.n249 VTAIL.n244 5.81868
R1605 VTAIL.n288 VTAIL.n224 5.81868
R1606 VTAIL.n27 VTAIL.n22 5.81868
R1607 VTAIL.n66 VTAIL.n2 5.81868
R1608 VTAIL.n214 VTAIL.n150 5.81868
R1609 VTAIL.n177 VTAIL.n172 5.81868
R1610 VTAIL.n140 VTAIL.n76 5.81868
R1611 VTAIL.n103 VTAIL.n98 5.81868
R1612 VTAIL.n250 VTAIL.n242 5.04292
R1613 VTAIL.n287 VTAIL.n226 5.04292
R1614 VTAIL.n28 VTAIL.n20 5.04292
R1615 VTAIL.n65 VTAIL.n4 5.04292
R1616 VTAIL.n213 VTAIL.n152 5.04292
R1617 VTAIL.n178 VTAIL.n170 5.04292
R1618 VTAIL.n139 VTAIL.n78 5.04292
R1619 VTAIL.n104 VTAIL.n96 5.04292
R1620 VTAIL.n254 VTAIL.n253 4.26717
R1621 VTAIL.n284 VTAIL.n283 4.26717
R1622 VTAIL.n32 VTAIL.n31 4.26717
R1623 VTAIL.n62 VTAIL.n61 4.26717
R1624 VTAIL.n210 VTAIL.n209 4.26717
R1625 VTAIL.n182 VTAIL.n181 4.26717
R1626 VTAIL.n136 VTAIL.n135 4.26717
R1627 VTAIL.n108 VTAIL.n107 4.26717
R1628 VTAIL.n257 VTAIL.n240 3.49141
R1629 VTAIL.n280 VTAIL.n228 3.49141
R1630 VTAIL.n35 VTAIL.n18 3.49141
R1631 VTAIL.n58 VTAIL.n6 3.49141
R1632 VTAIL.n206 VTAIL.n154 3.49141
R1633 VTAIL.n185 VTAIL.n168 3.49141
R1634 VTAIL.n132 VTAIL.n80 3.49141
R1635 VTAIL.n111 VTAIL.n94 3.49141
R1636 VTAIL.n245 VTAIL.n243 2.84303
R1637 VTAIL.n23 VTAIL.n21 2.84303
R1638 VTAIL.n173 VTAIL.n171 2.84303
R1639 VTAIL.n99 VTAIL.n97 2.84303
R1640 VTAIL.n258 VTAIL.n238 2.71565
R1641 VTAIL.n279 VTAIL.n230 2.71565
R1642 VTAIL.n36 VTAIL.n16 2.71565
R1643 VTAIL.n57 VTAIL.n8 2.71565
R1644 VTAIL.n205 VTAIL.n156 2.71565
R1645 VTAIL.n186 VTAIL.n166 2.71565
R1646 VTAIL.n131 VTAIL.n82 2.71565
R1647 VTAIL.n112 VTAIL.n92 2.71565
R1648 VTAIL.n263 VTAIL.n261 1.93989
R1649 VTAIL.n276 VTAIL.n275 1.93989
R1650 VTAIL.n41 VTAIL.n39 1.93989
R1651 VTAIL.n54 VTAIL.n53 1.93989
R1652 VTAIL.n202 VTAIL.n201 1.93989
R1653 VTAIL.n190 VTAIL.n189 1.93989
R1654 VTAIL.n128 VTAIL.n127 1.93989
R1655 VTAIL.n116 VTAIL.n115 1.93989
R1656 VTAIL.n221 VTAIL.n147 1.64705
R1657 VTAIL.n262 VTAIL.n236 1.16414
R1658 VTAIL.n272 VTAIL.n232 1.16414
R1659 VTAIL.n40 VTAIL.n14 1.16414
R1660 VTAIL.n50 VTAIL.n10 1.16414
R1661 VTAIL.n198 VTAIL.n158 1.16414
R1662 VTAIL.n193 VTAIL.n163 1.16414
R1663 VTAIL.n124 VTAIL.n84 1.16414
R1664 VTAIL.n119 VTAIL.n89 1.16414
R1665 VTAIL VTAIL.n73 1.11688
R1666 VTAIL VTAIL.n295 0.530672
R1667 VTAIL.n268 VTAIL.n267 0.388379
R1668 VTAIL.n271 VTAIL.n234 0.388379
R1669 VTAIL.n46 VTAIL.n45 0.388379
R1670 VTAIL.n49 VTAIL.n12 0.388379
R1671 VTAIL.n197 VTAIL.n160 0.388379
R1672 VTAIL.n194 VTAIL.n162 0.388379
R1673 VTAIL.n123 VTAIL.n86 0.388379
R1674 VTAIL.n120 VTAIL.n88 0.388379
R1675 VTAIL.n251 VTAIL.n243 0.155672
R1676 VTAIL.n252 VTAIL.n251 0.155672
R1677 VTAIL.n252 VTAIL.n239 0.155672
R1678 VTAIL.n259 VTAIL.n239 0.155672
R1679 VTAIL.n260 VTAIL.n259 0.155672
R1680 VTAIL.n260 VTAIL.n235 0.155672
R1681 VTAIL.n269 VTAIL.n235 0.155672
R1682 VTAIL.n270 VTAIL.n269 0.155672
R1683 VTAIL.n270 VTAIL.n231 0.155672
R1684 VTAIL.n277 VTAIL.n231 0.155672
R1685 VTAIL.n278 VTAIL.n277 0.155672
R1686 VTAIL.n278 VTAIL.n227 0.155672
R1687 VTAIL.n285 VTAIL.n227 0.155672
R1688 VTAIL.n286 VTAIL.n285 0.155672
R1689 VTAIL.n286 VTAIL.n223 0.155672
R1690 VTAIL.n293 VTAIL.n223 0.155672
R1691 VTAIL.n29 VTAIL.n21 0.155672
R1692 VTAIL.n30 VTAIL.n29 0.155672
R1693 VTAIL.n30 VTAIL.n17 0.155672
R1694 VTAIL.n37 VTAIL.n17 0.155672
R1695 VTAIL.n38 VTAIL.n37 0.155672
R1696 VTAIL.n38 VTAIL.n13 0.155672
R1697 VTAIL.n47 VTAIL.n13 0.155672
R1698 VTAIL.n48 VTAIL.n47 0.155672
R1699 VTAIL.n48 VTAIL.n9 0.155672
R1700 VTAIL.n55 VTAIL.n9 0.155672
R1701 VTAIL.n56 VTAIL.n55 0.155672
R1702 VTAIL.n56 VTAIL.n5 0.155672
R1703 VTAIL.n63 VTAIL.n5 0.155672
R1704 VTAIL.n64 VTAIL.n63 0.155672
R1705 VTAIL.n64 VTAIL.n1 0.155672
R1706 VTAIL.n71 VTAIL.n1 0.155672
R1707 VTAIL.n219 VTAIL.n149 0.155672
R1708 VTAIL.n212 VTAIL.n149 0.155672
R1709 VTAIL.n212 VTAIL.n211 0.155672
R1710 VTAIL.n211 VTAIL.n153 0.155672
R1711 VTAIL.n204 VTAIL.n153 0.155672
R1712 VTAIL.n204 VTAIL.n203 0.155672
R1713 VTAIL.n203 VTAIL.n157 0.155672
R1714 VTAIL.n196 VTAIL.n157 0.155672
R1715 VTAIL.n196 VTAIL.n195 0.155672
R1716 VTAIL.n195 VTAIL.n161 0.155672
R1717 VTAIL.n188 VTAIL.n161 0.155672
R1718 VTAIL.n188 VTAIL.n187 0.155672
R1719 VTAIL.n187 VTAIL.n167 0.155672
R1720 VTAIL.n180 VTAIL.n167 0.155672
R1721 VTAIL.n180 VTAIL.n179 0.155672
R1722 VTAIL.n179 VTAIL.n171 0.155672
R1723 VTAIL.n145 VTAIL.n75 0.155672
R1724 VTAIL.n138 VTAIL.n75 0.155672
R1725 VTAIL.n138 VTAIL.n137 0.155672
R1726 VTAIL.n137 VTAIL.n79 0.155672
R1727 VTAIL.n130 VTAIL.n79 0.155672
R1728 VTAIL.n130 VTAIL.n129 0.155672
R1729 VTAIL.n129 VTAIL.n83 0.155672
R1730 VTAIL.n122 VTAIL.n83 0.155672
R1731 VTAIL.n122 VTAIL.n121 0.155672
R1732 VTAIL.n121 VTAIL.n87 0.155672
R1733 VTAIL.n114 VTAIL.n87 0.155672
R1734 VTAIL.n114 VTAIL.n113 0.155672
R1735 VTAIL.n113 VTAIL.n93 0.155672
R1736 VTAIL.n106 VTAIL.n93 0.155672
R1737 VTAIL.n106 VTAIL.n105 0.155672
R1738 VTAIL.n105 VTAIL.n97 0.155672
R1739 VDD1.n68 VDD1.n0 289.615
R1740 VDD1.n141 VDD1.n73 289.615
R1741 VDD1.n69 VDD1.n68 185
R1742 VDD1.n67 VDD1.n66 185
R1743 VDD1.n4 VDD1.n3 185
R1744 VDD1.n61 VDD1.n60 185
R1745 VDD1.n59 VDD1.n58 185
R1746 VDD1.n8 VDD1.n7 185
R1747 VDD1.n53 VDD1.n52 185
R1748 VDD1.n51 VDD1.n50 185
R1749 VDD1.n12 VDD1.n11 185
R1750 VDD1.n16 VDD1.n14 185
R1751 VDD1.n45 VDD1.n44 185
R1752 VDD1.n43 VDD1.n42 185
R1753 VDD1.n18 VDD1.n17 185
R1754 VDD1.n37 VDD1.n36 185
R1755 VDD1.n35 VDD1.n34 185
R1756 VDD1.n22 VDD1.n21 185
R1757 VDD1.n29 VDD1.n28 185
R1758 VDD1.n27 VDD1.n26 185
R1759 VDD1.n98 VDD1.n97 185
R1760 VDD1.n100 VDD1.n99 185
R1761 VDD1.n93 VDD1.n92 185
R1762 VDD1.n106 VDD1.n105 185
R1763 VDD1.n108 VDD1.n107 185
R1764 VDD1.n89 VDD1.n88 185
R1765 VDD1.n115 VDD1.n114 185
R1766 VDD1.n116 VDD1.n87 185
R1767 VDD1.n118 VDD1.n117 185
R1768 VDD1.n85 VDD1.n84 185
R1769 VDD1.n124 VDD1.n123 185
R1770 VDD1.n126 VDD1.n125 185
R1771 VDD1.n81 VDD1.n80 185
R1772 VDD1.n132 VDD1.n131 185
R1773 VDD1.n134 VDD1.n133 185
R1774 VDD1.n77 VDD1.n76 185
R1775 VDD1.n140 VDD1.n139 185
R1776 VDD1.n142 VDD1.n141 185
R1777 VDD1.n25 VDD1.t0 149.524
R1778 VDD1.n96 VDD1.t1 149.524
R1779 VDD1.n68 VDD1.n67 104.615
R1780 VDD1.n67 VDD1.n3 104.615
R1781 VDD1.n60 VDD1.n3 104.615
R1782 VDD1.n60 VDD1.n59 104.615
R1783 VDD1.n59 VDD1.n7 104.615
R1784 VDD1.n52 VDD1.n7 104.615
R1785 VDD1.n52 VDD1.n51 104.615
R1786 VDD1.n51 VDD1.n11 104.615
R1787 VDD1.n16 VDD1.n11 104.615
R1788 VDD1.n44 VDD1.n16 104.615
R1789 VDD1.n44 VDD1.n43 104.615
R1790 VDD1.n43 VDD1.n17 104.615
R1791 VDD1.n36 VDD1.n17 104.615
R1792 VDD1.n36 VDD1.n35 104.615
R1793 VDD1.n35 VDD1.n21 104.615
R1794 VDD1.n28 VDD1.n21 104.615
R1795 VDD1.n28 VDD1.n27 104.615
R1796 VDD1.n99 VDD1.n98 104.615
R1797 VDD1.n99 VDD1.n92 104.615
R1798 VDD1.n106 VDD1.n92 104.615
R1799 VDD1.n107 VDD1.n106 104.615
R1800 VDD1.n107 VDD1.n88 104.615
R1801 VDD1.n115 VDD1.n88 104.615
R1802 VDD1.n116 VDD1.n115 104.615
R1803 VDD1.n117 VDD1.n116 104.615
R1804 VDD1.n117 VDD1.n84 104.615
R1805 VDD1.n124 VDD1.n84 104.615
R1806 VDD1.n125 VDD1.n124 104.615
R1807 VDD1.n125 VDD1.n80 104.615
R1808 VDD1.n132 VDD1.n80 104.615
R1809 VDD1.n133 VDD1.n132 104.615
R1810 VDD1.n133 VDD1.n76 104.615
R1811 VDD1.n140 VDD1.n76 104.615
R1812 VDD1.n141 VDD1.n140 104.615
R1813 VDD1 VDD1.n145 89.4256
R1814 VDD1.n27 VDD1.t0 52.3082
R1815 VDD1.n98 VDD1.t1 52.3082
R1816 VDD1 VDD1.n72 48.9289
R1817 VDD1.n14 VDD1.n12 13.1884
R1818 VDD1.n118 VDD1.n85 13.1884
R1819 VDD1.n50 VDD1.n49 12.8005
R1820 VDD1.n46 VDD1.n45 12.8005
R1821 VDD1.n119 VDD1.n87 12.8005
R1822 VDD1.n123 VDD1.n122 12.8005
R1823 VDD1.n53 VDD1.n10 12.0247
R1824 VDD1.n42 VDD1.n15 12.0247
R1825 VDD1.n114 VDD1.n113 12.0247
R1826 VDD1.n126 VDD1.n83 12.0247
R1827 VDD1.n54 VDD1.n8 11.249
R1828 VDD1.n41 VDD1.n18 11.249
R1829 VDD1.n112 VDD1.n89 11.249
R1830 VDD1.n127 VDD1.n81 11.249
R1831 VDD1.n58 VDD1.n57 10.4732
R1832 VDD1.n38 VDD1.n37 10.4732
R1833 VDD1.n109 VDD1.n108 10.4732
R1834 VDD1.n131 VDD1.n130 10.4732
R1835 VDD1.n26 VDD1.n25 10.2747
R1836 VDD1.n97 VDD1.n96 10.2747
R1837 VDD1.n61 VDD1.n6 9.69747
R1838 VDD1.n34 VDD1.n20 9.69747
R1839 VDD1.n105 VDD1.n91 9.69747
R1840 VDD1.n134 VDD1.n79 9.69747
R1841 VDD1.n72 VDD1.n71 9.45567
R1842 VDD1.n145 VDD1.n144 9.45567
R1843 VDD1.n24 VDD1.n23 9.3005
R1844 VDD1.n31 VDD1.n30 9.3005
R1845 VDD1.n33 VDD1.n32 9.3005
R1846 VDD1.n20 VDD1.n19 9.3005
R1847 VDD1.n39 VDD1.n38 9.3005
R1848 VDD1.n41 VDD1.n40 9.3005
R1849 VDD1.n15 VDD1.n13 9.3005
R1850 VDD1.n47 VDD1.n46 9.3005
R1851 VDD1.n71 VDD1.n70 9.3005
R1852 VDD1.n2 VDD1.n1 9.3005
R1853 VDD1.n65 VDD1.n64 9.3005
R1854 VDD1.n63 VDD1.n62 9.3005
R1855 VDD1.n6 VDD1.n5 9.3005
R1856 VDD1.n57 VDD1.n56 9.3005
R1857 VDD1.n55 VDD1.n54 9.3005
R1858 VDD1.n10 VDD1.n9 9.3005
R1859 VDD1.n49 VDD1.n48 9.3005
R1860 VDD1.n144 VDD1.n143 9.3005
R1861 VDD1.n138 VDD1.n137 9.3005
R1862 VDD1.n136 VDD1.n135 9.3005
R1863 VDD1.n79 VDD1.n78 9.3005
R1864 VDD1.n130 VDD1.n129 9.3005
R1865 VDD1.n128 VDD1.n127 9.3005
R1866 VDD1.n83 VDD1.n82 9.3005
R1867 VDD1.n122 VDD1.n121 9.3005
R1868 VDD1.n95 VDD1.n94 9.3005
R1869 VDD1.n102 VDD1.n101 9.3005
R1870 VDD1.n104 VDD1.n103 9.3005
R1871 VDD1.n91 VDD1.n90 9.3005
R1872 VDD1.n110 VDD1.n109 9.3005
R1873 VDD1.n112 VDD1.n111 9.3005
R1874 VDD1.n113 VDD1.n86 9.3005
R1875 VDD1.n120 VDD1.n119 9.3005
R1876 VDD1.n75 VDD1.n74 9.3005
R1877 VDD1.n62 VDD1.n4 8.92171
R1878 VDD1.n33 VDD1.n22 8.92171
R1879 VDD1.n104 VDD1.n93 8.92171
R1880 VDD1.n135 VDD1.n77 8.92171
R1881 VDD1.n66 VDD1.n65 8.14595
R1882 VDD1.n30 VDD1.n29 8.14595
R1883 VDD1.n101 VDD1.n100 8.14595
R1884 VDD1.n139 VDD1.n138 8.14595
R1885 VDD1.n72 VDD1.n0 7.3702
R1886 VDD1.n69 VDD1.n2 7.3702
R1887 VDD1.n26 VDD1.n24 7.3702
R1888 VDD1.n97 VDD1.n95 7.3702
R1889 VDD1.n142 VDD1.n75 7.3702
R1890 VDD1.n145 VDD1.n73 7.3702
R1891 VDD1.n70 VDD1.n0 6.59444
R1892 VDD1.n70 VDD1.n69 6.59444
R1893 VDD1.n143 VDD1.n142 6.59444
R1894 VDD1.n143 VDD1.n73 6.59444
R1895 VDD1.n66 VDD1.n2 5.81868
R1896 VDD1.n29 VDD1.n24 5.81868
R1897 VDD1.n100 VDD1.n95 5.81868
R1898 VDD1.n139 VDD1.n75 5.81868
R1899 VDD1.n65 VDD1.n4 5.04292
R1900 VDD1.n30 VDD1.n22 5.04292
R1901 VDD1.n101 VDD1.n93 5.04292
R1902 VDD1.n138 VDD1.n77 5.04292
R1903 VDD1.n62 VDD1.n61 4.26717
R1904 VDD1.n34 VDD1.n33 4.26717
R1905 VDD1.n105 VDD1.n104 4.26717
R1906 VDD1.n135 VDD1.n134 4.26717
R1907 VDD1.n58 VDD1.n6 3.49141
R1908 VDD1.n37 VDD1.n20 3.49141
R1909 VDD1.n108 VDD1.n91 3.49141
R1910 VDD1.n131 VDD1.n79 3.49141
R1911 VDD1.n25 VDD1.n23 2.84303
R1912 VDD1.n96 VDD1.n94 2.84303
R1913 VDD1.n57 VDD1.n8 2.71565
R1914 VDD1.n38 VDD1.n18 2.71565
R1915 VDD1.n109 VDD1.n89 2.71565
R1916 VDD1.n130 VDD1.n81 2.71565
R1917 VDD1.n54 VDD1.n53 1.93989
R1918 VDD1.n42 VDD1.n41 1.93989
R1919 VDD1.n114 VDD1.n112 1.93989
R1920 VDD1.n127 VDD1.n126 1.93989
R1921 VDD1.n50 VDD1.n10 1.16414
R1922 VDD1.n45 VDD1.n15 1.16414
R1923 VDD1.n113 VDD1.n87 1.16414
R1924 VDD1.n123 VDD1.n83 1.16414
R1925 VDD1.n49 VDD1.n12 0.388379
R1926 VDD1.n46 VDD1.n14 0.388379
R1927 VDD1.n119 VDD1.n118 0.388379
R1928 VDD1.n122 VDD1.n85 0.388379
R1929 VDD1.n71 VDD1.n1 0.155672
R1930 VDD1.n64 VDD1.n1 0.155672
R1931 VDD1.n64 VDD1.n63 0.155672
R1932 VDD1.n63 VDD1.n5 0.155672
R1933 VDD1.n56 VDD1.n5 0.155672
R1934 VDD1.n56 VDD1.n55 0.155672
R1935 VDD1.n55 VDD1.n9 0.155672
R1936 VDD1.n48 VDD1.n9 0.155672
R1937 VDD1.n48 VDD1.n47 0.155672
R1938 VDD1.n47 VDD1.n13 0.155672
R1939 VDD1.n40 VDD1.n13 0.155672
R1940 VDD1.n40 VDD1.n39 0.155672
R1941 VDD1.n39 VDD1.n19 0.155672
R1942 VDD1.n32 VDD1.n19 0.155672
R1943 VDD1.n32 VDD1.n31 0.155672
R1944 VDD1.n31 VDD1.n23 0.155672
R1945 VDD1.n102 VDD1.n94 0.155672
R1946 VDD1.n103 VDD1.n102 0.155672
R1947 VDD1.n103 VDD1.n90 0.155672
R1948 VDD1.n110 VDD1.n90 0.155672
R1949 VDD1.n111 VDD1.n110 0.155672
R1950 VDD1.n111 VDD1.n86 0.155672
R1951 VDD1.n120 VDD1.n86 0.155672
R1952 VDD1.n121 VDD1.n120 0.155672
R1953 VDD1.n121 VDD1.n82 0.155672
R1954 VDD1.n128 VDD1.n82 0.155672
R1955 VDD1.n129 VDD1.n128 0.155672
R1956 VDD1.n129 VDD1.n78 0.155672
R1957 VDD1.n136 VDD1.n78 0.155672
R1958 VDD1.n137 VDD1.n136 0.155672
R1959 VDD1.n137 VDD1.n74 0.155672
R1960 VDD1.n144 VDD1.n74 0.155672
R1961 VN VN.t1 230.417
R1962 VN VN.t0 185.37
R1963 VDD2.n141 VDD2.n73 289.615
R1964 VDD2.n68 VDD2.n0 289.615
R1965 VDD2.n142 VDD2.n141 185
R1966 VDD2.n140 VDD2.n139 185
R1967 VDD2.n77 VDD2.n76 185
R1968 VDD2.n134 VDD2.n133 185
R1969 VDD2.n132 VDD2.n131 185
R1970 VDD2.n81 VDD2.n80 185
R1971 VDD2.n126 VDD2.n125 185
R1972 VDD2.n124 VDD2.n123 185
R1973 VDD2.n85 VDD2.n84 185
R1974 VDD2.n89 VDD2.n87 185
R1975 VDD2.n118 VDD2.n117 185
R1976 VDD2.n116 VDD2.n115 185
R1977 VDD2.n91 VDD2.n90 185
R1978 VDD2.n110 VDD2.n109 185
R1979 VDD2.n108 VDD2.n107 185
R1980 VDD2.n95 VDD2.n94 185
R1981 VDD2.n102 VDD2.n101 185
R1982 VDD2.n100 VDD2.n99 185
R1983 VDD2.n25 VDD2.n24 185
R1984 VDD2.n27 VDD2.n26 185
R1985 VDD2.n20 VDD2.n19 185
R1986 VDD2.n33 VDD2.n32 185
R1987 VDD2.n35 VDD2.n34 185
R1988 VDD2.n16 VDD2.n15 185
R1989 VDD2.n42 VDD2.n41 185
R1990 VDD2.n43 VDD2.n14 185
R1991 VDD2.n45 VDD2.n44 185
R1992 VDD2.n12 VDD2.n11 185
R1993 VDD2.n51 VDD2.n50 185
R1994 VDD2.n53 VDD2.n52 185
R1995 VDD2.n8 VDD2.n7 185
R1996 VDD2.n59 VDD2.n58 185
R1997 VDD2.n61 VDD2.n60 185
R1998 VDD2.n4 VDD2.n3 185
R1999 VDD2.n67 VDD2.n66 185
R2000 VDD2.n69 VDD2.n68 185
R2001 VDD2.n98 VDD2.t0 149.524
R2002 VDD2.n23 VDD2.t1 149.524
R2003 VDD2.n141 VDD2.n140 104.615
R2004 VDD2.n140 VDD2.n76 104.615
R2005 VDD2.n133 VDD2.n76 104.615
R2006 VDD2.n133 VDD2.n132 104.615
R2007 VDD2.n132 VDD2.n80 104.615
R2008 VDD2.n125 VDD2.n80 104.615
R2009 VDD2.n125 VDD2.n124 104.615
R2010 VDD2.n124 VDD2.n84 104.615
R2011 VDD2.n89 VDD2.n84 104.615
R2012 VDD2.n117 VDD2.n89 104.615
R2013 VDD2.n117 VDD2.n116 104.615
R2014 VDD2.n116 VDD2.n90 104.615
R2015 VDD2.n109 VDD2.n90 104.615
R2016 VDD2.n109 VDD2.n108 104.615
R2017 VDD2.n108 VDD2.n94 104.615
R2018 VDD2.n101 VDD2.n94 104.615
R2019 VDD2.n101 VDD2.n100 104.615
R2020 VDD2.n26 VDD2.n25 104.615
R2021 VDD2.n26 VDD2.n19 104.615
R2022 VDD2.n33 VDD2.n19 104.615
R2023 VDD2.n34 VDD2.n33 104.615
R2024 VDD2.n34 VDD2.n15 104.615
R2025 VDD2.n42 VDD2.n15 104.615
R2026 VDD2.n43 VDD2.n42 104.615
R2027 VDD2.n44 VDD2.n43 104.615
R2028 VDD2.n44 VDD2.n11 104.615
R2029 VDD2.n51 VDD2.n11 104.615
R2030 VDD2.n52 VDD2.n51 104.615
R2031 VDD2.n52 VDD2.n7 104.615
R2032 VDD2.n59 VDD2.n7 104.615
R2033 VDD2.n60 VDD2.n59 104.615
R2034 VDD2.n60 VDD2.n3 104.615
R2035 VDD2.n67 VDD2.n3 104.615
R2036 VDD2.n68 VDD2.n67 104.615
R2037 VDD2.n146 VDD2.n72 88.3125
R2038 VDD2.n100 VDD2.t0 52.3082
R2039 VDD2.n25 VDD2.t1 52.3082
R2040 VDD2.n146 VDD2.n145 48.2823
R2041 VDD2.n87 VDD2.n85 13.1884
R2042 VDD2.n45 VDD2.n12 13.1884
R2043 VDD2.n123 VDD2.n122 12.8005
R2044 VDD2.n119 VDD2.n118 12.8005
R2045 VDD2.n46 VDD2.n14 12.8005
R2046 VDD2.n50 VDD2.n49 12.8005
R2047 VDD2.n126 VDD2.n83 12.0247
R2048 VDD2.n115 VDD2.n88 12.0247
R2049 VDD2.n41 VDD2.n40 12.0247
R2050 VDD2.n53 VDD2.n10 12.0247
R2051 VDD2.n127 VDD2.n81 11.249
R2052 VDD2.n114 VDD2.n91 11.249
R2053 VDD2.n39 VDD2.n16 11.249
R2054 VDD2.n54 VDD2.n8 11.249
R2055 VDD2.n131 VDD2.n130 10.4732
R2056 VDD2.n111 VDD2.n110 10.4732
R2057 VDD2.n36 VDD2.n35 10.4732
R2058 VDD2.n58 VDD2.n57 10.4732
R2059 VDD2.n99 VDD2.n98 10.2747
R2060 VDD2.n24 VDD2.n23 10.2747
R2061 VDD2.n134 VDD2.n79 9.69747
R2062 VDD2.n107 VDD2.n93 9.69747
R2063 VDD2.n32 VDD2.n18 9.69747
R2064 VDD2.n61 VDD2.n6 9.69747
R2065 VDD2.n145 VDD2.n144 9.45567
R2066 VDD2.n72 VDD2.n71 9.45567
R2067 VDD2.n97 VDD2.n96 9.3005
R2068 VDD2.n104 VDD2.n103 9.3005
R2069 VDD2.n106 VDD2.n105 9.3005
R2070 VDD2.n93 VDD2.n92 9.3005
R2071 VDD2.n112 VDD2.n111 9.3005
R2072 VDD2.n114 VDD2.n113 9.3005
R2073 VDD2.n88 VDD2.n86 9.3005
R2074 VDD2.n120 VDD2.n119 9.3005
R2075 VDD2.n144 VDD2.n143 9.3005
R2076 VDD2.n75 VDD2.n74 9.3005
R2077 VDD2.n138 VDD2.n137 9.3005
R2078 VDD2.n136 VDD2.n135 9.3005
R2079 VDD2.n79 VDD2.n78 9.3005
R2080 VDD2.n130 VDD2.n129 9.3005
R2081 VDD2.n128 VDD2.n127 9.3005
R2082 VDD2.n83 VDD2.n82 9.3005
R2083 VDD2.n122 VDD2.n121 9.3005
R2084 VDD2.n71 VDD2.n70 9.3005
R2085 VDD2.n65 VDD2.n64 9.3005
R2086 VDD2.n63 VDD2.n62 9.3005
R2087 VDD2.n6 VDD2.n5 9.3005
R2088 VDD2.n57 VDD2.n56 9.3005
R2089 VDD2.n55 VDD2.n54 9.3005
R2090 VDD2.n10 VDD2.n9 9.3005
R2091 VDD2.n49 VDD2.n48 9.3005
R2092 VDD2.n22 VDD2.n21 9.3005
R2093 VDD2.n29 VDD2.n28 9.3005
R2094 VDD2.n31 VDD2.n30 9.3005
R2095 VDD2.n18 VDD2.n17 9.3005
R2096 VDD2.n37 VDD2.n36 9.3005
R2097 VDD2.n39 VDD2.n38 9.3005
R2098 VDD2.n40 VDD2.n13 9.3005
R2099 VDD2.n47 VDD2.n46 9.3005
R2100 VDD2.n2 VDD2.n1 9.3005
R2101 VDD2.n135 VDD2.n77 8.92171
R2102 VDD2.n106 VDD2.n95 8.92171
R2103 VDD2.n31 VDD2.n20 8.92171
R2104 VDD2.n62 VDD2.n4 8.92171
R2105 VDD2.n139 VDD2.n138 8.14595
R2106 VDD2.n103 VDD2.n102 8.14595
R2107 VDD2.n28 VDD2.n27 8.14595
R2108 VDD2.n66 VDD2.n65 8.14595
R2109 VDD2.n145 VDD2.n73 7.3702
R2110 VDD2.n142 VDD2.n75 7.3702
R2111 VDD2.n99 VDD2.n97 7.3702
R2112 VDD2.n24 VDD2.n22 7.3702
R2113 VDD2.n69 VDD2.n2 7.3702
R2114 VDD2.n72 VDD2.n0 7.3702
R2115 VDD2.n143 VDD2.n73 6.59444
R2116 VDD2.n143 VDD2.n142 6.59444
R2117 VDD2.n70 VDD2.n69 6.59444
R2118 VDD2.n70 VDD2.n0 6.59444
R2119 VDD2.n139 VDD2.n75 5.81868
R2120 VDD2.n102 VDD2.n97 5.81868
R2121 VDD2.n27 VDD2.n22 5.81868
R2122 VDD2.n66 VDD2.n2 5.81868
R2123 VDD2.n138 VDD2.n77 5.04292
R2124 VDD2.n103 VDD2.n95 5.04292
R2125 VDD2.n28 VDD2.n20 5.04292
R2126 VDD2.n65 VDD2.n4 5.04292
R2127 VDD2.n135 VDD2.n134 4.26717
R2128 VDD2.n107 VDD2.n106 4.26717
R2129 VDD2.n32 VDD2.n31 4.26717
R2130 VDD2.n62 VDD2.n61 4.26717
R2131 VDD2.n131 VDD2.n79 3.49141
R2132 VDD2.n110 VDD2.n93 3.49141
R2133 VDD2.n35 VDD2.n18 3.49141
R2134 VDD2.n58 VDD2.n6 3.49141
R2135 VDD2.n98 VDD2.n96 2.84303
R2136 VDD2.n23 VDD2.n21 2.84303
R2137 VDD2.n130 VDD2.n81 2.71565
R2138 VDD2.n111 VDD2.n91 2.71565
R2139 VDD2.n36 VDD2.n16 2.71565
R2140 VDD2.n57 VDD2.n8 2.71565
R2141 VDD2.n127 VDD2.n126 1.93989
R2142 VDD2.n115 VDD2.n114 1.93989
R2143 VDD2.n41 VDD2.n39 1.93989
R2144 VDD2.n54 VDD2.n53 1.93989
R2145 VDD2.n123 VDD2.n83 1.16414
R2146 VDD2.n118 VDD2.n88 1.16414
R2147 VDD2.n40 VDD2.n14 1.16414
R2148 VDD2.n50 VDD2.n10 1.16414
R2149 VDD2 VDD2.n146 0.647052
R2150 VDD2.n122 VDD2.n85 0.388379
R2151 VDD2.n119 VDD2.n87 0.388379
R2152 VDD2.n46 VDD2.n45 0.388379
R2153 VDD2.n49 VDD2.n12 0.388379
R2154 VDD2.n144 VDD2.n74 0.155672
R2155 VDD2.n137 VDD2.n74 0.155672
R2156 VDD2.n137 VDD2.n136 0.155672
R2157 VDD2.n136 VDD2.n78 0.155672
R2158 VDD2.n129 VDD2.n78 0.155672
R2159 VDD2.n129 VDD2.n128 0.155672
R2160 VDD2.n128 VDD2.n82 0.155672
R2161 VDD2.n121 VDD2.n82 0.155672
R2162 VDD2.n121 VDD2.n120 0.155672
R2163 VDD2.n120 VDD2.n86 0.155672
R2164 VDD2.n113 VDD2.n86 0.155672
R2165 VDD2.n113 VDD2.n112 0.155672
R2166 VDD2.n112 VDD2.n92 0.155672
R2167 VDD2.n105 VDD2.n92 0.155672
R2168 VDD2.n105 VDD2.n104 0.155672
R2169 VDD2.n104 VDD2.n96 0.155672
R2170 VDD2.n29 VDD2.n21 0.155672
R2171 VDD2.n30 VDD2.n29 0.155672
R2172 VDD2.n30 VDD2.n17 0.155672
R2173 VDD2.n37 VDD2.n17 0.155672
R2174 VDD2.n38 VDD2.n37 0.155672
R2175 VDD2.n38 VDD2.n13 0.155672
R2176 VDD2.n47 VDD2.n13 0.155672
R2177 VDD2.n48 VDD2.n47 0.155672
R2178 VDD2.n48 VDD2.n9 0.155672
R2179 VDD2.n55 VDD2.n9 0.155672
R2180 VDD2.n56 VDD2.n55 0.155672
R2181 VDD2.n56 VDD2.n5 0.155672
R2182 VDD2.n63 VDD2.n5 0.155672
R2183 VDD2.n64 VDD2.n63 0.155672
R2184 VDD2.n64 VDD2.n1 0.155672
R2185 VDD2.n71 VDD2.n1 0.155672
C0 VN VP 5.64488f
C1 VTAIL VP 2.65647f
C2 VN VDD2 3.06335f
C3 VN VDD1 0.14803f
C4 VTAIL VDD2 5.50063f
C5 VTAIL VDD1 5.451971f
C6 VP VDD2 0.324804f
C7 VP VDD1 3.2372f
C8 VDD2 VDD1 0.650872f
C9 VTAIL VN 2.64214f
C10 VDD2 B 4.635581f
C11 VDD1 B 7.43492f
C12 VTAIL B 7.90085f
C13 VN B 10.83943f
C14 VP B 6.252493f
C15 VDD2.n0 B 0.029095f
C16 VDD2.n1 B 0.020215f
C17 VDD2.n2 B 0.010862f
C18 VDD2.n3 B 0.025675f
C19 VDD2.n4 B 0.011501f
C20 VDD2.n5 B 0.020215f
C21 VDD2.n6 B 0.010862f
C22 VDD2.n7 B 0.025675f
C23 VDD2.n8 B 0.011501f
C24 VDD2.n9 B 0.020215f
C25 VDD2.n10 B 0.010862f
C26 VDD2.n11 B 0.025675f
C27 VDD2.n12 B 0.011182f
C28 VDD2.n13 B 0.020215f
C29 VDD2.n14 B 0.011501f
C30 VDD2.n15 B 0.025675f
C31 VDD2.n16 B 0.011501f
C32 VDD2.n17 B 0.020215f
C33 VDD2.n18 B 0.010862f
C34 VDD2.n19 B 0.025675f
C35 VDD2.n20 B 0.011501f
C36 VDD2.n21 B 1.15735f
C37 VDD2.n22 B 0.010862f
C38 VDD2.t1 B 0.043529f
C39 VDD2.n23 B 0.157618f
C40 VDD2.n24 B 0.01815f
C41 VDD2.n25 B 0.019256f
C42 VDD2.n26 B 0.025675f
C43 VDD2.n27 B 0.011501f
C44 VDD2.n28 B 0.010862f
C45 VDD2.n29 B 0.020215f
C46 VDD2.n30 B 0.020215f
C47 VDD2.n31 B 0.010862f
C48 VDD2.n32 B 0.011501f
C49 VDD2.n33 B 0.025675f
C50 VDD2.n34 B 0.025675f
C51 VDD2.n35 B 0.011501f
C52 VDD2.n36 B 0.010862f
C53 VDD2.n37 B 0.020215f
C54 VDD2.n38 B 0.020215f
C55 VDD2.n39 B 0.010862f
C56 VDD2.n40 B 0.010862f
C57 VDD2.n41 B 0.011501f
C58 VDD2.n42 B 0.025675f
C59 VDD2.n43 B 0.025675f
C60 VDD2.n44 B 0.025675f
C61 VDD2.n45 B 0.011182f
C62 VDD2.n46 B 0.010862f
C63 VDD2.n47 B 0.020215f
C64 VDD2.n48 B 0.020215f
C65 VDD2.n49 B 0.010862f
C66 VDD2.n50 B 0.011501f
C67 VDD2.n51 B 0.025675f
C68 VDD2.n52 B 0.025675f
C69 VDD2.n53 B 0.011501f
C70 VDD2.n54 B 0.010862f
C71 VDD2.n55 B 0.020215f
C72 VDD2.n56 B 0.020215f
C73 VDD2.n57 B 0.010862f
C74 VDD2.n58 B 0.011501f
C75 VDD2.n59 B 0.025675f
C76 VDD2.n60 B 0.025675f
C77 VDD2.n61 B 0.011501f
C78 VDD2.n62 B 0.010862f
C79 VDD2.n63 B 0.020215f
C80 VDD2.n64 B 0.020215f
C81 VDD2.n65 B 0.010862f
C82 VDD2.n66 B 0.011501f
C83 VDD2.n67 B 0.025675f
C84 VDD2.n68 B 0.056787f
C85 VDD2.n69 B 0.011501f
C86 VDD2.n70 B 0.010862f
C87 VDD2.n71 B 0.045897f
C88 VDD2.n72 B 0.632405f
C89 VDD2.n73 B 0.029095f
C90 VDD2.n74 B 0.020215f
C91 VDD2.n75 B 0.010862f
C92 VDD2.n76 B 0.025675f
C93 VDD2.n77 B 0.011501f
C94 VDD2.n78 B 0.020215f
C95 VDD2.n79 B 0.010862f
C96 VDD2.n80 B 0.025675f
C97 VDD2.n81 B 0.011501f
C98 VDD2.n82 B 0.020215f
C99 VDD2.n83 B 0.010862f
C100 VDD2.n84 B 0.025675f
C101 VDD2.n85 B 0.011182f
C102 VDD2.n86 B 0.020215f
C103 VDD2.n87 B 0.011182f
C104 VDD2.n88 B 0.010862f
C105 VDD2.n89 B 0.025675f
C106 VDD2.n90 B 0.025675f
C107 VDD2.n91 B 0.011501f
C108 VDD2.n92 B 0.020215f
C109 VDD2.n93 B 0.010862f
C110 VDD2.n94 B 0.025675f
C111 VDD2.n95 B 0.011501f
C112 VDD2.n96 B 1.15735f
C113 VDD2.n97 B 0.010862f
C114 VDD2.t0 B 0.043529f
C115 VDD2.n98 B 0.157618f
C116 VDD2.n99 B 0.01815f
C117 VDD2.n100 B 0.019256f
C118 VDD2.n101 B 0.025675f
C119 VDD2.n102 B 0.011501f
C120 VDD2.n103 B 0.010862f
C121 VDD2.n104 B 0.020215f
C122 VDD2.n105 B 0.020215f
C123 VDD2.n106 B 0.010862f
C124 VDD2.n107 B 0.011501f
C125 VDD2.n108 B 0.025675f
C126 VDD2.n109 B 0.025675f
C127 VDD2.n110 B 0.011501f
C128 VDD2.n111 B 0.010862f
C129 VDD2.n112 B 0.020215f
C130 VDD2.n113 B 0.020215f
C131 VDD2.n114 B 0.010862f
C132 VDD2.n115 B 0.011501f
C133 VDD2.n116 B 0.025675f
C134 VDD2.n117 B 0.025675f
C135 VDD2.n118 B 0.011501f
C136 VDD2.n119 B 0.010862f
C137 VDD2.n120 B 0.020215f
C138 VDD2.n121 B 0.020215f
C139 VDD2.n122 B 0.010862f
C140 VDD2.n123 B 0.011501f
C141 VDD2.n124 B 0.025675f
C142 VDD2.n125 B 0.025675f
C143 VDD2.n126 B 0.011501f
C144 VDD2.n127 B 0.010862f
C145 VDD2.n128 B 0.020215f
C146 VDD2.n129 B 0.020215f
C147 VDD2.n130 B 0.010862f
C148 VDD2.n131 B 0.011501f
C149 VDD2.n132 B 0.025675f
C150 VDD2.n133 B 0.025675f
C151 VDD2.n134 B 0.011501f
C152 VDD2.n135 B 0.010862f
C153 VDD2.n136 B 0.020215f
C154 VDD2.n137 B 0.020215f
C155 VDD2.n138 B 0.010862f
C156 VDD2.n139 B 0.011501f
C157 VDD2.n140 B 0.025675f
C158 VDD2.n141 B 0.056787f
C159 VDD2.n142 B 0.011501f
C160 VDD2.n143 B 0.010862f
C161 VDD2.n144 B 0.045897f
C162 VDD2.n145 B 0.045838f
C163 VDD2.n146 B 2.55994f
C164 VN.t0 B 3.13521f
C165 VN.t1 B 3.62436f
C166 VDD1.n0 B 0.02918f
C167 VDD1.n1 B 0.020274f
C168 VDD1.n2 B 0.010894f
C169 VDD1.n3 B 0.02575f
C170 VDD1.n4 B 0.011535f
C171 VDD1.n5 B 0.020274f
C172 VDD1.n6 B 0.010894f
C173 VDD1.n7 B 0.02575f
C174 VDD1.n8 B 0.011535f
C175 VDD1.n9 B 0.020274f
C176 VDD1.n10 B 0.010894f
C177 VDD1.n11 B 0.02575f
C178 VDD1.n12 B 0.011215f
C179 VDD1.n13 B 0.020274f
C180 VDD1.n14 B 0.011215f
C181 VDD1.n15 B 0.010894f
C182 VDD1.n16 B 0.02575f
C183 VDD1.n17 B 0.02575f
C184 VDD1.n18 B 0.011535f
C185 VDD1.n19 B 0.020274f
C186 VDD1.n20 B 0.010894f
C187 VDD1.n21 B 0.02575f
C188 VDD1.n22 B 0.011535f
C189 VDD1.n23 B 1.16073f
C190 VDD1.n24 B 0.010894f
C191 VDD1.t0 B 0.043657f
C192 VDD1.n25 B 0.158079f
C193 VDD1.n26 B 0.018203f
C194 VDD1.n27 B 0.019312f
C195 VDD1.n28 B 0.02575f
C196 VDD1.n29 B 0.011535f
C197 VDD1.n30 B 0.010894f
C198 VDD1.n31 B 0.020274f
C199 VDD1.n32 B 0.020274f
C200 VDD1.n33 B 0.010894f
C201 VDD1.n34 B 0.011535f
C202 VDD1.n35 B 0.02575f
C203 VDD1.n36 B 0.02575f
C204 VDD1.n37 B 0.011535f
C205 VDD1.n38 B 0.010894f
C206 VDD1.n39 B 0.020274f
C207 VDD1.n40 B 0.020274f
C208 VDD1.n41 B 0.010894f
C209 VDD1.n42 B 0.011535f
C210 VDD1.n43 B 0.02575f
C211 VDD1.n44 B 0.02575f
C212 VDD1.n45 B 0.011535f
C213 VDD1.n46 B 0.010894f
C214 VDD1.n47 B 0.020274f
C215 VDD1.n48 B 0.020274f
C216 VDD1.n49 B 0.010894f
C217 VDD1.n50 B 0.011535f
C218 VDD1.n51 B 0.02575f
C219 VDD1.n52 B 0.02575f
C220 VDD1.n53 B 0.011535f
C221 VDD1.n54 B 0.010894f
C222 VDD1.n55 B 0.020274f
C223 VDD1.n56 B 0.020274f
C224 VDD1.n57 B 0.010894f
C225 VDD1.n58 B 0.011535f
C226 VDD1.n59 B 0.02575f
C227 VDD1.n60 B 0.02575f
C228 VDD1.n61 B 0.011535f
C229 VDD1.n62 B 0.010894f
C230 VDD1.n63 B 0.020274f
C231 VDD1.n64 B 0.020274f
C232 VDD1.n65 B 0.010894f
C233 VDD1.n66 B 0.011535f
C234 VDD1.n67 B 0.02575f
C235 VDD1.n68 B 0.056953f
C236 VDD1.n69 B 0.011535f
C237 VDD1.n70 B 0.010894f
C238 VDD1.n71 B 0.04603f
C239 VDD1.n72 B 0.047039f
C240 VDD1.n73 B 0.02918f
C241 VDD1.n74 B 0.020274f
C242 VDD1.n75 B 0.010894f
C243 VDD1.n76 B 0.02575f
C244 VDD1.n77 B 0.011535f
C245 VDD1.n78 B 0.020274f
C246 VDD1.n79 B 0.010894f
C247 VDD1.n80 B 0.02575f
C248 VDD1.n81 B 0.011535f
C249 VDD1.n82 B 0.020274f
C250 VDD1.n83 B 0.010894f
C251 VDD1.n84 B 0.02575f
C252 VDD1.n85 B 0.011215f
C253 VDD1.n86 B 0.020274f
C254 VDD1.n87 B 0.011535f
C255 VDD1.n88 B 0.02575f
C256 VDD1.n89 B 0.011535f
C257 VDD1.n90 B 0.020274f
C258 VDD1.n91 B 0.010894f
C259 VDD1.n92 B 0.02575f
C260 VDD1.n93 B 0.011535f
C261 VDD1.n94 B 1.16073f
C262 VDD1.n95 B 0.010894f
C263 VDD1.t1 B 0.043657f
C264 VDD1.n96 B 0.158079f
C265 VDD1.n97 B 0.018203f
C266 VDD1.n98 B 0.019312f
C267 VDD1.n99 B 0.02575f
C268 VDD1.n100 B 0.011535f
C269 VDD1.n101 B 0.010894f
C270 VDD1.n102 B 0.020274f
C271 VDD1.n103 B 0.020274f
C272 VDD1.n104 B 0.010894f
C273 VDD1.n105 B 0.011535f
C274 VDD1.n106 B 0.02575f
C275 VDD1.n107 B 0.02575f
C276 VDD1.n108 B 0.011535f
C277 VDD1.n109 B 0.010894f
C278 VDD1.n110 B 0.020274f
C279 VDD1.n111 B 0.020274f
C280 VDD1.n112 B 0.010894f
C281 VDD1.n113 B 0.010894f
C282 VDD1.n114 B 0.011535f
C283 VDD1.n115 B 0.02575f
C284 VDD1.n116 B 0.02575f
C285 VDD1.n117 B 0.02575f
C286 VDD1.n118 B 0.011215f
C287 VDD1.n119 B 0.010894f
C288 VDD1.n120 B 0.020274f
C289 VDD1.n121 B 0.020274f
C290 VDD1.n122 B 0.010894f
C291 VDD1.n123 B 0.011535f
C292 VDD1.n124 B 0.02575f
C293 VDD1.n125 B 0.02575f
C294 VDD1.n126 B 0.011535f
C295 VDD1.n127 B 0.010894f
C296 VDD1.n128 B 0.020274f
C297 VDD1.n129 B 0.020274f
C298 VDD1.n130 B 0.010894f
C299 VDD1.n131 B 0.011535f
C300 VDD1.n132 B 0.02575f
C301 VDD1.n133 B 0.02575f
C302 VDD1.n134 B 0.011535f
C303 VDD1.n135 B 0.010894f
C304 VDD1.n136 B 0.020274f
C305 VDD1.n137 B 0.020274f
C306 VDD1.n138 B 0.010894f
C307 VDD1.n139 B 0.011535f
C308 VDD1.n140 B 0.02575f
C309 VDD1.n141 B 0.056953f
C310 VDD1.n142 B 0.011535f
C311 VDD1.n143 B 0.010894f
C312 VDD1.n144 B 0.04603f
C313 VDD1.n145 B 0.673822f
C314 VTAIL.n0 B 0.029337f
C315 VTAIL.n1 B 0.020382f
C316 VTAIL.n2 B 0.010953f
C317 VTAIL.n3 B 0.025888f
C318 VTAIL.n4 B 0.011597f
C319 VTAIL.n5 B 0.020382f
C320 VTAIL.n6 B 0.010953f
C321 VTAIL.n7 B 0.025888f
C322 VTAIL.n8 B 0.011597f
C323 VTAIL.n9 B 0.020382f
C324 VTAIL.n10 B 0.010953f
C325 VTAIL.n11 B 0.025888f
C326 VTAIL.n12 B 0.011275f
C327 VTAIL.n13 B 0.020382f
C328 VTAIL.n14 B 0.011597f
C329 VTAIL.n15 B 0.025888f
C330 VTAIL.n16 B 0.011597f
C331 VTAIL.n17 B 0.020382f
C332 VTAIL.n18 B 0.010953f
C333 VTAIL.n19 B 0.025888f
C334 VTAIL.n20 B 0.011597f
C335 VTAIL.n21 B 1.16697f
C336 VTAIL.n22 B 0.010953f
C337 VTAIL.t2 B 0.043891f
C338 VTAIL.n23 B 0.158928f
C339 VTAIL.n24 B 0.018301f
C340 VTAIL.n25 B 0.019416f
C341 VTAIL.n26 B 0.025888f
C342 VTAIL.n27 B 0.011597f
C343 VTAIL.n28 B 0.010953f
C344 VTAIL.n29 B 0.020382f
C345 VTAIL.n30 B 0.020382f
C346 VTAIL.n31 B 0.010953f
C347 VTAIL.n32 B 0.011597f
C348 VTAIL.n33 B 0.025888f
C349 VTAIL.n34 B 0.025888f
C350 VTAIL.n35 B 0.011597f
C351 VTAIL.n36 B 0.010953f
C352 VTAIL.n37 B 0.020382f
C353 VTAIL.n38 B 0.020382f
C354 VTAIL.n39 B 0.010953f
C355 VTAIL.n40 B 0.010953f
C356 VTAIL.n41 B 0.011597f
C357 VTAIL.n42 B 0.025888f
C358 VTAIL.n43 B 0.025888f
C359 VTAIL.n44 B 0.025888f
C360 VTAIL.n45 B 0.011275f
C361 VTAIL.n46 B 0.010953f
C362 VTAIL.n47 B 0.020382f
C363 VTAIL.n48 B 0.020382f
C364 VTAIL.n49 B 0.010953f
C365 VTAIL.n50 B 0.011597f
C366 VTAIL.n51 B 0.025888f
C367 VTAIL.n52 B 0.025888f
C368 VTAIL.n53 B 0.011597f
C369 VTAIL.n54 B 0.010953f
C370 VTAIL.n55 B 0.020382f
C371 VTAIL.n56 B 0.020382f
C372 VTAIL.n57 B 0.010953f
C373 VTAIL.n58 B 0.011597f
C374 VTAIL.n59 B 0.025888f
C375 VTAIL.n60 B 0.025888f
C376 VTAIL.n61 B 0.011597f
C377 VTAIL.n62 B 0.010953f
C378 VTAIL.n63 B 0.020382f
C379 VTAIL.n64 B 0.020382f
C380 VTAIL.n65 B 0.010953f
C381 VTAIL.n66 B 0.011597f
C382 VTAIL.n67 B 0.025888f
C383 VTAIL.n68 B 0.057259f
C384 VTAIL.n69 B 0.011597f
C385 VTAIL.n70 B 0.010953f
C386 VTAIL.n71 B 0.046278f
C387 VTAIL.n72 B 0.032138f
C388 VTAIL.n73 B 1.4423f
C389 VTAIL.n74 B 0.029337f
C390 VTAIL.n75 B 0.020382f
C391 VTAIL.n76 B 0.010953f
C392 VTAIL.n77 B 0.025888f
C393 VTAIL.n78 B 0.011597f
C394 VTAIL.n79 B 0.020382f
C395 VTAIL.n80 B 0.010953f
C396 VTAIL.n81 B 0.025888f
C397 VTAIL.n82 B 0.011597f
C398 VTAIL.n83 B 0.020382f
C399 VTAIL.n84 B 0.010953f
C400 VTAIL.n85 B 0.025888f
C401 VTAIL.n86 B 0.011275f
C402 VTAIL.n87 B 0.020382f
C403 VTAIL.n88 B 0.011275f
C404 VTAIL.n89 B 0.010953f
C405 VTAIL.n90 B 0.025888f
C406 VTAIL.n91 B 0.025888f
C407 VTAIL.n92 B 0.011597f
C408 VTAIL.n93 B 0.020382f
C409 VTAIL.n94 B 0.010953f
C410 VTAIL.n95 B 0.025888f
C411 VTAIL.n96 B 0.011597f
C412 VTAIL.n97 B 1.16697f
C413 VTAIL.n98 B 0.010953f
C414 VTAIL.t0 B 0.043891f
C415 VTAIL.n99 B 0.158928f
C416 VTAIL.n100 B 0.018301f
C417 VTAIL.n101 B 0.019416f
C418 VTAIL.n102 B 0.025888f
C419 VTAIL.n103 B 0.011597f
C420 VTAIL.n104 B 0.010953f
C421 VTAIL.n105 B 0.020382f
C422 VTAIL.n106 B 0.020382f
C423 VTAIL.n107 B 0.010953f
C424 VTAIL.n108 B 0.011597f
C425 VTAIL.n109 B 0.025888f
C426 VTAIL.n110 B 0.025888f
C427 VTAIL.n111 B 0.011597f
C428 VTAIL.n112 B 0.010953f
C429 VTAIL.n113 B 0.020382f
C430 VTAIL.n114 B 0.020382f
C431 VTAIL.n115 B 0.010953f
C432 VTAIL.n116 B 0.011597f
C433 VTAIL.n117 B 0.025888f
C434 VTAIL.n118 B 0.025888f
C435 VTAIL.n119 B 0.011597f
C436 VTAIL.n120 B 0.010953f
C437 VTAIL.n121 B 0.020382f
C438 VTAIL.n122 B 0.020382f
C439 VTAIL.n123 B 0.010953f
C440 VTAIL.n124 B 0.011597f
C441 VTAIL.n125 B 0.025888f
C442 VTAIL.n126 B 0.025888f
C443 VTAIL.n127 B 0.011597f
C444 VTAIL.n128 B 0.010953f
C445 VTAIL.n129 B 0.020382f
C446 VTAIL.n130 B 0.020382f
C447 VTAIL.n131 B 0.010953f
C448 VTAIL.n132 B 0.011597f
C449 VTAIL.n133 B 0.025888f
C450 VTAIL.n134 B 0.025888f
C451 VTAIL.n135 B 0.011597f
C452 VTAIL.n136 B 0.010953f
C453 VTAIL.n137 B 0.020382f
C454 VTAIL.n138 B 0.020382f
C455 VTAIL.n139 B 0.010953f
C456 VTAIL.n140 B 0.011597f
C457 VTAIL.n141 B 0.025888f
C458 VTAIL.n142 B 0.057259f
C459 VTAIL.n143 B 0.011597f
C460 VTAIL.n144 B 0.010953f
C461 VTAIL.n145 B 0.046278f
C462 VTAIL.n146 B 0.032138f
C463 VTAIL.n147 B 1.47712f
C464 VTAIL.n148 B 0.029337f
C465 VTAIL.n149 B 0.020382f
C466 VTAIL.n150 B 0.010953f
C467 VTAIL.n151 B 0.025888f
C468 VTAIL.n152 B 0.011597f
C469 VTAIL.n153 B 0.020382f
C470 VTAIL.n154 B 0.010953f
C471 VTAIL.n155 B 0.025888f
C472 VTAIL.n156 B 0.011597f
C473 VTAIL.n157 B 0.020382f
C474 VTAIL.n158 B 0.010953f
C475 VTAIL.n159 B 0.025888f
C476 VTAIL.n160 B 0.011275f
C477 VTAIL.n161 B 0.020382f
C478 VTAIL.n162 B 0.011275f
C479 VTAIL.n163 B 0.010953f
C480 VTAIL.n164 B 0.025888f
C481 VTAIL.n165 B 0.025888f
C482 VTAIL.n166 B 0.011597f
C483 VTAIL.n167 B 0.020382f
C484 VTAIL.n168 B 0.010953f
C485 VTAIL.n169 B 0.025888f
C486 VTAIL.n170 B 0.011597f
C487 VTAIL.n171 B 1.16697f
C488 VTAIL.n172 B 0.010953f
C489 VTAIL.t3 B 0.043891f
C490 VTAIL.n173 B 0.158928f
C491 VTAIL.n174 B 0.018301f
C492 VTAIL.n175 B 0.019416f
C493 VTAIL.n176 B 0.025888f
C494 VTAIL.n177 B 0.011597f
C495 VTAIL.n178 B 0.010953f
C496 VTAIL.n179 B 0.020382f
C497 VTAIL.n180 B 0.020382f
C498 VTAIL.n181 B 0.010953f
C499 VTAIL.n182 B 0.011597f
C500 VTAIL.n183 B 0.025888f
C501 VTAIL.n184 B 0.025888f
C502 VTAIL.n185 B 0.011597f
C503 VTAIL.n186 B 0.010953f
C504 VTAIL.n187 B 0.020382f
C505 VTAIL.n188 B 0.020382f
C506 VTAIL.n189 B 0.010953f
C507 VTAIL.n190 B 0.011597f
C508 VTAIL.n191 B 0.025888f
C509 VTAIL.n192 B 0.025888f
C510 VTAIL.n193 B 0.011597f
C511 VTAIL.n194 B 0.010953f
C512 VTAIL.n195 B 0.020382f
C513 VTAIL.n196 B 0.020382f
C514 VTAIL.n197 B 0.010953f
C515 VTAIL.n198 B 0.011597f
C516 VTAIL.n199 B 0.025888f
C517 VTAIL.n200 B 0.025888f
C518 VTAIL.n201 B 0.011597f
C519 VTAIL.n202 B 0.010953f
C520 VTAIL.n203 B 0.020382f
C521 VTAIL.n204 B 0.020382f
C522 VTAIL.n205 B 0.010953f
C523 VTAIL.n206 B 0.011597f
C524 VTAIL.n207 B 0.025888f
C525 VTAIL.n208 B 0.025888f
C526 VTAIL.n209 B 0.011597f
C527 VTAIL.n210 B 0.010953f
C528 VTAIL.n211 B 0.020382f
C529 VTAIL.n212 B 0.020382f
C530 VTAIL.n213 B 0.010953f
C531 VTAIL.n214 B 0.011597f
C532 VTAIL.n215 B 0.025888f
C533 VTAIL.n216 B 0.057259f
C534 VTAIL.n217 B 0.011597f
C535 VTAIL.n218 B 0.010953f
C536 VTAIL.n219 B 0.046278f
C537 VTAIL.n220 B 0.032138f
C538 VTAIL.n221 B 1.32256f
C539 VTAIL.n222 B 0.029337f
C540 VTAIL.n223 B 0.020382f
C541 VTAIL.n224 B 0.010953f
C542 VTAIL.n225 B 0.025888f
C543 VTAIL.n226 B 0.011597f
C544 VTAIL.n227 B 0.020382f
C545 VTAIL.n228 B 0.010953f
C546 VTAIL.n229 B 0.025888f
C547 VTAIL.n230 B 0.011597f
C548 VTAIL.n231 B 0.020382f
C549 VTAIL.n232 B 0.010953f
C550 VTAIL.n233 B 0.025888f
C551 VTAIL.n234 B 0.011275f
C552 VTAIL.n235 B 0.020382f
C553 VTAIL.n236 B 0.011597f
C554 VTAIL.n237 B 0.025888f
C555 VTAIL.n238 B 0.011597f
C556 VTAIL.n239 B 0.020382f
C557 VTAIL.n240 B 0.010953f
C558 VTAIL.n241 B 0.025888f
C559 VTAIL.n242 B 0.011597f
C560 VTAIL.n243 B 1.16697f
C561 VTAIL.n244 B 0.010953f
C562 VTAIL.t1 B 0.043891f
C563 VTAIL.n245 B 0.158928f
C564 VTAIL.n246 B 0.018301f
C565 VTAIL.n247 B 0.019416f
C566 VTAIL.n248 B 0.025888f
C567 VTAIL.n249 B 0.011597f
C568 VTAIL.n250 B 0.010953f
C569 VTAIL.n251 B 0.020382f
C570 VTAIL.n252 B 0.020382f
C571 VTAIL.n253 B 0.010953f
C572 VTAIL.n254 B 0.011597f
C573 VTAIL.n255 B 0.025888f
C574 VTAIL.n256 B 0.025888f
C575 VTAIL.n257 B 0.011597f
C576 VTAIL.n258 B 0.010953f
C577 VTAIL.n259 B 0.020382f
C578 VTAIL.n260 B 0.020382f
C579 VTAIL.n261 B 0.010953f
C580 VTAIL.n262 B 0.010953f
C581 VTAIL.n263 B 0.011597f
C582 VTAIL.n264 B 0.025888f
C583 VTAIL.n265 B 0.025888f
C584 VTAIL.n266 B 0.025888f
C585 VTAIL.n267 B 0.011275f
C586 VTAIL.n268 B 0.010953f
C587 VTAIL.n269 B 0.020382f
C588 VTAIL.n270 B 0.020382f
C589 VTAIL.n271 B 0.010953f
C590 VTAIL.n272 B 0.011597f
C591 VTAIL.n273 B 0.025888f
C592 VTAIL.n274 B 0.025888f
C593 VTAIL.n275 B 0.011597f
C594 VTAIL.n276 B 0.010953f
C595 VTAIL.n277 B 0.020382f
C596 VTAIL.n278 B 0.020382f
C597 VTAIL.n279 B 0.010953f
C598 VTAIL.n280 B 0.011597f
C599 VTAIL.n281 B 0.025888f
C600 VTAIL.n282 B 0.025888f
C601 VTAIL.n283 B 0.011597f
C602 VTAIL.n284 B 0.010953f
C603 VTAIL.n285 B 0.020382f
C604 VTAIL.n286 B 0.020382f
C605 VTAIL.n287 B 0.010953f
C606 VTAIL.n288 B 0.011597f
C607 VTAIL.n289 B 0.025888f
C608 VTAIL.n290 B 0.057259f
C609 VTAIL.n291 B 0.011597f
C610 VTAIL.n292 B 0.010953f
C611 VTAIL.n293 B 0.046278f
C612 VTAIL.n294 B 0.032138f
C613 VTAIL.n295 B 1.24924f
C614 VP.t1 B 3.70005f
C615 VP.t0 B 3.20148f
C616 VP.n0 B 4.52676f
.ends

