* NGSPICE file created from diff_pair_sample_1281.ext - technology: sky130A

.subckt diff_pair_sample_1281 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X1 VTAIL.t14 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X2 VDD1.t7 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X3 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X4 VDD2.t7 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=4.4616 ps=23.66 w=11.44 l=3.81
X5 VTAIL.t12 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=1.8876 ps=11.77 w=11.44 l=3.81
X6 VDD1.t5 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=4.4616 ps=23.66 w=11.44 l=3.81
X7 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=0 ps=0 w=11.44 l=3.81
X8 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=0 ps=0 w=11.44 l=3.81
X9 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=0 ps=0 w=11.44 l=3.81
X10 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=1.8876 ps=11.77 w=11.44 l=3.81
X11 VTAIL.t7 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=1.8876 ps=11.77 w=11.44 l=3.81
X12 VDD2.t1 VN.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=4.4616 ps=23.66 w=11.44 l=3.81
X13 VDD2.t0 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X14 VTAIL.t9 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=1.8876 ps=11.77 w=11.44 l=3.81
X15 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=4.4616 ps=23.66 w=11.44 l=3.81
X16 VDD2.t2 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X17 VDD1.t1 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X18 VTAIL.t1 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8876 pd=11.77 as=1.8876 ps=11.77 w=11.44 l=3.81
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4616 pd=23.66 as=0 ps=0 w=11.44 l=3.81
R0 VN.n71 VN.n37 161.3
R1 VN.n70 VN.n69 161.3
R2 VN.n68 VN.n38 161.3
R3 VN.n67 VN.n66 161.3
R4 VN.n65 VN.n39 161.3
R5 VN.n64 VN.n63 161.3
R6 VN.n62 VN.n40 161.3
R7 VN.n61 VN.n60 161.3
R8 VN.n58 VN.n41 161.3
R9 VN.n57 VN.n56 161.3
R10 VN.n55 VN.n42 161.3
R11 VN.n54 VN.n53 161.3
R12 VN.n52 VN.n43 161.3
R13 VN.n51 VN.n50 161.3
R14 VN.n49 VN.n44 161.3
R15 VN.n48 VN.n47 161.3
R16 VN.n34 VN.n0 161.3
R17 VN.n33 VN.n32 161.3
R18 VN.n31 VN.n1 161.3
R19 VN.n30 VN.n29 161.3
R20 VN.n28 VN.n2 161.3
R21 VN.n27 VN.n26 161.3
R22 VN.n25 VN.n3 161.3
R23 VN.n24 VN.n23 161.3
R24 VN.n21 VN.n4 161.3
R25 VN.n20 VN.n19 161.3
R26 VN.n18 VN.n5 161.3
R27 VN.n17 VN.n16 161.3
R28 VN.n15 VN.n6 161.3
R29 VN.n14 VN.n13 161.3
R30 VN.n12 VN.n7 161.3
R31 VN.n11 VN.n10 161.3
R32 VN.n8 VN.t6 104.632
R33 VN.n45 VN.t4 104.632
R34 VN.n9 VN.t7 72.3638
R35 VN.n22 VN.t1 72.3638
R36 VN.n35 VN.t2 72.3638
R37 VN.n46 VN.t0 72.3638
R38 VN.n59 VN.t5 72.3638
R39 VN.n72 VN.t3 72.3638
R40 VN.n36 VN.n35 59.7554
R41 VN.n73 VN.n72 59.7554
R42 VN.n9 VN.n8 59.5587
R43 VN.n46 VN.n45 59.5587
R44 VN.n16 VN.n15 56.5617
R45 VN.n53 VN.n52 56.5617
R46 VN VN.n73 56.4059
R47 VN.n29 VN.n28 51.2335
R48 VN.n66 VN.n65 51.2335
R49 VN.n29 VN.n1 29.9206
R50 VN.n66 VN.n38 29.9206
R51 VN.n10 VN.n7 24.5923
R52 VN.n14 VN.n7 24.5923
R53 VN.n15 VN.n14 24.5923
R54 VN.n16 VN.n5 24.5923
R55 VN.n20 VN.n5 24.5923
R56 VN.n21 VN.n20 24.5923
R57 VN.n23 VN.n3 24.5923
R58 VN.n27 VN.n3 24.5923
R59 VN.n28 VN.n27 24.5923
R60 VN.n33 VN.n1 24.5923
R61 VN.n34 VN.n33 24.5923
R62 VN.n52 VN.n51 24.5923
R63 VN.n51 VN.n44 24.5923
R64 VN.n47 VN.n44 24.5923
R65 VN.n65 VN.n64 24.5923
R66 VN.n64 VN.n40 24.5923
R67 VN.n60 VN.n40 24.5923
R68 VN.n58 VN.n57 24.5923
R69 VN.n57 VN.n42 24.5923
R70 VN.n53 VN.n42 24.5923
R71 VN.n71 VN.n70 24.5923
R72 VN.n70 VN.n38 24.5923
R73 VN.n35 VN.n34 22.625
R74 VN.n72 VN.n71 22.625
R75 VN.n10 VN.n9 15.7393
R76 VN.n22 VN.n21 15.7393
R77 VN.n47 VN.n46 15.7393
R78 VN.n59 VN.n58 15.7393
R79 VN.n23 VN.n22 8.85356
R80 VN.n60 VN.n59 8.85356
R81 VN.n48 VN.n45 2.58852
R82 VN.n11 VN.n8 2.58852
R83 VN.n73 VN.n37 0.417304
R84 VN.n36 VN.n0 0.417304
R85 VN VN.n36 0.394524
R86 VN.n69 VN.n37 0.189894
R87 VN.n69 VN.n68 0.189894
R88 VN.n68 VN.n67 0.189894
R89 VN.n67 VN.n39 0.189894
R90 VN.n63 VN.n39 0.189894
R91 VN.n63 VN.n62 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n41 0.189894
R94 VN.n56 VN.n41 0.189894
R95 VN.n56 VN.n55 0.189894
R96 VN.n55 VN.n54 0.189894
R97 VN.n54 VN.n43 0.189894
R98 VN.n50 VN.n43 0.189894
R99 VN.n50 VN.n49 0.189894
R100 VN.n49 VN.n48 0.189894
R101 VN.n12 VN.n11 0.189894
R102 VN.n13 VN.n12 0.189894
R103 VN.n13 VN.n6 0.189894
R104 VN.n17 VN.n6 0.189894
R105 VN.n18 VN.n17 0.189894
R106 VN.n19 VN.n18 0.189894
R107 VN.n19 VN.n4 0.189894
R108 VN.n24 VN.n4 0.189894
R109 VN.n25 VN.n24 0.189894
R110 VN.n26 VN.n25 0.189894
R111 VN.n26 VN.n2 0.189894
R112 VN.n30 VN.n2 0.189894
R113 VN.n31 VN.n30 0.189894
R114 VN.n32 VN.n31 0.189894
R115 VN.n32 VN.n0 0.189894
R116 VDD2.n2 VDD2.n1 64.5946
R117 VDD2.n2 VDD2.n0 64.5946
R118 VDD2 VDD2.n5 64.5918
R119 VDD2.n4 VDD2.n3 62.8657
R120 VDD2.n4 VDD2.n2 49.6377
R121 VDD2 VDD2.n4 1.84317
R122 VDD2.n5 VDD2.t5 1.73127
R123 VDD2.n5 VDD2.t1 1.73127
R124 VDD2.n3 VDD2.t6 1.73127
R125 VDD2.n3 VDD2.t0 1.73127
R126 VDD2.n1 VDD2.t4 1.73127
R127 VDD2.n1 VDD2.t7 1.73127
R128 VDD2.n0 VDD2.t3 1.73127
R129 VDD2.n0 VDD2.t2 1.73127
R130 VTAIL.n498 VTAIL.n442 289.615
R131 VTAIL.n58 VTAIL.n2 289.615
R132 VTAIL.n120 VTAIL.n64 289.615
R133 VTAIL.n184 VTAIL.n128 289.615
R134 VTAIL.n436 VTAIL.n380 289.615
R135 VTAIL.n372 VTAIL.n316 289.615
R136 VTAIL.n310 VTAIL.n254 289.615
R137 VTAIL.n246 VTAIL.n190 289.615
R138 VTAIL.n463 VTAIL.n462 185
R139 VTAIL.n465 VTAIL.n464 185
R140 VTAIL.n458 VTAIL.n457 185
R141 VTAIL.n471 VTAIL.n470 185
R142 VTAIL.n473 VTAIL.n472 185
R143 VTAIL.n454 VTAIL.n453 185
R144 VTAIL.n480 VTAIL.n479 185
R145 VTAIL.n481 VTAIL.n452 185
R146 VTAIL.n483 VTAIL.n482 185
R147 VTAIL.n450 VTAIL.n449 185
R148 VTAIL.n489 VTAIL.n488 185
R149 VTAIL.n491 VTAIL.n490 185
R150 VTAIL.n446 VTAIL.n445 185
R151 VTAIL.n497 VTAIL.n496 185
R152 VTAIL.n499 VTAIL.n498 185
R153 VTAIL.n23 VTAIL.n22 185
R154 VTAIL.n25 VTAIL.n24 185
R155 VTAIL.n18 VTAIL.n17 185
R156 VTAIL.n31 VTAIL.n30 185
R157 VTAIL.n33 VTAIL.n32 185
R158 VTAIL.n14 VTAIL.n13 185
R159 VTAIL.n40 VTAIL.n39 185
R160 VTAIL.n41 VTAIL.n12 185
R161 VTAIL.n43 VTAIL.n42 185
R162 VTAIL.n10 VTAIL.n9 185
R163 VTAIL.n49 VTAIL.n48 185
R164 VTAIL.n51 VTAIL.n50 185
R165 VTAIL.n6 VTAIL.n5 185
R166 VTAIL.n57 VTAIL.n56 185
R167 VTAIL.n59 VTAIL.n58 185
R168 VTAIL.n85 VTAIL.n84 185
R169 VTAIL.n87 VTAIL.n86 185
R170 VTAIL.n80 VTAIL.n79 185
R171 VTAIL.n93 VTAIL.n92 185
R172 VTAIL.n95 VTAIL.n94 185
R173 VTAIL.n76 VTAIL.n75 185
R174 VTAIL.n102 VTAIL.n101 185
R175 VTAIL.n103 VTAIL.n74 185
R176 VTAIL.n105 VTAIL.n104 185
R177 VTAIL.n72 VTAIL.n71 185
R178 VTAIL.n111 VTAIL.n110 185
R179 VTAIL.n113 VTAIL.n112 185
R180 VTAIL.n68 VTAIL.n67 185
R181 VTAIL.n119 VTAIL.n118 185
R182 VTAIL.n121 VTAIL.n120 185
R183 VTAIL.n149 VTAIL.n148 185
R184 VTAIL.n151 VTAIL.n150 185
R185 VTAIL.n144 VTAIL.n143 185
R186 VTAIL.n157 VTAIL.n156 185
R187 VTAIL.n159 VTAIL.n158 185
R188 VTAIL.n140 VTAIL.n139 185
R189 VTAIL.n166 VTAIL.n165 185
R190 VTAIL.n167 VTAIL.n138 185
R191 VTAIL.n169 VTAIL.n168 185
R192 VTAIL.n136 VTAIL.n135 185
R193 VTAIL.n175 VTAIL.n174 185
R194 VTAIL.n177 VTAIL.n176 185
R195 VTAIL.n132 VTAIL.n131 185
R196 VTAIL.n183 VTAIL.n182 185
R197 VTAIL.n185 VTAIL.n184 185
R198 VTAIL.n437 VTAIL.n436 185
R199 VTAIL.n435 VTAIL.n434 185
R200 VTAIL.n384 VTAIL.n383 185
R201 VTAIL.n429 VTAIL.n428 185
R202 VTAIL.n427 VTAIL.n426 185
R203 VTAIL.n388 VTAIL.n387 185
R204 VTAIL.n392 VTAIL.n390 185
R205 VTAIL.n421 VTAIL.n420 185
R206 VTAIL.n419 VTAIL.n418 185
R207 VTAIL.n394 VTAIL.n393 185
R208 VTAIL.n413 VTAIL.n412 185
R209 VTAIL.n411 VTAIL.n410 185
R210 VTAIL.n398 VTAIL.n397 185
R211 VTAIL.n405 VTAIL.n404 185
R212 VTAIL.n403 VTAIL.n402 185
R213 VTAIL.n373 VTAIL.n372 185
R214 VTAIL.n371 VTAIL.n370 185
R215 VTAIL.n320 VTAIL.n319 185
R216 VTAIL.n365 VTAIL.n364 185
R217 VTAIL.n363 VTAIL.n362 185
R218 VTAIL.n324 VTAIL.n323 185
R219 VTAIL.n328 VTAIL.n326 185
R220 VTAIL.n357 VTAIL.n356 185
R221 VTAIL.n355 VTAIL.n354 185
R222 VTAIL.n330 VTAIL.n329 185
R223 VTAIL.n349 VTAIL.n348 185
R224 VTAIL.n347 VTAIL.n346 185
R225 VTAIL.n334 VTAIL.n333 185
R226 VTAIL.n341 VTAIL.n340 185
R227 VTAIL.n339 VTAIL.n338 185
R228 VTAIL.n311 VTAIL.n310 185
R229 VTAIL.n309 VTAIL.n308 185
R230 VTAIL.n258 VTAIL.n257 185
R231 VTAIL.n303 VTAIL.n302 185
R232 VTAIL.n301 VTAIL.n300 185
R233 VTAIL.n262 VTAIL.n261 185
R234 VTAIL.n266 VTAIL.n264 185
R235 VTAIL.n295 VTAIL.n294 185
R236 VTAIL.n293 VTAIL.n292 185
R237 VTAIL.n268 VTAIL.n267 185
R238 VTAIL.n287 VTAIL.n286 185
R239 VTAIL.n285 VTAIL.n284 185
R240 VTAIL.n272 VTAIL.n271 185
R241 VTAIL.n279 VTAIL.n278 185
R242 VTAIL.n277 VTAIL.n276 185
R243 VTAIL.n247 VTAIL.n246 185
R244 VTAIL.n245 VTAIL.n244 185
R245 VTAIL.n194 VTAIL.n193 185
R246 VTAIL.n239 VTAIL.n238 185
R247 VTAIL.n237 VTAIL.n236 185
R248 VTAIL.n198 VTAIL.n197 185
R249 VTAIL.n202 VTAIL.n200 185
R250 VTAIL.n231 VTAIL.n230 185
R251 VTAIL.n229 VTAIL.n228 185
R252 VTAIL.n204 VTAIL.n203 185
R253 VTAIL.n223 VTAIL.n222 185
R254 VTAIL.n221 VTAIL.n220 185
R255 VTAIL.n208 VTAIL.n207 185
R256 VTAIL.n215 VTAIL.n214 185
R257 VTAIL.n213 VTAIL.n212 185
R258 VTAIL.n461 VTAIL.t13 149.524
R259 VTAIL.n21 VTAIL.t9 149.524
R260 VTAIL.n83 VTAIL.t2 149.524
R261 VTAIL.n147 VTAIL.t7 149.524
R262 VTAIL.n401 VTAIL.t3 149.524
R263 VTAIL.n337 VTAIL.t0 149.524
R264 VTAIL.n275 VTAIL.t11 149.524
R265 VTAIL.n211 VTAIL.t12 149.524
R266 VTAIL.n464 VTAIL.n463 104.615
R267 VTAIL.n464 VTAIL.n457 104.615
R268 VTAIL.n471 VTAIL.n457 104.615
R269 VTAIL.n472 VTAIL.n471 104.615
R270 VTAIL.n472 VTAIL.n453 104.615
R271 VTAIL.n480 VTAIL.n453 104.615
R272 VTAIL.n481 VTAIL.n480 104.615
R273 VTAIL.n482 VTAIL.n481 104.615
R274 VTAIL.n482 VTAIL.n449 104.615
R275 VTAIL.n489 VTAIL.n449 104.615
R276 VTAIL.n490 VTAIL.n489 104.615
R277 VTAIL.n490 VTAIL.n445 104.615
R278 VTAIL.n497 VTAIL.n445 104.615
R279 VTAIL.n498 VTAIL.n497 104.615
R280 VTAIL.n24 VTAIL.n23 104.615
R281 VTAIL.n24 VTAIL.n17 104.615
R282 VTAIL.n31 VTAIL.n17 104.615
R283 VTAIL.n32 VTAIL.n31 104.615
R284 VTAIL.n32 VTAIL.n13 104.615
R285 VTAIL.n40 VTAIL.n13 104.615
R286 VTAIL.n41 VTAIL.n40 104.615
R287 VTAIL.n42 VTAIL.n41 104.615
R288 VTAIL.n42 VTAIL.n9 104.615
R289 VTAIL.n49 VTAIL.n9 104.615
R290 VTAIL.n50 VTAIL.n49 104.615
R291 VTAIL.n50 VTAIL.n5 104.615
R292 VTAIL.n57 VTAIL.n5 104.615
R293 VTAIL.n58 VTAIL.n57 104.615
R294 VTAIL.n86 VTAIL.n85 104.615
R295 VTAIL.n86 VTAIL.n79 104.615
R296 VTAIL.n93 VTAIL.n79 104.615
R297 VTAIL.n94 VTAIL.n93 104.615
R298 VTAIL.n94 VTAIL.n75 104.615
R299 VTAIL.n102 VTAIL.n75 104.615
R300 VTAIL.n103 VTAIL.n102 104.615
R301 VTAIL.n104 VTAIL.n103 104.615
R302 VTAIL.n104 VTAIL.n71 104.615
R303 VTAIL.n111 VTAIL.n71 104.615
R304 VTAIL.n112 VTAIL.n111 104.615
R305 VTAIL.n112 VTAIL.n67 104.615
R306 VTAIL.n119 VTAIL.n67 104.615
R307 VTAIL.n120 VTAIL.n119 104.615
R308 VTAIL.n150 VTAIL.n149 104.615
R309 VTAIL.n150 VTAIL.n143 104.615
R310 VTAIL.n157 VTAIL.n143 104.615
R311 VTAIL.n158 VTAIL.n157 104.615
R312 VTAIL.n158 VTAIL.n139 104.615
R313 VTAIL.n166 VTAIL.n139 104.615
R314 VTAIL.n167 VTAIL.n166 104.615
R315 VTAIL.n168 VTAIL.n167 104.615
R316 VTAIL.n168 VTAIL.n135 104.615
R317 VTAIL.n175 VTAIL.n135 104.615
R318 VTAIL.n176 VTAIL.n175 104.615
R319 VTAIL.n176 VTAIL.n131 104.615
R320 VTAIL.n183 VTAIL.n131 104.615
R321 VTAIL.n184 VTAIL.n183 104.615
R322 VTAIL.n436 VTAIL.n435 104.615
R323 VTAIL.n435 VTAIL.n383 104.615
R324 VTAIL.n428 VTAIL.n383 104.615
R325 VTAIL.n428 VTAIL.n427 104.615
R326 VTAIL.n427 VTAIL.n387 104.615
R327 VTAIL.n392 VTAIL.n387 104.615
R328 VTAIL.n420 VTAIL.n392 104.615
R329 VTAIL.n420 VTAIL.n419 104.615
R330 VTAIL.n419 VTAIL.n393 104.615
R331 VTAIL.n412 VTAIL.n393 104.615
R332 VTAIL.n412 VTAIL.n411 104.615
R333 VTAIL.n411 VTAIL.n397 104.615
R334 VTAIL.n404 VTAIL.n397 104.615
R335 VTAIL.n404 VTAIL.n403 104.615
R336 VTAIL.n372 VTAIL.n371 104.615
R337 VTAIL.n371 VTAIL.n319 104.615
R338 VTAIL.n364 VTAIL.n319 104.615
R339 VTAIL.n364 VTAIL.n363 104.615
R340 VTAIL.n363 VTAIL.n323 104.615
R341 VTAIL.n328 VTAIL.n323 104.615
R342 VTAIL.n356 VTAIL.n328 104.615
R343 VTAIL.n356 VTAIL.n355 104.615
R344 VTAIL.n355 VTAIL.n329 104.615
R345 VTAIL.n348 VTAIL.n329 104.615
R346 VTAIL.n348 VTAIL.n347 104.615
R347 VTAIL.n347 VTAIL.n333 104.615
R348 VTAIL.n340 VTAIL.n333 104.615
R349 VTAIL.n340 VTAIL.n339 104.615
R350 VTAIL.n310 VTAIL.n309 104.615
R351 VTAIL.n309 VTAIL.n257 104.615
R352 VTAIL.n302 VTAIL.n257 104.615
R353 VTAIL.n302 VTAIL.n301 104.615
R354 VTAIL.n301 VTAIL.n261 104.615
R355 VTAIL.n266 VTAIL.n261 104.615
R356 VTAIL.n294 VTAIL.n266 104.615
R357 VTAIL.n294 VTAIL.n293 104.615
R358 VTAIL.n293 VTAIL.n267 104.615
R359 VTAIL.n286 VTAIL.n267 104.615
R360 VTAIL.n286 VTAIL.n285 104.615
R361 VTAIL.n285 VTAIL.n271 104.615
R362 VTAIL.n278 VTAIL.n271 104.615
R363 VTAIL.n278 VTAIL.n277 104.615
R364 VTAIL.n246 VTAIL.n245 104.615
R365 VTAIL.n245 VTAIL.n193 104.615
R366 VTAIL.n238 VTAIL.n193 104.615
R367 VTAIL.n238 VTAIL.n237 104.615
R368 VTAIL.n237 VTAIL.n197 104.615
R369 VTAIL.n202 VTAIL.n197 104.615
R370 VTAIL.n230 VTAIL.n202 104.615
R371 VTAIL.n230 VTAIL.n229 104.615
R372 VTAIL.n229 VTAIL.n203 104.615
R373 VTAIL.n222 VTAIL.n203 104.615
R374 VTAIL.n222 VTAIL.n221 104.615
R375 VTAIL.n221 VTAIL.n207 104.615
R376 VTAIL.n214 VTAIL.n207 104.615
R377 VTAIL.n214 VTAIL.n213 104.615
R378 VTAIL.n463 VTAIL.t13 52.3082
R379 VTAIL.n23 VTAIL.t9 52.3082
R380 VTAIL.n85 VTAIL.t2 52.3082
R381 VTAIL.n149 VTAIL.t7 52.3082
R382 VTAIL.n403 VTAIL.t3 52.3082
R383 VTAIL.n339 VTAIL.t0 52.3082
R384 VTAIL.n277 VTAIL.t11 52.3082
R385 VTAIL.n213 VTAIL.t12 52.3082
R386 VTAIL.n379 VTAIL.n378 46.1869
R387 VTAIL.n253 VTAIL.n252 46.1869
R388 VTAIL.n1 VTAIL.n0 46.1867
R389 VTAIL.n127 VTAIL.n126 46.1867
R390 VTAIL.n503 VTAIL.n502 32.9611
R391 VTAIL.n63 VTAIL.n62 32.9611
R392 VTAIL.n125 VTAIL.n124 32.9611
R393 VTAIL.n189 VTAIL.n188 32.9611
R394 VTAIL.n441 VTAIL.n440 32.9611
R395 VTAIL.n377 VTAIL.n376 32.9611
R396 VTAIL.n315 VTAIL.n314 32.9611
R397 VTAIL.n251 VTAIL.n250 32.9611
R398 VTAIL.n503 VTAIL.n441 25.7979
R399 VTAIL.n251 VTAIL.n189 25.7979
R400 VTAIL.n483 VTAIL.n450 13.1884
R401 VTAIL.n43 VTAIL.n10 13.1884
R402 VTAIL.n105 VTAIL.n72 13.1884
R403 VTAIL.n169 VTAIL.n136 13.1884
R404 VTAIL.n390 VTAIL.n388 13.1884
R405 VTAIL.n326 VTAIL.n324 13.1884
R406 VTAIL.n264 VTAIL.n262 13.1884
R407 VTAIL.n200 VTAIL.n198 13.1884
R408 VTAIL.n484 VTAIL.n452 12.8005
R409 VTAIL.n488 VTAIL.n487 12.8005
R410 VTAIL.n44 VTAIL.n12 12.8005
R411 VTAIL.n48 VTAIL.n47 12.8005
R412 VTAIL.n106 VTAIL.n74 12.8005
R413 VTAIL.n110 VTAIL.n109 12.8005
R414 VTAIL.n170 VTAIL.n138 12.8005
R415 VTAIL.n174 VTAIL.n173 12.8005
R416 VTAIL.n426 VTAIL.n425 12.8005
R417 VTAIL.n422 VTAIL.n421 12.8005
R418 VTAIL.n362 VTAIL.n361 12.8005
R419 VTAIL.n358 VTAIL.n357 12.8005
R420 VTAIL.n300 VTAIL.n299 12.8005
R421 VTAIL.n296 VTAIL.n295 12.8005
R422 VTAIL.n236 VTAIL.n235 12.8005
R423 VTAIL.n232 VTAIL.n231 12.8005
R424 VTAIL.n479 VTAIL.n478 12.0247
R425 VTAIL.n491 VTAIL.n448 12.0247
R426 VTAIL.n39 VTAIL.n38 12.0247
R427 VTAIL.n51 VTAIL.n8 12.0247
R428 VTAIL.n101 VTAIL.n100 12.0247
R429 VTAIL.n113 VTAIL.n70 12.0247
R430 VTAIL.n165 VTAIL.n164 12.0247
R431 VTAIL.n177 VTAIL.n134 12.0247
R432 VTAIL.n429 VTAIL.n386 12.0247
R433 VTAIL.n418 VTAIL.n391 12.0247
R434 VTAIL.n365 VTAIL.n322 12.0247
R435 VTAIL.n354 VTAIL.n327 12.0247
R436 VTAIL.n303 VTAIL.n260 12.0247
R437 VTAIL.n292 VTAIL.n265 12.0247
R438 VTAIL.n239 VTAIL.n196 12.0247
R439 VTAIL.n228 VTAIL.n201 12.0247
R440 VTAIL.n477 VTAIL.n454 11.249
R441 VTAIL.n492 VTAIL.n446 11.249
R442 VTAIL.n37 VTAIL.n14 11.249
R443 VTAIL.n52 VTAIL.n6 11.249
R444 VTAIL.n99 VTAIL.n76 11.249
R445 VTAIL.n114 VTAIL.n68 11.249
R446 VTAIL.n163 VTAIL.n140 11.249
R447 VTAIL.n178 VTAIL.n132 11.249
R448 VTAIL.n430 VTAIL.n384 11.249
R449 VTAIL.n417 VTAIL.n394 11.249
R450 VTAIL.n366 VTAIL.n320 11.249
R451 VTAIL.n353 VTAIL.n330 11.249
R452 VTAIL.n304 VTAIL.n258 11.249
R453 VTAIL.n291 VTAIL.n268 11.249
R454 VTAIL.n240 VTAIL.n194 11.249
R455 VTAIL.n227 VTAIL.n204 11.249
R456 VTAIL.n474 VTAIL.n473 10.4732
R457 VTAIL.n496 VTAIL.n495 10.4732
R458 VTAIL.n34 VTAIL.n33 10.4732
R459 VTAIL.n56 VTAIL.n55 10.4732
R460 VTAIL.n96 VTAIL.n95 10.4732
R461 VTAIL.n118 VTAIL.n117 10.4732
R462 VTAIL.n160 VTAIL.n159 10.4732
R463 VTAIL.n182 VTAIL.n181 10.4732
R464 VTAIL.n434 VTAIL.n433 10.4732
R465 VTAIL.n414 VTAIL.n413 10.4732
R466 VTAIL.n370 VTAIL.n369 10.4732
R467 VTAIL.n350 VTAIL.n349 10.4732
R468 VTAIL.n308 VTAIL.n307 10.4732
R469 VTAIL.n288 VTAIL.n287 10.4732
R470 VTAIL.n244 VTAIL.n243 10.4732
R471 VTAIL.n224 VTAIL.n223 10.4732
R472 VTAIL.n462 VTAIL.n461 10.2747
R473 VTAIL.n22 VTAIL.n21 10.2747
R474 VTAIL.n84 VTAIL.n83 10.2747
R475 VTAIL.n148 VTAIL.n147 10.2747
R476 VTAIL.n402 VTAIL.n401 10.2747
R477 VTAIL.n338 VTAIL.n337 10.2747
R478 VTAIL.n276 VTAIL.n275 10.2747
R479 VTAIL.n212 VTAIL.n211 10.2747
R480 VTAIL.n470 VTAIL.n456 9.69747
R481 VTAIL.n499 VTAIL.n444 9.69747
R482 VTAIL.n30 VTAIL.n16 9.69747
R483 VTAIL.n59 VTAIL.n4 9.69747
R484 VTAIL.n92 VTAIL.n78 9.69747
R485 VTAIL.n121 VTAIL.n66 9.69747
R486 VTAIL.n156 VTAIL.n142 9.69747
R487 VTAIL.n185 VTAIL.n130 9.69747
R488 VTAIL.n437 VTAIL.n382 9.69747
R489 VTAIL.n410 VTAIL.n396 9.69747
R490 VTAIL.n373 VTAIL.n318 9.69747
R491 VTAIL.n346 VTAIL.n332 9.69747
R492 VTAIL.n311 VTAIL.n256 9.69747
R493 VTAIL.n284 VTAIL.n270 9.69747
R494 VTAIL.n247 VTAIL.n192 9.69747
R495 VTAIL.n220 VTAIL.n206 9.69747
R496 VTAIL.n502 VTAIL.n501 9.45567
R497 VTAIL.n62 VTAIL.n61 9.45567
R498 VTAIL.n124 VTAIL.n123 9.45567
R499 VTAIL.n188 VTAIL.n187 9.45567
R500 VTAIL.n440 VTAIL.n439 9.45567
R501 VTAIL.n376 VTAIL.n375 9.45567
R502 VTAIL.n314 VTAIL.n313 9.45567
R503 VTAIL.n250 VTAIL.n249 9.45567
R504 VTAIL.n501 VTAIL.n500 9.3005
R505 VTAIL.n444 VTAIL.n443 9.3005
R506 VTAIL.n495 VTAIL.n494 9.3005
R507 VTAIL.n493 VTAIL.n492 9.3005
R508 VTAIL.n448 VTAIL.n447 9.3005
R509 VTAIL.n487 VTAIL.n486 9.3005
R510 VTAIL.n460 VTAIL.n459 9.3005
R511 VTAIL.n467 VTAIL.n466 9.3005
R512 VTAIL.n469 VTAIL.n468 9.3005
R513 VTAIL.n456 VTAIL.n455 9.3005
R514 VTAIL.n475 VTAIL.n474 9.3005
R515 VTAIL.n477 VTAIL.n476 9.3005
R516 VTAIL.n478 VTAIL.n451 9.3005
R517 VTAIL.n485 VTAIL.n484 9.3005
R518 VTAIL.n61 VTAIL.n60 9.3005
R519 VTAIL.n4 VTAIL.n3 9.3005
R520 VTAIL.n55 VTAIL.n54 9.3005
R521 VTAIL.n53 VTAIL.n52 9.3005
R522 VTAIL.n8 VTAIL.n7 9.3005
R523 VTAIL.n47 VTAIL.n46 9.3005
R524 VTAIL.n20 VTAIL.n19 9.3005
R525 VTAIL.n27 VTAIL.n26 9.3005
R526 VTAIL.n29 VTAIL.n28 9.3005
R527 VTAIL.n16 VTAIL.n15 9.3005
R528 VTAIL.n35 VTAIL.n34 9.3005
R529 VTAIL.n37 VTAIL.n36 9.3005
R530 VTAIL.n38 VTAIL.n11 9.3005
R531 VTAIL.n45 VTAIL.n44 9.3005
R532 VTAIL.n123 VTAIL.n122 9.3005
R533 VTAIL.n66 VTAIL.n65 9.3005
R534 VTAIL.n117 VTAIL.n116 9.3005
R535 VTAIL.n115 VTAIL.n114 9.3005
R536 VTAIL.n70 VTAIL.n69 9.3005
R537 VTAIL.n109 VTAIL.n108 9.3005
R538 VTAIL.n82 VTAIL.n81 9.3005
R539 VTAIL.n89 VTAIL.n88 9.3005
R540 VTAIL.n91 VTAIL.n90 9.3005
R541 VTAIL.n78 VTAIL.n77 9.3005
R542 VTAIL.n97 VTAIL.n96 9.3005
R543 VTAIL.n99 VTAIL.n98 9.3005
R544 VTAIL.n100 VTAIL.n73 9.3005
R545 VTAIL.n107 VTAIL.n106 9.3005
R546 VTAIL.n187 VTAIL.n186 9.3005
R547 VTAIL.n130 VTAIL.n129 9.3005
R548 VTAIL.n181 VTAIL.n180 9.3005
R549 VTAIL.n179 VTAIL.n178 9.3005
R550 VTAIL.n134 VTAIL.n133 9.3005
R551 VTAIL.n173 VTAIL.n172 9.3005
R552 VTAIL.n146 VTAIL.n145 9.3005
R553 VTAIL.n153 VTAIL.n152 9.3005
R554 VTAIL.n155 VTAIL.n154 9.3005
R555 VTAIL.n142 VTAIL.n141 9.3005
R556 VTAIL.n161 VTAIL.n160 9.3005
R557 VTAIL.n163 VTAIL.n162 9.3005
R558 VTAIL.n164 VTAIL.n137 9.3005
R559 VTAIL.n171 VTAIL.n170 9.3005
R560 VTAIL.n400 VTAIL.n399 9.3005
R561 VTAIL.n407 VTAIL.n406 9.3005
R562 VTAIL.n409 VTAIL.n408 9.3005
R563 VTAIL.n396 VTAIL.n395 9.3005
R564 VTAIL.n415 VTAIL.n414 9.3005
R565 VTAIL.n417 VTAIL.n416 9.3005
R566 VTAIL.n391 VTAIL.n389 9.3005
R567 VTAIL.n423 VTAIL.n422 9.3005
R568 VTAIL.n439 VTAIL.n438 9.3005
R569 VTAIL.n382 VTAIL.n381 9.3005
R570 VTAIL.n433 VTAIL.n432 9.3005
R571 VTAIL.n431 VTAIL.n430 9.3005
R572 VTAIL.n386 VTAIL.n385 9.3005
R573 VTAIL.n425 VTAIL.n424 9.3005
R574 VTAIL.n336 VTAIL.n335 9.3005
R575 VTAIL.n343 VTAIL.n342 9.3005
R576 VTAIL.n345 VTAIL.n344 9.3005
R577 VTAIL.n332 VTAIL.n331 9.3005
R578 VTAIL.n351 VTAIL.n350 9.3005
R579 VTAIL.n353 VTAIL.n352 9.3005
R580 VTAIL.n327 VTAIL.n325 9.3005
R581 VTAIL.n359 VTAIL.n358 9.3005
R582 VTAIL.n375 VTAIL.n374 9.3005
R583 VTAIL.n318 VTAIL.n317 9.3005
R584 VTAIL.n369 VTAIL.n368 9.3005
R585 VTAIL.n367 VTAIL.n366 9.3005
R586 VTAIL.n322 VTAIL.n321 9.3005
R587 VTAIL.n361 VTAIL.n360 9.3005
R588 VTAIL.n274 VTAIL.n273 9.3005
R589 VTAIL.n281 VTAIL.n280 9.3005
R590 VTAIL.n283 VTAIL.n282 9.3005
R591 VTAIL.n270 VTAIL.n269 9.3005
R592 VTAIL.n289 VTAIL.n288 9.3005
R593 VTAIL.n291 VTAIL.n290 9.3005
R594 VTAIL.n265 VTAIL.n263 9.3005
R595 VTAIL.n297 VTAIL.n296 9.3005
R596 VTAIL.n313 VTAIL.n312 9.3005
R597 VTAIL.n256 VTAIL.n255 9.3005
R598 VTAIL.n307 VTAIL.n306 9.3005
R599 VTAIL.n305 VTAIL.n304 9.3005
R600 VTAIL.n260 VTAIL.n259 9.3005
R601 VTAIL.n299 VTAIL.n298 9.3005
R602 VTAIL.n210 VTAIL.n209 9.3005
R603 VTAIL.n217 VTAIL.n216 9.3005
R604 VTAIL.n219 VTAIL.n218 9.3005
R605 VTAIL.n206 VTAIL.n205 9.3005
R606 VTAIL.n225 VTAIL.n224 9.3005
R607 VTAIL.n227 VTAIL.n226 9.3005
R608 VTAIL.n201 VTAIL.n199 9.3005
R609 VTAIL.n233 VTAIL.n232 9.3005
R610 VTAIL.n249 VTAIL.n248 9.3005
R611 VTAIL.n192 VTAIL.n191 9.3005
R612 VTAIL.n243 VTAIL.n242 9.3005
R613 VTAIL.n241 VTAIL.n240 9.3005
R614 VTAIL.n196 VTAIL.n195 9.3005
R615 VTAIL.n235 VTAIL.n234 9.3005
R616 VTAIL.n469 VTAIL.n458 8.92171
R617 VTAIL.n500 VTAIL.n442 8.92171
R618 VTAIL.n29 VTAIL.n18 8.92171
R619 VTAIL.n60 VTAIL.n2 8.92171
R620 VTAIL.n91 VTAIL.n80 8.92171
R621 VTAIL.n122 VTAIL.n64 8.92171
R622 VTAIL.n155 VTAIL.n144 8.92171
R623 VTAIL.n186 VTAIL.n128 8.92171
R624 VTAIL.n438 VTAIL.n380 8.92171
R625 VTAIL.n409 VTAIL.n398 8.92171
R626 VTAIL.n374 VTAIL.n316 8.92171
R627 VTAIL.n345 VTAIL.n334 8.92171
R628 VTAIL.n312 VTAIL.n254 8.92171
R629 VTAIL.n283 VTAIL.n272 8.92171
R630 VTAIL.n248 VTAIL.n190 8.92171
R631 VTAIL.n219 VTAIL.n208 8.92171
R632 VTAIL.n466 VTAIL.n465 8.14595
R633 VTAIL.n26 VTAIL.n25 8.14595
R634 VTAIL.n88 VTAIL.n87 8.14595
R635 VTAIL.n152 VTAIL.n151 8.14595
R636 VTAIL.n406 VTAIL.n405 8.14595
R637 VTAIL.n342 VTAIL.n341 8.14595
R638 VTAIL.n280 VTAIL.n279 8.14595
R639 VTAIL.n216 VTAIL.n215 8.14595
R640 VTAIL.n462 VTAIL.n460 7.3702
R641 VTAIL.n22 VTAIL.n20 7.3702
R642 VTAIL.n84 VTAIL.n82 7.3702
R643 VTAIL.n148 VTAIL.n146 7.3702
R644 VTAIL.n402 VTAIL.n400 7.3702
R645 VTAIL.n338 VTAIL.n336 7.3702
R646 VTAIL.n276 VTAIL.n274 7.3702
R647 VTAIL.n212 VTAIL.n210 7.3702
R648 VTAIL.n465 VTAIL.n460 5.81868
R649 VTAIL.n25 VTAIL.n20 5.81868
R650 VTAIL.n87 VTAIL.n82 5.81868
R651 VTAIL.n151 VTAIL.n146 5.81868
R652 VTAIL.n405 VTAIL.n400 5.81868
R653 VTAIL.n341 VTAIL.n336 5.81868
R654 VTAIL.n279 VTAIL.n274 5.81868
R655 VTAIL.n215 VTAIL.n210 5.81868
R656 VTAIL.n466 VTAIL.n458 5.04292
R657 VTAIL.n502 VTAIL.n442 5.04292
R658 VTAIL.n26 VTAIL.n18 5.04292
R659 VTAIL.n62 VTAIL.n2 5.04292
R660 VTAIL.n88 VTAIL.n80 5.04292
R661 VTAIL.n124 VTAIL.n64 5.04292
R662 VTAIL.n152 VTAIL.n144 5.04292
R663 VTAIL.n188 VTAIL.n128 5.04292
R664 VTAIL.n440 VTAIL.n380 5.04292
R665 VTAIL.n406 VTAIL.n398 5.04292
R666 VTAIL.n376 VTAIL.n316 5.04292
R667 VTAIL.n342 VTAIL.n334 5.04292
R668 VTAIL.n314 VTAIL.n254 5.04292
R669 VTAIL.n280 VTAIL.n272 5.04292
R670 VTAIL.n250 VTAIL.n190 5.04292
R671 VTAIL.n216 VTAIL.n208 5.04292
R672 VTAIL.n470 VTAIL.n469 4.26717
R673 VTAIL.n500 VTAIL.n499 4.26717
R674 VTAIL.n30 VTAIL.n29 4.26717
R675 VTAIL.n60 VTAIL.n59 4.26717
R676 VTAIL.n92 VTAIL.n91 4.26717
R677 VTAIL.n122 VTAIL.n121 4.26717
R678 VTAIL.n156 VTAIL.n155 4.26717
R679 VTAIL.n186 VTAIL.n185 4.26717
R680 VTAIL.n438 VTAIL.n437 4.26717
R681 VTAIL.n410 VTAIL.n409 4.26717
R682 VTAIL.n374 VTAIL.n373 4.26717
R683 VTAIL.n346 VTAIL.n345 4.26717
R684 VTAIL.n312 VTAIL.n311 4.26717
R685 VTAIL.n284 VTAIL.n283 4.26717
R686 VTAIL.n248 VTAIL.n247 4.26717
R687 VTAIL.n220 VTAIL.n219 4.26717
R688 VTAIL.n253 VTAIL.n251 3.56947
R689 VTAIL.n315 VTAIL.n253 3.56947
R690 VTAIL.n379 VTAIL.n377 3.56947
R691 VTAIL.n441 VTAIL.n379 3.56947
R692 VTAIL.n189 VTAIL.n127 3.56947
R693 VTAIL.n127 VTAIL.n125 3.56947
R694 VTAIL.n63 VTAIL.n1 3.56947
R695 VTAIL VTAIL.n503 3.51128
R696 VTAIL.n473 VTAIL.n456 3.49141
R697 VTAIL.n496 VTAIL.n444 3.49141
R698 VTAIL.n33 VTAIL.n16 3.49141
R699 VTAIL.n56 VTAIL.n4 3.49141
R700 VTAIL.n95 VTAIL.n78 3.49141
R701 VTAIL.n118 VTAIL.n66 3.49141
R702 VTAIL.n159 VTAIL.n142 3.49141
R703 VTAIL.n182 VTAIL.n130 3.49141
R704 VTAIL.n434 VTAIL.n382 3.49141
R705 VTAIL.n413 VTAIL.n396 3.49141
R706 VTAIL.n370 VTAIL.n318 3.49141
R707 VTAIL.n349 VTAIL.n332 3.49141
R708 VTAIL.n308 VTAIL.n256 3.49141
R709 VTAIL.n287 VTAIL.n270 3.49141
R710 VTAIL.n244 VTAIL.n192 3.49141
R711 VTAIL.n223 VTAIL.n206 3.49141
R712 VTAIL.n461 VTAIL.n459 2.84303
R713 VTAIL.n21 VTAIL.n19 2.84303
R714 VTAIL.n83 VTAIL.n81 2.84303
R715 VTAIL.n147 VTAIL.n145 2.84303
R716 VTAIL.n401 VTAIL.n399 2.84303
R717 VTAIL.n337 VTAIL.n335 2.84303
R718 VTAIL.n275 VTAIL.n273 2.84303
R719 VTAIL.n211 VTAIL.n209 2.84303
R720 VTAIL.n474 VTAIL.n454 2.71565
R721 VTAIL.n495 VTAIL.n446 2.71565
R722 VTAIL.n34 VTAIL.n14 2.71565
R723 VTAIL.n55 VTAIL.n6 2.71565
R724 VTAIL.n96 VTAIL.n76 2.71565
R725 VTAIL.n117 VTAIL.n68 2.71565
R726 VTAIL.n160 VTAIL.n140 2.71565
R727 VTAIL.n181 VTAIL.n132 2.71565
R728 VTAIL.n433 VTAIL.n384 2.71565
R729 VTAIL.n414 VTAIL.n394 2.71565
R730 VTAIL.n369 VTAIL.n320 2.71565
R731 VTAIL.n350 VTAIL.n330 2.71565
R732 VTAIL.n307 VTAIL.n258 2.71565
R733 VTAIL.n288 VTAIL.n268 2.71565
R734 VTAIL.n243 VTAIL.n194 2.71565
R735 VTAIL.n224 VTAIL.n204 2.71565
R736 VTAIL.n479 VTAIL.n477 1.93989
R737 VTAIL.n492 VTAIL.n491 1.93989
R738 VTAIL.n39 VTAIL.n37 1.93989
R739 VTAIL.n52 VTAIL.n51 1.93989
R740 VTAIL.n101 VTAIL.n99 1.93989
R741 VTAIL.n114 VTAIL.n113 1.93989
R742 VTAIL.n165 VTAIL.n163 1.93989
R743 VTAIL.n178 VTAIL.n177 1.93989
R744 VTAIL.n430 VTAIL.n429 1.93989
R745 VTAIL.n418 VTAIL.n417 1.93989
R746 VTAIL.n366 VTAIL.n365 1.93989
R747 VTAIL.n354 VTAIL.n353 1.93989
R748 VTAIL.n304 VTAIL.n303 1.93989
R749 VTAIL.n292 VTAIL.n291 1.93989
R750 VTAIL.n240 VTAIL.n239 1.93989
R751 VTAIL.n228 VTAIL.n227 1.93989
R752 VTAIL.n0 VTAIL.t8 1.73127
R753 VTAIL.n0 VTAIL.t14 1.73127
R754 VTAIL.n126 VTAIL.t5 1.73127
R755 VTAIL.n126 VTAIL.t1 1.73127
R756 VTAIL.n378 VTAIL.t6 1.73127
R757 VTAIL.n378 VTAIL.t4 1.73127
R758 VTAIL.n252 VTAIL.t10 1.73127
R759 VTAIL.n252 VTAIL.t15 1.73127
R760 VTAIL.n478 VTAIL.n452 1.16414
R761 VTAIL.n488 VTAIL.n448 1.16414
R762 VTAIL.n38 VTAIL.n12 1.16414
R763 VTAIL.n48 VTAIL.n8 1.16414
R764 VTAIL.n100 VTAIL.n74 1.16414
R765 VTAIL.n110 VTAIL.n70 1.16414
R766 VTAIL.n164 VTAIL.n138 1.16414
R767 VTAIL.n174 VTAIL.n134 1.16414
R768 VTAIL.n426 VTAIL.n386 1.16414
R769 VTAIL.n421 VTAIL.n391 1.16414
R770 VTAIL.n362 VTAIL.n322 1.16414
R771 VTAIL.n357 VTAIL.n327 1.16414
R772 VTAIL.n300 VTAIL.n260 1.16414
R773 VTAIL.n295 VTAIL.n265 1.16414
R774 VTAIL.n236 VTAIL.n196 1.16414
R775 VTAIL.n231 VTAIL.n201 1.16414
R776 VTAIL.n377 VTAIL.n315 0.470328
R777 VTAIL.n125 VTAIL.n63 0.470328
R778 VTAIL.n484 VTAIL.n483 0.388379
R779 VTAIL.n487 VTAIL.n450 0.388379
R780 VTAIL.n44 VTAIL.n43 0.388379
R781 VTAIL.n47 VTAIL.n10 0.388379
R782 VTAIL.n106 VTAIL.n105 0.388379
R783 VTAIL.n109 VTAIL.n72 0.388379
R784 VTAIL.n170 VTAIL.n169 0.388379
R785 VTAIL.n173 VTAIL.n136 0.388379
R786 VTAIL.n425 VTAIL.n388 0.388379
R787 VTAIL.n422 VTAIL.n390 0.388379
R788 VTAIL.n361 VTAIL.n324 0.388379
R789 VTAIL.n358 VTAIL.n326 0.388379
R790 VTAIL.n299 VTAIL.n262 0.388379
R791 VTAIL.n296 VTAIL.n264 0.388379
R792 VTAIL.n235 VTAIL.n198 0.388379
R793 VTAIL.n232 VTAIL.n200 0.388379
R794 VTAIL.n467 VTAIL.n459 0.155672
R795 VTAIL.n468 VTAIL.n467 0.155672
R796 VTAIL.n468 VTAIL.n455 0.155672
R797 VTAIL.n475 VTAIL.n455 0.155672
R798 VTAIL.n476 VTAIL.n475 0.155672
R799 VTAIL.n476 VTAIL.n451 0.155672
R800 VTAIL.n485 VTAIL.n451 0.155672
R801 VTAIL.n486 VTAIL.n485 0.155672
R802 VTAIL.n486 VTAIL.n447 0.155672
R803 VTAIL.n493 VTAIL.n447 0.155672
R804 VTAIL.n494 VTAIL.n493 0.155672
R805 VTAIL.n494 VTAIL.n443 0.155672
R806 VTAIL.n501 VTAIL.n443 0.155672
R807 VTAIL.n27 VTAIL.n19 0.155672
R808 VTAIL.n28 VTAIL.n27 0.155672
R809 VTAIL.n28 VTAIL.n15 0.155672
R810 VTAIL.n35 VTAIL.n15 0.155672
R811 VTAIL.n36 VTAIL.n35 0.155672
R812 VTAIL.n36 VTAIL.n11 0.155672
R813 VTAIL.n45 VTAIL.n11 0.155672
R814 VTAIL.n46 VTAIL.n45 0.155672
R815 VTAIL.n46 VTAIL.n7 0.155672
R816 VTAIL.n53 VTAIL.n7 0.155672
R817 VTAIL.n54 VTAIL.n53 0.155672
R818 VTAIL.n54 VTAIL.n3 0.155672
R819 VTAIL.n61 VTAIL.n3 0.155672
R820 VTAIL.n89 VTAIL.n81 0.155672
R821 VTAIL.n90 VTAIL.n89 0.155672
R822 VTAIL.n90 VTAIL.n77 0.155672
R823 VTAIL.n97 VTAIL.n77 0.155672
R824 VTAIL.n98 VTAIL.n97 0.155672
R825 VTAIL.n98 VTAIL.n73 0.155672
R826 VTAIL.n107 VTAIL.n73 0.155672
R827 VTAIL.n108 VTAIL.n107 0.155672
R828 VTAIL.n108 VTAIL.n69 0.155672
R829 VTAIL.n115 VTAIL.n69 0.155672
R830 VTAIL.n116 VTAIL.n115 0.155672
R831 VTAIL.n116 VTAIL.n65 0.155672
R832 VTAIL.n123 VTAIL.n65 0.155672
R833 VTAIL.n153 VTAIL.n145 0.155672
R834 VTAIL.n154 VTAIL.n153 0.155672
R835 VTAIL.n154 VTAIL.n141 0.155672
R836 VTAIL.n161 VTAIL.n141 0.155672
R837 VTAIL.n162 VTAIL.n161 0.155672
R838 VTAIL.n162 VTAIL.n137 0.155672
R839 VTAIL.n171 VTAIL.n137 0.155672
R840 VTAIL.n172 VTAIL.n171 0.155672
R841 VTAIL.n172 VTAIL.n133 0.155672
R842 VTAIL.n179 VTAIL.n133 0.155672
R843 VTAIL.n180 VTAIL.n179 0.155672
R844 VTAIL.n180 VTAIL.n129 0.155672
R845 VTAIL.n187 VTAIL.n129 0.155672
R846 VTAIL.n439 VTAIL.n381 0.155672
R847 VTAIL.n432 VTAIL.n381 0.155672
R848 VTAIL.n432 VTAIL.n431 0.155672
R849 VTAIL.n431 VTAIL.n385 0.155672
R850 VTAIL.n424 VTAIL.n385 0.155672
R851 VTAIL.n424 VTAIL.n423 0.155672
R852 VTAIL.n423 VTAIL.n389 0.155672
R853 VTAIL.n416 VTAIL.n389 0.155672
R854 VTAIL.n416 VTAIL.n415 0.155672
R855 VTAIL.n415 VTAIL.n395 0.155672
R856 VTAIL.n408 VTAIL.n395 0.155672
R857 VTAIL.n408 VTAIL.n407 0.155672
R858 VTAIL.n407 VTAIL.n399 0.155672
R859 VTAIL.n375 VTAIL.n317 0.155672
R860 VTAIL.n368 VTAIL.n317 0.155672
R861 VTAIL.n368 VTAIL.n367 0.155672
R862 VTAIL.n367 VTAIL.n321 0.155672
R863 VTAIL.n360 VTAIL.n321 0.155672
R864 VTAIL.n360 VTAIL.n359 0.155672
R865 VTAIL.n359 VTAIL.n325 0.155672
R866 VTAIL.n352 VTAIL.n325 0.155672
R867 VTAIL.n352 VTAIL.n351 0.155672
R868 VTAIL.n351 VTAIL.n331 0.155672
R869 VTAIL.n344 VTAIL.n331 0.155672
R870 VTAIL.n344 VTAIL.n343 0.155672
R871 VTAIL.n343 VTAIL.n335 0.155672
R872 VTAIL.n313 VTAIL.n255 0.155672
R873 VTAIL.n306 VTAIL.n255 0.155672
R874 VTAIL.n306 VTAIL.n305 0.155672
R875 VTAIL.n305 VTAIL.n259 0.155672
R876 VTAIL.n298 VTAIL.n259 0.155672
R877 VTAIL.n298 VTAIL.n297 0.155672
R878 VTAIL.n297 VTAIL.n263 0.155672
R879 VTAIL.n290 VTAIL.n263 0.155672
R880 VTAIL.n290 VTAIL.n289 0.155672
R881 VTAIL.n289 VTAIL.n269 0.155672
R882 VTAIL.n282 VTAIL.n269 0.155672
R883 VTAIL.n282 VTAIL.n281 0.155672
R884 VTAIL.n281 VTAIL.n273 0.155672
R885 VTAIL.n249 VTAIL.n191 0.155672
R886 VTAIL.n242 VTAIL.n191 0.155672
R887 VTAIL.n242 VTAIL.n241 0.155672
R888 VTAIL.n241 VTAIL.n195 0.155672
R889 VTAIL.n234 VTAIL.n195 0.155672
R890 VTAIL.n234 VTAIL.n233 0.155672
R891 VTAIL.n233 VTAIL.n199 0.155672
R892 VTAIL.n226 VTAIL.n199 0.155672
R893 VTAIL.n226 VTAIL.n225 0.155672
R894 VTAIL.n225 VTAIL.n205 0.155672
R895 VTAIL.n218 VTAIL.n205 0.155672
R896 VTAIL.n218 VTAIL.n217 0.155672
R897 VTAIL.n217 VTAIL.n209 0.155672
R898 VTAIL VTAIL.n1 0.0586897
R899 B.n1015 B.n1014 585
R900 B.n353 B.n170 585
R901 B.n352 B.n351 585
R902 B.n350 B.n349 585
R903 B.n348 B.n347 585
R904 B.n346 B.n345 585
R905 B.n344 B.n343 585
R906 B.n342 B.n341 585
R907 B.n340 B.n339 585
R908 B.n338 B.n337 585
R909 B.n336 B.n335 585
R910 B.n334 B.n333 585
R911 B.n332 B.n331 585
R912 B.n330 B.n329 585
R913 B.n328 B.n327 585
R914 B.n326 B.n325 585
R915 B.n324 B.n323 585
R916 B.n322 B.n321 585
R917 B.n320 B.n319 585
R918 B.n318 B.n317 585
R919 B.n316 B.n315 585
R920 B.n314 B.n313 585
R921 B.n312 B.n311 585
R922 B.n310 B.n309 585
R923 B.n308 B.n307 585
R924 B.n306 B.n305 585
R925 B.n304 B.n303 585
R926 B.n302 B.n301 585
R927 B.n300 B.n299 585
R928 B.n298 B.n297 585
R929 B.n296 B.n295 585
R930 B.n294 B.n293 585
R931 B.n292 B.n291 585
R932 B.n290 B.n289 585
R933 B.n288 B.n287 585
R934 B.n286 B.n285 585
R935 B.n284 B.n283 585
R936 B.n282 B.n281 585
R937 B.n280 B.n279 585
R938 B.n278 B.n277 585
R939 B.n276 B.n275 585
R940 B.n274 B.n273 585
R941 B.n272 B.n271 585
R942 B.n270 B.n269 585
R943 B.n268 B.n267 585
R944 B.n266 B.n265 585
R945 B.n264 B.n263 585
R946 B.n262 B.n261 585
R947 B.n260 B.n259 585
R948 B.n258 B.n257 585
R949 B.n256 B.n255 585
R950 B.n254 B.n253 585
R951 B.n252 B.n251 585
R952 B.n250 B.n249 585
R953 B.n248 B.n247 585
R954 B.n246 B.n245 585
R955 B.n244 B.n243 585
R956 B.n242 B.n241 585
R957 B.n240 B.n239 585
R958 B.n238 B.n237 585
R959 B.n236 B.n235 585
R960 B.n234 B.n233 585
R961 B.n232 B.n231 585
R962 B.n230 B.n229 585
R963 B.n228 B.n227 585
R964 B.n226 B.n225 585
R965 B.n224 B.n223 585
R966 B.n222 B.n221 585
R967 B.n220 B.n219 585
R968 B.n218 B.n217 585
R969 B.n216 B.n215 585
R970 B.n214 B.n213 585
R971 B.n212 B.n211 585
R972 B.n210 B.n209 585
R973 B.n208 B.n207 585
R974 B.n206 B.n205 585
R975 B.n204 B.n203 585
R976 B.n202 B.n201 585
R977 B.n200 B.n199 585
R978 B.n198 B.n197 585
R979 B.n196 B.n195 585
R980 B.n194 B.n193 585
R981 B.n192 B.n191 585
R982 B.n190 B.n189 585
R983 B.n188 B.n187 585
R984 B.n186 B.n185 585
R985 B.n184 B.n183 585
R986 B.n182 B.n181 585
R987 B.n180 B.n179 585
R988 B.n178 B.n177 585
R989 B.n1013 B.n125 585
R990 B.n1018 B.n125 585
R991 B.n1012 B.n124 585
R992 B.n1019 B.n124 585
R993 B.n1011 B.n1010 585
R994 B.n1010 B.n120 585
R995 B.n1009 B.n119 585
R996 B.n1025 B.n119 585
R997 B.n1008 B.n118 585
R998 B.n1026 B.n118 585
R999 B.n1007 B.n117 585
R1000 B.n1027 B.n117 585
R1001 B.n1006 B.n1005 585
R1002 B.n1005 B.n113 585
R1003 B.n1004 B.n112 585
R1004 B.n1033 B.n112 585
R1005 B.n1003 B.n111 585
R1006 B.n1034 B.n111 585
R1007 B.n1002 B.n110 585
R1008 B.n1035 B.n110 585
R1009 B.n1001 B.n1000 585
R1010 B.n1000 B.n106 585
R1011 B.n999 B.n105 585
R1012 B.n1041 B.n105 585
R1013 B.n998 B.n104 585
R1014 B.n1042 B.n104 585
R1015 B.n997 B.n103 585
R1016 B.n1043 B.n103 585
R1017 B.n996 B.n995 585
R1018 B.n995 B.n99 585
R1019 B.n994 B.n98 585
R1020 B.n1049 B.n98 585
R1021 B.n993 B.n97 585
R1022 B.n1050 B.n97 585
R1023 B.n992 B.n96 585
R1024 B.n1051 B.n96 585
R1025 B.n991 B.n990 585
R1026 B.n990 B.n92 585
R1027 B.n989 B.n91 585
R1028 B.n1057 B.n91 585
R1029 B.n988 B.n90 585
R1030 B.n1058 B.n90 585
R1031 B.n987 B.n89 585
R1032 B.n1059 B.n89 585
R1033 B.n986 B.n985 585
R1034 B.n985 B.n85 585
R1035 B.n984 B.n84 585
R1036 B.n1065 B.n84 585
R1037 B.n983 B.n83 585
R1038 B.n1066 B.n83 585
R1039 B.n982 B.n82 585
R1040 B.n1067 B.n82 585
R1041 B.n981 B.n980 585
R1042 B.n980 B.n78 585
R1043 B.n979 B.n77 585
R1044 B.n1073 B.n77 585
R1045 B.n978 B.n76 585
R1046 B.n1074 B.n76 585
R1047 B.n977 B.n75 585
R1048 B.n1075 B.n75 585
R1049 B.n976 B.n975 585
R1050 B.n975 B.n71 585
R1051 B.n974 B.n70 585
R1052 B.n1081 B.n70 585
R1053 B.n973 B.n69 585
R1054 B.n1082 B.n69 585
R1055 B.n972 B.n68 585
R1056 B.n1083 B.n68 585
R1057 B.n971 B.n970 585
R1058 B.n970 B.n64 585
R1059 B.n969 B.n63 585
R1060 B.n1089 B.n63 585
R1061 B.n968 B.n62 585
R1062 B.n1090 B.n62 585
R1063 B.n967 B.n61 585
R1064 B.n1091 B.n61 585
R1065 B.n966 B.n965 585
R1066 B.n965 B.n57 585
R1067 B.n964 B.n56 585
R1068 B.n1097 B.n56 585
R1069 B.n963 B.n55 585
R1070 B.n1098 B.n55 585
R1071 B.n962 B.n54 585
R1072 B.n1099 B.n54 585
R1073 B.n961 B.n960 585
R1074 B.n960 B.n50 585
R1075 B.n959 B.n49 585
R1076 B.n1105 B.n49 585
R1077 B.n958 B.n48 585
R1078 B.n1106 B.n48 585
R1079 B.n957 B.n47 585
R1080 B.n1107 B.n47 585
R1081 B.n956 B.n955 585
R1082 B.n955 B.n43 585
R1083 B.n954 B.n42 585
R1084 B.n1113 B.n42 585
R1085 B.n953 B.n41 585
R1086 B.n1114 B.n41 585
R1087 B.n952 B.n40 585
R1088 B.n1115 B.n40 585
R1089 B.n951 B.n950 585
R1090 B.n950 B.n36 585
R1091 B.n949 B.n35 585
R1092 B.n1121 B.n35 585
R1093 B.n948 B.n34 585
R1094 B.n1122 B.n34 585
R1095 B.n947 B.n33 585
R1096 B.n1123 B.n33 585
R1097 B.n946 B.n945 585
R1098 B.n945 B.n29 585
R1099 B.n944 B.n28 585
R1100 B.n1129 B.n28 585
R1101 B.n943 B.n27 585
R1102 B.n1130 B.n27 585
R1103 B.n942 B.n26 585
R1104 B.n1131 B.n26 585
R1105 B.n941 B.n940 585
R1106 B.n940 B.n22 585
R1107 B.n939 B.n21 585
R1108 B.n1137 B.n21 585
R1109 B.n938 B.n20 585
R1110 B.n1138 B.n20 585
R1111 B.n937 B.n19 585
R1112 B.n1139 B.n19 585
R1113 B.n936 B.n935 585
R1114 B.n935 B.n15 585
R1115 B.n934 B.n14 585
R1116 B.n1145 B.n14 585
R1117 B.n933 B.n13 585
R1118 B.n1146 B.n13 585
R1119 B.n932 B.n12 585
R1120 B.n1147 B.n12 585
R1121 B.n931 B.n930 585
R1122 B.n930 B.n8 585
R1123 B.n929 B.n7 585
R1124 B.n1153 B.n7 585
R1125 B.n928 B.n6 585
R1126 B.n1154 B.n6 585
R1127 B.n927 B.n5 585
R1128 B.n1155 B.n5 585
R1129 B.n926 B.n925 585
R1130 B.n925 B.n4 585
R1131 B.n924 B.n354 585
R1132 B.n924 B.n923 585
R1133 B.n914 B.n355 585
R1134 B.n356 B.n355 585
R1135 B.n916 B.n915 585
R1136 B.n917 B.n916 585
R1137 B.n913 B.n361 585
R1138 B.n361 B.n360 585
R1139 B.n912 B.n911 585
R1140 B.n911 B.n910 585
R1141 B.n363 B.n362 585
R1142 B.n364 B.n363 585
R1143 B.n903 B.n902 585
R1144 B.n904 B.n903 585
R1145 B.n901 B.n369 585
R1146 B.n369 B.n368 585
R1147 B.n900 B.n899 585
R1148 B.n899 B.n898 585
R1149 B.n371 B.n370 585
R1150 B.n372 B.n371 585
R1151 B.n891 B.n890 585
R1152 B.n892 B.n891 585
R1153 B.n889 B.n377 585
R1154 B.n377 B.n376 585
R1155 B.n888 B.n887 585
R1156 B.n887 B.n886 585
R1157 B.n379 B.n378 585
R1158 B.n380 B.n379 585
R1159 B.n879 B.n878 585
R1160 B.n880 B.n879 585
R1161 B.n877 B.n385 585
R1162 B.n385 B.n384 585
R1163 B.n876 B.n875 585
R1164 B.n875 B.n874 585
R1165 B.n387 B.n386 585
R1166 B.n388 B.n387 585
R1167 B.n867 B.n866 585
R1168 B.n868 B.n867 585
R1169 B.n865 B.n393 585
R1170 B.n393 B.n392 585
R1171 B.n864 B.n863 585
R1172 B.n863 B.n862 585
R1173 B.n395 B.n394 585
R1174 B.n396 B.n395 585
R1175 B.n855 B.n854 585
R1176 B.n856 B.n855 585
R1177 B.n853 B.n401 585
R1178 B.n401 B.n400 585
R1179 B.n852 B.n851 585
R1180 B.n851 B.n850 585
R1181 B.n403 B.n402 585
R1182 B.n404 B.n403 585
R1183 B.n843 B.n842 585
R1184 B.n844 B.n843 585
R1185 B.n841 B.n409 585
R1186 B.n409 B.n408 585
R1187 B.n840 B.n839 585
R1188 B.n839 B.n838 585
R1189 B.n411 B.n410 585
R1190 B.n412 B.n411 585
R1191 B.n831 B.n830 585
R1192 B.n832 B.n831 585
R1193 B.n829 B.n416 585
R1194 B.n420 B.n416 585
R1195 B.n828 B.n827 585
R1196 B.n827 B.n826 585
R1197 B.n418 B.n417 585
R1198 B.n419 B.n418 585
R1199 B.n819 B.n818 585
R1200 B.n820 B.n819 585
R1201 B.n817 B.n425 585
R1202 B.n425 B.n424 585
R1203 B.n816 B.n815 585
R1204 B.n815 B.n814 585
R1205 B.n427 B.n426 585
R1206 B.n428 B.n427 585
R1207 B.n807 B.n806 585
R1208 B.n808 B.n807 585
R1209 B.n805 B.n433 585
R1210 B.n433 B.n432 585
R1211 B.n804 B.n803 585
R1212 B.n803 B.n802 585
R1213 B.n435 B.n434 585
R1214 B.n436 B.n435 585
R1215 B.n795 B.n794 585
R1216 B.n796 B.n795 585
R1217 B.n793 B.n440 585
R1218 B.n444 B.n440 585
R1219 B.n792 B.n791 585
R1220 B.n791 B.n790 585
R1221 B.n442 B.n441 585
R1222 B.n443 B.n442 585
R1223 B.n783 B.n782 585
R1224 B.n784 B.n783 585
R1225 B.n781 B.n449 585
R1226 B.n449 B.n448 585
R1227 B.n780 B.n779 585
R1228 B.n779 B.n778 585
R1229 B.n451 B.n450 585
R1230 B.n452 B.n451 585
R1231 B.n771 B.n770 585
R1232 B.n772 B.n771 585
R1233 B.n769 B.n457 585
R1234 B.n457 B.n456 585
R1235 B.n768 B.n767 585
R1236 B.n767 B.n766 585
R1237 B.n459 B.n458 585
R1238 B.n460 B.n459 585
R1239 B.n759 B.n758 585
R1240 B.n760 B.n759 585
R1241 B.n757 B.n465 585
R1242 B.n465 B.n464 585
R1243 B.n756 B.n755 585
R1244 B.n755 B.n754 585
R1245 B.n467 B.n466 585
R1246 B.n468 B.n467 585
R1247 B.n747 B.n746 585
R1248 B.n748 B.n747 585
R1249 B.n745 B.n473 585
R1250 B.n473 B.n472 585
R1251 B.n744 B.n743 585
R1252 B.n743 B.n742 585
R1253 B.n475 B.n474 585
R1254 B.n476 B.n475 585
R1255 B.n735 B.n734 585
R1256 B.n736 B.n735 585
R1257 B.n733 B.n481 585
R1258 B.n481 B.n480 585
R1259 B.n732 B.n731 585
R1260 B.n731 B.n730 585
R1261 B.n483 B.n482 585
R1262 B.n484 B.n483 585
R1263 B.n723 B.n722 585
R1264 B.n724 B.n723 585
R1265 B.n721 B.n489 585
R1266 B.n489 B.n488 585
R1267 B.n716 B.n715 585
R1268 B.n714 B.n536 585
R1269 B.n713 B.n535 585
R1270 B.n718 B.n535 585
R1271 B.n712 B.n711 585
R1272 B.n710 B.n709 585
R1273 B.n708 B.n707 585
R1274 B.n706 B.n705 585
R1275 B.n704 B.n703 585
R1276 B.n702 B.n701 585
R1277 B.n700 B.n699 585
R1278 B.n698 B.n697 585
R1279 B.n696 B.n695 585
R1280 B.n694 B.n693 585
R1281 B.n692 B.n691 585
R1282 B.n690 B.n689 585
R1283 B.n688 B.n687 585
R1284 B.n686 B.n685 585
R1285 B.n684 B.n683 585
R1286 B.n682 B.n681 585
R1287 B.n680 B.n679 585
R1288 B.n678 B.n677 585
R1289 B.n676 B.n675 585
R1290 B.n674 B.n673 585
R1291 B.n672 B.n671 585
R1292 B.n670 B.n669 585
R1293 B.n668 B.n667 585
R1294 B.n666 B.n665 585
R1295 B.n664 B.n663 585
R1296 B.n662 B.n661 585
R1297 B.n660 B.n659 585
R1298 B.n658 B.n657 585
R1299 B.n656 B.n655 585
R1300 B.n654 B.n653 585
R1301 B.n652 B.n651 585
R1302 B.n650 B.n649 585
R1303 B.n648 B.n647 585
R1304 B.n646 B.n645 585
R1305 B.n644 B.n643 585
R1306 B.n642 B.n641 585
R1307 B.n640 B.n639 585
R1308 B.n637 B.n636 585
R1309 B.n635 B.n634 585
R1310 B.n633 B.n632 585
R1311 B.n631 B.n630 585
R1312 B.n629 B.n628 585
R1313 B.n627 B.n626 585
R1314 B.n625 B.n624 585
R1315 B.n623 B.n622 585
R1316 B.n621 B.n620 585
R1317 B.n619 B.n618 585
R1318 B.n616 B.n615 585
R1319 B.n614 B.n613 585
R1320 B.n612 B.n611 585
R1321 B.n610 B.n609 585
R1322 B.n608 B.n607 585
R1323 B.n606 B.n605 585
R1324 B.n604 B.n603 585
R1325 B.n602 B.n601 585
R1326 B.n600 B.n599 585
R1327 B.n598 B.n597 585
R1328 B.n596 B.n595 585
R1329 B.n594 B.n593 585
R1330 B.n592 B.n591 585
R1331 B.n590 B.n589 585
R1332 B.n588 B.n587 585
R1333 B.n586 B.n585 585
R1334 B.n584 B.n583 585
R1335 B.n582 B.n581 585
R1336 B.n580 B.n579 585
R1337 B.n578 B.n577 585
R1338 B.n576 B.n575 585
R1339 B.n574 B.n573 585
R1340 B.n572 B.n571 585
R1341 B.n570 B.n569 585
R1342 B.n568 B.n567 585
R1343 B.n566 B.n565 585
R1344 B.n564 B.n563 585
R1345 B.n562 B.n561 585
R1346 B.n560 B.n559 585
R1347 B.n558 B.n557 585
R1348 B.n556 B.n555 585
R1349 B.n554 B.n553 585
R1350 B.n552 B.n551 585
R1351 B.n550 B.n549 585
R1352 B.n548 B.n547 585
R1353 B.n546 B.n545 585
R1354 B.n544 B.n543 585
R1355 B.n542 B.n541 585
R1356 B.n491 B.n490 585
R1357 B.n720 B.n719 585
R1358 B.n719 B.n718 585
R1359 B.n487 B.n486 585
R1360 B.n488 B.n487 585
R1361 B.n726 B.n725 585
R1362 B.n725 B.n724 585
R1363 B.n727 B.n485 585
R1364 B.n485 B.n484 585
R1365 B.n729 B.n728 585
R1366 B.n730 B.n729 585
R1367 B.n479 B.n478 585
R1368 B.n480 B.n479 585
R1369 B.n738 B.n737 585
R1370 B.n737 B.n736 585
R1371 B.n739 B.n477 585
R1372 B.n477 B.n476 585
R1373 B.n741 B.n740 585
R1374 B.n742 B.n741 585
R1375 B.n471 B.n470 585
R1376 B.n472 B.n471 585
R1377 B.n750 B.n749 585
R1378 B.n749 B.n748 585
R1379 B.n751 B.n469 585
R1380 B.n469 B.n468 585
R1381 B.n753 B.n752 585
R1382 B.n754 B.n753 585
R1383 B.n463 B.n462 585
R1384 B.n464 B.n463 585
R1385 B.n762 B.n761 585
R1386 B.n761 B.n760 585
R1387 B.n763 B.n461 585
R1388 B.n461 B.n460 585
R1389 B.n765 B.n764 585
R1390 B.n766 B.n765 585
R1391 B.n455 B.n454 585
R1392 B.n456 B.n455 585
R1393 B.n774 B.n773 585
R1394 B.n773 B.n772 585
R1395 B.n775 B.n453 585
R1396 B.n453 B.n452 585
R1397 B.n777 B.n776 585
R1398 B.n778 B.n777 585
R1399 B.n447 B.n446 585
R1400 B.n448 B.n447 585
R1401 B.n786 B.n785 585
R1402 B.n785 B.n784 585
R1403 B.n787 B.n445 585
R1404 B.n445 B.n443 585
R1405 B.n789 B.n788 585
R1406 B.n790 B.n789 585
R1407 B.n439 B.n438 585
R1408 B.n444 B.n439 585
R1409 B.n798 B.n797 585
R1410 B.n797 B.n796 585
R1411 B.n799 B.n437 585
R1412 B.n437 B.n436 585
R1413 B.n801 B.n800 585
R1414 B.n802 B.n801 585
R1415 B.n431 B.n430 585
R1416 B.n432 B.n431 585
R1417 B.n810 B.n809 585
R1418 B.n809 B.n808 585
R1419 B.n811 B.n429 585
R1420 B.n429 B.n428 585
R1421 B.n813 B.n812 585
R1422 B.n814 B.n813 585
R1423 B.n423 B.n422 585
R1424 B.n424 B.n423 585
R1425 B.n822 B.n821 585
R1426 B.n821 B.n820 585
R1427 B.n823 B.n421 585
R1428 B.n421 B.n419 585
R1429 B.n825 B.n824 585
R1430 B.n826 B.n825 585
R1431 B.n415 B.n414 585
R1432 B.n420 B.n415 585
R1433 B.n834 B.n833 585
R1434 B.n833 B.n832 585
R1435 B.n835 B.n413 585
R1436 B.n413 B.n412 585
R1437 B.n837 B.n836 585
R1438 B.n838 B.n837 585
R1439 B.n407 B.n406 585
R1440 B.n408 B.n407 585
R1441 B.n846 B.n845 585
R1442 B.n845 B.n844 585
R1443 B.n847 B.n405 585
R1444 B.n405 B.n404 585
R1445 B.n849 B.n848 585
R1446 B.n850 B.n849 585
R1447 B.n399 B.n398 585
R1448 B.n400 B.n399 585
R1449 B.n858 B.n857 585
R1450 B.n857 B.n856 585
R1451 B.n859 B.n397 585
R1452 B.n397 B.n396 585
R1453 B.n861 B.n860 585
R1454 B.n862 B.n861 585
R1455 B.n391 B.n390 585
R1456 B.n392 B.n391 585
R1457 B.n870 B.n869 585
R1458 B.n869 B.n868 585
R1459 B.n871 B.n389 585
R1460 B.n389 B.n388 585
R1461 B.n873 B.n872 585
R1462 B.n874 B.n873 585
R1463 B.n383 B.n382 585
R1464 B.n384 B.n383 585
R1465 B.n882 B.n881 585
R1466 B.n881 B.n880 585
R1467 B.n883 B.n381 585
R1468 B.n381 B.n380 585
R1469 B.n885 B.n884 585
R1470 B.n886 B.n885 585
R1471 B.n375 B.n374 585
R1472 B.n376 B.n375 585
R1473 B.n894 B.n893 585
R1474 B.n893 B.n892 585
R1475 B.n895 B.n373 585
R1476 B.n373 B.n372 585
R1477 B.n897 B.n896 585
R1478 B.n898 B.n897 585
R1479 B.n367 B.n366 585
R1480 B.n368 B.n367 585
R1481 B.n906 B.n905 585
R1482 B.n905 B.n904 585
R1483 B.n907 B.n365 585
R1484 B.n365 B.n364 585
R1485 B.n909 B.n908 585
R1486 B.n910 B.n909 585
R1487 B.n359 B.n358 585
R1488 B.n360 B.n359 585
R1489 B.n919 B.n918 585
R1490 B.n918 B.n917 585
R1491 B.n920 B.n357 585
R1492 B.n357 B.n356 585
R1493 B.n922 B.n921 585
R1494 B.n923 B.n922 585
R1495 B.n2 B.n0 585
R1496 B.n4 B.n2 585
R1497 B.n3 B.n1 585
R1498 B.n1154 B.n3 585
R1499 B.n1152 B.n1151 585
R1500 B.n1153 B.n1152 585
R1501 B.n1150 B.n9 585
R1502 B.n9 B.n8 585
R1503 B.n1149 B.n1148 585
R1504 B.n1148 B.n1147 585
R1505 B.n11 B.n10 585
R1506 B.n1146 B.n11 585
R1507 B.n1144 B.n1143 585
R1508 B.n1145 B.n1144 585
R1509 B.n1142 B.n16 585
R1510 B.n16 B.n15 585
R1511 B.n1141 B.n1140 585
R1512 B.n1140 B.n1139 585
R1513 B.n18 B.n17 585
R1514 B.n1138 B.n18 585
R1515 B.n1136 B.n1135 585
R1516 B.n1137 B.n1136 585
R1517 B.n1134 B.n23 585
R1518 B.n23 B.n22 585
R1519 B.n1133 B.n1132 585
R1520 B.n1132 B.n1131 585
R1521 B.n25 B.n24 585
R1522 B.n1130 B.n25 585
R1523 B.n1128 B.n1127 585
R1524 B.n1129 B.n1128 585
R1525 B.n1126 B.n30 585
R1526 B.n30 B.n29 585
R1527 B.n1125 B.n1124 585
R1528 B.n1124 B.n1123 585
R1529 B.n32 B.n31 585
R1530 B.n1122 B.n32 585
R1531 B.n1120 B.n1119 585
R1532 B.n1121 B.n1120 585
R1533 B.n1118 B.n37 585
R1534 B.n37 B.n36 585
R1535 B.n1117 B.n1116 585
R1536 B.n1116 B.n1115 585
R1537 B.n39 B.n38 585
R1538 B.n1114 B.n39 585
R1539 B.n1112 B.n1111 585
R1540 B.n1113 B.n1112 585
R1541 B.n1110 B.n44 585
R1542 B.n44 B.n43 585
R1543 B.n1109 B.n1108 585
R1544 B.n1108 B.n1107 585
R1545 B.n46 B.n45 585
R1546 B.n1106 B.n46 585
R1547 B.n1104 B.n1103 585
R1548 B.n1105 B.n1104 585
R1549 B.n1102 B.n51 585
R1550 B.n51 B.n50 585
R1551 B.n1101 B.n1100 585
R1552 B.n1100 B.n1099 585
R1553 B.n53 B.n52 585
R1554 B.n1098 B.n53 585
R1555 B.n1096 B.n1095 585
R1556 B.n1097 B.n1096 585
R1557 B.n1094 B.n58 585
R1558 B.n58 B.n57 585
R1559 B.n1093 B.n1092 585
R1560 B.n1092 B.n1091 585
R1561 B.n60 B.n59 585
R1562 B.n1090 B.n60 585
R1563 B.n1088 B.n1087 585
R1564 B.n1089 B.n1088 585
R1565 B.n1086 B.n65 585
R1566 B.n65 B.n64 585
R1567 B.n1085 B.n1084 585
R1568 B.n1084 B.n1083 585
R1569 B.n67 B.n66 585
R1570 B.n1082 B.n67 585
R1571 B.n1080 B.n1079 585
R1572 B.n1081 B.n1080 585
R1573 B.n1078 B.n72 585
R1574 B.n72 B.n71 585
R1575 B.n1077 B.n1076 585
R1576 B.n1076 B.n1075 585
R1577 B.n74 B.n73 585
R1578 B.n1074 B.n74 585
R1579 B.n1072 B.n1071 585
R1580 B.n1073 B.n1072 585
R1581 B.n1070 B.n79 585
R1582 B.n79 B.n78 585
R1583 B.n1069 B.n1068 585
R1584 B.n1068 B.n1067 585
R1585 B.n81 B.n80 585
R1586 B.n1066 B.n81 585
R1587 B.n1064 B.n1063 585
R1588 B.n1065 B.n1064 585
R1589 B.n1062 B.n86 585
R1590 B.n86 B.n85 585
R1591 B.n1061 B.n1060 585
R1592 B.n1060 B.n1059 585
R1593 B.n88 B.n87 585
R1594 B.n1058 B.n88 585
R1595 B.n1056 B.n1055 585
R1596 B.n1057 B.n1056 585
R1597 B.n1054 B.n93 585
R1598 B.n93 B.n92 585
R1599 B.n1053 B.n1052 585
R1600 B.n1052 B.n1051 585
R1601 B.n95 B.n94 585
R1602 B.n1050 B.n95 585
R1603 B.n1048 B.n1047 585
R1604 B.n1049 B.n1048 585
R1605 B.n1046 B.n100 585
R1606 B.n100 B.n99 585
R1607 B.n1045 B.n1044 585
R1608 B.n1044 B.n1043 585
R1609 B.n102 B.n101 585
R1610 B.n1042 B.n102 585
R1611 B.n1040 B.n1039 585
R1612 B.n1041 B.n1040 585
R1613 B.n1038 B.n107 585
R1614 B.n107 B.n106 585
R1615 B.n1037 B.n1036 585
R1616 B.n1036 B.n1035 585
R1617 B.n109 B.n108 585
R1618 B.n1034 B.n109 585
R1619 B.n1032 B.n1031 585
R1620 B.n1033 B.n1032 585
R1621 B.n1030 B.n114 585
R1622 B.n114 B.n113 585
R1623 B.n1029 B.n1028 585
R1624 B.n1028 B.n1027 585
R1625 B.n116 B.n115 585
R1626 B.n1026 B.n116 585
R1627 B.n1024 B.n1023 585
R1628 B.n1025 B.n1024 585
R1629 B.n1022 B.n121 585
R1630 B.n121 B.n120 585
R1631 B.n1021 B.n1020 585
R1632 B.n1020 B.n1019 585
R1633 B.n123 B.n122 585
R1634 B.n1018 B.n123 585
R1635 B.n1157 B.n1156 585
R1636 B.n1156 B.n1155 585
R1637 B.n716 B.n487 458.866
R1638 B.n177 B.n123 458.866
R1639 B.n719 B.n489 458.866
R1640 B.n1015 B.n125 458.866
R1641 B.n539 B.t14 352.913
R1642 B.n171 B.t17 352.913
R1643 B.n537 B.t11 352.913
R1644 B.n174 B.t20 352.913
R1645 B.n539 B.t12 281.714
R1646 B.n537 B.t8 281.714
R1647 B.n174 B.t19 281.714
R1648 B.n171 B.t15 281.714
R1649 B.n540 B.t13 272.623
R1650 B.n172 B.t18 272.623
R1651 B.n538 B.t10 272.623
R1652 B.n175 B.t21 272.623
R1653 B.n1017 B.n1016 256.663
R1654 B.n1017 B.n169 256.663
R1655 B.n1017 B.n168 256.663
R1656 B.n1017 B.n167 256.663
R1657 B.n1017 B.n166 256.663
R1658 B.n1017 B.n165 256.663
R1659 B.n1017 B.n164 256.663
R1660 B.n1017 B.n163 256.663
R1661 B.n1017 B.n162 256.663
R1662 B.n1017 B.n161 256.663
R1663 B.n1017 B.n160 256.663
R1664 B.n1017 B.n159 256.663
R1665 B.n1017 B.n158 256.663
R1666 B.n1017 B.n157 256.663
R1667 B.n1017 B.n156 256.663
R1668 B.n1017 B.n155 256.663
R1669 B.n1017 B.n154 256.663
R1670 B.n1017 B.n153 256.663
R1671 B.n1017 B.n152 256.663
R1672 B.n1017 B.n151 256.663
R1673 B.n1017 B.n150 256.663
R1674 B.n1017 B.n149 256.663
R1675 B.n1017 B.n148 256.663
R1676 B.n1017 B.n147 256.663
R1677 B.n1017 B.n146 256.663
R1678 B.n1017 B.n145 256.663
R1679 B.n1017 B.n144 256.663
R1680 B.n1017 B.n143 256.663
R1681 B.n1017 B.n142 256.663
R1682 B.n1017 B.n141 256.663
R1683 B.n1017 B.n140 256.663
R1684 B.n1017 B.n139 256.663
R1685 B.n1017 B.n138 256.663
R1686 B.n1017 B.n137 256.663
R1687 B.n1017 B.n136 256.663
R1688 B.n1017 B.n135 256.663
R1689 B.n1017 B.n134 256.663
R1690 B.n1017 B.n133 256.663
R1691 B.n1017 B.n132 256.663
R1692 B.n1017 B.n131 256.663
R1693 B.n1017 B.n130 256.663
R1694 B.n1017 B.n129 256.663
R1695 B.n1017 B.n128 256.663
R1696 B.n1017 B.n127 256.663
R1697 B.n1017 B.n126 256.663
R1698 B.n718 B.n717 256.663
R1699 B.n718 B.n492 256.663
R1700 B.n718 B.n493 256.663
R1701 B.n718 B.n494 256.663
R1702 B.n718 B.n495 256.663
R1703 B.n718 B.n496 256.663
R1704 B.n718 B.n497 256.663
R1705 B.n718 B.n498 256.663
R1706 B.n718 B.n499 256.663
R1707 B.n718 B.n500 256.663
R1708 B.n718 B.n501 256.663
R1709 B.n718 B.n502 256.663
R1710 B.n718 B.n503 256.663
R1711 B.n718 B.n504 256.663
R1712 B.n718 B.n505 256.663
R1713 B.n718 B.n506 256.663
R1714 B.n718 B.n507 256.663
R1715 B.n718 B.n508 256.663
R1716 B.n718 B.n509 256.663
R1717 B.n718 B.n510 256.663
R1718 B.n718 B.n511 256.663
R1719 B.n718 B.n512 256.663
R1720 B.n718 B.n513 256.663
R1721 B.n718 B.n514 256.663
R1722 B.n718 B.n515 256.663
R1723 B.n718 B.n516 256.663
R1724 B.n718 B.n517 256.663
R1725 B.n718 B.n518 256.663
R1726 B.n718 B.n519 256.663
R1727 B.n718 B.n520 256.663
R1728 B.n718 B.n521 256.663
R1729 B.n718 B.n522 256.663
R1730 B.n718 B.n523 256.663
R1731 B.n718 B.n524 256.663
R1732 B.n718 B.n525 256.663
R1733 B.n718 B.n526 256.663
R1734 B.n718 B.n527 256.663
R1735 B.n718 B.n528 256.663
R1736 B.n718 B.n529 256.663
R1737 B.n718 B.n530 256.663
R1738 B.n718 B.n531 256.663
R1739 B.n718 B.n532 256.663
R1740 B.n718 B.n533 256.663
R1741 B.n718 B.n534 256.663
R1742 B.n725 B.n487 163.367
R1743 B.n725 B.n485 163.367
R1744 B.n729 B.n485 163.367
R1745 B.n729 B.n479 163.367
R1746 B.n737 B.n479 163.367
R1747 B.n737 B.n477 163.367
R1748 B.n741 B.n477 163.367
R1749 B.n741 B.n471 163.367
R1750 B.n749 B.n471 163.367
R1751 B.n749 B.n469 163.367
R1752 B.n753 B.n469 163.367
R1753 B.n753 B.n463 163.367
R1754 B.n761 B.n463 163.367
R1755 B.n761 B.n461 163.367
R1756 B.n765 B.n461 163.367
R1757 B.n765 B.n455 163.367
R1758 B.n773 B.n455 163.367
R1759 B.n773 B.n453 163.367
R1760 B.n777 B.n453 163.367
R1761 B.n777 B.n447 163.367
R1762 B.n785 B.n447 163.367
R1763 B.n785 B.n445 163.367
R1764 B.n789 B.n445 163.367
R1765 B.n789 B.n439 163.367
R1766 B.n797 B.n439 163.367
R1767 B.n797 B.n437 163.367
R1768 B.n801 B.n437 163.367
R1769 B.n801 B.n431 163.367
R1770 B.n809 B.n431 163.367
R1771 B.n809 B.n429 163.367
R1772 B.n813 B.n429 163.367
R1773 B.n813 B.n423 163.367
R1774 B.n821 B.n423 163.367
R1775 B.n821 B.n421 163.367
R1776 B.n825 B.n421 163.367
R1777 B.n825 B.n415 163.367
R1778 B.n833 B.n415 163.367
R1779 B.n833 B.n413 163.367
R1780 B.n837 B.n413 163.367
R1781 B.n837 B.n407 163.367
R1782 B.n845 B.n407 163.367
R1783 B.n845 B.n405 163.367
R1784 B.n849 B.n405 163.367
R1785 B.n849 B.n399 163.367
R1786 B.n857 B.n399 163.367
R1787 B.n857 B.n397 163.367
R1788 B.n861 B.n397 163.367
R1789 B.n861 B.n391 163.367
R1790 B.n869 B.n391 163.367
R1791 B.n869 B.n389 163.367
R1792 B.n873 B.n389 163.367
R1793 B.n873 B.n383 163.367
R1794 B.n881 B.n383 163.367
R1795 B.n881 B.n381 163.367
R1796 B.n885 B.n381 163.367
R1797 B.n885 B.n375 163.367
R1798 B.n893 B.n375 163.367
R1799 B.n893 B.n373 163.367
R1800 B.n897 B.n373 163.367
R1801 B.n897 B.n367 163.367
R1802 B.n905 B.n367 163.367
R1803 B.n905 B.n365 163.367
R1804 B.n909 B.n365 163.367
R1805 B.n909 B.n359 163.367
R1806 B.n918 B.n359 163.367
R1807 B.n918 B.n357 163.367
R1808 B.n922 B.n357 163.367
R1809 B.n922 B.n2 163.367
R1810 B.n1156 B.n2 163.367
R1811 B.n1156 B.n3 163.367
R1812 B.n1152 B.n3 163.367
R1813 B.n1152 B.n9 163.367
R1814 B.n1148 B.n9 163.367
R1815 B.n1148 B.n11 163.367
R1816 B.n1144 B.n11 163.367
R1817 B.n1144 B.n16 163.367
R1818 B.n1140 B.n16 163.367
R1819 B.n1140 B.n18 163.367
R1820 B.n1136 B.n18 163.367
R1821 B.n1136 B.n23 163.367
R1822 B.n1132 B.n23 163.367
R1823 B.n1132 B.n25 163.367
R1824 B.n1128 B.n25 163.367
R1825 B.n1128 B.n30 163.367
R1826 B.n1124 B.n30 163.367
R1827 B.n1124 B.n32 163.367
R1828 B.n1120 B.n32 163.367
R1829 B.n1120 B.n37 163.367
R1830 B.n1116 B.n37 163.367
R1831 B.n1116 B.n39 163.367
R1832 B.n1112 B.n39 163.367
R1833 B.n1112 B.n44 163.367
R1834 B.n1108 B.n44 163.367
R1835 B.n1108 B.n46 163.367
R1836 B.n1104 B.n46 163.367
R1837 B.n1104 B.n51 163.367
R1838 B.n1100 B.n51 163.367
R1839 B.n1100 B.n53 163.367
R1840 B.n1096 B.n53 163.367
R1841 B.n1096 B.n58 163.367
R1842 B.n1092 B.n58 163.367
R1843 B.n1092 B.n60 163.367
R1844 B.n1088 B.n60 163.367
R1845 B.n1088 B.n65 163.367
R1846 B.n1084 B.n65 163.367
R1847 B.n1084 B.n67 163.367
R1848 B.n1080 B.n67 163.367
R1849 B.n1080 B.n72 163.367
R1850 B.n1076 B.n72 163.367
R1851 B.n1076 B.n74 163.367
R1852 B.n1072 B.n74 163.367
R1853 B.n1072 B.n79 163.367
R1854 B.n1068 B.n79 163.367
R1855 B.n1068 B.n81 163.367
R1856 B.n1064 B.n81 163.367
R1857 B.n1064 B.n86 163.367
R1858 B.n1060 B.n86 163.367
R1859 B.n1060 B.n88 163.367
R1860 B.n1056 B.n88 163.367
R1861 B.n1056 B.n93 163.367
R1862 B.n1052 B.n93 163.367
R1863 B.n1052 B.n95 163.367
R1864 B.n1048 B.n95 163.367
R1865 B.n1048 B.n100 163.367
R1866 B.n1044 B.n100 163.367
R1867 B.n1044 B.n102 163.367
R1868 B.n1040 B.n102 163.367
R1869 B.n1040 B.n107 163.367
R1870 B.n1036 B.n107 163.367
R1871 B.n1036 B.n109 163.367
R1872 B.n1032 B.n109 163.367
R1873 B.n1032 B.n114 163.367
R1874 B.n1028 B.n114 163.367
R1875 B.n1028 B.n116 163.367
R1876 B.n1024 B.n116 163.367
R1877 B.n1024 B.n121 163.367
R1878 B.n1020 B.n121 163.367
R1879 B.n1020 B.n123 163.367
R1880 B.n536 B.n535 163.367
R1881 B.n711 B.n535 163.367
R1882 B.n709 B.n708 163.367
R1883 B.n705 B.n704 163.367
R1884 B.n701 B.n700 163.367
R1885 B.n697 B.n696 163.367
R1886 B.n693 B.n692 163.367
R1887 B.n689 B.n688 163.367
R1888 B.n685 B.n684 163.367
R1889 B.n681 B.n680 163.367
R1890 B.n677 B.n676 163.367
R1891 B.n673 B.n672 163.367
R1892 B.n669 B.n668 163.367
R1893 B.n665 B.n664 163.367
R1894 B.n661 B.n660 163.367
R1895 B.n657 B.n656 163.367
R1896 B.n653 B.n652 163.367
R1897 B.n649 B.n648 163.367
R1898 B.n645 B.n644 163.367
R1899 B.n641 B.n640 163.367
R1900 B.n636 B.n635 163.367
R1901 B.n632 B.n631 163.367
R1902 B.n628 B.n627 163.367
R1903 B.n624 B.n623 163.367
R1904 B.n620 B.n619 163.367
R1905 B.n615 B.n614 163.367
R1906 B.n611 B.n610 163.367
R1907 B.n607 B.n606 163.367
R1908 B.n603 B.n602 163.367
R1909 B.n599 B.n598 163.367
R1910 B.n595 B.n594 163.367
R1911 B.n591 B.n590 163.367
R1912 B.n587 B.n586 163.367
R1913 B.n583 B.n582 163.367
R1914 B.n579 B.n578 163.367
R1915 B.n575 B.n574 163.367
R1916 B.n571 B.n570 163.367
R1917 B.n567 B.n566 163.367
R1918 B.n563 B.n562 163.367
R1919 B.n559 B.n558 163.367
R1920 B.n555 B.n554 163.367
R1921 B.n551 B.n550 163.367
R1922 B.n547 B.n546 163.367
R1923 B.n543 B.n542 163.367
R1924 B.n719 B.n491 163.367
R1925 B.n723 B.n489 163.367
R1926 B.n723 B.n483 163.367
R1927 B.n731 B.n483 163.367
R1928 B.n731 B.n481 163.367
R1929 B.n735 B.n481 163.367
R1930 B.n735 B.n475 163.367
R1931 B.n743 B.n475 163.367
R1932 B.n743 B.n473 163.367
R1933 B.n747 B.n473 163.367
R1934 B.n747 B.n467 163.367
R1935 B.n755 B.n467 163.367
R1936 B.n755 B.n465 163.367
R1937 B.n759 B.n465 163.367
R1938 B.n759 B.n459 163.367
R1939 B.n767 B.n459 163.367
R1940 B.n767 B.n457 163.367
R1941 B.n771 B.n457 163.367
R1942 B.n771 B.n451 163.367
R1943 B.n779 B.n451 163.367
R1944 B.n779 B.n449 163.367
R1945 B.n783 B.n449 163.367
R1946 B.n783 B.n442 163.367
R1947 B.n791 B.n442 163.367
R1948 B.n791 B.n440 163.367
R1949 B.n795 B.n440 163.367
R1950 B.n795 B.n435 163.367
R1951 B.n803 B.n435 163.367
R1952 B.n803 B.n433 163.367
R1953 B.n807 B.n433 163.367
R1954 B.n807 B.n427 163.367
R1955 B.n815 B.n427 163.367
R1956 B.n815 B.n425 163.367
R1957 B.n819 B.n425 163.367
R1958 B.n819 B.n418 163.367
R1959 B.n827 B.n418 163.367
R1960 B.n827 B.n416 163.367
R1961 B.n831 B.n416 163.367
R1962 B.n831 B.n411 163.367
R1963 B.n839 B.n411 163.367
R1964 B.n839 B.n409 163.367
R1965 B.n843 B.n409 163.367
R1966 B.n843 B.n403 163.367
R1967 B.n851 B.n403 163.367
R1968 B.n851 B.n401 163.367
R1969 B.n855 B.n401 163.367
R1970 B.n855 B.n395 163.367
R1971 B.n863 B.n395 163.367
R1972 B.n863 B.n393 163.367
R1973 B.n867 B.n393 163.367
R1974 B.n867 B.n387 163.367
R1975 B.n875 B.n387 163.367
R1976 B.n875 B.n385 163.367
R1977 B.n879 B.n385 163.367
R1978 B.n879 B.n379 163.367
R1979 B.n887 B.n379 163.367
R1980 B.n887 B.n377 163.367
R1981 B.n891 B.n377 163.367
R1982 B.n891 B.n371 163.367
R1983 B.n899 B.n371 163.367
R1984 B.n899 B.n369 163.367
R1985 B.n903 B.n369 163.367
R1986 B.n903 B.n363 163.367
R1987 B.n911 B.n363 163.367
R1988 B.n911 B.n361 163.367
R1989 B.n916 B.n361 163.367
R1990 B.n916 B.n355 163.367
R1991 B.n924 B.n355 163.367
R1992 B.n925 B.n924 163.367
R1993 B.n925 B.n5 163.367
R1994 B.n6 B.n5 163.367
R1995 B.n7 B.n6 163.367
R1996 B.n930 B.n7 163.367
R1997 B.n930 B.n12 163.367
R1998 B.n13 B.n12 163.367
R1999 B.n14 B.n13 163.367
R2000 B.n935 B.n14 163.367
R2001 B.n935 B.n19 163.367
R2002 B.n20 B.n19 163.367
R2003 B.n21 B.n20 163.367
R2004 B.n940 B.n21 163.367
R2005 B.n940 B.n26 163.367
R2006 B.n27 B.n26 163.367
R2007 B.n28 B.n27 163.367
R2008 B.n945 B.n28 163.367
R2009 B.n945 B.n33 163.367
R2010 B.n34 B.n33 163.367
R2011 B.n35 B.n34 163.367
R2012 B.n950 B.n35 163.367
R2013 B.n950 B.n40 163.367
R2014 B.n41 B.n40 163.367
R2015 B.n42 B.n41 163.367
R2016 B.n955 B.n42 163.367
R2017 B.n955 B.n47 163.367
R2018 B.n48 B.n47 163.367
R2019 B.n49 B.n48 163.367
R2020 B.n960 B.n49 163.367
R2021 B.n960 B.n54 163.367
R2022 B.n55 B.n54 163.367
R2023 B.n56 B.n55 163.367
R2024 B.n965 B.n56 163.367
R2025 B.n965 B.n61 163.367
R2026 B.n62 B.n61 163.367
R2027 B.n63 B.n62 163.367
R2028 B.n970 B.n63 163.367
R2029 B.n970 B.n68 163.367
R2030 B.n69 B.n68 163.367
R2031 B.n70 B.n69 163.367
R2032 B.n975 B.n70 163.367
R2033 B.n975 B.n75 163.367
R2034 B.n76 B.n75 163.367
R2035 B.n77 B.n76 163.367
R2036 B.n980 B.n77 163.367
R2037 B.n980 B.n82 163.367
R2038 B.n83 B.n82 163.367
R2039 B.n84 B.n83 163.367
R2040 B.n985 B.n84 163.367
R2041 B.n985 B.n89 163.367
R2042 B.n90 B.n89 163.367
R2043 B.n91 B.n90 163.367
R2044 B.n990 B.n91 163.367
R2045 B.n990 B.n96 163.367
R2046 B.n97 B.n96 163.367
R2047 B.n98 B.n97 163.367
R2048 B.n995 B.n98 163.367
R2049 B.n995 B.n103 163.367
R2050 B.n104 B.n103 163.367
R2051 B.n105 B.n104 163.367
R2052 B.n1000 B.n105 163.367
R2053 B.n1000 B.n110 163.367
R2054 B.n111 B.n110 163.367
R2055 B.n112 B.n111 163.367
R2056 B.n1005 B.n112 163.367
R2057 B.n1005 B.n117 163.367
R2058 B.n118 B.n117 163.367
R2059 B.n119 B.n118 163.367
R2060 B.n1010 B.n119 163.367
R2061 B.n1010 B.n124 163.367
R2062 B.n125 B.n124 163.367
R2063 B.n181 B.n180 163.367
R2064 B.n185 B.n184 163.367
R2065 B.n189 B.n188 163.367
R2066 B.n193 B.n192 163.367
R2067 B.n197 B.n196 163.367
R2068 B.n201 B.n200 163.367
R2069 B.n205 B.n204 163.367
R2070 B.n209 B.n208 163.367
R2071 B.n213 B.n212 163.367
R2072 B.n217 B.n216 163.367
R2073 B.n221 B.n220 163.367
R2074 B.n225 B.n224 163.367
R2075 B.n229 B.n228 163.367
R2076 B.n233 B.n232 163.367
R2077 B.n237 B.n236 163.367
R2078 B.n241 B.n240 163.367
R2079 B.n245 B.n244 163.367
R2080 B.n249 B.n248 163.367
R2081 B.n253 B.n252 163.367
R2082 B.n257 B.n256 163.367
R2083 B.n261 B.n260 163.367
R2084 B.n265 B.n264 163.367
R2085 B.n269 B.n268 163.367
R2086 B.n273 B.n272 163.367
R2087 B.n277 B.n276 163.367
R2088 B.n281 B.n280 163.367
R2089 B.n285 B.n284 163.367
R2090 B.n289 B.n288 163.367
R2091 B.n293 B.n292 163.367
R2092 B.n297 B.n296 163.367
R2093 B.n301 B.n300 163.367
R2094 B.n305 B.n304 163.367
R2095 B.n309 B.n308 163.367
R2096 B.n313 B.n312 163.367
R2097 B.n317 B.n316 163.367
R2098 B.n321 B.n320 163.367
R2099 B.n325 B.n324 163.367
R2100 B.n329 B.n328 163.367
R2101 B.n333 B.n332 163.367
R2102 B.n337 B.n336 163.367
R2103 B.n341 B.n340 163.367
R2104 B.n345 B.n344 163.367
R2105 B.n349 B.n348 163.367
R2106 B.n351 B.n170 163.367
R2107 B.n718 B.n488 80.9458
R2108 B.n1018 B.n1017 80.9458
R2109 B.n540 B.n539 80.2914
R2110 B.n538 B.n537 80.2914
R2111 B.n175 B.n174 80.2914
R2112 B.n172 B.n171 80.2914
R2113 B.n717 B.n716 71.676
R2114 B.n711 B.n492 71.676
R2115 B.n708 B.n493 71.676
R2116 B.n704 B.n494 71.676
R2117 B.n700 B.n495 71.676
R2118 B.n696 B.n496 71.676
R2119 B.n692 B.n497 71.676
R2120 B.n688 B.n498 71.676
R2121 B.n684 B.n499 71.676
R2122 B.n680 B.n500 71.676
R2123 B.n676 B.n501 71.676
R2124 B.n672 B.n502 71.676
R2125 B.n668 B.n503 71.676
R2126 B.n664 B.n504 71.676
R2127 B.n660 B.n505 71.676
R2128 B.n656 B.n506 71.676
R2129 B.n652 B.n507 71.676
R2130 B.n648 B.n508 71.676
R2131 B.n644 B.n509 71.676
R2132 B.n640 B.n510 71.676
R2133 B.n635 B.n511 71.676
R2134 B.n631 B.n512 71.676
R2135 B.n627 B.n513 71.676
R2136 B.n623 B.n514 71.676
R2137 B.n619 B.n515 71.676
R2138 B.n614 B.n516 71.676
R2139 B.n610 B.n517 71.676
R2140 B.n606 B.n518 71.676
R2141 B.n602 B.n519 71.676
R2142 B.n598 B.n520 71.676
R2143 B.n594 B.n521 71.676
R2144 B.n590 B.n522 71.676
R2145 B.n586 B.n523 71.676
R2146 B.n582 B.n524 71.676
R2147 B.n578 B.n525 71.676
R2148 B.n574 B.n526 71.676
R2149 B.n570 B.n527 71.676
R2150 B.n566 B.n528 71.676
R2151 B.n562 B.n529 71.676
R2152 B.n558 B.n530 71.676
R2153 B.n554 B.n531 71.676
R2154 B.n550 B.n532 71.676
R2155 B.n546 B.n533 71.676
R2156 B.n542 B.n534 71.676
R2157 B.n177 B.n126 71.676
R2158 B.n181 B.n127 71.676
R2159 B.n185 B.n128 71.676
R2160 B.n189 B.n129 71.676
R2161 B.n193 B.n130 71.676
R2162 B.n197 B.n131 71.676
R2163 B.n201 B.n132 71.676
R2164 B.n205 B.n133 71.676
R2165 B.n209 B.n134 71.676
R2166 B.n213 B.n135 71.676
R2167 B.n217 B.n136 71.676
R2168 B.n221 B.n137 71.676
R2169 B.n225 B.n138 71.676
R2170 B.n229 B.n139 71.676
R2171 B.n233 B.n140 71.676
R2172 B.n237 B.n141 71.676
R2173 B.n241 B.n142 71.676
R2174 B.n245 B.n143 71.676
R2175 B.n249 B.n144 71.676
R2176 B.n253 B.n145 71.676
R2177 B.n257 B.n146 71.676
R2178 B.n261 B.n147 71.676
R2179 B.n265 B.n148 71.676
R2180 B.n269 B.n149 71.676
R2181 B.n273 B.n150 71.676
R2182 B.n277 B.n151 71.676
R2183 B.n281 B.n152 71.676
R2184 B.n285 B.n153 71.676
R2185 B.n289 B.n154 71.676
R2186 B.n293 B.n155 71.676
R2187 B.n297 B.n156 71.676
R2188 B.n301 B.n157 71.676
R2189 B.n305 B.n158 71.676
R2190 B.n309 B.n159 71.676
R2191 B.n313 B.n160 71.676
R2192 B.n317 B.n161 71.676
R2193 B.n321 B.n162 71.676
R2194 B.n325 B.n163 71.676
R2195 B.n329 B.n164 71.676
R2196 B.n333 B.n165 71.676
R2197 B.n337 B.n166 71.676
R2198 B.n341 B.n167 71.676
R2199 B.n345 B.n168 71.676
R2200 B.n349 B.n169 71.676
R2201 B.n1016 B.n170 71.676
R2202 B.n1016 B.n1015 71.676
R2203 B.n351 B.n169 71.676
R2204 B.n348 B.n168 71.676
R2205 B.n344 B.n167 71.676
R2206 B.n340 B.n166 71.676
R2207 B.n336 B.n165 71.676
R2208 B.n332 B.n164 71.676
R2209 B.n328 B.n163 71.676
R2210 B.n324 B.n162 71.676
R2211 B.n320 B.n161 71.676
R2212 B.n316 B.n160 71.676
R2213 B.n312 B.n159 71.676
R2214 B.n308 B.n158 71.676
R2215 B.n304 B.n157 71.676
R2216 B.n300 B.n156 71.676
R2217 B.n296 B.n155 71.676
R2218 B.n292 B.n154 71.676
R2219 B.n288 B.n153 71.676
R2220 B.n284 B.n152 71.676
R2221 B.n280 B.n151 71.676
R2222 B.n276 B.n150 71.676
R2223 B.n272 B.n149 71.676
R2224 B.n268 B.n148 71.676
R2225 B.n264 B.n147 71.676
R2226 B.n260 B.n146 71.676
R2227 B.n256 B.n145 71.676
R2228 B.n252 B.n144 71.676
R2229 B.n248 B.n143 71.676
R2230 B.n244 B.n142 71.676
R2231 B.n240 B.n141 71.676
R2232 B.n236 B.n140 71.676
R2233 B.n232 B.n139 71.676
R2234 B.n228 B.n138 71.676
R2235 B.n224 B.n137 71.676
R2236 B.n220 B.n136 71.676
R2237 B.n216 B.n135 71.676
R2238 B.n212 B.n134 71.676
R2239 B.n208 B.n133 71.676
R2240 B.n204 B.n132 71.676
R2241 B.n200 B.n131 71.676
R2242 B.n196 B.n130 71.676
R2243 B.n192 B.n129 71.676
R2244 B.n188 B.n128 71.676
R2245 B.n184 B.n127 71.676
R2246 B.n180 B.n126 71.676
R2247 B.n717 B.n536 71.676
R2248 B.n709 B.n492 71.676
R2249 B.n705 B.n493 71.676
R2250 B.n701 B.n494 71.676
R2251 B.n697 B.n495 71.676
R2252 B.n693 B.n496 71.676
R2253 B.n689 B.n497 71.676
R2254 B.n685 B.n498 71.676
R2255 B.n681 B.n499 71.676
R2256 B.n677 B.n500 71.676
R2257 B.n673 B.n501 71.676
R2258 B.n669 B.n502 71.676
R2259 B.n665 B.n503 71.676
R2260 B.n661 B.n504 71.676
R2261 B.n657 B.n505 71.676
R2262 B.n653 B.n506 71.676
R2263 B.n649 B.n507 71.676
R2264 B.n645 B.n508 71.676
R2265 B.n641 B.n509 71.676
R2266 B.n636 B.n510 71.676
R2267 B.n632 B.n511 71.676
R2268 B.n628 B.n512 71.676
R2269 B.n624 B.n513 71.676
R2270 B.n620 B.n514 71.676
R2271 B.n615 B.n515 71.676
R2272 B.n611 B.n516 71.676
R2273 B.n607 B.n517 71.676
R2274 B.n603 B.n518 71.676
R2275 B.n599 B.n519 71.676
R2276 B.n595 B.n520 71.676
R2277 B.n591 B.n521 71.676
R2278 B.n587 B.n522 71.676
R2279 B.n583 B.n523 71.676
R2280 B.n579 B.n524 71.676
R2281 B.n575 B.n525 71.676
R2282 B.n571 B.n526 71.676
R2283 B.n567 B.n527 71.676
R2284 B.n563 B.n528 71.676
R2285 B.n559 B.n529 71.676
R2286 B.n555 B.n530 71.676
R2287 B.n551 B.n531 71.676
R2288 B.n547 B.n532 71.676
R2289 B.n543 B.n533 71.676
R2290 B.n534 B.n491 71.676
R2291 B.n617 B.n540 59.5399
R2292 B.n638 B.n538 59.5399
R2293 B.n176 B.n175 59.5399
R2294 B.n173 B.n172 59.5399
R2295 B.n724 B.n488 44.7507
R2296 B.n724 B.n484 44.7507
R2297 B.n730 B.n484 44.7507
R2298 B.n730 B.n480 44.7507
R2299 B.n736 B.n480 44.7507
R2300 B.n736 B.n476 44.7507
R2301 B.n742 B.n476 44.7507
R2302 B.n742 B.n472 44.7507
R2303 B.n748 B.n472 44.7507
R2304 B.n754 B.n468 44.7507
R2305 B.n754 B.n464 44.7507
R2306 B.n760 B.n464 44.7507
R2307 B.n760 B.n460 44.7507
R2308 B.n766 B.n460 44.7507
R2309 B.n766 B.n456 44.7507
R2310 B.n772 B.n456 44.7507
R2311 B.n772 B.n452 44.7507
R2312 B.n778 B.n452 44.7507
R2313 B.n778 B.n448 44.7507
R2314 B.n784 B.n448 44.7507
R2315 B.n784 B.n443 44.7507
R2316 B.n790 B.n443 44.7507
R2317 B.n790 B.n444 44.7507
R2318 B.n796 B.n436 44.7507
R2319 B.n802 B.n436 44.7507
R2320 B.n802 B.n432 44.7507
R2321 B.n808 B.n432 44.7507
R2322 B.n808 B.n428 44.7507
R2323 B.n814 B.n428 44.7507
R2324 B.n814 B.n424 44.7507
R2325 B.n820 B.n424 44.7507
R2326 B.n820 B.n419 44.7507
R2327 B.n826 B.n419 44.7507
R2328 B.n826 B.n420 44.7507
R2329 B.n832 B.n412 44.7507
R2330 B.n838 B.n412 44.7507
R2331 B.n838 B.n408 44.7507
R2332 B.n844 B.n408 44.7507
R2333 B.n844 B.n404 44.7507
R2334 B.n850 B.n404 44.7507
R2335 B.n850 B.n400 44.7507
R2336 B.n856 B.n400 44.7507
R2337 B.n856 B.n396 44.7507
R2338 B.n862 B.n396 44.7507
R2339 B.n862 B.n392 44.7507
R2340 B.n868 B.n392 44.7507
R2341 B.n874 B.n388 44.7507
R2342 B.n874 B.n384 44.7507
R2343 B.n880 B.n384 44.7507
R2344 B.n880 B.n380 44.7507
R2345 B.n886 B.n380 44.7507
R2346 B.n886 B.n376 44.7507
R2347 B.n892 B.n376 44.7507
R2348 B.n892 B.n372 44.7507
R2349 B.n898 B.n372 44.7507
R2350 B.n898 B.n368 44.7507
R2351 B.n904 B.n368 44.7507
R2352 B.n910 B.n364 44.7507
R2353 B.n910 B.n360 44.7507
R2354 B.n917 B.n360 44.7507
R2355 B.n917 B.n356 44.7507
R2356 B.n923 B.n356 44.7507
R2357 B.n923 B.n4 44.7507
R2358 B.n1155 B.n4 44.7507
R2359 B.n1155 B.n1154 44.7507
R2360 B.n1154 B.n1153 44.7507
R2361 B.n1153 B.n8 44.7507
R2362 B.n1147 B.n8 44.7507
R2363 B.n1147 B.n1146 44.7507
R2364 B.n1146 B.n1145 44.7507
R2365 B.n1145 B.n15 44.7507
R2366 B.n1139 B.n1138 44.7507
R2367 B.n1138 B.n1137 44.7507
R2368 B.n1137 B.n22 44.7507
R2369 B.n1131 B.n22 44.7507
R2370 B.n1131 B.n1130 44.7507
R2371 B.n1130 B.n1129 44.7507
R2372 B.n1129 B.n29 44.7507
R2373 B.n1123 B.n29 44.7507
R2374 B.n1123 B.n1122 44.7507
R2375 B.n1122 B.n1121 44.7507
R2376 B.n1121 B.n36 44.7507
R2377 B.n1115 B.n1114 44.7507
R2378 B.n1114 B.n1113 44.7507
R2379 B.n1113 B.n43 44.7507
R2380 B.n1107 B.n43 44.7507
R2381 B.n1107 B.n1106 44.7507
R2382 B.n1106 B.n1105 44.7507
R2383 B.n1105 B.n50 44.7507
R2384 B.n1099 B.n50 44.7507
R2385 B.n1099 B.n1098 44.7507
R2386 B.n1098 B.n1097 44.7507
R2387 B.n1097 B.n57 44.7507
R2388 B.n1091 B.n57 44.7507
R2389 B.n1090 B.n1089 44.7507
R2390 B.n1089 B.n64 44.7507
R2391 B.n1083 B.n64 44.7507
R2392 B.n1083 B.n1082 44.7507
R2393 B.n1082 B.n1081 44.7507
R2394 B.n1081 B.n71 44.7507
R2395 B.n1075 B.n71 44.7507
R2396 B.n1075 B.n1074 44.7507
R2397 B.n1074 B.n1073 44.7507
R2398 B.n1073 B.n78 44.7507
R2399 B.n1067 B.n78 44.7507
R2400 B.n1066 B.n1065 44.7507
R2401 B.n1065 B.n85 44.7507
R2402 B.n1059 B.n85 44.7507
R2403 B.n1059 B.n1058 44.7507
R2404 B.n1058 B.n1057 44.7507
R2405 B.n1057 B.n92 44.7507
R2406 B.n1051 B.n92 44.7507
R2407 B.n1051 B.n1050 44.7507
R2408 B.n1050 B.n1049 44.7507
R2409 B.n1049 B.n99 44.7507
R2410 B.n1043 B.n99 44.7507
R2411 B.n1043 B.n1042 44.7507
R2412 B.n1042 B.n1041 44.7507
R2413 B.n1041 B.n106 44.7507
R2414 B.n1035 B.n1034 44.7507
R2415 B.n1034 B.n1033 44.7507
R2416 B.n1033 B.n113 44.7507
R2417 B.n1027 B.n113 44.7507
R2418 B.n1027 B.n1026 44.7507
R2419 B.n1026 B.n1025 44.7507
R2420 B.n1025 B.n120 44.7507
R2421 B.n1019 B.n120 44.7507
R2422 B.n1019 B.n1018 44.7507
R2423 B.n420 B.t5 42.7764
R2424 B.t4 B.n1090 42.7764
R2425 B.t1 B.n388 38.8279
R2426 B.t6 B.n36 38.8279
R2427 B.n444 B.t7 34.8794
R2428 B.t3 B.n1066 34.8794
R2429 B.t2 B.n364 30.9308
R2430 B.t0 B.n15 30.9308
R2431 B.n1014 B.n1013 29.8151
R2432 B.n178 B.n122 29.8151
R2433 B.n721 B.n720 29.8151
R2434 B.n715 B.n486 29.8151
R2435 B.t9 B.n468 26.9823
R2436 B.t16 B.n106 26.9823
R2437 B B.n1157 18.0485
R2438 B.n748 B.t9 17.769
R2439 B.n1035 B.t16 17.769
R2440 B.n904 B.t2 13.8204
R2441 B.n1139 B.t0 13.8204
R2442 B.n179 B.n178 10.6151
R2443 B.n182 B.n179 10.6151
R2444 B.n183 B.n182 10.6151
R2445 B.n186 B.n183 10.6151
R2446 B.n187 B.n186 10.6151
R2447 B.n190 B.n187 10.6151
R2448 B.n191 B.n190 10.6151
R2449 B.n194 B.n191 10.6151
R2450 B.n195 B.n194 10.6151
R2451 B.n198 B.n195 10.6151
R2452 B.n199 B.n198 10.6151
R2453 B.n202 B.n199 10.6151
R2454 B.n203 B.n202 10.6151
R2455 B.n206 B.n203 10.6151
R2456 B.n207 B.n206 10.6151
R2457 B.n210 B.n207 10.6151
R2458 B.n211 B.n210 10.6151
R2459 B.n214 B.n211 10.6151
R2460 B.n215 B.n214 10.6151
R2461 B.n218 B.n215 10.6151
R2462 B.n219 B.n218 10.6151
R2463 B.n222 B.n219 10.6151
R2464 B.n223 B.n222 10.6151
R2465 B.n226 B.n223 10.6151
R2466 B.n227 B.n226 10.6151
R2467 B.n230 B.n227 10.6151
R2468 B.n231 B.n230 10.6151
R2469 B.n234 B.n231 10.6151
R2470 B.n235 B.n234 10.6151
R2471 B.n238 B.n235 10.6151
R2472 B.n239 B.n238 10.6151
R2473 B.n242 B.n239 10.6151
R2474 B.n243 B.n242 10.6151
R2475 B.n246 B.n243 10.6151
R2476 B.n247 B.n246 10.6151
R2477 B.n250 B.n247 10.6151
R2478 B.n251 B.n250 10.6151
R2479 B.n254 B.n251 10.6151
R2480 B.n255 B.n254 10.6151
R2481 B.n259 B.n258 10.6151
R2482 B.n262 B.n259 10.6151
R2483 B.n263 B.n262 10.6151
R2484 B.n266 B.n263 10.6151
R2485 B.n267 B.n266 10.6151
R2486 B.n270 B.n267 10.6151
R2487 B.n271 B.n270 10.6151
R2488 B.n274 B.n271 10.6151
R2489 B.n275 B.n274 10.6151
R2490 B.n279 B.n278 10.6151
R2491 B.n282 B.n279 10.6151
R2492 B.n283 B.n282 10.6151
R2493 B.n286 B.n283 10.6151
R2494 B.n287 B.n286 10.6151
R2495 B.n290 B.n287 10.6151
R2496 B.n291 B.n290 10.6151
R2497 B.n294 B.n291 10.6151
R2498 B.n295 B.n294 10.6151
R2499 B.n298 B.n295 10.6151
R2500 B.n299 B.n298 10.6151
R2501 B.n302 B.n299 10.6151
R2502 B.n303 B.n302 10.6151
R2503 B.n306 B.n303 10.6151
R2504 B.n307 B.n306 10.6151
R2505 B.n310 B.n307 10.6151
R2506 B.n311 B.n310 10.6151
R2507 B.n314 B.n311 10.6151
R2508 B.n315 B.n314 10.6151
R2509 B.n318 B.n315 10.6151
R2510 B.n319 B.n318 10.6151
R2511 B.n322 B.n319 10.6151
R2512 B.n323 B.n322 10.6151
R2513 B.n326 B.n323 10.6151
R2514 B.n327 B.n326 10.6151
R2515 B.n330 B.n327 10.6151
R2516 B.n331 B.n330 10.6151
R2517 B.n334 B.n331 10.6151
R2518 B.n335 B.n334 10.6151
R2519 B.n338 B.n335 10.6151
R2520 B.n339 B.n338 10.6151
R2521 B.n342 B.n339 10.6151
R2522 B.n343 B.n342 10.6151
R2523 B.n346 B.n343 10.6151
R2524 B.n347 B.n346 10.6151
R2525 B.n350 B.n347 10.6151
R2526 B.n352 B.n350 10.6151
R2527 B.n353 B.n352 10.6151
R2528 B.n1014 B.n353 10.6151
R2529 B.n722 B.n721 10.6151
R2530 B.n722 B.n482 10.6151
R2531 B.n732 B.n482 10.6151
R2532 B.n733 B.n732 10.6151
R2533 B.n734 B.n733 10.6151
R2534 B.n734 B.n474 10.6151
R2535 B.n744 B.n474 10.6151
R2536 B.n745 B.n744 10.6151
R2537 B.n746 B.n745 10.6151
R2538 B.n746 B.n466 10.6151
R2539 B.n756 B.n466 10.6151
R2540 B.n757 B.n756 10.6151
R2541 B.n758 B.n757 10.6151
R2542 B.n758 B.n458 10.6151
R2543 B.n768 B.n458 10.6151
R2544 B.n769 B.n768 10.6151
R2545 B.n770 B.n769 10.6151
R2546 B.n770 B.n450 10.6151
R2547 B.n780 B.n450 10.6151
R2548 B.n781 B.n780 10.6151
R2549 B.n782 B.n781 10.6151
R2550 B.n782 B.n441 10.6151
R2551 B.n792 B.n441 10.6151
R2552 B.n793 B.n792 10.6151
R2553 B.n794 B.n793 10.6151
R2554 B.n794 B.n434 10.6151
R2555 B.n804 B.n434 10.6151
R2556 B.n805 B.n804 10.6151
R2557 B.n806 B.n805 10.6151
R2558 B.n806 B.n426 10.6151
R2559 B.n816 B.n426 10.6151
R2560 B.n817 B.n816 10.6151
R2561 B.n818 B.n817 10.6151
R2562 B.n818 B.n417 10.6151
R2563 B.n828 B.n417 10.6151
R2564 B.n829 B.n828 10.6151
R2565 B.n830 B.n829 10.6151
R2566 B.n830 B.n410 10.6151
R2567 B.n840 B.n410 10.6151
R2568 B.n841 B.n840 10.6151
R2569 B.n842 B.n841 10.6151
R2570 B.n842 B.n402 10.6151
R2571 B.n852 B.n402 10.6151
R2572 B.n853 B.n852 10.6151
R2573 B.n854 B.n853 10.6151
R2574 B.n854 B.n394 10.6151
R2575 B.n864 B.n394 10.6151
R2576 B.n865 B.n864 10.6151
R2577 B.n866 B.n865 10.6151
R2578 B.n866 B.n386 10.6151
R2579 B.n876 B.n386 10.6151
R2580 B.n877 B.n876 10.6151
R2581 B.n878 B.n877 10.6151
R2582 B.n878 B.n378 10.6151
R2583 B.n888 B.n378 10.6151
R2584 B.n889 B.n888 10.6151
R2585 B.n890 B.n889 10.6151
R2586 B.n890 B.n370 10.6151
R2587 B.n900 B.n370 10.6151
R2588 B.n901 B.n900 10.6151
R2589 B.n902 B.n901 10.6151
R2590 B.n902 B.n362 10.6151
R2591 B.n912 B.n362 10.6151
R2592 B.n913 B.n912 10.6151
R2593 B.n915 B.n913 10.6151
R2594 B.n915 B.n914 10.6151
R2595 B.n914 B.n354 10.6151
R2596 B.n926 B.n354 10.6151
R2597 B.n927 B.n926 10.6151
R2598 B.n928 B.n927 10.6151
R2599 B.n929 B.n928 10.6151
R2600 B.n931 B.n929 10.6151
R2601 B.n932 B.n931 10.6151
R2602 B.n933 B.n932 10.6151
R2603 B.n934 B.n933 10.6151
R2604 B.n936 B.n934 10.6151
R2605 B.n937 B.n936 10.6151
R2606 B.n938 B.n937 10.6151
R2607 B.n939 B.n938 10.6151
R2608 B.n941 B.n939 10.6151
R2609 B.n942 B.n941 10.6151
R2610 B.n943 B.n942 10.6151
R2611 B.n944 B.n943 10.6151
R2612 B.n946 B.n944 10.6151
R2613 B.n947 B.n946 10.6151
R2614 B.n948 B.n947 10.6151
R2615 B.n949 B.n948 10.6151
R2616 B.n951 B.n949 10.6151
R2617 B.n952 B.n951 10.6151
R2618 B.n953 B.n952 10.6151
R2619 B.n954 B.n953 10.6151
R2620 B.n956 B.n954 10.6151
R2621 B.n957 B.n956 10.6151
R2622 B.n958 B.n957 10.6151
R2623 B.n959 B.n958 10.6151
R2624 B.n961 B.n959 10.6151
R2625 B.n962 B.n961 10.6151
R2626 B.n963 B.n962 10.6151
R2627 B.n964 B.n963 10.6151
R2628 B.n966 B.n964 10.6151
R2629 B.n967 B.n966 10.6151
R2630 B.n968 B.n967 10.6151
R2631 B.n969 B.n968 10.6151
R2632 B.n971 B.n969 10.6151
R2633 B.n972 B.n971 10.6151
R2634 B.n973 B.n972 10.6151
R2635 B.n974 B.n973 10.6151
R2636 B.n976 B.n974 10.6151
R2637 B.n977 B.n976 10.6151
R2638 B.n978 B.n977 10.6151
R2639 B.n979 B.n978 10.6151
R2640 B.n981 B.n979 10.6151
R2641 B.n982 B.n981 10.6151
R2642 B.n983 B.n982 10.6151
R2643 B.n984 B.n983 10.6151
R2644 B.n986 B.n984 10.6151
R2645 B.n987 B.n986 10.6151
R2646 B.n988 B.n987 10.6151
R2647 B.n989 B.n988 10.6151
R2648 B.n991 B.n989 10.6151
R2649 B.n992 B.n991 10.6151
R2650 B.n993 B.n992 10.6151
R2651 B.n994 B.n993 10.6151
R2652 B.n996 B.n994 10.6151
R2653 B.n997 B.n996 10.6151
R2654 B.n998 B.n997 10.6151
R2655 B.n999 B.n998 10.6151
R2656 B.n1001 B.n999 10.6151
R2657 B.n1002 B.n1001 10.6151
R2658 B.n1003 B.n1002 10.6151
R2659 B.n1004 B.n1003 10.6151
R2660 B.n1006 B.n1004 10.6151
R2661 B.n1007 B.n1006 10.6151
R2662 B.n1008 B.n1007 10.6151
R2663 B.n1009 B.n1008 10.6151
R2664 B.n1011 B.n1009 10.6151
R2665 B.n1012 B.n1011 10.6151
R2666 B.n1013 B.n1012 10.6151
R2667 B.n715 B.n714 10.6151
R2668 B.n714 B.n713 10.6151
R2669 B.n713 B.n712 10.6151
R2670 B.n712 B.n710 10.6151
R2671 B.n710 B.n707 10.6151
R2672 B.n707 B.n706 10.6151
R2673 B.n706 B.n703 10.6151
R2674 B.n703 B.n702 10.6151
R2675 B.n702 B.n699 10.6151
R2676 B.n699 B.n698 10.6151
R2677 B.n698 B.n695 10.6151
R2678 B.n695 B.n694 10.6151
R2679 B.n694 B.n691 10.6151
R2680 B.n691 B.n690 10.6151
R2681 B.n690 B.n687 10.6151
R2682 B.n687 B.n686 10.6151
R2683 B.n686 B.n683 10.6151
R2684 B.n683 B.n682 10.6151
R2685 B.n682 B.n679 10.6151
R2686 B.n679 B.n678 10.6151
R2687 B.n678 B.n675 10.6151
R2688 B.n675 B.n674 10.6151
R2689 B.n674 B.n671 10.6151
R2690 B.n671 B.n670 10.6151
R2691 B.n670 B.n667 10.6151
R2692 B.n667 B.n666 10.6151
R2693 B.n666 B.n663 10.6151
R2694 B.n663 B.n662 10.6151
R2695 B.n662 B.n659 10.6151
R2696 B.n659 B.n658 10.6151
R2697 B.n658 B.n655 10.6151
R2698 B.n655 B.n654 10.6151
R2699 B.n654 B.n651 10.6151
R2700 B.n651 B.n650 10.6151
R2701 B.n650 B.n647 10.6151
R2702 B.n647 B.n646 10.6151
R2703 B.n646 B.n643 10.6151
R2704 B.n643 B.n642 10.6151
R2705 B.n642 B.n639 10.6151
R2706 B.n637 B.n634 10.6151
R2707 B.n634 B.n633 10.6151
R2708 B.n633 B.n630 10.6151
R2709 B.n630 B.n629 10.6151
R2710 B.n629 B.n626 10.6151
R2711 B.n626 B.n625 10.6151
R2712 B.n625 B.n622 10.6151
R2713 B.n622 B.n621 10.6151
R2714 B.n621 B.n618 10.6151
R2715 B.n616 B.n613 10.6151
R2716 B.n613 B.n612 10.6151
R2717 B.n612 B.n609 10.6151
R2718 B.n609 B.n608 10.6151
R2719 B.n608 B.n605 10.6151
R2720 B.n605 B.n604 10.6151
R2721 B.n604 B.n601 10.6151
R2722 B.n601 B.n600 10.6151
R2723 B.n600 B.n597 10.6151
R2724 B.n597 B.n596 10.6151
R2725 B.n596 B.n593 10.6151
R2726 B.n593 B.n592 10.6151
R2727 B.n592 B.n589 10.6151
R2728 B.n589 B.n588 10.6151
R2729 B.n588 B.n585 10.6151
R2730 B.n585 B.n584 10.6151
R2731 B.n584 B.n581 10.6151
R2732 B.n581 B.n580 10.6151
R2733 B.n580 B.n577 10.6151
R2734 B.n577 B.n576 10.6151
R2735 B.n576 B.n573 10.6151
R2736 B.n573 B.n572 10.6151
R2737 B.n572 B.n569 10.6151
R2738 B.n569 B.n568 10.6151
R2739 B.n568 B.n565 10.6151
R2740 B.n565 B.n564 10.6151
R2741 B.n564 B.n561 10.6151
R2742 B.n561 B.n560 10.6151
R2743 B.n560 B.n557 10.6151
R2744 B.n557 B.n556 10.6151
R2745 B.n556 B.n553 10.6151
R2746 B.n553 B.n552 10.6151
R2747 B.n552 B.n549 10.6151
R2748 B.n549 B.n548 10.6151
R2749 B.n548 B.n545 10.6151
R2750 B.n545 B.n544 10.6151
R2751 B.n544 B.n541 10.6151
R2752 B.n541 B.n490 10.6151
R2753 B.n720 B.n490 10.6151
R2754 B.n726 B.n486 10.6151
R2755 B.n727 B.n726 10.6151
R2756 B.n728 B.n727 10.6151
R2757 B.n728 B.n478 10.6151
R2758 B.n738 B.n478 10.6151
R2759 B.n739 B.n738 10.6151
R2760 B.n740 B.n739 10.6151
R2761 B.n740 B.n470 10.6151
R2762 B.n750 B.n470 10.6151
R2763 B.n751 B.n750 10.6151
R2764 B.n752 B.n751 10.6151
R2765 B.n752 B.n462 10.6151
R2766 B.n762 B.n462 10.6151
R2767 B.n763 B.n762 10.6151
R2768 B.n764 B.n763 10.6151
R2769 B.n764 B.n454 10.6151
R2770 B.n774 B.n454 10.6151
R2771 B.n775 B.n774 10.6151
R2772 B.n776 B.n775 10.6151
R2773 B.n776 B.n446 10.6151
R2774 B.n786 B.n446 10.6151
R2775 B.n787 B.n786 10.6151
R2776 B.n788 B.n787 10.6151
R2777 B.n788 B.n438 10.6151
R2778 B.n798 B.n438 10.6151
R2779 B.n799 B.n798 10.6151
R2780 B.n800 B.n799 10.6151
R2781 B.n800 B.n430 10.6151
R2782 B.n810 B.n430 10.6151
R2783 B.n811 B.n810 10.6151
R2784 B.n812 B.n811 10.6151
R2785 B.n812 B.n422 10.6151
R2786 B.n822 B.n422 10.6151
R2787 B.n823 B.n822 10.6151
R2788 B.n824 B.n823 10.6151
R2789 B.n824 B.n414 10.6151
R2790 B.n834 B.n414 10.6151
R2791 B.n835 B.n834 10.6151
R2792 B.n836 B.n835 10.6151
R2793 B.n836 B.n406 10.6151
R2794 B.n846 B.n406 10.6151
R2795 B.n847 B.n846 10.6151
R2796 B.n848 B.n847 10.6151
R2797 B.n848 B.n398 10.6151
R2798 B.n858 B.n398 10.6151
R2799 B.n859 B.n858 10.6151
R2800 B.n860 B.n859 10.6151
R2801 B.n860 B.n390 10.6151
R2802 B.n870 B.n390 10.6151
R2803 B.n871 B.n870 10.6151
R2804 B.n872 B.n871 10.6151
R2805 B.n872 B.n382 10.6151
R2806 B.n882 B.n382 10.6151
R2807 B.n883 B.n882 10.6151
R2808 B.n884 B.n883 10.6151
R2809 B.n884 B.n374 10.6151
R2810 B.n894 B.n374 10.6151
R2811 B.n895 B.n894 10.6151
R2812 B.n896 B.n895 10.6151
R2813 B.n896 B.n366 10.6151
R2814 B.n906 B.n366 10.6151
R2815 B.n907 B.n906 10.6151
R2816 B.n908 B.n907 10.6151
R2817 B.n908 B.n358 10.6151
R2818 B.n919 B.n358 10.6151
R2819 B.n920 B.n919 10.6151
R2820 B.n921 B.n920 10.6151
R2821 B.n921 B.n0 10.6151
R2822 B.n1151 B.n1 10.6151
R2823 B.n1151 B.n1150 10.6151
R2824 B.n1150 B.n1149 10.6151
R2825 B.n1149 B.n10 10.6151
R2826 B.n1143 B.n10 10.6151
R2827 B.n1143 B.n1142 10.6151
R2828 B.n1142 B.n1141 10.6151
R2829 B.n1141 B.n17 10.6151
R2830 B.n1135 B.n17 10.6151
R2831 B.n1135 B.n1134 10.6151
R2832 B.n1134 B.n1133 10.6151
R2833 B.n1133 B.n24 10.6151
R2834 B.n1127 B.n24 10.6151
R2835 B.n1127 B.n1126 10.6151
R2836 B.n1126 B.n1125 10.6151
R2837 B.n1125 B.n31 10.6151
R2838 B.n1119 B.n31 10.6151
R2839 B.n1119 B.n1118 10.6151
R2840 B.n1118 B.n1117 10.6151
R2841 B.n1117 B.n38 10.6151
R2842 B.n1111 B.n38 10.6151
R2843 B.n1111 B.n1110 10.6151
R2844 B.n1110 B.n1109 10.6151
R2845 B.n1109 B.n45 10.6151
R2846 B.n1103 B.n45 10.6151
R2847 B.n1103 B.n1102 10.6151
R2848 B.n1102 B.n1101 10.6151
R2849 B.n1101 B.n52 10.6151
R2850 B.n1095 B.n52 10.6151
R2851 B.n1095 B.n1094 10.6151
R2852 B.n1094 B.n1093 10.6151
R2853 B.n1093 B.n59 10.6151
R2854 B.n1087 B.n59 10.6151
R2855 B.n1087 B.n1086 10.6151
R2856 B.n1086 B.n1085 10.6151
R2857 B.n1085 B.n66 10.6151
R2858 B.n1079 B.n66 10.6151
R2859 B.n1079 B.n1078 10.6151
R2860 B.n1078 B.n1077 10.6151
R2861 B.n1077 B.n73 10.6151
R2862 B.n1071 B.n73 10.6151
R2863 B.n1071 B.n1070 10.6151
R2864 B.n1070 B.n1069 10.6151
R2865 B.n1069 B.n80 10.6151
R2866 B.n1063 B.n80 10.6151
R2867 B.n1063 B.n1062 10.6151
R2868 B.n1062 B.n1061 10.6151
R2869 B.n1061 B.n87 10.6151
R2870 B.n1055 B.n87 10.6151
R2871 B.n1055 B.n1054 10.6151
R2872 B.n1054 B.n1053 10.6151
R2873 B.n1053 B.n94 10.6151
R2874 B.n1047 B.n94 10.6151
R2875 B.n1047 B.n1046 10.6151
R2876 B.n1046 B.n1045 10.6151
R2877 B.n1045 B.n101 10.6151
R2878 B.n1039 B.n101 10.6151
R2879 B.n1039 B.n1038 10.6151
R2880 B.n1038 B.n1037 10.6151
R2881 B.n1037 B.n108 10.6151
R2882 B.n1031 B.n108 10.6151
R2883 B.n1031 B.n1030 10.6151
R2884 B.n1030 B.n1029 10.6151
R2885 B.n1029 B.n115 10.6151
R2886 B.n1023 B.n115 10.6151
R2887 B.n1023 B.n1022 10.6151
R2888 B.n1022 B.n1021 10.6151
R2889 B.n1021 B.n122 10.6151
R2890 B.n796 B.t7 9.87187
R2891 B.n1067 B.t3 9.87187
R2892 B.n255 B.n176 9.36635
R2893 B.n278 B.n173 9.36635
R2894 B.n639 B.n638 9.36635
R2895 B.n617 B.n616 9.36635
R2896 B.n868 B.t1 5.92332
R2897 B.n1115 B.t6 5.92332
R2898 B.n1157 B.n0 2.81026
R2899 B.n1157 B.n1 2.81026
R2900 B.n832 B.t5 1.97477
R2901 B.n1091 B.t4 1.97477
R2902 B.n258 B.n176 1.24928
R2903 B.n275 B.n173 1.24928
R2904 B.n638 B.n637 1.24928
R2905 B.n618 B.n617 1.24928
R2906 VP.n23 VP.n22 161.3
R2907 VP.n24 VP.n19 161.3
R2908 VP.n26 VP.n25 161.3
R2909 VP.n27 VP.n18 161.3
R2910 VP.n29 VP.n28 161.3
R2911 VP.n30 VP.n17 161.3
R2912 VP.n32 VP.n31 161.3
R2913 VP.n33 VP.n16 161.3
R2914 VP.n36 VP.n35 161.3
R2915 VP.n37 VP.n15 161.3
R2916 VP.n39 VP.n38 161.3
R2917 VP.n40 VP.n14 161.3
R2918 VP.n42 VP.n41 161.3
R2919 VP.n43 VP.n13 161.3
R2920 VP.n45 VP.n44 161.3
R2921 VP.n46 VP.n12 161.3
R2922 VP.n88 VP.n0 161.3
R2923 VP.n87 VP.n86 161.3
R2924 VP.n85 VP.n1 161.3
R2925 VP.n84 VP.n83 161.3
R2926 VP.n82 VP.n2 161.3
R2927 VP.n81 VP.n80 161.3
R2928 VP.n79 VP.n3 161.3
R2929 VP.n78 VP.n77 161.3
R2930 VP.n75 VP.n4 161.3
R2931 VP.n74 VP.n73 161.3
R2932 VP.n72 VP.n5 161.3
R2933 VP.n71 VP.n70 161.3
R2934 VP.n69 VP.n6 161.3
R2935 VP.n68 VP.n67 161.3
R2936 VP.n66 VP.n7 161.3
R2937 VP.n65 VP.n64 161.3
R2938 VP.n62 VP.n8 161.3
R2939 VP.n61 VP.n60 161.3
R2940 VP.n59 VP.n9 161.3
R2941 VP.n58 VP.n57 161.3
R2942 VP.n56 VP.n10 161.3
R2943 VP.n55 VP.n54 161.3
R2944 VP.n53 VP.n11 161.3
R2945 VP.n52 VP.n51 161.3
R2946 VP.n20 VP.t3 104.632
R2947 VP.n50 VP.t4 72.3638
R2948 VP.n63 VP.t0 72.3638
R2949 VP.n76 VP.t7 72.3638
R2950 VP.n89 VP.t5 72.3638
R2951 VP.n47 VP.t2 72.3638
R2952 VP.n34 VP.t1 72.3638
R2953 VP.n21 VP.t6 72.3638
R2954 VP.n50 VP.n49 59.7554
R2955 VP.n90 VP.n89 59.7554
R2956 VP.n48 VP.n47 59.7554
R2957 VP.n21 VP.n20 59.5588
R2958 VP.n70 VP.n69 56.5617
R2959 VP.n28 VP.n27 56.5617
R2960 VP.n49 VP.n48 56.3681
R2961 VP.n57 VP.n56 51.2335
R2962 VP.n83 VP.n82 51.2335
R2963 VP.n41 VP.n40 51.2335
R2964 VP.n56 VP.n55 29.9206
R2965 VP.n83 VP.n1 29.9206
R2966 VP.n41 VP.n13 29.9206
R2967 VP.n51 VP.n11 24.5923
R2968 VP.n55 VP.n11 24.5923
R2969 VP.n57 VP.n9 24.5923
R2970 VP.n61 VP.n9 24.5923
R2971 VP.n62 VP.n61 24.5923
R2972 VP.n64 VP.n7 24.5923
R2973 VP.n68 VP.n7 24.5923
R2974 VP.n69 VP.n68 24.5923
R2975 VP.n70 VP.n5 24.5923
R2976 VP.n74 VP.n5 24.5923
R2977 VP.n75 VP.n74 24.5923
R2978 VP.n77 VP.n3 24.5923
R2979 VP.n81 VP.n3 24.5923
R2980 VP.n82 VP.n81 24.5923
R2981 VP.n87 VP.n1 24.5923
R2982 VP.n88 VP.n87 24.5923
R2983 VP.n45 VP.n13 24.5923
R2984 VP.n46 VP.n45 24.5923
R2985 VP.n28 VP.n17 24.5923
R2986 VP.n32 VP.n17 24.5923
R2987 VP.n33 VP.n32 24.5923
R2988 VP.n35 VP.n15 24.5923
R2989 VP.n39 VP.n15 24.5923
R2990 VP.n40 VP.n39 24.5923
R2991 VP.n22 VP.n19 24.5923
R2992 VP.n26 VP.n19 24.5923
R2993 VP.n27 VP.n26 24.5923
R2994 VP.n51 VP.n50 22.625
R2995 VP.n89 VP.n88 22.625
R2996 VP.n47 VP.n46 22.625
R2997 VP.n64 VP.n63 15.7393
R2998 VP.n76 VP.n75 15.7393
R2999 VP.n34 VP.n33 15.7393
R3000 VP.n22 VP.n21 15.7393
R3001 VP.n63 VP.n62 8.85356
R3002 VP.n77 VP.n76 8.85356
R3003 VP.n35 VP.n34 8.85356
R3004 VP.n23 VP.n20 2.58849
R3005 VP.n48 VP.n12 0.417304
R3006 VP.n52 VP.n49 0.417304
R3007 VP.n90 VP.n0 0.417304
R3008 VP VP.n90 0.394524
R3009 VP.n24 VP.n23 0.189894
R3010 VP.n25 VP.n24 0.189894
R3011 VP.n25 VP.n18 0.189894
R3012 VP.n29 VP.n18 0.189894
R3013 VP.n30 VP.n29 0.189894
R3014 VP.n31 VP.n30 0.189894
R3015 VP.n31 VP.n16 0.189894
R3016 VP.n36 VP.n16 0.189894
R3017 VP.n37 VP.n36 0.189894
R3018 VP.n38 VP.n37 0.189894
R3019 VP.n38 VP.n14 0.189894
R3020 VP.n42 VP.n14 0.189894
R3021 VP.n43 VP.n42 0.189894
R3022 VP.n44 VP.n43 0.189894
R3023 VP.n44 VP.n12 0.189894
R3024 VP.n53 VP.n52 0.189894
R3025 VP.n54 VP.n53 0.189894
R3026 VP.n54 VP.n10 0.189894
R3027 VP.n58 VP.n10 0.189894
R3028 VP.n59 VP.n58 0.189894
R3029 VP.n60 VP.n59 0.189894
R3030 VP.n60 VP.n8 0.189894
R3031 VP.n65 VP.n8 0.189894
R3032 VP.n66 VP.n65 0.189894
R3033 VP.n67 VP.n66 0.189894
R3034 VP.n67 VP.n6 0.189894
R3035 VP.n71 VP.n6 0.189894
R3036 VP.n72 VP.n71 0.189894
R3037 VP.n73 VP.n72 0.189894
R3038 VP.n73 VP.n4 0.189894
R3039 VP.n78 VP.n4 0.189894
R3040 VP.n79 VP.n78 0.189894
R3041 VP.n80 VP.n79 0.189894
R3042 VP.n80 VP.n2 0.189894
R3043 VP.n84 VP.n2 0.189894
R3044 VP.n85 VP.n84 0.189894
R3045 VP.n86 VP.n85 0.189894
R3046 VP.n86 VP.n0 0.189894
R3047 VDD1 VDD1.n0 64.7083
R3048 VDD1.n3 VDD1.n2 64.5946
R3049 VDD1.n3 VDD1.n1 64.5946
R3050 VDD1.n5 VDD1.n4 62.8655
R3051 VDD1.n5 VDD1.n3 50.2207
R3052 VDD1.n4 VDD1.t6 1.73127
R3053 VDD1.n4 VDD1.t5 1.73127
R3054 VDD1.n0 VDD1.t4 1.73127
R3055 VDD1.n0 VDD1.t1 1.73127
R3056 VDD1.n2 VDD1.t0 1.73127
R3057 VDD1.n2 VDD1.t2 1.73127
R3058 VDD1.n1 VDD1.t3 1.73127
R3059 VDD1.n1 VDD1.t7 1.73127
R3060 VDD1 VDD1.n5 1.72679
C0 VTAIL VDD1 8.45586f
C1 VTAIL VDD2 8.51839f
C2 VTAIL VP 9.69066f
C3 VDD1 VDD2 2.40504f
C4 VDD1 VP 9.344299f
C5 VTAIL VN 9.67655f
C6 VP VDD2 0.648697f
C7 VDD1 VN 0.154185f
C8 VN VDD2 8.851789f
C9 VP VN 9.035179f
C10 VDD2 B 6.576238f
C11 VDD1 B 7.14492f
C12 VTAIL B 10.960874f
C13 VN B 20.154982f
C14 VP B 18.818071f
C15 VDD1.t4 B 0.251289f
C16 VDD1.t1 B 0.251289f
C17 VDD1.n0 B 2.25392f
C18 VDD1.t3 B 0.251289f
C19 VDD1.t7 B 0.251289f
C20 VDD1.n1 B 2.25241f
C21 VDD1.t0 B 0.251289f
C22 VDD1.t2 B 0.251289f
C23 VDD1.n2 B 2.25241f
C24 VDD1.n3 B 4.439529f
C25 VDD1.t6 B 0.251289f
C26 VDD1.t5 B 0.251289f
C27 VDD1.n4 B 2.23328f
C28 VDD1.n5 B 3.73473f
C29 VP.n0 B 0.033319f
C30 VP.t5 B 2.10127f
C31 VP.n1 B 0.035111f
C32 VP.n2 B 0.017719f
C33 VP.n3 B 0.032858f
C34 VP.n4 B 0.017719f
C35 VP.t7 B 2.10127f
C36 VP.n5 B 0.032858f
C37 VP.n6 B 0.017719f
C38 VP.n7 B 0.032858f
C39 VP.n8 B 0.017719f
C40 VP.t0 B 2.10127f
C41 VP.n9 B 0.032858f
C42 VP.n10 B 0.017719f
C43 VP.n11 B 0.032858f
C44 VP.n12 B 0.033319f
C45 VP.t2 B 2.10127f
C46 VP.n13 B 0.035111f
C47 VP.n14 B 0.017719f
C48 VP.n15 B 0.032858f
C49 VP.n16 B 0.017719f
C50 VP.t1 B 2.10127f
C51 VP.n17 B 0.032858f
C52 VP.n18 B 0.017719f
C53 VP.n19 B 0.032858f
C54 VP.t3 B 2.37137f
C55 VP.n20 B 0.765272f
C56 VP.t6 B 2.10127f
C57 VP.n21 B 0.803223f
C58 VP.n22 B 0.027018f
C59 VP.n23 B 0.230549f
C60 VP.n24 B 0.017719f
C61 VP.n25 B 0.017719f
C62 VP.n26 B 0.032858f
C63 VP.n27 B 0.025757f
C64 VP.n28 B 0.025757f
C65 VP.n29 B 0.017719f
C66 VP.n30 B 0.017719f
C67 VP.n31 B 0.017719f
C68 VP.n32 B 0.032858f
C69 VP.n33 B 0.027018f
C70 VP.n34 B 0.737667f
C71 VP.n35 B 0.022476f
C72 VP.n36 B 0.017719f
C73 VP.n37 B 0.017719f
C74 VP.n38 B 0.017719f
C75 VP.n39 B 0.032858f
C76 VP.n40 B 0.032014f
C77 VP.n41 B 0.017246f
C78 VP.n42 B 0.017719f
C79 VP.n43 B 0.017719f
C80 VP.n44 B 0.017719f
C81 VP.n45 B 0.032858f
C82 VP.n46 B 0.03156f
C83 VP.n47 B 0.815275f
C84 VP.n48 B 1.21181f
C85 VP.n49 B 1.22314f
C86 VP.t4 B 2.10127f
C87 VP.n50 B 0.815275f
C88 VP.n51 B 0.03156f
C89 VP.n52 B 0.033319f
C90 VP.n53 B 0.017719f
C91 VP.n54 B 0.017719f
C92 VP.n55 B 0.035111f
C93 VP.n56 B 0.017246f
C94 VP.n57 B 0.032014f
C95 VP.n58 B 0.017719f
C96 VP.n59 B 0.017719f
C97 VP.n60 B 0.017719f
C98 VP.n61 B 0.032858f
C99 VP.n62 B 0.022476f
C100 VP.n63 B 0.737667f
C101 VP.n64 B 0.027018f
C102 VP.n65 B 0.017719f
C103 VP.n66 B 0.017719f
C104 VP.n67 B 0.017719f
C105 VP.n68 B 0.032858f
C106 VP.n69 B 0.025757f
C107 VP.n70 B 0.025757f
C108 VP.n71 B 0.017719f
C109 VP.n72 B 0.017719f
C110 VP.n73 B 0.017719f
C111 VP.n74 B 0.032858f
C112 VP.n75 B 0.027018f
C113 VP.n76 B 0.737667f
C114 VP.n77 B 0.022476f
C115 VP.n78 B 0.017719f
C116 VP.n79 B 0.017719f
C117 VP.n80 B 0.017719f
C118 VP.n81 B 0.032858f
C119 VP.n82 B 0.032014f
C120 VP.n83 B 0.017246f
C121 VP.n84 B 0.017719f
C122 VP.n85 B 0.017719f
C123 VP.n86 B 0.017719f
C124 VP.n87 B 0.032858f
C125 VP.n88 B 0.03156f
C126 VP.n89 B 0.815275f
C127 VP.n90 B 0.052877f
C128 VTAIL.t8 B 0.189824f
C129 VTAIL.t14 B 0.189824f
C130 VTAIL.n0 B 1.62614f
C131 VTAIL.n1 B 0.450371f
C132 VTAIL.n2 B 0.029514f
C133 VTAIL.n3 B 0.020998f
C134 VTAIL.n4 B 0.011283f
C135 VTAIL.n5 B 0.02667f
C136 VTAIL.n6 B 0.011947f
C137 VTAIL.n7 B 0.020998f
C138 VTAIL.n8 B 0.011283f
C139 VTAIL.n9 B 0.02667f
C140 VTAIL.n10 B 0.011615f
C141 VTAIL.n11 B 0.020998f
C142 VTAIL.n12 B 0.011947f
C143 VTAIL.n13 B 0.02667f
C144 VTAIL.n14 B 0.011947f
C145 VTAIL.n15 B 0.020998f
C146 VTAIL.n16 B 0.011283f
C147 VTAIL.n17 B 0.02667f
C148 VTAIL.n18 B 0.011947f
C149 VTAIL.n19 B 1.007f
C150 VTAIL.n20 B 0.011283f
C151 VTAIL.t9 B 0.04498f
C152 VTAIL.n21 B 0.146877f
C153 VTAIL.n22 B 0.018853f
C154 VTAIL.n23 B 0.020002f
C155 VTAIL.n24 B 0.02667f
C156 VTAIL.n25 B 0.011947f
C157 VTAIL.n26 B 0.011283f
C158 VTAIL.n27 B 0.020998f
C159 VTAIL.n28 B 0.020998f
C160 VTAIL.n29 B 0.011283f
C161 VTAIL.n30 B 0.011947f
C162 VTAIL.n31 B 0.02667f
C163 VTAIL.n32 B 0.02667f
C164 VTAIL.n33 B 0.011947f
C165 VTAIL.n34 B 0.011283f
C166 VTAIL.n35 B 0.020998f
C167 VTAIL.n36 B 0.020998f
C168 VTAIL.n37 B 0.011283f
C169 VTAIL.n38 B 0.011283f
C170 VTAIL.n39 B 0.011947f
C171 VTAIL.n40 B 0.02667f
C172 VTAIL.n41 B 0.02667f
C173 VTAIL.n42 B 0.02667f
C174 VTAIL.n43 B 0.011615f
C175 VTAIL.n44 B 0.011283f
C176 VTAIL.n45 B 0.020998f
C177 VTAIL.n46 B 0.020998f
C178 VTAIL.n47 B 0.011283f
C179 VTAIL.n48 B 0.011947f
C180 VTAIL.n49 B 0.02667f
C181 VTAIL.n50 B 0.02667f
C182 VTAIL.n51 B 0.011947f
C183 VTAIL.n52 B 0.011283f
C184 VTAIL.n53 B 0.020998f
C185 VTAIL.n54 B 0.020998f
C186 VTAIL.n55 B 0.011283f
C187 VTAIL.n56 B 0.011947f
C188 VTAIL.n57 B 0.02667f
C189 VTAIL.n58 B 0.057735f
C190 VTAIL.n59 B 0.011947f
C191 VTAIL.n60 B 0.011283f
C192 VTAIL.n61 B 0.049683f
C193 VTAIL.n62 B 0.03234f
C194 VTAIL.n63 B 0.291844f
C195 VTAIL.n64 B 0.029514f
C196 VTAIL.n65 B 0.020998f
C197 VTAIL.n66 B 0.011283f
C198 VTAIL.n67 B 0.02667f
C199 VTAIL.n68 B 0.011947f
C200 VTAIL.n69 B 0.020998f
C201 VTAIL.n70 B 0.011283f
C202 VTAIL.n71 B 0.02667f
C203 VTAIL.n72 B 0.011615f
C204 VTAIL.n73 B 0.020998f
C205 VTAIL.n74 B 0.011947f
C206 VTAIL.n75 B 0.02667f
C207 VTAIL.n76 B 0.011947f
C208 VTAIL.n77 B 0.020998f
C209 VTAIL.n78 B 0.011283f
C210 VTAIL.n79 B 0.02667f
C211 VTAIL.n80 B 0.011947f
C212 VTAIL.n81 B 1.007f
C213 VTAIL.n82 B 0.011283f
C214 VTAIL.t2 B 0.04498f
C215 VTAIL.n83 B 0.146877f
C216 VTAIL.n84 B 0.018853f
C217 VTAIL.n85 B 0.020002f
C218 VTAIL.n86 B 0.02667f
C219 VTAIL.n87 B 0.011947f
C220 VTAIL.n88 B 0.011283f
C221 VTAIL.n89 B 0.020998f
C222 VTAIL.n90 B 0.020998f
C223 VTAIL.n91 B 0.011283f
C224 VTAIL.n92 B 0.011947f
C225 VTAIL.n93 B 0.02667f
C226 VTAIL.n94 B 0.02667f
C227 VTAIL.n95 B 0.011947f
C228 VTAIL.n96 B 0.011283f
C229 VTAIL.n97 B 0.020998f
C230 VTAIL.n98 B 0.020998f
C231 VTAIL.n99 B 0.011283f
C232 VTAIL.n100 B 0.011283f
C233 VTAIL.n101 B 0.011947f
C234 VTAIL.n102 B 0.02667f
C235 VTAIL.n103 B 0.02667f
C236 VTAIL.n104 B 0.02667f
C237 VTAIL.n105 B 0.011615f
C238 VTAIL.n106 B 0.011283f
C239 VTAIL.n107 B 0.020998f
C240 VTAIL.n108 B 0.020998f
C241 VTAIL.n109 B 0.011283f
C242 VTAIL.n110 B 0.011947f
C243 VTAIL.n111 B 0.02667f
C244 VTAIL.n112 B 0.02667f
C245 VTAIL.n113 B 0.011947f
C246 VTAIL.n114 B 0.011283f
C247 VTAIL.n115 B 0.020998f
C248 VTAIL.n116 B 0.020998f
C249 VTAIL.n117 B 0.011283f
C250 VTAIL.n118 B 0.011947f
C251 VTAIL.n119 B 0.02667f
C252 VTAIL.n120 B 0.057735f
C253 VTAIL.n121 B 0.011947f
C254 VTAIL.n122 B 0.011283f
C255 VTAIL.n123 B 0.049683f
C256 VTAIL.n124 B 0.03234f
C257 VTAIL.n125 B 0.291844f
C258 VTAIL.t5 B 0.189824f
C259 VTAIL.t1 B 0.189824f
C260 VTAIL.n126 B 1.62614f
C261 VTAIL.n127 B 0.687908f
C262 VTAIL.n128 B 0.029514f
C263 VTAIL.n129 B 0.020998f
C264 VTAIL.n130 B 0.011283f
C265 VTAIL.n131 B 0.02667f
C266 VTAIL.n132 B 0.011947f
C267 VTAIL.n133 B 0.020998f
C268 VTAIL.n134 B 0.011283f
C269 VTAIL.n135 B 0.02667f
C270 VTAIL.n136 B 0.011615f
C271 VTAIL.n137 B 0.020998f
C272 VTAIL.n138 B 0.011947f
C273 VTAIL.n139 B 0.02667f
C274 VTAIL.n140 B 0.011947f
C275 VTAIL.n141 B 0.020998f
C276 VTAIL.n142 B 0.011283f
C277 VTAIL.n143 B 0.02667f
C278 VTAIL.n144 B 0.011947f
C279 VTAIL.n145 B 1.007f
C280 VTAIL.n146 B 0.011283f
C281 VTAIL.t7 B 0.04498f
C282 VTAIL.n147 B 0.146877f
C283 VTAIL.n148 B 0.018853f
C284 VTAIL.n149 B 0.020002f
C285 VTAIL.n150 B 0.02667f
C286 VTAIL.n151 B 0.011947f
C287 VTAIL.n152 B 0.011283f
C288 VTAIL.n153 B 0.020998f
C289 VTAIL.n154 B 0.020998f
C290 VTAIL.n155 B 0.011283f
C291 VTAIL.n156 B 0.011947f
C292 VTAIL.n157 B 0.02667f
C293 VTAIL.n158 B 0.02667f
C294 VTAIL.n159 B 0.011947f
C295 VTAIL.n160 B 0.011283f
C296 VTAIL.n161 B 0.020998f
C297 VTAIL.n162 B 0.020998f
C298 VTAIL.n163 B 0.011283f
C299 VTAIL.n164 B 0.011283f
C300 VTAIL.n165 B 0.011947f
C301 VTAIL.n166 B 0.02667f
C302 VTAIL.n167 B 0.02667f
C303 VTAIL.n168 B 0.02667f
C304 VTAIL.n169 B 0.011615f
C305 VTAIL.n170 B 0.011283f
C306 VTAIL.n171 B 0.020998f
C307 VTAIL.n172 B 0.020998f
C308 VTAIL.n173 B 0.011283f
C309 VTAIL.n174 B 0.011947f
C310 VTAIL.n175 B 0.02667f
C311 VTAIL.n176 B 0.02667f
C312 VTAIL.n177 B 0.011947f
C313 VTAIL.n178 B 0.011283f
C314 VTAIL.n179 B 0.020998f
C315 VTAIL.n180 B 0.020998f
C316 VTAIL.n181 B 0.011283f
C317 VTAIL.n182 B 0.011947f
C318 VTAIL.n183 B 0.02667f
C319 VTAIL.n184 B 0.057735f
C320 VTAIL.n185 B 0.011947f
C321 VTAIL.n186 B 0.011283f
C322 VTAIL.n187 B 0.049683f
C323 VTAIL.n188 B 0.03234f
C324 VTAIL.n189 B 1.45402f
C325 VTAIL.n190 B 0.029514f
C326 VTAIL.n191 B 0.020998f
C327 VTAIL.n192 B 0.011283f
C328 VTAIL.n193 B 0.02667f
C329 VTAIL.n194 B 0.011947f
C330 VTAIL.n195 B 0.020998f
C331 VTAIL.n196 B 0.011283f
C332 VTAIL.n197 B 0.02667f
C333 VTAIL.n198 B 0.011615f
C334 VTAIL.n199 B 0.020998f
C335 VTAIL.n200 B 0.011615f
C336 VTAIL.n201 B 0.011283f
C337 VTAIL.n202 B 0.02667f
C338 VTAIL.n203 B 0.02667f
C339 VTAIL.n204 B 0.011947f
C340 VTAIL.n205 B 0.020998f
C341 VTAIL.n206 B 0.011283f
C342 VTAIL.n207 B 0.02667f
C343 VTAIL.n208 B 0.011947f
C344 VTAIL.n209 B 1.007f
C345 VTAIL.n210 B 0.011283f
C346 VTAIL.t12 B 0.04498f
C347 VTAIL.n211 B 0.146877f
C348 VTAIL.n212 B 0.018853f
C349 VTAIL.n213 B 0.020002f
C350 VTAIL.n214 B 0.02667f
C351 VTAIL.n215 B 0.011947f
C352 VTAIL.n216 B 0.011283f
C353 VTAIL.n217 B 0.020998f
C354 VTAIL.n218 B 0.020998f
C355 VTAIL.n219 B 0.011283f
C356 VTAIL.n220 B 0.011947f
C357 VTAIL.n221 B 0.02667f
C358 VTAIL.n222 B 0.02667f
C359 VTAIL.n223 B 0.011947f
C360 VTAIL.n224 B 0.011283f
C361 VTAIL.n225 B 0.020998f
C362 VTAIL.n226 B 0.020998f
C363 VTAIL.n227 B 0.011283f
C364 VTAIL.n228 B 0.011947f
C365 VTAIL.n229 B 0.02667f
C366 VTAIL.n230 B 0.02667f
C367 VTAIL.n231 B 0.011947f
C368 VTAIL.n232 B 0.011283f
C369 VTAIL.n233 B 0.020998f
C370 VTAIL.n234 B 0.020998f
C371 VTAIL.n235 B 0.011283f
C372 VTAIL.n236 B 0.011947f
C373 VTAIL.n237 B 0.02667f
C374 VTAIL.n238 B 0.02667f
C375 VTAIL.n239 B 0.011947f
C376 VTAIL.n240 B 0.011283f
C377 VTAIL.n241 B 0.020998f
C378 VTAIL.n242 B 0.020998f
C379 VTAIL.n243 B 0.011283f
C380 VTAIL.n244 B 0.011947f
C381 VTAIL.n245 B 0.02667f
C382 VTAIL.n246 B 0.057735f
C383 VTAIL.n247 B 0.011947f
C384 VTAIL.n248 B 0.011283f
C385 VTAIL.n249 B 0.049683f
C386 VTAIL.n250 B 0.03234f
C387 VTAIL.n251 B 1.45402f
C388 VTAIL.t10 B 0.189824f
C389 VTAIL.t15 B 0.189824f
C390 VTAIL.n252 B 1.62615f
C391 VTAIL.n253 B 0.687899f
C392 VTAIL.n254 B 0.029514f
C393 VTAIL.n255 B 0.020998f
C394 VTAIL.n256 B 0.011283f
C395 VTAIL.n257 B 0.02667f
C396 VTAIL.n258 B 0.011947f
C397 VTAIL.n259 B 0.020998f
C398 VTAIL.n260 B 0.011283f
C399 VTAIL.n261 B 0.02667f
C400 VTAIL.n262 B 0.011615f
C401 VTAIL.n263 B 0.020998f
C402 VTAIL.n264 B 0.011615f
C403 VTAIL.n265 B 0.011283f
C404 VTAIL.n266 B 0.02667f
C405 VTAIL.n267 B 0.02667f
C406 VTAIL.n268 B 0.011947f
C407 VTAIL.n269 B 0.020998f
C408 VTAIL.n270 B 0.011283f
C409 VTAIL.n271 B 0.02667f
C410 VTAIL.n272 B 0.011947f
C411 VTAIL.n273 B 1.007f
C412 VTAIL.n274 B 0.011283f
C413 VTAIL.t11 B 0.04498f
C414 VTAIL.n275 B 0.146877f
C415 VTAIL.n276 B 0.018853f
C416 VTAIL.n277 B 0.020002f
C417 VTAIL.n278 B 0.02667f
C418 VTAIL.n279 B 0.011947f
C419 VTAIL.n280 B 0.011283f
C420 VTAIL.n281 B 0.020998f
C421 VTAIL.n282 B 0.020998f
C422 VTAIL.n283 B 0.011283f
C423 VTAIL.n284 B 0.011947f
C424 VTAIL.n285 B 0.02667f
C425 VTAIL.n286 B 0.02667f
C426 VTAIL.n287 B 0.011947f
C427 VTAIL.n288 B 0.011283f
C428 VTAIL.n289 B 0.020998f
C429 VTAIL.n290 B 0.020998f
C430 VTAIL.n291 B 0.011283f
C431 VTAIL.n292 B 0.011947f
C432 VTAIL.n293 B 0.02667f
C433 VTAIL.n294 B 0.02667f
C434 VTAIL.n295 B 0.011947f
C435 VTAIL.n296 B 0.011283f
C436 VTAIL.n297 B 0.020998f
C437 VTAIL.n298 B 0.020998f
C438 VTAIL.n299 B 0.011283f
C439 VTAIL.n300 B 0.011947f
C440 VTAIL.n301 B 0.02667f
C441 VTAIL.n302 B 0.02667f
C442 VTAIL.n303 B 0.011947f
C443 VTAIL.n304 B 0.011283f
C444 VTAIL.n305 B 0.020998f
C445 VTAIL.n306 B 0.020998f
C446 VTAIL.n307 B 0.011283f
C447 VTAIL.n308 B 0.011947f
C448 VTAIL.n309 B 0.02667f
C449 VTAIL.n310 B 0.057735f
C450 VTAIL.n311 B 0.011947f
C451 VTAIL.n312 B 0.011283f
C452 VTAIL.n313 B 0.049683f
C453 VTAIL.n314 B 0.03234f
C454 VTAIL.n315 B 0.291844f
C455 VTAIL.n316 B 0.029514f
C456 VTAIL.n317 B 0.020998f
C457 VTAIL.n318 B 0.011283f
C458 VTAIL.n319 B 0.02667f
C459 VTAIL.n320 B 0.011947f
C460 VTAIL.n321 B 0.020998f
C461 VTAIL.n322 B 0.011283f
C462 VTAIL.n323 B 0.02667f
C463 VTAIL.n324 B 0.011615f
C464 VTAIL.n325 B 0.020998f
C465 VTAIL.n326 B 0.011615f
C466 VTAIL.n327 B 0.011283f
C467 VTAIL.n328 B 0.02667f
C468 VTAIL.n329 B 0.02667f
C469 VTAIL.n330 B 0.011947f
C470 VTAIL.n331 B 0.020998f
C471 VTAIL.n332 B 0.011283f
C472 VTAIL.n333 B 0.02667f
C473 VTAIL.n334 B 0.011947f
C474 VTAIL.n335 B 1.007f
C475 VTAIL.n336 B 0.011283f
C476 VTAIL.t0 B 0.04498f
C477 VTAIL.n337 B 0.146877f
C478 VTAIL.n338 B 0.018853f
C479 VTAIL.n339 B 0.020002f
C480 VTAIL.n340 B 0.02667f
C481 VTAIL.n341 B 0.011947f
C482 VTAIL.n342 B 0.011283f
C483 VTAIL.n343 B 0.020998f
C484 VTAIL.n344 B 0.020998f
C485 VTAIL.n345 B 0.011283f
C486 VTAIL.n346 B 0.011947f
C487 VTAIL.n347 B 0.02667f
C488 VTAIL.n348 B 0.02667f
C489 VTAIL.n349 B 0.011947f
C490 VTAIL.n350 B 0.011283f
C491 VTAIL.n351 B 0.020998f
C492 VTAIL.n352 B 0.020998f
C493 VTAIL.n353 B 0.011283f
C494 VTAIL.n354 B 0.011947f
C495 VTAIL.n355 B 0.02667f
C496 VTAIL.n356 B 0.02667f
C497 VTAIL.n357 B 0.011947f
C498 VTAIL.n358 B 0.011283f
C499 VTAIL.n359 B 0.020998f
C500 VTAIL.n360 B 0.020998f
C501 VTAIL.n361 B 0.011283f
C502 VTAIL.n362 B 0.011947f
C503 VTAIL.n363 B 0.02667f
C504 VTAIL.n364 B 0.02667f
C505 VTAIL.n365 B 0.011947f
C506 VTAIL.n366 B 0.011283f
C507 VTAIL.n367 B 0.020998f
C508 VTAIL.n368 B 0.020998f
C509 VTAIL.n369 B 0.011283f
C510 VTAIL.n370 B 0.011947f
C511 VTAIL.n371 B 0.02667f
C512 VTAIL.n372 B 0.057735f
C513 VTAIL.n373 B 0.011947f
C514 VTAIL.n374 B 0.011283f
C515 VTAIL.n375 B 0.049683f
C516 VTAIL.n376 B 0.03234f
C517 VTAIL.n377 B 0.291844f
C518 VTAIL.t6 B 0.189824f
C519 VTAIL.t4 B 0.189824f
C520 VTAIL.n378 B 1.62615f
C521 VTAIL.n379 B 0.687899f
C522 VTAIL.n380 B 0.029514f
C523 VTAIL.n381 B 0.020998f
C524 VTAIL.n382 B 0.011283f
C525 VTAIL.n383 B 0.02667f
C526 VTAIL.n384 B 0.011947f
C527 VTAIL.n385 B 0.020998f
C528 VTAIL.n386 B 0.011283f
C529 VTAIL.n387 B 0.02667f
C530 VTAIL.n388 B 0.011615f
C531 VTAIL.n389 B 0.020998f
C532 VTAIL.n390 B 0.011615f
C533 VTAIL.n391 B 0.011283f
C534 VTAIL.n392 B 0.02667f
C535 VTAIL.n393 B 0.02667f
C536 VTAIL.n394 B 0.011947f
C537 VTAIL.n395 B 0.020998f
C538 VTAIL.n396 B 0.011283f
C539 VTAIL.n397 B 0.02667f
C540 VTAIL.n398 B 0.011947f
C541 VTAIL.n399 B 1.007f
C542 VTAIL.n400 B 0.011283f
C543 VTAIL.t3 B 0.04498f
C544 VTAIL.n401 B 0.146877f
C545 VTAIL.n402 B 0.018853f
C546 VTAIL.n403 B 0.020002f
C547 VTAIL.n404 B 0.02667f
C548 VTAIL.n405 B 0.011947f
C549 VTAIL.n406 B 0.011283f
C550 VTAIL.n407 B 0.020998f
C551 VTAIL.n408 B 0.020998f
C552 VTAIL.n409 B 0.011283f
C553 VTAIL.n410 B 0.011947f
C554 VTAIL.n411 B 0.02667f
C555 VTAIL.n412 B 0.02667f
C556 VTAIL.n413 B 0.011947f
C557 VTAIL.n414 B 0.011283f
C558 VTAIL.n415 B 0.020998f
C559 VTAIL.n416 B 0.020998f
C560 VTAIL.n417 B 0.011283f
C561 VTAIL.n418 B 0.011947f
C562 VTAIL.n419 B 0.02667f
C563 VTAIL.n420 B 0.02667f
C564 VTAIL.n421 B 0.011947f
C565 VTAIL.n422 B 0.011283f
C566 VTAIL.n423 B 0.020998f
C567 VTAIL.n424 B 0.020998f
C568 VTAIL.n425 B 0.011283f
C569 VTAIL.n426 B 0.011947f
C570 VTAIL.n427 B 0.02667f
C571 VTAIL.n428 B 0.02667f
C572 VTAIL.n429 B 0.011947f
C573 VTAIL.n430 B 0.011283f
C574 VTAIL.n431 B 0.020998f
C575 VTAIL.n432 B 0.020998f
C576 VTAIL.n433 B 0.011283f
C577 VTAIL.n434 B 0.011947f
C578 VTAIL.n435 B 0.02667f
C579 VTAIL.n436 B 0.057735f
C580 VTAIL.n437 B 0.011947f
C581 VTAIL.n438 B 0.011283f
C582 VTAIL.n439 B 0.049683f
C583 VTAIL.n440 B 0.03234f
C584 VTAIL.n441 B 1.45402f
C585 VTAIL.n442 B 0.029514f
C586 VTAIL.n443 B 0.020998f
C587 VTAIL.n444 B 0.011283f
C588 VTAIL.n445 B 0.02667f
C589 VTAIL.n446 B 0.011947f
C590 VTAIL.n447 B 0.020998f
C591 VTAIL.n448 B 0.011283f
C592 VTAIL.n449 B 0.02667f
C593 VTAIL.n450 B 0.011615f
C594 VTAIL.n451 B 0.020998f
C595 VTAIL.n452 B 0.011947f
C596 VTAIL.n453 B 0.02667f
C597 VTAIL.n454 B 0.011947f
C598 VTAIL.n455 B 0.020998f
C599 VTAIL.n456 B 0.011283f
C600 VTAIL.n457 B 0.02667f
C601 VTAIL.n458 B 0.011947f
C602 VTAIL.n459 B 1.007f
C603 VTAIL.n460 B 0.011283f
C604 VTAIL.t13 B 0.04498f
C605 VTAIL.n461 B 0.146877f
C606 VTAIL.n462 B 0.018853f
C607 VTAIL.n463 B 0.020002f
C608 VTAIL.n464 B 0.02667f
C609 VTAIL.n465 B 0.011947f
C610 VTAIL.n466 B 0.011283f
C611 VTAIL.n467 B 0.020998f
C612 VTAIL.n468 B 0.020998f
C613 VTAIL.n469 B 0.011283f
C614 VTAIL.n470 B 0.011947f
C615 VTAIL.n471 B 0.02667f
C616 VTAIL.n472 B 0.02667f
C617 VTAIL.n473 B 0.011947f
C618 VTAIL.n474 B 0.011283f
C619 VTAIL.n475 B 0.020998f
C620 VTAIL.n476 B 0.020998f
C621 VTAIL.n477 B 0.011283f
C622 VTAIL.n478 B 0.011283f
C623 VTAIL.n479 B 0.011947f
C624 VTAIL.n480 B 0.02667f
C625 VTAIL.n481 B 0.02667f
C626 VTAIL.n482 B 0.02667f
C627 VTAIL.n483 B 0.011615f
C628 VTAIL.n484 B 0.011283f
C629 VTAIL.n485 B 0.020998f
C630 VTAIL.n486 B 0.020998f
C631 VTAIL.n487 B 0.011283f
C632 VTAIL.n488 B 0.011947f
C633 VTAIL.n489 B 0.02667f
C634 VTAIL.n490 B 0.02667f
C635 VTAIL.n491 B 0.011947f
C636 VTAIL.n492 B 0.011283f
C637 VTAIL.n493 B 0.020998f
C638 VTAIL.n494 B 0.020998f
C639 VTAIL.n495 B 0.011283f
C640 VTAIL.n496 B 0.011947f
C641 VTAIL.n497 B 0.02667f
C642 VTAIL.n498 B 0.057735f
C643 VTAIL.n499 B 0.011947f
C644 VTAIL.n500 B 0.011283f
C645 VTAIL.n501 B 0.049683f
C646 VTAIL.n502 B 0.03234f
C647 VTAIL.n503 B 1.45008f
C648 VDD2.t3 B 0.247571f
C649 VDD2.t2 B 0.247571f
C650 VDD2.n0 B 2.21908f
C651 VDD2.t4 B 0.247571f
C652 VDD2.t7 B 0.247571f
C653 VDD2.n1 B 2.21908f
C654 VDD2.n2 B 4.31747f
C655 VDD2.t6 B 0.247571f
C656 VDD2.t0 B 0.247571f
C657 VDD2.n3 B 2.20025f
C658 VDD2.n4 B 3.64496f
C659 VDD2.t5 B 0.247571f
C660 VDD2.t1 B 0.247571f
C661 VDD2.n5 B 2.21904f
C662 VN.n0 B 0.032814f
C663 VN.t2 B 2.06941f
C664 VN.n1 B 0.034579f
C665 VN.n2 B 0.01745f
C666 VN.n3 B 0.03236f
C667 VN.n4 B 0.01745f
C668 VN.t1 B 2.06941f
C669 VN.n5 B 0.03236f
C670 VN.n6 B 0.01745f
C671 VN.n7 B 0.03236f
C672 VN.t6 B 2.33542f
C673 VN.n8 B 0.753667f
C674 VN.t7 B 2.06941f
C675 VN.n9 B 0.791045f
C676 VN.n10 B 0.026609f
C677 VN.n11 B 0.227053f
C678 VN.n12 B 0.01745f
C679 VN.n13 B 0.01745f
C680 VN.n14 B 0.03236f
C681 VN.n15 B 0.025366f
C682 VN.n16 B 0.025366f
C683 VN.n17 B 0.01745f
C684 VN.n18 B 0.01745f
C685 VN.n19 B 0.01745f
C686 VN.n20 B 0.03236f
C687 VN.n21 B 0.026609f
C688 VN.n22 B 0.726482f
C689 VN.n23 B 0.022135f
C690 VN.n24 B 0.01745f
C691 VN.n25 B 0.01745f
C692 VN.n26 B 0.01745f
C693 VN.n27 B 0.03236f
C694 VN.n28 B 0.031529f
C695 VN.n29 B 0.016985f
C696 VN.n30 B 0.01745f
C697 VN.n31 B 0.01745f
C698 VN.n32 B 0.01745f
C699 VN.n33 B 0.03236f
C700 VN.n34 B 0.031082f
C701 VN.n35 B 0.802914f
C702 VN.n36 B 0.052076f
C703 VN.n37 B 0.032814f
C704 VN.t3 B 2.06941f
C705 VN.n38 B 0.034579f
C706 VN.n39 B 0.01745f
C707 VN.n40 B 0.03236f
C708 VN.n41 B 0.01745f
C709 VN.t5 B 2.06941f
C710 VN.n42 B 0.03236f
C711 VN.n43 B 0.01745f
C712 VN.n44 B 0.03236f
C713 VN.t4 B 2.33542f
C714 VN.n45 B 0.753667f
C715 VN.t0 B 2.06941f
C716 VN.n46 B 0.791045f
C717 VN.n47 B 0.026609f
C718 VN.n48 B 0.227053f
C719 VN.n49 B 0.01745f
C720 VN.n50 B 0.01745f
C721 VN.n51 B 0.03236f
C722 VN.n52 B 0.025366f
C723 VN.n53 B 0.025366f
C724 VN.n54 B 0.01745f
C725 VN.n55 B 0.01745f
C726 VN.n56 B 0.01745f
C727 VN.n57 B 0.03236f
C728 VN.n58 B 0.026609f
C729 VN.n59 B 0.726482f
C730 VN.n60 B 0.022135f
C731 VN.n61 B 0.01745f
C732 VN.n62 B 0.01745f
C733 VN.n63 B 0.01745f
C734 VN.n64 B 0.03236f
C735 VN.n65 B 0.031529f
C736 VN.n66 B 0.016985f
C737 VN.n67 B 0.01745f
C738 VN.n68 B 0.01745f
C739 VN.n69 B 0.01745f
C740 VN.n70 B 0.03236f
C741 VN.n71 B 0.031082f
C742 VN.n72 B 0.802914f
C743 VN.n73 B 1.19761f
.ends

