* NGSPICE file created from diff_pair_sample_0756.ext - technology: sky130A

.subckt diff_pair_sample_0756 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X1 VDD1.t6 VP.t1 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X2 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X3 VTAIL.t6 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X4 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=1.6269 ps=10.19 w=9.86 l=3.08
X5 VDD1.t5 VP.t2 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=3.8454 ps=20.5 w=9.86 l=3.08
X6 VTAIL.t3 VN.t3 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=1.6269 ps=10.19 w=9.86 l=3.08
X7 VTAIL.t7 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X8 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=0 ps=0 w=9.86 l=3.08
X9 VTAIL.t11 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=1.6269 ps=10.19 w=9.86 l=3.08
X10 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=0 ps=0 w=9.86 l=3.08
X11 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=3.8454 ps=20.5 w=9.86 l=3.08
X12 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X13 VDD1.t3 VP.t4 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=3.8454 ps=20.5 w=9.86 l=3.08
X14 VTAIL.t14 VP.t5 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
X15 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=3.8454 ps=20.5 w=9.86 l=3.08
X16 VTAIL.t12 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=1.6269 ps=10.19 w=9.86 l=3.08
X17 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=0 ps=0 w=9.86 l=3.08
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8454 pd=20.5 as=0 ps=0 w=9.86 l=3.08
X19 VTAIL.t15 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6269 pd=10.19 as=1.6269 ps=10.19 w=9.86 l=3.08
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n19 VP.t3 110.55
R34 VP.n43 VP.t6 77.1518
R35 VP.n55 VP.t0 77.1518
R36 VP.n4 VP.t7 77.1518
R37 VP.n0 VP.t4 77.1518
R38 VP.n11 VP.t2 77.1518
R39 VP.n15 VP.t5 77.1518
R40 VP.n20 VP.t1 77.1518
R41 VP.n43 VP.n42 72.2935
R42 VP.n76 VP.n0 72.2935
R43 VP.n41 VP.n11 72.2935
R44 VP.n61 VP.n6 56.5617
R45 VP.n26 VP.n17 56.5617
R46 VP.n49 VP.n48 56.0773
R47 VP.n72 VP.n2 56.0773
R48 VP.n37 VP.n13 56.0773
R49 VP.n20 VP.n19 51.6451
R50 VP.n42 VP.n41 51.6283
R51 VP.n50 VP.n49 25.0767
R52 VP.n68 VP.n2 25.0767
R53 VP.n33 VP.n13 25.0767
R54 VP.n44 VP.n10 24.5923
R55 VP.n48 VP.n10 24.5923
R56 VP.n50 VP.n8 24.5923
R57 VP.n54 VP.n8 24.5923
R58 VP.n57 VP.n56 24.5923
R59 VP.n57 VP.n6 24.5923
R60 VP.n62 VP.n61 24.5923
R61 VP.n63 VP.n62 24.5923
R62 VP.n67 VP.n66 24.5923
R63 VP.n68 VP.n67 24.5923
R64 VP.n73 VP.n72 24.5923
R65 VP.n74 VP.n73 24.5923
R66 VP.n38 VP.n37 24.5923
R67 VP.n39 VP.n38 24.5923
R68 VP.n27 VP.n26 24.5923
R69 VP.n28 VP.n27 24.5923
R70 VP.n32 VP.n31 24.5923
R71 VP.n33 VP.n32 24.5923
R72 VP.n22 VP.n21 24.5923
R73 VP.n22 VP.n17 24.5923
R74 VP.n56 VP.n55 22.3791
R75 VP.n63 VP.n4 22.3791
R76 VP.n28 VP.n15 22.3791
R77 VP.n21 VP.n20 22.3791
R78 VP.n44 VP.n43 17.9525
R79 VP.n74 VP.n0 17.9525
R80 VP.n39 VP.n11 17.9525
R81 VP.n19 VP.n18 4.00187
R82 VP.n55 VP.n54 2.21377
R83 VP.n66 VP.n4 2.21377
R84 VP.n31 VP.n15 2.21377
R85 VP.n41 VP.n40 0.354861
R86 VP.n45 VP.n42 0.354861
R87 VP.n76 VP.n75 0.354861
R88 VP VP.n76 0.267071
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VTAIL.n11 VTAIL.t11 46.6626
R121 VTAIL.n10 VTAIL.t4 46.6626
R122 VTAIL.n7 VTAIL.t3 46.6626
R123 VTAIL.n14 VTAIL.t10 46.6626
R124 VTAIL.n15 VTAIL.t0 46.6624
R125 VTAIL.n2 VTAIL.t5 46.6624
R126 VTAIL.n3 VTAIL.t13 46.6624
R127 VTAIL.n6 VTAIL.t12 46.6624
R128 VTAIL.n13 VTAIL.n12 44.6545
R129 VTAIL.n9 VTAIL.n8 44.6545
R130 VTAIL.n1 VTAIL.n0 44.6543
R131 VTAIL.n5 VTAIL.n4 44.6543
R132 VTAIL.n15 VTAIL.n14 23.8065
R133 VTAIL.n7 VTAIL.n6 23.8065
R134 VTAIL.n9 VTAIL.n7 2.94016
R135 VTAIL.n10 VTAIL.n9 2.94016
R136 VTAIL.n13 VTAIL.n11 2.94016
R137 VTAIL.n14 VTAIL.n13 2.94016
R138 VTAIL.n6 VTAIL.n5 2.94016
R139 VTAIL.n5 VTAIL.n3 2.94016
R140 VTAIL.n2 VTAIL.n1 2.94016
R141 VTAIL VTAIL.n15 2.88197
R142 VTAIL.n0 VTAIL.t2 2.00861
R143 VTAIL.n0 VTAIL.t7 2.00861
R144 VTAIL.n4 VTAIL.t9 2.00861
R145 VTAIL.n4 VTAIL.t15 2.00861
R146 VTAIL.n12 VTAIL.t8 2.00861
R147 VTAIL.n12 VTAIL.t14 2.00861
R148 VTAIL.n8 VTAIL.t1 2.00861
R149 VTAIL.n8 VTAIL.t6 2.00861
R150 VTAIL.n11 VTAIL.n10 0.470328
R151 VTAIL.n3 VTAIL.n2 0.470328
R152 VTAIL VTAIL.n1 0.0586897
R153 VDD1 VDD1.n0 62.8613
R154 VDD1.n3 VDD1.n2 62.7476
R155 VDD1.n3 VDD1.n1 62.7476
R156 VDD1.n5 VDD1.n4 61.3333
R157 VDD1.n5 VDD1.n3 46.0268
R158 VDD1.n4 VDD1.t2 2.00861
R159 VDD1.n4 VDD1.t5 2.00861
R160 VDD1.n0 VDD1.t4 2.00861
R161 VDD1.n0 VDD1.t6 2.00861
R162 VDD1.n2 VDD1.t0 2.00861
R163 VDD1.n2 VDD1.t3 2.00861
R164 VDD1.n1 VDD1.t1 2.00861
R165 VDD1.n1 VDD1.t7 2.00861
R166 VDD1 VDD1.n5 1.41214
R167 B.n719 B.n718 585
R168 B.n721 B.n151 585
R169 B.n724 B.n723 585
R170 B.n725 B.n150 585
R171 B.n727 B.n726 585
R172 B.n729 B.n149 585
R173 B.n732 B.n731 585
R174 B.n733 B.n148 585
R175 B.n735 B.n734 585
R176 B.n737 B.n147 585
R177 B.n740 B.n739 585
R178 B.n741 B.n146 585
R179 B.n743 B.n742 585
R180 B.n745 B.n145 585
R181 B.n748 B.n747 585
R182 B.n749 B.n144 585
R183 B.n751 B.n750 585
R184 B.n753 B.n143 585
R185 B.n756 B.n755 585
R186 B.n757 B.n142 585
R187 B.n759 B.n758 585
R188 B.n761 B.n141 585
R189 B.n764 B.n763 585
R190 B.n765 B.n140 585
R191 B.n767 B.n766 585
R192 B.n769 B.n139 585
R193 B.n772 B.n771 585
R194 B.n773 B.n138 585
R195 B.n775 B.n774 585
R196 B.n777 B.n137 585
R197 B.n780 B.n779 585
R198 B.n781 B.n136 585
R199 B.n783 B.n782 585
R200 B.n785 B.n135 585
R201 B.n788 B.n787 585
R202 B.n790 B.n132 585
R203 B.n792 B.n791 585
R204 B.n794 B.n131 585
R205 B.n797 B.n796 585
R206 B.n798 B.n130 585
R207 B.n800 B.n799 585
R208 B.n802 B.n129 585
R209 B.n805 B.n804 585
R210 B.n806 B.n125 585
R211 B.n808 B.n807 585
R212 B.n810 B.n124 585
R213 B.n813 B.n812 585
R214 B.n814 B.n123 585
R215 B.n816 B.n815 585
R216 B.n818 B.n122 585
R217 B.n821 B.n820 585
R218 B.n822 B.n121 585
R219 B.n824 B.n823 585
R220 B.n826 B.n120 585
R221 B.n829 B.n828 585
R222 B.n830 B.n119 585
R223 B.n832 B.n831 585
R224 B.n834 B.n118 585
R225 B.n837 B.n836 585
R226 B.n838 B.n117 585
R227 B.n840 B.n839 585
R228 B.n842 B.n116 585
R229 B.n845 B.n844 585
R230 B.n846 B.n115 585
R231 B.n848 B.n847 585
R232 B.n850 B.n114 585
R233 B.n853 B.n852 585
R234 B.n854 B.n113 585
R235 B.n856 B.n855 585
R236 B.n858 B.n112 585
R237 B.n861 B.n860 585
R238 B.n862 B.n111 585
R239 B.n864 B.n863 585
R240 B.n866 B.n110 585
R241 B.n869 B.n868 585
R242 B.n870 B.n109 585
R243 B.n872 B.n871 585
R244 B.n874 B.n108 585
R245 B.n877 B.n876 585
R246 B.n878 B.n107 585
R247 B.n717 B.n105 585
R248 B.n881 B.n105 585
R249 B.n716 B.n104 585
R250 B.n882 B.n104 585
R251 B.n715 B.n103 585
R252 B.n883 B.n103 585
R253 B.n714 B.n713 585
R254 B.n713 B.n99 585
R255 B.n712 B.n98 585
R256 B.n889 B.n98 585
R257 B.n711 B.n97 585
R258 B.n890 B.n97 585
R259 B.n710 B.n96 585
R260 B.n891 B.n96 585
R261 B.n709 B.n708 585
R262 B.n708 B.n92 585
R263 B.n707 B.n91 585
R264 B.n897 B.n91 585
R265 B.n706 B.n90 585
R266 B.n898 B.n90 585
R267 B.n705 B.n89 585
R268 B.n899 B.n89 585
R269 B.n704 B.n703 585
R270 B.n703 B.n85 585
R271 B.n702 B.n84 585
R272 B.n905 B.n84 585
R273 B.n701 B.n83 585
R274 B.n906 B.n83 585
R275 B.n700 B.n82 585
R276 B.n907 B.n82 585
R277 B.n699 B.n698 585
R278 B.n698 B.n78 585
R279 B.n697 B.n77 585
R280 B.n913 B.n77 585
R281 B.n696 B.n76 585
R282 B.n914 B.n76 585
R283 B.n695 B.n75 585
R284 B.n915 B.n75 585
R285 B.n694 B.n693 585
R286 B.n693 B.n71 585
R287 B.n692 B.n70 585
R288 B.n921 B.n70 585
R289 B.n691 B.n69 585
R290 B.n922 B.n69 585
R291 B.n690 B.n68 585
R292 B.n923 B.n68 585
R293 B.n689 B.n688 585
R294 B.n688 B.n64 585
R295 B.n687 B.n63 585
R296 B.n929 B.n63 585
R297 B.n686 B.n62 585
R298 B.n930 B.n62 585
R299 B.n685 B.n61 585
R300 B.n931 B.n61 585
R301 B.n684 B.n683 585
R302 B.n683 B.n57 585
R303 B.n682 B.n56 585
R304 B.n937 B.n56 585
R305 B.n681 B.n55 585
R306 B.n938 B.n55 585
R307 B.n680 B.n54 585
R308 B.n939 B.n54 585
R309 B.n679 B.n678 585
R310 B.n678 B.n53 585
R311 B.n677 B.n49 585
R312 B.n945 B.n49 585
R313 B.n676 B.n48 585
R314 B.n946 B.n48 585
R315 B.n675 B.n47 585
R316 B.n947 B.n47 585
R317 B.n674 B.n673 585
R318 B.n673 B.n43 585
R319 B.n672 B.n42 585
R320 B.n953 B.n42 585
R321 B.n671 B.n41 585
R322 B.n954 B.n41 585
R323 B.n670 B.n40 585
R324 B.n955 B.n40 585
R325 B.n669 B.n668 585
R326 B.n668 B.n36 585
R327 B.n667 B.n35 585
R328 B.n961 B.n35 585
R329 B.n666 B.n34 585
R330 B.n962 B.n34 585
R331 B.n665 B.n33 585
R332 B.n963 B.n33 585
R333 B.n664 B.n663 585
R334 B.n663 B.n29 585
R335 B.n662 B.n28 585
R336 B.n969 B.n28 585
R337 B.n661 B.n27 585
R338 B.n970 B.n27 585
R339 B.n660 B.n26 585
R340 B.n971 B.n26 585
R341 B.n659 B.n658 585
R342 B.n658 B.n22 585
R343 B.n657 B.n21 585
R344 B.n977 B.n21 585
R345 B.n656 B.n20 585
R346 B.n978 B.n20 585
R347 B.n655 B.n19 585
R348 B.n979 B.n19 585
R349 B.n654 B.n653 585
R350 B.n653 B.n18 585
R351 B.n652 B.n14 585
R352 B.n985 B.n14 585
R353 B.n651 B.n13 585
R354 B.n986 B.n13 585
R355 B.n650 B.n12 585
R356 B.n987 B.n12 585
R357 B.n649 B.n648 585
R358 B.n648 B.n8 585
R359 B.n647 B.n7 585
R360 B.n993 B.n7 585
R361 B.n646 B.n6 585
R362 B.n994 B.n6 585
R363 B.n645 B.n5 585
R364 B.n995 B.n5 585
R365 B.n644 B.n643 585
R366 B.n643 B.n4 585
R367 B.n642 B.n152 585
R368 B.n642 B.n641 585
R369 B.n632 B.n153 585
R370 B.n154 B.n153 585
R371 B.n634 B.n633 585
R372 B.n635 B.n634 585
R373 B.n631 B.n159 585
R374 B.n159 B.n158 585
R375 B.n630 B.n629 585
R376 B.n629 B.n628 585
R377 B.n161 B.n160 585
R378 B.n621 B.n161 585
R379 B.n620 B.n619 585
R380 B.n622 B.n620 585
R381 B.n618 B.n166 585
R382 B.n166 B.n165 585
R383 B.n617 B.n616 585
R384 B.n616 B.n615 585
R385 B.n168 B.n167 585
R386 B.n169 B.n168 585
R387 B.n608 B.n607 585
R388 B.n609 B.n608 585
R389 B.n606 B.n174 585
R390 B.n174 B.n173 585
R391 B.n605 B.n604 585
R392 B.n604 B.n603 585
R393 B.n176 B.n175 585
R394 B.n177 B.n176 585
R395 B.n596 B.n595 585
R396 B.n597 B.n596 585
R397 B.n594 B.n181 585
R398 B.n185 B.n181 585
R399 B.n593 B.n592 585
R400 B.n592 B.n591 585
R401 B.n183 B.n182 585
R402 B.n184 B.n183 585
R403 B.n584 B.n583 585
R404 B.n585 B.n584 585
R405 B.n582 B.n190 585
R406 B.n190 B.n189 585
R407 B.n581 B.n580 585
R408 B.n580 B.n579 585
R409 B.n192 B.n191 585
R410 B.n193 B.n192 585
R411 B.n572 B.n571 585
R412 B.n573 B.n572 585
R413 B.n570 B.n198 585
R414 B.n198 B.n197 585
R415 B.n569 B.n568 585
R416 B.n568 B.n567 585
R417 B.n200 B.n199 585
R418 B.n560 B.n200 585
R419 B.n559 B.n558 585
R420 B.n561 B.n559 585
R421 B.n557 B.n205 585
R422 B.n205 B.n204 585
R423 B.n556 B.n555 585
R424 B.n555 B.n554 585
R425 B.n207 B.n206 585
R426 B.n208 B.n207 585
R427 B.n547 B.n546 585
R428 B.n548 B.n547 585
R429 B.n545 B.n213 585
R430 B.n213 B.n212 585
R431 B.n544 B.n543 585
R432 B.n543 B.n542 585
R433 B.n215 B.n214 585
R434 B.n216 B.n215 585
R435 B.n535 B.n534 585
R436 B.n536 B.n535 585
R437 B.n533 B.n220 585
R438 B.n224 B.n220 585
R439 B.n532 B.n531 585
R440 B.n531 B.n530 585
R441 B.n222 B.n221 585
R442 B.n223 B.n222 585
R443 B.n523 B.n522 585
R444 B.n524 B.n523 585
R445 B.n521 B.n229 585
R446 B.n229 B.n228 585
R447 B.n520 B.n519 585
R448 B.n519 B.n518 585
R449 B.n231 B.n230 585
R450 B.n232 B.n231 585
R451 B.n511 B.n510 585
R452 B.n512 B.n511 585
R453 B.n509 B.n237 585
R454 B.n237 B.n236 585
R455 B.n508 B.n507 585
R456 B.n507 B.n506 585
R457 B.n239 B.n238 585
R458 B.n240 B.n239 585
R459 B.n499 B.n498 585
R460 B.n500 B.n499 585
R461 B.n497 B.n245 585
R462 B.n245 B.n244 585
R463 B.n496 B.n495 585
R464 B.n495 B.n494 585
R465 B.n247 B.n246 585
R466 B.n248 B.n247 585
R467 B.n487 B.n486 585
R468 B.n488 B.n487 585
R469 B.n485 B.n253 585
R470 B.n253 B.n252 585
R471 B.n484 B.n483 585
R472 B.n483 B.n482 585
R473 B.n255 B.n254 585
R474 B.n256 B.n255 585
R475 B.n475 B.n474 585
R476 B.n476 B.n475 585
R477 B.n473 B.n261 585
R478 B.n261 B.n260 585
R479 B.n472 B.n471 585
R480 B.n471 B.n470 585
R481 B.n467 B.n265 585
R482 B.n466 B.n465 585
R483 B.n463 B.n266 585
R484 B.n463 B.n264 585
R485 B.n462 B.n461 585
R486 B.n460 B.n459 585
R487 B.n458 B.n268 585
R488 B.n456 B.n455 585
R489 B.n454 B.n269 585
R490 B.n453 B.n452 585
R491 B.n450 B.n270 585
R492 B.n448 B.n447 585
R493 B.n446 B.n271 585
R494 B.n445 B.n444 585
R495 B.n442 B.n272 585
R496 B.n440 B.n439 585
R497 B.n438 B.n273 585
R498 B.n437 B.n436 585
R499 B.n434 B.n274 585
R500 B.n432 B.n431 585
R501 B.n430 B.n275 585
R502 B.n429 B.n428 585
R503 B.n426 B.n276 585
R504 B.n424 B.n423 585
R505 B.n422 B.n277 585
R506 B.n421 B.n420 585
R507 B.n418 B.n278 585
R508 B.n416 B.n415 585
R509 B.n414 B.n279 585
R510 B.n413 B.n412 585
R511 B.n410 B.n280 585
R512 B.n408 B.n407 585
R513 B.n406 B.n281 585
R514 B.n405 B.n404 585
R515 B.n402 B.n282 585
R516 B.n400 B.n399 585
R517 B.n397 B.n283 585
R518 B.n396 B.n395 585
R519 B.n393 B.n286 585
R520 B.n391 B.n390 585
R521 B.n389 B.n287 585
R522 B.n388 B.n387 585
R523 B.n385 B.n288 585
R524 B.n383 B.n382 585
R525 B.n381 B.n289 585
R526 B.n380 B.n379 585
R527 B.n377 B.n376 585
R528 B.n375 B.n374 585
R529 B.n373 B.n294 585
R530 B.n371 B.n370 585
R531 B.n369 B.n295 585
R532 B.n368 B.n367 585
R533 B.n365 B.n296 585
R534 B.n363 B.n362 585
R535 B.n361 B.n297 585
R536 B.n360 B.n359 585
R537 B.n357 B.n298 585
R538 B.n355 B.n354 585
R539 B.n353 B.n299 585
R540 B.n352 B.n351 585
R541 B.n349 B.n300 585
R542 B.n347 B.n346 585
R543 B.n345 B.n301 585
R544 B.n344 B.n343 585
R545 B.n341 B.n302 585
R546 B.n339 B.n338 585
R547 B.n337 B.n303 585
R548 B.n336 B.n335 585
R549 B.n333 B.n304 585
R550 B.n331 B.n330 585
R551 B.n329 B.n305 585
R552 B.n328 B.n327 585
R553 B.n325 B.n306 585
R554 B.n323 B.n322 585
R555 B.n321 B.n307 585
R556 B.n320 B.n319 585
R557 B.n317 B.n308 585
R558 B.n315 B.n314 585
R559 B.n313 B.n309 585
R560 B.n312 B.n311 585
R561 B.n263 B.n262 585
R562 B.n264 B.n263 585
R563 B.n469 B.n468 585
R564 B.n470 B.n469 585
R565 B.n259 B.n258 585
R566 B.n260 B.n259 585
R567 B.n478 B.n477 585
R568 B.n477 B.n476 585
R569 B.n479 B.n257 585
R570 B.n257 B.n256 585
R571 B.n481 B.n480 585
R572 B.n482 B.n481 585
R573 B.n251 B.n250 585
R574 B.n252 B.n251 585
R575 B.n490 B.n489 585
R576 B.n489 B.n488 585
R577 B.n491 B.n249 585
R578 B.n249 B.n248 585
R579 B.n493 B.n492 585
R580 B.n494 B.n493 585
R581 B.n243 B.n242 585
R582 B.n244 B.n243 585
R583 B.n502 B.n501 585
R584 B.n501 B.n500 585
R585 B.n503 B.n241 585
R586 B.n241 B.n240 585
R587 B.n505 B.n504 585
R588 B.n506 B.n505 585
R589 B.n235 B.n234 585
R590 B.n236 B.n235 585
R591 B.n514 B.n513 585
R592 B.n513 B.n512 585
R593 B.n515 B.n233 585
R594 B.n233 B.n232 585
R595 B.n517 B.n516 585
R596 B.n518 B.n517 585
R597 B.n227 B.n226 585
R598 B.n228 B.n227 585
R599 B.n526 B.n525 585
R600 B.n525 B.n524 585
R601 B.n527 B.n225 585
R602 B.n225 B.n223 585
R603 B.n529 B.n528 585
R604 B.n530 B.n529 585
R605 B.n219 B.n218 585
R606 B.n224 B.n219 585
R607 B.n538 B.n537 585
R608 B.n537 B.n536 585
R609 B.n539 B.n217 585
R610 B.n217 B.n216 585
R611 B.n541 B.n540 585
R612 B.n542 B.n541 585
R613 B.n211 B.n210 585
R614 B.n212 B.n211 585
R615 B.n550 B.n549 585
R616 B.n549 B.n548 585
R617 B.n551 B.n209 585
R618 B.n209 B.n208 585
R619 B.n553 B.n552 585
R620 B.n554 B.n553 585
R621 B.n203 B.n202 585
R622 B.n204 B.n203 585
R623 B.n563 B.n562 585
R624 B.n562 B.n561 585
R625 B.n564 B.n201 585
R626 B.n560 B.n201 585
R627 B.n566 B.n565 585
R628 B.n567 B.n566 585
R629 B.n196 B.n195 585
R630 B.n197 B.n196 585
R631 B.n575 B.n574 585
R632 B.n574 B.n573 585
R633 B.n576 B.n194 585
R634 B.n194 B.n193 585
R635 B.n578 B.n577 585
R636 B.n579 B.n578 585
R637 B.n188 B.n187 585
R638 B.n189 B.n188 585
R639 B.n587 B.n586 585
R640 B.n586 B.n585 585
R641 B.n588 B.n186 585
R642 B.n186 B.n184 585
R643 B.n590 B.n589 585
R644 B.n591 B.n590 585
R645 B.n180 B.n179 585
R646 B.n185 B.n180 585
R647 B.n599 B.n598 585
R648 B.n598 B.n597 585
R649 B.n600 B.n178 585
R650 B.n178 B.n177 585
R651 B.n602 B.n601 585
R652 B.n603 B.n602 585
R653 B.n172 B.n171 585
R654 B.n173 B.n172 585
R655 B.n611 B.n610 585
R656 B.n610 B.n609 585
R657 B.n612 B.n170 585
R658 B.n170 B.n169 585
R659 B.n614 B.n613 585
R660 B.n615 B.n614 585
R661 B.n164 B.n163 585
R662 B.n165 B.n164 585
R663 B.n624 B.n623 585
R664 B.n623 B.n622 585
R665 B.n625 B.n162 585
R666 B.n621 B.n162 585
R667 B.n627 B.n626 585
R668 B.n628 B.n627 585
R669 B.n157 B.n156 585
R670 B.n158 B.n157 585
R671 B.n637 B.n636 585
R672 B.n636 B.n635 585
R673 B.n638 B.n155 585
R674 B.n155 B.n154 585
R675 B.n640 B.n639 585
R676 B.n641 B.n640 585
R677 B.n2 B.n0 585
R678 B.n4 B.n2 585
R679 B.n3 B.n1 585
R680 B.n994 B.n3 585
R681 B.n992 B.n991 585
R682 B.n993 B.n992 585
R683 B.n990 B.n9 585
R684 B.n9 B.n8 585
R685 B.n989 B.n988 585
R686 B.n988 B.n987 585
R687 B.n11 B.n10 585
R688 B.n986 B.n11 585
R689 B.n984 B.n983 585
R690 B.n985 B.n984 585
R691 B.n982 B.n15 585
R692 B.n18 B.n15 585
R693 B.n981 B.n980 585
R694 B.n980 B.n979 585
R695 B.n17 B.n16 585
R696 B.n978 B.n17 585
R697 B.n976 B.n975 585
R698 B.n977 B.n976 585
R699 B.n974 B.n23 585
R700 B.n23 B.n22 585
R701 B.n973 B.n972 585
R702 B.n972 B.n971 585
R703 B.n25 B.n24 585
R704 B.n970 B.n25 585
R705 B.n968 B.n967 585
R706 B.n969 B.n968 585
R707 B.n966 B.n30 585
R708 B.n30 B.n29 585
R709 B.n965 B.n964 585
R710 B.n964 B.n963 585
R711 B.n32 B.n31 585
R712 B.n962 B.n32 585
R713 B.n960 B.n959 585
R714 B.n961 B.n960 585
R715 B.n958 B.n37 585
R716 B.n37 B.n36 585
R717 B.n957 B.n956 585
R718 B.n956 B.n955 585
R719 B.n39 B.n38 585
R720 B.n954 B.n39 585
R721 B.n952 B.n951 585
R722 B.n953 B.n952 585
R723 B.n950 B.n44 585
R724 B.n44 B.n43 585
R725 B.n949 B.n948 585
R726 B.n948 B.n947 585
R727 B.n46 B.n45 585
R728 B.n946 B.n46 585
R729 B.n944 B.n943 585
R730 B.n945 B.n944 585
R731 B.n942 B.n50 585
R732 B.n53 B.n50 585
R733 B.n941 B.n940 585
R734 B.n940 B.n939 585
R735 B.n52 B.n51 585
R736 B.n938 B.n52 585
R737 B.n936 B.n935 585
R738 B.n937 B.n936 585
R739 B.n934 B.n58 585
R740 B.n58 B.n57 585
R741 B.n933 B.n932 585
R742 B.n932 B.n931 585
R743 B.n60 B.n59 585
R744 B.n930 B.n60 585
R745 B.n928 B.n927 585
R746 B.n929 B.n928 585
R747 B.n926 B.n65 585
R748 B.n65 B.n64 585
R749 B.n925 B.n924 585
R750 B.n924 B.n923 585
R751 B.n67 B.n66 585
R752 B.n922 B.n67 585
R753 B.n920 B.n919 585
R754 B.n921 B.n920 585
R755 B.n918 B.n72 585
R756 B.n72 B.n71 585
R757 B.n917 B.n916 585
R758 B.n916 B.n915 585
R759 B.n74 B.n73 585
R760 B.n914 B.n74 585
R761 B.n912 B.n911 585
R762 B.n913 B.n912 585
R763 B.n910 B.n79 585
R764 B.n79 B.n78 585
R765 B.n909 B.n908 585
R766 B.n908 B.n907 585
R767 B.n81 B.n80 585
R768 B.n906 B.n81 585
R769 B.n904 B.n903 585
R770 B.n905 B.n904 585
R771 B.n902 B.n86 585
R772 B.n86 B.n85 585
R773 B.n901 B.n900 585
R774 B.n900 B.n899 585
R775 B.n88 B.n87 585
R776 B.n898 B.n88 585
R777 B.n896 B.n895 585
R778 B.n897 B.n896 585
R779 B.n894 B.n93 585
R780 B.n93 B.n92 585
R781 B.n893 B.n892 585
R782 B.n892 B.n891 585
R783 B.n95 B.n94 585
R784 B.n890 B.n95 585
R785 B.n888 B.n887 585
R786 B.n889 B.n888 585
R787 B.n886 B.n100 585
R788 B.n100 B.n99 585
R789 B.n885 B.n884 585
R790 B.n884 B.n883 585
R791 B.n102 B.n101 585
R792 B.n882 B.n102 585
R793 B.n880 B.n879 585
R794 B.n881 B.n880 585
R795 B.n997 B.n996 585
R796 B.n996 B.n995 585
R797 B.n469 B.n265 559.769
R798 B.n880 B.n107 559.769
R799 B.n471 B.n263 559.769
R800 B.n719 B.n105 559.769
R801 B.n290 B.t8 285.824
R802 B.n284 B.t16 285.824
R803 B.n126 B.t19 285.824
R804 B.n133 B.t12 285.824
R805 B.n720 B.n106 256.663
R806 B.n722 B.n106 256.663
R807 B.n728 B.n106 256.663
R808 B.n730 B.n106 256.663
R809 B.n736 B.n106 256.663
R810 B.n738 B.n106 256.663
R811 B.n744 B.n106 256.663
R812 B.n746 B.n106 256.663
R813 B.n752 B.n106 256.663
R814 B.n754 B.n106 256.663
R815 B.n760 B.n106 256.663
R816 B.n762 B.n106 256.663
R817 B.n768 B.n106 256.663
R818 B.n770 B.n106 256.663
R819 B.n776 B.n106 256.663
R820 B.n778 B.n106 256.663
R821 B.n784 B.n106 256.663
R822 B.n786 B.n106 256.663
R823 B.n793 B.n106 256.663
R824 B.n795 B.n106 256.663
R825 B.n801 B.n106 256.663
R826 B.n803 B.n106 256.663
R827 B.n809 B.n106 256.663
R828 B.n811 B.n106 256.663
R829 B.n817 B.n106 256.663
R830 B.n819 B.n106 256.663
R831 B.n825 B.n106 256.663
R832 B.n827 B.n106 256.663
R833 B.n833 B.n106 256.663
R834 B.n835 B.n106 256.663
R835 B.n841 B.n106 256.663
R836 B.n843 B.n106 256.663
R837 B.n849 B.n106 256.663
R838 B.n851 B.n106 256.663
R839 B.n857 B.n106 256.663
R840 B.n859 B.n106 256.663
R841 B.n865 B.n106 256.663
R842 B.n867 B.n106 256.663
R843 B.n873 B.n106 256.663
R844 B.n875 B.n106 256.663
R845 B.n464 B.n264 256.663
R846 B.n267 B.n264 256.663
R847 B.n457 B.n264 256.663
R848 B.n451 B.n264 256.663
R849 B.n449 B.n264 256.663
R850 B.n443 B.n264 256.663
R851 B.n441 B.n264 256.663
R852 B.n435 B.n264 256.663
R853 B.n433 B.n264 256.663
R854 B.n427 B.n264 256.663
R855 B.n425 B.n264 256.663
R856 B.n419 B.n264 256.663
R857 B.n417 B.n264 256.663
R858 B.n411 B.n264 256.663
R859 B.n409 B.n264 256.663
R860 B.n403 B.n264 256.663
R861 B.n401 B.n264 256.663
R862 B.n394 B.n264 256.663
R863 B.n392 B.n264 256.663
R864 B.n386 B.n264 256.663
R865 B.n384 B.n264 256.663
R866 B.n378 B.n264 256.663
R867 B.n293 B.n264 256.663
R868 B.n372 B.n264 256.663
R869 B.n366 B.n264 256.663
R870 B.n364 B.n264 256.663
R871 B.n358 B.n264 256.663
R872 B.n356 B.n264 256.663
R873 B.n350 B.n264 256.663
R874 B.n348 B.n264 256.663
R875 B.n342 B.n264 256.663
R876 B.n340 B.n264 256.663
R877 B.n334 B.n264 256.663
R878 B.n332 B.n264 256.663
R879 B.n326 B.n264 256.663
R880 B.n324 B.n264 256.663
R881 B.n318 B.n264 256.663
R882 B.n316 B.n264 256.663
R883 B.n310 B.n264 256.663
R884 B.n469 B.n259 163.367
R885 B.n477 B.n259 163.367
R886 B.n477 B.n257 163.367
R887 B.n481 B.n257 163.367
R888 B.n481 B.n251 163.367
R889 B.n489 B.n251 163.367
R890 B.n489 B.n249 163.367
R891 B.n493 B.n249 163.367
R892 B.n493 B.n243 163.367
R893 B.n501 B.n243 163.367
R894 B.n501 B.n241 163.367
R895 B.n505 B.n241 163.367
R896 B.n505 B.n235 163.367
R897 B.n513 B.n235 163.367
R898 B.n513 B.n233 163.367
R899 B.n517 B.n233 163.367
R900 B.n517 B.n227 163.367
R901 B.n525 B.n227 163.367
R902 B.n525 B.n225 163.367
R903 B.n529 B.n225 163.367
R904 B.n529 B.n219 163.367
R905 B.n537 B.n219 163.367
R906 B.n537 B.n217 163.367
R907 B.n541 B.n217 163.367
R908 B.n541 B.n211 163.367
R909 B.n549 B.n211 163.367
R910 B.n549 B.n209 163.367
R911 B.n553 B.n209 163.367
R912 B.n553 B.n203 163.367
R913 B.n562 B.n203 163.367
R914 B.n562 B.n201 163.367
R915 B.n566 B.n201 163.367
R916 B.n566 B.n196 163.367
R917 B.n574 B.n196 163.367
R918 B.n574 B.n194 163.367
R919 B.n578 B.n194 163.367
R920 B.n578 B.n188 163.367
R921 B.n586 B.n188 163.367
R922 B.n586 B.n186 163.367
R923 B.n590 B.n186 163.367
R924 B.n590 B.n180 163.367
R925 B.n598 B.n180 163.367
R926 B.n598 B.n178 163.367
R927 B.n602 B.n178 163.367
R928 B.n602 B.n172 163.367
R929 B.n610 B.n172 163.367
R930 B.n610 B.n170 163.367
R931 B.n614 B.n170 163.367
R932 B.n614 B.n164 163.367
R933 B.n623 B.n164 163.367
R934 B.n623 B.n162 163.367
R935 B.n627 B.n162 163.367
R936 B.n627 B.n157 163.367
R937 B.n636 B.n157 163.367
R938 B.n636 B.n155 163.367
R939 B.n640 B.n155 163.367
R940 B.n640 B.n2 163.367
R941 B.n996 B.n2 163.367
R942 B.n996 B.n3 163.367
R943 B.n992 B.n3 163.367
R944 B.n992 B.n9 163.367
R945 B.n988 B.n9 163.367
R946 B.n988 B.n11 163.367
R947 B.n984 B.n11 163.367
R948 B.n984 B.n15 163.367
R949 B.n980 B.n15 163.367
R950 B.n980 B.n17 163.367
R951 B.n976 B.n17 163.367
R952 B.n976 B.n23 163.367
R953 B.n972 B.n23 163.367
R954 B.n972 B.n25 163.367
R955 B.n968 B.n25 163.367
R956 B.n968 B.n30 163.367
R957 B.n964 B.n30 163.367
R958 B.n964 B.n32 163.367
R959 B.n960 B.n32 163.367
R960 B.n960 B.n37 163.367
R961 B.n956 B.n37 163.367
R962 B.n956 B.n39 163.367
R963 B.n952 B.n39 163.367
R964 B.n952 B.n44 163.367
R965 B.n948 B.n44 163.367
R966 B.n948 B.n46 163.367
R967 B.n944 B.n46 163.367
R968 B.n944 B.n50 163.367
R969 B.n940 B.n50 163.367
R970 B.n940 B.n52 163.367
R971 B.n936 B.n52 163.367
R972 B.n936 B.n58 163.367
R973 B.n932 B.n58 163.367
R974 B.n932 B.n60 163.367
R975 B.n928 B.n60 163.367
R976 B.n928 B.n65 163.367
R977 B.n924 B.n65 163.367
R978 B.n924 B.n67 163.367
R979 B.n920 B.n67 163.367
R980 B.n920 B.n72 163.367
R981 B.n916 B.n72 163.367
R982 B.n916 B.n74 163.367
R983 B.n912 B.n74 163.367
R984 B.n912 B.n79 163.367
R985 B.n908 B.n79 163.367
R986 B.n908 B.n81 163.367
R987 B.n904 B.n81 163.367
R988 B.n904 B.n86 163.367
R989 B.n900 B.n86 163.367
R990 B.n900 B.n88 163.367
R991 B.n896 B.n88 163.367
R992 B.n896 B.n93 163.367
R993 B.n892 B.n93 163.367
R994 B.n892 B.n95 163.367
R995 B.n888 B.n95 163.367
R996 B.n888 B.n100 163.367
R997 B.n884 B.n100 163.367
R998 B.n884 B.n102 163.367
R999 B.n880 B.n102 163.367
R1000 B.n465 B.n463 163.367
R1001 B.n463 B.n462 163.367
R1002 B.n459 B.n458 163.367
R1003 B.n456 B.n269 163.367
R1004 B.n452 B.n450 163.367
R1005 B.n448 B.n271 163.367
R1006 B.n444 B.n442 163.367
R1007 B.n440 B.n273 163.367
R1008 B.n436 B.n434 163.367
R1009 B.n432 B.n275 163.367
R1010 B.n428 B.n426 163.367
R1011 B.n424 B.n277 163.367
R1012 B.n420 B.n418 163.367
R1013 B.n416 B.n279 163.367
R1014 B.n412 B.n410 163.367
R1015 B.n408 B.n281 163.367
R1016 B.n404 B.n402 163.367
R1017 B.n400 B.n283 163.367
R1018 B.n395 B.n393 163.367
R1019 B.n391 B.n287 163.367
R1020 B.n387 B.n385 163.367
R1021 B.n383 B.n289 163.367
R1022 B.n379 B.n377 163.367
R1023 B.n374 B.n373 163.367
R1024 B.n371 B.n295 163.367
R1025 B.n367 B.n365 163.367
R1026 B.n363 B.n297 163.367
R1027 B.n359 B.n357 163.367
R1028 B.n355 B.n299 163.367
R1029 B.n351 B.n349 163.367
R1030 B.n347 B.n301 163.367
R1031 B.n343 B.n341 163.367
R1032 B.n339 B.n303 163.367
R1033 B.n335 B.n333 163.367
R1034 B.n331 B.n305 163.367
R1035 B.n327 B.n325 163.367
R1036 B.n323 B.n307 163.367
R1037 B.n319 B.n317 163.367
R1038 B.n315 B.n309 163.367
R1039 B.n311 B.n263 163.367
R1040 B.n471 B.n261 163.367
R1041 B.n475 B.n261 163.367
R1042 B.n475 B.n255 163.367
R1043 B.n483 B.n255 163.367
R1044 B.n483 B.n253 163.367
R1045 B.n487 B.n253 163.367
R1046 B.n487 B.n247 163.367
R1047 B.n495 B.n247 163.367
R1048 B.n495 B.n245 163.367
R1049 B.n499 B.n245 163.367
R1050 B.n499 B.n239 163.367
R1051 B.n507 B.n239 163.367
R1052 B.n507 B.n237 163.367
R1053 B.n511 B.n237 163.367
R1054 B.n511 B.n231 163.367
R1055 B.n519 B.n231 163.367
R1056 B.n519 B.n229 163.367
R1057 B.n523 B.n229 163.367
R1058 B.n523 B.n222 163.367
R1059 B.n531 B.n222 163.367
R1060 B.n531 B.n220 163.367
R1061 B.n535 B.n220 163.367
R1062 B.n535 B.n215 163.367
R1063 B.n543 B.n215 163.367
R1064 B.n543 B.n213 163.367
R1065 B.n547 B.n213 163.367
R1066 B.n547 B.n207 163.367
R1067 B.n555 B.n207 163.367
R1068 B.n555 B.n205 163.367
R1069 B.n559 B.n205 163.367
R1070 B.n559 B.n200 163.367
R1071 B.n568 B.n200 163.367
R1072 B.n568 B.n198 163.367
R1073 B.n572 B.n198 163.367
R1074 B.n572 B.n192 163.367
R1075 B.n580 B.n192 163.367
R1076 B.n580 B.n190 163.367
R1077 B.n584 B.n190 163.367
R1078 B.n584 B.n183 163.367
R1079 B.n592 B.n183 163.367
R1080 B.n592 B.n181 163.367
R1081 B.n596 B.n181 163.367
R1082 B.n596 B.n176 163.367
R1083 B.n604 B.n176 163.367
R1084 B.n604 B.n174 163.367
R1085 B.n608 B.n174 163.367
R1086 B.n608 B.n168 163.367
R1087 B.n616 B.n168 163.367
R1088 B.n616 B.n166 163.367
R1089 B.n620 B.n166 163.367
R1090 B.n620 B.n161 163.367
R1091 B.n629 B.n161 163.367
R1092 B.n629 B.n159 163.367
R1093 B.n634 B.n159 163.367
R1094 B.n634 B.n153 163.367
R1095 B.n642 B.n153 163.367
R1096 B.n643 B.n642 163.367
R1097 B.n643 B.n5 163.367
R1098 B.n6 B.n5 163.367
R1099 B.n7 B.n6 163.367
R1100 B.n648 B.n7 163.367
R1101 B.n648 B.n12 163.367
R1102 B.n13 B.n12 163.367
R1103 B.n14 B.n13 163.367
R1104 B.n653 B.n14 163.367
R1105 B.n653 B.n19 163.367
R1106 B.n20 B.n19 163.367
R1107 B.n21 B.n20 163.367
R1108 B.n658 B.n21 163.367
R1109 B.n658 B.n26 163.367
R1110 B.n27 B.n26 163.367
R1111 B.n28 B.n27 163.367
R1112 B.n663 B.n28 163.367
R1113 B.n663 B.n33 163.367
R1114 B.n34 B.n33 163.367
R1115 B.n35 B.n34 163.367
R1116 B.n668 B.n35 163.367
R1117 B.n668 B.n40 163.367
R1118 B.n41 B.n40 163.367
R1119 B.n42 B.n41 163.367
R1120 B.n673 B.n42 163.367
R1121 B.n673 B.n47 163.367
R1122 B.n48 B.n47 163.367
R1123 B.n49 B.n48 163.367
R1124 B.n678 B.n49 163.367
R1125 B.n678 B.n54 163.367
R1126 B.n55 B.n54 163.367
R1127 B.n56 B.n55 163.367
R1128 B.n683 B.n56 163.367
R1129 B.n683 B.n61 163.367
R1130 B.n62 B.n61 163.367
R1131 B.n63 B.n62 163.367
R1132 B.n688 B.n63 163.367
R1133 B.n688 B.n68 163.367
R1134 B.n69 B.n68 163.367
R1135 B.n70 B.n69 163.367
R1136 B.n693 B.n70 163.367
R1137 B.n693 B.n75 163.367
R1138 B.n76 B.n75 163.367
R1139 B.n77 B.n76 163.367
R1140 B.n698 B.n77 163.367
R1141 B.n698 B.n82 163.367
R1142 B.n83 B.n82 163.367
R1143 B.n84 B.n83 163.367
R1144 B.n703 B.n84 163.367
R1145 B.n703 B.n89 163.367
R1146 B.n90 B.n89 163.367
R1147 B.n91 B.n90 163.367
R1148 B.n708 B.n91 163.367
R1149 B.n708 B.n96 163.367
R1150 B.n97 B.n96 163.367
R1151 B.n98 B.n97 163.367
R1152 B.n713 B.n98 163.367
R1153 B.n713 B.n103 163.367
R1154 B.n104 B.n103 163.367
R1155 B.n105 B.n104 163.367
R1156 B.n876 B.n874 163.367
R1157 B.n872 B.n109 163.367
R1158 B.n868 B.n866 163.367
R1159 B.n864 B.n111 163.367
R1160 B.n860 B.n858 163.367
R1161 B.n856 B.n113 163.367
R1162 B.n852 B.n850 163.367
R1163 B.n848 B.n115 163.367
R1164 B.n844 B.n842 163.367
R1165 B.n840 B.n117 163.367
R1166 B.n836 B.n834 163.367
R1167 B.n832 B.n119 163.367
R1168 B.n828 B.n826 163.367
R1169 B.n824 B.n121 163.367
R1170 B.n820 B.n818 163.367
R1171 B.n816 B.n123 163.367
R1172 B.n812 B.n810 163.367
R1173 B.n808 B.n125 163.367
R1174 B.n804 B.n802 163.367
R1175 B.n800 B.n130 163.367
R1176 B.n796 B.n794 163.367
R1177 B.n792 B.n132 163.367
R1178 B.n787 B.n785 163.367
R1179 B.n783 B.n136 163.367
R1180 B.n779 B.n777 163.367
R1181 B.n775 B.n138 163.367
R1182 B.n771 B.n769 163.367
R1183 B.n767 B.n140 163.367
R1184 B.n763 B.n761 163.367
R1185 B.n759 B.n142 163.367
R1186 B.n755 B.n753 163.367
R1187 B.n751 B.n144 163.367
R1188 B.n747 B.n745 163.367
R1189 B.n743 B.n146 163.367
R1190 B.n739 B.n737 163.367
R1191 B.n735 B.n148 163.367
R1192 B.n731 B.n729 163.367
R1193 B.n727 B.n150 163.367
R1194 B.n723 B.n721 163.367
R1195 B.n290 B.t11 140.871
R1196 B.n133 B.t14 140.871
R1197 B.n284 B.t18 140.861
R1198 B.n126 B.t20 140.861
R1199 B.n470 B.n264 102.478
R1200 B.n881 B.n106 102.478
R1201 B.n291 B.t10 74.7385
R1202 B.n134 B.t15 74.7385
R1203 B.n285 B.t17 74.7268
R1204 B.n127 B.t21 74.7268
R1205 B.n464 B.n265 71.676
R1206 B.n462 B.n267 71.676
R1207 B.n458 B.n457 71.676
R1208 B.n451 B.n269 71.676
R1209 B.n450 B.n449 71.676
R1210 B.n443 B.n271 71.676
R1211 B.n442 B.n441 71.676
R1212 B.n435 B.n273 71.676
R1213 B.n434 B.n433 71.676
R1214 B.n427 B.n275 71.676
R1215 B.n426 B.n425 71.676
R1216 B.n419 B.n277 71.676
R1217 B.n418 B.n417 71.676
R1218 B.n411 B.n279 71.676
R1219 B.n410 B.n409 71.676
R1220 B.n403 B.n281 71.676
R1221 B.n402 B.n401 71.676
R1222 B.n394 B.n283 71.676
R1223 B.n393 B.n392 71.676
R1224 B.n386 B.n287 71.676
R1225 B.n385 B.n384 71.676
R1226 B.n378 B.n289 71.676
R1227 B.n377 B.n293 71.676
R1228 B.n373 B.n372 71.676
R1229 B.n366 B.n295 71.676
R1230 B.n365 B.n364 71.676
R1231 B.n358 B.n297 71.676
R1232 B.n357 B.n356 71.676
R1233 B.n350 B.n299 71.676
R1234 B.n349 B.n348 71.676
R1235 B.n342 B.n301 71.676
R1236 B.n341 B.n340 71.676
R1237 B.n334 B.n303 71.676
R1238 B.n333 B.n332 71.676
R1239 B.n326 B.n305 71.676
R1240 B.n325 B.n324 71.676
R1241 B.n318 B.n307 71.676
R1242 B.n317 B.n316 71.676
R1243 B.n310 B.n309 71.676
R1244 B.n875 B.n107 71.676
R1245 B.n874 B.n873 71.676
R1246 B.n867 B.n109 71.676
R1247 B.n866 B.n865 71.676
R1248 B.n859 B.n111 71.676
R1249 B.n858 B.n857 71.676
R1250 B.n851 B.n113 71.676
R1251 B.n850 B.n849 71.676
R1252 B.n843 B.n115 71.676
R1253 B.n842 B.n841 71.676
R1254 B.n835 B.n117 71.676
R1255 B.n834 B.n833 71.676
R1256 B.n827 B.n119 71.676
R1257 B.n826 B.n825 71.676
R1258 B.n819 B.n121 71.676
R1259 B.n818 B.n817 71.676
R1260 B.n811 B.n123 71.676
R1261 B.n810 B.n809 71.676
R1262 B.n803 B.n125 71.676
R1263 B.n802 B.n801 71.676
R1264 B.n795 B.n130 71.676
R1265 B.n794 B.n793 71.676
R1266 B.n786 B.n132 71.676
R1267 B.n785 B.n784 71.676
R1268 B.n778 B.n136 71.676
R1269 B.n777 B.n776 71.676
R1270 B.n770 B.n138 71.676
R1271 B.n769 B.n768 71.676
R1272 B.n762 B.n140 71.676
R1273 B.n761 B.n760 71.676
R1274 B.n754 B.n142 71.676
R1275 B.n753 B.n752 71.676
R1276 B.n746 B.n144 71.676
R1277 B.n745 B.n744 71.676
R1278 B.n738 B.n146 71.676
R1279 B.n737 B.n736 71.676
R1280 B.n730 B.n148 71.676
R1281 B.n729 B.n728 71.676
R1282 B.n722 B.n150 71.676
R1283 B.n721 B.n720 71.676
R1284 B.n720 B.n719 71.676
R1285 B.n723 B.n722 71.676
R1286 B.n728 B.n727 71.676
R1287 B.n731 B.n730 71.676
R1288 B.n736 B.n735 71.676
R1289 B.n739 B.n738 71.676
R1290 B.n744 B.n743 71.676
R1291 B.n747 B.n746 71.676
R1292 B.n752 B.n751 71.676
R1293 B.n755 B.n754 71.676
R1294 B.n760 B.n759 71.676
R1295 B.n763 B.n762 71.676
R1296 B.n768 B.n767 71.676
R1297 B.n771 B.n770 71.676
R1298 B.n776 B.n775 71.676
R1299 B.n779 B.n778 71.676
R1300 B.n784 B.n783 71.676
R1301 B.n787 B.n786 71.676
R1302 B.n793 B.n792 71.676
R1303 B.n796 B.n795 71.676
R1304 B.n801 B.n800 71.676
R1305 B.n804 B.n803 71.676
R1306 B.n809 B.n808 71.676
R1307 B.n812 B.n811 71.676
R1308 B.n817 B.n816 71.676
R1309 B.n820 B.n819 71.676
R1310 B.n825 B.n824 71.676
R1311 B.n828 B.n827 71.676
R1312 B.n833 B.n832 71.676
R1313 B.n836 B.n835 71.676
R1314 B.n841 B.n840 71.676
R1315 B.n844 B.n843 71.676
R1316 B.n849 B.n848 71.676
R1317 B.n852 B.n851 71.676
R1318 B.n857 B.n856 71.676
R1319 B.n860 B.n859 71.676
R1320 B.n865 B.n864 71.676
R1321 B.n868 B.n867 71.676
R1322 B.n873 B.n872 71.676
R1323 B.n876 B.n875 71.676
R1324 B.n465 B.n464 71.676
R1325 B.n459 B.n267 71.676
R1326 B.n457 B.n456 71.676
R1327 B.n452 B.n451 71.676
R1328 B.n449 B.n448 71.676
R1329 B.n444 B.n443 71.676
R1330 B.n441 B.n440 71.676
R1331 B.n436 B.n435 71.676
R1332 B.n433 B.n432 71.676
R1333 B.n428 B.n427 71.676
R1334 B.n425 B.n424 71.676
R1335 B.n420 B.n419 71.676
R1336 B.n417 B.n416 71.676
R1337 B.n412 B.n411 71.676
R1338 B.n409 B.n408 71.676
R1339 B.n404 B.n403 71.676
R1340 B.n401 B.n400 71.676
R1341 B.n395 B.n394 71.676
R1342 B.n392 B.n391 71.676
R1343 B.n387 B.n386 71.676
R1344 B.n384 B.n383 71.676
R1345 B.n379 B.n378 71.676
R1346 B.n374 B.n293 71.676
R1347 B.n372 B.n371 71.676
R1348 B.n367 B.n366 71.676
R1349 B.n364 B.n363 71.676
R1350 B.n359 B.n358 71.676
R1351 B.n356 B.n355 71.676
R1352 B.n351 B.n350 71.676
R1353 B.n348 B.n347 71.676
R1354 B.n343 B.n342 71.676
R1355 B.n340 B.n339 71.676
R1356 B.n335 B.n334 71.676
R1357 B.n332 B.n331 71.676
R1358 B.n327 B.n326 71.676
R1359 B.n324 B.n323 71.676
R1360 B.n319 B.n318 71.676
R1361 B.n316 B.n315 71.676
R1362 B.n311 B.n310 71.676
R1363 B.n291 B.n290 66.1338
R1364 B.n285 B.n284 66.1338
R1365 B.n127 B.n126 66.1338
R1366 B.n134 B.n133 66.1338
R1367 B.n292 B.n291 59.5399
R1368 B.n398 B.n285 59.5399
R1369 B.n128 B.n127 59.5399
R1370 B.n789 B.n134 59.5399
R1371 B.n470 B.n260 49.4224
R1372 B.n476 B.n260 49.4224
R1373 B.n476 B.n256 49.4224
R1374 B.n482 B.n256 49.4224
R1375 B.n482 B.n252 49.4224
R1376 B.n488 B.n252 49.4224
R1377 B.n488 B.n248 49.4224
R1378 B.n494 B.n248 49.4224
R1379 B.n500 B.n244 49.4224
R1380 B.n500 B.n240 49.4224
R1381 B.n506 B.n240 49.4224
R1382 B.n506 B.n236 49.4224
R1383 B.n512 B.n236 49.4224
R1384 B.n512 B.n232 49.4224
R1385 B.n518 B.n232 49.4224
R1386 B.n518 B.n228 49.4224
R1387 B.n524 B.n228 49.4224
R1388 B.n524 B.n223 49.4224
R1389 B.n530 B.n223 49.4224
R1390 B.n530 B.n224 49.4224
R1391 B.n536 B.n216 49.4224
R1392 B.n542 B.n216 49.4224
R1393 B.n542 B.n212 49.4224
R1394 B.n548 B.n212 49.4224
R1395 B.n548 B.n208 49.4224
R1396 B.n554 B.n208 49.4224
R1397 B.n554 B.n204 49.4224
R1398 B.n561 B.n204 49.4224
R1399 B.n561 B.n560 49.4224
R1400 B.n567 B.n197 49.4224
R1401 B.n573 B.n197 49.4224
R1402 B.n573 B.n193 49.4224
R1403 B.n579 B.n193 49.4224
R1404 B.n579 B.n189 49.4224
R1405 B.n585 B.n189 49.4224
R1406 B.n585 B.n184 49.4224
R1407 B.n591 B.n184 49.4224
R1408 B.n591 B.n185 49.4224
R1409 B.n597 B.n177 49.4224
R1410 B.n603 B.n177 49.4224
R1411 B.n603 B.n173 49.4224
R1412 B.n609 B.n173 49.4224
R1413 B.n609 B.n169 49.4224
R1414 B.n615 B.n169 49.4224
R1415 B.n615 B.n165 49.4224
R1416 B.n622 B.n165 49.4224
R1417 B.n622 B.n621 49.4224
R1418 B.n628 B.n158 49.4224
R1419 B.n635 B.n158 49.4224
R1420 B.n635 B.n154 49.4224
R1421 B.n641 B.n154 49.4224
R1422 B.n641 B.n4 49.4224
R1423 B.n995 B.n4 49.4224
R1424 B.n995 B.n994 49.4224
R1425 B.n994 B.n993 49.4224
R1426 B.n993 B.n8 49.4224
R1427 B.n987 B.n8 49.4224
R1428 B.n987 B.n986 49.4224
R1429 B.n986 B.n985 49.4224
R1430 B.n979 B.n18 49.4224
R1431 B.n979 B.n978 49.4224
R1432 B.n978 B.n977 49.4224
R1433 B.n977 B.n22 49.4224
R1434 B.n971 B.n22 49.4224
R1435 B.n971 B.n970 49.4224
R1436 B.n970 B.n969 49.4224
R1437 B.n969 B.n29 49.4224
R1438 B.n963 B.n29 49.4224
R1439 B.n962 B.n961 49.4224
R1440 B.n961 B.n36 49.4224
R1441 B.n955 B.n36 49.4224
R1442 B.n955 B.n954 49.4224
R1443 B.n954 B.n953 49.4224
R1444 B.n953 B.n43 49.4224
R1445 B.n947 B.n43 49.4224
R1446 B.n947 B.n946 49.4224
R1447 B.n946 B.n945 49.4224
R1448 B.n939 B.n53 49.4224
R1449 B.n939 B.n938 49.4224
R1450 B.n938 B.n937 49.4224
R1451 B.n937 B.n57 49.4224
R1452 B.n931 B.n57 49.4224
R1453 B.n931 B.n930 49.4224
R1454 B.n930 B.n929 49.4224
R1455 B.n929 B.n64 49.4224
R1456 B.n923 B.n64 49.4224
R1457 B.n922 B.n921 49.4224
R1458 B.n921 B.n71 49.4224
R1459 B.n915 B.n71 49.4224
R1460 B.n915 B.n914 49.4224
R1461 B.n914 B.n913 49.4224
R1462 B.n913 B.n78 49.4224
R1463 B.n907 B.n78 49.4224
R1464 B.n907 B.n906 49.4224
R1465 B.n906 B.n905 49.4224
R1466 B.n905 B.n85 49.4224
R1467 B.n899 B.n85 49.4224
R1468 B.n899 B.n898 49.4224
R1469 B.n897 B.n92 49.4224
R1470 B.n891 B.n92 49.4224
R1471 B.n891 B.n890 49.4224
R1472 B.n890 B.n889 49.4224
R1473 B.n889 B.n99 49.4224
R1474 B.n883 B.n99 49.4224
R1475 B.n883 B.n882 49.4224
R1476 B.n882 B.n881 49.4224
R1477 B.t9 B.n244 46.5152
R1478 B.n898 B.t13 46.5152
R1479 B.n718 B.n717 36.3712
R1480 B.n879 B.n878 36.3712
R1481 B.n472 B.n262 36.3712
R1482 B.n468 B.n467 36.3712
R1483 B.n536 B.t3 34.8865
R1484 B.n923 B.t0 34.8865
R1485 B.n567 B.t1 33.4329
R1486 B.n945 B.t7 33.4329
R1487 B.n597 B.t6 31.9794
R1488 B.n963 B.t2 31.9794
R1489 B.n628 B.t4 30.5258
R1490 B.n985 B.t5 30.5258
R1491 B.n621 B.t4 18.8971
R1492 B.n18 B.t5 18.8971
R1493 B B.n997 18.0485
R1494 B.n185 B.t6 17.4435
R1495 B.t2 B.n962 17.4435
R1496 B.n560 B.t1 15.9899
R1497 B.n53 B.t7 15.9899
R1498 B.n224 B.t3 14.5363
R1499 B.t0 B.n922 14.5363
R1500 B.n878 B.n877 10.6151
R1501 B.n877 B.n108 10.6151
R1502 B.n871 B.n108 10.6151
R1503 B.n871 B.n870 10.6151
R1504 B.n870 B.n869 10.6151
R1505 B.n869 B.n110 10.6151
R1506 B.n863 B.n110 10.6151
R1507 B.n863 B.n862 10.6151
R1508 B.n862 B.n861 10.6151
R1509 B.n861 B.n112 10.6151
R1510 B.n855 B.n112 10.6151
R1511 B.n855 B.n854 10.6151
R1512 B.n854 B.n853 10.6151
R1513 B.n853 B.n114 10.6151
R1514 B.n847 B.n114 10.6151
R1515 B.n847 B.n846 10.6151
R1516 B.n846 B.n845 10.6151
R1517 B.n845 B.n116 10.6151
R1518 B.n839 B.n116 10.6151
R1519 B.n839 B.n838 10.6151
R1520 B.n838 B.n837 10.6151
R1521 B.n837 B.n118 10.6151
R1522 B.n831 B.n118 10.6151
R1523 B.n831 B.n830 10.6151
R1524 B.n830 B.n829 10.6151
R1525 B.n829 B.n120 10.6151
R1526 B.n823 B.n120 10.6151
R1527 B.n823 B.n822 10.6151
R1528 B.n822 B.n821 10.6151
R1529 B.n821 B.n122 10.6151
R1530 B.n815 B.n122 10.6151
R1531 B.n815 B.n814 10.6151
R1532 B.n814 B.n813 10.6151
R1533 B.n813 B.n124 10.6151
R1534 B.n807 B.n806 10.6151
R1535 B.n806 B.n805 10.6151
R1536 B.n805 B.n129 10.6151
R1537 B.n799 B.n129 10.6151
R1538 B.n799 B.n798 10.6151
R1539 B.n798 B.n797 10.6151
R1540 B.n797 B.n131 10.6151
R1541 B.n791 B.n131 10.6151
R1542 B.n791 B.n790 10.6151
R1543 B.n788 B.n135 10.6151
R1544 B.n782 B.n135 10.6151
R1545 B.n782 B.n781 10.6151
R1546 B.n781 B.n780 10.6151
R1547 B.n780 B.n137 10.6151
R1548 B.n774 B.n137 10.6151
R1549 B.n774 B.n773 10.6151
R1550 B.n773 B.n772 10.6151
R1551 B.n772 B.n139 10.6151
R1552 B.n766 B.n139 10.6151
R1553 B.n766 B.n765 10.6151
R1554 B.n765 B.n764 10.6151
R1555 B.n764 B.n141 10.6151
R1556 B.n758 B.n141 10.6151
R1557 B.n758 B.n757 10.6151
R1558 B.n757 B.n756 10.6151
R1559 B.n756 B.n143 10.6151
R1560 B.n750 B.n143 10.6151
R1561 B.n750 B.n749 10.6151
R1562 B.n749 B.n748 10.6151
R1563 B.n748 B.n145 10.6151
R1564 B.n742 B.n145 10.6151
R1565 B.n742 B.n741 10.6151
R1566 B.n741 B.n740 10.6151
R1567 B.n740 B.n147 10.6151
R1568 B.n734 B.n147 10.6151
R1569 B.n734 B.n733 10.6151
R1570 B.n733 B.n732 10.6151
R1571 B.n732 B.n149 10.6151
R1572 B.n726 B.n149 10.6151
R1573 B.n726 B.n725 10.6151
R1574 B.n725 B.n724 10.6151
R1575 B.n724 B.n151 10.6151
R1576 B.n718 B.n151 10.6151
R1577 B.n473 B.n472 10.6151
R1578 B.n474 B.n473 10.6151
R1579 B.n474 B.n254 10.6151
R1580 B.n484 B.n254 10.6151
R1581 B.n485 B.n484 10.6151
R1582 B.n486 B.n485 10.6151
R1583 B.n486 B.n246 10.6151
R1584 B.n496 B.n246 10.6151
R1585 B.n497 B.n496 10.6151
R1586 B.n498 B.n497 10.6151
R1587 B.n498 B.n238 10.6151
R1588 B.n508 B.n238 10.6151
R1589 B.n509 B.n508 10.6151
R1590 B.n510 B.n509 10.6151
R1591 B.n510 B.n230 10.6151
R1592 B.n520 B.n230 10.6151
R1593 B.n521 B.n520 10.6151
R1594 B.n522 B.n521 10.6151
R1595 B.n522 B.n221 10.6151
R1596 B.n532 B.n221 10.6151
R1597 B.n533 B.n532 10.6151
R1598 B.n534 B.n533 10.6151
R1599 B.n534 B.n214 10.6151
R1600 B.n544 B.n214 10.6151
R1601 B.n545 B.n544 10.6151
R1602 B.n546 B.n545 10.6151
R1603 B.n546 B.n206 10.6151
R1604 B.n556 B.n206 10.6151
R1605 B.n557 B.n556 10.6151
R1606 B.n558 B.n557 10.6151
R1607 B.n558 B.n199 10.6151
R1608 B.n569 B.n199 10.6151
R1609 B.n570 B.n569 10.6151
R1610 B.n571 B.n570 10.6151
R1611 B.n571 B.n191 10.6151
R1612 B.n581 B.n191 10.6151
R1613 B.n582 B.n581 10.6151
R1614 B.n583 B.n582 10.6151
R1615 B.n583 B.n182 10.6151
R1616 B.n593 B.n182 10.6151
R1617 B.n594 B.n593 10.6151
R1618 B.n595 B.n594 10.6151
R1619 B.n595 B.n175 10.6151
R1620 B.n605 B.n175 10.6151
R1621 B.n606 B.n605 10.6151
R1622 B.n607 B.n606 10.6151
R1623 B.n607 B.n167 10.6151
R1624 B.n617 B.n167 10.6151
R1625 B.n618 B.n617 10.6151
R1626 B.n619 B.n618 10.6151
R1627 B.n619 B.n160 10.6151
R1628 B.n630 B.n160 10.6151
R1629 B.n631 B.n630 10.6151
R1630 B.n633 B.n631 10.6151
R1631 B.n633 B.n632 10.6151
R1632 B.n632 B.n152 10.6151
R1633 B.n644 B.n152 10.6151
R1634 B.n645 B.n644 10.6151
R1635 B.n646 B.n645 10.6151
R1636 B.n647 B.n646 10.6151
R1637 B.n649 B.n647 10.6151
R1638 B.n650 B.n649 10.6151
R1639 B.n651 B.n650 10.6151
R1640 B.n652 B.n651 10.6151
R1641 B.n654 B.n652 10.6151
R1642 B.n655 B.n654 10.6151
R1643 B.n656 B.n655 10.6151
R1644 B.n657 B.n656 10.6151
R1645 B.n659 B.n657 10.6151
R1646 B.n660 B.n659 10.6151
R1647 B.n661 B.n660 10.6151
R1648 B.n662 B.n661 10.6151
R1649 B.n664 B.n662 10.6151
R1650 B.n665 B.n664 10.6151
R1651 B.n666 B.n665 10.6151
R1652 B.n667 B.n666 10.6151
R1653 B.n669 B.n667 10.6151
R1654 B.n670 B.n669 10.6151
R1655 B.n671 B.n670 10.6151
R1656 B.n672 B.n671 10.6151
R1657 B.n674 B.n672 10.6151
R1658 B.n675 B.n674 10.6151
R1659 B.n676 B.n675 10.6151
R1660 B.n677 B.n676 10.6151
R1661 B.n679 B.n677 10.6151
R1662 B.n680 B.n679 10.6151
R1663 B.n681 B.n680 10.6151
R1664 B.n682 B.n681 10.6151
R1665 B.n684 B.n682 10.6151
R1666 B.n685 B.n684 10.6151
R1667 B.n686 B.n685 10.6151
R1668 B.n687 B.n686 10.6151
R1669 B.n689 B.n687 10.6151
R1670 B.n690 B.n689 10.6151
R1671 B.n691 B.n690 10.6151
R1672 B.n692 B.n691 10.6151
R1673 B.n694 B.n692 10.6151
R1674 B.n695 B.n694 10.6151
R1675 B.n696 B.n695 10.6151
R1676 B.n697 B.n696 10.6151
R1677 B.n699 B.n697 10.6151
R1678 B.n700 B.n699 10.6151
R1679 B.n701 B.n700 10.6151
R1680 B.n702 B.n701 10.6151
R1681 B.n704 B.n702 10.6151
R1682 B.n705 B.n704 10.6151
R1683 B.n706 B.n705 10.6151
R1684 B.n707 B.n706 10.6151
R1685 B.n709 B.n707 10.6151
R1686 B.n710 B.n709 10.6151
R1687 B.n711 B.n710 10.6151
R1688 B.n712 B.n711 10.6151
R1689 B.n714 B.n712 10.6151
R1690 B.n715 B.n714 10.6151
R1691 B.n716 B.n715 10.6151
R1692 B.n717 B.n716 10.6151
R1693 B.n467 B.n466 10.6151
R1694 B.n466 B.n266 10.6151
R1695 B.n461 B.n266 10.6151
R1696 B.n461 B.n460 10.6151
R1697 B.n460 B.n268 10.6151
R1698 B.n455 B.n268 10.6151
R1699 B.n455 B.n454 10.6151
R1700 B.n454 B.n453 10.6151
R1701 B.n453 B.n270 10.6151
R1702 B.n447 B.n270 10.6151
R1703 B.n447 B.n446 10.6151
R1704 B.n446 B.n445 10.6151
R1705 B.n445 B.n272 10.6151
R1706 B.n439 B.n272 10.6151
R1707 B.n439 B.n438 10.6151
R1708 B.n438 B.n437 10.6151
R1709 B.n437 B.n274 10.6151
R1710 B.n431 B.n274 10.6151
R1711 B.n431 B.n430 10.6151
R1712 B.n430 B.n429 10.6151
R1713 B.n429 B.n276 10.6151
R1714 B.n423 B.n276 10.6151
R1715 B.n423 B.n422 10.6151
R1716 B.n422 B.n421 10.6151
R1717 B.n421 B.n278 10.6151
R1718 B.n415 B.n278 10.6151
R1719 B.n415 B.n414 10.6151
R1720 B.n414 B.n413 10.6151
R1721 B.n413 B.n280 10.6151
R1722 B.n407 B.n280 10.6151
R1723 B.n407 B.n406 10.6151
R1724 B.n406 B.n405 10.6151
R1725 B.n405 B.n282 10.6151
R1726 B.n399 B.n282 10.6151
R1727 B.n397 B.n396 10.6151
R1728 B.n396 B.n286 10.6151
R1729 B.n390 B.n286 10.6151
R1730 B.n390 B.n389 10.6151
R1731 B.n389 B.n388 10.6151
R1732 B.n388 B.n288 10.6151
R1733 B.n382 B.n288 10.6151
R1734 B.n382 B.n381 10.6151
R1735 B.n381 B.n380 10.6151
R1736 B.n376 B.n375 10.6151
R1737 B.n375 B.n294 10.6151
R1738 B.n370 B.n294 10.6151
R1739 B.n370 B.n369 10.6151
R1740 B.n369 B.n368 10.6151
R1741 B.n368 B.n296 10.6151
R1742 B.n362 B.n296 10.6151
R1743 B.n362 B.n361 10.6151
R1744 B.n361 B.n360 10.6151
R1745 B.n360 B.n298 10.6151
R1746 B.n354 B.n298 10.6151
R1747 B.n354 B.n353 10.6151
R1748 B.n353 B.n352 10.6151
R1749 B.n352 B.n300 10.6151
R1750 B.n346 B.n300 10.6151
R1751 B.n346 B.n345 10.6151
R1752 B.n345 B.n344 10.6151
R1753 B.n344 B.n302 10.6151
R1754 B.n338 B.n302 10.6151
R1755 B.n338 B.n337 10.6151
R1756 B.n337 B.n336 10.6151
R1757 B.n336 B.n304 10.6151
R1758 B.n330 B.n304 10.6151
R1759 B.n330 B.n329 10.6151
R1760 B.n329 B.n328 10.6151
R1761 B.n328 B.n306 10.6151
R1762 B.n322 B.n306 10.6151
R1763 B.n322 B.n321 10.6151
R1764 B.n321 B.n320 10.6151
R1765 B.n320 B.n308 10.6151
R1766 B.n314 B.n308 10.6151
R1767 B.n314 B.n313 10.6151
R1768 B.n313 B.n312 10.6151
R1769 B.n312 B.n262 10.6151
R1770 B.n468 B.n258 10.6151
R1771 B.n478 B.n258 10.6151
R1772 B.n479 B.n478 10.6151
R1773 B.n480 B.n479 10.6151
R1774 B.n480 B.n250 10.6151
R1775 B.n490 B.n250 10.6151
R1776 B.n491 B.n490 10.6151
R1777 B.n492 B.n491 10.6151
R1778 B.n492 B.n242 10.6151
R1779 B.n502 B.n242 10.6151
R1780 B.n503 B.n502 10.6151
R1781 B.n504 B.n503 10.6151
R1782 B.n504 B.n234 10.6151
R1783 B.n514 B.n234 10.6151
R1784 B.n515 B.n514 10.6151
R1785 B.n516 B.n515 10.6151
R1786 B.n516 B.n226 10.6151
R1787 B.n526 B.n226 10.6151
R1788 B.n527 B.n526 10.6151
R1789 B.n528 B.n527 10.6151
R1790 B.n528 B.n218 10.6151
R1791 B.n538 B.n218 10.6151
R1792 B.n539 B.n538 10.6151
R1793 B.n540 B.n539 10.6151
R1794 B.n540 B.n210 10.6151
R1795 B.n550 B.n210 10.6151
R1796 B.n551 B.n550 10.6151
R1797 B.n552 B.n551 10.6151
R1798 B.n552 B.n202 10.6151
R1799 B.n563 B.n202 10.6151
R1800 B.n564 B.n563 10.6151
R1801 B.n565 B.n564 10.6151
R1802 B.n565 B.n195 10.6151
R1803 B.n575 B.n195 10.6151
R1804 B.n576 B.n575 10.6151
R1805 B.n577 B.n576 10.6151
R1806 B.n577 B.n187 10.6151
R1807 B.n587 B.n187 10.6151
R1808 B.n588 B.n587 10.6151
R1809 B.n589 B.n588 10.6151
R1810 B.n589 B.n179 10.6151
R1811 B.n599 B.n179 10.6151
R1812 B.n600 B.n599 10.6151
R1813 B.n601 B.n600 10.6151
R1814 B.n601 B.n171 10.6151
R1815 B.n611 B.n171 10.6151
R1816 B.n612 B.n611 10.6151
R1817 B.n613 B.n612 10.6151
R1818 B.n613 B.n163 10.6151
R1819 B.n624 B.n163 10.6151
R1820 B.n625 B.n624 10.6151
R1821 B.n626 B.n625 10.6151
R1822 B.n626 B.n156 10.6151
R1823 B.n637 B.n156 10.6151
R1824 B.n638 B.n637 10.6151
R1825 B.n639 B.n638 10.6151
R1826 B.n639 B.n0 10.6151
R1827 B.n991 B.n1 10.6151
R1828 B.n991 B.n990 10.6151
R1829 B.n990 B.n989 10.6151
R1830 B.n989 B.n10 10.6151
R1831 B.n983 B.n10 10.6151
R1832 B.n983 B.n982 10.6151
R1833 B.n982 B.n981 10.6151
R1834 B.n981 B.n16 10.6151
R1835 B.n975 B.n16 10.6151
R1836 B.n975 B.n974 10.6151
R1837 B.n974 B.n973 10.6151
R1838 B.n973 B.n24 10.6151
R1839 B.n967 B.n24 10.6151
R1840 B.n967 B.n966 10.6151
R1841 B.n966 B.n965 10.6151
R1842 B.n965 B.n31 10.6151
R1843 B.n959 B.n31 10.6151
R1844 B.n959 B.n958 10.6151
R1845 B.n958 B.n957 10.6151
R1846 B.n957 B.n38 10.6151
R1847 B.n951 B.n38 10.6151
R1848 B.n951 B.n950 10.6151
R1849 B.n950 B.n949 10.6151
R1850 B.n949 B.n45 10.6151
R1851 B.n943 B.n45 10.6151
R1852 B.n943 B.n942 10.6151
R1853 B.n942 B.n941 10.6151
R1854 B.n941 B.n51 10.6151
R1855 B.n935 B.n51 10.6151
R1856 B.n935 B.n934 10.6151
R1857 B.n934 B.n933 10.6151
R1858 B.n933 B.n59 10.6151
R1859 B.n927 B.n59 10.6151
R1860 B.n927 B.n926 10.6151
R1861 B.n926 B.n925 10.6151
R1862 B.n925 B.n66 10.6151
R1863 B.n919 B.n66 10.6151
R1864 B.n919 B.n918 10.6151
R1865 B.n918 B.n917 10.6151
R1866 B.n917 B.n73 10.6151
R1867 B.n911 B.n73 10.6151
R1868 B.n911 B.n910 10.6151
R1869 B.n910 B.n909 10.6151
R1870 B.n909 B.n80 10.6151
R1871 B.n903 B.n80 10.6151
R1872 B.n903 B.n902 10.6151
R1873 B.n902 B.n901 10.6151
R1874 B.n901 B.n87 10.6151
R1875 B.n895 B.n87 10.6151
R1876 B.n895 B.n894 10.6151
R1877 B.n894 B.n893 10.6151
R1878 B.n893 B.n94 10.6151
R1879 B.n887 B.n94 10.6151
R1880 B.n887 B.n886 10.6151
R1881 B.n886 B.n885 10.6151
R1882 B.n885 B.n101 10.6151
R1883 B.n879 B.n101 10.6151
R1884 B.n128 B.n124 9.36635
R1885 B.n789 B.n788 9.36635
R1886 B.n399 B.n398 9.36635
R1887 B.n376 B.n292 9.36635
R1888 B.n494 B.t9 2.90767
R1889 B.t13 B.n897 2.90767
R1890 B.n997 B.n0 2.81026
R1891 B.n997 B.n1 2.81026
R1892 B.n807 B.n128 1.24928
R1893 B.n790 B.n789 1.24928
R1894 B.n398 B.n397 1.24928
R1895 B.n380 B.n292 1.24928
R1896 VN.n60 VN.n59 161.3
R1897 VN.n58 VN.n32 161.3
R1898 VN.n57 VN.n56 161.3
R1899 VN.n55 VN.n33 161.3
R1900 VN.n54 VN.n53 161.3
R1901 VN.n52 VN.n34 161.3
R1902 VN.n51 VN.n50 161.3
R1903 VN.n49 VN.n48 161.3
R1904 VN.n47 VN.n36 161.3
R1905 VN.n46 VN.n45 161.3
R1906 VN.n44 VN.n37 161.3
R1907 VN.n43 VN.n42 161.3
R1908 VN.n41 VN.n38 161.3
R1909 VN.n29 VN.n28 161.3
R1910 VN.n27 VN.n1 161.3
R1911 VN.n26 VN.n25 161.3
R1912 VN.n24 VN.n2 161.3
R1913 VN.n23 VN.n22 161.3
R1914 VN.n21 VN.n3 161.3
R1915 VN.n20 VN.n19 161.3
R1916 VN.n18 VN.n17 161.3
R1917 VN.n16 VN.n5 161.3
R1918 VN.n15 VN.n14 161.3
R1919 VN.n13 VN.n6 161.3
R1920 VN.n12 VN.n11 161.3
R1921 VN.n10 VN.n7 161.3
R1922 VN.n39 VN.t5 110.55
R1923 VN.n8 VN.t2 110.55
R1924 VN.n9 VN.t6 77.1518
R1925 VN.n4 VN.t4 77.1518
R1926 VN.n0 VN.t7 77.1518
R1927 VN.n40 VN.t1 77.1518
R1928 VN.n35 VN.t0 77.1518
R1929 VN.n31 VN.t3 77.1518
R1930 VN.n30 VN.n0 72.2935
R1931 VN.n61 VN.n31 72.2935
R1932 VN.n15 VN.n6 56.5617
R1933 VN.n46 VN.n37 56.5617
R1934 VN.n26 VN.n2 56.0773
R1935 VN.n57 VN.n33 56.0773
R1936 VN VN.n61 51.7936
R1937 VN.n9 VN.n8 51.645
R1938 VN.n40 VN.n39 51.645
R1939 VN.n22 VN.n2 25.0767
R1940 VN.n53 VN.n33 25.0767
R1941 VN.n11 VN.n10 24.5923
R1942 VN.n11 VN.n6 24.5923
R1943 VN.n16 VN.n15 24.5923
R1944 VN.n17 VN.n16 24.5923
R1945 VN.n21 VN.n20 24.5923
R1946 VN.n22 VN.n21 24.5923
R1947 VN.n27 VN.n26 24.5923
R1948 VN.n28 VN.n27 24.5923
R1949 VN.n42 VN.n37 24.5923
R1950 VN.n42 VN.n41 24.5923
R1951 VN.n53 VN.n52 24.5923
R1952 VN.n52 VN.n51 24.5923
R1953 VN.n48 VN.n47 24.5923
R1954 VN.n47 VN.n46 24.5923
R1955 VN.n59 VN.n58 24.5923
R1956 VN.n58 VN.n57 24.5923
R1957 VN.n10 VN.n9 22.3791
R1958 VN.n17 VN.n4 22.3791
R1959 VN.n41 VN.n40 22.3791
R1960 VN.n48 VN.n35 22.3791
R1961 VN.n28 VN.n0 17.9525
R1962 VN.n59 VN.n31 17.9525
R1963 VN.n39 VN.n38 4.00189
R1964 VN.n8 VN.n7 4.00189
R1965 VN.n20 VN.n4 2.21377
R1966 VN.n51 VN.n35 2.21377
R1967 VN.n61 VN.n60 0.354861
R1968 VN.n30 VN.n29 0.354861
R1969 VN VN.n30 0.267071
R1970 VN.n60 VN.n32 0.189894
R1971 VN.n56 VN.n32 0.189894
R1972 VN.n56 VN.n55 0.189894
R1973 VN.n55 VN.n54 0.189894
R1974 VN.n54 VN.n34 0.189894
R1975 VN.n50 VN.n34 0.189894
R1976 VN.n50 VN.n49 0.189894
R1977 VN.n49 VN.n36 0.189894
R1978 VN.n45 VN.n36 0.189894
R1979 VN.n45 VN.n44 0.189894
R1980 VN.n44 VN.n43 0.189894
R1981 VN.n43 VN.n38 0.189894
R1982 VN.n12 VN.n7 0.189894
R1983 VN.n13 VN.n12 0.189894
R1984 VN.n14 VN.n13 0.189894
R1985 VN.n14 VN.n5 0.189894
R1986 VN.n18 VN.n5 0.189894
R1987 VN.n19 VN.n18 0.189894
R1988 VN.n19 VN.n3 0.189894
R1989 VN.n23 VN.n3 0.189894
R1990 VN.n24 VN.n23 0.189894
R1991 VN.n25 VN.n24 0.189894
R1992 VN.n25 VN.n1 0.189894
R1993 VN.n29 VN.n1 0.189894
R1994 VDD2.n2 VDD2.n1 62.7476
R1995 VDD2.n2 VDD2.n0 62.7476
R1996 VDD2 VDD2.n5 62.7449
R1997 VDD2.n4 VDD2.n3 61.3333
R1998 VDD2.n4 VDD2.n2 45.4437
R1999 VDD2.n5 VDD2.t6 2.00861
R2000 VDD2.n5 VDD2.t2 2.00861
R2001 VDD2.n3 VDD2.t4 2.00861
R2002 VDD2.n3 VDD2.t7 2.00861
R2003 VDD2.n1 VDD2.t3 2.00861
R2004 VDD2.n1 VDD2.t0 2.00861
R2005 VDD2.n0 VDD2.t5 2.00861
R2006 VDD2.n0 VDD2.t1 2.00861
R2007 VDD2 VDD2.n4 1.52852
C0 VDD1 VTAIL 7.56706f
C1 VP VN 7.84913f
C2 VP VTAIL 8.11543f
C3 VN VDD2 7.44421f
C4 VP VDD1 7.86073f
C5 VDD2 VTAIL 7.6247f
C6 VDD1 VDD2 2.02805f
C7 VP VDD2 0.571168f
C8 VN VTAIL 8.101319f
C9 VDD1 VN 0.153016f
C10 VDD2 B 5.743533f
C11 VDD1 B 6.242458f
C12 VTAIL B 9.531887f
C13 VN B 17.183971f
C14 VP B 15.83495f
C15 VDD2.t5 B 0.212178f
C16 VDD2.t1 B 0.212178f
C17 VDD2.n0 B 1.87002f
C18 VDD2.t3 B 0.212178f
C19 VDD2.t0 B 0.212178f
C20 VDD2.n1 B 1.87002f
C21 VDD2.n2 B 3.74271f
C22 VDD2.t4 B 0.212178f
C23 VDD2.t7 B 0.212178f
C24 VDD2.n3 B 1.85592f
C25 VDD2.n4 B 3.225f
C26 VDD2.t6 B 0.212178f
C27 VDD2.t2 B 0.212178f
C28 VDD2.n5 B 1.86998f
C29 VN.t7 B 1.67505f
C30 VN.n0 B 0.675434f
C31 VN.n1 B 0.02037f
C32 VN.n2 B 0.024236f
C33 VN.n3 B 0.02037f
C34 VN.t4 B 1.67505f
C35 VN.n4 B 0.596536f
C36 VN.n5 B 0.02037f
C37 VN.n6 B 0.029611f
C38 VN.n7 B 0.232655f
C39 VN.t6 B 1.67505f
C40 VN.t2 B 1.89806f
C41 VN.n8 B 0.63268f
C42 VN.n9 B 0.67006f
C43 VN.n10 B 0.036096f
C44 VN.n11 B 0.037775f
C45 VN.n12 B 0.02037f
C46 VN.n13 B 0.02037f
C47 VN.n14 B 0.02037f
C48 VN.n15 B 0.029611f
C49 VN.n16 B 0.037775f
C50 VN.n17 B 0.036096f
C51 VN.n18 B 0.02037f
C52 VN.n19 B 0.02037f
C53 VN.n20 B 0.020805f
C54 VN.n21 B 0.037775f
C55 VN.n22 B 0.038128f
C56 VN.n23 B 0.02037f
C57 VN.n24 B 0.02037f
C58 VN.n25 B 0.02037f
C59 VN.n26 B 0.034634f
C60 VN.n27 B 0.037775f
C61 VN.n28 B 0.03274f
C62 VN.n29 B 0.032872f
C63 VN.n30 B 0.044836f
C64 VN.t3 B 1.67505f
C65 VN.n31 B 0.675434f
C66 VN.n32 B 0.02037f
C67 VN.n33 B 0.024236f
C68 VN.n34 B 0.02037f
C69 VN.t0 B 1.67505f
C70 VN.n35 B 0.596536f
C71 VN.n36 B 0.02037f
C72 VN.n37 B 0.029611f
C73 VN.n38 B 0.232655f
C74 VN.t1 B 1.67505f
C75 VN.t5 B 1.89806f
C76 VN.n39 B 0.63268f
C77 VN.n40 B 0.67006f
C78 VN.n41 B 0.036096f
C79 VN.n42 B 0.037775f
C80 VN.n43 B 0.02037f
C81 VN.n44 B 0.02037f
C82 VN.n45 B 0.02037f
C83 VN.n46 B 0.029611f
C84 VN.n47 B 0.037775f
C85 VN.n48 B 0.036096f
C86 VN.n49 B 0.02037f
C87 VN.n50 B 0.02037f
C88 VN.n51 B 0.020805f
C89 VN.n52 B 0.037775f
C90 VN.n53 B 0.038128f
C91 VN.n54 B 0.02037f
C92 VN.n55 B 0.02037f
C93 VN.n56 B 0.02037f
C94 VN.n57 B 0.034634f
C95 VN.n58 B 0.037775f
C96 VN.n59 B 0.03274f
C97 VN.n60 B 0.032872f
C98 VN.n61 B 1.21623f
C99 VDD1.t4 B 0.217134f
C100 VDD1.t6 B 0.217134f
C101 VDD1.n0 B 1.91507f
C102 VDD1.t1 B 0.217134f
C103 VDD1.t7 B 0.217134f
C104 VDD1.n1 B 1.91369f
C105 VDD1.t0 B 0.217134f
C106 VDD1.t3 B 0.217134f
C107 VDD1.n2 B 1.91369f
C108 VDD1.n3 B 3.88796f
C109 VDD1.t2 B 0.217134f
C110 VDD1.t5 B 0.217134f
C111 VDD1.n4 B 1.89927f
C112 VDD1.n5 B 3.33497f
C113 VTAIL.t2 B 0.163584f
C114 VTAIL.t7 B 0.163584f
C115 VTAIL.n0 B 1.36546f
C116 VTAIL.n1 B 0.418751f
C117 VTAIL.t5 B 1.74068f
C118 VTAIL.n2 B 0.517522f
C119 VTAIL.t13 B 1.74068f
C120 VTAIL.n3 B 0.517522f
C121 VTAIL.t9 B 0.163584f
C122 VTAIL.t15 B 0.163584f
C123 VTAIL.n4 B 1.36546f
C124 VTAIL.n5 B 0.613682f
C125 VTAIL.t12 B 1.74068f
C126 VTAIL.n6 B 1.54481f
C127 VTAIL.t3 B 1.74068f
C128 VTAIL.n7 B 1.54481f
C129 VTAIL.t1 B 0.163584f
C130 VTAIL.t6 B 0.163584f
C131 VTAIL.n8 B 1.36547f
C132 VTAIL.n9 B 0.613674f
C133 VTAIL.t4 B 1.74068f
C134 VTAIL.n10 B 0.517515f
C135 VTAIL.t11 B 1.74068f
C136 VTAIL.n11 B 0.517515f
C137 VTAIL.t8 B 0.163584f
C138 VTAIL.t14 B 0.163584f
C139 VTAIL.n12 B 1.36547f
C140 VTAIL.n13 B 0.613674f
C141 VTAIL.t10 B 1.74069f
C142 VTAIL.n14 B 1.54481f
C143 VTAIL.t0 B 1.74068f
C144 VTAIL.n15 B 1.54088f
C145 VP.t4 B 1.7131f
C146 VP.n0 B 0.690777f
C147 VP.n1 B 0.020833f
C148 VP.n2 B 0.024787f
C149 VP.n3 B 0.020833f
C150 VP.t7 B 1.7131f
C151 VP.n4 B 0.610087f
C152 VP.n5 B 0.020833f
C153 VP.n6 B 0.030284f
C154 VP.n7 B 0.020833f
C155 VP.t0 B 1.7131f
C156 VP.n8 B 0.038633f
C157 VP.n9 B 0.020833f
C158 VP.n10 B 0.038633f
C159 VP.t2 B 1.7131f
C160 VP.n11 B 0.690777f
C161 VP.n12 B 0.020833f
C162 VP.n13 B 0.024787f
C163 VP.n14 B 0.020833f
C164 VP.t5 B 1.7131f
C165 VP.n15 B 0.610087f
C166 VP.n16 B 0.020833f
C167 VP.n17 B 0.030284f
C168 VP.n18 B 0.237941f
C169 VP.t1 B 1.7131f
C170 VP.t3 B 1.94117f
C171 VP.n19 B 0.647053f
C172 VP.n20 B 0.685281f
C173 VP.n21 B 0.036916f
C174 VP.n22 B 0.038633f
C175 VP.n23 B 0.020833f
C176 VP.n24 B 0.020833f
C177 VP.n25 B 0.020833f
C178 VP.n26 B 0.030284f
C179 VP.n27 B 0.038633f
C180 VP.n28 B 0.036916f
C181 VP.n29 B 0.020833f
C182 VP.n30 B 0.020833f
C183 VP.n31 B 0.021277f
C184 VP.n32 B 0.038633f
C185 VP.n33 B 0.038994f
C186 VP.n34 B 0.020833f
C187 VP.n35 B 0.020833f
C188 VP.n36 B 0.020833f
C189 VP.n37 B 0.03542f
C190 VP.n38 B 0.038633f
C191 VP.n39 B 0.033483f
C192 VP.n40 B 0.033619f
C193 VP.n41 B 1.23543f
C194 VP.n42 B 1.24998f
C195 VP.t6 B 1.7131f
C196 VP.n43 B 0.690777f
C197 VP.n44 B 0.033483f
C198 VP.n45 B 0.033619f
C199 VP.n46 B 0.020833f
C200 VP.n47 B 0.020833f
C201 VP.n48 B 0.03542f
C202 VP.n49 B 0.024787f
C203 VP.n50 B 0.038994f
C204 VP.n51 B 0.020833f
C205 VP.n52 B 0.020833f
C206 VP.n53 B 0.020833f
C207 VP.n54 B 0.021277f
C208 VP.n55 B 0.610087f
C209 VP.n56 B 0.036916f
C210 VP.n57 B 0.038633f
C211 VP.n58 B 0.020833f
C212 VP.n59 B 0.020833f
C213 VP.n60 B 0.020833f
C214 VP.n61 B 0.030284f
C215 VP.n62 B 0.038633f
C216 VP.n63 B 0.036916f
C217 VP.n64 B 0.020833f
C218 VP.n65 B 0.020833f
C219 VP.n66 B 0.021277f
C220 VP.n67 B 0.038633f
C221 VP.n68 B 0.038994f
C222 VP.n69 B 0.020833f
C223 VP.n70 B 0.020833f
C224 VP.n71 B 0.020833f
C225 VP.n72 B 0.03542f
C226 VP.n73 B 0.038633f
C227 VP.n74 B 0.033483f
C228 VP.n75 B 0.033619f
C229 VP.n76 B 0.045855f
.ends

