* NGSPICE file created from diff_pair_sample_0721.ext - technology: sky130A

.subckt diff_pair_sample_0721 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VP.t0 VDD1.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X1 VDD2.t9 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0.5115 ps=3.43 w=3.1 l=0.76
X2 VTAIL.t19 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X3 VTAIL.t17 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X4 VTAIL.t15 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0 ps=0 w=3.1 l=0.76
X6 VDD2.t6 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=1.209 ps=6.98 w=3.1 l=0.76
X7 VTAIL.t18 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X8 VDD1.t8 VP.t2 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0.5115 ps=3.43 w=3.1 l=0.76
X9 VTAIL.t6 VN.t5 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X10 VDD2.t3 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X11 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0 ps=0 w=3.1 l=0.76
X12 VTAIL.t13 VP.t3 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X13 VDD1.t1 VP.t4 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=1.209 ps=6.98 w=3.1 l=0.76
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0 ps=0 w=3.1 l=0.76
X15 VTAIL.t11 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X16 VDD1.t7 VP.t6 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=1.209 ps=6.98 w=3.1 l=0.76
X17 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=1.209 ps=6.98 w=3.1 l=0.76
X18 VDD1.t2 VP.t7 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X19 VDD1.t0 VP.t8 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0.5115 ps=3.43 w=3.1 l=0.76
X20 VDD1.t9 VP.t9 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X21 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5115 pd=3.43 as=0.5115 ps=3.43 w=3.1 l=0.76
X22 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0.5115 ps=3.43 w=3.1 l=0.76
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.209 pd=6.98 as=0 ps=0 w=3.1 l=0.76
R0 VP.n6 VP.t2 170.805
R1 VP.n23 VP.n22 161.3
R2 VP.n10 VP.n3 161.3
R3 VP.n12 VP.n11 161.3
R4 VP.n21 VP.n0 161.3
R5 VP.n15 VP.n2 161.3
R6 VP.n14 VP.n13 161.3
R7 VP.n14 VP.t8 149.992
R8 VP.n16 VP.t5 149.992
R9 VP.n1 VP.t7 149.992
R10 VP.n20 VP.t3 149.992
R11 VP.n22 VP.t4 149.992
R12 VP.n11 VP.t6 149.992
R13 VP.n9 VP.t1 149.992
R14 VP.n8 VP.t9 149.992
R15 VP.n7 VP.t0 149.992
R16 VP.n8 VP.n5 80.6037
R17 VP.n9 VP.n4 80.6037
R18 VP.n20 VP.n19 80.6037
R19 VP.n18 VP.n1 80.6037
R20 VP.n17 VP.n16 80.6037
R21 VP.n16 VP.n1 48.2005
R22 VP.n20 VP.n1 48.2005
R23 VP.n9 VP.n8 48.2005
R24 VP.n8 VP.n7 48.2005
R25 VP.n16 VP.n15 40.8975
R26 VP.n21 VP.n20 40.8975
R27 VP.n10 VP.n9 40.8975
R28 VP.n13 VP.n12 36.2846
R29 VP.n6 VP.n5 31.6317
R30 VP.n7 VP.n6 17.5473
R31 VP.n15 VP.n14 7.30353
R32 VP.n22 VP.n21 7.30353
R33 VP.n11 VP.n10 7.30353
R34 VP.n5 VP.n4 0.380177
R35 VP.n18 VP.n17 0.380177
R36 VP.n19 VP.n18 0.380177
R37 VP.n4 VP.n3 0.285035
R38 VP.n17 VP.n2 0.285035
R39 VP.n19 VP.n0 0.285035
R40 VP.n12 VP.n3 0.189894
R41 VP.n13 VP.n2 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VDD1.n10 VDD1.n0 289.615
R45 VDD1.n27 VDD1.n17 289.615
R46 VDD1.n11 VDD1.n10 185
R47 VDD1.n9 VDD1.n8 185
R48 VDD1.n4 VDD1.n3 185
R49 VDD1.n21 VDD1.n20 185
R50 VDD1.n26 VDD1.n25 185
R51 VDD1.n28 VDD1.n27 185
R52 VDD1.n5 VDD1.t8 148.606
R53 VDD1.n22 VDD1.t0 148.606
R54 VDD1.n10 VDD1.n9 104.615
R55 VDD1.n9 VDD1.n3 104.615
R56 VDD1.n26 VDD1.n20 104.615
R57 VDD1.n27 VDD1.n26 104.615
R58 VDD1.n35 VDD1.n34 78.0106
R59 VDD1.n16 VDD1.n15 77.3613
R60 VDD1.n37 VDD1.n36 77.3612
R61 VDD1.n33 VDD1.n32 77.3612
R62 VDD1.t8 VDD1.n3 52.3082
R63 VDD1.t0 VDD1.n20 52.3082
R64 VDD1.n16 VDD1.n14 49.4159
R65 VDD1.n33 VDD1.n31 49.4159
R66 VDD1.n37 VDD1.n35 31.9039
R67 VDD1.n5 VDD1.n4 15.5966
R68 VDD1.n22 VDD1.n21 15.5966
R69 VDD1.n8 VDD1.n7 12.8005
R70 VDD1.n25 VDD1.n24 12.8005
R71 VDD1.n11 VDD1.n2 12.0247
R72 VDD1.n28 VDD1.n19 12.0247
R73 VDD1.n12 VDD1.n0 11.249
R74 VDD1.n29 VDD1.n17 11.249
R75 VDD1.n14 VDD1.n13 9.45567
R76 VDD1.n31 VDD1.n30 9.45567
R77 VDD1.n13 VDD1.n12 9.3005
R78 VDD1.n2 VDD1.n1 9.3005
R79 VDD1.n7 VDD1.n6 9.3005
R80 VDD1.n30 VDD1.n29 9.3005
R81 VDD1.n19 VDD1.n18 9.3005
R82 VDD1.n24 VDD1.n23 9.3005
R83 VDD1.n36 VDD1.t6 6.3876
R84 VDD1.n36 VDD1.t7 6.3876
R85 VDD1.n15 VDD1.t3 6.3876
R86 VDD1.n15 VDD1.t9 6.3876
R87 VDD1.n34 VDD1.t5 6.3876
R88 VDD1.n34 VDD1.t1 6.3876
R89 VDD1.n32 VDD1.t4 6.3876
R90 VDD1.n32 VDD1.t2 6.3876
R91 VDD1.n6 VDD1.n5 4.46457
R92 VDD1.n23 VDD1.n22 4.46457
R93 VDD1.n14 VDD1.n0 2.71565
R94 VDD1.n31 VDD1.n17 2.71565
R95 VDD1.n12 VDD1.n11 1.93989
R96 VDD1.n29 VDD1.n28 1.93989
R97 VDD1.n8 VDD1.n2 1.16414
R98 VDD1.n25 VDD1.n19 1.16414
R99 VDD1 VDD1.n37 0.647052
R100 VDD1.n7 VDD1.n4 0.388379
R101 VDD1.n24 VDD1.n21 0.388379
R102 VDD1 VDD1.n16 0.293603
R103 VDD1.n35 VDD1.n33 0.180068
R104 VDD1.n13 VDD1.n1 0.155672
R105 VDD1.n6 VDD1.n1 0.155672
R106 VDD1.n23 VDD1.n18 0.155672
R107 VDD1.n30 VDD1.n18 0.155672
R108 VTAIL.n72 VTAIL.n62 289.615
R109 VTAIL.n12 VTAIL.n2 289.615
R110 VTAIL.n56 VTAIL.n46 289.615
R111 VTAIL.n36 VTAIL.n26 289.615
R112 VTAIL.n66 VTAIL.n65 185
R113 VTAIL.n71 VTAIL.n70 185
R114 VTAIL.n73 VTAIL.n72 185
R115 VTAIL.n6 VTAIL.n5 185
R116 VTAIL.n11 VTAIL.n10 185
R117 VTAIL.n13 VTAIL.n12 185
R118 VTAIL.n57 VTAIL.n56 185
R119 VTAIL.n55 VTAIL.n54 185
R120 VTAIL.n50 VTAIL.n49 185
R121 VTAIL.n37 VTAIL.n36 185
R122 VTAIL.n35 VTAIL.n34 185
R123 VTAIL.n30 VTAIL.n29 185
R124 VTAIL.n67 VTAIL.t5 148.606
R125 VTAIL.n7 VTAIL.t12 148.606
R126 VTAIL.n51 VTAIL.t10 148.606
R127 VTAIL.n31 VTAIL.t2 148.606
R128 VTAIL.n71 VTAIL.n65 104.615
R129 VTAIL.n72 VTAIL.n71 104.615
R130 VTAIL.n11 VTAIL.n5 104.615
R131 VTAIL.n12 VTAIL.n11 104.615
R132 VTAIL.n56 VTAIL.n55 104.615
R133 VTAIL.n55 VTAIL.n49 104.615
R134 VTAIL.n36 VTAIL.n35 104.615
R135 VTAIL.n35 VTAIL.n29 104.615
R136 VTAIL.n45 VTAIL.n44 60.6825
R137 VTAIL.n43 VTAIL.n42 60.6825
R138 VTAIL.n25 VTAIL.n24 60.6825
R139 VTAIL.n23 VTAIL.n22 60.6825
R140 VTAIL.n79 VTAIL.n78 60.6824
R141 VTAIL.n1 VTAIL.n0 60.6824
R142 VTAIL.n19 VTAIL.n18 60.6824
R143 VTAIL.n21 VTAIL.n20 60.6824
R144 VTAIL.t5 VTAIL.n65 52.3082
R145 VTAIL.t12 VTAIL.n5 52.3082
R146 VTAIL.t10 VTAIL.n49 52.3082
R147 VTAIL.t2 VTAIL.n29 52.3082
R148 VTAIL.n77 VTAIL.n76 31.7975
R149 VTAIL.n17 VTAIL.n16 31.7975
R150 VTAIL.n61 VTAIL.n60 31.7975
R151 VTAIL.n41 VTAIL.n40 31.7975
R152 VTAIL.n23 VTAIL.n21 16.9186
R153 VTAIL.n77 VTAIL.n61 15.9789
R154 VTAIL.n67 VTAIL.n66 15.5966
R155 VTAIL.n7 VTAIL.n6 15.5966
R156 VTAIL.n51 VTAIL.n50 15.5966
R157 VTAIL.n31 VTAIL.n30 15.5966
R158 VTAIL.n70 VTAIL.n69 12.8005
R159 VTAIL.n10 VTAIL.n9 12.8005
R160 VTAIL.n54 VTAIL.n53 12.8005
R161 VTAIL.n34 VTAIL.n33 12.8005
R162 VTAIL.n73 VTAIL.n64 12.0247
R163 VTAIL.n13 VTAIL.n4 12.0247
R164 VTAIL.n57 VTAIL.n48 12.0247
R165 VTAIL.n37 VTAIL.n28 12.0247
R166 VTAIL.n74 VTAIL.n62 11.249
R167 VTAIL.n14 VTAIL.n2 11.249
R168 VTAIL.n58 VTAIL.n46 11.249
R169 VTAIL.n38 VTAIL.n26 11.249
R170 VTAIL.n76 VTAIL.n75 9.45567
R171 VTAIL.n16 VTAIL.n15 9.45567
R172 VTAIL.n60 VTAIL.n59 9.45567
R173 VTAIL.n40 VTAIL.n39 9.45567
R174 VTAIL.n75 VTAIL.n74 9.3005
R175 VTAIL.n64 VTAIL.n63 9.3005
R176 VTAIL.n69 VTAIL.n68 9.3005
R177 VTAIL.n15 VTAIL.n14 9.3005
R178 VTAIL.n4 VTAIL.n3 9.3005
R179 VTAIL.n9 VTAIL.n8 9.3005
R180 VTAIL.n59 VTAIL.n58 9.3005
R181 VTAIL.n48 VTAIL.n47 9.3005
R182 VTAIL.n53 VTAIL.n52 9.3005
R183 VTAIL.n39 VTAIL.n38 9.3005
R184 VTAIL.n28 VTAIL.n27 9.3005
R185 VTAIL.n33 VTAIL.n32 9.3005
R186 VTAIL.n78 VTAIL.t1 6.3876
R187 VTAIL.n78 VTAIL.t6 6.3876
R188 VTAIL.n0 VTAIL.t0 6.3876
R189 VTAIL.n0 VTAIL.t17 6.3876
R190 VTAIL.n18 VTAIL.t9 6.3876
R191 VTAIL.n18 VTAIL.t13 6.3876
R192 VTAIL.n20 VTAIL.t8 6.3876
R193 VTAIL.n20 VTAIL.t11 6.3876
R194 VTAIL.n44 VTAIL.t7 6.3876
R195 VTAIL.n44 VTAIL.t15 6.3876
R196 VTAIL.n42 VTAIL.t14 6.3876
R197 VTAIL.n42 VTAIL.t16 6.3876
R198 VTAIL.n24 VTAIL.t3 6.3876
R199 VTAIL.n24 VTAIL.t19 6.3876
R200 VTAIL.n22 VTAIL.t4 6.3876
R201 VTAIL.n22 VTAIL.t18 6.3876
R202 VTAIL.n68 VTAIL.n67 4.46457
R203 VTAIL.n8 VTAIL.n7 4.46457
R204 VTAIL.n52 VTAIL.n51 4.46457
R205 VTAIL.n32 VTAIL.n31 4.46457
R206 VTAIL.n76 VTAIL.n62 2.71565
R207 VTAIL.n16 VTAIL.n2 2.71565
R208 VTAIL.n60 VTAIL.n46 2.71565
R209 VTAIL.n40 VTAIL.n26 2.71565
R210 VTAIL.n74 VTAIL.n73 1.93989
R211 VTAIL.n14 VTAIL.n13 1.93989
R212 VTAIL.n58 VTAIL.n57 1.93989
R213 VTAIL.n38 VTAIL.n37 1.93989
R214 VTAIL.n70 VTAIL.n64 1.16414
R215 VTAIL.n10 VTAIL.n4 1.16414
R216 VTAIL.n54 VTAIL.n48 1.16414
R217 VTAIL.n34 VTAIL.n28 1.16414
R218 VTAIL.n25 VTAIL.n23 0.940155
R219 VTAIL.n41 VTAIL.n25 0.940155
R220 VTAIL.n43 VTAIL.n41 0.940155
R221 VTAIL.n45 VTAIL.n43 0.940155
R222 VTAIL.n61 VTAIL.n45 0.940155
R223 VTAIL.n21 VTAIL.n19 0.940155
R224 VTAIL.n19 VTAIL.n17 0.940155
R225 VTAIL.n17 VTAIL.n1 0.940155
R226 VTAIL.n79 VTAIL.n77 0.940155
R227 VTAIL VTAIL.n1 0.763431
R228 VTAIL.n69 VTAIL.n66 0.388379
R229 VTAIL.n9 VTAIL.n6 0.388379
R230 VTAIL.n53 VTAIL.n50 0.388379
R231 VTAIL.n33 VTAIL.n30 0.388379
R232 VTAIL VTAIL.n79 0.177224
R233 VTAIL.n68 VTAIL.n63 0.155672
R234 VTAIL.n75 VTAIL.n63 0.155672
R235 VTAIL.n8 VTAIL.n3 0.155672
R236 VTAIL.n15 VTAIL.n3 0.155672
R237 VTAIL.n59 VTAIL.n47 0.155672
R238 VTAIL.n52 VTAIL.n47 0.155672
R239 VTAIL.n39 VTAIL.n27 0.155672
R240 VTAIL.n32 VTAIL.n27 0.155672
R241 B.n429 B.n428 585
R242 B.n153 B.n73 585
R243 B.n152 B.n151 585
R244 B.n150 B.n149 585
R245 B.n148 B.n147 585
R246 B.n146 B.n145 585
R247 B.n144 B.n143 585
R248 B.n142 B.n141 585
R249 B.n140 B.n139 585
R250 B.n138 B.n137 585
R251 B.n136 B.n135 585
R252 B.n134 B.n133 585
R253 B.n132 B.n131 585
R254 B.n130 B.n129 585
R255 B.n128 B.n127 585
R256 B.n125 B.n124 585
R257 B.n123 B.n122 585
R258 B.n121 B.n120 585
R259 B.n119 B.n118 585
R260 B.n117 B.n116 585
R261 B.n115 B.n114 585
R262 B.n113 B.n112 585
R263 B.n111 B.n110 585
R264 B.n109 B.n108 585
R265 B.n107 B.n106 585
R266 B.n104 B.n103 585
R267 B.n102 B.n101 585
R268 B.n100 B.n99 585
R269 B.n98 B.n97 585
R270 B.n96 B.n95 585
R271 B.n94 B.n93 585
R272 B.n92 B.n91 585
R273 B.n90 B.n89 585
R274 B.n88 B.n87 585
R275 B.n86 B.n85 585
R276 B.n84 B.n83 585
R277 B.n82 B.n81 585
R278 B.n80 B.n79 585
R279 B.n54 B.n53 585
R280 B.n434 B.n433 585
R281 B.n427 B.n74 585
R282 B.n74 B.n51 585
R283 B.n426 B.n50 585
R284 B.n438 B.n50 585
R285 B.n425 B.n49 585
R286 B.n439 B.n49 585
R287 B.n424 B.n48 585
R288 B.n440 B.n48 585
R289 B.n423 B.n422 585
R290 B.n422 B.n44 585
R291 B.n421 B.n43 585
R292 B.n446 B.n43 585
R293 B.n420 B.n42 585
R294 B.n447 B.n42 585
R295 B.n419 B.n41 585
R296 B.n448 B.n41 585
R297 B.n418 B.n417 585
R298 B.n417 B.n37 585
R299 B.n416 B.n36 585
R300 B.n454 B.n36 585
R301 B.n415 B.n35 585
R302 B.n455 B.n35 585
R303 B.n414 B.n34 585
R304 B.n456 B.n34 585
R305 B.n413 B.n412 585
R306 B.n412 B.n30 585
R307 B.n411 B.n29 585
R308 B.n462 B.n29 585
R309 B.n410 B.n28 585
R310 B.n463 B.n28 585
R311 B.n409 B.n27 585
R312 B.n464 B.n27 585
R313 B.n408 B.n407 585
R314 B.n407 B.n23 585
R315 B.n406 B.n22 585
R316 B.n470 B.n22 585
R317 B.n405 B.n21 585
R318 B.n471 B.n21 585
R319 B.n404 B.n20 585
R320 B.n472 B.n20 585
R321 B.n403 B.n402 585
R322 B.n402 B.n16 585
R323 B.n401 B.n15 585
R324 B.n478 B.n15 585
R325 B.n400 B.n14 585
R326 B.n479 B.n14 585
R327 B.n399 B.n13 585
R328 B.n480 B.n13 585
R329 B.n398 B.n397 585
R330 B.n397 B.n12 585
R331 B.n396 B.n395 585
R332 B.n396 B.n8 585
R333 B.n394 B.n7 585
R334 B.n487 B.n7 585
R335 B.n393 B.n6 585
R336 B.n488 B.n6 585
R337 B.n392 B.n5 585
R338 B.n489 B.n5 585
R339 B.n391 B.n390 585
R340 B.n390 B.n4 585
R341 B.n389 B.n154 585
R342 B.n389 B.n388 585
R343 B.n378 B.n155 585
R344 B.n381 B.n155 585
R345 B.n380 B.n379 585
R346 B.n382 B.n380 585
R347 B.n377 B.n160 585
R348 B.n160 B.n159 585
R349 B.n376 B.n375 585
R350 B.n375 B.n374 585
R351 B.n162 B.n161 585
R352 B.n163 B.n162 585
R353 B.n367 B.n366 585
R354 B.n368 B.n367 585
R355 B.n365 B.n168 585
R356 B.n168 B.n167 585
R357 B.n364 B.n363 585
R358 B.n363 B.n362 585
R359 B.n170 B.n169 585
R360 B.n171 B.n170 585
R361 B.n355 B.n354 585
R362 B.n356 B.n355 585
R363 B.n353 B.n175 585
R364 B.n179 B.n175 585
R365 B.n352 B.n351 585
R366 B.n351 B.n350 585
R367 B.n177 B.n176 585
R368 B.n178 B.n177 585
R369 B.n343 B.n342 585
R370 B.n344 B.n343 585
R371 B.n341 B.n184 585
R372 B.n184 B.n183 585
R373 B.n340 B.n339 585
R374 B.n339 B.n338 585
R375 B.n186 B.n185 585
R376 B.n187 B.n186 585
R377 B.n331 B.n330 585
R378 B.n332 B.n331 585
R379 B.n329 B.n192 585
R380 B.n192 B.n191 585
R381 B.n328 B.n327 585
R382 B.n327 B.n326 585
R383 B.n194 B.n193 585
R384 B.n195 B.n194 585
R385 B.n319 B.n318 585
R386 B.n320 B.n319 585
R387 B.n317 B.n200 585
R388 B.n200 B.n199 585
R389 B.n316 B.n315 585
R390 B.n315 B.n314 585
R391 B.n202 B.n201 585
R392 B.n203 B.n202 585
R393 B.n310 B.n309 585
R394 B.n206 B.n205 585
R395 B.n306 B.n305 585
R396 B.n307 B.n306 585
R397 B.n304 B.n226 585
R398 B.n303 B.n302 585
R399 B.n301 B.n300 585
R400 B.n299 B.n298 585
R401 B.n297 B.n296 585
R402 B.n295 B.n294 585
R403 B.n293 B.n292 585
R404 B.n291 B.n290 585
R405 B.n289 B.n288 585
R406 B.n287 B.n286 585
R407 B.n285 B.n284 585
R408 B.n283 B.n282 585
R409 B.n281 B.n280 585
R410 B.n279 B.n278 585
R411 B.n277 B.n276 585
R412 B.n275 B.n274 585
R413 B.n273 B.n272 585
R414 B.n271 B.n270 585
R415 B.n269 B.n268 585
R416 B.n267 B.n266 585
R417 B.n265 B.n264 585
R418 B.n263 B.n262 585
R419 B.n261 B.n260 585
R420 B.n259 B.n258 585
R421 B.n257 B.n256 585
R422 B.n255 B.n254 585
R423 B.n253 B.n252 585
R424 B.n251 B.n250 585
R425 B.n249 B.n248 585
R426 B.n247 B.n246 585
R427 B.n245 B.n244 585
R428 B.n243 B.n242 585
R429 B.n241 B.n240 585
R430 B.n239 B.n238 585
R431 B.n237 B.n236 585
R432 B.n235 B.n234 585
R433 B.n233 B.n225 585
R434 B.n307 B.n225 585
R435 B.n311 B.n204 585
R436 B.n204 B.n203 585
R437 B.n313 B.n312 585
R438 B.n314 B.n313 585
R439 B.n198 B.n197 585
R440 B.n199 B.n198 585
R441 B.n322 B.n321 585
R442 B.n321 B.n320 585
R443 B.n323 B.n196 585
R444 B.n196 B.n195 585
R445 B.n325 B.n324 585
R446 B.n326 B.n325 585
R447 B.n190 B.n189 585
R448 B.n191 B.n190 585
R449 B.n334 B.n333 585
R450 B.n333 B.n332 585
R451 B.n335 B.n188 585
R452 B.n188 B.n187 585
R453 B.n337 B.n336 585
R454 B.n338 B.n337 585
R455 B.n182 B.n181 585
R456 B.n183 B.n182 585
R457 B.n346 B.n345 585
R458 B.n345 B.n344 585
R459 B.n347 B.n180 585
R460 B.n180 B.n178 585
R461 B.n349 B.n348 585
R462 B.n350 B.n349 585
R463 B.n174 B.n173 585
R464 B.n179 B.n174 585
R465 B.n358 B.n357 585
R466 B.n357 B.n356 585
R467 B.n359 B.n172 585
R468 B.n172 B.n171 585
R469 B.n361 B.n360 585
R470 B.n362 B.n361 585
R471 B.n166 B.n165 585
R472 B.n167 B.n166 585
R473 B.n370 B.n369 585
R474 B.n369 B.n368 585
R475 B.n371 B.n164 585
R476 B.n164 B.n163 585
R477 B.n373 B.n372 585
R478 B.n374 B.n373 585
R479 B.n158 B.n157 585
R480 B.n159 B.n158 585
R481 B.n384 B.n383 585
R482 B.n383 B.n382 585
R483 B.n385 B.n156 585
R484 B.n381 B.n156 585
R485 B.n387 B.n386 585
R486 B.n388 B.n387 585
R487 B.n3 B.n0 585
R488 B.n4 B.n3 585
R489 B.n486 B.n1 585
R490 B.n487 B.n486 585
R491 B.n485 B.n484 585
R492 B.n485 B.n8 585
R493 B.n483 B.n9 585
R494 B.n12 B.n9 585
R495 B.n482 B.n481 585
R496 B.n481 B.n480 585
R497 B.n11 B.n10 585
R498 B.n479 B.n11 585
R499 B.n477 B.n476 585
R500 B.n478 B.n477 585
R501 B.n475 B.n17 585
R502 B.n17 B.n16 585
R503 B.n474 B.n473 585
R504 B.n473 B.n472 585
R505 B.n19 B.n18 585
R506 B.n471 B.n19 585
R507 B.n469 B.n468 585
R508 B.n470 B.n469 585
R509 B.n467 B.n24 585
R510 B.n24 B.n23 585
R511 B.n466 B.n465 585
R512 B.n465 B.n464 585
R513 B.n26 B.n25 585
R514 B.n463 B.n26 585
R515 B.n461 B.n460 585
R516 B.n462 B.n461 585
R517 B.n459 B.n31 585
R518 B.n31 B.n30 585
R519 B.n458 B.n457 585
R520 B.n457 B.n456 585
R521 B.n33 B.n32 585
R522 B.n455 B.n33 585
R523 B.n453 B.n452 585
R524 B.n454 B.n453 585
R525 B.n451 B.n38 585
R526 B.n38 B.n37 585
R527 B.n450 B.n449 585
R528 B.n449 B.n448 585
R529 B.n40 B.n39 585
R530 B.n447 B.n40 585
R531 B.n445 B.n444 585
R532 B.n446 B.n445 585
R533 B.n443 B.n45 585
R534 B.n45 B.n44 585
R535 B.n442 B.n441 585
R536 B.n441 B.n440 585
R537 B.n47 B.n46 585
R538 B.n439 B.n47 585
R539 B.n437 B.n436 585
R540 B.n438 B.n437 585
R541 B.n435 B.n52 585
R542 B.n52 B.n51 585
R543 B.n490 B.n489 585
R544 B.n488 B.n2 585
R545 B.n433 B.n52 511.721
R546 B.n429 B.n74 511.721
R547 B.n225 B.n202 511.721
R548 B.n309 B.n204 511.721
R549 B.n77 B.t10 300.589
R550 B.n75 B.t18 300.589
R551 B.n230 B.t14 300.589
R552 B.n227 B.t21 300.589
R553 B.n431 B.n430 256.663
R554 B.n431 B.n72 256.663
R555 B.n431 B.n71 256.663
R556 B.n431 B.n70 256.663
R557 B.n431 B.n69 256.663
R558 B.n431 B.n68 256.663
R559 B.n431 B.n67 256.663
R560 B.n431 B.n66 256.663
R561 B.n431 B.n65 256.663
R562 B.n431 B.n64 256.663
R563 B.n431 B.n63 256.663
R564 B.n431 B.n62 256.663
R565 B.n431 B.n61 256.663
R566 B.n431 B.n60 256.663
R567 B.n431 B.n59 256.663
R568 B.n431 B.n58 256.663
R569 B.n431 B.n57 256.663
R570 B.n431 B.n56 256.663
R571 B.n431 B.n55 256.663
R572 B.n432 B.n431 256.663
R573 B.n308 B.n307 256.663
R574 B.n307 B.n207 256.663
R575 B.n307 B.n208 256.663
R576 B.n307 B.n209 256.663
R577 B.n307 B.n210 256.663
R578 B.n307 B.n211 256.663
R579 B.n307 B.n212 256.663
R580 B.n307 B.n213 256.663
R581 B.n307 B.n214 256.663
R582 B.n307 B.n215 256.663
R583 B.n307 B.n216 256.663
R584 B.n307 B.n217 256.663
R585 B.n307 B.n218 256.663
R586 B.n307 B.n219 256.663
R587 B.n307 B.n220 256.663
R588 B.n307 B.n221 256.663
R589 B.n307 B.n222 256.663
R590 B.n307 B.n223 256.663
R591 B.n307 B.n224 256.663
R592 B.n492 B.n491 256.663
R593 B.n79 B.n54 163.367
R594 B.n83 B.n82 163.367
R595 B.n87 B.n86 163.367
R596 B.n91 B.n90 163.367
R597 B.n95 B.n94 163.367
R598 B.n99 B.n98 163.367
R599 B.n103 B.n102 163.367
R600 B.n108 B.n107 163.367
R601 B.n112 B.n111 163.367
R602 B.n116 B.n115 163.367
R603 B.n120 B.n119 163.367
R604 B.n124 B.n123 163.367
R605 B.n129 B.n128 163.367
R606 B.n133 B.n132 163.367
R607 B.n137 B.n136 163.367
R608 B.n141 B.n140 163.367
R609 B.n145 B.n144 163.367
R610 B.n149 B.n148 163.367
R611 B.n151 B.n73 163.367
R612 B.n315 B.n202 163.367
R613 B.n315 B.n200 163.367
R614 B.n319 B.n200 163.367
R615 B.n319 B.n194 163.367
R616 B.n327 B.n194 163.367
R617 B.n327 B.n192 163.367
R618 B.n331 B.n192 163.367
R619 B.n331 B.n186 163.367
R620 B.n339 B.n186 163.367
R621 B.n339 B.n184 163.367
R622 B.n343 B.n184 163.367
R623 B.n343 B.n177 163.367
R624 B.n351 B.n177 163.367
R625 B.n351 B.n175 163.367
R626 B.n355 B.n175 163.367
R627 B.n355 B.n170 163.367
R628 B.n363 B.n170 163.367
R629 B.n363 B.n168 163.367
R630 B.n367 B.n168 163.367
R631 B.n367 B.n162 163.367
R632 B.n375 B.n162 163.367
R633 B.n375 B.n160 163.367
R634 B.n380 B.n160 163.367
R635 B.n380 B.n155 163.367
R636 B.n389 B.n155 163.367
R637 B.n390 B.n389 163.367
R638 B.n390 B.n5 163.367
R639 B.n6 B.n5 163.367
R640 B.n7 B.n6 163.367
R641 B.n396 B.n7 163.367
R642 B.n397 B.n396 163.367
R643 B.n397 B.n13 163.367
R644 B.n14 B.n13 163.367
R645 B.n15 B.n14 163.367
R646 B.n402 B.n15 163.367
R647 B.n402 B.n20 163.367
R648 B.n21 B.n20 163.367
R649 B.n22 B.n21 163.367
R650 B.n407 B.n22 163.367
R651 B.n407 B.n27 163.367
R652 B.n28 B.n27 163.367
R653 B.n29 B.n28 163.367
R654 B.n412 B.n29 163.367
R655 B.n412 B.n34 163.367
R656 B.n35 B.n34 163.367
R657 B.n36 B.n35 163.367
R658 B.n417 B.n36 163.367
R659 B.n417 B.n41 163.367
R660 B.n42 B.n41 163.367
R661 B.n43 B.n42 163.367
R662 B.n422 B.n43 163.367
R663 B.n422 B.n48 163.367
R664 B.n49 B.n48 163.367
R665 B.n50 B.n49 163.367
R666 B.n74 B.n50 163.367
R667 B.n306 B.n206 163.367
R668 B.n306 B.n226 163.367
R669 B.n302 B.n301 163.367
R670 B.n298 B.n297 163.367
R671 B.n294 B.n293 163.367
R672 B.n290 B.n289 163.367
R673 B.n286 B.n285 163.367
R674 B.n282 B.n281 163.367
R675 B.n278 B.n277 163.367
R676 B.n274 B.n273 163.367
R677 B.n270 B.n269 163.367
R678 B.n266 B.n265 163.367
R679 B.n262 B.n261 163.367
R680 B.n258 B.n257 163.367
R681 B.n254 B.n253 163.367
R682 B.n250 B.n249 163.367
R683 B.n246 B.n245 163.367
R684 B.n242 B.n241 163.367
R685 B.n238 B.n237 163.367
R686 B.n234 B.n225 163.367
R687 B.n313 B.n204 163.367
R688 B.n313 B.n198 163.367
R689 B.n321 B.n198 163.367
R690 B.n321 B.n196 163.367
R691 B.n325 B.n196 163.367
R692 B.n325 B.n190 163.367
R693 B.n333 B.n190 163.367
R694 B.n333 B.n188 163.367
R695 B.n337 B.n188 163.367
R696 B.n337 B.n182 163.367
R697 B.n345 B.n182 163.367
R698 B.n345 B.n180 163.367
R699 B.n349 B.n180 163.367
R700 B.n349 B.n174 163.367
R701 B.n357 B.n174 163.367
R702 B.n357 B.n172 163.367
R703 B.n361 B.n172 163.367
R704 B.n361 B.n166 163.367
R705 B.n369 B.n166 163.367
R706 B.n369 B.n164 163.367
R707 B.n373 B.n164 163.367
R708 B.n373 B.n158 163.367
R709 B.n383 B.n158 163.367
R710 B.n383 B.n156 163.367
R711 B.n387 B.n156 163.367
R712 B.n387 B.n3 163.367
R713 B.n490 B.n3 163.367
R714 B.n486 B.n2 163.367
R715 B.n486 B.n485 163.367
R716 B.n485 B.n9 163.367
R717 B.n481 B.n9 163.367
R718 B.n481 B.n11 163.367
R719 B.n477 B.n11 163.367
R720 B.n477 B.n17 163.367
R721 B.n473 B.n17 163.367
R722 B.n473 B.n19 163.367
R723 B.n469 B.n19 163.367
R724 B.n469 B.n24 163.367
R725 B.n465 B.n24 163.367
R726 B.n465 B.n26 163.367
R727 B.n461 B.n26 163.367
R728 B.n461 B.n31 163.367
R729 B.n457 B.n31 163.367
R730 B.n457 B.n33 163.367
R731 B.n453 B.n33 163.367
R732 B.n453 B.n38 163.367
R733 B.n449 B.n38 163.367
R734 B.n449 B.n40 163.367
R735 B.n445 B.n40 163.367
R736 B.n445 B.n45 163.367
R737 B.n441 B.n45 163.367
R738 B.n441 B.n47 163.367
R739 B.n437 B.n47 163.367
R740 B.n437 B.n52 163.367
R741 B.n75 B.t19 151.38
R742 B.n230 B.t17 151.38
R743 B.n77 B.t12 151.38
R744 B.n227 B.t23 151.38
R745 B.n307 B.n203 148.418
R746 B.n431 B.n51 148.418
R747 B.n76 B.t20 130.239
R748 B.n231 B.t16 130.239
R749 B.n78 B.t13 130.239
R750 B.n228 B.t22 130.239
R751 B.n314 B.n203 89.3139
R752 B.n314 B.n199 89.3139
R753 B.n320 B.n199 89.3139
R754 B.n320 B.n195 89.3139
R755 B.n326 B.n195 89.3139
R756 B.n332 B.n191 89.3139
R757 B.n332 B.n187 89.3139
R758 B.n338 B.n187 89.3139
R759 B.n338 B.n183 89.3139
R760 B.n344 B.n183 89.3139
R761 B.n350 B.n178 89.3139
R762 B.n350 B.n179 89.3139
R763 B.n356 B.n171 89.3139
R764 B.n362 B.n171 89.3139
R765 B.n368 B.n167 89.3139
R766 B.n368 B.n163 89.3139
R767 B.n374 B.n163 89.3139
R768 B.n382 B.n159 89.3139
R769 B.n382 B.n381 89.3139
R770 B.n388 B.n4 89.3139
R771 B.n489 B.n4 89.3139
R772 B.n489 B.n488 89.3139
R773 B.n488 B.n487 89.3139
R774 B.n487 B.n8 89.3139
R775 B.n480 B.n12 89.3139
R776 B.n480 B.n479 89.3139
R777 B.n478 B.n16 89.3139
R778 B.n472 B.n16 89.3139
R779 B.n472 B.n471 89.3139
R780 B.n470 B.n23 89.3139
R781 B.n464 B.n23 89.3139
R782 B.n463 B.n462 89.3139
R783 B.n462 B.n30 89.3139
R784 B.n456 B.n455 89.3139
R785 B.n455 B.n454 89.3139
R786 B.n454 B.n37 89.3139
R787 B.n448 B.n37 89.3139
R788 B.n448 B.n447 89.3139
R789 B.n446 B.n44 89.3139
R790 B.n440 B.n44 89.3139
R791 B.n440 B.n439 89.3139
R792 B.n439 B.n438 89.3139
R793 B.n438 B.n51 89.3139
R794 B.t15 B.n191 84.0602
R795 B.n447 B.t11 84.0602
R796 B.t8 B.n159 81.4333
R797 B.n479 B.t9 81.4333
R798 B.n362 B.t3 78.8065
R799 B.t1 B.n470 78.8065
R800 B.n433 B.n432 71.676
R801 B.n79 B.n55 71.676
R802 B.n83 B.n56 71.676
R803 B.n87 B.n57 71.676
R804 B.n91 B.n58 71.676
R805 B.n95 B.n59 71.676
R806 B.n99 B.n60 71.676
R807 B.n103 B.n61 71.676
R808 B.n108 B.n62 71.676
R809 B.n112 B.n63 71.676
R810 B.n116 B.n64 71.676
R811 B.n120 B.n65 71.676
R812 B.n124 B.n66 71.676
R813 B.n129 B.n67 71.676
R814 B.n133 B.n68 71.676
R815 B.n137 B.n69 71.676
R816 B.n141 B.n70 71.676
R817 B.n145 B.n71 71.676
R818 B.n149 B.n72 71.676
R819 B.n430 B.n73 71.676
R820 B.n430 B.n429 71.676
R821 B.n151 B.n72 71.676
R822 B.n148 B.n71 71.676
R823 B.n144 B.n70 71.676
R824 B.n140 B.n69 71.676
R825 B.n136 B.n68 71.676
R826 B.n132 B.n67 71.676
R827 B.n128 B.n66 71.676
R828 B.n123 B.n65 71.676
R829 B.n119 B.n64 71.676
R830 B.n115 B.n63 71.676
R831 B.n111 B.n62 71.676
R832 B.n107 B.n61 71.676
R833 B.n102 B.n60 71.676
R834 B.n98 B.n59 71.676
R835 B.n94 B.n58 71.676
R836 B.n90 B.n57 71.676
R837 B.n86 B.n56 71.676
R838 B.n82 B.n55 71.676
R839 B.n432 B.n54 71.676
R840 B.n309 B.n308 71.676
R841 B.n226 B.n207 71.676
R842 B.n301 B.n208 71.676
R843 B.n297 B.n209 71.676
R844 B.n293 B.n210 71.676
R845 B.n289 B.n211 71.676
R846 B.n285 B.n212 71.676
R847 B.n281 B.n213 71.676
R848 B.n277 B.n214 71.676
R849 B.n273 B.n215 71.676
R850 B.n269 B.n216 71.676
R851 B.n265 B.n217 71.676
R852 B.n261 B.n218 71.676
R853 B.n257 B.n219 71.676
R854 B.n253 B.n220 71.676
R855 B.n249 B.n221 71.676
R856 B.n245 B.n222 71.676
R857 B.n241 B.n223 71.676
R858 B.n237 B.n224 71.676
R859 B.n308 B.n206 71.676
R860 B.n302 B.n207 71.676
R861 B.n298 B.n208 71.676
R862 B.n294 B.n209 71.676
R863 B.n290 B.n210 71.676
R864 B.n286 B.n211 71.676
R865 B.n282 B.n212 71.676
R866 B.n278 B.n213 71.676
R867 B.n274 B.n214 71.676
R868 B.n270 B.n215 71.676
R869 B.n266 B.n216 71.676
R870 B.n262 B.n217 71.676
R871 B.n258 B.n218 71.676
R872 B.n254 B.n219 71.676
R873 B.n250 B.n220 71.676
R874 B.n246 B.n221 71.676
R875 B.n242 B.n222 71.676
R876 B.n238 B.n223 71.676
R877 B.n234 B.n224 71.676
R878 B.n491 B.n490 71.676
R879 B.n491 B.n2 71.676
R880 B.n388 B.t2 63.0453
R881 B.t0 B.n8 63.0453
R882 B.n179 B.t7 60.4184
R883 B.t6 B.n463 60.4184
R884 B.n105 B.n78 59.5399
R885 B.n126 B.n76 59.5399
R886 B.n232 B.n231 59.5399
R887 B.n229 B.n228 59.5399
R888 B.t4 B.n178 47.2841
R889 B.t5 B.n30 47.2841
R890 B.n344 B.t4 42.0304
R891 B.n456 B.t5 42.0304
R892 B.n311 B.n310 33.2493
R893 B.n233 B.n201 33.2493
R894 B.n428 B.n427 33.2493
R895 B.n435 B.n434 33.2493
R896 B.n356 B.t7 28.896
R897 B.n464 B.t6 28.896
R898 B.n381 B.t2 26.2692
R899 B.n12 B.t0 26.2692
R900 B.n78 B.n77 21.1399
R901 B.n76 B.n75 21.1399
R902 B.n231 B.n230 21.1399
R903 B.n228 B.n227 21.1399
R904 B B.n492 18.0485
R905 B.n312 B.n311 10.6151
R906 B.n312 B.n197 10.6151
R907 B.n322 B.n197 10.6151
R908 B.n323 B.n322 10.6151
R909 B.n324 B.n323 10.6151
R910 B.n324 B.n189 10.6151
R911 B.n334 B.n189 10.6151
R912 B.n335 B.n334 10.6151
R913 B.n336 B.n335 10.6151
R914 B.n336 B.n181 10.6151
R915 B.n346 B.n181 10.6151
R916 B.n347 B.n346 10.6151
R917 B.n348 B.n347 10.6151
R918 B.n348 B.n173 10.6151
R919 B.n358 B.n173 10.6151
R920 B.n359 B.n358 10.6151
R921 B.n360 B.n359 10.6151
R922 B.n360 B.n165 10.6151
R923 B.n370 B.n165 10.6151
R924 B.n371 B.n370 10.6151
R925 B.n372 B.n371 10.6151
R926 B.n372 B.n157 10.6151
R927 B.n384 B.n157 10.6151
R928 B.n385 B.n384 10.6151
R929 B.n386 B.n385 10.6151
R930 B.n386 B.n0 10.6151
R931 B.n310 B.n205 10.6151
R932 B.n305 B.n205 10.6151
R933 B.n305 B.n304 10.6151
R934 B.n304 B.n303 10.6151
R935 B.n303 B.n300 10.6151
R936 B.n300 B.n299 10.6151
R937 B.n299 B.n296 10.6151
R938 B.n296 B.n295 10.6151
R939 B.n295 B.n292 10.6151
R940 B.n292 B.n291 10.6151
R941 B.n291 B.n288 10.6151
R942 B.n288 B.n287 10.6151
R943 B.n287 B.n284 10.6151
R944 B.n284 B.n283 10.6151
R945 B.n280 B.n279 10.6151
R946 B.n279 B.n276 10.6151
R947 B.n276 B.n275 10.6151
R948 B.n275 B.n272 10.6151
R949 B.n272 B.n271 10.6151
R950 B.n271 B.n268 10.6151
R951 B.n268 B.n267 10.6151
R952 B.n267 B.n264 10.6151
R953 B.n264 B.n263 10.6151
R954 B.n260 B.n259 10.6151
R955 B.n259 B.n256 10.6151
R956 B.n256 B.n255 10.6151
R957 B.n255 B.n252 10.6151
R958 B.n252 B.n251 10.6151
R959 B.n251 B.n248 10.6151
R960 B.n248 B.n247 10.6151
R961 B.n247 B.n244 10.6151
R962 B.n244 B.n243 10.6151
R963 B.n243 B.n240 10.6151
R964 B.n240 B.n239 10.6151
R965 B.n239 B.n236 10.6151
R966 B.n236 B.n235 10.6151
R967 B.n235 B.n233 10.6151
R968 B.n316 B.n201 10.6151
R969 B.n317 B.n316 10.6151
R970 B.n318 B.n317 10.6151
R971 B.n318 B.n193 10.6151
R972 B.n328 B.n193 10.6151
R973 B.n329 B.n328 10.6151
R974 B.n330 B.n329 10.6151
R975 B.n330 B.n185 10.6151
R976 B.n340 B.n185 10.6151
R977 B.n341 B.n340 10.6151
R978 B.n342 B.n341 10.6151
R979 B.n342 B.n176 10.6151
R980 B.n352 B.n176 10.6151
R981 B.n353 B.n352 10.6151
R982 B.n354 B.n353 10.6151
R983 B.n354 B.n169 10.6151
R984 B.n364 B.n169 10.6151
R985 B.n365 B.n364 10.6151
R986 B.n366 B.n365 10.6151
R987 B.n366 B.n161 10.6151
R988 B.n376 B.n161 10.6151
R989 B.n377 B.n376 10.6151
R990 B.n379 B.n377 10.6151
R991 B.n379 B.n378 10.6151
R992 B.n378 B.n154 10.6151
R993 B.n391 B.n154 10.6151
R994 B.n392 B.n391 10.6151
R995 B.n393 B.n392 10.6151
R996 B.n394 B.n393 10.6151
R997 B.n395 B.n394 10.6151
R998 B.n398 B.n395 10.6151
R999 B.n399 B.n398 10.6151
R1000 B.n400 B.n399 10.6151
R1001 B.n401 B.n400 10.6151
R1002 B.n403 B.n401 10.6151
R1003 B.n404 B.n403 10.6151
R1004 B.n405 B.n404 10.6151
R1005 B.n406 B.n405 10.6151
R1006 B.n408 B.n406 10.6151
R1007 B.n409 B.n408 10.6151
R1008 B.n410 B.n409 10.6151
R1009 B.n411 B.n410 10.6151
R1010 B.n413 B.n411 10.6151
R1011 B.n414 B.n413 10.6151
R1012 B.n415 B.n414 10.6151
R1013 B.n416 B.n415 10.6151
R1014 B.n418 B.n416 10.6151
R1015 B.n419 B.n418 10.6151
R1016 B.n420 B.n419 10.6151
R1017 B.n421 B.n420 10.6151
R1018 B.n423 B.n421 10.6151
R1019 B.n424 B.n423 10.6151
R1020 B.n425 B.n424 10.6151
R1021 B.n426 B.n425 10.6151
R1022 B.n427 B.n426 10.6151
R1023 B.n484 B.n1 10.6151
R1024 B.n484 B.n483 10.6151
R1025 B.n483 B.n482 10.6151
R1026 B.n482 B.n10 10.6151
R1027 B.n476 B.n10 10.6151
R1028 B.n476 B.n475 10.6151
R1029 B.n475 B.n474 10.6151
R1030 B.n474 B.n18 10.6151
R1031 B.n468 B.n18 10.6151
R1032 B.n468 B.n467 10.6151
R1033 B.n467 B.n466 10.6151
R1034 B.n466 B.n25 10.6151
R1035 B.n460 B.n25 10.6151
R1036 B.n460 B.n459 10.6151
R1037 B.n459 B.n458 10.6151
R1038 B.n458 B.n32 10.6151
R1039 B.n452 B.n32 10.6151
R1040 B.n452 B.n451 10.6151
R1041 B.n451 B.n450 10.6151
R1042 B.n450 B.n39 10.6151
R1043 B.n444 B.n39 10.6151
R1044 B.n444 B.n443 10.6151
R1045 B.n443 B.n442 10.6151
R1046 B.n442 B.n46 10.6151
R1047 B.n436 B.n46 10.6151
R1048 B.n436 B.n435 10.6151
R1049 B.n434 B.n53 10.6151
R1050 B.n80 B.n53 10.6151
R1051 B.n81 B.n80 10.6151
R1052 B.n84 B.n81 10.6151
R1053 B.n85 B.n84 10.6151
R1054 B.n88 B.n85 10.6151
R1055 B.n89 B.n88 10.6151
R1056 B.n92 B.n89 10.6151
R1057 B.n93 B.n92 10.6151
R1058 B.n96 B.n93 10.6151
R1059 B.n97 B.n96 10.6151
R1060 B.n100 B.n97 10.6151
R1061 B.n101 B.n100 10.6151
R1062 B.n104 B.n101 10.6151
R1063 B.n109 B.n106 10.6151
R1064 B.n110 B.n109 10.6151
R1065 B.n113 B.n110 10.6151
R1066 B.n114 B.n113 10.6151
R1067 B.n117 B.n114 10.6151
R1068 B.n118 B.n117 10.6151
R1069 B.n121 B.n118 10.6151
R1070 B.n122 B.n121 10.6151
R1071 B.n125 B.n122 10.6151
R1072 B.n130 B.n127 10.6151
R1073 B.n131 B.n130 10.6151
R1074 B.n134 B.n131 10.6151
R1075 B.n135 B.n134 10.6151
R1076 B.n138 B.n135 10.6151
R1077 B.n139 B.n138 10.6151
R1078 B.n142 B.n139 10.6151
R1079 B.n143 B.n142 10.6151
R1080 B.n146 B.n143 10.6151
R1081 B.n147 B.n146 10.6151
R1082 B.n150 B.n147 10.6151
R1083 B.n152 B.n150 10.6151
R1084 B.n153 B.n152 10.6151
R1085 B.n428 B.n153 10.6151
R1086 B.t3 B.n167 10.508
R1087 B.n471 B.t1 10.508
R1088 B.n283 B.n229 9.36635
R1089 B.n260 B.n232 9.36635
R1090 B.n105 B.n104 9.36635
R1091 B.n127 B.n126 9.36635
R1092 B.n492 B.n0 8.11757
R1093 B.n492 B.n1 8.11757
R1094 B.n374 B.t8 7.8811
R1095 B.t9 B.n478 7.8811
R1096 B.n326 B.t15 5.25423
R1097 B.t11 B.n446 5.25423
R1098 B.n280 B.n229 1.24928
R1099 B.n263 B.n232 1.24928
R1100 B.n106 B.n105 1.24928
R1101 B.n126 B.n125 1.24928
R1102 VN.n3 VN.t9 170.805
R1103 VN.n13 VN.t7 170.805
R1104 VN.n9 VN.n8 161.3
R1105 VN.n19 VN.n18 161.3
R1106 VN.n17 VN.n10 161.3
R1107 VN.n7 VN.n0 161.3
R1108 VN.n2 VN.t2 149.992
R1109 VN.n1 VN.t6 149.992
R1110 VN.n6 VN.t5 149.992
R1111 VN.n8 VN.t3 149.992
R1112 VN.n12 VN.t1 149.992
R1113 VN.n11 VN.t8 149.992
R1114 VN.n16 VN.t4 149.992
R1115 VN.n18 VN.t0 149.992
R1116 VN.n16 VN.n15 80.6037
R1117 VN.n14 VN.n11 80.6037
R1118 VN.n6 VN.n5 80.6037
R1119 VN.n4 VN.n1 80.6037
R1120 VN.n2 VN.n1 48.2005
R1121 VN.n6 VN.n1 48.2005
R1122 VN.n12 VN.n11 48.2005
R1123 VN.n16 VN.n11 48.2005
R1124 VN.n7 VN.n6 40.8975
R1125 VN.n17 VN.n16 40.8975
R1126 VN VN.n19 36.6653
R1127 VN.n14 VN.n13 31.6317
R1128 VN.n4 VN.n3 31.6317
R1129 VN.n3 VN.n2 17.5473
R1130 VN.n13 VN.n12 17.5473
R1131 VN.n8 VN.n7 7.30353
R1132 VN.n18 VN.n17 7.30353
R1133 VN.n15 VN.n14 0.380177
R1134 VN.n5 VN.n4 0.380177
R1135 VN.n15 VN.n10 0.285035
R1136 VN.n5 VN.n0 0.285035
R1137 VN.n19 VN.n10 0.189894
R1138 VN.n9 VN.n0 0.189894
R1139 VN VN.n9 0.0516364
R1140 VDD2.n29 VDD2.n19 289.615
R1141 VDD2.n10 VDD2.n0 289.615
R1142 VDD2.n30 VDD2.n29 185
R1143 VDD2.n28 VDD2.n27 185
R1144 VDD2.n23 VDD2.n22 185
R1145 VDD2.n4 VDD2.n3 185
R1146 VDD2.n9 VDD2.n8 185
R1147 VDD2.n11 VDD2.n10 185
R1148 VDD2.n24 VDD2.t9 148.606
R1149 VDD2.n5 VDD2.t0 148.606
R1150 VDD2.n29 VDD2.n28 104.615
R1151 VDD2.n28 VDD2.n22 104.615
R1152 VDD2.n9 VDD2.n3 104.615
R1153 VDD2.n10 VDD2.n9 104.615
R1154 VDD2.n18 VDD2.n17 78.0106
R1155 VDD2 VDD2.n37 78.0077
R1156 VDD2.n36 VDD2.n35 77.3613
R1157 VDD2.n16 VDD2.n15 77.3612
R1158 VDD2.t9 VDD2.n22 52.3082
R1159 VDD2.t0 VDD2.n3 52.3082
R1160 VDD2.n16 VDD2.n14 49.4159
R1161 VDD2.n34 VDD2.n33 48.4763
R1162 VDD2.n34 VDD2.n18 30.8511
R1163 VDD2.n24 VDD2.n23 15.5966
R1164 VDD2.n5 VDD2.n4 15.5966
R1165 VDD2.n27 VDD2.n26 12.8005
R1166 VDD2.n8 VDD2.n7 12.8005
R1167 VDD2.n30 VDD2.n21 12.0247
R1168 VDD2.n11 VDD2.n2 12.0247
R1169 VDD2.n31 VDD2.n19 11.249
R1170 VDD2.n12 VDD2.n0 11.249
R1171 VDD2.n33 VDD2.n32 9.45567
R1172 VDD2.n14 VDD2.n13 9.45567
R1173 VDD2.n32 VDD2.n31 9.3005
R1174 VDD2.n21 VDD2.n20 9.3005
R1175 VDD2.n26 VDD2.n25 9.3005
R1176 VDD2.n13 VDD2.n12 9.3005
R1177 VDD2.n2 VDD2.n1 9.3005
R1178 VDD2.n7 VDD2.n6 9.3005
R1179 VDD2.n37 VDD2.t8 6.3876
R1180 VDD2.n37 VDD2.t2 6.3876
R1181 VDD2.n35 VDD2.t5 6.3876
R1182 VDD2.n35 VDD2.t1 6.3876
R1183 VDD2.n17 VDD2.t4 6.3876
R1184 VDD2.n17 VDD2.t6 6.3876
R1185 VDD2.n15 VDD2.t7 6.3876
R1186 VDD2.n15 VDD2.t3 6.3876
R1187 VDD2.n25 VDD2.n24 4.46457
R1188 VDD2.n6 VDD2.n5 4.46457
R1189 VDD2.n33 VDD2.n19 2.71565
R1190 VDD2.n14 VDD2.n0 2.71565
R1191 VDD2.n31 VDD2.n30 1.93989
R1192 VDD2.n12 VDD2.n11 1.93989
R1193 VDD2.n27 VDD2.n21 1.16414
R1194 VDD2.n8 VDD2.n2 1.16414
R1195 VDD2.n36 VDD2.n34 0.940155
R1196 VDD2.n26 VDD2.n23 0.388379
R1197 VDD2.n7 VDD2.n4 0.388379
R1198 VDD2 VDD2.n36 0.293603
R1199 VDD2.n18 VDD2.n16 0.180068
R1200 VDD2.n32 VDD2.n20 0.155672
R1201 VDD2.n25 VDD2.n20 0.155672
R1202 VDD2.n6 VDD2.n1 0.155672
R1203 VDD2.n13 VDD2.n1 0.155672
C0 VDD2 VP 0.353895f
C1 VN VP 4.04454f
C2 VDD1 VTAIL 5.46491f
C3 VDD2 VTAIL 5.50452f
C4 VN VTAIL 2.44545f
C5 VDD2 VDD1 1.00788f
C6 VN VDD1 0.154611f
C7 VP VTAIL 2.45969f
C8 VDD2 VN 2.12707f
C9 VP VDD1 2.32409f
C10 VDD2 B 3.4321f
C11 VDD1 B 3.379079f
C12 VTAIL B 3.128718f
C13 VN B 8.59223f
C14 VP B 7.046414f
C15 VDD2.n0 B 0.031158f
C16 VDD2.n1 B 0.024264f
C17 VDD2.n2 B 0.013038f
C18 VDD2.n3 B 0.023113f
C19 VDD2.n4 B 0.01797f
C20 VDD2.t0 B 0.051408f
C21 VDD2.n5 B 0.088035f
C22 VDD2.n6 B 0.251814f
C23 VDD2.n7 B 0.013038f
C24 VDD2.n8 B 0.013805f
C25 VDD2.n9 B 0.030818f
C26 VDD2.n10 B 0.061504f
C27 VDD2.n11 B 0.013805f
C28 VDD2.n12 B 0.013038f
C29 VDD2.n13 B 0.055421f
C30 VDD2.n14 B 0.052895f
C31 VDD2.t7 B 0.059439f
C32 VDD2.t3 B 0.059439f
C33 VDD2.n15 B 0.445757f
C34 VDD2.n16 B 0.389717f
C35 VDD2.t4 B 0.059439f
C36 VDD2.t6 B 0.059439f
C37 VDD2.n17 B 0.448391f
C38 VDD2.n18 B 1.35347f
C39 VDD2.n19 B 0.031158f
C40 VDD2.n20 B 0.024264f
C41 VDD2.n21 B 0.013038f
C42 VDD2.n22 B 0.023113f
C43 VDD2.n23 B 0.01797f
C44 VDD2.t9 B 0.051408f
C45 VDD2.n24 B 0.088035f
C46 VDD2.n25 B 0.251814f
C47 VDD2.n26 B 0.013038f
C48 VDD2.n27 B 0.013805f
C49 VDD2.n28 B 0.030818f
C50 VDD2.n29 B 0.061504f
C51 VDD2.n30 B 0.013805f
C52 VDD2.n31 B 0.013038f
C53 VDD2.n32 B 0.055421f
C54 VDD2.n33 B 0.050617f
C55 VDD2.n34 B 1.42094f
C56 VDD2.t5 B 0.059439f
C57 VDD2.t1 B 0.059439f
C58 VDD2.n35 B 0.445759f
C59 VDD2.n36 B 0.27793f
C60 VDD2.t8 B 0.059439f
C61 VDD2.t2 B 0.059439f
C62 VDD2.n37 B 0.448371f
C63 VN.n0 B 0.057619f
C64 VN.t6 B 0.304418f
C65 VN.n1 B 0.184835f
C66 VN.t9 B 0.325793f
C67 VN.t2 B 0.304418f
C68 VN.n2 B 0.18429f
C69 VN.n3 B 0.157753f
C70 VN.n4 B 0.259744f
C71 VN.n5 B 0.071923f
C72 VN.t5 B 0.304418f
C73 VN.n6 B 0.183504f
C74 VN.n7 B 0.009799f
C75 VN.t3 B 0.304418f
C76 VN.n8 B 0.167582f
C77 VN.n9 B 0.033463f
C78 VN.n10 B 0.057619f
C79 VN.t8 B 0.304418f
C80 VN.n11 B 0.184835f
C81 VN.t4 B 0.304418f
C82 VN.t7 B 0.325793f
C83 VN.t1 B 0.304418f
C84 VN.n12 B 0.18429f
C85 VN.n13 B 0.157753f
C86 VN.n14 B 0.259744f
C87 VN.n15 B 0.071923f
C88 VN.n16 B 0.183504f
C89 VN.n17 B 0.009799f
C90 VN.t0 B 0.304418f
C91 VN.n18 B 0.167582f
C92 VN.n19 B 1.40631f
C93 VTAIL.t0 B 0.073859f
C94 VTAIL.t17 B 0.073859f
C95 VTAIL.n0 B 0.493475f
C96 VTAIL.n1 B 0.410456f
C97 VTAIL.n2 B 0.038717f
C98 VTAIL.n3 B 0.03015f
C99 VTAIL.n4 B 0.016201f
C100 VTAIL.n5 B 0.028721f
C101 VTAIL.n6 B 0.02233f
C102 VTAIL.t12 B 0.06388f
C103 VTAIL.n7 B 0.109393f
C104 VTAIL.n8 B 0.312908f
C105 VTAIL.n9 B 0.016201f
C106 VTAIL.n10 B 0.017154f
C107 VTAIL.n11 B 0.038294f
C108 VTAIL.n12 B 0.076426f
C109 VTAIL.n13 B 0.017154f
C110 VTAIL.n14 B 0.016201f
C111 VTAIL.n15 B 0.068867f
C112 VTAIL.n16 B 0.042072f
C113 VTAIL.n17 B 0.207862f
C114 VTAIL.t9 B 0.073859f
C115 VTAIL.t13 B 0.073859f
C116 VTAIL.n18 B 0.493475f
C117 VTAIL.n19 B 0.427625f
C118 VTAIL.t8 B 0.073859f
C119 VTAIL.t11 B 0.073859f
C120 VTAIL.n20 B 0.493475f
C121 VTAIL.n21 B 1.1881f
C122 VTAIL.t4 B 0.073859f
C123 VTAIL.t18 B 0.073859f
C124 VTAIL.n22 B 0.493478f
C125 VTAIL.n23 B 1.18809f
C126 VTAIL.t3 B 0.073859f
C127 VTAIL.t19 B 0.073859f
C128 VTAIL.n24 B 0.493478f
C129 VTAIL.n25 B 0.427622f
C130 VTAIL.n26 B 0.038717f
C131 VTAIL.n27 B 0.03015f
C132 VTAIL.n28 B 0.016201f
C133 VTAIL.n29 B 0.028721f
C134 VTAIL.n30 B 0.02233f
C135 VTAIL.t2 B 0.06388f
C136 VTAIL.n31 B 0.109393f
C137 VTAIL.n32 B 0.312908f
C138 VTAIL.n33 B 0.016201f
C139 VTAIL.n34 B 0.017154f
C140 VTAIL.n35 B 0.038294f
C141 VTAIL.n36 B 0.076426f
C142 VTAIL.n37 B 0.017154f
C143 VTAIL.n38 B 0.016201f
C144 VTAIL.n39 B 0.068867f
C145 VTAIL.n40 B 0.042072f
C146 VTAIL.n41 B 0.207862f
C147 VTAIL.t14 B 0.073859f
C148 VTAIL.t16 B 0.073859f
C149 VTAIL.n42 B 0.493478f
C150 VTAIL.n43 B 0.427622f
C151 VTAIL.t7 B 0.073859f
C152 VTAIL.t15 B 0.073859f
C153 VTAIL.n44 B 0.493478f
C154 VTAIL.n45 B 0.427622f
C155 VTAIL.n46 B 0.038717f
C156 VTAIL.n47 B 0.03015f
C157 VTAIL.n48 B 0.016201f
C158 VTAIL.n49 B 0.028721f
C159 VTAIL.n50 B 0.02233f
C160 VTAIL.t10 B 0.06388f
C161 VTAIL.n51 B 0.109393f
C162 VTAIL.n52 B 0.312908f
C163 VTAIL.n53 B 0.016201f
C164 VTAIL.n54 B 0.017154f
C165 VTAIL.n55 B 0.038294f
C166 VTAIL.n56 B 0.076426f
C167 VTAIL.n57 B 0.017154f
C168 VTAIL.n58 B 0.016201f
C169 VTAIL.n59 B 0.068867f
C170 VTAIL.n60 B 0.042072f
C171 VTAIL.n61 B 0.877046f
C172 VTAIL.n62 B 0.038717f
C173 VTAIL.n63 B 0.03015f
C174 VTAIL.n64 B 0.016201f
C175 VTAIL.n65 B 0.028721f
C176 VTAIL.n66 B 0.02233f
C177 VTAIL.t5 B 0.06388f
C178 VTAIL.n67 B 0.109393f
C179 VTAIL.n68 B 0.312908f
C180 VTAIL.n69 B 0.016201f
C181 VTAIL.n70 B 0.017154f
C182 VTAIL.n71 B 0.038294f
C183 VTAIL.n72 B 0.076426f
C184 VTAIL.n73 B 0.017154f
C185 VTAIL.n74 B 0.016201f
C186 VTAIL.n75 B 0.068867f
C187 VTAIL.n76 B 0.042072f
C188 VTAIL.n77 B 0.877046f
C189 VTAIL.t1 B 0.073859f
C190 VTAIL.t6 B 0.073859f
C191 VTAIL.n78 B 0.493475f
C192 VTAIL.n79 B 0.353506f
C193 VDD1.n0 B 0.031605f
C194 VDD1.n1 B 0.024612f
C195 VDD1.n2 B 0.013225f
C196 VDD1.n3 B 0.023445f
C197 VDD1.n4 B 0.018228f
C198 VDD1.t8 B 0.052146f
C199 VDD1.n5 B 0.089299f
C200 VDD1.n6 B 0.255429f
C201 VDD1.n7 B 0.013225f
C202 VDD1.n8 B 0.014003f
C203 VDD1.n9 B 0.03126f
C204 VDD1.n10 B 0.062387f
C205 VDD1.n11 B 0.014003f
C206 VDD1.n12 B 0.013225f
C207 VDD1.n13 B 0.056217f
C208 VDD1.n14 B 0.053654f
C209 VDD1.t3 B 0.060292f
C210 VDD1.t9 B 0.060292f
C211 VDD1.n15 B 0.452158f
C212 VDD1.n16 B 0.401135f
C213 VDD1.n17 B 0.031605f
C214 VDD1.n18 B 0.024612f
C215 VDD1.n19 B 0.013225f
C216 VDD1.n20 B 0.023445f
C217 VDD1.n21 B 0.018228f
C218 VDD1.t0 B 0.052146f
C219 VDD1.n22 B 0.089299f
C220 VDD1.n23 B 0.255429f
C221 VDD1.n24 B 0.013225f
C222 VDD1.n25 B 0.014003f
C223 VDD1.n26 B 0.03126f
C224 VDD1.n27 B 0.062387f
C225 VDD1.n28 B 0.014003f
C226 VDD1.n29 B 0.013225f
C227 VDD1.n30 B 0.056217f
C228 VDD1.n31 B 0.053654f
C229 VDD1.t4 B 0.060292f
C230 VDD1.t2 B 0.060292f
C231 VDD1.n32 B 0.452156f
C232 VDD1.n33 B 0.395311f
C233 VDD1.t5 B 0.060292f
C234 VDD1.t1 B 0.060292f
C235 VDD1.n34 B 0.454828f
C236 VDD1.n35 B 1.44586f
C237 VDD1.t6 B 0.060292f
C238 VDD1.t7 B 0.060292f
C239 VDD1.n36 B 0.452156f
C240 VDD1.n37 B 1.65762f
C241 VP.n0 B 0.060082f
C242 VP.t7 B 0.317429f
C243 VP.n1 B 0.192735f
C244 VP.n2 B 0.060082f
C245 VP.n3 B 0.060082f
C246 VP.t6 B 0.317429f
C247 VP.t1 B 0.317429f
C248 VP.n4 B 0.074997f
C249 VP.t9 B 0.317429f
C250 VP.n5 B 0.270845f
C251 VP.t0 B 0.317429f
C252 VP.t2 B 0.339718f
C253 VP.n6 B 0.164496f
C254 VP.n7 B 0.192167f
C255 VP.n8 B 0.192735f
C256 VP.n9 B 0.191347f
C257 VP.n10 B 0.010217f
C258 VP.n11 B 0.174745f
C259 VP.n12 B 1.43657f
C260 VP.n13 B 1.4813f
C261 VP.t8 B 0.317429f
C262 VP.n14 B 0.174745f
C263 VP.n15 B 0.010217f
C264 VP.t5 B 0.317429f
C265 VP.n16 B 0.191347f
C266 VP.n17 B 0.074997f
C267 VP.n18 B 0.090052f
C268 VP.n19 B 0.074997f
C269 VP.t3 B 0.317429f
C270 VP.n20 B 0.191347f
C271 VP.n21 B 0.010217f
C272 VP.t4 B 0.317429f
C273 VP.n22 B 0.174745f
C274 VP.n23 B 0.034894f
.ends

