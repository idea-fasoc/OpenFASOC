* NGSPICE file created from diff_pair_sample_1139.ext - technology: sky130A

.subckt diff_pair_sample_1139 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0.9405 ps=6.03 w=5.7 l=2.05
X1 VDD1.t9 VP.t0 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0.9405 ps=6.03 w=5.7 l=2.05
X2 VDD2.t8 VN.t1 VTAIL.t19 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X3 VDD1.t8 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0.9405 ps=6.03 w=5.7 l=2.05
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0 ps=0 w=5.7 l=2.05
X5 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0 ps=0 w=5.7 l=2.05
X6 VTAIL.t4 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X7 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0 ps=0 w=5.7 l=2.05
X8 VDD1.t6 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=2.223 ps=12.18 w=5.7 l=2.05
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0 ps=0 w=5.7 l=2.05
X10 VTAIL.t11 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X11 VDD2.t6 VN.t3 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.223 pd=12.18 as=0.9405 ps=6.03 w=5.7 l=2.05
X12 VTAIL.t16 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X13 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X14 VDD1.t4 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X15 VDD2.t4 VN.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=2.223 ps=12.18 w=5.7 l=2.05
X16 VTAIL.t5 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X17 VDD2.t3 VN.t6 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X18 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=2.223 ps=12.18 w=5.7 l=2.05
X19 VTAIL.t9 VP.t8 VDD1.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X20 VTAIL.t7 VP.t9 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X21 VTAIL.t15 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X22 VTAIL.t13 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=0.9405 ps=6.03 w=5.7 l=2.05
X23 VDD2.t0 VN.t9 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9405 pd=6.03 as=2.223 ps=12.18 w=5.7 l=2.05
R0 VN.n35 VN.n34 185.4
R1 VN.n71 VN.n70 185.4
R2 VN.n69 VN.n36 161.3
R3 VN.n68 VN.n67 161.3
R4 VN.n66 VN.n37 161.3
R5 VN.n65 VN.n64 161.3
R6 VN.n63 VN.n38 161.3
R7 VN.n61 VN.n60 161.3
R8 VN.n59 VN.n39 161.3
R9 VN.n58 VN.n57 161.3
R10 VN.n56 VN.n40 161.3
R11 VN.n55 VN.n54 161.3
R12 VN.n53 VN.n52 161.3
R13 VN.n51 VN.n42 161.3
R14 VN.n50 VN.n49 161.3
R15 VN.n48 VN.n43 161.3
R16 VN.n47 VN.n46 161.3
R17 VN.n33 VN.n0 161.3
R18 VN.n32 VN.n31 161.3
R19 VN.n30 VN.n1 161.3
R20 VN.n29 VN.n28 161.3
R21 VN.n27 VN.n2 161.3
R22 VN.n25 VN.n24 161.3
R23 VN.n23 VN.n3 161.3
R24 VN.n22 VN.n21 161.3
R25 VN.n20 VN.n4 161.3
R26 VN.n19 VN.n18 161.3
R27 VN.n17 VN.n16 161.3
R28 VN.n15 VN.n6 161.3
R29 VN.n14 VN.n13 161.3
R30 VN.n12 VN.n7 161.3
R31 VN.n11 VN.n10 161.3
R32 VN.n8 VN.t0 98.5
R33 VN.n44 VN.t5 98.5
R34 VN.n9 VN.t4 67.0103
R35 VN.n5 VN.t6 67.0103
R36 VN.n26 VN.t7 67.0103
R37 VN.n34 VN.t9 67.0103
R38 VN.n45 VN.t8 67.0103
R39 VN.n41 VN.t1 67.0103
R40 VN.n62 VN.t2 67.0103
R41 VN.n70 VN.t3 67.0103
R42 VN.n9 VN.n8 64.2931
R43 VN.n45 VN.n44 64.2931
R44 VN.n28 VN.n1 56.5617
R45 VN.n64 VN.n37 56.5617
R46 VN.n15 VN.n14 46.3896
R47 VN.n21 VN.n20 46.3896
R48 VN.n51 VN.n50 46.3896
R49 VN.n57 VN.n56 46.3896
R50 VN VN.n71 45.6463
R51 VN.n14 VN.n7 34.7644
R52 VN.n21 VN.n3 34.7644
R53 VN.n50 VN.n43 34.7644
R54 VN.n57 VN.n39 34.7644
R55 VN.n10 VN.n7 24.5923
R56 VN.n16 VN.n15 24.5923
R57 VN.n20 VN.n19 24.5923
R58 VN.n25 VN.n3 24.5923
R59 VN.n28 VN.n27 24.5923
R60 VN.n32 VN.n1 24.5923
R61 VN.n33 VN.n32 24.5923
R62 VN.n46 VN.n43 24.5923
R63 VN.n56 VN.n55 24.5923
R64 VN.n52 VN.n51 24.5923
R65 VN.n64 VN.n63 24.5923
R66 VN.n61 VN.n39 24.5923
R67 VN.n69 VN.n68 24.5923
R68 VN.n68 VN.n37 24.5923
R69 VN.n27 VN.n26 18.1985
R70 VN.n63 VN.n62 18.1985
R71 VN.n47 VN.n44 12.6154
R72 VN.n11 VN.n8 12.6154
R73 VN.n16 VN.n5 12.2964
R74 VN.n19 VN.n5 12.2964
R75 VN.n55 VN.n41 12.2964
R76 VN.n52 VN.n41 12.2964
R77 VN.n10 VN.n9 6.39438
R78 VN.n26 VN.n25 6.39438
R79 VN.n46 VN.n45 6.39438
R80 VN.n62 VN.n61 6.39438
R81 VN.n34 VN.n33 0.492337
R82 VN.n70 VN.n69 0.492337
R83 VN.n71 VN.n36 0.189894
R84 VN.n67 VN.n36 0.189894
R85 VN.n67 VN.n66 0.189894
R86 VN.n66 VN.n65 0.189894
R87 VN.n65 VN.n38 0.189894
R88 VN.n60 VN.n38 0.189894
R89 VN.n60 VN.n59 0.189894
R90 VN.n59 VN.n58 0.189894
R91 VN.n58 VN.n40 0.189894
R92 VN.n54 VN.n40 0.189894
R93 VN.n54 VN.n53 0.189894
R94 VN.n53 VN.n42 0.189894
R95 VN.n49 VN.n42 0.189894
R96 VN.n49 VN.n48 0.189894
R97 VN.n48 VN.n47 0.189894
R98 VN.n12 VN.n11 0.189894
R99 VN.n13 VN.n12 0.189894
R100 VN.n13 VN.n6 0.189894
R101 VN.n17 VN.n6 0.189894
R102 VN.n18 VN.n17 0.189894
R103 VN.n18 VN.n4 0.189894
R104 VN.n22 VN.n4 0.189894
R105 VN.n23 VN.n22 0.189894
R106 VN.n24 VN.n23 0.189894
R107 VN.n24 VN.n2 0.189894
R108 VN.n29 VN.n2 0.189894
R109 VN.n30 VN.n29 0.189894
R110 VN.n31 VN.n30 0.189894
R111 VN.n31 VN.n0 0.189894
R112 VN.n35 VN.n0 0.189894
R113 VN VN.n35 0.0516364
R114 VTAIL.n11 VTAIL.t10 55.8285
R115 VTAIL.n17 VTAIL.t12 55.8283
R116 VTAIL.n2 VTAIL.t6 55.8283
R117 VTAIL.n16 VTAIL.t1 55.8283
R118 VTAIL.n15 VTAIL.n14 52.3549
R119 VTAIL.n13 VTAIL.n12 52.3549
R120 VTAIL.n10 VTAIL.n9 52.3549
R121 VTAIL.n8 VTAIL.n7 52.3549
R122 VTAIL.n19 VTAIL.n18 52.3547
R123 VTAIL.n1 VTAIL.n0 52.3547
R124 VTAIL.n4 VTAIL.n3 52.3547
R125 VTAIL.n6 VTAIL.n5 52.3547
R126 VTAIL.n8 VTAIL.n6 21.3841
R127 VTAIL.n17 VTAIL.n16 19.3324
R128 VTAIL.n18 VTAIL.t17 3.47418
R129 VTAIL.n18 VTAIL.t15 3.47418
R130 VTAIL.n0 VTAIL.t18 3.47418
R131 VTAIL.n0 VTAIL.t16 3.47418
R132 VTAIL.n3 VTAIL.t2 3.47418
R133 VTAIL.n3 VTAIL.t7 3.47418
R134 VTAIL.n5 VTAIL.t0 3.47418
R135 VTAIL.n5 VTAIL.t9 3.47418
R136 VTAIL.n14 VTAIL.t3 3.47418
R137 VTAIL.n14 VTAIL.t5 3.47418
R138 VTAIL.n12 VTAIL.t8 3.47418
R139 VTAIL.n12 VTAIL.t4 3.47418
R140 VTAIL.n9 VTAIL.t19 3.47418
R141 VTAIL.n9 VTAIL.t13 3.47418
R142 VTAIL.n7 VTAIL.t14 3.47418
R143 VTAIL.n7 VTAIL.t11 3.47418
R144 VTAIL.n10 VTAIL.n8 2.05222
R145 VTAIL.n11 VTAIL.n10 2.05222
R146 VTAIL.n15 VTAIL.n13 2.05222
R147 VTAIL.n16 VTAIL.n15 2.05222
R148 VTAIL.n6 VTAIL.n4 2.05222
R149 VTAIL.n4 VTAIL.n2 2.05222
R150 VTAIL.n19 VTAIL.n17 2.05222
R151 VTAIL VTAIL.n1 1.59748
R152 VTAIL.n13 VTAIL.n11 1.49619
R153 VTAIL.n2 VTAIL.n1 1.49619
R154 VTAIL VTAIL.n19 0.455241
R155 VDD2.n1 VDD2.t9 74.5589
R156 VDD2.n4 VDD2.t6 72.5073
R157 VDD2.n3 VDD2.n2 70.5169
R158 VDD2 VDD2.n7 70.5141
R159 VDD2.n6 VDD2.n5 69.0337
R160 VDD2.n1 VDD2.n0 69.0334
R161 VDD2.n4 VDD2.n3 38.3748
R162 VDD2.n7 VDD2.t1 3.47418
R163 VDD2.n7 VDD2.t4 3.47418
R164 VDD2.n5 VDD2.t7 3.47418
R165 VDD2.n5 VDD2.t8 3.47418
R166 VDD2.n2 VDD2.t2 3.47418
R167 VDD2.n2 VDD2.t0 3.47418
R168 VDD2.n0 VDD2.t5 3.47418
R169 VDD2.n0 VDD2.t3 3.47418
R170 VDD2.n6 VDD2.n4 2.05222
R171 VDD2 VDD2.n6 0.571621
R172 VDD2.n3 VDD2.n1 0.458085
R173 B.n583 B.n582 585
R174 B.n585 B.n125 585
R175 B.n588 B.n587 585
R176 B.n589 B.n124 585
R177 B.n591 B.n590 585
R178 B.n593 B.n123 585
R179 B.n596 B.n595 585
R180 B.n597 B.n122 585
R181 B.n599 B.n598 585
R182 B.n601 B.n121 585
R183 B.n604 B.n603 585
R184 B.n605 B.n120 585
R185 B.n607 B.n606 585
R186 B.n609 B.n119 585
R187 B.n612 B.n611 585
R188 B.n613 B.n118 585
R189 B.n615 B.n614 585
R190 B.n617 B.n117 585
R191 B.n620 B.n619 585
R192 B.n621 B.n116 585
R193 B.n623 B.n622 585
R194 B.n625 B.n115 585
R195 B.n628 B.n627 585
R196 B.n630 B.n112 585
R197 B.n632 B.n631 585
R198 B.n634 B.n111 585
R199 B.n637 B.n636 585
R200 B.n638 B.n110 585
R201 B.n640 B.n639 585
R202 B.n642 B.n109 585
R203 B.n645 B.n644 585
R204 B.n646 B.n105 585
R205 B.n648 B.n647 585
R206 B.n650 B.n104 585
R207 B.n653 B.n652 585
R208 B.n654 B.n103 585
R209 B.n656 B.n655 585
R210 B.n658 B.n102 585
R211 B.n661 B.n660 585
R212 B.n662 B.n101 585
R213 B.n664 B.n663 585
R214 B.n666 B.n100 585
R215 B.n669 B.n668 585
R216 B.n670 B.n99 585
R217 B.n672 B.n671 585
R218 B.n674 B.n98 585
R219 B.n677 B.n676 585
R220 B.n678 B.n97 585
R221 B.n680 B.n679 585
R222 B.n682 B.n96 585
R223 B.n685 B.n684 585
R224 B.n686 B.n95 585
R225 B.n688 B.n687 585
R226 B.n690 B.n94 585
R227 B.n693 B.n692 585
R228 B.n694 B.n93 585
R229 B.n581 B.n91 585
R230 B.n697 B.n91 585
R231 B.n580 B.n90 585
R232 B.n698 B.n90 585
R233 B.n579 B.n89 585
R234 B.n699 B.n89 585
R235 B.n578 B.n577 585
R236 B.n577 B.n85 585
R237 B.n576 B.n84 585
R238 B.n705 B.n84 585
R239 B.n575 B.n83 585
R240 B.n706 B.n83 585
R241 B.n574 B.n82 585
R242 B.n707 B.n82 585
R243 B.n573 B.n572 585
R244 B.n572 B.n78 585
R245 B.n571 B.n77 585
R246 B.n713 B.n77 585
R247 B.n570 B.n76 585
R248 B.n714 B.n76 585
R249 B.n569 B.n75 585
R250 B.n715 B.n75 585
R251 B.n568 B.n567 585
R252 B.n567 B.n71 585
R253 B.n566 B.n70 585
R254 B.n721 B.n70 585
R255 B.n565 B.n69 585
R256 B.n722 B.n69 585
R257 B.n564 B.n68 585
R258 B.n723 B.n68 585
R259 B.n563 B.n562 585
R260 B.n562 B.n64 585
R261 B.n561 B.n63 585
R262 B.n729 B.n63 585
R263 B.n560 B.n62 585
R264 B.n730 B.n62 585
R265 B.n559 B.n61 585
R266 B.n731 B.n61 585
R267 B.n558 B.n557 585
R268 B.n557 B.n57 585
R269 B.n556 B.n56 585
R270 B.n737 B.n56 585
R271 B.n555 B.n55 585
R272 B.n738 B.n55 585
R273 B.n554 B.n54 585
R274 B.n739 B.n54 585
R275 B.n553 B.n552 585
R276 B.n552 B.n53 585
R277 B.n551 B.n49 585
R278 B.n745 B.n49 585
R279 B.n550 B.n48 585
R280 B.n746 B.n48 585
R281 B.n549 B.n47 585
R282 B.n747 B.n47 585
R283 B.n548 B.n547 585
R284 B.n547 B.n43 585
R285 B.n546 B.n42 585
R286 B.n753 B.n42 585
R287 B.n545 B.n41 585
R288 B.n754 B.n41 585
R289 B.n544 B.n40 585
R290 B.n755 B.n40 585
R291 B.n543 B.n542 585
R292 B.n542 B.n36 585
R293 B.n541 B.n35 585
R294 B.n761 B.n35 585
R295 B.n540 B.n34 585
R296 B.n762 B.n34 585
R297 B.n539 B.n33 585
R298 B.n763 B.n33 585
R299 B.n538 B.n537 585
R300 B.n537 B.n29 585
R301 B.n536 B.n28 585
R302 B.n769 B.n28 585
R303 B.n535 B.n27 585
R304 B.n770 B.n27 585
R305 B.n534 B.n26 585
R306 B.n771 B.n26 585
R307 B.n533 B.n532 585
R308 B.n532 B.n22 585
R309 B.n531 B.n21 585
R310 B.n777 B.n21 585
R311 B.n530 B.n20 585
R312 B.n778 B.n20 585
R313 B.n529 B.n19 585
R314 B.n779 B.n19 585
R315 B.n528 B.n527 585
R316 B.n527 B.n15 585
R317 B.n526 B.n14 585
R318 B.n785 B.n14 585
R319 B.n525 B.n13 585
R320 B.n786 B.n13 585
R321 B.n524 B.n12 585
R322 B.n787 B.n12 585
R323 B.n523 B.n522 585
R324 B.n522 B.n8 585
R325 B.n521 B.n7 585
R326 B.n793 B.n7 585
R327 B.n520 B.n6 585
R328 B.n794 B.n6 585
R329 B.n519 B.n5 585
R330 B.n795 B.n5 585
R331 B.n518 B.n517 585
R332 B.n517 B.n4 585
R333 B.n516 B.n126 585
R334 B.n516 B.n515 585
R335 B.n506 B.n127 585
R336 B.n128 B.n127 585
R337 B.n508 B.n507 585
R338 B.n509 B.n508 585
R339 B.n505 B.n133 585
R340 B.n133 B.n132 585
R341 B.n504 B.n503 585
R342 B.n503 B.n502 585
R343 B.n135 B.n134 585
R344 B.n136 B.n135 585
R345 B.n495 B.n494 585
R346 B.n496 B.n495 585
R347 B.n493 B.n141 585
R348 B.n141 B.n140 585
R349 B.n492 B.n491 585
R350 B.n491 B.n490 585
R351 B.n143 B.n142 585
R352 B.n144 B.n143 585
R353 B.n483 B.n482 585
R354 B.n484 B.n483 585
R355 B.n481 B.n148 585
R356 B.n152 B.n148 585
R357 B.n480 B.n479 585
R358 B.n479 B.n478 585
R359 B.n150 B.n149 585
R360 B.n151 B.n150 585
R361 B.n471 B.n470 585
R362 B.n472 B.n471 585
R363 B.n469 B.n157 585
R364 B.n157 B.n156 585
R365 B.n468 B.n467 585
R366 B.n467 B.n466 585
R367 B.n159 B.n158 585
R368 B.n160 B.n159 585
R369 B.n459 B.n458 585
R370 B.n460 B.n459 585
R371 B.n457 B.n165 585
R372 B.n165 B.n164 585
R373 B.n456 B.n455 585
R374 B.n455 B.n454 585
R375 B.n167 B.n166 585
R376 B.n168 B.n167 585
R377 B.n447 B.n446 585
R378 B.n448 B.n447 585
R379 B.n445 B.n173 585
R380 B.n173 B.n172 585
R381 B.n444 B.n443 585
R382 B.n443 B.n442 585
R383 B.n175 B.n174 585
R384 B.n435 B.n175 585
R385 B.n434 B.n433 585
R386 B.n436 B.n434 585
R387 B.n432 B.n180 585
R388 B.n180 B.n179 585
R389 B.n431 B.n430 585
R390 B.n430 B.n429 585
R391 B.n182 B.n181 585
R392 B.n183 B.n182 585
R393 B.n422 B.n421 585
R394 B.n423 B.n422 585
R395 B.n420 B.n188 585
R396 B.n188 B.n187 585
R397 B.n419 B.n418 585
R398 B.n418 B.n417 585
R399 B.n190 B.n189 585
R400 B.n191 B.n190 585
R401 B.n410 B.n409 585
R402 B.n411 B.n410 585
R403 B.n408 B.n196 585
R404 B.n196 B.n195 585
R405 B.n407 B.n406 585
R406 B.n406 B.n405 585
R407 B.n198 B.n197 585
R408 B.n199 B.n198 585
R409 B.n398 B.n397 585
R410 B.n399 B.n398 585
R411 B.n396 B.n204 585
R412 B.n204 B.n203 585
R413 B.n395 B.n394 585
R414 B.n394 B.n393 585
R415 B.n206 B.n205 585
R416 B.n207 B.n206 585
R417 B.n386 B.n385 585
R418 B.n387 B.n386 585
R419 B.n384 B.n212 585
R420 B.n212 B.n211 585
R421 B.n383 B.n382 585
R422 B.n382 B.n381 585
R423 B.n214 B.n213 585
R424 B.n215 B.n214 585
R425 B.n374 B.n373 585
R426 B.n375 B.n374 585
R427 B.n372 B.n220 585
R428 B.n220 B.n219 585
R429 B.n371 B.n370 585
R430 B.n370 B.n369 585
R431 B.n366 B.n224 585
R432 B.n365 B.n364 585
R433 B.n362 B.n225 585
R434 B.n362 B.n223 585
R435 B.n361 B.n360 585
R436 B.n359 B.n358 585
R437 B.n357 B.n227 585
R438 B.n355 B.n354 585
R439 B.n353 B.n228 585
R440 B.n352 B.n351 585
R441 B.n349 B.n229 585
R442 B.n347 B.n346 585
R443 B.n345 B.n230 585
R444 B.n344 B.n343 585
R445 B.n341 B.n231 585
R446 B.n339 B.n338 585
R447 B.n337 B.n232 585
R448 B.n336 B.n335 585
R449 B.n333 B.n233 585
R450 B.n331 B.n330 585
R451 B.n329 B.n234 585
R452 B.n328 B.n327 585
R453 B.n325 B.n235 585
R454 B.n323 B.n322 585
R455 B.n320 B.n236 585
R456 B.n319 B.n318 585
R457 B.n316 B.n239 585
R458 B.n314 B.n313 585
R459 B.n312 B.n240 585
R460 B.n311 B.n310 585
R461 B.n308 B.n241 585
R462 B.n306 B.n305 585
R463 B.n304 B.n242 585
R464 B.n303 B.n302 585
R465 B.n300 B.n299 585
R466 B.n298 B.n297 585
R467 B.n296 B.n247 585
R468 B.n294 B.n293 585
R469 B.n292 B.n248 585
R470 B.n291 B.n290 585
R471 B.n288 B.n249 585
R472 B.n286 B.n285 585
R473 B.n284 B.n250 585
R474 B.n283 B.n282 585
R475 B.n280 B.n251 585
R476 B.n278 B.n277 585
R477 B.n276 B.n252 585
R478 B.n275 B.n274 585
R479 B.n272 B.n253 585
R480 B.n270 B.n269 585
R481 B.n268 B.n254 585
R482 B.n267 B.n266 585
R483 B.n264 B.n255 585
R484 B.n262 B.n261 585
R485 B.n260 B.n256 585
R486 B.n259 B.n258 585
R487 B.n222 B.n221 585
R488 B.n223 B.n222 585
R489 B.n368 B.n367 585
R490 B.n369 B.n368 585
R491 B.n218 B.n217 585
R492 B.n219 B.n218 585
R493 B.n377 B.n376 585
R494 B.n376 B.n375 585
R495 B.n378 B.n216 585
R496 B.n216 B.n215 585
R497 B.n380 B.n379 585
R498 B.n381 B.n380 585
R499 B.n210 B.n209 585
R500 B.n211 B.n210 585
R501 B.n389 B.n388 585
R502 B.n388 B.n387 585
R503 B.n390 B.n208 585
R504 B.n208 B.n207 585
R505 B.n392 B.n391 585
R506 B.n393 B.n392 585
R507 B.n202 B.n201 585
R508 B.n203 B.n202 585
R509 B.n401 B.n400 585
R510 B.n400 B.n399 585
R511 B.n402 B.n200 585
R512 B.n200 B.n199 585
R513 B.n404 B.n403 585
R514 B.n405 B.n404 585
R515 B.n194 B.n193 585
R516 B.n195 B.n194 585
R517 B.n413 B.n412 585
R518 B.n412 B.n411 585
R519 B.n414 B.n192 585
R520 B.n192 B.n191 585
R521 B.n416 B.n415 585
R522 B.n417 B.n416 585
R523 B.n186 B.n185 585
R524 B.n187 B.n186 585
R525 B.n425 B.n424 585
R526 B.n424 B.n423 585
R527 B.n426 B.n184 585
R528 B.n184 B.n183 585
R529 B.n428 B.n427 585
R530 B.n429 B.n428 585
R531 B.n178 B.n177 585
R532 B.n179 B.n178 585
R533 B.n438 B.n437 585
R534 B.n437 B.n436 585
R535 B.n439 B.n176 585
R536 B.n435 B.n176 585
R537 B.n441 B.n440 585
R538 B.n442 B.n441 585
R539 B.n171 B.n170 585
R540 B.n172 B.n171 585
R541 B.n450 B.n449 585
R542 B.n449 B.n448 585
R543 B.n451 B.n169 585
R544 B.n169 B.n168 585
R545 B.n453 B.n452 585
R546 B.n454 B.n453 585
R547 B.n163 B.n162 585
R548 B.n164 B.n163 585
R549 B.n462 B.n461 585
R550 B.n461 B.n460 585
R551 B.n463 B.n161 585
R552 B.n161 B.n160 585
R553 B.n465 B.n464 585
R554 B.n466 B.n465 585
R555 B.n155 B.n154 585
R556 B.n156 B.n155 585
R557 B.n474 B.n473 585
R558 B.n473 B.n472 585
R559 B.n475 B.n153 585
R560 B.n153 B.n151 585
R561 B.n477 B.n476 585
R562 B.n478 B.n477 585
R563 B.n147 B.n146 585
R564 B.n152 B.n147 585
R565 B.n486 B.n485 585
R566 B.n485 B.n484 585
R567 B.n487 B.n145 585
R568 B.n145 B.n144 585
R569 B.n489 B.n488 585
R570 B.n490 B.n489 585
R571 B.n139 B.n138 585
R572 B.n140 B.n139 585
R573 B.n498 B.n497 585
R574 B.n497 B.n496 585
R575 B.n499 B.n137 585
R576 B.n137 B.n136 585
R577 B.n501 B.n500 585
R578 B.n502 B.n501 585
R579 B.n131 B.n130 585
R580 B.n132 B.n131 585
R581 B.n511 B.n510 585
R582 B.n510 B.n509 585
R583 B.n512 B.n129 585
R584 B.n129 B.n128 585
R585 B.n514 B.n513 585
R586 B.n515 B.n514 585
R587 B.n2 B.n0 585
R588 B.n4 B.n2 585
R589 B.n3 B.n1 585
R590 B.n794 B.n3 585
R591 B.n792 B.n791 585
R592 B.n793 B.n792 585
R593 B.n790 B.n9 585
R594 B.n9 B.n8 585
R595 B.n789 B.n788 585
R596 B.n788 B.n787 585
R597 B.n11 B.n10 585
R598 B.n786 B.n11 585
R599 B.n784 B.n783 585
R600 B.n785 B.n784 585
R601 B.n782 B.n16 585
R602 B.n16 B.n15 585
R603 B.n781 B.n780 585
R604 B.n780 B.n779 585
R605 B.n18 B.n17 585
R606 B.n778 B.n18 585
R607 B.n776 B.n775 585
R608 B.n777 B.n776 585
R609 B.n774 B.n23 585
R610 B.n23 B.n22 585
R611 B.n773 B.n772 585
R612 B.n772 B.n771 585
R613 B.n25 B.n24 585
R614 B.n770 B.n25 585
R615 B.n768 B.n767 585
R616 B.n769 B.n768 585
R617 B.n766 B.n30 585
R618 B.n30 B.n29 585
R619 B.n765 B.n764 585
R620 B.n764 B.n763 585
R621 B.n32 B.n31 585
R622 B.n762 B.n32 585
R623 B.n760 B.n759 585
R624 B.n761 B.n760 585
R625 B.n758 B.n37 585
R626 B.n37 B.n36 585
R627 B.n757 B.n756 585
R628 B.n756 B.n755 585
R629 B.n39 B.n38 585
R630 B.n754 B.n39 585
R631 B.n752 B.n751 585
R632 B.n753 B.n752 585
R633 B.n750 B.n44 585
R634 B.n44 B.n43 585
R635 B.n749 B.n748 585
R636 B.n748 B.n747 585
R637 B.n46 B.n45 585
R638 B.n746 B.n46 585
R639 B.n744 B.n743 585
R640 B.n745 B.n744 585
R641 B.n742 B.n50 585
R642 B.n53 B.n50 585
R643 B.n741 B.n740 585
R644 B.n740 B.n739 585
R645 B.n52 B.n51 585
R646 B.n738 B.n52 585
R647 B.n736 B.n735 585
R648 B.n737 B.n736 585
R649 B.n734 B.n58 585
R650 B.n58 B.n57 585
R651 B.n733 B.n732 585
R652 B.n732 B.n731 585
R653 B.n60 B.n59 585
R654 B.n730 B.n60 585
R655 B.n728 B.n727 585
R656 B.n729 B.n728 585
R657 B.n726 B.n65 585
R658 B.n65 B.n64 585
R659 B.n725 B.n724 585
R660 B.n724 B.n723 585
R661 B.n67 B.n66 585
R662 B.n722 B.n67 585
R663 B.n720 B.n719 585
R664 B.n721 B.n720 585
R665 B.n718 B.n72 585
R666 B.n72 B.n71 585
R667 B.n717 B.n716 585
R668 B.n716 B.n715 585
R669 B.n74 B.n73 585
R670 B.n714 B.n74 585
R671 B.n712 B.n711 585
R672 B.n713 B.n712 585
R673 B.n710 B.n79 585
R674 B.n79 B.n78 585
R675 B.n709 B.n708 585
R676 B.n708 B.n707 585
R677 B.n81 B.n80 585
R678 B.n706 B.n81 585
R679 B.n704 B.n703 585
R680 B.n705 B.n704 585
R681 B.n702 B.n86 585
R682 B.n86 B.n85 585
R683 B.n701 B.n700 585
R684 B.n700 B.n699 585
R685 B.n88 B.n87 585
R686 B.n698 B.n88 585
R687 B.n696 B.n695 585
R688 B.n697 B.n696 585
R689 B.n797 B.n796 585
R690 B.n796 B.n795 585
R691 B.n368 B.n224 497.305
R692 B.n696 B.n93 497.305
R693 B.n370 B.n222 497.305
R694 B.n583 B.n91 497.305
R695 B.n243 B.t18 274.043
R696 B.n237 B.t14 274.043
R697 B.n106 B.t10 274.043
R698 B.n113 B.t21 274.043
R699 B.n584 B.n92 256.663
R700 B.n586 B.n92 256.663
R701 B.n592 B.n92 256.663
R702 B.n594 B.n92 256.663
R703 B.n600 B.n92 256.663
R704 B.n602 B.n92 256.663
R705 B.n608 B.n92 256.663
R706 B.n610 B.n92 256.663
R707 B.n616 B.n92 256.663
R708 B.n618 B.n92 256.663
R709 B.n624 B.n92 256.663
R710 B.n626 B.n92 256.663
R711 B.n633 B.n92 256.663
R712 B.n635 B.n92 256.663
R713 B.n641 B.n92 256.663
R714 B.n643 B.n92 256.663
R715 B.n649 B.n92 256.663
R716 B.n651 B.n92 256.663
R717 B.n657 B.n92 256.663
R718 B.n659 B.n92 256.663
R719 B.n665 B.n92 256.663
R720 B.n667 B.n92 256.663
R721 B.n673 B.n92 256.663
R722 B.n675 B.n92 256.663
R723 B.n681 B.n92 256.663
R724 B.n683 B.n92 256.663
R725 B.n689 B.n92 256.663
R726 B.n691 B.n92 256.663
R727 B.n363 B.n223 256.663
R728 B.n226 B.n223 256.663
R729 B.n356 B.n223 256.663
R730 B.n350 B.n223 256.663
R731 B.n348 B.n223 256.663
R732 B.n342 B.n223 256.663
R733 B.n340 B.n223 256.663
R734 B.n334 B.n223 256.663
R735 B.n332 B.n223 256.663
R736 B.n326 B.n223 256.663
R737 B.n324 B.n223 256.663
R738 B.n317 B.n223 256.663
R739 B.n315 B.n223 256.663
R740 B.n309 B.n223 256.663
R741 B.n307 B.n223 256.663
R742 B.n301 B.n223 256.663
R743 B.n246 B.n223 256.663
R744 B.n295 B.n223 256.663
R745 B.n289 B.n223 256.663
R746 B.n287 B.n223 256.663
R747 B.n281 B.n223 256.663
R748 B.n279 B.n223 256.663
R749 B.n273 B.n223 256.663
R750 B.n271 B.n223 256.663
R751 B.n265 B.n223 256.663
R752 B.n263 B.n223 256.663
R753 B.n257 B.n223 256.663
R754 B.n368 B.n218 163.367
R755 B.n376 B.n218 163.367
R756 B.n376 B.n216 163.367
R757 B.n380 B.n216 163.367
R758 B.n380 B.n210 163.367
R759 B.n388 B.n210 163.367
R760 B.n388 B.n208 163.367
R761 B.n392 B.n208 163.367
R762 B.n392 B.n202 163.367
R763 B.n400 B.n202 163.367
R764 B.n400 B.n200 163.367
R765 B.n404 B.n200 163.367
R766 B.n404 B.n194 163.367
R767 B.n412 B.n194 163.367
R768 B.n412 B.n192 163.367
R769 B.n416 B.n192 163.367
R770 B.n416 B.n186 163.367
R771 B.n424 B.n186 163.367
R772 B.n424 B.n184 163.367
R773 B.n428 B.n184 163.367
R774 B.n428 B.n178 163.367
R775 B.n437 B.n178 163.367
R776 B.n437 B.n176 163.367
R777 B.n441 B.n176 163.367
R778 B.n441 B.n171 163.367
R779 B.n449 B.n171 163.367
R780 B.n449 B.n169 163.367
R781 B.n453 B.n169 163.367
R782 B.n453 B.n163 163.367
R783 B.n461 B.n163 163.367
R784 B.n461 B.n161 163.367
R785 B.n465 B.n161 163.367
R786 B.n465 B.n155 163.367
R787 B.n473 B.n155 163.367
R788 B.n473 B.n153 163.367
R789 B.n477 B.n153 163.367
R790 B.n477 B.n147 163.367
R791 B.n485 B.n147 163.367
R792 B.n485 B.n145 163.367
R793 B.n489 B.n145 163.367
R794 B.n489 B.n139 163.367
R795 B.n497 B.n139 163.367
R796 B.n497 B.n137 163.367
R797 B.n501 B.n137 163.367
R798 B.n501 B.n131 163.367
R799 B.n510 B.n131 163.367
R800 B.n510 B.n129 163.367
R801 B.n514 B.n129 163.367
R802 B.n514 B.n2 163.367
R803 B.n796 B.n2 163.367
R804 B.n796 B.n3 163.367
R805 B.n792 B.n3 163.367
R806 B.n792 B.n9 163.367
R807 B.n788 B.n9 163.367
R808 B.n788 B.n11 163.367
R809 B.n784 B.n11 163.367
R810 B.n784 B.n16 163.367
R811 B.n780 B.n16 163.367
R812 B.n780 B.n18 163.367
R813 B.n776 B.n18 163.367
R814 B.n776 B.n23 163.367
R815 B.n772 B.n23 163.367
R816 B.n772 B.n25 163.367
R817 B.n768 B.n25 163.367
R818 B.n768 B.n30 163.367
R819 B.n764 B.n30 163.367
R820 B.n764 B.n32 163.367
R821 B.n760 B.n32 163.367
R822 B.n760 B.n37 163.367
R823 B.n756 B.n37 163.367
R824 B.n756 B.n39 163.367
R825 B.n752 B.n39 163.367
R826 B.n752 B.n44 163.367
R827 B.n748 B.n44 163.367
R828 B.n748 B.n46 163.367
R829 B.n744 B.n46 163.367
R830 B.n744 B.n50 163.367
R831 B.n740 B.n50 163.367
R832 B.n740 B.n52 163.367
R833 B.n736 B.n52 163.367
R834 B.n736 B.n58 163.367
R835 B.n732 B.n58 163.367
R836 B.n732 B.n60 163.367
R837 B.n728 B.n60 163.367
R838 B.n728 B.n65 163.367
R839 B.n724 B.n65 163.367
R840 B.n724 B.n67 163.367
R841 B.n720 B.n67 163.367
R842 B.n720 B.n72 163.367
R843 B.n716 B.n72 163.367
R844 B.n716 B.n74 163.367
R845 B.n712 B.n74 163.367
R846 B.n712 B.n79 163.367
R847 B.n708 B.n79 163.367
R848 B.n708 B.n81 163.367
R849 B.n704 B.n81 163.367
R850 B.n704 B.n86 163.367
R851 B.n700 B.n86 163.367
R852 B.n700 B.n88 163.367
R853 B.n696 B.n88 163.367
R854 B.n364 B.n362 163.367
R855 B.n362 B.n361 163.367
R856 B.n358 B.n357 163.367
R857 B.n355 B.n228 163.367
R858 B.n351 B.n349 163.367
R859 B.n347 B.n230 163.367
R860 B.n343 B.n341 163.367
R861 B.n339 B.n232 163.367
R862 B.n335 B.n333 163.367
R863 B.n331 B.n234 163.367
R864 B.n327 B.n325 163.367
R865 B.n323 B.n236 163.367
R866 B.n318 B.n316 163.367
R867 B.n314 B.n240 163.367
R868 B.n310 B.n308 163.367
R869 B.n306 B.n242 163.367
R870 B.n302 B.n300 163.367
R871 B.n297 B.n296 163.367
R872 B.n294 B.n248 163.367
R873 B.n290 B.n288 163.367
R874 B.n286 B.n250 163.367
R875 B.n282 B.n280 163.367
R876 B.n278 B.n252 163.367
R877 B.n274 B.n272 163.367
R878 B.n270 B.n254 163.367
R879 B.n266 B.n264 163.367
R880 B.n262 B.n256 163.367
R881 B.n258 B.n222 163.367
R882 B.n370 B.n220 163.367
R883 B.n374 B.n220 163.367
R884 B.n374 B.n214 163.367
R885 B.n382 B.n214 163.367
R886 B.n382 B.n212 163.367
R887 B.n386 B.n212 163.367
R888 B.n386 B.n206 163.367
R889 B.n394 B.n206 163.367
R890 B.n394 B.n204 163.367
R891 B.n398 B.n204 163.367
R892 B.n398 B.n198 163.367
R893 B.n406 B.n198 163.367
R894 B.n406 B.n196 163.367
R895 B.n410 B.n196 163.367
R896 B.n410 B.n190 163.367
R897 B.n418 B.n190 163.367
R898 B.n418 B.n188 163.367
R899 B.n422 B.n188 163.367
R900 B.n422 B.n182 163.367
R901 B.n430 B.n182 163.367
R902 B.n430 B.n180 163.367
R903 B.n434 B.n180 163.367
R904 B.n434 B.n175 163.367
R905 B.n443 B.n175 163.367
R906 B.n443 B.n173 163.367
R907 B.n447 B.n173 163.367
R908 B.n447 B.n167 163.367
R909 B.n455 B.n167 163.367
R910 B.n455 B.n165 163.367
R911 B.n459 B.n165 163.367
R912 B.n459 B.n159 163.367
R913 B.n467 B.n159 163.367
R914 B.n467 B.n157 163.367
R915 B.n471 B.n157 163.367
R916 B.n471 B.n150 163.367
R917 B.n479 B.n150 163.367
R918 B.n479 B.n148 163.367
R919 B.n483 B.n148 163.367
R920 B.n483 B.n143 163.367
R921 B.n491 B.n143 163.367
R922 B.n491 B.n141 163.367
R923 B.n495 B.n141 163.367
R924 B.n495 B.n135 163.367
R925 B.n503 B.n135 163.367
R926 B.n503 B.n133 163.367
R927 B.n508 B.n133 163.367
R928 B.n508 B.n127 163.367
R929 B.n516 B.n127 163.367
R930 B.n517 B.n516 163.367
R931 B.n517 B.n5 163.367
R932 B.n6 B.n5 163.367
R933 B.n7 B.n6 163.367
R934 B.n522 B.n7 163.367
R935 B.n522 B.n12 163.367
R936 B.n13 B.n12 163.367
R937 B.n14 B.n13 163.367
R938 B.n527 B.n14 163.367
R939 B.n527 B.n19 163.367
R940 B.n20 B.n19 163.367
R941 B.n21 B.n20 163.367
R942 B.n532 B.n21 163.367
R943 B.n532 B.n26 163.367
R944 B.n27 B.n26 163.367
R945 B.n28 B.n27 163.367
R946 B.n537 B.n28 163.367
R947 B.n537 B.n33 163.367
R948 B.n34 B.n33 163.367
R949 B.n35 B.n34 163.367
R950 B.n542 B.n35 163.367
R951 B.n542 B.n40 163.367
R952 B.n41 B.n40 163.367
R953 B.n42 B.n41 163.367
R954 B.n547 B.n42 163.367
R955 B.n547 B.n47 163.367
R956 B.n48 B.n47 163.367
R957 B.n49 B.n48 163.367
R958 B.n552 B.n49 163.367
R959 B.n552 B.n54 163.367
R960 B.n55 B.n54 163.367
R961 B.n56 B.n55 163.367
R962 B.n557 B.n56 163.367
R963 B.n557 B.n61 163.367
R964 B.n62 B.n61 163.367
R965 B.n63 B.n62 163.367
R966 B.n562 B.n63 163.367
R967 B.n562 B.n68 163.367
R968 B.n69 B.n68 163.367
R969 B.n70 B.n69 163.367
R970 B.n567 B.n70 163.367
R971 B.n567 B.n75 163.367
R972 B.n76 B.n75 163.367
R973 B.n77 B.n76 163.367
R974 B.n572 B.n77 163.367
R975 B.n572 B.n82 163.367
R976 B.n83 B.n82 163.367
R977 B.n84 B.n83 163.367
R978 B.n577 B.n84 163.367
R979 B.n577 B.n89 163.367
R980 B.n90 B.n89 163.367
R981 B.n91 B.n90 163.367
R982 B.n692 B.n690 163.367
R983 B.n688 B.n95 163.367
R984 B.n684 B.n682 163.367
R985 B.n680 B.n97 163.367
R986 B.n676 B.n674 163.367
R987 B.n672 B.n99 163.367
R988 B.n668 B.n666 163.367
R989 B.n664 B.n101 163.367
R990 B.n660 B.n658 163.367
R991 B.n656 B.n103 163.367
R992 B.n652 B.n650 163.367
R993 B.n648 B.n105 163.367
R994 B.n644 B.n642 163.367
R995 B.n640 B.n110 163.367
R996 B.n636 B.n634 163.367
R997 B.n632 B.n112 163.367
R998 B.n627 B.n625 163.367
R999 B.n623 B.n116 163.367
R1000 B.n619 B.n617 163.367
R1001 B.n615 B.n118 163.367
R1002 B.n611 B.n609 163.367
R1003 B.n607 B.n120 163.367
R1004 B.n603 B.n601 163.367
R1005 B.n599 B.n122 163.367
R1006 B.n595 B.n593 163.367
R1007 B.n591 B.n124 163.367
R1008 B.n587 B.n585 163.367
R1009 B.n369 B.n223 131.298
R1010 B.n697 B.n92 131.298
R1011 B.n243 B.t20 120.838
R1012 B.n113 B.t22 120.838
R1013 B.n237 B.t17 120.832
R1014 B.n106 B.t12 120.832
R1015 B.n244 B.t19 74.6805
R1016 B.n114 B.t23 74.6805
R1017 B.n238 B.t16 74.6747
R1018 B.n107 B.t13 74.6747
R1019 B.n363 B.n224 71.676
R1020 B.n361 B.n226 71.676
R1021 B.n357 B.n356 71.676
R1022 B.n350 B.n228 71.676
R1023 B.n349 B.n348 71.676
R1024 B.n342 B.n230 71.676
R1025 B.n341 B.n340 71.676
R1026 B.n334 B.n232 71.676
R1027 B.n333 B.n332 71.676
R1028 B.n326 B.n234 71.676
R1029 B.n325 B.n324 71.676
R1030 B.n317 B.n236 71.676
R1031 B.n316 B.n315 71.676
R1032 B.n309 B.n240 71.676
R1033 B.n308 B.n307 71.676
R1034 B.n301 B.n242 71.676
R1035 B.n300 B.n246 71.676
R1036 B.n296 B.n295 71.676
R1037 B.n289 B.n248 71.676
R1038 B.n288 B.n287 71.676
R1039 B.n281 B.n250 71.676
R1040 B.n280 B.n279 71.676
R1041 B.n273 B.n252 71.676
R1042 B.n272 B.n271 71.676
R1043 B.n265 B.n254 71.676
R1044 B.n264 B.n263 71.676
R1045 B.n257 B.n256 71.676
R1046 B.n691 B.n93 71.676
R1047 B.n690 B.n689 71.676
R1048 B.n683 B.n95 71.676
R1049 B.n682 B.n681 71.676
R1050 B.n675 B.n97 71.676
R1051 B.n674 B.n673 71.676
R1052 B.n667 B.n99 71.676
R1053 B.n666 B.n665 71.676
R1054 B.n659 B.n101 71.676
R1055 B.n658 B.n657 71.676
R1056 B.n651 B.n103 71.676
R1057 B.n650 B.n649 71.676
R1058 B.n643 B.n105 71.676
R1059 B.n642 B.n641 71.676
R1060 B.n635 B.n110 71.676
R1061 B.n634 B.n633 71.676
R1062 B.n626 B.n112 71.676
R1063 B.n625 B.n624 71.676
R1064 B.n618 B.n116 71.676
R1065 B.n617 B.n616 71.676
R1066 B.n610 B.n118 71.676
R1067 B.n609 B.n608 71.676
R1068 B.n602 B.n120 71.676
R1069 B.n601 B.n600 71.676
R1070 B.n594 B.n122 71.676
R1071 B.n593 B.n592 71.676
R1072 B.n586 B.n124 71.676
R1073 B.n585 B.n584 71.676
R1074 B.n584 B.n583 71.676
R1075 B.n587 B.n586 71.676
R1076 B.n592 B.n591 71.676
R1077 B.n595 B.n594 71.676
R1078 B.n600 B.n599 71.676
R1079 B.n603 B.n602 71.676
R1080 B.n608 B.n607 71.676
R1081 B.n611 B.n610 71.676
R1082 B.n616 B.n615 71.676
R1083 B.n619 B.n618 71.676
R1084 B.n624 B.n623 71.676
R1085 B.n627 B.n626 71.676
R1086 B.n633 B.n632 71.676
R1087 B.n636 B.n635 71.676
R1088 B.n641 B.n640 71.676
R1089 B.n644 B.n643 71.676
R1090 B.n649 B.n648 71.676
R1091 B.n652 B.n651 71.676
R1092 B.n657 B.n656 71.676
R1093 B.n660 B.n659 71.676
R1094 B.n665 B.n664 71.676
R1095 B.n668 B.n667 71.676
R1096 B.n673 B.n672 71.676
R1097 B.n676 B.n675 71.676
R1098 B.n681 B.n680 71.676
R1099 B.n684 B.n683 71.676
R1100 B.n689 B.n688 71.676
R1101 B.n692 B.n691 71.676
R1102 B.n364 B.n363 71.676
R1103 B.n358 B.n226 71.676
R1104 B.n356 B.n355 71.676
R1105 B.n351 B.n350 71.676
R1106 B.n348 B.n347 71.676
R1107 B.n343 B.n342 71.676
R1108 B.n340 B.n339 71.676
R1109 B.n335 B.n334 71.676
R1110 B.n332 B.n331 71.676
R1111 B.n327 B.n326 71.676
R1112 B.n324 B.n323 71.676
R1113 B.n318 B.n317 71.676
R1114 B.n315 B.n314 71.676
R1115 B.n310 B.n309 71.676
R1116 B.n307 B.n306 71.676
R1117 B.n302 B.n301 71.676
R1118 B.n297 B.n246 71.676
R1119 B.n295 B.n294 71.676
R1120 B.n290 B.n289 71.676
R1121 B.n287 B.n286 71.676
R1122 B.n282 B.n281 71.676
R1123 B.n279 B.n278 71.676
R1124 B.n274 B.n273 71.676
R1125 B.n271 B.n270 71.676
R1126 B.n266 B.n265 71.676
R1127 B.n263 B.n262 71.676
R1128 B.n258 B.n257 71.676
R1129 B.n369 B.n219 68.1554
R1130 B.n375 B.n219 68.1554
R1131 B.n375 B.n215 68.1554
R1132 B.n381 B.n215 68.1554
R1133 B.n381 B.n211 68.1554
R1134 B.n387 B.n211 68.1554
R1135 B.n393 B.n207 68.1554
R1136 B.n393 B.n203 68.1554
R1137 B.n399 B.n203 68.1554
R1138 B.n399 B.n199 68.1554
R1139 B.n405 B.n199 68.1554
R1140 B.n405 B.n195 68.1554
R1141 B.n411 B.n195 68.1554
R1142 B.n411 B.n191 68.1554
R1143 B.n417 B.n191 68.1554
R1144 B.n423 B.n187 68.1554
R1145 B.n423 B.n183 68.1554
R1146 B.n429 B.n183 68.1554
R1147 B.n429 B.n179 68.1554
R1148 B.n436 B.n179 68.1554
R1149 B.n436 B.n435 68.1554
R1150 B.n442 B.n172 68.1554
R1151 B.n448 B.n172 68.1554
R1152 B.n448 B.n168 68.1554
R1153 B.n454 B.n168 68.1554
R1154 B.n454 B.n164 68.1554
R1155 B.n460 B.n164 68.1554
R1156 B.n466 B.n160 68.1554
R1157 B.n466 B.n156 68.1554
R1158 B.n472 B.n156 68.1554
R1159 B.n472 B.n151 68.1554
R1160 B.n478 B.n151 68.1554
R1161 B.n478 B.n152 68.1554
R1162 B.n484 B.n144 68.1554
R1163 B.n490 B.n144 68.1554
R1164 B.n490 B.n140 68.1554
R1165 B.n496 B.n140 68.1554
R1166 B.n496 B.n136 68.1554
R1167 B.n502 B.n136 68.1554
R1168 B.n509 B.n132 68.1554
R1169 B.n509 B.n128 68.1554
R1170 B.n515 B.n128 68.1554
R1171 B.n515 B.n4 68.1554
R1172 B.n795 B.n4 68.1554
R1173 B.n795 B.n794 68.1554
R1174 B.n794 B.n793 68.1554
R1175 B.n793 B.n8 68.1554
R1176 B.n787 B.n8 68.1554
R1177 B.n787 B.n786 68.1554
R1178 B.n785 B.n15 68.1554
R1179 B.n779 B.n15 68.1554
R1180 B.n779 B.n778 68.1554
R1181 B.n778 B.n777 68.1554
R1182 B.n777 B.n22 68.1554
R1183 B.n771 B.n22 68.1554
R1184 B.n770 B.n769 68.1554
R1185 B.n769 B.n29 68.1554
R1186 B.n763 B.n29 68.1554
R1187 B.n763 B.n762 68.1554
R1188 B.n762 B.n761 68.1554
R1189 B.n761 B.n36 68.1554
R1190 B.n755 B.n754 68.1554
R1191 B.n754 B.n753 68.1554
R1192 B.n753 B.n43 68.1554
R1193 B.n747 B.n43 68.1554
R1194 B.n747 B.n746 68.1554
R1195 B.n746 B.n745 68.1554
R1196 B.n739 B.n53 68.1554
R1197 B.n739 B.n738 68.1554
R1198 B.n738 B.n737 68.1554
R1199 B.n737 B.n57 68.1554
R1200 B.n731 B.n57 68.1554
R1201 B.n731 B.n730 68.1554
R1202 B.n729 B.n64 68.1554
R1203 B.n723 B.n64 68.1554
R1204 B.n723 B.n722 68.1554
R1205 B.n722 B.n721 68.1554
R1206 B.n721 B.n71 68.1554
R1207 B.n715 B.n71 68.1554
R1208 B.n715 B.n714 68.1554
R1209 B.n714 B.n713 68.1554
R1210 B.n713 B.n78 68.1554
R1211 B.n707 B.n706 68.1554
R1212 B.n706 B.n705 68.1554
R1213 B.n705 B.n85 68.1554
R1214 B.n699 B.n85 68.1554
R1215 B.n699 B.n698 68.1554
R1216 B.n698 B.n697 68.1554
R1217 B.n417 B.t0 61.1395
R1218 B.n435 B.t9 61.1395
R1219 B.n460 B.t2 61.1395
R1220 B.n152 B.t7 61.1395
R1221 B.n502 B.t6 61.1395
R1222 B.t8 B.n785 61.1395
R1223 B.t4 B.n770 61.1395
R1224 B.n755 B.t3 61.1395
R1225 B.n53 B.t5 61.1395
R1226 B.t1 B.n729 61.1395
R1227 B.n245 B.n244 59.5399
R1228 B.n321 B.n238 59.5399
R1229 B.n108 B.n107 59.5399
R1230 B.n629 B.n114 59.5399
R1231 B.n387 B.t15 47.1076
R1232 B.n707 B.t11 47.1076
R1233 B.n244 B.n243 46.1581
R1234 B.n238 B.n237 46.1581
R1235 B.n107 B.n106 46.1581
R1236 B.n114 B.n113 46.1581
R1237 B.n695 B.n694 32.3127
R1238 B.n582 B.n581 32.3127
R1239 B.n371 B.n221 32.3127
R1240 B.n367 B.n366 32.3127
R1241 B.t15 B.n207 21.0483
R1242 B.t11 B.n78 21.0483
R1243 B B.n797 18.0485
R1244 B.n694 B.n693 10.6151
R1245 B.n693 B.n94 10.6151
R1246 B.n687 B.n94 10.6151
R1247 B.n687 B.n686 10.6151
R1248 B.n686 B.n685 10.6151
R1249 B.n685 B.n96 10.6151
R1250 B.n679 B.n96 10.6151
R1251 B.n679 B.n678 10.6151
R1252 B.n678 B.n677 10.6151
R1253 B.n677 B.n98 10.6151
R1254 B.n671 B.n98 10.6151
R1255 B.n671 B.n670 10.6151
R1256 B.n670 B.n669 10.6151
R1257 B.n669 B.n100 10.6151
R1258 B.n663 B.n100 10.6151
R1259 B.n663 B.n662 10.6151
R1260 B.n662 B.n661 10.6151
R1261 B.n661 B.n102 10.6151
R1262 B.n655 B.n102 10.6151
R1263 B.n655 B.n654 10.6151
R1264 B.n654 B.n653 10.6151
R1265 B.n653 B.n104 10.6151
R1266 B.n647 B.n646 10.6151
R1267 B.n646 B.n645 10.6151
R1268 B.n645 B.n109 10.6151
R1269 B.n639 B.n109 10.6151
R1270 B.n639 B.n638 10.6151
R1271 B.n638 B.n637 10.6151
R1272 B.n637 B.n111 10.6151
R1273 B.n631 B.n111 10.6151
R1274 B.n631 B.n630 10.6151
R1275 B.n628 B.n115 10.6151
R1276 B.n622 B.n115 10.6151
R1277 B.n622 B.n621 10.6151
R1278 B.n621 B.n620 10.6151
R1279 B.n620 B.n117 10.6151
R1280 B.n614 B.n117 10.6151
R1281 B.n614 B.n613 10.6151
R1282 B.n613 B.n612 10.6151
R1283 B.n612 B.n119 10.6151
R1284 B.n606 B.n119 10.6151
R1285 B.n606 B.n605 10.6151
R1286 B.n605 B.n604 10.6151
R1287 B.n604 B.n121 10.6151
R1288 B.n598 B.n121 10.6151
R1289 B.n598 B.n597 10.6151
R1290 B.n597 B.n596 10.6151
R1291 B.n596 B.n123 10.6151
R1292 B.n590 B.n123 10.6151
R1293 B.n590 B.n589 10.6151
R1294 B.n589 B.n588 10.6151
R1295 B.n588 B.n125 10.6151
R1296 B.n582 B.n125 10.6151
R1297 B.n372 B.n371 10.6151
R1298 B.n373 B.n372 10.6151
R1299 B.n373 B.n213 10.6151
R1300 B.n383 B.n213 10.6151
R1301 B.n384 B.n383 10.6151
R1302 B.n385 B.n384 10.6151
R1303 B.n385 B.n205 10.6151
R1304 B.n395 B.n205 10.6151
R1305 B.n396 B.n395 10.6151
R1306 B.n397 B.n396 10.6151
R1307 B.n397 B.n197 10.6151
R1308 B.n407 B.n197 10.6151
R1309 B.n408 B.n407 10.6151
R1310 B.n409 B.n408 10.6151
R1311 B.n409 B.n189 10.6151
R1312 B.n419 B.n189 10.6151
R1313 B.n420 B.n419 10.6151
R1314 B.n421 B.n420 10.6151
R1315 B.n421 B.n181 10.6151
R1316 B.n431 B.n181 10.6151
R1317 B.n432 B.n431 10.6151
R1318 B.n433 B.n432 10.6151
R1319 B.n433 B.n174 10.6151
R1320 B.n444 B.n174 10.6151
R1321 B.n445 B.n444 10.6151
R1322 B.n446 B.n445 10.6151
R1323 B.n446 B.n166 10.6151
R1324 B.n456 B.n166 10.6151
R1325 B.n457 B.n456 10.6151
R1326 B.n458 B.n457 10.6151
R1327 B.n458 B.n158 10.6151
R1328 B.n468 B.n158 10.6151
R1329 B.n469 B.n468 10.6151
R1330 B.n470 B.n469 10.6151
R1331 B.n470 B.n149 10.6151
R1332 B.n480 B.n149 10.6151
R1333 B.n481 B.n480 10.6151
R1334 B.n482 B.n481 10.6151
R1335 B.n482 B.n142 10.6151
R1336 B.n492 B.n142 10.6151
R1337 B.n493 B.n492 10.6151
R1338 B.n494 B.n493 10.6151
R1339 B.n494 B.n134 10.6151
R1340 B.n504 B.n134 10.6151
R1341 B.n505 B.n504 10.6151
R1342 B.n507 B.n505 10.6151
R1343 B.n507 B.n506 10.6151
R1344 B.n506 B.n126 10.6151
R1345 B.n518 B.n126 10.6151
R1346 B.n519 B.n518 10.6151
R1347 B.n520 B.n519 10.6151
R1348 B.n521 B.n520 10.6151
R1349 B.n523 B.n521 10.6151
R1350 B.n524 B.n523 10.6151
R1351 B.n525 B.n524 10.6151
R1352 B.n526 B.n525 10.6151
R1353 B.n528 B.n526 10.6151
R1354 B.n529 B.n528 10.6151
R1355 B.n530 B.n529 10.6151
R1356 B.n531 B.n530 10.6151
R1357 B.n533 B.n531 10.6151
R1358 B.n534 B.n533 10.6151
R1359 B.n535 B.n534 10.6151
R1360 B.n536 B.n535 10.6151
R1361 B.n538 B.n536 10.6151
R1362 B.n539 B.n538 10.6151
R1363 B.n540 B.n539 10.6151
R1364 B.n541 B.n540 10.6151
R1365 B.n543 B.n541 10.6151
R1366 B.n544 B.n543 10.6151
R1367 B.n545 B.n544 10.6151
R1368 B.n546 B.n545 10.6151
R1369 B.n548 B.n546 10.6151
R1370 B.n549 B.n548 10.6151
R1371 B.n550 B.n549 10.6151
R1372 B.n551 B.n550 10.6151
R1373 B.n553 B.n551 10.6151
R1374 B.n554 B.n553 10.6151
R1375 B.n555 B.n554 10.6151
R1376 B.n556 B.n555 10.6151
R1377 B.n558 B.n556 10.6151
R1378 B.n559 B.n558 10.6151
R1379 B.n560 B.n559 10.6151
R1380 B.n561 B.n560 10.6151
R1381 B.n563 B.n561 10.6151
R1382 B.n564 B.n563 10.6151
R1383 B.n565 B.n564 10.6151
R1384 B.n566 B.n565 10.6151
R1385 B.n568 B.n566 10.6151
R1386 B.n569 B.n568 10.6151
R1387 B.n570 B.n569 10.6151
R1388 B.n571 B.n570 10.6151
R1389 B.n573 B.n571 10.6151
R1390 B.n574 B.n573 10.6151
R1391 B.n575 B.n574 10.6151
R1392 B.n576 B.n575 10.6151
R1393 B.n578 B.n576 10.6151
R1394 B.n579 B.n578 10.6151
R1395 B.n580 B.n579 10.6151
R1396 B.n581 B.n580 10.6151
R1397 B.n366 B.n365 10.6151
R1398 B.n365 B.n225 10.6151
R1399 B.n360 B.n225 10.6151
R1400 B.n360 B.n359 10.6151
R1401 B.n359 B.n227 10.6151
R1402 B.n354 B.n227 10.6151
R1403 B.n354 B.n353 10.6151
R1404 B.n353 B.n352 10.6151
R1405 B.n352 B.n229 10.6151
R1406 B.n346 B.n229 10.6151
R1407 B.n346 B.n345 10.6151
R1408 B.n345 B.n344 10.6151
R1409 B.n344 B.n231 10.6151
R1410 B.n338 B.n231 10.6151
R1411 B.n338 B.n337 10.6151
R1412 B.n337 B.n336 10.6151
R1413 B.n336 B.n233 10.6151
R1414 B.n330 B.n233 10.6151
R1415 B.n330 B.n329 10.6151
R1416 B.n329 B.n328 10.6151
R1417 B.n328 B.n235 10.6151
R1418 B.n322 B.n235 10.6151
R1419 B.n320 B.n319 10.6151
R1420 B.n319 B.n239 10.6151
R1421 B.n313 B.n239 10.6151
R1422 B.n313 B.n312 10.6151
R1423 B.n312 B.n311 10.6151
R1424 B.n311 B.n241 10.6151
R1425 B.n305 B.n241 10.6151
R1426 B.n305 B.n304 10.6151
R1427 B.n304 B.n303 10.6151
R1428 B.n299 B.n298 10.6151
R1429 B.n298 B.n247 10.6151
R1430 B.n293 B.n247 10.6151
R1431 B.n293 B.n292 10.6151
R1432 B.n292 B.n291 10.6151
R1433 B.n291 B.n249 10.6151
R1434 B.n285 B.n249 10.6151
R1435 B.n285 B.n284 10.6151
R1436 B.n284 B.n283 10.6151
R1437 B.n283 B.n251 10.6151
R1438 B.n277 B.n251 10.6151
R1439 B.n277 B.n276 10.6151
R1440 B.n276 B.n275 10.6151
R1441 B.n275 B.n253 10.6151
R1442 B.n269 B.n253 10.6151
R1443 B.n269 B.n268 10.6151
R1444 B.n268 B.n267 10.6151
R1445 B.n267 B.n255 10.6151
R1446 B.n261 B.n255 10.6151
R1447 B.n261 B.n260 10.6151
R1448 B.n260 B.n259 10.6151
R1449 B.n259 B.n221 10.6151
R1450 B.n367 B.n217 10.6151
R1451 B.n377 B.n217 10.6151
R1452 B.n378 B.n377 10.6151
R1453 B.n379 B.n378 10.6151
R1454 B.n379 B.n209 10.6151
R1455 B.n389 B.n209 10.6151
R1456 B.n390 B.n389 10.6151
R1457 B.n391 B.n390 10.6151
R1458 B.n391 B.n201 10.6151
R1459 B.n401 B.n201 10.6151
R1460 B.n402 B.n401 10.6151
R1461 B.n403 B.n402 10.6151
R1462 B.n403 B.n193 10.6151
R1463 B.n413 B.n193 10.6151
R1464 B.n414 B.n413 10.6151
R1465 B.n415 B.n414 10.6151
R1466 B.n415 B.n185 10.6151
R1467 B.n425 B.n185 10.6151
R1468 B.n426 B.n425 10.6151
R1469 B.n427 B.n426 10.6151
R1470 B.n427 B.n177 10.6151
R1471 B.n438 B.n177 10.6151
R1472 B.n439 B.n438 10.6151
R1473 B.n440 B.n439 10.6151
R1474 B.n440 B.n170 10.6151
R1475 B.n450 B.n170 10.6151
R1476 B.n451 B.n450 10.6151
R1477 B.n452 B.n451 10.6151
R1478 B.n452 B.n162 10.6151
R1479 B.n462 B.n162 10.6151
R1480 B.n463 B.n462 10.6151
R1481 B.n464 B.n463 10.6151
R1482 B.n464 B.n154 10.6151
R1483 B.n474 B.n154 10.6151
R1484 B.n475 B.n474 10.6151
R1485 B.n476 B.n475 10.6151
R1486 B.n476 B.n146 10.6151
R1487 B.n486 B.n146 10.6151
R1488 B.n487 B.n486 10.6151
R1489 B.n488 B.n487 10.6151
R1490 B.n488 B.n138 10.6151
R1491 B.n498 B.n138 10.6151
R1492 B.n499 B.n498 10.6151
R1493 B.n500 B.n499 10.6151
R1494 B.n500 B.n130 10.6151
R1495 B.n511 B.n130 10.6151
R1496 B.n512 B.n511 10.6151
R1497 B.n513 B.n512 10.6151
R1498 B.n513 B.n0 10.6151
R1499 B.n791 B.n1 10.6151
R1500 B.n791 B.n790 10.6151
R1501 B.n790 B.n789 10.6151
R1502 B.n789 B.n10 10.6151
R1503 B.n783 B.n10 10.6151
R1504 B.n783 B.n782 10.6151
R1505 B.n782 B.n781 10.6151
R1506 B.n781 B.n17 10.6151
R1507 B.n775 B.n17 10.6151
R1508 B.n775 B.n774 10.6151
R1509 B.n774 B.n773 10.6151
R1510 B.n773 B.n24 10.6151
R1511 B.n767 B.n24 10.6151
R1512 B.n767 B.n766 10.6151
R1513 B.n766 B.n765 10.6151
R1514 B.n765 B.n31 10.6151
R1515 B.n759 B.n31 10.6151
R1516 B.n759 B.n758 10.6151
R1517 B.n758 B.n757 10.6151
R1518 B.n757 B.n38 10.6151
R1519 B.n751 B.n38 10.6151
R1520 B.n751 B.n750 10.6151
R1521 B.n750 B.n749 10.6151
R1522 B.n749 B.n45 10.6151
R1523 B.n743 B.n45 10.6151
R1524 B.n743 B.n742 10.6151
R1525 B.n742 B.n741 10.6151
R1526 B.n741 B.n51 10.6151
R1527 B.n735 B.n51 10.6151
R1528 B.n735 B.n734 10.6151
R1529 B.n734 B.n733 10.6151
R1530 B.n733 B.n59 10.6151
R1531 B.n727 B.n59 10.6151
R1532 B.n727 B.n726 10.6151
R1533 B.n726 B.n725 10.6151
R1534 B.n725 B.n66 10.6151
R1535 B.n719 B.n66 10.6151
R1536 B.n719 B.n718 10.6151
R1537 B.n718 B.n717 10.6151
R1538 B.n717 B.n73 10.6151
R1539 B.n711 B.n73 10.6151
R1540 B.n711 B.n710 10.6151
R1541 B.n710 B.n709 10.6151
R1542 B.n709 B.n80 10.6151
R1543 B.n703 B.n80 10.6151
R1544 B.n703 B.n702 10.6151
R1545 B.n702 B.n701 10.6151
R1546 B.n701 B.n87 10.6151
R1547 B.n695 B.n87 10.6151
R1548 B.n108 B.n104 9.36635
R1549 B.n629 B.n628 9.36635
R1550 B.n322 B.n321 9.36635
R1551 B.n299 B.n245 9.36635
R1552 B.t0 B.n187 7.01645
R1553 B.n442 B.t9 7.01645
R1554 B.t2 B.n160 7.01645
R1555 B.n484 B.t7 7.01645
R1556 B.t6 B.n132 7.01645
R1557 B.n786 B.t8 7.01645
R1558 B.n771 B.t4 7.01645
R1559 B.t3 B.n36 7.01645
R1560 B.n745 B.t5 7.01645
R1561 B.n730 B.t1 7.01645
R1562 B.n797 B.n0 2.81026
R1563 B.n797 B.n1 2.81026
R1564 B.n647 B.n108 1.24928
R1565 B.n630 B.n629 1.24928
R1566 B.n321 B.n320 1.24928
R1567 B.n303 B.n245 1.24928
R1568 VP.n48 VP.n47 185.4
R1569 VP.n82 VP.n81 185.4
R1570 VP.n46 VP.n45 185.4
R1571 VP.n22 VP.n21 161.3
R1572 VP.n23 VP.n18 161.3
R1573 VP.n25 VP.n24 161.3
R1574 VP.n26 VP.n17 161.3
R1575 VP.n28 VP.n27 161.3
R1576 VP.n30 VP.n29 161.3
R1577 VP.n31 VP.n15 161.3
R1578 VP.n33 VP.n32 161.3
R1579 VP.n34 VP.n14 161.3
R1580 VP.n36 VP.n35 161.3
R1581 VP.n38 VP.n13 161.3
R1582 VP.n40 VP.n39 161.3
R1583 VP.n41 VP.n12 161.3
R1584 VP.n43 VP.n42 161.3
R1585 VP.n44 VP.n11 161.3
R1586 VP.n80 VP.n0 161.3
R1587 VP.n79 VP.n78 161.3
R1588 VP.n77 VP.n1 161.3
R1589 VP.n76 VP.n75 161.3
R1590 VP.n74 VP.n2 161.3
R1591 VP.n72 VP.n71 161.3
R1592 VP.n70 VP.n3 161.3
R1593 VP.n69 VP.n68 161.3
R1594 VP.n67 VP.n4 161.3
R1595 VP.n66 VP.n65 161.3
R1596 VP.n64 VP.n63 161.3
R1597 VP.n62 VP.n6 161.3
R1598 VP.n61 VP.n60 161.3
R1599 VP.n59 VP.n7 161.3
R1600 VP.n58 VP.n57 161.3
R1601 VP.n55 VP.n8 161.3
R1602 VP.n54 VP.n53 161.3
R1603 VP.n52 VP.n9 161.3
R1604 VP.n51 VP.n50 161.3
R1605 VP.n49 VP.n10 161.3
R1606 VP.n19 VP.t0 98.5
R1607 VP.n48 VP.t1 67.0103
R1608 VP.n56 VP.t8 67.0103
R1609 VP.n5 VP.t4 67.0103
R1610 VP.n73 VP.t9 67.0103
R1611 VP.n81 VP.t3 67.0103
R1612 VP.n45 VP.t7 67.0103
R1613 VP.n37 VP.t6 67.0103
R1614 VP.n16 VP.t5 67.0103
R1615 VP.n20 VP.t2 67.0103
R1616 VP.n20 VP.n19 64.2931
R1617 VP.n54 VP.n9 56.5617
R1618 VP.n75 VP.n1 56.5617
R1619 VP.n39 VP.n12 56.5617
R1620 VP.n62 VP.n61 46.3896
R1621 VP.n68 VP.n67 46.3896
R1622 VP.n32 VP.n31 46.3896
R1623 VP.n26 VP.n25 46.3896
R1624 VP.n47 VP.n46 45.2656
R1625 VP.n61 VP.n7 34.7644
R1626 VP.n68 VP.n3 34.7644
R1627 VP.n32 VP.n14 34.7644
R1628 VP.n25 VP.n18 34.7644
R1629 VP.n50 VP.n49 24.5923
R1630 VP.n50 VP.n9 24.5923
R1631 VP.n55 VP.n54 24.5923
R1632 VP.n57 VP.n7 24.5923
R1633 VP.n63 VP.n62 24.5923
R1634 VP.n67 VP.n66 24.5923
R1635 VP.n72 VP.n3 24.5923
R1636 VP.n75 VP.n74 24.5923
R1637 VP.n79 VP.n1 24.5923
R1638 VP.n80 VP.n79 24.5923
R1639 VP.n43 VP.n12 24.5923
R1640 VP.n44 VP.n43 24.5923
R1641 VP.n36 VP.n14 24.5923
R1642 VP.n39 VP.n38 24.5923
R1643 VP.n27 VP.n26 24.5923
R1644 VP.n31 VP.n30 24.5923
R1645 VP.n21 VP.n18 24.5923
R1646 VP.n56 VP.n55 18.1985
R1647 VP.n74 VP.n73 18.1985
R1648 VP.n38 VP.n37 18.1985
R1649 VP.n22 VP.n19 12.6154
R1650 VP.n63 VP.n5 12.2964
R1651 VP.n66 VP.n5 12.2964
R1652 VP.n27 VP.n16 12.2964
R1653 VP.n30 VP.n16 12.2964
R1654 VP.n57 VP.n56 6.39438
R1655 VP.n73 VP.n72 6.39438
R1656 VP.n37 VP.n36 6.39438
R1657 VP.n21 VP.n20 6.39438
R1658 VP.n49 VP.n48 0.492337
R1659 VP.n81 VP.n80 0.492337
R1660 VP.n45 VP.n44 0.492337
R1661 VP.n23 VP.n22 0.189894
R1662 VP.n24 VP.n23 0.189894
R1663 VP.n24 VP.n17 0.189894
R1664 VP.n28 VP.n17 0.189894
R1665 VP.n29 VP.n28 0.189894
R1666 VP.n29 VP.n15 0.189894
R1667 VP.n33 VP.n15 0.189894
R1668 VP.n34 VP.n33 0.189894
R1669 VP.n35 VP.n34 0.189894
R1670 VP.n35 VP.n13 0.189894
R1671 VP.n40 VP.n13 0.189894
R1672 VP.n41 VP.n40 0.189894
R1673 VP.n42 VP.n41 0.189894
R1674 VP.n42 VP.n11 0.189894
R1675 VP.n46 VP.n11 0.189894
R1676 VP.n47 VP.n10 0.189894
R1677 VP.n51 VP.n10 0.189894
R1678 VP.n52 VP.n51 0.189894
R1679 VP.n53 VP.n52 0.189894
R1680 VP.n53 VP.n8 0.189894
R1681 VP.n58 VP.n8 0.189894
R1682 VP.n59 VP.n58 0.189894
R1683 VP.n60 VP.n59 0.189894
R1684 VP.n60 VP.n6 0.189894
R1685 VP.n64 VP.n6 0.189894
R1686 VP.n65 VP.n64 0.189894
R1687 VP.n65 VP.n4 0.189894
R1688 VP.n69 VP.n4 0.189894
R1689 VP.n70 VP.n69 0.189894
R1690 VP.n71 VP.n70 0.189894
R1691 VP.n71 VP.n2 0.189894
R1692 VP.n76 VP.n2 0.189894
R1693 VP.n77 VP.n76 0.189894
R1694 VP.n78 VP.n77 0.189894
R1695 VP.n78 VP.n0 0.189894
R1696 VP.n82 VP.n0 0.189894
R1697 VP VP.n82 0.0516364
R1698 VDD1.n1 VDD1.t9 74.5591
R1699 VDD1.n3 VDD1.t8 74.5589
R1700 VDD1.n5 VDD1.n4 70.5169
R1701 VDD1.n1 VDD1.n0 69.0337
R1702 VDD1.n7 VDD1.n6 69.0335
R1703 VDD1.n3 VDD1.n2 69.0334
R1704 VDD1.n7 VDD1.n5 39.9837
R1705 VDD1.n6 VDD1.t3 3.47418
R1706 VDD1.n6 VDD1.t2 3.47418
R1707 VDD1.n0 VDD1.t7 3.47418
R1708 VDD1.n0 VDD1.t4 3.47418
R1709 VDD1.n4 VDD1.t0 3.47418
R1710 VDD1.n4 VDD1.t6 3.47418
R1711 VDD1.n2 VDD1.t1 3.47418
R1712 VDD1.n2 VDD1.t5 3.47418
R1713 VDD1 VDD1.n7 1.4811
R1714 VDD1 VDD1.n1 0.571621
R1715 VDD1.n5 VDD1.n3 0.458085
C0 VN VP 6.41251f
C1 VTAIL VP 5.9336f
C2 VTAIL VN 5.91939f
C3 VDD1 VP 5.42828f
C4 VDD2 VP 0.513142f
C5 VDD1 VN 0.15239f
C6 VDD2 VN 5.07012f
C7 VDD1 VTAIL 7.14208f
C8 VDD2 VTAIL 7.19046f
C9 VDD2 VDD1 1.81535f
C10 VDD2 B 5.42448f
C11 VDD1 B 5.408313f
C12 VTAIL B 4.938972f
C13 VN B 14.83876f
C14 VP B 13.381405f
C15 VDD1.t9 B 1.0971f
C16 VDD1.t7 B 0.103086f
C17 VDD1.t4 B 0.103086f
C18 VDD1.n0 B 0.854568f
C19 VDD1.n1 B 0.761651f
C20 VDD1.t8 B 1.0971f
C21 VDD1.t1 B 0.103086f
C22 VDD1.t5 B 0.103086f
C23 VDD1.n2 B 0.854565f
C24 VDD1.n3 B 0.754444f
C25 VDD1.t0 B 0.103086f
C26 VDD1.t6 B 0.103086f
C27 VDD1.n4 B 0.864133f
C28 VDD1.n5 B 2.14146f
C29 VDD1.t3 B 0.103086f
C30 VDD1.t2 B 0.103086f
C31 VDD1.n6 B 0.854564f
C32 VDD1.n7 B 2.24443f
C33 VP.n0 B 0.027937f
C34 VP.t3 B 0.861341f
C35 VP.n1 B 0.0352f
C36 VP.n2 B 0.027937f
C37 VP.t9 B 0.861341f
C38 VP.n3 B 0.056146f
C39 VP.n4 B 0.027937f
C40 VP.t4 B 0.861341f
C41 VP.n5 B 0.330522f
C42 VP.n6 B 0.027937f
C43 VP.n7 B 0.056146f
C44 VP.n8 B 0.027937f
C45 VP.t8 B 0.861341f
C46 VP.n9 B 0.0352f
C47 VP.n10 B 0.027937f
C48 VP.t1 B 0.861341f
C49 VP.n11 B 0.027937f
C50 VP.t7 B 0.861341f
C51 VP.n12 B 0.0352f
C52 VP.n13 B 0.027937f
C53 VP.t6 B 0.861341f
C54 VP.n14 B 0.056146f
C55 VP.n15 B 0.027937f
C56 VP.t5 B 0.861341f
C57 VP.n16 B 0.330522f
C58 VP.n17 B 0.027937f
C59 VP.n18 B 0.056146f
C60 VP.t0 B 1.01298f
C61 VP.n19 B 0.397353f
C62 VP.t2 B 0.861341f
C63 VP.n20 B 0.392639f
C64 VP.n21 B 0.03288f
C65 VP.n22 B 0.210162f
C66 VP.n23 B 0.027937f
C67 VP.n24 B 0.027937f
C68 VP.n25 B 0.023872f
C69 VP.n26 B 0.053008f
C70 VP.n27 B 0.039019f
C71 VP.n28 B 0.027937f
C72 VP.n29 B 0.027937f
C73 VP.n30 B 0.039019f
C74 VP.n31 B 0.053008f
C75 VP.n32 B 0.023872f
C76 VP.n33 B 0.027937f
C77 VP.n34 B 0.027937f
C78 VP.n35 B 0.027937f
C79 VP.n36 B 0.03288f
C80 VP.n37 B 0.330522f
C81 VP.n38 B 0.045157f
C82 VP.n39 B 0.046021f
C83 VP.n40 B 0.027937f
C84 VP.n41 B 0.027937f
C85 VP.n42 B 0.027937f
C86 VP.n43 B 0.051806f
C87 VP.n44 B 0.026742f
C88 VP.n45 B 0.400515f
C89 VP.n46 B 1.31293f
C90 VP.n47 B 1.33518f
C91 VP.n48 B 0.400515f
C92 VP.n49 B 0.026742f
C93 VP.n50 B 0.051806f
C94 VP.n51 B 0.027937f
C95 VP.n52 B 0.027937f
C96 VP.n53 B 0.027937f
C97 VP.n54 B 0.046021f
C98 VP.n55 B 0.045157f
C99 VP.n56 B 0.330522f
C100 VP.n57 B 0.03288f
C101 VP.n58 B 0.027937f
C102 VP.n59 B 0.027937f
C103 VP.n60 B 0.027937f
C104 VP.n61 B 0.023872f
C105 VP.n62 B 0.053008f
C106 VP.n63 B 0.039019f
C107 VP.n64 B 0.027937f
C108 VP.n65 B 0.027937f
C109 VP.n66 B 0.039019f
C110 VP.n67 B 0.053008f
C111 VP.n68 B 0.023872f
C112 VP.n69 B 0.027937f
C113 VP.n70 B 0.027937f
C114 VP.n71 B 0.027937f
C115 VP.n72 B 0.03288f
C116 VP.n73 B 0.330522f
C117 VP.n74 B 0.045157f
C118 VP.n75 B 0.046021f
C119 VP.n76 B 0.027937f
C120 VP.n77 B 0.027937f
C121 VP.n78 B 0.027937f
C122 VP.n79 B 0.051806f
C123 VP.n80 B 0.026742f
C124 VP.n81 B 0.400515f
C125 VP.n82 B 0.032108f
C126 VDD2.t9 B 1.08689f
C127 VDD2.t5 B 0.102128f
C128 VDD2.t3 B 0.102128f
C129 VDD2.n0 B 0.846617f
C130 VDD2.n1 B 0.747427f
C131 VDD2.t2 B 0.102128f
C132 VDD2.t0 B 0.102128f
C133 VDD2.n2 B 0.856096f
C134 VDD2.n3 B 2.02553f
C135 VDD2.t6 B 1.07614f
C136 VDD2.n4 B 2.17666f
C137 VDD2.t7 B 0.102128f
C138 VDD2.t8 B 0.102128f
C139 VDD2.n5 B 0.84662f
C140 VDD2.n6 B 0.374452f
C141 VDD2.t1 B 0.102128f
C142 VDD2.t4 B 0.102128f
C143 VDD2.n7 B 0.856066f
C144 VTAIL.t18 B 0.126122f
C145 VTAIL.t16 B 0.126122f
C146 VTAIL.n0 B 0.975294f
C147 VTAIL.n1 B 0.536998f
C148 VTAIL.t6 B 1.24503f
C149 VTAIL.n2 B 0.652265f
C150 VTAIL.t2 B 0.126122f
C151 VTAIL.t7 B 0.126122f
C152 VTAIL.n3 B 0.975294f
C153 VTAIL.n4 B 0.628193f
C154 VTAIL.t0 B 0.126122f
C155 VTAIL.t9 B 0.126122f
C156 VTAIL.n5 B 0.975294f
C157 VTAIL.n6 B 1.637f
C158 VTAIL.t14 B 0.126122f
C159 VTAIL.t11 B 0.126122f
C160 VTAIL.n7 B 0.9753f
C161 VTAIL.n8 B 1.63699f
C162 VTAIL.t19 B 0.126122f
C163 VTAIL.t13 B 0.126122f
C164 VTAIL.n9 B 0.9753f
C165 VTAIL.n10 B 0.628188f
C166 VTAIL.t10 B 1.24503f
C167 VTAIL.n11 B 0.65226f
C168 VTAIL.t8 B 0.126122f
C169 VTAIL.t4 B 0.126122f
C170 VTAIL.n12 B 0.9753f
C171 VTAIL.n13 B 0.578021f
C172 VTAIL.t3 B 0.126122f
C173 VTAIL.t5 B 0.126122f
C174 VTAIL.n14 B 0.9753f
C175 VTAIL.n15 B 0.628188f
C176 VTAIL.t1 B 1.24502f
C177 VTAIL.n16 B 1.52612f
C178 VTAIL.t12 B 1.24503f
C179 VTAIL.n17 B 1.52612f
C180 VTAIL.t17 B 0.126122f
C181 VTAIL.t15 B 0.126122f
C182 VTAIL.n18 B 0.975294f
C183 VTAIL.n19 B 0.484108f
C184 VN.n0 B 0.027402f
C185 VN.t9 B 0.844867f
C186 VN.n1 B 0.034527f
C187 VN.n2 B 0.027402f
C188 VN.t7 B 0.844867f
C189 VN.n3 B 0.055073f
C190 VN.n4 B 0.027402f
C191 VN.t6 B 0.844867f
C192 VN.n5 B 0.324201f
C193 VN.n6 B 0.027402f
C194 VN.n7 B 0.055073f
C195 VN.t0 B 0.993608f
C196 VN.n8 B 0.389753f
C197 VN.t4 B 0.844867f
C198 VN.n9 B 0.38513f
C199 VN.n10 B 0.032251f
C200 VN.n11 B 0.206143f
C201 VN.n12 B 0.027402f
C202 VN.n13 B 0.027402f
C203 VN.n14 B 0.023416f
C204 VN.n15 B 0.051994f
C205 VN.n16 B 0.038272f
C206 VN.n17 B 0.027402f
C207 VN.n18 B 0.027402f
C208 VN.n19 B 0.038272f
C209 VN.n20 B 0.051994f
C210 VN.n21 B 0.023416f
C211 VN.n22 B 0.027402f
C212 VN.n23 B 0.027402f
C213 VN.n24 B 0.027402f
C214 VN.n25 B 0.032251f
C215 VN.n26 B 0.324201f
C216 VN.n27 B 0.044293f
C217 VN.n28 B 0.045141f
C218 VN.n29 B 0.027402f
C219 VN.n30 B 0.027402f
C220 VN.n31 B 0.027402f
C221 VN.n32 B 0.050815f
C222 VN.n33 B 0.026231f
C223 VN.n34 B 0.392855f
C224 VN.n35 B 0.031493f
C225 VN.n36 B 0.027402f
C226 VN.t3 B 0.844867f
C227 VN.n37 B 0.034527f
C228 VN.n38 B 0.027402f
C229 VN.t2 B 0.844867f
C230 VN.n39 B 0.055073f
C231 VN.n40 B 0.027402f
C232 VN.t1 B 0.844867f
C233 VN.n41 B 0.324201f
C234 VN.n42 B 0.027402f
C235 VN.n43 B 0.055073f
C236 VN.t5 B 0.993608f
C237 VN.n44 B 0.389753f
C238 VN.t8 B 0.844867f
C239 VN.n45 B 0.38513f
C240 VN.n46 B 0.032251f
C241 VN.n47 B 0.206143f
C242 VN.n48 B 0.027402f
C243 VN.n49 B 0.027402f
C244 VN.n50 B 0.023416f
C245 VN.n51 B 0.051994f
C246 VN.n52 B 0.038272f
C247 VN.n53 B 0.027402f
C248 VN.n54 B 0.027402f
C249 VN.n55 B 0.038272f
C250 VN.n56 B 0.051994f
C251 VN.n57 B 0.023416f
C252 VN.n58 B 0.027402f
C253 VN.n59 B 0.027402f
C254 VN.n60 B 0.027402f
C255 VN.n61 B 0.032251f
C256 VN.n62 B 0.324201f
C257 VN.n63 B 0.044293f
C258 VN.n64 B 0.045141f
C259 VN.n65 B 0.027402f
C260 VN.n66 B 0.027402f
C261 VN.n67 B 0.027402f
C262 VN.n68 B 0.050815f
C263 VN.n69 B 0.026231f
C264 VN.n70 B 0.392855f
C265 VN.n71 B 1.30573f
.ends

