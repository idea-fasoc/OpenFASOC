* NGSPICE file created from diff_pair_sample_0324.ext - technology: sky130A

.subckt diff_pair_sample_0324 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0 ps=0 w=0.58 l=3.64
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0.2262 ps=1.94 w=0.58 l=3.64
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0 ps=0 w=0.58 l=3.64
X3 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0.2262 ps=1.94 w=0.58 l=3.64
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0 ps=0 w=0.58 l=3.64
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0.2262 ps=1.94 w=0.58 l=3.64
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0.2262 ps=1.94 w=0.58 l=3.64
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2262 pd=1.94 as=0 ps=0 w=0.58 l=3.64
R0 B.n391 B.n390 585
R1 B.n125 B.n73 585
R2 B.n124 B.n123 585
R3 B.n122 B.n121 585
R4 B.n120 B.n119 585
R5 B.n118 B.n117 585
R6 B.n116 B.n115 585
R7 B.n114 B.n113 585
R8 B.n112 B.n111 585
R9 B.n110 B.n109 585
R10 B.n108 B.n107 585
R11 B.n106 B.n105 585
R12 B.n104 B.n103 585
R13 B.n102 B.n101 585
R14 B.n100 B.n99 585
R15 B.n98 B.n97 585
R16 B.n96 B.n95 585
R17 B.n94 B.n93 585
R18 B.n92 B.n91 585
R19 B.n90 B.n89 585
R20 B.n88 B.n87 585
R21 B.n86 B.n85 585
R22 B.n84 B.n83 585
R23 B.n82 B.n81 585
R24 B.n61 B.n60 585
R25 B.n396 B.n395 585
R26 B.n389 B.n74 585
R27 B.n74 B.n58 585
R28 B.n388 B.n57 585
R29 B.n400 B.n57 585
R30 B.n387 B.n56 585
R31 B.n401 B.n56 585
R32 B.n386 B.n55 585
R33 B.n402 B.n55 585
R34 B.n385 B.n384 585
R35 B.n384 B.n51 585
R36 B.n383 B.n50 585
R37 B.n408 B.n50 585
R38 B.n382 B.n49 585
R39 B.n409 B.n49 585
R40 B.n381 B.n48 585
R41 B.n410 B.n48 585
R42 B.n380 B.n379 585
R43 B.n379 B.n44 585
R44 B.n378 B.n43 585
R45 B.n416 B.n43 585
R46 B.n377 B.n42 585
R47 B.n417 B.n42 585
R48 B.n376 B.n41 585
R49 B.n418 B.n41 585
R50 B.n375 B.n374 585
R51 B.n374 B.n37 585
R52 B.n373 B.n36 585
R53 B.n424 B.n36 585
R54 B.n372 B.n35 585
R55 B.n425 B.n35 585
R56 B.n371 B.n34 585
R57 B.n426 B.n34 585
R58 B.n370 B.n369 585
R59 B.n369 B.n30 585
R60 B.n368 B.n29 585
R61 B.n432 B.n29 585
R62 B.n367 B.n28 585
R63 B.n433 B.n28 585
R64 B.n366 B.n27 585
R65 B.n434 B.n27 585
R66 B.n365 B.n364 585
R67 B.n364 B.n23 585
R68 B.n363 B.n22 585
R69 B.n440 B.n22 585
R70 B.n362 B.n21 585
R71 B.n441 B.n21 585
R72 B.n361 B.n20 585
R73 B.n442 B.n20 585
R74 B.n360 B.n359 585
R75 B.n359 B.n19 585
R76 B.n358 B.n15 585
R77 B.n448 B.n15 585
R78 B.n357 B.n14 585
R79 B.n449 B.n14 585
R80 B.n356 B.n13 585
R81 B.n450 B.n13 585
R82 B.n355 B.n354 585
R83 B.n354 B.n12 585
R84 B.n353 B.n352 585
R85 B.n353 B.n8 585
R86 B.n351 B.n7 585
R87 B.n457 B.n7 585
R88 B.n350 B.n6 585
R89 B.n458 B.n6 585
R90 B.n349 B.n5 585
R91 B.n459 B.n5 585
R92 B.n348 B.n347 585
R93 B.n347 B.n4 585
R94 B.n346 B.n126 585
R95 B.n346 B.n345 585
R96 B.n336 B.n127 585
R97 B.n128 B.n127 585
R98 B.n338 B.n337 585
R99 B.n339 B.n338 585
R100 B.n335 B.n133 585
R101 B.n133 B.n132 585
R102 B.n334 B.n333 585
R103 B.n333 B.n332 585
R104 B.n135 B.n134 585
R105 B.n325 B.n135 585
R106 B.n324 B.n323 585
R107 B.n326 B.n324 585
R108 B.n322 B.n140 585
R109 B.n140 B.n139 585
R110 B.n321 B.n320 585
R111 B.n320 B.n319 585
R112 B.n142 B.n141 585
R113 B.n143 B.n142 585
R114 B.n312 B.n311 585
R115 B.n313 B.n312 585
R116 B.n310 B.n148 585
R117 B.n148 B.n147 585
R118 B.n309 B.n308 585
R119 B.n308 B.n307 585
R120 B.n150 B.n149 585
R121 B.n151 B.n150 585
R122 B.n300 B.n299 585
R123 B.n301 B.n300 585
R124 B.n298 B.n156 585
R125 B.n156 B.n155 585
R126 B.n297 B.n296 585
R127 B.n296 B.n295 585
R128 B.n158 B.n157 585
R129 B.n159 B.n158 585
R130 B.n288 B.n287 585
R131 B.n289 B.n288 585
R132 B.n286 B.n164 585
R133 B.n164 B.n163 585
R134 B.n285 B.n284 585
R135 B.n284 B.n283 585
R136 B.n166 B.n165 585
R137 B.n167 B.n166 585
R138 B.n276 B.n275 585
R139 B.n277 B.n276 585
R140 B.n274 B.n172 585
R141 B.n172 B.n171 585
R142 B.n273 B.n272 585
R143 B.n272 B.n271 585
R144 B.n174 B.n173 585
R145 B.n175 B.n174 585
R146 B.n264 B.n263 585
R147 B.n265 B.n264 585
R148 B.n262 B.n180 585
R149 B.n180 B.n179 585
R150 B.n261 B.n260 585
R151 B.n260 B.n259 585
R152 B.n182 B.n181 585
R153 B.n183 B.n182 585
R154 B.n255 B.n254 585
R155 B.n186 B.n185 585
R156 B.n251 B.n250 585
R157 B.n252 B.n251 585
R158 B.n249 B.n199 585
R159 B.n248 B.n247 585
R160 B.n246 B.n245 585
R161 B.n244 B.n243 585
R162 B.n242 B.n241 585
R163 B.n239 B.n238 585
R164 B.n237 B.n236 585
R165 B.n235 B.n234 585
R166 B.n233 B.n232 585
R167 B.n231 B.n230 585
R168 B.n229 B.n228 585
R169 B.n227 B.n226 585
R170 B.n225 B.n224 585
R171 B.n223 B.n222 585
R172 B.n221 B.n220 585
R173 B.n218 B.n217 585
R174 B.n216 B.n215 585
R175 B.n214 B.n213 585
R176 B.n212 B.n211 585
R177 B.n210 B.n209 585
R178 B.n208 B.n207 585
R179 B.n206 B.n205 585
R180 B.n204 B.n198 585
R181 B.n252 B.n198 585
R182 B.n256 B.n184 585
R183 B.n184 B.n183 585
R184 B.n258 B.n257 585
R185 B.n259 B.n258 585
R186 B.n178 B.n177 585
R187 B.n179 B.n178 585
R188 B.n267 B.n266 585
R189 B.n266 B.n265 585
R190 B.n268 B.n176 585
R191 B.n176 B.n175 585
R192 B.n270 B.n269 585
R193 B.n271 B.n270 585
R194 B.n170 B.n169 585
R195 B.n171 B.n170 585
R196 B.n279 B.n278 585
R197 B.n278 B.n277 585
R198 B.n280 B.n168 585
R199 B.n168 B.n167 585
R200 B.n282 B.n281 585
R201 B.n283 B.n282 585
R202 B.n162 B.n161 585
R203 B.n163 B.n162 585
R204 B.n291 B.n290 585
R205 B.n290 B.n289 585
R206 B.n292 B.n160 585
R207 B.n160 B.n159 585
R208 B.n294 B.n293 585
R209 B.n295 B.n294 585
R210 B.n154 B.n153 585
R211 B.n155 B.n154 585
R212 B.n303 B.n302 585
R213 B.n302 B.n301 585
R214 B.n304 B.n152 585
R215 B.n152 B.n151 585
R216 B.n306 B.n305 585
R217 B.n307 B.n306 585
R218 B.n146 B.n145 585
R219 B.n147 B.n146 585
R220 B.n315 B.n314 585
R221 B.n314 B.n313 585
R222 B.n316 B.n144 585
R223 B.n144 B.n143 585
R224 B.n318 B.n317 585
R225 B.n319 B.n318 585
R226 B.n138 B.n137 585
R227 B.n139 B.n138 585
R228 B.n328 B.n327 585
R229 B.n327 B.n326 585
R230 B.n329 B.n136 585
R231 B.n325 B.n136 585
R232 B.n331 B.n330 585
R233 B.n332 B.n331 585
R234 B.n131 B.n130 585
R235 B.n132 B.n131 585
R236 B.n341 B.n340 585
R237 B.n340 B.n339 585
R238 B.n342 B.n129 585
R239 B.n129 B.n128 585
R240 B.n344 B.n343 585
R241 B.n345 B.n344 585
R242 B.n3 B.n0 585
R243 B.n4 B.n3 585
R244 B.n456 B.n1 585
R245 B.n457 B.n456 585
R246 B.n455 B.n454 585
R247 B.n455 B.n8 585
R248 B.n453 B.n9 585
R249 B.n12 B.n9 585
R250 B.n452 B.n451 585
R251 B.n451 B.n450 585
R252 B.n11 B.n10 585
R253 B.n449 B.n11 585
R254 B.n447 B.n446 585
R255 B.n448 B.n447 585
R256 B.n445 B.n16 585
R257 B.n19 B.n16 585
R258 B.n444 B.n443 585
R259 B.n443 B.n442 585
R260 B.n18 B.n17 585
R261 B.n441 B.n18 585
R262 B.n439 B.n438 585
R263 B.n440 B.n439 585
R264 B.n437 B.n24 585
R265 B.n24 B.n23 585
R266 B.n436 B.n435 585
R267 B.n435 B.n434 585
R268 B.n26 B.n25 585
R269 B.n433 B.n26 585
R270 B.n431 B.n430 585
R271 B.n432 B.n431 585
R272 B.n429 B.n31 585
R273 B.n31 B.n30 585
R274 B.n428 B.n427 585
R275 B.n427 B.n426 585
R276 B.n33 B.n32 585
R277 B.n425 B.n33 585
R278 B.n423 B.n422 585
R279 B.n424 B.n423 585
R280 B.n421 B.n38 585
R281 B.n38 B.n37 585
R282 B.n420 B.n419 585
R283 B.n419 B.n418 585
R284 B.n40 B.n39 585
R285 B.n417 B.n40 585
R286 B.n415 B.n414 585
R287 B.n416 B.n415 585
R288 B.n413 B.n45 585
R289 B.n45 B.n44 585
R290 B.n412 B.n411 585
R291 B.n411 B.n410 585
R292 B.n47 B.n46 585
R293 B.n409 B.n47 585
R294 B.n407 B.n406 585
R295 B.n408 B.n407 585
R296 B.n405 B.n52 585
R297 B.n52 B.n51 585
R298 B.n404 B.n403 585
R299 B.n403 B.n402 585
R300 B.n54 B.n53 585
R301 B.n401 B.n54 585
R302 B.n399 B.n398 585
R303 B.n400 B.n399 585
R304 B.n397 B.n59 585
R305 B.n59 B.n58 585
R306 B.n460 B.n459 585
R307 B.n458 B.n2 585
R308 B.n395 B.n59 463.671
R309 B.n391 B.n74 463.671
R310 B.n198 B.n182 463.671
R311 B.n254 B.n184 463.671
R312 B.n78 B.t14 317.077
R313 B.n75 B.t8 317.077
R314 B.n202 B.t12 317.077
R315 B.n200 B.t5 317.077
R316 B.n393 B.n392 256.663
R317 B.n393 B.n72 256.663
R318 B.n393 B.n71 256.663
R319 B.n393 B.n70 256.663
R320 B.n393 B.n69 256.663
R321 B.n393 B.n68 256.663
R322 B.n393 B.n67 256.663
R323 B.n393 B.n66 256.663
R324 B.n393 B.n65 256.663
R325 B.n393 B.n64 256.663
R326 B.n393 B.n63 256.663
R327 B.n393 B.n62 256.663
R328 B.n394 B.n393 256.663
R329 B.n253 B.n252 256.663
R330 B.n252 B.n187 256.663
R331 B.n252 B.n188 256.663
R332 B.n252 B.n189 256.663
R333 B.n252 B.n190 256.663
R334 B.n252 B.n191 256.663
R335 B.n252 B.n192 256.663
R336 B.n252 B.n193 256.663
R337 B.n252 B.n194 256.663
R338 B.n252 B.n195 256.663
R339 B.n252 B.n196 256.663
R340 B.n252 B.n197 256.663
R341 B.n462 B.n461 256.663
R342 B.n79 B.t15 240.083
R343 B.n76 B.t9 240.083
R344 B.n203 B.t11 240.083
R345 B.n201 B.t4 240.083
R346 B.n252 B.n183 227.327
R347 B.n393 B.n58 227.327
R348 B.n78 B.t13 210.222
R349 B.n75 B.t6 210.222
R350 B.n202 B.t10 210.222
R351 B.n200 B.t2 210.222
R352 B.n81 B.n61 163.367
R353 B.n85 B.n84 163.367
R354 B.n89 B.n88 163.367
R355 B.n93 B.n92 163.367
R356 B.n97 B.n96 163.367
R357 B.n101 B.n100 163.367
R358 B.n105 B.n104 163.367
R359 B.n109 B.n108 163.367
R360 B.n113 B.n112 163.367
R361 B.n117 B.n116 163.367
R362 B.n121 B.n120 163.367
R363 B.n123 B.n73 163.367
R364 B.n260 B.n182 163.367
R365 B.n260 B.n180 163.367
R366 B.n264 B.n180 163.367
R367 B.n264 B.n174 163.367
R368 B.n272 B.n174 163.367
R369 B.n272 B.n172 163.367
R370 B.n276 B.n172 163.367
R371 B.n276 B.n166 163.367
R372 B.n284 B.n166 163.367
R373 B.n284 B.n164 163.367
R374 B.n288 B.n164 163.367
R375 B.n288 B.n158 163.367
R376 B.n296 B.n158 163.367
R377 B.n296 B.n156 163.367
R378 B.n300 B.n156 163.367
R379 B.n300 B.n150 163.367
R380 B.n308 B.n150 163.367
R381 B.n308 B.n148 163.367
R382 B.n312 B.n148 163.367
R383 B.n312 B.n142 163.367
R384 B.n320 B.n142 163.367
R385 B.n320 B.n140 163.367
R386 B.n324 B.n140 163.367
R387 B.n324 B.n135 163.367
R388 B.n333 B.n135 163.367
R389 B.n333 B.n133 163.367
R390 B.n338 B.n133 163.367
R391 B.n338 B.n127 163.367
R392 B.n346 B.n127 163.367
R393 B.n347 B.n346 163.367
R394 B.n347 B.n5 163.367
R395 B.n6 B.n5 163.367
R396 B.n7 B.n6 163.367
R397 B.n353 B.n7 163.367
R398 B.n354 B.n353 163.367
R399 B.n354 B.n13 163.367
R400 B.n14 B.n13 163.367
R401 B.n15 B.n14 163.367
R402 B.n359 B.n15 163.367
R403 B.n359 B.n20 163.367
R404 B.n21 B.n20 163.367
R405 B.n22 B.n21 163.367
R406 B.n364 B.n22 163.367
R407 B.n364 B.n27 163.367
R408 B.n28 B.n27 163.367
R409 B.n29 B.n28 163.367
R410 B.n369 B.n29 163.367
R411 B.n369 B.n34 163.367
R412 B.n35 B.n34 163.367
R413 B.n36 B.n35 163.367
R414 B.n374 B.n36 163.367
R415 B.n374 B.n41 163.367
R416 B.n42 B.n41 163.367
R417 B.n43 B.n42 163.367
R418 B.n379 B.n43 163.367
R419 B.n379 B.n48 163.367
R420 B.n49 B.n48 163.367
R421 B.n50 B.n49 163.367
R422 B.n384 B.n50 163.367
R423 B.n384 B.n55 163.367
R424 B.n56 B.n55 163.367
R425 B.n57 B.n56 163.367
R426 B.n74 B.n57 163.367
R427 B.n251 B.n186 163.367
R428 B.n251 B.n199 163.367
R429 B.n247 B.n246 163.367
R430 B.n243 B.n242 163.367
R431 B.n238 B.n237 163.367
R432 B.n234 B.n233 163.367
R433 B.n230 B.n229 163.367
R434 B.n226 B.n225 163.367
R435 B.n222 B.n221 163.367
R436 B.n217 B.n216 163.367
R437 B.n213 B.n212 163.367
R438 B.n209 B.n208 163.367
R439 B.n205 B.n198 163.367
R440 B.n258 B.n184 163.367
R441 B.n258 B.n178 163.367
R442 B.n266 B.n178 163.367
R443 B.n266 B.n176 163.367
R444 B.n270 B.n176 163.367
R445 B.n270 B.n170 163.367
R446 B.n278 B.n170 163.367
R447 B.n278 B.n168 163.367
R448 B.n282 B.n168 163.367
R449 B.n282 B.n162 163.367
R450 B.n290 B.n162 163.367
R451 B.n290 B.n160 163.367
R452 B.n294 B.n160 163.367
R453 B.n294 B.n154 163.367
R454 B.n302 B.n154 163.367
R455 B.n302 B.n152 163.367
R456 B.n306 B.n152 163.367
R457 B.n306 B.n146 163.367
R458 B.n314 B.n146 163.367
R459 B.n314 B.n144 163.367
R460 B.n318 B.n144 163.367
R461 B.n318 B.n138 163.367
R462 B.n327 B.n138 163.367
R463 B.n327 B.n136 163.367
R464 B.n331 B.n136 163.367
R465 B.n331 B.n131 163.367
R466 B.n340 B.n131 163.367
R467 B.n340 B.n129 163.367
R468 B.n344 B.n129 163.367
R469 B.n344 B.n3 163.367
R470 B.n460 B.n3 163.367
R471 B.n456 B.n2 163.367
R472 B.n456 B.n455 163.367
R473 B.n455 B.n9 163.367
R474 B.n451 B.n9 163.367
R475 B.n451 B.n11 163.367
R476 B.n447 B.n11 163.367
R477 B.n447 B.n16 163.367
R478 B.n443 B.n16 163.367
R479 B.n443 B.n18 163.367
R480 B.n439 B.n18 163.367
R481 B.n439 B.n24 163.367
R482 B.n435 B.n24 163.367
R483 B.n435 B.n26 163.367
R484 B.n431 B.n26 163.367
R485 B.n431 B.n31 163.367
R486 B.n427 B.n31 163.367
R487 B.n427 B.n33 163.367
R488 B.n423 B.n33 163.367
R489 B.n423 B.n38 163.367
R490 B.n419 B.n38 163.367
R491 B.n419 B.n40 163.367
R492 B.n415 B.n40 163.367
R493 B.n415 B.n45 163.367
R494 B.n411 B.n45 163.367
R495 B.n411 B.n47 163.367
R496 B.n407 B.n47 163.367
R497 B.n407 B.n52 163.367
R498 B.n403 B.n52 163.367
R499 B.n403 B.n54 163.367
R500 B.n399 B.n54 163.367
R501 B.n399 B.n59 163.367
R502 B.n259 B.n183 127.754
R503 B.n259 B.n179 127.754
R504 B.n265 B.n179 127.754
R505 B.n265 B.n175 127.754
R506 B.n271 B.n175 127.754
R507 B.n271 B.n171 127.754
R508 B.n277 B.n171 127.754
R509 B.n277 B.n167 127.754
R510 B.n283 B.n167 127.754
R511 B.n289 B.n163 127.754
R512 B.n289 B.n159 127.754
R513 B.n295 B.n159 127.754
R514 B.n295 B.n155 127.754
R515 B.n301 B.n155 127.754
R516 B.n301 B.n151 127.754
R517 B.n307 B.n151 127.754
R518 B.n307 B.n147 127.754
R519 B.n313 B.n147 127.754
R520 B.n313 B.n143 127.754
R521 B.n319 B.n143 127.754
R522 B.n319 B.n139 127.754
R523 B.n326 B.n139 127.754
R524 B.n326 B.n325 127.754
R525 B.n332 B.n132 127.754
R526 B.n339 B.n132 127.754
R527 B.n339 B.n128 127.754
R528 B.n345 B.n128 127.754
R529 B.n345 B.n4 127.754
R530 B.n459 B.n4 127.754
R531 B.n459 B.n458 127.754
R532 B.n458 B.n457 127.754
R533 B.n457 B.n8 127.754
R534 B.n12 B.n8 127.754
R535 B.n450 B.n12 127.754
R536 B.n450 B.n449 127.754
R537 B.n449 B.n448 127.754
R538 B.n442 B.n19 127.754
R539 B.n442 B.n441 127.754
R540 B.n441 B.n440 127.754
R541 B.n440 B.n23 127.754
R542 B.n434 B.n23 127.754
R543 B.n434 B.n433 127.754
R544 B.n433 B.n432 127.754
R545 B.n432 B.n30 127.754
R546 B.n426 B.n30 127.754
R547 B.n426 B.n425 127.754
R548 B.n425 B.n424 127.754
R549 B.n424 B.n37 127.754
R550 B.n418 B.n37 127.754
R551 B.n418 B.n417 127.754
R552 B.n416 B.n44 127.754
R553 B.n410 B.n44 127.754
R554 B.n410 B.n409 127.754
R555 B.n409 B.n408 127.754
R556 B.n408 B.n51 127.754
R557 B.n402 B.n51 127.754
R558 B.n402 B.n401 127.754
R559 B.n401 B.n400 127.754
R560 B.n400 B.n58 127.754
R561 B.n332 B.t0 120.24
R562 B.n448 B.t1 120.24
R563 B.t3 B.n163 105.21
R564 B.n417 B.t7 105.21
R565 B.n79 B.n78 76.9944
R566 B.n76 B.n75 76.9944
R567 B.n203 B.n202 76.9944
R568 B.n201 B.n200 76.9944
R569 B.n395 B.n394 71.676
R570 B.n81 B.n62 71.676
R571 B.n85 B.n63 71.676
R572 B.n89 B.n64 71.676
R573 B.n93 B.n65 71.676
R574 B.n97 B.n66 71.676
R575 B.n101 B.n67 71.676
R576 B.n105 B.n68 71.676
R577 B.n109 B.n69 71.676
R578 B.n113 B.n70 71.676
R579 B.n117 B.n71 71.676
R580 B.n121 B.n72 71.676
R581 B.n392 B.n73 71.676
R582 B.n392 B.n391 71.676
R583 B.n123 B.n72 71.676
R584 B.n120 B.n71 71.676
R585 B.n116 B.n70 71.676
R586 B.n112 B.n69 71.676
R587 B.n108 B.n68 71.676
R588 B.n104 B.n67 71.676
R589 B.n100 B.n66 71.676
R590 B.n96 B.n65 71.676
R591 B.n92 B.n64 71.676
R592 B.n88 B.n63 71.676
R593 B.n84 B.n62 71.676
R594 B.n394 B.n61 71.676
R595 B.n254 B.n253 71.676
R596 B.n199 B.n187 71.676
R597 B.n246 B.n188 71.676
R598 B.n242 B.n189 71.676
R599 B.n237 B.n190 71.676
R600 B.n233 B.n191 71.676
R601 B.n229 B.n192 71.676
R602 B.n225 B.n193 71.676
R603 B.n221 B.n194 71.676
R604 B.n216 B.n195 71.676
R605 B.n212 B.n196 71.676
R606 B.n208 B.n197 71.676
R607 B.n253 B.n186 71.676
R608 B.n247 B.n187 71.676
R609 B.n243 B.n188 71.676
R610 B.n238 B.n189 71.676
R611 B.n234 B.n190 71.676
R612 B.n230 B.n191 71.676
R613 B.n226 B.n192 71.676
R614 B.n222 B.n193 71.676
R615 B.n217 B.n194 71.676
R616 B.n213 B.n195 71.676
R617 B.n209 B.n196 71.676
R618 B.n205 B.n197 71.676
R619 B.n461 B.n460 71.676
R620 B.n461 B.n2 71.676
R621 B.n80 B.n79 59.5399
R622 B.n77 B.n76 59.5399
R623 B.n219 B.n203 59.5399
R624 B.n240 B.n201 59.5399
R625 B.n256 B.n255 30.1273
R626 B.n204 B.n181 30.1273
R627 B.n390 B.n389 30.1273
R628 B.n397 B.n396 30.1273
R629 B.n283 B.t3 22.5453
R630 B.t7 B.n416 22.5453
R631 B B.n462 18.0485
R632 B.n257 B.n256 10.6151
R633 B.n257 B.n177 10.6151
R634 B.n267 B.n177 10.6151
R635 B.n268 B.n267 10.6151
R636 B.n269 B.n268 10.6151
R637 B.n269 B.n169 10.6151
R638 B.n279 B.n169 10.6151
R639 B.n280 B.n279 10.6151
R640 B.n281 B.n280 10.6151
R641 B.n281 B.n161 10.6151
R642 B.n291 B.n161 10.6151
R643 B.n292 B.n291 10.6151
R644 B.n293 B.n292 10.6151
R645 B.n293 B.n153 10.6151
R646 B.n303 B.n153 10.6151
R647 B.n304 B.n303 10.6151
R648 B.n305 B.n304 10.6151
R649 B.n305 B.n145 10.6151
R650 B.n315 B.n145 10.6151
R651 B.n316 B.n315 10.6151
R652 B.n317 B.n316 10.6151
R653 B.n317 B.n137 10.6151
R654 B.n328 B.n137 10.6151
R655 B.n329 B.n328 10.6151
R656 B.n330 B.n329 10.6151
R657 B.n330 B.n130 10.6151
R658 B.n341 B.n130 10.6151
R659 B.n342 B.n341 10.6151
R660 B.n343 B.n342 10.6151
R661 B.n343 B.n0 10.6151
R662 B.n255 B.n185 10.6151
R663 B.n250 B.n185 10.6151
R664 B.n250 B.n249 10.6151
R665 B.n249 B.n248 10.6151
R666 B.n248 B.n245 10.6151
R667 B.n245 B.n244 10.6151
R668 B.n244 B.n241 10.6151
R669 B.n239 B.n236 10.6151
R670 B.n236 B.n235 10.6151
R671 B.n235 B.n232 10.6151
R672 B.n232 B.n231 10.6151
R673 B.n231 B.n228 10.6151
R674 B.n228 B.n227 10.6151
R675 B.n227 B.n224 10.6151
R676 B.n224 B.n223 10.6151
R677 B.n223 B.n220 10.6151
R678 B.n218 B.n215 10.6151
R679 B.n215 B.n214 10.6151
R680 B.n214 B.n211 10.6151
R681 B.n211 B.n210 10.6151
R682 B.n210 B.n207 10.6151
R683 B.n207 B.n206 10.6151
R684 B.n206 B.n204 10.6151
R685 B.n261 B.n181 10.6151
R686 B.n262 B.n261 10.6151
R687 B.n263 B.n262 10.6151
R688 B.n263 B.n173 10.6151
R689 B.n273 B.n173 10.6151
R690 B.n274 B.n273 10.6151
R691 B.n275 B.n274 10.6151
R692 B.n275 B.n165 10.6151
R693 B.n285 B.n165 10.6151
R694 B.n286 B.n285 10.6151
R695 B.n287 B.n286 10.6151
R696 B.n287 B.n157 10.6151
R697 B.n297 B.n157 10.6151
R698 B.n298 B.n297 10.6151
R699 B.n299 B.n298 10.6151
R700 B.n299 B.n149 10.6151
R701 B.n309 B.n149 10.6151
R702 B.n310 B.n309 10.6151
R703 B.n311 B.n310 10.6151
R704 B.n311 B.n141 10.6151
R705 B.n321 B.n141 10.6151
R706 B.n322 B.n321 10.6151
R707 B.n323 B.n322 10.6151
R708 B.n323 B.n134 10.6151
R709 B.n334 B.n134 10.6151
R710 B.n335 B.n334 10.6151
R711 B.n337 B.n335 10.6151
R712 B.n337 B.n336 10.6151
R713 B.n336 B.n126 10.6151
R714 B.n348 B.n126 10.6151
R715 B.n349 B.n348 10.6151
R716 B.n350 B.n349 10.6151
R717 B.n351 B.n350 10.6151
R718 B.n352 B.n351 10.6151
R719 B.n355 B.n352 10.6151
R720 B.n356 B.n355 10.6151
R721 B.n357 B.n356 10.6151
R722 B.n358 B.n357 10.6151
R723 B.n360 B.n358 10.6151
R724 B.n361 B.n360 10.6151
R725 B.n362 B.n361 10.6151
R726 B.n363 B.n362 10.6151
R727 B.n365 B.n363 10.6151
R728 B.n366 B.n365 10.6151
R729 B.n367 B.n366 10.6151
R730 B.n368 B.n367 10.6151
R731 B.n370 B.n368 10.6151
R732 B.n371 B.n370 10.6151
R733 B.n372 B.n371 10.6151
R734 B.n373 B.n372 10.6151
R735 B.n375 B.n373 10.6151
R736 B.n376 B.n375 10.6151
R737 B.n377 B.n376 10.6151
R738 B.n378 B.n377 10.6151
R739 B.n380 B.n378 10.6151
R740 B.n381 B.n380 10.6151
R741 B.n382 B.n381 10.6151
R742 B.n383 B.n382 10.6151
R743 B.n385 B.n383 10.6151
R744 B.n386 B.n385 10.6151
R745 B.n387 B.n386 10.6151
R746 B.n388 B.n387 10.6151
R747 B.n389 B.n388 10.6151
R748 B.n454 B.n1 10.6151
R749 B.n454 B.n453 10.6151
R750 B.n453 B.n452 10.6151
R751 B.n452 B.n10 10.6151
R752 B.n446 B.n10 10.6151
R753 B.n446 B.n445 10.6151
R754 B.n445 B.n444 10.6151
R755 B.n444 B.n17 10.6151
R756 B.n438 B.n17 10.6151
R757 B.n438 B.n437 10.6151
R758 B.n437 B.n436 10.6151
R759 B.n436 B.n25 10.6151
R760 B.n430 B.n25 10.6151
R761 B.n430 B.n429 10.6151
R762 B.n429 B.n428 10.6151
R763 B.n428 B.n32 10.6151
R764 B.n422 B.n32 10.6151
R765 B.n422 B.n421 10.6151
R766 B.n421 B.n420 10.6151
R767 B.n420 B.n39 10.6151
R768 B.n414 B.n39 10.6151
R769 B.n414 B.n413 10.6151
R770 B.n413 B.n412 10.6151
R771 B.n412 B.n46 10.6151
R772 B.n406 B.n46 10.6151
R773 B.n406 B.n405 10.6151
R774 B.n405 B.n404 10.6151
R775 B.n404 B.n53 10.6151
R776 B.n398 B.n53 10.6151
R777 B.n398 B.n397 10.6151
R778 B.n396 B.n60 10.6151
R779 B.n82 B.n60 10.6151
R780 B.n83 B.n82 10.6151
R781 B.n86 B.n83 10.6151
R782 B.n87 B.n86 10.6151
R783 B.n90 B.n87 10.6151
R784 B.n91 B.n90 10.6151
R785 B.n95 B.n94 10.6151
R786 B.n98 B.n95 10.6151
R787 B.n99 B.n98 10.6151
R788 B.n102 B.n99 10.6151
R789 B.n103 B.n102 10.6151
R790 B.n106 B.n103 10.6151
R791 B.n107 B.n106 10.6151
R792 B.n110 B.n107 10.6151
R793 B.n111 B.n110 10.6151
R794 B.n115 B.n114 10.6151
R795 B.n118 B.n115 10.6151
R796 B.n119 B.n118 10.6151
R797 B.n122 B.n119 10.6151
R798 B.n124 B.n122 10.6151
R799 B.n125 B.n124 10.6151
R800 B.n390 B.n125 10.6151
R801 B.n241 B.n240 9.36635
R802 B.n219 B.n218 9.36635
R803 B.n91 B.n80 9.36635
R804 B.n114 B.n77 9.36635
R805 B.n462 B.n0 8.11757
R806 B.n462 B.n1 8.11757
R807 B.n325 B.t0 7.51544
R808 B.n19 B.t1 7.51544
R809 B.n240 B.n239 1.24928
R810 B.n220 B.n219 1.24928
R811 B.n94 B.n80 1.24928
R812 B.n111 B.n77 1.24928
R813 VP.n0 VP.t0 77.5867
R814 VP.n0 VP.t1 38.8237
R815 VP VP.n0 0.621233
R816 VTAIL.n3 VTAIL.t0 250.935
R817 VTAIL.n0 VTAIL.t3 250.935
R818 VTAIL.n2 VTAIL.t2 250.935
R819 VTAIL.n1 VTAIL.t1 250.935
R820 VTAIL.n1 VTAIL.n0 19.7117
R821 VTAIL.n3 VTAIL.n2 16.2893
R822 VTAIL.n2 VTAIL.n1 2.18153
R823 VTAIL VTAIL.n0 1.38412
R824 VTAIL VTAIL.n3 0.797914
R825 VDD1 VDD1.t0 299.998
R826 VDD1 VDD1.t1 268.527
R827 VN VN.t1 77.399
R828 VN VN.t0 39.4444
R829 VDD2.n0 VDD2.t1 298.618
R830 VDD2.n0 VDD2.t0 267.615
R831 VDD2 VDD2.n0 0.914293
C0 VDD2 VDD1 0.786817f
C1 VP VN 3.84695f
C2 VTAIL VP 1.06937f
C3 VP VDD2 0.385745f
C4 VP VDD1 0.621405f
C5 VTAIL VN 1.05525f
C6 VDD2 VN 0.394741f
C7 VDD1 VN 0.156646f
C8 VTAIL VDD2 2.4688f
C9 VTAIL VDD1 2.40849f
C10 VDD2 B 2.757202f
C11 VDD1 B 5.01424f
C12 VTAIL B 2.587028f
C13 VN B 8.92891f
C14 VP B 6.625517f
C15 VDD2.t1 B 0.141694f
C16 VDD2.t0 B 0.048599f
C17 VDD2.n0 B 2.12025f
C18 VN.t0 B 0.396095f
C19 VN.t1 B 1.12618f
C20 VDD1.t1 B 0.045597f
C21 VDD1.t0 B 0.142991f
C22 VTAIL.t3 B 0.05805f
C23 VTAIL.n0 B 1.25214f
C24 VTAIL.t1 B 0.05805f
C25 VTAIL.n1 B 1.32649f
C26 VTAIL.t2 B 0.05805f
C27 VTAIL.n2 B 1.00741f
C28 VTAIL.t0 B 0.05805f
C29 VTAIL.n3 B 0.878419f
C30 VP.t0 B 1.14009f
C31 VP.t1 B 0.396262f
C32 VP.n0 B 2.13282f
.ends

