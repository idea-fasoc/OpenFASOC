* NGSPICE file created from diff_pair_sample_0504.ext - technology: sky130A

.subckt diff_pair_sample_0504 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.15975 pd=19.48 as=7.4685 ps=39.08 w=19.15 l=3.76
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=0 ps=0 w=19.15 l=3.76
X2 VTAIL.t5 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=3.15975 ps=19.48 w=19.15 l=3.76
X3 VTAIL.t6 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=3.15975 ps=19.48 w=19.15 l=3.76
X4 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.15975 pd=19.48 as=7.4685 ps=39.08 w=19.15 l=3.76
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=0 ps=0 w=19.15 l=3.76
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=0 ps=0 w=19.15 l=3.76
X7 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.15975 pd=19.48 as=7.4685 ps=39.08 w=19.15 l=3.76
X8 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=3.15975 ps=19.48 w=19.15 l=3.76
X9 VDD2.t0 VN.t3 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.15975 pd=19.48 as=7.4685 ps=39.08 w=19.15 l=3.76
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=0 ps=0 w=19.15 l=3.76
X11 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.4685 pd=39.08 as=3.15975 ps=19.48 w=19.15 l=3.76
R0 VN.n1 VN.t3 156.429
R1 VN.n0 VN.t1 156.429
R2 VN.n0 VN.t0 155.089
R3 VN.n1 VN.t2 155.089
R4 VN VN.n1 57.3621
R5 VN VN.n0 1.88864
R6 VTAIL.n5 VTAIL.t1 48.2395
R7 VTAIL.n4 VTAIL.t7 48.2395
R8 VTAIL.n3 VTAIL.t6 48.2395
R9 VTAIL.n7 VTAIL.t4 48.2394
R10 VTAIL.n0 VTAIL.t5 48.2394
R11 VTAIL.n1 VTAIL.t0 48.2394
R12 VTAIL.n2 VTAIL.t3 48.2394
R13 VTAIL.n6 VTAIL.t2 48.2394
R14 VTAIL.n7 VTAIL.n6 32.4014
R15 VTAIL.n3 VTAIL.n2 32.4014
R16 VTAIL.n4 VTAIL.n3 3.52636
R17 VTAIL.n6 VTAIL.n5 3.52636
R18 VTAIL.n2 VTAIL.n1 3.52636
R19 VTAIL VTAIL.n0 1.82162
R20 VTAIL VTAIL.n7 1.70524
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 114.684
R24 VDD2.n2 VDD2.n1 63.8842
R25 VDD2.n1 VDD2.t1 1.03444
R26 VDD2.n1 VDD2.t0 1.03444
R27 VDD2.n0 VDD2.t2 1.03444
R28 VDD2.n0 VDD2.t3 1.03444
R29 VDD2 VDD2.n2 0.0586897
R30 B.n1040 B.n1039 585
R31 B.n1041 B.n1040 585
R32 B.n421 B.n150 585
R33 B.n420 B.n419 585
R34 B.n418 B.n417 585
R35 B.n416 B.n415 585
R36 B.n414 B.n413 585
R37 B.n412 B.n411 585
R38 B.n410 B.n409 585
R39 B.n408 B.n407 585
R40 B.n406 B.n405 585
R41 B.n404 B.n403 585
R42 B.n402 B.n401 585
R43 B.n400 B.n399 585
R44 B.n398 B.n397 585
R45 B.n396 B.n395 585
R46 B.n394 B.n393 585
R47 B.n392 B.n391 585
R48 B.n390 B.n389 585
R49 B.n388 B.n387 585
R50 B.n386 B.n385 585
R51 B.n384 B.n383 585
R52 B.n382 B.n381 585
R53 B.n380 B.n379 585
R54 B.n378 B.n377 585
R55 B.n376 B.n375 585
R56 B.n374 B.n373 585
R57 B.n372 B.n371 585
R58 B.n370 B.n369 585
R59 B.n368 B.n367 585
R60 B.n366 B.n365 585
R61 B.n364 B.n363 585
R62 B.n362 B.n361 585
R63 B.n360 B.n359 585
R64 B.n358 B.n357 585
R65 B.n356 B.n355 585
R66 B.n354 B.n353 585
R67 B.n352 B.n351 585
R68 B.n350 B.n349 585
R69 B.n348 B.n347 585
R70 B.n346 B.n345 585
R71 B.n344 B.n343 585
R72 B.n342 B.n341 585
R73 B.n340 B.n339 585
R74 B.n338 B.n337 585
R75 B.n336 B.n335 585
R76 B.n334 B.n333 585
R77 B.n332 B.n331 585
R78 B.n330 B.n329 585
R79 B.n328 B.n327 585
R80 B.n326 B.n325 585
R81 B.n324 B.n323 585
R82 B.n322 B.n321 585
R83 B.n320 B.n319 585
R84 B.n318 B.n317 585
R85 B.n316 B.n315 585
R86 B.n314 B.n313 585
R87 B.n312 B.n311 585
R88 B.n310 B.n309 585
R89 B.n308 B.n307 585
R90 B.n306 B.n305 585
R91 B.n304 B.n303 585
R92 B.n302 B.n301 585
R93 B.n300 B.n299 585
R94 B.n298 B.n297 585
R95 B.n296 B.n295 585
R96 B.n294 B.n293 585
R97 B.n292 B.n291 585
R98 B.n290 B.n289 585
R99 B.n288 B.n287 585
R100 B.n286 B.n285 585
R101 B.n284 B.n283 585
R102 B.n282 B.n281 585
R103 B.n279 B.n278 585
R104 B.n277 B.n276 585
R105 B.n275 B.n274 585
R106 B.n273 B.n272 585
R107 B.n271 B.n270 585
R108 B.n269 B.n268 585
R109 B.n267 B.n266 585
R110 B.n265 B.n264 585
R111 B.n263 B.n262 585
R112 B.n261 B.n260 585
R113 B.n259 B.n258 585
R114 B.n257 B.n256 585
R115 B.n255 B.n254 585
R116 B.n253 B.n252 585
R117 B.n251 B.n250 585
R118 B.n249 B.n248 585
R119 B.n247 B.n246 585
R120 B.n245 B.n244 585
R121 B.n243 B.n242 585
R122 B.n241 B.n240 585
R123 B.n239 B.n238 585
R124 B.n237 B.n236 585
R125 B.n235 B.n234 585
R126 B.n233 B.n232 585
R127 B.n231 B.n230 585
R128 B.n229 B.n228 585
R129 B.n227 B.n226 585
R130 B.n225 B.n224 585
R131 B.n223 B.n222 585
R132 B.n221 B.n220 585
R133 B.n219 B.n218 585
R134 B.n217 B.n216 585
R135 B.n215 B.n214 585
R136 B.n213 B.n212 585
R137 B.n211 B.n210 585
R138 B.n209 B.n208 585
R139 B.n207 B.n206 585
R140 B.n205 B.n204 585
R141 B.n203 B.n202 585
R142 B.n201 B.n200 585
R143 B.n199 B.n198 585
R144 B.n197 B.n196 585
R145 B.n195 B.n194 585
R146 B.n193 B.n192 585
R147 B.n191 B.n190 585
R148 B.n189 B.n188 585
R149 B.n187 B.n186 585
R150 B.n185 B.n184 585
R151 B.n183 B.n182 585
R152 B.n181 B.n180 585
R153 B.n179 B.n178 585
R154 B.n177 B.n176 585
R155 B.n175 B.n174 585
R156 B.n173 B.n172 585
R157 B.n171 B.n170 585
R158 B.n169 B.n168 585
R159 B.n167 B.n166 585
R160 B.n165 B.n164 585
R161 B.n163 B.n162 585
R162 B.n161 B.n160 585
R163 B.n159 B.n158 585
R164 B.n157 B.n156 585
R165 B.n81 B.n80 585
R166 B.n1038 B.n82 585
R167 B.n1042 B.n82 585
R168 B.n1037 B.n1036 585
R169 B.n1036 B.n78 585
R170 B.n1035 B.n77 585
R171 B.n1048 B.n77 585
R172 B.n1034 B.n76 585
R173 B.n1049 B.n76 585
R174 B.n1033 B.n75 585
R175 B.n1050 B.n75 585
R176 B.n1032 B.n1031 585
R177 B.n1031 B.n71 585
R178 B.n1030 B.n70 585
R179 B.n1056 B.n70 585
R180 B.n1029 B.n69 585
R181 B.n1057 B.n69 585
R182 B.n1028 B.n68 585
R183 B.n1058 B.n68 585
R184 B.n1027 B.n1026 585
R185 B.n1026 B.n67 585
R186 B.n1025 B.n63 585
R187 B.n1064 B.n63 585
R188 B.n1024 B.n62 585
R189 B.n1065 B.n62 585
R190 B.n1023 B.n61 585
R191 B.n1066 B.n61 585
R192 B.n1022 B.n1021 585
R193 B.n1021 B.n57 585
R194 B.n1020 B.n56 585
R195 B.n1072 B.n56 585
R196 B.n1019 B.n55 585
R197 B.n1073 B.n55 585
R198 B.n1018 B.n54 585
R199 B.n1074 B.n54 585
R200 B.n1017 B.n1016 585
R201 B.n1016 B.n50 585
R202 B.n1015 B.n49 585
R203 B.n1080 B.n49 585
R204 B.n1014 B.n48 585
R205 B.n1081 B.n48 585
R206 B.n1013 B.n47 585
R207 B.n1082 B.n47 585
R208 B.n1012 B.n1011 585
R209 B.n1011 B.n43 585
R210 B.n1010 B.n42 585
R211 B.n1088 B.n42 585
R212 B.n1009 B.n41 585
R213 B.n1089 B.n41 585
R214 B.n1008 B.n40 585
R215 B.n1090 B.n40 585
R216 B.n1007 B.n1006 585
R217 B.n1006 B.n36 585
R218 B.n1005 B.n35 585
R219 B.n1096 B.n35 585
R220 B.n1004 B.n34 585
R221 B.n1097 B.n34 585
R222 B.n1003 B.n33 585
R223 B.n1098 B.n33 585
R224 B.n1002 B.n1001 585
R225 B.n1001 B.n29 585
R226 B.n1000 B.n28 585
R227 B.n1104 B.n28 585
R228 B.n999 B.n27 585
R229 B.n1105 B.n27 585
R230 B.n998 B.n26 585
R231 B.n1106 B.n26 585
R232 B.n997 B.n996 585
R233 B.n996 B.n22 585
R234 B.n995 B.n21 585
R235 B.n1112 B.n21 585
R236 B.n994 B.n20 585
R237 B.n1113 B.n20 585
R238 B.n993 B.n19 585
R239 B.n1114 B.n19 585
R240 B.n992 B.n991 585
R241 B.n991 B.n15 585
R242 B.n990 B.n14 585
R243 B.n1120 B.n14 585
R244 B.n989 B.n13 585
R245 B.n1121 B.n13 585
R246 B.n988 B.n12 585
R247 B.n1122 B.n12 585
R248 B.n987 B.n986 585
R249 B.n986 B.n8 585
R250 B.n985 B.n7 585
R251 B.n1128 B.n7 585
R252 B.n984 B.n6 585
R253 B.n1129 B.n6 585
R254 B.n983 B.n5 585
R255 B.n1130 B.n5 585
R256 B.n982 B.n981 585
R257 B.n981 B.n4 585
R258 B.n980 B.n422 585
R259 B.n980 B.n979 585
R260 B.n970 B.n423 585
R261 B.n424 B.n423 585
R262 B.n972 B.n971 585
R263 B.n973 B.n972 585
R264 B.n969 B.n429 585
R265 B.n429 B.n428 585
R266 B.n968 B.n967 585
R267 B.n967 B.n966 585
R268 B.n431 B.n430 585
R269 B.n432 B.n431 585
R270 B.n959 B.n958 585
R271 B.n960 B.n959 585
R272 B.n957 B.n437 585
R273 B.n437 B.n436 585
R274 B.n956 B.n955 585
R275 B.n955 B.n954 585
R276 B.n439 B.n438 585
R277 B.n440 B.n439 585
R278 B.n947 B.n946 585
R279 B.n948 B.n947 585
R280 B.n945 B.n445 585
R281 B.n445 B.n444 585
R282 B.n944 B.n943 585
R283 B.n943 B.n942 585
R284 B.n447 B.n446 585
R285 B.n448 B.n447 585
R286 B.n935 B.n934 585
R287 B.n936 B.n935 585
R288 B.n933 B.n453 585
R289 B.n453 B.n452 585
R290 B.n932 B.n931 585
R291 B.n931 B.n930 585
R292 B.n455 B.n454 585
R293 B.n456 B.n455 585
R294 B.n923 B.n922 585
R295 B.n924 B.n923 585
R296 B.n921 B.n461 585
R297 B.n461 B.n460 585
R298 B.n920 B.n919 585
R299 B.n919 B.n918 585
R300 B.n463 B.n462 585
R301 B.n464 B.n463 585
R302 B.n911 B.n910 585
R303 B.n912 B.n911 585
R304 B.n909 B.n469 585
R305 B.n469 B.n468 585
R306 B.n908 B.n907 585
R307 B.n907 B.n906 585
R308 B.n471 B.n470 585
R309 B.n472 B.n471 585
R310 B.n899 B.n898 585
R311 B.n900 B.n899 585
R312 B.n897 B.n477 585
R313 B.n477 B.n476 585
R314 B.n896 B.n895 585
R315 B.n895 B.n894 585
R316 B.n479 B.n478 585
R317 B.n480 B.n479 585
R318 B.n887 B.n886 585
R319 B.n888 B.n887 585
R320 B.n885 B.n485 585
R321 B.n485 B.n484 585
R322 B.n884 B.n883 585
R323 B.n883 B.n882 585
R324 B.n487 B.n486 585
R325 B.n875 B.n487 585
R326 B.n874 B.n873 585
R327 B.n876 B.n874 585
R328 B.n872 B.n492 585
R329 B.n492 B.n491 585
R330 B.n871 B.n870 585
R331 B.n870 B.n869 585
R332 B.n494 B.n493 585
R333 B.n495 B.n494 585
R334 B.n862 B.n861 585
R335 B.n863 B.n862 585
R336 B.n860 B.n500 585
R337 B.n500 B.n499 585
R338 B.n859 B.n858 585
R339 B.n858 B.n857 585
R340 B.n502 B.n501 585
R341 B.n503 B.n502 585
R342 B.n850 B.n849 585
R343 B.n851 B.n850 585
R344 B.n506 B.n505 585
R345 B.n579 B.n578 585
R346 B.n580 B.n576 585
R347 B.n576 B.n507 585
R348 B.n582 B.n581 585
R349 B.n584 B.n575 585
R350 B.n587 B.n586 585
R351 B.n588 B.n574 585
R352 B.n590 B.n589 585
R353 B.n592 B.n573 585
R354 B.n595 B.n594 585
R355 B.n596 B.n572 585
R356 B.n598 B.n597 585
R357 B.n600 B.n571 585
R358 B.n603 B.n602 585
R359 B.n604 B.n570 585
R360 B.n606 B.n605 585
R361 B.n608 B.n569 585
R362 B.n611 B.n610 585
R363 B.n612 B.n568 585
R364 B.n614 B.n613 585
R365 B.n616 B.n567 585
R366 B.n619 B.n618 585
R367 B.n620 B.n566 585
R368 B.n622 B.n621 585
R369 B.n624 B.n565 585
R370 B.n627 B.n626 585
R371 B.n628 B.n564 585
R372 B.n630 B.n629 585
R373 B.n632 B.n563 585
R374 B.n635 B.n634 585
R375 B.n636 B.n562 585
R376 B.n638 B.n637 585
R377 B.n640 B.n561 585
R378 B.n643 B.n642 585
R379 B.n644 B.n560 585
R380 B.n646 B.n645 585
R381 B.n648 B.n559 585
R382 B.n651 B.n650 585
R383 B.n652 B.n558 585
R384 B.n654 B.n653 585
R385 B.n656 B.n557 585
R386 B.n659 B.n658 585
R387 B.n660 B.n556 585
R388 B.n662 B.n661 585
R389 B.n664 B.n555 585
R390 B.n667 B.n666 585
R391 B.n668 B.n554 585
R392 B.n670 B.n669 585
R393 B.n672 B.n553 585
R394 B.n675 B.n674 585
R395 B.n676 B.n552 585
R396 B.n678 B.n677 585
R397 B.n680 B.n551 585
R398 B.n683 B.n682 585
R399 B.n684 B.n550 585
R400 B.n686 B.n685 585
R401 B.n688 B.n549 585
R402 B.n691 B.n690 585
R403 B.n692 B.n548 585
R404 B.n694 B.n693 585
R405 B.n696 B.n547 585
R406 B.n699 B.n698 585
R407 B.n700 B.n544 585
R408 B.n703 B.n702 585
R409 B.n705 B.n543 585
R410 B.n708 B.n707 585
R411 B.n709 B.n542 585
R412 B.n711 B.n710 585
R413 B.n713 B.n541 585
R414 B.n716 B.n715 585
R415 B.n717 B.n540 585
R416 B.n722 B.n721 585
R417 B.n724 B.n539 585
R418 B.n727 B.n726 585
R419 B.n728 B.n538 585
R420 B.n730 B.n729 585
R421 B.n732 B.n537 585
R422 B.n735 B.n734 585
R423 B.n736 B.n536 585
R424 B.n738 B.n737 585
R425 B.n740 B.n535 585
R426 B.n743 B.n742 585
R427 B.n744 B.n534 585
R428 B.n746 B.n745 585
R429 B.n748 B.n533 585
R430 B.n751 B.n750 585
R431 B.n752 B.n532 585
R432 B.n754 B.n753 585
R433 B.n756 B.n531 585
R434 B.n759 B.n758 585
R435 B.n760 B.n530 585
R436 B.n762 B.n761 585
R437 B.n764 B.n529 585
R438 B.n767 B.n766 585
R439 B.n768 B.n528 585
R440 B.n770 B.n769 585
R441 B.n772 B.n527 585
R442 B.n775 B.n774 585
R443 B.n776 B.n526 585
R444 B.n778 B.n777 585
R445 B.n780 B.n525 585
R446 B.n783 B.n782 585
R447 B.n784 B.n524 585
R448 B.n786 B.n785 585
R449 B.n788 B.n523 585
R450 B.n791 B.n790 585
R451 B.n792 B.n522 585
R452 B.n794 B.n793 585
R453 B.n796 B.n521 585
R454 B.n799 B.n798 585
R455 B.n800 B.n520 585
R456 B.n802 B.n801 585
R457 B.n804 B.n519 585
R458 B.n807 B.n806 585
R459 B.n808 B.n518 585
R460 B.n810 B.n809 585
R461 B.n812 B.n517 585
R462 B.n815 B.n814 585
R463 B.n816 B.n516 585
R464 B.n818 B.n817 585
R465 B.n820 B.n515 585
R466 B.n823 B.n822 585
R467 B.n824 B.n514 585
R468 B.n826 B.n825 585
R469 B.n828 B.n513 585
R470 B.n831 B.n830 585
R471 B.n832 B.n512 585
R472 B.n834 B.n833 585
R473 B.n836 B.n511 585
R474 B.n839 B.n838 585
R475 B.n840 B.n510 585
R476 B.n842 B.n841 585
R477 B.n844 B.n509 585
R478 B.n847 B.n846 585
R479 B.n848 B.n508 585
R480 B.n853 B.n852 585
R481 B.n852 B.n851 585
R482 B.n854 B.n504 585
R483 B.n504 B.n503 585
R484 B.n856 B.n855 585
R485 B.n857 B.n856 585
R486 B.n498 B.n497 585
R487 B.n499 B.n498 585
R488 B.n865 B.n864 585
R489 B.n864 B.n863 585
R490 B.n866 B.n496 585
R491 B.n496 B.n495 585
R492 B.n868 B.n867 585
R493 B.n869 B.n868 585
R494 B.n490 B.n489 585
R495 B.n491 B.n490 585
R496 B.n878 B.n877 585
R497 B.n877 B.n876 585
R498 B.n879 B.n488 585
R499 B.n875 B.n488 585
R500 B.n881 B.n880 585
R501 B.n882 B.n881 585
R502 B.n483 B.n482 585
R503 B.n484 B.n483 585
R504 B.n890 B.n889 585
R505 B.n889 B.n888 585
R506 B.n891 B.n481 585
R507 B.n481 B.n480 585
R508 B.n893 B.n892 585
R509 B.n894 B.n893 585
R510 B.n475 B.n474 585
R511 B.n476 B.n475 585
R512 B.n902 B.n901 585
R513 B.n901 B.n900 585
R514 B.n903 B.n473 585
R515 B.n473 B.n472 585
R516 B.n905 B.n904 585
R517 B.n906 B.n905 585
R518 B.n467 B.n466 585
R519 B.n468 B.n467 585
R520 B.n914 B.n913 585
R521 B.n913 B.n912 585
R522 B.n915 B.n465 585
R523 B.n465 B.n464 585
R524 B.n917 B.n916 585
R525 B.n918 B.n917 585
R526 B.n459 B.n458 585
R527 B.n460 B.n459 585
R528 B.n926 B.n925 585
R529 B.n925 B.n924 585
R530 B.n927 B.n457 585
R531 B.n457 B.n456 585
R532 B.n929 B.n928 585
R533 B.n930 B.n929 585
R534 B.n451 B.n450 585
R535 B.n452 B.n451 585
R536 B.n938 B.n937 585
R537 B.n937 B.n936 585
R538 B.n939 B.n449 585
R539 B.n449 B.n448 585
R540 B.n941 B.n940 585
R541 B.n942 B.n941 585
R542 B.n443 B.n442 585
R543 B.n444 B.n443 585
R544 B.n950 B.n949 585
R545 B.n949 B.n948 585
R546 B.n951 B.n441 585
R547 B.n441 B.n440 585
R548 B.n953 B.n952 585
R549 B.n954 B.n953 585
R550 B.n435 B.n434 585
R551 B.n436 B.n435 585
R552 B.n962 B.n961 585
R553 B.n961 B.n960 585
R554 B.n963 B.n433 585
R555 B.n433 B.n432 585
R556 B.n965 B.n964 585
R557 B.n966 B.n965 585
R558 B.n427 B.n426 585
R559 B.n428 B.n427 585
R560 B.n975 B.n974 585
R561 B.n974 B.n973 585
R562 B.n976 B.n425 585
R563 B.n425 B.n424 585
R564 B.n978 B.n977 585
R565 B.n979 B.n978 585
R566 B.n2 B.n0 585
R567 B.n4 B.n2 585
R568 B.n3 B.n1 585
R569 B.n1129 B.n3 585
R570 B.n1127 B.n1126 585
R571 B.n1128 B.n1127 585
R572 B.n1125 B.n9 585
R573 B.n9 B.n8 585
R574 B.n1124 B.n1123 585
R575 B.n1123 B.n1122 585
R576 B.n11 B.n10 585
R577 B.n1121 B.n11 585
R578 B.n1119 B.n1118 585
R579 B.n1120 B.n1119 585
R580 B.n1117 B.n16 585
R581 B.n16 B.n15 585
R582 B.n1116 B.n1115 585
R583 B.n1115 B.n1114 585
R584 B.n18 B.n17 585
R585 B.n1113 B.n18 585
R586 B.n1111 B.n1110 585
R587 B.n1112 B.n1111 585
R588 B.n1109 B.n23 585
R589 B.n23 B.n22 585
R590 B.n1108 B.n1107 585
R591 B.n1107 B.n1106 585
R592 B.n25 B.n24 585
R593 B.n1105 B.n25 585
R594 B.n1103 B.n1102 585
R595 B.n1104 B.n1103 585
R596 B.n1101 B.n30 585
R597 B.n30 B.n29 585
R598 B.n1100 B.n1099 585
R599 B.n1099 B.n1098 585
R600 B.n32 B.n31 585
R601 B.n1097 B.n32 585
R602 B.n1095 B.n1094 585
R603 B.n1096 B.n1095 585
R604 B.n1093 B.n37 585
R605 B.n37 B.n36 585
R606 B.n1092 B.n1091 585
R607 B.n1091 B.n1090 585
R608 B.n39 B.n38 585
R609 B.n1089 B.n39 585
R610 B.n1087 B.n1086 585
R611 B.n1088 B.n1087 585
R612 B.n1085 B.n44 585
R613 B.n44 B.n43 585
R614 B.n1084 B.n1083 585
R615 B.n1083 B.n1082 585
R616 B.n46 B.n45 585
R617 B.n1081 B.n46 585
R618 B.n1079 B.n1078 585
R619 B.n1080 B.n1079 585
R620 B.n1077 B.n51 585
R621 B.n51 B.n50 585
R622 B.n1076 B.n1075 585
R623 B.n1075 B.n1074 585
R624 B.n53 B.n52 585
R625 B.n1073 B.n53 585
R626 B.n1071 B.n1070 585
R627 B.n1072 B.n1071 585
R628 B.n1069 B.n58 585
R629 B.n58 B.n57 585
R630 B.n1068 B.n1067 585
R631 B.n1067 B.n1066 585
R632 B.n60 B.n59 585
R633 B.n1065 B.n60 585
R634 B.n1063 B.n1062 585
R635 B.n1064 B.n1063 585
R636 B.n1061 B.n64 585
R637 B.n67 B.n64 585
R638 B.n1060 B.n1059 585
R639 B.n1059 B.n1058 585
R640 B.n66 B.n65 585
R641 B.n1057 B.n66 585
R642 B.n1055 B.n1054 585
R643 B.n1056 B.n1055 585
R644 B.n1053 B.n72 585
R645 B.n72 B.n71 585
R646 B.n1052 B.n1051 585
R647 B.n1051 B.n1050 585
R648 B.n74 B.n73 585
R649 B.n1049 B.n74 585
R650 B.n1047 B.n1046 585
R651 B.n1048 B.n1047 585
R652 B.n1045 B.n79 585
R653 B.n79 B.n78 585
R654 B.n1044 B.n1043 585
R655 B.n1043 B.n1042 585
R656 B.n1132 B.n1131 585
R657 B.n1131 B.n1130 585
R658 B.n852 B.n506 521.33
R659 B.n1043 B.n81 521.33
R660 B.n850 B.n508 521.33
R661 B.n1040 B.n82 521.33
R662 B.n718 B.t15 332.057
R663 B.n545 B.t4 332.057
R664 B.n154 B.t12 332.057
R665 B.n151 B.t8 332.057
R666 B.n1041 B.n149 256.663
R667 B.n1041 B.n148 256.663
R668 B.n1041 B.n147 256.663
R669 B.n1041 B.n146 256.663
R670 B.n1041 B.n145 256.663
R671 B.n1041 B.n144 256.663
R672 B.n1041 B.n143 256.663
R673 B.n1041 B.n142 256.663
R674 B.n1041 B.n141 256.663
R675 B.n1041 B.n140 256.663
R676 B.n1041 B.n139 256.663
R677 B.n1041 B.n138 256.663
R678 B.n1041 B.n137 256.663
R679 B.n1041 B.n136 256.663
R680 B.n1041 B.n135 256.663
R681 B.n1041 B.n134 256.663
R682 B.n1041 B.n133 256.663
R683 B.n1041 B.n132 256.663
R684 B.n1041 B.n131 256.663
R685 B.n1041 B.n130 256.663
R686 B.n1041 B.n129 256.663
R687 B.n1041 B.n128 256.663
R688 B.n1041 B.n127 256.663
R689 B.n1041 B.n126 256.663
R690 B.n1041 B.n125 256.663
R691 B.n1041 B.n124 256.663
R692 B.n1041 B.n123 256.663
R693 B.n1041 B.n122 256.663
R694 B.n1041 B.n121 256.663
R695 B.n1041 B.n120 256.663
R696 B.n1041 B.n119 256.663
R697 B.n1041 B.n118 256.663
R698 B.n1041 B.n117 256.663
R699 B.n1041 B.n116 256.663
R700 B.n1041 B.n115 256.663
R701 B.n1041 B.n114 256.663
R702 B.n1041 B.n113 256.663
R703 B.n1041 B.n112 256.663
R704 B.n1041 B.n111 256.663
R705 B.n1041 B.n110 256.663
R706 B.n1041 B.n109 256.663
R707 B.n1041 B.n108 256.663
R708 B.n1041 B.n107 256.663
R709 B.n1041 B.n106 256.663
R710 B.n1041 B.n105 256.663
R711 B.n1041 B.n104 256.663
R712 B.n1041 B.n103 256.663
R713 B.n1041 B.n102 256.663
R714 B.n1041 B.n101 256.663
R715 B.n1041 B.n100 256.663
R716 B.n1041 B.n99 256.663
R717 B.n1041 B.n98 256.663
R718 B.n1041 B.n97 256.663
R719 B.n1041 B.n96 256.663
R720 B.n1041 B.n95 256.663
R721 B.n1041 B.n94 256.663
R722 B.n1041 B.n93 256.663
R723 B.n1041 B.n92 256.663
R724 B.n1041 B.n91 256.663
R725 B.n1041 B.n90 256.663
R726 B.n1041 B.n89 256.663
R727 B.n1041 B.n88 256.663
R728 B.n1041 B.n87 256.663
R729 B.n1041 B.n86 256.663
R730 B.n1041 B.n85 256.663
R731 B.n1041 B.n84 256.663
R732 B.n1041 B.n83 256.663
R733 B.n577 B.n507 256.663
R734 B.n583 B.n507 256.663
R735 B.n585 B.n507 256.663
R736 B.n591 B.n507 256.663
R737 B.n593 B.n507 256.663
R738 B.n599 B.n507 256.663
R739 B.n601 B.n507 256.663
R740 B.n607 B.n507 256.663
R741 B.n609 B.n507 256.663
R742 B.n615 B.n507 256.663
R743 B.n617 B.n507 256.663
R744 B.n623 B.n507 256.663
R745 B.n625 B.n507 256.663
R746 B.n631 B.n507 256.663
R747 B.n633 B.n507 256.663
R748 B.n639 B.n507 256.663
R749 B.n641 B.n507 256.663
R750 B.n647 B.n507 256.663
R751 B.n649 B.n507 256.663
R752 B.n655 B.n507 256.663
R753 B.n657 B.n507 256.663
R754 B.n663 B.n507 256.663
R755 B.n665 B.n507 256.663
R756 B.n671 B.n507 256.663
R757 B.n673 B.n507 256.663
R758 B.n679 B.n507 256.663
R759 B.n681 B.n507 256.663
R760 B.n687 B.n507 256.663
R761 B.n689 B.n507 256.663
R762 B.n695 B.n507 256.663
R763 B.n697 B.n507 256.663
R764 B.n704 B.n507 256.663
R765 B.n706 B.n507 256.663
R766 B.n712 B.n507 256.663
R767 B.n714 B.n507 256.663
R768 B.n723 B.n507 256.663
R769 B.n725 B.n507 256.663
R770 B.n731 B.n507 256.663
R771 B.n733 B.n507 256.663
R772 B.n739 B.n507 256.663
R773 B.n741 B.n507 256.663
R774 B.n747 B.n507 256.663
R775 B.n749 B.n507 256.663
R776 B.n755 B.n507 256.663
R777 B.n757 B.n507 256.663
R778 B.n763 B.n507 256.663
R779 B.n765 B.n507 256.663
R780 B.n771 B.n507 256.663
R781 B.n773 B.n507 256.663
R782 B.n779 B.n507 256.663
R783 B.n781 B.n507 256.663
R784 B.n787 B.n507 256.663
R785 B.n789 B.n507 256.663
R786 B.n795 B.n507 256.663
R787 B.n797 B.n507 256.663
R788 B.n803 B.n507 256.663
R789 B.n805 B.n507 256.663
R790 B.n811 B.n507 256.663
R791 B.n813 B.n507 256.663
R792 B.n819 B.n507 256.663
R793 B.n821 B.n507 256.663
R794 B.n827 B.n507 256.663
R795 B.n829 B.n507 256.663
R796 B.n835 B.n507 256.663
R797 B.n837 B.n507 256.663
R798 B.n843 B.n507 256.663
R799 B.n845 B.n507 256.663
R800 B.n852 B.n504 163.367
R801 B.n856 B.n504 163.367
R802 B.n856 B.n498 163.367
R803 B.n864 B.n498 163.367
R804 B.n864 B.n496 163.367
R805 B.n868 B.n496 163.367
R806 B.n868 B.n490 163.367
R807 B.n877 B.n490 163.367
R808 B.n877 B.n488 163.367
R809 B.n881 B.n488 163.367
R810 B.n881 B.n483 163.367
R811 B.n889 B.n483 163.367
R812 B.n889 B.n481 163.367
R813 B.n893 B.n481 163.367
R814 B.n893 B.n475 163.367
R815 B.n901 B.n475 163.367
R816 B.n901 B.n473 163.367
R817 B.n905 B.n473 163.367
R818 B.n905 B.n467 163.367
R819 B.n913 B.n467 163.367
R820 B.n913 B.n465 163.367
R821 B.n917 B.n465 163.367
R822 B.n917 B.n459 163.367
R823 B.n925 B.n459 163.367
R824 B.n925 B.n457 163.367
R825 B.n929 B.n457 163.367
R826 B.n929 B.n451 163.367
R827 B.n937 B.n451 163.367
R828 B.n937 B.n449 163.367
R829 B.n941 B.n449 163.367
R830 B.n941 B.n443 163.367
R831 B.n949 B.n443 163.367
R832 B.n949 B.n441 163.367
R833 B.n953 B.n441 163.367
R834 B.n953 B.n435 163.367
R835 B.n961 B.n435 163.367
R836 B.n961 B.n433 163.367
R837 B.n965 B.n433 163.367
R838 B.n965 B.n427 163.367
R839 B.n974 B.n427 163.367
R840 B.n974 B.n425 163.367
R841 B.n978 B.n425 163.367
R842 B.n978 B.n2 163.367
R843 B.n1131 B.n2 163.367
R844 B.n1131 B.n3 163.367
R845 B.n1127 B.n3 163.367
R846 B.n1127 B.n9 163.367
R847 B.n1123 B.n9 163.367
R848 B.n1123 B.n11 163.367
R849 B.n1119 B.n11 163.367
R850 B.n1119 B.n16 163.367
R851 B.n1115 B.n16 163.367
R852 B.n1115 B.n18 163.367
R853 B.n1111 B.n18 163.367
R854 B.n1111 B.n23 163.367
R855 B.n1107 B.n23 163.367
R856 B.n1107 B.n25 163.367
R857 B.n1103 B.n25 163.367
R858 B.n1103 B.n30 163.367
R859 B.n1099 B.n30 163.367
R860 B.n1099 B.n32 163.367
R861 B.n1095 B.n32 163.367
R862 B.n1095 B.n37 163.367
R863 B.n1091 B.n37 163.367
R864 B.n1091 B.n39 163.367
R865 B.n1087 B.n39 163.367
R866 B.n1087 B.n44 163.367
R867 B.n1083 B.n44 163.367
R868 B.n1083 B.n46 163.367
R869 B.n1079 B.n46 163.367
R870 B.n1079 B.n51 163.367
R871 B.n1075 B.n51 163.367
R872 B.n1075 B.n53 163.367
R873 B.n1071 B.n53 163.367
R874 B.n1071 B.n58 163.367
R875 B.n1067 B.n58 163.367
R876 B.n1067 B.n60 163.367
R877 B.n1063 B.n60 163.367
R878 B.n1063 B.n64 163.367
R879 B.n1059 B.n64 163.367
R880 B.n1059 B.n66 163.367
R881 B.n1055 B.n66 163.367
R882 B.n1055 B.n72 163.367
R883 B.n1051 B.n72 163.367
R884 B.n1051 B.n74 163.367
R885 B.n1047 B.n74 163.367
R886 B.n1047 B.n79 163.367
R887 B.n1043 B.n79 163.367
R888 B.n578 B.n576 163.367
R889 B.n582 B.n576 163.367
R890 B.n586 B.n584 163.367
R891 B.n590 B.n574 163.367
R892 B.n594 B.n592 163.367
R893 B.n598 B.n572 163.367
R894 B.n602 B.n600 163.367
R895 B.n606 B.n570 163.367
R896 B.n610 B.n608 163.367
R897 B.n614 B.n568 163.367
R898 B.n618 B.n616 163.367
R899 B.n622 B.n566 163.367
R900 B.n626 B.n624 163.367
R901 B.n630 B.n564 163.367
R902 B.n634 B.n632 163.367
R903 B.n638 B.n562 163.367
R904 B.n642 B.n640 163.367
R905 B.n646 B.n560 163.367
R906 B.n650 B.n648 163.367
R907 B.n654 B.n558 163.367
R908 B.n658 B.n656 163.367
R909 B.n662 B.n556 163.367
R910 B.n666 B.n664 163.367
R911 B.n670 B.n554 163.367
R912 B.n674 B.n672 163.367
R913 B.n678 B.n552 163.367
R914 B.n682 B.n680 163.367
R915 B.n686 B.n550 163.367
R916 B.n690 B.n688 163.367
R917 B.n694 B.n548 163.367
R918 B.n698 B.n696 163.367
R919 B.n703 B.n544 163.367
R920 B.n707 B.n705 163.367
R921 B.n711 B.n542 163.367
R922 B.n715 B.n713 163.367
R923 B.n722 B.n540 163.367
R924 B.n726 B.n724 163.367
R925 B.n730 B.n538 163.367
R926 B.n734 B.n732 163.367
R927 B.n738 B.n536 163.367
R928 B.n742 B.n740 163.367
R929 B.n746 B.n534 163.367
R930 B.n750 B.n748 163.367
R931 B.n754 B.n532 163.367
R932 B.n758 B.n756 163.367
R933 B.n762 B.n530 163.367
R934 B.n766 B.n764 163.367
R935 B.n770 B.n528 163.367
R936 B.n774 B.n772 163.367
R937 B.n778 B.n526 163.367
R938 B.n782 B.n780 163.367
R939 B.n786 B.n524 163.367
R940 B.n790 B.n788 163.367
R941 B.n794 B.n522 163.367
R942 B.n798 B.n796 163.367
R943 B.n802 B.n520 163.367
R944 B.n806 B.n804 163.367
R945 B.n810 B.n518 163.367
R946 B.n814 B.n812 163.367
R947 B.n818 B.n516 163.367
R948 B.n822 B.n820 163.367
R949 B.n826 B.n514 163.367
R950 B.n830 B.n828 163.367
R951 B.n834 B.n512 163.367
R952 B.n838 B.n836 163.367
R953 B.n842 B.n510 163.367
R954 B.n846 B.n844 163.367
R955 B.n850 B.n502 163.367
R956 B.n858 B.n502 163.367
R957 B.n858 B.n500 163.367
R958 B.n862 B.n500 163.367
R959 B.n862 B.n494 163.367
R960 B.n870 B.n494 163.367
R961 B.n870 B.n492 163.367
R962 B.n874 B.n492 163.367
R963 B.n874 B.n487 163.367
R964 B.n883 B.n487 163.367
R965 B.n883 B.n485 163.367
R966 B.n887 B.n485 163.367
R967 B.n887 B.n479 163.367
R968 B.n895 B.n479 163.367
R969 B.n895 B.n477 163.367
R970 B.n899 B.n477 163.367
R971 B.n899 B.n471 163.367
R972 B.n907 B.n471 163.367
R973 B.n907 B.n469 163.367
R974 B.n911 B.n469 163.367
R975 B.n911 B.n463 163.367
R976 B.n919 B.n463 163.367
R977 B.n919 B.n461 163.367
R978 B.n923 B.n461 163.367
R979 B.n923 B.n455 163.367
R980 B.n931 B.n455 163.367
R981 B.n931 B.n453 163.367
R982 B.n935 B.n453 163.367
R983 B.n935 B.n447 163.367
R984 B.n943 B.n447 163.367
R985 B.n943 B.n445 163.367
R986 B.n947 B.n445 163.367
R987 B.n947 B.n439 163.367
R988 B.n955 B.n439 163.367
R989 B.n955 B.n437 163.367
R990 B.n959 B.n437 163.367
R991 B.n959 B.n431 163.367
R992 B.n967 B.n431 163.367
R993 B.n967 B.n429 163.367
R994 B.n972 B.n429 163.367
R995 B.n972 B.n423 163.367
R996 B.n980 B.n423 163.367
R997 B.n981 B.n980 163.367
R998 B.n981 B.n5 163.367
R999 B.n6 B.n5 163.367
R1000 B.n7 B.n6 163.367
R1001 B.n986 B.n7 163.367
R1002 B.n986 B.n12 163.367
R1003 B.n13 B.n12 163.367
R1004 B.n14 B.n13 163.367
R1005 B.n991 B.n14 163.367
R1006 B.n991 B.n19 163.367
R1007 B.n20 B.n19 163.367
R1008 B.n21 B.n20 163.367
R1009 B.n996 B.n21 163.367
R1010 B.n996 B.n26 163.367
R1011 B.n27 B.n26 163.367
R1012 B.n28 B.n27 163.367
R1013 B.n1001 B.n28 163.367
R1014 B.n1001 B.n33 163.367
R1015 B.n34 B.n33 163.367
R1016 B.n35 B.n34 163.367
R1017 B.n1006 B.n35 163.367
R1018 B.n1006 B.n40 163.367
R1019 B.n41 B.n40 163.367
R1020 B.n42 B.n41 163.367
R1021 B.n1011 B.n42 163.367
R1022 B.n1011 B.n47 163.367
R1023 B.n48 B.n47 163.367
R1024 B.n49 B.n48 163.367
R1025 B.n1016 B.n49 163.367
R1026 B.n1016 B.n54 163.367
R1027 B.n55 B.n54 163.367
R1028 B.n56 B.n55 163.367
R1029 B.n1021 B.n56 163.367
R1030 B.n1021 B.n61 163.367
R1031 B.n62 B.n61 163.367
R1032 B.n63 B.n62 163.367
R1033 B.n1026 B.n63 163.367
R1034 B.n1026 B.n68 163.367
R1035 B.n69 B.n68 163.367
R1036 B.n70 B.n69 163.367
R1037 B.n1031 B.n70 163.367
R1038 B.n1031 B.n75 163.367
R1039 B.n76 B.n75 163.367
R1040 B.n77 B.n76 163.367
R1041 B.n1036 B.n77 163.367
R1042 B.n1036 B.n82 163.367
R1043 B.n158 B.n157 163.367
R1044 B.n162 B.n161 163.367
R1045 B.n166 B.n165 163.367
R1046 B.n170 B.n169 163.367
R1047 B.n174 B.n173 163.367
R1048 B.n178 B.n177 163.367
R1049 B.n182 B.n181 163.367
R1050 B.n186 B.n185 163.367
R1051 B.n190 B.n189 163.367
R1052 B.n194 B.n193 163.367
R1053 B.n198 B.n197 163.367
R1054 B.n202 B.n201 163.367
R1055 B.n206 B.n205 163.367
R1056 B.n210 B.n209 163.367
R1057 B.n214 B.n213 163.367
R1058 B.n218 B.n217 163.367
R1059 B.n222 B.n221 163.367
R1060 B.n226 B.n225 163.367
R1061 B.n230 B.n229 163.367
R1062 B.n234 B.n233 163.367
R1063 B.n238 B.n237 163.367
R1064 B.n242 B.n241 163.367
R1065 B.n246 B.n245 163.367
R1066 B.n250 B.n249 163.367
R1067 B.n254 B.n253 163.367
R1068 B.n258 B.n257 163.367
R1069 B.n262 B.n261 163.367
R1070 B.n266 B.n265 163.367
R1071 B.n270 B.n269 163.367
R1072 B.n274 B.n273 163.367
R1073 B.n278 B.n277 163.367
R1074 B.n283 B.n282 163.367
R1075 B.n287 B.n286 163.367
R1076 B.n291 B.n290 163.367
R1077 B.n295 B.n294 163.367
R1078 B.n299 B.n298 163.367
R1079 B.n303 B.n302 163.367
R1080 B.n307 B.n306 163.367
R1081 B.n311 B.n310 163.367
R1082 B.n315 B.n314 163.367
R1083 B.n319 B.n318 163.367
R1084 B.n323 B.n322 163.367
R1085 B.n327 B.n326 163.367
R1086 B.n331 B.n330 163.367
R1087 B.n335 B.n334 163.367
R1088 B.n339 B.n338 163.367
R1089 B.n343 B.n342 163.367
R1090 B.n347 B.n346 163.367
R1091 B.n351 B.n350 163.367
R1092 B.n355 B.n354 163.367
R1093 B.n359 B.n358 163.367
R1094 B.n363 B.n362 163.367
R1095 B.n367 B.n366 163.367
R1096 B.n371 B.n370 163.367
R1097 B.n375 B.n374 163.367
R1098 B.n379 B.n378 163.367
R1099 B.n383 B.n382 163.367
R1100 B.n387 B.n386 163.367
R1101 B.n391 B.n390 163.367
R1102 B.n395 B.n394 163.367
R1103 B.n399 B.n398 163.367
R1104 B.n403 B.n402 163.367
R1105 B.n407 B.n406 163.367
R1106 B.n411 B.n410 163.367
R1107 B.n415 B.n414 163.367
R1108 B.n419 B.n418 163.367
R1109 B.n1040 B.n150 163.367
R1110 B.n718 B.t17 148.638
R1111 B.n151 B.t10 148.638
R1112 B.n545 B.t7 148.613
R1113 B.n154 B.t13 148.613
R1114 B.n719 B.n718 79.3217
R1115 B.n546 B.n545 79.3217
R1116 B.n155 B.n154 79.3217
R1117 B.n152 B.n151 79.3217
R1118 B.n577 B.n506 71.676
R1119 B.n583 B.n582 71.676
R1120 B.n586 B.n585 71.676
R1121 B.n591 B.n590 71.676
R1122 B.n594 B.n593 71.676
R1123 B.n599 B.n598 71.676
R1124 B.n602 B.n601 71.676
R1125 B.n607 B.n606 71.676
R1126 B.n610 B.n609 71.676
R1127 B.n615 B.n614 71.676
R1128 B.n618 B.n617 71.676
R1129 B.n623 B.n622 71.676
R1130 B.n626 B.n625 71.676
R1131 B.n631 B.n630 71.676
R1132 B.n634 B.n633 71.676
R1133 B.n639 B.n638 71.676
R1134 B.n642 B.n641 71.676
R1135 B.n647 B.n646 71.676
R1136 B.n650 B.n649 71.676
R1137 B.n655 B.n654 71.676
R1138 B.n658 B.n657 71.676
R1139 B.n663 B.n662 71.676
R1140 B.n666 B.n665 71.676
R1141 B.n671 B.n670 71.676
R1142 B.n674 B.n673 71.676
R1143 B.n679 B.n678 71.676
R1144 B.n682 B.n681 71.676
R1145 B.n687 B.n686 71.676
R1146 B.n690 B.n689 71.676
R1147 B.n695 B.n694 71.676
R1148 B.n698 B.n697 71.676
R1149 B.n704 B.n703 71.676
R1150 B.n707 B.n706 71.676
R1151 B.n712 B.n711 71.676
R1152 B.n715 B.n714 71.676
R1153 B.n723 B.n722 71.676
R1154 B.n726 B.n725 71.676
R1155 B.n731 B.n730 71.676
R1156 B.n734 B.n733 71.676
R1157 B.n739 B.n738 71.676
R1158 B.n742 B.n741 71.676
R1159 B.n747 B.n746 71.676
R1160 B.n750 B.n749 71.676
R1161 B.n755 B.n754 71.676
R1162 B.n758 B.n757 71.676
R1163 B.n763 B.n762 71.676
R1164 B.n766 B.n765 71.676
R1165 B.n771 B.n770 71.676
R1166 B.n774 B.n773 71.676
R1167 B.n779 B.n778 71.676
R1168 B.n782 B.n781 71.676
R1169 B.n787 B.n786 71.676
R1170 B.n790 B.n789 71.676
R1171 B.n795 B.n794 71.676
R1172 B.n798 B.n797 71.676
R1173 B.n803 B.n802 71.676
R1174 B.n806 B.n805 71.676
R1175 B.n811 B.n810 71.676
R1176 B.n814 B.n813 71.676
R1177 B.n819 B.n818 71.676
R1178 B.n822 B.n821 71.676
R1179 B.n827 B.n826 71.676
R1180 B.n830 B.n829 71.676
R1181 B.n835 B.n834 71.676
R1182 B.n838 B.n837 71.676
R1183 B.n843 B.n842 71.676
R1184 B.n846 B.n845 71.676
R1185 B.n83 B.n81 71.676
R1186 B.n158 B.n84 71.676
R1187 B.n162 B.n85 71.676
R1188 B.n166 B.n86 71.676
R1189 B.n170 B.n87 71.676
R1190 B.n174 B.n88 71.676
R1191 B.n178 B.n89 71.676
R1192 B.n182 B.n90 71.676
R1193 B.n186 B.n91 71.676
R1194 B.n190 B.n92 71.676
R1195 B.n194 B.n93 71.676
R1196 B.n198 B.n94 71.676
R1197 B.n202 B.n95 71.676
R1198 B.n206 B.n96 71.676
R1199 B.n210 B.n97 71.676
R1200 B.n214 B.n98 71.676
R1201 B.n218 B.n99 71.676
R1202 B.n222 B.n100 71.676
R1203 B.n226 B.n101 71.676
R1204 B.n230 B.n102 71.676
R1205 B.n234 B.n103 71.676
R1206 B.n238 B.n104 71.676
R1207 B.n242 B.n105 71.676
R1208 B.n246 B.n106 71.676
R1209 B.n250 B.n107 71.676
R1210 B.n254 B.n108 71.676
R1211 B.n258 B.n109 71.676
R1212 B.n262 B.n110 71.676
R1213 B.n266 B.n111 71.676
R1214 B.n270 B.n112 71.676
R1215 B.n274 B.n113 71.676
R1216 B.n278 B.n114 71.676
R1217 B.n283 B.n115 71.676
R1218 B.n287 B.n116 71.676
R1219 B.n291 B.n117 71.676
R1220 B.n295 B.n118 71.676
R1221 B.n299 B.n119 71.676
R1222 B.n303 B.n120 71.676
R1223 B.n307 B.n121 71.676
R1224 B.n311 B.n122 71.676
R1225 B.n315 B.n123 71.676
R1226 B.n319 B.n124 71.676
R1227 B.n323 B.n125 71.676
R1228 B.n327 B.n126 71.676
R1229 B.n331 B.n127 71.676
R1230 B.n335 B.n128 71.676
R1231 B.n339 B.n129 71.676
R1232 B.n343 B.n130 71.676
R1233 B.n347 B.n131 71.676
R1234 B.n351 B.n132 71.676
R1235 B.n355 B.n133 71.676
R1236 B.n359 B.n134 71.676
R1237 B.n363 B.n135 71.676
R1238 B.n367 B.n136 71.676
R1239 B.n371 B.n137 71.676
R1240 B.n375 B.n138 71.676
R1241 B.n379 B.n139 71.676
R1242 B.n383 B.n140 71.676
R1243 B.n387 B.n141 71.676
R1244 B.n391 B.n142 71.676
R1245 B.n395 B.n143 71.676
R1246 B.n399 B.n144 71.676
R1247 B.n403 B.n145 71.676
R1248 B.n407 B.n146 71.676
R1249 B.n411 B.n147 71.676
R1250 B.n415 B.n148 71.676
R1251 B.n419 B.n149 71.676
R1252 B.n150 B.n149 71.676
R1253 B.n418 B.n148 71.676
R1254 B.n414 B.n147 71.676
R1255 B.n410 B.n146 71.676
R1256 B.n406 B.n145 71.676
R1257 B.n402 B.n144 71.676
R1258 B.n398 B.n143 71.676
R1259 B.n394 B.n142 71.676
R1260 B.n390 B.n141 71.676
R1261 B.n386 B.n140 71.676
R1262 B.n382 B.n139 71.676
R1263 B.n378 B.n138 71.676
R1264 B.n374 B.n137 71.676
R1265 B.n370 B.n136 71.676
R1266 B.n366 B.n135 71.676
R1267 B.n362 B.n134 71.676
R1268 B.n358 B.n133 71.676
R1269 B.n354 B.n132 71.676
R1270 B.n350 B.n131 71.676
R1271 B.n346 B.n130 71.676
R1272 B.n342 B.n129 71.676
R1273 B.n338 B.n128 71.676
R1274 B.n334 B.n127 71.676
R1275 B.n330 B.n126 71.676
R1276 B.n326 B.n125 71.676
R1277 B.n322 B.n124 71.676
R1278 B.n318 B.n123 71.676
R1279 B.n314 B.n122 71.676
R1280 B.n310 B.n121 71.676
R1281 B.n306 B.n120 71.676
R1282 B.n302 B.n119 71.676
R1283 B.n298 B.n118 71.676
R1284 B.n294 B.n117 71.676
R1285 B.n290 B.n116 71.676
R1286 B.n286 B.n115 71.676
R1287 B.n282 B.n114 71.676
R1288 B.n277 B.n113 71.676
R1289 B.n273 B.n112 71.676
R1290 B.n269 B.n111 71.676
R1291 B.n265 B.n110 71.676
R1292 B.n261 B.n109 71.676
R1293 B.n257 B.n108 71.676
R1294 B.n253 B.n107 71.676
R1295 B.n249 B.n106 71.676
R1296 B.n245 B.n105 71.676
R1297 B.n241 B.n104 71.676
R1298 B.n237 B.n103 71.676
R1299 B.n233 B.n102 71.676
R1300 B.n229 B.n101 71.676
R1301 B.n225 B.n100 71.676
R1302 B.n221 B.n99 71.676
R1303 B.n217 B.n98 71.676
R1304 B.n213 B.n97 71.676
R1305 B.n209 B.n96 71.676
R1306 B.n205 B.n95 71.676
R1307 B.n201 B.n94 71.676
R1308 B.n197 B.n93 71.676
R1309 B.n193 B.n92 71.676
R1310 B.n189 B.n91 71.676
R1311 B.n185 B.n90 71.676
R1312 B.n181 B.n89 71.676
R1313 B.n177 B.n88 71.676
R1314 B.n173 B.n87 71.676
R1315 B.n169 B.n86 71.676
R1316 B.n165 B.n85 71.676
R1317 B.n161 B.n84 71.676
R1318 B.n157 B.n83 71.676
R1319 B.n578 B.n577 71.676
R1320 B.n584 B.n583 71.676
R1321 B.n585 B.n574 71.676
R1322 B.n592 B.n591 71.676
R1323 B.n593 B.n572 71.676
R1324 B.n600 B.n599 71.676
R1325 B.n601 B.n570 71.676
R1326 B.n608 B.n607 71.676
R1327 B.n609 B.n568 71.676
R1328 B.n616 B.n615 71.676
R1329 B.n617 B.n566 71.676
R1330 B.n624 B.n623 71.676
R1331 B.n625 B.n564 71.676
R1332 B.n632 B.n631 71.676
R1333 B.n633 B.n562 71.676
R1334 B.n640 B.n639 71.676
R1335 B.n641 B.n560 71.676
R1336 B.n648 B.n647 71.676
R1337 B.n649 B.n558 71.676
R1338 B.n656 B.n655 71.676
R1339 B.n657 B.n556 71.676
R1340 B.n664 B.n663 71.676
R1341 B.n665 B.n554 71.676
R1342 B.n672 B.n671 71.676
R1343 B.n673 B.n552 71.676
R1344 B.n680 B.n679 71.676
R1345 B.n681 B.n550 71.676
R1346 B.n688 B.n687 71.676
R1347 B.n689 B.n548 71.676
R1348 B.n696 B.n695 71.676
R1349 B.n697 B.n544 71.676
R1350 B.n705 B.n704 71.676
R1351 B.n706 B.n542 71.676
R1352 B.n713 B.n712 71.676
R1353 B.n714 B.n540 71.676
R1354 B.n724 B.n723 71.676
R1355 B.n725 B.n538 71.676
R1356 B.n732 B.n731 71.676
R1357 B.n733 B.n536 71.676
R1358 B.n740 B.n739 71.676
R1359 B.n741 B.n534 71.676
R1360 B.n748 B.n747 71.676
R1361 B.n749 B.n532 71.676
R1362 B.n756 B.n755 71.676
R1363 B.n757 B.n530 71.676
R1364 B.n764 B.n763 71.676
R1365 B.n765 B.n528 71.676
R1366 B.n772 B.n771 71.676
R1367 B.n773 B.n526 71.676
R1368 B.n780 B.n779 71.676
R1369 B.n781 B.n524 71.676
R1370 B.n788 B.n787 71.676
R1371 B.n789 B.n522 71.676
R1372 B.n796 B.n795 71.676
R1373 B.n797 B.n520 71.676
R1374 B.n804 B.n803 71.676
R1375 B.n805 B.n518 71.676
R1376 B.n812 B.n811 71.676
R1377 B.n813 B.n516 71.676
R1378 B.n820 B.n819 71.676
R1379 B.n821 B.n514 71.676
R1380 B.n828 B.n827 71.676
R1381 B.n829 B.n512 71.676
R1382 B.n836 B.n835 71.676
R1383 B.n837 B.n510 71.676
R1384 B.n844 B.n843 71.676
R1385 B.n845 B.n508 71.676
R1386 B.n719 B.t16 69.3177
R1387 B.n152 B.t11 69.3177
R1388 B.n546 B.t6 69.2919
R1389 B.n155 B.t14 69.2919
R1390 B.n851 B.n507 61.6996
R1391 B.n1042 B.n1041 61.6996
R1392 B.n720 B.n719 59.5399
R1393 B.n701 B.n546 59.5399
R1394 B.n280 B.n155 59.5399
R1395 B.n153 B.n152 59.5399
R1396 B.n1044 B.n80 33.8737
R1397 B.n1039 B.n1038 33.8737
R1398 B.n849 B.n848 33.8737
R1399 B.n853 B.n505 33.8737
R1400 B.n851 B.n503 30.6249
R1401 B.n857 B.n503 30.6249
R1402 B.n857 B.n499 30.6249
R1403 B.n863 B.n499 30.6249
R1404 B.n863 B.n495 30.6249
R1405 B.n869 B.n495 30.6249
R1406 B.n869 B.n491 30.6249
R1407 B.n876 B.n491 30.6249
R1408 B.n876 B.n875 30.6249
R1409 B.n882 B.n484 30.6249
R1410 B.n888 B.n484 30.6249
R1411 B.n888 B.n480 30.6249
R1412 B.n894 B.n480 30.6249
R1413 B.n894 B.n476 30.6249
R1414 B.n900 B.n476 30.6249
R1415 B.n900 B.n472 30.6249
R1416 B.n906 B.n472 30.6249
R1417 B.n906 B.n468 30.6249
R1418 B.n912 B.n468 30.6249
R1419 B.n912 B.n464 30.6249
R1420 B.n918 B.n464 30.6249
R1421 B.n918 B.n460 30.6249
R1422 B.n924 B.n460 30.6249
R1423 B.n930 B.n456 30.6249
R1424 B.n930 B.n452 30.6249
R1425 B.n936 B.n452 30.6249
R1426 B.n936 B.n448 30.6249
R1427 B.n942 B.n448 30.6249
R1428 B.n942 B.n444 30.6249
R1429 B.n948 B.n444 30.6249
R1430 B.n948 B.n440 30.6249
R1431 B.n954 B.n440 30.6249
R1432 B.n954 B.n436 30.6249
R1433 B.n960 B.n436 30.6249
R1434 B.n966 B.n432 30.6249
R1435 B.n966 B.n428 30.6249
R1436 B.n973 B.n428 30.6249
R1437 B.n973 B.n424 30.6249
R1438 B.n979 B.n424 30.6249
R1439 B.n979 B.n4 30.6249
R1440 B.n1130 B.n4 30.6249
R1441 B.n1130 B.n1129 30.6249
R1442 B.n1129 B.n1128 30.6249
R1443 B.n1128 B.n8 30.6249
R1444 B.n1122 B.n8 30.6249
R1445 B.n1122 B.n1121 30.6249
R1446 B.n1121 B.n1120 30.6249
R1447 B.n1120 B.n15 30.6249
R1448 B.n1114 B.n1113 30.6249
R1449 B.n1113 B.n1112 30.6249
R1450 B.n1112 B.n22 30.6249
R1451 B.n1106 B.n22 30.6249
R1452 B.n1106 B.n1105 30.6249
R1453 B.n1105 B.n1104 30.6249
R1454 B.n1104 B.n29 30.6249
R1455 B.n1098 B.n29 30.6249
R1456 B.n1098 B.n1097 30.6249
R1457 B.n1097 B.n1096 30.6249
R1458 B.n1096 B.n36 30.6249
R1459 B.n1090 B.n1089 30.6249
R1460 B.n1089 B.n1088 30.6249
R1461 B.n1088 B.n43 30.6249
R1462 B.n1082 B.n43 30.6249
R1463 B.n1082 B.n1081 30.6249
R1464 B.n1081 B.n1080 30.6249
R1465 B.n1080 B.n50 30.6249
R1466 B.n1074 B.n50 30.6249
R1467 B.n1074 B.n1073 30.6249
R1468 B.n1073 B.n1072 30.6249
R1469 B.n1072 B.n57 30.6249
R1470 B.n1066 B.n57 30.6249
R1471 B.n1066 B.n1065 30.6249
R1472 B.n1065 B.n1064 30.6249
R1473 B.n1058 B.n67 30.6249
R1474 B.n1058 B.n1057 30.6249
R1475 B.n1057 B.n1056 30.6249
R1476 B.n1056 B.n71 30.6249
R1477 B.n1050 B.n71 30.6249
R1478 B.n1050 B.n1049 30.6249
R1479 B.n1049 B.n1048 30.6249
R1480 B.n1048 B.n78 30.6249
R1481 B.n1042 B.n78 30.6249
R1482 B.n882 B.t5 27.022
R1483 B.n1064 B.t9 27.022
R1484 B.t3 B.n456 19.8163
R1485 B.t2 B.n36 19.8163
R1486 B.t0 B.n432 18.9155
R1487 B.t1 B.n15 18.9155
R1488 B B.n1132 18.0485
R1489 B.n960 B.t0 11.7098
R1490 B.n1114 B.t1 11.7098
R1491 B.n924 B.t3 10.8091
R1492 B.n1090 B.t2 10.8091
R1493 B.n156 B.n80 10.6151
R1494 B.n159 B.n156 10.6151
R1495 B.n160 B.n159 10.6151
R1496 B.n163 B.n160 10.6151
R1497 B.n164 B.n163 10.6151
R1498 B.n167 B.n164 10.6151
R1499 B.n168 B.n167 10.6151
R1500 B.n171 B.n168 10.6151
R1501 B.n172 B.n171 10.6151
R1502 B.n175 B.n172 10.6151
R1503 B.n176 B.n175 10.6151
R1504 B.n179 B.n176 10.6151
R1505 B.n180 B.n179 10.6151
R1506 B.n183 B.n180 10.6151
R1507 B.n184 B.n183 10.6151
R1508 B.n187 B.n184 10.6151
R1509 B.n188 B.n187 10.6151
R1510 B.n191 B.n188 10.6151
R1511 B.n192 B.n191 10.6151
R1512 B.n195 B.n192 10.6151
R1513 B.n196 B.n195 10.6151
R1514 B.n199 B.n196 10.6151
R1515 B.n200 B.n199 10.6151
R1516 B.n203 B.n200 10.6151
R1517 B.n204 B.n203 10.6151
R1518 B.n207 B.n204 10.6151
R1519 B.n208 B.n207 10.6151
R1520 B.n211 B.n208 10.6151
R1521 B.n212 B.n211 10.6151
R1522 B.n215 B.n212 10.6151
R1523 B.n216 B.n215 10.6151
R1524 B.n219 B.n216 10.6151
R1525 B.n220 B.n219 10.6151
R1526 B.n223 B.n220 10.6151
R1527 B.n224 B.n223 10.6151
R1528 B.n227 B.n224 10.6151
R1529 B.n228 B.n227 10.6151
R1530 B.n231 B.n228 10.6151
R1531 B.n232 B.n231 10.6151
R1532 B.n235 B.n232 10.6151
R1533 B.n236 B.n235 10.6151
R1534 B.n239 B.n236 10.6151
R1535 B.n240 B.n239 10.6151
R1536 B.n243 B.n240 10.6151
R1537 B.n244 B.n243 10.6151
R1538 B.n247 B.n244 10.6151
R1539 B.n248 B.n247 10.6151
R1540 B.n251 B.n248 10.6151
R1541 B.n252 B.n251 10.6151
R1542 B.n255 B.n252 10.6151
R1543 B.n256 B.n255 10.6151
R1544 B.n259 B.n256 10.6151
R1545 B.n260 B.n259 10.6151
R1546 B.n263 B.n260 10.6151
R1547 B.n264 B.n263 10.6151
R1548 B.n267 B.n264 10.6151
R1549 B.n268 B.n267 10.6151
R1550 B.n271 B.n268 10.6151
R1551 B.n272 B.n271 10.6151
R1552 B.n275 B.n272 10.6151
R1553 B.n276 B.n275 10.6151
R1554 B.n279 B.n276 10.6151
R1555 B.n284 B.n281 10.6151
R1556 B.n285 B.n284 10.6151
R1557 B.n288 B.n285 10.6151
R1558 B.n289 B.n288 10.6151
R1559 B.n292 B.n289 10.6151
R1560 B.n293 B.n292 10.6151
R1561 B.n296 B.n293 10.6151
R1562 B.n297 B.n296 10.6151
R1563 B.n301 B.n300 10.6151
R1564 B.n304 B.n301 10.6151
R1565 B.n305 B.n304 10.6151
R1566 B.n308 B.n305 10.6151
R1567 B.n309 B.n308 10.6151
R1568 B.n312 B.n309 10.6151
R1569 B.n313 B.n312 10.6151
R1570 B.n316 B.n313 10.6151
R1571 B.n317 B.n316 10.6151
R1572 B.n320 B.n317 10.6151
R1573 B.n321 B.n320 10.6151
R1574 B.n324 B.n321 10.6151
R1575 B.n325 B.n324 10.6151
R1576 B.n328 B.n325 10.6151
R1577 B.n329 B.n328 10.6151
R1578 B.n332 B.n329 10.6151
R1579 B.n333 B.n332 10.6151
R1580 B.n336 B.n333 10.6151
R1581 B.n337 B.n336 10.6151
R1582 B.n340 B.n337 10.6151
R1583 B.n341 B.n340 10.6151
R1584 B.n344 B.n341 10.6151
R1585 B.n345 B.n344 10.6151
R1586 B.n348 B.n345 10.6151
R1587 B.n349 B.n348 10.6151
R1588 B.n352 B.n349 10.6151
R1589 B.n353 B.n352 10.6151
R1590 B.n356 B.n353 10.6151
R1591 B.n357 B.n356 10.6151
R1592 B.n360 B.n357 10.6151
R1593 B.n361 B.n360 10.6151
R1594 B.n364 B.n361 10.6151
R1595 B.n365 B.n364 10.6151
R1596 B.n368 B.n365 10.6151
R1597 B.n369 B.n368 10.6151
R1598 B.n372 B.n369 10.6151
R1599 B.n373 B.n372 10.6151
R1600 B.n376 B.n373 10.6151
R1601 B.n377 B.n376 10.6151
R1602 B.n380 B.n377 10.6151
R1603 B.n381 B.n380 10.6151
R1604 B.n384 B.n381 10.6151
R1605 B.n385 B.n384 10.6151
R1606 B.n388 B.n385 10.6151
R1607 B.n389 B.n388 10.6151
R1608 B.n392 B.n389 10.6151
R1609 B.n393 B.n392 10.6151
R1610 B.n396 B.n393 10.6151
R1611 B.n397 B.n396 10.6151
R1612 B.n400 B.n397 10.6151
R1613 B.n401 B.n400 10.6151
R1614 B.n404 B.n401 10.6151
R1615 B.n405 B.n404 10.6151
R1616 B.n408 B.n405 10.6151
R1617 B.n409 B.n408 10.6151
R1618 B.n412 B.n409 10.6151
R1619 B.n413 B.n412 10.6151
R1620 B.n416 B.n413 10.6151
R1621 B.n417 B.n416 10.6151
R1622 B.n420 B.n417 10.6151
R1623 B.n421 B.n420 10.6151
R1624 B.n1039 B.n421 10.6151
R1625 B.n849 B.n501 10.6151
R1626 B.n859 B.n501 10.6151
R1627 B.n860 B.n859 10.6151
R1628 B.n861 B.n860 10.6151
R1629 B.n861 B.n493 10.6151
R1630 B.n871 B.n493 10.6151
R1631 B.n872 B.n871 10.6151
R1632 B.n873 B.n872 10.6151
R1633 B.n873 B.n486 10.6151
R1634 B.n884 B.n486 10.6151
R1635 B.n885 B.n884 10.6151
R1636 B.n886 B.n885 10.6151
R1637 B.n886 B.n478 10.6151
R1638 B.n896 B.n478 10.6151
R1639 B.n897 B.n896 10.6151
R1640 B.n898 B.n897 10.6151
R1641 B.n898 B.n470 10.6151
R1642 B.n908 B.n470 10.6151
R1643 B.n909 B.n908 10.6151
R1644 B.n910 B.n909 10.6151
R1645 B.n910 B.n462 10.6151
R1646 B.n920 B.n462 10.6151
R1647 B.n921 B.n920 10.6151
R1648 B.n922 B.n921 10.6151
R1649 B.n922 B.n454 10.6151
R1650 B.n932 B.n454 10.6151
R1651 B.n933 B.n932 10.6151
R1652 B.n934 B.n933 10.6151
R1653 B.n934 B.n446 10.6151
R1654 B.n944 B.n446 10.6151
R1655 B.n945 B.n944 10.6151
R1656 B.n946 B.n945 10.6151
R1657 B.n946 B.n438 10.6151
R1658 B.n956 B.n438 10.6151
R1659 B.n957 B.n956 10.6151
R1660 B.n958 B.n957 10.6151
R1661 B.n958 B.n430 10.6151
R1662 B.n968 B.n430 10.6151
R1663 B.n969 B.n968 10.6151
R1664 B.n971 B.n969 10.6151
R1665 B.n971 B.n970 10.6151
R1666 B.n970 B.n422 10.6151
R1667 B.n982 B.n422 10.6151
R1668 B.n983 B.n982 10.6151
R1669 B.n984 B.n983 10.6151
R1670 B.n985 B.n984 10.6151
R1671 B.n987 B.n985 10.6151
R1672 B.n988 B.n987 10.6151
R1673 B.n989 B.n988 10.6151
R1674 B.n990 B.n989 10.6151
R1675 B.n992 B.n990 10.6151
R1676 B.n993 B.n992 10.6151
R1677 B.n994 B.n993 10.6151
R1678 B.n995 B.n994 10.6151
R1679 B.n997 B.n995 10.6151
R1680 B.n998 B.n997 10.6151
R1681 B.n999 B.n998 10.6151
R1682 B.n1000 B.n999 10.6151
R1683 B.n1002 B.n1000 10.6151
R1684 B.n1003 B.n1002 10.6151
R1685 B.n1004 B.n1003 10.6151
R1686 B.n1005 B.n1004 10.6151
R1687 B.n1007 B.n1005 10.6151
R1688 B.n1008 B.n1007 10.6151
R1689 B.n1009 B.n1008 10.6151
R1690 B.n1010 B.n1009 10.6151
R1691 B.n1012 B.n1010 10.6151
R1692 B.n1013 B.n1012 10.6151
R1693 B.n1014 B.n1013 10.6151
R1694 B.n1015 B.n1014 10.6151
R1695 B.n1017 B.n1015 10.6151
R1696 B.n1018 B.n1017 10.6151
R1697 B.n1019 B.n1018 10.6151
R1698 B.n1020 B.n1019 10.6151
R1699 B.n1022 B.n1020 10.6151
R1700 B.n1023 B.n1022 10.6151
R1701 B.n1024 B.n1023 10.6151
R1702 B.n1025 B.n1024 10.6151
R1703 B.n1027 B.n1025 10.6151
R1704 B.n1028 B.n1027 10.6151
R1705 B.n1029 B.n1028 10.6151
R1706 B.n1030 B.n1029 10.6151
R1707 B.n1032 B.n1030 10.6151
R1708 B.n1033 B.n1032 10.6151
R1709 B.n1034 B.n1033 10.6151
R1710 B.n1035 B.n1034 10.6151
R1711 B.n1037 B.n1035 10.6151
R1712 B.n1038 B.n1037 10.6151
R1713 B.n579 B.n505 10.6151
R1714 B.n580 B.n579 10.6151
R1715 B.n581 B.n580 10.6151
R1716 B.n581 B.n575 10.6151
R1717 B.n587 B.n575 10.6151
R1718 B.n588 B.n587 10.6151
R1719 B.n589 B.n588 10.6151
R1720 B.n589 B.n573 10.6151
R1721 B.n595 B.n573 10.6151
R1722 B.n596 B.n595 10.6151
R1723 B.n597 B.n596 10.6151
R1724 B.n597 B.n571 10.6151
R1725 B.n603 B.n571 10.6151
R1726 B.n604 B.n603 10.6151
R1727 B.n605 B.n604 10.6151
R1728 B.n605 B.n569 10.6151
R1729 B.n611 B.n569 10.6151
R1730 B.n612 B.n611 10.6151
R1731 B.n613 B.n612 10.6151
R1732 B.n613 B.n567 10.6151
R1733 B.n619 B.n567 10.6151
R1734 B.n620 B.n619 10.6151
R1735 B.n621 B.n620 10.6151
R1736 B.n621 B.n565 10.6151
R1737 B.n627 B.n565 10.6151
R1738 B.n628 B.n627 10.6151
R1739 B.n629 B.n628 10.6151
R1740 B.n629 B.n563 10.6151
R1741 B.n635 B.n563 10.6151
R1742 B.n636 B.n635 10.6151
R1743 B.n637 B.n636 10.6151
R1744 B.n637 B.n561 10.6151
R1745 B.n643 B.n561 10.6151
R1746 B.n644 B.n643 10.6151
R1747 B.n645 B.n644 10.6151
R1748 B.n645 B.n559 10.6151
R1749 B.n651 B.n559 10.6151
R1750 B.n652 B.n651 10.6151
R1751 B.n653 B.n652 10.6151
R1752 B.n653 B.n557 10.6151
R1753 B.n659 B.n557 10.6151
R1754 B.n660 B.n659 10.6151
R1755 B.n661 B.n660 10.6151
R1756 B.n661 B.n555 10.6151
R1757 B.n667 B.n555 10.6151
R1758 B.n668 B.n667 10.6151
R1759 B.n669 B.n668 10.6151
R1760 B.n669 B.n553 10.6151
R1761 B.n675 B.n553 10.6151
R1762 B.n676 B.n675 10.6151
R1763 B.n677 B.n676 10.6151
R1764 B.n677 B.n551 10.6151
R1765 B.n683 B.n551 10.6151
R1766 B.n684 B.n683 10.6151
R1767 B.n685 B.n684 10.6151
R1768 B.n685 B.n549 10.6151
R1769 B.n691 B.n549 10.6151
R1770 B.n692 B.n691 10.6151
R1771 B.n693 B.n692 10.6151
R1772 B.n693 B.n547 10.6151
R1773 B.n699 B.n547 10.6151
R1774 B.n700 B.n699 10.6151
R1775 B.n702 B.n543 10.6151
R1776 B.n708 B.n543 10.6151
R1777 B.n709 B.n708 10.6151
R1778 B.n710 B.n709 10.6151
R1779 B.n710 B.n541 10.6151
R1780 B.n716 B.n541 10.6151
R1781 B.n717 B.n716 10.6151
R1782 B.n721 B.n717 10.6151
R1783 B.n727 B.n539 10.6151
R1784 B.n728 B.n727 10.6151
R1785 B.n729 B.n728 10.6151
R1786 B.n729 B.n537 10.6151
R1787 B.n735 B.n537 10.6151
R1788 B.n736 B.n735 10.6151
R1789 B.n737 B.n736 10.6151
R1790 B.n737 B.n535 10.6151
R1791 B.n743 B.n535 10.6151
R1792 B.n744 B.n743 10.6151
R1793 B.n745 B.n744 10.6151
R1794 B.n745 B.n533 10.6151
R1795 B.n751 B.n533 10.6151
R1796 B.n752 B.n751 10.6151
R1797 B.n753 B.n752 10.6151
R1798 B.n753 B.n531 10.6151
R1799 B.n759 B.n531 10.6151
R1800 B.n760 B.n759 10.6151
R1801 B.n761 B.n760 10.6151
R1802 B.n761 B.n529 10.6151
R1803 B.n767 B.n529 10.6151
R1804 B.n768 B.n767 10.6151
R1805 B.n769 B.n768 10.6151
R1806 B.n769 B.n527 10.6151
R1807 B.n775 B.n527 10.6151
R1808 B.n776 B.n775 10.6151
R1809 B.n777 B.n776 10.6151
R1810 B.n777 B.n525 10.6151
R1811 B.n783 B.n525 10.6151
R1812 B.n784 B.n783 10.6151
R1813 B.n785 B.n784 10.6151
R1814 B.n785 B.n523 10.6151
R1815 B.n791 B.n523 10.6151
R1816 B.n792 B.n791 10.6151
R1817 B.n793 B.n792 10.6151
R1818 B.n793 B.n521 10.6151
R1819 B.n799 B.n521 10.6151
R1820 B.n800 B.n799 10.6151
R1821 B.n801 B.n800 10.6151
R1822 B.n801 B.n519 10.6151
R1823 B.n807 B.n519 10.6151
R1824 B.n808 B.n807 10.6151
R1825 B.n809 B.n808 10.6151
R1826 B.n809 B.n517 10.6151
R1827 B.n815 B.n517 10.6151
R1828 B.n816 B.n815 10.6151
R1829 B.n817 B.n816 10.6151
R1830 B.n817 B.n515 10.6151
R1831 B.n823 B.n515 10.6151
R1832 B.n824 B.n823 10.6151
R1833 B.n825 B.n824 10.6151
R1834 B.n825 B.n513 10.6151
R1835 B.n831 B.n513 10.6151
R1836 B.n832 B.n831 10.6151
R1837 B.n833 B.n832 10.6151
R1838 B.n833 B.n511 10.6151
R1839 B.n839 B.n511 10.6151
R1840 B.n840 B.n839 10.6151
R1841 B.n841 B.n840 10.6151
R1842 B.n841 B.n509 10.6151
R1843 B.n847 B.n509 10.6151
R1844 B.n848 B.n847 10.6151
R1845 B.n854 B.n853 10.6151
R1846 B.n855 B.n854 10.6151
R1847 B.n855 B.n497 10.6151
R1848 B.n865 B.n497 10.6151
R1849 B.n866 B.n865 10.6151
R1850 B.n867 B.n866 10.6151
R1851 B.n867 B.n489 10.6151
R1852 B.n878 B.n489 10.6151
R1853 B.n879 B.n878 10.6151
R1854 B.n880 B.n879 10.6151
R1855 B.n880 B.n482 10.6151
R1856 B.n890 B.n482 10.6151
R1857 B.n891 B.n890 10.6151
R1858 B.n892 B.n891 10.6151
R1859 B.n892 B.n474 10.6151
R1860 B.n902 B.n474 10.6151
R1861 B.n903 B.n902 10.6151
R1862 B.n904 B.n903 10.6151
R1863 B.n904 B.n466 10.6151
R1864 B.n914 B.n466 10.6151
R1865 B.n915 B.n914 10.6151
R1866 B.n916 B.n915 10.6151
R1867 B.n916 B.n458 10.6151
R1868 B.n926 B.n458 10.6151
R1869 B.n927 B.n926 10.6151
R1870 B.n928 B.n927 10.6151
R1871 B.n928 B.n450 10.6151
R1872 B.n938 B.n450 10.6151
R1873 B.n939 B.n938 10.6151
R1874 B.n940 B.n939 10.6151
R1875 B.n940 B.n442 10.6151
R1876 B.n950 B.n442 10.6151
R1877 B.n951 B.n950 10.6151
R1878 B.n952 B.n951 10.6151
R1879 B.n952 B.n434 10.6151
R1880 B.n962 B.n434 10.6151
R1881 B.n963 B.n962 10.6151
R1882 B.n964 B.n963 10.6151
R1883 B.n964 B.n426 10.6151
R1884 B.n975 B.n426 10.6151
R1885 B.n976 B.n975 10.6151
R1886 B.n977 B.n976 10.6151
R1887 B.n977 B.n0 10.6151
R1888 B.n1126 B.n1 10.6151
R1889 B.n1126 B.n1125 10.6151
R1890 B.n1125 B.n1124 10.6151
R1891 B.n1124 B.n10 10.6151
R1892 B.n1118 B.n10 10.6151
R1893 B.n1118 B.n1117 10.6151
R1894 B.n1117 B.n1116 10.6151
R1895 B.n1116 B.n17 10.6151
R1896 B.n1110 B.n17 10.6151
R1897 B.n1110 B.n1109 10.6151
R1898 B.n1109 B.n1108 10.6151
R1899 B.n1108 B.n24 10.6151
R1900 B.n1102 B.n24 10.6151
R1901 B.n1102 B.n1101 10.6151
R1902 B.n1101 B.n1100 10.6151
R1903 B.n1100 B.n31 10.6151
R1904 B.n1094 B.n31 10.6151
R1905 B.n1094 B.n1093 10.6151
R1906 B.n1093 B.n1092 10.6151
R1907 B.n1092 B.n38 10.6151
R1908 B.n1086 B.n38 10.6151
R1909 B.n1086 B.n1085 10.6151
R1910 B.n1085 B.n1084 10.6151
R1911 B.n1084 B.n45 10.6151
R1912 B.n1078 B.n45 10.6151
R1913 B.n1078 B.n1077 10.6151
R1914 B.n1077 B.n1076 10.6151
R1915 B.n1076 B.n52 10.6151
R1916 B.n1070 B.n52 10.6151
R1917 B.n1070 B.n1069 10.6151
R1918 B.n1069 B.n1068 10.6151
R1919 B.n1068 B.n59 10.6151
R1920 B.n1062 B.n59 10.6151
R1921 B.n1062 B.n1061 10.6151
R1922 B.n1061 B.n1060 10.6151
R1923 B.n1060 B.n65 10.6151
R1924 B.n1054 B.n65 10.6151
R1925 B.n1054 B.n1053 10.6151
R1926 B.n1053 B.n1052 10.6151
R1927 B.n1052 B.n73 10.6151
R1928 B.n1046 B.n73 10.6151
R1929 B.n1046 B.n1045 10.6151
R1930 B.n1045 B.n1044 10.6151
R1931 B.n281 B.n280 6.5566
R1932 B.n297 B.n153 6.5566
R1933 B.n702 B.n701 6.5566
R1934 B.n721 B.n720 6.5566
R1935 B.n280 B.n279 4.05904
R1936 B.n300 B.n153 4.05904
R1937 B.n701 B.n700 4.05904
R1938 B.n720 B.n539 4.05904
R1939 B.n875 B.t5 3.60337
R1940 B.n67 B.t9 3.60337
R1941 B.n1132 B.n0 2.81026
R1942 B.n1132 B.n1 2.81026
R1943 VP.n21 VP.n20 161.3
R1944 VP.n19 VP.n1 161.3
R1945 VP.n18 VP.n17 161.3
R1946 VP.n16 VP.n2 161.3
R1947 VP.n15 VP.n14 161.3
R1948 VP.n13 VP.n3 161.3
R1949 VP.n12 VP.n11 161.3
R1950 VP.n10 VP.n4 161.3
R1951 VP.n9 VP.n8 161.3
R1952 VP.n5 VP.t2 156.429
R1953 VP.n5 VP.t0 155.089
R1954 VP.n7 VP.t3 122.743
R1955 VP.n0 VP.t1 122.743
R1956 VP.n7 VP.n6 87.8654
R1957 VP.n22 VP.n0 87.8654
R1958 VP.n6 VP.n5 57.1968
R1959 VP.n14 VP.n13 40.4934
R1960 VP.n14 VP.n2 40.4934
R1961 VP.n8 VP.n4 24.4675
R1962 VP.n12 VP.n4 24.4675
R1963 VP.n13 VP.n12 24.4675
R1964 VP.n18 VP.n2 24.4675
R1965 VP.n19 VP.n18 24.4675
R1966 VP.n20 VP.n19 24.4675
R1967 VP.n8 VP.n7 2.20253
R1968 VP.n20 VP.n0 2.20253
R1969 VP.n9 VP.n6 0.354971
R1970 VP.n22 VP.n21 0.354971
R1971 VP VP.n22 0.26696
R1972 VP.n10 VP.n9 0.189894
R1973 VP.n11 VP.n10 0.189894
R1974 VP.n11 VP.n3 0.189894
R1975 VP.n15 VP.n3 0.189894
R1976 VP.n16 VP.n15 0.189894
R1977 VP.n17 VP.n16 0.189894
R1978 VP.n17 VP.n1 0.189894
R1979 VP.n21 VP.n1 0.189894
R1980 VDD1 VDD1.n1 115.21
R1981 VDD1 VDD1.n0 63.9424
R1982 VDD1.n0 VDD1.t1 1.03444
R1983 VDD1.n0 VDD1.t3 1.03444
R1984 VDD1.n1 VDD1.t0 1.03444
R1985 VDD1.n1 VDD1.t2 1.03444
C0 VDD2 VP 0.467972f
C1 VDD2 VTAIL 7.28849f
C2 VDD2 VDD1 1.30724f
C3 VP VN 8.352849f
C4 VN VTAIL 7.56603f
C5 VDD1 VN 0.149902f
C6 VP VTAIL 7.58013f
C7 VP VDD1 8.146441f
C8 VDD1 VTAIL 7.22651f
C9 VDD2 VN 7.8294f
C10 VDD2 B 4.973081f
C11 VDD1 B 10.22117f
C12 VTAIL B 15.063789f
C13 VN B 13.50509f
C14 VP B 11.887332f
C15 VDD1.t1 B 0.406092f
C16 VDD1.t3 B 0.406092f
C17 VDD1.n0 B 3.71867f
C18 VDD1.t0 B 0.406092f
C19 VDD1.t2 B 0.406092f
C20 VDD1.n1 B 4.73669f
C21 VP.t1 B 3.75175f
C22 VP.n0 B 1.35979f
C23 VP.n1 B 0.018922f
C24 VP.n2 B 0.037607f
C25 VP.n3 B 0.018922f
C26 VP.n4 B 0.035265f
C27 VP.t2 B 4.06302f
C28 VP.t0 B 4.05113f
C29 VP.n5 B 3.88775f
C30 VP.n6 B 1.31506f
C31 VP.t3 B 3.75175f
C32 VP.n7 B 1.35979f
C33 VP.n8 B 0.019421f
C34 VP.n9 B 0.030539f
C35 VP.n10 B 0.018922f
C36 VP.n11 B 0.018922f
C37 VP.n12 B 0.035265f
C38 VP.n13 B 0.037607f
C39 VP.n14 B 0.015297f
C40 VP.n15 B 0.018922f
C41 VP.n16 B 0.018922f
C42 VP.n17 B 0.018922f
C43 VP.n18 B 0.035265f
C44 VP.n19 B 0.035265f
C45 VP.n20 B 0.019421f
C46 VP.n21 B 0.030539f
C47 VP.n22 B 0.058078f
C48 VDD2.t2 B 0.403397f
C49 VDD2.t3 B 0.403397f
C50 VDD2.n0 B 4.67653f
C51 VDD2.t1 B 0.403397f
C52 VDD2.t0 B 0.403397f
C53 VDD2.n1 B 3.69351f
C54 VDD2.n2 B 4.80779f
C55 VTAIL.t5 B 2.71217f
C56 VTAIL.n0 B 0.315974f
C57 VTAIL.t0 B 2.71217f
C58 VTAIL.n1 B 0.40179f
C59 VTAIL.t3 B 2.71217f
C60 VTAIL.n2 B 1.59888f
C61 VTAIL.t6 B 2.71218f
C62 VTAIL.n3 B 1.59886f
C63 VTAIL.t7 B 2.71218f
C64 VTAIL.n4 B 0.401771f
C65 VTAIL.t1 B 2.71218f
C66 VTAIL.n5 B 0.401771f
C67 VTAIL.t2 B 2.71217f
C68 VTAIL.n6 B 1.59888f
C69 VTAIL.t4 B 2.71217f
C70 VTAIL.n7 B 1.50721f
C71 VN.t0 B 3.99629f
C72 VN.t1 B 4.00802f
C73 VN.n0 B 2.45468f
C74 VN.t2 B 3.99629f
C75 VN.t3 B 4.00802f
C76 VN.n1 B 3.8424f
.ends

