* NGSPICE file created from diff_pair_sample_1413.ext - technology: sky130A

.subckt diff_pair_sample_1413 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.36
X1 B.t8 B.t6 B.t7 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.36
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=4.4889 ps=23.8 w=11.51 l=1.36
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=4.4889 ps=23.8 w=11.51 l=1.36
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=4.4889 ps=23.8 w=11.51 l=1.36
X5 B.t5 B.t3 B.t4 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.36
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=4.4889 ps=23.8 w=11.51 l=1.36
X7 B.t2 B.t0 B.t1 w_n1646_n3270# sky130_fd_pr__pfet_01v8 ad=4.4889 pd=23.8 as=0 ps=0 w=11.51 l=1.36
R0 B.n355 B.n60 585
R1 B.n357 B.n356 585
R2 B.n358 B.n59 585
R3 B.n360 B.n359 585
R4 B.n361 B.n58 585
R5 B.n363 B.n362 585
R6 B.n364 B.n57 585
R7 B.n366 B.n365 585
R8 B.n367 B.n56 585
R9 B.n369 B.n368 585
R10 B.n370 B.n55 585
R11 B.n372 B.n371 585
R12 B.n373 B.n54 585
R13 B.n375 B.n374 585
R14 B.n376 B.n53 585
R15 B.n378 B.n377 585
R16 B.n379 B.n52 585
R17 B.n381 B.n380 585
R18 B.n382 B.n51 585
R19 B.n384 B.n383 585
R20 B.n385 B.n50 585
R21 B.n387 B.n386 585
R22 B.n388 B.n49 585
R23 B.n390 B.n389 585
R24 B.n391 B.n48 585
R25 B.n393 B.n392 585
R26 B.n394 B.n47 585
R27 B.n396 B.n395 585
R28 B.n397 B.n46 585
R29 B.n399 B.n398 585
R30 B.n400 B.n45 585
R31 B.n402 B.n401 585
R32 B.n403 B.n44 585
R33 B.n405 B.n404 585
R34 B.n406 B.n43 585
R35 B.n408 B.n407 585
R36 B.n409 B.n42 585
R37 B.n411 B.n410 585
R38 B.n412 B.n41 585
R39 B.n414 B.n413 585
R40 B.n416 B.n415 585
R41 B.n417 B.n37 585
R42 B.n419 B.n418 585
R43 B.n420 B.n36 585
R44 B.n422 B.n421 585
R45 B.n423 B.n35 585
R46 B.n425 B.n424 585
R47 B.n426 B.n34 585
R48 B.n428 B.n427 585
R49 B.n429 B.n31 585
R50 B.n432 B.n431 585
R51 B.n433 B.n30 585
R52 B.n435 B.n434 585
R53 B.n436 B.n29 585
R54 B.n438 B.n437 585
R55 B.n439 B.n28 585
R56 B.n441 B.n440 585
R57 B.n442 B.n27 585
R58 B.n444 B.n443 585
R59 B.n445 B.n26 585
R60 B.n447 B.n446 585
R61 B.n448 B.n25 585
R62 B.n450 B.n449 585
R63 B.n451 B.n24 585
R64 B.n453 B.n452 585
R65 B.n454 B.n23 585
R66 B.n456 B.n455 585
R67 B.n457 B.n22 585
R68 B.n459 B.n458 585
R69 B.n460 B.n21 585
R70 B.n462 B.n461 585
R71 B.n463 B.n20 585
R72 B.n465 B.n464 585
R73 B.n466 B.n19 585
R74 B.n468 B.n467 585
R75 B.n469 B.n18 585
R76 B.n471 B.n470 585
R77 B.n472 B.n17 585
R78 B.n474 B.n473 585
R79 B.n475 B.n16 585
R80 B.n477 B.n476 585
R81 B.n478 B.n15 585
R82 B.n480 B.n479 585
R83 B.n481 B.n14 585
R84 B.n483 B.n482 585
R85 B.n484 B.n13 585
R86 B.n486 B.n485 585
R87 B.n487 B.n12 585
R88 B.n489 B.n488 585
R89 B.n490 B.n11 585
R90 B.n354 B.n353 585
R91 B.n352 B.n61 585
R92 B.n351 B.n350 585
R93 B.n349 B.n62 585
R94 B.n348 B.n347 585
R95 B.n346 B.n63 585
R96 B.n345 B.n344 585
R97 B.n343 B.n64 585
R98 B.n342 B.n341 585
R99 B.n340 B.n65 585
R100 B.n339 B.n338 585
R101 B.n337 B.n66 585
R102 B.n336 B.n335 585
R103 B.n334 B.n67 585
R104 B.n333 B.n332 585
R105 B.n331 B.n68 585
R106 B.n330 B.n329 585
R107 B.n328 B.n69 585
R108 B.n327 B.n326 585
R109 B.n325 B.n70 585
R110 B.n324 B.n323 585
R111 B.n322 B.n71 585
R112 B.n321 B.n320 585
R113 B.n319 B.n72 585
R114 B.n318 B.n317 585
R115 B.n316 B.n73 585
R116 B.n315 B.n314 585
R117 B.n313 B.n74 585
R118 B.n312 B.n311 585
R119 B.n310 B.n75 585
R120 B.n309 B.n308 585
R121 B.n307 B.n76 585
R122 B.n306 B.n305 585
R123 B.n304 B.n77 585
R124 B.n303 B.n302 585
R125 B.n301 B.n78 585
R126 B.n300 B.n299 585
R127 B.n163 B.n128 585
R128 B.n165 B.n164 585
R129 B.n166 B.n127 585
R130 B.n168 B.n167 585
R131 B.n169 B.n126 585
R132 B.n171 B.n170 585
R133 B.n172 B.n125 585
R134 B.n174 B.n173 585
R135 B.n175 B.n124 585
R136 B.n177 B.n176 585
R137 B.n178 B.n123 585
R138 B.n180 B.n179 585
R139 B.n181 B.n122 585
R140 B.n183 B.n182 585
R141 B.n184 B.n121 585
R142 B.n186 B.n185 585
R143 B.n187 B.n120 585
R144 B.n189 B.n188 585
R145 B.n190 B.n119 585
R146 B.n192 B.n191 585
R147 B.n193 B.n118 585
R148 B.n195 B.n194 585
R149 B.n196 B.n117 585
R150 B.n198 B.n197 585
R151 B.n199 B.n116 585
R152 B.n201 B.n200 585
R153 B.n202 B.n115 585
R154 B.n204 B.n203 585
R155 B.n205 B.n114 585
R156 B.n207 B.n206 585
R157 B.n208 B.n113 585
R158 B.n210 B.n209 585
R159 B.n211 B.n112 585
R160 B.n213 B.n212 585
R161 B.n214 B.n111 585
R162 B.n216 B.n215 585
R163 B.n217 B.n110 585
R164 B.n219 B.n218 585
R165 B.n220 B.n109 585
R166 B.n222 B.n221 585
R167 B.n224 B.n223 585
R168 B.n225 B.n105 585
R169 B.n227 B.n226 585
R170 B.n228 B.n104 585
R171 B.n230 B.n229 585
R172 B.n231 B.n103 585
R173 B.n233 B.n232 585
R174 B.n234 B.n102 585
R175 B.n236 B.n235 585
R176 B.n237 B.n99 585
R177 B.n240 B.n239 585
R178 B.n241 B.n98 585
R179 B.n243 B.n242 585
R180 B.n244 B.n97 585
R181 B.n246 B.n245 585
R182 B.n247 B.n96 585
R183 B.n249 B.n248 585
R184 B.n250 B.n95 585
R185 B.n252 B.n251 585
R186 B.n253 B.n94 585
R187 B.n255 B.n254 585
R188 B.n256 B.n93 585
R189 B.n258 B.n257 585
R190 B.n259 B.n92 585
R191 B.n261 B.n260 585
R192 B.n262 B.n91 585
R193 B.n264 B.n263 585
R194 B.n265 B.n90 585
R195 B.n267 B.n266 585
R196 B.n268 B.n89 585
R197 B.n270 B.n269 585
R198 B.n271 B.n88 585
R199 B.n273 B.n272 585
R200 B.n274 B.n87 585
R201 B.n276 B.n275 585
R202 B.n277 B.n86 585
R203 B.n279 B.n278 585
R204 B.n280 B.n85 585
R205 B.n282 B.n281 585
R206 B.n283 B.n84 585
R207 B.n285 B.n284 585
R208 B.n286 B.n83 585
R209 B.n288 B.n287 585
R210 B.n289 B.n82 585
R211 B.n291 B.n290 585
R212 B.n292 B.n81 585
R213 B.n294 B.n293 585
R214 B.n295 B.n80 585
R215 B.n297 B.n296 585
R216 B.n298 B.n79 585
R217 B.n162 B.n161 585
R218 B.n160 B.n129 585
R219 B.n159 B.n158 585
R220 B.n157 B.n130 585
R221 B.n156 B.n155 585
R222 B.n154 B.n131 585
R223 B.n153 B.n152 585
R224 B.n151 B.n132 585
R225 B.n150 B.n149 585
R226 B.n148 B.n133 585
R227 B.n147 B.n146 585
R228 B.n145 B.n134 585
R229 B.n144 B.n143 585
R230 B.n142 B.n135 585
R231 B.n141 B.n140 585
R232 B.n139 B.n136 585
R233 B.n138 B.n137 585
R234 B.n2 B.n0 585
R235 B.n517 B.n1 585
R236 B.n516 B.n515 585
R237 B.n514 B.n3 585
R238 B.n513 B.n512 585
R239 B.n511 B.n4 585
R240 B.n510 B.n509 585
R241 B.n508 B.n5 585
R242 B.n507 B.n506 585
R243 B.n505 B.n6 585
R244 B.n504 B.n503 585
R245 B.n502 B.n7 585
R246 B.n501 B.n500 585
R247 B.n499 B.n8 585
R248 B.n498 B.n497 585
R249 B.n496 B.n9 585
R250 B.n495 B.n494 585
R251 B.n493 B.n10 585
R252 B.n492 B.n491 585
R253 B.n519 B.n518 585
R254 B.n163 B.n162 502.111
R255 B.n492 B.n11 502.111
R256 B.n300 B.n79 502.111
R257 B.n355 B.n354 502.111
R258 B.n100 B.t9 408.841
R259 B.n106 B.t3 408.841
R260 B.n32 B.t0 408.841
R261 B.n38 B.t6 408.841
R262 B.n100 B.t11 399.745
R263 B.n38 B.t7 399.745
R264 B.n106 B.t5 399.745
R265 B.n32 B.t1 399.745
R266 B.n101 B.t10 366.969
R267 B.n39 B.t8 366.969
R268 B.n107 B.t4 366.969
R269 B.n33 B.t2 366.969
R270 B.n162 B.n129 163.367
R271 B.n158 B.n129 163.367
R272 B.n158 B.n157 163.367
R273 B.n157 B.n156 163.367
R274 B.n156 B.n131 163.367
R275 B.n152 B.n131 163.367
R276 B.n152 B.n151 163.367
R277 B.n151 B.n150 163.367
R278 B.n150 B.n133 163.367
R279 B.n146 B.n133 163.367
R280 B.n146 B.n145 163.367
R281 B.n145 B.n144 163.367
R282 B.n144 B.n135 163.367
R283 B.n140 B.n135 163.367
R284 B.n140 B.n139 163.367
R285 B.n139 B.n138 163.367
R286 B.n138 B.n2 163.367
R287 B.n518 B.n2 163.367
R288 B.n518 B.n517 163.367
R289 B.n517 B.n516 163.367
R290 B.n516 B.n3 163.367
R291 B.n512 B.n3 163.367
R292 B.n512 B.n511 163.367
R293 B.n511 B.n510 163.367
R294 B.n510 B.n5 163.367
R295 B.n506 B.n5 163.367
R296 B.n506 B.n505 163.367
R297 B.n505 B.n504 163.367
R298 B.n504 B.n7 163.367
R299 B.n500 B.n7 163.367
R300 B.n500 B.n499 163.367
R301 B.n499 B.n498 163.367
R302 B.n498 B.n9 163.367
R303 B.n494 B.n9 163.367
R304 B.n494 B.n493 163.367
R305 B.n493 B.n492 163.367
R306 B.n164 B.n163 163.367
R307 B.n164 B.n127 163.367
R308 B.n168 B.n127 163.367
R309 B.n169 B.n168 163.367
R310 B.n170 B.n169 163.367
R311 B.n170 B.n125 163.367
R312 B.n174 B.n125 163.367
R313 B.n175 B.n174 163.367
R314 B.n176 B.n175 163.367
R315 B.n176 B.n123 163.367
R316 B.n180 B.n123 163.367
R317 B.n181 B.n180 163.367
R318 B.n182 B.n181 163.367
R319 B.n182 B.n121 163.367
R320 B.n186 B.n121 163.367
R321 B.n187 B.n186 163.367
R322 B.n188 B.n187 163.367
R323 B.n188 B.n119 163.367
R324 B.n192 B.n119 163.367
R325 B.n193 B.n192 163.367
R326 B.n194 B.n193 163.367
R327 B.n194 B.n117 163.367
R328 B.n198 B.n117 163.367
R329 B.n199 B.n198 163.367
R330 B.n200 B.n199 163.367
R331 B.n200 B.n115 163.367
R332 B.n204 B.n115 163.367
R333 B.n205 B.n204 163.367
R334 B.n206 B.n205 163.367
R335 B.n206 B.n113 163.367
R336 B.n210 B.n113 163.367
R337 B.n211 B.n210 163.367
R338 B.n212 B.n211 163.367
R339 B.n212 B.n111 163.367
R340 B.n216 B.n111 163.367
R341 B.n217 B.n216 163.367
R342 B.n218 B.n217 163.367
R343 B.n218 B.n109 163.367
R344 B.n222 B.n109 163.367
R345 B.n223 B.n222 163.367
R346 B.n223 B.n105 163.367
R347 B.n227 B.n105 163.367
R348 B.n228 B.n227 163.367
R349 B.n229 B.n228 163.367
R350 B.n229 B.n103 163.367
R351 B.n233 B.n103 163.367
R352 B.n234 B.n233 163.367
R353 B.n235 B.n234 163.367
R354 B.n235 B.n99 163.367
R355 B.n240 B.n99 163.367
R356 B.n241 B.n240 163.367
R357 B.n242 B.n241 163.367
R358 B.n242 B.n97 163.367
R359 B.n246 B.n97 163.367
R360 B.n247 B.n246 163.367
R361 B.n248 B.n247 163.367
R362 B.n248 B.n95 163.367
R363 B.n252 B.n95 163.367
R364 B.n253 B.n252 163.367
R365 B.n254 B.n253 163.367
R366 B.n254 B.n93 163.367
R367 B.n258 B.n93 163.367
R368 B.n259 B.n258 163.367
R369 B.n260 B.n259 163.367
R370 B.n260 B.n91 163.367
R371 B.n264 B.n91 163.367
R372 B.n265 B.n264 163.367
R373 B.n266 B.n265 163.367
R374 B.n266 B.n89 163.367
R375 B.n270 B.n89 163.367
R376 B.n271 B.n270 163.367
R377 B.n272 B.n271 163.367
R378 B.n272 B.n87 163.367
R379 B.n276 B.n87 163.367
R380 B.n277 B.n276 163.367
R381 B.n278 B.n277 163.367
R382 B.n278 B.n85 163.367
R383 B.n282 B.n85 163.367
R384 B.n283 B.n282 163.367
R385 B.n284 B.n283 163.367
R386 B.n284 B.n83 163.367
R387 B.n288 B.n83 163.367
R388 B.n289 B.n288 163.367
R389 B.n290 B.n289 163.367
R390 B.n290 B.n81 163.367
R391 B.n294 B.n81 163.367
R392 B.n295 B.n294 163.367
R393 B.n296 B.n295 163.367
R394 B.n296 B.n79 163.367
R395 B.n301 B.n300 163.367
R396 B.n302 B.n301 163.367
R397 B.n302 B.n77 163.367
R398 B.n306 B.n77 163.367
R399 B.n307 B.n306 163.367
R400 B.n308 B.n307 163.367
R401 B.n308 B.n75 163.367
R402 B.n312 B.n75 163.367
R403 B.n313 B.n312 163.367
R404 B.n314 B.n313 163.367
R405 B.n314 B.n73 163.367
R406 B.n318 B.n73 163.367
R407 B.n319 B.n318 163.367
R408 B.n320 B.n319 163.367
R409 B.n320 B.n71 163.367
R410 B.n324 B.n71 163.367
R411 B.n325 B.n324 163.367
R412 B.n326 B.n325 163.367
R413 B.n326 B.n69 163.367
R414 B.n330 B.n69 163.367
R415 B.n331 B.n330 163.367
R416 B.n332 B.n331 163.367
R417 B.n332 B.n67 163.367
R418 B.n336 B.n67 163.367
R419 B.n337 B.n336 163.367
R420 B.n338 B.n337 163.367
R421 B.n338 B.n65 163.367
R422 B.n342 B.n65 163.367
R423 B.n343 B.n342 163.367
R424 B.n344 B.n343 163.367
R425 B.n344 B.n63 163.367
R426 B.n348 B.n63 163.367
R427 B.n349 B.n348 163.367
R428 B.n350 B.n349 163.367
R429 B.n350 B.n61 163.367
R430 B.n354 B.n61 163.367
R431 B.n488 B.n11 163.367
R432 B.n488 B.n487 163.367
R433 B.n487 B.n486 163.367
R434 B.n486 B.n13 163.367
R435 B.n482 B.n13 163.367
R436 B.n482 B.n481 163.367
R437 B.n481 B.n480 163.367
R438 B.n480 B.n15 163.367
R439 B.n476 B.n15 163.367
R440 B.n476 B.n475 163.367
R441 B.n475 B.n474 163.367
R442 B.n474 B.n17 163.367
R443 B.n470 B.n17 163.367
R444 B.n470 B.n469 163.367
R445 B.n469 B.n468 163.367
R446 B.n468 B.n19 163.367
R447 B.n464 B.n19 163.367
R448 B.n464 B.n463 163.367
R449 B.n463 B.n462 163.367
R450 B.n462 B.n21 163.367
R451 B.n458 B.n21 163.367
R452 B.n458 B.n457 163.367
R453 B.n457 B.n456 163.367
R454 B.n456 B.n23 163.367
R455 B.n452 B.n23 163.367
R456 B.n452 B.n451 163.367
R457 B.n451 B.n450 163.367
R458 B.n450 B.n25 163.367
R459 B.n446 B.n25 163.367
R460 B.n446 B.n445 163.367
R461 B.n445 B.n444 163.367
R462 B.n444 B.n27 163.367
R463 B.n440 B.n27 163.367
R464 B.n440 B.n439 163.367
R465 B.n439 B.n438 163.367
R466 B.n438 B.n29 163.367
R467 B.n434 B.n29 163.367
R468 B.n434 B.n433 163.367
R469 B.n433 B.n432 163.367
R470 B.n432 B.n31 163.367
R471 B.n427 B.n31 163.367
R472 B.n427 B.n426 163.367
R473 B.n426 B.n425 163.367
R474 B.n425 B.n35 163.367
R475 B.n421 B.n35 163.367
R476 B.n421 B.n420 163.367
R477 B.n420 B.n419 163.367
R478 B.n419 B.n37 163.367
R479 B.n415 B.n37 163.367
R480 B.n415 B.n414 163.367
R481 B.n414 B.n41 163.367
R482 B.n410 B.n41 163.367
R483 B.n410 B.n409 163.367
R484 B.n409 B.n408 163.367
R485 B.n408 B.n43 163.367
R486 B.n404 B.n43 163.367
R487 B.n404 B.n403 163.367
R488 B.n403 B.n402 163.367
R489 B.n402 B.n45 163.367
R490 B.n398 B.n45 163.367
R491 B.n398 B.n397 163.367
R492 B.n397 B.n396 163.367
R493 B.n396 B.n47 163.367
R494 B.n392 B.n47 163.367
R495 B.n392 B.n391 163.367
R496 B.n391 B.n390 163.367
R497 B.n390 B.n49 163.367
R498 B.n386 B.n49 163.367
R499 B.n386 B.n385 163.367
R500 B.n385 B.n384 163.367
R501 B.n384 B.n51 163.367
R502 B.n380 B.n51 163.367
R503 B.n380 B.n379 163.367
R504 B.n379 B.n378 163.367
R505 B.n378 B.n53 163.367
R506 B.n374 B.n53 163.367
R507 B.n374 B.n373 163.367
R508 B.n373 B.n372 163.367
R509 B.n372 B.n55 163.367
R510 B.n368 B.n55 163.367
R511 B.n368 B.n367 163.367
R512 B.n367 B.n366 163.367
R513 B.n366 B.n57 163.367
R514 B.n362 B.n57 163.367
R515 B.n362 B.n361 163.367
R516 B.n361 B.n360 163.367
R517 B.n360 B.n59 163.367
R518 B.n356 B.n59 163.367
R519 B.n356 B.n355 163.367
R520 B.n238 B.n101 59.5399
R521 B.n108 B.n107 59.5399
R522 B.n430 B.n33 59.5399
R523 B.n40 B.n39 59.5399
R524 B.n101 B.n100 32.7763
R525 B.n107 B.n106 32.7763
R526 B.n33 B.n32 32.7763
R527 B.n39 B.n38 32.7763
R528 B.n491 B.n490 32.6249
R529 B.n353 B.n60 32.6249
R530 B.n299 B.n298 32.6249
R531 B.n161 B.n128 32.6249
R532 B B.n519 18.0485
R533 B.n490 B.n489 10.6151
R534 B.n489 B.n12 10.6151
R535 B.n485 B.n12 10.6151
R536 B.n485 B.n484 10.6151
R537 B.n484 B.n483 10.6151
R538 B.n483 B.n14 10.6151
R539 B.n479 B.n14 10.6151
R540 B.n479 B.n478 10.6151
R541 B.n478 B.n477 10.6151
R542 B.n477 B.n16 10.6151
R543 B.n473 B.n16 10.6151
R544 B.n473 B.n472 10.6151
R545 B.n472 B.n471 10.6151
R546 B.n471 B.n18 10.6151
R547 B.n467 B.n18 10.6151
R548 B.n467 B.n466 10.6151
R549 B.n466 B.n465 10.6151
R550 B.n465 B.n20 10.6151
R551 B.n461 B.n20 10.6151
R552 B.n461 B.n460 10.6151
R553 B.n460 B.n459 10.6151
R554 B.n459 B.n22 10.6151
R555 B.n455 B.n22 10.6151
R556 B.n455 B.n454 10.6151
R557 B.n454 B.n453 10.6151
R558 B.n453 B.n24 10.6151
R559 B.n449 B.n24 10.6151
R560 B.n449 B.n448 10.6151
R561 B.n448 B.n447 10.6151
R562 B.n447 B.n26 10.6151
R563 B.n443 B.n26 10.6151
R564 B.n443 B.n442 10.6151
R565 B.n442 B.n441 10.6151
R566 B.n441 B.n28 10.6151
R567 B.n437 B.n28 10.6151
R568 B.n437 B.n436 10.6151
R569 B.n436 B.n435 10.6151
R570 B.n435 B.n30 10.6151
R571 B.n431 B.n30 10.6151
R572 B.n429 B.n428 10.6151
R573 B.n428 B.n34 10.6151
R574 B.n424 B.n34 10.6151
R575 B.n424 B.n423 10.6151
R576 B.n423 B.n422 10.6151
R577 B.n422 B.n36 10.6151
R578 B.n418 B.n36 10.6151
R579 B.n418 B.n417 10.6151
R580 B.n417 B.n416 10.6151
R581 B.n413 B.n412 10.6151
R582 B.n412 B.n411 10.6151
R583 B.n411 B.n42 10.6151
R584 B.n407 B.n42 10.6151
R585 B.n407 B.n406 10.6151
R586 B.n406 B.n405 10.6151
R587 B.n405 B.n44 10.6151
R588 B.n401 B.n44 10.6151
R589 B.n401 B.n400 10.6151
R590 B.n400 B.n399 10.6151
R591 B.n399 B.n46 10.6151
R592 B.n395 B.n46 10.6151
R593 B.n395 B.n394 10.6151
R594 B.n394 B.n393 10.6151
R595 B.n393 B.n48 10.6151
R596 B.n389 B.n48 10.6151
R597 B.n389 B.n388 10.6151
R598 B.n388 B.n387 10.6151
R599 B.n387 B.n50 10.6151
R600 B.n383 B.n50 10.6151
R601 B.n383 B.n382 10.6151
R602 B.n382 B.n381 10.6151
R603 B.n381 B.n52 10.6151
R604 B.n377 B.n52 10.6151
R605 B.n377 B.n376 10.6151
R606 B.n376 B.n375 10.6151
R607 B.n375 B.n54 10.6151
R608 B.n371 B.n54 10.6151
R609 B.n371 B.n370 10.6151
R610 B.n370 B.n369 10.6151
R611 B.n369 B.n56 10.6151
R612 B.n365 B.n56 10.6151
R613 B.n365 B.n364 10.6151
R614 B.n364 B.n363 10.6151
R615 B.n363 B.n58 10.6151
R616 B.n359 B.n58 10.6151
R617 B.n359 B.n358 10.6151
R618 B.n358 B.n357 10.6151
R619 B.n357 B.n60 10.6151
R620 B.n299 B.n78 10.6151
R621 B.n303 B.n78 10.6151
R622 B.n304 B.n303 10.6151
R623 B.n305 B.n304 10.6151
R624 B.n305 B.n76 10.6151
R625 B.n309 B.n76 10.6151
R626 B.n310 B.n309 10.6151
R627 B.n311 B.n310 10.6151
R628 B.n311 B.n74 10.6151
R629 B.n315 B.n74 10.6151
R630 B.n316 B.n315 10.6151
R631 B.n317 B.n316 10.6151
R632 B.n317 B.n72 10.6151
R633 B.n321 B.n72 10.6151
R634 B.n322 B.n321 10.6151
R635 B.n323 B.n322 10.6151
R636 B.n323 B.n70 10.6151
R637 B.n327 B.n70 10.6151
R638 B.n328 B.n327 10.6151
R639 B.n329 B.n328 10.6151
R640 B.n329 B.n68 10.6151
R641 B.n333 B.n68 10.6151
R642 B.n334 B.n333 10.6151
R643 B.n335 B.n334 10.6151
R644 B.n335 B.n66 10.6151
R645 B.n339 B.n66 10.6151
R646 B.n340 B.n339 10.6151
R647 B.n341 B.n340 10.6151
R648 B.n341 B.n64 10.6151
R649 B.n345 B.n64 10.6151
R650 B.n346 B.n345 10.6151
R651 B.n347 B.n346 10.6151
R652 B.n347 B.n62 10.6151
R653 B.n351 B.n62 10.6151
R654 B.n352 B.n351 10.6151
R655 B.n353 B.n352 10.6151
R656 B.n165 B.n128 10.6151
R657 B.n166 B.n165 10.6151
R658 B.n167 B.n166 10.6151
R659 B.n167 B.n126 10.6151
R660 B.n171 B.n126 10.6151
R661 B.n172 B.n171 10.6151
R662 B.n173 B.n172 10.6151
R663 B.n173 B.n124 10.6151
R664 B.n177 B.n124 10.6151
R665 B.n178 B.n177 10.6151
R666 B.n179 B.n178 10.6151
R667 B.n179 B.n122 10.6151
R668 B.n183 B.n122 10.6151
R669 B.n184 B.n183 10.6151
R670 B.n185 B.n184 10.6151
R671 B.n185 B.n120 10.6151
R672 B.n189 B.n120 10.6151
R673 B.n190 B.n189 10.6151
R674 B.n191 B.n190 10.6151
R675 B.n191 B.n118 10.6151
R676 B.n195 B.n118 10.6151
R677 B.n196 B.n195 10.6151
R678 B.n197 B.n196 10.6151
R679 B.n197 B.n116 10.6151
R680 B.n201 B.n116 10.6151
R681 B.n202 B.n201 10.6151
R682 B.n203 B.n202 10.6151
R683 B.n203 B.n114 10.6151
R684 B.n207 B.n114 10.6151
R685 B.n208 B.n207 10.6151
R686 B.n209 B.n208 10.6151
R687 B.n209 B.n112 10.6151
R688 B.n213 B.n112 10.6151
R689 B.n214 B.n213 10.6151
R690 B.n215 B.n214 10.6151
R691 B.n215 B.n110 10.6151
R692 B.n219 B.n110 10.6151
R693 B.n220 B.n219 10.6151
R694 B.n221 B.n220 10.6151
R695 B.n225 B.n224 10.6151
R696 B.n226 B.n225 10.6151
R697 B.n226 B.n104 10.6151
R698 B.n230 B.n104 10.6151
R699 B.n231 B.n230 10.6151
R700 B.n232 B.n231 10.6151
R701 B.n232 B.n102 10.6151
R702 B.n236 B.n102 10.6151
R703 B.n237 B.n236 10.6151
R704 B.n239 B.n98 10.6151
R705 B.n243 B.n98 10.6151
R706 B.n244 B.n243 10.6151
R707 B.n245 B.n244 10.6151
R708 B.n245 B.n96 10.6151
R709 B.n249 B.n96 10.6151
R710 B.n250 B.n249 10.6151
R711 B.n251 B.n250 10.6151
R712 B.n251 B.n94 10.6151
R713 B.n255 B.n94 10.6151
R714 B.n256 B.n255 10.6151
R715 B.n257 B.n256 10.6151
R716 B.n257 B.n92 10.6151
R717 B.n261 B.n92 10.6151
R718 B.n262 B.n261 10.6151
R719 B.n263 B.n262 10.6151
R720 B.n263 B.n90 10.6151
R721 B.n267 B.n90 10.6151
R722 B.n268 B.n267 10.6151
R723 B.n269 B.n268 10.6151
R724 B.n269 B.n88 10.6151
R725 B.n273 B.n88 10.6151
R726 B.n274 B.n273 10.6151
R727 B.n275 B.n274 10.6151
R728 B.n275 B.n86 10.6151
R729 B.n279 B.n86 10.6151
R730 B.n280 B.n279 10.6151
R731 B.n281 B.n280 10.6151
R732 B.n281 B.n84 10.6151
R733 B.n285 B.n84 10.6151
R734 B.n286 B.n285 10.6151
R735 B.n287 B.n286 10.6151
R736 B.n287 B.n82 10.6151
R737 B.n291 B.n82 10.6151
R738 B.n292 B.n291 10.6151
R739 B.n293 B.n292 10.6151
R740 B.n293 B.n80 10.6151
R741 B.n297 B.n80 10.6151
R742 B.n298 B.n297 10.6151
R743 B.n161 B.n160 10.6151
R744 B.n160 B.n159 10.6151
R745 B.n159 B.n130 10.6151
R746 B.n155 B.n130 10.6151
R747 B.n155 B.n154 10.6151
R748 B.n154 B.n153 10.6151
R749 B.n153 B.n132 10.6151
R750 B.n149 B.n132 10.6151
R751 B.n149 B.n148 10.6151
R752 B.n148 B.n147 10.6151
R753 B.n147 B.n134 10.6151
R754 B.n143 B.n134 10.6151
R755 B.n143 B.n142 10.6151
R756 B.n142 B.n141 10.6151
R757 B.n141 B.n136 10.6151
R758 B.n137 B.n136 10.6151
R759 B.n137 B.n0 10.6151
R760 B.n515 B.n1 10.6151
R761 B.n515 B.n514 10.6151
R762 B.n514 B.n513 10.6151
R763 B.n513 B.n4 10.6151
R764 B.n509 B.n4 10.6151
R765 B.n509 B.n508 10.6151
R766 B.n508 B.n507 10.6151
R767 B.n507 B.n6 10.6151
R768 B.n503 B.n6 10.6151
R769 B.n503 B.n502 10.6151
R770 B.n502 B.n501 10.6151
R771 B.n501 B.n8 10.6151
R772 B.n497 B.n8 10.6151
R773 B.n497 B.n496 10.6151
R774 B.n496 B.n495 10.6151
R775 B.n495 B.n10 10.6151
R776 B.n491 B.n10 10.6151
R777 B.n431 B.n430 9.36635
R778 B.n413 B.n40 9.36635
R779 B.n221 B.n108 9.36635
R780 B.n239 B.n238 9.36635
R781 B.n519 B.n0 2.81026
R782 B.n519 B.n1 2.81026
R783 B.n430 B.n429 1.24928
R784 B.n416 B.n40 1.24928
R785 B.n224 B.n108 1.24928
R786 B.n238 B.n237 1.24928
R787 VN VN.t0 354.913
R788 VN VN.t1 313.776
R789 VTAIL.n242 VTAIL.n186 756.745
R790 VTAIL.n56 VTAIL.n0 756.745
R791 VTAIL.n180 VTAIL.n124 756.745
R792 VTAIL.n118 VTAIL.n62 756.745
R793 VTAIL.n207 VTAIL.n206 585
R794 VTAIL.n209 VTAIL.n208 585
R795 VTAIL.n202 VTAIL.n201 585
R796 VTAIL.n215 VTAIL.n214 585
R797 VTAIL.n217 VTAIL.n216 585
R798 VTAIL.n198 VTAIL.n197 585
R799 VTAIL.n224 VTAIL.n223 585
R800 VTAIL.n225 VTAIL.n196 585
R801 VTAIL.n227 VTAIL.n226 585
R802 VTAIL.n194 VTAIL.n193 585
R803 VTAIL.n233 VTAIL.n232 585
R804 VTAIL.n235 VTAIL.n234 585
R805 VTAIL.n190 VTAIL.n189 585
R806 VTAIL.n241 VTAIL.n240 585
R807 VTAIL.n243 VTAIL.n242 585
R808 VTAIL.n21 VTAIL.n20 585
R809 VTAIL.n23 VTAIL.n22 585
R810 VTAIL.n16 VTAIL.n15 585
R811 VTAIL.n29 VTAIL.n28 585
R812 VTAIL.n31 VTAIL.n30 585
R813 VTAIL.n12 VTAIL.n11 585
R814 VTAIL.n38 VTAIL.n37 585
R815 VTAIL.n39 VTAIL.n10 585
R816 VTAIL.n41 VTAIL.n40 585
R817 VTAIL.n8 VTAIL.n7 585
R818 VTAIL.n47 VTAIL.n46 585
R819 VTAIL.n49 VTAIL.n48 585
R820 VTAIL.n4 VTAIL.n3 585
R821 VTAIL.n55 VTAIL.n54 585
R822 VTAIL.n57 VTAIL.n56 585
R823 VTAIL.n181 VTAIL.n180 585
R824 VTAIL.n179 VTAIL.n178 585
R825 VTAIL.n128 VTAIL.n127 585
R826 VTAIL.n173 VTAIL.n172 585
R827 VTAIL.n171 VTAIL.n170 585
R828 VTAIL.n132 VTAIL.n131 585
R829 VTAIL.n136 VTAIL.n134 585
R830 VTAIL.n165 VTAIL.n164 585
R831 VTAIL.n163 VTAIL.n162 585
R832 VTAIL.n138 VTAIL.n137 585
R833 VTAIL.n157 VTAIL.n156 585
R834 VTAIL.n155 VTAIL.n154 585
R835 VTAIL.n142 VTAIL.n141 585
R836 VTAIL.n149 VTAIL.n148 585
R837 VTAIL.n147 VTAIL.n146 585
R838 VTAIL.n119 VTAIL.n118 585
R839 VTAIL.n117 VTAIL.n116 585
R840 VTAIL.n66 VTAIL.n65 585
R841 VTAIL.n111 VTAIL.n110 585
R842 VTAIL.n109 VTAIL.n108 585
R843 VTAIL.n70 VTAIL.n69 585
R844 VTAIL.n74 VTAIL.n72 585
R845 VTAIL.n103 VTAIL.n102 585
R846 VTAIL.n101 VTAIL.n100 585
R847 VTAIL.n76 VTAIL.n75 585
R848 VTAIL.n95 VTAIL.n94 585
R849 VTAIL.n93 VTAIL.n92 585
R850 VTAIL.n80 VTAIL.n79 585
R851 VTAIL.n87 VTAIL.n86 585
R852 VTAIL.n85 VTAIL.n84 585
R853 VTAIL.n205 VTAIL.t2 329.036
R854 VTAIL.n19 VTAIL.t1 329.036
R855 VTAIL.n145 VTAIL.t0 329.036
R856 VTAIL.n83 VTAIL.t3 329.036
R857 VTAIL.n208 VTAIL.n207 171.744
R858 VTAIL.n208 VTAIL.n201 171.744
R859 VTAIL.n215 VTAIL.n201 171.744
R860 VTAIL.n216 VTAIL.n215 171.744
R861 VTAIL.n216 VTAIL.n197 171.744
R862 VTAIL.n224 VTAIL.n197 171.744
R863 VTAIL.n225 VTAIL.n224 171.744
R864 VTAIL.n226 VTAIL.n225 171.744
R865 VTAIL.n226 VTAIL.n193 171.744
R866 VTAIL.n233 VTAIL.n193 171.744
R867 VTAIL.n234 VTAIL.n233 171.744
R868 VTAIL.n234 VTAIL.n189 171.744
R869 VTAIL.n241 VTAIL.n189 171.744
R870 VTAIL.n242 VTAIL.n241 171.744
R871 VTAIL.n22 VTAIL.n21 171.744
R872 VTAIL.n22 VTAIL.n15 171.744
R873 VTAIL.n29 VTAIL.n15 171.744
R874 VTAIL.n30 VTAIL.n29 171.744
R875 VTAIL.n30 VTAIL.n11 171.744
R876 VTAIL.n38 VTAIL.n11 171.744
R877 VTAIL.n39 VTAIL.n38 171.744
R878 VTAIL.n40 VTAIL.n39 171.744
R879 VTAIL.n40 VTAIL.n7 171.744
R880 VTAIL.n47 VTAIL.n7 171.744
R881 VTAIL.n48 VTAIL.n47 171.744
R882 VTAIL.n48 VTAIL.n3 171.744
R883 VTAIL.n55 VTAIL.n3 171.744
R884 VTAIL.n56 VTAIL.n55 171.744
R885 VTAIL.n180 VTAIL.n179 171.744
R886 VTAIL.n179 VTAIL.n127 171.744
R887 VTAIL.n172 VTAIL.n127 171.744
R888 VTAIL.n172 VTAIL.n171 171.744
R889 VTAIL.n171 VTAIL.n131 171.744
R890 VTAIL.n136 VTAIL.n131 171.744
R891 VTAIL.n164 VTAIL.n136 171.744
R892 VTAIL.n164 VTAIL.n163 171.744
R893 VTAIL.n163 VTAIL.n137 171.744
R894 VTAIL.n156 VTAIL.n137 171.744
R895 VTAIL.n156 VTAIL.n155 171.744
R896 VTAIL.n155 VTAIL.n141 171.744
R897 VTAIL.n148 VTAIL.n141 171.744
R898 VTAIL.n148 VTAIL.n147 171.744
R899 VTAIL.n118 VTAIL.n117 171.744
R900 VTAIL.n117 VTAIL.n65 171.744
R901 VTAIL.n110 VTAIL.n65 171.744
R902 VTAIL.n110 VTAIL.n109 171.744
R903 VTAIL.n109 VTAIL.n69 171.744
R904 VTAIL.n74 VTAIL.n69 171.744
R905 VTAIL.n102 VTAIL.n74 171.744
R906 VTAIL.n102 VTAIL.n101 171.744
R907 VTAIL.n101 VTAIL.n75 171.744
R908 VTAIL.n94 VTAIL.n75 171.744
R909 VTAIL.n94 VTAIL.n93 171.744
R910 VTAIL.n93 VTAIL.n79 171.744
R911 VTAIL.n86 VTAIL.n79 171.744
R912 VTAIL.n86 VTAIL.n85 171.744
R913 VTAIL.n207 VTAIL.t2 85.8723
R914 VTAIL.n21 VTAIL.t1 85.8723
R915 VTAIL.n147 VTAIL.t0 85.8723
R916 VTAIL.n85 VTAIL.t3 85.8723
R917 VTAIL.n247 VTAIL.n246 34.3187
R918 VTAIL.n61 VTAIL.n60 34.3187
R919 VTAIL.n185 VTAIL.n184 34.3187
R920 VTAIL.n123 VTAIL.n122 34.3187
R921 VTAIL.n123 VTAIL.n61 25.2031
R922 VTAIL.n247 VTAIL.n185 23.7462
R923 VTAIL.n227 VTAIL.n194 13.1884
R924 VTAIL.n41 VTAIL.n8 13.1884
R925 VTAIL.n134 VTAIL.n132 13.1884
R926 VTAIL.n72 VTAIL.n70 13.1884
R927 VTAIL.n228 VTAIL.n196 12.8005
R928 VTAIL.n232 VTAIL.n231 12.8005
R929 VTAIL.n42 VTAIL.n10 12.8005
R930 VTAIL.n46 VTAIL.n45 12.8005
R931 VTAIL.n170 VTAIL.n169 12.8005
R932 VTAIL.n166 VTAIL.n165 12.8005
R933 VTAIL.n108 VTAIL.n107 12.8005
R934 VTAIL.n104 VTAIL.n103 12.8005
R935 VTAIL.n223 VTAIL.n222 12.0247
R936 VTAIL.n235 VTAIL.n192 12.0247
R937 VTAIL.n37 VTAIL.n36 12.0247
R938 VTAIL.n49 VTAIL.n6 12.0247
R939 VTAIL.n173 VTAIL.n130 12.0247
R940 VTAIL.n162 VTAIL.n135 12.0247
R941 VTAIL.n111 VTAIL.n68 12.0247
R942 VTAIL.n100 VTAIL.n73 12.0247
R943 VTAIL.n221 VTAIL.n198 11.249
R944 VTAIL.n236 VTAIL.n190 11.249
R945 VTAIL.n35 VTAIL.n12 11.249
R946 VTAIL.n50 VTAIL.n4 11.249
R947 VTAIL.n174 VTAIL.n128 11.249
R948 VTAIL.n161 VTAIL.n138 11.249
R949 VTAIL.n112 VTAIL.n66 11.249
R950 VTAIL.n99 VTAIL.n76 11.249
R951 VTAIL.n206 VTAIL.n205 10.7239
R952 VTAIL.n20 VTAIL.n19 10.7239
R953 VTAIL.n146 VTAIL.n145 10.7239
R954 VTAIL.n84 VTAIL.n83 10.7239
R955 VTAIL.n218 VTAIL.n217 10.4732
R956 VTAIL.n240 VTAIL.n239 10.4732
R957 VTAIL.n32 VTAIL.n31 10.4732
R958 VTAIL.n54 VTAIL.n53 10.4732
R959 VTAIL.n178 VTAIL.n177 10.4732
R960 VTAIL.n158 VTAIL.n157 10.4732
R961 VTAIL.n116 VTAIL.n115 10.4732
R962 VTAIL.n96 VTAIL.n95 10.4732
R963 VTAIL.n214 VTAIL.n200 9.69747
R964 VTAIL.n243 VTAIL.n188 9.69747
R965 VTAIL.n28 VTAIL.n14 9.69747
R966 VTAIL.n57 VTAIL.n2 9.69747
R967 VTAIL.n181 VTAIL.n126 9.69747
R968 VTAIL.n154 VTAIL.n140 9.69747
R969 VTAIL.n119 VTAIL.n64 9.69747
R970 VTAIL.n92 VTAIL.n78 9.69747
R971 VTAIL.n246 VTAIL.n245 9.45567
R972 VTAIL.n60 VTAIL.n59 9.45567
R973 VTAIL.n184 VTAIL.n183 9.45567
R974 VTAIL.n122 VTAIL.n121 9.45567
R975 VTAIL.n245 VTAIL.n244 9.3005
R976 VTAIL.n188 VTAIL.n187 9.3005
R977 VTAIL.n239 VTAIL.n238 9.3005
R978 VTAIL.n237 VTAIL.n236 9.3005
R979 VTAIL.n192 VTAIL.n191 9.3005
R980 VTAIL.n231 VTAIL.n230 9.3005
R981 VTAIL.n204 VTAIL.n203 9.3005
R982 VTAIL.n211 VTAIL.n210 9.3005
R983 VTAIL.n213 VTAIL.n212 9.3005
R984 VTAIL.n200 VTAIL.n199 9.3005
R985 VTAIL.n219 VTAIL.n218 9.3005
R986 VTAIL.n221 VTAIL.n220 9.3005
R987 VTAIL.n222 VTAIL.n195 9.3005
R988 VTAIL.n229 VTAIL.n228 9.3005
R989 VTAIL.n59 VTAIL.n58 9.3005
R990 VTAIL.n2 VTAIL.n1 9.3005
R991 VTAIL.n53 VTAIL.n52 9.3005
R992 VTAIL.n51 VTAIL.n50 9.3005
R993 VTAIL.n6 VTAIL.n5 9.3005
R994 VTAIL.n45 VTAIL.n44 9.3005
R995 VTAIL.n18 VTAIL.n17 9.3005
R996 VTAIL.n25 VTAIL.n24 9.3005
R997 VTAIL.n27 VTAIL.n26 9.3005
R998 VTAIL.n14 VTAIL.n13 9.3005
R999 VTAIL.n33 VTAIL.n32 9.3005
R1000 VTAIL.n35 VTAIL.n34 9.3005
R1001 VTAIL.n36 VTAIL.n9 9.3005
R1002 VTAIL.n43 VTAIL.n42 9.3005
R1003 VTAIL.n144 VTAIL.n143 9.3005
R1004 VTAIL.n151 VTAIL.n150 9.3005
R1005 VTAIL.n153 VTAIL.n152 9.3005
R1006 VTAIL.n140 VTAIL.n139 9.3005
R1007 VTAIL.n159 VTAIL.n158 9.3005
R1008 VTAIL.n161 VTAIL.n160 9.3005
R1009 VTAIL.n135 VTAIL.n133 9.3005
R1010 VTAIL.n167 VTAIL.n166 9.3005
R1011 VTAIL.n183 VTAIL.n182 9.3005
R1012 VTAIL.n126 VTAIL.n125 9.3005
R1013 VTAIL.n177 VTAIL.n176 9.3005
R1014 VTAIL.n175 VTAIL.n174 9.3005
R1015 VTAIL.n130 VTAIL.n129 9.3005
R1016 VTAIL.n169 VTAIL.n168 9.3005
R1017 VTAIL.n82 VTAIL.n81 9.3005
R1018 VTAIL.n89 VTAIL.n88 9.3005
R1019 VTAIL.n91 VTAIL.n90 9.3005
R1020 VTAIL.n78 VTAIL.n77 9.3005
R1021 VTAIL.n97 VTAIL.n96 9.3005
R1022 VTAIL.n99 VTAIL.n98 9.3005
R1023 VTAIL.n73 VTAIL.n71 9.3005
R1024 VTAIL.n105 VTAIL.n104 9.3005
R1025 VTAIL.n121 VTAIL.n120 9.3005
R1026 VTAIL.n64 VTAIL.n63 9.3005
R1027 VTAIL.n115 VTAIL.n114 9.3005
R1028 VTAIL.n113 VTAIL.n112 9.3005
R1029 VTAIL.n68 VTAIL.n67 9.3005
R1030 VTAIL.n107 VTAIL.n106 9.3005
R1031 VTAIL.n213 VTAIL.n202 8.92171
R1032 VTAIL.n244 VTAIL.n186 8.92171
R1033 VTAIL.n27 VTAIL.n16 8.92171
R1034 VTAIL.n58 VTAIL.n0 8.92171
R1035 VTAIL.n182 VTAIL.n124 8.92171
R1036 VTAIL.n153 VTAIL.n142 8.92171
R1037 VTAIL.n120 VTAIL.n62 8.92171
R1038 VTAIL.n91 VTAIL.n80 8.92171
R1039 VTAIL.n210 VTAIL.n209 8.14595
R1040 VTAIL.n24 VTAIL.n23 8.14595
R1041 VTAIL.n150 VTAIL.n149 8.14595
R1042 VTAIL.n88 VTAIL.n87 8.14595
R1043 VTAIL.n206 VTAIL.n204 7.3702
R1044 VTAIL.n20 VTAIL.n18 7.3702
R1045 VTAIL.n146 VTAIL.n144 7.3702
R1046 VTAIL.n84 VTAIL.n82 7.3702
R1047 VTAIL.n209 VTAIL.n204 5.81868
R1048 VTAIL.n23 VTAIL.n18 5.81868
R1049 VTAIL.n149 VTAIL.n144 5.81868
R1050 VTAIL.n87 VTAIL.n82 5.81868
R1051 VTAIL.n210 VTAIL.n202 5.04292
R1052 VTAIL.n246 VTAIL.n186 5.04292
R1053 VTAIL.n24 VTAIL.n16 5.04292
R1054 VTAIL.n60 VTAIL.n0 5.04292
R1055 VTAIL.n184 VTAIL.n124 5.04292
R1056 VTAIL.n150 VTAIL.n142 5.04292
R1057 VTAIL.n122 VTAIL.n62 5.04292
R1058 VTAIL.n88 VTAIL.n80 5.04292
R1059 VTAIL.n214 VTAIL.n213 4.26717
R1060 VTAIL.n244 VTAIL.n243 4.26717
R1061 VTAIL.n28 VTAIL.n27 4.26717
R1062 VTAIL.n58 VTAIL.n57 4.26717
R1063 VTAIL.n182 VTAIL.n181 4.26717
R1064 VTAIL.n154 VTAIL.n153 4.26717
R1065 VTAIL.n120 VTAIL.n119 4.26717
R1066 VTAIL.n92 VTAIL.n91 4.26717
R1067 VTAIL.n217 VTAIL.n200 3.49141
R1068 VTAIL.n240 VTAIL.n188 3.49141
R1069 VTAIL.n31 VTAIL.n14 3.49141
R1070 VTAIL.n54 VTAIL.n2 3.49141
R1071 VTAIL.n178 VTAIL.n126 3.49141
R1072 VTAIL.n157 VTAIL.n140 3.49141
R1073 VTAIL.n116 VTAIL.n64 3.49141
R1074 VTAIL.n95 VTAIL.n78 3.49141
R1075 VTAIL.n218 VTAIL.n198 2.71565
R1076 VTAIL.n239 VTAIL.n190 2.71565
R1077 VTAIL.n32 VTAIL.n12 2.71565
R1078 VTAIL.n53 VTAIL.n4 2.71565
R1079 VTAIL.n177 VTAIL.n128 2.71565
R1080 VTAIL.n158 VTAIL.n138 2.71565
R1081 VTAIL.n115 VTAIL.n66 2.71565
R1082 VTAIL.n96 VTAIL.n76 2.71565
R1083 VTAIL.n205 VTAIL.n203 2.41282
R1084 VTAIL.n19 VTAIL.n17 2.41282
R1085 VTAIL.n145 VTAIL.n143 2.41282
R1086 VTAIL.n83 VTAIL.n81 2.41282
R1087 VTAIL.n223 VTAIL.n221 1.93989
R1088 VTAIL.n236 VTAIL.n235 1.93989
R1089 VTAIL.n37 VTAIL.n35 1.93989
R1090 VTAIL.n50 VTAIL.n49 1.93989
R1091 VTAIL.n174 VTAIL.n173 1.93989
R1092 VTAIL.n162 VTAIL.n161 1.93989
R1093 VTAIL.n112 VTAIL.n111 1.93989
R1094 VTAIL.n100 VTAIL.n99 1.93989
R1095 VTAIL.n185 VTAIL.n123 1.19878
R1096 VTAIL.n222 VTAIL.n196 1.16414
R1097 VTAIL.n232 VTAIL.n192 1.16414
R1098 VTAIL.n36 VTAIL.n10 1.16414
R1099 VTAIL.n46 VTAIL.n6 1.16414
R1100 VTAIL.n170 VTAIL.n130 1.16414
R1101 VTAIL.n165 VTAIL.n135 1.16414
R1102 VTAIL.n108 VTAIL.n68 1.16414
R1103 VTAIL.n103 VTAIL.n73 1.16414
R1104 VTAIL VTAIL.n61 0.892741
R1105 VTAIL.n228 VTAIL.n227 0.388379
R1106 VTAIL.n231 VTAIL.n194 0.388379
R1107 VTAIL.n42 VTAIL.n41 0.388379
R1108 VTAIL.n45 VTAIL.n8 0.388379
R1109 VTAIL.n169 VTAIL.n132 0.388379
R1110 VTAIL.n166 VTAIL.n134 0.388379
R1111 VTAIL.n107 VTAIL.n70 0.388379
R1112 VTAIL.n104 VTAIL.n72 0.388379
R1113 VTAIL VTAIL.n247 0.306534
R1114 VTAIL.n211 VTAIL.n203 0.155672
R1115 VTAIL.n212 VTAIL.n211 0.155672
R1116 VTAIL.n212 VTAIL.n199 0.155672
R1117 VTAIL.n219 VTAIL.n199 0.155672
R1118 VTAIL.n220 VTAIL.n219 0.155672
R1119 VTAIL.n220 VTAIL.n195 0.155672
R1120 VTAIL.n229 VTAIL.n195 0.155672
R1121 VTAIL.n230 VTAIL.n229 0.155672
R1122 VTAIL.n230 VTAIL.n191 0.155672
R1123 VTAIL.n237 VTAIL.n191 0.155672
R1124 VTAIL.n238 VTAIL.n237 0.155672
R1125 VTAIL.n238 VTAIL.n187 0.155672
R1126 VTAIL.n245 VTAIL.n187 0.155672
R1127 VTAIL.n25 VTAIL.n17 0.155672
R1128 VTAIL.n26 VTAIL.n25 0.155672
R1129 VTAIL.n26 VTAIL.n13 0.155672
R1130 VTAIL.n33 VTAIL.n13 0.155672
R1131 VTAIL.n34 VTAIL.n33 0.155672
R1132 VTAIL.n34 VTAIL.n9 0.155672
R1133 VTAIL.n43 VTAIL.n9 0.155672
R1134 VTAIL.n44 VTAIL.n43 0.155672
R1135 VTAIL.n44 VTAIL.n5 0.155672
R1136 VTAIL.n51 VTAIL.n5 0.155672
R1137 VTAIL.n52 VTAIL.n51 0.155672
R1138 VTAIL.n52 VTAIL.n1 0.155672
R1139 VTAIL.n59 VTAIL.n1 0.155672
R1140 VTAIL.n183 VTAIL.n125 0.155672
R1141 VTAIL.n176 VTAIL.n125 0.155672
R1142 VTAIL.n176 VTAIL.n175 0.155672
R1143 VTAIL.n175 VTAIL.n129 0.155672
R1144 VTAIL.n168 VTAIL.n129 0.155672
R1145 VTAIL.n168 VTAIL.n167 0.155672
R1146 VTAIL.n167 VTAIL.n133 0.155672
R1147 VTAIL.n160 VTAIL.n133 0.155672
R1148 VTAIL.n160 VTAIL.n159 0.155672
R1149 VTAIL.n159 VTAIL.n139 0.155672
R1150 VTAIL.n152 VTAIL.n139 0.155672
R1151 VTAIL.n152 VTAIL.n151 0.155672
R1152 VTAIL.n151 VTAIL.n143 0.155672
R1153 VTAIL.n121 VTAIL.n63 0.155672
R1154 VTAIL.n114 VTAIL.n63 0.155672
R1155 VTAIL.n114 VTAIL.n113 0.155672
R1156 VTAIL.n113 VTAIL.n67 0.155672
R1157 VTAIL.n106 VTAIL.n67 0.155672
R1158 VTAIL.n106 VTAIL.n105 0.155672
R1159 VTAIL.n105 VTAIL.n71 0.155672
R1160 VTAIL.n98 VTAIL.n71 0.155672
R1161 VTAIL.n98 VTAIL.n97 0.155672
R1162 VTAIL.n97 VTAIL.n77 0.155672
R1163 VTAIL.n90 VTAIL.n77 0.155672
R1164 VTAIL.n90 VTAIL.n89 0.155672
R1165 VTAIL.n89 VTAIL.n81 0.155672
R1166 VDD2.n117 VDD2.n61 756.745
R1167 VDD2.n56 VDD2.n0 756.745
R1168 VDD2.n118 VDD2.n117 585
R1169 VDD2.n116 VDD2.n115 585
R1170 VDD2.n65 VDD2.n64 585
R1171 VDD2.n110 VDD2.n109 585
R1172 VDD2.n108 VDD2.n107 585
R1173 VDD2.n69 VDD2.n68 585
R1174 VDD2.n73 VDD2.n71 585
R1175 VDD2.n102 VDD2.n101 585
R1176 VDD2.n100 VDD2.n99 585
R1177 VDD2.n75 VDD2.n74 585
R1178 VDD2.n94 VDD2.n93 585
R1179 VDD2.n92 VDD2.n91 585
R1180 VDD2.n79 VDD2.n78 585
R1181 VDD2.n86 VDD2.n85 585
R1182 VDD2.n84 VDD2.n83 585
R1183 VDD2.n21 VDD2.n20 585
R1184 VDD2.n23 VDD2.n22 585
R1185 VDD2.n16 VDD2.n15 585
R1186 VDD2.n29 VDD2.n28 585
R1187 VDD2.n31 VDD2.n30 585
R1188 VDD2.n12 VDD2.n11 585
R1189 VDD2.n38 VDD2.n37 585
R1190 VDD2.n39 VDD2.n10 585
R1191 VDD2.n41 VDD2.n40 585
R1192 VDD2.n8 VDD2.n7 585
R1193 VDD2.n47 VDD2.n46 585
R1194 VDD2.n49 VDD2.n48 585
R1195 VDD2.n4 VDD2.n3 585
R1196 VDD2.n55 VDD2.n54 585
R1197 VDD2.n57 VDD2.n56 585
R1198 VDD2.n82 VDD2.t1 329.036
R1199 VDD2.n19 VDD2.t0 329.036
R1200 VDD2.n117 VDD2.n116 171.744
R1201 VDD2.n116 VDD2.n64 171.744
R1202 VDD2.n109 VDD2.n64 171.744
R1203 VDD2.n109 VDD2.n108 171.744
R1204 VDD2.n108 VDD2.n68 171.744
R1205 VDD2.n73 VDD2.n68 171.744
R1206 VDD2.n101 VDD2.n73 171.744
R1207 VDD2.n101 VDD2.n100 171.744
R1208 VDD2.n100 VDD2.n74 171.744
R1209 VDD2.n93 VDD2.n74 171.744
R1210 VDD2.n93 VDD2.n92 171.744
R1211 VDD2.n92 VDD2.n78 171.744
R1212 VDD2.n85 VDD2.n78 171.744
R1213 VDD2.n85 VDD2.n84 171.744
R1214 VDD2.n22 VDD2.n21 171.744
R1215 VDD2.n22 VDD2.n15 171.744
R1216 VDD2.n29 VDD2.n15 171.744
R1217 VDD2.n30 VDD2.n29 171.744
R1218 VDD2.n30 VDD2.n11 171.744
R1219 VDD2.n38 VDD2.n11 171.744
R1220 VDD2.n39 VDD2.n38 171.744
R1221 VDD2.n40 VDD2.n39 171.744
R1222 VDD2.n40 VDD2.n7 171.744
R1223 VDD2.n47 VDD2.n7 171.744
R1224 VDD2.n48 VDD2.n47 171.744
R1225 VDD2.n48 VDD2.n3 171.744
R1226 VDD2.n55 VDD2.n3 171.744
R1227 VDD2.n56 VDD2.n55 171.744
R1228 VDD2.n122 VDD2.n60 87.4931
R1229 VDD2.n84 VDD2.t1 85.8723
R1230 VDD2.n21 VDD2.t0 85.8723
R1231 VDD2.n122 VDD2.n121 50.9975
R1232 VDD2.n71 VDD2.n69 13.1884
R1233 VDD2.n41 VDD2.n8 13.1884
R1234 VDD2.n107 VDD2.n106 12.8005
R1235 VDD2.n103 VDD2.n102 12.8005
R1236 VDD2.n42 VDD2.n10 12.8005
R1237 VDD2.n46 VDD2.n45 12.8005
R1238 VDD2.n110 VDD2.n67 12.0247
R1239 VDD2.n99 VDD2.n72 12.0247
R1240 VDD2.n37 VDD2.n36 12.0247
R1241 VDD2.n49 VDD2.n6 12.0247
R1242 VDD2.n111 VDD2.n65 11.249
R1243 VDD2.n98 VDD2.n75 11.249
R1244 VDD2.n35 VDD2.n12 11.249
R1245 VDD2.n50 VDD2.n4 11.249
R1246 VDD2.n83 VDD2.n82 10.7239
R1247 VDD2.n20 VDD2.n19 10.7239
R1248 VDD2.n115 VDD2.n114 10.4732
R1249 VDD2.n95 VDD2.n94 10.4732
R1250 VDD2.n32 VDD2.n31 10.4732
R1251 VDD2.n54 VDD2.n53 10.4732
R1252 VDD2.n118 VDD2.n63 9.69747
R1253 VDD2.n91 VDD2.n77 9.69747
R1254 VDD2.n28 VDD2.n14 9.69747
R1255 VDD2.n57 VDD2.n2 9.69747
R1256 VDD2.n121 VDD2.n120 9.45567
R1257 VDD2.n60 VDD2.n59 9.45567
R1258 VDD2.n81 VDD2.n80 9.3005
R1259 VDD2.n88 VDD2.n87 9.3005
R1260 VDD2.n90 VDD2.n89 9.3005
R1261 VDD2.n77 VDD2.n76 9.3005
R1262 VDD2.n96 VDD2.n95 9.3005
R1263 VDD2.n98 VDD2.n97 9.3005
R1264 VDD2.n72 VDD2.n70 9.3005
R1265 VDD2.n104 VDD2.n103 9.3005
R1266 VDD2.n120 VDD2.n119 9.3005
R1267 VDD2.n63 VDD2.n62 9.3005
R1268 VDD2.n114 VDD2.n113 9.3005
R1269 VDD2.n112 VDD2.n111 9.3005
R1270 VDD2.n67 VDD2.n66 9.3005
R1271 VDD2.n106 VDD2.n105 9.3005
R1272 VDD2.n59 VDD2.n58 9.3005
R1273 VDD2.n2 VDD2.n1 9.3005
R1274 VDD2.n53 VDD2.n52 9.3005
R1275 VDD2.n51 VDD2.n50 9.3005
R1276 VDD2.n6 VDD2.n5 9.3005
R1277 VDD2.n45 VDD2.n44 9.3005
R1278 VDD2.n18 VDD2.n17 9.3005
R1279 VDD2.n25 VDD2.n24 9.3005
R1280 VDD2.n27 VDD2.n26 9.3005
R1281 VDD2.n14 VDD2.n13 9.3005
R1282 VDD2.n33 VDD2.n32 9.3005
R1283 VDD2.n35 VDD2.n34 9.3005
R1284 VDD2.n36 VDD2.n9 9.3005
R1285 VDD2.n43 VDD2.n42 9.3005
R1286 VDD2.n119 VDD2.n61 8.92171
R1287 VDD2.n90 VDD2.n79 8.92171
R1288 VDD2.n27 VDD2.n16 8.92171
R1289 VDD2.n58 VDD2.n0 8.92171
R1290 VDD2.n87 VDD2.n86 8.14595
R1291 VDD2.n24 VDD2.n23 8.14595
R1292 VDD2.n83 VDD2.n81 7.3702
R1293 VDD2.n20 VDD2.n18 7.3702
R1294 VDD2.n86 VDD2.n81 5.81868
R1295 VDD2.n23 VDD2.n18 5.81868
R1296 VDD2.n121 VDD2.n61 5.04292
R1297 VDD2.n87 VDD2.n79 5.04292
R1298 VDD2.n24 VDD2.n16 5.04292
R1299 VDD2.n60 VDD2.n0 5.04292
R1300 VDD2.n119 VDD2.n118 4.26717
R1301 VDD2.n91 VDD2.n90 4.26717
R1302 VDD2.n28 VDD2.n27 4.26717
R1303 VDD2.n58 VDD2.n57 4.26717
R1304 VDD2.n115 VDD2.n63 3.49141
R1305 VDD2.n94 VDD2.n77 3.49141
R1306 VDD2.n31 VDD2.n14 3.49141
R1307 VDD2.n54 VDD2.n2 3.49141
R1308 VDD2.n114 VDD2.n65 2.71565
R1309 VDD2.n95 VDD2.n75 2.71565
R1310 VDD2.n32 VDD2.n12 2.71565
R1311 VDD2.n53 VDD2.n4 2.71565
R1312 VDD2.n82 VDD2.n80 2.41282
R1313 VDD2.n19 VDD2.n17 2.41282
R1314 VDD2.n111 VDD2.n110 1.93989
R1315 VDD2.n99 VDD2.n98 1.93989
R1316 VDD2.n37 VDD2.n35 1.93989
R1317 VDD2.n50 VDD2.n49 1.93989
R1318 VDD2.n107 VDD2.n67 1.16414
R1319 VDD2.n102 VDD2.n72 1.16414
R1320 VDD2.n36 VDD2.n10 1.16414
R1321 VDD2.n46 VDD2.n6 1.16414
R1322 VDD2 VDD2.n122 0.422914
R1323 VDD2.n106 VDD2.n69 0.388379
R1324 VDD2.n103 VDD2.n71 0.388379
R1325 VDD2.n42 VDD2.n41 0.388379
R1326 VDD2.n45 VDD2.n8 0.388379
R1327 VDD2.n120 VDD2.n62 0.155672
R1328 VDD2.n113 VDD2.n62 0.155672
R1329 VDD2.n113 VDD2.n112 0.155672
R1330 VDD2.n112 VDD2.n66 0.155672
R1331 VDD2.n105 VDD2.n66 0.155672
R1332 VDD2.n105 VDD2.n104 0.155672
R1333 VDD2.n104 VDD2.n70 0.155672
R1334 VDD2.n97 VDD2.n70 0.155672
R1335 VDD2.n97 VDD2.n96 0.155672
R1336 VDD2.n96 VDD2.n76 0.155672
R1337 VDD2.n89 VDD2.n76 0.155672
R1338 VDD2.n89 VDD2.n88 0.155672
R1339 VDD2.n88 VDD2.n80 0.155672
R1340 VDD2.n25 VDD2.n17 0.155672
R1341 VDD2.n26 VDD2.n25 0.155672
R1342 VDD2.n26 VDD2.n13 0.155672
R1343 VDD2.n33 VDD2.n13 0.155672
R1344 VDD2.n34 VDD2.n33 0.155672
R1345 VDD2.n34 VDD2.n9 0.155672
R1346 VDD2.n43 VDD2.n9 0.155672
R1347 VDD2.n44 VDD2.n43 0.155672
R1348 VDD2.n44 VDD2.n5 0.155672
R1349 VDD2.n51 VDD2.n5 0.155672
R1350 VDD2.n52 VDD2.n51 0.155672
R1351 VDD2.n52 VDD2.n1 0.155672
R1352 VDD2.n59 VDD2.n1 0.155672
R1353 VP.n0 VP.t0 354.627
R1354 VP.n0 VP.t1 313.63
R1355 VP VP.n0 0.146778
R1356 VDD1.n56 VDD1.n0 756.745
R1357 VDD1.n117 VDD1.n61 756.745
R1358 VDD1.n57 VDD1.n56 585
R1359 VDD1.n55 VDD1.n54 585
R1360 VDD1.n4 VDD1.n3 585
R1361 VDD1.n49 VDD1.n48 585
R1362 VDD1.n47 VDD1.n46 585
R1363 VDD1.n8 VDD1.n7 585
R1364 VDD1.n12 VDD1.n10 585
R1365 VDD1.n41 VDD1.n40 585
R1366 VDD1.n39 VDD1.n38 585
R1367 VDD1.n14 VDD1.n13 585
R1368 VDD1.n33 VDD1.n32 585
R1369 VDD1.n31 VDD1.n30 585
R1370 VDD1.n18 VDD1.n17 585
R1371 VDD1.n25 VDD1.n24 585
R1372 VDD1.n23 VDD1.n22 585
R1373 VDD1.n82 VDD1.n81 585
R1374 VDD1.n84 VDD1.n83 585
R1375 VDD1.n77 VDD1.n76 585
R1376 VDD1.n90 VDD1.n89 585
R1377 VDD1.n92 VDD1.n91 585
R1378 VDD1.n73 VDD1.n72 585
R1379 VDD1.n99 VDD1.n98 585
R1380 VDD1.n100 VDD1.n71 585
R1381 VDD1.n102 VDD1.n101 585
R1382 VDD1.n69 VDD1.n68 585
R1383 VDD1.n108 VDD1.n107 585
R1384 VDD1.n110 VDD1.n109 585
R1385 VDD1.n65 VDD1.n64 585
R1386 VDD1.n116 VDD1.n115 585
R1387 VDD1.n118 VDD1.n117 585
R1388 VDD1.n21 VDD1.t1 329.036
R1389 VDD1.n80 VDD1.t0 329.036
R1390 VDD1.n56 VDD1.n55 171.744
R1391 VDD1.n55 VDD1.n3 171.744
R1392 VDD1.n48 VDD1.n3 171.744
R1393 VDD1.n48 VDD1.n47 171.744
R1394 VDD1.n47 VDD1.n7 171.744
R1395 VDD1.n12 VDD1.n7 171.744
R1396 VDD1.n40 VDD1.n12 171.744
R1397 VDD1.n40 VDD1.n39 171.744
R1398 VDD1.n39 VDD1.n13 171.744
R1399 VDD1.n32 VDD1.n13 171.744
R1400 VDD1.n32 VDD1.n31 171.744
R1401 VDD1.n31 VDD1.n17 171.744
R1402 VDD1.n24 VDD1.n17 171.744
R1403 VDD1.n24 VDD1.n23 171.744
R1404 VDD1.n83 VDD1.n82 171.744
R1405 VDD1.n83 VDD1.n76 171.744
R1406 VDD1.n90 VDD1.n76 171.744
R1407 VDD1.n91 VDD1.n90 171.744
R1408 VDD1.n91 VDD1.n72 171.744
R1409 VDD1.n99 VDD1.n72 171.744
R1410 VDD1.n100 VDD1.n99 171.744
R1411 VDD1.n101 VDD1.n100 171.744
R1412 VDD1.n101 VDD1.n68 171.744
R1413 VDD1.n108 VDD1.n68 171.744
R1414 VDD1.n109 VDD1.n108 171.744
R1415 VDD1.n109 VDD1.n64 171.744
R1416 VDD1.n116 VDD1.n64 171.744
R1417 VDD1.n117 VDD1.n116 171.744
R1418 VDD1 VDD1.n121 88.3822
R1419 VDD1.n23 VDD1.t1 85.8723
R1420 VDD1.n82 VDD1.t0 85.8723
R1421 VDD1 VDD1.n60 51.4199
R1422 VDD1.n10 VDD1.n8 13.1884
R1423 VDD1.n102 VDD1.n69 13.1884
R1424 VDD1.n46 VDD1.n45 12.8005
R1425 VDD1.n42 VDD1.n41 12.8005
R1426 VDD1.n103 VDD1.n71 12.8005
R1427 VDD1.n107 VDD1.n106 12.8005
R1428 VDD1.n49 VDD1.n6 12.0247
R1429 VDD1.n38 VDD1.n11 12.0247
R1430 VDD1.n98 VDD1.n97 12.0247
R1431 VDD1.n110 VDD1.n67 12.0247
R1432 VDD1.n50 VDD1.n4 11.249
R1433 VDD1.n37 VDD1.n14 11.249
R1434 VDD1.n96 VDD1.n73 11.249
R1435 VDD1.n111 VDD1.n65 11.249
R1436 VDD1.n22 VDD1.n21 10.7239
R1437 VDD1.n81 VDD1.n80 10.7239
R1438 VDD1.n54 VDD1.n53 10.4732
R1439 VDD1.n34 VDD1.n33 10.4732
R1440 VDD1.n93 VDD1.n92 10.4732
R1441 VDD1.n115 VDD1.n114 10.4732
R1442 VDD1.n57 VDD1.n2 9.69747
R1443 VDD1.n30 VDD1.n16 9.69747
R1444 VDD1.n89 VDD1.n75 9.69747
R1445 VDD1.n118 VDD1.n63 9.69747
R1446 VDD1.n60 VDD1.n59 9.45567
R1447 VDD1.n121 VDD1.n120 9.45567
R1448 VDD1.n20 VDD1.n19 9.3005
R1449 VDD1.n27 VDD1.n26 9.3005
R1450 VDD1.n29 VDD1.n28 9.3005
R1451 VDD1.n16 VDD1.n15 9.3005
R1452 VDD1.n35 VDD1.n34 9.3005
R1453 VDD1.n37 VDD1.n36 9.3005
R1454 VDD1.n11 VDD1.n9 9.3005
R1455 VDD1.n43 VDD1.n42 9.3005
R1456 VDD1.n59 VDD1.n58 9.3005
R1457 VDD1.n2 VDD1.n1 9.3005
R1458 VDD1.n53 VDD1.n52 9.3005
R1459 VDD1.n51 VDD1.n50 9.3005
R1460 VDD1.n6 VDD1.n5 9.3005
R1461 VDD1.n45 VDD1.n44 9.3005
R1462 VDD1.n120 VDD1.n119 9.3005
R1463 VDD1.n63 VDD1.n62 9.3005
R1464 VDD1.n114 VDD1.n113 9.3005
R1465 VDD1.n112 VDD1.n111 9.3005
R1466 VDD1.n67 VDD1.n66 9.3005
R1467 VDD1.n106 VDD1.n105 9.3005
R1468 VDD1.n79 VDD1.n78 9.3005
R1469 VDD1.n86 VDD1.n85 9.3005
R1470 VDD1.n88 VDD1.n87 9.3005
R1471 VDD1.n75 VDD1.n74 9.3005
R1472 VDD1.n94 VDD1.n93 9.3005
R1473 VDD1.n96 VDD1.n95 9.3005
R1474 VDD1.n97 VDD1.n70 9.3005
R1475 VDD1.n104 VDD1.n103 9.3005
R1476 VDD1.n58 VDD1.n0 8.92171
R1477 VDD1.n29 VDD1.n18 8.92171
R1478 VDD1.n88 VDD1.n77 8.92171
R1479 VDD1.n119 VDD1.n61 8.92171
R1480 VDD1.n26 VDD1.n25 8.14595
R1481 VDD1.n85 VDD1.n84 8.14595
R1482 VDD1.n22 VDD1.n20 7.3702
R1483 VDD1.n81 VDD1.n79 7.3702
R1484 VDD1.n25 VDD1.n20 5.81868
R1485 VDD1.n84 VDD1.n79 5.81868
R1486 VDD1.n60 VDD1.n0 5.04292
R1487 VDD1.n26 VDD1.n18 5.04292
R1488 VDD1.n85 VDD1.n77 5.04292
R1489 VDD1.n121 VDD1.n61 5.04292
R1490 VDD1.n58 VDD1.n57 4.26717
R1491 VDD1.n30 VDD1.n29 4.26717
R1492 VDD1.n89 VDD1.n88 4.26717
R1493 VDD1.n119 VDD1.n118 4.26717
R1494 VDD1.n54 VDD1.n2 3.49141
R1495 VDD1.n33 VDD1.n16 3.49141
R1496 VDD1.n92 VDD1.n75 3.49141
R1497 VDD1.n115 VDD1.n63 3.49141
R1498 VDD1.n53 VDD1.n4 2.71565
R1499 VDD1.n34 VDD1.n14 2.71565
R1500 VDD1.n93 VDD1.n73 2.71565
R1501 VDD1.n114 VDD1.n65 2.71565
R1502 VDD1.n21 VDD1.n19 2.41282
R1503 VDD1.n80 VDD1.n78 2.41282
R1504 VDD1.n50 VDD1.n49 1.93989
R1505 VDD1.n38 VDD1.n37 1.93989
R1506 VDD1.n98 VDD1.n96 1.93989
R1507 VDD1.n111 VDD1.n110 1.93989
R1508 VDD1.n46 VDD1.n6 1.16414
R1509 VDD1.n41 VDD1.n11 1.16414
R1510 VDD1.n97 VDD1.n71 1.16414
R1511 VDD1.n107 VDD1.n67 1.16414
R1512 VDD1.n45 VDD1.n8 0.388379
R1513 VDD1.n42 VDD1.n10 0.388379
R1514 VDD1.n103 VDD1.n102 0.388379
R1515 VDD1.n106 VDD1.n69 0.388379
R1516 VDD1.n59 VDD1.n1 0.155672
R1517 VDD1.n52 VDD1.n1 0.155672
R1518 VDD1.n52 VDD1.n51 0.155672
R1519 VDD1.n51 VDD1.n5 0.155672
R1520 VDD1.n44 VDD1.n5 0.155672
R1521 VDD1.n44 VDD1.n43 0.155672
R1522 VDD1.n43 VDD1.n9 0.155672
R1523 VDD1.n36 VDD1.n9 0.155672
R1524 VDD1.n36 VDD1.n35 0.155672
R1525 VDD1.n35 VDD1.n15 0.155672
R1526 VDD1.n28 VDD1.n15 0.155672
R1527 VDD1.n28 VDD1.n27 0.155672
R1528 VDD1.n27 VDD1.n19 0.155672
R1529 VDD1.n86 VDD1.n78 0.155672
R1530 VDD1.n87 VDD1.n86 0.155672
R1531 VDD1.n87 VDD1.n74 0.155672
R1532 VDD1.n94 VDD1.n74 0.155672
R1533 VDD1.n95 VDD1.n94 0.155672
R1534 VDD1.n95 VDD1.n70 0.155672
R1535 VDD1.n104 VDD1.n70 0.155672
R1536 VDD1.n105 VDD1.n104 0.155672
R1537 VDD1.n105 VDD1.n66 0.155672
R1538 VDD1.n112 VDD1.n66 0.155672
R1539 VDD1.n113 VDD1.n112 0.155672
R1540 VDD1.n113 VDD1.n62 0.155672
R1541 VDD1.n120 VDD1.n62 0.155672
C0 VTAIL VDD1 4.95625f
C1 w_n1646_n3270# VN 2.15445f
C2 VDD2 B 1.50879f
C3 w_n1646_n3270# VP 2.36144f
C4 VN VP 4.78275f
C5 B VDD1 1.48945f
C6 VDD2 VDD1 0.530565f
C7 VTAIL w_n1646_n3270# 2.72641f
C8 VTAIL VN 1.95103f
C9 VTAIL VP 1.96546f
C10 w_n1646_n3270# B 7.33069f
C11 VN B 0.834393f
C12 w_n1646_n3270# VDD2 1.61911f
C13 VN VDD2 2.34853f
C14 B VP 1.16973f
C15 w_n1646_n3270# VDD1 1.60781f
C16 VDD2 VP 0.281086f
C17 VN VDD1 0.147554f
C18 VTAIL B 2.98381f
C19 VTAIL VDD2 4.99674f
C20 VP VDD1 2.47872f
C21 VDD2 VSUBS 0.777155f
C22 VDD1 VSUBS 3.282036f
C23 VTAIL VSUBS 0.812528f
C24 VN VSUBS 6.508309f
C25 VP VSUBS 1.28914f
C26 B VSUBS 2.936546f
C27 w_n1646_n3270# VSUBS 66.3075f
C28 VDD1.n0 VSUBS 0.02305f
C29 VDD1.n1 VSUBS 0.020502f
C30 VDD1.n2 VSUBS 0.011017f
C31 VDD1.n3 VSUBS 0.026039f
C32 VDD1.n4 VSUBS 0.011665f
C33 VDD1.n5 VSUBS 0.020502f
C34 VDD1.n6 VSUBS 0.011017f
C35 VDD1.n7 VSUBS 0.026039f
C36 VDD1.n8 VSUBS 0.011341f
C37 VDD1.n9 VSUBS 0.020502f
C38 VDD1.n10 VSUBS 0.011341f
C39 VDD1.n11 VSUBS 0.011017f
C40 VDD1.n12 VSUBS 0.026039f
C41 VDD1.n13 VSUBS 0.026039f
C42 VDD1.n14 VSUBS 0.011665f
C43 VDD1.n15 VSUBS 0.020502f
C44 VDD1.n16 VSUBS 0.011017f
C45 VDD1.n17 VSUBS 0.026039f
C46 VDD1.n18 VSUBS 0.011665f
C47 VDD1.n19 VSUBS 0.963288f
C48 VDD1.n20 VSUBS 0.011017f
C49 VDD1.t1 VSUBS 0.056083f
C50 VDD1.n21 VSUBS 0.156924f
C51 VDD1.n22 VSUBS 0.019588f
C52 VDD1.n23 VSUBS 0.01953f
C53 VDD1.n24 VSUBS 0.026039f
C54 VDD1.n25 VSUBS 0.011665f
C55 VDD1.n26 VSUBS 0.011017f
C56 VDD1.n27 VSUBS 0.020502f
C57 VDD1.n28 VSUBS 0.020502f
C58 VDD1.n29 VSUBS 0.011017f
C59 VDD1.n30 VSUBS 0.011665f
C60 VDD1.n31 VSUBS 0.026039f
C61 VDD1.n32 VSUBS 0.026039f
C62 VDD1.n33 VSUBS 0.011665f
C63 VDD1.n34 VSUBS 0.011017f
C64 VDD1.n35 VSUBS 0.020502f
C65 VDD1.n36 VSUBS 0.020502f
C66 VDD1.n37 VSUBS 0.011017f
C67 VDD1.n38 VSUBS 0.011665f
C68 VDD1.n39 VSUBS 0.026039f
C69 VDD1.n40 VSUBS 0.026039f
C70 VDD1.n41 VSUBS 0.011665f
C71 VDD1.n42 VSUBS 0.011017f
C72 VDD1.n43 VSUBS 0.020502f
C73 VDD1.n44 VSUBS 0.020502f
C74 VDD1.n45 VSUBS 0.011017f
C75 VDD1.n46 VSUBS 0.011665f
C76 VDD1.n47 VSUBS 0.026039f
C77 VDD1.n48 VSUBS 0.026039f
C78 VDD1.n49 VSUBS 0.011665f
C79 VDD1.n50 VSUBS 0.011017f
C80 VDD1.n51 VSUBS 0.020502f
C81 VDD1.n52 VSUBS 0.020502f
C82 VDD1.n53 VSUBS 0.011017f
C83 VDD1.n54 VSUBS 0.011665f
C84 VDD1.n55 VSUBS 0.026039f
C85 VDD1.n56 VSUBS 0.064819f
C86 VDD1.n57 VSUBS 0.011665f
C87 VDD1.n58 VSUBS 0.011017f
C88 VDD1.n59 VSUBS 0.05047f
C89 VDD1.n60 VSUBS 0.047469f
C90 VDD1.n61 VSUBS 0.02305f
C91 VDD1.n62 VSUBS 0.020502f
C92 VDD1.n63 VSUBS 0.011017f
C93 VDD1.n64 VSUBS 0.026039f
C94 VDD1.n65 VSUBS 0.011665f
C95 VDD1.n66 VSUBS 0.020502f
C96 VDD1.n67 VSUBS 0.011017f
C97 VDD1.n68 VSUBS 0.026039f
C98 VDD1.n69 VSUBS 0.011341f
C99 VDD1.n70 VSUBS 0.020502f
C100 VDD1.n71 VSUBS 0.011665f
C101 VDD1.n72 VSUBS 0.026039f
C102 VDD1.n73 VSUBS 0.011665f
C103 VDD1.n74 VSUBS 0.020502f
C104 VDD1.n75 VSUBS 0.011017f
C105 VDD1.n76 VSUBS 0.026039f
C106 VDD1.n77 VSUBS 0.011665f
C107 VDD1.n78 VSUBS 0.963288f
C108 VDD1.n79 VSUBS 0.011017f
C109 VDD1.t0 VSUBS 0.056083f
C110 VDD1.n80 VSUBS 0.156924f
C111 VDD1.n81 VSUBS 0.019588f
C112 VDD1.n82 VSUBS 0.01953f
C113 VDD1.n83 VSUBS 0.026039f
C114 VDD1.n84 VSUBS 0.011665f
C115 VDD1.n85 VSUBS 0.011017f
C116 VDD1.n86 VSUBS 0.020502f
C117 VDD1.n87 VSUBS 0.020502f
C118 VDD1.n88 VSUBS 0.011017f
C119 VDD1.n89 VSUBS 0.011665f
C120 VDD1.n90 VSUBS 0.026039f
C121 VDD1.n91 VSUBS 0.026039f
C122 VDD1.n92 VSUBS 0.011665f
C123 VDD1.n93 VSUBS 0.011017f
C124 VDD1.n94 VSUBS 0.020502f
C125 VDD1.n95 VSUBS 0.020502f
C126 VDD1.n96 VSUBS 0.011017f
C127 VDD1.n97 VSUBS 0.011017f
C128 VDD1.n98 VSUBS 0.011665f
C129 VDD1.n99 VSUBS 0.026039f
C130 VDD1.n100 VSUBS 0.026039f
C131 VDD1.n101 VSUBS 0.026039f
C132 VDD1.n102 VSUBS 0.011341f
C133 VDD1.n103 VSUBS 0.011017f
C134 VDD1.n104 VSUBS 0.020502f
C135 VDD1.n105 VSUBS 0.020502f
C136 VDD1.n106 VSUBS 0.011017f
C137 VDD1.n107 VSUBS 0.011665f
C138 VDD1.n108 VSUBS 0.026039f
C139 VDD1.n109 VSUBS 0.026039f
C140 VDD1.n110 VSUBS 0.011665f
C141 VDD1.n111 VSUBS 0.011017f
C142 VDD1.n112 VSUBS 0.020502f
C143 VDD1.n113 VSUBS 0.020502f
C144 VDD1.n114 VSUBS 0.011017f
C145 VDD1.n115 VSUBS 0.011665f
C146 VDD1.n116 VSUBS 0.026039f
C147 VDD1.n117 VSUBS 0.064819f
C148 VDD1.n118 VSUBS 0.011665f
C149 VDD1.n119 VSUBS 0.011017f
C150 VDD1.n120 VSUBS 0.05047f
C151 VDD1.n121 VSUBS 0.544584f
C152 VP.t0 VSUBS 2.60216f
C153 VP.t1 VSUBS 2.31102f
C154 VP.n0 VSUBS 4.74214f
C155 VDD2.n0 VSUBS 0.022664f
C156 VDD2.n1 VSUBS 0.020159f
C157 VDD2.n2 VSUBS 0.010832f
C158 VDD2.n3 VSUBS 0.025604f
C159 VDD2.n4 VSUBS 0.011469f
C160 VDD2.n5 VSUBS 0.020159f
C161 VDD2.n6 VSUBS 0.010832f
C162 VDD2.n7 VSUBS 0.025604f
C163 VDD2.n8 VSUBS 0.011151f
C164 VDD2.n9 VSUBS 0.020159f
C165 VDD2.n10 VSUBS 0.011469f
C166 VDD2.n11 VSUBS 0.025604f
C167 VDD2.n12 VSUBS 0.011469f
C168 VDD2.n13 VSUBS 0.020159f
C169 VDD2.n14 VSUBS 0.010832f
C170 VDD2.n15 VSUBS 0.025604f
C171 VDD2.n16 VSUBS 0.011469f
C172 VDD2.n17 VSUBS 0.947163f
C173 VDD2.n18 VSUBS 0.010832f
C174 VDD2.t0 VSUBS 0.055144f
C175 VDD2.n19 VSUBS 0.154298f
C176 VDD2.n20 VSUBS 0.01926f
C177 VDD2.n21 VSUBS 0.019203f
C178 VDD2.n22 VSUBS 0.025604f
C179 VDD2.n23 VSUBS 0.011469f
C180 VDD2.n24 VSUBS 0.010832f
C181 VDD2.n25 VSUBS 0.020159f
C182 VDD2.n26 VSUBS 0.020159f
C183 VDD2.n27 VSUBS 0.010832f
C184 VDD2.n28 VSUBS 0.011469f
C185 VDD2.n29 VSUBS 0.025604f
C186 VDD2.n30 VSUBS 0.025604f
C187 VDD2.n31 VSUBS 0.011469f
C188 VDD2.n32 VSUBS 0.010832f
C189 VDD2.n33 VSUBS 0.020159f
C190 VDD2.n34 VSUBS 0.020159f
C191 VDD2.n35 VSUBS 0.010832f
C192 VDD2.n36 VSUBS 0.010832f
C193 VDD2.n37 VSUBS 0.011469f
C194 VDD2.n38 VSUBS 0.025604f
C195 VDD2.n39 VSUBS 0.025604f
C196 VDD2.n40 VSUBS 0.025604f
C197 VDD2.n41 VSUBS 0.011151f
C198 VDD2.n42 VSUBS 0.010832f
C199 VDD2.n43 VSUBS 0.020159f
C200 VDD2.n44 VSUBS 0.020159f
C201 VDD2.n45 VSUBS 0.010832f
C202 VDD2.n46 VSUBS 0.011469f
C203 VDD2.n47 VSUBS 0.025604f
C204 VDD2.n48 VSUBS 0.025604f
C205 VDD2.n49 VSUBS 0.011469f
C206 VDD2.n50 VSUBS 0.010832f
C207 VDD2.n51 VSUBS 0.020159f
C208 VDD2.n52 VSUBS 0.020159f
C209 VDD2.n53 VSUBS 0.010832f
C210 VDD2.n54 VSUBS 0.011469f
C211 VDD2.n55 VSUBS 0.025604f
C212 VDD2.n56 VSUBS 0.063734f
C213 VDD2.n57 VSUBS 0.011469f
C214 VDD2.n58 VSUBS 0.010832f
C215 VDD2.n59 VSUBS 0.049625f
C216 VDD2.n60 VSUBS 0.505266f
C217 VDD2.n61 VSUBS 0.022664f
C218 VDD2.n62 VSUBS 0.020159f
C219 VDD2.n63 VSUBS 0.010832f
C220 VDD2.n64 VSUBS 0.025604f
C221 VDD2.n65 VSUBS 0.011469f
C222 VDD2.n66 VSUBS 0.020159f
C223 VDD2.n67 VSUBS 0.010832f
C224 VDD2.n68 VSUBS 0.025604f
C225 VDD2.n69 VSUBS 0.011151f
C226 VDD2.n70 VSUBS 0.020159f
C227 VDD2.n71 VSUBS 0.011151f
C228 VDD2.n72 VSUBS 0.010832f
C229 VDD2.n73 VSUBS 0.025604f
C230 VDD2.n74 VSUBS 0.025604f
C231 VDD2.n75 VSUBS 0.011469f
C232 VDD2.n76 VSUBS 0.020159f
C233 VDD2.n77 VSUBS 0.010832f
C234 VDD2.n78 VSUBS 0.025604f
C235 VDD2.n79 VSUBS 0.011469f
C236 VDD2.n80 VSUBS 0.947163f
C237 VDD2.n81 VSUBS 0.010832f
C238 VDD2.t1 VSUBS 0.055144f
C239 VDD2.n82 VSUBS 0.154298f
C240 VDD2.n83 VSUBS 0.01926f
C241 VDD2.n84 VSUBS 0.019203f
C242 VDD2.n85 VSUBS 0.025604f
C243 VDD2.n86 VSUBS 0.011469f
C244 VDD2.n87 VSUBS 0.010832f
C245 VDD2.n88 VSUBS 0.020159f
C246 VDD2.n89 VSUBS 0.020159f
C247 VDD2.n90 VSUBS 0.010832f
C248 VDD2.n91 VSUBS 0.011469f
C249 VDD2.n92 VSUBS 0.025604f
C250 VDD2.n93 VSUBS 0.025604f
C251 VDD2.n94 VSUBS 0.011469f
C252 VDD2.n95 VSUBS 0.010832f
C253 VDD2.n96 VSUBS 0.020159f
C254 VDD2.n97 VSUBS 0.020159f
C255 VDD2.n98 VSUBS 0.010832f
C256 VDD2.n99 VSUBS 0.011469f
C257 VDD2.n100 VSUBS 0.025604f
C258 VDD2.n101 VSUBS 0.025604f
C259 VDD2.n102 VSUBS 0.011469f
C260 VDD2.n103 VSUBS 0.010832f
C261 VDD2.n104 VSUBS 0.020159f
C262 VDD2.n105 VSUBS 0.020159f
C263 VDD2.n106 VSUBS 0.010832f
C264 VDD2.n107 VSUBS 0.011469f
C265 VDD2.n108 VSUBS 0.025604f
C266 VDD2.n109 VSUBS 0.025604f
C267 VDD2.n110 VSUBS 0.011469f
C268 VDD2.n111 VSUBS 0.010832f
C269 VDD2.n112 VSUBS 0.020159f
C270 VDD2.n113 VSUBS 0.020159f
C271 VDD2.n114 VSUBS 0.010832f
C272 VDD2.n115 VSUBS 0.011469f
C273 VDD2.n116 VSUBS 0.025604f
C274 VDD2.n117 VSUBS 0.063734f
C275 VDD2.n118 VSUBS 0.011469f
C276 VDD2.n119 VSUBS 0.010832f
C277 VDD2.n120 VSUBS 0.049625f
C278 VDD2.n121 VSUBS 0.046116f
C279 VDD2.n122 VSUBS 2.23845f
C280 VTAIL.n0 VSUBS 0.026112f
C281 VTAIL.n1 VSUBS 0.023225f
C282 VTAIL.n2 VSUBS 0.01248f
C283 VTAIL.n3 VSUBS 0.029499f
C284 VTAIL.n4 VSUBS 0.013215f
C285 VTAIL.n5 VSUBS 0.023225f
C286 VTAIL.n6 VSUBS 0.01248f
C287 VTAIL.n7 VSUBS 0.029499f
C288 VTAIL.n8 VSUBS 0.012847f
C289 VTAIL.n9 VSUBS 0.023225f
C290 VTAIL.n10 VSUBS 0.013215f
C291 VTAIL.n11 VSUBS 0.029499f
C292 VTAIL.n12 VSUBS 0.013215f
C293 VTAIL.n13 VSUBS 0.023225f
C294 VTAIL.n14 VSUBS 0.01248f
C295 VTAIL.n15 VSUBS 0.029499f
C296 VTAIL.n16 VSUBS 0.013215f
C297 VTAIL.n17 VSUBS 1.09127f
C298 VTAIL.n18 VSUBS 0.01248f
C299 VTAIL.t1 VSUBS 0.063534f
C300 VTAIL.n19 VSUBS 0.177773f
C301 VTAIL.n20 VSUBS 0.022191f
C302 VTAIL.n21 VSUBS 0.022124f
C303 VTAIL.n22 VSUBS 0.029499f
C304 VTAIL.n23 VSUBS 0.013215f
C305 VTAIL.n24 VSUBS 0.01248f
C306 VTAIL.n25 VSUBS 0.023225f
C307 VTAIL.n26 VSUBS 0.023225f
C308 VTAIL.n27 VSUBS 0.01248f
C309 VTAIL.n28 VSUBS 0.013215f
C310 VTAIL.n29 VSUBS 0.029499f
C311 VTAIL.n30 VSUBS 0.029499f
C312 VTAIL.n31 VSUBS 0.013215f
C313 VTAIL.n32 VSUBS 0.01248f
C314 VTAIL.n33 VSUBS 0.023225f
C315 VTAIL.n34 VSUBS 0.023225f
C316 VTAIL.n35 VSUBS 0.01248f
C317 VTAIL.n36 VSUBS 0.01248f
C318 VTAIL.n37 VSUBS 0.013215f
C319 VTAIL.n38 VSUBS 0.029499f
C320 VTAIL.n39 VSUBS 0.029499f
C321 VTAIL.n40 VSUBS 0.029499f
C322 VTAIL.n41 VSUBS 0.012847f
C323 VTAIL.n42 VSUBS 0.01248f
C324 VTAIL.n43 VSUBS 0.023225f
C325 VTAIL.n44 VSUBS 0.023225f
C326 VTAIL.n45 VSUBS 0.01248f
C327 VTAIL.n46 VSUBS 0.013215f
C328 VTAIL.n47 VSUBS 0.029499f
C329 VTAIL.n48 VSUBS 0.029499f
C330 VTAIL.n49 VSUBS 0.013215f
C331 VTAIL.n50 VSUBS 0.01248f
C332 VTAIL.n51 VSUBS 0.023225f
C333 VTAIL.n52 VSUBS 0.023225f
C334 VTAIL.n53 VSUBS 0.01248f
C335 VTAIL.n54 VSUBS 0.013215f
C336 VTAIL.n55 VSUBS 0.029499f
C337 VTAIL.n56 VSUBS 0.07343f
C338 VTAIL.n57 VSUBS 0.013215f
C339 VTAIL.n58 VSUBS 0.01248f
C340 VTAIL.n59 VSUBS 0.057175f
C341 VTAIL.n60 VSUBS 0.037121f
C342 VTAIL.n61 VSUBS 1.3647f
C343 VTAIL.n62 VSUBS 0.026112f
C344 VTAIL.n63 VSUBS 0.023225f
C345 VTAIL.n64 VSUBS 0.01248f
C346 VTAIL.n65 VSUBS 0.029499f
C347 VTAIL.n66 VSUBS 0.013215f
C348 VTAIL.n67 VSUBS 0.023225f
C349 VTAIL.n68 VSUBS 0.01248f
C350 VTAIL.n69 VSUBS 0.029499f
C351 VTAIL.n70 VSUBS 0.012847f
C352 VTAIL.n71 VSUBS 0.023225f
C353 VTAIL.n72 VSUBS 0.012847f
C354 VTAIL.n73 VSUBS 0.01248f
C355 VTAIL.n74 VSUBS 0.029499f
C356 VTAIL.n75 VSUBS 0.029499f
C357 VTAIL.n76 VSUBS 0.013215f
C358 VTAIL.n77 VSUBS 0.023225f
C359 VTAIL.n78 VSUBS 0.01248f
C360 VTAIL.n79 VSUBS 0.029499f
C361 VTAIL.n80 VSUBS 0.013215f
C362 VTAIL.n81 VSUBS 1.09127f
C363 VTAIL.n82 VSUBS 0.01248f
C364 VTAIL.t3 VSUBS 0.063534f
C365 VTAIL.n83 VSUBS 0.177773f
C366 VTAIL.n84 VSUBS 0.022191f
C367 VTAIL.n85 VSUBS 0.022124f
C368 VTAIL.n86 VSUBS 0.029499f
C369 VTAIL.n87 VSUBS 0.013215f
C370 VTAIL.n88 VSUBS 0.01248f
C371 VTAIL.n89 VSUBS 0.023225f
C372 VTAIL.n90 VSUBS 0.023225f
C373 VTAIL.n91 VSUBS 0.01248f
C374 VTAIL.n92 VSUBS 0.013215f
C375 VTAIL.n93 VSUBS 0.029499f
C376 VTAIL.n94 VSUBS 0.029499f
C377 VTAIL.n95 VSUBS 0.013215f
C378 VTAIL.n96 VSUBS 0.01248f
C379 VTAIL.n97 VSUBS 0.023225f
C380 VTAIL.n98 VSUBS 0.023225f
C381 VTAIL.n99 VSUBS 0.01248f
C382 VTAIL.n100 VSUBS 0.013215f
C383 VTAIL.n101 VSUBS 0.029499f
C384 VTAIL.n102 VSUBS 0.029499f
C385 VTAIL.n103 VSUBS 0.013215f
C386 VTAIL.n104 VSUBS 0.01248f
C387 VTAIL.n105 VSUBS 0.023225f
C388 VTAIL.n106 VSUBS 0.023225f
C389 VTAIL.n107 VSUBS 0.01248f
C390 VTAIL.n108 VSUBS 0.013215f
C391 VTAIL.n109 VSUBS 0.029499f
C392 VTAIL.n110 VSUBS 0.029499f
C393 VTAIL.n111 VSUBS 0.013215f
C394 VTAIL.n112 VSUBS 0.01248f
C395 VTAIL.n113 VSUBS 0.023225f
C396 VTAIL.n114 VSUBS 0.023225f
C397 VTAIL.n115 VSUBS 0.01248f
C398 VTAIL.n116 VSUBS 0.013215f
C399 VTAIL.n117 VSUBS 0.029499f
C400 VTAIL.n118 VSUBS 0.07343f
C401 VTAIL.n119 VSUBS 0.013215f
C402 VTAIL.n120 VSUBS 0.01248f
C403 VTAIL.n121 VSUBS 0.057175f
C404 VTAIL.n122 VSUBS 0.037121f
C405 VTAIL.n123 VSUBS 1.38761f
C406 VTAIL.n124 VSUBS 0.026112f
C407 VTAIL.n125 VSUBS 0.023225f
C408 VTAIL.n126 VSUBS 0.01248f
C409 VTAIL.n127 VSUBS 0.029499f
C410 VTAIL.n128 VSUBS 0.013215f
C411 VTAIL.n129 VSUBS 0.023225f
C412 VTAIL.n130 VSUBS 0.01248f
C413 VTAIL.n131 VSUBS 0.029499f
C414 VTAIL.n132 VSUBS 0.012847f
C415 VTAIL.n133 VSUBS 0.023225f
C416 VTAIL.n134 VSUBS 0.012847f
C417 VTAIL.n135 VSUBS 0.01248f
C418 VTAIL.n136 VSUBS 0.029499f
C419 VTAIL.n137 VSUBS 0.029499f
C420 VTAIL.n138 VSUBS 0.013215f
C421 VTAIL.n139 VSUBS 0.023225f
C422 VTAIL.n140 VSUBS 0.01248f
C423 VTAIL.n141 VSUBS 0.029499f
C424 VTAIL.n142 VSUBS 0.013215f
C425 VTAIL.n143 VSUBS 1.09127f
C426 VTAIL.n144 VSUBS 0.01248f
C427 VTAIL.t0 VSUBS 0.063534f
C428 VTAIL.n145 VSUBS 0.177773f
C429 VTAIL.n146 VSUBS 0.022191f
C430 VTAIL.n147 VSUBS 0.022124f
C431 VTAIL.n148 VSUBS 0.029499f
C432 VTAIL.n149 VSUBS 0.013215f
C433 VTAIL.n150 VSUBS 0.01248f
C434 VTAIL.n151 VSUBS 0.023225f
C435 VTAIL.n152 VSUBS 0.023225f
C436 VTAIL.n153 VSUBS 0.01248f
C437 VTAIL.n154 VSUBS 0.013215f
C438 VTAIL.n155 VSUBS 0.029499f
C439 VTAIL.n156 VSUBS 0.029499f
C440 VTAIL.n157 VSUBS 0.013215f
C441 VTAIL.n158 VSUBS 0.01248f
C442 VTAIL.n159 VSUBS 0.023225f
C443 VTAIL.n160 VSUBS 0.023225f
C444 VTAIL.n161 VSUBS 0.01248f
C445 VTAIL.n162 VSUBS 0.013215f
C446 VTAIL.n163 VSUBS 0.029499f
C447 VTAIL.n164 VSUBS 0.029499f
C448 VTAIL.n165 VSUBS 0.013215f
C449 VTAIL.n166 VSUBS 0.01248f
C450 VTAIL.n167 VSUBS 0.023225f
C451 VTAIL.n168 VSUBS 0.023225f
C452 VTAIL.n169 VSUBS 0.01248f
C453 VTAIL.n170 VSUBS 0.013215f
C454 VTAIL.n171 VSUBS 0.029499f
C455 VTAIL.n172 VSUBS 0.029499f
C456 VTAIL.n173 VSUBS 0.013215f
C457 VTAIL.n174 VSUBS 0.01248f
C458 VTAIL.n175 VSUBS 0.023225f
C459 VTAIL.n176 VSUBS 0.023225f
C460 VTAIL.n177 VSUBS 0.01248f
C461 VTAIL.n178 VSUBS 0.013215f
C462 VTAIL.n179 VSUBS 0.029499f
C463 VTAIL.n180 VSUBS 0.07343f
C464 VTAIL.n181 VSUBS 0.013215f
C465 VTAIL.n182 VSUBS 0.01248f
C466 VTAIL.n183 VSUBS 0.057175f
C467 VTAIL.n184 VSUBS 0.037121f
C468 VTAIL.n185 VSUBS 1.27857f
C469 VTAIL.n186 VSUBS 0.026112f
C470 VTAIL.n187 VSUBS 0.023225f
C471 VTAIL.n188 VSUBS 0.01248f
C472 VTAIL.n189 VSUBS 0.029499f
C473 VTAIL.n190 VSUBS 0.013215f
C474 VTAIL.n191 VSUBS 0.023225f
C475 VTAIL.n192 VSUBS 0.01248f
C476 VTAIL.n193 VSUBS 0.029499f
C477 VTAIL.n194 VSUBS 0.012847f
C478 VTAIL.n195 VSUBS 0.023225f
C479 VTAIL.n196 VSUBS 0.013215f
C480 VTAIL.n197 VSUBS 0.029499f
C481 VTAIL.n198 VSUBS 0.013215f
C482 VTAIL.n199 VSUBS 0.023225f
C483 VTAIL.n200 VSUBS 0.01248f
C484 VTAIL.n201 VSUBS 0.029499f
C485 VTAIL.n202 VSUBS 0.013215f
C486 VTAIL.n203 VSUBS 1.09127f
C487 VTAIL.n204 VSUBS 0.01248f
C488 VTAIL.t2 VSUBS 0.063534f
C489 VTAIL.n205 VSUBS 0.177773f
C490 VTAIL.n206 VSUBS 0.022191f
C491 VTAIL.n207 VSUBS 0.022124f
C492 VTAIL.n208 VSUBS 0.029499f
C493 VTAIL.n209 VSUBS 0.013215f
C494 VTAIL.n210 VSUBS 0.01248f
C495 VTAIL.n211 VSUBS 0.023225f
C496 VTAIL.n212 VSUBS 0.023225f
C497 VTAIL.n213 VSUBS 0.01248f
C498 VTAIL.n214 VSUBS 0.013215f
C499 VTAIL.n215 VSUBS 0.029499f
C500 VTAIL.n216 VSUBS 0.029499f
C501 VTAIL.n217 VSUBS 0.013215f
C502 VTAIL.n218 VSUBS 0.01248f
C503 VTAIL.n219 VSUBS 0.023225f
C504 VTAIL.n220 VSUBS 0.023225f
C505 VTAIL.n221 VSUBS 0.01248f
C506 VTAIL.n222 VSUBS 0.01248f
C507 VTAIL.n223 VSUBS 0.013215f
C508 VTAIL.n224 VSUBS 0.029499f
C509 VTAIL.n225 VSUBS 0.029499f
C510 VTAIL.n226 VSUBS 0.029499f
C511 VTAIL.n227 VSUBS 0.012847f
C512 VTAIL.n228 VSUBS 0.01248f
C513 VTAIL.n229 VSUBS 0.023225f
C514 VTAIL.n230 VSUBS 0.023225f
C515 VTAIL.n231 VSUBS 0.01248f
C516 VTAIL.n232 VSUBS 0.013215f
C517 VTAIL.n233 VSUBS 0.029499f
C518 VTAIL.n234 VSUBS 0.029499f
C519 VTAIL.n235 VSUBS 0.013215f
C520 VTAIL.n236 VSUBS 0.01248f
C521 VTAIL.n237 VSUBS 0.023225f
C522 VTAIL.n238 VSUBS 0.023225f
C523 VTAIL.n239 VSUBS 0.01248f
C524 VTAIL.n240 VSUBS 0.013215f
C525 VTAIL.n241 VSUBS 0.029499f
C526 VTAIL.n242 VSUBS 0.07343f
C527 VTAIL.n243 VSUBS 0.013215f
C528 VTAIL.n244 VSUBS 0.01248f
C529 VTAIL.n245 VSUBS 0.057175f
C530 VTAIL.n246 VSUBS 0.037121f
C531 VTAIL.n247 VSUBS 1.2118f
C532 VN.t1 VSUBS 2.20105f
C533 VN.t0 VSUBS 2.48263f
C534 B.n0 VSUBS 0.004354f
C535 B.n1 VSUBS 0.004354f
C536 B.n2 VSUBS 0.006885f
C537 B.n3 VSUBS 0.006885f
C538 B.n4 VSUBS 0.006885f
C539 B.n5 VSUBS 0.006885f
C540 B.n6 VSUBS 0.006885f
C541 B.n7 VSUBS 0.006885f
C542 B.n8 VSUBS 0.006885f
C543 B.n9 VSUBS 0.006885f
C544 B.n10 VSUBS 0.006885f
C545 B.n11 VSUBS 0.016546f
C546 B.n12 VSUBS 0.006885f
C547 B.n13 VSUBS 0.006885f
C548 B.n14 VSUBS 0.006885f
C549 B.n15 VSUBS 0.006885f
C550 B.n16 VSUBS 0.006885f
C551 B.n17 VSUBS 0.006885f
C552 B.n18 VSUBS 0.006885f
C553 B.n19 VSUBS 0.006885f
C554 B.n20 VSUBS 0.006885f
C555 B.n21 VSUBS 0.006885f
C556 B.n22 VSUBS 0.006885f
C557 B.n23 VSUBS 0.006885f
C558 B.n24 VSUBS 0.006885f
C559 B.n25 VSUBS 0.006885f
C560 B.n26 VSUBS 0.006885f
C561 B.n27 VSUBS 0.006885f
C562 B.n28 VSUBS 0.006885f
C563 B.n29 VSUBS 0.006885f
C564 B.n30 VSUBS 0.006885f
C565 B.n31 VSUBS 0.006885f
C566 B.t2 VSUBS 0.197082f
C567 B.t1 VSUBS 0.215604f
C568 B.t0 VSUBS 0.670239f
C569 B.n32 VSUBS 0.329463f
C570 B.n33 VSUBS 0.235717f
C571 B.n34 VSUBS 0.006885f
C572 B.n35 VSUBS 0.006885f
C573 B.n36 VSUBS 0.006885f
C574 B.n37 VSUBS 0.006885f
C575 B.t8 VSUBS 0.197085f
C576 B.t7 VSUBS 0.215607f
C577 B.t6 VSUBS 0.670239f
C578 B.n38 VSUBS 0.32946f
C579 B.n39 VSUBS 0.235714f
C580 B.n40 VSUBS 0.015953f
C581 B.n41 VSUBS 0.006885f
C582 B.n42 VSUBS 0.006885f
C583 B.n43 VSUBS 0.006885f
C584 B.n44 VSUBS 0.006885f
C585 B.n45 VSUBS 0.006885f
C586 B.n46 VSUBS 0.006885f
C587 B.n47 VSUBS 0.006885f
C588 B.n48 VSUBS 0.006885f
C589 B.n49 VSUBS 0.006885f
C590 B.n50 VSUBS 0.006885f
C591 B.n51 VSUBS 0.006885f
C592 B.n52 VSUBS 0.006885f
C593 B.n53 VSUBS 0.006885f
C594 B.n54 VSUBS 0.006885f
C595 B.n55 VSUBS 0.006885f
C596 B.n56 VSUBS 0.006885f
C597 B.n57 VSUBS 0.006885f
C598 B.n58 VSUBS 0.006885f
C599 B.n59 VSUBS 0.006885f
C600 B.n60 VSUBS 0.015732f
C601 B.n61 VSUBS 0.006885f
C602 B.n62 VSUBS 0.006885f
C603 B.n63 VSUBS 0.006885f
C604 B.n64 VSUBS 0.006885f
C605 B.n65 VSUBS 0.006885f
C606 B.n66 VSUBS 0.006885f
C607 B.n67 VSUBS 0.006885f
C608 B.n68 VSUBS 0.006885f
C609 B.n69 VSUBS 0.006885f
C610 B.n70 VSUBS 0.006885f
C611 B.n71 VSUBS 0.006885f
C612 B.n72 VSUBS 0.006885f
C613 B.n73 VSUBS 0.006885f
C614 B.n74 VSUBS 0.006885f
C615 B.n75 VSUBS 0.006885f
C616 B.n76 VSUBS 0.006885f
C617 B.n77 VSUBS 0.006885f
C618 B.n78 VSUBS 0.006885f
C619 B.n79 VSUBS 0.016546f
C620 B.n80 VSUBS 0.006885f
C621 B.n81 VSUBS 0.006885f
C622 B.n82 VSUBS 0.006885f
C623 B.n83 VSUBS 0.006885f
C624 B.n84 VSUBS 0.006885f
C625 B.n85 VSUBS 0.006885f
C626 B.n86 VSUBS 0.006885f
C627 B.n87 VSUBS 0.006885f
C628 B.n88 VSUBS 0.006885f
C629 B.n89 VSUBS 0.006885f
C630 B.n90 VSUBS 0.006885f
C631 B.n91 VSUBS 0.006885f
C632 B.n92 VSUBS 0.006885f
C633 B.n93 VSUBS 0.006885f
C634 B.n94 VSUBS 0.006885f
C635 B.n95 VSUBS 0.006885f
C636 B.n96 VSUBS 0.006885f
C637 B.n97 VSUBS 0.006885f
C638 B.n98 VSUBS 0.006885f
C639 B.n99 VSUBS 0.006885f
C640 B.t10 VSUBS 0.197085f
C641 B.t11 VSUBS 0.215607f
C642 B.t9 VSUBS 0.670239f
C643 B.n100 VSUBS 0.32946f
C644 B.n101 VSUBS 0.235714f
C645 B.n102 VSUBS 0.006885f
C646 B.n103 VSUBS 0.006885f
C647 B.n104 VSUBS 0.006885f
C648 B.n105 VSUBS 0.006885f
C649 B.t4 VSUBS 0.197082f
C650 B.t5 VSUBS 0.215604f
C651 B.t3 VSUBS 0.670239f
C652 B.n106 VSUBS 0.329463f
C653 B.n107 VSUBS 0.235717f
C654 B.n108 VSUBS 0.015953f
C655 B.n109 VSUBS 0.006885f
C656 B.n110 VSUBS 0.006885f
C657 B.n111 VSUBS 0.006885f
C658 B.n112 VSUBS 0.006885f
C659 B.n113 VSUBS 0.006885f
C660 B.n114 VSUBS 0.006885f
C661 B.n115 VSUBS 0.006885f
C662 B.n116 VSUBS 0.006885f
C663 B.n117 VSUBS 0.006885f
C664 B.n118 VSUBS 0.006885f
C665 B.n119 VSUBS 0.006885f
C666 B.n120 VSUBS 0.006885f
C667 B.n121 VSUBS 0.006885f
C668 B.n122 VSUBS 0.006885f
C669 B.n123 VSUBS 0.006885f
C670 B.n124 VSUBS 0.006885f
C671 B.n125 VSUBS 0.006885f
C672 B.n126 VSUBS 0.006885f
C673 B.n127 VSUBS 0.006885f
C674 B.n128 VSUBS 0.016546f
C675 B.n129 VSUBS 0.006885f
C676 B.n130 VSUBS 0.006885f
C677 B.n131 VSUBS 0.006885f
C678 B.n132 VSUBS 0.006885f
C679 B.n133 VSUBS 0.006885f
C680 B.n134 VSUBS 0.006885f
C681 B.n135 VSUBS 0.006885f
C682 B.n136 VSUBS 0.006885f
C683 B.n137 VSUBS 0.006885f
C684 B.n138 VSUBS 0.006885f
C685 B.n139 VSUBS 0.006885f
C686 B.n140 VSUBS 0.006885f
C687 B.n141 VSUBS 0.006885f
C688 B.n142 VSUBS 0.006885f
C689 B.n143 VSUBS 0.006885f
C690 B.n144 VSUBS 0.006885f
C691 B.n145 VSUBS 0.006885f
C692 B.n146 VSUBS 0.006885f
C693 B.n147 VSUBS 0.006885f
C694 B.n148 VSUBS 0.006885f
C695 B.n149 VSUBS 0.006885f
C696 B.n150 VSUBS 0.006885f
C697 B.n151 VSUBS 0.006885f
C698 B.n152 VSUBS 0.006885f
C699 B.n153 VSUBS 0.006885f
C700 B.n154 VSUBS 0.006885f
C701 B.n155 VSUBS 0.006885f
C702 B.n156 VSUBS 0.006885f
C703 B.n157 VSUBS 0.006885f
C704 B.n158 VSUBS 0.006885f
C705 B.n159 VSUBS 0.006885f
C706 B.n160 VSUBS 0.006885f
C707 B.n161 VSUBS 0.015653f
C708 B.n162 VSUBS 0.015653f
C709 B.n163 VSUBS 0.016546f
C710 B.n164 VSUBS 0.006885f
C711 B.n165 VSUBS 0.006885f
C712 B.n166 VSUBS 0.006885f
C713 B.n167 VSUBS 0.006885f
C714 B.n168 VSUBS 0.006885f
C715 B.n169 VSUBS 0.006885f
C716 B.n170 VSUBS 0.006885f
C717 B.n171 VSUBS 0.006885f
C718 B.n172 VSUBS 0.006885f
C719 B.n173 VSUBS 0.006885f
C720 B.n174 VSUBS 0.006885f
C721 B.n175 VSUBS 0.006885f
C722 B.n176 VSUBS 0.006885f
C723 B.n177 VSUBS 0.006885f
C724 B.n178 VSUBS 0.006885f
C725 B.n179 VSUBS 0.006885f
C726 B.n180 VSUBS 0.006885f
C727 B.n181 VSUBS 0.006885f
C728 B.n182 VSUBS 0.006885f
C729 B.n183 VSUBS 0.006885f
C730 B.n184 VSUBS 0.006885f
C731 B.n185 VSUBS 0.006885f
C732 B.n186 VSUBS 0.006885f
C733 B.n187 VSUBS 0.006885f
C734 B.n188 VSUBS 0.006885f
C735 B.n189 VSUBS 0.006885f
C736 B.n190 VSUBS 0.006885f
C737 B.n191 VSUBS 0.006885f
C738 B.n192 VSUBS 0.006885f
C739 B.n193 VSUBS 0.006885f
C740 B.n194 VSUBS 0.006885f
C741 B.n195 VSUBS 0.006885f
C742 B.n196 VSUBS 0.006885f
C743 B.n197 VSUBS 0.006885f
C744 B.n198 VSUBS 0.006885f
C745 B.n199 VSUBS 0.006885f
C746 B.n200 VSUBS 0.006885f
C747 B.n201 VSUBS 0.006885f
C748 B.n202 VSUBS 0.006885f
C749 B.n203 VSUBS 0.006885f
C750 B.n204 VSUBS 0.006885f
C751 B.n205 VSUBS 0.006885f
C752 B.n206 VSUBS 0.006885f
C753 B.n207 VSUBS 0.006885f
C754 B.n208 VSUBS 0.006885f
C755 B.n209 VSUBS 0.006885f
C756 B.n210 VSUBS 0.006885f
C757 B.n211 VSUBS 0.006885f
C758 B.n212 VSUBS 0.006885f
C759 B.n213 VSUBS 0.006885f
C760 B.n214 VSUBS 0.006885f
C761 B.n215 VSUBS 0.006885f
C762 B.n216 VSUBS 0.006885f
C763 B.n217 VSUBS 0.006885f
C764 B.n218 VSUBS 0.006885f
C765 B.n219 VSUBS 0.006885f
C766 B.n220 VSUBS 0.006885f
C767 B.n221 VSUBS 0.00648f
C768 B.n222 VSUBS 0.006885f
C769 B.n223 VSUBS 0.006885f
C770 B.n224 VSUBS 0.003848f
C771 B.n225 VSUBS 0.006885f
C772 B.n226 VSUBS 0.006885f
C773 B.n227 VSUBS 0.006885f
C774 B.n228 VSUBS 0.006885f
C775 B.n229 VSUBS 0.006885f
C776 B.n230 VSUBS 0.006885f
C777 B.n231 VSUBS 0.006885f
C778 B.n232 VSUBS 0.006885f
C779 B.n233 VSUBS 0.006885f
C780 B.n234 VSUBS 0.006885f
C781 B.n235 VSUBS 0.006885f
C782 B.n236 VSUBS 0.006885f
C783 B.n237 VSUBS 0.003848f
C784 B.n238 VSUBS 0.015953f
C785 B.n239 VSUBS 0.00648f
C786 B.n240 VSUBS 0.006885f
C787 B.n241 VSUBS 0.006885f
C788 B.n242 VSUBS 0.006885f
C789 B.n243 VSUBS 0.006885f
C790 B.n244 VSUBS 0.006885f
C791 B.n245 VSUBS 0.006885f
C792 B.n246 VSUBS 0.006885f
C793 B.n247 VSUBS 0.006885f
C794 B.n248 VSUBS 0.006885f
C795 B.n249 VSUBS 0.006885f
C796 B.n250 VSUBS 0.006885f
C797 B.n251 VSUBS 0.006885f
C798 B.n252 VSUBS 0.006885f
C799 B.n253 VSUBS 0.006885f
C800 B.n254 VSUBS 0.006885f
C801 B.n255 VSUBS 0.006885f
C802 B.n256 VSUBS 0.006885f
C803 B.n257 VSUBS 0.006885f
C804 B.n258 VSUBS 0.006885f
C805 B.n259 VSUBS 0.006885f
C806 B.n260 VSUBS 0.006885f
C807 B.n261 VSUBS 0.006885f
C808 B.n262 VSUBS 0.006885f
C809 B.n263 VSUBS 0.006885f
C810 B.n264 VSUBS 0.006885f
C811 B.n265 VSUBS 0.006885f
C812 B.n266 VSUBS 0.006885f
C813 B.n267 VSUBS 0.006885f
C814 B.n268 VSUBS 0.006885f
C815 B.n269 VSUBS 0.006885f
C816 B.n270 VSUBS 0.006885f
C817 B.n271 VSUBS 0.006885f
C818 B.n272 VSUBS 0.006885f
C819 B.n273 VSUBS 0.006885f
C820 B.n274 VSUBS 0.006885f
C821 B.n275 VSUBS 0.006885f
C822 B.n276 VSUBS 0.006885f
C823 B.n277 VSUBS 0.006885f
C824 B.n278 VSUBS 0.006885f
C825 B.n279 VSUBS 0.006885f
C826 B.n280 VSUBS 0.006885f
C827 B.n281 VSUBS 0.006885f
C828 B.n282 VSUBS 0.006885f
C829 B.n283 VSUBS 0.006885f
C830 B.n284 VSUBS 0.006885f
C831 B.n285 VSUBS 0.006885f
C832 B.n286 VSUBS 0.006885f
C833 B.n287 VSUBS 0.006885f
C834 B.n288 VSUBS 0.006885f
C835 B.n289 VSUBS 0.006885f
C836 B.n290 VSUBS 0.006885f
C837 B.n291 VSUBS 0.006885f
C838 B.n292 VSUBS 0.006885f
C839 B.n293 VSUBS 0.006885f
C840 B.n294 VSUBS 0.006885f
C841 B.n295 VSUBS 0.006885f
C842 B.n296 VSUBS 0.006885f
C843 B.n297 VSUBS 0.006885f
C844 B.n298 VSUBS 0.016546f
C845 B.n299 VSUBS 0.015653f
C846 B.n300 VSUBS 0.015653f
C847 B.n301 VSUBS 0.006885f
C848 B.n302 VSUBS 0.006885f
C849 B.n303 VSUBS 0.006885f
C850 B.n304 VSUBS 0.006885f
C851 B.n305 VSUBS 0.006885f
C852 B.n306 VSUBS 0.006885f
C853 B.n307 VSUBS 0.006885f
C854 B.n308 VSUBS 0.006885f
C855 B.n309 VSUBS 0.006885f
C856 B.n310 VSUBS 0.006885f
C857 B.n311 VSUBS 0.006885f
C858 B.n312 VSUBS 0.006885f
C859 B.n313 VSUBS 0.006885f
C860 B.n314 VSUBS 0.006885f
C861 B.n315 VSUBS 0.006885f
C862 B.n316 VSUBS 0.006885f
C863 B.n317 VSUBS 0.006885f
C864 B.n318 VSUBS 0.006885f
C865 B.n319 VSUBS 0.006885f
C866 B.n320 VSUBS 0.006885f
C867 B.n321 VSUBS 0.006885f
C868 B.n322 VSUBS 0.006885f
C869 B.n323 VSUBS 0.006885f
C870 B.n324 VSUBS 0.006885f
C871 B.n325 VSUBS 0.006885f
C872 B.n326 VSUBS 0.006885f
C873 B.n327 VSUBS 0.006885f
C874 B.n328 VSUBS 0.006885f
C875 B.n329 VSUBS 0.006885f
C876 B.n330 VSUBS 0.006885f
C877 B.n331 VSUBS 0.006885f
C878 B.n332 VSUBS 0.006885f
C879 B.n333 VSUBS 0.006885f
C880 B.n334 VSUBS 0.006885f
C881 B.n335 VSUBS 0.006885f
C882 B.n336 VSUBS 0.006885f
C883 B.n337 VSUBS 0.006885f
C884 B.n338 VSUBS 0.006885f
C885 B.n339 VSUBS 0.006885f
C886 B.n340 VSUBS 0.006885f
C887 B.n341 VSUBS 0.006885f
C888 B.n342 VSUBS 0.006885f
C889 B.n343 VSUBS 0.006885f
C890 B.n344 VSUBS 0.006885f
C891 B.n345 VSUBS 0.006885f
C892 B.n346 VSUBS 0.006885f
C893 B.n347 VSUBS 0.006885f
C894 B.n348 VSUBS 0.006885f
C895 B.n349 VSUBS 0.006885f
C896 B.n350 VSUBS 0.006885f
C897 B.n351 VSUBS 0.006885f
C898 B.n352 VSUBS 0.006885f
C899 B.n353 VSUBS 0.016467f
C900 B.n354 VSUBS 0.015653f
C901 B.n355 VSUBS 0.016546f
C902 B.n356 VSUBS 0.006885f
C903 B.n357 VSUBS 0.006885f
C904 B.n358 VSUBS 0.006885f
C905 B.n359 VSUBS 0.006885f
C906 B.n360 VSUBS 0.006885f
C907 B.n361 VSUBS 0.006885f
C908 B.n362 VSUBS 0.006885f
C909 B.n363 VSUBS 0.006885f
C910 B.n364 VSUBS 0.006885f
C911 B.n365 VSUBS 0.006885f
C912 B.n366 VSUBS 0.006885f
C913 B.n367 VSUBS 0.006885f
C914 B.n368 VSUBS 0.006885f
C915 B.n369 VSUBS 0.006885f
C916 B.n370 VSUBS 0.006885f
C917 B.n371 VSUBS 0.006885f
C918 B.n372 VSUBS 0.006885f
C919 B.n373 VSUBS 0.006885f
C920 B.n374 VSUBS 0.006885f
C921 B.n375 VSUBS 0.006885f
C922 B.n376 VSUBS 0.006885f
C923 B.n377 VSUBS 0.006885f
C924 B.n378 VSUBS 0.006885f
C925 B.n379 VSUBS 0.006885f
C926 B.n380 VSUBS 0.006885f
C927 B.n381 VSUBS 0.006885f
C928 B.n382 VSUBS 0.006885f
C929 B.n383 VSUBS 0.006885f
C930 B.n384 VSUBS 0.006885f
C931 B.n385 VSUBS 0.006885f
C932 B.n386 VSUBS 0.006885f
C933 B.n387 VSUBS 0.006885f
C934 B.n388 VSUBS 0.006885f
C935 B.n389 VSUBS 0.006885f
C936 B.n390 VSUBS 0.006885f
C937 B.n391 VSUBS 0.006885f
C938 B.n392 VSUBS 0.006885f
C939 B.n393 VSUBS 0.006885f
C940 B.n394 VSUBS 0.006885f
C941 B.n395 VSUBS 0.006885f
C942 B.n396 VSUBS 0.006885f
C943 B.n397 VSUBS 0.006885f
C944 B.n398 VSUBS 0.006885f
C945 B.n399 VSUBS 0.006885f
C946 B.n400 VSUBS 0.006885f
C947 B.n401 VSUBS 0.006885f
C948 B.n402 VSUBS 0.006885f
C949 B.n403 VSUBS 0.006885f
C950 B.n404 VSUBS 0.006885f
C951 B.n405 VSUBS 0.006885f
C952 B.n406 VSUBS 0.006885f
C953 B.n407 VSUBS 0.006885f
C954 B.n408 VSUBS 0.006885f
C955 B.n409 VSUBS 0.006885f
C956 B.n410 VSUBS 0.006885f
C957 B.n411 VSUBS 0.006885f
C958 B.n412 VSUBS 0.006885f
C959 B.n413 VSUBS 0.00648f
C960 B.n414 VSUBS 0.006885f
C961 B.n415 VSUBS 0.006885f
C962 B.n416 VSUBS 0.003848f
C963 B.n417 VSUBS 0.006885f
C964 B.n418 VSUBS 0.006885f
C965 B.n419 VSUBS 0.006885f
C966 B.n420 VSUBS 0.006885f
C967 B.n421 VSUBS 0.006885f
C968 B.n422 VSUBS 0.006885f
C969 B.n423 VSUBS 0.006885f
C970 B.n424 VSUBS 0.006885f
C971 B.n425 VSUBS 0.006885f
C972 B.n426 VSUBS 0.006885f
C973 B.n427 VSUBS 0.006885f
C974 B.n428 VSUBS 0.006885f
C975 B.n429 VSUBS 0.003848f
C976 B.n430 VSUBS 0.015953f
C977 B.n431 VSUBS 0.00648f
C978 B.n432 VSUBS 0.006885f
C979 B.n433 VSUBS 0.006885f
C980 B.n434 VSUBS 0.006885f
C981 B.n435 VSUBS 0.006885f
C982 B.n436 VSUBS 0.006885f
C983 B.n437 VSUBS 0.006885f
C984 B.n438 VSUBS 0.006885f
C985 B.n439 VSUBS 0.006885f
C986 B.n440 VSUBS 0.006885f
C987 B.n441 VSUBS 0.006885f
C988 B.n442 VSUBS 0.006885f
C989 B.n443 VSUBS 0.006885f
C990 B.n444 VSUBS 0.006885f
C991 B.n445 VSUBS 0.006885f
C992 B.n446 VSUBS 0.006885f
C993 B.n447 VSUBS 0.006885f
C994 B.n448 VSUBS 0.006885f
C995 B.n449 VSUBS 0.006885f
C996 B.n450 VSUBS 0.006885f
C997 B.n451 VSUBS 0.006885f
C998 B.n452 VSUBS 0.006885f
C999 B.n453 VSUBS 0.006885f
C1000 B.n454 VSUBS 0.006885f
C1001 B.n455 VSUBS 0.006885f
C1002 B.n456 VSUBS 0.006885f
C1003 B.n457 VSUBS 0.006885f
C1004 B.n458 VSUBS 0.006885f
C1005 B.n459 VSUBS 0.006885f
C1006 B.n460 VSUBS 0.006885f
C1007 B.n461 VSUBS 0.006885f
C1008 B.n462 VSUBS 0.006885f
C1009 B.n463 VSUBS 0.006885f
C1010 B.n464 VSUBS 0.006885f
C1011 B.n465 VSUBS 0.006885f
C1012 B.n466 VSUBS 0.006885f
C1013 B.n467 VSUBS 0.006885f
C1014 B.n468 VSUBS 0.006885f
C1015 B.n469 VSUBS 0.006885f
C1016 B.n470 VSUBS 0.006885f
C1017 B.n471 VSUBS 0.006885f
C1018 B.n472 VSUBS 0.006885f
C1019 B.n473 VSUBS 0.006885f
C1020 B.n474 VSUBS 0.006885f
C1021 B.n475 VSUBS 0.006885f
C1022 B.n476 VSUBS 0.006885f
C1023 B.n477 VSUBS 0.006885f
C1024 B.n478 VSUBS 0.006885f
C1025 B.n479 VSUBS 0.006885f
C1026 B.n480 VSUBS 0.006885f
C1027 B.n481 VSUBS 0.006885f
C1028 B.n482 VSUBS 0.006885f
C1029 B.n483 VSUBS 0.006885f
C1030 B.n484 VSUBS 0.006885f
C1031 B.n485 VSUBS 0.006885f
C1032 B.n486 VSUBS 0.006885f
C1033 B.n487 VSUBS 0.006885f
C1034 B.n488 VSUBS 0.006885f
C1035 B.n489 VSUBS 0.006885f
C1036 B.n490 VSUBS 0.016546f
C1037 B.n491 VSUBS 0.015653f
C1038 B.n492 VSUBS 0.015653f
C1039 B.n493 VSUBS 0.006885f
C1040 B.n494 VSUBS 0.006885f
C1041 B.n495 VSUBS 0.006885f
C1042 B.n496 VSUBS 0.006885f
C1043 B.n497 VSUBS 0.006885f
C1044 B.n498 VSUBS 0.006885f
C1045 B.n499 VSUBS 0.006885f
C1046 B.n500 VSUBS 0.006885f
C1047 B.n501 VSUBS 0.006885f
C1048 B.n502 VSUBS 0.006885f
C1049 B.n503 VSUBS 0.006885f
C1050 B.n504 VSUBS 0.006885f
C1051 B.n505 VSUBS 0.006885f
C1052 B.n506 VSUBS 0.006885f
C1053 B.n507 VSUBS 0.006885f
C1054 B.n508 VSUBS 0.006885f
C1055 B.n509 VSUBS 0.006885f
C1056 B.n510 VSUBS 0.006885f
C1057 B.n511 VSUBS 0.006885f
C1058 B.n512 VSUBS 0.006885f
C1059 B.n513 VSUBS 0.006885f
C1060 B.n514 VSUBS 0.006885f
C1061 B.n515 VSUBS 0.006885f
C1062 B.n516 VSUBS 0.006885f
C1063 B.n517 VSUBS 0.006885f
C1064 B.n518 VSUBS 0.006885f
C1065 B.n519 VSUBS 0.015591f
.ends

