* NGSPICE file created from diff_pair_sample_1304.ext - technology: sky130A

.subckt diff_pair_sample_1304 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=1.07415 ps=6.84 w=6.51 l=3.81
X1 VTAIL.t14 VN.t1 VDD2.t3 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X2 VDD2.t2 VN.t2 VTAIL.t13 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=2.5389 ps=13.8 w=6.51 l=3.81
X3 VDD1.t7 VP.t0 VTAIL.t3 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X4 B.t11 B.t9 B.t10 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=0 ps=0 w=6.51 l=3.81
X5 VDD1.t6 VP.t1 VTAIL.t5 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=2.5389 ps=13.8 w=6.51 l=3.81
X6 VTAIL.t1 VP.t2 VDD1.t5 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=1.07415 ps=6.84 w=6.51 l=3.81
X7 B.t8 B.t6 B.t7 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=0 ps=0 w=6.51 l=3.81
X8 B.t5 B.t3 B.t4 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=0 ps=0 w=6.51 l=3.81
X9 VDD2.t1 VN.t3 VTAIL.t12 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=2.5389 ps=13.8 w=6.51 l=3.81
X10 VTAIL.t2 VP.t3 VDD1.t4 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=1.07415 ps=6.84 w=6.51 l=3.81
X11 VDD2.t6 VN.t4 VTAIL.t11 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X12 VTAIL.t10 VN.t5 VDD2.t5 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=1.07415 ps=6.84 w=6.51 l=3.81
X13 VDD1.t3 VP.t4 VTAIL.t0 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X14 VDD1.t2 VP.t5 VTAIL.t7 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=2.5389 ps=13.8 w=6.51 l=3.81
X15 B.t2 B.t0 B.t1 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=2.5389 pd=13.8 as=0 ps=0 w=6.51 l=3.81
X16 VDD2.t4 VN.t6 VTAIL.t9 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X17 VTAIL.t6 VP.t6 VDD1.t1 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X18 VTAIL.t8 VN.t7 VDD2.t7 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
X19 VTAIL.t4 VP.t7 VDD1.t0 w_n5110_n2270# sky130_fd_pr__pfet_01v8 ad=1.07415 pd=6.84 as=1.07415 ps=6.84 w=6.51 l=3.81
R0 VN.n71 VN.n37 161.3
R1 VN.n70 VN.n69 161.3
R2 VN.n68 VN.n38 161.3
R3 VN.n67 VN.n66 161.3
R4 VN.n65 VN.n39 161.3
R5 VN.n64 VN.n63 161.3
R6 VN.n62 VN.n40 161.3
R7 VN.n61 VN.n60 161.3
R8 VN.n58 VN.n41 161.3
R9 VN.n57 VN.n56 161.3
R10 VN.n55 VN.n42 161.3
R11 VN.n54 VN.n53 161.3
R12 VN.n52 VN.n43 161.3
R13 VN.n51 VN.n50 161.3
R14 VN.n49 VN.n44 161.3
R15 VN.n48 VN.n47 161.3
R16 VN.n34 VN.n0 161.3
R17 VN.n33 VN.n32 161.3
R18 VN.n31 VN.n1 161.3
R19 VN.n30 VN.n29 161.3
R20 VN.n28 VN.n2 161.3
R21 VN.n27 VN.n26 161.3
R22 VN.n25 VN.n3 161.3
R23 VN.n24 VN.n23 161.3
R24 VN.n21 VN.n4 161.3
R25 VN.n20 VN.n19 161.3
R26 VN.n18 VN.n5 161.3
R27 VN.n17 VN.n16 161.3
R28 VN.n15 VN.n6 161.3
R29 VN.n14 VN.n13 161.3
R30 VN.n12 VN.n7 161.3
R31 VN.n11 VN.n10 161.3
R32 VN.n8 VN.t5 73.3701
R33 VN.n45 VN.t3 73.3701
R34 VN.n36 VN.n35 59.6721
R35 VN.n73 VN.n72 59.6721
R36 VN.n9 VN.n8 59.407
R37 VN.n46 VN.n45 59.407
R38 VN.n16 VN.n15 56.5193
R39 VN.n53 VN.n52 56.5193
R40 VN VN.n73 52.6708
R41 VN.n29 VN.n28 51.1773
R42 VN.n66 VN.n65 51.1773
R43 VN.n9 VN.t6 41.1792
R44 VN.n22 VN.t1 41.1792
R45 VN.n35 VN.t2 41.1792
R46 VN.n46 VN.t7 41.1792
R47 VN.n59 VN.t4 41.1792
R48 VN.n72 VN.t0 41.1792
R49 VN.n29 VN.n1 29.8095
R50 VN.n66 VN.n38 29.8095
R51 VN.n10 VN.n7 24.4675
R52 VN.n14 VN.n7 24.4675
R53 VN.n15 VN.n14 24.4675
R54 VN.n16 VN.n5 24.4675
R55 VN.n20 VN.n5 24.4675
R56 VN.n21 VN.n20 24.4675
R57 VN.n23 VN.n3 24.4675
R58 VN.n27 VN.n3 24.4675
R59 VN.n28 VN.n27 24.4675
R60 VN.n33 VN.n1 24.4675
R61 VN.n34 VN.n33 24.4675
R62 VN.n52 VN.n51 24.4675
R63 VN.n51 VN.n44 24.4675
R64 VN.n47 VN.n44 24.4675
R65 VN.n65 VN.n64 24.4675
R66 VN.n64 VN.n40 24.4675
R67 VN.n60 VN.n40 24.4675
R68 VN.n58 VN.n57 24.4675
R69 VN.n57 VN.n42 24.4675
R70 VN.n53 VN.n42 24.4675
R71 VN.n71 VN.n70 24.4675
R72 VN.n70 VN.n38 24.4675
R73 VN.n35 VN.n34 22.5101
R74 VN.n72 VN.n71 22.5101
R75 VN.n10 VN.n9 15.6594
R76 VN.n22 VN.n21 15.6594
R77 VN.n47 VN.n46 15.6594
R78 VN.n59 VN.n58 15.6594
R79 VN.n23 VN.n22 8.80862
R80 VN.n60 VN.n59 8.80862
R81 VN.n48 VN.n45 2.59964
R82 VN.n11 VN.n8 2.59964
R83 VN.n73 VN.n37 0.417535
R84 VN.n36 VN.n0 0.417535
R85 VN VN.n36 0.394291
R86 VN.n69 VN.n37 0.189894
R87 VN.n69 VN.n68 0.189894
R88 VN.n68 VN.n67 0.189894
R89 VN.n67 VN.n39 0.189894
R90 VN.n63 VN.n39 0.189894
R91 VN.n63 VN.n62 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n41 0.189894
R94 VN.n56 VN.n41 0.189894
R95 VN.n56 VN.n55 0.189894
R96 VN.n55 VN.n54 0.189894
R97 VN.n54 VN.n43 0.189894
R98 VN.n50 VN.n43 0.189894
R99 VN.n50 VN.n49 0.189894
R100 VN.n49 VN.n48 0.189894
R101 VN.n12 VN.n11 0.189894
R102 VN.n13 VN.n12 0.189894
R103 VN.n13 VN.n6 0.189894
R104 VN.n17 VN.n6 0.189894
R105 VN.n18 VN.n17 0.189894
R106 VN.n19 VN.n18 0.189894
R107 VN.n19 VN.n4 0.189894
R108 VN.n24 VN.n4 0.189894
R109 VN.n25 VN.n24 0.189894
R110 VN.n26 VN.n25 0.189894
R111 VN.n26 VN.n2 0.189894
R112 VN.n30 VN.n2 0.189894
R113 VN.n31 VN.n30 0.189894
R114 VN.n32 VN.n31 0.189894
R115 VN.n32 VN.n0 0.189894
R116 VDD2.n2 VDD2.n1 92.4935
R117 VDD2.n2 VDD2.n0 92.4935
R118 VDD2 VDD2.n5 92.4905
R119 VDD2.n4 VDD2.n3 90.7653
R120 VDD2.n4 VDD2.n2 45.3877
R121 VDD2.n5 VDD2.t7 4.99359
R122 VDD2.n5 VDD2.t1 4.99359
R123 VDD2.n3 VDD2.t0 4.99359
R124 VDD2.n3 VDD2.t6 4.99359
R125 VDD2.n1 VDD2.t3 4.99359
R126 VDD2.n1 VDD2.t2 4.99359
R127 VDD2.n0 VDD2.t5 4.99359
R128 VDD2.n0 VDD2.t4 4.99359
R129 VDD2 VDD2.n4 1.84317
R130 VTAIL.n278 VTAIL.n277 756.745
R131 VTAIL.n34 VTAIL.n33 756.745
R132 VTAIL.n68 VTAIL.n67 756.745
R133 VTAIL.n104 VTAIL.n103 756.745
R134 VTAIL.n244 VTAIL.n243 756.745
R135 VTAIL.n208 VTAIL.n207 756.745
R136 VTAIL.n174 VTAIL.n173 756.745
R137 VTAIL.n138 VTAIL.n137 756.745
R138 VTAIL.n256 VTAIL.n255 585
R139 VTAIL.n261 VTAIL.n260 585
R140 VTAIL.n263 VTAIL.n262 585
R141 VTAIL.n252 VTAIL.n251 585
R142 VTAIL.n269 VTAIL.n268 585
R143 VTAIL.n271 VTAIL.n270 585
R144 VTAIL.n248 VTAIL.n247 585
R145 VTAIL.n277 VTAIL.n276 585
R146 VTAIL.n12 VTAIL.n11 585
R147 VTAIL.n17 VTAIL.n16 585
R148 VTAIL.n19 VTAIL.n18 585
R149 VTAIL.n8 VTAIL.n7 585
R150 VTAIL.n25 VTAIL.n24 585
R151 VTAIL.n27 VTAIL.n26 585
R152 VTAIL.n4 VTAIL.n3 585
R153 VTAIL.n33 VTAIL.n32 585
R154 VTAIL.n46 VTAIL.n45 585
R155 VTAIL.n51 VTAIL.n50 585
R156 VTAIL.n53 VTAIL.n52 585
R157 VTAIL.n42 VTAIL.n41 585
R158 VTAIL.n59 VTAIL.n58 585
R159 VTAIL.n61 VTAIL.n60 585
R160 VTAIL.n38 VTAIL.n37 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n82 VTAIL.n81 585
R163 VTAIL.n87 VTAIL.n86 585
R164 VTAIL.n89 VTAIL.n88 585
R165 VTAIL.n78 VTAIL.n77 585
R166 VTAIL.n95 VTAIL.n94 585
R167 VTAIL.n97 VTAIL.n96 585
R168 VTAIL.n74 VTAIL.n73 585
R169 VTAIL.n103 VTAIL.n102 585
R170 VTAIL.n243 VTAIL.n242 585
R171 VTAIL.n214 VTAIL.n213 585
R172 VTAIL.n237 VTAIL.n236 585
R173 VTAIL.n235 VTAIL.n234 585
R174 VTAIL.n218 VTAIL.n217 585
R175 VTAIL.n229 VTAIL.n228 585
R176 VTAIL.n227 VTAIL.n226 585
R177 VTAIL.n222 VTAIL.n221 585
R178 VTAIL.n207 VTAIL.n206 585
R179 VTAIL.n178 VTAIL.n177 585
R180 VTAIL.n201 VTAIL.n200 585
R181 VTAIL.n199 VTAIL.n198 585
R182 VTAIL.n182 VTAIL.n181 585
R183 VTAIL.n193 VTAIL.n192 585
R184 VTAIL.n191 VTAIL.n190 585
R185 VTAIL.n186 VTAIL.n185 585
R186 VTAIL.n173 VTAIL.n172 585
R187 VTAIL.n144 VTAIL.n143 585
R188 VTAIL.n167 VTAIL.n166 585
R189 VTAIL.n165 VTAIL.n164 585
R190 VTAIL.n148 VTAIL.n147 585
R191 VTAIL.n159 VTAIL.n158 585
R192 VTAIL.n157 VTAIL.n156 585
R193 VTAIL.n152 VTAIL.n151 585
R194 VTAIL.n137 VTAIL.n136 585
R195 VTAIL.n108 VTAIL.n107 585
R196 VTAIL.n131 VTAIL.n130 585
R197 VTAIL.n129 VTAIL.n128 585
R198 VTAIL.n112 VTAIL.n111 585
R199 VTAIL.n123 VTAIL.n122 585
R200 VTAIL.n121 VTAIL.n120 585
R201 VTAIL.n116 VTAIL.n115 585
R202 VTAIL.n257 VTAIL.t13 329.084
R203 VTAIL.n13 VTAIL.t10 329.084
R204 VTAIL.n47 VTAIL.t7 329.084
R205 VTAIL.n83 VTAIL.t2 329.084
R206 VTAIL.n223 VTAIL.t5 329.084
R207 VTAIL.n187 VTAIL.t1 329.084
R208 VTAIL.n153 VTAIL.t12 329.084
R209 VTAIL.n117 VTAIL.t15 329.084
R210 VTAIL.n261 VTAIL.n255 171.744
R211 VTAIL.n262 VTAIL.n261 171.744
R212 VTAIL.n262 VTAIL.n251 171.744
R213 VTAIL.n269 VTAIL.n251 171.744
R214 VTAIL.n270 VTAIL.n269 171.744
R215 VTAIL.n270 VTAIL.n247 171.744
R216 VTAIL.n277 VTAIL.n247 171.744
R217 VTAIL.n17 VTAIL.n11 171.744
R218 VTAIL.n18 VTAIL.n17 171.744
R219 VTAIL.n18 VTAIL.n7 171.744
R220 VTAIL.n25 VTAIL.n7 171.744
R221 VTAIL.n26 VTAIL.n25 171.744
R222 VTAIL.n26 VTAIL.n3 171.744
R223 VTAIL.n33 VTAIL.n3 171.744
R224 VTAIL.n51 VTAIL.n45 171.744
R225 VTAIL.n52 VTAIL.n51 171.744
R226 VTAIL.n52 VTAIL.n41 171.744
R227 VTAIL.n59 VTAIL.n41 171.744
R228 VTAIL.n60 VTAIL.n59 171.744
R229 VTAIL.n60 VTAIL.n37 171.744
R230 VTAIL.n67 VTAIL.n37 171.744
R231 VTAIL.n87 VTAIL.n81 171.744
R232 VTAIL.n88 VTAIL.n87 171.744
R233 VTAIL.n88 VTAIL.n77 171.744
R234 VTAIL.n95 VTAIL.n77 171.744
R235 VTAIL.n96 VTAIL.n95 171.744
R236 VTAIL.n96 VTAIL.n73 171.744
R237 VTAIL.n103 VTAIL.n73 171.744
R238 VTAIL.n243 VTAIL.n213 171.744
R239 VTAIL.n236 VTAIL.n213 171.744
R240 VTAIL.n236 VTAIL.n235 171.744
R241 VTAIL.n235 VTAIL.n217 171.744
R242 VTAIL.n228 VTAIL.n217 171.744
R243 VTAIL.n228 VTAIL.n227 171.744
R244 VTAIL.n227 VTAIL.n221 171.744
R245 VTAIL.n207 VTAIL.n177 171.744
R246 VTAIL.n200 VTAIL.n177 171.744
R247 VTAIL.n200 VTAIL.n199 171.744
R248 VTAIL.n199 VTAIL.n181 171.744
R249 VTAIL.n192 VTAIL.n181 171.744
R250 VTAIL.n192 VTAIL.n191 171.744
R251 VTAIL.n191 VTAIL.n185 171.744
R252 VTAIL.n173 VTAIL.n143 171.744
R253 VTAIL.n166 VTAIL.n143 171.744
R254 VTAIL.n166 VTAIL.n165 171.744
R255 VTAIL.n165 VTAIL.n147 171.744
R256 VTAIL.n158 VTAIL.n147 171.744
R257 VTAIL.n158 VTAIL.n157 171.744
R258 VTAIL.n157 VTAIL.n151 171.744
R259 VTAIL.n137 VTAIL.n107 171.744
R260 VTAIL.n130 VTAIL.n107 171.744
R261 VTAIL.n130 VTAIL.n129 171.744
R262 VTAIL.n129 VTAIL.n111 171.744
R263 VTAIL.n122 VTAIL.n111 171.744
R264 VTAIL.n122 VTAIL.n121 171.744
R265 VTAIL.n121 VTAIL.n115 171.744
R266 VTAIL.t13 VTAIL.n255 85.8723
R267 VTAIL.t10 VTAIL.n11 85.8723
R268 VTAIL.t7 VTAIL.n45 85.8723
R269 VTAIL.t2 VTAIL.n81 85.8723
R270 VTAIL.t5 VTAIL.n221 85.8723
R271 VTAIL.t1 VTAIL.n185 85.8723
R272 VTAIL.t12 VTAIL.n151 85.8723
R273 VTAIL.t15 VTAIL.n115 85.8723
R274 VTAIL.n211 VTAIL.n210 74.0865
R275 VTAIL.n141 VTAIL.n140 74.0865
R276 VTAIL.n1 VTAIL.n0 74.0855
R277 VTAIL.n71 VTAIL.n70 74.0855
R278 VTAIL.n279 VTAIL.n278 34.7066
R279 VTAIL.n35 VTAIL.n34 34.7066
R280 VTAIL.n69 VTAIL.n68 34.7066
R281 VTAIL.n105 VTAIL.n104 34.7066
R282 VTAIL.n245 VTAIL.n244 34.7066
R283 VTAIL.n209 VTAIL.n208 34.7066
R284 VTAIL.n175 VTAIL.n174 34.7066
R285 VTAIL.n139 VTAIL.n138 34.7066
R286 VTAIL.n279 VTAIL.n245 21.5479
R287 VTAIL.n139 VTAIL.n105 21.5479
R288 VTAIL.n276 VTAIL.n246 12.8005
R289 VTAIL.n32 VTAIL.n2 12.8005
R290 VTAIL.n66 VTAIL.n36 12.8005
R291 VTAIL.n102 VTAIL.n72 12.8005
R292 VTAIL.n242 VTAIL.n212 12.8005
R293 VTAIL.n206 VTAIL.n176 12.8005
R294 VTAIL.n172 VTAIL.n142 12.8005
R295 VTAIL.n136 VTAIL.n106 12.8005
R296 VTAIL.n275 VTAIL.n248 12.0247
R297 VTAIL.n31 VTAIL.n4 12.0247
R298 VTAIL.n65 VTAIL.n38 12.0247
R299 VTAIL.n101 VTAIL.n74 12.0247
R300 VTAIL.n241 VTAIL.n214 12.0247
R301 VTAIL.n205 VTAIL.n178 12.0247
R302 VTAIL.n171 VTAIL.n144 12.0247
R303 VTAIL.n135 VTAIL.n108 12.0247
R304 VTAIL.n272 VTAIL.n271 11.249
R305 VTAIL.n28 VTAIL.n27 11.249
R306 VTAIL.n62 VTAIL.n61 11.249
R307 VTAIL.n98 VTAIL.n97 11.249
R308 VTAIL.n238 VTAIL.n237 11.249
R309 VTAIL.n202 VTAIL.n201 11.249
R310 VTAIL.n168 VTAIL.n167 11.249
R311 VTAIL.n132 VTAIL.n131 11.249
R312 VTAIL.n257 VTAIL.n256 10.7233
R313 VTAIL.n13 VTAIL.n12 10.7233
R314 VTAIL.n47 VTAIL.n46 10.7233
R315 VTAIL.n83 VTAIL.n82 10.7233
R316 VTAIL.n223 VTAIL.n222 10.7233
R317 VTAIL.n187 VTAIL.n186 10.7233
R318 VTAIL.n153 VTAIL.n152 10.7233
R319 VTAIL.n117 VTAIL.n116 10.7233
R320 VTAIL.n268 VTAIL.n250 10.4732
R321 VTAIL.n24 VTAIL.n6 10.4732
R322 VTAIL.n58 VTAIL.n40 10.4732
R323 VTAIL.n94 VTAIL.n76 10.4732
R324 VTAIL.n234 VTAIL.n216 10.4732
R325 VTAIL.n198 VTAIL.n180 10.4732
R326 VTAIL.n164 VTAIL.n146 10.4732
R327 VTAIL.n128 VTAIL.n110 10.4732
R328 VTAIL.n267 VTAIL.n252 9.69747
R329 VTAIL.n23 VTAIL.n8 9.69747
R330 VTAIL.n57 VTAIL.n42 9.69747
R331 VTAIL.n93 VTAIL.n78 9.69747
R332 VTAIL.n233 VTAIL.n218 9.69747
R333 VTAIL.n197 VTAIL.n182 9.69747
R334 VTAIL.n163 VTAIL.n148 9.69747
R335 VTAIL.n127 VTAIL.n112 9.69747
R336 VTAIL.n274 VTAIL.n246 9.45567
R337 VTAIL.n30 VTAIL.n2 9.45567
R338 VTAIL.n64 VTAIL.n36 9.45567
R339 VTAIL.n100 VTAIL.n72 9.45567
R340 VTAIL.n240 VTAIL.n212 9.45567
R341 VTAIL.n204 VTAIL.n176 9.45567
R342 VTAIL.n170 VTAIL.n142 9.45567
R343 VTAIL.n134 VTAIL.n106 9.45567
R344 VTAIL.n259 VTAIL.n258 9.3005
R345 VTAIL.n254 VTAIL.n253 9.3005
R346 VTAIL.n265 VTAIL.n264 9.3005
R347 VTAIL.n267 VTAIL.n266 9.3005
R348 VTAIL.n250 VTAIL.n249 9.3005
R349 VTAIL.n273 VTAIL.n272 9.3005
R350 VTAIL.n275 VTAIL.n274 9.3005
R351 VTAIL.n15 VTAIL.n14 9.3005
R352 VTAIL.n10 VTAIL.n9 9.3005
R353 VTAIL.n21 VTAIL.n20 9.3005
R354 VTAIL.n23 VTAIL.n22 9.3005
R355 VTAIL.n6 VTAIL.n5 9.3005
R356 VTAIL.n29 VTAIL.n28 9.3005
R357 VTAIL.n31 VTAIL.n30 9.3005
R358 VTAIL.n49 VTAIL.n48 9.3005
R359 VTAIL.n44 VTAIL.n43 9.3005
R360 VTAIL.n55 VTAIL.n54 9.3005
R361 VTAIL.n57 VTAIL.n56 9.3005
R362 VTAIL.n40 VTAIL.n39 9.3005
R363 VTAIL.n63 VTAIL.n62 9.3005
R364 VTAIL.n65 VTAIL.n64 9.3005
R365 VTAIL.n85 VTAIL.n84 9.3005
R366 VTAIL.n80 VTAIL.n79 9.3005
R367 VTAIL.n91 VTAIL.n90 9.3005
R368 VTAIL.n93 VTAIL.n92 9.3005
R369 VTAIL.n76 VTAIL.n75 9.3005
R370 VTAIL.n99 VTAIL.n98 9.3005
R371 VTAIL.n101 VTAIL.n100 9.3005
R372 VTAIL.n241 VTAIL.n240 9.3005
R373 VTAIL.n239 VTAIL.n238 9.3005
R374 VTAIL.n216 VTAIL.n215 9.3005
R375 VTAIL.n233 VTAIL.n232 9.3005
R376 VTAIL.n231 VTAIL.n230 9.3005
R377 VTAIL.n220 VTAIL.n219 9.3005
R378 VTAIL.n225 VTAIL.n224 9.3005
R379 VTAIL.n184 VTAIL.n183 9.3005
R380 VTAIL.n195 VTAIL.n194 9.3005
R381 VTAIL.n197 VTAIL.n196 9.3005
R382 VTAIL.n180 VTAIL.n179 9.3005
R383 VTAIL.n203 VTAIL.n202 9.3005
R384 VTAIL.n205 VTAIL.n204 9.3005
R385 VTAIL.n189 VTAIL.n188 9.3005
R386 VTAIL.n150 VTAIL.n149 9.3005
R387 VTAIL.n161 VTAIL.n160 9.3005
R388 VTAIL.n163 VTAIL.n162 9.3005
R389 VTAIL.n146 VTAIL.n145 9.3005
R390 VTAIL.n169 VTAIL.n168 9.3005
R391 VTAIL.n171 VTAIL.n170 9.3005
R392 VTAIL.n155 VTAIL.n154 9.3005
R393 VTAIL.n114 VTAIL.n113 9.3005
R394 VTAIL.n125 VTAIL.n124 9.3005
R395 VTAIL.n127 VTAIL.n126 9.3005
R396 VTAIL.n110 VTAIL.n109 9.3005
R397 VTAIL.n133 VTAIL.n132 9.3005
R398 VTAIL.n135 VTAIL.n134 9.3005
R399 VTAIL.n119 VTAIL.n118 9.3005
R400 VTAIL.n264 VTAIL.n263 8.92171
R401 VTAIL.n20 VTAIL.n19 8.92171
R402 VTAIL.n54 VTAIL.n53 8.92171
R403 VTAIL.n90 VTAIL.n89 8.92171
R404 VTAIL.n230 VTAIL.n229 8.92171
R405 VTAIL.n194 VTAIL.n193 8.92171
R406 VTAIL.n160 VTAIL.n159 8.92171
R407 VTAIL.n124 VTAIL.n123 8.92171
R408 VTAIL.n260 VTAIL.n254 8.14595
R409 VTAIL.n16 VTAIL.n10 8.14595
R410 VTAIL.n50 VTAIL.n44 8.14595
R411 VTAIL.n86 VTAIL.n80 8.14595
R412 VTAIL.n226 VTAIL.n220 8.14595
R413 VTAIL.n190 VTAIL.n184 8.14595
R414 VTAIL.n156 VTAIL.n150 8.14595
R415 VTAIL.n120 VTAIL.n114 8.14595
R416 VTAIL.n259 VTAIL.n256 7.3702
R417 VTAIL.n15 VTAIL.n12 7.3702
R418 VTAIL.n49 VTAIL.n46 7.3702
R419 VTAIL.n85 VTAIL.n82 7.3702
R420 VTAIL.n225 VTAIL.n222 7.3702
R421 VTAIL.n189 VTAIL.n186 7.3702
R422 VTAIL.n155 VTAIL.n152 7.3702
R423 VTAIL.n119 VTAIL.n116 7.3702
R424 VTAIL.n260 VTAIL.n259 5.81868
R425 VTAIL.n16 VTAIL.n15 5.81868
R426 VTAIL.n50 VTAIL.n49 5.81868
R427 VTAIL.n86 VTAIL.n85 5.81868
R428 VTAIL.n226 VTAIL.n225 5.81868
R429 VTAIL.n190 VTAIL.n189 5.81868
R430 VTAIL.n156 VTAIL.n155 5.81868
R431 VTAIL.n120 VTAIL.n119 5.81868
R432 VTAIL.n263 VTAIL.n254 5.04292
R433 VTAIL.n19 VTAIL.n10 5.04292
R434 VTAIL.n53 VTAIL.n44 5.04292
R435 VTAIL.n89 VTAIL.n80 5.04292
R436 VTAIL.n229 VTAIL.n220 5.04292
R437 VTAIL.n193 VTAIL.n184 5.04292
R438 VTAIL.n159 VTAIL.n150 5.04292
R439 VTAIL.n123 VTAIL.n114 5.04292
R440 VTAIL.n0 VTAIL.t9 4.99359
R441 VTAIL.n0 VTAIL.t14 4.99359
R442 VTAIL.n70 VTAIL.t3 4.99359
R443 VTAIL.n70 VTAIL.t6 4.99359
R444 VTAIL.n210 VTAIL.t0 4.99359
R445 VTAIL.n210 VTAIL.t4 4.99359
R446 VTAIL.n140 VTAIL.t11 4.99359
R447 VTAIL.n140 VTAIL.t8 4.99359
R448 VTAIL.n264 VTAIL.n252 4.26717
R449 VTAIL.n20 VTAIL.n8 4.26717
R450 VTAIL.n54 VTAIL.n42 4.26717
R451 VTAIL.n90 VTAIL.n78 4.26717
R452 VTAIL.n230 VTAIL.n218 4.26717
R453 VTAIL.n194 VTAIL.n182 4.26717
R454 VTAIL.n160 VTAIL.n148 4.26717
R455 VTAIL.n124 VTAIL.n112 4.26717
R456 VTAIL.n141 VTAIL.n139 3.56947
R457 VTAIL.n175 VTAIL.n141 3.56947
R458 VTAIL.n211 VTAIL.n209 3.56947
R459 VTAIL.n245 VTAIL.n211 3.56947
R460 VTAIL.n105 VTAIL.n71 3.56947
R461 VTAIL.n71 VTAIL.n69 3.56947
R462 VTAIL.n35 VTAIL.n1 3.56947
R463 VTAIL VTAIL.n279 3.51128
R464 VTAIL.n268 VTAIL.n267 3.49141
R465 VTAIL.n24 VTAIL.n23 3.49141
R466 VTAIL.n58 VTAIL.n57 3.49141
R467 VTAIL.n94 VTAIL.n93 3.49141
R468 VTAIL.n234 VTAIL.n233 3.49141
R469 VTAIL.n198 VTAIL.n197 3.49141
R470 VTAIL.n164 VTAIL.n163 3.49141
R471 VTAIL.n128 VTAIL.n127 3.49141
R472 VTAIL.n271 VTAIL.n250 2.71565
R473 VTAIL.n27 VTAIL.n6 2.71565
R474 VTAIL.n61 VTAIL.n40 2.71565
R475 VTAIL.n97 VTAIL.n76 2.71565
R476 VTAIL.n237 VTAIL.n216 2.71565
R477 VTAIL.n201 VTAIL.n180 2.71565
R478 VTAIL.n167 VTAIL.n146 2.71565
R479 VTAIL.n131 VTAIL.n110 2.71565
R480 VTAIL.n188 VTAIL.n187 2.41347
R481 VTAIL.n154 VTAIL.n153 2.41347
R482 VTAIL.n118 VTAIL.n117 2.41347
R483 VTAIL.n258 VTAIL.n257 2.41347
R484 VTAIL.n14 VTAIL.n13 2.41347
R485 VTAIL.n48 VTAIL.n47 2.41347
R486 VTAIL.n84 VTAIL.n83 2.41347
R487 VTAIL.n224 VTAIL.n223 2.41347
R488 VTAIL.n272 VTAIL.n248 1.93989
R489 VTAIL.n28 VTAIL.n4 1.93989
R490 VTAIL.n62 VTAIL.n38 1.93989
R491 VTAIL.n98 VTAIL.n74 1.93989
R492 VTAIL.n238 VTAIL.n214 1.93989
R493 VTAIL.n202 VTAIL.n178 1.93989
R494 VTAIL.n168 VTAIL.n144 1.93989
R495 VTAIL.n132 VTAIL.n108 1.93989
R496 VTAIL.n276 VTAIL.n275 1.16414
R497 VTAIL.n32 VTAIL.n31 1.16414
R498 VTAIL.n66 VTAIL.n65 1.16414
R499 VTAIL.n102 VTAIL.n101 1.16414
R500 VTAIL.n242 VTAIL.n241 1.16414
R501 VTAIL.n206 VTAIL.n205 1.16414
R502 VTAIL.n172 VTAIL.n171 1.16414
R503 VTAIL.n136 VTAIL.n135 1.16414
R504 VTAIL.n209 VTAIL.n175 0.470328
R505 VTAIL.n69 VTAIL.n35 0.470328
R506 VTAIL.n278 VTAIL.n246 0.388379
R507 VTAIL.n34 VTAIL.n2 0.388379
R508 VTAIL.n68 VTAIL.n36 0.388379
R509 VTAIL.n104 VTAIL.n72 0.388379
R510 VTAIL.n244 VTAIL.n212 0.388379
R511 VTAIL.n208 VTAIL.n176 0.388379
R512 VTAIL.n174 VTAIL.n142 0.388379
R513 VTAIL.n138 VTAIL.n106 0.388379
R514 VTAIL.n258 VTAIL.n253 0.155672
R515 VTAIL.n265 VTAIL.n253 0.155672
R516 VTAIL.n266 VTAIL.n265 0.155672
R517 VTAIL.n266 VTAIL.n249 0.155672
R518 VTAIL.n273 VTAIL.n249 0.155672
R519 VTAIL.n274 VTAIL.n273 0.155672
R520 VTAIL.n14 VTAIL.n9 0.155672
R521 VTAIL.n21 VTAIL.n9 0.155672
R522 VTAIL.n22 VTAIL.n21 0.155672
R523 VTAIL.n22 VTAIL.n5 0.155672
R524 VTAIL.n29 VTAIL.n5 0.155672
R525 VTAIL.n30 VTAIL.n29 0.155672
R526 VTAIL.n48 VTAIL.n43 0.155672
R527 VTAIL.n55 VTAIL.n43 0.155672
R528 VTAIL.n56 VTAIL.n55 0.155672
R529 VTAIL.n56 VTAIL.n39 0.155672
R530 VTAIL.n63 VTAIL.n39 0.155672
R531 VTAIL.n64 VTAIL.n63 0.155672
R532 VTAIL.n84 VTAIL.n79 0.155672
R533 VTAIL.n91 VTAIL.n79 0.155672
R534 VTAIL.n92 VTAIL.n91 0.155672
R535 VTAIL.n92 VTAIL.n75 0.155672
R536 VTAIL.n99 VTAIL.n75 0.155672
R537 VTAIL.n100 VTAIL.n99 0.155672
R538 VTAIL.n240 VTAIL.n239 0.155672
R539 VTAIL.n239 VTAIL.n215 0.155672
R540 VTAIL.n232 VTAIL.n215 0.155672
R541 VTAIL.n232 VTAIL.n231 0.155672
R542 VTAIL.n231 VTAIL.n219 0.155672
R543 VTAIL.n224 VTAIL.n219 0.155672
R544 VTAIL.n204 VTAIL.n203 0.155672
R545 VTAIL.n203 VTAIL.n179 0.155672
R546 VTAIL.n196 VTAIL.n179 0.155672
R547 VTAIL.n196 VTAIL.n195 0.155672
R548 VTAIL.n195 VTAIL.n183 0.155672
R549 VTAIL.n188 VTAIL.n183 0.155672
R550 VTAIL.n170 VTAIL.n169 0.155672
R551 VTAIL.n169 VTAIL.n145 0.155672
R552 VTAIL.n162 VTAIL.n145 0.155672
R553 VTAIL.n162 VTAIL.n161 0.155672
R554 VTAIL.n161 VTAIL.n149 0.155672
R555 VTAIL.n154 VTAIL.n149 0.155672
R556 VTAIL.n134 VTAIL.n133 0.155672
R557 VTAIL.n133 VTAIL.n109 0.155672
R558 VTAIL.n126 VTAIL.n109 0.155672
R559 VTAIL.n126 VTAIL.n125 0.155672
R560 VTAIL.n125 VTAIL.n113 0.155672
R561 VTAIL.n118 VTAIL.n113 0.155672
R562 VTAIL VTAIL.n1 0.0586897
R563 VP.n23 VP.n22 161.3
R564 VP.n24 VP.n19 161.3
R565 VP.n26 VP.n25 161.3
R566 VP.n27 VP.n18 161.3
R567 VP.n29 VP.n28 161.3
R568 VP.n30 VP.n17 161.3
R569 VP.n32 VP.n31 161.3
R570 VP.n33 VP.n16 161.3
R571 VP.n36 VP.n35 161.3
R572 VP.n37 VP.n15 161.3
R573 VP.n39 VP.n38 161.3
R574 VP.n40 VP.n14 161.3
R575 VP.n42 VP.n41 161.3
R576 VP.n43 VP.n13 161.3
R577 VP.n45 VP.n44 161.3
R578 VP.n46 VP.n12 161.3
R579 VP.n88 VP.n0 161.3
R580 VP.n87 VP.n86 161.3
R581 VP.n85 VP.n1 161.3
R582 VP.n84 VP.n83 161.3
R583 VP.n82 VP.n2 161.3
R584 VP.n81 VP.n80 161.3
R585 VP.n79 VP.n3 161.3
R586 VP.n78 VP.n77 161.3
R587 VP.n75 VP.n4 161.3
R588 VP.n74 VP.n73 161.3
R589 VP.n72 VP.n5 161.3
R590 VP.n71 VP.n70 161.3
R591 VP.n69 VP.n6 161.3
R592 VP.n68 VP.n67 161.3
R593 VP.n66 VP.n7 161.3
R594 VP.n65 VP.n64 161.3
R595 VP.n62 VP.n8 161.3
R596 VP.n61 VP.n60 161.3
R597 VP.n59 VP.n9 161.3
R598 VP.n58 VP.n57 161.3
R599 VP.n56 VP.n10 161.3
R600 VP.n55 VP.n54 161.3
R601 VP.n53 VP.n11 161.3
R602 VP.n52 VP.n51 161.3
R603 VP.n20 VP.t2 73.3697
R604 VP.n50 VP.n49 59.6721
R605 VP.n90 VP.n89 59.6721
R606 VP.n48 VP.n47 59.6721
R607 VP.n21 VP.n20 59.407
R608 VP.n70 VP.n69 56.5193
R609 VP.n28 VP.n27 56.5193
R610 VP.n49 VP.n48 52.6328
R611 VP.n57 VP.n56 51.1773
R612 VP.n83 VP.n82 51.1773
R613 VP.n41 VP.n40 51.1773
R614 VP.n50 VP.t3 41.1792
R615 VP.n63 VP.t0 41.1792
R616 VP.n76 VP.t6 41.1792
R617 VP.n89 VP.t5 41.1792
R618 VP.n47 VP.t1 41.1792
R619 VP.n34 VP.t7 41.1792
R620 VP.n21 VP.t4 41.1792
R621 VP.n56 VP.n55 29.8095
R622 VP.n83 VP.n1 29.8095
R623 VP.n41 VP.n13 29.8095
R624 VP.n51 VP.n11 24.4675
R625 VP.n55 VP.n11 24.4675
R626 VP.n57 VP.n9 24.4675
R627 VP.n61 VP.n9 24.4675
R628 VP.n62 VP.n61 24.4675
R629 VP.n64 VP.n7 24.4675
R630 VP.n68 VP.n7 24.4675
R631 VP.n69 VP.n68 24.4675
R632 VP.n70 VP.n5 24.4675
R633 VP.n74 VP.n5 24.4675
R634 VP.n75 VP.n74 24.4675
R635 VP.n77 VP.n3 24.4675
R636 VP.n81 VP.n3 24.4675
R637 VP.n82 VP.n81 24.4675
R638 VP.n87 VP.n1 24.4675
R639 VP.n88 VP.n87 24.4675
R640 VP.n45 VP.n13 24.4675
R641 VP.n46 VP.n45 24.4675
R642 VP.n28 VP.n17 24.4675
R643 VP.n32 VP.n17 24.4675
R644 VP.n33 VP.n32 24.4675
R645 VP.n35 VP.n15 24.4675
R646 VP.n39 VP.n15 24.4675
R647 VP.n40 VP.n39 24.4675
R648 VP.n22 VP.n19 24.4675
R649 VP.n26 VP.n19 24.4675
R650 VP.n27 VP.n26 24.4675
R651 VP.n51 VP.n50 22.5101
R652 VP.n89 VP.n88 22.5101
R653 VP.n47 VP.n46 22.5101
R654 VP.n64 VP.n63 15.6594
R655 VP.n76 VP.n75 15.6594
R656 VP.n34 VP.n33 15.6594
R657 VP.n22 VP.n21 15.6594
R658 VP.n63 VP.n62 8.80862
R659 VP.n77 VP.n76 8.80862
R660 VP.n35 VP.n34 8.80862
R661 VP.n23 VP.n20 2.59961
R662 VP.n48 VP.n12 0.417535
R663 VP.n52 VP.n49 0.417535
R664 VP.n90 VP.n0 0.417535
R665 VP VP.n90 0.394291
R666 VP.n24 VP.n23 0.189894
R667 VP.n25 VP.n24 0.189894
R668 VP.n25 VP.n18 0.189894
R669 VP.n29 VP.n18 0.189894
R670 VP.n30 VP.n29 0.189894
R671 VP.n31 VP.n30 0.189894
R672 VP.n31 VP.n16 0.189894
R673 VP.n36 VP.n16 0.189894
R674 VP.n37 VP.n36 0.189894
R675 VP.n38 VP.n37 0.189894
R676 VP.n38 VP.n14 0.189894
R677 VP.n42 VP.n14 0.189894
R678 VP.n43 VP.n42 0.189894
R679 VP.n44 VP.n43 0.189894
R680 VP.n44 VP.n12 0.189894
R681 VP.n53 VP.n52 0.189894
R682 VP.n54 VP.n53 0.189894
R683 VP.n54 VP.n10 0.189894
R684 VP.n58 VP.n10 0.189894
R685 VP.n59 VP.n58 0.189894
R686 VP.n60 VP.n59 0.189894
R687 VP.n60 VP.n8 0.189894
R688 VP.n65 VP.n8 0.189894
R689 VP.n66 VP.n65 0.189894
R690 VP.n67 VP.n66 0.189894
R691 VP.n67 VP.n6 0.189894
R692 VP.n71 VP.n6 0.189894
R693 VP.n72 VP.n71 0.189894
R694 VP.n73 VP.n72 0.189894
R695 VP.n73 VP.n4 0.189894
R696 VP.n78 VP.n4 0.189894
R697 VP.n79 VP.n78 0.189894
R698 VP.n80 VP.n79 0.189894
R699 VP.n80 VP.n2 0.189894
R700 VP.n84 VP.n2 0.189894
R701 VP.n85 VP.n84 0.189894
R702 VP.n86 VP.n85 0.189894
R703 VP.n86 VP.n0 0.189894
R704 VDD1 VDD1.n0 92.608
R705 VDD1.n3 VDD1.n2 92.4935
R706 VDD1.n3 VDD1.n1 92.4935
R707 VDD1.n5 VDD1.n4 90.7642
R708 VDD1.n5 VDD1.n3 45.9707
R709 VDD1.n4 VDD1.t0 4.99359
R710 VDD1.n4 VDD1.t6 4.99359
R711 VDD1.n0 VDD1.t5 4.99359
R712 VDD1.n0 VDD1.t3 4.99359
R713 VDD1.n2 VDD1.t1 4.99359
R714 VDD1.n2 VDD1.t2 4.99359
R715 VDD1.n1 VDD1.t4 4.99359
R716 VDD1.n1 VDD1.t7 4.99359
R717 VDD1 VDD1.n5 1.72679
R718 B.n612 B.n611 585
R719 B.n613 B.n70 585
R720 B.n615 B.n614 585
R721 B.n616 B.n69 585
R722 B.n618 B.n617 585
R723 B.n619 B.n68 585
R724 B.n621 B.n620 585
R725 B.n622 B.n67 585
R726 B.n624 B.n623 585
R727 B.n625 B.n66 585
R728 B.n627 B.n626 585
R729 B.n628 B.n65 585
R730 B.n630 B.n629 585
R731 B.n631 B.n64 585
R732 B.n633 B.n632 585
R733 B.n634 B.n63 585
R734 B.n636 B.n635 585
R735 B.n637 B.n62 585
R736 B.n639 B.n638 585
R737 B.n640 B.n61 585
R738 B.n642 B.n641 585
R739 B.n643 B.n60 585
R740 B.n645 B.n644 585
R741 B.n646 B.n59 585
R742 B.n648 B.n647 585
R743 B.n650 B.n649 585
R744 B.n651 B.n55 585
R745 B.n653 B.n652 585
R746 B.n654 B.n54 585
R747 B.n656 B.n655 585
R748 B.n657 B.n53 585
R749 B.n659 B.n658 585
R750 B.n660 B.n52 585
R751 B.n662 B.n661 585
R752 B.n663 B.n49 585
R753 B.n666 B.n665 585
R754 B.n667 B.n48 585
R755 B.n669 B.n668 585
R756 B.n670 B.n47 585
R757 B.n672 B.n671 585
R758 B.n673 B.n46 585
R759 B.n675 B.n674 585
R760 B.n676 B.n45 585
R761 B.n678 B.n677 585
R762 B.n679 B.n44 585
R763 B.n681 B.n680 585
R764 B.n682 B.n43 585
R765 B.n684 B.n683 585
R766 B.n685 B.n42 585
R767 B.n687 B.n686 585
R768 B.n688 B.n41 585
R769 B.n690 B.n689 585
R770 B.n691 B.n40 585
R771 B.n693 B.n692 585
R772 B.n694 B.n39 585
R773 B.n696 B.n695 585
R774 B.n697 B.n38 585
R775 B.n699 B.n698 585
R776 B.n700 B.n37 585
R777 B.n702 B.n701 585
R778 B.n610 B.n71 585
R779 B.n609 B.n608 585
R780 B.n607 B.n72 585
R781 B.n606 B.n605 585
R782 B.n604 B.n73 585
R783 B.n603 B.n602 585
R784 B.n601 B.n74 585
R785 B.n600 B.n599 585
R786 B.n598 B.n75 585
R787 B.n597 B.n596 585
R788 B.n595 B.n76 585
R789 B.n594 B.n593 585
R790 B.n592 B.n77 585
R791 B.n591 B.n590 585
R792 B.n589 B.n78 585
R793 B.n588 B.n587 585
R794 B.n586 B.n79 585
R795 B.n585 B.n584 585
R796 B.n583 B.n80 585
R797 B.n582 B.n581 585
R798 B.n580 B.n81 585
R799 B.n579 B.n578 585
R800 B.n577 B.n82 585
R801 B.n576 B.n575 585
R802 B.n574 B.n83 585
R803 B.n573 B.n572 585
R804 B.n571 B.n84 585
R805 B.n570 B.n569 585
R806 B.n568 B.n85 585
R807 B.n567 B.n566 585
R808 B.n565 B.n86 585
R809 B.n564 B.n563 585
R810 B.n562 B.n87 585
R811 B.n561 B.n560 585
R812 B.n559 B.n88 585
R813 B.n558 B.n557 585
R814 B.n556 B.n89 585
R815 B.n555 B.n554 585
R816 B.n553 B.n90 585
R817 B.n552 B.n551 585
R818 B.n550 B.n91 585
R819 B.n549 B.n548 585
R820 B.n547 B.n92 585
R821 B.n546 B.n545 585
R822 B.n544 B.n93 585
R823 B.n543 B.n542 585
R824 B.n541 B.n94 585
R825 B.n540 B.n539 585
R826 B.n538 B.n95 585
R827 B.n537 B.n536 585
R828 B.n535 B.n96 585
R829 B.n534 B.n533 585
R830 B.n532 B.n97 585
R831 B.n531 B.n530 585
R832 B.n529 B.n98 585
R833 B.n528 B.n527 585
R834 B.n526 B.n99 585
R835 B.n525 B.n524 585
R836 B.n523 B.n100 585
R837 B.n522 B.n521 585
R838 B.n520 B.n101 585
R839 B.n519 B.n518 585
R840 B.n517 B.n102 585
R841 B.n516 B.n515 585
R842 B.n514 B.n103 585
R843 B.n513 B.n512 585
R844 B.n511 B.n104 585
R845 B.n510 B.n509 585
R846 B.n508 B.n105 585
R847 B.n507 B.n506 585
R848 B.n505 B.n106 585
R849 B.n504 B.n503 585
R850 B.n502 B.n107 585
R851 B.n501 B.n500 585
R852 B.n499 B.n108 585
R853 B.n498 B.n497 585
R854 B.n496 B.n109 585
R855 B.n495 B.n494 585
R856 B.n493 B.n110 585
R857 B.n492 B.n491 585
R858 B.n490 B.n111 585
R859 B.n489 B.n488 585
R860 B.n487 B.n112 585
R861 B.n486 B.n485 585
R862 B.n484 B.n113 585
R863 B.n483 B.n482 585
R864 B.n481 B.n114 585
R865 B.n480 B.n479 585
R866 B.n478 B.n115 585
R867 B.n477 B.n476 585
R868 B.n475 B.n116 585
R869 B.n474 B.n473 585
R870 B.n472 B.n117 585
R871 B.n471 B.n470 585
R872 B.n469 B.n118 585
R873 B.n468 B.n467 585
R874 B.n466 B.n119 585
R875 B.n465 B.n464 585
R876 B.n463 B.n120 585
R877 B.n462 B.n461 585
R878 B.n460 B.n121 585
R879 B.n459 B.n458 585
R880 B.n457 B.n122 585
R881 B.n456 B.n455 585
R882 B.n454 B.n123 585
R883 B.n453 B.n452 585
R884 B.n451 B.n124 585
R885 B.n450 B.n449 585
R886 B.n448 B.n125 585
R887 B.n447 B.n446 585
R888 B.n445 B.n126 585
R889 B.n444 B.n443 585
R890 B.n442 B.n127 585
R891 B.n441 B.n440 585
R892 B.n439 B.n128 585
R893 B.n438 B.n437 585
R894 B.n436 B.n129 585
R895 B.n435 B.n434 585
R896 B.n433 B.n130 585
R897 B.n432 B.n431 585
R898 B.n430 B.n131 585
R899 B.n429 B.n428 585
R900 B.n427 B.n132 585
R901 B.n426 B.n425 585
R902 B.n424 B.n133 585
R903 B.n423 B.n422 585
R904 B.n421 B.n134 585
R905 B.n420 B.n419 585
R906 B.n418 B.n135 585
R907 B.n417 B.n416 585
R908 B.n415 B.n136 585
R909 B.n414 B.n413 585
R910 B.n412 B.n137 585
R911 B.n411 B.n410 585
R912 B.n409 B.n138 585
R913 B.n408 B.n407 585
R914 B.n406 B.n139 585
R915 B.n405 B.n404 585
R916 B.n403 B.n140 585
R917 B.n312 B.n311 585
R918 B.n313 B.n174 585
R919 B.n315 B.n314 585
R920 B.n316 B.n173 585
R921 B.n318 B.n317 585
R922 B.n319 B.n172 585
R923 B.n321 B.n320 585
R924 B.n322 B.n171 585
R925 B.n324 B.n323 585
R926 B.n325 B.n170 585
R927 B.n327 B.n326 585
R928 B.n328 B.n169 585
R929 B.n330 B.n329 585
R930 B.n331 B.n168 585
R931 B.n333 B.n332 585
R932 B.n334 B.n167 585
R933 B.n336 B.n335 585
R934 B.n337 B.n166 585
R935 B.n339 B.n338 585
R936 B.n340 B.n165 585
R937 B.n342 B.n341 585
R938 B.n343 B.n164 585
R939 B.n345 B.n344 585
R940 B.n346 B.n163 585
R941 B.n348 B.n347 585
R942 B.n350 B.n349 585
R943 B.n351 B.n159 585
R944 B.n353 B.n352 585
R945 B.n354 B.n158 585
R946 B.n356 B.n355 585
R947 B.n357 B.n157 585
R948 B.n359 B.n358 585
R949 B.n360 B.n156 585
R950 B.n362 B.n361 585
R951 B.n363 B.n153 585
R952 B.n366 B.n365 585
R953 B.n367 B.n152 585
R954 B.n369 B.n368 585
R955 B.n370 B.n151 585
R956 B.n372 B.n371 585
R957 B.n373 B.n150 585
R958 B.n375 B.n374 585
R959 B.n376 B.n149 585
R960 B.n378 B.n377 585
R961 B.n379 B.n148 585
R962 B.n381 B.n380 585
R963 B.n382 B.n147 585
R964 B.n384 B.n383 585
R965 B.n385 B.n146 585
R966 B.n387 B.n386 585
R967 B.n388 B.n145 585
R968 B.n390 B.n389 585
R969 B.n391 B.n144 585
R970 B.n393 B.n392 585
R971 B.n394 B.n143 585
R972 B.n396 B.n395 585
R973 B.n397 B.n142 585
R974 B.n399 B.n398 585
R975 B.n400 B.n141 585
R976 B.n402 B.n401 585
R977 B.n310 B.n175 585
R978 B.n309 B.n308 585
R979 B.n307 B.n176 585
R980 B.n306 B.n305 585
R981 B.n304 B.n177 585
R982 B.n303 B.n302 585
R983 B.n301 B.n178 585
R984 B.n300 B.n299 585
R985 B.n298 B.n179 585
R986 B.n297 B.n296 585
R987 B.n295 B.n180 585
R988 B.n294 B.n293 585
R989 B.n292 B.n181 585
R990 B.n291 B.n290 585
R991 B.n289 B.n182 585
R992 B.n288 B.n287 585
R993 B.n286 B.n183 585
R994 B.n285 B.n284 585
R995 B.n283 B.n184 585
R996 B.n282 B.n281 585
R997 B.n280 B.n185 585
R998 B.n279 B.n278 585
R999 B.n277 B.n186 585
R1000 B.n276 B.n275 585
R1001 B.n274 B.n187 585
R1002 B.n273 B.n272 585
R1003 B.n271 B.n188 585
R1004 B.n270 B.n269 585
R1005 B.n268 B.n189 585
R1006 B.n267 B.n266 585
R1007 B.n265 B.n190 585
R1008 B.n264 B.n263 585
R1009 B.n262 B.n191 585
R1010 B.n261 B.n260 585
R1011 B.n259 B.n192 585
R1012 B.n258 B.n257 585
R1013 B.n256 B.n193 585
R1014 B.n255 B.n254 585
R1015 B.n253 B.n194 585
R1016 B.n252 B.n251 585
R1017 B.n250 B.n195 585
R1018 B.n249 B.n248 585
R1019 B.n247 B.n196 585
R1020 B.n246 B.n245 585
R1021 B.n244 B.n197 585
R1022 B.n243 B.n242 585
R1023 B.n241 B.n198 585
R1024 B.n240 B.n239 585
R1025 B.n238 B.n199 585
R1026 B.n237 B.n236 585
R1027 B.n235 B.n200 585
R1028 B.n234 B.n233 585
R1029 B.n232 B.n201 585
R1030 B.n231 B.n230 585
R1031 B.n229 B.n202 585
R1032 B.n228 B.n227 585
R1033 B.n226 B.n203 585
R1034 B.n225 B.n224 585
R1035 B.n223 B.n204 585
R1036 B.n222 B.n221 585
R1037 B.n220 B.n205 585
R1038 B.n219 B.n218 585
R1039 B.n217 B.n206 585
R1040 B.n216 B.n215 585
R1041 B.n214 B.n207 585
R1042 B.n213 B.n212 585
R1043 B.n211 B.n208 585
R1044 B.n210 B.n209 585
R1045 B.n2 B.n0 585
R1046 B.n805 B.n1 585
R1047 B.n804 B.n803 585
R1048 B.n802 B.n3 585
R1049 B.n801 B.n800 585
R1050 B.n799 B.n4 585
R1051 B.n798 B.n797 585
R1052 B.n796 B.n5 585
R1053 B.n795 B.n794 585
R1054 B.n793 B.n6 585
R1055 B.n792 B.n791 585
R1056 B.n790 B.n7 585
R1057 B.n789 B.n788 585
R1058 B.n787 B.n8 585
R1059 B.n786 B.n785 585
R1060 B.n784 B.n9 585
R1061 B.n783 B.n782 585
R1062 B.n781 B.n10 585
R1063 B.n780 B.n779 585
R1064 B.n778 B.n11 585
R1065 B.n777 B.n776 585
R1066 B.n775 B.n12 585
R1067 B.n774 B.n773 585
R1068 B.n772 B.n13 585
R1069 B.n771 B.n770 585
R1070 B.n769 B.n14 585
R1071 B.n768 B.n767 585
R1072 B.n766 B.n15 585
R1073 B.n765 B.n764 585
R1074 B.n763 B.n16 585
R1075 B.n762 B.n761 585
R1076 B.n760 B.n17 585
R1077 B.n759 B.n758 585
R1078 B.n757 B.n18 585
R1079 B.n756 B.n755 585
R1080 B.n754 B.n19 585
R1081 B.n753 B.n752 585
R1082 B.n751 B.n20 585
R1083 B.n750 B.n749 585
R1084 B.n748 B.n21 585
R1085 B.n747 B.n746 585
R1086 B.n745 B.n22 585
R1087 B.n744 B.n743 585
R1088 B.n742 B.n23 585
R1089 B.n741 B.n740 585
R1090 B.n739 B.n24 585
R1091 B.n738 B.n737 585
R1092 B.n736 B.n25 585
R1093 B.n735 B.n734 585
R1094 B.n733 B.n26 585
R1095 B.n732 B.n731 585
R1096 B.n730 B.n27 585
R1097 B.n729 B.n728 585
R1098 B.n727 B.n28 585
R1099 B.n726 B.n725 585
R1100 B.n724 B.n29 585
R1101 B.n723 B.n722 585
R1102 B.n721 B.n30 585
R1103 B.n720 B.n719 585
R1104 B.n718 B.n31 585
R1105 B.n717 B.n716 585
R1106 B.n715 B.n32 585
R1107 B.n714 B.n713 585
R1108 B.n712 B.n33 585
R1109 B.n711 B.n710 585
R1110 B.n709 B.n34 585
R1111 B.n708 B.n707 585
R1112 B.n706 B.n35 585
R1113 B.n705 B.n704 585
R1114 B.n703 B.n36 585
R1115 B.n807 B.n806 585
R1116 B.n312 B.n175 540.549
R1117 B.n703 B.n702 540.549
R1118 B.n403 B.n402 540.549
R1119 B.n612 B.n71 540.549
R1120 B.n154 B.t5 357.18
R1121 B.n56 B.t7 357.18
R1122 B.n160 B.t2 357.18
R1123 B.n50 B.t10 357.18
R1124 B.n155 B.t4 276.889
R1125 B.n57 B.t8 276.889
R1126 B.n161 B.t1 276.889
R1127 B.n51 B.t11 276.889
R1128 B.n154 B.t3 250.53
R1129 B.n160 B.t0 250.53
R1130 B.n50 B.t9 250.53
R1131 B.n56 B.t6 250.53
R1132 B.n308 B.n175 163.367
R1133 B.n308 B.n307 163.367
R1134 B.n307 B.n306 163.367
R1135 B.n306 B.n177 163.367
R1136 B.n302 B.n177 163.367
R1137 B.n302 B.n301 163.367
R1138 B.n301 B.n300 163.367
R1139 B.n300 B.n179 163.367
R1140 B.n296 B.n179 163.367
R1141 B.n296 B.n295 163.367
R1142 B.n295 B.n294 163.367
R1143 B.n294 B.n181 163.367
R1144 B.n290 B.n181 163.367
R1145 B.n290 B.n289 163.367
R1146 B.n289 B.n288 163.367
R1147 B.n288 B.n183 163.367
R1148 B.n284 B.n183 163.367
R1149 B.n284 B.n283 163.367
R1150 B.n283 B.n282 163.367
R1151 B.n282 B.n185 163.367
R1152 B.n278 B.n185 163.367
R1153 B.n278 B.n277 163.367
R1154 B.n277 B.n276 163.367
R1155 B.n276 B.n187 163.367
R1156 B.n272 B.n187 163.367
R1157 B.n272 B.n271 163.367
R1158 B.n271 B.n270 163.367
R1159 B.n270 B.n189 163.367
R1160 B.n266 B.n189 163.367
R1161 B.n266 B.n265 163.367
R1162 B.n265 B.n264 163.367
R1163 B.n264 B.n191 163.367
R1164 B.n260 B.n191 163.367
R1165 B.n260 B.n259 163.367
R1166 B.n259 B.n258 163.367
R1167 B.n258 B.n193 163.367
R1168 B.n254 B.n193 163.367
R1169 B.n254 B.n253 163.367
R1170 B.n253 B.n252 163.367
R1171 B.n252 B.n195 163.367
R1172 B.n248 B.n195 163.367
R1173 B.n248 B.n247 163.367
R1174 B.n247 B.n246 163.367
R1175 B.n246 B.n197 163.367
R1176 B.n242 B.n197 163.367
R1177 B.n242 B.n241 163.367
R1178 B.n241 B.n240 163.367
R1179 B.n240 B.n199 163.367
R1180 B.n236 B.n199 163.367
R1181 B.n236 B.n235 163.367
R1182 B.n235 B.n234 163.367
R1183 B.n234 B.n201 163.367
R1184 B.n230 B.n201 163.367
R1185 B.n230 B.n229 163.367
R1186 B.n229 B.n228 163.367
R1187 B.n228 B.n203 163.367
R1188 B.n224 B.n203 163.367
R1189 B.n224 B.n223 163.367
R1190 B.n223 B.n222 163.367
R1191 B.n222 B.n205 163.367
R1192 B.n218 B.n205 163.367
R1193 B.n218 B.n217 163.367
R1194 B.n217 B.n216 163.367
R1195 B.n216 B.n207 163.367
R1196 B.n212 B.n207 163.367
R1197 B.n212 B.n211 163.367
R1198 B.n211 B.n210 163.367
R1199 B.n210 B.n2 163.367
R1200 B.n806 B.n2 163.367
R1201 B.n806 B.n805 163.367
R1202 B.n805 B.n804 163.367
R1203 B.n804 B.n3 163.367
R1204 B.n800 B.n3 163.367
R1205 B.n800 B.n799 163.367
R1206 B.n799 B.n798 163.367
R1207 B.n798 B.n5 163.367
R1208 B.n794 B.n5 163.367
R1209 B.n794 B.n793 163.367
R1210 B.n793 B.n792 163.367
R1211 B.n792 B.n7 163.367
R1212 B.n788 B.n7 163.367
R1213 B.n788 B.n787 163.367
R1214 B.n787 B.n786 163.367
R1215 B.n786 B.n9 163.367
R1216 B.n782 B.n9 163.367
R1217 B.n782 B.n781 163.367
R1218 B.n781 B.n780 163.367
R1219 B.n780 B.n11 163.367
R1220 B.n776 B.n11 163.367
R1221 B.n776 B.n775 163.367
R1222 B.n775 B.n774 163.367
R1223 B.n774 B.n13 163.367
R1224 B.n770 B.n13 163.367
R1225 B.n770 B.n769 163.367
R1226 B.n769 B.n768 163.367
R1227 B.n768 B.n15 163.367
R1228 B.n764 B.n15 163.367
R1229 B.n764 B.n763 163.367
R1230 B.n763 B.n762 163.367
R1231 B.n762 B.n17 163.367
R1232 B.n758 B.n17 163.367
R1233 B.n758 B.n757 163.367
R1234 B.n757 B.n756 163.367
R1235 B.n756 B.n19 163.367
R1236 B.n752 B.n19 163.367
R1237 B.n752 B.n751 163.367
R1238 B.n751 B.n750 163.367
R1239 B.n750 B.n21 163.367
R1240 B.n746 B.n21 163.367
R1241 B.n746 B.n745 163.367
R1242 B.n745 B.n744 163.367
R1243 B.n744 B.n23 163.367
R1244 B.n740 B.n23 163.367
R1245 B.n740 B.n739 163.367
R1246 B.n739 B.n738 163.367
R1247 B.n738 B.n25 163.367
R1248 B.n734 B.n25 163.367
R1249 B.n734 B.n733 163.367
R1250 B.n733 B.n732 163.367
R1251 B.n732 B.n27 163.367
R1252 B.n728 B.n27 163.367
R1253 B.n728 B.n727 163.367
R1254 B.n727 B.n726 163.367
R1255 B.n726 B.n29 163.367
R1256 B.n722 B.n29 163.367
R1257 B.n722 B.n721 163.367
R1258 B.n721 B.n720 163.367
R1259 B.n720 B.n31 163.367
R1260 B.n716 B.n31 163.367
R1261 B.n716 B.n715 163.367
R1262 B.n715 B.n714 163.367
R1263 B.n714 B.n33 163.367
R1264 B.n710 B.n33 163.367
R1265 B.n710 B.n709 163.367
R1266 B.n709 B.n708 163.367
R1267 B.n708 B.n35 163.367
R1268 B.n704 B.n35 163.367
R1269 B.n704 B.n703 163.367
R1270 B.n313 B.n312 163.367
R1271 B.n314 B.n313 163.367
R1272 B.n314 B.n173 163.367
R1273 B.n318 B.n173 163.367
R1274 B.n319 B.n318 163.367
R1275 B.n320 B.n319 163.367
R1276 B.n320 B.n171 163.367
R1277 B.n324 B.n171 163.367
R1278 B.n325 B.n324 163.367
R1279 B.n326 B.n325 163.367
R1280 B.n326 B.n169 163.367
R1281 B.n330 B.n169 163.367
R1282 B.n331 B.n330 163.367
R1283 B.n332 B.n331 163.367
R1284 B.n332 B.n167 163.367
R1285 B.n336 B.n167 163.367
R1286 B.n337 B.n336 163.367
R1287 B.n338 B.n337 163.367
R1288 B.n338 B.n165 163.367
R1289 B.n342 B.n165 163.367
R1290 B.n343 B.n342 163.367
R1291 B.n344 B.n343 163.367
R1292 B.n344 B.n163 163.367
R1293 B.n348 B.n163 163.367
R1294 B.n349 B.n348 163.367
R1295 B.n349 B.n159 163.367
R1296 B.n353 B.n159 163.367
R1297 B.n354 B.n353 163.367
R1298 B.n355 B.n354 163.367
R1299 B.n355 B.n157 163.367
R1300 B.n359 B.n157 163.367
R1301 B.n360 B.n359 163.367
R1302 B.n361 B.n360 163.367
R1303 B.n361 B.n153 163.367
R1304 B.n366 B.n153 163.367
R1305 B.n367 B.n366 163.367
R1306 B.n368 B.n367 163.367
R1307 B.n368 B.n151 163.367
R1308 B.n372 B.n151 163.367
R1309 B.n373 B.n372 163.367
R1310 B.n374 B.n373 163.367
R1311 B.n374 B.n149 163.367
R1312 B.n378 B.n149 163.367
R1313 B.n379 B.n378 163.367
R1314 B.n380 B.n379 163.367
R1315 B.n380 B.n147 163.367
R1316 B.n384 B.n147 163.367
R1317 B.n385 B.n384 163.367
R1318 B.n386 B.n385 163.367
R1319 B.n386 B.n145 163.367
R1320 B.n390 B.n145 163.367
R1321 B.n391 B.n390 163.367
R1322 B.n392 B.n391 163.367
R1323 B.n392 B.n143 163.367
R1324 B.n396 B.n143 163.367
R1325 B.n397 B.n396 163.367
R1326 B.n398 B.n397 163.367
R1327 B.n398 B.n141 163.367
R1328 B.n402 B.n141 163.367
R1329 B.n404 B.n403 163.367
R1330 B.n404 B.n139 163.367
R1331 B.n408 B.n139 163.367
R1332 B.n409 B.n408 163.367
R1333 B.n410 B.n409 163.367
R1334 B.n410 B.n137 163.367
R1335 B.n414 B.n137 163.367
R1336 B.n415 B.n414 163.367
R1337 B.n416 B.n415 163.367
R1338 B.n416 B.n135 163.367
R1339 B.n420 B.n135 163.367
R1340 B.n421 B.n420 163.367
R1341 B.n422 B.n421 163.367
R1342 B.n422 B.n133 163.367
R1343 B.n426 B.n133 163.367
R1344 B.n427 B.n426 163.367
R1345 B.n428 B.n427 163.367
R1346 B.n428 B.n131 163.367
R1347 B.n432 B.n131 163.367
R1348 B.n433 B.n432 163.367
R1349 B.n434 B.n433 163.367
R1350 B.n434 B.n129 163.367
R1351 B.n438 B.n129 163.367
R1352 B.n439 B.n438 163.367
R1353 B.n440 B.n439 163.367
R1354 B.n440 B.n127 163.367
R1355 B.n444 B.n127 163.367
R1356 B.n445 B.n444 163.367
R1357 B.n446 B.n445 163.367
R1358 B.n446 B.n125 163.367
R1359 B.n450 B.n125 163.367
R1360 B.n451 B.n450 163.367
R1361 B.n452 B.n451 163.367
R1362 B.n452 B.n123 163.367
R1363 B.n456 B.n123 163.367
R1364 B.n457 B.n456 163.367
R1365 B.n458 B.n457 163.367
R1366 B.n458 B.n121 163.367
R1367 B.n462 B.n121 163.367
R1368 B.n463 B.n462 163.367
R1369 B.n464 B.n463 163.367
R1370 B.n464 B.n119 163.367
R1371 B.n468 B.n119 163.367
R1372 B.n469 B.n468 163.367
R1373 B.n470 B.n469 163.367
R1374 B.n470 B.n117 163.367
R1375 B.n474 B.n117 163.367
R1376 B.n475 B.n474 163.367
R1377 B.n476 B.n475 163.367
R1378 B.n476 B.n115 163.367
R1379 B.n480 B.n115 163.367
R1380 B.n481 B.n480 163.367
R1381 B.n482 B.n481 163.367
R1382 B.n482 B.n113 163.367
R1383 B.n486 B.n113 163.367
R1384 B.n487 B.n486 163.367
R1385 B.n488 B.n487 163.367
R1386 B.n488 B.n111 163.367
R1387 B.n492 B.n111 163.367
R1388 B.n493 B.n492 163.367
R1389 B.n494 B.n493 163.367
R1390 B.n494 B.n109 163.367
R1391 B.n498 B.n109 163.367
R1392 B.n499 B.n498 163.367
R1393 B.n500 B.n499 163.367
R1394 B.n500 B.n107 163.367
R1395 B.n504 B.n107 163.367
R1396 B.n505 B.n504 163.367
R1397 B.n506 B.n505 163.367
R1398 B.n506 B.n105 163.367
R1399 B.n510 B.n105 163.367
R1400 B.n511 B.n510 163.367
R1401 B.n512 B.n511 163.367
R1402 B.n512 B.n103 163.367
R1403 B.n516 B.n103 163.367
R1404 B.n517 B.n516 163.367
R1405 B.n518 B.n517 163.367
R1406 B.n518 B.n101 163.367
R1407 B.n522 B.n101 163.367
R1408 B.n523 B.n522 163.367
R1409 B.n524 B.n523 163.367
R1410 B.n524 B.n99 163.367
R1411 B.n528 B.n99 163.367
R1412 B.n529 B.n528 163.367
R1413 B.n530 B.n529 163.367
R1414 B.n530 B.n97 163.367
R1415 B.n534 B.n97 163.367
R1416 B.n535 B.n534 163.367
R1417 B.n536 B.n535 163.367
R1418 B.n536 B.n95 163.367
R1419 B.n540 B.n95 163.367
R1420 B.n541 B.n540 163.367
R1421 B.n542 B.n541 163.367
R1422 B.n542 B.n93 163.367
R1423 B.n546 B.n93 163.367
R1424 B.n547 B.n546 163.367
R1425 B.n548 B.n547 163.367
R1426 B.n548 B.n91 163.367
R1427 B.n552 B.n91 163.367
R1428 B.n553 B.n552 163.367
R1429 B.n554 B.n553 163.367
R1430 B.n554 B.n89 163.367
R1431 B.n558 B.n89 163.367
R1432 B.n559 B.n558 163.367
R1433 B.n560 B.n559 163.367
R1434 B.n560 B.n87 163.367
R1435 B.n564 B.n87 163.367
R1436 B.n565 B.n564 163.367
R1437 B.n566 B.n565 163.367
R1438 B.n566 B.n85 163.367
R1439 B.n570 B.n85 163.367
R1440 B.n571 B.n570 163.367
R1441 B.n572 B.n571 163.367
R1442 B.n572 B.n83 163.367
R1443 B.n576 B.n83 163.367
R1444 B.n577 B.n576 163.367
R1445 B.n578 B.n577 163.367
R1446 B.n578 B.n81 163.367
R1447 B.n582 B.n81 163.367
R1448 B.n583 B.n582 163.367
R1449 B.n584 B.n583 163.367
R1450 B.n584 B.n79 163.367
R1451 B.n588 B.n79 163.367
R1452 B.n589 B.n588 163.367
R1453 B.n590 B.n589 163.367
R1454 B.n590 B.n77 163.367
R1455 B.n594 B.n77 163.367
R1456 B.n595 B.n594 163.367
R1457 B.n596 B.n595 163.367
R1458 B.n596 B.n75 163.367
R1459 B.n600 B.n75 163.367
R1460 B.n601 B.n600 163.367
R1461 B.n602 B.n601 163.367
R1462 B.n602 B.n73 163.367
R1463 B.n606 B.n73 163.367
R1464 B.n607 B.n606 163.367
R1465 B.n608 B.n607 163.367
R1466 B.n608 B.n71 163.367
R1467 B.n702 B.n37 163.367
R1468 B.n698 B.n37 163.367
R1469 B.n698 B.n697 163.367
R1470 B.n697 B.n696 163.367
R1471 B.n696 B.n39 163.367
R1472 B.n692 B.n39 163.367
R1473 B.n692 B.n691 163.367
R1474 B.n691 B.n690 163.367
R1475 B.n690 B.n41 163.367
R1476 B.n686 B.n41 163.367
R1477 B.n686 B.n685 163.367
R1478 B.n685 B.n684 163.367
R1479 B.n684 B.n43 163.367
R1480 B.n680 B.n43 163.367
R1481 B.n680 B.n679 163.367
R1482 B.n679 B.n678 163.367
R1483 B.n678 B.n45 163.367
R1484 B.n674 B.n45 163.367
R1485 B.n674 B.n673 163.367
R1486 B.n673 B.n672 163.367
R1487 B.n672 B.n47 163.367
R1488 B.n668 B.n47 163.367
R1489 B.n668 B.n667 163.367
R1490 B.n667 B.n666 163.367
R1491 B.n666 B.n49 163.367
R1492 B.n661 B.n49 163.367
R1493 B.n661 B.n660 163.367
R1494 B.n660 B.n659 163.367
R1495 B.n659 B.n53 163.367
R1496 B.n655 B.n53 163.367
R1497 B.n655 B.n654 163.367
R1498 B.n654 B.n653 163.367
R1499 B.n653 B.n55 163.367
R1500 B.n649 B.n55 163.367
R1501 B.n649 B.n648 163.367
R1502 B.n648 B.n59 163.367
R1503 B.n644 B.n59 163.367
R1504 B.n644 B.n643 163.367
R1505 B.n643 B.n642 163.367
R1506 B.n642 B.n61 163.367
R1507 B.n638 B.n61 163.367
R1508 B.n638 B.n637 163.367
R1509 B.n637 B.n636 163.367
R1510 B.n636 B.n63 163.367
R1511 B.n632 B.n63 163.367
R1512 B.n632 B.n631 163.367
R1513 B.n631 B.n630 163.367
R1514 B.n630 B.n65 163.367
R1515 B.n626 B.n65 163.367
R1516 B.n626 B.n625 163.367
R1517 B.n625 B.n624 163.367
R1518 B.n624 B.n67 163.367
R1519 B.n620 B.n67 163.367
R1520 B.n620 B.n619 163.367
R1521 B.n619 B.n618 163.367
R1522 B.n618 B.n69 163.367
R1523 B.n614 B.n69 163.367
R1524 B.n614 B.n613 163.367
R1525 B.n613 B.n612 163.367
R1526 B.n155 B.n154 80.2914
R1527 B.n161 B.n160 80.2914
R1528 B.n51 B.n50 80.2914
R1529 B.n57 B.n56 80.2914
R1530 B.n364 B.n155 59.5399
R1531 B.n162 B.n161 59.5399
R1532 B.n664 B.n51 59.5399
R1533 B.n58 B.n57 59.5399
R1534 B.n701 B.n36 35.1225
R1535 B.n611 B.n610 35.1225
R1536 B.n401 B.n140 35.1225
R1537 B.n311 B.n310 35.1225
R1538 B B.n807 18.0485
R1539 B.n701 B.n700 10.6151
R1540 B.n700 B.n699 10.6151
R1541 B.n699 B.n38 10.6151
R1542 B.n695 B.n38 10.6151
R1543 B.n695 B.n694 10.6151
R1544 B.n694 B.n693 10.6151
R1545 B.n693 B.n40 10.6151
R1546 B.n689 B.n40 10.6151
R1547 B.n689 B.n688 10.6151
R1548 B.n688 B.n687 10.6151
R1549 B.n687 B.n42 10.6151
R1550 B.n683 B.n42 10.6151
R1551 B.n683 B.n682 10.6151
R1552 B.n682 B.n681 10.6151
R1553 B.n681 B.n44 10.6151
R1554 B.n677 B.n44 10.6151
R1555 B.n677 B.n676 10.6151
R1556 B.n676 B.n675 10.6151
R1557 B.n675 B.n46 10.6151
R1558 B.n671 B.n46 10.6151
R1559 B.n671 B.n670 10.6151
R1560 B.n670 B.n669 10.6151
R1561 B.n669 B.n48 10.6151
R1562 B.n665 B.n48 10.6151
R1563 B.n663 B.n662 10.6151
R1564 B.n662 B.n52 10.6151
R1565 B.n658 B.n52 10.6151
R1566 B.n658 B.n657 10.6151
R1567 B.n657 B.n656 10.6151
R1568 B.n656 B.n54 10.6151
R1569 B.n652 B.n54 10.6151
R1570 B.n652 B.n651 10.6151
R1571 B.n651 B.n650 10.6151
R1572 B.n647 B.n646 10.6151
R1573 B.n646 B.n645 10.6151
R1574 B.n645 B.n60 10.6151
R1575 B.n641 B.n60 10.6151
R1576 B.n641 B.n640 10.6151
R1577 B.n640 B.n639 10.6151
R1578 B.n639 B.n62 10.6151
R1579 B.n635 B.n62 10.6151
R1580 B.n635 B.n634 10.6151
R1581 B.n634 B.n633 10.6151
R1582 B.n633 B.n64 10.6151
R1583 B.n629 B.n64 10.6151
R1584 B.n629 B.n628 10.6151
R1585 B.n628 B.n627 10.6151
R1586 B.n627 B.n66 10.6151
R1587 B.n623 B.n66 10.6151
R1588 B.n623 B.n622 10.6151
R1589 B.n622 B.n621 10.6151
R1590 B.n621 B.n68 10.6151
R1591 B.n617 B.n68 10.6151
R1592 B.n617 B.n616 10.6151
R1593 B.n616 B.n615 10.6151
R1594 B.n615 B.n70 10.6151
R1595 B.n611 B.n70 10.6151
R1596 B.n405 B.n140 10.6151
R1597 B.n406 B.n405 10.6151
R1598 B.n407 B.n406 10.6151
R1599 B.n407 B.n138 10.6151
R1600 B.n411 B.n138 10.6151
R1601 B.n412 B.n411 10.6151
R1602 B.n413 B.n412 10.6151
R1603 B.n413 B.n136 10.6151
R1604 B.n417 B.n136 10.6151
R1605 B.n418 B.n417 10.6151
R1606 B.n419 B.n418 10.6151
R1607 B.n419 B.n134 10.6151
R1608 B.n423 B.n134 10.6151
R1609 B.n424 B.n423 10.6151
R1610 B.n425 B.n424 10.6151
R1611 B.n425 B.n132 10.6151
R1612 B.n429 B.n132 10.6151
R1613 B.n430 B.n429 10.6151
R1614 B.n431 B.n430 10.6151
R1615 B.n431 B.n130 10.6151
R1616 B.n435 B.n130 10.6151
R1617 B.n436 B.n435 10.6151
R1618 B.n437 B.n436 10.6151
R1619 B.n437 B.n128 10.6151
R1620 B.n441 B.n128 10.6151
R1621 B.n442 B.n441 10.6151
R1622 B.n443 B.n442 10.6151
R1623 B.n443 B.n126 10.6151
R1624 B.n447 B.n126 10.6151
R1625 B.n448 B.n447 10.6151
R1626 B.n449 B.n448 10.6151
R1627 B.n449 B.n124 10.6151
R1628 B.n453 B.n124 10.6151
R1629 B.n454 B.n453 10.6151
R1630 B.n455 B.n454 10.6151
R1631 B.n455 B.n122 10.6151
R1632 B.n459 B.n122 10.6151
R1633 B.n460 B.n459 10.6151
R1634 B.n461 B.n460 10.6151
R1635 B.n461 B.n120 10.6151
R1636 B.n465 B.n120 10.6151
R1637 B.n466 B.n465 10.6151
R1638 B.n467 B.n466 10.6151
R1639 B.n467 B.n118 10.6151
R1640 B.n471 B.n118 10.6151
R1641 B.n472 B.n471 10.6151
R1642 B.n473 B.n472 10.6151
R1643 B.n473 B.n116 10.6151
R1644 B.n477 B.n116 10.6151
R1645 B.n478 B.n477 10.6151
R1646 B.n479 B.n478 10.6151
R1647 B.n479 B.n114 10.6151
R1648 B.n483 B.n114 10.6151
R1649 B.n484 B.n483 10.6151
R1650 B.n485 B.n484 10.6151
R1651 B.n485 B.n112 10.6151
R1652 B.n489 B.n112 10.6151
R1653 B.n490 B.n489 10.6151
R1654 B.n491 B.n490 10.6151
R1655 B.n491 B.n110 10.6151
R1656 B.n495 B.n110 10.6151
R1657 B.n496 B.n495 10.6151
R1658 B.n497 B.n496 10.6151
R1659 B.n497 B.n108 10.6151
R1660 B.n501 B.n108 10.6151
R1661 B.n502 B.n501 10.6151
R1662 B.n503 B.n502 10.6151
R1663 B.n503 B.n106 10.6151
R1664 B.n507 B.n106 10.6151
R1665 B.n508 B.n507 10.6151
R1666 B.n509 B.n508 10.6151
R1667 B.n509 B.n104 10.6151
R1668 B.n513 B.n104 10.6151
R1669 B.n514 B.n513 10.6151
R1670 B.n515 B.n514 10.6151
R1671 B.n515 B.n102 10.6151
R1672 B.n519 B.n102 10.6151
R1673 B.n520 B.n519 10.6151
R1674 B.n521 B.n520 10.6151
R1675 B.n521 B.n100 10.6151
R1676 B.n525 B.n100 10.6151
R1677 B.n526 B.n525 10.6151
R1678 B.n527 B.n526 10.6151
R1679 B.n527 B.n98 10.6151
R1680 B.n531 B.n98 10.6151
R1681 B.n532 B.n531 10.6151
R1682 B.n533 B.n532 10.6151
R1683 B.n533 B.n96 10.6151
R1684 B.n537 B.n96 10.6151
R1685 B.n538 B.n537 10.6151
R1686 B.n539 B.n538 10.6151
R1687 B.n539 B.n94 10.6151
R1688 B.n543 B.n94 10.6151
R1689 B.n544 B.n543 10.6151
R1690 B.n545 B.n544 10.6151
R1691 B.n545 B.n92 10.6151
R1692 B.n549 B.n92 10.6151
R1693 B.n550 B.n549 10.6151
R1694 B.n551 B.n550 10.6151
R1695 B.n551 B.n90 10.6151
R1696 B.n555 B.n90 10.6151
R1697 B.n556 B.n555 10.6151
R1698 B.n557 B.n556 10.6151
R1699 B.n557 B.n88 10.6151
R1700 B.n561 B.n88 10.6151
R1701 B.n562 B.n561 10.6151
R1702 B.n563 B.n562 10.6151
R1703 B.n563 B.n86 10.6151
R1704 B.n567 B.n86 10.6151
R1705 B.n568 B.n567 10.6151
R1706 B.n569 B.n568 10.6151
R1707 B.n569 B.n84 10.6151
R1708 B.n573 B.n84 10.6151
R1709 B.n574 B.n573 10.6151
R1710 B.n575 B.n574 10.6151
R1711 B.n575 B.n82 10.6151
R1712 B.n579 B.n82 10.6151
R1713 B.n580 B.n579 10.6151
R1714 B.n581 B.n580 10.6151
R1715 B.n581 B.n80 10.6151
R1716 B.n585 B.n80 10.6151
R1717 B.n586 B.n585 10.6151
R1718 B.n587 B.n586 10.6151
R1719 B.n587 B.n78 10.6151
R1720 B.n591 B.n78 10.6151
R1721 B.n592 B.n591 10.6151
R1722 B.n593 B.n592 10.6151
R1723 B.n593 B.n76 10.6151
R1724 B.n597 B.n76 10.6151
R1725 B.n598 B.n597 10.6151
R1726 B.n599 B.n598 10.6151
R1727 B.n599 B.n74 10.6151
R1728 B.n603 B.n74 10.6151
R1729 B.n604 B.n603 10.6151
R1730 B.n605 B.n604 10.6151
R1731 B.n605 B.n72 10.6151
R1732 B.n609 B.n72 10.6151
R1733 B.n610 B.n609 10.6151
R1734 B.n311 B.n174 10.6151
R1735 B.n315 B.n174 10.6151
R1736 B.n316 B.n315 10.6151
R1737 B.n317 B.n316 10.6151
R1738 B.n317 B.n172 10.6151
R1739 B.n321 B.n172 10.6151
R1740 B.n322 B.n321 10.6151
R1741 B.n323 B.n322 10.6151
R1742 B.n323 B.n170 10.6151
R1743 B.n327 B.n170 10.6151
R1744 B.n328 B.n327 10.6151
R1745 B.n329 B.n328 10.6151
R1746 B.n329 B.n168 10.6151
R1747 B.n333 B.n168 10.6151
R1748 B.n334 B.n333 10.6151
R1749 B.n335 B.n334 10.6151
R1750 B.n335 B.n166 10.6151
R1751 B.n339 B.n166 10.6151
R1752 B.n340 B.n339 10.6151
R1753 B.n341 B.n340 10.6151
R1754 B.n341 B.n164 10.6151
R1755 B.n345 B.n164 10.6151
R1756 B.n346 B.n345 10.6151
R1757 B.n347 B.n346 10.6151
R1758 B.n351 B.n350 10.6151
R1759 B.n352 B.n351 10.6151
R1760 B.n352 B.n158 10.6151
R1761 B.n356 B.n158 10.6151
R1762 B.n357 B.n356 10.6151
R1763 B.n358 B.n357 10.6151
R1764 B.n358 B.n156 10.6151
R1765 B.n362 B.n156 10.6151
R1766 B.n363 B.n362 10.6151
R1767 B.n365 B.n152 10.6151
R1768 B.n369 B.n152 10.6151
R1769 B.n370 B.n369 10.6151
R1770 B.n371 B.n370 10.6151
R1771 B.n371 B.n150 10.6151
R1772 B.n375 B.n150 10.6151
R1773 B.n376 B.n375 10.6151
R1774 B.n377 B.n376 10.6151
R1775 B.n377 B.n148 10.6151
R1776 B.n381 B.n148 10.6151
R1777 B.n382 B.n381 10.6151
R1778 B.n383 B.n382 10.6151
R1779 B.n383 B.n146 10.6151
R1780 B.n387 B.n146 10.6151
R1781 B.n388 B.n387 10.6151
R1782 B.n389 B.n388 10.6151
R1783 B.n389 B.n144 10.6151
R1784 B.n393 B.n144 10.6151
R1785 B.n394 B.n393 10.6151
R1786 B.n395 B.n394 10.6151
R1787 B.n395 B.n142 10.6151
R1788 B.n399 B.n142 10.6151
R1789 B.n400 B.n399 10.6151
R1790 B.n401 B.n400 10.6151
R1791 B.n310 B.n309 10.6151
R1792 B.n309 B.n176 10.6151
R1793 B.n305 B.n176 10.6151
R1794 B.n305 B.n304 10.6151
R1795 B.n304 B.n303 10.6151
R1796 B.n303 B.n178 10.6151
R1797 B.n299 B.n178 10.6151
R1798 B.n299 B.n298 10.6151
R1799 B.n298 B.n297 10.6151
R1800 B.n297 B.n180 10.6151
R1801 B.n293 B.n180 10.6151
R1802 B.n293 B.n292 10.6151
R1803 B.n292 B.n291 10.6151
R1804 B.n291 B.n182 10.6151
R1805 B.n287 B.n182 10.6151
R1806 B.n287 B.n286 10.6151
R1807 B.n286 B.n285 10.6151
R1808 B.n285 B.n184 10.6151
R1809 B.n281 B.n184 10.6151
R1810 B.n281 B.n280 10.6151
R1811 B.n280 B.n279 10.6151
R1812 B.n279 B.n186 10.6151
R1813 B.n275 B.n186 10.6151
R1814 B.n275 B.n274 10.6151
R1815 B.n274 B.n273 10.6151
R1816 B.n273 B.n188 10.6151
R1817 B.n269 B.n188 10.6151
R1818 B.n269 B.n268 10.6151
R1819 B.n268 B.n267 10.6151
R1820 B.n267 B.n190 10.6151
R1821 B.n263 B.n190 10.6151
R1822 B.n263 B.n262 10.6151
R1823 B.n262 B.n261 10.6151
R1824 B.n261 B.n192 10.6151
R1825 B.n257 B.n192 10.6151
R1826 B.n257 B.n256 10.6151
R1827 B.n256 B.n255 10.6151
R1828 B.n255 B.n194 10.6151
R1829 B.n251 B.n194 10.6151
R1830 B.n251 B.n250 10.6151
R1831 B.n250 B.n249 10.6151
R1832 B.n249 B.n196 10.6151
R1833 B.n245 B.n196 10.6151
R1834 B.n245 B.n244 10.6151
R1835 B.n244 B.n243 10.6151
R1836 B.n243 B.n198 10.6151
R1837 B.n239 B.n198 10.6151
R1838 B.n239 B.n238 10.6151
R1839 B.n238 B.n237 10.6151
R1840 B.n237 B.n200 10.6151
R1841 B.n233 B.n200 10.6151
R1842 B.n233 B.n232 10.6151
R1843 B.n232 B.n231 10.6151
R1844 B.n231 B.n202 10.6151
R1845 B.n227 B.n202 10.6151
R1846 B.n227 B.n226 10.6151
R1847 B.n226 B.n225 10.6151
R1848 B.n225 B.n204 10.6151
R1849 B.n221 B.n204 10.6151
R1850 B.n221 B.n220 10.6151
R1851 B.n220 B.n219 10.6151
R1852 B.n219 B.n206 10.6151
R1853 B.n215 B.n206 10.6151
R1854 B.n215 B.n214 10.6151
R1855 B.n214 B.n213 10.6151
R1856 B.n213 B.n208 10.6151
R1857 B.n209 B.n208 10.6151
R1858 B.n209 B.n0 10.6151
R1859 B.n803 B.n1 10.6151
R1860 B.n803 B.n802 10.6151
R1861 B.n802 B.n801 10.6151
R1862 B.n801 B.n4 10.6151
R1863 B.n797 B.n4 10.6151
R1864 B.n797 B.n796 10.6151
R1865 B.n796 B.n795 10.6151
R1866 B.n795 B.n6 10.6151
R1867 B.n791 B.n6 10.6151
R1868 B.n791 B.n790 10.6151
R1869 B.n790 B.n789 10.6151
R1870 B.n789 B.n8 10.6151
R1871 B.n785 B.n8 10.6151
R1872 B.n785 B.n784 10.6151
R1873 B.n784 B.n783 10.6151
R1874 B.n783 B.n10 10.6151
R1875 B.n779 B.n10 10.6151
R1876 B.n779 B.n778 10.6151
R1877 B.n778 B.n777 10.6151
R1878 B.n777 B.n12 10.6151
R1879 B.n773 B.n12 10.6151
R1880 B.n773 B.n772 10.6151
R1881 B.n772 B.n771 10.6151
R1882 B.n771 B.n14 10.6151
R1883 B.n767 B.n14 10.6151
R1884 B.n767 B.n766 10.6151
R1885 B.n766 B.n765 10.6151
R1886 B.n765 B.n16 10.6151
R1887 B.n761 B.n16 10.6151
R1888 B.n761 B.n760 10.6151
R1889 B.n760 B.n759 10.6151
R1890 B.n759 B.n18 10.6151
R1891 B.n755 B.n18 10.6151
R1892 B.n755 B.n754 10.6151
R1893 B.n754 B.n753 10.6151
R1894 B.n753 B.n20 10.6151
R1895 B.n749 B.n20 10.6151
R1896 B.n749 B.n748 10.6151
R1897 B.n748 B.n747 10.6151
R1898 B.n747 B.n22 10.6151
R1899 B.n743 B.n22 10.6151
R1900 B.n743 B.n742 10.6151
R1901 B.n742 B.n741 10.6151
R1902 B.n741 B.n24 10.6151
R1903 B.n737 B.n24 10.6151
R1904 B.n737 B.n736 10.6151
R1905 B.n736 B.n735 10.6151
R1906 B.n735 B.n26 10.6151
R1907 B.n731 B.n26 10.6151
R1908 B.n731 B.n730 10.6151
R1909 B.n730 B.n729 10.6151
R1910 B.n729 B.n28 10.6151
R1911 B.n725 B.n28 10.6151
R1912 B.n725 B.n724 10.6151
R1913 B.n724 B.n723 10.6151
R1914 B.n723 B.n30 10.6151
R1915 B.n719 B.n30 10.6151
R1916 B.n719 B.n718 10.6151
R1917 B.n718 B.n717 10.6151
R1918 B.n717 B.n32 10.6151
R1919 B.n713 B.n32 10.6151
R1920 B.n713 B.n712 10.6151
R1921 B.n712 B.n711 10.6151
R1922 B.n711 B.n34 10.6151
R1923 B.n707 B.n34 10.6151
R1924 B.n707 B.n706 10.6151
R1925 B.n706 B.n705 10.6151
R1926 B.n705 B.n36 10.6151
R1927 B.n665 B.n664 9.36635
R1928 B.n647 B.n58 9.36635
R1929 B.n347 B.n162 9.36635
R1930 B.n365 B.n364 9.36635
R1931 B.n807 B.n0 2.81026
R1932 B.n807 B.n1 2.81026
R1933 B.n664 B.n663 1.24928
R1934 B.n650 B.n58 1.24928
R1935 B.n350 B.n162 1.24928
R1936 B.n364 B.n363 1.24928
C0 VTAIL w_n5110_n2270# 3.12753f
C1 w_n5110_n2270# VN 10.6468f
C2 VDD1 VDD2 2.40504f
C3 VP VDD2 0.648364f
C4 VDD1 VTAIL 7.09063f
C5 VDD1 VN 0.153851f
C6 VP VTAIL 6.55458f
C7 VDD1 w_n5110_n2270# 2.19481f
C8 VP VN 8.12994f
C9 VP w_n5110_n2270# 11.3138f
C10 VDD1 VP 5.73822f
C11 VDD2 B 2.00552f
C12 VTAIL B 3.56445f
C13 VN B 1.43899f
C14 w_n5110_n2270# B 10.4375f
C15 VTAIL VDD2 7.15316f
C16 VN VDD2 5.24572f
C17 VDD1 B 1.87143f
C18 w_n5110_n2270# VDD2 2.36028f
C19 VP B 2.56348f
C20 VTAIL VN 6.54047f
C21 VDD2 VSUBS 2.474257f
C22 VDD1 VSUBS 3.16451f
C23 VTAIL VSUBS 0.836469f
C24 VN VSUBS 8.148109f
C25 VP VSUBS 4.396927f
C26 B VSUBS 5.88997f
C27 w_n5110_n2270# VSUBS 0.144531p
C28 B.n0 VSUBS 0.006307f
C29 B.n1 VSUBS 0.006307f
C30 B.n2 VSUBS 0.009973f
C31 B.n3 VSUBS 0.009973f
C32 B.n4 VSUBS 0.009973f
C33 B.n5 VSUBS 0.009973f
C34 B.n6 VSUBS 0.009973f
C35 B.n7 VSUBS 0.009973f
C36 B.n8 VSUBS 0.009973f
C37 B.n9 VSUBS 0.009973f
C38 B.n10 VSUBS 0.009973f
C39 B.n11 VSUBS 0.009973f
C40 B.n12 VSUBS 0.009973f
C41 B.n13 VSUBS 0.009973f
C42 B.n14 VSUBS 0.009973f
C43 B.n15 VSUBS 0.009973f
C44 B.n16 VSUBS 0.009973f
C45 B.n17 VSUBS 0.009973f
C46 B.n18 VSUBS 0.009973f
C47 B.n19 VSUBS 0.009973f
C48 B.n20 VSUBS 0.009973f
C49 B.n21 VSUBS 0.009973f
C50 B.n22 VSUBS 0.009973f
C51 B.n23 VSUBS 0.009973f
C52 B.n24 VSUBS 0.009973f
C53 B.n25 VSUBS 0.009973f
C54 B.n26 VSUBS 0.009973f
C55 B.n27 VSUBS 0.009973f
C56 B.n28 VSUBS 0.009973f
C57 B.n29 VSUBS 0.009973f
C58 B.n30 VSUBS 0.009973f
C59 B.n31 VSUBS 0.009973f
C60 B.n32 VSUBS 0.009973f
C61 B.n33 VSUBS 0.009973f
C62 B.n34 VSUBS 0.009973f
C63 B.n35 VSUBS 0.009973f
C64 B.n36 VSUBS 0.024213f
C65 B.n37 VSUBS 0.009973f
C66 B.n38 VSUBS 0.009973f
C67 B.n39 VSUBS 0.009973f
C68 B.n40 VSUBS 0.009973f
C69 B.n41 VSUBS 0.009973f
C70 B.n42 VSUBS 0.009973f
C71 B.n43 VSUBS 0.009973f
C72 B.n44 VSUBS 0.009973f
C73 B.n45 VSUBS 0.009973f
C74 B.n46 VSUBS 0.009973f
C75 B.n47 VSUBS 0.009973f
C76 B.n48 VSUBS 0.009973f
C77 B.n49 VSUBS 0.009973f
C78 B.t11 VSUBS 0.139946f
C79 B.t10 VSUBS 0.191566f
C80 B.t9 VSUBS 1.69404f
C81 B.n50 VSUBS 0.315191f
C82 B.n51 VSUBS 0.243862f
C83 B.n52 VSUBS 0.009973f
C84 B.n53 VSUBS 0.009973f
C85 B.n54 VSUBS 0.009973f
C86 B.n55 VSUBS 0.009973f
C87 B.t8 VSUBS 0.139949f
C88 B.t7 VSUBS 0.191569f
C89 B.t6 VSUBS 1.69404f
C90 B.n56 VSUBS 0.315188f
C91 B.n57 VSUBS 0.243859f
C92 B.n58 VSUBS 0.023107f
C93 B.n59 VSUBS 0.009973f
C94 B.n60 VSUBS 0.009973f
C95 B.n61 VSUBS 0.009973f
C96 B.n62 VSUBS 0.009973f
C97 B.n63 VSUBS 0.009973f
C98 B.n64 VSUBS 0.009973f
C99 B.n65 VSUBS 0.009973f
C100 B.n66 VSUBS 0.009973f
C101 B.n67 VSUBS 0.009973f
C102 B.n68 VSUBS 0.009973f
C103 B.n69 VSUBS 0.009973f
C104 B.n70 VSUBS 0.009973f
C105 B.n71 VSUBS 0.024213f
C106 B.n72 VSUBS 0.009973f
C107 B.n73 VSUBS 0.009973f
C108 B.n74 VSUBS 0.009973f
C109 B.n75 VSUBS 0.009973f
C110 B.n76 VSUBS 0.009973f
C111 B.n77 VSUBS 0.009973f
C112 B.n78 VSUBS 0.009973f
C113 B.n79 VSUBS 0.009973f
C114 B.n80 VSUBS 0.009973f
C115 B.n81 VSUBS 0.009973f
C116 B.n82 VSUBS 0.009973f
C117 B.n83 VSUBS 0.009973f
C118 B.n84 VSUBS 0.009973f
C119 B.n85 VSUBS 0.009973f
C120 B.n86 VSUBS 0.009973f
C121 B.n87 VSUBS 0.009973f
C122 B.n88 VSUBS 0.009973f
C123 B.n89 VSUBS 0.009973f
C124 B.n90 VSUBS 0.009973f
C125 B.n91 VSUBS 0.009973f
C126 B.n92 VSUBS 0.009973f
C127 B.n93 VSUBS 0.009973f
C128 B.n94 VSUBS 0.009973f
C129 B.n95 VSUBS 0.009973f
C130 B.n96 VSUBS 0.009973f
C131 B.n97 VSUBS 0.009973f
C132 B.n98 VSUBS 0.009973f
C133 B.n99 VSUBS 0.009973f
C134 B.n100 VSUBS 0.009973f
C135 B.n101 VSUBS 0.009973f
C136 B.n102 VSUBS 0.009973f
C137 B.n103 VSUBS 0.009973f
C138 B.n104 VSUBS 0.009973f
C139 B.n105 VSUBS 0.009973f
C140 B.n106 VSUBS 0.009973f
C141 B.n107 VSUBS 0.009973f
C142 B.n108 VSUBS 0.009973f
C143 B.n109 VSUBS 0.009973f
C144 B.n110 VSUBS 0.009973f
C145 B.n111 VSUBS 0.009973f
C146 B.n112 VSUBS 0.009973f
C147 B.n113 VSUBS 0.009973f
C148 B.n114 VSUBS 0.009973f
C149 B.n115 VSUBS 0.009973f
C150 B.n116 VSUBS 0.009973f
C151 B.n117 VSUBS 0.009973f
C152 B.n118 VSUBS 0.009973f
C153 B.n119 VSUBS 0.009973f
C154 B.n120 VSUBS 0.009973f
C155 B.n121 VSUBS 0.009973f
C156 B.n122 VSUBS 0.009973f
C157 B.n123 VSUBS 0.009973f
C158 B.n124 VSUBS 0.009973f
C159 B.n125 VSUBS 0.009973f
C160 B.n126 VSUBS 0.009973f
C161 B.n127 VSUBS 0.009973f
C162 B.n128 VSUBS 0.009973f
C163 B.n129 VSUBS 0.009973f
C164 B.n130 VSUBS 0.009973f
C165 B.n131 VSUBS 0.009973f
C166 B.n132 VSUBS 0.009973f
C167 B.n133 VSUBS 0.009973f
C168 B.n134 VSUBS 0.009973f
C169 B.n135 VSUBS 0.009973f
C170 B.n136 VSUBS 0.009973f
C171 B.n137 VSUBS 0.009973f
C172 B.n138 VSUBS 0.009973f
C173 B.n139 VSUBS 0.009973f
C174 B.n140 VSUBS 0.024213f
C175 B.n141 VSUBS 0.009973f
C176 B.n142 VSUBS 0.009973f
C177 B.n143 VSUBS 0.009973f
C178 B.n144 VSUBS 0.009973f
C179 B.n145 VSUBS 0.009973f
C180 B.n146 VSUBS 0.009973f
C181 B.n147 VSUBS 0.009973f
C182 B.n148 VSUBS 0.009973f
C183 B.n149 VSUBS 0.009973f
C184 B.n150 VSUBS 0.009973f
C185 B.n151 VSUBS 0.009973f
C186 B.n152 VSUBS 0.009973f
C187 B.n153 VSUBS 0.009973f
C188 B.t4 VSUBS 0.139949f
C189 B.t5 VSUBS 0.191569f
C190 B.t3 VSUBS 1.69404f
C191 B.n154 VSUBS 0.315188f
C192 B.n155 VSUBS 0.243859f
C193 B.n156 VSUBS 0.009973f
C194 B.n157 VSUBS 0.009973f
C195 B.n158 VSUBS 0.009973f
C196 B.n159 VSUBS 0.009973f
C197 B.t1 VSUBS 0.139946f
C198 B.t2 VSUBS 0.191566f
C199 B.t0 VSUBS 1.69404f
C200 B.n160 VSUBS 0.315191f
C201 B.n161 VSUBS 0.243862f
C202 B.n162 VSUBS 0.023107f
C203 B.n163 VSUBS 0.009973f
C204 B.n164 VSUBS 0.009973f
C205 B.n165 VSUBS 0.009973f
C206 B.n166 VSUBS 0.009973f
C207 B.n167 VSUBS 0.009973f
C208 B.n168 VSUBS 0.009973f
C209 B.n169 VSUBS 0.009973f
C210 B.n170 VSUBS 0.009973f
C211 B.n171 VSUBS 0.009973f
C212 B.n172 VSUBS 0.009973f
C213 B.n173 VSUBS 0.009973f
C214 B.n174 VSUBS 0.009973f
C215 B.n175 VSUBS 0.024213f
C216 B.n176 VSUBS 0.009973f
C217 B.n177 VSUBS 0.009973f
C218 B.n178 VSUBS 0.009973f
C219 B.n179 VSUBS 0.009973f
C220 B.n180 VSUBS 0.009973f
C221 B.n181 VSUBS 0.009973f
C222 B.n182 VSUBS 0.009973f
C223 B.n183 VSUBS 0.009973f
C224 B.n184 VSUBS 0.009973f
C225 B.n185 VSUBS 0.009973f
C226 B.n186 VSUBS 0.009973f
C227 B.n187 VSUBS 0.009973f
C228 B.n188 VSUBS 0.009973f
C229 B.n189 VSUBS 0.009973f
C230 B.n190 VSUBS 0.009973f
C231 B.n191 VSUBS 0.009973f
C232 B.n192 VSUBS 0.009973f
C233 B.n193 VSUBS 0.009973f
C234 B.n194 VSUBS 0.009973f
C235 B.n195 VSUBS 0.009973f
C236 B.n196 VSUBS 0.009973f
C237 B.n197 VSUBS 0.009973f
C238 B.n198 VSUBS 0.009973f
C239 B.n199 VSUBS 0.009973f
C240 B.n200 VSUBS 0.009973f
C241 B.n201 VSUBS 0.009973f
C242 B.n202 VSUBS 0.009973f
C243 B.n203 VSUBS 0.009973f
C244 B.n204 VSUBS 0.009973f
C245 B.n205 VSUBS 0.009973f
C246 B.n206 VSUBS 0.009973f
C247 B.n207 VSUBS 0.009973f
C248 B.n208 VSUBS 0.009973f
C249 B.n209 VSUBS 0.009973f
C250 B.n210 VSUBS 0.009973f
C251 B.n211 VSUBS 0.009973f
C252 B.n212 VSUBS 0.009973f
C253 B.n213 VSUBS 0.009973f
C254 B.n214 VSUBS 0.009973f
C255 B.n215 VSUBS 0.009973f
C256 B.n216 VSUBS 0.009973f
C257 B.n217 VSUBS 0.009973f
C258 B.n218 VSUBS 0.009973f
C259 B.n219 VSUBS 0.009973f
C260 B.n220 VSUBS 0.009973f
C261 B.n221 VSUBS 0.009973f
C262 B.n222 VSUBS 0.009973f
C263 B.n223 VSUBS 0.009973f
C264 B.n224 VSUBS 0.009973f
C265 B.n225 VSUBS 0.009973f
C266 B.n226 VSUBS 0.009973f
C267 B.n227 VSUBS 0.009973f
C268 B.n228 VSUBS 0.009973f
C269 B.n229 VSUBS 0.009973f
C270 B.n230 VSUBS 0.009973f
C271 B.n231 VSUBS 0.009973f
C272 B.n232 VSUBS 0.009973f
C273 B.n233 VSUBS 0.009973f
C274 B.n234 VSUBS 0.009973f
C275 B.n235 VSUBS 0.009973f
C276 B.n236 VSUBS 0.009973f
C277 B.n237 VSUBS 0.009973f
C278 B.n238 VSUBS 0.009973f
C279 B.n239 VSUBS 0.009973f
C280 B.n240 VSUBS 0.009973f
C281 B.n241 VSUBS 0.009973f
C282 B.n242 VSUBS 0.009973f
C283 B.n243 VSUBS 0.009973f
C284 B.n244 VSUBS 0.009973f
C285 B.n245 VSUBS 0.009973f
C286 B.n246 VSUBS 0.009973f
C287 B.n247 VSUBS 0.009973f
C288 B.n248 VSUBS 0.009973f
C289 B.n249 VSUBS 0.009973f
C290 B.n250 VSUBS 0.009973f
C291 B.n251 VSUBS 0.009973f
C292 B.n252 VSUBS 0.009973f
C293 B.n253 VSUBS 0.009973f
C294 B.n254 VSUBS 0.009973f
C295 B.n255 VSUBS 0.009973f
C296 B.n256 VSUBS 0.009973f
C297 B.n257 VSUBS 0.009973f
C298 B.n258 VSUBS 0.009973f
C299 B.n259 VSUBS 0.009973f
C300 B.n260 VSUBS 0.009973f
C301 B.n261 VSUBS 0.009973f
C302 B.n262 VSUBS 0.009973f
C303 B.n263 VSUBS 0.009973f
C304 B.n264 VSUBS 0.009973f
C305 B.n265 VSUBS 0.009973f
C306 B.n266 VSUBS 0.009973f
C307 B.n267 VSUBS 0.009973f
C308 B.n268 VSUBS 0.009973f
C309 B.n269 VSUBS 0.009973f
C310 B.n270 VSUBS 0.009973f
C311 B.n271 VSUBS 0.009973f
C312 B.n272 VSUBS 0.009973f
C313 B.n273 VSUBS 0.009973f
C314 B.n274 VSUBS 0.009973f
C315 B.n275 VSUBS 0.009973f
C316 B.n276 VSUBS 0.009973f
C317 B.n277 VSUBS 0.009973f
C318 B.n278 VSUBS 0.009973f
C319 B.n279 VSUBS 0.009973f
C320 B.n280 VSUBS 0.009973f
C321 B.n281 VSUBS 0.009973f
C322 B.n282 VSUBS 0.009973f
C323 B.n283 VSUBS 0.009973f
C324 B.n284 VSUBS 0.009973f
C325 B.n285 VSUBS 0.009973f
C326 B.n286 VSUBS 0.009973f
C327 B.n287 VSUBS 0.009973f
C328 B.n288 VSUBS 0.009973f
C329 B.n289 VSUBS 0.009973f
C330 B.n290 VSUBS 0.009973f
C331 B.n291 VSUBS 0.009973f
C332 B.n292 VSUBS 0.009973f
C333 B.n293 VSUBS 0.009973f
C334 B.n294 VSUBS 0.009973f
C335 B.n295 VSUBS 0.009973f
C336 B.n296 VSUBS 0.009973f
C337 B.n297 VSUBS 0.009973f
C338 B.n298 VSUBS 0.009973f
C339 B.n299 VSUBS 0.009973f
C340 B.n300 VSUBS 0.009973f
C341 B.n301 VSUBS 0.009973f
C342 B.n302 VSUBS 0.009973f
C343 B.n303 VSUBS 0.009973f
C344 B.n304 VSUBS 0.009973f
C345 B.n305 VSUBS 0.009973f
C346 B.n306 VSUBS 0.009973f
C347 B.n307 VSUBS 0.009973f
C348 B.n308 VSUBS 0.009973f
C349 B.n309 VSUBS 0.009973f
C350 B.n310 VSUBS 0.024213f
C351 B.n311 VSUBS 0.024774f
C352 B.n312 VSUBS 0.024774f
C353 B.n313 VSUBS 0.009973f
C354 B.n314 VSUBS 0.009973f
C355 B.n315 VSUBS 0.009973f
C356 B.n316 VSUBS 0.009973f
C357 B.n317 VSUBS 0.009973f
C358 B.n318 VSUBS 0.009973f
C359 B.n319 VSUBS 0.009973f
C360 B.n320 VSUBS 0.009973f
C361 B.n321 VSUBS 0.009973f
C362 B.n322 VSUBS 0.009973f
C363 B.n323 VSUBS 0.009973f
C364 B.n324 VSUBS 0.009973f
C365 B.n325 VSUBS 0.009973f
C366 B.n326 VSUBS 0.009973f
C367 B.n327 VSUBS 0.009973f
C368 B.n328 VSUBS 0.009973f
C369 B.n329 VSUBS 0.009973f
C370 B.n330 VSUBS 0.009973f
C371 B.n331 VSUBS 0.009973f
C372 B.n332 VSUBS 0.009973f
C373 B.n333 VSUBS 0.009973f
C374 B.n334 VSUBS 0.009973f
C375 B.n335 VSUBS 0.009973f
C376 B.n336 VSUBS 0.009973f
C377 B.n337 VSUBS 0.009973f
C378 B.n338 VSUBS 0.009973f
C379 B.n339 VSUBS 0.009973f
C380 B.n340 VSUBS 0.009973f
C381 B.n341 VSUBS 0.009973f
C382 B.n342 VSUBS 0.009973f
C383 B.n343 VSUBS 0.009973f
C384 B.n344 VSUBS 0.009973f
C385 B.n345 VSUBS 0.009973f
C386 B.n346 VSUBS 0.009973f
C387 B.n347 VSUBS 0.009387f
C388 B.n348 VSUBS 0.009973f
C389 B.n349 VSUBS 0.009973f
C390 B.n350 VSUBS 0.005573f
C391 B.n351 VSUBS 0.009973f
C392 B.n352 VSUBS 0.009973f
C393 B.n353 VSUBS 0.009973f
C394 B.n354 VSUBS 0.009973f
C395 B.n355 VSUBS 0.009973f
C396 B.n356 VSUBS 0.009973f
C397 B.n357 VSUBS 0.009973f
C398 B.n358 VSUBS 0.009973f
C399 B.n359 VSUBS 0.009973f
C400 B.n360 VSUBS 0.009973f
C401 B.n361 VSUBS 0.009973f
C402 B.n362 VSUBS 0.009973f
C403 B.n363 VSUBS 0.005573f
C404 B.n364 VSUBS 0.023107f
C405 B.n365 VSUBS 0.009387f
C406 B.n366 VSUBS 0.009973f
C407 B.n367 VSUBS 0.009973f
C408 B.n368 VSUBS 0.009973f
C409 B.n369 VSUBS 0.009973f
C410 B.n370 VSUBS 0.009973f
C411 B.n371 VSUBS 0.009973f
C412 B.n372 VSUBS 0.009973f
C413 B.n373 VSUBS 0.009973f
C414 B.n374 VSUBS 0.009973f
C415 B.n375 VSUBS 0.009973f
C416 B.n376 VSUBS 0.009973f
C417 B.n377 VSUBS 0.009973f
C418 B.n378 VSUBS 0.009973f
C419 B.n379 VSUBS 0.009973f
C420 B.n380 VSUBS 0.009973f
C421 B.n381 VSUBS 0.009973f
C422 B.n382 VSUBS 0.009973f
C423 B.n383 VSUBS 0.009973f
C424 B.n384 VSUBS 0.009973f
C425 B.n385 VSUBS 0.009973f
C426 B.n386 VSUBS 0.009973f
C427 B.n387 VSUBS 0.009973f
C428 B.n388 VSUBS 0.009973f
C429 B.n389 VSUBS 0.009973f
C430 B.n390 VSUBS 0.009973f
C431 B.n391 VSUBS 0.009973f
C432 B.n392 VSUBS 0.009973f
C433 B.n393 VSUBS 0.009973f
C434 B.n394 VSUBS 0.009973f
C435 B.n395 VSUBS 0.009973f
C436 B.n396 VSUBS 0.009973f
C437 B.n397 VSUBS 0.009973f
C438 B.n398 VSUBS 0.009973f
C439 B.n399 VSUBS 0.009973f
C440 B.n400 VSUBS 0.009973f
C441 B.n401 VSUBS 0.024774f
C442 B.n402 VSUBS 0.024774f
C443 B.n403 VSUBS 0.024213f
C444 B.n404 VSUBS 0.009973f
C445 B.n405 VSUBS 0.009973f
C446 B.n406 VSUBS 0.009973f
C447 B.n407 VSUBS 0.009973f
C448 B.n408 VSUBS 0.009973f
C449 B.n409 VSUBS 0.009973f
C450 B.n410 VSUBS 0.009973f
C451 B.n411 VSUBS 0.009973f
C452 B.n412 VSUBS 0.009973f
C453 B.n413 VSUBS 0.009973f
C454 B.n414 VSUBS 0.009973f
C455 B.n415 VSUBS 0.009973f
C456 B.n416 VSUBS 0.009973f
C457 B.n417 VSUBS 0.009973f
C458 B.n418 VSUBS 0.009973f
C459 B.n419 VSUBS 0.009973f
C460 B.n420 VSUBS 0.009973f
C461 B.n421 VSUBS 0.009973f
C462 B.n422 VSUBS 0.009973f
C463 B.n423 VSUBS 0.009973f
C464 B.n424 VSUBS 0.009973f
C465 B.n425 VSUBS 0.009973f
C466 B.n426 VSUBS 0.009973f
C467 B.n427 VSUBS 0.009973f
C468 B.n428 VSUBS 0.009973f
C469 B.n429 VSUBS 0.009973f
C470 B.n430 VSUBS 0.009973f
C471 B.n431 VSUBS 0.009973f
C472 B.n432 VSUBS 0.009973f
C473 B.n433 VSUBS 0.009973f
C474 B.n434 VSUBS 0.009973f
C475 B.n435 VSUBS 0.009973f
C476 B.n436 VSUBS 0.009973f
C477 B.n437 VSUBS 0.009973f
C478 B.n438 VSUBS 0.009973f
C479 B.n439 VSUBS 0.009973f
C480 B.n440 VSUBS 0.009973f
C481 B.n441 VSUBS 0.009973f
C482 B.n442 VSUBS 0.009973f
C483 B.n443 VSUBS 0.009973f
C484 B.n444 VSUBS 0.009973f
C485 B.n445 VSUBS 0.009973f
C486 B.n446 VSUBS 0.009973f
C487 B.n447 VSUBS 0.009973f
C488 B.n448 VSUBS 0.009973f
C489 B.n449 VSUBS 0.009973f
C490 B.n450 VSUBS 0.009973f
C491 B.n451 VSUBS 0.009973f
C492 B.n452 VSUBS 0.009973f
C493 B.n453 VSUBS 0.009973f
C494 B.n454 VSUBS 0.009973f
C495 B.n455 VSUBS 0.009973f
C496 B.n456 VSUBS 0.009973f
C497 B.n457 VSUBS 0.009973f
C498 B.n458 VSUBS 0.009973f
C499 B.n459 VSUBS 0.009973f
C500 B.n460 VSUBS 0.009973f
C501 B.n461 VSUBS 0.009973f
C502 B.n462 VSUBS 0.009973f
C503 B.n463 VSUBS 0.009973f
C504 B.n464 VSUBS 0.009973f
C505 B.n465 VSUBS 0.009973f
C506 B.n466 VSUBS 0.009973f
C507 B.n467 VSUBS 0.009973f
C508 B.n468 VSUBS 0.009973f
C509 B.n469 VSUBS 0.009973f
C510 B.n470 VSUBS 0.009973f
C511 B.n471 VSUBS 0.009973f
C512 B.n472 VSUBS 0.009973f
C513 B.n473 VSUBS 0.009973f
C514 B.n474 VSUBS 0.009973f
C515 B.n475 VSUBS 0.009973f
C516 B.n476 VSUBS 0.009973f
C517 B.n477 VSUBS 0.009973f
C518 B.n478 VSUBS 0.009973f
C519 B.n479 VSUBS 0.009973f
C520 B.n480 VSUBS 0.009973f
C521 B.n481 VSUBS 0.009973f
C522 B.n482 VSUBS 0.009973f
C523 B.n483 VSUBS 0.009973f
C524 B.n484 VSUBS 0.009973f
C525 B.n485 VSUBS 0.009973f
C526 B.n486 VSUBS 0.009973f
C527 B.n487 VSUBS 0.009973f
C528 B.n488 VSUBS 0.009973f
C529 B.n489 VSUBS 0.009973f
C530 B.n490 VSUBS 0.009973f
C531 B.n491 VSUBS 0.009973f
C532 B.n492 VSUBS 0.009973f
C533 B.n493 VSUBS 0.009973f
C534 B.n494 VSUBS 0.009973f
C535 B.n495 VSUBS 0.009973f
C536 B.n496 VSUBS 0.009973f
C537 B.n497 VSUBS 0.009973f
C538 B.n498 VSUBS 0.009973f
C539 B.n499 VSUBS 0.009973f
C540 B.n500 VSUBS 0.009973f
C541 B.n501 VSUBS 0.009973f
C542 B.n502 VSUBS 0.009973f
C543 B.n503 VSUBS 0.009973f
C544 B.n504 VSUBS 0.009973f
C545 B.n505 VSUBS 0.009973f
C546 B.n506 VSUBS 0.009973f
C547 B.n507 VSUBS 0.009973f
C548 B.n508 VSUBS 0.009973f
C549 B.n509 VSUBS 0.009973f
C550 B.n510 VSUBS 0.009973f
C551 B.n511 VSUBS 0.009973f
C552 B.n512 VSUBS 0.009973f
C553 B.n513 VSUBS 0.009973f
C554 B.n514 VSUBS 0.009973f
C555 B.n515 VSUBS 0.009973f
C556 B.n516 VSUBS 0.009973f
C557 B.n517 VSUBS 0.009973f
C558 B.n518 VSUBS 0.009973f
C559 B.n519 VSUBS 0.009973f
C560 B.n520 VSUBS 0.009973f
C561 B.n521 VSUBS 0.009973f
C562 B.n522 VSUBS 0.009973f
C563 B.n523 VSUBS 0.009973f
C564 B.n524 VSUBS 0.009973f
C565 B.n525 VSUBS 0.009973f
C566 B.n526 VSUBS 0.009973f
C567 B.n527 VSUBS 0.009973f
C568 B.n528 VSUBS 0.009973f
C569 B.n529 VSUBS 0.009973f
C570 B.n530 VSUBS 0.009973f
C571 B.n531 VSUBS 0.009973f
C572 B.n532 VSUBS 0.009973f
C573 B.n533 VSUBS 0.009973f
C574 B.n534 VSUBS 0.009973f
C575 B.n535 VSUBS 0.009973f
C576 B.n536 VSUBS 0.009973f
C577 B.n537 VSUBS 0.009973f
C578 B.n538 VSUBS 0.009973f
C579 B.n539 VSUBS 0.009973f
C580 B.n540 VSUBS 0.009973f
C581 B.n541 VSUBS 0.009973f
C582 B.n542 VSUBS 0.009973f
C583 B.n543 VSUBS 0.009973f
C584 B.n544 VSUBS 0.009973f
C585 B.n545 VSUBS 0.009973f
C586 B.n546 VSUBS 0.009973f
C587 B.n547 VSUBS 0.009973f
C588 B.n548 VSUBS 0.009973f
C589 B.n549 VSUBS 0.009973f
C590 B.n550 VSUBS 0.009973f
C591 B.n551 VSUBS 0.009973f
C592 B.n552 VSUBS 0.009973f
C593 B.n553 VSUBS 0.009973f
C594 B.n554 VSUBS 0.009973f
C595 B.n555 VSUBS 0.009973f
C596 B.n556 VSUBS 0.009973f
C597 B.n557 VSUBS 0.009973f
C598 B.n558 VSUBS 0.009973f
C599 B.n559 VSUBS 0.009973f
C600 B.n560 VSUBS 0.009973f
C601 B.n561 VSUBS 0.009973f
C602 B.n562 VSUBS 0.009973f
C603 B.n563 VSUBS 0.009973f
C604 B.n564 VSUBS 0.009973f
C605 B.n565 VSUBS 0.009973f
C606 B.n566 VSUBS 0.009973f
C607 B.n567 VSUBS 0.009973f
C608 B.n568 VSUBS 0.009973f
C609 B.n569 VSUBS 0.009973f
C610 B.n570 VSUBS 0.009973f
C611 B.n571 VSUBS 0.009973f
C612 B.n572 VSUBS 0.009973f
C613 B.n573 VSUBS 0.009973f
C614 B.n574 VSUBS 0.009973f
C615 B.n575 VSUBS 0.009973f
C616 B.n576 VSUBS 0.009973f
C617 B.n577 VSUBS 0.009973f
C618 B.n578 VSUBS 0.009973f
C619 B.n579 VSUBS 0.009973f
C620 B.n580 VSUBS 0.009973f
C621 B.n581 VSUBS 0.009973f
C622 B.n582 VSUBS 0.009973f
C623 B.n583 VSUBS 0.009973f
C624 B.n584 VSUBS 0.009973f
C625 B.n585 VSUBS 0.009973f
C626 B.n586 VSUBS 0.009973f
C627 B.n587 VSUBS 0.009973f
C628 B.n588 VSUBS 0.009973f
C629 B.n589 VSUBS 0.009973f
C630 B.n590 VSUBS 0.009973f
C631 B.n591 VSUBS 0.009973f
C632 B.n592 VSUBS 0.009973f
C633 B.n593 VSUBS 0.009973f
C634 B.n594 VSUBS 0.009973f
C635 B.n595 VSUBS 0.009973f
C636 B.n596 VSUBS 0.009973f
C637 B.n597 VSUBS 0.009973f
C638 B.n598 VSUBS 0.009973f
C639 B.n599 VSUBS 0.009973f
C640 B.n600 VSUBS 0.009973f
C641 B.n601 VSUBS 0.009973f
C642 B.n602 VSUBS 0.009973f
C643 B.n603 VSUBS 0.009973f
C644 B.n604 VSUBS 0.009973f
C645 B.n605 VSUBS 0.009973f
C646 B.n606 VSUBS 0.009973f
C647 B.n607 VSUBS 0.009973f
C648 B.n608 VSUBS 0.009973f
C649 B.n609 VSUBS 0.009973f
C650 B.n610 VSUBS 0.025309f
C651 B.n611 VSUBS 0.023679f
C652 B.n612 VSUBS 0.024774f
C653 B.n613 VSUBS 0.009973f
C654 B.n614 VSUBS 0.009973f
C655 B.n615 VSUBS 0.009973f
C656 B.n616 VSUBS 0.009973f
C657 B.n617 VSUBS 0.009973f
C658 B.n618 VSUBS 0.009973f
C659 B.n619 VSUBS 0.009973f
C660 B.n620 VSUBS 0.009973f
C661 B.n621 VSUBS 0.009973f
C662 B.n622 VSUBS 0.009973f
C663 B.n623 VSUBS 0.009973f
C664 B.n624 VSUBS 0.009973f
C665 B.n625 VSUBS 0.009973f
C666 B.n626 VSUBS 0.009973f
C667 B.n627 VSUBS 0.009973f
C668 B.n628 VSUBS 0.009973f
C669 B.n629 VSUBS 0.009973f
C670 B.n630 VSUBS 0.009973f
C671 B.n631 VSUBS 0.009973f
C672 B.n632 VSUBS 0.009973f
C673 B.n633 VSUBS 0.009973f
C674 B.n634 VSUBS 0.009973f
C675 B.n635 VSUBS 0.009973f
C676 B.n636 VSUBS 0.009973f
C677 B.n637 VSUBS 0.009973f
C678 B.n638 VSUBS 0.009973f
C679 B.n639 VSUBS 0.009973f
C680 B.n640 VSUBS 0.009973f
C681 B.n641 VSUBS 0.009973f
C682 B.n642 VSUBS 0.009973f
C683 B.n643 VSUBS 0.009973f
C684 B.n644 VSUBS 0.009973f
C685 B.n645 VSUBS 0.009973f
C686 B.n646 VSUBS 0.009973f
C687 B.n647 VSUBS 0.009387f
C688 B.n648 VSUBS 0.009973f
C689 B.n649 VSUBS 0.009973f
C690 B.n650 VSUBS 0.005573f
C691 B.n651 VSUBS 0.009973f
C692 B.n652 VSUBS 0.009973f
C693 B.n653 VSUBS 0.009973f
C694 B.n654 VSUBS 0.009973f
C695 B.n655 VSUBS 0.009973f
C696 B.n656 VSUBS 0.009973f
C697 B.n657 VSUBS 0.009973f
C698 B.n658 VSUBS 0.009973f
C699 B.n659 VSUBS 0.009973f
C700 B.n660 VSUBS 0.009973f
C701 B.n661 VSUBS 0.009973f
C702 B.n662 VSUBS 0.009973f
C703 B.n663 VSUBS 0.005573f
C704 B.n664 VSUBS 0.023107f
C705 B.n665 VSUBS 0.009387f
C706 B.n666 VSUBS 0.009973f
C707 B.n667 VSUBS 0.009973f
C708 B.n668 VSUBS 0.009973f
C709 B.n669 VSUBS 0.009973f
C710 B.n670 VSUBS 0.009973f
C711 B.n671 VSUBS 0.009973f
C712 B.n672 VSUBS 0.009973f
C713 B.n673 VSUBS 0.009973f
C714 B.n674 VSUBS 0.009973f
C715 B.n675 VSUBS 0.009973f
C716 B.n676 VSUBS 0.009973f
C717 B.n677 VSUBS 0.009973f
C718 B.n678 VSUBS 0.009973f
C719 B.n679 VSUBS 0.009973f
C720 B.n680 VSUBS 0.009973f
C721 B.n681 VSUBS 0.009973f
C722 B.n682 VSUBS 0.009973f
C723 B.n683 VSUBS 0.009973f
C724 B.n684 VSUBS 0.009973f
C725 B.n685 VSUBS 0.009973f
C726 B.n686 VSUBS 0.009973f
C727 B.n687 VSUBS 0.009973f
C728 B.n688 VSUBS 0.009973f
C729 B.n689 VSUBS 0.009973f
C730 B.n690 VSUBS 0.009973f
C731 B.n691 VSUBS 0.009973f
C732 B.n692 VSUBS 0.009973f
C733 B.n693 VSUBS 0.009973f
C734 B.n694 VSUBS 0.009973f
C735 B.n695 VSUBS 0.009973f
C736 B.n696 VSUBS 0.009973f
C737 B.n697 VSUBS 0.009973f
C738 B.n698 VSUBS 0.009973f
C739 B.n699 VSUBS 0.009973f
C740 B.n700 VSUBS 0.009973f
C741 B.n701 VSUBS 0.024774f
C742 B.n702 VSUBS 0.024774f
C743 B.n703 VSUBS 0.024213f
C744 B.n704 VSUBS 0.009973f
C745 B.n705 VSUBS 0.009973f
C746 B.n706 VSUBS 0.009973f
C747 B.n707 VSUBS 0.009973f
C748 B.n708 VSUBS 0.009973f
C749 B.n709 VSUBS 0.009973f
C750 B.n710 VSUBS 0.009973f
C751 B.n711 VSUBS 0.009973f
C752 B.n712 VSUBS 0.009973f
C753 B.n713 VSUBS 0.009973f
C754 B.n714 VSUBS 0.009973f
C755 B.n715 VSUBS 0.009973f
C756 B.n716 VSUBS 0.009973f
C757 B.n717 VSUBS 0.009973f
C758 B.n718 VSUBS 0.009973f
C759 B.n719 VSUBS 0.009973f
C760 B.n720 VSUBS 0.009973f
C761 B.n721 VSUBS 0.009973f
C762 B.n722 VSUBS 0.009973f
C763 B.n723 VSUBS 0.009973f
C764 B.n724 VSUBS 0.009973f
C765 B.n725 VSUBS 0.009973f
C766 B.n726 VSUBS 0.009973f
C767 B.n727 VSUBS 0.009973f
C768 B.n728 VSUBS 0.009973f
C769 B.n729 VSUBS 0.009973f
C770 B.n730 VSUBS 0.009973f
C771 B.n731 VSUBS 0.009973f
C772 B.n732 VSUBS 0.009973f
C773 B.n733 VSUBS 0.009973f
C774 B.n734 VSUBS 0.009973f
C775 B.n735 VSUBS 0.009973f
C776 B.n736 VSUBS 0.009973f
C777 B.n737 VSUBS 0.009973f
C778 B.n738 VSUBS 0.009973f
C779 B.n739 VSUBS 0.009973f
C780 B.n740 VSUBS 0.009973f
C781 B.n741 VSUBS 0.009973f
C782 B.n742 VSUBS 0.009973f
C783 B.n743 VSUBS 0.009973f
C784 B.n744 VSUBS 0.009973f
C785 B.n745 VSUBS 0.009973f
C786 B.n746 VSUBS 0.009973f
C787 B.n747 VSUBS 0.009973f
C788 B.n748 VSUBS 0.009973f
C789 B.n749 VSUBS 0.009973f
C790 B.n750 VSUBS 0.009973f
C791 B.n751 VSUBS 0.009973f
C792 B.n752 VSUBS 0.009973f
C793 B.n753 VSUBS 0.009973f
C794 B.n754 VSUBS 0.009973f
C795 B.n755 VSUBS 0.009973f
C796 B.n756 VSUBS 0.009973f
C797 B.n757 VSUBS 0.009973f
C798 B.n758 VSUBS 0.009973f
C799 B.n759 VSUBS 0.009973f
C800 B.n760 VSUBS 0.009973f
C801 B.n761 VSUBS 0.009973f
C802 B.n762 VSUBS 0.009973f
C803 B.n763 VSUBS 0.009973f
C804 B.n764 VSUBS 0.009973f
C805 B.n765 VSUBS 0.009973f
C806 B.n766 VSUBS 0.009973f
C807 B.n767 VSUBS 0.009973f
C808 B.n768 VSUBS 0.009973f
C809 B.n769 VSUBS 0.009973f
C810 B.n770 VSUBS 0.009973f
C811 B.n771 VSUBS 0.009973f
C812 B.n772 VSUBS 0.009973f
C813 B.n773 VSUBS 0.009973f
C814 B.n774 VSUBS 0.009973f
C815 B.n775 VSUBS 0.009973f
C816 B.n776 VSUBS 0.009973f
C817 B.n777 VSUBS 0.009973f
C818 B.n778 VSUBS 0.009973f
C819 B.n779 VSUBS 0.009973f
C820 B.n780 VSUBS 0.009973f
C821 B.n781 VSUBS 0.009973f
C822 B.n782 VSUBS 0.009973f
C823 B.n783 VSUBS 0.009973f
C824 B.n784 VSUBS 0.009973f
C825 B.n785 VSUBS 0.009973f
C826 B.n786 VSUBS 0.009973f
C827 B.n787 VSUBS 0.009973f
C828 B.n788 VSUBS 0.009973f
C829 B.n789 VSUBS 0.009973f
C830 B.n790 VSUBS 0.009973f
C831 B.n791 VSUBS 0.009973f
C832 B.n792 VSUBS 0.009973f
C833 B.n793 VSUBS 0.009973f
C834 B.n794 VSUBS 0.009973f
C835 B.n795 VSUBS 0.009973f
C836 B.n796 VSUBS 0.009973f
C837 B.n797 VSUBS 0.009973f
C838 B.n798 VSUBS 0.009973f
C839 B.n799 VSUBS 0.009973f
C840 B.n800 VSUBS 0.009973f
C841 B.n801 VSUBS 0.009973f
C842 B.n802 VSUBS 0.009973f
C843 B.n803 VSUBS 0.009973f
C844 B.n804 VSUBS 0.009973f
C845 B.n805 VSUBS 0.009973f
C846 B.n806 VSUBS 0.009973f
C847 B.n807 VSUBS 0.022583f
C848 VDD1.t5 VSUBS 0.172182f
C849 VDD1.t3 VSUBS 0.172182f
C850 VDD1.n0 VSUBS 1.21245f
C851 VDD1.t4 VSUBS 0.172182f
C852 VDD1.t7 VSUBS 0.172182f
C853 VDD1.n1 VSUBS 1.21086f
C854 VDD1.t1 VSUBS 0.172182f
C855 VDD1.t2 VSUBS 0.172182f
C856 VDD1.n2 VSUBS 1.21086f
C857 VDD1.n3 VSUBS 5.45469f
C858 VDD1.t0 VSUBS 0.172182f
C859 VDD1.t6 VSUBS 0.172182f
C860 VDD1.n4 VSUBS 1.18994f
C861 VDD1.n5 VSUBS 4.25067f
C862 VP.n0 VSUBS 0.064059f
C863 VP.t5 VSUBS 2.24601f
C864 VP.n1 VSUBS 0.06785f
C865 VP.n2 VSUBS 0.034056f
C866 VP.n3 VSUBS 0.063472f
C867 VP.n4 VSUBS 0.034056f
C868 VP.t6 VSUBS 2.24601f
C869 VP.n5 VSUBS 0.063472f
C870 VP.n6 VSUBS 0.034056f
C871 VP.n7 VSUBS 0.063472f
C872 VP.n8 VSUBS 0.034056f
C873 VP.t0 VSUBS 2.24601f
C874 VP.n9 VSUBS 0.063472f
C875 VP.n10 VSUBS 0.034056f
C876 VP.n11 VSUBS 0.063472f
C877 VP.n12 VSUBS 0.064059f
C878 VP.t1 VSUBS 2.24601f
C879 VP.n13 VSUBS 0.06785f
C880 VP.n14 VSUBS 0.034056f
C881 VP.n15 VSUBS 0.063472f
C882 VP.n16 VSUBS 0.034056f
C883 VP.t7 VSUBS 2.24601f
C884 VP.n17 VSUBS 0.063472f
C885 VP.n18 VSUBS 0.034056f
C886 VP.n19 VSUBS 0.063472f
C887 VP.t2 VSUBS 2.72321f
C888 VP.n20 VSUBS 0.917526f
C889 VP.t4 VSUBS 2.24601f
C890 VP.n21 VSUBS 0.947261f
C891 VP.n22 VSUBS 0.052191f
C892 VP.n23 VSUBS 0.443564f
C893 VP.n24 VSUBS 0.034056f
C894 VP.n25 VSUBS 0.034056f
C895 VP.n26 VSUBS 0.063472f
C896 VP.n27 VSUBS 0.049716f
C897 VP.n28 VSUBS 0.049716f
C898 VP.n29 VSUBS 0.034056f
C899 VP.n30 VSUBS 0.034056f
C900 VP.n31 VSUBS 0.034056f
C901 VP.n32 VSUBS 0.063472f
C902 VP.n33 VSUBS 0.052191f
C903 VP.n34 VSUBS 0.82041f
C904 VP.n35 VSUBS 0.043416f
C905 VP.n36 VSUBS 0.034056f
C906 VP.n37 VSUBS 0.034056f
C907 VP.n38 VSUBS 0.034056f
C908 VP.n39 VSUBS 0.063472f
C909 VP.n40 VSUBS 0.061833f
C910 VP.n41 VSUBS 0.033219f
C911 VP.n42 VSUBS 0.034056f
C912 VP.n43 VSUBS 0.034056f
C913 VP.n44 VSUBS 0.034056f
C914 VP.n45 VSUBS 0.063472f
C915 VP.n46 VSUBS 0.060965f
C916 VP.n47 VSUBS 0.970581f
C917 VP.n48 VSUBS 2.12154f
C918 VP.n49 VSUBS 2.1448f
C919 VP.t3 VSUBS 2.24601f
C920 VP.n50 VSUBS 0.970581f
C921 VP.n51 VSUBS 0.060965f
C922 VP.n52 VSUBS 0.064059f
C923 VP.n53 VSUBS 0.034056f
C924 VP.n54 VSUBS 0.034056f
C925 VP.n55 VSUBS 0.06785f
C926 VP.n56 VSUBS 0.033219f
C927 VP.n57 VSUBS 0.061833f
C928 VP.n58 VSUBS 0.034056f
C929 VP.n59 VSUBS 0.034056f
C930 VP.n60 VSUBS 0.034056f
C931 VP.n61 VSUBS 0.063472f
C932 VP.n62 VSUBS 0.043416f
C933 VP.n63 VSUBS 0.82041f
C934 VP.n64 VSUBS 0.052191f
C935 VP.n65 VSUBS 0.034056f
C936 VP.n66 VSUBS 0.034056f
C937 VP.n67 VSUBS 0.034056f
C938 VP.n68 VSUBS 0.063472f
C939 VP.n69 VSUBS 0.049716f
C940 VP.n70 VSUBS 0.049716f
C941 VP.n71 VSUBS 0.034056f
C942 VP.n72 VSUBS 0.034056f
C943 VP.n73 VSUBS 0.034056f
C944 VP.n74 VSUBS 0.063472f
C945 VP.n75 VSUBS 0.052191f
C946 VP.n76 VSUBS 0.82041f
C947 VP.n77 VSUBS 0.043416f
C948 VP.n78 VSUBS 0.034056f
C949 VP.n79 VSUBS 0.034056f
C950 VP.n80 VSUBS 0.034056f
C951 VP.n81 VSUBS 0.063472f
C952 VP.n82 VSUBS 0.061833f
C953 VP.n83 VSUBS 0.033219f
C954 VP.n84 VSUBS 0.034056f
C955 VP.n85 VSUBS 0.034056f
C956 VP.n86 VSUBS 0.034056f
C957 VP.n87 VSUBS 0.063472f
C958 VP.n88 VSUBS 0.060965f
C959 VP.n89 VSUBS 0.970581f
C960 VP.n90 VSUBS 0.101754f
C961 VTAIL.t9 VSUBS 0.156945f
C962 VTAIL.t14 VSUBS 0.156945f
C963 VTAIL.n0 VSUBS 0.976461f
C964 VTAIL.n1 VSUBS 0.909619f
C965 VTAIL.n2 VSUBS 0.017166f
C966 VTAIL.n3 VSUBS 0.038749f
C967 VTAIL.n4 VSUBS 0.017358f
C968 VTAIL.n5 VSUBS 0.030508f
C969 VTAIL.n6 VSUBS 0.016394f
C970 VTAIL.n7 VSUBS 0.038749f
C971 VTAIL.n8 VSUBS 0.017358f
C972 VTAIL.n9 VSUBS 0.030508f
C973 VTAIL.n10 VSUBS 0.016394f
C974 VTAIL.n11 VSUBS 0.029062f
C975 VTAIL.n12 VSUBS 0.029145f
C976 VTAIL.t10 VSUBS 0.083291f
C977 VTAIL.n13 VSUBS 0.164826f
C978 VTAIL.n14 VSUBS 0.764436f
C979 VTAIL.n15 VSUBS 0.016394f
C980 VTAIL.n16 VSUBS 0.017358f
C981 VTAIL.n17 VSUBS 0.038749f
C982 VTAIL.n18 VSUBS 0.038749f
C983 VTAIL.n19 VSUBS 0.017358f
C984 VTAIL.n20 VSUBS 0.016394f
C985 VTAIL.n21 VSUBS 0.030508f
C986 VTAIL.n22 VSUBS 0.030508f
C987 VTAIL.n23 VSUBS 0.016394f
C988 VTAIL.n24 VSUBS 0.017358f
C989 VTAIL.n25 VSUBS 0.038749f
C990 VTAIL.n26 VSUBS 0.038749f
C991 VTAIL.n27 VSUBS 0.017358f
C992 VTAIL.n28 VSUBS 0.016394f
C993 VTAIL.n29 VSUBS 0.030508f
C994 VTAIL.n30 VSUBS 0.076769f
C995 VTAIL.n31 VSUBS 0.016394f
C996 VTAIL.n32 VSUBS 0.017358f
C997 VTAIL.n33 VSUBS 0.085883f
C998 VTAIL.n34 VSUBS 0.056561f
C999 VTAIL.n35 VSUBS 0.426147f
C1000 VTAIL.n36 VSUBS 0.017166f
C1001 VTAIL.n37 VSUBS 0.038749f
C1002 VTAIL.n38 VSUBS 0.017358f
C1003 VTAIL.n39 VSUBS 0.030508f
C1004 VTAIL.n40 VSUBS 0.016394f
C1005 VTAIL.n41 VSUBS 0.038749f
C1006 VTAIL.n42 VSUBS 0.017358f
C1007 VTAIL.n43 VSUBS 0.030508f
C1008 VTAIL.n44 VSUBS 0.016394f
C1009 VTAIL.n45 VSUBS 0.029062f
C1010 VTAIL.n46 VSUBS 0.029145f
C1011 VTAIL.t7 VSUBS 0.083291f
C1012 VTAIL.n47 VSUBS 0.164826f
C1013 VTAIL.n48 VSUBS 0.764436f
C1014 VTAIL.n49 VSUBS 0.016394f
C1015 VTAIL.n50 VSUBS 0.017358f
C1016 VTAIL.n51 VSUBS 0.038749f
C1017 VTAIL.n52 VSUBS 0.038749f
C1018 VTAIL.n53 VSUBS 0.017358f
C1019 VTAIL.n54 VSUBS 0.016394f
C1020 VTAIL.n55 VSUBS 0.030508f
C1021 VTAIL.n56 VSUBS 0.030508f
C1022 VTAIL.n57 VSUBS 0.016394f
C1023 VTAIL.n58 VSUBS 0.017358f
C1024 VTAIL.n59 VSUBS 0.038749f
C1025 VTAIL.n60 VSUBS 0.038749f
C1026 VTAIL.n61 VSUBS 0.017358f
C1027 VTAIL.n62 VSUBS 0.016394f
C1028 VTAIL.n63 VSUBS 0.030508f
C1029 VTAIL.n64 VSUBS 0.076769f
C1030 VTAIL.n65 VSUBS 0.016394f
C1031 VTAIL.n66 VSUBS 0.017358f
C1032 VTAIL.n67 VSUBS 0.085883f
C1033 VTAIL.n68 VSUBS 0.056561f
C1034 VTAIL.n69 VSUBS 0.426147f
C1035 VTAIL.t3 VSUBS 0.156945f
C1036 VTAIL.t6 VSUBS 0.156945f
C1037 VTAIL.n70 VSUBS 0.976461f
C1038 VTAIL.n71 VSUBS 1.25474f
C1039 VTAIL.n72 VSUBS 0.017166f
C1040 VTAIL.n73 VSUBS 0.038749f
C1041 VTAIL.n74 VSUBS 0.017358f
C1042 VTAIL.n75 VSUBS 0.030508f
C1043 VTAIL.n76 VSUBS 0.016394f
C1044 VTAIL.n77 VSUBS 0.038749f
C1045 VTAIL.n78 VSUBS 0.017358f
C1046 VTAIL.n79 VSUBS 0.030508f
C1047 VTAIL.n80 VSUBS 0.016394f
C1048 VTAIL.n81 VSUBS 0.029062f
C1049 VTAIL.n82 VSUBS 0.029145f
C1050 VTAIL.t2 VSUBS 0.083291f
C1051 VTAIL.n83 VSUBS 0.164826f
C1052 VTAIL.n84 VSUBS 0.764436f
C1053 VTAIL.n85 VSUBS 0.016394f
C1054 VTAIL.n86 VSUBS 0.017358f
C1055 VTAIL.n87 VSUBS 0.038749f
C1056 VTAIL.n88 VSUBS 0.038749f
C1057 VTAIL.n89 VSUBS 0.017358f
C1058 VTAIL.n90 VSUBS 0.016394f
C1059 VTAIL.n91 VSUBS 0.030508f
C1060 VTAIL.n92 VSUBS 0.030508f
C1061 VTAIL.n93 VSUBS 0.016394f
C1062 VTAIL.n94 VSUBS 0.017358f
C1063 VTAIL.n95 VSUBS 0.038749f
C1064 VTAIL.n96 VSUBS 0.038749f
C1065 VTAIL.n97 VSUBS 0.017358f
C1066 VTAIL.n98 VSUBS 0.016394f
C1067 VTAIL.n99 VSUBS 0.030508f
C1068 VTAIL.n100 VSUBS 0.076769f
C1069 VTAIL.n101 VSUBS 0.016394f
C1070 VTAIL.n102 VSUBS 0.017358f
C1071 VTAIL.n103 VSUBS 0.085883f
C1072 VTAIL.n104 VSUBS 0.056561f
C1073 VTAIL.n105 VSUBS 1.6969f
C1074 VTAIL.n106 VSUBS 0.017166f
C1075 VTAIL.n107 VSUBS 0.038749f
C1076 VTAIL.n108 VSUBS 0.017358f
C1077 VTAIL.n109 VSUBS 0.030508f
C1078 VTAIL.n110 VSUBS 0.016394f
C1079 VTAIL.n111 VSUBS 0.038749f
C1080 VTAIL.n112 VSUBS 0.017358f
C1081 VTAIL.n113 VSUBS 0.030508f
C1082 VTAIL.n114 VSUBS 0.016394f
C1083 VTAIL.n115 VSUBS 0.029062f
C1084 VTAIL.n116 VSUBS 0.029145f
C1085 VTAIL.t15 VSUBS 0.083291f
C1086 VTAIL.n117 VSUBS 0.164826f
C1087 VTAIL.n118 VSUBS 0.764436f
C1088 VTAIL.n119 VSUBS 0.016394f
C1089 VTAIL.n120 VSUBS 0.017358f
C1090 VTAIL.n121 VSUBS 0.038749f
C1091 VTAIL.n122 VSUBS 0.038749f
C1092 VTAIL.n123 VSUBS 0.017358f
C1093 VTAIL.n124 VSUBS 0.016394f
C1094 VTAIL.n125 VSUBS 0.030508f
C1095 VTAIL.n126 VSUBS 0.030508f
C1096 VTAIL.n127 VSUBS 0.016394f
C1097 VTAIL.n128 VSUBS 0.017358f
C1098 VTAIL.n129 VSUBS 0.038749f
C1099 VTAIL.n130 VSUBS 0.038749f
C1100 VTAIL.n131 VSUBS 0.017358f
C1101 VTAIL.n132 VSUBS 0.016394f
C1102 VTAIL.n133 VSUBS 0.030508f
C1103 VTAIL.n134 VSUBS 0.076769f
C1104 VTAIL.n135 VSUBS 0.016394f
C1105 VTAIL.n136 VSUBS 0.017358f
C1106 VTAIL.n137 VSUBS 0.085883f
C1107 VTAIL.n138 VSUBS 0.056561f
C1108 VTAIL.n139 VSUBS 1.6969f
C1109 VTAIL.t11 VSUBS 0.156945f
C1110 VTAIL.t8 VSUBS 0.156945f
C1111 VTAIL.n140 VSUBS 0.976465f
C1112 VTAIL.n141 VSUBS 1.25474f
C1113 VTAIL.n142 VSUBS 0.017166f
C1114 VTAIL.n143 VSUBS 0.038749f
C1115 VTAIL.n144 VSUBS 0.017358f
C1116 VTAIL.n145 VSUBS 0.030508f
C1117 VTAIL.n146 VSUBS 0.016394f
C1118 VTAIL.n147 VSUBS 0.038749f
C1119 VTAIL.n148 VSUBS 0.017358f
C1120 VTAIL.n149 VSUBS 0.030508f
C1121 VTAIL.n150 VSUBS 0.016394f
C1122 VTAIL.n151 VSUBS 0.029062f
C1123 VTAIL.n152 VSUBS 0.029145f
C1124 VTAIL.t12 VSUBS 0.083291f
C1125 VTAIL.n153 VSUBS 0.164826f
C1126 VTAIL.n154 VSUBS 0.764436f
C1127 VTAIL.n155 VSUBS 0.016394f
C1128 VTAIL.n156 VSUBS 0.017358f
C1129 VTAIL.n157 VSUBS 0.038749f
C1130 VTAIL.n158 VSUBS 0.038749f
C1131 VTAIL.n159 VSUBS 0.017358f
C1132 VTAIL.n160 VSUBS 0.016394f
C1133 VTAIL.n161 VSUBS 0.030508f
C1134 VTAIL.n162 VSUBS 0.030508f
C1135 VTAIL.n163 VSUBS 0.016394f
C1136 VTAIL.n164 VSUBS 0.017358f
C1137 VTAIL.n165 VSUBS 0.038749f
C1138 VTAIL.n166 VSUBS 0.038749f
C1139 VTAIL.n167 VSUBS 0.017358f
C1140 VTAIL.n168 VSUBS 0.016394f
C1141 VTAIL.n169 VSUBS 0.030508f
C1142 VTAIL.n170 VSUBS 0.076769f
C1143 VTAIL.n171 VSUBS 0.016394f
C1144 VTAIL.n172 VSUBS 0.017358f
C1145 VTAIL.n173 VSUBS 0.085883f
C1146 VTAIL.n174 VSUBS 0.056561f
C1147 VTAIL.n175 VSUBS 0.426147f
C1148 VTAIL.n176 VSUBS 0.017166f
C1149 VTAIL.n177 VSUBS 0.038749f
C1150 VTAIL.n178 VSUBS 0.017358f
C1151 VTAIL.n179 VSUBS 0.030508f
C1152 VTAIL.n180 VSUBS 0.016394f
C1153 VTAIL.n181 VSUBS 0.038749f
C1154 VTAIL.n182 VSUBS 0.017358f
C1155 VTAIL.n183 VSUBS 0.030508f
C1156 VTAIL.n184 VSUBS 0.016394f
C1157 VTAIL.n185 VSUBS 0.029062f
C1158 VTAIL.n186 VSUBS 0.029145f
C1159 VTAIL.t1 VSUBS 0.083291f
C1160 VTAIL.n187 VSUBS 0.164826f
C1161 VTAIL.n188 VSUBS 0.764436f
C1162 VTAIL.n189 VSUBS 0.016394f
C1163 VTAIL.n190 VSUBS 0.017358f
C1164 VTAIL.n191 VSUBS 0.038749f
C1165 VTAIL.n192 VSUBS 0.038749f
C1166 VTAIL.n193 VSUBS 0.017358f
C1167 VTAIL.n194 VSUBS 0.016394f
C1168 VTAIL.n195 VSUBS 0.030508f
C1169 VTAIL.n196 VSUBS 0.030508f
C1170 VTAIL.n197 VSUBS 0.016394f
C1171 VTAIL.n198 VSUBS 0.017358f
C1172 VTAIL.n199 VSUBS 0.038749f
C1173 VTAIL.n200 VSUBS 0.038749f
C1174 VTAIL.n201 VSUBS 0.017358f
C1175 VTAIL.n202 VSUBS 0.016394f
C1176 VTAIL.n203 VSUBS 0.030508f
C1177 VTAIL.n204 VSUBS 0.076769f
C1178 VTAIL.n205 VSUBS 0.016394f
C1179 VTAIL.n206 VSUBS 0.017358f
C1180 VTAIL.n207 VSUBS 0.085883f
C1181 VTAIL.n208 VSUBS 0.056561f
C1182 VTAIL.n209 VSUBS 0.426147f
C1183 VTAIL.t0 VSUBS 0.156945f
C1184 VTAIL.t4 VSUBS 0.156945f
C1185 VTAIL.n210 VSUBS 0.976465f
C1186 VTAIL.n211 VSUBS 1.25474f
C1187 VTAIL.n212 VSUBS 0.017166f
C1188 VTAIL.n213 VSUBS 0.038749f
C1189 VTAIL.n214 VSUBS 0.017358f
C1190 VTAIL.n215 VSUBS 0.030508f
C1191 VTAIL.n216 VSUBS 0.016394f
C1192 VTAIL.n217 VSUBS 0.038749f
C1193 VTAIL.n218 VSUBS 0.017358f
C1194 VTAIL.n219 VSUBS 0.030508f
C1195 VTAIL.n220 VSUBS 0.016394f
C1196 VTAIL.n221 VSUBS 0.029062f
C1197 VTAIL.n222 VSUBS 0.029145f
C1198 VTAIL.t5 VSUBS 0.083291f
C1199 VTAIL.n223 VSUBS 0.164826f
C1200 VTAIL.n224 VSUBS 0.764436f
C1201 VTAIL.n225 VSUBS 0.016394f
C1202 VTAIL.n226 VSUBS 0.017358f
C1203 VTAIL.n227 VSUBS 0.038749f
C1204 VTAIL.n228 VSUBS 0.038749f
C1205 VTAIL.n229 VSUBS 0.017358f
C1206 VTAIL.n230 VSUBS 0.016394f
C1207 VTAIL.n231 VSUBS 0.030508f
C1208 VTAIL.n232 VSUBS 0.030508f
C1209 VTAIL.n233 VSUBS 0.016394f
C1210 VTAIL.n234 VSUBS 0.017358f
C1211 VTAIL.n235 VSUBS 0.038749f
C1212 VTAIL.n236 VSUBS 0.038749f
C1213 VTAIL.n237 VSUBS 0.017358f
C1214 VTAIL.n238 VSUBS 0.016394f
C1215 VTAIL.n239 VSUBS 0.030508f
C1216 VTAIL.n240 VSUBS 0.076769f
C1217 VTAIL.n241 VSUBS 0.016394f
C1218 VTAIL.n242 VSUBS 0.017358f
C1219 VTAIL.n243 VSUBS 0.085883f
C1220 VTAIL.n244 VSUBS 0.056561f
C1221 VTAIL.n245 VSUBS 1.6969f
C1222 VTAIL.n246 VSUBS 0.017166f
C1223 VTAIL.n247 VSUBS 0.038749f
C1224 VTAIL.n248 VSUBS 0.017358f
C1225 VTAIL.n249 VSUBS 0.030508f
C1226 VTAIL.n250 VSUBS 0.016394f
C1227 VTAIL.n251 VSUBS 0.038749f
C1228 VTAIL.n252 VSUBS 0.017358f
C1229 VTAIL.n253 VSUBS 0.030508f
C1230 VTAIL.n254 VSUBS 0.016394f
C1231 VTAIL.n255 VSUBS 0.029062f
C1232 VTAIL.n256 VSUBS 0.029145f
C1233 VTAIL.t13 VSUBS 0.083291f
C1234 VTAIL.n257 VSUBS 0.164826f
C1235 VTAIL.n258 VSUBS 0.764436f
C1236 VTAIL.n259 VSUBS 0.016394f
C1237 VTAIL.n260 VSUBS 0.017358f
C1238 VTAIL.n261 VSUBS 0.038749f
C1239 VTAIL.n262 VSUBS 0.038749f
C1240 VTAIL.n263 VSUBS 0.017358f
C1241 VTAIL.n264 VSUBS 0.016394f
C1242 VTAIL.n265 VSUBS 0.030508f
C1243 VTAIL.n266 VSUBS 0.030508f
C1244 VTAIL.n267 VSUBS 0.016394f
C1245 VTAIL.n268 VSUBS 0.017358f
C1246 VTAIL.n269 VSUBS 0.038749f
C1247 VTAIL.n270 VSUBS 0.038749f
C1248 VTAIL.n271 VSUBS 0.017358f
C1249 VTAIL.n272 VSUBS 0.016394f
C1250 VTAIL.n273 VSUBS 0.030508f
C1251 VTAIL.n274 VSUBS 0.076769f
C1252 VTAIL.n275 VSUBS 0.016394f
C1253 VTAIL.n276 VSUBS 0.017358f
C1254 VTAIL.n277 VSUBS 0.085883f
C1255 VTAIL.n278 VSUBS 0.056561f
C1256 VTAIL.n279 VSUBS 1.69118f
C1257 VDD2.t5 VSUBS 0.191353f
C1258 VDD2.t4 VSUBS 0.191353f
C1259 VDD2.n0 VSUBS 1.34568f
C1260 VDD2.t3 VSUBS 0.191353f
C1261 VDD2.t2 VSUBS 0.191353f
C1262 VDD2.n1 VSUBS 1.34568f
C1263 VDD2.n2 VSUBS 5.98527f
C1264 VDD2.t0 VSUBS 0.191353f
C1265 VDD2.t6 VSUBS 0.191353f
C1266 VDD2.n3 VSUBS 1.32244f
C1267 VDD2.n4 VSUBS 4.67728f
C1268 VDD2.t7 VSUBS 0.191353f
C1269 VDD2.t1 VSUBS 0.191353f
C1270 VDD2.n5 VSUBS 1.34563f
C1271 VN.n0 VSUBS 0.056696f
C1272 VN.t2 VSUBS 1.98786f
C1273 VN.n1 VSUBS 0.060051f
C1274 VN.n2 VSUBS 0.030142f
C1275 VN.n3 VSUBS 0.056176f
C1276 VN.n4 VSUBS 0.030142f
C1277 VN.t1 VSUBS 1.98786f
C1278 VN.n5 VSUBS 0.056176f
C1279 VN.n6 VSUBS 0.030142f
C1280 VN.n7 VSUBS 0.056176f
C1281 VN.t5 VSUBS 2.41021f
C1282 VN.n8 VSUBS 0.812065f
C1283 VN.t6 VSUBS 1.98786f
C1284 VN.n9 VSUBS 0.838385f
C1285 VN.n10 VSUBS 0.046192f
C1286 VN.n11 VSUBS 0.39258f
C1287 VN.n12 VSUBS 0.030142f
C1288 VN.n13 VSUBS 0.030142f
C1289 VN.n14 VSUBS 0.056176f
C1290 VN.n15 VSUBS 0.044001f
C1291 VN.n16 VSUBS 0.044001f
C1292 VN.n17 VSUBS 0.030142f
C1293 VN.n18 VSUBS 0.030142f
C1294 VN.n19 VSUBS 0.030142f
C1295 VN.n20 VSUBS 0.056176f
C1296 VN.n21 VSUBS 0.046192f
C1297 VN.n22 VSUBS 0.726114f
C1298 VN.n23 VSUBS 0.038426f
C1299 VN.n24 VSUBS 0.030142f
C1300 VN.n25 VSUBS 0.030142f
C1301 VN.n26 VSUBS 0.030142f
C1302 VN.n27 VSUBS 0.056176f
C1303 VN.n28 VSUBS 0.054726f
C1304 VN.n29 VSUBS 0.029401f
C1305 VN.n30 VSUBS 0.030142f
C1306 VN.n31 VSUBS 0.030142f
C1307 VN.n32 VSUBS 0.030142f
C1308 VN.n33 VSUBS 0.056176f
C1309 VN.n34 VSUBS 0.053958f
C1310 VN.n35 VSUBS 0.859025f
C1311 VN.n36 VSUBS 0.090058f
C1312 VN.n37 VSUBS 0.056696f
C1313 VN.t0 VSUBS 1.98786f
C1314 VN.n38 VSUBS 0.060051f
C1315 VN.n39 VSUBS 0.030142f
C1316 VN.n40 VSUBS 0.056176f
C1317 VN.n41 VSUBS 0.030142f
C1318 VN.t4 VSUBS 1.98786f
C1319 VN.n42 VSUBS 0.056176f
C1320 VN.n43 VSUBS 0.030142f
C1321 VN.n44 VSUBS 0.056176f
C1322 VN.t3 VSUBS 2.41021f
C1323 VN.n45 VSUBS 0.812065f
C1324 VN.t7 VSUBS 1.98786f
C1325 VN.n46 VSUBS 0.838385f
C1326 VN.n47 VSUBS 0.046192f
C1327 VN.n48 VSUBS 0.39258f
C1328 VN.n49 VSUBS 0.030142f
C1329 VN.n50 VSUBS 0.030142f
C1330 VN.n51 VSUBS 0.056176f
C1331 VN.n52 VSUBS 0.044001f
C1332 VN.n53 VSUBS 0.044001f
C1333 VN.n54 VSUBS 0.030142f
C1334 VN.n55 VSUBS 0.030142f
C1335 VN.n56 VSUBS 0.030142f
C1336 VN.n57 VSUBS 0.056176f
C1337 VN.n58 VSUBS 0.046192f
C1338 VN.n59 VSUBS 0.726114f
C1339 VN.n60 VSUBS 0.038426f
C1340 VN.n61 VSUBS 0.030142f
C1341 VN.n62 VSUBS 0.030142f
C1342 VN.n63 VSUBS 0.030142f
C1343 VN.n64 VSUBS 0.056176f
C1344 VN.n65 VSUBS 0.054726f
C1345 VN.n66 VSUBS 0.029401f
C1346 VN.n67 VSUBS 0.030142f
C1347 VN.n68 VSUBS 0.030142f
C1348 VN.n69 VSUBS 0.030142f
C1349 VN.n70 VSUBS 0.056176f
C1350 VN.n71 VSUBS 0.053958f
C1351 VN.n72 VSUBS 0.859025f
C1352 VN.n73 VSUBS 1.88529f
.ends

