* NGSPICE file created from diff_pair_sample_1389.ext - technology: sky130A

.subckt diff_pair_sample_1389 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=1.8447 ps=10.24 w=4.73 l=2.24
X1 B.t11 B.t9 B.t10 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=2.24
X2 B.t8 B.t6 B.t7 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=2.24
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=1.8447 ps=10.24 w=4.73 l=2.24
X4 VDD1.t0 VP.t1 VTAIL.t3 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=1.8447 ps=10.24 w=4.73 l=2.24
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=1.8447 ps=10.24 w=4.73 l=2.24
X6 B.t5 B.t3 B.t4 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=2.24
X7 B.t2 B.t0 B.t1 w_n1998_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=2.24
R0 VP.n0 VP.t1 138.255
R1 VP.n0 VP.t0 100.061
R2 VP VP.n0 0.336784
R3 VTAIL.n90 VTAIL.n72 756.745
R4 VTAIL.n18 VTAIL.n0 756.745
R5 VTAIL.n66 VTAIL.n48 756.745
R6 VTAIL.n42 VTAIL.n24 756.745
R7 VTAIL.n81 VTAIL.n80 585
R8 VTAIL.n83 VTAIL.n82 585
R9 VTAIL.n76 VTAIL.n75 585
R10 VTAIL.n89 VTAIL.n88 585
R11 VTAIL.n91 VTAIL.n90 585
R12 VTAIL.n9 VTAIL.n8 585
R13 VTAIL.n11 VTAIL.n10 585
R14 VTAIL.n4 VTAIL.n3 585
R15 VTAIL.n17 VTAIL.n16 585
R16 VTAIL.n19 VTAIL.n18 585
R17 VTAIL.n67 VTAIL.n66 585
R18 VTAIL.n65 VTAIL.n64 585
R19 VTAIL.n52 VTAIL.n51 585
R20 VTAIL.n59 VTAIL.n58 585
R21 VTAIL.n57 VTAIL.n56 585
R22 VTAIL.n43 VTAIL.n42 585
R23 VTAIL.n41 VTAIL.n40 585
R24 VTAIL.n28 VTAIL.n27 585
R25 VTAIL.n35 VTAIL.n34 585
R26 VTAIL.n33 VTAIL.n32 585
R27 VTAIL.n79 VTAIL.t1 328.587
R28 VTAIL.n7 VTAIL.t2 328.587
R29 VTAIL.n55 VTAIL.t3 328.587
R30 VTAIL.n31 VTAIL.t0 328.587
R31 VTAIL.n82 VTAIL.n81 171.744
R32 VTAIL.n82 VTAIL.n75 171.744
R33 VTAIL.n89 VTAIL.n75 171.744
R34 VTAIL.n90 VTAIL.n89 171.744
R35 VTAIL.n10 VTAIL.n9 171.744
R36 VTAIL.n10 VTAIL.n3 171.744
R37 VTAIL.n17 VTAIL.n3 171.744
R38 VTAIL.n18 VTAIL.n17 171.744
R39 VTAIL.n66 VTAIL.n65 171.744
R40 VTAIL.n65 VTAIL.n51 171.744
R41 VTAIL.n58 VTAIL.n51 171.744
R42 VTAIL.n58 VTAIL.n57 171.744
R43 VTAIL.n42 VTAIL.n41 171.744
R44 VTAIL.n41 VTAIL.n27 171.744
R45 VTAIL.n34 VTAIL.n27 171.744
R46 VTAIL.n34 VTAIL.n33 171.744
R47 VTAIL.n81 VTAIL.t1 85.8723
R48 VTAIL.n9 VTAIL.t2 85.8723
R49 VTAIL.n57 VTAIL.t3 85.8723
R50 VTAIL.n33 VTAIL.t0 85.8723
R51 VTAIL.n95 VTAIL.n94 35.4823
R52 VTAIL.n23 VTAIL.n22 35.4823
R53 VTAIL.n71 VTAIL.n70 35.4823
R54 VTAIL.n47 VTAIL.n46 35.4823
R55 VTAIL.n47 VTAIL.n23 20.8755
R56 VTAIL.n95 VTAIL.n71 18.66
R57 VTAIL.n80 VTAIL.n79 16.3651
R58 VTAIL.n8 VTAIL.n7 16.3651
R59 VTAIL.n56 VTAIL.n55 16.3651
R60 VTAIL.n32 VTAIL.n31 16.3651
R61 VTAIL.n83 VTAIL.n78 12.8005
R62 VTAIL.n11 VTAIL.n6 12.8005
R63 VTAIL.n59 VTAIL.n54 12.8005
R64 VTAIL.n35 VTAIL.n30 12.8005
R65 VTAIL.n84 VTAIL.n76 12.0247
R66 VTAIL.n12 VTAIL.n4 12.0247
R67 VTAIL.n60 VTAIL.n52 12.0247
R68 VTAIL.n36 VTAIL.n28 12.0247
R69 VTAIL.n88 VTAIL.n87 11.249
R70 VTAIL.n16 VTAIL.n15 11.249
R71 VTAIL.n64 VTAIL.n63 11.249
R72 VTAIL.n40 VTAIL.n39 11.249
R73 VTAIL.n91 VTAIL.n74 10.4732
R74 VTAIL.n19 VTAIL.n2 10.4732
R75 VTAIL.n67 VTAIL.n50 10.4732
R76 VTAIL.n43 VTAIL.n26 10.4732
R77 VTAIL.n92 VTAIL.n72 9.69747
R78 VTAIL.n20 VTAIL.n0 9.69747
R79 VTAIL.n68 VTAIL.n48 9.69747
R80 VTAIL.n44 VTAIL.n24 9.69747
R81 VTAIL.n94 VTAIL.n93 9.45567
R82 VTAIL.n22 VTAIL.n21 9.45567
R83 VTAIL.n70 VTAIL.n69 9.45567
R84 VTAIL.n46 VTAIL.n45 9.45567
R85 VTAIL.n93 VTAIL.n92 9.3005
R86 VTAIL.n74 VTAIL.n73 9.3005
R87 VTAIL.n87 VTAIL.n86 9.3005
R88 VTAIL.n85 VTAIL.n84 9.3005
R89 VTAIL.n78 VTAIL.n77 9.3005
R90 VTAIL.n21 VTAIL.n20 9.3005
R91 VTAIL.n2 VTAIL.n1 9.3005
R92 VTAIL.n15 VTAIL.n14 9.3005
R93 VTAIL.n13 VTAIL.n12 9.3005
R94 VTAIL.n6 VTAIL.n5 9.3005
R95 VTAIL.n69 VTAIL.n68 9.3005
R96 VTAIL.n50 VTAIL.n49 9.3005
R97 VTAIL.n63 VTAIL.n62 9.3005
R98 VTAIL.n61 VTAIL.n60 9.3005
R99 VTAIL.n54 VTAIL.n53 9.3005
R100 VTAIL.n45 VTAIL.n44 9.3005
R101 VTAIL.n26 VTAIL.n25 9.3005
R102 VTAIL.n39 VTAIL.n38 9.3005
R103 VTAIL.n37 VTAIL.n36 9.3005
R104 VTAIL.n30 VTAIL.n29 9.3005
R105 VTAIL.n94 VTAIL.n72 4.26717
R106 VTAIL.n22 VTAIL.n0 4.26717
R107 VTAIL.n70 VTAIL.n48 4.26717
R108 VTAIL.n46 VTAIL.n24 4.26717
R109 VTAIL.n79 VTAIL.n77 3.73474
R110 VTAIL.n7 VTAIL.n5 3.73474
R111 VTAIL.n55 VTAIL.n53 3.73474
R112 VTAIL.n31 VTAIL.n29 3.73474
R113 VTAIL.n92 VTAIL.n91 3.49141
R114 VTAIL.n20 VTAIL.n19 3.49141
R115 VTAIL.n68 VTAIL.n67 3.49141
R116 VTAIL.n44 VTAIL.n43 3.49141
R117 VTAIL.n88 VTAIL.n74 2.71565
R118 VTAIL.n16 VTAIL.n2 2.71565
R119 VTAIL.n64 VTAIL.n50 2.71565
R120 VTAIL.n40 VTAIL.n26 2.71565
R121 VTAIL.n87 VTAIL.n76 1.93989
R122 VTAIL.n15 VTAIL.n4 1.93989
R123 VTAIL.n63 VTAIL.n52 1.93989
R124 VTAIL.n39 VTAIL.n28 1.93989
R125 VTAIL.n71 VTAIL.n47 1.57809
R126 VTAIL.n84 VTAIL.n83 1.16414
R127 VTAIL.n12 VTAIL.n11 1.16414
R128 VTAIL.n60 VTAIL.n59 1.16414
R129 VTAIL.n36 VTAIL.n35 1.16414
R130 VTAIL VTAIL.n23 1.0824
R131 VTAIL VTAIL.n95 0.49619
R132 VTAIL.n80 VTAIL.n78 0.388379
R133 VTAIL.n8 VTAIL.n6 0.388379
R134 VTAIL.n56 VTAIL.n54 0.388379
R135 VTAIL.n32 VTAIL.n30 0.388379
R136 VTAIL.n85 VTAIL.n77 0.155672
R137 VTAIL.n86 VTAIL.n85 0.155672
R138 VTAIL.n86 VTAIL.n73 0.155672
R139 VTAIL.n93 VTAIL.n73 0.155672
R140 VTAIL.n13 VTAIL.n5 0.155672
R141 VTAIL.n14 VTAIL.n13 0.155672
R142 VTAIL.n14 VTAIL.n1 0.155672
R143 VTAIL.n21 VTAIL.n1 0.155672
R144 VTAIL.n69 VTAIL.n49 0.155672
R145 VTAIL.n62 VTAIL.n49 0.155672
R146 VTAIL.n62 VTAIL.n61 0.155672
R147 VTAIL.n61 VTAIL.n53 0.155672
R148 VTAIL.n45 VTAIL.n25 0.155672
R149 VTAIL.n38 VTAIL.n25 0.155672
R150 VTAIL.n38 VTAIL.n37 0.155672
R151 VTAIL.n37 VTAIL.n29 0.155672
R152 VDD1.n18 VDD1.n0 756.745
R153 VDD1.n41 VDD1.n23 756.745
R154 VDD1.n19 VDD1.n18 585
R155 VDD1.n17 VDD1.n16 585
R156 VDD1.n4 VDD1.n3 585
R157 VDD1.n11 VDD1.n10 585
R158 VDD1.n9 VDD1.n8 585
R159 VDD1.n32 VDD1.n31 585
R160 VDD1.n34 VDD1.n33 585
R161 VDD1.n27 VDD1.n26 585
R162 VDD1.n40 VDD1.n39 585
R163 VDD1.n42 VDD1.n41 585
R164 VDD1.n7 VDD1.t0 328.587
R165 VDD1.n30 VDD1.t1 328.587
R166 VDD1.n18 VDD1.n17 171.744
R167 VDD1.n17 VDD1.n3 171.744
R168 VDD1.n10 VDD1.n3 171.744
R169 VDD1.n10 VDD1.n9 171.744
R170 VDD1.n33 VDD1.n32 171.744
R171 VDD1.n33 VDD1.n26 171.744
R172 VDD1.n40 VDD1.n26 171.744
R173 VDD1.n41 VDD1.n40 171.744
R174 VDD1.n9 VDD1.t0 85.8723
R175 VDD1.n32 VDD1.t1 85.8723
R176 VDD1 VDD1.n45 85.4079
R177 VDD1 VDD1.n22 52.7732
R178 VDD1.n8 VDD1.n7 16.3651
R179 VDD1.n31 VDD1.n30 16.3651
R180 VDD1.n11 VDD1.n6 12.8005
R181 VDD1.n34 VDD1.n29 12.8005
R182 VDD1.n12 VDD1.n4 12.0247
R183 VDD1.n35 VDD1.n27 12.0247
R184 VDD1.n16 VDD1.n15 11.249
R185 VDD1.n39 VDD1.n38 11.249
R186 VDD1.n19 VDD1.n2 10.4732
R187 VDD1.n42 VDD1.n25 10.4732
R188 VDD1.n20 VDD1.n0 9.69747
R189 VDD1.n43 VDD1.n23 9.69747
R190 VDD1.n22 VDD1.n21 9.45567
R191 VDD1.n45 VDD1.n44 9.45567
R192 VDD1.n21 VDD1.n20 9.3005
R193 VDD1.n2 VDD1.n1 9.3005
R194 VDD1.n15 VDD1.n14 9.3005
R195 VDD1.n13 VDD1.n12 9.3005
R196 VDD1.n6 VDD1.n5 9.3005
R197 VDD1.n44 VDD1.n43 9.3005
R198 VDD1.n25 VDD1.n24 9.3005
R199 VDD1.n38 VDD1.n37 9.3005
R200 VDD1.n36 VDD1.n35 9.3005
R201 VDD1.n29 VDD1.n28 9.3005
R202 VDD1.n22 VDD1.n0 4.26717
R203 VDD1.n45 VDD1.n23 4.26717
R204 VDD1.n7 VDD1.n5 3.73474
R205 VDD1.n30 VDD1.n28 3.73474
R206 VDD1.n20 VDD1.n19 3.49141
R207 VDD1.n43 VDD1.n42 3.49141
R208 VDD1.n16 VDD1.n2 2.71565
R209 VDD1.n39 VDD1.n25 2.71565
R210 VDD1.n15 VDD1.n4 1.93989
R211 VDD1.n38 VDD1.n27 1.93989
R212 VDD1.n12 VDD1.n11 1.16414
R213 VDD1.n35 VDD1.n34 1.16414
R214 VDD1.n8 VDD1.n6 0.388379
R215 VDD1.n31 VDD1.n29 0.388379
R216 VDD1.n21 VDD1.n1 0.155672
R217 VDD1.n14 VDD1.n1 0.155672
R218 VDD1.n14 VDD1.n13 0.155672
R219 VDD1.n13 VDD1.n5 0.155672
R220 VDD1.n36 VDD1.n28 0.155672
R221 VDD1.n37 VDD1.n36 0.155672
R222 VDD1.n37 VDD1.n24 0.155672
R223 VDD1.n44 VDD1.n24 0.155672
R224 B.n288 B.n43 585
R225 B.n290 B.n289 585
R226 B.n291 B.n42 585
R227 B.n293 B.n292 585
R228 B.n294 B.n41 585
R229 B.n296 B.n295 585
R230 B.n297 B.n40 585
R231 B.n299 B.n298 585
R232 B.n300 B.n39 585
R233 B.n302 B.n301 585
R234 B.n303 B.n38 585
R235 B.n305 B.n304 585
R236 B.n306 B.n37 585
R237 B.n308 B.n307 585
R238 B.n309 B.n36 585
R239 B.n311 B.n310 585
R240 B.n312 B.n35 585
R241 B.n314 B.n313 585
R242 B.n315 B.n31 585
R243 B.n317 B.n316 585
R244 B.n318 B.n30 585
R245 B.n320 B.n319 585
R246 B.n321 B.n29 585
R247 B.n323 B.n322 585
R248 B.n324 B.n28 585
R249 B.n326 B.n325 585
R250 B.n327 B.n27 585
R251 B.n329 B.n328 585
R252 B.n330 B.n26 585
R253 B.n332 B.n331 585
R254 B.n334 B.n23 585
R255 B.n336 B.n335 585
R256 B.n337 B.n22 585
R257 B.n339 B.n338 585
R258 B.n340 B.n21 585
R259 B.n342 B.n341 585
R260 B.n343 B.n20 585
R261 B.n345 B.n344 585
R262 B.n346 B.n19 585
R263 B.n348 B.n347 585
R264 B.n349 B.n18 585
R265 B.n351 B.n350 585
R266 B.n352 B.n17 585
R267 B.n354 B.n353 585
R268 B.n355 B.n16 585
R269 B.n357 B.n356 585
R270 B.n358 B.n15 585
R271 B.n360 B.n359 585
R272 B.n361 B.n14 585
R273 B.n363 B.n362 585
R274 B.n287 B.n286 585
R275 B.n285 B.n44 585
R276 B.n284 B.n283 585
R277 B.n282 B.n45 585
R278 B.n281 B.n280 585
R279 B.n279 B.n46 585
R280 B.n278 B.n277 585
R281 B.n276 B.n47 585
R282 B.n275 B.n274 585
R283 B.n273 B.n48 585
R284 B.n272 B.n271 585
R285 B.n270 B.n49 585
R286 B.n269 B.n268 585
R287 B.n267 B.n50 585
R288 B.n266 B.n265 585
R289 B.n264 B.n51 585
R290 B.n263 B.n262 585
R291 B.n261 B.n52 585
R292 B.n260 B.n259 585
R293 B.n258 B.n53 585
R294 B.n257 B.n256 585
R295 B.n255 B.n54 585
R296 B.n254 B.n253 585
R297 B.n252 B.n55 585
R298 B.n251 B.n250 585
R299 B.n249 B.n56 585
R300 B.n248 B.n247 585
R301 B.n246 B.n57 585
R302 B.n245 B.n244 585
R303 B.n243 B.n58 585
R304 B.n242 B.n241 585
R305 B.n240 B.n59 585
R306 B.n239 B.n238 585
R307 B.n237 B.n60 585
R308 B.n236 B.n235 585
R309 B.n234 B.n61 585
R310 B.n233 B.n232 585
R311 B.n231 B.n62 585
R312 B.n230 B.n229 585
R313 B.n228 B.n63 585
R314 B.n227 B.n226 585
R315 B.n225 B.n64 585
R316 B.n224 B.n223 585
R317 B.n222 B.n65 585
R318 B.n221 B.n220 585
R319 B.n219 B.n66 585
R320 B.n218 B.n217 585
R321 B.n141 B.n96 585
R322 B.n143 B.n142 585
R323 B.n144 B.n95 585
R324 B.n146 B.n145 585
R325 B.n147 B.n94 585
R326 B.n149 B.n148 585
R327 B.n150 B.n93 585
R328 B.n152 B.n151 585
R329 B.n153 B.n92 585
R330 B.n155 B.n154 585
R331 B.n156 B.n91 585
R332 B.n158 B.n157 585
R333 B.n159 B.n90 585
R334 B.n161 B.n160 585
R335 B.n162 B.n89 585
R336 B.n164 B.n163 585
R337 B.n165 B.n88 585
R338 B.n167 B.n166 585
R339 B.n168 B.n87 585
R340 B.n170 B.n169 585
R341 B.n172 B.n84 585
R342 B.n174 B.n173 585
R343 B.n175 B.n83 585
R344 B.n177 B.n176 585
R345 B.n178 B.n82 585
R346 B.n180 B.n179 585
R347 B.n181 B.n81 585
R348 B.n183 B.n182 585
R349 B.n184 B.n80 585
R350 B.n186 B.n185 585
R351 B.n188 B.n187 585
R352 B.n189 B.n76 585
R353 B.n191 B.n190 585
R354 B.n192 B.n75 585
R355 B.n194 B.n193 585
R356 B.n195 B.n74 585
R357 B.n197 B.n196 585
R358 B.n198 B.n73 585
R359 B.n200 B.n199 585
R360 B.n201 B.n72 585
R361 B.n203 B.n202 585
R362 B.n204 B.n71 585
R363 B.n206 B.n205 585
R364 B.n207 B.n70 585
R365 B.n209 B.n208 585
R366 B.n210 B.n69 585
R367 B.n212 B.n211 585
R368 B.n213 B.n68 585
R369 B.n215 B.n214 585
R370 B.n216 B.n67 585
R371 B.n140 B.n139 585
R372 B.n138 B.n97 585
R373 B.n137 B.n136 585
R374 B.n135 B.n98 585
R375 B.n134 B.n133 585
R376 B.n132 B.n99 585
R377 B.n131 B.n130 585
R378 B.n129 B.n100 585
R379 B.n128 B.n127 585
R380 B.n126 B.n101 585
R381 B.n125 B.n124 585
R382 B.n123 B.n102 585
R383 B.n122 B.n121 585
R384 B.n120 B.n103 585
R385 B.n119 B.n118 585
R386 B.n117 B.n104 585
R387 B.n116 B.n115 585
R388 B.n114 B.n105 585
R389 B.n113 B.n112 585
R390 B.n111 B.n106 585
R391 B.n110 B.n109 585
R392 B.n108 B.n107 585
R393 B.n2 B.n0 585
R394 B.n397 B.n1 585
R395 B.n396 B.n395 585
R396 B.n394 B.n3 585
R397 B.n393 B.n392 585
R398 B.n391 B.n4 585
R399 B.n390 B.n389 585
R400 B.n388 B.n5 585
R401 B.n387 B.n386 585
R402 B.n385 B.n6 585
R403 B.n384 B.n383 585
R404 B.n382 B.n7 585
R405 B.n381 B.n380 585
R406 B.n379 B.n8 585
R407 B.n378 B.n377 585
R408 B.n376 B.n9 585
R409 B.n375 B.n374 585
R410 B.n373 B.n10 585
R411 B.n372 B.n371 585
R412 B.n370 B.n11 585
R413 B.n369 B.n368 585
R414 B.n367 B.n12 585
R415 B.n366 B.n365 585
R416 B.n364 B.n13 585
R417 B.n399 B.n398 585
R418 B.n139 B.n96 540.549
R419 B.n362 B.n13 540.549
R420 B.n217 B.n216 540.549
R421 B.n288 B.n287 540.549
R422 B.n77 B.t11 296.709
R423 B.n32 B.t4 296.709
R424 B.n85 B.t2 296.709
R425 B.n24 B.t7 296.709
R426 B.n77 B.t9 258.32
R427 B.n85 B.t0 258.32
R428 B.n24 B.t6 258.32
R429 B.n32 B.t3 258.32
R430 B.n78 B.t10 246.865
R431 B.n33 B.t5 246.865
R432 B.n86 B.t1 246.865
R433 B.n25 B.t8 246.865
R434 B.n139 B.n138 163.367
R435 B.n138 B.n137 163.367
R436 B.n137 B.n98 163.367
R437 B.n133 B.n98 163.367
R438 B.n133 B.n132 163.367
R439 B.n132 B.n131 163.367
R440 B.n131 B.n100 163.367
R441 B.n127 B.n100 163.367
R442 B.n127 B.n126 163.367
R443 B.n126 B.n125 163.367
R444 B.n125 B.n102 163.367
R445 B.n121 B.n102 163.367
R446 B.n121 B.n120 163.367
R447 B.n120 B.n119 163.367
R448 B.n119 B.n104 163.367
R449 B.n115 B.n104 163.367
R450 B.n115 B.n114 163.367
R451 B.n114 B.n113 163.367
R452 B.n113 B.n106 163.367
R453 B.n109 B.n106 163.367
R454 B.n109 B.n108 163.367
R455 B.n108 B.n2 163.367
R456 B.n398 B.n2 163.367
R457 B.n398 B.n397 163.367
R458 B.n397 B.n396 163.367
R459 B.n396 B.n3 163.367
R460 B.n392 B.n3 163.367
R461 B.n392 B.n391 163.367
R462 B.n391 B.n390 163.367
R463 B.n390 B.n5 163.367
R464 B.n386 B.n5 163.367
R465 B.n386 B.n385 163.367
R466 B.n385 B.n384 163.367
R467 B.n384 B.n7 163.367
R468 B.n380 B.n7 163.367
R469 B.n380 B.n379 163.367
R470 B.n379 B.n378 163.367
R471 B.n378 B.n9 163.367
R472 B.n374 B.n9 163.367
R473 B.n374 B.n373 163.367
R474 B.n373 B.n372 163.367
R475 B.n372 B.n11 163.367
R476 B.n368 B.n11 163.367
R477 B.n368 B.n367 163.367
R478 B.n367 B.n366 163.367
R479 B.n366 B.n13 163.367
R480 B.n143 B.n96 163.367
R481 B.n144 B.n143 163.367
R482 B.n145 B.n144 163.367
R483 B.n145 B.n94 163.367
R484 B.n149 B.n94 163.367
R485 B.n150 B.n149 163.367
R486 B.n151 B.n150 163.367
R487 B.n151 B.n92 163.367
R488 B.n155 B.n92 163.367
R489 B.n156 B.n155 163.367
R490 B.n157 B.n156 163.367
R491 B.n157 B.n90 163.367
R492 B.n161 B.n90 163.367
R493 B.n162 B.n161 163.367
R494 B.n163 B.n162 163.367
R495 B.n163 B.n88 163.367
R496 B.n167 B.n88 163.367
R497 B.n168 B.n167 163.367
R498 B.n169 B.n168 163.367
R499 B.n169 B.n84 163.367
R500 B.n174 B.n84 163.367
R501 B.n175 B.n174 163.367
R502 B.n176 B.n175 163.367
R503 B.n176 B.n82 163.367
R504 B.n180 B.n82 163.367
R505 B.n181 B.n180 163.367
R506 B.n182 B.n181 163.367
R507 B.n182 B.n80 163.367
R508 B.n186 B.n80 163.367
R509 B.n187 B.n186 163.367
R510 B.n187 B.n76 163.367
R511 B.n191 B.n76 163.367
R512 B.n192 B.n191 163.367
R513 B.n193 B.n192 163.367
R514 B.n193 B.n74 163.367
R515 B.n197 B.n74 163.367
R516 B.n198 B.n197 163.367
R517 B.n199 B.n198 163.367
R518 B.n199 B.n72 163.367
R519 B.n203 B.n72 163.367
R520 B.n204 B.n203 163.367
R521 B.n205 B.n204 163.367
R522 B.n205 B.n70 163.367
R523 B.n209 B.n70 163.367
R524 B.n210 B.n209 163.367
R525 B.n211 B.n210 163.367
R526 B.n211 B.n68 163.367
R527 B.n215 B.n68 163.367
R528 B.n216 B.n215 163.367
R529 B.n217 B.n66 163.367
R530 B.n221 B.n66 163.367
R531 B.n222 B.n221 163.367
R532 B.n223 B.n222 163.367
R533 B.n223 B.n64 163.367
R534 B.n227 B.n64 163.367
R535 B.n228 B.n227 163.367
R536 B.n229 B.n228 163.367
R537 B.n229 B.n62 163.367
R538 B.n233 B.n62 163.367
R539 B.n234 B.n233 163.367
R540 B.n235 B.n234 163.367
R541 B.n235 B.n60 163.367
R542 B.n239 B.n60 163.367
R543 B.n240 B.n239 163.367
R544 B.n241 B.n240 163.367
R545 B.n241 B.n58 163.367
R546 B.n245 B.n58 163.367
R547 B.n246 B.n245 163.367
R548 B.n247 B.n246 163.367
R549 B.n247 B.n56 163.367
R550 B.n251 B.n56 163.367
R551 B.n252 B.n251 163.367
R552 B.n253 B.n252 163.367
R553 B.n253 B.n54 163.367
R554 B.n257 B.n54 163.367
R555 B.n258 B.n257 163.367
R556 B.n259 B.n258 163.367
R557 B.n259 B.n52 163.367
R558 B.n263 B.n52 163.367
R559 B.n264 B.n263 163.367
R560 B.n265 B.n264 163.367
R561 B.n265 B.n50 163.367
R562 B.n269 B.n50 163.367
R563 B.n270 B.n269 163.367
R564 B.n271 B.n270 163.367
R565 B.n271 B.n48 163.367
R566 B.n275 B.n48 163.367
R567 B.n276 B.n275 163.367
R568 B.n277 B.n276 163.367
R569 B.n277 B.n46 163.367
R570 B.n281 B.n46 163.367
R571 B.n282 B.n281 163.367
R572 B.n283 B.n282 163.367
R573 B.n283 B.n44 163.367
R574 B.n287 B.n44 163.367
R575 B.n362 B.n361 163.367
R576 B.n361 B.n360 163.367
R577 B.n360 B.n15 163.367
R578 B.n356 B.n15 163.367
R579 B.n356 B.n355 163.367
R580 B.n355 B.n354 163.367
R581 B.n354 B.n17 163.367
R582 B.n350 B.n17 163.367
R583 B.n350 B.n349 163.367
R584 B.n349 B.n348 163.367
R585 B.n348 B.n19 163.367
R586 B.n344 B.n19 163.367
R587 B.n344 B.n343 163.367
R588 B.n343 B.n342 163.367
R589 B.n342 B.n21 163.367
R590 B.n338 B.n21 163.367
R591 B.n338 B.n337 163.367
R592 B.n337 B.n336 163.367
R593 B.n336 B.n23 163.367
R594 B.n331 B.n23 163.367
R595 B.n331 B.n330 163.367
R596 B.n330 B.n329 163.367
R597 B.n329 B.n27 163.367
R598 B.n325 B.n27 163.367
R599 B.n325 B.n324 163.367
R600 B.n324 B.n323 163.367
R601 B.n323 B.n29 163.367
R602 B.n319 B.n29 163.367
R603 B.n319 B.n318 163.367
R604 B.n318 B.n317 163.367
R605 B.n317 B.n31 163.367
R606 B.n313 B.n31 163.367
R607 B.n313 B.n312 163.367
R608 B.n312 B.n311 163.367
R609 B.n311 B.n36 163.367
R610 B.n307 B.n36 163.367
R611 B.n307 B.n306 163.367
R612 B.n306 B.n305 163.367
R613 B.n305 B.n38 163.367
R614 B.n301 B.n38 163.367
R615 B.n301 B.n300 163.367
R616 B.n300 B.n299 163.367
R617 B.n299 B.n40 163.367
R618 B.n295 B.n40 163.367
R619 B.n295 B.n294 163.367
R620 B.n294 B.n293 163.367
R621 B.n293 B.n42 163.367
R622 B.n289 B.n42 163.367
R623 B.n289 B.n288 163.367
R624 B.n79 B.n78 59.5399
R625 B.n171 B.n86 59.5399
R626 B.n333 B.n25 59.5399
R627 B.n34 B.n33 59.5399
R628 B.n78 B.n77 49.8429
R629 B.n86 B.n85 49.8429
R630 B.n25 B.n24 49.8429
R631 B.n33 B.n32 49.8429
R632 B.n364 B.n363 35.1225
R633 B.n286 B.n43 35.1225
R634 B.n218 B.n67 35.1225
R635 B.n141 B.n140 35.1225
R636 B B.n399 18.0485
R637 B.n363 B.n14 10.6151
R638 B.n359 B.n14 10.6151
R639 B.n359 B.n358 10.6151
R640 B.n358 B.n357 10.6151
R641 B.n357 B.n16 10.6151
R642 B.n353 B.n16 10.6151
R643 B.n353 B.n352 10.6151
R644 B.n352 B.n351 10.6151
R645 B.n351 B.n18 10.6151
R646 B.n347 B.n18 10.6151
R647 B.n347 B.n346 10.6151
R648 B.n346 B.n345 10.6151
R649 B.n345 B.n20 10.6151
R650 B.n341 B.n20 10.6151
R651 B.n341 B.n340 10.6151
R652 B.n340 B.n339 10.6151
R653 B.n339 B.n22 10.6151
R654 B.n335 B.n22 10.6151
R655 B.n335 B.n334 10.6151
R656 B.n332 B.n26 10.6151
R657 B.n328 B.n26 10.6151
R658 B.n328 B.n327 10.6151
R659 B.n327 B.n326 10.6151
R660 B.n326 B.n28 10.6151
R661 B.n322 B.n28 10.6151
R662 B.n322 B.n321 10.6151
R663 B.n321 B.n320 10.6151
R664 B.n320 B.n30 10.6151
R665 B.n316 B.n315 10.6151
R666 B.n315 B.n314 10.6151
R667 B.n314 B.n35 10.6151
R668 B.n310 B.n35 10.6151
R669 B.n310 B.n309 10.6151
R670 B.n309 B.n308 10.6151
R671 B.n308 B.n37 10.6151
R672 B.n304 B.n37 10.6151
R673 B.n304 B.n303 10.6151
R674 B.n303 B.n302 10.6151
R675 B.n302 B.n39 10.6151
R676 B.n298 B.n39 10.6151
R677 B.n298 B.n297 10.6151
R678 B.n297 B.n296 10.6151
R679 B.n296 B.n41 10.6151
R680 B.n292 B.n41 10.6151
R681 B.n292 B.n291 10.6151
R682 B.n291 B.n290 10.6151
R683 B.n290 B.n43 10.6151
R684 B.n219 B.n218 10.6151
R685 B.n220 B.n219 10.6151
R686 B.n220 B.n65 10.6151
R687 B.n224 B.n65 10.6151
R688 B.n225 B.n224 10.6151
R689 B.n226 B.n225 10.6151
R690 B.n226 B.n63 10.6151
R691 B.n230 B.n63 10.6151
R692 B.n231 B.n230 10.6151
R693 B.n232 B.n231 10.6151
R694 B.n232 B.n61 10.6151
R695 B.n236 B.n61 10.6151
R696 B.n237 B.n236 10.6151
R697 B.n238 B.n237 10.6151
R698 B.n238 B.n59 10.6151
R699 B.n242 B.n59 10.6151
R700 B.n243 B.n242 10.6151
R701 B.n244 B.n243 10.6151
R702 B.n244 B.n57 10.6151
R703 B.n248 B.n57 10.6151
R704 B.n249 B.n248 10.6151
R705 B.n250 B.n249 10.6151
R706 B.n250 B.n55 10.6151
R707 B.n254 B.n55 10.6151
R708 B.n255 B.n254 10.6151
R709 B.n256 B.n255 10.6151
R710 B.n256 B.n53 10.6151
R711 B.n260 B.n53 10.6151
R712 B.n261 B.n260 10.6151
R713 B.n262 B.n261 10.6151
R714 B.n262 B.n51 10.6151
R715 B.n266 B.n51 10.6151
R716 B.n267 B.n266 10.6151
R717 B.n268 B.n267 10.6151
R718 B.n268 B.n49 10.6151
R719 B.n272 B.n49 10.6151
R720 B.n273 B.n272 10.6151
R721 B.n274 B.n273 10.6151
R722 B.n274 B.n47 10.6151
R723 B.n278 B.n47 10.6151
R724 B.n279 B.n278 10.6151
R725 B.n280 B.n279 10.6151
R726 B.n280 B.n45 10.6151
R727 B.n284 B.n45 10.6151
R728 B.n285 B.n284 10.6151
R729 B.n286 B.n285 10.6151
R730 B.n142 B.n141 10.6151
R731 B.n142 B.n95 10.6151
R732 B.n146 B.n95 10.6151
R733 B.n147 B.n146 10.6151
R734 B.n148 B.n147 10.6151
R735 B.n148 B.n93 10.6151
R736 B.n152 B.n93 10.6151
R737 B.n153 B.n152 10.6151
R738 B.n154 B.n153 10.6151
R739 B.n154 B.n91 10.6151
R740 B.n158 B.n91 10.6151
R741 B.n159 B.n158 10.6151
R742 B.n160 B.n159 10.6151
R743 B.n160 B.n89 10.6151
R744 B.n164 B.n89 10.6151
R745 B.n165 B.n164 10.6151
R746 B.n166 B.n165 10.6151
R747 B.n166 B.n87 10.6151
R748 B.n170 B.n87 10.6151
R749 B.n173 B.n172 10.6151
R750 B.n173 B.n83 10.6151
R751 B.n177 B.n83 10.6151
R752 B.n178 B.n177 10.6151
R753 B.n179 B.n178 10.6151
R754 B.n179 B.n81 10.6151
R755 B.n183 B.n81 10.6151
R756 B.n184 B.n183 10.6151
R757 B.n185 B.n184 10.6151
R758 B.n189 B.n188 10.6151
R759 B.n190 B.n189 10.6151
R760 B.n190 B.n75 10.6151
R761 B.n194 B.n75 10.6151
R762 B.n195 B.n194 10.6151
R763 B.n196 B.n195 10.6151
R764 B.n196 B.n73 10.6151
R765 B.n200 B.n73 10.6151
R766 B.n201 B.n200 10.6151
R767 B.n202 B.n201 10.6151
R768 B.n202 B.n71 10.6151
R769 B.n206 B.n71 10.6151
R770 B.n207 B.n206 10.6151
R771 B.n208 B.n207 10.6151
R772 B.n208 B.n69 10.6151
R773 B.n212 B.n69 10.6151
R774 B.n213 B.n212 10.6151
R775 B.n214 B.n213 10.6151
R776 B.n214 B.n67 10.6151
R777 B.n140 B.n97 10.6151
R778 B.n136 B.n97 10.6151
R779 B.n136 B.n135 10.6151
R780 B.n135 B.n134 10.6151
R781 B.n134 B.n99 10.6151
R782 B.n130 B.n99 10.6151
R783 B.n130 B.n129 10.6151
R784 B.n129 B.n128 10.6151
R785 B.n128 B.n101 10.6151
R786 B.n124 B.n101 10.6151
R787 B.n124 B.n123 10.6151
R788 B.n123 B.n122 10.6151
R789 B.n122 B.n103 10.6151
R790 B.n118 B.n103 10.6151
R791 B.n118 B.n117 10.6151
R792 B.n117 B.n116 10.6151
R793 B.n116 B.n105 10.6151
R794 B.n112 B.n105 10.6151
R795 B.n112 B.n111 10.6151
R796 B.n111 B.n110 10.6151
R797 B.n110 B.n107 10.6151
R798 B.n107 B.n0 10.6151
R799 B.n395 B.n1 10.6151
R800 B.n395 B.n394 10.6151
R801 B.n394 B.n393 10.6151
R802 B.n393 B.n4 10.6151
R803 B.n389 B.n4 10.6151
R804 B.n389 B.n388 10.6151
R805 B.n388 B.n387 10.6151
R806 B.n387 B.n6 10.6151
R807 B.n383 B.n6 10.6151
R808 B.n383 B.n382 10.6151
R809 B.n382 B.n381 10.6151
R810 B.n381 B.n8 10.6151
R811 B.n377 B.n8 10.6151
R812 B.n377 B.n376 10.6151
R813 B.n376 B.n375 10.6151
R814 B.n375 B.n10 10.6151
R815 B.n371 B.n10 10.6151
R816 B.n371 B.n370 10.6151
R817 B.n370 B.n369 10.6151
R818 B.n369 B.n12 10.6151
R819 B.n365 B.n12 10.6151
R820 B.n365 B.n364 10.6151
R821 B.n334 B.n333 9.36635
R822 B.n316 B.n34 9.36635
R823 B.n171 B.n170 9.36635
R824 B.n188 B.n79 9.36635
R825 B.n399 B.n0 2.81026
R826 B.n399 B.n1 2.81026
R827 B.n333 B.n332 1.24928
R828 B.n34 B.n30 1.24928
R829 B.n172 B.n171 1.24928
R830 B.n185 B.n79 1.24928
R831 VN VN.t0 138.351
R832 VN VN.t1 100.397
R833 VDD2.n41 VDD2.n23 756.745
R834 VDD2.n18 VDD2.n0 756.745
R835 VDD2.n42 VDD2.n41 585
R836 VDD2.n40 VDD2.n39 585
R837 VDD2.n27 VDD2.n26 585
R838 VDD2.n34 VDD2.n33 585
R839 VDD2.n32 VDD2.n31 585
R840 VDD2.n9 VDD2.n8 585
R841 VDD2.n11 VDD2.n10 585
R842 VDD2.n4 VDD2.n3 585
R843 VDD2.n17 VDD2.n16 585
R844 VDD2.n19 VDD2.n18 585
R845 VDD2.n30 VDD2.t1 328.587
R846 VDD2.n7 VDD2.t0 328.587
R847 VDD2.n41 VDD2.n40 171.744
R848 VDD2.n40 VDD2.n26 171.744
R849 VDD2.n33 VDD2.n26 171.744
R850 VDD2.n33 VDD2.n32 171.744
R851 VDD2.n10 VDD2.n9 171.744
R852 VDD2.n10 VDD2.n3 171.744
R853 VDD2.n17 VDD2.n3 171.744
R854 VDD2.n18 VDD2.n17 171.744
R855 VDD2.n32 VDD2.t1 85.8723
R856 VDD2.n9 VDD2.t0 85.8723
R857 VDD2.n46 VDD2.n22 84.3292
R858 VDD2.n46 VDD2.n45 52.1611
R859 VDD2.n31 VDD2.n30 16.3651
R860 VDD2.n8 VDD2.n7 16.3651
R861 VDD2.n34 VDD2.n29 12.8005
R862 VDD2.n11 VDD2.n6 12.8005
R863 VDD2.n35 VDD2.n27 12.0247
R864 VDD2.n12 VDD2.n4 12.0247
R865 VDD2.n39 VDD2.n38 11.249
R866 VDD2.n16 VDD2.n15 11.249
R867 VDD2.n42 VDD2.n25 10.4732
R868 VDD2.n19 VDD2.n2 10.4732
R869 VDD2.n43 VDD2.n23 9.69747
R870 VDD2.n20 VDD2.n0 9.69747
R871 VDD2.n45 VDD2.n44 9.45567
R872 VDD2.n22 VDD2.n21 9.45567
R873 VDD2.n44 VDD2.n43 9.3005
R874 VDD2.n25 VDD2.n24 9.3005
R875 VDD2.n38 VDD2.n37 9.3005
R876 VDD2.n36 VDD2.n35 9.3005
R877 VDD2.n29 VDD2.n28 9.3005
R878 VDD2.n21 VDD2.n20 9.3005
R879 VDD2.n2 VDD2.n1 9.3005
R880 VDD2.n15 VDD2.n14 9.3005
R881 VDD2.n13 VDD2.n12 9.3005
R882 VDD2.n6 VDD2.n5 9.3005
R883 VDD2.n45 VDD2.n23 4.26717
R884 VDD2.n22 VDD2.n0 4.26717
R885 VDD2.n30 VDD2.n28 3.73474
R886 VDD2.n7 VDD2.n5 3.73474
R887 VDD2.n43 VDD2.n42 3.49141
R888 VDD2.n20 VDD2.n19 3.49141
R889 VDD2.n39 VDD2.n25 2.71565
R890 VDD2.n16 VDD2.n2 2.71565
R891 VDD2.n38 VDD2.n27 1.93989
R892 VDD2.n15 VDD2.n4 1.93989
R893 VDD2.n35 VDD2.n34 1.16414
R894 VDD2.n12 VDD2.n11 1.16414
R895 VDD2 VDD2.n46 0.612569
R896 VDD2.n31 VDD2.n29 0.388379
R897 VDD2.n8 VDD2.n6 0.388379
R898 VDD2.n44 VDD2.n24 0.155672
R899 VDD2.n37 VDD2.n24 0.155672
R900 VDD2.n37 VDD2.n36 0.155672
R901 VDD2.n36 VDD2.n28 0.155672
R902 VDD2.n13 VDD2.n5 0.155672
R903 VDD2.n14 VDD2.n13 0.155672
R904 VDD2.n14 VDD2.n1 0.155672
R905 VDD2.n21 VDD2.n1 0.155672
C0 VTAIL B 1.9001f
C1 w_n1998_n1914# VN 2.59668f
C2 VTAIL VP 1.28722f
C3 w_n1998_n1914# B 6.39261f
C4 w_n1998_n1914# VP 2.85031f
C5 VDD2 VTAIL 3.10282f
C6 VDD2 w_n1998_n1914# 1.25232f
C7 VN B 0.902242f
C8 VP VN 3.9427f
C9 VP B 1.31786f
C10 VDD2 VN 1.2227f
C11 VDD2 B 1.11479f
C12 VDD2 VP 0.321505f
C13 VTAIL VDD1 3.05311f
C14 VDD1 w_n1998_n1914# 1.23109f
C15 VTAIL w_n1998_n1914# 1.71054f
C16 VDD1 VN 0.151829f
C17 VDD1 B 1.0878f
C18 VDD1 VP 1.39072f
C19 VDD2 VDD1 0.630651f
C20 VTAIL VN 1.27303f
C21 VDD2 VSUBS 0.591839f
C22 VDD1 VSUBS 2.19299f
C23 VTAIL VSUBS 0.445466f
C24 VN VSUBS 5.13029f
C25 VP VSUBS 1.203605f
C26 B VSUBS 2.878292f
C27 w_n1998_n1914# VSUBS 47.976f
C28 VDD2.n0 VSUBS 0.01719f
C29 VDD2.n1 VSUBS 0.015175f
C30 VDD2.n2 VSUBS 0.008155f
C31 VDD2.n3 VSUBS 0.019274f
C32 VDD2.n4 VSUBS 0.008634f
C33 VDD2.n5 VSUBS 0.258914f
C34 VDD2.n6 VSUBS 0.008155f
C35 VDD2.t0 VSUBS 0.04226f
C36 VDD2.n7 VSUBS 0.062211f
C37 VDD2.n8 VSUBS 0.012211f
C38 VDD2.n9 VSUBS 0.014456f
C39 VDD2.n10 VSUBS 0.019274f
C40 VDD2.n11 VSUBS 0.008634f
C41 VDD2.n12 VSUBS 0.008155f
C42 VDD2.n13 VSUBS 0.015175f
C43 VDD2.n14 VSUBS 0.015175f
C44 VDD2.n15 VSUBS 0.008155f
C45 VDD2.n16 VSUBS 0.008634f
C46 VDD2.n17 VSUBS 0.019274f
C47 VDD2.n18 VSUBS 0.048417f
C48 VDD2.n19 VSUBS 0.008634f
C49 VDD2.n20 VSUBS 0.008155f
C50 VDD2.n21 VSUBS 0.038601f
C51 VDD2.n22 VSUBS 0.280833f
C52 VDD2.n23 VSUBS 0.01719f
C53 VDD2.n24 VSUBS 0.015175f
C54 VDD2.n25 VSUBS 0.008155f
C55 VDD2.n26 VSUBS 0.019274f
C56 VDD2.n27 VSUBS 0.008634f
C57 VDD2.n28 VSUBS 0.258914f
C58 VDD2.n29 VSUBS 0.008155f
C59 VDD2.t1 VSUBS 0.04226f
C60 VDD2.n30 VSUBS 0.062211f
C61 VDD2.n31 VSUBS 0.012211f
C62 VDD2.n32 VSUBS 0.014456f
C63 VDD2.n33 VSUBS 0.019274f
C64 VDD2.n34 VSUBS 0.008634f
C65 VDD2.n35 VSUBS 0.008155f
C66 VDD2.n36 VSUBS 0.015175f
C67 VDD2.n37 VSUBS 0.015175f
C68 VDD2.n38 VSUBS 0.008155f
C69 VDD2.n39 VSUBS 0.008634f
C70 VDD2.n40 VSUBS 0.019274f
C71 VDD2.n41 VSUBS 0.048417f
C72 VDD2.n42 VSUBS 0.008634f
C73 VDD2.n43 VSUBS 0.008155f
C74 VDD2.n44 VSUBS 0.038601f
C75 VDD2.n45 VSUBS 0.034984f
C76 VDD2.n46 VSUBS 1.35383f
C77 VN.t1 VSUBS 1.38407f
C78 VN.t0 VSUBS 1.89095f
C79 B.n0 VSUBS 0.004212f
C80 B.n1 VSUBS 0.004212f
C81 B.n2 VSUBS 0.006661f
C82 B.n3 VSUBS 0.006661f
C83 B.n4 VSUBS 0.006661f
C84 B.n5 VSUBS 0.006661f
C85 B.n6 VSUBS 0.006661f
C86 B.n7 VSUBS 0.006661f
C87 B.n8 VSUBS 0.006661f
C88 B.n9 VSUBS 0.006661f
C89 B.n10 VSUBS 0.006661f
C90 B.n11 VSUBS 0.006661f
C91 B.n12 VSUBS 0.006661f
C92 B.n13 VSUBS 0.015885f
C93 B.n14 VSUBS 0.006661f
C94 B.n15 VSUBS 0.006661f
C95 B.n16 VSUBS 0.006661f
C96 B.n17 VSUBS 0.006661f
C97 B.n18 VSUBS 0.006661f
C98 B.n19 VSUBS 0.006661f
C99 B.n20 VSUBS 0.006661f
C100 B.n21 VSUBS 0.006661f
C101 B.n22 VSUBS 0.006661f
C102 B.n23 VSUBS 0.006661f
C103 B.t8 VSUBS 0.065551f
C104 B.t7 VSUBS 0.084676f
C105 B.t6 VSUBS 0.478729f
C106 B.n24 VSUBS 0.14772f
C107 B.n25 VSUBS 0.12335f
C108 B.n26 VSUBS 0.006661f
C109 B.n27 VSUBS 0.006661f
C110 B.n28 VSUBS 0.006661f
C111 B.n29 VSUBS 0.006661f
C112 B.n30 VSUBS 0.003722f
C113 B.n31 VSUBS 0.006661f
C114 B.t5 VSUBS 0.065552f
C115 B.t4 VSUBS 0.084677f
C116 B.t3 VSUBS 0.478729f
C117 B.n32 VSUBS 0.147719f
C118 B.n33 VSUBS 0.123349f
C119 B.n34 VSUBS 0.015432f
C120 B.n35 VSUBS 0.006661f
C121 B.n36 VSUBS 0.006661f
C122 B.n37 VSUBS 0.006661f
C123 B.n38 VSUBS 0.006661f
C124 B.n39 VSUBS 0.006661f
C125 B.n40 VSUBS 0.006661f
C126 B.n41 VSUBS 0.006661f
C127 B.n42 VSUBS 0.006661f
C128 B.n43 VSUBS 0.016099f
C129 B.n44 VSUBS 0.006661f
C130 B.n45 VSUBS 0.006661f
C131 B.n46 VSUBS 0.006661f
C132 B.n47 VSUBS 0.006661f
C133 B.n48 VSUBS 0.006661f
C134 B.n49 VSUBS 0.006661f
C135 B.n50 VSUBS 0.006661f
C136 B.n51 VSUBS 0.006661f
C137 B.n52 VSUBS 0.006661f
C138 B.n53 VSUBS 0.006661f
C139 B.n54 VSUBS 0.006661f
C140 B.n55 VSUBS 0.006661f
C141 B.n56 VSUBS 0.006661f
C142 B.n57 VSUBS 0.006661f
C143 B.n58 VSUBS 0.006661f
C144 B.n59 VSUBS 0.006661f
C145 B.n60 VSUBS 0.006661f
C146 B.n61 VSUBS 0.006661f
C147 B.n62 VSUBS 0.006661f
C148 B.n63 VSUBS 0.006661f
C149 B.n64 VSUBS 0.006661f
C150 B.n65 VSUBS 0.006661f
C151 B.n66 VSUBS 0.006661f
C152 B.n67 VSUBS 0.016831f
C153 B.n68 VSUBS 0.006661f
C154 B.n69 VSUBS 0.006661f
C155 B.n70 VSUBS 0.006661f
C156 B.n71 VSUBS 0.006661f
C157 B.n72 VSUBS 0.006661f
C158 B.n73 VSUBS 0.006661f
C159 B.n74 VSUBS 0.006661f
C160 B.n75 VSUBS 0.006661f
C161 B.n76 VSUBS 0.006661f
C162 B.t10 VSUBS 0.065552f
C163 B.t11 VSUBS 0.084677f
C164 B.t9 VSUBS 0.478729f
C165 B.n77 VSUBS 0.147719f
C166 B.n78 VSUBS 0.123349f
C167 B.n79 VSUBS 0.015432f
C168 B.n80 VSUBS 0.006661f
C169 B.n81 VSUBS 0.006661f
C170 B.n82 VSUBS 0.006661f
C171 B.n83 VSUBS 0.006661f
C172 B.n84 VSUBS 0.006661f
C173 B.t1 VSUBS 0.065551f
C174 B.t2 VSUBS 0.084676f
C175 B.t0 VSUBS 0.478729f
C176 B.n85 VSUBS 0.14772f
C177 B.n86 VSUBS 0.12335f
C178 B.n87 VSUBS 0.006661f
C179 B.n88 VSUBS 0.006661f
C180 B.n89 VSUBS 0.006661f
C181 B.n90 VSUBS 0.006661f
C182 B.n91 VSUBS 0.006661f
C183 B.n92 VSUBS 0.006661f
C184 B.n93 VSUBS 0.006661f
C185 B.n94 VSUBS 0.006661f
C186 B.n95 VSUBS 0.006661f
C187 B.n96 VSUBS 0.016831f
C188 B.n97 VSUBS 0.006661f
C189 B.n98 VSUBS 0.006661f
C190 B.n99 VSUBS 0.006661f
C191 B.n100 VSUBS 0.006661f
C192 B.n101 VSUBS 0.006661f
C193 B.n102 VSUBS 0.006661f
C194 B.n103 VSUBS 0.006661f
C195 B.n104 VSUBS 0.006661f
C196 B.n105 VSUBS 0.006661f
C197 B.n106 VSUBS 0.006661f
C198 B.n107 VSUBS 0.006661f
C199 B.n108 VSUBS 0.006661f
C200 B.n109 VSUBS 0.006661f
C201 B.n110 VSUBS 0.006661f
C202 B.n111 VSUBS 0.006661f
C203 B.n112 VSUBS 0.006661f
C204 B.n113 VSUBS 0.006661f
C205 B.n114 VSUBS 0.006661f
C206 B.n115 VSUBS 0.006661f
C207 B.n116 VSUBS 0.006661f
C208 B.n117 VSUBS 0.006661f
C209 B.n118 VSUBS 0.006661f
C210 B.n119 VSUBS 0.006661f
C211 B.n120 VSUBS 0.006661f
C212 B.n121 VSUBS 0.006661f
C213 B.n122 VSUBS 0.006661f
C214 B.n123 VSUBS 0.006661f
C215 B.n124 VSUBS 0.006661f
C216 B.n125 VSUBS 0.006661f
C217 B.n126 VSUBS 0.006661f
C218 B.n127 VSUBS 0.006661f
C219 B.n128 VSUBS 0.006661f
C220 B.n129 VSUBS 0.006661f
C221 B.n130 VSUBS 0.006661f
C222 B.n131 VSUBS 0.006661f
C223 B.n132 VSUBS 0.006661f
C224 B.n133 VSUBS 0.006661f
C225 B.n134 VSUBS 0.006661f
C226 B.n135 VSUBS 0.006661f
C227 B.n136 VSUBS 0.006661f
C228 B.n137 VSUBS 0.006661f
C229 B.n138 VSUBS 0.006661f
C230 B.n139 VSUBS 0.015885f
C231 B.n140 VSUBS 0.015885f
C232 B.n141 VSUBS 0.016831f
C233 B.n142 VSUBS 0.006661f
C234 B.n143 VSUBS 0.006661f
C235 B.n144 VSUBS 0.006661f
C236 B.n145 VSUBS 0.006661f
C237 B.n146 VSUBS 0.006661f
C238 B.n147 VSUBS 0.006661f
C239 B.n148 VSUBS 0.006661f
C240 B.n149 VSUBS 0.006661f
C241 B.n150 VSUBS 0.006661f
C242 B.n151 VSUBS 0.006661f
C243 B.n152 VSUBS 0.006661f
C244 B.n153 VSUBS 0.006661f
C245 B.n154 VSUBS 0.006661f
C246 B.n155 VSUBS 0.006661f
C247 B.n156 VSUBS 0.006661f
C248 B.n157 VSUBS 0.006661f
C249 B.n158 VSUBS 0.006661f
C250 B.n159 VSUBS 0.006661f
C251 B.n160 VSUBS 0.006661f
C252 B.n161 VSUBS 0.006661f
C253 B.n162 VSUBS 0.006661f
C254 B.n163 VSUBS 0.006661f
C255 B.n164 VSUBS 0.006661f
C256 B.n165 VSUBS 0.006661f
C257 B.n166 VSUBS 0.006661f
C258 B.n167 VSUBS 0.006661f
C259 B.n168 VSUBS 0.006661f
C260 B.n169 VSUBS 0.006661f
C261 B.n170 VSUBS 0.006269f
C262 B.n171 VSUBS 0.015432f
C263 B.n172 VSUBS 0.003722f
C264 B.n173 VSUBS 0.006661f
C265 B.n174 VSUBS 0.006661f
C266 B.n175 VSUBS 0.006661f
C267 B.n176 VSUBS 0.006661f
C268 B.n177 VSUBS 0.006661f
C269 B.n178 VSUBS 0.006661f
C270 B.n179 VSUBS 0.006661f
C271 B.n180 VSUBS 0.006661f
C272 B.n181 VSUBS 0.006661f
C273 B.n182 VSUBS 0.006661f
C274 B.n183 VSUBS 0.006661f
C275 B.n184 VSUBS 0.006661f
C276 B.n185 VSUBS 0.003722f
C277 B.n186 VSUBS 0.006661f
C278 B.n187 VSUBS 0.006661f
C279 B.n188 VSUBS 0.006269f
C280 B.n189 VSUBS 0.006661f
C281 B.n190 VSUBS 0.006661f
C282 B.n191 VSUBS 0.006661f
C283 B.n192 VSUBS 0.006661f
C284 B.n193 VSUBS 0.006661f
C285 B.n194 VSUBS 0.006661f
C286 B.n195 VSUBS 0.006661f
C287 B.n196 VSUBS 0.006661f
C288 B.n197 VSUBS 0.006661f
C289 B.n198 VSUBS 0.006661f
C290 B.n199 VSUBS 0.006661f
C291 B.n200 VSUBS 0.006661f
C292 B.n201 VSUBS 0.006661f
C293 B.n202 VSUBS 0.006661f
C294 B.n203 VSUBS 0.006661f
C295 B.n204 VSUBS 0.006661f
C296 B.n205 VSUBS 0.006661f
C297 B.n206 VSUBS 0.006661f
C298 B.n207 VSUBS 0.006661f
C299 B.n208 VSUBS 0.006661f
C300 B.n209 VSUBS 0.006661f
C301 B.n210 VSUBS 0.006661f
C302 B.n211 VSUBS 0.006661f
C303 B.n212 VSUBS 0.006661f
C304 B.n213 VSUBS 0.006661f
C305 B.n214 VSUBS 0.006661f
C306 B.n215 VSUBS 0.006661f
C307 B.n216 VSUBS 0.016831f
C308 B.n217 VSUBS 0.015885f
C309 B.n218 VSUBS 0.015885f
C310 B.n219 VSUBS 0.006661f
C311 B.n220 VSUBS 0.006661f
C312 B.n221 VSUBS 0.006661f
C313 B.n222 VSUBS 0.006661f
C314 B.n223 VSUBS 0.006661f
C315 B.n224 VSUBS 0.006661f
C316 B.n225 VSUBS 0.006661f
C317 B.n226 VSUBS 0.006661f
C318 B.n227 VSUBS 0.006661f
C319 B.n228 VSUBS 0.006661f
C320 B.n229 VSUBS 0.006661f
C321 B.n230 VSUBS 0.006661f
C322 B.n231 VSUBS 0.006661f
C323 B.n232 VSUBS 0.006661f
C324 B.n233 VSUBS 0.006661f
C325 B.n234 VSUBS 0.006661f
C326 B.n235 VSUBS 0.006661f
C327 B.n236 VSUBS 0.006661f
C328 B.n237 VSUBS 0.006661f
C329 B.n238 VSUBS 0.006661f
C330 B.n239 VSUBS 0.006661f
C331 B.n240 VSUBS 0.006661f
C332 B.n241 VSUBS 0.006661f
C333 B.n242 VSUBS 0.006661f
C334 B.n243 VSUBS 0.006661f
C335 B.n244 VSUBS 0.006661f
C336 B.n245 VSUBS 0.006661f
C337 B.n246 VSUBS 0.006661f
C338 B.n247 VSUBS 0.006661f
C339 B.n248 VSUBS 0.006661f
C340 B.n249 VSUBS 0.006661f
C341 B.n250 VSUBS 0.006661f
C342 B.n251 VSUBS 0.006661f
C343 B.n252 VSUBS 0.006661f
C344 B.n253 VSUBS 0.006661f
C345 B.n254 VSUBS 0.006661f
C346 B.n255 VSUBS 0.006661f
C347 B.n256 VSUBS 0.006661f
C348 B.n257 VSUBS 0.006661f
C349 B.n258 VSUBS 0.006661f
C350 B.n259 VSUBS 0.006661f
C351 B.n260 VSUBS 0.006661f
C352 B.n261 VSUBS 0.006661f
C353 B.n262 VSUBS 0.006661f
C354 B.n263 VSUBS 0.006661f
C355 B.n264 VSUBS 0.006661f
C356 B.n265 VSUBS 0.006661f
C357 B.n266 VSUBS 0.006661f
C358 B.n267 VSUBS 0.006661f
C359 B.n268 VSUBS 0.006661f
C360 B.n269 VSUBS 0.006661f
C361 B.n270 VSUBS 0.006661f
C362 B.n271 VSUBS 0.006661f
C363 B.n272 VSUBS 0.006661f
C364 B.n273 VSUBS 0.006661f
C365 B.n274 VSUBS 0.006661f
C366 B.n275 VSUBS 0.006661f
C367 B.n276 VSUBS 0.006661f
C368 B.n277 VSUBS 0.006661f
C369 B.n278 VSUBS 0.006661f
C370 B.n279 VSUBS 0.006661f
C371 B.n280 VSUBS 0.006661f
C372 B.n281 VSUBS 0.006661f
C373 B.n282 VSUBS 0.006661f
C374 B.n283 VSUBS 0.006661f
C375 B.n284 VSUBS 0.006661f
C376 B.n285 VSUBS 0.006661f
C377 B.n286 VSUBS 0.016617f
C378 B.n287 VSUBS 0.015885f
C379 B.n288 VSUBS 0.016831f
C380 B.n289 VSUBS 0.006661f
C381 B.n290 VSUBS 0.006661f
C382 B.n291 VSUBS 0.006661f
C383 B.n292 VSUBS 0.006661f
C384 B.n293 VSUBS 0.006661f
C385 B.n294 VSUBS 0.006661f
C386 B.n295 VSUBS 0.006661f
C387 B.n296 VSUBS 0.006661f
C388 B.n297 VSUBS 0.006661f
C389 B.n298 VSUBS 0.006661f
C390 B.n299 VSUBS 0.006661f
C391 B.n300 VSUBS 0.006661f
C392 B.n301 VSUBS 0.006661f
C393 B.n302 VSUBS 0.006661f
C394 B.n303 VSUBS 0.006661f
C395 B.n304 VSUBS 0.006661f
C396 B.n305 VSUBS 0.006661f
C397 B.n306 VSUBS 0.006661f
C398 B.n307 VSUBS 0.006661f
C399 B.n308 VSUBS 0.006661f
C400 B.n309 VSUBS 0.006661f
C401 B.n310 VSUBS 0.006661f
C402 B.n311 VSUBS 0.006661f
C403 B.n312 VSUBS 0.006661f
C404 B.n313 VSUBS 0.006661f
C405 B.n314 VSUBS 0.006661f
C406 B.n315 VSUBS 0.006661f
C407 B.n316 VSUBS 0.006269f
C408 B.n317 VSUBS 0.006661f
C409 B.n318 VSUBS 0.006661f
C410 B.n319 VSUBS 0.006661f
C411 B.n320 VSUBS 0.006661f
C412 B.n321 VSUBS 0.006661f
C413 B.n322 VSUBS 0.006661f
C414 B.n323 VSUBS 0.006661f
C415 B.n324 VSUBS 0.006661f
C416 B.n325 VSUBS 0.006661f
C417 B.n326 VSUBS 0.006661f
C418 B.n327 VSUBS 0.006661f
C419 B.n328 VSUBS 0.006661f
C420 B.n329 VSUBS 0.006661f
C421 B.n330 VSUBS 0.006661f
C422 B.n331 VSUBS 0.006661f
C423 B.n332 VSUBS 0.003722f
C424 B.n333 VSUBS 0.015432f
C425 B.n334 VSUBS 0.006269f
C426 B.n335 VSUBS 0.006661f
C427 B.n336 VSUBS 0.006661f
C428 B.n337 VSUBS 0.006661f
C429 B.n338 VSUBS 0.006661f
C430 B.n339 VSUBS 0.006661f
C431 B.n340 VSUBS 0.006661f
C432 B.n341 VSUBS 0.006661f
C433 B.n342 VSUBS 0.006661f
C434 B.n343 VSUBS 0.006661f
C435 B.n344 VSUBS 0.006661f
C436 B.n345 VSUBS 0.006661f
C437 B.n346 VSUBS 0.006661f
C438 B.n347 VSUBS 0.006661f
C439 B.n348 VSUBS 0.006661f
C440 B.n349 VSUBS 0.006661f
C441 B.n350 VSUBS 0.006661f
C442 B.n351 VSUBS 0.006661f
C443 B.n352 VSUBS 0.006661f
C444 B.n353 VSUBS 0.006661f
C445 B.n354 VSUBS 0.006661f
C446 B.n355 VSUBS 0.006661f
C447 B.n356 VSUBS 0.006661f
C448 B.n357 VSUBS 0.006661f
C449 B.n358 VSUBS 0.006661f
C450 B.n359 VSUBS 0.006661f
C451 B.n360 VSUBS 0.006661f
C452 B.n361 VSUBS 0.006661f
C453 B.n362 VSUBS 0.016831f
C454 B.n363 VSUBS 0.016831f
C455 B.n364 VSUBS 0.015885f
C456 B.n365 VSUBS 0.006661f
C457 B.n366 VSUBS 0.006661f
C458 B.n367 VSUBS 0.006661f
C459 B.n368 VSUBS 0.006661f
C460 B.n369 VSUBS 0.006661f
C461 B.n370 VSUBS 0.006661f
C462 B.n371 VSUBS 0.006661f
C463 B.n372 VSUBS 0.006661f
C464 B.n373 VSUBS 0.006661f
C465 B.n374 VSUBS 0.006661f
C466 B.n375 VSUBS 0.006661f
C467 B.n376 VSUBS 0.006661f
C468 B.n377 VSUBS 0.006661f
C469 B.n378 VSUBS 0.006661f
C470 B.n379 VSUBS 0.006661f
C471 B.n380 VSUBS 0.006661f
C472 B.n381 VSUBS 0.006661f
C473 B.n382 VSUBS 0.006661f
C474 B.n383 VSUBS 0.006661f
C475 B.n384 VSUBS 0.006661f
C476 B.n385 VSUBS 0.006661f
C477 B.n386 VSUBS 0.006661f
C478 B.n387 VSUBS 0.006661f
C479 B.n388 VSUBS 0.006661f
C480 B.n389 VSUBS 0.006661f
C481 B.n390 VSUBS 0.006661f
C482 B.n391 VSUBS 0.006661f
C483 B.n392 VSUBS 0.006661f
C484 B.n393 VSUBS 0.006661f
C485 B.n394 VSUBS 0.006661f
C486 B.n395 VSUBS 0.006661f
C487 B.n396 VSUBS 0.006661f
C488 B.n397 VSUBS 0.006661f
C489 B.n398 VSUBS 0.006661f
C490 B.n399 VSUBS 0.015082f
C491 VDD1.n0 VSUBS 0.016885f
C492 VDD1.n1 VSUBS 0.014906f
C493 VDD1.n2 VSUBS 0.00801f
C494 VDD1.n3 VSUBS 0.018932f
C495 VDD1.n4 VSUBS 0.008481f
C496 VDD1.n5 VSUBS 0.254316f
C497 VDD1.n6 VSUBS 0.00801f
C498 VDD1.t0 VSUBS 0.041509f
C499 VDD1.n7 VSUBS 0.061106f
C500 VDD1.n8 VSUBS 0.011994f
C501 VDD1.n9 VSUBS 0.014199f
C502 VDD1.n10 VSUBS 0.018932f
C503 VDD1.n11 VSUBS 0.008481f
C504 VDD1.n12 VSUBS 0.00801f
C505 VDD1.n13 VSUBS 0.014906f
C506 VDD1.n14 VSUBS 0.014906f
C507 VDD1.n15 VSUBS 0.00801f
C508 VDD1.n16 VSUBS 0.008481f
C509 VDD1.n17 VSUBS 0.018932f
C510 VDD1.n18 VSUBS 0.047557f
C511 VDD1.n19 VSUBS 0.008481f
C512 VDD1.n20 VSUBS 0.00801f
C513 VDD1.n21 VSUBS 0.037916f
C514 VDD1.n22 VSUBS 0.035059f
C515 VDD1.n23 VSUBS 0.016885f
C516 VDD1.n24 VSUBS 0.014906f
C517 VDD1.n25 VSUBS 0.00801f
C518 VDD1.n26 VSUBS 0.018932f
C519 VDD1.n27 VSUBS 0.008481f
C520 VDD1.n28 VSUBS 0.254316f
C521 VDD1.n29 VSUBS 0.00801f
C522 VDD1.t1 VSUBS 0.041509f
C523 VDD1.n30 VSUBS 0.061106f
C524 VDD1.n31 VSUBS 0.011994f
C525 VDD1.n32 VSUBS 0.014199f
C526 VDD1.n33 VSUBS 0.018932f
C527 VDD1.n34 VSUBS 0.008481f
C528 VDD1.n35 VSUBS 0.00801f
C529 VDD1.n36 VSUBS 0.014906f
C530 VDD1.n37 VSUBS 0.014906f
C531 VDD1.n38 VSUBS 0.00801f
C532 VDD1.n39 VSUBS 0.008481f
C533 VDD1.n40 VSUBS 0.018932f
C534 VDD1.n41 VSUBS 0.047557f
C535 VDD1.n42 VSUBS 0.008481f
C536 VDD1.n43 VSUBS 0.00801f
C537 VDD1.n44 VSUBS 0.037916f
C538 VDD1.n45 VSUBS 0.298558f
C539 VTAIL.n0 VSUBS 0.019627f
C540 VTAIL.n1 VSUBS 0.017326f
C541 VTAIL.n2 VSUBS 0.00931f
C542 VTAIL.n3 VSUBS 0.022006f
C543 VTAIL.n4 VSUBS 0.009858f
C544 VTAIL.n5 VSUBS 0.295614f
C545 VTAIL.n6 VSUBS 0.00931f
C546 VTAIL.t2 VSUBS 0.04825f
C547 VTAIL.n7 VSUBS 0.071029f
C548 VTAIL.n8 VSUBS 0.013941f
C549 VTAIL.n9 VSUBS 0.016505f
C550 VTAIL.n10 VSUBS 0.022006f
C551 VTAIL.n11 VSUBS 0.009858f
C552 VTAIL.n12 VSUBS 0.00931f
C553 VTAIL.n13 VSUBS 0.017326f
C554 VTAIL.n14 VSUBS 0.017326f
C555 VTAIL.n15 VSUBS 0.00931f
C556 VTAIL.n16 VSUBS 0.009858f
C557 VTAIL.n17 VSUBS 0.022006f
C558 VTAIL.n18 VSUBS 0.05528f
C559 VTAIL.n19 VSUBS 0.009858f
C560 VTAIL.n20 VSUBS 0.00931f
C561 VTAIL.n21 VSUBS 0.044073f
C562 VTAIL.n22 VSUBS 0.028007f
C563 VTAIL.n23 VSUBS 0.787863f
C564 VTAIL.n24 VSUBS 0.019627f
C565 VTAIL.n25 VSUBS 0.017326f
C566 VTAIL.n26 VSUBS 0.00931f
C567 VTAIL.n27 VSUBS 0.022006f
C568 VTAIL.n28 VSUBS 0.009858f
C569 VTAIL.n29 VSUBS 0.295614f
C570 VTAIL.n30 VSUBS 0.00931f
C571 VTAIL.t0 VSUBS 0.04825f
C572 VTAIL.n31 VSUBS 0.071029f
C573 VTAIL.n32 VSUBS 0.013941f
C574 VTAIL.n33 VSUBS 0.016505f
C575 VTAIL.n34 VSUBS 0.022006f
C576 VTAIL.n35 VSUBS 0.009858f
C577 VTAIL.n36 VSUBS 0.00931f
C578 VTAIL.n37 VSUBS 0.017326f
C579 VTAIL.n38 VSUBS 0.017326f
C580 VTAIL.n39 VSUBS 0.00931f
C581 VTAIL.n40 VSUBS 0.009858f
C582 VTAIL.n41 VSUBS 0.022006f
C583 VTAIL.n42 VSUBS 0.05528f
C584 VTAIL.n43 VSUBS 0.009858f
C585 VTAIL.n44 VSUBS 0.00931f
C586 VTAIL.n45 VSUBS 0.044073f
C587 VTAIL.n46 VSUBS 0.028007f
C588 VTAIL.n47 VSUBS 0.815537f
C589 VTAIL.n48 VSUBS 0.019627f
C590 VTAIL.n49 VSUBS 0.017326f
C591 VTAIL.n50 VSUBS 0.00931f
C592 VTAIL.n51 VSUBS 0.022006f
C593 VTAIL.n52 VSUBS 0.009858f
C594 VTAIL.n53 VSUBS 0.295614f
C595 VTAIL.n54 VSUBS 0.00931f
C596 VTAIL.t3 VSUBS 0.04825f
C597 VTAIL.n55 VSUBS 0.071029f
C598 VTAIL.n56 VSUBS 0.013941f
C599 VTAIL.n57 VSUBS 0.016505f
C600 VTAIL.n58 VSUBS 0.022006f
C601 VTAIL.n59 VSUBS 0.009858f
C602 VTAIL.n60 VSUBS 0.00931f
C603 VTAIL.n61 VSUBS 0.017326f
C604 VTAIL.n62 VSUBS 0.017326f
C605 VTAIL.n63 VSUBS 0.00931f
C606 VTAIL.n64 VSUBS 0.009858f
C607 VTAIL.n65 VSUBS 0.022006f
C608 VTAIL.n66 VSUBS 0.05528f
C609 VTAIL.n67 VSUBS 0.009858f
C610 VTAIL.n68 VSUBS 0.00931f
C611 VTAIL.n69 VSUBS 0.044073f
C612 VTAIL.n70 VSUBS 0.028007f
C613 VTAIL.n71 VSUBS 0.691846f
C614 VTAIL.n72 VSUBS 0.019627f
C615 VTAIL.n73 VSUBS 0.017326f
C616 VTAIL.n74 VSUBS 0.00931f
C617 VTAIL.n75 VSUBS 0.022006f
C618 VTAIL.n76 VSUBS 0.009858f
C619 VTAIL.n77 VSUBS 0.295614f
C620 VTAIL.n78 VSUBS 0.00931f
C621 VTAIL.t1 VSUBS 0.04825f
C622 VTAIL.n79 VSUBS 0.071029f
C623 VTAIL.n80 VSUBS 0.013941f
C624 VTAIL.n81 VSUBS 0.016505f
C625 VTAIL.n82 VSUBS 0.022006f
C626 VTAIL.n83 VSUBS 0.009858f
C627 VTAIL.n84 VSUBS 0.00931f
C628 VTAIL.n85 VSUBS 0.017326f
C629 VTAIL.n86 VSUBS 0.017326f
C630 VTAIL.n87 VSUBS 0.00931f
C631 VTAIL.n88 VSUBS 0.009858f
C632 VTAIL.n89 VSUBS 0.022006f
C633 VTAIL.n90 VSUBS 0.05528f
C634 VTAIL.n91 VSUBS 0.009858f
C635 VTAIL.n92 VSUBS 0.00931f
C636 VTAIL.n93 VSUBS 0.044073f
C637 VTAIL.n94 VSUBS 0.028007f
C638 VTAIL.n95 VSUBS 0.631445f
C639 VP.t1 VSUBS 1.98955f
C640 VP.t0 VSUBS 1.45846f
C641 VP.n0 VSUBS 3.26804f
.ends

