* NGSPICE file created from diff_pair_sample_1296.ext - technology: sky130A

.subckt diff_pair_sample_1296 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.75
X1 VDD1.t5 VP.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.75
X2 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.75
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.75
X4 VTAIL.t2 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.75
X5 VTAIL.t11 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.75
X6 VDD1.t3 VP.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.75
X7 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.75
X8 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.75
X9 VTAIL.t4 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.75
X10 VDD2.t1 VN.t4 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.75
X11 VDD2.t0 VN.t5 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.75
X12 VDD1.t2 VP.t3 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.75
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.75
X14 VDD1.t1 VP.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.75
X15 VTAIL.t8 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.75
R0 B.n673 B.n672 585
R1 B.n674 B.n673 585
R2 B.n237 B.n114 585
R3 B.n236 B.n235 585
R4 B.n234 B.n233 585
R5 B.n232 B.n231 585
R6 B.n230 B.n229 585
R7 B.n228 B.n227 585
R8 B.n226 B.n225 585
R9 B.n224 B.n223 585
R10 B.n222 B.n221 585
R11 B.n220 B.n219 585
R12 B.n218 B.n217 585
R13 B.n216 B.n215 585
R14 B.n214 B.n213 585
R15 B.n212 B.n211 585
R16 B.n210 B.n209 585
R17 B.n208 B.n207 585
R18 B.n206 B.n205 585
R19 B.n204 B.n203 585
R20 B.n202 B.n201 585
R21 B.n200 B.n199 585
R22 B.n198 B.n197 585
R23 B.n196 B.n195 585
R24 B.n194 B.n193 585
R25 B.n192 B.n191 585
R26 B.n190 B.n189 585
R27 B.n187 B.n186 585
R28 B.n185 B.n184 585
R29 B.n183 B.n182 585
R30 B.n181 B.n180 585
R31 B.n179 B.n178 585
R32 B.n177 B.n176 585
R33 B.n175 B.n174 585
R34 B.n173 B.n172 585
R35 B.n171 B.n170 585
R36 B.n169 B.n168 585
R37 B.n167 B.n166 585
R38 B.n165 B.n164 585
R39 B.n163 B.n162 585
R40 B.n161 B.n160 585
R41 B.n159 B.n158 585
R42 B.n157 B.n156 585
R43 B.n155 B.n154 585
R44 B.n153 B.n152 585
R45 B.n151 B.n150 585
R46 B.n149 B.n148 585
R47 B.n147 B.n146 585
R48 B.n145 B.n144 585
R49 B.n143 B.n142 585
R50 B.n141 B.n140 585
R51 B.n139 B.n138 585
R52 B.n137 B.n136 585
R53 B.n135 B.n134 585
R54 B.n133 B.n132 585
R55 B.n131 B.n130 585
R56 B.n129 B.n128 585
R57 B.n127 B.n126 585
R58 B.n125 B.n124 585
R59 B.n123 B.n122 585
R60 B.n121 B.n120 585
R61 B.n82 B.n81 585
R62 B.n671 B.n83 585
R63 B.n675 B.n83 585
R64 B.n670 B.n669 585
R65 B.n669 B.n79 585
R66 B.n668 B.n78 585
R67 B.n681 B.n78 585
R68 B.n667 B.n77 585
R69 B.n682 B.n77 585
R70 B.n666 B.n76 585
R71 B.n683 B.n76 585
R72 B.n665 B.n664 585
R73 B.n664 B.n72 585
R74 B.n663 B.n71 585
R75 B.n689 B.n71 585
R76 B.n662 B.n70 585
R77 B.n690 B.n70 585
R78 B.n661 B.n69 585
R79 B.n691 B.n69 585
R80 B.n660 B.n659 585
R81 B.n659 B.n65 585
R82 B.n658 B.n64 585
R83 B.n697 B.n64 585
R84 B.n657 B.n63 585
R85 B.n698 B.n63 585
R86 B.n656 B.n62 585
R87 B.n699 B.n62 585
R88 B.n655 B.n654 585
R89 B.n654 B.n58 585
R90 B.n653 B.n57 585
R91 B.n705 B.n57 585
R92 B.n652 B.n56 585
R93 B.n706 B.n56 585
R94 B.n651 B.n55 585
R95 B.n707 B.n55 585
R96 B.n650 B.n649 585
R97 B.n649 B.n51 585
R98 B.n648 B.n50 585
R99 B.n713 B.n50 585
R100 B.n647 B.n49 585
R101 B.n714 B.n49 585
R102 B.n646 B.n48 585
R103 B.n715 B.n48 585
R104 B.n645 B.n644 585
R105 B.n644 B.n44 585
R106 B.n643 B.n43 585
R107 B.n721 B.n43 585
R108 B.n642 B.n42 585
R109 B.n722 B.n42 585
R110 B.n641 B.n41 585
R111 B.n723 B.n41 585
R112 B.n640 B.n639 585
R113 B.n639 B.n37 585
R114 B.n638 B.n36 585
R115 B.n729 B.n36 585
R116 B.n637 B.n35 585
R117 B.n730 B.n35 585
R118 B.n636 B.n34 585
R119 B.n731 B.n34 585
R120 B.n635 B.n634 585
R121 B.n634 B.n33 585
R122 B.n633 B.n29 585
R123 B.n737 B.n29 585
R124 B.n632 B.n28 585
R125 B.n738 B.n28 585
R126 B.n631 B.n27 585
R127 B.n739 B.n27 585
R128 B.n630 B.n629 585
R129 B.n629 B.n23 585
R130 B.n628 B.n22 585
R131 B.n745 B.n22 585
R132 B.n627 B.n21 585
R133 B.n746 B.n21 585
R134 B.n626 B.n20 585
R135 B.n747 B.n20 585
R136 B.n625 B.n624 585
R137 B.n624 B.n16 585
R138 B.n623 B.n15 585
R139 B.n753 B.n15 585
R140 B.n622 B.n14 585
R141 B.n754 B.n14 585
R142 B.n621 B.n13 585
R143 B.n755 B.n13 585
R144 B.n620 B.n619 585
R145 B.n619 B.n12 585
R146 B.n618 B.n617 585
R147 B.n618 B.n8 585
R148 B.n616 B.n7 585
R149 B.n762 B.n7 585
R150 B.n615 B.n6 585
R151 B.n763 B.n6 585
R152 B.n614 B.n5 585
R153 B.n764 B.n5 585
R154 B.n613 B.n612 585
R155 B.n612 B.n4 585
R156 B.n611 B.n238 585
R157 B.n611 B.n610 585
R158 B.n601 B.n239 585
R159 B.n240 B.n239 585
R160 B.n603 B.n602 585
R161 B.n604 B.n603 585
R162 B.n600 B.n245 585
R163 B.n245 B.n244 585
R164 B.n599 B.n598 585
R165 B.n598 B.n597 585
R166 B.n247 B.n246 585
R167 B.n248 B.n247 585
R168 B.n590 B.n589 585
R169 B.n591 B.n590 585
R170 B.n588 B.n253 585
R171 B.n253 B.n252 585
R172 B.n587 B.n586 585
R173 B.n586 B.n585 585
R174 B.n255 B.n254 585
R175 B.n256 B.n255 585
R176 B.n578 B.n577 585
R177 B.n579 B.n578 585
R178 B.n576 B.n261 585
R179 B.n261 B.n260 585
R180 B.n575 B.n574 585
R181 B.n574 B.n573 585
R182 B.n263 B.n262 585
R183 B.n566 B.n263 585
R184 B.n565 B.n564 585
R185 B.n567 B.n565 585
R186 B.n563 B.n268 585
R187 B.n268 B.n267 585
R188 B.n562 B.n561 585
R189 B.n561 B.n560 585
R190 B.n270 B.n269 585
R191 B.n271 B.n270 585
R192 B.n553 B.n552 585
R193 B.n554 B.n553 585
R194 B.n551 B.n276 585
R195 B.n276 B.n275 585
R196 B.n550 B.n549 585
R197 B.n549 B.n548 585
R198 B.n278 B.n277 585
R199 B.n279 B.n278 585
R200 B.n541 B.n540 585
R201 B.n542 B.n541 585
R202 B.n539 B.n284 585
R203 B.n284 B.n283 585
R204 B.n538 B.n537 585
R205 B.n537 B.n536 585
R206 B.n286 B.n285 585
R207 B.n287 B.n286 585
R208 B.n529 B.n528 585
R209 B.n530 B.n529 585
R210 B.n527 B.n292 585
R211 B.n292 B.n291 585
R212 B.n526 B.n525 585
R213 B.n525 B.n524 585
R214 B.n294 B.n293 585
R215 B.n295 B.n294 585
R216 B.n517 B.n516 585
R217 B.n518 B.n517 585
R218 B.n515 B.n300 585
R219 B.n300 B.n299 585
R220 B.n514 B.n513 585
R221 B.n513 B.n512 585
R222 B.n302 B.n301 585
R223 B.n303 B.n302 585
R224 B.n505 B.n504 585
R225 B.n506 B.n505 585
R226 B.n503 B.n307 585
R227 B.n311 B.n307 585
R228 B.n502 B.n501 585
R229 B.n501 B.n500 585
R230 B.n309 B.n308 585
R231 B.n310 B.n309 585
R232 B.n493 B.n492 585
R233 B.n494 B.n493 585
R234 B.n491 B.n316 585
R235 B.n316 B.n315 585
R236 B.n490 B.n489 585
R237 B.n489 B.n488 585
R238 B.n318 B.n317 585
R239 B.n319 B.n318 585
R240 B.n481 B.n480 585
R241 B.n482 B.n481 585
R242 B.n322 B.n321 585
R243 B.n359 B.n357 585
R244 B.n360 B.n356 585
R245 B.n360 B.n323 585
R246 B.n363 B.n362 585
R247 B.n364 B.n355 585
R248 B.n366 B.n365 585
R249 B.n368 B.n354 585
R250 B.n371 B.n370 585
R251 B.n372 B.n353 585
R252 B.n374 B.n373 585
R253 B.n376 B.n352 585
R254 B.n379 B.n378 585
R255 B.n380 B.n351 585
R256 B.n382 B.n381 585
R257 B.n384 B.n350 585
R258 B.n387 B.n386 585
R259 B.n388 B.n349 585
R260 B.n390 B.n389 585
R261 B.n392 B.n348 585
R262 B.n395 B.n394 585
R263 B.n396 B.n347 585
R264 B.n398 B.n397 585
R265 B.n400 B.n346 585
R266 B.n403 B.n402 585
R267 B.n404 B.n345 585
R268 B.n409 B.n408 585
R269 B.n411 B.n344 585
R270 B.n414 B.n413 585
R271 B.n415 B.n343 585
R272 B.n417 B.n416 585
R273 B.n419 B.n342 585
R274 B.n422 B.n421 585
R275 B.n423 B.n341 585
R276 B.n425 B.n424 585
R277 B.n427 B.n340 585
R278 B.n430 B.n429 585
R279 B.n431 B.n336 585
R280 B.n433 B.n432 585
R281 B.n435 B.n335 585
R282 B.n438 B.n437 585
R283 B.n439 B.n334 585
R284 B.n441 B.n440 585
R285 B.n443 B.n333 585
R286 B.n446 B.n445 585
R287 B.n447 B.n332 585
R288 B.n449 B.n448 585
R289 B.n451 B.n331 585
R290 B.n454 B.n453 585
R291 B.n455 B.n330 585
R292 B.n457 B.n456 585
R293 B.n459 B.n329 585
R294 B.n462 B.n461 585
R295 B.n463 B.n328 585
R296 B.n465 B.n464 585
R297 B.n467 B.n327 585
R298 B.n470 B.n469 585
R299 B.n471 B.n326 585
R300 B.n473 B.n472 585
R301 B.n475 B.n325 585
R302 B.n478 B.n477 585
R303 B.n479 B.n324 585
R304 B.n484 B.n483 585
R305 B.n483 B.n482 585
R306 B.n485 B.n320 585
R307 B.n320 B.n319 585
R308 B.n487 B.n486 585
R309 B.n488 B.n487 585
R310 B.n314 B.n313 585
R311 B.n315 B.n314 585
R312 B.n496 B.n495 585
R313 B.n495 B.n494 585
R314 B.n497 B.n312 585
R315 B.n312 B.n310 585
R316 B.n499 B.n498 585
R317 B.n500 B.n499 585
R318 B.n306 B.n305 585
R319 B.n311 B.n306 585
R320 B.n508 B.n507 585
R321 B.n507 B.n506 585
R322 B.n509 B.n304 585
R323 B.n304 B.n303 585
R324 B.n511 B.n510 585
R325 B.n512 B.n511 585
R326 B.n298 B.n297 585
R327 B.n299 B.n298 585
R328 B.n520 B.n519 585
R329 B.n519 B.n518 585
R330 B.n521 B.n296 585
R331 B.n296 B.n295 585
R332 B.n523 B.n522 585
R333 B.n524 B.n523 585
R334 B.n290 B.n289 585
R335 B.n291 B.n290 585
R336 B.n532 B.n531 585
R337 B.n531 B.n530 585
R338 B.n533 B.n288 585
R339 B.n288 B.n287 585
R340 B.n535 B.n534 585
R341 B.n536 B.n535 585
R342 B.n282 B.n281 585
R343 B.n283 B.n282 585
R344 B.n544 B.n543 585
R345 B.n543 B.n542 585
R346 B.n545 B.n280 585
R347 B.n280 B.n279 585
R348 B.n547 B.n546 585
R349 B.n548 B.n547 585
R350 B.n274 B.n273 585
R351 B.n275 B.n274 585
R352 B.n556 B.n555 585
R353 B.n555 B.n554 585
R354 B.n557 B.n272 585
R355 B.n272 B.n271 585
R356 B.n559 B.n558 585
R357 B.n560 B.n559 585
R358 B.n266 B.n265 585
R359 B.n267 B.n266 585
R360 B.n569 B.n568 585
R361 B.n568 B.n567 585
R362 B.n570 B.n264 585
R363 B.n566 B.n264 585
R364 B.n572 B.n571 585
R365 B.n573 B.n572 585
R366 B.n259 B.n258 585
R367 B.n260 B.n259 585
R368 B.n581 B.n580 585
R369 B.n580 B.n579 585
R370 B.n582 B.n257 585
R371 B.n257 B.n256 585
R372 B.n584 B.n583 585
R373 B.n585 B.n584 585
R374 B.n251 B.n250 585
R375 B.n252 B.n251 585
R376 B.n593 B.n592 585
R377 B.n592 B.n591 585
R378 B.n594 B.n249 585
R379 B.n249 B.n248 585
R380 B.n596 B.n595 585
R381 B.n597 B.n596 585
R382 B.n243 B.n242 585
R383 B.n244 B.n243 585
R384 B.n606 B.n605 585
R385 B.n605 B.n604 585
R386 B.n607 B.n241 585
R387 B.n241 B.n240 585
R388 B.n609 B.n608 585
R389 B.n610 B.n609 585
R390 B.n3 B.n0 585
R391 B.n4 B.n3 585
R392 B.n761 B.n1 585
R393 B.n762 B.n761 585
R394 B.n760 B.n759 585
R395 B.n760 B.n8 585
R396 B.n758 B.n9 585
R397 B.n12 B.n9 585
R398 B.n757 B.n756 585
R399 B.n756 B.n755 585
R400 B.n11 B.n10 585
R401 B.n754 B.n11 585
R402 B.n752 B.n751 585
R403 B.n753 B.n752 585
R404 B.n750 B.n17 585
R405 B.n17 B.n16 585
R406 B.n749 B.n748 585
R407 B.n748 B.n747 585
R408 B.n19 B.n18 585
R409 B.n746 B.n19 585
R410 B.n744 B.n743 585
R411 B.n745 B.n744 585
R412 B.n742 B.n24 585
R413 B.n24 B.n23 585
R414 B.n741 B.n740 585
R415 B.n740 B.n739 585
R416 B.n26 B.n25 585
R417 B.n738 B.n26 585
R418 B.n736 B.n735 585
R419 B.n737 B.n736 585
R420 B.n734 B.n30 585
R421 B.n33 B.n30 585
R422 B.n733 B.n732 585
R423 B.n732 B.n731 585
R424 B.n32 B.n31 585
R425 B.n730 B.n32 585
R426 B.n728 B.n727 585
R427 B.n729 B.n728 585
R428 B.n726 B.n38 585
R429 B.n38 B.n37 585
R430 B.n725 B.n724 585
R431 B.n724 B.n723 585
R432 B.n40 B.n39 585
R433 B.n722 B.n40 585
R434 B.n720 B.n719 585
R435 B.n721 B.n720 585
R436 B.n718 B.n45 585
R437 B.n45 B.n44 585
R438 B.n717 B.n716 585
R439 B.n716 B.n715 585
R440 B.n47 B.n46 585
R441 B.n714 B.n47 585
R442 B.n712 B.n711 585
R443 B.n713 B.n712 585
R444 B.n710 B.n52 585
R445 B.n52 B.n51 585
R446 B.n709 B.n708 585
R447 B.n708 B.n707 585
R448 B.n54 B.n53 585
R449 B.n706 B.n54 585
R450 B.n704 B.n703 585
R451 B.n705 B.n704 585
R452 B.n702 B.n59 585
R453 B.n59 B.n58 585
R454 B.n701 B.n700 585
R455 B.n700 B.n699 585
R456 B.n61 B.n60 585
R457 B.n698 B.n61 585
R458 B.n696 B.n695 585
R459 B.n697 B.n696 585
R460 B.n694 B.n66 585
R461 B.n66 B.n65 585
R462 B.n693 B.n692 585
R463 B.n692 B.n691 585
R464 B.n68 B.n67 585
R465 B.n690 B.n68 585
R466 B.n688 B.n687 585
R467 B.n689 B.n688 585
R468 B.n686 B.n73 585
R469 B.n73 B.n72 585
R470 B.n685 B.n684 585
R471 B.n684 B.n683 585
R472 B.n75 B.n74 585
R473 B.n682 B.n75 585
R474 B.n680 B.n679 585
R475 B.n681 B.n680 585
R476 B.n678 B.n80 585
R477 B.n80 B.n79 585
R478 B.n677 B.n676 585
R479 B.n676 B.n675 585
R480 B.n765 B.n764 585
R481 B.n763 B.n2 585
R482 B.n676 B.n82 502.111
R483 B.n673 B.n83 502.111
R484 B.n481 B.n324 502.111
R485 B.n483 B.n322 502.111
R486 B.n117 B.t14 266.541
R487 B.n115 B.t6 266.541
R488 B.n337 B.t17 266.541
R489 B.n405 B.t10 266.541
R490 B.n674 B.n113 256.663
R491 B.n674 B.n112 256.663
R492 B.n674 B.n111 256.663
R493 B.n674 B.n110 256.663
R494 B.n674 B.n109 256.663
R495 B.n674 B.n108 256.663
R496 B.n674 B.n107 256.663
R497 B.n674 B.n106 256.663
R498 B.n674 B.n105 256.663
R499 B.n674 B.n104 256.663
R500 B.n674 B.n103 256.663
R501 B.n674 B.n102 256.663
R502 B.n674 B.n101 256.663
R503 B.n674 B.n100 256.663
R504 B.n674 B.n99 256.663
R505 B.n674 B.n98 256.663
R506 B.n674 B.n97 256.663
R507 B.n674 B.n96 256.663
R508 B.n674 B.n95 256.663
R509 B.n674 B.n94 256.663
R510 B.n674 B.n93 256.663
R511 B.n674 B.n92 256.663
R512 B.n674 B.n91 256.663
R513 B.n674 B.n90 256.663
R514 B.n674 B.n89 256.663
R515 B.n674 B.n88 256.663
R516 B.n674 B.n87 256.663
R517 B.n674 B.n86 256.663
R518 B.n674 B.n85 256.663
R519 B.n674 B.n84 256.663
R520 B.n358 B.n323 256.663
R521 B.n361 B.n323 256.663
R522 B.n367 B.n323 256.663
R523 B.n369 B.n323 256.663
R524 B.n375 B.n323 256.663
R525 B.n377 B.n323 256.663
R526 B.n383 B.n323 256.663
R527 B.n385 B.n323 256.663
R528 B.n391 B.n323 256.663
R529 B.n393 B.n323 256.663
R530 B.n399 B.n323 256.663
R531 B.n401 B.n323 256.663
R532 B.n410 B.n323 256.663
R533 B.n412 B.n323 256.663
R534 B.n418 B.n323 256.663
R535 B.n420 B.n323 256.663
R536 B.n426 B.n323 256.663
R537 B.n428 B.n323 256.663
R538 B.n434 B.n323 256.663
R539 B.n436 B.n323 256.663
R540 B.n442 B.n323 256.663
R541 B.n444 B.n323 256.663
R542 B.n450 B.n323 256.663
R543 B.n452 B.n323 256.663
R544 B.n458 B.n323 256.663
R545 B.n460 B.n323 256.663
R546 B.n466 B.n323 256.663
R547 B.n468 B.n323 256.663
R548 B.n474 B.n323 256.663
R549 B.n476 B.n323 256.663
R550 B.n767 B.n766 256.663
R551 B.n115 B.t8 249.816
R552 B.n337 B.t19 249.816
R553 B.n117 B.t15 249.816
R554 B.n405 B.t13 249.816
R555 B.n116 B.t9 190.083
R556 B.n338 B.t18 190.083
R557 B.n118 B.t16 190.083
R558 B.n406 B.t12 190.083
R559 B.n122 B.n121 163.367
R560 B.n126 B.n125 163.367
R561 B.n130 B.n129 163.367
R562 B.n134 B.n133 163.367
R563 B.n138 B.n137 163.367
R564 B.n142 B.n141 163.367
R565 B.n146 B.n145 163.367
R566 B.n150 B.n149 163.367
R567 B.n154 B.n153 163.367
R568 B.n158 B.n157 163.367
R569 B.n162 B.n161 163.367
R570 B.n166 B.n165 163.367
R571 B.n170 B.n169 163.367
R572 B.n174 B.n173 163.367
R573 B.n178 B.n177 163.367
R574 B.n182 B.n181 163.367
R575 B.n186 B.n185 163.367
R576 B.n191 B.n190 163.367
R577 B.n195 B.n194 163.367
R578 B.n199 B.n198 163.367
R579 B.n203 B.n202 163.367
R580 B.n207 B.n206 163.367
R581 B.n211 B.n210 163.367
R582 B.n215 B.n214 163.367
R583 B.n219 B.n218 163.367
R584 B.n223 B.n222 163.367
R585 B.n227 B.n226 163.367
R586 B.n231 B.n230 163.367
R587 B.n235 B.n234 163.367
R588 B.n673 B.n114 163.367
R589 B.n481 B.n318 163.367
R590 B.n489 B.n318 163.367
R591 B.n489 B.n316 163.367
R592 B.n493 B.n316 163.367
R593 B.n493 B.n309 163.367
R594 B.n501 B.n309 163.367
R595 B.n501 B.n307 163.367
R596 B.n505 B.n307 163.367
R597 B.n505 B.n302 163.367
R598 B.n513 B.n302 163.367
R599 B.n513 B.n300 163.367
R600 B.n517 B.n300 163.367
R601 B.n517 B.n294 163.367
R602 B.n525 B.n294 163.367
R603 B.n525 B.n292 163.367
R604 B.n529 B.n292 163.367
R605 B.n529 B.n286 163.367
R606 B.n537 B.n286 163.367
R607 B.n537 B.n284 163.367
R608 B.n541 B.n284 163.367
R609 B.n541 B.n278 163.367
R610 B.n549 B.n278 163.367
R611 B.n549 B.n276 163.367
R612 B.n553 B.n276 163.367
R613 B.n553 B.n270 163.367
R614 B.n561 B.n270 163.367
R615 B.n561 B.n268 163.367
R616 B.n565 B.n268 163.367
R617 B.n565 B.n263 163.367
R618 B.n574 B.n263 163.367
R619 B.n574 B.n261 163.367
R620 B.n578 B.n261 163.367
R621 B.n578 B.n255 163.367
R622 B.n586 B.n255 163.367
R623 B.n586 B.n253 163.367
R624 B.n590 B.n253 163.367
R625 B.n590 B.n247 163.367
R626 B.n598 B.n247 163.367
R627 B.n598 B.n245 163.367
R628 B.n603 B.n245 163.367
R629 B.n603 B.n239 163.367
R630 B.n611 B.n239 163.367
R631 B.n612 B.n611 163.367
R632 B.n612 B.n5 163.367
R633 B.n6 B.n5 163.367
R634 B.n7 B.n6 163.367
R635 B.n618 B.n7 163.367
R636 B.n619 B.n618 163.367
R637 B.n619 B.n13 163.367
R638 B.n14 B.n13 163.367
R639 B.n15 B.n14 163.367
R640 B.n624 B.n15 163.367
R641 B.n624 B.n20 163.367
R642 B.n21 B.n20 163.367
R643 B.n22 B.n21 163.367
R644 B.n629 B.n22 163.367
R645 B.n629 B.n27 163.367
R646 B.n28 B.n27 163.367
R647 B.n29 B.n28 163.367
R648 B.n634 B.n29 163.367
R649 B.n634 B.n34 163.367
R650 B.n35 B.n34 163.367
R651 B.n36 B.n35 163.367
R652 B.n639 B.n36 163.367
R653 B.n639 B.n41 163.367
R654 B.n42 B.n41 163.367
R655 B.n43 B.n42 163.367
R656 B.n644 B.n43 163.367
R657 B.n644 B.n48 163.367
R658 B.n49 B.n48 163.367
R659 B.n50 B.n49 163.367
R660 B.n649 B.n50 163.367
R661 B.n649 B.n55 163.367
R662 B.n56 B.n55 163.367
R663 B.n57 B.n56 163.367
R664 B.n654 B.n57 163.367
R665 B.n654 B.n62 163.367
R666 B.n63 B.n62 163.367
R667 B.n64 B.n63 163.367
R668 B.n659 B.n64 163.367
R669 B.n659 B.n69 163.367
R670 B.n70 B.n69 163.367
R671 B.n71 B.n70 163.367
R672 B.n664 B.n71 163.367
R673 B.n664 B.n76 163.367
R674 B.n77 B.n76 163.367
R675 B.n78 B.n77 163.367
R676 B.n669 B.n78 163.367
R677 B.n669 B.n83 163.367
R678 B.n360 B.n359 163.367
R679 B.n362 B.n360 163.367
R680 B.n366 B.n355 163.367
R681 B.n370 B.n368 163.367
R682 B.n374 B.n353 163.367
R683 B.n378 B.n376 163.367
R684 B.n382 B.n351 163.367
R685 B.n386 B.n384 163.367
R686 B.n390 B.n349 163.367
R687 B.n394 B.n392 163.367
R688 B.n398 B.n347 163.367
R689 B.n402 B.n400 163.367
R690 B.n409 B.n345 163.367
R691 B.n413 B.n411 163.367
R692 B.n417 B.n343 163.367
R693 B.n421 B.n419 163.367
R694 B.n425 B.n341 163.367
R695 B.n429 B.n427 163.367
R696 B.n433 B.n336 163.367
R697 B.n437 B.n435 163.367
R698 B.n441 B.n334 163.367
R699 B.n445 B.n443 163.367
R700 B.n449 B.n332 163.367
R701 B.n453 B.n451 163.367
R702 B.n457 B.n330 163.367
R703 B.n461 B.n459 163.367
R704 B.n465 B.n328 163.367
R705 B.n469 B.n467 163.367
R706 B.n473 B.n326 163.367
R707 B.n477 B.n475 163.367
R708 B.n483 B.n320 163.367
R709 B.n487 B.n320 163.367
R710 B.n487 B.n314 163.367
R711 B.n495 B.n314 163.367
R712 B.n495 B.n312 163.367
R713 B.n499 B.n312 163.367
R714 B.n499 B.n306 163.367
R715 B.n507 B.n306 163.367
R716 B.n507 B.n304 163.367
R717 B.n511 B.n304 163.367
R718 B.n511 B.n298 163.367
R719 B.n519 B.n298 163.367
R720 B.n519 B.n296 163.367
R721 B.n523 B.n296 163.367
R722 B.n523 B.n290 163.367
R723 B.n531 B.n290 163.367
R724 B.n531 B.n288 163.367
R725 B.n535 B.n288 163.367
R726 B.n535 B.n282 163.367
R727 B.n543 B.n282 163.367
R728 B.n543 B.n280 163.367
R729 B.n547 B.n280 163.367
R730 B.n547 B.n274 163.367
R731 B.n555 B.n274 163.367
R732 B.n555 B.n272 163.367
R733 B.n559 B.n272 163.367
R734 B.n559 B.n266 163.367
R735 B.n568 B.n266 163.367
R736 B.n568 B.n264 163.367
R737 B.n572 B.n264 163.367
R738 B.n572 B.n259 163.367
R739 B.n580 B.n259 163.367
R740 B.n580 B.n257 163.367
R741 B.n584 B.n257 163.367
R742 B.n584 B.n251 163.367
R743 B.n592 B.n251 163.367
R744 B.n592 B.n249 163.367
R745 B.n596 B.n249 163.367
R746 B.n596 B.n243 163.367
R747 B.n605 B.n243 163.367
R748 B.n605 B.n241 163.367
R749 B.n609 B.n241 163.367
R750 B.n609 B.n3 163.367
R751 B.n765 B.n3 163.367
R752 B.n761 B.n2 163.367
R753 B.n761 B.n760 163.367
R754 B.n760 B.n9 163.367
R755 B.n756 B.n9 163.367
R756 B.n756 B.n11 163.367
R757 B.n752 B.n11 163.367
R758 B.n752 B.n17 163.367
R759 B.n748 B.n17 163.367
R760 B.n748 B.n19 163.367
R761 B.n744 B.n19 163.367
R762 B.n744 B.n24 163.367
R763 B.n740 B.n24 163.367
R764 B.n740 B.n26 163.367
R765 B.n736 B.n26 163.367
R766 B.n736 B.n30 163.367
R767 B.n732 B.n30 163.367
R768 B.n732 B.n32 163.367
R769 B.n728 B.n32 163.367
R770 B.n728 B.n38 163.367
R771 B.n724 B.n38 163.367
R772 B.n724 B.n40 163.367
R773 B.n720 B.n40 163.367
R774 B.n720 B.n45 163.367
R775 B.n716 B.n45 163.367
R776 B.n716 B.n47 163.367
R777 B.n712 B.n47 163.367
R778 B.n712 B.n52 163.367
R779 B.n708 B.n52 163.367
R780 B.n708 B.n54 163.367
R781 B.n704 B.n54 163.367
R782 B.n704 B.n59 163.367
R783 B.n700 B.n59 163.367
R784 B.n700 B.n61 163.367
R785 B.n696 B.n61 163.367
R786 B.n696 B.n66 163.367
R787 B.n692 B.n66 163.367
R788 B.n692 B.n68 163.367
R789 B.n688 B.n68 163.367
R790 B.n688 B.n73 163.367
R791 B.n684 B.n73 163.367
R792 B.n684 B.n75 163.367
R793 B.n680 B.n75 163.367
R794 B.n680 B.n80 163.367
R795 B.n676 B.n80 163.367
R796 B.n482 B.n323 104.236
R797 B.n675 B.n674 104.236
R798 B.n84 B.n82 71.676
R799 B.n122 B.n85 71.676
R800 B.n126 B.n86 71.676
R801 B.n130 B.n87 71.676
R802 B.n134 B.n88 71.676
R803 B.n138 B.n89 71.676
R804 B.n142 B.n90 71.676
R805 B.n146 B.n91 71.676
R806 B.n150 B.n92 71.676
R807 B.n154 B.n93 71.676
R808 B.n158 B.n94 71.676
R809 B.n162 B.n95 71.676
R810 B.n166 B.n96 71.676
R811 B.n170 B.n97 71.676
R812 B.n174 B.n98 71.676
R813 B.n178 B.n99 71.676
R814 B.n182 B.n100 71.676
R815 B.n186 B.n101 71.676
R816 B.n191 B.n102 71.676
R817 B.n195 B.n103 71.676
R818 B.n199 B.n104 71.676
R819 B.n203 B.n105 71.676
R820 B.n207 B.n106 71.676
R821 B.n211 B.n107 71.676
R822 B.n215 B.n108 71.676
R823 B.n219 B.n109 71.676
R824 B.n223 B.n110 71.676
R825 B.n227 B.n111 71.676
R826 B.n231 B.n112 71.676
R827 B.n235 B.n113 71.676
R828 B.n114 B.n113 71.676
R829 B.n234 B.n112 71.676
R830 B.n230 B.n111 71.676
R831 B.n226 B.n110 71.676
R832 B.n222 B.n109 71.676
R833 B.n218 B.n108 71.676
R834 B.n214 B.n107 71.676
R835 B.n210 B.n106 71.676
R836 B.n206 B.n105 71.676
R837 B.n202 B.n104 71.676
R838 B.n198 B.n103 71.676
R839 B.n194 B.n102 71.676
R840 B.n190 B.n101 71.676
R841 B.n185 B.n100 71.676
R842 B.n181 B.n99 71.676
R843 B.n177 B.n98 71.676
R844 B.n173 B.n97 71.676
R845 B.n169 B.n96 71.676
R846 B.n165 B.n95 71.676
R847 B.n161 B.n94 71.676
R848 B.n157 B.n93 71.676
R849 B.n153 B.n92 71.676
R850 B.n149 B.n91 71.676
R851 B.n145 B.n90 71.676
R852 B.n141 B.n89 71.676
R853 B.n137 B.n88 71.676
R854 B.n133 B.n87 71.676
R855 B.n129 B.n86 71.676
R856 B.n125 B.n85 71.676
R857 B.n121 B.n84 71.676
R858 B.n358 B.n322 71.676
R859 B.n362 B.n361 71.676
R860 B.n367 B.n366 71.676
R861 B.n370 B.n369 71.676
R862 B.n375 B.n374 71.676
R863 B.n378 B.n377 71.676
R864 B.n383 B.n382 71.676
R865 B.n386 B.n385 71.676
R866 B.n391 B.n390 71.676
R867 B.n394 B.n393 71.676
R868 B.n399 B.n398 71.676
R869 B.n402 B.n401 71.676
R870 B.n410 B.n409 71.676
R871 B.n413 B.n412 71.676
R872 B.n418 B.n417 71.676
R873 B.n421 B.n420 71.676
R874 B.n426 B.n425 71.676
R875 B.n429 B.n428 71.676
R876 B.n434 B.n433 71.676
R877 B.n437 B.n436 71.676
R878 B.n442 B.n441 71.676
R879 B.n445 B.n444 71.676
R880 B.n450 B.n449 71.676
R881 B.n453 B.n452 71.676
R882 B.n458 B.n457 71.676
R883 B.n461 B.n460 71.676
R884 B.n466 B.n465 71.676
R885 B.n469 B.n468 71.676
R886 B.n474 B.n473 71.676
R887 B.n477 B.n476 71.676
R888 B.n359 B.n358 71.676
R889 B.n361 B.n355 71.676
R890 B.n368 B.n367 71.676
R891 B.n369 B.n353 71.676
R892 B.n376 B.n375 71.676
R893 B.n377 B.n351 71.676
R894 B.n384 B.n383 71.676
R895 B.n385 B.n349 71.676
R896 B.n392 B.n391 71.676
R897 B.n393 B.n347 71.676
R898 B.n400 B.n399 71.676
R899 B.n401 B.n345 71.676
R900 B.n411 B.n410 71.676
R901 B.n412 B.n343 71.676
R902 B.n419 B.n418 71.676
R903 B.n420 B.n341 71.676
R904 B.n427 B.n426 71.676
R905 B.n428 B.n336 71.676
R906 B.n435 B.n434 71.676
R907 B.n436 B.n334 71.676
R908 B.n443 B.n442 71.676
R909 B.n444 B.n332 71.676
R910 B.n451 B.n450 71.676
R911 B.n452 B.n330 71.676
R912 B.n459 B.n458 71.676
R913 B.n460 B.n328 71.676
R914 B.n467 B.n466 71.676
R915 B.n468 B.n326 71.676
R916 B.n475 B.n474 71.676
R917 B.n476 B.n324 71.676
R918 B.n766 B.n765 71.676
R919 B.n766 B.n2 71.676
R920 B.n482 B.n319 62.7259
R921 B.n488 B.n319 62.7259
R922 B.n488 B.n315 62.7259
R923 B.n494 B.n315 62.7259
R924 B.n494 B.n310 62.7259
R925 B.n500 B.n310 62.7259
R926 B.n500 B.n311 62.7259
R927 B.n506 B.n303 62.7259
R928 B.n512 B.n303 62.7259
R929 B.n512 B.n299 62.7259
R930 B.n518 B.n299 62.7259
R931 B.n518 B.n295 62.7259
R932 B.n524 B.n295 62.7259
R933 B.n524 B.n291 62.7259
R934 B.n530 B.n291 62.7259
R935 B.n530 B.n287 62.7259
R936 B.n536 B.n287 62.7259
R937 B.n536 B.n283 62.7259
R938 B.n542 B.n283 62.7259
R939 B.n548 B.n279 62.7259
R940 B.n548 B.n275 62.7259
R941 B.n554 B.n275 62.7259
R942 B.n554 B.n271 62.7259
R943 B.n560 B.n271 62.7259
R944 B.n560 B.n267 62.7259
R945 B.n567 B.n267 62.7259
R946 B.n567 B.n566 62.7259
R947 B.n573 B.n260 62.7259
R948 B.n579 B.n260 62.7259
R949 B.n579 B.n256 62.7259
R950 B.n585 B.n256 62.7259
R951 B.n585 B.n252 62.7259
R952 B.n591 B.n252 62.7259
R953 B.n591 B.n248 62.7259
R954 B.n597 B.n248 62.7259
R955 B.n604 B.n244 62.7259
R956 B.n604 B.n240 62.7259
R957 B.n610 B.n240 62.7259
R958 B.n610 B.n4 62.7259
R959 B.n764 B.n4 62.7259
R960 B.n764 B.n763 62.7259
R961 B.n763 B.n762 62.7259
R962 B.n762 B.n8 62.7259
R963 B.n12 B.n8 62.7259
R964 B.n755 B.n12 62.7259
R965 B.n755 B.n754 62.7259
R966 B.n753 B.n16 62.7259
R967 B.n747 B.n16 62.7259
R968 B.n747 B.n746 62.7259
R969 B.n746 B.n745 62.7259
R970 B.n745 B.n23 62.7259
R971 B.n739 B.n23 62.7259
R972 B.n739 B.n738 62.7259
R973 B.n738 B.n737 62.7259
R974 B.n731 B.n33 62.7259
R975 B.n731 B.n730 62.7259
R976 B.n730 B.n729 62.7259
R977 B.n729 B.n37 62.7259
R978 B.n723 B.n37 62.7259
R979 B.n723 B.n722 62.7259
R980 B.n722 B.n721 62.7259
R981 B.n721 B.n44 62.7259
R982 B.n715 B.n714 62.7259
R983 B.n714 B.n713 62.7259
R984 B.n713 B.n51 62.7259
R985 B.n707 B.n51 62.7259
R986 B.n707 B.n706 62.7259
R987 B.n706 B.n705 62.7259
R988 B.n705 B.n58 62.7259
R989 B.n699 B.n58 62.7259
R990 B.n699 B.n698 62.7259
R991 B.n698 B.n697 62.7259
R992 B.n697 B.n65 62.7259
R993 B.n691 B.n65 62.7259
R994 B.n690 B.n689 62.7259
R995 B.n689 B.n72 62.7259
R996 B.n683 B.n72 62.7259
R997 B.n683 B.n682 62.7259
R998 B.n682 B.n681 62.7259
R999 B.n681 B.n79 62.7259
R1000 B.n675 B.n79 62.7259
R1001 B.n311 B.t11 61.8034
R1002 B.t7 B.n690 61.8034
R1003 B.n118 B.n117 59.7338
R1004 B.n116 B.n115 59.7338
R1005 B.n338 B.n337 59.7338
R1006 B.n406 B.n405 59.7338
R1007 B.n119 B.n118 59.5399
R1008 B.n188 B.n116 59.5399
R1009 B.n339 B.n338 59.5399
R1010 B.n407 B.n406 59.5399
R1011 B.t5 B.n279 47.0445
R1012 B.t0 B.n44 47.0445
R1013 B.n573 B.t3 43.3548
R1014 B.n737 B.t2 43.3548
R1015 B.t1 B.n244 39.6651
R1016 B.n754 B.t4 39.6651
R1017 B.n484 B.n321 32.6249
R1018 B.n480 B.n479 32.6249
R1019 B.n672 B.n671 32.6249
R1020 B.n677 B.n81 32.6249
R1021 B.n597 B.t1 23.0613
R1022 B.t4 B.n753 23.0613
R1023 B.n566 B.t3 19.3716
R1024 B.n33 B.t2 19.3716
R1025 B B.n767 18.0485
R1026 B.n542 B.t5 15.6818
R1027 B.n715 B.t0 15.6818
R1028 B.n485 B.n484 10.6151
R1029 B.n486 B.n485 10.6151
R1030 B.n486 B.n313 10.6151
R1031 B.n496 B.n313 10.6151
R1032 B.n497 B.n496 10.6151
R1033 B.n498 B.n497 10.6151
R1034 B.n498 B.n305 10.6151
R1035 B.n508 B.n305 10.6151
R1036 B.n509 B.n508 10.6151
R1037 B.n510 B.n509 10.6151
R1038 B.n510 B.n297 10.6151
R1039 B.n520 B.n297 10.6151
R1040 B.n521 B.n520 10.6151
R1041 B.n522 B.n521 10.6151
R1042 B.n522 B.n289 10.6151
R1043 B.n532 B.n289 10.6151
R1044 B.n533 B.n532 10.6151
R1045 B.n534 B.n533 10.6151
R1046 B.n534 B.n281 10.6151
R1047 B.n544 B.n281 10.6151
R1048 B.n545 B.n544 10.6151
R1049 B.n546 B.n545 10.6151
R1050 B.n546 B.n273 10.6151
R1051 B.n556 B.n273 10.6151
R1052 B.n557 B.n556 10.6151
R1053 B.n558 B.n557 10.6151
R1054 B.n558 B.n265 10.6151
R1055 B.n569 B.n265 10.6151
R1056 B.n570 B.n569 10.6151
R1057 B.n571 B.n570 10.6151
R1058 B.n571 B.n258 10.6151
R1059 B.n581 B.n258 10.6151
R1060 B.n582 B.n581 10.6151
R1061 B.n583 B.n582 10.6151
R1062 B.n583 B.n250 10.6151
R1063 B.n593 B.n250 10.6151
R1064 B.n594 B.n593 10.6151
R1065 B.n595 B.n594 10.6151
R1066 B.n595 B.n242 10.6151
R1067 B.n606 B.n242 10.6151
R1068 B.n607 B.n606 10.6151
R1069 B.n608 B.n607 10.6151
R1070 B.n608 B.n0 10.6151
R1071 B.n357 B.n321 10.6151
R1072 B.n357 B.n356 10.6151
R1073 B.n363 B.n356 10.6151
R1074 B.n364 B.n363 10.6151
R1075 B.n365 B.n364 10.6151
R1076 B.n365 B.n354 10.6151
R1077 B.n371 B.n354 10.6151
R1078 B.n372 B.n371 10.6151
R1079 B.n373 B.n372 10.6151
R1080 B.n373 B.n352 10.6151
R1081 B.n379 B.n352 10.6151
R1082 B.n380 B.n379 10.6151
R1083 B.n381 B.n380 10.6151
R1084 B.n381 B.n350 10.6151
R1085 B.n387 B.n350 10.6151
R1086 B.n388 B.n387 10.6151
R1087 B.n389 B.n388 10.6151
R1088 B.n389 B.n348 10.6151
R1089 B.n395 B.n348 10.6151
R1090 B.n396 B.n395 10.6151
R1091 B.n397 B.n396 10.6151
R1092 B.n397 B.n346 10.6151
R1093 B.n403 B.n346 10.6151
R1094 B.n404 B.n403 10.6151
R1095 B.n408 B.n404 10.6151
R1096 B.n414 B.n344 10.6151
R1097 B.n415 B.n414 10.6151
R1098 B.n416 B.n415 10.6151
R1099 B.n416 B.n342 10.6151
R1100 B.n422 B.n342 10.6151
R1101 B.n423 B.n422 10.6151
R1102 B.n424 B.n423 10.6151
R1103 B.n424 B.n340 10.6151
R1104 B.n431 B.n430 10.6151
R1105 B.n432 B.n431 10.6151
R1106 B.n432 B.n335 10.6151
R1107 B.n438 B.n335 10.6151
R1108 B.n439 B.n438 10.6151
R1109 B.n440 B.n439 10.6151
R1110 B.n440 B.n333 10.6151
R1111 B.n446 B.n333 10.6151
R1112 B.n447 B.n446 10.6151
R1113 B.n448 B.n447 10.6151
R1114 B.n448 B.n331 10.6151
R1115 B.n454 B.n331 10.6151
R1116 B.n455 B.n454 10.6151
R1117 B.n456 B.n455 10.6151
R1118 B.n456 B.n329 10.6151
R1119 B.n462 B.n329 10.6151
R1120 B.n463 B.n462 10.6151
R1121 B.n464 B.n463 10.6151
R1122 B.n464 B.n327 10.6151
R1123 B.n470 B.n327 10.6151
R1124 B.n471 B.n470 10.6151
R1125 B.n472 B.n471 10.6151
R1126 B.n472 B.n325 10.6151
R1127 B.n478 B.n325 10.6151
R1128 B.n479 B.n478 10.6151
R1129 B.n480 B.n317 10.6151
R1130 B.n490 B.n317 10.6151
R1131 B.n491 B.n490 10.6151
R1132 B.n492 B.n491 10.6151
R1133 B.n492 B.n308 10.6151
R1134 B.n502 B.n308 10.6151
R1135 B.n503 B.n502 10.6151
R1136 B.n504 B.n503 10.6151
R1137 B.n504 B.n301 10.6151
R1138 B.n514 B.n301 10.6151
R1139 B.n515 B.n514 10.6151
R1140 B.n516 B.n515 10.6151
R1141 B.n516 B.n293 10.6151
R1142 B.n526 B.n293 10.6151
R1143 B.n527 B.n526 10.6151
R1144 B.n528 B.n527 10.6151
R1145 B.n528 B.n285 10.6151
R1146 B.n538 B.n285 10.6151
R1147 B.n539 B.n538 10.6151
R1148 B.n540 B.n539 10.6151
R1149 B.n540 B.n277 10.6151
R1150 B.n550 B.n277 10.6151
R1151 B.n551 B.n550 10.6151
R1152 B.n552 B.n551 10.6151
R1153 B.n552 B.n269 10.6151
R1154 B.n562 B.n269 10.6151
R1155 B.n563 B.n562 10.6151
R1156 B.n564 B.n563 10.6151
R1157 B.n564 B.n262 10.6151
R1158 B.n575 B.n262 10.6151
R1159 B.n576 B.n575 10.6151
R1160 B.n577 B.n576 10.6151
R1161 B.n577 B.n254 10.6151
R1162 B.n587 B.n254 10.6151
R1163 B.n588 B.n587 10.6151
R1164 B.n589 B.n588 10.6151
R1165 B.n589 B.n246 10.6151
R1166 B.n599 B.n246 10.6151
R1167 B.n600 B.n599 10.6151
R1168 B.n602 B.n600 10.6151
R1169 B.n602 B.n601 10.6151
R1170 B.n601 B.n238 10.6151
R1171 B.n613 B.n238 10.6151
R1172 B.n614 B.n613 10.6151
R1173 B.n615 B.n614 10.6151
R1174 B.n616 B.n615 10.6151
R1175 B.n617 B.n616 10.6151
R1176 B.n620 B.n617 10.6151
R1177 B.n621 B.n620 10.6151
R1178 B.n622 B.n621 10.6151
R1179 B.n623 B.n622 10.6151
R1180 B.n625 B.n623 10.6151
R1181 B.n626 B.n625 10.6151
R1182 B.n627 B.n626 10.6151
R1183 B.n628 B.n627 10.6151
R1184 B.n630 B.n628 10.6151
R1185 B.n631 B.n630 10.6151
R1186 B.n632 B.n631 10.6151
R1187 B.n633 B.n632 10.6151
R1188 B.n635 B.n633 10.6151
R1189 B.n636 B.n635 10.6151
R1190 B.n637 B.n636 10.6151
R1191 B.n638 B.n637 10.6151
R1192 B.n640 B.n638 10.6151
R1193 B.n641 B.n640 10.6151
R1194 B.n642 B.n641 10.6151
R1195 B.n643 B.n642 10.6151
R1196 B.n645 B.n643 10.6151
R1197 B.n646 B.n645 10.6151
R1198 B.n647 B.n646 10.6151
R1199 B.n648 B.n647 10.6151
R1200 B.n650 B.n648 10.6151
R1201 B.n651 B.n650 10.6151
R1202 B.n652 B.n651 10.6151
R1203 B.n653 B.n652 10.6151
R1204 B.n655 B.n653 10.6151
R1205 B.n656 B.n655 10.6151
R1206 B.n657 B.n656 10.6151
R1207 B.n658 B.n657 10.6151
R1208 B.n660 B.n658 10.6151
R1209 B.n661 B.n660 10.6151
R1210 B.n662 B.n661 10.6151
R1211 B.n663 B.n662 10.6151
R1212 B.n665 B.n663 10.6151
R1213 B.n666 B.n665 10.6151
R1214 B.n667 B.n666 10.6151
R1215 B.n668 B.n667 10.6151
R1216 B.n670 B.n668 10.6151
R1217 B.n671 B.n670 10.6151
R1218 B.n759 B.n1 10.6151
R1219 B.n759 B.n758 10.6151
R1220 B.n758 B.n757 10.6151
R1221 B.n757 B.n10 10.6151
R1222 B.n751 B.n10 10.6151
R1223 B.n751 B.n750 10.6151
R1224 B.n750 B.n749 10.6151
R1225 B.n749 B.n18 10.6151
R1226 B.n743 B.n18 10.6151
R1227 B.n743 B.n742 10.6151
R1228 B.n742 B.n741 10.6151
R1229 B.n741 B.n25 10.6151
R1230 B.n735 B.n25 10.6151
R1231 B.n735 B.n734 10.6151
R1232 B.n734 B.n733 10.6151
R1233 B.n733 B.n31 10.6151
R1234 B.n727 B.n31 10.6151
R1235 B.n727 B.n726 10.6151
R1236 B.n726 B.n725 10.6151
R1237 B.n725 B.n39 10.6151
R1238 B.n719 B.n39 10.6151
R1239 B.n719 B.n718 10.6151
R1240 B.n718 B.n717 10.6151
R1241 B.n717 B.n46 10.6151
R1242 B.n711 B.n46 10.6151
R1243 B.n711 B.n710 10.6151
R1244 B.n710 B.n709 10.6151
R1245 B.n709 B.n53 10.6151
R1246 B.n703 B.n53 10.6151
R1247 B.n703 B.n702 10.6151
R1248 B.n702 B.n701 10.6151
R1249 B.n701 B.n60 10.6151
R1250 B.n695 B.n60 10.6151
R1251 B.n695 B.n694 10.6151
R1252 B.n694 B.n693 10.6151
R1253 B.n693 B.n67 10.6151
R1254 B.n687 B.n67 10.6151
R1255 B.n687 B.n686 10.6151
R1256 B.n686 B.n685 10.6151
R1257 B.n685 B.n74 10.6151
R1258 B.n679 B.n74 10.6151
R1259 B.n679 B.n678 10.6151
R1260 B.n678 B.n677 10.6151
R1261 B.n120 B.n81 10.6151
R1262 B.n123 B.n120 10.6151
R1263 B.n124 B.n123 10.6151
R1264 B.n127 B.n124 10.6151
R1265 B.n128 B.n127 10.6151
R1266 B.n131 B.n128 10.6151
R1267 B.n132 B.n131 10.6151
R1268 B.n135 B.n132 10.6151
R1269 B.n136 B.n135 10.6151
R1270 B.n139 B.n136 10.6151
R1271 B.n140 B.n139 10.6151
R1272 B.n143 B.n140 10.6151
R1273 B.n144 B.n143 10.6151
R1274 B.n147 B.n144 10.6151
R1275 B.n148 B.n147 10.6151
R1276 B.n151 B.n148 10.6151
R1277 B.n152 B.n151 10.6151
R1278 B.n155 B.n152 10.6151
R1279 B.n156 B.n155 10.6151
R1280 B.n159 B.n156 10.6151
R1281 B.n160 B.n159 10.6151
R1282 B.n163 B.n160 10.6151
R1283 B.n164 B.n163 10.6151
R1284 B.n167 B.n164 10.6151
R1285 B.n168 B.n167 10.6151
R1286 B.n172 B.n171 10.6151
R1287 B.n175 B.n172 10.6151
R1288 B.n176 B.n175 10.6151
R1289 B.n179 B.n176 10.6151
R1290 B.n180 B.n179 10.6151
R1291 B.n183 B.n180 10.6151
R1292 B.n184 B.n183 10.6151
R1293 B.n187 B.n184 10.6151
R1294 B.n192 B.n189 10.6151
R1295 B.n193 B.n192 10.6151
R1296 B.n196 B.n193 10.6151
R1297 B.n197 B.n196 10.6151
R1298 B.n200 B.n197 10.6151
R1299 B.n201 B.n200 10.6151
R1300 B.n204 B.n201 10.6151
R1301 B.n205 B.n204 10.6151
R1302 B.n208 B.n205 10.6151
R1303 B.n209 B.n208 10.6151
R1304 B.n212 B.n209 10.6151
R1305 B.n213 B.n212 10.6151
R1306 B.n216 B.n213 10.6151
R1307 B.n217 B.n216 10.6151
R1308 B.n220 B.n217 10.6151
R1309 B.n221 B.n220 10.6151
R1310 B.n224 B.n221 10.6151
R1311 B.n225 B.n224 10.6151
R1312 B.n228 B.n225 10.6151
R1313 B.n229 B.n228 10.6151
R1314 B.n232 B.n229 10.6151
R1315 B.n233 B.n232 10.6151
R1316 B.n236 B.n233 10.6151
R1317 B.n237 B.n236 10.6151
R1318 B.n672 B.n237 10.6151
R1319 B.n767 B.n0 8.11757
R1320 B.n767 B.n1 8.11757
R1321 B.n407 B.n344 6.5566
R1322 B.n340 B.n339 6.5566
R1323 B.n171 B.n119 6.5566
R1324 B.n188 B.n187 6.5566
R1325 B.n408 B.n407 4.05904
R1326 B.n430 B.n339 4.05904
R1327 B.n168 B.n119 4.05904
R1328 B.n189 B.n188 4.05904
R1329 B.n506 B.t11 0.922932
R1330 B.n691 B.t7 0.922932
R1331 VP.n13 VP.n12 161.3
R1332 VP.n14 VP.n9 161.3
R1333 VP.n16 VP.n15 161.3
R1334 VP.n17 VP.n8 161.3
R1335 VP.n19 VP.n18 161.3
R1336 VP.n20 VP.n7 161.3
R1337 VP.n43 VP.n0 161.3
R1338 VP.n42 VP.n41 161.3
R1339 VP.n40 VP.n1 161.3
R1340 VP.n39 VP.n38 161.3
R1341 VP.n37 VP.n2 161.3
R1342 VP.n36 VP.n35 161.3
R1343 VP.n34 VP.n3 161.3
R1344 VP.n33 VP.n32 161.3
R1345 VP.n31 VP.n4 161.3
R1346 VP.n30 VP.n29 161.3
R1347 VP.n28 VP.n5 161.3
R1348 VP.n27 VP.n26 161.3
R1349 VP.n25 VP.n6 161.3
R1350 VP.n24 VP.n23 106.841
R1351 VP.n45 VP.n44 106.841
R1352 VP.n22 VP.n21 106.841
R1353 VP.n11 VP.t3 91.9343
R1354 VP.n3 VP.t1 58.2787
R1355 VP.n24 VP.t2 58.2787
R1356 VP.n44 VP.t0 58.2787
R1357 VP.n10 VP.t5 58.2787
R1358 VP.n21 VP.t4 58.2787
R1359 VP.n11 VP.n10 48.924
R1360 VP.n23 VP.n22 45.1738
R1361 VP.n30 VP.n5 44.3785
R1362 VP.n38 VP.n1 44.3785
R1363 VP.n15 VP.n8 44.3785
R1364 VP.n31 VP.n30 36.6083
R1365 VP.n38 VP.n37 36.6083
R1366 VP.n15 VP.n14 36.6083
R1367 VP.n26 VP.n25 24.4675
R1368 VP.n26 VP.n5 24.4675
R1369 VP.n32 VP.n31 24.4675
R1370 VP.n32 VP.n3 24.4675
R1371 VP.n36 VP.n3 24.4675
R1372 VP.n37 VP.n36 24.4675
R1373 VP.n42 VP.n1 24.4675
R1374 VP.n43 VP.n42 24.4675
R1375 VP.n19 VP.n8 24.4675
R1376 VP.n20 VP.n19 24.4675
R1377 VP.n13 VP.n10 24.4675
R1378 VP.n14 VP.n13 24.4675
R1379 VP.n12 VP.n11 5.02272
R1380 VP.n25 VP.n24 3.91522
R1381 VP.n44 VP.n43 3.91522
R1382 VP.n21 VP.n20 3.91522
R1383 VP.n22 VP.n7 0.278367
R1384 VP.n23 VP.n6 0.278367
R1385 VP.n45 VP.n0 0.278367
R1386 VP.n12 VP.n9 0.189894
R1387 VP.n16 VP.n9 0.189894
R1388 VP.n17 VP.n16 0.189894
R1389 VP.n18 VP.n17 0.189894
R1390 VP.n18 VP.n7 0.189894
R1391 VP.n27 VP.n6 0.189894
R1392 VP.n28 VP.n27 0.189894
R1393 VP.n29 VP.n28 0.189894
R1394 VP.n29 VP.n4 0.189894
R1395 VP.n33 VP.n4 0.189894
R1396 VP.n34 VP.n33 0.189894
R1397 VP.n35 VP.n34 0.189894
R1398 VP.n35 VP.n2 0.189894
R1399 VP.n39 VP.n2 0.189894
R1400 VP.n40 VP.n39 0.189894
R1401 VP.n41 VP.n40 0.189894
R1402 VP.n41 VP.n0 0.189894
R1403 VP VP.n45 0.153454
R1404 VTAIL.n146 VTAIL.n116 289.615
R1405 VTAIL.n32 VTAIL.n2 289.615
R1406 VTAIL.n110 VTAIL.n80 289.615
R1407 VTAIL.n72 VTAIL.n42 289.615
R1408 VTAIL.n129 VTAIL.n128 185
R1409 VTAIL.n131 VTAIL.n130 185
R1410 VTAIL.n124 VTAIL.n123 185
R1411 VTAIL.n137 VTAIL.n136 185
R1412 VTAIL.n139 VTAIL.n138 185
R1413 VTAIL.n120 VTAIL.n119 185
R1414 VTAIL.n145 VTAIL.n144 185
R1415 VTAIL.n147 VTAIL.n146 185
R1416 VTAIL.n15 VTAIL.n14 185
R1417 VTAIL.n17 VTAIL.n16 185
R1418 VTAIL.n10 VTAIL.n9 185
R1419 VTAIL.n23 VTAIL.n22 185
R1420 VTAIL.n25 VTAIL.n24 185
R1421 VTAIL.n6 VTAIL.n5 185
R1422 VTAIL.n31 VTAIL.n30 185
R1423 VTAIL.n33 VTAIL.n32 185
R1424 VTAIL.n111 VTAIL.n110 185
R1425 VTAIL.n109 VTAIL.n108 185
R1426 VTAIL.n84 VTAIL.n83 185
R1427 VTAIL.n103 VTAIL.n102 185
R1428 VTAIL.n101 VTAIL.n100 185
R1429 VTAIL.n88 VTAIL.n87 185
R1430 VTAIL.n95 VTAIL.n94 185
R1431 VTAIL.n93 VTAIL.n92 185
R1432 VTAIL.n73 VTAIL.n72 185
R1433 VTAIL.n71 VTAIL.n70 185
R1434 VTAIL.n46 VTAIL.n45 185
R1435 VTAIL.n65 VTAIL.n64 185
R1436 VTAIL.n63 VTAIL.n62 185
R1437 VTAIL.n50 VTAIL.n49 185
R1438 VTAIL.n57 VTAIL.n56 185
R1439 VTAIL.n55 VTAIL.n54 185
R1440 VTAIL.n127 VTAIL.t0 147.659
R1441 VTAIL.n13 VTAIL.t10 147.659
R1442 VTAIL.n91 VTAIL.t6 147.659
R1443 VTAIL.n53 VTAIL.t1 147.659
R1444 VTAIL.n130 VTAIL.n129 104.615
R1445 VTAIL.n130 VTAIL.n123 104.615
R1446 VTAIL.n137 VTAIL.n123 104.615
R1447 VTAIL.n138 VTAIL.n137 104.615
R1448 VTAIL.n138 VTAIL.n119 104.615
R1449 VTAIL.n145 VTAIL.n119 104.615
R1450 VTAIL.n146 VTAIL.n145 104.615
R1451 VTAIL.n16 VTAIL.n15 104.615
R1452 VTAIL.n16 VTAIL.n9 104.615
R1453 VTAIL.n23 VTAIL.n9 104.615
R1454 VTAIL.n24 VTAIL.n23 104.615
R1455 VTAIL.n24 VTAIL.n5 104.615
R1456 VTAIL.n31 VTAIL.n5 104.615
R1457 VTAIL.n32 VTAIL.n31 104.615
R1458 VTAIL.n110 VTAIL.n109 104.615
R1459 VTAIL.n109 VTAIL.n83 104.615
R1460 VTAIL.n102 VTAIL.n83 104.615
R1461 VTAIL.n102 VTAIL.n101 104.615
R1462 VTAIL.n101 VTAIL.n87 104.615
R1463 VTAIL.n94 VTAIL.n87 104.615
R1464 VTAIL.n94 VTAIL.n93 104.615
R1465 VTAIL.n72 VTAIL.n71 104.615
R1466 VTAIL.n71 VTAIL.n45 104.615
R1467 VTAIL.n64 VTAIL.n45 104.615
R1468 VTAIL.n64 VTAIL.n63 104.615
R1469 VTAIL.n63 VTAIL.n49 104.615
R1470 VTAIL.n56 VTAIL.n49 104.615
R1471 VTAIL.n56 VTAIL.n55 104.615
R1472 VTAIL.n129 VTAIL.t0 52.3082
R1473 VTAIL.n15 VTAIL.t10 52.3082
R1474 VTAIL.n93 VTAIL.t6 52.3082
R1475 VTAIL.n55 VTAIL.t1 52.3082
R1476 VTAIL.n79 VTAIL.n78 48.0378
R1477 VTAIL.n41 VTAIL.n40 48.0378
R1478 VTAIL.n1 VTAIL.n0 48.0376
R1479 VTAIL.n39 VTAIL.n38 48.0376
R1480 VTAIL.n151 VTAIL.n150 30.8278
R1481 VTAIL.n37 VTAIL.n36 30.8278
R1482 VTAIL.n115 VTAIL.n114 30.8278
R1483 VTAIL.n77 VTAIL.n76 30.8278
R1484 VTAIL.n41 VTAIL.n39 23.41
R1485 VTAIL.n151 VTAIL.n115 20.7548
R1486 VTAIL.n128 VTAIL.n127 15.6676
R1487 VTAIL.n14 VTAIL.n13 15.6676
R1488 VTAIL.n92 VTAIL.n91 15.6676
R1489 VTAIL.n54 VTAIL.n53 15.6676
R1490 VTAIL.n131 VTAIL.n126 12.8005
R1491 VTAIL.n17 VTAIL.n12 12.8005
R1492 VTAIL.n95 VTAIL.n90 12.8005
R1493 VTAIL.n57 VTAIL.n52 12.8005
R1494 VTAIL.n132 VTAIL.n124 12.0247
R1495 VTAIL.n18 VTAIL.n10 12.0247
R1496 VTAIL.n96 VTAIL.n88 12.0247
R1497 VTAIL.n58 VTAIL.n50 12.0247
R1498 VTAIL.n136 VTAIL.n135 11.249
R1499 VTAIL.n22 VTAIL.n21 11.249
R1500 VTAIL.n100 VTAIL.n99 11.249
R1501 VTAIL.n62 VTAIL.n61 11.249
R1502 VTAIL.n139 VTAIL.n122 10.4732
R1503 VTAIL.n25 VTAIL.n8 10.4732
R1504 VTAIL.n103 VTAIL.n86 10.4732
R1505 VTAIL.n65 VTAIL.n48 10.4732
R1506 VTAIL.n140 VTAIL.n120 9.69747
R1507 VTAIL.n26 VTAIL.n6 9.69747
R1508 VTAIL.n104 VTAIL.n84 9.69747
R1509 VTAIL.n66 VTAIL.n46 9.69747
R1510 VTAIL.n150 VTAIL.n149 9.45567
R1511 VTAIL.n36 VTAIL.n35 9.45567
R1512 VTAIL.n114 VTAIL.n113 9.45567
R1513 VTAIL.n76 VTAIL.n75 9.45567
R1514 VTAIL.n118 VTAIL.n117 9.3005
R1515 VTAIL.n143 VTAIL.n142 9.3005
R1516 VTAIL.n141 VTAIL.n140 9.3005
R1517 VTAIL.n122 VTAIL.n121 9.3005
R1518 VTAIL.n135 VTAIL.n134 9.3005
R1519 VTAIL.n133 VTAIL.n132 9.3005
R1520 VTAIL.n126 VTAIL.n125 9.3005
R1521 VTAIL.n149 VTAIL.n148 9.3005
R1522 VTAIL.n4 VTAIL.n3 9.3005
R1523 VTAIL.n29 VTAIL.n28 9.3005
R1524 VTAIL.n27 VTAIL.n26 9.3005
R1525 VTAIL.n8 VTAIL.n7 9.3005
R1526 VTAIL.n21 VTAIL.n20 9.3005
R1527 VTAIL.n19 VTAIL.n18 9.3005
R1528 VTAIL.n12 VTAIL.n11 9.3005
R1529 VTAIL.n35 VTAIL.n34 9.3005
R1530 VTAIL.n113 VTAIL.n112 9.3005
R1531 VTAIL.n82 VTAIL.n81 9.3005
R1532 VTAIL.n107 VTAIL.n106 9.3005
R1533 VTAIL.n105 VTAIL.n104 9.3005
R1534 VTAIL.n86 VTAIL.n85 9.3005
R1535 VTAIL.n99 VTAIL.n98 9.3005
R1536 VTAIL.n97 VTAIL.n96 9.3005
R1537 VTAIL.n90 VTAIL.n89 9.3005
R1538 VTAIL.n75 VTAIL.n74 9.3005
R1539 VTAIL.n44 VTAIL.n43 9.3005
R1540 VTAIL.n69 VTAIL.n68 9.3005
R1541 VTAIL.n67 VTAIL.n66 9.3005
R1542 VTAIL.n48 VTAIL.n47 9.3005
R1543 VTAIL.n61 VTAIL.n60 9.3005
R1544 VTAIL.n59 VTAIL.n58 9.3005
R1545 VTAIL.n52 VTAIL.n51 9.3005
R1546 VTAIL.n144 VTAIL.n143 8.92171
R1547 VTAIL.n30 VTAIL.n29 8.92171
R1548 VTAIL.n108 VTAIL.n107 8.92171
R1549 VTAIL.n70 VTAIL.n69 8.92171
R1550 VTAIL.n147 VTAIL.n118 8.14595
R1551 VTAIL.n33 VTAIL.n4 8.14595
R1552 VTAIL.n111 VTAIL.n82 8.14595
R1553 VTAIL.n73 VTAIL.n44 8.14595
R1554 VTAIL.n148 VTAIL.n116 7.3702
R1555 VTAIL.n34 VTAIL.n2 7.3702
R1556 VTAIL.n112 VTAIL.n80 7.3702
R1557 VTAIL.n74 VTAIL.n42 7.3702
R1558 VTAIL.n150 VTAIL.n116 6.59444
R1559 VTAIL.n36 VTAIL.n2 6.59444
R1560 VTAIL.n114 VTAIL.n80 6.59444
R1561 VTAIL.n76 VTAIL.n42 6.59444
R1562 VTAIL.n148 VTAIL.n147 5.81868
R1563 VTAIL.n34 VTAIL.n33 5.81868
R1564 VTAIL.n112 VTAIL.n111 5.81868
R1565 VTAIL.n74 VTAIL.n73 5.81868
R1566 VTAIL.n144 VTAIL.n118 5.04292
R1567 VTAIL.n30 VTAIL.n4 5.04292
R1568 VTAIL.n108 VTAIL.n82 5.04292
R1569 VTAIL.n70 VTAIL.n44 5.04292
R1570 VTAIL.n127 VTAIL.n125 4.38571
R1571 VTAIL.n13 VTAIL.n11 4.38571
R1572 VTAIL.n91 VTAIL.n89 4.38571
R1573 VTAIL.n53 VTAIL.n51 4.38571
R1574 VTAIL.n143 VTAIL.n120 4.26717
R1575 VTAIL.n29 VTAIL.n6 4.26717
R1576 VTAIL.n107 VTAIL.n84 4.26717
R1577 VTAIL.n69 VTAIL.n46 4.26717
R1578 VTAIL.n140 VTAIL.n139 3.49141
R1579 VTAIL.n26 VTAIL.n25 3.49141
R1580 VTAIL.n104 VTAIL.n103 3.49141
R1581 VTAIL.n66 VTAIL.n65 3.49141
R1582 VTAIL.n0 VTAIL.t5 2.97794
R1583 VTAIL.n0 VTAIL.t2 2.97794
R1584 VTAIL.n38 VTAIL.t9 2.97794
R1585 VTAIL.n38 VTAIL.t11 2.97794
R1586 VTAIL.n78 VTAIL.t7 2.97794
R1587 VTAIL.n78 VTAIL.t8 2.97794
R1588 VTAIL.n40 VTAIL.t3 2.97794
R1589 VTAIL.n40 VTAIL.t4 2.97794
R1590 VTAIL.n136 VTAIL.n122 2.71565
R1591 VTAIL.n22 VTAIL.n8 2.71565
R1592 VTAIL.n100 VTAIL.n86 2.71565
R1593 VTAIL.n62 VTAIL.n48 2.71565
R1594 VTAIL.n77 VTAIL.n41 2.65567
R1595 VTAIL.n115 VTAIL.n79 2.65567
R1596 VTAIL.n39 VTAIL.n37 2.65567
R1597 VTAIL.n135 VTAIL.n124 1.93989
R1598 VTAIL.n21 VTAIL.n10 1.93989
R1599 VTAIL.n99 VTAIL.n88 1.93989
R1600 VTAIL.n61 VTAIL.n50 1.93989
R1601 VTAIL VTAIL.n151 1.93369
R1602 VTAIL.n79 VTAIL.n77 1.79791
R1603 VTAIL.n37 VTAIL.n1 1.79791
R1604 VTAIL.n132 VTAIL.n131 1.16414
R1605 VTAIL.n18 VTAIL.n17 1.16414
R1606 VTAIL.n96 VTAIL.n95 1.16414
R1607 VTAIL.n58 VTAIL.n57 1.16414
R1608 VTAIL VTAIL.n1 0.722483
R1609 VTAIL.n128 VTAIL.n126 0.388379
R1610 VTAIL.n14 VTAIL.n12 0.388379
R1611 VTAIL.n92 VTAIL.n90 0.388379
R1612 VTAIL.n54 VTAIL.n52 0.388379
R1613 VTAIL.n133 VTAIL.n125 0.155672
R1614 VTAIL.n134 VTAIL.n133 0.155672
R1615 VTAIL.n134 VTAIL.n121 0.155672
R1616 VTAIL.n141 VTAIL.n121 0.155672
R1617 VTAIL.n142 VTAIL.n141 0.155672
R1618 VTAIL.n142 VTAIL.n117 0.155672
R1619 VTAIL.n149 VTAIL.n117 0.155672
R1620 VTAIL.n19 VTAIL.n11 0.155672
R1621 VTAIL.n20 VTAIL.n19 0.155672
R1622 VTAIL.n20 VTAIL.n7 0.155672
R1623 VTAIL.n27 VTAIL.n7 0.155672
R1624 VTAIL.n28 VTAIL.n27 0.155672
R1625 VTAIL.n28 VTAIL.n3 0.155672
R1626 VTAIL.n35 VTAIL.n3 0.155672
R1627 VTAIL.n113 VTAIL.n81 0.155672
R1628 VTAIL.n106 VTAIL.n81 0.155672
R1629 VTAIL.n106 VTAIL.n105 0.155672
R1630 VTAIL.n105 VTAIL.n85 0.155672
R1631 VTAIL.n98 VTAIL.n85 0.155672
R1632 VTAIL.n98 VTAIL.n97 0.155672
R1633 VTAIL.n97 VTAIL.n89 0.155672
R1634 VTAIL.n75 VTAIL.n43 0.155672
R1635 VTAIL.n68 VTAIL.n43 0.155672
R1636 VTAIL.n68 VTAIL.n67 0.155672
R1637 VTAIL.n67 VTAIL.n47 0.155672
R1638 VTAIL.n60 VTAIL.n47 0.155672
R1639 VTAIL.n60 VTAIL.n59 0.155672
R1640 VTAIL.n59 VTAIL.n51 0.155672
R1641 VDD1.n30 VDD1.n0 289.615
R1642 VDD1.n65 VDD1.n35 289.615
R1643 VDD1.n31 VDD1.n30 185
R1644 VDD1.n29 VDD1.n28 185
R1645 VDD1.n4 VDD1.n3 185
R1646 VDD1.n23 VDD1.n22 185
R1647 VDD1.n21 VDD1.n20 185
R1648 VDD1.n8 VDD1.n7 185
R1649 VDD1.n15 VDD1.n14 185
R1650 VDD1.n13 VDD1.n12 185
R1651 VDD1.n48 VDD1.n47 185
R1652 VDD1.n50 VDD1.n49 185
R1653 VDD1.n43 VDD1.n42 185
R1654 VDD1.n56 VDD1.n55 185
R1655 VDD1.n58 VDD1.n57 185
R1656 VDD1.n39 VDD1.n38 185
R1657 VDD1.n64 VDD1.n63 185
R1658 VDD1.n66 VDD1.n65 185
R1659 VDD1.n11 VDD1.t2 147.659
R1660 VDD1.n46 VDD1.t3 147.659
R1661 VDD1.n30 VDD1.n29 104.615
R1662 VDD1.n29 VDD1.n3 104.615
R1663 VDD1.n22 VDD1.n3 104.615
R1664 VDD1.n22 VDD1.n21 104.615
R1665 VDD1.n21 VDD1.n7 104.615
R1666 VDD1.n14 VDD1.n7 104.615
R1667 VDD1.n14 VDD1.n13 104.615
R1668 VDD1.n49 VDD1.n48 104.615
R1669 VDD1.n49 VDD1.n42 104.615
R1670 VDD1.n56 VDD1.n42 104.615
R1671 VDD1.n57 VDD1.n56 104.615
R1672 VDD1.n57 VDD1.n38 104.615
R1673 VDD1.n64 VDD1.n38 104.615
R1674 VDD1.n65 VDD1.n64 104.615
R1675 VDD1.n71 VDD1.n70 65.3248
R1676 VDD1.n73 VDD1.n72 64.7164
R1677 VDD1.n13 VDD1.t2 52.3082
R1678 VDD1.n48 VDD1.t3 52.3082
R1679 VDD1 VDD1.n34 49.5561
R1680 VDD1.n71 VDD1.n69 49.4426
R1681 VDD1.n73 VDD1.n71 39.988
R1682 VDD1.n12 VDD1.n11 15.6676
R1683 VDD1.n47 VDD1.n46 15.6676
R1684 VDD1.n15 VDD1.n10 12.8005
R1685 VDD1.n50 VDD1.n45 12.8005
R1686 VDD1.n16 VDD1.n8 12.0247
R1687 VDD1.n51 VDD1.n43 12.0247
R1688 VDD1.n20 VDD1.n19 11.249
R1689 VDD1.n55 VDD1.n54 11.249
R1690 VDD1.n23 VDD1.n6 10.4732
R1691 VDD1.n58 VDD1.n41 10.4732
R1692 VDD1.n24 VDD1.n4 9.69747
R1693 VDD1.n59 VDD1.n39 9.69747
R1694 VDD1.n34 VDD1.n33 9.45567
R1695 VDD1.n69 VDD1.n68 9.45567
R1696 VDD1.n33 VDD1.n32 9.3005
R1697 VDD1.n2 VDD1.n1 9.3005
R1698 VDD1.n27 VDD1.n26 9.3005
R1699 VDD1.n25 VDD1.n24 9.3005
R1700 VDD1.n6 VDD1.n5 9.3005
R1701 VDD1.n19 VDD1.n18 9.3005
R1702 VDD1.n17 VDD1.n16 9.3005
R1703 VDD1.n10 VDD1.n9 9.3005
R1704 VDD1.n37 VDD1.n36 9.3005
R1705 VDD1.n62 VDD1.n61 9.3005
R1706 VDD1.n60 VDD1.n59 9.3005
R1707 VDD1.n41 VDD1.n40 9.3005
R1708 VDD1.n54 VDD1.n53 9.3005
R1709 VDD1.n52 VDD1.n51 9.3005
R1710 VDD1.n45 VDD1.n44 9.3005
R1711 VDD1.n68 VDD1.n67 9.3005
R1712 VDD1.n28 VDD1.n27 8.92171
R1713 VDD1.n63 VDD1.n62 8.92171
R1714 VDD1.n31 VDD1.n2 8.14595
R1715 VDD1.n66 VDD1.n37 8.14595
R1716 VDD1.n32 VDD1.n0 7.3702
R1717 VDD1.n67 VDD1.n35 7.3702
R1718 VDD1.n34 VDD1.n0 6.59444
R1719 VDD1.n69 VDD1.n35 6.59444
R1720 VDD1.n32 VDD1.n31 5.81868
R1721 VDD1.n67 VDD1.n66 5.81868
R1722 VDD1.n28 VDD1.n2 5.04292
R1723 VDD1.n63 VDD1.n37 5.04292
R1724 VDD1.n11 VDD1.n9 4.38571
R1725 VDD1.n46 VDD1.n44 4.38571
R1726 VDD1.n27 VDD1.n4 4.26717
R1727 VDD1.n62 VDD1.n39 4.26717
R1728 VDD1.n24 VDD1.n23 3.49141
R1729 VDD1.n59 VDD1.n58 3.49141
R1730 VDD1.n72 VDD1.t0 2.97794
R1731 VDD1.n72 VDD1.t1 2.97794
R1732 VDD1.n70 VDD1.t4 2.97794
R1733 VDD1.n70 VDD1.t5 2.97794
R1734 VDD1.n20 VDD1.n6 2.71565
R1735 VDD1.n55 VDD1.n41 2.71565
R1736 VDD1.n19 VDD1.n8 1.93989
R1737 VDD1.n54 VDD1.n43 1.93989
R1738 VDD1.n16 VDD1.n15 1.16414
R1739 VDD1.n51 VDD1.n50 1.16414
R1740 VDD1 VDD1.n73 0.606103
R1741 VDD1.n12 VDD1.n10 0.388379
R1742 VDD1.n47 VDD1.n45 0.388379
R1743 VDD1.n33 VDD1.n1 0.155672
R1744 VDD1.n26 VDD1.n1 0.155672
R1745 VDD1.n26 VDD1.n25 0.155672
R1746 VDD1.n25 VDD1.n5 0.155672
R1747 VDD1.n18 VDD1.n5 0.155672
R1748 VDD1.n18 VDD1.n17 0.155672
R1749 VDD1.n17 VDD1.n9 0.155672
R1750 VDD1.n52 VDD1.n44 0.155672
R1751 VDD1.n53 VDD1.n52 0.155672
R1752 VDD1.n53 VDD1.n40 0.155672
R1753 VDD1.n60 VDD1.n40 0.155672
R1754 VDD1.n61 VDD1.n60 0.155672
R1755 VDD1.n61 VDD1.n36 0.155672
R1756 VDD1.n68 VDD1.n36 0.155672
R1757 VN.n29 VN.n16 161.3
R1758 VN.n28 VN.n27 161.3
R1759 VN.n26 VN.n17 161.3
R1760 VN.n25 VN.n24 161.3
R1761 VN.n23 VN.n18 161.3
R1762 VN.n22 VN.n21 161.3
R1763 VN.n13 VN.n0 161.3
R1764 VN.n12 VN.n11 161.3
R1765 VN.n10 VN.n1 161.3
R1766 VN.n9 VN.n8 161.3
R1767 VN.n7 VN.n2 161.3
R1768 VN.n6 VN.n5 161.3
R1769 VN.n15 VN.n14 106.841
R1770 VN.n31 VN.n30 106.841
R1771 VN.n4 VN.t4 91.9343
R1772 VN.n20 VN.t2 91.9343
R1773 VN.n3 VN.t0 58.2787
R1774 VN.n14 VN.t1 58.2787
R1775 VN.n19 VN.t3 58.2787
R1776 VN.n30 VN.t5 58.2787
R1777 VN.n20 VN.n19 48.924
R1778 VN.n4 VN.n3 48.924
R1779 VN VN.n31 45.4527
R1780 VN.n8 VN.n1 44.3785
R1781 VN.n24 VN.n17 44.3785
R1782 VN.n8 VN.n7 36.6083
R1783 VN.n24 VN.n23 36.6083
R1784 VN.n6 VN.n3 24.4675
R1785 VN.n7 VN.n6 24.4675
R1786 VN.n12 VN.n1 24.4675
R1787 VN.n13 VN.n12 24.4675
R1788 VN.n23 VN.n22 24.4675
R1789 VN.n22 VN.n19 24.4675
R1790 VN.n29 VN.n28 24.4675
R1791 VN.n28 VN.n17 24.4675
R1792 VN.n21 VN.n20 5.02272
R1793 VN.n5 VN.n4 5.02272
R1794 VN.n14 VN.n13 3.91522
R1795 VN.n30 VN.n29 3.91522
R1796 VN.n31 VN.n16 0.278367
R1797 VN.n15 VN.n0 0.278367
R1798 VN.n27 VN.n16 0.189894
R1799 VN.n27 VN.n26 0.189894
R1800 VN.n26 VN.n25 0.189894
R1801 VN.n25 VN.n18 0.189894
R1802 VN.n21 VN.n18 0.189894
R1803 VN.n5 VN.n2 0.189894
R1804 VN.n9 VN.n2 0.189894
R1805 VN.n10 VN.n9 0.189894
R1806 VN.n11 VN.n10 0.189894
R1807 VN.n11 VN.n0 0.189894
R1808 VN VN.n15 0.153454
R1809 VDD2.n67 VDD2.n37 289.615
R1810 VDD2.n30 VDD2.n0 289.615
R1811 VDD2.n68 VDD2.n67 185
R1812 VDD2.n66 VDD2.n65 185
R1813 VDD2.n41 VDD2.n40 185
R1814 VDD2.n60 VDD2.n59 185
R1815 VDD2.n58 VDD2.n57 185
R1816 VDD2.n45 VDD2.n44 185
R1817 VDD2.n52 VDD2.n51 185
R1818 VDD2.n50 VDD2.n49 185
R1819 VDD2.n13 VDD2.n12 185
R1820 VDD2.n15 VDD2.n14 185
R1821 VDD2.n8 VDD2.n7 185
R1822 VDD2.n21 VDD2.n20 185
R1823 VDD2.n23 VDD2.n22 185
R1824 VDD2.n4 VDD2.n3 185
R1825 VDD2.n29 VDD2.n28 185
R1826 VDD2.n31 VDD2.n30 185
R1827 VDD2.n48 VDD2.t0 147.659
R1828 VDD2.n11 VDD2.t1 147.659
R1829 VDD2.n67 VDD2.n66 104.615
R1830 VDD2.n66 VDD2.n40 104.615
R1831 VDD2.n59 VDD2.n40 104.615
R1832 VDD2.n59 VDD2.n58 104.615
R1833 VDD2.n58 VDD2.n44 104.615
R1834 VDD2.n51 VDD2.n44 104.615
R1835 VDD2.n51 VDD2.n50 104.615
R1836 VDD2.n14 VDD2.n13 104.615
R1837 VDD2.n14 VDD2.n7 104.615
R1838 VDD2.n21 VDD2.n7 104.615
R1839 VDD2.n22 VDD2.n21 104.615
R1840 VDD2.n22 VDD2.n3 104.615
R1841 VDD2.n29 VDD2.n3 104.615
R1842 VDD2.n30 VDD2.n29 104.615
R1843 VDD2.n36 VDD2.n35 65.3248
R1844 VDD2 VDD2.n73 65.322
R1845 VDD2.n50 VDD2.t0 52.3082
R1846 VDD2.n13 VDD2.t1 52.3082
R1847 VDD2.n36 VDD2.n34 49.4426
R1848 VDD2.n72 VDD2.n71 47.5066
R1849 VDD2.n72 VDD2.n36 38.0774
R1850 VDD2.n49 VDD2.n48 15.6676
R1851 VDD2.n12 VDD2.n11 15.6676
R1852 VDD2.n52 VDD2.n47 12.8005
R1853 VDD2.n15 VDD2.n10 12.8005
R1854 VDD2.n53 VDD2.n45 12.0247
R1855 VDD2.n16 VDD2.n8 12.0247
R1856 VDD2.n57 VDD2.n56 11.249
R1857 VDD2.n20 VDD2.n19 11.249
R1858 VDD2.n60 VDD2.n43 10.4732
R1859 VDD2.n23 VDD2.n6 10.4732
R1860 VDD2.n61 VDD2.n41 9.69747
R1861 VDD2.n24 VDD2.n4 9.69747
R1862 VDD2.n71 VDD2.n70 9.45567
R1863 VDD2.n34 VDD2.n33 9.45567
R1864 VDD2.n70 VDD2.n69 9.3005
R1865 VDD2.n39 VDD2.n38 9.3005
R1866 VDD2.n64 VDD2.n63 9.3005
R1867 VDD2.n62 VDD2.n61 9.3005
R1868 VDD2.n43 VDD2.n42 9.3005
R1869 VDD2.n56 VDD2.n55 9.3005
R1870 VDD2.n54 VDD2.n53 9.3005
R1871 VDD2.n47 VDD2.n46 9.3005
R1872 VDD2.n2 VDD2.n1 9.3005
R1873 VDD2.n27 VDD2.n26 9.3005
R1874 VDD2.n25 VDD2.n24 9.3005
R1875 VDD2.n6 VDD2.n5 9.3005
R1876 VDD2.n19 VDD2.n18 9.3005
R1877 VDD2.n17 VDD2.n16 9.3005
R1878 VDD2.n10 VDD2.n9 9.3005
R1879 VDD2.n33 VDD2.n32 9.3005
R1880 VDD2.n65 VDD2.n64 8.92171
R1881 VDD2.n28 VDD2.n27 8.92171
R1882 VDD2.n68 VDD2.n39 8.14595
R1883 VDD2.n31 VDD2.n2 8.14595
R1884 VDD2.n69 VDD2.n37 7.3702
R1885 VDD2.n32 VDD2.n0 7.3702
R1886 VDD2.n71 VDD2.n37 6.59444
R1887 VDD2.n34 VDD2.n0 6.59444
R1888 VDD2.n69 VDD2.n68 5.81868
R1889 VDD2.n32 VDD2.n31 5.81868
R1890 VDD2.n65 VDD2.n39 5.04292
R1891 VDD2.n28 VDD2.n2 5.04292
R1892 VDD2.n48 VDD2.n46 4.38571
R1893 VDD2.n11 VDD2.n9 4.38571
R1894 VDD2.n64 VDD2.n41 4.26717
R1895 VDD2.n27 VDD2.n4 4.26717
R1896 VDD2.n61 VDD2.n60 3.49141
R1897 VDD2.n24 VDD2.n23 3.49141
R1898 VDD2.n73 VDD2.t2 2.97794
R1899 VDD2.n73 VDD2.t3 2.97794
R1900 VDD2.n35 VDD2.t5 2.97794
R1901 VDD2.n35 VDD2.t4 2.97794
R1902 VDD2.n57 VDD2.n43 2.71565
R1903 VDD2.n20 VDD2.n6 2.71565
R1904 VDD2 VDD2.n72 2.05007
R1905 VDD2.n56 VDD2.n45 1.93989
R1906 VDD2.n19 VDD2.n8 1.93989
R1907 VDD2.n53 VDD2.n52 1.16414
R1908 VDD2.n16 VDD2.n15 1.16414
R1909 VDD2.n49 VDD2.n47 0.388379
R1910 VDD2.n12 VDD2.n10 0.388379
R1911 VDD2.n70 VDD2.n38 0.155672
R1912 VDD2.n63 VDD2.n38 0.155672
R1913 VDD2.n63 VDD2.n62 0.155672
R1914 VDD2.n62 VDD2.n42 0.155672
R1915 VDD2.n55 VDD2.n42 0.155672
R1916 VDD2.n55 VDD2.n54 0.155672
R1917 VDD2.n54 VDD2.n46 0.155672
R1918 VDD2.n17 VDD2.n9 0.155672
R1919 VDD2.n18 VDD2.n17 0.155672
R1920 VDD2.n18 VDD2.n5 0.155672
R1921 VDD2.n25 VDD2.n5 0.155672
R1922 VDD2.n26 VDD2.n25 0.155672
R1923 VDD2.n26 VDD2.n1 0.155672
R1924 VDD2.n33 VDD2.n1 0.155672
C0 VN VP 6.08227f
C1 VTAIL VP 4.534431f
C2 VDD1 VP 4.26056f
C3 VTAIL VN 4.52023f
C4 VDD1 VN 0.150798f
C5 VDD1 VTAIL 5.85995f
C6 VDD2 VP 0.47048f
C7 VDD2 VN 3.94314f
C8 VDD2 VTAIL 5.91312f
C9 VDD2 VDD1 1.46384f
C10 VDD2 B 5.147177f
C11 VDD1 B 5.284004f
C12 VTAIL B 5.437437f
C13 VN B 12.75181f
C14 VP B 11.436545f
C15 VDD2.n0 B 0.029994f
C16 VDD2.n1 B 0.021651f
C17 VDD2.n2 B 0.011634f
C18 VDD2.n3 B 0.027499f
C19 VDD2.n4 B 0.012318f
C20 VDD2.n5 B 0.021651f
C21 VDD2.n6 B 0.011634f
C22 VDD2.n7 B 0.027499f
C23 VDD2.n8 B 0.012318f
C24 VDD2.n9 B 0.579887f
C25 VDD2.n10 B 0.011634f
C26 VDD2.t1 B 0.04479f
C27 VDD2.n11 B 0.096024f
C28 VDD2.n12 B 0.016244f
C29 VDD2.n13 B 0.020624f
C30 VDD2.n14 B 0.027499f
C31 VDD2.n15 B 0.012318f
C32 VDD2.n16 B 0.011634f
C33 VDD2.n17 B 0.021651f
C34 VDD2.n18 B 0.021651f
C35 VDD2.n19 B 0.011634f
C36 VDD2.n20 B 0.012318f
C37 VDD2.n21 B 0.027499f
C38 VDD2.n22 B 0.027499f
C39 VDD2.n23 B 0.012318f
C40 VDD2.n24 B 0.011634f
C41 VDD2.n25 B 0.021651f
C42 VDD2.n26 B 0.021651f
C43 VDD2.n27 B 0.011634f
C44 VDD2.n28 B 0.012318f
C45 VDD2.n29 B 0.027499f
C46 VDD2.n30 B 0.058756f
C47 VDD2.n31 B 0.012318f
C48 VDD2.n32 B 0.011634f
C49 VDD2.n33 B 0.047974f
C50 VDD2.n34 B 0.054583f
C51 VDD2.t5 B 0.113775f
C52 VDD2.t4 B 0.113775f
C53 VDD2.n35 B 0.96351f
C54 VDD2.n36 B 2.0924f
C55 VDD2.n37 B 0.029994f
C56 VDD2.n38 B 0.021651f
C57 VDD2.n39 B 0.011634f
C58 VDD2.n40 B 0.027499f
C59 VDD2.n41 B 0.012318f
C60 VDD2.n42 B 0.021651f
C61 VDD2.n43 B 0.011634f
C62 VDD2.n44 B 0.027499f
C63 VDD2.n45 B 0.012318f
C64 VDD2.n46 B 0.579887f
C65 VDD2.n47 B 0.011634f
C66 VDD2.t0 B 0.04479f
C67 VDD2.n48 B 0.096024f
C68 VDD2.n49 B 0.016244f
C69 VDD2.n50 B 0.020624f
C70 VDD2.n51 B 0.027499f
C71 VDD2.n52 B 0.012318f
C72 VDD2.n53 B 0.011634f
C73 VDD2.n54 B 0.021651f
C74 VDD2.n55 B 0.021651f
C75 VDD2.n56 B 0.011634f
C76 VDD2.n57 B 0.012318f
C77 VDD2.n58 B 0.027499f
C78 VDD2.n59 B 0.027499f
C79 VDD2.n60 B 0.012318f
C80 VDD2.n61 B 0.011634f
C81 VDD2.n62 B 0.021651f
C82 VDD2.n63 B 0.021651f
C83 VDD2.n64 B 0.011634f
C84 VDD2.n65 B 0.012318f
C85 VDD2.n66 B 0.027499f
C86 VDD2.n67 B 0.058756f
C87 VDD2.n68 B 0.012318f
C88 VDD2.n69 B 0.011634f
C89 VDD2.n70 B 0.047974f
C90 VDD2.n71 B 0.047698f
C91 VDD2.n72 B 1.89059f
C92 VDD2.t2 B 0.113775f
C93 VDD2.t3 B 0.113775f
C94 VDD2.n73 B 0.963482f
C95 VN.n0 B 0.032693f
C96 VN.t1 B 1.20718f
C97 VN.n1 B 0.048058f
C98 VN.n2 B 0.024798f
C99 VN.t0 B 1.20718f
C100 VN.n3 B 0.534576f
C101 VN.t4 B 1.43064f
C102 VN.n4 B 0.499095f
C103 VN.n5 B 0.259006f
C104 VN.n6 B 0.046217f
C105 VN.n7 B 0.049999f
C106 VN.n8 B 0.020561f
C107 VN.n9 B 0.024798f
C108 VN.n10 B 0.024798f
C109 VN.n11 B 0.024798f
C110 VN.n12 B 0.046217f
C111 VN.n13 B 0.02705f
C112 VN.n14 B 0.526355f
C113 VN.n15 B 0.045219f
C114 VN.n16 B 0.032693f
C115 VN.t5 B 1.20718f
C116 VN.n17 B 0.048058f
C117 VN.n18 B 0.024798f
C118 VN.t3 B 1.20718f
C119 VN.n19 B 0.534576f
C120 VN.t2 B 1.43064f
C121 VN.n20 B 0.499095f
C122 VN.n21 B 0.259006f
C123 VN.n22 B 0.046217f
C124 VN.n23 B 0.049999f
C125 VN.n24 B 0.020561f
C126 VN.n25 B 0.024798f
C127 VN.n26 B 0.024798f
C128 VN.n27 B 0.024798f
C129 VN.n28 B 0.046217f
C130 VN.n29 B 0.02705f
C131 VN.n30 B 0.526355f
C132 VN.n31 B 1.20224f
C133 VDD1.n0 B 0.030965f
C134 VDD1.n1 B 0.022352f
C135 VDD1.n2 B 0.012011f
C136 VDD1.n3 B 0.02839f
C137 VDD1.n4 B 0.012718f
C138 VDD1.n5 B 0.022352f
C139 VDD1.n6 B 0.012011f
C140 VDD1.n7 B 0.02839f
C141 VDD1.n8 B 0.012718f
C142 VDD1.n9 B 0.598671f
C143 VDD1.n10 B 0.012011f
C144 VDD1.t2 B 0.046241f
C145 VDD1.n11 B 0.099134f
C146 VDD1.n12 B 0.01677f
C147 VDD1.n13 B 0.021292f
C148 VDD1.n14 B 0.02839f
C149 VDD1.n15 B 0.012718f
C150 VDD1.n16 B 0.012011f
C151 VDD1.n17 B 0.022352f
C152 VDD1.n18 B 0.022352f
C153 VDD1.n19 B 0.012011f
C154 VDD1.n20 B 0.012718f
C155 VDD1.n21 B 0.02839f
C156 VDD1.n22 B 0.02839f
C157 VDD1.n23 B 0.012718f
C158 VDD1.n24 B 0.012011f
C159 VDD1.n25 B 0.022352f
C160 VDD1.n26 B 0.022352f
C161 VDD1.n27 B 0.012011f
C162 VDD1.n28 B 0.012718f
C163 VDD1.n29 B 0.02839f
C164 VDD1.n30 B 0.060659f
C165 VDD1.n31 B 0.012718f
C166 VDD1.n32 B 0.012011f
C167 VDD1.n33 B 0.049528f
C168 VDD1.n34 B 0.057078f
C169 VDD1.n35 B 0.030965f
C170 VDD1.n36 B 0.022352f
C171 VDD1.n37 B 0.012011f
C172 VDD1.n38 B 0.02839f
C173 VDD1.n39 B 0.012718f
C174 VDD1.n40 B 0.022352f
C175 VDD1.n41 B 0.012011f
C176 VDD1.n42 B 0.02839f
C177 VDD1.n43 B 0.012718f
C178 VDD1.n44 B 0.598671f
C179 VDD1.n45 B 0.012011f
C180 VDD1.t3 B 0.046241f
C181 VDD1.n46 B 0.099134f
C182 VDD1.n47 B 0.01677f
C183 VDD1.n48 B 0.021292f
C184 VDD1.n49 B 0.02839f
C185 VDD1.n50 B 0.012718f
C186 VDD1.n51 B 0.012011f
C187 VDD1.n52 B 0.022352f
C188 VDD1.n53 B 0.022352f
C189 VDD1.n54 B 0.012011f
C190 VDD1.n55 B 0.012718f
C191 VDD1.n56 B 0.02839f
C192 VDD1.n57 B 0.02839f
C193 VDD1.n58 B 0.012718f
C194 VDD1.n59 B 0.012011f
C195 VDD1.n60 B 0.022352f
C196 VDD1.n61 B 0.022352f
C197 VDD1.n62 B 0.012011f
C198 VDD1.n63 B 0.012718f
C199 VDD1.n64 B 0.02839f
C200 VDD1.n65 B 0.060659f
C201 VDD1.n66 B 0.012718f
C202 VDD1.n67 B 0.012011f
C203 VDD1.n68 B 0.049528f
C204 VDD1.n69 B 0.056351f
C205 VDD1.t4 B 0.117461f
C206 VDD1.t5 B 0.117461f
C207 VDD1.n70 B 0.99472f
C208 VDD1.n71 B 2.27018f
C209 VDD1.t0 B 0.117461f
C210 VDD1.t1 B 0.117461f
C211 VDD1.n72 B 0.990727f
C212 VDD1.n73 B 2.16262f
C213 VTAIL.t5 B 0.140127f
C214 VTAIL.t2 B 0.140127f
C215 VTAIL.n0 B 1.10754f
C216 VTAIL.n1 B 0.473874f
C217 VTAIL.n2 B 0.036941f
C218 VTAIL.n3 B 0.026665f
C219 VTAIL.n4 B 0.014329f
C220 VTAIL.n5 B 0.033868f
C221 VTAIL.n6 B 0.015172f
C222 VTAIL.n7 B 0.026665f
C223 VTAIL.n8 B 0.014329f
C224 VTAIL.n9 B 0.033868f
C225 VTAIL.n10 B 0.015172f
C226 VTAIL.n11 B 0.714196f
C227 VTAIL.n12 B 0.014329f
C228 VTAIL.t10 B 0.055164f
C229 VTAIL.n13 B 0.118264f
C230 VTAIL.n14 B 0.020007f
C231 VTAIL.n15 B 0.025401f
C232 VTAIL.n16 B 0.033868f
C233 VTAIL.n17 B 0.015172f
C234 VTAIL.n18 B 0.014329f
C235 VTAIL.n19 B 0.026665f
C236 VTAIL.n20 B 0.026665f
C237 VTAIL.n21 B 0.014329f
C238 VTAIL.n22 B 0.015172f
C239 VTAIL.n23 B 0.033868f
C240 VTAIL.n24 B 0.033868f
C241 VTAIL.n25 B 0.015172f
C242 VTAIL.n26 B 0.014329f
C243 VTAIL.n27 B 0.026665f
C244 VTAIL.n28 B 0.026665f
C245 VTAIL.n29 B 0.014329f
C246 VTAIL.n30 B 0.015172f
C247 VTAIL.n31 B 0.033868f
C248 VTAIL.n32 B 0.072364f
C249 VTAIL.n33 B 0.015172f
C250 VTAIL.n34 B 0.014329f
C251 VTAIL.n35 B 0.059086f
C252 VTAIL.n36 B 0.040313f
C253 VTAIL.n37 B 0.40391f
C254 VTAIL.t9 B 0.140127f
C255 VTAIL.t11 B 0.140127f
C256 VTAIL.n38 B 1.10754f
C257 VTAIL.n39 B 1.7966f
C258 VTAIL.t3 B 0.140127f
C259 VTAIL.t4 B 0.140127f
C260 VTAIL.n40 B 1.10754f
C261 VTAIL.n41 B 1.79659f
C262 VTAIL.n42 B 0.036941f
C263 VTAIL.n43 B 0.026665f
C264 VTAIL.n44 B 0.014329f
C265 VTAIL.n45 B 0.033868f
C266 VTAIL.n46 B 0.015172f
C267 VTAIL.n47 B 0.026665f
C268 VTAIL.n48 B 0.014329f
C269 VTAIL.n49 B 0.033868f
C270 VTAIL.n50 B 0.015172f
C271 VTAIL.n51 B 0.714196f
C272 VTAIL.n52 B 0.014329f
C273 VTAIL.t1 B 0.055164f
C274 VTAIL.n53 B 0.118264f
C275 VTAIL.n54 B 0.020007f
C276 VTAIL.n55 B 0.025401f
C277 VTAIL.n56 B 0.033868f
C278 VTAIL.n57 B 0.015172f
C279 VTAIL.n58 B 0.014329f
C280 VTAIL.n59 B 0.026665f
C281 VTAIL.n60 B 0.026665f
C282 VTAIL.n61 B 0.014329f
C283 VTAIL.n62 B 0.015172f
C284 VTAIL.n63 B 0.033868f
C285 VTAIL.n64 B 0.033868f
C286 VTAIL.n65 B 0.015172f
C287 VTAIL.n66 B 0.014329f
C288 VTAIL.n67 B 0.026665f
C289 VTAIL.n68 B 0.026665f
C290 VTAIL.n69 B 0.014329f
C291 VTAIL.n70 B 0.015172f
C292 VTAIL.n71 B 0.033868f
C293 VTAIL.n72 B 0.072364f
C294 VTAIL.n73 B 0.015172f
C295 VTAIL.n74 B 0.014329f
C296 VTAIL.n75 B 0.059086f
C297 VTAIL.n76 B 0.040313f
C298 VTAIL.n77 B 0.40391f
C299 VTAIL.t7 B 0.140127f
C300 VTAIL.t8 B 0.140127f
C301 VTAIL.n78 B 1.10754f
C302 VTAIL.n79 B 0.63997f
C303 VTAIL.n80 B 0.036941f
C304 VTAIL.n81 B 0.026665f
C305 VTAIL.n82 B 0.014329f
C306 VTAIL.n83 B 0.033868f
C307 VTAIL.n84 B 0.015172f
C308 VTAIL.n85 B 0.026665f
C309 VTAIL.n86 B 0.014329f
C310 VTAIL.n87 B 0.033868f
C311 VTAIL.n88 B 0.015172f
C312 VTAIL.n89 B 0.714196f
C313 VTAIL.n90 B 0.014329f
C314 VTAIL.t6 B 0.055164f
C315 VTAIL.n91 B 0.118264f
C316 VTAIL.n92 B 0.020007f
C317 VTAIL.n93 B 0.025401f
C318 VTAIL.n94 B 0.033868f
C319 VTAIL.n95 B 0.015172f
C320 VTAIL.n96 B 0.014329f
C321 VTAIL.n97 B 0.026665f
C322 VTAIL.n98 B 0.026665f
C323 VTAIL.n99 B 0.014329f
C324 VTAIL.n100 B 0.015172f
C325 VTAIL.n101 B 0.033868f
C326 VTAIL.n102 B 0.033868f
C327 VTAIL.n103 B 0.015172f
C328 VTAIL.n104 B 0.014329f
C329 VTAIL.n105 B 0.026665f
C330 VTAIL.n106 B 0.026665f
C331 VTAIL.n107 B 0.014329f
C332 VTAIL.n108 B 0.015172f
C333 VTAIL.n109 B 0.033868f
C334 VTAIL.n110 B 0.072364f
C335 VTAIL.n111 B 0.015172f
C336 VTAIL.n112 B 0.014329f
C337 VTAIL.n113 B 0.059086f
C338 VTAIL.n114 B 0.040313f
C339 VTAIL.n115 B 1.3324f
C340 VTAIL.n116 B 0.036941f
C341 VTAIL.n117 B 0.026665f
C342 VTAIL.n118 B 0.014329f
C343 VTAIL.n119 B 0.033868f
C344 VTAIL.n120 B 0.015172f
C345 VTAIL.n121 B 0.026665f
C346 VTAIL.n122 B 0.014329f
C347 VTAIL.n123 B 0.033868f
C348 VTAIL.n124 B 0.015172f
C349 VTAIL.n125 B 0.714196f
C350 VTAIL.n126 B 0.014329f
C351 VTAIL.t0 B 0.055164f
C352 VTAIL.n127 B 0.118264f
C353 VTAIL.n128 B 0.020007f
C354 VTAIL.n129 B 0.025401f
C355 VTAIL.n130 B 0.033868f
C356 VTAIL.n131 B 0.015172f
C357 VTAIL.n132 B 0.014329f
C358 VTAIL.n133 B 0.026665f
C359 VTAIL.n134 B 0.026665f
C360 VTAIL.n135 B 0.014329f
C361 VTAIL.n136 B 0.015172f
C362 VTAIL.n137 B 0.033868f
C363 VTAIL.n138 B 0.033868f
C364 VTAIL.n139 B 0.015172f
C365 VTAIL.n140 B 0.014329f
C366 VTAIL.n141 B 0.026665f
C367 VTAIL.n142 B 0.026665f
C368 VTAIL.n143 B 0.014329f
C369 VTAIL.n144 B 0.015172f
C370 VTAIL.n145 B 0.033868f
C371 VTAIL.n146 B 0.072364f
C372 VTAIL.n147 B 0.015172f
C373 VTAIL.n148 B 0.014329f
C374 VTAIL.n149 B 0.059086f
C375 VTAIL.n150 B 0.040313f
C376 VTAIL.n151 B 1.27036f
C377 VP.n0 B 0.033676f
C378 VP.t0 B 1.24347f
C379 VP.n1 B 0.049502f
C380 VP.n2 B 0.025543f
C381 VP.t1 B 1.24347f
C382 VP.n3 B 0.48397f
C383 VP.n4 B 0.025543f
C384 VP.n5 B 0.049502f
C385 VP.n6 B 0.033676f
C386 VP.t2 B 1.24347f
C387 VP.n7 B 0.033676f
C388 VP.t4 B 1.24347f
C389 VP.n8 B 0.049502f
C390 VP.n9 B 0.025543f
C391 VP.t5 B 1.24347f
C392 VP.n10 B 0.550646f
C393 VP.t3 B 1.47364f
C394 VP.n11 B 0.514099f
C395 VP.n12 B 0.266793f
C396 VP.n13 B 0.047606f
C397 VP.n14 B 0.051502f
C398 VP.n15 B 0.021179f
C399 VP.n16 B 0.025543f
C400 VP.n17 B 0.025543f
C401 VP.n18 B 0.025543f
C402 VP.n19 B 0.047606f
C403 VP.n20 B 0.027863f
C404 VP.n21 B 0.542178f
C405 VP.n22 B 1.22442f
C406 VP.n23 B 1.24475f
C407 VP.n24 B 0.542178f
C408 VP.n25 B 0.027863f
C409 VP.n26 B 0.047606f
C410 VP.n27 B 0.025543f
C411 VP.n28 B 0.025543f
C412 VP.n29 B 0.025543f
C413 VP.n30 B 0.021179f
C414 VP.n31 B 0.051502f
C415 VP.n32 B 0.047606f
C416 VP.n33 B 0.025543f
C417 VP.n34 B 0.025543f
C418 VP.n35 B 0.025543f
C419 VP.n36 B 0.047606f
C420 VP.n37 B 0.051502f
C421 VP.n38 B 0.021179f
C422 VP.n39 B 0.025543f
C423 VP.n40 B 0.025543f
C424 VP.n41 B 0.025543f
C425 VP.n42 B 0.047606f
C426 VP.n43 B 0.027863f
C427 VP.n44 B 0.542178f
C428 VP.n45 B 0.046578f
.ends

