* NGSPICE file created from diff_pair_sample_0709.ext - technology: sky130A

.subckt diff_pair_sample_0709 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=3.2058 ps=17.22 w=8.22 l=1.04
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=0 ps=0 w=8.22 l=1.04
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=0 ps=0 w=8.22 l=1.04
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=0 ps=0 w=8.22 l=1.04
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=3.2058 ps=17.22 w=8.22 l=1.04
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=3.2058 ps=17.22 w=8.22 l=1.04
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=0 ps=0 w=8.22 l=1.04
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2058 pd=17.22 as=3.2058 ps=17.22 w=8.22 l=1.04
R0 VN VN.t0 428.07
R1 VN VN.t1 390.07
R2 VTAIL.n1 VTAIL.t2 50.5892
R3 VTAIL.n3 VTAIL.t3 50.5892
R4 VTAIL.n0 VTAIL.t0 50.5892
R5 VTAIL.n2 VTAIL.t1 50.5892
R6 VTAIL.n1 VTAIL.n0 21.8324
R7 VTAIL.n3 VTAIL.n2 20.6514
R8 VTAIL.n2 VTAIL.n1 1.06084
R9 VTAIL VTAIL.n0 0.823776
R10 VTAIL VTAIL.n3 0.237569
R11 VDD2.n0 VDD2.t0 100.392
R12 VDD2.n0 VDD2.t1 67.268
R13 VDD2 VDD2.n0 0.353948
R14 B.n496 B.n495 585
R15 B.n497 B.n496 585
R16 B.n212 B.n69 585
R17 B.n211 B.n210 585
R18 B.n209 B.n208 585
R19 B.n207 B.n206 585
R20 B.n205 B.n204 585
R21 B.n203 B.n202 585
R22 B.n201 B.n200 585
R23 B.n199 B.n198 585
R24 B.n197 B.n196 585
R25 B.n195 B.n194 585
R26 B.n193 B.n192 585
R27 B.n191 B.n190 585
R28 B.n189 B.n188 585
R29 B.n187 B.n186 585
R30 B.n185 B.n184 585
R31 B.n183 B.n182 585
R32 B.n181 B.n180 585
R33 B.n179 B.n178 585
R34 B.n177 B.n176 585
R35 B.n175 B.n174 585
R36 B.n173 B.n172 585
R37 B.n171 B.n170 585
R38 B.n169 B.n168 585
R39 B.n167 B.n166 585
R40 B.n165 B.n164 585
R41 B.n163 B.n162 585
R42 B.n161 B.n160 585
R43 B.n159 B.n158 585
R44 B.n157 B.n156 585
R45 B.n155 B.n154 585
R46 B.n153 B.n152 585
R47 B.n151 B.n150 585
R48 B.n149 B.n148 585
R49 B.n147 B.n146 585
R50 B.n145 B.n144 585
R51 B.n143 B.n142 585
R52 B.n141 B.n140 585
R53 B.n139 B.n138 585
R54 B.n137 B.n136 585
R55 B.n134 B.n133 585
R56 B.n132 B.n131 585
R57 B.n130 B.n129 585
R58 B.n128 B.n127 585
R59 B.n126 B.n125 585
R60 B.n124 B.n123 585
R61 B.n122 B.n121 585
R62 B.n120 B.n119 585
R63 B.n118 B.n117 585
R64 B.n116 B.n115 585
R65 B.n114 B.n113 585
R66 B.n112 B.n111 585
R67 B.n110 B.n109 585
R68 B.n108 B.n107 585
R69 B.n106 B.n105 585
R70 B.n104 B.n103 585
R71 B.n102 B.n101 585
R72 B.n100 B.n99 585
R73 B.n98 B.n97 585
R74 B.n96 B.n95 585
R75 B.n94 B.n93 585
R76 B.n92 B.n91 585
R77 B.n90 B.n89 585
R78 B.n88 B.n87 585
R79 B.n86 B.n85 585
R80 B.n84 B.n83 585
R81 B.n82 B.n81 585
R82 B.n80 B.n79 585
R83 B.n78 B.n77 585
R84 B.n76 B.n75 585
R85 B.n32 B.n31 585
R86 B.n494 B.n33 585
R87 B.n498 B.n33 585
R88 B.n493 B.n492 585
R89 B.n492 B.n29 585
R90 B.n491 B.n28 585
R91 B.n504 B.n28 585
R92 B.n490 B.n27 585
R93 B.n505 B.n27 585
R94 B.n489 B.n26 585
R95 B.n506 B.n26 585
R96 B.n488 B.n487 585
R97 B.n487 B.n25 585
R98 B.n486 B.n21 585
R99 B.n512 B.n21 585
R100 B.n485 B.n20 585
R101 B.n513 B.n20 585
R102 B.n484 B.n19 585
R103 B.n514 B.n19 585
R104 B.n483 B.n482 585
R105 B.n482 B.n15 585
R106 B.n481 B.n14 585
R107 B.n520 B.n14 585
R108 B.n480 B.n13 585
R109 B.n521 B.n13 585
R110 B.n479 B.n12 585
R111 B.n522 B.n12 585
R112 B.n478 B.n477 585
R113 B.n477 B.n8 585
R114 B.n476 B.n7 585
R115 B.n528 B.n7 585
R116 B.n475 B.n6 585
R117 B.n529 B.n6 585
R118 B.n474 B.n5 585
R119 B.n530 B.n5 585
R120 B.n473 B.n472 585
R121 B.n472 B.n4 585
R122 B.n471 B.n213 585
R123 B.n471 B.n470 585
R124 B.n461 B.n214 585
R125 B.n215 B.n214 585
R126 B.n463 B.n462 585
R127 B.n464 B.n463 585
R128 B.n460 B.n220 585
R129 B.n220 B.n219 585
R130 B.n459 B.n458 585
R131 B.n458 B.n457 585
R132 B.n222 B.n221 585
R133 B.n223 B.n222 585
R134 B.n450 B.n449 585
R135 B.n451 B.n450 585
R136 B.n448 B.n228 585
R137 B.n228 B.n227 585
R138 B.n447 B.n446 585
R139 B.n446 B.n445 585
R140 B.n230 B.n229 585
R141 B.n438 B.n230 585
R142 B.n437 B.n436 585
R143 B.n439 B.n437 585
R144 B.n435 B.n235 585
R145 B.n235 B.n234 585
R146 B.n434 B.n433 585
R147 B.n433 B.n432 585
R148 B.n237 B.n236 585
R149 B.n238 B.n237 585
R150 B.n425 B.n424 585
R151 B.n426 B.n425 585
R152 B.n241 B.n240 585
R153 B.n282 B.n281 585
R154 B.n283 B.n279 585
R155 B.n279 B.n242 585
R156 B.n285 B.n284 585
R157 B.n287 B.n278 585
R158 B.n290 B.n289 585
R159 B.n291 B.n277 585
R160 B.n293 B.n292 585
R161 B.n295 B.n276 585
R162 B.n298 B.n297 585
R163 B.n299 B.n275 585
R164 B.n301 B.n300 585
R165 B.n303 B.n274 585
R166 B.n306 B.n305 585
R167 B.n307 B.n273 585
R168 B.n309 B.n308 585
R169 B.n311 B.n272 585
R170 B.n314 B.n313 585
R171 B.n315 B.n271 585
R172 B.n317 B.n316 585
R173 B.n319 B.n270 585
R174 B.n322 B.n321 585
R175 B.n323 B.n269 585
R176 B.n325 B.n324 585
R177 B.n327 B.n268 585
R178 B.n330 B.n329 585
R179 B.n331 B.n267 585
R180 B.n333 B.n332 585
R181 B.n335 B.n266 585
R182 B.n338 B.n337 585
R183 B.n339 B.n263 585
R184 B.n342 B.n341 585
R185 B.n344 B.n262 585
R186 B.n347 B.n346 585
R187 B.n348 B.n261 585
R188 B.n350 B.n349 585
R189 B.n352 B.n260 585
R190 B.n355 B.n354 585
R191 B.n356 B.n259 585
R192 B.n361 B.n360 585
R193 B.n363 B.n258 585
R194 B.n366 B.n365 585
R195 B.n367 B.n257 585
R196 B.n369 B.n368 585
R197 B.n371 B.n256 585
R198 B.n374 B.n373 585
R199 B.n375 B.n255 585
R200 B.n377 B.n376 585
R201 B.n379 B.n254 585
R202 B.n382 B.n381 585
R203 B.n383 B.n253 585
R204 B.n385 B.n384 585
R205 B.n387 B.n252 585
R206 B.n390 B.n389 585
R207 B.n391 B.n251 585
R208 B.n393 B.n392 585
R209 B.n395 B.n250 585
R210 B.n398 B.n397 585
R211 B.n399 B.n249 585
R212 B.n401 B.n400 585
R213 B.n403 B.n248 585
R214 B.n406 B.n405 585
R215 B.n407 B.n247 585
R216 B.n409 B.n408 585
R217 B.n411 B.n246 585
R218 B.n414 B.n413 585
R219 B.n415 B.n245 585
R220 B.n417 B.n416 585
R221 B.n419 B.n244 585
R222 B.n422 B.n421 585
R223 B.n423 B.n243 585
R224 B.n428 B.n427 585
R225 B.n427 B.n426 585
R226 B.n429 B.n239 585
R227 B.n239 B.n238 585
R228 B.n431 B.n430 585
R229 B.n432 B.n431 585
R230 B.n233 B.n232 585
R231 B.n234 B.n233 585
R232 B.n441 B.n440 585
R233 B.n440 B.n439 585
R234 B.n442 B.n231 585
R235 B.n438 B.n231 585
R236 B.n444 B.n443 585
R237 B.n445 B.n444 585
R238 B.n226 B.n225 585
R239 B.n227 B.n226 585
R240 B.n453 B.n452 585
R241 B.n452 B.n451 585
R242 B.n454 B.n224 585
R243 B.n224 B.n223 585
R244 B.n456 B.n455 585
R245 B.n457 B.n456 585
R246 B.n218 B.n217 585
R247 B.n219 B.n218 585
R248 B.n466 B.n465 585
R249 B.n465 B.n464 585
R250 B.n467 B.n216 585
R251 B.n216 B.n215 585
R252 B.n469 B.n468 585
R253 B.n470 B.n469 585
R254 B.n2 B.n0 585
R255 B.n4 B.n2 585
R256 B.n3 B.n1 585
R257 B.n529 B.n3 585
R258 B.n527 B.n526 585
R259 B.n528 B.n527 585
R260 B.n525 B.n9 585
R261 B.n9 B.n8 585
R262 B.n524 B.n523 585
R263 B.n523 B.n522 585
R264 B.n11 B.n10 585
R265 B.n521 B.n11 585
R266 B.n519 B.n518 585
R267 B.n520 B.n519 585
R268 B.n517 B.n16 585
R269 B.n16 B.n15 585
R270 B.n516 B.n515 585
R271 B.n515 B.n514 585
R272 B.n18 B.n17 585
R273 B.n513 B.n18 585
R274 B.n511 B.n510 585
R275 B.n512 B.n511 585
R276 B.n509 B.n22 585
R277 B.n25 B.n22 585
R278 B.n508 B.n507 585
R279 B.n507 B.n506 585
R280 B.n24 B.n23 585
R281 B.n505 B.n24 585
R282 B.n503 B.n502 585
R283 B.n504 B.n503 585
R284 B.n501 B.n30 585
R285 B.n30 B.n29 585
R286 B.n500 B.n499 585
R287 B.n499 B.n498 585
R288 B.n532 B.n531 585
R289 B.n531 B.n530 585
R290 B.n427 B.n241 502.111
R291 B.n499 B.n32 502.111
R292 B.n425 B.n243 502.111
R293 B.n496 B.n33 502.111
R294 B.n357 B.t13 393.673
R295 B.n264 B.t9 393.673
R296 B.n73 B.t2 393.673
R297 B.n70 B.t6 393.673
R298 B.n497 B.n68 256.663
R299 B.n497 B.n67 256.663
R300 B.n497 B.n66 256.663
R301 B.n497 B.n65 256.663
R302 B.n497 B.n64 256.663
R303 B.n497 B.n63 256.663
R304 B.n497 B.n62 256.663
R305 B.n497 B.n61 256.663
R306 B.n497 B.n60 256.663
R307 B.n497 B.n59 256.663
R308 B.n497 B.n58 256.663
R309 B.n497 B.n57 256.663
R310 B.n497 B.n56 256.663
R311 B.n497 B.n55 256.663
R312 B.n497 B.n54 256.663
R313 B.n497 B.n53 256.663
R314 B.n497 B.n52 256.663
R315 B.n497 B.n51 256.663
R316 B.n497 B.n50 256.663
R317 B.n497 B.n49 256.663
R318 B.n497 B.n48 256.663
R319 B.n497 B.n47 256.663
R320 B.n497 B.n46 256.663
R321 B.n497 B.n45 256.663
R322 B.n497 B.n44 256.663
R323 B.n497 B.n43 256.663
R324 B.n497 B.n42 256.663
R325 B.n497 B.n41 256.663
R326 B.n497 B.n40 256.663
R327 B.n497 B.n39 256.663
R328 B.n497 B.n38 256.663
R329 B.n497 B.n37 256.663
R330 B.n497 B.n36 256.663
R331 B.n497 B.n35 256.663
R332 B.n497 B.n34 256.663
R333 B.n280 B.n242 256.663
R334 B.n286 B.n242 256.663
R335 B.n288 B.n242 256.663
R336 B.n294 B.n242 256.663
R337 B.n296 B.n242 256.663
R338 B.n302 B.n242 256.663
R339 B.n304 B.n242 256.663
R340 B.n310 B.n242 256.663
R341 B.n312 B.n242 256.663
R342 B.n318 B.n242 256.663
R343 B.n320 B.n242 256.663
R344 B.n326 B.n242 256.663
R345 B.n328 B.n242 256.663
R346 B.n334 B.n242 256.663
R347 B.n336 B.n242 256.663
R348 B.n343 B.n242 256.663
R349 B.n345 B.n242 256.663
R350 B.n351 B.n242 256.663
R351 B.n353 B.n242 256.663
R352 B.n362 B.n242 256.663
R353 B.n364 B.n242 256.663
R354 B.n370 B.n242 256.663
R355 B.n372 B.n242 256.663
R356 B.n378 B.n242 256.663
R357 B.n380 B.n242 256.663
R358 B.n386 B.n242 256.663
R359 B.n388 B.n242 256.663
R360 B.n394 B.n242 256.663
R361 B.n396 B.n242 256.663
R362 B.n402 B.n242 256.663
R363 B.n404 B.n242 256.663
R364 B.n410 B.n242 256.663
R365 B.n412 B.n242 256.663
R366 B.n418 B.n242 256.663
R367 B.n420 B.n242 256.663
R368 B.n427 B.n239 163.367
R369 B.n431 B.n239 163.367
R370 B.n431 B.n233 163.367
R371 B.n440 B.n233 163.367
R372 B.n440 B.n231 163.367
R373 B.n444 B.n231 163.367
R374 B.n444 B.n226 163.367
R375 B.n452 B.n226 163.367
R376 B.n452 B.n224 163.367
R377 B.n456 B.n224 163.367
R378 B.n456 B.n218 163.367
R379 B.n465 B.n218 163.367
R380 B.n465 B.n216 163.367
R381 B.n469 B.n216 163.367
R382 B.n469 B.n2 163.367
R383 B.n531 B.n2 163.367
R384 B.n531 B.n3 163.367
R385 B.n527 B.n3 163.367
R386 B.n527 B.n9 163.367
R387 B.n523 B.n9 163.367
R388 B.n523 B.n11 163.367
R389 B.n519 B.n11 163.367
R390 B.n519 B.n16 163.367
R391 B.n515 B.n16 163.367
R392 B.n515 B.n18 163.367
R393 B.n511 B.n18 163.367
R394 B.n511 B.n22 163.367
R395 B.n507 B.n22 163.367
R396 B.n507 B.n24 163.367
R397 B.n503 B.n24 163.367
R398 B.n503 B.n30 163.367
R399 B.n499 B.n30 163.367
R400 B.n281 B.n279 163.367
R401 B.n285 B.n279 163.367
R402 B.n289 B.n287 163.367
R403 B.n293 B.n277 163.367
R404 B.n297 B.n295 163.367
R405 B.n301 B.n275 163.367
R406 B.n305 B.n303 163.367
R407 B.n309 B.n273 163.367
R408 B.n313 B.n311 163.367
R409 B.n317 B.n271 163.367
R410 B.n321 B.n319 163.367
R411 B.n325 B.n269 163.367
R412 B.n329 B.n327 163.367
R413 B.n333 B.n267 163.367
R414 B.n337 B.n335 163.367
R415 B.n342 B.n263 163.367
R416 B.n346 B.n344 163.367
R417 B.n350 B.n261 163.367
R418 B.n354 B.n352 163.367
R419 B.n361 B.n259 163.367
R420 B.n365 B.n363 163.367
R421 B.n369 B.n257 163.367
R422 B.n373 B.n371 163.367
R423 B.n377 B.n255 163.367
R424 B.n381 B.n379 163.367
R425 B.n385 B.n253 163.367
R426 B.n389 B.n387 163.367
R427 B.n393 B.n251 163.367
R428 B.n397 B.n395 163.367
R429 B.n401 B.n249 163.367
R430 B.n405 B.n403 163.367
R431 B.n409 B.n247 163.367
R432 B.n413 B.n411 163.367
R433 B.n417 B.n245 163.367
R434 B.n421 B.n419 163.367
R435 B.n425 B.n237 163.367
R436 B.n433 B.n237 163.367
R437 B.n433 B.n235 163.367
R438 B.n437 B.n235 163.367
R439 B.n437 B.n230 163.367
R440 B.n446 B.n230 163.367
R441 B.n446 B.n228 163.367
R442 B.n450 B.n228 163.367
R443 B.n450 B.n222 163.367
R444 B.n458 B.n222 163.367
R445 B.n458 B.n220 163.367
R446 B.n463 B.n220 163.367
R447 B.n463 B.n214 163.367
R448 B.n471 B.n214 163.367
R449 B.n472 B.n471 163.367
R450 B.n472 B.n5 163.367
R451 B.n6 B.n5 163.367
R452 B.n7 B.n6 163.367
R453 B.n477 B.n7 163.367
R454 B.n477 B.n12 163.367
R455 B.n13 B.n12 163.367
R456 B.n14 B.n13 163.367
R457 B.n482 B.n14 163.367
R458 B.n482 B.n19 163.367
R459 B.n20 B.n19 163.367
R460 B.n21 B.n20 163.367
R461 B.n487 B.n21 163.367
R462 B.n487 B.n26 163.367
R463 B.n27 B.n26 163.367
R464 B.n28 B.n27 163.367
R465 B.n492 B.n28 163.367
R466 B.n492 B.n33 163.367
R467 B.n77 B.n76 163.367
R468 B.n81 B.n80 163.367
R469 B.n85 B.n84 163.367
R470 B.n89 B.n88 163.367
R471 B.n93 B.n92 163.367
R472 B.n97 B.n96 163.367
R473 B.n101 B.n100 163.367
R474 B.n105 B.n104 163.367
R475 B.n109 B.n108 163.367
R476 B.n113 B.n112 163.367
R477 B.n117 B.n116 163.367
R478 B.n121 B.n120 163.367
R479 B.n125 B.n124 163.367
R480 B.n129 B.n128 163.367
R481 B.n133 B.n132 163.367
R482 B.n138 B.n137 163.367
R483 B.n142 B.n141 163.367
R484 B.n146 B.n145 163.367
R485 B.n150 B.n149 163.367
R486 B.n154 B.n153 163.367
R487 B.n158 B.n157 163.367
R488 B.n162 B.n161 163.367
R489 B.n166 B.n165 163.367
R490 B.n170 B.n169 163.367
R491 B.n174 B.n173 163.367
R492 B.n178 B.n177 163.367
R493 B.n182 B.n181 163.367
R494 B.n186 B.n185 163.367
R495 B.n190 B.n189 163.367
R496 B.n194 B.n193 163.367
R497 B.n198 B.n197 163.367
R498 B.n202 B.n201 163.367
R499 B.n206 B.n205 163.367
R500 B.n210 B.n209 163.367
R501 B.n496 B.n69 163.367
R502 B.n426 B.n242 109.879
R503 B.n498 B.n497 109.879
R504 B.n357 B.t15 96.277
R505 B.n70 B.t7 96.277
R506 B.n264 B.t12 96.2672
R507 B.n73 B.t4 96.2672
R508 B.n280 B.n241 71.676
R509 B.n286 B.n285 71.676
R510 B.n289 B.n288 71.676
R511 B.n294 B.n293 71.676
R512 B.n297 B.n296 71.676
R513 B.n302 B.n301 71.676
R514 B.n305 B.n304 71.676
R515 B.n310 B.n309 71.676
R516 B.n313 B.n312 71.676
R517 B.n318 B.n317 71.676
R518 B.n321 B.n320 71.676
R519 B.n326 B.n325 71.676
R520 B.n329 B.n328 71.676
R521 B.n334 B.n333 71.676
R522 B.n337 B.n336 71.676
R523 B.n343 B.n342 71.676
R524 B.n346 B.n345 71.676
R525 B.n351 B.n350 71.676
R526 B.n354 B.n353 71.676
R527 B.n362 B.n361 71.676
R528 B.n365 B.n364 71.676
R529 B.n370 B.n369 71.676
R530 B.n373 B.n372 71.676
R531 B.n378 B.n377 71.676
R532 B.n381 B.n380 71.676
R533 B.n386 B.n385 71.676
R534 B.n389 B.n388 71.676
R535 B.n394 B.n393 71.676
R536 B.n397 B.n396 71.676
R537 B.n402 B.n401 71.676
R538 B.n405 B.n404 71.676
R539 B.n410 B.n409 71.676
R540 B.n413 B.n412 71.676
R541 B.n418 B.n417 71.676
R542 B.n421 B.n420 71.676
R543 B.n34 B.n32 71.676
R544 B.n77 B.n35 71.676
R545 B.n81 B.n36 71.676
R546 B.n85 B.n37 71.676
R547 B.n89 B.n38 71.676
R548 B.n93 B.n39 71.676
R549 B.n97 B.n40 71.676
R550 B.n101 B.n41 71.676
R551 B.n105 B.n42 71.676
R552 B.n109 B.n43 71.676
R553 B.n113 B.n44 71.676
R554 B.n117 B.n45 71.676
R555 B.n121 B.n46 71.676
R556 B.n125 B.n47 71.676
R557 B.n129 B.n48 71.676
R558 B.n133 B.n49 71.676
R559 B.n138 B.n50 71.676
R560 B.n142 B.n51 71.676
R561 B.n146 B.n52 71.676
R562 B.n150 B.n53 71.676
R563 B.n154 B.n54 71.676
R564 B.n158 B.n55 71.676
R565 B.n162 B.n56 71.676
R566 B.n166 B.n57 71.676
R567 B.n170 B.n58 71.676
R568 B.n174 B.n59 71.676
R569 B.n178 B.n60 71.676
R570 B.n182 B.n61 71.676
R571 B.n186 B.n62 71.676
R572 B.n190 B.n63 71.676
R573 B.n194 B.n64 71.676
R574 B.n198 B.n65 71.676
R575 B.n202 B.n66 71.676
R576 B.n206 B.n67 71.676
R577 B.n210 B.n68 71.676
R578 B.n69 B.n68 71.676
R579 B.n209 B.n67 71.676
R580 B.n205 B.n66 71.676
R581 B.n201 B.n65 71.676
R582 B.n197 B.n64 71.676
R583 B.n193 B.n63 71.676
R584 B.n189 B.n62 71.676
R585 B.n185 B.n61 71.676
R586 B.n181 B.n60 71.676
R587 B.n177 B.n59 71.676
R588 B.n173 B.n58 71.676
R589 B.n169 B.n57 71.676
R590 B.n165 B.n56 71.676
R591 B.n161 B.n55 71.676
R592 B.n157 B.n54 71.676
R593 B.n153 B.n53 71.676
R594 B.n149 B.n52 71.676
R595 B.n145 B.n51 71.676
R596 B.n141 B.n50 71.676
R597 B.n137 B.n49 71.676
R598 B.n132 B.n48 71.676
R599 B.n128 B.n47 71.676
R600 B.n124 B.n46 71.676
R601 B.n120 B.n45 71.676
R602 B.n116 B.n44 71.676
R603 B.n112 B.n43 71.676
R604 B.n108 B.n42 71.676
R605 B.n104 B.n41 71.676
R606 B.n100 B.n40 71.676
R607 B.n96 B.n39 71.676
R608 B.n92 B.n38 71.676
R609 B.n88 B.n37 71.676
R610 B.n84 B.n36 71.676
R611 B.n80 B.n35 71.676
R612 B.n76 B.n34 71.676
R613 B.n281 B.n280 71.676
R614 B.n287 B.n286 71.676
R615 B.n288 B.n277 71.676
R616 B.n295 B.n294 71.676
R617 B.n296 B.n275 71.676
R618 B.n303 B.n302 71.676
R619 B.n304 B.n273 71.676
R620 B.n311 B.n310 71.676
R621 B.n312 B.n271 71.676
R622 B.n319 B.n318 71.676
R623 B.n320 B.n269 71.676
R624 B.n327 B.n326 71.676
R625 B.n328 B.n267 71.676
R626 B.n335 B.n334 71.676
R627 B.n336 B.n263 71.676
R628 B.n344 B.n343 71.676
R629 B.n345 B.n261 71.676
R630 B.n352 B.n351 71.676
R631 B.n353 B.n259 71.676
R632 B.n363 B.n362 71.676
R633 B.n364 B.n257 71.676
R634 B.n371 B.n370 71.676
R635 B.n372 B.n255 71.676
R636 B.n379 B.n378 71.676
R637 B.n380 B.n253 71.676
R638 B.n387 B.n386 71.676
R639 B.n388 B.n251 71.676
R640 B.n395 B.n394 71.676
R641 B.n396 B.n249 71.676
R642 B.n403 B.n402 71.676
R643 B.n404 B.n247 71.676
R644 B.n411 B.n410 71.676
R645 B.n412 B.n245 71.676
R646 B.n419 B.n418 71.676
R647 B.n420 B.n243 71.676
R648 B.n358 B.t14 69.7073
R649 B.n71 B.t8 69.7073
R650 B.n265 B.t11 69.6975
R651 B.n74 B.t5 69.6975
R652 B.n359 B.n358 59.5399
R653 B.n340 B.n265 59.5399
R654 B.n135 B.n74 59.5399
R655 B.n72 B.n71 59.5399
R656 B.n426 B.n238 55.3464
R657 B.n432 B.n238 55.3464
R658 B.n432 B.n234 55.3464
R659 B.n439 B.n234 55.3464
R660 B.n439 B.n438 55.3464
R661 B.n445 B.n227 55.3464
R662 B.n451 B.n227 55.3464
R663 B.n451 B.n223 55.3464
R664 B.n457 B.n223 55.3464
R665 B.n457 B.n219 55.3464
R666 B.n464 B.n219 55.3464
R667 B.n470 B.n215 55.3464
R668 B.n470 B.n4 55.3464
R669 B.n530 B.n4 55.3464
R670 B.n530 B.n529 55.3464
R671 B.n529 B.n528 55.3464
R672 B.n528 B.n8 55.3464
R673 B.n522 B.n521 55.3464
R674 B.n521 B.n520 55.3464
R675 B.n520 B.n15 55.3464
R676 B.n514 B.n15 55.3464
R677 B.n514 B.n513 55.3464
R678 B.n513 B.n512 55.3464
R679 B.n506 B.n25 55.3464
R680 B.n506 B.n505 55.3464
R681 B.n505 B.n504 55.3464
R682 B.n504 B.n29 55.3464
R683 B.n498 B.n29 55.3464
R684 B.n445 B.t10 47.2073
R685 B.n512 B.t3 47.2073
R686 B.t0 B.n215 34.1847
R687 B.t1 B.n8 34.1847
R688 B.n500 B.n31 32.6249
R689 B.n495 B.n494 32.6249
R690 B.n424 B.n423 32.6249
R691 B.n428 B.n240 32.6249
R692 B.n358 B.n357 26.5702
R693 B.n265 B.n264 26.5702
R694 B.n74 B.n73 26.5702
R695 B.n71 B.n70 26.5702
R696 B.n464 B.t0 21.1622
R697 B.n522 B.t1 21.1622
R698 B B.n532 18.0485
R699 B.n75 B.n31 10.6151
R700 B.n78 B.n75 10.6151
R701 B.n79 B.n78 10.6151
R702 B.n82 B.n79 10.6151
R703 B.n83 B.n82 10.6151
R704 B.n86 B.n83 10.6151
R705 B.n87 B.n86 10.6151
R706 B.n90 B.n87 10.6151
R707 B.n91 B.n90 10.6151
R708 B.n94 B.n91 10.6151
R709 B.n95 B.n94 10.6151
R710 B.n98 B.n95 10.6151
R711 B.n99 B.n98 10.6151
R712 B.n102 B.n99 10.6151
R713 B.n103 B.n102 10.6151
R714 B.n106 B.n103 10.6151
R715 B.n107 B.n106 10.6151
R716 B.n110 B.n107 10.6151
R717 B.n111 B.n110 10.6151
R718 B.n114 B.n111 10.6151
R719 B.n115 B.n114 10.6151
R720 B.n118 B.n115 10.6151
R721 B.n119 B.n118 10.6151
R722 B.n122 B.n119 10.6151
R723 B.n123 B.n122 10.6151
R724 B.n126 B.n123 10.6151
R725 B.n127 B.n126 10.6151
R726 B.n130 B.n127 10.6151
R727 B.n131 B.n130 10.6151
R728 B.n134 B.n131 10.6151
R729 B.n139 B.n136 10.6151
R730 B.n140 B.n139 10.6151
R731 B.n143 B.n140 10.6151
R732 B.n144 B.n143 10.6151
R733 B.n147 B.n144 10.6151
R734 B.n148 B.n147 10.6151
R735 B.n151 B.n148 10.6151
R736 B.n152 B.n151 10.6151
R737 B.n156 B.n155 10.6151
R738 B.n159 B.n156 10.6151
R739 B.n160 B.n159 10.6151
R740 B.n163 B.n160 10.6151
R741 B.n164 B.n163 10.6151
R742 B.n167 B.n164 10.6151
R743 B.n168 B.n167 10.6151
R744 B.n171 B.n168 10.6151
R745 B.n172 B.n171 10.6151
R746 B.n175 B.n172 10.6151
R747 B.n176 B.n175 10.6151
R748 B.n179 B.n176 10.6151
R749 B.n180 B.n179 10.6151
R750 B.n183 B.n180 10.6151
R751 B.n184 B.n183 10.6151
R752 B.n187 B.n184 10.6151
R753 B.n188 B.n187 10.6151
R754 B.n191 B.n188 10.6151
R755 B.n192 B.n191 10.6151
R756 B.n195 B.n192 10.6151
R757 B.n196 B.n195 10.6151
R758 B.n199 B.n196 10.6151
R759 B.n200 B.n199 10.6151
R760 B.n203 B.n200 10.6151
R761 B.n204 B.n203 10.6151
R762 B.n207 B.n204 10.6151
R763 B.n208 B.n207 10.6151
R764 B.n211 B.n208 10.6151
R765 B.n212 B.n211 10.6151
R766 B.n495 B.n212 10.6151
R767 B.n424 B.n236 10.6151
R768 B.n434 B.n236 10.6151
R769 B.n435 B.n434 10.6151
R770 B.n436 B.n435 10.6151
R771 B.n436 B.n229 10.6151
R772 B.n447 B.n229 10.6151
R773 B.n448 B.n447 10.6151
R774 B.n449 B.n448 10.6151
R775 B.n449 B.n221 10.6151
R776 B.n459 B.n221 10.6151
R777 B.n460 B.n459 10.6151
R778 B.n462 B.n460 10.6151
R779 B.n462 B.n461 10.6151
R780 B.n461 B.n213 10.6151
R781 B.n473 B.n213 10.6151
R782 B.n474 B.n473 10.6151
R783 B.n475 B.n474 10.6151
R784 B.n476 B.n475 10.6151
R785 B.n478 B.n476 10.6151
R786 B.n479 B.n478 10.6151
R787 B.n480 B.n479 10.6151
R788 B.n481 B.n480 10.6151
R789 B.n483 B.n481 10.6151
R790 B.n484 B.n483 10.6151
R791 B.n485 B.n484 10.6151
R792 B.n486 B.n485 10.6151
R793 B.n488 B.n486 10.6151
R794 B.n489 B.n488 10.6151
R795 B.n490 B.n489 10.6151
R796 B.n491 B.n490 10.6151
R797 B.n493 B.n491 10.6151
R798 B.n494 B.n493 10.6151
R799 B.n282 B.n240 10.6151
R800 B.n283 B.n282 10.6151
R801 B.n284 B.n283 10.6151
R802 B.n284 B.n278 10.6151
R803 B.n290 B.n278 10.6151
R804 B.n291 B.n290 10.6151
R805 B.n292 B.n291 10.6151
R806 B.n292 B.n276 10.6151
R807 B.n298 B.n276 10.6151
R808 B.n299 B.n298 10.6151
R809 B.n300 B.n299 10.6151
R810 B.n300 B.n274 10.6151
R811 B.n306 B.n274 10.6151
R812 B.n307 B.n306 10.6151
R813 B.n308 B.n307 10.6151
R814 B.n308 B.n272 10.6151
R815 B.n314 B.n272 10.6151
R816 B.n315 B.n314 10.6151
R817 B.n316 B.n315 10.6151
R818 B.n316 B.n270 10.6151
R819 B.n322 B.n270 10.6151
R820 B.n323 B.n322 10.6151
R821 B.n324 B.n323 10.6151
R822 B.n324 B.n268 10.6151
R823 B.n330 B.n268 10.6151
R824 B.n331 B.n330 10.6151
R825 B.n332 B.n331 10.6151
R826 B.n332 B.n266 10.6151
R827 B.n338 B.n266 10.6151
R828 B.n339 B.n338 10.6151
R829 B.n341 B.n262 10.6151
R830 B.n347 B.n262 10.6151
R831 B.n348 B.n347 10.6151
R832 B.n349 B.n348 10.6151
R833 B.n349 B.n260 10.6151
R834 B.n355 B.n260 10.6151
R835 B.n356 B.n355 10.6151
R836 B.n360 B.n356 10.6151
R837 B.n366 B.n258 10.6151
R838 B.n367 B.n366 10.6151
R839 B.n368 B.n367 10.6151
R840 B.n368 B.n256 10.6151
R841 B.n374 B.n256 10.6151
R842 B.n375 B.n374 10.6151
R843 B.n376 B.n375 10.6151
R844 B.n376 B.n254 10.6151
R845 B.n382 B.n254 10.6151
R846 B.n383 B.n382 10.6151
R847 B.n384 B.n383 10.6151
R848 B.n384 B.n252 10.6151
R849 B.n390 B.n252 10.6151
R850 B.n391 B.n390 10.6151
R851 B.n392 B.n391 10.6151
R852 B.n392 B.n250 10.6151
R853 B.n398 B.n250 10.6151
R854 B.n399 B.n398 10.6151
R855 B.n400 B.n399 10.6151
R856 B.n400 B.n248 10.6151
R857 B.n406 B.n248 10.6151
R858 B.n407 B.n406 10.6151
R859 B.n408 B.n407 10.6151
R860 B.n408 B.n246 10.6151
R861 B.n414 B.n246 10.6151
R862 B.n415 B.n414 10.6151
R863 B.n416 B.n415 10.6151
R864 B.n416 B.n244 10.6151
R865 B.n422 B.n244 10.6151
R866 B.n423 B.n422 10.6151
R867 B.n429 B.n428 10.6151
R868 B.n430 B.n429 10.6151
R869 B.n430 B.n232 10.6151
R870 B.n441 B.n232 10.6151
R871 B.n442 B.n441 10.6151
R872 B.n443 B.n442 10.6151
R873 B.n443 B.n225 10.6151
R874 B.n453 B.n225 10.6151
R875 B.n454 B.n453 10.6151
R876 B.n455 B.n454 10.6151
R877 B.n455 B.n217 10.6151
R878 B.n466 B.n217 10.6151
R879 B.n467 B.n466 10.6151
R880 B.n468 B.n467 10.6151
R881 B.n468 B.n0 10.6151
R882 B.n526 B.n1 10.6151
R883 B.n526 B.n525 10.6151
R884 B.n525 B.n524 10.6151
R885 B.n524 B.n10 10.6151
R886 B.n518 B.n10 10.6151
R887 B.n518 B.n517 10.6151
R888 B.n517 B.n516 10.6151
R889 B.n516 B.n17 10.6151
R890 B.n510 B.n17 10.6151
R891 B.n510 B.n509 10.6151
R892 B.n509 B.n508 10.6151
R893 B.n508 B.n23 10.6151
R894 B.n502 B.n23 10.6151
R895 B.n502 B.n501 10.6151
R896 B.n501 B.n500 10.6151
R897 B.n438 B.t10 8.1396
R898 B.n25 B.t3 8.1396
R899 B.n136 B.n135 7.18099
R900 B.n152 B.n72 7.18099
R901 B.n341 B.n340 7.18099
R902 B.n360 B.n359 7.18099
R903 B.n135 B.n134 3.43465
R904 B.n155 B.n72 3.43465
R905 B.n340 B.n339 3.43465
R906 B.n359 B.n258 3.43465
R907 B.n532 B.n0 2.81026
R908 B.n532 B.n1 2.81026
R909 VP.n0 VP.t0 427.69
R910 VP.n0 VP.t1 390.019
R911 VP VP.n0 0.0516364
R912 VDD1 VDD1.t0 101.213
R913 VDD1 VDD1.t1 67.6214
C0 VDD2 VTAIL 4.07443f
C1 VDD2 VN 1.62438f
C2 VDD1 VTAIL 4.03538f
C3 VDD1 VN 0.14841f
C4 VN VTAIL 1.33097f
C5 VP VDD2 0.2683f
C6 VP VDD1 1.74156f
C7 VDD2 VDD1 0.495395f
C8 VP VTAIL 1.34536f
C9 VP VN 4.01751f
C10 VDD2 B 3.181767f
C11 VDD1 B 4.95749f
C12 VTAIL B 5.083787f
C13 VN B 6.51986f
C14 VP B 4.17336f
C15 VDD1.t1 B 1.02474f
C16 VDD1.t0 B 1.29596f
C17 VP.t0 B 0.927884f
C18 VP.t1 B 0.825663f
C19 VP.n0 B 2.23047f
C20 VDD2.t0 B 1.32873f
C21 VDD2.t1 B 1.06347f
C22 VDD2.n0 B 1.66225f
C23 VTAIL.t0 B 1.09508f
C24 VTAIL.n0 B 0.948178f
C25 VTAIL.t2 B 1.09509f
C26 VTAIL.n1 B 0.960417f
C27 VTAIL.t1 B 1.09508f
C28 VTAIL.n2 B 0.899412f
C29 VTAIL.t3 B 1.09508f
C30 VTAIL.n3 B 0.856882f
C31 VN.t1 B 0.817462f
C32 VN.t0 B 0.921236f
.ends

