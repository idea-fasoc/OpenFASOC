* NGSPICE file created from diff_pair_sample_0402.ext - technology: sky130A

.subckt diff_pair_sample_0402 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0.50655 ps=3.4 w=3.07 l=1.13
X1 VTAIL.t6 VN.t1 VDD2.t2 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0.50655 ps=3.4 w=3.07 l=1.13
X2 B.t11 B.t9 B.t10 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.13
X3 VTAIL.t1 VP.t0 VDD1.t3 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0.50655 ps=3.4 w=3.07 l=1.13
X4 VDD1.t2 VP.t1 VTAIL.t3 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=0.50655 pd=3.4 as=1.1973 ps=6.92 w=3.07 l=1.13
X5 B.t8 B.t6 B.t7 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.13
X6 VDD2.t0 VN.t2 VTAIL.t5 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=0.50655 pd=3.4 as=1.1973 ps=6.92 w=3.07 l=1.13
X7 VDD2.t1 VN.t3 VTAIL.t4 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=0.50655 pd=3.4 as=1.1973 ps=6.92 w=3.07 l=1.13
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0.50655 ps=3.4 w=3.07 l=1.13
X9 B.t5 B.t3 B.t4 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.13
X10 B.t2 B.t0 B.t1 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.13
X11 VDD1.t0 VP.t3 VTAIL.t2 w_n1846_n1582# sky130_fd_pr__pfet_01v8 ad=0.50655 pd=3.4 as=1.1973 ps=6.92 w=3.07 l=1.13
R0 VN.n0 VN.t0 119.059
R1 VN.n1 VN.t2 119.059
R2 VN.n1 VN.t1 118.972
R3 VN.n0 VN.t3 118.972
R4 VN VN.n1 66.6751
R5 VN VN.n0 31.2622
R6 VDD2.n2 VDD2.n0 157.018
R7 VDD2.n2 VDD2.n1 126.882
R8 VDD2.n1 VDD2.t2 10.5884
R9 VDD2.n1 VDD2.t0 10.5884
R10 VDD2.n0 VDD2.t3 10.5884
R11 VDD2.n0 VDD2.t1 10.5884
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n122 VTAIL.n112 756.745
R14 VTAIL.n10 VTAIL.n0 756.745
R15 VTAIL.n26 VTAIL.n16 756.745
R16 VTAIL.n42 VTAIL.n32 756.745
R17 VTAIL.n106 VTAIL.n96 756.745
R18 VTAIL.n90 VTAIL.n80 756.745
R19 VTAIL.n74 VTAIL.n64 756.745
R20 VTAIL.n58 VTAIL.n48 756.745
R21 VTAIL.n116 VTAIL.n115 585
R22 VTAIL.n121 VTAIL.n120 585
R23 VTAIL.n123 VTAIL.n122 585
R24 VTAIL.n4 VTAIL.n3 585
R25 VTAIL.n9 VTAIL.n8 585
R26 VTAIL.n11 VTAIL.n10 585
R27 VTAIL.n20 VTAIL.n19 585
R28 VTAIL.n25 VTAIL.n24 585
R29 VTAIL.n27 VTAIL.n26 585
R30 VTAIL.n36 VTAIL.n35 585
R31 VTAIL.n41 VTAIL.n40 585
R32 VTAIL.n43 VTAIL.n42 585
R33 VTAIL.n107 VTAIL.n106 585
R34 VTAIL.n105 VTAIL.n104 585
R35 VTAIL.n100 VTAIL.n99 585
R36 VTAIL.n91 VTAIL.n90 585
R37 VTAIL.n89 VTAIL.n88 585
R38 VTAIL.n84 VTAIL.n83 585
R39 VTAIL.n75 VTAIL.n74 585
R40 VTAIL.n73 VTAIL.n72 585
R41 VTAIL.n68 VTAIL.n67 585
R42 VTAIL.n59 VTAIL.n58 585
R43 VTAIL.n57 VTAIL.n56 585
R44 VTAIL.n52 VTAIL.n51 585
R45 VTAIL.n117 VTAIL.t4 336.901
R46 VTAIL.n5 VTAIL.t7 336.901
R47 VTAIL.n21 VTAIL.t3 336.901
R48 VTAIL.n37 VTAIL.t0 336.901
R49 VTAIL.n101 VTAIL.t2 336.901
R50 VTAIL.n85 VTAIL.t1 336.901
R51 VTAIL.n69 VTAIL.t5 336.901
R52 VTAIL.n53 VTAIL.t6 336.901
R53 VTAIL.n121 VTAIL.n115 171.744
R54 VTAIL.n122 VTAIL.n121 171.744
R55 VTAIL.n9 VTAIL.n3 171.744
R56 VTAIL.n10 VTAIL.n9 171.744
R57 VTAIL.n25 VTAIL.n19 171.744
R58 VTAIL.n26 VTAIL.n25 171.744
R59 VTAIL.n41 VTAIL.n35 171.744
R60 VTAIL.n42 VTAIL.n41 171.744
R61 VTAIL.n106 VTAIL.n105 171.744
R62 VTAIL.n105 VTAIL.n99 171.744
R63 VTAIL.n90 VTAIL.n89 171.744
R64 VTAIL.n89 VTAIL.n83 171.744
R65 VTAIL.n74 VTAIL.n73 171.744
R66 VTAIL.n73 VTAIL.n67 171.744
R67 VTAIL.n58 VTAIL.n57 171.744
R68 VTAIL.n57 VTAIL.n51 171.744
R69 VTAIL.t4 VTAIL.n115 85.8723
R70 VTAIL.t7 VTAIL.n3 85.8723
R71 VTAIL.t3 VTAIL.n19 85.8723
R72 VTAIL.t0 VTAIL.n35 85.8723
R73 VTAIL.t2 VTAIL.n99 85.8723
R74 VTAIL.t1 VTAIL.n83 85.8723
R75 VTAIL.t5 VTAIL.n67 85.8723
R76 VTAIL.t6 VTAIL.n51 85.8723
R77 VTAIL.n127 VTAIL.n126 31.2157
R78 VTAIL.n15 VTAIL.n14 31.2157
R79 VTAIL.n31 VTAIL.n30 31.2157
R80 VTAIL.n47 VTAIL.n46 31.2157
R81 VTAIL.n111 VTAIL.n110 31.2157
R82 VTAIL.n95 VTAIL.n94 31.2157
R83 VTAIL.n79 VTAIL.n78 31.2157
R84 VTAIL.n63 VTAIL.n62 31.2157
R85 VTAIL.n127 VTAIL.n111 16.2721
R86 VTAIL.n63 VTAIL.n47 16.2721
R87 VTAIL.n117 VTAIL.n116 16.193
R88 VTAIL.n5 VTAIL.n4 16.193
R89 VTAIL.n21 VTAIL.n20 16.193
R90 VTAIL.n37 VTAIL.n36 16.193
R91 VTAIL.n101 VTAIL.n100 16.193
R92 VTAIL.n85 VTAIL.n84 16.193
R93 VTAIL.n69 VTAIL.n68 16.193
R94 VTAIL.n53 VTAIL.n52 16.193
R95 VTAIL.n120 VTAIL.n119 12.8005
R96 VTAIL.n8 VTAIL.n7 12.8005
R97 VTAIL.n24 VTAIL.n23 12.8005
R98 VTAIL.n40 VTAIL.n39 12.8005
R99 VTAIL.n104 VTAIL.n103 12.8005
R100 VTAIL.n88 VTAIL.n87 12.8005
R101 VTAIL.n72 VTAIL.n71 12.8005
R102 VTAIL.n56 VTAIL.n55 12.8005
R103 VTAIL.n123 VTAIL.n114 12.0247
R104 VTAIL.n11 VTAIL.n2 12.0247
R105 VTAIL.n27 VTAIL.n18 12.0247
R106 VTAIL.n43 VTAIL.n34 12.0247
R107 VTAIL.n107 VTAIL.n98 12.0247
R108 VTAIL.n91 VTAIL.n82 12.0247
R109 VTAIL.n75 VTAIL.n66 12.0247
R110 VTAIL.n59 VTAIL.n50 12.0247
R111 VTAIL.n124 VTAIL.n112 11.249
R112 VTAIL.n12 VTAIL.n0 11.249
R113 VTAIL.n28 VTAIL.n16 11.249
R114 VTAIL.n44 VTAIL.n32 11.249
R115 VTAIL.n108 VTAIL.n96 11.249
R116 VTAIL.n92 VTAIL.n80 11.249
R117 VTAIL.n76 VTAIL.n64 11.249
R118 VTAIL.n60 VTAIL.n48 11.249
R119 VTAIL.n126 VTAIL.n125 9.45567
R120 VTAIL.n14 VTAIL.n13 9.45567
R121 VTAIL.n30 VTAIL.n29 9.45567
R122 VTAIL.n46 VTAIL.n45 9.45567
R123 VTAIL.n110 VTAIL.n109 9.45567
R124 VTAIL.n94 VTAIL.n93 9.45567
R125 VTAIL.n78 VTAIL.n77 9.45567
R126 VTAIL.n62 VTAIL.n61 9.45567
R127 VTAIL.n125 VTAIL.n124 9.3005
R128 VTAIL.n114 VTAIL.n113 9.3005
R129 VTAIL.n119 VTAIL.n118 9.3005
R130 VTAIL.n13 VTAIL.n12 9.3005
R131 VTAIL.n2 VTAIL.n1 9.3005
R132 VTAIL.n7 VTAIL.n6 9.3005
R133 VTAIL.n29 VTAIL.n28 9.3005
R134 VTAIL.n18 VTAIL.n17 9.3005
R135 VTAIL.n23 VTAIL.n22 9.3005
R136 VTAIL.n45 VTAIL.n44 9.3005
R137 VTAIL.n34 VTAIL.n33 9.3005
R138 VTAIL.n39 VTAIL.n38 9.3005
R139 VTAIL.n109 VTAIL.n108 9.3005
R140 VTAIL.n98 VTAIL.n97 9.3005
R141 VTAIL.n103 VTAIL.n102 9.3005
R142 VTAIL.n93 VTAIL.n92 9.3005
R143 VTAIL.n82 VTAIL.n81 9.3005
R144 VTAIL.n87 VTAIL.n86 9.3005
R145 VTAIL.n77 VTAIL.n76 9.3005
R146 VTAIL.n66 VTAIL.n65 9.3005
R147 VTAIL.n71 VTAIL.n70 9.3005
R148 VTAIL.n61 VTAIL.n60 9.3005
R149 VTAIL.n50 VTAIL.n49 9.3005
R150 VTAIL.n55 VTAIL.n54 9.3005
R151 VTAIL.n102 VTAIL.n101 3.91276
R152 VTAIL.n86 VTAIL.n85 3.91276
R153 VTAIL.n70 VTAIL.n69 3.91276
R154 VTAIL.n54 VTAIL.n53 3.91276
R155 VTAIL.n118 VTAIL.n117 3.91276
R156 VTAIL.n6 VTAIL.n5 3.91276
R157 VTAIL.n22 VTAIL.n21 3.91276
R158 VTAIL.n38 VTAIL.n37 3.91276
R159 VTAIL.n126 VTAIL.n112 2.71565
R160 VTAIL.n14 VTAIL.n0 2.71565
R161 VTAIL.n30 VTAIL.n16 2.71565
R162 VTAIL.n46 VTAIL.n32 2.71565
R163 VTAIL.n110 VTAIL.n96 2.71565
R164 VTAIL.n94 VTAIL.n80 2.71565
R165 VTAIL.n78 VTAIL.n64 2.71565
R166 VTAIL.n62 VTAIL.n48 2.71565
R167 VTAIL.n124 VTAIL.n123 1.93989
R168 VTAIL.n12 VTAIL.n11 1.93989
R169 VTAIL.n28 VTAIL.n27 1.93989
R170 VTAIL.n44 VTAIL.n43 1.93989
R171 VTAIL.n108 VTAIL.n107 1.93989
R172 VTAIL.n92 VTAIL.n91 1.93989
R173 VTAIL.n76 VTAIL.n75 1.93989
R174 VTAIL.n60 VTAIL.n59 1.93989
R175 VTAIL.n79 VTAIL.n63 1.25912
R176 VTAIL.n111 VTAIL.n95 1.25912
R177 VTAIL.n47 VTAIL.n31 1.25912
R178 VTAIL.n120 VTAIL.n114 1.16414
R179 VTAIL.n8 VTAIL.n2 1.16414
R180 VTAIL.n24 VTAIL.n18 1.16414
R181 VTAIL.n40 VTAIL.n34 1.16414
R182 VTAIL.n104 VTAIL.n98 1.16414
R183 VTAIL.n88 VTAIL.n82 1.16414
R184 VTAIL.n72 VTAIL.n66 1.16414
R185 VTAIL.n56 VTAIL.n50 1.16414
R186 VTAIL VTAIL.n15 0.688
R187 VTAIL VTAIL.n127 0.571621
R188 VTAIL.n95 VTAIL.n79 0.470328
R189 VTAIL.n31 VTAIL.n15 0.470328
R190 VTAIL.n119 VTAIL.n116 0.388379
R191 VTAIL.n7 VTAIL.n4 0.388379
R192 VTAIL.n23 VTAIL.n20 0.388379
R193 VTAIL.n39 VTAIL.n36 0.388379
R194 VTAIL.n103 VTAIL.n100 0.388379
R195 VTAIL.n87 VTAIL.n84 0.388379
R196 VTAIL.n71 VTAIL.n68 0.388379
R197 VTAIL.n55 VTAIL.n52 0.388379
R198 VTAIL.n118 VTAIL.n113 0.155672
R199 VTAIL.n125 VTAIL.n113 0.155672
R200 VTAIL.n6 VTAIL.n1 0.155672
R201 VTAIL.n13 VTAIL.n1 0.155672
R202 VTAIL.n22 VTAIL.n17 0.155672
R203 VTAIL.n29 VTAIL.n17 0.155672
R204 VTAIL.n38 VTAIL.n33 0.155672
R205 VTAIL.n45 VTAIL.n33 0.155672
R206 VTAIL.n109 VTAIL.n97 0.155672
R207 VTAIL.n102 VTAIL.n97 0.155672
R208 VTAIL.n93 VTAIL.n81 0.155672
R209 VTAIL.n86 VTAIL.n81 0.155672
R210 VTAIL.n77 VTAIL.n65 0.155672
R211 VTAIL.n70 VTAIL.n65 0.155672
R212 VTAIL.n61 VTAIL.n49 0.155672
R213 VTAIL.n54 VTAIL.n49 0.155672
R214 B.n250 B.n249 585
R215 B.n251 B.n36 585
R216 B.n253 B.n252 585
R217 B.n254 B.n35 585
R218 B.n256 B.n255 585
R219 B.n257 B.n34 585
R220 B.n259 B.n258 585
R221 B.n260 B.n33 585
R222 B.n262 B.n261 585
R223 B.n263 B.n32 585
R224 B.n265 B.n264 585
R225 B.n266 B.n31 585
R226 B.n268 B.n267 585
R227 B.n269 B.n30 585
R228 B.n271 B.n270 585
R229 B.n273 B.n27 585
R230 B.n275 B.n274 585
R231 B.n276 B.n26 585
R232 B.n278 B.n277 585
R233 B.n279 B.n25 585
R234 B.n281 B.n280 585
R235 B.n282 B.n24 585
R236 B.n284 B.n283 585
R237 B.n285 B.n23 585
R238 B.n287 B.n286 585
R239 B.n289 B.n288 585
R240 B.n290 B.n19 585
R241 B.n292 B.n291 585
R242 B.n293 B.n18 585
R243 B.n295 B.n294 585
R244 B.n296 B.n17 585
R245 B.n298 B.n297 585
R246 B.n299 B.n16 585
R247 B.n301 B.n300 585
R248 B.n302 B.n15 585
R249 B.n304 B.n303 585
R250 B.n305 B.n14 585
R251 B.n307 B.n306 585
R252 B.n308 B.n13 585
R253 B.n310 B.n309 585
R254 B.n248 B.n37 585
R255 B.n247 B.n246 585
R256 B.n245 B.n38 585
R257 B.n244 B.n243 585
R258 B.n242 B.n39 585
R259 B.n241 B.n240 585
R260 B.n239 B.n40 585
R261 B.n238 B.n237 585
R262 B.n236 B.n41 585
R263 B.n235 B.n234 585
R264 B.n233 B.n42 585
R265 B.n232 B.n231 585
R266 B.n230 B.n43 585
R267 B.n229 B.n228 585
R268 B.n227 B.n44 585
R269 B.n226 B.n225 585
R270 B.n224 B.n45 585
R271 B.n223 B.n222 585
R272 B.n221 B.n46 585
R273 B.n220 B.n219 585
R274 B.n218 B.n47 585
R275 B.n217 B.n216 585
R276 B.n215 B.n48 585
R277 B.n214 B.n213 585
R278 B.n212 B.n49 585
R279 B.n211 B.n210 585
R280 B.n209 B.n50 585
R281 B.n208 B.n207 585
R282 B.n206 B.n51 585
R283 B.n205 B.n204 585
R284 B.n203 B.n52 585
R285 B.n202 B.n201 585
R286 B.n200 B.n53 585
R287 B.n199 B.n198 585
R288 B.n197 B.n54 585
R289 B.n196 B.n195 585
R290 B.n194 B.n55 585
R291 B.n193 B.n192 585
R292 B.n191 B.n56 585
R293 B.n190 B.n189 585
R294 B.n188 B.n57 585
R295 B.n187 B.n186 585
R296 B.n185 B.n58 585
R297 B.n124 B.n123 585
R298 B.n125 B.n82 585
R299 B.n127 B.n126 585
R300 B.n128 B.n81 585
R301 B.n130 B.n129 585
R302 B.n131 B.n80 585
R303 B.n133 B.n132 585
R304 B.n134 B.n79 585
R305 B.n136 B.n135 585
R306 B.n137 B.n78 585
R307 B.n139 B.n138 585
R308 B.n140 B.n77 585
R309 B.n142 B.n141 585
R310 B.n143 B.n76 585
R311 B.n145 B.n144 585
R312 B.n147 B.n73 585
R313 B.n149 B.n148 585
R314 B.n150 B.n72 585
R315 B.n152 B.n151 585
R316 B.n153 B.n71 585
R317 B.n155 B.n154 585
R318 B.n156 B.n70 585
R319 B.n158 B.n157 585
R320 B.n159 B.n69 585
R321 B.n161 B.n160 585
R322 B.n163 B.n162 585
R323 B.n164 B.n65 585
R324 B.n166 B.n165 585
R325 B.n167 B.n64 585
R326 B.n169 B.n168 585
R327 B.n170 B.n63 585
R328 B.n172 B.n171 585
R329 B.n173 B.n62 585
R330 B.n175 B.n174 585
R331 B.n176 B.n61 585
R332 B.n178 B.n177 585
R333 B.n179 B.n60 585
R334 B.n181 B.n180 585
R335 B.n182 B.n59 585
R336 B.n184 B.n183 585
R337 B.n122 B.n83 585
R338 B.n121 B.n120 585
R339 B.n119 B.n84 585
R340 B.n118 B.n117 585
R341 B.n116 B.n85 585
R342 B.n115 B.n114 585
R343 B.n113 B.n86 585
R344 B.n112 B.n111 585
R345 B.n110 B.n87 585
R346 B.n109 B.n108 585
R347 B.n107 B.n88 585
R348 B.n106 B.n105 585
R349 B.n104 B.n89 585
R350 B.n103 B.n102 585
R351 B.n101 B.n90 585
R352 B.n100 B.n99 585
R353 B.n98 B.n91 585
R354 B.n97 B.n96 585
R355 B.n95 B.n92 585
R356 B.n94 B.n93 585
R357 B.n2 B.n0 585
R358 B.n341 B.n1 585
R359 B.n340 B.n339 585
R360 B.n338 B.n3 585
R361 B.n337 B.n336 585
R362 B.n335 B.n4 585
R363 B.n334 B.n333 585
R364 B.n332 B.n5 585
R365 B.n331 B.n330 585
R366 B.n329 B.n6 585
R367 B.n328 B.n327 585
R368 B.n326 B.n7 585
R369 B.n325 B.n324 585
R370 B.n323 B.n8 585
R371 B.n322 B.n321 585
R372 B.n320 B.n9 585
R373 B.n319 B.n318 585
R374 B.n317 B.n10 585
R375 B.n316 B.n315 585
R376 B.n314 B.n11 585
R377 B.n313 B.n312 585
R378 B.n311 B.n12 585
R379 B.n343 B.n342 585
R380 B.n124 B.n83 521.33
R381 B.n311 B.n310 521.33
R382 B.n185 B.n184 521.33
R383 B.n250 B.n37 521.33
R384 B.n66 B.t0 269.211
R385 B.n74 B.t6 269.211
R386 B.n20 B.t9 269.211
R387 B.n28 B.t3 269.211
R388 B.n66 B.t2 251.355
R389 B.n28 B.t4 251.355
R390 B.n74 B.t8 251.355
R391 B.n20 B.t10 251.355
R392 B.n67 B.t1 223.04
R393 B.n29 B.t5 223.04
R394 B.n75 B.t7 223.04
R395 B.n21 B.t11 223.04
R396 B.n120 B.n83 163.367
R397 B.n120 B.n119 163.367
R398 B.n119 B.n118 163.367
R399 B.n118 B.n85 163.367
R400 B.n114 B.n85 163.367
R401 B.n114 B.n113 163.367
R402 B.n113 B.n112 163.367
R403 B.n112 B.n87 163.367
R404 B.n108 B.n87 163.367
R405 B.n108 B.n107 163.367
R406 B.n107 B.n106 163.367
R407 B.n106 B.n89 163.367
R408 B.n102 B.n89 163.367
R409 B.n102 B.n101 163.367
R410 B.n101 B.n100 163.367
R411 B.n100 B.n91 163.367
R412 B.n96 B.n91 163.367
R413 B.n96 B.n95 163.367
R414 B.n95 B.n94 163.367
R415 B.n94 B.n2 163.367
R416 B.n342 B.n2 163.367
R417 B.n342 B.n341 163.367
R418 B.n341 B.n340 163.367
R419 B.n340 B.n3 163.367
R420 B.n336 B.n3 163.367
R421 B.n336 B.n335 163.367
R422 B.n335 B.n334 163.367
R423 B.n334 B.n5 163.367
R424 B.n330 B.n5 163.367
R425 B.n330 B.n329 163.367
R426 B.n329 B.n328 163.367
R427 B.n328 B.n7 163.367
R428 B.n324 B.n7 163.367
R429 B.n324 B.n323 163.367
R430 B.n323 B.n322 163.367
R431 B.n322 B.n9 163.367
R432 B.n318 B.n9 163.367
R433 B.n318 B.n317 163.367
R434 B.n317 B.n316 163.367
R435 B.n316 B.n11 163.367
R436 B.n312 B.n11 163.367
R437 B.n312 B.n311 163.367
R438 B.n125 B.n124 163.367
R439 B.n126 B.n125 163.367
R440 B.n126 B.n81 163.367
R441 B.n130 B.n81 163.367
R442 B.n131 B.n130 163.367
R443 B.n132 B.n131 163.367
R444 B.n132 B.n79 163.367
R445 B.n136 B.n79 163.367
R446 B.n137 B.n136 163.367
R447 B.n138 B.n137 163.367
R448 B.n138 B.n77 163.367
R449 B.n142 B.n77 163.367
R450 B.n143 B.n142 163.367
R451 B.n144 B.n143 163.367
R452 B.n144 B.n73 163.367
R453 B.n149 B.n73 163.367
R454 B.n150 B.n149 163.367
R455 B.n151 B.n150 163.367
R456 B.n151 B.n71 163.367
R457 B.n155 B.n71 163.367
R458 B.n156 B.n155 163.367
R459 B.n157 B.n156 163.367
R460 B.n157 B.n69 163.367
R461 B.n161 B.n69 163.367
R462 B.n162 B.n161 163.367
R463 B.n162 B.n65 163.367
R464 B.n166 B.n65 163.367
R465 B.n167 B.n166 163.367
R466 B.n168 B.n167 163.367
R467 B.n168 B.n63 163.367
R468 B.n172 B.n63 163.367
R469 B.n173 B.n172 163.367
R470 B.n174 B.n173 163.367
R471 B.n174 B.n61 163.367
R472 B.n178 B.n61 163.367
R473 B.n179 B.n178 163.367
R474 B.n180 B.n179 163.367
R475 B.n180 B.n59 163.367
R476 B.n184 B.n59 163.367
R477 B.n186 B.n185 163.367
R478 B.n186 B.n57 163.367
R479 B.n190 B.n57 163.367
R480 B.n191 B.n190 163.367
R481 B.n192 B.n191 163.367
R482 B.n192 B.n55 163.367
R483 B.n196 B.n55 163.367
R484 B.n197 B.n196 163.367
R485 B.n198 B.n197 163.367
R486 B.n198 B.n53 163.367
R487 B.n202 B.n53 163.367
R488 B.n203 B.n202 163.367
R489 B.n204 B.n203 163.367
R490 B.n204 B.n51 163.367
R491 B.n208 B.n51 163.367
R492 B.n209 B.n208 163.367
R493 B.n210 B.n209 163.367
R494 B.n210 B.n49 163.367
R495 B.n214 B.n49 163.367
R496 B.n215 B.n214 163.367
R497 B.n216 B.n215 163.367
R498 B.n216 B.n47 163.367
R499 B.n220 B.n47 163.367
R500 B.n221 B.n220 163.367
R501 B.n222 B.n221 163.367
R502 B.n222 B.n45 163.367
R503 B.n226 B.n45 163.367
R504 B.n227 B.n226 163.367
R505 B.n228 B.n227 163.367
R506 B.n228 B.n43 163.367
R507 B.n232 B.n43 163.367
R508 B.n233 B.n232 163.367
R509 B.n234 B.n233 163.367
R510 B.n234 B.n41 163.367
R511 B.n238 B.n41 163.367
R512 B.n239 B.n238 163.367
R513 B.n240 B.n239 163.367
R514 B.n240 B.n39 163.367
R515 B.n244 B.n39 163.367
R516 B.n245 B.n244 163.367
R517 B.n246 B.n245 163.367
R518 B.n246 B.n37 163.367
R519 B.n310 B.n13 163.367
R520 B.n306 B.n13 163.367
R521 B.n306 B.n305 163.367
R522 B.n305 B.n304 163.367
R523 B.n304 B.n15 163.367
R524 B.n300 B.n15 163.367
R525 B.n300 B.n299 163.367
R526 B.n299 B.n298 163.367
R527 B.n298 B.n17 163.367
R528 B.n294 B.n17 163.367
R529 B.n294 B.n293 163.367
R530 B.n293 B.n292 163.367
R531 B.n292 B.n19 163.367
R532 B.n288 B.n19 163.367
R533 B.n288 B.n287 163.367
R534 B.n287 B.n23 163.367
R535 B.n283 B.n23 163.367
R536 B.n283 B.n282 163.367
R537 B.n282 B.n281 163.367
R538 B.n281 B.n25 163.367
R539 B.n277 B.n25 163.367
R540 B.n277 B.n276 163.367
R541 B.n276 B.n275 163.367
R542 B.n275 B.n27 163.367
R543 B.n270 B.n27 163.367
R544 B.n270 B.n269 163.367
R545 B.n269 B.n268 163.367
R546 B.n268 B.n31 163.367
R547 B.n264 B.n31 163.367
R548 B.n264 B.n263 163.367
R549 B.n263 B.n262 163.367
R550 B.n262 B.n33 163.367
R551 B.n258 B.n33 163.367
R552 B.n258 B.n257 163.367
R553 B.n257 B.n256 163.367
R554 B.n256 B.n35 163.367
R555 B.n252 B.n35 163.367
R556 B.n252 B.n251 163.367
R557 B.n251 B.n250 163.367
R558 B.n68 B.n67 59.5399
R559 B.n146 B.n75 59.5399
R560 B.n22 B.n21 59.5399
R561 B.n272 B.n29 59.5399
R562 B.n309 B.n12 33.8737
R563 B.n249 B.n248 33.8737
R564 B.n183 B.n58 33.8737
R565 B.n123 B.n122 33.8737
R566 B.n67 B.n66 28.3157
R567 B.n75 B.n74 28.3157
R568 B.n21 B.n20 28.3157
R569 B.n29 B.n28 28.3157
R570 B B.n343 18.0485
R571 B.n309 B.n308 10.6151
R572 B.n308 B.n307 10.6151
R573 B.n307 B.n14 10.6151
R574 B.n303 B.n14 10.6151
R575 B.n303 B.n302 10.6151
R576 B.n302 B.n301 10.6151
R577 B.n301 B.n16 10.6151
R578 B.n297 B.n16 10.6151
R579 B.n297 B.n296 10.6151
R580 B.n296 B.n295 10.6151
R581 B.n295 B.n18 10.6151
R582 B.n291 B.n18 10.6151
R583 B.n291 B.n290 10.6151
R584 B.n290 B.n289 10.6151
R585 B.n286 B.n285 10.6151
R586 B.n285 B.n284 10.6151
R587 B.n284 B.n24 10.6151
R588 B.n280 B.n24 10.6151
R589 B.n280 B.n279 10.6151
R590 B.n279 B.n278 10.6151
R591 B.n278 B.n26 10.6151
R592 B.n274 B.n26 10.6151
R593 B.n274 B.n273 10.6151
R594 B.n271 B.n30 10.6151
R595 B.n267 B.n30 10.6151
R596 B.n267 B.n266 10.6151
R597 B.n266 B.n265 10.6151
R598 B.n265 B.n32 10.6151
R599 B.n261 B.n32 10.6151
R600 B.n261 B.n260 10.6151
R601 B.n260 B.n259 10.6151
R602 B.n259 B.n34 10.6151
R603 B.n255 B.n34 10.6151
R604 B.n255 B.n254 10.6151
R605 B.n254 B.n253 10.6151
R606 B.n253 B.n36 10.6151
R607 B.n249 B.n36 10.6151
R608 B.n187 B.n58 10.6151
R609 B.n188 B.n187 10.6151
R610 B.n189 B.n188 10.6151
R611 B.n189 B.n56 10.6151
R612 B.n193 B.n56 10.6151
R613 B.n194 B.n193 10.6151
R614 B.n195 B.n194 10.6151
R615 B.n195 B.n54 10.6151
R616 B.n199 B.n54 10.6151
R617 B.n200 B.n199 10.6151
R618 B.n201 B.n200 10.6151
R619 B.n201 B.n52 10.6151
R620 B.n205 B.n52 10.6151
R621 B.n206 B.n205 10.6151
R622 B.n207 B.n206 10.6151
R623 B.n207 B.n50 10.6151
R624 B.n211 B.n50 10.6151
R625 B.n212 B.n211 10.6151
R626 B.n213 B.n212 10.6151
R627 B.n213 B.n48 10.6151
R628 B.n217 B.n48 10.6151
R629 B.n218 B.n217 10.6151
R630 B.n219 B.n218 10.6151
R631 B.n219 B.n46 10.6151
R632 B.n223 B.n46 10.6151
R633 B.n224 B.n223 10.6151
R634 B.n225 B.n224 10.6151
R635 B.n225 B.n44 10.6151
R636 B.n229 B.n44 10.6151
R637 B.n230 B.n229 10.6151
R638 B.n231 B.n230 10.6151
R639 B.n231 B.n42 10.6151
R640 B.n235 B.n42 10.6151
R641 B.n236 B.n235 10.6151
R642 B.n237 B.n236 10.6151
R643 B.n237 B.n40 10.6151
R644 B.n241 B.n40 10.6151
R645 B.n242 B.n241 10.6151
R646 B.n243 B.n242 10.6151
R647 B.n243 B.n38 10.6151
R648 B.n247 B.n38 10.6151
R649 B.n248 B.n247 10.6151
R650 B.n123 B.n82 10.6151
R651 B.n127 B.n82 10.6151
R652 B.n128 B.n127 10.6151
R653 B.n129 B.n128 10.6151
R654 B.n129 B.n80 10.6151
R655 B.n133 B.n80 10.6151
R656 B.n134 B.n133 10.6151
R657 B.n135 B.n134 10.6151
R658 B.n135 B.n78 10.6151
R659 B.n139 B.n78 10.6151
R660 B.n140 B.n139 10.6151
R661 B.n141 B.n140 10.6151
R662 B.n141 B.n76 10.6151
R663 B.n145 B.n76 10.6151
R664 B.n148 B.n147 10.6151
R665 B.n148 B.n72 10.6151
R666 B.n152 B.n72 10.6151
R667 B.n153 B.n152 10.6151
R668 B.n154 B.n153 10.6151
R669 B.n154 B.n70 10.6151
R670 B.n158 B.n70 10.6151
R671 B.n159 B.n158 10.6151
R672 B.n160 B.n159 10.6151
R673 B.n164 B.n163 10.6151
R674 B.n165 B.n164 10.6151
R675 B.n165 B.n64 10.6151
R676 B.n169 B.n64 10.6151
R677 B.n170 B.n169 10.6151
R678 B.n171 B.n170 10.6151
R679 B.n171 B.n62 10.6151
R680 B.n175 B.n62 10.6151
R681 B.n176 B.n175 10.6151
R682 B.n177 B.n176 10.6151
R683 B.n177 B.n60 10.6151
R684 B.n181 B.n60 10.6151
R685 B.n182 B.n181 10.6151
R686 B.n183 B.n182 10.6151
R687 B.n122 B.n121 10.6151
R688 B.n121 B.n84 10.6151
R689 B.n117 B.n84 10.6151
R690 B.n117 B.n116 10.6151
R691 B.n116 B.n115 10.6151
R692 B.n115 B.n86 10.6151
R693 B.n111 B.n86 10.6151
R694 B.n111 B.n110 10.6151
R695 B.n110 B.n109 10.6151
R696 B.n109 B.n88 10.6151
R697 B.n105 B.n88 10.6151
R698 B.n105 B.n104 10.6151
R699 B.n104 B.n103 10.6151
R700 B.n103 B.n90 10.6151
R701 B.n99 B.n90 10.6151
R702 B.n99 B.n98 10.6151
R703 B.n98 B.n97 10.6151
R704 B.n97 B.n92 10.6151
R705 B.n93 B.n92 10.6151
R706 B.n93 B.n0 10.6151
R707 B.n339 B.n1 10.6151
R708 B.n339 B.n338 10.6151
R709 B.n338 B.n337 10.6151
R710 B.n337 B.n4 10.6151
R711 B.n333 B.n4 10.6151
R712 B.n333 B.n332 10.6151
R713 B.n332 B.n331 10.6151
R714 B.n331 B.n6 10.6151
R715 B.n327 B.n6 10.6151
R716 B.n327 B.n326 10.6151
R717 B.n326 B.n325 10.6151
R718 B.n325 B.n8 10.6151
R719 B.n321 B.n8 10.6151
R720 B.n321 B.n320 10.6151
R721 B.n320 B.n319 10.6151
R722 B.n319 B.n10 10.6151
R723 B.n315 B.n10 10.6151
R724 B.n315 B.n314 10.6151
R725 B.n314 B.n313 10.6151
R726 B.n313 B.n12 10.6151
R727 B.n289 B.n22 9.36635
R728 B.n272 B.n271 9.36635
R729 B.n146 B.n145 9.36635
R730 B.n163 B.n68 9.36635
R731 B.n343 B.n0 2.81026
R732 B.n343 B.n1 2.81026
R733 B.n286 B.n22 1.24928
R734 B.n273 B.n272 1.24928
R735 B.n147 B.n146 1.24928
R736 B.n160 B.n68 1.24928
R737 VP.n0 VP.t0 119.059
R738 VP.n0 VP.t3 118.972
R739 VP.n2 VP.t2 100.453
R740 VP.n3 VP.t1 100.453
R741 VP.n4 VP.n3 80.6037
R742 VP.n2 VP.n1 80.6037
R743 VP.n1 VP.n0 66.3895
R744 VP.n3 VP.n2 48.2005
R745 VP.n4 VP.n1 0.380177
R746 VP VP.n4 0.146778
R747 VDD1 VDD1.n1 157.543
R748 VDD1 VDD1.n0 126.939
R749 VDD1.n0 VDD1.t3 10.5884
R750 VDD1.n0 VDD1.t0 10.5884
R751 VDD1.n1 VDD1.t1 10.5884
R752 VDD1.n1 VDD1.t2 10.5884
C0 VN VDD1 0.152634f
C1 VP VDD1 1.35138f
C2 B VDD2 0.789325f
C3 VN w_n1846_n1582# 2.65986f
C4 VP w_n1846_n1582# 2.89124f
C5 VTAIL VDD1 2.76885f
C6 VN VP 3.48074f
C7 VTAIL w_n1846_n1582# 1.84356f
C8 VDD2 VDD1 0.669657f
C9 B VDD1 0.760998f
C10 VDD2 w_n1846_n1582# 0.941227f
C11 B w_n1846_n1582# 4.93315f
C12 VN VTAIL 1.34404f
C13 VP VTAIL 1.35815f
C14 VN VDD2 1.19868f
C15 B VN 0.716874f
C16 VP VDD2 0.306219f
C17 B VP 1.09726f
C18 VDD1 w_n1846_n1582# 0.918163f
C19 VTAIL VDD2 2.81321f
C20 B VTAIL 1.53095f
C21 VDD2 VSUBS 0.474237f
C22 VDD1 VSUBS 2.626815f
C23 VTAIL VSUBS 0.377409f
C24 VN VSUBS 4.13643f
C25 VP VSUBS 1.100072f
C26 B VSUBS 2.136547f
C27 w_n1846_n1582# VSUBS 36.9717f
C28 VDD1.t3 VSUBS 0.044794f
C29 VDD1.t0 VSUBS 0.044794f
C30 VDD1.n0 VSUBS 0.238831f
C31 VDD1.t1 VSUBS 0.044794f
C32 VDD1.t2 VSUBS 0.044794f
C33 VDD1.n1 VSUBS 0.396944f
C34 VP.t3 VSUBS 0.545128f
C35 VP.t0 VSUBS 0.545388f
C36 VP.n0 VSUBS 1.3335f
C37 VP.n1 VSUBS 2.29051f
C38 VP.t2 VSUBS 0.500755f
C39 VP.n2 VSUBS 0.285059f
C40 VP.t1 VSUBS 0.500755f
C41 VP.n3 VSUBS 0.285059f
C42 VP.n4 VSUBS 0.061208f
C43 B.n0 VSUBS 0.004995f
C44 B.n1 VSUBS 0.004995f
C45 B.n2 VSUBS 0.007899f
C46 B.n3 VSUBS 0.007899f
C47 B.n4 VSUBS 0.007899f
C48 B.n5 VSUBS 0.007899f
C49 B.n6 VSUBS 0.007899f
C50 B.n7 VSUBS 0.007899f
C51 B.n8 VSUBS 0.007899f
C52 B.n9 VSUBS 0.007899f
C53 B.n10 VSUBS 0.007899f
C54 B.n11 VSUBS 0.007899f
C55 B.n12 VSUBS 0.018616f
C56 B.n13 VSUBS 0.007899f
C57 B.n14 VSUBS 0.007899f
C58 B.n15 VSUBS 0.007899f
C59 B.n16 VSUBS 0.007899f
C60 B.n17 VSUBS 0.007899f
C61 B.n18 VSUBS 0.007899f
C62 B.n19 VSUBS 0.007899f
C63 B.t11 VSUBS 0.050746f
C64 B.t10 VSUBS 0.060782f
C65 B.t9 VSUBS 0.184053f
C66 B.n20 VSUBS 0.111401f
C67 B.n21 VSUBS 0.100358f
C68 B.n22 VSUBS 0.018301f
C69 B.n23 VSUBS 0.007899f
C70 B.n24 VSUBS 0.007899f
C71 B.n25 VSUBS 0.007899f
C72 B.n26 VSUBS 0.007899f
C73 B.n27 VSUBS 0.007899f
C74 B.t5 VSUBS 0.050746f
C75 B.t4 VSUBS 0.060783f
C76 B.t3 VSUBS 0.184053f
C77 B.n28 VSUBS 0.1114f
C78 B.n29 VSUBS 0.100358f
C79 B.n30 VSUBS 0.007899f
C80 B.n31 VSUBS 0.007899f
C81 B.n32 VSUBS 0.007899f
C82 B.n33 VSUBS 0.007899f
C83 B.n34 VSUBS 0.007899f
C84 B.n35 VSUBS 0.007899f
C85 B.n36 VSUBS 0.007899f
C86 B.n37 VSUBS 0.018616f
C87 B.n38 VSUBS 0.007899f
C88 B.n39 VSUBS 0.007899f
C89 B.n40 VSUBS 0.007899f
C90 B.n41 VSUBS 0.007899f
C91 B.n42 VSUBS 0.007899f
C92 B.n43 VSUBS 0.007899f
C93 B.n44 VSUBS 0.007899f
C94 B.n45 VSUBS 0.007899f
C95 B.n46 VSUBS 0.007899f
C96 B.n47 VSUBS 0.007899f
C97 B.n48 VSUBS 0.007899f
C98 B.n49 VSUBS 0.007899f
C99 B.n50 VSUBS 0.007899f
C100 B.n51 VSUBS 0.007899f
C101 B.n52 VSUBS 0.007899f
C102 B.n53 VSUBS 0.007899f
C103 B.n54 VSUBS 0.007899f
C104 B.n55 VSUBS 0.007899f
C105 B.n56 VSUBS 0.007899f
C106 B.n57 VSUBS 0.007899f
C107 B.n58 VSUBS 0.018616f
C108 B.n59 VSUBS 0.007899f
C109 B.n60 VSUBS 0.007899f
C110 B.n61 VSUBS 0.007899f
C111 B.n62 VSUBS 0.007899f
C112 B.n63 VSUBS 0.007899f
C113 B.n64 VSUBS 0.007899f
C114 B.n65 VSUBS 0.007899f
C115 B.t1 VSUBS 0.050746f
C116 B.t2 VSUBS 0.060783f
C117 B.t0 VSUBS 0.184053f
C118 B.n66 VSUBS 0.1114f
C119 B.n67 VSUBS 0.100358f
C120 B.n68 VSUBS 0.018301f
C121 B.n69 VSUBS 0.007899f
C122 B.n70 VSUBS 0.007899f
C123 B.n71 VSUBS 0.007899f
C124 B.n72 VSUBS 0.007899f
C125 B.n73 VSUBS 0.007899f
C126 B.t7 VSUBS 0.050746f
C127 B.t8 VSUBS 0.060782f
C128 B.t6 VSUBS 0.184053f
C129 B.n74 VSUBS 0.111401f
C130 B.n75 VSUBS 0.100358f
C131 B.n76 VSUBS 0.007899f
C132 B.n77 VSUBS 0.007899f
C133 B.n78 VSUBS 0.007899f
C134 B.n79 VSUBS 0.007899f
C135 B.n80 VSUBS 0.007899f
C136 B.n81 VSUBS 0.007899f
C137 B.n82 VSUBS 0.007899f
C138 B.n83 VSUBS 0.018616f
C139 B.n84 VSUBS 0.007899f
C140 B.n85 VSUBS 0.007899f
C141 B.n86 VSUBS 0.007899f
C142 B.n87 VSUBS 0.007899f
C143 B.n88 VSUBS 0.007899f
C144 B.n89 VSUBS 0.007899f
C145 B.n90 VSUBS 0.007899f
C146 B.n91 VSUBS 0.007899f
C147 B.n92 VSUBS 0.007899f
C148 B.n93 VSUBS 0.007899f
C149 B.n94 VSUBS 0.007899f
C150 B.n95 VSUBS 0.007899f
C151 B.n96 VSUBS 0.007899f
C152 B.n97 VSUBS 0.007899f
C153 B.n98 VSUBS 0.007899f
C154 B.n99 VSUBS 0.007899f
C155 B.n100 VSUBS 0.007899f
C156 B.n101 VSUBS 0.007899f
C157 B.n102 VSUBS 0.007899f
C158 B.n103 VSUBS 0.007899f
C159 B.n104 VSUBS 0.007899f
C160 B.n105 VSUBS 0.007899f
C161 B.n106 VSUBS 0.007899f
C162 B.n107 VSUBS 0.007899f
C163 B.n108 VSUBS 0.007899f
C164 B.n109 VSUBS 0.007899f
C165 B.n110 VSUBS 0.007899f
C166 B.n111 VSUBS 0.007899f
C167 B.n112 VSUBS 0.007899f
C168 B.n113 VSUBS 0.007899f
C169 B.n114 VSUBS 0.007899f
C170 B.n115 VSUBS 0.007899f
C171 B.n116 VSUBS 0.007899f
C172 B.n117 VSUBS 0.007899f
C173 B.n118 VSUBS 0.007899f
C174 B.n119 VSUBS 0.007899f
C175 B.n120 VSUBS 0.007899f
C176 B.n121 VSUBS 0.007899f
C177 B.n122 VSUBS 0.018616f
C178 B.n123 VSUBS 0.019253f
C179 B.n124 VSUBS 0.019253f
C180 B.n125 VSUBS 0.007899f
C181 B.n126 VSUBS 0.007899f
C182 B.n127 VSUBS 0.007899f
C183 B.n128 VSUBS 0.007899f
C184 B.n129 VSUBS 0.007899f
C185 B.n130 VSUBS 0.007899f
C186 B.n131 VSUBS 0.007899f
C187 B.n132 VSUBS 0.007899f
C188 B.n133 VSUBS 0.007899f
C189 B.n134 VSUBS 0.007899f
C190 B.n135 VSUBS 0.007899f
C191 B.n136 VSUBS 0.007899f
C192 B.n137 VSUBS 0.007899f
C193 B.n138 VSUBS 0.007899f
C194 B.n139 VSUBS 0.007899f
C195 B.n140 VSUBS 0.007899f
C196 B.n141 VSUBS 0.007899f
C197 B.n142 VSUBS 0.007899f
C198 B.n143 VSUBS 0.007899f
C199 B.n144 VSUBS 0.007899f
C200 B.n145 VSUBS 0.007434f
C201 B.n146 VSUBS 0.018301f
C202 B.n147 VSUBS 0.004414f
C203 B.n148 VSUBS 0.007899f
C204 B.n149 VSUBS 0.007899f
C205 B.n150 VSUBS 0.007899f
C206 B.n151 VSUBS 0.007899f
C207 B.n152 VSUBS 0.007899f
C208 B.n153 VSUBS 0.007899f
C209 B.n154 VSUBS 0.007899f
C210 B.n155 VSUBS 0.007899f
C211 B.n156 VSUBS 0.007899f
C212 B.n157 VSUBS 0.007899f
C213 B.n158 VSUBS 0.007899f
C214 B.n159 VSUBS 0.007899f
C215 B.n160 VSUBS 0.004414f
C216 B.n161 VSUBS 0.007899f
C217 B.n162 VSUBS 0.007899f
C218 B.n163 VSUBS 0.007434f
C219 B.n164 VSUBS 0.007899f
C220 B.n165 VSUBS 0.007899f
C221 B.n166 VSUBS 0.007899f
C222 B.n167 VSUBS 0.007899f
C223 B.n168 VSUBS 0.007899f
C224 B.n169 VSUBS 0.007899f
C225 B.n170 VSUBS 0.007899f
C226 B.n171 VSUBS 0.007899f
C227 B.n172 VSUBS 0.007899f
C228 B.n173 VSUBS 0.007899f
C229 B.n174 VSUBS 0.007899f
C230 B.n175 VSUBS 0.007899f
C231 B.n176 VSUBS 0.007899f
C232 B.n177 VSUBS 0.007899f
C233 B.n178 VSUBS 0.007899f
C234 B.n179 VSUBS 0.007899f
C235 B.n180 VSUBS 0.007899f
C236 B.n181 VSUBS 0.007899f
C237 B.n182 VSUBS 0.007899f
C238 B.n183 VSUBS 0.019253f
C239 B.n184 VSUBS 0.019253f
C240 B.n185 VSUBS 0.018616f
C241 B.n186 VSUBS 0.007899f
C242 B.n187 VSUBS 0.007899f
C243 B.n188 VSUBS 0.007899f
C244 B.n189 VSUBS 0.007899f
C245 B.n190 VSUBS 0.007899f
C246 B.n191 VSUBS 0.007899f
C247 B.n192 VSUBS 0.007899f
C248 B.n193 VSUBS 0.007899f
C249 B.n194 VSUBS 0.007899f
C250 B.n195 VSUBS 0.007899f
C251 B.n196 VSUBS 0.007899f
C252 B.n197 VSUBS 0.007899f
C253 B.n198 VSUBS 0.007899f
C254 B.n199 VSUBS 0.007899f
C255 B.n200 VSUBS 0.007899f
C256 B.n201 VSUBS 0.007899f
C257 B.n202 VSUBS 0.007899f
C258 B.n203 VSUBS 0.007899f
C259 B.n204 VSUBS 0.007899f
C260 B.n205 VSUBS 0.007899f
C261 B.n206 VSUBS 0.007899f
C262 B.n207 VSUBS 0.007899f
C263 B.n208 VSUBS 0.007899f
C264 B.n209 VSUBS 0.007899f
C265 B.n210 VSUBS 0.007899f
C266 B.n211 VSUBS 0.007899f
C267 B.n212 VSUBS 0.007899f
C268 B.n213 VSUBS 0.007899f
C269 B.n214 VSUBS 0.007899f
C270 B.n215 VSUBS 0.007899f
C271 B.n216 VSUBS 0.007899f
C272 B.n217 VSUBS 0.007899f
C273 B.n218 VSUBS 0.007899f
C274 B.n219 VSUBS 0.007899f
C275 B.n220 VSUBS 0.007899f
C276 B.n221 VSUBS 0.007899f
C277 B.n222 VSUBS 0.007899f
C278 B.n223 VSUBS 0.007899f
C279 B.n224 VSUBS 0.007899f
C280 B.n225 VSUBS 0.007899f
C281 B.n226 VSUBS 0.007899f
C282 B.n227 VSUBS 0.007899f
C283 B.n228 VSUBS 0.007899f
C284 B.n229 VSUBS 0.007899f
C285 B.n230 VSUBS 0.007899f
C286 B.n231 VSUBS 0.007899f
C287 B.n232 VSUBS 0.007899f
C288 B.n233 VSUBS 0.007899f
C289 B.n234 VSUBS 0.007899f
C290 B.n235 VSUBS 0.007899f
C291 B.n236 VSUBS 0.007899f
C292 B.n237 VSUBS 0.007899f
C293 B.n238 VSUBS 0.007899f
C294 B.n239 VSUBS 0.007899f
C295 B.n240 VSUBS 0.007899f
C296 B.n241 VSUBS 0.007899f
C297 B.n242 VSUBS 0.007899f
C298 B.n243 VSUBS 0.007899f
C299 B.n244 VSUBS 0.007899f
C300 B.n245 VSUBS 0.007899f
C301 B.n246 VSUBS 0.007899f
C302 B.n247 VSUBS 0.007899f
C303 B.n248 VSUBS 0.019516f
C304 B.n249 VSUBS 0.018353f
C305 B.n250 VSUBS 0.019253f
C306 B.n251 VSUBS 0.007899f
C307 B.n252 VSUBS 0.007899f
C308 B.n253 VSUBS 0.007899f
C309 B.n254 VSUBS 0.007899f
C310 B.n255 VSUBS 0.007899f
C311 B.n256 VSUBS 0.007899f
C312 B.n257 VSUBS 0.007899f
C313 B.n258 VSUBS 0.007899f
C314 B.n259 VSUBS 0.007899f
C315 B.n260 VSUBS 0.007899f
C316 B.n261 VSUBS 0.007899f
C317 B.n262 VSUBS 0.007899f
C318 B.n263 VSUBS 0.007899f
C319 B.n264 VSUBS 0.007899f
C320 B.n265 VSUBS 0.007899f
C321 B.n266 VSUBS 0.007899f
C322 B.n267 VSUBS 0.007899f
C323 B.n268 VSUBS 0.007899f
C324 B.n269 VSUBS 0.007899f
C325 B.n270 VSUBS 0.007899f
C326 B.n271 VSUBS 0.007434f
C327 B.n272 VSUBS 0.018301f
C328 B.n273 VSUBS 0.004414f
C329 B.n274 VSUBS 0.007899f
C330 B.n275 VSUBS 0.007899f
C331 B.n276 VSUBS 0.007899f
C332 B.n277 VSUBS 0.007899f
C333 B.n278 VSUBS 0.007899f
C334 B.n279 VSUBS 0.007899f
C335 B.n280 VSUBS 0.007899f
C336 B.n281 VSUBS 0.007899f
C337 B.n282 VSUBS 0.007899f
C338 B.n283 VSUBS 0.007899f
C339 B.n284 VSUBS 0.007899f
C340 B.n285 VSUBS 0.007899f
C341 B.n286 VSUBS 0.004414f
C342 B.n287 VSUBS 0.007899f
C343 B.n288 VSUBS 0.007899f
C344 B.n289 VSUBS 0.007434f
C345 B.n290 VSUBS 0.007899f
C346 B.n291 VSUBS 0.007899f
C347 B.n292 VSUBS 0.007899f
C348 B.n293 VSUBS 0.007899f
C349 B.n294 VSUBS 0.007899f
C350 B.n295 VSUBS 0.007899f
C351 B.n296 VSUBS 0.007899f
C352 B.n297 VSUBS 0.007899f
C353 B.n298 VSUBS 0.007899f
C354 B.n299 VSUBS 0.007899f
C355 B.n300 VSUBS 0.007899f
C356 B.n301 VSUBS 0.007899f
C357 B.n302 VSUBS 0.007899f
C358 B.n303 VSUBS 0.007899f
C359 B.n304 VSUBS 0.007899f
C360 B.n305 VSUBS 0.007899f
C361 B.n306 VSUBS 0.007899f
C362 B.n307 VSUBS 0.007899f
C363 B.n308 VSUBS 0.007899f
C364 B.n309 VSUBS 0.019253f
C365 B.n310 VSUBS 0.019253f
C366 B.n311 VSUBS 0.018616f
C367 B.n312 VSUBS 0.007899f
C368 B.n313 VSUBS 0.007899f
C369 B.n314 VSUBS 0.007899f
C370 B.n315 VSUBS 0.007899f
C371 B.n316 VSUBS 0.007899f
C372 B.n317 VSUBS 0.007899f
C373 B.n318 VSUBS 0.007899f
C374 B.n319 VSUBS 0.007899f
C375 B.n320 VSUBS 0.007899f
C376 B.n321 VSUBS 0.007899f
C377 B.n322 VSUBS 0.007899f
C378 B.n323 VSUBS 0.007899f
C379 B.n324 VSUBS 0.007899f
C380 B.n325 VSUBS 0.007899f
C381 B.n326 VSUBS 0.007899f
C382 B.n327 VSUBS 0.007899f
C383 B.n328 VSUBS 0.007899f
C384 B.n329 VSUBS 0.007899f
C385 B.n330 VSUBS 0.007899f
C386 B.n331 VSUBS 0.007899f
C387 B.n332 VSUBS 0.007899f
C388 B.n333 VSUBS 0.007899f
C389 B.n334 VSUBS 0.007899f
C390 B.n335 VSUBS 0.007899f
C391 B.n336 VSUBS 0.007899f
C392 B.n337 VSUBS 0.007899f
C393 B.n338 VSUBS 0.007899f
C394 B.n339 VSUBS 0.007899f
C395 B.n340 VSUBS 0.007899f
C396 B.n341 VSUBS 0.007899f
C397 B.n342 VSUBS 0.007899f
C398 B.n343 VSUBS 0.017886f
C399 VTAIL.n0 VSUBS 0.01443f
C400 VTAIL.n1 VSUBS 0.01435f
C401 VTAIL.n2 VSUBS 0.007711f
C402 VTAIL.n3 VSUBS 0.013669f
C403 VTAIL.n4 VSUBS 0.011252f
C404 VTAIL.t7 VSUBS 0.039803f
C405 VTAIL.n5 VSUBS 0.050766f
C406 VTAIL.n6 VSUBS 0.138117f
C407 VTAIL.n7 VSUBS 0.007711f
C408 VTAIL.n8 VSUBS 0.008164f
C409 VTAIL.n9 VSUBS 0.018226f
C410 VTAIL.n10 VSUBS 0.039567f
C411 VTAIL.n11 VSUBS 0.008164f
C412 VTAIL.n12 VSUBS 0.007711f
C413 VTAIL.n13 VSUBS 0.032188f
C414 VTAIL.n14 VSUBS 0.019665f
C415 VTAIL.n15 VSUBS 0.065215f
C416 VTAIL.n16 VSUBS 0.01443f
C417 VTAIL.n17 VSUBS 0.01435f
C418 VTAIL.n18 VSUBS 0.007711f
C419 VTAIL.n19 VSUBS 0.013669f
C420 VTAIL.n20 VSUBS 0.011252f
C421 VTAIL.t3 VSUBS 0.039803f
C422 VTAIL.n21 VSUBS 0.050766f
C423 VTAIL.n22 VSUBS 0.138117f
C424 VTAIL.n23 VSUBS 0.007711f
C425 VTAIL.n24 VSUBS 0.008164f
C426 VTAIL.n25 VSUBS 0.018226f
C427 VTAIL.n26 VSUBS 0.039567f
C428 VTAIL.n27 VSUBS 0.008164f
C429 VTAIL.n28 VSUBS 0.007711f
C430 VTAIL.n29 VSUBS 0.032188f
C431 VTAIL.n30 VSUBS 0.019665f
C432 VTAIL.n31 VSUBS 0.091622f
C433 VTAIL.n32 VSUBS 0.01443f
C434 VTAIL.n33 VSUBS 0.01435f
C435 VTAIL.n34 VSUBS 0.007711f
C436 VTAIL.n35 VSUBS 0.013669f
C437 VTAIL.n36 VSUBS 0.011252f
C438 VTAIL.t0 VSUBS 0.039803f
C439 VTAIL.n37 VSUBS 0.050766f
C440 VTAIL.n38 VSUBS 0.138117f
C441 VTAIL.n39 VSUBS 0.007711f
C442 VTAIL.n40 VSUBS 0.008164f
C443 VTAIL.n41 VSUBS 0.018226f
C444 VTAIL.n42 VSUBS 0.039567f
C445 VTAIL.n43 VSUBS 0.008164f
C446 VTAIL.n44 VSUBS 0.007711f
C447 VTAIL.n45 VSUBS 0.032188f
C448 VTAIL.n46 VSUBS 0.019665f
C449 VTAIL.n47 VSUBS 0.445389f
C450 VTAIL.n48 VSUBS 0.01443f
C451 VTAIL.n49 VSUBS 0.01435f
C452 VTAIL.n50 VSUBS 0.007711f
C453 VTAIL.n51 VSUBS 0.013669f
C454 VTAIL.n52 VSUBS 0.011252f
C455 VTAIL.t6 VSUBS 0.039803f
C456 VTAIL.n53 VSUBS 0.050766f
C457 VTAIL.n54 VSUBS 0.138117f
C458 VTAIL.n55 VSUBS 0.007711f
C459 VTAIL.n56 VSUBS 0.008164f
C460 VTAIL.n57 VSUBS 0.018226f
C461 VTAIL.n58 VSUBS 0.039567f
C462 VTAIL.n59 VSUBS 0.008164f
C463 VTAIL.n60 VSUBS 0.007711f
C464 VTAIL.n61 VSUBS 0.032188f
C465 VTAIL.n62 VSUBS 0.019665f
C466 VTAIL.n63 VSUBS 0.445389f
C467 VTAIL.n64 VSUBS 0.01443f
C468 VTAIL.n65 VSUBS 0.01435f
C469 VTAIL.n66 VSUBS 0.007711f
C470 VTAIL.n67 VSUBS 0.013669f
C471 VTAIL.n68 VSUBS 0.011252f
C472 VTAIL.t5 VSUBS 0.039803f
C473 VTAIL.n69 VSUBS 0.050766f
C474 VTAIL.n70 VSUBS 0.138117f
C475 VTAIL.n71 VSUBS 0.007711f
C476 VTAIL.n72 VSUBS 0.008164f
C477 VTAIL.n73 VSUBS 0.018226f
C478 VTAIL.n74 VSUBS 0.039567f
C479 VTAIL.n75 VSUBS 0.008164f
C480 VTAIL.n76 VSUBS 0.007711f
C481 VTAIL.n77 VSUBS 0.032188f
C482 VTAIL.n78 VSUBS 0.019665f
C483 VTAIL.n79 VSUBS 0.091622f
C484 VTAIL.n80 VSUBS 0.01443f
C485 VTAIL.n81 VSUBS 0.01435f
C486 VTAIL.n82 VSUBS 0.007711f
C487 VTAIL.n83 VSUBS 0.013669f
C488 VTAIL.n84 VSUBS 0.011252f
C489 VTAIL.t1 VSUBS 0.039803f
C490 VTAIL.n85 VSUBS 0.050766f
C491 VTAIL.n86 VSUBS 0.138117f
C492 VTAIL.n87 VSUBS 0.007711f
C493 VTAIL.n88 VSUBS 0.008164f
C494 VTAIL.n89 VSUBS 0.018226f
C495 VTAIL.n90 VSUBS 0.039567f
C496 VTAIL.n91 VSUBS 0.008164f
C497 VTAIL.n92 VSUBS 0.007711f
C498 VTAIL.n93 VSUBS 0.032188f
C499 VTAIL.n94 VSUBS 0.019665f
C500 VTAIL.n95 VSUBS 0.091622f
C501 VTAIL.n96 VSUBS 0.01443f
C502 VTAIL.n97 VSUBS 0.01435f
C503 VTAIL.n98 VSUBS 0.007711f
C504 VTAIL.n99 VSUBS 0.013669f
C505 VTAIL.n100 VSUBS 0.011252f
C506 VTAIL.t2 VSUBS 0.039803f
C507 VTAIL.n101 VSUBS 0.050766f
C508 VTAIL.n102 VSUBS 0.138117f
C509 VTAIL.n103 VSUBS 0.007711f
C510 VTAIL.n104 VSUBS 0.008164f
C511 VTAIL.n105 VSUBS 0.018226f
C512 VTAIL.n106 VSUBS 0.039567f
C513 VTAIL.n107 VSUBS 0.008164f
C514 VTAIL.n108 VSUBS 0.007711f
C515 VTAIL.n109 VSUBS 0.032188f
C516 VTAIL.n110 VSUBS 0.019665f
C517 VTAIL.n111 VSUBS 0.445389f
C518 VTAIL.n112 VSUBS 0.01443f
C519 VTAIL.n113 VSUBS 0.01435f
C520 VTAIL.n114 VSUBS 0.007711f
C521 VTAIL.n115 VSUBS 0.013669f
C522 VTAIL.n116 VSUBS 0.011252f
C523 VTAIL.t4 VSUBS 0.039803f
C524 VTAIL.n117 VSUBS 0.050766f
C525 VTAIL.n118 VSUBS 0.138117f
C526 VTAIL.n119 VSUBS 0.007711f
C527 VTAIL.n120 VSUBS 0.008164f
C528 VTAIL.n121 VSUBS 0.018226f
C529 VTAIL.n122 VSUBS 0.039567f
C530 VTAIL.n123 VSUBS 0.008164f
C531 VTAIL.n124 VSUBS 0.007711f
C532 VTAIL.n125 VSUBS 0.032188f
C533 VTAIL.n126 VSUBS 0.019665f
C534 VTAIL.n127 VSUBS 0.4136f
C535 VDD2.t3 VSUBS 0.045913f
C536 VDD2.t1 VSUBS 0.045913f
C537 VDD2.n0 VSUBS 0.397143f
C538 VDD2.t2 VSUBS 0.045913f
C539 VDD2.t0 VSUBS 0.045913f
C540 VDD2.n1 VSUBS 0.244643f
C541 VDD2.n2 VSUBS 1.89374f
C542 VN.t0 VSUBS 0.522815f
C543 VN.t3 VSUBS 0.522565f
C544 VN.n0 VSUBS 0.462492f
C545 VN.t2 VSUBS 0.522815f
C546 VN.t1 VSUBS 0.522565f
C547 VN.n1 VSUBS 1.29567f
.ends

