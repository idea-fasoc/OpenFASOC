* NGSPICE file created from diff_pair_sample_0332.ext - technology: sky130A

.subckt diff_pair_sample_0332 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=0 ps=0 w=13.87 l=0.24
X1 VTAIL.t15 VN.t0 VDD2.t3 B.t20 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=2.28855 ps=14.2 w=13.87 l=0.24
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=0 ps=0 w=13.87 l=0.24
X3 VTAIL.t14 VN.t1 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=2.28855 ps=14.2 w=13.87 l=0.24
X4 VTAIL.t13 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=0 ps=0 w=13.87 l=0.24
X6 VDD1.t7 VP.t0 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=5.4093 ps=28.52 w=13.87 l=0.24
X7 VDD1.t6 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X8 VDD2.t5 VN.t3 VTAIL.t12 B.t21 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=5.4093 ps=28.52 w=13.87 l=0.24
X9 VTAIL.t4 VP.t2 VDD1.t5 B.t20 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=2.28855 ps=14.2 w=13.87 l=0.24
X10 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X11 VDD1.t3 VP.t4 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=5.4093 ps=28.52 w=13.87 l=0.24
X12 VDD2.t1 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=5.4093 ps=28.52 w=13.87 l=0.24
X13 VDD2.t2 VN.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X14 VTAIL.t1 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X15 VTAIL.t9 VN.t6 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X16 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=0 ps=0 w=13.87 l=0.24
X17 VTAIL.t3 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=5.4093 pd=28.52 as=2.28855 ps=14.2 w=13.87 l=0.24
X18 VDD2.t4 VN.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
X19 VDD1.t0 VP.t7 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.28855 pd=14.2 as=2.28855 ps=14.2 w=13.87 l=0.24
R0 B.n61 B.t10 1619.09
R1 B.n68 B.t6 1619.09
R2 B.n147 B.t13 1619.09
R3 B.n156 B.t17 1619.09
R4 B.n458 B.n457 585
R5 B.n460 B.n92 585
R6 B.n463 B.n462 585
R7 B.n464 B.n91 585
R8 B.n466 B.n465 585
R9 B.n468 B.n90 585
R10 B.n471 B.n470 585
R11 B.n472 B.n89 585
R12 B.n474 B.n473 585
R13 B.n476 B.n88 585
R14 B.n479 B.n478 585
R15 B.n480 B.n87 585
R16 B.n482 B.n481 585
R17 B.n484 B.n86 585
R18 B.n487 B.n486 585
R19 B.n488 B.n85 585
R20 B.n490 B.n489 585
R21 B.n492 B.n84 585
R22 B.n495 B.n494 585
R23 B.n496 B.n83 585
R24 B.n498 B.n497 585
R25 B.n500 B.n82 585
R26 B.n503 B.n502 585
R27 B.n504 B.n81 585
R28 B.n506 B.n505 585
R29 B.n508 B.n80 585
R30 B.n511 B.n510 585
R31 B.n512 B.n79 585
R32 B.n514 B.n513 585
R33 B.n516 B.n78 585
R34 B.n519 B.n518 585
R35 B.n520 B.n77 585
R36 B.n522 B.n521 585
R37 B.n524 B.n76 585
R38 B.n527 B.n526 585
R39 B.n528 B.n75 585
R40 B.n530 B.n529 585
R41 B.n532 B.n74 585
R42 B.n535 B.n534 585
R43 B.n536 B.n73 585
R44 B.n538 B.n537 585
R45 B.n540 B.n72 585
R46 B.n543 B.n542 585
R47 B.n544 B.n71 585
R48 B.n546 B.n545 585
R49 B.n548 B.n70 585
R50 B.n551 B.n550 585
R51 B.n553 B.n67 585
R52 B.n555 B.n554 585
R53 B.n557 B.n66 585
R54 B.n560 B.n559 585
R55 B.n561 B.n65 585
R56 B.n563 B.n562 585
R57 B.n565 B.n64 585
R58 B.n568 B.n567 585
R59 B.n569 B.n60 585
R60 B.n571 B.n570 585
R61 B.n573 B.n59 585
R62 B.n576 B.n575 585
R63 B.n577 B.n58 585
R64 B.n579 B.n578 585
R65 B.n581 B.n57 585
R66 B.n584 B.n583 585
R67 B.n585 B.n56 585
R68 B.n587 B.n586 585
R69 B.n589 B.n55 585
R70 B.n592 B.n591 585
R71 B.n593 B.n54 585
R72 B.n595 B.n594 585
R73 B.n597 B.n53 585
R74 B.n600 B.n599 585
R75 B.n601 B.n52 585
R76 B.n603 B.n602 585
R77 B.n605 B.n51 585
R78 B.n608 B.n607 585
R79 B.n609 B.n50 585
R80 B.n611 B.n610 585
R81 B.n613 B.n49 585
R82 B.n616 B.n615 585
R83 B.n617 B.n48 585
R84 B.n619 B.n618 585
R85 B.n621 B.n47 585
R86 B.n624 B.n623 585
R87 B.n625 B.n46 585
R88 B.n627 B.n626 585
R89 B.n629 B.n45 585
R90 B.n632 B.n631 585
R91 B.n633 B.n44 585
R92 B.n635 B.n634 585
R93 B.n637 B.n43 585
R94 B.n640 B.n639 585
R95 B.n641 B.n42 585
R96 B.n643 B.n642 585
R97 B.n645 B.n41 585
R98 B.n648 B.n647 585
R99 B.n649 B.n40 585
R100 B.n651 B.n650 585
R101 B.n653 B.n39 585
R102 B.n656 B.n655 585
R103 B.n657 B.n38 585
R104 B.n659 B.n658 585
R105 B.n661 B.n37 585
R106 B.n664 B.n663 585
R107 B.n665 B.n36 585
R108 B.n456 B.n34 585
R109 B.n668 B.n34 585
R110 B.n455 B.n33 585
R111 B.n669 B.n33 585
R112 B.n454 B.n32 585
R113 B.n670 B.n32 585
R114 B.n453 B.n452 585
R115 B.n452 B.n28 585
R116 B.n451 B.n27 585
R117 B.n676 B.n27 585
R118 B.n450 B.n26 585
R119 B.n677 B.n26 585
R120 B.n449 B.n25 585
R121 B.n678 B.n25 585
R122 B.n448 B.n447 585
R123 B.n447 B.n21 585
R124 B.n446 B.n20 585
R125 B.n684 B.n20 585
R126 B.n445 B.n19 585
R127 B.n685 B.n19 585
R128 B.n444 B.n18 585
R129 B.n686 B.n18 585
R130 B.n443 B.n442 585
R131 B.n442 B.n13 585
R132 B.n441 B.n12 585
R133 B.n692 B.n12 585
R134 B.n440 B.n11 585
R135 B.n693 B.n11 585
R136 B.n439 B.n10 585
R137 B.n694 B.n10 585
R138 B.n438 B.n7 585
R139 B.n697 B.n7 585
R140 B.n437 B.n6 585
R141 B.n698 B.n6 585
R142 B.n436 B.n5 585
R143 B.n699 B.n5 585
R144 B.n435 B.n434 585
R145 B.n434 B.n4 585
R146 B.n433 B.n93 585
R147 B.n433 B.n432 585
R148 B.n423 B.n94 585
R149 B.n95 B.n94 585
R150 B.n425 B.n424 585
R151 B.n426 B.n425 585
R152 B.n422 B.n100 585
R153 B.n100 B.n99 585
R154 B.n421 B.n420 585
R155 B.n420 B.n419 585
R156 B.n102 B.n101 585
R157 B.n412 B.n102 585
R158 B.n411 B.n410 585
R159 B.n413 B.n411 585
R160 B.n409 B.n107 585
R161 B.n107 B.n106 585
R162 B.n408 B.n407 585
R163 B.n407 B.n406 585
R164 B.n109 B.n108 585
R165 B.n110 B.n109 585
R166 B.n399 B.n398 585
R167 B.n400 B.n399 585
R168 B.n397 B.n115 585
R169 B.n115 B.n114 585
R170 B.n396 B.n395 585
R171 B.n395 B.n394 585
R172 B.n117 B.n116 585
R173 B.n118 B.n117 585
R174 B.n387 B.n386 585
R175 B.n388 B.n387 585
R176 B.n121 B.n120 585
R177 B.n182 B.n181 585
R178 B.n183 B.n179 585
R179 B.n179 B.n122 585
R180 B.n185 B.n184 585
R181 B.n187 B.n178 585
R182 B.n190 B.n189 585
R183 B.n191 B.n177 585
R184 B.n193 B.n192 585
R185 B.n195 B.n176 585
R186 B.n198 B.n197 585
R187 B.n199 B.n175 585
R188 B.n201 B.n200 585
R189 B.n203 B.n174 585
R190 B.n206 B.n205 585
R191 B.n207 B.n173 585
R192 B.n209 B.n208 585
R193 B.n211 B.n172 585
R194 B.n214 B.n213 585
R195 B.n215 B.n171 585
R196 B.n217 B.n216 585
R197 B.n219 B.n170 585
R198 B.n222 B.n221 585
R199 B.n223 B.n169 585
R200 B.n225 B.n224 585
R201 B.n227 B.n168 585
R202 B.n230 B.n229 585
R203 B.n231 B.n167 585
R204 B.n233 B.n232 585
R205 B.n235 B.n166 585
R206 B.n238 B.n237 585
R207 B.n239 B.n165 585
R208 B.n241 B.n240 585
R209 B.n243 B.n164 585
R210 B.n246 B.n245 585
R211 B.n247 B.n163 585
R212 B.n249 B.n248 585
R213 B.n251 B.n162 585
R214 B.n254 B.n253 585
R215 B.n255 B.n161 585
R216 B.n257 B.n256 585
R217 B.n259 B.n160 585
R218 B.n262 B.n261 585
R219 B.n263 B.n159 585
R220 B.n265 B.n264 585
R221 B.n267 B.n158 585
R222 B.n270 B.n269 585
R223 B.n271 B.n155 585
R224 B.n274 B.n273 585
R225 B.n276 B.n154 585
R226 B.n279 B.n278 585
R227 B.n280 B.n153 585
R228 B.n282 B.n281 585
R229 B.n284 B.n152 585
R230 B.n287 B.n286 585
R231 B.n288 B.n151 585
R232 B.n290 B.n289 585
R233 B.n292 B.n150 585
R234 B.n295 B.n294 585
R235 B.n296 B.n146 585
R236 B.n298 B.n297 585
R237 B.n300 B.n145 585
R238 B.n303 B.n302 585
R239 B.n304 B.n144 585
R240 B.n306 B.n305 585
R241 B.n308 B.n143 585
R242 B.n311 B.n310 585
R243 B.n312 B.n142 585
R244 B.n314 B.n313 585
R245 B.n316 B.n141 585
R246 B.n319 B.n318 585
R247 B.n320 B.n140 585
R248 B.n322 B.n321 585
R249 B.n324 B.n139 585
R250 B.n327 B.n326 585
R251 B.n328 B.n138 585
R252 B.n330 B.n329 585
R253 B.n332 B.n137 585
R254 B.n335 B.n334 585
R255 B.n336 B.n136 585
R256 B.n338 B.n337 585
R257 B.n340 B.n135 585
R258 B.n343 B.n342 585
R259 B.n344 B.n134 585
R260 B.n346 B.n345 585
R261 B.n348 B.n133 585
R262 B.n351 B.n350 585
R263 B.n352 B.n132 585
R264 B.n354 B.n353 585
R265 B.n356 B.n131 585
R266 B.n359 B.n358 585
R267 B.n360 B.n130 585
R268 B.n362 B.n361 585
R269 B.n364 B.n129 585
R270 B.n367 B.n366 585
R271 B.n368 B.n128 585
R272 B.n370 B.n369 585
R273 B.n372 B.n127 585
R274 B.n375 B.n374 585
R275 B.n376 B.n126 585
R276 B.n378 B.n377 585
R277 B.n380 B.n125 585
R278 B.n381 B.n124 585
R279 B.n384 B.n383 585
R280 B.n385 B.n123 585
R281 B.n123 B.n122 585
R282 B.n390 B.n389 585
R283 B.n389 B.n388 585
R284 B.n391 B.n119 585
R285 B.n119 B.n118 585
R286 B.n393 B.n392 585
R287 B.n394 B.n393 585
R288 B.n113 B.n112 585
R289 B.n114 B.n113 585
R290 B.n402 B.n401 585
R291 B.n401 B.n400 585
R292 B.n403 B.n111 585
R293 B.n111 B.n110 585
R294 B.n405 B.n404 585
R295 B.n406 B.n405 585
R296 B.n105 B.n104 585
R297 B.n106 B.n105 585
R298 B.n415 B.n414 585
R299 B.n414 B.n413 585
R300 B.n416 B.n103 585
R301 B.n412 B.n103 585
R302 B.n418 B.n417 585
R303 B.n419 B.n418 585
R304 B.n98 B.n97 585
R305 B.n99 B.n98 585
R306 B.n428 B.n427 585
R307 B.n427 B.n426 585
R308 B.n429 B.n96 585
R309 B.n96 B.n95 585
R310 B.n431 B.n430 585
R311 B.n432 B.n431 585
R312 B.n3 B.n0 585
R313 B.n4 B.n3 585
R314 B.n696 B.n1 585
R315 B.n697 B.n696 585
R316 B.n695 B.n9 585
R317 B.n695 B.n694 585
R318 B.n15 B.n8 585
R319 B.n693 B.n8 585
R320 B.n691 B.n690 585
R321 B.n692 B.n691 585
R322 B.n689 B.n14 585
R323 B.n14 B.n13 585
R324 B.n688 B.n687 585
R325 B.n687 B.n686 585
R326 B.n17 B.n16 585
R327 B.n685 B.n17 585
R328 B.n683 B.n682 585
R329 B.n684 B.n683 585
R330 B.n681 B.n22 585
R331 B.n22 B.n21 585
R332 B.n680 B.n679 585
R333 B.n679 B.n678 585
R334 B.n24 B.n23 585
R335 B.n677 B.n24 585
R336 B.n675 B.n674 585
R337 B.n676 B.n675 585
R338 B.n673 B.n29 585
R339 B.n29 B.n28 585
R340 B.n672 B.n671 585
R341 B.n671 B.n670 585
R342 B.n31 B.n30 585
R343 B.n669 B.n31 585
R344 B.n667 B.n666 585
R345 B.n668 B.n667 585
R346 B.n700 B.n699 585
R347 B.n698 B.n2 585
R348 B.n667 B.n36 482.89
R349 B.n458 B.n34 482.89
R350 B.n387 B.n123 482.89
R351 B.n389 B.n121 482.89
R352 B.n459 B.n35 256.663
R353 B.n461 B.n35 256.663
R354 B.n467 B.n35 256.663
R355 B.n469 B.n35 256.663
R356 B.n475 B.n35 256.663
R357 B.n477 B.n35 256.663
R358 B.n483 B.n35 256.663
R359 B.n485 B.n35 256.663
R360 B.n491 B.n35 256.663
R361 B.n493 B.n35 256.663
R362 B.n499 B.n35 256.663
R363 B.n501 B.n35 256.663
R364 B.n507 B.n35 256.663
R365 B.n509 B.n35 256.663
R366 B.n515 B.n35 256.663
R367 B.n517 B.n35 256.663
R368 B.n523 B.n35 256.663
R369 B.n525 B.n35 256.663
R370 B.n531 B.n35 256.663
R371 B.n533 B.n35 256.663
R372 B.n539 B.n35 256.663
R373 B.n541 B.n35 256.663
R374 B.n547 B.n35 256.663
R375 B.n549 B.n35 256.663
R376 B.n556 B.n35 256.663
R377 B.n558 B.n35 256.663
R378 B.n564 B.n35 256.663
R379 B.n566 B.n35 256.663
R380 B.n572 B.n35 256.663
R381 B.n574 B.n35 256.663
R382 B.n580 B.n35 256.663
R383 B.n582 B.n35 256.663
R384 B.n588 B.n35 256.663
R385 B.n590 B.n35 256.663
R386 B.n596 B.n35 256.663
R387 B.n598 B.n35 256.663
R388 B.n604 B.n35 256.663
R389 B.n606 B.n35 256.663
R390 B.n612 B.n35 256.663
R391 B.n614 B.n35 256.663
R392 B.n620 B.n35 256.663
R393 B.n622 B.n35 256.663
R394 B.n628 B.n35 256.663
R395 B.n630 B.n35 256.663
R396 B.n636 B.n35 256.663
R397 B.n638 B.n35 256.663
R398 B.n644 B.n35 256.663
R399 B.n646 B.n35 256.663
R400 B.n652 B.n35 256.663
R401 B.n654 B.n35 256.663
R402 B.n660 B.n35 256.663
R403 B.n662 B.n35 256.663
R404 B.n180 B.n122 256.663
R405 B.n186 B.n122 256.663
R406 B.n188 B.n122 256.663
R407 B.n194 B.n122 256.663
R408 B.n196 B.n122 256.663
R409 B.n202 B.n122 256.663
R410 B.n204 B.n122 256.663
R411 B.n210 B.n122 256.663
R412 B.n212 B.n122 256.663
R413 B.n218 B.n122 256.663
R414 B.n220 B.n122 256.663
R415 B.n226 B.n122 256.663
R416 B.n228 B.n122 256.663
R417 B.n234 B.n122 256.663
R418 B.n236 B.n122 256.663
R419 B.n242 B.n122 256.663
R420 B.n244 B.n122 256.663
R421 B.n250 B.n122 256.663
R422 B.n252 B.n122 256.663
R423 B.n258 B.n122 256.663
R424 B.n260 B.n122 256.663
R425 B.n266 B.n122 256.663
R426 B.n268 B.n122 256.663
R427 B.n275 B.n122 256.663
R428 B.n277 B.n122 256.663
R429 B.n283 B.n122 256.663
R430 B.n285 B.n122 256.663
R431 B.n291 B.n122 256.663
R432 B.n293 B.n122 256.663
R433 B.n299 B.n122 256.663
R434 B.n301 B.n122 256.663
R435 B.n307 B.n122 256.663
R436 B.n309 B.n122 256.663
R437 B.n315 B.n122 256.663
R438 B.n317 B.n122 256.663
R439 B.n323 B.n122 256.663
R440 B.n325 B.n122 256.663
R441 B.n331 B.n122 256.663
R442 B.n333 B.n122 256.663
R443 B.n339 B.n122 256.663
R444 B.n341 B.n122 256.663
R445 B.n347 B.n122 256.663
R446 B.n349 B.n122 256.663
R447 B.n355 B.n122 256.663
R448 B.n357 B.n122 256.663
R449 B.n363 B.n122 256.663
R450 B.n365 B.n122 256.663
R451 B.n371 B.n122 256.663
R452 B.n373 B.n122 256.663
R453 B.n379 B.n122 256.663
R454 B.n382 B.n122 256.663
R455 B.n702 B.n701 256.663
R456 B.n663 B.n661 163.367
R457 B.n659 B.n38 163.367
R458 B.n655 B.n653 163.367
R459 B.n651 B.n40 163.367
R460 B.n647 B.n645 163.367
R461 B.n643 B.n42 163.367
R462 B.n639 B.n637 163.367
R463 B.n635 B.n44 163.367
R464 B.n631 B.n629 163.367
R465 B.n627 B.n46 163.367
R466 B.n623 B.n621 163.367
R467 B.n619 B.n48 163.367
R468 B.n615 B.n613 163.367
R469 B.n611 B.n50 163.367
R470 B.n607 B.n605 163.367
R471 B.n603 B.n52 163.367
R472 B.n599 B.n597 163.367
R473 B.n595 B.n54 163.367
R474 B.n591 B.n589 163.367
R475 B.n587 B.n56 163.367
R476 B.n583 B.n581 163.367
R477 B.n579 B.n58 163.367
R478 B.n575 B.n573 163.367
R479 B.n571 B.n60 163.367
R480 B.n567 B.n565 163.367
R481 B.n563 B.n65 163.367
R482 B.n559 B.n557 163.367
R483 B.n555 B.n67 163.367
R484 B.n550 B.n548 163.367
R485 B.n546 B.n71 163.367
R486 B.n542 B.n540 163.367
R487 B.n538 B.n73 163.367
R488 B.n534 B.n532 163.367
R489 B.n530 B.n75 163.367
R490 B.n526 B.n524 163.367
R491 B.n522 B.n77 163.367
R492 B.n518 B.n516 163.367
R493 B.n514 B.n79 163.367
R494 B.n510 B.n508 163.367
R495 B.n506 B.n81 163.367
R496 B.n502 B.n500 163.367
R497 B.n498 B.n83 163.367
R498 B.n494 B.n492 163.367
R499 B.n490 B.n85 163.367
R500 B.n486 B.n484 163.367
R501 B.n482 B.n87 163.367
R502 B.n478 B.n476 163.367
R503 B.n474 B.n89 163.367
R504 B.n470 B.n468 163.367
R505 B.n466 B.n91 163.367
R506 B.n462 B.n460 163.367
R507 B.n387 B.n117 163.367
R508 B.n395 B.n117 163.367
R509 B.n395 B.n115 163.367
R510 B.n399 B.n115 163.367
R511 B.n399 B.n109 163.367
R512 B.n407 B.n109 163.367
R513 B.n407 B.n107 163.367
R514 B.n411 B.n107 163.367
R515 B.n411 B.n102 163.367
R516 B.n420 B.n102 163.367
R517 B.n420 B.n100 163.367
R518 B.n425 B.n100 163.367
R519 B.n425 B.n94 163.367
R520 B.n433 B.n94 163.367
R521 B.n434 B.n433 163.367
R522 B.n434 B.n5 163.367
R523 B.n6 B.n5 163.367
R524 B.n7 B.n6 163.367
R525 B.n10 B.n7 163.367
R526 B.n11 B.n10 163.367
R527 B.n12 B.n11 163.367
R528 B.n442 B.n12 163.367
R529 B.n442 B.n18 163.367
R530 B.n19 B.n18 163.367
R531 B.n20 B.n19 163.367
R532 B.n447 B.n20 163.367
R533 B.n447 B.n25 163.367
R534 B.n26 B.n25 163.367
R535 B.n27 B.n26 163.367
R536 B.n452 B.n27 163.367
R537 B.n452 B.n32 163.367
R538 B.n33 B.n32 163.367
R539 B.n34 B.n33 163.367
R540 B.n181 B.n179 163.367
R541 B.n185 B.n179 163.367
R542 B.n189 B.n187 163.367
R543 B.n193 B.n177 163.367
R544 B.n197 B.n195 163.367
R545 B.n201 B.n175 163.367
R546 B.n205 B.n203 163.367
R547 B.n209 B.n173 163.367
R548 B.n213 B.n211 163.367
R549 B.n217 B.n171 163.367
R550 B.n221 B.n219 163.367
R551 B.n225 B.n169 163.367
R552 B.n229 B.n227 163.367
R553 B.n233 B.n167 163.367
R554 B.n237 B.n235 163.367
R555 B.n241 B.n165 163.367
R556 B.n245 B.n243 163.367
R557 B.n249 B.n163 163.367
R558 B.n253 B.n251 163.367
R559 B.n257 B.n161 163.367
R560 B.n261 B.n259 163.367
R561 B.n265 B.n159 163.367
R562 B.n269 B.n267 163.367
R563 B.n274 B.n155 163.367
R564 B.n278 B.n276 163.367
R565 B.n282 B.n153 163.367
R566 B.n286 B.n284 163.367
R567 B.n290 B.n151 163.367
R568 B.n294 B.n292 163.367
R569 B.n298 B.n146 163.367
R570 B.n302 B.n300 163.367
R571 B.n306 B.n144 163.367
R572 B.n310 B.n308 163.367
R573 B.n314 B.n142 163.367
R574 B.n318 B.n316 163.367
R575 B.n322 B.n140 163.367
R576 B.n326 B.n324 163.367
R577 B.n330 B.n138 163.367
R578 B.n334 B.n332 163.367
R579 B.n338 B.n136 163.367
R580 B.n342 B.n340 163.367
R581 B.n346 B.n134 163.367
R582 B.n350 B.n348 163.367
R583 B.n354 B.n132 163.367
R584 B.n358 B.n356 163.367
R585 B.n362 B.n130 163.367
R586 B.n366 B.n364 163.367
R587 B.n370 B.n128 163.367
R588 B.n374 B.n372 163.367
R589 B.n378 B.n126 163.367
R590 B.n381 B.n380 163.367
R591 B.n383 B.n123 163.367
R592 B.n389 B.n119 163.367
R593 B.n393 B.n119 163.367
R594 B.n393 B.n113 163.367
R595 B.n401 B.n113 163.367
R596 B.n401 B.n111 163.367
R597 B.n405 B.n111 163.367
R598 B.n405 B.n105 163.367
R599 B.n414 B.n105 163.367
R600 B.n414 B.n103 163.367
R601 B.n418 B.n103 163.367
R602 B.n418 B.n98 163.367
R603 B.n427 B.n98 163.367
R604 B.n427 B.n96 163.367
R605 B.n431 B.n96 163.367
R606 B.n431 B.n3 163.367
R607 B.n700 B.n3 163.367
R608 B.n696 B.n2 163.367
R609 B.n696 B.n695 163.367
R610 B.n695 B.n8 163.367
R611 B.n691 B.n8 163.367
R612 B.n691 B.n14 163.367
R613 B.n687 B.n14 163.367
R614 B.n687 B.n17 163.367
R615 B.n683 B.n17 163.367
R616 B.n683 B.n22 163.367
R617 B.n679 B.n22 163.367
R618 B.n679 B.n24 163.367
R619 B.n675 B.n24 163.367
R620 B.n675 B.n29 163.367
R621 B.n671 B.n29 163.367
R622 B.n671 B.n31 163.367
R623 B.n667 B.n31 163.367
R624 B.n68 B.t8 83.8608
R625 B.n147 B.t16 83.8608
R626 B.n61 B.t11 83.8431
R627 B.n156 B.t19 83.8431
R628 B.n69 B.t9 72.8063
R629 B.n148 B.t15 72.8063
R630 B.n62 B.t12 72.7886
R631 B.n157 B.t18 72.7886
R632 B.n662 B.n36 71.676
R633 B.n661 B.n660 71.676
R634 B.n654 B.n38 71.676
R635 B.n653 B.n652 71.676
R636 B.n646 B.n40 71.676
R637 B.n645 B.n644 71.676
R638 B.n638 B.n42 71.676
R639 B.n637 B.n636 71.676
R640 B.n630 B.n44 71.676
R641 B.n629 B.n628 71.676
R642 B.n622 B.n46 71.676
R643 B.n621 B.n620 71.676
R644 B.n614 B.n48 71.676
R645 B.n613 B.n612 71.676
R646 B.n606 B.n50 71.676
R647 B.n605 B.n604 71.676
R648 B.n598 B.n52 71.676
R649 B.n597 B.n596 71.676
R650 B.n590 B.n54 71.676
R651 B.n589 B.n588 71.676
R652 B.n582 B.n56 71.676
R653 B.n581 B.n580 71.676
R654 B.n574 B.n58 71.676
R655 B.n573 B.n572 71.676
R656 B.n566 B.n60 71.676
R657 B.n565 B.n564 71.676
R658 B.n558 B.n65 71.676
R659 B.n557 B.n556 71.676
R660 B.n549 B.n67 71.676
R661 B.n548 B.n547 71.676
R662 B.n541 B.n71 71.676
R663 B.n540 B.n539 71.676
R664 B.n533 B.n73 71.676
R665 B.n532 B.n531 71.676
R666 B.n525 B.n75 71.676
R667 B.n524 B.n523 71.676
R668 B.n517 B.n77 71.676
R669 B.n516 B.n515 71.676
R670 B.n509 B.n79 71.676
R671 B.n508 B.n507 71.676
R672 B.n501 B.n81 71.676
R673 B.n500 B.n499 71.676
R674 B.n493 B.n83 71.676
R675 B.n492 B.n491 71.676
R676 B.n485 B.n85 71.676
R677 B.n484 B.n483 71.676
R678 B.n477 B.n87 71.676
R679 B.n476 B.n475 71.676
R680 B.n469 B.n89 71.676
R681 B.n468 B.n467 71.676
R682 B.n461 B.n91 71.676
R683 B.n460 B.n459 71.676
R684 B.n459 B.n458 71.676
R685 B.n462 B.n461 71.676
R686 B.n467 B.n466 71.676
R687 B.n470 B.n469 71.676
R688 B.n475 B.n474 71.676
R689 B.n478 B.n477 71.676
R690 B.n483 B.n482 71.676
R691 B.n486 B.n485 71.676
R692 B.n491 B.n490 71.676
R693 B.n494 B.n493 71.676
R694 B.n499 B.n498 71.676
R695 B.n502 B.n501 71.676
R696 B.n507 B.n506 71.676
R697 B.n510 B.n509 71.676
R698 B.n515 B.n514 71.676
R699 B.n518 B.n517 71.676
R700 B.n523 B.n522 71.676
R701 B.n526 B.n525 71.676
R702 B.n531 B.n530 71.676
R703 B.n534 B.n533 71.676
R704 B.n539 B.n538 71.676
R705 B.n542 B.n541 71.676
R706 B.n547 B.n546 71.676
R707 B.n550 B.n549 71.676
R708 B.n556 B.n555 71.676
R709 B.n559 B.n558 71.676
R710 B.n564 B.n563 71.676
R711 B.n567 B.n566 71.676
R712 B.n572 B.n571 71.676
R713 B.n575 B.n574 71.676
R714 B.n580 B.n579 71.676
R715 B.n583 B.n582 71.676
R716 B.n588 B.n587 71.676
R717 B.n591 B.n590 71.676
R718 B.n596 B.n595 71.676
R719 B.n599 B.n598 71.676
R720 B.n604 B.n603 71.676
R721 B.n607 B.n606 71.676
R722 B.n612 B.n611 71.676
R723 B.n615 B.n614 71.676
R724 B.n620 B.n619 71.676
R725 B.n623 B.n622 71.676
R726 B.n628 B.n627 71.676
R727 B.n631 B.n630 71.676
R728 B.n636 B.n635 71.676
R729 B.n639 B.n638 71.676
R730 B.n644 B.n643 71.676
R731 B.n647 B.n646 71.676
R732 B.n652 B.n651 71.676
R733 B.n655 B.n654 71.676
R734 B.n660 B.n659 71.676
R735 B.n663 B.n662 71.676
R736 B.n180 B.n121 71.676
R737 B.n186 B.n185 71.676
R738 B.n189 B.n188 71.676
R739 B.n194 B.n193 71.676
R740 B.n197 B.n196 71.676
R741 B.n202 B.n201 71.676
R742 B.n205 B.n204 71.676
R743 B.n210 B.n209 71.676
R744 B.n213 B.n212 71.676
R745 B.n218 B.n217 71.676
R746 B.n221 B.n220 71.676
R747 B.n226 B.n225 71.676
R748 B.n229 B.n228 71.676
R749 B.n234 B.n233 71.676
R750 B.n237 B.n236 71.676
R751 B.n242 B.n241 71.676
R752 B.n245 B.n244 71.676
R753 B.n250 B.n249 71.676
R754 B.n253 B.n252 71.676
R755 B.n258 B.n257 71.676
R756 B.n261 B.n260 71.676
R757 B.n266 B.n265 71.676
R758 B.n269 B.n268 71.676
R759 B.n275 B.n274 71.676
R760 B.n278 B.n277 71.676
R761 B.n283 B.n282 71.676
R762 B.n286 B.n285 71.676
R763 B.n291 B.n290 71.676
R764 B.n294 B.n293 71.676
R765 B.n299 B.n298 71.676
R766 B.n302 B.n301 71.676
R767 B.n307 B.n306 71.676
R768 B.n310 B.n309 71.676
R769 B.n315 B.n314 71.676
R770 B.n318 B.n317 71.676
R771 B.n323 B.n322 71.676
R772 B.n326 B.n325 71.676
R773 B.n331 B.n330 71.676
R774 B.n334 B.n333 71.676
R775 B.n339 B.n338 71.676
R776 B.n342 B.n341 71.676
R777 B.n347 B.n346 71.676
R778 B.n350 B.n349 71.676
R779 B.n355 B.n354 71.676
R780 B.n358 B.n357 71.676
R781 B.n363 B.n362 71.676
R782 B.n366 B.n365 71.676
R783 B.n371 B.n370 71.676
R784 B.n374 B.n373 71.676
R785 B.n379 B.n378 71.676
R786 B.n382 B.n381 71.676
R787 B.n181 B.n180 71.676
R788 B.n187 B.n186 71.676
R789 B.n188 B.n177 71.676
R790 B.n195 B.n194 71.676
R791 B.n196 B.n175 71.676
R792 B.n203 B.n202 71.676
R793 B.n204 B.n173 71.676
R794 B.n211 B.n210 71.676
R795 B.n212 B.n171 71.676
R796 B.n219 B.n218 71.676
R797 B.n220 B.n169 71.676
R798 B.n227 B.n226 71.676
R799 B.n228 B.n167 71.676
R800 B.n235 B.n234 71.676
R801 B.n236 B.n165 71.676
R802 B.n243 B.n242 71.676
R803 B.n244 B.n163 71.676
R804 B.n251 B.n250 71.676
R805 B.n252 B.n161 71.676
R806 B.n259 B.n258 71.676
R807 B.n260 B.n159 71.676
R808 B.n267 B.n266 71.676
R809 B.n268 B.n155 71.676
R810 B.n276 B.n275 71.676
R811 B.n277 B.n153 71.676
R812 B.n284 B.n283 71.676
R813 B.n285 B.n151 71.676
R814 B.n292 B.n291 71.676
R815 B.n293 B.n146 71.676
R816 B.n300 B.n299 71.676
R817 B.n301 B.n144 71.676
R818 B.n308 B.n307 71.676
R819 B.n309 B.n142 71.676
R820 B.n316 B.n315 71.676
R821 B.n317 B.n140 71.676
R822 B.n324 B.n323 71.676
R823 B.n325 B.n138 71.676
R824 B.n332 B.n331 71.676
R825 B.n333 B.n136 71.676
R826 B.n340 B.n339 71.676
R827 B.n341 B.n134 71.676
R828 B.n348 B.n347 71.676
R829 B.n349 B.n132 71.676
R830 B.n356 B.n355 71.676
R831 B.n357 B.n130 71.676
R832 B.n364 B.n363 71.676
R833 B.n365 B.n128 71.676
R834 B.n372 B.n371 71.676
R835 B.n373 B.n126 71.676
R836 B.n380 B.n379 71.676
R837 B.n383 B.n382 71.676
R838 B.n701 B.n700 71.676
R839 B.n701 B.n2 71.676
R840 B.n388 B.n122 70.6717
R841 B.n668 B.n35 70.6717
R842 B.n63 B.n62 59.5399
R843 B.n552 B.n69 59.5399
R844 B.n149 B.n148 59.5399
R845 B.n272 B.n157 59.5399
R846 B.n388 B.n118 39.0708
R847 B.n394 B.n118 39.0708
R848 B.n394 B.n114 39.0708
R849 B.n400 B.n114 39.0708
R850 B.n406 B.n110 39.0708
R851 B.n406 B.n106 39.0708
R852 B.n413 B.n106 39.0708
R853 B.n413 B.n412 39.0708
R854 B.n426 B.n99 39.0708
R855 B.n432 B.n95 39.0708
R856 B.n699 B.n4 39.0708
R857 B.n699 B.n698 39.0708
R858 B.n698 B.n697 39.0708
R859 B.n694 B.n693 39.0708
R860 B.n692 B.n13 39.0708
R861 B.n685 B.n684 39.0708
R862 B.n684 B.n21 39.0708
R863 B.n678 B.n21 39.0708
R864 B.n678 B.n677 39.0708
R865 B.n676 B.n28 39.0708
R866 B.n670 B.n28 39.0708
R867 B.n670 B.n669 39.0708
R868 B.n669 B.n668 39.0708
R869 B.n419 B.t20 37.9216
R870 B.n686 B.t21 37.9216
R871 B.t5 B.n4 36.7725
R872 B.n697 B.t4 36.7725
R873 B.t14 B.n110 33.3251
R874 B.n677 B.t7 33.3251
R875 B.n390 B.n120 31.3761
R876 B.n386 B.n385 31.3761
R877 B.n457 B.n456 31.3761
R878 B.n666 B.n665 31.3761
R879 B.n419 B.t2 27.5795
R880 B.n686 B.t0 27.5795
R881 B.t3 B.n95 24.1321
R882 B.n693 B.t1 24.1321
R883 B B.n702 18.0485
R884 B.n426 B.t3 14.9391
R885 B.t1 B.n692 14.9391
R886 B.t2 B.n99 11.4918
R887 B.t0 B.n13 11.4918
R888 B.n62 B.n61 11.055
R889 B.n69 B.n68 11.055
R890 B.n148 B.n147 11.055
R891 B.n157 B.n156 11.055
R892 B.n391 B.n390 10.6151
R893 B.n392 B.n391 10.6151
R894 B.n392 B.n112 10.6151
R895 B.n402 B.n112 10.6151
R896 B.n403 B.n402 10.6151
R897 B.n404 B.n403 10.6151
R898 B.n404 B.n104 10.6151
R899 B.n415 B.n104 10.6151
R900 B.n416 B.n415 10.6151
R901 B.n417 B.n416 10.6151
R902 B.n417 B.n97 10.6151
R903 B.n428 B.n97 10.6151
R904 B.n429 B.n428 10.6151
R905 B.n430 B.n429 10.6151
R906 B.n430 B.n0 10.6151
R907 B.n182 B.n120 10.6151
R908 B.n183 B.n182 10.6151
R909 B.n184 B.n183 10.6151
R910 B.n184 B.n178 10.6151
R911 B.n190 B.n178 10.6151
R912 B.n191 B.n190 10.6151
R913 B.n192 B.n191 10.6151
R914 B.n192 B.n176 10.6151
R915 B.n198 B.n176 10.6151
R916 B.n199 B.n198 10.6151
R917 B.n200 B.n199 10.6151
R918 B.n200 B.n174 10.6151
R919 B.n206 B.n174 10.6151
R920 B.n207 B.n206 10.6151
R921 B.n208 B.n207 10.6151
R922 B.n208 B.n172 10.6151
R923 B.n214 B.n172 10.6151
R924 B.n215 B.n214 10.6151
R925 B.n216 B.n215 10.6151
R926 B.n216 B.n170 10.6151
R927 B.n222 B.n170 10.6151
R928 B.n223 B.n222 10.6151
R929 B.n224 B.n223 10.6151
R930 B.n224 B.n168 10.6151
R931 B.n230 B.n168 10.6151
R932 B.n231 B.n230 10.6151
R933 B.n232 B.n231 10.6151
R934 B.n232 B.n166 10.6151
R935 B.n238 B.n166 10.6151
R936 B.n239 B.n238 10.6151
R937 B.n240 B.n239 10.6151
R938 B.n240 B.n164 10.6151
R939 B.n246 B.n164 10.6151
R940 B.n247 B.n246 10.6151
R941 B.n248 B.n247 10.6151
R942 B.n248 B.n162 10.6151
R943 B.n254 B.n162 10.6151
R944 B.n255 B.n254 10.6151
R945 B.n256 B.n255 10.6151
R946 B.n256 B.n160 10.6151
R947 B.n262 B.n160 10.6151
R948 B.n263 B.n262 10.6151
R949 B.n264 B.n263 10.6151
R950 B.n264 B.n158 10.6151
R951 B.n270 B.n158 10.6151
R952 B.n271 B.n270 10.6151
R953 B.n273 B.n154 10.6151
R954 B.n279 B.n154 10.6151
R955 B.n280 B.n279 10.6151
R956 B.n281 B.n280 10.6151
R957 B.n281 B.n152 10.6151
R958 B.n287 B.n152 10.6151
R959 B.n288 B.n287 10.6151
R960 B.n289 B.n288 10.6151
R961 B.n289 B.n150 10.6151
R962 B.n296 B.n295 10.6151
R963 B.n297 B.n296 10.6151
R964 B.n297 B.n145 10.6151
R965 B.n303 B.n145 10.6151
R966 B.n304 B.n303 10.6151
R967 B.n305 B.n304 10.6151
R968 B.n305 B.n143 10.6151
R969 B.n311 B.n143 10.6151
R970 B.n312 B.n311 10.6151
R971 B.n313 B.n312 10.6151
R972 B.n313 B.n141 10.6151
R973 B.n319 B.n141 10.6151
R974 B.n320 B.n319 10.6151
R975 B.n321 B.n320 10.6151
R976 B.n321 B.n139 10.6151
R977 B.n327 B.n139 10.6151
R978 B.n328 B.n327 10.6151
R979 B.n329 B.n328 10.6151
R980 B.n329 B.n137 10.6151
R981 B.n335 B.n137 10.6151
R982 B.n336 B.n335 10.6151
R983 B.n337 B.n336 10.6151
R984 B.n337 B.n135 10.6151
R985 B.n343 B.n135 10.6151
R986 B.n344 B.n343 10.6151
R987 B.n345 B.n344 10.6151
R988 B.n345 B.n133 10.6151
R989 B.n351 B.n133 10.6151
R990 B.n352 B.n351 10.6151
R991 B.n353 B.n352 10.6151
R992 B.n353 B.n131 10.6151
R993 B.n359 B.n131 10.6151
R994 B.n360 B.n359 10.6151
R995 B.n361 B.n360 10.6151
R996 B.n361 B.n129 10.6151
R997 B.n367 B.n129 10.6151
R998 B.n368 B.n367 10.6151
R999 B.n369 B.n368 10.6151
R1000 B.n369 B.n127 10.6151
R1001 B.n375 B.n127 10.6151
R1002 B.n376 B.n375 10.6151
R1003 B.n377 B.n376 10.6151
R1004 B.n377 B.n125 10.6151
R1005 B.n125 B.n124 10.6151
R1006 B.n384 B.n124 10.6151
R1007 B.n385 B.n384 10.6151
R1008 B.n386 B.n116 10.6151
R1009 B.n396 B.n116 10.6151
R1010 B.n397 B.n396 10.6151
R1011 B.n398 B.n397 10.6151
R1012 B.n398 B.n108 10.6151
R1013 B.n408 B.n108 10.6151
R1014 B.n409 B.n408 10.6151
R1015 B.n410 B.n409 10.6151
R1016 B.n410 B.n101 10.6151
R1017 B.n421 B.n101 10.6151
R1018 B.n422 B.n421 10.6151
R1019 B.n424 B.n422 10.6151
R1020 B.n424 B.n423 10.6151
R1021 B.n423 B.n93 10.6151
R1022 B.n435 B.n93 10.6151
R1023 B.n436 B.n435 10.6151
R1024 B.n437 B.n436 10.6151
R1025 B.n438 B.n437 10.6151
R1026 B.n439 B.n438 10.6151
R1027 B.n440 B.n439 10.6151
R1028 B.n441 B.n440 10.6151
R1029 B.n443 B.n441 10.6151
R1030 B.n444 B.n443 10.6151
R1031 B.n445 B.n444 10.6151
R1032 B.n446 B.n445 10.6151
R1033 B.n448 B.n446 10.6151
R1034 B.n449 B.n448 10.6151
R1035 B.n450 B.n449 10.6151
R1036 B.n451 B.n450 10.6151
R1037 B.n453 B.n451 10.6151
R1038 B.n454 B.n453 10.6151
R1039 B.n455 B.n454 10.6151
R1040 B.n456 B.n455 10.6151
R1041 B.n9 B.n1 10.6151
R1042 B.n15 B.n9 10.6151
R1043 B.n690 B.n15 10.6151
R1044 B.n690 B.n689 10.6151
R1045 B.n689 B.n688 10.6151
R1046 B.n688 B.n16 10.6151
R1047 B.n682 B.n16 10.6151
R1048 B.n682 B.n681 10.6151
R1049 B.n681 B.n680 10.6151
R1050 B.n680 B.n23 10.6151
R1051 B.n674 B.n23 10.6151
R1052 B.n674 B.n673 10.6151
R1053 B.n673 B.n672 10.6151
R1054 B.n672 B.n30 10.6151
R1055 B.n666 B.n30 10.6151
R1056 B.n665 B.n664 10.6151
R1057 B.n664 B.n37 10.6151
R1058 B.n658 B.n37 10.6151
R1059 B.n658 B.n657 10.6151
R1060 B.n657 B.n656 10.6151
R1061 B.n656 B.n39 10.6151
R1062 B.n650 B.n39 10.6151
R1063 B.n650 B.n649 10.6151
R1064 B.n649 B.n648 10.6151
R1065 B.n648 B.n41 10.6151
R1066 B.n642 B.n41 10.6151
R1067 B.n642 B.n641 10.6151
R1068 B.n641 B.n640 10.6151
R1069 B.n640 B.n43 10.6151
R1070 B.n634 B.n43 10.6151
R1071 B.n634 B.n633 10.6151
R1072 B.n633 B.n632 10.6151
R1073 B.n632 B.n45 10.6151
R1074 B.n626 B.n45 10.6151
R1075 B.n626 B.n625 10.6151
R1076 B.n625 B.n624 10.6151
R1077 B.n624 B.n47 10.6151
R1078 B.n618 B.n47 10.6151
R1079 B.n618 B.n617 10.6151
R1080 B.n617 B.n616 10.6151
R1081 B.n616 B.n49 10.6151
R1082 B.n610 B.n49 10.6151
R1083 B.n610 B.n609 10.6151
R1084 B.n609 B.n608 10.6151
R1085 B.n608 B.n51 10.6151
R1086 B.n602 B.n51 10.6151
R1087 B.n602 B.n601 10.6151
R1088 B.n601 B.n600 10.6151
R1089 B.n600 B.n53 10.6151
R1090 B.n594 B.n53 10.6151
R1091 B.n594 B.n593 10.6151
R1092 B.n593 B.n592 10.6151
R1093 B.n592 B.n55 10.6151
R1094 B.n586 B.n55 10.6151
R1095 B.n586 B.n585 10.6151
R1096 B.n585 B.n584 10.6151
R1097 B.n584 B.n57 10.6151
R1098 B.n578 B.n57 10.6151
R1099 B.n578 B.n577 10.6151
R1100 B.n577 B.n576 10.6151
R1101 B.n576 B.n59 10.6151
R1102 B.n570 B.n569 10.6151
R1103 B.n569 B.n568 10.6151
R1104 B.n568 B.n64 10.6151
R1105 B.n562 B.n64 10.6151
R1106 B.n562 B.n561 10.6151
R1107 B.n561 B.n560 10.6151
R1108 B.n560 B.n66 10.6151
R1109 B.n554 B.n66 10.6151
R1110 B.n554 B.n553 10.6151
R1111 B.n551 B.n70 10.6151
R1112 B.n545 B.n70 10.6151
R1113 B.n545 B.n544 10.6151
R1114 B.n544 B.n543 10.6151
R1115 B.n543 B.n72 10.6151
R1116 B.n537 B.n72 10.6151
R1117 B.n537 B.n536 10.6151
R1118 B.n536 B.n535 10.6151
R1119 B.n535 B.n74 10.6151
R1120 B.n529 B.n74 10.6151
R1121 B.n529 B.n528 10.6151
R1122 B.n528 B.n527 10.6151
R1123 B.n527 B.n76 10.6151
R1124 B.n521 B.n76 10.6151
R1125 B.n521 B.n520 10.6151
R1126 B.n520 B.n519 10.6151
R1127 B.n519 B.n78 10.6151
R1128 B.n513 B.n78 10.6151
R1129 B.n513 B.n512 10.6151
R1130 B.n512 B.n511 10.6151
R1131 B.n511 B.n80 10.6151
R1132 B.n505 B.n80 10.6151
R1133 B.n505 B.n504 10.6151
R1134 B.n504 B.n503 10.6151
R1135 B.n503 B.n82 10.6151
R1136 B.n497 B.n82 10.6151
R1137 B.n497 B.n496 10.6151
R1138 B.n496 B.n495 10.6151
R1139 B.n495 B.n84 10.6151
R1140 B.n489 B.n84 10.6151
R1141 B.n489 B.n488 10.6151
R1142 B.n488 B.n487 10.6151
R1143 B.n487 B.n86 10.6151
R1144 B.n481 B.n86 10.6151
R1145 B.n481 B.n480 10.6151
R1146 B.n480 B.n479 10.6151
R1147 B.n479 B.n88 10.6151
R1148 B.n473 B.n88 10.6151
R1149 B.n473 B.n472 10.6151
R1150 B.n472 B.n471 10.6151
R1151 B.n471 B.n90 10.6151
R1152 B.n465 B.n90 10.6151
R1153 B.n465 B.n464 10.6151
R1154 B.n464 B.n463 10.6151
R1155 B.n463 B.n92 10.6151
R1156 B.n457 B.n92 10.6151
R1157 B.n272 B.n271 9.36635
R1158 B.n295 B.n149 9.36635
R1159 B.n63 B.n59 9.36635
R1160 B.n552 B.n551 9.36635
R1161 B.n702 B.n0 8.11757
R1162 B.n702 B.n1 8.11757
R1163 B.n400 B.t14 5.74613
R1164 B.t7 B.n676 5.74613
R1165 B.n432 B.t5 2.29875
R1166 B.n694 B.t4 2.29875
R1167 B.n273 B.n272 1.24928
R1168 B.n150 B.n149 1.24928
R1169 B.n570 B.n63 1.24928
R1170 B.n553 B.n552 1.24928
R1171 B.n412 B.t20 1.14963
R1172 B.t21 B.n685 1.14963
R1173 VN.n5 VN.t3 1576.18
R1174 VN.n1 VN.t1 1576.18
R1175 VN.n12 VN.t0 1576.18
R1176 VN.n8 VN.t4 1576.18
R1177 VN.n4 VN.t2 1524.32
R1178 VN.n2 VN.t5 1524.32
R1179 VN.n11 VN.t7 1524.32
R1180 VN.n9 VN.t6 1524.32
R1181 VN.n8 VN.n7 161.489
R1182 VN.n1 VN.n0 161.489
R1183 VN.n6 VN.n5 161.3
R1184 VN.n13 VN.n12 161.3
R1185 VN.n10 VN.n7 161.3
R1186 VN.n3 VN.n0 161.3
R1187 VN VN.n13 41.76
R1188 VN.n3 VN.n2 41.6278
R1189 VN.n4 VN.n3 41.6278
R1190 VN.n11 VN.n10 41.6278
R1191 VN.n10 VN.n9 41.6278
R1192 VN.n2 VN.n1 31.4035
R1193 VN.n5 VN.n4 31.4035
R1194 VN.n12 VN.n11 31.4035
R1195 VN.n9 VN.n8 31.4035
R1196 VN.n13 VN.n7 0.189894
R1197 VN.n6 VN.n0 0.189894
R1198 VN VN.n6 0.0516364
R1199 VDD2.n2 VDD2.n1 60.7089
R1200 VDD2.n2 VDD2.n0 60.7089
R1201 VDD2 VDD2.n5 60.7061
R1202 VDD2.n4 VDD2.n3 60.5186
R1203 VDD2.n4 VDD2.n2 37.8834
R1204 VDD2.n5 VDD2.t6 1.42804
R1205 VDD2.n5 VDD2.t1 1.42804
R1206 VDD2.n3 VDD2.t3 1.42804
R1207 VDD2.n3 VDD2.t4 1.42804
R1208 VDD2.n1 VDD2.t7 1.42804
R1209 VDD2.n1 VDD2.t5 1.42804
R1210 VDD2.n0 VDD2.t0 1.42804
R1211 VDD2.n0 VDD2.t2 1.42804
R1212 VDD2 VDD2.n4 0.304379
R1213 VTAIL.n14 VTAIL.t7 45.2674
R1214 VTAIL.n11 VTAIL.t3 45.2673
R1215 VTAIL.n10 VTAIL.t11 45.2673
R1216 VTAIL.n7 VTAIL.t15 45.2673
R1217 VTAIL.n15 VTAIL.t12 45.2672
R1218 VTAIL.n2 VTAIL.t14 45.2672
R1219 VTAIL.n3 VTAIL.t2 45.2672
R1220 VTAIL.n6 VTAIL.t4 45.2672
R1221 VTAIL.n13 VTAIL.n12 43.8398
R1222 VTAIL.n9 VTAIL.n8 43.8398
R1223 VTAIL.n1 VTAIL.n0 43.8398
R1224 VTAIL.n5 VTAIL.n4 43.8398
R1225 VTAIL.n15 VTAIL.n14 24.8152
R1226 VTAIL.n7 VTAIL.n6 24.8152
R1227 VTAIL.n0 VTAIL.t10 1.42804
R1228 VTAIL.n0 VTAIL.t13 1.42804
R1229 VTAIL.n4 VTAIL.t5 1.42804
R1230 VTAIL.n4 VTAIL.t1 1.42804
R1231 VTAIL.n12 VTAIL.t6 1.42804
R1232 VTAIL.n12 VTAIL.t0 1.42804
R1233 VTAIL.n8 VTAIL.t8 1.42804
R1234 VTAIL.n8 VTAIL.t9 1.42804
R1235 VTAIL.n9 VTAIL.n7 0.491879
R1236 VTAIL.n10 VTAIL.n9 0.491879
R1237 VTAIL.n13 VTAIL.n11 0.491879
R1238 VTAIL.n14 VTAIL.n13 0.491879
R1239 VTAIL.n6 VTAIL.n5 0.491879
R1240 VTAIL.n5 VTAIL.n3 0.491879
R1241 VTAIL.n2 VTAIL.n1 0.491879
R1242 VTAIL.n11 VTAIL.n10 0.470328
R1243 VTAIL.n3 VTAIL.n2 0.470328
R1244 VTAIL VTAIL.n15 0.43369
R1245 VTAIL VTAIL.n1 0.0586897
R1246 VP.n13 VP.t0 1576.18
R1247 VP.n9 VP.t2 1576.18
R1248 VP.n2 VP.t6 1576.18
R1249 VP.n6 VP.t4 1576.18
R1250 VP.n12 VP.t5 1524.32
R1251 VP.n10 VP.t7 1524.32
R1252 VP.n3 VP.t1 1524.32
R1253 VP.n5 VP.t3 1524.32
R1254 VP.n2 VP.n1 161.489
R1255 VP.n14 VP.n13 161.3
R1256 VP.n4 VP.n1 161.3
R1257 VP.n7 VP.n6 161.3
R1258 VP.n11 VP.n0 161.3
R1259 VP.n9 VP.n8 161.3
R1260 VP.n11 VP.n10 41.6278
R1261 VP.n12 VP.n11 41.6278
R1262 VP.n4 VP.n3 41.6278
R1263 VP.n5 VP.n4 41.6278
R1264 VP.n8 VP.n7 41.3793
R1265 VP.n10 VP.n9 31.4035
R1266 VP.n13 VP.n12 31.4035
R1267 VP.n3 VP.n2 31.4035
R1268 VP.n6 VP.n5 31.4035
R1269 VP.n7 VP.n1 0.189894
R1270 VP.n8 VP.n0 0.189894
R1271 VP.n14 VP.n0 0.189894
R1272 VP VP.n14 0.0516364
R1273 VDD1 VDD1.n0 60.8225
R1274 VDD1.n3 VDD1.n2 60.7089
R1275 VDD1.n3 VDD1.n1 60.7089
R1276 VDD1.n5 VDD1.n4 60.5186
R1277 VDD1.n5 VDD1.n3 38.4664
R1278 VDD1.n4 VDD1.t4 1.42804
R1279 VDD1.n4 VDD1.t3 1.42804
R1280 VDD1.n0 VDD1.t1 1.42804
R1281 VDD1.n0 VDD1.t6 1.42804
R1282 VDD1.n2 VDD1.t2 1.42804
R1283 VDD1.n2 VDD1.t7 1.42804
R1284 VDD1.n1 VDD1.t5 1.42804
R1285 VDD1.n1 VDD1.t0 1.42804
R1286 VDD1 VDD1.n5 0.188
C0 VDD1 VDD2 0.602088f
C1 VTAIL VDD2 20.6841f
C2 VDD1 VN 0.147137f
C3 VN VTAIL 2.77126f
C4 VP VDD2 0.268217f
C5 VN VP 5.12081f
C6 VDD1 VTAIL 20.6455f
C7 VDD1 VP 3.43411f
C8 VTAIL VP 2.78537f
C9 VN VDD2 3.31324f
C10 VDD2 B 3.256206f
C11 VDD1 B 3.427243f
C12 VTAIL B 9.382847f
C13 VN B 7.39499f
C14 VP B 4.958063f
C15 VDD1.t1 B 0.392622f
C16 VDD1.t6 B 0.392622f
C17 VDD1.n0 B 3.52716f
C18 VDD1.t5 B 0.392622f
C19 VDD1.t0 B 0.392622f
C20 VDD1.n1 B 3.52637f
C21 VDD1.t2 B 0.392622f
C22 VDD1.t7 B 0.392622f
C23 VDD1.n2 B 3.52637f
C24 VDD1.n3 B 2.98102f
C25 VDD1.t4 B 0.392622f
C26 VDD1.t3 B 0.392622f
C27 VDD1.n4 B 3.52512f
C28 VDD1.n5 B 3.31019f
C29 VP.n0 B 0.058456f
C30 VP.t5 B 0.549392f
C31 VP.t7 B 0.549392f
C32 VP.t2 B 0.556642f
C33 VP.n1 B 0.133043f
C34 VP.t3 B 0.549392f
C35 VP.t1 B 0.549392f
C36 VP.t6 B 0.556642f
C37 VP.n2 B 0.235141f
C38 VP.n3 B 0.216965f
C39 VP.n4 B 0.021915f
C40 VP.n5 B 0.216965f
C41 VP.t4 B 0.556642f
C42 VP.n6 B 0.235054f
C43 VP.n7 B 2.35346f
C44 VP.n8 B 2.40424f
C45 VP.n9 B 0.235054f
C46 VP.n10 B 0.216965f
C47 VP.n11 B 0.021915f
C48 VP.n12 B 0.216965f
C49 VP.t0 B 0.556642f
C50 VP.n13 B 0.235054f
C51 VP.n14 B 0.045301f
C52 VTAIL.t10 B 0.27957f
C53 VTAIL.t13 B 0.27957f
C54 VTAIL.n0 B 2.43016f
C55 VTAIL.n1 B 0.305401f
C56 VTAIL.t14 B 3.10074f
C57 VTAIL.n2 B 0.431114f
C58 VTAIL.t2 B 3.10074f
C59 VTAIL.n3 B 0.431114f
C60 VTAIL.t5 B 0.27957f
C61 VTAIL.t1 B 0.27957f
C62 VTAIL.n4 B 2.43016f
C63 VTAIL.n5 B 0.341004f
C64 VTAIL.t4 B 3.10074f
C65 VTAIL.n6 B 1.7621f
C66 VTAIL.t15 B 3.10076f
C67 VTAIL.n7 B 1.76208f
C68 VTAIL.t8 B 0.27957f
C69 VTAIL.t9 B 0.27957f
C70 VTAIL.n8 B 2.43016f
C71 VTAIL.n9 B 0.341006f
C72 VTAIL.t11 B 3.10076f
C73 VTAIL.n10 B 0.431096f
C74 VTAIL.t3 B 3.10076f
C75 VTAIL.n11 B 0.431096f
C76 VTAIL.t6 B 0.27957f
C77 VTAIL.t0 B 0.27957f
C78 VTAIL.n12 B 2.43016f
C79 VTAIL.n13 B 0.341006f
C80 VTAIL.t7 B 3.10075f
C81 VTAIL.n14 B 1.76209f
C82 VTAIL.t12 B 3.10074f
C83 VTAIL.n15 B 1.75732f
C84 VDD2.t0 B 0.394799f
C85 VDD2.t2 B 0.394799f
C86 VDD2.n0 B 3.54592f
C87 VDD2.t7 B 0.394799f
C88 VDD2.t5 B 0.394799f
C89 VDD2.n1 B 3.54592f
C90 VDD2.n2 B 2.92029f
C91 VDD2.t3 B 0.394799f
C92 VDD2.t4 B 0.394799f
C93 VDD2.n3 B 3.54466f
C94 VDD2.n4 B 3.28627f
C95 VDD2.t6 B 0.394799f
C96 VDD2.t1 B 0.394799f
C97 VDD2.n5 B 3.54588f
C98 VN.n0 B 0.130914f
C99 VN.t2 B 0.540599f
C100 VN.t5 B 0.540599f
C101 VN.t1 B 0.547733f
C102 VN.n1 B 0.231378f
C103 VN.n2 B 0.213493f
C104 VN.n3 B 0.021564f
C105 VN.n4 B 0.213493f
C106 VN.t3 B 0.547733f
C107 VN.n5 B 0.231292f
C108 VN.n6 B 0.044576f
C109 VN.n7 B 0.130914f
C110 VN.t0 B 0.547733f
C111 VN.t7 B 0.540599f
C112 VN.t6 B 0.540599f
C113 VN.t4 B 0.547733f
C114 VN.n8 B 0.231378f
C115 VN.n9 B 0.213493f
C116 VN.n10 B 0.021564f
C117 VN.n11 B 0.213493f
C118 VN.n12 B 0.231292f
C119 VN.n13 B 2.35358f
.ends

