* NGSPICE file created from diff_pair_sample_1511.ext - technology: sky130A

.subckt diff_pair_sample_1511 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X1 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X2 VTAIL.t18 VN.t1 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X3 VDD1.t8 VP.t1 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X4 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.9321 ps=5.56 w=2.39 l=2.63
X5 VTAIL.t6 VP.t3 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X6 VDD2.t1 VN.t2 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X7 VDD2.t2 VN.t3 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X8 VDD2.t3 VN.t4 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0.39435 ps=2.72 w=2.39 l=2.63
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0 ps=0 w=2.39 l=2.63
X10 VDD1.t5 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0.39435 ps=2.72 w=2.39 l=2.63
X11 VTAIL.t14 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X12 VTAIL.t2 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X13 VDD1.t3 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.9321 ps=5.56 w=2.39 l=2.63
X14 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0 ps=0 w=2.39 l=2.63
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0 ps=0 w=2.39 l=2.63
X16 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0.39435 ps=2.72 w=2.39 l=2.63
X17 VDD2.t7 VN.t6 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.9321 ps=5.56 w=2.39 l=2.63
X18 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X19 VDD2.t8 VN.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.9321 ps=5.56 w=2.39 l=2.63
X20 VDD2.t9 VN.t8 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0.39435 ps=2.72 w=2.39 l=2.63
X21 VTAIL.t10 VN.t9 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9321 pd=5.56 as=0 ps=0 w=2.39 l=2.63
X23 VTAIL.t3 VP.t9 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.39435 pd=2.72 as=0.39435 ps=2.72 w=2.39 l=2.63
R0 VN.n81 VN.n42 161.3
R1 VN.n80 VN.n79 161.3
R2 VN.n78 VN.n43 161.3
R3 VN.n77 VN.n76 161.3
R4 VN.n75 VN.n44 161.3
R5 VN.n74 VN.n73 161.3
R6 VN.n72 VN.n71 161.3
R7 VN.n70 VN.n46 161.3
R8 VN.n69 VN.n68 161.3
R9 VN.n67 VN.n47 161.3
R10 VN.n66 VN.n65 161.3
R11 VN.n64 VN.n48 161.3
R12 VN.n62 VN.n61 161.3
R13 VN.n60 VN.n49 161.3
R14 VN.n59 VN.n58 161.3
R15 VN.n57 VN.n50 161.3
R16 VN.n56 VN.n55 161.3
R17 VN.n54 VN.n51 161.3
R18 VN.n39 VN.n0 161.3
R19 VN.n38 VN.n37 161.3
R20 VN.n36 VN.n1 161.3
R21 VN.n35 VN.n34 161.3
R22 VN.n33 VN.n2 161.3
R23 VN.n32 VN.n31 161.3
R24 VN.n30 VN.n29 161.3
R25 VN.n28 VN.n4 161.3
R26 VN.n27 VN.n26 161.3
R27 VN.n25 VN.n5 161.3
R28 VN.n24 VN.n23 161.3
R29 VN.n22 VN.n6 161.3
R30 VN.n20 VN.n19 161.3
R31 VN.n18 VN.n7 161.3
R32 VN.n17 VN.n16 161.3
R33 VN.n15 VN.n8 161.3
R34 VN.n14 VN.n13 161.3
R35 VN.n12 VN.n9 161.3
R36 VN.n41 VN.n40 102.438
R37 VN.n83 VN.n82 102.438
R38 VN.n11 VN.n10 62.0711
R39 VN.n53 VN.n52 62.0711
R40 VN.n16 VN.n15 56.5193
R41 VN.n27 VN.n5 56.5193
R42 VN.n34 VN.n1 56.5193
R43 VN.n58 VN.n57 56.5193
R44 VN.n69 VN.n47 56.5193
R45 VN.n76 VN.n43 56.5193
R46 VN.n11 VN.t4 55.0181
R47 VN.n53 VN.t6 55.0181
R48 VN VN.n83 46.2785
R49 VN.n14 VN.n9 24.4675
R50 VN.n15 VN.n14 24.4675
R51 VN.n16 VN.n7 24.4675
R52 VN.n20 VN.n7 24.4675
R53 VN.n23 VN.n22 24.4675
R54 VN.n23 VN.n5 24.4675
R55 VN.n28 VN.n27 24.4675
R56 VN.n29 VN.n28 24.4675
R57 VN.n33 VN.n32 24.4675
R58 VN.n34 VN.n33 24.4675
R59 VN.n38 VN.n1 24.4675
R60 VN.n39 VN.n38 24.4675
R61 VN.n57 VN.n56 24.4675
R62 VN.n56 VN.n51 24.4675
R63 VN.n65 VN.n47 24.4675
R64 VN.n65 VN.n64 24.4675
R65 VN.n62 VN.n49 24.4675
R66 VN.n58 VN.n49 24.4675
R67 VN.n76 VN.n75 24.4675
R68 VN.n75 VN.n74 24.4675
R69 VN.n71 VN.n70 24.4675
R70 VN.n70 VN.n69 24.4675
R71 VN.n81 VN.n80 24.4675
R72 VN.n80 VN.n43 24.4675
R73 VN.n10 VN.t9 21.9013
R74 VN.n21 VN.t2 21.9013
R75 VN.n3 VN.t0 21.9013
R76 VN.n40 VN.t7 21.9013
R77 VN.n52 VN.t5 21.9013
R78 VN.n63 VN.t3 21.9013
R79 VN.n45 VN.t1 21.9013
R80 VN.n82 VN.t8 21.9013
R81 VN.n32 VN.n3 14.1914
R82 VN.n74 VN.n45 14.1914
R83 VN.n21 VN.n20 12.234
R84 VN.n22 VN.n21 12.234
R85 VN.n64 VN.n63 12.234
R86 VN.n63 VN.n62 12.234
R87 VN.n10 VN.n9 10.2766
R88 VN.n29 VN.n3 10.2766
R89 VN.n52 VN.n51 10.2766
R90 VN.n71 VN.n45 10.2766
R91 VN.n40 VN.n39 8.31928
R92 VN.n82 VN.n81 8.31928
R93 VN.n54 VN.n53 6.95571
R94 VN.n12 VN.n11 6.95571
R95 VN.n83 VN.n42 0.278367
R96 VN.n41 VN.n0 0.278367
R97 VN.n79 VN.n42 0.189894
R98 VN.n79 VN.n78 0.189894
R99 VN.n78 VN.n77 0.189894
R100 VN.n77 VN.n44 0.189894
R101 VN.n73 VN.n44 0.189894
R102 VN.n73 VN.n72 0.189894
R103 VN.n72 VN.n46 0.189894
R104 VN.n68 VN.n46 0.189894
R105 VN.n68 VN.n67 0.189894
R106 VN.n67 VN.n66 0.189894
R107 VN.n66 VN.n48 0.189894
R108 VN.n61 VN.n48 0.189894
R109 VN.n61 VN.n60 0.189894
R110 VN.n60 VN.n59 0.189894
R111 VN.n59 VN.n50 0.189894
R112 VN.n55 VN.n50 0.189894
R113 VN.n55 VN.n54 0.189894
R114 VN.n13 VN.n12 0.189894
R115 VN.n13 VN.n8 0.189894
R116 VN.n17 VN.n8 0.189894
R117 VN.n18 VN.n17 0.189894
R118 VN.n19 VN.n18 0.189894
R119 VN.n19 VN.n6 0.189894
R120 VN.n24 VN.n6 0.189894
R121 VN.n25 VN.n24 0.189894
R122 VN.n26 VN.n25 0.189894
R123 VN.n26 VN.n4 0.189894
R124 VN.n30 VN.n4 0.189894
R125 VN.n31 VN.n30 0.189894
R126 VN.n31 VN.n2 0.189894
R127 VN.n35 VN.n2 0.189894
R128 VN.n36 VN.n35 0.189894
R129 VN.n37 VN.n36 0.189894
R130 VN.n37 VN.n0 0.189894
R131 VN VN.n41 0.153454
R132 VDD2.n21 VDD2.n15 289.615
R133 VDD2.n6 VDD2.n0 289.615
R134 VDD2.n22 VDD2.n21 185
R135 VDD2.n20 VDD2.n19 185
R136 VDD2.n5 VDD2.n4 185
R137 VDD2.n7 VDD2.n6 185
R138 VDD2.n18 VDD2.t9 151.613
R139 VDD2.n3 VDD2.t3 151.613
R140 VDD2.n21 VDD2.n20 104.615
R141 VDD2.n6 VDD2.n5 104.615
R142 VDD2.n14 VDD2.n13 86.6237
R143 VDD2 VDD2.n29 86.6208
R144 VDD2.n28 VDD2.n27 84.7653
R145 VDD2.n12 VDD2.n11 84.7652
R146 VDD2.n20 VDD2.t9 52.3082
R147 VDD2.n5 VDD2.t3 52.3082
R148 VDD2.n12 VDD2.n10 51.2219
R149 VDD2.n26 VDD2.n25 48.6702
R150 VDD2.n26 VDD2.n14 37.8963
R151 VDD2.n19 VDD2.n18 15.3979
R152 VDD2.n4 VDD2.n3 15.3979
R153 VDD2.n22 VDD2.n17 12.8005
R154 VDD2.n7 VDD2.n2 12.8005
R155 VDD2.n23 VDD2.n15 12.0247
R156 VDD2.n8 VDD2.n0 12.0247
R157 VDD2.n25 VDD2.n24 9.45567
R158 VDD2.n10 VDD2.n9 9.45567
R159 VDD2.n24 VDD2.n23 9.3005
R160 VDD2.n17 VDD2.n16 9.3005
R161 VDD2.n9 VDD2.n8 9.3005
R162 VDD2.n2 VDD2.n1 9.3005
R163 VDD2.n29 VDD2.t4 8.28502
R164 VDD2.n29 VDD2.t7 8.28502
R165 VDD2.n27 VDD2.t0 8.28502
R166 VDD2.n27 VDD2.t2 8.28502
R167 VDD2.n13 VDD2.t5 8.28502
R168 VDD2.n13 VDD2.t8 8.28502
R169 VDD2.n11 VDD2.t6 8.28502
R170 VDD2.n11 VDD2.t1 8.28502
R171 VDD2.n18 VDD2.n16 4.69785
R172 VDD2.n3 VDD2.n1 4.69785
R173 VDD2.n28 VDD2.n26 2.55222
R174 VDD2.n25 VDD2.n15 1.93989
R175 VDD2.n10 VDD2.n0 1.93989
R176 VDD2.n23 VDD2.n22 1.16414
R177 VDD2.n8 VDD2.n7 1.16414
R178 VDD2 VDD2.n28 0.696621
R179 VDD2.n14 VDD2.n12 0.583085
R180 VDD2.n19 VDD2.n17 0.388379
R181 VDD2.n4 VDD2.n2 0.388379
R182 VDD2.n24 VDD2.n16 0.155672
R183 VDD2.n9 VDD2.n1 0.155672
R184 VTAIL.n56 VTAIL.n50 289.615
R185 VTAIL.n8 VTAIL.n2 289.615
R186 VTAIL.n44 VTAIL.n38 289.615
R187 VTAIL.n28 VTAIL.n22 289.615
R188 VTAIL.n55 VTAIL.n54 185
R189 VTAIL.n57 VTAIL.n56 185
R190 VTAIL.n7 VTAIL.n6 185
R191 VTAIL.n9 VTAIL.n8 185
R192 VTAIL.n45 VTAIL.n44 185
R193 VTAIL.n43 VTAIL.n42 185
R194 VTAIL.n29 VTAIL.n28 185
R195 VTAIL.n27 VTAIL.n26 185
R196 VTAIL.n53 VTAIL.t12 151.613
R197 VTAIL.n5 VTAIL.t4 151.613
R198 VTAIL.n41 VTAIL.t8 151.613
R199 VTAIL.n25 VTAIL.t13 151.613
R200 VTAIL.n56 VTAIL.n55 104.615
R201 VTAIL.n8 VTAIL.n7 104.615
R202 VTAIL.n44 VTAIL.n43 104.615
R203 VTAIL.n28 VTAIL.n27 104.615
R204 VTAIL.n37 VTAIL.n36 68.0866
R205 VTAIL.n35 VTAIL.n34 68.0866
R206 VTAIL.n21 VTAIL.n20 68.0866
R207 VTAIL.n19 VTAIL.n18 68.0866
R208 VTAIL.n63 VTAIL.n62 68.0865
R209 VTAIL.n1 VTAIL.n0 68.0865
R210 VTAIL.n15 VTAIL.n14 68.0865
R211 VTAIL.n17 VTAIL.n16 68.0865
R212 VTAIL.n55 VTAIL.t12 52.3082
R213 VTAIL.n7 VTAIL.t4 52.3082
R214 VTAIL.n43 VTAIL.t8 52.3082
R215 VTAIL.n27 VTAIL.t13 52.3082
R216 VTAIL.n61 VTAIL.n60 31.9914
R217 VTAIL.n13 VTAIL.n12 31.9914
R218 VTAIL.n49 VTAIL.n48 31.9914
R219 VTAIL.n33 VTAIL.n32 31.9914
R220 VTAIL.n19 VTAIL.n17 19.5307
R221 VTAIL.n61 VTAIL.n49 16.9789
R222 VTAIL.n54 VTAIL.n53 15.3979
R223 VTAIL.n6 VTAIL.n5 15.3979
R224 VTAIL.n42 VTAIL.n41 15.3979
R225 VTAIL.n26 VTAIL.n25 15.3979
R226 VTAIL.n57 VTAIL.n52 12.8005
R227 VTAIL.n9 VTAIL.n4 12.8005
R228 VTAIL.n45 VTAIL.n40 12.8005
R229 VTAIL.n29 VTAIL.n24 12.8005
R230 VTAIL.n58 VTAIL.n50 12.0247
R231 VTAIL.n10 VTAIL.n2 12.0247
R232 VTAIL.n46 VTAIL.n38 12.0247
R233 VTAIL.n30 VTAIL.n22 12.0247
R234 VTAIL.n60 VTAIL.n59 9.45567
R235 VTAIL.n12 VTAIL.n11 9.45567
R236 VTAIL.n48 VTAIL.n47 9.45567
R237 VTAIL.n32 VTAIL.n31 9.45567
R238 VTAIL.n59 VTAIL.n58 9.3005
R239 VTAIL.n52 VTAIL.n51 9.3005
R240 VTAIL.n11 VTAIL.n10 9.3005
R241 VTAIL.n4 VTAIL.n3 9.3005
R242 VTAIL.n47 VTAIL.n46 9.3005
R243 VTAIL.n40 VTAIL.n39 9.3005
R244 VTAIL.n31 VTAIL.n30 9.3005
R245 VTAIL.n24 VTAIL.n23 9.3005
R246 VTAIL.n62 VTAIL.t17 8.28502
R247 VTAIL.n62 VTAIL.t19 8.28502
R248 VTAIL.n0 VTAIL.t15 8.28502
R249 VTAIL.n0 VTAIL.t10 8.28502
R250 VTAIL.n14 VTAIL.t9 8.28502
R251 VTAIL.n14 VTAIL.t3 8.28502
R252 VTAIL.n16 VTAIL.t5 8.28502
R253 VTAIL.n16 VTAIL.t2 8.28502
R254 VTAIL.n36 VTAIL.t7 8.28502
R255 VTAIL.n36 VTAIL.t1 8.28502
R256 VTAIL.n34 VTAIL.t0 8.28502
R257 VTAIL.n34 VTAIL.t6 8.28502
R258 VTAIL.n20 VTAIL.t16 8.28502
R259 VTAIL.n20 VTAIL.t14 8.28502
R260 VTAIL.n18 VTAIL.t11 8.28502
R261 VTAIL.n18 VTAIL.t18 8.28502
R262 VTAIL.n53 VTAIL.n51 4.69785
R263 VTAIL.n5 VTAIL.n3 4.69785
R264 VTAIL.n41 VTAIL.n39 4.69785
R265 VTAIL.n25 VTAIL.n23 4.69785
R266 VTAIL.n21 VTAIL.n19 2.55222
R267 VTAIL.n33 VTAIL.n21 2.55222
R268 VTAIL.n37 VTAIL.n35 2.55222
R269 VTAIL.n49 VTAIL.n37 2.55222
R270 VTAIL.n17 VTAIL.n15 2.55222
R271 VTAIL.n15 VTAIL.n13 2.55222
R272 VTAIL.n63 VTAIL.n61 2.55222
R273 VTAIL VTAIL.n1 1.97248
R274 VTAIL.n60 VTAIL.n50 1.93989
R275 VTAIL.n12 VTAIL.n2 1.93989
R276 VTAIL.n48 VTAIL.n38 1.93989
R277 VTAIL.n32 VTAIL.n22 1.93989
R278 VTAIL.n35 VTAIL.n33 1.74619
R279 VTAIL.n13 VTAIL.n1 1.74619
R280 VTAIL.n58 VTAIL.n57 1.16414
R281 VTAIL.n10 VTAIL.n9 1.16414
R282 VTAIL.n46 VTAIL.n45 1.16414
R283 VTAIL.n30 VTAIL.n29 1.16414
R284 VTAIL VTAIL.n63 0.580241
R285 VTAIL.n54 VTAIL.n52 0.388379
R286 VTAIL.n6 VTAIL.n4 0.388379
R287 VTAIL.n42 VTAIL.n40 0.388379
R288 VTAIL.n26 VTAIL.n24 0.388379
R289 VTAIL.n59 VTAIL.n51 0.155672
R290 VTAIL.n11 VTAIL.n3 0.155672
R291 VTAIL.n47 VTAIL.n39 0.155672
R292 VTAIL.n31 VTAIL.n23 0.155672
R293 B.n675 B.n674 585
R294 B.n202 B.n129 585
R295 B.n201 B.n200 585
R296 B.n199 B.n198 585
R297 B.n197 B.n196 585
R298 B.n195 B.n194 585
R299 B.n193 B.n192 585
R300 B.n191 B.n190 585
R301 B.n189 B.n188 585
R302 B.n187 B.n186 585
R303 B.n185 B.n184 585
R304 B.n183 B.n182 585
R305 B.n181 B.n180 585
R306 B.n178 B.n177 585
R307 B.n176 B.n175 585
R308 B.n174 B.n173 585
R309 B.n172 B.n171 585
R310 B.n170 B.n169 585
R311 B.n168 B.n167 585
R312 B.n166 B.n165 585
R313 B.n164 B.n163 585
R314 B.n162 B.n161 585
R315 B.n160 B.n159 585
R316 B.n157 B.n156 585
R317 B.n155 B.n154 585
R318 B.n153 B.n152 585
R319 B.n151 B.n150 585
R320 B.n149 B.n148 585
R321 B.n147 B.n146 585
R322 B.n145 B.n144 585
R323 B.n143 B.n142 585
R324 B.n141 B.n140 585
R325 B.n139 B.n138 585
R326 B.n137 B.n136 585
R327 B.n135 B.n134 585
R328 B.n110 B.n109 585
R329 B.n673 B.n111 585
R330 B.n678 B.n111 585
R331 B.n672 B.n671 585
R332 B.n671 B.n107 585
R333 B.n670 B.n106 585
R334 B.n684 B.n106 585
R335 B.n669 B.n105 585
R336 B.n685 B.n105 585
R337 B.n668 B.n104 585
R338 B.n686 B.n104 585
R339 B.n667 B.n666 585
R340 B.n666 B.n100 585
R341 B.n665 B.n99 585
R342 B.n692 B.n99 585
R343 B.n664 B.n98 585
R344 B.n693 B.n98 585
R345 B.n663 B.n97 585
R346 B.n694 B.n97 585
R347 B.n662 B.n661 585
R348 B.n661 B.n93 585
R349 B.n660 B.n92 585
R350 B.n700 B.n92 585
R351 B.n659 B.n91 585
R352 B.n701 B.n91 585
R353 B.n658 B.n90 585
R354 B.n702 B.n90 585
R355 B.n657 B.n656 585
R356 B.n656 B.n86 585
R357 B.n655 B.n85 585
R358 B.n708 B.n85 585
R359 B.n654 B.n84 585
R360 B.n709 B.n84 585
R361 B.n653 B.n83 585
R362 B.n710 B.n83 585
R363 B.n652 B.n651 585
R364 B.n651 B.n79 585
R365 B.n650 B.n78 585
R366 B.n716 B.n78 585
R367 B.n649 B.n77 585
R368 B.n717 B.n77 585
R369 B.n648 B.n76 585
R370 B.n718 B.n76 585
R371 B.n647 B.n646 585
R372 B.n646 B.n72 585
R373 B.n645 B.n71 585
R374 B.n724 B.n71 585
R375 B.n644 B.n70 585
R376 B.n725 B.n70 585
R377 B.n643 B.n69 585
R378 B.n726 B.n69 585
R379 B.n642 B.n641 585
R380 B.n641 B.n65 585
R381 B.n640 B.n64 585
R382 B.n732 B.n64 585
R383 B.n639 B.n63 585
R384 B.n733 B.n63 585
R385 B.n638 B.n62 585
R386 B.n734 B.n62 585
R387 B.n637 B.n636 585
R388 B.n636 B.n58 585
R389 B.n635 B.n57 585
R390 B.n740 B.n57 585
R391 B.n634 B.n56 585
R392 B.n741 B.n56 585
R393 B.n633 B.n55 585
R394 B.n742 B.n55 585
R395 B.n632 B.n631 585
R396 B.n631 B.n51 585
R397 B.n630 B.n50 585
R398 B.n748 B.n50 585
R399 B.n629 B.n49 585
R400 B.n749 B.n49 585
R401 B.n628 B.n48 585
R402 B.n750 B.n48 585
R403 B.n627 B.n626 585
R404 B.n626 B.n47 585
R405 B.n625 B.n43 585
R406 B.n756 B.n43 585
R407 B.n624 B.n42 585
R408 B.n757 B.n42 585
R409 B.n623 B.n41 585
R410 B.n758 B.n41 585
R411 B.n622 B.n621 585
R412 B.n621 B.n37 585
R413 B.n620 B.n36 585
R414 B.n764 B.n36 585
R415 B.n619 B.n35 585
R416 B.n765 B.n35 585
R417 B.n618 B.n34 585
R418 B.n766 B.n34 585
R419 B.n617 B.n616 585
R420 B.n616 B.n33 585
R421 B.n615 B.n29 585
R422 B.n772 B.n29 585
R423 B.n614 B.n28 585
R424 B.n773 B.n28 585
R425 B.n613 B.n27 585
R426 B.n774 B.n27 585
R427 B.n612 B.n611 585
R428 B.n611 B.n23 585
R429 B.n610 B.n22 585
R430 B.n780 B.n22 585
R431 B.n609 B.n21 585
R432 B.n781 B.n21 585
R433 B.n608 B.n20 585
R434 B.n782 B.n20 585
R435 B.n607 B.n606 585
R436 B.n606 B.n16 585
R437 B.n605 B.n15 585
R438 B.n788 B.n15 585
R439 B.n604 B.n14 585
R440 B.n789 B.n14 585
R441 B.n603 B.n13 585
R442 B.n790 B.n13 585
R443 B.n602 B.n601 585
R444 B.n601 B.n12 585
R445 B.n600 B.n599 585
R446 B.n600 B.n8 585
R447 B.n598 B.n7 585
R448 B.n797 B.n7 585
R449 B.n597 B.n6 585
R450 B.n798 B.n6 585
R451 B.n596 B.n5 585
R452 B.n799 B.n5 585
R453 B.n595 B.n594 585
R454 B.n594 B.n4 585
R455 B.n593 B.n203 585
R456 B.n593 B.n592 585
R457 B.n583 B.n204 585
R458 B.n205 B.n204 585
R459 B.n585 B.n584 585
R460 B.n586 B.n585 585
R461 B.n582 B.n210 585
R462 B.n210 B.n209 585
R463 B.n581 B.n580 585
R464 B.n580 B.n579 585
R465 B.n212 B.n211 585
R466 B.n213 B.n212 585
R467 B.n572 B.n571 585
R468 B.n573 B.n572 585
R469 B.n570 B.n218 585
R470 B.n218 B.n217 585
R471 B.n569 B.n568 585
R472 B.n568 B.n567 585
R473 B.n220 B.n219 585
R474 B.n221 B.n220 585
R475 B.n560 B.n559 585
R476 B.n561 B.n560 585
R477 B.n558 B.n226 585
R478 B.n226 B.n225 585
R479 B.n557 B.n556 585
R480 B.n556 B.n555 585
R481 B.n228 B.n227 585
R482 B.n548 B.n228 585
R483 B.n547 B.n546 585
R484 B.n549 B.n547 585
R485 B.n545 B.n233 585
R486 B.n233 B.n232 585
R487 B.n544 B.n543 585
R488 B.n543 B.n542 585
R489 B.n235 B.n234 585
R490 B.n236 B.n235 585
R491 B.n535 B.n534 585
R492 B.n536 B.n535 585
R493 B.n533 B.n241 585
R494 B.n241 B.n240 585
R495 B.n532 B.n531 585
R496 B.n531 B.n530 585
R497 B.n243 B.n242 585
R498 B.n523 B.n243 585
R499 B.n522 B.n521 585
R500 B.n524 B.n522 585
R501 B.n520 B.n248 585
R502 B.n248 B.n247 585
R503 B.n519 B.n518 585
R504 B.n518 B.n517 585
R505 B.n250 B.n249 585
R506 B.n251 B.n250 585
R507 B.n510 B.n509 585
R508 B.n511 B.n510 585
R509 B.n508 B.n256 585
R510 B.n256 B.n255 585
R511 B.n507 B.n506 585
R512 B.n506 B.n505 585
R513 B.n258 B.n257 585
R514 B.n259 B.n258 585
R515 B.n498 B.n497 585
R516 B.n499 B.n498 585
R517 B.n496 B.n264 585
R518 B.n264 B.n263 585
R519 B.n495 B.n494 585
R520 B.n494 B.n493 585
R521 B.n266 B.n265 585
R522 B.n267 B.n266 585
R523 B.n486 B.n485 585
R524 B.n487 B.n486 585
R525 B.n484 B.n272 585
R526 B.n272 B.n271 585
R527 B.n483 B.n482 585
R528 B.n482 B.n481 585
R529 B.n274 B.n273 585
R530 B.n275 B.n274 585
R531 B.n474 B.n473 585
R532 B.n475 B.n474 585
R533 B.n472 B.n279 585
R534 B.n283 B.n279 585
R535 B.n471 B.n470 585
R536 B.n470 B.n469 585
R537 B.n281 B.n280 585
R538 B.n282 B.n281 585
R539 B.n462 B.n461 585
R540 B.n463 B.n462 585
R541 B.n460 B.n288 585
R542 B.n288 B.n287 585
R543 B.n459 B.n458 585
R544 B.n458 B.n457 585
R545 B.n290 B.n289 585
R546 B.n291 B.n290 585
R547 B.n450 B.n449 585
R548 B.n451 B.n450 585
R549 B.n448 B.n296 585
R550 B.n296 B.n295 585
R551 B.n447 B.n446 585
R552 B.n446 B.n445 585
R553 B.n298 B.n297 585
R554 B.n299 B.n298 585
R555 B.n438 B.n437 585
R556 B.n439 B.n438 585
R557 B.n436 B.n303 585
R558 B.n307 B.n303 585
R559 B.n435 B.n434 585
R560 B.n434 B.n433 585
R561 B.n305 B.n304 585
R562 B.n306 B.n305 585
R563 B.n426 B.n425 585
R564 B.n427 B.n426 585
R565 B.n424 B.n312 585
R566 B.n312 B.n311 585
R567 B.n423 B.n422 585
R568 B.n422 B.n421 585
R569 B.n314 B.n313 585
R570 B.n315 B.n314 585
R571 B.n414 B.n413 585
R572 B.n415 B.n414 585
R573 B.n318 B.n317 585
R574 B.n345 B.n344 585
R575 B.n346 B.n342 585
R576 B.n342 B.n319 585
R577 B.n348 B.n347 585
R578 B.n350 B.n341 585
R579 B.n353 B.n352 585
R580 B.n354 B.n340 585
R581 B.n356 B.n355 585
R582 B.n358 B.n339 585
R583 B.n361 B.n360 585
R584 B.n362 B.n338 585
R585 B.n364 B.n363 585
R586 B.n366 B.n337 585
R587 B.n369 B.n368 585
R588 B.n370 B.n333 585
R589 B.n372 B.n371 585
R590 B.n374 B.n332 585
R591 B.n377 B.n376 585
R592 B.n378 B.n331 585
R593 B.n380 B.n379 585
R594 B.n382 B.n330 585
R595 B.n385 B.n384 585
R596 B.n386 B.n327 585
R597 B.n389 B.n388 585
R598 B.n391 B.n326 585
R599 B.n394 B.n393 585
R600 B.n395 B.n325 585
R601 B.n397 B.n396 585
R602 B.n399 B.n324 585
R603 B.n402 B.n401 585
R604 B.n403 B.n323 585
R605 B.n405 B.n404 585
R606 B.n407 B.n322 585
R607 B.n408 B.n321 585
R608 B.n411 B.n410 585
R609 B.n412 B.n320 585
R610 B.n320 B.n319 585
R611 B.n417 B.n416 585
R612 B.n416 B.n415 585
R613 B.n418 B.n316 585
R614 B.n316 B.n315 585
R615 B.n420 B.n419 585
R616 B.n421 B.n420 585
R617 B.n310 B.n309 585
R618 B.n311 B.n310 585
R619 B.n429 B.n428 585
R620 B.n428 B.n427 585
R621 B.n430 B.n308 585
R622 B.n308 B.n306 585
R623 B.n432 B.n431 585
R624 B.n433 B.n432 585
R625 B.n302 B.n301 585
R626 B.n307 B.n302 585
R627 B.n441 B.n440 585
R628 B.n440 B.n439 585
R629 B.n442 B.n300 585
R630 B.n300 B.n299 585
R631 B.n444 B.n443 585
R632 B.n445 B.n444 585
R633 B.n294 B.n293 585
R634 B.n295 B.n294 585
R635 B.n453 B.n452 585
R636 B.n452 B.n451 585
R637 B.n454 B.n292 585
R638 B.n292 B.n291 585
R639 B.n456 B.n455 585
R640 B.n457 B.n456 585
R641 B.n286 B.n285 585
R642 B.n287 B.n286 585
R643 B.n465 B.n464 585
R644 B.n464 B.n463 585
R645 B.n466 B.n284 585
R646 B.n284 B.n282 585
R647 B.n468 B.n467 585
R648 B.n469 B.n468 585
R649 B.n278 B.n277 585
R650 B.n283 B.n278 585
R651 B.n477 B.n476 585
R652 B.n476 B.n475 585
R653 B.n478 B.n276 585
R654 B.n276 B.n275 585
R655 B.n480 B.n479 585
R656 B.n481 B.n480 585
R657 B.n270 B.n269 585
R658 B.n271 B.n270 585
R659 B.n489 B.n488 585
R660 B.n488 B.n487 585
R661 B.n490 B.n268 585
R662 B.n268 B.n267 585
R663 B.n492 B.n491 585
R664 B.n493 B.n492 585
R665 B.n262 B.n261 585
R666 B.n263 B.n262 585
R667 B.n501 B.n500 585
R668 B.n500 B.n499 585
R669 B.n502 B.n260 585
R670 B.n260 B.n259 585
R671 B.n504 B.n503 585
R672 B.n505 B.n504 585
R673 B.n254 B.n253 585
R674 B.n255 B.n254 585
R675 B.n513 B.n512 585
R676 B.n512 B.n511 585
R677 B.n514 B.n252 585
R678 B.n252 B.n251 585
R679 B.n516 B.n515 585
R680 B.n517 B.n516 585
R681 B.n246 B.n245 585
R682 B.n247 B.n246 585
R683 B.n526 B.n525 585
R684 B.n525 B.n524 585
R685 B.n527 B.n244 585
R686 B.n523 B.n244 585
R687 B.n529 B.n528 585
R688 B.n530 B.n529 585
R689 B.n239 B.n238 585
R690 B.n240 B.n239 585
R691 B.n538 B.n537 585
R692 B.n537 B.n536 585
R693 B.n539 B.n237 585
R694 B.n237 B.n236 585
R695 B.n541 B.n540 585
R696 B.n542 B.n541 585
R697 B.n231 B.n230 585
R698 B.n232 B.n231 585
R699 B.n551 B.n550 585
R700 B.n550 B.n549 585
R701 B.n552 B.n229 585
R702 B.n548 B.n229 585
R703 B.n554 B.n553 585
R704 B.n555 B.n554 585
R705 B.n224 B.n223 585
R706 B.n225 B.n224 585
R707 B.n563 B.n562 585
R708 B.n562 B.n561 585
R709 B.n564 B.n222 585
R710 B.n222 B.n221 585
R711 B.n566 B.n565 585
R712 B.n567 B.n566 585
R713 B.n216 B.n215 585
R714 B.n217 B.n216 585
R715 B.n575 B.n574 585
R716 B.n574 B.n573 585
R717 B.n576 B.n214 585
R718 B.n214 B.n213 585
R719 B.n578 B.n577 585
R720 B.n579 B.n578 585
R721 B.n208 B.n207 585
R722 B.n209 B.n208 585
R723 B.n588 B.n587 585
R724 B.n587 B.n586 585
R725 B.n589 B.n206 585
R726 B.n206 B.n205 585
R727 B.n591 B.n590 585
R728 B.n592 B.n591 585
R729 B.n3 B.n0 585
R730 B.n4 B.n3 585
R731 B.n796 B.n1 585
R732 B.n797 B.n796 585
R733 B.n795 B.n794 585
R734 B.n795 B.n8 585
R735 B.n793 B.n9 585
R736 B.n12 B.n9 585
R737 B.n792 B.n791 585
R738 B.n791 B.n790 585
R739 B.n11 B.n10 585
R740 B.n789 B.n11 585
R741 B.n787 B.n786 585
R742 B.n788 B.n787 585
R743 B.n785 B.n17 585
R744 B.n17 B.n16 585
R745 B.n784 B.n783 585
R746 B.n783 B.n782 585
R747 B.n19 B.n18 585
R748 B.n781 B.n19 585
R749 B.n779 B.n778 585
R750 B.n780 B.n779 585
R751 B.n777 B.n24 585
R752 B.n24 B.n23 585
R753 B.n776 B.n775 585
R754 B.n775 B.n774 585
R755 B.n26 B.n25 585
R756 B.n773 B.n26 585
R757 B.n771 B.n770 585
R758 B.n772 B.n771 585
R759 B.n769 B.n30 585
R760 B.n33 B.n30 585
R761 B.n768 B.n767 585
R762 B.n767 B.n766 585
R763 B.n32 B.n31 585
R764 B.n765 B.n32 585
R765 B.n763 B.n762 585
R766 B.n764 B.n763 585
R767 B.n761 B.n38 585
R768 B.n38 B.n37 585
R769 B.n760 B.n759 585
R770 B.n759 B.n758 585
R771 B.n40 B.n39 585
R772 B.n757 B.n40 585
R773 B.n755 B.n754 585
R774 B.n756 B.n755 585
R775 B.n753 B.n44 585
R776 B.n47 B.n44 585
R777 B.n752 B.n751 585
R778 B.n751 B.n750 585
R779 B.n46 B.n45 585
R780 B.n749 B.n46 585
R781 B.n747 B.n746 585
R782 B.n748 B.n747 585
R783 B.n745 B.n52 585
R784 B.n52 B.n51 585
R785 B.n744 B.n743 585
R786 B.n743 B.n742 585
R787 B.n54 B.n53 585
R788 B.n741 B.n54 585
R789 B.n739 B.n738 585
R790 B.n740 B.n739 585
R791 B.n737 B.n59 585
R792 B.n59 B.n58 585
R793 B.n736 B.n735 585
R794 B.n735 B.n734 585
R795 B.n61 B.n60 585
R796 B.n733 B.n61 585
R797 B.n731 B.n730 585
R798 B.n732 B.n731 585
R799 B.n729 B.n66 585
R800 B.n66 B.n65 585
R801 B.n728 B.n727 585
R802 B.n727 B.n726 585
R803 B.n68 B.n67 585
R804 B.n725 B.n68 585
R805 B.n723 B.n722 585
R806 B.n724 B.n723 585
R807 B.n721 B.n73 585
R808 B.n73 B.n72 585
R809 B.n720 B.n719 585
R810 B.n719 B.n718 585
R811 B.n75 B.n74 585
R812 B.n717 B.n75 585
R813 B.n715 B.n714 585
R814 B.n716 B.n715 585
R815 B.n713 B.n80 585
R816 B.n80 B.n79 585
R817 B.n712 B.n711 585
R818 B.n711 B.n710 585
R819 B.n82 B.n81 585
R820 B.n709 B.n82 585
R821 B.n707 B.n706 585
R822 B.n708 B.n707 585
R823 B.n705 B.n87 585
R824 B.n87 B.n86 585
R825 B.n704 B.n703 585
R826 B.n703 B.n702 585
R827 B.n89 B.n88 585
R828 B.n701 B.n89 585
R829 B.n699 B.n698 585
R830 B.n700 B.n699 585
R831 B.n697 B.n94 585
R832 B.n94 B.n93 585
R833 B.n696 B.n695 585
R834 B.n695 B.n694 585
R835 B.n96 B.n95 585
R836 B.n693 B.n96 585
R837 B.n691 B.n690 585
R838 B.n692 B.n691 585
R839 B.n689 B.n101 585
R840 B.n101 B.n100 585
R841 B.n688 B.n687 585
R842 B.n687 B.n686 585
R843 B.n103 B.n102 585
R844 B.n685 B.n103 585
R845 B.n683 B.n682 585
R846 B.n684 B.n683 585
R847 B.n681 B.n108 585
R848 B.n108 B.n107 585
R849 B.n680 B.n679 585
R850 B.n679 B.n678 585
R851 B.n800 B.n799 585
R852 B.n798 B.n2 585
R853 B.n679 B.n110 497.305
R854 B.n675 B.n111 497.305
R855 B.n414 B.n320 497.305
R856 B.n416 B.n318 497.305
R857 B.n677 B.n676 256.663
R858 B.n677 B.n128 256.663
R859 B.n677 B.n127 256.663
R860 B.n677 B.n126 256.663
R861 B.n677 B.n125 256.663
R862 B.n677 B.n124 256.663
R863 B.n677 B.n123 256.663
R864 B.n677 B.n122 256.663
R865 B.n677 B.n121 256.663
R866 B.n677 B.n120 256.663
R867 B.n677 B.n119 256.663
R868 B.n677 B.n118 256.663
R869 B.n677 B.n117 256.663
R870 B.n677 B.n116 256.663
R871 B.n677 B.n115 256.663
R872 B.n677 B.n114 256.663
R873 B.n677 B.n113 256.663
R874 B.n677 B.n112 256.663
R875 B.n343 B.n319 256.663
R876 B.n349 B.n319 256.663
R877 B.n351 B.n319 256.663
R878 B.n357 B.n319 256.663
R879 B.n359 B.n319 256.663
R880 B.n365 B.n319 256.663
R881 B.n367 B.n319 256.663
R882 B.n373 B.n319 256.663
R883 B.n375 B.n319 256.663
R884 B.n381 B.n319 256.663
R885 B.n383 B.n319 256.663
R886 B.n390 B.n319 256.663
R887 B.n392 B.n319 256.663
R888 B.n398 B.n319 256.663
R889 B.n400 B.n319 256.663
R890 B.n406 B.n319 256.663
R891 B.n409 B.n319 256.663
R892 B.n802 B.n801 256.663
R893 B.n132 B.t14 229.993
R894 B.n130 B.t21 229.993
R895 B.n328 B.t18 229.993
R896 B.n334 B.t10 229.993
R897 B.n130 B.t22 177.971
R898 B.n328 B.t20 177.971
R899 B.n132 B.t16 177.971
R900 B.n334 B.t13 177.971
R901 B.n136 B.n135 163.367
R902 B.n140 B.n139 163.367
R903 B.n144 B.n143 163.367
R904 B.n148 B.n147 163.367
R905 B.n152 B.n151 163.367
R906 B.n156 B.n155 163.367
R907 B.n161 B.n160 163.367
R908 B.n165 B.n164 163.367
R909 B.n169 B.n168 163.367
R910 B.n173 B.n172 163.367
R911 B.n177 B.n176 163.367
R912 B.n182 B.n181 163.367
R913 B.n186 B.n185 163.367
R914 B.n190 B.n189 163.367
R915 B.n194 B.n193 163.367
R916 B.n198 B.n197 163.367
R917 B.n200 B.n129 163.367
R918 B.n414 B.n314 163.367
R919 B.n422 B.n314 163.367
R920 B.n422 B.n312 163.367
R921 B.n426 B.n312 163.367
R922 B.n426 B.n305 163.367
R923 B.n434 B.n305 163.367
R924 B.n434 B.n303 163.367
R925 B.n438 B.n303 163.367
R926 B.n438 B.n298 163.367
R927 B.n446 B.n298 163.367
R928 B.n446 B.n296 163.367
R929 B.n450 B.n296 163.367
R930 B.n450 B.n290 163.367
R931 B.n458 B.n290 163.367
R932 B.n458 B.n288 163.367
R933 B.n462 B.n288 163.367
R934 B.n462 B.n281 163.367
R935 B.n470 B.n281 163.367
R936 B.n470 B.n279 163.367
R937 B.n474 B.n279 163.367
R938 B.n474 B.n274 163.367
R939 B.n482 B.n274 163.367
R940 B.n482 B.n272 163.367
R941 B.n486 B.n272 163.367
R942 B.n486 B.n266 163.367
R943 B.n494 B.n266 163.367
R944 B.n494 B.n264 163.367
R945 B.n498 B.n264 163.367
R946 B.n498 B.n258 163.367
R947 B.n506 B.n258 163.367
R948 B.n506 B.n256 163.367
R949 B.n510 B.n256 163.367
R950 B.n510 B.n250 163.367
R951 B.n518 B.n250 163.367
R952 B.n518 B.n248 163.367
R953 B.n522 B.n248 163.367
R954 B.n522 B.n243 163.367
R955 B.n531 B.n243 163.367
R956 B.n531 B.n241 163.367
R957 B.n535 B.n241 163.367
R958 B.n535 B.n235 163.367
R959 B.n543 B.n235 163.367
R960 B.n543 B.n233 163.367
R961 B.n547 B.n233 163.367
R962 B.n547 B.n228 163.367
R963 B.n556 B.n228 163.367
R964 B.n556 B.n226 163.367
R965 B.n560 B.n226 163.367
R966 B.n560 B.n220 163.367
R967 B.n568 B.n220 163.367
R968 B.n568 B.n218 163.367
R969 B.n572 B.n218 163.367
R970 B.n572 B.n212 163.367
R971 B.n580 B.n212 163.367
R972 B.n580 B.n210 163.367
R973 B.n585 B.n210 163.367
R974 B.n585 B.n204 163.367
R975 B.n593 B.n204 163.367
R976 B.n594 B.n593 163.367
R977 B.n594 B.n5 163.367
R978 B.n6 B.n5 163.367
R979 B.n7 B.n6 163.367
R980 B.n600 B.n7 163.367
R981 B.n601 B.n600 163.367
R982 B.n601 B.n13 163.367
R983 B.n14 B.n13 163.367
R984 B.n15 B.n14 163.367
R985 B.n606 B.n15 163.367
R986 B.n606 B.n20 163.367
R987 B.n21 B.n20 163.367
R988 B.n22 B.n21 163.367
R989 B.n611 B.n22 163.367
R990 B.n611 B.n27 163.367
R991 B.n28 B.n27 163.367
R992 B.n29 B.n28 163.367
R993 B.n616 B.n29 163.367
R994 B.n616 B.n34 163.367
R995 B.n35 B.n34 163.367
R996 B.n36 B.n35 163.367
R997 B.n621 B.n36 163.367
R998 B.n621 B.n41 163.367
R999 B.n42 B.n41 163.367
R1000 B.n43 B.n42 163.367
R1001 B.n626 B.n43 163.367
R1002 B.n626 B.n48 163.367
R1003 B.n49 B.n48 163.367
R1004 B.n50 B.n49 163.367
R1005 B.n631 B.n50 163.367
R1006 B.n631 B.n55 163.367
R1007 B.n56 B.n55 163.367
R1008 B.n57 B.n56 163.367
R1009 B.n636 B.n57 163.367
R1010 B.n636 B.n62 163.367
R1011 B.n63 B.n62 163.367
R1012 B.n64 B.n63 163.367
R1013 B.n641 B.n64 163.367
R1014 B.n641 B.n69 163.367
R1015 B.n70 B.n69 163.367
R1016 B.n71 B.n70 163.367
R1017 B.n646 B.n71 163.367
R1018 B.n646 B.n76 163.367
R1019 B.n77 B.n76 163.367
R1020 B.n78 B.n77 163.367
R1021 B.n651 B.n78 163.367
R1022 B.n651 B.n83 163.367
R1023 B.n84 B.n83 163.367
R1024 B.n85 B.n84 163.367
R1025 B.n656 B.n85 163.367
R1026 B.n656 B.n90 163.367
R1027 B.n91 B.n90 163.367
R1028 B.n92 B.n91 163.367
R1029 B.n661 B.n92 163.367
R1030 B.n661 B.n97 163.367
R1031 B.n98 B.n97 163.367
R1032 B.n99 B.n98 163.367
R1033 B.n666 B.n99 163.367
R1034 B.n666 B.n104 163.367
R1035 B.n105 B.n104 163.367
R1036 B.n106 B.n105 163.367
R1037 B.n671 B.n106 163.367
R1038 B.n671 B.n111 163.367
R1039 B.n344 B.n342 163.367
R1040 B.n348 B.n342 163.367
R1041 B.n352 B.n350 163.367
R1042 B.n356 B.n340 163.367
R1043 B.n360 B.n358 163.367
R1044 B.n364 B.n338 163.367
R1045 B.n368 B.n366 163.367
R1046 B.n372 B.n333 163.367
R1047 B.n376 B.n374 163.367
R1048 B.n380 B.n331 163.367
R1049 B.n384 B.n382 163.367
R1050 B.n389 B.n327 163.367
R1051 B.n393 B.n391 163.367
R1052 B.n397 B.n325 163.367
R1053 B.n401 B.n399 163.367
R1054 B.n405 B.n323 163.367
R1055 B.n408 B.n407 163.367
R1056 B.n410 B.n320 163.367
R1057 B.n416 B.n316 163.367
R1058 B.n420 B.n316 163.367
R1059 B.n420 B.n310 163.367
R1060 B.n428 B.n310 163.367
R1061 B.n428 B.n308 163.367
R1062 B.n432 B.n308 163.367
R1063 B.n432 B.n302 163.367
R1064 B.n440 B.n302 163.367
R1065 B.n440 B.n300 163.367
R1066 B.n444 B.n300 163.367
R1067 B.n444 B.n294 163.367
R1068 B.n452 B.n294 163.367
R1069 B.n452 B.n292 163.367
R1070 B.n456 B.n292 163.367
R1071 B.n456 B.n286 163.367
R1072 B.n464 B.n286 163.367
R1073 B.n464 B.n284 163.367
R1074 B.n468 B.n284 163.367
R1075 B.n468 B.n278 163.367
R1076 B.n476 B.n278 163.367
R1077 B.n476 B.n276 163.367
R1078 B.n480 B.n276 163.367
R1079 B.n480 B.n270 163.367
R1080 B.n488 B.n270 163.367
R1081 B.n488 B.n268 163.367
R1082 B.n492 B.n268 163.367
R1083 B.n492 B.n262 163.367
R1084 B.n500 B.n262 163.367
R1085 B.n500 B.n260 163.367
R1086 B.n504 B.n260 163.367
R1087 B.n504 B.n254 163.367
R1088 B.n512 B.n254 163.367
R1089 B.n512 B.n252 163.367
R1090 B.n516 B.n252 163.367
R1091 B.n516 B.n246 163.367
R1092 B.n525 B.n246 163.367
R1093 B.n525 B.n244 163.367
R1094 B.n529 B.n244 163.367
R1095 B.n529 B.n239 163.367
R1096 B.n537 B.n239 163.367
R1097 B.n537 B.n237 163.367
R1098 B.n541 B.n237 163.367
R1099 B.n541 B.n231 163.367
R1100 B.n550 B.n231 163.367
R1101 B.n550 B.n229 163.367
R1102 B.n554 B.n229 163.367
R1103 B.n554 B.n224 163.367
R1104 B.n562 B.n224 163.367
R1105 B.n562 B.n222 163.367
R1106 B.n566 B.n222 163.367
R1107 B.n566 B.n216 163.367
R1108 B.n574 B.n216 163.367
R1109 B.n574 B.n214 163.367
R1110 B.n578 B.n214 163.367
R1111 B.n578 B.n208 163.367
R1112 B.n587 B.n208 163.367
R1113 B.n587 B.n206 163.367
R1114 B.n591 B.n206 163.367
R1115 B.n591 B.n3 163.367
R1116 B.n800 B.n3 163.367
R1117 B.n796 B.n2 163.367
R1118 B.n796 B.n795 163.367
R1119 B.n795 B.n9 163.367
R1120 B.n791 B.n9 163.367
R1121 B.n791 B.n11 163.367
R1122 B.n787 B.n11 163.367
R1123 B.n787 B.n17 163.367
R1124 B.n783 B.n17 163.367
R1125 B.n783 B.n19 163.367
R1126 B.n779 B.n19 163.367
R1127 B.n779 B.n24 163.367
R1128 B.n775 B.n24 163.367
R1129 B.n775 B.n26 163.367
R1130 B.n771 B.n26 163.367
R1131 B.n771 B.n30 163.367
R1132 B.n767 B.n30 163.367
R1133 B.n767 B.n32 163.367
R1134 B.n763 B.n32 163.367
R1135 B.n763 B.n38 163.367
R1136 B.n759 B.n38 163.367
R1137 B.n759 B.n40 163.367
R1138 B.n755 B.n40 163.367
R1139 B.n755 B.n44 163.367
R1140 B.n751 B.n44 163.367
R1141 B.n751 B.n46 163.367
R1142 B.n747 B.n46 163.367
R1143 B.n747 B.n52 163.367
R1144 B.n743 B.n52 163.367
R1145 B.n743 B.n54 163.367
R1146 B.n739 B.n54 163.367
R1147 B.n739 B.n59 163.367
R1148 B.n735 B.n59 163.367
R1149 B.n735 B.n61 163.367
R1150 B.n731 B.n61 163.367
R1151 B.n731 B.n66 163.367
R1152 B.n727 B.n66 163.367
R1153 B.n727 B.n68 163.367
R1154 B.n723 B.n68 163.367
R1155 B.n723 B.n73 163.367
R1156 B.n719 B.n73 163.367
R1157 B.n719 B.n75 163.367
R1158 B.n715 B.n75 163.367
R1159 B.n715 B.n80 163.367
R1160 B.n711 B.n80 163.367
R1161 B.n711 B.n82 163.367
R1162 B.n707 B.n82 163.367
R1163 B.n707 B.n87 163.367
R1164 B.n703 B.n87 163.367
R1165 B.n703 B.n89 163.367
R1166 B.n699 B.n89 163.367
R1167 B.n699 B.n94 163.367
R1168 B.n695 B.n94 163.367
R1169 B.n695 B.n96 163.367
R1170 B.n691 B.n96 163.367
R1171 B.n691 B.n101 163.367
R1172 B.n687 B.n101 163.367
R1173 B.n687 B.n103 163.367
R1174 B.n683 B.n103 163.367
R1175 B.n683 B.n108 163.367
R1176 B.n679 B.n108 163.367
R1177 B.n415 B.n319 162.167
R1178 B.n678 B.n677 162.167
R1179 B.n131 B.t23 120.566
R1180 B.n329 B.t19 120.566
R1181 B.n133 B.t17 120.566
R1182 B.n335 B.t12 120.566
R1183 B.n415 B.n315 97.5869
R1184 B.n421 B.n315 97.5869
R1185 B.n421 B.n311 97.5869
R1186 B.n427 B.n311 97.5869
R1187 B.n427 B.n306 97.5869
R1188 B.n433 B.n306 97.5869
R1189 B.n433 B.n307 97.5869
R1190 B.n439 B.n299 97.5869
R1191 B.n445 B.n299 97.5869
R1192 B.n445 B.n295 97.5869
R1193 B.n451 B.n295 97.5869
R1194 B.n451 B.n291 97.5869
R1195 B.n457 B.n291 97.5869
R1196 B.n457 B.n287 97.5869
R1197 B.n463 B.n287 97.5869
R1198 B.n463 B.n282 97.5869
R1199 B.n469 B.n282 97.5869
R1200 B.n469 B.n283 97.5869
R1201 B.n475 B.n275 97.5869
R1202 B.n481 B.n275 97.5869
R1203 B.n481 B.n271 97.5869
R1204 B.n487 B.n271 97.5869
R1205 B.n487 B.n267 97.5869
R1206 B.n493 B.n267 97.5869
R1207 B.n493 B.n263 97.5869
R1208 B.n499 B.n263 97.5869
R1209 B.n505 B.n259 97.5869
R1210 B.n505 B.n255 97.5869
R1211 B.n511 B.n255 97.5869
R1212 B.n511 B.n251 97.5869
R1213 B.n517 B.n251 97.5869
R1214 B.n517 B.n247 97.5869
R1215 B.n524 B.n247 97.5869
R1216 B.n524 B.n523 97.5869
R1217 B.n530 B.n240 97.5869
R1218 B.n536 B.n240 97.5869
R1219 B.n536 B.n236 97.5869
R1220 B.n542 B.n236 97.5869
R1221 B.n542 B.n232 97.5869
R1222 B.n549 B.n232 97.5869
R1223 B.n549 B.n548 97.5869
R1224 B.n555 B.n225 97.5869
R1225 B.n561 B.n225 97.5869
R1226 B.n561 B.n221 97.5869
R1227 B.n567 B.n221 97.5869
R1228 B.n567 B.n217 97.5869
R1229 B.n573 B.n217 97.5869
R1230 B.n573 B.n213 97.5869
R1231 B.n579 B.n213 97.5869
R1232 B.n586 B.n209 97.5869
R1233 B.n586 B.n205 97.5869
R1234 B.n592 B.n205 97.5869
R1235 B.n592 B.n4 97.5869
R1236 B.n799 B.n4 97.5869
R1237 B.n799 B.n798 97.5869
R1238 B.n798 B.n797 97.5869
R1239 B.n797 B.n8 97.5869
R1240 B.n12 B.n8 97.5869
R1241 B.n790 B.n12 97.5869
R1242 B.n790 B.n789 97.5869
R1243 B.n788 B.n16 97.5869
R1244 B.n782 B.n16 97.5869
R1245 B.n782 B.n781 97.5869
R1246 B.n781 B.n780 97.5869
R1247 B.n780 B.n23 97.5869
R1248 B.n774 B.n23 97.5869
R1249 B.n774 B.n773 97.5869
R1250 B.n773 B.n772 97.5869
R1251 B.n766 B.n33 97.5869
R1252 B.n766 B.n765 97.5869
R1253 B.n765 B.n764 97.5869
R1254 B.n764 B.n37 97.5869
R1255 B.n758 B.n37 97.5869
R1256 B.n758 B.n757 97.5869
R1257 B.n757 B.n756 97.5869
R1258 B.n750 B.n47 97.5869
R1259 B.n750 B.n749 97.5869
R1260 B.n749 B.n748 97.5869
R1261 B.n748 B.n51 97.5869
R1262 B.n742 B.n51 97.5869
R1263 B.n742 B.n741 97.5869
R1264 B.n741 B.n740 97.5869
R1265 B.n740 B.n58 97.5869
R1266 B.n734 B.n733 97.5869
R1267 B.n733 B.n732 97.5869
R1268 B.n732 B.n65 97.5869
R1269 B.n726 B.n65 97.5869
R1270 B.n726 B.n725 97.5869
R1271 B.n725 B.n724 97.5869
R1272 B.n724 B.n72 97.5869
R1273 B.n718 B.n72 97.5869
R1274 B.n717 B.n716 97.5869
R1275 B.n716 B.n79 97.5869
R1276 B.n710 B.n79 97.5869
R1277 B.n710 B.n709 97.5869
R1278 B.n709 B.n708 97.5869
R1279 B.n708 B.n86 97.5869
R1280 B.n702 B.n86 97.5869
R1281 B.n702 B.n701 97.5869
R1282 B.n701 B.n700 97.5869
R1283 B.n700 B.n93 97.5869
R1284 B.n694 B.n93 97.5869
R1285 B.n693 B.n692 97.5869
R1286 B.n692 B.n100 97.5869
R1287 B.n686 B.n100 97.5869
R1288 B.n686 B.n685 97.5869
R1289 B.n685 B.n684 97.5869
R1290 B.n684 B.n107 97.5869
R1291 B.n678 B.n107 97.5869
R1292 B.n530 B.t9 84.6711
R1293 B.n756 B.t7 84.6711
R1294 B.n548 B.t3 81.8009
R1295 B.n33 B.t6 81.8009
R1296 B.n307 B.t11 78.9307
R1297 B.t15 B.n693 78.9307
R1298 B.n112 B.n110 71.676
R1299 B.n136 B.n113 71.676
R1300 B.n140 B.n114 71.676
R1301 B.n144 B.n115 71.676
R1302 B.n148 B.n116 71.676
R1303 B.n152 B.n117 71.676
R1304 B.n156 B.n118 71.676
R1305 B.n161 B.n119 71.676
R1306 B.n165 B.n120 71.676
R1307 B.n169 B.n121 71.676
R1308 B.n173 B.n122 71.676
R1309 B.n177 B.n123 71.676
R1310 B.n182 B.n124 71.676
R1311 B.n186 B.n125 71.676
R1312 B.n190 B.n126 71.676
R1313 B.n194 B.n127 71.676
R1314 B.n198 B.n128 71.676
R1315 B.n676 B.n129 71.676
R1316 B.n676 B.n675 71.676
R1317 B.n200 B.n128 71.676
R1318 B.n197 B.n127 71.676
R1319 B.n193 B.n126 71.676
R1320 B.n189 B.n125 71.676
R1321 B.n185 B.n124 71.676
R1322 B.n181 B.n123 71.676
R1323 B.n176 B.n122 71.676
R1324 B.n172 B.n121 71.676
R1325 B.n168 B.n120 71.676
R1326 B.n164 B.n119 71.676
R1327 B.n160 B.n118 71.676
R1328 B.n155 B.n117 71.676
R1329 B.n151 B.n116 71.676
R1330 B.n147 B.n115 71.676
R1331 B.n143 B.n114 71.676
R1332 B.n139 B.n113 71.676
R1333 B.n135 B.n112 71.676
R1334 B.n343 B.n318 71.676
R1335 B.n349 B.n348 71.676
R1336 B.n352 B.n351 71.676
R1337 B.n357 B.n356 71.676
R1338 B.n360 B.n359 71.676
R1339 B.n365 B.n364 71.676
R1340 B.n368 B.n367 71.676
R1341 B.n373 B.n372 71.676
R1342 B.n376 B.n375 71.676
R1343 B.n381 B.n380 71.676
R1344 B.n384 B.n383 71.676
R1345 B.n390 B.n389 71.676
R1346 B.n393 B.n392 71.676
R1347 B.n398 B.n397 71.676
R1348 B.n401 B.n400 71.676
R1349 B.n406 B.n405 71.676
R1350 B.n409 B.n408 71.676
R1351 B.n344 B.n343 71.676
R1352 B.n350 B.n349 71.676
R1353 B.n351 B.n340 71.676
R1354 B.n358 B.n357 71.676
R1355 B.n359 B.n338 71.676
R1356 B.n366 B.n365 71.676
R1357 B.n367 B.n333 71.676
R1358 B.n374 B.n373 71.676
R1359 B.n375 B.n331 71.676
R1360 B.n382 B.n381 71.676
R1361 B.n383 B.n327 71.676
R1362 B.n391 B.n390 71.676
R1363 B.n392 B.n325 71.676
R1364 B.n399 B.n398 71.676
R1365 B.n400 B.n323 71.676
R1366 B.n407 B.n406 71.676
R1367 B.n410 B.n409 71.676
R1368 B.n801 B.n800 71.676
R1369 B.n801 B.n2 71.676
R1370 B.n283 B.t5 70.3201
R1371 B.t8 B.n717 70.3201
R1372 B.n158 B.n133 59.5399
R1373 B.n179 B.n131 59.5399
R1374 B.n387 B.n329 59.5399
R1375 B.n336 B.n335 59.5399
R1376 B.n133 B.n132 57.4066
R1377 B.n131 B.n130 57.4066
R1378 B.n329 B.n328 57.4066
R1379 B.n335 B.n334 57.4066
R1380 B.t2 B.n259 55.9692
R1381 B.t1 B.n58 55.9692
R1382 B.n579 B.t4 53.099
R1383 B.t0 B.n788 53.099
R1384 B.t4 B.n209 44.4884
R1385 B.n789 B.t0 44.4884
R1386 B.n499 B.t2 41.6182
R1387 B.n734 B.t1 41.6182
R1388 B.n417 B.n317 32.3127
R1389 B.n413 B.n412 32.3127
R1390 B.n674 B.n673 32.3127
R1391 B.n680 B.n109 32.3127
R1392 B.n475 B.t5 27.2673
R1393 B.n718 B.t8 27.2673
R1394 B.n439 B.t11 18.6567
R1395 B.n694 B.t15 18.6567
R1396 B B.n802 18.0485
R1397 B.n555 B.t3 15.7865
R1398 B.n772 B.t6 15.7865
R1399 B.n523 B.t9 12.9164
R1400 B.n47 B.t7 12.9164
R1401 B.n418 B.n417 10.6151
R1402 B.n419 B.n418 10.6151
R1403 B.n419 B.n309 10.6151
R1404 B.n429 B.n309 10.6151
R1405 B.n430 B.n429 10.6151
R1406 B.n431 B.n430 10.6151
R1407 B.n431 B.n301 10.6151
R1408 B.n441 B.n301 10.6151
R1409 B.n442 B.n441 10.6151
R1410 B.n443 B.n442 10.6151
R1411 B.n443 B.n293 10.6151
R1412 B.n453 B.n293 10.6151
R1413 B.n454 B.n453 10.6151
R1414 B.n455 B.n454 10.6151
R1415 B.n455 B.n285 10.6151
R1416 B.n465 B.n285 10.6151
R1417 B.n466 B.n465 10.6151
R1418 B.n467 B.n466 10.6151
R1419 B.n467 B.n277 10.6151
R1420 B.n477 B.n277 10.6151
R1421 B.n478 B.n477 10.6151
R1422 B.n479 B.n478 10.6151
R1423 B.n479 B.n269 10.6151
R1424 B.n489 B.n269 10.6151
R1425 B.n490 B.n489 10.6151
R1426 B.n491 B.n490 10.6151
R1427 B.n491 B.n261 10.6151
R1428 B.n501 B.n261 10.6151
R1429 B.n502 B.n501 10.6151
R1430 B.n503 B.n502 10.6151
R1431 B.n503 B.n253 10.6151
R1432 B.n513 B.n253 10.6151
R1433 B.n514 B.n513 10.6151
R1434 B.n515 B.n514 10.6151
R1435 B.n515 B.n245 10.6151
R1436 B.n526 B.n245 10.6151
R1437 B.n527 B.n526 10.6151
R1438 B.n528 B.n527 10.6151
R1439 B.n528 B.n238 10.6151
R1440 B.n538 B.n238 10.6151
R1441 B.n539 B.n538 10.6151
R1442 B.n540 B.n539 10.6151
R1443 B.n540 B.n230 10.6151
R1444 B.n551 B.n230 10.6151
R1445 B.n552 B.n551 10.6151
R1446 B.n553 B.n552 10.6151
R1447 B.n553 B.n223 10.6151
R1448 B.n563 B.n223 10.6151
R1449 B.n564 B.n563 10.6151
R1450 B.n565 B.n564 10.6151
R1451 B.n565 B.n215 10.6151
R1452 B.n575 B.n215 10.6151
R1453 B.n576 B.n575 10.6151
R1454 B.n577 B.n576 10.6151
R1455 B.n577 B.n207 10.6151
R1456 B.n588 B.n207 10.6151
R1457 B.n589 B.n588 10.6151
R1458 B.n590 B.n589 10.6151
R1459 B.n590 B.n0 10.6151
R1460 B.n345 B.n317 10.6151
R1461 B.n346 B.n345 10.6151
R1462 B.n347 B.n346 10.6151
R1463 B.n347 B.n341 10.6151
R1464 B.n353 B.n341 10.6151
R1465 B.n354 B.n353 10.6151
R1466 B.n355 B.n354 10.6151
R1467 B.n355 B.n339 10.6151
R1468 B.n361 B.n339 10.6151
R1469 B.n362 B.n361 10.6151
R1470 B.n363 B.n362 10.6151
R1471 B.n363 B.n337 10.6151
R1472 B.n370 B.n369 10.6151
R1473 B.n371 B.n370 10.6151
R1474 B.n371 B.n332 10.6151
R1475 B.n377 B.n332 10.6151
R1476 B.n378 B.n377 10.6151
R1477 B.n379 B.n378 10.6151
R1478 B.n379 B.n330 10.6151
R1479 B.n385 B.n330 10.6151
R1480 B.n386 B.n385 10.6151
R1481 B.n388 B.n326 10.6151
R1482 B.n394 B.n326 10.6151
R1483 B.n395 B.n394 10.6151
R1484 B.n396 B.n395 10.6151
R1485 B.n396 B.n324 10.6151
R1486 B.n402 B.n324 10.6151
R1487 B.n403 B.n402 10.6151
R1488 B.n404 B.n403 10.6151
R1489 B.n404 B.n322 10.6151
R1490 B.n322 B.n321 10.6151
R1491 B.n411 B.n321 10.6151
R1492 B.n412 B.n411 10.6151
R1493 B.n413 B.n313 10.6151
R1494 B.n423 B.n313 10.6151
R1495 B.n424 B.n423 10.6151
R1496 B.n425 B.n424 10.6151
R1497 B.n425 B.n304 10.6151
R1498 B.n435 B.n304 10.6151
R1499 B.n436 B.n435 10.6151
R1500 B.n437 B.n436 10.6151
R1501 B.n437 B.n297 10.6151
R1502 B.n447 B.n297 10.6151
R1503 B.n448 B.n447 10.6151
R1504 B.n449 B.n448 10.6151
R1505 B.n449 B.n289 10.6151
R1506 B.n459 B.n289 10.6151
R1507 B.n460 B.n459 10.6151
R1508 B.n461 B.n460 10.6151
R1509 B.n461 B.n280 10.6151
R1510 B.n471 B.n280 10.6151
R1511 B.n472 B.n471 10.6151
R1512 B.n473 B.n472 10.6151
R1513 B.n473 B.n273 10.6151
R1514 B.n483 B.n273 10.6151
R1515 B.n484 B.n483 10.6151
R1516 B.n485 B.n484 10.6151
R1517 B.n485 B.n265 10.6151
R1518 B.n495 B.n265 10.6151
R1519 B.n496 B.n495 10.6151
R1520 B.n497 B.n496 10.6151
R1521 B.n497 B.n257 10.6151
R1522 B.n507 B.n257 10.6151
R1523 B.n508 B.n507 10.6151
R1524 B.n509 B.n508 10.6151
R1525 B.n509 B.n249 10.6151
R1526 B.n519 B.n249 10.6151
R1527 B.n520 B.n519 10.6151
R1528 B.n521 B.n520 10.6151
R1529 B.n521 B.n242 10.6151
R1530 B.n532 B.n242 10.6151
R1531 B.n533 B.n532 10.6151
R1532 B.n534 B.n533 10.6151
R1533 B.n534 B.n234 10.6151
R1534 B.n544 B.n234 10.6151
R1535 B.n545 B.n544 10.6151
R1536 B.n546 B.n545 10.6151
R1537 B.n546 B.n227 10.6151
R1538 B.n557 B.n227 10.6151
R1539 B.n558 B.n557 10.6151
R1540 B.n559 B.n558 10.6151
R1541 B.n559 B.n219 10.6151
R1542 B.n569 B.n219 10.6151
R1543 B.n570 B.n569 10.6151
R1544 B.n571 B.n570 10.6151
R1545 B.n571 B.n211 10.6151
R1546 B.n581 B.n211 10.6151
R1547 B.n582 B.n581 10.6151
R1548 B.n584 B.n582 10.6151
R1549 B.n584 B.n583 10.6151
R1550 B.n583 B.n203 10.6151
R1551 B.n595 B.n203 10.6151
R1552 B.n596 B.n595 10.6151
R1553 B.n597 B.n596 10.6151
R1554 B.n598 B.n597 10.6151
R1555 B.n599 B.n598 10.6151
R1556 B.n602 B.n599 10.6151
R1557 B.n603 B.n602 10.6151
R1558 B.n604 B.n603 10.6151
R1559 B.n605 B.n604 10.6151
R1560 B.n607 B.n605 10.6151
R1561 B.n608 B.n607 10.6151
R1562 B.n609 B.n608 10.6151
R1563 B.n610 B.n609 10.6151
R1564 B.n612 B.n610 10.6151
R1565 B.n613 B.n612 10.6151
R1566 B.n614 B.n613 10.6151
R1567 B.n615 B.n614 10.6151
R1568 B.n617 B.n615 10.6151
R1569 B.n618 B.n617 10.6151
R1570 B.n619 B.n618 10.6151
R1571 B.n620 B.n619 10.6151
R1572 B.n622 B.n620 10.6151
R1573 B.n623 B.n622 10.6151
R1574 B.n624 B.n623 10.6151
R1575 B.n625 B.n624 10.6151
R1576 B.n627 B.n625 10.6151
R1577 B.n628 B.n627 10.6151
R1578 B.n629 B.n628 10.6151
R1579 B.n630 B.n629 10.6151
R1580 B.n632 B.n630 10.6151
R1581 B.n633 B.n632 10.6151
R1582 B.n634 B.n633 10.6151
R1583 B.n635 B.n634 10.6151
R1584 B.n637 B.n635 10.6151
R1585 B.n638 B.n637 10.6151
R1586 B.n639 B.n638 10.6151
R1587 B.n640 B.n639 10.6151
R1588 B.n642 B.n640 10.6151
R1589 B.n643 B.n642 10.6151
R1590 B.n644 B.n643 10.6151
R1591 B.n645 B.n644 10.6151
R1592 B.n647 B.n645 10.6151
R1593 B.n648 B.n647 10.6151
R1594 B.n649 B.n648 10.6151
R1595 B.n650 B.n649 10.6151
R1596 B.n652 B.n650 10.6151
R1597 B.n653 B.n652 10.6151
R1598 B.n654 B.n653 10.6151
R1599 B.n655 B.n654 10.6151
R1600 B.n657 B.n655 10.6151
R1601 B.n658 B.n657 10.6151
R1602 B.n659 B.n658 10.6151
R1603 B.n660 B.n659 10.6151
R1604 B.n662 B.n660 10.6151
R1605 B.n663 B.n662 10.6151
R1606 B.n664 B.n663 10.6151
R1607 B.n665 B.n664 10.6151
R1608 B.n667 B.n665 10.6151
R1609 B.n668 B.n667 10.6151
R1610 B.n669 B.n668 10.6151
R1611 B.n670 B.n669 10.6151
R1612 B.n672 B.n670 10.6151
R1613 B.n673 B.n672 10.6151
R1614 B.n794 B.n1 10.6151
R1615 B.n794 B.n793 10.6151
R1616 B.n793 B.n792 10.6151
R1617 B.n792 B.n10 10.6151
R1618 B.n786 B.n10 10.6151
R1619 B.n786 B.n785 10.6151
R1620 B.n785 B.n784 10.6151
R1621 B.n784 B.n18 10.6151
R1622 B.n778 B.n18 10.6151
R1623 B.n778 B.n777 10.6151
R1624 B.n777 B.n776 10.6151
R1625 B.n776 B.n25 10.6151
R1626 B.n770 B.n25 10.6151
R1627 B.n770 B.n769 10.6151
R1628 B.n769 B.n768 10.6151
R1629 B.n768 B.n31 10.6151
R1630 B.n762 B.n31 10.6151
R1631 B.n762 B.n761 10.6151
R1632 B.n761 B.n760 10.6151
R1633 B.n760 B.n39 10.6151
R1634 B.n754 B.n39 10.6151
R1635 B.n754 B.n753 10.6151
R1636 B.n753 B.n752 10.6151
R1637 B.n752 B.n45 10.6151
R1638 B.n746 B.n45 10.6151
R1639 B.n746 B.n745 10.6151
R1640 B.n745 B.n744 10.6151
R1641 B.n744 B.n53 10.6151
R1642 B.n738 B.n53 10.6151
R1643 B.n738 B.n737 10.6151
R1644 B.n737 B.n736 10.6151
R1645 B.n736 B.n60 10.6151
R1646 B.n730 B.n60 10.6151
R1647 B.n730 B.n729 10.6151
R1648 B.n729 B.n728 10.6151
R1649 B.n728 B.n67 10.6151
R1650 B.n722 B.n67 10.6151
R1651 B.n722 B.n721 10.6151
R1652 B.n721 B.n720 10.6151
R1653 B.n720 B.n74 10.6151
R1654 B.n714 B.n74 10.6151
R1655 B.n714 B.n713 10.6151
R1656 B.n713 B.n712 10.6151
R1657 B.n712 B.n81 10.6151
R1658 B.n706 B.n81 10.6151
R1659 B.n706 B.n705 10.6151
R1660 B.n705 B.n704 10.6151
R1661 B.n704 B.n88 10.6151
R1662 B.n698 B.n88 10.6151
R1663 B.n698 B.n697 10.6151
R1664 B.n697 B.n696 10.6151
R1665 B.n696 B.n95 10.6151
R1666 B.n690 B.n95 10.6151
R1667 B.n690 B.n689 10.6151
R1668 B.n689 B.n688 10.6151
R1669 B.n688 B.n102 10.6151
R1670 B.n682 B.n102 10.6151
R1671 B.n682 B.n681 10.6151
R1672 B.n681 B.n680 10.6151
R1673 B.n134 B.n109 10.6151
R1674 B.n137 B.n134 10.6151
R1675 B.n138 B.n137 10.6151
R1676 B.n141 B.n138 10.6151
R1677 B.n142 B.n141 10.6151
R1678 B.n145 B.n142 10.6151
R1679 B.n146 B.n145 10.6151
R1680 B.n149 B.n146 10.6151
R1681 B.n150 B.n149 10.6151
R1682 B.n153 B.n150 10.6151
R1683 B.n154 B.n153 10.6151
R1684 B.n157 B.n154 10.6151
R1685 B.n162 B.n159 10.6151
R1686 B.n163 B.n162 10.6151
R1687 B.n166 B.n163 10.6151
R1688 B.n167 B.n166 10.6151
R1689 B.n170 B.n167 10.6151
R1690 B.n171 B.n170 10.6151
R1691 B.n174 B.n171 10.6151
R1692 B.n175 B.n174 10.6151
R1693 B.n178 B.n175 10.6151
R1694 B.n183 B.n180 10.6151
R1695 B.n184 B.n183 10.6151
R1696 B.n187 B.n184 10.6151
R1697 B.n188 B.n187 10.6151
R1698 B.n191 B.n188 10.6151
R1699 B.n192 B.n191 10.6151
R1700 B.n195 B.n192 10.6151
R1701 B.n196 B.n195 10.6151
R1702 B.n199 B.n196 10.6151
R1703 B.n201 B.n199 10.6151
R1704 B.n202 B.n201 10.6151
R1705 B.n674 B.n202 10.6151
R1706 B.n337 B.n336 9.36635
R1707 B.n388 B.n387 9.36635
R1708 B.n158 B.n157 9.36635
R1709 B.n180 B.n179 9.36635
R1710 B.n802 B.n0 8.11757
R1711 B.n802 B.n1 8.11757
R1712 B.n369 B.n336 1.24928
R1713 B.n387 B.n386 1.24928
R1714 B.n159 B.n158 1.24928
R1715 B.n179 B.n178 1.24928
R1716 VP.n25 VP.n22 161.3
R1717 VP.n27 VP.n26 161.3
R1718 VP.n28 VP.n21 161.3
R1719 VP.n30 VP.n29 161.3
R1720 VP.n31 VP.n20 161.3
R1721 VP.n33 VP.n32 161.3
R1722 VP.n35 VP.n19 161.3
R1723 VP.n37 VP.n36 161.3
R1724 VP.n38 VP.n18 161.3
R1725 VP.n40 VP.n39 161.3
R1726 VP.n41 VP.n17 161.3
R1727 VP.n43 VP.n42 161.3
R1728 VP.n45 VP.n44 161.3
R1729 VP.n46 VP.n15 161.3
R1730 VP.n48 VP.n47 161.3
R1731 VP.n49 VP.n14 161.3
R1732 VP.n51 VP.n50 161.3
R1733 VP.n52 VP.n13 161.3
R1734 VP.n94 VP.n0 161.3
R1735 VP.n93 VP.n92 161.3
R1736 VP.n91 VP.n1 161.3
R1737 VP.n90 VP.n89 161.3
R1738 VP.n88 VP.n2 161.3
R1739 VP.n87 VP.n86 161.3
R1740 VP.n85 VP.n84 161.3
R1741 VP.n83 VP.n4 161.3
R1742 VP.n82 VP.n81 161.3
R1743 VP.n80 VP.n5 161.3
R1744 VP.n79 VP.n78 161.3
R1745 VP.n77 VP.n6 161.3
R1746 VP.n75 VP.n74 161.3
R1747 VP.n73 VP.n7 161.3
R1748 VP.n72 VP.n71 161.3
R1749 VP.n70 VP.n8 161.3
R1750 VP.n69 VP.n68 161.3
R1751 VP.n67 VP.n9 161.3
R1752 VP.n66 VP.n65 161.3
R1753 VP.n63 VP.n10 161.3
R1754 VP.n62 VP.n61 161.3
R1755 VP.n60 VP.n11 161.3
R1756 VP.n59 VP.n58 161.3
R1757 VP.n57 VP.n12 161.3
R1758 VP.n56 VP.n55 102.438
R1759 VP.n96 VP.n95 102.438
R1760 VP.n54 VP.n53 102.438
R1761 VP.n24 VP.n23 62.0711
R1762 VP.n62 VP.n11 56.5193
R1763 VP.n71 VP.n70 56.5193
R1764 VP.n82 VP.n5 56.5193
R1765 VP.n89 VP.n1 56.5193
R1766 VP.n47 VP.n14 56.5193
R1767 VP.n40 VP.n18 56.5193
R1768 VP.n29 VP.n28 56.5193
R1769 VP.n24 VP.t7 55.0181
R1770 VP.n55 VP.n54 45.9996
R1771 VP.n58 VP.n57 24.4675
R1772 VP.n58 VP.n11 24.4675
R1773 VP.n63 VP.n62 24.4675
R1774 VP.n65 VP.n63 24.4675
R1775 VP.n69 VP.n9 24.4675
R1776 VP.n70 VP.n69 24.4675
R1777 VP.n71 VP.n7 24.4675
R1778 VP.n75 VP.n7 24.4675
R1779 VP.n78 VP.n77 24.4675
R1780 VP.n78 VP.n5 24.4675
R1781 VP.n83 VP.n82 24.4675
R1782 VP.n84 VP.n83 24.4675
R1783 VP.n88 VP.n87 24.4675
R1784 VP.n89 VP.n88 24.4675
R1785 VP.n93 VP.n1 24.4675
R1786 VP.n94 VP.n93 24.4675
R1787 VP.n51 VP.n14 24.4675
R1788 VP.n52 VP.n51 24.4675
R1789 VP.n41 VP.n40 24.4675
R1790 VP.n42 VP.n41 24.4675
R1791 VP.n46 VP.n45 24.4675
R1792 VP.n47 VP.n46 24.4675
R1793 VP.n29 VP.n20 24.4675
R1794 VP.n33 VP.n20 24.4675
R1795 VP.n36 VP.n35 24.4675
R1796 VP.n36 VP.n18 24.4675
R1797 VP.n27 VP.n22 24.4675
R1798 VP.n28 VP.n27 24.4675
R1799 VP.n56 VP.t4 21.9013
R1800 VP.n64 VP.t5 21.9013
R1801 VP.n76 VP.t1 21.9013
R1802 VP.n3 VP.t9 21.9013
R1803 VP.n95 VP.t6 21.9013
R1804 VP.n53 VP.t2 21.9013
R1805 VP.n16 VP.t8 21.9013
R1806 VP.n34 VP.t0 21.9013
R1807 VP.n23 VP.t3 21.9013
R1808 VP.n65 VP.n64 14.1914
R1809 VP.n87 VP.n3 14.1914
R1810 VP.n45 VP.n16 14.1914
R1811 VP.n76 VP.n75 12.234
R1812 VP.n77 VP.n76 12.234
R1813 VP.n34 VP.n33 12.234
R1814 VP.n35 VP.n34 12.234
R1815 VP.n64 VP.n9 10.2766
R1816 VP.n84 VP.n3 10.2766
R1817 VP.n42 VP.n16 10.2766
R1818 VP.n23 VP.n22 10.2766
R1819 VP.n57 VP.n56 8.31928
R1820 VP.n95 VP.n94 8.31928
R1821 VP.n53 VP.n52 8.31928
R1822 VP.n25 VP.n24 6.95571
R1823 VP.n54 VP.n13 0.278367
R1824 VP.n55 VP.n12 0.278367
R1825 VP.n96 VP.n0 0.278367
R1826 VP.n26 VP.n25 0.189894
R1827 VP.n26 VP.n21 0.189894
R1828 VP.n30 VP.n21 0.189894
R1829 VP.n31 VP.n30 0.189894
R1830 VP.n32 VP.n31 0.189894
R1831 VP.n32 VP.n19 0.189894
R1832 VP.n37 VP.n19 0.189894
R1833 VP.n38 VP.n37 0.189894
R1834 VP.n39 VP.n38 0.189894
R1835 VP.n39 VP.n17 0.189894
R1836 VP.n43 VP.n17 0.189894
R1837 VP.n44 VP.n43 0.189894
R1838 VP.n44 VP.n15 0.189894
R1839 VP.n48 VP.n15 0.189894
R1840 VP.n49 VP.n48 0.189894
R1841 VP.n50 VP.n49 0.189894
R1842 VP.n50 VP.n13 0.189894
R1843 VP.n59 VP.n12 0.189894
R1844 VP.n60 VP.n59 0.189894
R1845 VP.n61 VP.n60 0.189894
R1846 VP.n61 VP.n10 0.189894
R1847 VP.n66 VP.n10 0.189894
R1848 VP.n67 VP.n66 0.189894
R1849 VP.n68 VP.n67 0.189894
R1850 VP.n68 VP.n8 0.189894
R1851 VP.n72 VP.n8 0.189894
R1852 VP.n73 VP.n72 0.189894
R1853 VP.n74 VP.n73 0.189894
R1854 VP.n74 VP.n6 0.189894
R1855 VP.n79 VP.n6 0.189894
R1856 VP.n80 VP.n79 0.189894
R1857 VP.n81 VP.n80 0.189894
R1858 VP.n81 VP.n4 0.189894
R1859 VP.n85 VP.n4 0.189894
R1860 VP.n86 VP.n85 0.189894
R1861 VP.n86 VP.n2 0.189894
R1862 VP.n90 VP.n2 0.189894
R1863 VP.n91 VP.n90 0.189894
R1864 VP.n92 VP.n91 0.189894
R1865 VP.n92 VP.n0 0.189894
R1866 VP VP.n96 0.153454
R1867 VDD1.n6 VDD1.n0 289.615
R1868 VDD1.n19 VDD1.n13 289.615
R1869 VDD1.n7 VDD1.n6 185
R1870 VDD1.n5 VDD1.n4 185
R1871 VDD1.n18 VDD1.n17 185
R1872 VDD1.n20 VDD1.n19 185
R1873 VDD1.n3 VDD1.t2 151.613
R1874 VDD1.n16 VDD1.t5 151.613
R1875 VDD1.n6 VDD1.n5 104.615
R1876 VDD1.n19 VDD1.n18 104.615
R1877 VDD1.n27 VDD1.n26 86.6237
R1878 VDD1.n12 VDD1.n11 84.7653
R1879 VDD1.n29 VDD1.n28 84.7652
R1880 VDD1.n25 VDD1.n24 84.7652
R1881 VDD1.n5 VDD1.t2 52.3082
R1882 VDD1.n18 VDD1.t5 52.3082
R1883 VDD1.n12 VDD1.n10 51.2219
R1884 VDD1.n25 VDD1.n23 51.2219
R1885 VDD1.n29 VDD1.n27 39.7552
R1886 VDD1.n4 VDD1.n3 15.3979
R1887 VDD1.n17 VDD1.n16 15.3979
R1888 VDD1.n7 VDD1.n2 12.8005
R1889 VDD1.n20 VDD1.n15 12.8005
R1890 VDD1.n8 VDD1.n0 12.0247
R1891 VDD1.n21 VDD1.n13 12.0247
R1892 VDD1.n10 VDD1.n9 9.45567
R1893 VDD1.n23 VDD1.n22 9.45567
R1894 VDD1.n9 VDD1.n8 9.3005
R1895 VDD1.n2 VDD1.n1 9.3005
R1896 VDD1.n22 VDD1.n21 9.3005
R1897 VDD1.n15 VDD1.n14 9.3005
R1898 VDD1.n28 VDD1.t1 8.28502
R1899 VDD1.n28 VDD1.t7 8.28502
R1900 VDD1.n11 VDD1.t6 8.28502
R1901 VDD1.n11 VDD1.t9 8.28502
R1902 VDD1.n26 VDD1.t0 8.28502
R1903 VDD1.n26 VDD1.t3 8.28502
R1904 VDD1.n24 VDD1.t4 8.28502
R1905 VDD1.n24 VDD1.t8 8.28502
R1906 VDD1.n3 VDD1.n1 4.69785
R1907 VDD1.n16 VDD1.n14 4.69785
R1908 VDD1.n10 VDD1.n0 1.93989
R1909 VDD1.n23 VDD1.n13 1.93989
R1910 VDD1 VDD1.n29 1.8561
R1911 VDD1.n8 VDD1.n7 1.16414
R1912 VDD1.n21 VDD1.n20 1.16414
R1913 VDD1 VDD1.n12 0.696621
R1914 VDD1.n27 VDD1.n25 0.583085
R1915 VDD1.n4 VDD1.n2 0.388379
R1916 VDD1.n17 VDD1.n15 0.388379
R1917 VDD1.n9 VDD1.n1 0.155672
R1918 VDD1.n22 VDD1.n14 0.155672
C0 VTAIL VDD2 6.04412f
C1 VN VDD1 0.159493f
C2 VP VDD2 0.593868f
C3 VP VTAIL 3.94513f
C4 VDD2 VDD1 2.19394f
C5 VTAIL VDD1 5.99074f
C6 VN VDD2 2.54322f
C7 VP VDD1 2.97393f
C8 VN VTAIL 3.93099f
C9 VN VP 6.66973f
C10 VDD2 B 5.653098f
C11 VDD1 B 5.544736f
C12 VTAIL B 3.910884f
C13 VN B 17.44759f
C14 VP B 15.883682f
C15 VDD1.n0 B 0.03778f
C16 VDD1.n1 B 0.213772f
C17 VDD1.n2 B 0.016062f
C18 VDD1.t2 B 0.064181f
C19 VDD1.n3 B 0.102045f
C20 VDD1.n4 B 0.021492f
C21 VDD1.n5 B 0.028474f
C22 VDD1.n6 B 0.0747f
C23 VDD1.n7 B 0.017007f
C24 VDD1.n8 B 0.016062f
C25 VDD1.n9 B 0.068685f
C26 VDD1.n10 B 0.076758f
C27 VDD1.t6 B 0.056455f
C28 VDD1.t9 B 0.056455f
C29 VDD1.n11 B 0.398755f
C30 VDD1.n12 B 0.815306f
C31 VDD1.n13 B 0.03778f
C32 VDD1.n14 B 0.213772f
C33 VDD1.n15 B 0.016062f
C34 VDD1.t5 B 0.064181f
C35 VDD1.n16 B 0.102045f
C36 VDD1.n17 B 0.021492f
C37 VDD1.n18 B 0.028474f
C38 VDD1.n19 B 0.0747f
C39 VDD1.n20 B 0.017007f
C40 VDD1.n21 B 0.016062f
C41 VDD1.n22 B 0.068685f
C42 VDD1.n23 B 0.076758f
C43 VDD1.t4 B 0.056455f
C44 VDD1.t8 B 0.056455f
C45 VDD1.n24 B 0.398754f
C46 VDD1.n25 B 0.805562f
C47 VDD1.t0 B 0.056455f
C48 VDD1.t3 B 0.056455f
C49 VDD1.n26 B 0.412735f
C50 VDD1.n27 B 2.91474f
C51 VDD1.t1 B 0.056455f
C52 VDD1.t7 B 0.056455f
C53 VDD1.n28 B 0.398754f
C54 VDD1.n29 B 2.88394f
C55 VP.n0 B 0.038809f
C56 VP.t6 B 0.446211f
C57 VP.n1 B 0.047893f
C58 VP.n2 B 0.029436f
C59 VP.t9 B 0.446211f
C60 VP.n3 B 0.199929f
C61 VP.n4 B 0.029436f
C62 VP.n5 B 0.041331f
C63 VP.n6 B 0.029436f
C64 VP.t1 B 0.446211f
C65 VP.n7 B 0.054862f
C66 VP.n8 B 0.029436f
C67 VP.n9 B 0.039152f
C68 VP.n10 B 0.029436f
C69 VP.n11 B 0.047893f
C70 VP.n12 B 0.038809f
C71 VP.t4 B 0.446211f
C72 VP.n13 B 0.038809f
C73 VP.t2 B 0.446211f
C74 VP.n14 B 0.047893f
C75 VP.n15 B 0.029436f
C76 VP.t8 B 0.446211f
C77 VP.n16 B 0.199929f
C78 VP.n17 B 0.029436f
C79 VP.n18 B 0.041331f
C80 VP.n19 B 0.029436f
C81 VP.t0 B 0.446211f
C82 VP.n20 B 0.054862f
C83 VP.n21 B 0.029436f
C84 VP.n22 B 0.039152f
C85 VP.t7 B 0.676774f
C86 VP.t3 B 0.446211f
C87 VP.n23 B 0.283181f
C88 VP.n24 B 0.276272f
C89 VP.n25 B 0.285407f
C90 VP.n26 B 0.029436f
C91 VP.n27 B 0.054862f
C92 VP.n28 B 0.044612f
C93 VP.n29 B 0.041331f
C94 VP.n30 B 0.029436f
C95 VP.n31 B 0.029436f
C96 VP.n32 B 0.029436f
C97 VP.n33 B 0.041319f
C98 VP.n34 B 0.199929f
C99 VP.n35 B 0.041319f
C100 VP.n36 B 0.054862f
C101 VP.n37 B 0.029436f
C102 VP.n38 B 0.029436f
C103 VP.n39 B 0.029436f
C104 VP.n40 B 0.044612f
C105 VP.n41 B 0.054862f
C106 VP.n42 B 0.039152f
C107 VP.n43 B 0.029436f
C108 VP.n44 B 0.029436f
C109 VP.n45 B 0.043486f
C110 VP.n46 B 0.054862f
C111 VP.n47 B 0.03805f
C112 VP.n48 B 0.029436f
C113 VP.n49 B 0.029436f
C114 VP.n50 B 0.029436f
C115 VP.n51 B 0.054862f
C116 VP.n52 B 0.036985f
C117 VP.n53 B 0.297133f
C118 VP.n54 B 1.44683f
C119 VP.n55 B 1.46984f
C120 VP.n56 B 0.297133f
C121 VP.n57 B 0.036985f
C122 VP.n58 B 0.054862f
C123 VP.n59 B 0.029436f
C124 VP.n60 B 0.029436f
C125 VP.n61 B 0.029436f
C126 VP.n62 B 0.03805f
C127 VP.n63 B 0.054862f
C128 VP.t5 B 0.446211f
C129 VP.n64 B 0.199929f
C130 VP.n65 B 0.043486f
C131 VP.n66 B 0.029436f
C132 VP.n67 B 0.029436f
C133 VP.n68 B 0.029436f
C134 VP.n69 B 0.054862f
C135 VP.n70 B 0.044612f
C136 VP.n71 B 0.041331f
C137 VP.n72 B 0.029436f
C138 VP.n73 B 0.029436f
C139 VP.n74 B 0.029436f
C140 VP.n75 B 0.041319f
C141 VP.n76 B 0.199929f
C142 VP.n77 B 0.041319f
C143 VP.n78 B 0.054862f
C144 VP.n79 B 0.029436f
C145 VP.n80 B 0.029436f
C146 VP.n81 B 0.029436f
C147 VP.n82 B 0.044612f
C148 VP.n83 B 0.054862f
C149 VP.n84 B 0.039152f
C150 VP.n85 B 0.029436f
C151 VP.n86 B 0.029436f
C152 VP.n87 B 0.043486f
C153 VP.n88 B 0.054862f
C154 VP.n89 B 0.03805f
C155 VP.n90 B 0.029436f
C156 VP.n91 B 0.029436f
C157 VP.n92 B 0.029436f
C158 VP.n93 B 0.054862f
C159 VP.n94 B 0.036985f
C160 VP.n95 B 0.297133f
C161 VP.n96 B 0.049418f
C162 VTAIL.t15 B 0.066189f
C163 VTAIL.t10 B 0.066189f
C164 VTAIL.n0 B 0.407544f
C165 VTAIL.n1 B 0.683617f
C166 VTAIL.n2 B 0.044294f
C167 VTAIL.n3 B 0.250632f
C168 VTAIL.n4 B 0.018832f
C169 VTAIL.t4 B 0.075248f
C170 VTAIL.n5 B 0.119641f
C171 VTAIL.n6 B 0.025197f
C172 VTAIL.n7 B 0.033384f
C173 VTAIL.n8 B 0.08758f
C174 VTAIL.n9 B 0.01994f
C175 VTAIL.n10 B 0.018832f
C176 VTAIL.n11 B 0.080528f
C177 VTAIL.n12 B 0.048087f
C178 VTAIL.n13 B 0.514948f
C179 VTAIL.t9 B 0.066189f
C180 VTAIL.t3 B 0.066189f
C181 VTAIL.n14 B 0.407544f
C182 VTAIL.n15 B 0.840107f
C183 VTAIL.t5 B 0.066189f
C184 VTAIL.t2 B 0.066189f
C185 VTAIL.n16 B 0.407544f
C186 VTAIL.n17 B 1.83698f
C187 VTAIL.t11 B 0.066189f
C188 VTAIL.t18 B 0.066189f
C189 VTAIL.n18 B 0.407547f
C190 VTAIL.n19 B 1.83698f
C191 VTAIL.t16 B 0.066189f
C192 VTAIL.t14 B 0.066189f
C193 VTAIL.n20 B 0.407547f
C194 VTAIL.n21 B 0.840104f
C195 VTAIL.n22 B 0.044294f
C196 VTAIL.n23 B 0.250632f
C197 VTAIL.n24 B 0.018832f
C198 VTAIL.t13 B 0.075248f
C199 VTAIL.n25 B 0.119641f
C200 VTAIL.n26 B 0.025197f
C201 VTAIL.n27 B 0.033384f
C202 VTAIL.n28 B 0.08758f
C203 VTAIL.n29 B 0.01994f
C204 VTAIL.n30 B 0.018832f
C205 VTAIL.n31 B 0.080528f
C206 VTAIL.n32 B 0.048087f
C207 VTAIL.n33 B 0.514948f
C208 VTAIL.t0 B 0.066189f
C209 VTAIL.t6 B 0.066189f
C210 VTAIL.n34 B 0.407547f
C211 VTAIL.n35 B 0.749082f
C212 VTAIL.t7 B 0.066189f
C213 VTAIL.t1 B 0.066189f
C214 VTAIL.n36 B 0.407547f
C215 VTAIL.n37 B 0.840104f
C216 VTAIL.n38 B 0.044294f
C217 VTAIL.n39 B 0.250632f
C218 VTAIL.n40 B 0.018832f
C219 VTAIL.t8 B 0.075248f
C220 VTAIL.n41 B 0.119641f
C221 VTAIL.n42 B 0.025197f
C222 VTAIL.n43 B 0.033384f
C223 VTAIL.n44 B 0.08758f
C224 VTAIL.n45 B 0.01994f
C225 VTAIL.n46 B 0.018832f
C226 VTAIL.n47 B 0.080528f
C227 VTAIL.n48 B 0.048087f
C228 VTAIL.n49 B 1.31469f
C229 VTAIL.n50 B 0.044294f
C230 VTAIL.n51 B 0.250632f
C231 VTAIL.n52 B 0.018832f
C232 VTAIL.t12 B 0.075248f
C233 VTAIL.n53 B 0.119641f
C234 VTAIL.n54 B 0.025197f
C235 VTAIL.n55 B 0.033384f
C236 VTAIL.n56 B 0.08758f
C237 VTAIL.n57 B 0.01994f
C238 VTAIL.n58 B 0.018832f
C239 VTAIL.n59 B 0.080528f
C240 VTAIL.n60 B 0.048087f
C241 VTAIL.n61 B 1.31469f
C242 VTAIL.t17 B 0.066189f
C243 VTAIL.t19 B 0.066189f
C244 VTAIL.n62 B 0.407544f
C245 VTAIL.n63 B 0.61742f
C246 VDD2.n0 B 0.036453f
C247 VDD2.n1 B 0.206262f
C248 VDD2.n2 B 0.015498f
C249 VDD2.t3 B 0.061926f
C250 VDD2.n3 B 0.09846f
C251 VDD2.n4 B 0.020737f
C252 VDD2.n5 B 0.027474f
C253 VDD2.n6 B 0.072076f
C254 VDD2.n7 B 0.01641f
C255 VDD2.n8 B 0.015498f
C256 VDD2.n9 B 0.066272f
C257 VDD2.n10 B 0.074061f
C258 VDD2.t6 B 0.054472f
C259 VDD2.t1 B 0.054472f
C260 VDD2.n11 B 0.384745f
C261 VDD2.n12 B 0.777261f
C262 VDD2.t5 B 0.054472f
C263 VDD2.t8 B 0.054472f
C264 VDD2.n13 B 0.398235f
C265 VDD2.n14 B 2.67726f
C266 VDD2.n15 B 0.036453f
C267 VDD2.n16 B 0.206262f
C268 VDD2.n17 B 0.015498f
C269 VDD2.t9 B 0.061926f
C270 VDD2.n18 B 0.09846f
C271 VDD2.n19 B 0.020737f
C272 VDD2.n20 B 0.027474f
C273 VDD2.n21 B 0.072076f
C274 VDD2.n22 B 0.01641f
C275 VDD2.n23 B 0.015498f
C276 VDD2.n24 B 0.066272f
C277 VDD2.n25 B 0.059492f
C278 VDD2.n26 B 2.47548f
C279 VDD2.t0 B 0.054472f
C280 VDD2.t2 B 0.054472f
C281 VDD2.n27 B 0.384747f
C282 VDD2.n28 B 0.50878f
C283 VDD2.t4 B 0.054472f
C284 VDD2.t7 B 0.054472f
C285 VDD2.n29 B 0.398201f
C286 VN.n0 B 0.037268f
C287 VN.t7 B 0.428503f
C288 VN.n1 B 0.045992f
C289 VN.n2 B 0.028268f
C290 VN.t0 B 0.428503f
C291 VN.n3 B 0.191995f
C292 VN.n4 B 0.028268f
C293 VN.n5 B 0.039691f
C294 VN.n6 B 0.028268f
C295 VN.t2 B 0.428503f
C296 VN.n7 B 0.052684f
C297 VN.n8 B 0.028268f
C298 VN.n9 B 0.037598f
C299 VN.t4 B 0.649916f
C300 VN.t9 B 0.428503f
C301 VN.n10 B 0.271943f
C302 VN.n11 B 0.265308f
C303 VN.n12 B 0.27408f
C304 VN.n13 B 0.028268f
C305 VN.n14 B 0.052684f
C306 VN.n15 B 0.042841f
C307 VN.n16 B 0.039691f
C308 VN.n17 B 0.028268f
C309 VN.n18 B 0.028268f
C310 VN.n19 B 0.028268f
C311 VN.n20 B 0.039679f
C312 VN.n21 B 0.191995f
C313 VN.n22 B 0.039679f
C314 VN.n23 B 0.052684f
C315 VN.n24 B 0.028268f
C316 VN.n25 B 0.028268f
C317 VN.n26 B 0.028268f
C318 VN.n27 B 0.042841f
C319 VN.n28 B 0.052684f
C320 VN.n29 B 0.037598f
C321 VN.n30 B 0.028268f
C322 VN.n31 B 0.028268f
C323 VN.n32 B 0.04176f
C324 VN.n33 B 0.052684f
C325 VN.n34 B 0.03654f
C326 VN.n35 B 0.028268f
C327 VN.n36 B 0.028268f
C328 VN.n37 B 0.028268f
C329 VN.n38 B 0.052684f
C330 VN.n39 B 0.035517f
C331 VN.n40 B 0.285341f
C332 VN.n41 B 0.047457f
C333 VN.n42 B 0.037268f
C334 VN.t8 B 0.428503f
C335 VN.n43 B 0.045992f
C336 VN.n44 B 0.028268f
C337 VN.t1 B 0.428503f
C338 VN.n45 B 0.191995f
C339 VN.n46 B 0.028268f
C340 VN.n47 B 0.039691f
C341 VN.n48 B 0.028268f
C342 VN.t3 B 0.428503f
C343 VN.n49 B 0.052684f
C344 VN.n50 B 0.028268f
C345 VN.n51 B 0.037598f
C346 VN.t6 B 0.649916f
C347 VN.t5 B 0.428503f
C348 VN.n52 B 0.271943f
C349 VN.n53 B 0.265308f
C350 VN.n54 B 0.27408f
C351 VN.n55 B 0.028268f
C352 VN.n56 B 0.052684f
C353 VN.n57 B 0.042841f
C354 VN.n58 B 0.039691f
C355 VN.n59 B 0.028268f
C356 VN.n60 B 0.028268f
C357 VN.n61 B 0.028268f
C358 VN.n62 B 0.039679f
C359 VN.n63 B 0.191995f
C360 VN.n64 B 0.039679f
C361 VN.n65 B 0.052684f
C362 VN.n66 B 0.028268f
C363 VN.n67 B 0.028268f
C364 VN.n68 B 0.028268f
C365 VN.n69 B 0.042841f
C366 VN.n70 B 0.052684f
C367 VN.n71 B 0.037598f
C368 VN.n72 B 0.028268f
C369 VN.n73 B 0.028268f
C370 VN.n74 B 0.04176f
C371 VN.n75 B 0.052684f
C372 VN.n76 B 0.03654f
C373 VN.n77 B 0.028268f
C374 VN.n78 B 0.028268f
C375 VN.n79 B 0.028268f
C376 VN.n80 B 0.052684f
C377 VN.n81 B 0.035517f
C378 VN.n82 B 0.285341f
C379 VN.n83 B 1.40481f
.ends

