* NGSPICE file created from diff_pair_sample_1381.ext - technology: sky130A

.subckt diff_pair_sample_1381 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X1 VTAIL.t8 VP.t1 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X2 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=1
X3 VTAIL.t15 VP.t2 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X4 VDD2.t9 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=1
X5 VTAIL.t14 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X6 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=1
X7 VTAIL.t10 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X8 VDD1.t4 VP.t5 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=1
X9 VDD1.t3 VP.t6 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=1
X10 VTAIL.t18 VN.t2 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X11 VDD2.t6 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=1
X12 VTAIL.t17 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X13 VDD1.t2 VP.t7 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X14 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=1
X15 VDD2.t4 VN.t5 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X16 VDD2.t3 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=1.7979 ps=10 w=4.61 l=1
X17 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=1
X18 VDD2.t2 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0 ps=0 w=4.61 l=1
X20 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X21 VDD1.t1 VP.t8 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=1
X22 VTAIL.t5 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76065 pd=4.94 as=0.76065 ps=4.94 w=4.61 l=1
X23 VDD1.t0 VP.t9 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7979 pd=10 as=0.76065 ps=4.94 w=4.61 l=1
R0 VP.n9 VP.t9 164.95
R1 VP.n10 VP.n7 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n13 VP.n6 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n5 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n21 VP.n4 161.3
R8 VP.n40 VP.n0 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n36 VP.n1 161.3
R11 VP.n35 VP.n34 161.3
R12 VP.n32 VP.n2 161.3
R13 VP.n31 VP.n30 161.3
R14 VP.n29 VP.n3 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n25 VP.t8 150.625
R17 VP.n41 VP.t5 150.625
R18 VP.n22 VP.t6 150.625
R19 VP.n26 VP.t3 111.102
R20 VP.n33 VP.t7 111.102
R21 VP.n39 VP.t4 111.102
R22 VP.n20 VP.t2 111.102
R23 VP.n14 VP.t0 111.102
R24 VP.n8 VP.t1 111.102
R25 VP.n23 VP.n22 80.6037
R26 VP.n42 VP.n41 80.6037
R27 VP.n25 VP.n24 80.6037
R28 VP.n27 VP.n25 52.1152
R29 VP.n41 VP.n40 52.1152
R30 VP.n22 VP.n21 52.1152
R31 VP.n9 VP.n8 49.1161
R32 VP.n32 VP.n31 48.7492
R33 VP.n34 VP.n1 48.7492
R34 VP.n15 VP.n5 48.7492
R35 VP.n13 VP.n12 48.7492
R36 VP.n10 VP.n9 44.523
R37 VP.n24 VP.n23 38.9673
R38 VP.n31 VP.n3 32.2376
R39 VP.n38 VP.n1 32.2376
R40 VP.n19 VP.n5 32.2376
R41 VP.n12 VP.n7 32.2376
R42 VP.n27 VP.n26 20.5528
R43 VP.n40 VP.n39 20.5528
R44 VP.n21 VP.n20 20.5528
R45 VP.n33 VP.n32 12.234
R46 VP.n34 VP.n33 12.234
R47 VP.n14 VP.n13 12.234
R48 VP.n15 VP.n14 12.234
R49 VP.n26 VP.n3 3.91522
R50 VP.n39 VP.n38 3.91522
R51 VP.n20 VP.n19 3.91522
R52 VP.n8 VP.n7 3.91522
R53 VP.n23 VP.n4 0.285035
R54 VP.n28 VP.n24 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n11 VP.n10 0.189894
R57 VP.n11 VP.n6 0.189894
R58 VP.n16 VP.n6 0.189894
R59 VP.n17 VP.n16 0.189894
R60 VP.n18 VP.n17 0.189894
R61 VP.n18 VP.n4 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n30 VP.n29 0.189894
R64 VP.n30 VP.n2 0.189894
R65 VP.n35 VP.n2 0.189894
R66 VP.n36 VP.n35 0.189894
R67 VP.n37 VP.n36 0.189894
R68 VP.n37 VP.n0 0.189894
R69 VP VP.n42 0.146778
R70 VTAIL.n104 VTAIL.n86 289.615
R71 VTAIL.n20 VTAIL.n2 289.615
R72 VTAIL.n80 VTAIL.n62 289.615
R73 VTAIL.n52 VTAIL.n34 289.615
R74 VTAIL.n95 VTAIL.n94 185
R75 VTAIL.n97 VTAIL.n96 185
R76 VTAIL.n90 VTAIL.n89 185
R77 VTAIL.n103 VTAIL.n102 185
R78 VTAIL.n105 VTAIL.n104 185
R79 VTAIL.n11 VTAIL.n10 185
R80 VTAIL.n13 VTAIL.n12 185
R81 VTAIL.n6 VTAIL.n5 185
R82 VTAIL.n19 VTAIL.n18 185
R83 VTAIL.n21 VTAIL.n20 185
R84 VTAIL.n81 VTAIL.n80 185
R85 VTAIL.n79 VTAIL.n78 185
R86 VTAIL.n66 VTAIL.n65 185
R87 VTAIL.n73 VTAIL.n72 185
R88 VTAIL.n71 VTAIL.n70 185
R89 VTAIL.n53 VTAIL.n52 185
R90 VTAIL.n51 VTAIL.n50 185
R91 VTAIL.n38 VTAIL.n37 185
R92 VTAIL.n45 VTAIL.n44 185
R93 VTAIL.n43 VTAIL.n42 185
R94 VTAIL.n93 VTAIL.t3 147.714
R95 VTAIL.n9 VTAIL.t16 147.714
R96 VTAIL.n69 VTAIL.t7 147.714
R97 VTAIL.n41 VTAIL.t1 147.714
R98 VTAIL.n96 VTAIL.n95 104.615
R99 VTAIL.n96 VTAIL.n89 104.615
R100 VTAIL.n103 VTAIL.n89 104.615
R101 VTAIL.n104 VTAIL.n103 104.615
R102 VTAIL.n12 VTAIL.n11 104.615
R103 VTAIL.n12 VTAIL.n5 104.615
R104 VTAIL.n19 VTAIL.n5 104.615
R105 VTAIL.n20 VTAIL.n19 104.615
R106 VTAIL.n80 VTAIL.n79 104.615
R107 VTAIL.n79 VTAIL.n65 104.615
R108 VTAIL.n72 VTAIL.n65 104.615
R109 VTAIL.n72 VTAIL.n71 104.615
R110 VTAIL.n52 VTAIL.n51 104.615
R111 VTAIL.n51 VTAIL.n37 104.615
R112 VTAIL.n44 VTAIL.n37 104.615
R113 VTAIL.n44 VTAIL.n43 104.615
R114 VTAIL.n61 VTAIL.n60 54.9327
R115 VTAIL.n59 VTAIL.n58 54.9327
R116 VTAIL.n33 VTAIL.n32 54.9327
R117 VTAIL.n31 VTAIL.n30 54.9327
R118 VTAIL.n111 VTAIL.n110 54.9326
R119 VTAIL.n1 VTAIL.n0 54.9326
R120 VTAIL.n27 VTAIL.n26 54.9326
R121 VTAIL.n29 VTAIL.n28 54.9326
R122 VTAIL.n95 VTAIL.t3 52.3082
R123 VTAIL.n11 VTAIL.t16 52.3082
R124 VTAIL.n71 VTAIL.t7 52.3082
R125 VTAIL.n43 VTAIL.t1 52.3082
R126 VTAIL.n109 VTAIL.n108 33.155
R127 VTAIL.n25 VTAIL.n24 33.155
R128 VTAIL.n85 VTAIL.n84 33.155
R129 VTAIL.n57 VTAIL.n56 33.155
R130 VTAIL.n31 VTAIL.n29 18.6341
R131 VTAIL.n109 VTAIL.n85 17.4876
R132 VTAIL.n94 VTAIL.n93 15.6631
R133 VTAIL.n10 VTAIL.n9 15.6631
R134 VTAIL.n70 VTAIL.n69 15.6631
R135 VTAIL.n42 VTAIL.n41 15.6631
R136 VTAIL.n97 VTAIL.n92 12.8005
R137 VTAIL.n13 VTAIL.n8 12.8005
R138 VTAIL.n73 VTAIL.n68 12.8005
R139 VTAIL.n45 VTAIL.n40 12.8005
R140 VTAIL.n98 VTAIL.n90 12.0247
R141 VTAIL.n14 VTAIL.n6 12.0247
R142 VTAIL.n74 VTAIL.n66 12.0247
R143 VTAIL.n46 VTAIL.n38 12.0247
R144 VTAIL.n102 VTAIL.n101 11.249
R145 VTAIL.n18 VTAIL.n17 11.249
R146 VTAIL.n78 VTAIL.n77 11.249
R147 VTAIL.n50 VTAIL.n49 11.249
R148 VTAIL.n105 VTAIL.n88 10.4732
R149 VTAIL.n21 VTAIL.n4 10.4732
R150 VTAIL.n81 VTAIL.n64 10.4732
R151 VTAIL.n53 VTAIL.n36 10.4732
R152 VTAIL.n106 VTAIL.n86 9.69747
R153 VTAIL.n22 VTAIL.n2 9.69747
R154 VTAIL.n82 VTAIL.n62 9.69747
R155 VTAIL.n54 VTAIL.n34 9.69747
R156 VTAIL.n108 VTAIL.n107 9.45567
R157 VTAIL.n24 VTAIL.n23 9.45567
R158 VTAIL.n84 VTAIL.n83 9.45567
R159 VTAIL.n56 VTAIL.n55 9.45567
R160 VTAIL.n107 VTAIL.n106 9.3005
R161 VTAIL.n88 VTAIL.n87 9.3005
R162 VTAIL.n101 VTAIL.n100 9.3005
R163 VTAIL.n99 VTAIL.n98 9.3005
R164 VTAIL.n92 VTAIL.n91 9.3005
R165 VTAIL.n23 VTAIL.n22 9.3005
R166 VTAIL.n4 VTAIL.n3 9.3005
R167 VTAIL.n17 VTAIL.n16 9.3005
R168 VTAIL.n15 VTAIL.n14 9.3005
R169 VTAIL.n8 VTAIL.n7 9.3005
R170 VTAIL.n83 VTAIL.n82 9.3005
R171 VTAIL.n64 VTAIL.n63 9.3005
R172 VTAIL.n77 VTAIL.n76 9.3005
R173 VTAIL.n75 VTAIL.n74 9.3005
R174 VTAIL.n68 VTAIL.n67 9.3005
R175 VTAIL.n55 VTAIL.n54 9.3005
R176 VTAIL.n36 VTAIL.n35 9.3005
R177 VTAIL.n49 VTAIL.n48 9.3005
R178 VTAIL.n47 VTAIL.n46 9.3005
R179 VTAIL.n40 VTAIL.n39 9.3005
R180 VTAIL.n93 VTAIL.n91 4.39059
R181 VTAIL.n9 VTAIL.n7 4.39059
R182 VTAIL.n69 VTAIL.n67 4.39059
R183 VTAIL.n41 VTAIL.n39 4.39059
R184 VTAIL.n110 VTAIL.t19 4.29551
R185 VTAIL.n110 VTAIL.t17 4.29551
R186 VTAIL.n0 VTAIL.t2 4.29551
R187 VTAIL.n0 VTAIL.t18 4.29551
R188 VTAIL.n26 VTAIL.t13 4.29551
R189 VTAIL.n26 VTAIL.t10 4.29551
R190 VTAIL.n28 VTAIL.t11 4.29551
R191 VTAIL.n28 VTAIL.t14 4.29551
R192 VTAIL.n60 VTAIL.t12 4.29551
R193 VTAIL.n60 VTAIL.t15 4.29551
R194 VTAIL.n58 VTAIL.t9 4.29551
R195 VTAIL.n58 VTAIL.t8 4.29551
R196 VTAIL.n32 VTAIL.t4 4.29551
R197 VTAIL.n32 VTAIL.t0 4.29551
R198 VTAIL.n30 VTAIL.t6 4.29551
R199 VTAIL.n30 VTAIL.t5 4.29551
R200 VTAIL.n108 VTAIL.n86 4.26717
R201 VTAIL.n24 VTAIL.n2 4.26717
R202 VTAIL.n84 VTAIL.n62 4.26717
R203 VTAIL.n56 VTAIL.n34 4.26717
R204 VTAIL.n106 VTAIL.n105 3.49141
R205 VTAIL.n22 VTAIL.n21 3.49141
R206 VTAIL.n82 VTAIL.n81 3.49141
R207 VTAIL.n54 VTAIL.n53 3.49141
R208 VTAIL.n102 VTAIL.n88 2.71565
R209 VTAIL.n18 VTAIL.n4 2.71565
R210 VTAIL.n78 VTAIL.n64 2.71565
R211 VTAIL.n50 VTAIL.n36 2.71565
R212 VTAIL.n101 VTAIL.n90 1.93989
R213 VTAIL.n17 VTAIL.n6 1.93989
R214 VTAIL.n77 VTAIL.n66 1.93989
R215 VTAIL.n49 VTAIL.n38 1.93989
R216 VTAIL.n98 VTAIL.n97 1.16414
R217 VTAIL.n14 VTAIL.n13 1.16414
R218 VTAIL.n74 VTAIL.n73 1.16414
R219 VTAIL.n46 VTAIL.n45 1.16414
R220 VTAIL.n33 VTAIL.n31 1.14705
R221 VTAIL.n57 VTAIL.n33 1.14705
R222 VTAIL.n61 VTAIL.n59 1.14705
R223 VTAIL.n85 VTAIL.n61 1.14705
R224 VTAIL.n29 VTAIL.n27 1.14705
R225 VTAIL.n27 VTAIL.n25 1.14705
R226 VTAIL.n111 VTAIL.n109 1.14705
R227 VTAIL.n59 VTAIL.n57 1.0436
R228 VTAIL.n25 VTAIL.n1 1.0436
R229 VTAIL VTAIL.n1 0.918603
R230 VTAIL.n94 VTAIL.n92 0.388379
R231 VTAIL.n10 VTAIL.n8 0.388379
R232 VTAIL.n70 VTAIL.n68 0.388379
R233 VTAIL.n42 VTAIL.n40 0.388379
R234 VTAIL VTAIL.n111 0.228948
R235 VTAIL.n99 VTAIL.n91 0.155672
R236 VTAIL.n100 VTAIL.n99 0.155672
R237 VTAIL.n100 VTAIL.n87 0.155672
R238 VTAIL.n107 VTAIL.n87 0.155672
R239 VTAIL.n15 VTAIL.n7 0.155672
R240 VTAIL.n16 VTAIL.n15 0.155672
R241 VTAIL.n16 VTAIL.n3 0.155672
R242 VTAIL.n23 VTAIL.n3 0.155672
R243 VTAIL.n83 VTAIL.n63 0.155672
R244 VTAIL.n76 VTAIL.n63 0.155672
R245 VTAIL.n76 VTAIL.n75 0.155672
R246 VTAIL.n75 VTAIL.n67 0.155672
R247 VTAIL.n55 VTAIL.n35 0.155672
R248 VTAIL.n48 VTAIL.n35 0.155672
R249 VTAIL.n48 VTAIL.n47 0.155672
R250 VTAIL.n47 VTAIL.n39 0.155672
R251 VDD1.n18 VDD1.n0 289.615
R252 VDD1.n43 VDD1.n25 289.615
R253 VDD1.n19 VDD1.n18 185
R254 VDD1.n17 VDD1.n16 185
R255 VDD1.n4 VDD1.n3 185
R256 VDD1.n11 VDD1.n10 185
R257 VDD1.n9 VDD1.n8 185
R258 VDD1.n34 VDD1.n33 185
R259 VDD1.n36 VDD1.n35 185
R260 VDD1.n29 VDD1.n28 185
R261 VDD1.n42 VDD1.n41 185
R262 VDD1.n44 VDD1.n43 185
R263 VDD1.n7 VDD1.t0 147.714
R264 VDD1.n32 VDD1.t1 147.714
R265 VDD1.n18 VDD1.n17 104.615
R266 VDD1.n17 VDD1.n3 104.615
R267 VDD1.n10 VDD1.n3 104.615
R268 VDD1.n10 VDD1.n9 104.615
R269 VDD1.n35 VDD1.n34 104.615
R270 VDD1.n35 VDD1.n28 104.615
R271 VDD1.n42 VDD1.n28 104.615
R272 VDD1.n43 VDD1.n42 104.615
R273 VDD1.n51 VDD1.n50 72.4159
R274 VDD1.n24 VDD1.n23 71.6115
R275 VDD1.n53 VDD1.n52 71.6113
R276 VDD1.n49 VDD1.n48 71.6113
R277 VDD1.n9 VDD1.t0 52.3082
R278 VDD1.n34 VDD1.t1 52.3082
R279 VDD1.n24 VDD1.n22 50.9804
R280 VDD1.n49 VDD1.n47 50.9804
R281 VDD1.n53 VDD1.n51 34.2918
R282 VDD1.n8 VDD1.n7 15.6631
R283 VDD1.n33 VDD1.n32 15.6631
R284 VDD1.n11 VDD1.n6 12.8005
R285 VDD1.n36 VDD1.n31 12.8005
R286 VDD1.n12 VDD1.n4 12.0247
R287 VDD1.n37 VDD1.n29 12.0247
R288 VDD1.n16 VDD1.n15 11.249
R289 VDD1.n41 VDD1.n40 11.249
R290 VDD1.n19 VDD1.n2 10.4732
R291 VDD1.n44 VDD1.n27 10.4732
R292 VDD1.n20 VDD1.n0 9.69747
R293 VDD1.n45 VDD1.n25 9.69747
R294 VDD1.n22 VDD1.n21 9.45567
R295 VDD1.n47 VDD1.n46 9.45567
R296 VDD1.n21 VDD1.n20 9.3005
R297 VDD1.n2 VDD1.n1 9.3005
R298 VDD1.n15 VDD1.n14 9.3005
R299 VDD1.n13 VDD1.n12 9.3005
R300 VDD1.n6 VDD1.n5 9.3005
R301 VDD1.n46 VDD1.n45 9.3005
R302 VDD1.n27 VDD1.n26 9.3005
R303 VDD1.n40 VDD1.n39 9.3005
R304 VDD1.n38 VDD1.n37 9.3005
R305 VDD1.n31 VDD1.n30 9.3005
R306 VDD1.n7 VDD1.n5 4.39059
R307 VDD1.n32 VDD1.n30 4.39059
R308 VDD1.n52 VDD1.t7 4.29551
R309 VDD1.n52 VDD1.t3 4.29551
R310 VDD1.n23 VDD1.t8 4.29551
R311 VDD1.n23 VDD1.t9 4.29551
R312 VDD1.n50 VDD1.t5 4.29551
R313 VDD1.n50 VDD1.t4 4.29551
R314 VDD1.n48 VDD1.t6 4.29551
R315 VDD1.n48 VDD1.t2 4.29551
R316 VDD1.n22 VDD1.n0 4.26717
R317 VDD1.n47 VDD1.n25 4.26717
R318 VDD1.n20 VDD1.n19 3.49141
R319 VDD1.n45 VDD1.n44 3.49141
R320 VDD1.n16 VDD1.n2 2.71565
R321 VDD1.n41 VDD1.n27 2.71565
R322 VDD1.n15 VDD1.n4 1.93989
R323 VDD1.n40 VDD1.n29 1.93989
R324 VDD1.n12 VDD1.n11 1.16414
R325 VDD1.n37 VDD1.n36 1.16414
R326 VDD1 VDD1.n53 0.802224
R327 VDD1.n8 VDD1.n6 0.388379
R328 VDD1.n33 VDD1.n31 0.388379
R329 VDD1 VDD1.n24 0.345328
R330 VDD1.n51 VDD1.n49 0.231792
R331 VDD1.n21 VDD1.n1 0.155672
R332 VDD1.n14 VDD1.n1 0.155672
R333 VDD1.n14 VDD1.n13 0.155672
R334 VDD1.n13 VDD1.n5 0.155672
R335 VDD1.n38 VDD1.n30 0.155672
R336 VDD1.n39 VDD1.n38 0.155672
R337 VDD1.n39 VDD1.n26 0.155672
R338 VDD1.n46 VDD1.n26 0.155672
R339 B.n507 B.n506 585
R340 B.n508 B.n507 585
R341 B.n182 B.n84 585
R342 B.n181 B.n180 585
R343 B.n179 B.n178 585
R344 B.n177 B.n176 585
R345 B.n175 B.n174 585
R346 B.n173 B.n172 585
R347 B.n171 B.n170 585
R348 B.n169 B.n168 585
R349 B.n167 B.n166 585
R350 B.n165 B.n164 585
R351 B.n163 B.n162 585
R352 B.n161 B.n160 585
R353 B.n159 B.n158 585
R354 B.n157 B.n156 585
R355 B.n155 B.n154 585
R356 B.n153 B.n152 585
R357 B.n151 B.n150 585
R358 B.n149 B.n148 585
R359 B.n147 B.n146 585
R360 B.n144 B.n143 585
R361 B.n142 B.n141 585
R362 B.n140 B.n139 585
R363 B.n138 B.n137 585
R364 B.n136 B.n135 585
R365 B.n134 B.n133 585
R366 B.n132 B.n131 585
R367 B.n130 B.n129 585
R368 B.n128 B.n127 585
R369 B.n126 B.n125 585
R370 B.n124 B.n123 585
R371 B.n122 B.n121 585
R372 B.n120 B.n119 585
R373 B.n118 B.n117 585
R374 B.n116 B.n115 585
R375 B.n114 B.n113 585
R376 B.n112 B.n111 585
R377 B.n110 B.n109 585
R378 B.n108 B.n107 585
R379 B.n106 B.n105 585
R380 B.n104 B.n103 585
R381 B.n102 B.n101 585
R382 B.n100 B.n99 585
R383 B.n98 B.n97 585
R384 B.n96 B.n95 585
R385 B.n94 B.n93 585
R386 B.n92 B.n91 585
R387 B.n60 B.n59 585
R388 B.n511 B.n510 585
R389 B.n505 B.n85 585
R390 B.n85 B.n57 585
R391 B.n504 B.n56 585
R392 B.n515 B.n56 585
R393 B.n503 B.n55 585
R394 B.n516 B.n55 585
R395 B.n502 B.n54 585
R396 B.n517 B.n54 585
R397 B.n501 B.n500 585
R398 B.n500 B.n50 585
R399 B.n499 B.n49 585
R400 B.n523 B.n49 585
R401 B.n498 B.n48 585
R402 B.n524 B.n48 585
R403 B.n497 B.n47 585
R404 B.n525 B.n47 585
R405 B.n496 B.n495 585
R406 B.n495 B.n43 585
R407 B.n494 B.n42 585
R408 B.n531 B.n42 585
R409 B.n493 B.n41 585
R410 B.n532 B.n41 585
R411 B.n492 B.n40 585
R412 B.n533 B.n40 585
R413 B.n491 B.n490 585
R414 B.n490 B.n39 585
R415 B.n489 B.n35 585
R416 B.n539 B.n35 585
R417 B.n488 B.n34 585
R418 B.n540 B.n34 585
R419 B.n487 B.n33 585
R420 B.n541 B.n33 585
R421 B.n486 B.n485 585
R422 B.n485 B.n32 585
R423 B.n484 B.n28 585
R424 B.n547 B.n28 585
R425 B.n483 B.n27 585
R426 B.n548 B.n27 585
R427 B.n482 B.n26 585
R428 B.n549 B.n26 585
R429 B.n481 B.n480 585
R430 B.n480 B.n25 585
R431 B.n479 B.n21 585
R432 B.n555 B.n21 585
R433 B.n478 B.n20 585
R434 B.n556 B.n20 585
R435 B.n477 B.n19 585
R436 B.n557 B.n19 585
R437 B.n476 B.n475 585
R438 B.n475 B.n18 585
R439 B.n474 B.n14 585
R440 B.n563 B.n14 585
R441 B.n473 B.n13 585
R442 B.n564 B.n13 585
R443 B.n472 B.n12 585
R444 B.n565 B.n12 585
R445 B.n471 B.n470 585
R446 B.n470 B.n469 585
R447 B.n468 B.n467 585
R448 B.n468 B.n8 585
R449 B.n466 B.n7 585
R450 B.n572 B.n7 585
R451 B.n465 B.n6 585
R452 B.n573 B.n6 585
R453 B.n464 B.n5 585
R454 B.n574 B.n5 585
R455 B.n463 B.n462 585
R456 B.n462 B.n4 585
R457 B.n461 B.n183 585
R458 B.n461 B.n460 585
R459 B.n451 B.n184 585
R460 B.n185 B.n184 585
R461 B.n453 B.n452 585
R462 B.n454 B.n453 585
R463 B.n450 B.n190 585
R464 B.n190 B.n189 585
R465 B.n449 B.n448 585
R466 B.n448 B.n447 585
R467 B.n192 B.n191 585
R468 B.n440 B.n192 585
R469 B.n439 B.n438 585
R470 B.n441 B.n439 585
R471 B.n437 B.n197 585
R472 B.n197 B.n196 585
R473 B.n436 B.n435 585
R474 B.n435 B.n434 585
R475 B.n199 B.n198 585
R476 B.n427 B.n199 585
R477 B.n426 B.n425 585
R478 B.n428 B.n426 585
R479 B.n424 B.n204 585
R480 B.n204 B.n203 585
R481 B.n423 B.n422 585
R482 B.n422 B.n421 585
R483 B.n206 B.n205 585
R484 B.n414 B.n206 585
R485 B.n413 B.n412 585
R486 B.n415 B.n413 585
R487 B.n411 B.n211 585
R488 B.n211 B.n210 585
R489 B.n410 B.n409 585
R490 B.n409 B.n408 585
R491 B.n213 B.n212 585
R492 B.n401 B.n213 585
R493 B.n400 B.n399 585
R494 B.n402 B.n400 585
R495 B.n398 B.n218 585
R496 B.n218 B.n217 585
R497 B.n397 B.n396 585
R498 B.n396 B.n395 585
R499 B.n220 B.n219 585
R500 B.n221 B.n220 585
R501 B.n388 B.n387 585
R502 B.n389 B.n388 585
R503 B.n386 B.n226 585
R504 B.n226 B.n225 585
R505 B.n385 B.n384 585
R506 B.n384 B.n383 585
R507 B.n228 B.n227 585
R508 B.n229 B.n228 585
R509 B.n376 B.n375 585
R510 B.n377 B.n376 585
R511 B.n374 B.n234 585
R512 B.n234 B.n233 585
R513 B.n373 B.n372 585
R514 B.n372 B.n371 585
R515 B.n236 B.n235 585
R516 B.n237 B.n236 585
R517 B.n367 B.n366 585
R518 B.n240 B.n239 585
R519 B.n363 B.n362 585
R520 B.n364 B.n363 585
R521 B.n361 B.n264 585
R522 B.n360 B.n359 585
R523 B.n358 B.n357 585
R524 B.n356 B.n355 585
R525 B.n354 B.n353 585
R526 B.n352 B.n351 585
R527 B.n350 B.n349 585
R528 B.n348 B.n347 585
R529 B.n346 B.n345 585
R530 B.n344 B.n343 585
R531 B.n342 B.n341 585
R532 B.n340 B.n339 585
R533 B.n338 B.n337 585
R534 B.n336 B.n335 585
R535 B.n334 B.n333 585
R536 B.n332 B.n331 585
R537 B.n330 B.n329 585
R538 B.n327 B.n326 585
R539 B.n325 B.n324 585
R540 B.n323 B.n322 585
R541 B.n321 B.n320 585
R542 B.n319 B.n318 585
R543 B.n317 B.n316 585
R544 B.n315 B.n314 585
R545 B.n313 B.n312 585
R546 B.n311 B.n310 585
R547 B.n309 B.n308 585
R548 B.n307 B.n306 585
R549 B.n305 B.n304 585
R550 B.n303 B.n302 585
R551 B.n301 B.n300 585
R552 B.n299 B.n298 585
R553 B.n297 B.n296 585
R554 B.n295 B.n294 585
R555 B.n293 B.n292 585
R556 B.n291 B.n290 585
R557 B.n289 B.n288 585
R558 B.n287 B.n286 585
R559 B.n285 B.n284 585
R560 B.n283 B.n282 585
R561 B.n281 B.n280 585
R562 B.n279 B.n278 585
R563 B.n277 B.n276 585
R564 B.n275 B.n274 585
R565 B.n273 B.n272 585
R566 B.n271 B.n270 585
R567 B.n368 B.n238 585
R568 B.n238 B.n237 585
R569 B.n370 B.n369 585
R570 B.n371 B.n370 585
R571 B.n232 B.n231 585
R572 B.n233 B.n232 585
R573 B.n379 B.n378 585
R574 B.n378 B.n377 585
R575 B.n380 B.n230 585
R576 B.n230 B.n229 585
R577 B.n382 B.n381 585
R578 B.n383 B.n382 585
R579 B.n224 B.n223 585
R580 B.n225 B.n224 585
R581 B.n391 B.n390 585
R582 B.n390 B.n389 585
R583 B.n392 B.n222 585
R584 B.n222 B.n221 585
R585 B.n394 B.n393 585
R586 B.n395 B.n394 585
R587 B.n216 B.n215 585
R588 B.n217 B.n216 585
R589 B.n404 B.n403 585
R590 B.n403 B.n402 585
R591 B.n405 B.n214 585
R592 B.n401 B.n214 585
R593 B.n407 B.n406 585
R594 B.n408 B.n407 585
R595 B.n209 B.n208 585
R596 B.n210 B.n209 585
R597 B.n417 B.n416 585
R598 B.n416 B.n415 585
R599 B.n418 B.n207 585
R600 B.n414 B.n207 585
R601 B.n420 B.n419 585
R602 B.n421 B.n420 585
R603 B.n202 B.n201 585
R604 B.n203 B.n202 585
R605 B.n430 B.n429 585
R606 B.n429 B.n428 585
R607 B.n431 B.n200 585
R608 B.n427 B.n200 585
R609 B.n433 B.n432 585
R610 B.n434 B.n433 585
R611 B.n195 B.n194 585
R612 B.n196 B.n195 585
R613 B.n443 B.n442 585
R614 B.n442 B.n441 585
R615 B.n444 B.n193 585
R616 B.n440 B.n193 585
R617 B.n446 B.n445 585
R618 B.n447 B.n446 585
R619 B.n188 B.n187 585
R620 B.n189 B.n188 585
R621 B.n456 B.n455 585
R622 B.n455 B.n454 585
R623 B.n457 B.n186 585
R624 B.n186 B.n185 585
R625 B.n459 B.n458 585
R626 B.n460 B.n459 585
R627 B.n3 B.n0 585
R628 B.n4 B.n3 585
R629 B.n571 B.n1 585
R630 B.n572 B.n571 585
R631 B.n570 B.n569 585
R632 B.n570 B.n8 585
R633 B.n568 B.n9 585
R634 B.n469 B.n9 585
R635 B.n567 B.n566 585
R636 B.n566 B.n565 585
R637 B.n11 B.n10 585
R638 B.n564 B.n11 585
R639 B.n562 B.n561 585
R640 B.n563 B.n562 585
R641 B.n560 B.n15 585
R642 B.n18 B.n15 585
R643 B.n559 B.n558 585
R644 B.n558 B.n557 585
R645 B.n17 B.n16 585
R646 B.n556 B.n17 585
R647 B.n554 B.n553 585
R648 B.n555 B.n554 585
R649 B.n552 B.n22 585
R650 B.n25 B.n22 585
R651 B.n551 B.n550 585
R652 B.n550 B.n549 585
R653 B.n24 B.n23 585
R654 B.n548 B.n24 585
R655 B.n546 B.n545 585
R656 B.n547 B.n546 585
R657 B.n544 B.n29 585
R658 B.n32 B.n29 585
R659 B.n543 B.n542 585
R660 B.n542 B.n541 585
R661 B.n31 B.n30 585
R662 B.n540 B.n31 585
R663 B.n538 B.n537 585
R664 B.n539 B.n538 585
R665 B.n536 B.n36 585
R666 B.n39 B.n36 585
R667 B.n535 B.n534 585
R668 B.n534 B.n533 585
R669 B.n38 B.n37 585
R670 B.n532 B.n38 585
R671 B.n530 B.n529 585
R672 B.n531 B.n530 585
R673 B.n528 B.n44 585
R674 B.n44 B.n43 585
R675 B.n527 B.n526 585
R676 B.n526 B.n525 585
R677 B.n46 B.n45 585
R678 B.n524 B.n46 585
R679 B.n522 B.n521 585
R680 B.n523 B.n522 585
R681 B.n520 B.n51 585
R682 B.n51 B.n50 585
R683 B.n519 B.n518 585
R684 B.n518 B.n517 585
R685 B.n53 B.n52 585
R686 B.n516 B.n53 585
R687 B.n514 B.n513 585
R688 B.n515 B.n514 585
R689 B.n512 B.n58 585
R690 B.n58 B.n57 585
R691 B.n575 B.n574 585
R692 B.n573 B.n2 585
R693 B.n510 B.n58 540.549
R694 B.n507 B.n85 540.549
R695 B.n270 B.n236 540.549
R696 B.n366 B.n238 540.549
R697 B.n88 B.t10 314.026
R698 B.n86 B.t14 314.026
R699 B.n267 B.t21 314.026
R700 B.n265 B.t17 314.026
R701 B.n508 B.n83 256.663
R702 B.n508 B.n82 256.663
R703 B.n508 B.n81 256.663
R704 B.n508 B.n80 256.663
R705 B.n508 B.n79 256.663
R706 B.n508 B.n78 256.663
R707 B.n508 B.n77 256.663
R708 B.n508 B.n76 256.663
R709 B.n508 B.n75 256.663
R710 B.n508 B.n74 256.663
R711 B.n508 B.n73 256.663
R712 B.n508 B.n72 256.663
R713 B.n508 B.n71 256.663
R714 B.n508 B.n70 256.663
R715 B.n508 B.n69 256.663
R716 B.n508 B.n68 256.663
R717 B.n508 B.n67 256.663
R718 B.n508 B.n66 256.663
R719 B.n508 B.n65 256.663
R720 B.n508 B.n64 256.663
R721 B.n508 B.n63 256.663
R722 B.n508 B.n62 256.663
R723 B.n508 B.n61 256.663
R724 B.n509 B.n508 256.663
R725 B.n365 B.n364 256.663
R726 B.n364 B.n241 256.663
R727 B.n364 B.n242 256.663
R728 B.n364 B.n243 256.663
R729 B.n364 B.n244 256.663
R730 B.n364 B.n245 256.663
R731 B.n364 B.n246 256.663
R732 B.n364 B.n247 256.663
R733 B.n364 B.n248 256.663
R734 B.n364 B.n249 256.663
R735 B.n364 B.n250 256.663
R736 B.n364 B.n251 256.663
R737 B.n364 B.n252 256.663
R738 B.n364 B.n253 256.663
R739 B.n364 B.n254 256.663
R740 B.n364 B.n255 256.663
R741 B.n364 B.n256 256.663
R742 B.n364 B.n257 256.663
R743 B.n364 B.n258 256.663
R744 B.n364 B.n259 256.663
R745 B.n364 B.n260 256.663
R746 B.n364 B.n261 256.663
R747 B.n364 B.n262 256.663
R748 B.n364 B.n263 256.663
R749 B.n577 B.n576 256.663
R750 B.n86 B.t15 181.018
R751 B.n267 B.t23 181.018
R752 B.n88 B.t12 181.018
R753 B.n265 B.t20 181.018
R754 B.n91 B.n60 163.367
R755 B.n95 B.n94 163.367
R756 B.n99 B.n98 163.367
R757 B.n103 B.n102 163.367
R758 B.n107 B.n106 163.367
R759 B.n111 B.n110 163.367
R760 B.n115 B.n114 163.367
R761 B.n119 B.n118 163.367
R762 B.n123 B.n122 163.367
R763 B.n127 B.n126 163.367
R764 B.n131 B.n130 163.367
R765 B.n135 B.n134 163.367
R766 B.n139 B.n138 163.367
R767 B.n143 B.n142 163.367
R768 B.n148 B.n147 163.367
R769 B.n152 B.n151 163.367
R770 B.n156 B.n155 163.367
R771 B.n160 B.n159 163.367
R772 B.n164 B.n163 163.367
R773 B.n168 B.n167 163.367
R774 B.n172 B.n171 163.367
R775 B.n176 B.n175 163.367
R776 B.n180 B.n179 163.367
R777 B.n507 B.n84 163.367
R778 B.n372 B.n236 163.367
R779 B.n372 B.n234 163.367
R780 B.n376 B.n234 163.367
R781 B.n376 B.n228 163.367
R782 B.n384 B.n228 163.367
R783 B.n384 B.n226 163.367
R784 B.n388 B.n226 163.367
R785 B.n388 B.n220 163.367
R786 B.n396 B.n220 163.367
R787 B.n396 B.n218 163.367
R788 B.n400 B.n218 163.367
R789 B.n400 B.n213 163.367
R790 B.n409 B.n213 163.367
R791 B.n409 B.n211 163.367
R792 B.n413 B.n211 163.367
R793 B.n413 B.n206 163.367
R794 B.n422 B.n206 163.367
R795 B.n422 B.n204 163.367
R796 B.n426 B.n204 163.367
R797 B.n426 B.n199 163.367
R798 B.n435 B.n199 163.367
R799 B.n435 B.n197 163.367
R800 B.n439 B.n197 163.367
R801 B.n439 B.n192 163.367
R802 B.n448 B.n192 163.367
R803 B.n448 B.n190 163.367
R804 B.n453 B.n190 163.367
R805 B.n453 B.n184 163.367
R806 B.n461 B.n184 163.367
R807 B.n462 B.n461 163.367
R808 B.n462 B.n5 163.367
R809 B.n6 B.n5 163.367
R810 B.n7 B.n6 163.367
R811 B.n468 B.n7 163.367
R812 B.n470 B.n468 163.367
R813 B.n470 B.n12 163.367
R814 B.n13 B.n12 163.367
R815 B.n14 B.n13 163.367
R816 B.n475 B.n14 163.367
R817 B.n475 B.n19 163.367
R818 B.n20 B.n19 163.367
R819 B.n21 B.n20 163.367
R820 B.n480 B.n21 163.367
R821 B.n480 B.n26 163.367
R822 B.n27 B.n26 163.367
R823 B.n28 B.n27 163.367
R824 B.n485 B.n28 163.367
R825 B.n485 B.n33 163.367
R826 B.n34 B.n33 163.367
R827 B.n35 B.n34 163.367
R828 B.n490 B.n35 163.367
R829 B.n490 B.n40 163.367
R830 B.n41 B.n40 163.367
R831 B.n42 B.n41 163.367
R832 B.n495 B.n42 163.367
R833 B.n495 B.n47 163.367
R834 B.n48 B.n47 163.367
R835 B.n49 B.n48 163.367
R836 B.n500 B.n49 163.367
R837 B.n500 B.n54 163.367
R838 B.n55 B.n54 163.367
R839 B.n56 B.n55 163.367
R840 B.n85 B.n56 163.367
R841 B.n363 B.n240 163.367
R842 B.n363 B.n264 163.367
R843 B.n359 B.n358 163.367
R844 B.n355 B.n354 163.367
R845 B.n351 B.n350 163.367
R846 B.n347 B.n346 163.367
R847 B.n343 B.n342 163.367
R848 B.n339 B.n338 163.367
R849 B.n335 B.n334 163.367
R850 B.n331 B.n330 163.367
R851 B.n326 B.n325 163.367
R852 B.n322 B.n321 163.367
R853 B.n318 B.n317 163.367
R854 B.n314 B.n313 163.367
R855 B.n310 B.n309 163.367
R856 B.n306 B.n305 163.367
R857 B.n302 B.n301 163.367
R858 B.n298 B.n297 163.367
R859 B.n294 B.n293 163.367
R860 B.n290 B.n289 163.367
R861 B.n286 B.n285 163.367
R862 B.n282 B.n281 163.367
R863 B.n278 B.n277 163.367
R864 B.n274 B.n273 163.367
R865 B.n370 B.n238 163.367
R866 B.n370 B.n232 163.367
R867 B.n378 B.n232 163.367
R868 B.n378 B.n230 163.367
R869 B.n382 B.n230 163.367
R870 B.n382 B.n224 163.367
R871 B.n390 B.n224 163.367
R872 B.n390 B.n222 163.367
R873 B.n394 B.n222 163.367
R874 B.n394 B.n216 163.367
R875 B.n403 B.n216 163.367
R876 B.n403 B.n214 163.367
R877 B.n407 B.n214 163.367
R878 B.n407 B.n209 163.367
R879 B.n416 B.n209 163.367
R880 B.n416 B.n207 163.367
R881 B.n420 B.n207 163.367
R882 B.n420 B.n202 163.367
R883 B.n429 B.n202 163.367
R884 B.n429 B.n200 163.367
R885 B.n433 B.n200 163.367
R886 B.n433 B.n195 163.367
R887 B.n442 B.n195 163.367
R888 B.n442 B.n193 163.367
R889 B.n446 B.n193 163.367
R890 B.n446 B.n188 163.367
R891 B.n455 B.n188 163.367
R892 B.n455 B.n186 163.367
R893 B.n459 B.n186 163.367
R894 B.n459 B.n3 163.367
R895 B.n575 B.n3 163.367
R896 B.n571 B.n2 163.367
R897 B.n571 B.n570 163.367
R898 B.n570 B.n9 163.367
R899 B.n566 B.n9 163.367
R900 B.n566 B.n11 163.367
R901 B.n562 B.n11 163.367
R902 B.n562 B.n15 163.367
R903 B.n558 B.n15 163.367
R904 B.n558 B.n17 163.367
R905 B.n554 B.n17 163.367
R906 B.n554 B.n22 163.367
R907 B.n550 B.n22 163.367
R908 B.n550 B.n24 163.367
R909 B.n546 B.n24 163.367
R910 B.n546 B.n29 163.367
R911 B.n542 B.n29 163.367
R912 B.n542 B.n31 163.367
R913 B.n538 B.n31 163.367
R914 B.n538 B.n36 163.367
R915 B.n534 B.n36 163.367
R916 B.n534 B.n38 163.367
R917 B.n530 B.n38 163.367
R918 B.n530 B.n44 163.367
R919 B.n526 B.n44 163.367
R920 B.n526 B.n46 163.367
R921 B.n522 B.n46 163.367
R922 B.n522 B.n51 163.367
R923 B.n518 B.n51 163.367
R924 B.n518 B.n53 163.367
R925 B.n514 B.n53 163.367
R926 B.n514 B.n58 163.367
R927 B.n87 B.t16 155.225
R928 B.n268 B.t22 155.225
R929 B.n89 B.t13 155.225
R930 B.n266 B.t19 155.225
R931 B.n364 B.n237 143.552
R932 B.n508 B.n57 143.552
R933 B.n371 B.n237 75.6707
R934 B.n371 B.n233 75.6707
R935 B.n377 B.n233 75.6707
R936 B.n377 B.n229 75.6707
R937 B.n383 B.n229 75.6707
R938 B.n389 B.n225 75.6707
R939 B.n389 B.n221 75.6707
R940 B.n395 B.n221 75.6707
R941 B.n395 B.n217 75.6707
R942 B.n402 B.n217 75.6707
R943 B.n402 B.n401 75.6707
R944 B.n408 B.n210 75.6707
R945 B.n415 B.n210 75.6707
R946 B.n415 B.n414 75.6707
R947 B.n421 B.n203 75.6707
R948 B.n428 B.n203 75.6707
R949 B.n428 B.n427 75.6707
R950 B.n434 B.n196 75.6707
R951 B.n441 B.n196 75.6707
R952 B.n441 B.n440 75.6707
R953 B.n447 B.n189 75.6707
R954 B.n454 B.n189 75.6707
R955 B.n460 B.n185 75.6707
R956 B.n460 B.n4 75.6707
R957 B.n574 B.n4 75.6707
R958 B.n574 B.n573 75.6707
R959 B.n573 B.n572 75.6707
R960 B.n572 B.n8 75.6707
R961 B.n469 B.n8 75.6707
R962 B.n565 B.n564 75.6707
R963 B.n564 B.n563 75.6707
R964 B.n557 B.n18 75.6707
R965 B.n557 B.n556 75.6707
R966 B.n556 B.n555 75.6707
R967 B.n549 B.n25 75.6707
R968 B.n549 B.n548 75.6707
R969 B.n548 B.n547 75.6707
R970 B.n541 B.n32 75.6707
R971 B.n541 B.n540 75.6707
R972 B.n540 B.n539 75.6707
R973 B.n533 B.n39 75.6707
R974 B.n533 B.n532 75.6707
R975 B.n532 B.n531 75.6707
R976 B.n531 B.n43 75.6707
R977 B.n525 B.n43 75.6707
R978 B.n525 B.n524 75.6707
R979 B.n523 B.n50 75.6707
R980 B.n517 B.n50 75.6707
R981 B.n517 B.n516 75.6707
R982 B.n516 B.n515 75.6707
R983 B.n515 B.n57 75.6707
R984 B.n447 B.t0 73.4451
R985 B.n563 B.t8 73.4451
R986 B.n510 B.n509 71.676
R987 B.n91 B.n61 71.676
R988 B.n95 B.n62 71.676
R989 B.n99 B.n63 71.676
R990 B.n103 B.n64 71.676
R991 B.n107 B.n65 71.676
R992 B.n111 B.n66 71.676
R993 B.n115 B.n67 71.676
R994 B.n119 B.n68 71.676
R995 B.n123 B.n69 71.676
R996 B.n127 B.n70 71.676
R997 B.n131 B.n71 71.676
R998 B.n135 B.n72 71.676
R999 B.n139 B.n73 71.676
R1000 B.n143 B.n74 71.676
R1001 B.n148 B.n75 71.676
R1002 B.n152 B.n76 71.676
R1003 B.n156 B.n77 71.676
R1004 B.n160 B.n78 71.676
R1005 B.n164 B.n79 71.676
R1006 B.n168 B.n80 71.676
R1007 B.n172 B.n81 71.676
R1008 B.n176 B.n82 71.676
R1009 B.n180 B.n83 71.676
R1010 B.n84 B.n83 71.676
R1011 B.n179 B.n82 71.676
R1012 B.n175 B.n81 71.676
R1013 B.n171 B.n80 71.676
R1014 B.n167 B.n79 71.676
R1015 B.n163 B.n78 71.676
R1016 B.n159 B.n77 71.676
R1017 B.n155 B.n76 71.676
R1018 B.n151 B.n75 71.676
R1019 B.n147 B.n74 71.676
R1020 B.n142 B.n73 71.676
R1021 B.n138 B.n72 71.676
R1022 B.n134 B.n71 71.676
R1023 B.n130 B.n70 71.676
R1024 B.n126 B.n69 71.676
R1025 B.n122 B.n68 71.676
R1026 B.n118 B.n67 71.676
R1027 B.n114 B.n66 71.676
R1028 B.n110 B.n65 71.676
R1029 B.n106 B.n64 71.676
R1030 B.n102 B.n63 71.676
R1031 B.n98 B.n62 71.676
R1032 B.n94 B.n61 71.676
R1033 B.n509 B.n60 71.676
R1034 B.n366 B.n365 71.676
R1035 B.n264 B.n241 71.676
R1036 B.n358 B.n242 71.676
R1037 B.n354 B.n243 71.676
R1038 B.n350 B.n244 71.676
R1039 B.n346 B.n245 71.676
R1040 B.n342 B.n246 71.676
R1041 B.n338 B.n247 71.676
R1042 B.n334 B.n248 71.676
R1043 B.n330 B.n249 71.676
R1044 B.n325 B.n250 71.676
R1045 B.n321 B.n251 71.676
R1046 B.n317 B.n252 71.676
R1047 B.n313 B.n253 71.676
R1048 B.n309 B.n254 71.676
R1049 B.n305 B.n255 71.676
R1050 B.n301 B.n256 71.676
R1051 B.n297 B.n257 71.676
R1052 B.n293 B.n258 71.676
R1053 B.n289 B.n259 71.676
R1054 B.n285 B.n260 71.676
R1055 B.n281 B.n261 71.676
R1056 B.n277 B.n262 71.676
R1057 B.n273 B.n263 71.676
R1058 B.n365 B.n240 71.676
R1059 B.n359 B.n241 71.676
R1060 B.n355 B.n242 71.676
R1061 B.n351 B.n243 71.676
R1062 B.n347 B.n244 71.676
R1063 B.n343 B.n245 71.676
R1064 B.n339 B.n246 71.676
R1065 B.n335 B.n247 71.676
R1066 B.n331 B.n248 71.676
R1067 B.n326 B.n249 71.676
R1068 B.n322 B.n250 71.676
R1069 B.n318 B.n251 71.676
R1070 B.n314 B.n252 71.676
R1071 B.n310 B.n253 71.676
R1072 B.n306 B.n254 71.676
R1073 B.n302 B.n255 71.676
R1074 B.n298 B.n256 71.676
R1075 B.n294 B.n257 71.676
R1076 B.n290 B.n258 71.676
R1077 B.n286 B.n259 71.676
R1078 B.n282 B.n260 71.676
R1079 B.n278 B.n261 71.676
R1080 B.n274 B.n262 71.676
R1081 B.n270 B.n263 71.676
R1082 B.n576 B.n575 71.676
R1083 B.n576 B.n2 71.676
R1084 B.n454 B.t1 71.2195
R1085 B.n565 B.t2 71.2195
R1086 B.n434 B.t4 66.7683
R1087 B.n555 B.t9 66.7683
R1088 B.t18 B.n225 62.3171
R1089 B.n524 B.t11 62.3171
R1090 B.n421 B.t5 60.0915
R1091 B.n547 B.t7 60.0915
R1092 B.n90 B.n89 59.5399
R1093 B.n145 B.n87 59.5399
R1094 B.n269 B.n268 59.5399
R1095 B.n328 B.n266 59.5399
R1096 B.n408 B.t6 53.4148
R1097 B.n539 B.t3 53.4148
R1098 B.n368 B.n367 35.1225
R1099 B.n271 B.n235 35.1225
R1100 B.n512 B.n511 35.1225
R1101 B.n506 B.n505 35.1224
R1102 B.n89 B.n88 25.7944
R1103 B.n87 B.n86 25.7944
R1104 B.n268 B.n267 25.7944
R1105 B.n266 B.n265 25.7944
R1106 B.n401 B.t6 22.2564
R1107 B.n39 B.t3 22.2564
R1108 B B.n577 18.0485
R1109 B.n414 B.t5 15.5797
R1110 B.n32 B.t7 15.5797
R1111 B.n383 B.t18 13.3541
R1112 B.t11 B.n523 13.3541
R1113 B.n369 B.n368 10.6151
R1114 B.n369 B.n231 10.6151
R1115 B.n379 B.n231 10.6151
R1116 B.n380 B.n379 10.6151
R1117 B.n381 B.n380 10.6151
R1118 B.n381 B.n223 10.6151
R1119 B.n391 B.n223 10.6151
R1120 B.n392 B.n391 10.6151
R1121 B.n393 B.n392 10.6151
R1122 B.n393 B.n215 10.6151
R1123 B.n404 B.n215 10.6151
R1124 B.n405 B.n404 10.6151
R1125 B.n406 B.n405 10.6151
R1126 B.n406 B.n208 10.6151
R1127 B.n417 B.n208 10.6151
R1128 B.n418 B.n417 10.6151
R1129 B.n419 B.n418 10.6151
R1130 B.n419 B.n201 10.6151
R1131 B.n430 B.n201 10.6151
R1132 B.n431 B.n430 10.6151
R1133 B.n432 B.n431 10.6151
R1134 B.n432 B.n194 10.6151
R1135 B.n443 B.n194 10.6151
R1136 B.n444 B.n443 10.6151
R1137 B.n445 B.n444 10.6151
R1138 B.n445 B.n187 10.6151
R1139 B.n456 B.n187 10.6151
R1140 B.n457 B.n456 10.6151
R1141 B.n458 B.n457 10.6151
R1142 B.n458 B.n0 10.6151
R1143 B.n367 B.n239 10.6151
R1144 B.n362 B.n239 10.6151
R1145 B.n362 B.n361 10.6151
R1146 B.n361 B.n360 10.6151
R1147 B.n360 B.n357 10.6151
R1148 B.n357 B.n356 10.6151
R1149 B.n356 B.n353 10.6151
R1150 B.n353 B.n352 10.6151
R1151 B.n352 B.n349 10.6151
R1152 B.n349 B.n348 10.6151
R1153 B.n348 B.n345 10.6151
R1154 B.n345 B.n344 10.6151
R1155 B.n344 B.n341 10.6151
R1156 B.n341 B.n340 10.6151
R1157 B.n340 B.n337 10.6151
R1158 B.n337 B.n336 10.6151
R1159 B.n336 B.n333 10.6151
R1160 B.n333 B.n332 10.6151
R1161 B.n332 B.n329 10.6151
R1162 B.n327 B.n324 10.6151
R1163 B.n324 B.n323 10.6151
R1164 B.n323 B.n320 10.6151
R1165 B.n320 B.n319 10.6151
R1166 B.n319 B.n316 10.6151
R1167 B.n316 B.n315 10.6151
R1168 B.n315 B.n312 10.6151
R1169 B.n312 B.n311 10.6151
R1170 B.n308 B.n307 10.6151
R1171 B.n307 B.n304 10.6151
R1172 B.n304 B.n303 10.6151
R1173 B.n303 B.n300 10.6151
R1174 B.n300 B.n299 10.6151
R1175 B.n299 B.n296 10.6151
R1176 B.n296 B.n295 10.6151
R1177 B.n295 B.n292 10.6151
R1178 B.n292 B.n291 10.6151
R1179 B.n291 B.n288 10.6151
R1180 B.n288 B.n287 10.6151
R1181 B.n287 B.n284 10.6151
R1182 B.n284 B.n283 10.6151
R1183 B.n283 B.n280 10.6151
R1184 B.n280 B.n279 10.6151
R1185 B.n279 B.n276 10.6151
R1186 B.n276 B.n275 10.6151
R1187 B.n275 B.n272 10.6151
R1188 B.n272 B.n271 10.6151
R1189 B.n373 B.n235 10.6151
R1190 B.n374 B.n373 10.6151
R1191 B.n375 B.n374 10.6151
R1192 B.n375 B.n227 10.6151
R1193 B.n385 B.n227 10.6151
R1194 B.n386 B.n385 10.6151
R1195 B.n387 B.n386 10.6151
R1196 B.n387 B.n219 10.6151
R1197 B.n397 B.n219 10.6151
R1198 B.n398 B.n397 10.6151
R1199 B.n399 B.n398 10.6151
R1200 B.n399 B.n212 10.6151
R1201 B.n410 B.n212 10.6151
R1202 B.n411 B.n410 10.6151
R1203 B.n412 B.n411 10.6151
R1204 B.n412 B.n205 10.6151
R1205 B.n423 B.n205 10.6151
R1206 B.n424 B.n423 10.6151
R1207 B.n425 B.n424 10.6151
R1208 B.n425 B.n198 10.6151
R1209 B.n436 B.n198 10.6151
R1210 B.n437 B.n436 10.6151
R1211 B.n438 B.n437 10.6151
R1212 B.n438 B.n191 10.6151
R1213 B.n449 B.n191 10.6151
R1214 B.n450 B.n449 10.6151
R1215 B.n452 B.n450 10.6151
R1216 B.n452 B.n451 10.6151
R1217 B.n451 B.n183 10.6151
R1218 B.n463 B.n183 10.6151
R1219 B.n464 B.n463 10.6151
R1220 B.n465 B.n464 10.6151
R1221 B.n466 B.n465 10.6151
R1222 B.n467 B.n466 10.6151
R1223 B.n471 B.n467 10.6151
R1224 B.n472 B.n471 10.6151
R1225 B.n473 B.n472 10.6151
R1226 B.n474 B.n473 10.6151
R1227 B.n476 B.n474 10.6151
R1228 B.n477 B.n476 10.6151
R1229 B.n478 B.n477 10.6151
R1230 B.n479 B.n478 10.6151
R1231 B.n481 B.n479 10.6151
R1232 B.n482 B.n481 10.6151
R1233 B.n483 B.n482 10.6151
R1234 B.n484 B.n483 10.6151
R1235 B.n486 B.n484 10.6151
R1236 B.n487 B.n486 10.6151
R1237 B.n488 B.n487 10.6151
R1238 B.n489 B.n488 10.6151
R1239 B.n491 B.n489 10.6151
R1240 B.n492 B.n491 10.6151
R1241 B.n493 B.n492 10.6151
R1242 B.n494 B.n493 10.6151
R1243 B.n496 B.n494 10.6151
R1244 B.n497 B.n496 10.6151
R1245 B.n498 B.n497 10.6151
R1246 B.n499 B.n498 10.6151
R1247 B.n501 B.n499 10.6151
R1248 B.n502 B.n501 10.6151
R1249 B.n503 B.n502 10.6151
R1250 B.n504 B.n503 10.6151
R1251 B.n505 B.n504 10.6151
R1252 B.n569 B.n1 10.6151
R1253 B.n569 B.n568 10.6151
R1254 B.n568 B.n567 10.6151
R1255 B.n567 B.n10 10.6151
R1256 B.n561 B.n10 10.6151
R1257 B.n561 B.n560 10.6151
R1258 B.n560 B.n559 10.6151
R1259 B.n559 B.n16 10.6151
R1260 B.n553 B.n16 10.6151
R1261 B.n553 B.n552 10.6151
R1262 B.n552 B.n551 10.6151
R1263 B.n551 B.n23 10.6151
R1264 B.n545 B.n23 10.6151
R1265 B.n545 B.n544 10.6151
R1266 B.n544 B.n543 10.6151
R1267 B.n543 B.n30 10.6151
R1268 B.n537 B.n30 10.6151
R1269 B.n537 B.n536 10.6151
R1270 B.n536 B.n535 10.6151
R1271 B.n535 B.n37 10.6151
R1272 B.n529 B.n37 10.6151
R1273 B.n529 B.n528 10.6151
R1274 B.n528 B.n527 10.6151
R1275 B.n527 B.n45 10.6151
R1276 B.n521 B.n45 10.6151
R1277 B.n521 B.n520 10.6151
R1278 B.n520 B.n519 10.6151
R1279 B.n519 B.n52 10.6151
R1280 B.n513 B.n52 10.6151
R1281 B.n513 B.n512 10.6151
R1282 B.n511 B.n59 10.6151
R1283 B.n92 B.n59 10.6151
R1284 B.n93 B.n92 10.6151
R1285 B.n96 B.n93 10.6151
R1286 B.n97 B.n96 10.6151
R1287 B.n100 B.n97 10.6151
R1288 B.n101 B.n100 10.6151
R1289 B.n104 B.n101 10.6151
R1290 B.n105 B.n104 10.6151
R1291 B.n108 B.n105 10.6151
R1292 B.n109 B.n108 10.6151
R1293 B.n112 B.n109 10.6151
R1294 B.n113 B.n112 10.6151
R1295 B.n116 B.n113 10.6151
R1296 B.n117 B.n116 10.6151
R1297 B.n120 B.n117 10.6151
R1298 B.n121 B.n120 10.6151
R1299 B.n124 B.n121 10.6151
R1300 B.n125 B.n124 10.6151
R1301 B.n129 B.n128 10.6151
R1302 B.n132 B.n129 10.6151
R1303 B.n133 B.n132 10.6151
R1304 B.n136 B.n133 10.6151
R1305 B.n137 B.n136 10.6151
R1306 B.n140 B.n137 10.6151
R1307 B.n141 B.n140 10.6151
R1308 B.n144 B.n141 10.6151
R1309 B.n149 B.n146 10.6151
R1310 B.n150 B.n149 10.6151
R1311 B.n153 B.n150 10.6151
R1312 B.n154 B.n153 10.6151
R1313 B.n157 B.n154 10.6151
R1314 B.n158 B.n157 10.6151
R1315 B.n161 B.n158 10.6151
R1316 B.n162 B.n161 10.6151
R1317 B.n165 B.n162 10.6151
R1318 B.n166 B.n165 10.6151
R1319 B.n169 B.n166 10.6151
R1320 B.n170 B.n169 10.6151
R1321 B.n173 B.n170 10.6151
R1322 B.n174 B.n173 10.6151
R1323 B.n177 B.n174 10.6151
R1324 B.n178 B.n177 10.6151
R1325 B.n181 B.n178 10.6151
R1326 B.n182 B.n181 10.6151
R1327 B.n506 B.n182 10.6151
R1328 B.n427 B.t4 8.90288
R1329 B.n25 B.t9 8.90288
R1330 B.n577 B.n0 8.11757
R1331 B.n577 B.n1 8.11757
R1332 B.n328 B.n327 6.5566
R1333 B.n311 B.n269 6.5566
R1334 B.n128 B.n90 6.5566
R1335 B.n145 B.n144 6.5566
R1336 B.t1 B.n185 4.45169
R1337 B.n469 B.t2 4.45169
R1338 B.n329 B.n328 4.05904
R1339 B.n308 B.n269 4.05904
R1340 B.n125 B.n90 4.05904
R1341 B.n146 B.n145 4.05904
R1342 B.n440 B.t0 2.22609
R1343 B.n18 B.t8 2.22609
R1344 VN.n5 VN.t3 164.95
R1345 VN.n25 VN.t6 164.95
R1346 VN.n37 VN.n20 161.3
R1347 VN.n35 VN.n34 161.3
R1348 VN.n33 VN.n21 161.3
R1349 VN.n32 VN.n31 161.3
R1350 VN.n29 VN.n22 161.3
R1351 VN.n28 VN.n27 161.3
R1352 VN.n26 VN.n23 161.3
R1353 VN.n17 VN.n0 161.3
R1354 VN.n15 VN.n14 161.3
R1355 VN.n13 VN.n1 161.3
R1356 VN.n12 VN.n11 161.3
R1357 VN.n9 VN.n2 161.3
R1358 VN.n8 VN.n7 161.3
R1359 VN.n6 VN.n3 161.3
R1360 VN.n18 VN.t0 150.625
R1361 VN.n38 VN.t1 150.625
R1362 VN.n4 VN.t2 111.102
R1363 VN.n10 VN.t5 111.102
R1364 VN.n16 VN.t4 111.102
R1365 VN.n24 VN.t8 111.102
R1366 VN.n30 VN.t7 111.102
R1367 VN.n36 VN.t9 111.102
R1368 VN.n39 VN.n38 80.6037
R1369 VN.n19 VN.n18 80.6037
R1370 VN.n18 VN.n17 52.1152
R1371 VN.n38 VN.n37 52.1152
R1372 VN.n5 VN.n4 49.1161
R1373 VN.n25 VN.n24 49.1161
R1374 VN.n9 VN.n8 48.7492
R1375 VN.n11 VN.n1 48.7492
R1376 VN.n29 VN.n28 48.7492
R1377 VN.n31 VN.n21 48.7492
R1378 VN.n26 VN.n25 44.523
R1379 VN.n6 VN.n5 44.523
R1380 VN VN.n39 39.2528
R1381 VN.n8 VN.n3 32.2376
R1382 VN.n15 VN.n1 32.2376
R1383 VN.n28 VN.n23 32.2376
R1384 VN.n35 VN.n21 32.2376
R1385 VN.n17 VN.n16 20.5528
R1386 VN.n37 VN.n36 20.5528
R1387 VN.n10 VN.n9 12.234
R1388 VN.n11 VN.n10 12.234
R1389 VN.n31 VN.n30 12.234
R1390 VN.n30 VN.n29 12.234
R1391 VN.n4 VN.n3 3.91522
R1392 VN.n16 VN.n15 3.91522
R1393 VN.n24 VN.n23 3.91522
R1394 VN.n36 VN.n35 3.91522
R1395 VN.n39 VN.n20 0.285035
R1396 VN.n19 VN.n0 0.285035
R1397 VN.n34 VN.n20 0.189894
R1398 VN.n34 VN.n33 0.189894
R1399 VN.n33 VN.n32 0.189894
R1400 VN.n32 VN.n22 0.189894
R1401 VN.n27 VN.n22 0.189894
R1402 VN.n27 VN.n26 0.189894
R1403 VN.n7 VN.n6 0.189894
R1404 VN.n7 VN.n2 0.189894
R1405 VN.n12 VN.n2 0.189894
R1406 VN.n13 VN.n12 0.189894
R1407 VN.n14 VN.n13 0.189894
R1408 VN.n14 VN.n0 0.189894
R1409 VN VN.n19 0.146778
R1410 VDD2.n45 VDD2.n27 289.615
R1411 VDD2.n18 VDD2.n0 289.615
R1412 VDD2.n46 VDD2.n45 185
R1413 VDD2.n44 VDD2.n43 185
R1414 VDD2.n31 VDD2.n30 185
R1415 VDD2.n38 VDD2.n37 185
R1416 VDD2.n36 VDD2.n35 185
R1417 VDD2.n9 VDD2.n8 185
R1418 VDD2.n11 VDD2.n10 185
R1419 VDD2.n4 VDD2.n3 185
R1420 VDD2.n17 VDD2.n16 185
R1421 VDD2.n19 VDD2.n18 185
R1422 VDD2.n34 VDD2.t8 147.714
R1423 VDD2.n7 VDD2.t6 147.714
R1424 VDD2.n45 VDD2.n44 104.615
R1425 VDD2.n44 VDD2.n30 104.615
R1426 VDD2.n37 VDD2.n30 104.615
R1427 VDD2.n37 VDD2.n36 104.615
R1428 VDD2.n10 VDD2.n9 104.615
R1429 VDD2.n10 VDD2.n3 104.615
R1430 VDD2.n17 VDD2.n3 104.615
R1431 VDD2.n18 VDD2.n17 104.615
R1432 VDD2.n26 VDD2.n25 72.4159
R1433 VDD2 VDD2.n53 72.4131
R1434 VDD2.n52 VDD2.n51 71.6115
R1435 VDD2.n24 VDD2.n23 71.6113
R1436 VDD2.n36 VDD2.t8 52.3082
R1437 VDD2.n9 VDD2.t6 52.3082
R1438 VDD2.n24 VDD2.n22 50.9804
R1439 VDD2.n50 VDD2.n49 49.8338
R1440 VDD2.n50 VDD2.n26 33.1356
R1441 VDD2.n35 VDD2.n34 15.6631
R1442 VDD2.n8 VDD2.n7 15.6631
R1443 VDD2.n38 VDD2.n33 12.8005
R1444 VDD2.n11 VDD2.n6 12.8005
R1445 VDD2.n39 VDD2.n31 12.0247
R1446 VDD2.n12 VDD2.n4 12.0247
R1447 VDD2.n43 VDD2.n42 11.249
R1448 VDD2.n16 VDD2.n15 11.249
R1449 VDD2.n46 VDD2.n29 10.4732
R1450 VDD2.n19 VDD2.n2 10.4732
R1451 VDD2.n47 VDD2.n27 9.69747
R1452 VDD2.n20 VDD2.n0 9.69747
R1453 VDD2.n49 VDD2.n48 9.45567
R1454 VDD2.n22 VDD2.n21 9.45567
R1455 VDD2.n48 VDD2.n47 9.3005
R1456 VDD2.n29 VDD2.n28 9.3005
R1457 VDD2.n42 VDD2.n41 9.3005
R1458 VDD2.n40 VDD2.n39 9.3005
R1459 VDD2.n33 VDD2.n32 9.3005
R1460 VDD2.n21 VDD2.n20 9.3005
R1461 VDD2.n2 VDD2.n1 9.3005
R1462 VDD2.n15 VDD2.n14 9.3005
R1463 VDD2.n13 VDD2.n12 9.3005
R1464 VDD2.n6 VDD2.n5 9.3005
R1465 VDD2.n34 VDD2.n32 4.39059
R1466 VDD2.n7 VDD2.n5 4.39059
R1467 VDD2.n53 VDD2.t1 4.29551
R1468 VDD2.n53 VDD2.t3 4.29551
R1469 VDD2.n51 VDD2.t0 4.29551
R1470 VDD2.n51 VDD2.t2 4.29551
R1471 VDD2.n25 VDD2.t5 4.29551
R1472 VDD2.n25 VDD2.t9 4.29551
R1473 VDD2.n23 VDD2.t7 4.29551
R1474 VDD2.n23 VDD2.t4 4.29551
R1475 VDD2.n49 VDD2.n27 4.26717
R1476 VDD2.n22 VDD2.n0 4.26717
R1477 VDD2.n47 VDD2.n46 3.49141
R1478 VDD2.n20 VDD2.n19 3.49141
R1479 VDD2.n43 VDD2.n29 2.71565
R1480 VDD2.n16 VDD2.n2 2.71565
R1481 VDD2.n42 VDD2.n31 1.93989
R1482 VDD2.n15 VDD2.n4 1.93989
R1483 VDD2.n39 VDD2.n38 1.16414
R1484 VDD2.n12 VDD2.n11 1.16414
R1485 VDD2.n52 VDD2.n50 1.14705
R1486 VDD2.n35 VDD2.n33 0.388379
R1487 VDD2.n8 VDD2.n6 0.388379
R1488 VDD2 VDD2.n52 0.345328
R1489 VDD2.n26 VDD2.n24 0.231792
R1490 VDD2.n48 VDD2.n28 0.155672
R1491 VDD2.n41 VDD2.n28 0.155672
R1492 VDD2.n41 VDD2.n40 0.155672
R1493 VDD2.n40 VDD2.n32 0.155672
R1494 VDD2.n13 VDD2.n5 0.155672
R1495 VDD2.n14 VDD2.n13 0.155672
R1496 VDD2.n14 VDD2.n1 0.155672
R1497 VDD2.n21 VDD2.n1 0.155672
C0 VDD1 VTAIL 6.50221f
C1 VDD1 VDD2 1.15947f
C2 VTAIL VP 3.71214f
C3 VDD2 VP 0.383074f
C4 VTAIL VDD2 6.54295f
C5 VDD1 VN 0.153679f
C6 VP VN 4.6772f
C7 VDD1 VP 3.55844f
C8 VTAIL VN 3.69787f
C9 VDD2 VN 3.33162f
C10 VDD2 B 3.989209f
C11 VDD1 B 3.942739f
C12 VTAIL B 3.860196f
C13 VN B 9.89332f
C14 VP B 8.321318f
C15 VDD2.n0 B 0.032418f
C16 VDD2.n1 B 0.0234f
C17 VDD2.n2 B 0.012574f
C18 VDD2.n3 B 0.029721f
C19 VDD2.n4 B 0.013314f
C20 VDD2.n5 B 0.406481f
C21 VDD2.n6 B 0.012574f
C22 VDD2.t6 B 0.048772f
C23 VDD2.n7 B 0.092798f
C24 VDD2.n8 B 0.01754f
C25 VDD2.n9 B 0.022291f
C26 VDD2.n10 B 0.029721f
C27 VDD2.n11 B 0.013314f
C28 VDD2.n12 B 0.012574f
C29 VDD2.n13 B 0.0234f
C30 VDD2.n14 B 0.0234f
C31 VDD2.n15 B 0.012574f
C32 VDD2.n16 B 0.013314f
C33 VDD2.n17 B 0.029721f
C34 VDD2.n18 B 0.063504f
C35 VDD2.n19 B 0.013314f
C36 VDD2.n20 B 0.012574f
C37 VDD2.n21 B 0.055688f
C38 VDD2.n22 B 0.054619f
C39 VDD2.t7 B 0.085247f
C40 VDD2.t4 B 0.085247f
C41 VDD2.n23 B 0.685899f
C42 VDD2.n24 B 0.420471f
C43 VDD2.t5 B 0.085247f
C44 VDD2.t9 B 0.085247f
C45 VDD2.n25 B 0.689699f
C46 VDD2.n26 B 1.51314f
C47 VDD2.n27 B 0.032418f
C48 VDD2.n28 B 0.0234f
C49 VDD2.n29 B 0.012574f
C50 VDD2.n30 B 0.029721f
C51 VDD2.n31 B 0.013314f
C52 VDD2.n32 B 0.406481f
C53 VDD2.n33 B 0.012574f
C54 VDD2.t8 B 0.048772f
C55 VDD2.n34 B 0.092798f
C56 VDD2.n35 B 0.01754f
C57 VDD2.n36 B 0.022291f
C58 VDD2.n37 B 0.029721f
C59 VDD2.n38 B 0.013314f
C60 VDD2.n39 B 0.012574f
C61 VDD2.n40 B 0.0234f
C62 VDD2.n41 B 0.0234f
C63 VDD2.n42 B 0.012574f
C64 VDD2.n43 B 0.013314f
C65 VDD2.n44 B 0.029721f
C66 VDD2.n45 B 0.063504f
C67 VDD2.n46 B 0.013314f
C68 VDD2.n47 B 0.012574f
C69 VDD2.n48 B 0.055688f
C70 VDD2.n49 B 0.051641f
C71 VDD2.n50 B 1.57598f
C72 VDD2.t0 B 0.085247f
C73 VDD2.t2 B 0.085247f
C74 VDD2.n51 B 0.685903f
C75 VDD2.n52 B 0.297234f
C76 VDD2.t1 B 0.085247f
C77 VDD2.t3 B 0.085247f
C78 VDD2.n53 B 0.689676f
C79 VN.n0 B 0.051996f
C80 VN.t4 B 0.46702f
C81 VN.n1 B 0.035275f
C82 VN.n2 B 0.038966f
C83 VN.t5 B 0.46702f
C84 VN.n3 B 0.048382f
C85 VN.t3 B 0.549518f
C86 VN.t2 B 0.46702f
C87 VN.n4 B 0.232395f
C88 VN.n5 B 0.260969f
C89 VN.n6 B 0.162769f
C90 VN.n7 B 0.038966f
C91 VN.n8 B 0.035275f
C92 VN.n9 B 0.054696f
C93 VN.n10 B 0.203662f
C94 VN.n11 B 0.054696f
C95 VN.n12 B 0.038966f
C96 VN.n13 B 0.038966f
C97 VN.n14 B 0.038966f
C98 VN.n15 B 0.048382f
C99 VN.n16 B 0.203662f
C100 VN.n17 B 0.049407f
C101 VN.t0 B 0.526717f
C102 VN.n18 B 0.262311f
C103 VN.n19 B 0.036494f
C104 VN.n20 B 0.051996f
C105 VN.t9 B 0.46702f
C106 VN.n21 B 0.035275f
C107 VN.n22 B 0.038966f
C108 VN.t7 B 0.46702f
C109 VN.n23 B 0.048382f
C110 VN.t6 B 0.549518f
C111 VN.t8 B 0.46702f
C112 VN.n24 B 0.232395f
C113 VN.n25 B 0.260969f
C114 VN.n26 B 0.162769f
C115 VN.n27 B 0.038966f
C116 VN.n28 B 0.035275f
C117 VN.n29 B 0.054696f
C118 VN.n30 B 0.203662f
C119 VN.n31 B 0.054696f
C120 VN.n32 B 0.038966f
C121 VN.n33 B 0.038966f
C122 VN.n34 B 0.038966f
C123 VN.n35 B 0.048382f
C124 VN.n36 B 0.203662f
C125 VN.n37 B 0.049407f
C126 VN.t1 B 0.526717f
C127 VN.n38 B 0.262311f
C128 VN.n39 B 1.45079f
C129 VDD1.n0 B 0.033118f
C130 VDD1.n1 B 0.023906f
C131 VDD1.n2 B 0.012846f
C132 VDD1.n3 B 0.030363f
C133 VDD1.n4 B 0.013602f
C134 VDD1.n5 B 0.415262f
C135 VDD1.n6 B 0.012846f
C136 VDD1.t0 B 0.049826f
C137 VDD1.n7 B 0.094803f
C138 VDD1.n8 B 0.017919f
C139 VDD1.n9 B 0.022773f
C140 VDD1.n10 B 0.030363f
C141 VDD1.n11 B 0.013602f
C142 VDD1.n12 B 0.012846f
C143 VDD1.n13 B 0.023906f
C144 VDD1.n14 B 0.023906f
C145 VDD1.n15 B 0.012846f
C146 VDD1.n16 B 0.013602f
C147 VDD1.n17 B 0.030363f
C148 VDD1.n18 B 0.064876f
C149 VDD1.n19 B 0.013602f
C150 VDD1.n20 B 0.012846f
C151 VDD1.n21 B 0.056891f
C152 VDD1.n22 B 0.055799f
C153 VDD1.t8 B 0.087089f
C154 VDD1.t9 B 0.087089f
C155 VDD1.n23 B 0.70072f
C156 VDD1.n24 B 0.4359f
C157 VDD1.n25 B 0.033118f
C158 VDD1.n26 B 0.023906f
C159 VDD1.n27 B 0.012846f
C160 VDD1.n28 B 0.030363f
C161 VDD1.n29 B 0.013602f
C162 VDD1.n30 B 0.415262f
C163 VDD1.n31 B 0.012846f
C164 VDD1.t1 B 0.049826f
C165 VDD1.n32 B 0.094803f
C166 VDD1.n33 B 0.017919f
C167 VDD1.n34 B 0.022773f
C168 VDD1.n35 B 0.030363f
C169 VDD1.n36 B 0.013602f
C170 VDD1.n37 B 0.012846f
C171 VDD1.n38 B 0.023906f
C172 VDD1.n39 B 0.023906f
C173 VDD1.n40 B 0.012846f
C174 VDD1.n41 B 0.013602f
C175 VDD1.n42 B 0.030363f
C176 VDD1.n43 B 0.064876f
C177 VDD1.n44 B 0.013602f
C178 VDD1.n45 B 0.012846f
C179 VDD1.n46 B 0.056891f
C180 VDD1.n47 B 0.055799f
C181 VDD1.t6 B 0.087089f
C182 VDD1.t2 B 0.087089f
C183 VDD1.n48 B 0.700716f
C184 VDD1.n49 B 0.429554f
C185 VDD1.t5 B 0.087089f
C186 VDD1.t4 B 0.087089f
C187 VDD1.n50 B 0.704598f
C188 VDD1.n51 B 1.62256f
C189 VDD1.t7 B 0.087089f
C190 VDD1.t3 B 0.087089f
C191 VDD1.n52 B 0.700716f
C192 VDD1.n53 B 1.83478f
C193 VTAIL.t2 B 0.102014f
C194 VTAIL.t18 B 0.102014f
C195 VTAIL.n0 B 0.755282f
C196 VTAIL.n1 B 0.425553f
C197 VTAIL.n2 B 0.038794f
C198 VTAIL.n3 B 0.028003f
C199 VTAIL.n4 B 0.015048f
C200 VTAIL.n5 B 0.035567f
C201 VTAIL.n6 B 0.015933f
C202 VTAIL.n7 B 0.486429f
C203 VTAIL.n8 B 0.015048f
C204 VTAIL.t16 B 0.058365f
C205 VTAIL.n9 B 0.11105f
C206 VTAIL.n10 B 0.02099f
C207 VTAIL.n11 B 0.026675f
C208 VTAIL.n12 B 0.035567f
C209 VTAIL.n13 B 0.015933f
C210 VTAIL.n14 B 0.015048f
C211 VTAIL.n15 B 0.028003f
C212 VTAIL.n16 B 0.028003f
C213 VTAIL.n17 B 0.015048f
C214 VTAIL.n18 B 0.015933f
C215 VTAIL.n19 B 0.035567f
C216 VTAIL.n20 B 0.075994f
C217 VTAIL.n21 B 0.015933f
C218 VTAIL.n22 B 0.015048f
C219 VTAIL.n23 B 0.06664f
C220 VTAIL.n24 B 0.042477f
C221 VTAIL.n25 B 0.222574f
C222 VTAIL.t13 B 0.102014f
C223 VTAIL.t10 B 0.102014f
C224 VTAIL.n26 B 0.755282f
C225 VTAIL.n27 B 0.4555f
C226 VTAIL.t11 B 0.102014f
C227 VTAIL.t14 B 0.102014f
C228 VTAIL.n28 B 0.755282f
C229 VTAIL.n29 B 1.29794f
C230 VTAIL.t6 B 0.102014f
C231 VTAIL.t5 B 0.102014f
C232 VTAIL.n30 B 0.755288f
C233 VTAIL.n31 B 1.29793f
C234 VTAIL.t4 B 0.102014f
C235 VTAIL.t0 B 0.102014f
C236 VTAIL.n32 B 0.755288f
C237 VTAIL.n33 B 0.455495f
C238 VTAIL.n34 B 0.038794f
C239 VTAIL.n35 B 0.028003f
C240 VTAIL.n36 B 0.015048f
C241 VTAIL.n37 B 0.035567f
C242 VTAIL.n38 B 0.015933f
C243 VTAIL.n39 B 0.486429f
C244 VTAIL.n40 B 0.015048f
C245 VTAIL.t1 B 0.058365f
C246 VTAIL.n41 B 0.11105f
C247 VTAIL.n42 B 0.02099f
C248 VTAIL.n43 B 0.026675f
C249 VTAIL.n44 B 0.035567f
C250 VTAIL.n45 B 0.015933f
C251 VTAIL.n46 B 0.015048f
C252 VTAIL.n47 B 0.028003f
C253 VTAIL.n48 B 0.028003f
C254 VTAIL.n49 B 0.015048f
C255 VTAIL.n50 B 0.015933f
C256 VTAIL.n51 B 0.035567f
C257 VTAIL.n52 B 0.075994f
C258 VTAIL.n53 B 0.015933f
C259 VTAIL.n54 B 0.015048f
C260 VTAIL.n55 B 0.06664f
C261 VTAIL.n56 B 0.042477f
C262 VTAIL.n57 B 0.222574f
C263 VTAIL.t9 B 0.102014f
C264 VTAIL.t8 B 0.102014f
C265 VTAIL.n58 B 0.755288f
C266 VTAIL.n59 B 0.446161f
C267 VTAIL.t12 B 0.102014f
C268 VTAIL.t15 B 0.102014f
C269 VTAIL.n60 B 0.755288f
C270 VTAIL.n61 B 0.455495f
C271 VTAIL.n62 B 0.038794f
C272 VTAIL.n63 B 0.028003f
C273 VTAIL.n64 B 0.015048f
C274 VTAIL.n65 B 0.035567f
C275 VTAIL.n66 B 0.015933f
C276 VTAIL.n67 B 0.486429f
C277 VTAIL.n68 B 0.015048f
C278 VTAIL.t7 B 0.058365f
C279 VTAIL.n69 B 0.11105f
C280 VTAIL.n70 B 0.02099f
C281 VTAIL.n71 B 0.026675f
C282 VTAIL.n72 B 0.035567f
C283 VTAIL.n73 B 0.015933f
C284 VTAIL.n74 B 0.015048f
C285 VTAIL.n75 B 0.028003f
C286 VTAIL.n76 B 0.028003f
C287 VTAIL.n77 B 0.015048f
C288 VTAIL.n78 B 0.015933f
C289 VTAIL.n79 B 0.035567f
C290 VTAIL.n80 B 0.075994f
C291 VTAIL.n81 B 0.015933f
C292 VTAIL.n82 B 0.015048f
C293 VTAIL.n83 B 0.06664f
C294 VTAIL.n84 B 0.042477f
C295 VTAIL.n85 B 0.970891f
C296 VTAIL.n86 B 0.038794f
C297 VTAIL.n87 B 0.028003f
C298 VTAIL.n88 B 0.015048f
C299 VTAIL.n89 B 0.035567f
C300 VTAIL.n90 B 0.015933f
C301 VTAIL.n91 B 0.486429f
C302 VTAIL.n92 B 0.015048f
C303 VTAIL.t3 B 0.058365f
C304 VTAIL.n93 B 0.11105f
C305 VTAIL.n94 B 0.02099f
C306 VTAIL.n95 B 0.026675f
C307 VTAIL.n96 B 0.035567f
C308 VTAIL.n97 B 0.015933f
C309 VTAIL.n98 B 0.015048f
C310 VTAIL.n99 B 0.028003f
C311 VTAIL.n100 B 0.028003f
C312 VTAIL.n101 B 0.015048f
C313 VTAIL.n102 B 0.015933f
C314 VTAIL.n103 B 0.035567f
C315 VTAIL.n104 B 0.075994f
C316 VTAIL.n105 B 0.015933f
C317 VTAIL.n106 B 0.015048f
C318 VTAIL.n107 B 0.06664f
C319 VTAIL.n108 B 0.042477f
C320 VTAIL.n109 B 0.970891f
C321 VTAIL.t19 B 0.102014f
C322 VTAIL.t17 B 0.102014f
C323 VTAIL.n110 B 0.755282f
C324 VTAIL.n111 B 0.372658f
C325 VP.n0 B 0.05358f
C326 VP.t4 B 0.481248f
C327 VP.n1 B 0.03635f
C328 VP.n2 B 0.040153f
C329 VP.t7 B 0.481248f
C330 VP.n3 B 0.049856f
C331 VP.n4 B 0.05358f
C332 VP.t6 B 0.542764f
C333 VP.t2 B 0.481248f
C334 VP.n5 B 0.03635f
C335 VP.n6 B 0.040153f
C336 VP.t0 B 0.481248f
C337 VP.n7 B 0.049856f
C338 VP.t1 B 0.481248f
C339 VP.n8 B 0.239475f
C340 VP.t9 B 0.56626f
C341 VP.n9 B 0.268919f
C342 VP.n10 B 0.167728f
C343 VP.n11 B 0.040153f
C344 VP.n12 B 0.03635f
C345 VP.n13 B 0.056362f
C346 VP.n14 B 0.209866f
C347 VP.n15 B 0.056362f
C348 VP.n16 B 0.040153f
C349 VP.n17 B 0.040153f
C350 VP.n18 B 0.040153f
C351 VP.n19 B 0.049856f
C352 VP.n20 B 0.209866f
C353 VP.n21 B 0.050912f
C354 VP.n22 B 0.270303f
C355 VP.n23 B 1.47216f
C356 VP.n24 B 1.5092f
C357 VP.t8 B 0.542764f
C358 VP.n25 B 0.270303f
C359 VP.t3 B 0.481248f
C360 VP.n26 B 0.209866f
C361 VP.n27 B 0.050912f
C362 VP.n28 B 0.05358f
C363 VP.n29 B 0.040153f
C364 VP.n30 B 0.040153f
C365 VP.n31 B 0.03635f
C366 VP.n32 B 0.056362f
C367 VP.n33 B 0.209866f
C368 VP.n34 B 0.056362f
C369 VP.n35 B 0.040153f
C370 VP.n36 B 0.040153f
C371 VP.n37 B 0.040153f
C372 VP.n38 B 0.049856f
C373 VP.n39 B 0.209866f
C374 VP.n40 B 0.050912f
C375 VP.t5 B 0.542764f
C376 VP.n41 B 0.270303f
C377 VP.n42 B 0.037605f
.ends

