* NGSPICE file created from diff_pair_sample_1344.ext - technology: sky130A

.subckt diff_pair_sample_1344 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=0 ps=0 w=9.01 l=2.12
X1 VTAIL.t7 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=1.48665 ps=9.34 w=9.01 l=2.12
X2 VDD1.t0 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48665 pd=9.34 as=3.5139 ps=18.8 w=9.01 l=2.12
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=1.48665 ps=9.34 w=9.01 l=2.12
X4 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48665 pd=9.34 as=3.5139 ps=18.8 w=9.01 l=2.12
X5 VDD1.t2 VP.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.48665 pd=9.34 as=3.5139 ps=18.8 w=9.01 l=2.12
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=0 ps=0 w=9.01 l=2.12
X7 VTAIL.t4 VP.t3 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=1.48665 ps=9.34 w=9.01 l=2.12
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.48665 pd=9.34 as=3.5139 ps=18.8 w=9.01 l=2.12
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=1.48665 ps=9.34 w=9.01 l=2.12
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=0 ps=0 w=9.01 l=2.12
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5139 pd=18.8 as=0 ps=0 w=9.01 l=2.12
R0 B.n624 B.n623 585
R1 B.n625 B.n624 585
R2 B.n247 B.n94 585
R3 B.n246 B.n245 585
R4 B.n244 B.n243 585
R5 B.n242 B.n241 585
R6 B.n240 B.n239 585
R7 B.n238 B.n237 585
R8 B.n236 B.n235 585
R9 B.n234 B.n233 585
R10 B.n232 B.n231 585
R11 B.n230 B.n229 585
R12 B.n228 B.n227 585
R13 B.n226 B.n225 585
R14 B.n224 B.n223 585
R15 B.n222 B.n221 585
R16 B.n220 B.n219 585
R17 B.n218 B.n217 585
R18 B.n216 B.n215 585
R19 B.n214 B.n213 585
R20 B.n212 B.n211 585
R21 B.n210 B.n209 585
R22 B.n208 B.n207 585
R23 B.n206 B.n205 585
R24 B.n204 B.n203 585
R25 B.n202 B.n201 585
R26 B.n200 B.n199 585
R27 B.n198 B.n197 585
R28 B.n196 B.n195 585
R29 B.n194 B.n193 585
R30 B.n192 B.n191 585
R31 B.n190 B.n189 585
R32 B.n188 B.n187 585
R33 B.n186 B.n185 585
R34 B.n184 B.n183 585
R35 B.n182 B.n181 585
R36 B.n180 B.n179 585
R37 B.n178 B.n177 585
R38 B.n176 B.n175 585
R39 B.n174 B.n173 585
R40 B.n172 B.n171 585
R41 B.n170 B.n169 585
R42 B.n168 B.n167 585
R43 B.n165 B.n164 585
R44 B.n163 B.n162 585
R45 B.n161 B.n160 585
R46 B.n159 B.n158 585
R47 B.n157 B.n156 585
R48 B.n155 B.n154 585
R49 B.n153 B.n152 585
R50 B.n151 B.n150 585
R51 B.n149 B.n148 585
R52 B.n147 B.n146 585
R53 B.n145 B.n144 585
R54 B.n143 B.n142 585
R55 B.n141 B.n140 585
R56 B.n139 B.n138 585
R57 B.n137 B.n136 585
R58 B.n135 B.n134 585
R59 B.n133 B.n132 585
R60 B.n131 B.n130 585
R61 B.n129 B.n128 585
R62 B.n127 B.n126 585
R63 B.n125 B.n124 585
R64 B.n123 B.n122 585
R65 B.n121 B.n120 585
R66 B.n119 B.n118 585
R67 B.n117 B.n116 585
R68 B.n115 B.n114 585
R69 B.n113 B.n112 585
R70 B.n111 B.n110 585
R71 B.n109 B.n108 585
R72 B.n107 B.n106 585
R73 B.n105 B.n104 585
R74 B.n103 B.n102 585
R75 B.n101 B.n100 585
R76 B.n622 B.n56 585
R77 B.n626 B.n56 585
R78 B.n621 B.n55 585
R79 B.n627 B.n55 585
R80 B.n620 B.n619 585
R81 B.n619 B.n51 585
R82 B.n618 B.n50 585
R83 B.n633 B.n50 585
R84 B.n617 B.n49 585
R85 B.n634 B.n49 585
R86 B.n616 B.n48 585
R87 B.n635 B.n48 585
R88 B.n615 B.n614 585
R89 B.n614 B.n47 585
R90 B.n613 B.n43 585
R91 B.n641 B.n43 585
R92 B.n612 B.n42 585
R93 B.n642 B.n42 585
R94 B.n611 B.n41 585
R95 B.n643 B.n41 585
R96 B.n610 B.n609 585
R97 B.n609 B.n37 585
R98 B.n608 B.n36 585
R99 B.n649 B.n36 585
R100 B.n607 B.n35 585
R101 B.n650 B.n35 585
R102 B.n606 B.n34 585
R103 B.n651 B.n34 585
R104 B.n605 B.n604 585
R105 B.n604 B.n30 585
R106 B.n603 B.n29 585
R107 B.n657 B.n29 585
R108 B.n602 B.n28 585
R109 B.n658 B.n28 585
R110 B.n601 B.n27 585
R111 B.n659 B.n27 585
R112 B.n600 B.n599 585
R113 B.n599 B.n23 585
R114 B.n598 B.n22 585
R115 B.n665 B.n22 585
R116 B.n597 B.n21 585
R117 B.n666 B.n21 585
R118 B.n596 B.n20 585
R119 B.n667 B.n20 585
R120 B.n595 B.n594 585
R121 B.n594 B.n16 585
R122 B.n593 B.n15 585
R123 B.n673 B.n15 585
R124 B.n592 B.n14 585
R125 B.n674 B.n14 585
R126 B.n591 B.n13 585
R127 B.n675 B.n13 585
R128 B.n590 B.n589 585
R129 B.n589 B.n12 585
R130 B.n588 B.n587 585
R131 B.n588 B.n8 585
R132 B.n586 B.n7 585
R133 B.n682 B.n7 585
R134 B.n585 B.n6 585
R135 B.n683 B.n6 585
R136 B.n584 B.n5 585
R137 B.n684 B.n5 585
R138 B.n583 B.n582 585
R139 B.n582 B.n4 585
R140 B.n581 B.n248 585
R141 B.n581 B.n580 585
R142 B.n571 B.n249 585
R143 B.n250 B.n249 585
R144 B.n573 B.n572 585
R145 B.n574 B.n573 585
R146 B.n570 B.n254 585
R147 B.n258 B.n254 585
R148 B.n569 B.n568 585
R149 B.n568 B.n567 585
R150 B.n256 B.n255 585
R151 B.n257 B.n256 585
R152 B.n560 B.n559 585
R153 B.n561 B.n560 585
R154 B.n558 B.n263 585
R155 B.n263 B.n262 585
R156 B.n557 B.n556 585
R157 B.n556 B.n555 585
R158 B.n265 B.n264 585
R159 B.n266 B.n265 585
R160 B.n548 B.n547 585
R161 B.n549 B.n548 585
R162 B.n546 B.n271 585
R163 B.n271 B.n270 585
R164 B.n545 B.n544 585
R165 B.n544 B.n543 585
R166 B.n273 B.n272 585
R167 B.n274 B.n273 585
R168 B.n536 B.n535 585
R169 B.n537 B.n536 585
R170 B.n534 B.n279 585
R171 B.n279 B.n278 585
R172 B.n533 B.n532 585
R173 B.n532 B.n531 585
R174 B.n281 B.n280 585
R175 B.n282 B.n281 585
R176 B.n524 B.n523 585
R177 B.n525 B.n524 585
R178 B.n522 B.n287 585
R179 B.n287 B.n286 585
R180 B.n521 B.n520 585
R181 B.n520 B.n519 585
R182 B.n289 B.n288 585
R183 B.n512 B.n289 585
R184 B.n511 B.n510 585
R185 B.n513 B.n511 585
R186 B.n509 B.n294 585
R187 B.n294 B.n293 585
R188 B.n508 B.n507 585
R189 B.n507 B.n506 585
R190 B.n296 B.n295 585
R191 B.n297 B.n296 585
R192 B.n499 B.n498 585
R193 B.n500 B.n499 585
R194 B.n497 B.n302 585
R195 B.n302 B.n301 585
R196 B.n491 B.n490 585
R197 B.n489 B.n341 585
R198 B.n488 B.n340 585
R199 B.n493 B.n340 585
R200 B.n487 B.n486 585
R201 B.n485 B.n484 585
R202 B.n483 B.n482 585
R203 B.n481 B.n480 585
R204 B.n479 B.n478 585
R205 B.n477 B.n476 585
R206 B.n475 B.n474 585
R207 B.n473 B.n472 585
R208 B.n471 B.n470 585
R209 B.n469 B.n468 585
R210 B.n467 B.n466 585
R211 B.n465 B.n464 585
R212 B.n463 B.n462 585
R213 B.n461 B.n460 585
R214 B.n459 B.n458 585
R215 B.n457 B.n456 585
R216 B.n455 B.n454 585
R217 B.n453 B.n452 585
R218 B.n451 B.n450 585
R219 B.n449 B.n448 585
R220 B.n447 B.n446 585
R221 B.n445 B.n444 585
R222 B.n443 B.n442 585
R223 B.n441 B.n440 585
R224 B.n439 B.n438 585
R225 B.n437 B.n436 585
R226 B.n435 B.n434 585
R227 B.n433 B.n432 585
R228 B.n431 B.n430 585
R229 B.n429 B.n428 585
R230 B.n427 B.n426 585
R231 B.n425 B.n424 585
R232 B.n423 B.n422 585
R233 B.n421 B.n420 585
R234 B.n419 B.n418 585
R235 B.n417 B.n416 585
R236 B.n415 B.n414 585
R237 B.n413 B.n412 585
R238 B.n411 B.n410 585
R239 B.n408 B.n407 585
R240 B.n406 B.n405 585
R241 B.n404 B.n403 585
R242 B.n402 B.n401 585
R243 B.n400 B.n399 585
R244 B.n398 B.n397 585
R245 B.n396 B.n395 585
R246 B.n394 B.n393 585
R247 B.n392 B.n391 585
R248 B.n390 B.n389 585
R249 B.n388 B.n387 585
R250 B.n386 B.n385 585
R251 B.n384 B.n383 585
R252 B.n382 B.n381 585
R253 B.n380 B.n379 585
R254 B.n378 B.n377 585
R255 B.n376 B.n375 585
R256 B.n374 B.n373 585
R257 B.n372 B.n371 585
R258 B.n370 B.n369 585
R259 B.n368 B.n367 585
R260 B.n366 B.n365 585
R261 B.n364 B.n363 585
R262 B.n362 B.n361 585
R263 B.n360 B.n359 585
R264 B.n358 B.n357 585
R265 B.n356 B.n355 585
R266 B.n354 B.n353 585
R267 B.n352 B.n351 585
R268 B.n350 B.n349 585
R269 B.n348 B.n347 585
R270 B.n304 B.n303 585
R271 B.n496 B.n495 585
R272 B.n300 B.n299 585
R273 B.n301 B.n300 585
R274 B.n502 B.n501 585
R275 B.n501 B.n500 585
R276 B.n503 B.n298 585
R277 B.n298 B.n297 585
R278 B.n505 B.n504 585
R279 B.n506 B.n505 585
R280 B.n292 B.n291 585
R281 B.n293 B.n292 585
R282 B.n515 B.n514 585
R283 B.n514 B.n513 585
R284 B.n516 B.n290 585
R285 B.n512 B.n290 585
R286 B.n518 B.n517 585
R287 B.n519 B.n518 585
R288 B.n285 B.n284 585
R289 B.n286 B.n285 585
R290 B.n527 B.n526 585
R291 B.n526 B.n525 585
R292 B.n528 B.n283 585
R293 B.n283 B.n282 585
R294 B.n530 B.n529 585
R295 B.n531 B.n530 585
R296 B.n277 B.n276 585
R297 B.n278 B.n277 585
R298 B.n539 B.n538 585
R299 B.n538 B.n537 585
R300 B.n540 B.n275 585
R301 B.n275 B.n274 585
R302 B.n542 B.n541 585
R303 B.n543 B.n542 585
R304 B.n269 B.n268 585
R305 B.n270 B.n269 585
R306 B.n551 B.n550 585
R307 B.n550 B.n549 585
R308 B.n552 B.n267 585
R309 B.n267 B.n266 585
R310 B.n554 B.n553 585
R311 B.n555 B.n554 585
R312 B.n261 B.n260 585
R313 B.n262 B.n261 585
R314 B.n563 B.n562 585
R315 B.n562 B.n561 585
R316 B.n564 B.n259 585
R317 B.n259 B.n257 585
R318 B.n566 B.n565 585
R319 B.n567 B.n566 585
R320 B.n253 B.n252 585
R321 B.n258 B.n253 585
R322 B.n576 B.n575 585
R323 B.n575 B.n574 585
R324 B.n577 B.n251 585
R325 B.n251 B.n250 585
R326 B.n579 B.n578 585
R327 B.n580 B.n579 585
R328 B.n3 B.n0 585
R329 B.n4 B.n3 585
R330 B.n681 B.n1 585
R331 B.n682 B.n681 585
R332 B.n680 B.n679 585
R333 B.n680 B.n8 585
R334 B.n678 B.n9 585
R335 B.n12 B.n9 585
R336 B.n677 B.n676 585
R337 B.n676 B.n675 585
R338 B.n11 B.n10 585
R339 B.n674 B.n11 585
R340 B.n672 B.n671 585
R341 B.n673 B.n672 585
R342 B.n670 B.n17 585
R343 B.n17 B.n16 585
R344 B.n669 B.n668 585
R345 B.n668 B.n667 585
R346 B.n19 B.n18 585
R347 B.n666 B.n19 585
R348 B.n664 B.n663 585
R349 B.n665 B.n664 585
R350 B.n662 B.n24 585
R351 B.n24 B.n23 585
R352 B.n661 B.n660 585
R353 B.n660 B.n659 585
R354 B.n26 B.n25 585
R355 B.n658 B.n26 585
R356 B.n656 B.n655 585
R357 B.n657 B.n656 585
R358 B.n654 B.n31 585
R359 B.n31 B.n30 585
R360 B.n653 B.n652 585
R361 B.n652 B.n651 585
R362 B.n33 B.n32 585
R363 B.n650 B.n33 585
R364 B.n648 B.n647 585
R365 B.n649 B.n648 585
R366 B.n646 B.n38 585
R367 B.n38 B.n37 585
R368 B.n645 B.n644 585
R369 B.n644 B.n643 585
R370 B.n40 B.n39 585
R371 B.n642 B.n40 585
R372 B.n640 B.n639 585
R373 B.n641 B.n640 585
R374 B.n638 B.n44 585
R375 B.n47 B.n44 585
R376 B.n637 B.n636 585
R377 B.n636 B.n635 585
R378 B.n46 B.n45 585
R379 B.n634 B.n46 585
R380 B.n632 B.n631 585
R381 B.n633 B.n632 585
R382 B.n630 B.n52 585
R383 B.n52 B.n51 585
R384 B.n629 B.n628 585
R385 B.n628 B.n627 585
R386 B.n54 B.n53 585
R387 B.n626 B.n54 585
R388 B.n685 B.n684 585
R389 B.n683 B.n2 585
R390 B.n100 B.n54 554.963
R391 B.n624 B.n56 554.963
R392 B.n495 B.n302 554.963
R393 B.n491 B.n300 554.963
R394 B.n98 B.t11 309.611
R395 B.n95 B.t15 309.611
R396 B.n345 B.t8 309.611
R397 B.n342 B.t4 309.611
R398 B.n625 B.n93 256.663
R399 B.n625 B.n92 256.663
R400 B.n625 B.n91 256.663
R401 B.n625 B.n90 256.663
R402 B.n625 B.n89 256.663
R403 B.n625 B.n88 256.663
R404 B.n625 B.n87 256.663
R405 B.n625 B.n86 256.663
R406 B.n625 B.n85 256.663
R407 B.n625 B.n84 256.663
R408 B.n625 B.n83 256.663
R409 B.n625 B.n82 256.663
R410 B.n625 B.n81 256.663
R411 B.n625 B.n80 256.663
R412 B.n625 B.n79 256.663
R413 B.n625 B.n78 256.663
R414 B.n625 B.n77 256.663
R415 B.n625 B.n76 256.663
R416 B.n625 B.n75 256.663
R417 B.n625 B.n74 256.663
R418 B.n625 B.n73 256.663
R419 B.n625 B.n72 256.663
R420 B.n625 B.n71 256.663
R421 B.n625 B.n70 256.663
R422 B.n625 B.n69 256.663
R423 B.n625 B.n68 256.663
R424 B.n625 B.n67 256.663
R425 B.n625 B.n66 256.663
R426 B.n625 B.n65 256.663
R427 B.n625 B.n64 256.663
R428 B.n625 B.n63 256.663
R429 B.n625 B.n62 256.663
R430 B.n625 B.n61 256.663
R431 B.n625 B.n60 256.663
R432 B.n625 B.n59 256.663
R433 B.n625 B.n58 256.663
R434 B.n625 B.n57 256.663
R435 B.n493 B.n492 256.663
R436 B.n493 B.n305 256.663
R437 B.n493 B.n306 256.663
R438 B.n493 B.n307 256.663
R439 B.n493 B.n308 256.663
R440 B.n493 B.n309 256.663
R441 B.n493 B.n310 256.663
R442 B.n493 B.n311 256.663
R443 B.n493 B.n312 256.663
R444 B.n493 B.n313 256.663
R445 B.n493 B.n314 256.663
R446 B.n493 B.n315 256.663
R447 B.n493 B.n316 256.663
R448 B.n493 B.n317 256.663
R449 B.n493 B.n318 256.663
R450 B.n493 B.n319 256.663
R451 B.n493 B.n320 256.663
R452 B.n493 B.n321 256.663
R453 B.n493 B.n322 256.663
R454 B.n493 B.n323 256.663
R455 B.n493 B.n324 256.663
R456 B.n493 B.n325 256.663
R457 B.n493 B.n326 256.663
R458 B.n493 B.n327 256.663
R459 B.n493 B.n328 256.663
R460 B.n493 B.n329 256.663
R461 B.n493 B.n330 256.663
R462 B.n493 B.n331 256.663
R463 B.n493 B.n332 256.663
R464 B.n493 B.n333 256.663
R465 B.n493 B.n334 256.663
R466 B.n493 B.n335 256.663
R467 B.n493 B.n336 256.663
R468 B.n493 B.n337 256.663
R469 B.n493 B.n338 256.663
R470 B.n493 B.n339 256.663
R471 B.n494 B.n493 256.663
R472 B.n687 B.n686 256.663
R473 B.n104 B.n103 163.367
R474 B.n108 B.n107 163.367
R475 B.n112 B.n111 163.367
R476 B.n116 B.n115 163.367
R477 B.n120 B.n119 163.367
R478 B.n124 B.n123 163.367
R479 B.n128 B.n127 163.367
R480 B.n132 B.n131 163.367
R481 B.n136 B.n135 163.367
R482 B.n140 B.n139 163.367
R483 B.n144 B.n143 163.367
R484 B.n148 B.n147 163.367
R485 B.n152 B.n151 163.367
R486 B.n156 B.n155 163.367
R487 B.n160 B.n159 163.367
R488 B.n164 B.n163 163.367
R489 B.n169 B.n168 163.367
R490 B.n173 B.n172 163.367
R491 B.n177 B.n176 163.367
R492 B.n181 B.n180 163.367
R493 B.n185 B.n184 163.367
R494 B.n189 B.n188 163.367
R495 B.n193 B.n192 163.367
R496 B.n197 B.n196 163.367
R497 B.n201 B.n200 163.367
R498 B.n205 B.n204 163.367
R499 B.n209 B.n208 163.367
R500 B.n213 B.n212 163.367
R501 B.n217 B.n216 163.367
R502 B.n221 B.n220 163.367
R503 B.n225 B.n224 163.367
R504 B.n229 B.n228 163.367
R505 B.n233 B.n232 163.367
R506 B.n237 B.n236 163.367
R507 B.n241 B.n240 163.367
R508 B.n245 B.n244 163.367
R509 B.n624 B.n94 163.367
R510 B.n499 B.n302 163.367
R511 B.n499 B.n296 163.367
R512 B.n507 B.n296 163.367
R513 B.n507 B.n294 163.367
R514 B.n511 B.n294 163.367
R515 B.n511 B.n289 163.367
R516 B.n520 B.n289 163.367
R517 B.n520 B.n287 163.367
R518 B.n524 B.n287 163.367
R519 B.n524 B.n281 163.367
R520 B.n532 B.n281 163.367
R521 B.n532 B.n279 163.367
R522 B.n536 B.n279 163.367
R523 B.n536 B.n273 163.367
R524 B.n544 B.n273 163.367
R525 B.n544 B.n271 163.367
R526 B.n548 B.n271 163.367
R527 B.n548 B.n265 163.367
R528 B.n556 B.n265 163.367
R529 B.n556 B.n263 163.367
R530 B.n560 B.n263 163.367
R531 B.n560 B.n256 163.367
R532 B.n568 B.n256 163.367
R533 B.n568 B.n254 163.367
R534 B.n573 B.n254 163.367
R535 B.n573 B.n249 163.367
R536 B.n581 B.n249 163.367
R537 B.n582 B.n581 163.367
R538 B.n582 B.n5 163.367
R539 B.n6 B.n5 163.367
R540 B.n7 B.n6 163.367
R541 B.n588 B.n7 163.367
R542 B.n589 B.n588 163.367
R543 B.n589 B.n13 163.367
R544 B.n14 B.n13 163.367
R545 B.n15 B.n14 163.367
R546 B.n594 B.n15 163.367
R547 B.n594 B.n20 163.367
R548 B.n21 B.n20 163.367
R549 B.n22 B.n21 163.367
R550 B.n599 B.n22 163.367
R551 B.n599 B.n27 163.367
R552 B.n28 B.n27 163.367
R553 B.n29 B.n28 163.367
R554 B.n604 B.n29 163.367
R555 B.n604 B.n34 163.367
R556 B.n35 B.n34 163.367
R557 B.n36 B.n35 163.367
R558 B.n609 B.n36 163.367
R559 B.n609 B.n41 163.367
R560 B.n42 B.n41 163.367
R561 B.n43 B.n42 163.367
R562 B.n614 B.n43 163.367
R563 B.n614 B.n48 163.367
R564 B.n49 B.n48 163.367
R565 B.n50 B.n49 163.367
R566 B.n619 B.n50 163.367
R567 B.n619 B.n55 163.367
R568 B.n56 B.n55 163.367
R569 B.n341 B.n340 163.367
R570 B.n486 B.n340 163.367
R571 B.n484 B.n483 163.367
R572 B.n480 B.n479 163.367
R573 B.n476 B.n475 163.367
R574 B.n472 B.n471 163.367
R575 B.n468 B.n467 163.367
R576 B.n464 B.n463 163.367
R577 B.n460 B.n459 163.367
R578 B.n456 B.n455 163.367
R579 B.n452 B.n451 163.367
R580 B.n448 B.n447 163.367
R581 B.n444 B.n443 163.367
R582 B.n440 B.n439 163.367
R583 B.n436 B.n435 163.367
R584 B.n432 B.n431 163.367
R585 B.n428 B.n427 163.367
R586 B.n424 B.n423 163.367
R587 B.n420 B.n419 163.367
R588 B.n416 B.n415 163.367
R589 B.n412 B.n411 163.367
R590 B.n407 B.n406 163.367
R591 B.n403 B.n402 163.367
R592 B.n399 B.n398 163.367
R593 B.n395 B.n394 163.367
R594 B.n391 B.n390 163.367
R595 B.n387 B.n386 163.367
R596 B.n383 B.n382 163.367
R597 B.n379 B.n378 163.367
R598 B.n375 B.n374 163.367
R599 B.n371 B.n370 163.367
R600 B.n367 B.n366 163.367
R601 B.n363 B.n362 163.367
R602 B.n359 B.n358 163.367
R603 B.n355 B.n354 163.367
R604 B.n351 B.n350 163.367
R605 B.n347 B.n304 163.367
R606 B.n501 B.n300 163.367
R607 B.n501 B.n298 163.367
R608 B.n505 B.n298 163.367
R609 B.n505 B.n292 163.367
R610 B.n514 B.n292 163.367
R611 B.n514 B.n290 163.367
R612 B.n518 B.n290 163.367
R613 B.n518 B.n285 163.367
R614 B.n526 B.n285 163.367
R615 B.n526 B.n283 163.367
R616 B.n530 B.n283 163.367
R617 B.n530 B.n277 163.367
R618 B.n538 B.n277 163.367
R619 B.n538 B.n275 163.367
R620 B.n542 B.n275 163.367
R621 B.n542 B.n269 163.367
R622 B.n550 B.n269 163.367
R623 B.n550 B.n267 163.367
R624 B.n554 B.n267 163.367
R625 B.n554 B.n261 163.367
R626 B.n562 B.n261 163.367
R627 B.n562 B.n259 163.367
R628 B.n566 B.n259 163.367
R629 B.n566 B.n253 163.367
R630 B.n575 B.n253 163.367
R631 B.n575 B.n251 163.367
R632 B.n579 B.n251 163.367
R633 B.n579 B.n3 163.367
R634 B.n685 B.n3 163.367
R635 B.n681 B.n2 163.367
R636 B.n681 B.n680 163.367
R637 B.n680 B.n9 163.367
R638 B.n676 B.n9 163.367
R639 B.n676 B.n11 163.367
R640 B.n672 B.n11 163.367
R641 B.n672 B.n17 163.367
R642 B.n668 B.n17 163.367
R643 B.n668 B.n19 163.367
R644 B.n664 B.n19 163.367
R645 B.n664 B.n24 163.367
R646 B.n660 B.n24 163.367
R647 B.n660 B.n26 163.367
R648 B.n656 B.n26 163.367
R649 B.n656 B.n31 163.367
R650 B.n652 B.n31 163.367
R651 B.n652 B.n33 163.367
R652 B.n648 B.n33 163.367
R653 B.n648 B.n38 163.367
R654 B.n644 B.n38 163.367
R655 B.n644 B.n40 163.367
R656 B.n640 B.n40 163.367
R657 B.n640 B.n44 163.367
R658 B.n636 B.n44 163.367
R659 B.n636 B.n46 163.367
R660 B.n632 B.n46 163.367
R661 B.n632 B.n52 163.367
R662 B.n628 B.n52 163.367
R663 B.n628 B.n54 163.367
R664 B.n95 B.t16 119.145
R665 B.n345 B.t10 119.145
R666 B.n98 B.t13 119.135
R667 B.n342 B.t7 119.135
R668 B.n493 B.n301 107.035
R669 B.n626 B.n625 107.035
R670 B.n100 B.n57 71.676
R671 B.n104 B.n58 71.676
R672 B.n108 B.n59 71.676
R673 B.n112 B.n60 71.676
R674 B.n116 B.n61 71.676
R675 B.n120 B.n62 71.676
R676 B.n124 B.n63 71.676
R677 B.n128 B.n64 71.676
R678 B.n132 B.n65 71.676
R679 B.n136 B.n66 71.676
R680 B.n140 B.n67 71.676
R681 B.n144 B.n68 71.676
R682 B.n148 B.n69 71.676
R683 B.n152 B.n70 71.676
R684 B.n156 B.n71 71.676
R685 B.n160 B.n72 71.676
R686 B.n164 B.n73 71.676
R687 B.n169 B.n74 71.676
R688 B.n173 B.n75 71.676
R689 B.n177 B.n76 71.676
R690 B.n181 B.n77 71.676
R691 B.n185 B.n78 71.676
R692 B.n189 B.n79 71.676
R693 B.n193 B.n80 71.676
R694 B.n197 B.n81 71.676
R695 B.n201 B.n82 71.676
R696 B.n205 B.n83 71.676
R697 B.n209 B.n84 71.676
R698 B.n213 B.n85 71.676
R699 B.n217 B.n86 71.676
R700 B.n221 B.n87 71.676
R701 B.n225 B.n88 71.676
R702 B.n229 B.n89 71.676
R703 B.n233 B.n90 71.676
R704 B.n237 B.n91 71.676
R705 B.n241 B.n92 71.676
R706 B.n245 B.n93 71.676
R707 B.n94 B.n93 71.676
R708 B.n244 B.n92 71.676
R709 B.n240 B.n91 71.676
R710 B.n236 B.n90 71.676
R711 B.n232 B.n89 71.676
R712 B.n228 B.n88 71.676
R713 B.n224 B.n87 71.676
R714 B.n220 B.n86 71.676
R715 B.n216 B.n85 71.676
R716 B.n212 B.n84 71.676
R717 B.n208 B.n83 71.676
R718 B.n204 B.n82 71.676
R719 B.n200 B.n81 71.676
R720 B.n196 B.n80 71.676
R721 B.n192 B.n79 71.676
R722 B.n188 B.n78 71.676
R723 B.n184 B.n77 71.676
R724 B.n180 B.n76 71.676
R725 B.n176 B.n75 71.676
R726 B.n172 B.n74 71.676
R727 B.n168 B.n73 71.676
R728 B.n163 B.n72 71.676
R729 B.n159 B.n71 71.676
R730 B.n155 B.n70 71.676
R731 B.n151 B.n69 71.676
R732 B.n147 B.n68 71.676
R733 B.n143 B.n67 71.676
R734 B.n139 B.n66 71.676
R735 B.n135 B.n65 71.676
R736 B.n131 B.n64 71.676
R737 B.n127 B.n63 71.676
R738 B.n123 B.n62 71.676
R739 B.n119 B.n61 71.676
R740 B.n115 B.n60 71.676
R741 B.n111 B.n59 71.676
R742 B.n107 B.n58 71.676
R743 B.n103 B.n57 71.676
R744 B.n492 B.n491 71.676
R745 B.n486 B.n305 71.676
R746 B.n483 B.n306 71.676
R747 B.n479 B.n307 71.676
R748 B.n475 B.n308 71.676
R749 B.n471 B.n309 71.676
R750 B.n467 B.n310 71.676
R751 B.n463 B.n311 71.676
R752 B.n459 B.n312 71.676
R753 B.n455 B.n313 71.676
R754 B.n451 B.n314 71.676
R755 B.n447 B.n315 71.676
R756 B.n443 B.n316 71.676
R757 B.n439 B.n317 71.676
R758 B.n435 B.n318 71.676
R759 B.n431 B.n319 71.676
R760 B.n427 B.n320 71.676
R761 B.n423 B.n321 71.676
R762 B.n419 B.n322 71.676
R763 B.n415 B.n323 71.676
R764 B.n411 B.n324 71.676
R765 B.n406 B.n325 71.676
R766 B.n402 B.n326 71.676
R767 B.n398 B.n327 71.676
R768 B.n394 B.n328 71.676
R769 B.n390 B.n329 71.676
R770 B.n386 B.n330 71.676
R771 B.n382 B.n331 71.676
R772 B.n378 B.n332 71.676
R773 B.n374 B.n333 71.676
R774 B.n370 B.n334 71.676
R775 B.n366 B.n335 71.676
R776 B.n362 B.n336 71.676
R777 B.n358 B.n337 71.676
R778 B.n354 B.n338 71.676
R779 B.n350 B.n339 71.676
R780 B.n494 B.n304 71.676
R781 B.n492 B.n341 71.676
R782 B.n484 B.n305 71.676
R783 B.n480 B.n306 71.676
R784 B.n476 B.n307 71.676
R785 B.n472 B.n308 71.676
R786 B.n468 B.n309 71.676
R787 B.n464 B.n310 71.676
R788 B.n460 B.n311 71.676
R789 B.n456 B.n312 71.676
R790 B.n452 B.n313 71.676
R791 B.n448 B.n314 71.676
R792 B.n444 B.n315 71.676
R793 B.n440 B.n316 71.676
R794 B.n436 B.n317 71.676
R795 B.n432 B.n318 71.676
R796 B.n428 B.n319 71.676
R797 B.n424 B.n320 71.676
R798 B.n420 B.n321 71.676
R799 B.n416 B.n322 71.676
R800 B.n412 B.n323 71.676
R801 B.n407 B.n324 71.676
R802 B.n403 B.n325 71.676
R803 B.n399 B.n326 71.676
R804 B.n395 B.n327 71.676
R805 B.n391 B.n328 71.676
R806 B.n387 B.n329 71.676
R807 B.n383 B.n330 71.676
R808 B.n379 B.n331 71.676
R809 B.n375 B.n332 71.676
R810 B.n371 B.n333 71.676
R811 B.n367 B.n334 71.676
R812 B.n363 B.n335 71.676
R813 B.n359 B.n336 71.676
R814 B.n355 B.n337 71.676
R815 B.n351 B.n338 71.676
R816 B.n347 B.n339 71.676
R817 B.n495 B.n494 71.676
R818 B.n686 B.n685 71.676
R819 B.n686 B.n2 71.676
R820 B.n96 B.t17 71.6301
R821 B.n346 B.t9 71.6301
R822 B.n99 B.t14 71.6194
R823 B.n343 B.t6 71.6194
R824 B.n166 B.n99 59.5399
R825 B.n97 B.n96 59.5399
R826 B.n409 B.n346 59.5399
R827 B.n344 B.n343 59.5399
R828 B.n500 B.n301 52.3631
R829 B.n500 B.n297 52.3631
R830 B.n506 B.n297 52.3631
R831 B.n506 B.n293 52.3631
R832 B.n513 B.n293 52.3631
R833 B.n513 B.n512 52.3631
R834 B.n519 B.n286 52.3631
R835 B.n525 B.n286 52.3631
R836 B.n525 B.n282 52.3631
R837 B.n531 B.n282 52.3631
R838 B.n531 B.n278 52.3631
R839 B.n537 B.n278 52.3631
R840 B.n537 B.n274 52.3631
R841 B.n543 B.n274 52.3631
R842 B.n543 B.n270 52.3631
R843 B.n549 B.n270 52.3631
R844 B.n555 B.n266 52.3631
R845 B.n555 B.n262 52.3631
R846 B.n561 B.n262 52.3631
R847 B.n561 B.n257 52.3631
R848 B.n567 B.n257 52.3631
R849 B.n567 B.n258 52.3631
R850 B.n574 B.n250 52.3631
R851 B.n580 B.n250 52.3631
R852 B.n580 B.n4 52.3631
R853 B.n684 B.n4 52.3631
R854 B.n684 B.n683 52.3631
R855 B.n683 B.n682 52.3631
R856 B.n682 B.n8 52.3631
R857 B.n12 B.n8 52.3631
R858 B.n675 B.n12 52.3631
R859 B.n674 B.n673 52.3631
R860 B.n673 B.n16 52.3631
R861 B.n667 B.n16 52.3631
R862 B.n667 B.n666 52.3631
R863 B.n666 B.n665 52.3631
R864 B.n665 B.n23 52.3631
R865 B.n659 B.n658 52.3631
R866 B.n658 B.n657 52.3631
R867 B.n657 B.n30 52.3631
R868 B.n651 B.n30 52.3631
R869 B.n651 B.n650 52.3631
R870 B.n650 B.n649 52.3631
R871 B.n649 B.n37 52.3631
R872 B.n643 B.n37 52.3631
R873 B.n643 B.n642 52.3631
R874 B.n642 B.n641 52.3631
R875 B.n635 B.n47 52.3631
R876 B.n635 B.n634 52.3631
R877 B.n634 B.n633 52.3631
R878 B.n633 B.n51 52.3631
R879 B.n627 B.n51 52.3631
R880 B.n627 B.n626 52.3631
R881 B.t0 B.n266 47.7429
R882 B.t1 B.n23 47.7429
R883 B.n99 B.n98 47.5157
R884 B.n96 B.n95 47.5157
R885 B.n346 B.n345 47.5157
R886 B.n343 B.n342 47.5157
R887 B.n574 B.t2 36.9623
R888 B.n675 B.t3 36.9623
R889 B.n623 B.n622 36.059
R890 B.n490 B.n299 36.059
R891 B.n497 B.n496 36.059
R892 B.n101 B.n53 36.059
R893 B.n512 B.t5 35.4223
R894 B.n47 B.t12 35.4223
R895 B B.n687 18.0485
R896 B.n519 B.t5 16.9413
R897 B.n641 B.t12 16.9413
R898 B.n258 B.t2 15.4013
R899 B.t3 B.n674 15.4013
R900 B.n502 B.n299 10.6151
R901 B.n503 B.n502 10.6151
R902 B.n504 B.n503 10.6151
R903 B.n504 B.n291 10.6151
R904 B.n515 B.n291 10.6151
R905 B.n516 B.n515 10.6151
R906 B.n517 B.n516 10.6151
R907 B.n517 B.n284 10.6151
R908 B.n527 B.n284 10.6151
R909 B.n528 B.n527 10.6151
R910 B.n529 B.n528 10.6151
R911 B.n529 B.n276 10.6151
R912 B.n539 B.n276 10.6151
R913 B.n540 B.n539 10.6151
R914 B.n541 B.n540 10.6151
R915 B.n541 B.n268 10.6151
R916 B.n551 B.n268 10.6151
R917 B.n552 B.n551 10.6151
R918 B.n553 B.n552 10.6151
R919 B.n553 B.n260 10.6151
R920 B.n563 B.n260 10.6151
R921 B.n564 B.n563 10.6151
R922 B.n565 B.n564 10.6151
R923 B.n565 B.n252 10.6151
R924 B.n576 B.n252 10.6151
R925 B.n577 B.n576 10.6151
R926 B.n578 B.n577 10.6151
R927 B.n578 B.n0 10.6151
R928 B.n490 B.n489 10.6151
R929 B.n489 B.n488 10.6151
R930 B.n488 B.n487 10.6151
R931 B.n487 B.n485 10.6151
R932 B.n485 B.n482 10.6151
R933 B.n482 B.n481 10.6151
R934 B.n481 B.n478 10.6151
R935 B.n478 B.n477 10.6151
R936 B.n477 B.n474 10.6151
R937 B.n474 B.n473 10.6151
R938 B.n473 B.n470 10.6151
R939 B.n470 B.n469 10.6151
R940 B.n469 B.n466 10.6151
R941 B.n466 B.n465 10.6151
R942 B.n465 B.n462 10.6151
R943 B.n462 B.n461 10.6151
R944 B.n461 B.n458 10.6151
R945 B.n458 B.n457 10.6151
R946 B.n457 B.n454 10.6151
R947 B.n454 B.n453 10.6151
R948 B.n453 B.n450 10.6151
R949 B.n450 B.n449 10.6151
R950 B.n449 B.n446 10.6151
R951 B.n446 B.n445 10.6151
R952 B.n445 B.n442 10.6151
R953 B.n442 B.n441 10.6151
R954 B.n441 B.n438 10.6151
R955 B.n438 B.n437 10.6151
R956 B.n437 B.n434 10.6151
R957 B.n434 B.n433 10.6151
R958 B.n433 B.n430 10.6151
R959 B.n430 B.n429 10.6151
R960 B.n426 B.n425 10.6151
R961 B.n425 B.n422 10.6151
R962 B.n422 B.n421 10.6151
R963 B.n421 B.n418 10.6151
R964 B.n418 B.n417 10.6151
R965 B.n417 B.n414 10.6151
R966 B.n414 B.n413 10.6151
R967 B.n413 B.n410 10.6151
R968 B.n408 B.n405 10.6151
R969 B.n405 B.n404 10.6151
R970 B.n404 B.n401 10.6151
R971 B.n401 B.n400 10.6151
R972 B.n400 B.n397 10.6151
R973 B.n397 B.n396 10.6151
R974 B.n396 B.n393 10.6151
R975 B.n393 B.n392 10.6151
R976 B.n392 B.n389 10.6151
R977 B.n389 B.n388 10.6151
R978 B.n388 B.n385 10.6151
R979 B.n385 B.n384 10.6151
R980 B.n384 B.n381 10.6151
R981 B.n381 B.n380 10.6151
R982 B.n380 B.n377 10.6151
R983 B.n377 B.n376 10.6151
R984 B.n376 B.n373 10.6151
R985 B.n373 B.n372 10.6151
R986 B.n372 B.n369 10.6151
R987 B.n369 B.n368 10.6151
R988 B.n368 B.n365 10.6151
R989 B.n365 B.n364 10.6151
R990 B.n364 B.n361 10.6151
R991 B.n361 B.n360 10.6151
R992 B.n360 B.n357 10.6151
R993 B.n357 B.n356 10.6151
R994 B.n356 B.n353 10.6151
R995 B.n353 B.n352 10.6151
R996 B.n352 B.n349 10.6151
R997 B.n349 B.n348 10.6151
R998 B.n348 B.n303 10.6151
R999 B.n496 B.n303 10.6151
R1000 B.n498 B.n497 10.6151
R1001 B.n498 B.n295 10.6151
R1002 B.n508 B.n295 10.6151
R1003 B.n509 B.n508 10.6151
R1004 B.n510 B.n509 10.6151
R1005 B.n510 B.n288 10.6151
R1006 B.n521 B.n288 10.6151
R1007 B.n522 B.n521 10.6151
R1008 B.n523 B.n522 10.6151
R1009 B.n523 B.n280 10.6151
R1010 B.n533 B.n280 10.6151
R1011 B.n534 B.n533 10.6151
R1012 B.n535 B.n534 10.6151
R1013 B.n535 B.n272 10.6151
R1014 B.n545 B.n272 10.6151
R1015 B.n546 B.n545 10.6151
R1016 B.n547 B.n546 10.6151
R1017 B.n547 B.n264 10.6151
R1018 B.n557 B.n264 10.6151
R1019 B.n558 B.n557 10.6151
R1020 B.n559 B.n558 10.6151
R1021 B.n559 B.n255 10.6151
R1022 B.n569 B.n255 10.6151
R1023 B.n570 B.n569 10.6151
R1024 B.n572 B.n570 10.6151
R1025 B.n572 B.n571 10.6151
R1026 B.n571 B.n248 10.6151
R1027 B.n583 B.n248 10.6151
R1028 B.n584 B.n583 10.6151
R1029 B.n585 B.n584 10.6151
R1030 B.n586 B.n585 10.6151
R1031 B.n587 B.n586 10.6151
R1032 B.n590 B.n587 10.6151
R1033 B.n591 B.n590 10.6151
R1034 B.n592 B.n591 10.6151
R1035 B.n593 B.n592 10.6151
R1036 B.n595 B.n593 10.6151
R1037 B.n596 B.n595 10.6151
R1038 B.n597 B.n596 10.6151
R1039 B.n598 B.n597 10.6151
R1040 B.n600 B.n598 10.6151
R1041 B.n601 B.n600 10.6151
R1042 B.n602 B.n601 10.6151
R1043 B.n603 B.n602 10.6151
R1044 B.n605 B.n603 10.6151
R1045 B.n606 B.n605 10.6151
R1046 B.n607 B.n606 10.6151
R1047 B.n608 B.n607 10.6151
R1048 B.n610 B.n608 10.6151
R1049 B.n611 B.n610 10.6151
R1050 B.n612 B.n611 10.6151
R1051 B.n613 B.n612 10.6151
R1052 B.n615 B.n613 10.6151
R1053 B.n616 B.n615 10.6151
R1054 B.n617 B.n616 10.6151
R1055 B.n618 B.n617 10.6151
R1056 B.n620 B.n618 10.6151
R1057 B.n621 B.n620 10.6151
R1058 B.n622 B.n621 10.6151
R1059 B.n679 B.n1 10.6151
R1060 B.n679 B.n678 10.6151
R1061 B.n678 B.n677 10.6151
R1062 B.n677 B.n10 10.6151
R1063 B.n671 B.n10 10.6151
R1064 B.n671 B.n670 10.6151
R1065 B.n670 B.n669 10.6151
R1066 B.n669 B.n18 10.6151
R1067 B.n663 B.n18 10.6151
R1068 B.n663 B.n662 10.6151
R1069 B.n662 B.n661 10.6151
R1070 B.n661 B.n25 10.6151
R1071 B.n655 B.n25 10.6151
R1072 B.n655 B.n654 10.6151
R1073 B.n654 B.n653 10.6151
R1074 B.n653 B.n32 10.6151
R1075 B.n647 B.n32 10.6151
R1076 B.n647 B.n646 10.6151
R1077 B.n646 B.n645 10.6151
R1078 B.n645 B.n39 10.6151
R1079 B.n639 B.n39 10.6151
R1080 B.n639 B.n638 10.6151
R1081 B.n638 B.n637 10.6151
R1082 B.n637 B.n45 10.6151
R1083 B.n631 B.n45 10.6151
R1084 B.n631 B.n630 10.6151
R1085 B.n630 B.n629 10.6151
R1086 B.n629 B.n53 10.6151
R1087 B.n102 B.n101 10.6151
R1088 B.n105 B.n102 10.6151
R1089 B.n106 B.n105 10.6151
R1090 B.n109 B.n106 10.6151
R1091 B.n110 B.n109 10.6151
R1092 B.n113 B.n110 10.6151
R1093 B.n114 B.n113 10.6151
R1094 B.n117 B.n114 10.6151
R1095 B.n118 B.n117 10.6151
R1096 B.n121 B.n118 10.6151
R1097 B.n122 B.n121 10.6151
R1098 B.n125 B.n122 10.6151
R1099 B.n126 B.n125 10.6151
R1100 B.n129 B.n126 10.6151
R1101 B.n130 B.n129 10.6151
R1102 B.n133 B.n130 10.6151
R1103 B.n134 B.n133 10.6151
R1104 B.n137 B.n134 10.6151
R1105 B.n138 B.n137 10.6151
R1106 B.n141 B.n138 10.6151
R1107 B.n142 B.n141 10.6151
R1108 B.n145 B.n142 10.6151
R1109 B.n146 B.n145 10.6151
R1110 B.n149 B.n146 10.6151
R1111 B.n150 B.n149 10.6151
R1112 B.n153 B.n150 10.6151
R1113 B.n154 B.n153 10.6151
R1114 B.n157 B.n154 10.6151
R1115 B.n158 B.n157 10.6151
R1116 B.n161 B.n158 10.6151
R1117 B.n162 B.n161 10.6151
R1118 B.n165 B.n162 10.6151
R1119 B.n170 B.n167 10.6151
R1120 B.n171 B.n170 10.6151
R1121 B.n174 B.n171 10.6151
R1122 B.n175 B.n174 10.6151
R1123 B.n178 B.n175 10.6151
R1124 B.n179 B.n178 10.6151
R1125 B.n182 B.n179 10.6151
R1126 B.n183 B.n182 10.6151
R1127 B.n187 B.n186 10.6151
R1128 B.n190 B.n187 10.6151
R1129 B.n191 B.n190 10.6151
R1130 B.n194 B.n191 10.6151
R1131 B.n195 B.n194 10.6151
R1132 B.n198 B.n195 10.6151
R1133 B.n199 B.n198 10.6151
R1134 B.n202 B.n199 10.6151
R1135 B.n203 B.n202 10.6151
R1136 B.n206 B.n203 10.6151
R1137 B.n207 B.n206 10.6151
R1138 B.n210 B.n207 10.6151
R1139 B.n211 B.n210 10.6151
R1140 B.n214 B.n211 10.6151
R1141 B.n215 B.n214 10.6151
R1142 B.n218 B.n215 10.6151
R1143 B.n219 B.n218 10.6151
R1144 B.n222 B.n219 10.6151
R1145 B.n223 B.n222 10.6151
R1146 B.n226 B.n223 10.6151
R1147 B.n227 B.n226 10.6151
R1148 B.n230 B.n227 10.6151
R1149 B.n231 B.n230 10.6151
R1150 B.n234 B.n231 10.6151
R1151 B.n235 B.n234 10.6151
R1152 B.n238 B.n235 10.6151
R1153 B.n239 B.n238 10.6151
R1154 B.n242 B.n239 10.6151
R1155 B.n243 B.n242 10.6151
R1156 B.n246 B.n243 10.6151
R1157 B.n247 B.n246 10.6151
R1158 B.n623 B.n247 10.6151
R1159 B.n687 B.n0 8.11757
R1160 B.n687 B.n1 8.11757
R1161 B.n426 B.n344 6.5566
R1162 B.n410 B.n409 6.5566
R1163 B.n167 B.n166 6.5566
R1164 B.n183 B.n97 6.5566
R1165 B.n549 B.t0 4.62073
R1166 B.n659 B.t1 4.62073
R1167 B.n429 B.n344 4.05904
R1168 B.n409 B.n408 4.05904
R1169 B.n166 B.n165 4.05904
R1170 B.n186 B.n97 4.05904
R1171 VP.n10 VP.n0 161.3
R1172 VP.n9 VP.n8 161.3
R1173 VP.n7 VP.n1 161.3
R1174 VP.n6 VP.n5 161.3
R1175 VP.n2 VP.t3 138.625
R1176 VP.n2 VP.t1 138.075
R1177 VP.n4 VP.t0 102.425
R1178 VP.n11 VP.t2 102.425
R1179 VP.n4 VP.n3 87.5128
R1180 VP.n12 VP.n11 87.5128
R1181 VP.n9 VP.n1 56.5193
R1182 VP.n3 VP.n2 49.4585
R1183 VP.n5 VP.n1 24.4675
R1184 VP.n10 VP.n9 24.4675
R1185 VP.n5 VP.n4 23.2442
R1186 VP.n11 VP.n10 23.2442
R1187 VP.n6 VP.n3 0.278367
R1188 VP.n12 VP.n0 0.278367
R1189 VP.n7 VP.n6 0.189894
R1190 VP.n8 VP.n7 0.189894
R1191 VP.n8 VP.n0 0.189894
R1192 VP VP.n12 0.153454
R1193 VDD1 VDD1.n1 104.075
R1194 VDD1 VDD1.n0 65.7896
R1195 VDD1.n0 VDD1.t3 2.19806
R1196 VDD1.n0 VDD1.t0 2.19806
R1197 VDD1.n1 VDD1.t1 2.19806
R1198 VDD1.n1 VDD1.t2 2.19806
R1199 VTAIL.n5 VTAIL.t4 51.2503
R1200 VTAIL.n4 VTAIL.t2 51.2503
R1201 VTAIL.n3 VTAIL.t0 51.2503
R1202 VTAIL.n7 VTAIL.t1 51.25
R1203 VTAIL.n0 VTAIL.t3 51.25
R1204 VTAIL.n1 VTAIL.t5 51.25
R1205 VTAIL.n2 VTAIL.t7 51.25
R1206 VTAIL.n6 VTAIL.t6 51.25
R1207 VTAIL.n7 VTAIL.n6 22.2462
R1208 VTAIL.n3 VTAIL.n2 22.2462
R1209 VTAIL.n4 VTAIL.n3 2.11257
R1210 VTAIL.n6 VTAIL.n5 2.11257
R1211 VTAIL.n2 VTAIL.n1 2.11257
R1212 VTAIL VTAIL.n0 1.11472
R1213 VTAIL VTAIL.n7 0.998345
R1214 VTAIL.n5 VTAIL.n4 0.470328
R1215 VTAIL.n1 VTAIL.n0 0.470328
R1216 VN.n0 VN.t3 138.625
R1217 VN.n1 VN.t2 138.625
R1218 VN.n0 VN.t1 138.075
R1219 VN.n1 VN.t0 138.075
R1220 VN VN.n1 49.7374
R1221 VN VN.n0 6.83209
R1222 VDD2.n2 VDD2.n0 103.549
R1223 VDD2.n2 VDD2.n1 65.7314
R1224 VDD2.n1 VDD2.t3 2.19806
R1225 VDD2.n1 VDD2.t1 2.19806
R1226 VDD2.n0 VDD2.t0 2.19806
R1227 VDD2.n0 VDD2.t2 2.19806
R1228 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 4.60138f
C1 VDD1 VP 3.71388f
C2 VN VDD1 0.148694f
C3 VDD2 VTAIL 4.65236f
C4 VDD2 VP 0.36389f
C5 VTAIL VP 3.48817f
C6 VN VDD2 3.4993f
C7 VN VTAIL 3.47407f
C8 VN VP 5.28871f
C9 VDD2 VDD1 0.913864f
C10 VDD2 B 3.263415f
C11 VDD1 B 6.92305f
C12 VTAIL B 8.016685f
C13 VN B 9.55246f
C14 VP B 7.713583f
C15 VDD2.t0 B 0.19281f
C16 VDD2.t2 B 0.19281f
C17 VDD2.n0 B 2.21641f
C18 VDD2.t3 B 0.19281f
C19 VDD2.t1 B 0.19281f
C20 VDD2.n1 B 1.68672f
C21 VDD2.n2 B 3.3355f
C22 VN.t3 B 1.73224f
C23 VN.t1 B 1.72939f
C24 VN.n0 B 1.15954f
C25 VN.t2 B 1.73224f
C26 VN.t0 B 1.72939f
C27 VN.n1 B 2.46757f
C28 VTAIL.t3 B 1.30477f
C29 VTAIL.n0 B 0.300454f
C30 VTAIL.t5 B 1.30477f
C31 VTAIL.n1 B 0.355681f
C32 VTAIL.t7 B 1.30477f
C33 VTAIL.n2 B 1.10978f
C34 VTAIL.t0 B 1.30477f
C35 VTAIL.n3 B 1.10978f
C36 VTAIL.t2 B 1.30477f
C37 VTAIL.n4 B 0.355678f
C38 VTAIL.t4 B 1.30477f
C39 VTAIL.n5 B 0.355678f
C40 VTAIL.t6 B 1.30477f
C41 VTAIL.n6 B 1.10978f
C42 VTAIL.t1 B 1.30477f
C43 VTAIL.n7 B 1.04811f
C44 VDD1.t3 B 0.19281f
C45 VDD1.t0 B 0.19281f
C46 VDD1.n0 B 1.68709f
C47 VDD1.t1 B 0.19281f
C48 VDD1.t2 B 0.19281f
C49 VDD1.n1 B 2.24111f
C50 VP.n0 B 0.040199f
C51 VP.t2 B 1.57179f
C52 VP.n1 B 0.044511f
C53 VP.t1 B 1.76354f
C54 VP.t3 B 1.76644f
C55 VP.n2 B 2.50057f
C56 VP.n3 B 1.55363f
C57 VP.t0 B 1.57179f
C58 VP.n4 B 0.677898f
C59 VP.n5 B 0.055423f
C60 VP.n6 B 0.040199f
C61 VP.n7 B 0.030491f
C62 VP.n8 B 0.030491f
C63 VP.n9 B 0.044511f
C64 VP.n10 B 0.055423f
C65 VP.n11 B 0.677898f
C66 VP.n12 B 0.034093f
.ends

