* NGSPICE file created from diff_pair_sample_0436.ext - technology: sky130A

.subckt diff_pair_sample_0436 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=2.47
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=2.47
X2 VTAIL.t7 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=2.47
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=2.47
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=2.47
X5 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=2.47
X6 VTAIL.t2 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=2.47
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=2.47
X8 VDD1.t1 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=2.47
X9 VTAIL.t1 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=2.47
X10 VDD1.t0 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=2.47
X11 VTAIL.t4 VP.t3 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=2.47
R0 B.n937 B.n936 585
R1 B.n395 B.n128 585
R2 B.n394 B.n393 585
R3 B.n392 B.n391 585
R4 B.n390 B.n389 585
R5 B.n388 B.n387 585
R6 B.n386 B.n385 585
R7 B.n384 B.n383 585
R8 B.n382 B.n381 585
R9 B.n380 B.n379 585
R10 B.n378 B.n377 585
R11 B.n376 B.n375 585
R12 B.n374 B.n373 585
R13 B.n372 B.n371 585
R14 B.n370 B.n369 585
R15 B.n368 B.n367 585
R16 B.n366 B.n365 585
R17 B.n364 B.n363 585
R18 B.n362 B.n361 585
R19 B.n360 B.n359 585
R20 B.n358 B.n357 585
R21 B.n356 B.n355 585
R22 B.n354 B.n353 585
R23 B.n352 B.n351 585
R24 B.n350 B.n349 585
R25 B.n348 B.n347 585
R26 B.n346 B.n345 585
R27 B.n344 B.n343 585
R28 B.n342 B.n341 585
R29 B.n340 B.n339 585
R30 B.n338 B.n337 585
R31 B.n336 B.n335 585
R32 B.n334 B.n333 585
R33 B.n332 B.n331 585
R34 B.n330 B.n329 585
R35 B.n328 B.n327 585
R36 B.n326 B.n325 585
R37 B.n324 B.n323 585
R38 B.n322 B.n321 585
R39 B.n320 B.n319 585
R40 B.n318 B.n317 585
R41 B.n316 B.n315 585
R42 B.n314 B.n313 585
R43 B.n312 B.n311 585
R44 B.n310 B.n309 585
R45 B.n308 B.n307 585
R46 B.n306 B.n305 585
R47 B.n304 B.n303 585
R48 B.n302 B.n301 585
R49 B.n300 B.n299 585
R50 B.n298 B.n297 585
R51 B.n296 B.n295 585
R52 B.n294 B.n293 585
R53 B.n292 B.n291 585
R54 B.n290 B.n289 585
R55 B.n288 B.n287 585
R56 B.n286 B.n285 585
R57 B.n284 B.n283 585
R58 B.n282 B.n281 585
R59 B.n280 B.n279 585
R60 B.n278 B.n277 585
R61 B.n275 B.n274 585
R62 B.n273 B.n272 585
R63 B.n271 B.n270 585
R64 B.n269 B.n268 585
R65 B.n267 B.n266 585
R66 B.n265 B.n264 585
R67 B.n263 B.n262 585
R68 B.n261 B.n260 585
R69 B.n259 B.n258 585
R70 B.n257 B.n256 585
R71 B.n254 B.n253 585
R72 B.n252 B.n251 585
R73 B.n250 B.n249 585
R74 B.n248 B.n247 585
R75 B.n246 B.n245 585
R76 B.n244 B.n243 585
R77 B.n242 B.n241 585
R78 B.n240 B.n239 585
R79 B.n238 B.n237 585
R80 B.n236 B.n235 585
R81 B.n234 B.n233 585
R82 B.n232 B.n231 585
R83 B.n230 B.n229 585
R84 B.n228 B.n227 585
R85 B.n226 B.n225 585
R86 B.n224 B.n223 585
R87 B.n222 B.n221 585
R88 B.n220 B.n219 585
R89 B.n218 B.n217 585
R90 B.n216 B.n215 585
R91 B.n214 B.n213 585
R92 B.n212 B.n211 585
R93 B.n210 B.n209 585
R94 B.n208 B.n207 585
R95 B.n206 B.n205 585
R96 B.n204 B.n203 585
R97 B.n202 B.n201 585
R98 B.n200 B.n199 585
R99 B.n198 B.n197 585
R100 B.n196 B.n195 585
R101 B.n194 B.n193 585
R102 B.n192 B.n191 585
R103 B.n190 B.n189 585
R104 B.n188 B.n187 585
R105 B.n186 B.n185 585
R106 B.n184 B.n183 585
R107 B.n182 B.n181 585
R108 B.n180 B.n179 585
R109 B.n178 B.n177 585
R110 B.n176 B.n175 585
R111 B.n174 B.n173 585
R112 B.n172 B.n171 585
R113 B.n170 B.n169 585
R114 B.n168 B.n167 585
R115 B.n166 B.n165 585
R116 B.n164 B.n163 585
R117 B.n162 B.n161 585
R118 B.n160 B.n159 585
R119 B.n158 B.n157 585
R120 B.n156 B.n155 585
R121 B.n154 B.n153 585
R122 B.n152 B.n151 585
R123 B.n150 B.n149 585
R124 B.n148 B.n147 585
R125 B.n146 B.n145 585
R126 B.n144 B.n143 585
R127 B.n142 B.n141 585
R128 B.n140 B.n139 585
R129 B.n138 B.n137 585
R130 B.n136 B.n135 585
R131 B.n134 B.n133 585
R132 B.n935 B.n62 585
R133 B.n940 B.n62 585
R134 B.n934 B.n61 585
R135 B.n941 B.n61 585
R136 B.n933 B.n932 585
R137 B.n932 B.n57 585
R138 B.n931 B.n56 585
R139 B.n947 B.n56 585
R140 B.n930 B.n55 585
R141 B.n948 B.n55 585
R142 B.n929 B.n54 585
R143 B.n949 B.n54 585
R144 B.n928 B.n927 585
R145 B.n927 B.n50 585
R146 B.n926 B.n49 585
R147 B.n955 B.n49 585
R148 B.n925 B.n48 585
R149 B.n956 B.n48 585
R150 B.n924 B.n47 585
R151 B.n957 B.n47 585
R152 B.n923 B.n922 585
R153 B.n922 B.n43 585
R154 B.n921 B.n42 585
R155 B.n963 B.n42 585
R156 B.n920 B.n41 585
R157 B.n964 B.n41 585
R158 B.n919 B.n40 585
R159 B.n965 B.n40 585
R160 B.n918 B.n917 585
R161 B.n917 B.n36 585
R162 B.n916 B.n35 585
R163 B.n971 B.n35 585
R164 B.n915 B.n34 585
R165 B.n972 B.n34 585
R166 B.n914 B.n33 585
R167 B.n973 B.n33 585
R168 B.n913 B.n912 585
R169 B.n912 B.n29 585
R170 B.n911 B.n28 585
R171 B.n979 B.n28 585
R172 B.n910 B.n27 585
R173 B.n980 B.n27 585
R174 B.n909 B.n26 585
R175 B.n981 B.n26 585
R176 B.n908 B.n907 585
R177 B.n907 B.n22 585
R178 B.n906 B.n21 585
R179 B.n987 B.n21 585
R180 B.n905 B.n20 585
R181 B.n988 B.n20 585
R182 B.n904 B.n19 585
R183 B.n989 B.n19 585
R184 B.n903 B.n902 585
R185 B.n902 B.n15 585
R186 B.n901 B.n14 585
R187 B.n995 B.n14 585
R188 B.n900 B.n13 585
R189 B.n996 B.n13 585
R190 B.n899 B.n12 585
R191 B.n997 B.n12 585
R192 B.n898 B.n897 585
R193 B.n897 B.n8 585
R194 B.n896 B.n7 585
R195 B.n1003 B.n7 585
R196 B.n895 B.n6 585
R197 B.n1004 B.n6 585
R198 B.n894 B.n5 585
R199 B.n1005 B.n5 585
R200 B.n893 B.n892 585
R201 B.n892 B.n4 585
R202 B.n891 B.n396 585
R203 B.n891 B.n890 585
R204 B.n881 B.n397 585
R205 B.n398 B.n397 585
R206 B.n883 B.n882 585
R207 B.n884 B.n883 585
R208 B.n880 B.n403 585
R209 B.n403 B.n402 585
R210 B.n879 B.n878 585
R211 B.n878 B.n877 585
R212 B.n405 B.n404 585
R213 B.n406 B.n405 585
R214 B.n870 B.n869 585
R215 B.n871 B.n870 585
R216 B.n868 B.n411 585
R217 B.n411 B.n410 585
R218 B.n867 B.n866 585
R219 B.n866 B.n865 585
R220 B.n413 B.n412 585
R221 B.n414 B.n413 585
R222 B.n858 B.n857 585
R223 B.n859 B.n858 585
R224 B.n856 B.n419 585
R225 B.n419 B.n418 585
R226 B.n855 B.n854 585
R227 B.n854 B.n853 585
R228 B.n421 B.n420 585
R229 B.n422 B.n421 585
R230 B.n846 B.n845 585
R231 B.n847 B.n846 585
R232 B.n844 B.n427 585
R233 B.n427 B.n426 585
R234 B.n843 B.n842 585
R235 B.n842 B.n841 585
R236 B.n429 B.n428 585
R237 B.n430 B.n429 585
R238 B.n834 B.n833 585
R239 B.n835 B.n834 585
R240 B.n832 B.n435 585
R241 B.n435 B.n434 585
R242 B.n831 B.n830 585
R243 B.n830 B.n829 585
R244 B.n437 B.n436 585
R245 B.n438 B.n437 585
R246 B.n822 B.n821 585
R247 B.n823 B.n822 585
R248 B.n820 B.n443 585
R249 B.n443 B.n442 585
R250 B.n819 B.n818 585
R251 B.n818 B.n817 585
R252 B.n445 B.n444 585
R253 B.n446 B.n445 585
R254 B.n810 B.n809 585
R255 B.n811 B.n810 585
R256 B.n808 B.n451 585
R257 B.n451 B.n450 585
R258 B.n807 B.n806 585
R259 B.n806 B.n805 585
R260 B.n453 B.n452 585
R261 B.n454 B.n453 585
R262 B.n798 B.n797 585
R263 B.n799 B.n798 585
R264 B.n796 B.n459 585
R265 B.n459 B.n458 585
R266 B.n791 B.n790 585
R267 B.n789 B.n527 585
R268 B.n788 B.n526 585
R269 B.n793 B.n526 585
R270 B.n787 B.n786 585
R271 B.n785 B.n784 585
R272 B.n783 B.n782 585
R273 B.n781 B.n780 585
R274 B.n779 B.n778 585
R275 B.n777 B.n776 585
R276 B.n775 B.n774 585
R277 B.n773 B.n772 585
R278 B.n771 B.n770 585
R279 B.n769 B.n768 585
R280 B.n767 B.n766 585
R281 B.n765 B.n764 585
R282 B.n763 B.n762 585
R283 B.n761 B.n760 585
R284 B.n759 B.n758 585
R285 B.n757 B.n756 585
R286 B.n755 B.n754 585
R287 B.n753 B.n752 585
R288 B.n751 B.n750 585
R289 B.n749 B.n748 585
R290 B.n747 B.n746 585
R291 B.n745 B.n744 585
R292 B.n743 B.n742 585
R293 B.n741 B.n740 585
R294 B.n739 B.n738 585
R295 B.n737 B.n736 585
R296 B.n735 B.n734 585
R297 B.n733 B.n732 585
R298 B.n731 B.n730 585
R299 B.n729 B.n728 585
R300 B.n727 B.n726 585
R301 B.n725 B.n724 585
R302 B.n723 B.n722 585
R303 B.n721 B.n720 585
R304 B.n719 B.n718 585
R305 B.n717 B.n716 585
R306 B.n715 B.n714 585
R307 B.n713 B.n712 585
R308 B.n711 B.n710 585
R309 B.n709 B.n708 585
R310 B.n707 B.n706 585
R311 B.n705 B.n704 585
R312 B.n703 B.n702 585
R313 B.n701 B.n700 585
R314 B.n699 B.n698 585
R315 B.n697 B.n696 585
R316 B.n695 B.n694 585
R317 B.n693 B.n692 585
R318 B.n691 B.n690 585
R319 B.n689 B.n688 585
R320 B.n687 B.n686 585
R321 B.n685 B.n684 585
R322 B.n683 B.n682 585
R323 B.n681 B.n680 585
R324 B.n679 B.n678 585
R325 B.n677 B.n676 585
R326 B.n675 B.n674 585
R327 B.n673 B.n672 585
R328 B.n671 B.n670 585
R329 B.n669 B.n668 585
R330 B.n667 B.n666 585
R331 B.n665 B.n664 585
R332 B.n663 B.n662 585
R333 B.n661 B.n660 585
R334 B.n659 B.n658 585
R335 B.n657 B.n656 585
R336 B.n655 B.n654 585
R337 B.n653 B.n652 585
R338 B.n651 B.n650 585
R339 B.n649 B.n648 585
R340 B.n647 B.n646 585
R341 B.n645 B.n644 585
R342 B.n643 B.n642 585
R343 B.n641 B.n640 585
R344 B.n639 B.n638 585
R345 B.n637 B.n636 585
R346 B.n635 B.n634 585
R347 B.n633 B.n632 585
R348 B.n631 B.n630 585
R349 B.n629 B.n628 585
R350 B.n627 B.n626 585
R351 B.n625 B.n624 585
R352 B.n623 B.n622 585
R353 B.n621 B.n620 585
R354 B.n619 B.n618 585
R355 B.n617 B.n616 585
R356 B.n615 B.n614 585
R357 B.n613 B.n612 585
R358 B.n611 B.n610 585
R359 B.n609 B.n608 585
R360 B.n607 B.n606 585
R361 B.n605 B.n604 585
R362 B.n603 B.n602 585
R363 B.n601 B.n600 585
R364 B.n599 B.n598 585
R365 B.n597 B.n596 585
R366 B.n595 B.n594 585
R367 B.n593 B.n592 585
R368 B.n591 B.n590 585
R369 B.n589 B.n588 585
R370 B.n587 B.n586 585
R371 B.n585 B.n584 585
R372 B.n583 B.n582 585
R373 B.n581 B.n580 585
R374 B.n579 B.n578 585
R375 B.n577 B.n576 585
R376 B.n575 B.n574 585
R377 B.n573 B.n572 585
R378 B.n571 B.n570 585
R379 B.n569 B.n568 585
R380 B.n567 B.n566 585
R381 B.n565 B.n564 585
R382 B.n563 B.n562 585
R383 B.n561 B.n560 585
R384 B.n559 B.n558 585
R385 B.n557 B.n556 585
R386 B.n555 B.n554 585
R387 B.n553 B.n552 585
R388 B.n551 B.n550 585
R389 B.n549 B.n548 585
R390 B.n547 B.n546 585
R391 B.n545 B.n544 585
R392 B.n543 B.n542 585
R393 B.n541 B.n540 585
R394 B.n539 B.n538 585
R395 B.n537 B.n536 585
R396 B.n535 B.n534 585
R397 B.n461 B.n460 585
R398 B.n795 B.n794 585
R399 B.n794 B.n793 585
R400 B.n457 B.n456 585
R401 B.n458 B.n457 585
R402 B.n801 B.n800 585
R403 B.n800 B.n799 585
R404 B.n802 B.n455 585
R405 B.n455 B.n454 585
R406 B.n804 B.n803 585
R407 B.n805 B.n804 585
R408 B.n449 B.n448 585
R409 B.n450 B.n449 585
R410 B.n813 B.n812 585
R411 B.n812 B.n811 585
R412 B.n814 B.n447 585
R413 B.n447 B.n446 585
R414 B.n816 B.n815 585
R415 B.n817 B.n816 585
R416 B.n441 B.n440 585
R417 B.n442 B.n441 585
R418 B.n825 B.n824 585
R419 B.n824 B.n823 585
R420 B.n826 B.n439 585
R421 B.n439 B.n438 585
R422 B.n828 B.n827 585
R423 B.n829 B.n828 585
R424 B.n433 B.n432 585
R425 B.n434 B.n433 585
R426 B.n837 B.n836 585
R427 B.n836 B.n835 585
R428 B.n838 B.n431 585
R429 B.n431 B.n430 585
R430 B.n840 B.n839 585
R431 B.n841 B.n840 585
R432 B.n425 B.n424 585
R433 B.n426 B.n425 585
R434 B.n849 B.n848 585
R435 B.n848 B.n847 585
R436 B.n850 B.n423 585
R437 B.n423 B.n422 585
R438 B.n852 B.n851 585
R439 B.n853 B.n852 585
R440 B.n417 B.n416 585
R441 B.n418 B.n417 585
R442 B.n861 B.n860 585
R443 B.n860 B.n859 585
R444 B.n862 B.n415 585
R445 B.n415 B.n414 585
R446 B.n864 B.n863 585
R447 B.n865 B.n864 585
R448 B.n409 B.n408 585
R449 B.n410 B.n409 585
R450 B.n873 B.n872 585
R451 B.n872 B.n871 585
R452 B.n874 B.n407 585
R453 B.n407 B.n406 585
R454 B.n876 B.n875 585
R455 B.n877 B.n876 585
R456 B.n401 B.n400 585
R457 B.n402 B.n401 585
R458 B.n886 B.n885 585
R459 B.n885 B.n884 585
R460 B.n887 B.n399 585
R461 B.n399 B.n398 585
R462 B.n889 B.n888 585
R463 B.n890 B.n889 585
R464 B.n2 B.n0 585
R465 B.n4 B.n2 585
R466 B.n3 B.n1 585
R467 B.n1004 B.n3 585
R468 B.n1002 B.n1001 585
R469 B.n1003 B.n1002 585
R470 B.n1000 B.n9 585
R471 B.n9 B.n8 585
R472 B.n999 B.n998 585
R473 B.n998 B.n997 585
R474 B.n11 B.n10 585
R475 B.n996 B.n11 585
R476 B.n994 B.n993 585
R477 B.n995 B.n994 585
R478 B.n992 B.n16 585
R479 B.n16 B.n15 585
R480 B.n991 B.n990 585
R481 B.n990 B.n989 585
R482 B.n18 B.n17 585
R483 B.n988 B.n18 585
R484 B.n986 B.n985 585
R485 B.n987 B.n986 585
R486 B.n984 B.n23 585
R487 B.n23 B.n22 585
R488 B.n983 B.n982 585
R489 B.n982 B.n981 585
R490 B.n25 B.n24 585
R491 B.n980 B.n25 585
R492 B.n978 B.n977 585
R493 B.n979 B.n978 585
R494 B.n976 B.n30 585
R495 B.n30 B.n29 585
R496 B.n975 B.n974 585
R497 B.n974 B.n973 585
R498 B.n32 B.n31 585
R499 B.n972 B.n32 585
R500 B.n970 B.n969 585
R501 B.n971 B.n970 585
R502 B.n968 B.n37 585
R503 B.n37 B.n36 585
R504 B.n967 B.n966 585
R505 B.n966 B.n965 585
R506 B.n39 B.n38 585
R507 B.n964 B.n39 585
R508 B.n962 B.n961 585
R509 B.n963 B.n962 585
R510 B.n960 B.n44 585
R511 B.n44 B.n43 585
R512 B.n959 B.n958 585
R513 B.n958 B.n957 585
R514 B.n46 B.n45 585
R515 B.n956 B.n46 585
R516 B.n954 B.n953 585
R517 B.n955 B.n954 585
R518 B.n952 B.n51 585
R519 B.n51 B.n50 585
R520 B.n951 B.n950 585
R521 B.n950 B.n949 585
R522 B.n53 B.n52 585
R523 B.n948 B.n53 585
R524 B.n946 B.n945 585
R525 B.n947 B.n946 585
R526 B.n944 B.n58 585
R527 B.n58 B.n57 585
R528 B.n943 B.n942 585
R529 B.n942 B.n941 585
R530 B.n60 B.n59 585
R531 B.n940 B.n60 585
R532 B.n1007 B.n1006 585
R533 B.n1006 B.n1005 585
R534 B.n791 B.n457 444.452
R535 B.n133 B.n60 444.452
R536 B.n794 B.n459 444.452
R537 B.n937 B.n62 444.452
R538 B.n531 B.t15 389.421
R539 B.n528 B.t8 389.421
R540 B.n131 B.t4 389.421
R541 B.n129 B.t12 389.421
R542 B.n939 B.n938 256.663
R543 B.n939 B.n127 256.663
R544 B.n939 B.n126 256.663
R545 B.n939 B.n125 256.663
R546 B.n939 B.n124 256.663
R547 B.n939 B.n123 256.663
R548 B.n939 B.n122 256.663
R549 B.n939 B.n121 256.663
R550 B.n939 B.n120 256.663
R551 B.n939 B.n119 256.663
R552 B.n939 B.n118 256.663
R553 B.n939 B.n117 256.663
R554 B.n939 B.n116 256.663
R555 B.n939 B.n115 256.663
R556 B.n939 B.n114 256.663
R557 B.n939 B.n113 256.663
R558 B.n939 B.n112 256.663
R559 B.n939 B.n111 256.663
R560 B.n939 B.n110 256.663
R561 B.n939 B.n109 256.663
R562 B.n939 B.n108 256.663
R563 B.n939 B.n107 256.663
R564 B.n939 B.n106 256.663
R565 B.n939 B.n105 256.663
R566 B.n939 B.n104 256.663
R567 B.n939 B.n103 256.663
R568 B.n939 B.n102 256.663
R569 B.n939 B.n101 256.663
R570 B.n939 B.n100 256.663
R571 B.n939 B.n99 256.663
R572 B.n939 B.n98 256.663
R573 B.n939 B.n97 256.663
R574 B.n939 B.n96 256.663
R575 B.n939 B.n95 256.663
R576 B.n939 B.n94 256.663
R577 B.n939 B.n93 256.663
R578 B.n939 B.n92 256.663
R579 B.n939 B.n91 256.663
R580 B.n939 B.n90 256.663
R581 B.n939 B.n89 256.663
R582 B.n939 B.n88 256.663
R583 B.n939 B.n87 256.663
R584 B.n939 B.n86 256.663
R585 B.n939 B.n85 256.663
R586 B.n939 B.n84 256.663
R587 B.n939 B.n83 256.663
R588 B.n939 B.n82 256.663
R589 B.n939 B.n81 256.663
R590 B.n939 B.n80 256.663
R591 B.n939 B.n79 256.663
R592 B.n939 B.n78 256.663
R593 B.n939 B.n77 256.663
R594 B.n939 B.n76 256.663
R595 B.n939 B.n75 256.663
R596 B.n939 B.n74 256.663
R597 B.n939 B.n73 256.663
R598 B.n939 B.n72 256.663
R599 B.n939 B.n71 256.663
R600 B.n939 B.n70 256.663
R601 B.n939 B.n69 256.663
R602 B.n939 B.n68 256.663
R603 B.n939 B.n67 256.663
R604 B.n939 B.n66 256.663
R605 B.n939 B.n65 256.663
R606 B.n939 B.n64 256.663
R607 B.n939 B.n63 256.663
R608 B.n793 B.n792 256.663
R609 B.n793 B.n462 256.663
R610 B.n793 B.n463 256.663
R611 B.n793 B.n464 256.663
R612 B.n793 B.n465 256.663
R613 B.n793 B.n466 256.663
R614 B.n793 B.n467 256.663
R615 B.n793 B.n468 256.663
R616 B.n793 B.n469 256.663
R617 B.n793 B.n470 256.663
R618 B.n793 B.n471 256.663
R619 B.n793 B.n472 256.663
R620 B.n793 B.n473 256.663
R621 B.n793 B.n474 256.663
R622 B.n793 B.n475 256.663
R623 B.n793 B.n476 256.663
R624 B.n793 B.n477 256.663
R625 B.n793 B.n478 256.663
R626 B.n793 B.n479 256.663
R627 B.n793 B.n480 256.663
R628 B.n793 B.n481 256.663
R629 B.n793 B.n482 256.663
R630 B.n793 B.n483 256.663
R631 B.n793 B.n484 256.663
R632 B.n793 B.n485 256.663
R633 B.n793 B.n486 256.663
R634 B.n793 B.n487 256.663
R635 B.n793 B.n488 256.663
R636 B.n793 B.n489 256.663
R637 B.n793 B.n490 256.663
R638 B.n793 B.n491 256.663
R639 B.n793 B.n492 256.663
R640 B.n793 B.n493 256.663
R641 B.n793 B.n494 256.663
R642 B.n793 B.n495 256.663
R643 B.n793 B.n496 256.663
R644 B.n793 B.n497 256.663
R645 B.n793 B.n498 256.663
R646 B.n793 B.n499 256.663
R647 B.n793 B.n500 256.663
R648 B.n793 B.n501 256.663
R649 B.n793 B.n502 256.663
R650 B.n793 B.n503 256.663
R651 B.n793 B.n504 256.663
R652 B.n793 B.n505 256.663
R653 B.n793 B.n506 256.663
R654 B.n793 B.n507 256.663
R655 B.n793 B.n508 256.663
R656 B.n793 B.n509 256.663
R657 B.n793 B.n510 256.663
R658 B.n793 B.n511 256.663
R659 B.n793 B.n512 256.663
R660 B.n793 B.n513 256.663
R661 B.n793 B.n514 256.663
R662 B.n793 B.n515 256.663
R663 B.n793 B.n516 256.663
R664 B.n793 B.n517 256.663
R665 B.n793 B.n518 256.663
R666 B.n793 B.n519 256.663
R667 B.n793 B.n520 256.663
R668 B.n793 B.n521 256.663
R669 B.n793 B.n522 256.663
R670 B.n793 B.n523 256.663
R671 B.n793 B.n524 256.663
R672 B.n793 B.n525 256.663
R673 B.n800 B.n457 163.367
R674 B.n800 B.n455 163.367
R675 B.n804 B.n455 163.367
R676 B.n804 B.n449 163.367
R677 B.n812 B.n449 163.367
R678 B.n812 B.n447 163.367
R679 B.n816 B.n447 163.367
R680 B.n816 B.n441 163.367
R681 B.n824 B.n441 163.367
R682 B.n824 B.n439 163.367
R683 B.n828 B.n439 163.367
R684 B.n828 B.n433 163.367
R685 B.n836 B.n433 163.367
R686 B.n836 B.n431 163.367
R687 B.n840 B.n431 163.367
R688 B.n840 B.n425 163.367
R689 B.n848 B.n425 163.367
R690 B.n848 B.n423 163.367
R691 B.n852 B.n423 163.367
R692 B.n852 B.n417 163.367
R693 B.n860 B.n417 163.367
R694 B.n860 B.n415 163.367
R695 B.n864 B.n415 163.367
R696 B.n864 B.n409 163.367
R697 B.n872 B.n409 163.367
R698 B.n872 B.n407 163.367
R699 B.n876 B.n407 163.367
R700 B.n876 B.n401 163.367
R701 B.n885 B.n401 163.367
R702 B.n885 B.n399 163.367
R703 B.n889 B.n399 163.367
R704 B.n889 B.n2 163.367
R705 B.n1006 B.n2 163.367
R706 B.n1006 B.n3 163.367
R707 B.n1002 B.n3 163.367
R708 B.n1002 B.n9 163.367
R709 B.n998 B.n9 163.367
R710 B.n998 B.n11 163.367
R711 B.n994 B.n11 163.367
R712 B.n994 B.n16 163.367
R713 B.n990 B.n16 163.367
R714 B.n990 B.n18 163.367
R715 B.n986 B.n18 163.367
R716 B.n986 B.n23 163.367
R717 B.n982 B.n23 163.367
R718 B.n982 B.n25 163.367
R719 B.n978 B.n25 163.367
R720 B.n978 B.n30 163.367
R721 B.n974 B.n30 163.367
R722 B.n974 B.n32 163.367
R723 B.n970 B.n32 163.367
R724 B.n970 B.n37 163.367
R725 B.n966 B.n37 163.367
R726 B.n966 B.n39 163.367
R727 B.n962 B.n39 163.367
R728 B.n962 B.n44 163.367
R729 B.n958 B.n44 163.367
R730 B.n958 B.n46 163.367
R731 B.n954 B.n46 163.367
R732 B.n954 B.n51 163.367
R733 B.n950 B.n51 163.367
R734 B.n950 B.n53 163.367
R735 B.n946 B.n53 163.367
R736 B.n946 B.n58 163.367
R737 B.n942 B.n58 163.367
R738 B.n942 B.n60 163.367
R739 B.n527 B.n526 163.367
R740 B.n786 B.n526 163.367
R741 B.n784 B.n783 163.367
R742 B.n780 B.n779 163.367
R743 B.n776 B.n775 163.367
R744 B.n772 B.n771 163.367
R745 B.n768 B.n767 163.367
R746 B.n764 B.n763 163.367
R747 B.n760 B.n759 163.367
R748 B.n756 B.n755 163.367
R749 B.n752 B.n751 163.367
R750 B.n748 B.n747 163.367
R751 B.n744 B.n743 163.367
R752 B.n740 B.n739 163.367
R753 B.n736 B.n735 163.367
R754 B.n732 B.n731 163.367
R755 B.n728 B.n727 163.367
R756 B.n724 B.n723 163.367
R757 B.n720 B.n719 163.367
R758 B.n716 B.n715 163.367
R759 B.n712 B.n711 163.367
R760 B.n708 B.n707 163.367
R761 B.n704 B.n703 163.367
R762 B.n700 B.n699 163.367
R763 B.n696 B.n695 163.367
R764 B.n692 B.n691 163.367
R765 B.n688 B.n687 163.367
R766 B.n684 B.n683 163.367
R767 B.n680 B.n679 163.367
R768 B.n676 B.n675 163.367
R769 B.n672 B.n671 163.367
R770 B.n668 B.n667 163.367
R771 B.n664 B.n663 163.367
R772 B.n660 B.n659 163.367
R773 B.n656 B.n655 163.367
R774 B.n652 B.n651 163.367
R775 B.n648 B.n647 163.367
R776 B.n644 B.n643 163.367
R777 B.n640 B.n639 163.367
R778 B.n636 B.n635 163.367
R779 B.n632 B.n631 163.367
R780 B.n628 B.n627 163.367
R781 B.n624 B.n623 163.367
R782 B.n620 B.n619 163.367
R783 B.n616 B.n615 163.367
R784 B.n612 B.n611 163.367
R785 B.n608 B.n607 163.367
R786 B.n604 B.n603 163.367
R787 B.n600 B.n599 163.367
R788 B.n596 B.n595 163.367
R789 B.n592 B.n591 163.367
R790 B.n588 B.n587 163.367
R791 B.n584 B.n583 163.367
R792 B.n580 B.n579 163.367
R793 B.n576 B.n575 163.367
R794 B.n572 B.n571 163.367
R795 B.n568 B.n567 163.367
R796 B.n564 B.n563 163.367
R797 B.n560 B.n559 163.367
R798 B.n556 B.n555 163.367
R799 B.n552 B.n551 163.367
R800 B.n548 B.n547 163.367
R801 B.n544 B.n543 163.367
R802 B.n540 B.n539 163.367
R803 B.n536 B.n535 163.367
R804 B.n794 B.n461 163.367
R805 B.n798 B.n459 163.367
R806 B.n798 B.n453 163.367
R807 B.n806 B.n453 163.367
R808 B.n806 B.n451 163.367
R809 B.n810 B.n451 163.367
R810 B.n810 B.n445 163.367
R811 B.n818 B.n445 163.367
R812 B.n818 B.n443 163.367
R813 B.n822 B.n443 163.367
R814 B.n822 B.n437 163.367
R815 B.n830 B.n437 163.367
R816 B.n830 B.n435 163.367
R817 B.n834 B.n435 163.367
R818 B.n834 B.n429 163.367
R819 B.n842 B.n429 163.367
R820 B.n842 B.n427 163.367
R821 B.n846 B.n427 163.367
R822 B.n846 B.n421 163.367
R823 B.n854 B.n421 163.367
R824 B.n854 B.n419 163.367
R825 B.n858 B.n419 163.367
R826 B.n858 B.n413 163.367
R827 B.n866 B.n413 163.367
R828 B.n866 B.n411 163.367
R829 B.n870 B.n411 163.367
R830 B.n870 B.n405 163.367
R831 B.n878 B.n405 163.367
R832 B.n878 B.n403 163.367
R833 B.n883 B.n403 163.367
R834 B.n883 B.n397 163.367
R835 B.n891 B.n397 163.367
R836 B.n892 B.n891 163.367
R837 B.n892 B.n5 163.367
R838 B.n6 B.n5 163.367
R839 B.n7 B.n6 163.367
R840 B.n897 B.n7 163.367
R841 B.n897 B.n12 163.367
R842 B.n13 B.n12 163.367
R843 B.n14 B.n13 163.367
R844 B.n902 B.n14 163.367
R845 B.n902 B.n19 163.367
R846 B.n20 B.n19 163.367
R847 B.n21 B.n20 163.367
R848 B.n907 B.n21 163.367
R849 B.n907 B.n26 163.367
R850 B.n27 B.n26 163.367
R851 B.n28 B.n27 163.367
R852 B.n912 B.n28 163.367
R853 B.n912 B.n33 163.367
R854 B.n34 B.n33 163.367
R855 B.n35 B.n34 163.367
R856 B.n917 B.n35 163.367
R857 B.n917 B.n40 163.367
R858 B.n41 B.n40 163.367
R859 B.n42 B.n41 163.367
R860 B.n922 B.n42 163.367
R861 B.n922 B.n47 163.367
R862 B.n48 B.n47 163.367
R863 B.n49 B.n48 163.367
R864 B.n927 B.n49 163.367
R865 B.n927 B.n54 163.367
R866 B.n55 B.n54 163.367
R867 B.n56 B.n55 163.367
R868 B.n932 B.n56 163.367
R869 B.n932 B.n61 163.367
R870 B.n62 B.n61 163.367
R871 B.n137 B.n136 163.367
R872 B.n141 B.n140 163.367
R873 B.n145 B.n144 163.367
R874 B.n149 B.n148 163.367
R875 B.n153 B.n152 163.367
R876 B.n157 B.n156 163.367
R877 B.n161 B.n160 163.367
R878 B.n165 B.n164 163.367
R879 B.n169 B.n168 163.367
R880 B.n173 B.n172 163.367
R881 B.n177 B.n176 163.367
R882 B.n181 B.n180 163.367
R883 B.n185 B.n184 163.367
R884 B.n189 B.n188 163.367
R885 B.n193 B.n192 163.367
R886 B.n197 B.n196 163.367
R887 B.n201 B.n200 163.367
R888 B.n205 B.n204 163.367
R889 B.n209 B.n208 163.367
R890 B.n213 B.n212 163.367
R891 B.n217 B.n216 163.367
R892 B.n221 B.n220 163.367
R893 B.n225 B.n224 163.367
R894 B.n229 B.n228 163.367
R895 B.n233 B.n232 163.367
R896 B.n237 B.n236 163.367
R897 B.n241 B.n240 163.367
R898 B.n245 B.n244 163.367
R899 B.n249 B.n248 163.367
R900 B.n253 B.n252 163.367
R901 B.n258 B.n257 163.367
R902 B.n262 B.n261 163.367
R903 B.n266 B.n265 163.367
R904 B.n270 B.n269 163.367
R905 B.n274 B.n273 163.367
R906 B.n279 B.n278 163.367
R907 B.n283 B.n282 163.367
R908 B.n287 B.n286 163.367
R909 B.n291 B.n290 163.367
R910 B.n295 B.n294 163.367
R911 B.n299 B.n298 163.367
R912 B.n303 B.n302 163.367
R913 B.n307 B.n306 163.367
R914 B.n311 B.n310 163.367
R915 B.n315 B.n314 163.367
R916 B.n319 B.n318 163.367
R917 B.n323 B.n322 163.367
R918 B.n327 B.n326 163.367
R919 B.n331 B.n330 163.367
R920 B.n335 B.n334 163.367
R921 B.n339 B.n338 163.367
R922 B.n343 B.n342 163.367
R923 B.n347 B.n346 163.367
R924 B.n351 B.n350 163.367
R925 B.n355 B.n354 163.367
R926 B.n359 B.n358 163.367
R927 B.n363 B.n362 163.367
R928 B.n367 B.n366 163.367
R929 B.n371 B.n370 163.367
R930 B.n375 B.n374 163.367
R931 B.n379 B.n378 163.367
R932 B.n383 B.n382 163.367
R933 B.n387 B.n386 163.367
R934 B.n391 B.n390 163.367
R935 B.n393 B.n128 163.367
R936 B.n531 B.t17 126.365
R937 B.n129 B.t13 126.365
R938 B.n528 B.t11 126.341
R939 B.n131 B.t6 126.341
R940 B.n532 B.t16 72.0618
R941 B.n130 B.t14 72.0618
R942 B.n529 B.t10 72.0371
R943 B.n132 B.t7 72.0371
R944 B.n792 B.n791 71.676
R945 B.n786 B.n462 71.676
R946 B.n783 B.n463 71.676
R947 B.n779 B.n464 71.676
R948 B.n775 B.n465 71.676
R949 B.n771 B.n466 71.676
R950 B.n767 B.n467 71.676
R951 B.n763 B.n468 71.676
R952 B.n759 B.n469 71.676
R953 B.n755 B.n470 71.676
R954 B.n751 B.n471 71.676
R955 B.n747 B.n472 71.676
R956 B.n743 B.n473 71.676
R957 B.n739 B.n474 71.676
R958 B.n735 B.n475 71.676
R959 B.n731 B.n476 71.676
R960 B.n727 B.n477 71.676
R961 B.n723 B.n478 71.676
R962 B.n719 B.n479 71.676
R963 B.n715 B.n480 71.676
R964 B.n711 B.n481 71.676
R965 B.n707 B.n482 71.676
R966 B.n703 B.n483 71.676
R967 B.n699 B.n484 71.676
R968 B.n695 B.n485 71.676
R969 B.n691 B.n486 71.676
R970 B.n687 B.n487 71.676
R971 B.n683 B.n488 71.676
R972 B.n679 B.n489 71.676
R973 B.n675 B.n490 71.676
R974 B.n671 B.n491 71.676
R975 B.n667 B.n492 71.676
R976 B.n663 B.n493 71.676
R977 B.n659 B.n494 71.676
R978 B.n655 B.n495 71.676
R979 B.n651 B.n496 71.676
R980 B.n647 B.n497 71.676
R981 B.n643 B.n498 71.676
R982 B.n639 B.n499 71.676
R983 B.n635 B.n500 71.676
R984 B.n631 B.n501 71.676
R985 B.n627 B.n502 71.676
R986 B.n623 B.n503 71.676
R987 B.n619 B.n504 71.676
R988 B.n615 B.n505 71.676
R989 B.n611 B.n506 71.676
R990 B.n607 B.n507 71.676
R991 B.n603 B.n508 71.676
R992 B.n599 B.n509 71.676
R993 B.n595 B.n510 71.676
R994 B.n591 B.n511 71.676
R995 B.n587 B.n512 71.676
R996 B.n583 B.n513 71.676
R997 B.n579 B.n514 71.676
R998 B.n575 B.n515 71.676
R999 B.n571 B.n516 71.676
R1000 B.n567 B.n517 71.676
R1001 B.n563 B.n518 71.676
R1002 B.n559 B.n519 71.676
R1003 B.n555 B.n520 71.676
R1004 B.n551 B.n521 71.676
R1005 B.n547 B.n522 71.676
R1006 B.n543 B.n523 71.676
R1007 B.n539 B.n524 71.676
R1008 B.n535 B.n525 71.676
R1009 B.n133 B.n63 71.676
R1010 B.n137 B.n64 71.676
R1011 B.n141 B.n65 71.676
R1012 B.n145 B.n66 71.676
R1013 B.n149 B.n67 71.676
R1014 B.n153 B.n68 71.676
R1015 B.n157 B.n69 71.676
R1016 B.n161 B.n70 71.676
R1017 B.n165 B.n71 71.676
R1018 B.n169 B.n72 71.676
R1019 B.n173 B.n73 71.676
R1020 B.n177 B.n74 71.676
R1021 B.n181 B.n75 71.676
R1022 B.n185 B.n76 71.676
R1023 B.n189 B.n77 71.676
R1024 B.n193 B.n78 71.676
R1025 B.n197 B.n79 71.676
R1026 B.n201 B.n80 71.676
R1027 B.n205 B.n81 71.676
R1028 B.n209 B.n82 71.676
R1029 B.n213 B.n83 71.676
R1030 B.n217 B.n84 71.676
R1031 B.n221 B.n85 71.676
R1032 B.n225 B.n86 71.676
R1033 B.n229 B.n87 71.676
R1034 B.n233 B.n88 71.676
R1035 B.n237 B.n89 71.676
R1036 B.n241 B.n90 71.676
R1037 B.n245 B.n91 71.676
R1038 B.n249 B.n92 71.676
R1039 B.n253 B.n93 71.676
R1040 B.n258 B.n94 71.676
R1041 B.n262 B.n95 71.676
R1042 B.n266 B.n96 71.676
R1043 B.n270 B.n97 71.676
R1044 B.n274 B.n98 71.676
R1045 B.n279 B.n99 71.676
R1046 B.n283 B.n100 71.676
R1047 B.n287 B.n101 71.676
R1048 B.n291 B.n102 71.676
R1049 B.n295 B.n103 71.676
R1050 B.n299 B.n104 71.676
R1051 B.n303 B.n105 71.676
R1052 B.n307 B.n106 71.676
R1053 B.n311 B.n107 71.676
R1054 B.n315 B.n108 71.676
R1055 B.n319 B.n109 71.676
R1056 B.n323 B.n110 71.676
R1057 B.n327 B.n111 71.676
R1058 B.n331 B.n112 71.676
R1059 B.n335 B.n113 71.676
R1060 B.n339 B.n114 71.676
R1061 B.n343 B.n115 71.676
R1062 B.n347 B.n116 71.676
R1063 B.n351 B.n117 71.676
R1064 B.n355 B.n118 71.676
R1065 B.n359 B.n119 71.676
R1066 B.n363 B.n120 71.676
R1067 B.n367 B.n121 71.676
R1068 B.n371 B.n122 71.676
R1069 B.n375 B.n123 71.676
R1070 B.n379 B.n124 71.676
R1071 B.n383 B.n125 71.676
R1072 B.n387 B.n126 71.676
R1073 B.n391 B.n127 71.676
R1074 B.n938 B.n128 71.676
R1075 B.n938 B.n937 71.676
R1076 B.n393 B.n127 71.676
R1077 B.n390 B.n126 71.676
R1078 B.n386 B.n125 71.676
R1079 B.n382 B.n124 71.676
R1080 B.n378 B.n123 71.676
R1081 B.n374 B.n122 71.676
R1082 B.n370 B.n121 71.676
R1083 B.n366 B.n120 71.676
R1084 B.n362 B.n119 71.676
R1085 B.n358 B.n118 71.676
R1086 B.n354 B.n117 71.676
R1087 B.n350 B.n116 71.676
R1088 B.n346 B.n115 71.676
R1089 B.n342 B.n114 71.676
R1090 B.n338 B.n113 71.676
R1091 B.n334 B.n112 71.676
R1092 B.n330 B.n111 71.676
R1093 B.n326 B.n110 71.676
R1094 B.n322 B.n109 71.676
R1095 B.n318 B.n108 71.676
R1096 B.n314 B.n107 71.676
R1097 B.n310 B.n106 71.676
R1098 B.n306 B.n105 71.676
R1099 B.n302 B.n104 71.676
R1100 B.n298 B.n103 71.676
R1101 B.n294 B.n102 71.676
R1102 B.n290 B.n101 71.676
R1103 B.n286 B.n100 71.676
R1104 B.n282 B.n99 71.676
R1105 B.n278 B.n98 71.676
R1106 B.n273 B.n97 71.676
R1107 B.n269 B.n96 71.676
R1108 B.n265 B.n95 71.676
R1109 B.n261 B.n94 71.676
R1110 B.n257 B.n93 71.676
R1111 B.n252 B.n92 71.676
R1112 B.n248 B.n91 71.676
R1113 B.n244 B.n90 71.676
R1114 B.n240 B.n89 71.676
R1115 B.n236 B.n88 71.676
R1116 B.n232 B.n87 71.676
R1117 B.n228 B.n86 71.676
R1118 B.n224 B.n85 71.676
R1119 B.n220 B.n84 71.676
R1120 B.n216 B.n83 71.676
R1121 B.n212 B.n82 71.676
R1122 B.n208 B.n81 71.676
R1123 B.n204 B.n80 71.676
R1124 B.n200 B.n79 71.676
R1125 B.n196 B.n78 71.676
R1126 B.n192 B.n77 71.676
R1127 B.n188 B.n76 71.676
R1128 B.n184 B.n75 71.676
R1129 B.n180 B.n74 71.676
R1130 B.n176 B.n73 71.676
R1131 B.n172 B.n72 71.676
R1132 B.n168 B.n71 71.676
R1133 B.n164 B.n70 71.676
R1134 B.n160 B.n69 71.676
R1135 B.n156 B.n68 71.676
R1136 B.n152 B.n67 71.676
R1137 B.n148 B.n66 71.676
R1138 B.n144 B.n65 71.676
R1139 B.n140 B.n64 71.676
R1140 B.n136 B.n63 71.676
R1141 B.n792 B.n527 71.676
R1142 B.n784 B.n462 71.676
R1143 B.n780 B.n463 71.676
R1144 B.n776 B.n464 71.676
R1145 B.n772 B.n465 71.676
R1146 B.n768 B.n466 71.676
R1147 B.n764 B.n467 71.676
R1148 B.n760 B.n468 71.676
R1149 B.n756 B.n469 71.676
R1150 B.n752 B.n470 71.676
R1151 B.n748 B.n471 71.676
R1152 B.n744 B.n472 71.676
R1153 B.n740 B.n473 71.676
R1154 B.n736 B.n474 71.676
R1155 B.n732 B.n475 71.676
R1156 B.n728 B.n476 71.676
R1157 B.n724 B.n477 71.676
R1158 B.n720 B.n478 71.676
R1159 B.n716 B.n479 71.676
R1160 B.n712 B.n480 71.676
R1161 B.n708 B.n481 71.676
R1162 B.n704 B.n482 71.676
R1163 B.n700 B.n483 71.676
R1164 B.n696 B.n484 71.676
R1165 B.n692 B.n485 71.676
R1166 B.n688 B.n486 71.676
R1167 B.n684 B.n487 71.676
R1168 B.n680 B.n488 71.676
R1169 B.n676 B.n489 71.676
R1170 B.n672 B.n490 71.676
R1171 B.n668 B.n491 71.676
R1172 B.n664 B.n492 71.676
R1173 B.n660 B.n493 71.676
R1174 B.n656 B.n494 71.676
R1175 B.n652 B.n495 71.676
R1176 B.n648 B.n496 71.676
R1177 B.n644 B.n497 71.676
R1178 B.n640 B.n498 71.676
R1179 B.n636 B.n499 71.676
R1180 B.n632 B.n500 71.676
R1181 B.n628 B.n501 71.676
R1182 B.n624 B.n502 71.676
R1183 B.n620 B.n503 71.676
R1184 B.n616 B.n504 71.676
R1185 B.n612 B.n505 71.676
R1186 B.n608 B.n506 71.676
R1187 B.n604 B.n507 71.676
R1188 B.n600 B.n508 71.676
R1189 B.n596 B.n509 71.676
R1190 B.n592 B.n510 71.676
R1191 B.n588 B.n511 71.676
R1192 B.n584 B.n512 71.676
R1193 B.n580 B.n513 71.676
R1194 B.n576 B.n514 71.676
R1195 B.n572 B.n515 71.676
R1196 B.n568 B.n516 71.676
R1197 B.n564 B.n517 71.676
R1198 B.n560 B.n518 71.676
R1199 B.n556 B.n519 71.676
R1200 B.n552 B.n520 71.676
R1201 B.n548 B.n521 71.676
R1202 B.n544 B.n522 71.676
R1203 B.n540 B.n523 71.676
R1204 B.n536 B.n524 71.676
R1205 B.n525 B.n461 71.676
R1206 B.n533 B.n532 59.5399
R1207 B.n530 B.n529 59.5399
R1208 B.n255 B.n132 59.5399
R1209 B.n276 B.n130 59.5399
R1210 B.n532 B.n531 54.3035
R1211 B.n529 B.n528 54.3035
R1212 B.n132 B.n131 54.3035
R1213 B.n130 B.n129 54.3035
R1214 B.n793 B.n458 51.1204
R1215 B.n940 B.n939 51.1204
R1216 B.n799 B.n458 31.3172
R1217 B.n799 B.n454 31.3172
R1218 B.n805 B.n454 31.3172
R1219 B.n805 B.n450 31.3172
R1220 B.n811 B.n450 31.3172
R1221 B.n811 B.n446 31.3172
R1222 B.n817 B.n446 31.3172
R1223 B.n823 B.n442 31.3172
R1224 B.n823 B.n438 31.3172
R1225 B.n829 B.n438 31.3172
R1226 B.n829 B.n434 31.3172
R1227 B.n835 B.n434 31.3172
R1228 B.n835 B.n430 31.3172
R1229 B.n841 B.n430 31.3172
R1230 B.n841 B.n426 31.3172
R1231 B.n847 B.n426 31.3172
R1232 B.n847 B.n422 31.3172
R1233 B.n853 B.n422 31.3172
R1234 B.n859 B.n418 31.3172
R1235 B.n859 B.n414 31.3172
R1236 B.n865 B.n414 31.3172
R1237 B.n865 B.n410 31.3172
R1238 B.n871 B.n410 31.3172
R1239 B.n871 B.n406 31.3172
R1240 B.n877 B.n406 31.3172
R1241 B.n884 B.n402 31.3172
R1242 B.n884 B.n398 31.3172
R1243 B.n890 B.n398 31.3172
R1244 B.n890 B.n4 31.3172
R1245 B.n1005 B.n4 31.3172
R1246 B.n1005 B.n1004 31.3172
R1247 B.n1004 B.n1003 31.3172
R1248 B.n1003 B.n8 31.3172
R1249 B.n997 B.n8 31.3172
R1250 B.n997 B.n996 31.3172
R1251 B.n995 B.n15 31.3172
R1252 B.n989 B.n15 31.3172
R1253 B.n989 B.n988 31.3172
R1254 B.n988 B.n987 31.3172
R1255 B.n987 B.n22 31.3172
R1256 B.n981 B.n22 31.3172
R1257 B.n981 B.n980 31.3172
R1258 B.n979 B.n29 31.3172
R1259 B.n973 B.n29 31.3172
R1260 B.n973 B.n972 31.3172
R1261 B.n972 B.n971 31.3172
R1262 B.n971 B.n36 31.3172
R1263 B.n965 B.n36 31.3172
R1264 B.n965 B.n964 31.3172
R1265 B.n964 B.n963 31.3172
R1266 B.n963 B.n43 31.3172
R1267 B.n957 B.n43 31.3172
R1268 B.n957 B.n956 31.3172
R1269 B.n955 B.n50 31.3172
R1270 B.n949 B.n50 31.3172
R1271 B.n949 B.n948 31.3172
R1272 B.n948 B.n947 31.3172
R1273 B.n947 B.n57 31.3172
R1274 B.n941 B.n57 31.3172
R1275 B.n941 B.n940 31.3172
R1276 B.t2 B.n418 29.9356
R1277 B.n980 B.t1 29.9356
R1278 B.n134 B.n59 28.8785
R1279 B.n796 B.n795 28.8785
R1280 B.n790 B.n456 28.8785
R1281 B.n936 B.n935 28.8785
R1282 B.t3 B.n402 22.567
R1283 B.n996 B.t0 22.567
R1284 B.n817 B.t9 18.8826
R1285 B.t5 B.n955 18.8826
R1286 B B.n1007 18.0485
R1287 B.t9 B.n442 12.4351
R1288 B.n956 B.t5 12.4351
R1289 B.n135 B.n134 10.6151
R1290 B.n138 B.n135 10.6151
R1291 B.n139 B.n138 10.6151
R1292 B.n142 B.n139 10.6151
R1293 B.n143 B.n142 10.6151
R1294 B.n146 B.n143 10.6151
R1295 B.n147 B.n146 10.6151
R1296 B.n150 B.n147 10.6151
R1297 B.n151 B.n150 10.6151
R1298 B.n154 B.n151 10.6151
R1299 B.n155 B.n154 10.6151
R1300 B.n158 B.n155 10.6151
R1301 B.n159 B.n158 10.6151
R1302 B.n162 B.n159 10.6151
R1303 B.n163 B.n162 10.6151
R1304 B.n166 B.n163 10.6151
R1305 B.n167 B.n166 10.6151
R1306 B.n170 B.n167 10.6151
R1307 B.n171 B.n170 10.6151
R1308 B.n174 B.n171 10.6151
R1309 B.n175 B.n174 10.6151
R1310 B.n178 B.n175 10.6151
R1311 B.n179 B.n178 10.6151
R1312 B.n182 B.n179 10.6151
R1313 B.n183 B.n182 10.6151
R1314 B.n186 B.n183 10.6151
R1315 B.n187 B.n186 10.6151
R1316 B.n190 B.n187 10.6151
R1317 B.n191 B.n190 10.6151
R1318 B.n194 B.n191 10.6151
R1319 B.n195 B.n194 10.6151
R1320 B.n198 B.n195 10.6151
R1321 B.n199 B.n198 10.6151
R1322 B.n202 B.n199 10.6151
R1323 B.n203 B.n202 10.6151
R1324 B.n206 B.n203 10.6151
R1325 B.n207 B.n206 10.6151
R1326 B.n210 B.n207 10.6151
R1327 B.n211 B.n210 10.6151
R1328 B.n214 B.n211 10.6151
R1329 B.n215 B.n214 10.6151
R1330 B.n218 B.n215 10.6151
R1331 B.n219 B.n218 10.6151
R1332 B.n222 B.n219 10.6151
R1333 B.n223 B.n222 10.6151
R1334 B.n226 B.n223 10.6151
R1335 B.n227 B.n226 10.6151
R1336 B.n230 B.n227 10.6151
R1337 B.n231 B.n230 10.6151
R1338 B.n234 B.n231 10.6151
R1339 B.n235 B.n234 10.6151
R1340 B.n238 B.n235 10.6151
R1341 B.n239 B.n238 10.6151
R1342 B.n242 B.n239 10.6151
R1343 B.n243 B.n242 10.6151
R1344 B.n246 B.n243 10.6151
R1345 B.n247 B.n246 10.6151
R1346 B.n250 B.n247 10.6151
R1347 B.n251 B.n250 10.6151
R1348 B.n254 B.n251 10.6151
R1349 B.n259 B.n256 10.6151
R1350 B.n260 B.n259 10.6151
R1351 B.n263 B.n260 10.6151
R1352 B.n264 B.n263 10.6151
R1353 B.n267 B.n264 10.6151
R1354 B.n268 B.n267 10.6151
R1355 B.n271 B.n268 10.6151
R1356 B.n272 B.n271 10.6151
R1357 B.n275 B.n272 10.6151
R1358 B.n280 B.n277 10.6151
R1359 B.n281 B.n280 10.6151
R1360 B.n284 B.n281 10.6151
R1361 B.n285 B.n284 10.6151
R1362 B.n288 B.n285 10.6151
R1363 B.n289 B.n288 10.6151
R1364 B.n292 B.n289 10.6151
R1365 B.n293 B.n292 10.6151
R1366 B.n296 B.n293 10.6151
R1367 B.n297 B.n296 10.6151
R1368 B.n300 B.n297 10.6151
R1369 B.n301 B.n300 10.6151
R1370 B.n304 B.n301 10.6151
R1371 B.n305 B.n304 10.6151
R1372 B.n308 B.n305 10.6151
R1373 B.n309 B.n308 10.6151
R1374 B.n312 B.n309 10.6151
R1375 B.n313 B.n312 10.6151
R1376 B.n316 B.n313 10.6151
R1377 B.n317 B.n316 10.6151
R1378 B.n320 B.n317 10.6151
R1379 B.n321 B.n320 10.6151
R1380 B.n324 B.n321 10.6151
R1381 B.n325 B.n324 10.6151
R1382 B.n328 B.n325 10.6151
R1383 B.n329 B.n328 10.6151
R1384 B.n332 B.n329 10.6151
R1385 B.n333 B.n332 10.6151
R1386 B.n336 B.n333 10.6151
R1387 B.n337 B.n336 10.6151
R1388 B.n340 B.n337 10.6151
R1389 B.n341 B.n340 10.6151
R1390 B.n344 B.n341 10.6151
R1391 B.n345 B.n344 10.6151
R1392 B.n348 B.n345 10.6151
R1393 B.n349 B.n348 10.6151
R1394 B.n352 B.n349 10.6151
R1395 B.n353 B.n352 10.6151
R1396 B.n356 B.n353 10.6151
R1397 B.n357 B.n356 10.6151
R1398 B.n360 B.n357 10.6151
R1399 B.n361 B.n360 10.6151
R1400 B.n364 B.n361 10.6151
R1401 B.n365 B.n364 10.6151
R1402 B.n368 B.n365 10.6151
R1403 B.n369 B.n368 10.6151
R1404 B.n372 B.n369 10.6151
R1405 B.n373 B.n372 10.6151
R1406 B.n376 B.n373 10.6151
R1407 B.n377 B.n376 10.6151
R1408 B.n380 B.n377 10.6151
R1409 B.n381 B.n380 10.6151
R1410 B.n384 B.n381 10.6151
R1411 B.n385 B.n384 10.6151
R1412 B.n388 B.n385 10.6151
R1413 B.n389 B.n388 10.6151
R1414 B.n392 B.n389 10.6151
R1415 B.n394 B.n392 10.6151
R1416 B.n395 B.n394 10.6151
R1417 B.n936 B.n395 10.6151
R1418 B.n797 B.n796 10.6151
R1419 B.n797 B.n452 10.6151
R1420 B.n807 B.n452 10.6151
R1421 B.n808 B.n807 10.6151
R1422 B.n809 B.n808 10.6151
R1423 B.n809 B.n444 10.6151
R1424 B.n819 B.n444 10.6151
R1425 B.n820 B.n819 10.6151
R1426 B.n821 B.n820 10.6151
R1427 B.n821 B.n436 10.6151
R1428 B.n831 B.n436 10.6151
R1429 B.n832 B.n831 10.6151
R1430 B.n833 B.n832 10.6151
R1431 B.n833 B.n428 10.6151
R1432 B.n843 B.n428 10.6151
R1433 B.n844 B.n843 10.6151
R1434 B.n845 B.n844 10.6151
R1435 B.n845 B.n420 10.6151
R1436 B.n855 B.n420 10.6151
R1437 B.n856 B.n855 10.6151
R1438 B.n857 B.n856 10.6151
R1439 B.n857 B.n412 10.6151
R1440 B.n867 B.n412 10.6151
R1441 B.n868 B.n867 10.6151
R1442 B.n869 B.n868 10.6151
R1443 B.n869 B.n404 10.6151
R1444 B.n879 B.n404 10.6151
R1445 B.n880 B.n879 10.6151
R1446 B.n882 B.n880 10.6151
R1447 B.n882 B.n881 10.6151
R1448 B.n881 B.n396 10.6151
R1449 B.n893 B.n396 10.6151
R1450 B.n894 B.n893 10.6151
R1451 B.n895 B.n894 10.6151
R1452 B.n896 B.n895 10.6151
R1453 B.n898 B.n896 10.6151
R1454 B.n899 B.n898 10.6151
R1455 B.n900 B.n899 10.6151
R1456 B.n901 B.n900 10.6151
R1457 B.n903 B.n901 10.6151
R1458 B.n904 B.n903 10.6151
R1459 B.n905 B.n904 10.6151
R1460 B.n906 B.n905 10.6151
R1461 B.n908 B.n906 10.6151
R1462 B.n909 B.n908 10.6151
R1463 B.n910 B.n909 10.6151
R1464 B.n911 B.n910 10.6151
R1465 B.n913 B.n911 10.6151
R1466 B.n914 B.n913 10.6151
R1467 B.n915 B.n914 10.6151
R1468 B.n916 B.n915 10.6151
R1469 B.n918 B.n916 10.6151
R1470 B.n919 B.n918 10.6151
R1471 B.n920 B.n919 10.6151
R1472 B.n921 B.n920 10.6151
R1473 B.n923 B.n921 10.6151
R1474 B.n924 B.n923 10.6151
R1475 B.n925 B.n924 10.6151
R1476 B.n926 B.n925 10.6151
R1477 B.n928 B.n926 10.6151
R1478 B.n929 B.n928 10.6151
R1479 B.n930 B.n929 10.6151
R1480 B.n931 B.n930 10.6151
R1481 B.n933 B.n931 10.6151
R1482 B.n934 B.n933 10.6151
R1483 B.n935 B.n934 10.6151
R1484 B.n790 B.n789 10.6151
R1485 B.n789 B.n788 10.6151
R1486 B.n788 B.n787 10.6151
R1487 B.n787 B.n785 10.6151
R1488 B.n785 B.n782 10.6151
R1489 B.n782 B.n781 10.6151
R1490 B.n781 B.n778 10.6151
R1491 B.n778 B.n777 10.6151
R1492 B.n777 B.n774 10.6151
R1493 B.n774 B.n773 10.6151
R1494 B.n773 B.n770 10.6151
R1495 B.n770 B.n769 10.6151
R1496 B.n769 B.n766 10.6151
R1497 B.n766 B.n765 10.6151
R1498 B.n765 B.n762 10.6151
R1499 B.n762 B.n761 10.6151
R1500 B.n761 B.n758 10.6151
R1501 B.n758 B.n757 10.6151
R1502 B.n757 B.n754 10.6151
R1503 B.n754 B.n753 10.6151
R1504 B.n753 B.n750 10.6151
R1505 B.n750 B.n749 10.6151
R1506 B.n749 B.n746 10.6151
R1507 B.n746 B.n745 10.6151
R1508 B.n745 B.n742 10.6151
R1509 B.n742 B.n741 10.6151
R1510 B.n741 B.n738 10.6151
R1511 B.n738 B.n737 10.6151
R1512 B.n737 B.n734 10.6151
R1513 B.n734 B.n733 10.6151
R1514 B.n733 B.n730 10.6151
R1515 B.n730 B.n729 10.6151
R1516 B.n729 B.n726 10.6151
R1517 B.n726 B.n725 10.6151
R1518 B.n725 B.n722 10.6151
R1519 B.n722 B.n721 10.6151
R1520 B.n721 B.n718 10.6151
R1521 B.n718 B.n717 10.6151
R1522 B.n717 B.n714 10.6151
R1523 B.n714 B.n713 10.6151
R1524 B.n713 B.n710 10.6151
R1525 B.n710 B.n709 10.6151
R1526 B.n709 B.n706 10.6151
R1527 B.n706 B.n705 10.6151
R1528 B.n705 B.n702 10.6151
R1529 B.n702 B.n701 10.6151
R1530 B.n701 B.n698 10.6151
R1531 B.n698 B.n697 10.6151
R1532 B.n697 B.n694 10.6151
R1533 B.n694 B.n693 10.6151
R1534 B.n693 B.n690 10.6151
R1535 B.n690 B.n689 10.6151
R1536 B.n689 B.n686 10.6151
R1537 B.n686 B.n685 10.6151
R1538 B.n685 B.n682 10.6151
R1539 B.n682 B.n681 10.6151
R1540 B.n681 B.n678 10.6151
R1541 B.n678 B.n677 10.6151
R1542 B.n677 B.n674 10.6151
R1543 B.n674 B.n673 10.6151
R1544 B.n670 B.n669 10.6151
R1545 B.n669 B.n666 10.6151
R1546 B.n666 B.n665 10.6151
R1547 B.n665 B.n662 10.6151
R1548 B.n662 B.n661 10.6151
R1549 B.n661 B.n658 10.6151
R1550 B.n658 B.n657 10.6151
R1551 B.n657 B.n654 10.6151
R1552 B.n654 B.n653 10.6151
R1553 B.n650 B.n649 10.6151
R1554 B.n649 B.n646 10.6151
R1555 B.n646 B.n645 10.6151
R1556 B.n645 B.n642 10.6151
R1557 B.n642 B.n641 10.6151
R1558 B.n641 B.n638 10.6151
R1559 B.n638 B.n637 10.6151
R1560 B.n637 B.n634 10.6151
R1561 B.n634 B.n633 10.6151
R1562 B.n633 B.n630 10.6151
R1563 B.n630 B.n629 10.6151
R1564 B.n629 B.n626 10.6151
R1565 B.n626 B.n625 10.6151
R1566 B.n625 B.n622 10.6151
R1567 B.n622 B.n621 10.6151
R1568 B.n621 B.n618 10.6151
R1569 B.n618 B.n617 10.6151
R1570 B.n617 B.n614 10.6151
R1571 B.n614 B.n613 10.6151
R1572 B.n613 B.n610 10.6151
R1573 B.n610 B.n609 10.6151
R1574 B.n609 B.n606 10.6151
R1575 B.n606 B.n605 10.6151
R1576 B.n605 B.n602 10.6151
R1577 B.n602 B.n601 10.6151
R1578 B.n601 B.n598 10.6151
R1579 B.n598 B.n597 10.6151
R1580 B.n597 B.n594 10.6151
R1581 B.n594 B.n593 10.6151
R1582 B.n593 B.n590 10.6151
R1583 B.n590 B.n589 10.6151
R1584 B.n589 B.n586 10.6151
R1585 B.n586 B.n585 10.6151
R1586 B.n585 B.n582 10.6151
R1587 B.n582 B.n581 10.6151
R1588 B.n581 B.n578 10.6151
R1589 B.n578 B.n577 10.6151
R1590 B.n577 B.n574 10.6151
R1591 B.n574 B.n573 10.6151
R1592 B.n573 B.n570 10.6151
R1593 B.n570 B.n569 10.6151
R1594 B.n569 B.n566 10.6151
R1595 B.n566 B.n565 10.6151
R1596 B.n565 B.n562 10.6151
R1597 B.n562 B.n561 10.6151
R1598 B.n561 B.n558 10.6151
R1599 B.n558 B.n557 10.6151
R1600 B.n557 B.n554 10.6151
R1601 B.n554 B.n553 10.6151
R1602 B.n553 B.n550 10.6151
R1603 B.n550 B.n549 10.6151
R1604 B.n549 B.n546 10.6151
R1605 B.n546 B.n545 10.6151
R1606 B.n545 B.n542 10.6151
R1607 B.n542 B.n541 10.6151
R1608 B.n541 B.n538 10.6151
R1609 B.n538 B.n537 10.6151
R1610 B.n537 B.n534 10.6151
R1611 B.n534 B.n460 10.6151
R1612 B.n795 B.n460 10.6151
R1613 B.n801 B.n456 10.6151
R1614 B.n802 B.n801 10.6151
R1615 B.n803 B.n802 10.6151
R1616 B.n803 B.n448 10.6151
R1617 B.n813 B.n448 10.6151
R1618 B.n814 B.n813 10.6151
R1619 B.n815 B.n814 10.6151
R1620 B.n815 B.n440 10.6151
R1621 B.n825 B.n440 10.6151
R1622 B.n826 B.n825 10.6151
R1623 B.n827 B.n826 10.6151
R1624 B.n827 B.n432 10.6151
R1625 B.n837 B.n432 10.6151
R1626 B.n838 B.n837 10.6151
R1627 B.n839 B.n838 10.6151
R1628 B.n839 B.n424 10.6151
R1629 B.n849 B.n424 10.6151
R1630 B.n850 B.n849 10.6151
R1631 B.n851 B.n850 10.6151
R1632 B.n851 B.n416 10.6151
R1633 B.n861 B.n416 10.6151
R1634 B.n862 B.n861 10.6151
R1635 B.n863 B.n862 10.6151
R1636 B.n863 B.n408 10.6151
R1637 B.n873 B.n408 10.6151
R1638 B.n874 B.n873 10.6151
R1639 B.n875 B.n874 10.6151
R1640 B.n875 B.n400 10.6151
R1641 B.n886 B.n400 10.6151
R1642 B.n887 B.n886 10.6151
R1643 B.n888 B.n887 10.6151
R1644 B.n888 B.n0 10.6151
R1645 B.n1001 B.n1 10.6151
R1646 B.n1001 B.n1000 10.6151
R1647 B.n1000 B.n999 10.6151
R1648 B.n999 B.n10 10.6151
R1649 B.n993 B.n10 10.6151
R1650 B.n993 B.n992 10.6151
R1651 B.n992 B.n991 10.6151
R1652 B.n991 B.n17 10.6151
R1653 B.n985 B.n17 10.6151
R1654 B.n985 B.n984 10.6151
R1655 B.n984 B.n983 10.6151
R1656 B.n983 B.n24 10.6151
R1657 B.n977 B.n24 10.6151
R1658 B.n977 B.n976 10.6151
R1659 B.n976 B.n975 10.6151
R1660 B.n975 B.n31 10.6151
R1661 B.n969 B.n31 10.6151
R1662 B.n969 B.n968 10.6151
R1663 B.n968 B.n967 10.6151
R1664 B.n967 B.n38 10.6151
R1665 B.n961 B.n38 10.6151
R1666 B.n961 B.n960 10.6151
R1667 B.n960 B.n959 10.6151
R1668 B.n959 B.n45 10.6151
R1669 B.n953 B.n45 10.6151
R1670 B.n953 B.n952 10.6151
R1671 B.n952 B.n951 10.6151
R1672 B.n951 B.n52 10.6151
R1673 B.n945 B.n52 10.6151
R1674 B.n945 B.n944 10.6151
R1675 B.n944 B.n943 10.6151
R1676 B.n943 B.n59 10.6151
R1677 B.n255 B.n254 9.36635
R1678 B.n277 B.n276 9.36635
R1679 B.n673 B.n530 9.36635
R1680 B.n650 B.n533 9.36635
R1681 B.n877 B.t3 8.75076
R1682 B.t0 B.n995 8.75076
R1683 B.n1007 B.n0 2.81026
R1684 B.n1007 B.n1 2.81026
R1685 B.n853 B.t2 1.38212
R1686 B.t1 B.n979 1.38212
R1687 B.n256 B.n255 1.24928
R1688 B.n276 B.n275 1.24928
R1689 B.n670 B.n530 1.24928
R1690 B.n653 B.n533 1.24928
R1691 VP.n4 VP.t3 216.762
R1692 VP.n4 VP.t2 216.01
R1693 VP.n3 VP.t0 181.579
R1694 VP.n15 VP.t1 181.579
R1695 VP.n14 VP.n0 161.3
R1696 VP.n13 VP.n12 161.3
R1697 VP.n11 VP.n1 161.3
R1698 VP.n10 VP.n9 161.3
R1699 VP.n8 VP.n2 161.3
R1700 VP.n7 VP.n6 161.3
R1701 VP.n5 VP.n3 103.416
R1702 VP.n16 VP.n15 103.416
R1703 VP.n9 VP.n1 56.5193
R1704 VP.n5 VP.n4 55.4351
R1705 VP.n8 VP.n7 24.4675
R1706 VP.n9 VP.n8 24.4675
R1707 VP.n13 VP.n1 24.4675
R1708 VP.n14 VP.n13 24.4675
R1709 VP.n7 VP.n3 7.3406
R1710 VP.n15 VP.n14 7.3406
R1711 VP.n6 VP.n5 0.278367
R1712 VP.n16 VP.n0 0.278367
R1713 VP.n6 VP.n2 0.189894
R1714 VP.n10 VP.n2 0.189894
R1715 VP.n11 VP.n10 0.189894
R1716 VP.n12 VP.n11 0.189894
R1717 VP.n12 VP.n0 0.189894
R1718 VP VP.n16 0.153454
R1719 VDD1 VDD1.n1 108.352
R1720 VDD1 VDD1.n0 60.886
R1721 VDD1.n0 VDD1.t3 1.06444
R1722 VDD1.n0 VDD1.t0 1.06444
R1723 VDD1.n1 VDD1.t2 1.06444
R1724 VDD1.n1 VDD1.t1 1.06444
R1725 VTAIL.n5 VTAIL.t4 45.2131
R1726 VTAIL.n4 VTAIL.t3 45.2131
R1727 VTAIL.n3 VTAIL.t1 45.2131
R1728 VTAIL.n7 VTAIL.t0 45.213
R1729 VTAIL.n0 VTAIL.t2 45.213
R1730 VTAIL.n1 VTAIL.t6 45.213
R1731 VTAIL.n2 VTAIL.t7 45.213
R1732 VTAIL.n6 VTAIL.t5 45.213
R1733 VTAIL.n7 VTAIL.n6 30.8238
R1734 VTAIL.n3 VTAIL.n2 30.8238
R1735 VTAIL.n4 VTAIL.n3 2.41429
R1736 VTAIL.n6 VTAIL.n5 2.41429
R1737 VTAIL.n2 VTAIL.n1 2.41429
R1738 VTAIL VTAIL.n0 1.26559
R1739 VTAIL VTAIL.n7 1.14921
R1740 VTAIL.n5 VTAIL.n4 0.470328
R1741 VTAIL.n1 VTAIL.n0 0.470328
R1742 VN.n0 VN.t1 216.762
R1743 VN.n1 VN.t0 216.762
R1744 VN.n0 VN.t2 216.01
R1745 VN.n1 VN.t3 216.01
R1746 VN VN.n1 55.714
R1747 VN VN.n0 4.58899
R1748 VDD2.n2 VDD2.n0 107.828
R1749 VDD2.n2 VDD2.n1 60.8278
R1750 VDD2.n1 VDD2.t0 1.06444
R1751 VDD2.n1 VDD2.t3 1.06444
R1752 VDD2.n0 VDD2.t2 1.06444
R1753 VDD2.n0 VDD2.t1 1.06444
R1754 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 6.99317f
C1 VDD1 VN 0.149016f
C2 VTAIL VN 6.72613f
C3 VDD2 VDD1 1.00199f
C4 VP VDD1 7.35892f
C5 VDD2 VTAIL 7.04651f
C6 VDD2 VN 7.12248f
C7 VP VTAIL 6.74023f
C8 VP VN 7.32389f
C9 VDD2 VP 0.386166f
C10 VDD2 B 4.201078f
C11 VDD1 B 8.97934f
C12 VTAIL B 13.966022f
C13 VN B 11.022519f
C14 VP B 9.107763f
C15 VDD2.t2 B 0.387068f
C16 VDD2.t1 B 0.387068f
C17 VDD2.n0 B 4.4351f
C18 VDD2.t0 B 0.387068f
C19 VDD2.t3 B 0.387068f
C20 VDD2.n1 B 3.53064f
C21 VDD2.n2 B 4.37561f
C22 VN.t1 B 3.35303f
C23 VN.t2 B 3.34875f
C24 VN.n0 B 2.18708f
C25 VN.t0 B 3.35303f
C26 VN.t3 B 3.34875f
C27 VN.n1 B 3.70338f
C28 VTAIL.t2 B 2.53509f
C29 VTAIL.n0 B 0.292474f
C30 VTAIL.t6 B 2.53509f
C31 VTAIL.n1 B 0.348497f
C32 VTAIL.t7 B 2.53509f
C33 VTAIL.n2 B 1.43133f
C34 VTAIL.t1 B 2.5351f
C35 VTAIL.n3 B 1.43132f
C36 VTAIL.t3 B 2.5351f
C37 VTAIL.n4 B 0.348482f
C38 VTAIL.t4 B 2.5351f
C39 VTAIL.n5 B 0.348482f
C40 VTAIL.t5 B 2.53509f
C41 VTAIL.n6 B 1.43133f
C42 VTAIL.t0 B 2.53509f
C43 VTAIL.n7 B 1.36963f
C44 VDD1.t3 B 0.392597f
C45 VDD1.t0 B 0.392597f
C46 VDD1.n0 B 3.58149f
C47 VDD1.t2 B 0.392597f
C48 VDD1.t1 B 0.392597f
C49 VDD1.n1 B 4.52722f
C50 VP.n0 B 0.033356f
C51 VP.t1 B 3.20083f
C52 VP.n1 B 0.036934f
C53 VP.n2 B 0.0253f
C54 VP.t0 B 3.20083f
C55 VP.n3 B 1.18647f
C56 VP.t2 B 3.40201f
C57 VP.t3 B 3.40636f
C58 VP.n4 B 3.74913f
C59 VP.n5 B 1.60024f
C60 VP.n6 B 0.033356f
C61 VP.n7 B 0.030858f
C62 VP.n8 B 0.047154f
C63 VP.n9 B 0.036934f
C64 VP.n10 B 0.0253f
C65 VP.n11 B 0.0253f
C66 VP.n12 B 0.0253f
C67 VP.n13 B 0.047154f
C68 VP.n14 B 0.030858f
C69 VP.n15 B 1.18647f
C70 VP.n16 B 0.041671f
.ends

