* NGSPICE file created from diff_pair_sample_1244.ext - technology: sky130A

.subckt diff_pair_sample_1244 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=0 ps=0 w=16.67 l=0.24
X1 VTAIL.t9 VN.t0 VDD2.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=2.75055 ps=17 w=16.67 l=0.24
X2 VTAIL.t10 VP.t0 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=2.75055 ps=17 w=16.67 l=0.24
X3 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=0 ps=0 w=16.67 l=0.24
X4 VTAIL.t11 VP.t1 VDD1.t4 B.t19 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=2.75055 ps=17 w=16.67 l=0.24
X5 VDD1.t3 VP.t2 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=2.75055 ps=17 w=16.67 l=0.24
X6 VDD1.t2 VP.t3 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=6.5013 ps=34.12 w=16.67 l=0.24
X7 VDD2.t3 VN.t1 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=2.75055 ps=17 w=16.67 l=0.24
X8 VDD2.t1 VN.t2 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=6.5013 ps=34.12 w=16.67 l=0.24
X9 VDD2.t0 VN.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=6.5013 ps=34.12 w=16.67 l=0.24
X10 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=6.5013 ps=34.12 w=16.67 l=0.24
X11 VTAIL.t5 VN.t4 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.75055 pd=17 as=2.75055 ps=17 w=16.67 l=0.24
X12 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=0 ps=0 w=16.67 l=0.24
X13 VDD1.t0 VP.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=2.75055 ps=17 w=16.67 l=0.24
X14 VDD2.t5 VN.t5 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=2.75055 ps=17 w=16.67 l=0.24
X15 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=6.5013 pd=34.12 as=0 ps=0 w=16.67 l=0.24
R0 B.n423 B.t16 1900.25
R1 B.n420 B.t9 1900.25
R2 B.n95 B.t13 1900.25
R3 B.n93 B.t5 1900.25
R4 B.n730 B.n729 585
R5 B.n331 B.n91 585
R6 B.n330 B.n329 585
R7 B.n328 B.n327 585
R8 B.n326 B.n325 585
R9 B.n324 B.n323 585
R10 B.n322 B.n321 585
R11 B.n320 B.n319 585
R12 B.n318 B.n317 585
R13 B.n316 B.n315 585
R14 B.n314 B.n313 585
R15 B.n312 B.n311 585
R16 B.n310 B.n309 585
R17 B.n308 B.n307 585
R18 B.n306 B.n305 585
R19 B.n304 B.n303 585
R20 B.n302 B.n301 585
R21 B.n300 B.n299 585
R22 B.n298 B.n297 585
R23 B.n296 B.n295 585
R24 B.n294 B.n293 585
R25 B.n292 B.n291 585
R26 B.n290 B.n289 585
R27 B.n288 B.n287 585
R28 B.n286 B.n285 585
R29 B.n284 B.n283 585
R30 B.n282 B.n281 585
R31 B.n280 B.n279 585
R32 B.n278 B.n277 585
R33 B.n276 B.n275 585
R34 B.n274 B.n273 585
R35 B.n272 B.n271 585
R36 B.n270 B.n269 585
R37 B.n268 B.n267 585
R38 B.n266 B.n265 585
R39 B.n264 B.n263 585
R40 B.n262 B.n261 585
R41 B.n260 B.n259 585
R42 B.n258 B.n257 585
R43 B.n256 B.n255 585
R44 B.n254 B.n253 585
R45 B.n252 B.n251 585
R46 B.n250 B.n249 585
R47 B.n248 B.n247 585
R48 B.n246 B.n245 585
R49 B.n244 B.n243 585
R50 B.n242 B.n241 585
R51 B.n240 B.n239 585
R52 B.n238 B.n237 585
R53 B.n236 B.n235 585
R54 B.n234 B.n233 585
R55 B.n232 B.n231 585
R56 B.n230 B.n229 585
R57 B.n228 B.n227 585
R58 B.n226 B.n225 585
R59 B.n223 B.n222 585
R60 B.n221 B.n220 585
R61 B.n219 B.n218 585
R62 B.n217 B.n216 585
R63 B.n215 B.n214 585
R64 B.n213 B.n212 585
R65 B.n211 B.n210 585
R66 B.n209 B.n208 585
R67 B.n207 B.n206 585
R68 B.n205 B.n204 585
R69 B.n202 B.n201 585
R70 B.n200 B.n199 585
R71 B.n198 B.n197 585
R72 B.n196 B.n195 585
R73 B.n194 B.n193 585
R74 B.n192 B.n191 585
R75 B.n190 B.n189 585
R76 B.n188 B.n187 585
R77 B.n186 B.n185 585
R78 B.n184 B.n183 585
R79 B.n182 B.n181 585
R80 B.n180 B.n179 585
R81 B.n178 B.n177 585
R82 B.n176 B.n175 585
R83 B.n174 B.n173 585
R84 B.n172 B.n171 585
R85 B.n170 B.n169 585
R86 B.n168 B.n167 585
R87 B.n166 B.n165 585
R88 B.n164 B.n163 585
R89 B.n162 B.n161 585
R90 B.n160 B.n159 585
R91 B.n158 B.n157 585
R92 B.n156 B.n155 585
R93 B.n154 B.n153 585
R94 B.n152 B.n151 585
R95 B.n150 B.n149 585
R96 B.n148 B.n147 585
R97 B.n146 B.n145 585
R98 B.n144 B.n143 585
R99 B.n142 B.n141 585
R100 B.n140 B.n139 585
R101 B.n138 B.n137 585
R102 B.n136 B.n135 585
R103 B.n134 B.n133 585
R104 B.n132 B.n131 585
R105 B.n130 B.n129 585
R106 B.n128 B.n127 585
R107 B.n126 B.n125 585
R108 B.n124 B.n123 585
R109 B.n122 B.n121 585
R110 B.n120 B.n119 585
R111 B.n118 B.n117 585
R112 B.n116 B.n115 585
R113 B.n114 B.n113 585
R114 B.n112 B.n111 585
R115 B.n110 B.n109 585
R116 B.n108 B.n107 585
R117 B.n106 B.n105 585
R118 B.n104 B.n103 585
R119 B.n102 B.n101 585
R120 B.n100 B.n99 585
R121 B.n98 B.n97 585
R122 B.n32 B.n31 585
R123 B.n735 B.n734 585
R124 B.n728 B.n92 585
R125 B.n92 B.n29 585
R126 B.n727 B.n28 585
R127 B.n739 B.n28 585
R128 B.n726 B.n27 585
R129 B.n740 B.n27 585
R130 B.n725 B.n26 585
R131 B.n741 B.n26 585
R132 B.n724 B.n723 585
R133 B.n723 B.n25 585
R134 B.n722 B.n21 585
R135 B.n747 B.n21 585
R136 B.n721 B.n20 585
R137 B.n748 B.n20 585
R138 B.n720 B.n19 585
R139 B.n749 B.n19 585
R140 B.n719 B.n718 585
R141 B.n718 B.n15 585
R142 B.n717 B.n14 585
R143 B.n755 B.n14 585
R144 B.n716 B.n13 585
R145 B.n756 B.n13 585
R146 B.n715 B.n12 585
R147 B.n757 B.n12 585
R148 B.n714 B.n713 585
R149 B.n713 B.n11 585
R150 B.n712 B.n7 585
R151 B.n763 B.n7 585
R152 B.n711 B.n6 585
R153 B.n764 B.n6 585
R154 B.n710 B.n5 585
R155 B.n765 B.n5 585
R156 B.n709 B.n708 585
R157 B.n708 B.n4 585
R158 B.n707 B.n332 585
R159 B.n707 B.n706 585
R160 B.n696 B.n333 585
R161 B.n699 B.n333 585
R162 B.n698 B.n697 585
R163 B.n700 B.n698 585
R164 B.n695 B.n337 585
R165 B.n341 B.n337 585
R166 B.n694 B.n693 585
R167 B.n693 B.n692 585
R168 B.n339 B.n338 585
R169 B.n340 B.n339 585
R170 B.n685 B.n684 585
R171 B.n686 B.n685 585
R172 B.n683 B.n346 585
R173 B.n346 B.n345 585
R174 B.n682 B.n681 585
R175 B.n681 B.n680 585
R176 B.n348 B.n347 585
R177 B.n673 B.n348 585
R178 B.n672 B.n671 585
R179 B.n674 B.n672 585
R180 B.n670 B.n353 585
R181 B.n353 B.n352 585
R182 B.n669 B.n668 585
R183 B.n668 B.n667 585
R184 B.n355 B.n354 585
R185 B.n356 B.n355 585
R186 B.n663 B.n662 585
R187 B.n359 B.n358 585
R188 B.n659 B.n658 585
R189 B.n660 B.n659 585
R190 B.n657 B.n419 585
R191 B.n656 B.n655 585
R192 B.n654 B.n653 585
R193 B.n652 B.n651 585
R194 B.n650 B.n649 585
R195 B.n648 B.n647 585
R196 B.n646 B.n645 585
R197 B.n644 B.n643 585
R198 B.n642 B.n641 585
R199 B.n640 B.n639 585
R200 B.n638 B.n637 585
R201 B.n636 B.n635 585
R202 B.n634 B.n633 585
R203 B.n632 B.n631 585
R204 B.n630 B.n629 585
R205 B.n628 B.n627 585
R206 B.n626 B.n625 585
R207 B.n624 B.n623 585
R208 B.n622 B.n621 585
R209 B.n620 B.n619 585
R210 B.n618 B.n617 585
R211 B.n616 B.n615 585
R212 B.n614 B.n613 585
R213 B.n612 B.n611 585
R214 B.n610 B.n609 585
R215 B.n608 B.n607 585
R216 B.n606 B.n605 585
R217 B.n604 B.n603 585
R218 B.n602 B.n601 585
R219 B.n600 B.n599 585
R220 B.n598 B.n597 585
R221 B.n596 B.n595 585
R222 B.n594 B.n593 585
R223 B.n592 B.n591 585
R224 B.n590 B.n589 585
R225 B.n588 B.n587 585
R226 B.n586 B.n585 585
R227 B.n584 B.n583 585
R228 B.n582 B.n581 585
R229 B.n580 B.n579 585
R230 B.n578 B.n577 585
R231 B.n576 B.n575 585
R232 B.n574 B.n573 585
R233 B.n572 B.n571 585
R234 B.n570 B.n569 585
R235 B.n568 B.n567 585
R236 B.n566 B.n565 585
R237 B.n564 B.n563 585
R238 B.n562 B.n561 585
R239 B.n560 B.n559 585
R240 B.n558 B.n557 585
R241 B.n556 B.n555 585
R242 B.n554 B.n553 585
R243 B.n552 B.n551 585
R244 B.n550 B.n549 585
R245 B.n548 B.n547 585
R246 B.n546 B.n545 585
R247 B.n544 B.n543 585
R248 B.n542 B.n541 585
R249 B.n540 B.n539 585
R250 B.n538 B.n537 585
R251 B.n536 B.n535 585
R252 B.n534 B.n533 585
R253 B.n532 B.n531 585
R254 B.n530 B.n529 585
R255 B.n528 B.n527 585
R256 B.n526 B.n525 585
R257 B.n524 B.n523 585
R258 B.n522 B.n521 585
R259 B.n520 B.n519 585
R260 B.n518 B.n517 585
R261 B.n516 B.n515 585
R262 B.n514 B.n513 585
R263 B.n512 B.n511 585
R264 B.n510 B.n509 585
R265 B.n508 B.n507 585
R266 B.n506 B.n505 585
R267 B.n504 B.n503 585
R268 B.n502 B.n501 585
R269 B.n500 B.n499 585
R270 B.n498 B.n497 585
R271 B.n496 B.n495 585
R272 B.n494 B.n493 585
R273 B.n492 B.n491 585
R274 B.n490 B.n489 585
R275 B.n488 B.n487 585
R276 B.n486 B.n485 585
R277 B.n484 B.n483 585
R278 B.n482 B.n481 585
R279 B.n480 B.n479 585
R280 B.n478 B.n477 585
R281 B.n476 B.n475 585
R282 B.n474 B.n473 585
R283 B.n472 B.n471 585
R284 B.n470 B.n469 585
R285 B.n468 B.n467 585
R286 B.n466 B.n465 585
R287 B.n464 B.n463 585
R288 B.n462 B.n461 585
R289 B.n460 B.n459 585
R290 B.n458 B.n457 585
R291 B.n456 B.n455 585
R292 B.n454 B.n453 585
R293 B.n452 B.n451 585
R294 B.n450 B.n449 585
R295 B.n448 B.n447 585
R296 B.n446 B.n445 585
R297 B.n444 B.n443 585
R298 B.n442 B.n441 585
R299 B.n440 B.n439 585
R300 B.n438 B.n437 585
R301 B.n436 B.n435 585
R302 B.n434 B.n433 585
R303 B.n432 B.n431 585
R304 B.n430 B.n429 585
R305 B.n428 B.n427 585
R306 B.n426 B.n418 585
R307 B.n660 B.n418 585
R308 B.n664 B.n357 585
R309 B.n357 B.n356 585
R310 B.n666 B.n665 585
R311 B.n667 B.n666 585
R312 B.n351 B.n350 585
R313 B.n352 B.n351 585
R314 B.n676 B.n675 585
R315 B.n675 B.n674 585
R316 B.n677 B.n349 585
R317 B.n673 B.n349 585
R318 B.n679 B.n678 585
R319 B.n680 B.n679 585
R320 B.n344 B.n343 585
R321 B.n345 B.n344 585
R322 B.n688 B.n687 585
R323 B.n687 B.n686 585
R324 B.n689 B.n342 585
R325 B.n342 B.n340 585
R326 B.n691 B.n690 585
R327 B.n692 B.n691 585
R328 B.n336 B.n335 585
R329 B.n341 B.n336 585
R330 B.n702 B.n701 585
R331 B.n701 B.n700 585
R332 B.n703 B.n334 585
R333 B.n699 B.n334 585
R334 B.n705 B.n704 585
R335 B.n706 B.n705 585
R336 B.n2 B.n0 585
R337 B.n4 B.n2 585
R338 B.n3 B.n1 585
R339 B.n764 B.n3 585
R340 B.n762 B.n761 585
R341 B.n763 B.n762 585
R342 B.n760 B.n8 585
R343 B.n11 B.n8 585
R344 B.n759 B.n758 585
R345 B.n758 B.n757 585
R346 B.n10 B.n9 585
R347 B.n756 B.n10 585
R348 B.n754 B.n753 585
R349 B.n755 B.n754 585
R350 B.n752 B.n16 585
R351 B.n16 B.n15 585
R352 B.n751 B.n750 585
R353 B.n750 B.n749 585
R354 B.n18 B.n17 585
R355 B.n748 B.n18 585
R356 B.n746 B.n745 585
R357 B.n747 B.n746 585
R358 B.n744 B.n22 585
R359 B.n25 B.n22 585
R360 B.n743 B.n742 585
R361 B.n742 B.n741 585
R362 B.n24 B.n23 585
R363 B.n740 B.n24 585
R364 B.n738 B.n737 585
R365 B.n739 B.n738 585
R366 B.n736 B.n30 585
R367 B.n30 B.n29 585
R368 B.n767 B.n766 585
R369 B.n766 B.n765 585
R370 B.n662 B.n357 492.5
R371 B.n734 B.n30 492.5
R372 B.n418 B.n355 492.5
R373 B.n730 B.n92 492.5
R374 B.n423 B.t18 373.305
R375 B.n93 B.t7 373.305
R376 B.n420 B.t12 373.305
R377 B.n95 B.t14 373.305
R378 B.n424 B.t17 362.25
R379 B.n94 B.t8 362.25
R380 B.n421 B.t11 362.25
R381 B.n96 B.t15 362.25
R382 B.n732 B.n731 256.663
R383 B.n732 B.n90 256.663
R384 B.n732 B.n89 256.663
R385 B.n732 B.n88 256.663
R386 B.n732 B.n87 256.663
R387 B.n732 B.n86 256.663
R388 B.n732 B.n85 256.663
R389 B.n732 B.n84 256.663
R390 B.n732 B.n83 256.663
R391 B.n732 B.n82 256.663
R392 B.n732 B.n81 256.663
R393 B.n732 B.n80 256.663
R394 B.n732 B.n79 256.663
R395 B.n732 B.n78 256.663
R396 B.n732 B.n77 256.663
R397 B.n732 B.n76 256.663
R398 B.n732 B.n75 256.663
R399 B.n732 B.n74 256.663
R400 B.n732 B.n73 256.663
R401 B.n732 B.n72 256.663
R402 B.n732 B.n71 256.663
R403 B.n732 B.n70 256.663
R404 B.n732 B.n69 256.663
R405 B.n732 B.n68 256.663
R406 B.n732 B.n67 256.663
R407 B.n732 B.n66 256.663
R408 B.n732 B.n65 256.663
R409 B.n732 B.n64 256.663
R410 B.n732 B.n63 256.663
R411 B.n732 B.n62 256.663
R412 B.n732 B.n61 256.663
R413 B.n732 B.n60 256.663
R414 B.n732 B.n59 256.663
R415 B.n732 B.n58 256.663
R416 B.n732 B.n57 256.663
R417 B.n732 B.n56 256.663
R418 B.n732 B.n55 256.663
R419 B.n732 B.n54 256.663
R420 B.n732 B.n53 256.663
R421 B.n732 B.n52 256.663
R422 B.n732 B.n51 256.663
R423 B.n732 B.n50 256.663
R424 B.n732 B.n49 256.663
R425 B.n732 B.n48 256.663
R426 B.n732 B.n47 256.663
R427 B.n732 B.n46 256.663
R428 B.n732 B.n45 256.663
R429 B.n732 B.n44 256.663
R430 B.n732 B.n43 256.663
R431 B.n732 B.n42 256.663
R432 B.n732 B.n41 256.663
R433 B.n732 B.n40 256.663
R434 B.n732 B.n39 256.663
R435 B.n732 B.n38 256.663
R436 B.n732 B.n37 256.663
R437 B.n732 B.n36 256.663
R438 B.n732 B.n35 256.663
R439 B.n732 B.n34 256.663
R440 B.n732 B.n33 256.663
R441 B.n733 B.n732 256.663
R442 B.n661 B.n660 256.663
R443 B.n660 B.n360 256.663
R444 B.n660 B.n361 256.663
R445 B.n660 B.n362 256.663
R446 B.n660 B.n363 256.663
R447 B.n660 B.n364 256.663
R448 B.n660 B.n365 256.663
R449 B.n660 B.n366 256.663
R450 B.n660 B.n367 256.663
R451 B.n660 B.n368 256.663
R452 B.n660 B.n369 256.663
R453 B.n660 B.n370 256.663
R454 B.n660 B.n371 256.663
R455 B.n660 B.n372 256.663
R456 B.n660 B.n373 256.663
R457 B.n660 B.n374 256.663
R458 B.n660 B.n375 256.663
R459 B.n660 B.n376 256.663
R460 B.n660 B.n377 256.663
R461 B.n660 B.n378 256.663
R462 B.n660 B.n379 256.663
R463 B.n660 B.n380 256.663
R464 B.n660 B.n381 256.663
R465 B.n660 B.n382 256.663
R466 B.n660 B.n383 256.663
R467 B.n660 B.n384 256.663
R468 B.n660 B.n385 256.663
R469 B.n660 B.n386 256.663
R470 B.n660 B.n387 256.663
R471 B.n660 B.n388 256.663
R472 B.n660 B.n389 256.663
R473 B.n660 B.n390 256.663
R474 B.n660 B.n391 256.663
R475 B.n660 B.n392 256.663
R476 B.n660 B.n393 256.663
R477 B.n660 B.n394 256.663
R478 B.n660 B.n395 256.663
R479 B.n660 B.n396 256.663
R480 B.n660 B.n397 256.663
R481 B.n660 B.n398 256.663
R482 B.n660 B.n399 256.663
R483 B.n660 B.n400 256.663
R484 B.n660 B.n401 256.663
R485 B.n660 B.n402 256.663
R486 B.n660 B.n403 256.663
R487 B.n660 B.n404 256.663
R488 B.n660 B.n405 256.663
R489 B.n660 B.n406 256.663
R490 B.n660 B.n407 256.663
R491 B.n660 B.n408 256.663
R492 B.n660 B.n409 256.663
R493 B.n660 B.n410 256.663
R494 B.n660 B.n411 256.663
R495 B.n660 B.n412 256.663
R496 B.n660 B.n413 256.663
R497 B.n660 B.n414 256.663
R498 B.n660 B.n415 256.663
R499 B.n660 B.n416 256.663
R500 B.n660 B.n417 256.663
R501 B.n666 B.n357 163.367
R502 B.n666 B.n351 163.367
R503 B.n675 B.n351 163.367
R504 B.n675 B.n349 163.367
R505 B.n679 B.n349 163.367
R506 B.n679 B.n344 163.367
R507 B.n687 B.n344 163.367
R508 B.n687 B.n342 163.367
R509 B.n691 B.n342 163.367
R510 B.n691 B.n336 163.367
R511 B.n701 B.n336 163.367
R512 B.n701 B.n334 163.367
R513 B.n705 B.n334 163.367
R514 B.n705 B.n2 163.367
R515 B.n766 B.n2 163.367
R516 B.n766 B.n3 163.367
R517 B.n762 B.n3 163.367
R518 B.n762 B.n8 163.367
R519 B.n758 B.n8 163.367
R520 B.n758 B.n10 163.367
R521 B.n754 B.n10 163.367
R522 B.n754 B.n16 163.367
R523 B.n750 B.n16 163.367
R524 B.n750 B.n18 163.367
R525 B.n746 B.n18 163.367
R526 B.n746 B.n22 163.367
R527 B.n742 B.n22 163.367
R528 B.n742 B.n24 163.367
R529 B.n738 B.n24 163.367
R530 B.n738 B.n30 163.367
R531 B.n659 B.n359 163.367
R532 B.n659 B.n419 163.367
R533 B.n655 B.n654 163.367
R534 B.n651 B.n650 163.367
R535 B.n647 B.n646 163.367
R536 B.n643 B.n642 163.367
R537 B.n639 B.n638 163.367
R538 B.n635 B.n634 163.367
R539 B.n631 B.n630 163.367
R540 B.n627 B.n626 163.367
R541 B.n623 B.n622 163.367
R542 B.n619 B.n618 163.367
R543 B.n615 B.n614 163.367
R544 B.n611 B.n610 163.367
R545 B.n607 B.n606 163.367
R546 B.n603 B.n602 163.367
R547 B.n599 B.n598 163.367
R548 B.n595 B.n594 163.367
R549 B.n591 B.n590 163.367
R550 B.n587 B.n586 163.367
R551 B.n583 B.n582 163.367
R552 B.n579 B.n578 163.367
R553 B.n575 B.n574 163.367
R554 B.n571 B.n570 163.367
R555 B.n567 B.n566 163.367
R556 B.n563 B.n562 163.367
R557 B.n559 B.n558 163.367
R558 B.n555 B.n554 163.367
R559 B.n551 B.n550 163.367
R560 B.n547 B.n546 163.367
R561 B.n543 B.n542 163.367
R562 B.n539 B.n538 163.367
R563 B.n535 B.n534 163.367
R564 B.n531 B.n530 163.367
R565 B.n527 B.n526 163.367
R566 B.n523 B.n522 163.367
R567 B.n519 B.n518 163.367
R568 B.n515 B.n514 163.367
R569 B.n511 B.n510 163.367
R570 B.n507 B.n506 163.367
R571 B.n503 B.n502 163.367
R572 B.n499 B.n498 163.367
R573 B.n495 B.n494 163.367
R574 B.n491 B.n490 163.367
R575 B.n487 B.n486 163.367
R576 B.n483 B.n482 163.367
R577 B.n479 B.n478 163.367
R578 B.n475 B.n474 163.367
R579 B.n471 B.n470 163.367
R580 B.n467 B.n466 163.367
R581 B.n463 B.n462 163.367
R582 B.n459 B.n458 163.367
R583 B.n455 B.n454 163.367
R584 B.n451 B.n450 163.367
R585 B.n447 B.n446 163.367
R586 B.n443 B.n442 163.367
R587 B.n439 B.n438 163.367
R588 B.n435 B.n434 163.367
R589 B.n431 B.n430 163.367
R590 B.n427 B.n418 163.367
R591 B.n668 B.n355 163.367
R592 B.n668 B.n353 163.367
R593 B.n672 B.n353 163.367
R594 B.n672 B.n348 163.367
R595 B.n681 B.n348 163.367
R596 B.n681 B.n346 163.367
R597 B.n685 B.n346 163.367
R598 B.n685 B.n339 163.367
R599 B.n693 B.n339 163.367
R600 B.n693 B.n337 163.367
R601 B.n698 B.n337 163.367
R602 B.n698 B.n333 163.367
R603 B.n707 B.n333 163.367
R604 B.n708 B.n707 163.367
R605 B.n708 B.n5 163.367
R606 B.n6 B.n5 163.367
R607 B.n7 B.n6 163.367
R608 B.n713 B.n7 163.367
R609 B.n713 B.n12 163.367
R610 B.n13 B.n12 163.367
R611 B.n14 B.n13 163.367
R612 B.n718 B.n14 163.367
R613 B.n718 B.n19 163.367
R614 B.n20 B.n19 163.367
R615 B.n21 B.n20 163.367
R616 B.n723 B.n21 163.367
R617 B.n723 B.n26 163.367
R618 B.n27 B.n26 163.367
R619 B.n28 B.n27 163.367
R620 B.n92 B.n28 163.367
R621 B.n97 B.n32 163.367
R622 B.n101 B.n100 163.367
R623 B.n105 B.n104 163.367
R624 B.n109 B.n108 163.367
R625 B.n113 B.n112 163.367
R626 B.n117 B.n116 163.367
R627 B.n121 B.n120 163.367
R628 B.n125 B.n124 163.367
R629 B.n129 B.n128 163.367
R630 B.n133 B.n132 163.367
R631 B.n137 B.n136 163.367
R632 B.n141 B.n140 163.367
R633 B.n145 B.n144 163.367
R634 B.n149 B.n148 163.367
R635 B.n153 B.n152 163.367
R636 B.n157 B.n156 163.367
R637 B.n161 B.n160 163.367
R638 B.n165 B.n164 163.367
R639 B.n169 B.n168 163.367
R640 B.n173 B.n172 163.367
R641 B.n177 B.n176 163.367
R642 B.n181 B.n180 163.367
R643 B.n185 B.n184 163.367
R644 B.n189 B.n188 163.367
R645 B.n193 B.n192 163.367
R646 B.n197 B.n196 163.367
R647 B.n201 B.n200 163.367
R648 B.n206 B.n205 163.367
R649 B.n210 B.n209 163.367
R650 B.n214 B.n213 163.367
R651 B.n218 B.n217 163.367
R652 B.n222 B.n221 163.367
R653 B.n227 B.n226 163.367
R654 B.n231 B.n230 163.367
R655 B.n235 B.n234 163.367
R656 B.n239 B.n238 163.367
R657 B.n243 B.n242 163.367
R658 B.n247 B.n246 163.367
R659 B.n251 B.n250 163.367
R660 B.n255 B.n254 163.367
R661 B.n259 B.n258 163.367
R662 B.n263 B.n262 163.367
R663 B.n267 B.n266 163.367
R664 B.n271 B.n270 163.367
R665 B.n275 B.n274 163.367
R666 B.n279 B.n278 163.367
R667 B.n283 B.n282 163.367
R668 B.n287 B.n286 163.367
R669 B.n291 B.n290 163.367
R670 B.n295 B.n294 163.367
R671 B.n299 B.n298 163.367
R672 B.n303 B.n302 163.367
R673 B.n307 B.n306 163.367
R674 B.n311 B.n310 163.367
R675 B.n315 B.n314 163.367
R676 B.n319 B.n318 163.367
R677 B.n323 B.n322 163.367
R678 B.n327 B.n326 163.367
R679 B.n329 B.n91 163.367
R680 B.n662 B.n661 71.676
R681 B.n419 B.n360 71.676
R682 B.n654 B.n361 71.676
R683 B.n650 B.n362 71.676
R684 B.n646 B.n363 71.676
R685 B.n642 B.n364 71.676
R686 B.n638 B.n365 71.676
R687 B.n634 B.n366 71.676
R688 B.n630 B.n367 71.676
R689 B.n626 B.n368 71.676
R690 B.n622 B.n369 71.676
R691 B.n618 B.n370 71.676
R692 B.n614 B.n371 71.676
R693 B.n610 B.n372 71.676
R694 B.n606 B.n373 71.676
R695 B.n602 B.n374 71.676
R696 B.n598 B.n375 71.676
R697 B.n594 B.n376 71.676
R698 B.n590 B.n377 71.676
R699 B.n586 B.n378 71.676
R700 B.n582 B.n379 71.676
R701 B.n578 B.n380 71.676
R702 B.n574 B.n381 71.676
R703 B.n570 B.n382 71.676
R704 B.n566 B.n383 71.676
R705 B.n562 B.n384 71.676
R706 B.n558 B.n385 71.676
R707 B.n554 B.n386 71.676
R708 B.n550 B.n387 71.676
R709 B.n546 B.n388 71.676
R710 B.n542 B.n389 71.676
R711 B.n538 B.n390 71.676
R712 B.n534 B.n391 71.676
R713 B.n530 B.n392 71.676
R714 B.n526 B.n393 71.676
R715 B.n522 B.n394 71.676
R716 B.n518 B.n395 71.676
R717 B.n514 B.n396 71.676
R718 B.n510 B.n397 71.676
R719 B.n506 B.n398 71.676
R720 B.n502 B.n399 71.676
R721 B.n498 B.n400 71.676
R722 B.n494 B.n401 71.676
R723 B.n490 B.n402 71.676
R724 B.n486 B.n403 71.676
R725 B.n482 B.n404 71.676
R726 B.n478 B.n405 71.676
R727 B.n474 B.n406 71.676
R728 B.n470 B.n407 71.676
R729 B.n466 B.n408 71.676
R730 B.n462 B.n409 71.676
R731 B.n458 B.n410 71.676
R732 B.n454 B.n411 71.676
R733 B.n450 B.n412 71.676
R734 B.n446 B.n413 71.676
R735 B.n442 B.n414 71.676
R736 B.n438 B.n415 71.676
R737 B.n434 B.n416 71.676
R738 B.n430 B.n417 71.676
R739 B.n734 B.n733 71.676
R740 B.n97 B.n33 71.676
R741 B.n101 B.n34 71.676
R742 B.n105 B.n35 71.676
R743 B.n109 B.n36 71.676
R744 B.n113 B.n37 71.676
R745 B.n117 B.n38 71.676
R746 B.n121 B.n39 71.676
R747 B.n125 B.n40 71.676
R748 B.n129 B.n41 71.676
R749 B.n133 B.n42 71.676
R750 B.n137 B.n43 71.676
R751 B.n141 B.n44 71.676
R752 B.n145 B.n45 71.676
R753 B.n149 B.n46 71.676
R754 B.n153 B.n47 71.676
R755 B.n157 B.n48 71.676
R756 B.n161 B.n49 71.676
R757 B.n165 B.n50 71.676
R758 B.n169 B.n51 71.676
R759 B.n173 B.n52 71.676
R760 B.n177 B.n53 71.676
R761 B.n181 B.n54 71.676
R762 B.n185 B.n55 71.676
R763 B.n189 B.n56 71.676
R764 B.n193 B.n57 71.676
R765 B.n197 B.n58 71.676
R766 B.n201 B.n59 71.676
R767 B.n206 B.n60 71.676
R768 B.n210 B.n61 71.676
R769 B.n214 B.n62 71.676
R770 B.n218 B.n63 71.676
R771 B.n222 B.n64 71.676
R772 B.n227 B.n65 71.676
R773 B.n231 B.n66 71.676
R774 B.n235 B.n67 71.676
R775 B.n239 B.n68 71.676
R776 B.n243 B.n69 71.676
R777 B.n247 B.n70 71.676
R778 B.n251 B.n71 71.676
R779 B.n255 B.n72 71.676
R780 B.n259 B.n73 71.676
R781 B.n263 B.n74 71.676
R782 B.n267 B.n75 71.676
R783 B.n271 B.n76 71.676
R784 B.n275 B.n77 71.676
R785 B.n279 B.n78 71.676
R786 B.n283 B.n79 71.676
R787 B.n287 B.n80 71.676
R788 B.n291 B.n81 71.676
R789 B.n295 B.n82 71.676
R790 B.n299 B.n83 71.676
R791 B.n303 B.n84 71.676
R792 B.n307 B.n85 71.676
R793 B.n311 B.n86 71.676
R794 B.n315 B.n87 71.676
R795 B.n319 B.n88 71.676
R796 B.n323 B.n89 71.676
R797 B.n327 B.n90 71.676
R798 B.n731 B.n91 71.676
R799 B.n731 B.n730 71.676
R800 B.n329 B.n90 71.676
R801 B.n326 B.n89 71.676
R802 B.n322 B.n88 71.676
R803 B.n318 B.n87 71.676
R804 B.n314 B.n86 71.676
R805 B.n310 B.n85 71.676
R806 B.n306 B.n84 71.676
R807 B.n302 B.n83 71.676
R808 B.n298 B.n82 71.676
R809 B.n294 B.n81 71.676
R810 B.n290 B.n80 71.676
R811 B.n286 B.n79 71.676
R812 B.n282 B.n78 71.676
R813 B.n278 B.n77 71.676
R814 B.n274 B.n76 71.676
R815 B.n270 B.n75 71.676
R816 B.n266 B.n74 71.676
R817 B.n262 B.n73 71.676
R818 B.n258 B.n72 71.676
R819 B.n254 B.n71 71.676
R820 B.n250 B.n70 71.676
R821 B.n246 B.n69 71.676
R822 B.n242 B.n68 71.676
R823 B.n238 B.n67 71.676
R824 B.n234 B.n66 71.676
R825 B.n230 B.n65 71.676
R826 B.n226 B.n64 71.676
R827 B.n221 B.n63 71.676
R828 B.n217 B.n62 71.676
R829 B.n213 B.n61 71.676
R830 B.n209 B.n60 71.676
R831 B.n205 B.n59 71.676
R832 B.n200 B.n58 71.676
R833 B.n196 B.n57 71.676
R834 B.n192 B.n56 71.676
R835 B.n188 B.n55 71.676
R836 B.n184 B.n54 71.676
R837 B.n180 B.n53 71.676
R838 B.n176 B.n52 71.676
R839 B.n172 B.n51 71.676
R840 B.n168 B.n50 71.676
R841 B.n164 B.n49 71.676
R842 B.n160 B.n48 71.676
R843 B.n156 B.n47 71.676
R844 B.n152 B.n46 71.676
R845 B.n148 B.n45 71.676
R846 B.n144 B.n44 71.676
R847 B.n140 B.n43 71.676
R848 B.n136 B.n42 71.676
R849 B.n132 B.n41 71.676
R850 B.n128 B.n40 71.676
R851 B.n124 B.n39 71.676
R852 B.n120 B.n38 71.676
R853 B.n116 B.n37 71.676
R854 B.n112 B.n36 71.676
R855 B.n108 B.n35 71.676
R856 B.n104 B.n34 71.676
R857 B.n100 B.n33 71.676
R858 B.n733 B.n32 71.676
R859 B.n661 B.n359 71.676
R860 B.n655 B.n360 71.676
R861 B.n651 B.n361 71.676
R862 B.n647 B.n362 71.676
R863 B.n643 B.n363 71.676
R864 B.n639 B.n364 71.676
R865 B.n635 B.n365 71.676
R866 B.n631 B.n366 71.676
R867 B.n627 B.n367 71.676
R868 B.n623 B.n368 71.676
R869 B.n619 B.n369 71.676
R870 B.n615 B.n370 71.676
R871 B.n611 B.n371 71.676
R872 B.n607 B.n372 71.676
R873 B.n603 B.n373 71.676
R874 B.n599 B.n374 71.676
R875 B.n595 B.n375 71.676
R876 B.n591 B.n376 71.676
R877 B.n587 B.n377 71.676
R878 B.n583 B.n378 71.676
R879 B.n579 B.n379 71.676
R880 B.n575 B.n380 71.676
R881 B.n571 B.n381 71.676
R882 B.n567 B.n382 71.676
R883 B.n563 B.n383 71.676
R884 B.n559 B.n384 71.676
R885 B.n555 B.n385 71.676
R886 B.n551 B.n386 71.676
R887 B.n547 B.n387 71.676
R888 B.n543 B.n388 71.676
R889 B.n539 B.n389 71.676
R890 B.n535 B.n390 71.676
R891 B.n531 B.n391 71.676
R892 B.n527 B.n392 71.676
R893 B.n523 B.n393 71.676
R894 B.n519 B.n394 71.676
R895 B.n515 B.n395 71.676
R896 B.n511 B.n396 71.676
R897 B.n507 B.n397 71.676
R898 B.n503 B.n398 71.676
R899 B.n499 B.n399 71.676
R900 B.n495 B.n400 71.676
R901 B.n491 B.n401 71.676
R902 B.n487 B.n402 71.676
R903 B.n483 B.n403 71.676
R904 B.n479 B.n404 71.676
R905 B.n475 B.n405 71.676
R906 B.n471 B.n406 71.676
R907 B.n467 B.n407 71.676
R908 B.n463 B.n408 71.676
R909 B.n459 B.n409 71.676
R910 B.n455 B.n410 71.676
R911 B.n451 B.n411 71.676
R912 B.n447 B.n412 71.676
R913 B.n443 B.n413 71.676
R914 B.n439 B.n414 71.676
R915 B.n435 B.n415 71.676
R916 B.n431 B.n416 71.676
R917 B.n427 B.n417 71.676
R918 B.n425 B.n424 59.5399
R919 B.n422 B.n421 59.5399
R920 B.n203 B.n96 59.5399
R921 B.n224 B.n94 59.5399
R922 B.n660 B.n356 55.6396
R923 B.n732 B.n29 55.6396
R924 B.n667 B.n356 34.0857
R925 B.n667 B.n352 34.0857
R926 B.n674 B.n352 34.0857
R927 B.n674 B.n673 34.0857
R928 B.n680 B.n345 34.0857
R929 B.n686 B.n345 34.0857
R930 B.n686 B.n340 34.0857
R931 B.n692 B.n340 34.0857
R932 B.n700 B.n699 34.0857
R933 B.n706 B.n4 34.0857
R934 B.n765 B.n4 34.0857
R935 B.n765 B.n764 34.0857
R936 B.n764 B.n763 34.0857
R937 B.n757 B.n11 34.0857
R938 B.n755 B.n15 34.0857
R939 B.n749 B.n15 34.0857
R940 B.n749 B.n748 34.0857
R941 B.n748 B.n747 34.0857
R942 B.n741 B.n25 34.0857
R943 B.n741 B.n740 34.0857
R944 B.n740 B.n739 34.0857
R945 B.n739 B.n29 34.0857
R946 B.n736 B.n735 32.0005
R947 B.n729 B.n728 32.0005
R948 B.n426 B.n354 32.0005
R949 B.n664 B.n663 32.0005
R950 B.n341 B.t0 30.0757
R951 B.t19 B.n756 30.0757
R952 B.t1 B.n341 27.0682
R953 B.n756 B.t4 27.0682
R954 B.n680 B.t10 23.0581
R955 B.n747 B.t6 23.0581
R956 B.n699 B.t3 19.0481
R957 B.n11 B.t2 19.0481
R958 B B.n767 18.0485
R959 B.n706 B.t3 15.0381
R960 B.n763 B.t2 15.0381
R961 B.n424 B.n423 11.055
R962 B.n421 B.n420 11.055
R963 B.n96 B.n95 11.055
R964 B.n94 B.n93 11.055
R965 B.n673 B.t10 11.0281
R966 B.n25 B.t6 11.0281
R967 B.n735 B.n31 10.6151
R968 B.n98 B.n31 10.6151
R969 B.n99 B.n98 10.6151
R970 B.n102 B.n99 10.6151
R971 B.n103 B.n102 10.6151
R972 B.n106 B.n103 10.6151
R973 B.n107 B.n106 10.6151
R974 B.n110 B.n107 10.6151
R975 B.n111 B.n110 10.6151
R976 B.n114 B.n111 10.6151
R977 B.n115 B.n114 10.6151
R978 B.n118 B.n115 10.6151
R979 B.n119 B.n118 10.6151
R980 B.n122 B.n119 10.6151
R981 B.n123 B.n122 10.6151
R982 B.n126 B.n123 10.6151
R983 B.n127 B.n126 10.6151
R984 B.n130 B.n127 10.6151
R985 B.n131 B.n130 10.6151
R986 B.n134 B.n131 10.6151
R987 B.n135 B.n134 10.6151
R988 B.n138 B.n135 10.6151
R989 B.n139 B.n138 10.6151
R990 B.n142 B.n139 10.6151
R991 B.n143 B.n142 10.6151
R992 B.n146 B.n143 10.6151
R993 B.n147 B.n146 10.6151
R994 B.n150 B.n147 10.6151
R995 B.n151 B.n150 10.6151
R996 B.n154 B.n151 10.6151
R997 B.n155 B.n154 10.6151
R998 B.n158 B.n155 10.6151
R999 B.n159 B.n158 10.6151
R1000 B.n162 B.n159 10.6151
R1001 B.n163 B.n162 10.6151
R1002 B.n166 B.n163 10.6151
R1003 B.n167 B.n166 10.6151
R1004 B.n170 B.n167 10.6151
R1005 B.n171 B.n170 10.6151
R1006 B.n174 B.n171 10.6151
R1007 B.n175 B.n174 10.6151
R1008 B.n178 B.n175 10.6151
R1009 B.n179 B.n178 10.6151
R1010 B.n182 B.n179 10.6151
R1011 B.n183 B.n182 10.6151
R1012 B.n186 B.n183 10.6151
R1013 B.n187 B.n186 10.6151
R1014 B.n190 B.n187 10.6151
R1015 B.n191 B.n190 10.6151
R1016 B.n194 B.n191 10.6151
R1017 B.n195 B.n194 10.6151
R1018 B.n198 B.n195 10.6151
R1019 B.n199 B.n198 10.6151
R1020 B.n202 B.n199 10.6151
R1021 B.n207 B.n204 10.6151
R1022 B.n208 B.n207 10.6151
R1023 B.n211 B.n208 10.6151
R1024 B.n212 B.n211 10.6151
R1025 B.n215 B.n212 10.6151
R1026 B.n216 B.n215 10.6151
R1027 B.n219 B.n216 10.6151
R1028 B.n220 B.n219 10.6151
R1029 B.n223 B.n220 10.6151
R1030 B.n228 B.n225 10.6151
R1031 B.n229 B.n228 10.6151
R1032 B.n232 B.n229 10.6151
R1033 B.n233 B.n232 10.6151
R1034 B.n236 B.n233 10.6151
R1035 B.n237 B.n236 10.6151
R1036 B.n240 B.n237 10.6151
R1037 B.n241 B.n240 10.6151
R1038 B.n244 B.n241 10.6151
R1039 B.n245 B.n244 10.6151
R1040 B.n248 B.n245 10.6151
R1041 B.n249 B.n248 10.6151
R1042 B.n252 B.n249 10.6151
R1043 B.n253 B.n252 10.6151
R1044 B.n256 B.n253 10.6151
R1045 B.n257 B.n256 10.6151
R1046 B.n260 B.n257 10.6151
R1047 B.n261 B.n260 10.6151
R1048 B.n264 B.n261 10.6151
R1049 B.n265 B.n264 10.6151
R1050 B.n268 B.n265 10.6151
R1051 B.n269 B.n268 10.6151
R1052 B.n272 B.n269 10.6151
R1053 B.n273 B.n272 10.6151
R1054 B.n276 B.n273 10.6151
R1055 B.n277 B.n276 10.6151
R1056 B.n280 B.n277 10.6151
R1057 B.n281 B.n280 10.6151
R1058 B.n284 B.n281 10.6151
R1059 B.n285 B.n284 10.6151
R1060 B.n288 B.n285 10.6151
R1061 B.n289 B.n288 10.6151
R1062 B.n292 B.n289 10.6151
R1063 B.n293 B.n292 10.6151
R1064 B.n296 B.n293 10.6151
R1065 B.n297 B.n296 10.6151
R1066 B.n300 B.n297 10.6151
R1067 B.n301 B.n300 10.6151
R1068 B.n304 B.n301 10.6151
R1069 B.n305 B.n304 10.6151
R1070 B.n308 B.n305 10.6151
R1071 B.n309 B.n308 10.6151
R1072 B.n312 B.n309 10.6151
R1073 B.n313 B.n312 10.6151
R1074 B.n316 B.n313 10.6151
R1075 B.n317 B.n316 10.6151
R1076 B.n320 B.n317 10.6151
R1077 B.n321 B.n320 10.6151
R1078 B.n324 B.n321 10.6151
R1079 B.n325 B.n324 10.6151
R1080 B.n328 B.n325 10.6151
R1081 B.n330 B.n328 10.6151
R1082 B.n331 B.n330 10.6151
R1083 B.n729 B.n331 10.6151
R1084 B.n669 B.n354 10.6151
R1085 B.n670 B.n669 10.6151
R1086 B.n671 B.n670 10.6151
R1087 B.n671 B.n347 10.6151
R1088 B.n682 B.n347 10.6151
R1089 B.n683 B.n682 10.6151
R1090 B.n684 B.n683 10.6151
R1091 B.n684 B.n338 10.6151
R1092 B.n694 B.n338 10.6151
R1093 B.n695 B.n694 10.6151
R1094 B.n697 B.n695 10.6151
R1095 B.n697 B.n696 10.6151
R1096 B.n696 B.n332 10.6151
R1097 B.n709 B.n332 10.6151
R1098 B.n710 B.n709 10.6151
R1099 B.n711 B.n710 10.6151
R1100 B.n712 B.n711 10.6151
R1101 B.n714 B.n712 10.6151
R1102 B.n715 B.n714 10.6151
R1103 B.n716 B.n715 10.6151
R1104 B.n717 B.n716 10.6151
R1105 B.n719 B.n717 10.6151
R1106 B.n720 B.n719 10.6151
R1107 B.n721 B.n720 10.6151
R1108 B.n722 B.n721 10.6151
R1109 B.n724 B.n722 10.6151
R1110 B.n725 B.n724 10.6151
R1111 B.n726 B.n725 10.6151
R1112 B.n727 B.n726 10.6151
R1113 B.n728 B.n727 10.6151
R1114 B.n663 B.n358 10.6151
R1115 B.n658 B.n358 10.6151
R1116 B.n658 B.n657 10.6151
R1117 B.n657 B.n656 10.6151
R1118 B.n656 B.n653 10.6151
R1119 B.n653 B.n652 10.6151
R1120 B.n652 B.n649 10.6151
R1121 B.n649 B.n648 10.6151
R1122 B.n648 B.n645 10.6151
R1123 B.n645 B.n644 10.6151
R1124 B.n644 B.n641 10.6151
R1125 B.n641 B.n640 10.6151
R1126 B.n640 B.n637 10.6151
R1127 B.n637 B.n636 10.6151
R1128 B.n636 B.n633 10.6151
R1129 B.n633 B.n632 10.6151
R1130 B.n632 B.n629 10.6151
R1131 B.n629 B.n628 10.6151
R1132 B.n628 B.n625 10.6151
R1133 B.n625 B.n624 10.6151
R1134 B.n624 B.n621 10.6151
R1135 B.n621 B.n620 10.6151
R1136 B.n620 B.n617 10.6151
R1137 B.n617 B.n616 10.6151
R1138 B.n616 B.n613 10.6151
R1139 B.n613 B.n612 10.6151
R1140 B.n612 B.n609 10.6151
R1141 B.n609 B.n608 10.6151
R1142 B.n608 B.n605 10.6151
R1143 B.n605 B.n604 10.6151
R1144 B.n604 B.n601 10.6151
R1145 B.n601 B.n600 10.6151
R1146 B.n600 B.n597 10.6151
R1147 B.n597 B.n596 10.6151
R1148 B.n596 B.n593 10.6151
R1149 B.n593 B.n592 10.6151
R1150 B.n592 B.n589 10.6151
R1151 B.n589 B.n588 10.6151
R1152 B.n588 B.n585 10.6151
R1153 B.n585 B.n584 10.6151
R1154 B.n584 B.n581 10.6151
R1155 B.n581 B.n580 10.6151
R1156 B.n580 B.n577 10.6151
R1157 B.n577 B.n576 10.6151
R1158 B.n576 B.n573 10.6151
R1159 B.n573 B.n572 10.6151
R1160 B.n572 B.n569 10.6151
R1161 B.n569 B.n568 10.6151
R1162 B.n568 B.n565 10.6151
R1163 B.n565 B.n564 10.6151
R1164 B.n564 B.n561 10.6151
R1165 B.n561 B.n560 10.6151
R1166 B.n560 B.n557 10.6151
R1167 B.n557 B.n556 10.6151
R1168 B.n553 B.n552 10.6151
R1169 B.n552 B.n549 10.6151
R1170 B.n549 B.n548 10.6151
R1171 B.n548 B.n545 10.6151
R1172 B.n545 B.n544 10.6151
R1173 B.n544 B.n541 10.6151
R1174 B.n541 B.n540 10.6151
R1175 B.n540 B.n537 10.6151
R1176 B.n537 B.n536 10.6151
R1177 B.n533 B.n532 10.6151
R1178 B.n532 B.n529 10.6151
R1179 B.n529 B.n528 10.6151
R1180 B.n528 B.n525 10.6151
R1181 B.n525 B.n524 10.6151
R1182 B.n524 B.n521 10.6151
R1183 B.n521 B.n520 10.6151
R1184 B.n520 B.n517 10.6151
R1185 B.n517 B.n516 10.6151
R1186 B.n516 B.n513 10.6151
R1187 B.n513 B.n512 10.6151
R1188 B.n512 B.n509 10.6151
R1189 B.n509 B.n508 10.6151
R1190 B.n508 B.n505 10.6151
R1191 B.n505 B.n504 10.6151
R1192 B.n504 B.n501 10.6151
R1193 B.n501 B.n500 10.6151
R1194 B.n500 B.n497 10.6151
R1195 B.n497 B.n496 10.6151
R1196 B.n496 B.n493 10.6151
R1197 B.n493 B.n492 10.6151
R1198 B.n492 B.n489 10.6151
R1199 B.n489 B.n488 10.6151
R1200 B.n488 B.n485 10.6151
R1201 B.n485 B.n484 10.6151
R1202 B.n484 B.n481 10.6151
R1203 B.n481 B.n480 10.6151
R1204 B.n480 B.n477 10.6151
R1205 B.n477 B.n476 10.6151
R1206 B.n476 B.n473 10.6151
R1207 B.n473 B.n472 10.6151
R1208 B.n472 B.n469 10.6151
R1209 B.n469 B.n468 10.6151
R1210 B.n468 B.n465 10.6151
R1211 B.n465 B.n464 10.6151
R1212 B.n464 B.n461 10.6151
R1213 B.n461 B.n460 10.6151
R1214 B.n460 B.n457 10.6151
R1215 B.n457 B.n456 10.6151
R1216 B.n456 B.n453 10.6151
R1217 B.n453 B.n452 10.6151
R1218 B.n452 B.n449 10.6151
R1219 B.n449 B.n448 10.6151
R1220 B.n448 B.n445 10.6151
R1221 B.n445 B.n444 10.6151
R1222 B.n444 B.n441 10.6151
R1223 B.n441 B.n440 10.6151
R1224 B.n440 B.n437 10.6151
R1225 B.n437 B.n436 10.6151
R1226 B.n436 B.n433 10.6151
R1227 B.n433 B.n432 10.6151
R1228 B.n432 B.n429 10.6151
R1229 B.n429 B.n428 10.6151
R1230 B.n428 B.n426 10.6151
R1231 B.n665 B.n664 10.6151
R1232 B.n665 B.n350 10.6151
R1233 B.n676 B.n350 10.6151
R1234 B.n677 B.n676 10.6151
R1235 B.n678 B.n677 10.6151
R1236 B.n678 B.n343 10.6151
R1237 B.n688 B.n343 10.6151
R1238 B.n689 B.n688 10.6151
R1239 B.n690 B.n689 10.6151
R1240 B.n690 B.n335 10.6151
R1241 B.n702 B.n335 10.6151
R1242 B.n703 B.n702 10.6151
R1243 B.n704 B.n703 10.6151
R1244 B.n704 B.n0 10.6151
R1245 B.n761 B.n1 10.6151
R1246 B.n761 B.n760 10.6151
R1247 B.n760 B.n759 10.6151
R1248 B.n759 B.n9 10.6151
R1249 B.n753 B.n9 10.6151
R1250 B.n753 B.n752 10.6151
R1251 B.n752 B.n751 10.6151
R1252 B.n751 B.n17 10.6151
R1253 B.n745 B.n17 10.6151
R1254 B.n745 B.n744 10.6151
R1255 B.n744 B.n743 10.6151
R1256 B.n743 B.n23 10.6151
R1257 B.n737 B.n23 10.6151
R1258 B.n737 B.n736 10.6151
R1259 B.n203 B.n202 9.36635
R1260 B.n225 B.n224 9.36635
R1261 B.n556 B.n422 9.36635
R1262 B.n533 B.n425 9.36635
R1263 B.n692 B.t1 7.01804
R1264 B.t4 B.n755 7.01804
R1265 B.n700 B.t0 4.01053
R1266 B.n757 B.t19 4.01053
R1267 B.n767 B.n0 2.81026
R1268 B.n767 B.n1 2.81026
R1269 B.n204 B.n203 1.24928
R1270 B.n224 B.n223 1.24928
R1271 B.n553 B.n422 1.24928
R1272 B.n536 B.n425 1.24928
R1273 VN.n2 VN.t2 1852.23
R1274 VN.n0 VN.t1 1852.23
R1275 VN.n6 VN.t5 1852.23
R1276 VN.n4 VN.t3 1852.23
R1277 VN.n1 VN.t0 1805.49
R1278 VN.n5 VN.t4 1805.49
R1279 VN.n7 VN.n4 161.489
R1280 VN.n3 VN.n0 161.489
R1281 VN.n3 VN.n2 161.3
R1282 VN.n7 VN.n6 161.3
R1283 VN VN.n7 43.4228
R1284 VN.n1 VN.n0 36.5157
R1285 VN.n2 VN.n1 36.5157
R1286 VN.n6 VN.n5 36.5157
R1287 VN.n5 VN.n4 36.5157
R1288 VN VN.n3 0.0516364
R1289 VDD2.n183 VDD2.n182 289.615
R1290 VDD2.n90 VDD2.n89 289.615
R1291 VDD2.n182 VDD2.n181 185
R1292 VDD2.n95 VDD2.n94 185
R1293 VDD2.n176 VDD2.n175 185
R1294 VDD2.n174 VDD2.n173 185
R1295 VDD2.n99 VDD2.n98 185
R1296 VDD2.n168 VDD2.n167 185
R1297 VDD2.n166 VDD2.n165 185
R1298 VDD2.n103 VDD2.n102 185
R1299 VDD2.n160 VDD2.n159 185
R1300 VDD2.n158 VDD2.n157 185
R1301 VDD2.n107 VDD2.n106 185
R1302 VDD2.n152 VDD2.n151 185
R1303 VDD2.n150 VDD2.n149 185
R1304 VDD2.n111 VDD2.n110 185
R1305 VDD2.n115 VDD2.n113 185
R1306 VDD2.n144 VDD2.n143 185
R1307 VDD2.n142 VDD2.n141 185
R1308 VDD2.n117 VDD2.n116 185
R1309 VDD2.n136 VDD2.n135 185
R1310 VDD2.n134 VDD2.n133 185
R1311 VDD2.n121 VDD2.n120 185
R1312 VDD2.n128 VDD2.n127 185
R1313 VDD2.n126 VDD2.n125 185
R1314 VDD2.n31 VDD2.n30 185
R1315 VDD2.n33 VDD2.n32 185
R1316 VDD2.n26 VDD2.n25 185
R1317 VDD2.n39 VDD2.n38 185
R1318 VDD2.n41 VDD2.n40 185
R1319 VDD2.n22 VDD2.n21 185
R1320 VDD2.n48 VDD2.n47 185
R1321 VDD2.n49 VDD2.n20 185
R1322 VDD2.n51 VDD2.n50 185
R1323 VDD2.n18 VDD2.n17 185
R1324 VDD2.n57 VDD2.n56 185
R1325 VDD2.n59 VDD2.n58 185
R1326 VDD2.n14 VDD2.n13 185
R1327 VDD2.n65 VDD2.n64 185
R1328 VDD2.n67 VDD2.n66 185
R1329 VDD2.n10 VDD2.n9 185
R1330 VDD2.n73 VDD2.n72 185
R1331 VDD2.n75 VDD2.n74 185
R1332 VDD2.n6 VDD2.n5 185
R1333 VDD2.n81 VDD2.n80 185
R1334 VDD2.n83 VDD2.n82 185
R1335 VDD2.n2 VDD2.n1 185
R1336 VDD2.n89 VDD2.n88 185
R1337 VDD2.n124 VDD2.t5 149.524
R1338 VDD2.n29 VDD2.t3 149.524
R1339 VDD2.n182 VDD2.n94 104.615
R1340 VDD2.n175 VDD2.n94 104.615
R1341 VDD2.n175 VDD2.n174 104.615
R1342 VDD2.n174 VDD2.n98 104.615
R1343 VDD2.n167 VDD2.n98 104.615
R1344 VDD2.n167 VDD2.n166 104.615
R1345 VDD2.n166 VDD2.n102 104.615
R1346 VDD2.n159 VDD2.n102 104.615
R1347 VDD2.n159 VDD2.n158 104.615
R1348 VDD2.n158 VDD2.n106 104.615
R1349 VDD2.n151 VDD2.n106 104.615
R1350 VDD2.n151 VDD2.n150 104.615
R1351 VDD2.n150 VDD2.n110 104.615
R1352 VDD2.n115 VDD2.n110 104.615
R1353 VDD2.n143 VDD2.n115 104.615
R1354 VDD2.n143 VDD2.n142 104.615
R1355 VDD2.n142 VDD2.n116 104.615
R1356 VDD2.n135 VDD2.n116 104.615
R1357 VDD2.n135 VDD2.n134 104.615
R1358 VDD2.n134 VDD2.n120 104.615
R1359 VDD2.n127 VDD2.n120 104.615
R1360 VDD2.n127 VDD2.n126 104.615
R1361 VDD2.n32 VDD2.n31 104.615
R1362 VDD2.n32 VDD2.n25 104.615
R1363 VDD2.n39 VDD2.n25 104.615
R1364 VDD2.n40 VDD2.n39 104.615
R1365 VDD2.n40 VDD2.n21 104.615
R1366 VDD2.n48 VDD2.n21 104.615
R1367 VDD2.n49 VDD2.n48 104.615
R1368 VDD2.n50 VDD2.n49 104.615
R1369 VDD2.n50 VDD2.n17 104.615
R1370 VDD2.n57 VDD2.n17 104.615
R1371 VDD2.n58 VDD2.n57 104.615
R1372 VDD2.n58 VDD2.n13 104.615
R1373 VDD2.n65 VDD2.n13 104.615
R1374 VDD2.n66 VDD2.n65 104.615
R1375 VDD2.n66 VDD2.n9 104.615
R1376 VDD2.n73 VDD2.n9 104.615
R1377 VDD2.n74 VDD2.n73 104.615
R1378 VDD2.n74 VDD2.n5 104.615
R1379 VDD2.n81 VDD2.n5 104.615
R1380 VDD2.n82 VDD2.n81 104.615
R1381 VDD2.n82 VDD2.n1 104.615
R1382 VDD2.n89 VDD2.n1 104.615
R1383 VDD2.n92 VDD2.n91 64.5153
R1384 VDD2 VDD2.n185 64.5115
R1385 VDD2.n126 VDD2.t5 52.3082
R1386 VDD2.n31 VDD2.t3 52.3082
R1387 VDD2.n92 VDD2.n90 50.9228
R1388 VDD2.n184 VDD2.n183 50.6096
R1389 VDD2.n184 VDD2.n92 39.683
R1390 VDD2.n113 VDD2.n111 13.1884
R1391 VDD2.n51 VDD2.n18 13.1884
R1392 VDD2.n149 VDD2.n148 12.8005
R1393 VDD2.n145 VDD2.n144 12.8005
R1394 VDD2.n52 VDD2.n20 12.8005
R1395 VDD2.n56 VDD2.n55 12.8005
R1396 VDD2.n152 VDD2.n109 12.0247
R1397 VDD2.n141 VDD2.n114 12.0247
R1398 VDD2.n47 VDD2.n46 12.0247
R1399 VDD2.n59 VDD2.n16 12.0247
R1400 VDD2.n153 VDD2.n107 11.249
R1401 VDD2.n140 VDD2.n117 11.249
R1402 VDD2.n45 VDD2.n22 11.249
R1403 VDD2.n60 VDD2.n14 11.249
R1404 VDD2.n181 VDD2.n93 10.4732
R1405 VDD2.n157 VDD2.n156 10.4732
R1406 VDD2.n137 VDD2.n136 10.4732
R1407 VDD2.n42 VDD2.n41 10.4732
R1408 VDD2.n64 VDD2.n63 10.4732
R1409 VDD2.n88 VDD2.n0 10.4732
R1410 VDD2.n125 VDD2.n124 10.2747
R1411 VDD2.n30 VDD2.n29 10.2747
R1412 VDD2.n180 VDD2.n95 9.69747
R1413 VDD2.n160 VDD2.n105 9.69747
R1414 VDD2.n133 VDD2.n119 9.69747
R1415 VDD2.n38 VDD2.n24 9.69747
R1416 VDD2.n67 VDD2.n12 9.69747
R1417 VDD2.n87 VDD2.n2 9.69747
R1418 VDD2.n179 VDD2.n93 9.45567
R1419 VDD2.n86 VDD2.n0 9.45567
R1420 VDD2.n123 VDD2.n122 9.3005
R1421 VDD2.n130 VDD2.n129 9.3005
R1422 VDD2.n132 VDD2.n131 9.3005
R1423 VDD2.n119 VDD2.n118 9.3005
R1424 VDD2.n138 VDD2.n137 9.3005
R1425 VDD2.n140 VDD2.n139 9.3005
R1426 VDD2.n114 VDD2.n112 9.3005
R1427 VDD2.n146 VDD2.n145 9.3005
R1428 VDD2.n172 VDD2.n171 9.3005
R1429 VDD2.n97 VDD2.n96 9.3005
R1430 VDD2.n178 VDD2.n177 9.3005
R1431 VDD2.n180 VDD2.n179 9.3005
R1432 VDD2.n170 VDD2.n169 9.3005
R1433 VDD2.n101 VDD2.n100 9.3005
R1434 VDD2.n164 VDD2.n163 9.3005
R1435 VDD2.n162 VDD2.n161 9.3005
R1436 VDD2.n105 VDD2.n104 9.3005
R1437 VDD2.n156 VDD2.n155 9.3005
R1438 VDD2.n154 VDD2.n153 9.3005
R1439 VDD2.n109 VDD2.n108 9.3005
R1440 VDD2.n148 VDD2.n147 9.3005
R1441 VDD2.n77 VDD2.n76 9.3005
R1442 VDD2.n79 VDD2.n78 9.3005
R1443 VDD2.n4 VDD2.n3 9.3005
R1444 VDD2.n85 VDD2.n84 9.3005
R1445 VDD2.n87 VDD2.n86 9.3005
R1446 VDD2.n71 VDD2.n70 9.3005
R1447 VDD2.n69 VDD2.n68 9.3005
R1448 VDD2.n12 VDD2.n11 9.3005
R1449 VDD2.n63 VDD2.n62 9.3005
R1450 VDD2.n61 VDD2.n60 9.3005
R1451 VDD2.n16 VDD2.n15 9.3005
R1452 VDD2.n55 VDD2.n54 9.3005
R1453 VDD2.n28 VDD2.n27 9.3005
R1454 VDD2.n35 VDD2.n34 9.3005
R1455 VDD2.n37 VDD2.n36 9.3005
R1456 VDD2.n24 VDD2.n23 9.3005
R1457 VDD2.n43 VDD2.n42 9.3005
R1458 VDD2.n45 VDD2.n44 9.3005
R1459 VDD2.n46 VDD2.n19 9.3005
R1460 VDD2.n53 VDD2.n52 9.3005
R1461 VDD2.n8 VDD2.n7 9.3005
R1462 VDD2.n177 VDD2.n176 8.92171
R1463 VDD2.n161 VDD2.n103 8.92171
R1464 VDD2.n132 VDD2.n121 8.92171
R1465 VDD2.n37 VDD2.n26 8.92171
R1466 VDD2.n68 VDD2.n10 8.92171
R1467 VDD2.n84 VDD2.n83 8.92171
R1468 VDD2.n173 VDD2.n97 8.14595
R1469 VDD2.n165 VDD2.n164 8.14595
R1470 VDD2.n129 VDD2.n128 8.14595
R1471 VDD2.n34 VDD2.n33 8.14595
R1472 VDD2.n72 VDD2.n71 8.14595
R1473 VDD2.n80 VDD2.n4 8.14595
R1474 VDD2.n172 VDD2.n99 7.3702
R1475 VDD2.n168 VDD2.n101 7.3702
R1476 VDD2.n125 VDD2.n123 7.3702
R1477 VDD2.n30 VDD2.n28 7.3702
R1478 VDD2.n75 VDD2.n8 7.3702
R1479 VDD2.n79 VDD2.n6 7.3702
R1480 VDD2.n169 VDD2.n99 6.59444
R1481 VDD2.n169 VDD2.n168 6.59444
R1482 VDD2.n76 VDD2.n75 6.59444
R1483 VDD2.n76 VDD2.n6 6.59444
R1484 VDD2.n173 VDD2.n172 5.81868
R1485 VDD2.n165 VDD2.n101 5.81868
R1486 VDD2.n128 VDD2.n123 5.81868
R1487 VDD2.n33 VDD2.n28 5.81868
R1488 VDD2.n72 VDD2.n8 5.81868
R1489 VDD2.n80 VDD2.n79 5.81868
R1490 VDD2.n176 VDD2.n97 5.04292
R1491 VDD2.n164 VDD2.n103 5.04292
R1492 VDD2.n129 VDD2.n121 5.04292
R1493 VDD2.n34 VDD2.n26 5.04292
R1494 VDD2.n71 VDD2.n10 5.04292
R1495 VDD2.n83 VDD2.n4 5.04292
R1496 VDD2.n177 VDD2.n95 4.26717
R1497 VDD2.n161 VDD2.n160 4.26717
R1498 VDD2.n133 VDD2.n132 4.26717
R1499 VDD2.n38 VDD2.n37 4.26717
R1500 VDD2.n68 VDD2.n67 4.26717
R1501 VDD2.n84 VDD2.n2 4.26717
R1502 VDD2.n181 VDD2.n180 3.49141
R1503 VDD2.n157 VDD2.n105 3.49141
R1504 VDD2.n136 VDD2.n119 3.49141
R1505 VDD2.n41 VDD2.n24 3.49141
R1506 VDD2.n64 VDD2.n12 3.49141
R1507 VDD2.n88 VDD2.n87 3.49141
R1508 VDD2.n29 VDD2.n27 2.84303
R1509 VDD2.n124 VDD2.n122 2.84303
R1510 VDD2.n183 VDD2.n93 2.71565
R1511 VDD2.n156 VDD2.n107 2.71565
R1512 VDD2.n137 VDD2.n117 2.71565
R1513 VDD2.n42 VDD2.n22 2.71565
R1514 VDD2.n63 VDD2.n14 2.71565
R1515 VDD2.n90 VDD2.n0 2.71565
R1516 VDD2.n153 VDD2.n152 1.93989
R1517 VDD2.n141 VDD2.n140 1.93989
R1518 VDD2.n47 VDD2.n45 1.93989
R1519 VDD2.n60 VDD2.n59 1.93989
R1520 VDD2.n185 VDD2.t4 1.18826
R1521 VDD2.n185 VDD2.t0 1.18826
R1522 VDD2.n91 VDD2.t2 1.18826
R1523 VDD2.n91 VDD2.t1 1.18826
R1524 VDD2.n149 VDD2.n109 1.16414
R1525 VDD2.n144 VDD2.n114 1.16414
R1526 VDD2.n46 VDD2.n20 1.16414
R1527 VDD2.n56 VDD2.n16 1.16414
R1528 VDD2 VDD2.n184 0.427224
R1529 VDD2.n148 VDD2.n111 0.388379
R1530 VDD2.n145 VDD2.n113 0.388379
R1531 VDD2.n52 VDD2.n51 0.388379
R1532 VDD2.n55 VDD2.n18 0.388379
R1533 VDD2.n179 VDD2.n178 0.155672
R1534 VDD2.n178 VDD2.n96 0.155672
R1535 VDD2.n171 VDD2.n96 0.155672
R1536 VDD2.n171 VDD2.n170 0.155672
R1537 VDD2.n170 VDD2.n100 0.155672
R1538 VDD2.n163 VDD2.n100 0.155672
R1539 VDD2.n163 VDD2.n162 0.155672
R1540 VDD2.n162 VDD2.n104 0.155672
R1541 VDD2.n155 VDD2.n104 0.155672
R1542 VDD2.n155 VDD2.n154 0.155672
R1543 VDD2.n154 VDD2.n108 0.155672
R1544 VDD2.n147 VDD2.n108 0.155672
R1545 VDD2.n147 VDD2.n146 0.155672
R1546 VDD2.n146 VDD2.n112 0.155672
R1547 VDD2.n139 VDD2.n112 0.155672
R1548 VDD2.n139 VDD2.n138 0.155672
R1549 VDD2.n138 VDD2.n118 0.155672
R1550 VDD2.n131 VDD2.n118 0.155672
R1551 VDD2.n131 VDD2.n130 0.155672
R1552 VDD2.n130 VDD2.n122 0.155672
R1553 VDD2.n35 VDD2.n27 0.155672
R1554 VDD2.n36 VDD2.n35 0.155672
R1555 VDD2.n36 VDD2.n23 0.155672
R1556 VDD2.n43 VDD2.n23 0.155672
R1557 VDD2.n44 VDD2.n43 0.155672
R1558 VDD2.n44 VDD2.n19 0.155672
R1559 VDD2.n53 VDD2.n19 0.155672
R1560 VDD2.n54 VDD2.n53 0.155672
R1561 VDD2.n54 VDD2.n15 0.155672
R1562 VDD2.n61 VDD2.n15 0.155672
R1563 VDD2.n62 VDD2.n61 0.155672
R1564 VDD2.n62 VDD2.n11 0.155672
R1565 VDD2.n69 VDD2.n11 0.155672
R1566 VDD2.n70 VDD2.n69 0.155672
R1567 VDD2.n70 VDD2.n7 0.155672
R1568 VDD2.n77 VDD2.n7 0.155672
R1569 VDD2.n78 VDD2.n77 0.155672
R1570 VDD2.n78 VDD2.n3 0.155672
R1571 VDD2.n85 VDD2.n3 0.155672
R1572 VDD2.n86 VDD2.n85 0.155672
R1573 VTAIL.n374 VTAIL.n373 289.615
R1574 VTAIL.n92 VTAIL.n91 289.615
R1575 VTAIL.n282 VTAIL.n281 289.615
R1576 VTAIL.n188 VTAIL.n187 289.615
R1577 VTAIL.n315 VTAIL.n314 185
R1578 VTAIL.n317 VTAIL.n316 185
R1579 VTAIL.n310 VTAIL.n309 185
R1580 VTAIL.n323 VTAIL.n322 185
R1581 VTAIL.n325 VTAIL.n324 185
R1582 VTAIL.n306 VTAIL.n305 185
R1583 VTAIL.n332 VTAIL.n331 185
R1584 VTAIL.n333 VTAIL.n304 185
R1585 VTAIL.n335 VTAIL.n334 185
R1586 VTAIL.n302 VTAIL.n301 185
R1587 VTAIL.n341 VTAIL.n340 185
R1588 VTAIL.n343 VTAIL.n342 185
R1589 VTAIL.n298 VTAIL.n297 185
R1590 VTAIL.n349 VTAIL.n348 185
R1591 VTAIL.n351 VTAIL.n350 185
R1592 VTAIL.n294 VTAIL.n293 185
R1593 VTAIL.n357 VTAIL.n356 185
R1594 VTAIL.n359 VTAIL.n358 185
R1595 VTAIL.n290 VTAIL.n289 185
R1596 VTAIL.n365 VTAIL.n364 185
R1597 VTAIL.n367 VTAIL.n366 185
R1598 VTAIL.n286 VTAIL.n285 185
R1599 VTAIL.n373 VTAIL.n372 185
R1600 VTAIL.n33 VTAIL.n32 185
R1601 VTAIL.n35 VTAIL.n34 185
R1602 VTAIL.n28 VTAIL.n27 185
R1603 VTAIL.n41 VTAIL.n40 185
R1604 VTAIL.n43 VTAIL.n42 185
R1605 VTAIL.n24 VTAIL.n23 185
R1606 VTAIL.n50 VTAIL.n49 185
R1607 VTAIL.n51 VTAIL.n22 185
R1608 VTAIL.n53 VTAIL.n52 185
R1609 VTAIL.n20 VTAIL.n19 185
R1610 VTAIL.n59 VTAIL.n58 185
R1611 VTAIL.n61 VTAIL.n60 185
R1612 VTAIL.n16 VTAIL.n15 185
R1613 VTAIL.n67 VTAIL.n66 185
R1614 VTAIL.n69 VTAIL.n68 185
R1615 VTAIL.n12 VTAIL.n11 185
R1616 VTAIL.n75 VTAIL.n74 185
R1617 VTAIL.n77 VTAIL.n76 185
R1618 VTAIL.n8 VTAIL.n7 185
R1619 VTAIL.n83 VTAIL.n82 185
R1620 VTAIL.n85 VTAIL.n84 185
R1621 VTAIL.n4 VTAIL.n3 185
R1622 VTAIL.n91 VTAIL.n90 185
R1623 VTAIL.n281 VTAIL.n280 185
R1624 VTAIL.n194 VTAIL.n193 185
R1625 VTAIL.n275 VTAIL.n274 185
R1626 VTAIL.n273 VTAIL.n272 185
R1627 VTAIL.n198 VTAIL.n197 185
R1628 VTAIL.n267 VTAIL.n266 185
R1629 VTAIL.n265 VTAIL.n264 185
R1630 VTAIL.n202 VTAIL.n201 185
R1631 VTAIL.n259 VTAIL.n258 185
R1632 VTAIL.n257 VTAIL.n256 185
R1633 VTAIL.n206 VTAIL.n205 185
R1634 VTAIL.n251 VTAIL.n250 185
R1635 VTAIL.n249 VTAIL.n248 185
R1636 VTAIL.n210 VTAIL.n209 185
R1637 VTAIL.n214 VTAIL.n212 185
R1638 VTAIL.n243 VTAIL.n242 185
R1639 VTAIL.n241 VTAIL.n240 185
R1640 VTAIL.n216 VTAIL.n215 185
R1641 VTAIL.n235 VTAIL.n234 185
R1642 VTAIL.n233 VTAIL.n232 185
R1643 VTAIL.n220 VTAIL.n219 185
R1644 VTAIL.n227 VTAIL.n226 185
R1645 VTAIL.n225 VTAIL.n224 185
R1646 VTAIL.n187 VTAIL.n186 185
R1647 VTAIL.n100 VTAIL.n99 185
R1648 VTAIL.n181 VTAIL.n180 185
R1649 VTAIL.n179 VTAIL.n178 185
R1650 VTAIL.n104 VTAIL.n103 185
R1651 VTAIL.n173 VTAIL.n172 185
R1652 VTAIL.n171 VTAIL.n170 185
R1653 VTAIL.n108 VTAIL.n107 185
R1654 VTAIL.n165 VTAIL.n164 185
R1655 VTAIL.n163 VTAIL.n162 185
R1656 VTAIL.n112 VTAIL.n111 185
R1657 VTAIL.n157 VTAIL.n156 185
R1658 VTAIL.n155 VTAIL.n154 185
R1659 VTAIL.n116 VTAIL.n115 185
R1660 VTAIL.n120 VTAIL.n118 185
R1661 VTAIL.n149 VTAIL.n148 185
R1662 VTAIL.n147 VTAIL.n146 185
R1663 VTAIL.n122 VTAIL.n121 185
R1664 VTAIL.n141 VTAIL.n140 185
R1665 VTAIL.n139 VTAIL.n138 185
R1666 VTAIL.n126 VTAIL.n125 185
R1667 VTAIL.n133 VTAIL.n132 185
R1668 VTAIL.n131 VTAIL.n130 185
R1669 VTAIL.n313 VTAIL.t7 149.524
R1670 VTAIL.n31 VTAIL.t3 149.524
R1671 VTAIL.n223 VTAIL.t1 149.524
R1672 VTAIL.n129 VTAIL.t6 149.524
R1673 VTAIL.n316 VTAIL.n315 104.615
R1674 VTAIL.n316 VTAIL.n309 104.615
R1675 VTAIL.n323 VTAIL.n309 104.615
R1676 VTAIL.n324 VTAIL.n323 104.615
R1677 VTAIL.n324 VTAIL.n305 104.615
R1678 VTAIL.n332 VTAIL.n305 104.615
R1679 VTAIL.n333 VTAIL.n332 104.615
R1680 VTAIL.n334 VTAIL.n333 104.615
R1681 VTAIL.n334 VTAIL.n301 104.615
R1682 VTAIL.n341 VTAIL.n301 104.615
R1683 VTAIL.n342 VTAIL.n341 104.615
R1684 VTAIL.n342 VTAIL.n297 104.615
R1685 VTAIL.n349 VTAIL.n297 104.615
R1686 VTAIL.n350 VTAIL.n349 104.615
R1687 VTAIL.n350 VTAIL.n293 104.615
R1688 VTAIL.n357 VTAIL.n293 104.615
R1689 VTAIL.n358 VTAIL.n357 104.615
R1690 VTAIL.n358 VTAIL.n289 104.615
R1691 VTAIL.n365 VTAIL.n289 104.615
R1692 VTAIL.n366 VTAIL.n365 104.615
R1693 VTAIL.n366 VTAIL.n285 104.615
R1694 VTAIL.n373 VTAIL.n285 104.615
R1695 VTAIL.n34 VTAIL.n33 104.615
R1696 VTAIL.n34 VTAIL.n27 104.615
R1697 VTAIL.n41 VTAIL.n27 104.615
R1698 VTAIL.n42 VTAIL.n41 104.615
R1699 VTAIL.n42 VTAIL.n23 104.615
R1700 VTAIL.n50 VTAIL.n23 104.615
R1701 VTAIL.n51 VTAIL.n50 104.615
R1702 VTAIL.n52 VTAIL.n51 104.615
R1703 VTAIL.n52 VTAIL.n19 104.615
R1704 VTAIL.n59 VTAIL.n19 104.615
R1705 VTAIL.n60 VTAIL.n59 104.615
R1706 VTAIL.n60 VTAIL.n15 104.615
R1707 VTAIL.n67 VTAIL.n15 104.615
R1708 VTAIL.n68 VTAIL.n67 104.615
R1709 VTAIL.n68 VTAIL.n11 104.615
R1710 VTAIL.n75 VTAIL.n11 104.615
R1711 VTAIL.n76 VTAIL.n75 104.615
R1712 VTAIL.n76 VTAIL.n7 104.615
R1713 VTAIL.n83 VTAIL.n7 104.615
R1714 VTAIL.n84 VTAIL.n83 104.615
R1715 VTAIL.n84 VTAIL.n3 104.615
R1716 VTAIL.n91 VTAIL.n3 104.615
R1717 VTAIL.n281 VTAIL.n193 104.615
R1718 VTAIL.n274 VTAIL.n193 104.615
R1719 VTAIL.n274 VTAIL.n273 104.615
R1720 VTAIL.n273 VTAIL.n197 104.615
R1721 VTAIL.n266 VTAIL.n197 104.615
R1722 VTAIL.n266 VTAIL.n265 104.615
R1723 VTAIL.n265 VTAIL.n201 104.615
R1724 VTAIL.n258 VTAIL.n201 104.615
R1725 VTAIL.n258 VTAIL.n257 104.615
R1726 VTAIL.n257 VTAIL.n205 104.615
R1727 VTAIL.n250 VTAIL.n205 104.615
R1728 VTAIL.n250 VTAIL.n249 104.615
R1729 VTAIL.n249 VTAIL.n209 104.615
R1730 VTAIL.n214 VTAIL.n209 104.615
R1731 VTAIL.n242 VTAIL.n214 104.615
R1732 VTAIL.n242 VTAIL.n241 104.615
R1733 VTAIL.n241 VTAIL.n215 104.615
R1734 VTAIL.n234 VTAIL.n215 104.615
R1735 VTAIL.n234 VTAIL.n233 104.615
R1736 VTAIL.n233 VTAIL.n219 104.615
R1737 VTAIL.n226 VTAIL.n219 104.615
R1738 VTAIL.n226 VTAIL.n225 104.615
R1739 VTAIL.n187 VTAIL.n99 104.615
R1740 VTAIL.n180 VTAIL.n99 104.615
R1741 VTAIL.n180 VTAIL.n179 104.615
R1742 VTAIL.n179 VTAIL.n103 104.615
R1743 VTAIL.n172 VTAIL.n103 104.615
R1744 VTAIL.n172 VTAIL.n171 104.615
R1745 VTAIL.n171 VTAIL.n107 104.615
R1746 VTAIL.n164 VTAIL.n107 104.615
R1747 VTAIL.n164 VTAIL.n163 104.615
R1748 VTAIL.n163 VTAIL.n111 104.615
R1749 VTAIL.n156 VTAIL.n111 104.615
R1750 VTAIL.n156 VTAIL.n155 104.615
R1751 VTAIL.n155 VTAIL.n115 104.615
R1752 VTAIL.n120 VTAIL.n115 104.615
R1753 VTAIL.n148 VTAIL.n120 104.615
R1754 VTAIL.n148 VTAIL.n147 104.615
R1755 VTAIL.n147 VTAIL.n121 104.615
R1756 VTAIL.n140 VTAIL.n121 104.615
R1757 VTAIL.n140 VTAIL.n139 104.615
R1758 VTAIL.n139 VTAIL.n125 104.615
R1759 VTAIL.n132 VTAIL.n125 104.615
R1760 VTAIL.n132 VTAIL.n131 104.615
R1761 VTAIL.n315 VTAIL.t7 52.3082
R1762 VTAIL.n33 VTAIL.t3 52.3082
R1763 VTAIL.n225 VTAIL.t1 52.3082
R1764 VTAIL.n131 VTAIL.t6 52.3082
R1765 VTAIL.n191 VTAIL.n190 47.7692
R1766 VTAIL.n97 VTAIL.n96 47.7692
R1767 VTAIL.n1 VTAIL.n0 47.769
R1768 VTAIL.n95 VTAIL.n94 47.769
R1769 VTAIL.n375 VTAIL.n374 33.9308
R1770 VTAIL.n93 VTAIL.n92 33.9308
R1771 VTAIL.n283 VTAIL.n282 33.9308
R1772 VTAIL.n189 VTAIL.n188 33.9308
R1773 VTAIL.n97 VTAIL.n95 27.7203
R1774 VTAIL.n375 VTAIL.n283 27.2289
R1775 VTAIL.n335 VTAIL.n302 13.1884
R1776 VTAIL.n53 VTAIL.n20 13.1884
R1777 VTAIL.n212 VTAIL.n210 13.1884
R1778 VTAIL.n118 VTAIL.n116 13.1884
R1779 VTAIL.n336 VTAIL.n304 12.8005
R1780 VTAIL.n340 VTAIL.n339 12.8005
R1781 VTAIL.n54 VTAIL.n22 12.8005
R1782 VTAIL.n58 VTAIL.n57 12.8005
R1783 VTAIL.n248 VTAIL.n247 12.8005
R1784 VTAIL.n244 VTAIL.n243 12.8005
R1785 VTAIL.n154 VTAIL.n153 12.8005
R1786 VTAIL.n150 VTAIL.n149 12.8005
R1787 VTAIL.n331 VTAIL.n330 12.0247
R1788 VTAIL.n343 VTAIL.n300 12.0247
R1789 VTAIL.n49 VTAIL.n48 12.0247
R1790 VTAIL.n61 VTAIL.n18 12.0247
R1791 VTAIL.n251 VTAIL.n208 12.0247
R1792 VTAIL.n240 VTAIL.n213 12.0247
R1793 VTAIL.n157 VTAIL.n114 12.0247
R1794 VTAIL.n146 VTAIL.n119 12.0247
R1795 VTAIL.n329 VTAIL.n306 11.249
R1796 VTAIL.n344 VTAIL.n298 11.249
R1797 VTAIL.n47 VTAIL.n24 11.249
R1798 VTAIL.n62 VTAIL.n16 11.249
R1799 VTAIL.n252 VTAIL.n206 11.249
R1800 VTAIL.n239 VTAIL.n216 11.249
R1801 VTAIL.n158 VTAIL.n112 11.249
R1802 VTAIL.n145 VTAIL.n122 11.249
R1803 VTAIL.n326 VTAIL.n325 10.4732
R1804 VTAIL.n348 VTAIL.n347 10.4732
R1805 VTAIL.n372 VTAIL.n284 10.4732
R1806 VTAIL.n44 VTAIL.n43 10.4732
R1807 VTAIL.n66 VTAIL.n65 10.4732
R1808 VTAIL.n90 VTAIL.n2 10.4732
R1809 VTAIL.n280 VTAIL.n192 10.4732
R1810 VTAIL.n256 VTAIL.n255 10.4732
R1811 VTAIL.n236 VTAIL.n235 10.4732
R1812 VTAIL.n186 VTAIL.n98 10.4732
R1813 VTAIL.n162 VTAIL.n161 10.4732
R1814 VTAIL.n142 VTAIL.n141 10.4732
R1815 VTAIL.n314 VTAIL.n313 10.2747
R1816 VTAIL.n32 VTAIL.n31 10.2747
R1817 VTAIL.n224 VTAIL.n223 10.2747
R1818 VTAIL.n130 VTAIL.n129 10.2747
R1819 VTAIL.n322 VTAIL.n308 9.69747
R1820 VTAIL.n351 VTAIL.n296 9.69747
R1821 VTAIL.n371 VTAIL.n286 9.69747
R1822 VTAIL.n40 VTAIL.n26 9.69747
R1823 VTAIL.n69 VTAIL.n14 9.69747
R1824 VTAIL.n89 VTAIL.n4 9.69747
R1825 VTAIL.n279 VTAIL.n194 9.69747
R1826 VTAIL.n259 VTAIL.n204 9.69747
R1827 VTAIL.n232 VTAIL.n218 9.69747
R1828 VTAIL.n185 VTAIL.n100 9.69747
R1829 VTAIL.n165 VTAIL.n110 9.69747
R1830 VTAIL.n138 VTAIL.n124 9.69747
R1831 VTAIL.n370 VTAIL.n284 9.45567
R1832 VTAIL.n88 VTAIL.n2 9.45567
R1833 VTAIL.n278 VTAIL.n192 9.45567
R1834 VTAIL.n184 VTAIL.n98 9.45567
R1835 VTAIL.n361 VTAIL.n360 9.3005
R1836 VTAIL.n363 VTAIL.n362 9.3005
R1837 VTAIL.n288 VTAIL.n287 9.3005
R1838 VTAIL.n369 VTAIL.n368 9.3005
R1839 VTAIL.n371 VTAIL.n370 9.3005
R1840 VTAIL.n355 VTAIL.n354 9.3005
R1841 VTAIL.n353 VTAIL.n352 9.3005
R1842 VTAIL.n296 VTAIL.n295 9.3005
R1843 VTAIL.n347 VTAIL.n346 9.3005
R1844 VTAIL.n345 VTAIL.n344 9.3005
R1845 VTAIL.n300 VTAIL.n299 9.3005
R1846 VTAIL.n339 VTAIL.n338 9.3005
R1847 VTAIL.n312 VTAIL.n311 9.3005
R1848 VTAIL.n319 VTAIL.n318 9.3005
R1849 VTAIL.n321 VTAIL.n320 9.3005
R1850 VTAIL.n308 VTAIL.n307 9.3005
R1851 VTAIL.n327 VTAIL.n326 9.3005
R1852 VTAIL.n329 VTAIL.n328 9.3005
R1853 VTAIL.n330 VTAIL.n303 9.3005
R1854 VTAIL.n337 VTAIL.n336 9.3005
R1855 VTAIL.n292 VTAIL.n291 9.3005
R1856 VTAIL.n79 VTAIL.n78 9.3005
R1857 VTAIL.n81 VTAIL.n80 9.3005
R1858 VTAIL.n6 VTAIL.n5 9.3005
R1859 VTAIL.n87 VTAIL.n86 9.3005
R1860 VTAIL.n89 VTAIL.n88 9.3005
R1861 VTAIL.n73 VTAIL.n72 9.3005
R1862 VTAIL.n71 VTAIL.n70 9.3005
R1863 VTAIL.n14 VTAIL.n13 9.3005
R1864 VTAIL.n65 VTAIL.n64 9.3005
R1865 VTAIL.n63 VTAIL.n62 9.3005
R1866 VTAIL.n18 VTAIL.n17 9.3005
R1867 VTAIL.n57 VTAIL.n56 9.3005
R1868 VTAIL.n30 VTAIL.n29 9.3005
R1869 VTAIL.n37 VTAIL.n36 9.3005
R1870 VTAIL.n39 VTAIL.n38 9.3005
R1871 VTAIL.n26 VTAIL.n25 9.3005
R1872 VTAIL.n45 VTAIL.n44 9.3005
R1873 VTAIL.n47 VTAIL.n46 9.3005
R1874 VTAIL.n48 VTAIL.n21 9.3005
R1875 VTAIL.n55 VTAIL.n54 9.3005
R1876 VTAIL.n10 VTAIL.n9 9.3005
R1877 VTAIL.n279 VTAIL.n278 9.3005
R1878 VTAIL.n277 VTAIL.n276 9.3005
R1879 VTAIL.n196 VTAIL.n195 9.3005
R1880 VTAIL.n271 VTAIL.n270 9.3005
R1881 VTAIL.n269 VTAIL.n268 9.3005
R1882 VTAIL.n200 VTAIL.n199 9.3005
R1883 VTAIL.n263 VTAIL.n262 9.3005
R1884 VTAIL.n261 VTAIL.n260 9.3005
R1885 VTAIL.n204 VTAIL.n203 9.3005
R1886 VTAIL.n255 VTAIL.n254 9.3005
R1887 VTAIL.n253 VTAIL.n252 9.3005
R1888 VTAIL.n208 VTAIL.n207 9.3005
R1889 VTAIL.n247 VTAIL.n246 9.3005
R1890 VTAIL.n245 VTAIL.n244 9.3005
R1891 VTAIL.n213 VTAIL.n211 9.3005
R1892 VTAIL.n239 VTAIL.n238 9.3005
R1893 VTAIL.n237 VTAIL.n236 9.3005
R1894 VTAIL.n218 VTAIL.n217 9.3005
R1895 VTAIL.n231 VTAIL.n230 9.3005
R1896 VTAIL.n229 VTAIL.n228 9.3005
R1897 VTAIL.n222 VTAIL.n221 9.3005
R1898 VTAIL.n128 VTAIL.n127 9.3005
R1899 VTAIL.n135 VTAIL.n134 9.3005
R1900 VTAIL.n137 VTAIL.n136 9.3005
R1901 VTAIL.n124 VTAIL.n123 9.3005
R1902 VTAIL.n143 VTAIL.n142 9.3005
R1903 VTAIL.n145 VTAIL.n144 9.3005
R1904 VTAIL.n119 VTAIL.n117 9.3005
R1905 VTAIL.n151 VTAIL.n150 9.3005
R1906 VTAIL.n177 VTAIL.n176 9.3005
R1907 VTAIL.n102 VTAIL.n101 9.3005
R1908 VTAIL.n183 VTAIL.n182 9.3005
R1909 VTAIL.n185 VTAIL.n184 9.3005
R1910 VTAIL.n175 VTAIL.n174 9.3005
R1911 VTAIL.n106 VTAIL.n105 9.3005
R1912 VTAIL.n169 VTAIL.n168 9.3005
R1913 VTAIL.n167 VTAIL.n166 9.3005
R1914 VTAIL.n110 VTAIL.n109 9.3005
R1915 VTAIL.n161 VTAIL.n160 9.3005
R1916 VTAIL.n159 VTAIL.n158 9.3005
R1917 VTAIL.n114 VTAIL.n113 9.3005
R1918 VTAIL.n153 VTAIL.n152 9.3005
R1919 VTAIL.n321 VTAIL.n310 8.92171
R1920 VTAIL.n352 VTAIL.n294 8.92171
R1921 VTAIL.n368 VTAIL.n367 8.92171
R1922 VTAIL.n39 VTAIL.n28 8.92171
R1923 VTAIL.n70 VTAIL.n12 8.92171
R1924 VTAIL.n86 VTAIL.n85 8.92171
R1925 VTAIL.n276 VTAIL.n275 8.92171
R1926 VTAIL.n260 VTAIL.n202 8.92171
R1927 VTAIL.n231 VTAIL.n220 8.92171
R1928 VTAIL.n182 VTAIL.n181 8.92171
R1929 VTAIL.n166 VTAIL.n108 8.92171
R1930 VTAIL.n137 VTAIL.n126 8.92171
R1931 VTAIL.n318 VTAIL.n317 8.14595
R1932 VTAIL.n356 VTAIL.n355 8.14595
R1933 VTAIL.n364 VTAIL.n288 8.14595
R1934 VTAIL.n36 VTAIL.n35 8.14595
R1935 VTAIL.n74 VTAIL.n73 8.14595
R1936 VTAIL.n82 VTAIL.n6 8.14595
R1937 VTAIL.n272 VTAIL.n196 8.14595
R1938 VTAIL.n264 VTAIL.n263 8.14595
R1939 VTAIL.n228 VTAIL.n227 8.14595
R1940 VTAIL.n178 VTAIL.n102 8.14595
R1941 VTAIL.n170 VTAIL.n169 8.14595
R1942 VTAIL.n134 VTAIL.n133 8.14595
R1943 VTAIL.n314 VTAIL.n312 7.3702
R1944 VTAIL.n359 VTAIL.n292 7.3702
R1945 VTAIL.n363 VTAIL.n290 7.3702
R1946 VTAIL.n32 VTAIL.n30 7.3702
R1947 VTAIL.n77 VTAIL.n10 7.3702
R1948 VTAIL.n81 VTAIL.n8 7.3702
R1949 VTAIL.n271 VTAIL.n198 7.3702
R1950 VTAIL.n267 VTAIL.n200 7.3702
R1951 VTAIL.n224 VTAIL.n222 7.3702
R1952 VTAIL.n177 VTAIL.n104 7.3702
R1953 VTAIL.n173 VTAIL.n106 7.3702
R1954 VTAIL.n130 VTAIL.n128 7.3702
R1955 VTAIL.n360 VTAIL.n359 6.59444
R1956 VTAIL.n360 VTAIL.n290 6.59444
R1957 VTAIL.n78 VTAIL.n77 6.59444
R1958 VTAIL.n78 VTAIL.n8 6.59444
R1959 VTAIL.n268 VTAIL.n198 6.59444
R1960 VTAIL.n268 VTAIL.n267 6.59444
R1961 VTAIL.n174 VTAIL.n104 6.59444
R1962 VTAIL.n174 VTAIL.n173 6.59444
R1963 VTAIL.n317 VTAIL.n312 5.81868
R1964 VTAIL.n356 VTAIL.n292 5.81868
R1965 VTAIL.n364 VTAIL.n363 5.81868
R1966 VTAIL.n35 VTAIL.n30 5.81868
R1967 VTAIL.n74 VTAIL.n10 5.81868
R1968 VTAIL.n82 VTAIL.n81 5.81868
R1969 VTAIL.n272 VTAIL.n271 5.81868
R1970 VTAIL.n264 VTAIL.n200 5.81868
R1971 VTAIL.n227 VTAIL.n222 5.81868
R1972 VTAIL.n178 VTAIL.n177 5.81868
R1973 VTAIL.n170 VTAIL.n106 5.81868
R1974 VTAIL.n133 VTAIL.n128 5.81868
R1975 VTAIL.n318 VTAIL.n310 5.04292
R1976 VTAIL.n355 VTAIL.n294 5.04292
R1977 VTAIL.n367 VTAIL.n288 5.04292
R1978 VTAIL.n36 VTAIL.n28 5.04292
R1979 VTAIL.n73 VTAIL.n12 5.04292
R1980 VTAIL.n85 VTAIL.n6 5.04292
R1981 VTAIL.n275 VTAIL.n196 5.04292
R1982 VTAIL.n263 VTAIL.n202 5.04292
R1983 VTAIL.n228 VTAIL.n220 5.04292
R1984 VTAIL.n181 VTAIL.n102 5.04292
R1985 VTAIL.n169 VTAIL.n108 5.04292
R1986 VTAIL.n134 VTAIL.n126 5.04292
R1987 VTAIL.n322 VTAIL.n321 4.26717
R1988 VTAIL.n352 VTAIL.n351 4.26717
R1989 VTAIL.n368 VTAIL.n286 4.26717
R1990 VTAIL.n40 VTAIL.n39 4.26717
R1991 VTAIL.n70 VTAIL.n69 4.26717
R1992 VTAIL.n86 VTAIL.n4 4.26717
R1993 VTAIL.n276 VTAIL.n194 4.26717
R1994 VTAIL.n260 VTAIL.n259 4.26717
R1995 VTAIL.n232 VTAIL.n231 4.26717
R1996 VTAIL.n182 VTAIL.n100 4.26717
R1997 VTAIL.n166 VTAIL.n165 4.26717
R1998 VTAIL.n138 VTAIL.n137 4.26717
R1999 VTAIL.n325 VTAIL.n308 3.49141
R2000 VTAIL.n348 VTAIL.n296 3.49141
R2001 VTAIL.n372 VTAIL.n371 3.49141
R2002 VTAIL.n43 VTAIL.n26 3.49141
R2003 VTAIL.n66 VTAIL.n14 3.49141
R2004 VTAIL.n90 VTAIL.n89 3.49141
R2005 VTAIL.n280 VTAIL.n279 3.49141
R2006 VTAIL.n256 VTAIL.n204 3.49141
R2007 VTAIL.n235 VTAIL.n218 3.49141
R2008 VTAIL.n186 VTAIL.n185 3.49141
R2009 VTAIL.n162 VTAIL.n110 3.49141
R2010 VTAIL.n141 VTAIL.n124 3.49141
R2011 VTAIL.n313 VTAIL.n311 2.84303
R2012 VTAIL.n31 VTAIL.n29 2.84303
R2013 VTAIL.n223 VTAIL.n221 2.84303
R2014 VTAIL.n129 VTAIL.n127 2.84303
R2015 VTAIL.n326 VTAIL.n306 2.71565
R2016 VTAIL.n347 VTAIL.n298 2.71565
R2017 VTAIL.n374 VTAIL.n284 2.71565
R2018 VTAIL.n44 VTAIL.n24 2.71565
R2019 VTAIL.n65 VTAIL.n16 2.71565
R2020 VTAIL.n92 VTAIL.n2 2.71565
R2021 VTAIL.n282 VTAIL.n192 2.71565
R2022 VTAIL.n255 VTAIL.n206 2.71565
R2023 VTAIL.n236 VTAIL.n216 2.71565
R2024 VTAIL.n188 VTAIL.n98 2.71565
R2025 VTAIL.n161 VTAIL.n112 2.71565
R2026 VTAIL.n142 VTAIL.n122 2.71565
R2027 VTAIL.n331 VTAIL.n329 1.93989
R2028 VTAIL.n344 VTAIL.n343 1.93989
R2029 VTAIL.n49 VTAIL.n47 1.93989
R2030 VTAIL.n62 VTAIL.n61 1.93989
R2031 VTAIL.n252 VTAIL.n251 1.93989
R2032 VTAIL.n240 VTAIL.n239 1.93989
R2033 VTAIL.n158 VTAIL.n157 1.93989
R2034 VTAIL.n146 VTAIL.n145 1.93989
R2035 VTAIL.n0 VTAIL.t8 1.18826
R2036 VTAIL.n0 VTAIL.t9 1.18826
R2037 VTAIL.n94 VTAIL.t2 1.18826
R2038 VTAIL.n94 VTAIL.t10 1.18826
R2039 VTAIL.n190 VTAIL.t0 1.18826
R2040 VTAIL.n190 VTAIL.t11 1.18826
R2041 VTAIL.n96 VTAIL.t4 1.18826
R2042 VTAIL.n96 VTAIL.t5 1.18826
R2043 VTAIL.n330 VTAIL.n304 1.16414
R2044 VTAIL.n340 VTAIL.n300 1.16414
R2045 VTAIL.n48 VTAIL.n22 1.16414
R2046 VTAIL.n58 VTAIL.n18 1.16414
R2047 VTAIL.n248 VTAIL.n208 1.16414
R2048 VTAIL.n243 VTAIL.n213 1.16414
R2049 VTAIL.n154 VTAIL.n114 1.16414
R2050 VTAIL.n149 VTAIL.n119 1.16414
R2051 VTAIL.n191 VTAIL.n189 0.716017
R2052 VTAIL.n93 VTAIL.n1 0.716017
R2053 VTAIL.n189 VTAIL.n97 0.491879
R2054 VTAIL.n283 VTAIL.n191 0.491879
R2055 VTAIL.n95 VTAIL.n93 0.491879
R2056 VTAIL.n336 VTAIL.n335 0.388379
R2057 VTAIL.n339 VTAIL.n302 0.388379
R2058 VTAIL.n54 VTAIL.n53 0.388379
R2059 VTAIL.n57 VTAIL.n20 0.388379
R2060 VTAIL.n247 VTAIL.n210 0.388379
R2061 VTAIL.n244 VTAIL.n212 0.388379
R2062 VTAIL.n153 VTAIL.n116 0.388379
R2063 VTAIL.n150 VTAIL.n118 0.388379
R2064 VTAIL VTAIL.n375 0.310845
R2065 VTAIL VTAIL.n1 0.181534
R2066 VTAIL.n319 VTAIL.n311 0.155672
R2067 VTAIL.n320 VTAIL.n319 0.155672
R2068 VTAIL.n320 VTAIL.n307 0.155672
R2069 VTAIL.n327 VTAIL.n307 0.155672
R2070 VTAIL.n328 VTAIL.n327 0.155672
R2071 VTAIL.n328 VTAIL.n303 0.155672
R2072 VTAIL.n337 VTAIL.n303 0.155672
R2073 VTAIL.n338 VTAIL.n337 0.155672
R2074 VTAIL.n338 VTAIL.n299 0.155672
R2075 VTAIL.n345 VTAIL.n299 0.155672
R2076 VTAIL.n346 VTAIL.n345 0.155672
R2077 VTAIL.n346 VTAIL.n295 0.155672
R2078 VTAIL.n353 VTAIL.n295 0.155672
R2079 VTAIL.n354 VTAIL.n353 0.155672
R2080 VTAIL.n354 VTAIL.n291 0.155672
R2081 VTAIL.n361 VTAIL.n291 0.155672
R2082 VTAIL.n362 VTAIL.n361 0.155672
R2083 VTAIL.n362 VTAIL.n287 0.155672
R2084 VTAIL.n369 VTAIL.n287 0.155672
R2085 VTAIL.n370 VTAIL.n369 0.155672
R2086 VTAIL.n37 VTAIL.n29 0.155672
R2087 VTAIL.n38 VTAIL.n37 0.155672
R2088 VTAIL.n38 VTAIL.n25 0.155672
R2089 VTAIL.n45 VTAIL.n25 0.155672
R2090 VTAIL.n46 VTAIL.n45 0.155672
R2091 VTAIL.n46 VTAIL.n21 0.155672
R2092 VTAIL.n55 VTAIL.n21 0.155672
R2093 VTAIL.n56 VTAIL.n55 0.155672
R2094 VTAIL.n56 VTAIL.n17 0.155672
R2095 VTAIL.n63 VTAIL.n17 0.155672
R2096 VTAIL.n64 VTAIL.n63 0.155672
R2097 VTAIL.n64 VTAIL.n13 0.155672
R2098 VTAIL.n71 VTAIL.n13 0.155672
R2099 VTAIL.n72 VTAIL.n71 0.155672
R2100 VTAIL.n72 VTAIL.n9 0.155672
R2101 VTAIL.n79 VTAIL.n9 0.155672
R2102 VTAIL.n80 VTAIL.n79 0.155672
R2103 VTAIL.n80 VTAIL.n5 0.155672
R2104 VTAIL.n87 VTAIL.n5 0.155672
R2105 VTAIL.n88 VTAIL.n87 0.155672
R2106 VTAIL.n278 VTAIL.n277 0.155672
R2107 VTAIL.n277 VTAIL.n195 0.155672
R2108 VTAIL.n270 VTAIL.n195 0.155672
R2109 VTAIL.n270 VTAIL.n269 0.155672
R2110 VTAIL.n269 VTAIL.n199 0.155672
R2111 VTAIL.n262 VTAIL.n199 0.155672
R2112 VTAIL.n262 VTAIL.n261 0.155672
R2113 VTAIL.n261 VTAIL.n203 0.155672
R2114 VTAIL.n254 VTAIL.n203 0.155672
R2115 VTAIL.n254 VTAIL.n253 0.155672
R2116 VTAIL.n253 VTAIL.n207 0.155672
R2117 VTAIL.n246 VTAIL.n207 0.155672
R2118 VTAIL.n246 VTAIL.n245 0.155672
R2119 VTAIL.n245 VTAIL.n211 0.155672
R2120 VTAIL.n238 VTAIL.n211 0.155672
R2121 VTAIL.n238 VTAIL.n237 0.155672
R2122 VTAIL.n237 VTAIL.n217 0.155672
R2123 VTAIL.n230 VTAIL.n217 0.155672
R2124 VTAIL.n230 VTAIL.n229 0.155672
R2125 VTAIL.n229 VTAIL.n221 0.155672
R2126 VTAIL.n184 VTAIL.n183 0.155672
R2127 VTAIL.n183 VTAIL.n101 0.155672
R2128 VTAIL.n176 VTAIL.n101 0.155672
R2129 VTAIL.n176 VTAIL.n175 0.155672
R2130 VTAIL.n175 VTAIL.n105 0.155672
R2131 VTAIL.n168 VTAIL.n105 0.155672
R2132 VTAIL.n168 VTAIL.n167 0.155672
R2133 VTAIL.n167 VTAIL.n109 0.155672
R2134 VTAIL.n160 VTAIL.n109 0.155672
R2135 VTAIL.n160 VTAIL.n159 0.155672
R2136 VTAIL.n159 VTAIL.n113 0.155672
R2137 VTAIL.n152 VTAIL.n113 0.155672
R2138 VTAIL.n152 VTAIL.n151 0.155672
R2139 VTAIL.n151 VTAIL.n117 0.155672
R2140 VTAIL.n144 VTAIL.n117 0.155672
R2141 VTAIL.n144 VTAIL.n143 0.155672
R2142 VTAIL.n143 VTAIL.n123 0.155672
R2143 VTAIL.n136 VTAIL.n123 0.155672
R2144 VTAIL.n136 VTAIL.n135 0.155672
R2145 VTAIL.n135 VTAIL.n127 0.155672
R2146 VP.n7 VP.t4 1852.23
R2147 VP.n5 VP.t2 1852.23
R2148 VP.n0 VP.t5 1852.23
R2149 VP.n2 VP.t3 1852.23
R2150 VP.n6 VP.t0 1805.49
R2151 VP.n1 VP.t1 1805.49
R2152 VP.n3 VP.n0 161.489
R2153 VP.n8 VP.n7 161.3
R2154 VP.n3 VP.n2 161.3
R2155 VP.n5 VP.n4 161.3
R2156 VP.n4 VP.n3 43.0422
R2157 VP.n6 VP.n5 36.5157
R2158 VP.n7 VP.n6 36.5157
R2159 VP.n1 VP.n0 36.5157
R2160 VP.n2 VP.n1 36.5157
R2161 VP.n8 VP.n4 0.189894
R2162 VP VP.n8 0.0516364
R2163 VDD1.n90 VDD1.n89 289.615
R2164 VDD1.n181 VDD1.n180 289.615
R2165 VDD1.n89 VDD1.n88 185
R2166 VDD1.n2 VDD1.n1 185
R2167 VDD1.n83 VDD1.n82 185
R2168 VDD1.n81 VDD1.n80 185
R2169 VDD1.n6 VDD1.n5 185
R2170 VDD1.n75 VDD1.n74 185
R2171 VDD1.n73 VDD1.n72 185
R2172 VDD1.n10 VDD1.n9 185
R2173 VDD1.n67 VDD1.n66 185
R2174 VDD1.n65 VDD1.n64 185
R2175 VDD1.n14 VDD1.n13 185
R2176 VDD1.n59 VDD1.n58 185
R2177 VDD1.n57 VDD1.n56 185
R2178 VDD1.n18 VDD1.n17 185
R2179 VDD1.n22 VDD1.n20 185
R2180 VDD1.n51 VDD1.n50 185
R2181 VDD1.n49 VDD1.n48 185
R2182 VDD1.n24 VDD1.n23 185
R2183 VDD1.n43 VDD1.n42 185
R2184 VDD1.n41 VDD1.n40 185
R2185 VDD1.n28 VDD1.n27 185
R2186 VDD1.n35 VDD1.n34 185
R2187 VDD1.n33 VDD1.n32 185
R2188 VDD1.n122 VDD1.n121 185
R2189 VDD1.n124 VDD1.n123 185
R2190 VDD1.n117 VDD1.n116 185
R2191 VDD1.n130 VDD1.n129 185
R2192 VDD1.n132 VDD1.n131 185
R2193 VDD1.n113 VDD1.n112 185
R2194 VDD1.n139 VDD1.n138 185
R2195 VDD1.n140 VDD1.n111 185
R2196 VDD1.n142 VDD1.n141 185
R2197 VDD1.n109 VDD1.n108 185
R2198 VDD1.n148 VDD1.n147 185
R2199 VDD1.n150 VDD1.n149 185
R2200 VDD1.n105 VDD1.n104 185
R2201 VDD1.n156 VDD1.n155 185
R2202 VDD1.n158 VDD1.n157 185
R2203 VDD1.n101 VDD1.n100 185
R2204 VDD1.n164 VDD1.n163 185
R2205 VDD1.n166 VDD1.n165 185
R2206 VDD1.n97 VDD1.n96 185
R2207 VDD1.n172 VDD1.n171 185
R2208 VDD1.n174 VDD1.n173 185
R2209 VDD1.n93 VDD1.n92 185
R2210 VDD1.n180 VDD1.n179 185
R2211 VDD1.n31 VDD1.t0 149.524
R2212 VDD1.n120 VDD1.t3 149.524
R2213 VDD1.n89 VDD1.n1 104.615
R2214 VDD1.n82 VDD1.n1 104.615
R2215 VDD1.n82 VDD1.n81 104.615
R2216 VDD1.n81 VDD1.n5 104.615
R2217 VDD1.n74 VDD1.n5 104.615
R2218 VDD1.n74 VDD1.n73 104.615
R2219 VDD1.n73 VDD1.n9 104.615
R2220 VDD1.n66 VDD1.n9 104.615
R2221 VDD1.n66 VDD1.n65 104.615
R2222 VDD1.n65 VDD1.n13 104.615
R2223 VDD1.n58 VDD1.n13 104.615
R2224 VDD1.n58 VDD1.n57 104.615
R2225 VDD1.n57 VDD1.n17 104.615
R2226 VDD1.n22 VDD1.n17 104.615
R2227 VDD1.n50 VDD1.n22 104.615
R2228 VDD1.n50 VDD1.n49 104.615
R2229 VDD1.n49 VDD1.n23 104.615
R2230 VDD1.n42 VDD1.n23 104.615
R2231 VDD1.n42 VDD1.n41 104.615
R2232 VDD1.n41 VDD1.n27 104.615
R2233 VDD1.n34 VDD1.n27 104.615
R2234 VDD1.n34 VDD1.n33 104.615
R2235 VDD1.n123 VDD1.n122 104.615
R2236 VDD1.n123 VDD1.n116 104.615
R2237 VDD1.n130 VDD1.n116 104.615
R2238 VDD1.n131 VDD1.n130 104.615
R2239 VDD1.n131 VDD1.n112 104.615
R2240 VDD1.n139 VDD1.n112 104.615
R2241 VDD1.n140 VDD1.n139 104.615
R2242 VDD1.n141 VDD1.n140 104.615
R2243 VDD1.n141 VDD1.n108 104.615
R2244 VDD1.n148 VDD1.n108 104.615
R2245 VDD1.n149 VDD1.n148 104.615
R2246 VDD1.n149 VDD1.n104 104.615
R2247 VDD1.n156 VDD1.n104 104.615
R2248 VDD1.n157 VDD1.n156 104.615
R2249 VDD1.n157 VDD1.n100 104.615
R2250 VDD1.n164 VDD1.n100 104.615
R2251 VDD1.n165 VDD1.n164 104.615
R2252 VDD1.n165 VDD1.n96 104.615
R2253 VDD1.n172 VDD1.n96 104.615
R2254 VDD1.n173 VDD1.n172 104.615
R2255 VDD1.n173 VDD1.n92 104.615
R2256 VDD1.n180 VDD1.n92 104.615
R2257 VDD1.n183 VDD1.n182 64.5153
R2258 VDD1.n185 VDD1.n184 64.4468
R2259 VDD1.n33 VDD1.t0 52.3082
R2260 VDD1.n122 VDD1.t3 52.3082
R2261 VDD1 VDD1.n90 51.0363
R2262 VDD1.n183 VDD1.n181 50.9228
R2263 VDD1.n185 VDD1.n183 40.5117
R2264 VDD1.n20 VDD1.n18 13.1884
R2265 VDD1.n142 VDD1.n109 13.1884
R2266 VDD1.n56 VDD1.n55 12.8005
R2267 VDD1.n52 VDD1.n51 12.8005
R2268 VDD1.n143 VDD1.n111 12.8005
R2269 VDD1.n147 VDD1.n146 12.8005
R2270 VDD1.n59 VDD1.n16 12.0247
R2271 VDD1.n48 VDD1.n21 12.0247
R2272 VDD1.n138 VDD1.n137 12.0247
R2273 VDD1.n150 VDD1.n107 12.0247
R2274 VDD1.n60 VDD1.n14 11.249
R2275 VDD1.n47 VDD1.n24 11.249
R2276 VDD1.n136 VDD1.n113 11.249
R2277 VDD1.n151 VDD1.n105 11.249
R2278 VDD1.n88 VDD1.n0 10.4732
R2279 VDD1.n64 VDD1.n63 10.4732
R2280 VDD1.n44 VDD1.n43 10.4732
R2281 VDD1.n133 VDD1.n132 10.4732
R2282 VDD1.n155 VDD1.n154 10.4732
R2283 VDD1.n179 VDD1.n91 10.4732
R2284 VDD1.n32 VDD1.n31 10.2747
R2285 VDD1.n121 VDD1.n120 10.2747
R2286 VDD1.n87 VDD1.n2 9.69747
R2287 VDD1.n67 VDD1.n12 9.69747
R2288 VDD1.n40 VDD1.n26 9.69747
R2289 VDD1.n129 VDD1.n115 9.69747
R2290 VDD1.n158 VDD1.n103 9.69747
R2291 VDD1.n178 VDD1.n93 9.69747
R2292 VDD1.n86 VDD1.n0 9.45567
R2293 VDD1.n177 VDD1.n91 9.45567
R2294 VDD1.n30 VDD1.n29 9.3005
R2295 VDD1.n37 VDD1.n36 9.3005
R2296 VDD1.n39 VDD1.n38 9.3005
R2297 VDD1.n26 VDD1.n25 9.3005
R2298 VDD1.n45 VDD1.n44 9.3005
R2299 VDD1.n47 VDD1.n46 9.3005
R2300 VDD1.n21 VDD1.n19 9.3005
R2301 VDD1.n53 VDD1.n52 9.3005
R2302 VDD1.n79 VDD1.n78 9.3005
R2303 VDD1.n4 VDD1.n3 9.3005
R2304 VDD1.n85 VDD1.n84 9.3005
R2305 VDD1.n87 VDD1.n86 9.3005
R2306 VDD1.n77 VDD1.n76 9.3005
R2307 VDD1.n8 VDD1.n7 9.3005
R2308 VDD1.n71 VDD1.n70 9.3005
R2309 VDD1.n69 VDD1.n68 9.3005
R2310 VDD1.n12 VDD1.n11 9.3005
R2311 VDD1.n63 VDD1.n62 9.3005
R2312 VDD1.n61 VDD1.n60 9.3005
R2313 VDD1.n16 VDD1.n15 9.3005
R2314 VDD1.n55 VDD1.n54 9.3005
R2315 VDD1.n168 VDD1.n167 9.3005
R2316 VDD1.n170 VDD1.n169 9.3005
R2317 VDD1.n95 VDD1.n94 9.3005
R2318 VDD1.n176 VDD1.n175 9.3005
R2319 VDD1.n178 VDD1.n177 9.3005
R2320 VDD1.n162 VDD1.n161 9.3005
R2321 VDD1.n160 VDD1.n159 9.3005
R2322 VDD1.n103 VDD1.n102 9.3005
R2323 VDD1.n154 VDD1.n153 9.3005
R2324 VDD1.n152 VDD1.n151 9.3005
R2325 VDD1.n107 VDD1.n106 9.3005
R2326 VDD1.n146 VDD1.n145 9.3005
R2327 VDD1.n119 VDD1.n118 9.3005
R2328 VDD1.n126 VDD1.n125 9.3005
R2329 VDD1.n128 VDD1.n127 9.3005
R2330 VDD1.n115 VDD1.n114 9.3005
R2331 VDD1.n134 VDD1.n133 9.3005
R2332 VDD1.n136 VDD1.n135 9.3005
R2333 VDD1.n137 VDD1.n110 9.3005
R2334 VDD1.n144 VDD1.n143 9.3005
R2335 VDD1.n99 VDD1.n98 9.3005
R2336 VDD1.n84 VDD1.n83 8.92171
R2337 VDD1.n68 VDD1.n10 8.92171
R2338 VDD1.n39 VDD1.n28 8.92171
R2339 VDD1.n128 VDD1.n117 8.92171
R2340 VDD1.n159 VDD1.n101 8.92171
R2341 VDD1.n175 VDD1.n174 8.92171
R2342 VDD1.n80 VDD1.n4 8.14595
R2343 VDD1.n72 VDD1.n71 8.14595
R2344 VDD1.n36 VDD1.n35 8.14595
R2345 VDD1.n125 VDD1.n124 8.14595
R2346 VDD1.n163 VDD1.n162 8.14595
R2347 VDD1.n171 VDD1.n95 8.14595
R2348 VDD1.n79 VDD1.n6 7.3702
R2349 VDD1.n75 VDD1.n8 7.3702
R2350 VDD1.n32 VDD1.n30 7.3702
R2351 VDD1.n121 VDD1.n119 7.3702
R2352 VDD1.n166 VDD1.n99 7.3702
R2353 VDD1.n170 VDD1.n97 7.3702
R2354 VDD1.n76 VDD1.n6 6.59444
R2355 VDD1.n76 VDD1.n75 6.59444
R2356 VDD1.n167 VDD1.n166 6.59444
R2357 VDD1.n167 VDD1.n97 6.59444
R2358 VDD1.n80 VDD1.n79 5.81868
R2359 VDD1.n72 VDD1.n8 5.81868
R2360 VDD1.n35 VDD1.n30 5.81868
R2361 VDD1.n124 VDD1.n119 5.81868
R2362 VDD1.n163 VDD1.n99 5.81868
R2363 VDD1.n171 VDD1.n170 5.81868
R2364 VDD1.n83 VDD1.n4 5.04292
R2365 VDD1.n71 VDD1.n10 5.04292
R2366 VDD1.n36 VDD1.n28 5.04292
R2367 VDD1.n125 VDD1.n117 5.04292
R2368 VDD1.n162 VDD1.n101 5.04292
R2369 VDD1.n174 VDD1.n95 5.04292
R2370 VDD1.n84 VDD1.n2 4.26717
R2371 VDD1.n68 VDD1.n67 4.26717
R2372 VDD1.n40 VDD1.n39 4.26717
R2373 VDD1.n129 VDD1.n128 4.26717
R2374 VDD1.n159 VDD1.n158 4.26717
R2375 VDD1.n175 VDD1.n93 4.26717
R2376 VDD1.n88 VDD1.n87 3.49141
R2377 VDD1.n64 VDD1.n12 3.49141
R2378 VDD1.n43 VDD1.n26 3.49141
R2379 VDD1.n132 VDD1.n115 3.49141
R2380 VDD1.n155 VDD1.n103 3.49141
R2381 VDD1.n179 VDD1.n178 3.49141
R2382 VDD1.n120 VDD1.n118 2.84303
R2383 VDD1.n31 VDD1.n29 2.84303
R2384 VDD1.n90 VDD1.n0 2.71565
R2385 VDD1.n63 VDD1.n14 2.71565
R2386 VDD1.n44 VDD1.n24 2.71565
R2387 VDD1.n133 VDD1.n113 2.71565
R2388 VDD1.n154 VDD1.n105 2.71565
R2389 VDD1.n181 VDD1.n91 2.71565
R2390 VDD1.n60 VDD1.n59 1.93989
R2391 VDD1.n48 VDD1.n47 1.93989
R2392 VDD1.n138 VDD1.n136 1.93989
R2393 VDD1.n151 VDD1.n150 1.93989
R2394 VDD1.n184 VDD1.t4 1.18826
R2395 VDD1.n184 VDD1.t2 1.18826
R2396 VDD1.n182 VDD1.t5 1.18826
R2397 VDD1.n182 VDD1.t1 1.18826
R2398 VDD1.n56 VDD1.n16 1.16414
R2399 VDD1.n51 VDD1.n21 1.16414
R2400 VDD1.n137 VDD1.n111 1.16414
R2401 VDD1.n147 VDD1.n107 1.16414
R2402 VDD1.n55 VDD1.n18 0.388379
R2403 VDD1.n52 VDD1.n20 0.388379
R2404 VDD1.n143 VDD1.n142 0.388379
R2405 VDD1.n146 VDD1.n109 0.388379
R2406 VDD1.n86 VDD1.n85 0.155672
R2407 VDD1.n85 VDD1.n3 0.155672
R2408 VDD1.n78 VDD1.n3 0.155672
R2409 VDD1.n78 VDD1.n77 0.155672
R2410 VDD1.n77 VDD1.n7 0.155672
R2411 VDD1.n70 VDD1.n7 0.155672
R2412 VDD1.n70 VDD1.n69 0.155672
R2413 VDD1.n69 VDD1.n11 0.155672
R2414 VDD1.n62 VDD1.n11 0.155672
R2415 VDD1.n62 VDD1.n61 0.155672
R2416 VDD1.n61 VDD1.n15 0.155672
R2417 VDD1.n54 VDD1.n15 0.155672
R2418 VDD1.n54 VDD1.n53 0.155672
R2419 VDD1.n53 VDD1.n19 0.155672
R2420 VDD1.n46 VDD1.n19 0.155672
R2421 VDD1.n46 VDD1.n45 0.155672
R2422 VDD1.n45 VDD1.n25 0.155672
R2423 VDD1.n38 VDD1.n25 0.155672
R2424 VDD1.n38 VDD1.n37 0.155672
R2425 VDD1.n37 VDD1.n29 0.155672
R2426 VDD1.n126 VDD1.n118 0.155672
R2427 VDD1.n127 VDD1.n126 0.155672
R2428 VDD1.n127 VDD1.n114 0.155672
R2429 VDD1.n134 VDD1.n114 0.155672
R2430 VDD1.n135 VDD1.n134 0.155672
R2431 VDD1.n135 VDD1.n110 0.155672
R2432 VDD1.n144 VDD1.n110 0.155672
R2433 VDD1.n145 VDD1.n144 0.155672
R2434 VDD1.n145 VDD1.n106 0.155672
R2435 VDD1.n152 VDD1.n106 0.155672
R2436 VDD1.n153 VDD1.n152 0.155672
R2437 VDD1.n153 VDD1.n102 0.155672
R2438 VDD1.n160 VDD1.n102 0.155672
R2439 VDD1.n161 VDD1.n160 0.155672
R2440 VDD1.n161 VDD1.n98 0.155672
R2441 VDD1.n168 VDD1.n98 0.155672
R2442 VDD1.n169 VDD1.n168 0.155672
R2443 VDD1.n169 VDD1.n94 0.155672
R2444 VDD1.n176 VDD1.n94 0.155672
R2445 VDD1.n177 VDD1.n176 0.155672
R2446 VDD1 VDD1.n185 0.0651552
C0 VP VTAIL 2.50966f
C1 VTAIL VDD2 20.5207f
C2 VN VTAIL 2.49461f
C3 VTAIL VDD1 20.4954f
C4 VP VDD2 0.259576f
C5 VP VN 5.49758f
C6 VP VDD1 3.30524f
C7 VN VDD2 3.20019f
C8 VDD1 VDD2 0.550866f
C9 VN VDD1 0.147327f
C10 VDD2 B 4.991261f
C11 VDD1 B 4.940145f
C12 VTAIL B 7.607903f
C13 VN B 7.40075f
C14 VP B 4.69405f
C15 VDD1.n0 B 0.016771f
C16 VDD1.n1 B 0.037735f
C17 VDD1.n2 B 0.016904f
C18 VDD1.n3 B 0.02971f
C19 VDD1.n4 B 0.015965f
C20 VDD1.n5 B 0.037735f
C21 VDD1.n6 B 0.016904f
C22 VDD1.n7 B 0.02971f
C23 VDD1.n8 B 0.015965f
C24 VDD1.n9 B 0.037735f
C25 VDD1.n10 B 0.016904f
C26 VDD1.n11 B 0.02971f
C27 VDD1.n12 B 0.015965f
C28 VDD1.n13 B 0.037735f
C29 VDD1.n14 B 0.016904f
C30 VDD1.n15 B 0.02971f
C31 VDD1.n16 B 0.015965f
C32 VDD1.n17 B 0.037735f
C33 VDD1.n18 B 0.016434f
C34 VDD1.n19 B 0.02971f
C35 VDD1.n20 B 0.016434f
C36 VDD1.n21 B 0.015965f
C37 VDD1.n22 B 0.037735f
C38 VDD1.n23 B 0.037735f
C39 VDD1.n24 B 0.016904f
C40 VDD1.n25 B 0.02971f
C41 VDD1.n26 B 0.015965f
C42 VDD1.n27 B 0.037735f
C43 VDD1.n28 B 0.016904f
C44 VDD1.n29 B 2.11594f
C45 VDD1.n30 B 0.015965f
C46 VDD1.t0 B 0.064479f
C47 VDD1.n31 B 0.267472f
C48 VDD1.n32 B 0.026676f
C49 VDD1.n33 B 0.028301f
C50 VDD1.n34 B 0.037735f
C51 VDD1.n35 B 0.016904f
C52 VDD1.n36 B 0.015965f
C53 VDD1.n37 B 0.02971f
C54 VDD1.n38 B 0.02971f
C55 VDD1.n39 B 0.015965f
C56 VDD1.n40 B 0.016904f
C57 VDD1.n41 B 0.037735f
C58 VDD1.n42 B 0.037735f
C59 VDD1.n43 B 0.016904f
C60 VDD1.n44 B 0.015965f
C61 VDD1.n45 B 0.02971f
C62 VDD1.n46 B 0.02971f
C63 VDD1.n47 B 0.015965f
C64 VDD1.n48 B 0.016904f
C65 VDD1.n49 B 0.037735f
C66 VDD1.n50 B 0.037735f
C67 VDD1.n51 B 0.016904f
C68 VDD1.n52 B 0.015965f
C69 VDD1.n53 B 0.02971f
C70 VDD1.n54 B 0.02971f
C71 VDD1.n55 B 0.015965f
C72 VDD1.n56 B 0.016904f
C73 VDD1.n57 B 0.037735f
C74 VDD1.n58 B 0.037735f
C75 VDD1.n59 B 0.016904f
C76 VDD1.n60 B 0.015965f
C77 VDD1.n61 B 0.02971f
C78 VDD1.n62 B 0.02971f
C79 VDD1.n63 B 0.015965f
C80 VDD1.n64 B 0.016904f
C81 VDD1.n65 B 0.037735f
C82 VDD1.n66 B 0.037735f
C83 VDD1.n67 B 0.016904f
C84 VDD1.n68 B 0.015965f
C85 VDD1.n69 B 0.02971f
C86 VDD1.n70 B 0.02971f
C87 VDD1.n71 B 0.015965f
C88 VDD1.n72 B 0.016904f
C89 VDD1.n73 B 0.037735f
C90 VDD1.n74 B 0.037735f
C91 VDD1.n75 B 0.016904f
C92 VDD1.n76 B 0.015965f
C93 VDD1.n77 B 0.02971f
C94 VDD1.n78 B 0.02971f
C95 VDD1.n79 B 0.015965f
C96 VDD1.n80 B 0.016904f
C97 VDD1.n81 B 0.037735f
C98 VDD1.n82 B 0.037735f
C99 VDD1.n83 B 0.016904f
C100 VDD1.n84 B 0.015965f
C101 VDD1.n85 B 0.02971f
C102 VDD1.n86 B 0.078008f
C103 VDD1.n87 B 0.015965f
C104 VDD1.n88 B 0.016904f
C105 VDD1.n89 B 0.074246f
C106 VDD1.n90 B 0.085435f
C107 VDD1.n91 B 0.016771f
C108 VDD1.n92 B 0.037735f
C109 VDD1.n93 B 0.016904f
C110 VDD1.n94 B 0.02971f
C111 VDD1.n95 B 0.015965f
C112 VDD1.n96 B 0.037735f
C113 VDD1.n97 B 0.016904f
C114 VDD1.n98 B 0.02971f
C115 VDD1.n99 B 0.015965f
C116 VDD1.n100 B 0.037735f
C117 VDD1.n101 B 0.016904f
C118 VDD1.n102 B 0.02971f
C119 VDD1.n103 B 0.015965f
C120 VDD1.n104 B 0.037735f
C121 VDD1.n105 B 0.016904f
C122 VDD1.n106 B 0.02971f
C123 VDD1.n107 B 0.015965f
C124 VDD1.n108 B 0.037735f
C125 VDD1.n109 B 0.016434f
C126 VDD1.n110 B 0.02971f
C127 VDD1.n111 B 0.016904f
C128 VDD1.n112 B 0.037735f
C129 VDD1.n113 B 0.016904f
C130 VDD1.n114 B 0.02971f
C131 VDD1.n115 B 0.015965f
C132 VDD1.n116 B 0.037735f
C133 VDD1.n117 B 0.016904f
C134 VDD1.n118 B 2.11594f
C135 VDD1.n119 B 0.015965f
C136 VDD1.t3 B 0.064479f
C137 VDD1.n120 B 0.267472f
C138 VDD1.n121 B 0.026676f
C139 VDD1.n122 B 0.028301f
C140 VDD1.n123 B 0.037735f
C141 VDD1.n124 B 0.016904f
C142 VDD1.n125 B 0.015965f
C143 VDD1.n126 B 0.02971f
C144 VDD1.n127 B 0.02971f
C145 VDD1.n128 B 0.015965f
C146 VDD1.n129 B 0.016904f
C147 VDD1.n130 B 0.037735f
C148 VDD1.n131 B 0.037735f
C149 VDD1.n132 B 0.016904f
C150 VDD1.n133 B 0.015965f
C151 VDD1.n134 B 0.02971f
C152 VDD1.n135 B 0.02971f
C153 VDD1.n136 B 0.015965f
C154 VDD1.n137 B 0.015965f
C155 VDD1.n138 B 0.016904f
C156 VDD1.n139 B 0.037735f
C157 VDD1.n140 B 0.037735f
C158 VDD1.n141 B 0.037735f
C159 VDD1.n142 B 0.016434f
C160 VDD1.n143 B 0.015965f
C161 VDD1.n144 B 0.02971f
C162 VDD1.n145 B 0.02971f
C163 VDD1.n146 B 0.015965f
C164 VDD1.n147 B 0.016904f
C165 VDD1.n148 B 0.037735f
C166 VDD1.n149 B 0.037735f
C167 VDD1.n150 B 0.016904f
C168 VDD1.n151 B 0.015965f
C169 VDD1.n152 B 0.02971f
C170 VDD1.n153 B 0.02971f
C171 VDD1.n154 B 0.015965f
C172 VDD1.n155 B 0.016904f
C173 VDD1.n156 B 0.037735f
C174 VDD1.n157 B 0.037735f
C175 VDD1.n158 B 0.016904f
C176 VDD1.n159 B 0.015965f
C177 VDD1.n160 B 0.02971f
C178 VDD1.n161 B 0.02971f
C179 VDD1.n162 B 0.015965f
C180 VDD1.n163 B 0.016904f
C181 VDD1.n164 B 0.037735f
C182 VDD1.n165 B 0.037735f
C183 VDD1.n166 B 0.016904f
C184 VDD1.n167 B 0.015965f
C185 VDD1.n168 B 0.02971f
C186 VDD1.n169 B 0.02971f
C187 VDD1.n170 B 0.015965f
C188 VDD1.n171 B 0.016904f
C189 VDD1.n172 B 0.037735f
C190 VDD1.n173 B 0.037735f
C191 VDD1.n174 B 0.016904f
C192 VDD1.n175 B 0.015965f
C193 VDD1.n176 B 0.02971f
C194 VDD1.n177 B 0.078008f
C195 VDD1.n178 B 0.015965f
C196 VDD1.n179 B 0.016904f
C197 VDD1.n180 B 0.074246f
C198 VDD1.n181 B 0.08516f
C199 VDD1.t5 B 0.391374f
C200 VDD1.t1 B 0.391374f
C201 VDD1.n182 B 3.56794f
C202 VDD1.n183 B 2.37234f
C203 VDD1.t4 B 0.391374f
C204 VDD1.t2 B 0.391374f
C205 VDD1.n184 B 3.56762f
C206 VDD1.n185 B 2.9396f
C207 VP.t5 B 0.69718f
C208 VP.n0 B 0.284099f
C209 VP.t1 B 0.690421f
C210 VP.n1 B 0.265562f
C211 VP.t3 B 0.69718f
C212 VP.n2 B 0.284011f
C213 VP.n3 B 2.70599f
C214 VP.n4 B 2.68165f
C215 VP.t0 B 0.690421f
C216 VP.t2 B 0.69718f
C217 VP.n5 B 0.284011f
C218 VP.n6 B 0.265562f
C219 VP.t4 B 0.69718f
C220 VP.n7 B 0.284011f
C221 VP.n8 B 0.047427f
C222 VTAIL.t8 B 0.395467f
C223 VTAIL.t9 B 0.395467f
C224 VTAIL.n0 B 3.52509f
C225 VTAIL.n1 B 0.360151f
C226 VTAIL.n2 B 0.016946f
C227 VTAIL.n3 B 0.03813f
C228 VTAIL.n4 B 0.017081f
C229 VTAIL.n5 B 0.030021f
C230 VTAIL.n6 B 0.016132f
C231 VTAIL.n7 B 0.03813f
C232 VTAIL.n8 B 0.017081f
C233 VTAIL.n9 B 0.030021f
C234 VTAIL.n10 B 0.016132f
C235 VTAIL.n11 B 0.03813f
C236 VTAIL.n12 B 0.017081f
C237 VTAIL.n13 B 0.030021f
C238 VTAIL.n14 B 0.016132f
C239 VTAIL.n15 B 0.03813f
C240 VTAIL.n16 B 0.017081f
C241 VTAIL.n17 B 0.030021f
C242 VTAIL.n18 B 0.016132f
C243 VTAIL.n19 B 0.03813f
C244 VTAIL.n20 B 0.016606f
C245 VTAIL.n21 B 0.030021f
C246 VTAIL.n22 B 0.017081f
C247 VTAIL.n23 B 0.03813f
C248 VTAIL.n24 B 0.017081f
C249 VTAIL.n25 B 0.030021f
C250 VTAIL.n26 B 0.016132f
C251 VTAIL.n27 B 0.03813f
C252 VTAIL.n28 B 0.017081f
C253 VTAIL.n29 B 2.13807f
C254 VTAIL.n30 B 0.016132f
C255 VTAIL.t3 B 0.065154f
C256 VTAIL.n31 B 0.27027f
C257 VTAIL.n32 B 0.026955f
C258 VTAIL.n33 B 0.028597f
C259 VTAIL.n34 B 0.03813f
C260 VTAIL.n35 B 0.017081f
C261 VTAIL.n36 B 0.016132f
C262 VTAIL.n37 B 0.030021f
C263 VTAIL.n38 B 0.030021f
C264 VTAIL.n39 B 0.016132f
C265 VTAIL.n40 B 0.017081f
C266 VTAIL.n41 B 0.03813f
C267 VTAIL.n42 B 0.03813f
C268 VTAIL.n43 B 0.017081f
C269 VTAIL.n44 B 0.016132f
C270 VTAIL.n45 B 0.030021f
C271 VTAIL.n46 B 0.030021f
C272 VTAIL.n47 B 0.016132f
C273 VTAIL.n48 B 0.016132f
C274 VTAIL.n49 B 0.017081f
C275 VTAIL.n50 B 0.03813f
C276 VTAIL.n51 B 0.03813f
C277 VTAIL.n52 B 0.03813f
C278 VTAIL.n53 B 0.016606f
C279 VTAIL.n54 B 0.016132f
C280 VTAIL.n55 B 0.030021f
C281 VTAIL.n56 B 0.030021f
C282 VTAIL.n57 B 0.016132f
C283 VTAIL.n58 B 0.017081f
C284 VTAIL.n59 B 0.03813f
C285 VTAIL.n60 B 0.03813f
C286 VTAIL.n61 B 0.017081f
C287 VTAIL.n62 B 0.016132f
C288 VTAIL.n63 B 0.030021f
C289 VTAIL.n64 B 0.030021f
C290 VTAIL.n65 B 0.016132f
C291 VTAIL.n66 B 0.017081f
C292 VTAIL.n67 B 0.03813f
C293 VTAIL.n68 B 0.03813f
C294 VTAIL.n69 B 0.017081f
C295 VTAIL.n70 B 0.016132f
C296 VTAIL.n71 B 0.030021f
C297 VTAIL.n72 B 0.030021f
C298 VTAIL.n73 B 0.016132f
C299 VTAIL.n74 B 0.017081f
C300 VTAIL.n75 B 0.03813f
C301 VTAIL.n76 B 0.03813f
C302 VTAIL.n77 B 0.017081f
C303 VTAIL.n78 B 0.016132f
C304 VTAIL.n79 B 0.030021f
C305 VTAIL.n80 B 0.030021f
C306 VTAIL.n81 B 0.016132f
C307 VTAIL.n82 B 0.017081f
C308 VTAIL.n83 B 0.03813f
C309 VTAIL.n84 B 0.03813f
C310 VTAIL.n85 B 0.017081f
C311 VTAIL.n86 B 0.016132f
C312 VTAIL.n87 B 0.030021f
C313 VTAIL.n88 B 0.078824f
C314 VTAIL.n89 B 0.016132f
C315 VTAIL.n90 B 0.017081f
C316 VTAIL.n91 B 0.075023f
C317 VTAIL.n92 B 0.064781f
C318 VTAIL.n93 B 0.144473f
C319 VTAIL.t2 B 0.395467f
C320 VTAIL.t10 B 0.395467f
C321 VTAIL.n94 B 3.52509f
C322 VTAIL.n95 B 2.21394f
C323 VTAIL.t4 B 0.395467f
C324 VTAIL.t5 B 0.395467f
C325 VTAIL.n96 B 3.52509f
C326 VTAIL.n97 B 2.21394f
C327 VTAIL.n98 B 0.016946f
C328 VTAIL.n99 B 0.03813f
C329 VTAIL.n100 B 0.017081f
C330 VTAIL.n101 B 0.030021f
C331 VTAIL.n102 B 0.016132f
C332 VTAIL.n103 B 0.03813f
C333 VTAIL.n104 B 0.017081f
C334 VTAIL.n105 B 0.030021f
C335 VTAIL.n106 B 0.016132f
C336 VTAIL.n107 B 0.03813f
C337 VTAIL.n108 B 0.017081f
C338 VTAIL.n109 B 0.030021f
C339 VTAIL.n110 B 0.016132f
C340 VTAIL.n111 B 0.03813f
C341 VTAIL.n112 B 0.017081f
C342 VTAIL.n113 B 0.030021f
C343 VTAIL.n114 B 0.016132f
C344 VTAIL.n115 B 0.03813f
C345 VTAIL.n116 B 0.016606f
C346 VTAIL.n117 B 0.030021f
C347 VTAIL.n118 B 0.016606f
C348 VTAIL.n119 B 0.016132f
C349 VTAIL.n120 B 0.03813f
C350 VTAIL.n121 B 0.03813f
C351 VTAIL.n122 B 0.017081f
C352 VTAIL.n123 B 0.030021f
C353 VTAIL.n124 B 0.016132f
C354 VTAIL.n125 B 0.03813f
C355 VTAIL.n126 B 0.017081f
C356 VTAIL.n127 B 2.13807f
C357 VTAIL.n128 B 0.016132f
C358 VTAIL.t6 B 0.065154f
C359 VTAIL.n129 B 0.27027f
C360 VTAIL.n130 B 0.026955f
C361 VTAIL.n131 B 0.028597f
C362 VTAIL.n132 B 0.03813f
C363 VTAIL.n133 B 0.017081f
C364 VTAIL.n134 B 0.016132f
C365 VTAIL.n135 B 0.030021f
C366 VTAIL.n136 B 0.030021f
C367 VTAIL.n137 B 0.016132f
C368 VTAIL.n138 B 0.017081f
C369 VTAIL.n139 B 0.03813f
C370 VTAIL.n140 B 0.03813f
C371 VTAIL.n141 B 0.017081f
C372 VTAIL.n142 B 0.016132f
C373 VTAIL.n143 B 0.030021f
C374 VTAIL.n144 B 0.030021f
C375 VTAIL.n145 B 0.016132f
C376 VTAIL.n146 B 0.017081f
C377 VTAIL.n147 B 0.03813f
C378 VTAIL.n148 B 0.03813f
C379 VTAIL.n149 B 0.017081f
C380 VTAIL.n150 B 0.016132f
C381 VTAIL.n151 B 0.030021f
C382 VTAIL.n152 B 0.030021f
C383 VTAIL.n153 B 0.016132f
C384 VTAIL.n154 B 0.017081f
C385 VTAIL.n155 B 0.03813f
C386 VTAIL.n156 B 0.03813f
C387 VTAIL.n157 B 0.017081f
C388 VTAIL.n158 B 0.016132f
C389 VTAIL.n159 B 0.030021f
C390 VTAIL.n160 B 0.030021f
C391 VTAIL.n161 B 0.016132f
C392 VTAIL.n162 B 0.017081f
C393 VTAIL.n163 B 0.03813f
C394 VTAIL.n164 B 0.03813f
C395 VTAIL.n165 B 0.017081f
C396 VTAIL.n166 B 0.016132f
C397 VTAIL.n167 B 0.030021f
C398 VTAIL.n168 B 0.030021f
C399 VTAIL.n169 B 0.016132f
C400 VTAIL.n170 B 0.017081f
C401 VTAIL.n171 B 0.03813f
C402 VTAIL.n172 B 0.03813f
C403 VTAIL.n173 B 0.017081f
C404 VTAIL.n174 B 0.016132f
C405 VTAIL.n175 B 0.030021f
C406 VTAIL.n176 B 0.030021f
C407 VTAIL.n177 B 0.016132f
C408 VTAIL.n178 B 0.017081f
C409 VTAIL.n179 B 0.03813f
C410 VTAIL.n180 B 0.03813f
C411 VTAIL.n181 B 0.017081f
C412 VTAIL.n182 B 0.016132f
C413 VTAIL.n183 B 0.030021f
C414 VTAIL.n184 B 0.078824f
C415 VTAIL.n185 B 0.016132f
C416 VTAIL.n186 B 0.017081f
C417 VTAIL.n187 B 0.075023f
C418 VTAIL.n188 B 0.064781f
C419 VTAIL.n189 B 0.144473f
C420 VTAIL.t0 B 0.395467f
C421 VTAIL.t11 B 0.395467f
C422 VTAIL.n190 B 3.52509f
C423 VTAIL.n191 B 0.390164f
C424 VTAIL.n192 B 0.016946f
C425 VTAIL.n193 B 0.03813f
C426 VTAIL.n194 B 0.017081f
C427 VTAIL.n195 B 0.030021f
C428 VTAIL.n196 B 0.016132f
C429 VTAIL.n197 B 0.03813f
C430 VTAIL.n198 B 0.017081f
C431 VTAIL.n199 B 0.030021f
C432 VTAIL.n200 B 0.016132f
C433 VTAIL.n201 B 0.03813f
C434 VTAIL.n202 B 0.017081f
C435 VTAIL.n203 B 0.030021f
C436 VTAIL.n204 B 0.016132f
C437 VTAIL.n205 B 0.03813f
C438 VTAIL.n206 B 0.017081f
C439 VTAIL.n207 B 0.030021f
C440 VTAIL.n208 B 0.016132f
C441 VTAIL.n209 B 0.03813f
C442 VTAIL.n210 B 0.016606f
C443 VTAIL.n211 B 0.030021f
C444 VTAIL.n212 B 0.016606f
C445 VTAIL.n213 B 0.016132f
C446 VTAIL.n214 B 0.03813f
C447 VTAIL.n215 B 0.03813f
C448 VTAIL.n216 B 0.017081f
C449 VTAIL.n217 B 0.030021f
C450 VTAIL.n218 B 0.016132f
C451 VTAIL.n219 B 0.03813f
C452 VTAIL.n220 B 0.017081f
C453 VTAIL.n221 B 2.13807f
C454 VTAIL.n222 B 0.016132f
C455 VTAIL.t1 B 0.065154f
C456 VTAIL.n223 B 0.27027f
C457 VTAIL.n224 B 0.026955f
C458 VTAIL.n225 B 0.028597f
C459 VTAIL.n226 B 0.03813f
C460 VTAIL.n227 B 0.017081f
C461 VTAIL.n228 B 0.016132f
C462 VTAIL.n229 B 0.030021f
C463 VTAIL.n230 B 0.030021f
C464 VTAIL.n231 B 0.016132f
C465 VTAIL.n232 B 0.017081f
C466 VTAIL.n233 B 0.03813f
C467 VTAIL.n234 B 0.03813f
C468 VTAIL.n235 B 0.017081f
C469 VTAIL.n236 B 0.016132f
C470 VTAIL.n237 B 0.030021f
C471 VTAIL.n238 B 0.030021f
C472 VTAIL.n239 B 0.016132f
C473 VTAIL.n240 B 0.017081f
C474 VTAIL.n241 B 0.03813f
C475 VTAIL.n242 B 0.03813f
C476 VTAIL.n243 B 0.017081f
C477 VTAIL.n244 B 0.016132f
C478 VTAIL.n245 B 0.030021f
C479 VTAIL.n246 B 0.030021f
C480 VTAIL.n247 B 0.016132f
C481 VTAIL.n248 B 0.017081f
C482 VTAIL.n249 B 0.03813f
C483 VTAIL.n250 B 0.03813f
C484 VTAIL.n251 B 0.017081f
C485 VTAIL.n252 B 0.016132f
C486 VTAIL.n253 B 0.030021f
C487 VTAIL.n254 B 0.030021f
C488 VTAIL.n255 B 0.016132f
C489 VTAIL.n256 B 0.017081f
C490 VTAIL.n257 B 0.03813f
C491 VTAIL.n258 B 0.03813f
C492 VTAIL.n259 B 0.017081f
C493 VTAIL.n260 B 0.016132f
C494 VTAIL.n261 B 0.030021f
C495 VTAIL.n262 B 0.030021f
C496 VTAIL.n263 B 0.016132f
C497 VTAIL.n264 B 0.017081f
C498 VTAIL.n265 B 0.03813f
C499 VTAIL.n266 B 0.03813f
C500 VTAIL.n267 B 0.017081f
C501 VTAIL.n268 B 0.016132f
C502 VTAIL.n269 B 0.030021f
C503 VTAIL.n270 B 0.030021f
C504 VTAIL.n271 B 0.016132f
C505 VTAIL.n272 B 0.017081f
C506 VTAIL.n273 B 0.03813f
C507 VTAIL.n274 B 0.03813f
C508 VTAIL.n275 B 0.017081f
C509 VTAIL.n276 B 0.016132f
C510 VTAIL.n277 B 0.030021f
C511 VTAIL.n278 B 0.078824f
C512 VTAIL.n279 B 0.016132f
C513 VTAIL.n280 B 0.017081f
C514 VTAIL.n281 B 0.075023f
C515 VTAIL.n282 B 0.064781f
C516 VTAIL.n283 B 1.92071f
C517 VTAIL.n284 B 0.016946f
C518 VTAIL.n285 B 0.03813f
C519 VTAIL.n286 B 0.017081f
C520 VTAIL.n287 B 0.030021f
C521 VTAIL.n288 B 0.016132f
C522 VTAIL.n289 B 0.03813f
C523 VTAIL.n290 B 0.017081f
C524 VTAIL.n291 B 0.030021f
C525 VTAIL.n292 B 0.016132f
C526 VTAIL.n293 B 0.03813f
C527 VTAIL.n294 B 0.017081f
C528 VTAIL.n295 B 0.030021f
C529 VTAIL.n296 B 0.016132f
C530 VTAIL.n297 B 0.03813f
C531 VTAIL.n298 B 0.017081f
C532 VTAIL.n299 B 0.030021f
C533 VTAIL.n300 B 0.016132f
C534 VTAIL.n301 B 0.03813f
C535 VTAIL.n302 B 0.016606f
C536 VTAIL.n303 B 0.030021f
C537 VTAIL.n304 B 0.017081f
C538 VTAIL.n305 B 0.03813f
C539 VTAIL.n306 B 0.017081f
C540 VTAIL.n307 B 0.030021f
C541 VTAIL.n308 B 0.016132f
C542 VTAIL.n309 B 0.03813f
C543 VTAIL.n310 B 0.017081f
C544 VTAIL.n311 B 2.13807f
C545 VTAIL.n312 B 0.016132f
C546 VTAIL.t7 B 0.065154f
C547 VTAIL.n313 B 0.27027f
C548 VTAIL.n314 B 0.026955f
C549 VTAIL.n315 B 0.028597f
C550 VTAIL.n316 B 0.03813f
C551 VTAIL.n317 B 0.017081f
C552 VTAIL.n318 B 0.016132f
C553 VTAIL.n319 B 0.030021f
C554 VTAIL.n320 B 0.030021f
C555 VTAIL.n321 B 0.016132f
C556 VTAIL.n322 B 0.017081f
C557 VTAIL.n323 B 0.03813f
C558 VTAIL.n324 B 0.03813f
C559 VTAIL.n325 B 0.017081f
C560 VTAIL.n326 B 0.016132f
C561 VTAIL.n327 B 0.030021f
C562 VTAIL.n328 B 0.030021f
C563 VTAIL.n329 B 0.016132f
C564 VTAIL.n330 B 0.016132f
C565 VTAIL.n331 B 0.017081f
C566 VTAIL.n332 B 0.03813f
C567 VTAIL.n333 B 0.03813f
C568 VTAIL.n334 B 0.03813f
C569 VTAIL.n335 B 0.016606f
C570 VTAIL.n336 B 0.016132f
C571 VTAIL.n337 B 0.030021f
C572 VTAIL.n338 B 0.030021f
C573 VTAIL.n339 B 0.016132f
C574 VTAIL.n340 B 0.017081f
C575 VTAIL.n341 B 0.03813f
C576 VTAIL.n342 B 0.03813f
C577 VTAIL.n343 B 0.017081f
C578 VTAIL.n344 B 0.016132f
C579 VTAIL.n345 B 0.030021f
C580 VTAIL.n346 B 0.030021f
C581 VTAIL.n347 B 0.016132f
C582 VTAIL.n348 B 0.017081f
C583 VTAIL.n349 B 0.03813f
C584 VTAIL.n350 B 0.03813f
C585 VTAIL.n351 B 0.017081f
C586 VTAIL.n352 B 0.016132f
C587 VTAIL.n353 B 0.030021f
C588 VTAIL.n354 B 0.030021f
C589 VTAIL.n355 B 0.016132f
C590 VTAIL.n356 B 0.017081f
C591 VTAIL.n357 B 0.03813f
C592 VTAIL.n358 B 0.03813f
C593 VTAIL.n359 B 0.017081f
C594 VTAIL.n360 B 0.016132f
C595 VTAIL.n361 B 0.030021f
C596 VTAIL.n362 B 0.030021f
C597 VTAIL.n363 B 0.016132f
C598 VTAIL.n364 B 0.017081f
C599 VTAIL.n365 B 0.03813f
C600 VTAIL.n366 B 0.03813f
C601 VTAIL.n367 B 0.017081f
C602 VTAIL.n368 B 0.016132f
C603 VTAIL.n369 B 0.030021f
C604 VTAIL.n370 B 0.078824f
C605 VTAIL.n371 B 0.016132f
C606 VTAIL.n372 B 0.017081f
C607 VTAIL.n373 B 0.075023f
C608 VTAIL.n374 B 0.064781f
C609 VTAIL.n375 B 1.9032f
C610 VDD2.n0 B 0.016778f
C611 VDD2.n1 B 0.037751f
C612 VDD2.n2 B 0.016911f
C613 VDD2.n3 B 0.029722f
C614 VDD2.n4 B 0.015971f
C615 VDD2.n5 B 0.037751f
C616 VDD2.n6 B 0.016911f
C617 VDD2.n7 B 0.029722f
C618 VDD2.n8 B 0.015971f
C619 VDD2.n9 B 0.037751f
C620 VDD2.n10 B 0.016911f
C621 VDD2.n11 B 0.029722f
C622 VDD2.n12 B 0.015971f
C623 VDD2.n13 B 0.037751f
C624 VDD2.n14 B 0.016911f
C625 VDD2.n15 B 0.029722f
C626 VDD2.n16 B 0.015971f
C627 VDD2.n17 B 0.037751f
C628 VDD2.n18 B 0.016441f
C629 VDD2.n19 B 0.029722f
C630 VDD2.n20 B 0.016911f
C631 VDD2.n21 B 0.037751f
C632 VDD2.n22 B 0.016911f
C633 VDD2.n23 B 0.029722f
C634 VDD2.n24 B 0.015971f
C635 VDD2.n25 B 0.037751f
C636 VDD2.n26 B 0.016911f
C637 VDD2.n27 B 2.11681f
C638 VDD2.n28 B 0.015971f
C639 VDD2.t3 B 0.064506f
C640 VDD2.n29 B 0.267582f
C641 VDD2.n30 B 0.026687f
C642 VDD2.n31 B 0.028313f
C643 VDD2.n32 B 0.037751f
C644 VDD2.n33 B 0.016911f
C645 VDD2.n34 B 0.015971f
C646 VDD2.n35 B 0.029722f
C647 VDD2.n36 B 0.029722f
C648 VDD2.n37 B 0.015971f
C649 VDD2.n38 B 0.016911f
C650 VDD2.n39 B 0.037751f
C651 VDD2.n40 B 0.037751f
C652 VDD2.n41 B 0.016911f
C653 VDD2.n42 B 0.015971f
C654 VDD2.n43 B 0.029722f
C655 VDD2.n44 B 0.029722f
C656 VDD2.n45 B 0.015971f
C657 VDD2.n46 B 0.015971f
C658 VDD2.n47 B 0.016911f
C659 VDD2.n48 B 0.037751f
C660 VDD2.n49 B 0.037751f
C661 VDD2.n50 B 0.037751f
C662 VDD2.n51 B 0.016441f
C663 VDD2.n52 B 0.015971f
C664 VDD2.n53 B 0.029722f
C665 VDD2.n54 B 0.029722f
C666 VDD2.n55 B 0.015971f
C667 VDD2.n56 B 0.016911f
C668 VDD2.n57 B 0.037751f
C669 VDD2.n58 B 0.037751f
C670 VDD2.n59 B 0.016911f
C671 VDD2.n60 B 0.015971f
C672 VDD2.n61 B 0.029722f
C673 VDD2.n62 B 0.029722f
C674 VDD2.n63 B 0.015971f
C675 VDD2.n64 B 0.016911f
C676 VDD2.n65 B 0.037751f
C677 VDD2.n66 B 0.037751f
C678 VDD2.n67 B 0.016911f
C679 VDD2.n68 B 0.015971f
C680 VDD2.n69 B 0.029722f
C681 VDD2.n70 B 0.029722f
C682 VDD2.n71 B 0.015971f
C683 VDD2.n72 B 0.016911f
C684 VDD2.n73 B 0.037751f
C685 VDD2.n74 B 0.037751f
C686 VDD2.n75 B 0.016911f
C687 VDD2.n76 B 0.015971f
C688 VDD2.n77 B 0.029722f
C689 VDD2.n78 B 0.029722f
C690 VDD2.n79 B 0.015971f
C691 VDD2.n80 B 0.016911f
C692 VDD2.n81 B 0.037751f
C693 VDD2.n82 B 0.037751f
C694 VDD2.n83 B 0.016911f
C695 VDD2.n84 B 0.015971f
C696 VDD2.n85 B 0.029722f
C697 VDD2.n86 B 0.07804f
C698 VDD2.n87 B 0.015971f
C699 VDD2.n88 B 0.016911f
C700 VDD2.n89 B 0.074277f
C701 VDD2.n90 B 0.085195f
C702 VDD2.t2 B 0.391535f
C703 VDD2.t1 B 0.391535f
C704 VDD2.n91 B 3.56941f
C705 VDD2.n92 B 2.29335f
C706 VDD2.n93 B 0.016778f
C707 VDD2.n94 B 0.037751f
C708 VDD2.n95 B 0.016911f
C709 VDD2.n96 B 0.029722f
C710 VDD2.n97 B 0.015971f
C711 VDD2.n98 B 0.037751f
C712 VDD2.n99 B 0.016911f
C713 VDD2.n100 B 0.029722f
C714 VDD2.n101 B 0.015971f
C715 VDD2.n102 B 0.037751f
C716 VDD2.n103 B 0.016911f
C717 VDD2.n104 B 0.029722f
C718 VDD2.n105 B 0.015971f
C719 VDD2.n106 B 0.037751f
C720 VDD2.n107 B 0.016911f
C721 VDD2.n108 B 0.029722f
C722 VDD2.n109 B 0.015971f
C723 VDD2.n110 B 0.037751f
C724 VDD2.n111 B 0.016441f
C725 VDD2.n112 B 0.029722f
C726 VDD2.n113 B 0.016441f
C727 VDD2.n114 B 0.015971f
C728 VDD2.n115 B 0.037751f
C729 VDD2.n116 B 0.037751f
C730 VDD2.n117 B 0.016911f
C731 VDD2.n118 B 0.029722f
C732 VDD2.n119 B 0.015971f
C733 VDD2.n120 B 0.037751f
C734 VDD2.n121 B 0.016911f
C735 VDD2.n122 B 2.11681f
C736 VDD2.n123 B 0.015971f
C737 VDD2.t5 B 0.064506f
C738 VDD2.n124 B 0.267582f
C739 VDD2.n125 B 0.026687f
C740 VDD2.n126 B 0.028313f
C741 VDD2.n127 B 0.037751f
C742 VDD2.n128 B 0.016911f
C743 VDD2.n129 B 0.015971f
C744 VDD2.n130 B 0.029722f
C745 VDD2.n131 B 0.029722f
C746 VDD2.n132 B 0.015971f
C747 VDD2.n133 B 0.016911f
C748 VDD2.n134 B 0.037751f
C749 VDD2.n135 B 0.037751f
C750 VDD2.n136 B 0.016911f
C751 VDD2.n137 B 0.015971f
C752 VDD2.n138 B 0.029722f
C753 VDD2.n139 B 0.029722f
C754 VDD2.n140 B 0.015971f
C755 VDD2.n141 B 0.016911f
C756 VDD2.n142 B 0.037751f
C757 VDD2.n143 B 0.037751f
C758 VDD2.n144 B 0.016911f
C759 VDD2.n145 B 0.015971f
C760 VDD2.n146 B 0.029722f
C761 VDD2.n147 B 0.029722f
C762 VDD2.n148 B 0.015971f
C763 VDD2.n149 B 0.016911f
C764 VDD2.n150 B 0.037751f
C765 VDD2.n151 B 0.037751f
C766 VDD2.n152 B 0.016911f
C767 VDD2.n153 B 0.015971f
C768 VDD2.n154 B 0.029722f
C769 VDD2.n155 B 0.029722f
C770 VDD2.n156 B 0.015971f
C771 VDD2.n157 B 0.016911f
C772 VDD2.n158 B 0.037751f
C773 VDD2.n159 B 0.037751f
C774 VDD2.n160 B 0.016911f
C775 VDD2.n161 B 0.015971f
C776 VDD2.n162 B 0.029722f
C777 VDD2.n163 B 0.029722f
C778 VDD2.n164 B 0.015971f
C779 VDD2.n165 B 0.016911f
C780 VDD2.n166 B 0.037751f
C781 VDD2.n167 B 0.037751f
C782 VDD2.n168 B 0.016911f
C783 VDD2.n169 B 0.015971f
C784 VDD2.n170 B 0.029722f
C785 VDD2.n171 B 0.029722f
C786 VDD2.n172 B 0.015971f
C787 VDD2.n173 B 0.016911f
C788 VDD2.n174 B 0.037751f
C789 VDD2.n175 B 0.037751f
C790 VDD2.n176 B 0.016911f
C791 VDD2.n177 B 0.015971f
C792 VDD2.n178 B 0.029722f
C793 VDD2.n179 B 0.07804f
C794 VDD2.n180 B 0.015971f
C795 VDD2.n181 B 0.016911f
C796 VDD2.n182 B 0.074277f
C797 VDD2.n183 B 0.084632f
C798 VDD2.n184 B 2.71391f
C799 VDD2.t4 B 0.391535f
C800 VDD2.t0 B 0.391535f
C801 VDD2.n185 B 3.56938f
C802 VN.t1 B 0.685789f
C803 VN.n0 B 0.279458f
C804 VN.t0 B 0.679141f
C805 VN.n1 B 0.261224f
C806 VN.t2 B 0.685789f
C807 VN.n2 B 0.279371f
C808 VN.n3 B 0.120867f
C809 VN.t3 B 0.685789f
C810 VN.n4 B 0.279458f
C811 VN.t5 B 0.685789f
C812 VN.t4 B 0.679141f
C813 VN.n5 B 0.261224f
C814 VN.n6 B 0.279371f
C815 VN.n7 B 2.70124f
.ends

