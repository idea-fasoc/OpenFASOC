* NGSPICE file created from diff_pair_sample_0151.ext - technology: sky130A

.subckt diff_pair_sample_0151 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t7 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X1 B.t11 B.t9 B.t10 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0 ps=0 w=3.88 l=2.2
X2 VTAIL.t3 VP.t0 VDD1.t7 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0.6402 ps=4.21 w=3.88 l=2.2
X3 VTAIL.t4 VP.t1 VDD1.t6 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X4 VTAIL.t13 VN.t1 VDD2.t3 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0.6402 ps=4.21 w=3.88 l=2.2
X5 VTAIL.t2 VP.t2 VDD1.t5 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0.6402 ps=4.21 w=3.88 l=2.2
X6 B.t8 B.t6 B.t7 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0 ps=0 w=3.88 l=2.2
X7 VDD2.t0 VN.t2 VTAIL.t12 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=1.5132 ps=8.54 w=3.88 l=2.2
X8 VDD1.t4 VP.t3 VTAIL.t1 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=1.5132 ps=8.54 w=3.88 l=2.2
X9 VDD2.t1 VN.t3 VTAIL.t11 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X10 VTAIL.t0 VP.t4 VDD1.t3 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X11 VDD1.t2 VP.t5 VTAIL.t5 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X12 VDD2.t2 VN.t4 VTAIL.t10 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X13 VDD2.t4 VN.t5 VTAIL.t9 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=1.5132 ps=8.54 w=3.88 l=2.2
X14 VTAIL.t8 VN.t6 VDD2.t5 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0.6402 ps=4.21 w=3.88 l=2.2
X15 B.t5 B.t3 B.t4 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0 ps=0 w=3.88 l=2.2
X16 VDD1.t1 VP.t6 VTAIL.t15 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=1.5132 ps=8.54 w=3.88 l=2.2
X17 VDD1.t0 VP.t7 VTAIL.t6 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
X18 B.t2 B.t0 B.t1 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=1.5132 pd=8.54 as=0 ps=0 w=3.88 l=2.2
X19 VTAIL.t7 VN.t7 VDD2.t6 w_n3500_n1744# sky130_fd_pr__pfet_01v8 ad=0.6402 pd=4.21 as=0.6402 ps=4.21 w=3.88 l=2.2
R0 VN.n47 VN.n25 161.3
R1 VN.n46 VN.n45 161.3
R2 VN.n44 VN.n26 161.3
R3 VN.n43 VN.n42 161.3
R4 VN.n41 VN.n27 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n28 161.3
R7 VN.n36 VN.n35 161.3
R8 VN.n34 VN.n29 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n22 VN.n0 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n1 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n2 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n12 VN.n3 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n24 VN.n23 96.3991
R21 VN.n49 VN.n48 96.3991
R22 VN.n6 VN.t6 75.2438
R23 VN.n31 VN.t2 75.2438
R24 VN.n6 VN.n5 58.6104
R25 VN.n31 VN.n30 58.6104
R26 VN.n21 VN.n1 43.4833
R27 VN.n46 VN.n26 43.4833
R28 VN VN.n49 43.1421
R29 VN.n5 VN.t3 42.5041
R30 VN.n15 VN.t7 42.5041
R31 VN.n23 VN.t5 42.5041
R32 VN.n30 VN.t0 42.5041
R33 VN.n40 VN.t4 42.5041
R34 VN.n48 VN.t1 42.5041
R35 VN.n10 VN.n9 40.577
R36 VN.n10 VN.n3 40.577
R37 VN.n35 VN.n34 40.577
R38 VN.n35 VN.n28 40.577
R39 VN.n17 VN.n1 37.6707
R40 VN.n42 VN.n26 37.6707
R41 VN.n9 VN.n8 24.5923
R42 VN.n14 VN.n3 24.5923
R43 VN.n17 VN.n16 24.5923
R44 VN.n22 VN.n21 24.5923
R45 VN.n34 VN.n33 24.5923
R46 VN.n42 VN.n41 24.5923
R47 VN.n39 VN.n28 24.5923
R48 VN.n47 VN.n46 24.5923
R49 VN.n23 VN.n22 14.5097
R50 VN.n48 VN.n47 14.5097
R51 VN.n8 VN.n5 13.0342
R52 VN.n15 VN.n14 13.0342
R53 VN.n33 VN.n30 13.0342
R54 VN.n40 VN.n39 13.0342
R55 VN.n16 VN.n15 11.5587
R56 VN.n41 VN.n40 11.5587
R57 VN.n32 VN.n31 9.48651
R58 VN.n7 VN.n6 9.48651
R59 VN.n49 VN.n25 0.278335
R60 VN.n24 VN.n0 0.278335
R61 VN.n45 VN.n25 0.189894
R62 VN.n45 VN.n44 0.189894
R63 VN.n44 VN.n43 0.189894
R64 VN.n43 VN.n27 0.189894
R65 VN.n38 VN.n27 0.189894
R66 VN.n38 VN.n37 0.189894
R67 VN.n37 VN.n36 0.189894
R68 VN.n36 VN.n29 0.189894
R69 VN.n32 VN.n29 0.189894
R70 VN.n7 VN.n4 0.189894
R71 VN.n11 VN.n4 0.189894
R72 VN.n12 VN.n11 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n13 VN.n2 0.189894
R75 VN.n18 VN.n2 0.189894
R76 VN.n19 VN.n18 0.189894
R77 VN.n20 VN.n19 0.189894
R78 VN.n20 VN.n0 0.189894
R79 VN VN.n24 0.153485
R80 VDD2.n2 VDD2.n1 115.379
R81 VDD2.n2 VDD2.n0 115.379
R82 VDD2 VDD2.n5 115.376
R83 VDD2.n4 VDD2.n3 114.344
R84 VDD2.n4 VDD2.n2 36.8748
R85 VDD2.n5 VDD2.t7 8.37808
R86 VDD2.n5 VDD2.t0 8.37808
R87 VDD2.n3 VDD2.t3 8.37808
R88 VDD2.n3 VDD2.t2 8.37808
R89 VDD2.n1 VDD2.t6 8.37808
R90 VDD2.n1 VDD2.t4 8.37808
R91 VDD2.n0 VDD2.t5 8.37808
R92 VDD2.n0 VDD2.t1 8.37808
R93 VDD2 VDD2.n4 1.14921
R94 VTAIL.n162 VTAIL.n148 756.745
R95 VTAIL.n16 VTAIL.n2 756.745
R96 VTAIL.n36 VTAIL.n22 756.745
R97 VTAIL.n58 VTAIL.n44 756.745
R98 VTAIL.n142 VTAIL.n128 756.745
R99 VTAIL.n120 VTAIL.n106 756.745
R100 VTAIL.n100 VTAIL.n86 756.745
R101 VTAIL.n78 VTAIL.n64 756.745
R102 VTAIL.n155 VTAIL.n154 585
R103 VTAIL.n152 VTAIL.n151 585
R104 VTAIL.n161 VTAIL.n160 585
R105 VTAIL.n163 VTAIL.n162 585
R106 VTAIL.n9 VTAIL.n8 585
R107 VTAIL.n6 VTAIL.n5 585
R108 VTAIL.n15 VTAIL.n14 585
R109 VTAIL.n17 VTAIL.n16 585
R110 VTAIL.n29 VTAIL.n28 585
R111 VTAIL.n26 VTAIL.n25 585
R112 VTAIL.n35 VTAIL.n34 585
R113 VTAIL.n37 VTAIL.n36 585
R114 VTAIL.n51 VTAIL.n50 585
R115 VTAIL.n48 VTAIL.n47 585
R116 VTAIL.n57 VTAIL.n56 585
R117 VTAIL.n59 VTAIL.n58 585
R118 VTAIL.n143 VTAIL.n142 585
R119 VTAIL.n141 VTAIL.n140 585
R120 VTAIL.n132 VTAIL.n131 585
R121 VTAIL.n135 VTAIL.n134 585
R122 VTAIL.n121 VTAIL.n120 585
R123 VTAIL.n119 VTAIL.n118 585
R124 VTAIL.n110 VTAIL.n109 585
R125 VTAIL.n113 VTAIL.n112 585
R126 VTAIL.n101 VTAIL.n100 585
R127 VTAIL.n99 VTAIL.n98 585
R128 VTAIL.n90 VTAIL.n89 585
R129 VTAIL.n93 VTAIL.n92 585
R130 VTAIL.n79 VTAIL.n78 585
R131 VTAIL.n77 VTAIL.n76 585
R132 VTAIL.n68 VTAIL.n67 585
R133 VTAIL.n71 VTAIL.n70 585
R134 VTAIL.t9 VTAIL.n153 330.707
R135 VTAIL.t8 VTAIL.n7 330.707
R136 VTAIL.t15 VTAIL.n27 330.707
R137 VTAIL.t2 VTAIL.n49 330.707
R138 VTAIL.t1 VTAIL.n133 330.707
R139 VTAIL.t3 VTAIL.n111 330.707
R140 VTAIL.t12 VTAIL.n91 330.707
R141 VTAIL.t13 VTAIL.n69 330.707
R142 VTAIL.n154 VTAIL.n151 171.744
R143 VTAIL.n161 VTAIL.n151 171.744
R144 VTAIL.n162 VTAIL.n161 171.744
R145 VTAIL.n8 VTAIL.n5 171.744
R146 VTAIL.n15 VTAIL.n5 171.744
R147 VTAIL.n16 VTAIL.n15 171.744
R148 VTAIL.n28 VTAIL.n25 171.744
R149 VTAIL.n35 VTAIL.n25 171.744
R150 VTAIL.n36 VTAIL.n35 171.744
R151 VTAIL.n50 VTAIL.n47 171.744
R152 VTAIL.n57 VTAIL.n47 171.744
R153 VTAIL.n58 VTAIL.n57 171.744
R154 VTAIL.n142 VTAIL.n141 171.744
R155 VTAIL.n141 VTAIL.n131 171.744
R156 VTAIL.n134 VTAIL.n131 171.744
R157 VTAIL.n120 VTAIL.n119 171.744
R158 VTAIL.n119 VTAIL.n109 171.744
R159 VTAIL.n112 VTAIL.n109 171.744
R160 VTAIL.n100 VTAIL.n99 171.744
R161 VTAIL.n99 VTAIL.n89 171.744
R162 VTAIL.n92 VTAIL.n89 171.744
R163 VTAIL.n78 VTAIL.n77 171.744
R164 VTAIL.n77 VTAIL.n67 171.744
R165 VTAIL.n70 VTAIL.n67 171.744
R166 VTAIL.n127 VTAIL.n126 97.6653
R167 VTAIL.n85 VTAIL.n84 97.6653
R168 VTAIL.n1 VTAIL.n0 97.6651
R169 VTAIL.n43 VTAIL.n42 97.6651
R170 VTAIL.n154 VTAIL.t9 85.8723
R171 VTAIL.n8 VTAIL.t8 85.8723
R172 VTAIL.n28 VTAIL.t15 85.8723
R173 VTAIL.n50 VTAIL.t2 85.8723
R174 VTAIL.n134 VTAIL.t1 85.8723
R175 VTAIL.n112 VTAIL.t3 85.8723
R176 VTAIL.n92 VTAIL.t12 85.8723
R177 VTAIL.n70 VTAIL.t13 85.8723
R178 VTAIL.n167 VTAIL.n166 32.9611
R179 VTAIL.n21 VTAIL.n20 32.9611
R180 VTAIL.n41 VTAIL.n40 32.9611
R181 VTAIL.n63 VTAIL.n62 32.9611
R182 VTAIL.n147 VTAIL.n146 32.9611
R183 VTAIL.n125 VTAIL.n124 32.9611
R184 VTAIL.n105 VTAIL.n104 32.9611
R185 VTAIL.n83 VTAIL.n82 32.9611
R186 VTAIL.n167 VTAIL.n147 17.8927
R187 VTAIL.n83 VTAIL.n63 17.8927
R188 VTAIL.n155 VTAIL.n153 16.3201
R189 VTAIL.n9 VTAIL.n7 16.3201
R190 VTAIL.n29 VTAIL.n27 16.3201
R191 VTAIL.n51 VTAIL.n49 16.3201
R192 VTAIL.n135 VTAIL.n133 16.3201
R193 VTAIL.n113 VTAIL.n111 16.3201
R194 VTAIL.n93 VTAIL.n91 16.3201
R195 VTAIL.n71 VTAIL.n69 16.3201
R196 VTAIL.n156 VTAIL.n152 12.8005
R197 VTAIL.n10 VTAIL.n6 12.8005
R198 VTAIL.n30 VTAIL.n26 12.8005
R199 VTAIL.n52 VTAIL.n48 12.8005
R200 VTAIL.n136 VTAIL.n132 12.8005
R201 VTAIL.n114 VTAIL.n110 12.8005
R202 VTAIL.n94 VTAIL.n90 12.8005
R203 VTAIL.n72 VTAIL.n68 12.8005
R204 VTAIL.n160 VTAIL.n159 12.0247
R205 VTAIL.n14 VTAIL.n13 12.0247
R206 VTAIL.n34 VTAIL.n33 12.0247
R207 VTAIL.n56 VTAIL.n55 12.0247
R208 VTAIL.n140 VTAIL.n139 12.0247
R209 VTAIL.n118 VTAIL.n117 12.0247
R210 VTAIL.n98 VTAIL.n97 12.0247
R211 VTAIL.n76 VTAIL.n75 12.0247
R212 VTAIL.n163 VTAIL.n150 11.249
R213 VTAIL.n17 VTAIL.n4 11.249
R214 VTAIL.n37 VTAIL.n24 11.249
R215 VTAIL.n59 VTAIL.n46 11.249
R216 VTAIL.n143 VTAIL.n130 11.249
R217 VTAIL.n121 VTAIL.n108 11.249
R218 VTAIL.n101 VTAIL.n88 11.249
R219 VTAIL.n79 VTAIL.n66 11.249
R220 VTAIL.n164 VTAIL.n148 10.4732
R221 VTAIL.n18 VTAIL.n2 10.4732
R222 VTAIL.n38 VTAIL.n22 10.4732
R223 VTAIL.n60 VTAIL.n44 10.4732
R224 VTAIL.n144 VTAIL.n128 10.4732
R225 VTAIL.n122 VTAIL.n106 10.4732
R226 VTAIL.n102 VTAIL.n86 10.4732
R227 VTAIL.n80 VTAIL.n64 10.4732
R228 VTAIL.n166 VTAIL.n165 9.45567
R229 VTAIL.n20 VTAIL.n19 9.45567
R230 VTAIL.n40 VTAIL.n39 9.45567
R231 VTAIL.n62 VTAIL.n61 9.45567
R232 VTAIL.n146 VTAIL.n145 9.45567
R233 VTAIL.n124 VTAIL.n123 9.45567
R234 VTAIL.n104 VTAIL.n103 9.45567
R235 VTAIL.n82 VTAIL.n81 9.45567
R236 VTAIL.n165 VTAIL.n164 9.3005
R237 VTAIL.n150 VTAIL.n149 9.3005
R238 VTAIL.n159 VTAIL.n158 9.3005
R239 VTAIL.n157 VTAIL.n156 9.3005
R240 VTAIL.n19 VTAIL.n18 9.3005
R241 VTAIL.n4 VTAIL.n3 9.3005
R242 VTAIL.n13 VTAIL.n12 9.3005
R243 VTAIL.n11 VTAIL.n10 9.3005
R244 VTAIL.n39 VTAIL.n38 9.3005
R245 VTAIL.n24 VTAIL.n23 9.3005
R246 VTAIL.n33 VTAIL.n32 9.3005
R247 VTAIL.n31 VTAIL.n30 9.3005
R248 VTAIL.n61 VTAIL.n60 9.3005
R249 VTAIL.n46 VTAIL.n45 9.3005
R250 VTAIL.n55 VTAIL.n54 9.3005
R251 VTAIL.n53 VTAIL.n52 9.3005
R252 VTAIL.n145 VTAIL.n144 9.3005
R253 VTAIL.n130 VTAIL.n129 9.3005
R254 VTAIL.n139 VTAIL.n138 9.3005
R255 VTAIL.n137 VTAIL.n136 9.3005
R256 VTAIL.n123 VTAIL.n122 9.3005
R257 VTAIL.n108 VTAIL.n107 9.3005
R258 VTAIL.n117 VTAIL.n116 9.3005
R259 VTAIL.n115 VTAIL.n114 9.3005
R260 VTAIL.n103 VTAIL.n102 9.3005
R261 VTAIL.n88 VTAIL.n87 9.3005
R262 VTAIL.n97 VTAIL.n96 9.3005
R263 VTAIL.n95 VTAIL.n94 9.3005
R264 VTAIL.n81 VTAIL.n80 9.3005
R265 VTAIL.n66 VTAIL.n65 9.3005
R266 VTAIL.n75 VTAIL.n74 9.3005
R267 VTAIL.n73 VTAIL.n72 9.3005
R268 VTAIL.n0 VTAIL.t11 8.37808
R269 VTAIL.n0 VTAIL.t7 8.37808
R270 VTAIL.n42 VTAIL.t6 8.37808
R271 VTAIL.n42 VTAIL.t0 8.37808
R272 VTAIL.n126 VTAIL.t5 8.37808
R273 VTAIL.n126 VTAIL.t4 8.37808
R274 VTAIL.n84 VTAIL.t10 8.37808
R275 VTAIL.n84 VTAIL.t14 8.37808
R276 VTAIL.n157 VTAIL.n153 3.78097
R277 VTAIL.n11 VTAIL.n7 3.78097
R278 VTAIL.n31 VTAIL.n27 3.78097
R279 VTAIL.n53 VTAIL.n49 3.78097
R280 VTAIL.n137 VTAIL.n133 3.78097
R281 VTAIL.n115 VTAIL.n111 3.78097
R282 VTAIL.n95 VTAIL.n91 3.78097
R283 VTAIL.n73 VTAIL.n69 3.78097
R284 VTAIL.n166 VTAIL.n148 3.49141
R285 VTAIL.n20 VTAIL.n2 3.49141
R286 VTAIL.n40 VTAIL.n22 3.49141
R287 VTAIL.n62 VTAIL.n44 3.49141
R288 VTAIL.n146 VTAIL.n128 3.49141
R289 VTAIL.n124 VTAIL.n106 3.49141
R290 VTAIL.n104 VTAIL.n86 3.49141
R291 VTAIL.n82 VTAIL.n64 3.49141
R292 VTAIL.n164 VTAIL.n163 2.71565
R293 VTAIL.n18 VTAIL.n17 2.71565
R294 VTAIL.n38 VTAIL.n37 2.71565
R295 VTAIL.n60 VTAIL.n59 2.71565
R296 VTAIL.n144 VTAIL.n143 2.71565
R297 VTAIL.n122 VTAIL.n121 2.71565
R298 VTAIL.n102 VTAIL.n101 2.71565
R299 VTAIL.n80 VTAIL.n79 2.71565
R300 VTAIL.n85 VTAIL.n83 2.18153
R301 VTAIL.n105 VTAIL.n85 2.18153
R302 VTAIL.n127 VTAIL.n125 2.18153
R303 VTAIL.n147 VTAIL.n127 2.18153
R304 VTAIL.n63 VTAIL.n43 2.18153
R305 VTAIL.n43 VTAIL.n41 2.18153
R306 VTAIL.n21 VTAIL.n1 2.18153
R307 VTAIL VTAIL.n167 2.12334
R308 VTAIL.n160 VTAIL.n150 1.93989
R309 VTAIL.n14 VTAIL.n4 1.93989
R310 VTAIL.n34 VTAIL.n24 1.93989
R311 VTAIL.n56 VTAIL.n46 1.93989
R312 VTAIL.n140 VTAIL.n130 1.93989
R313 VTAIL.n118 VTAIL.n108 1.93989
R314 VTAIL.n98 VTAIL.n88 1.93989
R315 VTAIL.n76 VTAIL.n66 1.93989
R316 VTAIL.n159 VTAIL.n152 1.16414
R317 VTAIL.n13 VTAIL.n6 1.16414
R318 VTAIL.n33 VTAIL.n26 1.16414
R319 VTAIL.n55 VTAIL.n48 1.16414
R320 VTAIL.n139 VTAIL.n132 1.16414
R321 VTAIL.n117 VTAIL.n110 1.16414
R322 VTAIL.n97 VTAIL.n90 1.16414
R323 VTAIL.n75 VTAIL.n68 1.16414
R324 VTAIL.n125 VTAIL.n105 0.470328
R325 VTAIL.n41 VTAIL.n21 0.470328
R326 VTAIL.n156 VTAIL.n155 0.388379
R327 VTAIL.n10 VTAIL.n9 0.388379
R328 VTAIL.n30 VTAIL.n29 0.388379
R329 VTAIL.n52 VTAIL.n51 0.388379
R330 VTAIL.n136 VTAIL.n135 0.388379
R331 VTAIL.n114 VTAIL.n113 0.388379
R332 VTAIL.n94 VTAIL.n93 0.388379
R333 VTAIL.n72 VTAIL.n71 0.388379
R334 VTAIL.n158 VTAIL.n157 0.155672
R335 VTAIL.n158 VTAIL.n149 0.155672
R336 VTAIL.n165 VTAIL.n149 0.155672
R337 VTAIL.n12 VTAIL.n11 0.155672
R338 VTAIL.n12 VTAIL.n3 0.155672
R339 VTAIL.n19 VTAIL.n3 0.155672
R340 VTAIL.n32 VTAIL.n31 0.155672
R341 VTAIL.n32 VTAIL.n23 0.155672
R342 VTAIL.n39 VTAIL.n23 0.155672
R343 VTAIL.n54 VTAIL.n53 0.155672
R344 VTAIL.n54 VTAIL.n45 0.155672
R345 VTAIL.n61 VTAIL.n45 0.155672
R346 VTAIL.n145 VTAIL.n129 0.155672
R347 VTAIL.n138 VTAIL.n129 0.155672
R348 VTAIL.n138 VTAIL.n137 0.155672
R349 VTAIL.n123 VTAIL.n107 0.155672
R350 VTAIL.n116 VTAIL.n107 0.155672
R351 VTAIL.n116 VTAIL.n115 0.155672
R352 VTAIL.n103 VTAIL.n87 0.155672
R353 VTAIL.n96 VTAIL.n87 0.155672
R354 VTAIL.n96 VTAIL.n95 0.155672
R355 VTAIL.n81 VTAIL.n65 0.155672
R356 VTAIL.n74 VTAIL.n65 0.155672
R357 VTAIL.n74 VTAIL.n73 0.155672
R358 VTAIL VTAIL.n1 0.0586897
R359 B.n281 B.n280 585
R360 B.n279 B.n98 585
R361 B.n278 B.n277 585
R362 B.n276 B.n99 585
R363 B.n275 B.n274 585
R364 B.n273 B.n100 585
R365 B.n272 B.n271 585
R366 B.n270 B.n101 585
R367 B.n269 B.n268 585
R368 B.n267 B.n102 585
R369 B.n266 B.n265 585
R370 B.n264 B.n103 585
R371 B.n263 B.n262 585
R372 B.n261 B.n104 585
R373 B.n260 B.n259 585
R374 B.n258 B.n105 585
R375 B.n257 B.n256 585
R376 B.n255 B.n106 585
R377 B.n254 B.n253 585
R378 B.n249 B.n107 585
R379 B.n248 B.n247 585
R380 B.n246 B.n108 585
R381 B.n245 B.n244 585
R382 B.n243 B.n109 585
R383 B.n242 B.n241 585
R384 B.n240 B.n110 585
R385 B.n239 B.n238 585
R386 B.n236 B.n111 585
R387 B.n235 B.n234 585
R388 B.n233 B.n114 585
R389 B.n232 B.n231 585
R390 B.n230 B.n115 585
R391 B.n229 B.n228 585
R392 B.n227 B.n116 585
R393 B.n226 B.n225 585
R394 B.n224 B.n117 585
R395 B.n223 B.n222 585
R396 B.n221 B.n118 585
R397 B.n220 B.n219 585
R398 B.n218 B.n119 585
R399 B.n217 B.n216 585
R400 B.n215 B.n120 585
R401 B.n214 B.n213 585
R402 B.n212 B.n121 585
R403 B.n211 B.n210 585
R404 B.n282 B.n97 585
R405 B.n284 B.n283 585
R406 B.n285 B.n96 585
R407 B.n287 B.n286 585
R408 B.n288 B.n95 585
R409 B.n290 B.n289 585
R410 B.n291 B.n94 585
R411 B.n293 B.n292 585
R412 B.n294 B.n93 585
R413 B.n296 B.n295 585
R414 B.n297 B.n92 585
R415 B.n299 B.n298 585
R416 B.n300 B.n91 585
R417 B.n302 B.n301 585
R418 B.n303 B.n90 585
R419 B.n305 B.n304 585
R420 B.n306 B.n89 585
R421 B.n308 B.n307 585
R422 B.n309 B.n88 585
R423 B.n311 B.n310 585
R424 B.n312 B.n87 585
R425 B.n314 B.n313 585
R426 B.n315 B.n86 585
R427 B.n317 B.n316 585
R428 B.n318 B.n85 585
R429 B.n320 B.n319 585
R430 B.n321 B.n84 585
R431 B.n323 B.n322 585
R432 B.n324 B.n83 585
R433 B.n326 B.n325 585
R434 B.n327 B.n82 585
R435 B.n329 B.n328 585
R436 B.n330 B.n81 585
R437 B.n332 B.n331 585
R438 B.n333 B.n80 585
R439 B.n335 B.n334 585
R440 B.n336 B.n79 585
R441 B.n338 B.n337 585
R442 B.n339 B.n78 585
R443 B.n341 B.n340 585
R444 B.n342 B.n77 585
R445 B.n344 B.n343 585
R446 B.n345 B.n76 585
R447 B.n347 B.n346 585
R448 B.n348 B.n75 585
R449 B.n350 B.n349 585
R450 B.n351 B.n74 585
R451 B.n353 B.n352 585
R452 B.n354 B.n73 585
R453 B.n356 B.n355 585
R454 B.n357 B.n72 585
R455 B.n359 B.n358 585
R456 B.n360 B.n71 585
R457 B.n362 B.n361 585
R458 B.n363 B.n70 585
R459 B.n365 B.n364 585
R460 B.n366 B.n69 585
R461 B.n368 B.n367 585
R462 B.n369 B.n68 585
R463 B.n371 B.n370 585
R464 B.n372 B.n67 585
R465 B.n374 B.n373 585
R466 B.n375 B.n66 585
R467 B.n377 B.n376 585
R468 B.n378 B.n65 585
R469 B.n380 B.n379 585
R470 B.n381 B.n64 585
R471 B.n383 B.n382 585
R472 B.n384 B.n63 585
R473 B.n386 B.n385 585
R474 B.n387 B.n62 585
R475 B.n389 B.n388 585
R476 B.n390 B.n61 585
R477 B.n392 B.n391 585
R478 B.n393 B.n60 585
R479 B.n395 B.n394 585
R480 B.n396 B.n59 585
R481 B.n398 B.n397 585
R482 B.n399 B.n58 585
R483 B.n401 B.n400 585
R484 B.n402 B.n57 585
R485 B.n404 B.n403 585
R486 B.n405 B.n56 585
R487 B.n407 B.n406 585
R488 B.n408 B.n55 585
R489 B.n410 B.n409 585
R490 B.n411 B.n54 585
R491 B.n413 B.n412 585
R492 B.n414 B.n53 585
R493 B.n416 B.n415 585
R494 B.n417 B.n52 585
R495 B.n419 B.n418 585
R496 B.n488 B.n487 585
R497 B.n486 B.n25 585
R498 B.n485 B.n484 585
R499 B.n483 B.n26 585
R500 B.n482 B.n481 585
R501 B.n480 B.n27 585
R502 B.n479 B.n478 585
R503 B.n477 B.n28 585
R504 B.n476 B.n475 585
R505 B.n474 B.n29 585
R506 B.n473 B.n472 585
R507 B.n471 B.n30 585
R508 B.n470 B.n469 585
R509 B.n468 B.n31 585
R510 B.n467 B.n466 585
R511 B.n465 B.n32 585
R512 B.n464 B.n463 585
R513 B.n462 B.n33 585
R514 B.n460 B.n459 585
R515 B.n458 B.n36 585
R516 B.n457 B.n456 585
R517 B.n455 B.n37 585
R518 B.n454 B.n453 585
R519 B.n452 B.n38 585
R520 B.n451 B.n450 585
R521 B.n449 B.n39 585
R522 B.n448 B.n447 585
R523 B.n446 B.n445 585
R524 B.n444 B.n43 585
R525 B.n443 B.n442 585
R526 B.n441 B.n44 585
R527 B.n440 B.n439 585
R528 B.n438 B.n45 585
R529 B.n437 B.n436 585
R530 B.n435 B.n46 585
R531 B.n434 B.n433 585
R532 B.n432 B.n47 585
R533 B.n431 B.n430 585
R534 B.n429 B.n48 585
R535 B.n428 B.n427 585
R536 B.n426 B.n49 585
R537 B.n425 B.n424 585
R538 B.n423 B.n50 585
R539 B.n422 B.n421 585
R540 B.n420 B.n51 585
R541 B.n489 B.n24 585
R542 B.n491 B.n490 585
R543 B.n492 B.n23 585
R544 B.n494 B.n493 585
R545 B.n495 B.n22 585
R546 B.n497 B.n496 585
R547 B.n498 B.n21 585
R548 B.n500 B.n499 585
R549 B.n501 B.n20 585
R550 B.n503 B.n502 585
R551 B.n504 B.n19 585
R552 B.n506 B.n505 585
R553 B.n507 B.n18 585
R554 B.n509 B.n508 585
R555 B.n510 B.n17 585
R556 B.n512 B.n511 585
R557 B.n513 B.n16 585
R558 B.n515 B.n514 585
R559 B.n516 B.n15 585
R560 B.n518 B.n517 585
R561 B.n519 B.n14 585
R562 B.n521 B.n520 585
R563 B.n522 B.n13 585
R564 B.n524 B.n523 585
R565 B.n525 B.n12 585
R566 B.n527 B.n526 585
R567 B.n528 B.n11 585
R568 B.n530 B.n529 585
R569 B.n531 B.n10 585
R570 B.n533 B.n532 585
R571 B.n534 B.n9 585
R572 B.n536 B.n535 585
R573 B.n537 B.n8 585
R574 B.n539 B.n538 585
R575 B.n540 B.n7 585
R576 B.n542 B.n541 585
R577 B.n543 B.n6 585
R578 B.n545 B.n544 585
R579 B.n546 B.n5 585
R580 B.n548 B.n547 585
R581 B.n549 B.n4 585
R582 B.n551 B.n550 585
R583 B.n552 B.n3 585
R584 B.n554 B.n553 585
R585 B.n555 B.n0 585
R586 B.n2 B.n1 585
R587 B.n145 B.n144 585
R588 B.n146 B.n143 585
R589 B.n148 B.n147 585
R590 B.n149 B.n142 585
R591 B.n151 B.n150 585
R592 B.n152 B.n141 585
R593 B.n154 B.n153 585
R594 B.n155 B.n140 585
R595 B.n157 B.n156 585
R596 B.n158 B.n139 585
R597 B.n160 B.n159 585
R598 B.n161 B.n138 585
R599 B.n163 B.n162 585
R600 B.n164 B.n137 585
R601 B.n166 B.n165 585
R602 B.n167 B.n136 585
R603 B.n169 B.n168 585
R604 B.n170 B.n135 585
R605 B.n172 B.n171 585
R606 B.n173 B.n134 585
R607 B.n175 B.n174 585
R608 B.n176 B.n133 585
R609 B.n178 B.n177 585
R610 B.n179 B.n132 585
R611 B.n181 B.n180 585
R612 B.n182 B.n131 585
R613 B.n184 B.n183 585
R614 B.n185 B.n130 585
R615 B.n187 B.n186 585
R616 B.n188 B.n129 585
R617 B.n190 B.n189 585
R618 B.n191 B.n128 585
R619 B.n193 B.n192 585
R620 B.n194 B.n127 585
R621 B.n196 B.n195 585
R622 B.n197 B.n126 585
R623 B.n199 B.n198 585
R624 B.n200 B.n125 585
R625 B.n202 B.n201 585
R626 B.n203 B.n124 585
R627 B.n205 B.n204 585
R628 B.n206 B.n123 585
R629 B.n208 B.n207 585
R630 B.n209 B.n122 585
R631 B.n210 B.n209 473.281
R632 B.n280 B.n97 473.281
R633 B.n418 B.n51 473.281
R634 B.n489 B.n488 473.281
R635 B.n250 B.t7 282.368
R636 B.n40 B.t2 282.368
R637 B.n112 B.t4 282.368
R638 B.n34 B.t11 282.368
R639 B.n557 B.n556 256.663
R640 B.n112 B.t3 249.856
R641 B.n250 B.t6 249.856
R642 B.n40 B.t0 249.856
R643 B.n34 B.t9 249.856
R644 B.n556 B.n555 235.042
R645 B.n556 B.n2 235.042
R646 B.n251 B.t8 233.303
R647 B.n41 B.t1 233.303
R648 B.n113 B.t5 233.303
R649 B.n35 B.t10 233.303
R650 B.n210 B.n121 163.367
R651 B.n214 B.n121 163.367
R652 B.n215 B.n214 163.367
R653 B.n216 B.n215 163.367
R654 B.n216 B.n119 163.367
R655 B.n220 B.n119 163.367
R656 B.n221 B.n220 163.367
R657 B.n222 B.n221 163.367
R658 B.n222 B.n117 163.367
R659 B.n226 B.n117 163.367
R660 B.n227 B.n226 163.367
R661 B.n228 B.n227 163.367
R662 B.n228 B.n115 163.367
R663 B.n232 B.n115 163.367
R664 B.n233 B.n232 163.367
R665 B.n234 B.n233 163.367
R666 B.n234 B.n111 163.367
R667 B.n239 B.n111 163.367
R668 B.n240 B.n239 163.367
R669 B.n241 B.n240 163.367
R670 B.n241 B.n109 163.367
R671 B.n245 B.n109 163.367
R672 B.n246 B.n245 163.367
R673 B.n247 B.n246 163.367
R674 B.n247 B.n107 163.367
R675 B.n254 B.n107 163.367
R676 B.n255 B.n254 163.367
R677 B.n256 B.n255 163.367
R678 B.n256 B.n105 163.367
R679 B.n260 B.n105 163.367
R680 B.n261 B.n260 163.367
R681 B.n262 B.n261 163.367
R682 B.n262 B.n103 163.367
R683 B.n266 B.n103 163.367
R684 B.n267 B.n266 163.367
R685 B.n268 B.n267 163.367
R686 B.n268 B.n101 163.367
R687 B.n272 B.n101 163.367
R688 B.n273 B.n272 163.367
R689 B.n274 B.n273 163.367
R690 B.n274 B.n99 163.367
R691 B.n278 B.n99 163.367
R692 B.n279 B.n278 163.367
R693 B.n280 B.n279 163.367
R694 B.n418 B.n417 163.367
R695 B.n417 B.n416 163.367
R696 B.n416 B.n53 163.367
R697 B.n412 B.n53 163.367
R698 B.n412 B.n411 163.367
R699 B.n411 B.n410 163.367
R700 B.n410 B.n55 163.367
R701 B.n406 B.n55 163.367
R702 B.n406 B.n405 163.367
R703 B.n405 B.n404 163.367
R704 B.n404 B.n57 163.367
R705 B.n400 B.n57 163.367
R706 B.n400 B.n399 163.367
R707 B.n399 B.n398 163.367
R708 B.n398 B.n59 163.367
R709 B.n394 B.n59 163.367
R710 B.n394 B.n393 163.367
R711 B.n393 B.n392 163.367
R712 B.n392 B.n61 163.367
R713 B.n388 B.n61 163.367
R714 B.n388 B.n387 163.367
R715 B.n387 B.n386 163.367
R716 B.n386 B.n63 163.367
R717 B.n382 B.n63 163.367
R718 B.n382 B.n381 163.367
R719 B.n381 B.n380 163.367
R720 B.n380 B.n65 163.367
R721 B.n376 B.n65 163.367
R722 B.n376 B.n375 163.367
R723 B.n375 B.n374 163.367
R724 B.n374 B.n67 163.367
R725 B.n370 B.n67 163.367
R726 B.n370 B.n369 163.367
R727 B.n369 B.n368 163.367
R728 B.n368 B.n69 163.367
R729 B.n364 B.n69 163.367
R730 B.n364 B.n363 163.367
R731 B.n363 B.n362 163.367
R732 B.n362 B.n71 163.367
R733 B.n358 B.n71 163.367
R734 B.n358 B.n357 163.367
R735 B.n357 B.n356 163.367
R736 B.n356 B.n73 163.367
R737 B.n352 B.n73 163.367
R738 B.n352 B.n351 163.367
R739 B.n351 B.n350 163.367
R740 B.n350 B.n75 163.367
R741 B.n346 B.n75 163.367
R742 B.n346 B.n345 163.367
R743 B.n345 B.n344 163.367
R744 B.n344 B.n77 163.367
R745 B.n340 B.n77 163.367
R746 B.n340 B.n339 163.367
R747 B.n339 B.n338 163.367
R748 B.n338 B.n79 163.367
R749 B.n334 B.n79 163.367
R750 B.n334 B.n333 163.367
R751 B.n333 B.n332 163.367
R752 B.n332 B.n81 163.367
R753 B.n328 B.n81 163.367
R754 B.n328 B.n327 163.367
R755 B.n327 B.n326 163.367
R756 B.n326 B.n83 163.367
R757 B.n322 B.n83 163.367
R758 B.n322 B.n321 163.367
R759 B.n321 B.n320 163.367
R760 B.n320 B.n85 163.367
R761 B.n316 B.n85 163.367
R762 B.n316 B.n315 163.367
R763 B.n315 B.n314 163.367
R764 B.n314 B.n87 163.367
R765 B.n310 B.n87 163.367
R766 B.n310 B.n309 163.367
R767 B.n309 B.n308 163.367
R768 B.n308 B.n89 163.367
R769 B.n304 B.n89 163.367
R770 B.n304 B.n303 163.367
R771 B.n303 B.n302 163.367
R772 B.n302 B.n91 163.367
R773 B.n298 B.n91 163.367
R774 B.n298 B.n297 163.367
R775 B.n297 B.n296 163.367
R776 B.n296 B.n93 163.367
R777 B.n292 B.n93 163.367
R778 B.n292 B.n291 163.367
R779 B.n291 B.n290 163.367
R780 B.n290 B.n95 163.367
R781 B.n286 B.n95 163.367
R782 B.n286 B.n285 163.367
R783 B.n285 B.n284 163.367
R784 B.n284 B.n97 163.367
R785 B.n488 B.n25 163.367
R786 B.n484 B.n25 163.367
R787 B.n484 B.n483 163.367
R788 B.n483 B.n482 163.367
R789 B.n482 B.n27 163.367
R790 B.n478 B.n27 163.367
R791 B.n478 B.n477 163.367
R792 B.n477 B.n476 163.367
R793 B.n476 B.n29 163.367
R794 B.n472 B.n29 163.367
R795 B.n472 B.n471 163.367
R796 B.n471 B.n470 163.367
R797 B.n470 B.n31 163.367
R798 B.n466 B.n31 163.367
R799 B.n466 B.n465 163.367
R800 B.n465 B.n464 163.367
R801 B.n464 B.n33 163.367
R802 B.n459 B.n33 163.367
R803 B.n459 B.n458 163.367
R804 B.n458 B.n457 163.367
R805 B.n457 B.n37 163.367
R806 B.n453 B.n37 163.367
R807 B.n453 B.n452 163.367
R808 B.n452 B.n451 163.367
R809 B.n451 B.n39 163.367
R810 B.n447 B.n39 163.367
R811 B.n447 B.n446 163.367
R812 B.n446 B.n43 163.367
R813 B.n442 B.n43 163.367
R814 B.n442 B.n441 163.367
R815 B.n441 B.n440 163.367
R816 B.n440 B.n45 163.367
R817 B.n436 B.n45 163.367
R818 B.n436 B.n435 163.367
R819 B.n435 B.n434 163.367
R820 B.n434 B.n47 163.367
R821 B.n430 B.n47 163.367
R822 B.n430 B.n429 163.367
R823 B.n429 B.n428 163.367
R824 B.n428 B.n49 163.367
R825 B.n424 B.n49 163.367
R826 B.n424 B.n423 163.367
R827 B.n423 B.n422 163.367
R828 B.n422 B.n51 163.367
R829 B.n490 B.n489 163.367
R830 B.n490 B.n23 163.367
R831 B.n494 B.n23 163.367
R832 B.n495 B.n494 163.367
R833 B.n496 B.n495 163.367
R834 B.n496 B.n21 163.367
R835 B.n500 B.n21 163.367
R836 B.n501 B.n500 163.367
R837 B.n502 B.n501 163.367
R838 B.n502 B.n19 163.367
R839 B.n506 B.n19 163.367
R840 B.n507 B.n506 163.367
R841 B.n508 B.n507 163.367
R842 B.n508 B.n17 163.367
R843 B.n512 B.n17 163.367
R844 B.n513 B.n512 163.367
R845 B.n514 B.n513 163.367
R846 B.n514 B.n15 163.367
R847 B.n518 B.n15 163.367
R848 B.n519 B.n518 163.367
R849 B.n520 B.n519 163.367
R850 B.n520 B.n13 163.367
R851 B.n524 B.n13 163.367
R852 B.n525 B.n524 163.367
R853 B.n526 B.n525 163.367
R854 B.n526 B.n11 163.367
R855 B.n530 B.n11 163.367
R856 B.n531 B.n530 163.367
R857 B.n532 B.n531 163.367
R858 B.n532 B.n9 163.367
R859 B.n536 B.n9 163.367
R860 B.n537 B.n536 163.367
R861 B.n538 B.n537 163.367
R862 B.n538 B.n7 163.367
R863 B.n542 B.n7 163.367
R864 B.n543 B.n542 163.367
R865 B.n544 B.n543 163.367
R866 B.n544 B.n5 163.367
R867 B.n548 B.n5 163.367
R868 B.n549 B.n548 163.367
R869 B.n550 B.n549 163.367
R870 B.n550 B.n3 163.367
R871 B.n554 B.n3 163.367
R872 B.n555 B.n554 163.367
R873 B.n144 B.n2 163.367
R874 B.n144 B.n143 163.367
R875 B.n148 B.n143 163.367
R876 B.n149 B.n148 163.367
R877 B.n150 B.n149 163.367
R878 B.n150 B.n141 163.367
R879 B.n154 B.n141 163.367
R880 B.n155 B.n154 163.367
R881 B.n156 B.n155 163.367
R882 B.n156 B.n139 163.367
R883 B.n160 B.n139 163.367
R884 B.n161 B.n160 163.367
R885 B.n162 B.n161 163.367
R886 B.n162 B.n137 163.367
R887 B.n166 B.n137 163.367
R888 B.n167 B.n166 163.367
R889 B.n168 B.n167 163.367
R890 B.n168 B.n135 163.367
R891 B.n172 B.n135 163.367
R892 B.n173 B.n172 163.367
R893 B.n174 B.n173 163.367
R894 B.n174 B.n133 163.367
R895 B.n178 B.n133 163.367
R896 B.n179 B.n178 163.367
R897 B.n180 B.n179 163.367
R898 B.n180 B.n131 163.367
R899 B.n184 B.n131 163.367
R900 B.n185 B.n184 163.367
R901 B.n186 B.n185 163.367
R902 B.n186 B.n129 163.367
R903 B.n190 B.n129 163.367
R904 B.n191 B.n190 163.367
R905 B.n192 B.n191 163.367
R906 B.n192 B.n127 163.367
R907 B.n196 B.n127 163.367
R908 B.n197 B.n196 163.367
R909 B.n198 B.n197 163.367
R910 B.n198 B.n125 163.367
R911 B.n202 B.n125 163.367
R912 B.n203 B.n202 163.367
R913 B.n204 B.n203 163.367
R914 B.n204 B.n123 163.367
R915 B.n208 B.n123 163.367
R916 B.n209 B.n208 163.367
R917 B.n237 B.n113 59.5399
R918 B.n252 B.n251 59.5399
R919 B.n42 B.n41 59.5399
R920 B.n461 B.n35 59.5399
R921 B.n113 B.n112 49.0672
R922 B.n251 B.n250 49.0672
R923 B.n41 B.n40 49.0672
R924 B.n35 B.n34 49.0672
R925 B.n487 B.n24 30.7517
R926 B.n420 B.n419 30.7517
R927 B.n211 B.n122 30.7517
R928 B.n282 B.n281 30.7517
R929 B B.n557 18.0485
R930 B.n491 B.n24 10.6151
R931 B.n492 B.n491 10.6151
R932 B.n493 B.n492 10.6151
R933 B.n493 B.n22 10.6151
R934 B.n497 B.n22 10.6151
R935 B.n498 B.n497 10.6151
R936 B.n499 B.n498 10.6151
R937 B.n499 B.n20 10.6151
R938 B.n503 B.n20 10.6151
R939 B.n504 B.n503 10.6151
R940 B.n505 B.n504 10.6151
R941 B.n505 B.n18 10.6151
R942 B.n509 B.n18 10.6151
R943 B.n510 B.n509 10.6151
R944 B.n511 B.n510 10.6151
R945 B.n511 B.n16 10.6151
R946 B.n515 B.n16 10.6151
R947 B.n516 B.n515 10.6151
R948 B.n517 B.n516 10.6151
R949 B.n517 B.n14 10.6151
R950 B.n521 B.n14 10.6151
R951 B.n522 B.n521 10.6151
R952 B.n523 B.n522 10.6151
R953 B.n523 B.n12 10.6151
R954 B.n527 B.n12 10.6151
R955 B.n528 B.n527 10.6151
R956 B.n529 B.n528 10.6151
R957 B.n529 B.n10 10.6151
R958 B.n533 B.n10 10.6151
R959 B.n534 B.n533 10.6151
R960 B.n535 B.n534 10.6151
R961 B.n535 B.n8 10.6151
R962 B.n539 B.n8 10.6151
R963 B.n540 B.n539 10.6151
R964 B.n541 B.n540 10.6151
R965 B.n541 B.n6 10.6151
R966 B.n545 B.n6 10.6151
R967 B.n546 B.n545 10.6151
R968 B.n547 B.n546 10.6151
R969 B.n547 B.n4 10.6151
R970 B.n551 B.n4 10.6151
R971 B.n552 B.n551 10.6151
R972 B.n553 B.n552 10.6151
R973 B.n553 B.n0 10.6151
R974 B.n487 B.n486 10.6151
R975 B.n486 B.n485 10.6151
R976 B.n485 B.n26 10.6151
R977 B.n481 B.n26 10.6151
R978 B.n481 B.n480 10.6151
R979 B.n480 B.n479 10.6151
R980 B.n479 B.n28 10.6151
R981 B.n475 B.n28 10.6151
R982 B.n475 B.n474 10.6151
R983 B.n474 B.n473 10.6151
R984 B.n473 B.n30 10.6151
R985 B.n469 B.n30 10.6151
R986 B.n469 B.n468 10.6151
R987 B.n468 B.n467 10.6151
R988 B.n467 B.n32 10.6151
R989 B.n463 B.n32 10.6151
R990 B.n463 B.n462 10.6151
R991 B.n460 B.n36 10.6151
R992 B.n456 B.n36 10.6151
R993 B.n456 B.n455 10.6151
R994 B.n455 B.n454 10.6151
R995 B.n454 B.n38 10.6151
R996 B.n450 B.n38 10.6151
R997 B.n450 B.n449 10.6151
R998 B.n449 B.n448 10.6151
R999 B.n445 B.n444 10.6151
R1000 B.n444 B.n443 10.6151
R1001 B.n443 B.n44 10.6151
R1002 B.n439 B.n44 10.6151
R1003 B.n439 B.n438 10.6151
R1004 B.n438 B.n437 10.6151
R1005 B.n437 B.n46 10.6151
R1006 B.n433 B.n46 10.6151
R1007 B.n433 B.n432 10.6151
R1008 B.n432 B.n431 10.6151
R1009 B.n431 B.n48 10.6151
R1010 B.n427 B.n48 10.6151
R1011 B.n427 B.n426 10.6151
R1012 B.n426 B.n425 10.6151
R1013 B.n425 B.n50 10.6151
R1014 B.n421 B.n50 10.6151
R1015 B.n421 B.n420 10.6151
R1016 B.n419 B.n52 10.6151
R1017 B.n415 B.n52 10.6151
R1018 B.n415 B.n414 10.6151
R1019 B.n414 B.n413 10.6151
R1020 B.n413 B.n54 10.6151
R1021 B.n409 B.n54 10.6151
R1022 B.n409 B.n408 10.6151
R1023 B.n408 B.n407 10.6151
R1024 B.n407 B.n56 10.6151
R1025 B.n403 B.n56 10.6151
R1026 B.n403 B.n402 10.6151
R1027 B.n402 B.n401 10.6151
R1028 B.n401 B.n58 10.6151
R1029 B.n397 B.n58 10.6151
R1030 B.n397 B.n396 10.6151
R1031 B.n396 B.n395 10.6151
R1032 B.n395 B.n60 10.6151
R1033 B.n391 B.n60 10.6151
R1034 B.n391 B.n390 10.6151
R1035 B.n390 B.n389 10.6151
R1036 B.n389 B.n62 10.6151
R1037 B.n385 B.n62 10.6151
R1038 B.n385 B.n384 10.6151
R1039 B.n384 B.n383 10.6151
R1040 B.n383 B.n64 10.6151
R1041 B.n379 B.n64 10.6151
R1042 B.n379 B.n378 10.6151
R1043 B.n378 B.n377 10.6151
R1044 B.n377 B.n66 10.6151
R1045 B.n373 B.n66 10.6151
R1046 B.n373 B.n372 10.6151
R1047 B.n372 B.n371 10.6151
R1048 B.n371 B.n68 10.6151
R1049 B.n367 B.n68 10.6151
R1050 B.n367 B.n366 10.6151
R1051 B.n366 B.n365 10.6151
R1052 B.n365 B.n70 10.6151
R1053 B.n361 B.n70 10.6151
R1054 B.n361 B.n360 10.6151
R1055 B.n360 B.n359 10.6151
R1056 B.n359 B.n72 10.6151
R1057 B.n355 B.n72 10.6151
R1058 B.n355 B.n354 10.6151
R1059 B.n354 B.n353 10.6151
R1060 B.n353 B.n74 10.6151
R1061 B.n349 B.n74 10.6151
R1062 B.n349 B.n348 10.6151
R1063 B.n348 B.n347 10.6151
R1064 B.n347 B.n76 10.6151
R1065 B.n343 B.n76 10.6151
R1066 B.n343 B.n342 10.6151
R1067 B.n342 B.n341 10.6151
R1068 B.n341 B.n78 10.6151
R1069 B.n337 B.n78 10.6151
R1070 B.n337 B.n336 10.6151
R1071 B.n336 B.n335 10.6151
R1072 B.n335 B.n80 10.6151
R1073 B.n331 B.n80 10.6151
R1074 B.n331 B.n330 10.6151
R1075 B.n330 B.n329 10.6151
R1076 B.n329 B.n82 10.6151
R1077 B.n325 B.n82 10.6151
R1078 B.n325 B.n324 10.6151
R1079 B.n324 B.n323 10.6151
R1080 B.n323 B.n84 10.6151
R1081 B.n319 B.n84 10.6151
R1082 B.n319 B.n318 10.6151
R1083 B.n318 B.n317 10.6151
R1084 B.n317 B.n86 10.6151
R1085 B.n313 B.n86 10.6151
R1086 B.n313 B.n312 10.6151
R1087 B.n312 B.n311 10.6151
R1088 B.n311 B.n88 10.6151
R1089 B.n307 B.n88 10.6151
R1090 B.n307 B.n306 10.6151
R1091 B.n306 B.n305 10.6151
R1092 B.n305 B.n90 10.6151
R1093 B.n301 B.n90 10.6151
R1094 B.n301 B.n300 10.6151
R1095 B.n300 B.n299 10.6151
R1096 B.n299 B.n92 10.6151
R1097 B.n295 B.n92 10.6151
R1098 B.n295 B.n294 10.6151
R1099 B.n294 B.n293 10.6151
R1100 B.n293 B.n94 10.6151
R1101 B.n289 B.n94 10.6151
R1102 B.n289 B.n288 10.6151
R1103 B.n288 B.n287 10.6151
R1104 B.n287 B.n96 10.6151
R1105 B.n283 B.n96 10.6151
R1106 B.n283 B.n282 10.6151
R1107 B.n145 B.n1 10.6151
R1108 B.n146 B.n145 10.6151
R1109 B.n147 B.n146 10.6151
R1110 B.n147 B.n142 10.6151
R1111 B.n151 B.n142 10.6151
R1112 B.n152 B.n151 10.6151
R1113 B.n153 B.n152 10.6151
R1114 B.n153 B.n140 10.6151
R1115 B.n157 B.n140 10.6151
R1116 B.n158 B.n157 10.6151
R1117 B.n159 B.n158 10.6151
R1118 B.n159 B.n138 10.6151
R1119 B.n163 B.n138 10.6151
R1120 B.n164 B.n163 10.6151
R1121 B.n165 B.n164 10.6151
R1122 B.n165 B.n136 10.6151
R1123 B.n169 B.n136 10.6151
R1124 B.n170 B.n169 10.6151
R1125 B.n171 B.n170 10.6151
R1126 B.n171 B.n134 10.6151
R1127 B.n175 B.n134 10.6151
R1128 B.n176 B.n175 10.6151
R1129 B.n177 B.n176 10.6151
R1130 B.n177 B.n132 10.6151
R1131 B.n181 B.n132 10.6151
R1132 B.n182 B.n181 10.6151
R1133 B.n183 B.n182 10.6151
R1134 B.n183 B.n130 10.6151
R1135 B.n187 B.n130 10.6151
R1136 B.n188 B.n187 10.6151
R1137 B.n189 B.n188 10.6151
R1138 B.n189 B.n128 10.6151
R1139 B.n193 B.n128 10.6151
R1140 B.n194 B.n193 10.6151
R1141 B.n195 B.n194 10.6151
R1142 B.n195 B.n126 10.6151
R1143 B.n199 B.n126 10.6151
R1144 B.n200 B.n199 10.6151
R1145 B.n201 B.n200 10.6151
R1146 B.n201 B.n124 10.6151
R1147 B.n205 B.n124 10.6151
R1148 B.n206 B.n205 10.6151
R1149 B.n207 B.n206 10.6151
R1150 B.n207 B.n122 10.6151
R1151 B.n212 B.n211 10.6151
R1152 B.n213 B.n212 10.6151
R1153 B.n213 B.n120 10.6151
R1154 B.n217 B.n120 10.6151
R1155 B.n218 B.n217 10.6151
R1156 B.n219 B.n218 10.6151
R1157 B.n219 B.n118 10.6151
R1158 B.n223 B.n118 10.6151
R1159 B.n224 B.n223 10.6151
R1160 B.n225 B.n224 10.6151
R1161 B.n225 B.n116 10.6151
R1162 B.n229 B.n116 10.6151
R1163 B.n230 B.n229 10.6151
R1164 B.n231 B.n230 10.6151
R1165 B.n231 B.n114 10.6151
R1166 B.n235 B.n114 10.6151
R1167 B.n236 B.n235 10.6151
R1168 B.n238 B.n110 10.6151
R1169 B.n242 B.n110 10.6151
R1170 B.n243 B.n242 10.6151
R1171 B.n244 B.n243 10.6151
R1172 B.n244 B.n108 10.6151
R1173 B.n248 B.n108 10.6151
R1174 B.n249 B.n248 10.6151
R1175 B.n253 B.n249 10.6151
R1176 B.n257 B.n106 10.6151
R1177 B.n258 B.n257 10.6151
R1178 B.n259 B.n258 10.6151
R1179 B.n259 B.n104 10.6151
R1180 B.n263 B.n104 10.6151
R1181 B.n264 B.n263 10.6151
R1182 B.n265 B.n264 10.6151
R1183 B.n265 B.n102 10.6151
R1184 B.n269 B.n102 10.6151
R1185 B.n270 B.n269 10.6151
R1186 B.n271 B.n270 10.6151
R1187 B.n271 B.n100 10.6151
R1188 B.n275 B.n100 10.6151
R1189 B.n276 B.n275 10.6151
R1190 B.n277 B.n276 10.6151
R1191 B.n277 B.n98 10.6151
R1192 B.n281 B.n98 10.6151
R1193 B.n557 B.n0 8.11757
R1194 B.n557 B.n1 8.11757
R1195 B.n461 B.n460 6.5566
R1196 B.n448 B.n42 6.5566
R1197 B.n238 B.n237 6.5566
R1198 B.n253 B.n252 6.5566
R1199 B.n462 B.n461 4.05904
R1200 B.n445 B.n42 4.05904
R1201 B.n237 B.n236 4.05904
R1202 B.n252 B.n106 4.05904
R1203 VP.n16 VP.n15 161.3
R1204 VP.n17 VP.n12 161.3
R1205 VP.n19 VP.n18 161.3
R1206 VP.n20 VP.n11 161.3
R1207 VP.n22 VP.n21 161.3
R1208 VP.n24 VP.n10 161.3
R1209 VP.n26 VP.n25 161.3
R1210 VP.n27 VP.n9 161.3
R1211 VP.n29 VP.n28 161.3
R1212 VP.n30 VP.n8 161.3
R1213 VP.n58 VP.n0 161.3
R1214 VP.n57 VP.n56 161.3
R1215 VP.n55 VP.n1 161.3
R1216 VP.n54 VP.n53 161.3
R1217 VP.n52 VP.n2 161.3
R1218 VP.n50 VP.n49 161.3
R1219 VP.n48 VP.n3 161.3
R1220 VP.n47 VP.n46 161.3
R1221 VP.n45 VP.n4 161.3
R1222 VP.n44 VP.n43 161.3
R1223 VP.n42 VP.n41 161.3
R1224 VP.n40 VP.n6 161.3
R1225 VP.n39 VP.n38 161.3
R1226 VP.n37 VP.n7 161.3
R1227 VP.n36 VP.n35 161.3
R1228 VP.n34 VP.n33 96.3991
R1229 VP.n60 VP.n59 96.3991
R1230 VP.n32 VP.n31 96.3991
R1231 VP.n14 VP.t0 75.2438
R1232 VP.n14 VP.n13 58.6104
R1233 VP.n39 VP.n7 43.4833
R1234 VP.n57 VP.n1 43.4833
R1235 VP.n29 VP.n9 43.4833
R1236 VP.n33 VP.n32 42.8633
R1237 VP.n34 VP.t2 42.5041
R1238 VP.n5 VP.t7 42.5041
R1239 VP.n51 VP.t4 42.5041
R1240 VP.n59 VP.t6 42.5041
R1241 VP.n31 VP.t3 42.5041
R1242 VP.n23 VP.t1 42.5041
R1243 VP.n13 VP.t5 42.5041
R1244 VP.n46 VP.n45 40.577
R1245 VP.n46 VP.n3 40.577
R1246 VP.n18 VP.n11 40.577
R1247 VP.n18 VP.n17 40.577
R1248 VP.n40 VP.n39 37.6707
R1249 VP.n53 VP.n1 37.6707
R1250 VP.n25 VP.n9 37.6707
R1251 VP.n35 VP.n7 24.5923
R1252 VP.n41 VP.n40 24.5923
R1253 VP.n45 VP.n44 24.5923
R1254 VP.n50 VP.n3 24.5923
R1255 VP.n53 VP.n52 24.5923
R1256 VP.n58 VP.n57 24.5923
R1257 VP.n30 VP.n29 24.5923
R1258 VP.n22 VP.n11 24.5923
R1259 VP.n25 VP.n24 24.5923
R1260 VP.n17 VP.n16 24.5923
R1261 VP.n35 VP.n34 14.5097
R1262 VP.n59 VP.n58 14.5097
R1263 VP.n31 VP.n30 14.5097
R1264 VP.n44 VP.n5 13.0342
R1265 VP.n51 VP.n50 13.0342
R1266 VP.n23 VP.n22 13.0342
R1267 VP.n16 VP.n13 13.0342
R1268 VP.n41 VP.n5 11.5587
R1269 VP.n52 VP.n51 11.5587
R1270 VP.n24 VP.n23 11.5587
R1271 VP.n15 VP.n14 9.48651
R1272 VP.n32 VP.n8 0.278335
R1273 VP.n36 VP.n33 0.278335
R1274 VP.n60 VP.n0 0.278335
R1275 VP.n15 VP.n12 0.189894
R1276 VP.n19 VP.n12 0.189894
R1277 VP.n20 VP.n19 0.189894
R1278 VP.n21 VP.n20 0.189894
R1279 VP.n21 VP.n10 0.189894
R1280 VP.n26 VP.n10 0.189894
R1281 VP.n27 VP.n26 0.189894
R1282 VP.n28 VP.n27 0.189894
R1283 VP.n28 VP.n8 0.189894
R1284 VP.n37 VP.n36 0.189894
R1285 VP.n38 VP.n37 0.189894
R1286 VP.n38 VP.n6 0.189894
R1287 VP.n42 VP.n6 0.189894
R1288 VP.n43 VP.n42 0.189894
R1289 VP.n43 VP.n4 0.189894
R1290 VP.n47 VP.n4 0.189894
R1291 VP.n48 VP.n47 0.189894
R1292 VP.n49 VP.n48 0.189894
R1293 VP.n49 VP.n2 0.189894
R1294 VP.n54 VP.n2 0.189894
R1295 VP.n55 VP.n54 0.189894
R1296 VP.n56 VP.n55 0.189894
R1297 VP.n56 VP.n0 0.189894
R1298 VP VP.n60 0.153485
R1299 VDD1 VDD1.n0 115.493
R1300 VDD1.n3 VDD1.n2 115.379
R1301 VDD1.n3 VDD1.n1 115.379
R1302 VDD1.n5 VDD1.n4 114.344
R1303 VDD1.n5 VDD1.n3 37.4578
R1304 VDD1.n4 VDD1.t6 8.37808
R1305 VDD1.n4 VDD1.t4 8.37808
R1306 VDD1.n0 VDD1.t7 8.37808
R1307 VDD1.n0 VDD1.t2 8.37808
R1308 VDD1.n2 VDD1.t3 8.37808
R1309 VDD1.n2 VDD1.t1 8.37808
R1310 VDD1.n1 VDD1.t5 8.37808
R1311 VDD1.n1 VDD1.t0 8.37808
R1312 VDD1 VDD1.n5 1.03283
C0 B w_n3500_n1744# 7.24378f
C1 B VTAIL 2.16038f
C2 VDD1 B 1.30938f
C3 VDD2 w_n3500_n1744# 1.69648f
C4 VN w_n3500_n1744# 6.86759f
C5 VDD2 VTAIL 5.11426f
C6 VDD1 VDD2 1.5664f
C7 VN VTAIL 3.81509f
C8 VN VDD1 0.155313f
C9 w_n3500_n1744# VP 7.31974f
C10 VP VTAIL 3.8292f
C11 VDD1 VP 3.34605f
C12 B VDD2 1.39297f
C13 VN B 1.05835f
C14 VN VDD2 3.02124f
C15 B VP 1.8157f
C16 VDD2 VP 0.481973f
C17 VN VP 5.67226f
C18 w_n3500_n1744# VTAIL 2.30529f
C19 VDD1 w_n3500_n1744# 1.59894f
C20 VDD1 VTAIL 5.06253f
C21 VDD2 VSUBS 1.366239f
C22 VDD1 VSUBS 1.954783f
C23 VTAIL VSUBS 0.597761f
C24 VN VSUBS 5.96969f
C25 VP VSUBS 2.649658f
C26 B VSUBS 3.652218f
C27 w_n3500_n1744# VSUBS 76.902f
C28 VDD1.t7 VSUBS 0.076204f
C29 VDD1.t2 VSUBS 0.076204f
C30 VDD1.n0 VSUBS 0.447107f
C31 VDD1.t5 VSUBS 0.076204f
C32 VDD1.t0 VSUBS 0.076204f
C33 VDD1.n1 VSUBS 0.446421f
C34 VDD1.t3 VSUBS 0.076204f
C35 VDD1.t1 VSUBS 0.076204f
C36 VDD1.n2 VSUBS 0.446421f
C37 VDD1.n3 VSUBS 2.87861f
C38 VDD1.t6 VSUBS 0.076204f
C39 VDD1.t4 VSUBS 0.076204f
C40 VDD1.n4 VSUBS 0.440898f
C41 VDD1.n5 VSUBS 2.33835f
C42 VP.n0 VSUBS 0.061851f
C43 VP.t6 VSUBS 1.02591f
C44 VP.n1 VSUBS 0.038434f
C45 VP.n2 VSUBS 0.046916f
C46 VP.t4 VSUBS 1.02591f
C47 VP.n3 VSUBS 0.092755f
C48 VP.n4 VSUBS 0.046916f
C49 VP.t7 VSUBS 1.02591f
C50 VP.n5 VSUBS 0.417059f
C51 VP.n6 VSUBS 0.046916f
C52 VP.n7 VSUBS 0.091107f
C53 VP.n8 VSUBS 0.061851f
C54 VP.t3 VSUBS 1.02591f
C55 VP.n9 VSUBS 0.038434f
C56 VP.n10 VSUBS 0.046916f
C57 VP.t1 VSUBS 1.02591f
C58 VP.n11 VSUBS 0.092755f
C59 VP.n12 VSUBS 0.046916f
C60 VP.t5 VSUBS 1.02591f
C61 VP.n13 VSUBS 0.538536f
C62 VP.t0 VSUBS 1.31657f
C63 VP.n14 VSUBS 0.519853f
C64 VP.n15 VSUBS 0.399396f
C65 VP.n16 VSUBS 0.066815f
C66 VP.n17 VSUBS 0.092755f
C67 VP.n18 VSUBS 0.037893f
C68 VP.n19 VSUBS 0.046916f
C69 VP.n20 VSUBS 0.046916f
C70 VP.n21 VSUBS 0.046916f
C71 VP.n22 VSUBS 0.066815f
C72 VP.n23 VSUBS 0.417059f
C73 VP.n24 VSUBS 0.064238f
C74 VP.n25 VSUBS 0.093861f
C75 VP.n26 VSUBS 0.046916f
C76 VP.n27 VSUBS 0.046916f
C77 VP.n28 VSUBS 0.046916f
C78 VP.n29 VSUBS 0.091107f
C79 VP.n30 VSUBS 0.069392f
C80 VP.n31 VSUBS 0.559222f
C81 VP.n32 VSUBS 2.05067f
C82 VP.n33 VSUBS 2.09013f
C83 VP.t2 VSUBS 1.02591f
C84 VP.n34 VSUBS 0.559222f
C85 VP.n35 VSUBS 0.069392f
C86 VP.n36 VSUBS 0.061851f
C87 VP.n37 VSUBS 0.046916f
C88 VP.n38 VSUBS 0.046916f
C89 VP.n39 VSUBS 0.038434f
C90 VP.n40 VSUBS 0.093861f
C91 VP.n41 VSUBS 0.064238f
C92 VP.n42 VSUBS 0.046916f
C93 VP.n43 VSUBS 0.046916f
C94 VP.n44 VSUBS 0.066815f
C95 VP.n45 VSUBS 0.092755f
C96 VP.n46 VSUBS 0.037893f
C97 VP.n47 VSUBS 0.046916f
C98 VP.n48 VSUBS 0.046916f
C99 VP.n49 VSUBS 0.046916f
C100 VP.n50 VSUBS 0.066815f
C101 VP.n51 VSUBS 0.417059f
C102 VP.n52 VSUBS 0.064238f
C103 VP.n53 VSUBS 0.093861f
C104 VP.n54 VSUBS 0.046916f
C105 VP.n55 VSUBS 0.046916f
C106 VP.n56 VSUBS 0.046916f
C107 VP.n57 VSUBS 0.091107f
C108 VP.n58 VSUBS 0.069392f
C109 VP.n59 VSUBS 0.559222f
C110 VP.n60 VSUBS 0.06569f
C111 B.n0 VSUBS 0.008108f
C112 B.n1 VSUBS 0.008108f
C113 B.n2 VSUBS 0.011991f
C114 B.n3 VSUBS 0.009189f
C115 B.n4 VSUBS 0.009189f
C116 B.n5 VSUBS 0.009189f
C117 B.n6 VSUBS 0.009189f
C118 B.n7 VSUBS 0.009189f
C119 B.n8 VSUBS 0.009189f
C120 B.n9 VSUBS 0.009189f
C121 B.n10 VSUBS 0.009189f
C122 B.n11 VSUBS 0.009189f
C123 B.n12 VSUBS 0.009189f
C124 B.n13 VSUBS 0.009189f
C125 B.n14 VSUBS 0.009189f
C126 B.n15 VSUBS 0.009189f
C127 B.n16 VSUBS 0.009189f
C128 B.n17 VSUBS 0.009189f
C129 B.n18 VSUBS 0.009189f
C130 B.n19 VSUBS 0.009189f
C131 B.n20 VSUBS 0.009189f
C132 B.n21 VSUBS 0.009189f
C133 B.n22 VSUBS 0.009189f
C134 B.n23 VSUBS 0.009189f
C135 B.n24 VSUBS 0.020324f
C136 B.n25 VSUBS 0.009189f
C137 B.n26 VSUBS 0.009189f
C138 B.n27 VSUBS 0.009189f
C139 B.n28 VSUBS 0.009189f
C140 B.n29 VSUBS 0.009189f
C141 B.n30 VSUBS 0.009189f
C142 B.n31 VSUBS 0.009189f
C143 B.n32 VSUBS 0.009189f
C144 B.n33 VSUBS 0.009189f
C145 B.t10 VSUBS 0.073517f
C146 B.t11 VSUBS 0.096701f
C147 B.t9 VSUBS 0.536408f
C148 B.n34 VSUBS 0.171199f
C149 B.n35 VSUBS 0.146524f
C150 B.n36 VSUBS 0.009189f
C151 B.n37 VSUBS 0.009189f
C152 B.n38 VSUBS 0.009189f
C153 B.n39 VSUBS 0.009189f
C154 B.t1 VSUBS 0.073518f
C155 B.t2 VSUBS 0.096702f
C156 B.t0 VSUBS 0.536408f
C157 B.n40 VSUBS 0.171198f
C158 B.n41 VSUBS 0.146523f
C159 B.n42 VSUBS 0.02129f
C160 B.n43 VSUBS 0.009189f
C161 B.n44 VSUBS 0.009189f
C162 B.n45 VSUBS 0.009189f
C163 B.n46 VSUBS 0.009189f
C164 B.n47 VSUBS 0.009189f
C165 B.n48 VSUBS 0.009189f
C166 B.n49 VSUBS 0.009189f
C167 B.n50 VSUBS 0.009189f
C168 B.n51 VSUBS 0.021027f
C169 B.n52 VSUBS 0.009189f
C170 B.n53 VSUBS 0.009189f
C171 B.n54 VSUBS 0.009189f
C172 B.n55 VSUBS 0.009189f
C173 B.n56 VSUBS 0.009189f
C174 B.n57 VSUBS 0.009189f
C175 B.n58 VSUBS 0.009189f
C176 B.n59 VSUBS 0.009189f
C177 B.n60 VSUBS 0.009189f
C178 B.n61 VSUBS 0.009189f
C179 B.n62 VSUBS 0.009189f
C180 B.n63 VSUBS 0.009189f
C181 B.n64 VSUBS 0.009189f
C182 B.n65 VSUBS 0.009189f
C183 B.n66 VSUBS 0.009189f
C184 B.n67 VSUBS 0.009189f
C185 B.n68 VSUBS 0.009189f
C186 B.n69 VSUBS 0.009189f
C187 B.n70 VSUBS 0.009189f
C188 B.n71 VSUBS 0.009189f
C189 B.n72 VSUBS 0.009189f
C190 B.n73 VSUBS 0.009189f
C191 B.n74 VSUBS 0.009189f
C192 B.n75 VSUBS 0.009189f
C193 B.n76 VSUBS 0.009189f
C194 B.n77 VSUBS 0.009189f
C195 B.n78 VSUBS 0.009189f
C196 B.n79 VSUBS 0.009189f
C197 B.n80 VSUBS 0.009189f
C198 B.n81 VSUBS 0.009189f
C199 B.n82 VSUBS 0.009189f
C200 B.n83 VSUBS 0.009189f
C201 B.n84 VSUBS 0.009189f
C202 B.n85 VSUBS 0.009189f
C203 B.n86 VSUBS 0.009189f
C204 B.n87 VSUBS 0.009189f
C205 B.n88 VSUBS 0.009189f
C206 B.n89 VSUBS 0.009189f
C207 B.n90 VSUBS 0.009189f
C208 B.n91 VSUBS 0.009189f
C209 B.n92 VSUBS 0.009189f
C210 B.n93 VSUBS 0.009189f
C211 B.n94 VSUBS 0.009189f
C212 B.n95 VSUBS 0.009189f
C213 B.n96 VSUBS 0.009189f
C214 B.n97 VSUBS 0.020324f
C215 B.n98 VSUBS 0.009189f
C216 B.n99 VSUBS 0.009189f
C217 B.n100 VSUBS 0.009189f
C218 B.n101 VSUBS 0.009189f
C219 B.n102 VSUBS 0.009189f
C220 B.n103 VSUBS 0.009189f
C221 B.n104 VSUBS 0.009189f
C222 B.n105 VSUBS 0.009189f
C223 B.n106 VSUBS 0.006351f
C224 B.n107 VSUBS 0.009189f
C225 B.n108 VSUBS 0.009189f
C226 B.n109 VSUBS 0.009189f
C227 B.n110 VSUBS 0.009189f
C228 B.n111 VSUBS 0.009189f
C229 B.t5 VSUBS 0.073517f
C230 B.t4 VSUBS 0.096701f
C231 B.t3 VSUBS 0.536408f
C232 B.n112 VSUBS 0.171199f
C233 B.n113 VSUBS 0.146524f
C234 B.n114 VSUBS 0.009189f
C235 B.n115 VSUBS 0.009189f
C236 B.n116 VSUBS 0.009189f
C237 B.n117 VSUBS 0.009189f
C238 B.n118 VSUBS 0.009189f
C239 B.n119 VSUBS 0.009189f
C240 B.n120 VSUBS 0.009189f
C241 B.n121 VSUBS 0.009189f
C242 B.n122 VSUBS 0.020324f
C243 B.n123 VSUBS 0.009189f
C244 B.n124 VSUBS 0.009189f
C245 B.n125 VSUBS 0.009189f
C246 B.n126 VSUBS 0.009189f
C247 B.n127 VSUBS 0.009189f
C248 B.n128 VSUBS 0.009189f
C249 B.n129 VSUBS 0.009189f
C250 B.n130 VSUBS 0.009189f
C251 B.n131 VSUBS 0.009189f
C252 B.n132 VSUBS 0.009189f
C253 B.n133 VSUBS 0.009189f
C254 B.n134 VSUBS 0.009189f
C255 B.n135 VSUBS 0.009189f
C256 B.n136 VSUBS 0.009189f
C257 B.n137 VSUBS 0.009189f
C258 B.n138 VSUBS 0.009189f
C259 B.n139 VSUBS 0.009189f
C260 B.n140 VSUBS 0.009189f
C261 B.n141 VSUBS 0.009189f
C262 B.n142 VSUBS 0.009189f
C263 B.n143 VSUBS 0.009189f
C264 B.n144 VSUBS 0.009189f
C265 B.n145 VSUBS 0.009189f
C266 B.n146 VSUBS 0.009189f
C267 B.n147 VSUBS 0.009189f
C268 B.n148 VSUBS 0.009189f
C269 B.n149 VSUBS 0.009189f
C270 B.n150 VSUBS 0.009189f
C271 B.n151 VSUBS 0.009189f
C272 B.n152 VSUBS 0.009189f
C273 B.n153 VSUBS 0.009189f
C274 B.n154 VSUBS 0.009189f
C275 B.n155 VSUBS 0.009189f
C276 B.n156 VSUBS 0.009189f
C277 B.n157 VSUBS 0.009189f
C278 B.n158 VSUBS 0.009189f
C279 B.n159 VSUBS 0.009189f
C280 B.n160 VSUBS 0.009189f
C281 B.n161 VSUBS 0.009189f
C282 B.n162 VSUBS 0.009189f
C283 B.n163 VSUBS 0.009189f
C284 B.n164 VSUBS 0.009189f
C285 B.n165 VSUBS 0.009189f
C286 B.n166 VSUBS 0.009189f
C287 B.n167 VSUBS 0.009189f
C288 B.n168 VSUBS 0.009189f
C289 B.n169 VSUBS 0.009189f
C290 B.n170 VSUBS 0.009189f
C291 B.n171 VSUBS 0.009189f
C292 B.n172 VSUBS 0.009189f
C293 B.n173 VSUBS 0.009189f
C294 B.n174 VSUBS 0.009189f
C295 B.n175 VSUBS 0.009189f
C296 B.n176 VSUBS 0.009189f
C297 B.n177 VSUBS 0.009189f
C298 B.n178 VSUBS 0.009189f
C299 B.n179 VSUBS 0.009189f
C300 B.n180 VSUBS 0.009189f
C301 B.n181 VSUBS 0.009189f
C302 B.n182 VSUBS 0.009189f
C303 B.n183 VSUBS 0.009189f
C304 B.n184 VSUBS 0.009189f
C305 B.n185 VSUBS 0.009189f
C306 B.n186 VSUBS 0.009189f
C307 B.n187 VSUBS 0.009189f
C308 B.n188 VSUBS 0.009189f
C309 B.n189 VSUBS 0.009189f
C310 B.n190 VSUBS 0.009189f
C311 B.n191 VSUBS 0.009189f
C312 B.n192 VSUBS 0.009189f
C313 B.n193 VSUBS 0.009189f
C314 B.n194 VSUBS 0.009189f
C315 B.n195 VSUBS 0.009189f
C316 B.n196 VSUBS 0.009189f
C317 B.n197 VSUBS 0.009189f
C318 B.n198 VSUBS 0.009189f
C319 B.n199 VSUBS 0.009189f
C320 B.n200 VSUBS 0.009189f
C321 B.n201 VSUBS 0.009189f
C322 B.n202 VSUBS 0.009189f
C323 B.n203 VSUBS 0.009189f
C324 B.n204 VSUBS 0.009189f
C325 B.n205 VSUBS 0.009189f
C326 B.n206 VSUBS 0.009189f
C327 B.n207 VSUBS 0.009189f
C328 B.n208 VSUBS 0.009189f
C329 B.n209 VSUBS 0.020324f
C330 B.n210 VSUBS 0.021027f
C331 B.n211 VSUBS 0.021027f
C332 B.n212 VSUBS 0.009189f
C333 B.n213 VSUBS 0.009189f
C334 B.n214 VSUBS 0.009189f
C335 B.n215 VSUBS 0.009189f
C336 B.n216 VSUBS 0.009189f
C337 B.n217 VSUBS 0.009189f
C338 B.n218 VSUBS 0.009189f
C339 B.n219 VSUBS 0.009189f
C340 B.n220 VSUBS 0.009189f
C341 B.n221 VSUBS 0.009189f
C342 B.n222 VSUBS 0.009189f
C343 B.n223 VSUBS 0.009189f
C344 B.n224 VSUBS 0.009189f
C345 B.n225 VSUBS 0.009189f
C346 B.n226 VSUBS 0.009189f
C347 B.n227 VSUBS 0.009189f
C348 B.n228 VSUBS 0.009189f
C349 B.n229 VSUBS 0.009189f
C350 B.n230 VSUBS 0.009189f
C351 B.n231 VSUBS 0.009189f
C352 B.n232 VSUBS 0.009189f
C353 B.n233 VSUBS 0.009189f
C354 B.n234 VSUBS 0.009189f
C355 B.n235 VSUBS 0.009189f
C356 B.n236 VSUBS 0.006351f
C357 B.n237 VSUBS 0.02129f
C358 B.n238 VSUBS 0.007432f
C359 B.n239 VSUBS 0.009189f
C360 B.n240 VSUBS 0.009189f
C361 B.n241 VSUBS 0.009189f
C362 B.n242 VSUBS 0.009189f
C363 B.n243 VSUBS 0.009189f
C364 B.n244 VSUBS 0.009189f
C365 B.n245 VSUBS 0.009189f
C366 B.n246 VSUBS 0.009189f
C367 B.n247 VSUBS 0.009189f
C368 B.n248 VSUBS 0.009189f
C369 B.n249 VSUBS 0.009189f
C370 B.t8 VSUBS 0.073518f
C371 B.t7 VSUBS 0.096702f
C372 B.t6 VSUBS 0.536408f
C373 B.n250 VSUBS 0.171198f
C374 B.n251 VSUBS 0.146523f
C375 B.n252 VSUBS 0.02129f
C376 B.n253 VSUBS 0.007432f
C377 B.n254 VSUBS 0.009189f
C378 B.n255 VSUBS 0.009189f
C379 B.n256 VSUBS 0.009189f
C380 B.n257 VSUBS 0.009189f
C381 B.n258 VSUBS 0.009189f
C382 B.n259 VSUBS 0.009189f
C383 B.n260 VSUBS 0.009189f
C384 B.n261 VSUBS 0.009189f
C385 B.n262 VSUBS 0.009189f
C386 B.n263 VSUBS 0.009189f
C387 B.n264 VSUBS 0.009189f
C388 B.n265 VSUBS 0.009189f
C389 B.n266 VSUBS 0.009189f
C390 B.n267 VSUBS 0.009189f
C391 B.n268 VSUBS 0.009189f
C392 B.n269 VSUBS 0.009189f
C393 B.n270 VSUBS 0.009189f
C394 B.n271 VSUBS 0.009189f
C395 B.n272 VSUBS 0.009189f
C396 B.n273 VSUBS 0.009189f
C397 B.n274 VSUBS 0.009189f
C398 B.n275 VSUBS 0.009189f
C399 B.n276 VSUBS 0.009189f
C400 B.n277 VSUBS 0.009189f
C401 B.n278 VSUBS 0.009189f
C402 B.n279 VSUBS 0.009189f
C403 B.n280 VSUBS 0.021027f
C404 B.n281 VSUBS 0.019874f
C405 B.n282 VSUBS 0.021477f
C406 B.n283 VSUBS 0.009189f
C407 B.n284 VSUBS 0.009189f
C408 B.n285 VSUBS 0.009189f
C409 B.n286 VSUBS 0.009189f
C410 B.n287 VSUBS 0.009189f
C411 B.n288 VSUBS 0.009189f
C412 B.n289 VSUBS 0.009189f
C413 B.n290 VSUBS 0.009189f
C414 B.n291 VSUBS 0.009189f
C415 B.n292 VSUBS 0.009189f
C416 B.n293 VSUBS 0.009189f
C417 B.n294 VSUBS 0.009189f
C418 B.n295 VSUBS 0.009189f
C419 B.n296 VSUBS 0.009189f
C420 B.n297 VSUBS 0.009189f
C421 B.n298 VSUBS 0.009189f
C422 B.n299 VSUBS 0.009189f
C423 B.n300 VSUBS 0.009189f
C424 B.n301 VSUBS 0.009189f
C425 B.n302 VSUBS 0.009189f
C426 B.n303 VSUBS 0.009189f
C427 B.n304 VSUBS 0.009189f
C428 B.n305 VSUBS 0.009189f
C429 B.n306 VSUBS 0.009189f
C430 B.n307 VSUBS 0.009189f
C431 B.n308 VSUBS 0.009189f
C432 B.n309 VSUBS 0.009189f
C433 B.n310 VSUBS 0.009189f
C434 B.n311 VSUBS 0.009189f
C435 B.n312 VSUBS 0.009189f
C436 B.n313 VSUBS 0.009189f
C437 B.n314 VSUBS 0.009189f
C438 B.n315 VSUBS 0.009189f
C439 B.n316 VSUBS 0.009189f
C440 B.n317 VSUBS 0.009189f
C441 B.n318 VSUBS 0.009189f
C442 B.n319 VSUBS 0.009189f
C443 B.n320 VSUBS 0.009189f
C444 B.n321 VSUBS 0.009189f
C445 B.n322 VSUBS 0.009189f
C446 B.n323 VSUBS 0.009189f
C447 B.n324 VSUBS 0.009189f
C448 B.n325 VSUBS 0.009189f
C449 B.n326 VSUBS 0.009189f
C450 B.n327 VSUBS 0.009189f
C451 B.n328 VSUBS 0.009189f
C452 B.n329 VSUBS 0.009189f
C453 B.n330 VSUBS 0.009189f
C454 B.n331 VSUBS 0.009189f
C455 B.n332 VSUBS 0.009189f
C456 B.n333 VSUBS 0.009189f
C457 B.n334 VSUBS 0.009189f
C458 B.n335 VSUBS 0.009189f
C459 B.n336 VSUBS 0.009189f
C460 B.n337 VSUBS 0.009189f
C461 B.n338 VSUBS 0.009189f
C462 B.n339 VSUBS 0.009189f
C463 B.n340 VSUBS 0.009189f
C464 B.n341 VSUBS 0.009189f
C465 B.n342 VSUBS 0.009189f
C466 B.n343 VSUBS 0.009189f
C467 B.n344 VSUBS 0.009189f
C468 B.n345 VSUBS 0.009189f
C469 B.n346 VSUBS 0.009189f
C470 B.n347 VSUBS 0.009189f
C471 B.n348 VSUBS 0.009189f
C472 B.n349 VSUBS 0.009189f
C473 B.n350 VSUBS 0.009189f
C474 B.n351 VSUBS 0.009189f
C475 B.n352 VSUBS 0.009189f
C476 B.n353 VSUBS 0.009189f
C477 B.n354 VSUBS 0.009189f
C478 B.n355 VSUBS 0.009189f
C479 B.n356 VSUBS 0.009189f
C480 B.n357 VSUBS 0.009189f
C481 B.n358 VSUBS 0.009189f
C482 B.n359 VSUBS 0.009189f
C483 B.n360 VSUBS 0.009189f
C484 B.n361 VSUBS 0.009189f
C485 B.n362 VSUBS 0.009189f
C486 B.n363 VSUBS 0.009189f
C487 B.n364 VSUBS 0.009189f
C488 B.n365 VSUBS 0.009189f
C489 B.n366 VSUBS 0.009189f
C490 B.n367 VSUBS 0.009189f
C491 B.n368 VSUBS 0.009189f
C492 B.n369 VSUBS 0.009189f
C493 B.n370 VSUBS 0.009189f
C494 B.n371 VSUBS 0.009189f
C495 B.n372 VSUBS 0.009189f
C496 B.n373 VSUBS 0.009189f
C497 B.n374 VSUBS 0.009189f
C498 B.n375 VSUBS 0.009189f
C499 B.n376 VSUBS 0.009189f
C500 B.n377 VSUBS 0.009189f
C501 B.n378 VSUBS 0.009189f
C502 B.n379 VSUBS 0.009189f
C503 B.n380 VSUBS 0.009189f
C504 B.n381 VSUBS 0.009189f
C505 B.n382 VSUBS 0.009189f
C506 B.n383 VSUBS 0.009189f
C507 B.n384 VSUBS 0.009189f
C508 B.n385 VSUBS 0.009189f
C509 B.n386 VSUBS 0.009189f
C510 B.n387 VSUBS 0.009189f
C511 B.n388 VSUBS 0.009189f
C512 B.n389 VSUBS 0.009189f
C513 B.n390 VSUBS 0.009189f
C514 B.n391 VSUBS 0.009189f
C515 B.n392 VSUBS 0.009189f
C516 B.n393 VSUBS 0.009189f
C517 B.n394 VSUBS 0.009189f
C518 B.n395 VSUBS 0.009189f
C519 B.n396 VSUBS 0.009189f
C520 B.n397 VSUBS 0.009189f
C521 B.n398 VSUBS 0.009189f
C522 B.n399 VSUBS 0.009189f
C523 B.n400 VSUBS 0.009189f
C524 B.n401 VSUBS 0.009189f
C525 B.n402 VSUBS 0.009189f
C526 B.n403 VSUBS 0.009189f
C527 B.n404 VSUBS 0.009189f
C528 B.n405 VSUBS 0.009189f
C529 B.n406 VSUBS 0.009189f
C530 B.n407 VSUBS 0.009189f
C531 B.n408 VSUBS 0.009189f
C532 B.n409 VSUBS 0.009189f
C533 B.n410 VSUBS 0.009189f
C534 B.n411 VSUBS 0.009189f
C535 B.n412 VSUBS 0.009189f
C536 B.n413 VSUBS 0.009189f
C537 B.n414 VSUBS 0.009189f
C538 B.n415 VSUBS 0.009189f
C539 B.n416 VSUBS 0.009189f
C540 B.n417 VSUBS 0.009189f
C541 B.n418 VSUBS 0.020324f
C542 B.n419 VSUBS 0.020324f
C543 B.n420 VSUBS 0.021027f
C544 B.n421 VSUBS 0.009189f
C545 B.n422 VSUBS 0.009189f
C546 B.n423 VSUBS 0.009189f
C547 B.n424 VSUBS 0.009189f
C548 B.n425 VSUBS 0.009189f
C549 B.n426 VSUBS 0.009189f
C550 B.n427 VSUBS 0.009189f
C551 B.n428 VSUBS 0.009189f
C552 B.n429 VSUBS 0.009189f
C553 B.n430 VSUBS 0.009189f
C554 B.n431 VSUBS 0.009189f
C555 B.n432 VSUBS 0.009189f
C556 B.n433 VSUBS 0.009189f
C557 B.n434 VSUBS 0.009189f
C558 B.n435 VSUBS 0.009189f
C559 B.n436 VSUBS 0.009189f
C560 B.n437 VSUBS 0.009189f
C561 B.n438 VSUBS 0.009189f
C562 B.n439 VSUBS 0.009189f
C563 B.n440 VSUBS 0.009189f
C564 B.n441 VSUBS 0.009189f
C565 B.n442 VSUBS 0.009189f
C566 B.n443 VSUBS 0.009189f
C567 B.n444 VSUBS 0.009189f
C568 B.n445 VSUBS 0.006351f
C569 B.n446 VSUBS 0.009189f
C570 B.n447 VSUBS 0.009189f
C571 B.n448 VSUBS 0.007432f
C572 B.n449 VSUBS 0.009189f
C573 B.n450 VSUBS 0.009189f
C574 B.n451 VSUBS 0.009189f
C575 B.n452 VSUBS 0.009189f
C576 B.n453 VSUBS 0.009189f
C577 B.n454 VSUBS 0.009189f
C578 B.n455 VSUBS 0.009189f
C579 B.n456 VSUBS 0.009189f
C580 B.n457 VSUBS 0.009189f
C581 B.n458 VSUBS 0.009189f
C582 B.n459 VSUBS 0.009189f
C583 B.n460 VSUBS 0.007432f
C584 B.n461 VSUBS 0.02129f
C585 B.n462 VSUBS 0.006351f
C586 B.n463 VSUBS 0.009189f
C587 B.n464 VSUBS 0.009189f
C588 B.n465 VSUBS 0.009189f
C589 B.n466 VSUBS 0.009189f
C590 B.n467 VSUBS 0.009189f
C591 B.n468 VSUBS 0.009189f
C592 B.n469 VSUBS 0.009189f
C593 B.n470 VSUBS 0.009189f
C594 B.n471 VSUBS 0.009189f
C595 B.n472 VSUBS 0.009189f
C596 B.n473 VSUBS 0.009189f
C597 B.n474 VSUBS 0.009189f
C598 B.n475 VSUBS 0.009189f
C599 B.n476 VSUBS 0.009189f
C600 B.n477 VSUBS 0.009189f
C601 B.n478 VSUBS 0.009189f
C602 B.n479 VSUBS 0.009189f
C603 B.n480 VSUBS 0.009189f
C604 B.n481 VSUBS 0.009189f
C605 B.n482 VSUBS 0.009189f
C606 B.n483 VSUBS 0.009189f
C607 B.n484 VSUBS 0.009189f
C608 B.n485 VSUBS 0.009189f
C609 B.n486 VSUBS 0.009189f
C610 B.n487 VSUBS 0.021027f
C611 B.n488 VSUBS 0.021027f
C612 B.n489 VSUBS 0.020324f
C613 B.n490 VSUBS 0.009189f
C614 B.n491 VSUBS 0.009189f
C615 B.n492 VSUBS 0.009189f
C616 B.n493 VSUBS 0.009189f
C617 B.n494 VSUBS 0.009189f
C618 B.n495 VSUBS 0.009189f
C619 B.n496 VSUBS 0.009189f
C620 B.n497 VSUBS 0.009189f
C621 B.n498 VSUBS 0.009189f
C622 B.n499 VSUBS 0.009189f
C623 B.n500 VSUBS 0.009189f
C624 B.n501 VSUBS 0.009189f
C625 B.n502 VSUBS 0.009189f
C626 B.n503 VSUBS 0.009189f
C627 B.n504 VSUBS 0.009189f
C628 B.n505 VSUBS 0.009189f
C629 B.n506 VSUBS 0.009189f
C630 B.n507 VSUBS 0.009189f
C631 B.n508 VSUBS 0.009189f
C632 B.n509 VSUBS 0.009189f
C633 B.n510 VSUBS 0.009189f
C634 B.n511 VSUBS 0.009189f
C635 B.n512 VSUBS 0.009189f
C636 B.n513 VSUBS 0.009189f
C637 B.n514 VSUBS 0.009189f
C638 B.n515 VSUBS 0.009189f
C639 B.n516 VSUBS 0.009189f
C640 B.n517 VSUBS 0.009189f
C641 B.n518 VSUBS 0.009189f
C642 B.n519 VSUBS 0.009189f
C643 B.n520 VSUBS 0.009189f
C644 B.n521 VSUBS 0.009189f
C645 B.n522 VSUBS 0.009189f
C646 B.n523 VSUBS 0.009189f
C647 B.n524 VSUBS 0.009189f
C648 B.n525 VSUBS 0.009189f
C649 B.n526 VSUBS 0.009189f
C650 B.n527 VSUBS 0.009189f
C651 B.n528 VSUBS 0.009189f
C652 B.n529 VSUBS 0.009189f
C653 B.n530 VSUBS 0.009189f
C654 B.n531 VSUBS 0.009189f
C655 B.n532 VSUBS 0.009189f
C656 B.n533 VSUBS 0.009189f
C657 B.n534 VSUBS 0.009189f
C658 B.n535 VSUBS 0.009189f
C659 B.n536 VSUBS 0.009189f
C660 B.n537 VSUBS 0.009189f
C661 B.n538 VSUBS 0.009189f
C662 B.n539 VSUBS 0.009189f
C663 B.n540 VSUBS 0.009189f
C664 B.n541 VSUBS 0.009189f
C665 B.n542 VSUBS 0.009189f
C666 B.n543 VSUBS 0.009189f
C667 B.n544 VSUBS 0.009189f
C668 B.n545 VSUBS 0.009189f
C669 B.n546 VSUBS 0.009189f
C670 B.n547 VSUBS 0.009189f
C671 B.n548 VSUBS 0.009189f
C672 B.n549 VSUBS 0.009189f
C673 B.n550 VSUBS 0.009189f
C674 B.n551 VSUBS 0.009189f
C675 B.n552 VSUBS 0.009189f
C676 B.n553 VSUBS 0.009189f
C677 B.n554 VSUBS 0.009189f
C678 B.n555 VSUBS 0.011991f
C679 B.n556 VSUBS 0.012774f
C680 B.n557 VSUBS 0.025402f
C681 VTAIL.t11 VSUBS 0.097705f
C682 VTAIL.t7 VSUBS 0.097705f
C683 VTAIL.n0 VSUBS 0.490259f
C684 VTAIL.n1 VSUBS 0.707115f
C685 VTAIL.n2 VSUBS 0.0338f
C686 VTAIL.n3 VSUBS 0.031866f
C687 VTAIL.n4 VSUBS 0.017124f
C688 VTAIL.n5 VSUBS 0.040474f
C689 VTAIL.n6 VSUBS 0.018131f
C690 VTAIL.n7 VSUBS 0.122345f
C691 VTAIL.t8 VSUBS 0.088965f
C692 VTAIL.n8 VSUBS 0.030355f
C693 VTAIL.n9 VSUBS 0.025458f
C694 VTAIL.n10 VSUBS 0.017124f
C695 VTAIL.n11 VSUBS 0.420918f
C696 VTAIL.n12 VSUBS 0.031866f
C697 VTAIL.n13 VSUBS 0.017124f
C698 VTAIL.n14 VSUBS 0.018131f
C699 VTAIL.n15 VSUBS 0.040474f
C700 VTAIL.n16 VSUBS 0.093848f
C701 VTAIL.n17 VSUBS 0.018131f
C702 VTAIL.n18 VSUBS 0.017124f
C703 VTAIL.n19 VSUBS 0.075399f
C704 VTAIL.n20 VSUBS 0.047065f
C705 VTAIL.n21 VSUBS 0.300391f
C706 VTAIL.n22 VSUBS 0.0338f
C707 VTAIL.n23 VSUBS 0.031866f
C708 VTAIL.n24 VSUBS 0.017124f
C709 VTAIL.n25 VSUBS 0.040474f
C710 VTAIL.n26 VSUBS 0.018131f
C711 VTAIL.n27 VSUBS 0.122345f
C712 VTAIL.t15 VSUBS 0.088965f
C713 VTAIL.n28 VSUBS 0.030355f
C714 VTAIL.n29 VSUBS 0.025458f
C715 VTAIL.n30 VSUBS 0.017124f
C716 VTAIL.n31 VSUBS 0.420918f
C717 VTAIL.n32 VSUBS 0.031866f
C718 VTAIL.n33 VSUBS 0.017124f
C719 VTAIL.n34 VSUBS 0.018131f
C720 VTAIL.n35 VSUBS 0.040474f
C721 VTAIL.n36 VSUBS 0.093848f
C722 VTAIL.n37 VSUBS 0.018131f
C723 VTAIL.n38 VSUBS 0.017124f
C724 VTAIL.n39 VSUBS 0.075399f
C725 VTAIL.n40 VSUBS 0.047065f
C726 VTAIL.n41 VSUBS 0.300391f
C727 VTAIL.t6 VSUBS 0.097705f
C728 VTAIL.t0 VSUBS 0.097705f
C729 VTAIL.n42 VSUBS 0.490259f
C730 VTAIL.n43 VSUBS 0.925089f
C731 VTAIL.n44 VSUBS 0.0338f
C732 VTAIL.n45 VSUBS 0.031866f
C733 VTAIL.n46 VSUBS 0.017124f
C734 VTAIL.n47 VSUBS 0.040474f
C735 VTAIL.n48 VSUBS 0.018131f
C736 VTAIL.n49 VSUBS 0.122345f
C737 VTAIL.t2 VSUBS 0.088965f
C738 VTAIL.n50 VSUBS 0.030355f
C739 VTAIL.n51 VSUBS 0.025458f
C740 VTAIL.n52 VSUBS 0.017124f
C741 VTAIL.n53 VSUBS 0.420918f
C742 VTAIL.n54 VSUBS 0.031866f
C743 VTAIL.n55 VSUBS 0.017124f
C744 VTAIL.n56 VSUBS 0.018131f
C745 VTAIL.n57 VSUBS 0.040474f
C746 VTAIL.n58 VSUBS 0.093848f
C747 VTAIL.n59 VSUBS 0.018131f
C748 VTAIL.n60 VSUBS 0.017124f
C749 VTAIL.n61 VSUBS 0.075399f
C750 VTAIL.n62 VSUBS 0.047065f
C751 VTAIL.n63 VSUBS 1.25241f
C752 VTAIL.n64 VSUBS 0.0338f
C753 VTAIL.n65 VSUBS 0.031866f
C754 VTAIL.n66 VSUBS 0.017124f
C755 VTAIL.n67 VSUBS 0.040474f
C756 VTAIL.n68 VSUBS 0.018131f
C757 VTAIL.n69 VSUBS 0.122345f
C758 VTAIL.t13 VSUBS 0.088965f
C759 VTAIL.n70 VSUBS 0.030355f
C760 VTAIL.n71 VSUBS 0.025458f
C761 VTAIL.n72 VSUBS 0.017124f
C762 VTAIL.n73 VSUBS 0.420918f
C763 VTAIL.n74 VSUBS 0.031866f
C764 VTAIL.n75 VSUBS 0.017124f
C765 VTAIL.n76 VSUBS 0.018131f
C766 VTAIL.n77 VSUBS 0.040474f
C767 VTAIL.n78 VSUBS 0.093848f
C768 VTAIL.n79 VSUBS 0.018131f
C769 VTAIL.n80 VSUBS 0.017124f
C770 VTAIL.n81 VSUBS 0.075399f
C771 VTAIL.n82 VSUBS 0.047065f
C772 VTAIL.n83 VSUBS 1.25241f
C773 VTAIL.t10 VSUBS 0.097705f
C774 VTAIL.t14 VSUBS 0.097705f
C775 VTAIL.n84 VSUBS 0.490263f
C776 VTAIL.n85 VSUBS 0.925086f
C777 VTAIL.n86 VSUBS 0.0338f
C778 VTAIL.n87 VSUBS 0.031866f
C779 VTAIL.n88 VSUBS 0.017124f
C780 VTAIL.n89 VSUBS 0.040474f
C781 VTAIL.n90 VSUBS 0.018131f
C782 VTAIL.n91 VSUBS 0.122345f
C783 VTAIL.t12 VSUBS 0.088965f
C784 VTAIL.n92 VSUBS 0.030355f
C785 VTAIL.n93 VSUBS 0.025458f
C786 VTAIL.n94 VSUBS 0.017124f
C787 VTAIL.n95 VSUBS 0.420918f
C788 VTAIL.n96 VSUBS 0.031866f
C789 VTAIL.n97 VSUBS 0.017124f
C790 VTAIL.n98 VSUBS 0.018131f
C791 VTAIL.n99 VSUBS 0.040474f
C792 VTAIL.n100 VSUBS 0.093848f
C793 VTAIL.n101 VSUBS 0.018131f
C794 VTAIL.n102 VSUBS 0.017124f
C795 VTAIL.n103 VSUBS 0.075399f
C796 VTAIL.n104 VSUBS 0.047065f
C797 VTAIL.n105 VSUBS 0.300391f
C798 VTAIL.n106 VSUBS 0.0338f
C799 VTAIL.n107 VSUBS 0.031866f
C800 VTAIL.n108 VSUBS 0.017124f
C801 VTAIL.n109 VSUBS 0.040474f
C802 VTAIL.n110 VSUBS 0.018131f
C803 VTAIL.n111 VSUBS 0.122345f
C804 VTAIL.t3 VSUBS 0.088965f
C805 VTAIL.n112 VSUBS 0.030355f
C806 VTAIL.n113 VSUBS 0.025458f
C807 VTAIL.n114 VSUBS 0.017124f
C808 VTAIL.n115 VSUBS 0.420918f
C809 VTAIL.n116 VSUBS 0.031866f
C810 VTAIL.n117 VSUBS 0.017124f
C811 VTAIL.n118 VSUBS 0.018131f
C812 VTAIL.n119 VSUBS 0.040474f
C813 VTAIL.n120 VSUBS 0.093848f
C814 VTAIL.n121 VSUBS 0.018131f
C815 VTAIL.n122 VSUBS 0.017124f
C816 VTAIL.n123 VSUBS 0.075399f
C817 VTAIL.n124 VSUBS 0.047065f
C818 VTAIL.n125 VSUBS 0.300391f
C819 VTAIL.t5 VSUBS 0.097705f
C820 VTAIL.t4 VSUBS 0.097705f
C821 VTAIL.n126 VSUBS 0.490263f
C822 VTAIL.n127 VSUBS 0.925086f
C823 VTAIL.n128 VSUBS 0.0338f
C824 VTAIL.n129 VSUBS 0.031866f
C825 VTAIL.n130 VSUBS 0.017124f
C826 VTAIL.n131 VSUBS 0.040474f
C827 VTAIL.n132 VSUBS 0.018131f
C828 VTAIL.n133 VSUBS 0.122345f
C829 VTAIL.t1 VSUBS 0.088965f
C830 VTAIL.n134 VSUBS 0.030355f
C831 VTAIL.n135 VSUBS 0.025458f
C832 VTAIL.n136 VSUBS 0.017124f
C833 VTAIL.n137 VSUBS 0.420918f
C834 VTAIL.n138 VSUBS 0.031866f
C835 VTAIL.n139 VSUBS 0.017124f
C836 VTAIL.n140 VSUBS 0.018131f
C837 VTAIL.n141 VSUBS 0.040474f
C838 VTAIL.n142 VSUBS 0.093848f
C839 VTAIL.n143 VSUBS 0.018131f
C840 VTAIL.n144 VSUBS 0.017124f
C841 VTAIL.n145 VSUBS 0.075399f
C842 VTAIL.n146 VSUBS 0.047065f
C843 VTAIL.n147 VSUBS 1.25241f
C844 VTAIL.n148 VSUBS 0.0338f
C845 VTAIL.n149 VSUBS 0.031866f
C846 VTAIL.n150 VSUBS 0.017124f
C847 VTAIL.n151 VSUBS 0.040474f
C848 VTAIL.n152 VSUBS 0.018131f
C849 VTAIL.n153 VSUBS 0.122345f
C850 VTAIL.t9 VSUBS 0.088965f
C851 VTAIL.n154 VSUBS 0.030355f
C852 VTAIL.n155 VSUBS 0.025458f
C853 VTAIL.n156 VSUBS 0.017124f
C854 VTAIL.n157 VSUBS 0.420918f
C855 VTAIL.n158 VSUBS 0.031866f
C856 VTAIL.n159 VSUBS 0.017124f
C857 VTAIL.n160 VSUBS 0.018131f
C858 VTAIL.n161 VSUBS 0.040474f
C859 VTAIL.n162 VSUBS 0.093848f
C860 VTAIL.n163 VSUBS 0.018131f
C861 VTAIL.n164 VSUBS 0.017124f
C862 VTAIL.n165 VSUBS 0.075399f
C863 VTAIL.n166 VSUBS 0.047065f
C864 VTAIL.n167 VSUBS 1.24644f
C865 VDD2.t5 VSUBS 0.074294f
C866 VDD2.t1 VSUBS 0.074294f
C867 VDD2.n0 VSUBS 0.435233f
C868 VDD2.t6 VSUBS 0.074294f
C869 VDD2.t4 VSUBS 0.074294f
C870 VDD2.n1 VSUBS 0.435233f
C871 VDD2.n2 VSUBS 2.75556f
C872 VDD2.t3 VSUBS 0.074294f
C873 VDD2.t2 VSUBS 0.074294f
C874 VDD2.n3 VSUBS 0.429851f
C875 VDD2.n4 VSUBS 2.25025f
C876 VDD2.t7 VSUBS 0.074294f
C877 VDD2.t0 VSUBS 0.074294f
C878 VDD2.n5 VSUBS 0.435212f
C879 VN.n0 VSUBS 0.059502f
C880 VN.t5 VSUBS 0.98694f
C881 VN.n1 VSUBS 0.036974f
C882 VN.n2 VSUBS 0.045134f
C883 VN.t7 VSUBS 0.98694f
C884 VN.n3 VSUBS 0.089232f
C885 VN.n4 VSUBS 0.045134f
C886 VN.t3 VSUBS 0.98694f
C887 VN.n5 VSUBS 0.518081f
C888 VN.t6 VSUBS 1.26656f
C889 VN.n6 VSUBS 0.500108f
C890 VN.n7 VSUBS 0.384225f
C891 VN.n8 VSUBS 0.064277f
C892 VN.n9 VSUBS 0.089232f
C893 VN.n10 VSUBS 0.036454f
C894 VN.n11 VSUBS 0.045134f
C895 VN.n12 VSUBS 0.045134f
C896 VN.n13 VSUBS 0.045134f
C897 VN.n14 VSUBS 0.064277f
C898 VN.n15 VSUBS 0.401218f
C899 VN.n16 VSUBS 0.061798f
C900 VN.n17 VSUBS 0.090296f
C901 VN.n18 VSUBS 0.045134f
C902 VN.n19 VSUBS 0.045134f
C903 VN.n20 VSUBS 0.045134f
C904 VN.n21 VSUBS 0.087647f
C905 VN.n22 VSUBS 0.066757f
C906 VN.n23 VSUBS 0.537982f
C907 VN.n24 VSUBS 0.063195f
C908 VN.n25 VSUBS 0.059502f
C909 VN.t1 VSUBS 0.98694f
C910 VN.n26 VSUBS 0.036974f
C911 VN.n27 VSUBS 0.045134f
C912 VN.t4 VSUBS 0.98694f
C913 VN.n28 VSUBS 0.089232f
C914 VN.n29 VSUBS 0.045134f
C915 VN.t0 VSUBS 0.98694f
C916 VN.n30 VSUBS 0.518081f
C917 VN.t2 VSUBS 1.26656f
C918 VN.n31 VSUBS 0.500108f
C919 VN.n32 VSUBS 0.384225f
C920 VN.n33 VSUBS 0.064277f
C921 VN.n34 VSUBS 0.089232f
C922 VN.n35 VSUBS 0.036454f
C923 VN.n36 VSUBS 0.045134f
C924 VN.n37 VSUBS 0.045134f
C925 VN.n38 VSUBS 0.045134f
C926 VN.n39 VSUBS 0.064277f
C927 VN.n40 VSUBS 0.401218f
C928 VN.n41 VSUBS 0.061798f
C929 VN.n42 VSUBS 0.090296f
C930 VN.n43 VSUBS 0.045134f
C931 VN.n44 VSUBS 0.045134f
C932 VN.n45 VSUBS 0.045134f
C933 VN.n46 VSUBS 0.087647f
C934 VN.n47 VSUBS 0.066757f
C935 VN.n48 VSUBS 0.537982f
C936 VN.n49 VSUBS 1.99768f
.ends

