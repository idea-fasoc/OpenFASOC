* NGSPICE file created from diff_pair_sample_1221.ext - technology: sky130A

.subckt diff_pair_sample_1221 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=0.25
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=0.25
X2 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=0.25
X3 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=0.25
X4 VTAIL.t4 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=0.25
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=0.25
X6 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=0.25
X7 VTAIL.t5 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=0.25
X8 VDD2.t0 VN.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=0.25
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=0.25
X10 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=0.25
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=0.25
R0 VN.n0 VN.t3 1014.07
R1 VN.n0 VN.t1 1014.07
R2 VN.n1 VN.t2 1014.07
R3 VN.n1 VN.t0 1014.07
R4 VN VN.n1 198.333
R5 VN VN.n0 161.351
R6 VTAIL.n378 VTAIL.n336 289.615
R7 VTAIL.n42 VTAIL.n0 289.615
R8 VTAIL.n90 VTAIL.n48 289.615
R9 VTAIL.n138 VTAIL.n96 289.615
R10 VTAIL.n330 VTAIL.n288 289.615
R11 VTAIL.n282 VTAIL.n240 289.615
R12 VTAIL.n234 VTAIL.n192 289.615
R13 VTAIL.n186 VTAIL.n144 289.615
R14 VTAIL.n353 VTAIL.n352 185
R15 VTAIL.n355 VTAIL.n354 185
R16 VTAIL.n348 VTAIL.n347 185
R17 VTAIL.n361 VTAIL.n360 185
R18 VTAIL.n363 VTAIL.n362 185
R19 VTAIL.n344 VTAIL.n343 185
R20 VTAIL.n369 VTAIL.n368 185
R21 VTAIL.n371 VTAIL.n370 185
R22 VTAIL.n340 VTAIL.n339 185
R23 VTAIL.n377 VTAIL.n376 185
R24 VTAIL.n379 VTAIL.n378 185
R25 VTAIL.n17 VTAIL.n16 185
R26 VTAIL.n19 VTAIL.n18 185
R27 VTAIL.n12 VTAIL.n11 185
R28 VTAIL.n25 VTAIL.n24 185
R29 VTAIL.n27 VTAIL.n26 185
R30 VTAIL.n8 VTAIL.n7 185
R31 VTAIL.n33 VTAIL.n32 185
R32 VTAIL.n35 VTAIL.n34 185
R33 VTAIL.n4 VTAIL.n3 185
R34 VTAIL.n41 VTAIL.n40 185
R35 VTAIL.n43 VTAIL.n42 185
R36 VTAIL.n65 VTAIL.n64 185
R37 VTAIL.n67 VTAIL.n66 185
R38 VTAIL.n60 VTAIL.n59 185
R39 VTAIL.n73 VTAIL.n72 185
R40 VTAIL.n75 VTAIL.n74 185
R41 VTAIL.n56 VTAIL.n55 185
R42 VTAIL.n81 VTAIL.n80 185
R43 VTAIL.n83 VTAIL.n82 185
R44 VTAIL.n52 VTAIL.n51 185
R45 VTAIL.n89 VTAIL.n88 185
R46 VTAIL.n91 VTAIL.n90 185
R47 VTAIL.n113 VTAIL.n112 185
R48 VTAIL.n115 VTAIL.n114 185
R49 VTAIL.n108 VTAIL.n107 185
R50 VTAIL.n121 VTAIL.n120 185
R51 VTAIL.n123 VTAIL.n122 185
R52 VTAIL.n104 VTAIL.n103 185
R53 VTAIL.n129 VTAIL.n128 185
R54 VTAIL.n131 VTAIL.n130 185
R55 VTAIL.n100 VTAIL.n99 185
R56 VTAIL.n137 VTAIL.n136 185
R57 VTAIL.n139 VTAIL.n138 185
R58 VTAIL.n331 VTAIL.n330 185
R59 VTAIL.n329 VTAIL.n328 185
R60 VTAIL.n292 VTAIL.n291 185
R61 VTAIL.n323 VTAIL.n322 185
R62 VTAIL.n321 VTAIL.n320 185
R63 VTAIL.n296 VTAIL.n295 185
R64 VTAIL.n315 VTAIL.n314 185
R65 VTAIL.n313 VTAIL.n312 185
R66 VTAIL.n300 VTAIL.n299 185
R67 VTAIL.n307 VTAIL.n306 185
R68 VTAIL.n305 VTAIL.n304 185
R69 VTAIL.n283 VTAIL.n282 185
R70 VTAIL.n281 VTAIL.n280 185
R71 VTAIL.n244 VTAIL.n243 185
R72 VTAIL.n275 VTAIL.n274 185
R73 VTAIL.n273 VTAIL.n272 185
R74 VTAIL.n248 VTAIL.n247 185
R75 VTAIL.n267 VTAIL.n266 185
R76 VTAIL.n265 VTAIL.n264 185
R77 VTAIL.n252 VTAIL.n251 185
R78 VTAIL.n259 VTAIL.n258 185
R79 VTAIL.n257 VTAIL.n256 185
R80 VTAIL.n235 VTAIL.n234 185
R81 VTAIL.n233 VTAIL.n232 185
R82 VTAIL.n196 VTAIL.n195 185
R83 VTAIL.n227 VTAIL.n226 185
R84 VTAIL.n225 VTAIL.n224 185
R85 VTAIL.n200 VTAIL.n199 185
R86 VTAIL.n219 VTAIL.n218 185
R87 VTAIL.n217 VTAIL.n216 185
R88 VTAIL.n204 VTAIL.n203 185
R89 VTAIL.n211 VTAIL.n210 185
R90 VTAIL.n209 VTAIL.n208 185
R91 VTAIL.n187 VTAIL.n186 185
R92 VTAIL.n185 VTAIL.n184 185
R93 VTAIL.n148 VTAIL.n147 185
R94 VTAIL.n179 VTAIL.n178 185
R95 VTAIL.n177 VTAIL.n176 185
R96 VTAIL.n152 VTAIL.n151 185
R97 VTAIL.n171 VTAIL.n170 185
R98 VTAIL.n169 VTAIL.n168 185
R99 VTAIL.n156 VTAIL.n155 185
R100 VTAIL.n163 VTAIL.n162 185
R101 VTAIL.n161 VTAIL.n160 185
R102 VTAIL.n255 VTAIL.t0 147.659
R103 VTAIL.n207 VTAIL.t6 147.659
R104 VTAIL.n159 VTAIL.t5 147.659
R105 VTAIL.n351 VTAIL.t7 147.659
R106 VTAIL.n15 VTAIL.t4 147.659
R107 VTAIL.n63 VTAIL.t2 147.659
R108 VTAIL.n111 VTAIL.t1 147.659
R109 VTAIL.n303 VTAIL.t3 147.659
R110 VTAIL.n354 VTAIL.n353 104.615
R111 VTAIL.n354 VTAIL.n347 104.615
R112 VTAIL.n361 VTAIL.n347 104.615
R113 VTAIL.n362 VTAIL.n361 104.615
R114 VTAIL.n362 VTAIL.n343 104.615
R115 VTAIL.n369 VTAIL.n343 104.615
R116 VTAIL.n370 VTAIL.n369 104.615
R117 VTAIL.n370 VTAIL.n339 104.615
R118 VTAIL.n377 VTAIL.n339 104.615
R119 VTAIL.n378 VTAIL.n377 104.615
R120 VTAIL.n18 VTAIL.n17 104.615
R121 VTAIL.n18 VTAIL.n11 104.615
R122 VTAIL.n25 VTAIL.n11 104.615
R123 VTAIL.n26 VTAIL.n25 104.615
R124 VTAIL.n26 VTAIL.n7 104.615
R125 VTAIL.n33 VTAIL.n7 104.615
R126 VTAIL.n34 VTAIL.n33 104.615
R127 VTAIL.n34 VTAIL.n3 104.615
R128 VTAIL.n41 VTAIL.n3 104.615
R129 VTAIL.n42 VTAIL.n41 104.615
R130 VTAIL.n66 VTAIL.n65 104.615
R131 VTAIL.n66 VTAIL.n59 104.615
R132 VTAIL.n73 VTAIL.n59 104.615
R133 VTAIL.n74 VTAIL.n73 104.615
R134 VTAIL.n74 VTAIL.n55 104.615
R135 VTAIL.n81 VTAIL.n55 104.615
R136 VTAIL.n82 VTAIL.n81 104.615
R137 VTAIL.n82 VTAIL.n51 104.615
R138 VTAIL.n89 VTAIL.n51 104.615
R139 VTAIL.n90 VTAIL.n89 104.615
R140 VTAIL.n114 VTAIL.n113 104.615
R141 VTAIL.n114 VTAIL.n107 104.615
R142 VTAIL.n121 VTAIL.n107 104.615
R143 VTAIL.n122 VTAIL.n121 104.615
R144 VTAIL.n122 VTAIL.n103 104.615
R145 VTAIL.n129 VTAIL.n103 104.615
R146 VTAIL.n130 VTAIL.n129 104.615
R147 VTAIL.n130 VTAIL.n99 104.615
R148 VTAIL.n137 VTAIL.n99 104.615
R149 VTAIL.n138 VTAIL.n137 104.615
R150 VTAIL.n330 VTAIL.n329 104.615
R151 VTAIL.n329 VTAIL.n291 104.615
R152 VTAIL.n322 VTAIL.n291 104.615
R153 VTAIL.n322 VTAIL.n321 104.615
R154 VTAIL.n321 VTAIL.n295 104.615
R155 VTAIL.n314 VTAIL.n295 104.615
R156 VTAIL.n314 VTAIL.n313 104.615
R157 VTAIL.n313 VTAIL.n299 104.615
R158 VTAIL.n306 VTAIL.n299 104.615
R159 VTAIL.n306 VTAIL.n305 104.615
R160 VTAIL.n282 VTAIL.n281 104.615
R161 VTAIL.n281 VTAIL.n243 104.615
R162 VTAIL.n274 VTAIL.n243 104.615
R163 VTAIL.n274 VTAIL.n273 104.615
R164 VTAIL.n273 VTAIL.n247 104.615
R165 VTAIL.n266 VTAIL.n247 104.615
R166 VTAIL.n266 VTAIL.n265 104.615
R167 VTAIL.n265 VTAIL.n251 104.615
R168 VTAIL.n258 VTAIL.n251 104.615
R169 VTAIL.n258 VTAIL.n257 104.615
R170 VTAIL.n234 VTAIL.n233 104.615
R171 VTAIL.n233 VTAIL.n195 104.615
R172 VTAIL.n226 VTAIL.n195 104.615
R173 VTAIL.n226 VTAIL.n225 104.615
R174 VTAIL.n225 VTAIL.n199 104.615
R175 VTAIL.n218 VTAIL.n199 104.615
R176 VTAIL.n218 VTAIL.n217 104.615
R177 VTAIL.n217 VTAIL.n203 104.615
R178 VTAIL.n210 VTAIL.n203 104.615
R179 VTAIL.n210 VTAIL.n209 104.615
R180 VTAIL.n186 VTAIL.n185 104.615
R181 VTAIL.n185 VTAIL.n147 104.615
R182 VTAIL.n178 VTAIL.n147 104.615
R183 VTAIL.n178 VTAIL.n177 104.615
R184 VTAIL.n177 VTAIL.n151 104.615
R185 VTAIL.n170 VTAIL.n151 104.615
R186 VTAIL.n170 VTAIL.n169 104.615
R187 VTAIL.n169 VTAIL.n155 104.615
R188 VTAIL.n162 VTAIL.n155 104.615
R189 VTAIL.n162 VTAIL.n161 104.615
R190 VTAIL.n353 VTAIL.t7 52.3082
R191 VTAIL.n17 VTAIL.t4 52.3082
R192 VTAIL.n65 VTAIL.t2 52.3082
R193 VTAIL.n113 VTAIL.t1 52.3082
R194 VTAIL.n305 VTAIL.t3 52.3082
R195 VTAIL.n257 VTAIL.t0 52.3082
R196 VTAIL.n209 VTAIL.t6 52.3082
R197 VTAIL.n161 VTAIL.t5 52.3082
R198 VTAIL.n383 VTAIL.n382 30.052
R199 VTAIL.n47 VTAIL.n46 30.052
R200 VTAIL.n95 VTAIL.n94 30.052
R201 VTAIL.n143 VTAIL.n142 30.052
R202 VTAIL.n335 VTAIL.n334 30.052
R203 VTAIL.n287 VTAIL.n286 30.052
R204 VTAIL.n239 VTAIL.n238 30.052
R205 VTAIL.n191 VTAIL.n190 30.052
R206 VTAIL.n383 VTAIL.n335 20.4445
R207 VTAIL.n191 VTAIL.n143 20.4445
R208 VTAIL.n352 VTAIL.n351 15.6677
R209 VTAIL.n16 VTAIL.n15 15.6677
R210 VTAIL.n64 VTAIL.n63 15.6677
R211 VTAIL.n112 VTAIL.n111 15.6677
R212 VTAIL.n304 VTAIL.n303 15.6677
R213 VTAIL.n256 VTAIL.n255 15.6677
R214 VTAIL.n208 VTAIL.n207 15.6677
R215 VTAIL.n160 VTAIL.n159 15.6677
R216 VTAIL.n355 VTAIL.n350 12.8005
R217 VTAIL.n19 VTAIL.n14 12.8005
R218 VTAIL.n67 VTAIL.n62 12.8005
R219 VTAIL.n115 VTAIL.n110 12.8005
R220 VTAIL.n307 VTAIL.n302 12.8005
R221 VTAIL.n259 VTAIL.n254 12.8005
R222 VTAIL.n211 VTAIL.n206 12.8005
R223 VTAIL.n163 VTAIL.n158 12.8005
R224 VTAIL.n356 VTAIL.n348 12.0247
R225 VTAIL.n20 VTAIL.n12 12.0247
R226 VTAIL.n68 VTAIL.n60 12.0247
R227 VTAIL.n116 VTAIL.n108 12.0247
R228 VTAIL.n308 VTAIL.n300 12.0247
R229 VTAIL.n260 VTAIL.n252 12.0247
R230 VTAIL.n212 VTAIL.n204 12.0247
R231 VTAIL.n164 VTAIL.n156 12.0247
R232 VTAIL.n360 VTAIL.n359 11.249
R233 VTAIL.n24 VTAIL.n23 11.249
R234 VTAIL.n72 VTAIL.n71 11.249
R235 VTAIL.n120 VTAIL.n119 11.249
R236 VTAIL.n312 VTAIL.n311 11.249
R237 VTAIL.n264 VTAIL.n263 11.249
R238 VTAIL.n216 VTAIL.n215 11.249
R239 VTAIL.n168 VTAIL.n167 11.249
R240 VTAIL.n363 VTAIL.n346 10.4732
R241 VTAIL.n27 VTAIL.n10 10.4732
R242 VTAIL.n75 VTAIL.n58 10.4732
R243 VTAIL.n123 VTAIL.n106 10.4732
R244 VTAIL.n315 VTAIL.n298 10.4732
R245 VTAIL.n267 VTAIL.n250 10.4732
R246 VTAIL.n219 VTAIL.n202 10.4732
R247 VTAIL.n171 VTAIL.n154 10.4732
R248 VTAIL.n364 VTAIL.n344 9.69747
R249 VTAIL.n28 VTAIL.n8 9.69747
R250 VTAIL.n76 VTAIL.n56 9.69747
R251 VTAIL.n124 VTAIL.n104 9.69747
R252 VTAIL.n316 VTAIL.n296 9.69747
R253 VTAIL.n268 VTAIL.n248 9.69747
R254 VTAIL.n220 VTAIL.n200 9.69747
R255 VTAIL.n172 VTAIL.n152 9.69747
R256 VTAIL.n382 VTAIL.n381 9.45567
R257 VTAIL.n46 VTAIL.n45 9.45567
R258 VTAIL.n94 VTAIL.n93 9.45567
R259 VTAIL.n142 VTAIL.n141 9.45567
R260 VTAIL.n334 VTAIL.n333 9.45567
R261 VTAIL.n286 VTAIL.n285 9.45567
R262 VTAIL.n238 VTAIL.n237 9.45567
R263 VTAIL.n190 VTAIL.n189 9.45567
R264 VTAIL.n375 VTAIL.n374 9.3005
R265 VTAIL.n338 VTAIL.n337 9.3005
R266 VTAIL.n381 VTAIL.n380 9.3005
R267 VTAIL.n342 VTAIL.n341 9.3005
R268 VTAIL.n367 VTAIL.n366 9.3005
R269 VTAIL.n365 VTAIL.n364 9.3005
R270 VTAIL.n346 VTAIL.n345 9.3005
R271 VTAIL.n359 VTAIL.n358 9.3005
R272 VTAIL.n357 VTAIL.n356 9.3005
R273 VTAIL.n350 VTAIL.n349 9.3005
R274 VTAIL.n373 VTAIL.n372 9.3005
R275 VTAIL.n39 VTAIL.n38 9.3005
R276 VTAIL.n2 VTAIL.n1 9.3005
R277 VTAIL.n45 VTAIL.n44 9.3005
R278 VTAIL.n6 VTAIL.n5 9.3005
R279 VTAIL.n31 VTAIL.n30 9.3005
R280 VTAIL.n29 VTAIL.n28 9.3005
R281 VTAIL.n10 VTAIL.n9 9.3005
R282 VTAIL.n23 VTAIL.n22 9.3005
R283 VTAIL.n21 VTAIL.n20 9.3005
R284 VTAIL.n14 VTAIL.n13 9.3005
R285 VTAIL.n37 VTAIL.n36 9.3005
R286 VTAIL.n87 VTAIL.n86 9.3005
R287 VTAIL.n50 VTAIL.n49 9.3005
R288 VTAIL.n93 VTAIL.n92 9.3005
R289 VTAIL.n54 VTAIL.n53 9.3005
R290 VTAIL.n79 VTAIL.n78 9.3005
R291 VTAIL.n77 VTAIL.n76 9.3005
R292 VTAIL.n58 VTAIL.n57 9.3005
R293 VTAIL.n71 VTAIL.n70 9.3005
R294 VTAIL.n69 VTAIL.n68 9.3005
R295 VTAIL.n62 VTAIL.n61 9.3005
R296 VTAIL.n85 VTAIL.n84 9.3005
R297 VTAIL.n135 VTAIL.n134 9.3005
R298 VTAIL.n98 VTAIL.n97 9.3005
R299 VTAIL.n141 VTAIL.n140 9.3005
R300 VTAIL.n102 VTAIL.n101 9.3005
R301 VTAIL.n127 VTAIL.n126 9.3005
R302 VTAIL.n125 VTAIL.n124 9.3005
R303 VTAIL.n106 VTAIL.n105 9.3005
R304 VTAIL.n119 VTAIL.n118 9.3005
R305 VTAIL.n117 VTAIL.n116 9.3005
R306 VTAIL.n110 VTAIL.n109 9.3005
R307 VTAIL.n133 VTAIL.n132 9.3005
R308 VTAIL.n290 VTAIL.n289 9.3005
R309 VTAIL.n327 VTAIL.n326 9.3005
R310 VTAIL.n325 VTAIL.n324 9.3005
R311 VTAIL.n294 VTAIL.n293 9.3005
R312 VTAIL.n319 VTAIL.n318 9.3005
R313 VTAIL.n317 VTAIL.n316 9.3005
R314 VTAIL.n298 VTAIL.n297 9.3005
R315 VTAIL.n311 VTAIL.n310 9.3005
R316 VTAIL.n309 VTAIL.n308 9.3005
R317 VTAIL.n302 VTAIL.n301 9.3005
R318 VTAIL.n333 VTAIL.n332 9.3005
R319 VTAIL.n242 VTAIL.n241 9.3005
R320 VTAIL.n285 VTAIL.n284 9.3005
R321 VTAIL.n279 VTAIL.n278 9.3005
R322 VTAIL.n277 VTAIL.n276 9.3005
R323 VTAIL.n246 VTAIL.n245 9.3005
R324 VTAIL.n271 VTAIL.n270 9.3005
R325 VTAIL.n269 VTAIL.n268 9.3005
R326 VTAIL.n250 VTAIL.n249 9.3005
R327 VTAIL.n263 VTAIL.n262 9.3005
R328 VTAIL.n261 VTAIL.n260 9.3005
R329 VTAIL.n254 VTAIL.n253 9.3005
R330 VTAIL.n194 VTAIL.n193 9.3005
R331 VTAIL.n237 VTAIL.n236 9.3005
R332 VTAIL.n231 VTAIL.n230 9.3005
R333 VTAIL.n229 VTAIL.n228 9.3005
R334 VTAIL.n198 VTAIL.n197 9.3005
R335 VTAIL.n223 VTAIL.n222 9.3005
R336 VTAIL.n221 VTAIL.n220 9.3005
R337 VTAIL.n202 VTAIL.n201 9.3005
R338 VTAIL.n215 VTAIL.n214 9.3005
R339 VTAIL.n213 VTAIL.n212 9.3005
R340 VTAIL.n206 VTAIL.n205 9.3005
R341 VTAIL.n146 VTAIL.n145 9.3005
R342 VTAIL.n189 VTAIL.n188 9.3005
R343 VTAIL.n183 VTAIL.n182 9.3005
R344 VTAIL.n181 VTAIL.n180 9.3005
R345 VTAIL.n150 VTAIL.n149 9.3005
R346 VTAIL.n175 VTAIL.n174 9.3005
R347 VTAIL.n173 VTAIL.n172 9.3005
R348 VTAIL.n154 VTAIL.n153 9.3005
R349 VTAIL.n167 VTAIL.n166 9.3005
R350 VTAIL.n165 VTAIL.n164 9.3005
R351 VTAIL.n158 VTAIL.n157 9.3005
R352 VTAIL.n368 VTAIL.n367 8.92171
R353 VTAIL.n382 VTAIL.n336 8.92171
R354 VTAIL.n32 VTAIL.n31 8.92171
R355 VTAIL.n46 VTAIL.n0 8.92171
R356 VTAIL.n80 VTAIL.n79 8.92171
R357 VTAIL.n94 VTAIL.n48 8.92171
R358 VTAIL.n128 VTAIL.n127 8.92171
R359 VTAIL.n142 VTAIL.n96 8.92171
R360 VTAIL.n334 VTAIL.n288 8.92171
R361 VTAIL.n320 VTAIL.n319 8.92171
R362 VTAIL.n286 VTAIL.n240 8.92171
R363 VTAIL.n272 VTAIL.n271 8.92171
R364 VTAIL.n238 VTAIL.n192 8.92171
R365 VTAIL.n224 VTAIL.n223 8.92171
R366 VTAIL.n190 VTAIL.n144 8.92171
R367 VTAIL.n176 VTAIL.n175 8.92171
R368 VTAIL.n371 VTAIL.n342 8.14595
R369 VTAIL.n380 VTAIL.n379 8.14595
R370 VTAIL.n35 VTAIL.n6 8.14595
R371 VTAIL.n44 VTAIL.n43 8.14595
R372 VTAIL.n83 VTAIL.n54 8.14595
R373 VTAIL.n92 VTAIL.n91 8.14595
R374 VTAIL.n131 VTAIL.n102 8.14595
R375 VTAIL.n140 VTAIL.n139 8.14595
R376 VTAIL.n332 VTAIL.n331 8.14595
R377 VTAIL.n323 VTAIL.n294 8.14595
R378 VTAIL.n284 VTAIL.n283 8.14595
R379 VTAIL.n275 VTAIL.n246 8.14595
R380 VTAIL.n236 VTAIL.n235 8.14595
R381 VTAIL.n227 VTAIL.n198 8.14595
R382 VTAIL.n188 VTAIL.n187 8.14595
R383 VTAIL.n179 VTAIL.n150 8.14595
R384 VTAIL.n372 VTAIL.n340 7.3702
R385 VTAIL.n376 VTAIL.n338 7.3702
R386 VTAIL.n36 VTAIL.n4 7.3702
R387 VTAIL.n40 VTAIL.n2 7.3702
R388 VTAIL.n84 VTAIL.n52 7.3702
R389 VTAIL.n88 VTAIL.n50 7.3702
R390 VTAIL.n132 VTAIL.n100 7.3702
R391 VTAIL.n136 VTAIL.n98 7.3702
R392 VTAIL.n328 VTAIL.n290 7.3702
R393 VTAIL.n324 VTAIL.n292 7.3702
R394 VTAIL.n280 VTAIL.n242 7.3702
R395 VTAIL.n276 VTAIL.n244 7.3702
R396 VTAIL.n232 VTAIL.n194 7.3702
R397 VTAIL.n228 VTAIL.n196 7.3702
R398 VTAIL.n184 VTAIL.n146 7.3702
R399 VTAIL.n180 VTAIL.n148 7.3702
R400 VTAIL.n375 VTAIL.n340 6.59444
R401 VTAIL.n376 VTAIL.n375 6.59444
R402 VTAIL.n39 VTAIL.n4 6.59444
R403 VTAIL.n40 VTAIL.n39 6.59444
R404 VTAIL.n87 VTAIL.n52 6.59444
R405 VTAIL.n88 VTAIL.n87 6.59444
R406 VTAIL.n135 VTAIL.n100 6.59444
R407 VTAIL.n136 VTAIL.n135 6.59444
R408 VTAIL.n328 VTAIL.n327 6.59444
R409 VTAIL.n327 VTAIL.n292 6.59444
R410 VTAIL.n280 VTAIL.n279 6.59444
R411 VTAIL.n279 VTAIL.n244 6.59444
R412 VTAIL.n232 VTAIL.n231 6.59444
R413 VTAIL.n231 VTAIL.n196 6.59444
R414 VTAIL.n184 VTAIL.n183 6.59444
R415 VTAIL.n183 VTAIL.n148 6.59444
R416 VTAIL.n372 VTAIL.n371 5.81868
R417 VTAIL.n379 VTAIL.n338 5.81868
R418 VTAIL.n36 VTAIL.n35 5.81868
R419 VTAIL.n43 VTAIL.n2 5.81868
R420 VTAIL.n84 VTAIL.n83 5.81868
R421 VTAIL.n91 VTAIL.n50 5.81868
R422 VTAIL.n132 VTAIL.n131 5.81868
R423 VTAIL.n139 VTAIL.n98 5.81868
R424 VTAIL.n331 VTAIL.n290 5.81868
R425 VTAIL.n324 VTAIL.n323 5.81868
R426 VTAIL.n283 VTAIL.n242 5.81868
R427 VTAIL.n276 VTAIL.n275 5.81868
R428 VTAIL.n235 VTAIL.n194 5.81868
R429 VTAIL.n228 VTAIL.n227 5.81868
R430 VTAIL.n187 VTAIL.n146 5.81868
R431 VTAIL.n180 VTAIL.n179 5.81868
R432 VTAIL.n368 VTAIL.n342 5.04292
R433 VTAIL.n380 VTAIL.n336 5.04292
R434 VTAIL.n32 VTAIL.n6 5.04292
R435 VTAIL.n44 VTAIL.n0 5.04292
R436 VTAIL.n80 VTAIL.n54 5.04292
R437 VTAIL.n92 VTAIL.n48 5.04292
R438 VTAIL.n128 VTAIL.n102 5.04292
R439 VTAIL.n140 VTAIL.n96 5.04292
R440 VTAIL.n332 VTAIL.n288 5.04292
R441 VTAIL.n320 VTAIL.n294 5.04292
R442 VTAIL.n284 VTAIL.n240 5.04292
R443 VTAIL.n272 VTAIL.n246 5.04292
R444 VTAIL.n236 VTAIL.n192 5.04292
R445 VTAIL.n224 VTAIL.n198 5.04292
R446 VTAIL.n188 VTAIL.n144 5.04292
R447 VTAIL.n176 VTAIL.n150 5.04292
R448 VTAIL.n351 VTAIL.n349 4.38563
R449 VTAIL.n15 VTAIL.n13 4.38563
R450 VTAIL.n63 VTAIL.n61 4.38563
R451 VTAIL.n111 VTAIL.n109 4.38563
R452 VTAIL.n303 VTAIL.n301 4.38563
R453 VTAIL.n255 VTAIL.n253 4.38563
R454 VTAIL.n207 VTAIL.n205 4.38563
R455 VTAIL.n159 VTAIL.n157 4.38563
R456 VTAIL.n367 VTAIL.n344 4.26717
R457 VTAIL.n31 VTAIL.n8 4.26717
R458 VTAIL.n79 VTAIL.n56 4.26717
R459 VTAIL.n127 VTAIL.n104 4.26717
R460 VTAIL.n319 VTAIL.n296 4.26717
R461 VTAIL.n271 VTAIL.n248 4.26717
R462 VTAIL.n223 VTAIL.n200 4.26717
R463 VTAIL.n175 VTAIL.n152 4.26717
R464 VTAIL.n364 VTAIL.n363 3.49141
R465 VTAIL.n28 VTAIL.n27 3.49141
R466 VTAIL.n76 VTAIL.n75 3.49141
R467 VTAIL.n124 VTAIL.n123 3.49141
R468 VTAIL.n316 VTAIL.n315 3.49141
R469 VTAIL.n268 VTAIL.n267 3.49141
R470 VTAIL.n220 VTAIL.n219 3.49141
R471 VTAIL.n172 VTAIL.n171 3.49141
R472 VTAIL.n360 VTAIL.n346 2.71565
R473 VTAIL.n24 VTAIL.n10 2.71565
R474 VTAIL.n72 VTAIL.n58 2.71565
R475 VTAIL.n120 VTAIL.n106 2.71565
R476 VTAIL.n312 VTAIL.n298 2.71565
R477 VTAIL.n264 VTAIL.n250 2.71565
R478 VTAIL.n216 VTAIL.n202 2.71565
R479 VTAIL.n168 VTAIL.n154 2.71565
R480 VTAIL.n359 VTAIL.n348 1.93989
R481 VTAIL.n23 VTAIL.n12 1.93989
R482 VTAIL.n71 VTAIL.n60 1.93989
R483 VTAIL.n119 VTAIL.n108 1.93989
R484 VTAIL.n311 VTAIL.n300 1.93989
R485 VTAIL.n263 VTAIL.n252 1.93989
R486 VTAIL.n215 VTAIL.n204 1.93989
R487 VTAIL.n167 VTAIL.n156 1.93989
R488 VTAIL.n356 VTAIL.n355 1.16414
R489 VTAIL.n20 VTAIL.n19 1.16414
R490 VTAIL.n68 VTAIL.n67 1.16414
R491 VTAIL.n116 VTAIL.n115 1.16414
R492 VTAIL.n308 VTAIL.n307 1.16414
R493 VTAIL.n260 VTAIL.n259 1.16414
R494 VTAIL.n212 VTAIL.n211 1.16414
R495 VTAIL.n164 VTAIL.n163 1.16414
R496 VTAIL.n239 VTAIL.n191 0.5005
R497 VTAIL.n335 VTAIL.n287 0.5005
R498 VTAIL.n143 VTAIL.n95 0.5005
R499 VTAIL.n287 VTAIL.n239 0.470328
R500 VTAIL.n95 VTAIL.n47 0.470328
R501 VTAIL.n352 VTAIL.n350 0.388379
R502 VTAIL.n16 VTAIL.n14 0.388379
R503 VTAIL.n64 VTAIL.n62 0.388379
R504 VTAIL.n112 VTAIL.n110 0.388379
R505 VTAIL.n304 VTAIL.n302 0.388379
R506 VTAIL.n256 VTAIL.n254 0.388379
R507 VTAIL.n208 VTAIL.n206 0.388379
R508 VTAIL.n160 VTAIL.n158 0.388379
R509 VTAIL VTAIL.n47 0.30869
R510 VTAIL VTAIL.n383 0.19231
R511 VTAIL.n357 VTAIL.n349 0.155672
R512 VTAIL.n358 VTAIL.n357 0.155672
R513 VTAIL.n358 VTAIL.n345 0.155672
R514 VTAIL.n365 VTAIL.n345 0.155672
R515 VTAIL.n366 VTAIL.n365 0.155672
R516 VTAIL.n366 VTAIL.n341 0.155672
R517 VTAIL.n373 VTAIL.n341 0.155672
R518 VTAIL.n374 VTAIL.n373 0.155672
R519 VTAIL.n374 VTAIL.n337 0.155672
R520 VTAIL.n381 VTAIL.n337 0.155672
R521 VTAIL.n21 VTAIL.n13 0.155672
R522 VTAIL.n22 VTAIL.n21 0.155672
R523 VTAIL.n22 VTAIL.n9 0.155672
R524 VTAIL.n29 VTAIL.n9 0.155672
R525 VTAIL.n30 VTAIL.n29 0.155672
R526 VTAIL.n30 VTAIL.n5 0.155672
R527 VTAIL.n37 VTAIL.n5 0.155672
R528 VTAIL.n38 VTAIL.n37 0.155672
R529 VTAIL.n38 VTAIL.n1 0.155672
R530 VTAIL.n45 VTAIL.n1 0.155672
R531 VTAIL.n69 VTAIL.n61 0.155672
R532 VTAIL.n70 VTAIL.n69 0.155672
R533 VTAIL.n70 VTAIL.n57 0.155672
R534 VTAIL.n77 VTAIL.n57 0.155672
R535 VTAIL.n78 VTAIL.n77 0.155672
R536 VTAIL.n78 VTAIL.n53 0.155672
R537 VTAIL.n85 VTAIL.n53 0.155672
R538 VTAIL.n86 VTAIL.n85 0.155672
R539 VTAIL.n86 VTAIL.n49 0.155672
R540 VTAIL.n93 VTAIL.n49 0.155672
R541 VTAIL.n117 VTAIL.n109 0.155672
R542 VTAIL.n118 VTAIL.n117 0.155672
R543 VTAIL.n118 VTAIL.n105 0.155672
R544 VTAIL.n125 VTAIL.n105 0.155672
R545 VTAIL.n126 VTAIL.n125 0.155672
R546 VTAIL.n126 VTAIL.n101 0.155672
R547 VTAIL.n133 VTAIL.n101 0.155672
R548 VTAIL.n134 VTAIL.n133 0.155672
R549 VTAIL.n134 VTAIL.n97 0.155672
R550 VTAIL.n141 VTAIL.n97 0.155672
R551 VTAIL.n333 VTAIL.n289 0.155672
R552 VTAIL.n326 VTAIL.n289 0.155672
R553 VTAIL.n326 VTAIL.n325 0.155672
R554 VTAIL.n325 VTAIL.n293 0.155672
R555 VTAIL.n318 VTAIL.n293 0.155672
R556 VTAIL.n318 VTAIL.n317 0.155672
R557 VTAIL.n317 VTAIL.n297 0.155672
R558 VTAIL.n310 VTAIL.n297 0.155672
R559 VTAIL.n310 VTAIL.n309 0.155672
R560 VTAIL.n309 VTAIL.n301 0.155672
R561 VTAIL.n285 VTAIL.n241 0.155672
R562 VTAIL.n278 VTAIL.n241 0.155672
R563 VTAIL.n278 VTAIL.n277 0.155672
R564 VTAIL.n277 VTAIL.n245 0.155672
R565 VTAIL.n270 VTAIL.n245 0.155672
R566 VTAIL.n270 VTAIL.n269 0.155672
R567 VTAIL.n269 VTAIL.n249 0.155672
R568 VTAIL.n262 VTAIL.n249 0.155672
R569 VTAIL.n262 VTAIL.n261 0.155672
R570 VTAIL.n261 VTAIL.n253 0.155672
R571 VTAIL.n237 VTAIL.n193 0.155672
R572 VTAIL.n230 VTAIL.n193 0.155672
R573 VTAIL.n230 VTAIL.n229 0.155672
R574 VTAIL.n229 VTAIL.n197 0.155672
R575 VTAIL.n222 VTAIL.n197 0.155672
R576 VTAIL.n222 VTAIL.n221 0.155672
R577 VTAIL.n221 VTAIL.n201 0.155672
R578 VTAIL.n214 VTAIL.n201 0.155672
R579 VTAIL.n214 VTAIL.n213 0.155672
R580 VTAIL.n213 VTAIL.n205 0.155672
R581 VTAIL.n189 VTAIL.n145 0.155672
R582 VTAIL.n182 VTAIL.n145 0.155672
R583 VTAIL.n182 VTAIL.n181 0.155672
R584 VTAIL.n181 VTAIL.n149 0.155672
R585 VTAIL.n174 VTAIL.n149 0.155672
R586 VTAIL.n174 VTAIL.n173 0.155672
R587 VTAIL.n173 VTAIL.n153 0.155672
R588 VTAIL.n166 VTAIL.n153 0.155672
R589 VTAIL.n166 VTAIL.n165 0.155672
R590 VTAIL.n165 VTAIL.n157 0.155672
R591 VDD2.n2 VDD2.n0 94.597
R592 VDD2.n2 VDD2.n1 61.8048
R593 VDD2.n1 VDD2.t1 2.2582
R594 VDD2.n1 VDD2.t3 2.2582
R595 VDD2.n0 VDD2.t2 2.2582
R596 VDD2.n0 VDD2.t0 2.2582
R597 VDD2 VDD2.n2 0.0586897
R598 B.n280 B.t4 1069.73
R599 B.n278 B.t8 1069.73
R600 B.n68 B.t11 1069.73
R601 B.n65 B.t15 1069.73
R602 B.n487 B.n486 585
R603 B.n215 B.n64 585
R604 B.n214 B.n213 585
R605 B.n212 B.n211 585
R606 B.n210 B.n209 585
R607 B.n208 B.n207 585
R608 B.n206 B.n205 585
R609 B.n204 B.n203 585
R610 B.n202 B.n201 585
R611 B.n200 B.n199 585
R612 B.n198 B.n197 585
R613 B.n196 B.n195 585
R614 B.n194 B.n193 585
R615 B.n192 B.n191 585
R616 B.n190 B.n189 585
R617 B.n188 B.n187 585
R618 B.n186 B.n185 585
R619 B.n184 B.n183 585
R620 B.n182 B.n181 585
R621 B.n180 B.n179 585
R622 B.n178 B.n177 585
R623 B.n176 B.n175 585
R624 B.n174 B.n173 585
R625 B.n172 B.n171 585
R626 B.n170 B.n169 585
R627 B.n168 B.n167 585
R628 B.n166 B.n165 585
R629 B.n164 B.n163 585
R630 B.n162 B.n161 585
R631 B.n160 B.n159 585
R632 B.n158 B.n157 585
R633 B.n156 B.n155 585
R634 B.n154 B.n153 585
R635 B.n152 B.n151 585
R636 B.n150 B.n149 585
R637 B.n148 B.n147 585
R638 B.n146 B.n145 585
R639 B.n144 B.n143 585
R640 B.n142 B.n141 585
R641 B.n140 B.n139 585
R642 B.n138 B.n137 585
R643 B.n136 B.n135 585
R644 B.n134 B.n133 585
R645 B.n132 B.n131 585
R646 B.n130 B.n129 585
R647 B.n128 B.n127 585
R648 B.n126 B.n125 585
R649 B.n124 B.n123 585
R650 B.n122 B.n121 585
R651 B.n120 B.n119 585
R652 B.n118 B.n117 585
R653 B.n116 B.n115 585
R654 B.n114 B.n113 585
R655 B.n112 B.n111 585
R656 B.n110 B.n109 585
R657 B.n108 B.n107 585
R658 B.n106 B.n105 585
R659 B.n104 B.n103 585
R660 B.n102 B.n101 585
R661 B.n100 B.n99 585
R662 B.n98 B.n97 585
R663 B.n96 B.n95 585
R664 B.n94 B.n93 585
R665 B.n92 B.n91 585
R666 B.n90 B.n89 585
R667 B.n88 B.n87 585
R668 B.n86 B.n85 585
R669 B.n84 B.n83 585
R670 B.n82 B.n81 585
R671 B.n80 B.n79 585
R672 B.n78 B.n77 585
R673 B.n76 B.n75 585
R674 B.n74 B.n73 585
R675 B.n72 B.n71 585
R676 B.n485 B.n27 585
R677 B.n490 B.n27 585
R678 B.n484 B.n26 585
R679 B.n491 B.n26 585
R680 B.n483 B.n482 585
R681 B.n482 B.n22 585
R682 B.n481 B.n21 585
R683 B.n497 B.n21 585
R684 B.n480 B.n20 585
R685 B.n498 B.n20 585
R686 B.n479 B.n19 585
R687 B.n499 B.n19 585
R688 B.n478 B.n477 585
R689 B.n477 B.n15 585
R690 B.n476 B.n14 585
R691 B.n505 B.n14 585
R692 B.n475 B.n13 585
R693 B.n506 B.n13 585
R694 B.n474 B.n12 585
R695 B.n507 B.n12 585
R696 B.n473 B.n472 585
R697 B.n472 B.n11 585
R698 B.n471 B.n7 585
R699 B.n513 B.n7 585
R700 B.n470 B.n6 585
R701 B.n514 B.n6 585
R702 B.n469 B.n5 585
R703 B.n515 B.n5 585
R704 B.n468 B.n467 585
R705 B.n467 B.n4 585
R706 B.n466 B.n216 585
R707 B.n466 B.n465 585
R708 B.n455 B.n217 585
R709 B.n458 B.n217 585
R710 B.n457 B.n456 585
R711 B.n459 B.n457 585
R712 B.n454 B.n221 585
R713 B.n225 B.n221 585
R714 B.n453 B.n452 585
R715 B.n452 B.n451 585
R716 B.n223 B.n222 585
R717 B.n224 B.n223 585
R718 B.n444 B.n443 585
R719 B.n445 B.n444 585
R720 B.n442 B.n230 585
R721 B.n230 B.n229 585
R722 B.n441 B.n440 585
R723 B.n440 B.n439 585
R724 B.n232 B.n231 585
R725 B.n233 B.n232 585
R726 B.n432 B.n431 585
R727 B.n433 B.n432 585
R728 B.n430 B.n238 585
R729 B.n238 B.n237 585
R730 B.n425 B.n424 585
R731 B.n423 B.n277 585
R732 B.n422 B.n276 585
R733 B.n427 B.n276 585
R734 B.n421 B.n420 585
R735 B.n419 B.n418 585
R736 B.n417 B.n416 585
R737 B.n415 B.n414 585
R738 B.n413 B.n412 585
R739 B.n411 B.n410 585
R740 B.n409 B.n408 585
R741 B.n407 B.n406 585
R742 B.n405 B.n404 585
R743 B.n403 B.n402 585
R744 B.n401 B.n400 585
R745 B.n399 B.n398 585
R746 B.n397 B.n396 585
R747 B.n395 B.n394 585
R748 B.n393 B.n392 585
R749 B.n391 B.n390 585
R750 B.n389 B.n388 585
R751 B.n387 B.n386 585
R752 B.n385 B.n384 585
R753 B.n383 B.n382 585
R754 B.n381 B.n380 585
R755 B.n379 B.n378 585
R756 B.n377 B.n376 585
R757 B.n375 B.n374 585
R758 B.n373 B.n372 585
R759 B.n371 B.n370 585
R760 B.n369 B.n368 585
R761 B.n367 B.n366 585
R762 B.n365 B.n364 585
R763 B.n362 B.n361 585
R764 B.n360 B.n359 585
R765 B.n358 B.n357 585
R766 B.n356 B.n355 585
R767 B.n354 B.n353 585
R768 B.n352 B.n351 585
R769 B.n350 B.n349 585
R770 B.n348 B.n347 585
R771 B.n346 B.n345 585
R772 B.n344 B.n343 585
R773 B.n341 B.n340 585
R774 B.n339 B.n338 585
R775 B.n337 B.n336 585
R776 B.n335 B.n334 585
R777 B.n333 B.n332 585
R778 B.n331 B.n330 585
R779 B.n329 B.n328 585
R780 B.n327 B.n326 585
R781 B.n325 B.n324 585
R782 B.n323 B.n322 585
R783 B.n321 B.n320 585
R784 B.n319 B.n318 585
R785 B.n317 B.n316 585
R786 B.n315 B.n314 585
R787 B.n313 B.n312 585
R788 B.n311 B.n310 585
R789 B.n309 B.n308 585
R790 B.n307 B.n306 585
R791 B.n305 B.n304 585
R792 B.n303 B.n302 585
R793 B.n301 B.n300 585
R794 B.n299 B.n298 585
R795 B.n297 B.n296 585
R796 B.n295 B.n294 585
R797 B.n293 B.n292 585
R798 B.n291 B.n290 585
R799 B.n289 B.n288 585
R800 B.n287 B.n286 585
R801 B.n285 B.n284 585
R802 B.n283 B.n282 585
R803 B.n240 B.n239 585
R804 B.n429 B.n428 585
R805 B.n428 B.n427 585
R806 B.n236 B.n235 585
R807 B.n237 B.n236 585
R808 B.n435 B.n434 585
R809 B.n434 B.n433 585
R810 B.n436 B.n234 585
R811 B.n234 B.n233 585
R812 B.n438 B.n437 585
R813 B.n439 B.n438 585
R814 B.n228 B.n227 585
R815 B.n229 B.n228 585
R816 B.n447 B.n446 585
R817 B.n446 B.n445 585
R818 B.n448 B.n226 585
R819 B.n226 B.n224 585
R820 B.n450 B.n449 585
R821 B.n451 B.n450 585
R822 B.n220 B.n219 585
R823 B.n225 B.n220 585
R824 B.n461 B.n460 585
R825 B.n460 B.n459 585
R826 B.n462 B.n218 585
R827 B.n458 B.n218 585
R828 B.n464 B.n463 585
R829 B.n465 B.n464 585
R830 B.n2 B.n0 585
R831 B.n4 B.n2 585
R832 B.n3 B.n1 585
R833 B.n514 B.n3 585
R834 B.n512 B.n511 585
R835 B.n513 B.n512 585
R836 B.n510 B.n8 585
R837 B.n11 B.n8 585
R838 B.n509 B.n508 585
R839 B.n508 B.n507 585
R840 B.n10 B.n9 585
R841 B.n506 B.n10 585
R842 B.n504 B.n503 585
R843 B.n505 B.n504 585
R844 B.n502 B.n16 585
R845 B.n16 B.n15 585
R846 B.n501 B.n500 585
R847 B.n500 B.n499 585
R848 B.n18 B.n17 585
R849 B.n498 B.n18 585
R850 B.n496 B.n495 585
R851 B.n497 B.n496 585
R852 B.n494 B.n23 585
R853 B.n23 B.n22 585
R854 B.n493 B.n492 585
R855 B.n492 B.n491 585
R856 B.n25 B.n24 585
R857 B.n490 B.n25 585
R858 B.n517 B.n516 585
R859 B.n516 B.n515 585
R860 B.n425 B.n236 530.939
R861 B.n71 B.n25 530.939
R862 B.n428 B.n238 530.939
R863 B.n487 B.n27 530.939
R864 B.n489 B.n488 256.663
R865 B.n489 B.n63 256.663
R866 B.n489 B.n62 256.663
R867 B.n489 B.n61 256.663
R868 B.n489 B.n60 256.663
R869 B.n489 B.n59 256.663
R870 B.n489 B.n58 256.663
R871 B.n489 B.n57 256.663
R872 B.n489 B.n56 256.663
R873 B.n489 B.n55 256.663
R874 B.n489 B.n54 256.663
R875 B.n489 B.n53 256.663
R876 B.n489 B.n52 256.663
R877 B.n489 B.n51 256.663
R878 B.n489 B.n50 256.663
R879 B.n489 B.n49 256.663
R880 B.n489 B.n48 256.663
R881 B.n489 B.n47 256.663
R882 B.n489 B.n46 256.663
R883 B.n489 B.n45 256.663
R884 B.n489 B.n44 256.663
R885 B.n489 B.n43 256.663
R886 B.n489 B.n42 256.663
R887 B.n489 B.n41 256.663
R888 B.n489 B.n40 256.663
R889 B.n489 B.n39 256.663
R890 B.n489 B.n38 256.663
R891 B.n489 B.n37 256.663
R892 B.n489 B.n36 256.663
R893 B.n489 B.n35 256.663
R894 B.n489 B.n34 256.663
R895 B.n489 B.n33 256.663
R896 B.n489 B.n32 256.663
R897 B.n489 B.n31 256.663
R898 B.n489 B.n30 256.663
R899 B.n489 B.n29 256.663
R900 B.n489 B.n28 256.663
R901 B.n427 B.n426 256.663
R902 B.n427 B.n241 256.663
R903 B.n427 B.n242 256.663
R904 B.n427 B.n243 256.663
R905 B.n427 B.n244 256.663
R906 B.n427 B.n245 256.663
R907 B.n427 B.n246 256.663
R908 B.n427 B.n247 256.663
R909 B.n427 B.n248 256.663
R910 B.n427 B.n249 256.663
R911 B.n427 B.n250 256.663
R912 B.n427 B.n251 256.663
R913 B.n427 B.n252 256.663
R914 B.n427 B.n253 256.663
R915 B.n427 B.n254 256.663
R916 B.n427 B.n255 256.663
R917 B.n427 B.n256 256.663
R918 B.n427 B.n257 256.663
R919 B.n427 B.n258 256.663
R920 B.n427 B.n259 256.663
R921 B.n427 B.n260 256.663
R922 B.n427 B.n261 256.663
R923 B.n427 B.n262 256.663
R924 B.n427 B.n263 256.663
R925 B.n427 B.n264 256.663
R926 B.n427 B.n265 256.663
R927 B.n427 B.n266 256.663
R928 B.n427 B.n267 256.663
R929 B.n427 B.n268 256.663
R930 B.n427 B.n269 256.663
R931 B.n427 B.n270 256.663
R932 B.n427 B.n271 256.663
R933 B.n427 B.n272 256.663
R934 B.n427 B.n273 256.663
R935 B.n427 B.n274 256.663
R936 B.n427 B.n275 256.663
R937 B.n280 B.t7 237.994
R938 B.n65 B.t16 237.994
R939 B.n278 B.t10 237.994
R940 B.n68 B.t13 237.994
R941 B.n281 B.t6 226.745
R942 B.n66 B.t17 226.745
R943 B.n279 B.t9 226.745
R944 B.n69 B.t14 226.745
R945 B.n434 B.n236 163.367
R946 B.n434 B.n234 163.367
R947 B.n438 B.n234 163.367
R948 B.n438 B.n228 163.367
R949 B.n446 B.n228 163.367
R950 B.n446 B.n226 163.367
R951 B.n450 B.n226 163.367
R952 B.n450 B.n220 163.367
R953 B.n460 B.n220 163.367
R954 B.n460 B.n218 163.367
R955 B.n464 B.n218 163.367
R956 B.n464 B.n2 163.367
R957 B.n516 B.n2 163.367
R958 B.n516 B.n3 163.367
R959 B.n512 B.n3 163.367
R960 B.n512 B.n8 163.367
R961 B.n508 B.n8 163.367
R962 B.n508 B.n10 163.367
R963 B.n504 B.n10 163.367
R964 B.n504 B.n16 163.367
R965 B.n500 B.n16 163.367
R966 B.n500 B.n18 163.367
R967 B.n496 B.n18 163.367
R968 B.n496 B.n23 163.367
R969 B.n492 B.n23 163.367
R970 B.n492 B.n25 163.367
R971 B.n277 B.n276 163.367
R972 B.n420 B.n276 163.367
R973 B.n418 B.n417 163.367
R974 B.n414 B.n413 163.367
R975 B.n410 B.n409 163.367
R976 B.n406 B.n405 163.367
R977 B.n402 B.n401 163.367
R978 B.n398 B.n397 163.367
R979 B.n394 B.n393 163.367
R980 B.n390 B.n389 163.367
R981 B.n386 B.n385 163.367
R982 B.n382 B.n381 163.367
R983 B.n378 B.n377 163.367
R984 B.n374 B.n373 163.367
R985 B.n370 B.n369 163.367
R986 B.n366 B.n365 163.367
R987 B.n361 B.n360 163.367
R988 B.n357 B.n356 163.367
R989 B.n353 B.n352 163.367
R990 B.n349 B.n348 163.367
R991 B.n345 B.n344 163.367
R992 B.n340 B.n339 163.367
R993 B.n336 B.n335 163.367
R994 B.n332 B.n331 163.367
R995 B.n328 B.n327 163.367
R996 B.n324 B.n323 163.367
R997 B.n320 B.n319 163.367
R998 B.n316 B.n315 163.367
R999 B.n312 B.n311 163.367
R1000 B.n308 B.n307 163.367
R1001 B.n304 B.n303 163.367
R1002 B.n300 B.n299 163.367
R1003 B.n296 B.n295 163.367
R1004 B.n292 B.n291 163.367
R1005 B.n288 B.n287 163.367
R1006 B.n284 B.n283 163.367
R1007 B.n428 B.n240 163.367
R1008 B.n432 B.n238 163.367
R1009 B.n432 B.n232 163.367
R1010 B.n440 B.n232 163.367
R1011 B.n440 B.n230 163.367
R1012 B.n444 B.n230 163.367
R1013 B.n444 B.n223 163.367
R1014 B.n452 B.n223 163.367
R1015 B.n452 B.n221 163.367
R1016 B.n457 B.n221 163.367
R1017 B.n457 B.n217 163.367
R1018 B.n466 B.n217 163.367
R1019 B.n467 B.n466 163.367
R1020 B.n467 B.n5 163.367
R1021 B.n6 B.n5 163.367
R1022 B.n7 B.n6 163.367
R1023 B.n472 B.n7 163.367
R1024 B.n472 B.n12 163.367
R1025 B.n13 B.n12 163.367
R1026 B.n14 B.n13 163.367
R1027 B.n477 B.n14 163.367
R1028 B.n477 B.n19 163.367
R1029 B.n20 B.n19 163.367
R1030 B.n21 B.n20 163.367
R1031 B.n482 B.n21 163.367
R1032 B.n482 B.n26 163.367
R1033 B.n27 B.n26 163.367
R1034 B.n75 B.n74 163.367
R1035 B.n79 B.n78 163.367
R1036 B.n83 B.n82 163.367
R1037 B.n87 B.n86 163.367
R1038 B.n91 B.n90 163.367
R1039 B.n95 B.n94 163.367
R1040 B.n99 B.n98 163.367
R1041 B.n103 B.n102 163.367
R1042 B.n107 B.n106 163.367
R1043 B.n111 B.n110 163.367
R1044 B.n115 B.n114 163.367
R1045 B.n119 B.n118 163.367
R1046 B.n123 B.n122 163.367
R1047 B.n127 B.n126 163.367
R1048 B.n131 B.n130 163.367
R1049 B.n135 B.n134 163.367
R1050 B.n139 B.n138 163.367
R1051 B.n143 B.n142 163.367
R1052 B.n147 B.n146 163.367
R1053 B.n151 B.n150 163.367
R1054 B.n155 B.n154 163.367
R1055 B.n159 B.n158 163.367
R1056 B.n163 B.n162 163.367
R1057 B.n167 B.n166 163.367
R1058 B.n171 B.n170 163.367
R1059 B.n175 B.n174 163.367
R1060 B.n179 B.n178 163.367
R1061 B.n183 B.n182 163.367
R1062 B.n187 B.n186 163.367
R1063 B.n191 B.n190 163.367
R1064 B.n195 B.n194 163.367
R1065 B.n199 B.n198 163.367
R1066 B.n203 B.n202 163.367
R1067 B.n207 B.n206 163.367
R1068 B.n211 B.n210 163.367
R1069 B.n213 B.n64 163.367
R1070 B.n427 B.n237 108.71
R1071 B.n490 B.n489 108.71
R1072 B.n426 B.n425 71.676
R1073 B.n420 B.n241 71.676
R1074 B.n417 B.n242 71.676
R1075 B.n413 B.n243 71.676
R1076 B.n409 B.n244 71.676
R1077 B.n405 B.n245 71.676
R1078 B.n401 B.n246 71.676
R1079 B.n397 B.n247 71.676
R1080 B.n393 B.n248 71.676
R1081 B.n389 B.n249 71.676
R1082 B.n385 B.n250 71.676
R1083 B.n381 B.n251 71.676
R1084 B.n377 B.n252 71.676
R1085 B.n373 B.n253 71.676
R1086 B.n369 B.n254 71.676
R1087 B.n365 B.n255 71.676
R1088 B.n360 B.n256 71.676
R1089 B.n356 B.n257 71.676
R1090 B.n352 B.n258 71.676
R1091 B.n348 B.n259 71.676
R1092 B.n344 B.n260 71.676
R1093 B.n339 B.n261 71.676
R1094 B.n335 B.n262 71.676
R1095 B.n331 B.n263 71.676
R1096 B.n327 B.n264 71.676
R1097 B.n323 B.n265 71.676
R1098 B.n319 B.n266 71.676
R1099 B.n315 B.n267 71.676
R1100 B.n311 B.n268 71.676
R1101 B.n307 B.n269 71.676
R1102 B.n303 B.n270 71.676
R1103 B.n299 B.n271 71.676
R1104 B.n295 B.n272 71.676
R1105 B.n291 B.n273 71.676
R1106 B.n287 B.n274 71.676
R1107 B.n283 B.n275 71.676
R1108 B.n71 B.n28 71.676
R1109 B.n75 B.n29 71.676
R1110 B.n79 B.n30 71.676
R1111 B.n83 B.n31 71.676
R1112 B.n87 B.n32 71.676
R1113 B.n91 B.n33 71.676
R1114 B.n95 B.n34 71.676
R1115 B.n99 B.n35 71.676
R1116 B.n103 B.n36 71.676
R1117 B.n107 B.n37 71.676
R1118 B.n111 B.n38 71.676
R1119 B.n115 B.n39 71.676
R1120 B.n119 B.n40 71.676
R1121 B.n123 B.n41 71.676
R1122 B.n127 B.n42 71.676
R1123 B.n131 B.n43 71.676
R1124 B.n135 B.n44 71.676
R1125 B.n139 B.n45 71.676
R1126 B.n143 B.n46 71.676
R1127 B.n147 B.n47 71.676
R1128 B.n151 B.n48 71.676
R1129 B.n155 B.n49 71.676
R1130 B.n159 B.n50 71.676
R1131 B.n163 B.n51 71.676
R1132 B.n167 B.n52 71.676
R1133 B.n171 B.n53 71.676
R1134 B.n175 B.n54 71.676
R1135 B.n179 B.n55 71.676
R1136 B.n183 B.n56 71.676
R1137 B.n187 B.n57 71.676
R1138 B.n191 B.n58 71.676
R1139 B.n195 B.n59 71.676
R1140 B.n199 B.n60 71.676
R1141 B.n203 B.n61 71.676
R1142 B.n207 B.n62 71.676
R1143 B.n211 B.n63 71.676
R1144 B.n488 B.n64 71.676
R1145 B.n488 B.n487 71.676
R1146 B.n213 B.n63 71.676
R1147 B.n210 B.n62 71.676
R1148 B.n206 B.n61 71.676
R1149 B.n202 B.n60 71.676
R1150 B.n198 B.n59 71.676
R1151 B.n194 B.n58 71.676
R1152 B.n190 B.n57 71.676
R1153 B.n186 B.n56 71.676
R1154 B.n182 B.n55 71.676
R1155 B.n178 B.n54 71.676
R1156 B.n174 B.n53 71.676
R1157 B.n170 B.n52 71.676
R1158 B.n166 B.n51 71.676
R1159 B.n162 B.n50 71.676
R1160 B.n158 B.n49 71.676
R1161 B.n154 B.n48 71.676
R1162 B.n150 B.n47 71.676
R1163 B.n146 B.n46 71.676
R1164 B.n142 B.n45 71.676
R1165 B.n138 B.n44 71.676
R1166 B.n134 B.n43 71.676
R1167 B.n130 B.n42 71.676
R1168 B.n126 B.n41 71.676
R1169 B.n122 B.n40 71.676
R1170 B.n118 B.n39 71.676
R1171 B.n114 B.n38 71.676
R1172 B.n110 B.n37 71.676
R1173 B.n106 B.n36 71.676
R1174 B.n102 B.n35 71.676
R1175 B.n98 B.n34 71.676
R1176 B.n94 B.n33 71.676
R1177 B.n90 B.n32 71.676
R1178 B.n86 B.n31 71.676
R1179 B.n82 B.n30 71.676
R1180 B.n78 B.n29 71.676
R1181 B.n74 B.n28 71.676
R1182 B.n426 B.n277 71.676
R1183 B.n418 B.n241 71.676
R1184 B.n414 B.n242 71.676
R1185 B.n410 B.n243 71.676
R1186 B.n406 B.n244 71.676
R1187 B.n402 B.n245 71.676
R1188 B.n398 B.n246 71.676
R1189 B.n394 B.n247 71.676
R1190 B.n390 B.n248 71.676
R1191 B.n386 B.n249 71.676
R1192 B.n382 B.n250 71.676
R1193 B.n378 B.n251 71.676
R1194 B.n374 B.n252 71.676
R1195 B.n370 B.n253 71.676
R1196 B.n366 B.n254 71.676
R1197 B.n361 B.n255 71.676
R1198 B.n357 B.n256 71.676
R1199 B.n353 B.n257 71.676
R1200 B.n349 B.n258 71.676
R1201 B.n345 B.n259 71.676
R1202 B.n340 B.n260 71.676
R1203 B.n336 B.n261 71.676
R1204 B.n332 B.n262 71.676
R1205 B.n328 B.n263 71.676
R1206 B.n324 B.n264 71.676
R1207 B.n320 B.n265 71.676
R1208 B.n316 B.n266 71.676
R1209 B.n312 B.n267 71.676
R1210 B.n308 B.n268 71.676
R1211 B.n304 B.n269 71.676
R1212 B.n300 B.n270 71.676
R1213 B.n296 B.n271 71.676
R1214 B.n292 B.n272 71.676
R1215 B.n288 B.n273 71.676
R1216 B.n284 B.n274 71.676
R1217 B.n275 B.n240 71.676
R1218 B.n342 B.n281 59.5399
R1219 B.n363 B.n279 59.5399
R1220 B.n70 B.n69 59.5399
R1221 B.n67 B.n66 59.5399
R1222 B.n433 B.n237 53.1822
R1223 B.n433 B.n233 53.1822
R1224 B.n439 B.n233 53.1822
R1225 B.n445 B.n229 53.1822
R1226 B.n445 B.n224 53.1822
R1227 B.n451 B.n224 53.1822
R1228 B.n451 B.n225 53.1822
R1229 B.n459 B.n458 53.1822
R1230 B.n465 B.n4 53.1822
R1231 B.n515 B.n4 53.1822
R1232 B.n515 B.n514 53.1822
R1233 B.n514 B.n513 53.1822
R1234 B.n507 B.n11 53.1822
R1235 B.n506 B.n505 53.1822
R1236 B.n505 B.n15 53.1822
R1237 B.n499 B.n15 53.1822
R1238 B.n499 B.n498 53.1822
R1239 B.n497 B.n22 53.1822
R1240 B.n491 B.n22 53.1822
R1241 B.n491 B.n490 53.1822
R1242 B.n439 B.t5 49.2717
R1243 B.t12 B.n497 49.2717
R1244 B.n225 B.t1 44.5792
R1245 B.t3 B.n506 44.5792
R1246 B.n72 B.n24 34.4981
R1247 B.n486 B.n485 34.4981
R1248 B.n430 B.n429 34.4981
R1249 B.n424 B.n235 34.4981
R1250 B.n458 B.t2 28.9376
R1251 B.n11 B.t0 28.9376
R1252 B.n465 B.t2 24.2451
R1253 B.n513 B.t0 24.2451
R1254 B B.n517 18.0485
R1255 B.n281 B.n280 11.249
R1256 B.n279 B.n278 11.249
R1257 B.n69 B.n68 11.249
R1258 B.n66 B.n65 11.249
R1259 B.n73 B.n72 10.6151
R1260 B.n76 B.n73 10.6151
R1261 B.n77 B.n76 10.6151
R1262 B.n80 B.n77 10.6151
R1263 B.n81 B.n80 10.6151
R1264 B.n84 B.n81 10.6151
R1265 B.n85 B.n84 10.6151
R1266 B.n88 B.n85 10.6151
R1267 B.n89 B.n88 10.6151
R1268 B.n92 B.n89 10.6151
R1269 B.n93 B.n92 10.6151
R1270 B.n96 B.n93 10.6151
R1271 B.n97 B.n96 10.6151
R1272 B.n100 B.n97 10.6151
R1273 B.n101 B.n100 10.6151
R1274 B.n104 B.n101 10.6151
R1275 B.n105 B.n104 10.6151
R1276 B.n108 B.n105 10.6151
R1277 B.n109 B.n108 10.6151
R1278 B.n112 B.n109 10.6151
R1279 B.n113 B.n112 10.6151
R1280 B.n116 B.n113 10.6151
R1281 B.n117 B.n116 10.6151
R1282 B.n120 B.n117 10.6151
R1283 B.n121 B.n120 10.6151
R1284 B.n124 B.n121 10.6151
R1285 B.n125 B.n124 10.6151
R1286 B.n128 B.n125 10.6151
R1287 B.n129 B.n128 10.6151
R1288 B.n132 B.n129 10.6151
R1289 B.n133 B.n132 10.6151
R1290 B.n137 B.n136 10.6151
R1291 B.n140 B.n137 10.6151
R1292 B.n141 B.n140 10.6151
R1293 B.n144 B.n141 10.6151
R1294 B.n145 B.n144 10.6151
R1295 B.n148 B.n145 10.6151
R1296 B.n149 B.n148 10.6151
R1297 B.n152 B.n149 10.6151
R1298 B.n153 B.n152 10.6151
R1299 B.n157 B.n156 10.6151
R1300 B.n160 B.n157 10.6151
R1301 B.n161 B.n160 10.6151
R1302 B.n164 B.n161 10.6151
R1303 B.n165 B.n164 10.6151
R1304 B.n168 B.n165 10.6151
R1305 B.n169 B.n168 10.6151
R1306 B.n172 B.n169 10.6151
R1307 B.n173 B.n172 10.6151
R1308 B.n176 B.n173 10.6151
R1309 B.n177 B.n176 10.6151
R1310 B.n180 B.n177 10.6151
R1311 B.n181 B.n180 10.6151
R1312 B.n184 B.n181 10.6151
R1313 B.n185 B.n184 10.6151
R1314 B.n188 B.n185 10.6151
R1315 B.n189 B.n188 10.6151
R1316 B.n192 B.n189 10.6151
R1317 B.n193 B.n192 10.6151
R1318 B.n196 B.n193 10.6151
R1319 B.n197 B.n196 10.6151
R1320 B.n200 B.n197 10.6151
R1321 B.n201 B.n200 10.6151
R1322 B.n204 B.n201 10.6151
R1323 B.n205 B.n204 10.6151
R1324 B.n208 B.n205 10.6151
R1325 B.n209 B.n208 10.6151
R1326 B.n212 B.n209 10.6151
R1327 B.n214 B.n212 10.6151
R1328 B.n215 B.n214 10.6151
R1329 B.n486 B.n215 10.6151
R1330 B.n431 B.n430 10.6151
R1331 B.n431 B.n231 10.6151
R1332 B.n441 B.n231 10.6151
R1333 B.n442 B.n441 10.6151
R1334 B.n443 B.n442 10.6151
R1335 B.n443 B.n222 10.6151
R1336 B.n453 B.n222 10.6151
R1337 B.n454 B.n453 10.6151
R1338 B.n456 B.n454 10.6151
R1339 B.n456 B.n455 10.6151
R1340 B.n455 B.n216 10.6151
R1341 B.n468 B.n216 10.6151
R1342 B.n469 B.n468 10.6151
R1343 B.n470 B.n469 10.6151
R1344 B.n471 B.n470 10.6151
R1345 B.n473 B.n471 10.6151
R1346 B.n474 B.n473 10.6151
R1347 B.n475 B.n474 10.6151
R1348 B.n476 B.n475 10.6151
R1349 B.n478 B.n476 10.6151
R1350 B.n479 B.n478 10.6151
R1351 B.n480 B.n479 10.6151
R1352 B.n481 B.n480 10.6151
R1353 B.n483 B.n481 10.6151
R1354 B.n484 B.n483 10.6151
R1355 B.n485 B.n484 10.6151
R1356 B.n424 B.n423 10.6151
R1357 B.n423 B.n422 10.6151
R1358 B.n422 B.n421 10.6151
R1359 B.n421 B.n419 10.6151
R1360 B.n419 B.n416 10.6151
R1361 B.n416 B.n415 10.6151
R1362 B.n415 B.n412 10.6151
R1363 B.n412 B.n411 10.6151
R1364 B.n411 B.n408 10.6151
R1365 B.n408 B.n407 10.6151
R1366 B.n407 B.n404 10.6151
R1367 B.n404 B.n403 10.6151
R1368 B.n403 B.n400 10.6151
R1369 B.n400 B.n399 10.6151
R1370 B.n399 B.n396 10.6151
R1371 B.n396 B.n395 10.6151
R1372 B.n395 B.n392 10.6151
R1373 B.n392 B.n391 10.6151
R1374 B.n391 B.n388 10.6151
R1375 B.n388 B.n387 10.6151
R1376 B.n387 B.n384 10.6151
R1377 B.n384 B.n383 10.6151
R1378 B.n383 B.n380 10.6151
R1379 B.n380 B.n379 10.6151
R1380 B.n379 B.n376 10.6151
R1381 B.n376 B.n375 10.6151
R1382 B.n375 B.n372 10.6151
R1383 B.n372 B.n371 10.6151
R1384 B.n371 B.n368 10.6151
R1385 B.n368 B.n367 10.6151
R1386 B.n367 B.n364 10.6151
R1387 B.n362 B.n359 10.6151
R1388 B.n359 B.n358 10.6151
R1389 B.n358 B.n355 10.6151
R1390 B.n355 B.n354 10.6151
R1391 B.n354 B.n351 10.6151
R1392 B.n351 B.n350 10.6151
R1393 B.n350 B.n347 10.6151
R1394 B.n347 B.n346 10.6151
R1395 B.n346 B.n343 10.6151
R1396 B.n341 B.n338 10.6151
R1397 B.n338 B.n337 10.6151
R1398 B.n337 B.n334 10.6151
R1399 B.n334 B.n333 10.6151
R1400 B.n333 B.n330 10.6151
R1401 B.n330 B.n329 10.6151
R1402 B.n329 B.n326 10.6151
R1403 B.n326 B.n325 10.6151
R1404 B.n325 B.n322 10.6151
R1405 B.n322 B.n321 10.6151
R1406 B.n321 B.n318 10.6151
R1407 B.n318 B.n317 10.6151
R1408 B.n317 B.n314 10.6151
R1409 B.n314 B.n313 10.6151
R1410 B.n313 B.n310 10.6151
R1411 B.n310 B.n309 10.6151
R1412 B.n309 B.n306 10.6151
R1413 B.n306 B.n305 10.6151
R1414 B.n305 B.n302 10.6151
R1415 B.n302 B.n301 10.6151
R1416 B.n301 B.n298 10.6151
R1417 B.n298 B.n297 10.6151
R1418 B.n297 B.n294 10.6151
R1419 B.n294 B.n293 10.6151
R1420 B.n293 B.n290 10.6151
R1421 B.n290 B.n289 10.6151
R1422 B.n289 B.n286 10.6151
R1423 B.n286 B.n285 10.6151
R1424 B.n285 B.n282 10.6151
R1425 B.n282 B.n239 10.6151
R1426 B.n429 B.n239 10.6151
R1427 B.n435 B.n235 10.6151
R1428 B.n436 B.n435 10.6151
R1429 B.n437 B.n436 10.6151
R1430 B.n437 B.n227 10.6151
R1431 B.n447 B.n227 10.6151
R1432 B.n448 B.n447 10.6151
R1433 B.n449 B.n448 10.6151
R1434 B.n449 B.n219 10.6151
R1435 B.n461 B.n219 10.6151
R1436 B.n462 B.n461 10.6151
R1437 B.n463 B.n462 10.6151
R1438 B.n463 B.n0 10.6151
R1439 B.n511 B.n1 10.6151
R1440 B.n511 B.n510 10.6151
R1441 B.n510 B.n509 10.6151
R1442 B.n509 B.n9 10.6151
R1443 B.n503 B.n9 10.6151
R1444 B.n503 B.n502 10.6151
R1445 B.n502 B.n501 10.6151
R1446 B.n501 B.n17 10.6151
R1447 B.n495 B.n17 10.6151
R1448 B.n495 B.n494 10.6151
R1449 B.n494 B.n493 10.6151
R1450 B.n493 B.n24 10.6151
R1451 B.n133 B.n70 8.74196
R1452 B.n156 B.n67 8.74196
R1453 B.n364 B.n363 8.74196
R1454 B.n342 B.n341 8.74196
R1455 B.n459 B.t1 8.60341
R1456 B.n507 B.t3 8.60341
R1457 B.t5 B.n229 3.91092
R1458 B.n498 B.t12 3.91092
R1459 B.n517 B.n0 2.81026
R1460 B.n517 B.n1 2.81026
R1461 B.n136 B.n70 1.87367
R1462 B.n153 B.n67 1.87367
R1463 B.n363 B.n362 1.87367
R1464 B.n343 B.n342 1.87367
R1465 VP.n1 VP.t1 1014.07
R1466 VP.n1 VP.t0 1014.07
R1467 VP.n0 VP.t3 1014.07
R1468 VP.n0 VP.t2 1014.07
R1469 VP.n2 VP.n0 197.952
R1470 VP.n2 VP.n1 161.3
R1471 VP VP.n2 0.0516364
R1472 VDD1 VDD1.n1 95.1218
R1473 VDD1 VDD1.n0 61.863
R1474 VDD1.n0 VDD1.t0 2.2582
R1475 VDD1.n0 VDD1.t1 2.2582
R1476 VDD1.n1 VDD1.t3 2.2582
R1477 VDD1.n1 VDD1.t2 2.2582
C0 VDD2 VP 0.24591f
C1 VDD2 VTAIL 7.76851f
C2 VDD1 VP 1.55687f
C3 VDD1 VTAIL 7.73006f
C4 VN VP 3.89565f
C5 VN VTAIL 1.05863f
C6 VDD2 VDD1 0.468258f
C7 VP VTAIL 1.07274f
C8 VDD2 VN 1.45912f
C9 VN VDD1 0.148015f
C10 VDD2 B 2.186081f
C11 VDD1 B 5.3237f
C12 VTAIL B 6.309138f
C13 VN B 6.10357f
C14 VP B 3.719769f
C15 VDD1.t0 B 0.194094f
C16 VDD1.t1 B 0.194094f
C17 VDD1.n0 B 1.68151f
C18 VDD1.t3 B 0.194094f
C19 VDD1.t2 B 0.194094f
C20 VDD1.n1 B 2.18353f
C21 VP.t3 B 0.240146f
C22 VP.t2 B 0.240146f
C23 VP.n0 B 0.439633f
C24 VP.t0 B 0.240146f
C25 VP.t1 B 0.240146f
C26 VP.n1 B 0.20985f
C27 VP.n2 B 2.27367f
C28 VDD2.t2 B 0.199292f
C29 VDD2.t0 B 0.199292f
C30 VDD2.n0 B 2.21622f
C31 VDD2.t1 B 0.199292f
C32 VDD2.t3 B 0.199292f
C33 VDD2.n1 B 1.72626f
C34 VDD2.n2 B 3.00783f
C35 VTAIL.n0 B 0.025773f
C36 VTAIL.n1 B 0.017906f
C37 VTAIL.n2 B 0.009622f
C38 VTAIL.n3 B 0.022743f
C39 VTAIL.n4 B 0.010188f
C40 VTAIL.n5 B 0.017906f
C41 VTAIL.n6 B 0.009622f
C42 VTAIL.n7 B 0.022743f
C43 VTAIL.n8 B 0.010188f
C44 VTAIL.n9 B 0.017906f
C45 VTAIL.n10 B 0.009622f
C46 VTAIL.n11 B 0.022743f
C47 VTAIL.n12 B 0.010188f
C48 VTAIL.n13 B 0.653715f
C49 VTAIL.n14 B 0.009622f
C50 VTAIL.t4 B 0.037125f
C51 VTAIL.n15 B 0.088835f
C52 VTAIL.n16 B 0.013435f
C53 VTAIL.n17 B 0.017057f
C54 VTAIL.n18 B 0.022743f
C55 VTAIL.n19 B 0.010188f
C56 VTAIL.n20 B 0.009622f
C57 VTAIL.n21 B 0.017906f
C58 VTAIL.n22 B 0.017906f
C59 VTAIL.n23 B 0.009622f
C60 VTAIL.n24 B 0.010188f
C61 VTAIL.n25 B 0.022743f
C62 VTAIL.n26 B 0.022743f
C63 VTAIL.n27 B 0.010188f
C64 VTAIL.n28 B 0.009622f
C65 VTAIL.n29 B 0.017906f
C66 VTAIL.n30 B 0.017906f
C67 VTAIL.n31 B 0.009622f
C68 VTAIL.n32 B 0.010188f
C69 VTAIL.n33 B 0.022743f
C70 VTAIL.n34 B 0.022743f
C71 VTAIL.n35 B 0.010188f
C72 VTAIL.n36 B 0.009622f
C73 VTAIL.n37 B 0.017906f
C74 VTAIL.n38 B 0.017906f
C75 VTAIL.n39 B 0.009622f
C76 VTAIL.n40 B 0.010188f
C77 VTAIL.n41 B 0.022743f
C78 VTAIL.n42 B 0.050303f
C79 VTAIL.n43 B 0.010188f
C80 VTAIL.n44 B 0.009622f
C81 VTAIL.n45 B 0.038698f
C82 VTAIL.n46 B 0.028171f
C83 VTAIL.n47 B 0.058667f
C84 VTAIL.n48 B 0.025773f
C85 VTAIL.n49 B 0.017906f
C86 VTAIL.n50 B 0.009622f
C87 VTAIL.n51 B 0.022743f
C88 VTAIL.n52 B 0.010188f
C89 VTAIL.n53 B 0.017906f
C90 VTAIL.n54 B 0.009622f
C91 VTAIL.n55 B 0.022743f
C92 VTAIL.n56 B 0.010188f
C93 VTAIL.n57 B 0.017906f
C94 VTAIL.n58 B 0.009622f
C95 VTAIL.n59 B 0.022743f
C96 VTAIL.n60 B 0.010188f
C97 VTAIL.n61 B 0.653715f
C98 VTAIL.n62 B 0.009622f
C99 VTAIL.t2 B 0.037125f
C100 VTAIL.n63 B 0.088835f
C101 VTAIL.n64 B 0.013435f
C102 VTAIL.n65 B 0.017057f
C103 VTAIL.n66 B 0.022743f
C104 VTAIL.n67 B 0.010188f
C105 VTAIL.n68 B 0.009622f
C106 VTAIL.n69 B 0.017906f
C107 VTAIL.n70 B 0.017906f
C108 VTAIL.n71 B 0.009622f
C109 VTAIL.n72 B 0.010188f
C110 VTAIL.n73 B 0.022743f
C111 VTAIL.n74 B 0.022743f
C112 VTAIL.n75 B 0.010188f
C113 VTAIL.n76 B 0.009622f
C114 VTAIL.n77 B 0.017906f
C115 VTAIL.n78 B 0.017906f
C116 VTAIL.n79 B 0.009622f
C117 VTAIL.n80 B 0.010188f
C118 VTAIL.n81 B 0.022743f
C119 VTAIL.n82 B 0.022743f
C120 VTAIL.n83 B 0.010188f
C121 VTAIL.n84 B 0.009622f
C122 VTAIL.n85 B 0.017906f
C123 VTAIL.n86 B 0.017906f
C124 VTAIL.n87 B 0.009622f
C125 VTAIL.n88 B 0.010188f
C126 VTAIL.n89 B 0.022743f
C127 VTAIL.n90 B 0.050303f
C128 VTAIL.n91 B 0.010188f
C129 VTAIL.n92 B 0.009622f
C130 VTAIL.n93 B 0.038698f
C131 VTAIL.n94 B 0.028171f
C132 VTAIL.n95 B 0.069734f
C133 VTAIL.n96 B 0.025773f
C134 VTAIL.n97 B 0.017906f
C135 VTAIL.n98 B 0.009622f
C136 VTAIL.n99 B 0.022743f
C137 VTAIL.n100 B 0.010188f
C138 VTAIL.n101 B 0.017906f
C139 VTAIL.n102 B 0.009622f
C140 VTAIL.n103 B 0.022743f
C141 VTAIL.n104 B 0.010188f
C142 VTAIL.n105 B 0.017906f
C143 VTAIL.n106 B 0.009622f
C144 VTAIL.n107 B 0.022743f
C145 VTAIL.n108 B 0.010188f
C146 VTAIL.n109 B 0.653715f
C147 VTAIL.n110 B 0.009622f
C148 VTAIL.t1 B 0.037125f
C149 VTAIL.n111 B 0.088835f
C150 VTAIL.n112 B 0.013435f
C151 VTAIL.n113 B 0.017057f
C152 VTAIL.n114 B 0.022743f
C153 VTAIL.n115 B 0.010188f
C154 VTAIL.n116 B 0.009622f
C155 VTAIL.n117 B 0.017906f
C156 VTAIL.n118 B 0.017906f
C157 VTAIL.n119 B 0.009622f
C158 VTAIL.n120 B 0.010188f
C159 VTAIL.n121 B 0.022743f
C160 VTAIL.n122 B 0.022743f
C161 VTAIL.n123 B 0.010188f
C162 VTAIL.n124 B 0.009622f
C163 VTAIL.n125 B 0.017906f
C164 VTAIL.n126 B 0.017906f
C165 VTAIL.n127 B 0.009622f
C166 VTAIL.n128 B 0.010188f
C167 VTAIL.n129 B 0.022743f
C168 VTAIL.n130 B 0.022743f
C169 VTAIL.n131 B 0.010188f
C170 VTAIL.n132 B 0.009622f
C171 VTAIL.n133 B 0.017906f
C172 VTAIL.n134 B 0.017906f
C173 VTAIL.n135 B 0.009622f
C174 VTAIL.n136 B 0.010188f
C175 VTAIL.n137 B 0.022743f
C176 VTAIL.n138 B 0.050303f
C177 VTAIL.n139 B 0.010188f
C178 VTAIL.n140 B 0.009622f
C179 VTAIL.n141 B 0.038698f
C180 VTAIL.n142 B 0.028171f
C181 VTAIL.n143 B 0.751917f
C182 VTAIL.n144 B 0.025773f
C183 VTAIL.n145 B 0.017906f
C184 VTAIL.n146 B 0.009622f
C185 VTAIL.n147 B 0.022743f
C186 VTAIL.n148 B 0.010188f
C187 VTAIL.n149 B 0.017906f
C188 VTAIL.n150 B 0.009622f
C189 VTAIL.n151 B 0.022743f
C190 VTAIL.n152 B 0.010188f
C191 VTAIL.n153 B 0.017906f
C192 VTAIL.n154 B 0.009622f
C193 VTAIL.n155 B 0.022743f
C194 VTAIL.n156 B 0.010188f
C195 VTAIL.n157 B 0.653715f
C196 VTAIL.n158 B 0.009622f
C197 VTAIL.t5 B 0.037125f
C198 VTAIL.n159 B 0.088835f
C199 VTAIL.n160 B 0.013435f
C200 VTAIL.n161 B 0.017057f
C201 VTAIL.n162 B 0.022743f
C202 VTAIL.n163 B 0.010188f
C203 VTAIL.n164 B 0.009622f
C204 VTAIL.n165 B 0.017906f
C205 VTAIL.n166 B 0.017906f
C206 VTAIL.n167 B 0.009622f
C207 VTAIL.n168 B 0.010188f
C208 VTAIL.n169 B 0.022743f
C209 VTAIL.n170 B 0.022743f
C210 VTAIL.n171 B 0.010188f
C211 VTAIL.n172 B 0.009622f
C212 VTAIL.n173 B 0.017906f
C213 VTAIL.n174 B 0.017906f
C214 VTAIL.n175 B 0.009622f
C215 VTAIL.n176 B 0.010188f
C216 VTAIL.n177 B 0.022743f
C217 VTAIL.n178 B 0.022743f
C218 VTAIL.n179 B 0.010188f
C219 VTAIL.n180 B 0.009622f
C220 VTAIL.n181 B 0.017906f
C221 VTAIL.n182 B 0.017906f
C222 VTAIL.n183 B 0.009622f
C223 VTAIL.n184 B 0.010188f
C224 VTAIL.n185 B 0.022743f
C225 VTAIL.n186 B 0.050303f
C226 VTAIL.n187 B 0.010188f
C227 VTAIL.n188 B 0.009622f
C228 VTAIL.n189 B 0.038698f
C229 VTAIL.n190 B 0.028171f
C230 VTAIL.n191 B 0.751917f
C231 VTAIL.n192 B 0.025773f
C232 VTAIL.n193 B 0.017906f
C233 VTAIL.n194 B 0.009622f
C234 VTAIL.n195 B 0.022743f
C235 VTAIL.n196 B 0.010188f
C236 VTAIL.n197 B 0.017906f
C237 VTAIL.n198 B 0.009622f
C238 VTAIL.n199 B 0.022743f
C239 VTAIL.n200 B 0.010188f
C240 VTAIL.n201 B 0.017906f
C241 VTAIL.n202 B 0.009622f
C242 VTAIL.n203 B 0.022743f
C243 VTAIL.n204 B 0.010188f
C244 VTAIL.n205 B 0.653715f
C245 VTAIL.n206 B 0.009622f
C246 VTAIL.t6 B 0.037125f
C247 VTAIL.n207 B 0.088835f
C248 VTAIL.n208 B 0.013435f
C249 VTAIL.n209 B 0.017057f
C250 VTAIL.n210 B 0.022743f
C251 VTAIL.n211 B 0.010188f
C252 VTAIL.n212 B 0.009622f
C253 VTAIL.n213 B 0.017906f
C254 VTAIL.n214 B 0.017906f
C255 VTAIL.n215 B 0.009622f
C256 VTAIL.n216 B 0.010188f
C257 VTAIL.n217 B 0.022743f
C258 VTAIL.n218 B 0.022743f
C259 VTAIL.n219 B 0.010188f
C260 VTAIL.n220 B 0.009622f
C261 VTAIL.n221 B 0.017906f
C262 VTAIL.n222 B 0.017906f
C263 VTAIL.n223 B 0.009622f
C264 VTAIL.n224 B 0.010188f
C265 VTAIL.n225 B 0.022743f
C266 VTAIL.n226 B 0.022743f
C267 VTAIL.n227 B 0.010188f
C268 VTAIL.n228 B 0.009622f
C269 VTAIL.n229 B 0.017906f
C270 VTAIL.n230 B 0.017906f
C271 VTAIL.n231 B 0.009622f
C272 VTAIL.n232 B 0.010188f
C273 VTAIL.n233 B 0.022743f
C274 VTAIL.n234 B 0.050303f
C275 VTAIL.n235 B 0.010188f
C276 VTAIL.n236 B 0.009622f
C277 VTAIL.n237 B 0.038698f
C278 VTAIL.n238 B 0.028171f
C279 VTAIL.n239 B 0.069734f
C280 VTAIL.n240 B 0.025773f
C281 VTAIL.n241 B 0.017906f
C282 VTAIL.n242 B 0.009622f
C283 VTAIL.n243 B 0.022743f
C284 VTAIL.n244 B 0.010188f
C285 VTAIL.n245 B 0.017906f
C286 VTAIL.n246 B 0.009622f
C287 VTAIL.n247 B 0.022743f
C288 VTAIL.n248 B 0.010188f
C289 VTAIL.n249 B 0.017906f
C290 VTAIL.n250 B 0.009622f
C291 VTAIL.n251 B 0.022743f
C292 VTAIL.n252 B 0.010188f
C293 VTAIL.n253 B 0.653715f
C294 VTAIL.n254 B 0.009622f
C295 VTAIL.t0 B 0.037125f
C296 VTAIL.n255 B 0.088835f
C297 VTAIL.n256 B 0.013435f
C298 VTAIL.n257 B 0.017057f
C299 VTAIL.n258 B 0.022743f
C300 VTAIL.n259 B 0.010188f
C301 VTAIL.n260 B 0.009622f
C302 VTAIL.n261 B 0.017906f
C303 VTAIL.n262 B 0.017906f
C304 VTAIL.n263 B 0.009622f
C305 VTAIL.n264 B 0.010188f
C306 VTAIL.n265 B 0.022743f
C307 VTAIL.n266 B 0.022743f
C308 VTAIL.n267 B 0.010188f
C309 VTAIL.n268 B 0.009622f
C310 VTAIL.n269 B 0.017906f
C311 VTAIL.n270 B 0.017906f
C312 VTAIL.n271 B 0.009622f
C313 VTAIL.n272 B 0.010188f
C314 VTAIL.n273 B 0.022743f
C315 VTAIL.n274 B 0.022743f
C316 VTAIL.n275 B 0.010188f
C317 VTAIL.n276 B 0.009622f
C318 VTAIL.n277 B 0.017906f
C319 VTAIL.n278 B 0.017906f
C320 VTAIL.n279 B 0.009622f
C321 VTAIL.n280 B 0.010188f
C322 VTAIL.n281 B 0.022743f
C323 VTAIL.n282 B 0.050303f
C324 VTAIL.n283 B 0.010188f
C325 VTAIL.n284 B 0.009622f
C326 VTAIL.n285 B 0.038698f
C327 VTAIL.n286 B 0.028171f
C328 VTAIL.n287 B 0.069734f
C329 VTAIL.n288 B 0.025773f
C330 VTAIL.n289 B 0.017906f
C331 VTAIL.n290 B 0.009622f
C332 VTAIL.n291 B 0.022743f
C333 VTAIL.n292 B 0.010188f
C334 VTAIL.n293 B 0.017906f
C335 VTAIL.n294 B 0.009622f
C336 VTAIL.n295 B 0.022743f
C337 VTAIL.n296 B 0.010188f
C338 VTAIL.n297 B 0.017906f
C339 VTAIL.n298 B 0.009622f
C340 VTAIL.n299 B 0.022743f
C341 VTAIL.n300 B 0.010188f
C342 VTAIL.n301 B 0.653715f
C343 VTAIL.n302 B 0.009622f
C344 VTAIL.t3 B 0.037125f
C345 VTAIL.n303 B 0.088835f
C346 VTAIL.n304 B 0.013435f
C347 VTAIL.n305 B 0.017057f
C348 VTAIL.n306 B 0.022743f
C349 VTAIL.n307 B 0.010188f
C350 VTAIL.n308 B 0.009622f
C351 VTAIL.n309 B 0.017906f
C352 VTAIL.n310 B 0.017906f
C353 VTAIL.n311 B 0.009622f
C354 VTAIL.n312 B 0.010188f
C355 VTAIL.n313 B 0.022743f
C356 VTAIL.n314 B 0.022743f
C357 VTAIL.n315 B 0.010188f
C358 VTAIL.n316 B 0.009622f
C359 VTAIL.n317 B 0.017906f
C360 VTAIL.n318 B 0.017906f
C361 VTAIL.n319 B 0.009622f
C362 VTAIL.n320 B 0.010188f
C363 VTAIL.n321 B 0.022743f
C364 VTAIL.n322 B 0.022743f
C365 VTAIL.n323 B 0.010188f
C366 VTAIL.n324 B 0.009622f
C367 VTAIL.n325 B 0.017906f
C368 VTAIL.n326 B 0.017906f
C369 VTAIL.n327 B 0.009622f
C370 VTAIL.n328 B 0.010188f
C371 VTAIL.n329 B 0.022743f
C372 VTAIL.n330 B 0.050303f
C373 VTAIL.n331 B 0.010188f
C374 VTAIL.n332 B 0.009622f
C375 VTAIL.n333 B 0.038698f
C376 VTAIL.n334 B 0.028171f
C377 VTAIL.n335 B 0.751917f
C378 VTAIL.n336 B 0.025773f
C379 VTAIL.n337 B 0.017906f
C380 VTAIL.n338 B 0.009622f
C381 VTAIL.n339 B 0.022743f
C382 VTAIL.n340 B 0.010188f
C383 VTAIL.n341 B 0.017906f
C384 VTAIL.n342 B 0.009622f
C385 VTAIL.n343 B 0.022743f
C386 VTAIL.n344 B 0.010188f
C387 VTAIL.n345 B 0.017906f
C388 VTAIL.n346 B 0.009622f
C389 VTAIL.n347 B 0.022743f
C390 VTAIL.n348 B 0.010188f
C391 VTAIL.n349 B 0.653715f
C392 VTAIL.n350 B 0.009622f
C393 VTAIL.t7 B 0.037125f
C394 VTAIL.n351 B 0.088835f
C395 VTAIL.n352 B 0.013435f
C396 VTAIL.n353 B 0.017057f
C397 VTAIL.n354 B 0.022743f
C398 VTAIL.n355 B 0.010188f
C399 VTAIL.n356 B 0.009622f
C400 VTAIL.n357 B 0.017906f
C401 VTAIL.n358 B 0.017906f
C402 VTAIL.n359 B 0.009622f
C403 VTAIL.n360 B 0.010188f
C404 VTAIL.n361 B 0.022743f
C405 VTAIL.n362 B 0.022743f
C406 VTAIL.n363 B 0.010188f
C407 VTAIL.n364 B 0.009622f
C408 VTAIL.n365 B 0.017906f
C409 VTAIL.n366 B 0.017906f
C410 VTAIL.n367 B 0.009622f
C411 VTAIL.n368 B 0.010188f
C412 VTAIL.n369 B 0.022743f
C413 VTAIL.n370 B 0.022743f
C414 VTAIL.n371 B 0.010188f
C415 VTAIL.n372 B 0.009622f
C416 VTAIL.n373 B 0.017906f
C417 VTAIL.n374 B 0.017906f
C418 VTAIL.n375 B 0.009622f
C419 VTAIL.n376 B 0.010188f
C420 VTAIL.n377 B 0.022743f
C421 VTAIL.n378 B 0.050303f
C422 VTAIL.n379 B 0.010188f
C423 VTAIL.n380 B 0.009622f
C424 VTAIL.n381 B 0.038698f
C425 VTAIL.n382 B 0.028171f
C426 VTAIL.n383 B 0.734135f
C427 VN.t1 B 0.236906f
C428 VN.t3 B 0.236906f
C429 VN.n0 B 0.20703f
C430 VN.t2 B 0.236906f
C431 VN.t0 B 0.236906f
C432 VN.n1 B 0.440247f
.ends

