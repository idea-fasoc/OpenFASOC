* NGSPICE file created from diff_pair_sample_0275.ext - technology: sky130A

.subckt diff_pair_sample_0275 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=0 ps=0 w=13.12 l=2.79
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=5.1168 ps=27.02 w=13.12 l=2.79
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=5.1168 ps=27.02 w=13.12 l=2.79
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=0 ps=0 w=13.12 l=2.79
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=5.1168 ps=27.02 w=13.12 l=2.79
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=0 ps=0 w=13.12 l=2.79
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=5.1168 ps=27.02 w=13.12 l=2.79
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1168 pd=27.02 as=0 ps=0 w=13.12 l=2.79
R0 B.n523 B.n106 585
R1 B.n106 B.n51 585
R2 B.n525 B.n524 585
R3 B.n527 B.n105 585
R4 B.n530 B.n529 585
R5 B.n531 B.n104 585
R6 B.n533 B.n532 585
R7 B.n535 B.n103 585
R8 B.n538 B.n537 585
R9 B.n539 B.n102 585
R10 B.n541 B.n540 585
R11 B.n543 B.n101 585
R12 B.n546 B.n545 585
R13 B.n547 B.n100 585
R14 B.n549 B.n548 585
R15 B.n551 B.n99 585
R16 B.n554 B.n553 585
R17 B.n555 B.n98 585
R18 B.n557 B.n556 585
R19 B.n559 B.n97 585
R20 B.n562 B.n561 585
R21 B.n563 B.n96 585
R22 B.n565 B.n564 585
R23 B.n567 B.n95 585
R24 B.n570 B.n569 585
R25 B.n571 B.n94 585
R26 B.n573 B.n572 585
R27 B.n575 B.n93 585
R28 B.n578 B.n577 585
R29 B.n579 B.n92 585
R30 B.n581 B.n580 585
R31 B.n583 B.n91 585
R32 B.n586 B.n585 585
R33 B.n587 B.n90 585
R34 B.n589 B.n588 585
R35 B.n591 B.n89 585
R36 B.n594 B.n593 585
R37 B.n595 B.n88 585
R38 B.n597 B.n596 585
R39 B.n599 B.n87 585
R40 B.n602 B.n601 585
R41 B.n603 B.n86 585
R42 B.n605 B.n604 585
R43 B.n607 B.n85 585
R44 B.n609 B.n608 585
R45 B.n611 B.n610 585
R46 B.n614 B.n613 585
R47 B.n615 B.n80 585
R48 B.n617 B.n616 585
R49 B.n619 B.n79 585
R50 B.n622 B.n621 585
R51 B.n623 B.n78 585
R52 B.n625 B.n624 585
R53 B.n627 B.n77 585
R54 B.n630 B.n629 585
R55 B.n632 B.n74 585
R56 B.n634 B.n633 585
R57 B.n636 B.n73 585
R58 B.n639 B.n638 585
R59 B.n640 B.n72 585
R60 B.n642 B.n641 585
R61 B.n644 B.n71 585
R62 B.n647 B.n646 585
R63 B.n648 B.n70 585
R64 B.n650 B.n649 585
R65 B.n652 B.n69 585
R66 B.n655 B.n654 585
R67 B.n656 B.n68 585
R68 B.n658 B.n657 585
R69 B.n660 B.n67 585
R70 B.n663 B.n662 585
R71 B.n664 B.n66 585
R72 B.n666 B.n665 585
R73 B.n668 B.n65 585
R74 B.n671 B.n670 585
R75 B.n672 B.n64 585
R76 B.n674 B.n673 585
R77 B.n676 B.n63 585
R78 B.n679 B.n678 585
R79 B.n680 B.n62 585
R80 B.n682 B.n681 585
R81 B.n684 B.n61 585
R82 B.n687 B.n686 585
R83 B.n688 B.n60 585
R84 B.n690 B.n689 585
R85 B.n692 B.n59 585
R86 B.n695 B.n694 585
R87 B.n696 B.n58 585
R88 B.n698 B.n697 585
R89 B.n700 B.n57 585
R90 B.n703 B.n702 585
R91 B.n704 B.n56 585
R92 B.n706 B.n705 585
R93 B.n708 B.n55 585
R94 B.n711 B.n710 585
R95 B.n712 B.n54 585
R96 B.n714 B.n713 585
R97 B.n716 B.n53 585
R98 B.n719 B.n718 585
R99 B.n720 B.n52 585
R100 B.n522 B.n50 585
R101 B.n723 B.n50 585
R102 B.n521 B.n49 585
R103 B.n724 B.n49 585
R104 B.n520 B.n48 585
R105 B.n725 B.n48 585
R106 B.n519 B.n518 585
R107 B.n518 B.n44 585
R108 B.n517 B.n43 585
R109 B.n731 B.n43 585
R110 B.n516 B.n42 585
R111 B.n732 B.n42 585
R112 B.n515 B.n41 585
R113 B.n733 B.n41 585
R114 B.n514 B.n513 585
R115 B.n513 B.n40 585
R116 B.n512 B.n36 585
R117 B.n739 B.n36 585
R118 B.n511 B.n35 585
R119 B.n740 B.n35 585
R120 B.n510 B.n34 585
R121 B.n741 B.n34 585
R122 B.n509 B.n508 585
R123 B.n508 B.n30 585
R124 B.n507 B.n29 585
R125 B.n747 B.n29 585
R126 B.n506 B.n28 585
R127 B.n748 B.n28 585
R128 B.n505 B.n27 585
R129 B.n749 B.n27 585
R130 B.n504 B.n503 585
R131 B.n503 B.n23 585
R132 B.n502 B.n22 585
R133 B.n755 B.n22 585
R134 B.n501 B.n21 585
R135 B.n756 B.n21 585
R136 B.n500 B.n20 585
R137 B.n757 B.n20 585
R138 B.n499 B.n498 585
R139 B.n498 B.n16 585
R140 B.n497 B.n15 585
R141 B.n763 B.n15 585
R142 B.n496 B.n14 585
R143 B.n764 B.n14 585
R144 B.n495 B.n13 585
R145 B.n765 B.n13 585
R146 B.n494 B.n493 585
R147 B.n493 B.n12 585
R148 B.n492 B.n491 585
R149 B.n492 B.n8 585
R150 B.n490 B.n7 585
R151 B.n772 B.n7 585
R152 B.n489 B.n6 585
R153 B.n773 B.n6 585
R154 B.n488 B.n5 585
R155 B.n774 B.n5 585
R156 B.n487 B.n486 585
R157 B.n486 B.n4 585
R158 B.n485 B.n107 585
R159 B.n485 B.n484 585
R160 B.n475 B.n108 585
R161 B.n109 B.n108 585
R162 B.n477 B.n476 585
R163 B.n478 B.n477 585
R164 B.n474 B.n114 585
R165 B.n114 B.n113 585
R166 B.n473 B.n472 585
R167 B.n472 B.n471 585
R168 B.n116 B.n115 585
R169 B.n117 B.n116 585
R170 B.n464 B.n463 585
R171 B.n465 B.n464 585
R172 B.n462 B.n122 585
R173 B.n122 B.n121 585
R174 B.n461 B.n460 585
R175 B.n460 B.n459 585
R176 B.n124 B.n123 585
R177 B.n125 B.n124 585
R178 B.n452 B.n451 585
R179 B.n453 B.n452 585
R180 B.n450 B.n130 585
R181 B.n130 B.n129 585
R182 B.n449 B.n448 585
R183 B.n448 B.n447 585
R184 B.n132 B.n131 585
R185 B.n133 B.n132 585
R186 B.n440 B.n439 585
R187 B.n441 B.n440 585
R188 B.n438 B.n138 585
R189 B.n138 B.n137 585
R190 B.n437 B.n436 585
R191 B.n436 B.n435 585
R192 B.n140 B.n139 585
R193 B.n428 B.n140 585
R194 B.n427 B.n426 585
R195 B.n429 B.n427 585
R196 B.n425 B.n145 585
R197 B.n145 B.n144 585
R198 B.n424 B.n423 585
R199 B.n423 B.n422 585
R200 B.n147 B.n146 585
R201 B.n148 B.n147 585
R202 B.n415 B.n414 585
R203 B.n416 B.n415 585
R204 B.n413 B.n153 585
R205 B.n153 B.n152 585
R206 B.n412 B.n411 585
R207 B.n411 B.n410 585
R208 B.n407 B.n157 585
R209 B.n406 B.n405 585
R210 B.n403 B.n158 585
R211 B.n403 B.n156 585
R212 B.n402 B.n401 585
R213 B.n400 B.n399 585
R214 B.n398 B.n160 585
R215 B.n396 B.n395 585
R216 B.n394 B.n161 585
R217 B.n393 B.n392 585
R218 B.n390 B.n162 585
R219 B.n388 B.n387 585
R220 B.n386 B.n163 585
R221 B.n385 B.n384 585
R222 B.n382 B.n164 585
R223 B.n380 B.n379 585
R224 B.n378 B.n165 585
R225 B.n377 B.n376 585
R226 B.n374 B.n166 585
R227 B.n372 B.n371 585
R228 B.n370 B.n167 585
R229 B.n369 B.n368 585
R230 B.n366 B.n168 585
R231 B.n364 B.n363 585
R232 B.n362 B.n169 585
R233 B.n361 B.n360 585
R234 B.n358 B.n170 585
R235 B.n356 B.n355 585
R236 B.n354 B.n171 585
R237 B.n353 B.n352 585
R238 B.n350 B.n172 585
R239 B.n348 B.n347 585
R240 B.n346 B.n173 585
R241 B.n345 B.n344 585
R242 B.n342 B.n174 585
R243 B.n340 B.n339 585
R244 B.n338 B.n175 585
R245 B.n337 B.n336 585
R246 B.n334 B.n176 585
R247 B.n332 B.n331 585
R248 B.n330 B.n177 585
R249 B.n329 B.n328 585
R250 B.n326 B.n178 585
R251 B.n324 B.n323 585
R252 B.n322 B.n179 585
R253 B.n321 B.n320 585
R254 B.n318 B.n317 585
R255 B.n316 B.n315 585
R256 B.n314 B.n184 585
R257 B.n312 B.n311 585
R258 B.n310 B.n185 585
R259 B.n309 B.n308 585
R260 B.n306 B.n186 585
R261 B.n304 B.n303 585
R262 B.n302 B.n187 585
R263 B.n300 B.n299 585
R264 B.n297 B.n190 585
R265 B.n295 B.n294 585
R266 B.n293 B.n191 585
R267 B.n292 B.n291 585
R268 B.n289 B.n192 585
R269 B.n287 B.n286 585
R270 B.n285 B.n193 585
R271 B.n284 B.n283 585
R272 B.n281 B.n194 585
R273 B.n279 B.n278 585
R274 B.n277 B.n195 585
R275 B.n276 B.n275 585
R276 B.n273 B.n196 585
R277 B.n271 B.n270 585
R278 B.n269 B.n197 585
R279 B.n268 B.n267 585
R280 B.n265 B.n198 585
R281 B.n263 B.n262 585
R282 B.n261 B.n199 585
R283 B.n260 B.n259 585
R284 B.n257 B.n200 585
R285 B.n255 B.n254 585
R286 B.n253 B.n201 585
R287 B.n252 B.n251 585
R288 B.n249 B.n202 585
R289 B.n247 B.n246 585
R290 B.n245 B.n203 585
R291 B.n244 B.n243 585
R292 B.n241 B.n204 585
R293 B.n239 B.n238 585
R294 B.n237 B.n205 585
R295 B.n236 B.n235 585
R296 B.n233 B.n206 585
R297 B.n231 B.n230 585
R298 B.n229 B.n207 585
R299 B.n228 B.n227 585
R300 B.n225 B.n208 585
R301 B.n223 B.n222 585
R302 B.n221 B.n209 585
R303 B.n220 B.n219 585
R304 B.n217 B.n210 585
R305 B.n215 B.n214 585
R306 B.n213 B.n212 585
R307 B.n155 B.n154 585
R308 B.n409 B.n408 585
R309 B.n410 B.n409 585
R310 B.n151 B.n150 585
R311 B.n152 B.n151 585
R312 B.n418 B.n417 585
R313 B.n417 B.n416 585
R314 B.n419 B.n149 585
R315 B.n149 B.n148 585
R316 B.n421 B.n420 585
R317 B.n422 B.n421 585
R318 B.n143 B.n142 585
R319 B.n144 B.n143 585
R320 B.n431 B.n430 585
R321 B.n430 B.n429 585
R322 B.n432 B.n141 585
R323 B.n428 B.n141 585
R324 B.n434 B.n433 585
R325 B.n435 B.n434 585
R326 B.n136 B.n135 585
R327 B.n137 B.n136 585
R328 B.n443 B.n442 585
R329 B.n442 B.n441 585
R330 B.n444 B.n134 585
R331 B.n134 B.n133 585
R332 B.n446 B.n445 585
R333 B.n447 B.n446 585
R334 B.n128 B.n127 585
R335 B.n129 B.n128 585
R336 B.n455 B.n454 585
R337 B.n454 B.n453 585
R338 B.n456 B.n126 585
R339 B.n126 B.n125 585
R340 B.n458 B.n457 585
R341 B.n459 B.n458 585
R342 B.n120 B.n119 585
R343 B.n121 B.n120 585
R344 B.n467 B.n466 585
R345 B.n466 B.n465 585
R346 B.n468 B.n118 585
R347 B.n118 B.n117 585
R348 B.n470 B.n469 585
R349 B.n471 B.n470 585
R350 B.n112 B.n111 585
R351 B.n113 B.n112 585
R352 B.n480 B.n479 585
R353 B.n479 B.n478 585
R354 B.n481 B.n110 585
R355 B.n110 B.n109 585
R356 B.n483 B.n482 585
R357 B.n484 B.n483 585
R358 B.n3 B.n0 585
R359 B.n4 B.n3 585
R360 B.n771 B.n1 585
R361 B.n772 B.n771 585
R362 B.n770 B.n769 585
R363 B.n770 B.n8 585
R364 B.n768 B.n9 585
R365 B.n12 B.n9 585
R366 B.n767 B.n766 585
R367 B.n766 B.n765 585
R368 B.n11 B.n10 585
R369 B.n764 B.n11 585
R370 B.n762 B.n761 585
R371 B.n763 B.n762 585
R372 B.n760 B.n17 585
R373 B.n17 B.n16 585
R374 B.n759 B.n758 585
R375 B.n758 B.n757 585
R376 B.n19 B.n18 585
R377 B.n756 B.n19 585
R378 B.n754 B.n753 585
R379 B.n755 B.n754 585
R380 B.n752 B.n24 585
R381 B.n24 B.n23 585
R382 B.n751 B.n750 585
R383 B.n750 B.n749 585
R384 B.n26 B.n25 585
R385 B.n748 B.n26 585
R386 B.n746 B.n745 585
R387 B.n747 B.n746 585
R388 B.n744 B.n31 585
R389 B.n31 B.n30 585
R390 B.n743 B.n742 585
R391 B.n742 B.n741 585
R392 B.n33 B.n32 585
R393 B.n740 B.n33 585
R394 B.n738 B.n737 585
R395 B.n739 B.n738 585
R396 B.n736 B.n37 585
R397 B.n40 B.n37 585
R398 B.n735 B.n734 585
R399 B.n734 B.n733 585
R400 B.n39 B.n38 585
R401 B.n732 B.n39 585
R402 B.n730 B.n729 585
R403 B.n731 B.n730 585
R404 B.n728 B.n45 585
R405 B.n45 B.n44 585
R406 B.n727 B.n726 585
R407 B.n726 B.n725 585
R408 B.n47 B.n46 585
R409 B.n724 B.n47 585
R410 B.n722 B.n721 585
R411 B.n723 B.n722 585
R412 B.n775 B.n774 585
R413 B.n773 B.n2 585
R414 B.n722 B.n52 526.135
R415 B.n106 B.n50 526.135
R416 B.n411 B.n155 526.135
R417 B.n409 B.n157 526.135
R418 B.n75 B.t9 321.647
R419 B.n81 B.t13 321.647
R420 B.n188 B.t2 321.647
R421 B.n180 B.t6 321.647
R422 B.n526 B.n51 256.663
R423 B.n528 B.n51 256.663
R424 B.n534 B.n51 256.663
R425 B.n536 B.n51 256.663
R426 B.n542 B.n51 256.663
R427 B.n544 B.n51 256.663
R428 B.n550 B.n51 256.663
R429 B.n552 B.n51 256.663
R430 B.n558 B.n51 256.663
R431 B.n560 B.n51 256.663
R432 B.n566 B.n51 256.663
R433 B.n568 B.n51 256.663
R434 B.n574 B.n51 256.663
R435 B.n576 B.n51 256.663
R436 B.n582 B.n51 256.663
R437 B.n584 B.n51 256.663
R438 B.n590 B.n51 256.663
R439 B.n592 B.n51 256.663
R440 B.n598 B.n51 256.663
R441 B.n600 B.n51 256.663
R442 B.n606 B.n51 256.663
R443 B.n84 B.n51 256.663
R444 B.n612 B.n51 256.663
R445 B.n618 B.n51 256.663
R446 B.n620 B.n51 256.663
R447 B.n626 B.n51 256.663
R448 B.n628 B.n51 256.663
R449 B.n635 B.n51 256.663
R450 B.n637 B.n51 256.663
R451 B.n643 B.n51 256.663
R452 B.n645 B.n51 256.663
R453 B.n651 B.n51 256.663
R454 B.n653 B.n51 256.663
R455 B.n659 B.n51 256.663
R456 B.n661 B.n51 256.663
R457 B.n667 B.n51 256.663
R458 B.n669 B.n51 256.663
R459 B.n675 B.n51 256.663
R460 B.n677 B.n51 256.663
R461 B.n683 B.n51 256.663
R462 B.n685 B.n51 256.663
R463 B.n691 B.n51 256.663
R464 B.n693 B.n51 256.663
R465 B.n699 B.n51 256.663
R466 B.n701 B.n51 256.663
R467 B.n707 B.n51 256.663
R468 B.n709 B.n51 256.663
R469 B.n715 B.n51 256.663
R470 B.n717 B.n51 256.663
R471 B.n404 B.n156 256.663
R472 B.n159 B.n156 256.663
R473 B.n397 B.n156 256.663
R474 B.n391 B.n156 256.663
R475 B.n389 B.n156 256.663
R476 B.n383 B.n156 256.663
R477 B.n381 B.n156 256.663
R478 B.n375 B.n156 256.663
R479 B.n373 B.n156 256.663
R480 B.n367 B.n156 256.663
R481 B.n365 B.n156 256.663
R482 B.n359 B.n156 256.663
R483 B.n357 B.n156 256.663
R484 B.n351 B.n156 256.663
R485 B.n349 B.n156 256.663
R486 B.n343 B.n156 256.663
R487 B.n341 B.n156 256.663
R488 B.n335 B.n156 256.663
R489 B.n333 B.n156 256.663
R490 B.n327 B.n156 256.663
R491 B.n325 B.n156 256.663
R492 B.n319 B.n156 256.663
R493 B.n183 B.n156 256.663
R494 B.n313 B.n156 256.663
R495 B.n307 B.n156 256.663
R496 B.n305 B.n156 256.663
R497 B.n298 B.n156 256.663
R498 B.n296 B.n156 256.663
R499 B.n290 B.n156 256.663
R500 B.n288 B.n156 256.663
R501 B.n282 B.n156 256.663
R502 B.n280 B.n156 256.663
R503 B.n274 B.n156 256.663
R504 B.n272 B.n156 256.663
R505 B.n266 B.n156 256.663
R506 B.n264 B.n156 256.663
R507 B.n258 B.n156 256.663
R508 B.n256 B.n156 256.663
R509 B.n250 B.n156 256.663
R510 B.n248 B.n156 256.663
R511 B.n242 B.n156 256.663
R512 B.n240 B.n156 256.663
R513 B.n234 B.n156 256.663
R514 B.n232 B.n156 256.663
R515 B.n226 B.n156 256.663
R516 B.n224 B.n156 256.663
R517 B.n218 B.n156 256.663
R518 B.n216 B.n156 256.663
R519 B.n211 B.n156 256.663
R520 B.n777 B.n776 256.663
R521 B.n718 B.n716 163.367
R522 B.n714 B.n54 163.367
R523 B.n710 B.n708 163.367
R524 B.n706 B.n56 163.367
R525 B.n702 B.n700 163.367
R526 B.n698 B.n58 163.367
R527 B.n694 B.n692 163.367
R528 B.n690 B.n60 163.367
R529 B.n686 B.n684 163.367
R530 B.n682 B.n62 163.367
R531 B.n678 B.n676 163.367
R532 B.n674 B.n64 163.367
R533 B.n670 B.n668 163.367
R534 B.n666 B.n66 163.367
R535 B.n662 B.n660 163.367
R536 B.n658 B.n68 163.367
R537 B.n654 B.n652 163.367
R538 B.n650 B.n70 163.367
R539 B.n646 B.n644 163.367
R540 B.n642 B.n72 163.367
R541 B.n638 B.n636 163.367
R542 B.n634 B.n74 163.367
R543 B.n629 B.n627 163.367
R544 B.n625 B.n78 163.367
R545 B.n621 B.n619 163.367
R546 B.n617 B.n80 163.367
R547 B.n613 B.n611 163.367
R548 B.n608 B.n607 163.367
R549 B.n605 B.n86 163.367
R550 B.n601 B.n599 163.367
R551 B.n597 B.n88 163.367
R552 B.n593 B.n591 163.367
R553 B.n589 B.n90 163.367
R554 B.n585 B.n583 163.367
R555 B.n581 B.n92 163.367
R556 B.n577 B.n575 163.367
R557 B.n573 B.n94 163.367
R558 B.n569 B.n567 163.367
R559 B.n565 B.n96 163.367
R560 B.n561 B.n559 163.367
R561 B.n557 B.n98 163.367
R562 B.n553 B.n551 163.367
R563 B.n549 B.n100 163.367
R564 B.n545 B.n543 163.367
R565 B.n541 B.n102 163.367
R566 B.n537 B.n535 163.367
R567 B.n533 B.n104 163.367
R568 B.n529 B.n527 163.367
R569 B.n525 B.n106 163.367
R570 B.n411 B.n153 163.367
R571 B.n415 B.n153 163.367
R572 B.n415 B.n147 163.367
R573 B.n423 B.n147 163.367
R574 B.n423 B.n145 163.367
R575 B.n427 B.n145 163.367
R576 B.n427 B.n140 163.367
R577 B.n436 B.n140 163.367
R578 B.n436 B.n138 163.367
R579 B.n440 B.n138 163.367
R580 B.n440 B.n132 163.367
R581 B.n448 B.n132 163.367
R582 B.n448 B.n130 163.367
R583 B.n452 B.n130 163.367
R584 B.n452 B.n124 163.367
R585 B.n460 B.n124 163.367
R586 B.n460 B.n122 163.367
R587 B.n464 B.n122 163.367
R588 B.n464 B.n116 163.367
R589 B.n472 B.n116 163.367
R590 B.n472 B.n114 163.367
R591 B.n477 B.n114 163.367
R592 B.n477 B.n108 163.367
R593 B.n485 B.n108 163.367
R594 B.n486 B.n485 163.367
R595 B.n486 B.n5 163.367
R596 B.n6 B.n5 163.367
R597 B.n7 B.n6 163.367
R598 B.n492 B.n7 163.367
R599 B.n493 B.n492 163.367
R600 B.n493 B.n13 163.367
R601 B.n14 B.n13 163.367
R602 B.n15 B.n14 163.367
R603 B.n498 B.n15 163.367
R604 B.n498 B.n20 163.367
R605 B.n21 B.n20 163.367
R606 B.n22 B.n21 163.367
R607 B.n503 B.n22 163.367
R608 B.n503 B.n27 163.367
R609 B.n28 B.n27 163.367
R610 B.n29 B.n28 163.367
R611 B.n508 B.n29 163.367
R612 B.n508 B.n34 163.367
R613 B.n35 B.n34 163.367
R614 B.n36 B.n35 163.367
R615 B.n513 B.n36 163.367
R616 B.n513 B.n41 163.367
R617 B.n42 B.n41 163.367
R618 B.n43 B.n42 163.367
R619 B.n518 B.n43 163.367
R620 B.n518 B.n48 163.367
R621 B.n49 B.n48 163.367
R622 B.n50 B.n49 163.367
R623 B.n405 B.n403 163.367
R624 B.n403 B.n402 163.367
R625 B.n399 B.n398 163.367
R626 B.n396 B.n161 163.367
R627 B.n392 B.n390 163.367
R628 B.n388 B.n163 163.367
R629 B.n384 B.n382 163.367
R630 B.n380 B.n165 163.367
R631 B.n376 B.n374 163.367
R632 B.n372 B.n167 163.367
R633 B.n368 B.n366 163.367
R634 B.n364 B.n169 163.367
R635 B.n360 B.n358 163.367
R636 B.n356 B.n171 163.367
R637 B.n352 B.n350 163.367
R638 B.n348 B.n173 163.367
R639 B.n344 B.n342 163.367
R640 B.n340 B.n175 163.367
R641 B.n336 B.n334 163.367
R642 B.n332 B.n177 163.367
R643 B.n328 B.n326 163.367
R644 B.n324 B.n179 163.367
R645 B.n320 B.n318 163.367
R646 B.n315 B.n314 163.367
R647 B.n312 B.n185 163.367
R648 B.n308 B.n306 163.367
R649 B.n304 B.n187 163.367
R650 B.n299 B.n297 163.367
R651 B.n295 B.n191 163.367
R652 B.n291 B.n289 163.367
R653 B.n287 B.n193 163.367
R654 B.n283 B.n281 163.367
R655 B.n279 B.n195 163.367
R656 B.n275 B.n273 163.367
R657 B.n271 B.n197 163.367
R658 B.n267 B.n265 163.367
R659 B.n263 B.n199 163.367
R660 B.n259 B.n257 163.367
R661 B.n255 B.n201 163.367
R662 B.n251 B.n249 163.367
R663 B.n247 B.n203 163.367
R664 B.n243 B.n241 163.367
R665 B.n239 B.n205 163.367
R666 B.n235 B.n233 163.367
R667 B.n231 B.n207 163.367
R668 B.n227 B.n225 163.367
R669 B.n223 B.n209 163.367
R670 B.n219 B.n217 163.367
R671 B.n215 B.n212 163.367
R672 B.n409 B.n151 163.367
R673 B.n417 B.n151 163.367
R674 B.n417 B.n149 163.367
R675 B.n421 B.n149 163.367
R676 B.n421 B.n143 163.367
R677 B.n430 B.n143 163.367
R678 B.n430 B.n141 163.367
R679 B.n434 B.n141 163.367
R680 B.n434 B.n136 163.367
R681 B.n442 B.n136 163.367
R682 B.n442 B.n134 163.367
R683 B.n446 B.n134 163.367
R684 B.n446 B.n128 163.367
R685 B.n454 B.n128 163.367
R686 B.n454 B.n126 163.367
R687 B.n458 B.n126 163.367
R688 B.n458 B.n120 163.367
R689 B.n466 B.n120 163.367
R690 B.n466 B.n118 163.367
R691 B.n470 B.n118 163.367
R692 B.n470 B.n112 163.367
R693 B.n479 B.n112 163.367
R694 B.n479 B.n110 163.367
R695 B.n483 B.n110 163.367
R696 B.n483 B.n3 163.367
R697 B.n775 B.n3 163.367
R698 B.n771 B.n2 163.367
R699 B.n771 B.n770 163.367
R700 B.n770 B.n9 163.367
R701 B.n766 B.n9 163.367
R702 B.n766 B.n11 163.367
R703 B.n762 B.n11 163.367
R704 B.n762 B.n17 163.367
R705 B.n758 B.n17 163.367
R706 B.n758 B.n19 163.367
R707 B.n754 B.n19 163.367
R708 B.n754 B.n24 163.367
R709 B.n750 B.n24 163.367
R710 B.n750 B.n26 163.367
R711 B.n746 B.n26 163.367
R712 B.n746 B.n31 163.367
R713 B.n742 B.n31 163.367
R714 B.n742 B.n33 163.367
R715 B.n738 B.n33 163.367
R716 B.n738 B.n37 163.367
R717 B.n734 B.n37 163.367
R718 B.n734 B.n39 163.367
R719 B.n730 B.n39 163.367
R720 B.n730 B.n45 163.367
R721 B.n726 B.n45 163.367
R722 B.n726 B.n47 163.367
R723 B.n722 B.n47 163.367
R724 B.n81 B.t14 132.038
R725 B.n188 B.t5 132.038
R726 B.n75 B.t11 132.022
R727 B.n180 B.t8 132.022
R728 B.n410 B.n156 72.3571
R729 B.n723 B.n51 72.3571
R730 B.n717 B.n52 71.676
R731 B.n716 B.n715 71.676
R732 B.n709 B.n54 71.676
R733 B.n708 B.n707 71.676
R734 B.n701 B.n56 71.676
R735 B.n700 B.n699 71.676
R736 B.n693 B.n58 71.676
R737 B.n692 B.n691 71.676
R738 B.n685 B.n60 71.676
R739 B.n684 B.n683 71.676
R740 B.n677 B.n62 71.676
R741 B.n676 B.n675 71.676
R742 B.n669 B.n64 71.676
R743 B.n668 B.n667 71.676
R744 B.n661 B.n66 71.676
R745 B.n660 B.n659 71.676
R746 B.n653 B.n68 71.676
R747 B.n652 B.n651 71.676
R748 B.n645 B.n70 71.676
R749 B.n644 B.n643 71.676
R750 B.n637 B.n72 71.676
R751 B.n636 B.n635 71.676
R752 B.n628 B.n74 71.676
R753 B.n627 B.n626 71.676
R754 B.n620 B.n78 71.676
R755 B.n619 B.n618 71.676
R756 B.n612 B.n80 71.676
R757 B.n611 B.n84 71.676
R758 B.n607 B.n606 71.676
R759 B.n600 B.n86 71.676
R760 B.n599 B.n598 71.676
R761 B.n592 B.n88 71.676
R762 B.n591 B.n590 71.676
R763 B.n584 B.n90 71.676
R764 B.n583 B.n582 71.676
R765 B.n576 B.n92 71.676
R766 B.n575 B.n574 71.676
R767 B.n568 B.n94 71.676
R768 B.n567 B.n566 71.676
R769 B.n560 B.n96 71.676
R770 B.n559 B.n558 71.676
R771 B.n552 B.n98 71.676
R772 B.n551 B.n550 71.676
R773 B.n544 B.n100 71.676
R774 B.n543 B.n542 71.676
R775 B.n536 B.n102 71.676
R776 B.n535 B.n534 71.676
R777 B.n528 B.n104 71.676
R778 B.n527 B.n526 71.676
R779 B.n526 B.n525 71.676
R780 B.n529 B.n528 71.676
R781 B.n534 B.n533 71.676
R782 B.n537 B.n536 71.676
R783 B.n542 B.n541 71.676
R784 B.n545 B.n544 71.676
R785 B.n550 B.n549 71.676
R786 B.n553 B.n552 71.676
R787 B.n558 B.n557 71.676
R788 B.n561 B.n560 71.676
R789 B.n566 B.n565 71.676
R790 B.n569 B.n568 71.676
R791 B.n574 B.n573 71.676
R792 B.n577 B.n576 71.676
R793 B.n582 B.n581 71.676
R794 B.n585 B.n584 71.676
R795 B.n590 B.n589 71.676
R796 B.n593 B.n592 71.676
R797 B.n598 B.n597 71.676
R798 B.n601 B.n600 71.676
R799 B.n606 B.n605 71.676
R800 B.n608 B.n84 71.676
R801 B.n613 B.n612 71.676
R802 B.n618 B.n617 71.676
R803 B.n621 B.n620 71.676
R804 B.n626 B.n625 71.676
R805 B.n629 B.n628 71.676
R806 B.n635 B.n634 71.676
R807 B.n638 B.n637 71.676
R808 B.n643 B.n642 71.676
R809 B.n646 B.n645 71.676
R810 B.n651 B.n650 71.676
R811 B.n654 B.n653 71.676
R812 B.n659 B.n658 71.676
R813 B.n662 B.n661 71.676
R814 B.n667 B.n666 71.676
R815 B.n670 B.n669 71.676
R816 B.n675 B.n674 71.676
R817 B.n678 B.n677 71.676
R818 B.n683 B.n682 71.676
R819 B.n686 B.n685 71.676
R820 B.n691 B.n690 71.676
R821 B.n694 B.n693 71.676
R822 B.n699 B.n698 71.676
R823 B.n702 B.n701 71.676
R824 B.n707 B.n706 71.676
R825 B.n710 B.n709 71.676
R826 B.n715 B.n714 71.676
R827 B.n718 B.n717 71.676
R828 B.n404 B.n157 71.676
R829 B.n402 B.n159 71.676
R830 B.n398 B.n397 71.676
R831 B.n391 B.n161 71.676
R832 B.n390 B.n389 71.676
R833 B.n383 B.n163 71.676
R834 B.n382 B.n381 71.676
R835 B.n375 B.n165 71.676
R836 B.n374 B.n373 71.676
R837 B.n367 B.n167 71.676
R838 B.n366 B.n365 71.676
R839 B.n359 B.n169 71.676
R840 B.n358 B.n357 71.676
R841 B.n351 B.n171 71.676
R842 B.n350 B.n349 71.676
R843 B.n343 B.n173 71.676
R844 B.n342 B.n341 71.676
R845 B.n335 B.n175 71.676
R846 B.n334 B.n333 71.676
R847 B.n327 B.n177 71.676
R848 B.n326 B.n325 71.676
R849 B.n319 B.n179 71.676
R850 B.n318 B.n183 71.676
R851 B.n314 B.n313 71.676
R852 B.n307 B.n185 71.676
R853 B.n306 B.n305 71.676
R854 B.n298 B.n187 71.676
R855 B.n297 B.n296 71.676
R856 B.n290 B.n191 71.676
R857 B.n289 B.n288 71.676
R858 B.n282 B.n193 71.676
R859 B.n281 B.n280 71.676
R860 B.n274 B.n195 71.676
R861 B.n273 B.n272 71.676
R862 B.n266 B.n197 71.676
R863 B.n265 B.n264 71.676
R864 B.n258 B.n199 71.676
R865 B.n257 B.n256 71.676
R866 B.n250 B.n201 71.676
R867 B.n249 B.n248 71.676
R868 B.n242 B.n203 71.676
R869 B.n241 B.n240 71.676
R870 B.n234 B.n205 71.676
R871 B.n233 B.n232 71.676
R872 B.n226 B.n207 71.676
R873 B.n225 B.n224 71.676
R874 B.n218 B.n209 71.676
R875 B.n217 B.n216 71.676
R876 B.n212 B.n211 71.676
R877 B.n405 B.n404 71.676
R878 B.n399 B.n159 71.676
R879 B.n397 B.n396 71.676
R880 B.n392 B.n391 71.676
R881 B.n389 B.n388 71.676
R882 B.n384 B.n383 71.676
R883 B.n381 B.n380 71.676
R884 B.n376 B.n375 71.676
R885 B.n373 B.n372 71.676
R886 B.n368 B.n367 71.676
R887 B.n365 B.n364 71.676
R888 B.n360 B.n359 71.676
R889 B.n357 B.n356 71.676
R890 B.n352 B.n351 71.676
R891 B.n349 B.n348 71.676
R892 B.n344 B.n343 71.676
R893 B.n341 B.n340 71.676
R894 B.n336 B.n335 71.676
R895 B.n333 B.n332 71.676
R896 B.n328 B.n327 71.676
R897 B.n325 B.n324 71.676
R898 B.n320 B.n319 71.676
R899 B.n315 B.n183 71.676
R900 B.n313 B.n312 71.676
R901 B.n308 B.n307 71.676
R902 B.n305 B.n304 71.676
R903 B.n299 B.n298 71.676
R904 B.n296 B.n295 71.676
R905 B.n291 B.n290 71.676
R906 B.n288 B.n287 71.676
R907 B.n283 B.n282 71.676
R908 B.n280 B.n279 71.676
R909 B.n275 B.n274 71.676
R910 B.n272 B.n271 71.676
R911 B.n267 B.n266 71.676
R912 B.n264 B.n263 71.676
R913 B.n259 B.n258 71.676
R914 B.n256 B.n255 71.676
R915 B.n251 B.n250 71.676
R916 B.n248 B.n247 71.676
R917 B.n243 B.n242 71.676
R918 B.n240 B.n239 71.676
R919 B.n235 B.n234 71.676
R920 B.n232 B.n231 71.676
R921 B.n227 B.n226 71.676
R922 B.n224 B.n223 71.676
R923 B.n219 B.n218 71.676
R924 B.n216 B.n215 71.676
R925 B.n211 B.n155 71.676
R926 B.n776 B.n775 71.676
R927 B.n776 B.n2 71.676
R928 B.n82 B.t15 71.5293
R929 B.n189 B.t4 71.5293
R930 B.n76 B.t12 71.5126
R931 B.n181 B.t7 71.5126
R932 B.n76 B.n75 60.5096
R933 B.n82 B.n81 60.5096
R934 B.n189 B.n188 60.5096
R935 B.n181 B.n180 60.5096
R936 B.n631 B.n76 59.5399
R937 B.n83 B.n82 59.5399
R938 B.n301 B.n189 59.5399
R939 B.n182 B.n181 59.5399
R940 B.n410 B.n152 40.6637
R941 B.n416 B.n152 40.6637
R942 B.n416 B.n148 40.6637
R943 B.n422 B.n148 40.6637
R944 B.n422 B.n144 40.6637
R945 B.n429 B.n144 40.6637
R946 B.n429 B.n428 40.6637
R947 B.n435 B.n137 40.6637
R948 B.n441 B.n137 40.6637
R949 B.n441 B.n133 40.6637
R950 B.n447 B.n133 40.6637
R951 B.n447 B.n129 40.6637
R952 B.n453 B.n129 40.6637
R953 B.n453 B.n125 40.6637
R954 B.n459 B.n125 40.6637
R955 B.n459 B.n121 40.6637
R956 B.n465 B.n121 40.6637
R957 B.n465 B.n117 40.6637
R958 B.n471 B.n117 40.6637
R959 B.n478 B.n113 40.6637
R960 B.n478 B.n109 40.6637
R961 B.n484 B.n109 40.6637
R962 B.n484 B.n4 40.6637
R963 B.n774 B.n4 40.6637
R964 B.n774 B.n773 40.6637
R965 B.n773 B.n772 40.6637
R966 B.n772 B.n8 40.6637
R967 B.n12 B.n8 40.6637
R968 B.n765 B.n12 40.6637
R969 B.n765 B.n764 40.6637
R970 B.n763 B.n16 40.6637
R971 B.n757 B.n16 40.6637
R972 B.n757 B.n756 40.6637
R973 B.n756 B.n755 40.6637
R974 B.n755 B.n23 40.6637
R975 B.n749 B.n23 40.6637
R976 B.n749 B.n748 40.6637
R977 B.n748 B.n747 40.6637
R978 B.n747 B.n30 40.6637
R979 B.n741 B.n30 40.6637
R980 B.n741 B.n740 40.6637
R981 B.n740 B.n739 40.6637
R982 B.n733 B.n40 40.6637
R983 B.n733 B.n732 40.6637
R984 B.n732 B.n731 40.6637
R985 B.n731 B.n44 40.6637
R986 B.n725 B.n44 40.6637
R987 B.n725 B.n724 40.6637
R988 B.n724 B.n723 40.6637
R989 B.n428 B.t3 37.6738
R990 B.n40 B.t10 37.6738
R991 B.n408 B.n407 34.1859
R992 B.n412 B.n154 34.1859
R993 B.n523 B.n522 34.1859
R994 B.n721 B.n720 34.1859
R995 B.t0 B.n113 28.106
R996 B.n764 B.t1 28.106
R997 B B.n777 18.0485
R998 B.n471 B.t0 12.5583
R999 B.t1 B.n763 12.5583
R1000 B.n408 B.n150 10.6151
R1001 B.n418 B.n150 10.6151
R1002 B.n419 B.n418 10.6151
R1003 B.n420 B.n419 10.6151
R1004 B.n420 B.n142 10.6151
R1005 B.n431 B.n142 10.6151
R1006 B.n432 B.n431 10.6151
R1007 B.n433 B.n432 10.6151
R1008 B.n433 B.n135 10.6151
R1009 B.n443 B.n135 10.6151
R1010 B.n444 B.n443 10.6151
R1011 B.n445 B.n444 10.6151
R1012 B.n445 B.n127 10.6151
R1013 B.n455 B.n127 10.6151
R1014 B.n456 B.n455 10.6151
R1015 B.n457 B.n456 10.6151
R1016 B.n457 B.n119 10.6151
R1017 B.n467 B.n119 10.6151
R1018 B.n468 B.n467 10.6151
R1019 B.n469 B.n468 10.6151
R1020 B.n469 B.n111 10.6151
R1021 B.n480 B.n111 10.6151
R1022 B.n481 B.n480 10.6151
R1023 B.n482 B.n481 10.6151
R1024 B.n482 B.n0 10.6151
R1025 B.n407 B.n406 10.6151
R1026 B.n406 B.n158 10.6151
R1027 B.n401 B.n158 10.6151
R1028 B.n401 B.n400 10.6151
R1029 B.n400 B.n160 10.6151
R1030 B.n395 B.n160 10.6151
R1031 B.n395 B.n394 10.6151
R1032 B.n394 B.n393 10.6151
R1033 B.n393 B.n162 10.6151
R1034 B.n387 B.n162 10.6151
R1035 B.n387 B.n386 10.6151
R1036 B.n386 B.n385 10.6151
R1037 B.n385 B.n164 10.6151
R1038 B.n379 B.n164 10.6151
R1039 B.n379 B.n378 10.6151
R1040 B.n378 B.n377 10.6151
R1041 B.n377 B.n166 10.6151
R1042 B.n371 B.n166 10.6151
R1043 B.n371 B.n370 10.6151
R1044 B.n370 B.n369 10.6151
R1045 B.n369 B.n168 10.6151
R1046 B.n363 B.n168 10.6151
R1047 B.n363 B.n362 10.6151
R1048 B.n362 B.n361 10.6151
R1049 B.n361 B.n170 10.6151
R1050 B.n355 B.n170 10.6151
R1051 B.n355 B.n354 10.6151
R1052 B.n354 B.n353 10.6151
R1053 B.n353 B.n172 10.6151
R1054 B.n347 B.n172 10.6151
R1055 B.n347 B.n346 10.6151
R1056 B.n346 B.n345 10.6151
R1057 B.n345 B.n174 10.6151
R1058 B.n339 B.n174 10.6151
R1059 B.n339 B.n338 10.6151
R1060 B.n338 B.n337 10.6151
R1061 B.n337 B.n176 10.6151
R1062 B.n331 B.n176 10.6151
R1063 B.n331 B.n330 10.6151
R1064 B.n330 B.n329 10.6151
R1065 B.n329 B.n178 10.6151
R1066 B.n323 B.n178 10.6151
R1067 B.n323 B.n322 10.6151
R1068 B.n322 B.n321 10.6151
R1069 B.n317 B.n316 10.6151
R1070 B.n316 B.n184 10.6151
R1071 B.n311 B.n184 10.6151
R1072 B.n311 B.n310 10.6151
R1073 B.n310 B.n309 10.6151
R1074 B.n309 B.n186 10.6151
R1075 B.n303 B.n186 10.6151
R1076 B.n303 B.n302 10.6151
R1077 B.n300 B.n190 10.6151
R1078 B.n294 B.n190 10.6151
R1079 B.n294 B.n293 10.6151
R1080 B.n293 B.n292 10.6151
R1081 B.n292 B.n192 10.6151
R1082 B.n286 B.n192 10.6151
R1083 B.n286 B.n285 10.6151
R1084 B.n285 B.n284 10.6151
R1085 B.n284 B.n194 10.6151
R1086 B.n278 B.n194 10.6151
R1087 B.n278 B.n277 10.6151
R1088 B.n277 B.n276 10.6151
R1089 B.n276 B.n196 10.6151
R1090 B.n270 B.n196 10.6151
R1091 B.n270 B.n269 10.6151
R1092 B.n269 B.n268 10.6151
R1093 B.n268 B.n198 10.6151
R1094 B.n262 B.n198 10.6151
R1095 B.n262 B.n261 10.6151
R1096 B.n261 B.n260 10.6151
R1097 B.n260 B.n200 10.6151
R1098 B.n254 B.n200 10.6151
R1099 B.n254 B.n253 10.6151
R1100 B.n253 B.n252 10.6151
R1101 B.n252 B.n202 10.6151
R1102 B.n246 B.n202 10.6151
R1103 B.n246 B.n245 10.6151
R1104 B.n245 B.n244 10.6151
R1105 B.n244 B.n204 10.6151
R1106 B.n238 B.n204 10.6151
R1107 B.n238 B.n237 10.6151
R1108 B.n237 B.n236 10.6151
R1109 B.n236 B.n206 10.6151
R1110 B.n230 B.n206 10.6151
R1111 B.n230 B.n229 10.6151
R1112 B.n229 B.n228 10.6151
R1113 B.n228 B.n208 10.6151
R1114 B.n222 B.n208 10.6151
R1115 B.n222 B.n221 10.6151
R1116 B.n221 B.n220 10.6151
R1117 B.n220 B.n210 10.6151
R1118 B.n214 B.n210 10.6151
R1119 B.n214 B.n213 10.6151
R1120 B.n213 B.n154 10.6151
R1121 B.n413 B.n412 10.6151
R1122 B.n414 B.n413 10.6151
R1123 B.n414 B.n146 10.6151
R1124 B.n424 B.n146 10.6151
R1125 B.n425 B.n424 10.6151
R1126 B.n426 B.n425 10.6151
R1127 B.n426 B.n139 10.6151
R1128 B.n437 B.n139 10.6151
R1129 B.n438 B.n437 10.6151
R1130 B.n439 B.n438 10.6151
R1131 B.n439 B.n131 10.6151
R1132 B.n449 B.n131 10.6151
R1133 B.n450 B.n449 10.6151
R1134 B.n451 B.n450 10.6151
R1135 B.n451 B.n123 10.6151
R1136 B.n461 B.n123 10.6151
R1137 B.n462 B.n461 10.6151
R1138 B.n463 B.n462 10.6151
R1139 B.n463 B.n115 10.6151
R1140 B.n473 B.n115 10.6151
R1141 B.n474 B.n473 10.6151
R1142 B.n476 B.n474 10.6151
R1143 B.n476 B.n475 10.6151
R1144 B.n475 B.n107 10.6151
R1145 B.n487 B.n107 10.6151
R1146 B.n488 B.n487 10.6151
R1147 B.n489 B.n488 10.6151
R1148 B.n490 B.n489 10.6151
R1149 B.n491 B.n490 10.6151
R1150 B.n494 B.n491 10.6151
R1151 B.n495 B.n494 10.6151
R1152 B.n496 B.n495 10.6151
R1153 B.n497 B.n496 10.6151
R1154 B.n499 B.n497 10.6151
R1155 B.n500 B.n499 10.6151
R1156 B.n501 B.n500 10.6151
R1157 B.n502 B.n501 10.6151
R1158 B.n504 B.n502 10.6151
R1159 B.n505 B.n504 10.6151
R1160 B.n506 B.n505 10.6151
R1161 B.n507 B.n506 10.6151
R1162 B.n509 B.n507 10.6151
R1163 B.n510 B.n509 10.6151
R1164 B.n511 B.n510 10.6151
R1165 B.n512 B.n511 10.6151
R1166 B.n514 B.n512 10.6151
R1167 B.n515 B.n514 10.6151
R1168 B.n516 B.n515 10.6151
R1169 B.n517 B.n516 10.6151
R1170 B.n519 B.n517 10.6151
R1171 B.n520 B.n519 10.6151
R1172 B.n521 B.n520 10.6151
R1173 B.n522 B.n521 10.6151
R1174 B.n769 B.n1 10.6151
R1175 B.n769 B.n768 10.6151
R1176 B.n768 B.n767 10.6151
R1177 B.n767 B.n10 10.6151
R1178 B.n761 B.n10 10.6151
R1179 B.n761 B.n760 10.6151
R1180 B.n760 B.n759 10.6151
R1181 B.n759 B.n18 10.6151
R1182 B.n753 B.n18 10.6151
R1183 B.n753 B.n752 10.6151
R1184 B.n752 B.n751 10.6151
R1185 B.n751 B.n25 10.6151
R1186 B.n745 B.n25 10.6151
R1187 B.n745 B.n744 10.6151
R1188 B.n744 B.n743 10.6151
R1189 B.n743 B.n32 10.6151
R1190 B.n737 B.n32 10.6151
R1191 B.n737 B.n736 10.6151
R1192 B.n736 B.n735 10.6151
R1193 B.n735 B.n38 10.6151
R1194 B.n729 B.n38 10.6151
R1195 B.n729 B.n728 10.6151
R1196 B.n728 B.n727 10.6151
R1197 B.n727 B.n46 10.6151
R1198 B.n721 B.n46 10.6151
R1199 B.n720 B.n719 10.6151
R1200 B.n719 B.n53 10.6151
R1201 B.n713 B.n53 10.6151
R1202 B.n713 B.n712 10.6151
R1203 B.n712 B.n711 10.6151
R1204 B.n711 B.n55 10.6151
R1205 B.n705 B.n55 10.6151
R1206 B.n705 B.n704 10.6151
R1207 B.n704 B.n703 10.6151
R1208 B.n703 B.n57 10.6151
R1209 B.n697 B.n57 10.6151
R1210 B.n697 B.n696 10.6151
R1211 B.n696 B.n695 10.6151
R1212 B.n695 B.n59 10.6151
R1213 B.n689 B.n59 10.6151
R1214 B.n689 B.n688 10.6151
R1215 B.n688 B.n687 10.6151
R1216 B.n687 B.n61 10.6151
R1217 B.n681 B.n61 10.6151
R1218 B.n681 B.n680 10.6151
R1219 B.n680 B.n679 10.6151
R1220 B.n679 B.n63 10.6151
R1221 B.n673 B.n63 10.6151
R1222 B.n673 B.n672 10.6151
R1223 B.n672 B.n671 10.6151
R1224 B.n671 B.n65 10.6151
R1225 B.n665 B.n65 10.6151
R1226 B.n665 B.n664 10.6151
R1227 B.n664 B.n663 10.6151
R1228 B.n663 B.n67 10.6151
R1229 B.n657 B.n67 10.6151
R1230 B.n657 B.n656 10.6151
R1231 B.n656 B.n655 10.6151
R1232 B.n655 B.n69 10.6151
R1233 B.n649 B.n69 10.6151
R1234 B.n649 B.n648 10.6151
R1235 B.n648 B.n647 10.6151
R1236 B.n647 B.n71 10.6151
R1237 B.n641 B.n71 10.6151
R1238 B.n641 B.n640 10.6151
R1239 B.n640 B.n639 10.6151
R1240 B.n639 B.n73 10.6151
R1241 B.n633 B.n73 10.6151
R1242 B.n633 B.n632 10.6151
R1243 B.n630 B.n77 10.6151
R1244 B.n624 B.n77 10.6151
R1245 B.n624 B.n623 10.6151
R1246 B.n623 B.n622 10.6151
R1247 B.n622 B.n79 10.6151
R1248 B.n616 B.n79 10.6151
R1249 B.n616 B.n615 10.6151
R1250 B.n615 B.n614 10.6151
R1251 B.n610 B.n609 10.6151
R1252 B.n609 B.n85 10.6151
R1253 B.n604 B.n85 10.6151
R1254 B.n604 B.n603 10.6151
R1255 B.n603 B.n602 10.6151
R1256 B.n602 B.n87 10.6151
R1257 B.n596 B.n87 10.6151
R1258 B.n596 B.n595 10.6151
R1259 B.n595 B.n594 10.6151
R1260 B.n594 B.n89 10.6151
R1261 B.n588 B.n89 10.6151
R1262 B.n588 B.n587 10.6151
R1263 B.n587 B.n586 10.6151
R1264 B.n586 B.n91 10.6151
R1265 B.n580 B.n91 10.6151
R1266 B.n580 B.n579 10.6151
R1267 B.n579 B.n578 10.6151
R1268 B.n578 B.n93 10.6151
R1269 B.n572 B.n93 10.6151
R1270 B.n572 B.n571 10.6151
R1271 B.n571 B.n570 10.6151
R1272 B.n570 B.n95 10.6151
R1273 B.n564 B.n95 10.6151
R1274 B.n564 B.n563 10.6151
R1275 B.n563 B.n562 10.6151
R1276 B.n562 B.n97 10.6151
R1277 B.n556 B.n97 10.6151
R1278 B.n556 B.n555 10.6151
R1279 B.n555 B.n554 10.6151
R1280 B.n554 B.n99 10.6151
R1281 B.n548 B.n99 10.6151
R1282 B.n548 B.n547 10.6151
R1283 B.n547 B.n546 10.6151
R1284 B.n546 B.n101 10.6151
R1285 B.n540 B.n101 10.6151
R1286 B.n540 B.n539 10.6151
R1287 B.n539 B.n538 10.6151
R1288 B.n538 B.n103 10.6151
R1289 B.n532 B.n103 10.6151
R1290 B.n532 B.n531 10.6151
R1291 B.n531 B.n530 10.6151
R1292 B.n530 B.n105 10.6151
R1293 B.n524 B.n105 10.6151
R1294 B.n524 B.n523 10.6151
R1295 B.n777 B.n0 8.11757
R1296 B.n777 B.n1 8.11757
R1297 B.n317 B.n182 6.5566
R1298 B.n302 B.n301 6.5566
R1299 B.n631 B.n630 6.5566
R1300 B.n614 B.n83 6.5566
R1301 B.n321 B.n182 4.05904
R1302 B.n301 B.n300 4.05904
R1303 B.n632 B.n631 4.05904
R1304 B.n610 B.n83 4.05904
R1305 B.n435 B.t3 2.99044
R1306 B.n739 B.t10 2.99044
R1307 VP.n0 VP.t1 200.477
R1308 VP.n0 VP.t0 154.469
R1309 VP VP.n0 0.431812
R1310 VTAIL.n1 VTAIL.t1 44.9041
R1311 VTAIL.n3 VTAIL.t0 44.9039
R1312 VTAIL.n0 VTAIL.t2 44.9039
R1313 VTAIL.n2 VTAIL.t3 44.9039
R1314 VTAIL.n1 VTAIL.n0 29.0565
R1315 VTAIL.n3 VTAIL.n2 26.3669
R1316 VTAIL.n2 VTAIL.n1 1.81516
R1317 VTAIL VTAIL.n0 1.20093
R1318 VTAIL VTAIL.n3 0.614724
R1319 VDD1 VDD1.t1 103.129
R1320 VDD1 VDD1.t0 62.3133
R1321 VN VN.t1 200.48
R1322 VN VN.t0 154.9
R1323 VDD2.n0 VDD2.t1 101.931
R1324 VDD2.n0 VDD2.t0 61.5827
R1325 VDD2 VDD2.n0 0.731103
C0 VTAIL VDD1 5.38773f
C1 VP VDD1 3.23827f
C2 VN VDD2 3.04798f
C3 VTAIL VN 2.68033f
C4 VP VN 5.75089f
C5 VTAIL VDD2 5.43957f
C6 VP VDD2 0.341462f
C7 VN VDD1 0.148543f
C8 VP VTAIL 2.69461f
C9 VDD1 VDD2 0.697696f
C10 VDD2 B 4.696283f
C11 VDD1 B 7.92792f
C12 VTAIL B 7.901886f
C13 VN B 11.176901f
C14 VP B 6.717873f
C15 VDD2.t1 B 2.95481f
C16 VDD2.t0 B 2.36625f
C17 VDD2.n0 B 2.94467f
C18 VN.t0 B 3.25894f
C19 VN.t1 B 3.82266f
C20 VDD1.t0 B 2.40478f
C21 VDD1.t1 B 3.03782f
C22 VTAIL.t2 B 2.34949f
C23 VTAIL.n0 B 1.74891f
C24 VTAIL.t1 B 2.3495f
C25 VTAIL.n1 B 1.7896f
C26 VTAIL.t3 B 2.34949f
C27 VTAIL.n2 B 1.61142f
C28 VTAIL.t0 B 2.34949f
C29 VTAIL.n3 B 1.53189f
C30 VP.t0 B 3.32454f
C31 VP.t1 B 3.90144f
C32 VP.n0 B 4.39154f
.ends

