* NGSPICE file created from diff_pair_sample_1184.ext - technology: sky130A

.subckt diff_pair_sample_1184 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=3.2736 ps=20.17 w=19.84 l=0.7
X1 VDD1.t8 VP.t1 VTAIL.t14 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=7.7376 ps=40.46 w=19.84 l=0.7
X2 VTAIL.t3 VN.t0 VDD2.t9 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X3 VDD2.t8 VN.t1 VTAIL.t5 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X4 VTAIL.t17 VP.t2 VDD1.t7 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X5 B.t11 B.t9 B.t10 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=0 ps=0 w=19.84 l=0.7
X6 B.t8 B.t6 B.t7 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=0 ps=0 w=19.84 l=0.7
X7 VDD2.t7 VN.t2 VTAIL.t0 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=7.7376 ps=40.46 w=19.84 l=0.7
X8 VDD2.t6 VN.t3 VTAIL.t4 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=3.2736 ps=20.17 w=19.84 l=0.7
X9 B.t5 B.t3 B.t4 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=0 ps=0 w=19.84 l=0.7
X10 VDD2.t5 VN.t4 VTAIL.t7 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=3.2736 ps=20.17 w=19.84 l=0.7
X11 VDD2.t4 VN.t5 VTAIL.t1 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X12 VTAIL.t6 VN.t6 VDD2.t3 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X13 VTAIL.t13 VP.t3 VDD1.t6 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X14 VDD2.t2 VN.t7 VTAIL.t9 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=7.7376 ps=40.46 w=19.84 l=0.7
X15 VTAIL.t18 VP.t4 VDD1.t5 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X16 VTAIL.t11 VP.t5 VDD1.t4 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X17 VDD1.t3 VP.t6 VTAIL.t16 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=3.2736 ps=20.17 w=19.84 l=0.7
X18 VTAIL.t2 VN.t8 VDD2.t1 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X19 VDD1.t2 VP.t7 VTAIL.t19 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X20 VDD1.t1 VP.t8 VTAIL.t10 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X21 VTAIL.t8 VN.t9 VDD2.t0 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=3.2736 ps=20.17 w=19.84 l=0.7
X22 B.t2 B.t0 B.t1 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=7.7376 pd=40.46 as=0 ps=0 w=19.84 l=0.7
X23 VDD1.t0 VP.t9 VTAIL.t15 w_n2206_n4936# sky130_fd_pr__pfet_01v8 ad=3.2736 pd=20.17 as=7.7376 ps=40.46 w=19.84 l=0.7
R0 VP.n7 VP.t0 761.929
R1 VP.n18 VP.t6 739.182
R2 VP.n22 VP.t5 739.182
R3 VP.n24 VP.t7 739.182
R4 VP.n28 VP.t2 739.182
R5 VP.n30 VP.t1 739.182
R6 VP.n16 VP.t9 739.182
R7 VP.n14 VP.t3 739.182
R8 VP.n6 VP.t8 739.182
R9 VP.n8 VP.t4 739.182
R10 VP.n31 VP.n30 161.3
R11 VP.n10 VP.n9 161.3
R12 VP.n11 VP.n6 161.3
R13 VP.n13 VP.n12 161.3
R14 VP.n14 VP.n5 161.3
R15 VP.n15 VP.n4 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n29 VP.n0 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.n1 161.3
R20 VP.n25 VP.n24 161.3
R21 VP.n23 VP.n2 161.3
R22 VP.n22 VP.n21 161.3
R23 VP.n20 VP.n3 161.3
R24 VP.n19 VP.n18 161.3
R25 VP.n19 VP.n17 48.724
R26 VP.n10 VP.n7 44.8741
R27 VP.n18 VP.n3 30.6732
R28 VP.n30 VP.n29 30.6732
R29 VP.n16 VP.n15 30.6732
R30 VP.n23 VP.n22 26.2914
R31 VP.n28 VP.n1 26.2914
R32 VP.n14 VP.n13 26.2914
R33 VP.n9 VP.n8 26.2914
R34 VP.n24 VP.n23 21.9096
R35 VP.n24 VP.n1 21.9096
R36 VP.n13 VP.n6 21.9096
R37 VP.n9 VP.n6 21.9096
R38 VP.n8 VP.n7 19.0667
R39 VP.n22 VP.n3 17.5278
R40 VP.n29 VP.n28 17.5278
R41 VP.n15 VP.n14 17.5278
R42 VP.n11 VP.n10 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n5 0.189894
R45 VP.n5 VP.n4 0.189894
R46 VP.n17 VP.n4 0.189894
R47 VP.n20 VP.n19 0.189894
R48 VP.n21 VP.n20 0.189894
R49 VP.n21 VP.n2 0.189894
R50 VP.n25 VP.n2 0.189894
R51 VP.n26 VP.n25 0.189894
R52 VP.n27 VP.n26 0.189894
R53 VP.n27 VP.n0 0.189894
R54 VP.n31 VP.n0 0.189894
R55 VP VP.n31 0.0516364
R56 VTAIL.n11 VTAIL.t9 55.7848
R57 VTAIL.n17 VTAIL.t0 55.7846
R58 VTAIL.n2 VTAIL.t14 55.7846
R59 VTAIL.n16 VTAIL.t15 55.7846
R60 VTAIL.n15 VTAIL.n14 54.1464
R61 VTAIL.n13 VTAIL.n12 54.1464
R62 VTAIL.n10 VTAIL.n9 54.1464
R63 VTAIL.n8 VTAIL.n7 54.1464
R64 VTAIL.n19 VTAIL.n18 54.1462
R65 VTAIL.n1 VTAIL.n0 54.1462
R66 VTAIL.n4 VTAIL.n3 54.1462
R67 VTAIL.n6 VTAIL.n5 54.1462
R68 VTAIL.n8 VTAIL.n6 31.2462
R69 VTAIL.n17 VTAIL.n16 30.3583
R70 VTAIL.n18 VTAIL.t5 1.63886
R71 VTAIL.n18 VTAIL.t3 1.63886
R72 VTAIL.n0 VTAIL.t7 1.63886
R73 VTAIL.n0 VTAIL.t6 1.63886
R74 VTAIL.n3 VTAIL.t19 1.63886
R75 VTAIL.n3 VTAIL.t17 1.63886
R76 VTAIL.n5 VTAIL.t16 1.63886
R77 VTAIL.n5 VTAIL.t11 1.63886
R78 VTAIL.n14 VTAIL.t10 1.63886
R79 VTAIL.n14 VTAIL.t13 1.63886
R80 VTAIL.n12 VTAIL.t12 1.63886
R81 VTAIL.n12 VTAIL.t18 1.63886
R82 VTAIL.n9 VTAIL.t1 1.63886
R83 VTAIL.n9 VTAIL.t8 1.63886
R84 VTAIL.n7 VTAIL.t4 1.63886
R85 VTAIL.n7 VTAIL.t2 1.63886
R86 VTAIL.n13 VTAIL.n11 0.914293
R87 VTAIL.n2 VTAIL.n1 0.914293
R88 VTAIL.n10 VTAIL.n8 0.888431
R89 VTAIL.n11 VTAIL.n10 0.888431
R90 VTAIL.n15 VTAIL.n13 0.888431
R91 VTAIL.n16 VTAIL.n15 0.888431
R92 VTAIL.n6 VTAIL.n4 0.888431
R93 VTAIL.n4 VTAIL.n2 0.888431
R94 VTAIL.n19 VTAIL.n17 0.888431
R95 VTAIL VTAIL.n1 0.724638
R96 VTAIL VTAIL.n19 0.164293
R97 VDD1.n1 VDD1.t9 73.3515
R98 VDD1.n3 VDD1.t3 73.3513
R99 VDD1.n5 VDD1.n4 71.4356
R100 VDD1.n1 VDD1.n0 70.8252
R101 VDD1.n7 VDD1.n6 70.8251
R102 VDD1.n3 VDD1.n2 70.825
R103 VDD1.n7 VDD1.n5 46.0634
R104 VDD1.n6 VDD1.t6 1.63886
R105 VDD1.n6 VDD1.t0 1.63886
R106 VDD1.n0 VDD1.t5 1.63886
R107 VDD1.n0 VDD1.t1 1.63886
R108 VDD1.n4 VDD1.t7 1.63886
R109 VDD1.n4 VDD1.t8 1.63886
R110 VDD1.n2 VDD1.t4 1.63886
R111 VDD1.n2 VDD1.t2 1.63886
R112 VDD1 VDD1.n7 0.608259
R113 VDD1 VDD1.n1 0.280672
R114 VDD1.n5 VDD1.n3 0.167137
R115 VN.n3 VN.t4 761.929
R116 VN.n17 VN.t7 761.929
R117 VN.n4 VN.t6 739.182
R118 VN.n6 VN.t1 739.182
R119 VN.n10 VN.t0 739.182
R120 VN.n12 VN.t2 739.182
R121 VN.n18 VN.t9 739.182
R122 VN.n20 VN.t5 739.182
R123 VN.n24 VN.t8 739.182
R124 VN.n26 VN.t3 739.182
R125 VN.n13 VN.n12 161.3
R126 VN.n27 VN.n26 161.3
R127 VN.n25 VN.n14 161.3
R128 VN.n24 VN.n23 161.3
R129 VN.n22 VN.n15 161.3
R130 VN.n21 VN.n20 161.3
R131 VN.n19 VN.n16 161.3
R132 VN.n11 VN.n0 161.3
R133 VN.n10 VN.n9 161.3
R134 VN.n8 VN.n1 161.3
R135 VN.n7 VN.n6 161.3
R136 VN.n5 VN.n2 161.3
R137 VN VN.n27 49.1047
R138 VN.n17 VN.n16 44.8741
R139 VN.n3 VN.n2 44.8741
R140 VN.n12 VN.n11 30.6732
R141 VN.n26 VN.n25 30.6732
R142 VN.n5 VN.n4 26.2914
R143 VN.n10 VN.n1 26.2914
R144 VN.n19 VN.n18 26.2914
R145 VN.n24 VN.n15 26.2914
R146 VN.n6 VN.n5 21.9096
R147 VN.n6 VN.n1 21.9096
R148 VN.n20 VN.n19 21.9096
R149 VN.n20 VN.n15 21.9096
R150 VN.n4 VN.n3 19.0667
R151 VN.n18 VN.n17 19.0667
R152 VN.n11 VN.n10 17.5278
R153 VN.n25 VN.n24 17.5278
R154 VN.n27 VN.n14 0.189894
R155 VN.n23 VN.n14 0.189894
R156 VN.n23 VN.n22 0.189894
R157 VN.n22 VN.n21 0.189894
R158 VN.n21 VN.n16 0.189894
R159 VN.n7 VN.n2 0.189894
R160 VN.n8 VN.n7 0.189894
R161 VN.n9 VN.n8 0.189894
R162 VN.n9 VN.n0 0.189894
R163 VN.n13 VN.n0 0.189894
R164 VN VN.n13 0.0516364
R165 VDD2.n1 VDD2.t5 73.3513
R166 VDD2.n4 VDD2.t6 72.4636
R167 VDD2.n3 VDD2.n2 71.4356
R168 VDD2 VDD2.n7 71.4328
R169 VDD2.n6 VDD2.n5 70.8252
R170 VDD2.n1 VDD2.n0 70.825
R171 VDD2.n4 VDD2.n3 45.0364
R172 VDD2.n7 VDD2.t0 1.63886
R173 VDD2.n7 VDD2.t2 1.63886
R174 VDD2.n5 VDD2.t1 1.63886
R175 VDD2.n5 VDD2.t4 1.63886
R176 VDD2.n2 VDD2.t9 1.63886
R177 VDD2.n2 VDD2.t7 1.63886
R178 VDD2.n0 VDD2.t3 1.63886
R179 VDD2.n0 VDD2.t8 1.63886
R180 VDD2.n6 VDD2.n4 0.888431
R181 VDD2 VDD2.n6 0.280672
R182 VDD2.n3 VDD2.n1 0.167137
R183 B.n148 B.t6 886.029
R184 B.n156 B.t3 886.029
R185 B.n48 B.t0 886.029
R186 B.n54 B.t9 886.029
R187 B.n530 B.n529 585
R188 B.n531 B.n88 585
R189 B.n533 B.n532 585
R190 B.n534 B.n87 585
R191 B.n536 B.n535 585
R192 B.n537 B.n86 585
R193 B.n539 B.n538 585
R194 B.n540 B.n85 585
R195 B.n542 B.n541 585
R196 B.n543 B.n84 585
R197 B.n545 B.n544 585
R198 B.n546 B.n83 585
R199 B.n548 B.n547 585
R200 B.n549 B.n82 585
R201 B.n551 B.n550 585
R202 B.n552 B.n81 585
R203 B.n554 B.n553 585
R204 B.n555 B.n80 585
R205 B.n557 B.n556 585
R206 B.n558 B.n79 585
R207 B.n560 B.n559 585
R208 B.n561 B.n78 585
R209 B.n563 B.n562 585
R210 B.n564 B.n77 585
R211 B.n566 B.n565 585
R212 B.n567 B.n76 585
R213 B.n569 B.n568 585
R214 B.n570 B.n75 585
R215 B.n572 B.n571 585
R216 B.n573 B.n74 585
R217 B.n575 B.n574 585
R218 B.n576 B.n73 585
R219 B.n578 B.n577 585
R220 B.n579 B.n72 585
R221 B.n581 B.n580 585
R222 B.n582 B.n71 585
R223 B.n584 B.n583 585
R224 B.n585 B.n70 585
R225 B.n587 B.n586 585
R226 B.n588 B.n69 585
R227 B.n590 B.n589 585
R228 B.n591 B.n68 585
R229 B.n593 B.n592 585
R230 B.n594 B.n67 585
R231 B.n596 B.n595 585
R232 B.n597 B.n66 585
R233 B.n599 B.n598 585
R234 B.n600 B.n65 585
R235 B.n602 B.n601 585
R236 B.n603 B.n64 585
R237 B.n605 B.n604 585
R238 B.n606 B.n63 585
R239 B.n608 B.n607 585
R240 B.n609 B.n62 585
R241 B.n611 B.n610 585
R242 B.n612 B.n61 585
R243 B.n614 B.n613 585
R244 B.n615 B.n60 585
R245 B.n617 B.n616 585
R246 B.n618 B.n59 585
R247 B.n620 B.n619 585
R248 B.n621 B.n58 585
R249 B.n623 B.n622 585
R250 B.n624 B.n57 585
R251 B.n626 B.n625 585
R252 B.n628 B.n627 585
R253 B.n629 B.n53 585
R254 B.n631 B.n630 585
R255 B.n632 B.n52 585
R256 B.n634 B.n633 585
R257 B.n635 B.n51 585
R258 B.n637 B.n636 585
R259 B.n638 B.n50 585
R260 B.n640 B.n639 585
R261 B.n642 B.n47 585
R262 B.n644 B.n643 585
R263 B.n645 B.n46 585
R264 B.n647 B.n646 585
R265 B.n648 B.n45 585
R266 B.n650 B.n649 585
R267 B.n651 B.n44 585
R268 B.n653 B.n652 585
R269 B.n654 B.n43 585
R270 B.n656 B.n655 585
R271 B.n657 B.n42 585
R272 B.n659 B.n658 585
R273 B.n660 B.n41 585
R274 B.n662 B.n661 585
R275 B.n663 B.n40 585
R276 B.n665 B.n664 585
R277 B.n666 B.n39 585
R278 B.n668 B.n667 585
R279 B.n669 B.n38 585
R280 B.n671 B.n670 585
R281 B.n672 B.n37 585
R282 B.n674 B.n673 585
R283 B.n675 B.n36 585
R284 B.n677 B.n676 585
R285 B.n678 B.n35 585
R286 B.n680 B.n679 585
R287 B.n681 B.n34 585
R288 B.n683 B.n682 585
R289 B.n684 B.n33 585
R290 B.n686 B.n685 585
R291 B.n687 B.n32 585
R292 B.n689 B.n688 585
R293 B.n690 B.n31 585
R294 B.n692 B.n691 585
R295 B.n693 B.n30 585
R296 B.n695 B.n694 585
R297 B.n696 B.n29 585
R298 B.n698 B.n697 585
R299 B.n699 B.n28 585
R300 B.n701 B.n700 585
R301 B.n702 B.n27 585
R302 B.n704 B.n703 585
R303 B.n705 B.n26 585
R304 B.n707 B.n706 585
R305 B.n708 B.n25 585
R306 B.n710 B.n709 585
R307 B.n711 B.n24 585
R308 B.n713 B.n712 585
R309 B.n714 B.n23 585
R310 B.n716 B.n715 585
R311 B.n717 B.n22 585
R312 B.n719 B.n718 585
R313 B.n720 B.n21 585
R314 B.n722 B.n721 585
R315 B.n723 B.n20 585
R316 B.n725 B.n724 585
R317 B.n726 B.n19 585
R318 B.n728 B.n727 585
R319 B.n729 B.n18 585
R320 B.n731 B.n730 585
R321 B.n732 B.n17 585
R322 B.n734 B.n733 585
R323 B.n735 B.n16 585
R324 B.n737 B.n736 585
R325 B.n738 B.n15 585
R326 B.n528 B.n89 585
R327 B.n527 B.n526 585
R328 B.n525 B.n90 585
R329 B.n524 B.n523 585
R330 B.n522 B.n91 585
R331 B.n521 B.n520 585
R332 B.n519 B.n92 585
R333 B.n518 B.n517 585
R334 B.n516 B.n93 585
R335 B.n515 B.n514 585
R336 B.n513 B.n94 585
R337 B.n512 B.n511 585
R338 B.n510 B.n95 585
R339 B.n509 B.n508 585
R340 B.n507 B.n96 585
R341 B.n506 B.n505 585
R342 B.n504 B.n97 585
R343 B.n503 B.n502 585
R344 B.n501 B.n98 585
R345 B.n500 B.n499 585
R346 B.n498 B.n99 585
R347 B.n497 B.n496 585
R348 B.n495 B.n100 585
R349 B.n494 B.n493 585
R350 B.n492 B.n101 585
R351 B.n491 B.n490 585
R352 B.n489 B.n102 585
R353 B.n488 B.n487 585
R354 B.n486 B.n103 585
R355 B.n485 B.n484 585
R356 B.n483 B.n104 585
R357 B.n482 B.n481 585
R358 B.n480 B.n105 585
R359 B.n479 B.n478 585
R360 B.n477 B.n106 585
R361 B.n476 B.n475 585
R362 B.n474 B.n107 585
R363 B.n473 B.n472 585
R364 B.n471 B.n108 585
R365 B.n470 B.n469 585
R366 B.n468 B.n109 585
R367 B.n467 B.n466 585
R368 B.n465 B.n110 585
R369 B.n464 B.n463 585
R370 B.n462 B.n111 585
R371 B.n461 B.n460 585
R372 B.n459 B.n112 585
R373 B.n458 B.n457 585
R374 B.n456 B.n113 585
R375 B.n455 B.n454 585
R376 B.n453 B.n114 585
R377 B.n452 B.n451 585
R378 B.n450 B.n115 585
R379 B.n240 B.n189 585
R380 B.n242 B.n241 585
R381 B.n243 B.n188 585
R382 B.n245 B.n244 585
R383 B.n246 B.n187 585
R384 B.n248 B.n247 585
R385 B.n249 B.n186 585
R386 B.n251 B.n250 585
R387 B.n252 B.n185 585
R388 B.n254 B.n253 585
R389 B.n255 B.n184 585
R390 B.n257 B.n256 585
R391 B.n258 B.n183 585
R392 B.n260 B.n259 585
R393 B.n261 B.n182 585
R394 B.n263 B.n262 585
R395 B.n264 B.n181 585
R396 B.n266 B.n265 585
R397 B.n267 B.n180 585
R398 B.n269 B.n268 585
R399 B.n270 B.n179 585
R400 B.n272 B.n271 585
R401 B.n273 B.n178 585
R402 B.n275 B.n274 585
R403 B.n276 B.n177 585
R404 B.n278 B.n277 585
R405 B.n279 B.n176 585
R406 B.n281 B.n280 585
R407 B.n282 B.n175 585
R408 B.n284 B.n283 585
R409 B.n285 B.n174 585
R410 B.n287 B.n286 585
R411 B.n288 B.n173 585
R412 B.n290 B.n289 585
R413 B.n291 B.n172 585
R414 B.n293 B.n292 585
R415 B.n294 B.n171 585
R416 B.n296 B.n295 585
R417 B.n297 B.n170 585
R418 B.n299 B.n298 585
R419 B.n300 B.n169 585
R420 B.n302 B.n301 585
R421 B.n303 B.n168 585
R422 B.n305 B.n304 585
R423 B.n306 B.n167 585
R424 B.n308 B.n307 585
R425 B.n309 B.n166 585
R426 B.n311 B.n310 585
R427 B.n312 B.n165 585
R428 B.n314 B.n313 585
R429 B.n315 B.n164 585
R430 B.n317 B.n316 585
R431 B.n318 B.n163 585
R432 B.n320 B.n319 585
R433 B.n321 B.n162 585
R434 B.n323 B.n322 585
R435 B.n324 B.n161 585
R436 B.n326 B.n325 585
R437 B.n327 B.n160 585
R438 B.n329 B.n328 585
R439 B.n330 B.n159 585
R440 B.n332 B.n331 585
R441 B.n333 B.n158 585
R442 B.n335 B.n334 585
R443 B.n336 B.n155 585
R444 B.n339 B.n338 585
R445 B.n340 B.n154 585
R446 B.n342 B.n341 585
R447 B.n343 B.n153 585
R448 B.n345 B.n344 585
R449 B.n346 B.n152 585
R450 B.n348 B.n347 585
R451 B.n349 B.n151 585
R452 B.n351 B.n350 585
R453 B.n353 B.n352 585
R454 B.n354 B.n147 585
R455 B.n356 B.n355 585
R456 B.n357 B.n146 585
R457 B.n359 B.n358 585
R458 B.n360 B.n145 585
R459 B.n362 B.n361 585
R460 B.n363 B.n144 585
R461 B.n365 B.n364 585
R462 B.n366 B.n143 585
R463 B.n368 B.n367 585
R464 B.n369 B.n142 585
R465 B.n371 B.n370 585
R466 B.n372 B.n141 585
R467 B.n374 B.n373 585
R468 B.n375 B.n140 585
R469 B.n377 B.n376 585
R470 B.n378 B.n139 585
R471 B.n380 B.n379 585
R472 B.n381 B.n138 585
R473 B.n383 B.n382 585
R474 B.n384 B.n137 585
R475 B.n386 B.n385 585
R476 B.n387 B.n136 585
R477 B.n389 B.n388 585
R478 B.n390 B.n135 585
R479 B.n392 B.n391 585
R480 B.n393 B.n134 585
R481 B.n395 B.n394 585
R482 B.n396 B.n133 585
R483 B.n398 B.n397 585
R484 B.n399 B.n132 585
R485 B.n401 B.n400 585
R486 B.n402 B.n131 585
R487 B.n404 B.n403 585
R488 B.n405 B.n130 585
R489 B.n407 B.n406 585
R490 B.n408 B.n129 585
R491 B.n410 B.n409 585
R492 B.n411 B.n128 585
R493 B.n413 B.n412 585
R494 B.n414 B.n127 585
R495 B.n416 B.n415 585
R496 B.n417 B.n126 585
R497 B.n419 B.n418 585
R498 B.n420 B.n125 585
R499 B.n422 B.n421 585
R500 B.n423 B.n124 585
R501 B.n425 B.n424 585
R502 B.n426 B.n123 585
R503 B.n428 B.n427 585
R504 B.n429 B.n122 585
R505 B.n431 B.n430 585
R506 B.n432 B.n121 585
R507 B.n434 B.n433 585
R508 B.n435 B.n120 585
R509 B.n437 B.n436 585
R510 B.n438 B.n119 585
R511 B.n440 B.n439 585
R512 B.n441 B.n118 585
R513 B.n443 B.n442 585
R514 B.n444 B.n117 585
R515 B.n446 B.n445 585
R516 B.n447 B.n116 585
R517 B.n449 B.n448 585
R518 B.n239 B.n238 585
R519 B.n237 B.n190 585
R520 B.n236 B.n235 585
R521 B.n234 B.n191 585
R522 B.n233 B.n232 585
R523 B.n231 B.n192 585
R524 B.n230 B.n229 585
R525 B.n228 B.n193 585
R526 B.n227 B.n226 585
R527 B.n225 B.n194 585
R528 B.n224 B.n223 585
R529 B.n222 B.n195 585
R530 B.n221 B.n220 585
R531 B.n219 B.n196 585
R532 B.n218 B.n217 585
R533 B.n216 B.n197 585
R534 B.n215 B.n214 585
R535 B.n213 B.n198 585
R536 B.n212 B.n211 585
R537 B.n210 B.n199 585
R538 B.n209 B.n208 585
R539 B.n207 B.n200 585
R540 B.n206 B.n205 585
R541 B.n204 B.n201 585
R542 B.n203 B.n202 585
R543 B.n2 B.n0 585
R544 B.n777 B.n1 585
R545 B.n776 B.n775 585
R546 B.n774 B.n3 585
R547 B.n773 B.n772 585
R548 B.n771 B.n4 585
R549 B.n770 B.n769 585
R550 B.n768 B.n5 585
R551 B.n767 B.n766 585
R552 B.n765 B.n6 585
R553 B.n764 B.n763 585
R554 B.n762 B.n7 585
R555 B.n761 B.n760 585
R556 B.n759 B.n8 585
R557 B.n758 B.n757 585
R558 B.n756 B.n9 585
R559 B.n755 B.n754 585
R560 B.n753 B.n10 585
R561 B.n752 B.n751 585
R562 B.n750 B.n11 585
R563 B.n749 B.n748 585
R564 B.n747 B.n12 585
R565 B.n746 B.n745 585
R566 B.n744 B.n13 585
R567 B.n743 B.n742 585
R568 B.n741 B.n14 585
R569 B.n740 B.n739 585
R570 B.n779 B.n778 585
R571 B.n238 B.n189 540.549
R572 B.n740 B.n15 540.549
R573 B.n448 B.n115 540.549
R574 B.n530 B.n89 540.549
R575 B.n238 B.n237 163.367
R576 B.n237 B.n236 163.367
R577 B.n236 B.n191 163.367
R578 B.n232 B.n191 163.367
R579 B.n232 B.n231 163.367
R580 B.n231 B.n230 163.367
R581 B.n230 B.n193 163.367
R582 B.n226 B.n193 163.367
R583 B.n226 B.n225 163.367
R584 B.n225 B.n224 163.367
R585 B.n224 B.n195 163.367
R586 B.n220 B.n195 163.367
R587 B.n220 B.n219 163.367
R588 B.n219 B.n218 163.367
R589 B.n218 B.n197 163.367
R590 B.n214 B.n197 163.367
R591 B.n214 B.n213 163.367
R592 B.n213 B.n212 163.367
R593 B.n212 B.n199 163.367
R594 B.n208 B.n199 163.367
R595 B.n208 B.n207 163.367
R596 B.n207 B.n206 163.367
R597 B.n206 B.n201 163.367
R598 B.n202 B.n201 163.367
R599 B.n202 B.n2 163.367
R600 B.n778 B.n2 163.367
R601 B.n778 B.n777 163.367
R602 B.n777 B.n776 163.367
R603 B.n776 B.n3 163.367
R604 B.n772 B.n3 163.367
R605 B.n772 B.n771 163.367
R606 B.n771 B.n770 163.367
R607 B.n770 B.n5 163.367
R608 B.n766 B.n5 163.367
R609 B.n766 B.n765 163.367
R610 B.n765 B.n764 163.367
R611 B.n764 B.n7 163.367
R612 B.n760 B.n7 163.367
R613 B.n760 B.n759 163.367
R614 B.n759 B.n758 163.367
R615 B.n758 B.n9 163.367
R616 B.n754 B.n9 163.367
R617 B.n754 B.n753 163.367
R618 B.n753 B.n752 163.367
R619 B.n752 B.n11 163.367
R620 B.n748 B.n11 163.367
R621 B.n748 B.n747 163.367
R622 B.n747 B.n746 163.367
R623 B.n746 B.n13 163.367
R624 B.n742 B.n13 163.367
R625 B.n742 B.n741 163.367
R626 B.n741 B.n740 163.367
R627 B.n242 B.n189 163.367
R628 B.n243 B.n242 163.367
R629 B.n244 B.n243 163.367
R630 B.n244 B.n187 163.367
R631 B.n248 B.n187 163.367
R632 B.n249 B.n248 163.367
R633 B.n250 B.n249 163.367
R634 B.n250 B.n185 163.367
R635 B.n254 B.n185 163.367
R636 B.n255 B.n254 163.367
R637 B.n256 B.n255 163.367
R638 B.n256 B.n183 163.367
R639 B.n260 B.n183 163.367
R640 B.n261 B.n260 163.367
R641 B.n262 B.n261 163.367
R642 B.n262 B.n181 163.367
R643 B.n266 B.n181 163.367
R644 B.n267 B.n266 163.367
R645 B.n268 B.n267 163.367
R646 B.n268 B.n179 163.367
R647 B.n272 B.n179 163.367
R648 B.n273 B.n272 163.367
R649 B.n274 B.n273 163.367
R650 B.n274 B.n177 163.367
R651 B.n278 B.n177 163.367
R652 B.n279 B.n278 163.367
R653 B.n280 B.n279 163.367
R654 B.n280 B.n175 163.367
R655 B.n284 B.n175 163.367
R656 B.n285 B.n284 163.367
R657 B.n286 B.n285 163.367
R658 B.n286 B.n173 163.367
R659 B.n290 B.n173 163.367
R660 B.n291 B.n290 163.367
R661 B.n292 B.n291 163.367
R662 B.n292 B.n171 163.367
R663 B.n296 B.n171 163.367
R664 B.n297 B.n296 163.367
R665 B.n298 B.n297 163.367
R666 B.n298 B.n169 163.367
R667 B.n302 B.n169 163.367
R668 B.n303 B.n302 163.367
R669 B.n304 B.n303 163.367
R670 B.n304 B.n167 163.367
R671 B.n308 B.n167 163.367
R672 B.n309 B.n308 163.367
R673 B.n310 B.n309 163.367
R674 B.n310 B.n165 163.367
R675 B.n314 B.n165 163.367
R676 B.n315 B.n314 163.367
R677 B.n316 B.n315 163.367
R678 B.n316 B.n163 163.367
R679 B.n320 B.n163 163.367
R680 B.n321 B.n320 163.367
R681 B.n322 B.n321 163.367
R682 B.n322 B.n161 163.367
R683 B.n326 B.n161 163.367
R684 B.n327 B.n326 163.367
R685 B.n328 B.n327 163.367
R686 B.n328 B.n159 163.367
R687 B.n332 B.n159 163.367
R688 B.n333 B.n332 163.367
R689 B.n334 B.n333 163.367
R690 B.n334 B.n155 163.367
R691 B.n339 B.n155 163.367
R692 B.n340 B.n339 163.367
R693 B.n341 B.n340 163.367
R694 B.n341 B.n153 163.367
R695 B.n345 B.n153 163.367
R696 B.n346 B.n345 163.367
R697 B.n347 B.n346 163.367
R698 B.n347 B.n151 163.367
R699 B.n351 B.n151 163.367
R700 B.n352 B.n351 163.367
R701 B.n352 B.n147 163.367
R702 B.n356 B.n147 163.367
R703 B.n357 B.n356 163.367
R704 B.n358 B.n357 163.367
R705 B.n358 B.n145 163.367
R706 B.n362 B.n145 163.367
R707 B.n363 B.n362 163.367
R708 B.n364 B.n363 163.367
R709 B.n364 B.n143 163.367
R710 B.n368 B.n143 163.367
R711 B.n369 B.n368 163.367
R712 B.n370 B.n369 163.367
R713 B.n370 B.n141 163.367
R714 B.n374 B.n141 163.367
R715 B.n375 B.n374 163.367
R716 B.n376 B.n375 163.367
R717 B.n376 B.n139 163.367
R718 B.n380 B.n139 163.367
R719 B.n381 B.n380 163.367
R720 B.n382 B.n381 163.367
R721 B.n382 B.n137 163.367
R722 B.n386 B.n137 163.367
R723 B.n387 B.n386 163.367
R724 B.n388 B.n387 163.367
R725 B.n388 B.n135 163.367
R726 B.n392 B.n135 163.367
R727 B.n393 B.n392 163.367
R728 B.n394 B.n393 163.367
R729 B.n394 B.n133 163.367
R730 B.n398 B.n133 163.367
R731 B.n399 B.n398 163.367
R732 B.n400 B.n399 163.367
R733 B.n400 B.n131 163.367
R734 B.n404 B.n131 163.367
R735 B.n405 B.n404 163.367
R736 B.n406 B.n405 163.367
R737 B.n406 B.n129 163.367
R738 B.n410 B.n129 163.367
R739 B.n411 B.n410 163.367
R740 B.n412 B.n411 163.367
R741 B.n412 B.n127 163.367
R742 B.n416 B.n127 163.367
R743 B.n417 B.n416 163.367
R744 B.n418 B.n417 163.367
R745 B.n418 B.n125 163.367
R746 B.n422 B.n125 163.367
R747 B.n423 B.n422 163.367
R748 B.n424 B.n423 163.367
R749 B.n424 B.n123 163.367
R750 B.n428 B.n123 163.367
R751 B.n429 B.n428 163.367
R752 B.n430 B.n429 163.367
R753 B.n430 B.n121 163.367
R754 B.n434 B.n121 163.367
R755 B.n435 B.n434 163.367
R756 B.n436 B.n435 163.367
R757 B.n436 B.n119 163.367
R758 B.n440 B.n119 163.367
R759 B.n441 B.n440 163.367
R760 B.n442 B.n441 163.367
R761 B.n442 B.n117 163.367
R762 B.n446 B.n117 163.367
R763 B.n447 B.n446 163.367
R764 B.n448 B.n447 163.367
R765 B.n452 B.n115 163.367
R766 B.n453 B.n452 163.367
R767 B.n454 B.n453 163.367
R768 B.n454 B.n113 163.367
R769 B.n458 B.n113 163.367
R770 B.n459 B.n458 163.367
R771 B.n460 B.n459 163.367
R772 B.n460 B.n111 163.367
R773 B.n464 B.n111 163.367
R774 B.n465 B.n464 163.367
R775 B.n466 B.n465 163.367
R776 B.n466 B.n109 163.367
R777 B.n470 B.n109 163.367
R778 B.n471 B.n470 163.367
R779 B.n472 B.n471 163.367
R780 B.n472 B.n107 163.367
R781 B.n476 B.n107 163.367
R782 B.n477 B.n476 163.367
R783 B.n478 B.n477 163.367
R784 B.n478 B.n105 163.367
R785 B.n482 B.n105 163.367
R786 B.n483 B.n482 163.367
R787 B.n484 B.n483 163.367
R788 B.n484 B.n103 163.367
R789 B.n488 B.n103 163.367
R790 B.n489 B.n488 163.367
R791 B.n490 B.n489 163.367
R792 B.n490 B.n101 163.367
R793 B.n494 B.n101 163.367
R794 B.n495 B.n494 163.367
R795 B.n496 B.n495 163.367
R796 B.n496 B.n99 163.367
R797 B.n500 B.n99 163.367
R798 B.n501 B.n500 163.367
R799 B.n502 B.n501 163.367
R800 B.n502 B.n97 163.367
R801 B.n506 B.n97 163.367
R802 B.n507 B.n506 163.367
R803 B.n508 B.n507 163.367
R804 B.n508 B.n95 163.367
R805 B.n512 B.n95 163.367
R806 B.n513 B.n512 163.367
R807 B.n514 B.n513 163.367
R808 B.n514 B.n93 163.367
R809 B.n518 B.n93 163.367
R810 B.n519 B.n518 163.367
R811 B.n520 B.n519 163.367
R812 B.n520 B.n91 163.367
R813 B.n524 B.n91 163.367
R814 B.n525 B.n524 163.367
R815 B.n526 B.n525 163.367
R816 B.n526 B.n89 163.367
R817 B.n736 B.n15 163.367
R818 B.n736 B.n735 163.367
R819 B.n735 B.n734 163.367
R820 B.n734 B.n17 163.367
R821 B.n730 B.n17 163.367
R822 B.n730 B.n729 163.367
R823 B.n729 B.n728 163.367
R824 B.n728 B.n19 163.367
R825 B.n724 B.n19 163.367
R826 B.n724 B.n723 163.367
R827 B.n723 B.n722 163.367
R828 B.n722 B.n21 163.367
R829 B.n718 B.n21 163.367
R830 B.n718 B.n717 163.367
R831 B.n717 B.n716 163.367
R832 B.n716 B.n23 163.367
R833 B.n712 B.n23 163.367
R834 B.n712 B.n711 163.367
R835 B.n711 B.n710 163.367
R836 B.n710 B.n25 163.367
R837 B.n706 B.n25 163.367
R838 B.n706 B.n705 163.367
R839 B.n705 B.n704 163.367
R840 B.n704 B.n27 163.367
R841 B.n700 B.n27 163.367
R842 B.n700 B.n699 163.367
R843 B.n699 B.n698 163.367
R844 B.n698 B.n29 163.367
R845 B.n694 B.n29 163.367
R846 B.n694 B.n693 163.367
R847 B.n693 B.n692 163.367
R848 B.n692 B.n31 163.367
R849 B.n688 B.n31 163.367
R850 B.n688 B.n687 163.367
R851 B.n687 B.n686 163.367
R852 B.n686 B.n33 163.367
R853 B.n682 B.n33 163.367
R854 B.n682 B.n681 163.367
R855 B.n681 B.n680 163.367
R856 B.n680 B.n35 163.367
R857 B.n676 B.n35 163.367
R858 B.n676 B.n675 163.367
R859 B.n675 B.n674 163.367
R860 B.n674 B.n37 163.367
R861 B.n670 B.n37 163.367
R862 B.n670 B.n669 163.367
R863 B.n669 B.n668 163.367
R864 B.n668 B.n39 163.367
R865 B.n664 B.n39 163.367
R866 B.n664 B.n663 163.367
R867 B.n663 B.n662 163.367
R868 B.n662 B.n41 163.367
R869 B.n658 B.n41 163.367
R870 B.n658 B.n657 163.367
R871 B.n657 B.n656 163.367
R872 B.n656 B.n43 163.367
R873 B.n652 B.n43 163.367
R874 B.n652 B.n651 163.367
R875 B.n651 B.n650 163.367
R876 B.n650 B.n45 163.367
R877 B.n646 B.n45 163.367
R878 B.n646 B.n645 163.367
R879 B.n645 B.n644 163.367
R880 B.n644 B.n47 163.367
R881 B.n639 B.n47 163.367
R882 B.n639 B.n638 163.367
R883 B.n638 B.n637 163.367
R884 B.n637 B.n51 163.367
R885 B.n633 B.n51 163.367
R886 B.n633 B.n632 163.367
R887 B.n632 B.n631 163.367
R888 B.n631 B.n53 163.367
R889 B.n627 B.n53 163.367
R890 B.n627 B.n626 163.367
R891 B.n626 B.n57 163.367
R892 B.n622 B.n57 163.367
R893 B.n622 B.n621 163.367
R894 B.n621 B.n620 163.367
R895 B.n620 B.n59 163.367
R896 B.n616 B.n59 163.367
R897 B.n616 B.n615 163.367
R898 B.n615 B.n614 163.367
R899 B.n614 B.n61 163.367
R900 B.n610 B.n61 163.367
R901 B.n610 B.n609 163.367
R902 B.n609 B.n608 163.367
R903 B.n608 B.n63 163.367
R904 B.n604 B.n63 163.367
R905 B.n604 B.n603 163.367
R906 B.n603 B.n602 163.367
R907 B.n602 B.n65 163.367
R908 B.n598 B.n65 163.367
R909 B.n598 B.n597 163.367
R910 B.n597 B.n596 163.367
R911 B.n596 B.n67 163.367
R912 B.n592 B.n67 163.367
R913 B.n592 B.n591 163.367
R914 B.n591 B.n590 163.367
R915 B.n590 B.n69 163.367
R916 B.n586 B.n69 163.367
R917 B.n586 B.n585 163.367
R918 B.n585 B.n584 163.367
R919 B.n584 B.n71 163.367
R920 B.n580 B.n71 163.367
R921 B.n580 B.n579 163.367
R922 B.n579 B.n578 163.367
R923 B.n578 B.n73 163.367
R924 B.n574 B.n73 163.367
R925 B.n574 B.n573 163.367
R926 B.n573 B.n572 163.367
R927 B.n572 B.n75 163.367
R928 B.n568 B.n75 163.367
R929 B.n568 B.n567 163.367
R930 B.n567 B.n566 163.367
R931 B.n566 B.n77 163.367
R932 B.n562 B.n77 163.367
R933 B.n562 B.n561 163.367
R934 B.n561 B.n560 163.367
R935 B.n560 B.n79 163.367
R936 B.n556 B.n79 163.367
R937 B.n556 B.n555 163.367
R938 B.n555 B.n554 163.367
R939 B.n554 B.n81 163.367
R940 B.n550 B.n81 163.367
R941 B.n550 B.n549 163.367
R942 B.n549 B.n548 163.367
R943 B.n548 B.n83 163.367
R944 B.n544 B.n83 163.367
R945 B.n544 B.n543 163.367
R946 B.n543 B.n542 163.367
R947 B.n542 B.n85 163.367
R948 B.n538 B.n85 163.367
R949 B.n538 B.n537 163.367
R950 B.n537 B.n536 163.367
R951 B.n536 B.n87 163.367
R952 B.n532 B.n87 163.367
R953 B.n532 B.n531 163.367
R954 B.n531 B.n530 163.367
R955 B.n148 B.t8 128.343
R956 B.n54 B.t10 128.343
R957 B.n156 B.t5 128.316
R958 B.n48 B.t1 128.316
R959 B.n149 B.t7 108.367
R960 B.n55 B.t11 108.367
R961 B.n157 B.t4 108.341
R962 B.n49 B.t2 108.341
R963 B.n150 B.n149 59.5399
R964 B.n337 B.n157 59.5399
R965 B.n641 B.n49 59.5399
R966 B.n56 B.n55 59.5399
R967 B.n739 B.n738 35.1225
R968 B.n529 B.n528 35.1225
R969 B.n450 B.n449 35.1225
R970 B.n240 B.n239 35.1225
R971 B.n149 B.n148 19.9763
R972 B.n157 B.n156 19.9763
R973 B.n49 B.n48 19.9763
R974 B.n55 B.n54 19.9763
R975 B B.n779 18.0485
R976 B.n738 B.n737 10.6151
R977 B.n737 B.n16 10.6151
R978 B.n733 B.n16 10.6151
R979 B.n733 B.n732 10.6151
R980 B.n732 B.n731 10.6151
R981 B.n731 B.n18 10.6151
R982 B.n727 B.n18 10.6151
R983 B.n727 B.n726 10.6151
R984 B.n726 B.n725 10.6151
R985 B.n725 B.n20 10.6151
R986 B.n721 B.n20 10.6151
R987 B.n721 B.n720 10.6151
R988 B.n720 B.n719 10.6151
R989 B.n719 B.n22 10.6151
R990 B.n715 B.n22 10.6151
R991 B.n715 B.n714 10.6151
R992 B.n714 B.n713 10.6151
R993 B.n713 B.n24 10.6151
R994 B.n709 B.n24 10.6151
R995 B.n709 B.n708 10.6151
R996 B.n708 B.n707 10.6151
R997 B.n707 B.n26 10.6151
R998 B.n703 B.n26 10.6151
R999 B.n703 B.n702 10.6151
R1000 B.n702 B.n701 10.6151
R1001 B.n701 B.n28 10.6151
R1002 B.n697 B.n28 10.6151
R1003 B.n697 B.n696 10.6151
R1004 B.n696 B.n695 10.6151
R1005 B.n695 B.n30 10.6151
R1006 B.n691 B.n30 10.6151
R1007 B.n691 B.n690 10.6151
R1008 B.n690 B.n689 10.6151
R1009 B.n689 B.n32 10.6151
R1010 B.n685 B.n32 10.6151
R1011 B.n685 B.n684 10.6151
R1012 B.n684 B.n683 10.6151
R1013 B.n683 B.n34 10.6151
R1014 B.n679 B.n34 10.6151
R1015 B.n679 B.n678 10.6151
R1016 B.n678 B.n677 10.6151
R1017 B.n677 B.n36 10.6151
R1018 B.n673 B.n36 10.6151
R1019 B.n673 B.n672 10.6151
R1020 B.n672 B.n671 10.6151
R1021 B.n671 B.n38 10.6151
R1022 B.n667 B.n38 10.6151
R1023 B.n667 B.n666 10.6151
R1024 B.n666 B.n665 10.6151
R1025 B.n665 B.n40 10.6151
R1026 B.n661 B.n40 10.6151
R1027 B.n661 B.n660 10.6151
R1028 B.n660 B.n659 10.6151
R1029 B.n659 B.n42 10.6151
R1030 B.n655 B.n42 10.6151
R1031 B.n655 B.n654 10.6151
R1032 B.n654 B.n653 10.6151
R1033 B.n653 B.n44 10.6151
R1034 B.n649 B.n44 10.6151
R1035 B.n649 B.n648 10.6151
R1036 B.n648 B.n647 10.6151
R1037 B.n647 B.n46 10.6151
R1038 B.n643 B.n46 10.6151
R1039 B.n643 B.n642 10.6151
R1040 B.n640 B.n50 10.6151
R1041 B.n636 B.n50 10.6151
R1042 B.n636 B.n635 10.6151
R1043 B.n635 B.n634 10.6151
R1044 B.n634 B.n52 10.6151
R1045 B.n630 B.n52 10.6151
R1046 B.n630 B.n629 10.6151
R1047 B.n629 B.n628 10.6151
R1048 B.n625 B.n624 10.6151
R1049 B.n624 B.n623 10.6151
R1050 B.n623 B.n58 10.6151
R1051 B.n619 B.n58 10.6151
R1052 B.n619 B.n618 10.6151
R1053 B.n618 B.n617 10.6151
R1054 B.n617 B.n60 10.6151
R1055 B.n613 B.n60 10.6151
R1056 B.n613 B.n612 10.6151
R1057 B.n612 B.n611 10.6151
R1058 B.n611 B.n62 10.6151
R1059 B.n607 B.n62 10.6151
R1060 B.n607 B.n606 10.6151
R1061 B.n606 B.n605 10.6151
R1062 B.n605 B.n64 10.6151
R1063 B.n601 B.n64 10.6151
R1064 B.n601 B.n600 10.6151
R1065 B.n600 B.n599 10.6151
R1066 B.n599 B.n66 10.6151
R1067 B.n595 B.n66 10.6151
R1068 B.n595 B.n594 10.6151
R1069 B.n594 B.n593 10.6151
R1070 B.n593 B.n68 10.6151
R1071 B.n589 B.n68 10.6151
R1072 B.n589 B.n588 10.6151
R1073 B.n588 B.n587 10.6151
R1074 B.n587 B.n70 10.6151
R1075 B.n583 B.n70 10.6151
R1076 B.n583 B.n582 10.6151
R1077 B.n582 B.n581 10.6151
R1078 B.n581 B.n72 10.6151
R1079 B.n577 B.n72 10.6151
R1080 B.n577 B.n576 10.6151
R1081 B.n576 B.n575 10.6151
R1082 B.n575 B.n74 10.6151
R1083 B.n571 B.n74 10.6151
R1084 B.n571 B.n570 10.6151
R1085 B.n570 B.n569 10.6151
R1086 B.n569 B.n76 10.6151
R1087 B.n565 B.n76 10.6151
R1088 B.n565 B.n564 10.6151
R1089 B.n564 B.n563 10.6151
R1090 B.n563 B.n78 10.6151
R1091 B.n559 B.n78 10.6151
R1092 B.n559 B.n558 10.6151
R1093 B.n558 B.n557 10.6151
R1094 B.n557 B.n80 10.6151
R1095 B.n553 B.n80 10.6151
R1096 B.n553 B.n552 10.6151
R1097 B.n552 B.n551 10.6151
R1098 B.n551 B.n82 10.6151
R1099 B.n547 B.n82 10.6151
R1100 B.n547 B.n546 10.6151
R1101 B.n546 B.n545 10.6151
R1102 B.n545 B.n84 10.6151
R1103 B.n541 B.n84 10.6151
R1104 B.n541 B.n540 10.6151
R1105 B.n540 B.n539 10.6151
R1106 B.n539 B.n86 10.6151
R1107 B.n535 B.n86 10.6151
R1108 B.n535 B.n534 10.6151
R1109 B.n534 B.n533 10.6151
R1110 B.n533 B.n88 10.6151
R1111 B.n529 B.n88 10.6151
R1112 B.n451 B.n450 10.6151
R1113 B.n451 B.n114 10.6151
R1114 B.n455 B.n114 10.6151
R1115 B.n456 B.n455 10.6151
R1116 B.n457 B.n456 10.6151
R1117 B.n457 B.n112 10.6151
R1118 B.n461 B.n112 10.6151
R1119 B.n462 B.n461 10.6151
R1120 B.n463 B.n462 10.6151
R1121 B.n463 B.n110 10.6151
R1122 B.n467 B.n110 10.6151
R1123 B.n468 B.n467 10.6151
R1124 B.n469 B.n468 10.6151
R1125 B.n469 B.n108 10.6151
R1126 B.n473 B.n108 10.6151
R1127 B.n474 B.n473 10.6151
R1128 B.n475 B.n474 10.6151
R1129 B.n475 B.n106 10.6151
R1130 B.n479 B.n106 10.6151
R1131 B.n480 B.n479 10.6151
R1132 B.n481 B.n480 10.6151
R1133 B.n481 B.n104 10.6151
R1134 B.n485 B.n104 10.6151
R1135 B.n486 B.n485 10.6151
R1136 B.n487 B.n486 10.6151
R1137 B.n487 B.n102 10.6151
R1138 B.n491 B.n102 10.6151
R1139 B.n492 B.n491 10.6151
R1140 B.n493 B.n492 10.6151
R1141 B.n493 B.n100 10.6151
R1142 B.n497 B.n100 10.6151
R1143 B.n498 B.n497 10.6151
R1144 B.n499 B.n498 10.6151
R1145 B.n499 B.n98 10.6151
R1146 B.n503 B.n98 10.6151
R1147 B.n504 B.n503 10.6151
R1148 B.n505 B.n504 10.6151
R1149 B.n505 B.n96 10.6151
R1150 B.n509 B.n96 10.6151
R1151 B.n510 B.n509 10.6151
R1152 B.n511 B.n510 10.6151
R1153 B.n511 B.n94 10.6151
R1154 B.n515 B.n94 10.6151
R1155 B.n516 B.n515 10.6151
R1156 B.n517 B.n516 10.6151
R1157 B.n517 B.n92 10.6151
R1158 B.n521 B.n92 10.6151
R1159 B.n522 B.n521 10.6151
R1160 B.n523 B.n522 10.6151
R1161 B.n523 B.n90 10.6151
R1162 B.n527 B.n90 10.6151
R1163 B.n528 B.n527 10.6151
R1164 B.n241 B.n240 10.6151
R1165 B.n241 B.n188 10.6151
R1166 B.n245 B.n188 10.6151
R1167 B.n246 B.n245 10.6151
R1168 B.n247 B.n246 10.6151
R1169 B.n247 B.n186 10.6151
R1170 B.n251 B.n186 10.6151
R1171 B.n252 B.n251 10.6151
R1172 B.n253 B.n252 10.6151
R1173 B.n253 B.n184 10.6151
R1174 B.n257 B.n184 10.6151
R1175 B.n258 B.n257 10.6151
R1176 B.n259 B.n258 10.6151
R1177 B.n259 B.n182 10.6151
R1178 B.n263 B.n182 10.6151
R1179 B.n264 B.n263 10.6151
R1180 B.n265 B.n264 10.6151
R1181 B.n265 B.n180 10.6151
R1182 B.n269 B.n180 10.6151
R1183 B.n270 B.n269 10.6151
R1184 B.n271 B.n270 10.6151
R1185 B.n271 B.n178 10.6151
R1186 B.n275 B.n178 10.6151
R1187 B.n276 B.n275 10.6151
R1188 B.n277 B.n276 10.6151
R1189 B.n277 B.n176 10.6151
R1190 B.n281 B.n176 10.6151
R1191 B.n282 B.n281 10.6151
R1192 B.n283 B.n282 10.6151
R1193 B.n283 B.n174 10.6151
R1194 B.n287 B.n174 10.6151
R1195 B.n288 B.n287 10.6151
R1196 B.n289 B.n288 10.6151
R1197 B.n289 B.n172 10.6151
R1198 B.n293 B.n172 10.6151
R1199 B.n294 B.n293 10.6151
R1200 B.n295 B.n294 10.6151
R1201 B.n295 B.n170 10.6151
R1202 B.n299 B.n170 10.6151
R1203 B.n300 B.n299 10.6151
R1204 B.n301 B.n300 10.6151
R1205 B.n301 B.n168 10.6151
R1206 B.n305 B.n168 10.6151
R1207 B.n306 B.n305 10.6151
R1208 B.n307 B.n306 10.6151
R1209 B.n307 B.n166 10.6151
R1210 B.n311 B.n166 10.6151
R1211 B.n312 B.n311 10.6151
R1212 B.n313 B.n312 10.6151
R1213 B.n313 B.n164 10.6151
R1214 B.n317 B.n164 10.6151
R1215 B.n318 B.n317 10.6151
R1216 B.n319 B.n318 10.6151
R1217 B.n319 B.n162 10.6151
R1218 B.n323 B.n162 10.6151
R1219 B.n324 B.n323 10.6151
R1220 B.n325 B.n324 10.6151
R1221 B.n325 B.n160 10.6151
R1222 B.n329 B.n160 10.6151
R1223 B.n330 B.n329 10.6151
R1224 B.n331 B.n330 10.6151
R1225 B.n331 B.n158 10.6151
R1226 B.n335 B.n158 10.6151
R1227 B.n336 B.n335 10.6151
R1228 B.n338 B.n154 10.6151
R1229 B.n342 B.n154 10.6151
R1230 B.n343 B.n342 10.6151
R1231 B.n344 B.n343 10.6151
R1232 B.n344 B.n152 10.6151
R1233 B.n348 B.n152 10.6151
R1234 B.n349 B.n348 10.6151
R1235 B.n350 B.n349 10.6151
R1236 B.n354 B.n353 10.6151
R1237 B.n355 B.n354 10.6151
R1238 B.n355 B.n146 10.6151
R1239 B.n359 B.n146 10.6151
R1240 B.n360 B.n359 10.6151
R1241 B.n361 B.n360 10.6151
R1242 B.n361 B.n144 10.6151
R1243 B.n365 B.n144 10.6151
R1244 B.n366 B.n365 10.6151
R1245 B.n367 B.n366 10.6151
R1246 B.n367 B.n142 10.6151
R1247 B.n371 B.n142 10.6151
R1248 B.n372 B.n371 10.6151
R1249 B.n373 B.n372 10.6151
R1250 B.n373 B.n140 10.6151
R1251 B.n377 B.n140 10.6151
R1252 B.n378 B.n377 10.6151
R1253 B.n379 B.n378 10.6151
R1254 B.n379 B.n138 10.6151
R1255 B.n383 B.n138 10.6151
R1256 B.n384 B.n383 10.6151
R1257 B.n385 B.n384 10.6151
R1258 B.n385 B.n136 10.6151
R1259 B.n389 B.n136 10.6151
R1260 B.n390 B.n389 10.6151
R1261 B.n391 B.n390 10.6151
R1262 B.n391 B.n134 10.6151
R1263 B.n395 B.n134 10.6151
R1264 B.n396 B.n395 10.6151
R1265 B.n397 B.n396 10.6151
R1266 B.n397 B.n132 10.6151
R1267 B.n401 B.n132 10.6151
R1268 B.n402 B.n401 10.6151
R1269 B.n403 B.n402 10.6151
R1270 B.n403 B.n130 10.6151
R1271 B.n407 B.n130 10.6151
R1272 B.n408 B.n407 10.6151
R1273 B.n409 B.n408 10.6151
R1274 B.n409 B.n128 10.6151
R1275 B.n413 B.n128 10.6151
R1276 B.n414 B.n413 10.6151
R1277 B.n415 B.n414 10.6151
R1278 B.n415 B.n126 10.6151
R1279 B.n419 B.n126 10.6151
R1280 B.n420 B.n419 10.6151
R1281 B.n421 B.n420 10.6151
R1282 B.n421 B.n124 10.6151
R1283 B.n425 B.n124 10.6151
R1284 B.n426 B.n425 10.6151
R1285 B.n427 B.n426 10.6151
R1286 B.n427 B.n122 10.6151
R1287 B.n431 B.n122 10.6151
R1288 B.n432 B.n431 10.6151
R1289 B.n433 B.n432 10.6151
R1290 B.n433 B.n120 10.6151
R1291 B.n437 B.n120 10.6151
R1292 B.n438 B.n437 10.6151
R1293 B.n439 B.n438 10.6151
R1294 B.n439 B.n118 10.6151
R1295 B.n443 B.n118 10.6151
R1296 B.n444 B.n443 10.6151
R1297 B.n445 B.n444 10.6151
R1298 B.n445 B.n116 10.6151
R1299 B.n449 B.n116 10.6151
R1300 B.n239 B.n190 10.6151
R1301 B.n235 B.n190 10.6151
R1302 B.n235 B.n234 10.6151
R1303 B.n234 B.n233 10.6151
R1304 B.n233 B.n192 10.6151
R1305 B.n229 B.n192 10.6151
R1306 B.n229 B.n228 10.6151
R1307 B.n228 B.n227 10.6151
R1308 B.n227 B.n194 10.6151
R1309 B.n223 B.n194 10.6151
R1310 B.n223 B.n222 10.6151
R1311 B.n222 B.n221 10.6151
R1312 B.n221 B.n196 10.6151
R1313 B.n217 B.n196 10.6151
R1314 B.n217 B.n216 10.6151
R1315 B.n216 B.n215 10.6151
R1316 B.n215 B.n198 10.6151
R1317 B.n211 B.n198 10.6151
R1318 B.n211 B.n210 10.6151
R1319 B.n210 B.n209 10.6151
R1320 B.n209 B.n200 10.6151
R1321 B.n205 B.n200 10.6151
R1322 B.n205 B.n204 10.6151
R1323 B.n204 B.n203 10.6151
R1324 B.n203 B.n0 10.6151
R1325 B.n775 B.n1 10.6151
R1326 B.n775 B.n774 10.6151
R1327 B.n774 B.n773 10.6151
R1328 B.n773 B.n4 10.6151
R1329 B.n769 B.n4 10.6151
R1330 B.n769 B.n768 10.6151
R1331 B.n768 B.n767 10.6151
R1332 B.n767 B.n6 10.6151
R1333 B.n763 B.n6 10.6151
R1334 B.n763 B.n762 10.6151
R1335 B.n762 B.n761 10.6151
R1336 B.n761 B.n8 10.6151
R1337 B.n757 B.n8 10.6151
R1338 B.n757 B.n756 10.6151
R1339 B.n756 B.n755 10.6151
R1340 B.n755 B.n10 10.6151
R1341 B.n751 B.n10 10.6151
R1342 B.n751 B.n750 10.6151
R1343 B.n750 B.n749 10.6151
R1344 B.n749 B.n12 10.6151
R1345 B.n745 B.n12 10.6151
R1346 B.n745 B.n744 10.6151
R1347 B.n744 B.n743 10.6151
R1348 B.n743 B.n14 10.6151
R1349 B.n739 B.n14 10.6151
R1350 B.n641 B.n640 6.5566
R1351 B.n628 B.n56 6.5566
R1352 B.n338 B.n337 6.5566
R1353 B.n350 B.n150 6.5566
R1354 B.n642 B.n641 4.05904
R1355 B.n625 B.n56 4.05904
R1356 B.n337 B.n336 4.05904
R1357 B.n353 B.n150 4.05904
R1358 B.n779 B.n0 2.81026
R1359 B.n779 B.n1 2.81026
C0 B w_n2206_n4936# 9.55223f
C1 B VDD1 2.27387f
C2 w_n2206_n4936# VTAIL 4.21113f
C3 VDD1 VTAIL 21.8516f
C4 w_n2206_n4936# VN 4.29107f
C5 VP w_n2206_n4936# 4.57242f
C6 VDD1 VN 0.148983f
C7 VP VDD1 10.972401f
C8 B VTAIL 4.1292f
C9 w_n2206_n4936# VDD2 2.65805f
C10 B VN 0.892694f
C11 VP B 1.35531f
C12 VDD2 VDD1 0.972099f
C13 B VDD2 2.31815f
C14 VN VTAIL 10.323501f
C15 VP VTAIL 10.3385f
C16 VP VN 7.04646f
C17 w_n2206_n4936# VDD1 2.61344f
C18 VDD2 VTAIL 21.881401f
C19 VDD2 VN 10.786099f
C20 VP VDD2 0.342736f
C21 VDD2 VSUBS 1.755595f
C22 VDD1 VSUBS 1.413576f
C23 VTAIL VSUBS 0.988596f
C24 VN VSUBS 5.53811f
C25 VP VSUBS 2.108855f
C26 B VSUBS 3.675884f
C27 w_n2206_n4936# VSUBS 0.132969p
C28 B.n0 VSUBS 0.005658f
C29 B.n1 VSUBS 0.005658f
C30 B.n2 VSUBS 0.008948f
C31 B.n3 VSUBS 0.008948f
C32 B.n4 VSUBS 0.008948f
C33 B.n5 VSUBS 0.008948f
C34 B.n6 VSUBS 0.008948f
C35 B.n7 VSUBS 0.008948f
C36 B.n8 VSUBS 0.008948f
C37 B.n9 VSUBS 0.008948f
C38 B.n10 VSUBS 0.008948f
C39 B.n11 VSUBS 0.008948f
C40 B.n12 VSUBS 0.008948f
C41 B.n13 VSUBS 0.008948f
C42 B.n14 VSUBS 0.008948f
C43 B.n15 VSUBS 0.022707f
C44 B.n16 VSUBS 0.008948f
C45 B.n17 VSUBS 0.008948f
C46 B.n18 VSUBS 0.008948f
C47 B.n19 VSUBS 0.008948f
C48 B.n20 VSUBS 0.008948f
C49 B.n21 VSUBS 0.008948f
C50 B.n22 VSUBS 0.008948f
C51 B.n23 VSUBS 0.008948f
C52 B.n24 VSUBS 0.008948f
C53 B.n25 VSUBS 0.008948f
C54 B.n26 VSUBS 0.008948f
C55 B.n27 VSUBS 0.008948f
C56 B.n28 VSUBS 0.008948f
C57 B.n29 VSUBS 0.008948f
C58 B.n30 VSUBS 0.008948f
C59 B.n31 VSUBS 0.008948f
C60 B.n32 VSUBS 0.008948f
C61 B.n33 VSUBS 0.008948f
C62 B.n34 VSUBS 0.008948f
C63 B.n35 VSUBS 0.008948f
C64 B.n36 VSUBS 0.008948f
C65 B.n37 VSUBS 0.008948f
C66 B.n38 VSUBS 0.008948f
C67 B.n39 VSUBS 0.008948f
C68 B.n40 VSUBS 0.008948f
C69 B.n41 VSUBS 0.008948f
C70 B.n42 VSUBS 0.008948f
C71 B.n43 VSUBS 0.008948f
C72 B.n44 VSUBS 0.008948f
C73 B.n45 VSUBS 0.008948f
C74 B.n46 VSUBS 0.008948f
C75 B.n47 VSUBS 0.008948f
C76 B.t2 VSUBS 0.861755f
C77 B.t1 VSUBS 0.872566f
C78 B.t0 VSUBS 0.712146f
C79 B.n48 VSUBS 0.255875f
C80 B.n49 VSUBS 0.082212f
C81 B.n50 VSUBS 0.008948f
C82 B.n51 VSUBS 0.008948f
C83 B.n52 VSUBS 0.008948f
C84 B.n53 VSUBS 0.008948f
C85 B.t11 VSUBS 0.861718f
C86 B.t10 VSUBS 0.872533f
C87 B.t9 VSUBS 0.712146f
C88 B.n54 VSUBS 0.255909f
C89 B.n55 VSUBS 0.082249f
C90 B.n56 VSUBS 0.020732f
C91 B.n57 VSUBS 0.008948f
C92 B.n58 VSUBS 0.008948f
C93 B.n59 VSUBS 0.008948f
C94 B.n60 VSUBS 0.008948f
C95 B.n61 VSUBS 0.008948f
C96 B.n62 VSUBS 0.008948f
C97 B.n63 VSUBS 0.008948f
C98 B.n64 VSUBS 0.008948f
C99 B.n65 VSUBS 0.008948f
C100 B.n66 VSUBS 0.008948f
C101 B.n67 VSUBS 0.008948f
C102 B.n68 VSUBS 0.008948f
C103 B.n69 VSUBS 0.008948f
C104 B.n70 VSUBS 0.008948f
C105 B.n71 VSUBS 0.008948f
C106 B.n72 VSUBS 0.008948f
C107 B.n73 VSUBS 0.008948f
C108 B.n74 VSUBS 0.008948f
C109 B.n75 VSUBS 0.008948f
C110 B.n76 VSUBS 0.008948f
C111 B.n77 VSUBS 0.008948f
C112 B.n78 VSUBS 0.008948f
C113 B.n79 VSUBS 0.008948f
C114 B.n80 VSUBS 0.008948f
C115 B.n81 VSUBS 0.008948f
C116 B.n82 VSUBS 0.008948f
C117 B.n83 VSUBS 0.008948f
C118 B.n84 VSUBS 0.008948f
C119 B.n85 VSUBS 0.008948f
C120 B.n86 VSUBS 0.008948f
C121 B.n87 VSUBS 0.008948f
C122 B.n88 VSUBS 0.008948f
C123 B.n89 VSUBS 0.021244f
C124 B.n90 VSUBS 0.008948f
C125 B.n91 VSUBS 0.008948f
C126 B.n92 VSUBS 0.008948f
C127 B.n93 VSUBS 0.008948f
C128 B.n94 VSUBS 0.008948f
C129 B.n95 VSUBS 0.008948f
C130 B.n96 VSUBS 0.008948f
C131 B.n97 VSUBS 0.008948f
C132 B.n98 VSUBS 0.008948f
C133 B.n99 VSUBS 0.008948f
C134 B.n100 VSUBS 0.008948f
C135 B.n101 VSUBS 0.008948f
C136 B.n102 VSUBS 0.008948f
C137 B.n103 VSUBS 0.008948f
C138 B.n104 VSUBS 0.008948f
C139 B.n105 VSUBS 0.008948f
C140 B.n106 VSUBS 0.008948f
C141 B.n107 VSUBS 0.008948f
C142 B.n108 VSUBS 0.008948f
C143 B.n109 VSUBS 0.008948f
C144 B.n110 VSUBS 0.008948f
C145 B.n111 VSUBS 0.008948f
C146 B.n112 VSUBS 0.008948f
C147 B.n113 VSUBS 0.008948f
C148 B.n114 VSUBS 0.008948f
C149 B.n115 VSUBS 0.021244f
C150 B.n116 VSUBS 0.008948f
C151 B.n117 VSUBS 0.008948f
C152 B.n118 VSUBS 0.008948f
C153 B.n119 VSUBS 0.008948f
C154 B.n120 VSUBS 0.008948f
C155 B.n121 VSUBS 0.008948f
C156 B.n122 VSUBS 0.008948f
C157 B.n123 VSUBS 0.008948f
C158 B.n124 VSUBS 0.008948f
C159 B.n125 VSUBS 0.008948f
C160 B.n126 VSUBS 0.008948f
C161 B.n127 VSUBS 0.008948f
C162 B.n128 VSUBS 0.008948f
C163 B.n129 VSUBS 0.008948f
C164 B.n130 VSUBS 0.008948f
C165 B.n131 VSUBS 0.008948f
C166 B.n132 VSUBS 0.008948f
C167 B.n133 VSUBS 0.008948f
C168 B.n134 VSUBS 0.008948f
C169 B.n135 VSUBS 0.008948f
C170 B.n136 VSUBS 0.008948f
C171 B.n137 VSUBS 0.008948f
C172 B.n138 VSUBS 0.008948f
C173 B.n139 VSUBS 0.008948f
C174 B.n140 VSUBS 0.008948f
C175 B.n141 VSUBS 0.008948f
C176 B.n142 VSUBS 0.008948f
C177 B.n143 VSUBS 0.008948f
C178 B.n144 VSUBS 0.008948f
C179 B.n145 VSUBS 0.008948f
C180 B.n146 VSUBS 0.008948f
C181 B.n147 VSUBS 0.008948f
C182 B.t7 VSUBS 0.861718f
C183 B.t8 VSUBS 0.872533f
C184 B.t6 VSUBS 0.712146f
C185 B.n148 VSUBS 0.255909f
C186 B.n149 VSUBS 0.082249f
C187 B.n150 VSUBS 0.020732f
C188 B.n151 VSUBS 0.008948f
C189 B.n152 VSUBS 0.008948f
C190 B.n153 VSUBS 0.008948f
C191 B.n154 VSUBS 0.008948f
C192 B.n155 VSUBS 0.008948f
C193 B.t4 VSUBS 0.861755f
C194 B.t5 VSUBS 0.872566f
C195 B.t3 VSUBS 0.712146f
C196 B.n156 VSUBS 0.255875f
C197 B.n157 VSUBS 0.082212f
C198 B.n158 VSUBS 0.008948f
C199 B.n159 VSUBS 0.008948f
C200 B.n160 VSUBS 0.008948f
C201 B.n161 VSUBS 0.008948f
C202 B.n162 VSUBS 0.008948f
C203 B.n163 VSUBS 0.008948f
C204 B.n164 VSUBS 0.008948f
C205 B.n165 VSUBS 0.008948f
C206 B.n166 VSUBS 0.008948f
C207 B.n167 VSUBS 0.008948f
C208 B.n168 VSUBS 0.008948f
C209 B.n169 VSUBS 0.008948f
C210 B.n170 VSUBS 0.008948f
C211 B.n171 VSUBS 0.008948f
C212 B.n172 VSUBS 0.008948f
C213 B.n173 VSUBS 0.008948f
C214 B.n174 VSUBS 0.008948f
C215 B.n175 VSUBS 0.008948f
C216 B.n176 VSUBS 0.008948f
C217 B.n177 VSUBS 0.008948f
C218 B.n178 VSUBS 0.008948f
C219 B.n179 VSUBS 0.008948f
C220 B.n180 VSUBS 0.008948f
C221 B.n181 VSUBS 0.008948f
C222 B.n182 VSUBS 0.008948f
C223 B.n183 VSUBS 0.008948f
C224 B.n184 VSUBS 0.008948f
C225 B.n185 VSUBS 0.008948f
C226 B.n186 VSUBS 0.008948f
C227 B.n187 VSUBS 0.008948f
C228 B.n188 VSUBS 0.008948f
C229 B.n189 VSUBS 0.022707f
C230 B.n190 VSUBS 0.008948f
C231 B.n191 VSUBS 0.008948f
C232 B.n192 VSUBS 0.008948f
C233 B.n193 VSUBS 0.008948f
C234 B.n194 VSUBS 0.008948f
C235 B.n195 VSUBS 0.008948f
C236 B.n196 VSUBS 0.008948f
C237 B.n197 VSUBS 0.008948f
C238 B.n198 VSUBS 0.008948f
C239 B.n199 VSUBS 0.008948f
C240 B.n200 VSUBS 0.008948f
C241 B.n201 VSUBS 0.008948f
C242 B.n202 VSUBS 0.008948f
C243 B.n203 VSUBS 0.008948f
C244 B.n204 VSUBS 0.008948f
C245 B.n205 VSUBS 0.008948f
C246 B.n206 VSUBS 0.008948f
C247 B.n207 VSUBS 0.008948f
C248 B.n208 VSUBS 0.008948f
C249 B.n209 VSUBS 0.008948f
C250 B.n210 VSUBS 0.008948f
C251 B.n211 VSUBS 0.008948f
C252 B.n212 VSUBS 0.008948f
C253 B.n213 VSUBS 0.008948f
C254 B.n214 VSUBS 0.008948f
C255 B.n215 VSUBS 0.008948f
C256 B.n216 VSUBS 0.008948f
C257 B.n217 VSUBS 0.008948f
C258 B.n218 VSUBS 0.008948f
C259 B.n219 VSUBS 0.008948f
C260 B.n220 VSUBS 0.008948f
C261 B.n221 VSUBS 0.008948f
C262 B.n222 VSUBS 0.008948f
C263 B.n223 VSUBS 0.008948f
C264 B.n224 VSUBS 0.008948f
C265 B.n225 VSUBS 0.008948f
C266 B.n226 VSUBS 0.008948f
C267 B.n227 VSUBS 0.008948f
C268 B.n228 VSUBS 0.008948f
C269 B.n229 VSUBS 0.008948f
C270 B.n230 VSUBS 0.008948f
C271 B.n231 VSUBS 0.008948f
C272 B.n232 VSUBS 0.008948f
C273 B.n233 VSUBS 0.008948f
C274 B.n234 VSUBS 0.008948f
C275 B.n235 VSUBS 0.008948f
C276 B.n236 VSUBS 0.008948f
C277 B.n237 VSUBS 0.008948f
C278 B.n238 VSUBS 0.021244f
C279 B.n239 VSUBS 0.021244f
C280 B.n240 VSUBS 0.022707f
C281 B.n241 VSUBS 0.008948f
C282 B.n242 VSUBS 0.008948f
C283 B.n243 VSUBS 0.008948f
C284 B.n244 VSUBS 0.008948f
C285 B.n245 VSUBS 0.008948f
C286 B.n246 VSUBS 0.008948f
C287 B.n247 VSUBS 0.008948f
C288 B.n248 VSUBS 0.008948f
C289 B.n249 VSUBS 0.008948f
C290 B.n250 VSUBS 0.008948f
C291 B.n251 VSUBS 0.008948f
C292 B.n252 VSUBS 0.008948f
C293 B.n253 VSUBS 0.008948f
C294 B.n254 VSUBS 0.008948f
C295 B.n255 VSUBS 0.008948f
C296 B.n256 VSUBS 0.008948f
C297 B.n257 VSUBS 0.008948f
C298 B.n258 VSUBS 0.008948f
C299 B.n259 VSUBS 0.008948f
C300 B.n260 VSUBS 0.008948f
C301 B.n261 VSUBS 0.008948f
C302 B.n262 VSUBS 0.008948f
C303 B.n263 VSUBS 0.008948f
C304 B.n264 VSUBS 0.008948f
C305 B.n265 VSUBS 0.008948f
C306 B.n266 VSUBS 0.008948f
C307 B.n267 VSUBS 0.008948f
C308 B.n268 VSUBS 0.008948f
C309 B.n269 VSUBS 0.008948f
C310 B.n270 VSUBS 0.008948f
C311 B.n271 VSUBS 0.008948f
C312 B.n272 VSUBS 0.008948f
C313 B.n273 VSUBS 0.008948f
C314 B.n274 VSUBS 0.008948f
C315 B.n275 VSUBS 0.008948f
C316 B.n276 VSUBS 0.008948f
C317 B.n277 VSUBS 0.008948f
C318 B.n278 VSUBS 0.008948f
C319 B.n279 VSUBS 0.008948f
C320 B.n280 VSUBS 0.008948f
C321 B.n281 VSUBS 0.008948f
C322 B.n282 VSUBS 0.008948f
C323 B.n283 VSUBS 0.008948f
C324 B.n284 VSUBS 0.008948f
C325 B.n285 VSUBS 0.008948f
C326 B.n286 VSUBS 0.008948f
C327 B.n287 VSUBS 0.008948f
C328 B.n288 VSUBS 0.008948f
C329 B.n289 VSUBS 0.008948f
C330 B.n290 VSUBS 0.008948f
C331 B.n291 VSUBS 0.008948f
C332 B.n292 VSUBS 0.008948f
C333 B.n293 VSUBS 0.008948f
C334 B.n294 VSUBS 0.008948f
C335 B.n295 VSUBS 0.008948f
C336 B.n296 VSUBS 0.008948f
C337 B.n297 VSUBS 0.008948f
C338 B.n298 VSUBS 0.008948f
C339 B.n299 VSUBS 0.008948f
C340 B.n300 VSUBS 0.008948f
C341 B.n301 VSUBS 0.008948f
C342 B.n302 VSUBS 0.008948f
C343 B.n303 VSUBS 0.008948f
C344 B.n304 VSUBS 0.008948f
C345 B.n305 VSUBS 0.008948f
C346 B.n306 VSUBS 0.008948f
C347 B.n307 VSUBS 0.008948f
C348 B.n308 VSUBS 0.008948f
C349 B.n309 VSUBS 0.008948f
C350 B.n310 VSUBS 0.008948f
C351 B.n311 VSUBS 0.008948f
C352 B.n312 VSUBS 0.008948f
C353 B.n313 VSUBS 0.008948f
C354 B.n314 VSUBS 0.008948f
C355 B.n315 VSUBS 0.008948f
C356 B.n316 VSUBS 0.008948f
C357 B.n317 VSUBS 0.008948f
C358 B.n318 VSUBS 0.008948f
C359 B.n319 VSUBS 0.008948f
C360 B.n320 VSUBS 0.008948f
C361 B.n321 VSUBS 0.008948f
C362 B.n322 VSUBS 0.008948f
C363 B.n323 VSUBS 0.008948f
C364 B.n324 VSUBS 0.008948f
C365 B.n325 VSUBS 0.008948f
C366 B.n326 VSUBS 0.008948f
C367 B.n327 VSUBS 0.008948f
C368 B.n328 VSUBS 0.008948f
C369 B.n329 VSUBS 0.008948f
C370 B.n330 VSUBS 0.008948f
C371 B.n331 VSUBS 0.008948f
C372 B.n332 VSUBS 0.008948f
C373 B.n333 VSUBS 0.008948f
C374 B.n334 VSUBS 0.008948f
C375 B.n335 VSUBS 0.008948f
C376 B.n336 VSUBS 0.006185f
C377 B.n337 VSUBS 0.020732f
C378 B.n338 VSUBS 0.007238f
C379 B.n339 VSUBS 0.008948f
C380 B.n340 VSUBS 0.008948f
C381 B.n341 VSUBS 0.008948f
C382 B.n342 VSUBS 0.008948f
C383 B.n343 VSUBS 0.008948f
C384 B.n344 VSUBS 0.008948f
C385 B.n345 VSUBS 0.008948f
C386 B.n346 VSUBS 0.008948f
C387 B.n347 VSUBS 0.008948f
C388 B.n348 VSUBS 0.008948f
C389 B.n349 VSUBS 0.008948f
C390 B.n350 VSUBS 0.007238f
C391 B.n351 VSUBS 0.008948f
C392 B.n352 VSUBS 0.008948f
C393 B.n353 VSUBS 0.006185f
C394 B.n354 VSUBS 0.008948f
C395 B.n355 VSUBS 0.008948f
C396 B.n356 VSUBS 0.008948f
C397 B.n357 VSUBS 0.008948f
C398 B.n358 VSUBS 0.008948f
C399 B.n359 VSUBS 0.008948f
C400 B.n360 VSUBS 0.008948f
C401 B.n361 VSUBS 0.008948f
C402 B.n362 VSUBS 0.008948f
C403 B.n363 VSUBS 0.008948f
C404 B.n364 VSUBS 0.008948f
C405 B.n365 VSUBS 0.008948f
C406 B.n366 VSUBS 0.008948f
C407 B.n367 VSUBS 0.008948f
C408 B.n368 VSUBS 0.008948f
C409 B.n369 VSUBS 0.008948f
C410 B.n370 VSUBS 0.008948f
C411 B.n371 VSUBS 0.008948f
C412 B.n372 VSUBS 0.008948f
C413 B.n373 VSUBS 0.008948f
C414 B.n374 VSUBS 0.008948f
C415 B.n375 VSUBS 0.008948f
C416 B.n376 VSUBS 0.008948f
C417 B.n377 VSUBS 0.008948f
C418 B.n378 VSUBS 0.008948f
C419 B.n379 VSUBS 0.008948f
C420 B.n380 VSUBS 0.008948f
C421 B.n381 VSUBS 0.008948f
C422 B.n382 VSUBS 0.008948f
C423 B.n383 VSUBS 0.008948f
C424 B.n384 VSUBS 0.008948f
C425 B.n385 VSUBS 0.008948f
C426 B.n386 VSUBS 0.008948f
C427 B.n387 VSUBS 0.008948f
C428 B.n388 VSUBS 0.008948f
C429 B.n389 VSUBS 0.008948f
C430 B.n390 VSUBS 0.008948f
C431 B.n391 VSUBS 0.008948f
C432 B.n392 VSUBS 0.008948f
C433 B.n393 VSUBS 0.008948f
C434 B.n394 VSUBS 0.008948f
C435 B.n395 VSUBS 0.008948f
C436 B.n396 VSUBS 0.008948f
C437 B.n397 VSUBS 0.008948f
C438 B.n398 VSUBS 0.008948f
C439 B.n399 VSUBS 0.008948f
C440 B.n400 VSUBS 0.008948f
C441 B.n401 VSUBS 0.008948f
C442 B.n402 VSUBS 0.008948f
C443 B.n403 VSUBS 0.008948f
C444 B.n404 VSUBS 0.008948f
C445 B.n405 VSUBS 0.008948f
C446 B.n406 VSUBS 0.008948f
C447 B.n407 VSUBS 0.008948f
C448 B.n408 VSUBS 0.008948f
C449 B.n409 VSUBS 0.008948f
C450 B.n410 VSUBS 0.008948f
C451 B.n411 VSUBS 0.008948f
C452 B.n412 VSUBS 0.008948f
C453 B.n413 VSUBS 0.008948f
C454 B.n414 VSUBS 0.008948f
C455 B.n415 VSUBS 0.008948f
C456 B.n416 VSUBS 0.008948f
C457 B.n417 VSUBS 0.008948f
C458 B.n418 VSUBS 0.008948f
C459 B.n419 VSUBS 0.008948f
C460 B.n420 VSUBS 0.008948f
C461 B.n421 VSUBS 0.008948f
C462 B.n422 VSUBS 0.008948f
C463 B.n423 VSUBS 0.008948f
C464 B.n424 VSUBS 0.008948f
C465 B.n425 VSUBS 0.008948f
C466 B.n426 VSUBS 0.008948f
C467 B.n427 VSUBS 0.008948f
C468 B.n428 VSUBS 0.008948f
C469 B.n429 VSUBS 0.008948f
C470 B.n430 VSUBS 0.008948f
C471 B.n431 VSUBS 0.008948f
C472 B.n432 VSUBS 0.008948f
C473 B.n433 VSUBS 0.008948f
C474 B.n434 VSUBS 0.008948f
C475 B.n435 VSUBS 0.008948f
C476 B.n436 VSUBS 0.008948f
C477 B.n437 VSUBS 0.008948f
C478 B.n438 VSUBS 0.008948f
C479 B.n439 VSUBS 0.008948f
C480 B.n440 VSUBS 0.008948f
C481 B.n441 VSUBS 0.008948f
C482 B.n442 VSUBS 0.008948f
C483 B.n443 VSUBS 0.008948f
C484 B.n444 VSUBS 0.008948f
C485 B.n445 VSUBS 0.008948f
C486 B.n446 VSUBS 0.008948f
C487 B.n447 VSUBS 0.008948f
C488 B.n448 VSUBS 0.022707f
C489 B.n449 VSUBS 0.022707f
C490 B.n450 VSUBS 0.021244f
C491 B.n451 VSUBS 0.008948f
C492 B.n452 VSUBS 0.008948f
C493 B.n453 VSUBS 0.008948f
C494 B.n454 VSUBS 0.008948f
C495 B.n455 VSUBS 0.008948f
C496 B.n456 VSUBS 0.008948f
C497 B.n457 VSUBS 0.008948f
C498 B.n458 VSUBS 0.008948f
C499 B.n459 VSUBS 0.008948f
C500 B.n460 VSUBS 0.008948f
C501 B.n461 VSUBS 0.008948f
C502 B.n462 VSUBS 0.008948f
C503 B.n463 VSUBS 0.008948f
C504 B.n464 VSUBS 0.008948f
C505 B.n465 VSUBS 0.008948f
C506 B.n466 VSUBS 0.008948f
C507 B.n467 VSUBS 0.008948f
C508 B.n468 VSUBS 0.008948f
C509 B.n469 VSUBS 0.008948f
C510 B.n470 VSUBS 0.008948f
C511 B.n471 VSUBS 0.008948f
C512 B.n472 VSUBS 0.008948f
C513 B.n473 VSUBS 0.008948f
C514 B.n474 VSUBS 0.008948f
C515 B.n475 VSUBS 0.008948f
C516 B.n476 VSUBS 0.008948f
C517 B.n477 VSUBS 0.008948f
C518 B.n478 VSUBS 0.008948f
C519 B.n479 VSUBS 0.008948f
C520 B.n480 VSUBS 0.008948f
C521 B.n481 VSUBS 0.008948f
C522 B.n482 VSUBS 0.008948f
C523 B.n483 VSUBS 0.008948f
C524 B.n484 VSUBS 0.008948f
C525 B.n485 VSUBS 0.008948f
C526 B.n486 VSUBS 0.008948f
C527 B.n487 VSUBS 0.008948f
C528 B.n488 VSUBS 0.008948f
C529 B.n489 VSUBS 0.008948f
C530 B.n490 VSUBS 0.008948f
C531 B.n491 VSUBS 0.008948f
C532 B.n492 VSUBS 0.008948f
C533 B.n493 VSUBS 0.008948f
C534 B.n494 VSUBS 0.008948f
C535 B.n495 VSUBS 0.008948f
C536 B.n496 VSUBS 0.008948f
C537 B.n497 VSUBS 0.008948f
C538 B.n498 VSUBS 0.008948f
C539 B.n499 VSUBS 0.008948f
C540 B.n500 VSUBS 0.008948f
C541 B.n501 VSUBS 0.008948f
C542 B.n502 VSUBS 0.008948f
C543 B.n503 VSUBS 0.008948f
C544 B.n504 VSUBS 0.008948f
C545 B.n505 VSUBS 0.008948f
C546 B.n506 VSUBS 0.008948f
C547 B.n507 VSUBS 0.008948f
C548 B.n508 VSUBS 0.008948f
C549 B.n509 VSUBS 0.008948f
C550 B.n510 VSUBS 0.008948f
C551 B.n511 VSUBS 0.008948f
C552 B.n512 VSUBS 0.008948f
C553 B.n513 VSUBS 0.008948f
C554 B.n514 VSUBS 0.008948f
C555 B.n515 VSUBS 0.008948f
C556 B.n516 VSUBS 0.008948f
C557 B.n517 VSUBS 0.008948f
C558 B.n518 VSUBS 0.008948f
C559 B.n519 VSUBS 0.008948f
C560 B.n520 VSUBS 0.008948f
C561 B.n521 VSUBS 0.008948f
C562 B.n522 VSUBS 0.008948f
C563 B.n523 VSUBS 0.008948f
C564 B.n524 VSUBS 0.008948f
C565 B.n525 VSUBS 0.008948f
C566 B.n526 VSUBS 0.008948f
C567 B.n527 VSUBS 0.008948f
C568 B.n528 VSUBS 0.022228f
C569 B.n529 VSUBS 0.021724f
C570 B.n530 VSUBS 0.022707f
C571 B.n531 VSUBS 0.008948f
C572 B.n532 VSUBS 0.008948f
C573 B.n533 VSUBS 0.008948f
C574 B.n534 VSUBS 0.008948f
C575 B.n535 VSUBS 0.008948f
C576 B.n536 VSUBS 0.008948f
C577 B.n537 VSUBS 0.008948f
C578 B.n538 VSUBS 0.008948f
C579 B.n539 VSUBS 0.008948f
C580 B.n540 VSUBS 0.008948f
C581 B.n541 VSUBS 0.008948f
C582 B.n542 VSUBS 0.008948f
C583 B.n543 VSUBS 0.008948f
C584 B.n544 VSUBS 0.008948f
C585 B.n545 VSUBS 0.008948f
C586 B.n546 VSUBS 0.008948f
C587 B.n547 VSUBS 0.008948f
C588 B.n548 VSUBS 0.008948f
C589 B.n549 VSUBS 0.008948f
C590 B.n550 VSUBS 0.008948f
C591 B.n551 VSUBS 0.008948f
C592 B.n552 VSUBS 0.008948f
C593 B.n553 VSUBS 0.008948f
C594 B.n554 VSUBS 0.008948f
C595 B.n555 VSUBS 0.008948f
C596 B.n556 VSUBS 0.008948f
C597 B.n557 VSUBS 0.008948f
C598 B.n558 VSUBS 0.008948f
C599 B.n559 VSUBS 0.008948f
C600 B.n560 VSUBS 0.008948f
C601 B.n561 VSUBS 0.008948f
C602 B.n562 VSUBS 0.008948f
C603 B.n563 VSUBS 0.008948f
C604 B.n564 VSUBS 0.008948f
C605 B.n565 VSUBS 0.008948f
C606 B.n566 VSUBS 0.008948f
C607 B.n567 VSUBS 0.008948f
C608 B.n568 VSUBS 0.008948f
C609 B.n569 VSUBS 0.008948f
C610 B.n570 VSUBS 0.008948f
C611 B.n571 VSUBS 0.008948f
C612 B.n572 VSUBS 0.008948f
C613 B.n573 VSUBS 0.008948f
C614 B.n574 VSUBS 0.008948f
C615 B.n575 VSUBS 0.008948f
C616 B.n576 VSUBS 0.008948f
C617 B.n577 VSUBS 0.008948f
C618 B.n578 VSUBS 0.008948f
C619 B.n579 VSUBS 0.008948f
C620 B.n580 VSUBS 0.008948f
C621 B.n581 VSUBS 0.008948f
C622 B.n582 VSUBS 0.008948f
C623 B.n583 VSUBS 0.008948f
C624 B.n584 VSUBS 0.008948f
C625 B.n585 VSUBS 0.008948f
C626 B.n586 VSUBS 0.008948f
C627 B.n587 VSUBS 0.008948f
C628 B.n588 VSUBS 0.008948f
C629 B.n589 VSUBS 0.008948f
C630 B.n590 VSUBS 0.008948f
C631 B.n591 VSUBS 0.008948f
C632 B.n592 VSUBS 0.008948f
C633 B.n593 VSUBS 0.008948f
C634 B.n594 VSUBS 0.008948f
C635 B.n595 VSUBS 0.008948f
C636 B.n596 VSUBS 0.008948f
C637 B.n597 VSUBS 0.008948f
C638 B.n598 VSUBS 0.008948f
C639 B.n599 VSUBS 0.008948f
C640 B.n600 VSUBS 0.008948f
C641 B.n601 VSUBS 0.008948f
C642 B.n602 VSUBS 0.008948f
C643 B.n603 VSUBS 0.008948f
C644 B.n604 VSUBS 0.008948f
C645 B.n605 VSUBS 0.008948f
C646 B.n606 VSUBS 0.008948f
C647 B.n607 VSUBS 0.008948f
C648 B.n608 VSUBS 0.008948f
C649 B.n609 VSUBS 0.008948f
C650 B.n610 VSUBS 0.008948f
C651 B.n611 VSUBS 0.008948f
C652 B.n612 VSUBS 0.008948f
C653 B.n613 VSUBS 0.008948f
C654 B.n614 VSUBS 0.008948f
C655 B.n615 VSUBS 0.008948f
C656 B.n616 VSUBS 0.008948f
C657 B.n617 VSUBS 0.008948f
C658 B.n618 VSUBS 0.008948f
C659 B.n619 VSUBS 0.008948f
C660 B.n620 VSUBS 0.008948f
C661 B.n621 VSUBS 0.008948f
C662 B.n622 VSUBS 0.008948f
C663 B.n623 VSUBS 0.008948f
C664 B.n624 VSUBS 0.008948f
C665 B.n625 VSUBS 0.006185f
C666 B.n626 VSUBS 0.008948f
C667 B.n627 VSUBS 0.008948f
C668 B.n628 VSUBS 0.007238f
C669 B.n629 VSUBS 0.008948f
C670 B.n630 VSUBS 0.008948f
C671 B.n631 VSUBS 0.008948f
C672 B.n632 VSUBS 0.008948f
C673 B.n633 VSUBS 0.008948f
C674 B.n634 VSUBS 0.008948f
C675 B.n635 VSUBS 0.008948f
C676 B.n636 VSUBS 0.008948f
C677 B.n637 VSUBS 0.008948f
C678 B.n638 VSUBS 0.008948f
C679 B.n639 VSUBS 0.008948f
C680 B.n640 VSUBS 0.007238f
C681 B.n641 VSUBS 0.020732f
C682 B.n642 VSUBS 0.006185f
C683 B.n643 VSUBS 0.008948f
C684 B.n644 VSUBS 0.008948f
C685 B.n645 VSUBS 0.008948f
C686 B.n646 VSUBS 0.008948f
C687 B.n647 VSUBS 0.008948f
C688 B.n648 VSUBS 0.008948f
C689 B.n649 VSUBS 0.008948f
C690 B.n650 VSUBS 0.008948f
C691 B.n651 VSUBS 0.008948f
C692 B.n652 VSUBS 0.008948f
C693 B.n653 VSUBS 0.008948f
C694 B.n654 VSUBS 0.008948f
C695 B.n655 VSUBS 0.008948f
C696 B.n656 VSUBS 0.008948f
C697 B.n657 VSUBS 0.008948f
C698 B.n658 VSUBS 0.008948f
C699 B.n659 VSUBS 0.008948f
C700 B.n660 VSUBS 0.008948f
C701 B.n661 VSUBS 0.008948f
C702 B.n662 VSUBS 0.008948f
C703 B.n663 VSUBS 0.008948f
C704 B.n664 VSUBS 0.008948f
C705 B.n665 VSUBS 0.008948f
C706 B.n666 VSUBS 0.008948f
C707 B.n667 VSUBS 0.008948f
C708 B.n668 VSUBS 0.008948f
C709 B.n669 VSUBS 0.008948f
C710 B.n670 VSUBS 0.008948f
C711 B.n671 VSUBS 0.008948f
C712 B.n672 VSUBS 0.008948f
C713 B.n673 VSUBS 0.008948f
C714 B.n674 VSUBS 0.008948f
C715 B.n675 VSUBS 0.008948f
C716 B.n676 VSUBS 0.008948f
C717 B.n677 VSUBS 0.008948f
C718 B.n678 VSUBS 0.008948f
C719 B.n679 VSUBS 0.008948f
C720 B.n680 VSUBS 0.008948f
C721 B.n681 VSUBS 0.008948f
C722 B.n682 VSUBS 0.008948f
C723 B.n683 VSUBS 0.008948f
C724 B.n684 VSUBS 0.008948f
C725 B.n685 VSUBS 0.008948f
C726 B.n686 VSUBS 0.008948f
C727 B.n687 VSUBS 0.008948f
C728 B.n688 VSUBS 0.008948f
C729 B.n689 VSUBS 0.008948f
C730 B.n690 VSUBS 0.008948f
C731 B.n691 VSUBS 0.008948f
C732 B.n692 VSUBS 0.008948f
C733 B.n693 VSUBS 0.008948f
C734 B.n694 VSUBS 0.008948f
C735 B.n695 VSUBS 0.008948f
C736 B.n696 VSUBS 0.008948f
C737 B.n697 VSUBS 0.008948f
C738 B.n698 VSUBS 0.008948f
C739 B.n699 VSUBS 0.008948f
C740 B.n700 VSUBS 0.008948f
C741 B.n701 VSUBS 0.008948f
C742 B.n702 VSUBS 0.008948f
C743 B.n703 VSUBS 0.008948f
C744 B.n704 VSUBS 0.008948f
C745 B.n705 VSUBS 0.008948f
C746 B.n706 VSUBS 0.008948f
C747 B.n707 VSUBS 0.008948f
C748 B.n708 VSUBS 0.008948f
C749 B.n709 VSUBS 0.008948f
C750 B.n710 VSUBS 0.008948f
C751 B.n711 VSUBS 0.008948f
C752 B.n712 VSUBS 0.008948f
C753 B.n713 VSUBS 0.008948f
C754 B.n714 VSUBS 0.008948f
C755 B.n715 VSUBS 0.008948f
C756 B.n716 VSUBS 0.008948f
C757 B.n717 VSUBS 0.008948f
C758 B.n718 VSUBS 0.008948f
C759 B.n719 VSUBS 0.008948f
C760 B.n720 VSUBS 0.008948f
C761 B.n721 VSUBS 0.008948f
C762 B.n722 VSUBS 0.008948f
C763 B.n723 VSUBS 0.008948f
C764 B.n724 VSUBS 0.008948f
C765 B.n725 VSUBS 0.008948f
C766 B.n726 VSUBS 0.008948f
C767 B.n727 VSUBS 0.008948f
C768 B.n728 VSUBS 0.008948f
C769 B.n729 VSUBS 0.008948f
C770 B.n730 VSUBS 0.008948f
C771 B.n731 VSUBS 0.008948f
C772 B.n732 VSUBS 0.008948f
C773 B.n733 VSUBS 0.008948f
C774 B.n734 VSUBS 0.008948f
C775 B.n735 VSUBS 0.008948f
C776 B.n736 VSUBS 0.008948f
C777 B.n737 VSUBS 0.008948f
C778 B.n738 VSUBS 0.022707f
C779 B.n739 VSUBS 0.021244f
C780 B.n740 VSUBS 0.021244f
C781 B.n741 VSUBS 0.008948f
C782 B.n742 VSUBS 0.008948f
C783 B.n743 VSUBS 0.008948f
C784 B.n744 VSUBS 0.008948f
C785 B.n745 VSUBS 0.008948f
C786 B.n746 VSUBS 0.008948f
C787 B.n747 VSUBS 0.008948f
C788 B.n748 VSUBS 0.008948f
C789 B.n749 VSUBS 0.008948f
C790 B.n750 VSUBS 0.008948f
C791 B.n751 VSUBS 0.008948f
C792 B.n752 VSUBS 0.008948f
C793 B.n753 VSUBS 0.008948f
C794 B.n754 VSUBS 0.008948f
C795 B.n755 VSUBS 0.008948f
C796 B.n756 VSUBS 0.008948f
C797 B.n757 VSUBS 0.008948f
C798 B.n758 VSUBS 0.008948f
C799 B.n759 VSUBS 0.008948f
C800 B.n760 VSUBS 0.008948f
C801 B.n761 VSUBS 0.008948f
C802 B.n762 VSUBS 0.008948f
C803 B.n763 VSUBS 0.008948f
C804 B.n764 VSUBS 0.008948f
C805 B.n765 VSUBS 0.008948f
C806 B.n766 VSUBS 0.008948f
C807 B.n767 VSUBS 0.008948f
C808 B.n768 VSUBS 0.008948f
C809 B.n769 VSUBS 0.008948f
C810 B.n770 VSUBS 0.008948f
C811 B.n771 VSUBS 0.008948f
C812 B.n772 VSUBS 0.008948f
C813 B.n773 VSUBS 0.008948f
C814 B.n774 VSUBS 0.008948f
C815 B.n775 VSUBS 0.008948f
C816 B.n776 VSUBS 0.008948f
C817 B.n777 VSUBS 0.008948f
C818 B.n778 VSUBS 0.008948f
C819 B.n779 VSUBS 0.020262f
C820 VDD2.t5 VSUBS 4.85431f
C821 VDD2.t3 VSUBS 0.442355f
C822 VDD2.t8 VSUBS 0.442355f
C823 VDD2.n0 VSUBS 3.74086f
C824 VDD2.n1 VSUBS 1.36487f
C825 VDD2.t9 VSUBS 0.442355f
C826 VDD2.t7 VSUBS 0.442355f
C827 VDD2.n2 VSUBS 3.74674f
C828 VDD2.n3 VSUBS 3.00329f
C829 VDD2.t6 VSUBS 4.84542f
C830 VDD2.n4 VSUBS 3.70968f
C831 VDD2.t1 VSUBS 0.442355f
C832 VDD2.t4 VSUBS 0.442355f
C833 VDD2.n5 VSUBS 3.74086f
C834 VDD2.n6 VSUBS 0.646203f
C835 VDD2.t0 VSUBS 0.442355f
C836 VDD2.t2 VSUBS 0.442355f
C837 VDD2.n7 VSUBS 3.7467f
C838 VN.n0 VSUBS 0.048735f
C839 VN.n1 VSUBS 0.011059f
C840 VN.n2 VSUBS 0.203558f
C841 VN.t4 VSUBS 1.93825f
C842 VN.n3 VSUBS 0.698499f
C843 VN.t6 VSUBS 1.9169f
C844 VN.n4 VSUBS 0.72032f
C845 VN.n5 VSUBS 0.011059f
C846 VN.t1 VSUBS 1.9169f
C847 VN.n6 VSUBS 0.71541f
C848 VN.n7 VSUBS 0.048735f
C849 VN.n8 VSUBS 0.048735f
C850 VN.n9 VSUBS 0.048735f
C851 VN.t0 VSUBS 1.9169f
C852 VN.n10 VSUBS 0.71541f
C853 VN.n11 VSUBS 0.011059f
C854 VN.t2 VSUBS 1.9169f
C855 VN.n12 VSUBS 0.712706f
C856 VN.n13 VSUBS 0.037768f
C857 VN.n14 VSUBS 0.048735f
C858 VN.n15 VSUBS 0.011059f
C859 VN.t8 VSUBS 1.9169f
C860 VN.n16 VSUBS 0.203558f
C861 VN.t7 VSUBS 1.93825f
C862 VN.n17 VSUBS 0.698499f
C863 VN.t9 VSUBS 1.9169f
C864 VN.n18 VSUBS 0.72032f
C865 VN.n19 VSUBS 0.011059f
C866 VN.t5 VSUBS 1.9169f
C867 VN.n20 VSUBS 0.71541f
C868 VN.n21 VSUBS 0.048735f
C869 VN.n22 VSUBS 0.048735f
C870 VN.n23 VSUBS 0.048735f
C871 VN.n24 VSUBS 0.71541f
C872 VN.n25 VSUBS 0.011059f
C873 VN.t3 VSUBS 1.9169f
C874 VN.n26 VSUBS 0.712706f
C875 VN.n27 VSUBS 2.57959f
C876 VDD1.t9 VSUBS 4.85377f
C877 VDD1.t5 VSUBS 0.442305f
C878 VDD1.t1 VSUBS 0.442305f
C879 VDD1.n0 VSUBS 3.74044f
C880 VDD1.n1 VSUBS 1.37112f
C881 VDD1.t3 VSUBS 4.85377f
C882 VDD1.t4 VSUBS 0.442305f
C883 VDD1.t2 VSUBS 0.442305f
C884 VDD1.n2 VSUBS 3.74044f
C885 VDD1.n3 VSUBS 1.36472f
C886 VDD1.t7 VSUBS 0.442305f
C887 VDD1.t8 VSUBS 0.442305f
C888 VDD1.n4 VSUBS 3.74633f
C889 VDD1.n5 VSUBS 3.09197f
C890 VDD1.t6 VSUBS 0.442305f
C891 VDD1.t0 VSUBS 0.442305f
C892 VDD1.n6 VSUBS 3.74043f
C893 VDD1.n7 VSUBS 3.67786f
C894 VTAIL.t7 VSUBS 0.442509f
C895 VTAIL.t6 VSUBS 0.442509f
C896 VTAIL.n0 VSUBS 3.57742f
C897 VTAIL.n1 VSUBS 0.815539f
C898 VTAIL.t14 VSUBS 4.65675f
C899 VTAIL.n2 VSUBS 0.957951f
C900 VTAIL.t19 VSUBS 0.442509f
C901 VTAIL.t17 VSUBS 0.442509f
C902 VTAIL.n3 VSUBS 3.57742f
C903 VTAIL.n4 VSUBS 0.828083f
C904 VTAIL.t16 VSUBS 0.442509f
C905 VTAIL.t11 VSUBS 0.442509f
C906 VTAIL.n5 VSUBS 3.57742f
C907 VTAIL.n6 VSUBS 2.84772f
C908 VTAIL.t4 VSUBS 0.442509f
C909 VTAIL.t2 VSUBS 0.442509f
C910 VTAIL.n7 VSUBS 3.57742f
C911 VTAIL.n8 VSUBS 2.84772f
C912 VTAIL.t1 VSUBS 0.442509f
C913 VTAIL.t8 VSUBS 0.442509f
C914 VTAIL.n9 VSUBS 3.57742f
C915 VTAIL.n10 VSUBS 0.828082f
C916 VTAIL.t9 VSUBS 4.65675f
C917 VTAIL.n11 VSUBS 0.957949f
C918 VTAIL.t12 VSUBS 0.442509f
C919 VTAIL.t18 VSUBS 0.442509f
C920 VTAIL.n12 VSUBS 3.57742f
C921 VTAIL.n13 VSUBS 0.830434f
C922 VTAIL.t10 VSUBS 0.442509f
C923 VTAIL.t13 VSUBS 0.442509f
C924 VTAIL.n14 VSUBS 3.57742f
C925 VTAIL.n15 VSUBS 0.828082f
C926 VTAIL.t15 VSUBS 4.65675f
C927 VTAIL.n16 VSUBS 2.89448f
C928 VTAIL.t0 VSUBS 4.65675f
C929 VTAIL.n17 VSUBS 2.89448f
C930 VTAIL.t5 VSUBS 0.442509f
C931 VTAIL.t3 VSUBS 0.442509f
C932 VTAIL.n18 VSUBS 3.57742f
C933 VTAIL.n19 VSUBS 0.762226f
C934 VP.n0 VSUBS 0.049592f
C935 VP.n1 VSUBS 0.011254f
C936 VP.n2 VSUBS 0.049592f
C937 VP.n3 VSUBS 0.011254f
C938 VP.n4 VSUBS 0.049592f
C939 VP.t9 VSUBS 1.9506f
C940 VP.t3 VSUBS 1.9506f
C941 VP.n5 VSUBS 0.049592f
C942 VP.t8 VSUBS 1.9506f
C943 VP.n6 VSUBS 0.727989f
C944 VP.t0 VSUBS 1.97233f
C945 VP.n7 VSUBS 0.710781f
C946 VP.t4 VSUBS 1.9506f
C947 VP.n8 VSUBS 0.732986f
C948 VP.n9 VSUBS 0.011254f
C949 VP.n10 VSUBS 0.207138f
C950 VP.n11 VSUBS 0.049592f
C951 VP.n12 VSUBS 0.049592f
C952 VP.n13 VSUBS 0.011254f
C953 VP.n14 VSUBS 0.727989f
C954 VP.n15 VSUBS 0.011254f
C955 VP.n16 VSUBS 0.725237f
C956 VP.n17 VSUBS 2.59266f
C957 VP.t6 VSUBS 1.9506f
C958 VP.n18 VSUBS 0.725237f
C959 VP.n19 VSUBS 2.62935f
C960 VP.n20 VSUBS 0.049592f
C961 VP.n21 VSUBS 0.049592f
C962 VP.t5 VSUBS 1.9506f
C963 VP.n22 VSUBS 0.727989f
C964 VP.n23 VSUBS 0.011254f
C965 VP.t7 VSUBS 1.9506f
C966 VP.n24 VSUBS 0.727989f
C967 VP.n25 VSUBS 0.049592f
C968 VP.n26 VSUBS 0.049592f
C969 VP.n27 VSUBS 0.049592f
C970 VP.t2 VSUBS 1.9506f
C971 VP.n28 VSUBS 0.727989f
C972 VP.n29 VSUBS 0.011254f
C973 VP.t1 VSUBS 1.9506f
C974 VP.n30 VSUBS 0.725237f
C975 VP.n31 VSUBS 0.038432f
.ends

