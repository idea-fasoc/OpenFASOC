* NGSPICE file created from diff_pair_sample_0473.ext - technology: sky130A

.subckt diff_pair_sample_0473 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X1 VTAIL.t11 VP.t1 VDD1.t6 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=3.1944 ps=19.69 w=19.36 l=0.26
X2 VDD2.t7 VN.t0 VTAIL.t0 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X3 VDD1.t5 VP.t2 VTAIL.t13 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=7.5504 ps=39.5 w=19.36 l=0.26
X4 VTAIL.t7 VN.t1 VDD2.t6 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=3.1944 ps=19.69 w=19.36 l=0.26
X5 VTAIL.t1 VN.t2 VDD2.t5 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X6 VTAIL.t14 VP.t3 VDD1.t4 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X7 B.t11 B.t9 B.t10 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=0 ps=0 w=19.36 l=0.26
X8 VTAIL.t10 VP.t4 VDD1.t3 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=3.1944 ps=19.69 w=19.36 l=0.26
X9 VDD2.t4 VN.t3 VTAIL.t2 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=7.5504 ps=39.5 w=19.36 l=0.26
X10 VDD1.t2 VP.t5 VTAIL.t12 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X11 B.t8 B.t6 B.t7 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=0 ps=0 w=19.36 l=0.26
X12 VDD2.t3 VN.t4 VTAIL.t4 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X13 B.t5 B.t3 B.t4 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=0 ps=0 w=19.36 l=0.26
X14 VDD1.t1 VP.t6 VTAIL.t8 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=7.5504 ps=39.5 w=19.36 l=0.26
X15 VTAIL.t15 VP.t7 VDD1.t0 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X16 B.t2 B.t0 B.t1 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=0 ps=0 w=19.36 l=0.26
X17 VDD2.t2 VN.t5 VTAIL.t3 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=7.5504 ps=39.5 w=19.36 l=0.26
X18 VTAIL.t5 VN.t6 VDD2.t1 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=3.1944 pd=19.69 as=3.1944 ps=19.69 w=19.36 l=0.26
X19 VTAIL.t6 VN.t7 VDD2.t0 w_n1560_n4840# sky130_fd_pr__pfet_01v8 ad=7.5504 pd=39.5 as=3.1944 ps=19.69 w=19.36 l=0.26
R0 VP.n13 VP.t6 1971.26
R1 VP.n9 VP.t1 1971.26
R2 VP.n2 VP.t4 1971.26
R3 VP.n6 VP.t2 1971.26
R4 VP.n12 VP.t7 1915.02
R5 VP.n10 VP.t0 1915.02
R6 VP.n3 VP.t5 1915.02
R7 VP.n5 VP.t3 1915.02
R8 VP.n2 VP.n1 161.489
R9 VP.n14 VP.n13 161.3
R10 VP.n4 VP.n1 161.3
R11 VP.n7 VP.n6 161.3
R12 VP.n11 VP.n0 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n8 VP.n7 45.6596
R15 VP.n11 VP.n10 43.0884
R16 VP.n12 VP.n11 43.0884
R17 VP.n4 VP.n3 43.0884
R18 VP.n5 VP.n4 43.0884
R19 VP.n10 VP.n9 29.9429
R20 VP.n13 VP.n12 29.9429
R21 VP.n3 VP.n2 29.9429
R22 VP.n6 VP.n5 29.9429
R23 VP.n7 VP.n1 0.189894
R24 VP.n8 VP.n0 0.189894
R25 VP.n14 VP.n0 0.189894
R26 VP VP.n14 0.0516364
R27 VTAIL.n11 VTAIL.t10 54.0198
R28 VTAIL.n10 VTAIL.t2 54.0198
R29 VTAIL.n7 VTAIL.t6 54.0198
R30 VTAIL.n15 VTAIL.t3 54.0196
R31 VTAIL.n2 VTAIL.t7 54.0196
R32 VTAIL.n3 VTAIL.t8 54.0196
R33 VTAIL.n6 VTAIL.t11 54.0196
R34 VTAIL.n14 VTAIL.t13 54.0196
R35 VTAIL.n13 VTAIL.n12 52.3409
R36 VTAIL.n9 VTAIL.n8 52.3409
R37 VTAIL.n1 VTAIL.n0 52.3408
R38 VTAIL.n5 VTAIL.n4 52.3408
R39 VTAIL.n15 VTAIL.n14 29.5652
R40 VTAIL.n7 VTAIL.n6 29.5652
R41 VTAIL.n0 VTAIL.t4 1.67948
R42 VTAIL.n0 VTAIL.t5 1.67948
R43 VTAIL.n4 VTAIL.t9 1.67948
R44 VTAIL.n4 VTAIL.t15 1.67948
R45 VTAIL.n12 VTAIL.t12 1.67948
R46 VTAIL.n12 VTAIL.t14 1.67948
R47 VTAIL.n8 VTAIL.t0 1.67948
R48 VTAIL.n8 VTAIL.t1 1.67948
R49 VTAIL.n9 VTAIL.n7 0.509121
R50 VTAIL.n10 VTAIL.n9 0.509121
R51 VTAIL.n13 VTAIL.n11 0.509121
R52 VTAIL.n14 VTAIL.n13 0.509121
R53 VTAIL.n6 VTAIL.n5 0.509121
R54 VTAIL.n5 VTAIL.n3 0.509121
R55 VTAIL.n2 VTAIL.n1 0.509121
R56 VTAIL.n11 VTAIL.n10 0.470328
R57 VTAIL.n3 VTAIL.n2 0.470328
R58 VTAIL VTAIL.n15 0.450931
R59 VTAIL VTAIL.n1 0.0586897
R60 VDD1 VDD1.n0 69.3322
R61 VDD1.n3 VDD1.n2 69.2186
R62 VDD1.n3 VDD1.n1 69.2186
R63 VDD1.n5 VDD1.n4 69.0195
R64 VDD1.n5 VDD1.n3 43.2768
R65 VDD1.n4 VDD1.t4 1.67948
R66 VDD1.n4 VDD1.t5 1.67948
R67 VDD1.n0 VDD1.t3 1.67948
R68 VDD1.n0 VDD1.t2 1.67948
R69 VDD1.n2 VDD1.t0 1.67948
R70 VDD1.n2 VDD1.t1 1.67948
R71 VDD1.n1 VDD1.t6 1.67948
R72 VDD1.n1 VDD1.t7 1.67948
R73 VDD1 VDD1.n5 0.196621
R74 VN.n5 VN.t5 1971.26
R75 VN.n1 VN.t1 1971.26
R76 VN.n12 VN.t7 1971.26
R77 VN.n8 VN.t3 1971.26
R78 VN.n4 VN.t6 1915.02
R79 VN.n2 VN.t4 1915.02
R80 VN.n11 VN.t0 1915.02
R81 VN.n9 VN.t2 1915.02
R82 VN.n8 VN.n7 161.489
R83 VN.n1 VN.n0 161.489
R84 VN.n6 VN.n5 161.3
R85 VN.n13 VN.n12 161.3
R86 VN.n10 VN.n7 161.3
R87 VN.n3 VN.n0 161.3
R88 VN VN.n13 46.0403
R89 VN.n3 VN.n2 43.0884
R90 VN.n4 VN.n3 43.0884
R91 VN.n11 VN.n10 43.0884
R92 VN.n10 VN.n9 43.0884
R93 VN.n2 VN.n1 29.9429
R94 VN.n5 VN.n4 29.9429
R95 VN.n12 VN.n11 29.9429
R96 VN.n9 VN.n8 29.9429
R97 VN.n13 VN.n7 0.189894
R98 VN.n6 VN.n0 0.189894
R99 VN VN.n6 0.0516364
R100 VDD2.n2 VDD2.n1 69.2186
R101 VDD2.n2 VDD2.n0 69.2186
R102 VDD2 VDD2.n5 69.2156
R103 VDD2.n4 VDD2.n3 69.0197
R104 VDD2.n4 VDD2.n2 42.6937
R105 VDD2.n5 VDD2.t5 1.67948
R106 VDD2.n5 VDD2.t4 1.67948
R107 VDD2.n3 VDD2.t0 1.67948
R108 VDD2.n3 VDD2.t7 1.67948
R109 VDD2.n1 VDD2.t1 1.67948
R110 VDD2.n1 VDD2.t2 1.67948
R111 VDD2.n0 VDD2.t6 1.67948
R112 VDD2.n0 VDD2.t3 1.67948
R113 VDD2 VDD2.n4 0.313
R114 B.n132 B.t9 2016.97
R115 B.n140 B.t3 2016.97
R116 B.n42 B.t6 2016.97
R117 B.n50 B.t0 2016.97
R118 B.n464 B.n463 585
R119 B.n465 B.n82 585
R120 B.n467 B.n466 585
R121 B.n468 B.n81 585
R122 B.n470 B.n469 585
R123 B.n471 B.n80 585
R124 B.n473 B.n472 585
R125 B.n474 B.n79 585
R126 B.n476 B.n475 585
R127 B.n477 B.n78 585
R128 B.n479 B.n478 585
R129 B.n480 B.n77 585
R130 B.n482 B.n481 585
R131 B.n483 B.n76 585
R132 B.n485 B.n484 585
R133 B.n486 B.n75 585
R134 B.n488 B.n487 585
R135 B.n489 B.n74 585
R136 B.n491 B.n490 585
R137 B.n492 B.n73 585
R138 B.n494 B.n493 585
R139 B.n495 B.n72 585
R140 B.n497 B.n496 585
R141 B.n498 B.n71 585
R142 B.n500 B.n499 585
R143 B.n501 B.n70 585
R144 B.n503 B.n502 585
R145 B.n504 B.n69 585
R146 B.n506 B.n505 585
R147 B.n507 B.n68 585
R148 B.n509 B.n508 585
R149 B.n510 B.n67 585
R150 B.n512 B.n511 585
R151 B.n513 B.n66 585
R152 B.n515 B.n514 585
R153 B.n516 B.n65 585
R154 B.n518 B.n517 585
R155 B.n519 B.n64 585
R156 B.n521 B.n520 585
R157 B.n522 B.n63 585
R158 B.n524 B.n523 585
R159 B.n525 B.n62 585
R160 B.n527 B.n526 585
R161 B.n528 B.n61 585
R162 B.n530 B.n529 585
R163 B.n531 B.n60 585
R164 B.n533 B.n532 585
R165 B.n534 B.n59 585
R166 B.n536 B.n535 585
R167 B.n537 B.n58 585
R168 B.n539 B.n538 585
R169 B.n540 B.n57 585
R170 B.n542 B.n541 585
R171 B.n543 B.n56 585
R172 B.n545 B.n544 585
R173 B.n546 B.n55 585
R174 B.n548 B.n547 585
R175 B.n549 B.n54 585
R176 B.n551 B.n550 585
R177 B.n552 B.n53 585
R178 B.n554 B.n553 585
R179 B.n555 B.n52 585
R180 B.n557 B.n556 585
R181 B.n559 B.n49 585
R182 B.n561 B.n560 585
R183 B.n562 B.n48 585
R184 B.n564 B.n563 585
R185 B.n565 B.n47 585
R186 B.n567 B.n566 585
R187 B.n568 B.n46 585
R188 B.n570 B.n569 585
R189 B.n571 B.n45 585
R190 B.n573 B.n572 585
R191 B.n575 B.n574 585
R192 B.n576 B.n41 585
R193 B.n578 B.n577 585
R194 B.n579 B.n40 585
R195 B.n581 B.n580 585
R196 B.n582 B.n39 585
R197 B.n584 B.n583 585
R198 B.n585 B.n38 585
R199 B.n587 B.n586 585
R200 B.n588 B.n37 585
R201 B.n590 B.n589 585
R202 B.n591 B.n36 585
R203 B.n593 B.n592 585
R204 B.n594 B.n35 585
R205 B.n596 B.n595 585
R206 B.n597 B.n34 585
R207 B.n599 B.n598 585
R208 B.n600 B.n33 585
R209 B.n602 B.n601 585
R210 B.n603 B.n32 585
R211 B.n605 B.n604 585
R212 B.n606 B.n31 585
R213 B.n608 B.n607 585
R214 B.n609 B.n30 585
R215 B.n611 B.n610 585
R216 B.n612 B.n29 585
R217 B.n614 B.n613 585
R218 B.n615 B.n28 585
R219 B.n617 B.n616 585
R220 B.n618 B.n27 585
R221 B.n620 B.n619 585
R222 B.n621 B.n26 585
R223 B.n623 B.n622 585
R224 B.n624 B.n25 585
R225 B.n626 B.n625 585
R226 B.n627 B.n24 585
R227 B.n629 B.n628 585
R228 B.n630 B.n23 585
R229 B.n632 B.n631 585
R230 B.n633 B.n22 585
R231 B.n635 B.n634 585
R232 B.n636 B.n21 585
R233 B.n638 B.n637 585
R234 B.n639 B.n20 585
R235 B.n641 B.n640 585
R236 B.n642 B.n19 585
R237 B.n644 B.n643 585
R238 B.n645 B.n18 585
R239 B.n647 B.n646 585
R240 B.n648 B.n17 585
R241 B.n650 B.n649 585
R242 B.n651 B.n16 585
R243 B.n653 B.n652 585
R244 B.n654 B.n15 585
R245 B.n656 B.n655 585
R246 B.n657 B.n14 585
R247 B.n659 B.n658 585
R248 B.n660 B.n13 585
R249 B.n662 B.n661 585
R250 B.n663 B.n12 585
R251 B.n665 B.n664 585
R252 B.n666 B.n11 585
R253 B.n668 B.n667 585
R254 B.n462 B.n83 585
R255 B.n461 B.n460 585
R256 B.n459 B.n84 585
R257 B.n458 B.n457 585
R258 B.n456 B.n85 585
R259 B.n455 B.n454 585
R260 B.n453 B.n86 585
R261 B.n452 B.n451 585
R262 B.n450 B.n87 585
R263 B.n449 B.n448 585
R264 B.n447 B.n88 585
R265 B.n446 B.n445 585
R266 B.n444 B.n89 585
R267 B.n443 B.n442 585
R268 B.n441 B.n90 585
R269 B.n440 B.n439 585
R270 B.n438 B.n91 585
R271 B.n437 B.n436 585
R272 B.n435 B.n92 585
R273 B.n434 B.n433 585
R274 B.n432 B.n93 585
R275 B.n431 B.n430 585
R276 B.n429 B.n94 585
R277 B.n428 B.n427 585
R278 B.n426 B.n95 585
R279 B.n425 B.n424 585
R280 B.n423 B.n96 585
R281 B.n422 B.n421 585
R282 B.n420 B.n97 585
R283 B.n419 B.n418 585
R284 B.n417 B.n98 585
R285 B.n416 B.n415 585
R286 B.n414 B.n99 585
R287 B.n413 B.n412 585
R288 B.n411 B.n100 585
R289 B.n206 B.n205 585
R290 B.n207 B.n172 585
R291 B.n209 B.n208 585
R292 B.n210 B.n171 585
R293 B.n212 B.n211 585
R294 B.n213 B.n170 585
R295 B.n215 B.n214 585
R296 B.n216 B.n169 585
R297 B.n218 B.n217 585
R298 B.n219 B.n168 585
R299 B.n221 B.n220 585
R300 B.n222 B.n167 585
R301 B.n224 B.n223 585
R302 B.n225 B.n166 585
R303 B.n227 B.n226 585
R304 B.n228 B.n165 585
R305 B.n230 B.n229 585
R306 B.n231 B.n164 585
R307 B.n233 B.n232 585
R308 B.n234 B.n163 585
R309 B.n236 B.n235 585
R310 B.n237 B.n162 585
R311 B.n239 B.n238 585
R312 B.n240 B.n161 585
R313 B.n242 B.n241 585
R314 B.n243 B.n160 585
R315 B.n245 B.n244 585
R316 B.n246 B.n159 585
R317 B.n248 B.n247 585
R318 B.n249 B.n158 585
R319 B.n251 B.n250 585
R320 B.n252 B.n157 585
R321 B.n254 B.n253 585
R322 B.n255 B.n156 585
R323 B.n257 B.n256 585
R324 B.n258 B.n155 585
R325 B.n260 B.n259 585
R326 B.n261 B.n154 585
R327 B.n263 B.n262 585
R328 B.n264 B.n153 585
R329 B.n266 B.n265 585
R330 B.n267 B.n152 585
R331 B.n269 B.n268 585
R332 B.n270 B.n151 585
R333 B.n272 B.n271 585
R334 B.n273 B.n150 585
R335 B.n275 B.n274 585
R336 B.n276 B.n149 585
R337 B.n278 B.n277 585
R338 B.n279 B.n148 585
R339 B.n281 B.n280 585
R340 B.n282 B.n147 585
R341 B.n284 B.n283 585
R342 B.n285 B.n146 585
R343 B.n287 B.n286 585
R344 B.n288 B.n145 585
R345 B.n290 B.n289 585
R346 B.n291 B.n144 585
R347 B.n293 B.n292 585
R348 B.n294 B.n143 585
R349 B.n296 B.n295 585
R350 B.n297 B.n142 585
R351 B.n299 B.n298 585
R352 B.n301 B.n139 585
R353 B.n303 B.n302 585
R354 B.n304 B.n138 585
R355 B.n306 B.n305 585
R356 B.n307 B.n137 585
R357 B.n309 B.n308 585
R358 B.n310 B.n136 585
R359 B.n312 B.n311 585
R360 B.n313 B.n135 585
R361 B.n315 B.n314 585
R362 B.n317 B.n316 585
R363 B.n318 B.n131 585
R364 B.n320 B.n319 585
R365 B.n321 B.n130 585
R366 B.n323 B.n322 585
R367 B.n324 B.n129 585
R368 B.n326 B.n325 585
R369 B.n327 B.n128 585
R370 B.n329 B.n328 585
R371 B.n330 B.n127 585
R372 B.n332 B.n331 585
R373 B.n333 B.n126 585
R374 B.n335 B.n334 585
R375 B.n336 B.n125 585
R376 B.n338 B.n337 585
R377 B.n339 B.n124 585
R378 B.n341 B.n340 585
R379 B.n342 B.n123 585
R380 B.n344 B.n343 585
R381 B.n345 B.n122 585
R382 B.n347 B.n346 585
R383 B.n348 B.n121 585
R384 B.n350 B.n349 585
R385 B.n351 B.n120 585
R386 B.n353 B.n352 585
R387 B.n354 B.n119 585
R388 B.n356 B.n355 585
R389 B.n357 B.n118 585
R390 B.n359 B.n358 585
R391 B.n360 B.n117 585
R392 B.n362 B.n361 585
R393 B.n363 B.n116 585
R394 B.n365 B.n364 585
R395 B.n366 B.n115 585
R396 B.n368 B.n367 585
R397 B.n369 B.n114 585
R398 B.n371 B.n370 585
R399 B.n372 B.n113 585
R400 B.n374 B.n373 585
R401 B.n375 B.n112 585
R402 B.n377 B.n376 585
R403 B.n378 B.n111 585
R404 B.n380 B.n379 585
R405 B.n381 B.n110 585
R406 B.n383 B.n382 585
R407 B.n384 B.n109 585
R408 B.n386 B.n385 585
R409 B.n387 B.n108 585
R410 B.n389 B.n388 585
R411 B.n390 B.n107 585
R412 B.n392 B.n391 585
R413 B.n393 B.n106 585
R414 B.n395 B.n394 585
R415 B.n396 B.n105 585
R416 B.n398 B.n397 585
R417 B.n399 B.n104 585
R418 B.n401 B.n400 585
R419 B.n402 B.n103 585
R420 B.n404 B.n403 585
R421 B.n405 B.n102 585
R422 B.n407 B.n406 585
R423 B.n408 B.n101 585
R424 B.n410 B.n409 585
R425 B.n204 B.n173 585
R426 B.n203 B.n202 585
R427 B.n201 B.n174 585
R428 B.n200 B.n199 585
R429 B.n198 B.n175 585
R430 B.n197 B.n196 585
R431 B.n195 B.n176 585
R432 B.n194 B.n193 585
R433 B.n192 B.n177 585
R434 B.n191 B.n190 585
R435 B.n189 B.n178 585
R436 B.n188 B.n187 585
R437 B.n186 B.n179 585
R438 B.n185 B.n184 585
R439 B.n183 B.n180 585
R440 B.n182 B.n181 585
R441 B.n2 B.n0 585
R442 B.n693 B.n1 585
R443 B.n692 B.n691 585
R444 B.n690 B.n3 585
R445 B.n689 B.n688 585
R446 B.n687 B.n4 585
R447 B.n686 B.n685 585
R448 B.n684 B.n5 585
R449 B.n683 B.n682 585
R450 B.n681 B.n6 585
R451 B.n680 B.n679 585
R452 B.n678 B.n7 585
R453 B.n677 B.n676 585
R454 B.n675 B.n8 585
R455 B.n674 B.n673 585
R456 B.n672 B.n9 585
R457 B.n671 B.n670 585
R458 B.n669 B.n10 585
R459 B.n695 B.n694 585
R460 B.n206 B.n173 473.281
R461 B.n669 B.n668 473.281
R462 B.n411 B.n410 473.281
R463 B.n464 B.n83 473.281
R464 B.n202 B.n173 163.367
R465 B.n202 B.n201 163.367
R466 B.n201 B.n200 163.367
R467 B.n200 B.n175 163.367
R468 B.n196 B.n175 163.367
R469 B.n196 B.n195 163.367
R470 B.n195 B.n194 163.367
R471 B.n194 B.n177 163.367
R472 B.n190 B.n177 163.367
R473 B.n190 B.n189 163.367
R474 B.n189 B.n188 163.367
R475 B.n188 B.n179 163.367
R476 B.n184 B.n179 163.367
R477 B.n184 B.n183 163.367
R478 B.n183 B.n182 163.367
R479 B.n182 B.n2 163.367
R480 B.n694 B.n2 163.367
R481 B.n694 B.n693 163.367
R482 B.n693 B.n692 163.367
R483 B.n692 B.n3 163.367
R484 B.n688 B.n3 163.367
R485 B.n688 B.n687 163.367
R486 B.n687 B.n686 163.367
R487 B.n686 B.n5 163.367
R488 B.n682 B.n5 163.367
R489 B.n682 B.n681 163.367
R490 B.n681 B.n680 163.367
R491 B.n680 B.n7 163.367
R492 B.n676 B.n7 163.367
R493 B.n676 B.n675 163.367
R494 B.n675 B.n674 163.367
R495 B.n674 B.n9 163.367
R496 B.n670 B.n9 163.367
R497 B.n670 B.n669 163.367
R498 B.n207 B.n206 163.367
R499 B.n208 B.n207 163.367
R500 B.n208 B.n171 163.367
R501 B.n212 B.n171 163.367
R502 B.n213 B.n212 163.367
R503 B.n214 B.n213 163.367
R504 B.n214 B.n169 163.367
R505 B.n218 B.n169 163.367
R506 B.n219 B.n218 163.367
R507 B.n220 B.n219 163.367
R508 B.n220 B.n167 163.367
R509 B.n224 B.n167 163.367
R510 B.n225 B.n224 163.367
R511 B.n226 B.n225 163.367
R512 B.n226 B.n165 163.367
R513 B.n230 B.n165 163.367
R514 B.n231 B.n230 163.367
R515 B.n232 B.n231 163.367
R516 B.n232 B.n163 163.367
R517 B.n236 B.n163 163.367
R518 B.n237 B.n236 163.367
R519 B.n238 B.n237 163.367
R520 B.n238 B.n161 163.367
R521 B.n242 B.n161 163.367
R522 B.n243 B.n242 163.367
R523 B.n244 B.n243 163.367
R524 B.n244 B.n159 163.367
R525 B.n248 B.n159 163.367
R526 B.n249 B.n248 163.367
R527 B.n250 B.n249 163.367
R528 B.n250 B.n157 163.367
R529 B.n254 B.n157 163.367
R530 B.n255 B.n254 163.367
R531 B.n256 B.n255 163.367
R532 B.n256 B.n155 163.367
R533 B.n260 B.n155 163.367
R534 B.n261 B.n260 163.367
R535 B.n262 B.n261 163.367
R536 B.n262 B.n153 163.367
R537 B.n266 B.n153 163.367
R538 B.n267 B.n266 163.367
R539 B.n268 B.n267 163.367
R540 B.n268 B.n151 163.367
R541 B.n272 B.n151 163.367
R542 B.n273 B.n272 163.367
R543 B.n274 B.n273 163.367
R544 B.n274 B.n149 163.367
R545 B.n278 B.n149 163.367
R546 B.n279 B.n278 163.367
R547 B.n280 B.n279 163.367
R548 B.n280 B.n147 163.367
R549 B.n284 B.n147 163.367
R550 B.n285 B.n284 163.367
R551 B.n286 B.n285 163.367
R552 B.n286 B.n145 163.367
R553 B.n290 B.n145 163.367
R554 B.n291 B.n290 163.367
R555 B.n292 B.n291 163.367
R556 B.n292 B.n143 163.367
R557 B.n296 B.n143 163.367
R558 B.n297 B.n296 163.367
R559 B.n298 B.n297 163.367
R560 B.n298 B.n139 163.367
R561 B.n303 B.n139 163.367
R562 B.n304 B.n303 163.367
R563 B.n305 B.n304 163.367
R564 B.n305 B.n137 163.367
R565 B.n309 B.n137 163.367
R566 B.n310 B.n309 163.367
R567 B.n311 B.n310 163.367
R568 B.n311 B.n135 163.367
R569 B.n315 B.n135 163.367
R570 B.n316 B.n315 163.367
R571 B.n316 B.n131 163.367
R572 B.n320 B.n131 163.367
R573 B.n321 B.n320 163.367
R574 B.n322 B.n321 163.367
R575 B.n322 B.n129 163.367
R576 B.n326 B.n129 163.367
R577 B.n327 B.n326 163.367
R578 B.n328 B.n327 163.367
R579 B.n328 B.n127 163.367
R580 B.n332 B.n127 163.367
R581 B.n333 B.n332 163.367
R582 B.n334 B.n333 163.367
R583 B.n334 B.n125 163.367
R584 B.n338 B.n125 163.367
R585 B.n339 B.n338 163.367
R586 B.n340 B.n339 163.367
R587 B.n340 B.n123 163.367
R588 B.n344 B.n123 163.367
R589 B.n345 B.n344 163.367
R590 B.n346 B.n345 163.367
R591 B.n346 B.n121 163.367
R592 B.n350 B.n121 163.367
R593 B.n351 B.n350 163.367
R594 B.n352 B.n351 163.367
R595 B.n352 B.n119 163.367
R596 B.n356 B.n119 163.367
R597 B.n357 B.n356 163.367
R598 B.n358 B.n357 163.367
R599 B.n358 B.n117 163.367
R600 B.n362 B.n117 163.367
R601 B.n363 B.n362 163.367
R602 B.n364 B.n363 163.367
R603 B.n364 B.n115 163.367
R604 B.n368 B.n115 163.367
R605 B.n369 B.n368 163.367
R606 B.n370 B.n369 163.367
R607 B.n370 B.n113 163.367
R608 B.n374 B.n113 163.367
R609 B.n375 B.n374 163.367
R610 B.n376 B.n375 163.367
R611 B.n376 B.n111 163.367
R612 B.n380 B.n111 163.367
R613 B.n381 B.n380 163.367
R614 B.n382 B.n381 163.367
R615 B.n382 B.n109 163.367
R616 B.n386 B.n109 163.367
R617 B.n387 B.n386 163.367
R618 B.n388 B.n387 163.367
R619 B.n388 B.n107 163.367
R620 B.n392 B.n107 163.367
R621 B.n393 B.n392 163.367
R622 B.n394 B.n393 163.367
R623 B.n394 B.n105 163.367
R624 B.n398 B.n105 163.367
R625 B.n399 B.n398 163.367
R626 B.n400 B.n399 163.367
R627 B.n400 B.n103 163.367
R628 B.n404 B.n103 163.367
R629 B.n405 B.n404 163.367
R630 B.n406 B.n405 163.367
R631 B.n406 B.n101 163.367
R632 B.n410 B.n101 163.367
R633 B.n412 B.n411 163.367
R634 B.n412 B.n99 163.367
R635 B.n416 B.n99 163.367
R636 B.n417 B.n416 163.367
R637 B.n418 B.n417 163.367
R638 B.n418 B.n97 163.367
R639 B.n422 B.n97 163.367
R640 B.n423 B.n422 163.367
R641 B.n424 B.n423 163.367
R642 B.n424 B.n95 163.367
R643 B.n428 B.n95 163.367
R644 B.n429 B.n428 163.367
R645 B.n430 B.n429 163.367
R646 B.n430 B.n93 163.367
R647 B.n434 B.n93 163.367
R648 B.n435 B.n434 163.367
R649 B.n436 B.n435 163.367
R650 B.n436 B.n91 163.367
R651 B.n440 B.n91 163.367
R652 B.n441 B.n440 163.367
R653 B.n442 B.n441 163.367
R654 B.n442 B.n89 163.367
R655 B.n446 B.n89 163.367
R656 B.n447 B.n446 163.367
R657 B.n448 B.n447 163.367
R658 B.n448 B.n87 163.367
R659 B.n452 B.n87 163.367
R660 B.n453 B.n452 163.367
R661 B.n454 B.n453 163.367
R662 B.n454 B.n85 163.367
R663 B.n458 B.n85 163.367
R664 B.n459 B.n458 163.367
R665 B.n460 B.n459 163.367
R666 B.n460 B.n83 163.367
R667 B.n668 B.n11 163.367
R668 B.n664 B.n11 163.367
R669 B.n664 B.n663 163.367
R670 B.n663 B.n662 163.367
R671 B.n662 B.n13 163.367
R672 B.n658 B.n13 163.367
R673 B.n658 B.n657 163.367
R674 B.n657 B.n656 163.367
R675 B.n656 B.n15 163.367
R676 B.n652 B.n15 163.367
R677 B.n652 B.n651 163.367
R678 B.n651 B.n650 163.367
R679 B.n650 B.n17 163.367
R680 B.n646 B.n17 163.367
R681 B.n646 B.n645 163.367
R682 B.n645 B.n644 163.367
R683 B.n644 B.n19 163.367
R684 B.n640 B.n19 163.367
R685 B.n640 B.n639 163.367
R686 B.n639 B.n638 163.367
R687 B.n638 B.n21 163.367
R688 B.n634 B.n21 163.367
R689 B.n634 B.n633 163.367
R690 B.n633 B.n632 163.367
R691 B.n632 B.n23 163.367
R692 B.n628 B.n23 163.367
R693 B.n628 B.n627 163.367
R694 B.n627 B.n626 163.367
R695 B.n626 B.n25 163.367
R696 B.n622 B.n25 163.367
R697 B.n622 B.n621 163.367
R698 B.n621 B.n620 163.367
R699 B.n620 B.n27 163.367
R700 B.n616 B.n27 163.367
R701 B.n616 B.n615 163.367
R702 B.n615 B.n614 163.367
R703 B.n614 B.n29 163.367
R704 B.n610 B.n29 163.367
R705 B.n610 B.n609 163.367
R706 B.n609 B.n608 163.367
R707 B.n608 B.n31 163.367
R708 B.n604 B.n31 163.367
R709 B.n604 B.n603 163.367
R710 B.n603 B.n602 163.367
R711 B.n602 B.n33 163.367
R712 B.n598 B.n33 163.367
R713 B.n598 B.n597 163.367
R714 B.n597 B.n596 163.367
R715 B.n596 B.n35 163.367
R716 B.n592 B.n35 163.367
R717 B.n592 B.n591 163.367
R718 B.n591 B.n590 163.367
R719 B.n590 B.n37 163.367
R720 B.n586 B.n37 163.367
R721 B.n586 B.n585 163.367
R722 B.n585 B.n584 163.367
R723 B.n584 B.n39 163.367
R724 B.n580 B.n39 163.367
R725 B.n580 B.n579 163.367
R726 B.n579 B.n578 163.367
R727 B.n578 B.n41 163.367
R728 B.n574 B.n41 163.367
R729 B.n574 B.n573 163.367
R730 B.n573 B.n45 163.367
R731 B.n569 B.n45 163.367
R732 B.n569 B.n568 163.367
R733 B.n568 B.n567 163.367
R734 B.n567 B.n47 163.367
R735 B.n563 B.n47 163.367
R736 B.n563 B.n562 163.367
R737 B.n562 B.n561 163.367
R738 B.n561 B.n49 163.367
R739 B.n556 B.n49 163.367
R740 B.n556 B.n555 163.367
R741 B.n555 B.n554 163.367
R742 B.n554 B.n53 163.367
R743 B.n550 B.n53 163.367
R744 B.n550 B.n549 163.367
R745 B.n549 B.n548 163.367
R746 B.n548 B.n55 163.367
R747 B.n544 B.n55 163.367
R748 B.n544 B.n543 163.367
R749 B.n543 B.n542 163.367
R750 B.n542 B.n57 163.367
R751 B.n538 B.n57 163.367
R752 B.n538 B.n537 163.367
R753 B.n537 B.n536 163.367
R754 B.n536 B.n59 163.367
R755 B.n532 B.n59 163.367
R756 B.n532 B.n531 163.367
R757 B.n531 B.n530 163.367
R758 B.n530 B.n61 163.367
R759 B.n526 B.n61 163.367
R760 B.n526 B.n525 163.367
R761 B.n525 B.n524 163.367
R762 B.n524 B.n63 163.367
R763 B.n520 B.n63 163.367
R764 B.n520 B.n519 163.367
R765 B.n519 B.n518 163.367
R766 B.n518 B.n65 163.367
R767 B.n514 B.n65 163.367
R768 B.n514 B.n513 163.367
R769 B.n513 B.n512 163.367
R770 B.n512 B.n67 163.367
R771 B.n508 B.n67 163.367
R772 B.n508 B.n507 163.367
R773 B.n507 B.n506 163.367
R774 B.n506 B.n69 163.367
R775 B.n502 B.n69 163.367
R776 B.n502 B.n501 163.367
R777 B.n501 B.n500 163.367
R778 B.n500 B.n71 163.367
R779 B.n496 B.n71 163.367
R780 B.n496 B.n495 163.367
R781 B.n495 B.n494 163.367
R782 B.n494 B.n73 163.367
R783 B.n490 B.n73 163.367
R784 B.n490 B.n489 163.367
R785 B.n489 B.n488 163.367
R786 B.n488 B.n75 163.367
R787 B.n484 B.n75 163.367
R788 B.n484 B.n483 163.367
R789 B.n483 B.n482 163.367
R790 B.n482 B.n77 163.367
R791 B.n478 B.n77 163.367
R792 B.n478 B.n477 163.367
R793 B.n477 B.n476 163.367
R794 B.n476 B.n79 163.367
R795 B.n472 B.n79 163.367
R796 B.n472 B.n471 163.367
R797 B.n471 B.n470 163.367
R798 B.n470 B.n81 163.367
R799 B.n466 B.n81 163.367
R800 B.n466 B.n465 163.367
R801 B.n465 B.n464 163.367
R802 B.n132 B.t11 123.728
R803 B.n50 B.t1 123.728
R804 B.n140 B.t5 123.703
R805 B.n42 B.t7 123.703
R806 B.n133 B.t10 112.284
R807 B.n51 B.t2 112.284
R808 B.n141 B.t4 112.26
R809 B.n43 B.t8 112.26
R810 B.n134 B.n133 59.5399
R811 B.n300 B.n141 59.5399
R812 B.n44 B.n43 59.5399
R813 B.n558 B.n51 59.5399
R814 B.n667 B.n10 30.7517
R815 B.n463 B.n462 30.7517
R816 B.n409 B.n100 30.7517
R817 B.n205 B.n204 30.7517
R818 B B.n695 18.0485
R819 B.n133 B.n132 11.4429
R820 B.n141 B.n140 11.4429
R821 B.n43 B.n42 11.4429
R822 B.n51 B.n50 11.4429
R823 B.n667 B.n666 10.6151
R824 B.n666 B.n665 10.6151
R825 B.n665 B.n12 10.6151
R826 B.n661 B.n12 10.6151
R827 B.n661 B.n660 10.6151
R828 B.n660 B.n659 10.6151
R829 B.n659 B.n14 10.6151
R830 B.n655 B.n14 10.6151
R831 B.n655 B.n654 10.6151
R832 B.n654 B.n653 10.6151
R833 B.n653 B.n16 10.6151
R834 B.n649 B.n16 10.6151
R835 B.n649 B.n648 10.6151
R836 B.n648 B.n647 10.6151
R837 B.n647 B.n18 10.6151
R838 B.n643 B.n18 10.6151
R839 B.n643 B.n642 10.6151
R840 B.n642 B.n641 10.6151
R841 B.n641 B.n20 10.6151
R842 B.n637 B.n20 10.6151
R843 B.n637 B.n636 10.6151
R844 B.n636 B.n635 10.6151
R845 B.n635 B.n22 10.6151
R846 B.n631 B.n22 10.6151
R847 B.n631 B.n630 10.6151
R848 B.n630 B.n629 10.6151
R849 B.n629 B.n24 10.6151
R850 B.n625 B.n24 10.6151
R851 B.n625 B.n624 10.6151
R852 B.n624 B.n623 10.6151
R853 B.n623 B.n26 10.6151
R854 B.n619 B.n26 10.6151
R855 B.n619 B.n618 10.6151
R856 B.n618 B.n617 10.6151
R857 B.n617 B.n28 10.6151
R858 B.n613 B.n28 10.6151
R859 B.n613 B.n612 10.6151
R860 B.n612 B.n611 10.6151
R861 B.n611 B.n30 10.6151
R862 B.n607 B.n30 10.6151
R863 B.n607 B.n606 10.6151
R864 B.n606 B.n605 10.6151
R865 B.n605 B.n32 10.6151
R866 B.n601 B.n32 10.6151
R867 B.n601 B.n600 10.6151
R868 B.n600 B.n599 10.6151
R869 B.n599 B.n34 10.6151
R870 B.n595 B.n34 10.6151
R871 B.n595 B.n594 10.6151
R872 B.n594 B.n593 10.6151
R873 B.n593 B.n36 10.6151
R874 B.n589 B.n36 10.6151
R875 B.n589 B.n588 10.6151
R876 B.n588 B.n587 10.6151
R877 B.n587 B.n38 10.6151
R878 B.n583 B.n38 10.6151
R879 B.n583 B.n582 10.6151
R880 B.n582 B.n581 10.6151
R881 B.n581 B.n40 10.6151
R882 B.n577 B.n40 10.6151
R883 B.n577 B.n576 10.6151
R884 B.n576 B.n575 10.6151
R885 B.n572 B.n571 10.6151
R886 B.n571 B.n570 10.6151
R887 B.n570 B.n46 10.6151
R888 B.n566 B.n46 10.6151
R889 B.n566 B.n565 10.6151
R890 B.n565 B.n564 10.6151
R891 B.n564 B.n48 10.6151
R892 B.n560 B.n48 10.6151
R893 B.n560 B.n559 10.6151
R894 B.n557 B.n52 10.6151
R895 B.n553 B.n52 10.6151
R896 B.n553 B.n552 10.6151
R897 B.n552 B.n551 10.6151
R898 B.n551 B.n54 10.6151
R899 B.n547 B.n54 10.6151
R900 B.n547 B.n546 10.6151
R901 B.n546 B.n545 10.6151
R902 B.n545 B.n56 10.6151
R903 B.n541 B.n56 10.6151
R904 B.n541 B.n540 10.6151
R905 B.n540 B.n539 10.6151
R906 B.n539 B.n58 10.6151
R907 B.n535 B.n58 10.6151
R908 B.n535 B.n534 10.6151
R909 B.n534 B.n533 10.6151
R910 B.n533 B.n60 10.6151
R911 B.n529 B.n60 10.6151
R912 B.n529 B.n528 10.6151
R913 B.n528 B.n527 10.6151
R914 B.n527 B.n62 10.6151
R915 B.n523 B.n62 10.6151
R916 B.n523 B.n522 10.6151
R917 B.n522 B.n521 10.6151
R918 B.n521 B.n64 10.6151
R919 B.n517 B.n64 10.6151
R920 B.n517 B.n516 10.6151
R921 B.n516 B.n515 10.6151
R922 B.n515 B.n66 10.6151
R923 B.n511 B.n66 10.6151
R924 B.n511 B.n510 10.6151
R925 B.n510 B.n509 10.6151
R926 B.n509 B.n68 10.6151
R927 B.n505 B.n68 10.6151
R928 B.n505 B.n504 10.6151
R929 B.n504 B.n503 10.6151
R930 B.n503 B.n70 10.6151
R931 B.n499 B.n70 10.6151
R932 B.n499 B.n498 10.6151
R933 B.n498 B.n497 10.6151
R934 B.n497 B.n72 10.6151
R935 B.n493 B.n72 10.6151
R936 B.n493 B.n492 10.6151
R937 B.n492 B.n491 10.6151
R938 B.n491 B.n74 10.6151
R939 B.n487 B.n74 10.6151
R940 B.n487 B.n486 10.6151
R941 B.n486 B.n485 10.6151
R942 B.n485 B.n76 10.6151
R943 B.n481 B.n76 10.6151
R944 B.n481 B.n480 10.6151
R945 B.n480 B.n479 10.6151
R946 B.n479 B.n78 10.6151
R947 B.n475 B.n78 10.6151
R948 B.n475 B.n474 10.6151
R949 B.n474 B.n473 10.6151
R950 B.n473 B.n80 10.6151
R951 B.n469 B.n80 10.6151
R952 B.n469 B.n468 10.6151
R953 B.n468 B.n467 10.6151
R954 B.n467 B.n82 10.6151
R955 B.n463 B.n82 10.6151
R956 B.n413 B.n100 10.6151
R957 B.n414 B.n413 10.6151
R958 B.n415 B.n414 10.6151
R959 B.n415 B.n98 10.6151
R960 B.n419 B.n98 10.6151
R961 B.n420 B.n419 10.6151
R962 B.n421 B.n420 10.6151
R963 B.n421 B.n96 10.6151
R964 B.n425 B.n96 10.6151
R965 B.n426 B.n425 10.6151
R966 B.n427 B.n426 10.6151
R967 B.n427 B.n94 10.6151
R968 B.n431 B.n94 10.6151
R969 B.n432 B.n431 10.6151
R970 B.n433 B.n432 10.6151
R971 B.n433 B.n92 10.6151
R972 B.n437 B.n92 10.6151
R973 B.n438 B.n437 10.6151
R974 B.n439 B.n438 10.6151
R975 B.n439 B.n90 10.6151
R976 B.n443 B.n90 10.6151
R977 B.n444 B.n443 10.6151
R978 B.n445 B.n444 10.6151
R979 B.n445 B.n88 10.6151
R980 B.n449 B.n88 10.6151
R981 B.n450 B.n449 10.6151
R982 B.n451 B.n450 10.6151
R983 B.n451 B.n86 10.6151
R984 B.n455 B.n86 10.6151
R985 B.n456 B.n455 10.6151
R986 B.n457 B.n456 10.6151
R987 B.n457 B.n84 10.6151
R988 B.n461 B.n84 10.6151
R989 B.n462 B.n461 10.6151
R990 B.n205 B.n172 10.6151
R991 B.n209 B.n172 10.6151
R992 B.n210 B.n209 10.6151
R993 B.n211 B.n210 10.6151
R994 B.n211 B.n170 10.6151
R995 B.n215 B.n170 10.6151
R996 B.n216 B.n215 10.6151
R997 B.n217 B.n216 10.6151
R998 B.n217 B.n168 10.6151
R999 B.n221 B.n168 10.6151
R1000 B.n222 B.n221 10.6151
R1001 B.n223 B.n222 10.6151
R1002 B.n223 B.n166 10.6151
R1003 B.n227 B.n166 10.6151
R1004 B.n228 B.n227 10.6151
R1005 B.n229 B.n228 10.6151
R1006 B.n229 B.n164 10.6151
R1007 B.n233 B.n164 10.6151
R1008 B.n234 B.n233 10.6151
R1009 B.n235 B.n234 10.6151
R1010 B.n235 B.n162 10.6151
R1011 B.n239 B.n162 10.6151
R1012 B.n240 B.n239 10.6151
R1013 B.n241 B.n240 10.6151
R1014 B.n241 B.n160 10.6151
R1015 B.n245 B.n160 10.6151
R1016 B.n246 B.n245 10.6151
R1017 B.n247 B.n246 10.6151
R1018 B.n247 B.n158 10.6151
R1019 B.n251 B.n158 10.6151
R1020 B.n252 B.n251 10.6151
R1021 B.n253 B.n252 10.6151
R1022 B.n253 B.n156 10.6151
R1023 B.n257 B.n156 10.6151
R1024 B.n258 B.n257 10.6151
R1025 B.n259 B.n258 10.6151
R1026 B.n259 B.n154 10.6151
R1027 B.n263 B.n154 10.6151
R1028 B.n264 B.n263 10.6151
R1029 B.n265 B.n264 10.6151
R1030 B.n265 B.n152 10.6151
R1031 B.n269 B.n152 10.6151
R1032 B.n270 B.n269 10.6151
R1033 B.n271 B.n270 10.6151
R1034 B.n271 B.n150 10.6151
R1035 B.n275 B.n150 10.6151
R1036 B.n276 B.n275 10.6151
R1037 B.n277 B.n276 10.6151
R1038 B.n277 B.n148 10.6151
R1039 B.n281 B.n148 10.6151
R1040 B.n282 B.n281 10.6151
R1041 B.n283 B.n282 10.6151
R1042 B.n283 B.n146 10.6151
R1043 B.n287 B.n146 10.6151
R1044 B.n288 B.n287 10.6151
R1045 B.n289 B.n288 10.6151
R1046 B.n289 B.n144 10.6151
R1047 B.n293 B.n144 10.6151
R1048 B.n294 B.n293 10.6151
R1049 B.n295 B.n294 10.6151
R1050 B.n295 B.n142 10.6151
R1051 B.n299 B.n142 10.6151
R1052 B.n302 B.n301 10.6151
R1053 B.n302 B.n138 10.6151
R1054 B.n306 B.n138 10.6151
R1055 B.n307 B.n306 10.6151
R1056 B.n308 B.n307 10.6151
R1057 B.n308 B.n136 10.6151
R1058 B.n312 B.n136 10.6151
R1059 B.n313 B.n312 10.6151
R1060 B.n314 B.n313 10.6151
R1061 B.n318 B.n317 10.6151
R1062 B.n319 B.n318 10.6151
R1063 B.n319 B.n130 10.6151
R1064 B.n323 B.n130 10.6151
R1065 B.n324 B.n323 10.6151
R1066 B.n325 B.n324 10.6151
R1067 B.n325 B.n128 10.6151
R1068 B.n329 B.n128 10.6151
R1069 B.n330 B.n329 10.6151
R1070 B.n331 B.n330 10.6151
R1071 B.n331 B.n126 10.6151
R1072 B.n335 B.n126 10.6151
R1073 B.n336 B.n335 10.6151
R1074 B.n337 B.n336 10.6151
R1075 B.n337 B.n124 10.6151
R1076 B.n341 B.n124 10.6151
R1077 B.n342 B.n341 10.6151
R1078 B.n343 B.n342 10.6151
R1079 B.n343 B.n122 10.6151
R1080 B.n347 B.n122 10.6151
R1081 B.n348 B.n347 10.6151
R1082 B.n349 B.n348 10.6151
R1083 B.n349 B.n120 10.6151
R1084 B.n353 B.n120 10.6151
R1085 B.n354 B.n353 10.6151
R1086 B.n355 B.n354 10.6151
R1087 B.n355 B.n118 10.6151
R1088 B.n359 B.n118 10.6151
R1089 B.n360 B.n359 10.6151
R1090 B.n361 B.n360 10.6151
R1091 B.n361 B.n116 10.6151
R1092 B.n365 B.n116 10.6151
R1093 B.n366 B.n365 10.6151
R1094 B.n367 B.n366 10.6151
R1095 B.n367 B.n114 10.6151
R1096 B.n371 B.n114 10.6151
R1097 B.n372 B.n371 10.6151
R1098 B.n373 B.n372 10.6151
R1099 B.n373 B.n112 10.6151
R1100 B.n377 B.n112 10.6151
R1101 B.n378 B.n377 10.6151
R1102 B.n379 B.n378 10.6151
R1103 B.n379 B.n110 10.6151
R1104 B.n383 B.n110 10.6151
R1105 B.n384 B.n383 10.6151
R1106 B.n385 B.n384 10.6151
R1107 B.n385 B.n108 10.6151
R1108 B.n389 B.n108 10.6151
R1109 B.n390 B.n389 10.6151
R1110 B.n391 B.n390 10.6151
R1111 B.n391 B.n106 10.6151
R1112 B.n395 B.n106 10.6151
R1113 B.n396 B.n395 10.6151
R1114 B.n397 B.n396 10.6151
R1115 B.n397 B.n104 10.6151
R1116 B.n401 B.n104 10.6151
R1117 B.n402 B.n401 10.6151
R1118 B.n403 B.n402 10.6151
R1119 B.n403 B.n102 10.6151
R1120 B.n407 B.n102 10.6151
R1121 B.n408 B.n407 10.6151
R1122 B.n409 B.n408 10.6151
R1123 B.n204 B.n203 10.6151
R1124 B.n203 B.n174 10.6151
R1125 B.n199 B.n174 10.6151
R1126 B.n199 B.n198 10.6151
R1127 B.n198 B.n197 10.6151
R1128 B.n197 B.n176 10.6151
R1129 B.n193 B.n176 10.6151
R1130 B.n193 B.n192 10.6151
R1131 B.n192 B.n191 10.6151
R1132 B.n191 B.n178 10.6151
R1133 B.n187 B.n178 10.6151
R1134 B.n187 B.n186 10.6151
R1135 B.n186 B.n185 10.6151
R1136 B.n185 B.n180 10.6151
R1137 B.n181 B.n180 10.6151
R1138 B.n181 B.n0 10.6151
R1139 B.n691 B.n1 10.6151
R1140 B.n691 B.n690 10.6151
R1141 B.n690 B.n689 10.6151
R1142 B.n689 B.n4 10.6151
R1143 B.n685 B.n4 10.6151
R1144 B.n685 B.n684 10.6151
R1145 B.n684 B.n683 10.6151
R1146 B.n683 B.n6 10.6151
R1147 B.n679 B.n6 10.6151
R1148 B.n679 B.n678 10.6151
R1149 B.n678 B.n677 10.6151
R1150 B.n677 B.n8 10.6151
R1151 B.n673 B.n8 10.6151
R1152 B.n673 B.n672 10.6151
R1153 B.n672 B.n671 10.6151
R1154 B.n671 B.n10 10.6151
R1155 B.n575 B.n44 9.36635
R1156 B.n558 B.n557 9.36635
R1157 B.n300 B.n299 9.36635
R1158 B.n317 B.n134 9.36635
R1159 B.n695 B.n0 2.81026
R1160 B.n695 B.n1 2.81026
R1161 B.n572 B.n44 1.24928
R1162 B.n559 B.n558 1.24928
R1163 B.n301 B.n300 1.24928
R1164 B.n314 B.n134 1.24928
C0 w_n1560_n4840# VN 2.651f
C1 VN VP 6.15816f
C2 VN VDD1 0.147577f
C3 w_n1560_n4840# VP 2.84662f
C4 w_n1560_n4840# VDD1 1.31232f
C5 VP VDD1 4.8498f
C6 VN VTAIL 3.96982f
C7 B VN 0.764194f
C8 w_n1560_n4840# VTAIL 6.21134f
C9 B w_n1560_n4840# 8.632f
C10 VTAIL VP 3.98392f
C11 VTAIL VDD1 27.138f
C12 B VP 1.07965f
C13 B VDD1 1.13389f
C14 VDD2 VN 4.72684f
C15 VDD2 w_n1560_n4840# 1.32918f
C16 VDD2 VP 0.270749f
C17 VDD2 VDD1 0.6119f
C18 B VTAIL 5.27196f
C19 VDD2 VTAIL 27.1767f
C20 B VDD2 1.15724f
C21 VDD2 VSUBS 1.61473f
C22 VDD1 VSUBS 1.826384f
C23 VTAIL VSUBS 0.922057f
C24 VN VSUBS 5.31183f
C25 VP VSUBS 1.485857f
C26 B VSUBS 3.002973f
C27 w_n1560_n4840# VSUBS 92.2334f
C28 B.n0 VSUBS 0.005233f
C29 B.n1 VSUBS 0.005233f
C30 B.n2 VSUBS 0.008275f
C31 B.n3 VSUBS 0.008275f
C32 B.n4 VSUBS 0.008275f
C33 B.n5 VSUBS 0.008275f
C34 B.n6 VSUBS 0.008275f
C35 B.n7 VSUBS 0.008275f
C36 B.n8 VSUBS 0.008275f
C37 B.n9 VSUBS 0.008275f
C38 B.n10 VSUBS 0.018353f
C39 B.n11 VSUBS 0.008275f
C40 B.n12 VSUBS 0.008275f
C41 B.n13 VSUBS 0.008275f
C42 B.n14 VSUBS 0.008275f
C43 B.n15 VSUBS 0.008275f
C44 B.n16 VSUBS 0.008275f
C45 B.n17 VSUBS 0.008275f
C46 B.n18 VSUBS 0.008275f
C47 B.n19 VSUBS 0.008275f
C48 B.n20 VSUBS 0.008275f
C49 B.n21 VSUBS 0.008275f
C50 B.n22 VSUBS 0.008275f
C51 B.n23 VSUBS 0.008275f
C52 B.n24 VSUBS 0.008275f
C53 B.n25 VSUBS 0.008275f
C54 B.n26 VSUBS 0.008275f
C55 B.n27 VSUBS 0.008275f
C56 B.n28 VSUBS 0.008275f
C57 B.n29 VSUBS 0.008275f
C58 B.n30 VSUBS 0.008275f
C59 B.n31 VSUBS 0.008275f
C60 B.n32 VSUBS 0.008275f
C61 B.n33 VSUBS 0.008275f
C62 B.n34 VSUBS 0.008275f
C63 B.n35 VSUBS 0.008275f
C64 B.n36 VSUBS 0.008275f
C65 B.n37 VSUBS 0.008275f
C66 B.n38 VSUBS 0.008275f
C67 B.n39 VSUBS 0.008275f
C68 B.n40 VSUBS 0.008275f
C69 B.n41 VSUBS 0.008275f
C70 B.t8 VSUBS 0.776471f
C71 B.t7 VSUBS 0.782208f
C72 B.t6 VSUBS 0.229374f
C73 B.n42 VSUBS 0.137957f
C74 B.n43 VSUBS 0.073818f
C75 B.n44 VSUBS 0.019173f
C76 B.n45 VSUBS 0.008275f
C77 B.n46 VSUBS 0.008275f
C78 B.n47 VSUBS 0.008275f
C79 B.n48 VSUBS 0.008275f
C80 B.n49 VSUBS 0.008275f
C81 B.t2 VSUBS 0.77644f
C82 B.t1 VSUBS 0.782179f
C83 B.t0 VSUBS 0.229374f
C84 B.n50 VSUBS 0.137986f
C85 B.n51 VSUBS 0.073849f
C86 B.n52 VSUBS 0.008275f
C87 B.n53 VSUBS 0.008275f
C88 B.n54 VSUBS 0.008275f
C89 B.n55 VSUBS 0.008275f
C90 B.n56 VSUBS 0.008275f
C91 B.n57 VSUBS 0.008275f
C92 B.n58 VSUBS 0.008275f
C93 B.n59 VSUBS 0.008275f
C94 B.n60 VSUBS 0.008275f
C95 B.n61 VSUBS 0.008275f
C96 B.n62 VSUBS 0.008275f
C97 B.n63 VSUBS 0.008275f
C98 B.n64 VSUBS 0.008275f
C99 B.n65 VSUBS 0.008275f
C100 B.n66 VSUBS 0.008275f
C101 B.n67 VSUBS 0.008275f
C102 B.n68 VSUBS 0.008275f
C103 B.n69 VSUBS 0.008275f
C104 B.n70 VSUBS 0.008275f
C105 B.n71 VSUBS 0.008275f
C106 B.n72 VSUBS 0.008275f
C107 B.n73 VSUBS 0.008275f
C108 B.n74 VSUBS 0.008275f
C109 B.n75 VSUBS 0.008275f
C110 B.n76 VSUBS 0.008275f
C111 B.n77 VSUBS 0.008275f
C112 B.n78 VSUBS 0.008275f
C113 B.n79 VSUBS 0.008275f
C114 B.n80 VSUBS 0.008275f
C115 B.n81 VSUBS 0.008275f
C116 B.n82 VSUBS 0.008275f
C117 B.n83 VSUBS 0.018353f
C118 B.n84 VSUBS 0.008275f
C119 B.n85 VSUBS 0.008275f
C120 B.n86 VSUBS 0.008275f
C121 B.n87 VSUBS 0.008275f
C122 B.n88 VSUBS 0.008275f
C123 B.n89 VSUBS 0.008275f
C124 B.n90 VSUBS 0.008275f
C125 B.n91 VSUBS 0.008275f
C126 B.n92 VSUBS 0.008275f
C127 B.n93 VSUBS 0.008275f
C128 B.n94 VSUBS 0.008275f
C129 B.n95 VSUBS 0.008275f
C130 B.n96 VSUBS 0.008275f
C131 B.n97 VSUBS 0.008275f
C132 B.n98 VSUBS 0.008275f
C133 B.n99 VSUBS 0.008275f
C134 B.n100 VSUBS 0.018353f
C135 B.n101 VSUBS 0.008275f
C136 B.n102 VSUBS 0.008275f
C137 B.n103 VSUBS 0.008275f
C138 B.n104 VSUBS 0.008275f
C139 B.n105 VSUBS 0.008275f
C140 B.n106 VSUBS 0.008275f
C141 B.n107 VSUBS 0.008275f
C142 B.n108 VSUBS 0.008275f
C143 B.n109 VSUBS 0.008275f
C144 B.n110 VSUBS 0.008275f
C145 B.n111 VSUBS 0.008275f
C146 B.n112 VSUBS 0.008275f
C147 B.n113 VSUBS 0.008275f
C148 B.n114 VSUBS 0.008275f
C149 B.n115 VSUBS 0.008275f
C150 B.n116 VSUBS 0.008275f
C151 B.n117 VSUBS 0.008275f
C152 B.n118 VSUBS 0.008275f
C153 B.n119 VSUBS 0.008275f
C154 B.n120 VSUBS 0.008275f
C155 B.n121 VSUBS 0.008275f
C156 B.n122 VSUBS 0.008275f
C157 B.n123 VSUBS 0.008275f
C158 B.n124 VSUBS 0.008275f
C159 B.n125 VSUBS 0.008275f
C160 B.n126 VSUBS 0.008275f
C161 B.n127 VSUBS 0.008275f
C162 B.n128 VSUBS 0.008275f
C163 B.n129 VSUBS 0.008275f
C164 B.n130 VSUBS 0.008275f
C165 B.n131 VSUBS 0.008275f
C166 B.t10 VSUBS 0.77644f
C167 B.t11 VSUBS 0.782179f
C168 B.t9 VSUBS 0.229374f
C169 B.n132 VSUBS 0.137986f
C170 B.n133 VSUBS 0.073849f
C171 B.n134 VSUBS 0.019173f
C172 B.n135 VSUBS 0.008275f
C173 B.n136 VSUBS 0.008275f
C174 B.n137 VSUBS 0.008275f
C175 B.n138 VSUBS 0.008275f
C176 B.n139 VSUBS 0.008275f
C177 B.t4 VSUBS 0.776471f
C178 B.t5 VSUBS 0.782208f
C179 B.t3 VSUBS 0.229374f
C180 B.n140 VSUBS 0.137957f
C181 B.n141 VSUBS 0.073818f
C182 B.n142 VSUBS 0.008275f
C183 B.n143 VSUBS 0.008275f
C184 B.n144 VSUBS 0.008275f
C185 B.n145 VSUBS 0.008275f
C186 B.n146 VSUBS 0.008275f
C187 B.n147 VSUBS 0.008275f
C188 B.n148 VSUBS 0.008275f
C189 B.n149 VSUBS 0.008275f
C190 B.n150 VSUBS 0.008275f
C191 B.n151 VSUBS 0.008275f
C192 B.n152 VSUBS 0.008275f
C193 B.n153 VSUBS 0.008275f
C194 B.n154 VSUBS 0.008275f
C195 B.n155 VSUBS 0.008275f
C196 B.n156 VSUBS 0.008275f
C197 B.n157 VSUBS 0.008275f
C198 B.n158 VSUBS 0.008275f
C199 B.n159 VSUBS 0.008275f
C200 B.n160 VSUBS 0.008275f
C201 B.n161 VSUBS 0.008275f
C202 B.n162 VSUBS 0.008275f
C203 B.n163 VSUBS 0.008275f
C204 B.n164 VSUBS 0.008275f
C205 B.n165 VSUBS 0.008275f
C206 B.n166 VSUBS 0.008275f
C207 B.n167 VSUBS 0.008275f
C208 B.n168 VSUBS 0.008275f
C209 B.n169 VSUBS 0.008275f
C210 B.n170 VSUBS 0.008275f
C211 B.n171 VSUBS 0.008275f
C212 B.n172 VSUBS 0.008275f
C213 B.n173 VSUBS 0.018353f
C214 B.n174 VSUBS 0.008275f
C215 B.n175 VSUBS 0.008275f
C216 B.n176 VSUBS 0.008275f
C217 B.n177 VSUBS 0.008275f
C218 B.n178 VSUBS 0.008275f
C219 B.n179 VSUBS 0.008275f
C220 B.n180 VSUBS 0.008275f
C221 B.n181 VSUBS 0.008275f
C222 B.n182 VSUBS 0.008275f
C223 B.n183 VSUBS 0.008275f
C224 B.n184 VSUBS 0.008275f
C225 B.n185 VSUBS 0.008275f
C226 B.n186 VSUBS 0.008275f
C227 B.n187 VSUBS 0.008275f
C228 B.n188 VSUBS 0.008275f
C229 B.n189 VSUBS 0.008275f
C230 B.n190 VSUBS 0.008275f
C231 B.n191 VSUBS 0.008275f
C232 B.n192 VSUBS 0.008275f
C233 B.n193 VSUBS 0.008275f
C234 B.n194 VSUBS 0.008275f
C235 B.n195 VSUBS 0.008275f
C236 B.n196 VSUBS 0.008275f
C237 B.n197 VSUBS 0.008275f
C238 B.n198 VSUBS 0.008275f
C239 B.n199 VSUBS 0.008275f
C240 B.n200 VSUBS 0.008275f
C241 B.n201 VSUBS 0.008275f
C242 B.n202 VSUBS 0.008275f
C243 B.n203 VSUBS 0.008275f
C244 B.n204 VSUBS 0.018353f
C245 B.n205 VSUBS 0.018885f
C246 B.n206 VSUBS 0.018885f
C247 B.n207 VSUBS 0.008275f
C248 B.n208 VSUBS 0.008275f
C249 B.n209 VSUBS 0.008275f
C250 B.n210 VSUBS 0.008275f
C251 B.n211 VSUBS 0.008275f
C252 B.n212 VSUBS 0.008275f
C253 B.n213 VSUBS 0.008275f
C254 B.n214 VSUBS 0.008275f
C255 B.n215 VSUBS 0.008275f
C256 B.n216 VSUBS 0.008275f
C257 B.n217 VSUBS 0.008275f
C258 B.n218 VSUBS 0.008275f
C259 B.n219 VSUBS 0.008275f
C260 B.n220 VSUBS 0.008275f
C261 B.n221 VSUBS 0.008275f
C262 B.n222 VSUBS 0.008275f
C263 B.n223 VSUBS 0.008275f
C264 B.n224 VSUBS 0.008275f
C265 B.n225 VSUBS 0.008275f
C266 B.n226 VSUBS 0.008275f
C267 B.n227 VSUBS 0.008275f
C268 B.n228 VSUBS 0.008275f
C269 B.n229 VSUBS 0.008275f
C270 B.n230 VSUBS 0.008275f
C271 B.n231 VSUBS 0.008275f
C272 B.n232 VSUBS 0.008275f
C273 B.n233 VSUBS 0.008275f
C274 B.n234 VSUBS 0.008275f
C275 B.n235 VSUBS 0.008275f
C276 B.n236 VSUBS 0.008275f
C277 B.n237 VSUBS 0.008275f
C278 B.n238 VSUBS 0.008275f
C279 B.n239 VSUBS 0.008275f
C280 B.n240 VSUBS 0.008275f
C281 B.n241 VSUBS 0.008275f
C282 B.n242 VSUBS 0.008275f
C283 B.n243 VSUBS 0.008275f
C284 B.n244 VSUBS 0.008275f
C285 B.n245 VSUBS 0.008275f
C286 B.n246 VSUBS 0.008275f
C287 B.n247 VSUBS 0.008275f
C288 B.n248 VSUBS 0.008275f
C289 B.n249 VSUBS 0.008275f
C290 B.n250 VSUBS 0.008275f
C291 B.n251 VSUBS 0.008275f
C292 B.n252 VSUBS 0.008275f
C293 B.n253 VSUBS 0.008275f
C294 B.n254 VSUBS 0.008275f
C295 B.n255 VSUBS 0.008275f
C296 B.n256 VSUBS 0.008275f
C297 B.n257 VSUBS 0.008275f
C298 B.n258 VSUBS 0.008275f
C299 B.n259 VSUBS 0.008275f
C300 B.n260 VSUBS 0.008275f
C301 B.n261 VSUBS 0.008275f
C302 B.n262 VSUBS 0.008275f
C303 B.n263 VSUBS 0.008275f
C304 B.n264 VSUBS 0.008275f
C305 B.n265 VSUBS 0.008275f
C306 B.n266 VSUBS 0.008275f
C307 B.n267 VSUBS 0.008275f
C308 B.n268 VSUBS 0.008275f
C309 B.n269 VSUBS 0.008275f
C310 B.n270 VSUBS 0.008275f
C311 B.n271 VSUBS 0.008275f
C312 B.n272 VSUBS 0.008275f
C313 B.n273 VSUBS 0.008275f
C314 B.n274 VSUBS 0.008275f
C315 B.n275 VSUBS 0.008275f
C316 B.n276 VSUBS 0.008275f
C317 B.n277 VSUBS 0.008275f
C318 B.n278 VSUBS 0.008275f
C319 B.n279 VSUBS 0.008275f
C320 B.n280 VSUBS 0.008275f
C321 B.n281 VSUBS 0.008275f
C322 B.n282 VSUBS 0.008275f
C323 B.n283 VSUBS 0.008275f
C324 B.n284 VSUBS 0.008275f
C325 B.n285 VSUBS 0.008275f
C326 B.n286 VSUBS 0.008275f
C327 B.n287 VSUBS 0.008275f
C328 B.n288 VSUBS 0.008275f
C329 B.n289 VSUBS 0.008275f
C330 B.n290 VSUBS 0.008275f
C331 B.n291 VSUBS 0.008275f
C332 B.n292 VSUBS 0.008275f
C333 B.n293 VSUBS 0.008275f
C334 B.n294 VSUBS 0.008275f
C335 B.n295 VSUBS 0.008275f
C336 B.n296 VSUBS 0.008275f
C337 B.n297 VSUBS 0.008275f
C338 B.n298 VSUBS 0.008275f
C339 B.n299 VSUBS 0.007788f
C340 B.n300 VSUBS 0.019173f
C341 B.n301 VSUBS 0.004624f
C342 B.n302 VSUBS 0.008275f
C343 B.n303 VSUBS 0.008275f
C344 B.n304 VSUBS 0.008275f
C345 B.n305 VSUBS 0.008275f
C346 B.n306 VSUBS 0.008275f
C347 B.n307 VSUBS 0.008275f
C348 B.n308 VSUBS 0.008275f
C349 B.n309 VSUBS 0.008275f
C350 B.n310 VSUBS 0.008275f
C351 B.n311 VSUBS 0.008275f
C352 B.n312 VSUBS 0.008275f
C353 B.n313 VSUBS 0.008275f
C354 B.n314 VSUBS 0.004624f
C355 B.n315 VSUBS 0.008275f
C356 B.n316 VSUBS 0.008275f
C357 B.n317 VSUBS 0.007788f
C358 B.n318 VSUBS 0.008275f
C359 B.n319 VSUBS 0.008275f
C360 B.n320 VSUBS 0.008275f
C361 B.n321 VSUBS 0.008275f
C362 B.n322 VSUBS 0.008275f
C363 B.n323 VSUBS 0.008275f
C364 B.n324 VSUBS 0.008275f
C365 B.n325 VSUBS 0.008275f
C366 B.n326 VSUBS 0.008275f
C367 B.n327 VSUBS 0.008275f
C368 B.n328 VSUBS 0.008275f
C369 B.n329 VSUBS 0.008275f
C370 B.n330 VSUBS 0.008275f
C371 B.n331 VSUBS 0.008275f
C372 B.n332 VSUBS 0.008275f
C373 B.n333 VSUBS 0.008275f
C374 B.n334 VSUBS 0.008275f
C375 B.n335 VSUBS 0.008275f
C376 B.n336 VSUBS 0.008275f
C377 B.n337 VSUBS 0.008275f
C378 B.n338 VSUBS 0.008275f
C379 B.n339 VSUBS 0.008275f
C380 B.n340 VSUBS 0.008275f
C381 B.n341 VSUBS 0.008275f
C382 B.n342 VSUBS 0.008275f
C383 B.n343 VSUBS 0.008275f
C384 B.n344 VSUBS 0.008275f
C385 B.n345 VSUBS 0.008275f
C386 B.n346 VSUBS 0.008275f
C387 B.n347 VSUBS 0.008275f
C388 B.n348 VSUBS 0.008275f
C389 B.n349 VSUBS 0.008275f
C390 B.n350 VSUBS 0.008275f
C391 B.n351 VSUBS 0.008275f
C392 B.n352 VSUBS 0.008275f
C393 B.n353 VSUBS 0.008275f
C394 B.n354 VSUBS 0.008275f
C395 B.n355 VSUBS 0.008275f
C396 B.n356 VSUBS 0.008275f
C397 B.n357 VSUBS 0.008275f
C398 B.n358 VSUBS 0.008275f
C399 B.n359 VSUBS 0.008275f
C400 B.n360 VSUBS 0.008275f
C401 B.n361 VSUBS 0.008275f
C402 B.n362 VSUBS 0.008275f
C403 B.n363 VSUBS 0.008275f
C404 B.n364 VSUBS 0.008275f
C405 B.n365 VSUBS 0.008275f
C406 B.n366 VSUBS 0.008275f
C407 B.n367 VSUBS 0.008275f
C408 B.n368 VSUBS 0.008275f
C409 B.n369 VSUBS 0.008275f
C410 B.n370 VSUBS 0.008275f
C411 B.n371 VSUBS 0.008275f
C412 B.n372 VSUBS 0.008275f
C413 B.n373 VSUBS 0.008275f
C414 B.n374 VSUBS 0.008275f
C415 B.n375 VSUBS 0.008275f
C416 B.n376 VSUBS 0.008275f
C417 B.n377 VSUBS 0.008275f
C418 B.n378 VSUBS 0.008275f
C419 B.n379 VSUBS 0.008275f
C420 B.n380 VSUBS 0.008275f
C421 B.n381 VSUBS 0.008275f
C422 B.n382 VSUBS 0.008275f
C423 B.n383 VSUBS 0.008275f
C424 B.n384 VSUBS 0.008275f
C425 B.n385 VSUBS 0.008275f
C426 B.n386 VSUBS 0.008275f
C427 B.n387 VSUBS 0.008275f
C428 B.n388 VSUBS 0.008275f
C429 B.n389 VSUBS 0.008275f
C430 B.n390 VSUBS 0.008275f
C431 B.n391 VSUBS 0.008275f
C432 B.n392 VSUBS 0.008275f
C433 B.n393 VSUBS 0.008275f
C434 B.n394 VSUBS 0.008275f
C435 B.n395 VSUBS 0.008275f
C436 B.n396 VSUBS 0.008275f
C437 B.n397 VSUBS 0.008275f
C438 B.n398 VSUBS 0.008275f
C439 B.n399 VSUBS 0.008275f
C440 B.n400 VSUBS 0.008275f
C441 B.n401 VSUBS 0.008275f
C442 B.n402 VSUBS 0.008275f
C443 B.n403 VSUBS 0.008275f
C444 B.n404 VSUBS 0.008275f
C445 B.n405 VSUBS 0.008275f
C446 B.n406 VSUBS 0.008275f
C447 B.n407 VSUBS 0.008275f
C448 B.n408 VSUBS 0.008275f
C449 B.n409 VSUBS 0.018885f
C450 B.n410 VSUBS 0.018885f
C451 B.n411 VSUBS 0.018353f
C452 B.n412 VSUBS 0.008275f
C453 B.n413 VSUBS 0.008275f
C454 B.n414 VSUBS 0.008275f
C455 B.n415 VSUBS 0.008275f
C456 B.n416 VSUBS 0.008275f
C457 B.n417 VSUBS 0.008275f
C458 B.n418 VSUBS 0.008275f
C459 B.n419 VSUBS 0.008275f
C460 B.n420 VSUBS 0.008275f
C461 B.n421 VSUBS 0.008275f
C462 B.n422 VSUBS 0.008275f
C463 B.n423 VSUBS 0.008275f
C464 B.n424 VSUBS 0.008275f
C465 B.n425 VSUBS 0.008275f
C466 B.n426 VSUBS 0.008275f
C467 B.n427 VSUBS 0.008275f
C468 B.n428 VSUBS 0.008275f
C469 B.n429 VSUBS 0.008275f
C470 B.n430 VSUBS 0.008275f
C471 B.n431 VSUBS 0.008275f
C472 B.n432 VSUBS 0.008275f
C473 B.n433 VSUBS 0.008275f
C474 B.n434 VSUBS 0.008275f
C475 B.n435 VSUBS 0.008275f
C476 B.n436 VSUBS 0.008275f
C477 B.n437 VSUBS 0.008275f
C478 B.n438 VSUBS 0.008275f
C479 B.n439 VSUBS 0.008275f
C480 B.n440 VSUBS 0.008275f
C481 B.n441 VSUBS 0.008275f
C482 B.n442 VSUBS 0.008275f
C483 B.n443 VSUBS 0.008275f
C484 B.n444 VSUBS 0.008275f
C485 B.n445 VSUBS 0.008275f
C486 B.n446 VSUBS 0.008275f
C487 B.n447 VSUBS 0.008275f
C488 B.n448 VSUBS 0.008275f
C489 B.n449 VSUBS 0.008275f
C490 B.n450 VSUBS 0.008275f
C491 B.n451 VSUBS 0.008275f
C492 B.n452 VSUBS 0.008275f
C493 B.n453 VSUBS 0.008275f
C494 B.n454 VSUBS 0.008275f
C495 B.n455 VSUBS 0.008275f
C496 B.n456 VSUBS 0.008275f
C497 B.n457 VSUBS 0.008275f
C498 B.n458 VSUBS 0.008275f
C499 B.n459 VSUBS 0.008275f
C500 B.n460 VSUBS 0.008275f
C501 B.n461 VSUBS 0.008275f
C502 B.n462 VSUBS 0.019392f
C503 B.n463 VSUBS 0.017847f
C504 B.n464 VSUBS 0.018885f
C505 B.n465 VSUBS 0.008275f
C506 B.n466 VSUBS 0.008275f
C507 B.n467 VSUBS 0.008275f
C508 B.n468 VSUBS 0.008275f
C509 B.n469 VSUBS 0.008275f
C510 B.n470 VSUBS 0.008275f
C511 B.n471 VSUBS 0.008275f
C512 B.n472 VSUBS 0.008275f
C513 B.n473 VSUBS 0.008275f
C514 B.n474 VSUBS 0.008275f
C515 B.n475 VSUBS 0.008275f
C516 B.n476 VSUBS 0.008275f
C517 B.n477 VSUBS 0.008275f
C518 B.n478 VSUBS 0.008275f
C519 B.n479 VSUBS 0.008275f
C520 B.n480 VSUBS 0.008275f
C521 B.n481 VSUBS 0.008275f
C522 B.n482 VSUBS 0.008275f
C523 B.n483 VSUBS 0.008275f
C524 B.n484 VSUBS 0.008275f
C525 B.n485 VSUBS 0.008275f
C526 B.n486 VSUBS 0.008275f
C527 B.n487 VSUBS 0.008275f
C528 B.n488 VSUBS 0.008275f
C529 B.n489 VSUBS 0.008275f
C530 B.n490 VSUBS 0.008275f
C531 B.n491 VSUBS 0.008275f
C532 B.n492 VSUBS 0.008275f
C533 B.n493 VSUBS 0.008275f
C534 B.n494 VSUBS 0.008275f
C535 B.n495 VSUBS 0.008275f
C536 B.n496 VSUBS 0.008275f
C537 B.n497 VSUBS 0.008275f
C538 B.n498 VSUBS 0.008275f
C539 B.n499 VSUBS 0.008275f
C540 B.n500 VSUBS 0.008275f
C541 B.n501 VSUBS 0.008275f
C542 B.n502 VSUBS 0.008275f
C543 B.n503 VSUBS 0.008275f
C544 B.n504 VSUBS 0.008275f
C545 B.n505 VSUBS 0.008275f
C546 B.n506 VSUBS 0.008275f
C547 B.n507 VSUBS 0.008275f
C548 B.n508 VSUBS 0.008275f
C549 B.n509 VSUBS 0.008275f
C550 B.n510 VSUBS 0.008275f
C551 B.n511 VSUBS 0.008275f
C552 B.n512 VSUBS 0.008275f
C553 B.n513 VSUBS 0.008275f
C554 B.n514 VSUBS 0.008275f
C555 B.n515 VSUBS 0.008275f
C556 B.n516 VSUBS 0.008275f
C557 B.n517 VSUBS 0.008275f
C558 B.n518 VSUBS 0.008275f
C559 B.n519 VSUBS 0.008275f
C560 B.n520 VSUBS 0.008275f
C561 B.n521 VSUBS 0.008275f
C562 B.n522 VSUBS 0.008275f
C563 B.n523 VSUBS 0.008275f
C564 B.n524 VSUBS 0.008275f
C565 B.n525 VSUBS 0.008275f
C566 B.n526 VSUBS 0.008275f
C567 B.n527 VSUBS 0.008275f
C568 B.n528 VSUBS 0.008275f
C569 B.n529 VSUBS 0.008275f
C570 B.n530 VSUBS 0.008275f
C571 B.n531 VSUBS 0.008275f
C572 B.n532 VSUBS 0.008275f
C573 B.n533 VSUBS 0.008275f
C574 B.n534 VSUBS 0.008275f
C575 B.n535 VSUBS 0.008275f
C576 B.n536 VSUBS 0.008275f
C577 B.n537 VSUBS 0.008275f
C578 B.n538 VSUBS 0.008275f
C579 B.n539 VSUBS 0.008275f
C580 B.n540 VSUBS 0.008275f
C581 B.n541 VSUBS 0.008275f
C582 B.n542 VSUBS 0.008275f
C583 B.n543 VSUBS 0.008275f
C584 B.n544 VSUBS 0.008275f
C585 B.n545 VSUBS 0.008275f
C586 B.n546 VSUBS 0.008275f
C587 B.n547 VSUBS 0.008275f
C588 B.n548 VSUBS 0.008275f
C589 B.n549 VSUBS 0.008275f
C590 B.n550 VSUBS 0.008275f
C591 B.n551 VSUBS 0.008275f
C592 B.n552 VSUBS 0.008275f
C593 B.n553 VSUBS 0.008275f
C594 B.n554 VSUBS 0.008275f
C595 B.n555 VSUBS 0.008275f
C596 B.n556 VSUBS 0.008275f
C597 B.n557 VSUBS 0.007788f
C598 B.n558 VSUBS 0.019173f
C599 B.n559 VSUBS 0.004624f
C600 B.n560 VSUBS 0.008275f
C601 B.n561 VSUBS 0.008275f
C602 B.n562 VSUBS 0.008275f
C603 B.n563 VSUBS 0.008275f
C604 B.n564 VSUBS 0.008275f
C605 B.n565 VSUBS 0.008275f
C606 B.n566 VSUBS 0.008275f
C607 B.n567 VSUBS 0.008275f
C608 B.n568 VSUBS 0.008275f
C609 B.n569 VSUBS 0.008275f
C610 B.n570 VSUBS 0.008275f
C611 B.n571 VSUBS 0.008275f
C612 B.n572 VSUBS 0.004624f
C613 B.n573 VSUBS 0.008275f
C614 B.n574 VSUBS 0.008275f
C615 B.n575 VSUBS 0.007788f
C616 B.n576 VSUBS 0.008275f
C617 B.n577 VSUBS 0.008275f
C618 B.n578 VSUBS 0.008275f
C619 B.n579 VSUBS 0.008275f
C620 B.n580 VSUBS 0.008275f
C621 B.n581 VSUBS 0.008275f
C622 B.n582 VSUBS 0.008275f
C623 B.n583 VSUBS 0.008275f
C624 B.n584 VSUBS 0.008275f
C625 B.n585 VSUBS 0.008275f
C626 B.n586 VSUBS 0.008275f
C627 B.n587 VSUBS 0.008275f
C628 B.n588 VSUBS 0.008275f
C629 B.n589 VSUBS 0.008275f
C630 B.n590 VSUBS 0.008275f
C631 B.n591 VSUBS 0.008275f
C632 B.n592 VSUBS 0.008275f
C633 B.n593 VSUBS 0.008275f
C634 B.n594 VSUBS 0.008275f
C635 B.n595 VSUBS 0.008275f
C636 B.n596 VSUBS 0.008275f
C637 B.n597 VSUBS 0.008275f
C638 B.n598 VSUBS 0.008275f
C639 B.n599 VSUBS 0.008275f
C640 B.n600 VSUBS 0.008275f
C641 B.n601 VSUBS 0.008275f
C642 B.n602 VSUBS 0.008275f
C643 B.n603 VSUBS 0.008275f
C644 B.n604 VSUBS 0.008275f
C645 B.n605 VSUBS 0.008275f
C646 B.n606 VSUBS 0.008275f
C647 B.n607 VSUBS 0.008275f
C648 B.n608 VSUBS 0.008275f
C649 B.n609 VSUBS 0.008275f
C650 B.n610 VSUBS 0.008275f
C651 B.n611 VSUBS 0.008275f
C652 B.n612 VSUBS 0.008275f
C653 B.n613 VSUBS 0.008275f
C654 B.n614 VSUBS 0.008275f
C655 B.n615 VSUBS 0.008275f
C656 B.n616 VSUBS 0.008275f
C657 B.n617 VSUBS 0.008275f
C658 B.n618 VSUBS 0.008275f
C659 B.n619 VSUBS 0.008275f
C660 B.n620 VSUBS 0.008275f
C661 B.n621 VSUBS 0.008275f
C662 B.n622 VSUBS 0.008275f
C663 B.n623 VSUBS 0.008275f
C664 B.n624 VSUBS 0.008275f
C665 B.n625 VSUBS 0.008275f
C666 B.n626 VSUBS 0.008275f
C667 B.n627 VSUBS 0.008275f
C668 B.n628 VSUBS 0.008275f
C669 B.n629 VSUBS 0.008275f
C670 B.n630 VSUBS 0.008275f
C671 B.n631 VSUBS 0.008275f
C672 B.n632 VSUBS 0.008275f
C673 B.n633 VSUBS 0.008275f
C674 B.n634 VSUBS 0.008275f
C675 B.n635 VSUBS 0.008275f
C676 B.n636 VSUBS 0.008275f
C677 B.n637 VSUBS 0.008275f
C678 B.n638 VSUBS 0.008275f
C679 B.n639 VSUBS 0.008275f
C680 B.n640 VSUBS 0.008275f
C681 B.n641 VSUBS 0.008275f
C682 B.n642 VSUBS 0.008275f
C683 B.n643 VSUBS 0.008275f
C684 B.n644 VSUBS 0.008275f
C685 B.n645 VSUBS 0.008275f
C686 B.n646 VSUBS 0.008275f
C687 B.n647 VSUBS 0.008275f
C688 B.n648 VSUBS 0.008275f
C689 B.n649 VSUBS 0.008275f
C690 B.n650 VSUBS 0.008275f
C691 B.n651 VSUBS 0.008275f
C692 B.n652 VSUBS 0.008275f
C693 B.n653 VSUBS 0.008275f
C694 B.n654 VSUBS 0.008275f
C695 B.n655 VSUBS 0.008275f
C696 B.n656 VSUBS 0.008275f
C697 B.n657 VSUBS 0.008275f
C698 B.n658 VSUBS 0.008275f
C699 B.n659 VSUBS 0.008275f
C700 B.n660 VSUBS 0.008275f
C701 B.n661 VSUBS 0.008275f
C702 B.n662 VSUBS 0.008275f
C703 B.n663 VSUBS 0.008275f
C704 B.n664 VSUBS 0.008275f
C705 B.n665 VSUBS 0.008275f
C706 B.n666 VSUBS 0.008275f
C707 B.n667 VSUBS 0.018885f
C708 B.n668 VSUBS 0.018885f
C709 B.n669 VSUBS 0.018353f
C710 B.n670 VSUBS 0.008275f
C711 B.n671 VSUBS 0.008275f
C712 B.n672 VSUBS 0.008275f
C713 B.n673 VSUBS 0.008275f
C714 B.n674 VSUBS 0.008275f
C715 B.n675 VSUBS 0.008275f
C716 B.n676 VSUBS 0.008275f
C717 B.n677 VSUBS 0.008275f
C718 B.n678 VSUBS 0.008275f
C719 B.n679 VSUBS 0.008275f
C720 B.n680 VSUBS 0.008275f
C721 B.n681 VSUBS 0.008275f
C722 B.n682 VSUBS 0.008275f
C723 B.n683 VSUBS 0.008275f
C724 B.n684 VSUBS 0.008275f
C725 B.n685 VSUBS 0.008275f
C726 B.n686 VSUBS 0.008275f
C727 B.n687 VSUBS 0.008275f
C728 B.n688 VSUBS 0.008275f
C729 B.n689 VSUBS 0.008275f
C730 B.n690 VSUBS 0.008275f
C731 B.n691 VSUBS 0.008275f
C732 B.n692 VSUBS 0.008275f
C733 B.n693 VSUBS 0.008275f
C734 B.n694 VSUBS 0.008275f
C735 B.n695 VSUBS 0.018738f
C736 VDD2.t6 VSUBS 0.543764f
C737 VDD2.t3 VSUBS 0.543764f
C738 VDD2.n0 VSUBS 4.56231f
C739 VDD2.t1 VSUBS 0.543764f
C740 VDD2.t2 VSUBS 0.543764f
C741 VDD2.n1 VSUBS 4.56231f
C742 VDD2.n2 VSUBS 4.19302f
C743 VDD2.t0 VSUBS 0.543764f
C744 VDD2.t7 VSUBS 0.543764f
C745 VDD2.n3 VSUBS 4.56f
C746 VDD2.n4 VSUBS 4.25454f
C747 VDD2.t5 VSUBS 0.543764f
C748 VDD2.t4 VSUBS 0.543764f
C749 VDD2.n5 VSUBS 4.56224f
C750 VN.n0 VSUBS 0.157334f
C751 VN.t6 VSUBS 0.959437f
C752 VN.t4 VSUBS 0.959437f
C753 VN.t1 VSUBS 0.969891f
C754 VN.n1 VSUBS 0.382295f
C755 VN.n2 VSUBS 0.360393f
C756 VN.n3 VSUBS 0.026201f
C757 VN.n4 VSUBS 0.360393f
C758 VN.t5 VSUBS 0.969891f
C759 VN.n5 VSUBS 0.382189f
C760 VN.n6 VSUBS 0.052437f
C761 VN.n7 VSUBS 0.157334f
C762 VN.t7 VSUBS 0.969891f
C763 VN.t0 VSUBS 0.959437f
C764 VN.t2 VSUBS 0.959437f
C765 VN.t3 VSUBS 0.969891f
C766 VN.n8 VSUBS 0.382295f
C767 VN.n9 VSUBS 0.360393f
C768 VN.n10 VSUBS 0.026201f
C769 VN.n11 VSUBS 0.360393f
C770 VN.n12 VSUBS 0.382189f
C771 VN.n13 VSUBS 3.24247f
C772 VDD1.t3 VSUBS 0.541535f
C773 VDD1.t2 VSUBS 0.541535f
C774 VDD1.n0 VSUBS 4.54496f
C775 VDD1.t6 VSUBS 0.541535f
C776 VDD1.t7 VSUBS 0.541535f
C777 VDD1.n1 VSUBS 4.54361f
C778 VDD1.t0 VSUBS 0.541535f
C779 VDD1.t1 VSUBS 0.541535f
C780 VDD1.n2 VSUBS 4.54361f
C781 VDD1.n3 VSUBS 4.2512f
C782 VDD1.t4 VSUBS 0.541535f
C783 VDD1.t5 VSUBS 0.541535f
C784 VDD1.n4 VSUBS 4.54129f
C785 VDD1.n5 VSUBS 4.27922f
C786 VTAIL.t4 VSUBS 0.447055f
C787 VTAIL.t5 VSUBS 0.447055f
C788 VTAIL.n0 VSUBS 3.56622f
C789 VTAIL.n1 VSUBS 0.775586f
C790 VTAIL.t7 VSUBS 4.65061f
C791 VTAIL.n2 VSUBS 0.949196f
C792 VTAIL.t8 VSUBS 4.65061f
C793 VTAIL.n3 VSUBS 0.949196f
C794 VTAIL.t9 VSUBS 0.447055f
C795 VTAIL.t15 VSUBS 0.447055f
C796 VTAIL.n4 VSUBS 3.56622f
C797 VTAIL.n5 VSUBS 0.817998f
C798 VTAIL.t11 VSUBS 4.65061f
C799 VTAIL.n6 VSUBS 2.92125f
C800 VTAIL.t6 VSUBS 4.65062f
C801 VTAIL.n7 VSUBS 2.92125f
C802 VTAIL.t0 VSUBS 0.447055f
C803 VTAIL.t1 VSUBS 0.447055f
C804 VTAIL.n8 VSUBS 3.56622f
C805 VTAIL.n9 VSUBS 0.817998f
C806 VTAIL.t2 VSUBS 4.65062f
C807 VTAIL.n10 VSUBS 0.949187f
C808 VTAIL.t10 VSUBS 4.65062f
C809 VTAIL.n11 VSUBS 0.949187f
C810 VTAIL.t12 VSUBS 0.447055f
C811 VTAIL.t14 VSUBS 0.447055f
C812 VTAIL.n12 VSUBS 3.56622f
C813 VTAIL.n13 VSUBS 0.817998f
C814 VTAIL.t13 VSUBS 4.65061f
C815 VTAIL.n14 VSUBS 2.92125f
C816 VTAIL.t3 VSUBS 4.65061f
C817 VTAIL.n15 VSUBS 2.91578f
C818 VP.n0 VSUBS 0.068805f
C819 VP.t7 VSUBS 0.975613f
C820 VP.t0 VSUBS 0.975613f
C821 VP.t1 VSUBS 0.986242f
C822 VP.n1 VSUBS 0.159986f
C823 VP.t3 VSUBS 0.975613f
C824 VP.t5 VSUBS 0.975613f
C825 VP.t4 VSUBS 0.986242f
C826 VP.n2 VSUBS 0.38874f
C827 VP.n3 VSUBS 0.366469f
C828 VP.n4 VSUBS 0.026643f
C829 VP.n5 VSUBS 0.366469f
C830 VP.t2 VSUBS 0.986242f
C831 VP.n6 VSUBS 0.388633f
C832 VP.n7 VSUBS 3.25219f
C833 VP.n8 VSUBS 3.30651f
C834 VP.n9 VSUBS 0.388633f
C835 VP.n10 VSUBS 0.366469f
C836 VP.n11 VSUBS 0.026643f
C837 VP.n12 VSUBS 0.366469f
C838 VP.t6 VSUBS 0.986242f
C839 VP.n13 VSUBS 0.388633f
C840 VP.n14 VSUBS 0.053321f
.ends

