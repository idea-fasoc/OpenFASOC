* NGSPICE file created from diff_pair_sample_1776.ext - technology: sky130A

.subckt diff_pair_sample_1776 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=5.4951 ps=28.96 w=14.09 l=2.52
X1 VDD1.t6 VP.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=5.4951 ps=28.96 w=14.09 l=2.52
X2 VTAIL.t11 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=2.32485 ps=14.42 w=14.09 l=2.52
X3 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=0 ps=0 w=14.09 l=2.52
X4 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=0 ps=0 w=14.09 l=2.52
X5 VTAIL.t13 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X6 VTAIL.t9 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X7 VTAIL.t7 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=2.32485 ps=14.42 w=14.09 l=2.52
X8 VDD2.t6 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X9 VTAIL.t3 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X10 VDD1.t2 VP.t5 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X11 VDD2.t4 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=5.4951 ps=28.96 w=14.09 l=2.52
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=0 ps=0 w=14.09 l=2.52
X13 VTAIL.t10 VP.t6 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=2.32485 ps=14.42 w=14.09 l=2.52
X14 VTAIL.t1 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X15 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=2.32485 ps=14.42 w=14.09 l=2.52
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4951 pd=28.96 as=0 ps=0 w=14.09 l=2.52
X17 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=5.4951 ps=28.96 w=14.09 l=2.52
X18 VDD2.t0 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
X19 VDD1.t0 VP.t7 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.32485 pd=14.42 as=2.32485 ps=14.42 w=14.09 l=2.52
R0 VP.n16 VP.t6 169.323
R1 VP.n19 VP.n18 161.3
R2 VP.n20 VP.n15 161.3
R3 VP.n22 VP.n21 161.3
R4 VP.n23 VP.n14 161.3
R5 VP.n25 VP.n24 161.3
R6 VP.n27 VP.n26 161.3
R7 VP.n28 VP.n12 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n31 VP.n11 161.3
R10 VP.n33 VP.n32 161.3
R11 VP.n34 VP.n10 161.3
R12 VP.n64 VP.n0 161.3
R13 VP.n63 VP.n62 161.3
R14 VP.n61 VP.n1 161.3
R15 VP.n60 VP.n59 161.3
R16 VP.n58 VP.n2 161.3
R17 VP.n57 VP.n56 161.3
R18 VP.n55 VP.n54 161.3
R19 VP.n53 VP.n4 161.3
R20 VP.n52 VP.n51 161.3
R21 VP.n50 VP.n5 161.3
R22 VP.n49 VP.n48 161.3
R23 VP.n46 VP.n6 161.3
R24 VP.n45 VP.n44 161.3
R25 VP.n43 VP.n7 161.3
R26 VP.n42 VP.n41 161.3
R27 VP.n40 VP.n8 161.3
R28 VP.n39 VP.n38 161.3
R29 VP.n9 VP.t2 134.75
R30 VP.n47 VP.t7 134.75
R31 VP.n3 VP.t3 134.75
R32 VP.n65 VP.t1 134.75
R33 VP.n35 VP.t0 134.75
R34 VP.n13 VP.t4 134.75
R35 VP.n17 VP.t5 134.75
R36 VP.n37 VP.n9 97.2996
R37 VP.n66 VP.n65 97.2996
R38 VP.n36 VP.n35 97.2996
R39 VP.n41 VP.n7 55.0624
R40 VP.n59 VP.n1 55.0624
R41 VP.n29 VP.n11 55.0624
R42 VP.n37 VP.n36 52.1587
R43 VP.n17 VP.n16 51.8291
R44 VP.n52 VP.n5 40.4934
R45 VP.n53 VP.n52 40.4934
R46 VP.n23 VP.n22 40.4934
R47 VP.n22 VP.n15 40.4934
R48 VP.n41 VP.n40 25.9244
R49 VP.n63 VP.n1 25.9244
R50 VP.n33 VP.n11 25.9244
R51 VP.n40 VP.n39 24.4675
R52 VP.n45 VP.n7 24.4675
R53 VP.n46 VP.n45 24.4675
R54 VP.n48 VP.n5 24.4675
R55 VP.n54 VP.n53 24.4675
R56 VP.n58 VP.n57 24.4675
R57 VP.n59 VP.n58 24.4675
R58 VP.n64 VP.n63 24.4675
R59 VP.n34 VP.n33 24.4675
R60 VP.n24 VP.n23 24.4675
R61 VP.n28 VP.n27 24.4675
R62 VP.n29 VP.n28 24.4675
R63 VP.n18 VP.n15 24.4675
R64 VP.n48 VP.n47 20.7975
R65 VP.n54 VP.n3 20.7975
R66 VP.n24 VP.n13 20.7975
R67 VP.n18 VP.n17 20.7975
R68 VP.n39 VP.n9 13.4574
R69 VP.n65 VP.n64 13.4574
R70 VP.n35 VP.n34 13.4574
R71 VP.n19 VP.n16 6.62497
R72 VP.n47 VP.n46 3.67055
R73 VP.n57 VP.n3 3.67055
R74 VP.n27 VP.n13 3.67055
R75 VP.n36 VP.n10 0.278367
R76 VP.n38 VP.n37 0.278367
R77 VP.n66 VP.n0 0.278367
R78 VP.n20 VP.n19 0.189894
R79 VP.n21 VP.n20 0.189894
R80 VP.n21 VP.n14 0.189894
R81 VP.n25 VP.n14 0.189894
R82 VP.n26 VP.n25 0.189894
R83 VP.n26 VP.n12 0.189894
R84 VP.n30 VP.n12 0.189894
R85 VP.n31 VP.n30 0.189894
R86 VP.n32 VP.n31 0.189894
R87 VP.n32 VP.n10 0.189894
R88 VP.n38 VP.n8 0.189894
R89 VP.n42 VP.n8 0.189894
R90 VP.n43 VP.n42 0.189894
R91 VP.n44 VP.n43 0.189894
R92 VP.n44 VP.n6 0.189894
R93 VP.n49 VP.n6 0.189894
R94 VP.n50 VP.n49 0.189894
R95 VP.n51 VP.n50 0.189894
R96 VP.n51 VP.n4 0.189894
R97 VP.n55 VP.n4 0.189894
R98 VP.n56 VP.n55 0.189894
R99 VP.n56 VP.n2 0.189894
R100 VP.n60 VP.n2 0.189894
R101 VP.n61 VP.n60 0.189894
R102 VP.n62 VP.n61 0.189894
R103 VP.n62 VP.n0 0.189894
R104 VP VP.n66 0.153454
R105 VTAIL.n626 VTAIL.n554 289.615
R106 VTAIL.n74 VTAIL.n2 289.615
R107 VTAIL.n152 VTAIL.n80 289.615
R108 VTAIL.n232 VTAIL.n160 289.615
R109 VTAIL.n548 VTAIL.n476 289.615
R110 VTAIL.n468 VTAIL.n396 289.615
R111 VTAIL.n390 VTAIL.n318 289.615
R112 VTAIL.n310 VTAIL.n238 289.615
R113 VTAIL.n578 VTAIL.n577 185
R114 VTAIL.n583 VTAIL.n582 185
R115 VTAIL.n585 VTAIL.n584 185
R116 VTAIL.n574 VTAIL.n573 185
R117 VTAIL.n591 VTAIL.n590 185
R118 VTAIL.n593 VTAIL.n592 185
R119 VTAIL.n570 VTAIL.n569 185
R120 VTAIL.n599 VTAIL.n598 185
R121 VTAIL.n601 VTAIL.n600 185
R122 VTAIL.n566 VTAIL.n565 185
R123 VTAIL.n607 VTAIL.n606 185
R124 VTAIL.n609 VTAIL.n608 185
R125 VTAIL.n562 VTAIL.n561 185
R126 VTAIL.n615 VTAIL.n614 185
R127 VTAIL.n617 VTAIL.n616 185
R128 VTAIL.n558 VTAIL.n557 185
R129 VTAIL.n624 VTAIL.n623 185
R130 VTAIL.n625 VTAIL.n556 185
R131 VTAIL.n627 VTAIL.n626 185
R132 VTAIL.n26 VTAIL.n25 185
R133 VTAIL.n31 VTAIL.n30 185
R134 VTAIL.n33 VTAIL.n32 185
R135 VTAIL.n22 VTAIL.n21 185
R136 VTAIL.n39 VTAIL.n38 185
R137 VTAIL.n41 VTAIL.n40 185
R138 VTAIL.n18 VTAIL.n17 185
R139 VTAIL.n47 VTAIL.n46 185
R140 VTAIL.n49 VTAIL.n48 185
R141 VTAIL.n14 VTAIL.n13 185
R142 VTAIL.n55 VTAIL.n54 185
R143 VTAIL.n57 VTAIL.n56 185
R144 VTAIL.n10 VTAIL.n9 185
R145 VTAIL.n63 VTAIL.n62 185
R146 VTAIL.n65 VTAIL.n64 185
R147 VTAIL.n6 VTAIL.n5 185
R148 VTAIL.n72 VTAIL.n71 185
R149 VTAIL.n73 VTAIL.n4 185
R150 VTAIL.n75 VTAIL.n74 185
R151 VTAIL.n104 VTAIL.n103 185
R152 VTAIL.n109 VTAIL.n108 185
R153 VTAIL.n111 VTAIL.n110 185
R154 VTAIL.n100 VTAIL.n99 185
R155 VTAIL.n117 VTAIL.n116 185
R156 VTAIL.n119 VTAIL.n118 185
R157 VTAIL.n96 VTAIL.n95 185
R158 VTAIL.n125 VTAIL.n124 185
R159 VTAIL.n127 VTAIL.n126 185
R160 VTAIL.n92 VTAIL.n91 185
R161 VTAIL.n133 VTAIL.n132 185
R162 VTAIL.n135 VTAIL.n134 185
R163 VTAIL.n88 VTAIL.n87 185
R164 VTAIL.n141 VTAIL.n140 185
R165 VTAIL.n143 VTAIL.n142 185
R166 VTAIL.n84 VTAIL.n83 185
R167 VTAIL.n150 VTAIL.n149 185
R168 VTAIL.n151 VTAIL.n82 185
R169 VTAIL.n153 VTAIL.n152 185
R170 VTAIL.n184 VTAIL.n183 185
R171 VTAIL.n189 VTAIL.n188 185
R172 VTAIL.n191 VTAIL.n190 185
R173 VTAIL.n180 VTAIL.n179 185
R174 VTAIL.n197 VTAIL.n196 185
R175 VTAIL.n199 VTAIL.n198 185
R176 VTAIL.n176 VTAIL.n175 185
R177 VTAIL.n205 VTAIL.n204 185
R178 VTAIL.n207 VTAIL.n206 185
R179 VTAIL.n172 VTAIL.n171 185
R180 VTAIL.n213 VTAIL.n212 185
R181 VTAIL.n215 VTAIL.n214 185
R182 VTAIL.n168 VTAIL.n167 185
R183 VTAIL.n221 VTAIL.n220 185
R184 VTAIL.n223 VTAIL.n222 185
R185 VTAIL.n164 VTAIL.n163 185
R186 VTAIL.n230 VTAIL.n229 185
R187 VTAIL.n231 VTAIL.n162 185
R188 VTAIL.n233 VTAIL.n232 185
R189 VTAIL.n549 VTAIL.n548 185
R190 VTAIL.n547 VTAIL.n478 185
R191 VTAIL.n546 VTAIL.n545 185
R192 VTAIL.n481 VTAIL.n479 185
R193 VTAIL.n540 VTAIL.n539 185
R194 VTAIL.n538 VTAIL.n537 185
R195 VTAIL.n485 VTAIL.n484 185
R196 VTAIL.n532 VTAIL.n531 185
R197 VTAIL.n530 VTAIL.n529 185
R198 VTAIL.n489 VTAIL.n488 185
R199 VTAIL.n524 VTAIL.n523 185
R200 VTAIL.n522 VTAIL.n521 185
R201 VTAIL.n493 VTAIL.n492 185
R202 VTAIL.n516 VTAIL.n515 185
R203 VTAIL.n514 VTAIL.n513 185
R204 VTAIL.n497 VTAIL.n496 185
R205 VTAIL.n508 VTAIL.n507 185
R206 VTAIL.n506 VTAIL.n505 185
R207 VTAIL.n501 VTAIL.n500 185
R208 VTAIL.n469 VTAIL.n468 185
R209 VTAIL.n467 VTAIL.n398 185
R210 VTAIL.n466 VTAIL.n465 185
R211 VTAIL.n401 VTAIL.n399 185
R212 VTAIL.n460 VTAIL.n459 185
R213 VTAIL.n458 VTAIL.n457 185
R214 VTAIL.n405 VTAIL.n404 185
R215 VTAIL.n452 VTAIL.n451 185
R216 VTAIL.n450 VTAIL.n449 185
R217 VTAIL.n409 VTAIL.n408 185
R218 VTAIL.n444 VTAIL.n443 185
R219 VTAIL.n442 VTAIL.n441 185
R220 VTAIL.n413 VTAIL.n412 185
R221 VTAIL.n436 VTAIL.n435 185
R222 VTAIL.n434 VTAIL.n433 185
R223 VTAIL.n417 VTAIL.n416 185
R224 VTAIL.n428 VTAIL.n427 185
R225 VTAIL.n426 VTAIL.n425 185
R226 VTAIL.n421 VTAIL.n420 185
R227 VTAIL.n391 VTAIL.n390 185
R228 VTAIL.n389 VTAIL.n320 185
R229 VTAIL.n388 VTAIL.n387 185
R230 VTAIL.n323 VTAIL.n321 185
R231 VTAIL.n382 VTAIL.n381 185
R232 VTAIL.n380 VTAIL.n379 185
R233 VTAIL.n327 VTAIL.n326 185
R234 VTAIL.n374 VTAIL.n373 185
R235 VTAIL.n372 VTAIL.n371 185
R236 VTAIL.n331 VTAIL.n330 185
R237 VTAIL.n366 VTAIL.n365 185
R238 VTAIL.n364 VTAIL.n363 185
R239 VTAIL.n335 VTAIL.n334 185
R240 VTAIL.n358 VTAIL.n357 185
R241 VTAIL.n356 VTAIL.n355 185
R242 VTAIL.n339 VTAIL.n338 185
R243 VTAIL.n350 VTAIL.n349 185
R244 VTAIL.n348 VTAIL.n347 185
R245 VTAIL.n343 VTAIL.n342 185
R246 VTAIL.n311 VTAIL.n310 185
R247 VTAIL.n309 VTAIL.n240 185
R248 VTAIL.n308 VTAIL.n307 185
R249 VTAIL.n243 VTAIL.n241 185
R250 VTAIL.n302 VTAIL.n301 185
R251 VTAIL.n300 VTAIL.n299 185
R252 VTAIL.n247 VTAIL.n246 185
R253 VTAIL.n294 VTAIL.n293 185
R254 VTAIL.n292 VTAIL.n291 185
R255 VTAIL.n251 VTAIL.n250 185
R256 VTAIL.n286 VTAIL.n285 185
R257 VTAIL.n284 VTAIL.n283 185
R258 VTAIL.n255 VTAIL.n254 185
R259 VTAIL.n278 VTAIL.n277 185
R260 VTAIL.n276 VTAIL.n275 185
R261 VTAIL.n259 VTAIL.n258 185
R262 VTAIL.n270 VTAIL.n269 185
R263 VTAIL.n268 VTAIL.n267 185
R264 VTAIL.n263 VTAIL.n262 185
R265 VTAIL.n579 VTAIL.t2 147.659
R266 VTAIL.n27 VTAIL.t0 147.659
R267 VTAIL.n105 VTAIL.t8 147.659
R268 VTAIL.n185 VTAIL.t11 147.659
R269 VTAIL.n502 VTAIL.t12 147.659
R270 VTAIL.n422 VTAIL.t10 147.659
R271 VTAIL.n344 VTAIL.t4 147.659
R272 VTAIL.n264 VTAIL.t7 147.659
R273 VTAIL.n583 VTAIL.n577 104.615
R274 VTAIL.n584 VTAIL.n583 104.615
R275 VTAIL.n584 VTAIL.n573 104.615
R276 VTAIL.n591 VTAIL.n573 104.615
R277 VTAIL.n592 VTAIL.n591 104.615
R278 VTAIL.n592 VTAIL.n569 104.615
R279 VTAIL.n599 VTAIL.n569 104.615
R280 VTAIL.n600 VTAIL.n599 104.615
R281 VTAIL.n600 VTAIL.n565 104.615
R282 VTAIL.n607 VTAIL.n565 104.615
R283 VTAIL.n608 VTAIL.n607 104.615
R284 VTAIL.n608 VTAIL.n561 104.615
R285 VTAIL.n615 VTAIL.n561 104.615
R286 VTAIL.n616 VTAIL.n615 104.615
R287 VTAIL.n616 VTAIL.n557 104.615
R288 VTAIL.n624 VTAIL.n557 104.615
R289 VTAIL.n625 VTAIL.n624 104.615
R290 VTAIL.n626 VTAIL.n625 104.615
R291 VTAIL.n31 VTAIL.n25 104.615
R292 VTAIL.n32 VTAIL.n31 104.615
R293 VTAIL.n32 VTAIL.n21 104.615
R294 VTAIL.n39 VTAIL.n21 104.615
R295 VTAIL.n40 VTAIL.n39 104.615
R296 VTAIL.n40 VTAIL.n17 104.615
R297 VTAIL.n47 VTAIL.n17 104.615
R298 VTAIL.n48 VTAIL.n47 104.615
R299 VTAIL.n48 VTAIL.n13 104.615
R300 VTAIL.n55 VTAIL.n13 104.615
R301 VTAIL.n56 VTAIL.n55 104.615
R302 VTAIL.n56 VTAIL.n9 104.615
R303 VTAIL.n63 VTAIL.n9 104.615
R304 VTAIL.n64 VTAIL.n63 104.615
R305 VTAIL.n64 VTAIL.n5 104.615
R306 VTAIL.n72 VTAIL.n5 104.615
R307 VTAIL.n73 VTAIL.n72 104.615
R308 VTAIL.n74 VTAIL.n73 104.615
R309 VTAIL.n109 VTAIL.n103 104.615
R310 VTAIL.n110 VTAIL.n109 104.615
R311 VTAIL.n110 VTAIL.n99 104.615
R312 VTAIL.n117 VTAIL.n99 104.615
R313 VTAIL.n118 VTAIL.n117 104.615
R314 VTAIL.n118 VTAIL.n95 104.615
R315 VTAIL.n125 VTAIL.n95 104.615
R316 VTAIL.n126 VTAIL.n125 104.615
R317 VTAIL.n126 VTAIL.n91 104.615
R318 VTAIL.n133 VTAIL.n91 104.615
R319 VTAIL.n134 VTAIL.n133 104.615
R320 VTAIL.n134 VTAIL.n87 104.615
R321 VTAIL.n141 VTAIL.n87 104.615
R322 VTAIL.n142 VTAIL.n141 104.615
R323 VTAIL.n142 VTAIL.n83 104.615
R324 VTAIL.n150 VTAIL.n83 104.615
R325 VTAIL.n151 VTAIL.n150 104.615
R326 VTAIL.n152 VTAIL.n151 104.615
R327 VTAIL.n189 VTAIL.n183 104.615
R328 VTAIL.n190 VTAIL.n189 104.615
R329 VTAIL.n190 VTAIL.n179 104.615
R330 VTAIL.n197 VTAIL.n179 104.615
R331 VTAIL.n198 VTAIL.n197 104.615
R332 VTAIL.n198 VTAIL.n175 104.615
R333 VTAIL.n205 VTAIL.n175 104.615
R334 VTAIL.n206 VTAIL.n205 104.615
R335 VTAIL.n206 VTAIL.n171 104.615
R336 VTAIL.n213 VTAIL.n171 104.615
R337 VTAIL.n214 VTAIL.n213 104.615
R338 VTAIL.n214 VTAIL.n167 104.615
R339 VTAIL.n221 VTAIL.n167 104.615
R340 VTAIL.n222 VTAIL.n221 104.615
R341 VTAIL.n222 VTAIL.n163 104.615
R342 VTAIL.n230 VTAIL.n163 104.615
R343 VTAIL.n231 VTAIL.n230 104.615
R344 VTAIL.n232 VTAIL.n231 104.615
R345 VTAIL.n548 VTAIL.n547 104.615
R346 VTAIL.n547 VTAIL.n546 104.615
R347 VTAIL.n546 VTAIL.n479 104.615
R348 VTAIL.n539 VTAIL.n479 104.615
R349 VTAIL.n539 VTAIL.n538 104.615
R350 VTAIL.n538 VTAIL.n484 104.615
R351 VTAIL.n531 VTAIL.n484 104.615
R352 VTAIL.n531 VTAIL.n530 104.615
R353 VTAIL.n530 VTAIL.n488 104.615
R354 VTAIL.n523 VTAIL.n488 104.615
R355 VTAIL.n523 VTAIL.n522 104.615
R356 VTAIL.n522 VTAIL.n492 104.615
R357 VTAIL.n515 VTAIL.n492 104.615
R358 VTAIL.n515 VTAIL.n514 104.615
R359 VTAIL.n514 VTAIL.n496 104.615
R360 VTAIL.n507 VTAIL.n496 104.615
R361 VTAIL.n507 VTAIL.n506 104.615
R362 VTAIL.n506 VTAIL.n500 104.615
R363 VTAIL.n468 VTAIL.n467 104.615
R364 VTAIL.n467 VTAIL.n466 104.615
R365 VTAIL.n466 VTAIL.n399 104.615
R366 VTAIL.n459 VTAIL.n399 104.615
R367 VTAIL.n459 VTAIL.n458 104.615
R368 VTAIL.n458 VTAIL.n404 104.615
R369 VTAIL.n451 VTAIL.n404 104.615
R370 VTAIL.n451 VTAIL.n450 104.615
R371 VTAIL.n450 VTAIL.n408 104.615
R372 VTAIL.n443 VTAIL.n408 104.615
R373 VTAIL.n443 VTAIL.n442 104.615
R374 VTAIL.n442 VTAIL.n412 104.615
R375 VTAIL.n435 VTAIL.n412 104.615
R376 VTAIL.n435 VTAIL.n434 104.615
R377 VTAIL.n434 VTAIL.n416 104.615
R378 VTAIL.n427 VTAIL.n416 104.615
R379 VTAIL.n427 VTAIL.n426 104.615
R380 VTAIL.n426 VTAIL.n420 104.615
R381 VTAIL.n390 VTAIL.n389 104.615
R382 VTAIL.n389 VTAIL.n388 104.615
R383 VTAIL.n388 VTAIL.n321 104.615
R384 VTAIL.n381 VTAIL.n321 104.615
R385 VTAIL.n381 VTAIL.n380 104.615
R386 VTAIL.n380 VTAIL.n326 104.615
R387 VTAIL.n373 VTAIL.n326 104.615
R388 VTAIL.n373 VTAIL.n372 104.615
R389 VTAIL.n372 VTAIL.n330 104.615
R390 VTAIL.n365 VTAIL.n330 104.615
R391 VTAIL.n365 VTAIL.n364 104.615
R392 VTAIL.n364 VTAIL.n334 104.615
R393 VTAIL.n357 VTAIL.n334 104.615
R394 VTAIL.n357 VTAIL.n356 104.615
R395 VTAIL.n356 VTAIL.n338 104.615
R396 VTAIL.n349 VTAIL.n338 104.615
R397 VTAIL.n349 VTAIL.n348 104.615
R398 VTAIL.n348 VTAIL.n342 104.615
R399 VTAIL.n310 VTAIL.n309 104.615
R400 VTAIL.n309 VTAIL.n308 104.615
R401 VTAIL.n308 VTAIL.n241 104.615
R402 VTAIL.n301 VTAIL.n241 104.615
R403 VTAIL.n301 VTAIL.n300 104.615
R404 VTAIL.n300 VTAIL.n246 104.615
R405 VTAIL.n293 VTAIL.n246 104.615
R406 VTAIL.n293 VTAIL.n292 104.615
R407 VTAIL.n292 VTAIL.n250 104.615
R408 VTAIL.n285 VTAIL.n250 104.615
R409 VTAIL.n285 VTAIL.n284 104.615
R410 VTAIL.n284 VTAIL.n254 104.615
R411 VTAIL.n277 VTAIL.n254 104.615
R412 VTAIL.n277 VTAIL.n276 104.615
R413 VTAIL.n276 VTAIL.n258 104.615
R414 VTAIL.n269 VTAIL.n258 104.615
R415 VTAIL.n269 VTAIL.n268 104.615
R416 VTAIL.n268 VTAIL.n262 104.615
R417 VTAIL.t2 VTAIL.n577 52.3082
R418 VTAIL.t0 VTAIL.n25 52.3082
R419 VTAIL.t8 VTAIL.n103 52.3082
R420 VTAIL.t11 VTAIL.n183 52.3082
R421 VTAIL.t12 VTAIL.n500 52.3082
R422 VTAIL.t10 VTAIL.n420 52.3082
R423 VTAIL.t4 VTAIL.n342 52.3082
R424 VTAIL.t7 VTAIL.n262 52.3082
R425 VTAIL.n475 VTAIL.n474 47.6326
R426 VTAIL.n317 VTAIL.n316 47.6326
R427 VTAIL.n1 VTAIL.n0 47.6324
R428 VTAIL.n159 VTAIL.n158 47.6324
R429 VTAIL.n631 VTAIL.n630 35.4823
R430 VTAIL.n79 VTAIL.n78 35.4823
R431 VTAIL.n157 VTAIL.n156 35.4823
R432 VTAIL.n237 VTAIL.n236 35.4823
R433 VTAIL.n553 VTAIL.n552 35.4823
R434 VTAIL.n473 VTAIL.n472 35.4823
R435 VTAIL.n395 VTAIL.n394 35.4823
R436 VTAIL.n315 VTAIL.n314 35.4823
R437 VTAIL.n631 VTAIL.n553 26.9703
R438 VTAIL.n315 VTAIL.n237 26.9703
R439 VTAIL.n579 VTAIL.n578 15.6677
R440 VTAIL.n27 VTAIL.n26 15.6677
R441 VTAIL.n105 VTAIL.n104 15.6677
R442 VTAIL.n185 VTAIL.n184 15.6677
R443 VTAIL.n502 VTAIL.n501 15.6677
R444 VTAIL.n422 VTAIL.n421 15.6677
R445 VTAIL.n344 VTAIL.n343 15.6677
R446 VTAIL.n264 VTAIL.n263 15.6677
R447 VTAIL.n627 VTAIL.n556 13.1884
R448 VTAIL.n75 VTAIL.n4 13.1884
R449 VTAIL.n153 VTAIL.n82 13.1884
R450 VTAIL.n233 VTAIL.n162 13.1884
R451 VTAIL.n549 VTAIL.n478 13.1884
R452 VTAIL.n469 VTAIL.n398 13.1884
R453 VTAIL.n391 VTAIL.n320 13.1884
R454 VTAIL.n311 VTAIL.n240 13.1884
R455 VTAIL.n582 VTAIL.n581 12.8005
R456 VTAIL.n623 VTAIL.n622 12.8005
R457 VTAIL.n628 VTAIL.n554 12.8005
R458 VTAIL.n30 VTAIL.n29 12.8005
R459 VTAIL.n71 VTAIL.n70 12.8005
R460 VTAIL.n76 VTAIL.n2 12.8005
R461 VTAIL.n108 VTAIL.n107 12.8005
R462 VTAIL.n149 VTAIL.n148 12.8005
R463 VTAIL.n154 VTAIL.n80 12.8005
R464 VTAIL.n188 VTAIL.n187 12.8005
R465 VTAIL.n229 VTAIL.n228 12.8005
R466 VTAIL.n234 VTAIL.n160 12.8005
R467 VTAIL.n550 VTAIL.n476 12.8005
R468 VTAIL.n545 VTAIL.n480 12.8005
R469 VTAIL.n505 VTAIL.n504 12.8005
R470 VTAIL.n470 VTAIL.n396 12.8005
R471 VTAIL.n465 VTAIL.n400 12.8005
R472 VTAIL.n425 VTAIL.n424 12.8005
R473 VTAIL.n392 VTAIL.n318 12.8005
R474 VTAIL.n387 VTAIL.n322 12.8005
R475 VTAIL.n347 VTAIL.n346 12.8005
R476 VTAIL.n312 VTAIL.n238 12.8005
R477 VTAIL.n307 VTAIL.n242 12.8005
R478 VTAIL.n267 VTAIL.n266 12.8005
R479 VTAIL.n585 VTAIL.n576 12.0247
R480 VTAIL.n621 VTAIL.n558 12.0247
R481 VTAIL.n33 VTAIL.n24 12.0247
R482 VTAIL.n69 VTAIL.n6 12.0247
R483 VTAIL.n111 VTAIL.n102 12.0247
R484 VTAIL.n147 VTAIL.n84 12.0247
R485 VTAIL.n191 VTAIL.n182 12.0247
R486 VTAIL.n227 VTAIL.n164 12.0247
R487 VTAIL.n544 VTAIL.n481 12.0247
R488 VTAIL.n508 VTAIL.n499 12.0247
R489 VTAIL.n464 VTAIL.n401 12.0247
R490 VTAIL.n428 VTAIL.n419 12.0247
R491 VTAIL.n386 VTAIL.n323 12.0247
R492 VTAIL.n350 VTAIL.n341 12.0247
R493 VTAIL.n306 VTAIL.n243 12.0247
R494 VTAIL.n270 VTAIL.n261 12.0247
R495 VTAIL.n586 VTAIL.n574 11.249
R496 VTAIL.n618 VTAIL.n617 11.249
R497 VTAIL.n34 VTAIL.n22 11.249
R498 VTAIL.n66 VTAIL.n65 11.249
R499 VTAIL.n112 VTAIL.n100 11.249
R500 VTAIL.n144 VTAIL.n143 11.249
R501 VTAIL.n192 VTAIL.n180 11.249
R502 VTAIL.n224 VTAIL.n223 11.249
R503 VTAIL.n541 VTAIL.n540 11.249
R504 VTAIL.n509 VTAIL.n497 11.249
R505 VTAIL.n461 VTAIL.n460 11.249
R506 VTAIL.n429 VTAIL.n417 11.249
R507 VTAIL.n383 VTAIL.n382 11.249
R508 VTAIL.n351 VTAIL.n339 11.249
R509 VTAIL.n303 VTAIL.n302 11.249
R510 VTAIL.n271 VTAIL.n259 11.249
R511 VTAIL.n590 VTAIL.n589 10.4732
R512 VTAIL.n614 VTAIL.n560 10.4732
R513 VTAIL.n38 VTAIL.n37 10.4732
R514 VTAIL.n62 VTAIL.n8 10.4732
R515 VTAIL.n116 VTAIL.n115 10.4732
R516 VTAIL.n140 VTAIL.n86 10.4732
R517 VTAIL.n196 VTAIL.n195 10.4732
R518 VTAIL.n220 VTAIL.n166 10.4732
R519 VTAIL.n537 VTAIL.n483 10.4732
R520 VTAIL.n513 VTAIL.n512 10.4732
R521 VTAIL.n457 VTAIL.n403 10.4732
R522 VTAIL.n433 VTAIL.n432 10.4732
R523 VTAIL.n379 VTAIL.n325 10.4732
R524 VTAIL.n355 VTAIL.n354 10.4732
R525 VTAIL.n299 VTAIL.n245 10.4732
R526 VTAIL.n275 VTAIL.n274 10.4732
R527 VTAIL.n593 VTAIL.n572 9.69747
R528 VTAIL.n613 VTAIL.n562 9.69747
R529 VTAIL.n41 VTAIL.n20 9.69747
R530 VTAIL.n61 VTAIL.n10 9.69747
R531 VTAIL.n119 VTAIL.n98 9.69747
R532 VTAIL.n139 VTAIL.n88 9.69747
R533 VTAIL.n199 VTAIL.n178 9.69747
R534 VTAIL.n219 VTAIL.n168 9.69747
R535 VTAIL.n536 VTAIL.n485 9.69747
R536 VTAIL.n516 VTAIL.n495 9.69747
R537 VTAIL.n456 VTAIL.n405 9.69747
R538 VTAIL.n436 VTAIL.n415 9.69747
R539 VTAIL.n378 VTAIL.n327 9.69747
R540 VTAIL.n358 VTAIL.n337 9.69747
R541 VTAIL.n298 VTAIL.n247 9.69747
R542 VTAIL.n278 VTAIL.n257 9.69747
R543 VTAIL.n630 VTAIL.n629 9.45567
R544 VTAIL.n78 VTAIL.n77 9.45567
R545 VTAIL.n156 VTAIL.n155 9.45567
R546 VTAIL.n236 VTAIL.n235 9.45567
R547 VTAIL.n552 VTAIL.n551 9.45567
R548 VTAIL.n472 VTAIL.n471 9.45567
R549 VTAIL.n394 VTAIL.n393 9.45567
R550 VTAIL.n314 VTAIL.n313 9.45567
R551 VTAIL.n629 VTAIL.n628 9.3005
R552 VTAIL.n568 VTAIL.n567 9.3005
R553 VTAIL.n597 VTAIL.n596 9.3005
R554 VTAIL.n595 VTAIL.n594 9.3005
R555 VTAIL.n572 VTAIL.n571 9.3005
R556 VTAIL.n589 VTAIL.n588 9.3005
R557 VTAIL.n587 VTAIL.n586 9.3005
R558 VTAIL.n576 VTAIL.n575 9.3005
R559 VTAIL.n581 VTAIL.n580 9.3005
R560 VTAIL.n603 VTAIL.n602 9.3005
R561 VTAIL.n605 VTAIL.n604 9.3005
R562 VTAIL.n564 VTAIL.n563 9.3005
R563 VTAIL.n611 VTAIL.n610 9.3005
R564 VTAIL.n613 VTAIL.n612 9.3005
R565 VTAIL.n560 VTAIL.n559 9.3005
R566 VTAIL.n619 VTAIL.n618 9.3005
R567 VTAIL.n621 VTAIL.n620 9.3005
R568 VTAIL.n622 VTAIL.n555 9.3005
R569 VTAIL.n77 VTAIL.n76 9.3005
R570 VTAIL.n16 VTAIL.n15 9.3005
R571 VTAIL.n45 VTAIL.n44 9.3005
R572 VTAIL.n43 VTAIL.n42 9.3005
R573 VTAIL.n20 VTAIL.n19 9.3005
R574 VTAIL.n37 VTAIL.n36 9.3005
R575 VTAIL.n35 VTAIL.n34 9.3005
R576 VTAIL.n24 VTAIL.n23 9.3005
R577 VTAIL.n29 VTAIL.n28 9.3005
R578 VTAIL.n51 VTAIL.n50 9.3005
R579 VTAIL.n53 VTAIL.n52 9.3005
R580 VTAIL.n12 VTAIL.n11 9.3005
R581 VTAIL.n59 VTAIL.n58 9.3005
R582 VTAIL.n61 VTAIL.n60 9.3005
R583 VTAIL.n8 VTAIL.n7 9.3005
R584 VTAIL.n67 VTAIL.n66 9.3005
R585 VTAIL.n69 VTAIL.n68 9.3005
R586 VTAIL.n70 VTAIL.n3 9.3005
R587 VTAIL.n155 VTAIL.n154 9.3005
R588 VTAIL.n94 VTAIL.n93 9.3005
R589 VTAIL.n123 VTAIL.n122 9.3005
R590 VTAIL.n121 VTAIL.n120 9.3005
R591 VTAIL.n98 VTAIL.n97 9.3005
R592 VTAIL.n115 VTAIL.n114 9.3005
R593 VTAIL.n113 VTAIL.n112 9.3005
R594 VTAIL.n102 VTAIL.n101 9.3005
R595 VTAIL.n107 VTAIL.n106 9.3005
R596 VTAIL.n129 VTAIL.n128 9.3005
R597 VTAIL.n131 VTAIL.n130 9.3005
R598 VTAIL.n90 VTAIL.n89 9.3005
R599 VTAIL.n137 VTAIL.n136 9.3005
R600 VTAIL.n139 VTAIL.n138 9.3005
R601 VTAIL.n86 VTAIL.n85 9.3005
R602 VTAIL.n145 VTAIL.n144 9.3005
R603 VTAIL.n147 VTAIL.n146 9.3005
R604 VTAIL.n148 VTAIL.n81 9.3005
R605 VTAIL.n235 VTAIL.n234 9.3005
R606 VTAIL.n174 VTAIL.n173 9.3005
R607 VTAIL.n203 VTAIL.n202 9.3005
R608 VTAIL.n201 VTAIL.n200 9.3005
R609 VTAIL.n178 VTAIL.n177 9.3005
R610 VTAIL.n195 VTAIL.n194 9.3005
R611 VTAIL.n193 VTAIL.n192 9.3005
R612 VTAIL.n182 VTAIL.n181 9.3005
R613 VTAIL.n187 VTAIL.n186 9.3005
R614 VTAIL.n209 VTAIL.n208 9.3005
R615 VTAIL.n211 VTAIL.n210 9.3005
R616 VTAIL.n170 VTAIL.n169 9.3005
R617 VTAIL.n217 VTAIL.n216 9.3005
R618 VTAIL.n219 VTAIL.n218 9.3005
R619 VTAIL.n166 VTAIL.n165 9.3005
R620 VTAIL.n225 VTAIL.n224 9.3005
R621 VTAIL.n227 VTAIL.n226 9.3005
R622 VTAIL.n228 VTAIL.n161 9.3005
R623 VTAIL.n528 VTAIL.n527 9.3005
R624 VTAIL.n487 VTAIL.n486 9.3005
R625 VTAIL.n534 VTAIL.n533 9.3005
R626 VTAIL.n536 VTAIL.n535 9.3005
R627 VTAIL.n483 VTAIL.n482 9.3005
R628 VTAIL.n542 VTAIL.n541 9.3005
R629 VTAIL.n544 VTAIL.n543 9.3005
R630 VTAIL.n480 VTAIL.n477 9.3005
R631 VTAIL.n551 VTAIL.n550 9.3005
R632 VTAIL.n526 VTAIL.n525 9.3005
R633 VTAIL.n491 VTAIL.n490 9.3005
R634 VTAIL.n520 VTAIL.n519 9.3005
R635 VTAIL.n518 VTAIL.n517 9.3005
R636 VTAIL.n495 VTAIL.n494 9.3005
R637 VTAIL.n512 VTAIL.n511 9.3005
R638 VTAIL.n510 VTAIL.n509 9.3005
R639 VTAIL.n499 VTAIL.n498 9.3005
R640 VTAIL.n504 VTAIL.n503 9.3005
R641 VTAIL.n448 VTAIL.n447 9.3005
R642 VTAIL.n407 VTAIL.n406 9.3005
R643 VTAIL.n454 VTAIL.n453 9.3005
R644 VTAIL.n456 VTAIL.n455 9.3005
R645 VTAIL.n403 VTAIL.n402 9.3005
R646 VTAIL.n462 VTAIL.n461 9.3005
R647 VTAIL.n464 VTAIL.n463 9.3005
R648 VTAIL.n400 VTAIL.n397 9.3005
R649 VTAIL.n471 VTAIL.n470 9.3005
R650 VTAIL.n446 VTAIL.n445 9.3005
R651 VTAIL.n411 VTAIL.n410 9.3005
R652 VTAIL.n440 VTAIL.n439 9.3005
R653 VTAIL.n438 VTAIL.n437 9.3005
R654 VTAIL.n415 VTAIL.n414 9.3005
R655 VTAIL.n432 VTAIL.n431 9.3005
R656 VTAIL.n430 VTAIL.n429 9.3005
R657 VTAIL.n419 VTAIL.n418 9.3005
R658 VTAIL.n424 VTAIL.n423 9.3005
R659 VTAIL.n370 VTAIL.n369 9.3005
R660 VTAIL.n329 VTAIL.n328 9.3005
R661 VTAIL.n376 VTAIL.n375 9.3005
R662 VTAIL.n378 VTAIL.n377 9.3005
R663 VTAIL.n325 VTAIL.n324 9.3005
R664 VTAIL.n384 VTAIL.n383 9.3005
R665 VTAIL.n386 VTAIL.n385 9.3005
R666 VTAIL.n322 VTAIL.n319 9.3005
R667 VTAIL.n393 VTAIL.n392 9.3005
R668 VTAIL.n368 VTAIL.n367 9.3005
R669 VTAIL.n333 VTAIL.n332 9.3005
R670 VTAIL.n362 VTAIL.n361 9.3005
R671 VTAIL.n360 VTAIL.n359 9.3005
R672 VTAIL.n337 VTAIL.n336 9.3005
R673 VTAIL.n354 VTAIL.n353 9.3005
R674 VTAIL.n352 VTAIL.n351 9.3005
R675 VTAIL.n341 VTAIL.n340 9.3005
R676 VTAIL.n346 VTAIL.n345 9.3005
R677 VTAIL.n290 VTAIL.n289 9.3005
R678 VTAIL.n249 VTAIL.n248 9.3005
R679 VTAIL.n296 VTAIL.n295 9.3005
R680 VTAIL.n298 VTAIL.n297 9.3005
R681 VTAIL.n245 VTAIL.n244 9.3005
R682 VTAIL.n304 VTAIL.n303 9.3005
R683 VTAIL.n306 VTAIL.n305 9.3005
R684 VTAIL.n242 VTAIL.n239 9.3005
R685 VTAIL.n313 VTAIL.n312 9.3005
R686 VTAIL.n288 VTAIL.n287 9.3005
R687 VTAIL.n253 VTAIL.n252 9.3005
R688 VTAIL.n282 VTAIL.n281 9.3005
R689 VTAIL.n280 VTAIL.n279 9.3005
R690 VTAIL.n257 VTAIL.n256 9.3005
R691 VTAIL.n274 VTAIL.n273 9.3005
R692 VTAIL.n272 VTAIL.n271 9.3005
R693 VTAIL.n261 VTAIL.n260 9.3005
R694 VTAIL.n266 VTAIL.n265 9.3005
R695 VTAIL.n594 VTAIL.n570 8.92171
R696 VTAIL.n610 VTAIL.n609 8.92171
R697 VTAIL.n42 VTAIL.n18 8.92171
R698 VTAIL.n58 VTAIL.n57 8.92171
R699 VTAIL.n120 VTAIL.n96 8.92171
R700 VTAIL.n136 VTAIL.n135 8.92171
R701 VTAIL.n200 VTAIL.n176 8.92171
R702 VTAIL.n216 VTAIL.n215 8.92171
R703 VTAIL.n533 VTAIL.n532 8.92171
R704 VTAIL.n517 VTAIL.n493 8.92171
R705 VTAIL.n453 VTAIL.n452 8.92171
R706 VTAIL.n437 VTAIL.n413 8.92171
R707 VTAIL.n375 VTAIL.n374 8.92171
R708 VTAIL.n359 VTAIL.n335 8.92171
R709 VTAIL.n295 VTAIL.n294 8.92171
R710 VTAIL.n279 VTAIL.n255 8.92171
R711 VTAIL.n598 VTAIL.n597 8.14595
R712 VTAIL.n606 VTAIL.n564 8.14595
R713 VTAIL.n46 VTAIL.n45 8.14595
R714 VTAIL.n54 VTAIL.n12 8.14595
R715 VTAIL.n124 VTAIL.n123 8.14595
R716 VTAIL.n132 VTAIL.n90 8.14595
R717 VTAIL.n204 VTAIL.n203 8.14595
R718 VTAIL.n212 VTAIL.n170 8.14595
R719 VTAIL.n529 VTAIL.n487 8.14595
R720 VTAIL.n521 VTAIL.n520 8.14595
R721 VTAIL.n449 VTAIL.n407 8.14595
R722 VTAIL.n441 VTAIL.n440 8.14595
R723 VTAIL.n371 VTAIL.n329 8.14595
R724 VTAIL.n363 VTAIL.n362 8.14595
R725 VTAIL.n291 VTAIL.n249 8.14595
R726 VTAIL.n283 VTAIL.n282 8.14595
R727 VTAIL.n601 VTAIL.n568 7.3702
R728 VTAIL.n605 VTAIL.n566 7.3702
R729 VTAIL.n49 VTAIL.n16 7.3702
R730 VTAIL.n53 VTAIL.n14 7.3702
R731 VTAIL.n127 VTAIL.n94 7.3702
R732 VTAIL.n131 VTAIL.n92 7.3702
R733 VTAIL.n207 VTAIL.n174 7.3702
R734 VTAIL.n211 VTAIL.n172 7.3702
R735 VTAIL.n528 VTAIL.n489 7.3702
R736 VTAIL.n524 VTAIL.n491 7.3702
R737 VTAIL.n448 VTAIL.n409 7.3702
R738 VTAIL.n444 VTAIL.n411 7.3702
R739 VTAIL.n370 VTAIL.n331 7.3702
R740 VTAIL.n366 VTAIL.n333 7.3702
R741 VTAIL.n290 VTAIL.n251 7.3702
R742 VTAIL.n286 VTAIL.n253 7.3702
R743 VTAIL.n602 VTAIL.n601 6.59444
R744 VTAIL.n602 VTAIL.n566 6.59444
R745 VTAIL.n50 VTAIL.n49 6.59444
R746 VTAIL.n50 VTAIL.n14 6.59444
R747 VTAIL.n128 VTAIL.n127 6.59444
R748 VTAIL.n128 VTAIL.n92 6.59444
R749 VTAIL.n208 VTAIL.n207 6.59444
R750 VTAIL.n208 VTAIL.n172 6.59444
R751 VTAIL.n525 VTAIL.n489 6.59444
R752 VTAIL.n525 VTAIL.n524 6.59444
R753 VTAIL.n445 VTAIL.n409 6.59444
R754 VTAIL.n445 VTAIL.n444 6.59444
R755 VTAIL.n367 VTAIL.n331 6.59444
R756 VTAIL.n367 VTAIL.n366 6.59444
R757 VTAIL.n287 VTAIL.n251 6.59444
R758 VTAIL.n287 VTAIL.n286 6.59444
R759 VTAIL.n598 VTAIL.n568 5.81868
R760 VTAIL.n606 VTAIL.n605 5.81868
R761 VTAIL.n46 VTAIL.n16 5.81868
R762 VTAIL.n54 VTAIL.n53 5.81868
R763 VTAIL.n124 VTAIL.n94 5.81868
R764 VTAIL.n132 VTAIL.n131 5.81868
R765 VTAIL.n204 VTAIL.n174 5.81868
R766 VTAIL.n212 VTAIL.n211 5.81868
R767 VTAIL.n529 VTAIL.n528 5.81868
R768 VTAIL.n521 VTAIL.n491 5.81868
R769 VTAIL.n449 VTAIL.n448 5.81868
R770 VTAIL.n441 VTAIL.n411 5.81868
R771 VTAIL.n371 VTAIL.n370 5.81868
R772 VTAIL.n363 VTAIL.n333 5.81868
R773 VTAIL.n291 VTAIL.n290 5.81868
R774 VTAIL.n283 VTAIL.n253 5.81868
R775 VTAIL.n597 VTAIL.n570 5.04292
R776 VTAIL.n609 VTAIL.n564 5.04292
R777 VTAIL.n45 VTAIL.n18 5.04292
R778 VTAIL.n57 VTAIL.n12 5.04292
R779 VTAIL.n123 VTAIL.n96 5.04292
R780 VTAIL.n135 VTAIL.n90 5.04292
R781 VTAIL.n203 VTAIL.n176 5.04292
R782 VTAIL.n215 VTAIL.n170 5.04292
R783 VTAIL.n532 VTAIL.n487 5.04292
R784 VTAIL.n520 VTAIL.n493 5.04292
R785 VTAIL.n452 VTAIL.n407 5.04292
R786 VTAIL.n440 VTAIL.n413 5.04292
R787 VTAIL.n374 VTAIL.n329 5.04292
R788 VTAIL.n362 VTAIL.n335 5.04292
R789 VTAIL.n294 VTAIL.n249 5.04292
R790 VTAIL.n282 VTAIL.n255 5.04292
R791 VTAIL.n580 VTAIL.n579 4.38563
R792 VTAIL.n28 VTAIL.n27 4.38563
R793 VTAIL.n106 VTAIL.n105 4.38563
R794 VTAIL.n186 VTAIL.n185 4.38563
R795 VTAIL.n503 VTAIL.n502 4.38563
R796 VTAIL.n423 VTAIL.n422 4.38563
R797 VTAIL.n345 VTAIL.n344 4.38563
R798 VTAIL.n265 VTAIL.n264 4.38563
R799 VTAIL.n594 VTAIL.n593 4.26717
R800 VTAIL.n610 VTAIL.n562 4.26717
R801 VTAIL.n42 VTAIL.n41 4.26717
R802 VTAIL.n58 VTAIL.n10 4.26717
R803 VTAIL.n120 VTAIL.n119 4.26717
R804 VTAIL.n136 VTAIL.n88 4.26717
R805 VTAIL.n200 VTAIL.n199 4.26717
R806 VTAIL.n216 VTAIL.n168 4.26717
R807 VTAIL.n533 VTAIL.n485 4.26717
R808 VTAIL.n517 VTAIL.n516 4.26717
R809 VTAIL.n453 VTAIL.n405 4.26717
R810 VTAIL.n437 VTAIL.n436 4.26717
R811 VTAIL.n375 VTAIL.n327 4.26717
R812 VTAIL.n359 VTAIL.n358 4.26717
R813 VTAIL.n295 VTAIL.n247 4.26717
R814 VTAIL.n279 VTAIL.n278 4.26717
R815 VTAIL.n590 VTAIL.n572 3.49141
R816 VTAIL.n614 VTAIL.n613 3.49141
R817 VTAIL.n38 VTAIL.n20 3.49141
R818 VTAIL.n62 VTAIL.n61 3.49141
R819 VTAIL.n116 VTAIL.n98 3.49141
R820 VTAIL.n140 VTAIL.n139 3.49141
R821 VTAIL.n196 VTAIL.n178 3.49141
R822 VTAIL.n220 VTAIL.n219 3.49141
R823 VTAIL.n537 VTAIL.n536 3.49141
R824 VTAIL.n513 VTAIL.n495 3.49141
R825 VTAIL.n457 VTAIL.n456 3.49141
R826 VTAIL.n433 VTAIL.n415 3.49141
R827 VTAIL.n379 VTAIL.n378 3.49141
R828 VTAIL.n355 VTAIL.n337 3.49141
R829 VTAIL.n299 VTAIL.n298 3.49141
R830 VTAIL.n275 VTAIL.n257 3.49141
R831 VTAIL.n589 VTAIL.n574 2.71565
R832 VTAIL.n617 VTAIL.n560 2.71565
R833 VTAIL.n37 VTAIL.n22 2.71565
R834 VTAIL.n65 VTAIL.n8 2.71565
R835 VTAIL.n115 VTAIL.n100 2.71565
R836 VTAIL.n143 VTAIL.n86 2.71565
R837 VTAIL.n195 VTAIL.n180 2.71565
R838 VTAIL.n223 VTAIL.n166 2.71565
R839 VTAIL.n540 VTAIL.n483 2.71565
R840 VTAIL.n512 VTAIL.n497 2.71565
R841 VTAIL.n460 VTAIL.n403 2.71565
R842 VTAIL.n432 VTAIL.n417 2.71565
R843 VTAIL.n382 VTAIL.n325 2.71565
R844 VTAIL.n354 VTAIL.n339 2.71565
R845 VTAIL.n302 VTAIL.n245 2.71565
R846 VTAIL.n274 VTAIL.n259 2.71565
R847 VTAIL.n317 VTAIL.n315 2.4574
R848 VTAIL.n395 VTAIL.n317 2.4574
R849 VTAIL.n475 VTAIL.n473 2.4574
R850 VTAIL.n553 VTAIL.n475 2.4574
R851 VTAIL.n237 VTAIL.n159 2.4574
R852 VTAIL.n159 VTAIL.n157 2.4574
R853 VTAIL.n79 VTAIL.n1 2.4574
R854 VTAIL VTAIL.n631 2.39921
R855 VTAIL.n586 VTAIL.n585 1.93989
R856 VTAIL.n618 VTAIL.n558 1.93989
R857 VTAIL.n34 VTAIL.n33 1.93989
R858 VTAIL.n66 VTAIL.n6 1.93989
R859 VTAIL.n112 VTAIL.n111 1.93989
R860 VTAIL.n144 VTAIL.n84 1.93989
R861 VTAIL.n192 VTAIL.n191 1.93989
R862 VTAIL.n224 VTAIL.n164 1.93989
R863 VTAIL.n541 VTAIL.n481 1.93989
R864 VTAIL.n509 VTAIL.n508 1.93989
R865 VTAIL.n461 VTAIL.n401 1.93989
R866 VTAIL.n429 VTAIL.n428 1.93989
R867 VTAIL.n383 VTAIL.n323 1.93989
R868 VTAIL.n351 VTAIL.n350 1.93989
R869 VTAIL.n303 VTAIL.n243 1.93989
R870 VTAIL.n271 VTAIL.n270 1.93989
R871 VTAIL.n0 VTAIL.t6 1.40575
R872 VTAIL.n0 VTAIL.t1 1.40575
R873 VTAIL.n158 VTAIL.t15 1.40575
R874 VTAIL.n158 VTAIL.t13 1.40575
R875 VTAIL.n474 VTAIL.t14 1.40575
R876 VTAIL.n474 VTAIL.t9 1.40575
R877 VTAIL.n316 VTAIL.t5 1.40575
R878 VTAIL.n316 VTAIL.t3 1.40575
R879 VTAIL.n582 VTAIL.n576 1.16414
R880 VTAIL.n623 VTAIL.n621 1.16414
R881 VTAIL.n630 VTAIL.n554 1.16414
R882 VTAIL.n30 VTAIL.n24 1.16414
R883 VTAIL.n71 VTAIL.n69 1.16414
R884 VTAIL.n78 VTAIL.n2 1.16414
R885 VTAIL.n108 VTAIL.n102 1.16414
R886 VTAIL.n149 VTAIL.n147 1.16414
R887 VTAIL.n156 VTAIL.n80 1.16414
R888 VTAIL.n188 VTAIL.n182 1.16414
R889 VTAIL.n229 VTAIL.n227 1.16414
R890 VTAIL.n236 VTAIL.n160 1.16414
R891 VTAIL.n552 VTAIL.n476 1.16414
R892 VTAIL.n545 VTAIL.n544 1.16414
R893 VTAIL.n505 VTAIL.n499 1.16414
R894 VTAIL.n472 VTAIL.n396 1.16414
R895 VTAIL.n465 VTAIL.n464 1.16414
R896 VTAIL.n425 VTAIL.n419 1.16414
R897 VTAIL.n394 VTAIL.n318 1.16414
R898 VTAIL.n387 VTAIL.n386 1.16414
R899 VTAIL.n347 VTAIL.n341 1.16414
R900 VTAIL.n314 VTAIL.n238 1.16414
R901 VTAIL.n307 VTAIL.n306 1.16414
R902 VTAIL.n267 VTAIL.n261 1.16414
R903 VTAIL.n473 VTAIL.n395 0.470328
R904 VTAIL.n157 VTAIL.n79 0.470328
R905 VTAIL.n581 VTAIL.n578 0.388379
R906 VTAIL.n622 VTAIL.n556 0.388379
R907 VTAIL.n628 VTAIL.n627 0.388379
R908 VTAIL.n29 VTAIL.n26 0.388379
R909 VTAIL.n70 VTAIL.n4 0.388379
R910 VTAIL.n76 VTAIL.n75 0.388379
R911 VTAIL.n107 VTAIL.n104 0.388379
R912 VTAIL.n148 VTAIL.n82 0.388379
R913 VTAIL.n154 VTAIL.n153 0.388379
R914 VTAIL.n187 VTAIL.n184 0.388379
R915 VTAIL.n228 VTAIL.n162 0.388379
R916 VTAIL.n234 VTAIL.n233 0.388379
R917 VTAIL.n550 VTAIL.n549 0.388379
R918 VTAIL.n480 VTAIL.n478 0.388379
R919 VTAIL.n504 VTAIL.n501 0.388379
R920 VTAIL.n470 VTAIL.n469 0.388379
R921 VTAIL.n400 VTAIL.n398 0.388379
R922 VTAIL.n424 VTAIL.n421 0.388379
R923 VTAIL.n392 VTAIL.n391 0.388379
R924 VTAIL.n322 VTAIL.n320 0.388379
R925 VTAIL.n346 VTAIL.n343 0.388379
R926 VTAIL.n312 VTAIL.n311 0.388379
R927 VTAIL.n242 VTAIL.n240 0.388379
R928 VTAIL.n266 VTAIL.n263 0.388379
R929 VTAIL.n580 VTAIL.n575 0.155672
R930 VTAIL.n587 VTAIL.n575 0.155672
R931 VTAIL.n588 VTAIL.n587 0.155672
R932 VTAIL.n588 VTAIL.n571 0.155672
R933 VTAIL.n595 VTAIL.n571 0.155672
R934 VTAIL.n596 VTAIL.n595 0.155672
R935 VTAIL.n596 VTAIL.n567 0.155672
R936 VTAIL.n603 VTAIL.n567 0.155672
R937 VTAIL.n604 VTAIL.n603 0.155672
R938 VTAIL.n604 VTAIL.n563 0.155672
R939 VTAIL.n611 VTAIL.n563 0.155672
R940 VTAIL.n612 VTAIL.n611 0.155672
R941 VTAIL.n612 VTAIL.n559 0.155672
R942 VTAIL.n619 VTAIL.n559 0.155672
R943 VTAIL.n620 VTAIL.n619 0.155672
R944 VTAIL.n620 VTAIL.n555 0.155672
R945 VTAIL.n629 VTAIL.n555 0.155672
R946 VTAIL.n28 VTAIL.n23 0.155672
R947 VTAIL.n35 VTAIL.n23 0.155672
R948 VTAIL.n36 VTAIL.n35 0.155672
R949 VTAIL.n36 VTAIL.n19 0.155672
R950 VTAIL.n43 VTAIL.n19 0.155672
R951 VTAIL.n44 VTAIL.n43 0.155672
R952 VTAIL.n44 VTAIL.n15 0.155672
R953 VTAIL.n51 VTAIL.n15 0.155672
R954 VTAIL.n52 VTAIL.n51 0.155672
R955 VTAIL.n52 VTAIL.n11 0.155672
R956 VTAIL.n59 VTAIL.n11 0.155672
R957 VTAIL.n60 VTAIL.n59 0.155672
R958 VTAIL.n60 VTAIL.n7 0.155672
R959 VTAIL.n67 VTAIL.n7 0.155672
R960 VTAIL.n68 VTAIL.n67 0.155672
R961 VTAIL.n68 VTAIL.n3 0.155672
R962 VTAIL.n77 VTAIL.n3 0.155672
R963 VTAIL.n106 VTAIL.n101 0.155672
R964 VTAIL.n113 VTAIL.n101 0.155672
R965 VTAIL.n114 VTAIL.n113 0.155672
R966 VTAIL.n114 VTAIL.n97 0.155672
R967 VTAIL.n121 VTAIL.n97 0.155672
R968 VTAIL.n122 VTAIL.n121 0.155672
R969 VTAIL.n122 VTAIL.n93 0.155672
R970 VTAIL.n129 VTAIL.n93 0.155672
R971 VTAIL.n130 VTAIL.n129 0.155672
R972 VTAIL.n130 VTAIL.n89 0.155672
R973 VTAIL.n137 VTAIL.n89 0.155672
R974 VTAIL.n138 VTAIL.n137 0.155672
R975 VTAIL.n138 VTAIL.n85 0.155672
R976 VTAIL.n145 VTAIL.n85 0.155672
R977 VTAIL.n146 VTAIL.n145 0.155672
R978 VTAIL.n146 VTAIL.n81 0.155672
R979 VTAIL.n155 VTAIL.n81 0.155672
R980 VTAIL.n186 VTAIL.n181 0.155672
R981 VTAIL.n193 VTAIL.n181 0.155672
R982 VTAIL.n194 VTAIL.n193 0.155672
R983 VTAIL.n194 VTAIL.n177 0.155672
R984 VTAIL.n201 VTAIL.n177 0.155672
R985 VTAIL.n202 VTAIL.n201 0.155672
R986 VTAIL.n202 VTAIL.n173 0.155672
R987 VTAIL.n209 VTAIL.n173 0.155672
R988 VTAIL.n210 VTAIL.n209 0.155672
R989 VTAIL.n210 VTAIL.n169 0.155672
R990 VTAIL.n217 VTAIL.n169 0.155672
R991 VTAIL.n218 VTAIL.n217 0.155672
R992 VTAIL.n218 VTAIL.n165 0.155672
R993 VTAIL.n225 VTAIL.n165 0.155672
R994 VTAIL.n226 VTAIL.n225 0.155672
R995 VTAIL.n226 VTAIL.n161 0.155672
R996 VTAIL.n235 VTAIL.n161 0.155672
R997 VTAIL.n551 VTAIL.n477 0.155672
R998 VTAIL.n543 VTAIL.n477 0.155672
R999 VTAIL.n543 VTAIL.n542 0.155672
R1000 VTAIL.n542 VTAIL.n482 0.155672
R1001 VTAIL.n535 VTAIL.n482 0.155672
R1002 VTAIL.n535 VTAIL.n534 0.155672
R1003 VTAIL.n534 VTAIL.n486 0.155672
R1004 VTAIL.n527 VTAIL.n486 0.155672
R1005 VTAIL.n527 VTAIL.n526 0.155672
R1006 VTAIL.n526 VTAIL.n490 0.155672
R1007 VTAIL.n519 VTAIL.n490 0.155672
R1008 VTAIL.n519 VTAIL.n518 0.155672
R1009 VTAIL.n518 VTAIL.n494 0.155672
R1010 VTAIL.n511 VTAIL.n494 0.155672
R1011 VTAIL.n511 VTAIL.n510 0.155672
R1012 VTAIL.n510 VTAIL.n498 0.155672
R1013 VTAIL.n503 VTAIL.n498 0.155672
R1014 VTAIL.n471 VTAIL.n397 0.155672
R1015 VTAIL.n463 VTAIL.n397 0.155672
R1016 VTAIL.n463 VTAIL.n462 0.155672
R1017 VTAIL.n462 VTAIL.n402 0.155672
R1018 VTAIL.n455 VTAIL.n402 0.155672
R1019 VTAIL.n455 VTAIL.n454 0.155672
R1020 VTAIL.n454 VTAIL.n406 0.155672
R1021 VTAIL.n447 VTAIL.n406 0.155672
R1022 VTAIL.n447 VTAIL.n446 0.155672
R1023 VTAIL.n446 VTAIL.n410 0.155672
R1024 VTAIL.n439 VTAIL.n410 0.155672
R1025 VTAIL.n439 VTAIL.n438 0.155672
R1026 VTAIL.n438 VTAIL.n414 0.155672
R1027 VTAIL.n431 VTAIL.n414 0.155672
R1028 VTAIL.n431 VTAIL.n430 0.155672
R1029 VTAIL.n430 VTAIL.n418 0.155672
R1030 VTAIL.n423 VTAIL.n418 0.155672
R1031 VTAIL.n393 VTAIL.n319 0.155672
R1032 VTAIL.n385 VTAIL.n319 0.155672
R1033 VTAIL.n385 VTAIL.n384 0.155672
R1034 VTAIL.n384 VTAIL.n324 0.155672
R1035 VTAIL.n377 VTAIL.n324 0.155672
R1036 VTAIL.n377 VTAIL.n376 0.155672
R1037 VTAIL.n376 VTAIL.n328 0.155672
R1038 VTAIL.n369 VTAIL.n328 0.155672
R1039 VTAIL.n369 VTAIL.n368 0.155672
R1040 VTAIL.n368 VTAIL.n332 0.155672
R1041 VTAIL.n361 VTAIL.n332 0.155672
R1042 VTAIL.n361 VTAIL.n360 0.155672
R1043 VTAIL.n360 VTAIL.n336 0.155672
R1044 VTAIL.n353 VTAIL.n336 0.155672
R1045 VTAIL.n353 VTAIL.n352 0.155672
R1046 VTAIL.n352 VTAIL.n340 0.155672
R1047 VTAIL.n345 VTAIL.n340 0.155672
R1048 VTAIL.n313 VTAIL.n239 0.155672
R1049 VTAIL.n305 VTAIL.n239 0.155672
R1050 VTAIL.n305 VTAIL.n304 0.155672
R1051 VTAIL.n304 VTAIL.n244 0.155672
R1052 VTAIL.n297 VTAIL.n244 0.155672
R1053 VTAIL.n297 VTAIL.n296 0.155672
R1054 VTAIL.n296 VTAIL.n248 0.155672
R1055 VTAIL.n289 VTAIL.n248 0.155672
R1056 VTAIL.n289 VTAIL.n288 0.155672
R1057 VTAIL.n288 VTAIL.n252 0.155672
R1058 VTAIL.n281 VTAIL.n252 0.155672
R1059 VTAIL.n281 VTAIL.n280 0.155672
R1060 VTAIL.n280 VTAIL.n256 0.155672
R1061 VTAIL.n273 VTAIL.n256 0.155672
R1062 VTAIL.n273 VTAIL.n272 0.155672
R1063 VTAIL.n272 VTAIL.n260 0.155672
R1064 VTAIL.n265 VTAIL.n260 0.155672
R1065 VTAIL VTAIL.n1 0.0586897
R1066 VDD1 VDD1.n0 65.598
R1067 VDD1.n3 VDD1.n2 65.4843
R1068 VDD1.n3 VDD1.n1 65.4843
R1069 VDD1.n5 VDD1.n4 64.3112
R1070 VDD1.n5 VDD1.n3 47.5009
R1071 VDD1.n4 VDD1.t3 1.40575
R1072 VDD1.n4 VDD1.t7 1.40575
R1073 VDD1.n0 VDD1.t1 1.40575
R1074 VDD1.n0 VDD1.t2 1.40575
R1075 VDD1.n2 VDD1.t4 1.40575
R1076 VDD1.n2 VDD1.t6 1.40575
R1077 VDD1.n1 VDD1.t5 1.40575
R1078 VDD1.n1 VDD1.t0 1.40575
R1079 VDD1 VDD1.n5 1.17076
R1080 B.n729 B.n149 585
R1081 B.n149 B.n92 585
R1082 B.n731 B.n730 585
R1083 B.n733 B.n148 585
R1084 B.n736 B.n735 585
R1085 B.n737 B.n147 585
R1086 B.n739 B.n738 585
R1087 B.n741 B.n146 585
R1088 B.n744 B.n743 585
R1089 B.n745 B.n145 585
R1090 B.n747 B.n746 585
R1091 B.n749 B.n144 585
R1092 B.n752 B.n751 585
R1093 B.n753 B.n143 585
R1094 B.n755 B.n754 585
R1095 B.n757 B.n142 585
R1096 B.n760 B.n759 585
R1097 B.n761 B.n141 585
R1098 B.n763 B.n762 585
R1099 B.n765 B.n140 585
R1100 B.n768 B.n767 585
R1101 B.n769 B.n139 585
R1102 B.n771 B.n770 585
R1103 B.n773 B.n138 585
R1104 B.n776 B.n775 585
R1105 B.n777 B.n137 585
R1106 B.n779 B.n778 585
R1107 B.n781 B.n136 585
R1108 B.n784 B.n783 585
R1109 B.n785 B.n135 585
R1110 B.n787 B.n786 585
R1111 B.n789 B.n134 585
R1112 B.n792 B.n791 585
R1113 B.n793 B.n133 585
R1114 B.n795 B.n794 585
R1115 B.n797 B.n132 585
R1116 B.n800 B.n799 585
R1117 B.n801 B.n131 585
R1118 B.n803 B.n802 585
R1119 B.n805 B.n130 585
R1120 B.n808 B.n807 585
R1121 B.n809 B.n129 585
R1122 B.n811 B.n810 585
R1123 B.n813 B.n128 585
R1124 B.n816 B.n815 585
R1125 B.n817 B.n127 585
R1126 B.n819 B.n818 585
R1127 B.n821 B.n126 585
R1128 B.n824 B.n823 585
R1129 B.n826 B.n123 585
R1130 B.n828 B.n827 585
R1131 B.n830 B.n122 585
R1132 B.n833 B.n832 585
R1133 B.n834 B.n121 585
R1134 B.n836 B.n835 585
R1135 B.n838 B.n120 585
R1136 B.n841 B.n840 585
R1137 B.n842 B.n117 585
R1138 B.n845 B.n844 585
R1139 B.n847 B.n116 585
R1140 B.n850 B.n849 585
R1141 B.n851 B.n115 585
R1142 B.n853 B.n852 585
R1143 B.n855 B.n114 585
R1144 B.n858 B.n857 585
R1145 B.n859 B.n113 585
R1146 B.n861 B.n860 585
R1147 B.n863 B.n112 585
R1148 B.n866 B.n865 585
R1149 B.n867 B.n111 585
R1150 B.n869 B.n868 585
R1151 B.n871 B.n110 585
R1152 B.n874 B.n873 585
R1153 B.n875 B.n109 585
R1154 B.n877 B.n876 585
R1155 B.n879 B.n108 585
R1156 B.n882 B.n881 585
R1157 B.n883 B.n107 585
R1158 B.n885 B.n884 585
R1159 B.n887 B.n106 585
R1160 B.n890 B.n889 585
R1161 B.n891 B.n105 585
R1162 B.n893 B.n892 585
R1163 B.n895 B.n104 585
R1164 B.n898 B.n897 585
R1165 B.n899 B.n103 585
R1166 B.n901 B.n900 585
R1167 B.n903 B.n102 585
R1168 B.n906 B.n905 585
R1169 B.n907 B.n101 585
R1170 B.n909 B.n908 585
R1171 B.n911 B.n100 585
R1172 B.n914 B.n913 585
R1173 B.n915 B.n99 585
R1174 B.n917 B.n916 585
R1175 B.n919 B.n98 585
R1176 B.n922 B.n921 585
R1177 B.n923 B.n97 585
R1178 B.n925 B.n924 585
R1179 B.n927 B.n96 585
R1180 B.n930 B.n929 585
R1181 B.n931 B.n95 585
R1182 B.n933 B.n932 585
R1183 B.n935 B.n94 585
R1184 B.n938 B.n937 585
R1185 B.n939 B.n93 585
R1186 B.n728 B.n91 585
R1187 B.n942 B.n91 585
R1188 B.n727 B.n90 585
R1189 B.n943 B.n90 585
R1190 B.n726 B.n89 585
R1191 B.n944 B.n89 585
R1192 B.n725 B.n724 585
R1193 B.n724 B.n85 585
R1194 B.n723 B.n84 585
R1195 B.n950 B.n84 585
R1196 B.n722 B.n83 585
R1197 B.n951 B.n83 585
R1198 B.n721 B.n82 585
R1199 B.n952 B.n82 585
R1200 B.n720 B.n719 585
R1201 B.n719 B.n81 585
R1202 B.n718 B.n77 585
R1203 B.n958 B.n77 585
R1204 B.n717 B.n76 585
R1205 B.n959 B.n76 585
R1206 B.n716 B.n75 585
R1207 B.n960 B.n75 585
R1208 B.n715 B.n714 585
R1209 B.n714 B.n71 585
R1210 B.n713 B.n70 585
R1211 B.n966 B.n70 585
R1212 B.n712 B.n69 585
R1213 B.n967 B.n69 585
R1214 B.n711 B.n68 585
R1215 B.n968 B.n68 585
R1216 B.n710 B.n709 585
R1217 B.n709 B.n64 585
R1218 B.n708 B.n63 585
R1219 B.n974 B.n63 585
R1220 B.n707 B.n62 585
R1221 B.n975 B.n62 585
R1222 B.n706 B.n61 585
R1223 B.n976 B.n61 585
R1224 B.n705 B.n704 585
R1225 B.n704 B.n60 585
R1226 B.n703 B.n56 585
R1227 B.n982 B.n56 585
R1228 B.n702 B.n55 585
R1229 B.n983 B.n55 585
R1230 B.n701 B.n54 585
R1231 B.n984 B.n54 585
R1232 B.n700 B.n699 585
R1233 B.n699 B.n50 585
R1234 B.n698 B.n49 585
R1235 B.n990 B.n49 585
R1236 B.n697 B.n48 585
R1237 B.n991 B.n48 585
R1238 B.n696 B.n47 585
R1239 B.n992 B.n47 585
R1240 B.n695 B.n694 585
R1241 B.n694 B.n46 585
R1242 B.n693 B.n42 585
R1243 B.n998 B.n42 585
R1244 B.n692 B.n41 585
R1245 B.n999 B.n41 585
R1246 B.n691 B.n40 585
R1247 B.n1000 B.n40 585
R1248 B.n690 B.n689 585
R1249 B.n689 B.n36 585
R1250 B.n688 B.n35 585
R1251 B.n1006 B.n35 585
R1252 B.n687 B.n34 585
R1253 B.n1007 B.n34 585
R1254 B.n686 B.n33 585
R1255 B.n1008 B.n33 585
R1256 B.n685 B.n684 585
R1257 B.n684 B.n32 585
R1258 B.n683 B.n28 585
R1259 B.n1014 B.n28 585
R1260 B.n682 B.n27 585
R1261 B.n1015 B.n27 585
R1262 B.n681 B.n26 585
R1263 B.n1016 B.n26 585
R1264 B.n680 B.n679 585
R1265 B.n679 B.n22 585
R1266 B.n678 B.n21 585
R1267 B.n1022 B.n21 585
R1268 B.n677 B.n20 585
R1269 B.n1023 B.n20 585
R1270 B.n676 B.n19 585
R1271 B.n1024 B.n19 585
R1272 B.n675 B.n674 585
R1273 B.n674 B.n15 585
R1274 B.n673 B.n14 585
R1275 B.n1030 B.n14 585
R1276 B.n672 B.n13 585
R1277 B.n1031 B.n13 585
R1278 B.n671 B.n12 585
R1279 B.n1032 B.n12 585
R1280 B.n670 B.n669 585
R1281 B.n669 B.n8 585
R1282 B.n668 B.n7 585
R1283 B.n1038 B.n7 585
R1284 B.n667 B.n6 585
R1285 B.n1039 B.n6 585
R1286 B.n666 B.n5 585
R1287 B.n1040 B.n5 585
R1288 B.n665 B.n664 585
R1289 B.n664 B.n4 585
R1290 B.n663 B.n150 585
R1291 B.n663 B.n662 585
R1292 B.n653 B.n151 585
R1293 B.n152 B.n151 585
R1294 B.n655 B.n654 585
R1295 B.n656 B.n655 585
R1296 B.n652 B.n157 585
R1297 B.n157 B.n156 585
R1298 B.n651 B.n650 585
R1299 B.n650 B.n649 585
R1300 B.n159 B.n158 585
R1301 B.n160 B.n159 585
R1302 B.n642 B.n641 585
R1303 B.n643 B.n642 585
R1304 B.n640 B.n165 585
R1305 B.n165 B.n164 585
R1306 B.n639 B.n638 585
R1307 B.n638 B.n637 585
R1308 B.n167 B.n166 585
R1309 B.n168 B.n167 585
R1310 B.n630 B.n629 585
R1311 B.n631 B.n630 585
R1312 B.n628 B.n173 585
R1313 B.n173 B.n172 585
R1314 B.n627 B.n626 585
R1315 B.n626 B.n625 585
R1316 B.n175 B.n174 585
R1317 B.n618 B.n175 585
R1318 B.n617 B.n616 585
R1319 B.n619 B.n617 585
R1320 B.n615 B.n180 585
R1321 B.n180 B.n179 585
R1322 B.n614 B.n613 585
R1323 B.n613 B.n612 585
R1324 B.n182 B.n181 585
R1325 B.n183 B.n182 585
R1326 B.n605 B.n604 585
R1327 B.n606 B.n605 585
R1328 B.n603 B.n188 585
R1329 B.n188 B.n187 585
R1330 B.n602 B.n601 585
R1331 B.n601 B.n600 585
R1332 B.n190 B.n189 585
R1333 B.n593 B.n190 585
R1334 B.n592 B.n591 585
R1335 B.n594 B.n592 585
R1336 B.n590 B.n195 585
R1337 B.n195 B.n194 585
R1338 B.n589 B.n588 585
R1339 B.n588 B.n587 585
R1340 B.n197 B.n196 585
R1341 B.n198 B.n197 585
R1342 B.n580 B.n579 585
R1343 B.n581 B.n580 585
R1344 B.n578 B.n203 585
R1345 B.n203 B.n202 585
R1346 B.n577 B.n576 585
R1347 B.n576 B.n575 585
R1348 B.n205 B.n204 585
R1349 B.n568 B.n205 585
R1350 B.n567 B.n566 585
R1351 B.n569 B.n567 585
R1352 B.n565 B.n210 585
R1353 B.n210 B.n209 585
R1354 B.n564 B.n563 585
R1355 B.n563 B.n562 585
R1356 B.n212 B.n211 585
R1357 B.n213 B.n212 585
R1358 B.n555 B.n554 585
R1359 B.n556 B.n555 585
R1360 B.n553 B.n218 585
R1361 B.n218 B.n217 585
R1362 B.n552 B.n551 585
R1363 B.n551 B.n550 585
R1364 B.n220 B.n219 585
R1365 B.n221 B.n220 585
R1366 B.n543 B.n542 585
R1367 B.n544 B.n543 585
R1368 B.n541 B.n226 585
R1369 B.n226 B.n225 585
R1370 B.n540 B.n539 585
R1371 B.n539 B.n538 585
R1372 B.n228 B.n227 585
R1373 B.n531 B.n228 585
R1374 B.n530 B.n529 585
R1375 B.n532 B.n530 585
R1376 B.n528 B.n233 585
R1377 B.n233 B.n232 585
R1378 B.n527 B.n526 585
R1379 B.n526 B.n525 585
R1380 B.n235 B.n234 585
R1381 B.n236 B.n235 585
R1382 B.n518 B.n517 585
R1383 B.n519 B.n518 585
R1384 B.n516 B.n241 585
R1385 B.n241 B.n240 585
R1386 B.n515 B.n514 585
R1387 B.n514 B.n513 585
R1388 B.n510 B.n245 585
R1389 B.n509 B.n508 585
R1390 B.n506 B.n246 585
R1391 B.n506 B.n244 585
R1392 B.n505 B.n504 585
R1393 B.n503 B.n502 585
R1394 B.n501 B.n248 585
R1395 B.n499 B.n498 585
R1396 B.n497 B.n249 585
R1397 B.n496 B.n495 585
R1398 B.n493 B.n250 585
R1399 B.n491 B.n490 585
R1400 B.n489 B.n251 585
R1401 B.n488 B.n487 585
R1402 B.n485 B.n252 585
R1403 B.n483 B.n482 585
R1404 B.n481 B.n253 585
R1405 B.n480 B.n479 585
R1406 B.n477 B.n254 585
R1407 B.n475 B.n474 585
R1408 B.n473 B.n255 585
R1409 B.n472 B.n471 585
R1410 B.n469 B.n256 585
R1411 B.n467 B.n466 585
R1412 B.n465 B.n257 585
R1413 B.n464 B.n463 585
R1414 B.n461 B.n258 585
R1415 B.n459 B.n458 585
R1416 B.n457 B.n259 585
R1417 B.n456 B.n455 585
R1418 B.n453 B.n260 585
R1419 B.n451 B.n450 585
R1420 B.n449 B.n261 585
R1421 B.n448 B.n447 585
R1422 B.n445 B.n262 585
R1423 B.n443 B.n442 585
R1424 B.n441 B.n263 585
R1425 B.n440 B.n439 585
R1426 B.n437 B.n264 585
R1427 B.n435 B.n434 585
R1428 B.n433 B.n265 585
R1429 B.n432 B.n431 585
R1430 B.n429 B.n266 585
R1431 B.n427 B.n426 585
R1432 B.n425 B.n267 585
R1433 B.n424 B.n423 585
R1434 B.n421 B.n268 585
R1435 B.n419 B.n418 585
R1436 B.n417 B.n269 585
R1437 B.n415 B.n414 585
R1438 B.n412 B.n272 585
R1439 B.n410 B.n409 585
R1440 B.n408 B.n273 585
R1441 B.n407 B.n406 585
R1442 B.n404 B.n274 585
R1443 B.n402 B.n401 585
R1444 B.n400 B.n275 585
R1445 B.n399 B.n398 585
R1446 B.n396 B.n395 585
R1447 B.n394 B.n393 585
R1448 B.n392 B.n280 585
R1449 B.n390 B.n389 585
R1450 B.n388 B.n281 585
R1451 B.n387 B.n386 585
R1452 B.n384 B.n282 585
R1453 B.n382 B.n381 585
R1454 B.n380 B.n283 585
R1455 B.n379 B.n378 585
R1456 B.n376 B.n284 585
R1457 B.n374 B.n373 585
R1458 B.n372 B.n285 585
R1459 B.n371 B.n370 585
R1460 B.n368 B.n286 585
R1461 B.n366 B.n365 585
R1462 B.n364 B.n287 585
R1463 B.n363 B.n362 585
R1464 B.n360 B.n288 585
R1465 B.n358 B.n357 585
R1466 B.n356 B.n289 585
R1467 B.n355 B.n354 585
R1468 B.n352 B.n290 585
R1469 B.n350 B.n349 585
R1470 B.n348 B.n291 585
R1471 B.n347 B.n346 585
R1472 B.n344 B.n292 585
R1473 B.n342 B.n341 585
R1474 B.n340 B.n293 585
R1475 B.n339 B.n338 585
R1476 B.n336 B.n294 585
R1477 B.n334 B.n333 585
R1478 B.n332 B.n295 585
R1479 B.n331 B.n330 585
R1480 B.n328 B.n296 585
R1481 B.n326 B.n325 585
R1482 B.n324 B.n297 585
R1483 B.n323 B.n322 585
R1484 B.n320 B.n298 585
R1485 B.n318 B.n317 585
R1486 B.n316 B.n299 585
R1487 B.n315 B.n314 585
R1488 B.n312 B.n300 585
R1489 B.n310 B.n309 585
R1490 B.n308 B.n301 585
R1491 B.n307 B.n306 585
R1492 B.n304 B.n302 585
R1493 B.n243 B.n242 585
R1494 B.n512 B.n511 585
R1495 B.n513 B.n512 585
R1496 B.n239 B.n238 585
R1497 B.n240 B.n239 585
R1498 B.n521 B.n520 585
R1499 B.n520 B.n519 585
R1500 B.n522 B.n237 585
R1501 B.n237 B.n236 585
R1502 B.n524 B.n523 585
R1503 B.n525 B.n524 585
R1504 B.n231 B.n230 585
R1505 B.n232 B.n231 585
R1506 B.n534 B.n533 585
R1507 B.n533 B.n532 585
R1508 B.n535 B.n229 585
R1509 B.n531 B.n229 585
R1510 B.n537 B.n536 585
R1511 B.n538 B.n537 585
R1512 B.n224 B.n223 585
R1513 B.n225 B.n224 585
R1514 B.n546 B.n545 585
R1515 B.n545 B.n544 585
R1516 B.n547 B.n222 585
R1517 B.n222 B.n221 585
R1518 B.n549 B.n548 585
R1519 B.n550 B.n549 585
R1520 B.n216 B.n215 585
R1521 B.n217 B.n216 585
R1522 B.n558 B.n557 585
R1523 B.n557 B.n556 585
R1524 B.n559 B.n214 585
R1525 B.n214 B.n213 585
R1526 B.n561 B.n560 585
R1527 B.n562 B.n561 585
R1528 B.n208 B.n207 585
R1529 B.n209 B.n208 585
R1530 B.n571 B.n570 585
R1531 B.n570 B.n569 585
R1532 B.n572 B.n206 585
R1533 B.n568 B.n206 585
R1534 B.n574 B.n573 585
R1535 B.n575 B.n574 585
R1536 B.n201 B.n200 585
R1537 B.n202 B.n201 585
R1538 B.n583 B.n582 585
R1539 B.n582 B.n581 585
R1540 B.n584 B.n199 585
R1541 B.n199 B.n198 585
R1542 B.n586 B.n585 585
R1543 B.n587 B.n586 585
R1544 B.n193 B.n192 585
R1545 B.n194 B.n193 585
R1546 B.n596 B.n595 585
R1547 B.n595 B.n594 585
R1548 B.n597 B.n191 585
R1549 B.n593 B.n191 585
R1550 B.n599 B.n598 585
R1551 B.n600 B.n599 585
R1552 B.n186 B.n185 585
R1553 B.n187 B.n186 585
R1554 B.n608 B.n607 585
R1555 B.n607 B.n606 585
R1556 B.n609 B.n184 585
R1557 B.n184 B.n183 585
R1558 B.n611 B.n610 585
R1559 B.n612 B.n611 585
R1560 B.n178 B.n177 585
R1561 B.n179 B.n178 585
R1562 B.n621 B.n620 585
R1563 B.n620 B.n619 585
R1564 B.n622 B.n176 585
R1565 B.n618 B.n176 585
R1566 B.n624 B.n623 585
R1567 B.n625 B.n624 585
R1568 B.n171 B.n170 585
R1569 B.n172 B.n171 585
R1570 B.n633 B.n632 585
R1571 B.n632 B.n631 585
R1572 B.n634 B.n169 585
R1573 B.n169 B.n168 585
R1574 B.n636 B.n635 585
R1575 B.n637 B.n636 585
R1576 B.n163 B.n162 585
R1577 B.n164 B.n163 585
R1578 B.n645 B.n644 585
R1579 B.n644 B.n643 585
R1580 B.n646 B.n161 585
R1581 B.n161 B.n160 585
R1582 B.n648 B.n647 585
R1583 B.n649 B.n648 585
R1584 B.n155 B.n154 585
R1585 B.n156 B.n155 585
R1586 B.n658 B.n657 585
R1587 B.n657 B.n656 585
R1588 B.n659 B.n153 585
R1589 B.n153 B.n152 585
R1590 B.n661 B.n660 585
R1591 B.n662 B.n661 585
R1592 B.n2 B.n0 585
R1593 B.n4 B.n2 585
R1594 B.n3 B.n1 585
R1595 B.n1039 B.n3 585
R1596 B.n1037 B.n1036 585
R1597 B.n1038 B.n1037 585
R1598 B.n1035 B.n9 585
R1599 B.n9 B.n8 585
R1600 B.n1034 B.n1033 585
R1601 B.n1033 B.n1032 585
R1602 B.n11 B.n10 585
R1603 B.n1031 B.n11 585
R1604 B.n1029 B.n1028 585
R1605 B.n1030 B.n1029 585
R1606 B.n1027 B.n16 585
R1607 B.n16 B.n15 585
R1608 B.n1026 B.n1025 585
R1609 B.n1025 B.n1024 585
R1610 B.n18 B.n17 585
R1611 B.n1023 B.n18 585
R1612 B.n1021 B.n1020 585
R1613 B.n1022 B.n1021 585
R1614 B.n1019 B.n23 585
R1615 B.n23 B.n22 585
R1616 B.n1018 B.n1017 585
R1617 B.n1017 B.n1016 585
R1618 B.n25 B.n24 585
R1619 B.n1015 B.n25 585
R1620 B.n1013 B.n1012 585
R1621 B.n1014 B.n1013 585
R1622 B.n1011 B.n29 585
R1623 B.n32 B.n29 585
R1624 B.n1010 B.n1009 585
R1625 B.n1009 B.n1008 585
R1626 B.n31 B.n30 585
R1627 B.n1007 B.n31 585
R1628 B.n1005 B.n1004 585
R1629 B.n1006 B.n1005 585
R1630 B.n1003 B.n37 585
R1631 B.n37 B.n36 585
R1632 B.n1002 B.n1001 585
R1633 B.n1001 B.n1000 585
R1634 B.n39 B.n38 585
R1635 B.n999 B.n39 585
R1636 B.n997 B.n996 585
R1637 B.n998 B.n997 585
R1638 B.n995 B.n43 585
R1639 B.n46 B.n43 585
R1640 B.n994 B.n993 585
R1641 B.n993 B.n992 585
R1642 B.n45 B.n44 585
R1643 B.n991 B.n45 585
R1644 B.n989 B.n988 585
R1645 B.n990 B.n989 585
R1646 B.n987 B.n51 585
R1647 B.n51 B.n50 585
R1648 B.n986 B.n985 585
R1649 B.n985 B.n984 585
R1650 B.n53 B.n52 585
R1651 B.n983 B.n53 585
R1652 B.n981 B.n980 585
R1653 B.n982 B.n981 585
R1654 B.n979 B.n57 585
R1655 B.n60 B.n57 585
R1656 B.n978 B.n977 585
R1657 B.n977 B.n976 585
R1658 B.n59 B.n58 585
R1659 B.n975 B.n59 585
R1660 B.n973 B.n972 585
R1661 B.n974 B.n973 585
R1662 B.n971 B.n65 585
R1663 B.n65 B.n64 585
R1664 B.n970 B.n969 585
R1665 B.n969 B.n968 585
R1666 B.n67 B.n66 585
R1667 B.n967 B.n67 585
R1668 B.n965 B.n964 585
R1669 B.n966 B.n965 585
R1670 B.n963 B.n72 585
R1671 B.n72 B.n71 585
R1672 B.n962 B.n961 585
R1673 B.n961 B.n960 585
R1674 B.n74 B.n73 585
R1675 B.n959 B.n74 585
R1676 B.n957 B.n956 585
R1677 B.n958 B.n957 585
R1678 B.n955 B.n78 585
R1679 B.n81 B.n78 585
R1680 B.n954 B.n953 585
R1681 B.n953 B.n952 585
R1682 B.n80 B.n79 585
R1683 B.n951 B.n80 585
R1684 B.n949 B.n948 585
R1685 B.n950 B.n949 585
R1686 B.n947 B.n86 585
R1687 B.n86 B.n85 585
R1688 B.n946 B.n945 585
R1689 B.n945 B.n944 585
R1690 B.n88 B.n87 585
R1691 B.n943 B.n88 585
R1692 B.n941 B.n940 585
R1693 B.n942 B.n941 585
R1694 B.n1042 B.n1041 585
R1695 B.n1041 B.n1040 585
R1696 B.n512 B.n245 511.721
R1697 B.n941 B.n93 511.721
R1698 B.n514 B.n243 511.721
R1699 B.n149 B.n91 511.721
R1700 B.n276 B.t21 373.387
R1701 B.n124 B.t10 373.387
R1702 B.n270 B.t15 373.387
R1703 B.n118 B.t17 373.387
R1704 B.n276 B.t19 342.673
R1705 B.n270 B.t12 342.673
R1706 B.n118 B.t16 342.673
R1707 B.n124 B.t8 342.673
R1708 B.n277 B.t20 318.115
R1709 B.n125 B.t11 318.115
R1710 B.n271 B.t14 318.115
R1711 B.n119 B.t18 318.115
R1712 B.n732 B.n92 256.663
R1713 B.n734 B.n92 256.663
R1714 B.n740 B.n92 256.663
R1715 B.n742 B.n92 256.663
R1716 B.n748 B.n92 256.663
R1717 B.n750 B.n92 256.663
R1718 B.n756 B.n92 256.663
R1719 B.n758 B.n92 256.663
R1720 B.n764 B.n92 256.663
R1721 B.n766 B.n92 256.663
R1722 B.n772 B.n92 256.663
R1723 B.n774 B.n92 256.663
R1724 B.n780 B.n92 256.663
R1725 B.n782 B.n92 256.663
R1726 B.n788 B.n92 256.663
R1727 B.n790 B.n92 256.663
R1728 B.n796 B.n92 256.663
R1729 B.n798 B.n92 256.663
R1730 B.n804 B.n92 256.663
R1731 B.n806 B.n92 256.663
R1732 B.n812 B.n92 256.663
R1733 B.n814 B.n92 256.663
R1734 B.n820 B.n92 256.663
R1735 B.n822 B.n92 256.663
R1736 B.n829 B.n92 256.663
R1737 B.n831 B.n92 256.663
R1738 B.n837 B.n92 256.663
R1739 B.n839 B.n92 256.663
R1740 B.n846 B.n92 256.663
R1741 B.n848 B.n92 256.663
R1742 B.n854 B.n92 256.663
R1743 B.n856 B.n92 256.663
R1744 B.n862 B.n92 256.663
R1745 B.n864 B.n92 256.663
R1746 B.n870 B.n92 256.663
R1747 B.n872 B.n92 256.663
R1748 B.n878 B.n92 256.663
R1749 B.n880 B.n92 256.663
R1750 B.n886 B.n92 256.663
R1751 B.n888 B.n92 256.663
R1752 B.n894 B.n92 256.663
R1753 B.n896 B.n92 256.663
R1754 B.n902 B.n92 256.663
R1755 B.n904 B.n92 256.663
R1756 B.n910 B.n92 256.663
R1757 B.n912 B.n92 256.663
R1758 B.n918 B.n92 256.663
R1759 B.n920 B.n92 256.663
R1760 B.n926 B.n92 256.663
R1761 B.n928 B.n92 256.663
R1762 B.n934 B.n92 256.663
R1763 B.n936 B.n92 256.663
R1764 B.n507 B.n244 256.663
R1765 B.n247 B.n244 256.663
R1766 B.n500 B.n244 256.663
R1767 B.n494 B.n244 256.663
R1768 B.n492 B.n244 256.663
R1769 B.n486 B.n244 256.663
R1770 B.n484 B.n244 256.663
R1771 B.n478 B.n244 256.663
R1772 B.n476 B.n244 256.663
R1773 B.n470 B.n244 256.663
R1774 B.n468 B.n244 256.663
R1775 B.n462 B.n244 256.663
R1776 B.n460 B.n244 256.663
R1777 B.n454 B.n244 256.663
R1778 B.n452 B.n244 256.663
R1779 B.n446 B.n244 256.663
R1780 B.n444 B.n244 256.663
R1781 B.n438 B.n244 256.663
R1782 B.n436 B.n244 256.663
R1783 B.n430 B.n244 256.663
R1784 B.n428 B.n244 256.663
R1785 B.n422 B.n244 256.663
R1786 B.n420 B.n244 256.663
R1787 B.n413 B.n244 256.663
R1788 B.n411 B.n244 256.663
R1789 B.n405 B.n244 256.663
R1790 B.n403 B.n244 256.663
R1791 B.n397 B.n244 256.663
R1792 B.n279 B.n244 256.663
R1793 B.n391 B.n244 256.663
R1794 B.n385 B.n244 256.663
R1795 B.n383 B.n244 256.663
R1796 B.n377 B.n244 256.663
R1797 B.n375 B.n244 256.663
R1798 B.n369 B.n244 256.663
R1799 B.n367 B.n244 256.663
R1800 B.n361 B.n244 256.663
R1801 B.n359 B.n244 256.663
R1802 B.n353 B.n244 256.663
R1803 B.n351 B.n244 256.663
R1804 B.n345 B.n244 256.663
R1805 B.n343 B.n244 256.663
R1806 B.n337 B.n244 256.663
R1807 B.n335 B.n244 256.663
R1808 B.n329 B.n244 256.663
R1809 B.n327 B.n244 256.663
R1810 B.n321 B.n244 256.663
R1811 B.n319 B.n244 256.663
R1812 B.n313 B.n244 256.663
R1813 B.n311 B.n244 256.663
R1814 B.n305 B.n244 256.663
R1815 B.n303 B.n244 256.663
R1816 B.n512 B.n239 163.367
R1817 B.n520 B.n239 163.367
R1818 B.n520 B.n237 163.367
R1819 B.n524 B.n237 163.367
R1820 B.n524 B.n231 163.367
R1821 B.n533 B.n231 163.367
R1822 B.n533 B.n229 163.367
R1823 B.n537 B.n229 163.367
R1824 B.n537 B.n224 163.367
R1825 B.n545 B.n224 163.367
R1826 B.n545 B.n222 163.367
R1827 B.n549 B.n222 163.367
R1828 B.n549 B.n216 163.367
R1829 B.n557 B.n216 163.367
R1830 B.n557 B.n214 163.367
R1831 B.n561 B.n214 163.367
R1832 B.n561 B.n208 163.367
R1833 B.n570 B.n208 163.367
R1834 B.n570 B.n206 163.367
R1835 B.n574 B.n206 163.367
R1836 B.n574 B.n201 163.367
R1837 B.n582 B.n201 163.367
R1838 B.n582 B.n199 163.367
R1839 B.n586 B.n199 163.367
R1840 B.n586 B.n193 163.367
R1841 B.n595 B.n193 163.367
R1842 B.n595 B.n191 163.367
R1843 B.n599 B.n191 163.367
R1844 B.n599 B.n186 163.367
R1845 B.n607 B.n186 163.367
R1846 B.n607 B.n184 163.367
R1847 B.n611 B.n184 163.367
R1848 B.n611 B.n178 163.367
R1849 B.n620 B.n178 163.367
R1850 B.n620 B.n176 163.367
R1851 B.n624 B.n176 163.367
R1852 B.n624 B.n171 163.367
R1853 B.n632 B.n171 163.367
R1854 B.n632 B.n169 163.367
R1855 B.n636 B.n169 163.367
R1856 B.n636 B.n163 163.367
R1857 B.n644 B.n163 163.367
R1858 B.n644 B.n161 163.367
R1859 B.n648 B.n161 163.367
R1860 B.n648 B.n155 163.367
R1861 B.n657 B.n155 163.367
R1862 B.n657 B.n153 163.367
R1863 B.n661 B.n153 163.367
R1864 B.n661 B.n2 163.367
R1865 B.n1041 B.n2 163.367
R1866 B.n1041 B.n3 163.367
R1867 B.n1037 B.n3 163.367
R1868 B.n1037 B.n9 163.367
R1869 B.n1033 B.n9 163.367
R1870 B.n1033 B.n11 163.367
R1871 B.n1029 B.n11 163.367
R1872 B.n1029 B.n16 163.367
R1873 B.n1025 B.n16 163.367
R1874 B.n1025 B.n18 163.367
R1875 B.n1021 B.n18 163.367
R1876 B.n1021 B.n23 163.367
R1877 B.n1017 B.n23 163.367
R1878 B.n1017 B.n25 163.367
R1879 B.n1013 B.n25 163.367
R1880 B.n1013 B.n29 163.367
R1881 B.n1009 B.n29 163.367
R1882 B.n1009 B.n31 163.367
R1883 B.n1005 B.n31 163.367
R1884 B.n1005 B.n37 163.367
R1885 B.n1001 B.n37 163.367
R1886 B.n1001 B.n39 163.367
R1887 B.n997 B.n39 163.367
R1888 B.n997 B.n43 163.367
R1889 B.n993 B.n43 163.367
R1890 B.n993 B.n45 163.367
R1891 B.n989 B.n45 163.367
R1892 B.n989 B.n51 163.367
R1893 B.n985 B.n51 163.367
R1894 B.n985 B.n53 163.367
R1895 B.n981 B.n53 163.367
R1896 B.n981 B.n57 163.367
R1897 B.n977 B.n57 163.367
R1898 B.n977 B.n59 163.367
R1899 B.n973 B.n59 163.367
R1900 B.n973 B.n65 163.367
R1901 B.n969 B.n65 163.367
R1902 B.n969 B.n67 163.367
R1903 B.n965 B.n67 163.367
R1904 B.n965 B.n72 163.367
R1905 B.n961 B.n72 163.367
R1906 B.n961 B.n74 163.367
R1907 B.n957 B.n74 163.367
R1908 B.n957 B.n78 163.367
R1909 B.n953 B.n78 163.367
R1910 B.n953 B.n80 163.367
R1911 B.n949 B.n80 163.367
R1912 B.n949 B.n86 163.367
R1913 B.n945 B.n86 163.367
R1914 B.n945 B.n88 163.367
R1915 B.n941 B.n88 163.367
R1916 B.n508 B.n506 163.367
R1917 B.n506 B.n505 163.367
R1918 B.n502 B.n501 163.367
R1919 B.n499 B.n249 163.367
R1920 B.n495 B.n493 163.367
R1921 B.n491 B.n251 163.367
R1922 B.n487 B.n485 163.367
R1923 B.n483 B.n253 163.367
R1924 B.n479 B.n477 163.367
R1925 B.n475 B.n255 163.367
R1926 B.n471 B.n469 163.367
R1927 B.n467 B.n257 163.367
R1928 B.n463 B.n461 163.367
R1929 B.n459 B.n259 163.367
R1930 B.n455 B.n453 163.367
R1931 B.n451 B.n261 163.367
R1932 B.n447 B.n445 163.367
R1933 B.n443 B.n263 163.367
R1934 B.n439 B.n437 163.367
R1935 B.n435 B.n265 163.367
R1936 B.n431 B.n429 163.367
R1937 B.n427 B.n267 163.367
R1938 B.n423 B.n421 163.367
R1939 B.n419 B.n269 163.367
R1940 B.n414 B.n412 163.367
R1941 B.n410 B.n273 163.367
R1942 B.n406 B.n404 163.367
R1943 B.n402 B.n275 163.367
R1944 B.n398 B.n396 163.367
R1945 B.n393 B.n392 163.367
R1946 B.n390 B.n281 163.367
R1947 B.n386 B.n384 163.367
R1948 B.n382 B.n283 163.367
R1949 B.n378 B.n376 163.367
R1950 B.n374 B.n285 163.367
R1951 B.n370 B.n368 163.367
R1952 B.n366 B.n287 163.367
R1953 B.n362 B.n360 163.367
R1954 B.n358 B.n289 163.367
R1955 B.n354 B.n352 163.367
R1956 B.n350 B.n291 163.367
R1957 B.n346 B.n344 163.367
R1958 B.n342 B.n293 163.367
R1959 B.n338 B.n336 163.367
R1960 B.n334 B.n295 163.367
R1961 B.n330 B.n328 163.367
R1962 B.n326 B.n297 163.367
R1963 B.n322 B.n320 163.367
R1964 B.n318 B.n299 163.367
R1965 B.n314 B.n312 163.367
R1966 B.n310 B.n301 163.367
R1967 B.n306 B.n304 163.367
R1968 B.n514 B.n241 163.367
R1969 B.n518 B.n241 163.367
R1970 B.n518 B.n235 163.367
R1971 B.n526 B.n235 163.367
R1972 B.n526 B.n233 163.367
R1973 B.n530 B.n233 163.367
R1974 B.n530 B.n228 163.367
R1975 B.n539 B.n228 163.367
R1976 B.n539 B.n226 163.367
R1977 B.n543 B.n226 163.367
R1978 B.n543 B.n220 163.367
R1979 B.n551 B.n220 163.367
R1980 B.n551 B.n218 163.367
R1981 B.n555 B.n218 163.367
R1982 B.n555 B.n212 163.367
R1983 B.n563 B.n212 163.367
R1984 B.n563 B.n210 163.367
R1985 B.n567 B.n210 163.367
R1986 B.n567 B.n205 163.367
R1987 B.n576 B.n205 163.367
R1988 B.n576 B.n203 163.367
R1989 B.n580 B.n203 163.367
R1990 B.n580 B.n197 163.367
R1991 B.n588 B.n197 163.367
R1992 B.n588 B.n195 163.367
R1993 B.n592 B.n195 163.367
R1994 B.n592 B.n190 163.367
R1995 B.n601 B.n190 163.367
R1996 B.n601 B.n188 163.367
R1997 B.n605 B.n188 163.367
R1998 B.n605 B.n182 163.367
R1999 B.n613 B.n182 163.367
R2000 B.n613 B.n180 163.367
R2001 B.n617 B.n180 163.367
R2002 B.n617 B.n175 163.367
R2003 B.n626 B.n175 163.367
R2004 B.n626 B.n173 163.367
R2005 B.n630 B.n173 163.367
R2006 B.n630 B.n167 163.367
R2007 B.n638 B.n167 163.367
R2008 B.n638 B.n165 163.367
R2009 B.n642 B.n165 163.367
R2010 B.n642 B.n159 163.367
R2011 B.n650 B.n159 163.367
R2012 B.n650 B.n157 163.367
R2013 B.n655 B.n157 163.367
R2014 B.n655 B.n151 163.367
R2015 B.n663 B.n151 163.367
R2016 B.n664 B.n663 163.367
R2017 B.n664 B.n5 163.367
R2018 B.n6 B.n5 163.367
R2019 B.n7 B.n6 163.367
R2020 B.n669 B.n7 163.367
R2021 B.n669 B.n12 163.367
R2022 B.n13 B.n12 163.367
R2023 B.n14 B.n13 163.367
R2024 B.n674 B.n14 163.367
R2025 B.n674 B.n19 163.367
R2026 B.n20 B.n19 163.367
R2027 B.n21 B.n20 163.367
R2028 B.n679 B.n21 163.367
R2029 B.n679 B.n26 163.367
R2030 B.n27 B.n26 163.367
R2031 B.n28 B.n27 163.367
R2032 B.n684 B.n28 163.367
R2033 B.n684 B.n33 163.367
R2034 B.n34 B.n33 163.367
R2035 B.n35 B.n34 163.367
R2036 B.n689 B.n35 163.367
R2037 B.n689 B.n40 163.367
R2038 B.n41 B.n40 163.367
R2039 B.n42 B.n41 163.367
R2040 B.n694 B.n42 163.367
R2041 B.n694 B.n47 163.367
R2042 B.n48 B.n47 163.367
R2043 B.n49 B.n48 163.367
R2044 B.n699 B.n49 163.367
R2045 B.n699 B.n54 163.367
R2046 B.n55 B.n54 163.367
R2047 B.n56 B.n55 163.367
R2048 B.n704 B.n56 163.367
R2049 B.n704 B.n61 163.367
R2050 B.n62 B.n61 163.367
R2051 B.n63 B.n62 163.367
R2052 B.n709 B.n63 163.367
R2053 B.n709 B.n68 163.367
R2054 B.n69 B.n68 163.367
R2055 B.n70 B.n69 163.367
R2056 B.n714 B.n70 163.367
R2057 B.n714 B.n75 163.367
R2058 B.n76 B.n75 163.367
R2059 B.n77 B.n76 163.367
R2060 B.n719 B.n77 163.367
R2061 B.n719 B.n82 163.367
R2062 B.n83 B.n82 163.367
R2063 B.n84 B.n83 163.367
R2064 B.n724 B.n84 163.367
R2065 B.n724 B.n89 163.367
R2066 B.n90 B.n89 163.367
R2067 B.n91 B.n90 163.367
R2068 B.n937 B.n935 163.367
R2069 B.n933 B.n95 163.367
R2070 B.n929 B.n927 163.367
R2071 B.n925 B.n97 163.367
R2072 B.n921 B.n919 163.367
R2073 B.n917 B.n99 163.367
R2074 B.n913 B.n911 163.367
R2075 B.n909 B.n101 163.367
R2076 B.n905 B.n903 163.367
R2077 B.n901 B.n103 163.367
R2078 B.n897 B.n895 163.367
R2079 B.n893 B.n105 163.367
R2080 B.n889 B.n887 163.367
R2081 B.n885 B.n107 163.367
R2082 B.n881 B.n879 163.367
R2083 B.n877 B.n109 163.367
R2084 B.n873 B.n871 163.367
R2085 B.n869 B.n111 163.367
R2086 B.n865 B.n863 163.367
R2087 B.n861 B.n113 163.367
R2088 B.n857 B.n855 163.367
R2089 B.n853 B.n115 163.367
R2090 B.n849 B.n847 163.367
R2091 B.n845 B.n117 163.367
R2092 B.n840 B.n838 163.367
R2093 B.n836 B.n121 163.367
R2094 B.n832 B.n830 163.367
R2095 B.n828 B.n123 163.367
R2096 B.n823 B.n821 163.367
R2097 B.n819 B.n127 163.367
R2098 B.n815 B.n813 163.367
R2099 B.n811 B.n129 163.367
R2100 B.n807 B.n805 163.367
R2101 B.n803 B.n131 163.367
R2102 B.n799 B.n797 163.367
R2103 B.n795 B.n133 163.367
R2104 B.n791 B.n789 163.367
R2105 B.n787 B.n135 163.367
R2106 B.n783 B.n781 163.367
R2107 B.n779 B.n137 163.367
R2108 B.n775 B.n773 163.367
R2109 B.n771 B.n139 163.367
R2110 B.n767 B.n765 163.367
R2111 B.n763 B.n141 163.367
R2112 B.n759 B.n757 163.367
R2113 B.n755 B.n143 163.367
R2114 B.n751 B.n749 163.367
R2115 B.n747 B.n145 163.367
R2116 B.n743 B.n741 163.367
R2117 B.n739 B.n147 163.367
R2118 B.n735 B.n733 163.367
R2119 B.n731 B.n149 163.367
R2120 B.n507 B.n245 71.676
R2121 B.n505 B.n247 71.676
R2122 B.n501 B.n500 71.676
R2123 B.n494 B.n249 71.676
R2124 B.n493 B.n492 71.676
R2125 B.n486 B.n251 71.676
R2126 B.n485 B.n484 71.676
R2127 B.n478 B.n253 71.676
R2128 B.n477 B.n476 71.676
R2129 B.n470 B.n255 71.676
R2130 B.n469 B.n468 71.676
R2131 B.n462 B.n257 71.676
R2132 B.n461 B.n460 71.676
R2133 B.n454 B.n259 71.676
R2134 B.n453 B.n452 71.676
R2135 B.n446 B.n261 71.676
R2136 B.n445 B.n444 71.676
R2137 B.n438 B.n263 71.676
R2138 B.n437 B.n436 71.676
R2139 B.n430 B.n265 71.676
R2140 B.n429 B.n428 71.676
R2141 B.n422 B.n267 71.676
R2142 B.n421 B.n420 71.676
R2143 B.n413 B.n269 71.676
R2144 B.n412 B.n411 71.676
R2145 B.n405 B.n273 71.676
R2146 B.n404 B.n403 71.676
R2147 B.n397 B.n275 71.676
R2148 B.n396 B.n279 71.676
R2149 B.n392 B.n391 71.676
R2150 B.n385 B.n281 71.676
R2151 B.n384 B.n383 71.676
R2152 B.n377 B.n283 71.676
R2153 B.n376 B.n375 71.676
R2154 B.n369 B.n285 71.676
R2155 B.n368 B.n367 71.676
R2156 B.n361 B.n287 71.676
R2157 B.n360 B.n359 71.676
R2158 B.n353 B.n289 71.676
R2159 B.n352 B.n351 71.676
R2160 B.n345 B.n291 71.676
R2161 B.n344 B.n343 71.676
R2162 B.n337 B.n293 71.676
R2163 B.n336 B.n335 71.676
R2164 B.n329 B.n295 71.676
R2165 B.n328 B.n327 71.676
R2166 B.n321 B.n297 71.676
R2167 B.n320 B.n319 71.676
R2168 B.n313 B.n299 71.676
R2169 B.n312 B.n311 71.676
R2170 B.n305 B.n301 71.676
R2171 B.n304 B.n303 71.676
R2172 B.n936 B.n93 71.676
R2173 B.n935 B.n934 71.676
R2174 B.n928 B.n95 71.676
R2175 B.n927 B.n926 71.676
R2176 B.n920 B.n97 71.676
R2177 B.n919 B.n918 71.676
R2178 B.n912 B.n99 71.676
R2179 B.n911 B.n910 71.676
R2180 B.n904 B.n101 71.676
R2181 B.n903 B.n902 71.676
R2182 B.n896 B.n103 71.676
R2183 B.n895 B.n894 71.676
R2184 B.n888 B.n105 71.676
R2185 B.n887 B.n886 71.676
R2186 B.n880 B.n107 71.676
R2187 B.n879 B.n878 71.676
R2188 B.n872 B.n109 71.676
R2189 B.n871 B.n870 71.676
R2190 B.n864 B.n111 71.676
R2191 B.n863 B.n862 71.676
R2192 B.n856 B.n113 71.676
R2193 B.n855 B.n854 71.676
R2194 B.n848 B.n115 71.676
R2195 B.n847 B.n846 71.676
R2196 B.n839 B.n117 71.676
R2197 B.n838 B.n837 71.676
R2198 B.n831 B.n121 71.676
R2199 B.n830 B.n829 71.676
R2200 B.n822 B.n123 71.676
R2201 B.n821 B.n820 71.676
R2202 B.n814 B.n127 71.676
R2203 B.n813 B.n812 71.676
R2204 B.n806 B.n129 71.676
R2205 B.n805 B.n804 71.676
R2206 B.n798 B.n131 71.676
R2207 B.n797 B.n796 71.676
R2208 B.n790 B.n133 71.676
R2209 B.n789 B.n788 71.676
R2210 B.n782 B.n135 71.676
R2211 B.n781 B.n780 71.676
R2212 B.n774 B.n137 71.676
R2213 B.n773 B.n772 71.676
R2214 B.n766 B.n139 71.676
R2215 B.n765 B.n764 71.676
R2216 B.n758 B.n141 71.676
R2217 B.n757 B.n756 71.676
R2218 B.n750 B.n143 71.676
R2219 B.n749 B.n748 71.676
R2220 B.n742 B.n145 71.676
R2221 B.n741 B.n740 71.676
R2222 B.n734 B.n147 71.676
R2223 B.n733 B.n732 71.676
R2224 B.n732 B.n731 71.676
R2225 B.n735 B.n734 71.676
R2226 B.n740 B.n739 71.676
R2227 B.n743 B.n742 71.676
R2228 B.n748 B.n747 71.676
R2229 B.n751 B.n750 71.676
R2230 B.n756 B.n755 71.676
R2231 B.n759 B.n758 71.676
R2232 B.n764 B.n763 71.676
R2233 B.n767 B.n766 71.676
R2234 B.n772 B.n771 71.676
R2235 B.n775 B.n774 71.676
R2236 B.n780 B.n779 71.676
R2237 B.n783 B.n782 71.676
R2238 B.n788 B.n787 71.676
R2239 B.n791 B.n790 71.676
R2240 B.n796 B.n795 71.676
R2241 B.n799 B.n798 71.676
R2242 B.n804 B.n803 71.676
R2243 B.n807 B.n806 71.676
R2244 B.n812 B.n811 71.676
R2245 B.n815 B.n814 71.676
R2246 B.n820 B.n819 71.676
R2247 B.n823 B.n822 71.676
R2248 B.n829 B.n828 71.676
R2249 B.n832 B.n831 71.676
R2250 B.n837 B.n836 71.676
R2251 B.n840 B.n839 71.676
R2252 B.n846 B.n845 71.676
R2253 B.n849 B.n848 71.676
R2254 B.n854 B.n853 71.676
R2255 B.n857 B.n856 71.676
R2256 B.n862 B.n861 71.676
R2257 B.n865 B.n864 71.676
R2258 B.n870 B.n869 71.676
R2259 B.n873 B.n872 71.676
R2260 B.n878 B.n877 71.676
R2261 B.n881 B.n880 71.676
R2262 B.n886 B.n885 71.676
R2263 B.n889 B.n888 71.676
R2264 B.n894 B.n893 71.676
R2265 B.n897 B.n896 71.676
R2266 B.n902 B.n901 71.676
R2267 B.n905 B.n904 71.676
R2268 B.n910 B.n909 71.676
R2269 B.n913 B.n912 71.676
R2270 B.n918 B.n917 71.676
R2271 B.n921 B.n920 71.676
R2272 B.n926 B.n925 71.676
R2273 B.n929 B.n928 71.676
R2274 B.n934 B.n933 71.676
R2275 B.n937 B.n936 71.676
R2276 B.n508 B.n507 71.676
R2277 B.n502 B.n247 71.676
R2278 B.n500 B.n499 71.676
R2279 B.n495 B.n494 71.676
R2280 B.n492 B.n491 71.676
R2281 B.n487 B.n486 71.676
R2282 B.n484 B.n483 71.676
R2283 B.n479 B.n478 71.676
R2284 B.n476 B.n475 71.676
R2285 B.n471 B.n470 71.676
R2286 B.n468 B.n467 71.676
R2287 B.n463 B.n462 71.676
R2288 B.n460 B.n459 71.676
R2289 B.n455 B.n454 71.676
R2290 B.n452 B.n451 71.676
R2291 B.n447 B.n446 71.676
R2292 B.n444 B.n443 71.676
R2293 B.n439 B.n438 71.676
R2294 B.n436 B.n435 71.676
R2295 B.n431 B.n430 71.676
R2296 B.n428 B.n427 71.676
R2297 B.n423 B.n422 71.676
R2298 B.n420 B.n419 71.676
R2299 B.n414 B.n413 71.676
R2300 B.n411 B.n410 71.676
R2301 B.n406 B.n405 71.676
R2302 B.n403 B.n402 71.676
R2303 B.n398 B.n397 71.676
R2304 B.n393 B.n279 71.676
R2305 B.n391 B.n390 71.676
R2306 B.n386 B.n385 71.676
R2307 B.n383 B.n382 71.676
R2308 B.n378 B.n377 71.676
R2309 B.n375 B.n374 71.676
R2310 B.n370 B.n369 71.676
R2311 B.n367 B.n366 71.676
R2312 B.n362 B.n361 71.676
R2313 B.n359 B.n358 71.676
R2314 B.n354 B.n353 71.676
R2315 B.n351 B.n350 71.676
R2316 B.n346 B.n345 71.676
R2317 B.n343 B.n342 71.676
R2318 B.n338 B.n337 71.676
R2319 B.n335 B.n334 71.676
R2320 B.n330 B.n329 71.676
R2321 B.n327 B.n326 71.676
R2322 B.n322 B.n321 71.676
R2323 B.n319 B.n318 71.676
R2324 B.n314 B.n313 71.676
R2325 B.n311 B.n310 71.676
R2326 B.n306 B.n305 71.676
R2327 B.n303 B.n243 71.676
R2328 B.n513 B.n244 71.0049
R2329 B.n942 B.n92 71.0049
R2330 B.n278 B.n277 59.5399
R2331 B.n416 B.n271 59.5399
R2332 B.n843 B.n119 59.5399
R2333 B.n825 B.n125 59.5399
R2334 B.n277 B.n276 55.2732
R2335 B.n271 B.n270 55.2732
R2336 B.n119 B.n118 55.2732
R2337 B.n125 B.n124 55.2732
R2338 B.n513 B.n240 38.6269
R2339 B.n519 B.n240 38.6269
R2340 B.n519 B.n236 38.6269
R2341 B.n525 B.n236 38.6269
R2342 B.n525 B.n232 38.6269
R2343 B.n532 B.n232 38.6269
R2344 B.n532 B.n531 38.6269
R2345 B.n538 B.n225 38.6269
R2346 B.n544 B.n225 38.6269
R2347 B.n544 B.n221 38.6269
R2348 B.n550 B.n221 38.6269
R2349 B.n550 B.n217 38.6269
R2350 B.n556 B.n217 38.6269
R2351 B.n556 B.n213 38.6269
R2352 B.n562 B.n213 38.6269
R2353 B.n562 B.n209 38.6269
R2354 B.n569 B.n209 38.6269
R2355 B.n569 B.n568 38.6269
R2356 B.n575 B.n202 38.6269
R2357 B.n581 B.n202 38.6269
R2358 B.n581 B.n198 38.6269
R2359 B.n587 B.n198 38.6269
R2360 B.n587 B.n194 38.6269
R2361 B.n594 B.n194 38.6269
R2362 B.n594 B.n593 38.6269
R2363 B.n600 B.n187 38.6269
R2364 B.n606 B.n187 38.6269
R2365 B.n606 B.n183 38.6269
R2366 B.n612 B.n183 38.6269
R2367 B.n612 B.n179 38.6269
R2368 B.n619 B.n179 38.6269
R2369 B.n619 B.n618 38.6269
R2370 B.n625 B.n172 38.6269
R2371 B.n631 B.n172 38.6269
R2372 B.n631 B.n168 38.6269
R2373 B.n637 B.n168 38.6269
R2374 B.n637 B.n164 38.6269
R2375 B.n643 B.n164 38.6269
R2376 B.n643 B.n160 38.6269
R2377 B.n649 B.n160 38.6269
R2378 B.n656 B.n156 38.6269
R2379 B.n656 B.n152 38.6269
R2380 B.n662 B.n152 38.6269
R2381 B.n662 B.n4 38.6269
R2382 B.n1040 B.n4 38.6269
R2383 B.n1040 B.n1039 38.6269
R2384 B.n1039 B.n1038 38.6269
R2385 B.n1038 B.n8 38.6269
R2386 B.n1032 B.n8 38.6269
R2387 B.n1032 B.n1031 38.6269
R2388 B.n1030 B.n15 38.6269
R2389 B.n1024 B.n15 38.6269
R2390 B.n1024 B.n1023 38.6269
R2391 B.n1023 B.n1022 38.6269
R2392 B.n1022 B.n22 38.6269
R2393 B.n1016 B.n22 38.6269
R2394 B.n1016 B.n1015 38.6269
R2395 B.n1015 B.n1014 38.6269
R2396 B.n1008 B.n32 38.6269
R2397 B.n1008 B.n1007 38.6269
R2398 B.n1007 B.n1006 38.6269
R2399 B.n1006 B.n36 38.6269
R2400 B.n1000 B.n36 38.6269
R2401 B.n1000 B.n999 38.6269
R2402 B.n999 B.n998 38.6269
R2403 B.n992 B.n46 38.6269
R2404 B.n992 B.n991 38.6269
R2405 B.n991 B.n990 38.6269
R2406 B.n990 B.n50 38.6269
R2407 B.n984 B.n50 38.6269
R2408 B.n984 B.n983 38.6269
R2409 B.n983 B.n982 38.6269
R2410 B.n976 B.n60 38.6269
R2411 B.n976 B.n975 38.6269
R2412 B.n975 B.n974 38.6269
R2413 B.n974 B.n64 38.6269
R2414 B.n968 B.n64 38.6269
R2415 B.n968 B.n967 38.6269
R2416 B.n967 B.n966 38.6269
R2417 B.n966 B.n71 38.6269
R2418 B.n960 B.n71 38.6269
R2419 B.n960 B.n959 38.6269
R2420 B.n959 B.n958 38.6269
R2421 B.n952 B.n81 38.6269
R2422 B.n952 B.n951 38.6269
R2423 B.n951 B.n950 38.6269
R2424 B.n950 B.n85 38.6269
R2425 B.n944 B.n85 38.6269
R2426 B.n944 B.n943 38.6269
R2427 B.n943 B.n942 38.6269
R2428 B.n575 B.t7 36.3547
R2429 B.n982 B.t2 36.3547
R2430 B.n940 B.n939 33.2493
R2431 B.n729 B.n728 33.2493
R2432 B.n515 B.n242 33.2493
R2433 B.n511 B.n510 33.2493
R2434 B.n618 B.t3 31.8105
R2435 B.n32 B.t6 31.8105
R2436 B.t4 B.n156 30.6744
R2437 B.n1031 B.t0 30.6744
R2438 B.n600 B.t5 21.5858
R2439 B.n998 B.t1 21.5858
R2440 B.n538 B.t13 20.4498
R2441 B.n958 B.t9 20.4498
R2442 B.n531 B.t13 18.1776
R2443 B.n81 B.t9 18.1776
R2444 B B.n1042 18.0485
R2445 B.n593 B.t5 17.0416
R2446 B.n46 B.t1 17.0416
R2447 B.n939 B.n938 10.6151
R2448 B.n938 B.n94 10.6151
R2449 B.n932 B.n94 10.6151
R2450 B.n932 B.n931 10.6151
R2451 B.n931 B.n930 10.6151
R2452 B.n930 B.n96 10.6151
R2453 B.n924 B.n96 10.6151
R2454 B.n924 B.n923 10.6151
R2455 B.n923 B.n922 10.6151
R2456 B.n922 B.n98 10.6151
R2457 B.n916 B.n98 10.6151
R2458 B.n916 B.n915 10.6151
R2459 B.n915 B.n914 10.6151
R2460 B.n914 B.n100 10.6151
R2461 B.n908 B.n100 10.6151
R2462 B.n908 B.n907 10.6151
R2463 B.n907 B.n906 10.6151
R2464 B.n906 B.n102 10.6151
R2465 B.n900 B.n102 10.6151
R2466 B.n900 B.n899 10.6151
R2467 B.n899 B.n898 10.6151
R2468 B.n898 B.n104 10.6151
R2469 B.n892 B.n104 10.6151
R2470 B.n892 B.n891 10.6151
R2471 B.n891 B.n890 10.6151
R2472 B.n890 B.n106 10.6151
R2473 B.n884 B.n106 10.6151
R2474 B.n884 B.n883 10.6151
R2475 B.n883 B.n882 10.6151
R2476 B.n882 B.n108 10.6151
R2477 B.n876 B.n108 10.6151
R2478 B.n876 B.n875 10.6151
R2479 B.n875 B.n874 10.6151
R2480 B.n874 B.n110 10.6151
R2481 B.n868 B.n110 10.6151
R2482 B.n868 B.n867 10.6151
R2483 B.n867 B.n866 10.6151
R2484 B.n866 B.n112 10.6151
R2485 B.n860 B.n112 10.6151
R2486 B.n860 B.n859 10.6151
R2487 B.n859 B.n858 10.6151
R2488 B.n858 B.n114 10.6151
R2489 B.n852 B.n114 10.6151
R2490 B.n852 B.n851 10.6151
R2491 B.n851 B.n850 10.6151
R2492 B.n850 B.n116 10.6151
R2493 B.n844 B.n116 10.6151
R2494 B.n842 B.n841 10.6151
R2495 B.n841 B.n120 10.6151
R2496 B.n835 B.n120 10.6151
R2497 B.n835 B.n834 10.6151
R2498 B.n834 B.n833 10.6151
R2499 B.n833 B.n122 10.6151
R2500 B.n827 B.n122 10.6151
R2501 B.n827 B.n826 10.6151
R2502 B.n824 B.n126 10.6151
R2503 B.n818 B.n126 10.6151
R2504 B.n818 B.n817 10.6151
R2505 B.n817 B.n816 10.6151
R2506 B.n816 B.n128 10.6151
R2507 B.n810 B.n128 10.6151
R2508 B.n810 B.n809 10.6151
R2509 B.n809 B.n808 10.6151
R2510 B.n808 B.n130 10.6151
R2511 B.n802 B.n130 10.6151
R2512 B.n802 B.n801 10.6151
R2513 B.n801 B.n800 10.6151
R2514 B.n800 B.n132 10.6151
R2515 B.n794 B.n132 10.6151
R2516 B.n794 B.n793 10.6151
R2517 B.n793 B.n792 10.6151
R2518 B.n792 B.n134 10.6151
R2519 B.n786 B.n134 10.6151
R2520 B.n786 B.n785 10.6151
R2521 B.n785 B.n784 10.6151
R2522 B.n784 B.n136 10.6151
R2523 B.n778 B.n136 10.6151
R2524 B.n778 B.n777 10.6151
R2525 B.n777 B.n776 10.6151
R2526 B.n776 B.n138 10.6151
R2527 B.n770 B.n138 10.6151
R2528 B.n770 B.n769 10.6151
R2529 B.n769 B.n768 10.6151
R2530 B.n768 B.n140 10.6151
R2531 B.n762 B.n140 10.6151
R2532 B.n762 B.n761 10.6151
R2533 B.n761 B.n760 10.6151
R2534 B.n760 B.n142 10.6151
R2535 B.n754 B.n142 10.6151
R2536 B.n754 B.n753 10.6151
R2537 B.n753 B.n752 10.6151
R2538 B.n752 B.n144 10.6151
R2539 B.n746 B.n144 10.6151
R2540 B.n746 B.n745 10.6151
R2541 B.n745 B.n744 10.6151
R2542 B.n744 B.n146 10.6151
R2543 B.n738 B.n146 10.6151
R2544 B.n738 B.n737 10.6151
R2545 B.n737 B.n736 10.6151
R2546 B.n736 B.n148 10.6151
R2547 B.n730 B.n148 10.6151
R2548 B.n730 B.n729 10.6151
R2549 B.n516 B.n515 10.6151
R2550 B.n517 B.n516 10.6151
R2551 B.n517 B.n234 10.6151
R2552 B.n527 B.n234 10.6151
R2553 B.n528 B.n527 10.6151
R2554 B.n529 B.n528 10.6151
R2555 B.n529 B.n227 10.6151
R2556 B.n540 B.n227 10.6151
R2557 B.n541 B.n540 10.6151
R2558 B.n542 B.n541 10.6151
R2559 B.n542 B.n219 10.6151
R2560 B.n552 B.n219 10.6151
R2561 B.n553 B.n552 10.6151
R2562 B.n554 B.n553 10.6151
R2563 B.n554 B.n211 10.6151
R2564 B.n564 B.n211 10.6151
R2565 B.n565 B.n564 10.6151
R2566 B.n566 B.n565 10.6151
R2567 B.n566 B.n204 10.6151
R2568 B.n577 B.n204 10.6151
R2569 B.n578 B.n577 10.6151
R2570 B.n579 B.n578 10.6151
R2571 B.n579 B.n196 10.6151
R2572 B.n589 B.n196 10.6151
R2573 B.n590 B.n589 10.6151
R2574 B.n591 B.n590 10.6151
R2575 B.n591 B.n189 10.6151
R2576 B.n602 B.n189 10.6151
R2577 B.n603 B.n602 10.6151
R2578 B.n604 B.n603 10.6151
R2579 B.n604 B.n181 10.6151
R2580 B.n614 B.n181 10.6151
R2581 B.n615 B.n614 10.6151
R2582 B.n616 B.n615 10.6151
R2583 B.n616 B.n174 10.6151
R2584 B.n627 B.n174 10.6151
R2585 B.n628 B.n627 10.6151
R2586 B.n629 B.n628 10.6151
R2587 B.n629 B.n166 10.6151
R2588 B.n639 B.n166 10.6151
R2589 B.n640 B.n639 10.6151
R2590 B.n641 B.n640 10.6151
R2591 B.n641 B.n158 10.6151
R2592 B.n651 B.n158 10.6151
R2593 B.n652 B.n651 10.6151
R2594 B.n654 B.n652 10.6151
R2595 B.n654 B.n653 10.6151
R2596 B.n653 B.n150 10.6151
R2597 B.n665 B.n150 10.6151
R2598 B.n666 B.n665 10.6151
R2599 B.n667 B.n666 10.6151
R2600 B.n668 B.n667 10.6151
R2601 B.n670 B.n668 10.6151
R2602 B.n671 B.n670 10.6151
R2603 B.n672 B.n671 10.6151
R2604 B.n673 B.n672 10.6151
R2605 B.n675 B.n673 10.6151
R2606 B.n676 B.n675 10.6151
R2607 B.n677 B.n676 10.6151
R2608 B.n678 B.n677 10.6151
R2609 B.n680 B.n678 10.6151
R2610 B.n681 B.n680 10.6151
R2611 B.n682 B.n681 10.6151
R2612 B.n683 B.n682 10.6151
R2613 B.n685 B.n683 10.6151
R2614 B.n686 B.n685 10.6151
R2615 B.n687 B.n686 10.6151
R2616 B.n688 B.n687 10.6151
R2617 B.n690 B.n688 10.6151
R2618 B.n691 B.n690 10.6151
R2619 B.n692 B.n691 10.6151
R2620 B.n693 B.n692 10.6151
R2621 B.n695 B.n693 10.6151
R2622 B.n696 B.n695 10.6151
R2623 B.n697 B.n696 10.6151
R2624 B.n698 B.n697 10.6151
R2625 B.n700 B.n698 10.6151
R2626 B.n701 B.n700 10.6151
R2627 B.n702 B.n701 10.6151
R2628 B.n703 B.n702 10.6151
R2629 B.n705 B.n703 10.6151
R2630 B.n706 B.n705 10.6151
R2631 B.n707 B.n706 10.6151
R2632 B.n708 B.n707 10.6151
R2633 B.n710 B.n708 10.6151
R2634 B.n711 B.n710 10.6151
R2635 B.n712 B.n711 10.6151
R2636 B.n713 B.n712 10.6151
R2637 B.n715 B.n713 10.6151
R2638 B.n716 B.n715 10.6151
R2639 B.n717 B.n716 10.6151
R2640 B.n718 B.n717 10.6151
R2641 B.n720 B.n718 10.6151
R2642 B.n721 B.n720 10.6151
R2643 B.n722 B.n721 10.6151
R2644 B.n723 B.n722 10.6151
R2645 B.n725 B.n723 10.6151
R2646 B.n726 B.n725 10.6151
R2647 B.n727 B.n726 10.6151
R2648 B.n728 B.n727 10.6151
R2649 B.n510 B.n509 10.6151
R2650 B.n509 B.n246 10.6151
R2651 B.n504 B.n246 10.6151
R2652 B.n504 B.n503 10.6151
R2653 B.n503 B.n248 10.6151
R2654 B.n498 B.n248 10.6151
R2655 B.n498 B.n497 10.6151
R2656 B.n497 B.n496 10.6151
R2657 B.n496 B.n250 10.6151
R2658 B.n490 B.n250 10.6151
R2659 B.n490 B.n489 10.6151
R2660 B.n489 B.n488 10.6151
R2661 B.n488 B.n252 10.6151
R2662 B.n482 B.n252 10.6151
R2663 B.n482 B.n481 10.6151
R2664 B.n481 B.n480 10.6151
R2665 B.n480 B.n254 10.6151
R2666 B.n474 B.n254 10.6151
R2667 B.n474 B.n473 10.6151
R2668 B.n473 B.n472 10.6151
R2669 B.n472 B.n256 10.6151
R2670 B.n466 B.n256 10.6151
R2671 B.n466 B.n465 10.6151
R2672 B.n465 B.n464 10.6151
R2673 B.n464 B.n258 10.6151
R2674 B.n458 B.n258 10.6151
R2675 B.n458 B.n457 10.6151
R2676 B.n457 B.n456 10.6151
R2677 B.n456 B.n260 10.6151
R2678 B.n450 B.n260 10.6151
R2679 B.n450 B.n449 10.6151
R2680 B.n449 B.n448 10.6151
R2681 B.n448 B.n262 10.6151
R2682 B.n442 B.n262 10.6151
R2683 B.n442 B.n441 10.6151
R2684 B.n441 B.n440 10.6151
R2685 B.n440 B.n264 10.6151
R2686 B.n434 B.n264 10.6151
R2687 B.n434 B.n433 10.6151
R2688 B.n433 B.n432 10.6151
R2689 B.n432 B.n266 10.6151
R2690 B.n426 B.n266 10.6151
R2691 B.n426 B.n425 10.6151
R2692 B.n425 B.n424 10.6151
R2693 B.n424 B.n268 10.6151
R2694 B.n418 B.n268 10.6151
R2695 B.n418 B.n417 10.6151
R2696 B.n415 B.n272 10.6151
R2697 B.n409 B.n272 10.6151
R2698 B.n409 B.n408 10.6151
R2699 B.n408 B.n407 10.6151
R2700 B.n407 B.n274 10.6151
R2701 B.n401 B.n274 10.6151
R2702 B.n401 B.n400 10.6151
R2703 B.n400 B.n399 10.6151
R2704 B.n395 B.n394 10.6151
R2705 B.n394 B.n280 10.6151
R2706 B.n389 B.n280 10.6151
R2707 B.n389 B.n388 10.6151
R2708 B.n388 B.n387 10.6151
R2709 B.n387 B.n282 10.6151
R2710 B.n381 B.n282 10.6151
R2711 B.n381 B.n380 10.6151
R2712 B.n380 B.n379 10.6151
R2713 B.n379 B.n284 10.6151
R2714 B.n373 B.n284 10.6151
R2715 B.n373 B.n372 10.6151
R2716 B.n372 B.n371 10.6151
R2717 B.n371 B.n286 10.6151
R2718 B.n365 B.n286 10.6151
R2719 B.n365 B.n364 10.6151
R2720 B.n364 B.n363 10.6151
R2721 B.n363 B.n288 10.6151
R2722 B.n357 B.n288 10.6151
R2723 B.n357 B.n356 10.6151
R2724 B.n356 B.n355 10.6151
R2725 B.n355 B.n290 10.6151
R2726 B.n349 B.n290 10.6151
R2727 B.n349 B.n348 10.6151
R2728 B.n348 B.n347 10.6151
R2729 B.n347 B.n292 10.6151
R2730 B.n341 B.n292 10.6151
R2731 B.n341 B.n340 10.6151
R2732 B.n340 B.n339 10.6151
R2733 B.n339 B.n294 10.6151
R2734 B.n333 B.n294 10.6151
R2735 B.n333 B.n332 10.6151
R2736 B.n332 B.n331 10.6151
R2737 B.n331 B.n296 10.6151
R2738 B.n325 B.n296 10.6151
R2739 B.n325 B.n324 10.6151
R2740 B.n324 B.n323 10.6151
R2741 B.n323 B.n298 10.6151
R2742 B.n317 B.n298 10.6151
R2743 B.n317 B.n316 10.6151
R2744 B.n316 B.n315 10.6151
R2745 B.n315 B.n300 10.6151
R2746 B.n309 B.n300 10.6151
R2747 B.n309 B.n308 10.6151
R2748 B.n308 B.n307 10.6151
R2749 B.n307 B.n302 10.6151
R2750 B.n302 B.n242 10.6151
R2751 B.n511 B.n238 10.6151
R2752 B.n521 B.n238 10.6151
R2753 B.n522 B.n521 10.6151
R2754 B.n523 B.n522 10.6151
R2755 B.n523 B.n230 10.6151
R2756 B.n534 B.n230 10.6151
R2757 B.n535 B.n534 10.6151
R2758 B.n536 B.n535 10.6151
R2759 B.n536 B.n223 10.6151
R2760 B.n546 B.n223 10.6151
R2761 B.n547 B.n546 10.6151
R2762 B.n548 B.n547 10.6151
R2763 B.n548 B.n215 10.6151
R2764 B.n558 B.n215 10.6151
R2765 B.n559 B.n558 10.6151
R2766 B.n560 B.n559 10.6151
R2767 B.n560 B.n207 10.6151
R2768 B.n571 B.n207 10.6151
R2769 B.n572 B.n571 10.6151
R2770 B.n573 B.n572 10.6151
R2771 B.n573 B.n200 10.6151
R2772 B.n583 B.n200 10.6151
R2773 B.n584 B.n583 10.6151
R2774 B.n585 B.n584 10.6151
R2775 B.n585 B.n192 10.6151
R2776 B.n596 B.n192 10.6151
R2777 B.n597 B.n596 10.6151
R2778 B.n598 B.n597 10.6151
R2779 B.n598 B.n185 10.6151
R2780 B.n608 B.n185 10.6151
R2781 B.n609 B.n608 10.6151
R2782 B.n610 B.n609 10.6151
R2783 B.n610 B.n177 10.6151
R2784 B.n621 B.n177 10.6151
R2785 B.n622 B.n621 10.6151
R2786 B.n623 B.n622 10.6151
R2787 B.n623 B.n170 10.6151
R2788 B.n633 B.n170 10.6151
R2789 B.n634 B.n633 10.6151
R2790 B.n635 B.n634 10.6151
R2791 B.n635 B.n162 10.6151
R2792 B.n645 B.n162 10.6151
R2793 B.n646 B.n645 10.6151
R2794 B.n647 B.n646 10.6151
R2795 B.n647 B.n154 10.6151
R2796 B.n658 B.n154 10.6151
R2797 B.n659 B.n658 10.6151
R2798 B.n660 B.n659 10.6151
R2799 B.n660 B.n0 10.6151
R2800 B.n1036 B.n1 10.6151
R2801 B.n1036 B.n1035 10.6151
R2802 B.n1035 B.n1034 10.6151
R2803 B.n1034 B.n10 10.6151
R2804 B.n1028 B.n10 10.6151
R2805 B.n1028 B.n1027 10.6151
R2806 B.n1027 B.n1026 10.6151
R2807 B.n1026 B.n17 10.6151
R2808 B.n1020 B.n17 10.6151
R2809 B.n1020 B.n1019 10.6151
R2810 B.n1019 B.n1018 10.6151
R2811 B.n1018 B.n24 10.6151
R2812 B.n1012 B.n24 10.6151
R2813 B.n1012 B.n1011 10.6151
R2814 B.n1011 B.n1010 10.6151
R2815 B.n1010 B.n30 10.6151
R2816 B.n1004 B.n30 10.6151
R2817 B.n1004 B.n1003 10.6151
R2818 B.n1003 B.n1002 10.6151
R2819 B.n1002 B.n38 10.6151
R2820 B.n996 B.n38 10.6151
R2821 B.n996 B.n995 10.6151
R2822 B.n995 B.n994 10.6151
R2823 B.n994 B.n44 10.6151
R2824 B.n988 B.n44 10.6151
R2825 B.n988 B.n987 10.6151
R2826 B.n987 B.n986 10.6151
R2827 B.n986 B.n52 10.6151
R2828 B.n980 B.n52 10.6151
R2829 B.n980 B.n979 10.6151
R2830 B.n979 B.n978 10.6151
R2831 B.n978 B.n58 10.6151
R2832 B.n972 B.n58 10.6151
R2833 B.n972 B.n971 10.6151
R2834 B.n971 B.n970 10.6151
R2835 B.n970 B.n66 10.6151
R2836 B.n964 B.n66 10.6151
R2837 B.n964 B.n963 10.6151
R2838 B.n963 B.n962 10.6151
R2839 B.n962 B.n73 10.6151
R2840 B.n956 B.n73 10.6151
R2841 B.n956 B.n955 10.6151
R2842 B.n955 B.n954 10.6151
R2843 B.n954 B.n79 10.6151
R2844 B.n948 B.n79 10.6151
R2845 B.n948 B.n947 10.6151
R2846 B.n947 B.n946 10.6151
R2847 B.n946 B.n87 10.6151
R2848 B.n940 B.n87 10.6151
R2849 B.n649 B.t4 7.95299
R2850 B.t0 B.n1030 7.95299
R2851 B.n625 B.t3 6.81692
R2852 B.n1014 B.t6 6.81692
R2853 B.n843 B.n842 6.5566
R2854 B.n826 B.n825 6.5566
R2855 B.n416 B.n415 6.5566
R2856 B.n399 B.n278 6.5566
R2857 B.n844 B.n843 4.05904
R2858 B.n825 B.n824 4.05904
R2859 B.n417 B.n416 4.05904
R2860 B.n395 B.n278 4.05904
R2861 B.n1042 B.n0 2.81026
R2862 B.n1042 B.n1 2.81026
R2863 B.n568 B.t7 2.27264
R2864 B.n60 B.t2 2.27264
R2865 VN.n6 VN.t5 169.323
R2866 VN.n33 VN.t3 169.323
R2867 VN.n51 VN.n27 161.3
R2868 VN.n50 VN.n49 161.3
R2869 VN.n48 VN.n28 161.3
R2870 VN.n47 VN.n46 161.3
R2871 VN.n45 VN.n29 161.3
R2872 VN.n44 VN.n43 161.3
R2873 VN.n42 VN.n41 161.3
R2874 VN.n40 VN.n31 161.3
R2875 VN.n39 VN.n38 161.3
R2876 VN.n37 VN.n32 161.3
R2877 VN.n36 VN.n35 161.3
R2878 VN.n24 VN.n0 161.3
R2879 VN.n23 VN.n22 161.3
R2880 VN.n21 VN.n1 161.3
R2881 VN.n20 VN.n19 161.3
R2882 VN.n18 VN.n2 161.3
R2883 VN.n17 VN.n16 161.3
R2884 VN.n15 VN.n14 161.3
R2885 VN.n13 VN.n4 161.3
R2886 VN.n12 VN.n11 161.3
R2887 VN.n10 VN.n5 161.3
R2888 VN.n9 VN.n8 161.3
R2889 VN.n7 VN.t7 134.75
R2890 VN.n3 VN.t4 134.75
R2891 VN.n25 VN.t6 134.75
R2892 VN.n34 VN.t2 134.75
R2893 VN.n30 VN.t1 134.75
R2894 VN.n52 VN.t0 134.75
R2895 VN.n26 VN.n25 97.2996
R2896 VN.n53 VN.n52 97.2996
R2897 VN.n19 VN.n1 55.0624
R2898 VN.n46 VN.n28 55.0624
R2899 VN VN.n53 52.4375
R2900 VN.n7 VN.n6 51.8291
R2901 VN.n34 VN.n33 51.8291
R2902 VN.n12 VN.n5 40.4934
R2903 VN.n13 VN.n12 40.4934
R2904 VN.n39 VN.n32 40.4934
R2905 VN.n40 VN.n39 40.4934
R2906 VN.n23 VN.n1 25.9244
R2907 VN.n50 VN.n28 25.9244
R2908 VN.n8 VN.n5 24.4675
R2909 VN.n14 VN.n13 24.4675
R2910 VN.n18 VN.n17 24.4675
R2911 VN.n19 VN.n18 24.4675
R2912 VN.n24 VN.n23 24.4675
R2913 VN.n35 VN.n32 24.4675
R2914 VN.n46 VN.n45 24.4675
R2915 VN.n45 VN.n44 24.4675
R2916 VN.n41 VN.n40 24.4675
R2917 VN.n51 VN.n50 24.4675
R2918 VN.n8 VN.n7 20.7975
R2919 VN.n14 VN.n3 20.7975
R2920 VN.n35 VN.n34 20.7975
R2921 VN.n41 VN.n30 20.7975
R2922 VN.n25 VN.n24 13.4574
R2923 VN.n52 VN.n51 13.4574
R2924 VN.n36 VN.n33 6.62497
R2925 VN.n9 VN.n6 6.62497
R2926 VN.n17 VN.n3 3.67055
R2927 VN.n44 VN.n30 3.67055
R2928 VN.n53 VN.n27 0.278367
R2929 VN.n26 VN.n0 0.278367
R2930 VN.n49 VN.n27 0.189894
R2931 VN.n49 VN.n48 0.189894
R2932 VN.n48 VN.n47 0.189894
R2933 VN.n47 VN.n29 0.189894
R2934 VN.n43 VN.n29 0.189894
R2935 VN.n43 VN.n42 0.189894
R2936 VN.n42 VN.n31 0.189894
R2937 VN.n38 VN.n31 0.189894
R2938 VN.n38 VN.n37 0.189894
R2939 VN.n37 VN.n36 0.189894
R2940 VN.n10 VN.n9 0.189894
R2941 VN.n11 VN.n10 0.189894
R2942 VN.n11 VN.n4 0.189894
R2943 VN.n15 VN.n4 0.189894
R2944 VN.n16 VN.n15 0.189894
R2945 VN.n16 VN.n2 0.189894
R2946 VN.n20 VN.n2 0.189894
R2947 VN.n21 VN.n20 0.189894
R2948 VN.n22 VN.n21 0.189894
R2949 VN.n22 VN.n0 0.189894
R2950 VN VN.n26 0.153454
R2951 VDD2.n2 VDD2.n1 65.4843
R2952 VDD2.n2 VDD2.n0 65.4843
R2953 VDD2 VDD2.n5 65.4815
R2954 VDD2.n4 VDD2.n3 64.3114
R2955 VDD2.n4 VDD2.n2 46.9179
R2956 VDD2.n5 VDD2.t5 1.40575
R2957 VDD2.n5 VDD2.t4 1.40575
R2958 VDD2.n3 VDD2.t7 1.40575
R2959 VDD2.n3 VDD2.t6 1.40575
R2960 VDD2.n1 VDD2.t3 1.40575
R2961 VDD2.n1 VDD2.t1 1.40575
R2962 VDD2.n0 VDD2.t2 1.40575
R2963 VDD2.n0 VDD2.t0 1.40575
R2964 VDD2 VDD2.n4 1.28714
C0 VDD2 VTAIL 8.834089f
C1 VP VTAIL 10.3618f
C2 VDD2 VDD1 1.73595f
C3 VP VDD1 10.4219f
C4 VN VTAIL 10.3477f
C5 VN VDD1 0.151616f
C6 VTAIL VDD1 8.78021f
C7 VDD2 VP 0.51119f
C8 VDD2 VN 10.0637f
C9 VP VN 7.94951f
C10 VDD2 B 5.426659f
C11 VDD1 B 5.854169f
C12 VTAIL B 11.674248f
C13 VN B 15.36585f
C14 VP B 13.912697f
C15 VDD2.t2 B 0.270885f
C16 VDD2.t0 B 0.270885f
C17 VDD2.n0 B 2.45332f
C18 VDD2.t3 B 0.270885f
C19 VDD2.t1 B 0.270885f
C20 VDD2.n1 B 2.45332f
C21 VDD2.n2 B 3.26227f
C22 VDD2.t7 B 0.270885f
C23 VDD2.t6 B 0.270885f
C24 VDD2.n3 B 2.44456f
C25 VDD2.n4 B 2.99328f
C26 VDD2.t5 B 0.270885f
C27 VDD2.t4 B 0.270885f
C28 VDD2.n5 B 2.45329f
C29 VN.n0 B 0.029192f
C30 VN.t6 B 2.15114f
C31 VN.n1 B 0.025249f
C32 VN.n2 B 0.022142f
C33 VN.t4 B 2.15114f
C34 VN.n3 B 0.754792f
C35 VN.n4 B 0.022142f
C36 VN.n5 B 0.044007f
C37 VN.t5 B 2.33314f
C38 VN.n6 B 0.794696f
C39 VN.t7 B 2.15114f
C40 VN.n7 B 0.825568f
C41 VN.n8 B 0.03821f
C42 VN.n9 B 0.212158f
C43 VN.n10 B 0.022142f
C44 VN.n11 B 0.022142f
C45 VN.n12 B 0.0179f
C46 VN.n13 B 0.044007f
C47 VN.n14 B 0.03821f
C48 VN.n15 B 0.022142f
C49 VN.n16 B 0.022142f
C50 VN.n17 B 0.023948f
C51 VN.n18 B 0.041267f
C52 VN.n19 B 0.038322f
C53 VN.n20 B 0.022142f
C54 VN.n21 B 0.022142f
C55 VN.n22 B 0.022142f
C56 VN.n23 B 0.042342f
C57 VN.n24 B 0.032098f
C58 VN.n25 B 0.831113f
C59 VN.n26 B 0.033407f
C60 VN.n27 B 0.029192f
C61 VN.t0 B 2.15114f
C62 VN.n28 B 0.025249f
C63 VN.n29 B 0.022142f
C64 VN.t1 B 2.15114f
C65 VN.n30 B 0.754792f
C66 VN.n31 B 0.022142f
C67 VN.n32 B 0.044007f
C68 VN.t3 B 2.33314f
C69 VN.n33 B 0.794696f
C70 VN.t2 B 2.15114f
C71 VN.n34 B 0.825568f
C72 VN.n35 B 0.03821f
C73 VN.n36 B 0.212158f
C74 VN.n37 B 0.022142f
C75 VN.n38 B 0.022142f
C76 VN.n39 B 0.0179f
C77 VN.n40 B 0.044007f
C78 VN.n41 B 0.03821f
C79 VN.n42 B 0.022142f
C80 VN.n43 B 0.022142f
C81 VN.n44 B 0.023948f
C82 VN.n45 B 0.041267f
C83 VN.n46 B 0.038322f
C84 VN.n47 B 0.022142f
C85 VN.n48 B 0.022142f
C86 VN.n49 B 0.022142f
C87 VN.n50 B 0.042342f
C88 VN.n51 B 0.032098f
C89 VN.n52 B 0.831113f
C90 VN.n53 B 1.31971f
C91 VDD1.t1 B 0.273883f
C92 VDD1.t2 B 0.273883f
C93 VDD1.n0 B 2.48149f
C94 VDD1.t5 B 0.273883f
C95 VDD1.t0 B 0.273883f
C96 VDD1.n1 B 2.48047f
C97 VDD1.t4 B 0.273883f
C98 VDD1.t6 B 0.273883f
C99 VDD1.n2 B 2.48047f
C100 VDD1.n3 B 3.34957f
C101 VDD1.t3 B 0.273883f
C102 VDD1.t7 B 0.273883f
C103 VDD1.n4 B 2.4716f
C104 VDD1.n5 B 3.05685f
C105 VTAIL.t6 B 0.213988f
C106 VTAIL.t1 B 0.213988f
C107 VTAIL.n0 B 1.87846f
C108 VTAIL.n1 B 0.336194f
C109 VTAIL.n2 B 0.026106f
C110 VTAIL.n3 B 0.019219f
C111 VTAIL.n4 B 0.010631f
C112 VTAIL.n5 B 0.02441f
C113 VTAIL.n6 B 0.010935f
C114 VTAIL.n7 B 0.019219f
C115 VTAIL.n8 B 0.010327f
C116 VTAIL.n9 B 0.02441f
C117 VTAIL.n10 B 0.010935f
C118 VTAIL.n11 B 0.019219f
C119 VTAIL.n12 B 0.010327f
C120 VTAIL.n13 B 0.02441f
C121 VTAIL.n14 B 0.010935f
C122 VTAIL.n15 B 0.019219f
C123 VTAIL.n16 B 0.010327f
C124 VTAIL.n17 B 0.02441f
C125 VTAIL.n18 B 0.010935f
C126 VTAIL.n19 B 0.019219f
C127 VTAIL.n20 B 0.010327f
C128 VTAIL.n21 B 0.02441f
C129 VTAIL.n22 B 0.010935f
C130 VTAIL.n23 B 0.019219f
C131 VTAIL.n24 B 0.010327f
C132 VTAIL.n25 B 0.018307f
C133 VTAIL.n26 B 0.01442f
C134 VTAIL.t0 B 0.040189f
C135 VTAIL.n27 B 0.120964f
C136 VTAIL.n28 B 1.17024f
C137 VTAIL.n29 B 0.010327f
C138 VTAIL.n30 B 0.010935f
C139 VTAIL.n31 B 0.02441f
C140 VTAIL.n32 B 0.02441f
C141 VTAIL.n33 B 0.010935f
C142 VTAIL.n34 B 0.010327f
C143 VTAIL.n35 B 0.019219f
C144 VTAIL.n36 B 0.019219f
C145 VTAIL.n37 B 0.010327f
C146 VTAIL.n38 B 0.010935f
C147 VTAIL.n39 B 0.02441f
C148 VTAIL.n40 B 0.02441f
C149 VTAIL.n41 B 0.010935f
C150 VTAIL.n42 B 0.010327f
C151 VTAIL.n43 B 0.019219f
C152 VTAIL.n44 B 0.019219f
C153 VTAIL.n45 B 0.010327f
C154 VTAIL.n46 B 0.010935f
C155 VTAIL.n47 B 0.02441f
C156 VTAIL.n48 B 0.02441f
C157 VTAIL.n49 B 0.010935f
C158 VTAIL.n50 B 0.010327f
C159 VTAIL.n51 B 0.019219f
C160 VTAIL.n52 B 0.019219f
C161 VTAIL.n53 B 0.010327f
C162 VTAIL.n54 B 0.010935f
C163 VTAIL.n55 B 0.02441f
C164 VTAIL.n56 B 0.02441f
C165 VTAIL.n57 B 0.010935f
C166 VTAIL.n58 B 0.010327f
C167 VTAIL.n59 B 0.019219f
C168 VTAIL.n60 B 0.019219f
C169 VTAIL.n61 B 0.010327f
C170 VTAIL.n62 B 0.010935f
C171 VTAIL.n63 B 0.02441f
C172 VTAIL.n64 B 0.02441f
C173 VTAIL.n65 B 0.010935f
C174 VTAIL.n66 B 0.010327f
C175 VTAIL.n67 B 0.019219f
C176 VTAIL.n68 B 0.019219f
C177 VTAIL.n69 B 0.010327f
C178 VTAIL.n70 B 0.010327f
C179 VTAIL.n71 B 0.010935f
C180 VTAIL.n72 B 0.02441f
C181 VTAIL.n73 B 0.02441f
C182 VTAIL.n74 B 0.051238f
C183 VTAIL.n75 B 0.010631f
C184 VTAIL.n76 B 0.010327f
C185 VTAIL.n77 B 0.048886f
C186 VTAIL.n78 B 0.028636f
C187 VTAIL.n79 B 0.200182f
C188 VTAIL.n80 B 0.026106f
C189 VTAIL.n81 B 0.019219f
C190 VTAIL.n82 B 0.010631f
C191 VTAIL.n83 B 0.02441f
C192 VTAIL.n84 B 0.010935f
C193 VTAIL.n85 B 0.019219f
C194 VTAIL.n86 B 0.010327f
C195 VTAIL.n87 B 0.02441f
C196 VTAIL.n88 B 0.010935f
C197 VTAIL.n89 B 0.019219f
C198 VTAIL.n90 B 0.010327f
C199 VTAIL.n91 B 0.02441f
C200 VTAIL.n92 B 0.010935f
C201 VTAIL.n93 B 0.019219f
C202 VTAIL.n94 B 0.010327f
C203 VTAIL.n95 B 0.02441f
C204 VTAIL.n96 B 0.010935f
C205 VTAIL.n97 B 0.019219f
C206 VTAIL.n98 B 0.010327f
C207 VTAIL.n99 B 0.02441f
C208 VTAIL.n100 B 0.010935f
C209 VTAIL.n101 B 0.019219f
C210 VTAIL.n102 B 0.010327f
C211 VTAIL.n103 B 0.018307f
C212 VTAIL.n104 B 0.01442f
C213 VTAIL.t8 B 0.040189f
C214 VTAIL.n105 B 0.120964f
C215 VTAIL.n106 B 1.17024f
C216 VTAIL.n107 B 0.010327f
C217 VTAIL.n108 B 0.010935f
C218 VTAIL.n109 B 0.02441f
C219 VTAIL.n110 B 0.02441f
C220 VTAIL.n111 B 0.010935f
C221 VTAIL.n112 B 0.010327f
C222 VTAIL.n113 B 0.019219f
C223 VTAIL.n114 B 0.019219f
C224 VTAIL.n115 B 0.010327f
C225 VTAIL.n116 B 0.010935f
C226 VTAIL.n117 B 0.02441f
C227 VTAIL.n118 B 0.02441f
C228 VTAIL.n119 B 0.010935f
C229 VTAIL.n120 B 0.010327f
C230 VTAIL.n121 B 0.019219f
C231 VTAIL.n122 B 0.019219f
C232 VTAIL.n123 B 0.010327f
C233 VTAIL.n124 B 0.010935f
C234 VTAIL.n125 B 0.02441f
C235 VTAIL.n126 B 0.02441f
C236 VTAIL.n127 B 0.010935f
C237 VTAIL.n128 B 0.010327f
C238 VTAIL.n129 B 0.019219f
C239 VTAIL.n130 B 0.019219f
C240 VTAIL.n131 B 0.010327f
C241 VTAIL.n132 B 0.010935f
C242 VTAIL.n133 B 0.02441f
C243 VTAIL.n134 B 0.02441f
C244 VTAIL.n135 B 0.010935f
C245 VTAIL.n136 B 0.010327f
C246 VTAIL.n137 B 0.019219f
C247 VTAIL.n138 B 0.019219f
C248 VTAIL.n139 B 0.010327f
C249 VTAIL.n140 B 0.010935f
C250 VTAIL.n141 B 0.02441f
C251 VTAIL.n142 B 0.02441f
C252 VTAIL.n143 B 0.010935f
C253 VTAIL.n144 B 0.010327f
C254 VTAIL.n145 B 0.019219f
C255 VTAIL.n146 B 0.019219f
C256 VTAIL.n147 B 0.010327f
C257 VTAIL.n148 B 0.010327f
C258 VTAIL.n149 B 0.010935f
C259 VTAIL.n150 B 0.02441f
C260 VTAIL.n151 B 0.02441f
C261 VTAIL.n152 B 0.051238f
C262 VTAIL.n153 B 0.010631f
C263 VTAIL.n154 B 0.010327f
C264 VTAIL.n155 B 0.048886f
C265 VTAIL.n156 B 0.028636f
C266 VTAIL.n157 B 0.200182f
C267 VTAIL.t15 B 0.213988f
C268 VTAIL.t13 B 0.213988f
C269 VTAIL.n158 B 1.87846f
C270 VTAIL.n159 B 0.484739f
C271 VTAIL.n160 B 0.026106f
C272 VTAIL.n161 B 0.019219f
C273 VTAIL.n162 B 0.010631f
C274 VTAIL.n163 B 0.02441f
C275 VTAIL.n164 B 0.010935f
C276 VTAIL.n165 B 0.019219f
C277 VTAIL.n166 B 0.010327f
C278 VTAIL.n167 B 0.02441f
C279 VTAIL.n168 B 0.010935f
C280 VTAIL.n169 B 0.019219f
C281 VTAIL.n170 B 0.010327f
C282 VTAIL.n171 B 0.02441f
C283 VTAIL.n172 B 0.010935f
C284 VTAIL.n173 B 0.019219f
C285 VTAIL.n174 B 0.010327f
C286 VTAIL.n175 B 0.02441f
C287 VTAIL.n176 B 0.010935f
C288 VTAIL.n177 B 0.019219f
C289 VTAIL.n178 B 0.010327f
C290 VTAIL.n179 B 0.02441f
C291 VTAIL.n180 B 0.010935f
C292 VTAIL.n181 B 0.019219f
C293 VTAIL.n182 B 0.010327f
C294 VTAIL.n183 B 0.018307f
C295 VTAIL.n184 B 0.01442f
C296 VTAIL.t11 B 0.040189f
C297 VTAIL.n185 B 0.120964f
C298 VTAIL.n186 B 1.17024f
C299 VTAIL.n187 B 0.010327f
C300 VTAIL.n188 B 0.010935f
C301 VTAIL.n189 B 0.02441f
C302 VTAIL.n190 B 0.02441f
C303 VTAIL.n191 B 0.010935f
C304 VTAIL.n192 B 0.010327f
C305 VTAIL.n193 B 0.019219f
C306 VTAIL.n194 B 0.019219f
C307 VTAIL.n195 B 0.010327f
C308 VTAIL.n196 B 0.010935f
C309 VTAIL.n197 B 0.02441f
C310 VTAIL.n198 B 0.02441f
C311 VTAIL.n199 B 0.010935f
C312 VTAIL.n200 B 0.010327f
C313 VTAIL.n201 B 0.019219f
C314 VTAIL.n202 B 0.019219f
C315 VTAIL.n203 B 0.010327f
C316 VTAIL.n204 B 0.010935f
C317 VTAIL.n205 B 0.02441f
C318 VTAIL.n206 B 0.02441f
C319 VTAIL.n207 B 0.010935f
C320 VTAIL.n208 B 0.010327f
C321 VTAIL.n209 B 0.019219f
C322 VTAIL.n210 B 0.019219f
C323 VTAIL.n211 B 0.010327f
C324 VTAIL.n212 B 0.010935f
C325 VTAIL.n213 B 0.02441f
C326 VTAIL.n214 B 0.02441f
C327 VTAIL.n215 B 0.010935f
C328 VTAIL.n216 B 0.010327f
C329 VTAIL.n217 B 0.019219f
C330 VTAIL.n218 B 0.019219f
C331 VTAIL.n219 B 0.010327f
C332 VTAIL.n220 B 0.010935f
C333 VTAIL.n221 B 0.02441f
C334 VTAIL.n222 B 0.02441f
C335 VTAIL.n223 B 0.010935f
C336 VTAIL.n224 B 0.010327f
C337 VTAIL.n225 B 0.019219f
C338 VTAIL.n226 B 0.019219f
C339 VTAIL.n227 B 0.010327f
C340 VTAIL.n228 B 0.010327f
C341 VTAIL.n229 B 0.010935f
C342 VTAIL.n230 B 0.02441f
C343 VTAIL.n231 B 0.02441f
C344 VTAIL.n232 B 0.051238f
C345 VTAIL.n233 B 0.010631f
C346 VTAIL.n234 B 0.010327f
C347 VTAIL.n235 B 0.048886f
C348 VTAIL.n236 B 0.028636f
C349 VTAIL.n237 B 1.3365f
C350 VTAIL.n238 B 0.026106f
C351 VTAIL.n239 B 0.019219f
C352 VTAIL.n240 B 0.010631f
C353 VTAIL.n241 B 0.02441f
C354 VTAIL.n242 B 0.010327f
C355 VTAIL.n243 B 0.010935f
C356 VTAIL.n244 B 0.019219f
C357 VTAIL.n245 B 0.010327f
C358 VTAIL.n246 B 0.02441f
C359 VTAIL.n247 B 0.010935f
C360 VTAIL.n248 B 0.019219f
C361 VTAIL.n249 B 0.010327f
C362 VTAIL.n250 B 0.02441f
C363 VTAIL.n251 B 0.010935f
C364 VTAIL.n252 B 0.019219f
C365 VTAIL.n253 B 0.010327f
C366 VTAIL.n254 B 0.02441f
C367 VTAIL.n255 B 0.010935f
C368 VTAIL.n256 B 0.019219f
C369 VTAIL.n257 B 0.010327f
C370 VTAIL.n258 B 0.02441f
C371 VTAIL.n259 B 0.010935f
C372 VTAIL.n260 B 0.019219f
C373 VTAIL.n261 B 0.010327f
C374 VTAIL.n262 B 0.018307f
C375 VTAIL.n263 B 0.01442f
C376 VTAIL.t7 B 0.040189f
C377 VTAIL.n264 B 0.120964f
C378 VTAIL.n265 B 1.17024f
C379 VTAIL.n266 B 0.010327f
C380 VTAIL.n267 B 0.010935f
C381 VTAIL.n268 B 0.02441f
C382 VTAIL.n269 B 0.02441f
C383 VTAIL.n270 B 0.010935f
C384 VTAIL.n271 B 0.010327f
C385 VTAIL.n272 B 0.019219f
C386 VTAIL.n273 B 0.019219f
C387 VTAIL.n274 B 0.010327f
C388 VTAIL.n275 B 0.010935f
C389 VTAIL.n276 B 0.02441f
C390 VTAIL.n277 B 0.02441f
C391 VTAIL.n278 B 0.010935f
C392 VTAIL.n279 B 0.010327f
C393 VTAIL.n280 B 0.019219f
C394 VTAIL.n281 B 0.019219f
C395 VTAIL.n282 B 0.010327f
C396 VTAIL.n283 B 0.010935f
C397 VTAIL.n284 B 0.02441f
C398 VTAIL.n285 B 0.02441f
C399 VTAIL.n286 B 0.010935f
C400 VTAIL.n287 B 0.010327f
C401 VTAIL.n288 B 0.019219f
C402 VTAIL.n289 B 0.019219f
C403 VTAIL.n290 B 0.010327f
C404 VTAIL.n291 B 0.010935f
C405 VTAIL.n292 B 0.02441f
C406 VTAIL.n293 B 0.02441f
C407 VTAIL.n294 B 0.010935f
C408 VTAIL.n295 B 0.010327f
C409 VTAIL.n296 B 0.019219f
C410 VTAIL.n297 B 0.019219f
C411 VTAIL.n298 B 0.010327f
C412 VTAIL.n299 B 0.010935f
C413 VTAIL.n300 B 0.02441f
C414 VTAIL.n301 B 0.02441f
C415 VTAIL.n302 B 0.010935f
C416 VTAIL.n303 B 0.010327f
C417 VTAIL.n304 B 0.019219f
C418 VTAIL.n305 B 0.019219f
C419 VTAIL.n306 B 0.010327f
C420 VTAIL.n307 B 0.010935f
C421 VTAIL.n308 B 0.02441f
C422 VTAIL.n309 B 0.02441f
C423 VTAIL.n310 B 0.051238f
C424 VTAIL.n311 B 0.010631f
C425 VTAIL.n312 B 0.010327f
C426 VTAIL.n313 B 0.048886f
C427 VTAIL.n314 B 0.028636f
C428 VTAIL.n315 B 1.3365f
C429 VTAIL.t5 B 0.213988f
C430 VTAIL.t3 B 0.213988f
C431 VTAIL.n316 B 1.87847f
C432 VTAIL.n317 B 0.48473f
C433 VTAIL.n318 B 0.026106f
C434 VTAIL.n319 B 0.019219f
C435 VTAIL.n320 B 0.010631f
C436 VTAIL.n321 B 0.02441f
C437 VTAIL.n322 B 0.010327f
C438 VTAIL.n323 B 0.010935f
C439 VTAIL.n324 B 0.019219f
C440 VTAIL.n325 B 0.010327f
C441 VTAIL.n326 B 0.02441f
C442 VTAIL.n327 B 0.010935f
C443 VTAIL.n328 B 0.019219f
C444 VTAIL.n329 B 0.010327f
C445 VTAIL.n330 B 0.02441f
C446 VTAIL.n331 B 0.010935f
C447 VTAIL.n332 B 0.019219f
C448 VTAIL.n333 B 0.010327f
C449 VTAIL.n334 B 0.02441f
C450 VTAIL.n335 B 0.010935f
C451 VTAIL.n336 B 0.019219f
C452 VTAIL.n337 B 0.010327f
C453 VTAIL.n338 B 0.02441f
C454 VTAIL.n339 B 0.010935f
C455 VTAIL.n340 B 0.019219f
C456 VTAIL.n341 B 0.010327f
C457 VTAIL.n342 B 0.018307f
C458 VTAIL.n343 B 0.01442f
C459 VTAIL.t4 B 0.040189f
C460 VTAIL.n344 B 0.120964f
C461 VTAIL.n345 B 1.17024f
C462 VTAIL.n346 B 0.010327f
C463 VTAIL.n347 B 0.010935f
C464 VTAIL.n348 B 0.02441f
C465 VTAIL.n349 B 0.02441f
C466 VTAIL.n350 B 0.010935f
C467 VTAIL.n351 B 0.010327f
C468 VTAIL.n352 B 0.019219f
C469 VTAIL.n353 B 0.019219f
C470 VTAIL.n354 B 0.010327f
C471 VTAIL.n355 B 0.010935f
C472 VTAIL.n356 B 0.02441f
C473 VTAIL.n357 B 0.02441f
C474 VTAIL.n358 B 0.010935f
C475 VTAIL.n359 B 0.010327f
C476 VTAIL.n360 B 0.019219f
C477 VTAIL.n361 B 0.019219f
C478 VTAIL.n362 B 0.010327f
C479 VTAIL.n363 B 0.010935f
C480 VTAIL.n364 B 0.02441f
C481 VTAIL.n365 B 0.02441f
C482 VTAIL.n366 B 0.010935f
C483 VTAIL.n367 B 0.010327f
C484 VTAIL.n368 B 0.019219f
C485 VTAIL.n369 B 0.019219f
C486 VTAIL.n370 B 0.010327f
C487 VTAIL.n371 B 0.010935f
C488 VTAIL.n372 B 0.02441f
C489 VTAIL.n373 B 0.02441f
C490 VTAIL.n374 B 0.010935f
C491 VTAIL.n375 B 0.010327f
C492 VTAIL.n376 B 0.019219f
C493 VTAIL.n377 B 0.019219f
C494 VTAIL.n378 B 0.010327f
C495 VTAIL.n379 B 0.010935f
C496 VTAIL.n380 B 0.02441f
C497 VTAIL.n381 B 0.02441f
C498 VTAIL.n382 B 0.010935f
C499 VTAIL.n383 B 0.010327f
C500 VTAIL.n384 B 0.019219f
C501 VTAIL.n385 B 0.019219f
C502 VTAIL.n386 B 0.010327f
C503 VTAIL.n387 B 0.010935f
C504 VTAIL.n388 B 0.02441f
C505 VTAIL.n389 B 0.02441f
C506 VTAIL.n390 B 0.051238f
C507 VTAIL.n391 B 0.010631f
C508 VTAIL.n392 B 0.010327f
C509 VTAIL.n393 B 0.048886f
C510 VTAIL.n394 B 0.028636f
C511 VTAIL.n395 B 0.200182f
C512 VTAIL.n396 B 0.026106f
C513 VTAIL.n397 B 0.019219f
C514 VTAIL.n398 B 0.010631f
C515 VTAIL.n399 B 0.02441f
C516 VTAIL.n400 B 0.010327f
C517 VTAIL.n401 B 0.010935f
C518 VTAIL.n402 B 0.019219f
C519 VTAIL.n403 B 0.010327f
C520 VTAIL.n404 B 0.02441f
C521 VTAIL.n405 B 0.010935f
C522 VTAIL.n406 B 0.019219f
C523 VTAIL.n407 B 0.010327f
C524 VTAIL.n408 B 0.02441f
C525 VTAIL.n409 B 0.010935f
C526 VTAIL.n410 B 0.019219f
C527 VTAIL.n411 B 0.010327f
C528 VTAIL.n412 B 0.02441f
C529 VTAIL.n413 B 0.010935f
C530 VTAIL.n414 B 0.019219f
C531 VTAIL.n415 B 0.010327f
C532 VTAIL.n416 B 0.02441f
C533 VTAIL.n417 B 0.010935f
C534 VTAIL.n418 B 0.019219f
C535 VTAIL.n419 B 0.010327f
C536 VTAIL.n420 B 0.018307f
C537 VTAIL.n421 B 0.01442f
C538 VTAIL.t10 B 0.040189f
C539 VTAIL.n422 B 0.120964f
C540 VTAIL.n423 B 1.17024f
C541 VTAIL.n424 B 0.010327f
C542 VTAIL.n425 B 0.010935f
C543 VTAIL.n426 B 0.02441f
C544 VTAIL.n427 B 0.02441f
C545 VTAIL.n428 B 0.010935f
C546 VTAIL.n429 B 0.010327f
C547 VTAIL.n430 B 0.019219f
C548 VTAIL.n431 B 0.019219f
C549 VTAIL.n432 B 0.010327f
C550 VTAIL.n433 B 0.010935f
C551 VTAIL.n434 B 0.02441f
C552 VTAIL.n435 B 0.02441f
C553 VTAIL.n436 B 0.010935f
C554 VTAIL.n437 B 0.010327f
C555 VTAIL.n438 B 0.019219f
C556 VTAIL.n439 B 0.019219f
C557 VTAIL.n440 B 0.010327f
C558 VTAIL.n441 B 0.010935f
C559 VTAIL.n442 B 0.02441f
C560 VTAIL.n443 B 0.02441f
C561 VTAIL.n444 B 0.010935f
C562 VTAIL.n445 B 0.010327f
C563 VTAIL.n446 B 0.019219f
C564 VTAIL.n447 B 0.019219f
C565 VTAIL.n448 B 0.010327f
C566 VTAIL.n449 B 0.010935f
C567 VTAIL.n450 B 0.02441f
C568 VTAIL.n451 B 0.02441f
C569 VTAIL.n452 B 0.010935f
C570 VTAIL.n453 B 0.010327f
C571 VTAIL.n454 B 0.019219f
C572 VTAIL.n455 B 0.019219f
C573 VTAIL.n456 B 0.010327f
C574 VTAIL.n457 B 0.010935f
C575 VTAIL.n458 B 0.02441f
C576 VTAIL.n459 B 0.02441f
C577 VTAIL.n460 B 0.010935f
C578 VTAIL.n461 B 0.010327f
C579 VTAIL.n462 B 0.019219f
C580 VTAIL.n463 B 0.019219f
C581 VTAIL.n464 B 0.010327f
C582 VTAIL.n465 B 0.010935f
C583 VTAIL.n466 B 0.02441f
C584 VTAIL.n467 B 0.02441f
C585 VTAIL.n468 B 0.051238f
C586 VTAIL.n469 B 0.010631f
C587 VTAIL.n470 B 0.010327f
C588 VTAIL.n471 B 0.048886f
C589 VTAIL.n472 B 0.028636f
C590 VTAIL.n473 B 0.200182f
C591 VTAIL.t14 B 0.213988f
C592 VTAIL.t9 B 0.213988f
C593 VTAIL.n474 B 1.87847f
C594 VTAIL.n475 B 0.48473f
C595 VTAIL.n476 B 0.026106f
C596 VTAIL.n477 B 0.019219f
C597 VTAIL.n478 B 0.010631f
C598 VTAIL.n479 B 0.02441f
C599 VTAIL.n480 B 0.010327f
C600 VTAIL.n481 B 0.010935f
C601 VTAIL.n482 B 0.019219f
C602 VTAIL.n483 B 0.010327f
C603 VTAIL.n484 B 0.02441f
C604 VTAIL.n485 B 0.010935f
C605 VTAIL.n486 B 0.019219f
C606 VTAIL.n487 B 0.010327f
C607 VTAIL.n488 B 0.02441f
C608 VTAIL.n489 B 0.010935f
C609 VTAIL.n490 B 0.019219f
C610 VTAIL.n491 B 0.010327f
C611 VTAIL.n492 B 0.02441f
C612 VTAIL.n493 B 0.010935f
C613 VTAIL.n494 B 0.019219f
C614 VTAIL.n495 B 0.010327f
C615 VTAIL.n496 B 0.02441f
C616 VTAIL.n497 B 0.010935f
C617 VTAIL.n498 B 0.019219f
C618 VTAIL.n499 B 0.010327f
C619 VTAIL.n500 B 0.018307f
C620 VTAIL.n501 B 0.01442f
C621 VTAIL.t12 B 0.040189f
C622 VTAIL.n502 B 0.120964f
C623 VTAIL.n503 B 1.17024f
C624 VTAIL.n504 B 0.010327f
C625 VTAIL.n505 B 0.010935f
C626 VTAIL.n506 B 0.02441f
C627 VTAIL.n507 B 0.02441f
C628 VTAIL.n508 B 0.010935f
C629 VTAIL.n509 B 0.010327f
C630 VTAIL.n510 B 0.019219f
C631 VTAIL.n511 B 0.019219f
C632 VTAIL.n512 B 0.010327f
C633 VTAIL.n513 B 0.010935f
C634 VTAIL.n514 B 0.02441f
C635 VTAIL.n515 B 0.02441f
C636 VTAIL.n516 B 0.010935f
C637 VTAIL.n517 B 0.010327f
C638 VTAIL.n518 B 0.019219f
C639 VTAIL.n519 B 0.019219f
C640 VTAIL.n520 B 0.010327f
C641 VTAIL.n521 B 0.010935f
C642 VTAIL.n522 B 0.02441f
C643 VTAIL.n523 B 0.02441f
C644 VTAIL.n524 B 0.010935f
C645 VTAIL.n525 B 0.010327f
C646 VTAIL.n526 B 0.019219f
C647 VTAIL.n527 B 0.019219f
C648 VTAIL.n528 B 0.010327f
C649 VTAIL.n529 B 0.010935f
C650 VTAIL.n530 B 0.02441f
C651 VTAIL.n531 B 0.02441f
C652 VTAIL.n532 B 0.010935f
C653 VTAIL.n533 B 0.010327f
C654 VTAIL.n534 B 0.019219f
C655 VTAIL.n535 B 0.019219f
C656 VTAIL.n536 B 0.010327f
C657 VTAIL.n537 B 0.010935f
C658 VTAIL.n538 B 0.02441f
C659 VTAIL.n539 B 0.02441f
C660 VTAIL.n540 B 0.010935f
C661 VTAIL.n541 B 0.010327f
C662 VTAIL.n542 B 0.019219f
C663 VTAIL.n543 B 0.019219f
C664 VTAIL.n544 B 0.010327f
C665 VTAIL.n545 B 0.010935f
C666 VTAIL.n546 B 0.02441f
C667 VTAIL.n547 B 0.02441f
C668 VTAIL.n548 B 0.051238f
C669 VTAIL.n549 B 0.010631f
C670 VTAIL.n550 B 0.010327f
C671 VTAIL.n551 B 0.048886f
C672 VTAIL.n552 B 0.028636f
C673 VTAIL.n553 B 1.3365f
C674 VTAIL.n554 B 0.026106f
C675 VTAIL.n555 B 0.019219f
C676 VTAIL.n556 B 0.010631f
C677 VTAIL.n557 B 0.02441f
C678 VTAIL.n558 B 0.010935f
C679 VTAIL.n559 B 0.019219f
C680 VTAIL.n560 B 0.010327f
C681 VTAIL.n561 B 0.02441f
C682 VTAIL.n562 B 0.010935f
C683 VTAIL.n563 B 0.019219f
C684 VTAIL.n564 B 0.010327f
C685 VTAIL.n565 B 0.02441f
C686 VTAIL.n566 B 0.010935f
C687 VTAIL.n567 B 0.019219f
C688 VTAIL.n568 B 0.010327f
C689 VTAIL.n569 B 0.02441f
C690 VTAIL.n570 B 0.010935f
C691 VTAIL.n571 B 0.019219f
C692 VTAIL.n572 B 0.010327f
C693 VTAIL.n573 B 0.02441f
C694 VTAIL.n574 B 0.010935f
C695 VTAIL.n575 B 0.019219f
C696 VTAIL.n576 B 0.010327f
C697 VTAIL.n577 B 0.018307f
C698 VTAIL.n578 B 0.01442f
C699 VTAIL.t2 B 0.040189f
C700 VTAIL.n579 B 0.120964f
C701 VTAIL.n580 B 1.17024f
C702 VTAIL.n581 B 0.010327f
C703 VTAIL.n582 B 0.010935f
C704 VTAIL.n583 B 0.02441f
C705 VTAIL.n584 B 0.02441f
C706 VTAIL.n585 B 0.010935f
C707 VTAIL.n586 B 0.010327f
C708 VTAIL.n587 B 0.019219f
C709 VTAIL.n588 B 0.019219f
C710 VTAIL.n589 B 0.010327f
C711 VTAIL.n590 B 0.010935f
C712 VTAIL.n591 B 0.02441f
C713 VTAIL.n592 B 0.02441f
C714 VTAIL.n593 B 0.010935f
C715 VTAIL.n594 B 0.010327f
C716 VTAIL.n595 B 0.019219f
C717 VTAIL.n596 B 0.019219f
C718 VTAIL.n597 B 0.010327f
C719 VTAIL.n598 B 0.010935f
C720 VTAIL.n599 B 0.02441f
C721 VTAIL.n600 B 0.02441f
C722 VTAIL.n601 B 0.010935f
C723 VTAIL.n602 B 0.010327f
C724 VTAIL.n603 B 0.019219f
C725 VTAIL.n604 B 0.019219f
C726 VTAIL.n605 B 0.010327f
C727 VTAIL.n606 B 0.010935f
C728 VTAIL.n607 B 0.02441f
C729 VTAIL.n608 B 0.02441f
C730 VTAIL.n609 B 0.010935f
C731 VTAIL.n610 B 0.010327f
C732 VTAIL.n611 B 0.019219f
C733 VTAIL.n612 B 0.019219f
C734 VTAIL.n613 B 0.010327f
C735 VTAIL.n614 B 0.010935f
C736 VTAIL.n615 B 0.02441f
C737 VTAIL.n616 B 0.02441f
C738 VTAIL.n617 B 0.010935f
C739 VTAIL.n618 B 0.010327f
C740 VTAIL.n619 B 0.019219f
C741 VTAIL.n620 B 0.019219f
C742 VTAIL.n621 B 0.010327f
C743 VTAIL.n622 B 0.010327f
C744 VTAIL.n623 B 0.010935f
C745 VTAIL.n624 B 0.02441f
C746 VTAIL.n625 B 0.02441f
C747 VTAIL.n626 B 0.051238f
C748 VTAIL.n627 B 0.010631f
C749 VTAIL.n628 B 0.010327f
C750 VTAIL.n629 B 0.048886f
C751 VTAIL.n630 B 0.028636f
C752 VTAIL.n631 B 1.3329f
C753 VP.n0 B 0.029637f
C754 VP.t1 B 2.18395f
C755 VP.n1 B 0.025635f
C756 VP.n2 B 0.02248f
C757 VP.t3 B 2.18395f
C758 VP.n3 B 0.766304f
C759 VP.n4 B 0.02248f
C760 VP.n5 B 0.044678f
C761 VP.n6 B 0.02248f
C762 VP.t7 B 2.18395f
C763 VP.n7 B 0.038906f
C764 VP.n8 B 0.02248f
C765 VP.t2 B 2.18395f
C766 VP.n9 B 0.843788f
C767 VP.n10 B 0.029637f
C768 VP.t0 B 2.18395f
C769 VP.n11 B 0.025635f
C770 VP.n12 B 0.02248f
C771 VP.t4 B 2.18395f
C772 VP.n13 B 0.766304f
C773 VP.n14 B 0.02248f
C774 VP.n15 B 0.044678f
C775 VP.t6 B 2.36872f
C776 VP.n16 B 0.806816f
C777 VP.t5 B 2.18395f
C778 VP.n17 B 0.838158f
C779 VP.n18 B 0.038793f
C780 VP.n19 B 0.215394f
C781 VP.n20 B 0.02248f
C782 VP.n21 B 0.02248f
C783 VP.n22 B 0.018173f
C784 VP.n23 B 0.044678f
C785 VP.n24 B 0.038793f
C786 VP.n25 B 0.02248f
C787 VP.n26 B 0.02248f
C788 VP.n27 B 0.024313f
C789 VP.n28 B 0.041896f
C790 VP.n29 B 0.038906f
C791 VP.n30 B 0.02248f
C792 VP.n31 B 0.02248f
C793 VP.n32 B 0.02248f
C794 VP.n33 B 0.042988f
C795 VP.n34 B 0.032587f
C796 VP.n35 B 0.843788f
C797 VP.n36 B 1.32784f
C798 VP.n37 B 1.34333f
C799 VP.n38 B 0.029637f
C800 VP.n39 B 0.032587f
C801 VP.n40 B 0.042988f
C802 VP.n41 B 0.025635f
C803 VP.n42 B 0.02248f
C804 VP.n43 B 0.02248f
C805 VP.n44 B 0.02248f
C806 VP.n45 B 0.041896f
C807 VP.n46 B 0.024313f
C808 VP.n47 B 0.766304f
C809 VP.n48 B 0.038793f
C810 VP.n49 B 0.02248f
C811 VP.n50 B 0.02248f
C812 VP.n51 B 0.02248f
C813 VP.n52 B 0.018173f
C814 VP.n53 B 0.044678f
C815 VP.n54 B 0.038793f
C816 VP.n55 B 0.02248f
C817 VP.n56 B 0.02248f
C818 VP.n57 B 0.024313f
C819 VP.n58 B 0.041896f
C820 VP.n59 B 0.038906f
C821 VP.n60 B 0.02248f
C822 VP.n61 B 0.02248f
C823 VP.n62 B 0.02248f
C824 VP.n63 B 0.042988f
C825 VP.n64 B 0.032587f
C826 VP.n65 B 0.843788f
C827 VP.n66 B 0.033916f
.ends

