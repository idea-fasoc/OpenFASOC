* NGSPICE file created from diff_pair_sample_1132.ext - technology: sky130A

.subckt diff_pair_sample_1132 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=0 ps=0 w=8.04 l=0.23
X1 B.t8 B.t6 B.t7 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=0 ps=0 w=8.04 l=0.23
X2 VDD1.t3 VP.t0 VTAIL.t6 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=1.3266 pd=8.37 as=3.1356 ps=16.86 w=8.04 l=0.23
X3 VTAIL.t4 VP.t1 VDD1.t2 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=1.3266 ps=8.37 w=8.04 l=0.23
X4 B.t5 B.t3 B.t4 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=0 ps=0 w=8.04 l=0.23
X5 VDD1.t1 VP.t2 VTAIL.t5 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=1.3266 pd=8.37 as=3.1356 ps=16.86 w=8.04 l=0.23
X6 VTAIL.t3 VN.t0 VDD2.t3 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=1.3266 ps=8.37 w=8.04 l=0.23
X7 VTAIL.t7 VP.t3 VDD1.t0 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=1.3266 ps=8.37 w=8.04 l=0.23
X8 VTAIL.t2 VN.t1 VDD2.t2 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=1.3266 ps=8.37 w=8.04 l=0.23
X9 VDD2.t1 VN.t2 VTAIL.t1 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=1.3266 pd=8.37 as=3.1356 ps=16.86 w=8.04 l=0.23
X10 VDD2.t0 VN.t3 VTAIL.t0 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=1.3266 pd=8.37 as=3.1356 ps=16.86 w=8.04 l=0.23
X11 B.t2 B.t0 B.t1 w_n1306_n2580# sky130_fd_pr__pfet_01v8 ad=3.1356 pd=16.86 as=0 ps=0 w=8.04 l=0.23
R0 B.n77 B.t3 1070.94
R1 B.n85 B.t0 1070.94
R2 B.n24 B.t9 1070.94
R3 B.n32 B.t6 1070.94
R4 B.n273 B.n48 585
R5 B.n275 B.n274 585
R6 B.n276 B.n47 585
R7 B.n278 B.n277 585
R8 B.n279 B.n46 585
R9 B.n281 B.n280 585
R10 B.n282 B.n45 585
R11 B.n284 B.n283 585
R12 B.n285 B.n44 585
R13 B.n287 B.n286 585
R14 B.n288 B.n43 585
R15 B.n290 B.n289 585
R16 B.n291 B.n42 585
R17 B.n293 B.n292 585
R18 B.n294 B.n41 585
R19 B.n296 B.n295 585
R20 B.n297 B.n40 585
R21 B.n299 B.n298 585
R22 B.n300 B.n39 585
R23 B.n302 B.n301 585
R24 B.n303 B.n38 585
R25 B.n305 B.n304 585
R26 B.n306 B.n37 585
R27 B.n308 B.n307 585
R28 B.n309 B.n36 585
R29 B.n311 B.n310 585
R30 B.n312 B.n35 585
R31 B.n314 B.n313 585
R32 B.n315 B.n31 585
R33 B.n317 B.n316 585
R34 B.n318 B.n30 585
R35 B.n320 B.n319 585
R36 B.n321 B.n29 585
R37 B.n323 B.n322 585
R38 B.n324 B.n28 585
R39 B.n326 B.n325 585
R40 B.n327 B.n27 585
R41 B.n329 B.n328 585
R42 B.n330 B.n26 585
R43 B.n332 B.n331 585
R44 B.n334 B.n23 585
R45 B.n336 B.n335 585
R46 B.n337 B.n22 585
R47 B.n339 B.n338 585
R48 B.n340 B.n21 585
R49 B.n342 B.n341 585
R50 B.n343 B.n20 585
R51 B.n345 B.n344 585
R52 B.n346 B.n19 585
R53 B.n348 B.n347 585
R54 B.n349 B.n18 585
R55 B.n351 B.n350 585
R56 B.n352 B.n17 585
R57 B.n354 B.n353 585
R58 B.n355 B.n16 585
R59 B.n357 B.n356 585
R60 B.n358 B.n15 585
R61 B.n360 B.n359 585
R62 B.n361 B.n14 585
R63 B.n363 B.n362 585
R64 B.n364 B.n13 585
R65 B.n366 B.n365 585
R66 B.n367 B.n12 585
R67 B.n369 B.n368 585
R68 B.n370 B.n11 585
R69 B.n372 B.n371 585
R70 B.n373 B.n10 585
R71 B.n375 B.n374 585
R72 B.n376 B.n9 585
R73 B.n378 B.n377 585
R74 B.n272 B.n271 585
R75 B.n270 B.n49 585
R76 B.n269 B.n268 585
R77 B.n267 B.n50 585
R78 B.n266 B.n265 585
R79 B.n264 B.n51 585
R80 B.n263 B.n262 585
R81 B.n261 B.n52 585
R82 B.n260 B.n259 585
R83 B.n258 B.n53 585
R84 B.n257 B.n256 585
R85 B.n255 B.n54 585
R86 B.n254 B.n253 585
R87 B.n252 B.n55 585
R88 B.n251 B.n250 585
R89 B.n249 B.n56 585
R90 B.n248 B.n247 585
R91 B.n246 B.n57 585
R92 B.n245 B.n244 585
R93 B.n243 B.n58 585
R94 B.n242 B.n241 585
R95 B.n240 B.n59 585
R96 B.n239 B.n238 585
R97 B.n237 B.n60 585
R98 B.n236 B.n235 585
R99 B.n234 B.n61 585
R100 B.n233 B.n232 585
R101 B.n126 B.n101 585
R102 B.n128 B.n127 585
R103 B.n129 B.n100 585
R104 B.n131 B.n130 585
R105 B.n132 B.n99 585
R106 B.n134 B.n133 585
R107 B.n135 B.n98 585
R108 B.n137 B.n136 585
R109 B.n138 B.n97 585
R110 B.n140 B.n139 585
R111 B.n141 B.n96 585
R112 B.n143 B.n142 585
R113 B.n144 B.n95 585
R114 B.n146 B.n145 585
R115 B.n147 B.n94 585
R116 B.n149 B.n148 585
R117 B.n150 B.n93 585
R118 B.n152 B.n151 585
R119 B.n153 B.n92 585
R120 B.n155 B.n154 585
R121 B.n156 B.n91 585
R122 B.n158 B.n157 585
R123 B.n159 B.n90 585
R124 B.n161 B.n160 585
R125 B.n162 B.n89 585
R126 B.n164 B.n163 585
R127 B.n165 B.n88 585
R128 B.n167 B.n166 585
R129 B.n168 B.n87 585
R130 B.n170 B.n169 585
R131 B.n172 B.n84 585
R132 B.n174 B.n173 585
R133 B.n175 B.n83 585
R134 B.n177 B.n176 585
R135 B.n178 B.n82 585
R136 B.n180 B.n179 585
R137 B.n181 B.n81 585
R138 B.n183 B.n182 585
R139 B.n184 B.n80 585
R140 B.n186 B.n185 585
R141 B.n188 B.n187 585
R142 B.n189 B.n76 585
R143 B.n191 B.n190 585
R144 B.n192 B.n75 585
R145 B.n194 B.n193 585
R146 B.n195 B.n74 585
R147 B.n197 B.n196 585
R148 B.n198 B.n73 585
R149 B.n200 B.n199 585
R150 B.n201 B.n72 585
R151 B.n203 B.n202 585
R152 B.n204 B.n71 585
R153 B.n206 B.n205 585
R154 B.n207 B.n70 585
R155 B.n209 B.n208 585
R156 B.n210 B.n69 585
R157 B.n212 B.n211 585
R158 B.n213 B.n68 585
R159 B.n215 B.n214 585
R160 B.n216 B.n67 585
R161 B.n218 B.n217 585
R162 B.n219 B.n66 585
R163 B.n221 B.n220 585
R164 B.n222 B.n65 585
R165 B.n224 B.n223 585
R166 B.n225 B.n64 585
R167 B.n227 B.n226 585
R168 B.n228 B.n63 585
R169 B.n230 B.n229 585
R170 B.n231 B.n62 585
R171 B.n125 B.n124 585
R172 B.n123 B.n102 585
R173 B.n122 B.n121 585
R174 B.n120 B.n103 585
R175 B.n119 B.n118 585
R176 B.n117 B.n104 585
R177 B.n116 B.n115 585
R178 B.n114 B.n105 585
R179 B.n113 B.n112 585
R180 B.n111 B.n106 585
R181 B.n110 B.n109 585
R182 B.n108 B.n107 585
R183 B.n2 B.n0 585
R184 B.n397 B.n1 585
R185 B.n396 B.n395 585
R186 B.n394 B.n3 585
R187 B.n393 B.n392 585
R188 B.n391 B.n4 585
R189 B.n390 B.n389 585
R190 B.n388 B.n5 585
R191 B.n387 B.n386 585
R192 B.n385 B.n6 585
R193 B.n384 B.n383 585
R194 B.n382 B.n7 585
R195 B.n381 B.n380 585
R196 B.n379 B.n8 585
R197 B.n399 B.n398 585
R198 B.n126 B.n125 478.086
R199 B.n379 B.n378 478.086
R200 B.n233 B.n62 478.086
R201 B.n271 B.n48 478.086
R202 B.n77 B.t5 315.327
R203 B.n32 B.t7 315.327
R204 B.n85 B.t2 315.327
R205 B.n24 B.t10 315.327
R206 B.n78 B.t4 304.466
R207 B.n33 B.t8 304.466
R208 B.n86 B.t1 304.466
R209 B.n25 B.t11 304.466
R210 B.n125 B.n102 163.367
R211 B.n121 B.n102 163.367
R212 B.n121 B.n120 163.367
R213 B.n120 B.n119 163.367
R214 B.n119 B.n104 163.367
R215 B.n115 B.n104 163.367
R216 B.n115 B.n114 163.367
R217 B.n114 B.n113 163.367
R218 B.n113 B.n106 163.367
R219 B.n109 B.n106 163.367
R220 B.n109 B.n108 163.367
R221 B.n108 B.n2 163.367
R222 B.n398 B.n2 163.367
R223 B.n398 B.n397 163.367
R224 B.n397 B.n396 163.367
R225 B.n396 B.n3 163.367
R226 B.n392 B.n3 163.367
R227 B.n392 B.n391 163.367
R228 B.n391 B.n390 163.367
R229 B.n390 B.n5 163.367
R230 B.n386 B.n5 163.367
R231 B.n386 B.n385 163.367
R232 B.n385 B.n384 163.367
R233 B.n384 B.n7 163.367
R234 B.n380 B.n7 163.367
R235 B.n380 B.n379 163.367
R236 B.n127 B.n126 163.367
R237 B.n127 B.n100 163.367
R238 B.n131 B.n100 163.367
R239 B.n132 B.n131 163.367
R240 B.n133 B.n132 163.367
R241 B.n133 B.n98 163.367
R242 B.n137 B.n98 163.367
R243 B.n138 B.n137 163.367
R244 B.n139 B.n138 163.367
R245 B.n139 B.n96 163.367
R246 B.n143 B.n96 163.367
R247 B.n144 B.n143 163.367
R248 B.n145 B.n144 163.367
R249 B.n145 B.n94 163.367
R250 B.n149 B.n94 163.367
R251 B.n150 B.n149 163.367
R252 B.n151 B.n150 163.367
R253 B.n151 B.n92 163.367
R254 B.n155 B.n92 163.367
R255 B.n156 B.n155 163.367
R256 B.n157 B.n156 163.367
R257 B.n157 B.n90 163.367
R258 B.n161 B.n90 163.367
R259 B.n162 B.n161 163.367
R260 B.n163 B.n162 163.367
R261 B.n163 B.n88 163.367
R262 B.n167 B.n88 163.367
R263 B.n168 B.n167 163.367
R264 B.n169 B.n168 163.367
R265 B.n169 B.n84 163.367
R266 B.n174 B.n84 163.367
R267 B.n175 B.n174 163.367
R268 B.n176 B.n175 163.367
R269 B.n176 B.n82 163.367
R270 B.n180 B.n82 163.367
R271 B.n181 B.n180 163.367
R272 B.n182 B.n181 163.367
R273 B.n182 B.n80 163.367
R274 B.n186 B.n80 163.367
R275 B.n187 B.n186 163.367
R276 B.n187 B.n76 163.367
R277 B.n191 B.n76 163.367
R278 B.n192 B.n191 163.367
R279 B.n193 B.n192 163.367
R280 B.n193 B.n74 163.367
R281 B.n197 B.n74 163.367
R282 B.n198 B.n197 163.367
R283 B.n199 B.n198 163.367
R284 B.n199 B.n72 163.367
R285 B.n203 B.n72 163.367
R286 B.n204 B.n203 163.367
R287 B.n205 B.n204 163.367
R288 B.n205 B.n70 163.367
R289 B.n209 B.n70 163.367
R290 B.n210 B.n209 163.367
R291 B.n211 B.n210 163.367
R292 B.n211 B.n68 163.367
R293 B.n215 B.n68 163.367
R294 B.n216 B.n215 163.367
R295 B.n217 B.n216 163.367
R296 B.n217 B.n66 163.367
R297 B.n221 B.n66 163.367
R298 B.n222 B.n221 163.367
R299 B.n223 B.n222 163.367
R300 B.n223 B.n64 163.367
R301 B.n227 B.n64 163.367
R302 B.n228 B.n227 163.367
R303 B.n229 B.n228 163.367
R304 B.n229 B.n62 163.367
R305 B.n234 B.n233 163.367
R306 B.n235 B.n234 163.367
R307 B.n235 B.n60 163.367
R308 B.n239 B.n60 163.367
R309 B.n240 B.n239 163.367
R310 B.n241 B.n240 163.367
R311 B.n241 B.n58 163.367
R312 B.n245 B.n58 163.367
R313 B.n246 B.n245 163.367
R314 B.n247 B.n246 163.367
R315 B.n247 B.n56 163.367
R316 B.n251 B.n56 163.367
R317 B.n252 B.n251 163.367
R318 B.n253 B.n252 163.367
R319 B.n253 B.n54 163.367
R320 B.n257 B.n54 163.367
R321 B.n258 B.n257 163.367
R322 B.n259 B.n258 163.367
R323 B.n259 B.n52 163.367
R324 B.n263 B.n52 163.367
R325 B.n264 B.n263 163.367
R326 B.n265 B.n264 163.367
R327 B.n265 B.n50 163.367
R328 B.n269 B.n50 163.367
R329 B.n270 B.n269 163.367
R330 B.n271 B.n270 163.367
R331 B.n378 B.n9 163.367
R332 B.n374 B.n9 163.367
R333 B.n374 B.n373 163.367
R334 B.n373 B.n372 163.367
R335 B.n372 B.n11 163.367
R336 B.n368 B.n11 163.367
R337 B.n368 B.n367 163.367
R338 B.n367 B.n366 163.367
R339 B.n366 B.n13 163.367
R340 B.n362 B.n13 163.367
R341 B.n362 B.n361 163.367
R342 B.n361 B.n360 163.367
R343 B.n360 B.n15 163.367
R344 B.n356 B.n15 163.367
R345 B.n356 B.n355 163.367
R346 B.n355 B.n354 163.367
R347 B.n354 B.n17 163.367
R348 B.n350 B.n17 163.367
R349 B.n350 B.n349 163.367
R350 B.n349 B.n348 163.367
R351 B.n348 B.n19 163.367
R352 B.n344 B.n19 163.367
R353 B.n344 B.n343 163.367
R354 B.n343 B.n342 163.367
R355 B.n342 B.n21 163.367
R356 B.n338 B.n21 163.367
R357 B.n338 B.n337 163.367
R358 B.n337 B.n336 163.367
R359 B.n336 B.n23 163.367
R360 B.n331 B.n23 163.367
R361 B.n331 B.n330 163.367
R362 B.n330 B.n329 163.367
R363 B.n329 B.n27 163.367
R364 B.n325 B.n27 163.367
R365 B.n325 B.n324 163.367
R366 B.n324 B.n323 163.367
R367 B.n323 B.n29 163.367
R368 B.n319 B.n29 163.367
R369 B.n319 B.n318 163.367
R370 B.n318 B.n317 163.367
R371 B.n317 B.n31 163.367
R372 B.n313 B.n31 163.367
R373 B.n313 B.n312 163.367
R374 B.n312 B.n311 163.367
R375 B.n311 B.n36 163.367
R376 B.n307 B.n36 163.367
R377 B.n307 B.n306 163.367
R378 B.n306 B.n305 163.367
R379 B.n305 B.n38 163.367
R380 B.n301 B.n38 163.367
R381 B.n301 B.n300 163.367
R382 B.n300 B.n299 163.367
R383 B.n299 B.n40 163.367
R384 B.n295 B.n40 163.367
R385 B.n295 B.n294 163.367
R386 B.n294 B.n293 163.367
R387 B.n293 B.n42 163.367
R388 B.n289 B.n42 163.367
R389 B.n289 B.n288 163.367
R390 B.n288 B.n287 163.367
R391 B.n287 B.n44 163.367
R392 B.n283 B.n44 163.367
R393 B.n283 B.n282 163.367
R394 B.n282 B.n281 163.367
R395 B.n281 B.n46 163.367
R396 B.n277 B.n46 163.367
R397 B.n277 B.n276 163.367
R398 B.n276 B.n275 163.367
R399 B.n275 B.n48 163.367
R400 B.n79 B.n78 59.5399
R401 B.n171 B.n86 59.5399
R402 B.n333 B.n25 59.5399
R403 B.n34 B.n33 59.5399
R404 B.n377 B.n8 31.0639
R405 B.n273 B.n272 31.0639
R406 B.n232 B.n231 31.0639
R407 B.n124 B.n101 31.0639
R408 B B.n399 18.0485
R409 B.n78 B.n77 10.8611
R410 B.n86 B.n85 10.8611
R411 B.n25 B.n24 10.8611
R412 B.n33 B.n32 10.8611
R413 B.n377 B.n376 10.6151
R414 B.n376 B.n375 10.6151
R415 B.n375 B.n10 10.6151
R416 B.n371 B.n10 10.6151
R417 B.n371 B.n370 10.6151
R418 B.n370 B.n369 10.6151
R419 B.n369 B.n12 10.6151
R420 B.n365 B.n12 10.6151
R421 B.n365 B.n364 10.6151
R422 B.n364 B.n363 10.6151
R423 B.n363 B.n14 10.6151
R424 B.n359 B.n14 10.6151
R425 B.n359 B.n358 10.6151
R426 B.n358 B.n357 10.6151
R427 B.n357 B.n16 10.6151
R428 B.n353 B.n16 10.6151
R429 B.n353 B.n352 10.6151
R430 B.n352 B.n351 10.6151
R431 B.n351 B.n18 10.6151
R432 B.n347 B.n18 10.6151
R433 B.n347 B.n346 10.6151
R434 B.n346 B.n345 10.6151
R435 B.n345 B.n20 10.6151
R436 B.n341 B.n20 10.6151
R437 B.n341 B.n340 10.6151
R438 B.n340 B.n339 10.6151
R439 B.n339 B.n22 10.6151
R440 B.n335 B.n22 10.6151
R441 B.n335 B.n334 10.6151
R442 B.n332 B.n26 10.6151
R443 B.n328 B.n26 10.6151
R444 B.n328 B.n327 10.6151
R445 B.n327 B.n326 10.6151
R446 B.n326 B.n28 10.6151
R447 B.n322 B.n28 10.6151
R448 B.n322 B.n321 10.6151
R449 B.n321 B.n320 10.6151
R450 B.n320 B.n30 10.6151
R451 B.n316 B.n315 10.6151
R452 B.n315 B.n314 10.6151
R453 B.n314 B.n35 10.6151
R454 B.n310 B.n35 10.6151
R455 B.n310 B.n309 10.6151
R456 B.n309 B.n308 10.6151
R457 B.n308 B.n37 10.6151
R458 B.n304 B.n37 10.6151
R459 B.n304 B.n303 10.6151
R460 B.n303 B.n302 10.6151
R461 B.n302 B.n39 10.6151
R462 B.n298 B.n39 10.6151
R463 B.n298 B.n297 10.6151
R464 B.n297 B.n296 10.6151
R465 B.n296 B.n41 10.6151
R466 B.n292 B.n41 10.6151
R467 B.n292 B.n291 10.6151
R468 B.n291 B.n290 10.6151
R469 B.n290 B.n43 10.6151
R470 B.n286 B.n43 10.6151
R471 B.n286 B.n285 10.6151
R472 B.n285 B.n284 10.6151
R473 B.n284 B.n45 10.6151
R474 B.n280 B.n45 10.6151
R475 B.n280 B.n279 10.6151
R476 B.n279 B.n278 10.6151
R477 B.n278 B.n47 10.6151
R478 B.n274 B.n47 10.6151
R479 B.n274 B.n273 10.6151
R480 B.n232 B.n61 10.6151
R481 B.n236 B.n61 10.6151
R482 B.n237 B.n236 10.6151
R483 B.n238 B.n237 10.6151
R484 B.n238 B.n59 10.6151
R485 B.n242 B.n59 10.6151
R486 B.n243 B.n242 10.6151
R487 B.n244 B.n243 10.6151
R488 B.n244 B.n57 10.6151
R489 B.n248 B.n57 10.6151
R490 B.n249 B.n248 10.6151
R491 B.n250 B.n249 10.6151
R492 B.n250 B.n55 10.6151
R493 B.n254 B.n55 10.6151
R494 B.n255 B.n254 10.6151
R495 B.n256 B.n255 10.6151
R496 B.n256 B.n53 10.6151
R497 B.n260 B.n53 10.6151
R498 B.n261 B.n260 10.6151
R499 B.n262 B.n261 10.6151
R500 B.n262 B.n51 10.6151
R501 B.n266 B.n51 10.6151
R502 B.n267 B.n266 10.6151
R503 B.n268 B.n267 10.6151
R504 B.n268 B.n49 10.6151
R505 B.n272 B.n49 10.6151
R506 B.n128 B.n101 10.6151
R507 B.n129 B.n128 10.6151
R508 B.n130 B.n129 10.6151
R509 B.n130 B.n99 10.6151
R510 B.n134 B.n99 10.6151
R511 B.n135 B.n134 10.6151
R512 B.n136 B.n135 10.6151
R513 B.n136 B.n97 10.6151
R514 B.n140 B.n97 10.6151
R515 B.n141 B.n140 10.6151
R516 B.n142 B.n141 10.6151
R517 B.n142 B.n95 10.6151
R518 B.n146 B.n95 10.6151
R519 B.n147 B.n146 10.6151
R520 B.n148 B.n147 10.6151
R521 B.n148 B.n93 10.6151
R522 B.n152 B.n93 10.6151
R523 B.n153 B.n152 10.6151
R524 B.n154 B.n153 10.6151
R525 B.n154 B.n91 10.6151
R526 B.n158 B.n91 10.6151
R527 B.n159 B.n158 10.6151
R528 B.n160 B.n159 10.6151
R529 B.n160 B.n89 10.6151
R530 B.n164 B.n89 10.6151
R531 B.n165 B.n164 10.6151
R532 B.n166 B.n165 10.6151
R533 B.n166 B.n87 10.6151
R534 B.n170 B.n87 10.6151
R535 B.n173 B.n172 10.6151
R536 B.n173 B.n83 10.6151
R537 B.n177 B.n83 10.6151
R538 B.n178 B.n177 10.6151
R539 B.n179 B.n178 10.6151
R540 B.n179 B.n81 10.6151
R541 B.n183 B.n81 10.6151
R542 B.n184 B.n183 10.6151
R543 B.n185 B.n184 10.6151
R544 B.n189 B.n188 10.6151
R545 B.n190 B.n189 10.6151
R546 B.n190 B.n75 10.6151
R547 B.n194 B.n75 10.6151
R548 B.n195 B.n194 10.6151
R549 B.n196 B.n195 10.6151
R550 B.n196 B.n73 10.6151
R551 B.n200 B.n73 10.6151
R552 B.n201 B.n200 10.6151
R553 B.n202 B.n201 10.6151
R554 B.n202 B.n71 10.6151
R555 B.n206 B.n71 10.6151
R556 B.n207 B.n206 10.6151
R557 B.n208 B.n207 10.6151
R558 B.n208 B.n69 10.6151
R559 B.n212 B.n69 10.6151
R560 B.n213 B.n212 10.6151
R561 B.n214 B.n213 10.6151
R562 B.n214 B.n67 10.6151
R563 B.n218 B.n67 10.6151
R564 B.n219 B.n218 10.6151
R565 B.n220 B.n219 10.6151
R566 B.n220 B.n65 10.6151
R567 B.n224 B.n65 10.6151
R568 B.n225 B.n224 10.6151
R569 B.n226 B.n225 10.6151
R570 B.n226 B.n63 10.6151
R571 B.n230 B.n63 10.6151
R572 B.n231 B.n230 10.6151
R573 B.n124 B.n123 10.6151
R574 B.n123 B.n122 10.6151
R575 B.n122 B.n103 10.6151
R576 B.n118 B.n103 10.6151
R577 B.n118 B.n117 10.6151
R578 B.n117 B.n116 10.6151
R579 B.n116 B.n105 10.6151
R580 B.n112 B.n105 10.6151
R581 B.n112 B.n111 10.6151
R582 B.n111 B.n110 10.6151
R583 B.n110 B.n107 10.6151
R584 B.n107 B.n0 10.6151
R585 B.n395 B.n1 10.6151
R586 B.n395 B.n394 10.6151
R587 B.n394 B.n393 10.6151
R588 B.n393 B.n4 10.6151
R589 B.n389 B.n4 10.6151
R590 B.n389 B.n388 10.6151
R591 B.n388 B.n387 10.6151
R592 B.n387 B.n6 10.6151
R593 B.n383 B.n6 10.6151
R594 B.n383 B.n382 10.6151
R595 B.n382 B.n381 10.6151
R596 B.n381 B.n8 10.6151
R597 B.n334 B.n333 8.74196
R598 B.n316 B.n34 8.74196
R599 B.n171 B.n170 8.74196
R600 B.n188 B.n79 8.74196
R601 B.n399 B.n0 2.81026
R602 B.n399 B.n1 2.81026
R603 B.n333 B.n332 1.87367
R604 B.n34 B.n30 1.87367
R605 B.n172 B.n171 1.87367
R606 B.n185 B.n79 1.87367
R607 VP.n1 VP.t0 1019.57
R608 VP.n1 VP.t1 1019.57
R609 VP.n0 VP.t3 1019.57
R610 VP.n0 VP.t2 1019.57
R611 VP.n2 VP.n0 197.323
R612 VP.n2 VP.n1 161.3
R613 VP VP.n2 0.0516364
R614 VTAIL.n330 VTAIL.n294 756.745
R615 VTAIL.n36 VTAIL.n0 756.745
R616 VTAIL.n78 VTAIL.n42 756.745
R617 VTAIL.n120 VTAIL.n84 756.745
R618 VTAIL.n288 VTAIL.n252 756.745
R619 VTAIL.n246 VTAIL.n210 756.745
R620 VTAIL.n204 VTAIL.n168 756.745
R621 VTAIL.n162 VTAIL.n126 756.745
R622 VTAIL.n306 VTAIL.n305 585
R623 VTAIL.n311 VTAIL.n310 585
R624 VTAIL.n313 VTAIL.n312 585
R625 VTAIL.n302 VTAIL.n301 585
R626 VTAIL.n319 VTAIL.n318 585
R627 VTAIL.n321 VTAIL.n320 585
R628 VTAIL.n298 VTAIL.n297 585
R629 VTAIL.n328 VTAIL.n327 585
R630 VTAIL.n329 VTAIL.n296 585
R631 VTAIL.n331 VTAIL.n330 585
R632 VTAIL.n12 VTAIL.n11 585
R633 VTAIL.n17 VTAIL.n16 585
R634 VTAIL.n19 VTAIL.n18 585
R635 VTAIL.n8 VTAIL.n7 585
R636 VTAIL.n25 VTAIL.n24 585
R637 VTAIL.n27 VTAIL.n26 585
R638 VTAIL.n4 VTAIL.n3 585
R639 VTAIL.n34 VTAIL.n33 585
R640 VTAIL.n35 VTAIL.n2 585
R641 VTAIL.n37 VTAIL.n36 585
R642 VTAIL.n54 VTAIL.n53 585
R643 VTAIL.n59 VTAIL.n58 585
R644 VTAIL.n61 VTAIL.n60 585
R645 VTAIL.n50 VTAIL.n49 585
R646 VTAIL.n67 VTAIL.n66 585
R647 VTAIL.n69 VTAIL.n68 585
R648 VTAIL.n46 VTAIL.n45 585
R649 VTAIL.n76 VTAIL.n75 585
R650 VTAIL.n77 VTAIL.n44 585
R651 VTAIL.n79 VTAIL.n78 585
R652 VTAIL.n96 VTAIL.n95 585
R653 VTAIL.n101 VTAIL.n100 585
R654 VTAIL.n103 VTAIL.n102 585
R655 VTAIL.n92 VTAIL.n91 585
R656 VTAIL.n109 VTAIL.n108 585
R657 VTAIL.n111 VTAIL.n110 585
R658 VTAIL.n88 VTAIL.n87 585
R659 VTAIL.n118 VTAIL.n117 585
R660 VTAIL.n119 VTAIL.n86 585
R661 VTAIL.n121 VTAIL.n120 585
R662 VTAIL.n289 VTAIL.n288 585
R663 VTAIL.n287 VTAIL.n254 585
R664 VTAIL.n286 VTAIL.n285 585
R665 VTAIL.n257 VTAIL.n255 585
R666 VTAIL.n280 VTAIL.n279 585
R667 VTAIL.n278 VTAIL.n277 585
R668 VTAIL.n261 VTAIL.n260 585
R669 VTAIL.n272 VTAIL.n271 585
R670 VTAIL.n270 VTAIL.n269 585
R671 VTAIL.n265 VTAIL.n264 585
R672 VTAIL.n247 VTAIL.n246 585
R673 VTAIL.n245 VTAIL.n212 585
R674 VTAIL.n244 VTAIL.n243 585
R675 VTAIL.n215 VTAIL.n213 585
R676 VTAIL.n238 VTAIL.n237 585
R677 VTAIL.n236 VTAIL.n235 585
R678 VTAIL.n219 VTAIL.n218 585
R679 VTAIL.n230 VTAIL.n229 585
R680 VTAIL.n228 VTAIL.n227 585
R681 VTAIL.n223 VTAIL.n222 585
R682 VTAIL.n205 VTAIL.n204 585
R683 VTAIL.n203 VTAIL.n170 585
R684 VTAIL.n202 VTAIL.n201 585
R685 VTAIL.n173 VTAIL.n171 585
R686 VTAIL.n196 VTAIL.n195 585
R687 VTAIL.n194 VTAIL.n193 585
R688 VTAIL.n177 VTAIL.n176 585
R689 VTAIL.n188 VTAIL.n187 585
R690 VTAIL.n186 VTAIL.n185 585
R691 VTAIL.n181 VTAIL.n180 585
R692 VTAIL.n163 VTAIL.n162 585
R693 VTAIL.n161 VTAIL.n128 585
R694 VTAIL.n160 VTAIL.n159 585
R695 VTAIL.n131 VTAIL.n129 585
R696 VTAIL.n154 VTAIL.n153 585
R697 VTAIL.n152 VTAIL.n151 585
R698 VTAIL.n135 VTAIL.n134 585
R699 VTAIL.n146 VTAIL.n145 585
R700 VTAIL.n144 VTAIL.n143 585
R701 VTAIL.n139 VTAIL.n138 585
R702 VTAIL.n307 VTAIL.t0 329.043
R703 VTAIL.n13 VTAIL.t2 329.043
R704 VTAIL.n55 VTAIL.t6 329.043
R705 VTAIL.n97 VTAIL.t4 329.043
R706 VTAIL.n266 VTAIL.t5 329.043
R707 VTAIL.n224 VTAIL.t7 329.043
R708 VTAIL.n182 VTAIL.t1 329.043
R709 VTAIL.n140 VTAIL.t3 329.043
R710 VTAIL.n311 VTAIL.n305 171.744
R711 VTAIL.n312 VTAIL.n311 171.744
R712 VTAIL.n312 VTAIL.n301 171.744
R713 VTAIL.n319 VTAIL.n301 171.744
R714 VTAIL.n320 VTAIL.n319 171.744
R715 VTAIL.n320 VTAIL.n297 171.744
R716 VTAIL.n328 VTAIL.n297 171.744
R717 VTAIL.n329 VTAIL.n328 171.744
R718 VTAIL.n330 VTAIL.n329 171.744
R719 VTAIL.n17 VTAIL.n11 171.744
R720 VTAIL.n18 VTAIL.n17 171.744
R721 VTAIL.n18 VTAIL.n7 171.744
R722 VTAIL.n25 VTAIL.n7 171.744
R723 VTAIL.n26 VTAIL.n25 171.744
R724 VTAIL.n26 VTAIL.n3 171.744
R725 VTAIL.n34 VTAIL.n3 171.744
R726 VTAIL.n35 VTAIL.n34 171.744
R727 VTAIL.n36 VTAIL.n35 171.744
R728 VTAIL.n59 VTAIL.n53 171.744
R729 VTAIL.n60 VTAIL.n59 171.744
R730 VTAIL.n60 VTAIL.n49 171.744
R731 VTAIL.n67 VTAIL.n49 171.744
R732 VTAIL.n68 VTAIL.n67 171.744
R733 VTAIL.n68 VTAIL.n45 171.744
R734 VTAIL.n76 VTAIL.n45 171.744
R735 VTAIL.n77 VTAIL.n76 171.744
R736 VTAIL.n78 VTAIL.n77 171.744
R737 VTAIL.n101 VTAIL.n95 171.744
R738 VTAIL.n102 VTAIL.n101 171.744
R739 VTAIL.n102 VTAIL.n91 171.744
R740 VTAIL.n109 VTAIL.n91 171.744
R741 VTAIL.n110 VTAIL.n109 171.744
R742 VTAIL.n110 VTAIL.n87 171.744
R743 VTAIL.n118 VTAIL.n87 171.744
R744 VTAIL.n119 VTAIL.n118 171.744
R745 VTAIL.n120 VTAIL.n119 171.744
R746 VTAIL.n288 VTAIL.n287 171.744
R747 VTAIL.n287 VTAIL.n286 171.744
R748 VTAIL.n286 VTAIL.n255 171.744
R749 VTAIL.n279 VTAIL.n255 171.744
R750 VTAIL.n279 VTAIL.n278 171.744
R751 VTAIL.n278 VTAIL.n260 171.744
R752 VTAIL.n271 VTAIL.n260 171.744
R753 VTAIL.n271 VTAIL.n270 171.744
R754 VTAIL.n270 VTAIL.n264 171.744
R755 VTAIL.n246 VTAIL.n245 171.744
R756 VTAIL.n245 VTAIL.n244 171.744
R757 VTAIL.n244 VTAIL.n213 171.744
R758 VTAIL.n237 VTAIL.n213 171.744
R759 VTAIL.n237 VTAIL.n236 171.744
R760 VTAIL.n236 VTAIL.n218 171.744
R761 VTAIL.n229 VTAIL.n218 171.744
R762 VTAIL.n229 VTAIL.n228 171.744
R763 VTAIL.n228 VTAIL.n222 171.744
R764 VTAIL.n204 VTAIL.n203 171.744
R765 VTAIL.n203 VTAIL.n202 171.744
R766 VTAIL.n202 VTAIL.n171 171.744
R767 VTAIL.n195 VTAIL.n171 171.744
R768 VTAIL.n195 VTAIL.n194 171.744
R769 VTAIL.n194 VTAIL.n176 171.744
R770 VTAIL.n187 VTAIL.n176 171.744
R771 VTAIL.n187 VTAIL.n186 171.744
R772 VTAIL.n186 VTAIL.n180 171.744
R773 VTAIL.n162 VTAIL.n161 171.744
R774 VTAIL.n161 VTAIL.n160 171.744
R775 VTAIL.n160 VTAIL.n129 171.744
R776 VTAIL.n153 VTAIL.n129 171.744
R777 VTAIL.n153 VTAIL.n152 171.744
R778 VTAIL.n152 VTAIL.n134 171.744
R779 VTAIL.n145 VTAIL.n134 171.744
R780 VTAIL.n145 VTAIL.n144 171.744
R781 VTAIL.n144 VTAIL.n138 171.744
R782 VTAIL.t0 VTAIL.n305 85.8723
R783 VTAIL.t2 VTAIL.n11 85.8723
R784 VTAIL.t6 VTAIL.n53 85.8723
R785 VTAIL.t4 VTAIL.n95 85.8723
R786 VTAIL.t5 VTAIL.n264 85.8723
R787 VTAIL.t7 VTAIL.n222 85.8723
R788 VTAIL.t1 VTAIL.n180 85.8723
R789 VTAIL.t3 VTAIL.n138 85.8723
R790 VTAIL.n335 VTAIL.n334 36.8399
R791 VTAIL.n41 VTAIL.n40 36.8399
R792 VTAIL.n83 VTAIL.n82 36.8399
R793 VTAIL.n125 VTAIL.n124 36.8399
R794 VTAIL.n293 VTAIL.n292 36.8399
R795 VTAIL.n251 VTAIL.n250 36.8399
R796 VTAIL.n209 VTAIL.n208 36.8399
R797 VTAIL.n167 VTAIL.n166 36.8399
R798 VTAIL.n335 VTAIL.n293 19.7979
R799 VTAIL.n167 VTAIL.n125 19.7979
R800 VTAIL.n331 VTAIL.n296 13.1884
R801 VTAIL.n37 VTAIL.n2 13.1884
R802 VTAIL.n79 VTAIL.n44 13.1884
R803 VTAIL.n121 VTAIL.n86 13.1884
R804 VTAIL.n289 VTAIL.n254 13.1884
R805 VTAIL.n247 VTAIL.n212 13.1884
R806 VTAIL.n205 VTAIL.n170 13.1884
R807 VTAIL.n163 VTAIL.n128 13.1884
R808 VTAIL.n327 VTAIL.n326 12.8005
R809 VTAIL.n332 VTAIL.n294 12.8005
R810 VTAIL.n33 VTAIL.n32 12.8005
R811 VTAIL.n38 VTAIL.n0 12.8005
R812 VTAIL.n75 VTAIL.n74 12.8005
R813 VTAIL.n80 VTAIL.n42 12.8005
R814 VTAIL.n117 VTAIL.n116 12.8005
R815 VTAIL.n122 VTAIL.n84 12.8005
R816 VTAIL.n290 VTAIL.n252 12.8005
R817 VTAIL.n285 VTAIL.n256 12.8005
R818 VTAIL.n248 VTAIL.n210 12.8005
R819 VTAIL.n243 VTAIL.n214 12.8005
R820 VTAIL.n206 VTAIL.n168 12.8005
R821 VTAIL.n201 VTAIL.n172 12.8005
R822 VTAIL.n164 VTAIL.n126 12.8005
R823 VTAIL.n159 VTAIL.n130 12.8005
R824 VTAIL.n325 VTAIL.n298 12.0247
R825 VTAIL.n31 VTAIL.n4 12.0247
R826 VTAIL.n73 VTAIL.n46 12.0247
R827 VTAIL.n115 VTAIL.n88 12.0247
R828 VTAIL.n284 VTAIL.n257 12.0247
R829 VTAIL.n242 VTAIL.n215 12.0247
R830 VTAIL.n200 VTAIL.n173 12.0247
R831 VTAIL.n158 VTAIL.n131 12.0247
R832 VTAIL.n322 VTAIL.n321 11.249
R833 VTAIL.n28 VTAIL.n27 11.249
R834 VTAIL.n70 VTAIL.n69 11.249
R835 VTAIL.n112 VTAIL.n111 11.249
R836 VTAIL.n281 VTAIL.n280 11.249
R837 VTAIL.n239 VTAIL.n238 11.249
R838 VTAIL.n197 VTAIL.n196 11.249
R839 VTAIL.n155 VTAIL.n154 11.249
R840 VTAIL.n307 VTAIL.n306 10.7238
R841 VTAIL.n13 VTAIL.n12 10.7238
R842 VTAIL.n55 VTAIL.n54 10.7238
R843 VTAIL.n97 VTAIL.n96 10.7238
R844 VTAIL.n266 VTAIL.n265 10.7238
R845 VTAIL.n224 VTAIL.n223 10.7238
R846 VTAIL.n182 VTAIL.n181 10.7238
R847 VTAIL.n140 VTAIL.n139 10.7238
R848 VTAIL.n318 VTAIL.n300 10.4732
R849 VTAIL.n24 VTAIL.n6 10.4732
R850 VTAIL.n66 VTAIL.n48 10.4732
R851 VTAIL.n108 VTAIL.n90 10.4732
R852 VTAIL.n277 VTAIL.n259 10.4732
R853 VTAIL.n235 VTAIL.n217 10.4732
R854 VTAIL.n193 VTAIL.n175 10.4732
R855 VTAIL.n151 VTAIL.n133 10.4732
R856 VTAIL.n317 VTAIL.n302 9.69747
R857 VTAIL.n23 VTAIL.n8 9.69747
R858 VTAIL.n65 VTAIL.n50 9.69747
R859 VTAIL.n107 VTAIL.n92 9.69747
R860 VTAIL.n276 VTAIL.n261 9.69747
R861 VTAIL.n234 VTAIL.n219 9.69747
R862 VTAIL.n192 VTAIL.n177 9.69747
R863 VTAIL.n150 VTAIL.n135 9.69747
R864 VTAIL.n334 VTAIL.n333 9.45567
R865 VTAIL.n40 VTAIL.n39 9.45567
R866 VTAIL.n82 VTAIL.n81 9.45567
R867 VTAIL.n124 VTAIL.n123 9.45567
R868 VTAIL.n292 VTAIL.n291 9.45567
R869 VTAIL.n250 VTAIL.n249 9.45567
R870 VTAIL.n208 VTAIL.n207 9.45567
R871 VTAIL.n166 VTAIL.n165 9.45567
R872 VTAIL.n333 VTAIL.n332 9.3005
R873 VTAIL.n309 VTAIL.n308 9.3005
R874 VTAIL.n304 VTAIL.n303 9.3005
R875 VTAIL.n315 VTAIL.n314 9.3005
R876 VTAIL.n317 VTAIL.n316 9.3005
R877 VTAIL.n300 VTAIL.n299 9.3005
R878 VTAIL.n323 VTAIL.n322 9.3005
R879 VTAIL.n325 VTAIL.n324 9.3005
R880 VTAIL.n326 VTAIL.n295 9.3005
R881 VTAIL.n39 VTAIL.n38 9.3005
R882 VTAIL.n15 VTAIL.n14 9.3005
R883 VTAIL.n10 VTAIL.n9 9.3005
R884 VTAIL.n21 VTAIL.n20 9.3005
R885 VTAIL.n23 VTAIL.n22 9.3005
R886 VTAIL.n6 VTAIL.n5 9.3005
R887 VTAIL.n29 VTAIL.n28 9.3005
R888 VTAIL.n31 VTAIL.n30 9.3005
R889 VTAIL.n32 VTAIL.n1 9.3005
R890 VTAIL.n81 VTAIL.n80 9.3005
R891 VTAIL.n57 VTAIL.n56 9.3005
R892 VTAIL.n52 VTAIL.n51 9.3005
R893 VTAIL.n63 VTAIL.n62 9.3005
R894 VTAIL.n65 VTAIL.n64 9.3005
R895 VTAIL.n48 VTAIL.n47 9.3005
R896 VTAIL.n71 VTAIL.n70 9.3005
R897 VTAIL.n73 VTAIL.n72 9.3005
R898 VTAIL.n74 VTAIL.n43 9.3005
R899 VTAIL.n123 VTAIL.n122 9.3005
R900 VTAIL.n99 VTAIL.n98 9.3005
R901 VTAIL.n94 VTAIL.n93 9.3005
R902 VTAIL.n105 VTAIL.n104 9.3005
R903 VTAIL.n107 VTAIL.n106 9.3005
R904 VTAIL.n90 VTAIL.n89 9.3005
R905 VTAIL.n113 VTAIL.n112 9.3005
R906 VTAIL.n115 VTAIL.n114 9.3005
R907 VTAIL.n116 VTAIL.n85 9.3005
R908 VTAIL.n268 VTAIL.n267 9.3005
R909 VTAIL.n263 VTAIL.n262 9.3005
R910 VTAIL.n274 VTAIL.n273 9.3005
R911 VTAIL.n276 VTAIL.n275 9.3005
R912 VTAIL.n259 VTAIL.n258 9.3005
R913 VTAIL.n282 VTAIL.n281 9.3005
R914 VTAIL.n284 VTAIL.n283 9.3005
R915 VTAIL.n256 VTAIL.n253 9.3005
R916 VTAIL.n291 VTAIL.n290 9.3005
R917 VTAIL.n226 VTAIL.n225 9.3005
R918 VTAIL.n221 VTAIL.n220 9.3005
R919 VTAIL.n232 VTAIL.n231 9.3005
R920 VTAIL.n234 VTAIL.n233 9.3005
R921 VTAIL.n217 VTAIL.n216 9.3005
R922 VTAIL.n240 VTAIL.n239 9.3005
R923 VTAIL.n242 VTAIL.n241 9.3005
R924 VTAIL.n214 VTAIL.n211 9.3005
R925 VTAIL.n249 VTAIL.n248 9.3005
R926 VTAIL.n184 VTAIL.n183 9.3005
R927 VTAIL.n179 VTAIL.n178 9.3005
R928 VTAIL.n190 VTAIL.n189 9.3005
R929 VTAIL.n192 VTAIL.n191 9.3005
R930 VTAIL.n175 VTAIL.n174 9.3005
R931 VTAIL.n198 VTAIL.n197 9.3005
R932 VTAIL.n200 VTAIL.n199 9.3005
R933 VTAIL.n172 VTAIL.n169 9.3005
R934 VTAIL.n207 VTAIL.n206 9.3005
R935 VTAIL.n142 VTAIL.n141 9.3005
R936 VTAIL.n137 VTAIL.n136 9.3005
R937 VTAIL.n148 VTAIL.n147 9.3005
R938 VTAIL.n150 VTAIL.n149 9.3005
R939 VTAIL.n133 VTAIL.n132 9.3005
R940 VTAIL.n156 VTAIL.n155 9.3005
R941 VTAIL.n158 VTAIL.n157 9.3005
R942 VTAIL.n130 VTAIL.n127 9.3005
R943 VTAIL.n165 VTAIL.n164 9.3005
R944 VTAIL.n314 VTAIL.n313 8.92171
R945 VTAIL.n20 VTAIL.n19 8.92171
R946 VTAIL.n62 VTAIL.n61 8.92171
R947 VTAIL.n104 VTAIL.n103 8.92171
R948 VTAIL.n273 VTAIL.n272 8.92171
R949 VTAIL.n231 VTAIL.n230 8.92171
R950 VTAIL.n189 VTAIL.n188 8.92171
R951 VTAIL.n147 VTAIL.n146 8.92171
R952 VTAIL.n310 VTAIL.n304 8.14595
R953 VTAIL.n16 VTAIL.n10 8.14595
R954 VTAIL.n58 VTAIL.n52 8.14595
R955 VTAIL.n100 VTAIL.n94 8.14595
R956 VTAIL.n269 VTAIL.n263 8.14595
R957 VTAIL.n227 VTAIL.n221 8.14595
R958 VTAIL.n185 VTAIL.n179 8.14595
R959 VTAIL.n143 VTAIL.n137 8.14595
R960 VTAIL.n309 VTAIL.n306 7.3702
R961 VTAIL.n15 VTAIL.n12 7.3702
R962 VTAIL.n57 VTAIL.n54 7.3702
R963 VTAIL.n99 VTAIL.n96 7.3702
R964 VTAIL.n268 VTAIL.n265 7.3702
R965 VTAIL.n226 VTAIL.n223 7.3702
R966 VTAIL.n184 VTAIL.n181 7.3702
R967 VTAIL.n142 VTAIL.n139 7.3702
R968 VTAIL.n310 VTAIL.n309 5.81868
R969 VTAIL.n16 VTAIL.n15 5.81868
R970 VTAIL.n58 VTAIL.n57 5.81868
R971 VTAIL.n100 VTAIL.n99 5.81868
R972 VTAIL.n269 VTAIL.n268 5.81868
R973 VTAIL.n227 VTAIL.n226 5.81868
R974 VTAIL.n185 VTAIL.n184 5.81868
R975 VTAIL.n143 VTAIL.n142 5.81868
R976 VTAIL.n313 VTAIL.n304 5.04292
R977 VTAIL.n19 VTAIL.n10 5.04292
R978 VTAIL.n61 VTAIL.n52 5.04292
R979 VTAIL.n103 VTAIL.n94 5.04292
R980 VTAIL.n272 VTAIL.n263 5.04292
R981 VTAIL.n230 VTAIL.n221 5.04292
R982 VTAIL.n188 VTAIL.n179 5.04292
R983 VTAIL.n146 VTAIL.n137 5.04292
R984 VTAIL.n314 VTAIL.n302 4.26717
R985 VTAIL.n20 VTAIL.n8 4.26717
R986 VTAIL.n62 VTAIL.n50 4.26717
R987 VTAIL.n104 VTAIL.n92 4.26717
R988 VTAIL.n273 VTAIL.n261 4.26717
R989 VTAIL.n231 VTAIL.n219 4.26717
R990 VTAIL.n189 VTAIL.n177 4.26717
R991 VTAIL.n147 VTAIL.n135 4.26717
R992 VTAIL.n318 VTAIL.n317 3.49141
R993 VTAIL.n24 VTAIL.n23 3.49141
R994 VTAIL.n66 VTAIL.n65 3.49141
R995 VTAIL.n108 VTAIL.n107 3.49141
R996 VTAIL.n277 VTAIL.n276 3.49141
R997 VTAIL.n235 VTAIL.n234 3.49141
R998 VTAIL.n193 VTAIL.n192 3.49141
R999 VTAIL.n151 VTAIL.n150 3.49141
R1000 VTAIL.n321 VTAIL.n300 2.71565
R1001 VTAIL.n27 VTAIL.n6 2.71565
R1002 VTAIL.n69 VTAIL.n48 2.71565
R1003 VTAIL.n111 VTAIL.n90 2.71565
R1004 VTAIL.n280 VTAIL.n259 2.71565
R1005 VTAIL.n238 VTAIL.n217 2.71565
R1006 VTAIL.n196 VTAIL.n175 2.71565
R1007 VTAIL.n154 VTAIL.n133 2.71565
R1008 VTAIL.n308 VTAIL.n307 2.4129
R1009 VTAIL.n14 VTAIL.n13 2.4129
R1010 VTAIL.n56 VTAIL.n55 2.4129
R1011 VTAIL.n98 VTAIL.n97 2.4129
R1012 VTAIL.n267 VTAIL.n266 2.4129
R1013 VTAIL.n225 VTAIL.n224 2.4129
R1014 VTAIL.n183 VTAIL.n182 2.4129
R1015 VTAIL.n141 VTAIL.n140 2.4129
R1016 VTAIL.n322 VTAIL.n298 1.93989
R1017 VTAIL.n28 VTAIL.n4 1.93989
R1018 VTAIL.n70 VTAIL.n46 1.93989
R1019 VTAIL.n112 VTAIL.n88 1.93989
R1020 VTAIL.n281 VTAIL.n257 1.93989
R1021 VTAIL.n239 VTAIL.n215 1.93989
R1022 VTAIL.n197 VTAIL.n173 1.93989
R1023 VTAIL.n155 VTAIL.n131 1.93989
R1024 VTAIL.n327 VTAIL.n325 1.16414
R1025 VTAIL.n334 VTAIL.n294 1.16414
R1026 VTAIL.n33 VTAIL.n31 1.16414
R1027 VTAIL.n40 VTAIL.n0 1.16414
R1028 VTAIL.n75 VTAIL.n73 1.16414
R1029 VTAIL.n82 VTAIL.n42 1.16414
R1030 VTAIL.n117 VTAIL.n115 1.16414
R1031 VTAIL.n124 VTAIL.n84 1.16414
R1032 VTAIL.n292 VTAIL.n252 1.16414
R1033 VTAIL.n285 VTAIL.n284 1.16414
R1034 VTAIL.n250 VTAIL.n210 1.16414
R1035 VTAIL.n243 VTAIL.n242 1.16414
R1036 VTAIL.n208 VTAIL.n168 1.16414
R1037 VTAIL.n201 VTAIL.n200 1.16414
R1038 VTAIL.n166 VTAIL.n126 1.16414
R1039 VTAIL.n159 VTAIL.n158 1.16414
R1040 VTAIL.n209 VTAIL.n167 0.483259
R1041 VTAIL.n293 VTAIL.n251 0.483259
R1042 VTAIL.n125 VTAIL.n83 0.483259
R1043 VTAIL.n251 VTAIL.n209 0.470328
R1044 VTAIL.n83 VTAIL.n41 0.470328
R1045 VTAIL.n326 VTAIL.n296 0.388379
R1046 VTAIL.n332 VTAIL.n331 0.388379
R1047 VTAIL.n32 VTAIL.n2 0.388379
R1048 VTAIL.n38 VTAIL.n37 0.388379
R1049 VTAIL.n74 VTAIL.n44 0.388379
R1050 VTAIL.n80 VTAIL.n79 0.388379
R1051 VTAIL.n116 VTAIL.n86 0.388379
R1052 VTAIL.n122 VTAIL.n121 0.388379
R1053 VTAIL.n290 VTAIL.n289 0.388379
R1054 VTAIL.n256 VTAIL.n254 0.388379
R1055 VTAIL.n248 VTAIL.n247 0.388379
R1056 VTAIL.n214 VTAIL.n212 0.388379
R1057 VTAIL.n206 VTAIL.n205 0.388379
R1058 VTAIL.n172 VTAIL.n170 0.388379
R1059 VTAIL.n164 VTAIL.n163 0.388379
R1060 VTAIL.n130 VTAIL.n128 0.388379
R1061 VTAIL VTAIL.n41 0.300069
R1062 VTAIL VTAIL.n335 0.18369
R1063 VTAIL.n308 VTAIL.n303 0.155672
R1064 VTAIL.n315 VTAIL.n303 0.155672
R1065 VTAIL.n316 VTAIL.n315 0.155672
R1066 VTAIL.n316 VTAIL.n299 0.155672
R1067 VTAIL.n323 VTAIL.n299 0.155672
R1068 VTAIL.n324 VTAIL.n323 0.155672
R1069 VTAIL.n324 VTAIL.n295 0.155672
R1070 VTAIL.n333 VTAIL.n295 0.155672
R1071 VTAIL.n14 VTAIL.n9 0.155672
R1072 VTAIL.n21 VTAIL.n9 0.155672
R1073 VTAIL.n22 VTAIL.n21 0.155672
R1074 VTAIL.n22 VTAIL.n5 0.155672
R1075 VTAIL.n29 VTAIL.n5 0.155672
R1076 VTAIL.n30 VTAIL.n29 0.155672
R1077 VTAIL.n30 VTAIL.n1 0.155672
R1078 VTAIL.n39 VTAIL.n1 0.155672
R1079 VTAIL.n56 VTAIL.n51 0.155672
R1080 VTAIL.n63 VTAIL.n51 0.155672
R1081 VTAIL.n64 VTAIL.n63 0.155672
R1082 VTAIL.n64 VTAIL.n47 0.155672
R1083 VTAIL.n71 VTAIL.n47 0.155672
R1084 VTAIL.n72 VTAIL.n71 0.155672
R1085 VTAIL.n72 VTAIL.n43 0.155672
R1086 VTAIL.n81 VTAIL.n43 0.155672
R1087 VTAIL.n98 VTAIL.n93 0.155672
R1088 VTAIL.n105 VTAIL.n93 0.155672
R1089 VTAIL.n106 VTAIL.n105 0.155672
R1090 VTAIL.n106 VTAIL.n89 0.155672
R1091 VTAIL.n113 VTAIL.n89 0.155672
R1092 VTAIL.n114 VTAIL.n113 0.155672
R1093 VTAIL.n114 VTAIL.n85 0.155672
R1094 VTAIL.n123 VTAIL.n85 0.155672
R1095 VTAIL.n291 VTAIL.n253 0.155672
R1096 VTAIL.n283 VTAIL.n253 0.155672
R1097 VTAIL.n283 VTAIL.n282 0.155672
R1098 VTAIL.n282 VTAIL.n258 0.155672
R1099 VTAIL.n275 VTAIL.n258 0.155672
R1100 VTAIL.n275 VTAIL.n274 0.155672
R1101 VTAIL.n274 VTAIL.n262 0.155672
R1102 VTAIL.n267 VTAIL.n262 0.155672
R1103 VTAIL.n249 VTAIL.n211 0.155672
R1104 VTAIL.n241 VTAIL.n211 0.155672
R1105 VTAIL.n241 VTAIL.n240 0.155672
R1106 VTAIL.n240 VTAIL.n216 0.155672
R1107 VTAIL.n233 VTAIL.n216 0.155672
R1108 VTAIL.n233 VTAIL.n232 0.155672
R1109 VTAIL.n232 VTAIL.n220 0.155672
R1110 VTAIL.n225 VTAIL.n220 0.155672
R1111 VTAIL.n207 VTAIL.n169 0.155672
R1112 VTAIL.n199 VTAIL.n169 0.155672
R1113 VTAIL.n199 VTAIL.n198 0.155672
R1114 VTAIL.n198 VTAIL.n174 0.155672
R1115 VTAIL.n191 VTAIL.n174 0.155672
R1116 VTAIL.n191 VTAIL.n190 0.155672
R1117 VTAIL.n190 VTAIL.n178 0.155672
R1118 VTAIL.n183 VTAIL.n178 0.155672
R1119 VTAIL.n165 VTAIL.n127 0.155672
R1120 VTAIL.n157 VTAIL.n127 0.155672
R1121 VTAIL.n157 VTAIL.n156 0.155672
R1122 VTAIL.n156 VTAIL.n132 0.155672
R1123 VTAIL.n149 VTAIL.n132 0.155672
R1124 VTAIL.n149 VTAIL.n148 0.155672
R1125 VTAIL.n148 VTAIL.n136 0.155672
R1126 VTAIL.n141 VTAIL.n136 0.155672
R1127 VDD1 VDD1.n1 119.65
R1128 VDD1 VDD1.n0 87.0718
R1129 VDD1.n0 VDD1.t0 4.04341
R1130 VDD1.n0 VDD1.t1 4.04341
R1131 VDD1.n1 VDD1.t2 4.04341
R1132 VDD1.n1 VDD1.t3 4.04341
R1133 VN.n0 VN.t3 1019.57
R1134 VN.n0 VN.t1 1019.57
R1135 VN.n1 VN.t0 1019.57
R1136 VN.n1 VN.t2 1019.57
R1137 VN VN.n1 197.703
R1138 VN VN.n0 161.351
R1139 VDD2.n2 VDD2.n0 119.124
R1140 VDD2.n2 VDD2.n1 87.0136
R1141 VDD2.n1 VDD2.t3 4.04341
R1142 VDD2.n1 VDD2.t1 4.04341
R1143 VDD2.n0 VDD2.t2 4.04341
R1144 VDD2.n0 VDD2.t0 4.04341
R1145 VDD2 VDD2.n2 0.0586897
C0 VP w_n1306_n2580# 1.86742f
C1 VN w_n1306_n2580# 1.70552f
C2 VDD1 VDD2 0.464214f
C3 w_n1306_n2580# B 5.26815f
C4 VN VP 3.74472f
C5 VP B 0.867064f
C6 VDD2 VTAIL 7.44021f
C7 VN B 0.609432f
C8 VDD1 w_n1306_n2580# 0.844837f
C9 VDD1 VP 1.40553f
C10 VTAIL w_n1306_n2580# 3.22889f
C11 VDD1 VN 0.14833f
C12 VTAIL VP 0.948809f
C13 VDD1 B 0.735889f
C14 VN VTAIL 0.934703f
C15 VTAIL B 2.46563f
C16 VDD2 w_n1306_n2580# 0.850297f
C17 VDD2 VP 0.244971f
C18 VN VDD2 1.30903f
C19 VDD2 B 0.75099f
C20 VDD1 VTAIL 7.40189f
C21 VDD2 VSUBS 0.516426f
C22 VDD1 VSUBS 4.171023f
C23 VTAIL VSUBS 0.228561f
C24 VN VSUBS 3.67963f
C25 VP VSUBS 0.894991f
C26 B VSUBS 1.88554f
C27 w_n1306_n2580# VSUBS 41.7972f
C28 VDD2.t2 VSUBS 0.185375f
C29 VDD2.t0 VSUBS 0.185375f
C30 VDD2.n0 VSUBS 1.78752f
C31 VDD2.t3 VSUBS 0.185375f
C32 VDD2.t1 VSUBS 0.185375f
C33 VDD2.n1 VSUBS 1.3497f
C34 VDD2.n2 VSUBS 3.46961f
C35 VN.t1 VSUBS 0.204264f
C36 VN.t3 VSUBS 0.204264f
C37 VN.n0 VSUBS 0.184575f
C38 VN.t0 VSUBS 0.204264f
C39 VN.t2 VSUBS 0.204264f
C40 VN.n1 VSUBS 0.412157f
C41 VDD1.t0 VSUBS 0.182714f
C42 VDD1.t1 VSUBS 0.182714f
C43 VDD1.n0 VSUBS 1.33069f
C44 VDD1.t2 VSUBS 0.182714f
C45 VDD1.t3 VSUBS 0.182714f
C46 VDD1.n1 VSUBS 1.78313f
C47 VTAIL.n0 VSUBS 0.028037f
C48 VTAIL.n1 VSUBS 0.025614f
C49 VTAIL.n2 VSUBS 0.014169f
C50 VTAIL.n3 VSUBS 0.032533f
C51 VTAIL.n4 VSUBS 0.014573f
C52 VTAIL.n5 VSUBS 0.025614f
C53 VTAIL.n6 VSUBS 0.013764f
C54 VTAIL.n7 VSUBS 0.032533f
C55 VTAIL.n8 VSUBS 0.014573f
C56 VTAIL.n9 VSUBS 0.025614f
C57 VTAIL.n10 VSUBS 0.013764f
C58 VTAIL.n11 VSUBS 0.024399f
C59 VTAIL.n12 VSUBS 0.024472f
C60 VTAIL.t2 VSUBS 0.069908f
C61 VTAIL.n13 VSUBS 0.155985f
C62 VTAIL.n14 VSUBS 0.813787f
C63 VTAIL.n15 VSUBS 0.013764f
C64 VTAIL.n16 VSUBS 0.014573f
C65 VTAIL.n17 VSUBS 0.032533f
C66 VTAIL.n18 VSUBS 0.032533f
C67 VTAIL.n19 VSUBS 0.014573f
C68 VTAIL.n20 VSUBS 0.013764f
C69 VTAIL.n21 VSUBS 0.025614f
C70 VTAIL.n22 VSUBS 0.025614f
C71 VTAIL.n23 VSUBS 0.013764f
C72 VTAIL.n24 VSUBS 0.014573f
C73 VTAIL.n25 VSUBS 0.032533f
C74 VTAIL.n26 VSUBS 0.032533f
C75 VTAIL.n27 VSUBS 0.014573f
C76 VTAIL.n28 VSUBS 0.013764f
C77 VTAIL.n29 VSUBS 0.025614f
C78 VTAIL.n30 VSUBS 0.025614f
C79 VTAIL.n31 VSUBS 0.013764f
C80 VTAIL.n32 VSUBS 0.013764f
C81 VTAIL.n33 VSUBS 0.014573f
C82 VTAIL.n34 VSUBS 0.032533f
C83 VTAIL.n35 VSUBS 0.032533f
C84 VTAIL.n36 VSUBS 0.078393f
C85 VTAIL.n37 VSUBS 0.014169f
C86 VTAIL.n38 VSUBS 0.013764f
C87 VTAIL.n39 VSUBS 0.067603f
C88 VTAIL.n40 VSUBS 0.03965f
C89 VTAIL.n41 VSUBS 0.090132f
C90 VTAIL.n42 VSUBS 0.028037f
C91 VTAIL.n43 VSUBS 0.025614f
C92 VTAIL.n44 VSUBS 0.014169f
C93 VTAIL.n45 VSUBS 0.032533f
C94 VTAIL.n46 VSUBS 0.014573f
C95 VTAIL.n47 VSUBS 0.025614f
C96 VTAIL.n48 VSUBS 0.013764f
C97 VTAIL.n49 VSUBS 0.032533f
C98 VTAIL.n50 VSUBS 0.014573f
C99 VTAIL.n51 VSUBS 0.025614f
C100 VTAIL.n52 VSUBS 0.013764f
C101 VTAIL.n53 VSUBS 0.024399f
C102 VTAIL.n54 VSUBS 0.024472f
C103 VTAIL.t6 VSUBS 0.069908f
C104 VTAIL.n55 VSUBS 0.155985f
C105 VTAIL.n56 VSUBS 0.813787f
C106 VTAIL.n57 VSUBS 0.013764f
C107 VTAIL.n58 VSUBS 0.014573f
C108 VTAIL.n59 VSUBS 0.032533f
C109 VTAIL.n60 VSUBS 0.032533f
C110 VTAIL.n61 VSUBS 0.014573f
C111 VTAIL.n62 VSUBS 0.013764f
C112 VTAIL.n63 VSUBS 0.025614f
C113 VTAIL.n64 VSUBS 0.025614f
C114 VTAIL.n65 VSUBS 0.013764f
C115 VTAIL.n66 VSUBS 0.014573f
C116 VTAIL.n67 VSUBS 0.032533f
C117 VTAIL.n68 VSUBS 0.032533f
C118 VTAIL.n69 VSUBS 0.014573f
C119 VTAIL.n70 VSUBS 0.013764f
C120 VTAIL.n71 VSUBS 0.025614f
C121 VTAIL.n72 VSUBS 0.025614f
C122 VTAIL.n73 VSUBS 0.013764f
C123 VTAIL.n74 VSUBS 0.013764f
C124 VTAIL.n75 VSUBS 0.014573f
C125 VTAIL.n76 VSUBS 0.032533f
C126 VTAIL.n77 VSUBS 0.032533f
C127 VTAIL.n78 VSUBS 0.078393f
C128 VTAIL.n79 VSUBS 0.014169f
C129 VTAIL.n80 VSUBS 0.013764f
C130 VTAIL.n81 VSUBS 0.067603f
C131 VTAIL.n82 VSUBS 0.03965f
C132 VTAIL.n83 VSUBS 0.105251f
C133 VTAIL.n84 VSUBS 0.028037f
C134 VTAIL.n85 VSUBS 0.025614f
C135 VTAIL.n86 VSUBS 0.014169f
C136 VTAIL.n87 VSUBS 0.032533f
C137 VTAIL.n88 VSUBS 0.014573f
C138 VTAIL.n89 VSUBS 0.025614f
C139 VTAIL.n90 VSUBS 0.013764f
C140 VTAIL.n91 VSUBS 0.032533f
C141 VTAIL.n92 VSUBS 0.014573f
C142 VTAIL.n93 VSUBS 0.025614f
C143 VTAIL.n94 VSUBS 0.013764f
C144 VTAIL.n95 VSUBS 0.024399f
C145 VTAIL.n96 VSUBS 0.024472f
C146 VTAIL.t4 VSUBS 0.069908f
C147 VTAIL.n97 VSUBS 0.155985f
C148 VTAIL.n98 VSUBS 0.813787f
C149 VTAIL.n99 VSUBS 0.013764f
C150 VTAIL.n100 VSUBS 0.014573f
C151 VTAIL.n101 VSUBS 0.032533f
C152 VTAIL.n102 VSUBS 0.032533f
C153 VTAIL.n103 VSUBS 0.014573f
C154 VTAIL.n104 VSUBS 0.013764f
C155 VTAIL.n105 VSUBS 0.025614f
C156 VTAIL.n106 VSUBS 0.025614f
C157 VTAIL.n107 VSUBS 0.013764f
C158 VTAIL.n108 VSUBS 0.014573f
C159 VTAIL.n109 VSUBS 0.032533f
C160 VTAIL.n110 VSUBS 0.032533f
C161 VTAIL.n111 VSUBS 0.014573f
C162 VTAIL.n112 VSUBS 0.013764f
C163 VTAIL.n113 VSUBS 0.025614f
C164 VTAIL.n114 VSUBS 0.025614f
C165 VTAIL.n115 VSUBS 0.013764f
C166 VTAIL.n116 VSUBS 0.013764f
C167 VTAIL.n117 VSUBS 0.014573f
C168 VTAIL.n118 VSUBS 0.032533f
C169 VTAIL.n119 VSUBS 0.032533f
C170 VTAIL.n120 VSUBS 0.078393f
C171 VTAIL.n121 VSUBS 0.014169f
C172 VTAIL.n122 VSUBS 0.013764f
C173 VTAIL.n123 VSUBS 0.067603f
C174 VTAIL.n124 VSUBS 0.03965f
C175 VTAIL.n125 VSUBS 1.02772f
C176 VTAIL.n126 VSUBS 0.028037f
C177 VTAIL.n127 VSUBS 0.025614f
C178 VTAIL.n128 VSUBS 0.014169f
C179 VTAIL.n129 VSUBS 0.032533f
C180 VTAIL.n130 VSUBS 0.013764f
C181 VTAIL.n131 VSUBS 0.014573f
C182 VTAIL.n132 VSUBS 0.025614f
C183 VTAIL.n133 VSUBS 0.013764f
C184 VTAIL.n134 VSUBS 0.032533f
C185 VTAIL.n135 VSUBS 0.014573f
C186 VTAIL.n136 VSUBS 0.025614f
C187 VTAIL.n137 VSUBS 0.013764f
C188 VTAIL.n138 VSUBS 0.024399f
C189 VTAIL.n139 VSUBS 0.024472f
C190 VTAIL.t3 VSUBS 0.069908f
C191 VTAIL.n140 VSUBS 0.155985f
C192 VTAIL.n141 VSUBS 0.813787f
C193 VTAIL.n142 VSUBS 0.013764f
C194 VTAIL.n143 VSUBS 0.014573f
C195 VTAIL.n144 VSUBS 0.032533f
C196 VTAIL.n145 VSUBS 0.032533f
C197 VTAIL.n146 VSUBS 0.014573f
C198 VTAIL.n147 VSUBS 0.013764f
C199 VTAIL.n148 VSUBS 0.025614f
C200 VTAIL.n149 VSUBS 0.025614f
C201 VTAIL.n150 VSUBS 0.013764f
C202 VTAIL.n151 VSUBS 0.014573f
C203 VTAIL.n152 VSUBS 0.032533f
C204 VTAIL.n153 VSUBS 0.032533f
C205 VTAIL.n154 VSUBS 0.014573f
C206 VTAIL.n155 VSUBS 0.013764f
C207 VTAIL.n156 VSUBS 0.025614f
C208 VTAIL.n157 VSUBS 0.025614f
C209 VTAIL.n158 VSUBS 0.013764f
C210 VTAIL.n159 VSUBS 0.014573f
C211 VTAIL.n160 VSUBS 0.032533f
C212 VTAIL.n161 VSUBS 0.032533f
C213 VTAIL.n162 VSUBS 0.078393f
C214 VTAIL.n163 VSUBS 0.014169f
C215 VTAIL.n164 VSUBS 0.013764f
C216 VTAIL.n165 VSUBS 0.067603f
C217 VTAIL.n166 VSUBS 0.03965f
C218 VTAIL.n167 VSUBS 1.02772f
C219 VTAIL.n168 VSUBS 0.028037f
C220 VTAIL.n169 VSUBS 0.025614f
C221 VTAIL.n170 VSUBS 0.014169f
C222 VTAIL.n171 VSUBS 0.032533f
C223 VTAIL.n172 VSUBS 0.013764f
C224 VTAIL.n173 VSUBS 0.014573f
C225 VTAIL.n174 VSUBS 0.025614f
C226 VTAIL.n175 VSUBS 0.013764f
C227 VTAIL.n176 VSUBS 0.032533f
C228 VTAIL.n177 VSUBS 0.014573f
C229 VTAIL.n178 VSUBS 0.025614f
C230 VTAIL.n179 VSUBS 0.013764f
C231 VTAIL.n180 VSUBS 0.024399f
C232 VTAIL.n181 VSUBS 0.024472f
C233 VTAIL.t1 VSUBS 0.069908f
C234 VTAIL.n182 VSUBS 0.155985f
C235 VTAIL.n183 VSUBS 0.813787f
C236 VTAIL.n184 VSUBS 0.013764f
C237 VTAIL.n185 VSUBS 0.014573f
C238 VTAIL.n186 VSUBS 0.032533f
C239 VTAIL.n187 VSUBS 0.032533f
C240 VTAIL.n188 VSUBS 0.014573f
C241 VTAIL.n189 VSUBS 0.013764f
C242 VTAIL.n190 VSUBS 0.025614f
C243 VTAIL.n191 VSUBS 0.025614f
C244 VTAIL.n192 VSUBS 0.013764f
C245 VTAIL.n193 VSUBS 0.014573f
C246 VTAIL.n194 VSUBS 0.032533f
C247 VTAIL.n195 VSUBS 0.032533f
C248 VTAIL.n196 VSUBS 0.014573f
C249 VTAIL.n197 VSUBS 0.013764f
C250 VTAIL.n198 VSUBS 0.025614f
C251 VTAIL.n199 VSUBS 0.025614f
C252 VTAIL.n200 VSUBS 0.013764f
C253 VTAIL.n201 VSUBS 0.014573f
C254 VTAIL.n202 VSUBS 0.032533f
C255 VTAIL.n203 VSUBS 0.032533f
C256 VTAIL.n204 VSUBS 0.078393f
C257 VTAIL.n205 VSUBS 0.014169f
C258 VTAIL.n206 VSUBS 0.013764f
C259 VTAIL.n207 VSUBS 0.067603f
C260 VTAIL.n208 VSUBS 0.03965f
C261 VTAIL.n209 VSUBS 0.105251f
C262 VTAIL.n210 VSUBS 0.028037f
C263 VTAIL.n211 VSUBS 0.025614f
C264 VTAIL.n212 VSUBS 0.014169f
C265 VTAIL.n213 VSUBS 0.032533f
C266 VTAIL.n214 VSUBS 0.013764f
C267 VTAIL.n215 VSUBS 0.014573f
C268 VTAIL.n216 VSUBS 0.025614f
C269 VTAIL.n217 VSUBS 0.013764f
C270 VTAIL.n218 VSUBS 0.032533f
C271 VTAIL.n219 VSUBS 0.014573f
C272 VTAIL.n220 VSUBS 0.025614f
C273 VTAIL.n221 VSUBS 0.013764f
C274 VTAIL.n222 VSUBS 0.024399f
C275 VTAIL.n223 VSUBS 0.024472f
C276 VTAIL.t7 VSUBS 0.069908f
C277 VTAIL.n224 VSUBS 0.155985f
C278 VTAIL.n225 VSUBS 0.813787f
C279 VTAIL.n226 VSUBS 0.013764f
C280 VTAIL.n227 VSUBS 0.014573f
C281 VTAIL.n228 VSUBS 0.032533f
C282 VTAIL.n229 VSUBS 0.032533f
C283 VTAIL.n230 VSUBS 0.014573f
C284 VTAIL.n231 VSUBS 0.013764f
C285 VTAIL.n232 VSUBS 0.025614f
C286 VTAIL.n233 VSUBS 0.025614f
C287 VTAIL.n234 VSUBS 0.013764f
C288 VTAIL.n235 VSUBS 0.014573f
C289 VTAIL.n236 VSUBS 0.032533f
C290 VTAIL.n237 VSUBS 0.032533f
C291 VTAIL.n238 VSUBS 0.014573f
C292 VTAIL.n239 VSUBS 0.013764f
C293 VTAIL.n240 VSUBS 0.025614f
C294 VTAIL.n241 VSUBS 0.025614f
C295 VTAIL.n242 VSUBS 0.013764f
C296 VTAIL.n243 VSUBS 0.014573f
C297 VTAIL.n244 VSUBS 0.032533f
C298 VTAIL.n245 VSUBS 0.032533f
C299 VTAIL.n246 VSUBS 0.078393f
C300 VTAIL.n247 VSUBS 0.014169f
C301 VTAIL.n248 VSUBS 0.013764f
C302 VTAIL.n249 VSUBS 0.067603f
C303 VTAIL.n250 VSUBS 0.03965f
C304 VTAIL.n251 VSUBS 0.105251f
C305 VTAIL.n252 VSUBS 0.028037f
C306 VTAIL.n253 VSUBS 0.025614f
C307 VTAIL.n254 VSUBS 0.014169f
C308 VTAIL.n255 VSUBS 0.032533f
C309 VTAIL.n256 VSUBS 0.013764f
C310 VTAIL.n257 VSUBS 0.014573f
C311 VTAIL.n258 VSUBS 0.025614f
C312 VTAIL.n259 VSUBS 0.013764f
C313 VTAIL.n260 VSUBS 0.032533f
C314 VTAIL.n261 VSUBS 0.014573f
C315 VTAIL.n262 VSUBS 0.025614f
C316 VTAIL.n263 VSUBS 0.013764f
C317 VTAIL.n264 VSUBS 0.024399f
C318 VTAIL.n265 VSUBS 0.024472f
C319 VTAIL.t5 VSUBS 0.069908f
C320 VTAIL.n266 VSUBS 0.155985f
C321 VTAIL.n267 VSUBS 0.813787f
C322 VTAIL.n268 VSUBS 0.013764f
C323 VTAIL.n269 VSUBS 0.014573f
C324 VTAIL.n270 VSUBS 0.032533f
C325 VTAIL.n271 VSUBS 0.032533f
C326 VTAIL.n272 VSUBS 0.014573f
C327 VTAIL.n273 VSUBS 0.013764f
C328 VTAIL.n274 VSUBS 0.025614f
C329 VTAIL.n275 VSUBS 0.025614f
C330 VTAIL.n276 VSUBS 0.013764f
C331 VTAIL.n277 VSUBS 0.014573f
C332 VTAIL.n278 VSUBS 0.032533f
C333 VTAIL.n279 VSUBS 0.032533f
C334 VTAIL.n280 VSUBS 0.014573f
C335 VTAIL.n281 VSUBS 0.013764f
C336 VTAIL.n282 VSUBS 0.025614f
C337 VTAIL.n283 VSUBS 0.025614f
C338 VTAIL.n284 VSUBS 0.013764f
C339 VTAIL.n285 VSUBS 0.014573f
C340 VTAIL.n286 VSUBS 0.032533f
C341 VTAIL.n287 VSUBS 0.032533f
C342 VTAIL.n288 VSUBS 0.078393f
C343 VTAIL.n289 VSUBS 0.014169f
C344 VTAIL.n290 VSUBS 0.013764f
C345 VTAIL.n291 VSUBS 0.067603f
C346 VTAIL.n292 VSUBS 0.03965f
C347 VTAIL.n293 VSUBS 1.02772f
C348 VTAIL.n294 VSUBS 0.028037f
C349 VTAIL.n295 VSUBS 0.025614f
C350 VTAIL.n296 VSUBS 0.014169f
C351 VTAIL.n297 VSUBS 0.032533f
C352 VTAIL.n298 VSUBS 0.014573f
C353 VTAIL.n299 VSUBS 0.025614f
C354 VTAIL.n300 VSUBS 0.013764f
C355 VTAIL.n301 VSUBS 0.032533f
C356 VTAIL.n302 VSUBS 0.014573f
C357 VTAIL.n303 VSUBS 0.025614f
C358 VTAIL.n304 VSUBS 0.013764f
C359 VTAIL.n305 VSUBS 0.024399f
C360 VTAIL.n306 VSUBS 0.024472f
C361 VTAIL.t0 VSUBS 0.069908f
C362 VTAIL.n307 VSUBS 0.155985f
C363 VTAIL.n308 VSUBS 0.813787f
C364 VTAIL.n309 VSUBS 0.013764f
C365 VTAIL.n310 VSUBS 0.014573f
C366 VTAIL.n311 VSUBS 0.032533f
C367 VTAIL.n312 VSUBS 0.032533f
C368 VTAIL.n313 VSUBS 0.014573f
C369 VTAIL.n314 VSUBS 0.013764f
C370 VTAIL.n315 VSUBS 0.025614f
C371 VTAIL.n316 VSUBS 0.025614f
C372 VTAIL.n317 VSUBS 0.013764f
C373 VTAIL.n318 VSUBS 0.014573f
C374 VTAIL.n319 VSUBS 0.032533f
C375 VTAIL.n320 VSUBS 0.032533f
C376 VTAIL.n321 VSUBS 0.014573f
C377 VTAIL.n322 VSUBS 0.013764f
C378 VTAIL.n323 VSUBS 0.025614f
C379 VTAIL.n324 VSUBS 0.025614f
C380 VTAIL.n325 VSUBS 0.013764f
C381 VTAIL.n326 VSUBS 0.013764f
C382 VTAIL.n327 VSUBS 0.014573f
C383 VTAIL.n328 VSUBS 0.032533f
C384 VTAIL.n329 VSUBS 0.032533f
C385 VTAIL.n330 VSUBS 0.078393f
C386 VTAIL.n331 VSUBS 0.014169f
C387 VTAIL.n332 VSUBS 0.013764f
C388 VTAIL.n333 VSUBS 0.067603f
C389 VTAIL.n334 VSUBS 0.03965f
C390 VTAIL.n335 VSUBS 1.00299f
C391 VP.t3 VSUBS 0.207276f
C392 VP.t2 VSUBS 0.207276f
C393 VP.n0 VSUBS 0.41156f
C394 VP.t1 VSUBS 0.207276f
C395 VP.t0 VSUBS 0.207276f
C396 VP.n1 VSUBS 0.187286f
C397 VP.n2 VSUBS 2.25637f
C398 B.n0 VSUBS 0.005982f
C399 B.n1 VSUBS 0.005982f
C400 B.n2 VSUBS 0.00946f
C401 B.n3 VSUBS 0.00946f
C402 B.n4 VSUBS 0.00946f
C403 B.n5 VSUBS 0.00946f
C404 B.n6 VSUBS 0.00946f
C405 B.n7 VSUBS 0.00946f
C406 B.n8 VSUBS 0.020635f
C407 B.n9 VSUBS 0.00946f
C408 B.n10 VSUBS 0.00946f
C409 B.n11 VSUBS 0.00946f
C410 B.n12 VSUBS 0.00946f
C411 B.n13 VSUBS 0.00946f
C412 B.n14 VSUBS 0.00946f
C413 B.n15 VSUBS 0.00946f
C414 B.n16 VSUBS 0.00946f
C415 B.n17 VSUBS 0.00946f
C416 B.n18 VSUBS 0.00946f
C417 B.n19 VSUBS 0.00946f
C418 B.n20 VSUBS 0.00946f
C419 B.n21 VSUBS 0.00946f
C420 B.n22 VSUBS 0.00946f
C421 B.n23 VSUBS 0.00946f
C422 B.t11 VSUBS 0.172302f
C423 B.t10 VSUBS 0.180326f
C424 B.t9 VSUBS 0.098733f
C425 B.n24 VSUBS 0.265338f
C426 B.n25 VSUBS 0.246441f
C427 B.n26 VSUBS 0.00946f
C428 B.n27 VSUBS 0.00946f
C429 B.n28 VSUBS 0.00946f
C430 B.n29 VSUBS 0.00946f
C431 B.n30 VSUBS 0.005564f
C432 B.n31 VSUBS 0.00946f
C433 B.t8 VSUBS 0.172305f
C434 B.t7 VSUBS 0.180329f
C435 B.t6 VSUBS 0.098733f
C436 B.n32 VSUBS 0.265335f
C437 B.n33 VSUBS 0.246438f
C438 B.n34 VSUBS 0.021917f
C439 B.n35 VSUBS 0.00946f
C440 B.n36 VSUBS 0.00946f
C441 B.n37 VSUBS 0.00946f
C442 B.n38 VSUBS 0.00946f
C443 B.n39 VSUBS 0.00946f
C444 B.n40 VSUBS 0.00946f
C445 B.n41 VSUBS 0.00946f
C446 B.n42 VSUBS 0.00946f
C447 B.n43 VSUBS 0.00946f
C448 B.n44 VSUBS 0.00946f
C449 B.n45 VSUBS 0.00946f
C450 B.n46 VSUBS 0.00946f
C451 B.n47 VSUBS 0.00946f
C452 B.n48 VSUBS 0.022211f
C453 B.n49 VSUBS 0.00946f
C454 B.n50 VSUBS 0.00946f
C455 B.n51 VSUBS 0.00946f
C456 B.n52 VSUBS 0.00946f
C457 B.n53 VSUBS 0.00946f
C458 B.n54 VSUBS 0.00946f
C459 B.n55 VSUBS 0.00946f
C460 B.n56 VSUBS 0.00946f
C461 B.n57 VSUBS 0.00946f
C462 B.n58 VSUBS 0.00946f
C463 B.n59 VSUBS 0.00946f
C464 B.n60 VSUBS 0.00946f
C465 B.n61 VSUBS 0.00946f
C466 B.n62 VSUBS 0.022211f
C467 B.n63 VSUBS 0.00946f
C468 B.n64 VSUBS 0.00946f
C469 B.n65 VSUBS 0.00946f
C470 B.n66 VSUBS 0.00946f
C471 B.n67 VSUBS 0.00946f
C472 B.n68 VSUBS 0.00946f
C473 B.n69 VSUBS 0.00946f
C474 B.n70 VSUBS 0.00946f
C475 B.n71 VSUBS 0.00946f
C476 B.n72 VSUBS 0.00946f
C477 B.n73 VSUBS 0.00946f
C478 B.n74 VSUBS 0.00946f
C479 B.n75 VSUBS 0.00946f
C480 B.n76 VSUBS 0.00946f
C481 B.t4 VSUBS 0.172305f
C482 B.t5 VSUBS 0.180329f
C483 B.t3 VSUBS 0.098733f
C484 B.n77 VSUBS 0.265335f
C485 B.n78 VSUBS 0.246438f
C486 B.n79 VSUBS 0.021917f
C487 B.n80 VSUBS 0.00946f
C488 B.n81 VSUBS 0.00946f
C489 B.n82 VSUBS 0.00946f
C490 B.n83 VSUBS 0.00946f
C491 B.n84 VSUBS 0.00946f
C492 B.t1 VSUBS 0.172302f
C493 B.t2 VSUBS 0.180326f
C494 B.t0 VSUBS 0.098733f
C495 B.n85 VSUBS 0.265338f
C496 B.n86 VSUBS 0.246441f
C497 B.n87 VSUBS 0.00946f
C498 B.n88 VSUBS 0.00946f
C499 B.n89 VSUBS 0.00946f
C500 B.n90 VSUBS 0.00946f
C501 B.n91 VSUBS 0.00946f
C502 B.n92 VSUBS 0.00946f
C503 B.n93 VSUBS 0.00946f
C504 B.n94 VSUBS 0.00946f
C505 B.n95 VSUBS 0.00946f
C506 B.n96 VSUBS 0.00946f
C507 B.n97 VSUBS 0.00946f
C508 B.n98 VSUBS 0.00946f
C509 B.n99 VSUBS 0.00946f
C510 B.n100 VSUBS 0.00946f
C511 B.n101 VSUBS 0.022211f
C512 B.n102 VSUBS 0.00946f
C513 B.n103 VSUBS 0.00946f
C514 B.n104 VSUBS 0.00946f
C515 B.n105 VSUBS 0.00946f
C516 B.n106 VSUBS 0.00946f
C517 B.n107 VSUBS 0.00946f
C518 B.n108 VSUBS 0.00946f
C519 B.n109 VSUBS 0.00946f
C520 B.n110 VSUBS 0.00946f
C521 B.n111 VSUBS 0.00946f
C522 B.n112 VSUBS 0.00946f
C523 B.n113 VSUBS 0.00946f
C524 B.n114 VSUBS 0.00946f
C525 B.n115 VSUBS 0.00946f
C526 B.n116 VSUBS 0.00946f
C527 B.n117 VSUBS 0.00946f
C528 B.n118 VSUBS 0.00946f
C529 B.n119 VSUBS 0.00946f
C530 B.n120 VSUBS 0.00946f
C531 B.n121 VSUBS 0.00946f
C532 B.n122 VSUBS 0.00946f
C533 B.n123 VSUBS 0.00946f
C534 B.n124 VSUBS 0.020635f
C535 B.n125 VSUBS 0.020635f
C536 B.n126 VSUBS 0.022211f
C537 B.n127 VSUBS 0.00946f
C538 B.n128 VSUBS 0.00946f
C539 B.n129 VSUBS 0.00946f
C540 B.n130 VSUBS 0.00946f
C541 B.n131 VSUBS 0.00946f
C542 B.n132 VSUBS 0.00946f
C543 B.n133 VSUBS 0.00946f
C544 B.n134 VSUBS 0.00946f
C545 B.n135 VSUBS 0.00946f
C546 B.n136 VSUBS 0.00946f
C547 B.n137 VSUBS 0.00946f
C548 B.n138 VSUBS 0.00946f
C549 B.n139 VSUBS 0.00946f
C550 B.n140 VSUBS 0.00946f
C551 B.n141 VSUBS 0.00946f
C552 B.n142 VSUBS 0.00946f
C553 B.n143 VSUBS 0.00946f
C554 B.n144 VSUBS 0.00946f
C555 B.n145 VSUBS 0.00946f
C556 B.n146 VSUBS 0.00946f
C557 B.n147 VSUBS 0.00946f
C558 B.n148 VSUBS 0.00946f
C559 B.n149 VSUBS 0.00946f
C560 B.n150 VSUBS 0.00946f
C561 B.n151 VSUBS 0.00946f
C562 B.n152 VSUBS 0.00946f
C563 B.n153 VSUBS 0.00946f
C564 B.n154 VSUBS 0.00946f
C565 B.n155 VSUBS 0.00946f
C566 B.n156 VSUBS 0.00946f
C567 B.n157 VSUBS 0.00946f
C568 B.n158 VSUBS 0.00946f
C569 B.n159 VSUBS 0.00946f
C570 B.n160 VSUBS 0.00946f
C571 B.n161 VSUBS 0.00946f
C572 B.n162 VSUBS 0.00946f
C573 B.n163 VSUBS 0.00946f
C574 B.n164 VSUBS 0.00946f
C575 B.n165 VSUBS 0.00946f
C576 B.n166 VSUBS 0.00946f
C577 B.n167 VSUBS 0.00946f
C578 B.n168 VSUBS 0.00946f
C579 B.n169 VSUBS 0.00946f
C580 B.n170 VSUBS 0.008625f
C581 B.n171 VSUBS 0.021917f
C582 B.n172 VSUBS 0.005564f
C583 B.n173 VSUBS 0.00946f
C584 B.n174 VSUBS 0.00946f
C585 B.n175 VSUBS 0.00946f
C586 B.n176 VSUBS 0.00946f
C587 B.n177 VSUBS 0.00946f
C588 B.n178 VSUBS 0.00946f
C589 B.n179 VSUBS 0.00946f
C590 B.n180 VSUBS 0.00946f
C591 B.n181 VSUBS 0.00946f
C592 B.n182 VSUBS 0.00946f
C593 B.n183 VSUBS 0.00946f
C594 B.n184 VSUBS 0.00946f
C595 B.n185 VSUBS 0.005564f
C596 B.n186 VSUBS 0.00946f
C597 B.n187 VSUBS 0.00946f
C598 B.n188 VSUBS 0.008625f
C599 B.n189 VSUBS 0.00946f
C600 B.n190 VSUBS 0.00946f
C601 B.n191 VSUBS 0.00946f
C602 B.n192 VSUBS 0.00946f
C603 B.n193 VSUBS 0.00946f
C604 B.n194 VSUBS 0.00946f
C605 B.n195 VSUBS 0.00946f
C606 B.n196 VSUBS 0.00946f
C607 B.n197 VSUBS 0.00946f
C608 B.n198 VSUBS 0.00946f
C609 B.n199 VSUBS 0.00946f
C610 B.n200 VSUBS 0.00946f
C611 B.n201 VSUBS 0.00946f
C612 B.n202 VSUBS 0.00946f
C613 B.n203 VSUBS 0.00946f
C614 B.n204 VSUBS 0.00946f
C615 B.n205 VSUBS 0.00946f
C616 B.n206 VSUBS 0.00946f
C617 B.n207 VSUBS 0.00946f
C618 B.n208 VSUBS 0.00946f
C619 B.n209 VSUBS 0.00946f
C620 B.n210 VSUBS 0.00946f
C621 B.n211 VSUBS 0.00946f
C622 B.n212 VSUBS 0.00946f
C623 B.n213 VSUBS 0.00946f
C624 B.n214 VSUBS 0.00946f
C625 B.n215 VSUBS 0.00946f
C626 B.n216 VSUBS 0.00946f
C627 B.n217 VSUBS 0.00946f
C628 B.n218 VSUBS 0.00946f
C629 B.n219 VSUBS 0.00946f
C630 B.n220 VSUBS 0.00946f
C631 B.n221 VSUBS 0.00946f
C632 B.n222 VSUBS 0.00946f
C633 B.n223 VSUBS 0.00946f
C634 B.n224 VSUBS 0.00946f
C635 B.n225 VSUBS 0.00946f
C636 B.n226 VSUBS 0.00946f
C637 B.n227 VSUBS 0.00946f
C638 B.n228 VSUBS 0.00946f
C639 B.n229 VSUBS 0.00946f
C640 B.n230 VSUBS 0.00946f
C641 B.n231 VSUBS 0.022211f
C642 B.n232 VSUBS 0.020635f
C643 B.n233 VSUBS 0.020635f
C644 B.n234 VSUBS 0.00946f
C645 B.n235 VSUBS 0.00946f
C646 B.n236 VSUBS 0.00946f
C647 B.n237 VSUBS 0.00946f
C648 B.n238 VSUBS 0.00946f
C649 B.n239 VSUBS 0.00946f
C650 B.n240 VSUBS 0.00946f
C651 B.n241 VSUBS 0.00946f
C652 B.n242 VSUBS 0.00946f
C653 B.n243 VSUBS 0.00946f
C654 B.n244 VSUBS 0.00946f
C655 B.n245 VSUBS 0.00946f
C656 B.n246 VSUBS 0.00946f
C657 B.n247 VSUBS 0.00946f
C658 B.n248 VSUBS 0.00946f
C659 B.n249 VSUBS 0.00946f
C660 B.n250 VSUBS 0.00946f
C661 B.n251 VSUBS 0.00946f
C662 B.n252 VSUBS 0.00946f
C663 B.n253 VSUBS 0.00946f
C664 B.n254 VSUBS 0.00946f
C665 B.n255 VSUBS 0.00946f
C666 B.n256 VSUBS 0.00946f
C667 B.n257 VSUBS 0.00946f
C668 B.n258 VSUBS 0.00946f
C669 B.n259 VSUBS 0.00946f
C670 B.n260 VSUBS 0.00946f
C671 B.n261 VSUBS 0.00946f
C672 B.n262 VSUBS 0.00946f
C673 B.n263 VSUBS 0.00946f
C674 B.n264 VSUBS 0.00946f
C675 B.n265 VSUBS 0.00946f
C676 B.n266 VSUBS 0.00946f
C677 B.n267 VSUBS 0.00946f
C678 B.n268 VSUBS 0.00946f
C679 B.n269 VSUBS 0.00946f
C680 B.n270 VSUBS 0.00946f
C681 B.n271 VSUBS 0.020635f
C682 B.n272 VSUBS 0.02181f
C683 B.n273 VSUBS 0.021036f
C684 B.n274 VSUBS 0.00946f
C685 B.n275 VSUBS 0.00946f
C686 B.n276 VSUBS 0.00946f
C687 B.n277 VSUBS 0.00946f
C688 B.n278 VSUBS 0.00946f
C689 B.n279 VSUBS 0.00946f
C690 B.n280 VSUBS 0.00946f
C691 B.n281 VSUBS 0.00946f
C692 B.n282 VSUBS 0.00946f
C693 B.n283 VSUBS 0.00946f
C694 B.n284 VSUBS 0.00946f
C695 B.n285 VSUBS 0.00946f
C696 B.n286 VSUBS 0.00946f
C697 B.n287 VSUBS 0.00946f
C698 B.n288 VSUBS 0.00946f
C699 B.n289 VSUBS 0.00946f
C700 B.n290 VSUBS 0.00946f
C701 B.n291 VSUBS 0.00946f
C702 B.n292 VSUBS 0.00946f
C703 B.n293 VSUBS 0.00946f
C704 B.n294 VSUBS 0.00946f
C705 B.n295 VSUBS 0.00946f
C706 B.n296 VSUBS 0.00946f
C707 B.n297 VSUBS 0.00946f
C708 B.n298 VSUBS 0.00946f
C709 B.n299 VSUBS 0.00946f
C710 B.n300 VSUBS 0.00946f
C711 B.n301 VSUBS 0.00946f
C712 B.n302 VSUBS 0.00946f
C713 B.n303 VSUBS 0.00946f
C714 B.n304 VSUBS 0.00946f
C715 B.n305 VSUBS 0.00946f
C716 B.n306 VSUBS 0.00946f
C717 B.n307 VSUBS 0.00946f
C718 B.n308 VSUBS 0.00946f
C719 B.n309 VSUBS 0.00946f
C720 B.n310 VSUBS 0.00946f
C721 B.n311 VSUBS 0.00946f
C722 B.n312 VSUBS 0.00946f
C723 B.n313 VSUBS 0.00946f
C724 B.n314 VSUBS 0.00946f
C725 B.n315 VSUBS 0.00946f
C726 B.n316 VSUBS 0.008625f
C727 B.n317 VSUBS 0.00946f
C728 B.n318 VSUBS 0.00946f
C729 B.n319 VSUBS 0.00946f
C730 B.n320 VSUBS 0.00946f
C731 B.n321 VSUBS 0.00946f
C732 B.n322 VSUBS 0.00946f
C733 B.n323 VSUBS 0.00946f
C734 B.n324 VSUBS 0.00946f
C735 B.n325 VSUBS 0.00946f
C736 B.n326 VSUBS 0.00946f
C737 B.n327 VSUBS 0.00946f
C738 B.n328 VSUBS 0.00946f
C739 B.n329 VSUBS 0.00946f
C740 B.n330 VSUBS 0.00946f
C741 B.n331 VSUBS 0.00946f
C742 B.n332 VSUBS 0.005564f
C743 B.n333 VSUBS 0.021917f
C744 B.n334 VSUBS 0.008625f
C745 B.n335 VSUBS 0.00946f
C746 B.n336 VSUBS 0.00946f
C747 B.n337 VSUBS 0.00946f
C748 B.n338 VSUBS 0.00946f
C749 B.n339 VSUBS 0.00946f
C750 B.n340 VSUBS 0.00946f
C751 B.n341 VSUBS 0.00946f
C752 B.n342 VSUBS 0.00946f
C753 B.n343 VSUBS 0.00946f
C754 B.n344 VSUBS 0.00946f
C755 B.n345 VSUBS 0.00946f
C756 B.n346 VSUBS 0.00946f
C757 B.n347 VSUBS 0.00946f
C758 B.n348 VSUBS 0.00946f
C759 B.n349 VSUBS 0.00946f
C760 B.n350 VSUBS 0.00946f
C761 B.n351 VSUBS 0.00946f
C762 B.n352 VSUBS 0.00946f
C763 B.n353 VSUBS 0.00946f
C764 B.n354 VSUBS 0.00946f
C765 B.n355 VSUBS 0.00946f
C766 B.n356 VSUBS 0.00946f
C767 B.n357 VSUBS 0.00946f
C768 B.n358 VSUBS 0.00946f
C769 B.n359 VSUBS 0.00946f
C770 B.n360 VSUBS 0.00946f
C771 B.n361 VSUBS 0.00946f
C772 B.n362 VSUBS 0.00946f
C773 B.n363 VSUBS 0.00946f
C774 B.n364 VSUBS 0.00946f
C775 B.n365 VSUBS 0.00946f
C776 B.n366 VSUBS 0.00946f
C777 B.n367 VSUBS 0.00946f
C778 B.n368 VSUBS 0.00946f
C779 B.n369 VSUBS 0.00946f
C780 B.n370 VSUBS 0.00946f
C781 B.n371 VSUBS 0.00946f
C782 B.n372 VSUBS 0.00946f
C783 B.n373 VSUBS 0.00946f
C784 B.n374 VSUBS 0.00946f
C785 B.n375 VSUBS 0.00946f
C786 B.n376 VSUBS 0.00946f
C787 B.n377 VSUBS 0.022211f
C788 B.n378 VSUBS 0.022211f
C789 B.n379 VSUBS 0.020635f
C790 B.n380 VSUBS 0.00946f
C791 B.n381 VSUBS 0.00946f
C792 B.n382 VSUBS 0.00946f
C793 B.n383 VSUBS 0.00946f
C794 B.n384 VSUBS 0.00946f
C795 B.n385 VSUBS 0.00946f
C796 B.n386 VSUBS 0.00946f
C797 B.n387 VSUBS 0.00946f
C798 B.n388 VSUBS 0.00946f
C799 B.n389 VSUBS 0.00946f
C800 B.n390 VSUBS 0.00946f
C801 B.n391 VSUBS 0.00946f
C802 B.n392 VSUBS 0.00946f
C803 B.n393 VSUBS 0.00946f
C804 B.n394 VSUBS 0.00946f
C805 B.n395 VSUBS 0.00946f
C806 B.n396 VSUBS 0.00946f
C807 B.n397 VSUBS 0.00946f
C808 B.n398 VSUBS 0.00946f
C809 B.n399 VSUBS 0.02142f
.ends

