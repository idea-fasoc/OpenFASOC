* NGSPICE file created from diff_pair_sample_0405.ext - technology: sky130A

.subckt diff_pair_sample_0405 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=2.4258 ps=13.22 w=6.22 l=1.54
X1 VTAIL.t3 VN.t0 VDD2.t5 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=1.0263 ps=6.55 w=6.22 l=1.54
X2 VTAIL.t9 VP.t1 VDD1.t4 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=1.0263 ps=6.55 w=6.22 l=1.54
X3 VDD2.t4 VN.t1 VTAIL.t5 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=1.0263 ps=6.55 w=6.22 l=1.54
X4 B.t11 B.t9 B.t10 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=0 ps=0 w=6.22 l=1.54
X5 VDD1.t3 VP.t2 VTAIL.t6 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=1.0263 ps=6.55 w=6.22 l=1.54
X6 VDD2.t3 VN.t2 VTAIL.t4 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=2.4258 ps=13.22 w=6.22 l=1.54
X7 VDD1.t2 VP.t3 VTAIL.t7 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=2.4258 ps=13.22 w=6.22 l=1.54
X8 B.t8 B.t6 B.t7 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=0 ps=0 w=6.22 l=1.54
X9 VTAIL.t8 VP.t4 VDD1.t1 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=1.0263 ps=6.55 w=6.22 l=1.54
X10 VDD2.t2 VN.t3 VTAIL.t0 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=1.0263 ps=6.55 w=6.22 l=1.54
X11 VTAIL.t1 VN.t4 VDD2.t1 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=1.0263 ps=6.55 w=6.22 l=1.54
X12 B.t5 B.t3 B.t4 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=0 ps=0 w=6.22 l=1.54
X13 VDD1.t0 VP.t5 VTAIL.t10 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=1.0263 ps=6.55 w=6.22 l=1.54
X14 VDD2.t0 VN.t5 VTAIL.t2 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=1.0263 pd=6.55 as=2.4258 ps=13.22 w=6.22 l=1.54
X15 B.t2 B.t0 B.t1 w_n2466_n2212# sky130_fd_pr__pfet_01v8 ad=2.4258 pd=13.22 as=0 ps=0 w=6.22 l=1.54
R0 VP.n17 VP.n16 179.99
R1 VP.n32 VP.n31 179.99
R2 VP.n15 VP.n14 179.99
R3 VP.n9 VP.n8 161.3
R4 VP.n10 VP.n5 161.3
R5 VP.n12 VP.n11 161.3
R6 VP.n13 VP.n4 161.3
R7 VP.n30 VP.n0 161.3
R8 VP.n29 VP.n28 161.3
R9 VP.n27 VP.n1 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n23 VP.n2 161.3
R12 VP.n22 VP.n21 161.3
R13 VP.n20 VP.n3 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n6 VP.t5 128.93
R16 VP.n17 VP.t2 97.3395
R17 VP.n24 VP.t4 97.3395
R18 VP.n31 VP.t3 97.3395
R19 VP.n14 VP.t0 97.3395
R20 VP.n7 VP.t1 97.3395
R21 VP.n22 VP.n3 56.5617
R22 VP.n29 VP.n1 56.5617
R23 VP.n12 VP.n5 56.5617
R24 VP.n7 VP.n6 53.8793
R25 VP.n16 VP.n15 40.0119
R26 VP.n18 VP.n3 24.5923
R27 VP.n23 VP.n22 24.5923
R28 VP.n25 VP.n1 24.5923
R29 VP.n30 VP.n29 24.5923
R30 VP.n13 VP.n12 24.5923
R31 VP.n8 VP.n5 24.5923
R32 VP.n9 VP.n6 18.1684
R33 VP.n24 VP.n23 12.2964
R34 VP.n25 VP.n24 12.2964
R35 VP.n8 VP.n7 12.2964
R36 VP.n18 VP.n17 5.90254
R37 VP.n31 VP.n30 5.90254
R38 VP.n14 VP.n13 5.90254
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VTAIL.n7 VTAIL.t4 82.4386
R54 VTAIL.n11 VTAIL.t2 82.4376
R55 VTAIL.n2 VTAIL.t7 82.4376
R56 VTAIL.n10 VTAIL.t11 82.4376
R57 VTAIL.n9 VTAIL.n8 77.2127
R58 VTAIL.n6 VTAIL.n5 77.2127
R59 VTAIL.n1 VTAIL.n0 77.2126
R60 VTAIL.n4 VTAIL.n3 77.2126
R61 VTAIL.n6 VTAIL.n4 20.9531
R62 VTAIL.n11 VTAIL.n10 19.341
R63 VTAIL.n0 VTAIL.t5 5.22638
R64 VTAIL.n0 VTAIL.t3 5.22638
R65 VTAIL.n3 VTAIL.t6 5.22638
R66 VTAIL.n3 VTAIL.t8 5.22638
R67 VTAIL.n8 VTAIL.t10 5.22638
R68 VTAIL.n8 VTAIL.t9 5.22638
R69 VTAIL.n5 VTAIL.t0 5.22638
R70 VTAIL.n5 VTAIL.t1 5.22638
R71 VTAIL.n7 VTAIL.n6 1.61257
R72 VTAIL.n10 VTAIL.n9 1.61257
R73 VTAIL.n4 VTAIL.n2 1.61257
R74 VTAIL.n9 VTAIL.n7 1.27636
R75 VTAIL.n2 VTAIL.n1 1.27636
R76 VTAIL VTAIL.n11 1.15136
R77 VTAIL VTAIL.n1 0.461707
R78 VDD1 VDD1.t0 100.385
R79 VDD1.n1 VDD1.t3 100.27
R80 VDD1.n1 VDD1.n0 94.239
R81 VDD1.n3 VDD1.n2 93.8905
R82 VDD1.n3 VDD1.n1 35.7056
R83 VDD1.n2 VDD1.t4 5.22638
R84 VDD1.n2 VDD1.t5 5.22638
R85 VDD1.n0 VDD1.t1 5.22638
R86 VDD1.n0 VDD1.t2 5.22638
R87 VDD1 VDD1.n3 0.345328
R88 VN.n11 VN.n10 179.99
R89 VN.n23 VN.n22 179.99
R90 VN.n21 VN.n12 161.3
R91 VN.n20 VN.n19 161.3
R92 VN.n18 VN.n13 161.3
R93 VN.n17 VN.n16 161.3
R94 VN.n9 VN.n0 161.3
R95 VN.n8 VN.n7 161.3
R96 VN.n6 VN.n1 161.3
R97 VN.n5 VN.n4 161.3
R98 VN.n2 VN.t1 128.93
R99 VN.n14 VN.t2 128.93
R100 VN.n3 VN.t0 97.3395
R101 VN.n10 VN.t5 97.3395
R102 VN.n15 VN.t4 97.3395
R103 VN.n22 VN.t3 97.3395
R104 VN.n8 VN.n1 56.5617
R105 VN.n20 VN.n13 56.5617
R106 VN.n3 VN.n2 53.8793
R107 VN.n15 VN.n14 53.8793
R108 VN VN.n23 40.3925
R109 VN.n4 VN.n1 24.5923
R110 VN.n9 VN.n8 24.5923
R111 VN.n16 VN.n13 24.5923
R112 VN.n21 VN.n20 24.5923
R113 VN.n17 VN.n14 18.1684
R114 VN.n5 VN.n2 18.1684
R115 VN.n4 VN.n3 12.2964
R116 VN.n16 VN.n15 12.2964
R117 VN.n10 VN.n9 5.90254
R118 VN.n22 VN.n21 5.90254
R119 VN.n23 VN.n12 0.189894
R120 VN.n19 VN.n12 0.189894
R121 VN.n19 VN.n18 0.189894
R122 VN.n18 VN.n17 0.189894
R123 VN.n6 VN.n5 0.189894
R124 VN.n7 VN.n6 0.189894
R125 VN.n7 VN.n0 0.189894
R126 VN.n11 VN.n0 0.189894
R127 VN VN.n11 0.0516364
R128 VDD2.n1 VDD2.t4 100.27
R129 VDD2.n2 VDD2.t2 99.1174
R130 VDD2.n1 VDD2.n0 94.239
R131 VDD2 VDD2.n3 94.2353
R132 VDD2.n2 VDD2.n1 34.3166
R133 VDD2.n3 VDD2.t1 5.22638
R134 VDD2.n3 VDD2.t3 5.22638
R135 VDD2.n0 VDD2.t5 5.22638
R136 VDD2.n0 VDD2.t0 5.22638
R137 VDD2 VDD2.n2 1.26774
R138 B.n356 B.n355 585
R139 B.n357 B.n50 585
R140 B.n359 B.n358 585
R141 B.n360 B.n49 585
R142 B.n362 B.n361 585
R143 B.n363 B.n48 585
R144 B.n365 B.n364 585
R145 B.n366 B.n47 585
R146 B.n368 B.n367 585
R147 B.n369 B.n46 585
R148 B.n371 B.n370 585
R149 B.n372 B.n45 585
R150 B.n374 B.n373 585
R151 B.n375 B.n44 585
R152 B.n377 B.n376 585
R153 B.n378 B.n43 585
R154 B.n380 B.n379 585
R155 B.n381 B.n42 585
R156 B.n383 B.n382 585
R157 B.n384 B.n41 585
R158 B.n386 B.n385 585
R159 B.n387 B.n40 585
R160 B.n389 B.n388 585
R161 B.n390 B.n39 585
R162 B.n392 B.n391 585
R163 B.n394 B.n393 585
R164 B.n395 B.n35 585
R165 B.n397 B.n396 585
R166 B.n398 B.n34 585
R167 B.n400 B.n399 585
R168 B.n401 B.n33 585
R169 B.n403 B.n402 585
R170 B.n404 B.n32 585
R171 B.n406 B.n405 585
R172 B.n408 B.n29 585
R173 B.n410 B.n409 585
R174 B.n411 B.n28 585
R175 B.n413 B.n412 585
R176 B.n414 B.n27 585
R177 B.n416 B.n415 585
R178 B.n417 B.n26 585
R179 B.n419 B.n418 585
R180 B.n420 B.n25 585
R181 B.n422 B.n421 585
R182 B.n423 B.n24 585
R183 B.n425 B.n424 585
R184 B.n426 B.n23 585
R185 B.n428 B.n427 585
R186 B.n429 B.n22 585
R187 B.n431 B.n430 585
R188 B.n432 B.n21 585
R189 B.n434 B.n433 585
R190 B.n435 B.n20 585
R191 B.n437 B.n436 585
R192 B.n438 B.n19 585
R193 B.n440 B.n439 585
R194 B.n441 B.n18 585
R195 B.n443 B.n442 585
R196 B.n444 B.n17 585
R197 B.n354 B.n51 585
R198 B.n353 B.n352 585
R199 B.n351 B.n52 585
R200 B.n350 B.n349 585
R201 B.n348 B.n53 585
R202 B.n347 B.n346 585
R203 B.n345 B.n54 585
R204 B.n344 B.n343 585
R205 B.n342 B.n55 585
R206 B.n341 B.n340 585
R207 B.n339 B.n56 585
R208 B.n338 B.n337 585
R209 B.n336 B.n57 585
R210 B.n335 B.n334 585
R211 B.n333 B.n58 585
R212 B.n332 B.n331 585
R213 B.n330 B.n59 585
R214 B.n329 B.n328 585
R215 B.n327 B.n60 585
R216 B.n326 B.n325 585
R217 B.n324 B.n61 585
R218 B.n323 B.n322 585
R219 B.n321 B.n62 585
R220 B.n320 B.n319 585
R221 B.n318 B.n63 585
R222 B.n317 B.n316 585
R223 B.n315 B.n64 585
R224 B.n314 B.n313 585
R225 B.n312 B.n65 585
R226 B.n311 B.n310 585
R227 B.n309 B.n66 585
R228 B.n308 B.n307 585
R229 B.n306 B.n67 585
R230 B.n305 B.n304 585
R231 B.n303 B.n68 585
R232 B.n302 B.n301 585
R233 B.n300 B.n69 585
R234 B.n299 B.n298 585
R235 B.n297 B.n70 585
R236 B.n296 B.n295 585
R237 B.n294 B.n71 585
R238 B.n293 B.n292 585
R239 B.n291 B.n72 585
R240 B.n290 B.n289 585
R241 B.n288 B.n73 585
R242 B.n287 B.n286 585
R243 B.n285 B.n74 585
R244 B.n284 B.n283 585
R245 B.n282 B.n75 585
R246 B.n281 B.n280 585
R247 B.n279 B.n76 585
R248 B.n278 B.n277 585
R249 B.n276 B.n77 585
R250 B.n275 B.n274 585
R251 B.n273 B.n78 585
R252 B.n272 B.n271 585
R253 B.n270 B.n79 585
R254 B.n269 B.n268 585
R255 B.n267 B.n80 585
R256 B.n266 B.n265 585
R257 B.n264 B.n81 585
R258 B.n174 B.n115 585
R259 B.n176 B.n175 585
R260 B.n177 B.n114 585
R261 B.n179 B.n178 585
R262 B.n180 B.n113 585
R263 B.n182 B.n181 585
R264 B.n183 B.n112 585
R265 B.n185 B.n184 585
R266 B.n186 B.n111 585
R267 B.n188 B.n187 585
R268 B.n189 B.n110 585
R269 B.n191 B.n190 585
R270 B.n192 B.n109 585
R271 B.n194 B.n193 585
R272 B.n195 B.n108 585
R273 B.n197 B.n196 585
R274 B.n198 B.n107 585
R275 B.n200 B.n199 585
R276 B.n201 B.n106 585
R277 B.n203 B.n202 585
R278 B.n204 B.n105 585
R279 B.n206 B.n205 585
R280 B.n207 B.n104 585
R281 B.n209 B.n208 585
R282 B.n210 B.n101 585
R283 B.n213 B.n212 585
R284 B.n214 B.n100 585
R285 B.n216 B.n215 585
R286 B.n217 B.n99 585
R287 B.n219 B.n218 585
R288 B.n220 B.n98 585
R289 B.n222 B.n221 585
R290 B.n223 B.n97 585
R291 B.n225 B.n224 585
R292 B.n227 B.n226 585
R293 B.n228 B.n93 585
R294 B.n230 B.n229 585
R295 B.n231 B.n92 585
R296 B.n233 B.n232 585
R297 B.n234 B.n91 585
R298 B.n236 B.n235 585
R299 B.n237 B.n90 585
R300 B.n239 B.n238 585
R301 B.n240 B.n89 585
R302 B.n242 B.n241 585
R303 B.n243 B.n88 585
R304 B.n245 B.n244 585
R305 B.n246 B.n87 585
R306 B.n248 B.n247 585
R307 B.n249 B.n86 585
R308 B.n251 B.n250 585
R309 B.n252 B.n85 585
R310 B.n254 B.n253 585
R311 B.n255 B.n84 585
R312 B.n257 B.n256 585
R313 B.n258 B.n83 585
R314 B.n260 B.n259 585
R315 B.n261 B.n82 585
R316 B.n263 B.n262 585
R317 B.n173 B.n172 585
R318 B.n171 B.n116 585
R319 B.n170 B.n169 585
R320 B.n168 B.n117 585
R321 B.n167 B.n166 585
R322 B.n165 B.n118 585
R323 B.n164 B.n163 585
R324 B.n162 B.n119 585
R325 B.n161 B.n160 585
R326 B.n159 B.n120 585
R327 B.n158 B.n157 585
R328 B.n156 B.n121 585
R329 B.n155 B.n154 585
R330 B.n153 B.n122 585
R331 B.n152 B.n151 585
R332 B.n150 B.n123 585
R333 B.n149 B.n148 585
R334 B.n147 B.n124 585
R335 B.n146 B.n145 585
R336 B.n144 B.n125 585
R337 B.n143 B.n142 585
R338 B.n141 B.n126 585
R339 B.n140 B.n139 585
R340 B.n138 B.n127 585
R341 B.n137 B.n136 585
R342 B.n135 B.n128 585
R343 B.n134 B.n133 585
R344 B.n132 B.n129 585
R345 B.n131 B.n130 585
R346 B.n2 B.n0 585
R347 B.n489 B.n1 585
R348 B.n488 B.n487 585
R349 B.n486 B.n3 585
R350 B.n485 B.n484 585
R351 B.n483 B.n4 585
R352 B.n482 B.n481 585
R353 B.n480 B.n5 585
R354 B.n479 B.n478 585
R355 B.n477 B.n6 585
R356 B.n476 B.n475 585
R357 B.n474 B.n7 585
R358 B.n473 B.n472 585
R359 B.n471 B.n8 585
R360 B.n470 B.n469 585
R361 B.n468 B.n9 585
R362 B.n467 B.n466 585
R363 B.n465 B.n10 585
R364 B.n464 B.n463 585
R365 B.n462 B.n11 585
R366 B.n461 B.n460 585
R367 B.n459 B.n12 585
R368 B.n458 B.n457 585
R369 B.n456 B.n13 585
R370 B.n455 B.n454 585
R371 B.n453 B.n14 585
R372 B.n452 B.n451 585
R373 B.n450 B.n15 585
R374 B.n449 B.n448 585
R375 B.n447 B.n16 585
R376 B.n446 B.n445 585
R377 B.n491 B.n490 585
R378 B.n172 B.n115 502.111
R379 B.n446 B.n17 502.111
R380 B.n262 B.n81 502.111
R381 B.n356 B.n51 502.111
R382 B.n94 B.t9 302.925
R383 B.n102 B.t6 302.925
R384 B.n30 B.t3 302.925
R385 B.n36 B.t0 302.925
R386 B.n172 B.n171 163.367
R387 B.n171 B.n170 163.367
R388 B.n170 B.n117 163.367
R389 B.n166 B.n117 163.367
R390 B.n166 B.n165 163.367
R391 B.n165 B.n164 163.367
R392 B.n164 B.n119 163.367
R393 B.n160 B.n119 163.367
R394 B.n160 B.n159 163.367
R395 B.n159 B.n158 163.367
R396 B.n158 B.n121 163.367
R397 B.n154 B.n121 163.367
R398 B.n154 B.n153 163.367
R399 B.n153 B.n152 163.367
R400 B.n152 B.n123 163.367
R401 B.n148 B.n123 163.367
R402 B.n148 B.n147 163.367
R403 B.n147 B.n146 163.367
R404 B.n146 B.n125 163.367
R405 B.n142 B.n125 163.367
R406 B.n142 B.n141 163.367
R407 B.n141 B.n140 163.367
R408 B.n140 B.n127 163.367
R409 B.n136 B.n127 163.367
R410 B.n136 B.n135 163.367
R411 B.n135 B.n134 163.367
R412 B.n134 B.n129 163.367
R413 B.n130 B.n129 163.367
R414 B.n130 B.n2 163.367
R415 B.n490 B.n2 163.367
R416 B.n490 B.n489 163.367
R417 B.n489 B.n488 163.367
R418 B.n488 B.n3 163.367
R419 B.n484 B.n3 163.367
R420 B.n484 B.n483 163.367
R421 B.n483 B.n482 163.367
R422 B.n482 B.n5 163.367
R423 B.n478 B.n5 163.367
R424 B.n478 B.n477 163.367
R425 B.n477 B.n476 163.367
R426 B.n476 B.n7 163.367
R427 B.n472 B.n7 163.367
R428 B.n472 B.n471 163.367
R429 B.n471 B.n470 163.367
R430 B.n470 B.n9 163.367
R431 B.n466 B.n9 163.367
R432 B.n466 B.n465 163.367
R433 B.n465 B.n464 163.367
R434 B.n464 B.n11 163.367
R435 B.n460 B.n11 163.367
R436 B.n460 B.n459 163.367
R437 B.n459 B.n458 163.367
R438 B.n458 B.n13 163.367
R439 B.n454 B.n13 163.367
R440 B.n454 B.n453 163.367
R441 B.n453 B.n452 163.367
R442 B.n452 B.n15 163.367
R443 B.n448 B.n15 163.367
R444 B.n448 B.n447 163.367
R445 B.n447 B.n446 163.367
R446 B.n176 B.n115 163.367
R447 B.n177 B.n176 163.367
R448 B.n178 B.n177 163.367
R449 B.n178 B.n113 163.367
R450 B.n182 B.n113 163.367
R451 B.n183 B.n182 163.367
R452 B.n184 B.n183 163.367
R453 B.n184 B.n111 163.367
R454 B.n188 B.n111 163.367
R455 B.n189 B.n188 163.367
R456 B.n190 B.n189 163.367
R457 B.n190 B.n109 163.367
R458 B.n194 B.n109 163.367
R459 B.n195 B.n194 163.367
R460 B.n196 B.n195 163.367
R461 B.n196 B.n107 163.367
R462 B.n200 B.n107 163.367
R463 B.n201 B.n200 163.367
R464 B.n202 B.n201 163.367
R465 B.n202 B.n105 163.367
R466 B.n206 B.n105 163.367
R467 B.n207 B.n206 163.367
R468 B.n208 B.n207 163.367
R469 B.n208 B.n101 163.367
R470 B.n213 B.n101 163.367
R471 B.n214 B.n213 163.367
R472 B.n215 B.n214 163.367
R473 B.n215 B.n99 163.367
R474 B.n219 B.n99 163.367
R475 B.n220 B.n219 163.367
R476 B.n221 B.n220 163.367
R477 B.n221 B.n97 163.367
R478 B.n225 B.n97 163.367
R479 B.n226 B.n225 163.367
R480 B.n226 B.n93 163.367
R481 B.n230 B.n93 163.367
R482 B.n231 B.n230 163.367
R483 B.n232 B.n231 163.367
R484 B.n232 B.n91 163.367
R485 B.n236 B.n91 163.367
R486 B.n237 B.n236 163.367
R487 B.n238 B.n237 163.367
R488 B.n238 B.n89 163.367
R489 B.n242 B.n89 163.367
R490 B.n243 B.n242 163.367
R491 B.n244 B.n243 163.367
R492 B.n244 B.n87 163.367
R493 B.n248 B.n87 163.367
R494 B.n249 B.n248 163.367
R495 B.n250 B.n249 163.367
R496 B.n250 B.n85 163.367
R497 B.n254 B.n85 163.367
R498 B.n255 B.n254 163.367
R499 B.n256 B.n255 163.367
R500 B.n256 B.n83 163.367
R501 B.n260 B.n83 163.367
R502 B.n261 B.n260 163.367
R503 B.n262 B.n261 163.367
R504 B.n266 B.n81 163.367
R505 B.n267 B.n266 163.367
R506 B.n268 B.n267 163.367
R507 B.n268 B.n79 163.367
R508 B.n272 B.n79 163.367
R509 B.n273 B.n272 163.367
R510 B.n274 B.n273 163.367
R511 B.n274 B.n77 163.367
R512 B.n278 B.n77 163.367
R513 B.n279 B.n278 163.367
R514 B.n280 B.n279 163.367
R515 B.n280 B.n75 163.367
R516 B.n284 B.n75 163.367
R517 B.n285 B.n284 163.367
R518 B.n286 B.n285 163.367
R519 B.n286 B.n73 163.367
R520 B.n290 B.n73 163.367
R521 B.n291 B.n290 163.367
R522 B.n292 B.n291 163.367
R523 B.n292 B.n71 163.367
R524 B.n296 B.n71 163.367
R525 B.n297 B.n296 163.367
R526 B.n298 B.n297 163.367
R527 B.n298 B.n69 163.367
R528 B.n302 B.n69 163.367
R529 B.n303 B.n302 163.367
R530 B.n304 B.n303 163.367
R531 B.n304 B.n67 163.367
R532 B.n308 B.n67 163.367
R533 B.n309 B.n308 163.367
R534 B.n310 B.n309 163.367
R535 B.n310 B.n65 163.367
R536 B.n314 B.n65 163.367
R537 B.n315 B.n314 163.367
R538 B.n316 B.n315 163.367
R539 B.n316 B.n63 163.367
R540 B.n320 B.n63 163.367
R541 B.n321 B.n320 163.367
R542 B.n322 B.n321 163.367
R543 B.n322 B.n61 163.367
R544 B.n326 B.n61 163.367
R545 B.n327 B.n326 163.367
R546 B.n328 B.n327 163.367
R547 B.n328 B.n59 163.367
R548 B.n332 B.n59 163.367
R549 B.n333 B.n332 163.367
R550 B.n334 B.n333 163.367
R551 B.n334 B.n57 163.367
R552 B.n338 B.n57 163.367
R553 B.n339 B.n338 163.367
R554 B.n340 B.n339 163.367
R555 B.n340 B.n55 163.367
R556 B.n344 B.n55 163.367
R557 B.n345 B.n344 163.367
R558 B.n346 B.n345 163.367
R559 B.n346 B.n53 163.367
R560 B.n350 B.n53 163.367
R561 B.n351 B.n350 163.367
R562 B.n352 B.n351 163.367
R563 B.n352 B.n51 163.367
R564 B.n442 B.n17 163.367
R565 B.n442 B.n441 163.367
R566 B.n441 B.n440 163.367
R567 B.n440 B.n19 163.367
R568 B.n436 B.n19 163.367
R569 B.n436 B.n435 163.367
R570 B.n435 B.n434 163.367
R571 B.n434 B.n21 163.367
R572 B.n430 B.n21 163.367
R573 B.n430 B.n429 163.367
R574 B.n429 B.n428 163.367
R575 B.n428 B.n23 163.367
R576 B.n424 B.n23 163.367
R577 B.n424 B.n423 163.367
R578 B.n423 B.n422 163.367
R579 B.n422 B.n25 163.367
R580 B.n418 B.n25 163.367
R581 B.n418 B.n417 163.367
R582 B.n417 B.n416 163.367
R583 B.n416 B.n27 163.367
R584 B.n412 B.n27 163.367
R585 B.n412 B.n411 163.367
R586 B.n411 B.n410 163.367
R587 B.n410 B.n29 163.367
R588 B.n405 B.n29 163.367
R589 B.n405 B.n404 163.367
R590 B.n404 B.n403 163.367
R591 B.n403 B.n33 163.367
R592 B.n399 B.n33 163.367
R593 B.n399 B.n398 163.367
R594 B.n398 B.n397 163.367
R595 B.n397 B.n35 163.367
R596 B.n393 B.n35 163.367
R597 B.n393 B.n392 163.367
R598 B.n392 B.n39 163.367
R599 B.n388 B.n39 163.367
R600 B.n388 B.n387 163.367
R601 B.n387 B.n386 163.367
R602 B.n386 B.n41 163.367
R603 B.n382 B.n41 163.367
R604 B.n382 B.n381 163.367
R605 B.n381 B.n380 163.367
R606 B.n380 B.n43 163.367
R607 B.n376 B.n43 163.367
R608 B.n376 B.n375 163.367
R609 B.n375 B.n374 163.367
R610 B.n374 B.n45 163.367
R611 B.n370 B.n45 163.367
R612 B.n370 B.n369 163.367
R613 B.n369 B.n368 163.367
R614 B.n368 B.n47 163.367
R615 B.n364 B.n47 163.367
R616 B.n364 B.n363 163.367
R617 B.n363 B.n362 163.367
R618 B.n362 B.n49 163.367
R619 B.n358 B.n49 163.367
R620 B.n358 B.n357 163.367
R621 B.n357 B.n356 163.367
R622 B.n94 B.t11 148.893
R623 B.n36 B.t1 148.893
R624 B.n102 B.t8 148.887
R625 B.n30 B.t4 148.887
R626 B.n95 B.t10 112.626
R627 B.n37 B.t2 112.626
R628 B.n103 B.t7 112.621
R629 B.n31 B.t5 112.621
R630 B.n96 B.n95 59.5399
R631 B.n211 B.n103 59.5399
R632 B.n407 B.n31 59.5399
R633 B.n38 B.n37 59.5399
R634 B.n95 B.n94 36.2672
R635 B.n103 B.n102 36.2672
R636 B.n31 B.n30 36.2672
R637 B.n37 B.n36 36.2672
R638 B.n445 B.n444 32.6249
R639 B.n355 B.n354 32.6249
R640 B.n264 B.n263 32.6249
R641 B.n174 B.n173 32.6249
R642 B B.n491 18.0485
R643 B.n444 B.n443 10.6151
R644 B.n443 B.n18 10.6151
R645 B.n439 B.n18 10.6151
R646 B.n439 B.n438 10.6151
R647 B.n438 B.n437 10.6151
R648 B.n437 B.n20 10.6151
R649 B.n433 B.n20 10.6151
R650 B.n433 B.n432 10.6151
R651 B.n432 B.n431 10.6151
R652 B.n431 B.n22 10.6151
R653 B.n427 B.n22 10.6151
R654 B.n427 B.n426 10.6151
R655 B.n426 B.n425 10.6151
R656 B.n425 B.n24 10.6151
R657 B.n421 B.n24 10.6151
R658 B.n421 B.n420 10.6151
R659 B.n420 B.n419 10.6151
R660 B.n419 B.n26 10.6151
R661 B.n415 B.n26 10.6151
R662 B.n415 B.n414 10.6151
R663 B.n414 B.n413 10.6151
R664 B.n413 B.n28 10.6151
R665 B.n409 B.n28 10.6151
R666 B.n409 B.n408 10.6151
R667 B.n406 B.n32 10.6151
R668 B.n402 B.n32 10.6151
R669 B.n402 B.n401 10.6151
R670 B.n401 B.n400 10.6151
R671 B.n400 B.n34 10.6151
R672 B.n396 B.n34 10.6151
R673 B.n396 B.n395 10.6151
R674 B.n395 B.n394 10.6151
R675 B.n391 B.n390 10.6151
R676 B.n390 B.n389 10.6151
R677 B.n389 B.n40 10.6151
R678 B.n385 B.n40 10.6151
R679 B.n385 B.n384 10.6151
R680 B.n384 B.n383 10.6151
R681 B.n383 B.n42 10.6151
R682 B.n379 B.n42 10.6151
R683 B.n379 B.n378 10.6151
R684 B.n378 B.n377 10.6151
R685 B.n377 B.n44 10.6151
R686 B.n373 B.n44 10.6151
R687 B.n373 B.n372 10.6151
R688 B.n372 B.n371 10.6151
R689 B.n371 B.n46 10.6151
R690 B.n367 B.n46 10.6151
R691 B.n367 B.n366 10.6151
R692 B.n366 B.n365 10.6151
R693 B.n365 B.n48 10.6151
R694 B.n361 B.n48 10.6151
R695 B.n361 B.n360 10.6151
R696 B.n360 B.n359 10.6151
R697 B.n359 B.n50 10.6151
R698 B.n355 B.n50 10.6151
R699 B.n265 B.n264 10.6151
R700 B.n265 B.n80 10.6151
R701 B.n269 B.n80 10.6151
R702 B.n270 B.n269 10.6151
R703 B.n271 B.n270 10.6151
R704 B.n271 B.n78 10.6151
R705 B.n275 B.n78 10.6151
R706 B.n276 B.n275 10.6151
R707 B.n277 B.n276 10.6151
R708 B.n277 B.n76 10.6151
R709 B.n281 B.n76 10.6151
R710 B.n282 B.n281 10.6151
R711 B.n283 B.n282 10.6151
R712 B.n283 B.n74 10.6151
R713 B.n287 B.n74 10.6151
R714 B.n288 B.n287 10.6151
R715 B.n289 B.n288 10.6151
R716 B.n289 B.n72 10.6151
R717 B.n293 B.n72 10.6151
R718 B.n294 B.n293 10.6151
R719 B.n295 B.n294 10.6151
R720 B.n295 B.n70 10.6151
R721 B.n299 B.n70 10.6151
R722 B.n300 B.n299 10.6151
R723 B.n301 B.n300 10.6151
R724 B.n301 B.n68 10.6151
R725 B.n305 B.n68 10.6151
R726 B.n306 B.n305 10.6151
R727 B.n307 B.n306 10.6151
R728 B.n307 B.n66 10.6151
R729 B.n311 B.n66 10.6151
R730 B.n312 B.n311 10.6151
R731 B.n313 B.n312 10.6151
R732 B.n313 B.n64 10.6151
R733 B.n317 B.n64 10.6151
R734 B.n318 B.n317 10.6151
R735 B.n319 B.n318 10.6151
R736 B.n319 B.n62 10.6151
R737 B.n323 B.n62 10.6151
R738 B.n324 B.n323 10.6151
R739 B.n325 B.n324 10.6151
R740 B.n325 B.n60 10.6151
R741 B.n329 B.n60 10.6151
R742 B.n330 B.n329 10.6151
R743 B.n331 B.n330 10.6151
R744 B.n331 B.n58 10.6151
R745 B.n335 B.n58 10.6151
R746 B.n336 B.n335 10.6151
R747 B.n337 B.n336 10.6151
R748 B.n337 B.n56 10.6151
R749 B.n341 B.n56 10.6151
R750 B.n342 B.n341 10.6151
R751 B.n343 B.n342 10.6151
R752 B.n343 B.n54 10.6151
R753 B.n347 B.n54 10.6151
R754 B.n348 B.n347 10.6151
R755 B.n349 B.n348 10.6151
R756 B.n349 B.n52 10.6151
R757 B.n353 B.n52 10.6151
R758 B.n354 B.n353 10.6151
R759 B.n175 B.n174 10.6151
R760 B.n175 B.n114 10.6151
R761 B.n179 B.n114 10.6151
R762 B.n180 B.n179 10.6151
R763 B.n181 B.n180 10.6151
R764 B.n181 B.n112 10.6151
R765 B.n185 B.n112 10.6151
R766 B.n186 B.n185 10.6151
R767 B.n187 B.n186 10.6151
R768 B.n187 B.n110 10.6151
R769 B.n191 B.n110 10.6151
R770 B.n192 B.n191 10.6151
R771 B.n193 B.n192 10.6151
R772 B.n193 B.n108 10.6151
R773 B.n197 B.n108 10.6151
R774 B.n198 B.n197 10.6151
R775 B.n199 B.n198 10.6151
R776 B.n199 B.n106 10.6151
R777 B.n203 B.n106 10.6151
R778 B.n204 B.n203 10.6151
R779 B.n205 B.n204 10.6151
R780 B.n205 B.n104 10.6151
R781 B.n209 B.n104 10.6151
R782 B.n210 B.n209 10.6151
R783 B.n212 B.n100 10.6151
R784 B.n216 B.n100 10.6151
R785 B.n217 B.n216 10.6151
R786 B.n218 B.n217 10.6151
R787 B.n218 B.n98 10.6151
R788 B.n222 B.n98 10.6151
R789 B.n223 B.n222 10.6151
R790 B.n224 B.n223 10.6151
R791 B.n228 B.n227 10.6151
R792 B.n229 B.n228 10.6151
R793 B.n229 B.n92 10.6151
R794 B.n233 B.n92 10.6151
R795 B.n234 B.n233 10.6151
R796 B.n235 B.n234 10.6151
R797 B.n235 B.n90 10.6151
R798 B.n239 B.n90 10.6151
R799 B.n240 B.n239 10.6151
R800 B.n241 B.n240 10.6151
R801 B.n241 B.n88 10.6151
R802 B.n245 B.n88 10.6151
R803 B.n246 B.n245 10.6151
R804 B.n247 B.n246 10.6151
R805 B.n247 B.n86 10.6151
R806 B.n251 B.n86 10.6151
R807 B.n252 B.n251 10.6151
R808 B.n253 B.n252 10.6151
R809 B.n253 B.n84 10.6151
R810 B.n257 B.n84 10.6151
R811 B.n258 B.n257 10.6151
R812 B.n259 B.n258 10.6151
R813 B.n259 B.n82 10.6151
R814 B.n263 B.n82 10.6151
R815 B.n173 B.n116 10.6151
R816 B.n169 B.n116 10.6151
R817 B.n169 B.n168 10.6151
R818 B.n168 B.n167 10.6151
R819 B.n167 B.n118 10.6151
R820 B.n163 B.n118 10.6151
R821 B.n163 B.n162 10.6151
R822 B.n162 B.n161 10.6151
R823 B.n161 B.n120 10.6151
R824 B.n157 B.n120 10.6151
R825 B.n157 B.n156 10.6151
R826 B.n156 B.n155 10.6151
R827 B.n155 B.n122 10.6151
R828 B.n151 B.n122 10.6151
R829 B.n151 B.n150 10.6151
R830 B.n150 B.n149 10.6151
R831 B.n149 B.n124 10.6151
R832 B.n145 B.n124 10.6151
R833 B.n145 B.n144 10.6151
R834 B.n144 B.n143 10.6151
R835 B.n143 B.n126 10.6151
R836 B.n139 B.n126 10.6151
R837 B.n139 B.n138 10.6151
R838 B.n138 B.n137 10.6151
R839 B.n137 B.n128 10.6151
R840 B.n133 B.n128 10.6151
R841 B.n133 B.n132 10.6151
R842 B.n132 B.n131 10.6151
R843 B.n131 B.n0 10.6151
R844 B.n487 B.n1 10.6151
R845 B.n487 B.n486 10.6151
R846 B.n486 B.n485 10.6151
R847 B.n485 B.n4 10.6151
R848 B.n481 B.n4 10.6151
R849 B.n481 B.n480 10.6151
R850 B.n480 B.n479 10.6151
R851 B.n479 B.n6 10.6151
R852 B.n475 B.n6 10.6151
R853 B.n475 B.n474 10.6151
R854 B.n474 B.n473 10.6151
R855 B.n473 B.n8 10.6151
R856 B.n469 B.n8 10.6151
R857 B.n469 B.n468 10.6151
R858 B.n468 B.n467 10.6151
R859 B.n467 B.n10 10.6151
R860 B.n463 B.n10 10.6151
R861 B.n463 B.n462 10.6151
R862 B.n462 B.n461 10.6151
R863 B.n461 B.n12 10.6151
R864 B.n457 B.n12 10.6151
R865 B.n457 B.n456 10.6151
R866 B.n456 B.n455 10.6151
R867 B.n455 B.n14 10.6151
R868 B.n451 B.n14 10.6151
R869 B.n451 B.n450 10.6151
R870 B.n450 B.n449 10.6151
R871 B.n449 B.n16 10.6151
R872 B.n445 B.n16 10.6151
R873 B.n407 B.n406 6.5566
R874 B.n394 B.n38 6.5566
R875 B.n212 B.n211 6.5566
R876 B.n224 B.n96 6.5566
R877 B.n408 B.n407 4.05904
R878 B.n391 B.n38 4.05904
R879 B.n211 B.n210 4.05904
R880 B.n227 B.n96 4.05904
R881 B.n491 B.n0 2.81026
R882 B.n491 B.n1 2.81026
C0 VDD2 VN 3.24516f
C1 VTAIL VN 3.48609f
C2 VDD2 VP 0.368322f
C3 VDD1 VN 0.14969f
C4 VTAIL VP 3.50035f
C5 VDD1 VP 3.46156f
C6 w_n2466_n2212# VDD2 1.67008f
C7 w_n2466_n2212# VTAIL 2.06196f
C8 w_n2466_n2212# VDD1 1.61909f
C9 VN B 0.875507f
C10 VP B 1.39754f
C11 VTAIL VDD2 5.38763f
C12 VDD1 VDD2 1.02165f
C13 w_n2466_n2212# B 6.59717f
C14 VTAIL VDD1 5.34341f
C15 VP VN 4.8244f
C16 VDD2 B 1.41362f
C17 VTAIL B 2.02582f
C18 VDD1 B 1.36484f
C19 w_n2466_n2212# VN 4.30519f
C20 w_n2466_n2212# VP 4.62105f
C21 VDD2 VSUBS 1.190777f
C22 VDD1 VSUBS 1.55942f
C23 VTAIL VSUBS 0.571721f
C24 VN VSUBS 4.544361f
C25 VP VSUBS 1.780393f
C26 B VSUBS 3.101338f
C27 w_n2466_n2212# VSUBS 68.032f
C28 B.n0 VSUBS 0.005051f
C29 B.n1 VSUBS 0.005051f
C30 B.n2 VSUBS 0.007987f
C31 B.n3 VSUBS 0.007987f
C32 B.n4 VSUBS 0.007987f
C33 B.n5 VSUBS 0.007987f
C34 B.n6 VSUBS 0.007987f
C35 B.n7 VSUBS 0.007987f
C36 B.n8 VSUBS 0.007987f
C37 B.n9 VSUBS 0.007987f
C38 B.n10 VSUBS 0.007987f
C39 B.n11 VSUBS 0.007987f
C40 B.n12 VSUBS 0.007987f
C41 B.n13 VSUBS 0.007987f
C42 B.n14 VSUBS 0.007987f
C43 B.n15 VSUBS 0.007987f
C44 B.n16 VSUBS 0.007987f
C45 B.n17 VSUBS 0.019286f
C46 B.n18 VSUBS 0.007987f
C47 B.n19 VSUBS 0.007987f
C48 B.n20 VSUBS 0.007987f
C49 B.n21 VSUBS 0.007987f
C50 B.n22 VSUBS 0.007987f
C51 B.n23 VSUBS 0.007987f
C52 B.n24 VSUBS 0.007987f
C53 B.n25 VSUBS 0.007987f
C54 B.n26 VSUBS 0.007987f
C55 B.n27 VSUBS 0.007987f
C56 B.n28 VSUBS 0.007987f
C57 B.n29 VSUBS 0.007987f
C58 B.t5 VSUBS 0.208807f
C59 B.t4 VSUBS 0.224512f
C60 B.t3 VSUBS 0.500543f
C61 B.n30 VSUBS 0.120973f
C62 B.n31 VSUBS 0.075866f
C63 B.n32 VSUBS 0.007987f
C64 B.n33 VSUBS 0.007987f
C65 B.n34 VSUBS 0.007987f
C66 B.n35 VSUBS 0.007987f
C67 B.t2 VSUBS 0.208806f
C68 B.t1 VSUBS 0.224511f
C69 B.t0 VSUBS 0.500543f
C70 B.n36 VSUBS 0.120974f
C71 B.n37 VSUBS 0.075867f
C72 B.n38 VSUBS 0.018505f
C73 B.n39 VSUBS 0.007987f
C74 B.n40 VSUBS 0.007987f
C75 B.n41 VSUBS 0.007987f
C76 B.n42 VSUBS 0.007987f
C77 B.n43 VSUBS 0.007987f
C78 B.n44 VSUBS 0.007987f
C79 B.n45 VSUBS 0.007987f
C80 B.n46 VSUBS 0.007987f
C81 B.n47 VSUBS 0.007987f
C82 B.n48 VSUBS 0.007987f
C83 B.n49 VSUBS 0.007987f
C84 B.n50 VSUBS 0.007987f
C85 B.n51 VSUBS 0.018065f
C86 B.n52 VSUBS 0.007987f
C87 B.n53 VSUBS 0.007987f
C88 B.n54 VSUBS 0.007987f
C89 B.n55 VSUBS 0.007987f
C90 B.n56 VSUBS 0.007987f
C91 B.n57 VSUBS 0.007987f
C92 B.n58 VSUBS 0.007987f
C93 B.n59 VSUBS 0.007987f
C94 B.n60 VSUBS 0.007987f
C95 B.n61 VSUBS 0.007987f
C96 B.n62 VSUBS 0.007987f
C97 B.n63 VSUBS 0.007987f
C98 B.n64 VSUBS 0.007987f
C99 B.n65 VSUBS 0.007987f
C100 B.n66 VSUBS 0.007987f
C101 B.n67 VSUBS 0.007987f
C102 B.n68 VSUBS 0.007987f
C103 B.n69 VSUBS 0.007987f
C104 B.n70 VSUBS 0.007987f
C105 B.n71 VSUBS 0.007987f
C106 B.n72 VSUBS 0.007987f
C107 B.n73 VSUBS 0.007987f
C108 B.n74 VSUBS 0.007987f
C109 B.n75 VSUBS 0.007987f
C110 B.n76 VSUBS 0.007987f
C111 B.n77 VSUBS 0.007987f
C112 B.n78 VSUBS 0.007987f
C113 B.n79 VSUBS 0.007987f
C114 B.n80 VSUBS 0.007987f
C115 B.n81 VSUBS 0.018065f
C116 B.n82 VSUBS 0.007987f
C117 B.n83 VSUBS 0.007987f
C118 B.n84 VSUBS 0.007987f
C119 B.n85 VSUBS 0.007987f
C120 B.n86 VSUBS 0.007987f
C121 B.n87 VSUBS 0.007987f
C122 B.n88 VSUBS 0.007987f
C123 B.n89 VSUBS 0.007987f
C124 B.n90 VSUBS 0.007987f
C125 B.n91 VSUBS 0.007987f
C126 B.n92 VSUBS 0.007987f
C127 B.n93 VSUBS 0.007987f
C128 B.t10 VSUBS 0.208806f
C129 B.t11 VSUBS 0.224511f
C130 B.t9 VSUBS 0.500543f
C131 B.n94 VSUBS 0.120974f
C132 B.n95 VSUBS 0.075867f
C133 B.n96 VSUBS 0.018505f
C134 B.n97 VSUBS 0.007987f
C135 B.n98 VSUBS 0.007987f
C136 B.n99 VSUBS 0.007987f
C137 B.n100 VSUBS 0.007987f
C138 B.n101 VSUBS 0.007987f
C139 B.t7 VSUBS 0.208807f
C140 B.t8 VSUBS 0.224512f
C141 B.t6 VSUBS 0.500543f
C142 B.n102 VSUBS 0.120973f
C143 B.n103 VSUBS 0.075866f
C144 B.n104 VSUBS 0.007987f
C145 B.n105 VSUBS 0.007987f
C146 B.n106 VSUBS 0.007987f
C147 B.n107 VSUBS 0.007987f
C148 B.n108 VSUBS 0.007987f
C149 B.n109 VSUBS 0.007987f
C150 B.n110 VSUBS 0.007987f
C151 B.n111 VSUBS 0.007987f
C152 B.n112 VSUBS 0.007987f
C153 B.n113 VSUBS 0.007987f
C154 B.n114 VSUBS 0.007987f
C155 B.n115 VSUBS 0.019286f
C156 B.n116 VSUBS 0.007987f
C157 B.n117 VSUBS 0.007987f
C158 B.n118 VSUBS 0.007987f
C159 B.n119 VSUBS 0.007987f
C160 B.n120 VSUBS 0.007987f
C161 B.n121 VSUBS 0.007987f
C162 B.n122 VSUBS 0.007987f
C163 B.n123 VSUBS 0.007987f
C164 B.n124 VSUBS 0.007987f
C165 B.n125 VSUBS 0.007987f
C166 B.n126 VSUBS 0.007987f
C167 B.n127 VSUBS 0.007987f
C168 B.n128 VSUBS 0.007987f
C169 B.n129 VSUBS 0.007987f
C170 B.n130 VSUBS 0.007987f
C171 B.n131 VSUBS 0.007987f
C172 B.n132 VSUBS 0.007987f
C173 B.n133 VSUBS 0.007987f
C174 B.n134 VSUBS 0.007987f
C175 B.n135 VSUBS 0.007987f
C176 B.n136 VSUBS 0.007987f
C177 B.n137 VSUBS 0.007987f
C178 B.n138 VSUBS 0.007987f
C179 B.n139 VSUBS 0.007987f
C180 B.n140 VSUBS 0.007987f
C181 B.n141 VSUBS 0.007987f
C182 B.n142 VSUBS 0.007987f
C183 B.n143 VSUBS 0.007987f
C184 B.n144 VSUBS 0.007987f
C185 B.n145 VSUBS 0.007987f
C186 B.n146 VSUBS 0.007987f
C187 B.n147 VSUBS 0.007987f
C188 B.n148 VSUBS 0.007987f
C189 B.n149 VSUBS 0.007987f
C190 B.n150 VSUBS 0.007987f
C191 B.n151 VSUBS 0.007987f
C192 B.n152 VSUBS 0.007987f
C193 B.n153 VSUBS 0.007987f
C194 B.n154 VSUBS 0.007987f
C195 B.n155 VSUBS 0.007987f
C196 B.n156 VSUBS 0.007987f
C197 B.n157 VSUBS 0.007987f
C198 B.n158 VSUBS 0.007987f
C199 B.n159 VSUBS 0.007987f
C200 B.n160 VSUBS 0.007987f
C201 B.n161 VSUBS 0.007987f
C202 B.n162 VSUBS 0.007987f
C203 B.n163 VSUBS 0.007987f
C204 B.n164 VSUBS 0.007987f
C205 B.n165 VSUBS 0.007987f
C206 B.n166 VSUBS 0.007987f
C207 B.n167 VSUBS 0.007987f
C208 B.n168 VSUBS 0.007987f
C209 B.n169 VSUBS 0.007987f
C210 B.n170 VSUBS 0.007987f
C211 B.n171 VSUBS 0.007987f
C212 B.n172 VSUBS 0.018065f
C213 B.n173 VSUBS 0.018065f
C214 B.n174 VSUBS 0.019286f
C215 B.n175 VSUBS 0.007987f
C216 B.n176 VSUBS 0.007987f
C217 B.n177 VSUBS 0.007987f
C218 B.n178 VSUBS 0.007987f
C219 B.n179 VSUBS 0.007987f
C220 B.n180 VSUBS 0.007987f
C221 B.n181 VSUBS 0.007987f
C222 B.n182 VSUBS 0.007987f
C223 B.n183 VSUBS 0.007987f
C224 B.n184 VSUBS 0.007987f
C225 B.n185 VSUBS 0.007987f
C226 B.n186 VSUBS 0.007987f
C227 B.n187 VSUBS 0.007987f
C228 B.n188 VSUBS 0.007987f
C229 B.n189 VSUBS 0.007987f
C230 B.n190 VSUBS 0.007987f
C231 B.n191 VSUBS 0.007987f
C232 B.n192 VSUBS 0.007987f
C233 B.n193 VSUBS 0.007987f
C234 B.n194 VSUBS 0.007987f
C235 B.n195 VSUBS 0.007987f
C236 B.n196 VSUBS 0.007987f
C237 B.n197 VSUBS 0.007987f
C238 B.n198 VSUBS 0.007987f
C239 B.n199 VSUBS 0.007987f
C240 B.n200 VSUBS 0.007987f
C241 B.n201 VSUBS 0.007987f
C242 B.n202 VSUBS 0.007987f
C243 B.n203 VSUBS 0.007987f
C244 B.n204 VSUBS 0.007987f
C245 B.n205 VSUBS 0.007987f
C246 B.n206 VSUBS 0.007987f
C247 B.n207 VSUBS 0.007987f
C248 B.n208 VSUBS 0.007987f
C249 B.n209 VSUBS 0.007987f
C250 B.n210 VSUBS 0.00552f
C251 B.n211 VSUBS 0.018505f
C252 B.n212 VSUBS 0.00646f
C253 B.n213 VSUBS 0.007987f
C254 B.n214 VSUBS 0.007987f
C255 B.n215 VSUBS 0.007987f
C256 B.n216 VSUBS 0.007987f
C257 B.n217 VSUBS 0.007987f
C258 B.n218 VSUBS 0.007987f
C259 B.n219 VSUBS 0.007987f
C260 B.n220 VSUBS 0.007987f
C261 B.n221 VSUBS 0.007987f
C262 B.n222 VSUBS 0.007987f
C263 B.n223 VSUBS 0.007987f
C264 B.n224 VSUBS 0.00646f
C265 B.n225 VSUBS 0.007987f
C266 B.n226 VSUBS 0.007987f
C267 B.n227 VSUBS 0.00552f
C268 B.n228 VSUBS 0.007987f
C269 B.n229 VSUBS 0.007987f
C270 B.n230 VSUBS 0.007987f
C271 B.n231 VSUBS 0.007987f
C272 B.n232 VSUBS 0.007987f
C273 B.n233 VSUBS 0.007987f
C274 B.n234 VSUBS 0.007987f
C275 B.n235 VSUBS 0.007987f
C276 B.n236 VSUBS 0.007987f
C277 B.n237 VSUBS 0.007987f
C278 B.n238 VSUBS 0.007987f
C279 B.n239 VSUBS 0.007987f
C280 B.n240 VSUBS 0.007987f
C281 B.n241 VSUBS 0.007987f
C282 B.n242 VSUBS 0.007987f
C283 B.n243 VSUBS 0.007987f
C284 B.n244 VSUBS 0.007987f
C285 B.n245 VSUBS 0.007987f
C286 B.n246 VSUBS 0.007987f
C287 B.n247 VSUBS 0.007987f
C288 B.n248 VSUBS 0.007987f
C289 B.n249 VSUBS 0.007987f
C290 B.n250 VSUBS 0.007987f
C291 B.n251 VSUBS 0.007987f
C292 B.n252 VSUBS 0.007987f
C293 B.n253 VSUBS 0.007987f
C294 B.n254 VSUBS 0.007987f
C295 B.n255 VSUBS 0.007987f
C296 B.n256 VSUBS 0.007987f
C297 B.n257 VSUBS 0.007987f
C298 B.n258 VSUBS 0.007987f
C299 B.n259 VSUBS 0.007987f
C300 B.n260 VSUBS 0.007987f
C301 B.n261 VSUBS 0.007987f
C302 B.n262 VSUBS 0.019286f
C303 B.n263 VSUBS 0.019286f
C304 B.n264 VSUBS 0.018065f
C305 B.n265 VSUBS 0.007987f
C306 B.n266 VSUBS 0.007987f
C307 B.n267 VSUBS 0.007987f
C308 B.n268 VSUBS 0.007987f
C309 B.n269 VSUBS 0.007987f
C310 B.n270 VSUBS 0.007987f
C311 B.n271 VSUBS 0.007987f
C312 B.n272 VSUBS 0.007987f
C313 B.n273 VSUBS 0.007987f
C314 B.n274 VSUBS 0.007987f
C315 B.n275 VSUBS 0.007987f
C316 B.n276 VSUBS 0.007987f
C317 B.n277 VSUBS 0.007987f
C318 B.n278 VSUBS 0.007987f
C319 B.n279 VSUBS 0.007987f
C320 B.n280 VSUBS 0.007987f
C321 B.n281 VSUBS 0.007987f
C322 B.n282 VSUBS 0.007987f
C323 B.n283 VSUBS 0.007987f
C324 B.n284 VSUBS 0.007987f
C325 B.n285 VSUBS 0.007987f
C326 B.n286 VSUBS 0.007987f
C327 B.n287 VSUBS 0.007987f
C328 B.n288 VSUBS 0.007987f
C329 B.n289 VSUBS 0.007987f
C330 B.n290 VSUBS 0.007987f
C331 B.n291 VSUBS 0.007987f
C332 B.n292 VSUBS 0.007987f
C333 B.n293 VSUBS 0.007987f
C334 B.n294 VSUBS 0.007987f
C335 B.n295 VSUBS 0.007987f
C336 B.n296 VSUBS 0.007987f
C337 B.n297 VSUBS 0.007987f
C338 B.n298 VSUBS 0.007987f
C339 B.n299 VSUBS 0.007987f
C340 B.n300 VSUBS 0.007987f
C341 B.n301 VSUBS 0.007987f
C342 B.n302 VSUBS 0.007987f
C343 B.n303 VSUBS 0.007987f
C344 B.n304 VSUBS 0.007987f
C345 B.n305 VSUBS 0.007987f
C346 B.n306 VSUBS 0.007987f
C347 B.n307 VSUBS 0.007987f
C348 B.n308 VSUBS 0.007987f
C349 B.n309 VSUBS 0.007987f
C350 B.n310 VSUBS 0.007987f
C351 B.n311 VSUBS 0.007987f
C352 B.n312 VSUBS 0.007987f
C353 B.n313 VSUBS 0.007987f
C354 B.n314 VSUBS 0.007987f
C355 B.n315 VSUBS 0.007987f
C356 B.n316 VSUBS 0.007987f
C357 B.n317 VSUBS 0.007987f
C358 B.n318 VSUBS 0.007987f
C359 B.n319 VSUBS 0.007987f
C360 B.n320 VSUBS 0.007987f
C361 B.n321 VSUBS 0.007987f
C362 B.n322 VSUBS 0.007987f
C363 B.n323 VSUBS 0.007987f
C364 B.n324 VSUBS 0.007987f
C365 B.n325 VSUBS 0.007987f
C366 B.n326 VSUBS 0.007987f
C367 B.n327 VSUBS 0.007987f
C368 B.n328 VSUBS 0.007987f
C369 B.n329 VSUBS 0.007987f
C370 B.n330 VSUBS 0.007987f
C371 B.n331 VSUBS 0.007987f
C372 B.n332 VSUBS 0.007987f
C373 B.n333 VSUBS 0.007987f
C374 B.n334 VSUBS 0.007987f
C375 B.n335 VSUBS 0.007987f
C376 B.n336 VSUBS 0.007987f
C377 B.n337 VSUBS 0.007987f
C378 B.n338 VSUBS 0.007987f
C379 B.n339 VSUBS 0.007987f
C380 B.n340 VSUBS 0.007987f
C381 B.n341 VSUBS 0.007987f
C382 B.n342 VSUBS 0.007987f
C383 B.n343 VSUBS 0.007987f
C384 B.n344 VSUBS 0.007987f
C385 B.n345 VSUBS 0.007987f
C386 B.n346 VSUBS 0.007987f
C387 B.n347 VSUBS 0.007987f
C388 B.n348 VSUBS 0.007987f
C389 B.n349 VSUBS 0.007987f
C390 B.n350 VSUBS 0.007987f
C391 B.n351 VSUBS 0.007987f
C392 B.n352 VSUBS 0.007987f
C393 B.n353 VSUBS 0.007987f
C394 B.n354 VSUBS 0.01901f
C395 B.n355 VSUBS 0.018342f
C396 B.n356 VSUBS 0.019286f
C397 B.n357 VSUBS 0.007987f
C398 B.n358 VSUBS 0.007987f
C399 B.n359 VSUBS 0.007987f
C400 B.n360 VSUBS 0.007987f
C401 B.n361 VSUBS 0.007987f
C402 B.n362 VSUBS 0.007987f
C403 B.n363 VSUBS 0.007987f
C404 B.n364 VSUBS 0.007987f
C405 B.n365 VSUBS 0.007987f
C406 B.n366 VSUBS 0.007987f
C407 B.n367 VSUBS 0.007987f
C408 B.n368 VSUBS 0.007987f
C409 B.n369 VSUBS 0.007987f
C410 B.n370 VSUBS 0.007987f
C411 B.n371 VSUBS 0.007987f
C412 B.n372 VSUBS 0.007987f
C413 B.n373 VSUBS 0.007987f
C414 B.n374 VSUBS 0.007987f
C415 B.n375 VSUBS 0.007987f
C416 B.n376 VSUBS 0.007987f
C417 B.n377 VSUBS 0.007987f
C418 B.n378 VSUBS 0.007987f
C419 B.n379 VSUBS 0.007987f
C420 B.n380 VSUBS 0.007987f
C421 B.n381 VSUBS 0.007987f
C422 B.n382 VSUBS 0.007987f
C423 B.n383 VSUBS 0.007987f
C424 B.n384 VSUBS 0.007987f
C425 B.n385 VSUBS 0.007987f
C426 B.n386 VSUBS 0.007987f
C427 B.n387 VSUBS 0.007987f
C428 B.n388 VSUBS 0.007987f
C429 B.n389 VSUBS 0.007987f
C430 B.n390 VSUBS 0.007987f
C431 B.n391 VSUBS 0.00552f
C432 B.n392 VSUBS 0.007987f
C433 B.n393 VSUBS 0.007987f
C434 B.n394 VSUBS 0.00646f
C435 B.n395 VSUBS 0.007987f
C436 B.n396 VSUBS 0.007987f
C437 B.n397 VSUBS 0.007987f
C438 B.n398 VSUBS 0.007987f
C439 B.n399 VSUBS 0.007987f
C440 B.n400 VSUBS 0.007987f
C441 B.n401 VSUBS 0.007987f
C442 B.n402 VSUBS 0.007987f
C443 B.n403 VSUBS 0.007987f
C444 B.n404 VSUBS 0.007987f
C445 B.n405 VSUBS 0.007987f
C446 B.n406 VSUBS 0.00646f
C447 B.n407 VSUBS 0.018505f
C448 B.n408 VSUBS 0.00552f
C449 B.n409 VSUBS 0.007987f
C450 B.n410 VSUBS 0.007987f
C451 B.n411 VSUBS 0.007987f
C452 B.n412 VSUBS 0.007987f
C453 B.n413 VSUBS 0.007987f
C454 B.n414 VSUBS 0.007987f
C455 B.n415 VSUBS 0.007987f
C456 B.n416 VSUBS 0.007987f
C457 B.n417 VSUBS 0.007987f
C458 B.n418 VSUBS 0.007987f
C459 B.n419 VSUBS 0.007987f
C460 B.n420 VSUBS 0.007987f
C461 B.n421 VSUBS 0.007987f
C462 B.n422 VSUBS 0.007987f
C463 B.n423 VSUBS 0.007987f
C464 B.n424 VSUBS 0.007987f
C465 B.n425 VSUBS 0.007987f
C466 B.n426 VSUBS 0.007987f
C467 B.n427 VSUBS 0.007987f
C468 B.n428 VSUBS 0.007987f
C469 B.n429 VSUBS 0.007987f
C470 B.n430 VSUBS 0.007987f
C471 B.n431 VSUBS 0.007987f
C472 B.n432 VSUBS 0.007987f
C473 B.n433 VSUBS 0.007987f
C474 B.n434 VSUBS 0.007987f
C475 B.n435 VSUBS 0.007987f
C476 B.n436 VSUBS 0.007987f
C477 B.n437 VSUBS 0.007987f
C478 B.n438 VSUBS 0.007987f
C479 B.n439 VSUBS 0.007987f
C480 B.n440 VSUBS 0.007987f
C481 B.n441 VSUBS 0.007987f
C482 B.n442 VSUBS 0.007987f
C483 B.n443 VSUBS 0.007987f
C484 B.n444 VSUBS 0.019286f
C485 B.n445 VSUBS 0.018065f
C486 B.n446 VSUBS 0.018065f
C487 B.n447 VSUBS 0.007987f
C488 B.n448 VSUBS 0.007987f
C489 B.n449 VSUBS 0.007987f
C490 B.n450 VSUBS 0.007987f
C491 B.n451 VSUBS 0.007987f
C492 B.n452 VSUBS 0.007987f
C493 B.n453 VSUBS 0.007987f
C494 B.n454 VSUBS 0.007987f
C495 B.n455 VSUBS 0.007987f
C496 B.n456 VSUBS 0.007987f
C497 B.n457 VSUBS 0.007987f
C498 B.n458 VSUBS 0.007987f
C499 B.n459 VSUBS 0.007987f
C500 B.n460 VSUBS 0.007987f
C501 B.n461 VSUBS 0.007987f
C502 B.n462 VSUBS 0.007987f
C503 B.n463 VSUBS 0.007987f
C504 B.n464 VSUBS 0.007987f
C505 B.n465 VSUBS 0.007987f
C506 B.n466 VSUBS 0.007987f
C507 B.n467 VSUBS 0.007987f
C508 B.n468 VSUBS 0.007987f
C509 B.n469 VSUBS 0.007987f
C510 B.n470 VSUBS 0.007987f
C511 B.n471 VSUBS 0.007987f
C512 B.n472 VSUBS 0.007987f
C513 B.n473 VSUBS 0.007987f
C514 B.n474 VSUBS 0.007987f
C515 B.n475 VSUBS 0.007987f
C516 B.n476 VSUBS 0.007987f
C517 B.n477 VSUBS 0.007987f
C518 B.n478 VSUBS 0.007987f
C519 B.n479 VSUBS 0.007987f
C520 B.n480 VSUBS 0.007987f
C521 B.n481 VSUBS 0.007987f
C522 B.n482 VSUBS 0.007987f
C523 B.n483 VSUBS 0.007987f
C524 B.n484 VSUBS 0.007987f
C525 B.n485 VSUBS 0.007987f
C526 B.n486 VSUBS 0.007987f
C527 B.n487 VSUBS 0.007987f
C528 B.n488 VSUBS 0.007987f
C529 B.n489 VSUBS 0.007987f
C530 B.n490 VSUBS 0.007987f
C531 B.n491 VSUBS 0.018086f
C532 VDD2.t4 VSUBS 0.988899f
C533 VDD2.t5 VSUBS 0.107809f
C534 VDD2.t0 VSUBS 0.107809f
C535 VDD2.n0 VSUBS 0.739863f
C536 VDD2.n1 VSUBS 2.16153f
C537 VDD2.t2 VSUBS 0.983342f
C538 VDD2.n2 VSUBS 1.95243f
C539 VDD2.t1 VSUBS 0.107809f
C540 VDD2.t3 VSUBS 0.107809f
C541 VDD2.n3 VSUBS 0.73984f
C542 VN.n0 VSUBS 0.046643f
C543 VN.t5 VSUBS 1.18499f
C544 VN.n1 VSUBS 0.059415f
C545 VN.t1 VSUBS 1.34227f
C546 VN.n2 VSUBS 0.56441f
C547 VN.t0 VSUBS 1.18499f
C548 VN.n3 VSUBS 0.547877f
C549 VN.n4 VSUBS 0.065145f
C550 VN.n5 VSUBS 0.293432f
C551 VN.n6 VSUBS 0.046643f
C552 VN.n7 VSUBS 0.046643f
C553 VN.n8 VSUBS 0.076191f
C554 VN.n9 VSUBS 0.054043f
C555 VN.n10 VSUBS 0.549824f
C556 VN.n11 VSUBS 0.046547f
C557 VN.n12 VSUBS 0.046643f
C558 VN.t3 VSUBS 1.18499f
C559 VN.n13 VSUBS 0.059415f
C560 VN.t2 VSUBS 1.34227f
C561 VN.n14 VSUBS 0.56441f
C562 VN.t4 VSUBS 1.18499f
C563 VN.n15 VSUBS 0.547877f
C564 VN.n16 VSUBS 0.065145f
C565 VN.n17 VSUBS 0.293432f
C566 VN.n18 VSUBS 0.046643f
C567 VN.n19 VSUBS 0.046643f
C568 VN.n20 VSUBS 0.076191f
C569 VN.n21 VSUBS 0.054043f
C570 VN.n22 VSUBS 0.549824f
C571 VN.n23 VSUBS 1.8144f
C572 VDD1.t0 VSUBS 1.0031f
C573 VDD1.t3 VSUBS 1.00245f
C574 VDD1.t1 VSUBS 0.109287f
C575 VDD1.t2 VSUBS 0.109287f
C576 VDD1.n0 VSUBS 0.750004f
C577 VDD1.n1 VSUBS 2.27412f
C578 VDD1.t4 VSUBS 0.109287f
C579 VDD1.t5 VSUBS 0.109287f
C580 VDD1.n2 VSUBS 0.748161f
C581 VDD1.n3 VSUBS 1.97837f
C582 VTAIL.t5 VSUBS 0.155475f
C583 VTAIL.t3 VSUBS 0.155475f
C584 VTAIL.n0 VSUBS 0.958629f
C585 VTAIL.n1 VSUBS 0.73528f
C586 VTAIL.t7 VSUBS 1.30486f
C587 VTAIL.n2 VSUBS 0.930371f
C588 VTAIL.t6 VSUBS 0.155475f
C589 VTAIL.t8 VSUBS 0.155475f
C590 VTAIL.n3 VSUBS 0.958629f
C591 VTAIL.n4 VSUBS 2.02734f
C592 VTAIL.t0 VSUBS 0.155475f
C593 VTAIL.t1 VSUBS 0.155475f
C594 VTAIL.n5 VSUBS 0.958634f
C595 VTAIL.n6 VSUBS 2.02734f
C596 VTAIL.t4 VSUBS 1.30486f
C597 VTAIL.n7 VSUBS 0.930366f
C598 VTAIL.t10 VSUBS 0.155475f
C599 VTAIL.t9 VSUBS 0.155475f
C600 VTAIL.n8 VSUBS 0.958634f
C601 VTAIL.n9 VSUBS 0.852573f
C602 VTAIL.t11 VSUBS 1.30485f
C603 VTAIL.n10 VSUBS 1.94083f
C604 VTAIL.t2 VSUBS 1.30486f
C605 VTAIL.n11 VSUBS 1.89382f
C606 VP.n0 VSUBS 0.048616f
C607 VP.t3 VSUBS 1.23512f
C608 VP.n1 VSUBS 0.061928f
C609 VP.n2 VSUBS 0.048616f
C610 VP.t4 VSUBS 1.23512f
C611 VP.n3 VSUBS 0.079414f
C612 VP.n4 VSUBS 0.048616f
C613 VP.t0 VSUBS 1.23512f
C614 VP.n5 VSUBS 0.061928f
C615 VP.t5 VSUBS 1.39904f
C616 VP.n6 VSUBS 0.588284f
C617 VP.t1 VSUBS 1.23512f
C618 VP.n7 VSUBS 0.571053f
C619 VP.n8 VSUBS 0.0679f
C620 VP.n9 VSUBS 0.305844f
C621 VP.n10 VSUBS 0.048616f
C622 VP.n11 VSUBS 0.048616f
C623 VP.n12 VSUBS 0.079414f
C624 VP.n13 VSUBS 0.056329f
C625 VP.n14 VSUBS 0.573082f
C626 VP.n15 VSUBS 1.85913f
C627 VP.n16 VSUBS 1.90294f
C628 VP.t2 VSUBS 1.23512f
C629 VP.n17 VSUBS 0.573082f
C630 VP.n18 VSUBS 0.056329f
C631 VP.n19 VSUBS 0.048616f
C632 VP.n20 VSUBS 0.048616f
C633 VP.n21 VSUBS 0.048616f
C634 VP.n22 VSUBS 0.061928f
C635 VP.n23 VSUBS 0.0679f
C636 VP.n24 VSUBS 0.479526f
C637 VP.n25 VSUBS 0.0679f
C638 VP.n26 VSUBS 0.048616f
C639 VP.n27 VSUBS 0.048616f
C640 VP.n28 VSUBS 0.048616f
C641 VP.n29 VSUBS 0.079414f
C642 VP.n30 VSUBS 0.056329f
C643 VP.n31 VSUBS 0.573082f
C644 VP.n32 VSUBS 0.048516f
.ends

