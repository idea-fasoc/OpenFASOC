* NGSPICE file created from diff_pair_sample_1668.ext - technology: sky130A

.subckt diff_pair_sample_1668 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X1 B.t11 B.t9 B.t10 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.15
X2 VDD1.t6 VP.t1 VTAIL.t13 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X3 VDD2.t7 VN.t0 VTAIL.t7 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X4 VDD2.t6 VN.t1 VTAIL.t1 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.15
X5 VTAIL.t6 VN.t2 VDD2.t5 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X6 VTAIL.t14 VP.t2 VDD1.t5 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.15
X7 VTAIL.t5 VN.t3 VDD2.t4 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X8 VDD2.t3 VN.t4 VTAIL.t0 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.15
X9 VDD1.t4 VP.t3 VTAIL.t15 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.15
X10 VTAIL.t10 VP.t4 VDD1.t3 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X11 VDD1.t2 VP.t5 VTAIL.t11 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.15
X12 B.t8 B.t6 B.t7 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.15
X13 VDD2.t2 VN.t5 VTAIL.t4 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X14 VTAIL.t2 VN.t6 VDD2.t1 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.15
X15 VTAIL.t12 VP.t6 VDD1.t1 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.15
X16 B.t5 B.t3 B.t4 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.15
X17 VTAIL.t9 VP.t7 VDD1.t0 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=1.61535 pd=10.12 as=1.61535 ps=10.12 w=9.79 l=2.15
X18 VTAIL.t3 VN.t7 VDD2.t0 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.15
X19 B.t2 B.t0 B.t1 w_n3450_n2926# sky130_fd_pr__pfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.15
R0 VP.n15 VP.n12 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n18 VP.n11 161.3
R3 VP.n20 VP.n19 161.3
R4 VP.n22 VP.n10 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n9 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n28 VP.n8 161.3
R9 VP.n54 VP.n0 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n1 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n2 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n3 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n41 VP.n4 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n5 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n6 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n13 VP.t2 144.333
R24 VP.n7 VP.t6 109.74
R25 VP.n40 VP.t0 109.74
R26 VP.n47 VP.t4 109.74
R27 VP.n55 VP.t3 109.74
R28 VP.n29 VP.t5 109.74
R29 VP.n21 VP.t7 109.74
R30 VP.n14 VP.t1 109.74
R31 VP.n31 VP.n7 87.7575
R32 VP.n56 VP.n55 87.7575
R33 VP.n30 VP.n29 87.7575
R34 VP.n35 VP.n34 56.5193
R35 VP.n42 VP.n3 56.5193
R36 VP.n53 VP.n1 56.5193
R37 VP.n27 VP.n9 56.5193
R38 VP.n16 VP.n11 56.5193
R39 VP.n31 VP.n30 47.2269
R40 VP.n14 VP.n13 46.8391
R41 VP.n34 VP.n33 24.4675
R42 VP.n35 VP.n5 24.4675
R43 VP.n39 VP.n5 24.4675
R44 VP.n42 VP.n41 24.4675
R45 VP.n46 VP.n3 24.4675
R46 VP.n49 VP.n48 24.4675
R47 VP.n49 VP.n1 24.4675
R48 VP.n54 VP.n53 24.4675
R49 VP.n28 VP.n27 24.4675
R50 VP.n20 VP.n11 24.4675
R51 VP.n23 VP.n22 24.4675
R52 VP.n23 VP.n9 24.4675
R53 VP.n16 VP.n15 24.4675
R54 VP.n41 VP.n40 23.9782
R55 VP.n47 VP.n46 23.9782
R56 VP.n21 VP.n20 23.9782
R57 VP.n15 VP.n14 23.9782
R58 VP.n33 VP.n7 22.9995
R59 VP.n55 VP.n54 22.9995
R60 VP.n29 VP.n28 22.9995
R61 VP.n13 VP.n12 8.69054
R62 VP.n40 VP.n39 0.48984
R63 VP.n48 VP.n47 0.48984
R64 VP.n22 VP.n21 0.48984
R65 VP.n30 VP.n8 0.278367
R66 VP.n32 VP.n31 0.278367
R67 VP.n56 VP.n0 0.278367
R68 VP.n17 VP.n12 0.189894
R69 VP.n18 VP.n17 0.189894
R70 VP.n19 VP.n18 0.189894
R71 VP.n19 VP.n10 0.189894
R72 VP.n24 VP.n10 0.189894
R73 VP.n25 VP.n24 0.189894
R74 VP.n26 VP.n25 0.189894
R75 VP.n26 VP.n8 0.189894
R76 VP.n32 VP.n6 0.189894
R77 VP.n36 VP.n6 0.189894
R78 VP.n37 VP.n36 0.189894
R79 VP.n38 VP.n37 0.189894
R80 VP.n38 VP.n4 0.189894
R81 VP.n43 VP.n4 0.189894
R82 VP.n44 VP.n43 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n45 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VP VP.n56 0.153454
R90 VTAIL.n11 VTAIL.t14 68.1466
R91 VTAIL.n10 VTAIL.t0 68.1466
R92 VTAIL.n7 VTAIL.t3 68.1466
R93 VTAIL.n15 VTAIL.t1 68.1465
R94 VTAIL.n2 VTAIL.t2 68.1465
R95 VTAIL.n3 VTAIL.t15 68.1465
R96 VTAIL.n6 VTAIL.t12 68.1465
R97 VTAIL.n14 VTAIL.t11 68.1465
R98 VTAIL.n13 VTAIL.n12 64.8265
R99 VTAIL.n9 VTAIL.n8 64.8265
R100 VTAIL.n1 VTAIL.n0 64.8262
R101 VTAIL.n5 VTAIL.n4 64.8262
R102 VTAIL.n15 VTAIL.n14 22.9445
R103 VTAIL.n7 VTAIL.n6 22.9445
R104 VTAIL.n0 VTAIL.t4 3.32072
R105 VTAIL.n0 VTAIL.t5 3.32072
R106 VTAIL.n4 VTAIL.t8 3.32072
R107 VTAIL.n4 VTAIL.t10 3.32072
R108 VTAIL.n12 VTAIL.t13 3.32072
R109 VTAIL.n12 VTAIL.t9 3.32072
R110 VTAIL.n8 VTAIL.t7 3.32072
R111 VTAIL.n8 VTAIL.t6 3.32072
R112 VTAIL.n9 VTAIL.n7 2.13843
R113 VTAIL.n10 VTAIL.n9 2.13843
R114 VTAIL.n13 VTAIL.n11 2.13843
R115 VTAIL.n14 VTAIL.n13 2.13843
R116 VTAIL.n6 VTAIL.n5 2.13843
R117 VTAIL.n5 VTAIL.n3 2.13843
R118 VTAIL.n2 VTAIL.n1 2.13843
R119 VTAIL VTAIL.n15 2.08024
R120 VTAIL.n11 VTAIL.n10 0.470328
R121 VTAIL.n3 VTAIL.n2 0.470328
R122 VTAIL VTAIL.n1 0.0586897
R123 VDD1 VDD1.n0 82.6324
R124 VDD1.n3 VDD1.n2 82.5186
R125 VDD1.n3 VDD1.n1 82.5186
R126 VDD1.n5 VDD1.n4 81.505
R127 VDD1.n5 VDD1.n3 42.3586
R128 VDD1.n4 VDD1.t0 3.32072
R129 VDD1.n4 VDD1.t2 3.32072
R130 VDD1.n0 VDD1.t5 3.32072
R131 VDD1.n0 VDD1.t6 3.32072
R132 VDD1.n2 VDD1.t3 3.32072
R133 VDD1.n2 VDD1.t4 3.32072
R134 VDD1.n1 VDD1.t1 3.32072
R135 VDD1.n1 VDD1.t7 3.32072
R136 VDD1 VDD1.n5 1.01128
R137 B.n365 B.n114 585
R138 B.n364 B.n363 585
R139 B.n362 B.n115 585
R140 B.n361 B.n360 585
R141 B.n359 B.n116 585
R142 B.n358 B.n357 585
R143 B.n356 B.n117 585
R144 B.n355 B.n354 585
R145 B.n353 B.n118 585
R146 B.n352 B.n351 585
R147 B.n350 B.n119 585
R148 B.n349 B.n348 585
R149 B.n347 B.n120 585
R150 B.n346 B.n345 585
R151 B.n344 B.n121 585
R152 B.n343 B.n342 585
R153 B.n341 B.n122 585
R154 B.n340 B.n339 585
R155 B.n338 B.n123 585
R156 B.n337 B.n336 585
R157 B.n335 B.n124 585
R158 B.n334 B.n333 585
R159 B.n332 B.n125 585
R160 B.n331 B.n330 585
R161 B.n329 B.n126 585
R162 B.n328 B.n327 585
R163 B.n326 B.n127 585
R164 B.n325 B.n324 585
R165 B.n323 B.n128 585
R166 B.n322 B.n321 585
R167 B.n320 B.n129 585
R168 B.n319 B.n318 585
R169 B.n317 B.n130 585
R170 B.n316 B.n315 585
R171 B.n314 B.n131 585
R172 B.n313 B.n312 585
R173 B.n308 B.n132 585
R174 B.n307 B.n306 585
R175 B.n305 B.n133 585
R176 B.n304 B.n303 585
R177 B.n302 B.n134 585
R178 B.n301 B.n300 585
R179 B.n299 B.n135 585
R180 B.n298 B.n297 585
R181 B.n296 B.n136 585
R182 B.n294 B.n293 585
R183 B.n292 B.n139 585
R184 B.n291 B.n290 585
R185 B.n289 B.n140 585
R186 B.n288 B.n287 585
R187 B.n286 B.n141 585
R188 B.n285 B.n284 585
R189 B.n283 B.n142 585
R190 B.n282 B.n281 585
R191 B.n280 B.n143 585
R192 B.n279 B.n278 585
R193 B.n277 B.n144 585
R194 B.n276 B.n275 585
R195 B.n274 B.n145 585
R196 B.n273 B.n272 585
R197 B.n271 B.n146 585
R198 B.n270 B.n269 585
R199 B.n268 B.n147 585
R200 B.n267 B.n266 585
R201 B.n265 B.n148 585
R202 B.n264 B.n263 585
R203 B.n262 B.n149 585
R204 B.n261 B.n260 585
R205 B.n259 B.n150 585
R206 B.n258 B.n257 585
R207 B.n256 B.n151 585
R208 B.n255 B.n254 585
R209 B.n253 B.n152 585
R210 B.n252 B.n251 585
R211 B.n250 B.n153 585
R212 B.n249 B.n248 585
R213 B.n247 B.n154 585
R214 B.n246 B.n245 585
R215 B.n244 B.n155 585
R216 B.n243 B.n242 585
R217 B.n367 B.n366 585
R218 B.n368 B.n113 585
R219 B.n370 B.n369 585
R220 B.n371 B.n112 585
R221 B.n373 B.n372 585
R222 B.n374 B.n111 585
R223 B.n376 B.n375 585
R224 B.n377 B.n110 585
R225 B.n379 B.n378 585
R226 B.n380 B.n109 585
R227 B.n382 B.n381 585
R228 B.n383 B.n108 585
R229 B.n385 B.n384 585
R230 B.n386 B.n107 585
R231 B.n388 B.n387 585
R232 B.n389 B.n106 585
R233 B.n391 B.n390 585
R234 B.n392 B.n105 585
R235 B.n394 B.n393 585
R236 B.n395 B.n104 585
R237 B.n397 B.n396 585
R238 B.n398 B.n103 585
R239 B.n400 B.n399 585
R240 B.n401 B.n102 585
R241 B.n403 B.n402 585
R242 B.n404 B.n101 585
R243 B.n406 B.n405 585
R244 B.n407 B.n100 585
R245 B.n409 B.n408 585
R246 B.n410 B.n99 585
R247 B.n412 B.n411 585
R248 B.n413 B.n98 585
R249 B.n415 B.n414 585
R250 B.n416 B.n97 585
R251 B.n418 B.n417 585
R252 B.n419 B.n96 585
R253 B.n421 B.n420 585
R254 B.n422 B.n95 585
R255 B.n424 B.n423 585
R256 B.n425 B.n94 585
R257 B.n427 B.n426 585
R258 B.n428 B.n93 585
R259 B.n430 B.n429 585
R260 B.n431 B.n92 585
R261 B.n433 B.n432 585
R262 B.n434 B.n91 585
R263 B.n436 B.n435 585
R264 B.n437 B.n90 585
R265 B.n439 B.n438 585
R266 B.n440 B.n89 585
R267 B.n442 B.n441 585
R268 B.n443 B.n88 585
R269 B.n445 B.n444 585
R270 B.n446 B.n87 585
R271 B.n448 B.n447 585
R272 B.n449 B.n86 585
R273 B.n451 B.n450 585
R274 B.n452 B.n85 585
R275 B.n454 B.n453 585
R276 B.n455 B.n84 585
R277 B.n457 B.n456 585
R278 B.n458 B.n83 585
R279 B.n460 B.n459 585
R280 B.n461 B.n82 585
R281 B.n463 B.n462 585
R282 B.n464 B.n81 585
R283 B.n466 B.n465 585
R284 B.n467 B.n80 585
R285 B.n469 B.n468 585
R286 B.n470 B.n79 585
R287 B.n472 B.n471 585
R288 B.n473 B.n78 585
R289 B.n475 B.n474 585
R290 B.n476 B.n77 585
R291 B.n478 B.n477 585
R292 B.n479 B.n76 585
R293 B.n481 B.n480 585
R294 B.n482 B.n75 585
R295 B.n484 B.n483 585
R296 B.n485 B.n74 585
R297 B.n487 B.n486 585
R298 B.n488 B.n73 585
R299 B.n490 B.n489 585
R300 B.n491 B.n72 585
R301 B.n493 B.n492 585
R302 B.n494 B.n71 585
R303 B.n496 B.n495 585
R304 B.n497 B.n70 585
R305 B.n499 B.n498 585
R306 B.n500 B.n69 585
R307 B.n621 B.n24 585
R308 B.n620 B.n619 585
R309 B.n618 B.n25 585
R310 B.n617 B.n616 585
R311 B.n615 B.n26 585
R312 B.n614 B.n613 585
R313 B.n612 B.n27 585
R314 B.n611 B.n610 585
R315 B.n609 B.n28 585
R316 B.n608 B.n607 585
R317 B.n606 B.n29 585
R318 B.n605 B.n604 585
R319 B.n603 B.n30 585
R320 B.n602 B.n601 585
R321 B.n600 B.n31 585
R322 B.n599 B.n598 585
R323 B.n597 B.n32 585
R324 B.n596 B.n595 585
R325 B.n594 B.n33 585
R326 B.n593 B.n592 585
R327 B.n591 B.n34 585
R328 B.n590 B.n589 585
R329 B.n588 B.n35 585
R330 B.n587 B.n586 585
R331 B.n585 B.n36 585
R332 B.n584 B.n583 585
R333 B.n582 B.n37 585
R334 B.n581 B.n580 585
R335 B.n579 B.n38 585
R336 B.n578 B.n577 585
R337 B.n576 B.n39 585
R338 B.n575 B.n574 585
R339 B.n573 B.n40 585
R340 B.n572 B.n571 585
R341 B.n570 B.n41 585
R342 B.n568 B.n567 585
R343 B.n566 B.n44 585
R344 B.n565 B.n564 585
R345 B.n563 B.n45 585
R346 B.n562 B.n561 585
R347 B.n560 B.n46 585
R348 B.n559 B.n558 585
R349 B.n557 B.n47 585
R350 B.n556 B.n555 585
R351 B.n554 B.n48 585
R352 B.n553 B.n552 585
R353 B.n551 B.n49 585
R354 B.n550 B.n549 585
R355 B.n548 B.n53 585
R356 B.n547 B.n546 585
R357 B.n545 B.n54 585
R358 B.n544 B.n543 585
R359 B.n542 B.n55 585
R360 B.n541 B.n540 585
R361 B.n539 B.n56 585
R362 B.n538 B.n537 585
R363 B.n536 B.n57 585
R364 B.n535 B.n534 585
R365 B.n533 B.n58 585
R366 B.n532 B.n531 585
R367 B.n530 B.n59 585
R368 B.n529 B.n528 585
R369 B.n527 B.n60 585
R370 B.n526 B.n525 585
R371 B.n524 B.n61 585
R372 B.n523 B.n522 585
R373 B.n521 B.n62 585
R374 B.n520 B.n519 585
R375 B.n518 B.n63 585
R376 B.n517 B.n516 585
R377 B.n515 B.n64 585
R378 B.n514 B.n513 585
R379 B.n512 B.n65 585
R380 B.n511 B.n510 585
R381 B.n509 B.n66 585
R382 B.n508 B.n507 585
R383 B.n506 B.n67 585
R384 B.n505 B.n504 585
R385 B.n503 B.n68 585
R386 B.n502 B.n501 585
R387 B.n623 B.n622 585
R388 B.n624 B.n23 585
R389 B.n626 B.n625 585
R390 B.n627 B.n22 585
R391 B.n629 B.n628 585
R392 B.n630 B.n21 585
R393 B.n632 B.n631 585
R394 B.n633 B.n20 585
R395 B.n635 B.n634 585
R396 B.n636 B.n19 585
R397 B.n638 B.n637 585
R398 B.n639 B.n18 585
R399 B.n641 B.n640 585
R400 B.n642 B.n17 585
R401 B.n644 B.n643 585
R402 B.n645 B.n16 585
R403 B.n647 B.n646 585
R404 B.n648 B.n15 585
R405 B.n650 B.n649 585
R406 B.n651 B.n14 585
R407 B.n653 B.n652 585
R408 B.n654 B.n13 585
R409 B.n656 B.n655 585
R410 B.n657 B.n12 585
R411 B.n659 B.n658 585
R412 B.n660 B.n11 585
R413 B.n662 B.n661 585
R414 B.n663 B.n10 585
R415 B.n665 B.n664 585
R416 B.n666 B.n9 585
R417 B.n668 B.n667 585
R418 B.n669 B.n8 585
R419 B.n671 B.n670 585
R420 B.n672 B.n7 585
R421 B.n674 B.n673 585
R422 B.n675 B.n6 585
R423 B.n677 B.n676 585
R424 B.n678 B.n5 585
R425 B.n680 B.n679 585
R426 B.n681 B.n4 585
R427 B.n683 B.n682 585
R428 B.n684 B.n3 585
R429 B.n686 B.n685 585
R430 B.n687 B.n0 585
R431 B.n2 B.n1 585
R432 B.n178 B.n177 585
R433 B.n180 B.n179 585
R434 B.n181 B.n176 585
R435 B.n183 B.n182 585
R436 B.n184 B.n175 585
R437 B.n186 B.n185 585
R438 B.n187 B.n174 585
R439 B.n189 B.n188 585
R440 B.n190 B.n173 585
R441 B.n192 B.n191 585
R442 B.n193 B.n172 585
R443 B.n195 B.n194 585
R444 B.n196 B.n171 585
R445 B.n198 B.n197 585
R446 B.n199 B.n170 585
R447 B.n201 B.n200 585
R448 B.n202 B.n169 585
R449 B.n204 B.n203 585
R450 B.n205 B.n168 585
R451 B.n207 B.n206 585
R452 B.n208 B.n167 585
R453 B.n210 B.n209 585
R454 B.n211 B.n166 585
R455 B.n213 B.n212 585
R456 B.n214 B.n165 585
R457 B.n216 B.n215 585
R458 B.n217 B.n164 585
R459 B.n219 B.n218 585
R460 B.n220 B.n163 585
R461 B.n222 B.n221 585
R462 B.n223 B.n162 585
R463 B.n225 B.n224 585
R464 B.n226 B.n161 585
R465 B.n228 B.n227 585
R466 B.n229 B.n160 585
R467 B.n231 B.n230 585
R468 B.n232 B.n159 585
R469 B.n234 B.n233 585
R470 B.n235 B.n158 585
R471 B.n237 B.n236 585
R472 B.n238 B.n157 585
R473 B.n240 B.n239 585
R474 B.n241 B.n156 585
R475 B.n243 B.n156 497.305
R476 B.n367 B.n114 497.305
R477 B.n501 B.n500 497.305
R478 B.n622 B.n621 497.305
R479 B.n137 B.t3 316.988
R480 B.n309 B.t0 316.988
R481 B.n50 B.t6 316.988
R482 B.n42 B.t9 316.988
R483 B.n689 B.n688 256.663
R484 B.n688 B.n687 235.042
R485 B.n688 B.n2 235.042
R486 B.n244 B.n243 163.367
R487 B.n245 B.n244 163.367
R488 B.n245 B.n154 163.367
R489 B.n249 B.n154 163.367
R490 B.n250 B.n249 163.367
R491 B.n251 B.n250 163.367
R492 B.n251 B.n152 163.367
R493 B.n255 B.n152 163.367
R494 B.n256 B.n255 163.367
R495 B.n257 B.n256 163.367
R496 B.n257 B.n150 163.367
R497 B.n261 B.n150 163.367
R498 B.n262 B.n261 163.367
R499 B.n263 B.n262 163.367
R500 B.n263 B.n148 163.367
R501 B.n267 B.n148 163.367
R502 B.n268 B.n267 163.367
R503 B.n269 B.n268 163.367
R504 B.n269 B.n146 163.367
R505 B.n273 B.n146 163.367
R506 B.n274 B.n273 163.367
R507 B.n275 B.n274 163.367
R508 B.n275 B.n144 163.367
R509 B.n279 B.n144 163.367
R510 B.n280 B.n279 163.367
R511 B.n281 B.n280 163.367
R512 B.n281 B.n142 163.367
R513 B.n285 B.n142 163.367
R514 B.n286 B.n285 163.367
R515 B.n287 B.n286 163.367
R516 B.n287 B.n140 163.367
R517 B.n291 B.n140 163.367
R518 B.n292 B.n291 163.367
R519 B.n293 B.n292 163.367
R520 B.n293 B.n136 163.367
R521 B.n298 B.n136 163.367
R522 B.n299 B.n298 163.367
R523 B.n300 B.n299 163.367
R524 B.n300 B.n134 163.367
R525 B.n304 B.n134 163.367
R526 B.n305 B.n304 163.367
R527 B.n306 B.n305 163.367
R528 B.n306 B.n132 163.367
R529 B.n313 B.n132 163.367
R530 B.n314 B.n313 163.367
R531 B.n315 B.n314 163.367
R532 B.n315 B.n130 163.367
R533 B.n319 B.n130 163.367
R534 B.n320 B.n319 163.367
R535 B.n321 B.n320 163.367
R536 B.n321 B.n128 163.367
R537 B.n325 B.n128 163.367
R538 B.n326 B.n325 163.367
R539 B.n327 B.n326 163.367
R540 B.n327 B.n126 163.367
R541 B.n331 B.n126 163.367
R542 B.n332 B.n331 163.367
R543 B.n333 B.n332 163.367
R544 B.n333 B.n124 163.367
R545 B.n337 B.n124 163.367
R546 B.n338 B.n337 163.367
R547 B.n339 B.n338 163.367
R548 B.n339 B.n122 163.367
R549 B.n343 B.n122 163.367
R550 B.n344 B.n343 163.367
R551 B.n345 B.n344 163.367
R552 B.n345 B.n120 163.367
R553 B.n349 B.n120 163.367
R554 B.n350 B.n349 163.367
R555 B.n351 B.n350 163.367
R556 B.n351 B.n118 163.367
R557 B.n355 B.n118 163.367
R558 B.n356 B.n355 163.367
R559 B.n357 B.n356 163.367
R560 B.n357 B.n116 163.367
R561 B.n361 B.n116 163.367
R562 B.n362 B.n361 163.367
R563 B.n363 B.n362 163.367
R564 B.n363 B.n114 163.367
R565 B.n500 B.n499 163.367
R566 B.n499 B.n70 163.367
R567 B.n495 B.n70 163.367
R568 B.n495 B.n494 163.367
R569 B.n494 B.n493 163.367
R570 B.n493 B.n72 163.367
R571 B.n489 B.n72 163.367
R572 B.n489 B.n488 163.367
R573 B.n488 B.n487 163.367
R574 B.n487 B.n74 163.367
R575 B.n483 B.n74 163.367
R576 B.n483 B.n482 163.367
R577 B.n482 B.n481 163.367
R578 B.n481 B.n76 163.367
R579 B.n477 B.n76 163.367
R580 B.n477 B.n476 163.367
R581 B.n476 B.n475 163.367
R582 B.n475 B.n78 163.367
R583 B.n471 B.n78 163.367
R584 B.n471 B.n470 163.367
R585 B.n470 B.n469 163.367
R586 B.n469 B.n80 163.367
R587 B.n465 B.n80 163.367
R588 B.n465 B.n464 163.367
R589 B.n464 B.n463 163.367
R590 B.n463 B.n82 163.367
R591 B.n459 B.n82 163.367
R592 B.n459 B.n458 163.367
R593 B.n458 B.n457 163.367
R594 B.n457 B.n84 163.367
R595 B.n453 B.n84 163.367
R596 B.n453 B.n452 163.367
R597 B.n452 B.n451 163.367
R598 B.n451 B.n86 163.367
R599 B.n447 B.n86 163.367
R600 B.n447 B.n446 163.367
R601 B.n446 B.n445 163.367
R602 B.n445 B.n88 163.367
R603 B.n441 B.n88 163.367
R604 B.n441 B.n440 163.367
R605 B.n440 B.n439 163.367
R606 B.n439 B.n90 163.367
R607 B.n435 B.n90 163.367
R608 B.n435 B.n434 163.367
R609 B.n434 B.n433 163.367
R610 B.n433 B.n92 163.367
R611 B.n429 B.n92 163.367
R612 B.n429 B.n428 163.367
R613 B.n428 B.n427 163.367
R614 B.n427 B.n94 163.367
R615 B.n423 B.n94 163.367
R616 B.n423 B.n422 163.367
R617 B.n422 B.n421 163.367
R618 B.n421 B.n96 163.367
R619 B.n417 B.n96 163.367
R620 B.n417 B.n416 163.367
R621 B.n416 B.n415 163.367
R622 B.n415 B.n98 163.367
R623 B.n411 B.n98 163.367
R624 B.n411 B.n410 163.367
R625 B.n410 B.n409 163.367
R626 B.n409 B.n100 163.367
R627 B.n405 B.n100 163.367
R628 B.n405 B.n404 163.367
R629 B.n404 B.n403 163.367
R630 B.n403 B.n102 163.367
R631 B.n399 B.n102 163.367
R632 B.n399 B.n398 163.367
R633 B.n398 B.n397 163.367
R634 B.n397 B.n104 163.367
R635 B.n393 B.n104 163.367
R636 B.n393 B.n392 163.367
R637 B.n392 B.n391 163.367
R638 B.n391 B.n106 163.367
R639 B.n387 B.n106 163.367
R640 B.n387 B.n386 163.367
R641 B.n386 B.n385 163.367
R642 B.n385 B.n108 163.367
R643 B.n381 B.n108 163.367
R644 B.n381 B.n380 163.367
R645 B.n380 B.n379 163.367
R646 B.n379 B.n110 163.367
R647 B.n375 B.n110 163.367
R648 B.n375 B.n374 163.367
R649 B.n374 B.n373 163.367
R650 B.n373 B.n112 163.367
R651 B.n369 B.n112 163.367
R652 B.n369 B.n368 163.367
R653 B.n368 B.n367 163.367
R654 B.n621 B.n620 163.367
R655 B.n620 B.n25 163.367
R656 B.n616 B.n25 163.367
R657 B.n616 B.n615 163.367
R658 B.n615 B.n614 163.367
R659 B.n614 B.n27 163.367
R660 B.n610 B.n27 163.367
R661 B.n610 B.n609 163.367
R662 B.n609 B.n608 163.367
R663 B.n608 B.n29 163.367
R664 B.n604 B.n29 163.367
R665 B.n604 B.n603 163.367
R666 B.n603 B.n602 163.367
R667 B.n602 B.n31 163.367
R668 B.n598 B.n31 163.367
R669 B.n598 B.n597 163.367
R670 B.n597 B.n596 163.367
R671 B.n596 B.n33 163.367
R672 B.n592 B.n33 163.367
R673 B.n592 B.n591 163.367
R674 B.n591 B.n590 163.367
R675 B.n590 B.n35 163.367
R676 B.n586 B.n35 163.367
R677 B.n586 B.n585 163.367
R678 B.n585 B.n584 163.367
R679 B.n584 B.n37 163.367
R680 B.n580 B.n37 163.367
R681 B.n580 B.n579 163.367
R682 B.n579 B.n578 163.367
R683 B.n578 B.n39 163.367
R684 B.n574 B.n39 163.367
R685 B.n574 B.n573 163.367
R686 B.n573 B.n572 163.367
R687 B.n572 B.n41 163.367
R688 B.n567 B.n41 163.367
R689 B.n567 B.n566 163.367
R690 B.n566 B.n565 163.367
R691 B.n565 B.n45 163.367
R692 B.n561 B.n45 163.367
R693 B.n561 B.n560 163.367
R694 B.n560 B.n559 163.367
R695 B.n559 B.n47 163.367
R696 B.n555 B.n47 163.367
R697 B.n555 B.n554 163.367
R698 B.n554 B.n553 163.367
R699 B.n553 B.n49 163.367
R700 B.n549 B.n49 163.367
R701 B.n549 B.n548 163.367
R702 B.n548 B.n547 163.367
R703 B.n547 B.n54 163.367
R704 B.n543 B.n54 163.367
R705 B.n543 B.n542 163.367
R706 B.n542 B.n541 163.367
R707 B.n541 B.n56 163.367
R708 B.n537 B.n56 163.367
R709 B.n537 B.n536 163.367
R710 B.n536 B.n535 163.367
R711 B.n535 B.n58 163.367
R712 B.n531 B.n58 163.367
R713 B.n531 B.n530 163.367
R714 B.n530 B.n529 163.367
R715 B.n529 B.n60 163.367
R716 B.n525 B.n60 163.367
R717 B.n525 B.n524 163.367
R718 B.n524 B.n523 163.367
R719 B.n523 B.n62 163.367
R720 B.n519 B.n62 163.367
R721 B.n519 B.n518 163.367
R722 B.n518 B.n517 163.367
R723 B.n517 B.n64 163.367
R724 B.n513 B.n64 163.367
R725 B.n513 B.n512 163.367
R726 B.n512 B.n511 163.367
R727 B.n511 B.n66 163.367
R728 B.n507 B.n66 163.367
R729 B.n507 B.n506 163.367
R730 B.n506 B.n505 163.367
R731 B.n505 B.n68 163.367
R732 B.n501 B.n68 163.367
R733 B.n622 B.n23 163.367
R734 B.n626 B.n23 163.367
R735 B.n627 B.n626 163.367
R736 B.n628 B.n627 163.367
R737 B.n628 B.n21 163.367
R738 B.n632 B.n21 163.367
R739 B.n633 B.n632 163.367
R740 B.n634 B.n633 163.367
R741 B.n634 B.n19 163.367
R742 B.n638 B.n19 163.367
R743 B.n639 B.n638 163.367
R744 B.n640 B.n639 163.367
R745 B.n640 B.n17 163.367
R746 B.n644 B.n17 163.367
R747 B.n645 B.n644 163.367
R748 B.n646 B.n645 163.367
R749 B.n646 B.n15 163.367
R750 B.n650 B.n15 163.367
R751 B.n651 B.n650 163.367
R752 B.n652 B.n651 163.367
R753 B.n652 B.n13 163.367
R754 B.n656 B.n13 163.367
R755 B.n657 B.n656 163.367
R756 B.n658 B.n657 163.367
R757 B.n658 B.n11 163.367
R758 B.n662 B.n11 163.367
R759 B.n663 B.n662 163.367
R760 B.n664 B.n663 163.367
R761 B.n664 B.n9 163.367
R762 B.n668 B.n9 163.367
R763 B.n669 B.n668 163.367
R764 B.n670 B.n669 163.367
R765 B.n670 B.n7 163.367
R766 B.n674 B.n7 163.367
R767 B.n675 B.n674 163.367
R768 B.n676 B.n675 163.367
R769 B.n676 B.n5 163.367
R770 B.n680 B.n5 163.367
R771 B.n681 B.n680 163.367
R772 B.n682 B.n681 163.367
R773 B.n682 B.n3 163.367
R774 B.n686 B.n3 163.367
R775 B.n687 B.n686 163.367
R776 B.n178 B.n2 163.367
R777 B.n179 B.n178 163.367
R778 B.n179 B.n176 163.367
R779 B.n183 B.n176 163.367
R780 B.n184 B.n183 163.367
R781 B.n185 B.n184 163.367
R782 B.n185 B.n174 163.367
R783 B.n189 B.n174 163.367
R784 B.n190 B.n189 163.367
R785 B.n191 B.n190 163.367
R786 B.n191 B.n172 163.367
R787 B.n195 B.n172 163.367
R788 B.n196 B.n195 163.367
R789 B.n197 B.n196 163.367
R790 B.n197 B.n170 163.367
R791 B.n201 B.n170 163.367
R792 B.n202 B.n201 163.367
R793 B.n203 B.n202 163.367
R794 B.n203 B.n168 163.367
R795 B.n207 B.n168 163.367
R796 B.n208 B.n207 163.367
R797 B.n209 B.n208 163.367
R798 B.n209 B.n166 163.367
R799 B.n213 B.n166 163.367
R800 B.n214 B.n213 163.367
R801 B.n215 B.n214 163.367
R802 B.n215 B.n164 163.367
R803 B.n219 B.n164 163.367
R804 B.n220 B.n219 163.367
R805 B.n221 B.n220 163.367
R806 B.n221 B.n162 163.367
R807 B.n225 B.n162 163.367
R808 B.n226 B.n225 163.367
R809 B.n227 B.n226 163.367
R810 B.n227 B.n160 163.367
R811 B.n231 B.n160 163.367
R812 B.n232 B.n231 163.367
R813 B.n233 B.n232 163.367
R814 B.n233 B.n158 163.367
R815 B.n237 B.n158 163.367
R816 B.n238 B.n237 163.367
R817 B.n239 B.n238 163.367
R818 B.n239 B.n156 163.367
R819 B.n309 B.t1 161.094
R820 B.n50 B.t8 161.094
R821 B.n137 B.t4 161.082
R822 B.n42 B.t11 161.082
R823 B.n310 B.t2 112.996
R824 B.n51 B.t7 112.996
R825 B.n138 B.t5 112.984
R826 B.n43 B.t10 112.984
R827 B.n295 B.n138 59.5399
R828 B.n311 B.n310 59.5399
R829 B.n52 B.n51 59.5399
R830 B.n569 B.n43 59.5399
R831 B.n138 B.n137 48.0975
R832 B.n310 B.n309 48.0975
R833 B.n51 B.n50 48.0975
R834 B.n43 B.n42 48.0975
R835 B.n623 B.n24 32.3127
R836 B.n502 B.n69 32.3127
R837 B.n366 B.n365 32.3127
R838 B.n242 B.n241 32.3127
R839 B B.n689 18.0485
R840 B.n624 B.n623 10.6151
R841 B.n625 B.n624 10.6151
R842 B.n625 B.n22 10.6151
R843 B.n629 B.n22 10.6151
R844 B.n630 B.n629 10.6151
R845 B.n631 B.n630 10.6151
R846 B.n631 B.n20 10.6151
R847 B.n635 B.n20 10.6151
R848 B.n636 B.n635 10.6151
R849 B.n637 B.n636 10.6151
R850 B.n637 B.n18 10.6151
R851 B.n641 B.n18 10.6151
R852 B.n642 B.n641 10.6151
R853 B.n643 B.n642 10.6151
R854 B.n643 B.n16 10.6151
R855 B.n647 B.n16 10.6151
R856 B.n648 B.n647 10.6151
R857 B.n649 B.n648 10.6151
R858 B.n649 B.n14 10.6151
R859 B.n653 B.n14 10.6151
R860 B.n654 B.n653 10.6151
R861 B.n655 B.n654 10.6151
R862 B.n655 B.n12 10.6151
R863 B.n659 B.n12 10.6151
R864 B.n660 B.n659 10.6151
R865 B.n661 B.n660 10.6151
R866 B.n661 B.n10 10.6151
R867 B.n665 B.n10 10.6151
R868 B.n666 B.n665 10.6151
R869 B.n667 B.n666 10.6151
R870 B.n667 B.n8 10.6151
R871 B.n671 B.n8 10.6151
R872 B.n672 B.n671 10.6151
R873 B.n673 B.n672 10.6151
R874 B.n673 B.n6 10.6151
R875 B.n677 B.n6 10.6151
R876 B.n678 B.n677 10.6151
R877 B.n679 B.n678 10.6151
R878 B.n679 B.n4 10.6151
R879 B.n683 B.n4 10.6151
R880 B.n684 B.n683 10.6151
R881 B.n685 B.n684 10.6151
R882 B.n685 B.n0 10.6151
R883 B.n619 B.n24 10.6151
R884 B.n619 B.n618 10.6151
R885 B.n618 B.n617 10.6151
R886 B.n617 B.n26 10.6151
R887 B.n613 B.n26 10.6151
R888 B.n613 B.n612 10.6151
R889 B.n612 B.n611 10.6151
R890 B.n611 B.n28 10.6151
R891 B.n607 B.n28 10.6151
R892 B.n607 B.n606 10.6151
R893 B.n606 B.n605 10.6151
R894 B.n605 B.n30 10.6151
R895 B.n601 B.n30 10.6151
R896 B.n601 B.n600 10.6151
R897 B.n600 B.n599 10.6151
R898 B.n599 B.n32 10.6151
R899 B.n595 B.n32 10.6151
R900 B.n595 B.n594 10.6151
R901 B.n594 B.n593 10.6151
R902 B.n593 B.n34 10.6151
R903 B.n589 B.n34 10.6151
R904 B.n589 B.n588 10.6151
R905 B.n588 B.n587 10.6151
R906 B.n587 B.n36 10.6151
R907 B.n583 B.n36 10.6151
R908 B.n583 B.n582 10.6151
R909 B.n582 B.n581 10.6151
R910 B.n581 B.n38 10.6151
R911 B.n577 B.n38 10.6151
R912 B.n577 B.n576 10.6151
R913 B.n576 B.n575 10.6151
R914 B.n575 B.n40 10.6151
R915 B.n571 B.n40 10.6151
R916 B.n571 B.n570 10.6151
R917 B.n568 B.n44 10.6151
R918 B.n564 B.n44 10.6151
R919 B.n564 B.n563 10.6151
R920 B.n563 B.n562 10.6151
R921 B.n562 B.n46 10.6151
R922 B.n558 B.n46 10.6151
R923 B.n558 B.n557 10.6151
R924 B.n557 B.n556 10.6151
R925 B.n556 B.n48 10.6151
R926 B.n552 B.n551 10.6151
R927 B.n551 B.n550 10.6151
R928 B.n550 B.n53 10.6151
R929 B.n546 B.n53 10.6151
R930 B.n546 B.n545 10.6151
R931 B.n545 B.n544 10.6151
R932 B.n544 B.n55 10.6151
R933 B.n540 B.n55 10.6151
R934 B.n540 B.n539 10.6151
R935 B.n539 B.n538 10.6151
R936 B.n538 B.n57 10.6151
R937 B.n534 B.n57 10.6151
R938 B.n534 B.n533 10.6151
R939 B.n533 B.n532 10.6151
R940 B.n532 B.n59 10.6151
R941 B.n528 B.n59 10.6151
R942 B.n528 B.n527 10.6151
R943 B.n527 B.n526 10.6151
R944 B.n526 B.n61 10.6151
R945 B.n522 B.n61 10.6151
R946 B.n522 B.n521 10.6151
R947 B.n521 B.n520 10.6151
R948 B.n520 B.n63 10.6151
R949 B.n516 B.n63 10.6151
R950 B.n516 B.n515 10.6151
R951 B.n515 B.n514 10.6151
R952 B.n514 B.n65 10.6151
R953 B.n510 B.n65 10.6151
R954 B.n510 B.n509 10.6151
R955 B.n509 B.n508 10.6151
R956 B.n508 B.n67 10.6151
R957 B.n504 B.n67 10.6151
R958 B.n504 B.n503 10.6151
R959 B.n503 B.n502 10.6151
R960 B.n498 B.n69 10.6151
R961 B.n498 B.n497 10.6151
R962 B.n497 B.n496 10.6151
R963 B.n496 B.n71 10.6151
R964 B.n492 B.n71 10.6151
R965 B.n492 B.n491 10.6151
R966 B.n491 B.n490 10.6151
R967 B.n490 B.n73 10.6151
R968 B.n486 B.n73 10.6151
R969 B.n486 B.n485 10.6151
R970 B.n485 B.n484 10.6151
R971 B.n484 B.n75 10.6151
R972 B.n480 B.n75 10.6151
R973 B.n480 B.n479 10.6151
R974 B.n479 B.n478 10.6151
R975 B.n478 B.n77 10.6151
R976 B.n474 B.n77 10.6151
R977 B.n474 B.n473 10.6151
R978 B.n473 B.n472 10.6151
R979 B.n472 B.n79 10.6151
R980 B.n468 B.n79 10.6151
R981 B.n468 B.n467 10.6151
R982 B.n467 B.n466 10.6151
R983 B.n466 B.n81 10.6151
R984 B.n462 B.n81 10.6151
R985 B.n462 B.n461 10.6151
R986 B.n461 B.n460 10.6151
R987 B.n460 B.n83 10.6151
R988 B.n456 B.n83 10.6151
R989 B.n456 B.n455 10.6151
R990 B.n455 B.n454 10.6151
R991 B.n454 B.n85 10.6151
R992 B.n450 B.n85 10.6151
R993 B.n450 B.n449 10.6151
R994 B.n449 B.n448 10.6151
R995 B.n448 B.n87 10.6151
R996 B.n444 B.n87 10.6151
R997 B.n444 B.n443 10.6151
R998 B.n443 B.n442 10.6151
R999 B.n442 B.n89 10.6151
R1000 B.n438 B.n89 10.6151
R1001 B.n438 B.n437 10.6151
R1002 B.n437 B.n436 10.6151
R1003 B.n436 B.n91 10.6151
R1004 B.n432 B.n91 10.6151
R1005 B.n432 B.n431 10.6151
R1006 B.n431 B.n430 10.6151
R1007 B.n430 B.n93 10.6151
R1008 B.n426 B.n93 10.6151
R1009 B.n426 B.n425 10.6151
R1010 B.n425 B.n424 10.6151
R1011 B.n424 B.n95 10.6151
R1012 B.n420 B.n95 10.6151
R1013 B.n420 B.n419 10.6151
R1014 B.n419 B.n418 10.6151
R1015 B.n418 B.n97 10.6151
R1016 B.n414 B.n97 10.6151
R1017 B.n414 B.n413 10.6151
R1018 B.n413 B.n412 10.6151
R1019 B.n412 B.n99 10.6151
R1020 B.n408 B.n99 10.6151
R1021 B.n408 B.n407 10.6151
R1022 B.n407 B.n406 10.6151
R1023 B.n406 B.n101 10.6151
R1024 B.n402 B.n101 10.6151
R1025 B.n402 B.n401 10.6151
R1026 B.n401 B.n400 10.6151
R1027 B.n400 B.n103 10.6151
R1028 B.n396 B.n103 10.6151
R1029 B.n396 B.n395 10.6151
R1030 B.n395 B.n394 10.6151
R1031 B.n394 B.n105 10.6151
R1032 B.n390 B.n105 10.6151
R1033 B.n390 B.n389 10.6151
R1034 B.n389 B.n388 10.6151
R1035 B.n388 B.n107 10.6151
R1036 B.n384 B.n107 10.6151
R1037 B.n384 B.n383 10.6151
R1038 B.n383 B.n382 10.6151
R1039 B.n382 B.n109 10.6151
R1040 B.n378 B.n109 10.6151
R1041 B.n378 B.n377 10.6151
R1042 B.n377 B.n376 10.6151
R1043 B.n376 B.n111 10.6151
R1044 B.n372 B.n111 10.6151
R1045 B.n372 B.n371 10.6151
R1046 B.n371 B.n370 10.6151
R1047 B.n370 B.n113 10.6151
R1048 B.n366 B.n113 10.6151
R1049 B.n177 B.n1 10.6151
R1050 B.n180 B.n177 10.6151
R1051 B.n181 B.n180 10.6151
R1052 B.n182 B.n181 10.6151
R1053 B.n182 B.n175 10.6151
R1054 B.n186 B.n175 10.6151
R1055 B.n187 B.n186 10.6151
R1056 B.n188 B.n187 10.6151
R1057 B.n188 B.n173 10.6151
R1058 B.n192 B.n173 10.6151
R1059 B.n193 B.n192 10.6151
R1060 B.n194 B.n193 10.6151
R1061 B.n194 B.n171 10.6151
R1062 B.n198 B.n171 10.6151
R1063 B.n199 B.n198 10.6151
R1064 B.n200 B.n199 10.6151
R1065 B.n200 B.n169 10.6151
R1066 B.n204 B.n169 10.6151
R1067 B.n205 B.n204 10.6151
R1068 B.n206 B.n205 10.6151
R1069 B.n206 B.n167 10.6151
R1070 B.n210 B.n167 10.6151
R1071 B.n211 B.n210 10.6151
R1072 B.n212 B.n211 10.6151
R1073 B.n212 B.n165 10.6151
R1074 B.n216 B.n165 10.6151
R1075 B.n217 B.n216 10.6151
R1076 B.n218 B.n217 10.6151
R1077 B.n218 B.n163 10.6151
R1078 B.n222 B.n163 10.6151
R1079 B.n223 B.n222 10.6151
R1080 B.n224 B.n223 10.6151
R1081 B.n224 B.n161 10.6151
R1082 B.n228 B.n161 10.6151
R1083 B.n229 B.n228 10.6151
R1084 B.n230 B.n229 10.6151
R1085 B.n230 B.n159 10.6151
R1086 B.n234 B.n159 10.6151
R1087 B.n235 B.n234 10.6151
R1088 B.n236 B.n235 10.6151
R1089 B.n236 B.n157 10.6151
R1090 B.n240 B.n157 10.6151
R1091 B.n241 B.n240 10.6151
R1092 B.n242 B.n155 10.6151
R1093 B.n246 B.n155 10.6151
R1094 B.n247 B.n246 10.6151
R1095 B.n248 B.n247 10.6151
R1096 B.n248 B.n153 10.6151
R1097 B.n252 B.n153 10.6151
R1098 B.n253 B.n252 10.6151
R1099 B.n254 B.n253 10.6151
R1100 B.n254 B.n151 10.6151
R1101 B.n258 B.n151 10.6151
R1102 B.n259 B.n258 10.6151
R1103 B.n260 B.n259 10.6151
R1104 B.n260 B.n149 10.6151
R1105 B.n264 B.n149 10.6151
R1106 B.n265 B.n264 10.6151
R1107 B.n266 B.n265 10.6151
R1108 B.n266 B.n147 10.6151
R1109 B.n270 B.n147 10.6151
R1110 B.n271 B.n270 10.6151
R1111 B.n272 B.n271 10.6151
R1112 B.n272 B.n145 10.6151
R1113 B.n276 B.n145 10.6151
R1114 B.n277 B.n276 10.6151
R1115 B.n278 B.n277 10.6151
R1116 B.n278 B.n143 10.6151
R1117 B.n282 B.n143 10.6151
R1118 B.n283 B.n282 10.6151
R1119 B.n284 B.n283 10.6151
R1120 B.n284 B.n141 10.6151
R1121 B.n288 B.n141 10.6151
R1122 B.n289 B.n288 10.6151
R1123 B.n290 B.n289 10.6151
R1124 B.n290 B.n139 10.6151
R1125 B.n294 B.n139 10.6151
R1126 B.n297 B.n296 10.6151
R1127 B.n297 B.n135 10.6151
R1128 B.n301 B.n135 10.6151
R1129 B.n302 B.n301 10.6151
R1130 B.n303 B.n302 10.6151
R1131 B.n303 B.n133 10.6151
R1132 B.n307 B.n133 10.6151
R1133 B.n308 B.n307 10.6151
R1134 B.n312 B.n308 10.6151
R1135 B.n316 B.n131 10.6151
R1136 B.n317 B.n316 10.6151
R1137 B.n318 B.n317 10.6151
R1138 B.n318 B.n129 10.6151
R1139 B.n322 B.n129 10.6151
R1140 B.n323 B.n322 10.6151
R1141 B.n324 B.n323 10.6151
R1142 B.n324 B.n127 10.6151
R1143 B.n328 B.n127 10.6151
R1144 B.n329 B.n328 10.6151
R1145 B.n330 B.n329 10.6151
R1146 B.n330 B.n125 10.6151
R1147 B.n334 B.n125 10.6151
R1148 B.n335 B.n334 10.6151
R1149 B.n336 B.n335 10.6151
R1150 B.n336 B.n123 10.6151
R1151 B.n340 B.n123 10.6151
R1152 B.n341 B.n340 10.6151
R1153 B.n342 B.n341 10.6151
R1154 B.n342 B.n121 10.6151
R1155 B.n346 B.n121 10.6151
R1156 B.n347 B.n346 10.6151
R1157 B.n348 B.n347 10.6151
R1158 B.n348 B.n119 10.6151
R1159 B.n352 B.n119 10.6151
R1160 B.n353 B.n352 10.6151
R1161 B.n354 B.n353 10.6151
R1162 B.n354 B.n117 10.6151
R1163 B.n358 B.n117 10.6151
R1164 B.n359 B.n358 10.6151
R1165 B.n360 B.n359 10.6151
R1166 B.n360 B.n115 10.6151
R1167 B.n364 B.n115 10.6151
R1168 B.n365 B.n364 10.6151
R1169 B.n570 B.n569 9.36635
R1170 B.n552 B.n52 9.36635
R1171 B.n295 B.n294 9.36635
R1172 B.n311 B.n131 9.36635
R1173 B.n689 B.n0 8.11757
R1174 B.n689 B.n1 8.11757
R1175 B.n569 B.n568 1.24928
R1176 B.n52 B.n48 1.24928
R1177 B.n296 B.n295 1.24928
R1178 B.n312 B.n311 1.24928
R1179 VN.n43 VN.n23 161.3
R1180 VN.n42 VN.n41 161.3
R1181 VN.n40 VN.n24 161.3
R1182 VN.n39 VN.n38 161.3
R1183 VN.n37 VN.n25 161.3
R1184 VN.n35 VN.n34 161.3
R1185 VN.n33 VN.n26 161.3
R1186 VN.n32 VN.n31 161.3
R1187 VN.n30 VN.n27 161.3
R1188 VN.n20 VN.n0 161.3
R1189 VN.n19 VN.n18 161.3
R1190 VN.n17 VN.n1 161.3
R1191 VN.n16 VN.n15 161.3
R1192 VN.n14 VN.n2 161.3
R1193 VN.n12 VN.n11 161.3
R1194 VN.n10 VN.n3 161.3
R1195 VN.n9 VN.n8 161.3
R1196 VN.n7 VN.n4 161.3
R1197 VN.n5 VN.t6 144.333
R1198 VN.n28 VN.t4 144.333
R1199 VN.n6 VN.t5 109.74
R1200 VN.n13 VN.t3 109.74
R1201 VN.n21 VN.t1 109.74
R1202 VN.n29 VN.t2 109.74
R1203 VN.n36 VN.t0 109.74
R1204 VN.n44 VN.t7 109.74
R1205 VN.n22 VN.n21 87.7575
R1206 VN.n45 VN.n44 87.7575
R1207 VN.n8 VN.n3 56.5193
R1208 VN.n19 VN.n1 56.5193
R1209 VN.n31 VN.n26 56.5193
R1210 VN.n42 VN.n24 56.5193
R1211 VN VN.n45 47.5057
R1212 VN.n6 VN.n5 46.8391
R1213 VN.n29 VN.n28 46.8391
R1214 VN.n8 VN.n7 24.4675
R1215 VN.n12 VN.n3 24.4675
R1216 VN.n15 VN.n14 24.4675
R1217 VN.n15 VN.n1 24.4675
R1218 VN.n20 VN.n19 24.4675
R1219 VN.n31 VN.n30 24.4675
R1220 VN.n38 VN.n24 24.4675
R1221 VN.n38 VN.n37 24.4675
R1222 VN.n35 VN.n26 24.4675
R1223 VN.n43 VN.n42 24.4675
R1224 VN.n7 VN.n6 23.9782
R1225 VN.n13 VN.n12 23.9782
R1226 VN.n30 VN.n29 23.9782
R1227 VN.n36 VN.n35 23.9782
R1228 VN.n21 VN.n20 22.9995
R1229 VN.n44 VN.n43 22.9995
R1230 VN.n28 VN.n27 8.69054
R1231 VN.n5 VN.n4 8.69054
R1232 VN.n14 VN.n13 0.48984
R1233 VN.n37 VN.n36 0.48984
R1234 VN.n45 VN.n23 0.278367
R1235 VN.n22 VN.n0 0.278367
R1236 VN.n41 VN.n23 0.189894
R1237 VN.n41 VN.n40 0.189894
R1238 VN.n40 VN.n39 0.189894
R1239 VN.n39 VN.n25 0.189894
R1240 VN.n34 VN.n25 0.189894
R1241 VN.n34 VN.n33 0.189894
R1242 VN.n33 VN.n32 0.189894
R1243 VN.n32 VN.n27 0.189894
R1244 VN.n9 VN.n4 0.189894
R1245 VN.n10 VN.n9 0.189894
R1246 VN.n11 VN.n10 0.189894
R1247 VN.n11 VN.n2 0.189894
R1248 VN.n16 VN.n2 0.189894
R1249 VN.n17 VN.n16 0.189894
R1250 VN.n18 VN.n17 0.189894
R1251 VN.n18 VN.n0 0.189894
R1252 VN VN.n22 0.153454
R1253 VDD2.n2 VDD2.n1 82.5186
R1254 VDD2.n2 VDD2.n0 82.5186
R1255 VDD2 VDD2.n5 82.5158
R1256 VDD2.n4 VDD2.n3 81.5052
R1257 VDD2.n4 VDD2.n2 41.7756
R1258 VDD2.n5 VDD2.t5 3.32072
R1259 VDD2.n5 VDD2.t3 3.32072
R1260 VDD2.n3 VDD2.t0 3.32072
R1261 VDD2.n3 VDD2.t7 3.32072
R1262 VDD2.n1 VDD2.t4 3.32072
R1263 VDD2.n1 VDD2.t6 3.32072
R1264 VDD2.n0 VDD2.t1 3.32072
R1265 VDD2.n0 VDD2.t2 3.32072
R1266 VDD2 VDD2.n4 1.12766
C0 VN B 1.0946f
C1 VTAIL VDD2 7.29191f
C2 VDD2 B 1.53553f
C3 w_n3450_n2926# VP 7.28898f
C4 VN VDD1 0.151005f
C5 VP VTAIL 7.24478f
C6 VP B 1.84078f
C7 VDD2 VDD1 1.54385f
C8 VP VDD1 7.20378f
C9 VN VDD2 6.88407f
C10 VP VN 6.70011f
C11 VP VDD2 0.471877f
C12 w_n3450_n2926# VTAIL 3.67977f
C13 w_n3450_n2926# B 8.806951f
C14 VTAIL B 4.06232f
C15 w_n3450_n2926# VDD1 1.75128f
C16 VTAIL VDD1 7.24051f
C17 VDD1 B 1.45366f
C18 w_n3450_n2926# VN 6.84243f
C19 VN VTAIL 7.23068f
C20 w_n3450_n2926# VDD2 1.84711f
C21 VDD2 VSUBS 1.592822f
C22 VDD1 VSUBS 2.158953f
C23 VTAIL VSUBS 1.156383f
C24 VN VSUBS 6.09186f
C25 VP VSUBS 3.053991f
C26 B VSUBS 4.311013f
C27 w_n3450_n2926# VSUBS 0.124738p
C28 VDD2.t1 VSUBS 0.189404f
C29 VDD2.t2 VSUBS 0.189404f
C30 VDD2.n0 VSUBS 1.44237f
C31 VDD2.t4 VSUBS 0.189404f
C32 VDD2.t6 VSUBS 0.189404f
C33 VDD2.n1 VSUBS 1.44237f
C34 VDD2.n2 VSUBS 3.27629f
C35 VDD2.t0 VSUBS 0.189404f
C36 VDD2.t7 VSUBS 0.189404f
C37 VDD2.n3 VSUBS 1.4339f
C38 VDD2.n4 VSUBS 2.79841f
C39 VDD2.t5 VSUBS 0.189404f
C40 VDD2.t3 VSUBS 0.189404f
C41 VDD2.n5 VSUBS 1.44234f
C42 VN.n0 VSUBS 0.044614f
C43 VN.t1 VSUBS 1.92814f
C44 VN.n1 VSUBS 0.047513f
C45 VN.n2 VSUBS 0.033839f
C46 VN.t3 VSUBS 1.92814f
C47 VN.n3 VSUBS 0.049399f
C48 VN.n4 VSUBS 0.285735f
C49 VN.t5 VSUBS 1.92814f
C50 VN.t6 VSUBS 2.14066f
C51 VN.n5 VSUBS 0.768045f
C52 VN.n6 VSUBS 0.798956f
C53 VN.n7 VSUBS 0.062445f
C54 VN.n8 VSUBS 0.049399f
C55 VN.n9 VSUBS 0.033839f
C56 VN.n10 VSUBS 0.033839f
C57 VN.n11 VSUBS 0.033839f
C58 VN.n12 VSUBS 0.062445f
C59 VN.n13 VSUBS 0.696504f
C60 VN.n14 VSUBS 0.032554f
C61 VN.n15 VSUBS 0.063068f
C62 VN.n16 VSUBS 0.033839f
C63 VN.n17 VSUBS 0.033839f
C64 VN.n18 VSUBS 0.033839f
C65 VN.n19 VSUBS 0.051285f
C66 VN.n20 VSUBS 0.0612f
C67 VN.n21 VSUBS 0.814951f
C68 VN.n22 VSUBS 0.038242f
C69 VN.n23 VSUBS 0.044614f
C70 VN.t7 VSUBS 1.92814f
C71 VN.n24 VSUBS 0.047513f
C72 VN.n25 VSUBS 0.033839f
C73 VN.t0 VSUBS 1.92814f
C74 VN.n26 VSUBS 0.049399f
C75 VN.n27 VSUBS 0.285735f
C76 VN.t2 VSUBS 1.92814f
C77 VN.t4 VSUBS 2.14066f
C78 VN.n28 VSUBS 0.768045f
C79 VN.n29 VSUBS 0.798956f
C80 VN.n30 VSUBS 0.062445f
C81 VN.n31 VSUBS 0.049399f
C82 VN.n32 VSUBS 0.033839f
C83 VN.n33 VSUBS 0.033839f
C84 VN.n34 VSUBS 0.033839f
C85 VN.n35 VSUBS 0.062445f
C86 VN.n36 VSUBS 0.696504f
C87 VN.n37 VSUBS 0.032554f
C88 VN.n38 VSUBS 0.063068f
C89 VN.n39 VSUBS 0.033839f
C90 VN.n40 VSUBS 0.033839f
C91 VN.n41 VSUBS 0.033839f
C92 VN.n42 VSUBS 0.051285f
C93 VN.n43 VSUBS 0.0612f
C94 VN.n44 VSUBS 0.814951f
C95 VN.n45 VSUBS 1.73163f
C96 B.n0 VSUBS 0.006471f
C97 B.n1 VSUBS 0.006471f
C98 B.n2 VSUBS 0.009571f
C99 B.n3 VSUBS 0.007334f
C100 B.n4 VSUBS 0.007334f
C101 B.n5 VSUBS 0.007334f
C102 B.n6 VSUBS 0.007334f
C103 B.n7 VSUBS 0.007334f
C104 B.n8 VSUBS 0.007334f
C105 B.n9 VSUBS 0.007334f
C106 B.n10 VSUBS 0.007334f
C107 B.n11 VSUBS 0.007334f
C108 B.n12 VSUBS 0.007334f
C109 B.n13 VSUBS 0.007334f
C110 B.n14 VSUBS 0.007334f
C111 B.n15 VSUBS 0.007334f
C112 B.n16 VSUBS 0.007334f
C113 B.n17 VSUBS 0.007334f
C114 B.n18 VSUBS 0.007334f
C115 B.n19 VSUBS 0.007334f
C116 B.n20 VSUBS 0.007334f
C117 B.n21 VSUBS 0.007334f
C118 B.n22 VSUBS 0.007334f
C119 B.n23 VSUBS 0.007334f
C120 B.n24 VSUBS 0.017586f
C121 B.n25 VSUBS 0.007334f
C122 B.n26 VSUBS 0.007334f
C123 B.n27 VSUBS 0.007334f
C124 B.n28 VSUBS 0.007334f
C125 B.n29 VSUBS 0.007334f
C126 B.n30 VSUBS 0.007334f
C127 B.n31 VSUBS 0.007334f
C128 B.n32 VSUBS 0.007334f
C129 B.n33 VSUBS 0.007334f
C130 B.n34 VSUBS 0.007334f
C131 B.n35 VSUBS 0.007334f
C132 B.n36 VSUBS 0.007334f
C133 B.n37 VSUBS 0.007334f
C134 B.n38 VSUBS 0.007334f
C135 B.n39 VSUBS 0.007334f
C136 B.n40 VSUBS 0.007334f
C137 B.n41 VSUBS 0.007334f
C138 B.t10 VSUBS 0.326185f
C139 B.t11 VSUBS 0.344888f
C140 B.t9 VSUBS 1.00419f
C141 B.n42 VSUBS 0.174407f
C142 B.n43 VSUBS 0.073096f
C143 B.n44 VSUBS 0.007334f
C144 B.n45 VSUBS 0.007334f
C145 B.n46 VSUBS 0.007334f
C146 B.n47 VSUBS 0.007334f
C147 B.n48 VSUBS 0.004098f
C148 B.n49 VSUBS 0.007334f
C149 B.t7 VSUBS 0.326181f
C150 B.t8 VSUBS 0.344883f
C151 B.t6 VSUBS 1.00419f
C152 B.n50 VSUBS 0.174411f
C153 B.n51 VSUBS 0.0731f
C154 B.n52 VSUBS 0.016992f
C155 B.n53 VSUBS 0.007334f
C156 B.n54 VSUBS 0.007334f
C157 B.n55 VSUBS 0.007334f
C158 B.n56 VSUBS 0.007334f
C159 B.n57 VSUBS 0.007334f
C160 B.n58 VSUBS 0.007334f
C161 B.n59 VSUBS 0.007334f
C162 B.n60 VSUBS 0.007334f
C163 B.n61 VSUBS 0.007334f
C164 B.n62 VSUBS 0.007334f
C165 B.n63 VSUBS 0.007334f
C166 B.n64 VSUBS 0.007334f
C167 B.n65 VSUBS 0.007334f
C168 B.n66 VSUBS 0.007334f
C169 B.n67 VSUBS 0.007334f
C170 B.n68 VSUBS 0.007334f
C171 B.n69 VSUBS 0.016496f
C172 B.n70 VSUBS 0.007334f
C173 B.n71 VSUBS 0.007334f
C174 B.n72 VSUBS 0.007334f
C175 B.n73 VSUBS 0.007334f
C176 B.n74 VSUBS 0.007334f
C177 B.n75 VSUBS 0.007334f
C178 B.n76 VSUBS 0.007334f
C179 B.n77 VSUBS 0.007334f
C180 B.n78 VSUBS 0.007334f
C181 B.n79 VSUBS 0.007334f
C182 B.n80 VSUBS 0.007334f
C183 B.n81 VSUBS 0.007334f
C184 B.n82 VSUBS 0.007334f
C185 B.n83 VSUBS 0.007334f
C186 B.n84 VSUBS 0.007334f
C187 B.n85 VSUBS 0.007334f
C188 B.n86 VSUBS 0.007334f
C189 B.n87 VSUBS 0.007334f
C190 B.n88 VSUBS 0.007334f
C191 B.n89 VSUBS 0.007334f
C192 B.n90 VSUBS 0.007334f
C193 B.n91 VSUBS 0.007334f
C194 B.n92 VSUBS 0.007334f
C195 B.n93 VSUBS 0.007334f
C196 B.n94 VSUBS 0.007334f
C197 B.n95 VSUBS 0.007334f
C198 B.n96 VSUBS 0.007334f
C199 B.n97 VSUBS 0.007334f
C200 B.n98 VSUBS 0.007334f
C201 B.n99 VSUBS 0.007334f
C202 B.n100 VSUBS 0.007334f
C203 B.n101 VSUBS 0.007334f
C204 B.n102 VSUBS 0.007334f
C205 B.n103 VSUBS 0.007334f
C206 B.n104 VSUBS 0.007334f
C207 B.n105 VSUBS 0.007334f
C208 B.n106 VSUBS 0.007334f
C209 B.n107 VSUBS 0.007334f
C210 B.n108 VSUBS 0.007334f
C211 B.n109 VSUBS 0.007334f
C212 B.n110 VSUBS 0.007334f
C213 B.n111 VSUBS 0.007334f
C214 B.n112 VSUBS 0.007334f
C215 B.n113 VSUBS 0.007334f
C216 B.n114 VSUBS 0.017586f
C217 B.n115 VSUBS 0.007334f
C218 B.n116 VSUBS 0.007334f
C219 B.n117 VSUBS 0.007334f
C220 B.n118 VSUBS 0.007334f
C221 B.n119 VSUBS 0.007334f
C222 B.n120 VSUBS 0.007334f
C223 B.n121 VSUBS 0.007334f
C224 B.n122 VSUBS 0.007334f
C225 B.n123 VSUBS 0.007334f
C226 B.n124 VSUBS 0.007334f
C227 B.n125 VSUBS 0.007334f
C228 B.n126 VSUBS 0.007334f
C229 B.n127 VSUBS 0.007334f
C230 B.n128 VSUBS 0.007334f
C231 B.n129 VSUBS 0.007334f
C232 B.n130 VSUBS 0.007334f
C233 B.n131 VSUBS 0.006903f
C234 B.n132 VSUBS 0.007334f
C235 B.n133 VSUBS 0.007334f
C236 B.n134 VSUBS 0.007334f
C237 B.n135 VSUBS 0.007334f
C238 B.n136 VSUBS 0.007334f
C239 B.t5 VSUBS 0.326185f
C240 B.t4 VSUBS 0.344888f
C241 B.t3 VSUBS 1.00419f
C242 B.n137 VSUBS 0.174407f
C243 B.n138 VSUBS 0.073096f
C244 B.n139 VSUBS 0.007334f
C245 B.n140 VSUBS 0.007334f
C246 B.n141 VSUBS 0.007334f
C247 B.n142 VSUBS 0.007334f
C248 B.n143 VSUBS 0.007334f
C249 B.n144 VSUBS 0.007334f
C250 B.n145 VSUBS 0.007334f
C251 B.n146 VSUBS 0.007334f
C252 B.n147 VSUBS 0.007334f
C253 B.n148 VSUBS 0.007334f
C254 B.n149 VSUBS 0.007334f
C255 B.n150 VSUBS 0.007334f
C256 B.n151 VSUBS 0.007334f
C257 B.n152 VSUBS 0.007334f
C258 B.n153 VSUBS 0.007334f
C259 B.n154 VSUBS 0.007334f
C260 B.n155 VSUBS 0.007334f
C261 B.n156 VSUBS 0.016496f
C262 B.n157 VSUBS 0.007334f
C263 B.n158 VSUBS 0.007334f
C264 B.n159 VSUBS 0.007334f
C265 B.n160 VSUBS 0.007334f
C266 B.n161 VSUBS 0.007334f
C267 B.n162 VSUBS 0.007334f
C268 B.n163 VSUBS 0.007334f
C269 B.n164 VSUBS 0.007334f
C270 B.n165 VSUBS 0.007334f
C271 B.n166 VSUBS 0.007334f
C272 B.n167 VSUBS 0.007334f
C273 B.n168 VSUBS 0.007334f
C274 B.n169 VSUBS 0.007334f
C275 B.n170 VSUBS 0.007334f
C276 B.n171 VSUBS 0.007334f
C277 B.n172 VSUBS 0.007334f
C278 B.n173 VSUBS 0.007334f
C279 B.n174 VSUBS 0.007334f
C280 B.n175 VSUBS 0.007334f
C281 B.n176 VSUBS 0.007334f
C282 B.n177 VSUBS 0.007334f
C283 B.n178 VSUBS 0.007334f
C284 B.n179 VSUBS 0.007334f
C285 B.n180 VSUBS 0.007334f
C286 B.n181 VSUBS 0.007334f
C287 B.n182 VSUBS 0.007334f
C288 B.n183 VSUBS 0.007334f
C289 B.n184 VSUBS 0.007334f
C290 B.n185 VSUBS 0.007334f
C291 B.n186 VSUBS 0.007334f
C292 B.n187 VSUBS 0.007334f
C293 B.n188 VSUBS 0.007334f
C294 B.n189 VSUBS 0.007334f
C295 B.n190 VSUBS 0.007334f
C296 B.n191 VSUBS 0.007334f
C297 B.n192 VSUBS 0.007334f
C298 B.n193 VSUBS 0.007334f
C299 B.n194 VSUBS 0.007334f
C300 B.n195 VSUBS 0.007334f
C301 B.n196 VSUBS 0.007334f
C302 B.n197 VSUBS 0.007334f
C303 B.n198 VSUBS 0.007334f
C304 B.n199 VSUBS 0.007334f
C305 B.n200 VSUBS 0.007334f
C306 B.n201 VSUBS 0.007334f
C307 B.n202 VSUBS 0.007334f
C308 B.n203 VSUBS 0.007334f
C309 B.n204 VSUBS 0.007334f
C310 B.n205 VSUBS 0.007334f
C311 B.n206 VSUBS 0.007334f
C312 B.n207 VSUBS 0.007334f
C313 B.n208 VSUBS 0.007334f
C314 B.n209 VSUBS 0.007334f
C315 B.n210 VSUBS 0.007334f
C316 B.n211 VSUBS 0.007334f
C317 B.n212 VSUBS 0.007334f
C318 B.n213 VSUBS 0.007334f
C319 B.n214 VSUBS 0.007334f
C320 B.n215 VSUBS 0.007334f
C321 B.n216 VSUBS 0.007334f
C322 B.n217 VSUBS 0.007334f
C323 B.n218 VSUBS 0.007334f
C324 B.n219 VSUBS 0.007334f
C325 B.n220 VSUBS 0.007334f
C326 B.n221 VSUBS 0.007334f
C327 B.n222 VSUBS 0.007334f
C328 B.n223 VSUBS 0.007334f
C329 B.n224 VSUBS 0.007334f
C330 B.n225 VSUBS 0.007334f
C331 B.n226 VSUBS 0.007334f
C332 B.n227 VSUBS 0.007334f
C333 B.n228 VSUBS 0.007334f
C334 B.n229 VSUBS 0.007334f
C335 B.n230 VSUBS 0.007334f
C336 B.n231 VSUBS 0.007334f
C337 B.n232 VSUBS 0.007334f
C338 B.n233 VSUBS 0.007334f
C339 B.n234 VSUBS 0.007334f
C340 B.n235 VSUBS 0.007334f
C341 B.n236 VSUBS 0.007334f
C342 B.n237 VSUBS 0.007334f
C343 B.n238 VSUBS 0.007334f
C344 B.n239 VSUBS 0.007334f
C345 B.n240 VSUBS 0.007334f
C346 B.n241 VSUBS 0.016496f
C347 B.n242 VSUBS 0.017586f
C348 B.n243 VSUBS 0.017586f
C349 B.n244 VSUBS 0.007334f
C350 B.n245 VSUBS 0.007334f
C351 B.n246 VSUBS 0.007334f
C352 B.n247 VSUBS 0.007334f
C353 B.n248 VSUBS 0.007334f
C354 B.n249 VSUBS 0.007334f
C355 B.n250 VSUBS 0.007334f
C356 B.n251 VSUBS 0.007334f
C357 B.n252 VSUBS 0.007334f
C358 B.n253 VSUBS 0.007334f
C359 B.n254 VSUBS 0.007334f
C360 B.n255 VSUBS 0.007334f
C361 B.n256 VSUBS 0.007334f
C362 B.n257 VSUBS 0.007334f
C363 B.n258 VSUBS 0.007334f
C364 B.n259 VSUBS 0.007334f
C365 B.n260 VSUBS 0.007334f
C366 B.n261 VSUBS 0.007334f
C367 B.n262 VSUBS 0.007334f
C368 B.n263 VSUBS 0.007334f
C369 B.n264 VSUBS 0.007334f
C370 B.n265 VSUBS 0.007334f
C371 B.n266 VSUBS 0.007334f
C372 B.n267 VSUBS 0.007334f
C373 B.n268 VSUBS 0.007334f
C374 B.n269 VSUBS 0.007334f
C375 B.n270 VSUBS 0.007334f
C376 B.n271 VSUBS 0.007334f
C377 B.n272 VSUBS 0.007334f
C378 B.n273 VSUBS 0.007334f
C379 B.n274 VSUBS 0.007334f
C380 B.n275 VSUBS 0.007334f
C381 B.n276 VSUBS 0.007334f
C382 B.n277 VSUBS 0.007334f
C383 B.n278 VSUBS 0.007334f
C384 B.n279 VSUBS 0.007334f
C385 B.n280 VSUBS 0.007334f
C386 B.n281 VSUBS 0.007334f
C387 B.n282 VSUBS 0.007334f
C388 B.n283 VSUBS 0.007334f
C389 B.n284 VSUBS 0.007334f
C390 B.n285 VSUBS 0.007334f
C391 B.n286 VSUBS 0.007334f
C392 B.n287 VSUBS 0.007334f
C393 B.n288 VSUBS 0.007334f
C394 B.n289 VSUBS 0.007334f
C395 B.n290 VSUBS 0.007334f
C396 B.n291 VSUBS 0.007334f
C397 B.n292 VSUBS 0.007334f
C398 B.n293 VSUBS 0.007334f
C399 B.n294 VSUBS 0.006903f
C400 B.n295 VSUBS 0.016992f
C401 B.n296 VSUBS 0.004098f
C402 B.n297 VSUBS 0.007334f
C403 B.n298 VSUBS 0.007334f
C404 B.n299 VSUBS 0.007334f
C405 B.n300 VSUBS 0.007334f
C406 B.n301 VSUBS 0.007334f
C407 B.n302 VSUBS 0.007334f
C408 B.n303 VSUBS 0.007334f
C409 B.n304 VSUBS 0.007334f
C410 B.n305 VSUBS 0.007334f
C411 B.n306 VSUBS 0.007334f
C412 B.n307 VSUBS 0.007334f
C413 B.n308 VSUBS 0.007334f
C414 B.t2 VSUBS 0.326181f
C415 B.t1 VSUBS 0.344883f
C416 B.t0 VSUBS 1.00419f
C417 B.n309 VSUBS 0.174411f
C418 B.n310 VSUBS 0.0731f
C419 B.n311 VSUBS 0.016992f
C420 B.n312 VSUBS 0.004098f
C421 B.n313 VSUBS 0.007334f
C422 B.n314 VSUBS 0.007334f
C423 B.n315 VSUBS 0.007334f
C424 B.n316 VSUBS 0.007334f
C425 B.n317 VSUBS 0.007334f
C426 B.n318 VSUBS 0.007334f
C427 B.n319 VSUBS 0.007334f
C428 B.n320 VSUBS 0.007334f
C429 B.n321 VSUBS 0.007334f
C430 B.n322 VSUBS 0.007334f
C431 B.n323 VSUBS 0.007334f
C432 B.n324 VSUBS 0.007334f
C433 B.n325 VSUBS 0.007334f
C434 B.n326 VSUBS 0.007334f
C435 B.n327 VSUBS 0.007334f
C436 B.n328 VSUBS 0.007334f
C437 B.n329 VSUBS 0.007334f
C438 B.n330 VSUBS 0.007334f
C439 B.n331 VSUBS 0.007334f
C440 B.n332 VSUBS 0.007334f
C441 B.n333 VSUBS 0.007334f
C442 B.n334 VSUBS 0.007334f
C443 B.n335 VSUBS 0.007334f
C444 B.n336 VSUBS 0.007334f
C445 B.n337 VSUBS 0.007334f
C446 B.n338 VSUBS 0.007334f
C447 B.n339 VSUBS 0.007334f
C448 B.n340 VSUBS 0.007334f
C449 B.n341 VSUBS 0.007334f
C450 B.n342 VSUBS 0.007334f
C451 B.n343 VSUBS 0.007334f
C452 B.n344 VSUBS 0.007334f
C453 B.n345 VSUBS 0.007334f
C454 B.n346 VSUBS 0.007334f
C455 B.n347 VSUBS 0.007334f
C456 B.n348 VSUBS 0.007334f
C457 B.n349 VSUBS 0.007334f
C458 B.n350 VSUBS 0.007334f
C459 B.n351 VSUBS 0.007334f
C460 B.n352 VSUBS 0.007334f
C461 B.n353 VSUBS 0.007334f
C462 B.n354 VSUBS 0.007334f
C463 B.n355 VSUBS 0.007334f
C464 B.n356 VSUBS 0.007334f
C465 B.n357 VSUBS 0.007334f
C466 B.n358 VSUBS 0.007334f
C467 B.n359 VSUBS 0.007334f
C468 B.n360 VSUBS 0.007334f
C469 B.n361 VSUBS 0.007334f
C470 B.n362 VSUBS 0.007334f
C471 B.n363 VSUBS 0.007334f
C472 B.n364 VSUBS 0.007334f
C473 B.n365 VSUBS 0.01671f
C474 B.n366 VSUBS 0.017372f
C475 B.n367 VSUBS 0.016496f
C476 B.n368 VSUBS 0.007334f
C477 B.n369 VSUBS 0.007334f
C478 B.n370 VSUBS 0.007334f
C479 B.n371 VSUBS 0.007334f
C480 B.n372 VSUBS 0.007334f
C481 B.n373 VSUBS 0.007334f
C482 B.n374 VSUBS 0.007334f
C483 B.n375 VSUBS 0.007334f
C484 B.n376 VSUBS 0.007334f
C485 B.n377 VSUBS 0.007334f
C486 B.n378 VSUBS 0.007334f
C487 B.n379 VSUBS 0.007334f
C488 B.n380 VSUBS 0.007334f
C489 B.n381 VSUBS 0.007334f
C490 B.n382 VSUBS 0.007334f
C491 B.n383 VSUBS 0.007334f
C492 B.n384 VSUBS 0.007334f
C493 B.n385 VSUBS 0.007334f
C494 B.n386 VSUBS 0.007334f
C495 B.n387 VSUBS 0.007334f
C496 B.n388 VSUBS 0.007334f
C497 B.n389 VSUBS 0.007334f
C498 B.n390 VSUBS 0.007334f
C499 B.n391 VSUBS 0.007334f
C500 B.n392 VSUBS 0.007334f
C501 B.n393 VSUBS 0.007334f
C502 B.n394 VSUBS 0.007334f
C503 B.n395 VSUBS 0.007334f
C504 B.n396 VSUBS 0.007334f
C505 B.n397 VSUBS 0.007334f
C506 B.n398 VSUBS 0.007334f
C507 B.n399 VSUBS 0.007334f
C508 B.n400 VSUBS 0.007334f
C509 B.n401 VSUBS 0.007334f
C510 B.n402 VSUBS 0.007334f
C511 B.n403 VSUBS 0.007334f
C512 B.n404 VSUBS 0.007334f
C513 B.n405 VSUBS 0.007334f
C514 B.n406 VSUBS 0.007334f
C515 B.n407 VSUBS 0.007334f
C516 B.n408 VSUBS 0.007334f
C517 B.n409 VSUBS 0.007334f
C518 B.n410 VSUBS 0.007334f
C519 B.n411 VSUBS 0.007334f
C520 B.n412 VSUBS 0.007334f
C521 B.n413 VSUBS 0.007334f
C522 B.n414 VSUBS 0.007334f
C523 B.n415 VSUBS 0.007334f
C524 B.n416 VSUBS 0.007334f
C525 B.n417 VSUBS 0.007334f
C526 B.n418 VSUBS 0.007334f
C527 B.n419 VSUBS 0.007334f
C528 B.n420 VSUBS 0.007334f
C529 B.n421 VSUBS 0.007334f
C530 B.n422 VSUBS 0.007334f
C531 B.n423 VSUBS 0.007334f
C532 B.n424 VSUBS 0.007334f
C533 B.n425 VSUBS 0.007334f
C534 B.n426 VSUBS 0.007334f
C535 B.n427 VSUBS 0.007334f
C536 B.n428 VSUBS 0.007334f
C537 B.n429 VSUBS 0.007334f
C538 B.n430 VSUBS 0.007334f
C539 B.n431 VSUBS 0.007334f
C540 B.n432 VSUBS 0.007334f
C541 B.n433 VSUBS 0.007334f
C542 B.n434 VSUBS 0.007334f
C543 B.n435 VSUBS 0.007334f
C544 B.n436 VSUBS 0.007334f
C545 B.n437 VSUBS 0.007334f
C546 B.n438 VSUBS 0.007334f
C547 B.n439 VSUBS 0.007334f
C548 B.n440 VSUBS 0.007334f
C549 B.n441 VSUBS 0.007334f
C550 B.n442 VSUBS 0.007334f
C551 B.n443 VSUBS 0.007334f
C552 B.n444 VSUBS 0.007334f
C553 B.n445 VSUBS 0.007334f
C554 B.n446 VSUBS 0.007334f
C555 B.n447 VSUBS 0.007334f
C556 B.n448 VSUBS 0.007334f
C557 B.n449 VSUBS 0.007334f
C558 B.n450 VSUBS 0.007334f
C559 B.n451 VSUBS 0.007334f
C560 B.n452 VSUBS 0.007334f
C561 B.n453 VSUBS 0.007334f
C562 B.n454 VSUBS 0.007334f
C563 B.n455 VSUBS 0.007334f
C564 B.n456 VSUBS 0.007334f
C565 B.n457 VSUBS 0.007334f
C566 B.n458 VSUBS 0.007334f
C567 B.n459 VSUBS 0.007334f
C568 B.n460 VSUBS 0.007334f
C569 B.n461 VSUBS 0.007334f
C570 B.n462 VSUBS 0.007334f
C571 B.n463 VSUBS 0.007334f
C572 B.n464 VSUBS 0.007334f
C573 B.n465 VSUBS 0.007334f
C574 B.n466 VSUBS 0.007334f
C575 B.n467 VSUBS 0.007334f
C576 B.n468 VSUBS 0.007334f
C577 B.n469 VSUBS 0.007334f
C578 B.n470 VSUBS 0.007334f
C579 B.n471 VSUBS 0.007334f
C580 B.n472 VSUBS 0.007334f
C581 B.n473 VSUBS 0.007334f
C582 B.n474 VSUBS 0.007334f
C583 B.n475 VSUBS 0.007334f
C584 B.n476 VSUBS 0.007334f
C585 B.n477 VSUBS 0.007334f
C586 B.n478 VSUBS 0.007334f
C587 B.n479 VSUBS 0.007334f
C588 B.n480 VSUBS 0.007334f
C589 B.n481 VSUBS 0.007334f
C590 B.n482 VSUBS 0.007334f
C591 B.n483 VSUBS 0.007334f
C592 B.n484 VSUBS 0.007334f
C593 B.n485 VSUBS 0.007334f
C594 B.n486 VSUBS 0.007334f
C595 B.n487 VSUBS 0.007334f
C596 B.n488 VSUBS 0.007334f
C597 B.n489 VSUBS 0.007334f
C598 B.n490 VSUBS 0.007334f
C599 B.n491 VSUBS 0.007334f
C600 B.n492 VSUBS 0.007334f
C601 B.n493 VSUBS 0.007334f
C602 B.n494 VSUBS 0.007334f
C603 B.n495 VSUBS 0.007334f
C604 B.n496 VSUBS 0.007334f
C605 B.n497 VSUBS 0.007334f
C606 B.n498 VSUBS 0.007334f
C607 B.n499 VSUBS 0.007334f
C608 B.n500 VSUBS 0.016496f
C609 B.n501 VSUBS 0.017586f
C610 B.n502 VSUBS 0.017586f
C611 B.n503 VSUBS 0.007334f
C612 B.n504 VSUBS 0.007334f
C613 B.n505 VSUBS 0.007334f
C614 B.n506 VSUBS 0.007334f
C615 B.n507 VSUBS 0.007334f
C616 B.n508 VSUBS 0.007334f
C617 B.n509 VSUBS 0.007334f
C618 B.n510 VSUBS 0.007334f
C619 B.n511 VSUBS 0.007334f
C620 B.n512 VSUBS 0.007334f
C621 B.n513 VSUBS 0.007334f
C622 B.n514 VSUBS 0.007334f
C623 B.n515 VSUBS 0.007334f
C624 B.n516 VSUBS 0.007334f
C625 B.n517 VSUBS 0.007334f
C626 B.n518 VSUBS 0.007334f
C627 B.n519 VSUBS 0.007334f
C628 B.n520 VSUBS 0.007334f
C629 B.n521 VSUBS 0.007334f
C630 B.n522 VSUBS 0.007334f
C631 B.n523 VSUBS 0.007334f
C632 B.n524 VSUBS 0.007334f
C633 B.n525 VSUBS 0.007334f
C634 B.n526 VSUBS 0.007334f
C635 B.n527 VSUBS 0.007334f
C636 B.n528 VSUBS 0.007334f
C637 B.n529 VSUBS 0.007334f
C638 B.n530 VSUBS 0.007334f
C639 B.n531 VSUBS 0.007334f
C640 B.n532 VSUBS 0.007334f
C641 B.n533 VSUBS 0.007334f
C642 B.n534 VSUBS 0.007334f
C643 B.n535 VSUBS 0.007334f
C644 B.n536 VSUBS 0.007334f
C645 B.n537 VSUBS 0.007334f
C646 B.n538 VSUBS 0.007334f
C647 B.n539 VSUBS 0.007334f
C648 B.n540 VSUBS 0.007334f
C649 B.n541 VSUBS 0.007334f
C650 B.n542 VSUBS 0.007334f
C651 B.n543 VSUBS 0.007334f
C652 B.n544 VSUBS 0.007334f
C653 B.n545 VSUBS 0.007334f
C654 B.n546 VSUBS 0.007334f
C655 B.n547 VSUBS 0.007334f
C656 B.n548 VSUBS 0.007334f
C657 B.n549 VSUBS 0.007334f
C658 B.n550 VSUBS 0.007334f
C659 B.n551 VSUBS 0.007334f
C660 B.n552 VSUBS 0.006903f
C661 B.n553 VSUBS 0.007334f
C662 B.n554 VSUBS 0.007334f
C663 B.n555 VSUBS 0.007334f
C664 B.n556 VSUBS 0.007334f
C665 B.n557 VSUBS 0.007334f
C666 B.n558 VSUBS 0.007334f
C667 B.n559 VSUBS 0.007334f
C668 B.n560 VSUBS 0.007334f
C669 B.n561 VSUBS 0.007334f
C670 B.n562 VSUBS 0.007334f
C671 B.n563 VSUBS 0.007334f
C672 B.n564 VSUBS 0.007334f
C673 B.n565 VSUBS 0.007334f
C674 B.n566 VSUBS 0.007334f
C675 B.n567 VSUBS 0.007334f
C676 B.n568 VSUBS 0.004098f
C677 B.n569 VSUBS 0.016992f
C678 B.n570 VSUBS 0.006903f
C679 B.n571 VSUBS 0.007334f
C680 B.n572 VSUBS 0.007334f
C681 B.n573 VSUBS 0.007334f
C682 B.n574 VSUBS 0.007334f
C683 B.n575 VSUBS 0.007334f
C684 B.n576 VSUBS 0.007334f
C685 B.n577 VSUBS 0.007334f
C686 B.n578 VSUBS 0.007334f
C687 B.n579 VSUBS 0.007334f
C688 B.n580 VSUBS 0.007334f
C689 B.n581 VSUBS 0.007334f
C690 B.n582 VSUBS 0.007334f
C691 B.n583 VSUBS 0.007334f
C692 B.n584 VSUBS 0.007334f
C693 B.n585 VSUBS 0.007334f
C694 B.n586 VSUBS 0.007334f
C695 B.n587 VSUBS 0.007334f
C696 B.n588 VSUBS 0.007334f
C697 B.n589 VSUBS 0.007334f
C698 B.n590 VSUBS 0.007334f
C699 B.n591 VSUBS 0.007334f
C700 B.n592 VSUBS 0.007334f
C701 B.n593 VSUBS 0.007334f
C702 B.n594 VSUBS 0.007334f
C703 B.n595 VSUBS 0.007334f
C704 B.n596 VSUBS 0.007334f
C705 B.n597 VSUBS 0.007334f
C706 B.n598 VSUBS 0.007334f
C707 B.n599 VSUBS 0.007334f
C708 B.n600 VSUBS 0.007334f
C709 B.n601 VSUBS 0.007334f
C710 B.n602 VSUBS 0.007334f
C711 B.n603 VSUBS 0.007334f
C712 B.n604 VSUBS 0.007334f
C713 B.n605 VSUBS 0.007334f
C714 B.n606 VSUBS 0.007334f
C715 B.n607 VSUBS 0.007334f
C716 B.n608 VSUBS 0.007334f
C717 B.n609 VSUBS 0.007334f
C718 B.n610 VSUBS 0.007334f
C719 B.n611 VSUBS 0.007334f
C720 B.n612 VSUBS 0.007334f
C721 B.n613 VSUBS 0.007334f
C722 B.n614 VSUBS 0.007334f
C723 B.n615 VSUBS 0.007334f
C724 B.n616 VSUBS 0.007334f
C725 B.n617 VSUBS 0.007334f
C726 B.n618 VSUBS 0.007334f
C727 B.n619 VSUBS 0.007334f
C728 B.n620 VSUBS 0.007334f
C729 B.n621 VSUBS 0.017586f
C730 B.n622 VSUBS 0.016496f
C731 B.n623 VSUBS 0.016496f
C732 B.n624 VSUBS 0.007334f
C733 B.n625 VSUBS 0.007334f
C734 B.n626 VSUBS 0.007334f
C735 B.n627 VSUBS 0.007334f
C736 B.n628 VSUBS 0.007334f
C737 B.n629 VSUBS 0.007334f
C738 B.n630 VSUBS 0.007334f
C739 B.n631 VSUBS 0.007334f
C740 B.n632 VSUBS 0.007334f
C741 B.n633 VSUBS 0.007334f
C742 B.n634 VSUBS 0.007334f
C743 B.n635 VSUBS 0.007334f
C744 B.n636 VSUBS 0.007334f
C745 B.n637 VSUBS 0.007334f
C746 B.n638 VSUBS 0.007334f
C747 B.n639 VSUBS 0.007334f
C748 B.n640 VSUBS 0.007334f
C749 B.n641 VSUBS 0.007334f
C750 B.n642 VSUBS 0.007334f
C751 B.n643 VSUBS 0.007334f
C752 B.n644 VSUBS 0.007334f
C753 B.n645 VSUBS 0.007334f
C754 B.n646 VSUBS 0.007334f
C755 B.n647 VSUBS 0.007334f
C756 B.n648 VSUBS 0.007334f
C757 B.n649 VSUBS 0.007334f
C758 B.n650 VSUBS 0.007334f
C759 B.n651 VSUBS 0.007334f
C760 B.n652 VSUBS 0.007334f
C761 B.n653 VSUBS 0.007334f
C762 B.n654 VSUBS 0.007334f
C763 B.n655 VSUBS 0.007334f
C764 B.n656 VSUBS 0.007334f
C765 B.n657 VSUBS 0.007334f
C766 B.n658 VSUBS 0.007334f
C767 B.n659 VSUBS 0.007334f
C768 B.n660 VSUBS 0.007334f
C769 B.n661 VSUBS 0.007334f
C770 B.n662 VSUBS 0.007334f
C771 B.n663 VSUBS 0.007334f
C772 B.n664 VSUBS 0.007334f
C773 B.n665 VSUBS 0.007334f
C774 B.n666 VSUBS 0.007334f
C775 B.n667 VSUBS 0.007334f
C776 B.n668 VSUBS 0.007334f
C777 B.n669 VSUBS 0.007334f
C778 B.n670 VSUBS 0.007334f
C779 B.n671 VSUBS 0.007334f
C780 B.n672 VSUBS 0.007334f
C781 B.n673 VSUBS 0.007334f
C782 B.n674 VSUBS 0.007334f
C783 B.n675 VSUBS 0.007334f
C784 B.n676 VSUBS 0.007334f
C785 B.n677 VSUBS 0.007334f
C786 B.n678 VSUBS 0.007334f
C787 B.n679 VSUBS 0.007334f
C788 B.n680 VSUBS 0.007334f
C789 B.n681 VSUBS 0.007334f
C790 B.n682 VSUBS 0.007334f
C791 B.n683 VSUBS 0.007334f
C792 B.n684 VSUBS 0.007334f
C793 B.n685 VSUBS 0.007334f
C794 B.n686 VSUBS 0.007334f
C795 B.n687 VSUBS 0.009571f
C796 B.n688 VSUBS 0.010195f
C797 B.n689 VSUBS 0.020274f
C798 VDD1.t5 VSUBS 0.190856f
C799 VDD1.t6 VSUBS 0.190856f
C800 VDD1.n0 VSUBS 1.45449f
C801 VDD1.t1 VSUBS 0.190856f
C802 VDD1.t7 VSUBS 0.190856f
C803 VDD1.n1 VSUBS 1.45343f
C804 VDD1.t3 VSUBS 0.190856f
C805 VDD1.t4 VSUBS 0.190856f
C806 VDD1.n2 VSUBS 1.45343f
C807 VDD1.n3 VSUBS 3.35314f
C808 VDD1.t0 VSUBS 0.190856f
C809 VDD1.t2 VSUBS 0.190856f
C810 VDD1.n4 VSUBS 1.44489f
C811 VDD1.n5 VSUBS 2.85002f
C812 VTAIL.t4 VSUBS 0.197828f
C813 VTAIL.t5 VSUBS 0.197828f
C814 VTAIL.n0 VSUBS 1.38321f
C815 VTAIL.n1 VSUBS 0.710415f
C816 VTAIL.t2 VSUBS 1.8387f
C817 VTAIL.n2 VSUBS 0.828378f
C818 VTAIL.t15 VSUBS 1.8387f
C819 VTAIL.n3 VSUBS 0.828378f
C820 VTAIL.t8 VSUBS 0.197828f
C821 VTAIL.t10 VSUBS 0.197828f
C822 VTAIL.n4 VSUBS 1.38321f
C823 VTAIL.n5 VSUBS 0.881778f
C824 VTAIL.t12 VSUBS 1.8387f
C825 VTAIL.n6 VSUBS 2.00858f
C826 VTAIL.t3 VSUBS 1.83871f
C827 VTAIL.n7 VSUBS 2.00856f
C828 VTAIL.t7 VSUBS 0.197828f
C829 VTAIL.t6 VSUBS 0.197828f
C830 VTAIL.n8 VSUBS 1.38322f
C831 VTAIL.n9 VSUBS 0.881773f
C832 VTAIL.t0 VSUBS 1.83871f
C833 VTAIL.n10 VSUBS 0.828366f
C834 VTAIL.t14 VSUBS 1.83871f
C835 VTAIL.n11 VSUBS 0.828366f
C836 VTAIL.t13 VSUBS 0.197828f
C837 VTAIL.t9 VSUBS 0.197828f
C838 VTAIL.n12 VSUBS 1.38322f
C839 VTAIL.n13 VSUBS 0.881773f
C840 VTAIL.t11 VSUBS 1.8387f
C841 VTAIL.n14 VSUBS 2.00857f
C842 VTAIL.t1 VSUBS 1.8387f
C843 VTAIL.n15 VSUBS 2.00378f
C844 VP.n0 VSUBS 0.045986f
C845 VP.t3 VSUBS 1.98745f
C846 VP.n1 VSUBS 0.048975f
C847 VP.n2 VSUBS 0.03488f
C848 VP.t4 VSUBS 1.98745f
C849 VP.n3 VSUBS 0.050919f
C850 VP.n4 VSUBS 0.03488f
C851 VP.t0 VSUBS 1.98745f
C852 VP.n5 VSUBS 0.065008f
C853 VP.n6 VSUBS 0.03488f
C854 VP.t6 VSUBS 1.98745f
C855 VP.n7 VSUBS 0.840021f
C856 VP.n8 VSUBS 0.045986f
C857 VP.t5 VSUBS 1.98745f
C858 VP.n9 VSUBS 0.048975f
C859 VP.n10 VSUBS 0.03488f
C860 VP.t7 VSUBS 1.98745f
C861 VP.n11 VSUBS 0.050919f
C862 VP.n12 VSUBS 0.294525f
C863 VP.t1 VSUBS 1.98745f
C864 VP.t2 VSUBS 2.20651f
C865 VP.n13 VSUBS 0.791671f
C866 VP.n14 VSUBS 0.823533f
C867 VP.n15 VSUBS 0.064366f
C868 VP.n16 VSUBS 0.050919f
C869 VP.n17 VSUBS 0.03488f
C870 VP.n18 VSUBS 0.03488f
C871 VP.n19 VSUBS 0.03488f
C872 VP.n20 VSUBS 0.064366f
C873 VP.n21 VSUBS 0.71793f
C874 VP.n22 VSUBS 0.033555f
C875 VP.n23 VSUBS 0.065008f
C876 VP.n24 VSUBS 0.03488f
C877 VP.n25 VSUBS 0.03488f
C878 VP.n26 VSUBS 0.03488f
C879 VP.n27 VSUBS 0.052863f
C880 VP.n28 VSUBS 0.063082f
C881 VP.n29 VSUBS 0.840021f
C882 VP.n30 VSUBS 1.76599f
C883 VP.n31 VSUBS 1.79254f
C884 VP.n32 VSUBS 0.045986f
C885 VP.n33 VSUBS 0.063082f
C886 VP.n34 VSUBS 0.052863f
C887 VP.n35 VSUBS 0.048975f
C888 VP.n36 VSUBS 0.03488f
C889 VP.n37 VSUBS 0.03488f
C890 VP.n38 VSUBS 0.03488f
C891 VP.n39 VSUBS 0.033555f
C892 VP.n40 VSUBS 0.71793f
C893 VP.n41 VSUBS 0.064366f
C894 VP.n42 VSUBS 0.050919f
C895 VP.n43 VSUBS 0.03488f
C896 VP.n44 VSUBS 0.03488f
C897 VP.n45 VSUBS 0.03488f
C898 VP.n46 VSUBS 0.064366f
C899 VP.n47 VSUBS 0.71793f
C900 VP.n48 VSUBS 0.033555f
C901 VP.n49 VSUBS 0.065008f
C902 VP.n50 VSUBS 0.03488f
C903 VP.n51 VSUBS 0.03488f
C904 VP.n52 VSUBS 0.03488f
C905 VP.n53 VSUBS 0.052863f
C906 VP.n54 VSUBS 0.063082f
C907 VP.n55 VSUBS 0.840021f
C908 VP.n56 VSUBS 0.039419f
.ends

