* NGSPICE file created from diff_pair_sample_0431.ext - technology: sky130A

.subckt diff_pair_sample_0431 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X1 VDD2.t9 VN.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=1.38
X2 VDD1.t2 VP.t1 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X3 VTAIL.t4 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=1.38
X5 VDD1.t7 VP.t2 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=1.38
X6 VTAIL.t3 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=1.38
X8 VDD1.t6 VP.t3 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=1.38
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=1.38
X10 VDD2.t6 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=1.38
X11 VDD1.t5 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=1.38
X12 VDD1.t4 VP.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=1.38
X13 VDD1.t9 VP.t6 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X14 VTAIL.t6 VN.t4 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X15 VTAIL.t12 VP.t7 VDD1.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X16 VDD2.t4 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=1.38
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=1.38
X18 VDD2.t3 VN.t6 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X19 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X20 VTAIL.t11 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X21 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X22 VTAIL.t10 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=1.38
X23 VDD2.t0 VN.t9 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=1.38
R0 VP.n14 VP.t5 326.76
R1 VP.n34 VP.t2 293.916
R2 VP.n5 VP.t0 293.916
R3 VP.n45 VP.t1 293.916
R4 VP.n52 VP.t7 293.916
R5 VP.n59 VP.t4 293.916
R6 VP.n32 VP.t3 293.916
R7 VP.n25 VP.t9 293.916
R8 VP.n18 VP.t6 293.916
R9 VP.n13 VP.t8 293.916
R10 VP.n35 VP.n34 177.448
R11 VP.n60 VP.n59 177.448
R12 VP.n33 VP.n32 177.448
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n12 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n11 161.3
R17 VP.n23 VP.n22 161.3
R18 VP.n24 VP.n10 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n28 VP.n9 161.3
R21 VP.n30 VP.n29 161.3
R22 VP.n31 VP.n8 161.3
R23 VP.n58 VP.n0 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n1 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n51 VP.n2 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n3 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n44 VP.n4 161.3
R32 VP.n43 VP.n42 161.3
R33 VP.n41 VP.n40 161.3
R34 VP.n39 VP.n6 161.3
R35 VP.n38 VP.n37 161.3
R36 VP.n36 VP.n7 161.3
R37 VP.n39 VP.n38 56.5193
R38 VP.n57 VP.n1 56.5193
R39 VP.n30 VP.n9 56.5193
R40 VP.n44 VP.n43 50.6917
R41 VP.n51 VP.n50 50.6917
R42 VP.n24 VP.n23 50.6917
R43 VP.n17 VP.n16 50.6917
R44 VP.n35 VP.n33 50.0119
R45 VP.n14 VP.n13 43.6963
R46 VP.n46 VP.n44 30.2951
R47 VP.n50 VP.n3 30.2951
R48 VP.n23 VP.n11 30.2951
R49 VP.n19 VP.n17 30.2951
R50 VP.n38 VP.n7 24.4675
R51 VP.n40 VP.n39 24.4675
R52 VP.n53 VP.n1 24.4675
R53 VP.n58 VP.n57 24.4675
R54 VP.n31 VP.n30 24.4675
R55 VP.n26 VP.n9 24.4675
R56 VP.n43 VP.n5 22.5101
R57 VP.n52 VP.n51 22.5101
R58 VP.n25 VP.n24 22.5101
R59 VP.n16 VP.n13 22.5101
R60 VP.n15 VP.n14 17.9509
R61 VP.n46 VP.n45 12.234
R62 VP.n45 VP.n3 12.234
R63 VP.n19 VP.n18 12.234
R64 VP.n18 VP.n11 12.234
R65 VP.n34 VP.n7 8.31928
R66 VP.n59 VP.n58 8.31928
R67 VP.n32 VP.n31 8.31928
R68 VP.n40 VP.n5 1.95786
R69 VP.n53 VP.n52 1.95786
R70 VP.n26 VP.n25 1.95786
R71 VP.n15 VP.n12 0.189894
R72 VP.n20 VP.n12 0.189894
R73 VP.n21 VP.n20 0.189894
R74 VP.n22 VP.n21 0.189894
R75 VP.n22 VP.n10 0.189894
R76 VP.n27 VP.n10 0.189894
R77 VP.n28 VP.n27 0.189894
R78 VP.n29 VP.n28 0.189894
R79 VP.n29 VP.n8 0.189894
R80 VP.n33 VP.n8 0.189894
R81 VP.n36 VP.n35 0.189894
R82 VP.n37 VP.n36 0.189894
R83 VP.n37 VP.n6 0.189894
R84 VP.n41 VP.n6 0.189894
R85 VP.n42 VP.n41 0.189894
R86 VP.n42 VP.n4 0.189894
R87 VP.n47 VP.n4 0.189894
R88 VP.n48 VP.n47 0.189894
R89 VP.n49 VP.n48 0.189894
R90 VP.n49 VP.n2 0.189894
R91 VP.n54 VP.n2 0.189894
R92 VP.n55 VP.n54 0.189894
R93 VP.n56 VP.n55 0.189894
R94 VP.n56 VP.n0 0.189894
R95 VP.n60 VP.n0 0.189894
R96 VP VP.n60 0.0516364
R97 VDD1.n88 VDD1.n0 289.615
R98 VDD1.n183 VDD1.n95 289.615
R99 VDD1.n89 VDD1.n88 185
R100 VDD1.n87 VDD1.n86 185
R101 VDD1.n4 VDD1.n3 185
R102 VDD1.n81 VDD1.n80 185
R103 VDD1.n79 VDD1.n78 185
R104 VDD1.n77 VDD1.n7 185
R105 VDD1.n11 VDD1.n8 185
R106 VDD1.n72 VDD1.n71 185
R107 VDD1.n70 VDD1.n69 185
R108 VDD1.n13 VDD1.n12 185
R109 VDD1.n64 VDD1.n63 185
R110 VDD1.n62 VDD1.n61 185
R111 VDD1.n17 VDD1.n16 185
R112 VDD1.n56 VDD1.n55 185
R113 VDD1.n54 VDD1.n53 185
R114 VDD1.n21 VDD1.n20 185
R115 VDD1.n48 VDD1.n47 185
R116 VDD1.n46 VDD1.n45 185
R117 VDD1.n25 VDD1.n24 185
R118 VDD1.n40 VDD1.n39 185
R119 VDD1.n38 VDD1.n37 185
R120 VDD1.n29 VDD1.n28 185
R121 VDD1.n32 VDD1.n31 185
R122 VDD1.n126 VDD1.n125 185
R123 VDD1.n123 VDD1.n122 185
R124 VDD1.n132 VDD1.n131 185
R125 VDD1.n134 VDD1.n133 185
R126 VDD1.n119 VDD1.n118 185
R127 VDD1.n140 VDD1.n139 185
R128 VDD1.n142 VDD1.n141 185
R129 VDD1.n115 VDD1.n114 185
R130 VDD1.n148 VDD1.n147 185
R131 VDD1.n150 VDD1.n149 185
R132 VDD1.n111 VDD1.n110 185
R133 VDD1.n156 VDD1.n155 185
R134 VDD1.n158 VDD1.n157 185
R135 VDD1.n107 VDD1.n106 185
R136 VDD1.n164 VDD1.n163 185
R137 VDD1.n167 VDD1.n166 185
R138 VDD1.n165 VDD1.n103 185
R139 VDD1.n172 VDD1.n102 185
R140 VDD1.n174 VDD1.n173 185
R141 VDD1.n176 VDD1.n175 185
R142 VDD1.n99 VDD1.n98 185
R143 VDD1.n182 VDD1.n181 185
R144 VDD1.n184 VDD1.n183 185
R145 VDD1.t4 VDD1.n30 147.659
R146 VDD1.t7 VDD1.n124 147.659
R147 VDD1.n88 VDD1.n87 104.615
R148 VDD1.n87 VDD1.n3 104.615
R149 VDD1.n80 VDD1.n3 104.615
R150 VDD1.n80 VDD1.n79 104.615
R151 VDD1.n79 VDD1.n7 104.615
R152 VDD1.n11 VDD1.n7 104.615
R153 VDD1.n71 VDD1.n11 104.615
R154 VDD1.n71 VDD1.n70 104.615
R155 VDD1.n70 VDD1.n12 104.615
R156 VDD1.n63 VDD1.n12 104.615
R157 VDD1.n63 VDD1.n62 104.615
R158 VDD1.n62 VDD1.n16 104.615
R159 VDD1.n55 VDD1.n16 104.615
R160 VDD1.n55 VDD1.n54 104.615
R161 VDD1.n54 VDD1.n20 104.615
R162 VDD1.n47 VDD1.n20 104.615
R163 VDD1.n47 VDD1.n46 104.615
R164 VDD1.n46 VDD1.n24 104.615
R165 VDD1.n39 VDD1.n24 104.615
R166 VDD1.n39 VDD1.n38 104.615
R167 VDD1.n38 VDD1.n28 104.615
R168 VDD1.n31 VDD1.n28 104.615
R169 VDD1.n125 VDD1.n122 104.615
R170 VDD1.n132 VDD1.n122 104.615
R171 VDD1.n133 VDD1.n132 104.615
R172 VDD1.n133 VDD1.n118 104.615
R173 VDD1.n140 VDD1.n118 104.615
R174 VDD1.n141 VDD1.n140 104.615
R175 VDD1.n141 VDD1.n114 104.615
R176 VDD1.n148 VDD1.n114 104.615
R177 VDD1.n149 VDD1.n148 104.615
R178 VDD1.n149 VDD1.n110 104.615
R179 VDD1.n156 VDD1.n110 104.615
R180 VDD1.n157 VDD1.n156 104.615
R181 VDD1.n157 VDD1.n106 104.615
R182 VDD1.n164 VDD1.n106 104.615
R183 VDD1.n166 VDD1.n164 104.615
R184 VDD1.n166 VDD1.n165 104.615
R185 VDD1.n165 VDD1.n102 104.615
R186 VDD1.n174 VDD1.n102 104.615
R187 VDD1.n175 VDD1.n174 104.615
R188 VDD1.n175 VDD1.n98 104.615
R189 VDD1.n182 VDD1.n98 104.615
R190 VDD1.n183 VDD1.n182 104.615
R191 VDD1.n191 VDD1.n190 62.3567
R192 VDD1.n94 VDD1.n93 61.3066
R193 VDD1.n193 VDD1.n192 61.3065
R194 VDD1.n189 VDD1.n188 61.3065
R195 VDD1.n31 VDD1.t4 52.3082
R196 VDD1.n125 VDD1.t7 52.3082
R197 VDD1.n94 VDD1.n92 50.9201
R198 VDD1.n189 VDD1.n187 50.9201
R199 VDD1.n193 VDD1.n191 46.5462
R200 VDD1.n32 VDD1.n30 15.6677
R201 VDD1.n126 VDD1.n124 15.6677
R202 VDD1.n78 VDD1.n77 13.1884
R203 VDD1.n173 VDD1.n172 13.1884
R204 VDD1.n81 VDD1.n6 12.8005
R205 VDD1.n76 VDD1.n8 12.8005
R206 VDD1.n33 VDD1.n29 12.8005
R207 VDD1.n127 VDD1.n123 12.8005
R208 VDD1.n171 VDD1.n103 12.8005
R209 VDD1.n176 VDD1.n101 12.8005
R210 VDD1.n82 VDD1.n4 12.0247
R211 VDD1.n73 VDD1.n72 12.0247
R212 VDD1.n37 VDD1.n36 12.0247
R213 VDD1.n131 VDD1.n130 12.0247
R214 VDD1.n168 VDD1.n167 12.0247
R215 VDD1.n177 VDD1.n99 12.0247
R216 VDD1.n86 VDD1.n85 11.249
R217 VDD1.n69 VDD1.n10 11.249
R218 VDD1.n40 VDD1.n27 11.249
R219 VDD1.n134 VDD1.n121 11.249
R220 VDD1.n163 VDD1.n105 11.249
R221 VDD1.n181 VDD1.n180 11.249
R222 VDD1.n89 VDD1.n2 10.4732
R223 VDD1.n68 VDD1.n13 10.4732
R224 VDD1.n41 VDD1.n25 10.4732
R225 VDD1.n135 VDD1.n119 10.4732
R226 VDD1.n162 VDD1.n107 10.4732
R227 VDD1.n184 VDD1.n97 10.4732
R228 VDD1.n90 VDD1.n0 9.69747
R229 VDD1.n65 VDD1.n64 9.69747
R230 VDD1.n45 VDD1.n44 9.69747
R231 VDD1.n139 VDD1.n138 9.69747
R232 VDD1.n159 VDD1.n158 9.69747
R233 VDD1.n185 VDD1.n95 9.69747
R234 VDD1.n92 VDD1.n91 9.45567
R235 VDD1.n187 VDD1.n186 9.45567
R236 VDD1.n58 VDD1.n57 9.3005
R237 VDD1.n60 VDD1.n59 9.3005
R238 VDD1.n15 VDD1.n14 9.3005
R239 VDD1.n66 VDD1.n65 9.3005
R240 VDD1.n68 VDD1.n67 9.3005
R241 VDD1.n10 VDD1.n9 9.3005
R242 VDD1.n74 VDD1.n73 9.3005
R243 VDD1.n76 VDD1.n75 9.3005
R244 VDD1.n91 VDD1.n90 9.3005
R245 VDD1.n2 VDD1.n1 9.3005
R246 VDD1.n85 VDD1.n84 9.3005
R247 VDD1.n83 VDD1.n82 9.3005
R248 VDD1.n6 VDD1.n5 9.3005
R249 VDD1.n19 VDD1.n18 9.3005
R250 VDD1.n52 VDD1.n51 9.3005
R251 VDD1.n50 VDD1.n49 9.3005
R252 VDD1.n23 VDD1.n22 9.3005
R253 VDD1.n44 VDD1.n43 9.3005
R254 VDD1.n42 VDD1.n41 9.3005
R255 VDD1.n27 VDD1.n26 9.3005
R256 VDD1.n36 VDD1.n35 9.3005
R257 VDD1.n34 VDD1.n33 9.3005
R258 VDD1.n186 VDD1.n185 9.3005
R259 VDD1.n97 VDD1.n96 9.3005
R260 VDD1.n180 VDD1.n179 9.3005
R261 VDD1.n178 VDD1.n177 9.3005
R262 VDD1.n101 VDD1.n100 9.3005
R263 VDD1.n146 VDD1.n145 9.3005
R264 VDD1.n144 VDD1.n143 9.3005
R265 VDD1.n117 VDD1.n116 9.3005
R266 VDD1.n138 VDD1.n137 9.3005
R267 VDD1.n136 VDD1.n135 9.3005
R268 VDD1.n121 VDD1.n120 9.3005
R269 VDD1.n130 VDD1.n129 9.3005
R270 VDD1.n128 VDD1.n127 9.3005
R271 VDD1.n113 VDD1.n112 9.3005
R272 VDD1.n152 VDD1.n151 9.3005
R273 VDD1.n154 VDD1.n153 9.3005
R274 VDD1.n109 VDD1.n108 9.3005
R275 VDD1.n160 VDD1.n159 9.3005
R276 VDD1.n162 VDD1.n161 9.3005
R277 VDD1.n105 VDD1.n104 9.3005
R278 VDD1.n169 VDD1.n168 9.3005
R279 VDD1.n171 VDD1.n170 9.3005
R280 VDD1.n61 VDD1.n15 8.92171
R281 VDD1.n48 VDD1.n23 8.92171
R282 VDD1.n142 VDD1.n117 8.92171
R283 VDD1.n155 VDD1.n109 8.92171
R284 VDD1.n60 VDD1.n17 8.14595
R285 VDD1.n49 VDD1.n21 8.14595
R286 VDD1.n143 VDD1.n115 8.14595
R287 VDD1.n154 VDD1.n111 8.14595
R288 VDD1.n57 VDD1.n56 7.3702
R289 VDD1.n53 VDD1.n52 7.3702
R290 VDD1.n147 VDD1.n146 7.3702
R291 VDD1.n151 VDD1.n150 7.3702
R292 VDD1.n56 VDD1.n19 6.59444
R293 VDD1.n53 VDD1.n19 6.59444
R294 VDD1.n147 VDD1.n113 6.59444
R295 VDD1.n150 VDD1.n113 6.59444
R296 VDD1.n57 VDD1.n17 5.81868
R297 VDD1.n52 VDD1.n21 5.81868
R298 VDD1.n146 VDD1.n115 5.81868
R299 VDD1.n151 VDD1.n111 5.81868
R300 VDD1.n61 VDD1.n60 5.04292
R301 VDD1.n49 VDD1.n48 5.04292
R302 VDD1.n143 VDD1.n142 5.04292
R303 VDD1.n155 VDD1.n154 5.04292
R304 VDD1.n34 VDD1.n30 4.38563
R305 VDD1.n128 VDD1.n124 4.38563
R306 VDD1.n92 VDD1.n0 4.26717
R307 VDD1.n64 VDD1.n15 4.26717
R308 VDD1.n45 VDD1.n23 4.26717
R309 VDD1.n139 VDD1.n117 4.26717
R310 VDD1.n158 VDD1.n109 4.26717
R311 VDD1.n187 VDD1.n95 4.26717
R312 VDD1.n90 VDD1.n89 3.49141
R313 VDD1.n65 VDD1.n13 3.49141
R314 VDD1.n44 VDD1.n25 3.49141
R315 VDD1.n138 VDD1.n119 3.49141
R316 VDD1.n159 VDD1.n107 3.49141
R317 VDD1.n185 VDD1.n184 3.49141
R318 VDD1.n86 VDD1.n2 2.71565
R319 VDD1.n69 VDD1.n68 2.71565
R320 VDD1.n41 VDD1.n40 2.71565
R321 VDD1.n135 VDD1.n134 2.71565
R322 VDD1.n163 VDD1.n162 2.71565
R323 VDD1.n181 VDD1.n97 2.71565
R324 VDD1.n85 VDD1.n4 1.93989
R325 VDD1.n72 VDD1.n10 1.93989
R326 VDD1.n37 VDD1.n27 1.93989
R327 VDD1.n131 VDD1.n121 1.93989
R328 VDD1.n167 VDD1.n105 1.93989
R329 VDD1.n180 VDD1.n99 1.93989
R330 VDD1.n192 VDD1.t0 1.17697
R331 VDD1.n192 VDD1.t6 1.17697
R332 VDD1.n93 VDD1.t1 1.17697
R333 VDD1.n93 VDD1.t9 1.17697
R334 VDD1.n190 VDD1.t8 1.17697
R335 VDD1.n190 VDD1.t5 1.17697
R336 VDD1.n188 VDD1.t3 1.17697
R337 VDD1.n188 VDD1.t2 1.17697
R338 VDD1.n82 VDD1.n81 1.16414
R339 VDD1.n73 VDD1.n8 1.16414
R340 VDD1.n36 VDD1.n29 1.16414
R341 VDD1.n130 VDD1.n123 1.16414
R342 VDD1.n168 VDD1.n103 1.16414
R343 VDD1.n177 VDD1.n176 1.16414
R344 VDD1 VDD1.n193 1.04791
R345 VDD1 VDD1.n94 0.427224
R346 VDD1.n78 VDD1.n6 0.388379
R347 VDD1.n77 VDD1.n76 0.388379
R348 VDD1.n33 VDD1.n32 0.388379
R349 VDD1.n127 VDD1.n126 0.388379
R350 VDD1.n172 VDD1.n171 0.388379
R351 VDD1.n173 VDD1.n101 0.388379
R352 VDD1.n191 VDD1.n189 0.313688
R353 VDD1.n91 VDD1.n1 0.155672
R354 VDD1.n84 VDD1.n1 0.155672
R355 VDD1.n84 VDD1.n83 0.155672
R356 VDD1.n83 VDD1.n5 0.155672
R357 VDD1.n75 VDD1.n5 0.155672
R358 VDD1.n75 VDD1.n74 0.155672
R359 VDD1.n74 VDD1.n9 0.155672
R360 VDD1.n67 VDD1.n9 0.155672
R361 VDD1.n67 VDD1.n66 0.155672
R362 VDD1.n66 VDD1.n14 0.155672
R363 VDD1.n59 VDD1.n14 0.155672
R364 VDD1.n59 VDD1.n58 0.155672
R365 VDD1.n58 VDD1.n18 0.155672
R366 VDD1.n51 VDD1.n18 0.155672
R367 VDD1.n51 VDD1.n50 0.155672
R368 VDD1.n50 VDD1.n22 0.155672
R369 VDD1.n43 VDD1.n22 0.155672
R370 VDD1.n43 VDD1.n42 0.155672
R371 VDD1.n42 VDD1.n26 0.155672
R372 VDD1.n35 VDD1.n26 0.155672
R373 VDD1.n35 VDD1.n34 0.155672
R374 VDD1.n129 VDD1.n128 0.155672
R375 VDD1.n129 VDD1.n120 0.155672
R376 VDD1.n136 VDD1.n120 0.155672
R377 VDD1.n137 VDD1.n136 0.155672
R378 VDD1.n137 VDD1.n116 0.155672
R379 VDD1.n144 VDD1.n116 0.155672
R380 VDD1.n145 VDD1.n144 0.155672
R381 VDD1.n145 VDD1.n112 0.155672
R382 VDD1.n152 VDD1.n112 0.155672
R383 VDD1.n153 VDD1.n152 0.155672
R384 VDD1.n153 VDD1.n108 0.155672
R385 VDD1.n160 VDD1.n108 0.155672
R386 VDD1.n161 VDD1.n160 0.155672
R387 VDD1.n161 VDD1.n104 0.155672
R388 VDD1.n169 VDD1.n104 0.155672
R389 VDD1.n170 VDD1.n169 0.155672
R390 VDD1.n170 VDD1.n100 0.155672
R391 VDD1.n178 VDD1.n100 0.155672
R392 VDD1.n179 VDD1.n178 0.155672
R393 VDD1.n179 VDD1.n96 0.155672
R394 VDD1.n186 VDD1.n96 0.155672
R395 VTAIL.n384 VTAIL.n296 289.615
R396 VTAIL.n90 VTAIL.n2 289.615
R397 VTAIL.n290 VTAIL.n202 289.615
R398 VTAIL.n192 VTAIL.n104 289.615
R399 VTAIL.n327 VTAIL.n326 185
R400 VTAIL.n324 VTAIL.n323 185
R401 VTAIL.n333 VTAIL.n332 185
R402 VTAIL.n335 VTAIL.n334 185
R403 VTAIL.n320 VTAIL.n319 185
R404 VTAIL.n341 VTAIL.n340 185
R405 VTAIL.n343 VTAIL.n342 185
R406 VTAIL.n316 VTAIL.n315 185
R407 VTAIL.n349 VTAIL.n348 185
R408 VTAIL.n351 VTAIL.n350 185
R409 VTAIL.n312 VTAIL.n311 185
R410 VTAIL.n357 VTAIL.n356 185
R411 VTAIL.n359 VTAIL.n358 185
R412 VTAIL.n308 VTAIL.n307 185
R413 VTAIL.n365 VTAIL.n364 185
R414 VTAIL.n368 VTAIL.n367 185
R415 VTAIL.n366 VTAIL.n304 185
R416 VTAIL.n373 VTAIL.n303 185
R417 VTAIL.n375 VTAIL.n374 185
R418 VTAIL.n377 VTAIL.n376 185
R419 VTAIL.n300 VTAIL.n299 185
R420 VTAIL.n383 VTAIL.n382 185
R421 VTAIL.n385 VTAIL.n384 185
R422 VTAIL.n33 VTAIL.n32 185
R423 VTAIL.n30 VTAIL.n29 185
R424 VTAIL.n39 VTAIL.n38 185
R425 VTAIL.n41 VTAIL.n40 185
R426 VTAIL.n26 VTAIL.n25 185
R427 VTAIL.n47 VTAIL.n46 185
R428 VTAIL.n49 VTAIL.n48 185
R429 VTAIL.n22 VTAIL.n21 185
R430 VTAIL.n55 VTAIL.n54 185
R431 VTAIL.n57 VTAIL.n56 185
R432 VTAIL.n18 VTAIL.n17 185
R433 VTAIL.n63 VTAIL.n62 185
R434 VTAIL.n65 VTAIL.n64 185
R435 VTAIL.n14 VTAIL.n13 185
R436 VTAIL.n71 VTAIL.n70 185
R437 VTAIL.n74 VTAIL.n73 185
R438 VTAIL.n72 VTAIL.n10 185
R439 VTAIL.n79 VTAIL.n9 185
R440 VTAIL.n81 VTAIL.n80 185
R441 VTAIL.n83 VTAIL.n82 185
R442 VTAIL.n6 VTAIL.n5 185
R443 VTAIL.n89 VTAIL.n88 185
R444 VTAIL.n91 VTAIL.n90 185
R445 VTAIL.n291 VTAIL.n290 185
R446 VTAIL.n289 VTAIL.n288 185
R447 VTAIL.n206 VTAIL.n205 185
R448 VTAIL.n283 VTAIL.n282 185
R449 VTAIL.n281 VTAIL.n280 185
R450 VTAIL.n279 VTAIL.n209 185
R451 VTAIL.n213 VTAIL.n210 185
R452 VTAIL.n274 VTAIL.n273 185
R453 VTAIL.n272 VTAIL.n271 185
R454 VTAIL.n215 VTAIL.n214 185
R455 VTAIL.n266 VTAIL.n265 185
R456 VTAIL.n264 VTAIL.n263 185
R457 VTAIL.n219 VTAIL.n218 185
R458 VTAIL.n258 VTAIL.n257 185
R459 VTAIL.n256 VTAIL.n255 185
R460 VTAIL.n223 VTAIL.n222 185
R461 VTAIL.n250 VTAIL.n249 185
R462 VTAIL.n248 VTAIL.n247 185
R463 VTAIL.n227 VTAIL.n226 185
R464 VTAIL.n242 VTAIL.n241 185
R465 VTAIL.n240 VTAIL.n239 185
R466 VTAIL.n231 VTAIL.n230 185
R467 VTAIL.n234 VTAIL.n233 185
R468 VTAIL.n193 VTAIL.n192 185
R469 VTAIL.n191 VTAIL.n190 185
R470 VTAIL.n108 VTAIL.n107 185
R471 VTAIL.n185 VTAIL.n184 185
R472 VTAIL.n183 VTAIL.n182 185
R473 VTAIL.n181 VTAIL.n111 185
R474 VTAIL.n115 VTAIL.n112 185
R475 VTAIL.n176 VTAIL.n175 185
R476 VTAIL.n174 VTAIL.n173 185
R477 VTAIL.n117 VTAIL.n116 185
R478 VTAIL.n168 VTAIL.n167 185
R479 VTAIL.n166 VTAIL.n165 185
R480 VTAIL.n121 VTAIL.n120 185
R481 VTAIL.n160 VTAIL.n159 185
R482 VTAIL.n158 VTAIL.n157 185
R483 VTAIL.n125 VTAIL.n124 185
R484 VTAIL.n152 VTAIL.n151 185
R485 VTAIL.n150 VTAIL.n149 185
R486 VTAIL.n129 VTAIL.n128 185
R487 VTAIL.n144 VTAIL.n143 185
R488 VTAIL.n142 VTAIL.n141 185
R489 VTAIL.n133 VTAIL.n132 185
R490 VTAIL.n136 VTAIL.n135 185
R491 VTAIL.t16 VTAIL.n232 147.659
R492 VTAIL.t5 VTAIL.n134 147.659
R493 VTAIL.t9 VTAIL.n325 147.659
R494 VTAIL.t15 VTAIL.n31 147.659
R495 VTAIL.n326 VTAIL.n323 104.615
R496 VTAIL.n333 VTAIL.n323 104.615
R497 VTAIL.n334 VTAIL.n333 104.615
R498 VTAIL.n334 VTAIL.n319 104.615
R499 VTAIL.n341 VTAIL.n319 104.615
R500 VTAIL.n342 VTAIL.n341 104.615
R501 VTAIL.n342 VTAIL.n315 104.615
R502 VTAIL.n349 VTAIL.n315 104.615
R503 VTAIL.n350 VTAIL.n349 104.615
R504 VTAIL.n350 VTAIL.n311 104.615
R505 VTAIL.n357 VTAIL.n311 104.615
R506 VTAIL.n358 VTAIL.n357 104.615
R507 VTAIL.n358 VTAIL.n307 104.615
R508 VTAIL.n365 VTAIL.n307 104.615
R509 VTAIL.n367 VTAIL.n365 104.615
R510 VTAIL.n367 VTAIL.n366 104.615
R511 VTAIL.n366 VTAIL.n303 104.615
R512 VTAIL.n375 VTAIL.n303 104.615
R513 VTAIL.n376 VTAIL.n375 104.615
R514 VTAIL.n376 VTAIL.n299 104.615
R515 VTAIL.n383 VTAIL.n299 104.615
R516 VTAIL.n384 VTAIL.n383 104.615
R517 VTAIL.n32 VTAIL.n29 104.615
R518 VTAIL.n39 VTAIL.n29 104.615
R519 VTAIL.n40 VTAIL.n39 104.615
R520 VTAIL.n40 VTAIL.n25 104.615
R521 VTAIL.n47 VTAIL.n25 104.615
R522 VTAIL.n48 VTAIL.n47 104.615
R523 VTAIL.n48 VTAIL.n21 104.615
R524 VTAIL.n55 VTAIL.n21 104.615
R525 VTAIL.n56 VTAIL.n55 104.615
R526 VTAIL.n56 VTAIL.n17 104.615
R527 VTAIL.n63 VTAIL.n17 104.615
R528 VTAIL.n64 VTAIL.n63 104.615
R529 VTAIL.n64 VTAIL.n13 104.615
R530 VTAIL.n71 VTAIL.n13 104.615
R531 VTAIL.n73 VTAIL.n71 104.615
R532 VTAIL.n73 VTAIL.n72 104.615
R533 VTAIL.n72 VTAIL.n9 104.615
R534 VTAIL.n81 VTAIL.n9 104.615
R535 VTAIL.n82 VTAIL.n81 104.615
R536 VTAIL.n82 VTAIL.n5 104.615
R537 VTAIL.n89 VTAIL.n5 104.615
R538 VTAIL.n90 VTAIL.n89 104.615
R539 VTAIL.n290 VTAIL.n289 104.615
R540 VTAIL.n289 VTAIL.n205 104.615
R541 VTAIL.n282 VTAIL.n205 104.615
R542 VTAIL.n282 VTAIL.n281 104.615
R543 VTAIL.n281 VTAIL.n209 104.615
R544 VTAIL.n213 VTAIL.n209 104.615
R545 VTAIL.n273 VTAIL.n213 104.615
R546 VTAIL.n273 VTAIL.n272 104.615
R547 VTAIL.n272 VTAIL.n214 104.615
R548 VTAIL.n265 VTAIL.n214 104.615
R549 VTAIL.n265 VTAIL.n264 104.615
R550 VTAIL.n264 VTAIL.n218 104.615
R551 VTAIL.n257 VTAIL.n218 104.615
R552 VTAIL.n257 VTAIL.n256 104.615
R553 VTAIL.n256 VTAIL.n222 104.615
R554 VTAIL.n249 VTAIL.n222 104.615
R555 VTAIL.n249 VTAIL.n248 104.615
R556 VTAIL.n248 VTAIL.n226 104.615
R557 VTAIL.n241 VTAIL.n226 104.615
R558 VTAIL.n241 VTAIL.n240 104.615
R559 VTAIL.n240 VTAIL.n230 104.615
R560 VTAIL.n233 VTAIL.n230 104.615
R561 VTAIL.n192 VTAIL.n191 104.615
R562 VTAIL.n191 VTAIL.n107 104.615
R563 VTAIL.n184 VTAIL.n107 104.615
R564 VTAIL.n184 VTAIL.n183 104.615
R565 VTAIL.n183 VTAIL.n111 104.615
R566 VTAIL.n115 VTAIL.n111 104.615
R567 VTAIL.n175 VTAIL.n115 104.615
R568 VTAIL.n175 VTAIL.n174 104.615
R569 VTAIL.n174 VTAIL.n116 104.615
R570 VTAIL.n167 VTAIL.n116 104.615
R571 VTAIL.n167 VTAIL.n166 104.615
R572 VTAIL.n166 VTAIL.n120 104.615
R573 VTAIL.n159 VTAIL.n120 104.615
R574 VTAIL.n159 VTAIL.n158 104.615
R575 VTAIL.n158 VTAIL.n124 104.615
R576 VTAIL.n151 VTAIL.n124 104.615
R577 VTAIL.n151 VTAIL.n150 104.615
R578 VTAIL.n150 VTAIL.n128 104.615
R579 VTAIL.n143 VTAIL.n128 104.615
R580 VTAIL.n143 VTAIL.n142 104.615
R581 VTAIL.n142 VTAIL.n132 104.615
R582 VTAIL.n135 VTAIL.n132 104.615
R583 VTAIL.n326 VTAIL.t9 52.3082
R584 VTAIL.n32 VTAIL.t15 52.3082
R585 VTAIL.n233 VTAIL.t16 52.3082
R586 VTAIL.n135 VTAIL.t5 52.3082
R587 VTAIL.n201 VTAIL.n200 44.6278
R588 VTAIL.n199 VTAIL.n198 44.6278
R589 VTAIL.n103 VTAIL.n102 44.6278
R590 VTAIL.n101 VTAIL.n100 44.6278
R591 VTAIL.n391 VTAIL.n390 44.6277
R592 VTAIL.n1 VTAIL.n0 44.6277
R593 VTAIL.n97 VTAIL.n96 44.6277
R594 VTAIL.n99 VTAIL.n98 44.6277
R595 VTAIL.n389 VTAIL.n388 32.7672
R596 VTAIL.n95 VTAIL.n94 32.7672
R597 VTAIL.n295 VTAIL.n294 32.7672
R598 VTAIL.n197 VTAIL.n196 32.7672
R599 VTAIL.n101 VTAIL.n99 29.8238
R600 VTAIL.n389 VTAIL.n295 28.3496
R601 VTAIL.n327 VTAIL.n325 15.6677
R602 VTAIL.n33 VTAIL.n31 15.6677
R603 VTAIL.n234 VTAIL.n232 15.6677
R604 VTAIL.n136 VTAIL.n134 15.6677
R605 VTAIL.n374 VTAIL.n373 13.1884
R606 VTAIL.n80 VTAIL.n79 13.1884
R607 VTAIL.n280 VTAIL.n279 13.1884
R608 VTAIL.n182 VTAIL.n181 13.1884
R609 VTAIL.n328 VTAIL.n324 12.8005
R610 VTAIL.n372 VTAIL.n304 12.8005
R611 VTAIL.n377 VTAIL.n302 12.8005
R612 VTAIL.n34 VTAIL.n30 12.8005
R613 VTAIL.n78 VTAIL.n10 12.8005
R614 VTAIL.n83 VTAIL.n8 12.8005
R615 VTAIL.n283 VTAIL.n208 12.8005
R616 VTAIL.n278 VTAIL.n210 12.8005
R617 VTAIL.n235 VTAIL.n231 12.8005
R618 VTAIL.n185 VTAIL.n110 12.8005
R619 VTAIL.n180 VTAIL.n112 12.8005
R620 VTAIL.n137 VTAIL.n133 12.8005
R621 VTAIL.n332 VTAIL.n331 12.0247
R622 VTAIL.n369 VTAIL.n368 12.0247
R623 VTAIL.n378 VTAIL.n300 12.0247
R624 VTAIL.n38 VTAIL.n37 12.0247
R625 VTAIL.n75 VTAIL.n74 12.0247
R626 VTAIL.n84 VTAIL.n6 12.0247
R627 VTAIL.n284 VTAIL.n206 12.0247
R628 VTAIL.n275 VTAIL.n274 12.0247
R629 VTAIL.n239 VTAIL.n238 12.0247
R630 VTAIL.n186 VTAIL.n108 12.0247
R631 VTAIL.n177 VTAIL.n176 12.0247
R632 VTAIL.n141 VTAIL.n140 12.0247
R633 VTAIL.n335 VTAIL.n322 11.249
R634 VTAIL.n364 VTAIL.n306 11.249
R635 VTAIL.n382 VTAIL.n381 11.249
R636 VTAIL.n41 VTAIL.n28 11.249
R637 VTAIL.n70 VTAIL.n12 11.249
R638 VTAIL.n88 VTAIL.n87 11.249
R639 VTAIL.n288 VTAIL.n287 11.249
R640 VTAIL.n271 VTAIL.n212 11.249
R641 VTAIL.n242 VTAIL.n229 11.249
R642 VTAIL.n190 VTAIL.n189 11.249
R643 VTAIL.n173 VTAIL.n114 11.249
R644 VTAIL.n144 VTAIL.n131 11.249
R645 VTAIL.n336 VTAIL.n320 10.4732
R646 VTAIL.n363 VTAIL.n308 10.4732
R647 VTAIL.n385 VTAIL.n298 10.4732
R648 VTAIL.n42 VTAIL.n26 10.4732
R649 VTAIL.n69 VTAIL.n14 10.4732
R650 VTAIL.n91 VTAIL.n4 10.4732
R651 VTAIL.n291 VTAIL.n204 10.4732
R652 VTAIL.n270 VTAIL.n215 10.4732
R653 VTAIL.n243 VTAIL.n227 10.4732
R654 VTAIL.n193 VTAIL.n106 10.4732
R655 VTAIL.n172 VTAIL.n117 10.4732
R656 VTAIL.n145 VTAIL.n129 10.4732
R657 VTAIL.n340 VTAIL.n339 9.69747
R658 VTAIL.n360 VTAIL.n359 9.69747
R659 VTAIL.n386 VTAIL.n296 9.69747
R660 VTAIL.n46 VTAIL.n45 9.69747
R661 VTAIL.n66 VTAIL.n65 9.69747
R662 VTAIL.n92 VTAIL.n2 9.69747
R663 VTAIL.n292 VTAIL.n202 9.69747
R664 VTAIL.n267 VTAIL.n266 9.69747
R665 VTAIL.n247 VTAIL.n246 9.69747
R666 VTAIL.n194 VTAIL.n104 9.69747
R667 VTAIL.n169 VTAIL.n168 9.69747
R668 VTAIL.n149 VTAIL.n148 9.69747
R669 VTAIL.n388 VTAIL.n387 9.45567
R670 VTAIL.n94 VTAIL.n93 9.45567
R671 VTAIL.n294 VTAIL.n293 9.45567
R672 VTAIL.n196 VTAIL.n195 9.45567
R673 VTAIL.n387 VTAIL.n386 9.3005
R674 VTAIL.n298 VTAIL.n297 9.3005
R675 VTAIL.n381 VTAIL.n380 9.3005
R676 VTAIL.n379 VTAIL.n378 9.3005
R677 VTAIL.n302 VTAIL.n301 9.3005
R678 VTAIL.n347 VTAIL.n346 9.3005
R679 VTAIL.n345 VTAIL.n344 9.3005
R680 VTAIL.n318 VTAIL.n317 9.3005
R681 VTAIL.n339 VTAIL.n338 9.3005
R682 VTAIL.n337 VTAIL.n336 9.3005
R683 VTAIL.n322 VTAIL.n321 9.3005
R684 VTAIL.n331 VTAIL.n330 9.3005
R685 VTAIL.n329 VTAIL.n328 9.3005
R686 VTAIL.n314 VTAIL.n313 9.3005
R687 VTAIL.n353 VTAIL.n352 9.3005
R688 VTAIL.n355 VTAIL.n354 9.3005
R689 VTAIL.n310 VTAIL.n309 9.3005
R690 VTAIL.n361 VTAIL.n360 9.3005
R691 VTAIL.n363 VTAIL.n362 9.3005
R692 VTAIL.n306 VTAIL.n305 9.3005
R693 VTAIL.n370 VTAIL.n369 9.3005
R694 VTAIL.n372 VTAIL.n371 9.3005
R695 VTAIL.n93 VTAIL.n92 9.3005
R696 VTAIL.n4 VTAIL.n3 9.3005
R697 VTAIL.n87 VTAIL.n86 9.3005
R698 VTAIL.n85 VTAIL.n84 9.3005
R699 VTAIL.n8 VTAIL.n7 9.3005
R700 VTAIL.n53 VTAIL.n52 9.3005
R701 VTAIL.n51 VTAIL.n50 9.3005
R702 VTAIL.n24 VTAIL.n23 9.3005
R703 VTAIL.n45 VTAIL.n44 9.3005
R704 VTAIL.n43 VTAIL.n42 9.3005
R705 VTAIL.n28 VTAIL.n27 9.3005
R706 VTAIL.n37 VTAIL.n36 9.3005
R707 VTAIL.n35 VTAIL.n34 9.3005
R708 VTAIL.n20 VTAIL.n19 9.3005
R709 VTAIL.n59 VTAIL.n58 9.3005
R710 VTAIL.n61 VTAIL.n60 9.3005
R711 VTAIL.n16 VTAIL.n15 9.3005
R712 VTAIL.n67 VTAIL.n66 9.3005
R713 VTAIL.n69 VTAIL.n68 9.3005
R714 VTAIL.n12 VTAIL.n11 9.3005
R715 VTAIL.n76 VTAIL.n75 9.3005
R716 VTAIL.n78 VTAIL.n77 9.3005
R717 VTAIL.n260 VTAIL.n259 9.3005
R718 VTAIL.n262 VTAIL.n261 9.3005
R719 VTAIL.n217 VTAIL.n216 9.3005
R720 VTAIL.n268 VTAIL.n267 9.3005
R721 VTAIL.n270 VTAIL.n269 9.3005
R722 VTAIL.n212 VTAIL.n211 9.3005
R723 VTAIL.n276 VTAIL.n275 9.3005
R724 VTAIL.n278 VTAIL.n277 9.3005
R725 VTAIL.n293 VTAIL.n292 9.3005
R726 VTAIL.n204 VTAIL.n203 9.3005
R727 VTAIL.n287 VTAIL.n286 9.3005
R728 VTAIL.n285 VTAIL.n284 9.3005
R729 VTAIL.n208 VTAIL.n207 9.3005
R730 VTAIL.n221 VTAIL.n220 9.3005
R731 VTAIL.n254 VTAIL.n253 9.3005
R732 VTAIL.n252 VTAIL.n251 9.3005
R733 VTAIL.n225 VTAIL.n224 9.3005
R734 VTAIL.n246 VTAIL.n245 9.3005
R735 VTAIL.n244 VTAIL.n243 9.3005
R736 VTAIL.n229 VTAIL.n228 9.3005
R737 VTAIL.n238 VTAIL.n237 9.3005
R738 VTAIL.n236 VTAIL.n235 9.3005
R739 VTAIL.n162 VTAIL.n161 9.3005
R740 VTAIL.n164 VTAIL.n163 9.3005
R741 VTAIL.n119 VTAIL.n118 9.3005
R742 VTAIL.n170 VTAIL.n169 9.3005
R743 VTAIL.n172 VTAIL.n171 9.3005
R744 VTAIL.n114 VTAIL.n113 9.3005
R745 VTAIL.n178 VTAIL.n177 9.3005
R746 VTAIL.n180 VTAIL.n179 9.3005
R747 VTAIL.n195 VTAIL.n194 9.3005
R748 VTAIL.n106 VTAIL.n105 9.3005
R749 VTAIL.n189 VTAIL.n188 9.3005
R750 VTAIL.n187 VTAIL.n186 9.3005
R751 VTAIL.n110 VTAIL.n109 9.3005
R752 VTAIL.n123 VTAIL.n122 9.3005
R753 VTAIL.n156 VTAIL.n155 9.3005
R754 VTAIL.n154 VTAIL.n153 9.3005
R755 VTAIL.n127 VTAIL.n126 9.3005
R756 VTAIL.n148 VTAIL.n147 9.3005
R757 VTAIL.n146 VTAIL.n145 9.3005
R758 VTAIL.n131 VTAIL.n130 9.3005
R759 VTAIL.n140 VTAIL.n139 9.3005
R760 VTAIL.n138 VTAIL.n137 9.3005
R761 VTAIL.n343 VTAIL.n318 8.92171
R762 VTAIL.n356 VTAIL.n310 8.92171
R763 VTAIL.n49 VTAIL.n24 8.92171
R764 VTAIL.n62 VTAIL.n16 8.92171
R765 VTAIL.n263 VTAIL.n217 8.92171
R766 VTAIL.n250 VTAIL.n225 8.92171
R767 VTAIL.n165 VTAIL.n119 8.92171
R768 VTAIL.n152 VTAIL.n127 8.92171
R769 VTAIL.n344 VTAIL.n316 8.14595
R770 VTAIL.n355 VTAIL.n312 8.14595
R771 VTAIL.n50 VTAIL.n22 8.14595
R772 VTAIL.n61 VTAIL.n18 8.14595
R773 VTAIL.n262 VTAIL.n219 8.14595
R774 VTAIL.n251 VTAIL.n223 8.14595
R775 VTAIL.n164 VTAIL.n121 8.14595
R776 VTAIL.n153 VTAIL.n125 8.14595
R777 VTAIL.n348 VTAIL.n347 7.3702
R778 VTAIL.n352 VTAIL.n351 7.3702
R779 VTAIL.n54 VTAIL.n53 7.3702
R780 VTAIL.n58 VTAIL.n57 7.3702
R781 VTAIL.n259 VTAIL.n258 7.3702
R782 VTAIL.n255 VTAIL.n254 7.3702
R783 VTAIL.n161 VTAIL.n160 7.3702
R784 VTAIL.n157 VTAIL.n156 7.3702
R785 VTAIL.n348 VTAIL.n314 6.59444
R786 VTAIL.n351 VTAIL.n314 6.59444
R787 VTAIL.n54 VTAIL.n20 6.59444
R788 VTAIL.n57 VTAIL.n20 6.59444
R789 VTAIL.n258 VTAIL.n221 6.59444
R790 VTAIL.n255 VTAIL.n221 6.59444
R791 VTAIL.n160 VTAIL.n123 6.59444
R792 VTAIL.n157 VTAIL.n123 6.59444
R793 VTAIL.n347 VTAIL.n316 5.81868
R794 VTAIL.n352 VTAIL.n312 5.81868
R795 VTAIL.n53 VTAIL.n22 5.81868
R796 VTAIL.n58 VTAIL.n18 5.81868
R797 VTAIL.n259 VTAIL.n219 5.81868
R798 VTAIL.n254 VTAIL.n223 5.81868
R799 VTAIL.n161 VTAIL.n121 5.81868
R800 VTAIL.n156 VTAIL.n125 5.81868
R801 VTAIL.n344 VTAIL.n343 5.04292
R802 VTAIL.n356 VTAIL.n355 5.04292
R803 VTAIL.n50 VTAIL.n49 5.04292
R804 VTAIL.n62 VTAIL.n61 5.04292
R805 VTAIL.n263 VTAIL.n262 5.04292
R806 VTAIL.n251 VTAIL.n250 5.04292
R807 VTAIL.n165 VTAIL.n164 5.04292
R808 VTAIL.n153 VTAIL.n152 5.04292
R809 VTAIL.n236 VTAIL.n232 4.38563
R810 VTAIL.n138 VTAIL.n134 4.38563
R811 VTAIL.n329 VTAIL.n325 4.38563
R812 VTAIL.n35 VTAIL.n31 4.38563
R813 VTAIL.n340 VTAIL.n318 4.26717
R814 VTAIL.n359 VTAIL.n310 4.26717
R815 VTAIL.n388 VTAIL.n296 4.26717
R816 VTAIL.n46 VTAIL.n24 4.26717
R817 VTAIL.n65 VTAIL.n16 4.26717
R818 VTAIL.n94 VTAIL.n2 4.26717
R819 VTAIL.n294 VTAIL.n202 4.26717
R820 VTAIL.n266 VTAIL.n217 4.26717
R821 VTAIL.n247 VTAIL.n225 4.26717
R822 VTAIL.n196 VTAIL.n104 4.26717
R823 VTAIL.n168 VTAIL.n119 4.26717
R824 VTAIL.n149 VTAIL.n127 4.26717
R825 VTAIL.n339 VTAIL.n320 3.49141
R826 VTAIL.n360 VTAIL.n308 3.49141
R827 VTAIL.n386 VTAIL.n385 3.49141
R828 VTAIL.n45 VTAIL.n26 3.49141
R829 VTAIL.n66 VTAIL.n14 3.49141
R830 VTAIL.n92 VTAIL.n91 3.49141
R831 VTAIL.n292 VTAIL.n291 3.49141
R832 VTAIL.n267 VTAIL.n215 3.49141
R833 VTAIL.n246 VTAIL.n227 3.49141
R834 VTAIL.n194 VTAIL.n193 3.49141
R835 VTAIL.n169 VTAIL.n117 3.49141
R836 VTAIL.n148 VTAIL.n129 3.49141
R837 VTAIL.n336 VTAIL.n335 2.71565
R838 VTAIL.n364 VTAIL.n363 2.71565
R839 VTAIL.n382 VTAIL.n298 2.71565
R840 VTAIL.n42 VTAIL.n41 2.71565
R841 VTAIL.n70 VTAIL.n69 2.71565
R842 VTAIL.n88 VTAIL.n4 2.71565
R843 VTAIL.n288 VTAIL.n204 2.71565
R844 VTAIL.n271 VTAIL.n270 2.71565
R845 VTAIL.n243 VTAIL.n242 2.71565
R846 VTAIL.n190 VTAIL.n106 2.71565
R847 VTAIL.n173 VTAIL.n172 2.71565
R848 VTAIL.n145 VTAIL.n144 2.71565
R849 VTAIL.n332 VTAIL.n322 1.93989
R850 VTAIL.n368 VTAIL.n306 1.93989
R851 VTAIL.n381 VTAIL.n300 1.93989
R852 VTAIL.n38 VTAIL.n28 1.93989
R853 VTAIL.n74 VTAIL.n12 1.93989
R854 VTAIL.n87 VTAIL.n6 1.93989
R855 VTAIL.n287 VTAIL.n206 1.93989
R856 VTAIL.n274 VTAIL.n212 1.93989
R857 VTAIL.n239 VTAIL.n229 1.93989
R858 VTAIL.n189 VTAIL.n108 1.93989
R859 VTAIL.n176 VTAIL.n114 1.93989
R860 VTAIL.n141 VTAIL.n131 1.93989
R861 VTAIL.n103 VTAIL.n101 1.47464
R862 VTAIL.n197 VTAIL.n103 1.47464
R863 VTAIL.n201 VTAIL.n199 1.47464
R864 VTAIL.n295 VTAIL.n201 1.47464
R865 VTAIL.n99 VTAIL.n97 1.47464
R866 VTAIL.n97 VTAIL.n95 1.47464
R867 VTAIL.n391 VTAIL.n389 1.47464
R868 VTAIL.n199 VTAIL.n197 1.2074
R869 VTAIL.n95 VTAIL.n1 1.2074
R870 VTAIL.n390 VTAIL.t8 1.17697
R871 VTAIL.n390 VTAIL.t0 1.17697
R872 VTAIL.n0 VTAIL.t1 1.17697
R873 VTAIL.n0 VTAIL.t6 1.17697
R874 VTAIL.n96 VTAIL.t18 1.17697
R875 VTAIL.n96 VTAIL.t12 1.17697
R876 VTAIL.n98 VTAIL.t17 1.17697
R877 VTAIL.n98 VTAIL.t19 1.17697
R878 VTAIL.n200 VTAIL.t13 1.17697
R879 VTAIL.n200 VTAIL.t10 1.17697
R880 VTAIL.n198 VTAIL.t14 1.17697
R881 VTAIL.n198 VTAIL.t11 1.17697
R882 VTAIL.n102 VTAIL.t7 1.17697
R883 VTAIL.n102 VTAIL.t4 1.17697
R884 VTAIL.n100 VTAIL.t2 1.17697
R885 VTAIL.n100 VTAIL.t3 1.17697
R886 VTAIL VTAIL.n1 1.16429
R887 VTAIL.n331 VTAIL.n324 1.16414
R888 VTAIL.n369 VTAIL.n304 1.16414
R889 VTAIL.n378 VTAIL.n377 1.16414
R890 VTAIL.n37 VTAIL.n30 1.16414
R891 VTAIL.n75 VTAIL.n10 1.16414
R892 VTAIL.n84 VTAIL.n83 1.16414
R893 VTAIL.n284 VTAIL.n283 1.16414
R894 VTAIL.n275 VTAIL.n210 1.16414
R895 VTAIL.n238 VTAIL.n231 1.16414
R896 VTAIL.n186 VTAIL.n185 1.16414
R897 VTAIL.n177 VTAIL.n112 1.16414
R898 VTAIL.n140 VTAIL.n133 1.16414
R899 VTAIL.n328 VTAIL.n327 0.388379
R900 VTAIL.n373 VTAIL.n372 0.388379
R901 VTAIL.n374 VTAIL.n302 0.388379
R902 VTAIL.n34 VTAIL.n33 0.388379
R903 VTAIL.n79 VTAIL.n78 0.388379
R904 VTAIL.n80 VTAIL.n8 0.388379
R905 VTAIL.n280 VTAIL.n208 0.388379
R906 VTAIL.n279 VTAIL.n278 0.388379
R907 VTAIL.n235 VTAIL.n234 0.388379
R908 VTAIL.n182 VTAIL.n110 0.388379
R909 VTAIL.n181 VTAIL.n180 0.388379
R910 VTAIL.n137 VTAIL.n136 0.388379
R911 VTAIL VTAIL.n391 0.310845
R912 VTAIL.n330 VTAIL.n329 0.155672
R913 VTAIL.n330 VTAIL.n321 0.155672
R914 VTAIL.n337 VTAIL.n321 0.155672
R915 VTAIL.n338 VTAIL.n337 0.155672
R916 VTAIL.n338 VTAIL.n317 0.155672
R917 VTAIL.n345 VTAIL.n317 0.155672
R918 VTAIL.n346 VTAIL.n345 0.155672
R919 VTAIL.n346 VTAIL.n313 0.155672
R920 VTAIL.n353 VTAIL.n313 0.155672
R921 VTAIL.n354 VTAIL.n353 0.155672
R922 VTAIL.n354 VTAIL.n309 0.155672
R923 VTAIL.n361 VTAIL.n309 0.155672
R924 VTAIL.n362 VTAIL.n361 0.155672
R925 VTAIL.n362 VTAIL.n305 0.155672
R926 VTAIL.n370 VTAIL.n305 0.155672
R927 VTAIL.n371 VTAIL.n370 0.155672
R928 VTAIL.n371 VTAIL.n301 0.155672
R929 VTAIL.n379 VTAIL.n301 0.155672
R930 VTAIL.n380 VTAIL.n379 0.155672
R931 VTAIL.n380 VTAIL.n297 0.155672
R932 VTAIL.n387 VTAIL.n297 0.155672
R933 VTAIL.n36 VTAIL.n35 0.155672
R934 VTAIL.n36 VTAIL.n27 0.155672
R935 VTAIL.n43 VTAIL.n27 0.155672
R936 VTAIL.n44 VTAIL.n43 0.155672
R937 VTAIL.n44 VTAIL.n23 0.155672
R938 VTAIL.n51 VTAIL.n23 0.155672
R939 VTAIL.n52 VTAIL.n51 0.155672
R940 VTAIL.n52 VTAIL.n19 0.155672
R941 VTAIL.n59 VTAIL.n19 0.155672
R942 VTAIL.n60 VTAIL.n59 0.155672
R943 VTAIL.n60 VTAIL.n15 0.155672
R944 VTAIL.n67 VTAIL.n15 0.155672
R945 VTAIL.n68 VTAIL.n67 0.155672
R946 VTAIL.n68 VTAIL.n11 0.155672
R947 VTAIL.n76 VTAIL.n11 0.155672
R948 VTAIL.n77 VTAIL.n76 0.155672
R949 VTAIL.n77 VTAIL.n7 0.155672
R950 VTAIL.n85 VTAIL.n7 0.155672
R951 VTAIL.n86 VTAIL.n85 0.155672
R952 VTAIL.n86 VTAIL.n3 0.155672
R953 VTAIL.n93 VTAIL.n3 0.155672
R954 VTAIL.n293 VTAIL.n203 0.155672
R955 VTAIL.n286 VTAIL.n203 0.155672
R956 VTAIL.n286 VTAIL.n285 0.155672
R957 VTAIL.n285 VTAIL.n207 0.155672
R958 VTAIL.n277 VTAIL.n207 0.155672
R959 VTAIL.n277 VTAIL.n276 0.155672
R960 VTAIL.n276 VTAIL.n211 0.155672
R961 VTAIL.n269 VTAIL.n211 0.155672
R962 VTAIL.n269 VTAIL.n268 0.155672
R963 VTAIL.n268 VTAIL.n216 0.155672
R964 VTAIL.n261 VTAIL.n216 0.155672
R965 VTAIL.n261 VTAIL.n260 0.155672
R966 VTAIL.n260 VTAIL.n220 0.155672
R967 VTAIL.n253 VTAIL.n220 0.155672
R968 VTAIL.n253 VTAIL.n252 0.155672
R969 VTAIL.n252 VTAIL.n224 0.155672
R970 VTAIL.n245 VTAIL.n224 0.155672
R971 VTAIL.n245 VTAIL.n244 0.155672
R972 VTAIL.n244 VTAIL.n228 0.155672
R973 VTAIL.n237 VTAIL.n228 0.155672
R974 VTAIL.n237 VTAIL.n236 0.155672
R975 VTAIL.n195 VTAIL.n105 0.155672
R976 VTAIL.n188 VTAIL.n105 0.155672
R977 VTAIL.n188 VTAIL.n187 0.155672
R978 VTAIL.n187 VTAIL.n109 0.155672
R979 VTAIL.n179 VTAIL.n109 0.155672
R980 VTAIL.n179 VTAIL.n178 0.155672
R981 VTAIL.n178 VTAIL.n113 0.155672
R982 VTAIL.n171 VTAIL.n113 0.155672
R983 VTAIL.n171 VTAIL.n170 0.155672
R984 VTAIL.n170 VTAIL.n118 0.155672
R985 VTAIL.n163 VTAIL.n118 0.155672
R986 VTAIL.n163 VTAIL.n162 0.155672
R987 VTAIL.n162 VTAIL.n122 0.155672
R988 VTAIL.n155 VTAIL.n122 0.155672
R989 VTAIL.n155 VTAIL.n154 0.155672
R990 VTAIL.n154 VTAIL.n126 0.155672
R991 VTAIL.n147 VTAIL.n126 0.155672
R992 VTAIL.n147 VTAIL.n146 0.155672
R993 VTAIL.n146 VTAIL.n130 0.155672
R994 VTAIL.n139 VTAIL.n130 0.155672
R995 VTAIL.n139 VTAIL.n138 0.155672
R996 B.n681 B.n136 585
R997 B.n136 B.n71 585
R998 B.n683 B.n682 585
R999 B.n685 B.n135 585
R1000 B.n688 B.n687 585
R1001 B.n689 B.n134 585
R1002 B.n691 B.n690 585
R1003 B.n693 B.n133 585
R1004 B.n696 B.n695 585
R1005 B.n697 B.n132 585
R1006 B.n699 B.n698 585
R1007 B.n701 B.n131 585
R1008 B.n704 B.n703 585
R1009 B.n705 B.n130 585
R1010 B.n707 B.n706 585
R1011 B.n709 B.n129 585
R1012 B.n712 B.n711 585
R1013 B.n713 B.n128 585
R1014 B.n715 B.n714 585
R1015 B.n717 B.n127 585
R1016 B.n720 B.n719 585
R1017 B.n721 B.n126 585
R1018 B.n723 B.n722 585
R1019 B.n725 B.n125 585
R1020 B.n728 B.n727 585
R1021 B.n729 B.n124 585
R1022 B.n731 B.n730 585
R1023 B.n733 B.n123 585
R1024 B.n736 B.n735 585
R1025 B.n737 B.n122 585
R1026 B.n739 B.n738 585
R1027 B.n741 B.n121 585
R1028 B.n744 B.n743 585
R1029 B.n745 B.n120 585
R1030 B.n747 B.n746 585
R1031 B.n749 B.n119 585
R1032 B.n752 B.n751 585
R1033 B.n753 B.n118 585
R1034 B.n755 B.n754 585
R1035 B.n757 B.n117 585
R1036 B.n760 B.n759 585
R1037 B.n761 B.n116 585
R1038 B.n763 B.n762 585
R1039 B.n765 B.n115 585
R1040 B.n768 B.n767 585
R1041 B.n769 B.n114 585
R1042 B.n771 B.n770 585
R1043 B.n773 B.n113 585
R1044 B.n776 B.n775 585
R1045 B.n777 B.n112 585
R1046 B.n779 B.n778 585
R1047 B.n781 B.n111 585
R1048 B.n784 B.n783 585
R1049 B.n785 B.n110 585
R1050 B.n787 B.n786 585
R1051 B.n789 B.n109 585
R1052 B.n792 B.n791 585
R1053 B.n794 B.n106 585
R1054 B.n796 B.n795 585
R1055 B.n798 B.n105 585
R1056 B.n801 B.n800 585
R1057 B.n802 B.n104 585
R1058 B.n804 B.n803 585
R1059 B.n806 B.n103 585
R1060 B.n809 B.n808 585
R1061 B.n810 B.n100 585
R1062 B.n813 B.n812 585
R1063 B.n815 B.n99 585
R1064 B.n818 B.n817 585
R1065 B.n819 B.n98 585
R1066 B.n821 B.n820 585
R1067 B.n823 B.n97 585
R1068 B.n826 B.n825 585
R1069 B.n827 B.n96 585
R1070 B.n829 B.n828 585
R1071 B.n831 B.n95 585
R1072 B.n834 B.n833 585
R1073 B.n835 B.n94 585
R1074 B.n837 B.n836 585
R1075 B.n839 B.n93 585
R1076 B.n842 B.n841 585
R1077 B.n843 B.n92 585
R1078 B.n845 B.n844 585
R1079 B.n847 B.n91 585
R1080 B.n850 B.n849 585
R1081 B.n851 B.n90 585
R1082 B.n853 B.n852 585
R1083 B.n855 B.n89 585
R1084 B.n858 B.n857 585
R1085 B.n859 B.n88 585
R1086 B.n861 B.n860 585
R1087 B.n863 B.n87 585
R1088 B.n866 B.n865 585
R1089 B.n867 B.n86 585
R1090 B.n869 B.n868 585
R1091 B.n871 B.n85 585
R1092 B.n874 B.n873 585
R1093 B.n875 B.n84 585
R1094 B.n877 B.n876 585
R1095 B.n879 B.n83 585
R1096 B.n882 B.n881 585
R1097 B.n883 B.n82 585
R1098 B.n885 B.n884 585
R1099 B.n887 B.n81 585
R1100 B.n890 B.n889 585
R1101 B.n891 B.n80 585
R1102 B.n893 B.n892 585
R1103 B.n895 B.n79 585
R1104 B.n898 B.n897 585
R1105 B.n899 B.n78 585
R1106 B.n901 B.n900 585
R1107 B.n903 B.n77 585
R1108 B.n906 B.n905 585
R1109 B.n907 B.n76 585
R1110 B.n909 B.n908 585
R1111 B.n911 B.n75 585
R1112 B.n914 B.n913 585
R1113 B.n915 B.n74 585
R1114 B.n917 B.n916 585
R1115 B.n919 B.n73 585
R1116 B.n922 B.n921 585
R1117 B.n923 B.n72 585
R1118 B.n680 B.n70 585
R1119 B.n926 B.n70 585
R1120 B.n679 B.n69 585
R1121 B.n927 B.n69 585
R1122 B.n678 B.n68 585
R1123 B.n928 B.n68 585
R1124 B.n677 B.n676 585
R1125 B.n676 B.n64 585
R1126 B.n675 B.n63 585
R1127 B.n934 B.n63 585
R1128 B.n674 B.n62 585
R1129 B.n935 B.n62 585
R1130 B.n673 B.n61 585
R1131 B.n936 B.n61 585
R1132 B.n672 B.n671 585
R1133 B.n671 B.n57 585
R1134 B.n670 B.n56 585
R1135 B.n942 B.n56 585
R1136 B.n669 B.n55 585
R1137 B.n943 B.n55 585
R1138 B.n668 B.n54 585
R1139 B.n944 B.n54 585
R1140 B.n667 B.n666 585
R1141 B.n666 B.n50 585
R1142 B.n665 B.n49 585
R1143 B.n950 B.n49 585
R1144 B.n664 B.n48 585
R1145 B.n951 B.n48 585
R1146 B.n663 B.n47 585
R1147 B.n952 B.n47 585
R1148 B.n662 B.n661 585
R1149 B.n661 B.n43 585
R1150 B.n660 B.n42 585
R1151 B.n958 B.n42 585
R1152 B.n659 B.n41 585
R1153 B.n959 B.n41 585
R1154 B.n658 B.n40 585
R1155 B.n960 B.n40 585
R1156 B.n657 B.n656 585
R1157 B.n656 B.n36 585
R1158 B.n655 B.n35 585
R1159 B.n966 B.n35 585
R1160 B.n654 B.n34 585
R1161 B.n967 B.n34 585
R1162 B.n653 B.n33 585
R1163 B.n968 B.n33 585
R1164 B.n652 B.n651 585
R1165 B.n651 B.n32 585
R1166 B.n650 B.n28 585
R1167 B.n974 B.n28 585
R1168 B.n649 B.n27 585
R1169 B.n975 B.n27 585
R1170 B.n648 B.n26 585
R1171 B.n976 B.n26 585
R1172 B.n647 B.n646 585
R1173 B.n646 B.n22 585
R1174 B.n645 B.n21 585
R1175 B.n982 B.n21 585
R1176 B.n644 B.n20 585
R1177 B.n983 B.n20 585
R1178 B.n643 B.n19 585
R1179 B.n984 B.n19 585
R1180 B.n642 B.n641 585
R1181 B.n641 B.n15 585
R1182 B.n640 B.n14 585
R1183 B.n990 B.n14 585
R1184 B.n639 B.n13 585
R1185 B.n991 B.n13 585
R1186 B.n638 B.n12 585
R1187 B.n992 B.n12 585
R1188 B.n637 B.n636 585
R1189 B.n636 B.n8 585
R1190 B.n635 B.n7 585
R1191 B.n998 B.n7 585
R1192 B.n634 B.n6 585
R1193 B.n999 B.n6 585
R1194 B.n633 B.n5 585
R1195 B.n1000 B.n5 585
R1196 B.n632 B.n631 585
R1197 B.n631 B.n4 585
R1198 B.n630 B.n137 585
R1199 B.n630 B.n629 585
R1200 B.n620 B.n138 585
R1201 B.n139 B.n138 585
R1202 B.n622 B.n621 585
R1203 B.n623 B.n622 585
R1204 B.n619 B.n143 585
R1205 B.n147 B.n143 585
R1206 B.n618 B.n617 585
R1207 B.n617 B.n616 585
R1208 B.n145 B.n144 585
R1209 B.n146 B.n145 585
R1210 B.n609 B.n608 585
R1211 B.n610 B.n609 585
R1212 B.n607 B.n152 585
R1213 B.n152 B.n151 585
R1214 B.n606 B.n605 585
R1215 B.n605 B.n604 585
R1216 B.n154 B.n153 585
R1217 B.n155 B.n154 585
R1218 B.n597 B.n596 585
R1219 B.n598 B.n597 585
R1220 B.n595 B.n160 585
R1221 B.n160 B.n159 585
R1222 B.n594 B.n593 585
R1223 B.n593 B.n592 585
R1224 B.n162 B.n161 585
R1225 B.n585 B.n162 585
R1226 B.n584 B.n583 585
R1227 B.n586 B.n584 585
R1228 B.n582 B.n167 585
R1229 B.n167 B.n166 585
R1230 B.n581 B.n580 585
R1231 B.n580 B.n579 585
R1232 B.n169 B.n168 585
R1233 B.n170 B.n169 585
R1234 B.n572 B.n571 585
R1235 B.n573 B.n572 585
R1236 B.n570 B.n175 585
R1237 B.n175 B.n174 585
R1238 B.n569 B.n568 585
R1239 B.n568 B.n567 585
R1240 B.n177 B.n176 585
R1241 B.n178 B.n177 585
R1242 B.n560 B.n559 585
R1243 B.n561 B.n560 585
R1244 B.n558 B.n182 585
R1245 B.n186 B.n182 585
R1246 B.n557 B.n556 585
R1247 B.n556 B.n555 585
R1248 B.n184 B.n183 585
R1249 B.n185 B.n184 585
R1250 B.n548 B.n547 585
R1251 B.n549 B.n548 585
R1252 B.n546 B.n191 585
R1253 B.n191 B.n190 585
R1254 B.n545 B.n544 585
R1255 B.n544 B.n543 585
R1256 B.n193 B.n192 585
R1257 B.n194 B.n193 585
R1258 B.n536 B.n535 585
R1259 B.n537 B.n536 585
R1260 B.n534 B.n198 585
R1261 B.n202 B.n198 585
R1262 B.n533 B.n532 585
R1263 B.n532 B.n531 585
R1264 B.n200 B.n199 585
R1265 B.n201 B.n200 585
R1266 B.n524 B.n523 585
R1267 B.n525 B.n524 585
R1268 B.n522 B.n207 585
R1269 B.n207 B.n206 585
R1270 B.n521 B.n520 585
R1271 B.n520 B.n519 585
R1272 B.n516 B.n211 585
R1273 B.n515 B.n514 585
R1274 B.n512 B.n212 585
R1275 B.n512 B.n210 585
R1276 B.n511 B.n510 585
R1277 B.n509 B.n508 585
R1278 B.n507 B.n214 585
R1279 B.n505 B.n504 585
R1280 B.n503 B.n215 585
R1281 B.n502 B.n501 585
R1282 B.n499 B.n216 585
R1283 B.n497 B.n496 585
R1284 B.n495 B.n217 585
R1285 B.n494 B.n493 585
R1286 B.n491 B.n218 585
R1287 B.n489 B.n488 585
R1288 B.n487 B.n219 585
R1289 B.n486 B.n485 585
R1290 B.n483 B.n220 585
R1291 B.n481 B.n480 585
R1292 B.n479 B.n221 585
R1293 B.n478 B.n477 585
R1294 B.n475 B.n222 585
R1295 B.n473 B.n472 585
R1296 B.n471 B.n223 585
R1297 B.n470 B.n469 585
R1298 B.n467 B.n224 585
R1299 B.n465 B.n464 585
R1300 B.n463 B.n225 585
R1301 B.n462 B.n461 585
R1302 B.n459 B.n226 585
R1303 B.n457 B.n456 585
R1304 B.n455 B.n227 585
R1305 B.n454 B.n453 585
R1306 B.n451 B.n228 585
R1307 B.n449 B.n448 585
R1308 B.n447 B.n229 585
R1309 B.n446 B.n445 585
R1310 B.n443 B.n230 585
R1311 B.n441 B.n440 585
R1312 B.n439 B.n231 585
R1313 B.n438 B.n437 585
R1314 B.n435 B.n232 585
R1315 B.n433 B.n432 585
R1316 B.n431 B.n233 585
R1317 B.n430 B.n429 585
R1318 B.n427 B.n234 585
R1319 B.n425 B.n424 585
R1320 B.n423 B.n235 585
R1321 B.n422 B.n421 585
R1322 B.n419 B.n236 585
R1323 B.n417 B.n416 585
R1324 B.n415 B.n237 585
R1325 B.n414 B.n413 585
R1326 B.n411 B.n238 585
R1327 B.n409 B.n408 585
R1328 B.n407 B.n239 585
R1329 B.n405 B.n404 585
R1330 B.n402 B.n242 585
R1331 B.n400 B.n399 585
R1332 B.n398 B.n243 585
R1333 B.n397 B.n396 585
R1334 B.n394 B.n244 585
R1335 B.n392 B.n391 585
R1336 B.n390 B.n245 585
R1337 B.n389 B.n388 585
R1338 B.n386 B.n385 585
R1339 B.n384 B.n383 585
R1340 B.n382 B.n250 585
R1341 B.n380 B.n379 585
R1342 B.n378 B.n251 585
R1343 B.n377 B.n376 585
R1344 B.n374 B.n252 585
R1345 B.n372 B.n371 585
R1346 B.n370 B.n253 585
R1347 B.n369 B.n368 585
R1348 B.n366 B.n254 585
R1349 B.n364 B.n363 585
R1350 B.n362 B.n255 585
R1351 B.n361 B.n360 585
R1352 B.n358 B.n256 585
R1353 B.n356 B.n355 585
R1354 B.n354 B.n257 585
R1355 B.n353 B.n352 585
R1356 B.n350 B.n258 585
R1357 B.n348 B.n347 585
R1358 B.n346 B.n259 585
R1359 B.n345 B.n344 585
R1360 B.n342 B.n260 585
R1361 B.n340 B.n339 585
R1362 B.n338 B.n261 585
R1363 B.n337 B.n336 585
R1364 B.n334 B.n262 585
R1365 B.n332 B.n331 585
R1366 B.n330 B.n263 585
R1367 B.n329 B.n328 585
R1368 B.n326 B.n264 585
R1369 B.n324 B.n323 585
R1370 B.n322 B.n265 585
R1371 B.n321 B.n320 585
R1372 B.n318 B.n266 585
R1373 B.n316 B.n315 585
R1374 B.n314 B.n267 585
R1375 B.n313 B.n312 585
R1376 B.n310 B.n268 585
R1377 B.n308 B.n307 585
R1378 B.n306 B.n269 585
R1379 B.n305 B.n304 585
R1380 B.n302 B.n270 585
R1381 B.n300 B.n299 585
R1382 B.n298 B.n271 585
R1383 B.n297 B.n296 585
R1384 B.n294 B.n272 585
R1385 B.n292 B.n291 585
R1386 B.n290 B.n273 585
R1387 B.n289 B.n288 585
R1388 B.n286 B.n274 585
R1389 B.n284 B.n283 585
R1390 B.n282 B.n275 585
R1391 B.n281 B.n280 585
R1392 B.n278 B.n276 585
R1393 B.n209 B.n208 585
R1394 B.n518 B.n517 585
R1395 B.n519 B.n518 585
R1396 B.n205 B.n204 585
R1397 B.n206 B.n205 585
R1398 B.n527 B.n526 585
R1399 B.n526 B.n525 585
R1400 B.n528 B.n203 585
R1401 B.n203 B.n201 585
R1402 B.n530 B.n529 585
R1403 B.n531 B.n530 585
R1404 B.n197 B.n196 585
R1405 B.n202 B.n197 585
R1406 B.n539 B.n538 585
R1407 B.n538 B.n537 585
R1408 B.n540 B.n195 585
R1409 B.n195 B.n194 585
R1410 B.n542 B.n541 585
R1411 B.n543 B.n542 585
R1412 B.n189 B.n188 585
R1413 B.n190 B.n189 585
R1414 B.n551 B.n550 585
R1415 B.n550 B.n549 585
R1416 B.n552 B.n187 585
R1417 B.n187 B.n185 585
R1418 B.n554 B.n553 585
R1419 B.n555 B.n554 585
R1420 B.n181 B.n180 585
R1421 B.n186 B.n181 585
R1422 B.n563 B.n562 585
R1423 B.n562 B.n561 585
R1424 B.n564 B.n179 585
R1425 B.n179 B.n178 585
R1426 B.n566 B.n565 585
R1427 B.n567 B.n566 585
R1428 B.n173 B.n172 585
R1429 B.n174 B.n173 585
R1430 B.n575 B.n574 585
R1431 B.n574 B.n573 585
R1432 B.n576 B.n171 585
R1433 B.n171 B.n170 585
R1434 B.n578 B.n577 585
R1435 B.n579 B.n578 585
R1436 B.n165 B.n164 585
R1437 B.n166 B.n165 585
R1438 B.n588 B.n587 585
R1439 B.n587 B.n586 585
R1440 B.n589 B.n163 585
R1441 B.n585 B.n163 585
R1442 B.n591 B.n590 585
R1443 B.n592 B.n591 585
R1444 B.n158 B.n157 585
R1445 B.n159 B.n158 585
R1446 B.n600 B.n599 585
R1447 B.n599 B.n598 585
R1448 B.n601 B.n156 585
R1449 B.n156 B.n155 585
R1450 B.n603 B.n602 585
R1451 B.n604 B.n603 585
R1452 B.n150 B.n149 585
R1453 B.n151 B.n150 585
R1454 B.n612 B.n611 585
R1455 B.n611 B.n610 585
R1456 B.n613 B.n148 585
R1457 B.n148 B.n146 585
R1458 B.n615 B.n614 585
R1459 B.n616 B.n615 585
R1460 B.n142 B.n141 585
R1461 B.n147 B.n142 585
R1462 B.n625 B.n624 585
R1463 B.n624 B.n623 585
R1464 B.n626 B.n140 585
R1465 B.n140 B.n139 585
R1466 B.n628 B.n627 585
R1467 B.n629 B.n628 585
R1468 B.n2 B.n0 585
R1469 B.n4 B.n2 585
R1470 B.n3 B.n1 585
R1471 B.n999 B.n3 585
R1472 B.n997 B.n996 585
R1473 B.n998 B.n997 585
R1474 B.n995 B.n9 585
R1475 B.n9 B.n8 585
R1476 B.n994 B.n993 585
R1477 B.n993 B.n992 585
R1478 B.n11 B.n10 585
R1479 B.n991 B.n11 585
R1480 B.n989 B.n988 585
R1481 B.n990 B.n989 585
R1482 B.n987 B.n16 585
R1483 B.n16 B.n15 585
R1484 B.n986 B.n985 585
R1485 B.n985 B.n984 585
R1486 B.n18 B.n17 585
R1487 B.n983 B.n18 585
R1488 B.n981 B.n980 585
R1489 B.n982 B.n981 585
R1490 B.n979 B.n23 585
R1491 B.n23 B.n22 585
R1492 B.n978 B.n977 585
R1493 B.n977 B.n976 585
R1494 B.n25 B.n24 585
R1495 B.n975 B.n25 585
R1496 B.n973 B.n972 585
R1497 B.n974 B.n973 585
R1498 B.n971 B.n29 585
R1499 B.n32 B.n29 585
R1500 B.n970 B.n969 585
R1501 B.n969 B.n968 585
R1502 B.n31 B.n30 585
R1503 B.n967 B.n31 585
R1504 B.n965 B.n964 585
R1505 B.n966 B.n965 585
R1506 B.n963 B.n37 585
R1507 B.n37 B.n36 585
R1508 B.n962 B.n961 585
R1509 B.n961 B.n960 585
R1510 B.n39 B.n38 585
R1511 B.n959 B.n39 585
R1512 B.n957 B.n956 585
R1513 B.n958 B.n957 585
R1514 B.n955 B.n44 585
R1515 B.n44 B.n43 585
R1516 B.n954 B.n953 585
R1517 B.n953 B.n952 585
R1518 B.n46 B.n45 585
R1519 B.n951 B.n46 585
R1520 B.n949 B.n948 585
R1521 B.n950 B.n949 585
R1522 B.n947 B.n51 585
R1523 B.n51 B.n50 585
R1524 B.n946 B.n945 585
R1525 B.n945 B.n944 585
R1526 B.n53 B.n52 585
R1527 B.n943 B.n53 585
R1528 B.n941 B.n940 585
R1529 B.n942 B.n941 585
R1530 B.n939 B.n58 585
R1531 B.n58 B.n57 585
R1532 B.n938 B.n937 585
R1533 B.n937 B.n936 585
R1534 B.n60 B.n59 585
R1535 B.n935 B.n60 585
R1536 B.n933 B.n932 585
R1537 B.n934 B.n933 585
R1538 B.n931 B.n65 585
R1539 B.n65 B.n64 585
R1540 B.n930 B.n929 585
R1541 B.n929 B.n928 585
R1542 B.n67 B.n66 585
R1543 B.n927 B.n67 585
R1544 B.n925 B.n924 585
R1545 B.n926 B.n925 585
R1546 B.n1002 B.n1001 585
R1547 B.n1001 B.n1000 585
R1548 B.n518 B.n211 564.573
R1549 B.n925 B.n72 564.573
R1550 B.n520 B.n209 564.573
R1551 B.n136 B.n70 564.573
R1552 B.n246 B.t21 498.878
R1553 B.n240 B.t10 498.878
R1554 B.n101 B.t18 498.878
R1555 B.n107 B.t14 498.878
R1556 B.n246 B.t23 398.517
R1557 B.n240 B.t13 398.517
R1558 B.n101 B.t19 398.517
R1559 B.n107 B.t16 398.517
R1560 B.n247 B.t22 365.353
R1561 B.n108 B.t17 365.353
R1562 B.n241 B.t12 365.353
R1563 B.n102 B.t20 365.353
R1564 B.n684 B.n71 256.663
R1565 B.n686 B.n71 256.663
R1566 B.n692 B.n71 256.663
R1567 B.n694 B.n71 256.663
R1568 B.n700 B.n71 256.663
R1569 B.n702 B.n71 256.663
R1570 B.n708 B.n71 256.663
R1571 B.n710 B.n71 256.663
R1572 B.n716 B.n71 256.663
R1573 B.n718 B.n71 256.663
R1574 B.n724 B.n71 256.663
R1575 B.n726 B.n71 256.663
R1576 B.n732 B.n71 256.663
R1577 B.n734 B.n71 256.663
R1578 B.n740 B.n71 256.663
R1579 B.n742 B.n71 256.663
R1580 B.n748 B.n71 256.663
R1581 B.n750 B.n71 256.663
R1582 B.n756 B.n71 256.663
R1583 B.n758 B.n71 256.663
R1584 B.n764 B.n71 256.663
R1585 B.n766 B.n71 256.663
R1586 B.n772 B.n71 256.663
R1587 B.n774 B.n71 256.663
R1588 B.n780 B.n71 256.663
R1589 B.n782 B.n71 256.663
R1590 B.n788 B.n71 256.663
R1591 B.n790 B.n71 256.663
R1592 B.n797 B.n71 256.663
R1593 B.n799 B.n71 256.663
R1594 B.n805 B.n71 256.663
R1595 B.n807 B.n71 256.663
R1596 B.n814 B.n71 256.663
R1597 B.n816 B.n71 256.663
R1598 B.n822 B.n71 256.663
R1599 B.n824 B.n71 256.663
R1600 B.n830 B.n71 256.663
R1601 B.n832 B.n71 256.663
R1602 B.n838 B.n71 256.663
R1603 B.n840 B.n71 256.663
R1604 B.n846 B.n71 256.663
R1605 B.n848 B.n71 256.663
R1606 B.n854 B.n71 256.663
R1607 B.n856 B.n71 256.663
R1608 B.n862 B.n71 256.663
R1609 B.n864 B.n71 256.663
R1610 B.n870 B.n71 256.663
R1611 B.n872 B.n71 256.663
R1612 B.n878 B.n71 256.663
R1613 B.n880 B.n71 256.663
R1614 B.n886 B.n71 256.663
R1615 B.n888 B.n71 256.663
R1616 B.n894 B.n71 256.663
R1617 B.n896 B.n71 256.663
R1618 B.n902 B.n71 256.663
R1619 B.n904 B.n71 256.663
R1620 B.n910 B.n71 256.663
R1621 B.n912 B.n71 256.663
R1622 B.n918 B.n71 256.663
R1623 B.n920 B.n71 256.663
R1624 B.n513 B.n210 256.663
R1625 B.n213 B.n210 256.663
R1626 B.n506 B.n210 256.663
R1627 B.n500 B.n210 256.663
R1628 B.n498 B.n210 256.663
R1629 B.n492 B.n210 256.663
R1630 B.n490 B.n210 256.663
R1631 B.n484 B.n210 256.663
R1632 B.n482 B.n210 256.663
R1633 B.n476 B.n210 256.663
R1634 B.n474 B.n210 256.663
R1635 B.n468 B.n210 256.663
R1636 B.n466 B.n210 256.663
R1637 B.n460 B.n210 256.663
R1638 B.n458 B.n210 256.663
R1639 B.n452 B.n210 256.663
R1640 B.n450 B.n210 256.663
R1641 B.n444 B.n210 256.663
R1642 B.n442 B.n210 256.663
R1643 B.n436 B.n210 256.663
R1644 B.n434 B.n210 256.663
R1645 B.n428 B.n210 256.663
R1646 B.n426 B.n210 256.663
R1647 B.n420 B.n210 256.663
R1648 B.n418 B.n210 256.663
R1649 B.n412 B.n210 256.663
R1650 B.n410 B.n210 256.663
R1651 B.n403 B.n210 256.663
R1652 B.n401 B.n210 256.663
R1653 B.n395 B.n210 256.663
R1654 B.n393 B.n210 256.663
R1655 B.n387 B.n210 256.663
R1656 B.n249 B.n210 256.663
R1657 B.n381 B.n210 256.663
R1658 B.n375 B.n210 256.663
R1659 B.n373 B.n210 256.663
R1660 B.n367 B.n210 256.663
R1661 B.n365 B.n210 256.663
R1662 B.n359 B.n210 256.663
R1663 B.n357 B.n210 256.663
R1664 B.n351 B.n210 256.663
R1665 B.n349 B.n210 256.663
R1666 B.n343 B.n210 256.663
R1667 B.n341 B.n210 256.663
R1668 B.n335 B.n210 256.663
R1669 B.n333 B.n210 256.663
R1670 B.n327 B.n210 256.663
R1671 B.n325 B.n210 256.663
R1672 B.n319 B.n210 256.663
R1673 B.n317 B.n210 256.663
R1674 B.n311 B.n210 256.663
R1675 B.n309 B.n210 256.663
R1676 B.n303 B.n210 256.663
R1677 B.n301 B.n210 256.663
R1678 B.n295 B.n210 256.663
R1679 B.n293 B.n210 256.663
R1680 B.n287 B.n210 256.663
R1681 B.n285 B.n210 256.663
R1682 B.n279 B.n210 256.663
R1683 B.n277 B.n210 256.663
R1684 B.n518 B.n205 163.367
R1685 B.n526 B.n205 163.367
R1686 B.n526 B.n203 163.367
R1687 B.n530 B.n203 163.367
R1688 B.n530 B.n197 163.367
R1689 B.n538 B.n197 163.367
R1690 B.n538 B.n195 163.367
R1691 B.n542 B.n195 163.367
R1692 B.n542 B.n189 163.367
R1693 B.n550 B.n189 163.367
R1694 B.n550 B.n187 163.367
R1695 B.n554 B.n187 163.367
R1696 B.n554 B.n181 163.367
R1697 B.n562 B.n181 163.367
R1698 B.n562 B.n179 163.367
R1699 B.n566 B.n179 163.367
R1700 B.n566 B.n173 163.367
R1701 B.n574 B.n173 163.367
R1702 B.n574 B.n171 163.367
R1703 B.n578 B.n171 163.367
R1704 B.n578 B.n165 163.367
R1705 B.n587 B.n165 163.367
R1706 B.n587 B.n163 163.367
R1707 B.n591 B.n163 163.367
R1708 B.n591 B.n158 163.367
R1709 B.n599 B.n158 163.367
R1710 B.n599 B.n156 163.367
R1711 B.n603 B.n156 163.367
R1712 B.n603 B.n150 163.367
R1713 B.n611 B.n150 163.367
R1714 B.n611 B.n148 163.367
R1715 B.n615 B.n148 163.367
R1716 B.n615 B.n142 163.367
R1717 B.n624 B.n142 163.367
R1718 B.n624 B.n140 163.367
R1719 B.n628 B.n140 163.367
R1720 B.n628 B.n2 163.367
R1721 B.n1001 B.n2 163.367
R1722 B.n1001 B.n3 163.367
R1723 B.n997 B.n3 163.367
R1724 B.n997 B.n9 163.367
R1725 B.n993 B.n9 163.367
R1726 B.n993 B.n11 163.367
R1727 B.n989 B.n11 163.367
R1728 B.n989 B.n16 163.367
R1729 B.n985 B.n16 163.367
R1730 B.n985 B.n18 163.367
R1731 B.n981 B.n18 163.367
R1732 B.n981 B.n23 163.367
R1733 B.n977 B.n23 163.367
R1734 B.n977 B.n25 163.367
R1735 B.n973 B.n25 163.367
R1736 B.n973 B.n29 163.367
R1737 B.n969 B.n29 163.367
R1738 B.n969 B.n31 163.367
R1739 B.n965 B.n31 163.367
R1740 B.n965 B.n37 163.367
R1741 B.n961 B.n37 163.367
R1742 B.n961 B.n39 163.367
R1743 B.n957 B.n39 163.367
R1744 B.n957 B.n44 163.367
R1745 B.n953 B.n44 163.367
R1746 B.n953 B.n46 163.367
R1747 B.n949 B.n46 163.367
R1748 B.n949 B.n51 163.367
R1749 B.n945 B.n51 163.367
R1750 B.n945 B.n53 163.367
R1751 B.n941 B.n53 163.367
R1752 B.n941 B.n58 163.367
R1753 B.n937 B.n58 163.367
R1754 B.n937 B.n60 163.367
R1755 B.n933 B.n60 163.367
R1756 B.n933 B.n65 163.367
R1757 B.n929 B.n65 163.367
R1758 B.n929 B.n67 163.367
R1759 B.n925 B.n67 163.367
R1760 B.n514 B.n512 163.367
R1761 B.n512 B.n511 163.367
R1762 B.n508 B.n507 163.367
R1763 B.n505 B.n215 163.367
R1764 B.n501 B.n499 163.367
R1765 B.n497 B.n217 163.367
R1766 B.n493 B.n491 163.367
R1767 B.n489 B.n219 163.367
R1768 B.n485 B.n483 163.367
R1769 B.n481 B.n221 163.367
R1770 B.n477 B.n475 163.367
R1771 B.n473 B.n223 163.367
R1772 B.n469 B.n467 163.367
R1773 B.n465 B.n225 163.367
R1774 B.n461 B.n459 163.367
R1775 B.n457 B.n227 163.367
R1776 B.n453 B.n451 163.367
R1777 B.n449 B.n229 163.367
R1778 B.n445 B.n443 163.367
R1779 B.n441 B.n231 163.367
R1780 B.n437 B.n435 163.367
R1781 B.n433 B.n233 163.367
R1782 B.n429 B.n427 163.367
R1783 B.n425 B.n235 163.367
R1784 B.n421 B.n419 163.367
R1785 B.n417 B.n237 163.367
R1786 B.n413 B.n411 163.367
R1787 B.n409 B.n239 163.367
R1788 B.n404 B.n402 163.367
R1789 B.n400 B.n243 163.367
R1790 B.n396 B.n394 163.367
R1791 B.n392 B.n245 163.367
R1792 B.n388 B.n386 163.367
R1793 B.n383 B.n382 163.367
R1794 B.n380 B.n251 163.367
R1795 B.n376 B.n374 163.367
R1796 B.n372 B.n253 163.367
R1797 B.n368 B.n366 163.367
R1798 B.n364 B.n255 163.367
R1799 B.n360 B.n358 163.367
R1800 B.n356 B.n257 163.367
R1801 B.n352 B.n350 163.367
R1802 B.n348 B.n259 163.367
R1803 B.n344 B.n342 163.367
R1804 B.n340 B.n261 163.367
R1805 B.n336 B.n334 163.367
R1806 B.n332 B.n263 163.367
R1807 B.n328 B.n326 163.367
R1808 B.n324 B.n265 163.367
R1809 B.n320 B.n318 163.367
R1810 B.n316 B.n267 163.367
R1811 B.n312 B.n310 163.367
R1812 B.n308 B.n269 163.367
R1813 B.n304 B.n302 163.367
R1814 B.n300 B.n271 163.367
R1815 B.n296 B.n294 163.367
R1816 B.n292 B.n273 163.367
R1817 B.n288 B.n286 163.367
R1818 B.n284 B.n275 163.367
R1819 B.n280 B.n278 163.367
R1820 B.n520 B.n207 163.367
R1821 B.n524 B.n207 163.367
R1822 B.n524 B.n200 163.367
R1823 B.n532 B.n200 163.367
R1824 B.n532 B.n198 163.367
R1825 B.n536 B.n198 163.367
R1826 B.n536 B.n193 163.367
R1827 B.n544 B.n193 163.367
R1828 B.n544 B.n191 163.367
R1829 B.n548 B.n191 163.367
R1830 B.n548 B.n184 163.367
R1831 B.n556 B.n184 163.367
R1832 B.n556 B.n182 163.367
R1833 B.n560 B.n182 163.367
R1834 B.n560 B.n177 163.367
R1835 B.n568 B.n177 163.367
R1836 B.n568 B.n175 163.367
R1837 B.n572 B.n175 163.367
R1838 B.n572 B.n169 163.367
R1839 B.n580 B.n169 163.367
R1840 B.n580 B.n167 163.367
R1841 B.n584 B.n167 163.367
R1842 B.n584 B.n162 163.367
R1843 B.n593 B.n162 163.367
R1844 B.n593 B.n160 163.367
R1845 B.n597 B.n160 163.367
R1846 B.n597 B.n154 163.367
R1847 B.n605 B.n154 163.367
R1848 B.n605 B.n152 163.367
R1849 B.n609 B.n152 163.367
R1850 B.n609 B.n145 163.367
R1851 B.n617 B.n145 163.367
R1852 B.n617 B.n143 163.367
R1853 B.n622 B.n143 163.367
R1854 B.n622 B.n138 163.367
R1855 B.n630 B.n138 163.367
R1856 B.n631 B.n630 163.367
R1857 B.n631 B.n5 163.367
R1858 B.n6 B.n5 163.367
R1859 B.n7 B.n6 163.367
R1860 B.n636 B.n7 163.367
R1861 B.n636 B.n12 163.367
R1862 B.n13 B.n12 163.367
R1863 B.n14 B.n13 163.367
R1864 B.n641 B.n14 163.367
R1865 B.n641 B.n19 163.367
R1866 B.n20 B.n19 163.367
R1867 B.n21 B.n20 163.367
R1868 B.n646 B.n21 163.367
R1869 B.n646 B.n26 163.367
R1870 B.n27 B.n26 163.367
R1871 B.n28 B.n27 163.367
R1872 B.n651 B.n28 163.367
R1873 B.n651 B.n33 163.367
R1874 B.n34 B.n33 163.367
R1875 B.n35 B.n34 163.367
R1876 B.n656 B.n35 163.367
R1877 B.n656 B.n40 163.367
R1878 B.n41 B.n40 163.367
R1879 B.n42 B.n41 163.367
R1880 B.n661 B.n42 163.367
R1881 B.n661 B.n47 163.367
R1882 B.n48 B.n47 163.367
R1883 B.n49 B.n48 163.367
R1884 B.n666 B.n49 163.367
R1885 B.n666 B.n54 163.367
R1886 B.n55 B.n54 163.367
R1887 B.n56 B.n55 163.367
R1888 B.n671 B.n56 163.367
R1889 B.n671 B.n61 163.367
R1890 B.n62 B.n61 163.367
R1891 B.n63 B.n62 163.367
R1892 B.n676 B.n63 163.367
R1893 B.n676 B.n68 163.367
R1894 B.n69 B.n68 163.367
R1895 B.n70 B.n69 163.367
R1896 B.n921 B.n919 163.367
R1897 B.n917 B.n74 163.367
R1898 B.n913 B.n911 163.367
R1899 B.n909 B.n76 163.367
R1900 B.n905 B.n903 163.367
R1901 B.n901 B.n78 163.367
R1902 B.n897 B.n895 163.367
R1903 B.n893 B.n80 163.367
R1904 B.n889 B.n887 163.367
R1905 B.n885 B.n82 163.367
R1906 B.n881 B.n879 163.367
R1907 B.n877 B.n84 163.367
R1908 B.n873 B.n871 163.367
R1909 B.n869 B.n86 163.367
R1910 B.n865 B.n863 163.367
R1911 B.n861 B.n88 163.367
R1912 B.n857 B.n855 163.367
R1913 B.n853 B.n90 163.367
R1914 B.n849 B.n847 163.367
R1915 B.n845 B.n92 163.367
R1916 B.n841 B.n839 163.367
R1917 B.n837 B.n94 163.367
R1918 B.n833 B.n831 163.367
R1919 B.n829 B.n96 163.367
R1920 B.n825 B.n823 163.367
R1921 B.n821 B.n98 163.367
R1922 B.n817 B.n815 163.367
R1923 B.n813 B.n100 163.367
R1924 B.n808 B.n806 163.367
R1925 B.n804 B.n104 163.367
R1926 B.n800 B.n798 163.367
R1927 B.n796 B.n106 163.367
R1928 B.n791 B.n789 163.367
R1929 B.n787 B.n110 163.367
R1930 B.n783 B.n781 163.367
R1931 B.n779 B.n112 163.367
R1932 B.n775 B.n773 163.367
R1933 B.n771 B.n114 163.367
R1934 B.n767 B.n765 163.367
R1935 B.n763 B.n116 163.367
R1936 B.n759 B.n757 163.367
R1937 B.n755 B.n118 163.367
R1938 B.n751 B.n749 163.367
R1939 B.n747 B.n120 163.367
R1940 B.n743 B.n741 163.367
R1941 B.n739 B.n122 163.367
R1942 B.n735 B.n733 163.367
R1943 B.n731 B.n124 163.367
R1944 B.n727 B.n725 163.367
R1945 B.n723 B.n126 163.367
R1946 B.n719 B.n717 163.367
R1947 B.n715 B.n128 163.367
R1948 B.n711 B.n709 163.367
R1949 B.n707 B.n130 163.367
R1950 B.n703 B.n701 163.367
R1951 B.n699 B.n132 163.367
R1952 B.n695 B.n693 163.367
R1953 B.n691 B.n134 163.367
R1954 B.n687 B.n685 163.367
R1955 B.n683 B.n136 163.367
R1956 B.n513 B.n211 71.676
R1957 B.n511 B.n213 71.676
R1958 B.n507 B.n506 71.676
R1959 B.n500 B.n215 71.676
R1960 B.n499 B.n498 71.676
R1961 B.n492 B.n217 71.676
R1962 B.n491 B.n490 71.676
R1963 B.n484 B.n219 71.676
R1964 B.n483 B.n482 71.676
R1965 B.n476 B.n221 71.676
R1966 B.n475 B.n474 71.676
R1967 B.n468 B.n223 71.676
R1968 B.n467 B.n466 71.676
R1969 B.n460 B.n225 71.676
R1970 B.n459 B.n458 71.676
R1971 B.n452 B.n227 71.676
R1972 B.n451 B.n450 71.676
R1973 B.n444 B.n229 71.676
R1974 B.n443 B.n442 71.676
R1975 B.n436 B.n231 71.676
R1976 B.n435 B.n434 71.676
R1977 B.n428 B.n233 71.676
R1978 B.n427 B.n426 71.676
R1979 B.n420 B.n235 71.676
R1980 B.n419 B.n418 71.676
R1981 B.n412 B.n237 71.676
R1982 B.n411 B.n410 71.676
R1983 B.n403 B.n239 71.676
R1984 B.n402 B.n401 71.676
R1985 B.n395 B.n243 71.676
R1986 B.n394 B.n393 71.676
R1987 B.n387 B.n245 71.676
R1988 B.n386 B.n249 71.676
R1989 B.n382 B.n381 71.676
R1990 B.n375 B.n251 71.676
R1991 B.n374 B.n373 71.676
R1992 B.n367 B.n253 71.676
R1993 B.n366 B.n365 71.676
R1994 B.n359 B.n255 71.676
R1995 B.n358 B.n357 71.676
R1996 B.n351 B.n257 71.676
R1997 B.n350 B.n349 71.676
R1998 B.n343 B.n259 71.676
R1999 B.n342 B.n341 71.676
R2000 B.n335 B.n261 71.676
R2001 B.n334 B.n333 71.676
R2002 B.n327 B.n263 71.676
R2003 B.n326 B.n325 71.676
R2004 B.n319 B.n265 71.676
R2005 B.n318 B.n317 71.676
R2006 B.n311 B.n267 71.676
R2007 B.n310 B.n309 71.676
R2008 B.n303 B.n269 71.676
R2009 B.n302 B.n301 71.676
R2010 B.n295 B.n271 71.676
R2011 B.n294 B.n293 71.676
R2012 B.n287 B.n273 71.676
R2013 B.n286 B.n285 71.676
R2014 B.n279 B.n275 71.676
R2015 B.n278 B.n277 71.676
R2016 B.n920 B.n72 71.676
R2017 B.n919 B.n918 71.676
R2018 B.n912 B.n74 71.676
R2019 B.n911 B.n910 71.676
R2020 B.n904 B.n76 71.676
R2021 B.n903 B.n902 71.676
R2022 B.n896 B.n78 71.676
R2023 B.n895 B.n894 71.676
R2024 B.n888 B.n80 71.676
R2025 B.n887 B.n886 71.676
R2026 B.n880 B.n82 71.676
R2027 B.n879 B.n878 71.676
R2028 B.n872 B.n84 71.676
R2029 B.n871 B.n870 71.676
R2030 B.n864 B.n86 71.676
R2031 B.n863 B.n862 71.676
R2032 B.n856 B.n88 71.676
R2033 B.n855 B.n854 71.676
R2034 B.n848 B.n90 71.676
R2035 B.n847 B.n846 71.676
R2036 B.n840 B.n92 71.676
R2037 B.n839 B.n838 71.676
R2038 B.n832 B.n94 71.676
R2039 B.n831 B.n830 71.676
R2040 B.n824 B.n96 71.676
R2041 B.n823 B.n822 71.676
R2042 B.n816 B.n98 71.676
R2043 B.n815 B.n814 71.676
R2044 B.n807 B.n100 71.676
R2045 B.n806 B.n805 71.676
R2046 B.n799 B.n104 71.676
R2047 B.n798 B.n797 71.676
R2048 B.n790 B.n106 71.676
R2049 B.n789 B.n788 71.676
R2050 B.n782 B.n110 71.676
R2051 B.n781 B.n780 71.676
R2052 B.n774 B.n112 71.676
R2053 B.n773 B.n772 71.676
R2054 B.n766 B.n114 71.676
R2055 B.n765 B.n764 71.676
R2056 B.n758 B.n116 71.676
R2057 B.n757 B.n756 71.676
R2058 B.n750 B.n118 71.676
R2059 B.n749 B.n748 71.676
R2060 B.n742 B.n120 71.676
R2061 B.n741 B.n740 71.676
R2062 B.n734 B.n122 71.676
R2063 B.n733 B.n732 71.676
R2064 B.n726 B.n124 71.676
R2065 B.n725 B.n724 71.676
R2066 B.n718 B.n126 71.676
R2067 B.n717 B.n716 71.676
R2068 B.n710 B.n128 71.676
R2069 B.n709 B.n708 71.676
R2070 B.n702 B.n130 71.676
R2071 B.n701 B.n700 71.676
R2072 B.n694 B.n132 71.676
R2073 B.n693 B.n692 71.676
R2074 B.n686 B.n134 71.676
R2075 B.n685 B.n684 71.676
R2076 B.n684 B.n683 71.676
R2077 B.n687 B.n686 71.676
R2078 B.n692 B.n691 71.676
R2079 B.n695 B.n694 71.676
R2080 B.n700 B.n699 71.676
R2081 B.n703 B.n702 71.676
R2082 B.n708 B.n707 71.676
R2083 B.n711 B.n710 71.676
R2084 B.n716 B.n715 71.676
R2085 B.n719 B.n718 71.676
R2086 B.n724 B.n723 71.676
R2087 B.n727 B.n726 71.676
R2088 B.n732 B.n731 71.676
R2089 B.n735 B.n734 71.676
R2090 B.n740 B.n739 71.676
R2091 B.n743 B.n742 71.676
R2092 B.n748 B.n747 71.676
R2093 B.n751 B.n750 71.676
R2094 B.n756 B.n755 71.676
R2095 B.n759 B.n758 71.676
R2096 B.n764 B.n763 71.676
R2097 B.n767 B.n766 71.676
R2098 B.n772 B.n771 71.676
R2099 B.n775 B.n774 71.676
R2100 B.n780 B.n779 71.676
R2101 B.n783 B.n782 71.676
R2102 B.n788 B.n787 71.676
R2103 B.n791 B.n790 71.676
R2104 B.n797 B.n796 71.676
R2105 B.n800 B.n799 71.676
R2106 B.n805 B.n804 71.676
R2107 B.n808 B.n807 71.676
R2108 B.n814 B.n813 71.676
R2109 B.n817 B.n816 71.676
R2110 B.n822 B.n821 71.676
R2111 B.n825 B.n824 71.676
R2112 B.n830 B.n829 71.676
R2113 B.n833 B.n832 71.676
R2114 B.n838 B.n837 71.676
R2115 B.n841 B.n840 71.676
R2116 B.n846 B.n845 71.676
R2117 B.n849 B.n848 71.676
R2118 B.n854 B.n853 71.676
R2119 B.n857 B.n856 71.676
R2120 B.n862 B.n861 71.676
R2121 B.n865 B.n864 71.676
R2122 B.n870 B.n869 71.676
R2123 B.n873 B.n872 71.676
R2124 B.n878 B.n877 71.676
R2125 B.n881 B.n880 71.676
R2126 B.n886 B.n885 71.676
R2127 B.n889 B.n888 71.676
R2128 B.n894 B.n893 71.676
R2129 B.n897 B.n896 71.676
R2130 B.n902 B.n901 71.676
R2131 B.n905 B.n904 71.676
R2132 B.n910 B.n909 71.676
R2133 B.n913 B.n912 71.676
R2134 B.n918 B.n917 71.676
R2135 B.n921 B.n920 71.676
R2136 B.n514 B.n513 71.676
R2137 B.n508 B.n213 71.676
R2138 B.n506 B.n505 71.676
R2139 B.n501 B.n500 71.676
R2140 B.n498 B.n497 71.676
R2141 B.n493 B.n492 71.676
R2142 B.n490 B.n489 71.676
R2143 B.n485 B.n484 71.676
R2144 B.n482 B.n481 71.676
R2145 B.n477 B.n476 71.676
R2146 B.n474 B.n473 71.676
R2147 B.n469 B.n468 71.676
R2148 B.n466 B.n465 71.676
R2149 B.n461 B.n460 71.676
R2150 B.n458 B.n457 71.676
R2151 B.n453 B.n452 71.676
R2152 B.n450 B.n449 71.676
R2153 B.n445 B.n444 71.676
R2154 B.n442 B.n441 71.676
R2155 B.n437 B.n436 71.676
R2156 B.n434 B.n433 71.676
R2157 B.n429 B.n428 71.676
R2158 B.n426 B.n425 71.676
R2159 B.n421 B.n420 71.676
R2160 B.n418 B.n417 71.676
R2161 B.n413 B.n412 71.676
R2162 B.n410 B.n409 71.676
R2163 B.n404 B.n403 71.676
R2164 B.n401 B.n400 71.676
R2165 B.n396 B.n395 71.676
R2166 B.n393 B.n392 71.676
R2167 B.n388 B.n387 71.676
R2168 B.n383 B.n249 71.676
R2169 B.n381 B.n380 71.676
R2170 B.n376 B.n375 71.676
R2171 B.n373 B.n372 71.676
R2172 B.n368 B.n367 71.676
R2173 B.n365 B.n364 71.676
R2174 B.n360 B.n359 71.676
R2175 B.n357 B.n356 71.676
R2176 B.n352 B.n351 71.676
R2177 B.n349 B.n348 71.676
R2178 B.n344 B.n343 71.676
R2179 B.n341 B.n340 71.676
R2180 B.n336 B.n335 71.676
R2181 B.n333 B.n332 71.676
R2182 B.n328 B.n327 71.676
R2183 B.n325 B.n324 71.676
R2184 B.n320 B.n319 71.676
R2185 B.n317 B.n316 71.676
R2186 B.n312 B.n311 71.676
R2187 B.n309 B.n308 71.676
R2188 B.n304 B.n303 71.676
R2189 B.n301 B.n300 71.676
R2190 B.n296 B.n295 71.676
R2191 B.n293 B.n292 71.676
R2192 B.n288 B.n287 71.676
R2193 B.n285 B.n284 71.676
R2194 B.n280 B.n279 71.676
R2195 B.n277 B.n209 71.676
R2196 B.n519 B.n210 71.1609
R2197 B.n926 B.n71 71.1609
R2198 B.n248 B.n247 59.5399
R2199 B.n406 B.n241 59.5399
R2200 B.n811 B.n102 59.5399
R2201 B.n793 B.n108 59.5399
R2202 B.n681 B.n680 36.6834
R2203 B.n924 B.n923 36.6834
R2204 B.n521 B.n208 36.6834
R2205 B.n517 B.n516 36.6834
R2206 B.n519 B.n206 33.839
R2207 B.n525 B.n206 33.839
R2208 B.n525 B.n201 33.839
R2209 B.n531 B.n201 33.839
R2210 B.n531 B.n202 33.839
R2211 B.n537 B.n194 33.839
R2212 B.n543 B.n194 33.839
R2213 B.n543 B.n190 33.839
R2214 B.n549 B.n190 33.839
R2215 B.n549 B.n185 33.839
R2216 B.n555 B.n185 33.839
R2217 B.n555 B.n186 33.839
R2218 B.n561 B.n178 33.839
R2219 B.n567 B.n178 33.839
R2220 B.n567 B.n174 33.839
R2221 B.n573 B.n174 33.839
R2222 B.n579 B.n170 33.839
R2223 B.n579 B.n166 33.839
R2224 B.n586 B.n166 33.839
R2225 B.n586 B.n585 33.839
R2226 B.n592 B.n159 33.839
R2227 B.n598 B.n159 33.839
R2228 B.n598 B.n155 33.839
R2229 B.n604 B.n155 33.839
R2230 B.n610 B.n151 33.839
R2231 B.n610 B.n146 33.839
R2232 B.n616 B.n146 33.839
R2233 B.n616 B.n147 33.839
R2234 B.n623 B.n139 33.839
R2235 B.n629 B.n139 33.839
R2236 B.n629 B.n4 33.839
R2237 B.n1000 B.n4 33.839
R2238 B.n1000 B.n999 33.839
R2239 B.n999 B.n998 33.839
R2240 B.n998 B.n8 33.839
R2241 B.n992 B.n8 33.839
R2242 B.n991 B.n990 33.839
R2243 B.n990 B.n15 33.839
R2244 B.n984 B.n15 33.839
R2245 B.n984 B.n983 33.839
R2246 B.n982 B.n22 33.839
R2247 B.n976 B.n22 33.839
R2248 B.n976 B.n975 33.839
R2249 B.n975 B.n974 33.839
R2250 B.n968 B.n32 33.839
R2251 B.n968 B.n967 33.839
R2252 B.n967 B.n966 33.839
R2253 B.n966 B.n36 33.839
R2254 B.n960 B.n959 33.839
R2255 B.n959 B.n958 33.839
R2256 B.n958 B.n43 33.839
R2257 B.n952 B.n43 33.839
R2258 B.n951 B.n950 33.839
R2259 B.n950 B.n50 33.839
R2260 B.n944 B.n50 33.839
R2261 B.n944 B.n943 33.839
R2262 B.n943 B.n942 33.839
R2263 B.n942 B.n57 33.839
R2264 B.n936 B.n57 33.839
R2265 B.n935 B.n934 33.839
R2266 B.n934 B.n64 33.839
R2267 B.n928 B.n64 33.839
R2268 B.n928 B.n927 33.839
R2269 B.n927 B.n926 33.839
R2270 B.n247 B.n246 33.1641
R2271 B.n241 B.n240 33.1641
R2272 B.n102 B.n101 33.1641
R2273 B.n108 B.n107 33.1641
R2274 B.n147 B.t5 29.858
R2275 B.t1 B.n991 29.858
R2276 B.n604 B.t4 28.8627
R2277 B.t6 B.n982 28.8627
R2278 B.n585 B.t7 27.8675
R2279 B.n32 B.t8 27.8675
R2280 B.n573 B.t3 26.8722
R2281 B.n960 B.t0 26.8722
R2282 B.n186 B.t2 25.877
R2283 B.t9 B.n951 25.877
R2284 B B.n1002 18.0485
R2285 B.n202 B.t11 17.915
R2286 B.t15 B.n935 17.915
R2287 B.n537 B.t11 15.9245
R2288 B.n936 B.t15 15.9245
R2289 B.n923 B.n922 10.6151
R2290 B.n922 B.n73 10.6151
R2291 B.n916 B.n73 10.6151
R2292 B.n916 B.n915 10.6151
R2293 B.n915 B.n914 10.6151
R2294 B.n914 B.n75 10.6151
R2295 B.n908 B.n75 10.6151
R2296 B.n908 B.n907 10.6151
R2297 B.n907 B.n906 10.6151
R2298 B.n906 B.n77 10.6151
R2299 B.n900 B.n77 10.6151
R2300 B.n900 B.n899 10.6151
R2301 B.n899 B.n898 10.6151
R2302 B.n898 B.n79 10.6151
R2303 B.n892 B.n79 10.6151
R2304 B.n892 B.n891 10.6151
R2305 B.n891 B.n890 10.6151
R2306 B.n890 B.n81 10.6151
R2307 B.n884 B.n81 10.6151
R2308 B.n884 B.n883 10.6151
R2309 B.n883 B.n882 10.6151
R2310 B.n882 B.n83 10.6151
R2311 B.n876 B.n83 10.6151
R2312 B.n876 B.n875 10.6151
R2313 B.n875 B.n874 10.6151
R2314 B.n874 B.n85 10.6151
R2315 B.n868 B.n85 10.6151
R2316 B.n868 B.n867 10.6151
R2317 B.n867 B.n866 10.6151
R2318 B.n866 B.n87 10.6151
R2319 B.n860 B.n87 10.6151
R2320 B.n860 B.n859 10.6151
R2321 B.n859 B.n858 10.6151
R2322 B.n858 B.n89 10.6151
R2323 B.n852 B.n89 10.6151
R2324 B.n852 B.n851 10.6151
R2325 B.n851 B.n850 10.6151
R2326 B.n850 B.n91 10.6151
R2327 B.n844 B.n91 10.6151
R2328 B.n844 B.n843 10.6151
R2329 B.n843 B.n842 10.6151
R2330 B.n842 B.n93 10.6151
R2331 B.n836 B.n93 10.6151
R2332 B.n836 B.n835 10.6151
R2333 B.n835 B.n834 10.6151
R2334 B.n834 B.n95 10.6151
R2335 B.n828 B.n95 10.6151
R2336 B.n828 B.n827 10.6151
R2337 B.n827 B.n826 10.6151
R2338 B.n826 B.n97 10.6151
R2339 B.n820 B.n97 10.6151
R2340 B.n820 B.n819 10.6151
R2341 B.n819 B.n818 10.6151
R2342 B.n818 B.n99 10.6151
R2343 B.n812 B.n99 10.6151
R2344 B.n810 B.n809 10.6151
R2345 B.n809 B.n103 10.6151
R2346 B.n803 B.n103 10.6151
R2347 B.n803 B.n802 10.6151
R2348 B.n802 B.n801 10.6151
R2349 B.n801 B.n105 10.6151
R2350 B.n795 B.n105 10.6151
R2351 B.n795 B.n794 10.6151
R2352 B.n792 B.n109 10.6151
R2353 B.n786 B.n109 10.6151
R2354 B.n786 B.n785 10.6151
R2355 B.n785 B.n784 10.6151
R2356 B.n784 B.n111 10.6151
R2357 B.n778 B.n111 10.6151
R2358 B.n778 B.n777 10.6151
R2359 B.n777 B.n776 10.6151
R2360 B.n776 B.n113 10.6151
R2361 B.n770 B.n113 10.6151
R2362 B.n770 B.n769 10.6151
R2363 B.n769 B.n768 10.6151
R2364 B.n768 B.n115 10.6151
R2365 B.n762 B.n115 10.6151
R2366 B.n762 B.n761 10.6151
R2367 B.n761 B.n760 10.6151
R2368 B.n760 B.n117 10.6151
R2369 B.n754 B.n117 10.6151
R2370 B.n754 B.n753 10.6151
R2371 B.n753 B.n752 10.6151
R2372 B.n752 B.n119 10.6151
R2373 B.n746 B.n119 10.6151
R2374 B.n746 B.n745 10.6151
R2375 B.n745 B.n744 10.6151
R2376 B.n744 B.n121 10.6151
R2377 B.n738 B.n121 10.6151
R2378 B.n738 B.n737 10.6151
R2379 B.n737 B.n736 10.6151
R2380 B.n736 B.n123 10.6151
R2381 B.n730 B.n123 10.6151
R2382 B.n730 B.n729 10.6151
R2383 B.n729 B.n728 10.6151
R2384 B.n728 B.n125 10.6151
R2385 B.n722 B.n125 10.6151
R2386 B.n722 B.n721 10.6151
R2387 B.n721 B.n720 10.6151
R2388 B.n720 B.n127 10.6151
R2389 B.n714 B.n127 10.6151
R2390 B.n714 B.n713 10.6151
R2391 B.n713 B.n712 10.6151
R2392 B.n712 B.n129 10.6151
R2393 B.n706 B.n129 10.6151
R2394 B.n706 B.n705 10.6151
R2395 B.n705 B.n704 10.6151
R2396 B.n704 B.n131 10.6151
R2397 B.n698 B.n131 10.6151
R2398 B.n698 B.n697 10.6151
R2399 B.n697 B.n696 10.6151
R2400 B.n696 B.n133 10.6151
R2401 B.n690 B.n133 10.6151
R2402 B.n690 B.n689 10.6151
R2403 B.n689 B.n688 10.6151
R2404 B.n688 B.n135 10.6151
R2405 B.n682 B.n135 10.6151
R2406 B.n682 B.n681 10.6151
R2407 B.n522 B.n521 10.6151
R2408 B.n523 B.n522 10.6151
R2409 B.n523 B.n199 10.6151
R2410 B.n533 B.n199 10.6151
R2411 B.n534 B.n533 10.6151
R2412 B.n535 B.n534 10.6151
R2413 B.n535 B.n192 10.6151
R2414 B.n545 B.n192 10.6151
R2415 B.n546 B.n545 10.6151
R2416 B.n547 B.n546 10.6151
R2417 B.n547 B.n183 10.6151
R2418 B.n557 B.n183 10.6151
R2419 B.n558 B.n557 10.6151
R2420 B.n559 B.n558 10.6151
R2421 B.n559 B.n176 10.6151
R2422 B.n569 B.n176 10.6151
R2423 B.n570 B.n569 10.6151
R2424 B.n571 B.n570 10.6151
R2425 B.n571 B.n168 10.6151
R2426 B.n581 B.n168 10.6151
R2427 B.n582 B.n581 10.6151
R2428 B.n583 B.n582 10.6151
R2429 B.n583 B.n161 10.6151
R2430 B.n594 B.n161 10.6151
R2431 B.n595 B.n594 10.6151
R2432 B.n596 B.n595 10.6151
R2433 B.n596 B.n153 10.6151
R2434 B.n606 B.n153 10.6151
R2435 B.n607 B.n606 10.6151
R2436 B.n608 B.n607 10.6151
R2437 B.n608 B.n144 10.6151
R2438 B.n618 B.n144 10.6151
R2439 B.n619 B.n618 10.6151
R2440 B.n621 B.n619 10.6151
R2441 B.n621 B.n620 10.6151
R2442 B.n620 B.n137 10.6151
R2443 B.n632 B.n137 10.6151
R2444 B.n633 B.n632 10.6151
R2445 B.n634 B.n633 10.6151
R2446 B.n635 B.n634 10.6151
R2447 B.n637 B.n635 10.6151
R2448 B.n638 B.n637 10.6151
R2449 B.n639 B.n638 10.6151
R2450 B.n640 B.n639 10.6151
R2451 B.n642 B.n640 10.6151
R2452 B.n643 B.n642 10.6151
R2453 B.n644 B.n643 10.6151
R2454 B.n645 B.n644 10.6151
R2455 B.n647 B.n645 10.6151
R2456 B.n648 B.n647 10.6151
R2457 B.n649 B.n648 10.6151
R2458 B.n650 B.n649 10.6151
R2459 B.n652 B.n650 10.6151
R2460 B.n653 B.n652 10.6151
R2461 B.n654 B.n653 10.6151
R2462 B.n655 B.n654 10.6151
R2463 B.n657 B.n655 10.6151
R2464 B.n658 B.n657 10.6151
R2465 B.n659 B.n658 10.6151
R2466 B.n660 B.n659 10.6151
R2467 B.n662 B.n660 10.6151
R2468 B.n663 B.n662 10.6151
R2469 B.n664 B.n663 10.6151
R2470 B.n665 B.n664 10.6151
R2471 B.n667 B.n665 10.6151
R2472 B.n668 B.n667 10.6151
R2473 B.n669 B.n668 10.6151
R2474 B.n670 B.n669 10.6151
R2475 B.n672 B.n670 10.6151
R2476 B.n673 B.n672 10.6151
R2477 B.n674 B.n673 10.6151
R2478 B.n675 B.n674 10.6151
R2479 B.n677 B.n675 10.6151
R2480 B.n678 B.n677 10.6151
R2481 B.n679 B.n678 10.6151
R2482 B.n680 B.n679 10.6151
R2483 B.n516 B.n515 10.6151
R2484 B.n515 B.n212 10.6151
R2485 B.n510 B.n212 10.6151
R2486 B.n510 B.n509 10.6151
R2487 B.n509 B.n214 10.6151
R2488 B.n504 B.n214 10.6151
R2489 B.n504 B.n503 10.6151
R2490 B.n503 B.n502 10.6151
R2491 B.n502 B.n216 10.6151
R2492 B.n496 B.n216 10.6151
R2493 B.n496 B.n495 10.6151
R2494 B.n495 B.n494 10.6151
R2495 B.n494 B.n218 10.6151
R2496 B.n488 B.n218 10.6151
R2497 B.n488 B.n487 10.6151
R2498 B.n487 B.n486 10.6151
R2499 B.n486 B.n220 10.6151
R2500 B.n480 B.n220 10.6151
R2501 B.n480 B.n479 10.6151
R2502 B.n479 B.n478 10.6151
R2503 B.n478 B.n222 10.6151
R2504 B.n472 B.n222 10.6151
R2505 B.n472 B.n471 10.6151
R2506 B.n471 B.n470 10.6151
R2507 B.n470 B.n224 10.6151
R2508 B.n464 B.n224 10.6151
R2509 B.n464 B.n463 10.6151
R2510 B.n463 B.n462 10.6151
R2511 B.n462 B.n226 10.6151
R2512 B.n456 B.n226 10.6151
R2513 B.n456 B.n455 10.6151
R2514 B.n455 B.n454 10.6151
R2515 B.n454 B.n228 10.6151
R2516 B.n448 B.n228 10.6151
R2517 B.n448 B.n447 10.6151
R2518 B.n447 B.n446 10.6151
R2519 B.n446 B.n230 10.6151
R2520 B.n440 B.n230 10.6151
R2521 B.n440 B.n439 10.6151
R2522 B.n439 B.n438 10.6151
R2523 B.n438 B.n232 10.6151
R2524 B.n432 B.n232 10.6151
R2525 B.n432 B.n431 10.6151
R2526 B.n431 B.n430 10.6151
R2527 B.n430 B.n234 10.6151
R2528 B.n424 B.n234 10.6151
R2529 B.n424 B.n423 10.6151
R2530 B.n423 B.n422 10.6151
R2531 B.n422 B.n236 10.6151
R2532 B.n416 B.n236 10.6151
R2533 B.n416 B.n415 10.6151
R2534 B.n415 B.n414 10.6151
R2535 B.n414 B.n238 10.6151
R2536 B.n408 B.n238 10.6151
R2537 B.n408 B.n407 10.6151
R2538 B.n405 B.n242 10.6151
R2539 B.n399 B.n242 10.6151
R2540 B.n399 B.n398 10.6151
R2541 B.n398 B.n397 10.6151
R2542 B.n397 B.n244 10.6151
R2543 B.n391 B.n244 10.6151
R2544 B.n391 B.n390 10.6151
R2545 B.n390 B.n389 10.6151
R2546 B.n385 B.n384 10.6151
R2547 B.n384 B.n250 10.6151
R2548 B.n379 B.n250 10.6151
R2549 B.n379 B.n378 10.6151
R2550 B.n378 B.n377 10.6151
R2551 B.n377 B.n252 10.6151
R2552 B.n371 B.n252 10.6151
R2553 B.n371 B.n370 10.6151
R2554 B.n370 B.n369 10.6151
R2555 B.n369 B.n254 10.6151
R2556 B.n363 B.n254 10.6151
R2557 B.n363 B.n362 10.6151
R2558 B.n362 B.n361 10.6151
R2559 B.n361 B.n256 10.6151
R2560 B.n355 B.n256 10.6151
R2561 B.n355 B.n354 10.6151
R2562 B.n354 B.n353 10.6151
R2563 B.n353 B.n258 10.6151
R2564 B.n347 B.n258 10.6151
R2565 B.n347 B.n346 10.6151
R2566 B.n346 B.n345 10.6151
R2567 B.n345 B.n260 10.6151
R2568 B.n339 B.n260 10.6151
R2569 B.n339 B.n338 10.6151
R2570 B.n338 B.n337 10.6151
R2571 B.n337 B.n262 10.6151
R2572 B.n331 B.n262 10.6151
R2573 B.n331 B.n330 10.6151
R2574 B.n330 B.n329 10.6151
R2575 B.n329 B.n264 10.6151
R2576 B.n323 B.n264 10.6151
R2577 B.n323 B.n322 10.6151
R2578 B.n322 B.n321 10.6151
R2579 B.n321 B.n266 10.6151
R2580 B.n315 B.n266 10.6151
R2581 B.n315 B.n314 10.6151
R2582 B.n314 B.n313 10.6151
R2583 B.n313 B.n268 10.6151
R2584 B.n307 B.n268 10.6151
R2585 B.n307 B.n306 10.6151
R2586 B.n306 B.n305 10.6151
R2587 B.n305 B.n270 10.6151
R2588 B.n299 B.n270 10.6151
R2589 B.n299 B.n298 10.6151
R2590 B.n298 B.n297 10.6151
R2591 B.n297 B.n272 10.6151
R2592 B.n291 B.n272 10.6151
R2593 B.n291 B.n290 10.6151
R2594 B.n290 B.n289 10.6151
R2595 B.n289 B.n274 10.6151
R2596 B.n283 B.n274 10.6151
R2597 B.n283 B.n282 10.6151
R2598 B.n282 B.n281 10.6151
R2599 B.n281 B.n276 10.6151
R2600 B.n276 B.n208 10.6151
R2601 B.n517 B.n204 10.6151
R2602 B.n527 B.n204 10.6151
R2603 B.n528 B.n527 10.6151
R2604 B.n529 B.n528 10.6151
R2605 B.n529 B.n196 10.6151
R2606 B.n539 B.n196 10.6151
R2607 B.n540 B.n539 10.6151
R2608 B.n541 B.n540 10.6151
R2609 B.n541 B.n188 10.6151
R2610 B.n551 B.n188 10.6151
R2611 B.n552 B.n551 10.6151
R2612 B.n553 B.n552 10.6151
R2613 B.n553 B.n180 10.6151
R2614 B.n563 B.n180 10.6151
R2615 B.n564 B.n563 10.6151
R2616 B.n565 B.n564 10.6151
R2617 B.n565 B.n172 10.6151
R2618 B.n575 B.n172 10.6151
R2619 B.n576 B.n575 10.6151
R2620 B.n577 B.n576 10.6151
R2621 B.n577 B.n164 10.6151
R2622 B.n588 B.n164 10.6151
R2623 B.n589 B.n588 10.6151
R2624 B.n590 B.n589 10.6151
R2625 B.n590 B.n157 10.6151
R2626 B.n600 B.n157 10.6151
R2627 B.n601 B.n600 10.6151
R2628 B.n602 B.n601 10.6151
R2629 B.n602 B.n149 10.6151
R2630 B.n612 B.n149 10.6151
R2631 B.n613 B.n612 10.6151
R2632 B.n614 B.n613 10.6151
R2633 B.n614 B.n141 10.6151
R2634 B.n625 B.n141 10.6151
R2635 B.n626 B.n625 10.6151
R2636 B.n627 B.n626 10.6151
R2637 B.n627 B.n0 10.6151
R2638 B.n996 B.n1 10.6151
R2639 B.n996 B.n995 10.6151
R2640 B.n995 B.n994 10.6151
R2641 B.n994 B.n10 10.6151
R2642 B.n988 B.n10 10.6151
R2643 B.n988 B.n987 10.6151
R2644 B.n987 B.n986 10.6151
R2645 B.n986 B.n17 10.6151
R2646 B.n980 B.n17 10.6151
R2647 B.n980 B.n979 10.6151
R2648 B.n979 B.n978 10.6151
R2649 B.n978 B.n24 10.6151
R2650 B.n972 B.n24 10.6151
R2651 B.n972 B.n971 10.6151
R2652 B.n971 B.n970 10.6151
R2653 B.n970 B.n30 10.6151
R2654 B.n964 B.n30 10.6151
R2655 B.n964 B.n963 10.6151
R2656 B.n963 B.n962 10.6151
R2657 B.n962 B.n38 10.6151
R2658 B.n956 B.n38 10.6151
R2659 B.n956 B.n955 10.6151
R2660 B.n955 B.n954 10.6151
R2661 B.n954 B.n45 10.6151
R2662 B.n948 B.n45 10.6151
R2663 B.n948 B.n947 10.6151
R2664 B.n947 B.n946 10.6151
R2665 B.n946 B.n52 10.6151
R2666 B.n940 B.n52 10.6151
R2667 B.n940 B.n939 10.6151
R2668 B.n939 B.n938 10.6151
R2669 B.n938 B.n59 10.6151
R2670 B.n932 B.n59 10.6151
R2671 B.n932 B.n931 10.6151
R2672 B.n931 B.n930 10.6151
R2673 B.n930 B.n66 10.6151
R2674 B.n924 B.n66 10.6151
R2675 B.n561 B.t2 7.9625
R2676 B.n952 B.t9 7.9625
R2677 B.t3 B.n170 6.96725
R2678 B.t0 B.n36 6.96725
R2679 B.n811 B.n810 6.5566
R2680 B.n794 B.n793 6.5566
R2681 B.n406 B.n405 6.5566
R2682 B.n389 B.n248 6.5566
R2683 B.n592 B.t7 5.972
R2684 B.n974 B.t8 5.972
R2685 B.t4 B.n151 4.97675
R2686 B.n983 B.t6 4.97675
R2687 B.n812 B.n811 4.05904
R2688 B.n793 B.n792 4.05904
R2689 B.n407 B.n406 4.05904
R2690 B.n385 B.n248 4.05904
R2691 B.n623 B.t5 3.9815
R2692 B.n992 B.t1 3.9815
R2693 B.n1002 B.n0 2.81026
R2694 B.n1002 B.n1 2.81026
R2695 VN.n6 VN.t3 326.76
R2696 VN.n33 VN.t5 326.76
R2697 VN.n5 VN.t4 293.916
R2698 VN.n10 VN.t6 293.916
R2699 VN.n17 VN.t8 293.916
R2700 VN.n24 VN.t0 293.916
R2701 VN.n32 VN.t1 293.916
R2702 VN.n31 VN.t7 293.916
R2703 VN.n43 VN.t2 293.916
R2704 VN.n50 VN.t9 293.916
R2705 VN.n25 VN.n24 177.448
R2706 VN.n51 VN.n50 177.448
R2707 VN.n49 VN.n26 161.3
R2708 VN.n48 VN.n47 161.3
R2709 VN.n46 VN.n27 161.3
R2710 VN.n45 VN.n44 161.3
R2711 VN.n42 VN.n28 161.3
R2712 VN.n41 VN.n40 161.3
R2713 VN.n39 VN.n29 161.3
R2714 VN.n38 VN.n37 161.3
R2715 VN.n36 VN.n30 161.3
R2716 VN.n35 VN.n34 161.3
R2717 VN.n23 VN.n0 161.3
R2718 VN.n22 VN.n21 161.3
R2719 VN.n20 VN.n1 161.3
R2720 VN.n19 VN.n18 161.3
R2721 VN.n16 VN.n2 161.3
R2722 VN.n15 VN.n14 161.3
R2723 VN.n13 VN.n3 161.3
R2724 VN.n12 VN.n11 161.3
R2725 VN.n9 VN.n4 161.3
R2726 VN.n8 VN.n7 161.3
R2727 VN.n22 VN.n1 56.5193
R2728 VN.n48 VN.n27 56.5193
R2729 VN.n9 VN.n8 50.6917
R2730 VN.n16 VN.n15 50.6917
R2731 VN.n36 VN.n35 50.6917
R2732 VN.n42 VN.n41 50.6917
R2733 VN VN.n51 50.3925
R2734 VN.n6 VN.n5 43.6963
R2735 VN.n33 VN.n32 43.6963
R2736 VN.n11 VN.n9 30.2951
R2737 VN.n15 VN.n3 30.2951
R2738 VN.n37 VN.n36 30.2951
R2739 VN.n41 VN.n29 30.2951
R2740 VN.n18 VN.n1 24.4675
R2741 VN.n23 VN.n22 24.4675
R2742 VN.n44 VN.n27 24.4675
R2743 VN.n49 VN.n48 24.4675
R2744 VN.n8 VN.n5 22.5101
R2745 VN.n17 VN.n16 22.5101
R2746 VN.n35 VN.n32 22.5101
R2747 VN.n43 VN.n42 22.5101
R2748 VN.n34 VN.n33 17.9509
R2749 VN.n7 VN.n6 17.9509
R2750 VN.n11 VN.n10 12.234
R2751 VN.n10 VN.n3 12.234
R2752 VN.n31 VN.n29 12.234
R2753 VN.n37 VN.n31 12.234
R2754 VN.n24 VN.n23 8.31928
R2755 VN.n50 VN.n49 8.31928
R2756 VN.n18 VN.n17 1.95786
R2757 VN.n44 VN.n43 1.95786
R2758 VN.n51 VN.n26 0.189894
R2759 VN.n47 VN.n26 0.189894
R2760 VN.n47 VN.n46 0.189894
R2761 VN.n46 VN.n45 0.189894
R2762 VN.n45 VN.n28 0.189894
R2763 VN.n40 VN.n28 0.189894
R2764 VN.n40 VN.n39 0.189894
R2765 VN.n39 VN.n38 0.189894
R2766 VN.n38 VN.n30 0.189894
R2767 VN.n34 VN.n30 0.189894
R2768 VN.n7 VN.n4 0.189894
R2769 VN.n12 VN.n4 0.189894
R2770 VN.n13 VN.n12 0.189894
R2771 VN.n14 VN.n13 0.189894
R2772 VN.n14 VN.n2 0.189894
R2773 VN.n19 VN.n2 0.189894
R2774 VN.n20 VN.n19 0.189894
R2775 VN.n21 VN.n20 0.189894
R2776 VN.n21 VN.n0 0.189894
R2777 VN.n25 VN.n0 0.189894
R2778 VN VN.n25 0.0516364
R2779 VDD2.n185 VDD2.n97 289.615
R2780 VDD2.n88 VDD2.n0 289.615
R2781 VDD2.n186 VDD2.n185 185
R2782 VDD2.n184 VDD2.n183 185
R2783 VDD2.n101 VDD2.n100 185
R2784 VDD2.n178 VDD2.n177 185
R2785 VDD2.n176 VDD2.n175 185
R2786 VDD2.n174 VDD2.n104 185
R2787 VDD2.n108 VDD2.n105 185
R2788 VDD2.n169 VDD2.n168 185
R2789 VDD2.n167 VDD2.n166 185
R2790 VDD2.n110 VDD2.n109 185
R2791 VDD2.n161 VDD2.n160 185
R2792 VDD2.n159 VDD2.n158 185
R2793 VDD2.n114 VDD2.n113 185
R2794 VDD2.n153 VDD2.n152 185
R2795 VDD2.n151 VDD2.n150 185
R2796 VDD2.n118 VDD2.n117 185
R2797 VDD2.n145 VDD2.n144 185
R2798 VDD2.n143 VDD2.n142 185
R2799 VDD2.n122 VDD2.n121 185
R2800 VDD2.n137 VDD2.n136 185
R2801 VDD2.n135 VDD2.n134 185
R2802 VDD2.n126 VDD2.n125 185
R2803 VDD2.n129 VDD2.n128 185
R2804 VDD2.n31 VDD2.n30 185
R2805 VDD2.n28 VDD2.n27 185
R2806 VDD2.n37 VDD2.n36 185
R2807 VDD2.n39 VDD2.n38 185
R2808 VDD2.n24 VDD2.n23 185
R2809 VDD2.n45 VDD2.n44 185
R2810 VDD2.n47 VDD2.n46 185
R2811 VDD2.n20 VDD2.n19 185
R2812 VDD2.n53 VDD2.n52 185
R2813 VDD2.n55 VDD2.n54 185
R2814 VDD2.n16 VDD2.n15 185
R2815 VDD2.n61 VDD2.n60 185
R2816 VDD2.n63 VDD2.n62 185
R2817 VDD2.n12 VDD2.n11 185
R2818 VDD2.n69 VDD2.n68 185
R2819 VDD2.n72 VDD2.n71 185
R2820 VDD2.n70 VDD2.n8 185
R2821 VDD2.n77 VDD2.n7 185
R2822 VDD2.n79 VDD2.n78 185
R2823 VDD2.n81 VDD2.n80 185
R2824 VDD2.n4 VDD2.n3 185
R2825 VDD2.n87 VDD2.n86 185
R2826 VDD2.n89 VDD2.n88 185
R2827 VDD2.t0 VDD2.n127 147.659
R2828 VDD2.t6 VDD2.n29 147.659
R2829 VDD2.n185 VDD2.n184 104.615
R2830 VDD2.n184 VDD2.n100 104.615
R2831 VDD2.n177 VDD2.n100 104.615
R2832 VDD2.n177 VDD2.n176 104.615
R2833 VDD2.n176 VDD2.n104 104.615
R2834 VDD2.n108 VDD2.n104 104.615
R2835 VDD2.n168 VDD2.n108 104.615
R2836 VDD2.n168 VDD2.n167 104.615
R2837 VDD2.n167 VDD2.n109 104.615
R2838 VDD2.n160 VDD2.n109 104.615
R2839 VDD2.n160 VDD2.n159 104.615
R2840 VDD2.n159 VDD2.n113 104.615
R2841 VDD2.n152 VDD2.n113 104.615
R2842 VDD2.n152 VDD2.n151 104.615
R2843 VDD2.n151 VDD2.n117 104.615
R2844 VDD2.n144 VDD2.n117 104.615
R2845 VDD2.n144 VDD2.n143 104.615
R2846 VDD2.n143 VDD2.n121 104.615
R2847 VDD2.n136 VDD2.n121 104.615
R2848 VDD2.n136 VDD2.n135 104.615
R2849 VDD2.n135 VDD2.n125 104.615
R2850 VDD2.n128 VDD2.n125 104.615
R2851 VDD2.n30 VDD2.n27 104.615
R2852 VDD2.n37 VDD2.n27 104.615
R2853 VDD2.n38 VDD2.n37 104.615
R2854 VDD2.n38 VDD2.n23 104.615
R2855 VDD2.n45 VDD2.n23 104.615
R2856 VDD2.n46 VDD2.n45 104.615
R2857 VDD2.n46 VDD2.n19 104.615
R2858 VDD2.n53 VDD2.n19 104.615
R2859 VDD2.n54 VDD2.n53 104.615
R2860 VDD2.n54 VDD2.n15 104.615
R2861 VDD2.n61 VDD2.n15 104.615
R2862 VDD2.n62 VDD2.n61 104.615
R2863 VDD2.n62 VDD2.n11 104.615
R2864 VDD2.n69 VDD2.n11 104.615
R2865 VDD2.n71 VDD2.n69 104.615
R2866 VDD2.n71 VDD2.n70 104.615
R2867 VDD2.n70 VDD2.n7 104.615
R2868 VDD2.n79 VDD2.n7 104.615
R2869 VDD2.n80 VDD2.n79 104.615
R2870 VDD2.n80 VDD2.n3 104.615
R2871 VDD2.n87 VDD2.n3 104.615
R2872 VDD2.n88 VDD2.n87 104.615
R2873 VDD2.n96 VDD2.n95 62.3567
R2874 VDD2 VDD2.n193 62.3539
R2875 VDD2.n192 VDD2.n191 61.3066
R2876 VDD2.n94 VDD2.n93 61.3065
R2877 VDD2.n128 VDD2.t0 52.3082
R2878 VDD2.n30 VDD2.t6 52.3082
R2879 VDD2.n94 VDD2.n92 50.9201
R2880 VDD2.n190 VDD2.n189 49.446
R2881 VDD2.n190 VDD2.n96 45.2261
R2882 VDD2.n129 VDD2.n127 15.6677
R2883 VDD2.n31 VDD2.n29 15.6677
R2884 VDD2.n175 VDD2.n174 13.1884
R2885 VDD2.n78 VDD2.n77 13.1884
R2886 VDD2.n178 VDD2.n103 12.8005
R2887 VDD2.n173 VDD2.n105 12.8005
R2888 VDD2.n130 VDD2.n126 12.8005
R2889 VDD2.n32 VDD2.n28 12.8005
R2890 VDD2.n76 VDD2.n8 12.8005
R2891 VDD2.n81 VDD2.n6 12.8005
R2892 VDD2.n179 VDD2.n101 12.0247
R2893 VDD2.n170 VDD2.n169 12.0247
R2894 VDD2.n134 VDD2.n133 12.0247
R2895 VDD2.n36 VDD2.n35 12.0247
R2896 VDD2.n73 VDD2.n72 12.0247
R2897 VDD2.n82 VDD2.n4 12.0247
R2898 VDD2.n183 VDD2.n182 11.249
R2899 VDD2.n166 VDD2.n107 11.249
R2900 VDD2.n137 VDD2.n124 11.249
R2901 VDD2.n39 VDD2.n26 11.249
R2902 VDD2.n68 VDD2.n10 11.249
R2903 VDD2.n86 VDD2.n85 11.249
R2904 VDD2.n186 VDD2.n99 10.4732
R2905 VDD2.n165 VDD2.n110 10.4732
R2906 VDD2.n138 VDD2.n122 10.4732
R2907 VDD2.n40 VDD2.n24 10.4732
R2908 VDD2.n67 VDD2.n12 10.4732
R2909 VDD2.n89 VDD2.n2 10.4732
R2910 VDD2.n187 VDD2.n97 9.69747
R2911 VDD2.n162 VDD2.n161 9.69747
R2912 VDD2.n142 VDD2.n141 9.69747
R2913 VDD2.n44 VDD2.n43 9.69747
R2914 VDD2.n64 VDD2.n63 9.69747
R2915 VDD2.n90 VDD2.n0 9.69747
R2916 VDD2.n189 VDD2.n188 9.45567
R2917 VDD2.n92 VDD2.n91 9.45567
R2918 VDD2.n155 VDD2.n154 9.3005
R2919 VDD2.n157 VDD2.n156 9.3005
R2920 VDD2.n112 VDD2.n111 9.3005
R2921 VDD2.n163 VDD2.n162 9.3005
R2922 VDD2.n165 VDD2.n164 9.3005
R2923 VDD2.n107 VDD2.n106 9.3005
R2924 VDD2.n171 VDD2.n170 9.3005
R2925 VDD2.n173 VDD2.n172 9.3005
R2926 VDD2.n188 VDD2.n187 9.3005
R2927 VDD2.n99 VDD2.n98 9.3005
R2928 VDD2.n182 VDD2.n181 9.3005
R2929 VDD2.n180 VDD2.n179 9.3005
R2930 VDD2.n103 VDD2.n102 9.3005
R2931 VDD2.n116 VDD2.n115 9.3005
R2932 VDD2.n149 VDD2.n148 9.3005
R2933 VDD2.n147 VDD2.n146 9.3005
R2934 VDD2.n120 VDD2.n119 9.3005
R2935 VDD2.n141 VDD2.n140 9.3005
R2936 VDD2.n139 VDD2.n138 9.3005
R2937 VDD2.n124 VDD2.n123 9.3005
R2938 VDD2.n133 VDD2.n132 9.3005
R2939 VDD2.n131 VDD2.n130 9.3005
R2940 VDD2.n91 VDD2.n90 9.3005
R2941 VDD2.n2 VDD2.n1 9.3005
R2942 VDD2.n85 VDD2.n84 9.3005
R2943 VDD2.n83 VDD2.n82 9.3005
R2944 VDD2.n6 VDD2.n5 9.3005
R2945 VDD2.n51 VDD2.n50 9.3005
R2946 VDD2.n49 VDD2.n48 9.3005
R2947 VDD2.n22 VDD2.n21 9.3005
R2948 VDD2.n43 VDD2.n42 9.3005
R2949 VDD2.n41 VDD2.n40 9.3005
R2950 VDD2.n26 VDD2.n25 9.3005
R2951 VDD2.n35 VDD2.n34 9.3005
R2952 VDD2.n33 VDD2.n32 9.3005
R2953 VDD2.n18 VDD2.n17 9.3005
R2954 VDD2.n57 VDD2.n56 9.3005
R2955 VDD2.n59 VDD2.n58 9.3005
R2956 VDD2.n14 VDD2.n13 9.3005
R2957 VDD2.n65 VDD2.n64 9.3005
R2958 VDD2.n67 VDD2.n66 9.3005
R2959 VDD2.n10 VDD2.n9 9.3005
R2960 VDD2.n74 VDD2.n73 9.3005
R2961 VDD2.n76 VDD2.n75 9.3005
R2962 VDD2.n158 VDD2.n112 8.92171
R2963 VDD2.n145 VDD2.n120 8.92171
R2964 VDD2.n47 VDD2.n22 8.92171
R2965 VDD2.n60 VDD2.n14 8.92171
R2966 VDD2.n157 VDD2.n114 8.14595
R2967 VDD2.n146 VDD2.n118 8.14595
R2968 VDD2.n48 VDD2.n20 8.14595
R2969 VDD2.n59 VDD2.n16 8.14595
R2970 VDD2.n154 VDD2.n153 7.3702
R2971 VDD2.n150 VDD2.n149 7.3702
R2972 VDD2.n52 VDD2.n51 7.3702
R2973 VDD2.n56 VDD2.n55 7.3702
R2974 VDD2.n153 VDD2.n116 6.59444
R2975 VDD2.n150 VDD2.n116 6.59444
R2976 VDD2.n52 VDD2.n18 6.59444
R2977 VDD2.n55 VDD2.n18 6.59444
R2978 VDD2.n154 VDD2.n114 5.81868
R2979 VDD2.n149 VDD2.n118 5.81868
R2980 VDD2.n51 VDD2.n20 5.81868
R2981 VDD2.n56 VDD2.n16 5.81868
R2982 VDD2.n158 VDD2.n157 5.04292
R2983 VDD2.n146 VDD2.n145 5.04292
R2984 VDD2.n48 VDD2.n47 5.04292
R2985 VDD2.n60 VDD2.n59 5.04292
R2986 VDD2.n131 VDD2.n127 4.38563
R2987 VDD2.n33 VDD2.n29 4.38563
R2988 VDD2.n189 VDD2.n97 4.26717
R2989 VDD2.n161 VDD2.n112 4.26717
R2990 VDD2.n142 VDD2.n120 4.26717
R2991 VDD2.n44 VDD2.n22 4.26717
R2992 VDD2.n63 VDD2.n14 4.26717
R2993 VDD2.n92 VDD2.n0 4.26717
R2994 VDD2.n187 VDD2.n186 3.49141
R2995 VDD2.n162 VDD2.n110 3.49141
R2996 VDD2.n141 VDD2.n122 3.49141
R2997 VDD2.n43 VDD2.n24 3.49141
R2998 VDD2.n64 VDD2.n12 3.49141
R2999 VDD2.n90 VDD2.n89 3.49141
R3000 VDD2.n183 VDD2.n99 2.71565
R3001 VDD2.n166 VDD2.n165 2.71565
R3002 VDD2.n138 VDD2.n137 2.71565
R3003 VDD2.n40 VDD2.n39 2.71565
R3004 VDD2.n68 VDD2.n67 2.71565
R3005 VDD2.n86 VDD2.n2 2.71565
R3006 VDD2.n182 VDD2.n101 1.93989
R3007 VDD2.n169 VDD2.n107 1.93989
R3008 VDD2.n134 VDD2.n124 1.93989
R3009 VDD2.n36 VDD2.n26 1.93989
R3010 VDD2.n72 VDD2.n10 1.93989
R3011 VDD2.n85 VDD2.n4 1.93989
R3012 VDD2.n192 VDD2.n190 1.47464
R3013 VDD2.n193 VDD2.t8 1.17697
R3014 VDD2.n193 VDD2.t4 1.17697
R3015 VDD2.n191 VDD2.t7 1.17697
R3016 VDD2.n191 VDD2.t2 1.17697
R3017 VDD2.n95 VDD2.t1 1.17697
R3018 VDD2.n95 VDD2.t9 1.17697
R3019 VDD2.n93 VDD2.t5 1.17697
R3020 VDD2.n93 VDD2.t3 1.17697
R3021 VDD2.n179 VDD2.n178 1.16414
R3022 VDD2.n170 VDD2.n105 1.16414
R3023 VDD2.n133 VDD2.n126 1.16414
R3024 VDD2.n35 VDD2.n28 1.16414
R3025 VDD2.n73 VDD2.n8 1.16414
R3026 VDD2.n82 VDD2.n81 1.16414
R3027 VDD2 VDD2.n192 0.427224
R3028 VDD2.n175 VDD2.n103 0.388379
R3029 VDD2.n174 VDD2.n173 0.388379
R3030 VDD2.n130 VDD2.n129 0.388379
R3031 VDD2.n32 VDD2.n31 0.388379
R3032 VDD2.n77 VDD2.n76 0.388379
R3033 VDD2.n78 VDD2.n6 0.388379
R3034 VDD2.n96 VDD2.n94 0.313688
R3035 VDD2.n188 VDD2.n98 0.155672
R3036 VDD2.n181 VDD2.n98 0.155672
R3037 VDD2.n181 VDD2.n180 0.155672
R3038 VDD2.n180 VDD2.n102 0.155672
R3039 VDD2.n172 VDD2.n102 0.155672
R3040 VDD2.n172 VDD2.n171 0.155672
R3041 VDD2.n171 VDD2.n106 0.155672
R3042 VDD2.n164 VDD2.n106 0.155672
R3043 VDD2.n164 VDD2.n163 0.155672
R3044 VDD2.n163 VDD2.n111 0.155672
R3045 VDD2.n156 VDD2.n111 0.155672
R3046 VDD2.n156 VDD2.n155 0.155672
R3047 VDD2.n155 VDD2.n115 0.155672
R3048 VDD2.n148 VDD2.n115 0.155672
R3049 VDD2.n148 VDD2.n147 0.155672
R3050 VDD2.n147 VDD2.n119 0.155672
R3051 VDD2.n140 VDD2.n119 0.155672
R3052 VDD2.n140 VDD2.n139 0.155672
R3053 VDD2.n139 VDD2.n123 0.155672
R3054 VDD2.n132 VDD2.n123 0.155672
R3055 VDD2.n132 VDD2.n131 0.155672
R3056 VDD2.n34 VDD2.n33 0.155672
R3057 VDD2.n34 VDD2.n25 0.155672
R3058 VDD2.n41 VDD2.n25 0.155672
R3059 VDD2.n42 VDD2.n41 0.155672
R3060 VDD2.n42 VDD2.n21 0.155672
R3061 VDD2.n49 VDD2.n21 0.155672
R3062 VDD2.n50 VDD2.n49 0.155672
R3063 VDD2.n50 VDD2.n17 0.155672
R3064 VDD2.n57 VDD2.n17 0.155672
R3065 VDD2.n58 VDD2.n57 0.155672
R3066 VDD2.n58 VDD2.n13 0.155672
R3067 VDD2.n65 VDD2.n13 0.155672
R3068 VDD2.n66 VDD2.n65 0.155672
R3069 VDD2.n66 VDD2.n9 0.155672
R3070 VDD2.n74 VDD2.n9 0.155672
R3071 VDD2.n75 VDD2.n74 0.155672
R3072 VDD2.n75 VDD2.n5 0.155672
R3073 VDD2.n83 VDD2.n5 0.155672
R3074 VDD2.n84 VDD2.n83 0.155672
R3075 VDD2.n84 VDD2.n1 0.155672
R3076 VDD2.n91 VDD2.n1 0.155672
C0 VDD1 VN 0.150595f
C1 VDD1 VP 12.708401f
C2 VDD1 VTAIL 14.281401f
C3 VDD2 VN 12.4358f
C4 VDD2 VP 0.428681f
C5 VDD2 VTAIL 14.3204f
C6 VP VN 7.497089f
C7 VN VTAIL 12.378401f
C8 VDD1 VDD2 1.38251f
C9 VP VTAIL 12.393f
C10 VDD2 B 6.642107f
C11 VDD1 B 6.610085f
C12 VTAIL B 9.035049f
C13 VN B 12.93595f
C14 VP B 11.104903f
C15 VDD2.n0 B 0.030819f
C16 VDD2.n1 B 0.022465f
C17 VDD2.n2 B 0.012072f
C18 VDD2.n3 B 0.028534f
C19 VDD2.n4 B 0.012782f
C20 VDD2.n5 B 0.022465f
C21 VDD2.n6 B 0.012072f
C22 VDD2.n7 B 0.028534f
C23 VDD2.n8 B 0.012782f
C24 VDD2.n9 B 0.022465f
C25 VDD2.n10 B 0.012072f
C26 VDD2.n11 B 0.028534f
C27 VDD2.n12 B 0.012782f
C28 VDD2.n13 B 0.022465f
C29 VDD2.n14 B 0.012072f
C30 VDD2.n15 B 0.028534f
C31 VDD2.n16 B 0.012782f
C32 VDD2.n17 B 0.022465f
C33 VDD2.n18 B 0.012072f
C34 VDD2.n19 B 0.028534f
C35 VDD2.n20 B 0.012782f
C36 VDD2.n21 B 0.022465f
C37 VDD2.n22 B 0.012072f
C38 VDD2.n23 B 0.028534f
C39 VDD2.n24 B 0.012782f
C40 VDD2.n25 B 0.022465f
C41 VDD2.n26 B 0.012072f
C42 VDD2.n27 B 0.028534f
C43 VDD2.n28 B 0.012782f
C44 VDD2.n29 B 0.156832f
C45 VDD2.t6 B 0.04719f
C46 VDD2.n30 B 0.0214f
C47 VDD2.n31 B 0.016856f
C48 VDD2.n32 B 0.012072f
C49 VDD2.n33 B 1.65004f
C50 VDD2.n34 B 0.022465f
C51 VDD2.n35 B 0.012072f
C52 VDD2.n36 B 0.012782f
C53 VDD2.n37 B 0.028534f
C54 VDD2.n38 B 0.028534f
C55 VDD2.n39 B 0.012782f
C56 VDD2.n40 B 0.012072f
C57 VDD2.n41 B 0.022465f
C58 VDD2.n42 B 0.022465f
C59 VDD2.n43 B 0.012072f
C60 VDD2.n44 B 0.012782f
C61 VDD2.n45 B 0.028534f
C62 VDD2.n46 B 0.028534f
C63 VDD2.n47 B 0.012782f
C64 VDD2.n48 B 0.012072f
C65 VDD2.n49 B 0.022465f
C66 VDD2.n50 B 0.022465f
C67 VDD2.n51 B 0.012072f
C68 VDD2.n52 B 0.012782f
C69 VDD2.n53 B 0.028534f
C70 VDD2.n54 B 0.028534f
C71 VDD2.n55 B 0.012782f
C72 VDD2.n56 B 0.012072f
C73 VDD2.n57 B 0.022465f
C74 VDD2.n58 B 0.022465f
C75 VDD2.n59 B 0.012072f
C76 VDD2.n60 B 0.012782f
C77 VDD2.n61 B 0.028534f
C78 VDD2.n62 B 0.028534f
C79 VDD2.n63 B 0.012782f
C80 VDD2.n64 B 0.012072f
C81 VDD2.n65 B 0.022465f
C82 VDD2.n66 B 0.022465f
C83 VDD2.n67 B 0.012072f
C84 VDD2.n68 B 0.012782f
C85 VDD2.n69 B 0.028534f
C86 VDD2.n70 B 0.028534f
C87 VDD2.n71 B 0.028534f
C88 VDD2.n72 B 0.012782f
C89 VDD2.n73 B 0.012072f
C90 VDD2.n74 B 0.022465f
C91 VDD2.n75 B 0.022465f
C92 VDD2.n76 B 0.012072f
C93 VDD2.n77 B 0.012427f
C94 VDD2.n78 B 0.012427f
C95 VDD2.n79 B 0.028534f
C96 VDD2.n80 B 0.028534f
C97 VDD2.n81 B 0.012782f
C98 VDD2.n82 B 0.012072f
C99 VDD2.n83 B 0.022465f
C100 VDD2.n84 B 0.022465f
C101 VDD2.n85 B 0.012072f
C102 VDD2.n86 B 0.012782f
C103 VDD2.n87 B 0.028534f
C104 VDD2.n88 B 0.06043f
C105 VDD2.n89 B 0.012782f
C106 VDD2.n90 B 0.012072f
C107 VDD2.n91 B 0.052848f
C108 VDD2.n92 B 0.053565f
C109 VDD2.t5 B 0.29878f
C110 VDD2.t3 B 0.29878f
C111 VDD2.n93 B 2.7149f
C112 VDD2.n94 B 0.46238f
C113 VDD2.t1 B 0.29878f
C114 VDD2.t9 B 0.29878f
C115 VDD2.n95 B 2.72126f
C116 VDD2.n96 B 2.30421f
C117 VDD2.n97 B 0.030819f
C118 VDD2.n98 B 0.022465f
C119 VDD2.n99 B 0.012072f
C120 VDD2.n100 B 0.028534f
C121 VDD2.n101 B 0.012782f
C122 VDD2.n102 B 0.022465f
C123 VDD2.n103 B 0.012072f
C124 VDD2.n104 B 0.028534f
C125 VDD2.n105 B 0.012782f
C126 VDD2.n106 B 0.022465f
C127 VDD2.n107 B 0.012072f
C128 VDD2.n108 B 0.028534f
C129 VDD2.n109 B 0.028534f
C130 VDD2.n110 B 0.012782f
C131 VDD2.n111 B 0.022465f
C132 VDD2.n112 B 0.012072f
C133 VDD2.n113 B 0.028534f
C134 VDD2.n114 B 0.012782f
C135 VDD2.n115 B 0.022465f
C136 VDD2.n116 B 0.012072f
C137 VDD2.n117 B 0.028534f
C138 VDD2.n118 B 0.012782f
C139 VDD2.n119 B 0.022465f
C140 VDD2.n120 B 0.012072f
C141 VDD2.n121 B 0.028534f
C142 VDD2.n122 B 0.012782f
C143 VDD2.n123 B 0.022465f
C144 VDD2.n124 B 0.012072f
C145 VDD2.n125 B 0.028534f
C146 VDD2.n126 B 0.012782f
C147 VDD2.n127 B 0.156832f
C148 VDD2.t0 B 0.04719f
C149 VDD2.n128 B 0.0214f
C150 VDD2.n129 B 0.016856f
C151 VDD2.n130 B 0.012072f
C152 VDD2.n131 B 1.65004f
C153 VDD2.n132 B 0.022465f
C154 VDD2.n133 B 0.012072f
C155 VDD2.n134 B 0.012782f
C156 VDD2.n135 B 0.028534f
C157 VDD2.n136 B 0.028534f
C158 VDD2.n137 B 0.012782f
C159 VDD2.n138 B 0.012072f
C160 VDD2.n139 B 0.022465f
C161 VDD2.n140 B 0.022465f
C162 VDD2.n141 B 0.012072f
C163 VDD2.n142 B 0.012782f
C164 VDD2.n143 B 0.028534f
C165 VDD2.n144 B 0.028534f
C166 VDD2.n145 B 0.012782f
C167 VDD2.n146 B 0.012072f
C168 VDD2.n147 B 0.022465f
C169 VDD2.n148 B 0.022465f
C170 VDD2.n149 B 0.012072f
C171 VDD2.n150 B 0.012782f
C172 VDD2.n151 B 0.028534f
C173 VDD2.n152 B 0.028534f
C174 VDD2.n153 B 0.012782f
C175 VDD2.n154 B 0.012072f
C176 VDD2.n155 B 0.022465f
C177 VDD2.n156 B 0.022465f
C178 VDD2.n157 B 0.012072f
C179 VDD2.n158 B 0.012782f
C180 VDD2.n159 B 0.028534f
C181 VDD2.n160 B 0.028534f
C182 VDD2.n161 B 0.012782f
C183 VDD2.n162 B 0.012072f
C184 VDD2.n163 B 0.022465f
C185 VDD2.n164 B 0.022465f
C186 VDD2.n165 B 0.012072f
C187 VDD2.n166 B 0.012782f
C188 VDD2.n167 B 0.028534f
C189 VDD2.n168 B 0.028534f
C190 VDD2.n169 B 0.012782f
C191 VDD2.n170 B 0.012072f
C192 VDD2.n171 B 0.022465f
C193 VDD2.n172 B 0.022465f
C194 VDD2.n173 B 0.012072f
C195 VDD2.n174 B 0.012427f
C196 VDD2.n175 B 0.012427f
C197 VDD2.n176 B 0.028534f
C198 VDD2.n177 B 0.028534f
C199 VDD2.n178 B 0.012782f
C200 VDD2.n179 B 0.012072f
C201 VDD2.n180 B 0.022465f
C202 VDD2.n181 B 0.022465f
C203 VDD2.n182 B 0.012072f
C204 VDD2.n183 B 0.012782f
C205 VDD2.n184 B 0.028534f
C206 VDD2.n185 B 0.06043f
C207 VDD2.n186 B 0.012782f
C208 VDD2.n187 B 0.012072f
C209 VDD2.n188 B 0.052848f
C210 VDD2.n189 B 0.049208f
C211 VDD2.n190 B 2.50614f
C212 VDD2.t7 B 0.29878f
C213 VDD2.t2 B 0.29878f
C214 VDD2.n191 B 2.71491f
C215 VDD2.n192 B 0.322788f
C216 VDD2.t8 B 0.29878f
C217 VDD2.t4 B 0.29878f
C218 VDD2.n193 B 2.72123f
C219 VN.n0 B 0.030735f
C220 VN.t0 B 1.96087f
C221 VN.n1 B 0.050437f
C222 VN.n2 B 0.030735f
C223 VN.t8 B 1.96087f
C224 VN.n3 B 0.047277f
C225 VN.n4 B 0.030735f
C226 VN.t4 B 1.96087f
C227 VN.n5 B 0.761468f
C228 VN.t3 B 2.04181f
C229 VN.n6 B 0.765264f
C230 VN.n7 B 0.190856f
C231 VN.n8 B 0.053849f
C232 VN.n9 B 0.029494f
C233 VN.t6 B 1.96087f
C234 VN.n10 B 0.695111f
C235 VN.n11 B 0.047277f
C236 VN.n12 B 0.030735f
C237 VN.n13 B 0.030735f
C238 VN.n14 B 0.030735f
C239 VN.n15 B 0.029494f
C240 VN.n16 B 0.053849f
C241 VN.n17 B 0.695111f
C242 VN.n18 B 0.031264f
C243 VN.n19 B 0.030735f
C244 VN.n20 B 0.030735f
C245 VN.n21 B 0.030735f
C246 VN.n22 B 0.039304f
C247 VN.n23 B 0.038617f
C248 VN.n24 B 0.749751f
C249 VN.n25 B 0.029289f
C250 VN.n26 B 0.030735f
C251 VN.t9 B 1.96087f
C252 VN.n27 B 0.050437f
C253 VN.n28 B 0.030735f
C254 VN.t2 B 1.96087f
C255 VN.n29 B 0.047277f
C256 VN.n30 B 0.030735f
C257 VN.t7 B 1.96087f
C258 VN.n31 B 0.695111f
C259 VN.t1 B 1.96087f
C260 VN.n32 B 0.761468f
C261 VN.t5 B 2.04181f
C262 VN.n33 B 0.765264f
C263 VN.n34 B 0.190856f
C264 VN.n35 B 0.053849f
C265 VN.n36 B 0.029494f
C266 VN.n37 B 0.047277f
C267 VN.n38 B 0.030735f
C268 VN.n39 B 0.030735f
C269 VN.n40 B 0.030735f
C270 VN.n41 B 0.029494f
C271 VN.n42 B 0.053849f
C272 VN.n43 B 0.695111f
C273 VN.n44 B 0.031264f
C274 VN.n45 B 0.030735f
C275 VN.n46 B 0.030735f
C276 VN.n47 B 0.030735f
C277 VN.n48 B 0.039304f
C278 VN.n49 B 0.038617f
C279 VN.n50 B 0.749751f
C280 VN.n51 B 1.69701f
C281 VTAIL.t1 B 0.315354f
C282 VTAIL.t6 B 0.315354f
C283 VTAIL.n0 B 2.79414f
C284 VTAIL.n1 B 0.415738f
C285 VTAIL.n2 B 0.032529f
C286 VTAIL.n3 B 0.023712f
C287 VTAIL.n4 B 0.012742f
C288 VTAIL.n5 B 0.030116f
C289 VTAIL.n6 B 0.013491f
C290 VTAIL.n7 B 0.023712f
C291 VTAIL.n8 B 0.012742f
C292 VTAIL.n9 B 0.030116f
C293 VTAIL.n10 B 0.013491f
C294 VTAIL.n11 B 0.023712f
C295 VTAIL.n12 B 0.012742f
C296 VTAIL.n13 B 0.030116f
C297 VTAIL.n14 B 0.013491f
C298 VTAIL.n15 B 0.023712f
C299 VTAIL.n16 B 0.012742f
C300 VTAIL.n17 B 0.030116f
C301 VTAIL.n18 B 0.013491f
C302 VTAIL.n19 B 0.023712f
C303 VTAIL.n20 B 0.012742f
C304 VTAIL.n21 B 0.030116f
C305 VTAIL.n22 B 0.013491f
C306 VTAIL.n23 B 0.023712f
C307 VTAIL.n24 B 0.012742f
C308 VTAIL.n25 B 0.030116f
C309 VTAIL.n26 B 0.013491f
C310 VTAIL.n27 B 0.023712f
C311 VTAIL.n28 B 0.012742f
C312 VTAIL.n29 B 0.030116f
C313 VTAIL.n30 B 0.013491f
C314 VTAIL.n31 B 0.165531f
C315 VTAIL.t15 B 0.049807f
C316 VTAIL.n32 B 0.022587f
C317 VTAIL.n33 B 0.017791f
C318 VTAIL.n34 B 0.012742f
C319 VTAIL.n35 B 1.74158f
C320 VTAIL.n36 B 0.023712f
C321 VTAIL.n37 B 0.012742f
C322 VTAIL.n38 B 0.013491f
C323 VTAIL.n39 B 0.030116f
C324 VTAIL.n40 B 0.030116f
C325 VTAIL.n41 B 0.013491f
C326 VTAIL.n42 B 0.012742f
C327 VTAIL.n43 B 0.023712f
C328 VTAIL.n44 B 0.023712f
C329 VTAIL.n45 B 0.012742f
C330 VTAIL.n46 B 0.013491f
C331 VTAIL.n47 B 0.030116f
C332 VTAIL.n48 B 0.030116f
C333 VTAIL.n49 B 0.013491f
C334 VTAIL.n50 B 0.012742f
C335 VTAIL.n51 B 0.023712f
C336 VTAIL.n52 B 0.023712f
C337 VTAIL.n53 B 0.012742f
C338 VTAIL.n54 B 0.013491f
C339 VTAIL.n55 B 0.030116f
C340 VTAIL.n56 B 0.030116f
C341 VTAIL.n57 B 0.013491f
C342 VTAIL.n58 B 0.012742f
C343 VTAIL.n59 B 0.023712f
C344 VTAIL.n60 B 0.023712f
C345 VTAIL.n61 B 0.012742f
C346 VTAIL.n62 B 0.013491f
C347 VTAIL.n63 B 0.030116f
C348 VTAIL.n64 B 0.030116f
C349 VTAIL.n65 B 0.013491f
C350 VTAIL.n66 B 0.012742f
C351 VTAIL.n67 B 0.023712f
C352 VTAIL.n68 B 0.023712f
C353 VTAIL.n69 B 0.012742f
C354 VTAIL.n70 B 0.013491f
C355 VTAIL.n71 B 0.030116f
C356 VTAIL.n72 B 0.030116f
C357 VTAIL.n73 B 0.030116f
C358 VTAIL.n74 B 0.013491f
C359 VTAIL.n75 B 0.012742f
C360 VTAIL.n76 B 0.023712f
C361 VTAIL.n77 B 0.023712f
C362 VTAIL.n78 B 0.012742f
C363 VTAIL.n79 B 0.013116f
C364 VTAIL.n80 B 0.013116f
C365 VTAIL.n81 B 0.030116f
C366 VTAIL.n82 B 0.030116f
C367 VTAIL.n83 B 0.013491f
C368 VTAIL.n84 B 0.012742f
C369 VTAIL.n85 B 0.023712f
C370 VTAIL.n86 B 0.023712f
C371 VTAIL.n87 B 0.012742f
C372 VTAIL.n88 B 0.013491f
C373 VTAIL.n89 B 0.030116f
C374 VTAIL.n90 B 0.063782f
C375 VTAIL.n91 B 0.013491f
C376 VTAIL.n92 B 0.012742f
C377 VTAIL.n93 B 0.05578f
C378 VTAIL.n94 B 0.035573f
C379 VTAIL.n95 B 0.225642f
C380 VTAIL.t18 B 0.315354f
C381 VTAIL.t12 B 0.315354f
C382 VTAIL.n96 B 2.79414f
C383 VTAIL.n97 B 0.459867f
C384 VTAIL.t17 B 0.315354f
C385 VTAIL.t19 B 0.315354f
C386 VTAIL.n98 B 2.79414f
C387 VTAIL.n99 B 2.00311f
C388 VTAIL.t2 B 0.315354f
C389 VTAIL.t3 B 0.315354f
C390 VTAIL.n100 B 2.79415f
C391 VTAIL.n101 B 2.0031f
C392 VTAIL.t7 B 0.315354f
C393 VTAIL.t4 B 0.315354f
C394 VTAIL.n102 B 2.79415f
C395 VTAIL.n103 B 0.459854f
C396 VTAIL.n104 B 0.032529f
C397 VTAIL.n105 B 0.023712f
C398 VTAIL.n106 B 0.012742f
C399 VTAIL.n107 B 0.030116f
C400 VTAIL.n108 B 0.013491f
C401 VTAIL.n109 B 0.023712f
C402 VTAIL.n110 B 0.012742f
C403 VTAIL.n111 B 0.030116f
C404 VTAIL.n112 B 0.013491f
C405 VTAIL.n113 B 0.023712f
C406 VTAIL.n114 B 0.012742f
C407 VTAIL.n115 B 0.030116f
C408 VTAIL.n116 B 0.030116f
C409 VTAIL.n117 B 0.013491f
C410 VTAIL.n118 B 0.023712f
C411 VTAIL.n119 B 0.012742f
C412 VTAIL.n120 B 0.030116f
C413 VTAIL.n121 B 0.013491f
C414 VTAIL.n122 B 0.023712f
C415 VTAIL.n123 B 0.012742f
C416 VTAIL.n124 B 0.030116f
C417 VTAIL.n125 B 0.013491f
C418 VTAIL.n126 B 0.023712f
C419 VTAIL.n127 B 0.012742f
C420 VTAIL.n128 B 0.030116f
C421 VTAIL.n129 B 0.013491f
C422 VTAIL.n130 B 0.023712f
C423 VTAIL.n131 B 0.012742f
C424 VTAIL.n132 B 0.030116f
C425 VTAIL.n133 B 0.013491f
C426 VTAIL.n134 B 0.165531f
C427 VTAIL.t5 B 0.049807f
C428 VTAIL.n135 B 0.022587f
C429 VTAIL.n136 B 0.017791f
C430 VTAIL.n137 B 0.012742f
C431 VTAIL.n138 B 1.74158f
C432 VTAIL.n139 B 0.023712f
C433 VTAIL.n140 B 0.012742f
C434 VTAIL.n141 B 0.013491f
C435 VTAIL.n142 B 0.030116f
C436 VTAIL.n143 B 0.030116f
C437 VTAIL.n144 B 0.013491f
C438 VTAIL.n145 B 0.012742f
C439 VTAIL.n146 B 0.023712f
C440 VTAIL.n147 B 0.023712f
C441 VTAIL.n148 B 0.012742f
C442 VTAIL.n149 B 0.013491f
C443 VTAIL.n150 B 0.030116f
C444 VTAIL.n151 B 0.030116f
C445 VTAIL.n152 B 0.013491f
C446 VTAIL.n153 B 0.012742f
C447 VTAIL.n154 B 0.023712f
C448 VTAIL.n155 B 0.023712f
C449 VTAIL.n156 B 0.012742f
C450 VTAIL.n157 B 0.013491f
C451 VTAIL.n158 B 0.030116f
C452 VTAIL.n159 B 0.030116f
C453 VTAIL.n160 B 0.013491f
C454 VTAIL.n161 B 0.012742f
C455 VTAIL.n162 B 0.023712f
C456 VTAIL.n163 B 0.023712f
C457 VTAIL.n164 B 0.012742f
C458 VTAIL.n165 B 0.013491f
C459 VTAIL.n166 B 0.030116f
C460 VTAIL.n167 B 0.030116f
C461 VTAIL.n168 B 0.013491f
C462 VTAIL.n169 B 0.012742f
C463 VTAIL.n170 B 0.023712f
C464 VTAIL.n171 B 0.023712f
C465 VTAIL.n172 B 0.012742f
C466 VTAIL.n173 B 0.013491f
C467 VTAIL.n174 B 0.030116f
C468 VTAIL.n175 B 0.030116f
C469 VTAIL.n176 B 0.013491f
C470 VTAIL.n177 B 0.012742f
C471 VTAIL.n178 B 0.023712f
C472 VTAIL.n179 B 0.023712f
C473 VTAIL.n180 B 0.012742f
C474 VTAIL.n181 B 0.013116f
C475 VTAIL.n182 B 0.013116f
C476 VTAIL.n183 B 0.030116f
C477 VTAIL.n184 B 0.030116f
C478 VTAIL.n185 B 0.013491f
C479 VTAIL.n186 B 0.012742f
C480 VTAIL.n187 B 0.023712f
C481 VTAIL.n188 B 0.023712f
C482 VTAIL.n189 B 0.012742f
C483 VTAIL.n190 B 0.013491f
C484 VTAIL.n191 B 0.030116f
C485 VTAIL.n192 B 0.063782f
C486 VTAIL.n193 B 0.013491f
C487 VTAIL.n194 B 0.012742f
C488 VTAIL.n195 B 0.05578f
C489 VTAIL.n196 B 0.035573f
C490 VTAIL.n197 B 0.225642f
C491 VTAIL.t14 B 0.315354f
C492 VTAIL.t11 B 0.315354f
C493 VTAIL.n198 B 2.79415f
C494 VTAIL.n199 B 0.439436f
C495 VTAIL.t13 B 0.315354f
C496 VTAIL.t10 B 0.315354f
C497 VTAIL.n200 B 2.79415f
C498 VTAIL.n201 B 0.459854f
C499 VTAIL.n202 B 0.032529f
C500 VTAIL.n203 B 0.023712f
C501 VTAIL.n204 B 0.012742f
C502 VTAIL.n205 B 0.030116f
C503 VTAIL.n206 B 0.013491f
C504 VTAIL.n207 B 0.023712f
C505 VTAIL.n208 B 0.012742f
C506 VTAIL.n209 B 0.030116f
C507 VTAIL.n210 B 0.013491f
C508 VTAIL.n211 B 0.023712f
C509 VTAIL.n212 B 0.012742f
C510 VTAIL.n213 B 0.030116f
C511 VTAIL.n214 B 0.030116f
C512 VTAIL.n215 B 0.013491f
C513 VTAIL.n216 B 0.023712f
C514 VTAIL.n217 B 0.012742f
C515 VTAIL.n218 B 0.030116f
C516 VTAIL.n219 B 0.013491f
C517 VTAIL.n220 B 0.023712f
C518 VTAIL.n221 B 0.012742f
C519 VTAIL.n222 B 0.030116f
C520 VTAIL.n223 B 0.013491f
C521 VTAIL.n224 B 0.023712f
C522 VTAIL.n225 B 0.012742f
C523 VTAIL.n226 B 0.030116f
C524 VTAIL.n227 B 0.013491f
C525 VTAIL.n228 B 0.023712f
C526 VTAIL.n229 B 0.012742f
C527 VTAIL.n230 B 0.030116f
C528 VTAIL.n231 B 0.013491f
C529 VTAIL.n232 B 0.165531f
C530 VTAIL.t16 B 0.049807f
C531 VTAIL.n233 B 0.022587f
C532 VTAIL.n234 B 0.017791f
C533 VTAIL.n235 B 0.012742f
C534 VTAIL.n236 B 1.74158f
C535 VTAIL.n237 B 0.023712f
C536 VTAIL.n238 B 0.012742f
C537 VTAIL.n239 B 0.013491f
C538 VTAIL.n240 B 0.030116f
C539 VTAIL.n241 B 0.030116f
C540 VTAIL.n242 B 0.013491f
C541 VTAIL.n243 B 0.012742f
C542 VTAIL.n244 B 0.023712f
C543 VTAIL.n245 B 0.023712f
C544 VTAIL.n246 B 0.012742f
C545 VTAIL.n247 B 0.013491f
C546 VTAIL.n248 B 0.030116f
C547 VTAIL.n249 B 0.030116f
C548 VTAIL.n250 B 0.013491f
C549 VTAIL.n251 B 0.012742f
C550 VTAIL.n252 B 0.023712f
C551 VTAIL.n253 B 0.023712f
C552 VTAIL.n254 B 0.012742f
C553 VTAIL.n255 B 0.013491f
C554 VTAIL.n256 B 0.030116f
C555 VTAIL.n257 B 0.030116f
C556 VTAIL.n258 B 0.013491f
C557 VTAIL.n259 B 0.012742f
C558 VTAIL.n260 B 0.023712f
C559 VTAIL.n261 B 0.023712f
C560 VTAIL.n262 B 0.012742f
C561 VTAIL.n263 B 0.013491f
C562 VTAIL.n264 B 0.030116f
C563 VTAIL.n265 B 0.030116f
C564 VTAIL.n266 B 0.013491f
C565 VTAIL.n267 B 0.012742f
C566 VTAIL.n268 B 0.023712f
C567 VTAIL.n269 B 0.023712f
C568 VTAIL.n270 B 0.012742f
C569 VTAIL.n271 B 0.013491f
C570 VTAIL.n272 B 0.030116f
C571 VTAIL.n273 B 0.030116f
C572 VTAIL.n274 B 0.013491f
C573 VTAIL.n275 B 0.012742f
C574 VTAIL.n276 B 0.023712f
C575 VTAIL.n277 B 0.023712f
C576 VTAIL.n278 B 0.012742f
C577 VTAIL.n279 B 0.013116f
C578 VTAIL.n280 B 0.013116f
C579 VTAIL.n281 B 0.030116f
C580 VTAIL.n282 B 0.030116f
C581 VTAIL.n283 B 0.013491f
C582 VTAIL.n284 B 0.012742f
C583 VTAIL.n285 B 0.023712f
C584 VTAIL.n286 B 0.023712f
C585 VTAIL.n287 B 0.012742f
C586 VTAIL.n288 B 0.013491f
C587 VTAIL.n289 B 0.030116f
C588 VTAIL.n290 B 0.063782f
C589 VTAIL.n291 B 0.013491f
C590 VTAIL.n292 B 0.012742f
C591 VTAIL.n293 B 0.05578f
C592 VTAIL.n294 B 0.035573f
C593 VTAIL.n295 B 1.67667f
C594 VTAIL.n296 B 0.032529f
C595 VTAIL.n297 B 0.023712f
C596 VTAIL.n298 B 0.012742f
C597 VTAIL.n299 B 0.030116f
C598 VTAIL.n300 B 0.013491f
C599 VTAIL.n301 B 0.023712f
C600 VTAIL.n302 B 0.012742f
C601 VTAIL.n303 B 0.030116f
C602 VTAIL.n304 B 0.013491f
C603 VTAIL.n305 B 0.023712f
C604 VTAIL.n306 B 0.012742f
C605 VTAIL.n307 B 0.030116f
C606 VTAIL.n308 B 0.013491f
C607 VTAIL.n309 B 0.023712f
C608 VTAIL.n310 B 0.012742f
C609 VTAIL.n311 B 0.030116f
C610 VTAIL.n312 B 0.013491f
C611 VTAIL.n313 B 0.023712f
C612 VTAIL.n314 B 0.012742f
C613 VTAIL.n315 B 0.030116f
C614 VTAIL.n316 B 0.013491f
C615 VTAIL.n317 B 0.023712f
C616 VTAIL.n318 B 0.012742f
C617 VTAIL.n319 B 0.030116f
C618 VTAIL.n320 B 0.013491f
C619 VTAIL.n321 B 0.023712f
C620 VTAIL.n322 B 0.012742f
C621 VTAIL.n323 B 0.030116f
C622 VTAIL.n324 B 0.013491f
C623 VTAIL.n325 B 0.165531f
C624 VTAIL.t9 B 0.049807f
C625 VTAIL.n326 B 0.022587f
C626 VTAIL.n327 B 0.017791f
C627 VTAIL.n328 B 0.012742f
C628 VTAIL.n329 B 1.74158f
C629 VTAIL.n330 B 0.023712f
C630 VTAIL.n331 B 0.012742f
C631 VTAIL.n332 B 0.013491f
C632 VTAIL.n333 B 0.030116f
C633 VTAIL.n334 B 0.030116f
C634 VTAIL.n335 B 0.013491f
C635 VTAIL.n336 B 0.012742f
C636 VTAIL.n337 B 0.023712f
C637 VTAIL.n338 B 0.023712f
C638 VTAIL.n339 B 0.012742f
C639 VTAIL.n340 B 0.013491f
C640 VTAIL.n341 B 0.030116f
C641 VTAIL.n342 B 0.030116f
C642 VTAIL.n343 B 0.013491f
C643 VTAIL.n344 B 0.012742f
C644 VTAIL.n345 B 0.023712f
C645 VTAIL.n346 B 0.023712f
C646 VTAIL.n347 B 0.012742f
C647 VTAIL.n348 B 0.013491f
C648 VTAIL.n349 B 0.030116f
C649 VTAIL.n350 B 0.030116f
C650 VTAIL.n351 B 0.013491f
C651 VTAIL.n352 B 0.012742f
C652 VTAIL.n353 B 0.023712f
C653 VTAIL.n354 B 0.023712f
C654 VTAIL.n355 B 0.012742f
C655 VTAIL.n356 B 0.013491f
C656 VTAIL.n357 B 0.030116f
C657 VTAIL.n358 B 0.030116f
C658 VTAIL.n359 B 0.013491f
C659 VTAIL.n360 B 0.012742f
C660 VTAIL.n361 B 0.023712f
C661 VTAIL.n362 B 0.023712f
C662 VTAIL.n363 B 0.012742f
C663 VTAIL.n364 B 0.013491f
C664 VTAIL.n365 B 0.030116f
C665 VTAIL.n366 B 0.030116f
C666 VTAIL.n367 B 0.030116f
C667 VTAIL.n368 B 0.013491f
C668 VTAIL.n369 B 0.012742f
C669 VTAIL.n370 B 0.023712f
C670 VTAIL.n371 B 0.023712f
C671 VTAIL.n372 B 0.012742f
C672 VTAIL.n373 B 0.013116f
C673 VTAIL.n374 B 0.013116f
C674 VTAIL.n375 B 0.030116f
C675 VTAIL.n376 B 0.030116f
C676 VTAIL.n377 B 0.013491f
C677 VTAIL.n378 B 0.012742f
C678 VTAIL.n379 B 0.023712f
C679 VTAIL.n380 B 0.023712f
C680 VTAIL.n381 B 0.012742f
C681 VTAIL.n382 B 0.013491f
C682 VTAIL.n383 B 0.030116f
C683 VTAIL.n384 B 0.063782f
C684 VTAIL.n385 B 0.013491f
C685 VTAIL.n386 B 0.012742f
C686 VTAIL.n387 B 0.05578f
C687 VTAIL.n388 B 0.035573f
C688 VTAIL.n389 B 1.67667f
C689 VTAIL.t8 B 0.315354f
C690 VTAIL.t0 B 0.315354f
C691 VTAIL.n390 B 2.79414f
C692 VTAIL.n391 B 0.370949f
C693 VDD1.n0 B 0.031069f
C694 VDD1.n1 B 0.022647f
C695 VDD1.n2 B 0.01217f
C696 VDD1.n3 B 0.028765f
C697 VDD1.n4 B 0.012886f
C698 VDD1.n5 B 0.022647f
C699 VDD1.n6 B 0.01217f
C700 VDD1.n7 B 0.028765f
C701 VDD1.n8 B 0.012886f
C702 VDD1.n9 B 0.022647f
C703 VDD1.n10 B 0.01217f
C704 VDD1.n11 B 0.028765f
C705 VDD1.n12 B 0.028765f
C706 VDD1.n13 B 0.012886f
C707 VDD1.n14 B 0.022647f
C708 VDD1.n15 B 0.01217f
C709 VDD1.n16 B 0.028765f
C710 VDD1.n17 B 0.012886f
C711 VDD1.n18 B 0.022647f
C712 VDD1.n19 B 0.01217f
C713 VDD1.n20 B 0.028765f
C714 VDD1.n21 B 0.012886f
C715 VDD1.n22 B 0.022647f
C716 VDD1.n23 B 0.01217f
C717 VDD1.n24 B 0.028765f
C718 VDD1.n25 B 0.012886f
C719 VDD1.n26 B 0.022647f
C720 VDD1.n27 B 0.01217f
C721 VDD1.n28 B 0.028765f
C722 VDD1.n29 B 0.012886f
C723 VDD1.n30 B 0.158102f
C724 VDD1.t4 B 0.047572f
C725 VDD1.n31 B 0.021574f
C726 VDD1.n32 B 0.016992f
C727 VDD1.n33 B 0.01217f
C728 VDD1.n34 B 1.66341f
C729 VDD1.n35 B 0.022647f
C730 VDD1.n36 B 0.01217f
C731 VDD1.n37 B 0.012886f
C732 VDD1.n38 B 0.028765f
C733 VDD1.n39 B 0.028765f
C734 VDD1.n40 B 0.012886f
C735 VDD1.n41 B 0.01217f
C736 VDD1.n42 B 0.022647f
C737 VDD1.n43 B 0.022647f
C738 VDD1.n44 B 0.01217f
C739 VDD1.n45 B 0.012886f
C740 VDD1.n46 B 0.028765f
C741 VDD1.n47 B 0.028765f
C742 VDD1.n48 B 0.012886f
C743 VDD1.n49 B 0.01217f
C744 VDD1.n50 B 0.022647f
C745 VDD1.n51 B 0.022647f
C746 VDD1.n52 B 0.01217f
C747 VDD1.n53 B 0.012886f
C748 VDD1.n54 B 0.028765f
C749 VDD1.n55 B 0.028765f
C750 VDD1.n56 B 0.012886f
C751 VDD1.n57 B 0.01217f
C752 VDD1.n58 B 0.022647f
C753 VDD1.n59 B 0.022647f
C754 VDD1.n60 B 0.01217f
C755 VDD1.n61 B 0.012886f
C756 VDD1.n62 B 0.028765f
C757 VDD1.n63 B 0.028765f
C758 VDD1.n64 B 0.012886f
C759 VDD1.n65 B 0.01217f
C760 VDD1.n66 B 0.022647f
C761 VDD1.n67 B 0.022647f
C762 VDD1.n68 B 0.01217f
C763 VDD1.n69 B 0.012886f
C764 VDD1.n70 B 0.028765f
C765 VDD1.n71 B 0.028765f
C766 VDD1.n72 B 0.012886f
C767 VDD1.n73 B 0.01217f
C768 VDD1.n74 B 0.022647f
C769 VDD1.n75 B 0.022647f
C770 VDD1.n76 B 0.01217f
C771 VDD1.n77 B 0.012528f
C772 VDD1.n78 B 0.012528f
C773 VDD1.n79 B 0.028765f
C774 VDD1.n80 B 0.028765f
C775 VDD1.n81 B 0.012886f
C776 VDD1.n82 B 0.01217f
C777 VDD1.n83 B 0.022647f
C778 VDD1.n84 B 0.022647f
C779 VDD1.n85 B 0.01217f
C780 VDD1.n86 B 0.012886f
C781 VDD1.n87 B 0.028765f
C782 VDD1.n88 B 0.06092f
C783 VDD1.n89 B 0.012886f
C784 VDD1.n90 B 0.01217f
C785 VDD1.n91 B 0.053277f
C786 VDD1.n92 B 0.053999f
C787 VDD1.t1 B 0.301201f
C788 VDD1.t9 B 0.301201f
C789 VDD1.n93 B 2.73691f
C790 VDD1.n94 B 0.472727f
C791 VDD1.n95 B 0.031069f
C792 VDD1.n96 B 0.022647f
C793 VDD1.n97 B 0.01217f
C794 VDD1.n98 B 0.028765f
C795 VDD1.n99 B 0.012886f
C796 VDD1.n100 B 0.022647f
C797 VDD1.n101 B 0.01217f
C798 VDD1.n102 B 0.028765f
C799 VDD1.n103 B 0.012886f
C800 VDD1.n104 B 0.022647f
C801 VDD1.n105 B 0.01217f
C802 VDD1.n106 B 0.028765f
C803 VDD1.n107 B 0.012886f
C804 VDD1.n108 B 0.022647f
C805 VDD1.n109 B 0.01217f
C806 VDD1.n110 B 0.028765f
C807 VDD1.n111 B 0.012886f
C808 VDD1.n112 B 0.022647f
C809 VDD1.n113 B 0.01217f
C810 VDD1.n114 B 0.028765f
C811 VDD1.n115 B 0.012886f
C812 VDD1.n116 B 0.022647f
C813 VDD1.n117 B 0.01217f
C814 VDD1.n118 B 0.028765f
C815 VDD1.n119 B 0.012886f
C816 VDD1.n120 B 0.022647f
C817 VDD1.n121 B 0.01217f
C818 VDD1.n122 B 0.028765f
C819 VDD1.n123 B 0.012886f
C820 VDD1.n124 B 0.158102f
C821 VDD1.t7 B 0.047572f
C822 VDD1.n125 B 0.021574f
C823 VDD1.n126 B 0.016992f
C824 VDD1.n127 B 0.01217f
C825 VDD1.n128 B 1.66341f
C826 VDD1.n129 B 0.022647f
C827 VDD1.n130 B 0.01217f
C828 VDD1.n131 B 0.012886f
C829 VDD1.n132 B 0.028765f
C830 VDD1.n133 B 0.028765f
C831 VDD1.n134 B 0.012886f
C832 VDD1.n135 B 0.01217f
C833 VDD1.n136 B 0.022647f
C834 VDD1.n137 B 0.022647f
C835 VDD1.n138 B 0.01217f
C836 VDD1.n139 B 0.012886f
C837 VDD1.n140 B 0.028765f
C838 VDD1.n141 B 0.028765f
C839 VDD1.n142 B 0.012886f
C840 VDD1.n143 B 0.01217f
C841 VDD1.n144 B 0.022647f
C842 VDD1.n145 B 0.022647f
C843 VDD1.n146 B 0.01217f
C844 VDD1.n147 B 0.012886f
C845 VDD1.n148 B 0.028765f
C846 VDD1.n149 B 0.028765f
C847 VDD1.n150 B 0.012886f
C848 VDD1.n151 B 0.01217f
C849 VDD1.n152 B 0.022647f
C850 VDD1.n153 B 0.022647f
C851 VDD1.n154 B 0.01217f
C852 VDD1.n155 B 0.012886f
C853 VDD1.n156 B 0.028765f
C854 VDD1.n157 B 0.028765f
C855 VDD1.n158 B 0.012886f
C856 VDD1.n159 B 0.01217f
C857 VDD1.n160 B 0.022647f
C858 VDD1.n161 B 0.022647f
C859 VDD1.n162 B 0.01217f
C860 VDD1.n163 B 0.012886f
C861 VDD1.n164 B 0.028765f
C862 VDD1.n165 B 0.028765f
C863 VDD1.n166 B 0.028765f
C864 VDD1.n167 B 0.012886f
C865 VDD1.n168 B 0.01217f
C866 VDD1.n169 B 0.022647f
C867 VDD1.n170 B 0.022647f
C868 VDD1.n171 B 0.01217f
C869 VDD1.n172 B 0.012528f
C870 VDD1.n173 B 0.012528f
C871 VDD1.n174 B 0.028765f
C872 VDD1.n175 B 0.028765f
C873 VDD1.n176 B 0.012886f
C874 VDD1.n177 B 0.01217f
C875 VDD1.n178 B 0.022647f
C876 VDD1.n179 B 0.022647f
C877 VDD1.n180 B 0.01217f
C878 VDD1.n181 B 0.012886f
C879 VDD1.n182 B 0.028765f
C880 VDD1.n183 B 0.06092f
C881 VDD1.n184 B 0.012886f
C882 VDD1.n185 B 0.01217f
C883 VDD1.n186 B 0.053277f
C884 VDD1.n187 B 0.053999f
C885 VDD1.t3 B 0.301201f
C886 VDD1.t2 B 0.301201f
C887 VDD1.n188 B 2.7369f
C888 VDD1.n189 B 0.466127f
C889 VDD1.t8 B 0.301201f
C890 VDD1.t5 B 0.301201f
C891 VDD1.n190 B 2.74331f
C892 VDD1.n191 B 2.40936f
C893 VDD1.t0 B 0.301201f
C894 VDD1.t6 B 0.301201f
C895 VDD1.n192 B 2.7369f
C896 VDD1.n193 B 2.75172f
C897 VP.n0 B 0.031062f
C898 VP.t4 B 1.98173f
C899 VP.n1 B 0.050974f
C900 VP.n2 B 0.031062f
C901 VP.t7 B 1.98173f
C902 VP.n3 B 0.04778f
C903 VP.n4 B 0.031062f
C904 VP.t0 B 1.98173f
C905 VP.n5 B 0.702506f
C906 VP.n6 B 0.031062f
C907 VP.n7 B 0.039028f
C908 VP.n8 B 0.031062f
C909 VP.t3 B 1.98173f
C910 VP.n9 B 0.050974f
C911 VP.n10 B 0.031062f
C912 VP.t9 B 1.98173f
C913 VP.n11 B 0.04778f
C914 VP.n12 B 0.031062f
C915 VP.t8 B 1.98173f
C916 VP.n13 B 0.76957f
C917 VP.t5 B 2.06354f
C918 VP.n14 B 0.773407f
C919 VP.n15 B 0.192886f
C920 VP.n16 B 0.054422f
C921 VP.n17 B 0.029808f
C922 VP.t6 B 1.98173f
C923 VP.n18 B 0.702506f
C924 VP.n19 B 0.04778f
C925 VP.n20 B 0.031062f
C926 VP.n21 B 0.031062f
C927 VP.n22 B 0.031062f
C928 VP.n23 B 0.029808f
C929 VP.n24 B 0.054422f
C930 VP.n25 B 0.702506f
C931 VP.n26 B 0.031597f
C932 VP.n27 B 0.031062f
C933 VP.n28 B 0.031062f
C934 VP.n29 B 0.031062f
C935 VP.n30 B 0.039722f
C936 VP.n31 B 0.039028f
C937 VP.n32 B 0.757728f
C938 VP.n33 B 1.69487f
C939 VP.t2 B 1.98173f
C940 VP.n34 B 0.757728f
C941 VP.n35 B 1.7172f
C942 VP.n36 B 0.031062f
C943 VP.n37 B 0.031062f
C944 VP.n38 B 0.039722f
C945 VP.n39 B 0.050974f
C946 VP.n40 B 0.031597f
C947 VP.n41 B 0.031062f
C948 VP.n42 B 0.031062f
C949 VP.n43 B 0.054422f
C950 VP.n44 B 0.029808f
C951 VP.t1 B 1.98173f
C952 VP.n45 B 0.702506f
C953 VP.n46 B 0.04778f
C954 VP.n47 B 0.031062f
C955 VP.n48 B 0.031062f
C956 VP.n49 B 0.031062f
C957 VP.n50 B 0.029808f
C958 VP.n51 B 0.054422f
C959 VP.n52 B 0.702506f
C960 VP.n53 B 0.031597f
C961 VP.n54 B 0.031062f
C962 VP.n55 B 0.031062f
C963 VP.n56 B 0.031062f
C964 VP.n57 B 0.039722f
C965 VP.n58 B 0.039028f
C966 VP.n59 B 0.757728f
C967 VP.n60 B 0.0296f
.ends

