* NGSPICE file created from diff_pair_sample_0158.ext - technology: sky130A

.subckt diff_pair_sample_0158 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=2.0097 ps=12.51 w=12.18 l=3.97
X1 VTAIL.t3 VN.t0 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=2.0097 ps=12.51 w=12.18 l=3.97
X2 VDD1.t5 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=4.7502 ps=25.14 w=12.18 l=3.97
X3 VTAIL.t9 VP.t2 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=2.0097 ps=12.51 w=12.18 l=3.97
X4 VDD1.t4 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=2.0097 ps=12.51 w=12.18 l=3.97
X5 VDD2.t4 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=2.0097 ps=12.51 w=12.18 l=3.97
X6 VDD1.t0 VP.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=4.7502 ps=25.14 w=12.18 l=3.97
X7 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=0 ps=0 w=12.18 l=3.97
X8 VTAIL.t4 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=2.0097 ps=12.51 w=12.18 l=3.97
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=4.7502 ps=25.14 w=12.18 l=3.97
X10 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0097 pd=12.51 as=4.7502 ps=25.14 w=12.18 l=3.97
X11 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=2.0097 ps=12.51 w=12.18 l=3.97
X12 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=0 ps=0 w=12.18 l=3.97
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=0 ps=0 w=12.18 l=3.97
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=0 ps=0 w=12.18 l=3.97
X15 VDD1.t2 VP.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7502 pd=25.14 as=2.0097 ps=12.51 w=12.18 l=3.97
R0 VP.n18 VP.n17 161.3
R1 VP.n19 VP.n14 161.3
R2 VP.n21 VP.n20 161.3
R3 VP.n22 VP.n13 161.3
R4 VP.n24 VP.n23 161.3
R5 VP.n25 VP.n12 161.3
R6 VP.n27 VP.n26 161.3
R7 VP.n28 VP.n11 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n61 VP.n60 161.3
R10 VP.n59 VP.n1 161.3
R11 VP.n58 VP.n57 161.3
R12 VP.n56 VP.n2 161.3
R13 VP.n55 VP.n54 161.3
R14 VP.n53 VP.n3 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n50 VP.n4 161.3
R17 VP.n49 VP.n48 161.3
R18 VP.n46 VP.n5 161.3
R19 VP.n45 VP.n44 161.3
R20 VP.n43 VP.n6 161.3
R21 VP.n42 VP.n41 161.3
R22 VP.n40 VP.n7 161.3
R23 VP.n39 VP.n38 161.3
R24 VP.n37 VP.n8 161.3
R25 VP.n36 VP.n35 161.3
R26 VP.n34 VP.n9 161.3
R27 VP.n15 VP.t3 106.707
R28 VP.n33 VP.n32 87.7864
R29 VP.n62 VP.n0 87.7864
R30 VP.n31 VP.n10 87.7864
R31 VP.n33 VP.t5 73.9395
R32 VP.n47 VP.t0 73.9395
R33 VP.n0 VP.t1 73.9395
R34 VP.n10 VP.t4 73.9395
R35 VP.n16 VP.t2 73.9395
R36 VP.n16 VP.n15 63.107
R37 VP.n32 VP.n31 54.2723
R38 VP.n41 VP.n40 50.2647
R39 VP.n54 VP.n53 50.2647
R40 VP.n23 VP.n22 50.2647
R41 VP.n40 VP.n39 30.8893
R42 VP.n54 VP.n2 30.8893
R43 VP.n23 VP.n12 30.8893
R44 VP.n35 VP.n34 24.5923
R45 VP.n35 VP.n8 24.5923
R46 VP.n39 VP.n8 24.5923
R47 VP.n41 VP.n6 24.5923
R48 VP.n45 VP.n6 24.5923
R49 VP.n46 VP.n45 24.5923
R50 VP.n48 VP.n4 24.5923
R51 VP.n52 VP.n4 24.5923
R52 VP.n53 VP.n52 24.5923
R53 VP.n58 VP.n2 24.5923
R54 VP.n59 VP.n58 24.5923
R55 VP.n60 VP.n59 24.5923
R56 VP.n27 VP.n12 24.5923
R57 VP.n28 VP.n27 24.5923
R58 VP.n29 VP.n28 24.5923
R59 VP.n17 VP.n14 24.5923
R60 VP.n21 VP.n14 24.5923
R61 VP.n22 VP.n21 24.5923
R62 VP.n47 VP.n46 12.2964
R63 VP.n48 VP.n47 12.2964
R64 VP.n17 VP.n16 12.2964
R65 VP.n18 VP.n15 2.46666
R66 VP.n34 VP.n33 2.45968
R67 VP.n60 VP.n0 2.45968
R68 VP.n29 VP.n10 2.45968
R69 VP.n31 VP.n30 0.354861
R70 VP.n32 VP.n9 0.354861
R71 VP.n62 VP.n61 0.354861
R72 VP VP.n62 0.267071
R73 VP.n19 VP.n18 0.189894
R74 VP.n20 VP.n19 0.189894
R75 VP.n20 VP.n13 0.189894
R76 VP.n24 VP.n13 0.189894
R77 VP.n25 VP.n24 0.189894
R78 VP.n26 VP.n25 0.189894
R79 VP.n26 VP.n11 0.189894
R80 VP.n30 VP.n11 0.189894
R81 VP.n36 VP.n9 0.189894
R82 VP.n37 VP.n36 0.189894
R83 VP.n38 VP.n37 0.189894
R84 VP.n38 VP.n7 0.189894
R85 VP.n42 VP.n7 0.189894
R86 VP.n43 VP.n42 0.189894
R87 VP.n44 VP.n43 0.189894
R88 VP.n44 VP.n5 0.189894
R89 VP.n49 VP.n5 0.189894
R90 VP.n50 VP.n49 0.189894
R91 VP.n51 VP.n50 0.189894
R92 VP.n51 VP.n3 0.189894
R93 VP.n55 VP.n3 0.189894
R94 VP.n56 VP.n55 0.189894
R95 VP.n57 VP.n56 0.189894
R96 VP.n57 VP.n1 0.189894
R97 VP.n61 VP.n1 0.189894
R98 VDD1.n60 VDD1.n0 289.615
R99 VDD1.n125 VDD1.n65 289.615
R100 VDD1.n61 VDD1.n60 185
R101 VDD1.n59 VDD1.n58 185
R102 VDD1.n4 VDD1.n3 185
R103 VDD1.n53 VDD1.n52 185
R104 VDD1.n51 VDD1.n50 185
R105 VDD1.n8 VDD1.n7 185
R106 VDD1.n45 VDD1.n44 185
R107 VDD1.n43 VDD1.n10 185
R108 VDD1.n42 VDD1.n41 185
R109 VDD1.n13 VDD1.n11 185
R110 VDD1.n36 VDD1.n35 185
R111 VDD1.n34 VDD1.n33 185
R112 VDD1.n17 VDD1.n16 185
R113 VDD1.n28 VDD1.n27 185
R114 VDD1.n26 VDD1.n25 185
R115 VDD1.n21 VDD1.n20 185
R116 VDD1.n85 VDD1.n84 185
R117 VDD1.n90 VDD1.n89 185
R118 VDD1.n92 VDD1.n91 185
R119 VDD1.n81 VDD1.n80 185
R120 VDD1.n98 VDD1.n97 185
R121 VDD1.n100 VDD1.n99 185
R122 VDD1.n77 VDD1.n76 185
R123 VDD1.n107 VDD1.n106 185
R124 VDD1.n108 VDD1.n75 185
R125 VDD1.n110 VDD1.n109 185
R126 VDD1.n73 VDD1.n72 185
R127 VDD1.n116 VDD1.n115 185
R128 VDD1.n118 VDD1.n117 185
R129 VDD1.n69 VDD1.n68 185
R130 VDD1.n124 VDD1.n123 185
R131 VDD1.n126 VDD1.n125 185
R132 VDD1.n22 VDD1.t4 149.524
R133 VDD1.n86 VDD1.t2 149.524
R134 VDD1.n60 VDD1.n59 104.615
R135 VDD1.n59 VDD1.n3 104.615
R136 VDD1.n52 VDD1.n3 104.615
R137 VDD1.n52 VDD1.n51 104.615
R138 VDD1.n51 VDD1.n7 104.615
R139 VDD1.n44 VDD1.n7 104.615
R140 VDD1.n44 VDD1.n43 104.615
R141 VDD1.n43 VDD1.n42 104.615
R142 VDD1.n42 VDD1.n11 104.615
R143 VDD1.n35 VDD1.n11 104.615
R144 VDD1.n35 VDD1.n34 104.615
R145 VDD1.n34 VDD1.n16 104.615
R146 VDD1.n27 VDD1.n16 104.615
R147 VDD1.n27 VDD1.n26 104.615
R148 VDD1.n26 VDD1.n20 104.615
R149 VDD1.n90 VDD1.n84 104.615
R150 VDD1.n91 VDD1.n90 104.615
R151 VDD1.n91 VDD1.n80 104.615
R152 VDD1.n98 VDD1.n80 104.615
R153 VDD1.n99 VDD1.n98 104.615
R154 VDD1.n99 VDD1.n76 104.615
R155 VDD1.n107 VDD1.n76 104.615
R156 VDD1.n108 VDD1.n107 104.615
R157 VDD1.n109 VDD1.n108 104.615
R158 VDD1.n109 VDD1.n72 104.615
R159 VDD1.n116 VDD1.n72 104.615
R160 VDD1.n117 VDD1.n116 104.615
R161 VDD1.n117 VDD1.n68 104.615
R162 VDD1.n124 VDD1.n68 104.615
R163 VDD1.n125 VDD1.n124 104.615
R164 VDD1.n131 VDD1.n130 63.9148
R165 VDD1.n133 VDD1.n132 63.0434
R166 VDD1 VDD1.n64 52.8661
R167 VDD1.n131 VDD1.n129 52.7526
R168 VDD1.t4 VDD1.n20 52.3082
R169 VDD1.t2 VDD1.n84 52.3082
R170 VDD1.n133 VDD1.n131 48.6992
R171 VDD1.n45 VDD1.n10 13.1884
R172 VDD1.n110 VDD1.n75 13.1884
R173 VDD1.n46 VDD1.n8 12.8005
R174 VDD1.n41 VDD1.n12 12.8005
R175 VDD1.n106 VDD1.n105 12.8005
R176 VDD1.n111 VDD1.n73 12.8005
R177 VDD1.n50 VDD1.n49 12.0247
R178 VDD1.n40 VDD1.n13 12.0247
R179 VDD1.n104 VDD1.n77 12.0247
R180 VDD1.n115 VDD1.n114 12.0247
R181 VDD1.n53 VDD1.n6 11.249
R182 VDD1.n37 VDD1.n36 11.249
R183 VDD1.n101 VDD1.n100 11.249
R184 VDD1.n118 VDD1.n71 11.249
R185 VDD1.n54 VDD1.n4 10.4732
R186 VDD1.n33 VDD1.n15 10.4732
R187 VDD1.n97 VDD1.n79 10.4732
R188 VDD1.n119 VDD1.n69 10.4732
R189 VDD1.n22 VDD1.n21 10.2747
R190 VDD1.n86 VDD1.n85 10.2747
R191 VDD1.n58 VDD1.n57 9.69747
R192 VDD1.n32 VDD1.n17 9.69747
R193 VDD1.n96 VDD1.n81 9.69747
R194 VDD1.n123 VDD1.n122 9.69747
R195 VDD1.n64 VDD1.n63 9.45567
R196 VDD1.n129 VDD1.n128 9.45567
R197 VDD1.n24 VDD1.n23 9.3005
R198 VDD1.n19 VDD1.n18 9.3005
R199 VDD1.n30 VDD1.n29 9.3005
R200 VDD1.n32 VDD1.n31 9.3005
R201 VDD1.n15 VDD1.n14 9.3005
R202 VDD1.n38 VDD1.n37 9.3005
R203 VDD1.n40 VDD1.n39 9.3005
R204 VDD1.n12 VDD1.n9 9.3005
R205 VDD1.n63 VDD1.n62 9.3005
R206 VDD1.n2 VDD1.n1 9.3005
R207 VDD1.n57 VDD1.n56 9.3005
R208 VDD1.n55 VDD1.n54 9.3005
R209 VDD1.n6 VDD1.n5 9.3005
R210 VDD1.n49 VDD1.n48 9.3005
R211 VDD1.n47 VDD1.n46 9.3005
R212 VDD1.n128 VDD1.n127 9.3005
R213 VDD1.n67 VDD1.n66 9.3005
R214 VDD1.n122 VDD1.n121 9.3005
R215 VDD1.n120 VDD1.n119 9.3005
R216 VDD1.n71 VDD1.n70 9.3005
R217 VDD1.n114 VDD1.n113 9.3005
R218 VDD1.n112 VDD1.n111 9.3005
R219 VDD1.n88 VDD1.n87 9.3005
R220 VDD1.n83 VDD1.n82 9.3005
R221 VDD1.n94 VDD1.n93 9.3005
R222 VDD1.n96 VDD1.n95 9.3005
R223 VDD1.n79 VDD1.n78 9.3005
R224 VDD1.n102 VDD1.n101 9.3005
R225 VDD1.n104 VDD1.n103 9.3005
R226 VDD1.n105 VDD1.n74 9.3005
R227 VDD1.n61 VDD1.n2 8.92171
R228 VDD1.n29 VDD1.n28 8.92171
R229 VDD1.n93 VDD1.n92 8.92171
R230 VDD1.n126 VDD1.n67 8.92171
R231 VDD1.n62 VDD1.n0 8.14595
R232 VDD1.n25 VDD1.n19 8.14595
R233 VDD1.n89 VDD1.n83 8.14595
R234 VDD1.n127 VDD1.n65 8.14595
R235 VDD1.n24 VDD1.n21 7.3702
R236 VDD1.n88 VDD1.n85 7.3702
R237 VDD1.n64 VDD1.n0 5.81868
R238 VDD1.n25 VDD1.n24 5.81868
R239 VDD1.n89 VDD1.n88 5.81868
R240 VDD1.n129 VDD1.n65 5.81868
R241 VDD1.n62 VDD1.n61 5.04292
R242 VDD1.n28 VDD1.n19 5.04292
R243 VDD1.n92 VDD1.n83 5.04292
R244 VDD1.n127 VDD1.n126 5.04292
R245 VDD1.n58 VDD1.n2 4.26717
R246 VDD1.n29 VDD1.n17 4.26717
R247 VDD1.n93 VDD1.n81 4.26717
R248 VDD1.n123 VDD1.n67 4.26717
R249 VDD1.n57 VDD1.n4 3.49141
R250 VDD1.n33 VDD1.n32 3.49141
R251 VDD1.n97 VDD1.n96 3.49141
R252 VDD1.n122 VDD1.n69 3.49141
R253 VDD1.n23 VDD1.n22 2.84303
R254 VDD1.n87 VDD1.n86 2.84303
R255 VDD1.n54 VDD1.n53 2.71565
R256 VDD1.n36 VDD1.n15 2.71565
R257 VDD1.n100 VDD1.n79 2.71565
R258 VDD1.n119 VDD1.n118 2.71565
R259 VDD1.n50 VDD1.n6 1.93989
R260 VDD1.n37 VDD1.n13 1.93989
R261 VDD1.n101 VDD1.n77 1.93989
R262 VDD1.n115 VDD1.n71 1.93989
R263 VDD1.n132 VDD1.t1 1.62612
R264 VDD1.n132 VDD1.t0 1.62612
R265 VDD1.n130 VDD1.t3 1.62612
R266 VDD1.n130 VDD1.t5 1.62612
R267 VDD1.n49 VDD1.n8 1.16414
R268 VDD1.n41 VDD1.n40 1.16414
R269 VDD1.n106 VDD1.n104 1.16414
R270 VDD1.n114 VDD1.n73 1.16414
R271 VDD1 VDD1.n133 0.869035
R272 VDD1.n46 VDD1.n45 0.388379
R273 VDD1.n12 VDD1.n10 0.388379
R274 VDD1.n105 VDD1.n75 0.388379
R275 VDD1.n111 VDD1.n110 0.388379
R276 VDD1.n63 VDD1.n1 0.155672
R277 VDD1.n56 VDD1.n1 0.155672
R278 VDD1.n56 VDD1.n55 0.155672
R279 VDD1.n55 VDD1.n5 0.155672
R280 VDD1.n48 VDD1.n5 0.155672
R281 VDD1.n48 VDD1.n47 0.155672
R282 VDD1.n47 VDD1.n9 0.155672
R283 VDD1.n39 VDD1.n9 0.155672
R284 VDD1.n39 VDD1.n38 0.155672
R285 VDD1.n38 VDD1.n14 0.155672
R286 VDD1.n31 VDD1.n14 0.155672
R287 VDD1.n31 VDD1.n30 0.155672
R288 VDD1.n30 VDD1.n18 0.155672
R289 VDD1.n23 VDD1.n18 0.155672
R290 VDD1.n87 VDD1.n82 0.155672
R291 VDD1.n94 VDD1.n82 0.155672
R292 VDD1.n95 VDD1.n94 0.155672
R293 VDD1.n95 VDD1.n78 0.155672
R294 VDD1.n102 VDD1.n78 0.155672
R295 VDD1.n103 VDD1.n102 0.155672
R296 VDD1.n103 VDD1.n74 0.155672
R297 VDD1.n112 VDD1.n74 0.155672
R298 VDD1.n113 VDD1.n112 0.155672
R299 VDD1.n113 VDD1.n70 0.155672
R300 VDD1.n120 VDD1.n70 0.155672
R301 VDD1.n121 VDD1.n120 0.155672
R302 VDD1.n121 VDD1.n66 0.155672
R303 VDD1.n128 VDD1.n66 0.155672
R304 VTAIL.n266 VTAIL.n206 289.615
R305 VTAIL.n62 VTAIL.n2 289.615
R306 VTAIL.n200 VTAIL.n140 289.615
R307 VTAIL.n132 VTAIL.n72 289.615
R308 VTAIL.n226 VTAIL.n225 185
R309 VTAIL.n231 VTAIL.n230 185
R310 VTAIL.n233 VTAIL.n232 185
R311 VTAIL.n222 VTAIL.n221 185
R312 VTAIL.n239 VTAIL.n238 185
R313 VTAIL.n241 VTAIL.n240 185
R314 VTAIL.n218 VTAIL.n217 185
R315 VTAIL.n248 VTAIL.n247 185
R316 VTAIL.n249 VTAIL.n216 185
R317 VTAIL.n251 VTAIL.n250 185
R318 VTAIL.n214 VTAIL.n213 185
R319 VTAIL.n257 VTAIL.n256 185
R320 VTAIL.n259 VTAIL.n258 185
R321 VTAIL.n210 VTAIL.n209 185
R322 VTAIL.n265 VTAIL.n264 185
R323 VTAIL.n267 VTAIL.n266 185
R324 VTAIL.n22 VTAIL.n21 185
R325 VTAIL.n27 VTAIL.n26 185
R326 VTAIL.n29 VTAIL.n28 185
R327 VTAIL.n18 VTAIL.n17 185
R328 VTAIL.n35 VTAIL.n34 185
R329 VTAIL.n37 VTAIL.n36 185
R330 VTAIL.n14 VTAIL.n13 185
R331 VTAIL.n44 VTAIL.n43 185
R332 VTAIL.n45 VTAIL.n12 185
R333 VTAIL.n47 VTAIL.n46 185
R334 VTAIL.n10 VTAIL.n9 185
R335 VTAIL.n53 VTAIL.n52 185
R336 VTAIL.n55 VTAIL.n54 185
R337 VTAIL.n6 VTAIL.n5 185
R338 VTAIL.n61 VTAIL.n60 185
R339 VTAIL.n63 VTAIL.n62 185
R340 VTAIL.n201 VTAIL.n200 185
R341 VTAIL.n199 VTAIL.n198 185
R342 VTAIL.n144 VTAIL.n143 185
R343 VTAIL.n193 VTAIL.n192 185
R344 VTAIL.n191 VTAIL.n190 185
R345 VTAIL.n148 VTAIL.n147 185
R346 VTAIL.n185 VTAIL.n184 185
R347 VTAIL.n183 VTAIL.n150 185
R348 VTAIL.n182 VTAIL.n181 185
R349 VTAIL.n153 VTAIL.n151 185
R350 VTAIL.n176 VTAIL.n175 185
R351 VTAIL.n174 VTAIL.n173 185
R352 VTAIL.n157 VTAIL.n156 185
R353 VTAIL.n168 VTAIL.n167 185
R354 VTAIL.n166 VTAIL.n165 185
R355 VTAIL.n161 VTAIL.n160 185
R356 VTAIL.n133 VTAIL.n132 185
R357 VTAIL.n131 VTAIL.n130 185
R358 VTAIL.n76 VTAIL.n75 185
R359 VTAIL.n125 VTAIL.n124 185
R360 VTAIL.n123 VTAIL.n122 185
R361 VTAIL.n80 VTAIL.n79 185
R362 VTAIL.n117 VTAIL.n116 185
R363 VTAIL.n115 VTAIL.n82 185
R364 VTAIL.n114 VTAIL.n113 185
R365 VTAIL.n85 VTAIL.n83 185
R366 VTAIL.n108 VTAIL.n107 185
R367 VTAIL.n106 VTAIL.n105 185
R368 VTAIL.n89 VTAIL.n88 185
R369 VTAIL.n100 VTAIL.n99 185
R370 VTAIL.n98 VTAIL.n97 185
R371 VTAIL.n93 VTAIL.n92 185
R372 VTAIL.n227 VTAIL.t1 149.524
R373 VTAIL.n23 VTAIL.t10 149.524
R374 VTAIL.n162 VTAIL.t7 149.524
R375 VTAIL.n94 VTAIL.t0 149.524
R376 VTAIL.n231 VTAIL.n225 104.615
R377 VTAIL.n232 VTAIL.n231 104.615
R378 VTAIL.n232 VTAIL.n221 104.615
R379 VTAIL.n239 VTAIL.n221 104.615
R380 VTAIL.n240 VTAIL.n239 104.615
R381 VTAIL.n240 VTAIL.n217 104.615
R382 VTAIL.n248 VTAIL.n217 104.615
R383 VTAIL.n249 VTAIL.n248 104.615
R384 VTAIL.n250 VTAIL.n249 104.615
R385 VTAIL.n250 VTAIL.n213 104.615
R386 VTAIL.n257 VTAIL.n213 104.615
R387 VTAIL.n258 VTAIL.n257 104.615
R388 VTAIL.n258 VTAIL.n209 104.615
R389 VTAIL.n265 VTAIL.n209 104.615
R390 VTAIL.n266 VTAIL.n265 104.615
R391 VTAIL.n27 VTAIL.n21 104.615
R392 VTAIL.n28 VTAIL.n27 104.615
R393 VTAIL.n28 VTAIL.n17 104.615
R394 VTAIL.n35 VTAIL.n17 104.615
R395 VTAIL.n36 VTAIL.n35 104.615
R396 VTAIL.n36 VTAIL.n13 104.615
R397 VTAIL.n44 VTAIL.n13 104.615
R398 VTAIL.n45 VTAIL.n44 104.615
R399 VTAIL.n46 VTAIL.n45 104.615
R400 VTAIL.n46 VTAIL.n9 104.615
R401 VTAIL.n53 VTAIL.n9 104.615
R402 VTAIL.n54 VTAIL.n53 104.615
R403 VTAIL.n54 VTAIL.n5 104.615
R404 VTAIL.n61 VTAIL.n5 104.615
R405 VTAIL.n62 VTAIL.n61 104.615
R406 VTAIL.n200 VTAIL.n199 104.615
R407 VTAIL.n199 VTAIL.n143 104.615
R408 VTAIL.n192 VTAIL.n143 104.615
R409 VTAIL.n192 VTAIL.n191 104.615
R410 VTAIL.n191 VTAIL.n147 104.615
R411 VTAIL.n184 VTAIL.n147 104.615
R412 VTAIL.n184 VTAIL.n183 104.615
R413 VTAIL.n183 VTAIL.n182 104.615
R414 VTAIL.n182 VTAIL.n151 104.615
R415 VTAIL.n175 VTAIL.n151 104.615
R416 VTAIL.n175 VTAIL.n174 104.615
R417 VTAIL.n174 VTAIL.n156 104.615
R418 VTAIL.n167 VTAIL.n156 104.615
R419 VTAIL.n167 VTAIL.n166 104.615
R420 VTAIL.n166 VTAIL.n160 104.615
R421 VTAIL.n132 VTAIL.n131 104.615
R422 VTAIL.n131 VTAIL.n75 104.615
R423 VTAIL.n124 VTAIL.n75 104.615
R424 VTAIL.n124 VTAIL.n123 104.615
R425 VTAIL.n123 VTAIL.n79 104.615
R426 VTAIL.n116 VTAIL.n79 104.615
R427 VTAIL.n116 VTAIL.n115 104.615
R428 VTAIL.n115 VTAIL.n114 104.615
R429 VTAIL.n114 VTAIL.n83 104.615
R430 VTAIL.n107 VTAIL.n83 104.615
R431 VTAIL.n107 VTAIL.n106 104.615
R432 VTAIL.n106 VTAIL.n88 104.615
R433 VTAIL.n99 VTAIL.n88 104.615
R434 VTAIL.n99 VTAIL.n98 104.615
R435 VTAIL.n98 VTAIL.n92 104.615
R436 VTAIL.t1 VTAIL.n225 52.3082
R437 VTAIL.t10 VTAIL.n21 52.3082
R438 VTAIL.t7 VTAIL.n160 52.3082
R439 VTAIL.t0 VTAIL.n92 52.3082
R440 VTAIL.n139 VTAIL.n138 46.3648
R441 VTAIL.n71 VTAIL.n70 46.3648
R442 VTAIL.n1 VTAIL.n0 46.3646
R443 VTAIL.n69 VTAIL.n68 46.3646
R444 VTAIL.n271 VTAIL.n270 33.349
R445 VTAIL.n67 VTAIL.n66 33.349
R446 VTAIL.n205 VTAIL.n204 33.349
R447 VTAIL.n137 VTAIL.n136 33.349
R448 VTAIL.n71 VTAIL.n69 30.2807
R449 VTAIL.n271 VTAIL.n205 26.5738
R450 VTAIL.n251 VTAIL.n216 13.1884
R451 VTAIL.n47 VTAIL.n12 13.1884
R452 VTAIL.n185 VTAIL.n150 13.1884
R453 VTAIL.n117 VTAIL.n82 13.1884
R454 VTAIL.n247 VTAIL.n246 12.8005
R455 VTAIL.n252 VTAIL.n214 12.8005
R456 VTAIL.n43 VTAIL.n42 12.8005
R457 VTAIL.n48 VTAIL.n10 12.8005
R458 VTAIL.n186 VTAIL.n148 12.8005
R459 VTAIL.n181 VTAIL.n152 12.8005
R460 VTAIL.n118 VTAIL.n80 12.8005
R461 VTAIL.n113 VTAIL.n84 12.8005
R462 VTAIL.n245 VTAIL.n218 12.0247
R463 VTAIL.n256 VTAIL.n255 12.0247
R464 VTAIL.n41 VTAIL.n14 12.0247
R465 VTAIL.n52 VTAIL.n51 12.0247
R466 VTAIL.n190 VTAIL.n189 12.0247
R467 VTAIL.n180 VTAIL.n153 12.0247
R468 VTAIL.n122 VTAIL.n121 12.0247
R469 VTAIL.n112 VTAIL.n85 12.0247
R470 VTAIL.n242 VTAIL.n241 11.249
R471 VTAIL.n259 VTAIL.n212 11.249
R472 VTAIL.n38 VTAIL.n37 11.249
R473 VTAIL.n55 VTAIL.n8 11.249
R474 VTAIL.n193 VTAIL.n146 11.249
R475 VTAIL.n177 VTAIL.n176 11.249
R476 VTAIL.n125 VTAIL.n78 11.249
R477 VTAIL.n109 VTAIL.n108 11.249
R478 VTAIL.n238 VTAIL.n220 10.4732
R479 VTAIL.n260 VTAIL.n210 10.4732
R480 VTAIL.n34 VTAIL.n16 10.4732
R481 VTAIL.n56 VTAIL.n6 10.4732
R482 VTAIL.n194 VTAIL.n144 10.4732
R483 VTAIL.n173 VTAIL.n155 10.4732
R484 VTAIL.n126 VTAIL.n76 10.4732
R485 VTAIL.n105 VTAIL.n87 10.4732
R486 VTAIL.n227 VTAIL.n226 10.2747
R487 VTAIL.n23 VTAIL.n22 10.2747
R488 VTAIL.n162 VTAIL.n161 10.2747
R489 VTAIL.n94 VTAIL.n93 10.2747
R490 VTAIL.n237 VTAIL.n222 9.69747
R491 VTAIL.n264 VTAIL.n263 9.69747
R492 VTAIL.n33 VTAIL.n18 9.69747
R493 VTAIL.n60 VTAIL.n59 9.69747
R494 VTAIL.n198 VTAIL.n197 9.69747
R495 VTAIL.n172 VTAIL.n157 9.69747
R496 VTAIL.n130 VTAIL.n129 9.69747
R497 VTAIL.n104 VTAIL.n89 9.69747
R498 VTAIL.n270 VTAIL.n269 9.45567
R499 VTAIL.n66 VTAIL.n65 9.45567
R500 VTAIL.n204 VTAIL.n203 9.45567
R501 VTAIL.n136 VTAIL.n135 9.45567
R502 VTAIL.n269 VTAIL.n268 9.3005
R503 VTAIL.n208 VTAIL.n207 9.3005
R504 VTAIL.n263 VTAIL.n262 9.3005
R505 VTAIL.n261 VTAIL.n260 9.3005
R506 VTAIL.n212 VTAIL.n211 9.3005
R507 VTAIL.n255 VTAIL.n254 9.3005
R508 VTAIL.n253 VTAIL.n252 9.3005
R509 VTAIL.n229 VTAIL.n228 9.3005
R510 VTAIL.n224 VTAIL.n223 9.3005
R511 VTAIL.n235 VTAIL.n234 9.3005
R512 VTAIL.n237 VTAIL.n236 9.3005
R513 VTAIL.n220 VTAIL.n219 9.3005
R514 VTAIL.n243 VTAIL.n242 9.3005
R515 VTAIL.n245 VTAIL.n244 9.3005
R516 VTAIL.n246 VTAIL.n215 9.3005
R517 VTAIL.n65 VTAIL.n64 9.3005
R518 VTAIL.n4 VTAIL.n3 9.3005
R519 VTAIL.n59 VTAIL.n58 9.3005
R520 VTAIL.n57 VTAIL.n56 9.3005
R521 VTAIL.n8 VTAIL.n7 9.3005
R522 VTAIL.n51 VTAIL.n50 9.3005
R523 VTAIL.n49 VTAIL.n48 9.3005
R524 VTAIL.n25 VTAIL.n24 9.3005
R525 VTAIL.n20 VTAIL.n19 9.3005
R526 VTAIL.n31 VTAIL.n30 9.3005
R527 VTAIL.n33 VTAIL.n32 9.3005
R528 VTAIL.n16 VTAIL.n15 9.3005
R529 VTAIL.n39 VTAIL.n38 9.3005
R530 VTAIL.n41 VTAIL.n40 9.3005
R531 VTAIL.n42 VTAIL.n11 9.3005
R532 VTAIL.n164 VTAIL.n163 9.3005
R533 VTAIL.n159 VTAIL.n158 9.3005
R534 VTAIL.n170 VTAIL.n169 9.3005
R535 VTAIL.n172 VTAIL.n171 9.3005
R536 VTAIL.n155 VTAIL.n154 9.3005
R537 VTAIL.n178 VTAIL.n177 9.3005
R538 VTAIL.n180 VTAIL.n179 9.3005
R539 VTAIL.n152 VTAIL.n149 9.3005
R540 VTAIL.n203 VTAIL.n202 9.3005
R541 VTAIL.n142 VTAIL.n141 9.3005
R542 VTAIL.n197 VTAIL.n196 9.3005
R543 VTAIL.n195 VTAIL.n194 9.3005
R544 VTAIL.n146 VTAIL.n145 9.3005
R545 VTAIL.n189 VTAIL.n188 9.3005
R546 VTAIL.n187 VTAIL.n186 9.3005
R547 VTAIL.n96 VTAIL.n95 9.3005
R548 VTAIL.n91 VTAIL.n90 9.3005
R549 VTAIL.n102 VTAIL.n101 9.3005
R550 VTAIL.n104 VTAIL.n103 9.3005
R551 VTAIL.n87 VTAIL.n86 9.3005
R552 VTAIL.n110 VTAIL.n109 9.3005
R553 VTAIL.n112 VTAIL.n111 9.3005
R554 VTAIL.n84 VTAIL.n81 9.3005
R555 VTAIL.n135 VTAIL.n134 9.3005
R556 VTAIL.n74 VTAIL.n73 9.3005
R557 VTAIL.n129 VTAIL.n128 9.3005
R558 VTAIL.n127 VTAIL.n126 9.3005
R559 VTAIL.n78 VTAIL.n77 9.3005
R560 VTAIL.n121 VTAIL.n120 9.3005
R561 VTAIL.n119 VTAIL.n118 9.3005
R562 VTAIL.n234 VTAIL.n233 8.92171
R563 VTAIL.n267 VTAIL.n208 8.92171
R564 VTAIL.n30 VTAIL.n29 8.92171
R565 VTAIL.n63 VTAIL.n4 8.92171
R566 VTAIL.n201 VTAIL.n142 8.92171
R567 VTAIL.n169 VTAIL.n168 8.92171
R568 VTAIL.n133 VTAIL.n74 8.92171
R569 VTAIL.n101 VTAIL.n100 8.92171
R570 VTAIL.n230 VTAIL.n224 8.14595
R571 VTAIL.n268 VTAIL.n206 8.14595
R572 VTAIL.n26 VTAIL.n20 8.14595
R573 VTAIL.n64 VTAIL.n2 8.14595
R574 VTAIL.n202 VTAIL.n140 8.14595
R575 VTAIL.n165 VTAIL.n159 8.14595
R576 VTAIL.n134 VTAIL.n72 8.14595
R577 VTAIL.n97 VTAIL.n91 8.14595
R578 VTAIL.n229 VTAIL.n226 7.3702
R579 VTAIL.n25 VTAIL.n22 7.3702
R580 VTAIL.n164 VTAIL.n161 7.3702
R581 VTAIL.n96 VTAIL.n93 7.3702
R582 VTAIL.n230 VTAIL.n229 5.81868
R583 VTAIL.n270 VTAIL.n206 5.81868
R584 VTAIL.n26 VTAIL.n25 5.81868
R585 VTAIL.n66 VTAIL.n2 5.81868
R586 VTAIL.n204 VTAIL.n140 5.81868
R587 VTAIL.n165 VTAIL.n164 5.81868
R588 VTAIL.n136 VTAIL.n72 5.81868
R589 VTAIL.n97 VTAIL.n96 5.81868
R590 VTAIL.n233 VTAIL.n224 5.04292
R591 VTAIL.n268 VTAIL.n267 5.04292
R592 VTAIL.n29 VTAIL.n20 5.04292
R593 VTAIL.n64 VTAIL.n63 5.04292
R594 VTAIL.n202 VTAIL.n201 5.04292
R595 VTAIL.n168 VTAIL.n159 5.04292
R596 VTAIL.n134 VTAIL.n133 5.04292
R597 VTAIL.n100 VTAIL.n91 5.04292
R598 VTAIL.n234 VTAIL.n222 4.26717
R599 VTAIL.n264 VTAIL.n208 4.26717
R600 VTAIL.n30 VTAIL.n18 4.26717
R601 VTAIL.n60 VTAIL.n4 4.26717
R602 VTAIL.n198 VTAIL.n142 4.26717
R603 VTAIL.n169 VTAIL.n157 4.26717
R604 VTAIL.n130 VTAIL.n74 4.26717
R605 VTAIL.n101 VTAIL.n89 4.26717
R606 VTAIL.n137 VTAIL.n71 3.7074
R607 VTAIL.n205 VTAIL.n139 3.7074
R608 VTAIL.n69 VTAIL.n67 3.7074
R609 VTAIL.n238 VTAIL.n237 3.49141
R610 VTAIL.n263 VTAIL.n210 3.49141
R611 VTAIL.n34 VTAIL.n33 3.49141
R612 VTAIL.n59 VTAIL.n6 3.49141
R613 VTAIL.n197 VTAIL.n144 3.49141
R614 VTAIL.n173 VTAIL.n172 3.49141
R615 VTAIL.n129 VTAIL.n76 3.49141
R616 VTAIL.n105 VTAIL.n104 3.49141
R617 VTAIL.n228 VTAIL.n227 2.84303
R618 VTAIL.n24 VTAIL.n23 2.84303
R619 VTAIL.n163 VTAIL.n162 2.84303
R620 VTAIL.n95 VTAIL.n94 2.84303
R621 VTAIL VTAIL.n271 2.72248
R622 VTAIL.n241 VTAIL.n220 2.71565
R623 VTAIL.n260 VTAIL.n259 2.71565
R624 VTAIL.n37 VTAIL.n16 2.71565
R625 VTAIL.n56 VTAIL.n55 2.71565
R626 VTAIL.n194 VTAIL.n193 2.71565
R627 VTAIL.n176 VTAIL.n155 2.71565
R628 VTAIL.n126 VTAIL.n125 2.71565
R629 VTAIL.n108 VTAIL.n87 2.71565
R630 VTAIL.n139 VTAIL.n137 2.32378
R631 VTAIL.n67 VTAIL.n1 2.32378
R632 VTAIL.n242 VTAIL.n218 1.93989
R633 VTAIL.n256 VTAIL.n212 1.93989
R634 VTAIL.n38 VTAIL.n14 1.93989
R635 VTAIL.n52 VTAIL.n8 1.93989
R636 VTAIL.n190 VTAIL.n146 1.93989
R637 VTAIL.n177 VTAIL.n153 1.93989
R638 VTAIL.n122 VTAIL.n78 1.93989
R639 VTAIL.n109 VTAIL.n85 1.93989
R640 VTAIL.n0 VTAIL.t2 1.62612
R641 VTAIL.n0 VTAIL.t4 1.62612
R642 VTAIL.n68 VTAIL.t6 1.62612
R643 VTAIL.n68 VTAIL.t11 1.62612
R644 VTAIL.n138 VTAIL.t8 1.62612
R645 VTAIL.n138 VTAIL.t9 1.62612
R646 VTAIL.n70 VTAIL.t5 1.62612
R647 VTAIL.n70 VTAIL.t3 1.62612
R648 VTAIL.n247 VTAIL.n245 1.16414
R649 VTAIL.n255 VTAIL.n214 1.16414
R650 VTAIL.n43 VTAIL.n41 1.16414
R651 VTAIL.n51 VTAIL.n10 1.16414
R652 VTAIL.n189 VTAIL.n148 1.16414
R653 VTAIL.n181 VTAIL.n180 1.16414
R654 VTAIL.n121 VTAIL.n80 1.16414
R655 VTAIL.n113 VTAIL.n112 1.16414
R656 VTAIL VTAIL.n1 0.985414
R657 VTAIL.n246 VTAIL.n216 0.388379
R658 VTAIL.n252 VTAIL.n251 0.388379
R659 VTAIL.n42 VTAIL.n12 0.388379
R660 VTAIL.n48 VTAIL.n47 0.388379
R661 VTAIL.n186 VTAIL.n185 0.388379
R662 VTAIL.n152 VTAIL.n150 0.388379
R663 VTAIL.n118 VTAIL.n117 0.388379
R664 VTAIL.n84 VTAIL.n82 0.388379
R665 VTAIL.n228 VTAIL.n223 0.155672
R666 VTAIL.n235 VTAIL.n223 0.155672
R667 VTAIL.n236 VTAIL.n235 0.155672
R668 VTAIL.n236 VTAIL.n219 0.155672
R669 VTAIL.n243 VTAIL.n219 0.155672
R670 VTAIL.n244 VTAIL.n243 0.155672
R671 VTAIL.n244 VTAIL.n215 0.155672
R672 VTAIL.n253 VTAIL.n215 0.155672
R673 VTAIL.n254 VTAIL.n253 0.155672
R674 VTAIL.n254 VTAIL.n211 0.155672
R675 VTAIL.n261 VTAIL.n211 0.155672
R676 VTAIL.n262 VTAIL.n261 0.155672
R677 VTAIL.n262 VTAIL.n207 0.155672
R678 VTAIL.n269 VTAIL.n207 0.155672
R679 VTAIL.n24 VTAIL.n19 0.155672
R680 VTAIL.n31 VTAIL.n19 0.155672
R681 VTAIL.n32 VTAIL.n31 0.155672
R682 VTAIL.n32 VTAIL.n15 0.155672
R683 VTAIL.n39 VTAIL.n15 0.155672
R684 VTAIL.n40 VTAIL.n39 0.155672
R685 VTAIL.n40 VTAIL.n11 0.155672
R686 VTAIL.n49 VTAIL.n11 0.155672
R687 VTAIL.n50 VTAIL.n49 0.155672
R688 VTAIL.n50 VTAIL.n7 0.155672
R689 VTAIL.n57 VTAIL.n7 0.155672
R690 VTAIL.n58 VTAIL.n57 0.155672
R691 VTAIL.n58 VTAIL.n3 0.155672
R692 VTAIL.n65 VTAIL.n3 0.155672
R693 VTAIL.n203 VTAIL.n141 0.155672
R694 VTAIL.n196 VTAIL.n141 0.155672
R695 VTAIL.n196 VTAIL.n195 0.155672
R696 VTAIL.n195 VTAIL.n145 0.155672
R697 VTAIL.n188 VTAIL.n145 0.155672
R698 VTAIL.n188 VTAIL.n187 0.155672
R699 VTAIL.n187 VTAIL.n149 0.155672
R700 VTAIL.n179 VTAIL.n149 0.155672
R701 VTAIL.n179 VTAIL.n178 0.155672
R702 VTAIL.n178 VTAIL.n154 0.155672
R703 VTAIL.n171 VTAIL.n154 0.155672
R704 VTAIL.n171 VTAIL.n170 0.155672
R705 VTAIL.n170 VTAIL.n158 0.155672
R706 VTAIL.n163 VTAIL.n158 0.155672
R707 VTAIL.n135 VTAIL.n73 0.155672
R708 VTAIL.n128 VTAIL.n73 0.155672
R709 VTAIL.n128 VTAIL.n127 0.155672
R710 VTAIL.n127 VTAIL.n77 0.155672
R711 VTAIL.n120 VTAIL.n77 0.155672
R712 VTAIL.n120 VTAIL.n119 0.155672
R713 VTAIL.n119 VTAIL.n81 0.155672
R714 VTAIL.n111 VTAIL.n81 0.155672
R715 VTAIL.n111 VTAIL.n110 0.155672
R716 VTAIL.n110 VTAIL.n86 0.155672
R717 VTAIL.n103 VTAIL.n86 0.155672
R718 VTAIL.n103 VTAIL.n102 0.155672
R719 VTAIL.n102 VTAIL.n90 0.155672
R720 VTAIL.n95 VTAIL.n90 0.155672
R721 B.n766 B.n765 585
R722 B.n767 B.n160 585
R723 B.n769 B.n768 585
R724 B.n771 B.n159 585
R725 B.n774 B.n773 585
R726 B.n775 B.n158 585
R727 B.n777 B.n776 585
R728 B.n779 B.n157 585
R729 B.n782 B.n781 585
R730 B.n783 B.n156 585
R731 B.n785 B.n784 585
R732 B.n787 B.n155 585
R733 B.n790 B.n789 585
R734 B.n791 B.n154 585
R735 B.n793 B.n792 585
R736 B.n795 B.n153 585
R737 B.n798 B.n797 585
R738 B.n799 B.n152 585
R739 B.n801 B.n800 585
R740 B.n803 B.n151 585
R741 B.n806 B.n805 585
R742 B.n807 B.n150 585
R743 B.n809 B.n808 585
R744 B.n811 B.n149 585
R745 B.n814 B.n813 585
R746 B.n815 B.n148 585
R747 B.n817 B.n816 585
R748 B.n819 B.n147 585
R749 B.n822 B.n821 585
R750 B.n823 B.n146 585
R751 B.n825 B.n824 585
R752 B.n827 B.n145 585
R753 B.n830 B.n829 585
R754 B.n831 B.n144 585
R755 B.n833 B.n832 585
R756 B.n835 B.n143 585
R757 B.n838 B.n837 585
R758 B.n839 B.n142 585
R759 B.n841 B.n840 585
R760 B.n843 B.n141 585
R761 B.n845 B.n844 585
R762 B.n847 B.n846 585
R763 B.n850 B.n849 585
R764 B.n851 B.n136 585
R765 B.n853 B.n852 585
R766 B.n855 B.n135 585
R767 B.n858 B.n857 585
R768 B.n859 B.n134 585
R769 B.n861 B.n860 585
R770 B.n863 B.n133 585
R771 B.n865 B.n864 585
R772 B.n867 B.n866 585
R773 B.n870 B.n869 585
R774 B.n871 B.n128 585
R775 B.n873 B.n872 585
R776 B.n875 B.n127 585
R777 B.n878 B.n877 585
R778 B.n879 B.n126 585
R779 B.n881 B.n880 585
R780 B.n883 B.n125 585
R781 B.n886 B.n885 585
R782 B.n887 B.n124 585
R783 B.n889 B.n888 585
R784 B.n891 B.n123 585
R785 B.n894 B.n893 585
R786 B.n895 B.n122 585
R787 B.n897 B.n896 585
R788 B.n899 B.n121 585
R789 B.n902 B.n901 585
R790 B.n903 B.n120 585
R791 B.n905 B.n904 585
R792 B.n907 B.n119 585
R793 B.n910 B.n909 585
R794 B.n911 B.n118 585
R795 B.n913 B.n912 585
R796 B.n915 B.n117 585
R797 B.n918 B.n917 585
R798 B.n919 B.n116 585
R799 B.n921 B.n920 585
R800 B.n923 B.n115 585
R801 B.n926 B.n925 585
R802 B.n927 B.n114 585
R803 B.n929 B.n928 585
R804 B.n931 B.n113 585
R805 B.n934 B.n933 585
R806 B.n935 B.n112 585
R807 B.n937 B.n936 585
R808 B.n939 B.n111 585
R809 B.n942 B.n941 585
R810 B.n943 B.n110 585
R811 B.n945 B.n944 585
R812 B.n947 B.n109 585
R813 B.n950 B.n949 585
R814 B.n951 B.n108 585
R815 B.n763 B.n106 585
R816 B.n954 B.n106 585
R817 B.n762 B.n105 585
R818 B.n955 B.n105 585
R819 B.n761 B.n104 585
R820 B.n956 B.n104 585
R821 B.n760 B.n759 585
R822 B.n759 B.n100 585
R823 B.n758 B.n99 585
R824 B.n962 B.n99 585
R825 B.n757 B.n98 585
R826 B.n963 B.n98 585
R827 B.n756 B.n97 585
R828 B.n964 B.n97 585
R829 B.n755 B.n754 585
R830 B.n754 B.n93 585
R831 B.n753 B.n92 585
R832 B.n970 B.n92 585
R833 B.n752 B.n91 585
R834 B.n971 B.n91 585
R835 B.n751 B.n90 585
R836 B.n972 B.n90 585
R837 B.n750 B.n749 585
R838 B.n749 B.n86 585
R839 B.n748 B.n85 585
R840 B.n978 B.n85 585
R841 B.n747 B.n84 585
R842 B.n979 B.n84 585
R843 B.n746 B.n83 585
R844 B.n980 B.n83 585
R845 B.n745 B.n744 585
R846 B.n744 B.n79 585
R847 B.n743 B.n78 585
R848 B.n986 B.n78 585
R849 B.n742 B.n77 585
R850 B.n987 B.n77 585
R851 B.n741 B.n76 585
R852 B.n988 B.n76 585
R853 B.n740 B.n739 585
R854 B.n739 B.n72 585
R855 B.n738 B.n71 585
R856 B.n994 B.n71 585
R857 B.n737 B.n70 585
R858 B.n995 B.n70 585
R859 B.n736 B.n69 585
R860 B.n996 B.n69 585
R861 B.n735 B.n734 585
R862 B.n734 B.n65 585
R863 B.n733 B.n64 585
R864 B.n1002 B.n64 585
R865 B.n732 B.n63 585
R866 B.n1003 B.n63 585
R867 B.n731 B.n62 585
R868 B.n1004 B.n62 585
R869 B.n730 B.n729 585
R870 B.n729 B.n58 585
R871 B.n728 B.n57 585
R872 B.n1010 B.n57 585
R873 B.n727 B.n56 585
R874 B.n1011 B.n56 585
R875 B.n726 B.n55 585
R876 B.n1012 B.n55 585
R877 B.n725 B.n724 585
R878 B.n724 B.n51 585
R879 B.n723 B.n50 585
R880 B.n1018 B.n50 585
R881 B.n722 B.n49 585
R882 B.n1019 B.n49 585
R883 B.n721 B.n48 585
R884 B.n1020 B.n48 585
R885 B.n720 B.n719 585
R886 B.n719 B.n44 585
R887 B.n718 B.n43 585
R888 B.n1026 B.n43 585
R889 B.n717 B.n42 585
R890 B.n1027 B.n42 585
R891 B.n716 B.n41 585
R892 B.n1028 B.n41 585
R893 B.n715 B.n714 585
R894 B.n714 B.n37 585
R895 B.n713 B.n36 585
R896 B.n1034 B.n36 585
R897 B.n712 B.n35 585
R898 B.n1035 B.n35 585
R899 B.n711 B.n34 585
R900 B.n1036 B.n34 585
R901 B.n710 B.n709 585
R902 B.n709 B.n30 585
R903 B.n708 B.n29 585
R904 B.n1042 B.n29 585
R905 B.n707 B.n28 585
R906 B.n1043 B.n28 585
R907 B.n706 B.n27 585
R908 B.n1044 B.n27 585
R909 B.n705 B.n704 585
R910 B.n704 B.n23 585
R911 B.n703 B.n22 585
R912 B.n1050 B.n22 585
R913 B.n702 B.n21 585
R914 B.n1051 B.n21 585
R915 B.n701 B.n20 585
R916 B.n1052 B.n20 585
R917 B.n700 B.n699 585
R918 B.n699 B.n16 585
R919 B.n698 B.n15 585
R920 B.n1058 B.n15 585
R921 B.n697 B.n14 585
R922 B.n1059 B.n14 585
R923 B.n696 B.n13 585
R924 B.n1060 B.n13 585
R925 B.n695 B.n694 585
R926 B.n694 B.n12 585
R927 B.n693 B.n692 585
R928 B.n693 B.n8 585
R929 B.n691 B.n7 585
R930 B.n1067 B.n7 585
R931 B.n690 B.n6 585
R932 B.n1068 B.n6 585
R933 B.n689 B.n5 585
R934 B.n1069 B.n5 585
R935 B.n688 B.n687 585
R936 B.n687 B.n4 585
R937 B.n686 B.n161 585
R938 B.n686 B.n685 585
R939 B.n676 B.n162 585
R940 B.n163 B.n162 585
R941 B.n678 B.n677 585
R942 B.n679 B.n678 585
R943 B.n675 B.n168 585
R944 B.n168 B.n167 585
R945 B.n674 B.n673 585
R946 B.n673 B.n672 585
R947 B.n170 B.n169 585
R948 B.n171 B.n170 585
R949 B.n665 B.n664 585
R950 B.n666 B.n665 585
R951 B.n663 B.n176 585
R952 B.n176 B.n175 585
R953 B.n662 B.n661 585
R954 B.n661 B.n660 585
R955 B.n178 B.n177 585
R956 B.n179 B.n178 585
R957 B.n653 B.n652 585
R958 B.n654 B.n653 585
R959 B.n651 B.n184 585
R960 B.n184 B.n183 585
R961 B.n650 B.n649 585
R962 B.n649 B.n648 585
R963 B.n186 B.n185 585
R964 B.n187 B.n186 585
R965 B.n641 B.n640 585
R966 B.n642 B.n641 585
R967 B.n639 B.n192 585
R968 B.n192 B.n191 585
R969 B.n638 B.n637 585
R970 B.n637 B.n636 585
R971 B.n194 B.n193 585
R972 B.n195 B.n194 585
R973 B.n629 B.n628 585
R974 B.n630 B.n629 585
R975 B.n627 B.n199 585
R976 B.n203 B.n199 585
R977 B.n626 B.n625 585
R978 B.n625 B.n624 585
R979 B.n201 B.n200 585
R980 B.n202 B.n201 585
R981 B.n617 B.n616 585
R982 B.n618 B.n617 585
R983 B.n615 B.n208 585
R984 B.n208 B.n207 585
R985 B.n614 B.n613 585
R986 B.n613 B.n612 585
R987 B.n210 B.n209 585
R988 B.n211 B.n210 585
R989 B.n605 B.n604 585
R990 B.n606 B.n605 585
R991 B.n603 B.n216 585
R992 B.n216 B.n215 585
R993 B.n602 B.n601 585
R994 B.n601 B.n600 585
R995 B.n218 B.n217 585
R996 B.n219 B.n218 585
R997 B.n593 B.n592 585
R998 B.n594 B.n593 585
R999 B.n591 B.n223 585
R1000 B.n227 B.n223 585
R1001 B.n590 B.n589 585
R1002 B.n589 B.n588 585
R1003 B.n225 B.n224 585
R1004 B.n226 B.n225 585
R1005 B.n581 B.n580 585
R1006 B.n582 B.n581 585
R1007 B.n579 B.n232 585
R1008 B.n232 B.n231 585
R1009 B.n578 B.n577 585
R1010 B.n577 B.n576 585
R1011 B.n234 B.n233 585
R1012 B.n235 B.n234 585
R1013 B.n569 B.n568 585
R1014 B.n570 B.n569 585
R1015 B.n567 B.n240 585
R1016 B.n240 B.n239 585
R1017 B.n566 B.n565 585
R1018 B.n565 B.n564 585
R1019 B.n242 B.n241 585
R1020 B.n243 B.n242 585
R1021 B.n557 B.n556 585
R1022 B.n558 B.n557 585
R1023 B.n555 B.n248 585
R1024 B.n248 B.n247 585
R1025 B.n554 B.n553 585
R1026 B.n553 B.n552 585
R1027 B.n250 B.n249 585
R1028 B.n251 B.n250 585
R1029 B.n545 B.n544 585
R1030 B.n546 B.n545 585
R1031 B.n543 B.n255 585
R1032 B.n259 B.n255 585
R1033 B.n542 B.n541 585
R1034 B.n541 B.n540 585
R1035 B.n257 B.n256 585
R1036 B.n258 B.n257 585
R1037 B.n533 B.n532 585
R1038 B.n534 B.n533 585
R1039 B.n531 B.n264 585
R1040 B.n264 B.n263 585
R1041 B.n530 B.n529 585
R1042 B.n529 B.n528 585
R1043 B.n266 B.n265 585
R1044 B.n267 B.n266 585
R1045 B.n521 B.n520 585
R1046 B.n522 B.n521 585
R1047 B.n519 B.n272 585
R1048 B.n272 B.n271 585
R1049 B.n518 B.n517 585
R1050 B.n517 B.n516 585
R1051 B.n513 B.n276 585
R1052 B.n512 B.n511 585
R1053 B.n509 B.n277 585
R1054 B.n509 B.n275 585
R1055 B.n508 B.n507 585
R1056 B.n506 B.n505 585
R1057 B.n504 B.n279 585
R1058 B.n502 B.n501 585
R1059 B.n500 B.n280 585
R1060 B.n499 B.n498 585
R1061 B.n496 B.n281 585
R1062 B.n494 B.n493 585
R1063 B.n492 B.n282 585
R1064 B.n491 B.n490 585
R1065 B.n488 B.n283 585
R1066 B.n486 B.n485 585
R1067 B.n484 B.n284 585
R1068 B.n483 B.n482 585
R1069 B.n480 B.n285 585
R1070 B.n478 B.n477 585
R1071 B.n476 B.n286 585
R1072 B.n475 B.n474 585
R1073 B.n472 B.n287 585
R1074 B.n470 B.n469 585
R1075 B.n468 B.n288 585
R1076 B.n467 B.n466 585
R1077 B.n464 B.n289 585
R1078 B.n462 B.n461 585
R1079 B.n460 B.n290 585
R1080 B.n459 B.n458 585
R1081 B.n456 B.n291 585
R1082 B.n454 B.n453 585
R1083 B.n452 B.n292 585
R1084 B.n451 B.n450 585
R1085 B.n448 B.n293 585
R1086 B.n446 B.n445 585
R1087 B.n444 B.n294 585
R1088 B.n443 B.n442 585
R1089 B.n440 B.n295 585
R1090 B.n438 B.n437 585
R1091 B.n436 B.n296 585
R1092 B.n435 B.n434 585
R1093 B.n432 B.n297 585
R1094 B.n430 B.n429 585
R1095 B.n428 B.n298 585
R1096 B.n427 B.n426 585
R1097 B.n424 B.n302 585
R1098 B.n422 B.n421 585
R1099 B.n420 B.n303 585
R1100 B.n419 B.n418 585
R1101 B.n416 B.n304 585
R1102 B.n414 B.n413 585
R1103 B.n412 B.n305 585
R1104 B.n410 B.n409 585
R1105 B.n407 B.n308 585
R1106 B.n405 B.n404 585
R1107 B.n403 B.n309 585
R1108 B.n402 B.n401 585
R1109 B.n399 B.n310 585
R1110 B.n397 B.n396 585
R1111 B.n395 B.n311 585
R1112 B.n394 B.n393 585
R1113 B.n391 B.n312 585
R1114 B.n389 B.n388 585
R1115 B.n387 B.n313 585
R1116 B.n386 B.n385 585
R1117 B.n383 B.n314 585
R1118 B.n381 B.n380 585
R1119 B.n379 B.n315 585
R1120 B.n378 B.n377 585
R1121 B.n375 B.n316 585
R1122 B.n373 B.n372 585
R1123 B.n371 B.n317 585
R1124 B.n370 B.n369 585
R1125 B.n367 B.n318 585
R1126 B.n365 B.n364 585
R1127 B.n363 B.n319 585
R1128 B.n362 B.n361 585
R1129 B.n359 B.n320 585
R1130 B.n357 B.n356 585
R1131 B.n355 B.n321 585
R1132 B.n354 B.n353 585
R1133 B.n351 B.n322 585
R1134 B.n349 B.n348 585
R1135 B.n347 B.n323 585
R1136 B.n346 B.n345 585
R1137 B.n343 B.n324 585
R1138 B.n341 B.n340 585
R1139 B.n339 B.n325 585
R1140 B.n338 B.n337 585
R1141 B.n335 B.n326 585
R1142 B.n333 B.n332 585
R1143 B.n331 B.n327 585
R1144 B.n330 B.n329 585
R1145 B.n274 B.n273 585
R1146 B.n275 B.n274 585
R1147 B.n515 B.n514 585
R1148 B.n516 B.n515 585
R1149 B.n270 B.n269 585
R1150 B.n271 B.n270 585
R1151 B.n524 B.n523 585
R1152 B.n523 B.n522 585
R1153 B.n525 B.n268 585
R1154 B.n268 B.n267 585
R1155 B.n527 B.n526 585
R1156 B.n528 B.n527 585
R1157 B.n262 B.n261 585
R1158 B.n263 B.n262 585
R1159 B.n536 B.n535 585
R1160 B.n535 B.n534 585
R1161 B.n537 B.n260 585
R1162 B.n260 B.n258 585
R1163 B.n539 B.n538 585
R1164 B.n540 B.n539 585
R1165 B.n254 B.n253 585
R1166 B.n259 B.n254 585
R1167 B.n548 B.n547 585
R1168 B.n547 B.n546 585
R1169 B.n549 B.n252 585
R1170 B.n252 B.n251 585
R1171 B.n551 B.n550 585
R1172 B.n552 B.n551 585
R1173 B.n246 B.n245 585
R1174 B.n247 B.n246 585
R1175 B.n560 B.n559 585
R1176 B.n559 B.n558 585
R1177 B.n561 B.n244 585
R1178 B.n244 B.n243 585
R1179 B.n563 B.n562 585
R1180 B.n564 B.n563 585
R1181 B.n238 B.n237 585
R1182 B.n239 B.n238 585
R1183 B.n572 B.n571 585
R1184 B.n571 B.n570 585
R1185 B.n573 B.n236 585
R1186 B.n236 B.n235 585
R1187 B.n575 B.n574 585
R1188 B.n576 B.n575 585
R1189 B.n230 B.n229 585
R1190 B.n231 B.n230 585
R1191 B.n584 B.n583 585
R1192 B.n583 B.n582 585
R1193 B.n585 B.n228 585
R1194 B.n228 B.n226 585
R1195 B.n587 B.n586 585
R1196 B.n588 B.n587 585
R1197 B.n222 B.n221 585
R1198 B.n227 B.n222 585
R1199 B.n596 B.n595 585
R1200 B.n595 B.n594 585
R1201 B.n597 B.n220 585
R1202 B.n220 B.n219 585
R1203 B.n599 B.n598 585
R1204 B.n600 B.n599 585
R1205 B.n214 B.n213 585
R1206 B.n215 B.n214 585
R1207 B.n608 B.n607 585
R1208 B.n607 B.n606 585
R1209 B.n609 B.n212 585
R1210 B.n212 B.n211 585
R1211 B.n611 B.n610 585
R1212 B.n612 B.n611 585
R1213 B.n206 B.n205 585
R1214 B.n207 B.n206 585
R1215 B.n620 B.n619 585
R1216 B.n619 B.n618 585
R1217 B.n621 B.n204 585
R1218 B.n204 B.n202 585
R1219 B.n623 B.n622 585
R1220 B.n624 B.n623 585
R1221 B.n198 B.n197 585
R1222 B.n203 B.n198 585
R1223 B.n632 B.n631 585
R1224 B.n631 B.n630 585
R1225 B.n633 B.n196 585
R1226 B.n196 B.n195 585
R1227 B.n635 B.n634 585
R1228 B.n636 B.n635 585
R1229 B.n190 B.n189 585
R1230 B.n191 B.n190 585
R1231 B.n644 B.n643 585
R1232 B.n643 B.n642 585
R1233 B.n645 B.n188 585
R1234 B.n188 B.n187 585
R1235 B.n647 B.n646 585
R1236 B.n648 B.n647 585
R1237 B.n182 B.n181 585
R1238 B.n183 B.n182 585
R1239 B.n656 B.n655 585
R1240 B.n655 B.n654 585
R1241 B.n657 B.n180 585
R1242 B.n180 B.n179 585
R1243 B.n659 B.n658 585
R1244 B.n660 B.n659 585
R1245 B.n174 B.n173 585
R1246 B.n175 B.n174 585
R1247 B.n668 B.n667 585
R1248 B.n667 B.n666 585
R1249 B.n669 B.n172 585
R1250 B.n172 B.n171 585
R1251 B.n671 B.n670 585
R1252 B.n672 B.n671 585
R1253 B.n166 B.n165 585
R1254 B.n167 B.n166 585
R1255 B.n681 B.n680 585
R1256 B.n680 B.n679 585
R1257 B.n682 B.n164 585
R1258 B.n164 B.n163 585
R1259 B.n684 B.n683 585
R1260 B.n685 B.n684 585
R1261 B.n3 B.n0 585
R1262 B.n4 B.n3 585
R1263 B.n1066 B.n1 585
R1264 B.n1067 B.n1066 585
R1265 B.n1065 B.n1064 585
R1266 B.n1065 B.n8 585
R1267 B.n1063 B.n9 585
R1268 B.n12 B.n9 585
R1269 B.n1062 B.n1061 585
R1270 B.n1061 B.n1060 585
R1271 B.n11 B.n10 585
R1272 B.n1059 B.n11 585
R1273 B.n1057 B.n1056 585
R1274 B.n1058 B.n1057 585
R1275 B.n1055 B.n17 585
R1276 B.n17 B.n16 585
R1277 B.n1054 B.n1053 585
R1278 B.n1053 B.n1052 585
R1279 B.n19 B.n18 585
R1280 B.n1051 B.n19 585
R1281 B.n1049 B.n1048 585
R1282 B.n1050 B.n1049 585
R1283 B.n1047 B.n24 585
R1284 B.n24 B.n23 585
R1285 B.n1046 B.n1045 585
R1286 B.n1045 B.n1044 585
R1287 B.n26 B.n25 585
R1288 B.n1043 B.n26 585
R1289 B.n1041 B.n1040 585
R1290 B.n1042 B.n1041 585
R1291 B.n1039 B.n31 585
R1292 B.n31 B.n30 585
R1293 B.n1038 B.n1037 585
R1294 B.n1037 B.n1036 585
R1295 B.n33 B.n32 585
R1296 B.n1035 B.n33 585
R1297 B.n1033 B.n1032 585
R1298 B.n1034 B.n1033 585
R1299 B.n1031 B.n38 585
R1300 B.n38 B.n37 585
R1301 B.n1030 B.n1029 585
R1302 B.n1029 B.n1028 585
R1303 B.n40 B.n39 585
R1304 B.n1027 B.n40 585
R1305 B.n1025 B.n1024 585
R1306 B.n1026 B.n1025 585
R1307 B.n1023 B.n45 585
R1308 B.n45 B.n44 585
R1309 B.n1022 B.n1021 585
R1310 B.n1021 B.n1020 585
R1311 B.n47 B.n46 585
R1312 B.n1019 B.n47 585
R1313 B.n1017 B.n1016 585
R1314 B.n1018 B.n1017 585
R1315 B.n1015 B.n52 585
R1316 B.n52 B.n51 585
R1317 B.n1014 B.n1013 585
R1318 B.n1013 B.n1012 585
R1319 B.n54 B.n53 585
R1320 B.n1011 B.n54 585
R1321 B.n1009 B.n1008 585
R1322 B.n1010 B.n1009 585
R1323 B.n1007 B.n59 585
R1324 B.n59 B.n58 585
R1325 B.n1006 B.n1005 585
R1326 B.n1005 B.n1004 585
R1327 B.n61 B.n60 585
R1328 B.n1003 B.n61 585
R1329 B.n1001 B.n1000 585
R1330 B.n1002 B.n1001 585
R1331 B.n999 B.n66 585
R1332 B.n66 B.n65 585
R1333 B.n998 B.n997 585
R1334 B.n997 B.n996 585
R1335 B.n68 B.n67 585
R1336 B.n995 B.n68 585
R1337 B.n993 B.n992 585
R1338 B.n994 B.n993 585
R1339 B.n991 B.n73 585
R1340 B.n73 B.n72 585
R1341 B.n990 B.n989 585
R1342 B.n989 B.n988 585
R1343 B.n75 B.n74 585
R1344 B.n987 B.n75 585
R1345 B.n985 B.n984 585
R1346 B.n986 B.n985 585
R1347 B.n983 B.n80 585
R1348 B.n80 B.n79 585
R1349 B.n982 B.n981 585
R1350 B.n981 B.n980 585
R1351 B.n82 B.n81 585
R1352 B.n979 B.n82 585
R1353 B.n977 B.n976 585
R1354 B.n978 B.n977 585
R1355 B.n975 B.n87 585
R1356 B.n87 B.n86 585
R1357 B.n974 B.n973 585
R1358 B.n973 B.n972 585
R1359 B.n89 B.n88 585
R1360 B.n971 B.n89 585
R1361 B.n969 B.n968 585
R1362 B.n970 B.n969 585
R1363 B.n967 B.n94 585
R1364 B.n94 B.n93 585
R1365 B.n966 B.n965 585
R1366 B.n965 B.n964 585
R1367 B.n96 B.n95 585
R1368 B.n963 B.n96 585
R1369 B.n961 B.n960 585
R1370 B.n962 B.n961 585
R1371 B.n959 B.n101 585
R1372 B.n101 B.n100 585
R1373 B.n958 B.n957 585
R1374 B.n957 B.n956 585
R1375 B.n103 B.n102 585
R1376 B.n955 B.n103 585
R1377 B.n953 B.n952 585
R1378 B.n954 B.n953 585
R1379 B.n1070 B.n1069 585
R1380 B.n1068 B.n2 585
R1381 B.n953 B.n108 521.33
R1382 B.n765 B.n106 521.33
R1383 B.n517 B.n274 521.33
R1384 B.n515 B.n276 521.33
R1385 B.n129 B.t12 368.892
R1386 B.n137 B.t18 368.892
R1387 B.n306 B.t9 368.892
R1388 B.n299 B.t16 368.892
R1389 B.n138 B.t19 285.5
R1390 B.n307 B.t8 285.5
R1391 B.n130 B.t13 285.5
R1392 B.n300 B.t15 285.5
R1393 B.n129 B.t10 283.409
R1394 B.n137 B.t17 283.409
R1395 B.n306 B.t6 283.409
R1396 B.n299 B.t14 283.409
R1397 B.n764 B.n107 256.663
R1398 B.n770 B.n107 256.663
R1399 B.n772 B.n107 256.663
R1400 B.n778 B.n107 256.663
R1401 B.n780 B.n107 256.663
R1402 B.n786 B.n107 256.663
R1403 B.n788 B.n107 256.663
R1404 B.n794 B.n107 256.663
R1405 B.n796 B.n107 256.663
R1406 B.n802 B.n107 256.663
R1407 B.n804 B.n107 256.663
R1408 B.n810 B.n107 256.663
R1409 B.n812 B.n107 256.663
R1410 B.n818 B.n107 256.663
R1411 B.n820 B.n107 256.663
R1412 B.n826 B.n107 256.663
R1413 B.n828 B.n107 256.663
R1414 B.n834 B.n107 256.663
R1415 B.n836 B.n107 256.663
R1416 B.n842 B.n107 256.663
R1417 B.n140 B.n107 256.663
R1418 B.n848 B.n107 256.663
R1419 B.n854 B.n107 256.663
R1420 B.n856 B.n107 256.663
R1421 B.n862 B.n107 256.663
R1422 B.n132 B.n107 256.663
R1423 B.n868 B.n107 256.663
R1424 B.n874 B.n107 256.663
R1425 B.n876 B.n107 256.663
R1426 B.n882 B.n107 256.663
R1427 B.n884 B.n107 256.663
R1428 B.n890 B.n107 256.663
R1429 B.n892 B.n107 256.663
R1430 B.n898 B.n107 256.663
R1431 B.n900 B.n107 256.663
R1432 B.n906 B.n107 256.663
R1433 B.n908 B.n107 256.663
R1434 B.n914 B.n107 256.663
R1435 B.n916 B.n107 256.663
R1436 B.n922 B.n107 256.663
R1437 B.n924 B.n107 256.663
R1438 B.n930 B.n107 256.663
R1439 B.n932 B.n107 256.663
R1440 B.n938 B.n107 256.663
R1441 B.n940 B.n107 256.663
R1442 B.n946 B.n107 256.663
R1443 B.n948 B.n107 256.663
R1444 B.n510 B.n275 256.663
R1445 B.n278 B.n275 256.663
R1446 B.n503 B.n275 256.663
R1447 B.n497 B.n275 256.663
R1448 B.n495 B.n275 256.663
R1449 B.n489 B.n275 256.663
R1450 B.n487 B.n275 256.663
R1451 B.n481 B.n275 256.663
R1452 B.n479 B.n275 256.663
R1453 B.n473 B.n275 256.663
R1454 B.n471 B.n275 256.663
R1455 B.n465 B.n275 256.663
R1456 B.n463 B.n275 256.663
R1457 B.n457 B.n275 256.663
R1458 B.n455 B.n275 256.663
R1459 B.n449 B.n275 256.663
R1460 B.n447 B.n275 256.663
R1461 B.n441 B.n275 256.663
R1462 B.n439 B.n275 256.663
R1463 B.n433 B.n275 256.663
R1464 B.n431 B.n275 256.663
R1465 B.n425 B.n275 256.663
R1466 B.n423 B.n275 256.663
R1467 B.n417 B.n275 256.663
R1468 B.n415 B.n275 256.663
R1469 B.n408 B.n275 256.663
R1470 B.n406 B.n275 256.663
R1471 B.n400 B.n275 256.663
R1472 B.n398 B.n275 256.663
R1473 B.n392 B.n275 256.663
R1474 B.n390 B.n275 256.663
R1475 B.n384 B.n275 256.663
R1476 B.n382 B.n275 256.663
R1477 B.n376 B.n275 256.663
R1478 B.n374 B.n275 256.663
R1479 B.n368 B.n275 256.663
R1480 B.n366 B.n275 256.663
R1481 B.n360 B.n275 256.663
R1482 B.n358 B.n275 256.663
R1483 B.n352 B.n275 256.663
R1484 B.n350 B.n275 256.663
R1485 B.n344 B.n275 256.663
R1486 B.n342 B.n275 256.663
R1487 B.n336 B.n275 256.663
R1488 B.n334 B.n275 256.663
R1489 B.n328 B.n275 256.663
R1490 B.n1072 B.n1071 256.663
R1491 B.n949 B.n947 163.367
R1492 B.n945 B.n110 163.367
R1493 B.n941 B.n939 163.367
R1494 B.n937 B.n112 163.367
R1495 B.n933 B.n931 163.367
R1496 B.n929 B.n114 163.367
R1497 B.n925 B.n923 163.367
R1498 B.n921 B.n116 163.367
R1499 B.n917 B.n915 163.367
R1500 B.n913 B.n118 163.367
R1501 B.n909 B.n907 163.367
R1502 B.n905 B.n120 163.367
R1503 B.n901 B.n899 163.367
R1504 B.n897 B.n122 163.367
R1505 B.n893 B.n891 163.367
R1506 B.n889 B.n124 163.367
R1507 B.n885 B.n883 163.367
R1508 B.n881 B.n126 163.367
R1509 B.n877 B.n875 163.367
R1510 B.n873 B.n128 163.367
R1511 B.n869 B.n867 163.367
R1512 B.n864 B.n863 163.367
R1513 B.n861 B.n134 163.367
R1514 B.n857 B.n855 163.367
R1515 B.n853 B.n136 163.367
R1516 B.n849 B.n847 163.367
R1517 B.n844 B.n843 163.367
R1518 B.n841 B.n142 163.367
R1519 B.n837 B.n835 163.367
R1520 B.n833 B.n144 163.367
R1521 B.n829 B.n827 163.367
R1522 B.n825 B.n146 163.367
R1523 B.n821 B.n819 163.367
R1524 B.n817 B.n148 163.367
R1525 B.n813 B.n811 163.367
R1526 B.n809 B.n150 163.367
R1527 B.n805 B.n803 163.367
R1528 B.n801 B.n152 163.367
R1529 B.n797 B.n795 163.367
R1530 B.n793 B.n154 163.367
R1531 B.n789 B.n787 163.367
R1532 B.n785 B.n156 163.367
R1533 B.n781 B.n779 163.367
R1534 B.n777 B.n158 163.367
R1535 B.n773 B.n771 163.367
R1536 B.n769 B.n160 163.367
R1537 B.n517 B.n272 163.367
R1538 B.n521 B.n272 163.367
R1539 B.n521 B.n266 163.367
R1540 B.n529 B.n266 163.367
R1541 B.n529 B.n264 163.367
R1542 B.n533 B.n264 163.367
R1543 B.n533 B.n257 163.367
R1544 B.n541 B.n257 163.367
R1545 B.n541 B.n255 163.367
R1546 B.n545 B.n255 163.367
R1547 B.n545 B.n250 163.367
R1548 B.n553 B.n250 163.367
R1549 B.n553 B.n248 163.367
R1550 B.n557 B.n248 163.367
R1551 B.n557 B.n242 163.367
R1552 B.n565 B.n242 163.367
R1553 B.n565 B.n240 163.367
R1554 B.n569 B.n240 163.367
R1555 B.n569 B.n234 163.367
R1556 B.n577 B.n234 163.367
R1557 B.n577 B.n232 163.367
R1558 B.n581 B.n232 163.367
R1559 B.n581 B.n225 163.367
R1560 B.n589 B.n225 163.367
R1561 B.n589 B.n223 163.367
R1562 B.n593 B.n223 163.367
R1563 B.n593 B.n218 163.367
R1564 B.n601 B.n218 163.367
R1565 B.n601 B.n216 163.367
R1566 B.n605 B.n216 163.367
R1567 B.n605 B.n210 163.367
R1568 B.n613 B.n210 163.367
R1569 B.n613 B.n208 163.367
R1570 B.n617 B.n208 163.367
R1571 B.n617 B.n201 163.367
R1572 B.n625 B.n201 163.367
R1573 B.n625 B.n199 163.367
R1574 B.n629 B.n199 163.367
R1575 B.n629 B.n194 163.367
R1576 B.n637 B.n194 163.367
R1577 B.n637 B.n192 163.367
R1578 B.n641 B.n192 163.367
R1579 B.n641 B.n186 163.367
R1580 B.n649 B.n186 163.367
R1581 B.n649 B.n184 163.367
R1582 B.n653 B.n184 163.367
R1583 B.n653 B.n178 163.367
R1584 B.n661 B.n178 163.367
R1585 B.n661 B.n176 163.367
R1586 B.n665 B.n176 163.367
R1587 B.n665 B.n170 163.367
R1588 B.n673 B.n170 163.367
R1589 B.n673 B.n168 163.367
R1590 B.n678 B.n168 163.367
R1591 B.n678 B.n162 163.367
R1592 B.n686 B.n162 163.367
R1593 B.n687 B.n686 163.367
R1594 B.n687 B.n5 163.367
R1595 B.n6 B.n5 163.367
R1596 B.n7 B.n6 163.367
R1597 B.n693 B.n7 163.367
R1598 B.n694 B.n693 163.367
R1599 B.n694 B.n13 163.367
R1600 B.n14 B.n13 163.367
R1601 B.n15 B.n14 163.367
R1602 B.n699 B.n15 163.367
R1603 B.n699 B.n20 163.367
R1604 B.n21 B.n20 163.367
R1605 B.n22 B.n21 163.367
R1606 B.n704 B.n22 163.367
R1607 B.n704 B.n27 163.367
R1608 B.n28 B.n27 163.367
R1609 B.n29 B.n28 163.367
R1610 B.n709 B.n29 163.367
R1611 B.n709 B.n34 163.367
R1612 B.n35 B.n34 163.367
R1613 B.n36 B.n35 163.367
R1614 B.n714 B.n36 163.367
R1615 B.n714 B.n41 163.367
R1616 B.n42 B.n41 163.367
R1617 B.n43 B.n42 163.367
R1618 B.n719 B.n43 163.367
R1619 B.n719 B.n48 163.367
R1620 B.n49 B.n48 163.367
R1621 B.n50 B.n49 163.367
R1622 B.n724 B.n50 163.367
R1623 B.n724 B.n55 163.367
R1624 B.n56 B.n55 163.367
R1625 B.n57 B.n56 163.367
R1626 B.n729 B.n57 163.367
R1627 B.n729 B.n62 163.367
R1628 B.n63 B.n62 163.367
R1629 B.n64 B.n63 163.367
R1630 B.n734 B.n64 163.367
R1631 B.n734 B.n69 163.367
R1632 B.n70 B.n69 163.367
R1633 B.n71 B.n70 163.367
R1634 B.n739 B.n71 163.367
R1635 B.n739 B.n76 163.367
R1636 B.n77 B.n76 163.367
R1637 B.n78 B.n77 163.367
R1638 B.n744 B.n78 163.367
R1639 B.n744 B.n83 163.367
R1640 B.n84 B.n83 163.367
R1641 B.n85 B.n84 163.367
R1642 B.n749 B.n85 163.367
R1643 B.n749 B.n90 163.367
R1644 B.n91 B.n90 163.367
R1645 B.n92 B.n91 163.367
R1646 B.n754 B.n92 163.367
R1647 B.n754 B.n97 163.367
R1648 B.n98 B.n97 163.367
R1649 B.n99 B.n98 163.367
R1650 B.n759 B.n99 163.367
R1651 B.n759 B.n104 163.367
R1652 B.n105 B.n104 163.367
R1653 B.n106 B.n105 163.367
R1654 B.n511 B.n509 163.367
R1655 B.n509 B.n508 163.367
R1656 B.n505 B.n504 163.367
R1657 B.n502 B.n280 163.367
R1658 B.n498 B.n496 163.367
R1659 B.n494 B.n282 163.367
R1660 B.n490 B.n488 163.367
R1661 B.n486 B.n284 163.367
R1662 B.n482 B.n480 163.367
R1663 B.n478 B.n286 163.367
R1664 B.n474 B.n472 163.367
R1665 B.n470 B.n288 163.367
R1666 B.n466 B.n464 163.367
R1667 B.n462 B.n290 163.367
R1668 B.n458 B.n456 163.367
R1669 B.n454 B.n292 163.367
R1670 B.n450 B.n448 163.367
R1671 B.n446 B.n294 163.367
R1672 B.n442 B.n440 163.367
R1673 B.n438 B.n296 163.367
R1674 B.n434 B.n432 163.367
R1675 B.n430 B.n298 163.367
R1676 B.n426 B.n424 163.367
R1677 B.n422 B.n303 163.367
R1678 B.n418 B.n416 163.367
R1679 B.n414 B.n305 163.367
R1680 B.n409 B.n407 163.367
R1681 B.n405 B.n309 163.367
R1682 B.n401 B.n399 163.367
R1683 B.n397 B.n311 163.367
R1684 B.n393 B.n391 163.367
R1685 B.n389 B.n313 163.367
R1686 B.n385 B.n383 163.367
R1687 B.n381 B.n315 163.367
R1688 B.n377 B.n375 163.367
R1689 B.n373 B.n317 163.367
R1690 B.n369 B.n367 163.367
R1691 B.n365 B.n319 163.367
R1692 B.n361 B.n359 163.367
R1693 B.n357 B.n321 163.367
R1694 B.n353 B.n351 163.367
R1695 B.n349 B.n323 163.367
R1696 B.n345 B.n343 163.367
R1697 B.n341 B.n325 163.367
R1698 B.n337 B.n335 163.367
R1699 B.n333 B.n327 163.367
R1700 B.n329 B.n274 163.367
R1701 B.n515 B.n270 163.367
R1702 B.n523 B.n270 163.367
R1703 B.n523 B.n268 163.367
R1704 B.n527 B.n268 163.367
R1705 B.n527 B.n262 163.367
R1706 B.n535 B.n262 163.367
R1707 B.n535 B.n260 163.367
R1708 B.n539 B.n260 163.367
R1709 B.n539 B.n254 163.367
R1710 B.n547 B.n254 163.367
R1711 B.n547 B.n252 163.367
R1712 B.n551 B.n252 163.367
R1713 B.n551 B.n246 163.367
R1714 B.n559 B.n246 163.367
R1715 B.n559 B.n244 163.367
R1716 B.n563 B.n244 163.367
R1717 B.n563 B.n238 163.367
R1718 B.n571 B.n238 163.367
R1719 B.n571 B.n236 163.367
R1720 B.n575 B.n236 163.367
R1721 B.n575 B.n230 163.367
R1722 B.n583 B.n230 163.367
R1723 B.n583 B.n228 163.367
R1724 B.n587 B.n228 163.367
R1725 B.n587 B.n222 163.367
R1726 B.n595 B.n222 163.367
R1727 B.n595 B.n220 163.367
R1728 B.n599 B.n220 163.367
R1729 B.n599 B.n214 163.367
R1730 B.n607 B.n214 163.367
R1731 B.n607 B.n212 163.367
R1732 B.n611 B.n212 163.367
R1733 B.n611 B.n206 163.367
R1734 B.n619 B.n206 163.367
R1735 B.n619 B.n204 163.367
R1736 B.n623 B.n204 163.367
R1737 B.n623 B.n198 163.367
R1738 B.n631 B.n198 163.367
R1739 B.n631 B.n196 163.367
R1740 B.n635 B.n196 163.367
R1741 B.n635 B.n190 163.367
R1742 B.n643 B.n190 163.367
R1743 B.n643 B.n188 163.367
R1744 B.n647 B.n188 163.367
R1745 B.n647 B.n182 163.367
R1746 B.n655 B.n182 163.367
R1747 B.n655 B.n180 163.367
R1748 B.n659 B.n180 163.367
R1749 B.n659 B.n174 163.367
R1750 B.n667 B.n174 163.367
R1751 B.n667 B.n172 163.367
R1752 B.n671 B.n172 163.367
R1753 B.n671 B.n166 163.367
R1754 B.n680 B.n166 163.367
R1755 B.n680 B.n164 163.367
R1756 B.n684 B.n164 163.367
R1757 B.n684 B.n3 163.367
R1758 B.n1070 B.n3 163.367
R1759 B.n1066 B.n2 163.367
R1760 B.n1066 B.n1065 163.367
R1761 B.n1065 B.n9 163.367
R1762 B.n1061 B.n9 163.367
R1763 B.n1061 B.n11 163.367
R1764 B.n1057 B.n11 163.367
R1765 B.n1057 B.n17 163.367
R1766 B.n1053 B.n17 163.367
R1767 B.n1053 B.n19 163.367
R1768 B.n1049 B.n19 163.367
R1769 B.n1049 B.n24 163.367
R1770 B.n1045 B.n24 163.367
R1771 B.n1045 B.n26 163.367
R1772 B.n1041 B.n26 163.367
R1773 B.n1041 B.n31 163.367
R1774 B.n1037 B.n31 163.367
R1775 B.n1037 B.n33 163.367
R1776 B.n1033 B.n33 163.367
R1777 B.n1033 B.n38 163.367
R1778 B.n1029 B.n38 163.367
R1779 B.n1029 B.n40 163.367
R1780 B.n1025 B.n40 163.367
R1781 B.n1025 B.n45 163.367
R1782 B.n1021 B.n45 163.367
R1783 B.n1021 B.n47 163.367
R1784 B.n1017 B.n47 163.367
R1785 B.n1017 B.n52 163.367
R1786 B.n1013 B.n52 163.367
R1787 B.n1013 B.n54 163.367
R1788 B.n1009 B.n54 163.367
R1789 B.n1009 B.n59 163.367
R1790 B.n1005 B.n59 163.367
R1791 B.n1005 B.n61 163.367
R1792 B.n1001 B.n61 163.367
R1793 B.n1001 B.n66 163.367
R1794 B.n997 B.n66 163.367
R1795 B.n997 B.n68 163.367
R1796 B.n993 B.n68 163.367
R1797 B.n993 B.n73 163.367
R1798 B.n989 B.n73 163.367
R1799 B.n989 B.n75 163.367
R1800 B.n985 B.n75 163.367
R1801 B.n985 B.n80 163.367
R1802 B.n981 B.n80 163.367
R1803 B.n981 B.n82 163.367
R1804 B.n977 B.n82 163.367
R1805 B.n977 B.n87 163.367
R1806 B.n973 B.n87 163.367
R1807 B.n973 B.n89 163.367
R1808 B.n969 B.n89 163.367
R1809 B.n969 B.n94 163.367
R1810 B.n965 B.n94 163.367
R1811 B.n965 B.n96 163.367
R1812 B.n961 B.n96 163.367
R1813 B.n961 B.n101 163.367
R1814 B.n957 B.n101 163.367
R1815 B.n957 B.n103 163.367
R1816 B.n953 B.n103 163.367
R1817 B.n516 B.n275 86.3368
R1818 B.n954 B.n107 86.3368
R1819 B.n130 B.n129 83.3944
R1820 B.n138 B.n137 83.3944
R1821 B.n307 B.n306 83.3944
R1822 B.n300 B.n299 83.3944
R1823 B.n948 B.n108 71.676
R1824 B.n947 B.n946 71.676
R1825 B.n940 B.n110 71.676
R1826 B.n939 B.n938 71.676
R1827 B.n932 B.n112 71.676
R1828 B.n931 B.n930 71.676
R1829 B.n924 B.n114 71.676
R1830 B.n923 B.n922 71.676
R1831 B.n916 B.n116 71.676
R1832 B.n915 B.n914 71.676
R1833 B.n908 B.n118 71.676
R1834 B.n907 B.n906 71.676
R1835 B.n900 B.n120 71.676
R1836 B.n899 B.n898 71.676
R1837 B.n892 B.n122 71.676
R1838 B.n891 B.n890 71.676
R1839 B.n884 B.n124 71.676
R1840 B.n883 B.n882 71.676
R1841 B.n876 B.n126 71.676
R1842 B.n875 B.n874 71.676
R1843 B.n868 B.n128 71.676
R1844 B.n867 B.n132 71.676
R1845 B.n863 B.n862 71.676
R1846 B.n856 B.n134 71.676
R1847 B.n855 B.n854 71.676
R1848 B.n848 B.n136 71.676
R1849 B.n847 B.n140 71.676
R1850 B.n843 B.n842 71.676
R1851 B.n836 B.n142 71.676
R1852 B.n835 B.n834 71.676
R1853 B.n828 B.n144 71.676
R1854 B.n827 B.n826 71.676
R1855 B.n820 B.n146 71.676
R1856 B.n819 B.n818 71.676
R1857 B.n812 B.n148 71.676
R1858 B.n811 B.n810 71.676
R1859 B.n804 B.n150 71.676
R1860 B.n803 B.n802 71.676
R1861 B.n796 B.n152 71.676
R1862 B.n795 B.n794 71.676
R1863 B.n788 B.n154 71.676
R1864 B.n787 B.n786 71.676
R1865 B.n780 B.n156 71.676
R1866 B.n779 B.n778 71.676
R1867 B.n772 B.n158 71.676
R1868 B.n771 B.n770 71.676
R1869 B.n764 B.n160 71.676
R1870 B.n765 B.n764 71.676
R1871 B.n770 B.n769 71.676
R1872 B.n773 B.n772 71.676
R1873 B.n778 B.n777 71.676
R1874 B.n781 B.n780 71.676
R1875 B.n786 B.n785 71.676
R1876 B.n789 B.n788 71.676
R1877 B.n794 B.n793 71.676
R1878 B.n797 B.n796 71.676
R1879 B.n802 B.n801 71.676
R1880 B.n805 B.n804 71.676
R1881 B.n810 B.n809 71.676
R1882 B.n813 B.n812 71.676
R1883 B.n818 B.n817 71.676
R1884 B.n821 B.n820 71.676
R1885 B.n826 B.n825 71.676
R1886 B.n829 B.n828 71.676
R1887 B.n834 B.n833 71.676
R1888 B.n837 B.n836 71.676
R1889 B.n842 B.n841 71.676
R1890 B.n844 B.n140 71.676
R1891 B.n849 B.n848 71.676
R1892 B.n854 B.n853 71.676
R1893 B.n857 B.n856 71.676
R1894 B.n862 B.n861 71.676
R1895 B.n864 B.n132 71.676
R1896 B.n869 B.n868 71.676
R1897 B.n874 B.n873 71.676
R1898 B.n877 B.n876 71.676
R1899 B.n882 B.n881 71.676
R1900 B.n885 B.n884 71.676
R1901 B.n890 B.n889 71.676
R1902 B.n893 B.n892 71.676
R1903 B.n898 B.n897 71.676
R1904 B.n901 B.n900 71.676
R1905 B.n906 B.n905 71.676
R1906 B.n909 B.n908 71.676
R1907 B.n914 B.n913 71.676
R1908 B.n917 B.n916 71.676
R1909 B.n922 B.n921 71.676
R1910 B.n925 B.n924 71.676
R1911 B.n930 B.n929 71.676
R1912 B.n933 B.n932 71.676
R1913 B.n938 B.n937 71.676
R1914 B.n941 B.n940 71.676
R1915 B.n946 B.n945 71.676
R1916 B.n949 B.n948 71.676
R1917 B.n510 B.n276 71.676
R1918 B.n508 B.n278 71.676
R1919 B.n504 B.n503 71.676
R1920 B.n497 B.n280 71.676
R1921 B.n496 B.n495 71.676
R1922 B.n489 B.n282 71.676
R1923 B.n488 B.n487 71.676
R1924 B.n481 B.n284 71.676
R1925 B.n480 B.n479 71.676
R1926 B.n473 B.n286 71.676
R1927 B.n472 B.n471 71.676
R1928 B.n465 B.n288 71.676
R1929 B.n464 B.n463 71.676
R1930 B.n457 B.n290 71.676
R1931 B.n456 B.n455 71.676
R1932 B.n449 B.n292 71.676
R1933 B.n448 B.n447 71.676
R1934 B.n441 B.n294 71.676
R1935 B.n440 B.n439 71.676
R1936 B.n433 B.n296 71.676
R1937 B.n432 B.n431 71.676
R1938 B.n425 B.n298 71.676
R1939 B.n424 B.n423 71.676
R1940 B.n417 B.n303 71.676
R1941 B.n416 B.n415 71.676
R1942 B.n408 B.n305 71.676
R1943 B.n407 B.n406 71.676
R1944 B.n400 B.n309 71.676
R1945 B.n399 B.n398 71.676
R1946 B.n392 B.n311 71.676
R1947 B.n391 B.n390 71.676
R1948 B.n384 B.n313 71.676
R1949 B.n383 B.n382 71.676
R1950 B.n376 B.n315 71.676
R1951 B.n375 B.n374 71.676
R1952 B.n368 B.n317 71.676
R1953 B.n367 B.n366 71.676
R1954 B.n360 B.n319 71.676
R1955 B.n359 B.n358 71.676
R1956 B.n352 B.n321 71.676
R1957 B.n351 B.n350 71.676
R1958 B.n344 B.n323 71.676
R1959 B.n343 B.n342 71.676
R1960 B.n336 B.n325 71.676
R1961 B.n335 B.n334 71.676
R1962 B.n328 B.n327 71.676
R1963 B.n511 B.n510 71.676
R1964 B.n505 B.n278 71.676
R1965 B.n503 B.n502 71.676
R1966 B.n498 B.n497 71.676
R1967 B.n495 B.n494 71.676
R1968 B.n490 B.n489 71.676
R1969 B.n487 B.n486 71.676
R1970 B.n482 B.n481 71.676
R1971 B.n479 B.n478 71.676
R1972 B.n474 B.n473 71.676
R1973 B.n471 B.n470 71.676
R1974 B.n466 B.n465 71.676
R1975 B.n463 B.n462 71.676
R1976 B.n458 B.n457 71.676
R1977 B.n455 B.n454 71.676
R1978 B.n450 B.n449 71.676
R1979 B.n447 B.n446 71.676
R1980 B.n442 B.n441 71.676
R1981 B.n439 B.n438 71.676
R1982 B.n434 B.n433 71.676
R1983 B.n431 B.n430 71.676
R1984 B.n426 B.n425 71.676
R1985 B.n423 B.n422 71.676
R1986 B.n418 B.n417 71.676
R1987 B.n415 B.n414 71.676
R1988 B.n409 B.n408 71.676
R1989 B.n406 B.n405 71.676
R1990 B.n401 B.n400 71.676
R1991 B.n398 B.n397 71.676
R1992 B.n393 B.n392 71.676
R1993 B.n390 B.n389 71.676
R1994 B.n385 B.n384 71.676
R1995 B.n382 B.n381 71.676
R1996 B.n377 B.n376 71.676
R1997 B.n374 B.n373 71.676
R1998 B.n369 B.n368 71.676
R1999 B.n366 B.n365 71.676
R2000 B.n361 B.n360 71.676
R2001 B.n358 B.n357 71.676
R2002 B.n353 B.n352 71.676
R2003 B.n350 B.n349 71.676
R2004 B.n345 B.n344 71.676
R2005 B.n342 B.n341 71.676
R2006 B.n337 B.n336 71.676
R2007 B.n334 B.n333 71.676
R2008 B.n329 B.n328 71.676
R2009 B.n1071 B.n1070 71.676
R2010 B.n1071 B.n2 71.676
R2011 B.n131 B.n130 59.5399
R2012 B.n139 B.n138 59.5399
R2013 B.n411 B.n307 59.5399
R2014 B.n301 B.n300 59.5399
R2015 B.n516 B.n271 42.8536
R2016 B.n522 B.n271 42.8536
R2017 B.n522 B.n267 42.8536
R2018 B.n528 B.n267 42.8536
R2019 B.n528 B.n263 42.8536
R2020 B.n534 B.n263 42.8536
R2021 B.n534 B.n258 42.8536
R2022 B.n540 B.n258 42.8536
R2023 B.n540 B.n259 42.8536
R2024 B.n546 B.n251 42.8536
R2025 B.n552 B.n251 42.8536
R2026 B.n552 B.n247 42.8536
R2027 B.n558 B.n247 42.8536
R2028 B.n558 B.n243 42.8536
R2029 B.n564 B.n243 42.8536
R2030 B.n564 B.n239 42.8536
R2031 B.n570 B.n239 42.8536
R2032 B.n570 B.n235 42.8536
R2033 B.n576 B.n235 42.8536
R2034 B.n576 B.n231 42.8536
R2035 B.n582 B.n231 42.8536
R2036 B.n582 B.n226 42.8536
R2037 B.n588 B.n226 42.8536
R2038 B.n588 B.n227 42.8536
R2039 B.n594 B.n219 42.8536
R2040 B.n600 B.n219 42.8536
R2041 B.n600 B.n215 42.8536
R2042 B.n606 B.n215 42.8536
R2043 B.n606 B.n211 42.8536
R2044 B.n612 B.n211 42.8536
R2045 B.n612 B.n207 42.8536
R2046 B.n618 B.n207 42.8536
R2047 B.n618 B.n202 42.8536
R2048 B.n624 B.n202 42.8536
R2049 B.n624 B.n203 42.8536
R2050 B.n630 B.n195 42.8536
R2051 B.n636 B.n195 42.8536
R2052 B.n636 B.n191 42.8536
R2053 B.n642 B.n191 42.8536
R2054 B.n642 B.n187 42.8536
R2055 B.n648 B.n187 42.8536
R2056 B.n648 B.n183 42.8536
R2057 B.n654 B.n183 42.8536
R2058 B.n654 B.n179 42.8536
R2059 B.n660 B.n179 42.8536
R2060 B.n660 B.n175 42.8536
R2061 B.n666 B.n175 42.8536
R2062 B.n672 B.n171 42.8536
R2063 B.n672 B.n167 42.8536
R2064 B.n679 B.n167 42.8536
R2065 B.n679 B.n163 42.8536
R2066 B.n685 B.n163 42.8536
R2067 B.n685 B.n4 42.8536
R2068 B.n1069 B.n4 42.8536
R2069 B.n1069 B.n1068 42.8536
R2070 B.n1068 B.n1067 42.8536
R2071 B.n1067 B.n8 42.8536
R2072 B.n12 B.n8 42.8536
R2073 B.n1060 B.n12 42.8536
R2074 B.n1060 B.n1059 42.8536
R2075 B.n1059 B.n1058 42.8536
R2076 B.n1058 B.n16 42.8536
R2077 B.n1052 B.n1051 42.8536
R2078 B.n1051 B.n1050 42.8536
R2079 B.n1050 B.n23 42.8536
R2080 B.n1044 B.n23 42.8536
R2081 B.n1044 B.n1043 42.8536
R2082 B.n1043 B.n1042 42.8536
R2083 B.n1042 B.n30 42.8536
R2084 B.n1036 B.n30 42.8536
R2085 B.n1036 B.n1035 42.8536
R2086 B.n1035 B.n1034 42.8536
R2087 B.n1034 B.n37 42.8536
R2088 B.n1028 B.n37 42.8536
R2089 B.n1027 B.n1026 42.8536
R2090 B.n1026 B.n44 42.8536
R2091 B.n1020 B.n44 42.8536
R2092 B.n1020 B.n1019 42.8536
R2093 B.n1019 B.n1018 42.8536
R2094 B.n1018 B.n51 42.8536
R2095 B.n1012 B.n51 42.8536
R2096 B.n1012 B.n1011 42.8536
R2097 B.n1011 B.n1010 42.8536
R2098 B.n1010 B.n58 42.8536
R2099 B.n1004 B.n58 42.8536
R2100 B.n1003 B.n1002 42.8536
R2101 B.n1002 B.n65 42.8536
R2102 B.n996 B.n65 42.8536
R2103 B.n996 B.n995 42.8536
R2104 B.n995 B.n994 42.8536
R2105 B.n994 B.n72 42.8536
R2106 B.n988 B.n72 42.8536
R2107 B.n988 B.n987 42.8536
R2108 B.n987 B.n986 42.8536
R2109 B.n986 B.n79 42.8536
R2110 B.n980 B.n79 42.8536
R2111 B.n980 B.n979 42.8536
R2112 B.n979 B.n978 42.8536
R2113 B.n978 B.n86 42.8536
R2114 B.n972 B.n86 42.8536
R2115 B.n971 B.n970 42.8536
R2116 B.n970 B.n93 42.8536
R2117 B.n964 B.n93 42.8536
R2118 B.n964 B.n963 42.8536
R2119 B.n963 B.n962 42.8536
R2120 B.n962 B.n100 42.8536
R2121 B.n956 B.n100 42.8536
R2122 B.n956 B.n955 42.8536
R2123 B.n955 B.n954 42.8536
R2124 B.n203 B.t3 39.7026
R2125 B.t4 B.n1027 39.7026
R2126 B.n514 B.n513 33.8737
R2127 B.n518 B.n273 33.8737
R2128 B.n766 B.n763 33.8737
R2129 B.n952 B.n951 33.8737
R2130 B.n594 B.t5 30.8799
R2131 B.n1004 B.t1 30.8799
R2132 B.n546 B.t7 24.578
R2133 B.n666 B.t0 24.578
R2134 B.n1052 B.t2 24.578
R2135 B.n972 B.t11 24.578
R2136 B.n259 B.t7 18.2761
R2137 B.t0 B.n171 18.2761
R2138 B.t2 B.n16 18.2761
R2139 B.t11 B.n971 18.2761
R2140 B B.n1072 18.0485
R2141 B.n227 B.t5 11.9741
R2142 B.t1 B.n1003 11.9741
R2143 B.n514 B.n269 10.6151
R2144 B.n524 B.n269 10.6151
R2145 B.n525 B.n524 10.6151
R2146 B.n526 B.n525 10.6151
R2147 B.n526 B.n261 10.6151
R2148 B.n536 B.n261 10.6151
R2149 B.n537 B.n536 10.6151
R2150 B.n538 B.n537 10.6151
R2151 B.n538 B.n253 10.6151
R2152 B.n548 B.n253 10.6151
R2153 B.n549 B.n548 10.6151
R2154 B.n550 B.n549 10.6151
R2155 B.n550 B.n245 10.6151
R2156 B.n560 B.n245 10.6151
R2157 B.n561 B.n560 10.6151
R2158 B.n562 B.n561 10.6151
R2159 B.n562 B.n237 10.6151
R2160 B.n572 B.n237 10.6151
R2161 B.n573 B.n572 10.6151
R2162 B.n574 B.n573 10.6151
R2163 B.n574 B.n229 10.6151
R2164 B.n584 B.n229 10.6151
R2165 B.n585 B.n584 10.6151
R2166 B.n586 B.n585 10.6151
R2167 B.n586 B.n221 10.6151
R2168 B.n596 B.n221 10.6151
R2169 B.n597 B.n596 10.6151
R2170 B.n598 B.n597 10.6151
R2171 B.n598 B.n213 10.6151
R2172 B.n608 B.n213 10.6151
R2173 B.n609 B.n608 10.6151
R2174 B.n610 B.n609 10.6151
R2175 B.n610 B.n205 10.6151
R2176 B.n620 B.n205 10.6151
R2177 B.n621 B.n620 10.6151
R2178 B.n622 B.n621 10.6151
R2179 B.n622 B.n197 10.6151
R2180 B.n632 B.n197 10.6151
R2181 B.n633 B.n632 10.6151
R2182 B.n634 B.n633 10.6151
R2183 B.n634 B.n189 10.6151
R2184 B.n644 B.n189 10.6151
R2185 B.n645 B.n644 10.6151
R2186 B.n646 B.n645 10.6151
R2187 B.n646 B.n181 10.6151
R2188 B.n656 B.n181 10.6151
R2189 B.n657 B.n656 10.6151
R2190 B.n658 B.n657 10.6151
R2191 B.n658 B.n173 10.6151
R2192 B.n668 B.n173 10.6151
R2193 B.n669 B.n668 10.6151
R2194 B.n670 B.n669 10.6151
R2195 B.n670 B.n165 10.6151
R2196 B.n681 B.n165 10.6151
R2197 B.n682 B.n681 10.6151
R2198 B.n683 B.n682 10.6151
R2199 B.n683 B.n0 10.6151
R2200 B.n513 B.n512 10.6151
R2201 B.n512 B.n277 10.6151
R2202 B.n507 B.n277 10.6151
R2203 B.n507 B.n506 10.6151
R2204 B.n506 B.n279 10.6151
R2205 B.n501 B.n279 10.6151
R2206 B.n501 B.n500 10.6151
R2207 B.n500 B.n499 10.6151
R2208 B.n499 B.n281 10.6151
R2209 B.n493 B.n281 10.6151
R2210 B.n493 B.n492 10.6151
R2211 B.n492 B.n491 10.6151
R2212 B.n491 B.n283 10.6151
R2213 B.n485 B.n283 10.6151
R2214 B.n485 B.n484 10.6151
R2215 B.n484 B.n483 10.6151
R2216 B.n483 B.n285 10.6151
R2217 B.n477 B.n285 10.6151
R2218 B.n477 B.n476 10.6151
R2219 B.n476 B.n475 10.6151
R2220 B.n475 B.n287 10.6151
R2221 B.n469 B.n287 10.6151
R2222 B.n469 B.n468 10.6151
R2223 B.n468 B.n467 10.6151
R2224 B.n467 B.n289 10.6151
R2225 B.n461 B.n289 10.6151
R2226 B.n461 B.n460 10.6151
R2227 B.n460 B.n459 10.6151
R2228 B.n459 B.n291 10.6151
R2229 B.n453 B.n291 10.6151
R2230 B.n453 B.n452 10.6151
R2231 B.n452 B.n451 10.6151
R2232 B.n451 B.n293 10.6151
R2233 B.n445 B.n293 10.6151
R2234 B.n445 B.n444 10.6151
R2235 B.n444 B.n443 10.6151
R2236 B.n443 B.n295 10.6151
R2237 B.n437 B.n295 10.6151
R2238 B.n437 B.n436 10.6151
R2239 B.n436 B.n435 10.6151
R2240 B.n435 B.n297 10.6151
R2241 B.n429 B.n428 10.6151
R2242 B.n428 B.n427 10.6151
R2243 B.n427 B.n302 10.6151
R2244 B.n421 B.n302 10.6151
R2245 B.n421 B.n420 10.6151
R2246 B.n420 B.n419 10.6151
R2247 B.n419 B.n304 10.6151
R2248 B.n413 B.n304 10.6151
R2249 B.n413 B.n412 10.6151
R2250 B.n410 B.n308 10.6151
R2251 B.n404 B.n308 10.6151
R2252 B.n404 B.n403 10.6151
R2253 B.n403 B.n402 10.6151
R2254 B.n402 B.n310 10.6151
R2255 B.n396 B.n310 10.6151
R2256 B.n396 B.n395 10.6151
R2257 B.n395 B.n394 10.6151
R2258 B.n394 B.n312 10.6151
R2259 B.n388 B.n312 10.6151
R2260 B.n388 B.n387 10.6151
R2261 B.n387 B.n386 10.6151
R2262 B.n386 B.n314 10.6151
R2263 B.n380 B.n314 10.6151
R2264 B.n380 B.n379 10.6151
R2265 B.n379 B.n378 10.6151
R2266 B.n378 B.n316 10.6151
R2267 B.n372 B.n316 10.6151
R2268 B.n372 B.n371 10.6151
R2269 B.n371 B.n370 10.6151
R2270 B.n370 B.n318 10.6151
R2271 B.n364 B.n318 10.6151
R2272 B.n364 B.n363 10.6151
R2273 B.n363 B.n362 10.6151
R2274 B.n362 B.n320 10.6151
R2275 B.n356 B.n320 10.6151
R2276 B.n356 B.n355 10.6151
R2277 B.n355 B.n354 10.6151
R2278 B.n354 B.n322 10.6151
R2279 B.n348 B.n322 10.6151
R2280 B.n348 B.n347 10.6151
R2281 B.n347 B.n346 10.6151
R2282 B.n346 B.n324 10.6151
R2283 B.n340 B.n324 10.6151
R2284 B.n340 B.n339 10.6151
R2285 B.n339 B.n338 10.6151
R2286 B.n338 B.n326 10.6151
R2287 B.n332 B.n326 10.6151
R2288 B.n332 B.n331 10.6151
R2289 B.n331 B.n330 10.6151
R2290 B.n330 B.n273 10.6151
R2291 B.n519 B.n518 10.6151
R2292 B.n520 B.n519 10.6151
R2293 B.n520 B.n265 10.6151
R2294 B.n530 B.n265 10.6151
R2295 B.n531 B.n530 10.6151
R2296 B.n532 B.n531 10.6151
R2297 B.n532 B.n256 10.6151
R2298 B.n542 B.n256 10.6151
R2299 B.n543 B.n542 10.6151
R2300 B.n544 B.n543 10.6151
R2301 B.n544 B.n249 10.6151
R2302 B.n554 B.n249 10.6151
R2303 B.n555 B.n554 10.6151
R2304 B.n556 B.n555 10.6151
R2305 B.n556 B.n241 10.6151
R2306 B.n566 B.n241 10.6151
R2307 B.n567 B.n566 10.6151
R2308 B.n568 B.n567 10.6151
R2309 B.n568 B.n233 10.6151
R2310 B.n578 B.n233 10.6151
R2311 B.n579 B.n578 10.6151
R2312 B.n580 B.n579 10.6151
R2313 B.n580 B.n224 10.6151
R2314 B.n590 B.n224 10.6151
R2315 B.n591 B.n590 10.6151
R2316 B.n592 B.n591 10.6151
R2317 B.n592 B.n217 10.6151
R2318 B.n602 B.n217 10.6151
R2319 B.n603 B.n602 10.6151
R2320 B.n604 B.n603 10.6151
R2321 B.n604 B.n209 10.6151
R2322 B.n614 B.n209 10.6151
R2323 B.n615 B.n614 10.6151
R2324 B.n616 B.n615 10.6151
R2325 B.n616 B.n200 10.6151
R2326 B.n626 B.n200 10.6151
R2327 B.n627 B.n626 10.6151
R2328 B.n628 B.n627 10.6151
R2329 B.n628 B.n193 10.6151
R2330 B.n638 B.n193 10.6151
R2331 B.n639 B.n638 10.6151
R2332 B.n640 B.n639 10.6151
R2333 B.n640 B.n185 10.6151
R2334 B.n650 B.n185 10.6151
R2335 B.n651 B.n650 10.6151
R2336 B.n652 B.n651 10.6151
R2337 B.n652 B.n177 10.6151
R2338 B.n662 B.n177 10.6151
R2339 B.n663 B.n662 10.6151
R2340 B.n664 B.n663 10.6151
R2341 B.n664 B.n169 10.6151
R2342 B.n674 B.n169 10.6151
R2343 B.n675 B.n674 10.6151
R2344 B.n677 B.n675 10.6151
R2345 B.n677 B.n676 10.6151
R2346 B.n676 B.n161 10.6151
R2347 B.n688 B.n161 10.6151
R2348 B.n689 B.n688 10.6151
R2349 B.n690 B.n689 10.6151
R2350 B.n691 B.n690 10.6151
R2351 B.n692 B.n691 10.6151
R2352 B.n695 B.n692 10.6151
R2353 B.n696 B.n695 10.6151
R2354 B.n697 B.n696 10.6151
R2355 B.n698 B.n697 10.6151
R2356 B.n700 B.n698 10.6151
R2357 B.n701 B.n700 10.6151
R2358 B.n702 B.n701 10.6151
R2359 B.n703 B.n702 10.6151
R2360 B.n705 B.n703 10.6151
R2361 B.n706 B.n705 10.6151
R2362 B.n707 B.n706 10.6151
R2363 B.n708 B.n707 10.6151
R2364 B.n710 B.n708 10.6151
R2365 B.n711 B.n710 10.6151
R2366 B.n712 B.n711 10.6151
R2367 B.n713 B.n712 10.6151
R2368 B.n715 B.n713 10.6151
R2369 B.n716 B.n715 10.6151
R2370 B.n717 B.n716 10.6151
R2371 B.n718 B.n717 10.6151
R2372 B.n720 B.n718 10.6151
R2373 B.n721 B.n720 10.6151
R2374 B.n722 B.n721 10.6151
R2375 B.n723 B.n722 10.6151
R2376 B.n725 B.n723 10.6151
R2377 B.n726 B.n725 10.6151
R2378 B.n727 B.n726 10.6151
R2379 B.n728 B.n727 10.6151
R2380 B.n730 B.n728 10.6151
R2381 B.n731 B.n730 10.6151
R2382 B.n732 B.n731 10.6151
R2383 B.n733 B.n732 10.6151
R2384 B.n735 B.n733 10.6151
R2385 B.n736 B.n735 10.6151
R2386 B.n737 B.n736 10.6151
R2387 B.n738 B.n737 10.6151
R2388 B.n740 B.n738 10.6151
R2389 B.n741 B.n740 10.6151
R2390 B.n742 B.n741 10.6151
R2391 B.n743 B.n742 10.6151
R2392 B.n745 B.n743 10.6151
R2393 B.n746 B.n745 10.6151
R2394 B.n747 B.n746 10.6151
R2395 B.n748 B.n747 10.6151
R2396 B.n750 B.n748 10.6151
R2397 B.n751 B.n750 10.6151
R2398 B.n752 B.n751 10.6151
R2399 B.n753 B.n752 10.6151
R2400 B.n755 B.n753 10.6151
R2401 B.n756 B.n755 10.6151
R2402 B.n757 B.n756 10.6151
R2403 B.n758 B.n757 10.6151
R2404 B.n760 B.n758 10.6151
R2405 B.n761 B.n760 10.6151
R2406 B.n762 B.n761 10.6151
R2407 B.n763 B.n762 10.6151
R2408 B.n1064 B.n1 10.6151
R2409 B.n1064 B.n1063 10.6151
R2410 B.n1063 B.n1062 10.6151
R2411 B.n1062 B.n10 10.6151
R2412 B.n1056 B.n10 10.6151
R2413 B.n1056 B.n1055 10.6151
R2414 B.n1055 B.n1054 10.6151
R2415 B.n1054 B.n18 10.6151
R2416 B.n1048 B.n18 10.6151
R2417 B.n1048 B.n1047 10.6151
R2418 B.n1047 B.n1046 10.6151
R2419 B.n1046 B.n25 10.6151
R2420 B.n1040 B.n25 10.6151
R2421 B.n1040 B.n1039 10.6151
R2422 B.n1039 B.n1038 10.6151
R2423 B.n1038 B.n32 10.6151
R2424 B.n1032 B.n32 10.6151
R2425 B.n1032 B.n1031 10.6151
R2426 B.n1031 B.n1030 10.6151
R2427 B.n1030 B.n39 10.6151
R2428 B.n1024 B.n39 10.6151
R2429 B.n1024 B.n1023 10.6151
R2430 B.n1023 B.n1022 10.6151
R2431 B.n1022 B.n46 10.6151
R2432 B.n1016 B.n46 10.6151
R2433 B.n1016 B.n1015 10.6151
R2434 B.n1015 B.n1014 10.6151
R2435 B.n1014 B.n53 10.6151
R2436 B.n1008 B.n53 10.6151
R2437 B.n1008 B.n1007 10.6151
R2438 B.n1007 B.n1006 10.6151
R2439 B.n1006 B.n60 10.6151
R2440 B.n1000 B.n60 10.6151
R2441 B.n1000 B.n999 10.6151
R2442 B.n999 B.n998 10.6151
R2443 B.n998 B.n67 10.6151
R2444 B.n992 B.n67 10.6151
R2445 B.n992 B.n991 10.6151
R2446 B.n991 B.n990 10.6151
R2447 B.n990 B.n74 10.6151
R2448 B.n984 B.n74 10.6151
R2449 B.n984 B.n983 10.6151
R2450 B.n983 B.n982 10.6151
R2451 B.n982 B.n81 10.6151
R2452 B.n976 B.n81 10.6151
R2453 B.n976 B.n975 10.6151
R2454 B.n975 B.n974 10.6151
R2455 B.n974 B.n88 10.6151
R2456 B.n968 B.n88 10.6151
R2457 B.n968 B.n967 10.6151
R2458 B.n967 B.n966 10.6151
R2459 B.n966 B.n95 10.6151
R2460 B.n960 B.n95 10.6151
R2461 B.n960 B.n959 10.6151
R2462 B.n959 B.n958 10.6151
R2463 B.n958 B.n102 10.6151
R2464 B.n952 B.n102 10.6151
R2465 B.n951 B.n950 10.6151
R2466 B.n950 B.n109 10.6151
R2467 B.n944 B.n109 10.6151
R2468 B.n944 B.n943 10.6151
R2469 B.n943 B.n942 10.6151
R2470 B.n942 B.n111 10.6151
R2471 B.n936 B.n111 10.6151
R2472 B.n936 B.n935 10.6151
R2473 B.n935 B.n934 10.6151
R2474 B.n934 B.n113 10.6151
R2475 B.n928 B.n113 10.6151
R2476 B.n928 B.n927 10.6151
R2477 B.n927 B.n926 10.6151
R2478 B.n926 B.n115 10.6151
R2479 B.n920 B.n115 10.6151
R2480 B.n920 B.n919 10.6151
R2481 B.n919 B.n918 10.6151
R2482 B.n918 B.n117 10.6151
R2483 B.n912 B.n117 10.6151
R2484 B.n912 B.n911 10.6151
R2485 B.n911 B.n910 10.6151
R2486 B.n910 B.n119 10.6151
R2487 B.n904 B.n119 10.6151
R2488 B.n904 B.n903 10.6151
R2489 B.n903 B.n902 10.6151
R2490 B.n902 B.n121 10.6151
R2491 B.n896 B.n121 10.6151
R2492 B.n896 B.n895 10.6151
R2493 B.n895 B.n894 10.6151
R2494 B.n894 B.n123 10.6151
R2495 B.n888 B.n123 10.6151
R2496 B.n888 B.n887 10.6151
R2497 B.n887 B.n886 10.6151
R2498 B.n886 B.n125 10.6151
R2499 B.n880 B.n125 10.6151
R2500 B.n880 B.n879 10.6151
R2501 B.n879 B.n878 10.6151
R2502 B.n878 B.n127 10.6151
R2503 B.n872 B.n127 10.6151
R2504 B.n872 B.n871 10.6151
R2505 B.n871 B.n870 10.6151
R2506 B.n866 B.n865 10.6151
R2507 B.n865 B.n133 10.6151
R2508 B.n860 B.n133 10.6151
R2509 B.n860 B.n859 10.6151
R2510 B.n859 B.n858 10.6151
R2511 B.n858 B.n135 10.6151
R2512 B.n852 B.n135 10.6151
R2513 B.n852 B.n851 10.6151
R2514 B.n851 B.n850 10.6151
R2515 B.n846 B.n845 10.6151
R2516 B.n845 B.n141 10.6151
R2517 B.n840 B.n141 10.6151
R2518 B.n840 B.n839 10.6151
R2519 B.n839 B.n838 10.6151
R2520 B.n838 B.n143 10.6151
R2521 B.n832 B.n143 10.6151
R2522 B.n832 B.n831 10.6151
R2523 B.n831 B.n830 10.6151
R2524 B.n830 B.n145 10.6151
R2525 B.n824 B.n145 10.6151
R2526 B.n824 B.n823 10.6151
R2527 B.n823 B.n822 10.6151
R2528 B.n822 B.n147 10.6151
R2529 B.n816 B.n147 10.6151
R2530 B.n816 B.n815 10.6151
R2531 B.n815 B.n814 10.6151
R2532 B.n814 B.n149 10.6151
R2533 B.n808 B.n149 10.6151
R2534 B.n808 B.n807 10.6151
R2535 B.n807 B.n806 10.6151
R2536 B.n806 B.n151 10.6151
R2537 B.n800 B.n151 10.6151
R2538 B.n800 B.n799 10.6151
R2539 B.n799 B.n798 10.6151
R2540 B.n798 B.n153 10.6151
R2541 B.n792 B.n153 10.6151
R2542 B.n792 B.n791 10.6151
R2543 B.n791 B.n790 10.6151
R2544 B.n790 B.n155 10.6151
R2545 B.n784 B.n155 10.6151
R2546 B.n784 B.n783 10.6151
R2547 B.n783 B.n782 10.6151
R2548 B.n782 B.n157 10.6151
R2549 B.n776 B.n157 10.6151
R2550 B.n776 B.n775 10.6151
R2551 B.n775 B.n774 10.6151
R2552 B.n774 B.n159 10.6151
R2553 B.n768 B.n159 10.6151
R2554 B.n768 B.n767 10.6151
R2555 B.n767 B.n766 10.6151
R2556 B.n301 B.n297 9.36635
R2557 B.n411 B.n410 9.36635
R2558 B.n870 B.n131 9.36635
R2559 B.n846 B.n139 9.36635
R2560 B.n1072 B.n0 8.11757
R2561 B.n1072 B.n1 8.11757
R2562 B.n630 B.t3 3.15146
R2563 B.n1028 B.t4 3.15146
R2564 B.n429 B.n301 1.24928
R2565 B.n412 B.n411 1.24928
R2566 B.n866 B.n131 1.24928
R2567 B.n850 B.n139 1.24928
R2568 VN.n42 VN.n41 161.3
R2569 VN.n40 VN.n23 161.3
R2570 VN.n39 VN.n38 161.3
R2571 VN.n37 VN.n24 161.3
R2572 VN.n36 VN.n35 161.3
R2573 VN.n34 VN.n25 161.3
R2574 VN.n33 VN.n32 161.3
R2575 VN.n31 VN.n26 161.3
R2576 VN.n30 VN.n29 161.3
R2577 VN.n20 VN.n19 161.3
R2578 VN.n18 VN.n1 161.3
R2579 VN.n17 VN.n16 161.3
R2580 VN.n15 VN.n2 161.3
R2581 VN.n14 VN.n13 161.3
R2582 VN.n12 VN.n3 161.3
R2583 VN.n11 VN.n10 161.3
R2584 VN.n9 VN.n4 161.3
R2585 VN.n8 VN.n7 161.3
R2586 VN.n27 VN.t4 106.707
R2587 VN.n5 VN.t5 106.707
R2588 VN.n21 VN.n0 87.7864
R2589 VN.n43 VN.n22 87.7864
R2590 VN.n6 VN.t2 73.9395
R2591 VN.n0 VN.t3 73.9395
R2592 VN.n28 VN.t0 73.9395
R2593 VN.n22 VN.t1 73.9395
R2594 VN.n6 VN.n5 63.107
R2595 VN.n28 VN.n27 63.107
R2596 VN VN.n43 54.4375
R2597 VN.n13 VN.n12 50.2647
R2598 VN.n35 VN.n34 50.2647
R2599 VN.n13 VN.n2 30.8893
R2600 VN.n35 VN.n24 30.8893
R2601 VN.n7 VN.n4 24.5923
R2602 VN.n11 VN.n4 24.5923
R2603 VN.n12 VN.n11 24.5923
R2604 VN.n17 VN.n2 24.5923
R2605 VN.n18 VN.n17 24.5923
R2606 VN.n19 VN.n18 24.5923
R2607 VN.n34 VN.n33 24.5923
R2608 VN.n33 VN.n26 24.5923
R2609 VN.n29 VN.n26 24.5923
R2610 VN.n41 VN.n40 24.5923
R2611 VN.n40 VN.n39 24.5923
R2612 VN.n39 VN.n24 24.5923
R2613 VN.n7 VN.n6 12.2964
R2614 VN.n29 VN.n28 12.2964
R2615 VN.n8 VN.n5 2.46667
R2616 VN.n30 VN.n27 2.46667
R2617 VN.n19 VN.n0 2.45968
R2618 VN.n41 VN.n22 2.45968
R2619 VN.n43 VN.n42 0.354861
R2620 VN.n21 VN.n20 0.354861
R2621 VN VN.n21 0.267071
R2622 VN.n42 VN.n23 0.189894
R2623 VN.n38 VN.n23 0.189894
R2624 VN.n38 VN.n37 0.189894
R2625 VN.n37 VN.n36 0.189894
R2626 VN.n36 VN.n25 0.189894
R2627 VN.n32 VN.n25 0.189894
R2628 VN.n32 VN.n31 0.189894
R2629 VN.n31 VN.n30 0.189894
R2630 VN.n9 VN.n8 0.189894
R2631 VN.n10 VN.n9 0.189894
R2632 VN.n10 VN.n3 0.189894
R2633 VN.n14 VN.n3 0.189894
R2634 VN.n15 VN.n14 0.189894
R2635 VN.n16 VN.n15 0.189894
R2636 VN.n16 VN.n1 0.189894
R2637 VN.n20 VN.n1 0.189894
R2638 VDD2.n127 VDD2.n67 289.615
R2639 VDD2.n60 VDD2.n0 289.615
R2640 VDD2.n128 VDD2.n127 185
R2641 VDD2.n126 VDD2.n125 185
R2642 VDD2.n71 VDD2.n70 185
R2643 VDD2.n120 VDD2.n119 185
R2644 VDD2.n118 VDD2.n117 185
R2645 VDD2.n75 VDD2.n74 185
R2646 VDD2.n112 VDD2.n111 185
R2647 VDD2.n110 VDD2.n77 185
R2648 VDD2.n109 VDD2.n108 185
R2649 VDD2.n80 VDD2.n78 185
R2650 VDD2.n103 VDD2.n102 185
R2651 VDD2.n101 VDD2.n100 185
R2652 VDD2.n84 VDD2.n83 185
R2653 VDD2.n95 VDD2.n94 185
R2654 VDD2.n93 VDD2.n92 185
R2655 VDD2.n88 VDD2.n87 185
R2656 VDD2.n20 VDD2.n19 185
R2657 VDD2.n25 VDD2.n24 185
R2658 VDD2.n27 VDD2.n26 185
R2659 VDD2.n16 VDD2.n15 185
R2660 VDD2.n33 VDD2.n32 185
R2661 VDD2.n35 VDD2.n34 185
R2662 VDD2.n12 VDD2.n11 185
R2663 VDD2.n42 VDD2.n41 185
R2664 VDD2.n43 VDD2.n10 185
R2665 VDD2.n45 VDD2.n44 185
R2666 VDD2.n8 VDD2.n7 185
R2667 VDD2.n51 VDD2.n50 185
R2668 VDD2.n53 VDD2.n52 185
R2669 VDD2.n4 VDD2.n3 185
R2670 VDD2.n59 VDD2.n58 185
R2671 VDD2.n61 VDD2.n60 185
R2672 VDD2.n89 VDD2.t4 149.524
R2673 VDD2.n21 VDD2.t0 149.524
R2674 VDD2.n127 VDD2.n126 104.615
R2675 VDD2.n126 VDD2.n70 104.615
R2676 VDD2.n119 VDD2.n70 104.615
R2677 VDD2.n119 VDD2.n118 104.615
R2678 VDD2.n118 VDD2.n74 104.615
R2679 VDD2.n111 VDD2.n74 104.615
R2680 VDD2.n111 VDD2.n110 104.615
R2681 VDD2.n110 VDD2.n109 104.615
R2682 VDD2.n109 VDD2.n78 104.615
R2683 VDD2.n102 VDD2.n78 104.615
R2684 VDD2.n102 VDD2.n101 104.615
R2685 VDD2.n101 VDD2.n83 104.615
R2686 VDD2.n94 VDD2.n83 104.615
R2687 VDD2.n94 VDD2.n93 104.615
R2688 VDD2.n93 VDD2.n87 104.615
R2689 VDD2.n25 VDD2.n19 104.615
R2690 VDD2.n26 VDD2.n25 104.615
R2691 VDD2.n26 VDD2.n15 104.615
R2692 VDD2.n33 VDD2.n15 104.615
R2693 VDD2.n34 VDD2.n33 104.615
R2694 VDD2.n34 VDD2.n11 104.615
R2695 VDD2.n42 VDD2.n11 104.615
R2696 VDD2.n43 VDD2.n42 104.615
R2697 VDD2.n44 VDD2.n43 104.615
R2698 VDD2.n44 VDD2.n7 104.615
R2699 VDD2.n51 VDD2.n7 104.615
R2700 VDD2.n52 VDD2.n51 104.615
R2701 VDD2.n52 VDD2.n3 104.615
R2702 VDD2.n59 VDD2.n3 104.615
R2703 VDD2.n60 VDD2.n59 104.615
R2704 VDD2.n66 VDD2.n65 63.9148
R2705 VDD2 VDD2.n133 63.9119
R2706 VDD2.n66 VDD2.n64 52.7526
R2707 VDD2.t4 VDD2.n87 52.3082
R2708 VDD2.t0 VDD2.n19 52.3082
R2709 VDD2.n132 VDD2.n131 50.0278
R2710 VDD2.n132 VDD2.n66 46.2627
R2711 VDD2.n112 VDD2.n77 13.1884
R2712 VDD2.n45 VDD2.n10 13.1884
R2713 VDD2.n113 VDD2.n75 12.8005
R2714 VDD2.n108 VDD2.n79 12.8005
R2715 VDD2.n41 VDD2.n40 12.8005
R2716 VDD2.n46 VDD2.n8 12.8005
R2717 VDD2.n117 VDD2.n116 12.0247
R2718 VDD2.n107 VDD2.n80 12.0247
R2719 VDD2.n39 VDD2.n12 12.0247
R2720 VDD2.n50 VDD2.n49 12.0247
R2721 VDD2.n120 VDD2.n73 11.249
R2722 VDD2.n104 VDD2.n103 11.249
R2723 VDD2.n36 VDD2.n35 11.249
R2724 VDD2.n53 VDD2.n6 11.249
R2725 VDD2.n121 VDD2.n71 10.4732
R2726 VDD2.n100 VDD2.n82 10.4732
R2727 VDD2.n32 VDD2.n14 10.4732
R2728 VDD2.n54 VDD2.n4 10.4732
R2729 VDD2.n89 VDD2.n88 10.2747
R2730 VDD2.n21 VDD2.n20 10.2747
R2731 VDD2.n125 VDD2.n124 9.69747
R2732 VDD2.n99 VDD2.n84 9.69747
R2733 VDD2.n31 VDD2.n16 9.69747
R2734 VDD2.n58 VDD2.n57 9.69747
R2735 VDD2.n131 VDD2.n130 9.45567
R2736 VDD2.n64 VDD2.n63 9.45567
R2737 VDD2.n91 VDD2.n90 9.3005
R2738 VDD2.n86 VDD2.n85 9.3005
R2739 VDD2.n97 VDD2.n96 9.3005
R2740 VDD2.n99 VDD2.n98 9.3005
R2741 VDD2.n82 VDD2.n81 9.3005
R2742 VDD2.n105 VDD2.n104 9.3005
R2743 VDD2.n107 VDD2.n106 9.3005
R2744 VDD2.n79 VDD2.n76 9.3005
R2745 VDD2.n130 VDD2.n129 9.3005
R2746 VDD2.n69 VDD2.n68 9.3005
R2747 VDD2.n124 VDD2.n123 9.3005
R2748 VDD2.n122 VDD2.n121 9.3005
R2749 VDD2.n73 VDD2.n72 9.3005
R2750 VDD2.n116 VDD2.n115 9.3005
R2751 VDD2.n114 VDD2.n113 9.3005
R2752 VDD2.n63 VDD2.n62 9.3005
R2753 VDD2.n2 VDD2.n1 9.3005
R2754 VDD2.n57 VDD2.n56 9.3005
R2755 VDD2.n55 VDD2.n54 9.3005
R2756 VDD2.n6 VDD2.n5 9.3005
R2757 VDD2.n49 VDD2.n48 9.3005
R2758 VDD2.n47 VDD2.n46 9.3005
R2759 VDD2.n23 VDD2.n22 9.3005
R2760 VDD2.n18 VDD2.n17 9.3005
R2761 VDD2.n29 VDD2.n28 9.3005
R2762 VDD2.n31 VDD2.n30 9.3005
R2763 VDD2.n14 VDD2.n13 9.3005
R2764 VDD2.n37 VDD2.n36 9.3005
R2765 VDD2.n39 VDD2.n38 9.3005
R2766 VDD2.n40 VDD2.n9 9.3005
R2767 VDD2.n128 VDD2.n69 8.92171
R2768 VDD2.n96 VDD2.n95 8.92171
R2769 VDD2.n28 VDD2.n27 8.92171
R2770 VDD2.n61 VDD2.n2 8.92171
R2771 VDD2.n129 VDD2.n67 8.14595
R2772 VDD2.n92 VDD2.n86 8.14595
R2773 VDD2.n24 VDD2.n18 8.14595
R2774 VDD2.n62 VDD2.n0 8.14595
R2775 VDD2.n91 VDD2.n88 7.3702
R2776 VDD2.n23 VDD2.n20 7.3702
R2777 VDD2.n131 VDD2.n67 5.81868
R2778 VDD2.n92 VDD2.n91 5.81868
R2779 VDD2.n24 VDD2.n23 5.81868
R2780 VDD2.n64 VDD2.n0 5.81868
R2781 VDD2.n129 VDD2.n128 5.04292
R2782 VDD2.n95 VDD2.n86 5.04292
R2783 VDD2.n27 VDD2.n18 5.04292
R2784 VDD2.n62 VDD2.n61 5.04292
R2785 VDD2.n125 VDD2.n69 4.26717
R2786 VDD2.n96 VDD2.n84 4.26717
R2787 VDD2.n28 VDD2.n16 4.26717
R2788 VDD2.n58 VDD2.n2 4.26717
R2789 VDD2.n124 VDD2.n71 3.49141
R2790 VDD2.n100 VDD2.n99 3.49141
R2791 VDD2.n32 VDD2.n31 3.49141
R2792 VDD2.n57 VDD2.n4 3.49141
R2793 VDD2.n90 VDD2.n89 2.84303
R2794 VDD2.n22 VDD2.n21 2.84303
R2795 VDD2 VDD2.n132 2.83886
R2796 VDD2.n121 VDD2.n120 2.71565
R2797 VDD2.n103 VDD2.n82 2.71565
R2798 VDD2.n35 VDD2.n14 2.71565
R2799 VDD2.n54 VDD2.n53 2.71565
R2800 VDD2.n117 VDD2.n73 1.93989
R2801 VDD2.n104 VDD2.n80 1.93989
R2802 VDD2.n36 VDD2.n12 1.93989
R2803 VDD2.n50 VDD2.n6 1.93989
R2804 VDD2.n133 VDD2.t5 1.62612
R2805 VDD2.n133 VDD2.t1 1.62612
R2806 VDD2.n65 VDD2.t3 1.62612
R2807 VDD2.n65 VDD2.t2 1.62612
R2808 VDD2.n116 VDD2.n75 1.16414
R2809 VDD2.n108 VDD2.n107 1.16414
R2810 VDD2.n41 VDD2.n39 1.16414
R2811 VDD2.n49 VDD2.n8 1.16414
R2812 VDD2.n113 VDD2.n112 0.388379
R2813 VDD2.n79 VDD2.n77 0.388379
R2814 VDD2.n40 VDD2.n10 0.388379
R2815 VDD2.n46 VDD2.n45 0.388379
R2816 VDD2.n130 VDD2.n68 0.155672
R2817 VDD2.n123 VDD2.n68 0.155672
R2818 VDD2.n123 VDD2.n122 0.155672
R2819 VDD2.n122 VDD2.n72 0.155672
R2820 VDD2.n115 VDD2.n72 0.155672
R2821 VDD2.n115 VDD2.n114 0.155672
R2822 VDD2.n114 VDD2.n76 0.155672
R2823 VDD2.n106 VDD2.n76 0.155672
R2824 VDD2.n106 VDD2.n105 0.155672
R2825 VDD2.n105 VDD2.n81 0.155672
R2826 VDD2.n98 VDD2.n81 0.155672
R2827 VDD2.n98 VDD2.n97 0.155672
R2828 VDD2.n97 VDD2.n85 0.155672
R2829 VDD2.n90 VDD2.n85 0.155672
R2830 VDD2.n22 VDD2.n17 0.155672
R2831 VDD2.n29 VDD2.n17 0.155672
R2832 VDD2.n30 VDD2.n29 0.155672
R2833 VDD2.n30 VDD2.n13 0.155672
R2834 VDD2.n37 VDD2.n13 0.155672
R2835 VDD2.n38 VDD2.n37 0.155672
R2836 VDD2.n38 VDD2.n9 0.155672
R2837 VDD2.n47 VDD2.n9 0.155672
R2838 VDD2.n48 VDD2.n47 0.155672
R2839 VDD2.n48 VDD2.n5 0.155672
R2840 VDD2.n55 VDD2.n5 0.155672
R2841 VDD2.n56 VDD2.n55 0.155672
R2842 VDD2.n56 VDD2.n1 0.155672
R2843 VDD2.n63 VDD2.n1 0.155672
C0 VTAIL VDD2 8.366349f
C1 VN VDD2 7.29082f
C2 VDD1 VDD2 1.94155f
C3 VP VDD2 0.574169f
C4 VTAIL VN 7.77219f
C5 VTAIL VDD1 8.3053f
C6 VDD1 VN 0.152923f
C7 VTAIL VP 7.787069f
C8 VP VN 8.28347f
C9 VDD1 VP 7.70967f
C10 VDD2 B 7.067491f
C11 VDD1 B 7.260428f
C12 VTAIL B 8.748857f
C13 VN B 16.92957f
C14 VP B 15.658037f
C15 VDD2.n0 B 0.030958f
C16 VDD2.n1 B 0.021408f
C17 VDD2.n2 B 0.011504f
C18 VDD2.n3 B 0.027191f
C19 VDD2.n4 B 0.01218f
C20 VDD2.n5 B 0.021408f
C21 VDD2.n6 B 0.011504f
C22 VDD2.n7 B 0.027191f
C23 VDD2.n8 B 0.01218f
C24 VDD2.n9 B 0.021408f
C25 VDD2.n10 B 0.011842f
C26 VDD2.n11 B 0.027191f
C27 VDD2.n12 B 0.01218f
C28 VDD2.n13 B 0.021408f
C29 VDD2.n14 B 0.011504f
C30 VDD2.n15 B 0.027191f
C31 VDD2.n16 B 0.01218f
C32 VDD2.n17 B 0.021408f
C33 VDD2.n18 B 0.011504f
C34 VDD2.n19 B 0.020393f
C35 VDD2.n20 B 0.019222f
C36 VDD2.t0 B 0.045945f
C37 VDD2.n21 B 0.15583f
C38 VDD2.n22 B 1.09715f
C39 VDD2.n23 B 0.011504f
C40 VDD2.n24 B 0.01218f
C41 VDD2.n25 B 0.027191f
C42 VDD2.n26 B 0.027191f
C43 VDD2.n27 B 0.01218f
C44 VDD2.n28 B 0.011504f
C45 VDD2.n29 B 0.021408f
C46 VDD2.n30 B 0.021408f
C47 VDD2.n31 B 0.011504f
C48 VDD2.n32 B 0.01218f
C49 VDD2.n33 B 0.027191f
C50 VDD2.n34 B 0.027191f
C51 VDD2.n35 B 0.01218f
C52 VDD2.n36 B 0.011504f
C53 VDD2.n37 B 0.021408f
C54 VDD2.n38 B 0.021408f
C55 VDD2.n39 B 0.011504f
C56 VDD2.n40 B 0.011504f
C57 VDD2.n41 B 0.01218f
C58 VDD2.n42 B 0.027191f
C59 VDD2.n43 B 0.027191f
C60 VDD2.n44 B 0.027191f
C61 VDD2.n45 B 0.011842f
C62 VDD2.n46 B 0.011504f
C63 VDD2.n47 B 0.021408f
C64 VDD2.n48 B 0.021408f
C65 VDD2.n49 B 0.011504f
C66 VDD2.n50 B 0.01218f
C67 VDD2.n51 B 0.027191f
C68 VDD2.n52 B 0.027191f
C69 VDD2.n53 B 0.01218f
C70 VDD2.n54 B 0.011504f
C71 VDD2.n55 B 0.021408f
C72 VDD2.n56 B 0.021408f
C73 VDD2.n57 B 0.011504f
C74 VDD2.n58 B 0.01218f
C75 VDD2.n59 B 0.027191f
C76 VDD2.n60 B 0.060396f
C77 VDD2.n61 B 0.01218f
C78 VDD2.n62 B 0.011504f
C79 VDD2.n63 B 0.051239f
C80 VDD2.n64 B 0.060673f
C81 VDD2.t3 B 0.206054f
C82 VDD2.t2 B 0.206054f
C83 VDD2.n65 B 1.84542f
C84 VDD2.n66 B 2.8095f
C85 VDD2.n67 B 0.030958f
C86 VDD2.n68 B 0.021408f
C87 VDD2.n69 B 0.011504f
C88 VDD2.n70 B 0.027191f
C89 VDD2.n71 B 0.01218f
C90 VDD2.n72 B 0.021408f
C91 VDD2.n73 B 0.011504f
C92 VDD2.n74 B 0.027191f
C93 VDD2.n75 B 0.01218f
C94 VDD2.n76 B 0.021408f
C95 VDD2.n77 B 0.011842f
C96 VDD2.n78 B 0.027191f
C97 VDD2.n79 B 0.011504f
C98 VDD2.n80 B 0.01218f
C99 VDD2.n81 B 0.021408f
C100 VDD2.n82 B 0.011504f
C101 VDD2.n83 B 0.027191f
C102 VDD2.n84 B 0.01218f
C103 VDD2.n85 B 0.021408f
C104 VDD2.n86 B 0.011504f
C105 VDD2.n87 B 0.020393f
C106 VDD2.n88 B 0.019222f
C107 VDD2.t4 B 0.045945f
C108 VDD2.n89 B 0.15583f
C109 VDD2.n90 B 1.09715f
C110 VDD2.n91 B 0.011504f
C111 VDD2.n92 B 0.01218f
C112 VDD2.n93 B 0.027191f
C113 VDD2.n94 B 0.027191f
C114 VDD2.n95 B 0.01218f
C115 VDD2.n96 B 0.011504f
C116 VDD2.n97 B 0.021408f
C117 VDD2.n98 B 0.021408f
C118 VDD2.n99 B 0.011504f
C119 VDD2.n100 B 0.01218f
C120 VDD2.n101 B 0.027191f
C121 VDD2.n102 B 0.027191f
C122 VDD2.n103 B 0.01218f
C123 VDD2.n104 B 0.011504f
C124 VDD2.n105 B 0.021408f
C125 VDD2.n106 B 0.021408f
C126 VDD2.n107 B 0.011504f
C127 VDD2.n108 B 0.01218f
C128 VDD2.n109 B 0.027191f
C129 VDD2.n110 B 0.027191f
C130 VDD2.n111 B 0.027191f
C131 VDD2.n112 B 0.011842f
C132 VDD2.n113 B 0.011504f
C133 VDD2.n114 B 0.021408f
C134 VDD2.n115 B 0.021408f
C135 VDD2.n116 B 0.011504f
C136 VDD2.n117 B 0.01218f
C137 VDD2.n118 B 0.027191f
C138 VDD2.n119 B 0.027191f
C139 VDD2.n120 B 0.01218f
C140 VDD2.n121 B 0.011504f
C141 VDD2.n122 B 0.021408f
C142 VDD2.n123 B 0.021408f
C143 VDD2.n124 B 0.011504f
C144 VDD2.n125 B 0.01218f
C145 VDD2.n126 B 0.027191f
C146 VDD2.n127 B 0.060396f
C147 VDD2.n128 B 0.01218f
C148 VDD2.n129 B 0.011504f
C149 VDD2.n130 B 0.051239f
C150 VDD2.n131 B 0.048773f
C151 VDD2.n132 B 2.52696f
C152 VDD2.t5 B 0.206054f
C153 VDD2.t1 B 0.206054f
C154 VDD2.n133 B 1.84539f
C155 VN.t3 B 2.33317f
C156 VN.n0 B 0.884168f
C157 VN.n1 B 0.017702f
C158 VN.n2 B 0.035271f
C159 VN.n3 B 0.017702f
C160 VN.n4 B 0.032827f
C161 VN.t5 B 2.62771f
C162 VN.n5 B 0.836062f
C163 VN.t2 B 2.33317f
C164 VN.n6 B 0.879959f
C165 VN.n7 B 0.024724f
C166 VN.n8 B 0.231309f
C167 VN.n9 B 0.017702f
C168 VN.n10 B 0.017702f
C169 VN.n11 B 0.032827f
C170 VN.n12 B 0.03233f
C171 VN.n13 B 0.01669f
C172 VN.n14 B 0.017702f
C173 VN.n15 B 0.017702f
C174 VN.n16 B 0.017702f
C175 VN.n17 B 0.032827f
C176 VN.n18 B 0.032827f
C177 VN.n19 B 0.018242f
C178 VN.n20 B 0.028566f
C179 VN.n21 B 0.056217f
C180 VN.t1 B 2.33317f
C181 VN.n22 B 0.884168f
C182 VN.n23 B 0.017702f
C183 VN.n24 B 0.035271f
C184 VN.n25 B 0.017702f
C185 VN.n26 B 0.032827f
C186 VN.t4 B 2.62771f
C187 VN.n27 B 0.836062f
C188 VN.t0 B 2.33317f
C189 VN.n28 B 0.879959f
C190 VN.n29 B 0.024724f
C191 VN.n30 B 0.231309f
C192 VN.n31 B 0.017702f
C193 VN.n32 B 0.017702f
C194 VN.n33 B 0.032827f
C195 VN.n34 B 0.03233f
C196 VN.n35 B 0.01669f
C197 VN.n36 B 0.017702f
C198 VN.n37 B 0.017702f
C199 VN.n38 B 0.017702f
C200 VN.n39 B 0.032827f
C201 VN.n40 B 0.032827f
C202 VN.n41 B 0.018242f
C203 VN.n42 B 0.028566f
C204 VN.n43 B 1.15212f
C205 VTAIL.t2 B 0.23714f
C206 VTAIL.t4 B 0.23714f
C207 VTAIL.n0 B 2.04456f
C208 VTAIL.n1 B 0.503706f
C209 VTAIL.n2 B 0.035628f
C210 VTAIL.n3 B 0.024638f
C211 VTAIL.n4 B 0.013239f
C212 VTAIL.n5 B 0.031293f
C213 VTAIL.n6 B 0.014018f
C214 VTAIL.n7 B 0.024638f
C215 VTAIL.n8 B 0.013239f
C216 VTAIL.n9 B 0.031293f
C217 VTAIL.n10 B 0.014018f
C218 VTAIL.n11 B 0.024638f
C219 VTAIL.n12 B 0.013629f
C220 VTAIL.n13 B 0.031293f
C221 VTAIL.n14 B 0.014018f
C222 VTAIL.n15 B 0.024638f
C223 VTAIL.n16 B 0.013239f
C224 VTAIL.n17 B 0.031293f
C225 VTAIL.n18 B 0.014018f
C226 VTAIL.n19 B 0.024638f
C227 VTAIL.n20 B 0.013239f
C228 VTAIL.n21 B 0.02347f
C229 VTAIL.n22 B 0.022122f
C230 VTAIL.t10 B 0.052876f
C231 VTAIL.n23 B 0.17934f
C232 VTAIL.n24 B 1.26267f
C233 VTAIL.n25 B 0.013239f
C234 VTAIL.n26 B 0.014018f
C235 VTAIL.n27 B 0.031293f
C236 VTAIL.n28 B 0.031293f
C237 VTAIL.n29 B 0.014018f
C238 VTAIL.n30 B 0.013239f
C239 VTAIL.n31 B 0.024638f
C240 VTAIL.n32 B 0.024638f
C241 VTAIL.n33 B 0.013239f
C242 VTAIL.n34 B 0.014018f
C243 VTAIL.n35 B 0.031293f
C244 VTAIL.n36 B 0.031293f
C245 VTAIL.n37 B 0.014018f
C246 VTAIL.n38 B 0.013239f
C247 VTAIL.n39 B 0.024638f
C248 VTAIL.n40 B 0.024638f
C249 VTAIL.n41 B 0.013239f
C250 VTAIL.n42 B 0.013239f
C251 VTAIL.n43 B 0.014018f
C252 VTAIL.n44 B 0.031293f
C253 VTAIL.n45 B 0.031293f
C254 VTAIL.n46 B 0.031293f
C255 VTAIL.n47 B 0.013629f
C256 VTAIL.n48 B 0.013239f
C257 VTAIL.n49 B 0.024638f
C258 VTAIL.n50 B 0.024638f
C259 VTAIL.n51 B 0.013239f
C260 VTAIL.n52 B 0.014018f
C261 VTAIL.n53 B 0.031293f
C262 VTAIL.n54 B 0.031293f
C263 VTAIL.n55 B 0.014018f
C264 VTAIL.n56 B 0.013239f
C265 VTAIL.n57 B 0.024638f
C266 VTAIL.n58 B 0.024638f
C267 VTAIL.n59 B 0.013239f
C268 VTAIL.n60 B 0.014018f
C269 VTAIL.n61 B 0.031293f
C270 VTAIL.n62 B 0.069508f
C271 VTAIL.n63 B 0.014018f
C272 VTAIL.n64 B 0.013239f
C273 VTAIL.n65 B 0.058969f
C274 VTAIL.n66 B 0.039135f
C275 VTAIL.n67 B 0.500913f
C276 VTAIL.t6 B 0.23714f
C277 VTAIL.t11 B 0.23714f
C278 VTAIL.n68 B 2.04456f
C279 VTAIL.n69 B 2.29219f
C280 VTAIL.t5 B 0.23714f
C281 VTAIL.t3 B 0.23714f
C282 VTAIL.n70 B 2.04457f
C283 VTAIL.n71 B 2.29218f
C284 VTAIL.n72 B 0.035628f
C285 VTAIL.n73 B 0.024638f
C286 VTAIL.n74 B 0.013239f
C287 VTAIL.n75 B 0.031293f
C288 VTAIL.n76 B 0.014018f
C289 VTAIL.n77 B 0.024638f
C290 VTAIL.n78 B 0.013239f
C291 VTAIL.n79 B 0.031293f
C292 VTAIL.n80 B 0.014018f
C293 VTAIL.n81 B 0.024638f
C294 VTAIL.n82 B 0.013629f
C295 VTAIL.n83 B 0.031293f
C296 VTAIL.n84 B 0.013239f
C297 VTAIL.n85 B 0.014018f
C298 VTAIL.n86 B 0.024638f
C299 VTAIL.n87 B 0.013239f
C300 VTAIL.n88 B 0.031293f
C301 VTAIL.n89 B 0.014018f
C302 VTAIL.n90 B 0.024638f
C303 VTAIL.n91 B 0.013239f
C304 VTAIL.n92 B 0.02347f
C305 VTAIL.n93 B 0.022122f
C306 VTAIL.t0 B 0.052876f
C307 VTAIL.n94 B 0.17934f
C308 VTAIL.n95 B 1.26267f
C309 VTAIL.n96 B 0.013239f
C310 VTAIL.n97 B 0.014018f
C311 VTAIL.n98 B 0.031293f
C312 VTAIL.n99 B 0.031293f
C313 VTAIL.n100 B 0.014018f
C314 VTAIL.n101 B 0.013239f
C315 VTAIL.n102 B 0.024638f
C316 VTAIL.n103 B 0.024638f
C317 VTAIL.n104 B 0.013239f
C318 VTAIL.n105 B 0.014018f
C319 VTAIL.n106 B 0.031293f
C320 VTAIL.n107 B 0.031293f
C321 VTAIL.n108 B 0.014018f
C322 VTAIL.n109 B 0.013239f
C323 VTAIL.n110 B 0.024638f
C324 VTAIL.n111 B 0.024638f
C325 VTAIL.n112 B 0.013239f
C326 VTAIL.n113 B 0.014018f
C327 VTAIL.n114 B 0.031293f
C328 VTAIL.n115 B 0.031293f
C329 VTAIL.n116 B 0.031293f
C330 VTAIL.n117 B 0.013629f
C331 VTAIL.n118 B 0.013239f
C332 VTAIL.n119 B 0.024638f
C333 VTAIL.n120 B 0.024638f
C334 VTAIL.n121 B 0.013239f
C335 VTAIL.n122 B 0.014018f
C336 VTAIL.n123 B 0.031293f
C337 VTAIL.n124 B 0.031293f
C338 VTAIL.n125 B 0.014018f
C339 VTAIL.n126 B 0.013239f
C340 VTAIL.n127 B 0.024638f
C341 VTAIL.n128 B 0.024638f
C342 VTAIL.n129 B 0.013239f
C343 VTAIL.n130 B 0.014018f
C344 VTAIL.n131 B 0.031293f
C345 VTAIL.n132 B 0.069508f
C346 VTAIL.n133 B 0.014018f
C347 VTAIL.n134 B 0.013239f
C348 VTAIL.n135 B 0.058969f
C349 VTAIL.n136 B 0.039135f
C350 VTAIL.n137 B 0.500913f
C351 VTAIL.t8 B 0.23714f
C352 VTAIL.t9 B 0.23714f
C353 VTAIL.n138 B 2.04457f
C354 VTAIL.n139 B 0.71979f
C355 VTAIL.n140 B 0.035628f
C356 VTAIL.n141 B 0.024638f
C357 VTAIL.n142 B 0.013239f
C358 VTAIL.n143 B 0.031293f
C359 VTAIL.n144 B 0.014018f
C360 VTAIL.n145 B 0.024638f
C361 VTAIL.n146 B 0.013239f
C362 VTAIL.n147 B 0.031293f
C363 VTAIL.n148 B 0.014018f
C364 VTAIL.n149 B 0.024638f
C365 VTAIL.n150 B 0.013629f
C366 VTAIL.n151 B 0.031293f
C367 VTAIL.n152 B 0.013239f
C368 VTAIL.n153 B 0.014018f
C369 VTAIL.n154 B 0.024638f
C370 VTAIL.n155 B 0.013239f
C371 VTAIL.n156 B 0.031293f
C372 VTAIL.n157 B 0.014018f
C373 VTAIL.n158 B 0.024638f
C374 VTAIL.n159 B 0.013239f
C375 VTAIL.n160 B 0.02347f
C376 VTAIL.n161 B 0.022122f
C377 VTAIL.t7 B 0.052876f
C378 VTAIL.n162 B 0.17934f
C379 VTAIL.n163 B 1.26267f
C380 VTAIL.n164 B 0.013239f
C381 VTAIL.n165 B 0.014018f
C382 VTAIL.n166 B 0.031293f
C383 VTAIL.n167 B 0.031293f
C384 VTAIL.n168 B 0.014018f
C385 VTAIL.n169 B 0.013239f
C386 VTAIL.n170 B 0.024638f
C387 VTAIL.n171 B 0.024638f
C388 VTAIL.n172 B 0.013239f
C389 VTAIL.n173 B 0.014018f
C390 VTAIL.n174 B 0.031293f
C391 VTAIL.n175 B 0.031293f
C392 VTAIL.n176 B 0.014018f
C393 VTAIL.n177 B 0.013239f
C394 VTAIL.n178 B 0.024638f
C395 VTAIL.n179 B 0.024638f
C396 VTAIL.n180 B 0.013239f
C397 VTAIL.n181 B 0.014018f
C398 VTAIL.n182 B 0.031293f
C399 VTAIL.n183 B 0.031293f
C400 VTAIL.n184 B 0.031293f
C401 VTAIL.n185 B 0.013629f
C402 VTAIL.n186 B 0.013239f
C403 VTAIL.n187 B 0.024638f
C404 VTAIL.n188 B 0.024638f
C405 VTAIL.n189 B 0.013239f
C406 VTAIL.n190 B 0.014018f
C407 VTAIL.n191 B 0.031293f
C408 VTAIL.n192 B 0.031293f
C409 VTAIL.n193 B 0.014018f
C410 VTAIL.n194 B 0.013239f
C411 VTAIL.n195 B 0.024638f
C412 VTAIL.n196 B 0.024638f
C413 VTAIL.n197 B 0.013239f
C414 VTAIL.n198 B 0.014018f
C415 VTAIL.n199 B 0.031293f
C416 VTAIL.n200 B 0.069508f
C417 VTAIL.n201 B 0.014018f
C418 VTAIL.n202 B 0.013239f
C419 VTAIL.n203 B 0.058969f
C420 VTAIL.n204 B 0.039135f
C421 VTAIL.n205 B 1.77902f
C422 VTAIL.n206 B 0.035628f
C423 VTAIL.n207 B 0.024638f
C424 VTAIL.n208 B 0.013239f
C425 VTAIL.n209 B 0.031293f
C426 VTAIL.n210 B 0.014018f
C427 VTAIL.n211 B 0.024638f
C428 VTAIL.n212 B 0.013239f
C429 VTAIL.n213 B 0.031293f
C430 VTAIL.n214 B 0.014018f
C431 VTAIL.n215 B 0.024638f
C432 VTAIL.n216 B 0.013629f
C433 VTAIL.n217 B 0.031293f
C434 VTAIL.n218 B 0.014018f
C435 VTAIL.n219 B 0.024638f
C436 VTAIL.n220 B 0.013239f
C437 VTAIL.n221 B 0.031293f
C438 VTAIL.n222 B 0.014018f
C439 VTAIL.n223 B 0.024638f
C440 VTAIL.n224 B 0.013239f
C441 VTAIL.n225 B 0.02347f
C442 VTAIL.n226 B 0.022122f
C443 VTAIL.t1 B 0.052876f
C444 VTAIL.n227 B 0.17934f
C445 VTAIL.n228 B 1.26267f
C446 VTAIL.n229 B 0.013239f
C447 VTAIL.n230 B 0.014018f
C448 VTAIL.n231 B 0.031293f
C449 VTAIL.n232 B 0.031293f
C450 VTAIL.n233 B 0.014018f
C451 VTAIL.n234 B 0.013239f
C452 VTAIL.n235 B 0.024638f
C453 VTAIL.n236 B 0.024638f
C454 VTAIL.n237 B 0.013239f
C455 VTAIL.n238 B 0.014018f
C456 VTAIL.n239 B 0.031293f
C457 VTAIL.n240 B 0.031293f
C458 VTAIL.n241 B 0.014018f
C459 VTAIL.n242 B 0.013239f
C460 VTAIL.n243 B 0.024638f
C461 VTAIL.n244 B 0.024638f
C462 VTAIL.n245 B 0.013239f
C463 VTAIL.n246 B 0.013239f
C464 VTAIL.n247 B 0.014018f
C465 VTAIL.n248 B 0.031293f
C466 VTAIL.n249 B 0.031293f
C467 VTAIL.n250 B 0.031293f
C468 VTAIL.n251 B 0.013629f
C469 VTAIL.n252 B 0.013239f
C470 VTAIL.n253 B 0.024638f
C471 VTAIL.n254 B 0.024638f
C472 VTAIL.n255 B 0.013239f
C473 VTAIL.n256 B 0.014018f
C474 VTAIL.n257 B 0.031293f
C475 VTAIL.n258 B 0.031293f
C476 VTAIL.n259 B 0.014018f
C477 VTAIL.n260 B 0.013239f
C478 VTAIL.n261 B 0.024638f
C479 VTAIL.n262 B 0.024638f
C480 VTAIL.n263 B 0.013239f
C481 VTAIL.n264 B 0.014018f
C482 VTAIL.n265 B 0.031293f
C483 VTAIL.n266 B 0.069508f
C484 VTAIL.n267 B 0.014018f
C485 VTAIL.n268 B 0.013239f
C486 VTAIL.n269 B 0.058969f
C487 VTAIL.n270 B 0.039135f
C488 VTAIL.n271 B 1.70083f
C489 VDD1.n0 B 0.031391f
C490 VDD1.n1 B 0.021708f
C491 VDD1.n2 B 0.011665f
C492 VDD1.n3 B 0.027572f
C493 VDD1.n4 B 0.012351f
C494 VDD1.n5 B 0.021708f
C495 VDD1.n6 B 0.011665f
C496 VDD1.n7 B 0.027572f
C497 VDD1.n8 B 0.012351f
C498 VDD1.n9 B 0.021708f
C499 VDD1.n10 B 0.012008f
C500 VDD1.n11 B 0.027572f
C501 VDD1.n12 B 0.011665f
C502 VDD1.n13 B 0.012351f
C503 VDD1.n14 B 0.021708f
C504 VDD1.n15 B 0.011665f
C505 VDD1.n16 B 0.027572f
C506 VDD1.n17 B 0.012351f
C507 VDD1.n18 B 0.021708f
C508 VDD1.n19 B 0.011665f
C509 VDD1.n20 B 0.020679f
C510 VDD1.n21 B 0.019491f
C511 VDD1.t4 B 0.046588f
C512 VDD1.n22 B 0.158012f
C513 VDD1.n23 B 1.11251f
C514 VDD1.n24 B 0.011665f
C515 VDD1.n25 B 0.012351f
C516 VDD1.n26 B 0.027572f
C517 VDD1.n27 B 0.027572f
C518 VDD1.n28 B 0.012351f
C519 VDD1.n29 B 0.011665f
C520 VDD1.n30 B 0.021708f
C521 VDD1.n31 B 0.021708f
C522 VDD1.n32 B 0.011665f
C523 VDD1.n33 B 0.012351f
C524 VDD1.n34 B 0.027572f
C525 VDD1.n35 B 0.027572f
C526 VDD1.n36 B 0.012351f
C527 VDD1.n37 B 0.011665f
C528 VDD1.n38 B 0.021708f
C529 VDD1.n39 B 0.021708f
C530 VDD1.n40 B 0.011665f
C531 VDD1.n41 B 0.012351f
C532 VDD1.n42 B 0.027572f
C533 VDD1.n43 B 0.027572f
C534 VDD1.n44 B 0.027572f
C535 VDD1.n45 B 0.012008f
C536 VDD1.n46 B 0.011665f
C537 VDD1.n47 B 0.021708f
C538 VDD1.n48 B 0.021708f
C539 VDD1.n49 B 0.011665f
C540 VDD1.n50 B 0.012351f
C541 VDD1.n51 B 0.027572f
C542 VDD1.n52 B 0.027572f
C543 VDD1.n53 B 0.012351f
C544 VDD1.n54 B 0.011665f
C545 VDD1.n55 B 0.021708f
C546 VDD1.n56 B 0.021708f
C547 VDD1.n57 B 0.011665f
C548 VDD1.n58 B 0.012351f
C549 VDD1.n59 B 0.027572f
C550 VDD1.n60 B 0.061242f
C551 VDD1.n61 B 0.012351f
C552 VDD1.n62 B 0.011665f
C553 VDD1.n63 B 0.051956f
C554 VDD1.n64 B 0.062415f
C555 VDD1.n65 B 0.031391f
C556 VDD1.n66 B 0.021708f
C557 VDD1.n67 B 0.011665f
C558 VDD1.n68 B 0.027572f
C559 VDD1.n69 B 0.012351f
C560 VDD1.n70 B 0.021708f
C561 VDD1.n71 B 0.011665f
C562 VDD1.n72 B 0.027572f
C563 VDD1.n73 B 0.012351f
C564 VDD1.n74 B 0.021708f
C565 VDD1.n75 B 0.012008f
C566 VDD1.n76 B 0.027572f
C567 VDD1.n77 B 0.012351f
C568 VDD1.n78 B 0.021708f
C569 VDD1.n79 B 0.011665f
C570 VDD1.n80 B 0.027572f
C571 VDD1.n81 B 0.012351f
C572 VDD1.n82 B 0.021708f
C573 VDD1.n83 B 0.011665f
C574 VDD1.n84 B 0.020679f
C575 VDD1.n85 B 0.019491f
C576 VDD1.t2 B 0.046588f
C577 VDD1.n86 B 0.158012f
C578 VDD1.n87 B 1.11251f
C579 VDD1.n88 B 0.011665f
C580 VDD1.n89 B 0.012351f
C581 VDD1.n90 B 0.027572f
C582 VDD1.n91 B 0.027572f
C583 VDD1.n92 B 0.012351f
C584 VDD1.n93 B 0.011665f
C585 VDD1.n94 B 0.021708f
C586 VDD1.n95 B 0.021708f
C587 VDD1.n96 B 0.011665f
C588 VDD1.n97 B 0.012351f
C589 VDD1.n98 B 0.027572f
C590 VDD1.n99 B 0.027572f
C591 VDD1.n100 B 0.012351f
C592 VDD1.n101 B 0.011665f
C593 VDD1.n102 B 0.021708f
C594 VDD1.n103 B 0.021708f
C595 VDD1.n104 B 0.011665f
C596 VDD1.n105 B 0.011665f
C597 VDD1.n106 B 0.012351f
C598 VDD1.n107 B 0.027572f
C599 VDD1.n108 B 0.027572f
C600 VDD1.n109 B 0.027572f
C601 VDD1.n110 B 0.012008f
C602 VDD1.n111 B 0.011665f
C603 VDD1.n112 B 0.021708f
C604 VDD1.n113 B 0.021708f
C605 VDD1.n114 B 0.011665f
C606 VDD1.n115 B 0.012351f
C607 VDD1.n116 B 0.027572f
C608 VDD1.n117 B 0.027572f
C609 VDD1.n118 B 0.012351f
C610 VDD1.n119 B 0.011665f
C611 VDD1.n120 B 0.021708f
C612 VDD1.n121 B 0.021708f
C613 VDD1.n122 B 0.011665f
C614 VDD1.n123 B 0.012351f
C615 VDD1.n124 B 0.027572f
C616 VDD1.n125 B 0.061242f
C617 VDD1.n126 B 0.012351f
C618 VDD1.n127 B 0.011665f
C619 VDD1.n128 B 0.051956f
C620 VDD1.n129 B 0.061522f
C621 VDD1.t3 B 0.208939f
C622 VDD1.t5 B 0.208939f
C623 VDD1.n130 B 1.87126f
C624 VDD1.n131 B 2.98866f
C625 VDD1.t1 B 0.208939f
C626 VDD1.t0 B 0.208939f
C627 VDD1.n132 B 1.86432f
C628 VDD1.n133 B 2.76913f
C629 VP.t1 B 2.37558f
C630 VP.n0 B 0.900239f
C631 VP.n1 B 0.018024f
C632 VP.n2 B 0.035912f
C633 VP.n3 B 0.018024f
C634 VP.n4 B 0.033423f
C635 VP.n5 B 0.018024f
C636 VP.t0 B 2.37558f
C637 VP.n6 B 0.033423f
C638 VP.n7 B 0.018024f
C639 VP.n8 B 0.033423f
C640 VP.n9 B 0.029085f
C641 VP.t5 B 2.37558f
C642 VP.t4 B 2.37558f
C643 VP.n10 B 0.900239f
C644 VP.n11 B 0.018024f
C645 VP.n12 B 0.035912f
C646 VP.n13 B 0.018024f
C647 VP.n14 B 0.033423f
C648 VP.t3 B 2.67547f
C649 VP.n15 B 0.85126f
C650 VP.t2 B 2.37558f
C651 VP.n16 B 0.895954f
C652 VP.n17 B 0.025173f
C653 VP.n18 B 0.235514f
C654 VP.n19 B 0.018024f
C655 VP.n20 B 0.018024f
C656 VP.n21 B 0.033423f
C657 VP.n22 B 0.032918f
C658 VP.n23 B 0.016994f
C659 VP.n24 B 0.018024f
C660 VP.n25 B 0.018024f
C661 VP.n26 B 0.018024f
C662 VP.n27 B 0.033423f
C663 VP.n28 B 0.033423f
C664 VP.n29 B 0.018573f
C665 VP.n30 B 0.029085f
C666 VP.n31 B 1.16589f
C667 VP.n32 B 1.17787f
C668 VP.n33 B 0.900239f
C669 VP.n34 B 0.018573f
C670 VP.n35 B 0.033423f
C671 VP.n36 B 0.018024f
C672 VP.n37 B 0.018024f
C673 VP.n38 B 0.018024f
C674 VP.n39 B 0.035912f
C675 VP.n40 B 0.016994f
C676 VP.n41 B 0.032918f
C677 VP.n42 B 0.018024f
C678 VP.n43 B 0.018024f
C679 VP.n44 B 0.018024f
C680 VP.n45 B 0.033423f
C681 VP.n46 B 0.025173f
C682 VP.n47 B 0.830642f
C683 VP.n48 B 0.025173f
C684 VP.n49 B 0.018024f
C685 VP.n50 B 0.018024f
C686 VP.n51 B 0.018024f
C687 VP.n52 B 0.033423f
C688 VP.n53 B 0.032918f
C689 VP.n54 B 0.016994f
C690 VP.n55 B 0.018024f
C691 VP.n56 B 0.018024f
C692 VP.n57 B 0.018024f
C693 VP.n58 B 0.033423f
C694 VP.n59 B 0.033423f
C695 VP.n60 B 0.018573f
C696 VP.n61 B 0.029085f
C697 VP.n62 B 0.057238f
.ends

