* NGSPICE file created from diff_pair_sample_1549.ext - technology: sky130A

.subckt diff_pair_sample_1549 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=0 ps=0 w=5.94 l=2.56
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=2.3166 ps=12.66 w=5.94 l=2.56
X2 B.t8 B.t6 B.t7 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=0 ps=0 w=5.94 l=2.56
X3 B.t5 B.t3 B.t4 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=0 ps=0 w=5.94 l=2.56
X4 B.t2 B.t0 B.t1 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=0 ps=0 w=5.94 l=2.56
X5 VDD1.t1 VP.t0 VTAIL.t1 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=2.3166 ps=12.66 w=5.94 l=2.56
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=2.3166 ps=12.66 w=5.94 l=2.56
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n2126_n2156# sky130_fd_pr__pfet_01v8 ad=2.3166 pd=12.66 as=2.3166 ps=12.66 w=5.94 l=2.56
R0 B.n319 B.n318 585
R1 B.n320 B.n47 585
R2 B.n322 B.n321 585
R3 B.n323 B.n46 585
R4 B.n325 B.n324 585
R5 B.n326 B.n45 585
R6 B.n328 B.n327 585
R7 B.n329 B.n44 585
R8 B.n331 B.n330 585
R9 B.n332 B.n43 585
R10 B.n334 B.n333 585
R11 B.n335 B.n42 585
R12 B.n337 B.n336 585
R13 B.n338 B.n41 585
R14 B.n340 B.n339 585
R15 B.n341 B.n40 585
R16 B.n343 B.n342 585
R17 B.n344 B.n39 585
R18 B.n346 B.n345 585
R19 B.n347 B.n38 585
R20 B.n349 B.n348 585
R21 B.n350 B.n37 585
R22 B.n352 B.n351 585
R23 B.n353 B.n34 585
R24 B.n356 B.n355 585
R25 B.n357 B.n33 585
R26 B.n359 B.n358 585
R27 B.n360 B.n32 585
R28 B.n362 B.n361 585
R29 B.n363 B.n31 585
R30 B.n365 B.n364 585
R31 B.n366 B.n27 585
R32 B.n368 B.n367 585
R33 B.n369 B.n26 585
R34 B.n371 B.n370 585
R35 B.n372 B.n25 585
R36 B.n374 B.n373 585
R37 B.n375 B.n24 585
R38 B.n377 B.n376 585
R39 B.n378 B.n23 585
R40 B.n380 B.n379 585
R41 B.n381 B.n22 585
R42 B.n383 B.n382 585
R43 B.n384 B.n21 585
R44 B.n386 B.n385 585
R45 B.n387 B.n20 585
R46 B.n389 B.n388 585
R47 B.n390 B.n19 585
R48 B.n392 B.n391 585
R49 B.n393 B.n18 585
R50 B.n395 B.n394 585
R51 B.n396 B.n17 585
R52 B.n398 B.n397 585
R53 B.n399 B.n16 585
R54 B.n401 B.n400 585
R55 B.n402 B.n15 585
R56 B.n404 B.n403 585
R57 B.n317 B.n48 585
R58 B.n316 B.n315 585
R59 B.n314 B.n49 585
R60 B.n313 B.n312 585
R61 B.n311 B.n50 585
R62 B.n310 B.n309 585
R63 B.n308 B.n51 585
R64 B.n307 B.n306 585
R65 B.n305 B.n52 585
R66 B.n304 B.n303 585
R67 B.n302 B.n53 585
R68 B.n301 B.n300 585
R69 B.n299 B.n54 585
R70 B.n298 B.n297 585
R71 B.n296 B.n55 585
R72 B.n295 B.n294 585
R73 B.n293 B.n56 585
R74 B.n292 B.n291 585
R75 B.n290 B.n57 585
R76 B.n289 B.n288 585
R77 B.n287 B.n58 585
R78 B.n286 B.n285 585
R79 B.n284 B.n59 585
R80 B.n283 B.n282 585
R81 B.n281 B.n60 585
R82 B.n280 B.n279 585
R83 B.n278 B.n61 585
R84 B.n277 B.n276 585
R85 B.n275 B.n62 585
R86 B.n274 B.n273 585
R87 B.n272 B.n63 585
R88 B.n271 B.n270 585
R89 B.n269 B.n64 585
R90 B.n268 B.n267 585
R91 B.n266 B.n65 585
R92 B.n265 B.n264 585
R93 B.n263 B.n66 585
R94 B.n262 B.n261 585
R95 B.n260 B.n67 585
R96 B.n259 B.n258 585
R97 B.n257 B.n68 585
R98 B.n256 B.n255 585
R99 B.n254 B.n69 585
R100 B.n253 B.n252 585
R101 B.n251 B.n70 585
R102 B.n250 B.n249 585
R103 B.n248 B.n71 585
R104 B.n247 B.n246 585
R105 B.n245 B.n72 585
R106 B.n244 B.n243 585
R107 B.n242 B.n73 585
R108 B.n153 B.n152 585
R109 B.n154 B.n103 585
R110 B.n156 B.n155 585
R111 B.n157 B.n102 585
R112 B.n159 B.n158 585
R113 B.n160 B.n101 585
R114 B.n162 B.n161 585
R115 B.n163 B.n100 585
R116 B.n165 B.n164 585
R117 B.n166 B.n99 585
R118 B.n168 B.n167 585
R119 B.n169 B.n98 585
R120 B.n171 B.n170 585
R121 B.n172 B.n97 585
R122 B.n174 B.n173 585
R123 B.n175 B.n96 585
R124 B.n177 B.n176 585
R125 B.n178 B.n95 585
R126 B.n180 B.n179 585
R127 B.n181 B.n94 585
R128 B.n183 B.n182 585
R129 B.n184 B.n93 585
R130 B.n186 B.n185 585
R131 B.n187 B.n90 585
R132 B.n190 B.n189 585
R133 B.n191 B.n89 585
R134 B.n193 B.n192 585
R135 B.n194 B.n88 585
R136 B.n196 B.n195 585
R137 B.n197 B.n87 585
R138 B.n199 B.n198 585
R139 B.n200 B.n86 585
R140 B.n205 B.n204 585
R141 B.n206 B.n85 585
R142 B.n208 B.n207 585
R143 B.n209 B.n84 585
R144 B.n211 B.n210 585
R145 B.n212 B.n83 585
R146 B.n214 B.n213 585
R147 B.n215 B.n82 585
R148 B.n217 B.n216 585
R149 B.n218 B.n81 585
R150 B.n220 B.n219 585
R151 B.n221 B.n80 585
R152 B.n223 B.n222 585
R153 B.n224 B.n79 585
R154 B.n226 B.n225 585
R155 B.n227 B.n78 585
R156 B.n229 B.n228 585
R157 B.n230 B.n77 585
R158 B.n232 B.n231 585
R159 B.n233 B.n76 585
R160 B.n235 B.n234 585
R161 B.n236 B.n75 585
R162 B.n238 B.n237 585
R163 B.n239 B.n74 585
R164 B.n241 B.n240 585
R165 B.n151 B.n104 585
R166 B.n150 B.n149 585
R167 B.n148 B.n105 585
R168 B.n147 B.n146 585
R169 B.n145 B.n106 585
R170 B.n144 B.n143 585
R171 B.n142 B.n107 585
R172 B.n141 B.n140 585
R173 B.n139 B.n108 585
R174 B.n138 B.n137 585
R175 B.n136 B.n109 585
R176 B.n135 B.n134 585
R177 B.n133 B.n110 585
R178 B.n132 B.n131 585
R179 B.n130 B.n111 585
R180 B.n129 B.n128 585
R181 B.n127 B.n112 585
R182 B.n126 B.n125 585
R183 B.n124 B.n113 585
R184 B.n123 B.n122 585
R185 B.n121 B.n114 585
R186 B.n120 B.n119 585
R187 B.n118 B.n115 585
R188 B.n117 B.n116 585
R189 B.n2 B.n0 585
R190 B.n441 B.n1 585
R191 B.n440 B.n439 585
R192 B.n438 B.n3 585
R193 B.n437 B.n436 585
R194 B.n435 B.n4 585
R195 B.n434 B.n433 585
R196 B.n432 B.n5 585
R197 B.n431 B.n430 585
R198 B.n429 B.n6 585
R199 B.n428 B.n427 585
R200 B.n426 B.n7 585
R201 B.n425 B.n424 585
R202 B.n423 B.n8 585
R203 B.n422 B.n421 585
R204 B.n420 B.n9 585
R205 B.n419 B.n418 585
R206 B.n417 B.n10 585
R207 B.n416 B.n415 585
R208 B.n414 B.n11 585
R209 B.n413 B.n412 585
R210 B.n411 B.n12 585
R211 B.n410 B.n409 585
R212 B.n408 B.n13 585
R213 B.n407 B.n406 585
R214 B.n405 B.n14 585
R215 B.n443 B.n442 585
R216 B.n153 B.n104 530.939
R217 B.n405 B.n404 530.939
R218 B.n242 B.n241 530.939
R219 B.n319 B.n48 530.939
R220 B.n201 B.t5 323.077
R221 B.n35 B.t7 323.077
R222 B.n91 B.t11 323.077
R223 B.n28 B.t1 323.077
R224 B.n202 B.t4 267.029
R225 B.n36 B.t8 267.029
R226 B.n92 B.t10 267.029
R227 B.n29 B.t2 267.029
R228 B.n201 B.t3 263.906
R229 B.n91 B.t9 263.906
R230 B.n28 B.t0 263.906
R231 B.n35 B.t6 263.906
R232 B.n149 B.n104 163.367
R233 B.n149 B.n148 163.367
R234 B.n148 B.n147 163.367
R235 B.n147 B.n106 163.367
R236 B.n143 B.n106 163.367
R237 B.n143 B.n142 163.367
R238 B.n142 B.n141 163.367
R239 B.n141 B.n108 163.367
R240 B.n137 B.n108 163.367
R241 B.n137 B.n136 163.367
R242 B.n136 B.n135 163.367
R243 B.n135 B.n110 163.367
R244 B.n131 B.n110 163.367
R245 B.n131 B.n130 163.367
R246 B.n130 B.n129 163.367
R247 B.n129 B.n112 163.367
R248 B.n125 B.n112 163.367
R249 B.n125 B.n124 163.367
R250 B.n124 B.n123 163.367
R251 B.n123 B.n114 163.367
R252 B.n119 B.n114 163.367
R253 B.n119 B.n118 163.367
R254 B.n118 B.n117 163.367
R255 B.n117 B.n2 163.367
R256 B.n442 B.n2 163.367
R257 B.n442 B.n441 163.367
R258 B.n441 B.n440 163.367
R259 B.n440 B.n3 163.367
R260 B.n436 B.n3 163.367
R261 B.n436 B.n435 163.367
R262 B.n435 B.n434 163.367
R263 B.n434 B.n5 163.367
R264 B.n430 B.n5 163.367
R265 B.n430 B.n429 163.367
R266 B.n429 B.n428 163.367
R267 B.n428 B.n7 163.367
R268 B.n424 B.n7 163.367
R269 B.n424 B.n423 163.367
R270 B.n423 B.n422 163.367
R271 B.n422 B.n9 163.367
R272 B.n418 B.n9 163.367
R273 B.n418 B.n417 163.367
R274 B.n417 B.n416 163.367
R275 B.n416 B.n11 163.367
R276 B.n412 B.n11 163.367
R277 B.n412 B.n411 163.367
R278 B.n411 B.n410 163.367
R279 B.n410 B.n13 163.367
R280 B.n406 B.n13 163.367
R281 B.n406 B.n405 163.367
R282 B.n154 B.n153 163.367
R283 B.n155 B.n154 163.367
R284 B.n155 B.n102 163.367
R285 B.n159 B.n102 163.367
R286 B.n160 B.n159 163.367
R287 B.n161 B.n160 163.367
R288 B.n161 B.n100 163.367
R289 B.n165 B.n100 163.367
R290 B.n166 B.n165 163.367
R291 B.n167 B.n166 163.367
R292 B.n167 B.n98 163.367
R293 B.n171 B.n98 163.367
R294 B.n172 B.n171 163.367
R295 B.n173 B.n172 163.367
R296 B.n173 B.n96 163.367
R297 B.n177 B.n96 163.367
R298 B.n178 B.n177 163.367
R299 B.n179 B.n178 163.367
R300 B.n179 B.n94 163.367
R301 B.n183 B.n94 163.367
R302 B.n184 B.n183 163.367
R303 B.n185 B.n184 163.367
R304 B.n185 B.n90 163.367
R305 B.n190 B.n90 163.367
R306 B.n191 B.n190 163.367
R307 B.n192 B.n191 163.367
R308 B.n192 B.n88 163.367
R309 B.n196 B.n88 163.367
R310 B.n197 B.n196 163.367
R311 B.n198 B.n197 163.367
R312 B.n198 B.n86 163.367
R313 B.n205 B.n86 163.367
R314 B.n206 B.n205 163.367
R315 B.n207 B.n206 163.367
R316 B.n207 B.n84 163.367
R317 B.n211 B.n84 163.367
R318 B.n212 B.n211 163.367
R319 B.n213 B.n212 163.367
R320 B.n213 B.n82 163.367
R321 B.n217 B.n82 163.367
R322 B.n218 B.n217 163.367
R323 B.n219 B.n218 163.367
R324 B.n219 B.n80 163.367
R325 B.n223 B.n80 163.367
R326 B.n224 B.n223 163.367
R327 B.n225 B.n224 163.367
R328 B.n225 B.n78 163.367
R329 B.n229 B.n78 163.367
R330 B.n230 B.n229 163.367
R331 B.n231 B.n230 163.367
R332 B.n231 B.n76 163.367
R333 B.n235 B.n76 163.367
R334 B.n236 B.n235 163.367
R335 B.n237 B.n236 163.367
R336 B.n237 B.n74 163.367
R337 B.n241 B.n74 163.367
R338 B.n243 B.n242 163.367
R339 B.n243 B.n72 163.367
R340 B.n247 B.n72 163.367
R341 B.n248 B.n247 163.367
R342 B.n249 B.n248 163.367
R343 B.n249 B.n70 163.367
R344 B.n253 B.n70 163.367
R345 B.n254 B.n253 163.367
R346 B.n255 B.n254 163.367
R347 B.n255 B.n68 163.367
R348 B.n259 B.n68 163.367
R349 B.n260 B.n259 163.367
R350 B.n261 B.n260 163.367
R351 B.n261 B.n66 163.367
R352 B.n265 B.n66 163.367
R353 B.n266 B.n265 163.367
R354 B.n267 B.n266 163.367
R355 B.n267 B.n64 163.367
R356 B.n271 B.n64 163.367
R357 B.n272 B.n271 163.367
R358 B.n273 B.n272 163.367
R359 B.n273 B.n62 163.367
R360 B.n277 B.n62 163.367
R361 B.n278 B.n277 163.367
R362 B.n279 B.n278 163.367
R363 B.n279 B.n60 163.367
R364 B.n283 B.n60 163.367
R365 B.n284 B.n283 163.367
R366 B.n285 B.n284 163.367
R367 B.n285 B.n58 163.367
R368 B.n289 B.n58 163.367
R369 B.n290 B.n289 163.367
R370 B.n291 B.n290 163.367
R371 B.n291 B.n56 163.367
R372 B.n295 B.n56 163.367
R373 B.n296 B.n295 163.367
R374 B.n297 B.n296 163.367
R375 B.n297 B.n54 163.367
R376 B.n301 B.n54 163.367
R377 B.n302 B.n301 163.367
R378 B.n303 B.n302 163.367
R379 B.n303 B.n52 163.367
R380 B.n307 B.n52 163.367
R381 B.n308 B.n307 163.367
R382 B.n309 B.n308 163.367
R383 B.n309 B.n50 163.367
R384 B.n313 B.n50 163.367
R385 B.n314 B.n313 163.367
R386 B.n315 B.n314 163.367
R387 B.n315 B.n48 163.367
R388 B.n404 B.n15 163.367
R389 B.n400 B.n15 163.367
R390 B.n400 B.n399 163.367
R391 B.n399 B.n398 163.367
R392 B.n398 B.n17 163.367
R393 B.n394 B.n17 163.367
R394 B.n394 B.n393 163.367
R395 B.n393 B.n392 163.367
R396 B.n392 B.n19 163.367
R397 B.n388 B.n19 163.367
R398 B.n388 B.n387 163.367
R399 B.n387 B.n386 163.367
R400 B.n386 B.n21 163.367
R401 B.n382 B.n21 163.367
R402 B.n382 B.n381 163.367
R403 B.n381 B.n380 163.367
R404 B.n380 B.n23 163.367
R405 B.n376 B.n23 163.367
R406 B.n376 B.n375 163.367
R407 B.n375 B.n374 163.367
R408 B.n374 B.n25 163.367
R409 B.n370 B.n25 163.367
R410 B.n370 B.n369 163.367
R411 B.n369 B.n368 163.367
R412 B.n368 B.n27 163.367
R413 B.n364 B.n27 163.367
R414 B.n364 B.n363 163.367
R415 B.n363 B.n362 163.367
R416 B.n362 B.n32 163.367
R417 B.n358 B.n32 163.367
R418 B.n358 B.n357 163.367
R419 B.n357 B.n356 163.367
R420 B.n356 B.n34 163.367
R421 B.n351 B.n34 163.367
R422 B.n351 B.n350 163.367
R423 B.n350 B.n349 163.367
R424 B.n349 B.n38 163.367
R425 B.n345 B.n38 163.367
R426 B.n345 B.n344 163.367
R427 B.n344 B.n343 163.367
R428 B.n343 B.n40 163.367
R429 B.n339 B.n40 163.367
R430 B.n339 B.n338 163.367
R431 B.n338 B.n337 163.367
R432 B.n337 B.n42 163.367
R433 B.n333 B.n42 163.367
R434 B.n333 B.n332 163.367
R435 B.n332 B.n331 163.367
R436 B.n331 B.n44 163.367
R437 B.n327 B.n44 163.367
R438 B.n327 B.n326 163.367
R439 B.n326 B.n325 163.367
R440 B.n325 B.n46 163.367
R441 B.n321 B.n46 163.367
R442 B.n321 B.n320 163.367
R443 B.n320 B.n319 163.367
R444 B.n203 B.n202 59.5399
R445 B.n188 B.n92 59.5399
R446 B.n30 B.n29 59.5399
R447 B.n354 B.n36 59.5399
R448 B.n202 B.n201 56.049
R449 B.n92 B.n91 56.049
R450 B.n29 B.n28 56.049
R451 B.n36 B.n35 56.049
R452 B.n403 B.n14 34.4981
R453 B.n318 B.n317 34.4981
R454 B.n240 B.n73 34.4981
R455 B.n152 B.n151 34.4981
R456 B B.n443 18.0485
R457 B.n403 B.n402 10.6151
R458 B.n402 B.n401 10.6151
R459 B.n401 B.n16 10.6151
R460 B.n397 B.n16 10.6151
R461 B.n397 B.n396 10.6151
R462 B.n396 B.n395 10.6151
R463 B.n395 B.n18 10.6151
R464 B.n391 B.n18 10.6151
R465 B.n391 B.n390 10.6151
R466 B.n390 B.n389 10.6151
R467 B.n389 B.n20 10.6151
R468 B.n385 B.n20 10.6151
R469 B.n385 B.n384 10.6151
R470 B.n384 B.n383 10.6151
R471 B.n383 B.n22 10.6151
R472 B.n379 B.n22 10.6151
R473 B.n379 B.n378 10.6151
R474 B.n378 B.n377 10.6151
R475 B.n377 B.n24 10.6151
R476 B.n373 B.n24 10.6151
R477 B.n373 B.n372 10.6151
R478 B.n372 B.n371 10.6151
R479 B.n371 B.n26 10.6151
R480 B.n367 B.n366 10.6151
R481 B.n366 B.n365 10.6151
R482 B.n365 B.n31 10.6151
R483 B.n361 B.n31 10.6151
R484 B.n361 B.n360 10.6151
R485 B.n360 B.n359 10.6151
R486 B.n359 B.n33 10.6151
R487 B.n355 B.n33 10.6151
R488 B.n353 B.n352 10.6151
R489 B.n352 B.n37 10.6151
R490 B.n348 B.n37 10.6151
R491 B.n348 B.n347 10.6151
R492 B.n347 B.n346 10.6151
R493 B.n346 B.n39 10.6151
R494 B.n342 B.n39 10.6151
R495 B.n342 B.n341 10.6151
R496 B.n341 B.n340 10.6151
R497 B.n340 B.n41 10.6151
R498 B.n336 B.n41 10.6151
R499 B.n336 B.n335 10.6151
R500 B.n335 B.n334 10.6151
R501 B.n334 B.n43 10.6151
R502 B.n330 B.n43 10.6151
R503 B.n330 B.n329 10.6151
R504 B.n329 B.n328 10.6151
R505 B.n328 B.n45 10.6151
R506 B.n324 B.n45 10.6151
R507 B.n324 B.n323 10.6151
R508 B.n323 B.n322 10.6151
R509 B.n322 B.n47 10.6151
R510 B.n318 B.n47 10.6151
R511 B.n244 B.n73 10.6151
R512 B.n245 B.n244 10.6151
R513 B.n246 B.n245 10.6151
R514 B.n246 B.n71 10.6151
R515 B.n250 B.n71 10.6151
R516 B.n251 B.n250 10.6151
R517 B.n252 B.n251 10.6151
R518 B.n252 B.n69 10.6151
R519 B.n256 B.n69 10.6151
R520 B.n257 B.n256 10.6151
R521 B.n258 B.n257 10.6151
R522 B.n258 B.n67 10.6151
R523 B.n262 B.n67 10.6151
R524 B.n263 B.n262 10.6151
R525 B.n264 B.n263 10.6151
R526 B.n264 B.n65 10.6151
R527 B.n268 B.n65 10.6151
R528 B.n269 B.n268 10.6151
R529 B.n270 B.n269 10.6151
R530 B.n270 B.n63 10.6151
R531 B.n274 B.n63 10.6151
R532 B.n275 B.n274 10.6151
R533 B.n276 B.n275 10.6151
R534 B.n276 B.n61 10.6151
R535 B.n280 B.n61 10.6151
R536 B.n281 B.n280 10.6151
R537 B.n282 B.n281 10.6151
R538 B.n282 B.n59 10.6151
R539 B.n286 B.n59 10.6151
R540 B.n287 B.n286 10.6151
R541 B.n288 B.n287 10.6151
R542 B.n288 B.n57 10.6151
R543 B.n292 B.n57 10.6151
R544 B.n293 B.n292 10.6151
R545 B.n294 B.n293 10.6151
R546 B.n294 B.n55 10.6151
R547 B.n298 B.n55 10.6151
R548 B.n299 B.n298 10.6151
R549 B.n300 B.n299 10.6151
R550 B.n300 B.n53 10.6151
R551 B.n304 B.n53 10.6151
R552 B.n305 B.n304 10.6151
R553 B.n306 B.n305 10.6151
R554 B.n306 B.n51 10.6151
R555 B.n310 B.n51 10.6151
R556 B.n311 B.n310 10.6151
R557 B.n312 B.n311 10.6151
R558 B.n312 B.n49 10.6151
R559 B.n316 B.n49 10.6151
R560 B.n317 B.n316 10.6151
R561 B.n152 B.n103 10.6151
R562 B.n156 B.n103 10.6151
R563 B.n157 B.n156 10.6151
R564 B.n158 B.n157 10.6151
R565 B.n158 B.n101 10.6151
R566 B.n162 B.n101 10.6151
R567 B.n163 B.n162 10.6151
R568 B.n164 B.n163 10.6151
R569 B.n164 B.n99 10.6151
R570 B.n168 B.n99 10.6151
R571 B.n169 B.n168 10.6151
R572 B.n170 B.n169 10.6151
R573 B.n170 B.n97 10.6151
R574 B.n174 B.n97 10.6151
R575 B.n175 B.n174 10.6151
R576 B.n176 B.n175 10.6151
R577 B.n176 B.n95 10.6151
R578 B.n180 B.n95 10.6151
R579 B.n181 B.n180 10.6151
R580 B.n182 B.n181 10.6151
R581 B.n182 B.n93 10.6151
R582 B.n186 B.n93 10.6151
R583 B.n187 B.n186 10.6151
R584 B.n189 B.n89 10.6151
R585 B.n193 B.n89 10.6151
R586 B.n194 B.n193 10.6151
R587 B.n195 B.n194 10.6151
R588 B.n195 B.n87 10.6151
R589 B.n199 B.n87 10.6151
R590 B.n200 B.n199 10.6151
R591 B.n204 B.n200 10.6151
R592 B.n208 B.n85 10.6151
R593 B.n209 B.n208 10.6151
R594 B.n210 B.n209 10.6151
R595 B.n210 B.n83 10.6151
R596 B.n214 B.n83 10.6151
R597 B.n215 B.n214 10.6151
R598 B.n216 B.n215 10.6151
R599 B.n216 B.n81 10.6151
R600 B.n220 B.n81 10.6151
R601 B.n221 B.n220 10.6151
R602 B.n222 B.n221 10.6151
R603 B.n222 B.n79 10.6151
R604 B.n226 B.n79 10.6151
R605 B.n227 B.n226 10.6151
R606 B.n228 B.n227 10.6151
R607 B.n228 B.n77 10.6151
R608 B.n232 B.n77 10.6151
R609 B.n233 B.n232 10.6151
R610 B.n234 B.n233 10.6151
R611 B.n234 B.n75 10.6151
R612 B.n238 B.n75 10.6151
R613 B.n239 B.n238 10.6151
R614 B.n240 B.n239 10.6151
R615 B.n151 B.n150 10.6151
R616 B.n150 B.n105 10.6151
R617 B.n146 B.n105 10.6151
R618 B.n146 B.n145 10.6151
R619 B.n145 B.n144 10.6151
R620 B.n144 B.n107 10.6151
R621 B.n140 B.n107 10.6151
R622 B.n140 B.n139 10.6151
R623 B.n139 B.n138 10.6151
R624 B.n138 B.n109 10.6151
R625 B.n134 B.n109 10.6151
R626 B.n134 B.n133 10.6151
R627 B.n133 B.n132 10.6151
R628 B.n132 B.n111 10.6151
R629 B.n128 B.n111 10.6151
R630 B.n128 B.n127 10.6151
R631 B.n127 B.n126 10.6151
R632 B.n126 B.n113 10.6151
R633 B.n122 B.n113 10.6151
R634 B.n122 B.n121 10.6151
R635 B.n121 B.n120 10.6151
R636 B.n120 B.n115 10.6151
R637 B.n116 B.n115 10.6151
R638 B.n116 B.n0 10.6151
R639 B.n439 B.n1 10.6151
R640 B.n439 B.n438 10.6151
R641 B.n438 B.n437 10.6151
R642 B.n437 B.n4 10.6151
R643 B.n433 B.n4 10.6151
R644 B.n433 B.n432 10.6151
R645 B.n432 B.n431 10.6151
R646 B.n431 B.n6 10.6151
R647 B.n427 B.n6 10.6151
R648 B.n427 B.n426 10.6151
R649 B.n426 B.n425 10.6151
R650 B.n425 B.n8 10.6151
R651 B.n421 B.n8 10.6151
R652 B.n421 B.n420 10.6151
R653 B.n420 B.n419 10.6151
R654 B.n419 B.n10 10.6151
R655 B.n415 B.n10 10.6151
R656 B.n415 B.n414 10.6151
R657 B.n414 B.n413 10.6151
R658 B.n413 B.n12 10.6151
R659 B.n409 B.n12 10.6151
R660 B.n409 B.n408 10.6151
R661 B.n408 B.n407 10.6151
R662 B.n407 B.n14 10.6151
R663 B.n367 B.n30 6.5566
R664 B.n355 B.n354 6.5566
R665 B.n189 B.n188 6.5566
R666 B.n204 B.n203 6.5566
R667 B.n30 B.n26 4.05904
R668 B.n354 B.n353 4.05904
R669 B.n188 B.n187 4.05904
R670 B.n203 B.n85 4.05904
R671 B.n443 B.n0 2.81026
R672 B.n443 B.n1 2.81026
R673 VN VN.t0 145.191
R674 VN VN.t1 105.472
R675 VTAIL.n122 VTAIL.n96 756.745
R676 VTAIL.n26 VTAIL.n0 756.745
R677 VTAIL.n90 VTAIL.n64 756.745
R678 VTAIL.n58 VTAIL.n32 756.745
R679 VTAIL.n107 VTAIL.n106 585
R680 VTAIL.n104 VTAIL.n103 585
R681 VTAIL.n113 VTAIL.n112 585
R682 VTAIL.n115 VTAIL.n114 585
R683 VTAIL.n100 VTAIL.n99 585
R684 VTAIL.n121 VTAIL.n120 585
R685 VTAIL.n123 VTAIL.n122 585
R686 VTAIL.n11 VTAIL.n10 585
R687 VTAIL.n8 VTAIL.n7 585
R688 VTAIL.n17 VTAIL.n16 585
R689 VTAIL.n19 VTAIL.n18 585
R690 VTAIL.n4 VTAIL.n3 585
R691 VTAIL.n25 VTAIL.n24 585
R692 VTAIL.n27 VTAIL.n26 585
R693 VTAIL.n91 VTAIL.n90 585
R694 VTAIL.n89 VTAIL.n88 585
R695 VTAIL.n68 VTAIL.n67 585
R696 VTAIL.n83 VTAIL.n82 585
R697 VTAIL.n81 VTAIL.n80 585
R698 VTAIL.n72 VTAIL.n71 585
R699 VTAIL.n75 VTAIL.n74 585
R700 VTAIL.n59 VTAIL.n58 585
R701 VTAIL.n57 VTAIL.n56 585
R702 VTAIL.n36 VTAIL.n35 585
R703 VTAIL.n51 VTAIL.n50 585
R704 VTAIL.n49 VTAIL.n48 585
R705 VTAIL.n40 VTAIL.n39 585
R706 VTAIL.n43 VTAIL.n42 585
R707 VTAIL.t2 VTAIL.n105 327.601
R708 VTAIL.t0 VTAIL.n9 327.601
R709 VTAIL.t1 VTAIL.n73 327.601
R710 VTAIL.t3 VTAIL.n41 327.601
R711 VTAIL.n106 VTAIL.n103 171.744
R712 VTAIL.n113 VTAIL.n103 171.744
R713 VTAIL.n114 VTAIL.n113 171.744
R714 VTAIL.n114 VTAIL.n99 171.744
R715 VTAIL.n121 VTAIL.n99 171.744
R716 VTAIL.n122 VTAIL.n121 171.744
R717 VTAIL.n10 VTAIL.n7 171.744
R718 VTAIL.n17 VTAIL.n7 171.744
R719 VTAIL.n18 VTAIL.n17 171.744
R720 VTAIL.n18 VTAIL.n3 171.744
R721 VTAIL.n25 VTAIL.n3 171.744
R722 VTAIL.n26 VTAIL.n25 171.744
R723 VTAIL.n90 VTAIL.n89 171.744
R724 VTAIL.n89 VTAIL.n67 171.744
R725 VTAIL.n82 VTAIL.n67 171.744
R726 VTAIL.n82 VTAIL.n81 171.744
R727 VTAIL.n81 VTAIL.n71 171.744
R728 VTAIL.n74 VTAIL.n71 171.744
R729 VTAIL.n58 VTAIL.n57 171.744
R730 VTAIL.n57 VTAIL.n35 171.744
R731 VTAIL.n50 VTAIL.n35 171.744
R732 VTAIL.n50 VTAIL.n49 171.744
R733 VTAIL.n49 VTAIL.n39 171.744
R734 VTAIL.n42 VTAIL.n39 171.744
R735 VTAIL.n106 VTAIL.t2 85.8723
R736 VTAIL.n10 VTAIL.t0 85.8723
R737 VTAIL.n74 VTAIL.t1 85.8723
R738 VTAIL.n42 VTAIL.t3 85.8723
R739 VTAIL.n127 VTAIL.n126 31.0217
R740 VTAIL.n31 VTAIL.n30 31.0217
R741 VTAIL.n95 VTAIL.n94 31.0217
R742 VTAIL.n63 VTAIL.n62 31.0217
R743 VTAIL.n63 VTAIL.n31 22.4703
R744 VTAIL.n127 VTAIL.n95 19.9789
R745 VTAIL.n107 VTAIL.n105 16.3865
R746 VTAIL.n11 VTAIL.n9 16.3865
R747 VTAIL.n75 VTAIL.n73 16.3865
R748 VTAIL.n43 VTAIL.n41 16.3865
R749 VTAIL.n108 VTAIL.n104 12.8005
R750 VTAIL.n12 VTAIL.n8 12.8005
R751 VTAIL.n76 VTAIL.n72 12.8005
R752 VTAIL.n44 VTAIL.n40 12.8005
R753 VTAIL.n112 VTAIL.n111 12.0247
R754 VTAIL.n16 VTAIL.n15 12.0247
R755 VTAIL.n80 VTAIL.n79 12.0247
R756 VTAIL.n48 VTAIL.n47 12.0247
R757 VTAIL.n115 VTAIL.n102 11.249
R758 VTAIL.n19 VTAIL.n6 11.249
R759 VTAIL.n83 VTAIL.n70 11.249
R760 VTAIL.n51 VTAIL.n38 11.249
R761 VTAIL.n116 VTAIL.n100 10.4732
R762 VTAIL.n20 VTAIL.n4 10.4732
R763 VTAIL.n84 VTAIL.n68 10.4732
R764 VTAIL.n52 VTAIL.n36 10.4732
R765 VTAIL.n120 VTAIL.n119 9.69747
R766 VTAIL.n24 VTAIL.n23 9.69747
R767 VTAIL.n88 VTAIL.n87 9.69747
R768 VTAIL.n56 VTAIL.n55 9.69747
R769 VTAIL.n126 VTAIL.n125 9.45567
R770 VTAIL.n30 VTAIL.n29 9.45567
R771 VTAIL.n94 VTAIL.n93 9.45567
R772 VTAIL.n62 VTAIL.n61 9.45567
R773 VTAIL.n125 VTAIL.n124 9.3005
R774 VTAIL.n98 VTAIL.n97 9.3005
R775 VTAIL.n119 VTAIL.n118 9.3005
R776 VTAIL.n117 VTAIL.n116 9.3005
R777 VTAIL.n102 VTAIL.n101 9.3005
R778 VTAIL.n111 VTAIL.n110 9.3005
R779 VTAIL.n109 VTAIL.n108 9.3005
R780 VTAIL.n29 VTAIL.n28 9.3005
R781 VTAIL.n2 VTAIL.n1 9.3005
R782 VTAIL.n23 VTAIL.n22 9.3005
R783 VTAIL.n21 VTAIL.n20 9.3005
R784 VTAIL.n6 VTAIL.n5 9.3005
R785 VTAIL.n15 VTAIL.n14 9.3005
R786 VTAIL.n13 VTAIL.n12 9.3005
R787 VTAIL.n93 VTAIL.n92 9.3005
R788 VTAIL.n66 VTAIL.n65 9.3005
R789 VTAIL.n87 VTAIL.n86 9.3005
R790 VTAIL.n85 VTAIL.n84 9.3005
R791 VTAIL.n70 VTAIL.n69 9.3005
R792 VTAIL.n79 VTAIL.n78 9.3005
R793 VTAIL.n77 VTAIL.n76 9.3005
R794 VTAIL.n61 VTAIL.n60 9.3005
R795 VTAIL.n34 VTAIL.n33 9.3005
R796 VTAIL.n55 VTAIL.n54 9.3005
R797 VTAIL.n53 VTAIL.n52 9.3005
R798 VTAIL.n38 VTAIL.n37 9.3005
R799 VTAIL.n47 VTAIL.n46 9.3005
R800 VTAIL.n45 VTAIL.n44 9.3005
R801 VTAIL.n123 VTAIL.n98 8.92171
R802 VTAIL.n27 VTAIL.n2 8.92171
R803 VTAIL.n91 VTAIL.n66 8.92171
R804 VTAIL.n59 VTAIL.n34 8.92171
R805 VTAIL.n124 VTAIL.n96 8.14595
R806 VTAIL.n28 VTAIL.n0 8.14595
R807 VTAIL.n92 VTAIL.n64 8.14595
R808 VTAIL.n60 VTAIL.n32 8.14595
R809 VTAIL.n126 VTAIL.n96 5.81868
R810 VTAIL.n30 VTAIL.n0 5.81868
R811 VTAIL.n94 VTAIL.n64 5.81868
R812 VTAIL.n62 VTAIL.n32 5.81868
R813 VTAIL.n124 VTAIL.n123 5.04292
R814 VTAIL.n28 VTAIL.n27 5.04292
R815 VTAIL.n92 VTAIL.n91 5.04292
R816 VTAIL.n60 VTAIL.n59 5.04292
R817 VTAIL.n120 VTAIL.n98 4.26717
R818 VTAIL.n24 VTAIL.n2 4.26717
R819 VTAIL.n88 VTAIL.n66 4.26717
R820 VTAIL.n56 VTAIL.n34 4.26717
R821 VTAIL.n77 VTAIL.n73 3.71286
R822 VTAIL.n45 VTAIL.n41 3.71286
R823 VTAIL.n109 VTAIL.n105 3.71286
R824 VTAIL.n13 VTAIL.n9 3.71286
R825 VTAIL.n119 VTAIL.n100 3.49141
R826 VTAIL.n23 VTAIL.n4 3.49141
R827 VTAIL.n87 VTAIL.n68 3.49141
R828 VTAIL.n55 VTAIL.n36 3.49141
R829 VTAIL.n116 VTAIL.n115 2.71565
R830 VTAIL.n20 VTAIL.n19 2.71565
R831 VTAIL.n84 VTAIL.n83 2.71565
R832 VTAIL.n52 VTAIL.n51 2.71565
R833 VTAIL.n112 VTAIL.n102 1.93989
R834 VTAIL.n16 VTAIL.n6 1.93989
R835 VTAIL.n80 VTAIL.n70 1.93989
R836 VTAIL.n48 VTAIL.n38 1.93989
R837 VTAIL.n95 VTAIL.n63 1.71602
R838 VTAIL.n111 VTAIL.n104 1.16414
R839 VTAIL.n15 VTAIL.n8 1.16414
R840 VTAIL.n79 VTAIL.n72 1.16414
R841 VTAIL.n47 VTAIL.n40 1.16414
R842 VTAIL VTAIL.n31 1.15136
R843 VTAIL VTAIL.n127 0.565155
R844 VTAIL.n108 VTAIL.n107 0.388379
R845 VTAIL.n12 VTAIL.n11 0.388379
R846 VTAIL.n76 VTAIL.n75 0.388379
R847 VTAIL.n44 VTAIL.n43 0.388379
R848 VTAIL.n110 VTAIL.n109 0.155672
R849 VTAIL.n110 VTAIL.n101 0.155672
R850 VTAIL.n117 VTAIL.n101 0.155672
R851 VTAIL.n118 VTAIL.n117 0.155672
R852 VTAIL.n118 VTAIL.n97 0.155672
R853 VTAIL.n125 VTAIL.n97 0.155672
R854 VTAIL.n14 VTAIL.n13 0.155672
R855 VTAIL.n14 VTAIL.n5 0.155672
R856 VTAIL.n21 VTAIL.n5 0.155672
R857 VTAIL.n22 VTAIL.n21 0.155672
R858 VTAIL.n22 VTAIL.n1 0.155672
R859 VTAIL.n29 VTAIL.n1 0.155672
R860 VTAIL.n93 VTAIL.n65 0.155672
R861 VTAIL.n86 VTAIL.n65 0.155672
R862 VTAIL.n86 VTAIL.n85 0.155672
R863 VTAIL.n85 VTAIL.n69 0.155672
R864 VTAIL.n78 VTAIL.n69 0.155672
R865 VTAIL.n78 VTAIL.n77 0.155672
R866 VTAIL.n61 VTAIL.n33 0.155672
R867 VTAIL.n54 VTAIL.n33 0.155672
R868 VTAIL.n54 VTAIL.n53 0.155672
R869 VTAIL.n53 VTAIL.n37 0.155672
R870 VTAIL.n46 VTAIL.n37 0.155672
R871 VTAIL.n46 VTAIL.n45 0.155672
R872 VDD2.n57 VDD2.n31 756.745
R873 VDD2.n26 VDD2.n0 756.745
R874 VDD2.n58 VDD2.n57 585
R875 VDD2.n56 VDD2.n55 585
R876 VDD2.n35 VDD2.n34 585
R877 VDD2.n50 VDD2.n49 585
R878 VDD2.n48 VDD2.n47 585
R879 VDD2.n39 VDD2.n38 585
R880 VDD2.n42 VDD2.n41 585
R881 VDD2.n11 VDD2.n10 585
R882 VDD2.n8 VDD2.n7 585
R883 VDD2.n17 VDD2.n16 585
R884 VDD2.n19 VDD2.n18 585
R885 VDD2.n4 VDD2.n3 585
R886 VDD2.n25 VDD2.n24 585
R887 VDD2.n27 VDD2.n26 585
R888 VDD2.t1 VDD2.n40 327.601
R889 VDD2.t0 VDD2.n9 327.601
R890 VDD2.n57 VDD2.n56 171.744
R891 VDD2.n56 VDD2.n34 171.744
R892 VDD2.n49 VDD2.n34 171.744
R893 VDD2.n49 VDD2.n48 171.744
R894 VDD2.n48 VDD2.n38 171.744
R895 VDD2.n41 VDD2.n38 171.744
R896 VDD2.n10 VDD2.n7 171.744
R897 VDD2.n17 VDD2.n7 171.744
R898 VDD2.n18 VDD2.n17 171.744
R899 VDD2.n18 VDD2.n3 171.744
R900 VDD2.n25 VDD2.n3 171.744
R901 VDD2.n26 VDD2.n25 171.744
R902 VDD2.n41 VDD2.t1 85.8723
R903 VDD2.n10 VDD2.t0 85.8723
R904 VDD2.n62 VDD2.n30 81.4634
R905 VDD2.n62 VDD2.n61 47.7005
R906 VDD2.n42 VDD2.n40 16.3865
R907 VDD2.n11 VDD2.n9 16.3865
R908 VDD2.n43 VDD2.n39 12.8005
R909 VDD2.n12 VDD2.n8 12.8005
R910 VDD2.n47 VDD2.n46 12.0247
R911 VDD2.n16 VDD2.n15 12.0247
R912 VDD2.n50 VDD2.n37 11.249
R913 VDD2.n19 VDD2.n6 11.249
R914 VDD2.n51 VDD2.n35 10.4732
R915 VDD2.n20 VDD2.n4 10.4732
R916 VDD2.n55 VDD2.n54 9.69747
R917 VDD2.n24 VDD2.n23 9.69747
R918 VDD2.n61 VDD2.n60 9.45567
R919 VDD2.n30 VDD2.n29 9.45567
R920 VDD2.n60 VDD2.n59 9.3005
R921 VDD2.n33 VDD2.n32 9.3005
R922 VDD2.n54 VDD2.n53 9.3005
R923 VDD2.n52 VDD2.n51 9.3005
R924 VDD2.n37 VDD2.n36 9.3005
R925 VDD2.n46 VDD2.n45 9.3005
R926 VDD2.n44 VDD2.n43 9.3005
R927 VDD2.n29 VDD2.n28 9.3005
R928 VDD2.n2 VDD2.n1 9.3005
R929 VDD2.n23 VDD2.n22 9.3005
R930 VDD2.n21 VDD2.n20 9.3005
R931 VDD2.n6 VDD2.n5 9.3005
R932 VDD2.n15 VDD2.n14 9.3005
R933 VDD2.n13 VDD2.n12 9.3005
R934 VDD2.n58 VDD2.n33 8.92171
R935 VDD2.n27 VDD2.n2 8.92171
R936 VDD2.n59 VDD2.n31 8.14595
R937 VDD2.n28 VDD2.n0 8.14595
R938 VDD2.n61 VDD2.n31 5.81868
R939 VDD2.n30 VDD2.n0 5.81868
R940 VDD2.n59 VDD2.n58 5.04292
R941 VDD2.n28 VDD2.n27 5.04292
R942 VDD2.n55 VDD2.n33 4.26717
R943 VDD2.n24 VDD2.n2 4.26717
R944 VDD2.n44 VDD2.n40 3.71286
R945 VDD2.n13 VDD2.n9 3.71286
R946 VDD2.n54 VDD2.n35 3.49141
R947 VDD2.n23 VDD2.n4 3.49141
R948 VDD2.n51 VDD2.n50 2.71565
R949 VDD2.n20 VDD2.n19 2.71565
R950 VDD2.n47 VDD2.n37 1.93989
R951 VDD2.n16 VDD2.n6 1.93989
R952 VDD2.n46 VDD2.n39 1.16414
R953 VDD2.n15 VDD2.n8 1.16414
R954 VDD2 VDD2.n62 0.681535
R955 VDD2.n43 VDD2.n42 0.388379
R956 VDD2.n12 VDD2.n11 0.388379
R957 VDD2.n60 VDD2.n32 0.155672
R958 VDD2.n53 VDD2.n32 0.155672
R959 VDD2.n53 VDD2.n52 0.155672
R960 VDD2.n52 VDD2.n36 0.155672
R961 VDD2.n45 VDD2.n36 0.155672
R962 VDD2.n45 VDD2.n44 0.155672
R963 VDD2.n14 VDD2.n13 0.155672
R964 VDD2.n14 VDD2.n5 0.155672
R965 VDD2.n21 VDD2.n5 0.155672
R966 VDD2.n22 VDD2.n21 0.155672
R967 VDD2.n22 VDD2.n1 0.155672
R968 VDD2.n29 VDD2.n1 0.155672
R969 VP.n0 VP.t0 145.095
R970 VP.n0 VP.t1 105.135
R971 VP VP.n0 0.336784
R972 VDD1.n26 VDD1.n0 756.745
R973 VDD1.n57 VDD1.n31 756.745
R974 VDD1.n27 VDD1.n26 585
R975 VDD1.n25 VDD1.n24 585
R976 VDD1.n4 VDD1.n3 585
R977 VDD1.n19 VDD1.n18 585
R978 VDD1.n17 VDD1.n16 585
R979 VDD1.n8 VDD1.n7 585
R980 VDD1.n11 VDD1.n10 585
R981 VDD1.n42 VDD1.n41 585
R982 VDD1.n39 VDD1.n38 585
R983 VDD1.n48 VDD1.n47 585
R984 VDD1.n50 VDD1.n49 585
R985 VDD1.n35 VDD1.n34 585
R986 VDD1.n56 VDD1.n55 585
R987 VDD1.n58 VDD1.n57 585
R988 VDD1.t1 VDD1.n9 327.601
R989 VDD1.t0 VDD1.n40 327.601
R990 VDD1.n26 VDD1.n25 171.744
R991 VDD1.n25 VDD1.n3 171.744
R992 VDD1.n18 VDD1.n3 171.744
R993 VDD1.n18 VDD1.n17 171.744
R994 VDD1.n17 VDD1.n7 171.744
R995 VDD1.n10 VDD1.n7 171.744
R996 VDD1.n41 VDD1.n38 171.744
R997 VDD1.n48 VDD1.n38 171.744
R998 VDD1.n49 VDD1.n48 171.744
R999 VDD1.n49 VDD1.n34 171.744
R1000 VDD1.n56 VDD1.n34 171.744
R1001 VDD1.n57 VDD1.n56 171.744
R1002 VDD1.n10 VDD1.t1 85.8723
R1003 VDD1.n41 VDD1.t0 85.8723
R1004 VDD1 VDD1.n61 82.6111
R1005 VDD1 VDD1.n30 48.3815
R1006 VDD1.n11 VDD1.n9 16.3865
R1007 VDD1.n42 VDD1.n40 16.3865
R1008 VDD1.n12 VDD1.n8 12.8005
R1009 VDD1.n43 VDD1.n39 12.8005
R1010 VDD1.n16 VDD1.n15 12.0247
R1011 VDD1.n47 VDD1.n46 12.0247
R1012 VDD1.n19 VDD1.n6 11.249
R1013 VDD1.n50 VDD1.n37 11.249
R1014 VDD1.n20 VDD1.n4 10.4732
R1015 VDD1.n51 VDD1.n35 10.4732
R1016 VDD1.n24 VDD1.n23 9.69747
R1017 VDD1.n55 VDD1.n54 9.69747
R1018 VDD1.n30 VDD1.n29 9.45567
R1019 VDD1.n61 VDD1.n60 9.45567
R1020 VDD1.n29 VDD1.n28 9.3005
R1021 VDD1.n2 VDD1.n1 9.3005
R1022 VDD1.n23 VDD1.n22 9.3005
R1023 VDD1.n21 VDD1.n20 9.3005
R1024 VDD1.n6 VDD1.n5 9.3005
R1025 VDD1.n15 VDD1.n14 9.3005
R1026 VDD1.n13 VDD1.n12 9.3005
R1027 VDD1.n60 VDD1.n59 9.3005
R1028 VDD1.n33 VDD1.n32 9.3005
R1029 VDD1.n54 VDD1.n53 9.3005
R1030 VDD1.n52 VDD1.n51 9.3005
R1031 VDD1.n37 VDD1.n36 9.3005
R1032 VDD1.n46 VDD1.n45 9.3005
R1033 VDD1.n44 VDD1.n43 9.3005
R1034 VDD1.n27 VDD1.n2 8.92171
R1035 VDD1.n58 VDD1.n33 8.92171
R1036 VDD1.n28 VDD1.n0 8.14595
R1037 VDD1.n59 VDD1.n31 8.14595
R1038 VDD1.n30 VDD1.n0 5.81868
R1039 VDD1.n61 VDD1.n31 5.81868
R1040 VDD1.n28 VDD1.n27 5.04292
R1041 VDD1.n59 VDD1.n58 5.04292
R1042 VDD1.n24 VDD1.n2 4.26717
R1043 VDD1.n55 VDD1.n33 4.26717
R1044 VDD1.n13 VDD1.n9 3.71286
R1045 VDD1.n44 VDD1.n40 3.71286
R1046 VDD1.n23 VDD1.n4 3.49141
R1047 VDD1.n54 VDD1.n35 3.49141
R1048 VDD1.n20 VDD1.n19 2.71565
R1049 VDD1.n51 VDD1.n50 2.71565
R1050 VDD1.n16 VDD1.n6 1.93989
R1051 VDD1.n47 VDD1.n37 1.93989
R1052 VDD1.n15 VDD1.n8 1.16414
R1053 VDD1.n46 VDD1.n39 1.16414
R1054 VDD1.n12 VDD1.n11 0.388379
R1055 VDD1.n43 VDD1.n42 0.388379
R1056 VDD1.n29 VDD1.n1 0.155672
R1057 VDD1.n22 VDD1.n1 0.155672
R1058 VDD1.n22 VDD1.n21 0.155672
R1059 VDD1.n21 VDD1.n5 0.155672
R1060 VDD1.n14 VDD1.n5 0.155672
R1061 VDD1.n14 VDD1.n13 0.155672
R1062 VDD1.n45 VDD1.n44 0.155672
R1063 VDD1.n45 VDD1.n36 0.155672
R1064 VDD1.n52 VDD1.n36 0.155672
R1065 VDD1.n53 VDD1.n52 0.155672
R1066 VDD1.n53 VDD1.n32 0.155672
R1067 VDD1.n60 VDD1.n32 0.155672
C0 VDD2 VDD1 0.66908f
C1 VTAIL VDD2 3.50747f
C2 B w_n2126_n2156# 7.0777f
C3 VN VDD2 1.50186f
C4 VP w_n2126_n2156# 3.08304f
C5 B VDD1 1.22181f
C6 B VTAIL 2.27687f
C7 VP VDD1 1.68318f
C8 VP VTAIL 1.53668f
C9 VN B 0.970979f
C10 VN VP 4.30882f
C11 B VDD2 1.25153f
C12 VP VDD2 0.331232f
C13 VP B 1.4159f
C14 VDD1 w_n2126_n2156# 1.3549f
C15 VTAIL w_n2126_n2156# 1.89558f
C16 VTAIL VDD1 3.45574f
C17 VN w_n2126_n2156# 2.81231f
C18 VN VDD1 0.148438f
C19 VN VTAIL 1.52248f
C20 VDD2 w_n2126_n2156# 1.38029f
C21 VDD2 VSUBS 0.656363f
C22 VDD1 VSUBS 2.325111f
C23 VTAIL VSUBS 0.531008f
C24 VN VSUBS 5.2849f
C25 VP VSUBS 1.33842f
C26 B VSUBS 3.36886f
C27 w_n2126_n2156# VSUBS 57.223396f
C28 VDD1.n0 VSUBS 0.015456f
C29 VDD1.n1 VSUBS 0.014456f
C30 VDD1.n2 VSUBS 0.007768f
C31 VDD1.n3 VSUBS 0.018361f
C32 VDD1.n4 VSUBS 0.008225f
C33 VDD1.n5 VSUBS 0.014456f
C34 VDD1.n6 VSUBS 0.007768f
C35 VDD1.n7 VSUBS 0.018361f
C36 VDD1.n8 VSUBS 0.008225f
C37 VDD1.n9 VSUBS 0.063616f
C38 VDD1.t1 VSUBS 0.03935f
C39 VDD1.n10 VSUBS 0.013771f
C40 VDD1.n11 VSUBS 0.011674f
C41 VDD1.n12 VSUBS 0.007768f
C42 VDD1.n13 VSUBS 0.327776f
C43 VDD1.n14 VSUBS 0.014456f
C44 VDD1.n15 VSUBS 0.007768f
C45 VDD1.n16 VSUBS 0.008225f
C46 VDD1.n17 VSUBS 0.018361f
C47 VDD1.n18 VSUBS 0.018361f
C48 VDD1.n19 VSUBS 0.008225f
C49 VDD1.n20 VSUBS 0.007768f
C50 VDD1.n21 VSUBS 0.014456f
C51 VDD1.n22 VSUBS 0.014456f
C52 VDD1.n23 VSUBS 0.007768f
C53 VDD1.n24 VSUBS 0.008225f
C54 VDD1.n25 VSUBS 0.018361f
C55 VDD1.n26 VSUBS 0.042992f
C56 VDD1.n27 VSUBS 0.008225f
C57 VDD1.n28 VSUBS 0.007768f
C58 VDD1.n29 VSUBS 0.03223f
C59 VDD1.n30 VSUBS 0.032339f
C60 VDD1.n31 VSUBS 0.015456f
C61 VDD1.n32 VSUBS 0.014456f
C62 VDD1.n33 VSUBS 0.007768f
C63 VDD1.n34 VSUBS 0.018361f
C64 VDD1.n35 VSUBS 0.008225f
C65 VDD1.n36 VSUBS 0.014456f
C66 VDD1.n37 VSUBS 0.007768f
C67 VDD1.n38 VSUBS 0.018361f
C68 VDD1.n39 VSUBS 0.008225f
C69 VDD1.n40 VSUBS 0.063616f
C70 VDD1.t0 VSUBS 0.03935f
C71 VDD1.n41 VSUBS 0.013771f
C72 VDD1.n42 VSUBS 0.011674f
C73 VDD1.n43 VSUBS 0.007768f
C74 VDD1.n44 VSUBS 0.327776f
C75 VDD1.n45 VSUBS 0.014456f
C76 VDD1.n46 VSUBS 0.007768f
C77 VDD1.n47 VSUBS 0.008225f
C78 VDD1.n48 VSUBS 0.018361f
C79 VDD1.n49 VSUBS 0.018361f
C80 VDD1.n50 VSUBS 0.008225f
C81 VDD1.n51 VSUBS 0.007768f
C82 VDD1.n52 VSUBS 0.014456f
C83 VDD1.n53 VSUBS 0.014456f
C84 VDD1.n54 VSUBS 0.007768f
C85 VDD1.n55 VSUBS 0.008225f
C86 VDD1.n56 VSUBS 0.018361f
C87 VDD1.n57 VSUBS 0.042992f
C88 VDD1.n58 VSUBS 0.008225f
C89 VDD1.n59 VSUBS 0.007768f
C90 VDD1.n60 VSUBS 0.03223f
C91 VDD1.n61 VSUBS 0.33511f
C92 VP.t0 VSUBS 2.3076f
C93 VP.t1 VSUBS 1.78442f
C94 VP.n0 VSUBS 3.22457f
C95 VDD2.n0 VSUBS 0.015696f
C96 VDD2.n1 VSUBS 0.01468f
C97 VDD2.n2 VSUBS 0.007889f
C98 VDD2.n3 VSUBS 0.018646f
C99 VDD2.n4 VSUBS 0.008353f
C100 VDD2.n5 VSUBS 0.01468f
C101 VDD2.n6 VSUBS 0.007889f
C102 VDD2.n7 VSUBS 0.018646f
C103 VDD2.n8 VSUBS 0.008353f
C104 VDD2.n9 VSUBS 0.064602f
C105 VDD2.t0 VSUBS 0.039959f
C106 VDD2.n10 VSUBS 0.013984f
C107 VDD2.n11 VSUBS 0.011855f
C108 VDD2.n12 VSUBS 0.007889f
C109 VDD2.n13 VSUBS 0.332854f
C110 VDD2.n14 VSUBS 0.01468f
C111 VDD2.n15 VSUBS 0.007889f
C112 VDD2.n16 VSUBS 0.008353f
C113 VDD2.n17 VSUBS 0.018646f
C114 VDD2.n18 VSUBS 0.018646f
C115 VDD2.n19 VSUBS 0.008353f
C116 VDD2.n20 VSUBS 0.007889f
C117 VDD2.n21 VSUBS 0.01468f
C118 VDD2.n22 VSUBS 0.01468f
C119 VDD2.n23 VSUBS 0.007889f
C120 VDD2.n24 VSUBS 0.008353f
C121 VDD2.n25 VSUBS 0.018646f
C122 VDD2.n26 VSUBS 0.043658f
C123 VDD2.n27 VSUBS 0.008353f
C124 VDD2.n28 VSUBS 0.007889f
C125 VDD2.n29 VSUBS 0.03273f
C126 VDD2.n30 VSUBS 0.314712f
C127 VDD2.n31 VSUBS 0.015696f
C128 VDD2.n32 VSUBS 0.01468f
C129 VDD2.n33 VSUBS 0.007889f
C130 VDD2.n34 VSUBS 0.018646f
C131 VDD2.n35 VSUBS 0.008353f
C132 VDD2.n36 VSUBS 0.01468f
C133 VDD2.n37 VSUBS 0.007889f
C134 VDD2.n38 VSUBS 0.018646f
C135 VDD2.n39 VSUBS 0.008353f
C136 VDD2.n40 VSUBS 0.064602f
C137 VDD2.t1 VSUBS 0.039959f
C138 VDD2.n41 VSUBS 0.013984f
C139 VDD2.n42 VSUBS 0.011855f
C140 VDD2.n43 VSUBS 0.007889f
C141 VDD2.n44 VSUBS 0.332854f
C142 VDD2.n45 VSUBS 0.01468f
C143 VDD2.n46 VSUBS 0.007889f
C144 VDD2.n47 VSUBS 0.008353f
C145 VDD2.n48 VSUBS 0.018646f
C146 VDD2.n49 VSUBS 0.018646f
C147 VDD2.n50 VSUBS 0.008353f
C148 VDD2.n51 VSUBS 0.007889f
C149 VDD2.n52 VSUBS 0.01468f
C150 VDD2.n53 VSUBS 0.01468f
C151 VDD2.n54 VSUBS 0.007889f
C152 VDD2.n55 VSUBS 0.008353f
C153 VDD2.n56 VSUBS 0.018646f
C154 VDD2.n57 VSUBS 0.043658f
C155 VDD2.n58 VSUBS 0.008353f
C156 VDD2.n59 VSUBS 0.007889f
C157 VDD2.n60 VSUBS 0.03273f
C158 VDD2.n61 VSUBS 0.031999f
C159 VDD2.n62 VSUBS 1.40713f
C160 VTAIL.n0 VSUBS 0.023384f
C161 VTAIL.n1 VSUBS 0.021871f
C162 VTAIL.n2 VSUBS 0.011753f
C163 VTAIL.n3 VSUBS 0.027779f
C164 VTAIL.n4 VSUBS 0.012444f
C165 VTAIL.n5 VSUBS 0.021871f
C166 VTAIL.n6 VSUBS 0.011753f
C167 VTAIL.n7 VSUBS 0.027779f
C168 VTAIL.n8 VSUBS 0.012444f
C169 VTAIL.n9 VSUBS 0.096245f
C170 VTAIL.t0 VSUBS 0.059533f
C171 VTAIL.n10 VSUBS 0.020834f
C172 VTAIL.n11 VSUBS 0.017662f
C173 VTAIL.n12 VSUBS 0.011753f
C174 VTAIL.n13 VSUBS 0.495894f
C175 VTAIL.n14 VSUBS 0.021871f
C176 VTAIL.n15 VSUBS 0.011753f
C177 VTAIL.n16 VSUBS 0.012444f
C178 VTAIL.n17 VSUBS 0.027779f
C179 VTAIL.n18 VSUBS 0.027779f
C180 VTAIL.n19 VSUBS 0.012444f
C181 VTAIL.n20 VSUBS 0.011753f
C182 VTAIL.n21 VSUBS 0.021871f
C183 VTAIL.n22 VSUBS 0.021871f
C184 VTAIL.n23 VSUBS 0.011753f
C185 VTAIL.n24 VSUBS 0.012444f
C186 VTAIL.n25 VSUBS 0.027779f
C187 VTAIL.n26 VSUBS 0.065044f
C188 VTAIL.n27 VSUBS 0.012444f
C189 VTAIL.n28 VSUBS 0.011753f
C190 VTAIL.n29 VSUBS 0.048761f
C191 VTAIL.n30 VSUBS 0.032556f
C192 VTAIL.n31 VSUBS 1.1079f
C193 VTAIL.n32 VSUBS 0.023384f
C194 VTAIL.n33 VSUBS 0.021871f
C195 VTAIL.n34 VSUBS 0.011753f
C196 VTAIL.n35 VSUBS 0.027779f
C197 VTAIL.n36 VSUBS 0.012444f
C198 VTAIL.n37 VSUBS 0.021871f
C199 VTAIL.n38 VSUBS 0.011753f
C200 VTAIL.n39 VSUBS 0.027779f
C201 VTAIL.n40 VSUBS 0.012444f
C202 VTAIL.n41 VSUBS 0.096245f
C203 VTAIL.t3 VSUBS 0.059533f
C204 VTAIL.n42 VSUBS 0.020834f
C205 VTAIL.n43 VSUBS 0.017662f
C206 VTAIL.n44 VSUBS 0.011753f
C207 VTAIL.n45 VSUBS 0.495894f
C208 VTAIL.n46 VSUBS 0.021871f
C209 VTAIL.n47 VSUBS 0.011753f
C210 VTAIL.n48 VSUBS 0.012444f
C211 VTAIL.n49 VSUBS 0.027779f
C212 VTAIL.n50 VSUBS 0.027779f
C213 VTAIL.n51 VSUBS 0.012444f
C214 VTAIL.n52 VSUBS 0.011753f
C215 VTAIL.n53 VSUBS 0.021871f
C216 VTAIL.n54 VSUBS 0.021871f
C217 VTAIL.n55 VSUBS 0.011753f
C218 VTAIL.n56 VSUBS 0.012444f
C219 VTAIL.n57 VSUBS 0.027779f
C220 VTAIL.n58 VSUBS 0.065044f
C221 VTAIL.n59 VSUBS 0.012444f
C222 VTAIL.n60 VSUBS 0.011753f
C223 VTAIL.n61 VSUBS 0.048761f
C224 VTAIL.n62 VSUBS 0.032556f
C225 VTAIL.n63 VSUBS 1.14769f
C226 VTAIL.n64 VSUBS 0.023384f
C227 VTAIL.n65 VSUBS 0.021871f
C228 VTAIL.n66 VSUBS 0.011753f
C229 VTAIL.n67 VSUBS 0.027779f
C230 VTAIL.n68 VSUBS 0.012444f
C231 VTAIL.n69 VSUBS 0.021871f
C232 VTAIL.n70 VSUBS 0.011753f
C233 VTAIL.n71 VSUBS 0.027779f
C234 VTAIL.n72 VSUBS 0.012444f
C235 VTAIL.n73 VSUBS 0.096245f
C236 VTAIL.t1 VSUBS 0.059533f
C237 VTAIL.n74 VSUBS 0.020834f
C238 VTAIL.n75 VSUBS 0.017662f
C239 VTAIL.n76 VSUBS 0.011753f
C240 VTAIL.n77 VSUBS 0.495894f
C241 VTAIL.n78 VSUBS 0.021871f
C242 VTAIL.n79 VSUBS 0.011753f
C243 VTAIL.n80 VSUBS 0.012444f
C244 VTAIL.n81 VSUBS 0.027779f
C245 VTAIL.n82 VSUBS 0.027779f
C246 VTAIL.n83 VSUBS 0.012444f
C247 VTAIL.n84 VSUBS 0.011753f
C248 VTAIL.n85 VSUBS 0.021871f
C249 VTAIL.n86 VSUBS 0.021871f
C250 VTAIL.n87 VSUBS 0.011753f
C251 VTAIL.n88 VSUBS 0.012444f
C252 VTAIL.n89 VSUBS 0.027779f
C253 VTAIL.n90 VSUBS 0.065044f
C254 VTAIL.n91 VSUBS 0.012444f
C255 VTAIL.n92 VSUBS 0.011753f
C256 VTAIL.n93 VSUBS 0.048761f
C257 VTAIL.n94 VSUBS 0.032556f
C258 VTAIL.n95 VSUBS 0.972114f
C259 VTAIL.n96 VSUBS 0.023384f
C260 VTAIL.n97 VSUBS 0.021871f
C261 VTAIL.n98 VSUBS 0.011753f
C262 VTAIL.n99 VSUBS 0.027779f
C263 VTAIL.n100 VSUBS 0.012444f
C264 VTAIL.n101 VSUBS 0.021871f
C265 VTAIL.n102 VSUBS 0.011753f
C266 VTAIL.n103 VSUBS 0.027779f
C267 VTAIL.n104 VSUBS 0.012444f
C268 VTAIL.n105 VSUBS 0.096245f
C269 VTAIL.t2 VSUBS 0.059533f
C270 VTAIL.n106 VSUBS 0.020834f
C271 VTAIL.n107 VSUBS 0.017662f
C272 VTAIL.n108 VSUBS 0.011753f
C273 VTAIL.n109 VSUBS 0.495894f
C274 VTAIL.n110 VSUBS 0.021871f
C275 VTAIL.n111 VSUBS 0.011753f
C276 VTAIL.n112 VSUBS 0.012444f
C277 VTAIL.n113 VSUBS 0.027779f
C278 VTAIL.n114 VSUBS 0.027779f
C279 VTAIL.n115 VSUBS 0.012444f
C280 VTAIL.n116 VSUBS 0.011753f
C281 VTAIL.n117 VSUBS 0.021871f
C282 VTAIL.n118 VSUBS 0.021871f
C283 VTAIL.n119 VSUBS 0.011753f
C284 VTAIL.n120 VSUBS 0.012444f
C285 VTAIL.n121 VSUBS 0.027779f
C286 VTAIL.n122 VSUBS 0.065044f
C287 VTAIL.n123 VSUBS 0.012444f
C288 VTAIL.n124 VSUBS 0.011753f
C289 VTAIL.n125 VSUBS 0.048761f
C290 VTAIL.n126 VSUBS 0.032556f
C291 VTAIL.n127 VSUBS 0.891009f
C292 VN.t1 VSUBS 1.70235f
C293 VN.t0 VSUBS 2.20363f
C294 B.n0 VSUBS 0.004996f
C295 B.n1 VSUBS 0.004996f
C296 B.n2 VSUBS 0.007901f
C297 B.n3 VSUBS 0.007901f
C298 B.n4 VSUBS 0.007901f
C299 B.n5 VSUBS 0.007901f
C300 B.n6 VSUBS 0.007901f
C301 B.n7 VSUBS 0.007901f
C302 B.n8 VSUBS 0.007901f
C303 B.n9 VSUBS 0.007901f
C304 B.n10 VSUBS 0.007901f
C305 B.n11 VSUBS 0.007901f
C306 B.n12 VSUBS 0.007901f
C307 B.n13 VSUBS 0.007901f
C308 B.n14 VSUBS 0.01873f
C309 B.n15 VSUBS 0.007901f
C310 B.n16 VSUBS 0.007901f
C311 B.n17 VSUBS 0.007901f
C312 B.n18 VSUBS 0.007901f
C313 B.n19 VSUBS 0.007901f
C314 B.n20 VSUBS 0.007901f
C315 B.n21 VSUBS 0.007901f
C316 B.n22 VSUBS 0.007901f
C317 B.n23 VSUBS 0.007901f
C318 B.n24 VSUBS 0.007901f
C319 B.n25 VSUBS 0.007901f
C320 B.n26 VSUBS 0.005461f
C321 B.n27 VSUBS 0.007901f
C322 B.t2 VSUBS 0.099699f
C323 B.t1 VSUBS 0.128147f
C324 B.t0 VSUBS 0.811564f
C325 B.n28 VSUBS 0.21905f
C326 B.n29 VSUBS 0.17525f
C327 B.n30 VSUBS 0.018306f
C328 B.n31 VSUBS 0.007901f
C329 B.n32 VSUBS 0.007901f
C330 B.n33 VSUBS 0.007901f
C331 B.n34 VSUBS 0.007901f
C332 B.t8 VSUBS 0.099701f
C333 B.t7 VSUBS 0.128148f
C334 B.t6 VSUBS 0.811564f
C335 B.n35 VSUBS 0.219048f
C336 B.n36 VSUBS 0.175248f
C337 B.n37 VSUBS 0.007901f
C338 B.n38 VSUBS 0.007901f
C339 B.n39 VSUBS 0.007901f
C340 B.n40 VSUBS 0.007901f
C341 B.n41 VSUBS 0.007901f
C342 B.n42 VSUBS 0.007901f
C343 B.n43 VSUBS 0.007901f
C344 B.n44 VSUBS 0.007901f
C345 B.n45 VSUBS 0.007901f
C346 B.n46 VSUBS 0.007901f
C347 B.n47 VSUBS 0.007901f
C348 B.n48 VSUBS 0.01873f
C349 B.n49 VSUBS 0.007901f
C350 B.n50 VSUBS 0.007901f
C351 B.n51 VSUBS 0.007901f
C352 B.n52 VSUBS 0.007901f
C353 B.n53 VSUBS 0.007901f
C354 B.n54 VSUBS 0.007901f
C355 B.n55 VSUBS 0.007901f
C356 B.n56 VSUBS 0.007901f
C357 B.n57 VSUBS 0.007901f
C358 B.n58 VSUBS 0.007901f
C359 B.n59 VSUBS 0.007901f
C360 B.n60 VSUBS 0.007901f
C361 B.n61 VSUBS 0.007901f
C362 B.n62 VSUBS 0.007901f
C363 B.n63 VSUBS 0.007901f
C364 B.n64 VSUBS 0.007901f
C365 B.n65 VSUBS 0.007901f
C366 B.n66 VSUBS 0.007901f
C367 B.n67 VSUBS 0.007901f
C368 B.n68 VSUBS 0.007901f
C369 B.n69 VSUBS 0.007901f
C370 B.n70 VSUBS 0.007901f
C371 B.n71 VSUBS 0.007901f
C372 B.n72 VSUBS 0.007901f
C373 B.n73 VSUBS 0.01873f
C374 B.n74 VSUBS 0.007901f
C375 B.n75 VSUBS 0.007901f
C376 B.n76 VSUBS 0.007901f
C377 B.n77 VSUBS 0.007901f
C378 B.n78 VSUBS 0.007901f
C379 B.n79 VSUBS 0.007901f
C380 B.n80 VSUBS 0.007901f
C381 B.n81 VSUBS 0.007901f
C382 B.n82 VSUBS 0.007901f
C383 B.n83 VSUBS 0.007901f
C384 B.n84 VSUBS 0.007901f
C385 B.n85 VSUBS 0.005461f
C386 B.n86 VSUBS 0.007901f
C387 B.n87 VSUBS 0.007901f
C388 B.n88 VSUBS 0.007901f
C389 B.n89 VSUBS 0.007901f
C390 B.n90 VSUBS 0.007901f
C391 B.t10 VSUBS 0.099699f
C392 B.t11 VSUBS 0.128147f
C393 B.t9 VSUBS 0.811564f
C394 B.n91 VSUBS 0.21905f
C395 B.n92 VSUBS 0.17525f
C396 B.n93 VSUBS 0.007901f
C397 B.n94 VSUBS 0.007901f
C398 B.n95 VSUBS 0.007901f
C399 B.n96 VSUBS 0.007901f
C400 B.n97 VSUBS 0.007901f
C401 B.n98 VSUBS 0.007901f
C402 B.n99 VSUBS 0.007901f
C403 B.n100 VSUBS 0.007901f
C404 B.n101 VSUBS 0.007901f
C405 B.n102 VSUBS 0.007901f
C406 B.n103 VSUBS 0.007901f
C407 B.n104 VSUBS 0.01873f
C408 B.n105 VSUBS 0.007901f
C409 B.n106 VSUBS 0.007901f
C410 B.n107 VSUBS 0.007901f
C411 B.n108 VSUBS 0.007901f
C412 B.n109 VSUBS 0.007901f
C413 B.n110 VSUBS 0.007901f
C414 B.n111 VSUBS 0.007901f
C415 B.n112 VSUBS 0.007901f
C416 B.n113 VSUBS 0.007901f
C417 B.n114 VSUBS 0.007901f
C418 B.n115 VSUBS 0.007901f
C419 B.n116 VSUBS 0.007901f
C420 B.n117 VSUBS 0.007901f
C421 B.n118 VSUBS 0.007901f
C422 B.n119 VSUBS 0.007901f
C423 B.n120 VSUBS 0.007901f
C424 B.n121 VSUBS 0.007901f
C425 B.n122 VSUBS 0.007901f
C426 B.n123 VSUBS 0.007901f
C427 B.n124 VSUBS 0.007901f
C428 B.n125 VSUBS 0.007901f
C429 B.n126 VSUBS 0.007901f
C430 B.n127 VSUBS 0.007901f
C431 B.n128 VSUBS 0.007901f
C432 B.n129 VSUBS 0.007901f
C433 B.n130 VSUBS 0.007901f
C434 B.n131 VSUBS 0.007901f
C435 B.n132 VSUBS 0.007901f
C436 B.n133 VSUBS 0.007901f
C437 B.n134 VSUBS 0.007901f
C438 B.n135 VSUBS 0.007901f
C439 B.n136 VSUBS 0.007901f
C440 B.n137 VSUBS 0.007901f
C441 B.n138 VSUBS 0.007901f
C442 B.n139 VSUBS 0.007901f
C443 B.n140 VSUBS 0.007901f
C444 B.n141 VSUBS 0.007901f
C445 B.n142 VSUBS 0.007901f
C446 B.n143 VSUBS 0.007901f
C447 B.n144 VSUBS 0.007901f
C448 B.n145 VSUBS 0.007901f
C449 B.n146 VSUBS 0.007901f
C450 B.n147 VSUBS 0.007901f
C451 B.n148 VSUBS 0.007901f
C452 B.n149 VSUBS 0.007901f
C453 B.n150 VSUBS 0.007901f
C454 B.n151 VSUBS 0.01873f
C455 B.n152 VSUBS 0.019614f
C456 B.n153 VSUBS 0.019614f
C457 B.n154 VSUBS 0.007901f
C458 B.n155 VSUBS 0.007901f
C459 B.n156 VSUBS 0.007901f
C460 B.n157 VSUBS 0.007901f
C461 B.n158 VSUBS 0.007901f
C462 B.n159 VSUBS 0.007901f
C463 B.n160 VSUBS 0.007901f
C464 B.n161 VSUBS 0.007901f
C465 B.n162 VSUBS 0.007901f
C466 B.n163 VSUBS 0.007901f
C467 B.n164 VSUBS 0.007901f
C468 B.n165 VSUBS 0.007901f
C469 B.n166 VSUBS 0.007901f
C470 B.n167 VSUBS 0.007901f
C471 B.n168 VSUBS 0.007901f
C472 B.n169 VSUBS 0.007901f
C473 B.n170 VSUBS 0.007901f
C474 B.n171 VSUBS 0.007901f
C475 B.n172 VSUBS 0.007901f
C476 B.n173 VSUBS 0.007901f
C477 B.n174 VSUBS 0.007901f
C478 B.n175 VSUBS 0.007901f
C479 B.n176 VSUBS 0.007901f
C480 B.n177 VSUBS 0.007901f
C481 B.n178 VSUBS 0.007901f
C482 B.n179 VSUBS 0.007901f
C483 B.n180 VSUBS 0.007901f
C484 B.n181 VSUBS 0.007901f
C485 B.n182 VSUBS 0.007901f
C486 B.n183 VSUBS 0.007901f
C487 B.n184 VSUBS 0.007901f
C488 B.n185 VSUBS 0.007901f
C489 B.n186 VSUBS 0.007901f
C490 B.n187 VSUBS 0.005461f
C491 B.n188 VSUBS 0.018306f
C492 B.n189 VSUBS 0.006391f
C493 B.n190 VSUBS 0.007901f
C494 B.n191 VSUBS 0.007901f
C495 B.n192 VSUBS 0.007901f
C496 B.n193 VSUBS 0.007901f
C497 B.n194 VSUBS 0.007901f
C498 B.n195 VSUBS 0.007901f
C499 B.n196 VSUBS 0.007901f
C500 B.n197 VSUBS 0.007901f
C501 B.n198 VSUBS 0.007901f
C502 B.n199 VSUBS 0.007901f
C503 B.n200 VSUBS 0.007901f
C504 B.t4 VSUBS 0.099701f
C505 B.t5 VSUBS 0.128148f
C506 B.t3 VSUBS 0.811564f
C507 B.n201 VSUBS 0.219048f
C508 B.n202 VSUBS 0.175248f
C509 B.n203 VSUBS 0.018306f
C510 B.n204 VSUBS 0.006391f
C511 B.n205 VSUBS 0.007901f
C512 B.n206 VSUBS 0.007901f
C513 B.n207 VSUBS 0.007901f
C514 B.n208 VSUBS 0.007901f
C515 B.n209 VSUBS 0.007901f
C516 B.n210 VSUBS 0.007901f
C517 B.n211 VSUBS 0.007901f
C518 B.n212 VSUBS 0.007901f
C519 B.n213 VSUBS 0.007901f
C520 B.n214 VSUBS 0.007901f
C521 B.n215 VSUBS 0.007901f
C522 B.n216 VSUBS 0.007901f
C523 B.n217 VSUBS 0.007901f
C524 B.n218 VSUBS 0.007901f
C525 B.n219 VSUBS 0.007901f
C526 B.n220 VSUBS 0.007901f
C527 B.n221 VSUBS 0.007901f
C528 B.n222 VSUBS 0.007901f
C529 B.n223 VSUBS 0.007901f
C530 B.n224 VSUBS 0.007901f
C531 B.n225 VSUBS 0.007901f
C532 B.n226 VSUBS 0.007901f
C533 B.n227 VSUBS 0.007901f
C534 B.n228 VSUBS 0.007901f
C535 B.n229 VSUBS 0.007901f
C536 B.n230 VSUBS 0.007901f
C537 B.n231 VSUBS 0.007901f
C538 B.n232 VSUBS 0.007901f
C539 B.n233 VSUBS 0.007901f
C540 B.n234 VSUBS 0.007901f
C541 B.n235 VSUBS 0.007901f
C542 B.n236 VSUBS 0.007901f
C543 B.n237 VSUBS 0.007901f
C544 B.n238 VSUBS 0.007901f
C545 B.n239 VSUBS 0.007901f
C546 B.n240 VSUBS 0.019614f
C547 B.n241 VSUBS 0.019614f
C548 B.n242 VSUBS 0.01873f
C549 B.n243 VSUBS 0.007901f
C550 B.n244 VSUBS 0.007901f
C551 B.n245 VSUBS 0.007901f
C552 B.n246 VSUBS 0.007901f
C553 B.n247 VSUBS 0.007901f
C554 B.n248 VSUBS 0.007901f
C555 B.n249 VSUBS 0.007901f
C556 B.n250 VSUBS 0.007901f
C557 B.n251 VSUBS 0.007901f
C558 B.n252 VSUBS 0.007901f
C559 B.n253 VSUBS 0.007901f
C560 B.n254 VSUBS 0.007901f
C561 B.n255 VSUBS 0.007901f
C562 B.n256 VSUBS 0.007901f
C563 B.n257 VSUBS 0.007901f
C564 B.n258 VSUBS 0.007901f
C565 B.n259 VSUBS 0.007901f
C566 B.n260 VSUBS 0.007901f
C567 B.n261 VSUBS 0.007901f
C568 B.n262 VSUBS 0.007901f
C569 B.n263 VSUBS 0.007901f
C570 B.n264 VSUBS 0.007901f
C571 B.n265 VSUBS 0.007901f
C572 B.n266 VSUBS 0.007901f
C573 B.n267 VSUBS 0.007901f
C574 B.n268 VSUBS 0.007901f
C575 B.n269 VSUBS 0.007901f
C576 B.n270 VSUBS 0.007901f
C577 B.n271 VSUBS 0.007901f
C578 B.n272 VSUBS 0.007901f
C579 B.n273 VSUBS 0.007901f
C580 B.n274 VSUBS 0.007901f
C581 B.n275 VSUBS 0.007901f
C582 B.n276 VSUBS 0.007901f
C583 B.n277 VSUBS 0.007901f
C584 B.n278 VSUBS 0.007901f
C585 B.n279 VSUBS 0.007901f
C586 B.n280 VSUBS 0.007901f
C587 B.n281 VSUBS 0.007901f
C588 B.n282 VSUBS 0.007901f
C589 B.n283 VSUBS 0.007901f
C590 B.n284 VSUBS 0.007901f
C591 B.n285 VSUBS 0.007901f
C592 B.n286 VSUBS 0.007901f
C593 B.n287 VSUBS 0.007901f
C594 B.n288 VSUBS 0.007901f
C595 B.n289 VSUBS 0.007901f
C596 B.n290 VSUBS 0.007901f
C597 B.n291 VSUBS 0.007901f
C598 B.n292 VSUBS 0.007901f
C599 B.n293 VSUBS 0.007901f
C600 B.n294 VSUBS 0.007901f
C601 B.n295 VSUBS 0.007901f
C602 B.n296 VSUBS 0.007901f
C603 B.n297 VSUBS 0.007901f
C604 B.n298 VSUBS 0.007901f
C605 B.n299 VSUBS 0.007901f
C606 B.n300 VSUBS 0.007901f
C607 B.n301 VSUBS 0.007901f
C608 B.n302 VSUBS 0.007901f
C609 B.n303 VSUBS 0.007901f
C610 B.n304 VSUBS 0.007901f
C611 B.n305 VSUBS 0.007901f
C612 B.n306 VSUBS 0.007901f
C613 B.n307 VSUBS 0.007901f
C614 B.n308 VSUBS 0.007901f
C615 B.n309 VSUBS 0.007901f
C616 B.n310 VSUBS 0.007901f
C617 B.n311 VSUBS 0.007901f
C618 B.n312 VSUBS 0.007901f
C619 B.n313 VSUBS 0.007901f
C620 B.n314 VSUBS 0.007901f
C621 B.n315 VSUBS 0.007901f
C622 B.n316 VSUBS 0.007901f
C623 B.n317 VSUBS 0.019614f
C624 B.n318 VSUBS 0.01873f
C625 B.n319 VSUBS 0.019614f
C626 B.n320 VSUBS 0.007901f
C627 B.n321 VSUBS 0.007901f
C628 B.n322 VSUBS 0.007901f
C629 B.n323 VSUBS 0.007901f
C630 B.n324 VSUBS 0.007901f
C631 B.n325 VSUBS 0.007901f
C632 B.n326 VSUBS 0.007901f
C633 B.n327 VSUBS 0.007901f
C634 B.n328 VSUBS 0.007901f
C635 B.n329 VSUBS 0.007901f
C636 B.n330 VSUBS 0.007901f
C637 B.n331 VSUBS 0.007901f
C638 B.n332 VSUBS 0.007901f
C639 B.n333 VSUBS 0.007901f
C640 B.n334 VSUBS 0.007901f
C641 B.n335 VSUBS 0.007901f
C642 B.n336 VSUBS 0.007901f
C643 B.n337 VSUBS 0.007901f
C644 B.n338 VSUBS 0.007901f
C645 B.n339 VSUBS 0.007901f
C646 B.n340 VSUBS 0.007901f
C647 B.n341 VSUBS 0.007901f
C648 B.n342 VSUBS 0.007901f
C649 B.n343 VSUBS 0.007901f
C650 B.n344 VSUBS 0.007901f
C651 B.n345 VSUBS 0.007901f
C652 B.n346 VSUBS 0.007901f
C653 B.n347 VSUBS 0.007901f
C654 B.n348 VSUBS 0.007901f
C655 B.n349 VSUBS 0.007901f
C656 B.n350 VSUBS 0.007901f
C657 B.n351 VSUBS 0.007901f
C658 B.n352 VSUBS 0.007901f
C659 B.n353 VSUBS 0.005461f
C660 B.n354 VSUBS 0.018306f
C661 B.n355 VSUBS 0.006391f
C662 B.n356 VSUBS 0.007901f
C663 B.n357 VSUBS 0.007901f
C664 B.n358 VSUBS 0.007901f
C665 B.n359 VSUBS 0.007901f
C666 B.n360 VSUBS 0.007901f
C667 B.n361 VSUBS 0.007901f
C668 B.n362 VSUBS 0.007901f
C669 B.n363 VSUBS 0.007901f
C670 B.n364 VSUBS 0.007901f
C671 B.n365 VSUBS 0.007901f
C672 B.n366 VSUBS 0.007901f
C673 B.n367 VSUBS 0.006391f
C674 B.n368 VSUBS 0.007901f
C675 B.n369 VSUBS 0.007901f
C676 B.n370 VSUBS 0.007901f
C677 B.n371 VSUBS 0.007901f
C678 B.n372 VSUBS 0.007901f
C679 B.n373 VSUBS 0.007901f
C680 B.n374 VSUBS 0.007901f
C681 B.n375 VSUBS 0.007901f
C682 B.n376 VSUBS 0.007901f
C683 B.n377 VSUBS 0.007901f
C684 B.n378 VSUBS 0.007901f
C685 B.n379 VSUBS 0.007901f
C686 B.n380 VSUBS 0.007901f
C687 B.n381 VSUBS 0.007901f
C688 B.n382 VSUBS 0.007901f
C689 B.n383 VSUBS 0.007901f
C690 B.n384 VSUBS 0.007901f
C691 B.n385 VSUBS 0.007901f
C692 B.n386 VSUBS 0.007901f
C693 B.n387 VSUBS 0.007901f
C694 B.n388 VSUBS 0.007901f
C695 B.n389 VSUBS 0.007901f
C696 B.n390 VSUBS 0.007901f
C697 B.n391 VSUBS 0.007901f
C698 B.n392 VSUBS 0.007901f
C699 B.n393 VSUBS 0.007901f
C700 B.n394 VSUBS 0.007901f
C701 B.n395 VSUBS 0.007901f
C702 B.n396 VSUBS 0.007901f
C703 B.n397 VSUBS 0.007901f
C704 B.n398 VSUBS 0.007901f
C705 B.n399 VSUBS 0.007901f
C706 B.n400 VSUBS 0.007901f
C707 B.n401 VSUBS 0.007901f
C708 B.n402 VSUBS 0.007901f
C709 B.n403 VSUBS 0.019614f
C710 B.n404 VSUBS 0.019614f
C711 B.n405 VSUBS 0.01873f
C712 B.n406 VSUBS 0.007901f
C713 B.n407 VSUBS 0.007901f
C714 B.n408 VSUBS 0.007901f
C715 B.n409 VSUBS 0.007901f
C716 B.n410 VSUBS 0.007901f
C717 B.n411 VSUBS 0.007901f
C718 B.n412 VSUBS 0.007901f
C719 B.n413 VSUBS 0.007901f
C720 B.n414 VSUBS 0.007901f
C721 B.n415 VSUBS 0.007901f
C722 B.n416 VSUBS 0.007901f
C723 B.n417 VSUBS 0.007901f
C724 B.n418 VSUBS 0.007901f
C725 B.n419 VSUBS 0.007901f
C726 B.n420 VSUBS 0.007901f
C727 B.n421 VSUBS 0.007901f
C728 B.n422 VSUBS 0.007901f
C729 B.n423 VSUBS 0.007901f
C730 B.n424 VSUBS 0.007901f
C731 B.n425 VSUBS 0.007901f
C732 B.n426 VSUBS 0.007901f
C733 B.n427 VSUBS 0.007901f
C734 B.n428 VSUBS 0.007901f
C735 B.n429 VSUBS 0.007901f
C736 B.n430 VSUBS 0.007901f
C737 B.n431 VSUBS 0.007901f
C738 B.n432 VSUBS 0.007901f
C739 B.n433 VSUBS 0.007901f
C740 B.n434 VSUBS 0.007901f
C741 B.n435 VSUBS 0.007901f
C742 B.n436 VSUBS 0.007901f
C743 B.n437 VSUBS 0.007901f
C744 B.n438 VSUBS 0.007901f
C745 B.n439 VSUBS 0.007901f
C746 B.n440 VSUBS 0.007901f
C747 B.n441 VSUBS 0.007901f
C748 B.n442 VSUBS 0.007901f
C749 B.n443 VSUBS 0.017891f
.ends

