* NGSPICE file created from diff_pair_sample_1396.ext - technology: sky130A

.subckt diff_pair_sample_1396 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=2.4
X1 VTAIL.t4 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=2.4
X2 VTAIL.t7 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=2.4
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=2.4
X4 VDD1.t1 VP.t2 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=2.4
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=2.4
X6 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=2.4
X7 VTAIL.t6 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=2.4
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=2.4
X9 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=2.4
X10 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=2.4
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=2.4
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n3 105.252
R7 VP.n16 VP.n15 105.252
R8 VP.n4 VP.t3 95.7152
R9 VP.n4 VP.t0 94.9745
R10 VP.n3 VP.t1 61.0538
R11 VP.n15 VP.t2 61.0538
R12 VP.n9 VP.n1 56.5617
R13 VP.n5 VP.n4 45.8059
R14 VP.n8 VP.n7 24.5923
R15 VP.n9 VP.n8 24.5923
R16 VP.n13 VP.n1 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n3 5.65662
R19 VP.n15 VP.n14 5.65662
R20 VP.n6 VP.n5 0.278335
R21 VP.n16 VP.n0 0.278335
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153485
R28 VTAIL.n250 VTAIL.n224 289.615
R29 VTAIL.n26 VTAIL.n0 289.615
R30 VTAIL.n58 VTAIL.n32 289.615
R31 VTAIL.n90 VTAIL.n64 289.615
R32 VTAIL.n218 VTAIL.n192 289.615
R33 VTAIL.n186 VTAIL.n160 289.615
R34 VTAIL.n154 VTAIL.n128 289.615
R35 VTAIL.n122 VTAIL.n96 289.615
R36 VTAIL.n235 VTAIL.n234 185
R37 VTAIL.n232 VTAIL.n231 185
R38 VTAIL.n241 VTAIL.n240 185
R39 VTAIL.n243 VTAIL.n242 185
R40 VTAIL.n228 VTAIL.n227 185
R41 VTAIL.n249 VTAIL.n248 185
R42 VTAIL.n251 VTAIL.n250 185
R43 VTAIL.n11 VTAIL.n10 185
R44 VTAIL.n8 VTAIL.n7 185
R45 VTAIL.n17 VTAIL.n16 185
R46 VTAIL.n19 VTAIL.n18 185
R47 VTAIL.n4 VTAIL.n3 185
R48 VTAIL.n25 VTAIL.n24 185
R49 VTAIL.n27 VTAIL.n26 185
R50 VTAIL.n43 VTAIL.n42 185
R51 VTAIL.n40 VTAIL.n39 185
R52 VTAIL.n49 VTAIL.n48 185
R53 VTAIL.n51 VTAIL.n50 185
R54 VTAIL.n36 VTAIL.n35 185
R55 VTAIL.n57 VTAIL.n56 185
R56 VTAIL.n59 VTAIL.n58 185
R57 VTAIL.n75 VTAIL.n74 185
R58 VTAIL.n72 VTAIL.n71 185
R59 VTAIL.n81 VTAIL.n80 185
R60 VTAIL.n83 VTAIL.n82 185
R61 VTAIL.n68 VTAIL.n67 185
R62 VTAIL.n89 VTAIL.n88 185
R63 VTAIL.n91 VTAIL.n90 185
R64 VTAIL.n219 VTAIL.n218 185
R65 VTAIL.n217 VTAIL.n216 185
R66 VTAIL.n196 VTAIL.n195 185
R67 VTAIL.n211 VTAIL.n210 185
R68 VTAIL.n209 VTAIL.n208 185
R69 VTAIL.n200 VTAIL.n199 185
R70 VTAIL.n203 VTAIL.n202 185
R71 VTAIL.n187 VTAIL.n186 185
R72 VTAIL.n185 VTAIL.n184 185
R73 VTAIL.n164 VTAIL.n163 185
R74 VTAIL.n179 VTAIL.n178 185
R75 VTAIL.n177 VTAIL.n176 185
R76 VTAIL.n168 VTAIL.n167 185
R77 VTAIL.n171 VTAIL.n170 185
R78 VTAIL.n155 VTAIL.n154 185
R79 VTAIL.n153 VTAIL.n152 185
R80 VTAIL.n132 VTAIL.n131 185
R81 VTAIL.n147 VTAIL.n146 185
R82 VTAIL.n145 VTAIL.n144 185
R83 VTAIL.n136 VTAIL.n135 185
R84 VTAIL.n139 VTAIL.n138 185
R85 VTAIL.n123 VTAIL.n122 185
R86 VTAIL.n121 VTAIL.n120 185
R87 VTAIL.n100 VTAIL.n99 185
R88 VTAIL.n115 VTAIL.n114 185
R89 VTAIL.n113 VTAIL.n112 185
R90 VTAIL.n104 VTAIL.n103 185
R91 VTAIL.n107 VTAIL.n106 185
R92 VTAIL.t2 VTAIL.n233 147.661
R93 VTAIL.t1 VTAIL.n9 147.661
R94 VTAIL.t3 VTAIL.n41 147.661
R95 VTAIL.t4 VTAIL.n73 147.661
R96 VTAIL.t5 VTAIL.n201 147.661
R97 VTAIL.t6 VTAIL.n169 147.661
R98 VTAIL.t0 VTAIL.n137 147.661
R99 VTAIL.t7 VTAIL.n105 147.661
R100 VTAIL.n234 VTAIL.n231 104.615
R101 VTAIL.n241 VTAIL.n231 104.615
R102 VTAIL.n242 VTAIL.n241 104.615
R103 VTAIL.n242 VTAIL.n227 104.615
R104 VTAIL.n249 VTAIL.n227 104.615
R105 VTAIL.n250 VTAIL.n249 104.615
R106 VTAIL.n10 VTAIL.n7 104.615
R107 VTAIL.n17 VTAIL.n7 104.615
R108 VTAIL.n18 VTAIL.n17 104.615
R109 VTAIL.n18 VTAIL.n3 104.615
R110 VTAIL.n25 VTAIL.n3 104.615
R111 VTAIL.n26 VTAIL.n25 104.615
R112 VTAIL.n42 VTAIL.n39 104.615
R113 VTAIL.n49 VTAIL.n39 104.615
R114 VTAIL.n50 VTAIL.n49 104.615
R115 VTAIL.n50 VTAIL.n35 104.615
R116 VTAIL.n57 VTAIL.n35 104.615
R117 VTAIL.n58 VTAIL.n57 104.615
R118 VTAIL.n74 VTAIL.n71 104.615
R119 VTAIL.n81 VTAIL.n71 104.615
R120 VTAIL.n82 VTAIL.n81 104.615
R121 VTAIL.n82 VTAIL.n67 104.615
R122 VTAIL.n89 VTAIL.n67 104.615
R123 VTAIL.n90 VTAIL.n89 104.615
R124 VTAIL.n218 VTAIL.n217 104.615
R125 VTAIL.n217 VTAIL.n195 104.615
R126 VTAIL.n210 VTAIL.n195 104.615
R127 VTAIL.n210 VTAIL.n209 104.615
R128 VTAIL.n209 VTAIL.n199 104.615
R129 VTAIL.n202 VTAIL.n199 104.615
R130 VTAIL.n186 VTAIL.n185 104.615
R131 VTAIL.n185 VTAIL.n163 104.615
R132 VTAIL.n178 VTAIL.n163 104.615
R133 VTAIL.n178 VTAIL.n177 104.615
R134 VTAIL.n177 VTAIL.n167 104.615
R135 VTAIL.n170 VTAIL.n167 104.615
R136 VTAIL.n154 VTAIL.n153 104.615
R137 VTAIL.n153 VTAIL.n131 104.615
R138 VTAIL.n146 VTAIL.n131 104.615
R139 VTAIL.n146 VTAIL.n145 104.615
R140 VTAIL.n145 VTAIL.n135 104.615
R141 VTAIL.n138 VTAIL.n135 104.615
R142 VTAIL.n122 VTAIL.n121 104.615
R143 VTAIL.n121 VTAIL.n99 104.615
R144 VTAIL.n114 VTAIL.n99 104.615
R145 VTAIL.n114 VTAIL.n113 104.615
R146 VTAIL.n113 VTAIL.n103 104.615
R147 VTAIL.n106 VTAIL.n103 104.615
R148 VTAIL.n234 VTAIL.t2 52.3082
R149 VTAIL.n10 VTAIL.t1 52.3082
R150 VTAIL.n42 VTAIL.t3 52.3082
R151 VTAIL.n74 VTAIL.t4 52.3082
R152 VTAIL.n202 VTAIL.t5 52.3082
R153 VTAIL.n170 VTAIL.t6 52.3082
R154 VTAIL.n138 VTAIL.t0 52.3082
R155 VTAIL.n106 VTAIL.t7 52.3082
R156 VTAIL.n255 VTAIL.n254 33.7369
R157 VTAIL.n31 VTAIL.n30 33.7369
R158 VTAIL.n63 VTAIL.n62 33.7369
R159 VTAIL.n95 VTAIL.n94 33.7369
R160 VTAIL.n223 VTAIL.n222 33.7369
R161 VTAIL.n191 VTAIL.n190 33.7369
R162 VTAIL.n159 VTAIL.n158 33.7369
R163 VTAIL.n127 VTAIL.n126 33.7369
R164 VTAIL.n255 VTAIL.n223 19.9617
R165 VTAIL.n127 VTAIL.n95 19.9617
R166 VTAIL.n235 VTAIL.n233 15.6674
R167 VTAIL.n11 VTAIL.n9 15.6674
R168 VTAIL.n43 VTAIL.n41 15.6674
R169 VTAIL.n75 VTAIL.n73 15.6674
R170 VTAIL.n203 VTAIL.n201 15.6674
R171 VTAIL.n171 VTAIL.n169 15.6674
R172 VTAIL.n139 VTAIL.n137 15.6674
R173 VTAIL.n107 VTAIL.n105 15.6674
R174 VTAIL.n236 VTAIL.n232 12.8005
R175 VTAIL.n12 VTAIL.n8 12.8005
R176 VTAIL.n44 VTAIL.n40 12.8005
R177 VTAIL.n76 VTAIL.n72 12.8005
R178 VTAIL.n204 VTAIL.n200 12.8005
R179 VTAIL.n172 VTAIL.n168 12.8005
R180 VTAIL.n140 VTAIL.n136 12.8005
R181 VTAIL.n108 VTAIL.n104 12.8005
R182 VTAIL.n240 VTAIL.n239 12.0247
R183 VTAIL.n16 VTAIL.n15 12.0247
R184 VTAIL.n48 VTAIL.n47 12.0247
R185 VTAIL.n80 VTAIL.n79 12.0247
R186 VTAIL.n208 VTAIL.n207 12.0247
R187 VTAIL.n176 VTAIL.n175 12.0247
R188 VTAIL.n144 VTAIL.n143 12.0247
R189 VTAIL.n112 VTAIL.n111 12.0247
R190 VTAIL.n243 VTAIL.n230 11.249
R191 VTAIL.n19 VTAIL.n6 11.249
R192 VTAIL.n51 VTAIL.n38 11.249
R193 VTAIL.n83 VTAIL.n70 11.249
R194 VTAIL.n211 VTAIL.n198 11.249
R195 VTAIL.n179 VTAIL.n166 11.249
R196 VTAIL.n147 VTAIL.n134 11.249
R197 VTAIL.n115 VTAIL.n102 11.249
R198 VTAIL.n244 VTAIL.n228 10.4732
R199 VTAIL.n20 VTAIL.n4 10.4732
R200 VTAIL.n52 VTAIL.n36 10.4732
R201 VTAIL.n84 VTAIL.n68 10.4732
R202 VTAIL.n212 VTAIL.n196 10.4732
R203 VTAIL.n180 VTAIL.n164 10.4732
R204 VTAIL.n148 VTAIL.n132 10.4732
R205 VTAIL.n116 VTAIL.n100 10.4732
R206 VTAIL.n248 VTAIL.n247 9.69747
R207 VTAIL.n24 VTAIL.n23 9.69747
R208 VTAIL.n56 VTAIL.n55 9.69747
R209 VTAIL.n88 VTAIL.n87 9.69747
R210 VTAIL.n216 VTAIL.n215 9.69747
R211 VTAIL.n184 VTAIL.n183 9.69747
R212 VTAIL.n152 VTAIL.n151 9.69747
R213 VTAIL.n120 VTAIL.n119 9.69747
R214 VTAIL.n254 VTAIL.n253 9.45567
R215 VTAIL.n30 VTAIL.n29 9.45567
R216 VTAIL.n62 VTAIL.n61 9.45567
R217 VTAIL.n94 VTAIL.n93 9.45567
R218 VTAIL.n222 VTAIL.n221 9.45567
R219 VTAIL.n190 VTAIL.n189 9.45567
R220 VTAIL.n158 VTAIL.n157 9.45567
R221 VTAIL.n126 VTAIL.n125 9.45567
R222 VTAIL.n253 VTAIL.n252 9.3005
R223 VTAIL.n226 VTAIL.n225 9.3005
R224 VTAIL.n247 VTAIL.n246 9.3005
R225 VTAIL.n245 VTAIL.n244 9.3005
R226 VTAIL.n230 VTAIL.n229 9.3005
R227 VTAIL.n239 VTAIL.n238 9.3005
R228 VTAIL.n237 VTAIL.n236 9.3005
R229 VTAIL.n29 VTAIL.n28 9.3005
R230 VTAIL.n2 VTAIL.n1 9.3005
R231 VTAIL.n23 VTAIL.n22 9.3005
R232 VTAIL.n21 VTAIL.n20 9.3005
R233 VTAIL.n6 VTAIL.n5 9.3005
R234 VTAIL.n15 VTAIL.n14 9.3005
R235 VTAIL.n13 VTAIL.n12 9.3005
R236 VTAIL.n61 VTAIL.n60 9.3005
R237 VTAIL.n34 VTAIL.n33 9.3005
R238 VTAIL.n55 VTAIL.n54 9.3005
R239 VTAIL.n53 VTAIL.n52 9.3005
R240 VTAIL.n38 VTAIL.n37 9.3005
R241 VTAIL.n47 VTAIL.n46 9.3005
R242 VTAIL.n45 VTAIL.n44 9.3005
R243 VTAIL.n93 VTAIL.n92 9.3005
R244 VTAIL.n66 VTAIL.n65 9.3005
R245 VTAIL.n87 VTAIL.n86 9.3005
R246 VTAIL.n85 VTAIL.n84 9.3005
R247 VTAIL.n70 VTAIL.n69 9.3005
R248 VTAIL.n79 VTAIL.n78 9.3005
R249 VTAIL.n77 VTAIL.n76 9.3005
R250 VTAIL.n221 VTAIL.n220 9.3005
R251 VTAIL.n194 VTAIL.n193 9.3005
R252 VTAIL.n215 VTAIL.n214 9.3005
R253 VTAIL.n213 VTAIL.n212 9.3005
R254 VTAIL.n198 VTAIL.n197 9.3005
R255 VTAIL.n207 VTAIL.n206 9.3005
R256 VTAIL.n205 VTAIL.n204 9.3005
R257 VTAIL.n189 VTAIL.n188 9.3005
R258 VTAIL.n162 VTAIL.n161 9.3005
R259 VTAIL.n183 VTAIL.n182 9.3005
R260 VTAIL.n181 VTAIL.n180 9.3005
R261 VTAIL.n166 VTAIL.n165 9.3005
R262 VTAIL.n175 VTAIL.n174 9.3005
R263 VTAIL.n173 VTAIL.n172 9.3005
R264 VTAIL.n157 VTAIL.n156 9.3005
R265 VTAIL.n130 VTAIL.n129 9.3005
R266 VTAIL.n151 VTAIL.n150 9.3005
R267 VTAIL.n149 VTAIL.n148 9.3005
R268 VTAIL.n134 VTAIL.n133 9.3005
R269 VTAIL.n143 VTAIL.n142 9.3005
R270 VTAIL.n141 VTAIL.n140 9.3005
R271 VTAIL.n125 VTAIL.n124 9.3005
R272 VTAIL.n98 VTAIL.n97 9.3005
R273 VTAIL.n119 VTAIL.n118 9.3005
R274 VTAIL.n117 VTAIL.n116 9.3005
R275 VTAIL.n102 VTAIL.n101 9.3005
R276 VTAIL.n111 VTAIL.n110 9.3005
R277 VTAIL.n109 VTAIL.n108 9.3005
R278 VTAIL.n251 VTAIL.n226 8.92171
R279 VTAIL.n27 VTAIL.n2 8.92171
R280 VTAIL.n59 VTAIL.n34 8.92171
R281 VTAIL.n91 VTAIL.n66 8.92171
R282 VTAIL.n219 VTAIL.n194 8.92171
R283 VTAIL.n187 VTAIL.n162 8.92171
R284 VTAIL.n155 VTAIL.n130 8.92171
R285 VTAIL.n123 VTAIL.n98 8.92171
R286 VTAIL.n252 VTAIL.n224 8.14595
R287 VTAIL.n28 VTAIL.n0 8.14595
R288 VTAIL.n60 VTAIL.n32 8.14595
R289 VTAIL.n92 VTAIL.n64 8.14595
R290 VTAIL.n220 VTAIL.n192 8.14595
R291 VTAIL.n188 VTAIL.n160 8.14595
R292 VTAIL.n156 VTAIL.n128 8.14595
R293 VTAIL.n124 VTAIL.n96 8.14595
R294 VTAIL.n254 VTAIL.n224 5.81868
R295 VTAIL.n30 VTAIL.n0 5.81868
R296 VTAIL.n62 VTAIL.n32 5.81868
R297 VTAIL.n94 VTAIL.n64 5.81868
R298 VTAIL.n222 VTAIL.n192 5.81868
R299 VTAIL.n190 VTAIL.n160 5.81868
R300 VTAIL.n158 VTAIL.n128 5.81868
R301 VTAIL.n126 VTAIL.n96 5.81868
R302 VTAIL.n252 VTAIL.n251 5.04292
R303 VTAIL.n28 VTAIL.n27 5.04292
R304 VTAIL.n60 VTAIL.n59 5.04292
R305 VTAIL.n92 VTAIL.n91 5.04292
R306 VTAIL.n220 VTAIL.n219 5.04292
R307 VTAIL.n188 VTAIL.n187 5.04292
R308 VTAIL.n156 VTAIL.n155 5.04292
R309 VTAIL.n124 VTAIL.n123 5.04292
R310 VTAIL.n237 VTAIL.n233 4.38594
R311 VTAIL.n13 VTAIL.n9 4.38594
R312 VTAIL.n45 VTAIL.n41 4.38594
R313 VTAIL.n77 VTAIL.n73 4.38594
R314 VTAIL.n205 VTAIL.n201 4.38594
R315 VTAIL.n173 VTAIL.n169 4.38594
R316 VTAIL.n141 VTAIL.n137 4.38594
R317 VTAIL.n109 VTAIL.n105 4.38594
R318 VTAIL.n248 VTAIL.n226 4.26717
R319 VTAIL.n24 VTAIL.n2 4.26717
R320 VTAIL.n56 VTAIL.n34 4.26717
R321 VTAIL.n88 VTAIL.n66 4.26717
R322 VTAIL.n216 VTAIL.n194 4.26717
R323 VTAIL.n184 VTAIL.n162 4.26717
R324 VTAIL.n152 VTAIL.n130 4.26717
R325 VTAIL.n120 VTAIL.n98 4.26717
R326 VTAIL.n247 VTAIL.n228 3.49141
R327 VTAIL.n23 VTAIL.n4 3.49141
R328 VTAIL.n55 VTAIL.n36 3.49141
R329 VTAIL.n87 VTAIL.n68 3.49141
R330 VTAIL.n215 VTAIL.n196 3.49141
R331 VTAIL.n183 VTAIL.n164 3.49141
R332 VTAIL.n151 VTAIL.n132 3.49141
R333 VTAIL.n119 VTAIL.n100 3.49141
R334 VTAIL.n244 VTAIL.n243 2.71565
R335 VTAIL.n20 VTAIL.n19 2.71565
R336 VTAIL.n52 VTAIL.n51 2.71565
R337 VTAIL.n84 VTAIL.n83 2.71565
R338 VTAIL.n212 VTAIL.n211 2.71565
R339 VTAIL.n180 VTAIL.n179 2.71565
R340 VTAIL.n148 VTAIL.n147 2.71565
R341 VTAIL.n116 VTAIL.n115 2.71565
R342 VTAIL.n159 VTAIL.n127 2.35395
R343 VTAIL.n223 VTAIL.n191 2.35395
R344 VTAIL.n95 VTAIL.n63 2.35395
R345 VTAIL.n240 VTAIL.n230 1.93989
R346 VTAIL.n16 VTAIL.n6 1.93989
R347 VTAIL.n48 VTAIL.n38 1.93989
R348 VTAIL.n80 VTAIL.n70 1.93989
R349 VTAIL.n208 VTAIL.n198 1.93989
R350 VTAIL.n176 VTAIL.n166 1.93989
R351 VTAIL.n144 VTAIL.n134 1.93989
R352 VTAIL.n112 VTAIL.n102 1.93989
R353 VTAIL VTAIL.n31 1.23541
R354 VTAIL.n239 VTAIL.n232 1.16414
R355 VTAIL.n15 VTAIL.n8 1.16414
R356 VTAIL.n47 VTAIL.n40 1.16414
R357 VTAIL.n79 VTAIL.n72 1.16414
R358 VTAIL.n207 VTAIL.n200 1.16414
R359 VTAIL.n175 VTAIL.n168 1.16414
R360 VTAIL.n143 VTAIL.n136 1.16414
R361 VTAIL.n111 VTAIL.n104 1.16414
R362 VTAIL VTAIL.n255 1.11903
R363 VTAIL.n191 VTAIL.n159 0.470328
R364 VTAIL.n63 VTAIL.n31 0.470328
R365 VTAIL.n236 VTAIL.n235 0.388379
R366 VTAIL.n12 VTAIL.n11 0.388379
R367 VTAIL.n44 VTAIL.n43 0.388379
R368 VTAIL.n76 VTAIL.n75 0.388379
R369 VTAIL.n204 VTAIL.n203 0.388379
R370 VTAIL.n172 VTAIL.n171 0.388379
R371 VTAIL.n140 VTAIL.n139 0.388379
R372 VTAIL.n108 VTAIL.n107 0.388379
R373 VTAIL.n238 VTAIL.n237 0.155672
R374 VTAIL.n238 VTAIL.n229 0.155672
R375 VTAIL.n245 VTAIL.n229 0.155672
R376 VTAIL.n246 VTAIL.n245 0.155672
R377 VTAIL.n246 VTAIL.n225 0.155672
R378 VTAIL.n253 VTAIL.n225 0.155672
R379 VTAIL.n14 VTAIL.n13 0.155672
R380 VTAIL.n14 VTAIL.n5 0.155672
R381 VTAIL.n21 VTAIL.n5 0.155672
R382 VTAIL.n22 VTAIL.n21 0.155672
R383 VTAIL.n22 VTAIL.n1 0.155672
R384 VTAIL.n29 VTAIL.n1 0.155672
R385 VTAIL.n46 VTAIL.n45 0.155672
R386 VTAIL.n46 VTAIL.n37 0.155672
R387 VTAIL.n53 VTAIL.n37 0.155672
R388 VTAIL.n54 VTAIL.n53 0.155672
R389 VTAIL.n54 VTAIL.n33 0.155672
R390 VTAIL.n61 VTAIL.n33 0.155672
R391 VTAIL.n78 VTAIL.n77 0.155672
R392 VTAIL.n78 VTAIL.n69 0.155672
R393 VTAIL.n85 VTAIL.n69 0.155672
R394 VTAIL.n86 VTAIL.n85 0.155672
R395 VTAIL.n86 VTAIL.n65 0.155672
R396 VTAIL.n93 VTAIL.n65 0.155672
R397 VTAIL.n221 VTAIL.n193 0.155672
R398 VTAIL.n214 VTAIL.n193 0.155672
R399 VTAIL.n214 VTAIL.n213 0.155672
R400 VTAIL.n213 VTAIL.n197 0.155672
R401 VTAIL.n206 VTAIL.n197 0.155672
R402 VTAIL.n206 VTAIL.n205 0.155672
R403 VTAIL.n189 VTAIL.n161 0.155672
R404 VTAIL.n182 VTAIL.n161 0.155672
R405 VTAIL.n182 VTAIL.n181 0.155672
R406 VTAIL.n181 VTAIL.n165 0.155672
R407 VTAIL.n174 VTAIL.n165 0.155672
R408 VTAIL.n174 VTAIL.n173 0.155672
R409 VTAIL.n157 VTAIL.n129 0.155672
R410 VTAIL.n150 VTAIL.n129 0.155672
R411 VTAIL.n150 VTAIL.n149 0.155672
R412 VTAIL.n149 VTAIL.n133 0.155672
R413 VTAIL.n142 VTAIL.n133 0.155672
R414 VTAIL.n142 VTAIL.n141 0.155672
R415 VTAIL.n125 VTAIL.n97 0.155672
R416 VTAIL.n118 VTAIL.n97 0.155672
R417 VTAIL.n118 VTAIL.n117 0.155672
R418 VTAIL.n117 VTAIL.n101 0.155672
R419 VTAIL.n110 VTAIL.n101 0.155672
R420 VTAIL.n110 VTAIL.n109 0.155672
R421 VDD1 VDD1.n1 105.284
R422 VDD1 VDD1.n0 68.8004
R423 VDD1.n0 VDD1.t0 3.25708
R424 VDD1.n0 VDD1.t3 3.25708
R425 VDD1.n1 VDD1.t2 3.25708
R426 VDD1.n1 VDD1.t1 3.25708
R427 B.n558 B.n557 585
R428 B.n207 B.n90 585
R429 B.n206 B.n205 585
R430 B.n204 B.n203 585
R431 B.n202 B.n201 585
R432 B.n200 B.n199 585
R433 B.n198 B.n197 585
R434 B.n196 B.n195 585
R435 B.n194 B.n193 585
R436 B.n192 B.n191 585
R437 B.n190 B.n189 585
R438 B.n188 B.n187 585
R439 B.n186 B.n185 585
R440 B.n184 B.n183 585
R441 B.n182 B.n181 585
R442 B.n180 B.n179 585
R443 B.n178 B.n177 585
R444 B.n176 B.n175 585
R445 B.n174 B.n173 585
R446 B.n172 B.n171 585
R447 B.n170 B.n169 585
R448 B.n168 B.n167 585
R449 B.n166 B.n165 585
R450 B.n164 B.n163 585
R451 B.n162 B.n161 585
R452 B.n160 B.n159 585
R453 B.n158 B.n157 585
R454 B.n156 B.n155 585
R455 B.n154 B.n153 585
R456 B.n152 B.n151 585
R457 B.n150 B.n149 585
R458 B.n148 B.n147 585
R459 B.n146 B.n145 585
R460 B.n144 B.n143 585
R461 B.n142 B.n141 585
R462 B.n140 B.n139 585
R463 B.n138 B.n137 585
R464 B.n136 B.n135 585
R465 B.n134 B.n133 585
R466 B.n132 B.n131 585
R467 B.n130 B.n129 585
R468 B.n128 B.n127 585
R469 B.n126 B.n125 585
R470 B.n124 B.n123 585
R471 B.n122 B.n121 585
R472 B.n120 B.n119 585
R473 B.n118 B.n117 585
R474 B.n116 B.n115 585
R475 B.n114 B.n113 585
R476 B.n112 B.n111 585
R477 B.n110 B.n109 585
R478 B.n108 B.n107 585
R479 B.n106 B.n105 585
R480 B.n104 B.n103 585
R481 B.n102 B.n101 585
R482 B.n100 B.n99 585
R483 B.n98 B.n97 585
R484 B.n60 B.n59 585
R485 B.n556 B.n61 585
R486 B.n561 B.n61 585
R487 B.n555 B.n554 585
R488 B.n554 B.n57 585
R489 B.n553 B.n56 585
R490 B.n567 B.n56 585
R491 B.n552 B.n55 585
R492 B.n568 B.n55 585
R493 B.n551 B.n54 585
R494 B.n569 B.n54 585
R495 B.n550 B.n549 585
R496 B.n549 B.n50 585
R497 B.n548 B.n49 585
R498 B.n575 B.n49 585
R499 B.n547 B.n48 585
R500 B.n576 B.n48 585
R501 B.n546 B.n47 585
R502 B.n577 B.n47 585
R503 B.n545 B.n544 585
R504 B.n544 B.n43 585
R505 B.n543 B.n42 585
R506 B.n583 B.n42 585
R507 B.n542 B.n41 585
R508 B.n584 B.n41 585
R509 B.n541 B.n40 585
R510 B.n585 B.n40 585
R511 B.n540 B.n539 585
R512 B.n539 B.n36 585
R513 B.n538 B.n35 585
R514 B.n591 B.n35 585
R515 B.n537 B.n34 585
R516 B.n592 B.n34 585
R517 B.n536 B.n33 585
R518 B.n593 B.n33 585
R519 B.n535 B.n534 585
R520 B.n534 B.n29 585
R521 B.n533 B.n28 585
R522 B.n599 B.n28 585
R523 B.n532 B.n27 585
R524 B.n600 B.n27 585
R525 B.n531 B.n26 585
R526 B.n601 B.n26 585
R527 B.n530 B.n529 585
R528 B.n529 B.n22 585
R529 B.n528 B.n21 585
R530 B.n607 B.n21 585
R531 B.n527 B.n20 585
R532 B.n608 B.n20 585
R533 B.n526 B.n19 585
R534 B.n609 B.n19 585
R535 B.n525 B.n524 585
R536 B.n524 B.n15 585
R537 B.n523 B.n14 585
R538 B.n615 B.n14 585
R539 B.n522 B.n13 585
R540 B.n616 B.n13 585
R541 B.n521 B.n12 585
R542 B.n617 B.n12 585
R543 B.n520 B.n519 585
R544 B.n519 B.n8 585
R545 B.n518 B.n7 585
R546 B.n623 B.n7 585
R547 B.n517 B.n6 585
R548 B.n624 B.n6 585
R549 B.n516 B.n5 585
R550 B.n625 B.n5 585
R551 B.n515 B.n514 585
R552 B.n514 B.n4 585
R553 B.n513 B.n208 585
R554 B.n513 B.n512 585
R555 B.n503 B.n209 585
R556 B.n210 B.n209 585
R557 B.n505 B.n504 585
R558 B.n506 B.n505 585
R559 B.n502 B.n215 585
R560 B.n215 B.n214 585
R561 B.n501 B.n500 585
R562 B.n500 B.n499 585
R563 B.n217 B.n216 585
R564 B.n218 B.n217 585
R565 B.n492 B.n491 585
R566 B.n493 B.n492 585
R567 B.n490 B.n223 585
R568 B.n223 B.n222 585
R569 B.n489 B.n488 585
R570 B.n488 B.n487 585
R571 B.n225 B.n224 585
R572 B.n226 B.n225 585
R573 B.n480 B.n479 585
R574 B.n481 B.n480 585
R575 B.n478 B.n231 585
R576 B.n231 B.n230 585
R577 B.n477 B.n476 585
R578 B.n476 B.n475 585
R579 B.n233 B.n232 585
R580 B.n234 B.n233 585
R581 B.n468 B.n467 585
R582 B.n469 B.n468 585
R583 B.n466 B.n239 585
R584 B.n239 B.n238 585
R585 B.n465 B.n464 585
R586 B.n464 B.n463 585
R587 B.n241 B.n240 585
R588 B.n242 B.n241 585
R589 B.n456 B.n455 585
R590 B.n457 B.n456 585
R591 B.n454 B.n247 585
R592 B.n247 B.n246 585
R593 B.n453 B.n452 585
R594 B.n452 B.n451 585
R595 B.n249 B.n248 585
R596 B.n250 B.n249 585
R597 B.n444 B.n443 585
R598 B.n445 B.n444 585
R599 B.n442 B.n254 585
R600 B.n258 B.n254 585
R601 B.n441 B.n440 585
R602 B.n440 B.n439 585
R603 B.n256 B.n255 585
R604 B.n257 B.n256 585
R605 B.n432 B.n431 585
R606 B.n433 B.n432 585
R607 B.n430 B.n263 585
R608 B.n263 B.n262 585
R609 B.n429 B.n428 585
R610 B.n428 B.n427 585
R611 B.n265 B.n264 585
R612 B.n266 B.n265 585
R613 B.n420 B.n419 585
R614 B.n421 B.n420 585
R615 B.n269 B.n268 585
R616 B.n304 B.n302 585
R617 B.n305 B.n301 585
R618 B.n305 B.n270 585
R619 B.n308 B.n307 585
R620 B.n309 B.n300 585
R621 B.n311 B.n310 585
R622 B.n313 B.n299 585
R623 B.n316 B.n315 585
R624 B.n317 B.n298 585
R625 B.n319 B.n318 585
R626 B.n321 B.n297 585
R627 B.n324 B.n323 585
R628 B.n325 B.n296 585
R629 B.n327 B.n326 585
R630 B.n329 B.n295 585
R631 B.n332 B.n331 585
R632 B.n333 B.n294 585
R633 B.n335 B.n334 585
R634 B.n337 B.n293 585
R635 B.n340 B.n339 585
R636 B.n341 B.n292 585
R637 B.n343 B.n342 585
R638 B.n345 B.n291 585
R639 B.n348 B.n347 585
R640 B.n350 B.n288 585
R641 B.n352 B.n351 585
R642 B.n354 B.n287 585
R643 B.n357 B.n356 585
R644 B.n358 B.n286 585
R645 B.n360 B.n359 585
R646 B.n362 B.n285 585
R647 B.n365 B.n364 585
R648 B.n366 B.n284 585
R649 B.n371 B.n370 585
R650 B.n373 B.n283 585
R651 B.n376 B.n375 585
R652 B.n377 B.n282 585
R653 B.n379 B.n378 585
R654 B.n381 B.n281 585
R655 B.n384 B.n383 585
R656 B.n385 B.n280 585
R657 B.n387 B.n386 585
R658 B.n389 B.n279 585
R659 B.n392 B.n391 585
R660 B.n393 B.n278 585
R661 B.n395 B.n394 585
R662 B.n397 B.n277 585
R663 B.n400 B.n399 585
R664 B.n401 B.n276 585
R665 B.n403 B.n402 585
R666 B.n405 B.n275 585
R667 B.n408 B.n407 585
R668 B.n409 B.n274 585
R669 B.n411 B.n410 585
R670 B.n413 B.n273 585
R671 B.n414 B.n272 585
R672 B.n417 B.n416 585
R673 B.n418 B.n271 585
R674 B.n271 B.n270 585
R675 B.n423 B.n422 585
R676 B.n422 B.n421 585
R677 B.n424 B.n267 585
R678 B.n267 B.n266 585
R679 B.n426 B.n425 585
R680 B.n427 B.n426 585
R681 B.n261 B.n260 585
R682 B.n262 B.n261 585
R683 B.n435 B.n434 585
R684 B.n434 B.n433 585
R685 B.n436 B.n259 585
R686 B.n259 B.n257 585
R687 B.n438 B.n437 585
R688 B.n439 B.n438 585
R689 B.n253 B.n252 585
R690 B.n258 B.n253 585
R691 B.n447 B.n446 585
R692 B.n446 B.n445 585
R693 B.n448 B.n251 585
R694 B.n251 B.n250 585
R695 B.n450 B.n449 585
R696 B.n451 B.n450 585
R697 B.n245 B.n244 585
R698 B.n246 B.n245 585
R699 B.n459 B.n458 585
R700 B.n458 B.n457 585
R701 B.n460 B.n243 585
R702 B.n243 B.n242 585
R703 B.n462 B.n461 585
R704 B.n463 B.n462 585
R705 B.n237 B.n236 585
R706 B.n238 B.n237 585
R707 B.n471 B.n470 585
R708 B.n470 B.n469 585
R709 B.n472 B.n235 585
R710 B.n235 B.n234 585
R711 B.n474 B.n473 585
R712 B.n475 B.n474 585
R713 B.n229 B.n228 585
R714 B.n230 B.n229 585
R715 B.n483 B.n482 585
R716 B.n482 B.n481 585
R717 B.n484 B.n227 585
R718 B.n227 B.n226 585
R719 B.n486 B.n485 585
R720 B.n487 B.n486 585
R721 B.n221 B.n220 585
R722 B.n222 B.n221 585
R723 B.n495 B.n494 585
R724 B.n494 B.n493 585
R725 B.n496 B.n219 585
R726 B.n219 B.n218 585
R727 B.n498 B.n497 585
R728 B.n499 B.n498 585
R729 B.n213 B.n212 585
R730 B.n214 B.n213 585
R731 B.n508 B.n507 585
R732 B.n507 B.n506 585
R733 B.n509 B.n211 585
R734 B.n211 B.n210 585
R735 B.n511 B.n510 585
R736 B.n512 B.n511 585
R737 B.n2 B.n0 585
R738 B.n4 B.n2 585
R739 B.n3 B.n1 585
R740 B.n624 B.n3 585
R741 B.n622 B.n621 585
R742 B.n623 B.n622 585
R743 B.n620 B.n9 585
R744 B.n9 B.n8 585
R745 B.n619 B.n618 585
R746 B.n618 B.n617 585
R747 B.n11 B.n10 585
R748 B.n616 B.n11 585
R749 B.n614 B.n613 585
R750 B.n615 B.n614 585
R751 B.n612 B.n16 585
R752 B.n16 B.n15 585
R753 B.n611 B.n610 585
R754 B.n610 B.n609 585
R755 B.n18 B.n17 585
R756 B.n608 B.n18 585
R757 B.n606 B.n605 585
R758 B.n607 B.n606 585
R759 B.n604 B.n23 585
R760 B.n23 B.n22 585
R761 B.n603 B.n602 585
R762 B.n602 B.n601 585
R763 B.n25 B.n24 585
R764 B.n600 B.n25 585
R765 B.n598 B.n597 585
R766 B.n599 B.n598 585
R767 B.n596 B.n30 585
R768 B.n30 B.n29 585
R769 B.n595 B.n594 585
R770 B.n594 B.n593 585
R771 B.n32 B.n31 585
R772 B.n592 B.n32 585
R773 B.n590 B.n589 585
R774 B.n591 B.n590 585
R775 B.n588 B.n37 585
R776 B.n37 B.n36 585
R777 B.n587 B.n586 585
R778 B.n586 B.n585 585
R779 B.n39 B.n38 585
R780 B.n584 B.n39 585
R781 B.n582 B.n581 585
R782 B.n583 B.n582 585
R783 B.n580 B.n44 585
R784 B.n44 B.n43 585
R785 B.n579 B.n578 585
R786 B.n578 B.n577 585
R787 B.n46 B.n45 585
R788 B.n576 B.n46 585
R789 B.n574 B.n573 585
R790 B.n575 B.n574 585
R791 B.n572 B.n51 585
R792 B.n51 B.n50 585
R793 B.n571 B.n570 585
R794 B.n570 B.n569 585
R795 B.n53 B.n52 585
R796 B.n568 B.n53 585
R797 B.n566 B.n565 585
R798 B.n567 B.n566 585
R799 B.n564 B.n58 585
R800 B.n58 B.n57 585
R801 B.n563 B.n562 585
R802 B.n562 B.n561 585
R803 B.n627 B.n626 585
R804 B.n626 B.n625 585
R805 B.n422 B.n269 530.939
R806 B.n562 B.n60 530.939
R807 B.n420 B.n271 530.939
R808 B.n558 B.n61 530.939
R809 B.n367 B.t4 268.777
R810 B.n289 B.t8 268.777
R811 B.n94 B.t11 268.777
R812 B.n91 B.t15 268.777
R813 B.n560 B.n559 256.663
R814 B.n560 B.n89 256.663
R815 B.n560 B.n88 256.663
R816 B.n560 B.n87 256.663
R817 B.n560 B.n86 256.663
R818 B.n560 B.n85 256.663
R819 B.n560 B.n84 256.663
R820 B.n560 B.n83 256.663
R821 B.n560 B.n82 256.663
R822 B.n560 B.n81 256.663
R823 B.n560 B.n80 256.663
R824 B.n560 B.n79 256.663
R825 B.n560 B.n78 256.663
R826 B.n560 B.n77 256.663
R827 B.n560 B.n76 256.663
R828 B.n560 B.n75 256.663
R829 B.n560 B.n74 256.663
R830 B.n560 B.n73 256.663
R831 B.n560 B.n72 256.663
R832 B.n560 B.n71 256.663
R833 B.n560 B.n70 256.663
R834 B.n560 B.n69 256.663
R835 B.n560 B.n68 256.663
R836 B.n560 B.n67 256.663
R837 B.n560 B.n66 256.663
R838 B.n560 B.n65 256.663
R839 B.n560 B.n64 256.663
R840 B.n560 B.n63 256.663
R841 B.n560 B.n62 256.663
R842 B.n303 B.n270 256.663
R843 B.n306 B.n270 256.663
R844 B.n312 B.n270 256.663
R845 B.n314 B.n270 256.663
R846 B.n320 B.n270 256.663
R847 B.n322 B.n270 256.663
R848 B.n328 B.n270 256.663
R849 B.n330 B.n270 256.663
R850 B.n336 B.n270 256.663
R851 B.n338 B.n270 256.663
R852 B.n344 B.n270 256.663
R853 B.n346 B.n270 256.663
R854 B.n353 B.n270 256.663
R855 B.n355 B.n270 256.663
R856 B.n361 B.n270 256.663
R857 B.n363 B.n270 256.663
R858 B.n372 B.n270 256.663
R859 B.n374 B.n270 256.663
R860 B.n380 B.n270 256.663
R861 B.n382 B.n270 256.663
R862 B.n388 B.n270 256.663
R863 B.n390 B.n270 256.663
R864 B.n396 B.n270 256.663
R865 B.n398 B.n270 256.663
R866 B.n404 B.n270 256.663
R867 B.n406 B.n270 256.663
R868 B.n412 B.n270 256.663
R869 B.n415 B.n270 256.663
R870 B.n367 B.t7 233.483
R871 B.n91 B.t16 233.483
R872 B.n289 B.t10 233.483
R873 B.n94 B.t13 233.483
R874 B.n368 B.t6 180.538
R875 B.n92 B.t17 180.538
R876 B.n290 B.t9 180.538
R877 B.n95 B.t14 180.538
R878 B.n422 B.n267 163.367
R879 B.n426 B.n267 163.367
R880 B.n426 B.n261 163.367
R881 B.n434 B.n261 163.367
R882 B.n434 B.n259 163.367
R883 B.n438 B.n259 163.367
R884 B.n438 B.n253 163.367
R885 B.n446 B.n253 163.367
R886 B.n446 B.n251 163.367
R887 B.n450 B.n251 163.367
R888 B.n450 B.n245 163.367
R889 B.n458 B.n245 163.367
R890 B.n458 B.n243 163.367
R891 B.n462 B.n243 163.367
R892 B.n462 B.n237 163.367
R893 B.n470 B.n237 163.367
R894 B.n470 B.n235 163.367
R895 B.n474 B.n235 163.367
R896 B.n474 B.n229 163.367
R897 B.n482 B.n229 163.367
R898 B.n482 B.n227 163.367
R899 B.n486 B.n227 163.367
R900 B.n486 B.n221 163.367
R901 B.n494 B.n221 163.367
R902 B.n494 B.n219 163.367
R903 B.n498 B.n219 163.367
R904 B.n498 B.n213 163.367
R905 B.n507 B.n213 163.367
R906 B.n507 B.n211 163.367
R907 B.n511 B.n211 163.367
R908 B.n511 B.n2 163.367
R909 B.n626 B.n2 163.367
R910 B.n626 B.n3 163.367
R911 B.n622 B.n3 163.367
R912 B.n622 B.n9 163.367
R913 B.n618 B.n9 163.367
R914 B.n618 B.n11 163.367
R915 B.n614 B.n11 163.367
R916 B.n614 B.n16 163.367
R917 B.n610 B.n16 163.367
R918 B.n610 B.n18 163.367
R919 B.n606 B.n18 163.367
R920 B.n606 B.n23 163.367
R921 B.n602 B.n23 163.367
R922 B.n602 B.n25 163.367
R923 B.n598 B.n25 163.367
R924 B.n598 B.n30 163.367
R925 B.n594 B.n30 163.367
R926 B.n594 B.n32 163.367
R927 B.n590 B.n32 163.367
R928 B.n590 B.n37 163.367
R929 B.n586 B.n37 163.367
R930 B.n586 B.n39 163.367
R931 B.n582 B.n39 163.367
R932 B.n582 B.n44 163.367
R933 B.n578 B.n44 163.367
R934 B.n578 B.n46 163.367
R935 B.n574 B.n46 163.367
R936 B.n574 B.n51 163.367
R937 B.n570 B.n51 163.367
R938 B.n570 B.n53 163.367
R939 B.n566 B.n53 163.367
R940 B.n566 B.n58 163.367
R941 B.n562 B.n58 163.367
R942 B.n305 B.n304 163.367
R943 B.n307 B.n305 163.367
R944 B.n311 B.n300 163.367
R945 B.n315 B.n313 163.367
R946 B.n319 B.n298 163.367
R947 B.n323 B.n321 163.367
R948 B.n327 B.n296 163.367
R949 B.n331 B.n329 163.367
R950 B.n335 B.n294 163.367
R951 B.n339 B.n337 163.367
R952 B.n343 B.n292 163.367
R953 B.n347 B.n345 163.367
R954 B.n352 B.n288 163.367
R955 B.n356 B.n354 163.367
R956 B.n360 B.n286 163.367
R957 B.n364 B.n362 163.367
R958 B.n371 B.n284 163.367
R959 B.n375 B.n373 163.367
R960 B.n379 B.n282 163.367
R961 B.n383 B.n381 163.367
R962 B.n387 B.n280 163.367
R963 B.n391 B.n389 163.367
R964 B.n395 B.n278 163.367
R965 B.n399 B.n397 163.367
R966 B.n403 B.n276 163.367
R967 B.n407 B.n405 163.367
R968 B.n411 B.n274 163.367
R969 B.n414 B.n413 163.367
R970 B.n416 B.n271 163.367
R971 B.n420 B.n265 163.367
R972 B.n428 B.n265 163.367
R973 B.n428 B.n263 163.367
R974 B.n432 B.n263 163.367
R975 B.n432 B.n256 163.367
R976 B.n440 B.n256 163.367
R977 B.n440 B.n254 163.367
R978 B.n444 B.n254 163.367
R979 B.n444 B.n249 163.367
R980 B.n452 B.n249 163.367
R981 B.n452 B.n247 163.367
R982 B.n456 B.n247 163.367
R983 B.n456 B.n241 163.367
R984 B.n464 B.n241 163.367
R985 B.n464 B.n239 163.367
R986 B.n468 B.n239 163.367
R987 B.n468 B.n233 163.367
R988 B.n476 B.n233 163.367
R989 B.n476 B.n231 163.367
R990 B.n480 B.n231 163.367
R991 B.n480 B.n225 163.367
R992 B.n488 B.n225 163.367
R993 B.n488 B.n223 163.367
R994 B.n492 B.n223 163.367
R995 B.n492 B.n217 163.367
R996 B.n500 B.n217 163.367
R997 B.n500 B.n215 163.367
R998 B.n505 B.n215 163.367
R999 B.n505 B.n209 163.367
R1000 B.n513 B.n209 163.367
R1001 B.n514 B.n513 163.367
R1002 B.n514 B.n5 163.367
R1003 B.n6 B.n5 163.367
R1004 B.n7 B.n6 163.367
R1005 B.n519 B.n7 163.367
R1006 B.n519 B.n12 163.367
R1007 B.n13 B.n12 163.367
R1008 B.n14 B.n13 163.367
R1009 B.n524 B.n14 163.367
R1010 B.n524 B.n19 163.367
R1011 B.n20 B.n19 163.367
R1012 B.n21 B.n20 163.367
R1013 B.n529 B.n21 163.367
R1014 B.n529 B.n26 163.367
R1015 B.n27 B.n26 163.367
R1016 B.n28 B.n27 163.367
R1017 B.n534 B.n28 163.367
R1018 B.n534 B.n33 163.367
R1019 B.n34 B.n33 163.367
R1020 B.n35 B.n34 163.367
R1021 B.n539 B.n35 163.367
R1022 B.n539 B.n40 163.367
R1023 B.n41 B.n40 163.367
R1024 B.n42 B.n41 163.367
R1025 B.n544 B.n42 163.367
R1026 B.n544 B.n47 163.367
R1027 B.n48 B.n47 163.367
R1028 B.n49 B.n48 163.367
R1029 B.n549 B.n49 163.367
R1030 B.n549 B.n54 163.367
R1031 B.n55 B.n54 163.367
R1032 B.n56 B.n55 163.367
R1033 B.n554 B.n56 163.367
R1034 B.n554 B.n61 163.367
R1035 B.n99 B.n98 163.367
R1036 B.n103 B.n102 163.367
R1037 B.n107 B.n106 163.367
R1038 B.n111 B.n110 163.367
R1039 B.n115 B.n114 163.367
R1040 B.n119 B.n118 163.367
R1041 B.n123 B.n122 163.367
R1042 B.n127 B.n126 163.367
R1043 B.n131 B.n130 163.367
R1044 B.n135 B.n134 163.367
R1045 B.n139 B.n138 163.367
R1046 B.n143 B.n142 163.367
R1047 B.n147 B.n146 163.367
R1048 B.n151 B.n150 163.367
R1049 B.n155 B.n154 163.367
R1050 B.n159 B.n158 163.367
R1051 B.n163 B.n162 163.367
R1052 B.n167 B.n166 163.367
R1053 B.n171 B.n170 163.367
R1054 B.n175 B.n174 163.367
R1055 B.n179 B.n178 163.367
R1056 B.n183 B.n182 163.367
R1057 B.n187 B.n186 163.367
R1058 B.n191 B.n190 163.367
R1059 B.n195 B.n194 163.367
R1060 B.n199 B.n198 163.367
R1061 B.n203 B.n202 163.367
R1062 B.n205 B.n90 163.367
R1063 B.n421 B.n270 132.718
R1064 B.n561 B.n560 132.718
R1065 B.n303 B.n269 71.676
R1066 B.n307 B.n306 71.676
R1067 B.n312 B.n311 71.676
R1068 B.n315 B.n314 71.676
R1069 B.n320 B.n319 71.676
R1070 B.n323 B.n322 71.676
R1071 B.n328 B.n327 71.676
R1072 B.n331 B.n330 71.676
R1073 B.n336 B.n335 71.676
R1074 B.n339 B.n338 71.676
R1075 B.n344 B.n343 71.676
R1076 B.n347 B.n346 71.676
R1077 B.n353 B.n352 71.676
R1078 B.n356 B.n355 71.676
R1079 B.n361 B.n360 71.676
R1080 B.n364 B.n363 71.676
R1081 B.n372 B.n371 71.676
R1082 B.n375 B.n374 71.676
R1083 B.n380 B.n379 71.676
R1084 B.n383 B.n382 71.676
R1085 B.n388 B.n387 71.676
R1086 B.n391 B.n390 71.676
R1087 B.n396 B.n395 71.676
R1088 B.n399 B.n398 71.676
R1089 B.n404 B.n403 71.676
R1090 B.n407 B.n406 71.676
R1091 B.n412 B.n411 71.676
R1092 B.n415 B.n414 71.676
R1093 B.n62 B.n60 71.676
R1094 B.n99 B.n63 71.676
R1095 B.n103 B.n64 71.676
R1096 B.n107 B.n65 71.676
R1097 B.n111 B.n66 71.676
R1098 B.n115 B.n67 71.676
R1099 B.n119 B.n68 71.676
R1100 B.n123 B.n69 71.676
R1101 B.n127 B.n70 71.676
R1102 B.n131 B.n71 71.676
R1103 B.n135 B.n72 71.676
R1104 B.n139 B.n73 71.676
R1105 B.n143 B.n74 71.676
R1106 B.n147 B.n75 71.676
R1107 B.n151 B.n76 71.676
R1108 B.n155 B.n77 71.676
R1109 B.n159 B.n78 71.676
R1110 B.n163 B.n79 71.676
R1111 B.n167 B.n80 71.676
R1112 B.n171 B.n81 71.676
R1113 B.n175 B.n82 71.676
R1114 B.n179 B.n83 71.676
R1115 B.n183 B.n84 71.676
R1116 B.n187 B.n85 71.676
R1117 B.n191 B.n86 71.676
R1118 B.n195 B.n87 71.676
R1119 B.n199 B.n88 71.676
R1120 B.n203 B.n89 71.676
R1121 B.n559 B.n90 71.676
R1122 B.n559 B.n558 71.676
R1123 B.n205 B.n89 71.676
R1124 B.n202 B.n88 71.676
R1125 B.n198 B.n87 71.676
R1126 B.n194 B.n86 71.676
R1127 B.n190 B.n85 71.676
R1128 B.n186 B.n84 71.676
R1129 B.n182 B.n83 71.676
R1130 B.n178 B.n82 71.676
R1131 B.n174 B.n81 71.676
R1132 B.n170 B.n80 71.676
R1133 B.n166 B.n79 71.676
R1134 B.n162 B.n78 71.676
R1135 B.n158 B.n77 71.676
R1136 B.n154 B.n76 71.676
R1137 B.n150 B.n75 71.676
R1138 B.n146 B.n74 71.676
R1139 B.n142 B.n73 71.676
R1140 B.n138 B.n72 71.676
R1141 B.n134 B.n71 71.676
R1142 B.n130 B.n70 71.676
R1143 B.n126 B.n69 71.676
R1144 B.n122 B.n68 71.676
R1145 B.n118 B.n67 71.676
R1146 B.n114 B.n66 71.676
R1147 B.n110 B.n65 71.676
R1148 B.n106 B.n64 71.676
R1149 B.n102 B.n63 71.676
R1150 B.n98 B.n62 71.676
R1151 B.n304 B.n303 71.676
R1152 B.n306 B.n300 71.676
R1153 B.n313 B.n312 71.676
R1154 B.n314 B.n298 71.676
R1155 B.n321 B.n320 71.676
R1156 B.n322 B.n296 71.676
R1157 B.n329 B.n328 71.676
R1158 B.n330 B.n294 71.676
R1159 B.n337 B.n336 71.676
R1160 B.n338 B.n292 71.676
R1161 B.n345 B.n344 71.676
R1162 B.n346 B.n288 71.676
R1163 B.n354 B.n353 71.676
R1164 B.n355 B.n286 71.676
R1165 B.n362 B.n361 71.676
R1166 B.n363 B.n284 71.676
R1167 B.n373 B.n372 71.676
R1168 B.n374 B.n282 71.676
R1169 B.n381 B.n380 71.676
R1170 B.n382 B.n280 71.676
R1171 B.n389 B.n388 71.676
R1172 B.n390 B.n278 71.676
R1173 B.n397 B.n396 71.676
R1174 B.n398 B.n276 71.676
R1175 B.n405 B.n404 71.676
R1176 B.n406 B.n274 71.676
R1177 B.n413 B.n412 71.676
R1178 B.n416 B.n415 71.676
R1179 B.n421 B.n266 65.8746
R1180 B.n427 B.n266 65.8746
R1181 B.n427 B.n262 65.8746
R1182 B.n433 B.n262 65.8746
R1183 B.n433 B.n257 65.8746
R1184 B.n439 B.n257 65.8746
R1185 B.n439 B.n258 65.8746
R1186 B.n445 B.n250 65.8746
R1187 B.n451 B.n250 65.8746
R1188 B.n451 B.n246 65.8746
R1189 B.n457 B.n246 65.8746
R1190 B.n457 B.n242 65.8746
R1191 B.n463 B.n242 65.8746
R1192 B.n463 B.n238 65.8746
R1193 B.n469 B.n238 65.8746
R1194 B.n469 B.n234 65.8746
R1195 B.n475 B.n234 65.8746
R1196 B.n481 B.n230 65.8746
R1197 B.n481 B.n226 65.8746
R1198 B.n487 B.n226 65.8746
R1199 B.n487 B.n222 65.8746
R1200 B.n493 B.n222 65.8746
R1201 B.n493 B.n218 65.8746
R1202 B.n499 B.n218 65.8746
R1203 B.n506 B.n214 65.8746
R1204 B.n506 B.n210 65.8746
R1205 B.n512 B.n210 65.8746
R1206 B.n512 B.n4 65.8746
R1207 B.n625 B.n4 65.8746
R1208 B.n625 B.n624 65.8746
R1209 B.n624 B.n623 65.8746
R1210 B.n623 B.n8 65.8746
R1211 B.n617 B.n8 65.8746
R1212 B.n617 B.n616 65.8746
R1213 B.n615 B.n15 65.8746
R1214 B.n609 B.n15 65.8746
R1215 B.n609 B.n608 65.8746
R1216 B.n608 B.n607 65.8746
R1217 B.n607 B.n22 65.8746
R1218 B.n601 B.n22 65.8746
R1219 B.n601 B.n600 65.8746
R1220 B.n599 B.n29 65.8746
R1221 B.n593 B.n29 65.8746
R1222 B.n593 B.n592 65.8746
R1223 B.n592 B.n591 65.8746
R1224 B.n591 B.n36 65.8746
R1225 B.n585 B.n36 65.8746
R1226 B.n585 B.n584 65.8746
R1227 B.n584 B.n583 65.8746
R1228 B.n583 B.n43 65.8746
R1229 B.n577 B.n43 65.8746
R1230 B.n576 B.n575 65.8746
R1231 B.n575 B.n50 65.8746
R1232 B.n569 B.n50 65.8746
R1233 B.n569 B.n568 65.8746
R1234 B.n568 B.n567 65.8746
R1235 B.n567 B.n57 65.8746
R1236 B.n561 B.n57 65.8746
R1237 B.n369 B.n368 59.5399
R1238 B.n349 B.n290 59.5399
R1239 B.n96 B.n95 59.5399
R1240 B.n93 B.n92 59.5399
R1241 B.n445 B.t5 58.1247
R1242 B.n577 B.t12 58.1247
R1243 B.n368 B.n367 52.946
R1244 B.n290 B.n289 52.946
R1245 B.n95 B.n94 52.946
R1246 B.n92 B.n91 52.946
R1247 B.t3 B.n230 42.6249
R1248 B.n600 B.t2 42.6249
R1249 B.t0 B.n214 40.6874
R1250 B.n616 B.t1 40.6874
R1251 B.n563 B.n59 34.4981
R1252 B.n557 B.n556 34.4981
R1253 B.n419 B.n418 34.4981
R1254 B.n423 B.n268 34.4981
R1255 B.n499 B.t0 25.1876
R1256 B.t1 B.n615 25.1876
R1257 B.n475 B.t3 23.2502
R1258 B.t2 B.n599 23.2502
R1259 B B.n627 18.0485
R1260 B.n97 B.n59 10.6151
R1261 B.n100 B.n97 10.6151
R1262 B.n101 B.n100 10.6151
R1263 B.n104 B.n101 10.6151
R1264 B.n105 B.n104 10.6151
R1265 B.n108 B.n105 10.6151
R1266 B.n109 B.n108 10.6151
R1267 B.n112 B.n109 10.6151
R1268 B.n113 B.n112 10.6151
R1269 B.n116 B.n113 10.6151
R1270 B.n117 B.n116 10.6151
R1271 B.n120 B.n117 10.6151
R1272 B.n121 B.n120 10.6151
R1273 B.n124 B.n121 10.6151
R1274 B.n125 B.n124 10.6151
R1275 B.n128 B.n125 10.6151
R1276 B.n129 B.n128 10.6151
R1277 B.n132 B.n129 10.6151
R1278 B.n133 B.n132 10.6151
R1279 B.n136 B.n133 10.6151
R1280 B.n137 B.n136 10.6151
R1281 B.n140 B.n137 10.6151
R1282 B.n141 B.n140 10.6151
R1283 B.n145 B.n144 10.6151
R1284 B.n148 B.n145 10.6151
R1285 B.n149 B.n148 10.6151
R1286 B.n152 B.n149 10.6151
R1287 B.n153 B.n152 10.6151
R1288 B.n156 B.n153 10.6151
R1289 B.n157 B.n156 10.6151
R1290 B.n160 B.n157 10.6151
R1291 B.n161 B.n160 10.6151
R1292 B.n165 B.n164 10.6151
R1293 B.n168 B.n165 10.6151
R1294 B.n169 B.n168 10.6151
R1295 B.n172 B.n169 10.6151
R1296 B.n173 B.n172 10.6151
R1297 B.n176 B.n173 10.6151
R1298 B.n177 B.n176 10.6151
R1299 B.n180 B.n177 10.6151
R1300 B.n181 B.n180 10.6151
R1301 B.n184 B.n181 10.6151
R1302 B.n185 B.n184 10.6151
R1303 B.n188 B.n185 10.6151
R1304 B.n189 B.n188 10.6151
R1305 B.n192 B.n189 10.6151
R1306 B.n193 B.n192 10.6151
R1307 B.n196 B.n193 10.6151
R1308 B.n197 B.n196 10.6151
R1309 B.n200 B.n197 10.6151
R1310 B.n201 B.n200 10.6151
R1311 B.n204 B.n201 10.6151
R1312 B.n206 B.n204 10.6151
R1313 B.n207 B.n206 10.6151
R1314 B.n557 B.n207 10.6151
R1315 B.n419 B.n264 10.6151
R1316 B.n429 B.n264 10.6151
R1317 B.n430 B.n429 10.6151
R1318 B.n431 B.n430 10.6151
R1319 B.n431 B.n255 10.6151
R1320 B.n441 B.n255 10.6151
R1321 B.n442 B.n441 10.6151
R1322 B.n443 B.n442 10.6151
R1323 B.n443 B.n248 10.6151
R1324 B.n453 B.n248 10.6151
R1325 B.n454 B.n453 10.6151
R1326 B.n455 B.n454 10.6151
R1327 B.n455 B.n240 10.6151
R1328 B.n465 B.n240 10.6151
R1329 B.n466 B.n465 10.6151
R1330 B.n467 B.n466 10.6151
R1331 B.n467 B.n232 10.6151
R1332 B.n477 B.n232 10.6151
R1333 B.n478 B.n477 10.6151
R1334 B.n479 B.n478 10.6151
R1335 B.n479 B.n224 10.6151
R1336 B.n489 B.n224 10.6151
R1337 B.n490 B.n489 10.6151
R1338 B.n491 B.n490 10.6151
R1339 B.n491 B.n216 10.6151
R1340 B.n501 B.n216 10.6151
R1341 B.n502 B.n501 10.6151
R1342 B.n504 B.n502 10.6151
R1343 B.n504 B.n503 10.6151
R1344 B.n503 B.n208 10.6151
R1345 B.n515 B.n208 10.6151
R1346 B.n516 B.n515 10.6151
R1347 B.n517 B.n516 10.6151
R1348 B.n518 B.n517 10.6151
R1349 B.n520 B.n518 10.6151
R1350 B.n521 B.n520 10.6151
R1351 B.n522 B.n521 10.6151
R1352 B.n523 B.n522 10.6151
R1353 B.n525 B.n523 10.6151
R1354 B.n526 B.n525 10.6151
R1355 B.n527 B.n526 10.6151
R1356 B.n528 B.n527 10.6151
R1357 B.n530 B.n528 10.6151
R1358 B.n531 B.n530 10.6151
R1359 B.n532 B.n531 10.6151
R1360 B.n533 B.n532 10.6151
R1361 B.n535 B.n533 10.6151
R1362 B.n536 B.n535 10.6151
R1363 B.n537 B.n536 10.6151
R1364 B.n538 B.n537 10.6151
R1365 B.n540 B.n538 10.6151
R1366 B.n541 B.n540 10.6151
R1367 B.n542 B.n541 10.6151
R1368 B.n543 B.n542 10.6151
R1369 B.n545 B.n543 10.6151
R1370 B.n546 B.n545 10.6151
R1371 B.n547 B.n546 10.6151
R1372 B.n548 B.n547 10.6151
R1373 B.n550 B.n548 10.6151
R1374 B.n551 B.n550 10.6151
R1375 B.n552 B.n551 10.6151
R1376 B.n553 B.n552 10.6151
R1377 B.n555 B.n553 10.6151
R1378 B.n556 B.n555 10.6151
R1379 B.n302 B.n268 10.6151
R1380 B.n302 B.n301 10.6151
R1381 B.n308 B.n301 10.6151
R1382 B.n309 B.n308 10.6151
R1383 B.n310 B.n309 10.6151
R1384 B.n310 B.n299 10.6151
R1385 B.n316 B.n299 10.6151
R1386 B.n317 B.n316 10.6151
R1387 B.n318 B.n317 10.6151
R1388 B.n318 B.n297 10.6151
R1389 B.n324 B.n297 10.6151
R1390 B.n325 B.n324 10.6151
R1391 B.n326 B.n325 10.6151
R1392 B.n326 B.n295 10.6151
R1393 B.n332 B.n295 10.6151
R1394 B.n333 B.n332 10.6151
R1395 B.n334 B.n333 10.6151
R1396 B.n334 B.n293 10.6151
R1397 B.n340 B.n293 10.6151
R1398 B.n341 B.n340 10.6151
R1399 B.n342 B.n341 10.6151
R1400 B.n342 B.n291 10.6151
R1401 B.n348 B.n291 10.6151
R1402 B.n351 B.n350 10.6151
R1403 B.n351 B.n287 10.6151
R1404 B.n357 B.n287 10.6151
R1405 B.n358 B.n357 10.6151
R1406 B.n359 B.n358 10.6151
R1407 B.n359 B.n285 10.6151
R1408 B.n365 B.n285 10.6151
R1409 B.n366 B.n365 10.6151
R1410 B.n370 B.n366 10.6151
R1411 B.n376 B.n283 10.6151
R1412 B.n377 B.n376 10.6151
R1413 B.n378 B.n377 10.6151
R1414 B.n378 B.n281 10.6151
R1415 B.n384 B.n281 10.6151
R1416 B.n385 B.n384 10.6151
R1417 B.n386 B.n385 10.6151
R1418 B.n386 B.n279 10.6151
R1419 B.n392 B.n279 10.6151
R1420 B.n393 B.n392 10.6151
R1421 B.n394 B.n393 10.6151
R1422 B.n394 B.n277 10.6151
R1423 B.n400 B.n277 10.6151
R1424 B.n401 B.n400 10.6151
R1425 B.n402 B.n401 10.6151
R1426 B.n402 B.n275 10.6151
R1427 B.n408 B.n275 10.6151
R1428 B.n409 B.n408 10.6151
R1429 B.n410 B.n409 10.6151
R1430 B.n410 B.n273 10.6151
R1431 B.n273 B.n272 10.6151
R1432 B.n417 B.n272 10.6151
R1433 B.n418 B.n417 10.6151
R1434 B.n424 B.n423 10.6151
R1435 B.n425 B.n424 10.6151
R1436 B.n425 B.n260 10.6151
R1437 B.n435 B.n260 10.6151
R1438 B.n436 B.n435 10.6151
R1439 B.n437 B.n436 10.6151
R1440 B.n437 B.n252 10.6151
R1441 B.n447 B.n252 10.6151
R1442 B.n448 B.n447 10.6151
R1443 B.n449 B.n448 10.6151
R1444 B.n449 B.n244 10.6151
R1445 B.n459 B.n244 10.6151
R1446 B.n460 B.n459 10.6151
R1447 B.n461 B.n460 10.6151
R1448 B.n461 B.n236 10.6151
R1449 B.n471 B.n236 10.6151
R1450 B.n472 B.n471 10.6151
R1451 B.n473 B.n472 10.6151
R1452 B.n473 B.n228 10.6151
R1453 B.n483 B.n228 10.6151
R1454 B.n484 B.n483 10.6151
R1455 B.n485 B.n484 10.6151
R1456 B.n485 B.n220 10.6151
R1457 B.n495 B.n220 10.6151
R1458 B.n496 B.n495 10.6151
R1459 B.n497 B.n496 10.6151
R1460 B.n497 B.n212 10.6151
R1461 B.n508 B.n212 10.6151
R1462 B.n509 B.n508 10.6151
R1463 B.n510 B.n509 10.6151
R1464 B.n510 B.n0 10.6151
R1465 B.n621 B.n1 10.6151
R1466 B.n621 B.n620 10.6151
R1467 B.n620 B.n619 10.6151
R1468 B.n619 B.n10 10.6151
R1469 B.n613 B.n10 10.6151
R1470 B.n613 B.n612 10.6151
R1471 B.n612 B.n611 10.6151
R1472 B.n611 B.n17 10.6151
R1473 B.n605 B.n17 10.6151
R1474 B.n605 B.n604 10.6151
R1475 B.n604 B.n603 10.6151
R1476 B.n603 B.n24 10.6151
R1477 B.n597 B.n24 10.6151
R1478 B.n597 B.n596 10.6151
R1479 B.n596 B.n595 10.6151
R1480 B.n595 B.n31 10.6151
R1481 B.n589 B.n31 10.6151
R1482 B.n589 B.n588 10.6151
R1483 B.n588 B.n587 10.6151
R1484 B.n587 B.n38 10.6151
R1485 B.n581 B.n38 10.6151
R1486 B.n581 B.n580 10.6151
R1487 B.n580 B.n579 10.6151
R1488 B.n579 B.n45 10.6151
R1489 B.n573 B.n45 10.6151
R1490 B.n573 B.n572 10.6151
R1491 B.n572 B.n571 10.6151
R1492 B.n571 B.n52 10.6151
R1493 B.n565 B.n52 10.6151
R1494 B.n565 B.n564 10.6151
R1495 B.n564 B.n563 10.6151
R1496 B.n141 B.n96 9.36635
R1497 B.n164 B.n93 9.36635
R1498 B.n349 B.n348 9.36635
R1499 B.n369 B.n283 9.36635
R1500 B.n258 B.t5 7.75039
R1501 B.t12 B.n576 7.75039
R1502 B.n627 B.n0 2.81026
R1503 B.n627 B.n1 2.81026
R1504 B.n144 B.n96 1.24928
R1505 B.n161 B.n93 1.24928
R1506 B.n350 B.n349 1.24928
R1507 B.n370 B.n369 1.24928
R1508 VN.n0 VN.t3 95.7152
R1509 VN.n1 VN.t2 95.7152
R1510 VN.n0 VN.t1 94.9745
R1511 VN.n1 VN.t0 94.9745
R1512 VN VN.n1 46.0848
R1513 VN VN.n0 4.71735
R1514 VDD2.n2 VDD2.n0 104.758
R1515 VDD2.n2 VDD2.n1 68.7422
R1516 VDD2.n1 VDD2.t3 3.25708
R1517 VDD2.n1 VDD2.t1 3.25708
R1518 VDD2.n0 VDD2.t0 3.25708
R1519 VDD2.n0 VDD2.t2 3.25708
R1520 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 2.7901f
C1 VDD1 VTAIL 3.92936f
C2 VTAIL VDD2 3.98222f
C3 VN VP 4.95144f
C4 VDD1 VN 0.149285f
C5 VN VDD2 2.52575f
C6 VDD1 VP 2.75782f
C7 VP VDD2 0.382044f
C8 VDD1 VDD2 0.984365f
C9 VTAIL VN 2.77599f
C10 VDD2 B 3.187393f
C11 VDD1 B 6.69249f
C12 VTAIL B 6.182472f
C13 VN B 9.77882f
C14 VP B 7.994839f
C15 VDD2.t0 B 0.131721f
C16 VDD2.t2 B 0.131721f
C17 VDD2.n0 B 1.54578f
C18 VDD2.t3 B 0.131721f
C19 VDD2.t1 B 0.131721f
C20 VDD2.n1 B 1.10086f
C21 VDD2.n2 B 3.11268f
C22 VN.t3 B 1.37438f
C23 VN.t1 B 1.36965f
C24 VN.n0 B 0.893161f
C25 VN.t2 B 1.37438f
C26 VN.t0 B 1.36965f
C27 VN.n1 B 2.23947f
C28 VDD1.t0 B 0.133691f
C29 VDD1.t3 B 0.133691f
C30 VDD1.n0 B 1.11771f
C31 VDD1.t2 B 0.133691f
C32 VDD1.t1 B 0.133691f
C33 VDD1.n1 B 1.59267f
C34 VTAIL.n0 B 0.02819f
C35 VTAIL.n1 B 0.019314f
C36 VTAIL.n2 B 0.010378f
C37 VTAIL.n3 B 0.024531f
C38 VTAIL.n4 B 0.010989f
C39 VTAIL.n5 B 0.019314f
C40 VTAIL.n6 B 0.010378f
C41 VTAIL.n7 B 0.024531f
C42 VTAIL.n8 B 0.010989f
C43 VTAIL.n9 B 0.083077f
C44 VTAIL.t1 B 0.040007f
C45 VTAIL.n10 B 0.018398f
C46 VTAIL.n11 B 0.01449f
C47 VTAIL.n12 B 0.010378f
C48 VTAIL.n13 B 0.466569f
C49 VTAIL.n14 B 0.019314f
C50 VTAIL.n15 B 0.010378f
C51 VTAIL.n16 B 0.010989f
C52 VTAIL.n17 B 0.024531f
C53 VTAIL.n18 B 0.024531f
C54 VTAIL.n19 B 0.010989f
C55 VTAIL.n20 B 0.010378f
C56 VTAIL.n21 B 0.019314f
C57 VTAIL.n22 B 0.019314f
C58 VTAIL.n23 B 0.010378f
C59 VTAIL.n24 B 0.010989f
C60 VTAIL.n25 B 0.024531f
C61 VTAIL.n26 B 0.054948f
C62 VTAIL.n27 B 0.010989f
C63 VTAIL.n28 B 0.010378f
C64 VTAIL.n29 B 0.046753f
C65 VTAIL.n30 B 0.030999f
C66 VTAIL.n31 B 0.123779f
C67 VTAIL.n32 B 0.02819f
C68 VTAIL.n33 B 0.019314f
C69 VTAIL.n34 B 0.010378f
C70 VTAIL.n35 B 0.024531f
C71 VTAIL.n36 B 0.010989f
C72 VTAIL.n37 B 0.019314f
C73 VTAIL.n38 B 0.010378f
C74 VTAIL.n39 B 0.024531f
C75 VTAIL.n40 B 0.010989f
C76 VTAIL.n41 B 0.083077f
C77 VTAIL.t3 B 0.040007f
C78 VTAIL.n42 B 0.018398f
C79 VTAIL.n43 B 0.01449f
C80 VTAIL.n44 B 0.010378f
C81 VTAIL.n45 B 0.466569f
C82 VTAIL.n46 B 0.019314f
C83 VTAIL.n47 B 0.010378f
C84 VTAIL.n48 B 0.010989f
C85 VTAIL.n49 B 0.024531f
C86 VTAIL.n50 B 0.024531f
C87 VTAIL.n51 B 0.010989f
C88 VTAIL.n52 B 0.010378f
C89 VTAIL.n53 B 0.019314f
C90 VTAIL.n54 B 0.019314f
C91 VTAIL.n55 B 0.010378f
C92 VTAIL.n56 B 0.010989f
C93 VTAIL.n57 B 0.024531f
C94 VTAIL.n58 B 0.054948f
C95 VTAIL.n59 B 0.010989f
C96 VTAIL.n60 B 0.010378f
C97 VTAIL.n61 B 0.046753f
C98 VTAIL.n62 B 0.030999f
C99 VTAIL.n63 B 0.193388f
C100 VTAIL.n64 B 0.02819f
C101 VTAIL.n65 B 0.019314f
C102 VTAIL.n66 B 0.010378f
C103 VTAIL.n67 B 0.024531f
C104 VTAIL.n68 B 0.010989f
C105 VTAIL.n69 B 0.019314f
C106 VTAIL.n70 B 0.010378f
C107 VTAIL.n71 B 0.024531f
C108 VTAIL.n72 B 0.010989f
C109 VTAIL.n73 B 0.083077f
C110 VTAIL.t4 B 0.040007f
C111 VTAIL.n74 B 0.018398f
C112 VTAIL.n75 B 0.01449f
C113 VTAIL.n76 B 0.010378f
C114 VTAIL.n77 B 0.466569f
C115 VTAIL.n78 B 0.019314f
C116 VTAIL.n79 B 0.010378f
C117 VTAIL.n80 B 0.010989f
C118 VTAIL.n81 B 0.024531f
C119 VTAIL.n82 B 0.024531f
C120 VTAIL.n83 B 0.010989f
C121 VTAIL.n84 B 0.010378f
C122 VTAIL.n85 B 0.019314f
C123 VTAIL.n86 B 0.019314f
C124 VTAIL.n87 B 0.010378f
C125 VTAIL.n88 B 0.010989f
C126 VTAIL.n89 B 0.024531f
C127 VTAIL.n90 B 0.054948f
C128 VTAIL.n91 B 0.010989f
C129 VTAIL.n92 B 0.010378f
C130 VTAIL.n93 B 0.046753f
C131 VTAIL.n94 B 0.030999f
C132 VTAIL.n95 B 0.899149f
C133 VTAIL.n96 B 0.02819f
C134 VTAIL.n97 B 0.019314f
C135 VTAIL.n98 B 0.010378f
C136 VTAIL.n99 B 0.024531f
C137 VTAIL.n100 B 0.010989f
C138 VTAIL.n101 B 0.019314f
C139 VTAIL.n102 B 0.010378f
C140 VTAIL.n103 B 0.024531f
C141 VTAIL.n104 B 0.010989f
C142 VTAIL.n105 B 0.083077f
C143 VTAIL.t7 B 0.040007f
C144 VTAIL.n106 B 0.018398f
C145 VTAIL.n107 B 0.01449f
C146 VTAIL.n108 B 0.010378f
C147 VTAIL.n109 B 0.466569f
C148 VTAIL.n110 B 0.019314f
C149 VTAIL.n111 B 0.010378f
C150 VTAIL.n112 B 0.010989f
C151 VTAIL.n113 B 0.024531f
C152 VTAIL.n114 B 0.024531f
C153 VTAIL.n115 B 0.010989f
C154 VTAIL.n116 B 0.010378f
C155 VTAIL.n117 B 0.019314f
C156 VTAIL.n118 B 0.019314f
C157 VTAIL.n119 B 0.010378f
C158 VTAIL.n120 B 0.010989f
C159 VTAIL.n121 B 0.024531f
C160 VTAIL.n122 B 0.054948f
C161 VTAIL.n123 B 0.010989f
C162 VTAIL.n124 B 0.010378f
C163 VTAIL.n125 B 0.046753f
C164 VTAIL.n126 B 0.030999f
C165 VTAIL.n127 B 0.89915f
C166 VTAIL.n128 B 0.02819f
C167 VTAIL.n129 B 0.019314f
C168 VTAIL.n130 B 0.010378f
C169 VTAIL.n131 B 0.024531f
C170 VTAIL.n132 B 0.010989f
C171 VTAIL.n133 B 0.019314f
C172 VTAIL.n134 B 0.010378f
C173 VTAIL.n135 B 0.024531f
C174 VTAIL.n136 B 0.010989f
C175 VTAIL.n137 B 0.083077f
C176 VTAIL.t0 B 0.040007f
C177 VTAIL.n138 B 0.018398f
C178 VTAIL.n139 B 0.01449f
C179 VTAIL.n140 B 0.010378f
C180 VTAIL.n141 B 0.466569f
C181 VTAIL.n142 B 0.019314f
C182 VTAIL.n143 B 0.010378f
C183 VTAIL.n144 B 0.010989f
C184 VTAIL.n145 B 0.024531f
C185 VTAIL.n146 B 0.024531f
C186 VTAIL.n147 B 0.010989f
C187 VTAIL.n148 B 0.010378f
C188 VTAIL.n149 B 0.019314f
C189 VTAIL.n150 B 0.019314f
C190 VTAIL.n151 B 0.010378f
C191 VTAIL.n152 B 0.010989f
C192 VTAIL.n153 B 0.024531f
C193 VTAIL.n154 B 0.054948f
C194 VTAIL.n155 B 0.010989f
C195 VTAIL.n156 B 0.010378f
C196 VTAIL.n157 B 0.046753f
C197 VTAIL.n158 B 0.030999f
C198 VTAIL.n159 B 0.193388f
C199 VTAIL.n160 B 0.02819f
C200 VTAIL.n161 B 0.019314f
C201 VTAIL.n162 B 0.010378f
C202 VTAIL.n163 B 0.024531f
C203 VTAIL.n164 B 0.010989f
C204 VTAIL.n165 B 0.019314f
C205 VTAIL.n166 B 0.010378f
C206 VTAIL.n167 B 0.024531f
C207 VTAIL.n168 B 0.010989f
C208 VTAIL.n169 B 0.083077f
C209 VTAIL.t6 B 0.040007f
C210 VTAIL.n170 B 0.018398f
C211 VTAIL.n171 B 0.01449f
C212 VTAIL.n172 B 0.010378f
C213 VTAIL.n173 B 0.466569f
C214 VTAIL.n174 B 0.019314f
C215 VTAIL.n175 B 0.010378f
C216 VTAIL.n176 B 0.010989f
C217 VTAIL.n177 B 0.024531f
C218 VTAIL.n178 B 0.024531f
C219 VTAIL.n179 B 0.010989f
C220 VTAIL.n180 B 0.010378f
C221 VTAIL.n181 B 0.019314f
C222 VTAIL.n182 B 0.019314f
C223 VTAIL.n183 B 0.010378f
C224 VTAIL.n184 B 0.010989f
C225 VTAIL.n185 B 0.024531f
C226 VTAIL.n186 B 0.054948f
C227 VTAIL.n187 B 0.010989f
C228 VTAIL.n188 B 0.010378f
C229 VTAIL.n189 B 0.046753f
C230 VTAIL.n190 B 0.030999f
C231 VTAIL.n191 B 0.193388f
C232 VTAIL.n192 B 0.02819f
C233 VTAIL.n193 B 0.019314f
C234 VTAIL.n194 B 0.010378f
C235 VTAIL.n195 B 0.024531f
C236 VTAIL.n196 B 0.010989f
C237 VTAIL.n197 B 0.019314f
C238 VTAIL.n198 B 0.010378f
C239 VTAIL.n199 B 0.024531f
C240 VTAIL.n200 B 0.010989f
C241 VTAIL.n201 B 0.083077f
C242 VTAIL.t5 B 0.040007f
C243 VTAIL.n202 B 0.018398f
C244 VTAIL.n203 B 0.01449f
C245 VTAIL.n204 B 0.010378f
C246 VTAIL.n205 B 0.466569f
C247 VTAIL.n206 B 0.019314f
C248 VTAIL.n207 B 0.010378f
C249 VTAIL.n208 B 0.010989f
C250 VTAIL.n209 B 0.024531f
C251 VTAIL.n210 B 0.024531f
C252 VTAIL.n211 B 0.010989f
C253 VTAIL.n212 B 0.010378f
C254 VTAIL.n213 B 0.019314f
C255 VTAIL.n214 B 0.019314f
C256 VTAIL.n215 B 0.010378f
C257 VTAIL.n216 B 0.010989f
C258 VTAIL.n217 B 0.024531f
C259 VTAIL.n218 B 0.054948f
C260 VTAIL.n219 B 0.010989f
C261 VTAIL.n220 B 0.010378f
C262 VTAIL.n221 B 0.046753f
C263 VTAIL.n222 B 0.030999f
C264 VTAIL.n223 B 0.89915f
C265 VTAIL.n224 B 0.02819f
C266 VTAIL.n225 B 0.019314f
C267 VTAIL.n226 B 0.010378f
C268 VTAIL.n227 B 0.024531f
C269 VTAIL.n228 B 0.010989f
C270 VTAIL.n229 B 0.019314f
C271 VTAIL.n230 B 0.010378f
C272 VTAIL.n231 B 0.024531f
C273 VTAIL.n232 B 0.010989f
C274 VTAIL.n233 B 0.083077f
C275 VTAIL.t2 B 0.040007f
C276 VTAIL.n234 B 0.018398f
C277 VTAIL.n235 B 0.01449f
C278 VTAIL.n236 B 0.010378f
C279 VTAIL.n237 B 0.466569f
C280 VTAIL.n238 B 0.019314f
C281 VTAIL.n239 B 0.010378f
C282 VTAIL.n240 B 0.010989f
C283 VTAIL.n241 B 0.024531f
C284 VTAIL.n242 B 0.024531f
C285 VTAIL.n243 B 0.010989f
C286 VTAIL.n244 B 0.010378f
C287 VTAIL.n245 B 0.019314f
C288 VTAIL.n246 B 0.019314f
C289 VTAIL.n247 B 0.010378f
C290 VTAIL.n248 B 0.010989f
C291 VTAIL.n249 B 0.024531f
C292 VTAIL.n250 B 0.054948f
C293 VTAIL.n251 B 0.010989f
C294 VTAIL.n252 B 0.010378f
C295 VTAIL.n253 B 0.046753f
C296 VTAIL.n254 B 0.030999f
C297 VTAIL.n255 B 0.822297f
C298 VP.n0 B 0.040622f
C299 VP.t2 B 1.19098f
C300 VP.n1 B 0.044792f
C301 VP.n2 B 0.030813f
C302 VP.t1 B 1.19098f
C303 VP.n3 B 0.535649f
C304 VP.t0 B 1.4153f
C305 VP.t3 B 1.42019f
C306 VP.n4 B 2.29777f
C307 VP.n5 B 1.45229f
C308 VP.n6 B 0.040622f
C309 VP.n7 B 0.03542f
C310 VP.n8 B 0.05714f
C311 VP.n9 B 0.044792f
C312 VP.n10 B 0.030813f
C313 VP.n11 B 0.030813f
C314 VP.n12 B 0.030813f
C315 VP.n13 B 0.05714f
C316 VP.n14 B 0.03542f
C317 VP.n15 B 0.535649f
C318 VP.n16 B 0.051015f
.ends

