* NGSPICE file created from diff_pair_sample_1747.ext - technology: sky130A

.subckt diff_pair_sample_1747 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=0 ps=0 w=7.96 l=0.28
X1 VDD2.t9 VN.t0 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=1.3134 ps=8.29 w=7.96 l=0.28
X2 VTAIL.t6 VP.t0 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X3 VTAIL.t2 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X4 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=0 ps=0 w=7.96 l=0.28
X5 VTAIL.t13 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X6 VTAIL.t3 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X7 VTAIL.t4 VP.t3 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X8 VTAIL.t8 VN.t2 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X9 VDD1.t5 VP.t4 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=3.1044 ps=16.7 w=7.96 l=0.28
X10 VDD1.t4 VP.t5 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=1.3134 ps=8.29 w=7.96 l=0.28
X11 VDD2.t6 VN.t3 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=0 ps=0 w=7.96 l=0.28
X13 VTAIL.t9 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X14 VDD2.t4 VN.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=1.3134 ps=8.29 w=7.96 l=0.28
X15 VDD1.t3 VP.t6 VTAIL.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X16 VDD2.t3 VN.t6 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=3.1044 ps=16.7 w=7.96 l=0.28
X17 VDD1.t2 VP.t7 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=1.3134 ps=8.29 w=7.96 l=0.28
X18 VDD1.t1 VP.t8 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=3.1044 ps=16.7 w=7.96 l=0.28
X19 VTAIL.t12 VN.t7 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X20 VDD2.t1 VN.t8 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X21 VDD2.t0 VN.t9 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=3.1044 ps=16.7 w=7.96 l=0.28
X22 VDD1.t0 VP.t9 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3134 pd=8.29 as=1.3134 ps=8.29 w=7.96 l=0.28
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1044 pd=16.7 as=0 ps=0 w=7.96 l=0.28
R0 B.n282 B.t14 904.264
R1 B.n280 B.t18 904.264
R2 B.n76 B.t10 904.264
R3 B.n74 B.t21 904.264
R4 B.n508 B.n507 585
R5 B.n509 B.n508 585
R6 B.n210 B.n72 585
R7 B.n209 B.n208 585
R8 B.n207 B.n206 585
R9 B.n205 B.n204 585
R10 B.n203 B.n202 585
R11 B.n201 B.n200 585
R12 B.n199 B.n198 585
R13 B.n197 B.n196 585
R14 B.n195 B.n194 585
R15 B.n193 B.n192 585
R16 B.n191 B.n190 585
R17 B.n189 B.n188 585
R18 B.n187 B.n186 585
R19 B.n185 B.n184 585
R20 B.n183 B.n182 585
R21 B.n181 B.n180 585
R22 B.n179 B.n178 585
R23 B.n177 B.n176 585
R24 B.n175 B.n174 585
R25 B.n173 B.n172 585
R26 B.n171 B.n170 585
R27 B.n169 B.n168 585
R28 B.n167 B.n166 585
R29 B.n165 B.n164 585
R30 B.n163 B.n162 585
R31 B.n161 B.n160 585
R32 B.n159 B.n158 585
R33 B.n157 B.n156 585
R34 B.n155 B.n154 585
R35 B.n152 B.n151 585
R36 B.n150 B.n149 585
R37 B.n148 B.n147 585
R38 B.n146 B.n145 585
R39 B.n144 B.n143 585
R40 B.n142 B.n141 585
R41 B.n140 B.n139 585
R42 B.n138 B.n137 585
R43 B.n136 B.n135 585
R44 B.n134 B.n133 585
R45 B.n132 B.n131 585
R46 B.n130 B.n129 585
R47 B.n128 B.n127 585
R48 B.n126 B.n125 585
R49 B.n124 B.n123 585
R50 B.n122 B.n121 585
R51 B.n120 B.n119 585
R52 B.n118 B.n117 585
R53 B.n116 B.n115 585
R54 B.n114 B.n113 585
R55 B.n112 B.n111 585
R56 B.n110 B.n109 585
R57 B.n108 B.n107 585
R58 B.n106 B.n105 585
R59 B.n104 B.n103 585
R60 B.n102 B.n101 585
R61 B.n100 B.n99 585
R62 B.n98 B.n97 585
R63 B.n96 B.n95 585
R64 B.n94 B.n93 585
R65 B.n92 B.n91 585
R66 B.n90 B.n89 585
R67 B.n88 B.n87 585
R68 B.n86 B.n85 585
R69 B.n84 B.n83 585
R70 B.n82 B.n81 585
R71 B.n80 B.n79 585
R72 B.n38 B.n37 585
R73 B.n512 B.n511 585
R74 B.n506 B.n73 585
R75 B.n73 B.n35 585
R76 B.n505 B.n34 585
R77 B.n516 B.n34 585
R78 B.n504 B.n33 585
R79 B.n517 B.n33 585
R80 B.n503 B.n32 585
R81 B.n518 B.n32 585
R82 B.n502 B.n501 585
R83 B.n501 B.n31 585
R84 B.n500 B.n27 585
R85 B.n524 B.n27 585
R86 B.n499 B.n26 585
R87 B.n525 B.n26 585
R88 B.n498 B.n25 585
R89 B.n526 B.n25 585
R90 B.n497 B.n496 585
R91 B.n496 B.n21 585
R92 B.n495 B.n20 585
R93 B.n532 B.n20 585
R94 B.n494 B.n19 585
R95 B.n533 B.n19 585
R96 B.n493 B.n18 585
R97 B.n534 B.n18 585
R98 B.n492 B.n491 585
R99 B.n491 B.n490 585
R100 B.n489 B.n14 585
R101 B.n540 B.n14 585
R102 B.n488 B.n13 585
R103 B.n541 B.n13 585
R104 B.n487 B.n12 585
R105 B.n542 B.n12 585
R106 B.n486 B.n485 585
R107 B.n485 B.n11 585
R108 B.n484 B.n7 585
R109 B.n548 B.n7 585
R110 B.n483 B.n6 585
R111 B.n549 B.n6 585
R112 B.n482 B.n5 585
R113 B.n550 B.n5 585
R114 B.n481 B.n480 585
R115 B.n480 B.n4 585
R116 B.n479 B.n211 585
R117 B.n479 B.n478 585
R118 B.n468 B.n212 585
R119 B.n471 B.n212 585
R120 B.n470 B.n469 585
R121 B.n472 B.n470 585
R122 B.n467 B.n216 585
R123 B.n219 B.n216 585
R124 B.n466 B.n465 585
R125 B.n465 B.n464 585
R126 B.n218 B.n217 585
R127 B.n457 B.n218 585
R128 B.n456 B.n455 585
R129 B.n458 B.n456 585
R130 B.n454 B.n224 585
R131 B.n224 B.n223 585
R132 B.n453 B.n452 585
R133 B.n452 B.n451 585
R134 B.n226 B.n225 585
R135 B.n227 B.n226 585
R136 B.n444 B.n443 585
R137 B.n445 B.n444 585
R138 B.n442 B.n232 585
R139 B.n232 B.n231 585
R140 B.n441 B.n440 585
R141 B.n440 B.n439 585
R142 B.n234 B.n233 585
R143 B.n432 B.n234 585
R144 B.n431 B.n430 585
R145 B.n433 B.n431 585
R146 B.n429 B.n239 585
R147 B.n239 B.n238 585
R148 B.n428 B.n427 585
R149 B.n427 B.n426 585
R150 B.n241 B.n240 585
R151 B.n242 B.n241 585
R152 B.n422 B.n421 585
R153 B.n245 B.n244 585
R154 B.n418 B.n417 585
R155 B.n419 B.n418 585
R156 B.n416 B.n279 585
R157 B.n415 B.n414 585
R158 B.n413 B.n412 585
R159 B.n411 B.n410 585
R160 B.n409 B.n408 585
R161 B.n407 B.n406 585
R162 B.n405 B.n404 585
R163 B.n403 B.n402 585
R164 B.n401 B.n400 585
R165 B.n399 B.n398 585
R166 B.n397 B.n396 585
R167 B.n395 B.n394 585
R168 B.n393 B.n392 585
R169 B.n391 B.n390 585
R170 B.n389 B.n388 585
R171 B.n387 B.n386 585
R172 B.n385 B.n384 585
R173 B.n383 B.n382 585
R174 B.n381 B.n380 585
R175 B.n379 B.n378 585
R176 B.n377 B.n376 585
R177 B.n375 B.n374 585
R178 B.n373 B.n372 585
R179 B.n371 B.n370 585
R180 B.n369 B.n368 585
R181 B.n367 B.n366 585
R182 B.n365 B.n364 585
R183 B.n362 B.n361 585
R184 B.n360 B.n359 585
R185 B.n358 B.n357 585
R186 B.n356 B.n355 585
R187 B.n354 B.n353 585
R188 B.n352 B.n351 585
R189 B.n350 B.n349 585
R190 B.n348 B.n347 585
R191 B.n346 B.n345 585
R192 B.n344 B.n343 585
R193 B.n342 B.n341 585
R194 B.n340 B.n339 585
R195 B.n338 B.n337 585
R196 B.n336 B.n335 585
R197 B.n334 B.n333 585
R198 B.n332 B.n331 585
R199 B.n330 B.n329 585
R200 B.n328 B.n327 585
R201 B.n326 B.n325 585
R202 B.n324 B.n323 585
R203 B.n322 B.n321 585
R204 B.n320 B.n319 585
R205 B.n318 B.n317 585
R206 B.n316 B.n315 585
R207 B.n314 B.n313 585
R208 B.n312 B.n311 585
R209 B.n310 B.n309 585
R210 B.n308 B.n307 585
R211 B.n306 B.n305 585
R212 B.n304 B.n303 585
R213 B.n302 B.n301 585
R214 B.n300 B.n299 585
R215 B.n298 B.n297 585
R216 B.n296 B.n295 585
R217 B.n294 B.n293 585
R218 B.n292 B.n291 585
R219 B.n290 B.n289 585
R220 B.n288 B.n287 585
R221 B.n286 B.n285 585
R222 B.n423 B.n243 585
R223 B.n243 B.n242 585
R224 B.n425 B.n424 585
R225 B.n426 B.n425 585
R226 B.n237 B.n236 585
R227 B.n238 B.n237 585
R228 B.n435 B.n434 585
R229 B.n434 B.n433 585
R230 B.n436 B.n235 585
R231 B.n432 B.n235 585
R232 B.n438 B.n437 585
R233 B.n439 B.n438 585
R234 B.n230 B.n229 585
R235 B.n231 B.n230 585
R236 B.n447 B.n446 585
R237 B.n446 B.n445 585
R238 B.n448 B.n228 585
R239 B.n228 B.n227 585
R240 B.n450 B.n449 585
R241 B.n451 B.n450 585
R242 B.n222 B.n221 585
R243 B.n223 B.n222 585
R244 B.n460 B.n459 585
R245 B.n459 B.n458 585
R246 B.n461 B.n220 585
R247 B.n457 B.n220 585
R248 B.n463 B.n462 585
R249 B.n464 B.n463 585
R250 B.n215 B.n214 585
R251 B.n219 B.n215 585
R252 B.n474 B.n473 585
R253 B.n473 B.n472 585
R254 B.n475 B.n213 585
R255 B.n471 B.n213 585
R256 B.n477 B.n476 585
R257 B.n478 B.n477 585
R258 B.n2 B.n0 585
R259 B.n4 B.n2 585
R260 B.n3 B.n1 585
R261 B.n549 B.n3 585
R262 B.n547 B.n546 585
R263 B.n548 B.n547 585
R264 B.n545 B.n8 585
R265 B.n11 B.n8 585
R266 B.n544 B.n543 585
R267 B.n543 B.n542 585
R268 B.n10 B.n9 585
R269 B.n541 B.n10 585
R270 B.n539 B.n538 585
R271 B.n540 B.n539 585
R272 B.n537 B.n15 585
R273 B.n490 B.n15 585
R274 B.n536 B.n535 585
R275 B.n535 B.n534 585
R276 B.n17 B.n16 585
R277 B.n533 B.n17 585
R278 B.n531 B.n530 585
R279 B.n532 B.n531 585
R280 B.n529 B.n22 585
R281 B.n22 B.n21 585
R282 B.n528 B.n527 585
R283 B.n527 B.n526 585
R284 B.n24 B.n23 585
R285 B.n525 B.n24 585
R286 B.n523 B.n522 585
R287 B.n524 B.n523 585
R288 B.n521 B.n28 585
R289 B.n31 B.n28 585
R290 B.n520 B.n519 585
R291 B.n519 B.n518 585
R292 B.n30 B.n29 585
R293 B.n517 B.n30 585
R294 B.n515 B.n514 585
R295 B.n516 B.n515 585
R296 B.n513 B.n36 585
R297 B.n36 B.n35 585
R298 B.n552 B.n551 585
R299 B.n551 B.n550 585
R300 B.n421 B.n243 482.89
R301 B.n511 B.n36 482.89
R302 B.n285 B.n241 482.89
R303 B.n508 B.n73 482.89
R304 B.n509 B.n71 256.663
R305 B.n509 B.n70 256.663
R306 B.n509 B.n69 256.663
R307 B.n509 B.n68 256.663
R308 B.n509 B.n67 256.663
R309 B.n509 B.n66 256.663
R310 B.n509 B.n65 256.663
R311 B.n509 B.n64 256.663
R312 B.n509 B.n63 256.663
R313 B.n509 B.n62 256.663
R314 B.n509 B.n61 256.663
R315 B.n509 B.n60 256.663
R316 B.n509 B.n59 256.663
R317 B.n509 B.n58 256.663
R318 B.n509 B.n57 256.663
R319 B.n509 B.n56 256.663
R320 B.n509 B.n55 256.663
R321 B.n509 B.n54 256.663
R322 B.n509 B.n53 256.663
R323 B.n509 B.n52 256.663
R324 B.n509 B.n51 256.663
R325 B.n509 B.n50 256.663
R326 B.n509 B.n49 256.663
R327 B.n509 B.n48 256.663
R328 B.n509 B.n47 256.663
R329 B.n509 B.n46 256.663
R330 B.n509 B.n45 256.663
R331 B.n509 B.n44 256.663
R332 B.n509 B.n43 256.663
R333 B.n509 B.n42 256.663
R334 B.n509 B.n41 256.663
R335 B.n509 B.n40 256.663
R336 B.n509 B.n39 256.663
R337 B.n510 B.n509 256.663
R338 B.n420 B.n419 256.663
R339 B.n419 B.n246 256.663
R340 B.n419 B.n247 256.663
R341 B.n419 B.n248 256.663
R342 B.n419 B.n249 256.663
R343 B.n419 B.n250 256.663
R344 B.n419 B.n251 256.663
R345 B.n419 B.n252 256.663
R346 B.n419 B.n253 256.663
R347 B.n419 B.n254 256.663
R348 B.n419 B.n255 256.663
R349 B.n419 B.n256 256.663
R350 B.n419 B.n257 256.663
R351 B.n419 B.n258 256.663
R352 B.n419 B.n259 256.663
R353 B.n419 B.n260 256.663
R354 B.n419 B.n261 256.663
R355 B.n419 B.n262 256.663
R356 B.n419 B.n263 256.663
R357 B.n419 B.n264 256.663
R358 B.n419 B.n265 256.663
R359 B.n419 B.n266 256.663
R360 B.n419 B.n267 256.663
R361 B.n419 B.n268 256.663
R362 B.n419 B.n269 256.663
R363 B.n419 B.n270 256.663
R364 B.n419 B.n271 256.663
R365 B.n419 B.n272 256.663
R366 B.n419 B.n273 256.663
R367 B.n419 B.n274 256.663
R368 B.n419 B.n275 256.663
R369 B.n419 B.n276 256.663
R370 B.n419 B.n277 256.663
R371 B.n419 B.n278 256.663
R372 B.n282 B.t17 224.345
R373 B.n74 B.t22 224.345
R374 B.n280 B.t20 224.345
R375 B.n76 B.t12 224.345
R376 B.n283 B.t16 212.516
R377 B.n75 B.t23 212.516
R378 B.n281 B.t19 212.516
R379 B.n77 B.t13 212.516
R380 B.n425 B.n243 163.367
R381 B.n425 B.n237 163.367
R382 B.n434 B.n237 163.367
R383 B.n434 B.n235 163.367
R384 B.n438 B.n235 163.367
R385 B.n438 B.n230 163.367
R386 B.n446 B.n230 163.367
R387 B.n446 B.n228 163.367
R388 B.n450 B.n228 163.367
R389 B.n450 B.n222 163.367
R390 B.n459 B.n222 163.367
R391 B.n459 B.n220 163.367
R392 B.n463 B.n220 163.367
R393 B.n463 B.n215 163.367
R394 B.n473 B.n215 163.367
R395 B.n473 B.n213 163.367
R396 B.n477 B.n213 163.367
R397 B.n477 B.n2 163.367
R398 B.n551 B.n2 163.367
R399 B.n551 B.n3 163.367
R400 B.n547 B.n3 163.367
R401 B.n547 B.n8 163.367
R402 B.n543 B.n8 163.367
R403 B.n543 B.n10 163.367
R404 B.n539 B.n10 163.367
R405 B.n539 B.n15 163.367
R406 B.n535 B.n15 163.367
R407 B.n535 B.n17 163.367
R408 B.n531 B.n17 163.367
R409 B.n531 B.n22 163.367
R410 B.n527 B.n22 163.367
R411 B.n527 B.n24 163.367
R412 B.n523 B.n24 163.367
R413 B.n523 B.n28 163.367
R414 B.n519 B.n28 163.367
R415 B.n519 B.n30 163.367
R416 B.n515 B.n30 163.367
R417 B.n515 B.n36 163.367
R418 B.n418 B.n245 163.367
R419 B.n418 B.n279 163.367
R420 B.n414 B.n413 163.367
R421 B.n410 B.n409 163.367
R422 B.n406 B.n405 163.367
R423 B.n402 B.n401 163.367
R424 B.n398 B.n397 163.367
R425 B.n394 B.n393 163.367
R426 B.n390 B.n389 163.367
R427 B.n386 B.n385 163.367
R428 B.n382 B.n381 163.367
R429 B.n378 B.n377 163.367
R430 B.n374 B.n373 163.367
R431 B.n370 B.n369 163.367
R432 B.n366 B.n365 163.367
R433 B.n361 B.n360 163.367
R434 B.n357 B.n356 163.367
R435 B.n353 B.n352 163.367
R436 B.n349 B.n348 163.367
R437 B.n345 B.n344 163.367
R438 B.n341 B.n340 163.367
R439 B.n337 B.n336 163.367
R440 B.n333 B.n332 163.367
R441 B.n329 B.n328 163.367
R442 B.n325 B.n324 163.367
R443 B.n321 B.n320 163.367
R444 B.n317 B.n316 163.367
R445 B.n313 B.n312 163.367
R446 B.n309 B.n308 163.367
R447 B.n305 B.n304 163.367
R448 B.n301 B.n300 163.367
R449 B.n297 B.n296 163.367
R450 B.n293 B.n292 163.367
R451 B.n289 B.n288 163.367
R452 B.n427 B.n241 163.367
R453 B.n427 B.n239 163.367
R454 B.n431 B.n239 163.367
R455 B.n431 B.n234 163.367
R456 B.n440 B.n234 163.367
R457 B.n440 B.n232 163.367
R458 B.n444 B.n232 163.367
R459 B.n444 B.n226 163.367
R460 B.n452 B.n226 163.367
R461 B.n452 B.n224 163.367
R462 B.n456 B.n224 163.367
R463 B.n456 B.n218 163.367
R464 B.n465 B.n218 163.367
R465 B.n465 B.n216 163.367
R466 B.n470 B.n216 163.367
R467 B.n470 B.n212 163.367
R468 B.n479 B.n212 163.367
R469 B.n480 B.n479 163.367
R470 B.n480 B.n5 163.367
R471 B.n6 B.n5 163.367
R472 B.n7 B.n6 163.367
R473 B.n485 B.n7 163.367
R474 B.n485 B.n12 163.367
R475 B.n13 B.n12 163.367
R476 B.n14 B.n13 163.367
R477 B.n491 B.n14 163.367
R478 B.n491 B.n18 163.367
R479 B.n19 B.n18 163.367
R480 B.n20 B.n19 163.367
R481 B.n496 B.n20 163.367
R482 B.n496 B.n25 163.367
R483 B.n26 B.n25 163.367
R484 B.n27 B.n26 163.367
R485 B.n501 B.n27 163.367
R486 B.n501 B.n32 163.367
R487 B.n33 B.n32 163.367
R488 B.n34 B.n33 163.367
R489 B.n73 B.n34 163.367
R490 B.n79 B.n38 163.367
R491 B.n83 B.n82 163.367
R492 B.n87 B.n86 163.367
R493 B.n91 B.n90 163.367
R494 B.n95 B.n94 163.367
R495 B.n99 B.n98 163.367
R496 B.n103 B.n102 163.367
R497 B.n107 B.n106 163.367
R498 B.n111 B.n110 163.367
R499 B.n115 B.n114 163.367
R500 B.n119 B.n118 163.367
R501 B.n123 B.n122 163.367
R502 B.n127 B.n126 163.367
R503 B.n131 B.n130 163.367
R504 B.n135 B.n134 163.367
R505 B.n139 B.n138 163.367
R506 B.n143 B.n142 163.367
R507 B.n147 B.n146 163.367
R508 B.n151 B.n150 163.367
R509 B.n156 B.n155 163.367
R510 B.n160 B.n159 163.367
R511 B.n164 B.n163 163.367
R512 B.n168 B.n167 163.367
R513 B.n172 B.n171 163.367
R514 B.n176 B.n175 163.367
R515 B.n180 B.n179 163.367
R516 B.n184 B.n183 163.367
R517 B.n188 B.n187 163.367
R518 B.n192 B.n191 163.367
R519 B.n196 B.n195 163.367
R520 B.n200 B.n199 163.367
R521 B.n204 B.n203 163.367
R522 B.n208 B.n207 163.367
R523 B.n508 B.n72 163.367
R524 B.n419 B.n242 95.5804
R525 B.n509 B.n35 95.5804
R526 B.n421 B.n420 71.676
R527 B.n279 B.n246 71.676
R528 B.n413 B.n247 71.676
R529 B.n409 B.n248 71.676
R530 B.n405 B.n249 71.676
R531 B.n401 B.n250 71.676
R532 B.n397 B.n251 71.676
R533 B.n393 B.n252 71.676
R534 B.n389 B.n253 71.676
R535 B.n385 B.n254 71.676
R536 B.n381 B.n255 71.676
R537 B.n377 B.n256 71.676
R538 B.n373 B.n257 71.676
R539 B.n369 B.n258 71.676
R540 B.n365 B.n259 71.676
R541 B.n360 B.n260 71.676
R542 B.n356 B.n261 71.676
R543 B.n352 B.n262 71.676
R544 B.n348 B.n263 71.676
R545 B.n344 B.n264 71.676
R546 B.n340 B.n265 71.676
R547 B.n336 B.n266 71.676
R548 B.n332 B.n267 71.676
R549 B.n328 B.n268 71.676
R550 B.n324 B.n269 71.676
R551 B.n320 B.n270 71.676
R552 B.n316 B.n271 71.676
R553 B.n312 B.n272 71.676
R554 B.n308 B.n273 71.676
R555 B.n304 B.n274 71.676
R556 B.n300 B.n275 71.676
R557 B.n296 B.n276 71.676
R558 B.n292 B.n277 71.676
R559 B.n288 B.n278 71.676
R560 B.n511 B.n510 71.676
R561 B.n79 B.n39 71.676
R562 B.n83 B.n40 71.676
R563 B.n87 B.n41 71.676
R564 B.n91 B.n42 71.676
R565 B.n95 B.n43 71.676
R566 B.n99 B.n44 71.676
R567 B.n103 B.n45 71.676
R568 B.n107 B.n46 71.676
R569 B.n111 B.n47 71.676
R570 B.n115 B.n48 71.676
R571 B.n119 B.n49 71.676
R572 B.n123 B.n50 71.676
R573 B.n127 B.n51 71.676
R574 B.n131 B.n52 71.676
R575 B.n135 B.n53 71.676
R576 B.n139 B.n54 71.676
R577 B.n143 B.n55 71.676
R578 B.n147 B.n56 71.676
R579 B.n151 B.n57 71.676
R580 B.n156 B.n58 71.676
R581 B.n160 B.n59 71.676
R582 B.n164 B.n60 71.676
R583 B.n168 B.n61 71.676
R584 B.n172 B.n62 71.676
R585 B.n176 B.n63 71.676
R586 B.n180 B.n64 71.676
R587 B.n184 B.n65 71.676
R588 B.n188 B.n66 71.676
R589 B.n192 B.n67 71.676
R590 B.n196 B.n68 71.676
R591 B.n200 B.n69 71.676
R592 B.n204 B.n70 71.676
R593 B.n208 B.n71 71.676
R594 B.n72 B.n71 71.676
R595 B.n207 B.n70 71.676
R596 B.n203 B.n69 71.676
R597 B.n199 B.n68 71.676
R598 B.n195 B.n67 71.676
R599 B.n191 B.n66 71.676
R600 B.n187 B.n65 71.676
R601 B.n183 B.n64 71.676
R602 B.n179 B.n63 71.676
R603 B.n175 B.n62 71.676
R604 B.n171 B.n61 71.676
R605 B.n167 B.n60 71.676
R606 B.n163 B.n59 71.676
R607 B.n159 B.n58 71.676
R608 B.n155 B.n57 71.676
R609 B.n150 B.n56 71.676
R610 B.n146 B.n55 71.676
R611 B.n142 B.n54 71.676
R612 B.n138 B.n53 71.676
R613 B.n134 B.n52 71.676
R614 B.n130 B.n51 71.676
R615 B.n126 B.n50 71.676
R616 B.n122 B.n49 71.676
R617 B.n118 B.n48 71.676
R618 B.n114 B.n47 71.676
R619 B.n110 B.n46 71.676
R620 B.n106 B.n45 71.676
R621 B.n102 B.n44 71.676
R622 B.n98 B.n43 71.676
R623 B.n94 B.n42 71.676
R624 B.n90 B.n41 71.676
R625 B.n86 B.n40 71.676
R626 B.n82 B.n39 71.676
R627 B.n510 B.n38 71.676
R628 B.n420 B.n245 71.676
R629 B.n414 B.n246 71.676
R630 B.n410 B.n247 71.676
R631 B.n406 B.n248 71.676
R632 B.n402 B.n249 71.676
R633 B.n398 B.n250 71.676
R634 B.n394 B.n251 71.676
R635 B.n390 B.n252 71.676
R636 B.n386 B.n253 71.676
R637 B.n382 B.n254 71.676
R638 B.n378 B.n255 71.676
R639 B.n374 B.n256 71.676
R640 B.n370 B.n257 71.676
R641 B.n366 B.n258 71.676
R642 B.n361 B.n259 71.676
R643 B.n357 B.n260 71.676
R644 B.n353 B.n261 71.676
R645 B.n349 B.n262 71.676
R646 B.n345 B.n263 71.676
R647 B.n341 B.n264 71.676
R648 B.n337 B.n265 71.676
R649 B.n333 B.n266 71.676
R650 B.n329 B.n267 71.676
R651 B.n325 B.n268 71.676
R652 B.n321 B.n269 71.676
R653 B.n317 B.n270 71.676
R654 B.n313 B.n271 71.676
R655 B.n309 B.n272 71.676
R656 B.n305 B.n273 71.676
R657 B.n301 B.n274 71.676
R658 B.n297 B.n275 71.676
R659 B.n293 B.n276 71.676
R660 B.n289 B.n277 71.676
R661 B.n285 B.n278 71.676
R662 B.n284 B.n283 59.5399
R663 B.n363 B.n281 59.5399
R664 B.n78 B.n77 59.5399
R665 B.n153 B.n75 59.5399
R666 B.n426 B.n242 56.5173
R667 B.n426 B.n238 56.5173
R668 B.n433 B.n238 56.5173
R669 B.n433 B.n432 56.5173
R670 B.n439 B.n231 56.5173
R671 B.n445 B.n231 56.5173
R672 B.n445 B.n227 56.5173
R673 B.n451 B.n227 56.5173
R674 B.n458 B.n223 56.5173
R675 B.n464 B.n219 56.5173
R676 B.n472 B.n471 56.5173
R677 B.n478 B.n4 56.5173
R678 B.n550 B.n4 56.5173
R679 B.n550 B.n549 56.5173
R680 B.n549 B.n548 56.5173
R681 B.n542 B.n11 56.5173
R682 B.n541 B.n540 56.5173
R683 B.n534 B.n533 56.5173
R684 B.n532 B.n21 56.5173
R685 B.n526 B.n21 56.5173
R686 B.n526 B.n525 56.5173
R687 B.n525 B.n524 56.5173
R688 B.n518 B.n31 56.5173
R689 B.n518 B.n517 56.5173
R690 B.n517 B.n516 56.5173
R691 B.n516 B.n35 56.5173
R692 B.n457 B.t9 51.5305
R693 B.n490 B.t7 51.5305
R694 B.t4 B.n457 49.8683
R695 B.n490 B.t3 49.8683
R696 B.n219 B.t5 39.8947
R697 B.t0 B.n541 39.8947
R698 B.n439 B.t15 38.2325
R699 B.t6 B.n223 38.2325
R700 B.n533 B.t8 38.2325
R701 B.n524 B.t11 38.2325
R702 B.n513 B.n512 31.3761
R703 B.n507 B.n506 31.3761
R704 B.n286 B.n240 31.3761
R705 B.n423 B.n422 31.3761
R706 B.n471 B.t1 28.2589
R707 B.n478 B.t1 28.2589
R708 B.n548 B.t2 28.2589
R709 B.n11 B.t2 28.2589
R710 B.n432 B.t15 18.2854
R711 B.n451 B.t6 18.2854
R712 B.t8 B.n532 18.2854
R713 B.n31 B.t11 18.2854
R714 B B.n552 18.0485
R715 B.n472 B.t5 16.6231
R716 B.n542 B.t0 16.6231
R717 B.n283 B.n282 11.8308
R718 B.n281 B.n280 11.8308
R719 B.n77 B.n76 11.8308
R720 B.n75 B.n74 11.8308
R721 B.n512 B.n37 10.6151
R722 B.n80 B.n37 10.6151
R723 B.n81 B.n80 10.6151
R724 B.n84 B.n81 10.6151
R725 B.n85 B.n84 10.6151
R726 B.n88 B.n85 10.6151
R727 B.n89 B.n88 10.6151
R728 B.n92 B.n89 10.6151
R729 B.n93 B.n92 10.6151
R730 B.n96 B.n93 10.6151
R731 B.n97 B.n96 10.6151
R732 B.n100 B.n97 10.6151
R733 B.n101 B.n100 10.6151
R734 B.n104 B.n101 10.6151
R735 B.n105 B.n104 10.6151
R736 B.n108 B.n105 10.6151
R737 B.n109 B.n108 10.6151
R738 B.n112 B.n109 10.6151
R739 B.n113 B.n112 10.6151
R740 B.n116 B.n113 10.6151
R741 B.n117 B.n116 10.6151
R742 B.n120 B.n117 10.6151
R743 B.n121 B.n120 10.6151
R744 B.n124 B.n121 10.6151
R745 B.n125 B.n124 10.6151
R746 B.n128 B.n125 10.6151
R747 B.n129 B.n128 10.6151
R748 B.n132 B.n129 10.6151
R749 B.n133 B.n132 10.6151
R750 B.n137 B.n136 10.6151
R751 B.n140 B.n137 10.6151
R752 B.n141 B.n140 10.6151
R753 B.n144 B.n141 10.6151
R754 B.n145 B.n144 10.6151
R755 B.n148 B.n145 10.6151
R756 B.n149 B.n148 10.6151
R757 B.n152 B.n149 10.6151
R758 B.n157 B.n154 10.6151
R759 B.n158 B.n157 10.6151
R760 B.n161 B.n158 10.6151
R761 B.n162 B.n161 10.6151
R762 B.n165 B.n162 10.6151
R763 B.n166 B.n165 10.6151
R764 B.n169 B.n166 10.6151
R765 B.n170 B.n169 10.6151
R766 B.n173 B.n170 10.6151
R767 B.n174 B.n173 10.6151
R768 B.n177 B.n174 10.6151
R769 B.n178 B.n177 10.6151
R770 B.n181 B.n178 10.6151
R771 B.n182 B.n181 10.6151
R772 B.n185 B.n182 10.6151
R773 B.n186 B.n185 10.6151
R774 B.n189 B.n186 10.6151
R775 B.n190 B.n189 10.6151
R776 B.n193 B.n190 10.6151
R777 B.n194 B.n193 10.6151
R778 B.n197 B.n194 10.6151
R779 B.n198 B.n197 10.6151
R780 B.n201 B.n198 10.6151
R781 B.n202 B.n201 10.6151
R782 B.n205 B.n202 10.6151
R783 B.n206 B.n205 10.6151
R784 B.n209 B.n206 10.6151
R785 B.n210 B.n209 10.6151
R786 B.n507 B.n210 10.6151
R787 B.n428 B.n240 10.6151
R788 B.n429 B.n428 10.6151
R789 B.n430 B.n429 10.6151
R790 B.n430 B.n233 10.6151
R791 B.n441 B.n233 10.6151
R792 B.n442 B.n441 10.6151
R793 B.n443 B.n442 10.6151
R794 B.n443 B.n225 10.6151
R795 B.n453 B.n225 10.6151
R796 B.n454 B.n453 10.6151
R797 B.n455 B.n454 10.6151
R798 B.n455 B.n217 10.6151
R799 B.n466 B.n217 10.6151
R800 B.n467 B.n466 10.6151
R801 B.n469 B.n467 10.6151
R802 B.n469 B.n468 10.6151
R803 B.n468 B.n211 10.6151
R804 B.n481 B.n211 10.6151
R805 B.n482 B.n481 10.6151
R806 B.n483 B.n482 10.6151
R807 B.n484 B.n483 10.6151
R808 B.n486 B.n484 10.6151
R809 B.n487 B.n486 10.6151
R810 B.n488 B.n487 10.6151
R811 B.n489 B.n488 10.6151
R812 B.n492 B.n489 10.6151
R813 B.n493 B.n492 10.6151
R814 B.n494 B.n493 10.6151
R815 B.n495 B.n494 10.6151
R816 B.n497 B.n495 10.6151
R817 B.n498 B.n497 10.6151
R818 B.n499 B.n498 10.6151
R819 B.n500 B.n499 10.6151
R820 B.n502 B.n500 10.6151
R821 B.n503 B.n502 10.6151
R822 B.n504 B.n503 10.6151
R823 B.n505 B.n504 10.6151
R824 B.n506 B.n505 10.6151
R825 B.n422 B.n244 10.6151
R826 B.n417 B.n244 10.6151
R827 B.n417 B.n416 10.6151
R828 B.n416 B.n415 10.6151
R829 B.n415 B.n412 10.6151
R830 B.n412 B.n411 10.6151
R831 B.n411 B.n408 10.6151
R832 B.n408 B.n407 10.6151
R833 B.n407 B.n404 10.6151
R834 B.n404 B.n403 10.6151
R835 B.n403 B.n400 10.6151
R836 B.n400 B.n399 10.6151
R837 B.n399 B.n396 10.6151
R838 B.n396 B.n395 10.6151
R839 B.n395 B.n392 10.6151
R840 B.n392 B.n391 10.6151
R841 B.n391 B.n388 10.6151
R842 B.n388 B.n387 10.6151
R843 B.n387 B.n384 10.6151
R844 B.n384 B.n383 10.6151
R845 B.n383 B.n380 10.6151
R846 B.n380 B.n379 10.6151
R847 B.n379 B.n376 10.6151
R848 B.n376 B.n375 10.6151
R849 B.n375 B.n372 10.6151
R850 B.n372 B.n371 10.6151
R851 B.n371 B.n368 10.6151
R852 B.n368 B.n367 10.6151
R853 B.n367 B.n364 10.6151
R854 B.n362 B.n359 10.6151
R855 B.n359 B.n358 10.6151
R856 B.n358 B.n355 10.6151
R857 B.n355 B.n354 10.6151
R858 B.n354 B.n351 10.6151
R859 B.n351 B.n350 10.6151
R860 B.n350 B.n347 10.6151
R861 B.n347 B.n346 10.6151
R862 B.n343 B.n342 10.6151
R863 B.n342 B.n339 10.6151
R864 B.n339 B.n338 10.6151
R865 B.n338 B.n335 10.6151
R866 B.n335 B.n334 10.6151
R867 B.n334 B.n331 10.6151
R868 B.n331 B.n330 10.6151
R869 B.n330 B.n327 10.6151
R870 B.n327 B.n326 10.6151
R871 B.n326 B.n323 10.6151
R872 B.n323 B.n322 10.6151
R873 B.n322 B.n319 10.6151
R874 B.n319 B.n318 10.6151
R875 B.n318 B.n315 10.6151
R876 B.n315 B.n314 10.6151
R877 B.n314 B.n311 10.6151
R878 B.n311 B.n310 10.6151
R879 B.n310 B.n307 10.6151
R880 B.n307 B.n306 10.6151
R881 B.n306 B.n303 10.6151
R882 B.n303 B.n302 10.6151
R883 B.n302 B.n299 10.6151
R884 B.n299 B.n298 10.6151
R885 B.n298 B.n295 10.6151
R886 B.n295 B.n294 10.6151
R887 B.n294 B.n291 10.6151
R888 B.n291 B.n290 10.6151
R889 B.n290 B.n287 10.6151
R890 B.n287 B.n286 10.6151
R891 B.n424 B.n423 10.6151
R892 B.n424 B.n236 10.6151
R893 B.n435 B.n236 10.6151
R894 B.n436 B.n435 10.6151
R895 B.n437 B.n436 10.6151
R896 B.n437 B.n229 10.6151
R897 B.n447 B.n229 10.6151
R898 B.n448 B.n447 10.6151
R899 B.n449 B.n448 10.6151
R900 B.n449 B.n221 10.6151
R901 B.n460 B.n221 10.6151
R902 B.n461 B.n460 10.6151
R903 B.n462 B.n461 10.6151
R904 B.n462 B.n214 10.6151
R905 B.n474 B.n214 10.6151
R906 B.n475 B.n474 10.6151
R907 B.n476 B.n475 10.6151
R908 B.n476 B.n0 10.6151
R909 B.n546 B.n1 10.6151
R910 B.n546 B.n545 10.6151
R911 B.n545 B.n544 10.6151
R912 B.n544 B.n9 10.6151
R913 B.n538 B.n9 10.6151
R914 B.n538 B.n537 10.6151
R915 B.n537 B.n536 10.6151
R916 B.n536 B.n16 10.6151
R917 B.n530 B.n16 10.6151
R918 B.n530 B.n529 10.6151
R919 B.n529 B.n528 10.6151
R920 B.n528 B.n23 10.6151
R921 B.n522 B.n23 10.6151
R922 B.n522 B.n521 10.6151
R923 B.n521 B.n520 10.6151
R924 B.n520 B.n29 10.6151
R925 B.n514 B.n29 10.6151
R926 B.n514 B.n513 10.6151
R927 B.n458 B.t4 6.64954
R928 B.n534 B.t3 6.64954
R929 B.n136 B.n78 6.5566
R930 B.n153 B.n152 6.5566
R931 B.n363 B.n362 6.5566
R932 B.n346 B.n284 6.5566
R933 B.n464 B.t9 4.98728
R934 B.n540 B.t7 4.98728
R935 B.n133 B.n78 4.05904
R936 B.n154 B.n153 4.05904
R937 B.n364 B.n363 4.05904
R938 B.n343 B.n284 4.05904
R939 B.n552 B.n0 2.81026
R940 B.n552 B.n1 2.81026
R941 VN.n9 VN.t9 830.876
R942 VN.n3 VN.t5 830.876
R943 VN.n20 VN.t0 830.876
R944 VN.n14 VN.t6 830.876
R945 VN.n6 VN.t3 798.744
R946 VN.n8 VN.t1 798.744
R947 VN.n2 VN.t7 798.744
R948 VN.n17 VN.t8 798.744
R949 VN.n19 VN.t4 798.744
R950 VN.n13 VN.t2 798.744
R951 VN.n15 VN.n14 161.489
R952 VN.n4 VN.n3 161.489
R953 VN.n10 VN.n9 161.3
R954 VN.n21 VN.n20 161.3
R955 VN.n18 VN.n11 161.3
R956 VN.n17 VN.n16 161.3
R957 VN.n15 VN.n12 161.3
R958 VN.n7 VN.n0 161.3
R959 VN.n6 VN.n5 161.3
R960 VN.n4 VN.n1 161.3
R961 VN.n6 VN.n1 73.0308
R962 VN.n7 VN.n6 73.0308
R963 VN.n18 VN.n17 73.0308
R964 VN.n17 VN.n12 73.0308
R965 VN.n3 VN.n2 56.9641
R966 VN.n9 VN.n8 56.9641
R967 VN.n20 VN.n19 56.9641
R968 VN.n14 VN.n13 56.9641
R969 VN VN.n21 37.8395
R970 VN.n2 VN.n1 16.0672
R971 VN.n8 VN.n7 16.0672
R972 VN.n19 VN.n18 16.0672
R973 VN.n13 VN.n12 16.0672
R974 VN.n21 VN.n11 0.189894
R975 VN.n16 VN.n11 0.189894
R976 VN.n16 VN.n15 0.189894
R977 VN.n5 VN.n4 0.189894
R978 VN.n5 VN.n0 0.189894
R979 VN.n10 VN.n0 0.189894
R980 VN VN.n10 0.0516364
R981 VTAIL.n176 VTAIL.n140 289.615
R982 VTAIL.n38 VTAIL.n2 289.615
R983 VTAIL.n134 VTAIL.n98 289.615
R984 VTAIL.n88 VTAIL.n52 289.615
R985 VTAIL.n152 VTAIL.n151 185
R986 VTAIL.n157 VTAIL.n156 185
R987 VTAIL.n159 VTAIL.n158 185
R988 VTAIL.n148 VTAIL.n147 185
R989 VTAIL.n165 VTAIL.n164 185
R990 VTAIL.n167 VTAIL.n166 185
R991 VTAIL.n144 VTAIL.n143 185
R992 VTAIL.n174 VTAIL.n173 185
R993 VTAIL.n175 VTAIL.n142 185
R994 VTAIL.n177 VTAIL.n176 185
R995 VTAIL.n14 VTAIL.n13 185
R996 VTAIL.n19 VTAIL.n18 185
R997 VTAIL.n21 VTAIL.n20 185
R998 VTAIL.n10 VTAIL.n9 185
R999 VTAIL.n27 VTAIL.n26 185
R1000 VTAIL.n29 VTAIL.n28 185
R1001 VTAIL.n6 VTAIL.n5 185
R1002 VTAIL.n36 VTAIL.n35 185
R1003 VTAIL.n37 VTAIL.n4 185
R1004 VTAIL.n39 VTAIL.n38 185
R1005 VTAIL.n135 VTAIL.n134 185
R1006 VTAIL.n133 VTAIL.n100 185
R1007 VTAIL.n132 VTAIL.n131 185
R1008 VTAIL.n103 VTAIL.n101 185
R1009 VTAIL.n126 VTAIL.n125 185
R1010 VTAIL.n124 VTAIL.n123 185
R1011 VTAIL.n107 VTAIL.n106 185
R1012 VTAIL.n118 VTAIL.n117 185
R1013 VTAIL.n116 VTAIL.n115 185
R1014 VTAIL.n111 VTAIL.n110 185
R1015 VTAIL.n89 VTAIL.n88 185
R1016 VTAIL.n87 VTAIL.n54 185
R1017 VTAIL.n86 VTAIL.n85 185
R1018 VTAIL.n57 VTAIL.n55 185
R1019 VTAIL.n80 VTAIL.n79 185
R1020 VTAIL.n78 VTAIL.n77 185
R1021 VTAIL.n61 VTAIL.n60 185
R1022 VTAIL.n72 VTAIL.n71 185
R1023 VTAIL.n70 VTAIL.n69 185
R1024 VTAIL.n65 VTAIL.n64 185
R1025 VTAIL.n153 VTAIL.t16 149.524
R1026 VTAIL.n15 VTAIL.t0 149.524
R1027 VTAIL.n112 VTAIL.t18 149.524
R1028 VTAIL.n66 VTAIL.t7 149.524
R1029 VTAIL.n157 VTAIL.n151 104.615
R1030 VTAIL.n158 VTAIL.n157 104.615
R1031 VTAIL.n158 VTAIL.n147 104.615
R1032 VTAIL.n165 VTAIL.n147 104.615
R1033 VTAIL.n166 VTAIL.n165 104.615
R1034 VTAIL.n166 VTAIL.n143 104.615
R1035 VTAIL.n174 VTAIL.n143 104.615
R1036 VTAIL.n175 VTAIL.n174 104.615
R1037 VTAIL.n176 VTAIL.n175 104.615
R1038 VTAIL.n19 VTAIL.n13 104.615
R1039 VTAIL.n20 VTAIL.n19 104.615
R1040 VTAIL.n20 VTAIL.n9 104.615
R1041 VTAIL.n27 VTAIL.n9 104.615
R1042 VTAIL.n28 VTAIL.n27 104.615
R1043 VTAIL.n28 VTAIL.n5 104.615
R1044 VTAIL.n36 VTAIL.n5 104.615
R1045 VTAIL.n37 VTAIL.n36 104.615
R1046 VTAIL.n38 VTAIL.n37 104.615
R1047 VTAIL.n134 VTAIL.n133 104.615
R1048 VTAIL.n133 VTAIL.n132 104.615
R1049 VTAIL.n132 VTAIL.n101 104.615
R1050 VTAIL.n125 VTAIL.n101 104.615
R1051 VTAIL.n125 VTAIL.n124 104.615
R1052 VTAIL.n124 VTAIL.n106 104.615
R1053 VTAIL.n117 VTAIL.n106 104.615
R1054 VTAIL.n117 VTAIL.n116 104.615
R1055 VTAIL.n116 VTAIL.n110 104.615
R1056 VTAIL.n88 VTAIL.n87 104.615
R1057 VTAIL.n87 VTAIL.n86 104.615
R1058 VTAIL.n86 VTAIL.n55 104.615
R1059 VTAIL.n79 VTAIL.n55 104.615
R1060 VTAIL.n79 VTAIL.n78 104.615
R1061 VTAIL.n78 VTAIL.n60 104.615
R1062 VTAIL.n71 VTAIL.n60 104.615
R1063 VTAIL.n71 VTAIL.n70 104.615
R1064 VTAIL.n70 VTAIL.n64 104.615
R1065 VTAIL.t16 VTAIL.n151 52.3082
R1066 VTAIL.t0 VTAIL.n13 52.3082
R1067 VTAIL.t18 VTAIL.n110 52.3082
R1068 VTAIL.t7 VTAIL.n64 52.3082
R1069 VTAIL.n97 VTAIL.n96 50.4022
R1070 VTAIL.n95 VTAIL.n94 50.4022
R1071 VTAIL.n51 VTAIL.n50 50.4022
R1072 VTAIL.n49 VTAIL.n48 50.4022
R1073 VTAIL.n183 VTAIL.n182 50.402
R1074 VTAIL.n1 VTAIL.n0 50.402
R1075 VTAIL.n45 VTAIL.n44 50.402
R1076 VTAIL.n47 VTAIL.n46 50.402
R1077 VTAIL.n181 VTAIL.n180 35.2884
R1078 VTAIL.n43 VTAIL.n42 35.2884
R1079 VTAIL.n139 VTAIL.n138 35.2884
R1080 VTAIL.n93 VTAIL.n92 35.2884
R1081 VTAIL.n49 VTAIL.n47 20.2807
R1082 VTAIL.n181 VTAIL.n139 19.7548
R1083 VTAIL.n177 VTAIL.n142 13.1884
R1084 VTAIL.n39 VTAIL.n4 13.1884
R1085 VTAIL.n135 VTAIL.n100 13.1884
R1086 VTAIL.n89 VTAIL.n54 13.1884
R1087 VTAIL.n173 VTAIL.n172 12.8005
R1088 VTAIL.n178 VTAIL.n140 12.8005
R1089 VTAIL.n35 VTAIL.n34 12.8005
R1090 VTAIL.n40 VTAIL.n2 12.8005
R1091 VTAIL.n136 VTAIL.n98 12.8005
R1092 VTAIL.n131 VTAIL.n102 12.8005
R1093 VTAIL.n90 VTAIL.n52 12.8005
R1094 VTAIL.n85 VTAIL.n56 12.8005
R1095 VTAIL.n171 VTAIL.n144 12.0247
R1096 VTAIL.n33 VTAIL.n6 12.0247
R1097 VTAIL.n130 VTAIL.n103 12.0247
R1098 VTAIL.n84 VTAIL.n57 12.0247
R1099 VTAIL.n168 VTAIL.n167 11.249
R1100 VTAIL.n30 VTAIL.n29 11.249
R1101 VTAIL.n127 VTAIL.n126 11.249
R1102 VTAIL.n81 VTAIL.n80 11.249
R1103 VTAIL.n164 VTAIL.n146 10.4732
R1104 VTAIL.n26 VTAIL.n8 10.4732
R1105 VTAIL.n123 VTAIL.n105 10.4732
R1106 VTAIL.n77 VTAIL.n59 10.4732
R1107 VTAIL.n153 VTAIL.n152 10.2747
R1108 VTAIL.n15 VTAIL.n14 10.2747
R1109 VTAIL.n112 VTAIL.n111 10.2747
R1110 VTAIL.n66 VTAIL.n65 10.2747
R1111 VTAIL.n163 VTAIL.n148 9.69747
R1112 VTAIL.n25 VTAIL.n10 9.69747
R1113 VTAIL.n122 VTAIL.n107 9.69747
R1114 VTAIL.n76 VTAIL.n61 9.69747
R1115 VTAIL.n180 VTAIL.n179 9.45567
R1116 VTAIL.n42 VTAIL.n41 9.45567
R1117 VTAIL.n138 VTAIL.n137 9.45567
R1118 VTAIL.n92 VTAIL.n91 9.45567
R1119 VTAIL.n179 VTAIL.n178 9.3005
R1120 VTAIL.n155 VTAIL.n154 9.3005
R1121 VTAIL.n150 VTAIL.n149 9.3005
R1122 VTAIL.n161 VTAIL.n160 9.3005
R1123 VTAIL.n163 VTAIL.n162 9.3005
R1124 VTAIL.n146 VTAIL.n145 9.3005
R1125 VTAIL.n169 VTAIL.n168 9.3005
R1126 VTAIL.n171 VTAIL.n170 9.3005
R1127 VTAIL.n172 VTAIL.n141 9.3005
R1128 VTAIL.n41 VTAIL.n40 9.3005
R1129 VTAIL.n17 VTAIL.n16 9.3005
R1130 VTAIL.n12 VTAIL.n11 9.3005
R1131 VTAIL.n23 VTAIL.n22 9.3005
R1132 VTAIL.n25 VTAIL.n24 9.3005
R1133 VTAIL.n8 VTAIL.n7 9.3005
R1134 VTAIL.n31 VTAIL.n30 9.3005
R1135 VTAIL.n33 VTAIL.n32 9.3005
R1136 VTAIL.n34 VTAIL.n3 9.3005
R1137 VTAIL.n114 VTAIL.n113 9.3005
R1138 VTAIL.n109 VTAIL.n108 9.3005
R1139 VTAIL.n120 VTAIL.n119 9.3005
R1140 VTAIL.n122 VTAIL.n121 9.3005
R1141 VTAIL.n105 VTAIL.n104 9.3005
R1142 VTAIL.n128 VTAIL.n127 9.3005
R1143 VTAIL.n130 VTAIL.n129 9.3005
R1144 VTAIL.n102 VTAIL.n99 9.3005
R1145 VTAIL.n137 VTAIL.n136 9.3005
R1146 VTAIL.n68 VTAIL.n67 9.3005
R1147 VTAIL.n63 VTAIL.n62 9.3005
R1148 VTAIL.n74 VTAIL.n73 9.3005
R1149 VTAIL.n76 VTAIL.n75 9.3005
R1150 VTAIL.n59 VTAIL.n58 9.3005
R1151 VTAIL.n82 VTAIL.n81 9.3005
R1152 VTAIL.n84 VTAIL.n83 9.3005
R1153 VTAIL.n56 VTAIL.n53 9.3005
R1154 VTAIL.n91 VTAIL.n90 9.3005
R1155 VTAIL.n160 VTAIL.n159 8.92171
R1156 VTAIL.n22 VTAIL.n21 8.92171
R1157 VTAIL.n119 VTAIL.n118 8.92171
R1158 VTAIL.n73 VTAIL.n72 8.92171
R1159 VTAIL.n156 VTAIL.n150 8.14595
R1160 VTAIL.n18 VTAIL.n12 8.14595
R1161 VTAIL.n115 VTAIL.n109 8.14595
R1162 VTAIL.n69 VTAIL.n63 8.14595
R1163 VTAIL.n155 VTAIL.n152 7.3702
R1164 VTAIL.n17 VTAIL.n14 7.3702
R1165 VTAIL.n114 VTAIL.n111 7.3702
R1166 VTAIL.n68 VTAIL.n65 7.3702
R1167 VTAIL.n156 VTAIL.n155 5.81868
R1168 VTAIL.n18 VTAIL.n17 5.81868
R1169 VTAIL.n115 VTAIL.n114 5.81868
R1170 VTAIL.n69 VTAIL.n68 5.81868
R1171 VTAIL.n159 VTAIL.n150 5.04292
R1172 VTAIL.n21 VTAIL.n12 5.04292
R1173 VTAIL.n118 VTAIL.n109 5.04292
R1174 VTAIL.n72 VTAIL.n63 5.04292
R1175 VTAIL.n160 VTAIL.n148 4.26717
R1176 VTAIL.n22 VTAIL.n10 4.26717
R1177 VTAIL.n119 VTAIL.n107 4.26717
R1178 VTAIL.n73 VTAIL.n61 4.26717
R1179 VTAIL.n164 VTAIL.n163 3.49141
R1180 VTAIL.n26 VTAIL.n25 3.49141
R1181 VTAIL.n123 VTAIL.n122 3.49141
R1182 VTAIL.n77 VTAIL.n76 3.49141
R1183 VTAIL.n154 VTAIL.n153 2.84304
R1184 VTAIL.n16 VTAIL.n15 2.84304
R1185 VTAIL.n113 VTAIL.n112 2.84304
R1186 VTAIL.n67 VTAIL.n66 2.84304
R1187 VTAIL.n167 VTAIL.n146 2.71565
R1188 VTAIL.n29 VTAIL.n8 2.71565
R1189 VTAIL.n126 VTAIL.n105 2.71565
R1190 VTAIL.n80 VTAIL.n59 2.71565
R1191 VTAIL.n182 VTAIL.t14 2.48794
R1192 VTAIL.n182 VTAIL.t13 2.48794
R1193 VTAIL.n0 VTAIL.t10 2.48794
R1194 VTAIL.n0 VTAIL.t12 2.48794
R1195 VTAIL.n44 VTAIL.t19 2.48794
R1196 VTAIL.n44 VTAIL.t3 2.48794
R1197 VTAIL.n46 VTAIL.t17 2.48794
R1198 VTAIL.n46 VTAIL.t6 2.48794
R1199 VTAIL.n96 VTAIL.t5 2.48794
R1200 VTAIL.n96 VTAIL.t4 2.48794
R1201 VTAIL.n94 VTAIL.t1 2.48794
R1202 VTAIL.n94 VTAIL.t2 2.48794
R1203 VTAIL.n50 VTAIL.t15 2.48794
R1204 VTAIL.n50 VTAIL.t8 2.48794
R1205 VTAIL.n48 VTAIL.t11 2.48794
R1206 VTAIL.n48 VTAIL.t9 2.48794
R1207 VTAIL.n168 VTAIL.n144 1.93989
R1208 VTAIL.n30 VTAIL.n6 1.93989
R1209 VTAIL.n127 VTAIL.n103 1.93989
R1210 VTAIL.n81 VTAIL.n57 1.93989
R1211 VTAIL.n173 VTAIL.n171 1.16414
R1212 VTAIL.n180 VTAIL.n140 1.16414
R1213 VTAIL.n35 VTAIL.n33 1.16414
R1214 VTAIL.n42 VTAIL.n2 1.16414
R1215 VTAIL.n138 VTAIL.n98 1.16414
R1216 VTAIL.n131 VTAIL.n130 1.16414
R1217 VTAIL.n92 VTAIL.n52 1.16414
R1218 VTAIL.n85 VTAIL.n84 1.16414
R1219 VTAIL.n95 VTAIL.n93 0.733259
R1220 VTAIL.n43 VTAIL.n1 0.733259
R1221 VTAIL.n51 VTAIL.n49 0.526362
R1222 VTAIL.n93 VTAIL.n51 0.526362
R1223 VTAIL.n97 VTAIL.n95 0.526362
R1224 VTAIL.n139 VTAIL.n97 0.526362
R1225 VTAIL.n47 VTAIL.n45 0.526362
R1226 VTAIL.n45 VTAIL.n43 0.526362
R1227 VTAIL.n183 VTAIL.n181 0.526362
R1228 VTAIL VTAIL.n1 0.453086
R1229 VTAIL.n172 VTAIL.n142 0.388379
R1230 VTAIL.n178 VTAIL.n177 0.388379
R1231 VTAIL.n34 VTAIL.n4 0.388379
R1232 VTAIL.n40 VTAIL.n39 0.388379
R1233 VTAIL.n136 VTAIL.n135 0.388379
R1234 VTAIL.n102 VTAIL.n100 0.388379
R1235 VTAIL.n90 VTAIL.n89 0.388379
R1236 VTAIL.n56 VTAIL.n54 0.388379
R1237 VTAIL.n154 VTAIL.n149 0.155672
R1238 VTAIL.n161 VTAIL.n149 0.155672
R1239 VTAIL.n162 VTAIL.n161 0.155672
R1240 VTAIL.n162 VTAIL.n145 0.155672
R1241 VTAIL.n169 VTAIL.n145 0.155672
R1242 VTAIL.n170 VTAIL.n169 0.155672
R1243 VTAIL.n170 VTAIL.n141 0.155672
R1244 VTAIL.n179 VTAIL.n141 0.155672
R1245 VTAIL.n16 VTAIL.n11 0.155672
R1246 VTAIL.n23 VTAIL.n11 0.155672
R1247 VTAIL.n24 VTAIL.n23 0.155672
R1248 VTAIL.n24 VTAIL.n7 0.155672
R1249 VTAIL.n31 VTAIL.n7 0.155672
R1250 VTAIL.n32 VTAIL.n31 0.155672
R1251 VTAIL.n32 VTAIL.n3 0.155672
R1252 VTAIL.n41 VTAIL.n3 0.155672
R1253 VTAIL.n137 VTAIL.n99 0.155672
R1254 VTAIL.n129 VTAIL.n99 0.155672
R1255 VTAIL.n129 VTAIL.n128 0.155672
R1256 VTAIL.n128 VTAIL.n104 0.155672
R1257 VTAIL.n121 VTAIL.n104 0.155672
R1258 VTAIL.n121 VTAIL.n120 0.155672
R1259 VTAIL.n120 VTAIL.n108 0.155672
R1260 VTAIL.n113 VTAIL.n108 0.155672
R1261 VTAIL.n91 VTAIL.n53 0.155672
R1262 VTAIL.n83 VTAIL.n53 0.155672
R1263 VTAIL.n83 VTAIL.n82 0.155672
R1264 VTAIL.n82 VTAIL.n58 0.155672
R1265 VTAIL.n75 VTAIL.n58 0.155672
R1266 VTAIL.n75 VTAIL.n74 0.155672
R1267 VTAIL.n74 VTAIL.n62 0.155672
R1268 VTAIL.n67 VTAIL.n62 0.155672
R1269 VTAIL VTAIL.n183 0.0737759
R1270 VDD2.n81 VDD2.n45 289.615
R1271 VDD2.n36 VDD2.n0 289.615
R1272 VDD2.n82 VDD2.n81 185
R1273 VDD2.n80 VDD2.n47 185
R1274 VDD2.n79 VDD2.n78 185
R1275 VDD2.n50 VDD2.n48 185
R1276 VDD2.n73 VDD2.n72 185
R1277 VDD2.n71 VDD2.n70 185
R1278 VDD2.n54 VDD2.n53 185
R1279 VDD2.n65 VDD2.n64 185
R1280 VDD2.n63 VDD2.n62 185
R1281 VDD2.n58 VDD2.n57 185
R1282 VDD2.n12 VDD2.n11 185
R1283 VDD2.n17 VDD2.n16 185
R1284 VDD2.n19 VDD2.n18 185
R1285 VDD2.n8 VDD2.n7 185
R1286 VDD2.n25 VDD2.n24 185
R1287 VDD2.n27 VDD2.n26 185
R1288 VDD2.n4 VDD2.n3 185
R1289 VDD2.n34 VDD2.n33 185
R1290 VDD2.n35 VDD2.n2 185
R1291 VDD2.n37 VDD2.n36 185
R1292 VDD2.n59 VDD2.t9 149.524
R1293 VDD2.n13 VDD2.t4 149.524
R1294 VDD2.n81 VDD2.n80 104.615
R1295 VDD2.n80 VDD2.n79 104.615
R1296 VDD2.n79 VDD2.n48 104.615
R1297 VDD2.n72 VDD2.n48 104.615
R1298 VDD2.n72 VDD2.n71 104.615
R1299 VDD2.n71 VDD2.n53 104.615
R1300 VDD2.n64 VDD2.n53 104.615
R1301 VDD2.n64 VDD2.n63 104.615
R1302 VDD2.n63 VDD2.n57 104.615
R1303 VDD2.n17 VDD2.n11 104.615
R1304 VDD2.n18 VDD2.n17 104.615
R1305 VDD2.n18 VDD2.n7 104.615
R1306 VDD2.n25 VDD2.n7 104.615
R1307 VDD2.n26 VDD2.n25 104.615
R1308 VDD2.n26 VDD2.n3 104.615
R1309 VDD2.n34 VDD2.n3 104.615
R1310 VDD2.n35 VDD2.n34 104.615
R1311 VDD2.n36 VDD2.n35 104.615
R1312 VDD2.n44 VDD2.n43 67.4199
R1313 VDD2 VDD2.n89 67.417
R1314 VDD2.n88 VDD2.n87 67.081
R1315 VDD2.n42 VDD2.n41 67.0808
R1316 VDD2.n42 VDD2.n40 52.493
R1317 VDD2.t9 VDD2.n57 52.3082
R1318 VDD2.t4 VDD2.n11 52.3082
R1319 VDD2.n86 VDD2.n85 51.9672
R1320 VDD2.n86 VDD2.n44 33.0752
R1321 VDD2.n82 VDD2.n47 13.1884
R1322 VDD2.n37 VDD2.n2 13.1884
R1323 VDD2.n83 VDD2.n45 12.8005
R1324 VDD2.n78 VDD2.n49 12.8005
R1325 VDD2.n33 VDD2.n32 12.8005
R1326 VDD2.n38 VDD2.n0 12.8005
R1327 VDD2.n77 VDD2.n50 12.0247
R1328 VDD2.n31 VDD2.n4 12.0247
R1329 VDD2.n74 VDD2.n73 11.249
R1330 VDD2.n28 VDD2.n27 11.249
R1331 VDD2.n70 VDD2.n52 10.4732
R1332 VDD2.n24 VDD2.n6 10.4732
R1333 VDD2.n59 VDD2.n58 10.2747
R1334 VDD2.n13 VDD2.n12 10.2747
R1335 VDD2.n69 VDD2.n54 9.69747
R1336 VDD2.n23 VDD2.n8 9.69747
R1337 VDD2.n85 VDD2.n84 9.45567
R1338 VDD2.n40 VDD2.n39 9.45567
R1339 VDD2.n61 VDD2.n60 9.3005
R1340 VDD2.n56 VDD2.n55 9.3005
R1341 VDD2.n67 VDD2.n66 9.3005
R1342 VDD2.n69 VDD2.n68 9.3005
R1343 VDD2.n52 VDD2.n51 9.3005
R1344 VDD2.n75 VDD2.n74 9.3005
R1345 VDD2.n77 VDD2.n76 9.3005
R1346 VDD2.n49 VDD2.n46 9.3005
R1347 VDD2.n84 VDD2.n83 9.3005
R1348 VDD2.n39 VDD2.n38 9.3005
R1349 VDD2.n15 VDD2.n14 9.3005
R1350 VDD2.n10 VDD2.n9 9.3005
R1351 VDD2.n21 VDD2.n20 9.3005
R1352 VDD2.n23 VDD2.n22 9.3005
R1353 VDD2.n6 VDD2.n5 9.3005
R1354 VDD2.n29 VDD2.n28 9.3005
R1355 VDD2.n31 VDD2.n30 9.3005
R1356 VDD2.n32 VDD2.n1 9.3005
R1357 VDD2.n66 VDD2.n65 8.92171
R1358 VDD2.n20 VDD2.n19 8.92171
R1359 VDD2.n62 VDD2.n56 8.14595
R1360 VDD2.n16 VDD2.n10 8.14595
R1361 VDD2.n61 VDD2.n58 7.3702
R1362 VDD2.n15 VDD2.n12 7.3702
R1363 VDD2.n62 VDD2.n61 5.81868
R1364 VDD2.n16 VDD2.n15 5.81868
R1365 VDD2.n65 VDD2.n56 5.04292
R1366 VDD2.n19 VDD2.n10 5.04292
R1367 VDD2.n66 VDD2.n54 4.26717
R1368 VDD2.n20 VDD2.n8 4.26717
R1369 VDD2.n70 VDD2.n69 3.49141
R1370 VDD2.n24 VDD2.n23 3.49141
R1371 VDD2.n60 VDD2.n59 2.84304
R1372 VDD2.n14 VDD2.n13 2.84304
R1373 VDD2.n73 VDD2.n52 2.71565
R1374 VDD2.n27 VDD2.n6 2.71565
R1375 VDD2.n89 VDD2.t7 2.48794
R1376 VDD2.n89 VDD2.t3 2.48794
R1377 VDD2.n87 VDD2.t5 2.48794
R1378 VDD2.n87 VDD2.t1 2.48794
R1379 VDD2.n43 VDD2.t8 2.48794
R1380 VDD2.n43 VDD2.t0 2.48794
R1381 VDD2.n41 VDD2.t2 2.48794
R1382 VDD2.n41 VDD2.t6 2.48794
R1383 VDD2.n74 VDD2.n50 1.93989
R1384 VDD2.n28 VDD2.n4 1.93989
R1385 VDD2.n85 VDD2.n45 1.16414
R1386 VDD2.n78 VDD2.n77 1.16414
R1387 VDD2.n33 VDD2.n31 1.16414
R1388 VDD2.n40 VDD2.n0 1.16414
R1389 VDD2.n88 VDD2.n86 0.526362
R1390 VDD2.n83 VDD2.n82 0.388379
R1391 VDD2.n49 VDD2.n47 0.388379
R1392 VDD2.n32 VDD2.n2 0.388379
R1393 VDD2.n38 VDD2.n37 0.388379
R1394 VDD2 VDD2.n88 0.190155
R1395 VDD2.n84 VDD2.n46 0.155672
R1396 VDD2.n76 VDD2.n46 0.155672
R1397 VDD2.n76 VDD2.n75 0.155672
R1398 VDD2.n75 VDD2.n51 0.155672
R1399 VDD2.n68 VDD2.n51 0.155672
R1400 VDD2.n68 VDD2.n67 0.155672
R1401 VDD2.n67 VDD2.n55 0.155672
R1402 VDD2.n60 VDD2.n55 0.155672
R1403 VDD2.n14 VDD2.n9 0.155672
R1404 VDD2.n21 VDD2.n9 0.155672
R1405 VDD2.n22 VDD2.n21 0.155672
R1406 VDD2.n22 VDD2.n5 0.155672
R1407 VDD2.n29 VDD2.n5 0.155672
R1408 VDD2.n30 VDD2.n29 0.155672
R1409 VDD2.n30 VDD2.n1 0.155672
R1410 VDD2.n39 VDD2.n1 0.155672
R1411 VDD2.n44 VDD2.n42 0.0766195
R1412 VP.n21 VP.t4 830.876
R1413 VP.n14 VP.t7 830.876
R1414 VP.n5 VP.t5 830.876
R1415 VP.n11 VP.t8 830.876
R1416 VP.n18 VP.t9 798.744
R1417 VP.n20 VP.t2 798.744
R1418 VP.n13 VP.t0 798.744
R1419 VP.n8 VP.t6 798.744
R1420 VP.n4 VP.t1 798.744
R1421 VP.n10 VP.t3 798.744
R1422 VP.n6 VP.n5 161.489
R1423 VP.n22 VP.n21 161.3
R1424 VP.n6 VP.n3 161.3
R1425 VP.n8 VP.n7 161.3
R1426 VP.n9 VP.n2 161.3
R1427 VP.n12 VP.n11 161.3
R1428 VP.n19 VP.n0 161.3
R1429 VP.n18 VP.n17 161.3
R1430 VP.n16 VP.n1 161.3
R1431 VP.n15 VP.n14 161.3
R1432 VP.n18 VP.n1 73.0308
R1433 VP.n19 VP.n18 73.0308
R1434 VP.n8 VP.n3 73.0308
R1435 VP.n9 VP.n8 73.0308
R1436 VP.n14 VP.n13 56.9641
R1437 VP.n21 VP.n20 56.9641
R1438 VP.n5 VP.n4 56.9641
R1439 VP.n11 VP.n10 56.9641
R1440 VP.n15 VP.n12 37.4588
R1441 VP.n13 VP.n1 16.0672
R1442 VP.n20 VP.n19 16.0672
R1443 VP.n4 VP.n3 16.0672
R1444 VP.n10 VP.n9 16.0672
R1445 VP.n7 VP.n6 0.189894
R1446 VP.n7 VP.n2 0.189894
R1447 VP.n12 VP.n2 0.189894
R1448 VP.n16 VP.n15 0.189894
R1449 VP.n17 VP.n16 0.189894
R1450 VP.n17 VP.n0 0.189894
R1451 VP.n22 VP.n0 0.189894
R1452 VP VP.n22 0.0516364
R1453 VDD1.n36 VDD1.n0 289.615
R1454 VDD1.n79 VDD1.n43 289.615
R1455 VDD1.n37 VDD1.n36 185
R1456 VDD1.n35 VDD1.n2 185
R1457 VDD1.n34 VDD1.n33 185
R1458 VDD1.n5 VDD1.n3 185
R1459 VDD1.n28 VDD1.n27 185
R1460 VDD1.n26 VDD1.n25 185
R1461 VDD1.n9 VDD1.n8 185
R1462 VDD1.n20 VDD1.n19 185
R1463 VDD1.n18 VDD1.n17 185
R1464 VDD1.n13 VDD1.n12 185
R1465 VDD1.n55 VDD1.n54 185
R1466 VDD1.n60 VDD1.n59 185
R1467 VDD1.n62 VDD1.n61 185
R1468 VDD1.n51 VDD1.n50 185
R1469 VDD1.n68 VDD1.n67 185
R1470 VDD1.n70 VDD1.n69 185
R1471 VDD1.n47 VDD1.n46 185
R1472 VDD1.n77 VDD1.n76 185
R1473 VDD1.n78 VDD1.n45 185
R1474 VDD1.n80 VDD1.n79 185
R1475 VDD1.n14 VDD1.t4 149.524
R1476 VDD1.n56 VDD1.t2 149.524
R1477 VDD1.n36 VDD1.n35 104.615
R1478 VDD1.n35 VDD1.n34 104.615
R1479 VDD1.n34 VDD1.n3 104.615
R1480 VDD1.n27 VDD1.n3 104.615
R1481 VDD1.n27 VDD1.n26 104.615
R1482 VDD1.n26 VDD1.n8 104.615
R1483 VDD1.n19 VDD1.n8 104.615
R1484 VDD1.n19 VDD1.n18 104.615
R1485 VDD1.n18 VDD1.n12 104.615
R1486 VDD1.n60 VDD1.n54 104.615
R1487 VDD1.n61 VDD1.n60 104.615
R1488 VDD1.n61 VDD1.n50 104.615
R1489 VDD1.n68 VDD1.n50 104.615
R1490 VDD1.n69 VDD1.n68 104.615
R1491 VDD1.n69 VDD1.n46 104.615
R1492 VDD1.n77 VDD1.n46 104.615
R1493 VDD1.n78 VDD1.n77 104.615
R1494 VDD1.n79 VDD1.n78 104.615
R1495 VDD1.n87 VDD1.n86 67.4199
R1496 VDD1.n42 VDD1.n41 67.081
R1497 VDD1.n89 VDD1.n88 67.0808
R1498 VDD1.n85 VDD1.n84 67.0808
R1499 VDD1.n42 VDD1.n40 52.493
R1500 VDD1.n85 VDD1.n83 52.493
R1501 VDD1.t4 VDD1.n12 52.3082
R1502 VDD1.t2 VDD1.n54 52.3082
R1503 VDD1.n89 VDD1.n87 33.9212
R1504 VDD1.n37 VDD1.n2 13.1884
R1505 VDD1.n80 VDD1.n45 13.1884
R1506 VDD1.n38 VDD1.n0 12.8005
R1507 VDD1.n33 VDD1.n4 12.8005
R1508 VDD1.n76 VDD1.n75 12.8005
R1509 VDD1.n81 VDD1.n43 12.8005
R1510 VDD1.n32 VDD1.n5 12.0247
R1511 VDD1.n74 VDD1.n47 12.0247
R1512 VDD1.n29 VDD1.n28 11.249
R1513 VDD1.n71 VDD1.n70 11.249
R1514 VDD1.n25 VDD1.n7 10.4732
R1515 VDD1.n67 VDD1.n49 10.4732
R1516 VDD1.n14 VDD1.n13 10.2747
R1517 VDD1.n56 VDD1.n55 10.2747
R1518 VDD1.n24 VDD1.n9 9.69747
R1519 VDD1.n66 VDD1.n51 9.69747
R1520 VDD1.n40 VDD1.n39 9.45567
R1521 VDD1.n83 VDD1.n82 9.45567
R1522 VDD1.n16 VDD1.n15 9.3005
R1523 VDD1.n11 VDD1.n10 9.3005
R1524 VDD1.n22 VDD1.n21 9.3005
R1525 VDD1.n24 VDD1.n23 9.3005
R1526 VDD1.n7 VDD1.n6 9.3005
R1527 VDD1.n30 VDD1.n29 9.3005
R1528 VDD1.n32 VDD1.n31 9.3005
R1529 VDD1.n4 VDD1.n1 9.3005
R1530 VDD1.n39 VDD1.n38 9.3005
R1531 VDD1.n82 VDD1.n81 9.3005
R1532 VDD1.n58 VDD1.n57 9.3005
R1533 VDD1.n53 VDD1.n52 9.3005
R1534 VDD1.n64 VDD1.n63 9.3005
R1535 VDD1.n66 VDD1.n65 9.3005
R1536 VDD1.n49 VDD1.n48 9.3005
R1537 VDD1.n72 VDD1.n71 9.3005
R1538 VDD1.n74 VDD1.n73 9.3005
R1539 VDD1.n75 VDD1.n44 9.3005
R1540 VDD1.n21 VDD1.n20 8.92171
R1541 VDD1.n63 VDD1.n62 8.92171
R1542 VDD1.n17 VDD1.n11 8.14595
R1543 VDD1.n59 VDD1.n53 8.14595
R1544 VDD1.n16 VDD1.n13 7.3702
R1545 VDD1.n58 VDD1.n55 7.3702
R1546 VDD1.n17 VDD1.n16 5.81868
R1547 VDD1.n59 VDD1.n58 5.81868
R1548 VDD1.n20 VDD1.n11 5.04292
R1549 VDD1.n62 VDD1.n53 5.04292
R1550 VDD1.n21 VDD1.n9 4.26717
R1551 VDD1.n63 VDD1.n51 4.26717
R1552 VDD1.n25 VDD1.n24 3.49141
R1553 VDD1.n67 VDD1.n66 3.49141
R1554 VDD1.n15 VDD1.n14 2.84304
R1555 VDD1.n57 VDD1.n56 2.84304
R1556 VDD1.n28 VDD1.n7 2.71565
R1557 VDD1.n70 VDD1.n49 2.71565
R1558 VDD1.n88 VDD1.t6 2.48794
R1559 VDD1.n88 VDD1.t1 2.48794
R1560 VDD1.n41 VDD1.t8 2.48794
R1561 VDD1.n41 VDD1.t3 2.48794
R1562 VDD1.n86 VDD1.t7 2.48794
R1563 VDD1.n86 VDD1.t5 2.48794
R1564 VDD1.n84 VDD1.t9 2.48794
R1565 VDD1.n84 VDD1.t0 2.48794
R1566 VDD1.n29 VDD1.n5 1.93989
R1567 VDD1.n71 VDD1.n47 1.93989
R1568 VDD1.n40 VDD1.n0 1.16414
R1569 VDD1.n33 VDD1.n32 1.16414
R1570 VDD1.n76 VDD1.n74 1.16414
R1571 VDD1.n83 VDD1.n43 1.16414
R1572 VDD1.n38 VDD1.n37 0.388379
R1573 VDD1.n4 VDD1.n2 0.388379
R1574 VDD1.n75 VDD1.n45 0.388379
R1575 VDD1.n81 VDD1.n80 0.388379
R1576 VDD1 VDD1.n89 0.336707
R1577 VDD1 VDD1.n42 0.190155
R1578 VDD1.n39 VDD1.n1 0.155672
R1579 VDD1.n31 VDD1.n1 0.155672
R1580 VDD1.n31 VDD1.n30 0.155672
R1581 VDD1.n30 VDD1.n6 0.155672
R1582 VDD1.n23 VDD1.n6 0.155672
R1583 VDD1.n23 VDD1.n22 0.155672
R1584 VDD1.n22 VDD1.n10 0.155672
R1585 VDD1.n15 VDD1.n10 0.155672
R1586 VDD1.n57 VDD1.n52 0.155672
R1587 VDD1.n64 VDD1.n52 0.155672
R1588 VDD1.n65 VDD1.n64 0.155672
R1589 VDD1.n65 VDD1.n48 0.155672
R1590 VDD1.n72 VDD1.n48 0.155672
R1591 VDD1.n73 VDD1.n72 0.155672
R1592 VDD1.n73 VDD1.n44 0.155672
R1593 VDD1.n82 VDD1.n44 0.155672
R1594 VDD1.n87 VDD1.n85 0.0766195
C0 VP VTAIL 2.42886f
C1 VN VTAIL 2.41431f
C2 VP VDD2 0.287148f
C3 VDD2 VN 2.64938f
C4 VP VDD1 2.78531f
C5 VDD1 VN 0.147697f
C6 VDD2 VTAIL 15.0214f
C7 VDD1 VTAIL 14.989f
C8 VP VN 4.23482f
C9 VDD1 VDD2 0.712485f
C10 VDD2 B 3.788507f
C11 VDD1 B 3.65377f
C12 VTAIL B 4.638877f
C13 VN B 7.14291f
C14 VP B 5.204889f
C15 VDD1.n0 B 0.040857f
C16 VDD1.n1 B 0.030228f
C17 VDD1.n2 B 0.016721f
C18 VDD1.n3 B 0.038394f
C19 VDD1.n4 B 0.016243f
C20 VDD1.n5 B 0.017199f
C21 VDD1.n6 B 0.030228f
C22 VDD1.n7 B 0.016243f
C23 VDD1.n8 B 0.038394f
C24 VDD1.n9 B 0.017199f
C25 VDD1.n10 B 0.030228f
C26 VDD1.n11 B 0.016243f
C27 VDD1.n12 B 0.028795f
C28 VDD1.n13 B 0.027141f
C29 VDD1.t4 B 0.064209f
C30 VDD1.n14 B 0.171097f
C31 VDD1.n15 B 0.981723f
C32 VDD1.n16 B 0.016243f
C33 VDD1.n17 B 0.017199f
C34 VDD1.n18 B 0.038394f
C35 VDD1.n19 B 0.038394f
C36 VDD1.n20 B 0.017199f
C37 VDD1.n21 B 0.016243f
C38 VDD1.n22 B 0.030228f
C39 VDD1.n23 B 0.030228f
C40 VDD1.n24 B 0.016243f
C41 VDD1.n25 B 0.017199f
C42 VDD1.n26 B 0.038394f
C43 VDD1.n27 B 0.038394f
C44 VDD1.n28 B 0.017199f
C45 VDD1.n29 B 0.016243f
C46 VDD1.n30 B 0.030228f
C47 VDD1.n31 B 0.030228f
C48 VDD1.n32 B 0.016243f
C49 VDD1.n33 B 0.017199f
C50 VDD1.n34 B 0.038394f
C51 VDD1.n35 B 0.038394f
C52 VDD1.n36 B 0.08023f
C53 VDD1.n37 B 0.016721f
C54 VDD1.n38 B 0.016243f
C55 VDD1.n39 B 0.076479f
C56 VDD1.n40 B 0.066749f
C57 VDD1.t8 B 0.190143f
C58 VDD1.t3 B 0.190143f
C59 VDD1.n41 B 1.64704f
C60 VDD1.n42 B 0.420891f
C61 VDD1.n43 B 0.040857f
C62 VDD1.n44 B 0.030228f
C63 VDD1.n45 B 0.016721f
C64 VDD1.n46 B 0.038394f
C65 VDD1.n47 B 0.017199f
C66 VDD1.n48 B 0.030228f
C67 VDD1.n49 B 0.016243f
C68 VDD1.n50 B 0.038394f
C69 VDD1.n51 B 0.017199f
C70 VDD1.n52 B 0.030228f
C71 VDD1.n53 B 0.016243f
C72 VDD1.n54 B 0.028795f
C73 VDD1.n55 B 0.027141f
C74 VDD1.t2 B 0.064209f
C75 VDD1.n56 B 0.171097f
C76 VDD1.n57 B 0.981723f
C77 VDD1.n58 B 0.016243f
C78 VDD1.n59 B 0.017199f
C79 VDD1.n60 B 0.038394f
C80 VDD1.n61 B 0.038394f
C81 VDD1.n62 B 0.017199f
C82 VDD1.n63 B 0.016243f
C83 VDD1.n64 B 0.030228f
C84 VDD1.n65 B 0.030228f
C85 VDD1.n66 B 0.016243f
C86 VDD1.n67 B 0.017199f
C87 VDD1.n68 B 0.038394f
C88 VDD1.n69 B 0.038394f
C89 VDD1.n70 B 0.017199f
C90 VDD1.n71 B 0.016243f
C91 VDD1.n72 B 0.030228f
C92 VDD1.n73 B 0.030228f
C93 VDD1.n74 B 0.016243f
C94 VDD1.n75 B 0.016243f
C95 VDD1.n76 B 0.017199f
C96 VDD1.n77 B 0.038394f
C97 VDD1.n78 B 0.038394f
C98 VDD1.n79 B 0.08023f
C99 VDD1.n80 B 0.016721f
C100 VDD1.n81 B 0.016243f
C101 VDD1.n82 B 0.076479f
C102 VDD1.n83 B 0.066749f
C103 VDD1.t9 B 0.190143f
C104 VDD1.t0 B 0.190143f
C105 VDD1.n84 B 1.64703f
C106 VDD1.n85 B 0.419046f
C107 VDD1.t7 B 0.190143f
C108 VDD1.t5 B 0.190143f
C109 VDD1.n86 B 1.64873f
C110 VDD1.n87 B 1.80549f
C111 VDD1.t6 B 0.190143f
C112 VDD1.t1 B 0.190143f
C113 VDD1.n88 B 1.64703f
C114 VDD1.n89 B 2.28027f
C115 VP.n0 B 0.054839f
C116 VP.t2 B 0.34712f
C117 VP.t9 B 0.34712f
C118 VP.n1 B 0.021911f
C119 VP.n2 B 0.054839f
C120 VP.t3 B 0.34712f
C121 VP.t6 B 0.34712f
C122 VP.n3 B 0.021911f
C123 VP.t5 B 0.352922f
C124 VP.t1 B 0.34712f
C125 VP.n4 B 0.150016f
C126 VP.n5 B 0.166198f
C127 VP.n6 B 0.117042f
C128 VP.n7 B 0.054839f
C129 VP.n8 B 0.168207f
C130 VP.n9 B 0.021911f
C131 VP.n10 B 0.150016f
C132 VP.t8 B 0.352922f
C133 VP.n11 B 0.166125f
C134 VP.n12 B 1.85546f
C135 VP.t7 B 0.352922f
C136 VP.t0 B 0.34712f
C137 VP.n13 B 0.150016f
C138 VP.n14 B 0.166125f
C139 VP.n15 B 1.90793f
C140 VP.n16 B 0.054839f
C141 VP.n17 B 0.054839f
C142 VP.n18 B 0.168207f
C143 VP.n19 B 0.021911f
C144 VP.n20 B 0.150016f
C145 VP.t4 B 0.352922f
C146 VP.n21 B 0.166125f
C147 VP.n22 B 0.042498f
C148 VDD2.n0 B 0.040653f
C149 VDD2.n1 B 0.030077f
C150 VDD2.n2 B 0.016638f
C151 VDD2.n3 B 0.038202f
C152 VDD2.n4 B 0.017113f
C153 VDD2.n5 B 0.030077f
C154 VDD2.n6 B 0.016162f
C155 VDD2.n7 B 0.038202f
C156 VDD2.n8 B 0.017113f
C157 VDD2.n9 B 0.030077f
C158 VDD2.n10 B 0.016162f
C159 VDD2.n11 B 0.028651f
C160 VDD2.n12 B 0.027006f
C161 VDD2.t4 B 0.063888f
C162 VDD2.n13 B 0.170242f
C163 VDD2.n14 B 0.976819f
C164 VDD2.n15 B 0.016162f
C165 VDD2.n16 B 0.017113f
C166 VDD2.n17 B 0.038202f
C167 VDD2.n18 B 0.038202f
C168 VDD2.n19 B 0.017113f
C169 VDD2.n20 B 0.016162f
C170 VDD2.n21 B 0.030077f
C171 VDD2.n22 B 0.030077f
C172 VDD2.n23 B 0.016162f
C173 VDD2.n24 B 0.017113f
C174 VDD2.n25 B 0.038202f
C175 VDD2.n26 B 0.038202f
C176 VDD2.n27 B 0.017113f
C177 VDD2.n28 B 0.016162f
C178 VDD2.n29 B 0.030077f
C179 VDD2.n30 B 0.030077f
C180 VDD2.n31 B 0.016162f
C181 VDD2.n32 B 0.016162f
C182 VDD2.n33 B 0.017113f
C183 VDD2.n34 B 0.038202f
C184 VDD2.n35 B 0.038202f
C185 VDD2.n36 B 0.079829f
C186 VDD2.n37 B 0.016638f
C187 VDD2.n38 B 0.016162f
C188 VDD2.n39 B 0.076096f
C189 VDD2.n40 B 0.066416f
C190 VDD2.t2 B 0.189194f
C191 VDD2.t6 B 0.189194f
C192 VDD2.n41 B 1.6388f
C193 VDD2.n42 B 0.416953f
C194 VDD2.t8 B 0.189194f
C195 VDD2.t0 B 0.189194f
C196 VDD2.n43 B 1.64049f
C197 VDD2.n44 B 1.7165f
C198 VDD2.n45 B 0.040653f
C199 VDD2.n46 B 0.030077f
C200 VDD2.n47 B 0.016638f
C201 VDD2.n48 B 0.038202f
C202 VDD2.n49 B 0.016162f
C203 VDD2.n50 B 0.017113f
C204 VDD2.n51 B 0.030077f
C205 VDD2.n52 B 0.016162f
C206 VDD2.n53 B 0.038202f
C207 VDD2.n54 B 0.017113f
C208 VDD2.n55 B 0.030077f
C209 VDD2.n56 B 0.016162f
C210 VDD2.n57 B 0.028651f
C211 VDD2.n58 B 0.027006f
C212 VDD2.t9 B 0.063888f
C213 VDD2.n59 B 0.170242f
C214 VDD2.n60 B 0.976819f
C215 VDD2.n61 B 0.016162f
C216 VDD2.n62 B 0.017113f
C217 VDD2.n63 B 0.038202f
C218 VDD2.n64 B 0.038202f
C219 VDD2.n65 B 0.017113f
C220 VDD2.n66 B 0.016162f
C221 VDD2.n67 B 0.030077f
C222 VDD2.n68 B 0.030077f
C223 VDD2.n69 B 0.016162f
C224 VDD2.n70 B 0.017113f
C225 VDD2.n71 B 0.038202f
C226 VDD2.n72 B 0.038202f
C227 VDD2.n73 B 0.017113f
C228 VDD2.n74 B 0.016162f
C229 VDD2.n75 B 0.030077f
C230 VDD2.n76 B 0.030077f
C231 VDD2.n77 B 0.016162f
C232 VDD2.n78 B 0.017113f
C233 VDD2.n79 B 0.038202f
C234 VDD2.n80 B 0.038202f
C235 VDD2.n81 B 0.079829f
C236 VDD2.n82 B 0.016638f
C237 VDD2.n83 B 0.016162f
C238 VDD2.n84 B 0.076096f
C239 VDD2.n85 B 0.065288f
C240 VDD2.n86 B 2.01682f
C241 VDD2.t5 B 0.189194f
C242 VDD2.t1 B 0.189194f
C243 VDD2.n87 B 1.63881f
C244 VDD2.n88 B 0.307271f
C245 VDD2.t7 B 0.189194f
C246 VDD2.t3 B 0.189194f
C247 VDD2.n89 B 1.64047f
C248 VTAIL.t10 B 0.200601f
C249 VTAIL.t12 B 0.200601f
C250 VTAIL.n0 B 1.65614f
C251 VTAIL.n1 B 0.412214f
C252 VTAIL.n2 B 0.043104f
C253 VTAIL.n3 B 0.031891f
C254 VTAIL.n4 B 0.017641f
C255 VTAIL.n5 B 0.040505f
C256 VTAIL.n6 B 0.018145f
C257 VTAIL.n7 B 0.031891f
C258 VTAIL.n8 B 0.017137f
C259 VTAIL.n9 B 0.040505f
C260 VTAIL.n10 B 0.018145f
C261 VTAIL.n11 B 0.031891f
C262 VTAIL.n12 B 0.017137f
C263 VTAIL.n13 B 0.030379f
C264 VTAIL.n14 B 0.028634f
C265 VTAIL.t0 B 0.06774f
C266 VTAIL.n15 B 0.180507f
C267 VTAIL.n16 B 1.03572f
C268 VTAIL.n17 B 0.017137f
C269 VTAIL.n18 B 0.018145f
C270 VTAIL.n19 B 0.040505f
C271 VTAIL.n20 B 0.040505f
C272 VTAIL.n21 B 0.018145f
C273 VTAIL.n22 B 0.017137f
C274 VTAIL.n23 B 0.031891f
C275 VTAIL.n24 B 0.031891f
C276 VTAIL.n25 B 0.017137f
C277 VTAIL.n26 B 0.018145f
C278 VTAIL.n27 B 0.040505f
C279 VTAIL.n28 B 0.040505f
C280 VTAIL.n29 B 0.018145f
C281 VTAIL.n30 B 0.017137f
C282 VTAIL.n31 B 0.031891f
C283 VTAIL.n32 B 0.031891f
C284 VTAIL.n33 B 0.017137f
C285 VTAIL.n34 B 0.017137f
C286 VTAIL.n35 B 0.018145f
C287 VTAIL.n36 B 0.040505f
C288 VTAIL.n37 B 0.040505f
C289 VTAIL.n38 B 0.084643f
C290 VTAIL.n39 B 0.017641f
C291 VTAIL.n40 B 0.017137f
C292 VTAIL.n41 B 0.080685f
C293 VTAIL.n42 B 0.047254f
C294 VTAIL.n43 B 0.160515f
C295 VTAIL.t19 B 0.200601f
C296 VTAIL.t3 B 0.200601f
C297 VTAIL.n44 B 1.65614f
C298 VTAIL.n45 B 0.398483f
C299 VTAIL.t17 B 0.200601f
C300 VTAIL.t6 B 0.200601f
C301 VTAIL.n46 B 1.65614f
C302 VTAIL.n47 B 1.59086f
C303 VTAIL.t11 B 0.200601f
C304 VTAIL.t9 B 0.200601f
C305 VTAIL.n48 B 1.65615f
C306 VTAIL.n49 B 1.59085f
C307 VTAIL.t15 B 0.200601f
C308 VTAIL.t8 B 0.200601f
C309 VTAIL.n50 B 1.65615f
C310 VTAIL.n51 B 0.398473f
C311 VTAIL.n52 B 0.043104f
C312 VTAIL.n53 B 0.031891f
C313 VTAIL.n54 B 0.017641f
C314 VTAIL.n55 B 0.040505f
C315 VTAIL.n56 B 0.017137f
C316 VTAIL.n57 B 0.018145f
C317 VTAIL.n58 B 0.031891f
C318 VTAIL.n59 B 0.017137f
C319 VTAIL.n60 B 0.040505f
C320 VTAIL.n61 B 0.018145f
C321 VTAIL.n62 B 0.031891f
C322 VTAIL.n63 B 0.017137f
C323 VTAIL.n64 B 0.030379f
C324 VTAIL.n65 B 0.028634f
C325 VTAIL.t7 B 0.06774f
C326 VTAIL.n66 B 0.180507f
C327 VTAIL.n67 B 1.03572f
C328 VTAIL.n68 B 0.017137f
C329 VTAIL.n69 B 0.018145f
C330 VTAIL.n70 B 0.040505f
C331 VTAIL.n71 B 0.040505f
C332 VTAIL.n72 B 0.018145f
C333 VTAIL.n73 B 0.017137f
C334 VTAIL.n74 B 0.031891f
C335 VTAIL.n75 B 0.031891f
C336 VTAIL.n76 B 0.017137f
C337 VTAIL.n77 B 0.018145f
C338 VTAIL.n78 B 0.040505f
C339 VTAIL.n79 B 0.040505f
C340 VTAIL.n80 B 0.018145f
C341 VTAIL.n81 B 0.017137f
C342 VTAIL.n82 B 0.031891f
C343 VTAIL.n83 B 0.031891f
C344 VTAIL.n84 B 0.017137f
C345 VTAIL.n85 B 0.018145f
C346 VTAIL.n86 B 0.040505f
C347 VTAIL.n87 B 0.040505f
C348 VTAIL.n88 B 0.084643f
C349 VTAIL.n89 B 0.017641f
C350 VTAIL.n90 B 0.017137f
C351 VTAIL.n91 B 0.080685f
C352 VTAIL.n92 B 0.047254f
C353 VTAIL.n93 B 0.160515f
C354 VTAIL.t1 B 0.200601f
C355 VTAIL.t2 B 0.200601f
C356 VTAIL.n94 B 1.65615f
C357 VTAIL.n95 B 0.419734f
C358 VTAIL.t5 B 0.200601f
C359 VTAIL.t4 B 0.200601f
C360 VTAIL.n96 B 1.65615f
C361 VTAIL.n97 B 0.398473f
C362 VTAIL.n98 B 0.043104f
C363 VTAIL.n99 B 0.031891f
C364 VTAIL.n100 B 0.017641f
C365 VTAIL.n101 B 0.040505f
C366 VTAIL.n102 B 0.017137f
C367 VTAIL.n103 B 0.018145f
C368 VTAIL.n104 B 0.031891f
C369 VTAIL.n105 B 0.017137f
C370 VTAIL.n106 B 0.040505f
C371 VTAIL.n107 B 0.018145f
C372 VTAIL.n108 B 0.031891f
C373 VTAIL.n109 B 0.017137f
C374 VTAIL.n110 B 0.030379f
C375 VTAIL.n111 B 0.028634f
C376 VTAIL.t18 B 0.06774f
C377 VTAIL.n112 B 0.180507f
C378 VTAIL.n113 B 1.03572f
C379 VTAIL.n114 B 0.017137f
C380 VTAIL.n115 B 0.018145f
C381 VTAIL.n116 B 0.040505f
C382 VTAIL.n117 B 0.040505f
C383 VTAIL.n118 B 0.018145f
C384 VTAIL.n119 B 0.017137f
C385 VTAIL.n120 B 0.031891f
C386 VTAIL.n121 B 0.031891f
C387 VTAIL.n122 B 0.017137f
C388 VTAIL.n123 B 0.018145f
C389 VTAIL.n124 B 0.040505f
C390 VTAIL.n125 B 0.040505f
C391 VTAIL.n126 B 0.018145f
C392 VTAIL.n127 B 0.017137f
C393 VTAIL.n128 B 0.031891f
C394 VTAIL.n129 B 0.031891f
C395 VTAIL.n130 B 0.017137f
C396 VTAIL.n131 B 0.018145f
C397 VTAIL.n132 B 0.040505f
C398 VTAIL.n133 B 0.040505f
C399 VTAIL.n134 B 0.084643f
C400 VTAIL.n135 B 0.017641f
C401 VTAIL.n136 B 0.017137f
C402 VTAIL.n137 B 0.080685f
C403 VTAIL.n138 B 0.047254f
C404 VTAIL.n139 B 1.2776f
C405 VTAIL.n140 B 0.043104f
C406 VTAIL.n141 B 0.031891f
C407 VTAIL.n142 B 0.017641f
C408 VTAIL.n143 B 0.040505f
C409 VTAIL.n144 B 0.018145f
C410 VTAIL.n145 B 0.031891f
C411 VTAIL.n146 B 0.017137f
C412 VTAIL.n147 B 0.040505f
C413 VTAIL.n148 B 0.018145f
C414 VTAIL.n149 B 0.031891f
C415 VTAIL.n150 B 0.017137f
C416 VTAIL.n151 B 0.030379f
C417 VTAIL.n152 B 0.028634f
C418 VTAIL.t16 B 0.06774f
C419 VTAIL.n153 B 0.180507f
C420 VTAIL.n154 B 1.03572f
C421 VTAIL.n155 B 0.017137f
C422 VTAIL.n156 B 0.018145f
C423 VTAIL.n157 B 0.040505f
C424 VTAIL.n158 B 0.040505f
C425 VTAIL.n159 B 0.018145f
C426 VTAIL.n160 B 0.017137f
C427 VTAIL.n161 B 0.031891f
C428 VTAIL.n162 B 0.031891f
C429 VTAIL.n163 B 0.017137f
C430 VTAIL.n164 B 0.018145f
C431 VTAIL.n165 B 0.040505f
C432 VTAIL.n166 B 0.040505f
C433 VTAIL.n167 B 0.018145f
C434 VTAIL.n168 B 0.017137f
C435 VTAIL.n169 B 0.031891f
C436 VTAIL.n170 B 0.031891f
C437 VTAIL.n171 B 0.017137f
C438 VTAIL.n172 B 0.017137f
C439 VTAIL.n173 B 0.018145f
C440 VTAIL.n174 B 0.040505f
C441 VTAIL.n175 B 0.040505f
C442 VTAIL.n176 B 0.084643f
C443 VTAIL.n177 B 0.017641f
C444 VTAIL.n178 B 0.017137f
C445 VTAIL.n179 B 0.080685f
C446 VTAIL.n180 B 0.047254f
C447 VTAIL.n181 B 1.2776f
C448 VTAIL.t14 B 0.200601f
C449 VTAIL.t13 B 0.200601f
C450 VTAIL.n182 B 1.65614f
C451 VTAIL.n183 B 0.351975f
C452 VN.n0 B 0.053235f
C453 VN.t1 B 0.336971f
C454 VN.t3 B 0.336971f
C455 VN.n1 B 0.02127f
C456 VN.t5 B 0.342603f
C457 VN.t7 B 0.336971f
C458 VN.n2 B 0.14563f
C459 VN.n3 B 0.161339f
C460 VN.n4 B 0.11362f
C461 VN.n5 B 0.053235f
C462 VN.n6 B 0.163289f
C463 VN.n7 B 0.02127f
C464 VN.n8 B 0.14563f
C465 VN.t9 B 0.342603f
C466 VN.n9 B 0.161268f
C467 VN.n10 B 0.041255f
C468 VN.n11 B 0.053235f
C469 VN.t0 B 0.342603f
C470 VN.t4 B 0.336971f
C471 VN.t8 B 0.336971f
C472 VN.n12 B 0.02127f
C473 VN.t2 B 0.336971f
C474 VN.n13 B 0.14563f
C475 VN.t6 B 0.342603f
C476 VN.n14 B 0.161339f
C477 VN.n15 B 0.11362f
C478 VN.n16 B 0.053235f
C479 VN.n17 B 0.163289f
C480 VN.n18 B 0.02127f
C481 VN.n19 B 0.14563f
C482 VN.n20 B 0.161268f
C483 VN.n21 B 1.83642f
.ends

