* NGSPICE file created from diff_pair_sample_0749.ext - technology: sky130A

.subckt diff_pair_sample_0749 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X1 VTAIL.t3 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0.48015 ps=3.24 w=2.91 l=0.41
X2 VTAIL.t15 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0.48015 ps=3.24 w=2.91 l=0.41
X3 VDD1.t6 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X4 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0 ps=0 w=2.91 l=0.41
X5 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0 ps=0 w=2.91 l=0.41
X7 VDD2.t5 VN.t2 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X8 VTAIL.t5 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0.48015 ps=3.24 w=2.91 l=0.41
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0 ps=0 w=2.91 l=0.41
X10 VDD2.t4 VN.t3 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=1.1349 ps=6.6 w=2.91 l=0.41
X11 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X12 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=1.1349 ps=6.6 w=2.91 l=0.41
X13 VTAIL.t12 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0.48015 ps=3.24 w=2.91 l=0.41
X14 VDD1.t1 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=1.1349 ps=6.6 w=2.91 l=0.41
X15 VDD2.t2 VN.t5 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=1.1349 ps=6.6 w=2.91 l=0.41
X16 VTAIL.t9 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X17 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X18 VTAIL.t14 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.48015 pd=3.24 as=0.48015 ps=3.24 w=2.91 l=0.41
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1349 pd=6.6 as=0 ps=0 w=2.91 l=0.41
R0 VN.n2 VN.t4 288.433
R1 VN.n10 VN.t5 288.433
R2 VN.n1 VN.t2 267.452
R3 VN.n5 VN.t6 267.452
R4 VN.n6 VN.t3 267.452
R5 VN.n9 VN.t7 267.452
R6 VN.n13 VN.t0 267.452
R7 VN.n14 VN.t1 267.452
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.4033
R15 VN.n3 VN.n2 70.4033
R16 VN.n6 VN.n5 48.2005
R17 VN.n14 VN.n13 48.2005
R18 VN VN.n15 34.1085
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.9576
R24 VN.n2 VN.n1 20.9576
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VTAIL.n11 VTAIL.t3 73.863
R31 VTAIL.n10 VTAIL.t8 73.863
R32 VTAIL.n7 VTAIL.t15 73.863
R33 VTAIL.n15 VTAIL.t13 73.8628
R34 VTAIL.n2 VTAIL.t12 73.8628
R35 VTAIL.n3 VTAIL.t7 73.8628
R36 VTAIL.n6 VTAIL.t5 73.8628
R37 VTAIL.n14 VTAIL.t2 73.8628
R38 VTAIL.n13 VTAIL.n12 67.0589
R39 VTAIL.n9 VTAIL.n8 67.0589
R40 VTAIL.n1 VTAIL.n0 67.0587
R41 VTAIL.n5 VTAIL.n4 67.0587
R42 VTAIL.n15 VTAIL.n14 15.5134
R43 VTAIL.n7 VTAIL.n6 15.5134
R44 VTAIL.n0 VTAIL.t10 6.80462
R45 VTAIL.n0 VTAIL.t9 6.80462
R46 VTAIL.n4 VTAIL.t0 6.80462
R47 VTAIL.n4 VTAIL.t4 6.80462
R48 VTAIL.n12 VTAIL.t6 6.80462
R49 VTAIL.n12 VTAIL.t1 6.80462
R50 VTAIL.n8 VTAIL.t11 6.80462
R51 VTAIL.n8 VTAIL.t14 6.80462
R52 VTAIL.n9 VTAIL.n7 0.638431
R53 VTAIL.n10 VTAIL.n9 0.638431
R54 VTAIL.n13 VTAIL.n11 0.638431
R55 VTAIL.n14 VTAIL.n13 0.638431
R56 VTAIL.n6 VTAIL.n5 0.638431
R57 VTAIL.n5 VTAIL.n3 0.638431
R58 VTAIL.n2 VTAIL.n1 0.638431
R59 VTAIL VTAIL.n15 0.580241
R60 VTAIL.n11 VTAIL.n10 0.470328
R61 VTAIL.n3 VTAIL.n2 0.470328
R62 VTAIL VTAIL.n1 0.0586897
R63 VDD2.n2 VDD2.n1 84.0011
R64 VDD2.n2 VDD2.n0 84.0011
R65 VDD2 VDD2.n5 83.9983
R66 VDD2.n4 VDD2.n3 83.7377
R67 VDD2.n4 VDD2.n2 29.0946
R68 VDD2.n5 VDD2.t0 6.80462
R69 VDD2.n5 VDD2.t2 6.80462
R70 VDD2.n3 VDD2.t6 6.80462
R71 VDD2.n3 VDD2.t7 6.80462
R72 VDD2.n1 VDD2.t1 6.80462
R73 VDD2.n1 VDD2.t4 6.80462
R74 VDD2.n0 VDD2.t3 6.80462
R75 VDD2.n0 VDD2.t5 6.80462
R76 VDD2 VDD2.n4 0.377655
R77 B.n358 B.n357 585
R78 B.n359 B.n358 585
R79 B.n136 B.n58 585
R80 B.n135 B.n134 585
R81 B.n133 B.n132 585
R82 B.n131 B.n130 585
R83 B.n129 B.n128 585
R84 B.n127 B.n126 585
R85 B.n125 B.n124 585
R86 B.n123 B.n122 585
R87 B.n121 B.n120 585
R88 B.n119 B.n118 585
R89 B.n117 B.n116 585
R90 B.n115 B.n114 585
R91 B.n113 B.n112 585
R92 B.n111 B.n110 585
R93 B.n109 B.n108 585
R94 B.n107 B.n106 585
R95 B.n105 B.n104 585
R96 B.n103 B.n102 585
R97 B.n101 B.n100 585
R98 B.n99 B.n98 585
R99 B.n97 B.n96 585
R100 B.n95 B.n94 585
R101 B.n93 B.n92 585
R102 B.n90 B.n89 585
R103 B.n88 B.n87 585
R104 B.n86 B.n85 585
R105 B.n84 B.n83 585
R106 B.n82 B.n81 585
R107 B.n80 B.n79 585
R108 B.n78 B.n77 585
R109 B.n76 B.n75 585
R110 B.n74 B.n73 585
R111 B.n72 B.n71 585
R112 B.n70 B.n69 585
R113 B.n68 B.n67 585
R114 B.n66 B.n65 585
R115 B.n39 B.n38 585
R116 B.n362 B.n361 585
R117 B.n356 B.n59 585
R118 B.n59 B.n36 585
R119 B.n355 B.n35 585
R120 B.n366 B.n35 585
R121 B.n354 B.n34 585
R122 B.n367 B.n34 585
R123 B.n353 B.n33 585
R124 B.n368 B.n33 585
R125 B.n352 B.n351 585
R126 B.n351 B.n32 585
R127 B.n350 B.n28 585
R128 B.n374 B.n28 585
R129 B.n349 B.n27 585
R130 B.n375 B.n27 585
R131 B.n348 B.n26 585
R132 B.n376 B.n26 585
R133 B.n347 B.n346 585
R134 B.n346 B.n22 585
R135 B.n345 B.n21 585
R136 B.n382 B.n21 585
R137 B.n344 B.n20 585
R138 B.n383 B.n20 585
R139 B.n343 B.n19 585
R140 B.n384 B.n19 585
R141 B.n342 B.n341 585
R142 B.n341 B.n15 585
R143 B.n340 B.n14 585
R144 B.n390 B.n14 585
R145 B.n339 B.n13 585
R146 B.n391 B.n13 585
R147 B.n338 B.n12 585
R148 B.n392 B.n12 585
R149 B.n337 B.n336 585
R150 B.n336 B.n11 585
R151 B.n335 B.n7 585
R152 B.n398 B.n7 585
R153 B.n334 B.n6 585
R154 B.n399 B.n6 585
R155 B.n333 B.n5 585
R156 B.n400 B.n5 585
R157 B.n332 B.n331 585
R158 B.n331 B.n4 585
R159 B.n330 B.n137 585
R160 B.n330 B.n329 585
R161 B.n319 B.n138 585
R162 B.n322 B.n138 585
R163 B.n321 B.n320 585
R164 B.n323 B.n321 585
R165 B.n318 B.n142 585
R166 B.n146 B.n142 585
R167 B.n317 B.n316 585
R168 B.n316 B.n315 585
R169 B.n144 B.n143 585
R170 B.n145 B.n144 585
R171 B.n308 B.n307 585
R172 B.n309 B.n308 585
R173 B.n306 B.n151 585
R174 B.n151 B.n150 585
R175 B.n305 B.n304 585
R176 B.n304 B.n303 585
R177 B.n153 B.n152 585
R178 B.n154 B.n153 585
R179 B.n296 B.n295 585
R180 B.n297 B.n296 585
R181 B.n294 B.n159 585
R182 B.n159 B.n158 585
R183 B.n293 B.n292 585
R184 B.n292 B.n291 585
R185 B.n161 B.n160 585
R186 B.n284 B.n161 585
R187 B.n283 B.n282 585
R188 B.n285 B.n283 585
R189 B.n281 B.n166 585
R190 B.n166 B.n165 585
R191 B.n280 B.n279 585
R192 B.n279 B.n278 585
R193 B.n168 B.n167 585
R194 B.n169 B.n168 585
R195 B.n274 B.n273 585
R196 B.n172 B.n171 585
R197 B.n270 B.n269 585
R198 B.n271 B.n270 585
R199 B.n268 B.n191 585
R200 B.n267 B.n266 585
R201 B.n265 B.n264 585
R202 B.n263 B.n262 585
R203 B.n261 B.n260 585
R204 B.n259 B.n258 585
R205 B.n257 B.n256 585
R206 B.n255 B.n254 585
R207 B.n253 B.n252 585
R208 B.n251 B.n250 585
R209 B.n249 B.n248 585
R210 B.n247 B.n246 585
R211 B.n245 B.n244 585
R212 B.n243 B.n242 585
R213 B.n241 B.n240 585
R214 B.n239 B.n238 585
R215 B.n237 B.n236 585
R216 B.n235 B.n234 585
R217 B.n233 B.n232 585
R218 B.n231 B.n230 585
R219 B.n229 B.n228 585
R220 B.n226 B.n225 585
R221 B.n224 B.n223 585
R222 B.n222 B.n221 585
R223 B.n220 B.n219 585
R224 B.n218 B.n217 585
R225 B.n216 B.n215 585
R226 B.n214 B.n213 585
R227 B.n212 B.n211 585
R228 B.n210 B.n209 585
R229 B.n208 B.n207 585
R230 B.n206 B.n205 585
R231 B.n204 B.n203 585
R232 B.n202 B.n201 585
R233 B.n200 B.n199 585
R234 B.n198 B.n197 585
R235 B.n275 B.n170 585
R236 B.n170 B.n169 585
R237 B.n277 B.n276 585
R238 B.n278 B.n277 585
R239 B.n164 B.n163 585
R240 B.n165 B.n164 585
R241 B.n287 B.n286 585
R242 B.n286 B.n285 585
R243 B.n288 B.n162 585
R244 B.n284 B.n162 585
R245 B.n290 B.n289 585
R246 B.n291 B.n290 585
R247 B.n157 B.n156 585
R248 B.n158 B.n157 585
R249 B.n299 B.n298 585
R250 B.n298 B.n297 585
R251 B.n300 B.n155 585
R252 B.n155 B.n154 585
R253 B.n302 B.n301 585
R254 B.n303 B.n302 585
R255 B.n149 B.n148 585
R256 B.n150 B.n149 585
R257 B.n311 B.n310 585
R258 B.n310 B.n309 585
R259 B.n312 B.n147 585
R260 B.n147 B.n145 585
R261 B.n314 B.n313 585
R262 B.n315 B.n314 585
R263 B.n141 B.n140 585
R264 B.n146 B.n141 585
R265 B.n325 B.n324 585
R266 B.n324 B.n323 585
R267 B.n326 B.n139 585
R268 B.n322 B.n139 585
R269 B.n328 B.n327 585
R270 B.n329 B.n328 585
R271 B.n2 B.n0 585
R272 B.n4 B.n2 585
R273 B.n3 B.n1 585
R274 B.n399 B.n3 585
R275 B.n397 B.n396 585
R276 B.n398 B.n397 585
R277 B.n395 B.n8 585
R278 B.n11 B.n8 585
R279 B.n394 B.n393 585
R280 B.n393 B.n392 585
R281 B.n10 B.n9 585
R282 B.n391 B.n10 585
R283 B.n389 B.n388 585
R284 B.n390 B.n389 585
R285 B.n387 B.n16 585
R286 B.n16 B.n15 585
R287 B.n386 B.n385 585
R288 B.n385 B.n384 585
R289 B.n18 B.n17 585
R290 B.n383 B.n18 585
R291 B.n381 B.n380 585
R292 B.n382 B.n381 585
R293 B.n379 B.n23 585
R294 B.n23 B.n22 585
R295 B.n378 B.n377 585
R296 B.n377 B.n376 585
R297 B.n25 B.n24 585
R298 B.n375 B.n25 585
R299 B.n373 B.n372 585
R300 B.n374 B.n373 585
R301 B.n371 B.n29 585
R302 B.n32 B.n29 585
R303 B.n370 B.n369 585
R304 B.n369 B.n368 585
R305 B.n31 B.n30 585
R306 B.n367 B.n31 585
R307 B.n365 B.n364 585
R308 B.n366 B.n365 585
R309 B.n363 B.n37 585
R310 B.n37 B.n36 585
R311 B.n402 B.n401 585
R312 B.n401 B.n400 585
R313 B.n273 B.n170 526.135
R314 B.n361 B.n37 526.135
R315 B.n197 B.n168 526.135
R316 B.n358 B.n59 526.135
R317 B.n195 B.t16 380.104
R318 B.n192 B.t8 380.104
R319 B.n63 B.t19 380.104
R320 B.n60 B.t12 380.104
R321 B.n359 B.n57 256.663
R322 B.n359 B.n56 256.663
R323 B.n359 B.n55 256.663
R324 B.n359 B.n54 256.663
R325 B.n359 B.n53 256.663
R326 B.n359 B.n52 256.663
R327 B.n359 B.n51 256.663
R328 B.n359 B.n50 256.663
R329 B.n359 B.n49 256.663
R330 B.n359 B.n48 256.663
R331 B.n359 B.n47 256.663
R332 B.n359 B.n46 256.663
R333 B.n359 B.n45 256.663
R334 B.n359 B.n44 256.663
R335 B.n359 B.n43 256.663
R336 B.n359 B.n42 256.663
R337 B.n359 B.n41 256.663
R338 B.n359 B.n40 256.663
R339 B.n360 B.n359 256.663
R340 B.n272 B.n271 256.663
R341 B.n271 B.n173 256.663
R342 B.n271 B.n174 256.663
R343 B.n271 B.n175 256.663
R344 B.n271 B.n176 256.663
R345 B.n271 B.n177 256.663
R346 B.n271 B.n178 256.663
R347 B.n271 B.n179 256.663
R348 B.n271 B.n180 256.663
R349 B.n271 B.n181 256.663
R350 B.n271 B.n182 256.663
R351 B.n271 B.n183 256.663
R352 B.n271 B.n184 256.663
R353 B.n271 B.n185 256.663
R354 B.n271 B.n186 256.663
R355 B.n271 B.n187 256.663
R356 B.n271 B.n188 256.663
R357 B.n271 B.n189 256.663
R358 B.n271 B.n190 256.663
R359 B.n271 B.n169 165.303
R360 B.n359 B.n36 165.303
R361 B.n277 B.n170 163.367
R362 B.n277 B.n164 163.367
R363 B.n286 B.n164 163.367
R364 B.n286 B.n162 163.367
R365 B.n290 B.n162 163.367
R366 B.n290 B.n157 163.367
R367 B.n298 B.n157 163.367
R368 B.n298 B.n155 163.367
R369 B.n302 B.n155 163.367
R370 B.n302 B.n149 163.367
R371 B.n310 B.n149 163.367
R372 B.n310 B.n147 163.367
R373 B.n314 B.n147 163.367
R374 B.n314 B.n141 163.367
R375 B.n324 B.n141 163.367
R376 B.n324 B.n139 163.367
R377 B.n328 B.n139 163.367
R378 B.n328 B.n2 163.367
R379 B.n401 B.n2 163.367
R380 B.n401 B.n3 163.367
R381 B.n397 B.n3 163.367
R382 B.n397 B.n8 163.367
R383 B.n393 B.n8 163.367
R384 B.n393 B.n10 163.367
R385 B.n389 B.n10 163.367
R386 B.n389 B.n16 163.367
R387 B.n385 B.n16 163.367
R388 B.n385 B.n18 163.367
R389 B.n381 B.n18 163.367
R390 B.n381 B.n23 163.367
R391 B.n377 B.n23 163.367
R392 B.n377 B.n25 163.367
R393 B.n373 B.n25 163.367
R394 B.n373 B.n29 163.367
R395 B.n369 B.n29 163.367
R396 B.n369 B.n31 163.367
R397 B.n365 B.n31 163.367
R398 B.n365 B.n37 163.367
R399 B.n270 B.n172 163.367
R400 B.n270 B.n191 163.367
R401 B.n266 B.n265 163.367
R402 B.n262 B.n261 163.367
R403 B.n258 B.n257 163.367
R404 B.n254 B.n253 163.367
R405 B.n250 B.n249 163.367
R406 B.n246 B.n245 163.367
R407 B.n242 B.n241 163.367
R408 B.n238 B.n237 163.367
R409 B.n234 B.n233 163.367
R410 B.n230 B.n229 163.367
R411 B.n225 B.n224 163.367
R412 B.n221 B.n220 163.367
R413 B.n217 B.n216 163.367
R414 B.n213 B.n212 163.367
R415 B.n209 B.n208 163.367
R416 B.n205 B.n204 163.367
R417 B.n201 B.n200 163.367
R418 B.n279 B.n168 163.367
R419 B.n279 B.n166 163.367
R420 B.n283 B.n166 163.367
R421 B.n283 B.n161 163.367
R422 B.n292 B.n161 163.367
R423 B.n292 B.n159 163.367
R424 B.n296 B.n159 163.367
R425 B.n296 B.n153 163.367
R426 B.n304 B.n153 163.367
R427 B.n304 B.n151 163.367
R428 B.n308 B.n151 163.367
R429 B.n308 B.n144 163.367
R430 B.n316 B.n144 163.367
R431 B.n316 B.n142 163.367
R432 B.n321 B.n142 163.367
R433 B.n321 B.n138 163.367
R434 B.n330 B.n138 163.367
R435 B.n331 B.n330 163.367
R436 B.n331 B.n5 163.367
R437 B.n6 B.n5 163.367
R438 B.n7 B.n6 163.367
R439 B.n336 B.n7 163.367
R440 B.n336 B.n12 163.367
R441 B.n13 B.n12 163.367
R442 B.n14 B.n13 163.367
R443 B.n341 B.n14 163.367
R444 B.n341 B.n19 163.367
R445 B.n20 B.n19 163.367
R446 B.n21 B.n20 163.367
R447 B.n346 B.n21 163.367
R448 B.n346 B.n26 163.367
R449 B.n27 B.n26 163.367
R450 B.n28 B.n27 163.367
R451 B.n351 B.n28 163.367
R452 B.n351 B.n33 163.367
R453 B.n34 B.n33 163.367
R454 B.n35 B.n34 163.367
R455 B.n59 B.n35 163.367
R456 B.n65 B.n39 163.367
R457 B.n69 B.n68 163.367
R458 B.n73 B.n72 163.367
R459 B.n77 B.n76 163.367
R460 B.n81 B.n80 163.367
R461 B.n85 B.n84 163.367
R462 B.n89 B.n88 163.367
R463 B.n94 B.n93 163.367
R464 B.n98 B.n97 163.367
R465 B.n102 B.n101 163.367
R466 B.n106 B.n105 163.367
R467 B.n110 B.n109 163.367
R468 B.n114 B.n113 163.367
R469 B.n118 B.n117 163.367
R470 B.n122 B.n121 163.367
R471 B.n126 B.n125 163.367
R472 B.n130 B.n129 163.367
R473 B.n134 B.n133 163.367
R474 B.n358 B.n58 163.367
R475 B.n195 B.t18 93.425
R476 B.n60 B.t14 93.425
R477 B.n192 B.t11 93.4232
R478 B.n63 B.t20 93.4232
R479 B.n278 B.n169 91.3872
R480 B.n278 B.n165 91.3872
R481 B.n285 B.n165 91.3872
R482 B.n285 B.n284 91.3872
R483 B.n291 B.n158 91.3872
R484 B.n297 B.n158 91.3872
R485 B.n297 B.n154 91.3872
R486 B.n303 B.n154 91.3872
R487 B.n309 B.n150 91.3872
R488 B.n315 B.n145 91.3872
R489 B.n315 B.n146 91.3872
R490 B.n323 B.n322 91.3872
R491 B.n329 B.n4 91.3872
R492 B.n400 B.n4 91.3872
R493 B.n400 B.n399 91.3872
R494 B.n399 B.n398 91.3872
R495 B.n392 B.n11 91.3872
R496 B.n391 B.n390 91.3872
R497 B.n390 B.n15 91.3872
R498 B.n384 B.n383 91.3872
R499 B.n382 B.n22 91.3872
R500 B.n376 B.n22 91.3872
R501 B.n376 B.n375 91.3872
R502 B.n375 B.n374 91.3872
R503 B.n368 B.n32 91.3872
R504 B.n368 B.n367 91.3872
R505 B.n367 B.n366 91.3872
R506 B.n366 B.n36 91.3872
R507 B.n309 B.t0 87.3554
R508 B.n384 B.t1 87.3554
R509 B.n323 B.t4 79.2919
R510 B.n392 B.t6 79.2919
R511 B.n196 B.t17 79.0735
R512 B.n61 B.t15 79.0735
R513 B.n193 B.t10 79.0717
R514 B.n64 B.t21 79.0717
R515 B.n273 B.n272 71.676
R516 B.n191 B.n173 71.676
R517 B.n265 B.n174 71.676
R518 B.n261 B.n175 71.676
R519 B.n257 B.n176 71.676
R520 B.n253 B.n177 71.676
R521 B.n249 B.n178 71.676
R522 B.n245 B.n179 71.676
R523 B.n241 B.n180 71.676
R524 B.n237 B.n181 71.676
R525 B.n233 B.n182 71.676
R526 B.n229 B.n183 71.676
R527 B.n224 B.n184 71.676
R528 B.n220 B.n185 71.676
R529 B.n216 B.n186 71.676
R530 B.n212 B.n187 71.676
R531 B.n208 B.n188 71.676
R532 B.n204 B.n189 71.676
R533 B.n200 B.n190 71.676
R534 B.n361 B.n360 71.676
R535 B.n65 B.n40 71.676
R536 B.n69 B.n41 71.676
R537 B.n73 B.n42 71.676
R538 B.n77 B.n43 71.676
R539 B.n81 B.n44 71.676
R540 B.n85 B.n45 71.676
R541 B.n89 B.n46 71.676
R542 B.n94 B.n47 71.676
R543 B.n98 B.n48 71.676
R544 B.n102 B.n49 71.676
R545 B.n106 B.n50 71.676
R546 B.n110 B.n51 71.676
R547 B.n114 B.n52 71.676
R548 B.n118 B.n53 71.676
R549 B.n122 B.n54 71.676
R550 B.n126 B.n55 71.676
R551 B.n130 B.n56 71.676
R552 B.n134 B.n57 71.676
R553 B.n58 B.n57 71.676
R554 B.n133 B.n56 71.676
R555 B.n129 B.n55 71.676
R556 B.n125 B.n54 71.676
R557 B.n121 B.n53 71.676
R558 B.n117 B.n52 71.676
R559 B.n113 B.n51 71.676
R560 B.n109 B.n50 71.676
R561 B.n105 B.n49 71.676
R562 B.n101 B.n48 71.676
R563 B.n97 B.n47 71.676
R564 B.n93 B.n46 71.676
R565 B.n88 B.n45 71.676
R566 B.n84 B.n44 71.676
R567 B.n80 B.n43 71.676
R568 B.n76 B.n42 71.676
R569 B.n72 B.n41 71.676
R570 B.n68 B.n40 71.676
R571 B.n360 B.n39 71.676
R572 B.n272 B.n172 71.676
R573 B.n266 B.n173 71.676
R574 B.n262 B.n174 71.676
R575 B.n258 B.n175 71.676
R576 B.n254 B.n176 71.676
R577 B.n250 B.n177 71.676
R578 B.n246 B.n178 71.676
R579 B.n242 B.n179 71.676
R580 B.n238 B.n180 71.676
R581 B.n234 B.n181 71.676
R582 B.n230 B.n182 71.676
R583 B.n225 B.n183 71.676
R584 B.n221 B.n184 71.676
R585 B.n217 B.n185 71.676
R586 B.n213 B.n186 71.676
R587 B.n209 B.n187 71.676
R588 B.n205 B.n188 71.676
R589 B.n201 B.n189 71.676
R590 B.n197 B.n190 71.676
R591 B.n303 B.t5 71.2284
R592 B.t2 B.n382 71.2284
R593 B.n329 B.t7 63.1648
R594 B.n398 B.t3 63.1648
R595 B.n227 B.n196 59.5399
R596 B.n194 B.n193 59.5399
R597 B.n91 B.n64 59.5399
R598 B.n62 B.n61 59.5399
R599 B.n291 B.t9 55.1013
R600 B.n374 B.t13 55.1013
R601 B.n284 B.t9 36.2864
R602 B.n32 B.t13 36.2864
R603 B.n363 B.n362 34.1859
R604 B.n357 B.n356 34.1859
R605 B.n198 B.n167 34.1859
R606 B.n275 B.n274 34.1859
R607 B.n322 B.t7 28.2229
R608 B.n11 B.t3 28.2229
R609 B.t5 B.n150 20.1593
R610 B.n383 B.t2 20.1593
R611 B B.n402 18.0485
R612 B.n196 B.n195 14.352
R613 B.n193 B.n192 14.352
R614 B.n64 B.n63 14.352
R615 B.n61 B.n60 14.352
R616 B.n146 B.t4 12.0958
R617 B.t6 B.n391 12.0958
R618 B.n362 B.n38 10.6151
R619 B.n66 B.n38 10.6151
R620 B.n67 B.n66 10.6151
R621 B.n70 B.n67 10.6151
R622 B.n71 B.n70 10.6151
R623 B.n74 B.n71 10.6151
R624 B.n75 B.n74 10.6151
R625 B.n78 B.n75 10.6151
R626 B.n79 B.n78 10.6151
R627 B.n82 B.n79 10.6151
R628 B.n83 B.n82 10.6151
R629 B.n86 B.n83 10.6151
R630 B.n87 B.n86 10.6151
R631 B.n90 B.n87 10.6151
R632 B.n95 B.n92 10.6151
R633 B.n96 B.n95 10.6151
R634 B.n99 B.n96 10.6151
R635 B.n100 B.n99 10.6151
R636 B.n103 B.n100 10.6151
R637 B.n104 B.n103 10.6151
R638 B.n107 B.n104 10.6151
R639 B.n108 B.n107 10.6151
R640 B.n112 B.n111 10.6151
R641 B.n115 B.n112 10.6151
R642 B.n116 B.n115 10.6151
R643 B.n119 B.n116 10.6151
R644 B.n120 B.n119 10.6151
R645 B.n123 B.n120 10.6151
R646 B.n124 B.n123 10.6151
R647 B.n127 B.n124 10.6151
R648 B.n128 B.n127 10.6151
R649 B.n131 B.n128 10.6151
R650 B.n132 B.n131 10.6151
R651 B.n135 B.n132 10.6151
R652 B.n136 B.n135 10.6151
R653 B.n357 B.n136 10.6151
R654 B.n280 B.n167 10.6151
R655 B.n281 B.n280 10.6151
R656 B.n282 B.n281 10.6151
R657 B.n282 B.n160 10.6151
R658 B.n293 B.n160 10.6151
R659 B.n294 B.n293 10.6151
R660 B.n295 B.n294 10.6151
R661 B.n295 B.n152 10.6151
R662 B.n305 B.n152 10.6151
R663 B.n306 B.n305 10.6151
R664 B.n307 B.n306 10.6151
R665 B.n307 B.n143 10.6151
R666 B.n317 B.n143 10.6151
R667 B.n318 B.n317 10.6151
R668 B.n320 B.n318 10.6151
R669 B.n320 B.n319 10.6151
R670 B.n319 B.n137 10.6151
R671 B.n332 B.n137 10.6151
R672 B.n333 B.n332 10.6151
R673 B.n334 B.n333 10.6151
R674 B.n335 B.n334 10.6151
R675 B.n337 B.n335 10.6151
R676 B.n338 B.n337 10.6151
R677 B.n339 B.n338 10.6151
R678 B.n340 B.n339 10.6151
R679 B.n342 B.n340 10.6151
R680 B.n343 B.n342 10.6151
R681 B.n344 B.n343 10.6151
R682 B.n345 B.n344 10.6151
R683 B.n347 B.n345 10.6151
R684 B.n348 B.n347 10.6151
R685 B.n349 B.n348 10.6151
R686 B.n350 B.n349 10.6151
R687 B.n352 B.n350 10.6151
R688 B.n353 B.n352 10.6151
R689 B.n354 B.n353 10.6151
R690 B.n355 B.n354 10.6151
R691 B.n356 B.n355 10.6151
R692 B.n274 B.n171 10.6151
R693 B.n269 B.n171 10.6151
R694 B.n269 B.n268 10.6151
R695 B.n268 B.n267 10.6151
R696 B.n267 B.n264 10.6151
R697 B.n264 B.n263 10.6151
R698 B.n263 B.n260 10.6151
R699 B.n260 B.n259 10.6151
R700 B.n259 B.n256 10.6151
R701 B.n256 B.n255 10.6151
R702 B.n255 B.n252 10.6151
R703 B.n252 B.n251 10.6151
R704 B.n251 B.n248 10.6151
R705 B.n248 B.n247 10.6151
R706 B.n244 B.n243 10.6151
R707 B.n243 B.n240 10.6151
R708 B.n240 B.n239 10.6151
R709 B.n239 B.n236 10.6151
R710 B.n236 B.n235 10.6151
R711 B.n235 B.n232 10.6151
R712 B.n232 B.n231 10.6151
R713 B.n231 B.n228 10.6151
R714 B.n226 B.n223 10.6151
R715 B.n223 B.n222 10.6151
R716 B.n222 B.n219 10.6151
R717 B.n219 B.n218 10.6151
R718 B.n218 B.n215 10.6151
R719 B.n215 B.n214 10.6151
R720 B.n214 B.n211 10.6151
R721 B.n211 B.n210 10.6151
R722 B.n210 B.n207 10.6151
R723 B.n207 B.n206 10.6151
R724 B.n206 B.n203 10.6151
R725 B.n203 B.n202 10.6151
R726 B.n202 B.n199 10.6151
R727 B.n199 B.n198 10.6151
R728 B.n276 B.n275 10.6151
R729 B.n276 B.n163 10.6151
R730 B.n287 B.n163 10.6151
R731 B.n288 B.n287 10.6151
R732 B.n289 B.n288 10.6151
R733 B.n289 B.n156 10.6151
R734 B.n299 B.n156 10.6151
R735 B.n300 B.n299 10.6151
R736 B.n301 B.n300 10.6151
R737 B.n301 B.n148 10.6151
R738 B.n311 B.n148 10.6151
R739 B.n312 B.n311 10.6151
R740 B.n313 B.n312 10.6151
R741 B.n313 B.n140 10.6151
R742 B.n325 B.n140 10.6151
R743 B.n326 B.n325 10.6151
R744 B.n327 B.n326 10.6151
R745 B.n327 B.n0 10.6151
R746 B.n396 B.n1 10.6151
R747 B.n396 B.n395 10.6151
R748 B.n395 B.n394 10.6151
R749 B.n394 B.n9 10.6151
R750 B.n388 B.n9 10.6151
R751 B.n388 B.n387 10.6151
R752 B.n387 B.n386 10.6151
R753 B.n386 B.n17 10.6151
R754 B.n380 B.n17 10.6151
R755 B.n380 B.n379 10.6151
R756 B.n379 B.n378 10.6151
R757 B.n378 B.n24 10.6151
R758 B.n372 B.n24 10.6151
R759 B.n372 B.n371 10.6151
R760 B.n371 B.n370 10.6151
R761 B.n370 B.n30 10.6151
R762 B.n364 B.n30 10.6151
R763 B.n364 B.n363 10.6151
R764 B.n92 B.n91 6.5566
R765 B.n108 B.n62 6.5566
R766 B.n244 B.n194 6.5566
R767 B.n228 B.n227 6.5566
R768 B.n91 B.n90 4.05904
R769 B.n111 B.n62 4.05904
R770 B.n247 B.n194 4.05904
R771 B.n227 B.n226 4.05904
R772 B.t0 B.n145 4.03227
R773 B.t1 B.n15 4.03227
R774 B.n402 B.n0 2.81026
R775 B.n402 B.n1 2.81026
R776 VP.n4 VP.t0 288.433
R777 VP.n10 VP.t3 267.452
R778 VP.n1 VP.t7 267.452
R779 VP.n15 VP.t2 267.452
R780 VP.n16 VP.t6 267.452
R781 VP.n8 VP.t5 267.452
R782 VP.n7 VP.t4 267.452
R783 VP.n3 VP.t1 267.452
R784 VP.n17 VP.n16 161.3
R785 VP.n6 VP.n5 161.3
R786 VP.n7 VP.n2 161.3
R787 VP.n9 VP.n8 161.3
R788 VP.n15 VP.n0 161.3
R789 VP.n14 VP.n13 161.3
R790 VP.n12 VP.n1 161.3
R791 VP.n11 VP.n10 161.3
R792 VP.n5 VP.n4 70.4033
R793 VP.n10 VP.n1 48.2005
R794 VP.n16 VP.n15 48.2005
R795 VP.n8 VP.n7 48.2005
R796 VP.n11 VP.n9 33.7278
R797 VP.n14 VP.n1 24.1005
R798 VP.n15 VP.n14 24.1005
R799 VP.n6 VP.n3 24.1005
R800 VP.n7 VP.n6 24.1005
R801 VP.n4 VP.n3 20.9576
R802 VP.n5 VP.n2 0.189894
R803 VP.n9 VP.n2 0.189894
R804 VP.n12 VP.n11 0.189894
R805 VP.n13 VP.n12 0.189894
R806 VP.n13 VP.n0 0.189894
R807 VP.n17 VP.n0 0.189894
R808 VP VP.n17 0.0516364
R809 VDD1 VDD1.n0 84.1148
R810 VDD1.n3 VDD1.n2 84.0011
R811 VDD1.n3 VDD1.n1 84.0011
R812 VDD1.n5 VDD1.n4 83.7376
R813 VDD1.n5 VDD1.n3 29.6776
R814 VDD1.n4 VDD1.t3 6.80462
R815 VDD1.n4 VDD1.t2 6.80462
R816 VDD1.n0 VDD1.t7 6.80462
R817 VDD1.n0 VDD1.t6 6.80462
R818 VDD1.n2 VDD1.t5 6.80462
R819 VDD1.n2 VDD1.t1 6.80462
R820 VDD1.n1 VDD1.t4 6.80462
R821 VDD1.n1 VDD1.t0 6.80462
R822 VDD1 VDD1.n5 0.261276
C0 VDD2 VN 1.25477f
C1 VDD1 VN 0.15282f
C2 VP VN 3.31102f
C3 VDD2 VTAIL 4.89195f
C4 VDD1 VTAIL 4.85222f
C5 VTAIL VP 1.35156f
C6 VTAIL VN 1.33746f
C7 VDD2 VDD1 0.68501f
C8 VDD2 VP 0.292185f
C9 VDD1 VP 1.39333f
C10 VDD2 B 2.398495f
C11 VDD1 B 2.59672f
C12 VTAIL B 3.444218f
C13 VN B 5.71197f
C14 VP B 4.762352f
C15 VDD1.t7 B 0.051753f
C16 VDD1.t6 B 0.051753f
C17 VDD1.n0 B 0.381487f
C18 VDD1.t4 B 0.051753f
C19 VDD1.t0 B 0.051753f
C20 VDD1.n1 B 0.381127f
C21 VDD1.t5 B 0.051753f
C22 VDD1.t1 B 0.051753f
C23 VDD1.n2 B 0.381127f
C24 VDD1.n3 B 1.34006f
C25 VDD1.t3 B 0.051753f
C26 VDD1.t2 B 0.051753f
C27 VDD1.n4 B 0.380355f
C28 VDD1.n5 B 1.32467f
C29 VP.n0 B 0.029467f
C30 VP.t7 B 0.105749f
C31 VP.n1 B 0.068484f
C32 VP.n2 B 0.029467f
C33 VP.t5 B 0.105749f
C34 VP.t4 B 0.105749f
C35 VP.t1 B 0.105749f
C36 VP.n3 B 0.068484f
C37 VP.t0 B 0.110515f
C38 VP.n4 B 0.060922f
C39 VP.n5 B 0.09056f
C40 VP.n6 B 0.006687f
C41 VP.n7 B 0.068484f
C42 VP.n8 B 0.065486f
C43 VP.n9 B 0.816448f
C44 VP.t3 B 0.105749f
C45 VP.n10 B 0.065486f
C46 VP.n11 B 0.847854f
C47 VP.n12 B 0.029467f
C48 VP.n13 B 0.029467f
C49 VP.n14 B 0.006687f
C50 VP.t2 B 0.105749f
C51 VP.n15 B 0.068484f
C52 VP.t6 B 0.105749f
C53 VP.n16 B 0.065486f
C54 VP.n17 B 0.022836f
C55 VDD2.t3 B 0.052646f
C56 VDD2.t5 B 0.052646f
C57 VDD2.n0 B 0.387704f
C58 VDD2.t1 B 0.052646f
C59 VDD2.t4 B 0.052646f
C60 VDD2.n1 B 0.387704f
C61 VDD2.n2 B 1.3139f
C62 VDD2.t6 B 0.052646f
C63 VDD2.t7 B 0.052646f
C64 VDD2.n3 B 0.38692f
C65 VDD2.n4 B 1.32085f
C66 VDD2.t0 B 0.052646f
C67 VDD2.t2 B 0.052646f
C68 VDD2.n5 B 0.387688f
C69 VTAIL.t10 B 0.047028f
C70 VTAIL.t9 B 0.047028f
C71 VTAIL.n0 B 0.308327f
C72 VTAIL.n1 B 0.209267f
C73 VTAIL.t12 B 0.4007f
C74 VTAIL.n2 B 0.272278f
C75 VTAIL.t7 B 0.4007f
C76 VTAIL.n3 B 0.272278f
C77 VTAIL.t0 B 0.047028f
C78 VTAIL.t4 B 0.047028f
C79 VTAIL.n4 B 0.308327f
C80 VTAIL.n5 B 0.24747f
C81 VTAIL.t5 B 0.4007f
C82 VTAIL.n6 B 0.726468f
C83 VTAIL.t15 B 0.400702f
C84 VTAIL.n7 B 0.726466f
C85 VTAIL.t11 B 0.047028f
C86 VTAIL.t14 B 0.047028f
C87 VTAIL.n8 B 0.308329f
C88 VTAIL.n9 B 0.247469f
C89 VTAIL.t8 B 0.400702f
C90 VTAIL.n10 B 0.272277f
C91 VTAIL.t3 B 0.400702f
C92 VTAIL.n11 B 0.272277f
C93 VTAIL.t6 B 0.047028f
C94 VTAIL.t1 B 0.047028f
C95 VTAIL.n12 B 0.308329f
C96 VTAIL.n13 B 0.247469f
C97 VTAIL.t2 B 0.4007f
C98 VTAIL.n14 B 0.726467f
C99 VTAIL.t13 B 0.4007f
C100 VTAIL.n15 B 0.722633f
C101 VN.n0 B 0.029101f
C102 VN.t2 B 0.104438f
C103 VN.n1 B 0.067635f
C104 VN.t4 B 0.109145f
C105 VN.n2 B 0.060166f
C106 VN.n3 B 0.089437f
C107 VN.n4 B 0.006604f
C108 VN.t6 B 0.104438f
C109 VN.n5 B 0.067635f
C110 VN.t3 B 0.104438f
C111 VN.n6 B 0.064674f
C112 VN.n7 B 0.022552f
C113 VN.n8 B 0.029101f
C114 VN.t7 B 0.104438f
C115 VN.n9 B 0.067635f
C116 VN.t5 B 0.109145f
C117 VN.n10 B 0.060166f
C118 VN.n11 B 0.089437f
C119 VN.n12 B 0.006604f
C120 VN.t0 B 0.104438f
C121 VN.n13 B 0.067635f
C122 VN.t1 B 0.104438f
C123 VN.n14 B 0.064674f
C124 VN.n15 B 0.825725f
.ends

