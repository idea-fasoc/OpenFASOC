* NGSPICE file created from diff_pair_sample_0697.ext - technology: sky130A

.subckt diff_pair_sample_0697 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=0.81
X1 VDD2.t9 VN.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=0.81
X2 VDD2.t8 VN.t1 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=0.81
X3 VTAIL.t1 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X4 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=0.81
X5 VDD2.t7 VN.t2 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X6 VDD1.t8 VP.t1 VTAIL.t19 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X7 VDD1.t7 VP.t2 VTAIL.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=0.81
X8 VTAIL.t8 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X9 VTAIL.t7 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=0.81
X11 VDD2.t6 VN.t3 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=0.81
X12 VTAIL.t18 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X13 VTAIL.t3 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X14 VDD1.t3 VP.t6 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=0.81
X15 VDD2.t4 VN.t5 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=0.81
X16 VDD1.t2 VP.t7 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=7.761 ps=40.58 w=19.9 l=0.81
X17 VTAIL.t16 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X18 VDD2.t2 VN.t7 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=0 ps=0 w=19.9 l=0.81
X20 VTAIL.t15 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X21 VDD1.t1 VP.t8 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.761 pd=40.58 as=3.2835 ps=20.23 w=19.9 l=0.81
X22 VDD1.t0 VP.t9 VTAIL.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
X23 VTAIL.t9 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2835 pd=20.23 as=3.2835 ps=20.23 w=19.9 l=0.81
R0 B.n491 B.t10 793.883
R1 B.n497 B.t18 793.883
R2 B.n128 B.t14 793.883
R3 B.n125 B.t21 793.883
R4 B.n932 B.n931 585
R5 B.n933 B.n932 585
R6 B.n403 B.n124 585
R7 B.n402 B.n401 585
R8 B.n400 B.n399 585
R9 B.n398 B.n397 585
R10 B.n396 B.n395 585
R11 B.n394 B.n393 585
R12 B.n392 B.n391 585
R13 B.n390 B.n389 585
R14 B.n388 B.n387 585
R15 B.n386 B.n385 585
R16 B.n384 B.n383 585
R17 B.n382 B.n381 585
R18 B.n380 B.n379 585
R19 B.n378 B.n377 585
R20 B.n376 B.n375 585
R21 B.n374 B.n373 585
R22 B.n372 B.n371 585
R23 B.n370 B.n369 585
R24 B.n368 B.n367 585
R25 B.n366 B.n365 585
R26 B.n364 B.n363 585
R27 B.n362 B.n361 585
R28 B.n360 B.n359 585
R29 B.n358 B.n357 585
R30 B.n356 B.n355 585
R31 B.n354 B.n353 585
R32 B.n352 B.n351 585
R33 B.n350 B.n349 585
R34 B.n348 B.n347 585
R35 B.n346 B.n345 585
R36 B.n344 B.n343 585
R37 B.n342 B.n341 585
R38 B.n340 B.n339 585
R39 B.n338 B.n337 585
R40 B.n336 B.n335 585
R41 B.n334 B.n333 585
R42 B.n332 B.n331 585
R43 B.n330 B.n329 585
R44 B.n328 B.n327 585
R45 B.n326 B.n325 585
R46 B.n324 B.n323 585
R47 B.n322 B.n321 585
R48 B.n320 B.n319 585
R49 B.n318 B.n317 585
R50 B.n316 B.n315 585
R51 B.n314 B.n313 585
R52 B.n312 B.n311 585
R53 B.n310 B.n309 585
R54 B.n308 B.n307 585
R55 B.n306 B.n305 585
R56 B.n304 B.n303 585
R57 B.n302 B.n301 585
R58 B.n300 B.n299 585
R59 B.n298 B.n297 585
R60 B.n296 B.n295 585
R61 B.n294 B.n293 585
R62 B.n292 B.n291 585
R63 B.n290 B.n289 585
R64 B.n288 B.n287 585
R65 B.n286 B.n285 585
R66 B.n284 B.n283 585
R67 B.n282 B.n281 585
R68 B.n280 B.n279 585
R69 B.n278 B.n277 585
R70 B.n276 B.n275 585
R71 B.n274 B.n273 585
R72 B.n272 B.n271 585
R73 B.n270 B.n269 585
R74 B.n268 B.n267 585
R75 B.n266 B.n265 585
R76 B.n264 B.n263 585
R77 B.n262 B.n261 585
R78 B.n260 B.n259 585
R79 B.n257 B.n256 585
R80 B.n255 B.n254 585
R81 B.n253 B.n252 585
R82 B.n251 B.n250 585
R83 B.n249 B.n248 585
R84 B.n247 B.n246 585
R85 B.n245 B.n244 585
R86 B.n243 B.n242 585
R87 B.n241 B.n240 585
R88 B.n239 B.n238 585
R89 B.n237 B.n236 585
R90 B.n235 B.n234 585
R91 B.n233 B.n232 585
R92 B.n231 B.n230 585
R93 B.n229 B.n228 585
R94 B.n227 B.n226 585
R95 B.n225 B.n224 585
R96 B.n223 B.n222 585
R97 B.n221 B.n220 585
R98 B.n219 B.n218 585
R99 B.n217 B.n216 585
R100 B.n215 B.n214 585
R101 B.n213 B.n212 585
R102 B.n211 B.n210 585
R103 B.n209 B.n208 585
R104 B.n207 B.n206 585
R105 B.n205 B.n204 585
R106 B.n203 B.n202 585
R107 B.n201 B.n200 585
R108 B.n199 B.n198 585
R109 B.n197 B.n196 585
R110 B.n195 B.n194 585
R111 B.n193 B.n192 585
R112 B.n191 B.n190 585
R113 B.n189 B.n188 585
R114 B.n187 B.n186 585
R115 B.n185 B.n184 585
R116 B.n183 B.n182 585
R117 B.n181 B.n180 585
R118 B.n179 B.n178 585
R119 B.n177 B.n176 585
R120 B.n175 B.n174 585
R121 B.n173 B.n172 585
R122 B.n171 B.n170 585
R123 B.n169 B.n168 585
R124 B.n167 B.n166 585
R125 B.n165 B.n164 585
R126 B.n163 B.n162 585
R127 B.n161 B.n160 585
R128 B.n159 B.n158 585
R129 B.n157 B.n156 585
R130 B.n155 B.n154 585
R131 B.n153 B.n152 585
R132 B.n151 B.n150 585
R133 B.n149 B.n148 585
R134 B.n147 B.n146 585
R135 B.n145 B.n144 585
R136 B.n143 B.n142 585
R137 B.n141 B.n140 585
R138 B.n139 B.n138 585
R139 B.n137 B.n136 585
R140 B.n135 B.n134 585
R141 B.n133 B.n132 585
R142 B.n131 B.n130 585
R143 B.n53 B.n52 585
R144 B.n930 B.n54 585
R145 B.n934 B.n54 585
R146 B.n929 B.n928 585
R147 B.n928 B.n50 585
R148 B.n927 B.n49 585
R149 B.n940 B.n49 585
R150 B.n926 B.n48 585
R151 B.n941 B.n48 585
R152 B.n925 B.n47 585
R153 B.n942 B.n47 585
R154 B.n924 B.n923 585
R155 B.n923 B.n43 585
R156 B.n922 B.n42 585
R157 B.n948 B.n42 585
R158 B.n921 B.n41 585
R159 B.n949 B.n41 585
R160 B.n920 B.n40 585
R161 B.n950 B.n40 585
R162 B.n919 B.n918 585
R163 B.n918 B.n36 585
R164 B.n917 B.n35 585
R165 B.n956 B.n35 585
R166 B.n916 B.n34 585
R167 B.n957 B.n34 585
R168 B.n915 B.n33 585
R169 B.n958 B.n33 585
R170 B.n914 B.n913 585
R171 B.n913 B.n29 585
R172 B.n912 B.n28 585
R173 B.n964 B.n28 585
R174 B.n911 B.n27 585
R175 B.n965 B.n27 585
R176 B.n910 B.n26 585
R177 B.n966 B.n26 585
R178 B.n909 B.n908 585
R179 B.n908 B.n22 585
R180 B.n907 B.n21 585
R181 B.n972 B.n21 585
R182 B.n906 B.n20 585
R183 B.n973 B.n20 585
R184 B.n905 B.n19 585
R185 B.n974 B.n19 585
R186 B.n904 B.n903 585
R187 B.n903 B.n18 585
R188 B.n902 B.n14 585
R189 B.n980 B.n14 585
R190 B.n901 B.n13 585
R191 B.n981 B.n13 585
R192 B.n900 B.n12 585
R193 B.n982 B.n12 585
R194 B.n899 B.n898 585
R195 B.n898 B.n8 585
R196 B.n897 B.n7 585
R197 B.n988 B.n7 585
R198 B.n896 B.n6 585
R199 B.n989 B.n6 585
R200 B.n895 B.n5 585
R201 B.n990 B.n5 585
R202 B.n894 B.n893 585
R203 B.n893 B.n4 585
R204 B.n892 B.n404 585
R205 B.n892 B.n891 585
R206 B.n882 B.n405 585
R207 B.n406 B.n405 585
R208 B.n884 B.n883 585
R209 B.n885 B.n884 585
R210 B.n881 B.n411 585
R211 B.n411 B.n410 585
R212 B.n880 B.n879 585
R213 B.n879 B.n878 585
R214 B.n413 B.n412 585
R215 B.n871 B.n413 585
R216 B.n870 B.n869 585
R217 B.n872 B.n870 585
R218 B.n868 B.n418 585
R219 B.n418 B.n417 585
R220 B.n867 B.n866 585
R221 B.n866 B.n865 585
R222 B.n420 B.n419 585
R223 B.n421 B.n420 585
R224 B.n858 B.n857 585
R225 B.n859 B.n858 585
R226 B.n856 B.n426 585
R227 B.n426 B.n425 585
R228 B.n855 B.n854 585
R229 B.n854 B.n853 585
R230 B.n428 B.n427 585
R231 B.n429 B.n428 585
R232 B.n846 B.n845 585
R233 B.n847 B.n846 585
R234 B.n844 B.n433 585
R235 B.n437 B.n433 585
R236 B.n843 B.n842 585
R237 B.n842 B.n841 585
R238 B.n435 B.n434 585
R239 B.n436 B.n435 585
R240 B.n834 B.n833 585
R241 B.n835 B.n834 585
R242 B.n832 B.n442 585
R243 B.n442 B.n441 585
R244 B.n831 B.n830 585
R245 B.n830 B.n829 585
R246 B.n444 B.n443 585
R247 B.n445 B.n444 585
R248 B.n822 B.n821 585
R249 B.n823 B.n822 585
R250 B.n820 B.n450 585
R251 B.n450 B.n449 585
R252 B.n819 B.n818 585
R253 B.n818 B.n817 585
R254 B.n452 B.n451 585
R255 B.n453 B.n452 585
R256 B.n810 B.n809 585
R257 B.n811 B.n810 585
R258 B.n456 B.n455 585
R259 B.n534 B.n533 585
R260 B.n535 B.n531 585
R261 B.n531 B.n457 585
R262 B.n537 B.n536 585
R263 B.n539 B.n530 585
R264 B.n542 B.n541 585
R265 B.n543 B.n529 585
R266 B.n545 B.n544 585
R267 B.n547 B.n528 585
R268 B.n550 B.n549 585
R269 B.n551 B.n527 585
R270 B.n553 B.n552 585
R271 B.n555 B.n526 585
R272 B.n558 B.n557 585
R273 B.n559 B.n525 585
R274 B.n561 B.n560 585
R275 B.n563 B.n524 585
R276 B.n566 B.n565 585
R277 B.n567 B.n523 585
R278 B.n569 B.n568 585
R279 B.n571 B.n522 585
R280 B.n574 B.n573 585
R281 B.n575 B.n521 585
R282 B.n577 B.n576 585
R283 B.n579 B.n520 585
R284 B.n582 B.n581 585
R285 B.n583 B.n519 585
R286 B.n585 B.n584 585
R287 B.n587 B.n518 585
R288 B.n590 B.n589 585
R289 B.n591 B.n517 585
R290 B.n593 B.n592 585
R291 B.n595 B.n516 585
R292 B.n598 B.n597 585
R293 B.n599 B.n515 585
R294 B.n601 B.n600 585
R295 B.n603 B.n514 585
R296 B.n606 B.n605 585
R297 B.n607 B.n513 585
R298 B.n609 B.n608 585
R299 B.n611 B.n512 585
R300 B.n614 B.n613 585
R301 B.n615 B.n511 585
R302 B.n617 B.n616 585
R303 B.n619 B.n510 585
R304 B.n622 B.n621 585
R305 B.n623 B.n509 585
R306 B.n625 B.n624 585
R307 B.n627 B.n508 585
R308 B.n630 B.n629 585
R309 B.n631 B.n507 585
R310 B.n633 B.n632 585
R311 B.n635 B.n506 585
R312 B.n638 B.n637 585
R313 B.n639 B.n505 585
R314 B.n641 B.n640 585
R315 B.n643 B.n504 585
R316 B.n646 B.n645 585
R317 B.n647 B.n503 585
R318 B.n649 B.n648 585
R319 B.n651 B.n502 585
R320 B.n654 B.n653 585
R321 B.n655 B.n501 585
R322 B.n657 B.n656 585
R323 B.n659 B.n500 585
R324 B.n662 B.n661 585
R325 B.n663 B.n496 585
R326 B.n665 B.n664 585
R327 B.n667 B.n495 585
R328 B.n670 B.n669 585
R329 B.n671 B.n494 585
R330 B.n673 B.n672 585
R331 B.n675 B.n493 585
R332 B.n678 B.n677 585
R333 B.n680 B.n490 585
R334 B.n682 B.n681 585
R335 B.n684 B.n489 585
R336 B.n687 B.n686 585
R337 B.n688 B.n488 585
R338 B.n690 B.n689 585
R339 B.n692 B.n487 585
R340 B.n695 B.n694 585
R341 B.n696 B.n486 585
R342 B.n698 B.n697 585
R343 B.n700 B.n485 585
R344 B.n703 B.n702 585
R345 B.n704 B.n484 585
R346 B.n706 B.n705 585
R347 B.n708 B.n483 585
R348 B.n711 B.n710 585
R349 B.n712 B.n482 585
R350 B.n714 B.n713 585
R351 B.n716 B.n481 585
R352 B.n719 B.n718 585
R353 B.n720 B.n480 585
R354 B.n722 B.n721 585
R355 B.n724 B.n479 585
R356 B.n727 B.n726 585
R357 B.n728 B.n478 585
R358 B.n730 B.n729 585
R359 B.n732 B.n477 585
R360 B.n735 B.n734 585
R361 B.n736 B.n476 585
R362 B.n738 B.n737 585
R363 B.n740 B.n475 585
R364 B.n743 B.n742 585
R365 B.n744 B.n474 585
R366 B.n746 B.n745 585
R367 B.n748 B.n473 585
R368 B.n751 B.n750 585
R369 B.n752 B.n472 585
R370 B.n754 B.n753 585
R371 B.n756 B.n471 585
R372 B.n759 B.n758 585
R373 B.n760 B.n470 585
R374 B.n762 B.n761 585
R375 B.n764 B.n469 585
R376 B.n767 B.n766 585
R377 B.n768 B.n468 585
R378 B.n770 B.n769 585
R379 B.n772 B.n467 585
R380 B.n775 B.n774 585
R381 B.n776 B.n466 585
R382 B.n778 B.n777 585
R383 B.n780 B.n465 585
R384 B.n783 B.n782 585
R385 B.n784 B.n464 585
R386 B.n786 B.n785 585
R387 B.n788 B.n463 585
R388 B.n791 B.n790 585
R389 B.n792 B.n462 585
R390 B.n794 B.n793 585
R391 B.n796 B.n461 585
R392 B.n799 B.n798 585
R393 B.n800 B.n460 585
R394 B.n802 B.n801 585
R395 B.n804 B.n459 585
R396 B.n807 B.n806 585
R397 B.n808 B.n458 585
R398 B.n813 B.n812 585
R399 B.n812 B.n811 585
R400 B.n814 B.n454 585
R401 B.n454 B.n453 585
R402 B.n816 B.n815 585
R403 B.n817 B.n816 585
R404 B.n448 B.n447 585
R405 B.n449 B.n448 585
R406 B.n825 B.n824 585
R407 B.n824 B.n823 585
R408 B.n826 B.n446 585
R409 B.n446 B.n445 585
R410 B.n828 B.n827 585
R411 B.n829 B.n828 585
R412 B.n440 B.n439 585
R413 B.n441 B.n440 585
R414 B.n837 B.n836 585
R415 B.n836 B.n835 585
R416 B.n838 B.n438 585
R417 B.n438 B.n436 585
R418 B.n840 B.n839 585
R419 B.n841 B.n840 585
R420 B.n432 B.n431 585
R421 B.n437 B.n432 585
R422 B.n849 B.n848 585
R423 B.n848 B.n847 585
R424 B.n850 B.n430 585
R425 B.n430 B.n429 585
R426 B.n852 B.n851 585
R427 B.n853 B.n852 585
R428 B.n424 B.n423 585
R429 B.n425 B.n424 585
R430 B.n861 B.n860 585
R431 B.n860 B.n859 585
R432 B.n862 B.n422 585
R433 B.n422 B.n421 585
R434 B.n864 B.n863 585
R435 B.n865 B.n864 585
R436 B.n416 B.n415 585
R437 B.n417 B.n416 585
R438 B.n874 B.n873 585
R439 B.n873 B.n872 585
R440 B.n875 B.n414 585
R441 B.n871 B.n414 585
R442 B.n877 B.n876 585
R443 B.n878 B.n877 585
R444 B.n409 B.n408 585
R445 B.n410 B.n409 585
R446 B.n887 B.n886 585
R447 B.n886 B.n885 585
R448 B.n888 B.n407 585
R449 B.n407 B.n406 585
R450 B.n890 B.n889 585
R451 B.n891 B.n890 585
R452 B.n2 B.n0 585
R453 B.n4 B.n2 585
R454 B.n3 B.n1 585
R455 B.n989 B.n3 585
R456 B.n987 B.n986 585
R457 B.n988 B.n987 585
R458 B.n985 B.n9 585
R459 B.n9 B.n8 585
R460 B.n984 B.n983 585
R461 B.n983 B.n982 585
R462 B.n11 B.n10 585
R463 B.n981 B.n11 585
R464 B.n979 B.n978 585
R465 B.n980 B.n979 585
R466 B.n977 B.n15 585
R467 B.n18 B.n15 585
R468 B.n976 B.n975 585
R469 B.n975 B.n974 585
R470 B.n17 B.n16 585
R471 B.n973 B.n17 585
R472 B.n971 B.n970 585
R473 B.n972 B.n971 585
R474 B.n969 B.n23 585
R475 B.n23 B.n22 585
R476 B.n968 B.n967 585
R477 B.n967 B.n966 585
R478 B.n25 B.n24 585
R479 B.n965 B.n25 585
R480 B.n963 B.n962 585
R481 B.n964 B.n963 585
R482 B.n961 B.n30 585
R483 B.n30 B.n29 585
R484 B.n960 B.n959 585
R485 B.n959 B.n958 585
R486 B.n32 B.n31 585
R487 B.n957 B.n32 585
R488 B.n955 B.n954 585
R489 B.n956 B.n955 585
R490 B.n953 B.n37 585
R491 B.n37 B.n36 585
R492 B.n952 B.n951 585
R493 B.n951 B.n950 585
R494 B.n39 B.n38 585
R495 B.n949 B.n39 585
R496 B.n947 B.n946 585
R497 B.n948 B.n947 585
R498 B.n945 B.n44 585
R499 B.n44 B.n43 585
R500 B.n944 B.n943 585
R501 B.n943 B.n942 585
R502 B.n46 B.n45 585
R503 B.n941 B.n46 585
R504 B.n939 B.n938 585
R505 B.n940 B.n939 585
R506 B.n937 B.n51 585
R507 B.n51 B.n50 585
R508 B.n936 B.n935 585
R509 B.n935 B.n934 585
R510 B.n992 B.n991 585
R511 B.n991 B.n990 585
R512 B.n812 B.n456 559.769
R513 B.n935 B.n53 559.769
R514 B.n810 B.n458 559.769
R515 B.n932 B.n54 559.769
R516 B.n933 B.n123 256.663
R517 B.n933 B.n122 256.663
R518 B.n933 B.n121 256.663
R519 B.n933 B.n120 256.663
R520 B.n933 B.n119 256.663
R521 B.n933 B.n118 256.663
R522 B.n933 B.n117 256.663
R523 B.n933 B.n116 256.663
R524 B.n933 B.n115 256.663
R525 B.n933 B.n114 256.663
R526 B.n933 B.n113 256.663
R527 B.n933 B.n112 256.663
R528 B.n933 B.n111 256.663
R529 B.n933 B.n110 256.663
R530 B.n933 B.n109 256.663
R531 B.n933 B.n108 256.663
R532 B.n933 B.n107 256.663
R533 B.n933 B.n106 256.663
R534 B.n933 B.n105 256.663
R535 B.n933 B.n104 256.663
R536 B.n933 B.n103 256.663
R537 B.n933 B.n102 256.663
R538 B.n933 B.n101 256.663
R539 B.n933 B.n100 256.663
R540 B.n933 B.n99 256.663
R541 B.n933 B.n98 256.663
R542 B.n933 B.n97 256.663
R543 B.n933 B.n96 256.663
R544 B.n933 B.n95 256.663
R545 B.n933 B.n94 256.663
R546 B.n933 B.n93 256.663
R547 B.n933 B.n92 256.663
R548 B.n933 B.n91 256.663
R549 B.n933 B.n90 256.663
R550 B.n933 B.n89 256.663
R551 B.n933 B.n88 256.663
R552 B.n933 B.n87 256.663
R553 B.n933 B.n86 256.663
R554 B.n933 B.n85 256.663
R555 B.n933 B.n84 256.663
R556 B.n933 B.n83 256.663
R557 B.n933 B.n82 256.663
R558 B.n933 B.n81 256.663
R559 B.n933 B.n80 256.663
R560 B.n933 B.n79 256.663
R561 B.n933 B.n78 256.663
R562 B.n933 B.n77 256.663
R563 B.n933 B.n76 256.663
R564 B.n933 B.n75 256.663
R565 B.n933 B.n74 256.663
R566 B.n933 B.n73 256.663
R567 B.n933 B.n72 256.663
R568 B.n933 B.n71 256.663
R569 B.n933 B.n70 256.663
R570 B.n933 B.n69 256.663
R571 B.n933 B.n68 256.663
R572 B.n933 B.n67 256.663
R573 B.n933 B.n66 256.663
R574 B.n933 B.n65 256.663
R575 B.n933 B.n64 256.663
R576 B.n933 B.n63 256.663
R577 B.n933 B.n62 256.663
R578 B.n933 B.n61 256.663
R579 B.n933 B.n60 256.663
R580 B.n933 B.n59 256.663
R581 B.n933 B.n58 256.663
R582 B.n933 B.n57 256.663
R583 B.n933 B.n56 256.663
R584 B.n933 B.n55 256.663
R585 B.n532 B.n457 256.663
R586 B.n538 B.n457 256.663
R587 B.n540 B.n457 256.663
R588 B.n546 B.n457 256.663
R589 B.n548 B.n457 256.663
R590 B.n554 B.n457 256.663
R591 B.n556 B.n457 256.663
R592 B.n562 B.n457 256.663
R593 B.n564 B.n457 256.663
R594 B.n570 B.n457 256.663
R595 B.n572 B.n457 256.663
R596 B.n578 B.n457 256.663
R597 B.n580 B.n457 256.663
R598 B.n586 B.n457 256.663
R599 B.n588 B.n457 256.663
R600 B.n594 B.n457 256.663
R601 B.n596 B.n457 256.663
R602 B.n602 B.n457 256.663
R603 B.n604 B.n457 256.663
R604 B.n610 B.n457 256.663
R605 B.n612 B.n457 256.663
R606 B.n618 B.n457 256.663
R607 B.n620 B.n457 256.663
R608 B.n626 B.n457 256.663
R609 B.n628 B.n457 256.663
R610 B.n634 B.n457 256.663
R611 B.n636 B.n457 256.663
R612 B.n642 B.n457 256.663
R613 B.n644 B.n457 256.663
R614 B.n650 B.n457 256.663
R615 B.n652 B.n457 256.663
R616 B.n658 B.n457 256.663
R617 B.n660 B.n457 256.663
R618 B.n666 B.n457 256.663
R619 B.n668 B.n457 256.663
R620 B.n674 B.n457 256.663
R621 B.n676 B.n457 256.663
R622 B.n683 B.n457 256.663
R623 B.n685 B.n457 256.663
R624 B.n691 B.n457 256.663
R625 B.n693 B.n457 256.663
R626 B.n699 B.n457 256.663
R627 B.n701 B.n457 256.663
R628 B.n707 B.n457 256.663
R629 B.n709 B.n457 256.663
R630 B.n715 B.n457 256.663
R631 B.n717 B.n457 256.663
R632 B.n723 B.n457 256.663
R633 B.n725 B.n457 256.663
R634 B.n731 B.n457 256.663
R635 B.n733 B.n457 256.663
R636 B.n739 B.n457 256.663
R637 B.n741 B.n457 256.663
R638 B.n747 B.n457 256.663
R639 B.n749 B.n457 256.663
R640 B.n755 B.n457 256.663
R641 B.n757 B.n457 256.663
R642 B.n763 B.n457 256.663
R643 B.n765 B.n457 256.663
R644 B.n771 B.n457 256.663
R645 B.n773 B.n457 256.663
R646 B.n779 B.n457 256.663
R647 B.n781 B.n457 256.663
R648 B.n787 B.n457 256.663
R649 B.n789 B.n457 256.663
R650 B.n795 B.n457 256.663
R651 B.n797 B.n457 256.663
R652 B.n803 B.n457 256.663
R653 B.n805 B.n457 256.663
R654 B.n812 B.n454 163.367
R655 B.n816 B.n454 163.367
R656 B.n816 B.n448 163.367
R657 B.n824 B.n448 163.367
R658 B.n824 B.n446 163.367
R659 B.n828 B.n446 163.367
R660 B.n828 B.n440 163.367
R661 B.n836 B.n440 163.367
R662 B.n836 B.n438 163.367
R663 B.n840 B.n438 163.367
R664 B.n840 B.n432 163.367
R665 B.n848 B.n432 163.367
R666 B.n848 B.n430 163.367
R667 B.n852 B.n430 163.367
R668 B.n852 B.n424 163.367
R669 B.n860 B.n424 163.367
R670 B.n860 B.n422 163.367
R671 B.n864 B.n422 163.367
R672 B.n864 B.n416 163.367
R673 B.n873 B.n416 163.367
R674 B.n873 B.n414 163.367
R675 B.n877 B.n414 163.367
R676 B.n877 B.n409 163.367
R677 B.n886 B.n409 163.367
R678 B.n886 B.n407 163.367
R679 B.n890 B.n407 163.367
R680 B.n890 B.n2 163.367
R681 B.n991 B.n2 163.367
R682 B.n991 B.n3 163.367
R683 B.n987 B.n3 163.367
R684 B.n987 B.n9 163.367
R685 B.n983 B.n9 163.367
R686 B.n983 B.n11 163.367
R687 B.n979 B.n11 163.367
R688 B.n979 B.n15 163.367
R689 B.n975 B.n15 163.367
R690 B.n975 B.n17 163.367
R691 B.n971 B.n17 163.367
R692 B.n971 B.n23 163.367
R693 B.n967 B.n23 163.367
R694 B.n967 B.n25 163.367
R695 B.n963 B.n25 163.367
R696 B.n963 B.n30 163.367
R697 B.n959 B.n30 163.367
R698 B.n959 B.n32 163.367
R699 B.n955 B.n32 163.367
R700 B.n955 B.n37 163.367
R701 B.n951 B.n37 163.367
R702 B.n951 B.n39 163.367
R703 B.n947 B.n39 163.367
R704 B.n947 B.n44 163.367
R705 B.n943 B.n44 163.367
R706 B.n943 B.n46 163.367
R707 B.n939 B.n46 163.367
R708 B.n939 B.n51 163.367
R709 B.n935 B.n51 163.367
R710 B.n533 B.n531 163.367
R711 B.n537 B.n531 163.367
R712 B.n541 B.n539 163.367
R713 B.n545 B.n529 163.367
R714 B.n549 B.n547 163.367
R715 B.n553 B.n527 163.367
R716 B.n557 B.n555 163.367
R717 B.n561 B.n525 163.367
R718 B.n565 B.n563 163.367
R719 B.n569 B.n523 163.367
R720 B.n573 B.n571 163.367
R721 B.n577 B.n521 163.367
R722 B.n581 B.n579 163.367
R723 B.n585 B.n519 163.367
R724 B.n589 B.n587 163.367
R725 B.n593 B.n517 163.367
R726 B.n597 B.n595 163.367
R727 B.n601 B.n515 163.367
R728 B.n605 B.n603 163.367
R729 B.n609 B.n513 163.367
R730 B.n613 B.n611 163.367
R731 B.n617 B.n511 163.367
R732 B.n621 B.n619 163.367
R733 B.n625 B.n509 163.367
R734 B.n629 B.n627 163.367
R735 B.n633 B.n507 163.367
R736 B.n637 B.n635 163.367
R737 B.n641 B.n505 163.367
R738 B.n645 B.n643 163.367
R739 B.n649 B.n503 163.367
R740 B.n653 B.n651 163.367
R741 B.n657 B.n501 163.367
R742 B.n661 B.n659 163.367
R743 B.n665 B.n496 163.367
R744 B.n669 B.n667 163.367
R745 B.n673 B.n494 163.367
R746 B.n677 B.n675 163.367
R747 B.n682 B.n490 163.367
R748 B.n686 B.n684 163.367
R749 B.n690 B.n488 163.367
R750 B.n694 B.n692 163.367
R751 B.n698 B.n486 163.367
R752 B.n702 B.n700 163.367
R753 B.n706 B.n484 163.367
R754 B.n710 B.n708 163.367
R755 B.n714 B.n482 163.367
R756 B.n718 B.n716 163.367
R757 B.n722 B.n480 163.367
R758 B.n726 B.n724 163.367
R759 B.n730 B.n478 163.367
R760 B.n734 B.n732 163.367
R761 B.n738 B.n476 163.367
R762 B.n742 B.n740 163.367
R763 B.n746 B.n474 163.367
R764 B.n750 B.n748 163.367
R765 B.n754 B.n472 163.367
R766 B.n758 B.n756 163.367
R767 B.n762 B.n470 163.367
R768 B.n766 B.n764 163.367
R769 B.n770 B.n468 163.367
R770 B.n774 B.n772 163.367
R771 B.n778 B.n466 163.367
R772 B.n782 B.n780 163.367
R773 B.n786 B.n464 163.367
R774 B.n790 B.n788 163.367
R775 B.n794 B.n462 163.367
R776 B.n798 B.n796 163.367
R777 B.n802 B.n460 163.367
R778 B.n806 B.n804 163.367
R779 B.n810 B.n452 163.367
R780 B.n818 B.n452 163.367
R781 B.n818 B.n450 163.367
R782 B.n822 B.n450 163.367
R783 B.n822 B.n444 163.367
R784 B.n830 B.n444 163.367
R785 B.n830 B.n442 163.367
R786 B.n834 B.n442 163.367
R787 B.n834 B.n435 163.367
R788 B.n842 B.n435 163.367
R789 B.n842 B.n433 163.367
R790 B.n846 B.n433 163.367
R791 B.n846 B.n428 163.367
R792 B.n854 B.n428 163.367
R793 B.n854 B.n426 163.367
R794 B.n858 B.n426 163.367
R795 B.n858 B.n420 163.367
R796 B.n866 B.n420 163.367
R797 B.n866 B.n418 163.367
R798 B.n870 B.n418 163.367
R799 B.n870 B.n413 163.367
R800 B.n879 B.n413 163.367
R801 B.n879 B.n411 163.367
R802 B.n884 B.n411 163.367
R803 B.n884 B.n405 163.367
R804 B.n892 B.n405 163.367
R805 B.n893 B.n892 163.367
R806 B.n893 B.n5 163.367
R807 B.n6 B.n5 163.367
R808 B.n7 B.n6 163.367
R809 B.n898 B.n7 163.367
R810 B.n898 B.n12 163.367
R811 B.n13 B.n12 163.367
R812 B.n14 B.n13 163.367
R813 B.n903 B.n14 163.367
R814 B.n903 B.n19 163.367
R815 B.n20 B.n19 163.367
R816 B.n21 B.n20 163.367
R817 B.n908 B.n21 163.367
R818 B.n908 B.n26 163.367
R819 B.n27 B.n26 163.367
R820 B.n28 B.n27 163.367
R821 B.n913 B.n28 163.367
R822 B.n913 B.n33 163.367
R823 B.n34 B.n33 163.367
R824 B.n35 B.n34 163.367
R825 B.n918 B.n35 163.367
R826 B.n918 B.n40 163.367
R827 B.n41 B.n40 163.367
R828 B.n42 B.n41 163.367
R829 B.n923 B.n42 163.367
R830 B.n923 B.n47 163.367
R831 B.n48 B.n47 163.367
R832 B.n49 B.n48 163.367
R833 B.n928 B.n49 163.367
R834 B.n928 B.n54 163.367
R835 B.n132 B.n131 163.367
R836 B.n136 B.n135 163.367
R837 B.n140 B.n139 163.367
R838 B.n144 B.n143 163.367
R839 B.n148 B.n147 163.367
R840 B.n152 B.n151 163.367
R841 B.n156 B.n155 163.367
R842 B.n160 B.n159 163.367
R843 B.n164 B.n163 163.367
R844 B.n168 B.n167 163.367
R845 B.n172 B.n171 163.367
R846 B.n176 B.n175 163.367
R847 B.n180 B.n179 163.367
R848 B.n184 B.n183 163.367
R849 B.n188 B.n187 163.367
R850 B.n192 B.n191 163.367
R851 B.n196 B.n195 163.367
R852 B.n200 B.n199 163.367
R853 B.n204 B.n203 163.367
R854 B.n208 B.n207 163.367
R855 B.n212 B.n211 163.367
R856 B.n216 B.n215 163.367
R857 B.n220 B.n219 163.367
R858 B.n224 B.n223 163.367
R859 B.n228 B.n227 163.367
R860 B.n232 B.n231 163.367
R861 B.n236 B.n235 163.367
R862 B.n240 B.n239 163.367
R863 B.n244 B.n243 163.367
R864 B.n248 B.n247 163.367
R865 B.n252 B.n251 163.367
R866 B.n256 B.n255 163.367
R867 B.n261 B.n260 163.367
R868 B.n265 B.n264 163.367
R869 B.n269 B.n268 163.367
R870 B.n273 B.n272 163.367
R871 B.n277 B.n276 163.367
R872 B.n281 B.n280 163.367
R873 B.n285 B.n284 163.367
R874 B.n289 B.n288 163.367
R875 B.n293 B.n292 163.367
R876 B.n297 B.n296 163.367
R877 B.n301 B.n300 163.367
R878 B.n305 B.n304 163.367
R879 B.n309 B.n308 163.367
R880 B.n313 B.n312 163.367
R881 B.n317 B.n316 163.367
R882 B.n321 B.n320 163.367
R883 B.n325 B.n324 163.367
R884 B.n329 B.n328 163.367
R885 B.n333 B.n332 163.367
R886 B.n337 B.n336 163.367
R887 B.n341 B.n340 163.367
R888 B.n345 B.n344 163.367
R889 B.n349 B.n348 163.367
R890 B.n353 B.n352 163.367
R891 B.n357 B.n356 163.367
R892 B.n361 B.n360 163.367
R893 B.n365 B.n364 163.367
R894 B.n369 B.n368 163.367
R895 B.n373 B.n372 163.367
R896 B.n377 B.n376 163.367
R897 B.n381 B.n380 163.367
R898 B.n385 B.n384 163.367
R899 B.n389 B.n388 163.367
R900 B.n393 B.n392 163.367
R901 B.n397 B.n396 163.367
R902 B.n401 B.n400 163.367
R903 B.n932 B.n124 163.367
R904 B.n491 B.t13 92.7464
R905 B.n125 B.t22 92.7464
R906 B.n497 B.t20 92.7196
R907 B.n128 B.t16 92.7196
R908 B.n532 B.n456 71.676
R909 B.n538 B.n537 71.676
R910 B.n541 B.n540 71.676
R911 B.n546 B.n545 71.676
R912 B.n549 B.n548 71.676
R913 B.n554 B.n553 71.676
R914 B.n557 B.n556 71.676
R915 B.n562 B.n561 71.676
R916 B.n565 B.n564 71.676
R917 B.n570 B.n569 71.676
R918 B.n573 B.n572 71.676
R919 B.n578 B.n577 71.676
R920 B.n581 B.n580 71.676
R921 B.n586 B.n585 71.676
R922 B.n589 B.n588 71.676
R923 B.n594 B.n593 71.676
R924 B.n597 B.n596 71.676
R925 B.n602 B.n601 71.676
R926 B.n605 B.n604 71.676
R927 B.n610 B.n609 71.676
R928 B.n613 B.n612 71.676
R929 B.n618 B.n617 71.676
R930 B.n621 B.n620 71.676
R931 B.n626 B.n625 71.676
R932 B.n629 B.n628 71.676
R933 B.n634 B.n633 71.676
R934 B.n637 B.n636 71.676
R935 B.n642 B.n641 71.676
R936 B.n645 B.n644 71.676
R937 B.n650 B.n649 71.676
R938 B.n653 B.n652 71.676
R939 B.n658 B.n657 71.676
R940 B.n661 B.n660 71.676
R941 B.n666 B.n665 71.676
R942 B.n669 B.n668 71.676
R943 B.n674 B.n673 71.676
R944 B.n677 B.n676 71.676
R945 B.n683 B.n682 71.676
R946 B.n686 B.n685 71.676
R947 B.n691 B.n690 71.676
R948 B.n694 B.n693 71.676
R949 B.n699 B.n698 71.676
R950 B.n702 B.n701 71.676
R951 B.n707 B.n706 71.676
R952 B.n710 B.n709 71.676
R953 B.n715 B.n714 71.676
R954 B.n718 B.n717 71.676
R955 B.n723 B.n722 71.676
R956 B.n726 B.n725 71.676
R957 B.n731 B.n730 71.676
R958 B.n734 B.n733 71.676
R959 B.n739 B.n738 71.676
R960 B.n742 B.n741 71.676
R961 B.n747 B.n746 71.676
R962 B.n750 B.n749 71.676
R963 B.n755 B.n754 71.676
R964 B.n758 B.n757 71.676
R965 B.n763 B.n762 71.676
R966 B.n766 B.n765 71.676
R967 B.n771 B.n770 71.676
R968 B.n774 B.n773 71.676
R969 B.n779 B.n778 71.676
R970 B.n782 B.n781 71.676
R971 B.n787 B.n786 71.676
R972 B.n790 B.n789 71.676
R973 B.n795 B.n794 71.676
R974 B.n798 B.n797 71.676
R975 B.n803 B.n802 71.676
R976 B.n806 B.n805 71.676
R977 B.n55 B.n53 71.676
R978 B.n132 B.n56 71.676
R979 B.n136 B.n57 71.676
R980 B.n140 B.n58 71.676
R981 B.n144 B.n59 71.676
R982 B.n148 B.n60 71.676
R983 B.n152 B.n61 71.676
R984 B.n156 B.n62 71.676
R985 B.n160 B.n63 71.676
R986 B.n164 B.n64 71.676
R987 B.n168 B.n65 71.676
R988 B.n172 B.n66 71.676
R989 B.n176 B.n67 71.676
R990 B.n180 B.n68 71.676
R991 B.n184 B.n69 71.676
R992 B.n188 B.n70 71.676
R993 B.n192 B.n71 71.676
R994 B.n196 B.n72 71.676
R995 B.n200 B.n73 71.676
R996 B.n204 B.n74 71.676
R997 B.n208 B.n75 71.676
R998 B.n212 B.n76 71.676
R999 B.n216 B.n77 71.676
R1000 B.n220 B.n78 71.676
R1001 B.n224 B.n79 71.676
R1002 B.n228 B.n80 71.676
R1003 B.n232 B.n81 71.676
R1004 B.n236 B.n82 71.676
R1005 B.n240 B.n83 71.676
R1006 B.n244 B.n84 71.676
R1007 B.n248 B.n85 71.676
R1008 B.n252 B.n86 71.676
R1009 B.n256 B.n87 71.676
R1010 B.n261 B.n88 71.676
R1011 B.n265 B.n89 71.676
R1012 B.n269 B.n90 71.676
R1013 B.n273 B.n91 71.676
R1014 B.n277 B.n92 71.676
R1015 B.n281 B.n93 71.676
R1016 B.n285 B.n94 71.676
R1017 B.n289 B.n95 71.676
R1018 B.n293 B.n96 71.676
R1019 B.n297 B.n97 71.676
R1020 B.n301 B.n98 71.676
R1021 B.n305 B.n99 71.676
R1022 B.n309 B.n100 71.676
R1023 B.n313 B.n101 71.676
R1024 B.n317 B.n102 71.676
R1025 B.n321 B.n103 71.676
R1026 B.n325 B.n104 71.676
R1027 B.n329 B.n105 71.676
R1028 B.n333 B.n106 71.676
R1029 B.n337 B.n107 71.676
R1030 B.n341 B.n108 71.676
R1031 B.n345 B.n109 71.676
R1032 B.n349 B.n110 71.676
R1033 B.n353 B.n111 71.676
R1034 B.n357 B.n112 71.676
R1035 B.n361 B.n113 71.676
R1036 B.n365 B.n114 71.676
R1037 B.n369 B.n115 71.676
R1038 B.n373 B.n116 71.676
R1039 B.n377 B.n117 71.676
R1040 B.n381 B.n118 71.676
R1041 B.n385 B.n119 71.676
R1042 B.n389 B.n120 71.676
R1043 B.n393 B.n121 71.676
R1044 B.n397 B.n122 71.676
R1045 B.n401 B.n123 71.676
R1046 B.n124 B.n123 71.676
R1047 B.n400 B.n122 71.676
R1048 B.n396 B.n121 71.676
R1049 B.n392 B.n120 71.676
R1050 B.n388 B.n119 71.676
R1051 B.n384 B.n118 71.676
R1052 B.n380 B.n117 71.676
R1053 B.n376 B.n116 71.676
R1054 B.n372 B.n115 71.676
R1055 B.n368 B.n114 71.676
R1056 B.n364 B.n113 71.676
R1057 B.n360 B.n112 71.676
R1058 B.n356 B.n111 71.676
R1059 B.n352 B.n110 71.676
R1060 B.n348 B.n109 71.676
R1061 B.n344 B.n108 71.676
R1062 B.n340 B.n107 71.676
R1063 B.n336 B.n106 71.676
R1064 B.n332 B.n105 71.676
R1065 B.n328 B.n104 71.676
R1066 B.n324 B.n103 71.676
R1067 B.n320 B.n102 71.676
R1068 B.n316 B.n101 71.676
R1069 B.n312 B.n100 71.676
R1070 B.n308 B.n99 71.676
R1071 B.n304 B.n98 71.676
R1072 B.n300 B.n97 71.676
R1073 B.n296 B.n96 71.676
R1074 B.n292 B.n95 71.676
R1075 B.n288 B.n94 71.676
R1076 B.n284 B.n93 71.676
R1077 B.n280 B.n92 71.676
R1078 B.n276 B.n91 71.676
R1079 B.n272 B.n90 71.676
R1080 B.n268 B.n89 71.676
R1081 B.n264 B.n88 71.676
R1082 B.n260 B.n87 71.676
R1083 B.n255 B.n86 71.676
R1084 B.n251 B.n85 71.676
R1085 B.n247 B.n84 71.676
R1086 B.n243 B.n83 71.676
R1087 B.n239 B.n82 71.676
R1088 B.n235 B.n81 71.676
R1089 B.n231 B.n80 71.676
R1090 B.n227 B.n79 71.676
R1091 B.n223 B.n78 71.676
R1092 B.n219 B.n77 71.676
R1093 B.n215 B.n76 71.676
R1094 B.n211 B.n75 71.676
R1095 B.n207 B.n74 71.676
R1096 B.n203 B.n73 71.676
R1097 B.n199 B.n72 71.676
R1098 B.n195 B.n71 71.676
R1099 B.n191 B.n70 71.676
R1100 B.n187 B.n69 71.676
R1101 B.n183 B.n68 71.676
R1102 B.n179 B.n67 71.676
R1103 B.n175 B.n66 71.676
R1104 B.n171 B.n65 71.676
R1105 B.n167 B.n64 71.676
R1106 B.n163 B.n63 71.676
R1107 B.n159 B.n62 71.676
R1108 B.n155 B.n61 71.676
R1109 B.n151 B.n60 71.676
R1110 B.n147 B.n59 71.676
R1111 B.n143 B.n58 71.676
R1112 B.n139 B.n57 71.676
R1113 B.n135 B.n56 71.676
R1114 B.n131 B.n55 71.676
R1115 B.n533 B.n532 71.676
R1116 B.n539 B.n538 71.676
R1117 B.n540 B.n529 71.676
R1118 B.n547 B.n546 71.676
R1119 B.n548 B.n527 71.676
R1120 B.n555 B.n554 71.676
R1121 B.n556 B.n525 71.676
R1122 B.n563 B.n562 71.676
R1123 B.n564 B.n523 71.676
R1124 B.n571 B.n570 71.676
R1125 B.n572 B.n521 71.676
R1126 B.n579 B.n578 71.676
R1127 B.n580 B.n519 71.676
R1128 B.n587 B.n586 71.676
R1129 B.n588 B.n517 71.676
R1130 B.n595 B.n594 71.676
R1131 B.n596 B.n515 71.676
R1132 B.n603 B.n602 71.676
R1133 B.n604 B.n513 71.676
R1134 B.n611 B.n610 71.676
R1135 B.n612 B.n511 71.676
R1136 B.n619 B.n618 71.676
R1137 B.n620 B.n509 71.676
R1138 B.n627 B.n626 71.676
R1139 B.n628 B.n507 71.676
R1140 B.n635 B.n634 71.676
R1141 B.n636 B.n505 71.676
R1142 B.n643 B.n642 71.676
R1143 B.n644 B.n503 71.676
R1144 B.n651 B.n650 71.676
R1145 B.n652 B.n501 71.676
R1146 B.n659 B.n658 71.676
R1147 B.n660 B.n496 71.676
R1148 B.n667 B.n666 71.676
R1149 B.n668 B.n494 71.676
R1150 B.n675 B.n674 71.676
R1151 B.n676 B.n490 71.676
R1152 B.n684 B.n683 71.676
R1153 B.n685 B.n488 71.676
R1154 B.n692 B.n691 71.676
R1155 B.n693 B.n486 71.676
R1156 B.n700 B.n699 71.676
R1157 B.n701 B.n484 71.676
R1158 B.n708 B.n707 71.676
R1159 B.n709 B.n482 71.676
R1160 B.n716 B.n715 71.676
R1161 B.n717 B.n480 71.676
R1162 B.n724 B.n723 71.676
R1163 B.n725 B.n478 71.676
R1164 B.n732 B.n731 71.676
R1165 B.n733 B.n476 71.676
R1166 B.n740 B.n739 71.676
R1167 B.n741 B.n474 71.676
R1168 B.n748 B.n747 71.676
R1169 B.n749 B.n472 71.676
R1170 B.n756 B.n755 71.676
R1171 B.n757 B.n470 71.676
R1172 B.n764 B.n763 71.676
R1173 B.n765 B.n468 71.676
R1174 B.n772 B.n771 71.676
R1175 B.n773 B.n466 71.676
R1176 B.n780 B.n779 71.676
R1177 B.n781 B.n464 71.676
R1178 B.n788 B.n787 71.676
R1179 B.n789 B.n462 71.676
R1180 B.n796 B.n795 71.676
R1181 B.n797 B.n460 71.676
R1182 B.n804 B.n803 71.676
R1183 B.n805 B.n458 71.676
R1184 B.n492 B.t12 70.6373
R1185 B.n126 B.t23 70.6373
R1186 B.n498 B.t19 70.6105
R1187 B.n129 B.t17 70.6105
R1188 B.n811 B.n457 60.7354
R1189 B.n934 B.n933 60.7354
R1190 B.n679 B.n492 59.5399
R1191 B.n499 B.n498 59.5399
R1192 B.n258 B.n129 59.5399
R1193 B.n127 B.n126 59.5399
R1194 B.n936 B.n52 36.3712
R1195 B.n931 B.n930 36.3712
R1196 B.n809 B.n808 36.3712
R1197 B.n813 B.n455 36.3712
R1198 B.n811 B.n453 29.7125
R1199 B.n817 B.n453 29.7125
R1200 B.n817 B.n449 29.7125
R1201 B.n823 B.n449 29.7125
R1202 B.n829 B.n445 29.7125
R1203 B.n829 B.n441 29.7125
R1204 B.n835 B.n441 29.7125
R1205 B.n835 B.n436 29.7125
R1206 B.n841 B.n436 29.7125
R1207 B.n841 B.n437 29.7125
R1208 B.n847 B.n429 29.7125
R1209 B.n853 B.n429 29.7125
R1210 B.n859 B.n425 29.7125
R1211 B.n859 B.n421 29.7125
R1212 B.n865 B.n421 29.7125
R1213 B.n872 B.n417 29.7125
R1214 B.n872 B.n871 29.7125
R1215 B.n878 B.n410 29.7125
R1216 B.n885 B.n410 29.7125
R1217 B.n891 B.n406 29.7125
R1218 B.n891 B.n4 29.7125
R1219 B.n990 B.n4 29.7125
R1220 B.n990 B.n989 29.7125
R1221 B.n989 B.n988 29.7125
R1222 B.n988 B.n8 29.7125
R1223 B.n982 B.n981 29.7125
R1224 B.n981 B.n980 29.7125
R1225 B.n974 B.n18 29.7125
R1226 B.n974 B.n973 29.7125
R1227 B.n972 B.n22 29.7125
R1228 B.n966 B.n22 29.7125
R1229 B.n966 B.n965 29.7125
R1230 B.n964 B.n29 29.7125
R1231 B.n958 B.n29 29.7125
R1232 B.n957 B.n956 29.7125
R1233 B.n956 B.n36 29.7125
R1234 B.n950 B.n36 29.7125
R1235 B.n950 B.n949 29.7125
R1236 B.n949 B.n948 29.7125
R1237 B.n948 B.n43 29.7125
R1238 B.n942 B.n941 29.7125
R1239 B.n941 B.n940 29.7125
R1240 B.n940 B.n50 29.7125
R1241 B.n934 B.n50 29.7125
R1242 B.t4 B.n417 29.2756
R1243 B.n973 B.t9 29.2756
R1244 B.n823 B.t11 22.2845
R1245 B.n942 B.t15 22.2845
R1246 B.n492 B.n491 22.1096
R1247 B.n498 B.n497 22.1096
R1248 B.n129 B.n128 22.1096
R1249 B.n126 B.n125 22.1096
R1250 B.n885 B.t5 21.4106
R1251 B.n982 B.t6 21.4106
R1252 B.n847 B.t1 20.5367
R1253 B.n958 B.t8 20.5367
R1254 B.n853 B.t0 19.6629
R1255 B.t3 B.n964 19.6629
R1256 B.n878 B.t2 18.789
R1257 B.n980 B.t7 18.789
R1258 B B.n992 18.0485
R1259 B.n871 B.t2 10.924
R1260 B.n18 B.t7 10.924
R1261 B.n130 B.n52 10.6151
R1262 B.n133 B.n130 10.6151
R1263 B.n134 B.n133 10.6151
R1264 B.n137 B.n134 10.6151
R1265 B.n138 B.n137 10.6151
R1266 B.n141 B.n138 10.6151
R1267 B.n142 B.n141 10.6151
R1268 B.n145 B.n142 10.6151
R1269 B.n146 B.n145 10.6151
R1270 B.n149 B.n146 10.6151
R1271 B.n150 B.n149 10.6151
R1272 B.n153 B.n150 10.6151
R1273 B.n154 B.n153 10.6151
R1274 B.n157 B.n154 10.6151
R1275 B.n158 B.n157 10.6151
R1276 B.n161 B.n158 10.6151
R1277 B.n162 B.n161 10.6151
R1278 B.n165 B.n162 10.6151
R1279 B.n166 B.n165 10.6151
R1280 B.n169 B.n166 10.6151
R1281 B.n170 B.n169 10.6151
R1282 B.n173 B.n170 10.6151
R1283 B.n174 B.n173 10.6151
R1284 B.n177 B.n174 10.6151
R1285 B.n178 B.n177 10.6151
R1286 B.n181 B.n178 10.6151
R1287 B.n182 B.n181 10.6151
R1288 B.n185 B.n182 10.6151
R1289 B.n186 B.n185 10.6151
R1290 B.n189 B.n186 10.6151
R1291 B.n190 B.n189 10.6151
R1292 B.n193 B.n190 10.6151
R1293 B.n194 B.n193 10.6151
R1294 B.n197 B.n194 10.6151
R1295 B.n198 B.n197 10.6151
R1296 B.n201 B.n198 10.6151
R1297 B.n202 B.n201 10.6151
R1298 B.n205 B.n202 10.6151
R1299 B.n206 B.n205 10.6151
R1300 B.n209 B.n206 10.6151
R1301 B.n210 B.n209 10.6151
R1302 B.n213 B.n210 10.6151
R1303 B.n214 B.n213 10.6151
R1304 B.n217 B.n214 10.6151
R1305 B.n218 B.n217 10.6151
R1306 B.n221 B.n218 10.6151
R1307 B.n222 B.n221 10.6151
R1308 B.n225 B.n222 10.6151
R1309 B.n226 B.n225 10.6151
R1310 B.n229 B.n226 10.6151
R1311 B.n230 B.n229 10.6151
R1312 B.n233 B.n230 10.6151
R1313 B.n234 B.n233 10.6151
R1314 B.n237 B.n234 10.6151
R1315 B.n238 B.n237 10.6151
R1316 B.n241 B.n238 10.6151
R1317 B.n242 B.n241 10.6151
R1318 B.n245 B.n242 10.6151
R1319 B.n246 B.n245 10.6151
R1320 B.n249 B.n246 10.6151
R1321 B.n250 B.n249 10.6151
R1322 B.n253 B.n250 10.6151
R1323 B.n254 B.n253 10.6151
R1324 B.n257 B.n254 10.6151
R1325 B.n262 B.n259 10.6151
R1326 B.n263 B.n262 10.6151
R1327 B.n266 B.n263 10.6151
R1328 B.n267 B.n266 10.6151
R1329 B.n270 B.n267 10.6151
R1330 B.n271 B.n270 10.6151
R1331 B.n274 B.n271 10.6151
R1332 B.n275 B.n274 10.6151
R1333 B.n279 B.n278 10.6151
R1334 B.n282 B.n279 10.6151
R1335 B.n283 B.n282 10.6151
R1336 B.n286 B.n283 10.6151
R1337 B.n287 B.n286 10.6151
R1338 B.n290 B.n287 10.6151
R1339 B.n291 B.n290 10.6151
R1340 B.n294 B.n291 10.6151
R1341 B.n295 B.n294 10.6151
R1342 B.n298 B.n295 10.6151
R1343 B.n299 B.n298 10.6151
R1344 B.n302 B.n299 10.6151
R1345 B.n303 B.n302 10.6151
R1346 B.n306 B.n303 10.6151
R1347 B.n307 B.n306 10.6151
R1348 B.n310 B.n307 10.6151
R1349 B.n311 B.n310 10.6151
R1350 B.n314 B.n311 10.6151
R1351 B.n315 B.n314 10.6151
R1352 B.n318 B.n315 10.6151
R1353 B.n319 B.n318 10.6151
R1354 B.n322 B.n319 10.6151
R1355 B.n323 B.n322 10.6151
R1356 B.n326 B.n323 10.6151
R1357 B.n327 B.n326 10.6151
R1358 B.n330 B.n327 10.6151
R1359 B.n331 B.n330 10.6151
R1360 B.n334 B.n331 10.6151
R1361 B.n335 B.n334 10.6151
R1362 B.n338 B.n335 10.6151
R1363 B.n339 B.n338 10.6151
R1364 B.n342 B.n339 10.6151
R1365 B.n343 B.n342 10.6151
R1366 B.n346 B.n343 10.6151
R1367 B.n347 B.n346 10.6151
R1368 B.n350 B.n347 10.6151
R1369 B.n351 B.n350 10.6151
R1370 B.n354 B.n351 10.6151
R1371 B.n355 B.n354 10.6151
R1372 B.n358 B.n355 10.6151
R1373 B.n359 B.n358 10.6151
R1374 B.n362 B.n359 10.6151
R1375 B.n363 B.n362 10.6151
R1376 B.n366 B.n363 10.6151
R1377 B.n367 B.n366 10.6151
R1378 B.n370 B.n367 10.6151
R1379 B.n371 B.n370 10.6151
R1380 B.n374 B.n371 10.6151
R1381 B.n375 B.n374 10.6151
R1382 B.n378 B.n375 10.6151
R1383 B.n379 B.n378 10.6151
R1384 B.n382 B.n379 10.6151
R1385 B.n383 B.n382 10.6151
R1386 B.n386 B.n383 10.6151
R1387 B.n387 B.n386 10.6151
R1388 B.n390 B.n387 10.6151
R1389 B.n391 B.n390 10.6151
R1390 B.n394 B.n391 10.6151
R1391 B.n395 B.n394 10.6151
R1392 B.n398 B.n395 10.6151
R1393 B.n399 B.n398 10.6151
R1394 B.n402 B.n399 10.6151
R1395 B.n403 B.n402 10.6151
R1396 B.n931 B.n403 10.6151
R1397 B.n809 B.n451 10.6151
R1398 B.n819 B.n451 10.6151
R1399 B.n820 B.n819 10.6151
R1400 B.n821 B.n820 10.6151
R1401 B.n821 B.n443 10.6151
R1402 B.n831 B.n443 10.6151
R1403 B.n832 B.n831 10.6151
R1404 B.n833 B.n832 10.6151
R1405 B.n833 B.n434 10.6151
R1406 B.n843 B.n434 10.6151
R1407 B.n844 B.n843 10.6151
R1408 B.n845 B.n844 10.6151
R1409 B.n845 B.n427 10.6151
R1410 B.n855 B.n427 10.6151
R1411 B.n856 B.n855 10.6151
R1412 B.n857 B.n856 10.6151
R1413 B.n857 B.n419 10.6151
R1414 B.n867 B.n419 10.6151
R1415 B.n868 B.n867 10.6151
R1416 B.n869 B.n868 10.6151
R1417 B.n869 B.n412 10.6151
R1418 B.n880 B.n412 10.6151
R1419 B.n881 B.n880 10.6151
R1420 B.n883 B.n881 10.6151
R1421 B.n883 B.n882 10.6151
R1422 B.n882 B.n404 10.6151
R1423 B.n894 B.n404 10.6151
R1424 B.n895 B.n894 10.6151
R1425 B.n896 B.n895 10.6151
R1426 B.n897 B.n896 10.6151
R1427 B.n899 B.n897 10.6151
R1428 B.n900 B.n899 10.6151
R1429 B.n901 B.n900 10.6151
R1430 B.n902 B.n901 10.6151
R1431 B.n904 B.n902 10.6151
R1432 B.n905 B.n904 10.6151
R1433 B.n906 B.n905 10.6151
R1434 B.n907 B.n906 10.6151
R1435 B.n909 B.n907 10.6151
R1436 B.n910 B.n909 10.6151
R1437 B.n911 B.n910 10.6151
R1438 B.n912 B.n911 10.6151
R1439 B.n914 B.n912 10.6151
R1440 B.n915 B.n914 10.6151
R1441 B.n916 B.n915 10.6151
R1442 B.n917 B.n916 10.6151
R1443 B.n919 B.n917 10.6151
R1444 B.n920 B.n919 10.6151
R1445 B.n921 B.n920 10.6151
R1446 B.n922 B.n921 10.6151
R1447 B.n924 B.n922 10.6151
R1448 B.n925 B.n924 10.6151
R1449 B.n926 B.n925 10.6151
R1450 B.n927 B.n926 10.6151
R1451 B.n929 B.n927 10.6151
R1452 B.n930 B.n929 10.6151
R1453 B.n534 B.n455 10.6151
R1454 B.n535 B.n534 10.6151
R1455 B.n536 B.n535 10.6151
R1456 B.n536 B.n530 10.6151
R1457 B.n542 B.n530 10.6151
R1458 B.n543 B.n542 10.6151
R1459 B.n544 B.n543 10.6151
R1460 B.n544 B.n528 10.6151
R1461 B.n550 B.n528 10.6151
R1462 B.n551 B.n550 10.6151
R1463 B.n552 B.n551 10.6151
R1464 B.n552 B.n526 10.6151
R1465 B.n558 B.n526 10.6151
R1466 B.n559 B.n558 10.6151
R1467 B.n560 B.n559 10.6151
R1468 B.n560 B.n524 10.6151
R1469 B.n566 B.n524 10.6151
R1470 B.n567 B.n566 10.6151
R1471 B.n568 B.n567 10.6151
R1472 B.n568 B.n522 10.6151
R1473 B.n574 B.n522 10.6151
R1474 B.n575 B.n574 10.6151
R1475 B.n576 B.n575 10.6151
R1476 B.n576 B.n520 10.6151
R1477 B.n582 B.n520 10.6151
R1478 B.n583 B.n582 10.6151
R1479 B.n584 B.n583 10.6151
R1480 B.n584 B.n518 10.6151
R1481 B.n590 B.n518 10.6151
R1482 B.n591 B.n590 10.6151
R1483 B.n592 B.n591 10.6151
R1484 B.n592 B.n516 10.6151
R1485 B.n598 B.n516 10.6151
R1486 B.n599 B.n598 10.6151
R1487 B.n600 B.n599 10.6151
R1488 B.n600 B.n514 10.6151
R1489 B.n606 B.n514 10.6151
R1490 B.n607 B.n606 10.6151
R1491 B.n608 B.n607 10.6151
R1492 B.n608 B.n512 10.6151
R1493 B.n614 B.n512 10.6151
R1494 B.n615 B.n614 10.6151
R1495 B.n616 B.n615 10.6151
R1496 B.n616 B.n510 10.6151
R1497 B.n622 B.n510 10.6151
R1498 B.n623 B.n622 10.6151
R1499 B.n624 B.n623 10.6151
R1500 B.n624 B.n508 10.6151
R1501 B.n630 B.n508 10.6151
R1502 B.n631 B.n630 10.6151
R1503 B.n632 B.n631 10.6151
R1504 B.n632 B.n506 10.6151
R1505 B.n638 B.n506 10.6151
R1506 B.n639 B.n638 10.6151
R1507 B.n640 B.n639 10.6151
R1508 B.n640 B.n504 10.6151
R1509 B.n646 B.n504 10.6151
R1510 B.n647 B.n646 10.6151
R1511 B.n648 B.n647 10.6151
R1512 B.n648 B.n502 10.6151
R1513 B.n654 B.n502 10.6151
R1514 B.n655 B.n654 10.6151
R1515 B.n656 B.n655 10.6151
R1516 B.n656 B.n500 10.6151
R1517 B.n663 B.n662 10.6151
R1518 B.n664 B.n663 10.6151
R1519 B.n664 B.n495 10.6151
R1520 B.n670 B.n495 10.6151
R1521 B.n671 B.n670 10.6151
R1522 B.n672 B.n671 10.6151
R1523 B.n672 B.n493 10.6151
R1524 B.n678 B.n493 10.6151
R1525 B.n681 B.n680 10.6151
R1526 B.n681 B.n489 10.6151
R1527 B.n687 B.n489 10.6151
R1528 B.n688 B.n687 10.6151
R1529 B.n689 B.n688 10.6151
R1530 B.n689 B.n487 10.6151
R1531 B.n695 B.n487 10.6151
R1532 B.n696 B.n695 10.6151
R1533 B.n697 B.n696 10.6151
R1534 B.n697 B.n485 10.6151
R1535 B.n703 B.n485 10.6151
R1536 B.n704 B.n703 10.6151
R1537 B.n705 B.n704 10.6151
R1538 B.n705 B.n483 10.6151
R1539 B.n711 B.n483 10.6151
R1540 B.n712 B.n711 10.6151
R1541 B.n713 B.n712 10.6151
R1542 B.n713 B.n481 10.6151
R1543 B.n719 B.n481 10.6151
R1544 B.n720 B.n719 10.6151
R1545 B.n721 B.n720 10.6151
R1546 B.n721 B.n479 10.6151
R1547 B.n727 B.n479 10.6151
R1548 B.n728 B.n727 10.6151
R1549 B.n729 B.n728 10.6151
R1550 B.n729 B.n477 10.6151
R1551 B.n735 B.n477 10.6151
R1552 B.n736 B.n735 10.6151
R1553 B.n737 B.n736 10.6151
R1554 B.n737 B.n475 10.6151
R1555 B.n743 B.n475 10.6151
R1556 B.n744 B.n743 10.6151
R1557 B.n745 B.n744 10.6151
R1558 B.n745 B.n473 10.6151
R1559 B.n751 B.n473 10.6151
R1560 B.n752 B.n751 10.6151
R1561 B.n753 B.n752 10.6151
R1562 B.n753 B.n471 10.6151
R1563 B.n759 B.n471 10.6151
R1564 B.n760 B.n759 10.6151
R1565 B.n761 B.n760 10.6151
R1566 B.n761 B.n469 10.6151
R1567 B.n767 B.n469 10.6151
R1568 B.n768 B.n767 10.6151
R1569 B.n769 B.n768 10.6151
R1570 B.n769 B.n467 10.6151
R1571 B.n775 B.n467 10.6151
R1572 B.n776 B.n775 10.6151
R1573 B.n777 B.n776 10.6151
R1574 B.n777 B.n465 10.6151
R1575 B.n783 B.n465 10.6151
R1576 B.n784 B.n783 10.6151
R1577 B.n785 B.n784 10.6151
R1578 B.n785 B.n463 10.6151
R1579 B.n791 B.n463 10.6151
R1580 B.n792 B.n791 10.6151
R1581 B.n793 B.n792 10.6151
R1582 B.n793 B.n461 10.6151
R1583 B.n799 B.n461 10.6151
R1584 B.n800 B.n799 10.6151
R1585 B.n801 B.n800 10.6151
R1586 B.n801 B.n459 10.6151
R1587 B.n807 B.n459 10.6151
R1588 B.n808 B.n807 10.6151
R1589 B.n814 B.n813 10.6151
R1590 B.n815 B.n814 10.6151
R1591 B.n815 B.n447 10.6151
R1592 B.n825 B.n447 10.6151
R1593 B.n826 B.n825 10.6151
R1594 B.n827 B.n826 10.6151
R1595 B.n827 B.n439 10.6151
R1596 B.n837 B.n439 10.6151
R1597 B.n838 B.n837 10.6151
R1598 B.n839 B.n838 10.6151
R1599 B.n839 B.n431 10.6151
R1600 B.n849 B.n431 10.6151
R1601 B.n850 B.n849 10.6151
R1602 B.n851 B.n850 10.6151
R1603 B.n851 B.n423 10.6151
R1604 B.n861 B.n423 10.6151
R1605 B.n862 B.n861 10.6151
R1606 B.n863 B.n862 10.6151
R1607 B.n863 B.n415 10.6151
R1608 B.n874 B.n415 10.6151
R1609 B.n875 B.n874 10.6151
R1610 B.n876 B.n875 10.6151
R1611 B.n876 B.n408 10.6151
R1612 B.n887 B.n408 10.6151
R1613 B.n888 B.n887 10.6151
R1614 B.n889 B.n888 10.6151
R1615 B.n889 B.n0 10.6151
R1616 B.n986 B.n1 10.6151
R1617 B.n986 B.n985 10.6151
R1618 B.n985 B.n984 10.6151
R1619 B.n984 B.n10 10.6151
R1620 B.n978 B.n10 10.6151
R1621 B.n978 B.n977 10.6151
R1622 B.n977 B.n976 10.6151
R1623 B.n976 B.n16 10.6151
R1624 B.n970 B.n16 10.6151
R1625 B.n970 B.n969 10.6151
R1626 B.n969 B.n968 10.6151
R1627 B.n968 B.n24 10.6151
R1628 B.n962 B.n24 10.6151
R1629 B.n962 B.n961 10.6151
R1630 B.n961 B.n960 10.6151
R1631 B.n960 B.n31 10.6151
R1632 B.n954 B.n31 10.6151
R1633 B.n954 B.n953 10.6151
R1634 B.n953 B.n952 10.6151
R1635 B.n952 B.n38 10.6151
R1636 B.n946 B.n38 10.6151
R1637 B.n946 B.n945 10.6151
R1638 B.n945 B.n944 10.6151
R1639 B.n944 B.n45 10.6151
R1640 B.n938 B.n45 10.6151
R1641 B.n938 B.n937 10.6151
R1642 B.n937 B.n936 10.6151
R1643 B.t0 B.n425 10.0502
R1644 B.n965 B.t3 10.0502
R1645 B.n437 B.t1 9.17627
R1646 B.t8 B.n957 9.17627
R1647 B.t5 B.n406 8.30239
R1648 B.t6 B.n8 8.30239
R1649 B.t11 B.n445 7.4285
R1650 B.t15 B.n43 7.4285
R1651 B.n259 B.n258 6.5566
R1652 B.n275 B.n127 6.5566
R1653 B.n662 B.n499 6.5566
R1654 B.n679 B.n678 6.5566
R1655 B.n258 B.n257 4.05904
R1656 B.n278 B.n127 4.05904
R1657 B.n500 B.n499 4.05904
R1658 B.n680 B.n679 4.05904
R1659 B.n992 B.n0 2.81026
R1660 B.n992 B.n1 2.81026
R1661 B.n865 B.t4 0.437441
R1662 B.t9 B.n972 0.437441
R1663 VN.n3 VN.t1 664.332
R1664 VN.n13 VN.t5 664.332
R1665 VN.n2 VN.t8 640.585
R1666 VN.n1 VN.t7 640.585
R1667 VN.n6 VN.t4 640.585
R1668 VN.n8 VN.t3 640.585
R1669 VN.n12 VN.t9 640.585
R1670 VN.n11 VN.t2 640.585
R1671 VN.n16 VN.t6 640.585
R1672 VN.n18 VN.t0 640.585
R1673 VN.n9 VN.n8 161.3
R1674 VN.n19 VN.n18 161.3
R1675 VN.n17 VN.n10 161.3
R1676 VN.n7 VN.n0 161.3
R1677 VN.n16 VN.n15 80.6037
R1678 VN.n14 VN.n11 80.6037
R1679 VN.n6 VN.n5 80.6037
R1680 VN.n4 VN.n1 80.6037
R1681 VN VN.n19 49.7524
R1682 VN.n2 VN.n1 48.2005
R1683 VN.n6 VN.n1 48.2005
R1684 VN.n12 VN.n11 48.2005
R1685 VN.n16 VN.n11 48.2005
R1686 VN.n14 VN.n13 31.9326
R1687 VN.n4 VN.n3 31.9326
R1688 VN.n7 VN.n6 29.9429
R1689 VN.n17 VN.n16 29.9429
R1690 VN.n8 VN.n7 18.2581
R1691 VN.n18 VN.n17 18.2581
R1692 VN.n3 VN.n2 15.8785
R1693 VN.n13 VN.n12 15.8785
R1694 VN.n15 VN.n14 0.380177
R1695 VN.n5 VN.n4 0.380177
R1696 VN.n15 VN.n10 0.285035
R1697 VN.n5 VN.n0 0.285035
R1698 VN.n19 VN.n10 0.189894
R1699 VN.n9 VN.n0 0.189894
R1700 VN VN.n9 0.0516364
R1701 VTAIL.n11 VTAIL.t12 48.7877
R1702 VTAIL.n17 VTAIL.t13 48.7875
R1703 VTAIL.n2 VTAIL.t6 48.7875
R1704 VTAIL.n16 VTAIL.t5 48.7875
R1705 VTAIL.n15 VTAIL.n14 47.7927
R1706 VTAIL.n13 VTAIL.n12 47.7927
R1707 VTAIL.n10 VTAIL.n9 47.7927
R1708 VTAIL.n8 VTAIL.n7 47.7927
R1709 VTAIL.n19 VTAIL.n18 47.7925
R1710 VTAIL.n1 VTAIL.n0 47.7925
R1711 VTAIL.n4 VTAIL.n3 47.7925
R1712 VTAIL.n6 VTAIL.n5 47.7925
R1713 VTAIL.n8 VTAIL.n6 31.4876
R1714 VTAIL.n17 VTAIL.n16 30.5048
R1715 VTAIL.n18 VTAIL.t11 0.995475
R1716 VTAIL.n18 VTAIL.t18 0.995475
R1717 VTAIL.n0 VTAIL.t17 0.995475
R1718 VTAIL.n0 VTAIL.t15 0.995475
R1719 VTAIL.n3 VTAIL.t19 0.995475
R1720 VTAIL.n3 VTAIL.t7 0.995475
R1721 VTAIL.n5 VTAIL.t0 0.995475
R1722 VTAIL.n5 VTAIL.t8 0.995475
R1723 VTAIL.n14 VTAIL.t4 0.995475
R1724 VTAIL.n14 VTAIL.t1 0.995475
R1725 VTAIL.n12 VTAIL.t2 0.995475
R1726 VTAIL.n12 VTAIL.t3 0.995475
R1727 VTAIL.n9 VTAIL.t14 0.995475
R1728 VTAIL.n9 VTAIL.t9 0.995475
R1729 VTAIL.n7 VTAIL.t10 0.995475
R1730 VTAIL.n7 VTAIL.t16 0.995475
R1731 VTAIL.n10 VTAIL.n8 0.983259
R1732 VTAIL.n11 VTAIL.n10 0.983259
R1733 VTAIL.n15 VTAIL.n13 0.983259
R1734 VTAIL.n16 VTAIL.n15 0.983259
R1735 VTAIL.n6 VTAIL.n4 0.983259
R1736 VTAIL.n4 VTAIL.n2 0.983259
R1737 VTAIL.n19 VTAIL.n17 0.983259
R1738 VTAIL.n13 VTAIL.n11 0.961707
R1739 VTAIL.n2 VTAIL.n1 0.961707
R1740 VTAIL VTAIL.n1 0.795759
R1741 VTAIL VTAIL.n19 0.188
R1742 VDD2.n1 VDD2.t8 66.449
R1743 VDD2.n4 VDD2.t9 65.4665
R1744 VDD2.n3 VDD2.n2 65.153
R1745 VDD2 VDD2.n7 65.1502
R1746 VDD2.n6 VDD2.n5 64.4715
R1747 VDD2.n1 VDD2.n0 64.4713
R1748 VDD2.n4 VDD2.n3 45.5386
R1749 VDD2.n7 VDD2.t0 0.995475
R1750 VDD2.n7 VDD2.t4 0.995475
R1751 VDD2.n5 VDD2.t3 0.995475
R1752 VDD2.n5 VDD2.t7 0.995475
R1753 VDD2.n2 VDD2.t5 0.995475
R1754 VDD2.n2 VDD2.t6 0.995475
R1755 VDD2.n0 VDD2.t1 0.995475
R1756 VDD2.n0 VDD2.t2 0.995475
R1757 VDD2.n6 VDD2.n4 0.983259
R1758 VDD2 VDD2.n6 0.304379
R1759 VDD2.n3 VDD2.n1 0.190844
R1760 VP.n6 VP.t2 664.332
R1761 VP.n14 VP.t8 640.585
R1762 VP.n16 VP.t3 640.585
R1763 VP.n1 VP.t1 640.585
R1764 VP.n20 VP.t4 640.585
R1765 VP.n22 VP.t7 640.585
R1766 VP.n11 VP.t6 640.585
R1767 VP.n9 VP.t0 640.585
R1768 VP.n8 VP.t9 640.585
R1769 VP.n7 VP.t5 640.585
R1770 VP.n23 VP.n22 161.3
R1771 VP.n10 VP.n3 161.3
R1772 VP.n12 VP.n11 161.3
R1773 VP.n21 VP.n0 161.3
R1774 VP.n15 VP.n2 161.3
R1775 VP.n14 VP.n13 161.3
R1776 VP.n8 VP.n5 80.6037
R1777 VP.n9 VP.n4 80.6037
R1778 VP.n20 VP.n19 80.6037
R1779 VP.n18 VP.n1 80.6037
R1780 VP.n17 VP.n16 80.6037
R1781 VP.n13 VP.n12 49.3717
R1782 VP.n16 VP.n1 48.2005
R1783 VP.n20 VP.n1 48.2005
R1784 VP.n9 VP.n8 48.2005
R1785 VP.n8 VP.n7 48.2005
R1786 VP.n6 VP.n5 31.9325
R1787 VP.n16 VP.n15 29.9429
R1788 VP.n21 VP.n20 29.9429
R1789 VP.n10 VP.n9 29.9429
R1790 VP.n15 VP.n14 18.2581
R1791 VP.n22 VP.n21 18.2581
R1792 VP.n11 VP.n10 18.2581
R1793 VP.n7 VP.n6 15.8785
R1794 VP.n5 VP.n4 0.380177
R1795 VP.n18 VP.n17 0.380177
R1796 VP.n19 VP.n18 0.380177
R1797 VP.n4 VP.n3 0.285035
R1798 VP.n17 VP.n2 0.285035
R1799 VP.n19 VP.n0 0.285035
R1800 VP.n12 VP.n3 0.189894
R1801 VP.n13 VP.n2 0.189894
R1802 VP.n23 VP.n0 0.189894
R1803 VP VP.n23 0.0516364
R1804 VDD1.n1 VDD1.t7 66.4492
R1805 VDD1.n3 VDD1.t1 66.449
R1806 VDD1.n5 VDD1.n4 65.153
R1807 VDD1.n1 VDD1.n0 64.4715
R1808 VDD1.n7 VDD1.n6 64.4713
R1809 VDD1.n3 VDD1.n2 64.4713
R1810 VDD1.n7 VDD1.n5 46.613
R1811 VDD1.n6 VDD1.t9 0.995475
R1812 VDD1.n6 VDD1.t3 0.995475
R1813 VDD1.n0 VDD1.t4 0.995475
R1814 VDD1.n0 VDD1.t0 0.995475
R1815 VDD1.n4 VDD1.t5 0.995475
R1816 VDD1.n4 VDD1.t2 0.995475
R1817 VDD1.n2 VDD1.t6 0.995475
R1818 VDD1.n2 VDD1.t8 0.995475
R1819 VDD1 VDD1.n7 0.679379
R1820 VDD1 VDD1.n1 0.304379
R1821 VDD1.n5 VDD1.n3 0.190844
C0 VTAIL VDD1 20.413198f
C1 VN VTAIL 11.252f
C2 VDD2 VP 0.356943f
C3 VDD2 VDD1 1.0428f
C4 VP VDD1 11.8641f
C5 VN VDD2 11.663799f
C6 VN VP 7.21879f
C7 VN VDD1 0.149501f
C8 VDD2 VTAIL 20.4444f
C9 VTAIL VP 11.266799f
C10 VDD2 B 6.500072f
C11 VDD1 B 6.440493f
C12 VTAIL B 9.511022f
C13 VN B 10.83175f
C14 VP B 8.561701f
C15 VDD1.t7 B 4.42032f
C16 VDD1.t4 B 0.376385f
C17 VDD1.t0 B 0.376385f
C18 VDD1.n0 B 3.45113f
C19 VDD1.n1 B 0.624229f
C20 VDD1.t1 B 4.42032f
C21 VDD1.t6 B 0.376385f
C22 VDD1.t8 B 0.376385f
C23 VDD1.n2 B 3.45114f
C24 VDD1.n3 B 0.618388f
C25 VDD1.t5 B 0.376385f
C26 VDD1.t2 B 0.376385f
C27 VDD1.n4 B 3.45459f
C28 VDD1.n5 B 2.42122f
C29 VDD1.t9 B 0.376385f
C30 VDD1.t3 B 0.376385f
C31 VDD1.n6 B 3.45113f
C32 VDD1.n7 B 2.90067f
C33 VP.n0 B 0.0538f
C34 VP.t1 B 1.84054f
C35 VP.n1 B 0.69527f
C36 VP.n2 B 0.0538f
C37 VP.n3 B 0.0538f
C38 VP.t6 B 1.84054f
C39 VP.t0 B 1.84054f
C40 VP.n4 B 0.067156f
C41 VP.t9 B 1.84054f
C42 VP.n5 B 0.248648f
C43 VP.t5 B 1.84054f
C44 VP.t2 B 1.86506f
C45 VP.n6 B 0.666072f
C46 VP.n7 B 0.69421f
C47 VP.n8 B 0.69527f
C48 VP.n9 B 0.692162f
C49 VP.n10 B 0.009149f
C50 VP.n11 B 0.681025f
C51 VP.n12 B 2.15055f
C52 VP.n13 B 2.17999f
C53 VP.t8 B 1.84054f
C54 VP.n14 B 0.681025f
C55 VP.n15 B 0.009149f
C56 VP.t3 B 1.84054f
C57 VP.n16 B 0.692162f
C58 VP.n17 B 0.067156f
C59 VP.n18 B 0.080638f
C60 VP.n19 B 0.067156f
C61 VP.t4 B 1.84054f
C62 VP.n20 B 0.692162f
C63 VP.n21 B 0.009149f
C64 VP.t7 B 1.84054f
C65 VP.n22 B 0.681025f
C66 VP.n23 B 0.031246f
C67 VDD2.t8 B 4.405f
C68 VDD2.t1 B 0.375081f
C69 VDD2.t2 B 0.375081f
C70 VDD2.n0 B 3.43918f
C71 VDD2.n1 B 0.616246f
C72 VDD2.t5 B 0.375081f
C73 VDD2.t6 B 0.375081f
C74 VDD2.n2 B 3.44262f
C75 VDD2.n3 B 2.33489f
C76 VDD2.t9 B 4.40001f
C77 VDD2.n4 B 2.8904f
C78 VDD2.t3 B 0.375081f
C79 VDD2.t7 B 0.375081f
C80 VDD2.n5 B 3.43918f
C81 VDD2.n6 B 0.289346f
C82 VDD2.t0 B 0.375081f
C83 VDD2.t4 B 0.375081f
C84 VDD2.n7 B 3.44259f
C85 VTAIL.t17 B 0.384874f
C86 VTAIL.t15 B 0.384874f
C87 VTAIL.n0 B 3.4624f
C88 VTAIL.n1 B 0.367265f
C89 VTAIL.t6 B 4.42788f
C90 VTAIL.n2 B 0.466223f
C91 VTAIL.t19 B 0.384874f
C92 VTAIL.t7 B 0.384874f
C93 VTAIL.n3 B 3.4624f
C94 VTAIL.n4 B 0.383751f
C95 VTAIL.t0 B 0.384874f
C96 VTAIL.t8 B 0.384874f
C97 VTAIL.n5 B 3.4624f
C98 VTAIL.n6 B 2.1466f
C99 VTAIL.t10 B 0.384874f
C100 VTAIL.t16 B 0.384874f
C101 VTAIL.n7 B 3.4624f
C102 VTAIL.n8 B 2.1466f
C103 VTAIL.t14 B 0.384874f
C104 VTAIL.t9 B 0.384874f
C105 VTAIL.n9 B 3.4624f
C106 VTAIL.n10 B 0.383751f
C107 VTAIL.t12 B 4.42788f
C108 VTAIL.n11 B 0.466222f
C109 VTAIL.t2 B 0.384874f
C110 VTAIL.t3 B 0.384874f
C111 VTAIL.n12 B 3.4624f
C112 VTAIL.n13 B 0.382052f
C113 VTAIL.t4 B 0.384874f
C114 VTAIL.t1 B 0.384874f
C115 VTAIL.n14 B 3.4624f
C116 VTAIL.n15 B 0.383751f
C117 VTAIL.t5 B 4.42788f
C118 VTAIL.n16 B 2.15327f
C119 VTAIL.t13 B 4.42788f
C120 VTAIL.n17 B 2.15327f
C121 VTAIL.t11 B 0.384874f
C122 VTAIL.t18 B 0.384874f
C123 VTAIL.n18 B 3.4624f
C124 VTAIL.n19 B 0.321036f
C125 VN.n0 B 0.053347f
C126 VN.t7 B 1.82503f
C127 VN.n1 B 0.68941f
C128 VN.t1 B 1.84934f
C129 VN.t8 B 1.82503f
C130 VN.n2 B 0.68836f
C131 VN.n3 B 0.660459f
C132 VN.n4 B 0.246552f
C133 VN.n5 B 0.06659f
C134 VN.t4 B 1.82503f
C135 VN.n6 B 0.686329f
C136 VN.n7 B 0.009072f
C137 VN.t3 B 1.82503f
C138 VN.n8 B 0.675285f
C139 VN.n9 B 0.030982f
C140 VN.n10 B 0.053347f
C141 VN.t2 B 1.82503f
C142 VN.n11 B 0.68941f
C143 VN.t6 B 1.82503f
C144 VN.t5 B 1.84934f
C145 VN.t9 B 1.82503f
C146 VN.n12 B 0.68836f
C147 VN.n13 B 0.660459f
C148 VN.n14 B 0.246552f
C149 VN.n15 B 0.06659f
C150 VN.n16 B 0.686329f
C151 VN.n17 B 0.009072f
C152 VN.t0 B 1.82503f
C153 VN.n18 B 0.675285f
C154 VN.n19 B 2.15843f
.ends

