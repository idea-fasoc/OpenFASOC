* NGSPICE file created from diff_pair_sample_0895.ext - technology: sky130A

.subckt diff_pair_sample_0895 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=0 ps=0 w=9.8 l=3.87
X1 VDD1.t5 VP.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=1.617 ps=10.13 w=9.8 l=3.87
X2 VTAIL.t9 VP.t1 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=1.617 ps=10.13 w=9.8 l=3.87
X3 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=1.617 ps=10.13 w=9.8 l=3.87
X4 VTAIL.t4 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=1.617 ps=10.13 w=9.8 l=3.87
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=0 ps=0 w=9.8 l=3.87
X6 VDD1.t3 VP.t2 VTAIL.t8 B.t19 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=3.822 ps=20.38 w=9.8 l=3.87
X7 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=0 ps=0 w=9.8 l=3.87
X8 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=1.617 ps=10.13 w=9.8 l=3.87
X9 VDD1.t2 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=3.822 ps=20.38 w=9.8 l=3.87
X10 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=0 ps=0 w=9.8 l=3.87
X11 VDD1.t1 VP.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.822 pd=20.38 as=1.617 ps=10.13 w=9.8 l=3.87
X12 VDD2.t2 VN.t3 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=3.822 ps=20.38 w=9.8 l=3.87
X13 VTAIL.t10 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=1.617 ps=10.13 w=9.8 l=3.87
X14 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=1.617 ps=10.13 w=9.8 l=3.87
X15 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.617 pd=10.13 as=3.822 ps=20.38 w=9.8 l=3.87
R0 B.n872 B.n871 585
R1 B.n308 B.n145 585
R2 B.n307 B.n306 585
R3 B.n305 B.n304 585
R4 B.n303 B.n302 585
R5 B.n301 B.n300 585
R6 B.n299 B.n298 585
R7 B.n297 B.n296 585
R8 B.n295 B.n294 585
R9 B.n293 B.n292 585
R10 B.n291 B.n290 585
R11 B.n289 B.n288 585
R12 B.n287 B.n286 585
R13 B.n285 B.n284 585
R14 B.n283 B.n282 585
R15 B.n281 B.n280 585
R16 B.n279 B.n278 585
R17 B.n277 B.n276 585
R18 B.n275 B.n274 585
R19 B.n273 B.n272 585
R20 B.n271 B.n270 585
R21 B.n269 B.n268 585
R22 B.n267 B.n266 585
R23 B.n265 B.n264 585
R24 B.n263 B.n262 585
R25 B.n261 B.n260 585
R26 B.n259 B.n258 585
R27 B.n257 B.n256 585
R28 B.n255 B.n254 585
R29 B.n253 B.n252 585
R30 B.n251 B.n250 585
R31 B.n249 B.n248 585
R32 B.n247 B.n246 585
R33 B.n245 B.n244 585
R34 B.n243 B.n242 585
R35 B.n240 B.n239 585
R36 B.n238 B.n237 585
R37 B.n236 B.n235 585
R38 B.n234 B.n233 585
R39 B.n232 B.n231 585
R40 B.n230 B.n229 585
R41 B.n228 B.n227 585
R42 B.n226 B.n225 585
R43 B.n224 B.n223 585
R44 B.n222 B.n221 585
R45 B.n219 B.n218 585
R46 B.n217 B.n216 585
R47 B.n215 B.n214 585
R48 B.n213 B.n212 585
R49 B.n211 B.n210 585
R50 B.n209 B.n208 585
R51 B.n207 B.n206 585
R52 B.n205 B.n204 585
R53 B.n203 B.n202 585
R54 B.n201 B.n200 585
R55 B.n199 B.n198 585
R56 B.n197 B.n196 585
R57 B.n195 B.n194 585
R58 B.n193 B.n192 585
R59 B.n191 B.n190 585
R60 B.n189 B.n188 585
R61 B.n187 B.n186 585
R62 B.n185 B.n184 585
R63 B.n183 B.n182 585
R64 B.n181 B.n180 585
R65 B.n179 B.n178 585
R66 B.n177 B.n176 585
R67 B.n175 B.n174 585
R68 B.n173 B.n172 585
R69 B.n171 B.n170 585
R70 B.n169 B.n168 585
R71 B.n167 B.n166 585
R72 B.n165 B.n164 585
R73 B.n163 B.n162 585
R74 B.n161 B.n160 585
R75 B.n159 B.n158 585
R76 B.n157 B.n156 585
R77 B.n155 B.n154 585
R78 B.n153 B.n152 585
R79 B.n151 B.n150 585
R80 B.n870 B.n105 585
R81 B.n875 B.n105 585
R82 B.n869 B.n104 585
R83 B.n876 B.n104 585
R84 B.n868 B.n867 585
R85 B.n867 B.n100 585
R86 B.n866 B.n99 585
R87 B.n882 B.n99 585
R88 B.n865 B.n98 585
R89 B.n883 B.n98 585
R90 B.n864 B.n97 585
R91 B.n884 B.n97 585
R92 B.n863 B.n862 585
R93 B.n862 B.n93 585
R94 B.n861 B.n92 585
R95 B.n890 B.n92 585
R96 B.n860 B.n91 585
R97 B.n891 B.n91 585
R98 B.n859 B.n90 585
R99 B.n892 B.n90 585
R100 B.n858 B.n857 585
R101 B.n857 B.n86 585
R102 B.n856 B.n85 585
R103 B.n898 B.n85 585
R104 B.n855 B.n84 585
R105 B.n899 B.n84 585
R106 B.n854 B.n83 585
R107 B.n900 B.n83 585
R108 B.n853 B.n852 585
R109 B.n852 B.n79 585
R110 B.n851 B.n78 585
R111 B.n906 B.n78 585
R112 B.n850 B.n77 585
R113 B.n907 B.n77 585
R114 B.n849 B.n76 585
R115 B.n908 B.n76 585
R116 B.n848 B.n847 585
R117 B.n847 B.n72 585
R118 B.n846 B.n71 585
R119 B.n914 B.n71 585
R120 B.n845 B.n70 585
R121 B.n915 B.n70 585
R122 B.n844 B.n69 585
R123 B.n916 B.n69 585
R124 B.n843 B.n842 585
R125 B.n842 B.n65 585
R126 B.n841 B.n64 585
R127 B.n922 B.n64 585
R128 B.n840 B.n63 585
R129 B.n923 B.n63 585
R130 B.n839 B.n62 585
R131 B.n924 B.n62 585
R132 B.n838 B.n837 585
R133 B.n837 B.n58 585
R134 B.n836 B.n57 585
R135 B.n930 B.n57 585
R136 B.n835 B.n56 585
R137 B.n931 B.n56 585
R138 B.n834 B.n55 585
R139 B.n932 B.n55 585
R140 B.n833 B.n832 585
R141 B.n832 B.n51 585
R142 B.n831 B.n50 585
R143 B.n938 B.n50 585
R144 B.n830 B.n49 585
R145 B.n939 B.n49 585
R146 B.n829 B.n48 585
R147 B.n940 B.n48 585
R148 B.n828 B.n827 585
R149 B.n827 B.n44 585
R150 B.n826 B.n43 585
R151 B.n946 B.n43 585
R152 B.n825 B.n42 585
R153 B.n947 B.n42 585
R154 B.n824 B.n41 585
R155 B.n948 B.n41 585
R156 B.n823 B.n822 585
R157 B.n822 B.n37 585
R158 B.n821 B.n36 585
R159 B.n954 B.n36 585
R160 B.n820 B.n35 585
R161 B.n955 B.n35 585
R162 B.n819 B.n34 585
R163 B.n956 B.n34 585
R164 B.n818 B.n817 585
R165 B.n817 B.n30 585
R166 B.n816 B.n29 585
R167 B.n962 B.n29 585
R168 B.n815 B.n28 585
R169 B.n963 B.n28 585
R170 B.n814 B.n27 585
R171 B.n964 B.n27 585
R172 B.n813 B.n812 585
R173 B.n812 B.n23 585
R174 B.n811 B.n22 585
R175 B.n970 B.n22 585
R176 B.n810 B.n21 585
R177 B.n971 B.n21 585
R178 B.n809 B.n20 585
R179 B.n972 B.n20 585
R180 B.n808 B.n807 585
R181 B.n807 B.n16 585
R182 B.n806 B.n15 585
R183 B.n978 B.n15 585
R184 B.n805 B.n14 585
R185 B.n979 B.n14 585
R186 B.n804 B.n13 585
R187 B.n980 B.n13 585
R188 B.n803 B.n802 585
R189 B.n802 B.n12 585
R190 B.n801 B.n800 585
R191 B.n801 B.n8 585
R192 B.n799 B.n7 585
R193 B.n987 B.n7 585
R194 B.n798 B.n6 585
R195 B.n988 B.n6 585
R196 B.n797 B.n5 585
R197 B.n989 B.n5 585
R198 B.n796 B.n795 585
R199 B.n795 B.n4 585
R200 B.n794 B.n309 585
R201 B.n794 B.n793 585
R202 B.n784 B.n310 585
R203 B.n311 B.n310 585
R204 B.n786 B.n785 585
R205 B.n787 B.n786 585
R206 B.n783 B.n316 585
R207 B.n316 B.n315 585
R208 B.n782 B.n781 585
R209 B.n781 B.n780 585
R210 B.n318 B.n317 585
R211 B.n319 B.n318 585
R212 B.n773 B.n772 585
R213 B.n774 B.n773 585
R214 B.n771 B.n324 585
R215 B.n324 B.n323 585
R216 B.n770 B.n769 585
R217 B.n769 B.n768 585
R218 B.n326 B.n325 585
R219 B.n327 B.n326 585
R220 B.n761 B.n760 585
R221 B.n762 B.n761 585
R222 B.n759 B.n332 585
R223 B.n332 B.n331 585
R224 B.n758 B.n757 585
R225 B.n757 B.n756 585
R226 B.n334 B.n333 585
R227 B.n335 B.n334 585
R228 B.n749 B.n748 585
R229 B.n750 B.n749 585
R230 B.n747 B.n340 585
R231 B.n340 B.n339 585
R232 B.n746 B.n745 585
R233 B.n745 B.n744 585
R234 B.n342 B.n341 585
R235 B.n343 B.n342 585
R236 B.n737 B.n736 585
R237 B.n738 B.n737 585
R238 B.n735 B.n348 585
R239 B.n348 B.n347 585
R240 B.n734 B.n733 585
R241 B.n733 B.n732 585
R242 B.n350 B.n349 585
R243 B.n351 B.n350 585
R244 B.n725 B.n724 585
R245 B.n726 B.n725 585
R246 B.n723 B.n356 585
R247 B.n356 B.n355 585
R248 B.n722 B.n721 585
R249 B.n721 B.n720 585
R250 B.n358 B.n357 585
R251 B.n359 B.n358 585
R252 B.n713 B.n712 585
R253 B.n714 B.n713 585
R254 B.n711 B.n364 585
R255 B.n364 B.n363 585
R256 B.n710 B.n709 585
R257 B.n709 B.n708 585
R258 B.n366 B.n365 585
R259 B.n367 B.n366 585
R260 B.n701 B.n700 585
R261 B.n702 B.n701 585
R262 B.n699 B.n372 585
R263 B.n372 B.n371 585
R264 B.n698 B.n697 585
R265 B.n697 B.n696 585
R266 B.n374 B.n373 585
R267 B.n375 B.n374 585
R268 B.n689 B.n688 585
R269 B.n690 B.n689 585
R270 B.n687 B.n380 585
R271 B.n380 B.n379 585
R272 B.n686 B.n685 585
R273 B.n685 B.n684 585
R274 B.n382 B.n381 585
R275 B.n383 B.n382 585
R276 B.n677 B.n676 585
R277 B.n678 B.n677 585
R278 B.n675 B.n388 585
R279 B.n388 B.n387 585
R280 B.n674 B.n673 585
R281 B.n673 B.n672 585
R282 B.n390 B.n389 585
R283 B.n391 B.n390 585
R284 B.n665 B.n664 585
R285 B.n666 B.n665 585
R286 B.n663 B.n396 585
R287 B.n396 B.n395 585
R288 B.n662 B.n661 585
R289 B.n661 B.n660 585
R290 B.n398 B.n397 585
R291 B.n399 B.n398 585
R292 B.n653 B.n652 585
R293 B.n654 B.n653 585
R294 B.n651 B.n404 585
R295 B.n404 B.n403 585
R296 B.n650 B.n649 585
R297 B.n649 B.n648 585
R298 B.n406 B.n405 585
R299 B.n407 B.n406 585
R300 B.n641 B.n640 585
R301 B.n642 B.n641 585
R302 B.n639 B.n412 585
R303 B.n412 B.n411 585
R304 B.n638 B.n637 585
R305 B.n637 B.n636 585
R306 B.n414 B.n413 585
R307 B.n415 B.n414 585
R308 B.n629 B.n628 585
R309 B.n630 B.n629 585
R310 B.n627 B.n420 585
R311 B.n420 B.n419 585
R312 B.n622 B.n621 585
R313 B.n620 B.n462 585
R314 B.n619 B.n461 585
R315 B.n624 B.n461 585
R316 B.n618 B.n617 585
R317 B.n616 B.n615 585
R318 B.n614 B.n613 585
R319 B.n612 B.n611 585
R320 B.n610 B.n609 585
R321 B.n608 B.n607 585
R322 B.n606 B.n605 585
R323 B.n604 B.n603 585
R324 B.n602 B.n601 585
R325 B.n600 B.n599 585
R326 B.n598 B.n597 585
R327 B.n596 B.n595 585
R328 B.n594 B.n593 585
R329 B.n592 B.n591 585
R330 B.n590 B.n589 585
R331 B.n588 B.n587 585
R332 B.n586 B.n585 585
R333 B.n584 B.n583 585
R334 B.n582 B.n581 585
R335 B.n580 B.n579 585
R336 B.n578 B.n577 585
R337 B.n576 B.n575 585
R338 B.n574 B.n573 585
R339 B.n572 B.n571 585
R340 B.n570 B.n569 585
R341 B.n568 B.n567 585
R342 B.n566 B.n565 585
R343 B.n564 B.n563 585
R344 B.n562 B.n561 585
R345 B.n560 B.n559 585
R346 B.n558 B.n557 585
R347 B.n556 B.n555 585
R348 B.n554 B.n553 585
R349 B.n552 B.n551 585
R350 B.n550 B.n549 585
R351 B.n548 B.n547 585
R352 B.n546 B.n545 585
R353 B.n544 B.n543 585
R354 B.n542 B.n541 585
R355 B.n540 B.n539 585
R356 B.n538 B.n537 585
R357 B.n536 B.n535 585
R358 B.n534 B.n533 585
R359 B.n532 B.n531 585
R360 B.n530 B.n529 585
R361 B.n528 B.n527 585
R362 B.n526 B.n525 585
R363 B.n524 B.n523 585
R364 B.n522 B.n521 585
R365 B.n520 B.n519 585
R366 B.n518 B.n517 585
R367 B.n516 B.n515 585
R368 B.n514 B.n513 585
R369 B.n512 B.n511 585
R370 B.n510 B.n509 585
R371 B.n508 B.n507 585
R372 B.n506 B.n505 585
R373 B.n504 B.n503 585
R374 B.n502 B.n501 585
R375 B.n500 B.n499 585
R376 B.n498 B.n497 585
R377 B.n496 B.n495 585
R378 B.n494 B.n493 585
R379 B.n492 B.n491 585
R380 B.n490 B.n489 585
R381 B.n488 B.n487 585
R382 B.n486 B.n485 585
R383 B.n484 B.n483 585
R384 B.n482 B.n481 585
R385 B.n480 B.n479 585
R386 B.n478 B.n477 585
R387 B.n476 B.n475 585
R388 B.n474 B.n473 585
R389 B.n472 B.n471 585
R390 B.n470 B.n469 585
R391 B.n422 B.n421 585
R392 B.n626 B.n625 585
R393 B.n625 B.n624 585
R394 B.n418 B.n417 585
R395 B.n419 B.n418 585
R396 B.n632 B.n631 585
R397 B.n631 B.n630 585
R398 B.n633 B.n416 585
R399 B.n416 B.n415 585
R400 B.n635 B.n634 585
R401 B.n636 B.n635 585
R402 B.n410 B.n409 585
R403 B.n411 B.n410 585
R404 B.n644 B.n643 585
R405 B.n643 B.n642 585
R406 B.n645 B.n408 585
R407 B.n408 B.n407 585
R408 B.n647 B.n646 585
R409 B.n648 B.n647 585
R410 B.n402 B.n401 585
R411 B.n403 B.n402 585
R412 B.n656 B.n655 585
R413 B.n655 B.n654 585
R414 B.n657 B.n400 585
R415 B.n400 B.n399 585
R416 B.n659 B.n658 585
R417 B.n660 B.n659 585
R418 B.n394 B.n393 585
R419 B.n395 B.n394 585
R420 B.n668 B.n667 585
R421 B.n667 B.n666 585
R422 B.n669 B.n392 585
R423 B.n392 B.n391 585
R424 B.n671 B.n670 585
R425 B.n672 B.n671 585
R426 B.n386 B.n385 585
R427 B.n387 B.n386 585
R428 B.n680 B.n679 585
R429 B.n679 B.n678 585
R430 B.n681 B.n384 585
R431 B.n384 B.n383 585
R432 B.n683 B.n682 585
R433 B.n684 B.n683 585
R434 B.n378 B.n377 585
R435 B.n379 B.n378 585
R436 B.n692 B.n691 585
R437 B.n691 B.n690 585
R438 B.n693 B.n376 585
R439 B.n376 B.n375 585
R440 B.n695 B.n694 585
R441 B.n696 B.n695 585
R442 B.n370 B.n369 585
R443 B.n371 B.n370 585
R444 B.n704 B.n703 585
R445 B.n703 B.n702 585
R446 B.n705 B.n368 585
R447 B.n368 B.n367 585
R448 B.n707 B.n706 585
R449 B.n708 B.n707 585
R450 B.n362 B.n361 585
R451 B.n363 B.n362 585
R452 B.n716 B.n715 585
R453 B.n715 B.n714 585
R454 B.n717 B.n360 585
R455 B.n360 B.n359 585
R456 B.n719 B.n718 585
R457 B.n720 B.n719 585
R458 B.n354 B.n353 585
R459 B.n355 B.n354 585
R460 B.n728 B.n727 585
R461 B.n727 B.n726 585
R462 B.n729 B.n352 585
R463 B.n352 B.n351 585
R464 B.n731 B.n730 585
R465 B.n732 B.n731 585
R466 B.n346 B.n345 585
R467 B.n347 B.n346 585
R468 B.n740 B.n739 585
R469 B.n739 B.n738 585
R470 B.n741 B.n344 585
R471 B.n344 B.n343 585
R472 B.n743 B.n742 585
R473 B.n744 B.n743 585
R474 B.n338 B.n337 585
R475 B.n339 B.n338 585
R476 B.n752 B.n751 585
R477 B.n751 B.n750 585
R478 B.n753 B.n336 585
R479 B.n336 B.n335 585
R480 B.n755 B.n754 585
R481 B.n756 B.n755 585
R482 B.n330 B.n329 585
R483 B.n331 B.n330 585
R484 B.n764 B.n763 585
R485 B.n763 B.n762 585
R486 B.n765 B.n328 585
R487 B.n328 B.n327 585
R488 B.n767 B.n766 585
R489 B.n768 B.n767 585
R490 B.n322 B.n321 585
R491 B.n323 B.n322 585
R492 B.n776 B.n775 585
R493 B.n775 B.n774 585
R494 B.n777 B.n320 585
R495 B.n320 B.n319 585
R496 B.n779 B.n778 585
R497 B.n780 B.n779 585
R498 B.n314 B.n313 585
R499 B.n315 B.n314 585
R500 B.n789 B.n788 585
R501 B.n788 B.n787 585
R502 B.n790 B.n312 585
R503 B.n312 B.n311 585
R504 B.n792 B.n791 585
R505 B.n793 B.n792 585
R506 B.n3 B.n0 585
R507 B.n4 B.n3 585
R508 B.n986 B.n1 585
R509 B.n987 B.n986 585
R510 B.n985 B.n984 585
R511 B.n985 B.n8 585
R512 B.n983 B.n9 585
R513 B.n12 B.n9 585
R514 B.n982 B.n981 585
R515 B.n981 B.n980 585
R516 B.n11 B.n10 585
R517 B.n979 B.n11 585
R518 B.n977 B.n976 585
R519 B.n978 B.n977 585
R520 B.n975 B.n17 585
R521 B.n17 B.n16 585
R522 B.n974 B.n973 585
R523 B.n973 B.n972 585
R524 B.n19 B.n18 585
R525 B.n971 B.n19 585
R526 B.n969 B.n968 585
R527 B.n970 B.n969 585
R528 B.n967 B.n24 585
R529 B.n24 B.n23 585
R530 B.n966 B.n965 585
R531 B.n965 B.n964 585
R532 B.n26 B.n25 585
R533 B.n963 B.n26 585
R534 B.n961 B.n960 585
R535 B.n962 B.n961 585
R536 B.n959 B.n31 585
R537 B.n31 B.n30 585
R538 B.n958 B.n957 585
R539 B.n957 B.n956 585
R540 B.n33 B.n32 585
R541 B.n955 B.n33 585
R542 B.n953 B.n952 585
R543 B.n954 B.n953 585
R544 B.n951 B.n38 585
R545 B.n38 B.n37 585
R546 B.n950 B.n949 585
R547 B.n949 B.n948 585
R548 B.n40 B.n39 585
R549 B.n947 B.n40 585
R550 B.n945 B.n944 585
R551 B.n946 B.n945 585
R552 B.n943 B.n45 585
R553 B.n45 B.n44 585
R554 B.n942 B.n941 585
R555 B.n941 B.n940 585
R556 B.n47 B.n46 585
R557 B.n939 B.n47 585
R558 B.n937 B.n936 585
R559 B.n938 B.n937 585
R560 B.n935 B.n52 585
R561 B.n52 B.n51 585
R562 B.n934 B.n933 585
R563 B.n933 B.n932 585
R564 B.n54 B.n53 585
R565 B.n931 B.n54 585
R566 B.n929 B.n928 585
R567 B.n930 B.n929 585
R568 B.n927 B.n59 585
R569 B.n59 B.n58 585
R570 B.n926 B.n925 585
R571 B.n925 B.n924 585
R572 B.n61 B.n60 585
R573 B.n923 B.n61 585
R574 B.n921 B.n920 585
R575 B.n922 B.n921 585
R576 B.n919 B.n66 585
R577 B.n66 B.n65 585
R578 B.n918 B.n917 585
R579 B.n917 B.n916 585
R580 B.n68 B.n67 585
R581 B.n915 B.n68 585
R582 B.n913 B.n912 585
R583 B.n914 B.n913 585
R584 B.n911 B.n73 585
R585 B.n73 B.n72 585
R586 B.n910 B.n909 585
R587 B.n909 B.n908 585
R588 B.n75 B.n74 585
R589 B.n907 B.n75 585
R590 B.n905 B.n904 585
R591 B.n906 B.n905 585
R592 B.n903 B.n80 585
R593 B.n80 B.n79 585
R594 B.n902 B.n901 585
R595 B.n901 B.n900 585
R596 B.n82 B.n81 585
R597 B.n899 B.n82 585
R598 B.n897 B.n896 585
R599 B.n898 B.n897 585
R600 B.n895 B.n87 585
R601 B.n87 B.n86 585
R602 B.n894 B.n893 585
R603 B.n893 B.n892 585
R604 B.n89 B.n88 585
R605 B.n891 B.n89 585
R606 B.n889 B.n888 585
R607 B.n890 B.n889 585
R608 B.n887 B.n94 585
R609 B.n94 B.n93 585
R610 B.n886 B.n885 585
R611 B.n885 B.n884 585
R612 B.n96 B.n95 585
R613 B.n883 B.n96 585
R614 B.n881 B.n880 585
R615 B.n882 B.n881 585
R616 B.n879 B.n101 585
R617 B.n101 B.n100 585
R618 B.n878 B.n877 585
R619 B.n877 B.n876 585
R620 B.n103 B.n102 585
R621 B.n875 B.n103 585
R622 B.n990 B.n989 585
R623 B.n988 B.n2 585
R624 B.n150 B.n103 492.5
R625 B.n872 B.n105 492.5
R626 B.n625 B.n420 492.5
R627 B.n622 B.n418 492.5
R628 B.n148 B.t5 270.425
R629 B.n146 B.t9 270.425
R630 B.n466 B.t12 270.425
R631 B.n463 B.t16 270.425
R632 B.n874 B.n873 256.663
R633 B.n874 B.n144 256.663
R634 B.n874 B.n143 256.663
R635 B.n874 B.n142 256.663
R636 B.n874 B.n141 256.663
R637 B.n874 B.n140 256.663
R638 B.n874 B.n139 256.663
R639 B.n874 B.n138 256.663
R640 B.n874 B.n137 256.663
R641 B.n874 B.n136 256.663
R642 B.n874 B.n135 256.663
R643 B.n874 B.n134 256.663
R644 B.n874 B.n133 256.663
R645 B.n874 B.n132 256.663
R646 B.n874 B.n131 256.663
R647 B.n874 B.n130 256.663
R648 B.n874 B.n129 256.663
R649 B.n874 B.n128 256.663
R650 B.n874 B.n127 256.663
R651 B.n874 B.n126 256.663
R652 B.n874 B.n125 256.663
R653 B.n874 B.n124 256.663
R654 B.n874 B.n123 256.663
R655 B.n874 B.n122 256.663
R656 B.n874 B.n121 256.663
R657 B.n874 B.n120 256.663
R658 B.n874 B.n119 256.663
R659 B.n874 B.n118 256.663
R660 B.n874 B.n117 256.663
R661 B.n874 B.n116 256.663
R662 B.n874 B.n115 256.663
R663 B.n874 B.n114 256.663
R664 B.n874 B.n113 256.663
R665 B.n874 B.n112 256.663
R666 B.n874 B.n111 256.663
R667 B.n874 B.n110 256.663
R668 B.n874 B.n109 256.663
R669 B.n874 B.n108 256.663
R670 B.n874 B.n107 256.663
R671 B.n874 B.n106 256.663
R672 B.n624 B.n623 256.663
R673 B.n624 B.n423 256.663
R674 B.n624 B.n424 256.663
R675 B.n624 B.n425 256.663
R676 B.n624 B.n426 256.663
R677 B.n624 B.n427 256.663
R678 B.n624 B.n428 256.663
R679 B.n624 B.n429 256.663
R680 B.n624 B.n430 256.663
R681 B.n624 B.n431 256.663
R682 B.n624 B.n432 256.663
R683 B.n624 B.n433 256.663
R684 B.n624 B.n434 256.663
R685 B.n624 B.n435 256.663
R686 B.n624 B.n436 256.663
R687 B.n624 B.n437 256.663
R688 B.n624 B.n438 256.663
R689 B.n624 B.n439 256.663
R690 B.n624 B.n440 256.663
R691 B.n624 B.n441 256.663
R692 B.n624 B.n442 256.663
R693 B.n624 B.n443 256.663
R694 B.n624 B.n444 256.663
R695 B.n624 B.n445 256.663
R696 B.n624 B.n446 256.663
R697 B.n624 B.n447 256.663
R698 B.n624 B.n448 256.663
R699 B.n624 B.n449 256.663
R700 B.n624 B.n450 256.663
R701 B.n624 B.n451 256.663
R702 B.n624 B.n452 256.663
R703 B.n624 B.n453 256.663
R704 B.n624 B.n454 256.663
R705 B.n624 B.n455 256.663
R706 B.n624 B.n456 256.663
R707 B.n624 B.n457 256.663
R708 B.n624 B.n458 256.663
R709 B.n624 B.n459 256.663
R710 B.n624 B.n460 256.663
R711 B.n992 B.n991 256.663
R712 B.n154 B.n153 163.367
R713 B.n158 B.n157 163.367
R714 B.n162 B.n161 163.367
R715 B.n166 B.n165 163.367
R716 B.n170 B.n169 163.367
R717 B.n174 B.n173 163.367
R718 B.n178 B.n177 163.367
R719 B.n182 B.n181 163.367
R720 B.n186 B.n185 163.367
R721 B.n190 B.n189 163.367
R722 B.n194 B.n193 163.367
R723 B.n198 B.n197 163.367
R724 B.n202 B.n201 163.367
R725 B.n206 B.n205 163.367
R726 B.n210 B.n209 163.367
R727 B.n214 B.n213 163.367
R728 B.n218 B.n217 163.367
R729 B.n223 B.n222 163.367
R730 B.n227 B.n226 163.367
R731 B.n231 B.n230 163.367
R732 B.n235 B.n234 163.367
R733 B.n239 B.n238 163.367
R734 B.n244 B.n243 163.367
R735 B.n248 B.n247 163.367
R736 B.n252 B.n251 163.367
R737 B.n256 B.n255 163.367
R738 B.n260 B.n259 163.367
R739 B.n264 B.n263 163.367
R740 B.n268 B.n267 163.367
R741 B.n272 B.n271 163.367
R742 B.n276 B.n275 163.367
R743 B.n280 B.n279 163.367
R744 B.n284 B.n283 163.367
R745 B.n288 B.n287 163.367
R746 B.n292 B.n291 163.367
R747 B.n296 B.n295 163.367
R748 B.n300 B.n299 163.367
R749 B.n304 B.n303 163.367
R750 B.n306 B.n145 163.367
R751 B.n629 B.n420 163.367
R752 B.n629 B.n414 163.367
R753 B.n637 B.n414 163.367
R754 B.n637 B.n412 163.367
R755 B.n641 B.n412 163.367
R756 B.n641 B.n406 163.367
R757 B.n649 B.n406 163.367
R758 B.n649 B.n404 163.367
R759 B.n653 B.n404 163.367
R760 B.n653 B.n398 163.367
R761 B.n661 B.n398 163.367
R762 B.n661 B.n396 163.367
R763 B.n665 B.n396 163.367
R764 B.n665 B.n390 163.367
R765 B.n673 B.n390 163.367
R766 B.n673 B.n388 163.367
R767 B.n677 B.n388 163.367
R768 B.n677 B.n382 163.367
R769 B.n685 B.n382 163.367
R770 B.n685 B.n380 163.367
R771 B.n689 B.n380 163.367
R772 B.n689 B.n374 163.367
R773 B.n697 B.n374 163.367
R774 B.n697 B.n372 163.367
R775 B.n701 B.n372 163.367
R776 B.n701 B.n366 163.367
R777 B.n709 B.n366 163.367
R778 B.n709 B.n364 163.367
R779 B.n713 B.n364 163.367
R780 B.n713 B.n358 163.367
R781 B.n721 B.n358 163.367
R782 B.n721 B.n356 163.367
R783 B.n725 B.n356 163.367
R784 B.n725 B.n350 163.367
R785 B.n733 B.n350 163.367
R786 B.n733 B.n348 163.367
R787 B.n737 B.n348 163.367
R788 B.n737 B.n342 163.367
R789 B.n745 B.n342 163.367
R790 B.n745 B.n340 163.367
R791 B.n749 B.n340 163.367
R792 B.n749 B.n334 163.367
R793 B.n757 B.n334 163.367
R794 B.n757 B.n332 163.367
R795 B.n761 B.n332 163.367
R796 B.n761 B.n326 163.367
R797 B.n769 B.n326 163.367
R798 B.n769 B.n324 163.367
R799 B.n773 B.n324 163.367
R800 B.n773 B.n318 163.367
R801 B.n781 B.n318 163.367
R802 B.n781 B.n316 163.367
R803 B.n786 B.n316 163.367
R804 B.n786 B.n310 163.367
R805 B.n794 B.n310 163.367
R806 B.n795 B.n794 163.367
R807 B.n795 B.n5 163.367
R808 B.n6 B.n5 163.367
R809 B.n7 B.n6 163.367
R810 B.n801 B.n7 163.367
R811 B.n802 B.n801 163.367
R812 B.n802 B.n13 163.367
R813 B.n14 B.n13 163.367
R814 B.n15 B.n14 163.367
R815 B.n807 B.n15 163.367
R816 B.n807 B.n20 163.367
R817 B.n21 B.n20 163.367
R818 B.n22 B.n21 163.367
R819 B.n812 B.n22 163.367
R820 B.n812 B.n27 163.367
R821 B.n28 B.n27 163.367
R822 B.n29 B.n28 163.367
R823 B.n817 B.n29 163.367
R824 B.n817 B.n34 163.367
R825 B.n35 B.n34 163.367
R826 B.n36 B.n35 163.367
R827 B.n822 B.n36 163.367
R828 B.n822 B.n41 163.367
R829 B.n42 B.n41 163.367
R830 B.n43 B.n42 163.367
R831 B.n827 B.n43 163.367
R832 B.n827 B.n48 163.367
R833 B.n49 B.n48 163.367
R834 B.n50 B.n49 163.367
R835 B.n832 B.n50 163.367
R836 B.n832 B.n55 163.367
R837 B.n56 B.n55 163.367
R838 B.n57 B.n56 163.367
R839 B.n837 B.n57 163.367
R840 B.n837 B.n62 163.367
R841 B.n63 B.n62 163.367
R842 B.n64 B.n63 163.367
R843 B.n842 B.n64 163.367
R844 B.n842 B.n69 163.367
R845 B.n70 B.n69 163.367
R846 B.n71 B.n70 163.367
R847 B.n847 B.n71 163.367
R848 B.n847 B.n76 163.367
R849 B.n77 B.n76 163.367
R850 B.n78 B.n77 163.367
R851 B.n852 B.n78 163.367
R852 B.n852 B.n83 163.367
R853 B.n84 B.n83 163.367
R854 B.n85 B.n84 163.367
R855 B.n857 B.n85 163.367
R856 B.n857 B.n90 163.367
R857 B.n91 B.n90 163.367
R858 B.n92 B.n91 163.367
R859 B.n862 B.n92 163.367
R860 B.n862 B.n97 163.367
R861 B.n98 B.n97 163.367
R862 B.n99 B.n98 163.367
R863 B.n867 B.n99 163.367
R864 B.n867 B.n104 163.367
R865 B.n105 B.n104 163.367
R866 B.n462 B.n461 163.367
R867 B.n617 B.n461 163.367
R868 B.n615 B.n614 163.367
R869 B.n611 B.n610 163.367
R870 B.n607 B.n606 163.367
R871 B.n603 B.n602 163.367
R872 B.n599 B.n598 163.367
R873 B.n595 B.n594 163.367
R874 B.n591 B.n590 163.367
R875 B.n587 B.n586 163.367
R876 B.n583 B.n582 163.367
R877 B.n579 B.n578 163.367
R878 B.n575 B.n574 163.367
R879 B.n571 B.n570 163.367
R880 B.n567 B.n566 163.367
R881 B.n563 B.n562 163.367
R882 B.n559 B.n558 163.367
R883 B.n555 B.n554 163.367
R884 B.n551 B.n550 163.367
R885 B.n547 B.n546 163.367
R886 B.n543 B.n542 163.367
R887 B.n539 B.n538 163.367
R888 B.n535 B.n534 163.367
R889 B.n531 B.n530 163.367
R890 B.n527 B.n526 163.367
R891 B.n523 B.n522 163.367
R892 B.n519 B.n518 163.367
R893 B.n515 B.n514 163.367
R894 B.n511 B.n510 163.367
R895 B.n507 B.n506 163.367
R896 B.n503 B.n502 163.367
R897 B.n499 B.n498 163.367
R898 B.n495 B.n494 163.367
R899 B.n491 B.n490 163.367
R900 B.n487 B.n486 163.367
R901 B.n483 B.n482 163.367
R902 B.n479 B.n478 163.367
R903 B.n475 B.n474 163.367
R904 B.n471 B.n470 163.367
R905 B.n625 B.n422 163.367
R906 B.n631 B.n418 163.367
R907 B.n631 B.n416 163.367
R908 B.n635 B.n416 163.367
R909 B.n635 B.n410 163.367
R910 B.n643 B.n410 163.367
R911 B.n643 B.n408 163.367
R912 B.n647 B.n408 163.367
R913 B.n647 B.n402 163.367
R914 B.n655 B.n402 163.367
R915 B.n655 B.n400 163.367
R916 B.n659 B.n400 163.367
R917 B.n659 B.n394 163.367
R918 B.n667 B.n394 163.367
R919 B.n667 B.n392 163.367
R920 B.n671 B.n392 163.367
R921 B.n671 B.n386 163.367
R922 B.n679 B.n386 163.367
R923 B.n679 B.n384 163.367
R924 B.n683 B.n384 163.367
R925 B.n683 B.n378 163.367
R926 B.n691 B.n378 163.367
R927 B.n691 B.n376 163.367
R928 B.n695 B.n376 163.367
R929 B.n695 B.n370 163.367
R930 B.n703 B.n370 163.367
R931 B.n703 B.n368 163.367
R932 B.n707 B.n368 163.367
R933 B.n707 B.n362 163.367
R934 B.n715 B.n362 163.367
R935 B.n715 B.n360 163.367
R936 B.n719 B.n360 163.367
R937 B.n719 B.n354 163.367
R938 B.n727 B.n354 163.367
R939 B.n727 B.n352 163.367
R940 B.n731 B.n352 163.367
R941 B.n731 B.n346 163.367
R942 B.n739 B.n346 163.367
R943 B.n739 B.n344 163.367
R944 B.n743 B.n344 163.367
R945 B.n743 B.n338 163.367
R946 B.n751 B.n338 163.367
R947 B.n751 B.n336 163.367
R948 B.n755 B.n336 163.367
R949 B.n755 B.n330 163.367
R950 B.n763 B.n330 163.367
R951 B.n763 B.n328 163.367
R952 B.n767 B.n328 163.367
R953 B.n767 B.n322 163.367
R954 B.n775 B.n322 163.367
R955 B.n775 B.n320 163.367
R956 B.n779 B.n320 163.367
R957 B.n779 B.n314 163.367
R958 B.n788 B.n314 163.367
R959 B.n788 B.n312 163.367
R960 B.n792 B.n312 163.367
R961 B.n792 B.n3 163.367
R962 B.n990 B.n3 163.367
R963 B.n986 B.n2 163.367
R964 B.n986 B.n985 163.367
R965 B.n985 B.n9 163.367
R966 B.n981 B.n9 163.367
R967 B.n981 B.n11 163.367
R968 B.n977 B.n11 163.367
R969 B.n977 B.n17 163.367
R970 B.n973 B.n17 163.367
R971 B.n973 B.n19 163.367
R972 B.n969 B.n19 163.367
R973 B.n969 B.n24 163.367
R974 B.n965 B.n24 163.367
R975 B.n965 B.n26 163.367
R976 B.n961 B.n26 163.367
R977 B.n961 B.n31 163.367
R978 B.n957 B.n31 163.367
R979 B.n957 B.n33 163.367
R980 B.n953 B.n33 163.367
R981 B.n953 B.n38 163.367
R982 B.n949 B.n38 163.367
R983 B.n949 B.n40 163.367
R984 B.n945 B.n40 163.367
R985 B.n945 B.n45 163.367
R986 B.n941 B.n45 163.367
R987 B.n941 B.n47 163.367
R988 B.n937 B.n47 163.367
R989 B.n937 B.n52 163.367
R990 B.n933 B.n52 163.367
R991 B.n933 B.n54 163.367
R992 B.n929 B.n54 163.367
R993 B.n929 B.n59 163.367
R994 B.n925 B.n59 163.367
R995 B.n925 B.n61 163.367
R996 B.n921 B.n61 163.367
R997 B.n921 B.n66 163.367
R998 B.n917 B.n66 163.367
R999 B.n917 B.n68 163.367
R1000 B.n913 B.n68 163.367
R1001 B.n913 B.n73 163.367
R1002 B.n909 B.n73 163.367
R1003 B.n909 B.n75 163.367
R1004 B.n905 B.n75 163.367
R1005 B.n905 B.n80 163.367
R1006 B.n901 B.n80 163.367
R1007 B.n901 B.n82 163.367
R1008 B.n897 B.n82 163.367
R1009 B.n897 B.n87 163.367
R1010 B.n893 B.n87 163.367
R1011 B.n893 B.n89 163.367
R1012 B.n889 B.n89 163.367
R1013 B.n889 B.n94 163.367
R1014 B.n885 B.n94 163.367
R1015 B.n885 B.n96 163.367
R1016 B.n881 B.n96 163.367
R1017 B.n881 B.n101 163.367
R1018 B.n877 B.n101 163.367
R1019 B.n877 B.n103 163.367
R1020 B.n146 B.t10 155.042
R1021 B.n466 B.t15 155.042
R1022 B.n148 B.t7 155.03
R1023 B.n463 B.t18 155.03
R1024 B.n624 B.n419 91.2111
R1025 B.n875 B.n874 91.2111
R1026 B.n149 B.n148 81.455
R1027 B.n147 B.n146 81.455
R1028 B.n467 B.n466 81.455
R1029 B.n464 B.n463 81.455
R1030 B.n147 B.t11 73.5872
R1031 B.n467 B.t14 73.5872
R1032 B.n149 B.t8 73.5754
R1033 B.n464 B.t17 73.5754
R1034 B.n150 B.n106 71.676
R1035 B.n154 B.n107 71.676
R1036 B.n158 B.n108 71.676
R1037 B.n162 B.n109 71.676
R1038 B.n166 B.n110 71.676
R1039 B.n170 B.n111 71.676
R1040 B.n174 B.n112 71.676
R1041 B.n178 B.n113 71.676
R1042 B.n182 B.n114 71.676
R1043 B.n186 B.n115 71.676
R1044 B.n190 B.n116 71.676
R1045 B.n194 B.n117 71.676
R1046 B.n198 B.n118 71.676
R1047 B.n202 B.n119 71.676
R1048 B.n206 B.n120 71.676
R1049 B.n210 B.n121 71.676
R1050 B.n214 B.n122 71.676
R1051 B.n218 B.n123 71.676
R1052 B.n223 B.n124 71.676
R1053 B.n227 B.n125 71.676
R1054 B.n231 B.n126 71.676
R1055 B.n235 B.n127 71.676
R1056 B.n239 B.n128 71.676
R1057 B.n244 B.n129 71.676
R1058 B.n248 B.n130 71.676
R1059 B.n252 B.n131 71.676
R1060 B.n256 B.n132 71.676
R1061 B.n260 B.n133 71.676
R1062 B.n264 B.n134 71.676
R1063 B.n268 B.n135 71.676
R1064 B.n272 B.n136 71.676
R1065 B.n276 B.n137 71.676
R1066 B.n280 B.n138 71.676
R1067 B.n284 B.n139 71.676
R1068 B.n288 B.n140 71.676
R1069 B.n292 B.n141 71.676
R1070 B.n296 B.n142 71.676
R1071 B.n300 B.n143 71.676
R1072 B.n304 B.n144 71.676
R1073 B.n873 B.n145 71.676
R1074 B.n873 B.n872 71.676
R1075 B.n306 B.n144 71.676
R1076 B.n303 B.n143 71.676
R1077 B.n299 B.n142 71.676
R1078 B.n295 B.n141 71.676
R1079 B.n291 B.n140 71.676
R1080 B.n287 B.n139 71.676
R1081 B.n283 B.n138 71.676
R1082 B.n279 B.n137 71.676
R1083 B.n275 B.n136 71.676
R1084 B.n271 B.n135 71.676
R1085 B.n267 B.n134 71.676
R1086 B.n263 B.n133 71.676
R1087 B.n259 B.n132 71.676
R1088 B.n255 B.n131 71.676
R1089 B.n251 B.n130 71.676
R1090 B.n247 B.n129 71.676
R1091 B.n243 B.n128 71.676
R1092 B.n238 B.n127 71.676
R1093 B.n234 B.n126 71.676
R1094 B.n230 B.n125 71.676
R1095 B.n226 B.n124 71.676
R1096 B.n222 B.n123 71.676
R1097 B.n217 B.n122 71.676
R1098 B.n213 B.n121 71.676
R1099 B.n209 B.n120 71.676
R1100 B.n205 B.n119 71.676
R1101 B.n201 B.n118 71.676
R1102 B.n197 B.n117 71.676
R1103 B.n193 B.n116 71.676
R1104 B.n189 B.n115 71.676
R1105 B.n185 B.n114 71.676
R1106 B.n181 B.n113 71.676
R1107 B.n177 B.n112 71.676
R1108 B.n173 B.n111 71.676
R1109 B.n169 B.n110 71.676
R1110 B.n165 B.n109 71.676
R1111 B.n161 B.n108 71.676
R1112 B.n157 B.n107 71.676
R1113 B.n153 B.n106 71.676
R1114 B.n623 B.n622 71.676
R1115 B.n617 B.n423 71.676
R1116 B.n614 B.n424 71.676
R1117 B.n610 B.n425 71.676
R1118 B.n606 B.n426 71.676
R1119 B.n602 B.n427 71.676
R1120 B.n598 B.n428 71.676
R1121 B.n594 B.n429 71.676
R1122 B.n590 B.n430 71.676
R1123 B.n586 B.n431 71.676
R1124 B.n582 B.n432 71.676
R1125 B.n578 B.n433 71.676
R1126 B.n574 B.n434 71.676
R1127 B.n570 B.n435 71.676
R1128 B.n566 B.n436 71.676
R1129 B.n562 B.n437 71.676
R1130 B.n558 B.n438 71.676
R1131 B.n554 B.n439 71.676
R1132 B.n550 B.n440 71.676
R1133 B.n546 B.n441 71.676
R1134 B.n542 B.n442 71.676
R1135 B.n538 B.n443 71.676
R1136 B.n534 B.n444 71.676
R1137 B.n530 B.n445 71.676
R1138 B.n526 B.n446 71.676
R1139 B.n522 B.n447 71.676
R1140 B.n518 B.n448 71.676
R1141 B.n514 B.n449 71.676
R1142 B.n510 B.n450 71.676
R1143 B.n506 B.n451 71.676
R1144 B.n502 B.n452 71.676
R1145 B.n498 B.n453 71.676
R1146 B.n494 B.n454 71.676
R1147 B.n490 B.n455 71.676
R1148 B.n486 B.n456 71.676
R1149 B.n482 B.n457 71.676
R1150 B.n478 B.n458 71.676
R1151 B.n474 B.n459 71.676
R1152 B.n470 B.n460 71.676
R1153 B.n623 B.n462 71.676
R1154 B.n615 B.n423 71.676
R1155 B.n611 B.n424 71.676
R1156 B.n607 B.n425 71.676
R1157 B.n603 B.n426 71.676
R1158 B.n599 B.n427 71.676
R1159 B.n595 B.n428 71.676
R1160 B.n591 B.n429 71.676
R1161 B.n587 B.n430 71.676
R1162 B.n583 B.n431 71.676
R1163 B.n579 B.n432 71.676
R1164 B.n575 B.n433 71.676
R1165 B.n571 B.n434 71.676
R1166 B.n567 B.n435 71.676
R1167 B.n563 B.n436 71.676
R1168 B.n559 B.n437 71.676
R1169 B.n555 B.n438 71.676
R1170 B.n551 B.n439 71.676
R1171 B.n547 B.n440 71.676
R1172 B.n543 B.n441 71.676
R1173 B.n539 B.n442 71.676
R1174 B.n535 B.n443 71.676
R1175 B.n531 B.n444 71.676
R1176 B.n527 B.n445 71.676
R1177 B.n523 B.n446 71.676
R1178 B.n519 B.n447 71.676
R1179 B.n515 B.n448 71.676
R1180 B.n511 B.n449 71.676
R1181 B.n507 B.n450 71.676
R1182 B.n503 B.n451 71.676
R1183 B.n499 B.n452 71.676
R1184 B.n495 B.n453 71.676
R1185 B.n491 B.n454 71.676
R1186 B.n487 B.n455 71.676
R1187 B.n483 B.n456 71.676
R1188 B.n479 B.n457 71.676
R1189 B.n475 B.n458 71.676
R1190 B.n471 B.n459 71.676
R1191 B.n460 B.n422 71.676
R1192 B.n991 B.n990 71.676
R1193 B.n991 B.n2 71.676
R1194 B.n220 B.n149 59.5399
R1195 B.n241 B.n147 59.5399
R1196 B.n468 B.n467 59.5399
R1197 B.n465 B.n464 59.5399
R1198 B.n630 B.n419 49.6191
R1199 B.n630 B.n415 49.6191
R1200 B.n636 B.n415 49.6191
R1201 B.n636 B.n411 49.6191
R1202 B.n642 B.n411 49.6191
R1203 B.n642 B.n407 49.6191
R1204 B.n648 B.n407 49.6191
R1205 B.n648 B.n403 49.6191
R1206 B.n654 B.n403 49.6191
R1207 B.n660 B.n399 49.6191
R1208 B.n660 B.n395 49.6191
R1209 B.n666 B.n395 49.6191
R1210 B.n666 B.n391 49.6191
R1211 B.n672 B.n391 49.6191
R1212 B.n672 B.n387 49.6191
R1213 B.n678 B.n387 49.6191
R1214 B.n678 B.n383 49.6191
R1215 B.n684 B.n383 49.6191
R1216 B.n684 B.n379 49.6191
R1217 B.n690 B.n379 49.6191
R1218 B.n690 B.n375 49.6191
R1219 B.n696 B.n375 49.6191
R1220 B.n696 B.n371 49.6191
R1221 B.n702 B.n371 49.6191
R1222 B.n708 B.n367 49.6191
R1223 B.n708 B.n363 49.6191
R1224 B.n714 B.n363 49.6191
R1225 B.n714 B.n359 49.6191
R1226 B.n720 B.n359 49.6191
R1227 B.n720 B.n355 49.6191
R1228 B.n726 B.n355 49.6191
R1229 B.n726 B.n351 49.6191
R1230 B.n732 B.n351 49.6191
R1231 B.n732 B.n347 49.6191
R1232 B.n738 B.n347 49.6191
R1233 B.n744 B.n343 49.6191
R1234 B.n744 B.n339 49.6191
R1235 B.n750 B.n339 49.6191
R1236 B.n750 B.n335 49.6191
R1237 B.n756 B.n335 49.6191
R1238 B.n756 B.n331 49.6191
R1239 B.n762 B.n331 49.6191
R1240 B.n762 B.n327 49.6191
R1241 B.n768 B.n327 49.6191
R1242 B.n768 B.n323 49.6191
R1243 B.n774 B.n323 49.6191
R1244 B.n780 B.n319 49.6191
R1245 B.n780 B.n315 49.6191
R1246 B.n787 B.n315 49.6191
R1247 B.n787 B.n311 49.6191
R1248 B.n793 B.n311 49.6191
R1249 B.n793 B.n4 49.6191
R1250 B.n989 B.n4 49.6191
R1251 B.n989 B.n988 49.6191
R1252 B.n988 B.n987 49.6191
R1253 B.n987 B.n8 49.6191
R1254 B.n12 B.n8 49.6191
R1255 B.n980 B.n12 49.6191
R1256 B.n980 B.n979 49.6191
R1257 B.n979 B.n978 49.6191
R1258 B.n978 B.n16 49.6191
R1259 B.n972 B.n971 49.6191
R1260 B.n971 B.n970 49.6191
R1261 B.n970 B.n23 49.6191
R1262 B.n964 B.n23 49.6191
R1263 B.n964 B.n963 49.6191
R1264 B.n963 B.n962 49.6191
R1265 B.n962 B.n30 49.6191
R1266 B.n956 B.n30 49.6191
R1267 B.n956 B.n955 49.6191
R1268 B.n955 B.n954 49.6191
R1269 B.n954 B.n37 49.6191
R1270 B.n948 B.n947 49.6191
R1271 B.n947 B.n946 49.6191
R1272 B.n946 B.n44 49.6191
R1273 B.n940 B.n44 49.6191
R1274 B.n940 B.n939 49.6191
R1275 B.n939 B.n938 49.6191
R1276 B.n938 B.n51 49.6191
R1277 B.n932 B.n51 49.6191
R1278 B.n932 B.n931 49.6191
R1279 B.n931 B.n930 49.6191
R1280 B.n930 B.n58 49.6191
R1281 B.n924 B.n923 49.6191
R1282 B.n923 B.n922 49.6191
R1283 B.n922 B.n65 49.6191
R1284 B.n916 B.n65 49.6191
R1285 B.n916 B.n915 49.6191
R1286 B.n915 B.n914 49.6191
R1287 B.n914 B.n72 49.6191
R1288 B.n908 B.n72 49.6191
R1289 B.n908 B.n907 49.6191
R1290 B.n907 B.n906 49.6191
R1291 B.n906 B.n79 49.6191
R1292 B.n900 B.n79 49.6191
R1293 B.n900 B.n899 49.6191
R1294 B.n899 B.n898 49.6191
R1295 B.n898 B.n86 49.6191
R1296 B.n892 B.n891 49.6191
R1297 B.n891 B.n890 49.6191
R1298 B.n890 B.n93 49.6191
R1299 B.n884 B.n93 49.6191
R1300 B.n884 B.n883 49.6191
R1301 B.n883 B.n882 49.6191
R1302 B.n882 B.n100 49.6191
R1303 B.n876 B.n100 49.6191
R1304 B.n876 B.n875 49.6191
R1305 B.t0 B.n367 48.8894
R1306 B.t2 B.n58 48.8894
R1307 B.n774 B.t19 35.7551
R1308 B.n972 B.t3 35.7551
R1309 B.n621 B.n417 32.0005
R1310 B.n627 B.n626 32.0005
R1311 B.n871 B.n870 32.0005
R1312 B.n151 B.n102 32.0005
R1313 B.t4 B.n343 31.377
R1314 B.t1 B.n37 31.377
R1315 B.t13 B.n399 26.9988
R1316 B.t6 B.n86 26.9988
R1317 B.n654 B.t13 22.6207
R1318 B.n892 B.t6 22.6207
R1319 B.n738 B.t4 18.2426
R1320 B.n948 B.t1 18.2426
R1321 B B.n992 18.0485
R1322 B.t19 B.n319 13.8645
R1323 B.t3 B.n16 13.8645
R1324 B.n632 B.n417 10.6151
R1325 B.n633 B.n632 10.6151
R1326 B.n634 B.n633 10.6151
R1327 B.n634 B.n409 10.6151
R1328 B.n644 B.n409 10.6151
R1329 B.n645 B.n644 10.6151
R1330 B.n646 B.n645 10.6151
R1331 B.n646 B.n401 10.6151
R1332 B.n656 B.n401 10.6151
R1333 B.n657 B.n656 10.6151
R1334 B.n658 B.n657 10.6151
R1335 B.n658 B.n393 10.6151
R1336 B.n668 B.n393 10.6151
R1337 B.n669 B.n668 10.6151
R1338 B.n670 B.n669 10.6151
R1339 B.n670 B.n385 10.6151
R1340 B.n680 B.n385 10.6151
R1341 B.n681 B.n680 10.6151
R1342 B.n682 B.n681 10.6151
R1343 B.n682 B.n377 10.6151
R1344 B.n692 B.n377 10.6151
R1345 B.n693 B.n692 10.6151
R1346 B.n694 B.n693 10.6151
R1347 B.n694 B.n369 10.6151
R1348 B.n704 B.n369 10.6151
R1349 B.n705 B.n704 10.6151
R1350 B.n706 B.n705 10.6151
R1351 B.n706 B.n361 10.6151
R1352 B.n716 B.n361 10.6151
R1353 B.n717 B.n716 10.6151
R1354 B.n718 B.n717 10.6151
R1355 B.n718 B.n353 10.6151
R1356 B.n728 B.n353 10.6151
R1357 B.n729 B.n728 10.6151
R1358 B.n730 B.n729 10.6151
R1359 B.n730 B.n345 10.6151
R1360 B.n740 B.n345 10.6151
R1361 B.n741 B.n740 10.6151
R1362 B.n742 B.n741 10.6151
R1363 B.n742 B.n337 10.6151
R1364 B.n752 B.n337 10.6151
R1365 B.n753 B.n752 10.6151
R1366 B.n754 B.n753 10.6151
R1367 B.n754 B.n329 10.6151
R1368 B.n764 B.n329 10.6151
R1369 B.n765 B.n764 10.6151
R1370 B.n766 B.n765 10.6151
R1371 B.n766 B.n321 10.6151
R1372 B.n776 B.n321 10.6151
R1373 B.n777 B.n776 10.6151
R1374 B.n778 B.n777 10.6151
R1375 B.n778 B.n313 10.6151
R1376 B.n789 B.n313 10.6151
R1377 B.n790 B.n789 10.6151
R1378 B.n791 B.n790 10.6151
R1379 B.n791 B.n0 10.6151
R1380 B.n621 B.n620 10.6151
R1381 B.n620 B.n619 10.6151
R1382 B.n619 B.n618 10.6151
R1383 B.n618 B.n616 10.6151
R1384 B.n616 B.n613 10.6151
R1385 B.n613 B.n612 10.6151
R1386 B.n612 B.n609 10.6151
R1387 B.n609 B.n608 10.6151
R1388 B.n608 B.n605 10.6151
R1389 B.n605 B.n604 10.6151
R1390 B.n604 B.n601 10.6151
R1391 B.n601 B.n600 10.6151
R1392 B.n600 B.n597 10.6151
R1393 B.n597 B.n596 10.6151
R1394 B.n596 B.n593 10.6151
R1395 B.n593 B.n592 10.6151
R1396 B.n592 B.n589 10.6151
R1397 B.n589 B.n588 10.6151
R1398 B.n588 B.n585 10.6151
R1399 B.n585 B.n584 10.6151
R1400 B.n584 B.n581 10.6151
R1401 B.n581 B.n580 10.6151
R1402 B.n580 B.n577 10.6151
R1403 B.n577 B.n576 10.6151
R1404 B.n576 B.n573 10.6151
R1405 B.n573 B.n572 10.6151
R1406 B.n572 B.n569 10.6151
R1407 B.n569 B.n568 10.6151
R1408 B.n568 B.n565 10.6151
R1409 B.n565 B.n564 10.6151
R1410 B.n564 B.n561 10.6151
R1411 B.n561 B.n560 10.6151
R1412 B.n560 B.n557 10.6151
R1413 B.n557 B.n556 10.6151
R1414 B.n553 B.n552 10.6151
R1415 B.n552 B.n549 10.6151
R1416 B.n549 B.n548 10.6151
R1417 B.n548 B.n545 10.6151
R1418 B.n545 B.n544 10.6151
R1419 B.n544 B.n541 10.6151
R1420 B.n541 B.n540 10.6151
R1421 B.n540 B.n537 10.6151
R1422 B.n537 B.n536 10.6151
R1423 B.n533 B.n532 10.6151
R1424 B.n532 B.n529 10.6151
R1425 B.n529 B.n528 10.6151
R1426 B.n528 B.n525 10.6151
R1427 B.n525 B.n524 10.6151
R1428 B.n524 B.n521 10.6151
R1429 B.n521 B.n520 10.6151
R1430 B.n520 B.n517 10.6151
R1431 B.n517 B.n516 10.6151
R1432 B.n516 B.n513 10.6151
R1433 B.n513 B.n512 10.6151
R1434 B.n512 B.n509 10.6151
R1435 B.n509 B.n508 10.6151
R1436 B.n508 B.n505 10.6151
R1437 B.n505 B.n504 10.6151
R1438 B.n504 B.n501 10.6151
R1439 B.n501 B.n500 10.6151
R1440 B.n500 B.n497 10.6151
R1441 B.n497 B.n496 10.6151
R1442 B.n496 B.n493 10.6151
R1443 B.n493 B.n492 10.6151
R1444 B.n492 B.n489 10.6151
R1445 B.n489 B.n488 10.6151
R1446 B.n488 B.n485 10.6151
R1447 B.n485 B.n484 10.6151
R1448 B.n484 B.n481 10.6151
R1449 B.n481 B.n480 10.6151
R1450 B.n480 B.n477 10.6151
R1451 B.n477 B.n476 10.6151
R1452 B.n476 B.n473 10.6151
R1453 B.n473 B.n472 10.6151
R1454 B.n472 B.n469 10.6151
R1455 B.n469 B.n421 10.6151
R1456 B.n626 B.n421 10.6151
R1457 B.n628 B.n627 10.6151
R1458 B.n628 B.n413 10.6151
R1459 B.n638 B.n413 10.6151
R1460 B.n639 B.n638 10.6151
R1461 B.n640 B.n639 10.6151
R1462 B.n640 B.n405 10.6151
R1463 B.n650 B.n405 10.6151
R1464 B.n651 B.n650 10.6151
R1465 B.n652 B.n651 10.6151
R1466 B.n652 B.n397 10.6151
R1467 B.n662 B.n397 10.6151
R1468 B.n663 B.n662 10.6151
R1469 B.n664 B.n663 10.6151
R1470 B.n664 B.n389 10.6151
R1471 B.n674 B.n389 10.6151
R1472 B.n675 B.n674 10.6151
R1473 B.n676 B.n675 10.6151
R1474 B.n676 B.n381 10.6151
R1475 B.n686 B.n381 10.6151
R1476 B.n687 B.n686 10.6151
R1477 B.n688 B.n687 10.6151
R1478 B.n688 B.n373 10.6151
R1479 B.n698 B.n373 10.6151
R1480 B.n699 B.n698 10.6151
R1481 B.n700 B.n699 10.6151
R1482 B.n700 B.n365 10.6151
R1483 B.n710 B.n365 10.6151
R1484 B.n711 B.n710 10.6151
R1485 B.n712 B.n711 10.6151
R1486 B.n712 B.n357 10.6151
R1487 B.n722 B.n357 10.6151
R1488 B.n723 B.n722 10.6151
R1489 B.n724 B.n723 10.6151
R1490 B.n724 B.n349 10.6151
R1491 B.n734 B.n349 10.6151
R1492 B.n735 B.n734 10.6151
R1493 B.n736 B.n735 10.6151
R1494 B.n736 B.n341 10.6151
R1495 B.n746 B.n341 10.6151
R1496 B.n747 B.n746 10.6151
R1497 B.n748 B.n747 10.6151
R1498 B.n748 B.n333 10.6151
R1499 B.n758 B.n333 10.6151
R1500 B.n759 B.n758 10.6151
R1501 B.n760 B.n759 10.6151
R1502 B.n760 B.n325 10.6151
R1503 B.n770 B.n325 10.6151
R1504 B.n771 B.n770 10.6151
R1505 B.n772 B.n771 10.6151
R1506 B.n772 B.n317 10.6151
R1507 B.n782 B.n317 10.6151
R1508 B.n783 B.n782 10.6151
R1509 B.n785 B.n783 10.6151
R1510 B.n785 B.n784 10.6151
R1511 B.n784 B.n309 10.6151
R1512 B.n796 B.n309 10.6151
R1513 B.n797 B.n796 10.6151
R1514 B.n798 B.n797 10.6151
R1515 B.n799 B.n798 10.6151
R1516 B.n800 B.n799 10.6151
R1517 B.n803 B.n800 10.6151
R1518 B.n804 B.n803 10.6151
R1519 B.n805 B.n804 10.6151
R1520 B.n806 B.n805 10.6151
R1521 B.n808 B.n806 10.6151
R1522 B.n809 B.n808 10.6151
R1523 B.n810 B.n809 10.6151
R1524 B.n811 B.n810 10.6151
R1525 B.n813 B.n811 10.6151
R1526 B.n814 B.n813 10.6151
R1527 B.n815 B.n814 10.6151
R1528 B.n816 B.n815 10.6151
R1529 B.n818 B.n816 10.6151
R1530 B.n819 B.n818 10.6151
R1531 B.n820 B.n819 10.6151
R1532 B.n821 B.n820 10.6151
R1533 B.n823 B.n821 10.6151
R1534 B.n824 B.n823 10.6151
R1535 B.n825 B.n824 10.6151
R1536 B.n826 B.n825 10.6151
R1537 B.n828 B.n826 10.6151
R1538 B.n829 B.n828 10.6151
R1539 B.n830 B.n829 10.6151
R1540 B.n831 B.n830 10.6151
R1541 B.n833 B.n831 10.6151
R1542 B.n834 B.n833 10.6151
R1543 B.n835 B.n834 10.6151
R1544 B.n836 B.n835 10.6151
R1545 B.n838 B.n836 10.6151
R1546 B.n839 B.n838 10.6151
R1547 B.n840 B.n839 10.6151
R1548 B.n841 B.n840 10.6151
R1549 B.n843 B.n841 10.6151
R1550 B.n844 B.n843 10.6151
R1551 B.n845 B.n844 10.6151
R1552 B.n846 B.n845 10.6151
R1553 B.n848 B.n846 10.6151
R1554 B.n849 B.n848 10.6151
R1555 B.n850 B.n849 10.6151
R1556 B.n851 B.n850 10.6151
R1557 B.n853 B.n851 10.6151
R1558 B.n854 B.n853 10.6151
R1559 B.n855 B.n854 10.6151
R1560 B.n856 B.n855 10.6151
R1561 B.n858 B.n856 10.6151
R1562 B.n859 B.n858 10.6151
R1563 B.n860 B.n859 10.6151
R1564 B.n861 B.n860 10.6151
R1565 B.n863 B.n861 10.6151
R1566 B.n864 B.n863 10.6151
R1567 B.n865 B.n864 10.6151
R1568 B.n866 B.n865 10.6151
R1569 B.n868 B.n866 10.6151
R1570 B.n869 B.n868 10.6151
R1571 B.n870 B.n869 10.6151
R1572 B.n984 B.n1 10.6151
R1573 B.n984 B.n983 10.6151
R1574 B.n983 B.n982 10.6151
R1575 B.n982 B.n10 10.6151
R1576 B.n976 B.n10 10.6151
R1577 B.n976 B.n975 10.6151
R1578 B.n975 B.n974 10.6151
R1579 B.n974 B.n18 10.6151
R1580 B.n968 B.n18 10.6151
R1581 B.n968 B.n967 10.6151
R1582 B.n967 B.n966 10.6151
R1583 B.n966 B.n25 10.6151
R1584 B.n960 B.n25 10.6151
R1585 B.n960 B.n959 10.6151
R1586 B.n959 B.n958 10.6151
R1587 B.n958 B.n32 10.6151
R1588 B.n952 B.n32 10.6151
R1589 B.n952 B.n951 10.6151
R1590 B.n951 B.n950 10.6151
R1591 B.n950 B.n39 10.6151
R1592 B.n944 B.n39 10.6151
R1593 B.n944 B.n943 10.6151
R1594 B.n943 B.n942 10.6151
R1595 B.n942 B.n46 10.6151
R1596 B.n936 B.n46 10.6151
R1597 B.n936 B.n935 10.6151
R1598 B.n935 B.n934 10.6151
R1599 B.n934 B.n53 10.6151
R1600 B.n928 B.n53 10.6151
R1601 B.n928 B.n927 10.6151
R1602 B.n927 B.n926 10.6151
R1603 B.n926 B.n60 10.6151
R1604 B.n920 B.n60 10.6151
R1605 B.n920 B.n919 10.6151
R1606 B.n919 B.n918 10.6151
R1607 B.n918 B.n67 10.6151
R1608 B.n912 B.n67 10.6151
R1609 B.n912 B.n911 10.6151
R1610 B.n911 B.n910 10.6151
R1611 B.n910 B.n74 10.6151
R1612 B.n904 B.n74 10.6151
R1613 B.n904 B.n903 10.6151
R1614 B.n903 B.n902 10.6151
R1615 B.n902 B.n81 10.6151
R1616 B.n896 B.n81 10.6151
R1617 B.n896 B.n895 10.6151
R1618 B.n895 B.n894 10.6151
R1619 B.n894 B.n88 10.6151
R1620 B.n888 B.n88 10.6151
R1621 B.n888 B.n887 10.6151
R1622 B.n887 B.n886 10.6151
R1623 B.n886 B.n95 10.6151
R1624 B.n880 B.n95 10.6151
R1625 B.n880 B.n879 10.6151
R1626 B.n879 B.n878 10.6151
R1627 B.n878 B.n102 10.6151
R1628 B.n152 B.n151 10.6151
R1629 B.n155 B.n152 10.6151
R1630 B.n156 B.n155 10.6151
R1631 B.n159 B.n156 10.6151
R1632 B.n160 B.n159 10.6151
R1633 B.n163 B.n160 10.6151
R1634 B.n164 B.n163 10.6151
R1635 B.n167 B.n164 10.6151
R1636 B.n168 B.n167 10.6151
R1637 B.n171 B.n168 10.6151
R1638 B.n172 B.n171 10.6151
R1639 B.n175 B.n172 10.6151
R1640 B.n176 B.n175 10.6151
R1641 B.n179 B.n176 10.6151
R1642 B.n180 B.n179 10.6151
R1643 B.n183 B.n180 10.6151
R1644 B.n184 B.n183 10.6151
R1645 B.n187 B.n184 10.6151
R1646 B.n188 B.n187 10.6151
R1647 B.n191 B.n188 10.6151
R1648 B.n192 B.n191 10.6151
R1649 B.n195 B.n192 10.6151
R1650 B.n196 B.n195 10.6151
R1651 B.n199 B.n196 10.6151
R1652 B.n200 B.n199 10.6151
R1653 B.n203 B.n200 10.6151
R1654 B.n204 B.n203 10.6151
R1655 B.n207 B.n204 10.6151
R1656 B.n208 B.n207 10.6151
R1657 B.n211 B.n208 10.6151
R1658 B.n212 B.n211 10.6151
R1659 B.n215 B.n212 10.6151
R1660 B.n216 B.n215 10.6151
R1661 B.n219 B.n216 10.6151
R1662 B.n224 B.n221 10.6151
R1663 B.n225 B.n224 10.6151
R1664 B.n228 B.n225 10.6151
R1665 B.n229 B.n228 10.6151
R1666 B.n232 B.n229 10.6151
R1667 B.n233 B.n232 10.6151
R1668 B.n236 B.n233 10.6151
R1669 B.n237 B.n236 10.6151
R1670 B.n240 B.n237 10.6151
R1671 B.n245 B.n242 10.6151
R1672 B.n246 B.n245 10.6151
R1673 B.n249 B.n246 10.6151
R1674 B.n250 B.n249 10.6151
R1675 B.n253 B.n250 10.6151
R1676 B.n254 B.n253 10.6151
R1677 B.n257 B.n254 10.6151
R1678 B.n258 B.n257 10.6151
R1679 B.n261 B.n258 10.6151
R1680 B.n262 B.n261 10.6151
R1681 B.n265 B.n262 10.6151
R1682 B.n266 B.n265 10.6151
R1683 B.n269 B.n266 10.6151
R1684 B.n270 B.n269 10.6151
R1685 B.n273 B.n270 10.6151
R1686 B.n274 B.n273 10.6151
R1687 B.n277 B.n274 10.6151
R1688 B.n278 B.n277 10.6151
R1689 B.n281 B.n278 10.6151
R1690 B.n282 B.n281 10.6151
R1691 B.n285 B.n282 10.6151
R1692 B.n286 B.n285 10.6151
R1693 B.n289 B.n286 10.6151
R1694 B.n290 B.n289 10.6151
R1695 B.n293 B.n290 10.6151
R1696 B.n294 B.n293 10.6151
R1697 B.n297 B.n294 10.6151
R1698 B.n298 B.n297 10.6151
R1699 B.n301 B.n298 10.6151
R1700 B.n302 B.n301 10.6151
R1701 B.n305 B.n302 10.6151
R1702 B.n307 B.n305 10.6151
R1703 B.n308 B.n307 10.6151
R1704 B.n871 B.n308 10.6151
R1705 B.n556 B.n465 9.36635
R1706 B.n533 B.n468 9.36635
R1707 B.n220 B.n219 9.36635
R1708 B.n242 B.n241 9.36635
R1709 B.n992 B.n0 8.11757
R1710 B.n992 B.n1 8.11757
R1711 B.n553 B.n465 1.24928
R1712 B.n536 B.n468 1.24928
R1713 B.n221 B.n220 1.24928
R1714 B.n241 B.n240 1.24928
R1715 B.n702 B.t0 0.730185
R1716 B.n924 B.t2 0.730185
R1717 VP.n15 VP.n14 161.3
R1718 VP.n16 VP.n11 161.3
R1719 VP.n18 VP.n17 161.3
R1720 VP.n19 VP.n10 161.3
R1721 VP.n21 VP.n20 161.3
R1722 VP.n22 VP.n9 161.3
R1723 VP.n24 VP.n23 161.3
R1724 VP.n25 VP.n8 161.3
R1725 VP.n54 VP.n0 161.3
R1726 VP.n53 VP.n52 161.3
R1727 VP.n51 VP.n1 161.3
R1728 VP.n50 VP.n49 161.3
R1729 VP.n48 VP.n2 161.3
R1730 VP.n47 VP.n46 161.3
R1731 VP.n45 VP.n3 161.3
R1732 VP.n44 VP.n43 161.3
R1733 VP.n41 VP.n4 161.3
R1734 VP.n40 VP.n39 161.3
R1735 VP.n38 VP.n5 161.3
R1736 VP.n37 VP.n36 161.3
R1737 VP.n35 VP.n6 161.3
R1738 VP.n34 VP.n33 161.3
R1739 VP.n32 VP.n7 161.3
R1740 VP.n31 VP.n30 161.3
R1741 VP.n12 VP.t4 93.1314
R1742 VP.n13 VP.n12 62.7068
R1743 VP.n29 VP.t0 61.0289
R1744 VP.n42 VP.t5 61.0289
R1745 VP.n55 VP.t2 61.0289
R1746 VP.n26 VP.t3 61.0289
R1747 VP.n13 VP.t1 61.0289
R1748 VP.n29 VP.n28 60.0765
R1749 VP.n56 VP.n55 60.0765
R1750 VP.n27 VP.n26 60.0765
R1751 VP.n36 VP.n35 55.0167
R1752 VP.n49 VP.n48 55.0167
R1753 VP.n20 VP.n19 55.0167
R1754 VP.n28 VP.n27 52.2308
R1755 VP.n35 VP.n34 25.8045
R1756 VP.n49 VP.n1 25.8045
R1757 VP.n20 VP.n9 25.8045
R1758 VP.n30 VP.n7 24.3439
R1759 VP.n34 VP.n7 24.3439
R1760 VP.n36 VP.n5 24.3439
R1761 VP.n40 VP.n5 24.3439
R1762 VP.n41 VP.n40 24.3439
R1763 VP.n43 VP.n3 24.3439
R1764 VP.n47 VP.n3 24.3439
R1765 VP.n48 VP.n47 24.3439
R1766 VP.n53 VP.n1 24.3439
R1767 VP.n54 VP.n53 24.3439
R1768 VP.n24 VP.n9 24.3439
R1769 VP.n25 VP.n24 24.3439
R1770 VP.n14 VP.n11 24.3439
R1771 VP.n18 VP.n11 24.3439
R1772 VP.n19 VP.n18 24.3439
R1773 VP.n30 VP.n29 21.9096
R1774 VP.n55 VP.n54 21.9096
R1775 VP.n26 VP.n25 21.9096
R1776 VP.n42 VP.n41 12.1722
R1777 VP.n43 VP.n42 12.1722
R1778 VP.n14 VP.n13 12.1722
R1779 VP.n15 VP.n12 2.63302
R1780 VP.n27 VP.n8 0.417764
R1781 VP.n31 VP.n28 0.417764
R1782 VP.n56 VP.n0 0.417764
R1783 VP VP.n56 0.394061
R1784 VP.n16 VP.n15 0.189894
R1785 VP.n17 VP.n16 0.189894
R1786 VP.n17 VP.n10 0.189894
R1787 VP.n21 VP.n10 0.189894
R1788 VP.n22 VP.n21 0.189894
R1789 VP.n23 VP.n22 0.189894
R1790 VP.n23 VP.n8 0.189894
R1791 VP.n32 VP.n31 0.189894
R1792 VP.n33 VP.n32 0.189894
R1793 VP.n33 VP.n6 0.189894
R1794 VP.n37 VP.n6 0.189894
R1795 VP.n38 VP.n37 0.189894
R1796 VP.n39 VP.n38 0.189894
R1797 VP.n39 VP.n4 0.189894
R1798 VP.n44 VP.n4 0.189894
R1799 VP.n45 VP.n44 0.189894
R1800 VP.n46 VP.n45 0.189894
R1801 VP.n46 VP.n2 0.189894
R1802 VP.n50 VP.n2 0.189894
R1803 VP.n51 VP.n50 0.189894
R1804 VP.n52 VP.n51 0.189894
R1805 VP.n52 VP.n0 0.189894
R1806 VTAIL.n7 VTAIL.t11 52.0325
R1807 VTAIL.n10 VTAIL.t6 52.0324
R1808 VTAIL.n11 VTAIL.t2 52.0324
R1809 VTAIL.n2 VTAIL.t8 52.0324
R1810 VTAIL.n9 VTAIL.n8 50.0121
R1811 VTAIL.n6 VTAIL.n5 50.0121
R1812 VTAIL.n1 VTAIL.n0 50.0119
R1813 VTAIL.n4 VTAIL.n3 50.0119
R1814 VTAIL.n6 VTAIL.n4 28.0565
R1815 VTAIL.n11 VTAIL.n10 24.4358
R1816 VTAIL.n7 VTAIL.n6 3.62119
R1817 VTAIL.n10 VTAIL.n9 3.62119
R1818 VTAIL.n4 VTAIL.n2 3.62119
R1819 VTAIL VTAIL.n11 2.65783
R1820 VTAIL.n9 VTAIL.n7 2.28067
R1821 VTAIL.n2 VTAIL.n1 2.28067
R1822 VTAIL.n0 VTAIL.t3 2.02091
R1823 VTAIL.n0 VTAIL.t1 2.02091
R1824 VTAIL.n3 VTAIL.t5 2.02091
R1825 VTAIL.n3 VTAIL.t10 2.02091
R1826 VTAIL.n8 VTAIL.t7 2.02091
R1827 VTAIL.n8 VTAIL.t9 2.02091
R1828 VTAIL.n5 VTAIL.t0 2.02091
R1829 VTAIL.n5 VTAIL.t4 2.02091
R1830 VTAIL VTAIL.n1 0.963862
R1831 VDD1 VDD1.t1 71.4849
R1832 VDD1.n1 VDD1.t5 71.3713
R1833 VDD1.n1 VDD1.n0 67.5405
R1834 VDD1.n3 VDD1.n2 66.6907
R1835 VDD1.n3 VDD1.n1 46.3242
R1836 VDD1.n2 VDD1.t4 2.02091
R1837 VDD1.n2 VDD1.t2 2.02091
R1838 VDD1.n0 VDD1.t0 2.02091
R1839 VDD1.n0 VDD1.t3 2.02091
R1840 VDD1 VDD1.n3 0.847483
R1841 VN.n37 VN.n20 161.3
R1842 VN.n36 VN.n35 161.3
R1843 VN.n34 VN.n21 161.3
R1844 VN.n33 VN.n32 161.3
R1845 VN.n31 VN.n22 161.3
R1846 VN.n30 VN.n29 161.3
R1847 VN.n28 VN.n23 161.3
R1848 VN.n27 VN.n26 161.3
R1849 VN.n17 VN.n0 161.3
R1850 VN.n16 VN.n15 161.3
R1851 VN.n14 VN.n1 161.3
R1852 VN.n13 VN.n12 161.3
R1853 VN.n11 VN.n2 161.3
R1854 VN.n10 VN.n9 161.3
R1855 VN.n8 VN.n3 161.3
R1856 VN.n7 VN.n6 161.3
R1857 VN.n4 VN.t2 93.1318
R1858 VN.n24 VN.t3 93.1318
R1859 VN.n5 VN.n4 62.7067
R1860 VN.n25 VN.n24 62.7067
R1861 VN.n5 VN.t4 61.0289
R1862 VN.n18 VN.t5 61.0289
R1863 VN.n25 VN.t1 61.0289
R1864 VN.n38 VN.t0 61.0289
R1865 VN.n19 VN.n18 60.0765
R1866 VN.n39 VN.n38 60.0765
R1867 VN.n12 VN.n11 55.0167
R1868 VN.n32 VN.n31 55.0167
R1869 VN VN.n39 52.2691
R1870 VN.n12 VN.n1 25.8045
R1871 VN.n32 VN.n21 25.8045
R1872 VN.n6 VN.n3 24.3439
R1873 VN.n10 VN.n3 24.3439
R1874 VN.n11 VN.n10 24.3439
R1875 VN.n16 VN.n1 24.3439
R1876 VN.n17 VN.n16 24.3439
R1877 VN.n31 VN.n30 24.3439
R1878 VN.n30 VN.n23 24.3439
R1879 VN.n26 VN.n23 24.3439
R1880 VN.n37 VN.n36 24.3439
R1881 VN.n36 VN.n21 24.3439
R1882 VN.n18 VN.n17 21.9096
R1883 VN.n38 VN.n37 21.9096
R1884 VN.n6 VN.n5 12.1722
R1885 VN.n26 VN.n25 12.1722
R1886 VN.n27 VN.n24 2.63305
R1887 VN.n7 VN.n4 2.63305
R1888 VN.n39 VN.n20 0.417764
R1889 VN.n19 VN.n0 0.417764
R1890 VN VN.n19 0.394061
R1891 VN.n35 VN.n20 0.189894
R1892 VN.n35 VN.n34 0.189894
R1893 VN.n34 VN.n33 0.189894
R1894 VN.n33 VN.n22 0.189894
R1895 VN.n29 VN.n22 0.189894
R1896 VN.n29 VN.n28 0.189894
R1897 VN.n28 VN.n27 0.189894
R1898 VN.n8 VN.n7 0.189894
R1899 VN.n9 VN.n8 0.189894
R1900 VN.n9 VN.n2 0.189894
R1901 VN.n13 VN.n2 0.189894
R1902 VN.n14 VN.n13 0.189894
R1903 VN.n15 VN.n14 0.189894
R1904 VN.n15 VN.n0 0.189894
R1905 VDD2.n1 VDD2.t3 71.3713
R1906 VDD2.n2 VDD2.t5 68.7112
R1907 VDD2.n1 VDD2.n0 67.5405
R1908 VDD2 VDD2.n3 67.5377
R1909 VDD2.n2 VDD2.n1 43.9308
R1910 VDD2 VDD2.n2 2.77421
R1911 VDD2.n3 VDD2.t4 2.02091
R1912 VDD2.n3 VDD2.t2 2.02091
R1913 VDD2.n0 VDD2.t1 2.02091
R1914 VDD2.n0 VDD2.t0 2.02091
C0 VP VDD1 6.33354f
C1 VDD2 VTAIL 7.56217f
C2 VN VDD1 0.152207f
C3 VP VDD2 0.565121f
C4 VN VDD2 5.92288f
C5 VP VTAIL 6.50874f
C6 VN VTAIL 6.49403f
C7 VN VP 7.76348f
C8 VDD2 VDD1 1.90291f
C9 VDD1 VTAIL 7.50148f
C10 VDD2 B 6.569115f
C11 VDD1 B 6.950761f
C12 VTAIL B 7.72081f
C13 VN B 16.50189f
C14 VP B 15.235332f
C15 VDD2.t3 B 1.88639f
C16 VDD2.t1 B 0.166661f
C17 VDD2.t0 B 0.166661f
C18 VDD2.n0 B 1.47412f
C19 VDD2.n1 B 2.84257f
C20 VDD2.t5 B 1.87083f
C21 VDD2.n2 B 2.54933f
C22 VDD2.t4 B 0.166661f
C23 VDD2.t2 B 0.166661f
C24 VDD2.n3 B 1.47408f
C25 VN.n0 B 0.035209f
C26 VN.t5 B 1.92127f
C27 VN.n1 B 0.035972f
C28 VN.n2 B 0.018713f
C29 VN.n3 B 0.035051f
C30 VN.t2 B 2.2069f
C31 VN.n4 B 0.715759f
C32 VN.t4 B 1.92127f
C33 VN.n5 B 0.748364f
C34 VN.n6 B 0.026398f
C35 VN.n7 B 0.245954f
C36 VN.n8 B 0.018713f
C37 VN.n9 B 0.018713f
C38 VN.n10 B 0.035051f
C39 VN.n11 B 0.032542f
C40 VN.n12 B 0.021409f
C41 VN.n13 B 0.018713f
C42 VN.n14 B 0.018713f
C43 VN.n15 B 0.018713f
C44 VN.n16 B 0.035051f
C45 VN.n17 B 0.03332f
C46 VN.n18 B 0.763661f
C47 VN.n19 B 0.056991f
C48 VN.n20 B 0.035209f
C49 VN.t0 B 1.92127f
C50 VN.n21 B 0.035972f
C51 VN.n22 B 0.018713f
C52 VN.n23 B 0.035051f
C53 VN.t3 B 2.2069f
C54 VN.n24 B 0.715759f
C55 VN.t1 B 1.92127f
C56 VN.n25 B 0.748364f
C57 VN.n26 B 0.026398f
C58 VN.n27 B 0.245954f
C59 VN.n28 B 0.018713f
C60 VN.n29 B 0.018713f
C61 VN.n30 B 0.035051f
C62 VN.n31 B 0.032542f
C63 VN.n32 B 0.021409f
C64 VN.n33 B 0.018713f
C65 VN.n34 B 0.018713f
C66 VN.n35 B 0.018713f
C67 VN.n36 B 0.035051f
C68 VN.n37 B 0.03332f
C69 VN.n38 B 0.763661f
C70 VN.n39 B 1.15972f
C71 VDD1.t1 B 1.91798f
C72 VDD1.t5 B 1.91702f
C73 VDD1.t0 B 0.169368f
C74 VDD1.t3 B 0.169368f
C75 VDD1.n0 B 1.49805f
C76 VDD1.n1 B 3.02509f
C77 VDD1.t4 B 0.169368f
C78 VDD1.t2 B 0.169368f
C79 VDD1.n2 B 1.49176f
C80 VDD1.n3 B 2.60205f
C81 VTAIL.t3 B 0.197585f
C82 VTAIL.t1 B 0.197585f
C83 VTAIL.n0 B 1.67366f
C84 VTAIL.n1 B 0.503289f
C85 VTAIL.t8 B 2.13428f
C86 VTAIL.n2 B 0.799996f
C87 VTAIL.t5 B 0.197585f
C88 VTAIL.t10 B 0.197585f
C89 VTAIL.n3 B 1.67366f
C90 VTAIL.n4 B 2.17073f
C91 VTAIL.t0 B 0.197585f
C92 VTAIL.t4 B 0.197585f
C93 VTAIL.n5 B 1.67366f
C94 VTAIL.n6 B 2.17073f
C95 VTAIL.t11 B 2.13429f
C96 VTAIL.n7 B 0.799982f
C97 VTAIL.t7 B 0.197585f
C98 VTAIL.t9 B 0.197585f
C99 VTAIL.n8 B 1.67366f
C100 VTAIL.n9 B 0.721746f
C101 VTAIL.t6 B 2.13428f
C102 VTAIL.n10 B 1.95131f
C103 VTAIL.t2 B 2.13428f
C104 VTAIL.n11 B 1.87212f
C105 VP.n0 B 0.035953f
C106 VP.t2 B 1.96187f
C107 VP.n1 B 0.036732f
C108 VP.n2 B 0.019108f
C109 VP.n3 B 0.035792f
C110 VP.n4 B 0.019108f
C111 VP.t5 B 1.96187f
C112 VP.n5 B 0.035792f
C113 VP.n6 B 0.019108f
C114 VP.n7 B 0.035792f
C115 VP.n8 B 0.035953f
C116 VP.t3 B 1.96187f
C117 VP.n9 B 0.036732f
C118 VP.n10 B 0.019108f
C119 VP.n11 B 0.035792f
C120 VP.t4 B 2.25353f
C121 VP.n12 B 0.730886f
C122 VP.t1 B 1.96187f
C123 VP.n13 B 0.764178f
C124 VP.n14 B 0.026956f
C125 VP.n15 B 0.251152f
C126 VP.n16 B 0.019108f
C127 VP.n17 B 0.019108f
C128 VP.n18 B 0.035792f
C129 VP.n19 B 0.03323f
C130 VP.n20 B 0.021862f
C131 VP.n21 B 0.019108f
C132 VP.n22 B 0.019108f
C133 VP.n23 B 0.019108f
C134 VP.n24 B 0.035792f
C135 VP.n25 B 0.034024f
C136 VP.n26 B 0.779799f
C137 VP.n27 B 1.17939f
C138 VP.n28 B 1.1925f
C139 VP.t0 B 1.96187f
C140 VP.n29 B 0.779799f
C141 VP.n30 B 0.034024f
C142 VP.n31 B 0.035953f
C143 VP.n32 B 0.019108f
C144 VP.n33 B 0.019108f
C145 VP.n34 B 0.036732f
C146 VP.n35 B 0.021862f
C147 VP.n36 B 0.03323f
C148 VP.n37 B 0.019108f
C149 VP.n38 B 0.019108f
C150 VP.n39 B 0.019108f
C151 VP.n40 B 0.035792f
C152 VP.n41 B 0.026956f
C153 VP.n42 B 0.694654f
C154 VP.n43 B 0.026956f
C155 VP.n44 B 0.019108f
C156 VP.n45 B 0.019108f
C157 VP.n46 B 0.019108f
C158 VP.n47 B 0.035792f
C159 VP.n48 B 0.03323f
C160 VP.n49 B 0.021862f
C161 VP.n50 B 0.019108f
C162 VP.n51 B 0.019108f
C163 VP.n52 B 0.019108f
C164 VP.n53 B 0.035792f
C165 VP.n54 B 0.034024f
C166 VP.n55 B 0.779799f
C167 VP.n56 B 0.058196f
.ends

