* NGSPICE file created from diff_pair_sample_0742.ext - technology: sky130A

.subckt diff_pair_sample_0742 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=1.53945 ps=9.66 w=9.33 l=2.63
X1 VDD1.t3 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=3.6387 ps=19.44 w=9.33 l=2.63
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=0 ps=0 w=9.33 l=2.63
X3 VTAIL.t9 VP.t2 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=1.53945 ps=9.66 w=9.33 l=2.63
X4 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=1.53945 ps=9.66 w=9.33 l=2.63
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=0 ps=0 w=9.33 l=2.63
X6 VTAIL.t2 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=1.53945 ps=9.66 w=9.33 l=2.63
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=0 ps=0 w=9.33 l=2.63
X8 VDD2.t3 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=3.6387 ps=19.44 w=9.33 l=2.63
X9 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=1.53945 ps=9.66 w=9.33 l=2.63
X10 VDD1.t1 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=1.53945 ps=9.66 w=9.33 l=2.63
X11 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=1.53945 ps=9.66 w=9.33 l=2.63
X12 VDD2.t0 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=3.6387 ps=19.44 w=9.33 l=2.63
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=0 ps=0 w=9.33 l=2.63
X14 VDD1.t2 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.53945 pd=9.66 as=3.6387 ps=19.44 w=9.33 l=2.63
X15 VDD1.t4 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6387 pd=19.44 as=1.53945 ps=9.66 w=9.33 l=2.63
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n7 161.3
R6 VP.n42 VP.n0 161.3
R7 VP.n41 VP.n40 161.3
R8 VP.n39 VP.n1 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n36 VP.n2 161.3
R11 VP.n35 VP.n34 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n11 VP.t3 119.18
R19 VP.n24 VP.n23 100.481
R20 VP.n44 VP.n43 100.481
R21 VP.n22 VP.n21 100.481
R22 VP.n24 VP.t5 85.4959
R23 VP.n3 VP.t0 85.4959
R24 VP.n43 VP.t4 85.4959
R25 VP.n21 VP.t1 85.4959
R26 VP.n10 VP.t2 85.4959
R27 VP.n11 VP.n10 60.2369
R28 VP.n30 VP.n5 56.5193
R29 VP.n37 VP.n1 56.5193
R30 VP.n15 VP.n8 56.5193
R31 VP.n23 VP.n22 46.8026
R32 VP.n26 VP.n25 24.4675
R33 VP.n26 VP.n5 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n32 VP.n31 24.4675
R36 VP.n36 VP.n35 24.4675
R37 VP.n37 VP.n36 24.4675
R38 VP.n41 VP.n1 24.4675
R39 VP.n42 VP.n41 24.4675
R40 VP.n19 VP.n8 24.4675
R41 VP.n20 VP.n19 24.4675
R42 VP.n14 VP.n13 24.4675
R43 VP.n15 VP.n14 24.4675
R44 VP.n32 VP.n3 12.234
R45 VP.n35 VP.n3 12.234
R46 VP.n13 VP.n10 12.234
R47 VP.n25 VP.n24 10.2766
R48 VP.n43 VP.n42 10.2766
R49 VP.n21 VP.n20 10.2766
R50 VP.n12 VP.n11 6.83261
R51 VP.n22 VP.n7 0.278367
R52 VP.n23 VP.n6 0.278367
R53 VP.n44 VP.n0 0.278367
R54 VP.n12 VP.n9 0.189894
R55 VP.n16 VP.n9 0.189894
R56 VP.n17 VP.n16 0.189894
R57 VP.n18 VP.n17 0.189894
R58 VP.n18 VP.n7 0.189894
R59 VP.n27 VP.n6 0.189894
R60 VP.n28 VP.n27 0.189894
R61 VP.n29 VP.n28 0.189894
R62 VP.n29 VP.n4 0.189894
R63 VP.n33 VP.n4 0.189894
R64 VP.n34 VP.n33 0.189894
R65 VP.n34 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP VP.n44 0.153454
R71 VDD1.n44 VDD1.n0 289.615
R72 VDD1.n93 VDD1.n49 289.615
R73 VDD1.n45 VDD1.n44 185
R74 VDD1.n43 VDD1.n42 185
R75 VDD1.n4 VDD1.n3 185
R76 VDD1.n8 VDD1.n6 185
R77 VDD1.n37 VDD1.n36 185
R78 VDD1.n35 VDD1.n34 185
R79 VDD1.n10 VDD1.n9 185
R80 VDD1.n29 VDD1.n28 185
R81 VDD1.n27 VDD1.n26 185
R82 VDD1.n14 VDD1.n13 185
R83 VDD1.n21 VDD1.n20 185
R84 VDD1.n19 VDD1.n18 185
R85 VDD1.n66 VDD1.n65 185
R86 VDD1.n68 VDD1.n67 185
R87 VDD1.n61 VDD1.n60 185
R88 VDD1.n74 VDD1.n73 185
R89 VDD1.n76 VDD1.n75 185
R90 VDD1.n57 VDD1.n56 185
R91 VDD1.n83 VDD1.n82 185
R92 VDD1.n84 VDD1.n55 185
R93 VDD1.n86 VDD1.n85 185
R94 VDD1.n53 VDD1.n52 185
R95 VDD1.n92 VDD1.n91 185
R96 VDD1.n94 VDD1.n93 185
R97 VDD1.n17 VDD1.t1 149.524
R98 VDD1.n64 VDD1.t4 149.524
R99 VDD1.n44 VDD1.n43 104.615
R100 VDD1.n43 VDD1.n3 104.615
R101 VDD1.n8 VDD1.n3 104.615
R102 VDD1.n36 VDD1.n8 104.615
R103 VDD1.n36 VDD1.n35 104.615
R104 VDD1.n35 VDD1.n9 104.615
R105 VDD1.n28 VDD1.n9 104.615
R106 VDD1.n28 VDD1.n27 104.615
R107 VDD1.n27 VDD1.n13 104.615
R108 VDD1.n20 VDD1.n13 104.615
R109 VDD1.n20 VDD1.n19 104.615
R110 VDD1.n67 VDD1.n66 104.615
R111 VDD1.n67 VDD1.n60 104.615
R112 VDD1.n74 VDD1.n60 104.615
R113 VDD1.n75 VDD1.n74 104.615
R114 VDD1.n75 VDD1.n56 104.615
R115 VDD1.n83 VDD1.n56 104.615
R116 VDD1.n84 VDD1.n83 104.615
R117 VDD1.n85 VDD1.n84 104.615
R118 VDD1.n85 VDD1.n52 104.615
R119 VDD1.n92 VDD1.n52 104.615
R120 VDD1.n93 VDD1.n92 104.615
R121 VDD1.n99 VDD1.n98 65.3299
R122 VDD1.n101 VDD1.n100 64.7473
R123 VDD1 VDD1.n48 52.5816
R124 VDD1.n99 VDD1.n97 52.468
R125 VDD1.n19 VDD1.t1 52.3082
R126 VDD1.n66 VDD1.t4 52.3082
R127 VDD1.n101 VDD1.n99 41.9104
R128 VDD1.n6 VDD1.n4 13.1884
R129 VDD1.n86 VDD1.n53 13.1884
R130 VDD1.n42 VDD1.n41 12.8005
R131 VDD1.n38 VDD1.n37 12.8005
R132 VDD1.n87 VDD1.n55 12.8005
R133 VDD1.n91 VDD1.n90 12.8005
R134 VDD1.n45 VDD1.n2 12.0247
R135 VDD1.n34 VDD1.n7 12.0247
R136 VDD1.n82 VDD1.n81 12.0247
R137 VDD1.n94 VDD1.n51 12.0247
R138 VDD1.n46 VDD1.n0 11.249
R139 VDD1.n33 VDD1.n10 11.249
R140 VDD1.n80 VDD1.n57 11.249
R141 VDD1.n95 VDD1.n49 11.249
R142 VDD1.n30 VDD1.n29 10.4732
R143 VDD1.n77 VDD1.n76 10.4732
R144 VDD1.n18 VDD1.n17 10.2747
R145 VDD1.n65 VDD1.n64 10.2747
R146 VDD1.n26 VDD1.n12 9.69747
R147 VDD1.n73 VDD1.n59 9.69747
R148 VDD1.n48 VDD1.n47 9.45567
R149 VDD1.n97 VDD1.n96 9.45567
R150 VDD1.n16 VDD1.n15 9.3005
R151 VDD1.n23 VDD1.n22 9.3005
R152 VDD1.n25 VDD1.n24 9.3005
R153 VDD1.n12 VDD1.n11 9.3005
R154 VDD1.n31 VDD1.n30 9.3005
R155 VDD1.n33 VDD1.n32 9.3005
R156 VDD1.n7 VDD1.n5 9.3005
R157 VDD1.n39 VDD1.n38 9.3005
R158 VDD1.n47 VDD1.n46 9.3005
R159 VDD1.n2 VDD1.n1 9.3005
R160 VDD1.n41 VDD1.n40 9.3005
R161 VDD1.n96 VDD1.n95 9.3005
R162 VDD1.n51 VDD1.n50 9.3005
R163 VDD1.n90 VDD1.n89 9.3005
R164 VDD1.n63 VDD1.n62 9.3005
R165 VDD1.n70 VDD1.n69 9.3005
R166 VDD1.n72 VDD1.n71 9.3005
R167 VDD1.n59 VDD1.n58 9.3005
R168 VDD1.n78 VDD1.n77 9.3005
R169 VDD1.n80 VDD1.n79 9.3005
R170 VDD1.n81 VDD1.n54 9.3005
R171 VDD1.n88 VDD1.n87 9.3005
R172 VDD1.n25 VDD1.n14 8.92171
R173 VDD1.n72 VDD1.n61 8.92171
R174 VDD1.n22 VDD1.n21 8.14595
R175 VDD1.n69 VDD1.n68 8.14595
R176 VDD1.n18 VDD1.n16 7.3702
R177 VDD1.n65 VDD1.n63 7.3702
R178 VDD1.n21 VDD1.n16 5.81868
R179 VDD1.n68 VDD1.n63 5.81868
R180 VDD1.n22 VDD1.n14 5.04292
R181 VDD1.n69 VDD1.n61 5.04292
R182 VDD1.n26 VDD1.n25 4.26717
R183 VDD1.n73 VDD1.n72 4.26717
R184 VDD1.n29 VDD1.n12 3.49141
R185 VDD1.n76 VDD1.n59 3.49141
R186 VDD1.n17 VDD1.n15 2.84303
R187 VDD1.n64 VDD1.n62 2.84303
R188 VDD1.n48 VDD1.n0 2.71565
R189 VDD1.n30 VDD1.n10 2.71565
R190 VDD1.n77 VDD1.n57 2.71565
R191 VDD1.n97 VDD1.n49 2.71565
R192 VDD1.n100 VDD1.t0 2.12269
R193 VDD1.n100 VDD1.t3 2.12269
R194 VDD1.n98 VDD1.t5 2.12269
R195 VDD1.n98 VDD1.t2 2.12269
R196 VDD1.n46 VDD1.n45 1.93989
R197 VDD1.n34 VDD1.n33 1.93989
R198 VDD1.n82 VDD1.n80 1.93989
R199 VDD1.n95 VDD1.n94 1.93989
R200 VDD1.n42 VDD1.n2 1.16414
R201 VDD1.n37 VDD1.n7 1.16414
R202 VDD1.n81 VDD1.n55 1.16414
R203 VDD1.n91 VDD1.n51 1.16414
R204 VDD1 VDD1.n101 0.580241
R205 VDD1.n41 VDD1.n4 0.388379
R206 VDD1.n38 VDD1.n6 0.388379
R207 VDD1.n87 VDD1.n86 0.388379
R208 VDD1.n90 VDD1.n53 0.388379
R209 VDD1.n47 VDD1.n1 0.155672
R210 VDD1.n40 VDD1.n1 0.155672
R211 VDD1.n40 VDD1.n39 0.155672
R212 VDD1.n39 VDD1.n5 0.155672
R213 VDD1.n32 VDD1.n5 0.155672
R214 VDD1.n32 VDD1.n31 0.155672
R215 VDD1.n31 VDD1.n11 0.155672
R216 VDD1.n24 VDD1.n11 0.155672
R217 VDD1.n24 VDD1.n23 0.155672
R218 VDD1.n23 VDD1.n15 0.155672
R219 VDD1.n70 VDD1.n62 0.155672
R220 VDD1.n71 VDD1.n70 0.155672
R221 VDD1.n71 VDD1.n58 0.155672
R222 VDD1.n78 VDD1.n58 0.155672
R223 VDD1.n79 VDD1.n78 0.155672
R224 VDD1.n79 VDD1.n54 0.155672
R225 VDD1.n88 VDD1.n54 0.155672
R226 VDD1.n89 VDD1.n88 0.155672
R227 VDD1.n89 VDD1.n50 0.155672
R228 VDD1.n96 VDD1.n50 0.155672
R229 VTAIL.n202 VTAIL.n158 289.615
R230 VTAIL.n46 VTAIL.n2 289.615
R231 VTAIL.n152 VTAIL.n108 289.615
R232 VTAIL.n100 VTAIL.n56 289.615
R233 VTAIL.n175 VTAIL.n174 185
R234 VTAIL.n177 VTAIL.n176 185
R235 VTAIL.n170 VTAIL.n169 185
R236 VTAIL.n183 VTAIL.n182 185
R237 VTAIL.n185 VTAIL.n184 185
R238 VTAIL.n166 VTAIL.n165 185
R239 VTAIL.n192 VTAIL.n191 185
R240 VTAIL.n193 VTAIL.n164 185
R241 VTAIL.n195 VTAIL.n194 185
R242 VTAIL.n162 VTAIL.n161 185
R243 VTAIL.n201 VTAIL.n200 185
R244 VTAIL.n203 VTAIL.n202 185
R245 VTAIL.n19 VTAIL.n18 185
R246 VTAIL.n21 VTAIL.n20 185
R247 VTAIL.n14 VTAIL.n13 185
R248 VTAIL.n27 VTAIL.n26 185
R249 VTAIL.n29 VTAIL.n28 185
R250 VTAIL.n10 VTAIL.n9 185
R251 VTAIL.n36 VTAIL.n35 185
R252 VTAIL.n37 VTAIL.n8 185
R253 VTAIL.n39 VTAIL.n38 185
R254 VTAIL.n6 VTAIL.n5 185
R255 VTAIL.n45 VTAIL.n44 185
R256 VTAIL.n47 VTAIL.n46 185
R257 VTAIL.n153 VTAIL.n152 185
R258 VTAIL.n151 VTAIL.n150 185
R259 VTAIL.n112 VTAIL.n111 185
R260 VTAIL.n116 VTAIL.n114 185
R261 VTAIL.n145 VTAIL.n144 185
R262 VTAIL.n143 VTAIL.n142 185
R263 VTAIL.n118 VTAIL.n117 185
R264 VTAIL.n137 VTAIL.n136 185
R265 VTAIL.n135 VTAIL.n134 185
R266 VTAIL.n122 VTAIL.n121 185
R267 VTAIL.n129 VTAIL.n128 185
R268 VTAIL.n127 VTAIL.n126 185
R269 VTAIL.n101 VTAIL.n100 185
R270 VTAIL.n99 VTAIL.n98 185
R271 VTAIL.n60 VTAIL.n59 185
R272 VTAIL.n64 VTAIL.n62 185
R273 VTAIL.n93 VTAIL.n92 185
R274 VTAIL.n91 VTAIL.n90 185
R275 VTAIL.n66 VTAIL.n65 185
R276 VTAIL.n85 VTAIL.n84 185
R277 VTAIL.n83 VTAIL.n82 185
R278 VTAIL.n70 VTAIL.n69 185
R279 VTAIL.n77 VTAIL.n76 185
R280 VTAIL.n75 VTAIL.n74 185
R281 VTAIL.n173 VTAIL.t4 149.524
R282 VTAIL.n17 VTAIL.t7 149.524
R283 VTAIL.n125 VTAIL.t10 149.524
R284 VTAIL.n73 VTAIL.t5 149.524
R285 VTAIL.n176 VTAIL.n175 104.615
R286 VTAIL.n176 VTAIL.n169 104.615
R287 VTAIL.n183 VTAIL.n169 104.615
R288 VTAIL.n184 VTAIL.n183 104.615
R289 VTAIL.n184 VTAIL.n165 104.615
R290 VTAIL.n192 VTAIL.n165 104.615
R291 VTAIL.n193 VTAIL.n192 104.615
R292 VTAIL.n194 VTAIL.n193 104.615
R293 VTAIL.n194 VTAIL.n161 104.615
R294 VTAIL.n201 VTAIL.n161 104.615
R295 VTAIL.n202 VTAIL.n201 104.615
R296 VTAIL.n20 VTAIL.n19 104.615
R297 VTAIL.n20 VTAIL.n13 104.615
R298 VTAIL.n27 VTAIL.n13 104.615
R299 VTAIL.n28 VTAIL.n27 104.615
R300 VTAIL.n28 VTAIL.n9 104.615
R301 VTAIL.n36 VTAIL.n9 104.615
R302 VTAIL.n37 VTAIL.n36 104.615
R303 VTAIL.n38 VTAIL.n37 104.615
R304 VTAIL.n38 VTAIL.n5 104.615
R305 VTAIL.n45 VTAIL.n5 104.615
R306 VTAIL.n46 VTAIL.n45 104.615
R307 VTAIL.n152 VTAIL.n151 104.615
R308 VTAIL.n151 VTAIL.n111 104.615
R309 VTAIL.n116 VTAIL.n111 104.615
R310 VTAIL.n144 VTAIL.n116 104.615
R311 VTAIL.n144 VTAIL.n143 104.615
R312 VTAIL.n143 VTAIL.n117 104.615
R313 VTAIL.n136 VTAIL.n117 104.615
R314 VTAIL.n136 VTAIL.n135 104.615
R315 VTAIL.n135 VTAIL.n121 104.615
R316 VTAIL.n128 VTAIL.n121 104.615
R317 VTAIL.n128 VTAIL.n127 104.615
R318 VTAIL.n100 VTAIL.n99 104.615
R319 VTAIL.n99 VTAIL.n59 104.615
R320 VTAIL.n64 VTAIL.n59 104.615
R321 VTAIL.n92 VTAIL.n64 104.615
R322 VTAIL.n92 VTAIL.n91 104.615
R323 VTAIL.n91 VTAIL.n65 104.615
R324 VTAIL.n84 VTAIL.n65 104.615
R325 VTAIL.n84 VTAIL.n83 104.615
R326 VTAIL.n83 VTAIL.n69 104.615
R327 VTAIL.n76 VTAIL.n69 104.615
R328 VTAIL.n76 VTAIL.n75 104.615
R329 VTAIL.n175 VTAIL.t4 52.3082
R330 VTAIL.n19 VTAIL.t7 52.3082
R331 VTAIL.n127 VTAIL.t10 52.3082
R332 VTAIL.n75 VTAIL.t5 52.3082
R333 VTAIL.n107 VTAIL.n106 48.0687
R334 VTAIL.n55 VTAIL.n54 48.0687
R335 VTAIL.n1 VTAIL.n0 48.0685
R336 VTAIL.n53 VTAIL.n52 48.0685
R337 VTAIL.n207 VTAIL.n206 33.9308
R338 VTAIL.n51 VTAIL.n50 33.9308
R339 VTAIL.n157 VTAIL.n156 33.9308
R340 VTAIL.n105 VTAIL.n104 33.9308
R341 VTAIL.n55 VTAIL.n53 25.5134
R342 VTAIL.n207 VTAIL.n157 22.9617
R343 VTAIL.n195 VTAIL.n162 13.1884
R344 VTAIL.n39 VTAIL.n6 13.1884
R345 VTAIL.n114 VTAIL.n112 13.1884
R346 VTAIL.n62 VTAIL.n60 13.1884
R347 VTAIL.n196 VTAIL.n164 12.8005
R348 VTAIL.n200 VTAIL.n199 12.8005
R349 VTAIL.n40 VTAIL.n8 12.8005
R350 VTAIL.n44 VTAIL.n43 12.8005
R351 VTAIL.n150 VTAIL.n149 12.8005
R352 VTAIL.n146 VTAIL.n145 12.8005
R353 VTAIL.n98 VTAIL.n97 12.8005
R354 VTAIL.n94 VTAIL.n93 12.8005
R355 VTAIL.n191 VTAIL.n190 12.0247
R356 VTAIL.n203 VTAIL.n160 12.0247
R357 VTAIL.n35 VTAIL.n34 12.0247
R358 VTAIL.n47 VTAIL.n4 12.0247
R359 VTAIL.n153 VTAIL.n110 12.0247
R360 VTAIL.n142 VTAIL.n115 12.0247
R361 VTAIL.n101 VTAIL.n58 12.0247
R362 VTAIL.n90 VTAIL.n63 12.0247
R363 VTAIL.n189 VTAIL.n166 11.249
R364 VTAIL.n204 VTAIL.n158 11.249
R365 VTAIL.n33 VTAIL.n10 11.249
R366 VTAIL.n48 VTAIL.n2 11.249
R367 VTAIL.n154 VTAIL.n108 11.249
R368 VTAIL.n141 VTAIL.n118 11.249
R369 VTAIL.n102 VTAIL.n56 11.249
R370 VTAIL.n89 VTAIL.n66 11.249
R371 VTAIL.n186 VTAIL.n185 10.4732
R372 VTAIL.n30 VTAIL.n29 10.4732
R373 VTAIL.n138 VTAIL.n137 10.4732
R374 VTAIL.n86 VTAIL.n85 10.4732
R375 VTAIL.n174 VTAIL.n173 10.2747
R376 VTAIL.n18 VTAIL.n17 10.2747
R377 VTAIL.n126 VTAIL.n125 10.2747
R378 VTAIL.n74 VTAIL.n73 10.2747
R379 VTAIL.n182 VTAIL.n168 9.69747
R380 VTAIL.n26 VTAIL.n12 9.69747
R381 VTAIL.n134 VTAIL.n120 9.69747
R382 VTAIL.n82 VTAIL.n68 9.69747
R383 VTAIL.n206 VTAIL.n205 9.45567
R384 VTAIL.n50 VTAIL.n49 9.45567
R385 VTAIL.n156 VTAIL.n155 9.45567
R386 VTAIL.n104 VTAIL.n103 9.45567
R387 VTAIL.n205 VTAIL.n204 9.3005
R388 VTAIL.n160 VTAIL.n159 9.3005
R389 VTAIL.n199 VTAIL.n198 9.3005
R390 VTAIL.n172 VTAIL.n171 9.3005
R391 VTAIL.n179 VTAIL.n178 9.3005
R392 VTAIL.n181 VTAIL.n180 9.3005
R393 VTAIL.n168 VTAIL.n167 9.3005
R394 VTAIL.n187 VTAIL.n186 9.3005
R395 VTAIL.n189 VTAIL.n188 9.3005
R396 VTAIL.n190 VTAIL.n163 9.3005
R397 VTAIL.n197 VTAIL.n196 9.3005
R398 VTAIL.n49 VTAIL.n48 9.3005
R399 VTAIL.n4 VTAIL.n3 9.3005
R400 VTAIL.n43 VTAIL.n42 9.3005
R401 VTAIL.n16 VTAIL.n15 9.3005
R402 VTAIL.n23 VTAIL.n22 9.3005
R403 VTAIL.n25 VTAIL.n24 9.3005
R404 VTAIL.n12 VTAIL.n11 9.3005
R405 VTAIL.n31 VTAIL.n30 9.3005
R406 VTAIL.n33 VTAIL.n32 9.3005
R407 VTAIL.n34 VTAIL.n7 9.3005
R408 VTAIL.n41 VTAIL.n40 9.3005
R409 VTAIL.n124 VTAIL.n123 9.3005
R410 VTAIL.n131 VTAIL.n130 9.3005
R411 VTAIL.n133 VTAIL.n132 9.3005
R412 VTAIL.n120 VTAIL.n119 9.3005
R413 VTAIL.n139 VTAIL.n138 9.3005
R414 VTAIL.n141 VTAIL.n140 9.3005
R415 VTAIL.n115 VTAIL.n113 9.3005
R416 VTAIL.n147 VTAIL.n146 9.3005
R417 VTAIL.n155 VTAIL.n154 9.3005
R418 VTAIL.n110 VTAIL.n109 9.3005
R419 VTAIL.n149 VTAIL.n148 9.3005
R420 VTAIL.n72 VTAIL.n71 9.3005
R421 VTAIL.n79 VTAIL.n78 9.3005
R422 VTAIL.n81 VTAIL.n80 9.3005
R423 VTAIL.n68 VTAIL.n67 9.3005
R424 VTAIL.n87 VTAIL.n86 9.3005
R425 VTAIL.n89 VTAIL.n88 9.3005
R426 VTAIL.n63 VTAIL.n61 9.3005
R427 VTAIL.n95 VTAIL.n94 9.3005
R428 VTAIL.n103 VTAIL.n102 9.3005
R429 VTAIL.n58 VTAIL.n57 9.3005
R430 VTAIL.n97 VTAIL.n96 9.3005
R431 VTAIL.n181 VTAIL.n170 8.92171
R432 VTAIL.n25 VTAIL.n14 8.92171
R433 VTAIL.n133 VTAIL.n122 8.92171
R434 VTAIL.n81 VTAIL.n70 8.92171
R435 VTAIL.n178 VTAIL.n177 8.14595
R436 VTAIL.n22 VTAIL.n21 8.14595
R437 VTAIL.n130 VTAIL.n129 8.14595
R438 VTAIL.n78 VTAIL.n77 8.14595
R439 VTAIL.n174 VTAIL.n172 7.3702
R440 VTAIL.n18 VTAIL.n16 7.3702
R441 VTAIL.n126 VTAIL.n124 7.3702
R442 VTAIL.n74 VTAIL.n72 7.3702
R443 VTAIL.n177 VTAIL.n172 5.81868
R444 VTAIL.n21 VTAIL.n16 5.81868
R445 VTAIL.n129 VTAIL.n124 5.81868
R446 VTAIL.n77 VTAIL.n72 5.81868
R447 VTAIL.n178 VTAIL.n170 5.04292
R448 VTAIL.n22 VTAIL.n14 5.04292
R449 VTAIL.n130 VTAIL.n122 5.04292
R450 VTAIL.n78 VTAIL.n70 5.04292
R451 VTAIL.n182 VTAIL.n181 4.26717
R452 VTAIL.n26 VTAIL.n25 4.26717
R453 VTAIL.n134 VTAIL.n133 4.26717
R454 VTAIL.n82 VTAIL.n81 4.26717
R455 VTAIL.n185 VTAIL.n168 3.49141
R456 VTAIL.n29 VTAIL.n12 3.49141
R457 VTAIL.n137 VTAIL.n120 3.49141
R458 VTAIL.n85 VTAIL.n68 3.49141
R459 VTAIL.n173 VTAIL.n171 2.84303
R460 VTAIL.n17 VTAIL.n15 2.84303
R461 VTAIL.n125 VTAIL.n123 2.84303
R462 VTAIL.n73 VTAIL.n71 2.84303
R463 VTAIL.n186 VTAIL.n166 2.71565
R464 VTAIL.n206 VTAIL.n158 2.71565
R465 VTAIL.n30 VTAIL.n10 2.71565
R466 VTAIL.n50 VTAIL.n2 2.71565
R467 VTAIL.n156 VTAIL.n108 2.71565
R468 VTAIL.n138 VTAIL.n118 2.71565
R469 VTAIL.n104 VTAIL.n56 2.71565
R470 VTAIL.n86 VTAIL.n66 2.71565
R471 VTAIL.n105 VTAIL.n55 2.55222
R472 VTAIL.n157 VTAIL.n107 2.55222
R473 VTAIL.n53 VTAIL.n51 2.55222
R474 VTAIL.n0 VTAIL.t0 2.12269
R475 VTAIL.n0 VTAIL.t1 2.12269
R476 VTAIL.n52 VTAIL.t6 2.12269
R477 VTAIL.n52 VTAIL.t11 2.12269
R478 VTAIL.n106 VTAIL.t8 2.12269
R479 VTAIL.n106 VTAIL.t9 2.12269
R480 VTAIL.n54 VTAIL.t3 2.12269
R481 VTAIL.n54 VTAIL.t2 2.12269
R482 VTAIL.n191 VTAIL.n189 1.93989
R483 VTAIL.n204 VTAIL.n203 1.93989
R484 VTAIL.n35 VTAIL.n33 1.93989
R485 VTAIL.n48 VTAIL.n47 1.93989
R486 VTAIL.n154 VTAIL.n153 1.93989
R487 VTAIL.n142 VTAIL.n141 1.93989
R488 VTAIL.n102 VTAIL.n101 1.93989
R489 VTAIL.n90 VTAIL.n89 1.93989
R490 VTAIL VTAIL.n207 1.8561
R491 VTAIL.n107 VTAIL.n105 1.74619
R492 VTAIL.n51 VTAIL.n1 1.74619
R493 VTAIL.n190 VTAIL.n164 1.16414
R494 VTAIL.n200 VTAIL.n160 1.16414
R495 VTAIL.n34 VTAIL.n8 1.16414
R496 VTAIL.n44 VTAIL.n4 1.16414
R497 VTAIL.n150 VTAIL.n110 1.16414
R498 VTAIL.n145 VTAIL.n115 1.16414
R499 VTAIL.n98 VTAIL.n58 1.16414
R500 VTAIL.n93 VTAIL.n63 1.16414
R501 VTAIL VTAIL.n1 0.696621
R502 VTAIL.n196 VTAIL.n195 0.388379
R503 VTAIL.n199 VTAIL.n162 0.388379
R504 VTAIL.n40 VTAIL.n39 0.388379
R505 VTAIL.n43 VTAIL.n6 0.388379
R506 VTAIL.n149 VTAIL.n112 0.388379
R507 VTAIL.n146 VTAIL.n114 0.388379
R508 VTAIL.n97 VTAIL.n60 0.388379
R509 VTAIL.n94 VTAIL.n62 0.388379
R510 VTAIL.n179 VTAIL.n171 0.155672
R511 VTAIL.n180 VTAIL.n179 0.155672
R512 VTAIL.n180 VTAIL.n167 0.155672
R513 VTAIL.n187 VTAIL.n167 0.155672
R514 VTAIL.n188 VTAIL.n187 0.155672
R515 VTAIL.n188 VTAIL.n163 0.155672
R516 VTAIL.n197 VTAIL.n163 0.155672
R517 VTAIL.n198 VTAIL.n197 0.155672
R518 VTAIL.n198 VTAIL.n159 0.155672
R519 VTAIL.n205 VTAIL.n159 0.155672
R520 VTAIL.n23 VTAIL.n15 0.155672
R521 VTAIL.n24 VTAIL.n23 0.155672
R522 VTAIL.n24 VTAIL.n11 0.155672
R523 VTAIL.n31 VTAIL.n11 0.155672
R524 VTAIL.n32 VTAIL.n31 0.155672
R525 VTAIL.n32 VTAIL.n7 0.155672
R526 VTAIL.n41 VTAIL.n7 0.155672
R527 VTAIL.n42 VTAIL.n41 0.155672
R528 VTAIL.n42 VTAIL.n3 0.155672
R529 VTAIL.n49 VTAIL.n3 0.155672
R530 VTAIL.n155 VTAIL.n109 0.155672
R531 VTAIL.n148 VTAIL.n109 0.155672
R532 VTAIL.n148 VTAIL.n147 0.155672
R533 VTAIL.n147 VTAIL.n113 0.155672
R534 VTAIL.n140 VTAIL.n113 0.155672
R535 VTAIL.n140 VTAIL.n139 0.155672
R536 VTAIL.n139 VTAIL.n119 0.155672
R537 VTAIL.n132 VTAIL.n119 0.155672
R538 VTAIL.n132 VTAIL.n131 0.155672
R539 VTAIL.n131 VTAIL.n123 0.155672
R540 VTAIL.n103 VTAIL.n57 0.155672
R541 VTAIL.n96 VTAIL.n57 0.155672
R542 VTAIL.n96 VTAIL.n95 0.155672
R543 VTAIL.n95 VTAIL.n61 0.155672
R544 VTAIL.n88 VTAIL.n61 0.155672
R545 VTAIL.n88 VTAIL.n87 0.155672
R546 VTAIL.n87 VTAIL.n67 0.155672
R547 VTAIL.n80 VTAIL.n67 0.155672
R548 VTAIL.n80 VTAIL.n79 0.155672
R549 VTAIL.n79 VTAIL.n71 0.155672
R550 B.n740 B.n739 585
R551 B.n741 B.n740 585
R552 B.n273 B.n119 585
R553 B.n272 B.n271 585
R554 B.n270 B.n269 585
R555 B.n268 B.n267 585
R556 B.n266 B.n265 585
R557 B.n264 B.n263 585
R558 B.n262 B.n261 585
R559 B.n260 B.n259 585
R560 B.n258 B.n257 585
R561 B.n256 B.n255 585
R562 B.n254 B.n253 585
R563 B.n252 B.n251 585
R564 B.n250 B.n249 585
R565 B.n248 B.n247 585
R566 B.n246 B.n245 585
R567 B.n244 B.n243 585
R568 B.n242 B.n241 585
R569 B.n240 B.n239 585
R570 B.n238 B.n237 585
R571 B.n236 B.n235 585
R572 B.n234 B.n233 585
R573 B.n232 B.n231 585
R574 B.n230 B.n229 585
R575 B.n228 B.n227 585
R576 B.n226 B.n225 585
R577 B.n224 B.n223 585
R578 B.n222 B.n221 585
R579 B.n220 B.n219 585
R580 B.n218 B.n217 585
R581 B.n216 B.n215 585
R582 B.n214 B.n213 585
R583 B.n212 B.n211 585
R584 B.n210 B.n209 585
R585 B.n207 B.n206 585
R586 B.n205 B.n204 585
R587 B.n203 B.n202 585
R588 B.n201 B.n200 585
R589 B.n199 B.n198 585
R590 B.n197 B.n196 585
R591 B.n195 B.n194 585
R592 B.n193 B.n192 585
R593 B.n191 B.n190 585
R594 B.n189 B.n188 585
R595 B.n187 B.n186 585
R596 B.n185 B.n184 585
R597 B.n183 B.n182 585
R598 B.n181 B.n180 585
R599 B.n179 B.n178 585
R600 B.n177 B.n176 585
R601 B.n175 B.n174 585
R602 B.n173 B.n172 585
R603 B.n171 B.n170 585
R604 B.n169 B.n168 585
R605 B.n167 B.n166 585
R606 B.n165 B.n164 585
R607 B.n163 B.n162 585
R608 B.n161 B.n160 585
R609 B.n159 B.n158 585
R610 B.n157 B.n156 585
R611 B.n155 B.n154 585
R612 B.n153 B.n152 585
R613 B.n151 B.n150 585
R614 B.n149 B.n148 585
R615 B.n147 B.n146 585
R616 B.n145 B.n144 585
R617 B.n143 B.n142 585
R618 B.n141 B.n140 585
R619 B.n139 B.n138 585
R620 B.n137 B.n136 585
R621 B.n135 B.n134 585
R622 B.n133 B.n132 585
R623 B.n131 B.n130 585
R624 B.n129 B.n128 585
R625 B.n127 B.n126 585
R626 B.n81 B.n80 585
R627 B.n744 B.n743 585
R628 B.n738 B.n120 585
R629 B.n120 B.n78 585
R630 B.n737 B.n77 585
R631 B.n748 B.n77 585
R632 B.n736 B.n76 585
R633 B.n749 B.n76 585
R634 B.n735 B.n75 585
R635 B.n750 B.n75 585
R636 B.n734 B.n733 585
R637 B.n733 B.n71 585
R638 B.n732 B.n70 585
R639 B.n756 B.n70 585
R640 B.n731 B.n69 585
R641 B.n757 B.n69 585
R642 B.n730 B.n68 585
R643 B.n758 B.n68 585
R644 B.n729 B.n728 585
R645 B.n728 B.n64 585
R646 B.n727 B.n63 585
R647 B.n764 B.n63 585
R648 B.n726 B.n62 585
R649 B.n765 B.n62 585
R650 B.n725 B.n61 585
R651 B.n766 B.n61 585
R652 B.n724 B.n723 585
R653 B.n723 B.n57 585
R654 B.n722 B.n56 585
R655 B.n772 B.n56 585
R656 B.n721 B.n55 585
R657 B.n773 B.n55 585
R658 B.n720 B.n54 585
R659 B.n774 B.n54 585
R660 B.n719 B.n718 585
R661 B.n718 B.n50 585
R662 B.n717 B.n49 585
R663 B.n780 B.n49 585
R664 B.n716 B.n48 585
R665 B.n781 B.n48 585
R666 B.n715 B.n47 585
R667 B.n782 B.n47 585
R668 B.n714 B.n713 585
R669 B.n713 B.n43 585
R670 B.n712 B.n42 585
R671 B.n788 B.n42 585
R672 B.n711 B.n41 585
R673 B.n789 B.n41 585
R674 B.n710 B.n40 585
R675 B.n790 B.n40 585
R676 B.n709 B.n708 585
R677 B.n708 B.n36 585
R678 B.n707 B.n35 585
R679 B.n796 B.n35 585
R680 B.n706 B.n34 585
R681 B.n797 B.n34 585
R682 B.n705 B.n33 585
R683 B.n798 B.n33 585
R684 B.n704 B.n703 585
R685 B.n703 B.n32 585
R686 B.n702 B.n28 585
R687 B.n804 B.n28 585
R688 B.n701 B.n27 585
R689 B.n805 B.n27 585
R690 B.n700 B.n26 585
R691 B.n806 B.n26 585
R692 B.n699 B.n698 585
R693 B.n698 B.n22 585
R694 B.n697 B.n21 585
R695 B.n812 B.n21 585
R696 B.n696 B.n20 585
R697 B.n813 B.n20 585
R698 B.n695 B.n19 585
R699 B.n814 B.n19 585
R700 B.n694 B.n693 585
R701 B.n693 B.n15 585
R702 B.n692 B.n14 585
R703 B.n820 B.n14 585
R704 B.n691 B.n13 585
R705 B.n821 B.n13 585
R706 B.n690 B.n12 585
R707 B.n822 B.n12 585
R708 B.n689 B.n688 585
R709 B.n688 B.n8 585
R710 B.n687 B.n7 585
R711 B.n828 B.n7 585
R712 B.n686 B.n6 585
R713 B.n829 B.n6 585
R714 B.n685 B.n5 585
R715 B.n830 B.n5 585
R716 B.n684 B.n683 585
R717 B.n683 B.n4 585
R718 B.n682 B.n274 585
R719 B.n682 B.n681 585
R720 B.n672 B.n275 585
R721 B.n276 B.n275 585
R722 B.n674 B.n673 585
R723 B.n675 B.n674 585
R724 B.n671 B.n281 585
R725 B.n281 B.n280 585
R726 B.n670 B.n669 585
R727 B.n669 B.n668 585
R728 B.n283 B.n282 585
R729 B.n284 B.n283 585
R730 B.n661 B.n660 585
R731 B.n662 B.n661 585
R732 B.n659 B.n289 585
R733 B.n289 B.n288 585
R734 B.n658 B.n657 585
R735 B.n657 B.n656 585
R736 B.n291 B.n290 585
R737 B.n292 B.n291 585
R738 B.n649 B.n648 585
R739 B.n650 B.n649 585
R740 B.n647 B.n297 585
R741 B.n297 B.n296 585
R742 B.n646 B.n645 585
R743 B.n645 B.n644 585
R744 B.n299 B.n298 585
R745 B.n637 B.n299 585
R746 B.n636 B.n635 585
R747 B.n638 B.n636 585
R748 B.n634 B.n304 585
R749 B.n304 B.n303 585
R750 B.n633 B.n632 585
R751 B.n632 B.n631 585
R752 B.n306 B.n305 585
R753 B.n307 B.n306 585
R754 B.n624 B.n623 585
R755 B.n625 B.n624 585
R756 B.n622 B.n312 585
R757 B.n312 B.n311 585
R758 B.n621 B.n620 585
R759 B.n620 B.n619 585
R760 B.n314 B.n313 585
R761 B.n315 B.n314 585
R762 B.n612 B.n611 585
R763 B.n613 B.n612 585
R764 B.n610 B.n320 585
R765 B.n320 B.n319 585
R766 B.n609 B.n608 585
R767 B.n608 B.n607 585
R768 B.n322 B.n321 585
R769 B.n323 B.n322 585
R770 B.n600 B.n599 585
R771 B.n601 B.n600 585
R772 B.n598 B.n328 585
R773 B.n328 B.n327 585
R774 B.n597 B.n596 585
R775 B.n596 B.n595 585
R776 B.n330 B.n329 585
R777 B.n331 B.n330 585
R778 B.n588 B.n587 585
R779 B.n589 B.n588 585
R780 B.n586 B.n336 585
R781 B.n336 B.n335 585
R782 B.n585 B.n584 585
R783 B.n584 B.n583 585
R784 B.n338 B.n337 585
R785 B.n339 B.n338 585
R786 B.n576 B.n575 585
R787 B.n577 B.n576 585
R788 B.n574 B.n344 585
R789 B.n344 B.n343 585
R790 B.n573 B.n572 585
R791 B.n572 B.n571 585
R792 B.n346 B.n345 585
R793 B.n347 B.n346 585
R794 B.n564 B.n563 585
R795 B.n565 B.n564 585
R796 B.n562 B.n352 585
R797 B.n352 B.n351 585
R798 B.n561 B.n560 585
R799 B.n560 B.n559 585
R800 B.n354 B.n353 585
R801 B.n355 B.n354 585
R802 B.n555 B.n554 585
R803 B.n358 B.n357 585
R804 B.n551 B.n550 585
R805 B.n552 B.n551 585
R806 B.n549 B.n396 585
R807 B.n548 B.n547 585
R808 B.n546 B.n545 585
R809 B.n544 B.n543 585
R810 B.n542 B.n541 585
R811 B.n540 B.n539 585
R812 B.n538 B.n537 585
R813 B.n536 B.n535 585
R814 B.n534 B.n533 585
R815 B.n532 B.n531 585
R816 B.n530 B.n529 585
R817 B.n528 B.n527 585
R818 B.n526 B.n525 585
R819 B.n524 B.n523 585
R820 B.n522 B.n521 585
R821 B.n520 B.n519 585
R822 B.n518 B.n517 585
R823 B.n516 B.n515 585
R824 B.n514 B.n513 585
R825 B.n512 B.n511 585
R826 B.n510 B.n509 585
R827 B.n508 B.n507 585
R828 B.n506 B.n505 585
R829 B.n504 B.n503 585
R830 B.n502 B.n501 585
R831 B.n500 B.n499 585
R832 B.n498 B.n497 585
R833 B.n496 B.n495 585
R834 B.n494 B.n493 585
R835 B.n492 B.n491 585
R836 B.n490 B.n489 585
R837 B.n487 B.n486 585
R838 B.n485 B.n484 585
R839 B.n483 B.n482 585
R840 B.n481 B.n480 585
R841 B.n479 B.n478 585
R842 B.n477 B.n476 585
R843 B.n475 B.n474 585
R844 B.n473 B.n472 585
R845 B.n471 B.n470 585
R846 B.n469 B.n468 585
R847 B.n467 B.n466 585
R848 B.n465 B.n464 585
R849 B.n463 B.n462 585
R850 B.n461 B.n460 585
R851 B.n459 B.n458 585
R852 B.n457 B.n456 585
R853 B.n455 B.n454 585
R854 B.n453 B.n452 585
R855 B.n451 B.n450 585
R856 B.n449 B.n448 585
R857 B.n447 B.n446 585
R858 B.n445 B.n444 585
R859 B.n443 B.n442 585
R860 B.n441 B.n440 585
R861 B.n439 B.n438 585
R862 B.n437 B.n436 585
R863 B.n435 B.n434 585
R864 B.n433 B.n432 585
R865 B.n431 B.n430 585
R866 B.n429 B.n428 585
R867 B.n427 B.n426 585
R868 B.n425 B.n424 585
R869 B.n423 B.n422 585
R870 B.n421 B.n420 585
R871 B.n419 B.n418 585
R872 B.n417 B.n416 585
R873 B.n415 B.n414 585
R874 B.n413 B.n412 585
R875 B.n411 B.n410 585
R876 B.n409 B.n408 585
R877 B.n407 B.n406 585
R878 B.n405 B.n404 585
R879 B.n403 B.n402 585
R880 B.n556 B.n356 585
R881 B.n356 B.n355 585
R882 B.n558 B.n557 585
R883 B.n559 B.n558 585
R884 B.n350 B.n349 585
R885 B.n351 B.n350 585
R886 B.n567 B.n566 585
R887 B.n566 B.n565 585
R888 B.n568 B.n348 585
R889 B.n348 B.n347 585
R890 B.n570 B.n569 585
R891 B.n571 B.n570 585
R892 B.n342 B.n341 585
R893 B.n343 B.n342 585
R894 B.n579 B.n578 585
R895 B.n578 B.n577 585
R896 B.n580 B.n340 585
R897 B.n340 B.n339 585
R898 B.n582 B.n581 585
R899 B.n583 B.n582 585
R900 B.n334 B.n333 585
R901 B.n335 B.n334 585
R902 B.n591 B.n590 585
R903 B.n590 B.n589 585
R904 B.n592 B.n332 585
R905 B.n332 B.n331 585
R906 B.n594 B.n593 585
R907 B.n595 B.n594 585
R908 B.n326 B.n325 585
R909 B.n327 B.n326 585
R910 B.n603 B.n602 585
R911 B.n602 B.n601 585
R912 B.n604 B.n324 585
R913 B.n324 B.n323 585
R914 B.n606 B.n605 585
R915 B.n607 B.n606 585
R916 B.n318 B.n317 585
R917 B.n319 B.n318 585
R918 B.n615 B.n614 585
R919 B.n614 B.n613 585
R920 B.n616 B.n316 585
R921 B.n316 B.n315 585
R922 B.n618 B.n617 585
R923 B.n619 B.n618 585
R924 B.n310 B.n309 585
R925 B.n311 B.n310 585
R926 B.n627 B.n626 585
R927 B.n626 B.n625 585
R928 B.n628 B.n308 585
R929 B.n308 B.n307 585
R930 B.n630 B.n629 585
R931 B.n631 B.n630 585
R932 B.n302 B.n301 585
R933 B.n303 B.n302 585
R934 B.n640 B.n639 585
R935 B.n639 B.n638 585
R936 B.n641 B.n300 585
R937 B.n637 B.n300 585
R938 B.n643 B.n642 585
R939 B.n644 B.n643 585
R940 B.n295 B.n294 585
R941 B.n296 B.n295 585
R942 B.n652 B.n651 585
R943 B.n651 B.n650 585
R944 B.n653 B.n293 585
R945 B.n293 B.n292 585
R946 B.n655 B.n654 585
R947 B.n656 B.n655 585
R948 B.n287 B.n286 585
R949 B.n288 B.n287 585
R950 B.n664 B.n663 585
R951 B.n663 B.n662 585
R952 B.n665 B.n285 585
R953 B.n285 B.n284 585
R954 B.n667 B.n666 585
R955 B.n668 B.n667 585
R956 B.n279 B.n278 585
R957 B.n280 B.n279 585
R958 B.n677 B.n676 585
R959 B.n676 B.n675 585
R960 B.n678 B.n277 585
R961 B.n277 B.n276 585
R962 B.n680 B.n679 585
R963 B.n681 B.n680 585
R964 B.n2 B.n0 585
R965 B.n4 B.n2 585
R966 B.n3 B.n1 585
R967 B.n829 B.n3 585
R968 B.n827 B.n826 585
R969 B.n828 B.n827 585
R970 B.n825 B.n9 585
R971 B.n9 B.n8 585
R972 B.n824 B.n823 585
R973 B.n823 B.n822 585
R974 B.n11 B.n10 585
R975 B.n821 B.n11 585
R976 B.n819 B.n818 585
R977 B.n820 B.n819 585
R978 B.n817 B.n16 585
R979 B.n16 B.n15 585
R980 B.n816 B.n815 585
R981 B.n815 B.n814 585
R982 B.n18 B.n17 585
R983 B.n813 B.n18 585
R984 B.n811 B.n810 585
R985 B.n812 B.n811 585
R986 B.n809 B.n23 585
R987 B.n23 B.n22 585
R988 B.n808 B.n807 585
R989 B.n807 B.n806 585
R990 B.n25 B.n24 585
R991 B.n805 B.n25 585
R992 B.n803 B.n802 585
R993 B.n804 B.n803 585
R994 B.n801 B.n29 585
R995 B.n32 B.n29 585
R996 B.n800 B.n799 585
R997 B.n799 B.n798 585
R998 B.n31 B.n30 585
R999 B.n797 B.n31 585
R1000 B.n795 B.n794 585
R1001 B.n796 B.n795 585
R1002 B.n793 B.n37 585
R1003 B.n37 B.n36 585
R1004 B.n792 B.n791 585
R1005 B.n791 B.n790 585
R1006 B.n39 B.n38 585
R1007 B.n789 B.n39 585
R1008 B.n787 B.n786 585
R1009 B.n788 B.n787 585
R1010 B.n785 B.n44 585
R1011 B.n44 B.n43 585
R1012 B.n784 B.n783 585
R1013 B.n783 B.n782 585
R1014 B.n46 B.n45 585
R1015 B.n781 B.n46 585
R1016 B.n779 B.n778 585
R1017 B.n780 B.n779 585
R1018 B.n777 B.n51 585
R1019 B.n51 B.n50 585
R1020 B.n776 B.n775 585
R1021 B.n775 B.n774 585
R1022 B.n53 B.n52 585
R1023 B.n773 B.n53 585
R1024 B.n771 B.n770 585
R1025 B.n772 B.n771 585
R1026 B.n769 B.n58 585
R1027 B.n58 B.n57 585
R1028 B.n768 B.n767 585
R1029 B.n767 B.n766 585
R1030 B.n60 B.n59 585
R1031 B.n765 B.n60 585
R1032 B.n763 B.n762 585
R1033 B.n764 B.n763 585
R1034 B.n761 B.n65 585
R1035 B.n65 B.n64 585
R1036 B.n760 B.n759 585
R1037 B.n759 B.n758 585
R1038 B.n67 B.n66 585
R1039 B.n757 B.n67 585
R1040 B.n755 B.n754 585
R1041 B.n756 B.n755 585
R1042 B.n753 B.n72 585
R1043 B.n72 B.n71 585
R1044 B.n752 B.n751 585
R1045 B.n751 B.n750 585
R1046 B.n74 B.n73 585
R1047 B.n749 B.n74 585
R1048 B.n747 B.n746 585
R1049 B.n748 B.n747 585
R1050 B.n745 B.n79 585
R1051 B.n79 B.n78 585
R1052 B.n832 B.n831 585
R1053 B.n831 B.n830 585
R1054 B.n554 B.n356 497.305
R1055 B.n743 B.n79 497.305
R1056 B.n402 B.n354 497.305
R1057 B.n740 B.n120 497.305
R1058 B.n399 B.t6 293.587
R1059 B.n397 B.t10 293.587
R1060 B.n123 B.t17 293.587
R1061 B.n121 B.t13 293.587
R1062 B.n399 B.t9 293.536
R1063 B.n121 B.t15 293.536
R1064 B.n397 B.t12 293.536
R1065 B.n123 B.t18 293.536
R1066 B.n741 B.n118 256.663
R1067 B.n741 B.n117 256.663
R1068 B.n741 B.n116 256.663
R1069 B.n741 B.n115 256.663
R1070 B.n741 B.n114 256.663
R1071 B.n741 B.n113 256.663
R1072 B.n741 B.n112 256.663
R1073 B.n741 B.n111 256.663
R1074 B.n741 B.n110 256.663
R1075 B.n741 B.n109 256.663
R1076 B.n741 B.n108 256.663
R1077 B.n741 B.n107 256.663
R1078 B.n741 B.n106 256.663
R1079 B.n741 B.n105 256.663
R1080 B.n741 B.n104 256.663
R1081 B.n741 B.n103 256.663
R1082 B.n741 B.n102 256.663
R1083 B.n741 B.n101 256.663
R1084 B.n741 B.n100 256.663
R1085 B.n741 B.n99 256.663
R1086 B.n741 B.n98 256.663
R1087 B.n741 B.n97 256.663
R1088 B.n741 B.n96 256.663
R1089 B.n741 B.n95 256.663
R1090 B.n741 B.n94 256.663
R1091 B.n741 B.n93 256.663
R1092 B.n741 B.n92 256.663
R1093 B.n741 B.n91 256.663
R1094 B.n741 B.n90 256.663
R1095 B.n741 B.n89 256.663
R1096 B.n741 B.n88 256.663
R1097 B.n741 B.n87 256.663
R1098 B.n741 B.n86 256.663
R1099 B.n741 B.n85 256.663
R1100 B.n741 B.n84 256.663
R1101 B.n741 B.n83 256.663
R1102 B.n741 B.n82 256.663
R1103 B.n742 B.n741 256.663
R1104 B.n553 B.n552 256.663
R1105 B.n552 B.n359 256.663
R1106 B.n552 B.n360 256.663
R1107 B.n552 B.n361 256.663
R1108 B.n552 B.n362 256.663
R1109 B.n552 B.n363 256.663
R1110 B.n552 B.n364 256.663
R1111 B.n552 B.n365 256.663
R1112 B.n552 B.n366 256.663
R1113 B.n552 B.n367 256.663
R1114 B.n552 B.n368 256.663
R1115 B.n552 B.n369 256.663
R1116 B.n552 B.n370 256.663
R1117 B.n552 B.n371 256.663
R1118 B.n552 B.n372 256.663
R1119 B.n552 B.n373 256.663
R1120 B.n552 B.n374 256.663
R1121 B.n552 B.n375 256.663
R1122 B.n552 B.n376 256.663
R1123 B.n552 B.n377 256.663
R1124 B.n552 B.n378 256.663
R1125 B.n552 B.n379 256.663
R1126 B.n552 B.n380 256.663
R1127 B.n552 B.n381 256.663
R1128 B.n552 B.n382 256.663
R1129 B.n552 B.n383 256.663
R1130 B.n552 B.n384 256.663
R1131 B.n552 B.n385 256.663
R1132 B.n552 B.n386 256.663
R1133 B.n552 B.n387 256.663
R1134 B.n552 B.n388 256.663
R1135 B.n552 B.n389 256.663
R1136 B.n552 B.n390 256.663
R1137 B.n552 B.n391 256.663
R1138 B.n552 B.n392 256.663
R1139 B.n552 B.n393 256.663
R1140 B.n552 B.n394 256.663
R1141 B.n552 B.n395 256.663
R1142 B.n400 B.t8 236.13
R1143 B.n122 B.t16 236.13
R1144 B.n398 B.t11 236.13
R1145 B.n124 B.t19 236.13
R1146 B.n558 B.n356 163.367
R1147 B.n558 B.n350 163.367
R1148 B.n566 B.n350 163.367
R1149 B.n566 B.n348 163.367
R1150 B.n570 B.n348 163.367
R1151 B.n570 B.n342 163.367
R1152 B.n578 B.n342 163.367
R1153 B.n578 B.n340 163.367
R1154 B.n582 B.n340 163.367
R1155 B.n582 B.n334 163.367
R1156 B.n590 B.n334 163.367
R1157 B.n590 B.n332 163.367
R1158 B.n594 B.n332 163.367
R1159 B.n594 B.n326 163.367
R1160 B.n602 B.n326 163.367
R1161 B.n602 B.n324 163.367
R1162 B.n606 B.n324 163.367
R1163 B.n606 B.n318 163.367
R1164 B.n614 B.n318 163.367
R1165 B.n614 B.n316 163.367
R1166 B.n618 B.n316 163.367
R1167 B.n618 B.n310 163.367
R1168 B.n626 B.n310 163.367
R1169 B.n626 B.n308 163.367
R1170 B.n630 B.n308 163.367
R1171 B.n630 B.n302 163.367
R1172 B.n639 B.n302 163.367
R1173 B.n639 B.n300 163.367
R1174 B.n643 B.n300 163.367
R1175 B.n643 B.n295 163.367
R1176 B.n651 B.n295 163.367
R1177 B.n651 B.n293 163.367
R1178 B.n655 B.n293 163.367
R1179 B.n655 B.n287 163.367
R1180 B.n663 B.n287 163.367
R1181 B.n663 B.n285 163.367
R1182 B.n667 B.n285 163.367
R1183 B.n667 B.n279 163.367
R1184 B.n676 B.n279 163.367
R1185 B.n676 B.n277 163.367
R1186 B.n680 B.n277 163.367
R1187 B.n680 B.n2 163.367
R1188 B.n831 B.n2 163.367
R1189 B.n831 B.n3 163.367
R1190 B.n827 B.n3 163.367
R1191 B.n827 B.n9 163.367
R1192 B.n823 B.n9 163.367
R1193 B.n823 B.n11 163.367
R1194 B.n819 B.n11 163.367
R1195 B.n819 B.n16 163.367
R1196 B.n815 B.n16 163.367
R1197 B.n815 B.n18 163.367
R1198 B.n811 B.n18 163.367
R1199 B.n811 B.n23 163.367
R1200 B.n807 B.n23 163.367
R1201 B.n807 B.n25 163.367
R1202 B.n803 B.n25 163.367
R1203 B.n803 B.n29 163.367
R1204 B.n799 B.n29 163.367
R1205 B.n799 B.n31 163.367
R1206 B.n795 B.n31 163.367
R1207 B.n795 B.n37 163.367
R1208 B.n791 B.n37 163.367
R1209 B.n791 B.n39 163.367
R1210 B.n787 B.n39 163.367
R1211 B.n787 B.n44 163.367
R1212 B.n783 B.n44 163.367
R1213 B.n783 B.n46 163.367
R1214 B.n779 B.n46 163.367
R1215 B.n779 B.n51 163.367
R1216 B.n775 B.n51 163.367
R1217 B.n775 B.n53 163.367
R1218 B.n771 B.n53 163.367
R1219 B.n771 B.n58 163.367
R1220 B.n767 B.n58 163.367
R1221 B.n767 B.n60 163.367
R1222 B.n763 B.n60 163.367
R1223 B.n763 B.n65 163.367
R1224 B.n759 B.n65 163.367
R1225 B.n759 B.n67 163.367
R1226 B.n755 B.n67 163.367
R1227 B.n755 B.n72 163.367
R1228 B.n751 B.n72 163.367
R1229 B.n751 B.n74 163.367
R1230 B.n747 B.n74 163.367
R1231 B.n747 B.n79 163.367
R1232 B.n551 B.n358 163.367
R1233 B.n551 B.n396 163.367
R1234 B.n547 B.n546 163.367
R1235 B.n543 B.n542 163.367
R1236 B.n539 B.n538 163.367
R1237 B.n535 B.n534 163.367
R1238 B.n531 B.n530 163.367
R1239 B.n527 B.n526 163.367
R1240 B.n523 B.n522 163.367
R1241 B.n519 B.n518 163.367
R1242 B.n515 B.n514 163.367
R1243 B.n511 B.n510 163.367
R1244 B.n507 B.n506 163.367
R1245 B.n503 B.n502 163.367
R1246 B.n499 B.n498 163.367
R1247 B.n495 B.n494 163.367
R1248 B.n491 B.n490 163.367
R1249 B.n486 B.n485 163.367
R1250 B.n482 B.n481 163.367
R1251 B.n478 B.n477 163.367
R1252 B.n474 B.n473 163.367
R1253 B.n470 B.n469 163.367
R1254 B.n466 B.n465 163.367
R1255 B.n462 B.n461 163.367
R1256 B.n458 B.n457 163.367
R1257 B.n454 B.n453 163.367
R1258 B.n450 B.n449 163.367
R1259 B.n446 B.n445 163.367
R1260 B.n442 B.n441 163.367
R1261 B.n438 B.n437 163.367
R1262 B.n434 B.n433 163.367
R1263 B.n430 B.n429 163.367
R1264 B.n426 B.n425 163.367
R1265 B.n422 B.n421 163.367
R1266 B.n418 B.n417 163.367
R1267 B.n414 B.n413 163.367
R1268 B.n410 B.n409 163.367
R1269 B.n406 B.n405 163.367
R1270 B.n560 B.n354 163.367
R1271 B.n560 B.n352 163.367
R1272 B.n564 B.n352 163.367
R1273 B.n564 B.n346 163.367
R1274 B.n572 B.n346 163.367
R1275 B.n572 B.n344 163.367
R1276 B.n576 B.n344 163.367
R1277 B.n576 B.n338 163.367
R1278 B.n584 B.n338 163.367
R1279 B.n584 B.n336 163.367
R1280 B.n588 B.n336 163.367
R1281 B.n588 B.n330 163.367
R1282 B.n596 B.n330 163.367
R1283 B.n596 B.n328 163.367
R1284 B.n600 B.n328 163.367
R1285 B.n600 B.n322 163.367
R1286 B.n608 B.n322 163.367
R1287 B.n608 B.n320 163.367
R1288 B.n612 B.n320 163.367
R1289 B.n612 B.n314 163.367
R1290 B.n620 B.n314 163.367
R1291 B.n620 B.n312 163.367
R1292 B.n624 B.n312 163.367
R1293 B.n624 B.n306 163.367
R1294 B.n632 B.n306 163.367
R1295 B.n632 B.n304 163.367
R1296 B.n636 B.n304 163.367
R1297 B.n636 B.n299 163.367
R1298 B.n645 B.n299 163.367
R1299 B.n645 B.n297 163.367
R1300 B.n649 B.n297 163.367
R1301 B.n649 B.n291 163.367
R1302 B.n657 B.n291 163.367
R1303 B.n657 B.n289 163.367
R1304 B.n661 B.n289 163.367
R1305 B.n661 B.n283 163.367
R1306 B.n669 B.n283 163.367
R1307 B.n669 B.n281 163.367
R1308 B.n674 B.n281 163.367
R1309 B.n674 B.n275 163.367
R1310 B.n682 B.n275 163.367
R1311 B.n683 B.n682 163.367
R1312 B.n683 B.n5 163.367
R1313 B.n6 B.n5 163.367
R1314 B.n7 B.n6 163.367
R1315 B.n688 B.n7 163.367
R1316 B.n688 B.n12 163.367
R1317 B.n13 B.n12 163.367
R1318 B.n14 B.n13 163.367
R1319 B.n693 B.n14 163.367
R1320 B.n693 B.n19 163.367
R1321 B.n20 B.n19 163.367
R1322 B.n21 B.n20 163.367
R1323 B.n698 B.n21 163.367
R1324 B.n698 B.n26 163.367
R1325 B.n27 B.n26 163.367
R1326 B.n28 B.n27 163.367
R1327 B.n703 B.n28 163.367
R1328 B.n703 B.n33 163.367
R1329 B.n34 B.n33 163.367
R1330 B.n35 B.n34 163.367
R1331 B.n708 B.n35 163.367
R1332 B.n708 B.n40 163.367
R1333 B.n41 B.n40 163.367
R1334 B.n42 B.n41 163.367
R1335 B.n713 B.n42 163.367
R1336 B.n713 B.n47 163.367
R1337 B.n48 B.n47 163.367
R1338 B.n49 B.n48 163.367
R1339 B.n718 B.n49 163.367
R1340 B.n718 B.n54 163.367
R1341 B.n55 B.n54 163.367
R1342 B.n56 B.n55 163.367
R1343 B.n723 B.n56 163.367
R1344 B.n723 B.n61 163.367
R1345 B.n62 B.n61 163.367
R1346 B.n63 B.n62 163.367
R1347 B.n728 B.n63 163.367
R1348 B.n728 B.n68 163.367
R1349 B.n69 B.n68 163.367
R1350 B.n70 B.n69 163.367
R1351 B.n733 B.n70 163.367
R1352 B.n733 B.n75 163.367
R1353 B.n76 B.n75 163.367
R1354 B.n77 B.n76 163.367
R1355 B.n120 B.n77 163.367
R1356 B.n126 B.n81 163.367
R1357 B.n130 B.n129 163.367
R1358 B.n134 B.n133 163.367
R1359 B.n138 B.n137 163.367
R1360 B.n142 B.n141 163.367
R1361 B.n146 B.n145 163.367
R1362 B.n150 B.n149 163.367
R1363 B.n154 B.n153 163.367
R1364 B.n158 B.n157 163.367
R1365 B.n162 B.n161 163.367
R1366 B.n166 B.n165 163.367
R1367 B.n170 B.n169 163.367
R1368 B.n174 B.n173 163.367
R1369 B.n178 B.n177 163.367
R1370 B.n182 B.n181 163.367
R1371 B.n186 B.n185 163.367
R1372 B.n190 B.n189 163.367
R1373 B.n194 B.n193 163.367
R1374 B.n198 B.n197 163.367
R1375 B.n202 B.n201 163.367
R1376 B.n206 B.n205 163.367
R1377 B.n211 B.n210 163.367
R1378 B.n215 B.n214 163.367
R1379 B.n219 B.n218 163.367
R1380 B.n223 B.n222 163.367
R1381 B.n227 B.n226 163.367
R1382 B.n231 B.n230 163.367
R1383 B.n235 B.n234 163.367
R1384 B.n239 B.n238 163.367
R1385 B.n243 B.n242 163.367
R1386 B.n247 B.n246 163.367
R1387 B.n251 B.n250 163.367
R1388 B.n255 B.n254 163.367
R1389 B.n259 B.n258 163.367
R1390 B.n263 B.n262 163.367
R1391 B.n267 B.n266 163.367
R1392 B.n271 B.n270 163.367
R1393 B.n740 B.n119 163.367
R1394 B.n552 B.n355 89.6273
R1395 B.n741 B.n78 89.6273
R1396 B.n554 B.n553 71.676
R1397 B.n396 B.n359 71.676
R1398 B.n546 B.n360 71.676
R1399 B.n542 B.n361 71.676
R1400 B.n538 B.n362 71.676
R1401 B.n534 B.n363 71.676
R1402 B.n530 B.n364 71.676
R1403 B.n526 B.n365 71.676
R1404 B.n522 B.n366 71.676
R1405 B.n518 B.n367 71.676
R1406 B.n514 B.n368 71.676
R1407 B.n510 B.n369 71.676
R1408 B.n506 B.n370 71.676
R1409 B.n502 B.n371 71.676
R1410 B.n498 B.n372 71.676
R1411 B.n494 B.n373 71.676
R1412 B.n490 B.n374 71.676
R1413 B.n485 B.n375 71.676
R1414 B.n481 B.n376 71.676
R1415 B.n477 B.n377 71.676
R1416 B.n473 B.n378 71.676
R1417 B.n469 B.n379 71.676
R1418 B.n465 B.n380 71.676
R1419 B.n461 B.n381 71.676
R1420 B.n457 B.n382 71.676
R1421 B.n453 B.n383 71.676
R1422 B.n449 B.n384 71.676
R1423 B.n445 B.n385 71.676
R1424 B.n441 B.n386 71.676
R1425 B.n437 B.n387 71.676
R1426 B.n433 B.n388 71.676
R1427 B.n429 B.n389 71.676
R1428 B.n425 B.n390 71.676
R1429 B.n421 B.n391 71.676
R1430 B.n417 B.n392 71.676
R1431 B.n413 B.n393 71.676
R1432 B.n409 B.n394 71.676
R1433 B.n405 B.n395 71.676
R1434 B.n743 B.n742 71.676
R1435 B.n126 B.n82 71.676
R1436 B.n130 B.n83 71.676
R1437 B.n134 B.n84 71.676
R1438 B.n138 B.n85 71.676
R1439 B.n142 B.n86 71.676
R1440 B.n146 B.n87 71.676
R1441 B.n150 B.n88 71.676
R1442 B.n154 B.n89 71.676
R1443 B.n158 B.n90 71.676
R1444 B.n162 B.n91 71.676
R1445 B.n166 B.n92 71.676
R1446 B.n170 B.n93 71.676
R1447 B.n174 B.n94 71.676
R1448 B.n178 B.n95 71.676
R1449 B.n182 B.n96 71.676
R1450 B.n186 B.n97 71.676
R1451 B.n190 B.n98 71.676
R1452 B.n194 B.n99 71.676
R1453 B.n198 B.n100 71.676
R1454 B.n202 B.n101 71.676
R1455 B.n206 B.n102 71.676
R1456 B.n211 B.n103 71.676
R1457 B.n215 B.n104 71.676
R1458 B.n219 B.n105 71.676
R1459 B.n223 B.n106 71.676
R1460 B.n227 B.n107 71.676
R1461 B.n231 B.n108 71.676
R1462 B.n235 B.n109 71.676
R1463 B.n239 B.n110 71.676
R1464 B.n243 B.n111 71.676
R1465 B.n247 B.n112 71.676
R1466 B.n251 B.n113 71.676
R1467 B.n255 B.n114 71.676
R1468 B.n259 B.n115 71.676
R1469 B.n263 B.n116 71.676
R1470 B.n267 B.n117 71.676
R1471 B.n271 B.n118 71.676
R1472 B.n119 B.n118 71.676
R1473 B.n270 B.n117 71.676
R1474 B.n266 B.n116 71.676
R1475 B.n262 B.n115 71.676
R1476 B.n258 B.n114 71.676
R1477 B.n254 B.n113 71.676
R1478 B.n250 B.n112 71.676
R1479 B.n246 B.n111 71.676
R1480 B.n242 B.n110 71.676
R1481 B.n238 B.n109 71.676
R1482 B.n234 B.n108 71.676
R1483 B.n230 B.n107 71.676
R1484 B.n226 B.n106 71.676
R1485 B.n222 B.n105 71.676
R1486 B.n218 B.n104 71.676
R1487 B.n214 B.n103 71.676
R1488 B.n210 B.n102 71.676
R1489 B.n205 B.n101 71.676
R1490 B.n201 B.n100 71.676
R1491 B.n197 B.n99 71.676
R1492 B.n193 B.n98 71.676
R1493 B.n189 B.n97 71.676
R1494 B.n185 B.n96 71.676
R1495 B.n181 B.n95 71.676
R1496 B.n177 B.n94 71.676
R1497 B.n173 B.n93 71.676
R1498 B.n169 B.n92 71.676
R1499 B.n165 B.n91 71.676
R1500 B.n161 B.n90 71.676
R1501 B.n157 B.n89 71.676
R1502 B.n153 B.n88 71.676
R1503 B.n149 B.n87 71.676
R1504 B.n145 B.n86 71.676
R1505 B.n141 B.n85 71.676
R1506 B.n137 B.n84 71.676
R1507 B.n133 B.n83 71.676
R1508 B.n129 B.n82 71.676
R1509 B.n742 B.n81 71.676
R1510 B.n553 B.n358 71.676
R1511 B.n547 B.n359 71.676
R1512 B.n543 B.n360 71.676
R1513 B.n539 B.n361 71.676
R1514 B.n535 B.n362 71.676
R1515 B.n531 B.n363 71.676
R1516 B.n527 B.n364 71.676
R1517 B.n523 B.n365 71.676
R1518 B.n519 B.n366 71.676
R1519 B.n515 B.n367 71.676
R1520 B.n511 B.n368 71.676
R1521 B.n507 B.n369 71.676
R1522 B.n503 B.n370 71.676
R1523 B.n499 B.n371 71.676
R1524 B.n495 B.n372 71.676
R1525 B.n491 B.n373 71.676
R1526 B.n486 B.n374 71.676
R1527 B.n482 B.n375 71.676
R1528 B.n478 B.n376 71.676
R1529 B.n474 B.n377 71.676
R1530 B.n470 B.n378 71.676
R1531 B.n466 B.n379 71.676
R1532 B.n462 B.n380 71.676
R1533 B.n458 B.n381 71.676
R1534 B.n454 B.n382 71.676
R1535 B.n450 B.n383 71.676
R1536 B.n446 B.n384 71.676
R1537 B.n442 B.n385 71.676
R1538 B.n438 B.n386 71.676
R1539 B.n434 B.n387 71.676
R1540 B.n430 B.n388 71.676
R1541 B.n426 B.n389 71.676
R1542 B.n422 B.n390 71.676
R1543 B.n418 B.n391 71.676
R1544 B.n414 B.n392 71.676
R1545 B.n410 B.n393 71.676
R1546 B.n406 B.n394 71.676
R1547 B.n402 B.n395 71.676
R1548 B.n401 B.n400 59.5399
R1549 B.n488 B.n398 59.5399
R1550 B.n125 B.n124 59.5399
R1551 B.n208 B.n122 59.5399
R1552 B.n400 B.n399 57.4066
R1553 B.n398 B.n397 57.4066
R1554 B.n124 B.n123 57.4066
R1555 B.n122 B.n121 57.4066
R1556 B.n559 B.n355 51.2158
R1557 B.n559 B.n351 51.2158
R1558 B.n565 B.n351 51.2158
R1559 B.n565 B.n347 51.2158
R1560 B.n571 B.n347 51.2158
R1561 B.n571 B.n343 51.2158
R1562 B.n577 B.n343 51.2158
R1563 B.n583 B.n339 51.2158
R1564 B.n583 B.n335 51.2158
R1565 B.n589 B.n335 51.2158
R1566 B.n589 B.n331 51.2158
R1567 B.n595 B.n331 51.2158
R1568 B.n595 B.n327 51.2158
R1569 B.n601 B.n327 51.2158
R1570 B.n601 B.n323 51.2158
R1571 B.n607 B.n323 51.2158
R1572 B.n607 B.n319 51.2158
R1573 B.n613 B.n319 51.2158
R1574 B.n619 B.n315 51.2158
R1575 B.n619 B.n311 51.2158
R1576 B.n625 B.n311 51.2158
R1577 B.n625 B.n307 51.2158
R1578 B.n631 B.n307 51.2158
R1579 B.n631 B.n303 51.2158
R1580 B.n638 B.n303 51.2158
R1581 B.n638 B.n637 51.2158
R1582 B.n644 B.n296 51.2158
R1583 B.n650 B.n296 51.2158
R1584 B.n650 B.n292 51.2158
R1585 B.n656 B.n292 51.2158
R1586 B.n656 B.n288 51.2158
R1587 B.n662 B.n288 51.2158
R1588 B.n662 B.n284 51.2158
R1589 B.n668 B.n284 51.2158
R1590 B.n675 B.n280 51.2158
R1591 B.n675 B.n276 51.2158
R1592 B.n681 B.n276 51.2158
R1593 B.n681 B.n4 51.2158
R1594 B.n830 B.n4 51.2158
R1595 B.n830 B.n829 51.2158
R1596 B.n829 B.n828 51.2158
R1597 B.n828 B.n8 51.2158
R1598 B.n822 B.n8 51.2158
R1599 B.n822 B.n821 51.2158
R1600 B.n820 B.n15 51.2158
R1601 B.n814 B.n15 51.2158
R1602 B.n814 B.n813 51.2158
R1603 B.n813 B.n812 51.2158
R1604 B.n812 B.n22 51.2158
R1605 B.n806 B.n22 51.2158
R1606 B.n806 B.n805 51.2158
R1607 B.n805 B.n804 51.2158
R1608 B.n798 B.n32 51.2158
R1609 B.n798 B.n797 51.2158
R1610 B.n797 B.n796 51.2158
R1611 B.n796 B.n36 51.2158
R1612 B.n790 B.n36 51.2158
R1613 B.n790 B.n789 51.2158
R1614 B.n789 B.n788 51.2158
R1615 B.n788 B.n43 51.2158
R1616 B.n782 B.n781 51.2158
R1617 B.n781 B.n780 51.2158
R1618 B.n780 B.n50 51.2158
R1619 B.n774 B.n50 51.2158
R1620 B.n774 B.n773 51.2158
R1621 B.n773 B.n772 51.2158
R1622 B.n772 B.n57 51.2158
R1623 B.n766 B.n57 51.2158
R1624 B.n766 B.n765 51.2158
R1625 B.n765 B.n764 51.2158
R1626 B.n764 B.n64 51.2158
R1627 B.n758 B.n757 51.2158
R1628 B.n757 B.n756 51.2158
R1629 B.n756 B.n71 51.2158
R1630 B.n750 B.n71 51.2158
R1631 B.n750 B.n749 51.2158
R1632 B.n749 B.n748 51.2158
R1633 B.n748 B.n78 51.2158
R1634 B.t5 B.n280 48.9563
R1635 B.n821 B.t0 48.9563
R1636 B.n577 B.t7 36.9057
R1637 B.n758 B.t14 36.9057
R1638 B.n644 B.t2 33.893
R1639 B.n804 B.t1 33.893
R1640 B.n613 B.t3 32.3867
R1641 B.n782 B.t4 32.3867
R1642 B.n745 B.n744 32.3127
R1643 B.n739 B.n738 32.3127
R1644 B.n403 B.n353 32.3127
R1645 B.n556 B.n555 32.3127
R1646 B.t3 B.n315 18.8297
R1647 B.t4 B.n43 18.8297
R1648 B B.n832 18.0485
R1649 B.n637 B.t2 17.3233
R1650 B.n32 B.t1 17.3233
R1651 B.t7 B.n339 14.3107
R1652 B.t14 B.n64 14.3107
R1653 B.n744 B.n80 10.6151
R1654 B.n127 B.n80 10.6151
R1655 B.n128 B.n127 10.6151
R1656 B.n131 B.n128 10.6151
R1657 B.n132 B.n131 10.6151
R1658 B.n135 B.n132 10.6151
R1659 B.n136 B.n135 10.6151
R1660 B.n139 B.n136 10.6151
R1661 B.n140 B.n139 10.6151
R1662 B.n143 B.n140 10.6151
R1663 B.n144 B.n143 10.6151
R1664 B.n147 B.n144 10.6151
R1665 B.n148 B.n147 10.6151
R1666 B.n151 B.n148 10.6151
R1667 B.n152 B.n151 10.6151
R1668 B.n155 B.n152 10.6151
R1669 B.n156 B.n155 10.6151
R1670 B.n159 B.n156 10.6151
R1671 B.n160 B.n159 10.6151
R1672 B.n163 B.n160 10.6151
R1673 B.n164 B.n163 10.6151
R1674 B.n167 B.n164 10.6151
R1675 B.n168 B.n167 10.6151
R1676 B.n171 B.n168 10.6151
R1677 B.n172 B.n171 10.6151
R1678 B.n175 B.n172 10.6151
R1679 B.n176 B.n175 10.6151
R1680 B.n179 B.n176 10.6151
R1681 B.n180 B.n179 10.6151
R1682 B.n183 B.n180 10.6151
R1683 B.n184 B.n183 10.6151
R1684 B.n187 B.n184 10.6151
R1685 B.n188 B.n187 10.6151
R1686 B.n192 B.n191 10.6151
R1687 B.n195 B.n192 10.6151
R1688 B.n196 B.n195 10.6151
R1689 B.n199 B.n196 10.6151
R1690 B.n200 B.n199 10.6151
R1691 B.n203 B.n200 10.6151
R1692 B.n204 B.n203 10.6151
R1693 B.n207 B.n204 10.6151
R1694 B.n212 B.n209 10.6151
R1695 B.n213 B.n212 10.6151
R1696 B.n216 B.n213 10.6151
R1697 B.n217 B.n216 10.6151
R1698 B.n220 B.n217 10.6151
R1699 B.n221 B.n220 10.6151
R1700 B.n224 B.n221 10.6151
R1701 B.n225 B.n224 10.6151
R1702 B.n228 B.n225 10.6151
R1703 B.n229 B.n228 10.6151
R1704 B.n232 B.n229 10.6151
R1705 B.n233 B.n232 10.6151
R1706 B.n236 B.n233 10.6151
R1707 B.n237 B.n236 10.6151
R1708 B.n240 B.n237 10.6151
R1709 B.n241 B.n240 10.6151
R1710 B.n244 B.n241 10.6151
R1711 B.n245 B.n244 10.6151
R1712 B.n248 B.n245 10.6151
R1713 B.n249 B.n248 10.6151
R1714 B.n252 B.n249 10.6151
R1715 B.n253 B.n252 10.6151
R1716 B.n256 B.n253 10.6151
R1717 B.n257 B.n256 10.6151
R1718 B.n260 B.n257 10.6151
R1719 B.n261 B.n260 10.6151
R1720 B.n264 B.n261 10.6151
R1721 B.n265 B.n264 10.6151
R1722 B.n268 B.n265 10.6151
R1723 B.n269 B.n268 10.6151
R1724 B.n272 B.n269 10.6151
R1725 B.n273 B.n272 10.6151
R1726 B.n739 B.n273 10.6151
R1727 B.n561 B.n353 10.6151
R1728 B.n562 B.n561 10.6151
R1729 B.n563 B.n562 10.6151
R1730 B.n563 B.n345 10.6151
R1731 B.n573 B.n345 10.6151
R1732 B.n574 B.n573 10.6151
R1733 B.n575 B.n574 10.6151
R1734 B.n575 B.n337 10.6151
R1735 B.n585 B.n337 10.6151
R1736 B.n586 B.n585 10.6151
R1737 B.n587 B.n586 10.6151
R1738 B.n587 B.n329 10.6151
R1739 B.n597 B.n329 10.6151
R1740 B.n598 B.n597 10.6151
R1741 B.n599 B.n598 10.6151
R1742 B.n599 B.n321 10.6151
R1743 B.n609 B.n321 10.6151
R1744 B.n610 B.n609 10.6151
R1745 B.n611 B.n610 10.6151
R1746 B.n611 B.n313 10.6151
R1747 B.n621 B.n313 10.6151
R1748 B.n622 B.n621 10.6151
R1749 B.n623 B.n622 10.6151
R1750 B.n623 B.n305 10.6151
R1751 B.n633 B.n305 10.6151
R1752 B.n634 B.n633 10.6151
R1753 B.n635 B.n634 10.6151
R1754 B.n635 B.n298 10.6151
R1755 B.n646 B.n298 10.6151
R1756 B.n647 B.n646 10.6151
R1757 B.n648 B.n647 10.6151
R1758 B.n648 B.n290 10.6151
R1759 B.n658 B.n290 10.6151
R1760 B.n659 B.n658 10.6151
R1761 B.n660 B.n659 10.6151
R1762 B.n660 B.n282 10.6151
R1763 B.n670 B.n282 10.6151
R1764 B.n671 B.n670 10.6151
R1765 B.n673 B.n671 10.6151
R1766 B.n673 B.n672 10.6151
R1767 B.n672 B.n274 10.6151
R1768 B.n684 B.n274 10.6151
R1769 B.n685 B.n684 10.6151
R1770 B.n686 B.n685 10.6151
R1771 B.n687 B.n686 10.6151
R1772 B.n689 B.n687 10.6151
R1773 B.n690 B.n689 10.6151
R1774 B.n691 B.n690 10.6151
R1775 B.n692 B.n691 10.6151
R1776 B.n694 B.n692 10.6151
R1777 B.n695 B.n694 10.6151
R1778 B.n696 B.n695 10.6151
R1779 B.n697 B.n696 10.6151
R1780 B.n699 B.n697 10.6151
R1781 B.n700 B.n699 10.6151
R1782 B.n701 B.n700 10.6151
R1783 B.n702 B.n701 10.6151
R1784 B.n704 B.n702 10.6151
R1785 B.n705 B.n704 10.6151
R1786 B.n706 B.n705 10.6151
R1787 B.n707 B.n706 10.6151
R1788 B.n709 B.n707 10.6151
R1789 B.n710 B.n709 10.6151
R1790 B.n711 B.n710 10.6151
R1791 B.n712 B.n711 10.6151
R1792 B.n714 B.n712 10.6151
R1793 B.n715 B.n714 10.6151
R1794 B.n716 B.n715 10.6151
R1795 B.n717 B.n716 10.6151
R1796 B.n719 B.n717 10.6151
R1797 B.n720 B.n719 10.6151
R1798 B.n721 B.n720 10.6151
R1799 B.n722 B.n721 10.6151
R1800 B.n724 B.n722 10.6151
R1801 B.n725 B.n724 10.6151
R1802 B.n726 B.n725 10.6151
R1803 B.n727 B.n726 10.6151
R1804 B.n729 B.n727 10.6151
R1805 B.n730 B.n729 10.6151
R1806 B.n731 B.n730 10.6151
R1807 B.n732 B.n731 10.6151
R1808 B.n734 B.n732 10.6151
R1809 B.n735 B.n734 10.6151
R1810 B.n736 B.n735 10.6151
R1811 B.n737 B.n736 10.6151
R1812 B.n738 B.n737 10.6151
R1813 B.n555 B.n357 10.6151
R1814 B.n550 B.n357 10.6151
R1815 B.n550 B.n549 10.6151
R1816 B.n549 B.n548 10.6151
R1817 B.n548 B.n545 10.6151
R1818 B.n545 B.n544 10.6151
R1819 B.n544 B.n541 10.6151
R1820 B.n541 B.n540 10.6151
R1821 B.n540 B.n537 10.6151
R1822 B.n537 B.n536 10.6151
R1823 B.n536 B.n533 10.6151
R1824 B.n533 B.n532 10.6151
R1825 B.n532 B.n529 10.6151
R1826 B.n529 B.n528 10.6151
R1827 B.n528 B.n525 10.6151
R1828 B.n525 B.n524 10.6151
R1829 B.n524 B.n521 10.6151
R1830 B.n521 B.n520 10.6151
R1831 B.n520 B.n517 10.6151
R1832 B.n517 B.n516 10.6151
R1833 B.n516 B.n513 10.6151
R1834 B.n513 B.n512 10.6151
R1835 B.n512 B.n509 10.6151
R1836 B.n509 B.n508 10.6151
R1837 B.n508 B.n505 10.6151
R1838 B.n505 B.n504 10.6151
R1839 B.n504 B.n501 10.6151
R1840 B.n501 B.n500 10.6151
R1841 B.n500 B.n497 10.6151
R1842 B.n497 B.n496 10.6151
R1843 B.n496 B.n493 10.6151
R1844 B.n493 B.n492 10.6151
R1845 B.n492 B.n489 10.6151
R1846 B.n487 B.n484 10.6151
R1847 B.n484 B.n483 10.6151
R1848 B.n483 B.n480 10.6151
R1849 B.n480 B.n479 10.6151
R1850 B.n479 B.n476 10.6151
R1851 B.n476 B.n475 10.6151
R1852 B.n475 B.n472 10.6151
R1853 B.n472 B.n471 10.6151
R1854 B.n468 B.n467 10.6151
R1855 B.n467 B.n464 10.6151
R1856 B.n464 B.n463 10.6151
R1857 B.n463 B.n460 10.6151
R1858 B.n460 B.n459 10.6151
R1859 B.n459 B.n456 10.6151
R1860 B.n456 B.n455 10.6151
R1861 B.n455 B.n452 10.6151
R1862 B.n452 B.n451 10.6151
R1863 B.n451 B.n448 10.6151
R1864 B.n448 B.n447 10.6151
R1865 B.n447 B.n444 10.6151
R1866 B.n444 B.n443 10.6151
R1867 B.n443 B.n440 10.6151
R1868 B.n440 B.n439 10.6151
R1869 B.n439 B.n436 10.6151
R1870 B.n436 B.n435 10.6151
R1871 B.n435 B.n432 10.6151
R1872 B.n432 B.n431 10.6151
R1873 B.n431 B.n428 10.6151
R1874 B.n428 B.n427 10.6151
R1875 B.n427 B.n424 10.6151
R1876 B.n424 B.n423 10.6151
R1877 B.n423 B.n420 10.6151
R1878 B.n420 B.n419 10.6151
R1879 B.n419 B.n416 10.6151
R1880 B.n416 B.n415 10.6151
R1881 B.n415 B.n412 10.6151
R1882 B.n412 B.n411 10.6151
R1883 B.n411 B.n408 10.6151
R1884 B.n408 B.n407 10.6151
R1885 B.n407 B.n404 10.6151
R1886 B.n404 B.n403 10.6151
R1887 B.n557 B.n556 10.6151
R1888 B.n557 B.n349 10.6151
R1889 B.n567 B.n349 10.6151
R1890 B.n568 B.n567 10.6151
R1891 B.n569 B.n568 10.6151
R1892 B.n569 B.n341 10.6151
R1893 B.n579 B.n341 10.6151
R1894 B.n580 B.n579 10.6151
R1895 B.n581 B.n580 10.6151
R1896 B.n581 B.n333 10.6151
R1897 B.n591 B.n333 10.6151
R1898 B.n592 B.n591 10.6151
R1899 B.n593 B.n592 10.6151
R1900 B.n593 B.n325 10.6151
R1901 B.n603 B.n325 10.6151
R1902 B.n604 B.n603 10.6151
R1903 B.n605 B.n604 10.6151
R1904 B.n605 B.n317 10.6151
R1905 B.n615 B.n317 10.6151
R1906 B.n616 B.n615 10.6151
R1907 B.n617 B.n616 10.6151
R1908 B.n617 B.n309 10.6151
R1909 B.n627 B.n309 10.6151
R1910 B.n628 B.n627 10.6151
R1911 B.n629 B.n628 10.6151
R1912 B.n629 B.n301 10.6151
R1913 B.n640 B.n301 10.6151
R1914 B.n641 B.n640 10.6151
R1915 B.n642 B.n641 10.6151
R1916 B.n642 B.n294 10.6151
R1917 B.n652 B.n294 10.6151
R1918 B.n653 B.n652 10.6151
R1919 B.n654 B.n653 10.6151
R1920 B.n654 B.n286 10.6151
R1921 B.n664 B.n286 10.6151
R1922 B.n665 B.n664 10.6151
R1923 B.n666 B.n665 10.6151
R1924 B.n666 B.n278 10.6151
R1925 B.n677 B.n278 10.6151
R1926 B.n678 B.n677 10.6151
R1927 B.n679 B.n678 10.6151
R1928 B.n679 B.n0 10.6151
R1929 B.n826 B.n1 10.6151
R1930 B.n826 B.n825 10.6151
R1931 B.n825 B.n824 10.6151
R1932 B.n824 B.n10 10.6151
R1933 B.n818 B.n10 10.6151
R1934 B.n818 B.n817 10.6151
R1935 B.n817 B.n816 10.6151
R1936 B.n816 B.n17 10.6151
R1937 B.n810 B.n17 10.6151
R1938 B.n810 B.n809 10.6151
R1939 B.n809 B.n808 10.6151
R1940 B.n808 B.n24 10.6151
R1941 B.n802 B.n24 10.6151
R1942 B.n802 B.n801 10.6151
R1943 B.n801 B.n800 10.6151
R1944 B.n800 B.n30 10.6151
R1945 B.n794 B.n30 10.6151
R1946 B.n794 B.n793 10.6151
R1947 B.n793 B.n792 10.6151
R1948 B.n792 B.n38 10.6151
R1949 B.n786 B.n38 10.6151
R1950 B.n786 B.n785 10.6151
R1951 B.n785 B.n784 10.6151
R1952 B.n784 B.n45 10.6151
R1953 B.n778 B.n45 10.6151
R1954 B.n778 B.n777 10.6151
R1955 B.n777 B.n776 10.6151
R1956 B.n776 B.n52 10.6151
R1957 B.n770 B.n52 10.6151
R1958 B.n770 B.n769 10.6151
R1959 B.n769 B.n768 10.6151
R1960 B.n768 B.n59 10.6151
R1961 B.n762 B.n59 10.6151
R1962 B.n762 B.n761 10.6151
R1963 B.n761 B.n760 10.6151
R1964 B.n760 B.n66 10.6151
R1965 B.n754 B.n66 10.6151
R1966 B.n754 B.n753 10.6151
R1967 B.n753 B.n752 10.6151
R1968 B.n752 B.n73 10.6151
R1969 B.n746 B.n73 10.6151
R1970 B.n746 B.n745 10.6151
R1971 B.n191 B.n125 6.5566
R1972 B.n208 B.n207 6.5566
R1973 B.n488 B.n487 6.5566
R1974 B.n471 B.n401 6.5566
R1975 B.n188 B.n125 4.05904
R1976 B.n209 B.n208 4.05904
R1977 B.n489 B.n488 4.05904
R1978 B.n468 B.n401 4.05904
R1979 B.n832 B.n0 2.81026
R1980 B.n832 B.n1 2.81026
R1981 B.n668 B.t5 2.26
R1982 B.t0 B.n820 2.26
R1983 VN.n29 VN.n16 161.3
R1984 VN.n28 VN.n27 161.3
R1985 VN.n26 VN.n17 161.3
R1986 VN.n25 VN.n24 161.3
R1987 VN.n23 VN.n18 161.3
R1988 VN.n22 VN.n21 161.3
R1989 VN.n13 VN.n0 161.3
R1990 VN.n12 VN.n11 161.3
R1991 VN.n10 VN.n1 161.3
R1992 VN.n9 VN.n8 161.3
R1993 VN.n7 VN.n2 161.3
R1994 VN.n6 VN.n5 161.3
R1995 VN.n4 VN.t3 119.18
R1996 VN.n20 VN.t5 119.18
R1997 VN.n15 VN.n14 100.481
R1998 VN.n31 VN.n30 100.481
R1999 VN.n3 VN.t4 85.4959
R2000 VN.n14 VN.t2 85.4959
R2001 VN.n19 VN.t1 85.4959
R2002 VN.n30 VN.t0 85.4959
R2003 VN.n4 VN.n3 60.2369
R2004 VN.n20 VN.n19 60.2369
R2005 VN.n8 VN.n1 56.5193
R2006 VN.n24 VN.n17 56.5193
R2007 VN VN.n31 47.0815
R2008 VN.n7 VN.n6 24.4675
R2009 VN.n8 VN.n7 24.4675
R2010 VN.n12 VN.n1 24.4675
R2011 VN.n13 VN.n12 24.4675
R2012 VN.n24 VN.n23 24.4675
R2013 VN.n23 VN.n22 24.4675
R2014 VN.n29 VN.n28 24.4675
R2015 VN.n28 VN.n17 24.4675
R2016 VN.n6 VN.n3 12.234
R2017 VN.n22 VN.n19 12.234
R2018 VN.n14 VN.n13 10.2766
R2019 VN.n30 VN.n29 10.2766
R2020 VN.n21 VN.n20 6.83261
R2021 VN.n5 VN.n4 6.83261
R2022 VN.n31 VN.n16 0.278367
R2023 VN.n15 VN.n0 0.278367
R2024 VN.n27 VN.n16 0.189894
R2025 VN.n27 VN.n26 0.189894
R2026 VN.n26 VN.n25 0.189894
R2027 VN.n25 VN.n18 0.189894
R2028 VN.n21 VN.n18 0.189894
R2029 VN.n5 VN.n2 0.189894
R2030 VN.n9 VN.n2 0.189894
R2031 VN.n10 VN.n9 0.189894
R2032 VN.n11 VN.n10 0.189894
R2033 VN.n11 VN.n0 0.189894
R2034 VN VN.n15 0.153454
R2035 VDD2.n95 VDD2.n51 289.615
R2036 VDD2.n44 VDD2.n0 289.615
R2037 VDD2.n96 VDD2.n95 185
R2038 VDD2.n94 VDD2.n93 185
R2039 VDD2.n55 VDD2.n54 185
R2040 VDD2.n59 VDD2.n57 185
R2041 VDD2.n88 VDD2.n87 185
R2042 VDD2.n86 VDD2.n85 185
R2043 VDD2.n61 VDD2.n60 185
R2044 VDD2.n80 VDD2.n79 185
R2045 VDD2.n78 VDD2.n77 185
R2046 VDD2.n65 VDD2.n64 185
R2047 VDD2.n72 VDD2.n71 185
R2048 VDD2.n70 VDD2.n69 185
R2049 VDD2.n17 VDD2.n16 185
R2050 VDD2.n19 VDD2.n18 185
R2051 VDD2.n12 VDD2.n11 185
R2052 VDD2.n25 VDD2.n24 185
R2053 VDD2.n27 VDD2.n26 185
R2054 VDD2.n8 VDD2.n7 185
R2055 VDD2.n34 VDD2.n33 185
R2056 VDD2.n35 VDD2.n6 185
R2057 VDD2.n37 VDD2.n36 185
R2058 VDD2.n4 VDD2.n3 185
R2059 VDD2.n43 VDD2.n42 185
R2060 VDD2.n45 VDD2.n44 185
R2061 VDD2.n68 VDD2.t5 149.524
R2062 VDD2.n15 VDD2.t2 149.524
R2063 VDD2.n95 VDD2.n94 104.615
R2064 VDD2.n94 VDD2.n54 104.615
R2065 VDD2.n59 VDD2.n54 104.615
R2066 VDD2.n87 VDD2.n59 104.615
R2067 VDD2.n87 VDD2.n86 104.615
R2068 VDD2.n86 VDD2.n60 104.615
R2069 VDD2.n79 VDD2.n60 104.615
R2070 VDD2.n79 VDD2.n78 104.615
R2071 VDD2.n78 VDD2.n64 104.615
R2072 VDD2.n71 VDD2.n64 104.615
R2073 VDD2.n71 VDD2.n70 104.615
R2074 VDD2.n18 VDD2.n17 104.615
R2075 VDD2.n18 VDD2.n11 104.615
R2076 VDD2.n25 VDD2.n11 104.615
R2077 VDD2.n26 VDD2.n25 104.615
R2078 VDD2.n26 VDD2.n7 104.615
R2079 VDD2.n34 VDD2.n7 104.615
R2080 VDD2.n35 VDD2.n34 104.615
R2081 VDD2.n36 VDD2.n35 104.615
R2082 VDD2.n36 VDD2.n3 104.615
R2083 VDD2.n43 VDD2.n3 104.615
R2084 VDD2.n44 VDD2.n43 104.615
R2085 VDD2.n50 VDD2.n49 65.3299
R2086 VDD2 VDD2.n101 65.3271
R2087 VDD2.n50 VDD2.n48 52.468
R2088 VDD2.n70 VDD2.t5 52.3082
R2089 VDD2.n17 VDD2.t2 52.3082
R2090 VDD2.n100 VDD2.n99 50.6096
R2091 VDD2.n100 VDD2.n50 40.0515
R2092 VDD2.n57 VDD2.n55 13.1884
R2093 VDD2.n37 VDD2.n4 13.1884
R2094 VDD2.n93 VDD2.n92 12.8005
R2095 VDD2.n89 VDD2.n88 12.8005
R2096 VDD2.n38 VDD2.n6 12.8005
R2097 VDD2.n42 VDD2.n41 12.8005
R2098 VDD2.n96 VDD2.n53 12.0247
R2099 VDD2.n85 VDD2.n58 12.0247
R2100 VDD2.n33 VDD2.n32 12.0247
R2101 VDD2.n45 VDD2.n2 12.0247
R2102 VDD2.n97 VDD2.n51 11.249
R2103 VDD2.n84 VDD2.n61 11.249
R2104 VDD2.n31 VDD2.n8 11.249
R2105 VDD2.n46 VDD2.n0 11.249
R2106 VDD2.n81 VDD2.n80 10.4732
R2107 VDD2.n28 VDD2.n27 10.4732
R2108 VDD2.n69 VDD2.n68 10.2747
R2109 VDD2.n16 VDD2.n15 10.2747
R2110 VDD2.n77 VDD2.n63 9.69747
R2111 VDD2.n24 VDD2.n10 9.69747
R2112 VDD2.n99 VDD2.n98 9.45567
R2113 VDD2.n48 VDD2.n47 9.45567
R2114 VDD2.n67 VDD2.n66 9.3005
R2115 VDD2.n74 VDD2.n73 9.3005
R2116 VDD2.n76 VDD2.n75 9.3005
R2117 VDD2.n63 VDD2.n62 9.3005
R2118 VDD2.n82 VDD2.n81 9.3005
R2119 VDD2.n84 VDD2.n83 9.3005
R2120 VDD2.n58 VDD2.n56 9.3005
R2121 VDD2.n90 VDD2.n89 9.3005
R2122 VDD2.n98 VDD2.n97 9.3005
R2123 VDD2.n53 VDD2.n52 9.3005
R2124 VDD2.n92 VDD2.n91 9.3005
R2125 VDD2.n47 VDD2.n46 9.3005
R2126 VDD2.n2 VDD2.n1 9.3005
R2127 VDD2.n41 VDD2.n40 9.3005
R2128 VDD2.n14 VDD2.n13 9.3005
R2129 VDD2.n21 VDD2.n20 9.3005
R2130 VDD2.n23 VDD2.n22 9.3005
R2131 VDD2.n10 VDD2.n9 9.3005
R2132 VDD2.n29 VDD2.n28 9.3005
R2133 VDD2.n31 VDD2.n30 9.3005
R2134 VDD2.n32 VDD2.n5 9.3005
R2135 VDD2.n39 VDD2.n38 9.3005
R2136 VDD2.n76 VDD2.n65 8.92171
R2137 VDD2.n23 VDD2.n12 8.92171
R2138 VDD2.n73 VDD2.n72 8.14595
R2139 VDD2.n20 VDD2.n19 8.14595
R2140 VDD2.n69 VDD2.n67 7.3702
R2141 VDD2.n16 VDD2.n14 7.3702
R2142 VDD2.n72 VDD2.n67 5.81868
R2143 VDD2.n19 VDD2.n14 5.81868
R2144 VDD2.n73 VDD2.n65 5.04292
R2145 VDD2.n20 VDD2.n12 5.04292
R2146 VDD2.n77 VDD2.n76 4.26717
R2147 VDD2.n24 VDD2.n23 4.26717
R2148 VDD2.n80 VDD2.n63 3.49141
R2149 VDD2.n27 VDD2.n10 3.49141
R2150 VDD2.n68 VDD2.n66 2.84303
R2151 VDD2.n15 VDD2.n13 2.84303
R2152 VDD2.n99 VDD2.n51 2.71565
R2153 VDD2.n81 VDD2.n61 2.71565
R2154 VDD2.n28 VDD2.n8 2.71565
R2155 VDD2.n48 VDD2.n0 2.71565
R2156 VDD2.n101 VDD2.t4 2.12269
R2157 VDD2.n101 VDD2.t0 2.12269
R2158 VDD2.n49 VDD2.t1 2.12269
R2159 VDD2.n49 VDD2.t3 2.12269
R2160 VDD2 VDD2.n100 1.97248
R2161 VDD2.n97 VDD2.n96 1.93989
R2162 VDD2.n85 VDD2.n84 1.93989
R2163 VDD2.n33 VDD2.n31 1.93989
R2164 VDD2.n46 VDD2.n45 1.93989
R2165 VDD2.n93 VDD2.n53 1.16414
R2166 VDD2.n88 VDD2.n58 1.16414
R2167 VDD2.n32 VDD2.n6 1.16414
R2168 VDD2.n42 VDD2.n2 1.16414
R2169 VDD2.n92 VDD2.n55 0.388379
R2170 VDD2.n89 VDD2.n57 0.388379
R2171 VDD2.n38 VDD2.n37 0.388379
R2172 VDD2.n41 VDD2.n4 0.388379
R2173 VDD2.n98 VDD2.n52 0.155672
R2174 VDD2.n91 VDD2.n52 0.155672
R2175 VDD2.n91 VDD2.n90 0.155672
R2176 VDD2.n90 VDD2.n56 0.155672
R2177 VDD2.n83 VDD2.n56 0.155672
R2178 VDD2.n83 VDD2.n82 0.155672
R2179 VDD2.n82 VDD2.n62 0.155672
R2180 VDD2.n75 VDD2.n62 0.155672
R2181 VDD2.n75 VDD2.n74 0.155672
R2182 VDD2.n74 VDD2.n66 0.155672
R2183 VDD2.n21 VDD2.n13 0.155672
R2184 VDD2.n22 VDD2.n21 0.155672
R2185 VDD2.n22 VDD2.n9 0.155672
R2186 VDD2.n29 VDD2.n9 0.155672
R2187 VDD2.n30 VDD2.n29 0.155672
R2188 VDD2.n30 VDD2.n5 0.155672
R2189 VDD2.n39 VDD2.n5 0.155672
R2190 VDD2.n40 VDD2.n39 0.155672
R2191 VDD2.n40 VDD2.n1 0.155672
R2192 VDD2.n47 VDD2.n1 0.155672
C0 VDD2 VP 0.460734f
C1 VDD2 VN 5.32141f
C2 VDD1 VTAIL 6.77092f
C3 VP VN 6.45954f
C4 VDD2 VDD1 1.41894f
C5 VDD2 VTAIL 6.8226f
C6 VDD1 VP 5.62857f
C7 VDD1 VN 0.150862f
C8 VTAIL VP 5.61853f
C9 VTAIL VN 5.60428f
C10 VDD2 B 5.533466f
C11 VDD1 B 5.668161f
C12 VTAIL B 6.768637f
C13 VN B 12.749929f
C14 VP B 11.415327f
C15 VDD2.n0 B 0.029143f
C16 VDD2.n1 B 0.021454f
C17 VDD2.n2 B 0.011529f
C18 VDD2.n3 B 0.027249f
C19 VDD2.n4 B 0.011868f
C20 VDD2.n5 B 0.021454f
C21 VDD2.n6 B 0.012207f
C22 VDD2.n7 B 0.027249f
C23 VDD2.n8 B 0.012207f
C24 VDD2.n9 B 0.021454f
C25 VDD2.n10 B 0.011529f
C26 VDD2.n11 B 0.027249f
C27 VDD2.n12 B 0.012207f
C28 VDD2.n13 B 0.827534f
C29 VDD2.n14 B 0.011529f
C30 VDD2.t2 B 0.045717f
C31 VDD2.n15 B 0.132697f
C32 VDD2.n16 B 0.019263f
C33 VDD2.n17 B 0.020437f
C34 VDD2.n18 B 0.027249f
C35 VDD2.n19 B 0.012207f
C36 VDD2.n20 B 0.011529f
C37 VDD2.n21 B 0.021454f
C38 VDD2.n22 B 0.021454f
C39 VDD2.n23 B 0.011529f
C40 VDD2.n24 B 0.012207f
C41 VDD2.n25 B 0.027249f
C42 VDD2.n26 B 0.027249f
C43 VDD2.n27 B 0.012207f
C44 VDD2.n28 B 0.011529f
C45 VDD2.n29 B 0.021454f
C46 VDD2.n30 B 0.021454f
C47 VDD2.n31 B 0.011529f
C48 VDD2.n32 B 0.011529f
C49 VDD2.n33 B 0.012207f
C50 VDD2.n34 B 0.027249f
C51 VDD2.n35 B 0.027249f
C52 VDD2.n36 B 0.027249f
C53 VDD2.n37 B 0.011868f
C54 VDD2.n38 B 0.011529f
C55 VDD2.n39 B 0.021454f
C56 VDD2.n40 B 0.021454f
C57 VDD2.n41 B 0.011529f
C58 VDD2.n42 B 0.012207f
C59 VDD2.n43 B 0.027249f
C60 VDD2.n44 B 0.057199f
C61 VDD2.n45 B 0.012207f
C62 VDD2.n46 B 0.011529f
C63 VDD2.n47 B 0.052228f
C64 VDD2.n48 B 0.052771f
C65 VDD2.t1 B 0.158179f
C66 VDD2.t3 B 0.158179f
C67 VDD2.n49 B 1.39052f
C68 VDD2.n50 B 2.167f
C69 VDD2.n51 B 0.029143f
C70 VDD2.n52 B 0.021454f
C71 VDD2.n53 B 0.011529f
C72 VDD2.n54 B 0.027249f
C73 VDD2.n55 B 0.011868f
C74 VDD2.n56 B 0.021454f
C75 VDD2.n57 B 0.011868f
C76 VDD2.n58 B 0.011529f
C77 VDD2.n59 B 0.027249f
C78 VDD2.n60 B 0.027249f
C79 VDD2.n61 B 0.012207f
C80 VDD2.n62 B 0.021454f
C81 VDD2.n63 B 0.011529f
C82 VDD2.n64 B 0.027249f
C83 VDD2.n65 B 0.012207f
C84 VDD2.n66 B 0.827534f
C85 VDD2.n67 B 0.011529f
C86 VDD2.t5 B 0.045717f
C87 VDD2.n68 B 0.132697f
C88 VDD2.n69 B 0.019263f
C89 VDD2.n70 B 0.020437f
C90 VDD2.n71 B 0.027249f
C91 VDD2.n72 B 0.012207f
C92 VDD2.n73 B 0.011529f
C93 VDD2.n74 B 0.021454f
C94 VDD2.n75 B 0.021454f
C95 VDD2.n76 B 0.011529f
C96 VDD2.n77 B 0.012207f
C97 VDD2.n78 B 0.027249f
C98 VDD2.n79 B 0.027249f
C99 VDD2.n80 B 0.012207f
C100 VDD2.n81 B 0.011529f
C101 VDD2.n82 B 0.021454f
C102 VDD2.n83 B 0.021454f
C103 VDD2.n84 B 0.011529f
C104 VDD2.n85 B 0.012207f
C105 VDD2.n86 B 0.027249f
C106 VDD2.n87 B 0.027249f
C107 VDD2.n88 B 0.012207f
C108 VDD2.n89 B 0.011529f
C109 VDD2.n90 B 0.021454f
C110 VDD2.n91 B 0.021454f
C111 VDD2.n92 B 0.011529f
C112 VDD2.n93 B 0.012207f
C113 VDD2.n94 B 0.027249f
C114 VDD2.n95 B 0.057199f
C115 VDD2.n96 B 0.012207f
C116 VDD2.n97 B 0.011529f
C117 VDD2.n98 B 0.052228f
C118 VDD2.n99 B 0.046694f
C119 VDD2.n100 B 2.02867f
C120 VDD2.t4 B 0.158179f
C121 VDD2.t0 B 0.158179f
C122 VDD2.n101 B 1.39049f
C123 VN.n0 B 0.031584f
C124 VN.t2 B 1.58856f
C125 VN.n1 B 0.036307f
C126 VN.n2 B 0.023957f
C127 VN.t4 B 1.58856f
C128 VN.n3 B 0.6407f
C129 VN.t3 B 1.7924f
C130 VN.n4 B 0.61827f
C131 VN.n5 B 0.232299f
C132 VN.n6 B 0.033627f
C133 VN.n7 B 0.044649f
C134 VN.n8 B 0.033637f
C135 VN.n9 B 0.023957f
C136 VN.n10 B 0.023957f
C137 VN.n11 B 0.023957f
C138 VN.n12 B 0.044649f
C139 VN.n13 B 0.031864f
C140 VN.n14 B 0.652948f
C141 VN.n15 B 0.039016f
C142 VN.n16 B 0.031584f
C143 VN.t0 B 1.58856f
C144 VN.n17 B 0.036307f
C145 VN.n18 B 0.023957f
C146 VN.t1 B 1.58856f
C147 VN.n19 B 0.6407f
C148 VN.t5 B 1.7924f
C149 VN.n20 B 0.61827f
C150 VN.n21 B 0.232299f
C151 VN.n22 B 0.033627f
C152 VN.n23 B 0.044649f
C153 VN.n24 B 0.033637f
C154 VN.n25 B 0.023957f
C155 VN.n26 B 0.023957f
C156 VN.n27 B 0.023957f
C157 VN.n28 B 0.044649f
C158 VN.n29 B 0.031864f
C159 VN.n30 B 0.652948f
C160 VN.n31 B 1.2211f
C161 VTAIL.t0 B 0.181803f
C162 VTAIL.t1 B 0.181803f
C163 VTAIL.n0 B 1.52685f
C164 VTAIL.n1 B 0.426274f
C165 VTAIL.n2 B 0.033495f
C166 VTAIL.n3 B 0.024659f
C167 VTAIL.n4 B 0.01325f
C168 VTAIL.n5 B 0.031319f
C169 VTAIL.n6 B 0.01364f
C170 VTAIL.n7 B 0.024659f
C171 VTAIL.n8 B 0.01403f
C172 VTAIL.n9 B 0.031319f
C173 VTAIL.n10 B 0.01403f
C174 VTAIL.n11 B 0.024659f
C175 VTAIL.n12 B 0.01325f
C176 VTAIL.n13 B 0.031319f
C177 VTAIL.n14 B 0.01403f
C178 VTAIL.n15 B 0.951127f
C179 VTAIL.n16 B 0.01325f
C180 VTAIL.t7 B 0.052545f
C181 VTAIL.n17 B 0.152516f
C182 VTAIL.n18 B 0.02214f
C183 VTAIL.n19 B 0.023489f
C184 VTAIL.n20 B 0.031319f
C185 VTAIL.n21 B 0.01403f
C186 VTAIL.n22 B 0.01325f
C187 VTAIL.n23 B 0.024659f
C188 VTAIL.n24 B 0.024659f
C189 VTAIL.n25 B 0.01325f
C190 VTAIL.n26 B 0.01403f
C191 VTAIL.n27 B 0.031319f
C192 VTAIL.n28 B 0.031319f
C193 VTAIL.n29 B 0.01403f
C194 VTAIL.n30 B 0.01325f
C195 VTAIL.n31 B 0.024659f
C196 VTAIL.n32 B 0.024659f
C197 VTAIL.n33 B 0.01325f
C198 VTAIL.n34 B 0.01325f
C199 VTAIL.n35 B 0.01403f
C200 VTAIL.n36 B 0.031319f
C201 VTAIL.n37 B 0.031319f
C202 VTAIL.n38 B 0.031319f
C203 VTAIL.n39 B 0.01364f
C204 VTAIL.n40 B 0.01325f
C205 VTAIL.n41 B 0.024659f
C206 VTAIL.n42 B 0.024659f
C207 VTAIL.n43 B 0.01325f
C208 VTAIL.n44 B 0.01403f
C209 VTAIL.n45 B 0.031319f
C210 VTAIL.n46 B 0.065741f
C211 VTAIL.n47 B 0.01403f
C212 VTAIL.n48 B 0.01325f
C213 VTAIL.n49 B 0.060029f
C214 VTAIL.n50 B 0.036664f
C215 VTAIL.n51 B 0.364225f
C216 VTAIL.t6 B 0.181803f
C217 VTAIL.t11 B 0.181803f
C218 VTAIL.n52 B 1.52685f
C219 VTAIL.n53 B 1.81452f
C220 VTAIL.t3 B 0.181803f
C221 VTAIL.t2 B 0.181803f
C222 VTAIL.n54 B 1.52686f
C223 VTAIL.n55 B 1.81451f
C224 VTAIL.n56 B 0.033495f
C225 VTAIL.n57 B 0.024659f
C226 VTAIL.n58 B 0.01325f
C227 VTAIL.n59 B 0.031319f
C228 VTAIL.n60 B 0.01364f
C229 VTAIL.n61 B 0.024659f
C230 VTAIL.n62 B 0.01364f
C231 VTAIL.n63 B 0.01325f
C232 VTAIL.n64 B 0.031319f
C233 VTAIL.n65 B 0.031319f
C234 VTAIL.n66 B 0.01403f
C235 VTAIL.n67 B 0.024659f
C236 VTAIL.n68 B 0.01325f
C237 VTAIL.n69 B 0.031319f
C238 VTAIL.n70 B 0.01403f
C239 VTAIL.n71 B 0.951127f
C240 VTAIL.n72 B 0.01325f
C241 VTAIL.t5 B 0.052545f
C242 VTAIL.n73 B 0.152516f
C243 VTAIL.n74 B 0.02214f
C244 VTAIL.n75 B 0.023489f
C245 VTAIL.n76 B 0.031319f
C246 VTAIL.n77 B 0.01403f
C247 VTAIL.n78 B 0.01325f
C248 VTAIL.n79 B 0.024659f
C249 VTAIL.n80 B 0.024659f
C250 VTAIL.n81 B 0.01325f
C251 VTAIL.n82 B 0.01403f
C252 VTAIL.n83 B 0.031319f
C253 VTAIL.n84 B 0.031319f
C254 VTAIL.n85 B 0.01403f
C255 VTAIL.n86 B 0.01325f
C256 VTAIL.n87 B 0.024659f
C257 VTAIL.n88 B 0.024659f
C258 VTAIL.n89 B 0.01325f
C259 VTAIL.n90 B 0.01403f
C260 VTAIL.n91 B 0.031319f
C261 VTAIL.n92 B 0.031319f
C262 VTAIL.n93 B 0.01403f
C263 VTAIL.n94 B 0.01325f
C264 VTAIL.n95 B 0.024659f
C265 VTAIL.n96 B 0.024659f
C266 VTAIL.n97 B 0.01325f
C267 VTAIL.n98 B 0.01403f
C268 VTAIL.n99 B 0.031319f
C269 VTAIL.n100 B 0.065741f
C270 VTAIL.n101 B 0.01403f
C271 VTAIL.n102 B 0.01325f
C272 VTAIL.n103 B 0.060029f
C273 VTAIL.n104 B 0.036664f
C274 VTAIL.n105 B 0.364225f
C275 VTAIL.t8 B 0.181803f
C276 VTAIL.t9 B 0.181803f
C277 VTAIL.n106 B 1.52686f
C278 VTAIL.n107 B 0.573702f
C279 VTAIL.n108 B 0.033495f
C280 VTAIL.n109 B 0.024659f
C281 VTAIL.n110 B 0.01325f
C282 VTAIL.n111 B 0.031319f
C283 VTAIL.n112 B 0.01364f
C284 VTAIL.n113 B 0.024659f
C285 VTAIL.n114 B 0.01364f
C286 VTAIL.n115 B 0.01325f
C287 VTAIL.n116 B 0.031319f
C288 VTAIL.n117 B 0.031319f
C289 VTAIL.n118 B 0.01403f
C290 VTAIL.n119 B 0.024659f
C291 VTAIL.n120 B 0.01325f
C292 VTAIL.n121 B 0.031319f
C293 VTAIL.n122 B 0.01403f
C294 VTAIL.n123 B 0.951127f
C295 VTAIL.n124 B 0.01325f
C296 VTAIL.t10 B 0.052545f
C297 VTAIL.n125 B 0.152516f
C298 VTAIL.n126 B 0.02214f
C299 VTAIL.n127 B 0.023489f
C300 VTAIL.n128 B 0.031319f
C301 VTAIL.n129 B 0.01403f
C302 VTAIL.n130 B 0.01325f
C303 VTAIL.n131 B 0.024659f
C304 VTAIL.n132 B 0.024659f
C305 VTAIL.n133 B 0.01325f
C306 VTAIL.n134 B 0.01403f
C307 VTAIL.n135 B 0.031319f
C308 VTAIL.n136 B 0.031319f
C309 VTAIL.n137 B 0.01403f
C310 VTAIL.n138 B 0.01325f
C311 VTAIL.n139 B 0.024659f
C312 VTAIL.n140 B 0.024659f
C313 VTAIL.n141 B 0.01325f
C314 VTAIL.n142 B 0.01403f
C315 VTAIL.n143 B 0.031319f
C316 VTAIL.n144 B 0.031319f
C317 VTAIL.n145 B 0.01403f
C318 VTAIL.n146 B 0.01325f
C319 VTAIL.n147 B 0.024659f
C320 VTAIL.n148 B 0.024659f
C321 VTAIL.n149 B 0.01325f
C322 VTAIL.n150 B 0.01403f
C323 VTAIL.n151 B 0.031319f
C324 VTAIL.n152 B 0.065741f
C325 VTAIL.n153 B 0.01403f
C326 VTAIL.n154 B 0.01325f
C327 VTAIL.n155 B 0.060029f
C328 VTAIL.n156 B 0.036664f
C329 VTAIL.n157 B 1.40229f
C330 VTAIL.n158 B 0.033495f
C331 VTAIL.n159 B 0.024659f
C332 VTAIL.n160 B 0.01325f
C333 VTAIL.n161 B 0.031319f
C334 VTAIL.n162 B 0.01364f
C335 VTAIL.n163 B 0.024659f
C336 VTAIL.n164 B 0.01403f
C337 VTAIL.n165 B 0.031319f
C338 VTAIL.n166 B 0.01403f
C339 VTAIL.n167 B 0.024659f
C340 VTAIL.n168 B 0.01325f
C341 VTAIL.n169 B 0.031319f
C342 VTAIL.n170 B 0.01403f
C343 VTAIL.n171 B 0.951127f
C344 VTAIL.n172 B 0.01325f
C345 VTAIL.t4 B 0.052545f
C346 VTAIL.n173 B 0.152516f
C347 VTAIL.n174 B 0.02214f
C348 VTAIL.n175 B 0.023489f
C349 VTAIL.n176 B 0.031319f
C350 VTAIL.n177 B 0.01403f
C351 VTAIL.n178 B 0.01325f
C352 VTAIL.n179 B 0.024659f
C353 VTAIL.n180 B 0.024659f
C354 VTAIL.n181 B 0.01325f
C355 VTAIL.n182 B 0.01403f
C356 VTAIL.n183 B 0.031319f
C357 VTAIL.n184 B 0.031319f
C358 VTAIL.n185 B 0.01403f
C359 VTAIL.n186 B 0.01325f
C360 VTAIL.n187 B 0.024659f
C361 VTAIL.n188 B 0.024659f
C362 VTAIL.n189 B 0.01325f
C363 VTAIL.n190 B 0.01325f
C364 VTAIL.n191 B 0.01403f
C365 VTAIL.n192 B 0.031319f
C366 VTAIL.n193 B 0.031319f
C367 VTAIL.n194 B 0.031319f
C368 VTAIL.n195 B 0.01364f
C369 VTAIL.n196 B 0.01325f
C370 VTAIL.n197 B 0.024659f
C371 VTAIL.n198 B 0.024659f
C372 VTAIL.n199 B 0.01325f
C373 VTAIL.n200 B 0.01403f
C374 VTAIL.n201 B 0.031319f
C375 VTAIL.n202 B 0.065741f
C376 VTAIL.n203 B 0.01403f
C377 VTAIL.n204 B 0.01325f
C378 VTAIL.n205 B 0.060029f
C379 VTAIL.n206 B 0.036664f
C380 VTAIL.n207 B 1.34698f
C381 VDD1.n0 B 0.029671f
C382 VDD1.n1 B 0.021843f
C383 VDD1.n2 B 0.011738f
C384 VDD1.n3 B 0.027743f
C385 VDD1.n4 B 0.012083f
C386 VDD1.n5 B 0.021843f
C387 VDD1.n6 B 0.012083f
C388 VDD1.n7 B 0.011738f
C389 VDD1.n8 B 0.027743f
C390 VDD1.n9 B 0.027743f
C391 VDD1.n10 B 0.012428f
C392 VDD1.n11 B 0.021843f
C393 VDD1.n12 B 0.011738f
C394 VDD1.n13 B 0.027743f
C395 VDD1.n14 B 0.012428f
C396 VDD1.n15 B 0.842534f
C397 VDD1.n16 B 0.011738f
C398 VDD1.t1 B 0.046546f
C399 VDD1.n17 B 0.135102f
C400 VDD1.n18 B 0.019612f
C401 VDD1.n19 B 0.020808f
C402 VDD1.n20 B 0.027743f
C403 VDD1.n21 B 0.012428f
C404 VDD1.n22 B 0.011738f
C405 VDD1.n23 B 0.021843f
C406 VDD1.n24 B 0.021843f
C407 VDD1.n25 B 0.011738f
C408 VDD1.n26 B 0.012428f
C409 VDD1.n27 B 0.027743f
C410 VDD1.n28 B 0.027743f
C411 VDD1.n29 B 0.012428f
C412 VDD1.n30 B 0.011738f
C413 VDD1.n31 B 0.021843f
C414 VDD1.n32 B 0.021843f
C415 VDD1.n33 B 0.011738f
C416 VDD1.n34 B 0.012428f
C417 VDD1.n35 B 0.027743f
C418 VDD1.n36 B 0.027743f
C419 VDD1.n37 B 0.012428f
C420 VDD1.n38 B 0.011738f
C421 VDD1.n39 B 0.021843f
C422 VDD1.n40 B 0.021843f
C423 VDD1.n41 B 0.011738f
C424 VDD1.n42 B 0.012428f
C425 VDD1.n43 B 0.027743f
C426 VDD1.n44 B 0.058235f
C427 VDD1.n45 B 0.012428f
C428 VDD1.n46 B 0.011738f
C429 VDD1.n47 B 0.053175f
C430 VDD1.n48 B 0.054381f
C431 VDD1.n49 B 0.029671f
C432 VDD1.n50 B 0.021843f
C433 VDD1.n51 B 0.011738f
C434 VDD1.n52 B 0.027743f
C435 VDD1.n53 B 0.012083f
C436 VDD1.n54 B 0.021843f
C437 VDD1.n55 B 0.012428f
C438 VDD1.n56 B 0.027743f
C439 VDD1.n57 B 0.012428f
C440 VDD1.n58 B 0.021843f
C441 VDD1.n59 B 0.011738f
C442 VDD1.n60 B 0.027743f
C443 VDD1.n61 B 0.012428f
C444 VDD1.n62 B 0.842534f
C445 VDD1.n63 B 0.011738f
C446 VDD1.t4 B 0.046546f
C447 VDD1.n64 B 0.135102f
C448 VDD1.n65 B 0.019612f
C449 VDD1.n66 B 0.020808f
C450 VDD1.n67 B 0.027743f
C451 VDD1.n68 B 0.012428f
C452 VDD1.n69 B 0.011738f
C453 VDD1.n70 B 0.021843f
C454 VDD1.n71 B 0.021843f
C455 VDD1.n72 B 0.011738f
C456 VDD1.n73 B 0.012428f
C457 VDD1.n74 B 0.027743f
C458 VDD1.n75 B 0.027743f
C459 VDD1.n76 B 0.012428f
C460 VDD1.n77 B 0.011738f
C461 VDD1.n78 B 0.021843f
C462 VDD1.n79 B 0.021843f
C463 VDD1.n80 B 0.011738f
C464 VDD1.n81 B 0.011738f
C465 VDD1.n82 B 0.012428f
C466 VDD1.n83 B 0.027743f
C467 VDD1.n84 B 0.027743f
C468 VDD1.n85 B 0.027743f
C469 VDD1.n86 B 0.012083f
C470 VDD1.n87 B 0.011738f
C471 VDD1.n88 B 0.021843f
C472 VDD1.n89 B 0.021843f
C473 VDD1.n90 B 0.011738f
C474 VDD1.n91 B 0.012428f
C475 VDD1.n92 B 0.027743f
C476 VDD1.n93 B 0.058235f
C477 VDD1.n94 B 0.012428f
C478 VDD1.n95 B 0.011738f
C479 VDD1.n96 B 0.053175f
C480 VDD1.n97 B 0.053727f
C481 VDD1.t5 B 0.161046f
C482 VDD1.t2 B 0.161046f
C483 VDD1.n98 B 1.41572f
C484 VDD1.n99 B 2.31344f
C485 VDD1.t0 B 0.161046f
C486 VDD1.t3 B 0.161046f
C487 VDD1.n100 B 1.4121f
C488 VDD1.n101 B 2.26162f
C489 VP.n0 B 0.032191f
C490 VP.t4 B 1.61908f
C491 VP.n1 B 0.037005f
C492 VP.n2 B 0.024417f
C493 VP.t0 B 1.61908f
C494 VP.n3 B 0.582156f
C495 VP.n4 B 0.024417f
C496 VP.n5 B 0.037005f
C497 VP.n6 B 0.032191f
C498 VP.t5 B 1.61908f
C499 VP.n7 B 0.032191f
C500 VP.t1 B 1.61908f
C501 VP.n8 B 0.037005f
C502 VP.n9 B 0.024417f
C503 VP.t2 B 1.61908f
C504 VP.n10 B 0.65301f
C505 VP.t3 B 1.82684f
C506 VP.n11 B 0.630149f
C507 VP.n12 B 0.236762f
C508 VP.n13 B 0.034273f
C509 VP.n14 B 0.045507f
C510 VP.n15 B 0.034283f
C511 VP.n16 B 0.024417f
C512 VP.n17 B 0.024417f
C513 VP.n18 B 0.024417f
C514 VP.n19 B 0.045507f
C515 VP.n20 B 0.032476f
C516 VP.n21 B 0.665493f
C517 VP.n22 B 1.2313f
C518 VP.n23 B 1.25005f
C519 VP.n24 B 0.665493f
C520 VP.n25 B 0.032476f
C521 VP.n26 B 0.045507f
C522 VP.n27 B 0.024417f
C523 VP.n28 B 0.024417f
C524 VP.n29 B 0.024417f
C525 VP.n30 B 0.034283f
C526 VP.n31 B 0.045507f
C527 VP.n32 B 0.034273f
C528 VP.n33 B 0.024417f
C529 VP.n34 B 0.024417f
C530 VP.n35 B 0.034273f
C531 VP.n36 B 0.045507f
C532 VP.n37 B 0.034283f
C533 VP.n38 B 0.024417f
C534 VP.n39 B 0.024417f
C535 VP.n40 B 0.024417f
C536 VP.n41 B 0.045507f
C537 VP.n42 B 0.032476f
C538 VP.n43 B 0.665493f
C539 VP.n44 B 0.039766f
.ends

