* NGSPICE file created from diff_pair_sample_0649.ext - technology: sky130A

.subckt diff_pair_sample_0649 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0 ps=0 w=1.8 l=0.53
X1 VDD1.t9 VP.t0 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X2 VTAIL.t9 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X3 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0 ps=0 w=1.8 l=0.53
X4 VDD1.t7 VP.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.702 ps=4.38 w=1.8 l=0.53
X5 VTAIL.t12 VP.t3 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X6 VTAIL.t19 VN.t0 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X7 VDD1.t5 VP.t4 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.702 ps=4.38 w=1.8 l=0.53
X8 VDD1.t4 VP.t5 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X9 VDD1.t3 VP.t6 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0.297 ps=2.13 w=1.8 l=0.53
X10 VDD1.t2 VP.t7 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0.297 ps=2.13 w=1.8 l=0.53
X11 VDD2.t8 VN.t1 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X12 VDD2.t7 VN.t2 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0.297 ps=2.13 w=1.8 l=0.53
X13 VTAIL.t16 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X14 VDD2.t5 VN.t4 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0.297 ps=2.13 w=1.8 l=0.53
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0 ps=0 w=1.8 l=0.53
X16 VTAIL.t6 VP.t8 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.702 pd=4.38 as=0 ps=0 w=1.8 l=0.53
X18 VDD2.t4 VN.t5 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.702 ps=4.38 w=1.8 l=0.53
X19 VDD2.t3 VN.t6 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.702 ps=4.38 w=1.8 l=0.53
X20 VTAIL.t3 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X21 VTAIL.t7 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X22 VDD2.t1 VN.t8 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
X23 VTAIL.t2 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.297 pd=2.13 as=0.297 ps=2.13 w=1.8 l=0.53
R0 B.n363 B.n362 585
R1 B.n364 B.n363 585
R2 B.n129 B.n63 585
R3 B.n128 B.n127 585
R4 B.n126 B.n125 585
R5 B.n124 B.n123 585
R6 B.n122 B.n121 585
R7 B.n120 B.n119 585
R8 B.n118 B.n117 585
R9 B.n116 B.n115 585
R10 B.n114 B.n113 585
R11 B.n112 B.n111 585
R12 B.n110 B.n109 585
R13 B.n107 B.n106 585
R14 B.n105 B.n104 585
R15 B.n103 B.n102 585
R16 B.n101 B.n100 585
R17 B.n99 B.n98 585
R18 B.n97 B.n96 585
R19 B.n95 B.n94 585
R20 B.n93 B.n92 585
R21 B.n91 B.n90 585
R22 B.n89 B.n88 585
R23 B.n87 B.n86 585
R24 B.n85 B.n84 585
R25 B.n83 B.n82 585
R26 B.n81 B.n80 585
R27 B.n79 B.n78 585
R28 B.n77 B.n76 585
R29 B.n75 B.n74 585
R30 B.n73 B.n72 585
R31 B.n71 B.n70 585
R32 B.n47 B.n46 585
R33 B.n367 B.n366 585
R34 B.n361 B.n64 585
R35 B.n64 B.n44 585
R36 B.n360 B.n43 585
R37 B.n371 B.n43 585
R38 B.n359 B.n42 585
R39 B.n372 B.n42 585
R40 B.n358 B.n41 585
R41 B.n373 B.n41 585
R42 B.n357 B.n356 585
R43 B.n356 B.n40 585
R44 B.n355 B.n36 585
R45 B.n379 B.n36 585
R46 B.n354 B.n35 585
R47 B.n380 B.n35 585
R48 B.n353 B.n34 585
R49 B.n381 B.n34 585
R50 B.n352 B.n351 585
R51 B.n351 B.n30 585
R52 B.n350 B.n29 585
R53 B.n387 B.n29 585
R54 B.n349 B.n28 585
R55 B.n388 B.n28 585
R56 B.n348 B.n27 585
R57 B.n389 B.n27 585
R58 B.n347 B.n346 585
R59 B.n346 B.n23 585
R60 B.n345 B.n22 585
R61 B.n395 B.n22 585
R62 B.n344 B.n21 585
R63 B.n396 B.n21 585
R64 B.n343 B.n20 585
R65 B.n397 B.n20 585
R66 B.n342 B.n341 585
R67 B.n341 B.n16 585
R68 B.n340 B.n15 585
R69 B.n403 B.n15 585
R70 B.n339 B.n14 585
R71 B.n404 B.n14 585
R72 B.n338 B.n13 585
R73 B.n405 B.n13 585
R74 B.n337 B.n336 585
R75 B.n336 B.n12 585
R76 B.n335 B.n334 585
R77 B.n335 B.n8 585
R78 B.n333 B.n7 585
R79 B.n412 B.n7 585
R80 B.n332 B.n6 585
R81 B.n413 B.n6 585
R82 B.n331 B.n5 585
R83 B.n414 B.n5 585
R84 B.n330 B.n329 585
R85 B.n329 B.n4 585
R86 B.n328 B.n130 585
R87 B.n328 B.n327 585
R88 B.n317 B.n131 585
R89 B.n320 B.n131 585
R90 B.n319 B.n318 585
R91 B.n321 B.n319 585
R92 B.n316 B.n135 585
R93 B.n139 B.n135 585
R94 B.n315 B.n314 585
R95 B.n314 B.n313 585
R96 B.n137 B.n136 585
R97 B.n138 B.n137 585
R98 B.n306 B.n305 585
R99 B.n307 B.n306 585
R100 B.n304 B.n144 585
R101 B.n144 B.n143 585
R102 B.n303 B.n302 585
R103 B.n302 B.n301 585
R104 B.n146 B.n145 585
R105 B.n147 B.n146 585
R106 B.n294 B.n293 585
R107 B.n295 B.n294 585
R108 B.n292 B.n151 585
R109 B.n155 B.n151 585
R110 B.n291 B.n290 585
R111 B.n290 B.n289 585
R112 B.n153 B.n152 585
R113 B.n154 B.n153 585
R114 B.n282 B.n281 585
R115 B.n283 B.n282 585
R116 B.n280 B.n160 585
R117 B.n160 B.n159 585
R118 B.n279 B.n278 585
R119 B.n278 B.n277 585
R120 B.n162 B.n161 585
R121 B.n270 B.n162 585
R122 B.n269 B.n268 585
R123 B.n271 B.n269 585
R124 B.n267 B.n167 585
R125 B.n167 B.n166 585
R126 B.n266 B.n265 585
R127 B.n265 B.n264 585
R128 B.n169 B.n168 585
R129 B.n170 B.n169 585
R130 B.n260 B.n259 585
R131 B.n173 B.n172 585
R132 B.n256 B.n255 585
R133 B.n257 B.n256 585
R134 B.n254 B.n189 585
R135 B.n253 B.n252 585
R136 B.n251 B.n250 585
R137 B.n249 B.n248 585
R138 B.n247 B.n246 585
R139 B.n245 B.n244 585
R140 B.n243 B.n242 585
R141 B.n241 B.n240 585
R142 B.n239 B.n238 585
R143 B.n236 B.n235 585
R144 B.n234 B.n233 585
R145 B.n232 B.n231 585
R146 B.n230 B.n229 585
R147 B.n228 B.n227 585
R148 B.n226 B.n225 585
R149 B.n224 B.n223 585
R150 B.n222 B.n221 585
R151 B.n220 B.n219 585
R152 B.n218 B.n217 585
R153 B.n216 B.n215 585
R154 B.n214 B.n213 585
R155 B.n212 B.n211 585
R156 B.n210 B.n209 585
R157 B.n208 B.n207 585
R158 B.n206 B.n205 585
R159 B.n204 B.n203 585
R160 B.n202 B.n201 585
R161 B.n200 B.n199 585
R162 B.n198 B.n197 585
R163 B.n196 B.n195 585
R164 B.n261 B.n171 585
R165 B.n171 B.n170 585
R166 B.n263 B.n262 585
R167 B.n264 B.n263 585
R168 B.n165 B.n164 585
R169 B.n166 B.n165 585
R170 B.n273 B.n272 585
R171 B.n272 B.n271 585
R172 B.n274 B.n163 585
R173 B.n270 B.n163 585
R174 B.n276 B.n275 585
R175 B.n277 B.n276 585
R176 B.n158 B.n157 585
R177 B.n159 B.n158 585
R178 B.n285 B.n284 585
R179 B.n284 B.n283 585
R180 B.n286 B.n156 585
R181 B.n156 B.n154 585
R182 B.n288 B.n287 585
R183 B.n289 B.n288 585
R184 B.n150 B.n149 585
R185 B.n155 B.n150 585
R186 B.n297 B.n296 585
R187 B.n296 B.n295 585
R188 B.n298 B.n148 585
R189 B.n148 B.n147 585
R190 B.n300 B.n299 585
R191 B.n301 B.n300 585
R192 B.n142 B.n141 585
R193 B.n143 B.n142 585
R194 B.n309 B.n308 585
R195 B.n308 B.n307 585
R196 B.n310 B.n140 585
R197 B.n140 B.n138 585
R198 B.n312 B.n311 585
R199 B.n313 B.n312 585
R200 B.n134 B.n133 585
R201 B.n139 B.n134 585
R202 B.n323 B.n322 585
R203 B.n322 B.n321 585
R204 B.n324 B.n132 585
R205 B.n320 B.n132 585
R206 B.n326 B.n325 585
R207 B.n327 B.n326 585
R208 B.n3 B.n0 585
R209 B.n4 B.n3 585
R210 B.n411 B.n1 585
R211 B.n412 B.n411 585
R212 B.n410 B.n409 585
R213 B.n410 B.n8 585
R214 B.n408 B.n9 585
R215 B.n12 B.n9 585
R216 B.n407 B.n406 585
R217 B.n406 B.n405 585
R218 B.n11 B.n10 585
R219 B.n404 B.n11 585
R220 B.n402 B.n401 585
R221 B.n403 B.n402 585
R222 B.n400 B.n17 585
R223 B.n17 B.n16 585
R224 B.n399 B.n398 585
R225 B.n398 B.n397 585
R226 B.n19 B.n18 585
R227 B.n396 B.n19 585
R228 B.n394 B.n393 585
R229 B.n395 B.n394 585
R230 B.n392 B.n24 585
R231 B.n24 B.n23 585
R232 B.n391 B.n390 585
R233 B.n390 B.n389 585
R234 B.n26 B.n25 585
R235 B.n388 B.n26 585
R236 B.n386 B.n385 585
R237 B.n387 B.n386 585
R238 B.n384 B.n31 585
R239 B.n31 B.n30 585
R240 B.n383 B.n382 585
R241 B.n382 B.n381 585
R242 B.n33 B.n32 585
R243 B.n380 B.n33 585
R244 B.n378 B.n377 585
R245 B.n379 B.n378 585
R246 B.n376 B.n37 585
R247 B.n40 B.n37 585
R248 B.n375 B.n374 585
R249 B.n374 B.n373 585
R250 B.n39 B.n38 585
R251 B.n372 B.n39 585
R252 B.n370 B.n369 585
R253 B.n371 B.n370 585
R254 B.n368 B.n45 585
R255 B.n45 B.n44 585
R256 B.n415 B.n414 585
R257 B.n413 B.n2 585
R258 B.n366 B.n45 449.257
R259 B.n363 B.n64 449.257
R260 B.n195 B.n169 449.257
R261 B.n259 B.n171 449.257
R262 B.n67 B.t17 287.575
R263 B.n65 B.t21 287.575
R264 B.n192 B.t14 287.575
R265 B.n190 B.t10 287.575
R266 B.n364 B.n62 256.663
R267 B.n364 B.n61 256.663
R268 B.n364 B.n60 256.663
R269 B.n364 B.n59 256.663
R270 B.n364 B.n58 256.663
R271 B.n364 B.n57 256.663
R272 B.n364 B.n56 256.663
R273 B.n364 B.n55 256.663
R274 B.n364 B.n54 256.663
R275 B.n364 B.n53 256.663
R276 B.n364 B.n52 256.663
R277 B.n364 B.n51 256.663
R278 B.n364 B.n50 256.663
R279 B.n364 B.n49 256.663
R280 B.n364 B.n48 256.663
R281 B.n365 B.n364 256.663
R282 B.n258 B.n257 256.663
R283 B.n257 B.n174 256.663
R284 B.n257 B.n175 256.663
R285 B.n257 B.n176 256.663
R286 B.n257 B.n177 256.663
R287 B.n257 B.n178 256.663
R288 B.n257 B.n179 256.663
R289 B.n257 B.n180 256.663
R290 B.n257 B.n181 256.663
R291 B.n257 B.n182 256.663
R292 B.n257 B.n183 256.663
R293 B.n257 B.n184 256.663
R294 B.n257 B.n185 256.663
R295 B.n257 B.n186 256.663
R296 B.n257 B.n187 256.663
R297 B.n257 B.n188 256.663
R298 B.n417 B.n416 256.663
R299 B.n257 B.n170 169.47
R300 B.n364 B.n44 169.47
R301 B.n70 B.n47 163.367
R302 B.n74 B.n73 163.367
R303 B.n78 B.n77 163.367
R304 B.n82 B.n81 163.367
R305 B.n86 B.n85 163.367
R306 B.n90 B.n89 163.367
R307 B.n94 B.n93 163.367
R308 B.n98 B.n97 163.367
R309 B.n102 B.n101 163.367
R310 B.n106 B.n105 163.367
R311 B.n111 B.n110 163.367
R312 B.n115 B.n114 163.367
R313 B.n119 B.n118 163.367
R314 B.n123 B.n122 163.367
R315 B.n127 B.n126 163.367
R316 B.n363 B.n63 163.367
R317 B.n265 B.n169 163.367
R318 B.n265 B.n167 163.367
R319 B.n269 B.n167 163.367
R320 B.n269 B.n162 163.367
R321 B.n278 B.n162 163.367
R322 B.n278 B.n160 163.367
R323 B.n282 B.n160 163.367
R324 B.n282 B.n153 163.367
R325 B.n290 B.n153 163.367
R326 B.n290 B.n151 163.367
R327 B.n294 B.n151 163.367
R328 B.n294 B.n146 163.367
R329 B.n302 B.n146 163.367
R330 B.n302 B.n144 163.367
R331 B.n306 B.n144 163.367
R332 B.n306 B.n137 163.367
R333 B.n314 B.n137 163.367
R334 B.n314 B.n135 163.367
R335 B.n319 B.n135 163.367
R336 B.n319 B.n131 163.367
R337 B.n328 B.n131 163.367
R338 B.n329 B.n328 163.367
R339 B.n329 B.n5 163.367
R340 B.n6 B.n5 163.367
R341 B.n7 B.n6 163.367
R342 B.n335 B.n7 163.367
R343 B.n336 B.n335 163.367
R344 B.n336 B.n13 163.367
R345 B.n14 B.n13 163.367
R346 B.n15 B.n14 163.367
R347 B.n341 B.n15 163.367
R348 B.n341 B.n20 163.367
R349 B.n21 B.n20 163.367
R350 B.n22 B.n21 163.367
R351 B.n346 B.n22 163.367
R352 B.n346 B.n27 163.367
R353 B.n28 B.n27 163.367
R354 B.n29 B.n28 163.367
R355 B.n351 B.n29 163.367
R356 B.n351 B.n34 163.367
R357 B.n35 B.n34 163.367
R358 B.n36 B.n35 163.367
R359 B.n356 B.n36 163.367
R360 B.n356 B.n41 163.367
R361 B.n42 B.n41 163.367
R362 B.n43 B.n42 163.367
R363 B.n64 B.n43 163.367
R364 B.n256 B.n173 163.367
R365 B.n256 B.n189 163.367
R366 B.n252 B.n251 163.367
R367 B.n248 B.n247 163.367
R368 B.n244 B.n243 163.367
R369 B.n240 B.n239 163.367
R370 B.n235 B.n234 163.367
R371 B.n231 B.n230 163.367
R372 B.n227 B.n226 163.367
R373 B.n223 B.n222 163.367
R374 B.n219 B.n218 163.367
R375 B.n215 B.n214 163.367
R376 B.n211 B.n210 163.367
R377 B.n207 B.n206 163.367
R378 B.n203 B.n202 163.367
R379 B.n199 B.n198 163.367
R380 B.n263 B.n171 163.367
R381 B.n263 B.n165 163.367
R382 B.n272 B.n165 163.367
R383 B.n272 B.n163 163.367
R384 B.n276 B.n163 163.367
R385 B.n276 B.n158 163.367
R386 B.n284 B.n158 163.367
R387 B.n284 B.n156 163.367
R388 B.n288 B.n156 163.367
R389 B.n288 B.n150 163.367
R390 B.n296 B.n150 163.367
R391 B.n296 B.n148 163.367
R392 B.n300 B.n148 163.367
R393 B.n300 B.n142 163.367
R394 B.n308 B.n142 163.367
R395 B.n308 B.n140 163.367
R396 B.n312 B.n140 163.367
R397 B.n312 B.n134 163.367
R398 B.n322 B.n134 163.367
R399 B.n322 B.n132 163.367
R400 B.n326 B.n132 163.367
R401 B.n326 B.n3 163.367
R402 B.n415 B.n3 163.367
R403 B.n411 B.n2 163.367
R404 B.n411 B.n410 163.367
R405 B.n410 B.n9 163.367
R406 B.n406 B.n9 163.367
R407 B.n406 B.n11 163.367
R408 B.n402 B.n11 163.367
R409 B.n402 B.n17 163.367
R410 B.n398 B.n17 163.367
R411 B.n398 B.n19 163.367
R412 B.n394 B.n19 163.367
R413 B.n394 B.n24 163.367
R414 B.n390 B.n24 163.367
R415 B.n390 B.n26 163.367
R416 B.n386 B.n26 163.367
R417 B.n386 B.n31 163.367
R418 B.n382 B.n31 163.367
R419 B.n382 B.n33 163.367
R420 B.n378 B.n33 163.367
R421 B.n378 B.n37 163.367
R422 B.n374 B.n37 163.367
R423 B.n374 B.n39 163.367
R424 B.n370 B.n39 163.367
R425 B.n370 B.n45 163.367
R426 B.n65 B.t22 135.819
R427 B.n192 B.t16 135.819
R428 B.n67 B.t19 135.819
R429 B.n190 B.t13 135.819
R430 B.n66 B.t23 119.139
R431 B.n193 B.t15 119.139
R432 B.n68 B.t20 119.139
R433 B.n191 B.t12 119.139
R434 B.n264 B.n170 105.725
R435 B.n264 B.n166 105.725
R436 B.n271 B.n166 105.725
R437 B.n271 B.n270 105.725
R438 B.n277 B.n159 105.725
R439 B.n283 B.n159 105.725
R440 B.n283 B.n154 105.725
R441 B.n289 B.n154 105.725
R442 B.n289 B.n155 105.725
R443 B.n295 B.n147 105.725
R444 B.n301 B.n147 105.725
R445 B.n307 B.n143 105.725
R446 B.n313 B.n138 105.725
R447 B.n313 B.n139 105.725
R448 B.n321 B.n320 105.725
R449 B.n327 B.n4 105.725
R450 B.n414 B.n4 105.725
R451 B.n414 B.n413 105.725
R452 B.n413 B.n412 105.725
R453 B.n412 B.n8 105.725
R454 B.n405 B.n12 105.725
R455 B.n404 B.n403 105.725
R456 B.n403 B.n16 105.725
R457 B.n397 B.n396 105.725
R458 B.n395 B.n23 105.725
R459 B.n389 B.n23 105.725
R460 B.n388 B.n387 105.725
R461 B.n387 B.n30 105.725
R462 B.n381 B.n30 105.725
R463 B.n381 B.n380 105.725
R464 B.n380 B.n379 105.725
R465 B.n373 B.n40 105.725
R466 B.n373 B.n372 105.725
R467 B.n372 B.n371 105.725
R468 B.n371 B.n44 105.725
R469 B.t2 B.n143 101.061
R470 B.n396 B.t7 101.061
R471 B.n321 B.t0 94.8415
R472 B.n405 B.t9 94.8415
R473 B.n270 B.t11 82.4033
R474 B.n40 B.t18 82.4033
R475 B.n366 B.n365 71.676
R476 B.n70 B.n48 71.676
R477 B.n74 B.n49 71.676
R478 B.n78 B.n50 71.676
R479 B.n82 B.n51 71.676
R480 B.n86 B.n52 71.676
R481 B.n90 B.n53 71.676
R482 B.n94 B.n54 71.676
R483 B.n98 B.n55 71.676
R484 B.n102 B.n56 71.676
R485 B.n106 B.n57 71.676
R486 B.n111 B.n58 71.676
R487 B.n115 B.n59 71.676
R488 B.n119 B.n60 71.676
R489 B.n123 B.n61 71.676
R490 B.n127 B.n62 71.676
R491 B.n63 B.n62 71.676
R492 B.n126 B.n61 71.676
R493 B.n122 B.n60 71.676
R494 B.n118 B.n59 71.676
R495 B.n114 B.n58 71.676
R496 B.n110 B.n57 71.676
R497 B.n105 B.n56 71.676
R498 B.n101 B.n55 71.676
R499 B.n97 B.n54 71.676
R500 B.n93 B.n53 71.676
R501 B.n89 B.n52 71.676
R502 B.n85 B.n51 71.676
R503 B.n81 B.n50 71.676
R504 B.n77 B.n49 71.676
R505 B.n73 B.n48 71.676
R506 B.n365 B.n47 71.676
R507 B.n259 B.n258 71.676
R508 B.n189 B.n174 71.676
R509 B.n251 B.n175 71.676
R510 B.n247 B.n176 71.676
R511 B.n243 B.n177 71.676
R512 B.n239 B.n178 71.676
R513 B.n234 B.n179 71.676
R514 B.n230 B.n180 71.676
R515 B.n226 B.n181 71.676
R516 B.n222 B.n182 71.676
R517 B.n218 B.n183 71.676
R518 B.n214 B.n184 71.676
R519 B.n210 B.n185 71.676
R520 B.n206 B.n186 71.676
R521 B.n202 B.n187 71.676
R522 B.n198 B.n188 71.676
R523 B.n258 B.n173 71.676
R524 B.n252 B.n174 71.676
R525 B.n248 B.n175 71.676
R526 B.n244 B.n176 71.676
R527 B.n240 B.n177 71.676
R528 B.n235 B.n178 71.676
R529 B.n231 B.n179 71.676
R530 B.n227 B.n180 71.676
R531 B.n223 B.n181 71.676
R532 B.n219 B.n182 71.676
R533 B.n215 B.n183 71.676
R534 B.n211 B.n184 71.676
R535 B.n207 B.n185 71.676
R536 B.n203 B.n186 71.676
R537 B.n199 B.n187 71.676
R538 B.n195 B.n188 71.676
R539 B.n416 B.n415 71.676
R540 B.n416 B.n2 71.676
R541 B.n320 B.t5 66.8556
R542 B.n12 B.t8 66.8556
R543 B.n307 B.t4 60.6365
R544 B.n397 B.t6 60.6365
R545 B.n69 B.n68 59.5399
R546 B.n108 B.n66 59.5399
R547 B.n194 B.n193 59.5399
R548 B.n237 B.n191 59.5399
R549 B.n155 B.t3 54.4175
R550 B.t1 B.n388 54.4175
R551 B.n295 B.t3 51.3079
R552 B.n389 B.t1 51.3079
R553 B.t4 B.n138 45.0888
R554 B.t6 B.n16 45.0888
R555 B.n327 B.t5 38.8698
R556 B.t8 B.n8 38.8698
R557 B.n261 B.n260 29.1907
R558 B.n196 B.n168 29.1907
R559 B.n368 B.n367 29.1907
R560 B.n362 B.n361 29.1907
R561 B.n277 B.t11 23.3221
R562 B.n379 B.t18 23.3221
R563 B B.n417 18.0485
R564 B.n68 B.n67 16.6793
R565 B.n66 B.n65 16.6793
R566 B.n193 B.n192 16.6793
R567 B.n191 B.n190 16.6793
R568 B.n139 B.t0 10.8839
R569 B.t9 B.n404 10.8839
R570 B.n262 B.n261 10.6151
R571 B.n262 B.n164 10.6151
R572 B.n273 B.n164 10.6151
R573 B.n274 B.n273 10.6151
R574 B.n275 B.n274 10.6151
R575 B.n275 B.n157 10.6151
R576 B.n285 B.n157 10.6151
R577 B.n286 B.n285 10.6151
R578 B.n287 B.n286 10.6151
R579 B.n287 B.n149 10.6151
R580 B.n297 B.n149 10.6151
R581 B.n298 B.n297 10.6151
R582 B.n299 B.n298 10.6151
R583 B.n299 B.n141 10.6151
R584 B.n309 B.n141 10.6151
R585 B.n310 B.n309 10.6151
R586 B.n311 B.n310 10.6151
R587 B.n311 B.n133 10.6151
R588 B.n323 B.n133 10.6151
R589 B.n324 B.n323 10.6151
R590 B.n325 B.n324 10.6151
R591 B.n325 B.n0 10.6151
R592 B.n260 B.n172 10.6151
R593 B.n255 B.n172 10.6151
R594 B.n255 B.n254 10.6151
R595 B.n254 B.n253 10.6151
R596 B.n253 B.n250 10.6151
R597 B.n250 B.n249 10.6151
R598 B.n249 B.n246 10.6151
R599 B.n246 B.n245 10.6151
R600 B.n245 B.n242 10.6151
R601 B.n242 B.n241 10.6151
R602 B.n241 B.n238 10.6151
R603 B.n236 B.n233 10.6151
R604 B.n233 B.n232 10.6151
R605 B.n232 B.n229 10.6151
R606 B.n229 B.n228 10.6151
R607 B.n228 B.n225 10.6151
R608 B.n225 B.n224 10.6151
R609 B.n224 B.n221 10.6151
R610 B.n221 B.n220 10.6151
R611 B.n217 B.n216 10.6151
R612 B.n216 B.n213 10.6151
R613 B.n213 B.n212 10.6151
R614 B.n212 B.n209 10.6151
R615 B.n209 B.n208 10.6151
R616 B.n208 B.n205 10.6151
R617 B.n205 B.n204 10.6151
R618 B.n204 B.n201 10.6151
R619 B.n201 B.n200 10.6151
R620 B.n200 B.n197 10.6151
R621 B.n197 B.n196 10.6151
R622 B.n266 B.n168 10.6151
R623 B.n267 B.n266 10.6151
R624 B.n268 B.n267 10.6151
R625 B.n268 B.n161 10.6151
R626 B.n279 B.n161 10.6151
R627 B.n280 B.n279 10.6151
R628 B.n281 B.n280 10.6151
R629 B.n281 B.n152 10.6151
R630 B.n291 B.n152 10.6151
R631 B.n292 B.n291 10.6151
R632 B.n293 B.n292 10.6151
R633 B.n293 B.n145 10.6151
R634 B.n303 B.n145 10.6151
R635 B.n304 B.n303 10.6151
R636 B.n305 B.n304 10.6151
R637 B.n305 B.n136 10.6151
R638 B.n315 B.n136 10.6151
R639 B.n316 B.n315 10.6151
R640 B.n318 B.n316 10.6151
R641 B.n318 B.n317 10.6151
R642 B.n317 B.n130 10.6151
R643 B.n330 B.n130 10.6151
R644 B.n331 B.n330 10.6151
R645 B.n332 B.n331 10.6151
R646 B.n333 B.n332 10.6151
R647 B.n334 B.n333 10.6151
R648 B.n337 B.n334 10.6151
R649 B.n338 B.n337 10.6151
R650 B.n339 B.n338 10.6151
R651 B.n340 B.n339 10.6151
R652 B.n342 B.n340 10.6151
R653 B.n343 B.n342 10.6151
R654 B.n344 B.n343 10.6151
R655 B.n345 B.n344 10.6151
R656 B.n347 B.n345 10.6151
R657 B.n348 B.n347 10.6151
R658 B.n349 B.n348 10.6151
R659 B.n350 B.n349 10.6151
R660 B.n352 B.n350 10.6151
R661 B.n353 B.n352 10.6151
R662 B.n354 B.n353 10.6151
R663 B.n355 B.n354 10.6151
R664 B.n357 B.n355 10.6151
R665 B.n358 B.n357 10.6151
R666 B.n359 B.n358 10.6151
R667 B.n360 B.n359 10.6151
R668 B.n361 B.n360 10.6151
R669 B.n409 B.n1 10.6151
R670 B.n409 B.n408 10.6151
R671 B.n408 B.n407 10.6151
R672 B.n407 B.n10 10.6151
R673 B.n401 B.n10 10.6151
R674 B.n401 B.n400 10.6151
R675 B.n400 B.n399 10.6151
R676 B.n399 B.n18 10.6151
R677 B.n393 B.n18 10.6151
R678 B.n393 B.n392 10.6151
R679 B.n392 B.n391 10.6151
R680 B.n391 B.n25 10.6151
R681 B.n385 B.n25 10.6151
R682 B.n385 B.n384 10.6151
R683 B.n384 B.n383 10.6151
R684 B.n383 B.n32 10.6151
R685 B.n377 B.n32 10.6151
R686 B.n377 B.n376 10.6151
R687 B.n376 B.n375 10.6151
R688 B.n375 B.n38 10.6151
R689 B.n369 B.n38 10.6151
R690 B.n369 B.n368 10.6151
R691 B.n367 B.n46 10.6151
R692 B.n71 B.n46 10.6151
R693 B.n72 B.n71 10.6151
R694 B.n75 B.n72 10.6151
R695 B.n76 B.n75 10.6151
R696 B.n79 B.n76 10.6151
R697 B.n80 B.n79 10.6151
R698 B.n83 B.n80 10.6151
R699 B.n84 B.n83 10.6151
R700 B.n87 B.n84 10.6151
R701 B.n88 B.n87 10.6151
R702 B.n92 B.n91 10.6151
R703 B.n95 B.n92 10.6151
R704 B.n96 B.n95 10.6151
R705 B.n99 B.n96 10.6151
R706 B.n100 B.n99 10.6151
R707 B.n103 B.n100 10.6151
R708 B.n104 B.n103 10.6151
R709 B.n107 B.n104 10.6151
R710 B.n112 B.n109 10.6151
R711 B.n113 B.n112 10.6151
R712 B.n116 B.n113 10.6151
R713 B.n117 B.n116 10.6151
R714 B.n120 B.n117 10.6151
R715 B.n121 B.n120 10.6151
R716 B.n124 B.n121 10.6151
R717 B.n125 B.n124 10.6151
R718 B.n128 B.n125 10.6151
R719 B.n129 B.n128 10.6151
R720 B.n362 B.n129 10.6151
R721 B.n417 B.n0 8.11757
R722 B.n417 B.n1 8.11757
R723 B.n237 B.n236 6.5566
R724 B.n220 B.n194 6.5566
R725 B.n91 B.n69 6.5566
R726 B.n108 B.n107 6.5566
R727 B.n301 B.t2 4.66481
R728 B.t7 B.n395 4.66481
R729 B.n238 B.n237 4.05904
R730 B.n217 B.n194 4.05904
R731 B.n88 B.n69 4.05904
R732 B.n109 B.n108 4.05904
R733 VP.n5 VP.t7 176.951
R734 VP.n25 VP.n24 161.3
R735 VP.n8 VP.n7 161.3
R736 VP.n9 VP.n4 161.3
R737 VP.n11 VP.n10 161.3
R738 VP.n12 VP.n3 161.3
R739 VP.n14 VP.n13 161.3
R740 VP.n23 VP.n0 161.3
R741 VP.n22 VP.n21 161.3
R742 VP.n20 VP.n1 161.3
R743 VP.n19 VP.n18 161.3
R744 VP.n17 VP.n2 161.3
R745 VP.n16 VP.n15 161.3
R746 VP.n16 VP.t6 155.969
R747 VP.n17 VP.t3 155.969
R748 VP.n1 VP.t5 155.969
R749 VP.n23 VP.t1 155.969
R750 VP.n24 VP.t4 155.969
R751 VP.n13 VP.t2 155.969
R752 VP.n12 VP.t8 155.969
R753 VP.n4 VP.t0 155.969
R754 VP.n6 VP.t9 155.969
R755 VP.n8 VP.n5 70.4033
R756 VP.n17 VP.n16 48.2005
R757 VP.n24 VP.n23 48.2005
R758 VP.n13 VP.n12 48.2005
R759 VP.n18 VP.n1 34.3247
R760 VP.n22 VP.n1 34.3247
R761 VP.n11 VP.n4 34.3247
R762 VP.n7 VP.n4 34.3247
R763 VP.n15 VP.n14 34.2126
R764 VP.n6 VP.n5 20.9576
R765 VP.n18 VP.n17 13.8763
R766 VP.n23 VP.n22 13.8763
R767 VP.n12 VP.n11 13.8763
R768 VP.n7 VP.n6 13.8763
R769 VP.n9 VP.n8 0.189894
R770 VP.n10 VP.n9 0.189894
R771 VP.n10 VP.n3 0.189894
R772 VP.n14 VP.n3 0.189894
R773 VP.n15 VP.n2 0.189894
R774 VP.n19 VP.n2 0.189894
R775 VP.n20 VP.n19 0.189894
R776 VP.n21 VP.n20 0.189894
R777 VP.n21 VP.n0 0.189894
R778 VP.n25 VP.n0 0.189894
R779 VP VP.n25 0.0516364
R780 VTAIL.n40 VTAIL.n38 289.615
R781 VTAIL.n4 VTAIL.n2 289.615
R782 VTAIL.n32 VTAIL.n30 289.615
R783 VTAIL.n20 VTAIL.n18 289.615
R784 VTAIL.n41 VTAIL.n40 185
R785 VTAIL.n5 VTAIL.n4 185
R786 VTAIL.n33 VTAIL.n32 185
R787 VTAIL.n21 VTAIL.n20 185
R788 VTAIL.t14 VTAIL.n39 164.876
R789 VTAIL.t13 VTAIL.n3 164.876
R790 VTAIL.t10 VTAIL.n31 164.876
R791 VTAIL.t18 VTAIL.n19 164.876
R792 VTAIL.n29 VTAIL.n28 85.1322
R793 VTAIL.n27 VTAIL.n26 85.1322
R794 VTAIL.n17 VTAIL.n16 85.1322
R795 VTAIL.n15 VTAIL.n14 85.1322
R796 VTAIL.n47 VTAIL.n46 85.1321
R797 VTAIL.n1 VTAIL.n0 85.1321
R798 VTAIL.n11 VTAIL.n10 85.1321
R799 VTAIL.n13 VTAIL.n12 85.1321
R800 VTAIL.n40 VTAIL.t14 52.3082
R801 VTAIL.n4 VTAIL.t13 52.3082
R802 VTAIL.n32 VTAIL.t10 52.3082
R803 VTAIL.n20 VTAIL.t18 52.3082
R804 VTAIL.n45 VTAIL.n44 34.5126
R805 VTAIL.n9 VTAIL.n8 34.5126
R806 VTAIL.n37 VTAIL.n36 34.5126
R807 VTAIL.n25 VTAIL.n24 34.5126
R808 VTAIL.n15 VTAIL.n13 15.4014
R809 VTAIL.n41 VTAIL.n39 14.7318
R810 VTAIL.n5 VTAIL.n3 14.7318
R811 VTAIL.n33 VTAIL.n31 14.7318
R812 VTAIL.n21 VTAIL.n19 14.7318
R813 VTAIL.n45 VTAIL.n37 14.66
R814 VTAIL.n42 VTAIL.n38 12.8005
R815 VTAIL.n6 VTAIL.n2 12.8005
R816 VTAIL.n34 VTAIL.n30 12.8005
R817 VTAIL.n22 VTAIL.n18 12.8005
R818 VTAIL.n46 VTAIL.t15 11.0005
R819 VTAIL.n46 VTAIL.t3 11.0005
R820 VTAIL.n0 VTAIL.t17 11.0005
R821 VTAIL.n0 VTAIL.t16 11.0005
R822 VTAIL.n10 VTAIL.t11 11.0005
R823 VTAIL.n10 VTAIL.t9 11.0005
R824 VTAIL.n12 VTAIL.t4 11.0005
R825 VTAIL.n12 VTAIL.t12 11.0005
R826 VTAIL.n28 VTAIL.t8 11.0005
R827 VTAIL.n28 VTAIL.t6 11.0005
R828 VTAIL.n26 VTAIL.t5 11.0005
R829 VTAIL.n26 VTAIL.t7 11.0005
R830 VTAIL.n16 VTAIL.t1 11.0005
R831 VTAIL.n16 VTAIL.t19 11.0005
R832 VTAIL.n14 VTAIL.t0 11.0005
R833 VTAIL.n14 VTAIL.t2 11.0005
R834 VTAIL.n44 VTAIL.n43 9.45567
R835 VTAIL.n8 VTAIL.n7 9.45567
R836 VTAIL.n36 VTAIL.n35 9.45567
R837 VTAIL.n24 VTAIL.n23 9.45567
R838 VTAIL.n43 VTAIL.n42 9.3005
R839 VTAIL.n7 VTAIL.n6 9.3005
R840 VTAIL.n35 VTAIL.n34 9.3005
R841 VTAIL.n23 VTAIL.n22 9.3005
R842 VTAIL.n43 VTAIL.n39 5.62509
R843 VTAIL.n7 VTAIL.n3 5.62509
R844 VTAIL.n35 VTAIL.n31 5.62509
R845 VTAIL.n23 VTAIL.n19 5.62509
R846 VTAIL.n44 VTAIL.n38 1.16414
R847 VTAIL.n8 VTAIL.n2 1.16414
R848 VTAIL.n36 VTAIL.n30 1.16414
R849 VTAIL.n24 VTAIL.n18 1.16414
R850 VTAIL.n27 VTAIL.n25 0.841017
R851 VTAIL.n9 VTAIL.n1 0.841017
R852 VTAIL.n17 VTAIL.n15 0.741879
R853 VTAIL.n25 VTAIL.n17 0.741879
R854 VTAIL.n29 VTAIL.n27 0.741879
R855 VTAIL.n37 VTAIL.n29 0.741879
R856 VTAIL.n13 VTAIL.n11 0.741879
R857 VTAIL.n11 VTAIL.n9 0.741879
R858 VTAIL.n47 VTAIL.n45 0.741879
R859 VTAIL VTAIL.n1 0.614724
R860 VTAIL.n42 VTAIL.n41 0.388379
R861 VTAIL.n6 VTAIL.n5 0.388379
R862 VTAIL.n34 VTAIL.n33 0.388379
R863 VTAIL.n22 VTAIL.n21 0.388379
R864 VTAIL VTAIL.n47 0.127655
R865 VDD1.n2 VDD1.n0 289.615
R866 VDD1.n11 VDD1.n9 289.615
R867 VDD1.n3 VDD1.n2 185
R868 VDD1.n12 VDD1.n11 185
R869 VDD1.t2 VDD1.n1 164.876
R870 VDD1.t3 VDD1.n10 164.876
R871 VDD1.n19 VDD1.n18 102.311
R872 VDD1.n21 VDD1.n20 101.811
R873 VDD1.n8 VDD1.n7 101.811
R874 VDD1.n17 VDD1.n16 101.811
R875 VDD1.n2 VDD1.t2 52.3082
R876 VDD1.n11 VDD1.t3 52.3082
R877 VDD1.n8 VDD1.n6 51.9328
R878 VDD1.n17 VDD1.n15 51.9328
R879 VDD1.n21 VDD1.n19 29.7423
R880 VDD1.n3 VDD1.n1 14.7318
R881 VDD1.n12 VDD1.n10 14.7318
R882 VDD1.n4 VDD1.n0 12.8005
R883 VDD1.n13 VDD1.n9 12.8005
R884 VDD1.n20 VDD1.t1 11.0005
R885 VDD1.n20 VDD1.t7 11.0005
R886 VDD1.n7 VDD1.t0 11.0005
R887 VDD1.n7 VDD1.t9 11.0005
R888 VDD1.n18 VDD1.t8 11.0005
R889 VDD1.n18 VDD1.t5 11.0005
R890 VDD1.n16 VDD1.t6 11.0005
R891 VDD1.n16 VDD1.t4 11.0005
R892 VDD1.n6 VDD1.n5 9.45567
R893 VDD1.n15 VDD1.n14 9.45567
R894 VDD1.n5 VDD1.n4 9.3005
R895 VDD1.n14 VDD1.n13 9.3005
R896 VDD1.n5 VDD1.n1 5.62509
R897 VDD1.n14 VDD1.n10 5.62509
R898 VDD1.n6 VDD1.n0 1.16414
R899 VDD1.n15 VDD1.n9 1.16414
R900 VDD1 VDD1.n21 0.498345
R901 VDD1.n4 VDD1.n3 0.388379
R902 VDD1.n13 VDD1.n12 0.388379
R903 VDD1 VDD1.n8 0.244034
R904 VDD1.n19 VDD1.n17 0.130499
R905 VN.n2 VN.t4 176.951
R906 VN.n14 VN.t5 176.951
R907 VN.n11 VN.n10 161.3
R908 VN.n23 VN.n22 161.3
R909 VN.n21 VN.n12 161.3
R910 VN.n20 VN.n19 161.3
R911 VN.n18 VN.n13 161.3
R912 VN.n17 VN.n16 161.3
R913 VN.n9 VN.n0 161.3
R914 VN.n8 VN.n7 161.3
R915 VN.n6 VN.n1 161.3
R916 VN.n5 VN.n4 161.3
R917 VN.n3 VN.t3 155.969
R918 VN.n1 VN.t8 155.969
R919 VN.n9 VN.t7 155.969
R920 VN.n10 VN.t6 155.969
R921 VN.n15 VN.t0 155.969
R922 VN.n13 VN.t1 155.969
R923 VN.n21 VN.t9 155.969
R924 VN.n22 VN.t2 155.969
R925 VN.n17 VN.n14 70.4033
R926 VN.n5 VN.n2 70.4033
R927 VN.n10 VN.n9 48.2005
R928 VN.n22 VN.n21 48.2005
R929 VN VN.n23 34.5933
R930 VN.n4 VN.n1 34.3247
R931 VN.n8 VN.n1 34.3247
R932 VN.n16 VN.n13 34.3247
R933 VN.n20 VN.n13 34.3247
R934 VN.n15 VN.n14 20.9576
R935 VN.n3 VN.n2 20.9576
R936 VN.n4 VN.n3 13.8763
R937 VN.n9 VN.n8 13.8763
R938 VN.n16 VN.n15 13.8763
R939 VN.n21 VN.n20 13.8763
R940 VN.n23 VN.n12 0.189894
R941 VN.n19 VN.n12 0.189894
R942 VN.n19 VN.n18 0.189894
R943 VN.n18 VN.n17 0.189894
R944 VN.n6 VN.n5 0.189894
R945 VN.n7 VN.n6 0.189894
R946 VN.n7 VN.n0 0.189894
R947 VN.n11 VN.n0 0.189894
R948 VN VN.n11 0.0516364
R949 VDD2.n13 VDD2.n11 289.615
R950 VDD2.n2 VDD2.n0 289.615
R951 VDD2.n14 VDD2.n13 185
R952 VDD2.n3 VDD2.n2 185
R953 VDD2.t7 VDD2.n12 164.876
R954 VDD2.t5 VDD2.n1 164.876
R955 VDD2.n10 VDD2.n9 102.311
R956 VDD2 VDD2.n21 102.308
R957 VDD2.n20 VDD2.n19 101.811
R958 VDD2.n8 VDD2.n7 101.811
R959 VDD2.n13 VDD2.t7 52.3082
R960 VDD2.n2 VDD2.t5 52.3082
R961 VDD2.n8 VDD2.n6 51.9328
R962 VDD2.n18 VDD2.n17 51.1914
R963 VDD2.n18 VDD2.n10 28.7886
R964 VDD2.n14 VDD2.n12 14.7318
R965 VDD2.n3 VDD2.n1 14.7318
R966 VDD2.n15 VDD2.n11 12.8005
R967 VDD2.n4 VDD2.n0 12.8005
R968 VDD2.n21 VDD2.t9 11.0005
R969 VDD2.n21 VDD2.t4 11.0005
R970 VDD2.n19 VDD2.t0 11.0005
R971 VDD2.n19 VDD2.t8 11.0005
R972 VDD2.n9 VDD2.t2 11.0005
R973 VDD2.n9 VDD2.t3 11.0005
R974 VDD2.n7 VDD2.t6 11.0005
R975 VDD2.n7 VDD2.t1 11.0005
R976 VDD2.n17 VDD2.n16 9.45567
R977 VDD2.n6 VDD2.n5 9.45567
R978 VDD2.n16 VDD2.n15 9.3005
R979 VDD2.n5 VDD2.n4 9.3005
R980 VDD2.n16 VDD2.n12 5.62509
R981 VDD2.n5 VDD2.n1 5.62509
R982 VDD2.n17 VDD2.n11 1.16414
R983 VDD2.n6 VDD2.n0 1.16414
R984 VDD2.n20 VDD2.n18 0.741879
R985 VDD2.n15 VDD2.n14 0.388379
R986 VDD2.n4 VDD2.n3 0.388379
R987 VDD2 VDD2.n20 0.244034
R988 VDD2.n10 VDD2.n8 0.130499
C0 VDD1 VTAIL 4.3925f
C1 VP VTAIL 1.49587f
C2 VN VDD2 1.2135f
C3 VN VDD1 0.155657f
C4 VDD2 VDD1 0.863261f
C5 VN VP 3.46076f
C6 VP VDD2 0.326154f
C7 VN VTAIL 1.48168f
C8 VDD2 VTAIL 4.4311f
C9 VP VDD1 1.38203f
C10 VDD2 B 2.837882f
C11 VDD1 B 2.841364f
C12 VTAIL B 2.456654f
C13 VN B 6.768781f
C14 VP B 5.818003f
C15 VDD2.n0 B 0.026364f
C16 VDD2.n1 B 0.061784f
C17 VDD2.t5 B 0.044204f
C18 VDD2.n2 B 0.045555f
C19 VDD2.n3 B 0.013175f
C20 VDD2.n4 B 0.010695f
C21 VDD2.n5 B 0.120724f
C22 VDD2.n6 B 0.043801f
C23 VDD2.t6 B 0.02831f
C24 VDD2.t1 B 0.02831f
C25 VDD2.n7 B 0.181279f
C26 VDD2.n8 B 0.284656f
C27 VDD2.t2 B 0.02831f
C28 VDD2.t3 B 0.02831f
C29 VDD2.n9 B 0.182391f
C30 VDD2.n10 B 0.946618f
C31 VDD2.n11 B 0.026364f
C32 VDD2.n12 B 0.061784f
C33 VDD2.t7 B 0.044204f
C34 VDD2.n13 B 0.045555f
C35 VDD2.n14 B 0.013175f
C36 VDD2.n15 B 0.010695f
C37 VDD2.n16 B 0.120724f
C38 VDD2.n17 B 0.042549f
C39 VDD2.n18 B 1.00899f
C40 VDD2.t0 B 0.02831f
C41 VDD2.t8 B 0.02831f
C42 VDD2.n19 B 0.181279f
C43 VDD2.n20 B 0.201901f
C44 VDD2.t9 B 0.02831f
C45 VDD2.t4 B 0.02831f
C46 VDD2.n21 B 0.18238f
C47 VN.n0 B 0.027837f
C48 VN.t8 B 0.083106f
C49 VN.n1 B 0.065088f
C50 VN.t4 B 0.090544f
C51 VN.n2 B 0.055461f
C52 VN.t3 B 0.083106f
C53 VN.n3 B 0.064316f
C54 VN.n4 B 0.006317f
C55 VN.n5 B 0.091364f
C56 VN.n6 B 0.027837f
C57 VN.n7 B 0.027837f
C58 VN.n8 B 0.006317f
C59 VN.t7 B 0.083106f
C60 VN.n9 B 0.064316f
C61 VN.t6 B 0.083106f
C62 VN.n10 B 0.062686f
C63 VN.n11 B 0.021573f
C64 VN.n12 B 0.027837f
C65 VN.t1 B 0.083106f
C66 VN.n13 B 0.065088f
C67 VN.t5 B 0.090544f
C68 VN.n14 B 0.055461f
C69 VN.t0 B 0.083106f
C70 VN.n15 B 0.064316f
C71 VN.n16 B 0.006317f
C72 VN.n17 B 0.091364f
C73 VN.n18 B 0.027837f
C74 VN.n19 B 0.027837f
C75 VN.n20 B 0.006317f
C76 VN.t9 B 0.083106f
C77 VN.n21 B 0.064316f
C78 VN.t2 B 0.083106f
C79 VN.n22 B 0.062686f
C80 VN.n23 B 0.811961f
C81 VDD1.n0 B 0.025931f
C82 VDD1.n1 B 0.060769f
C83 VDD1.t2 B 0.043477f
C84 VDD1.n2 B 0.044807f
C85 VDD1.n3 B 0.012959f
C86 VDD1.n4 B 0.010519f
C87 VDD1.n5 B 0.118741f
C88 VDD1.n6 B 0.043082f
C89 VDD1.t0 B 0.027845f
C90 VDD1.t9 B 0.027845f
C91 VDD1.n7 B 0.178301f
C92 VDD1.n8 B 0.283648f
C93 VDD1.n9 B 0.025931f
C94 VDD1.n10 B 0.060769f
C95 VDD1.t3 B 0.043477f
C96 VDD1.n11 B 0.044807f
C97 VDD1.n12 B 0.012959f
C98 VDD1.n13 B 0.010519f
C99 VDD1.n14 B 0.118741f
C100 VDD1.n15 B 0.043082f
C101 VDD1.t6 B 0.027845f
C102 VDD1.t4 B 0.027845f
C103 VDD1.n16 B 0.1783f
C104 VDD1.n17 B 0.279978f
C105 VDD1.t8 B 0.027845f
C106 VDD1.t5 B 0.027845f
C107 VDD1.n18 B 0.179394f
C108 VDD1.n19 B 0.984847f
C109 VDD1.t1 B 0.027845f
C110 VDD1.t7 B 0.027845f
C111 VDD1.n20 B 0.178301f
C112 VDD1.n21 B 1.14714f
C113 VTAIL.t17 B 0.035496f
C114 VTAIL.t16 B 0.035496f
C115 VTAIL.n0 B 0.194144f
C116 VTAIL.n1 B 0.290162f
C117 VTAIL.n2 B 0.033056f
C118 VTAIL.n3 B 0.077467f
C119 VTAIL.t13 B 0.055424f
C120 VTAIL.n4 B 0.057119f
C121 VTAIL.n5 B 0.01652f
C122 VTAIL.n6 B 0.01341f
C123 VTAIL.n7 B 0.151368f
C124 VTAIL.n8 B 0.036148f
C125 VTAIL.n9 B 0.150826f
C126 VTAIL.t11 B 0.035496f
C127 VTAIL.t9 B 0.035496f
C128 VTAIL.n10 B 0.194144f
C129 VTAIL.n11 B 0.292415f
C130 VTAIL.t4 B 0.035496f
C131 VTAIL.t12 B 0.035496f
C132 VTAIL.n12 B 0.194144f
C133 VTAIL.n13 B 0.815784f
C134 VTAIL.t0 B 0.035496f
C135 VTAIL.t2 B 0.035496f
C136 VTAIL.n14 B 0.194145f
C137 VTAIL.n15 B 0.815783f
C138 VTAIL.t1 B 0.035496f
C139 VTAIL.t19 B 0.035496f
C140 VTAIL.n16 B 0.194145f
C141 VTAIL.n17 B 0.292414f
C142 VTAIL.n18 B 0.033056f
C143 VTAIL.n19 B 0.077467f
C144 VTAIL.t18 B 0.055424f
C145 VTAIL.n20 B 0.057119f
C146 VTAIL.n21 B 0.01652f
C147 VTAIL.n22 B 0.01341f
C148 VTAIL.n23 B 0.151368f
C149 VTAIL.n24 B 0.036148f
C150 VTAIL.n25 B 0.150826f
C151 VTAIL.t5 B 0.035496f
C152 VTAIL.t7 B 0.035496f
C153 VTAIL.n26 B 0.194145f
C154 VTAIL.n27 B 0.300385f
C155 VTAIL.t8 B 0.035496f
C156 VTAIL.t6 B 0.035496f
C157 VTAIL.n28 B 0.194145f
C158 VTAIL.n29 B 0.292414f
C159 VTAIL.n30 B 0.033056f
C160 VTAIL.n31 B 0.077467f
C161 VTAIL.t10 B 0.055424f
C162 VTAIL.n32 B 0.057119f
C163 VTAIL.n33 B 0.01652f
C164 VTAIL.n34 B 0.01341f
C165 VTAIL.n35 B 0.151368f
C166 VTAIL.n36 B 0.036148f
C167 VTAIL.n37 B 0.606609f
C168 VTAIL.n38 B 0.033056f
C169 VTAIL.n39 B 0.077467f
C170 VTAIL.t14 B 0.055424f
C171 VTAIL.n40 B 0.057119f
C172 VTAIL.n41 B 0.01652f
C173 VTAIL.n42 B 0.01341f
C174 VTAIL.n43 B 0.151368f
C175 VTAIL.n44 B 0.036148f
C176 VTAIL.n45 B 0.606609f
C177 VTAIL.t15 B 0.035496f
C178 VTAIL.t3 B 0.035496f
C179 VTAIL.n46 B 0.194144f
C180 VTAIL.n47 B 0.243025f
C181 VP.n0 B 0.028152f
C182 VP.t5 B 0.084046f
C183 VP.n1 B 0.065824f
C184 VP.n2 B 0.028152f
C185 VP.n3 B 0.028152f
C186 VP.t2 B 0.084046f
C187 VP.t8 B 0.084046f
C188 VP.t0 B 0.084046f
C189 VP.n4 B 0.065824f
C190 VP.t7 B 0.091568f
C191 VP.n5 B 0.056088f
C192 VP.t9 B 0.084046f
C193 VP.n6 B 0.065043f
C194 VP.n7 B 0.006388f
C195 VP.n8 B 0.092397f
C196 VP.n9 B 0.028152f
C197 VP.n10 B 0.028152f
C198 VP.n11 B 0.006388f
C199 VP.n12 B 0.065043f
C200 VP.n13 B 0.063394f
C201 VP.n14 B 0.802396f
C202 VP.n15 B 0.83206f
C203 VP.t6 B 0.084046f
C204 VP.n16 B 0.063394f
C205 VP.t3 B 0.084046f
C206 VP.n17 B 0.065043f
C207 VP.n18 B 0.006388f
C208 VP.n19 B 0.028152f
C209 VP.n20 B 0.028152f
C210 VP.n21 B 0.028152f
C211 VP.n22 B 0.006388f
C212 VP.t1 B 0.084046f
C213 VP.n23 B 0.065043f
C214 VP.t4 B 0.084046f
C215 VP.n24 B 0.063394f
C216 VP.n25 B 0.021816f
.ends

