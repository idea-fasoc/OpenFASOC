* NGSPICE file created from diff_pair_sample_0759.ext - technology: sky130A

.subckt diff_pair_sample_0759 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X1 B.t11 B.t9 B.t10 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0 ps=0 w=3.75 l=0.16
X2 VTAIL.t14 VP.t1 VDD1.t6 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X3 VDD2.t7 VN.t0 VTAIL.t7 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X4 B.t8 B.t6 B.t7 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0 ps=0 w=3.75 l=0.16
X5 VDD2.t6 VN.t1 VTAIL.t0 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X6 VDD1.t5 VP.t2 VTAIL.t15 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X7 VDD2.t5 VN.t2 VTAIL.t1 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=1.78125 ps=8.45 w=3.75 l=0.16
X8 VTAIL.t6 VN.t3 VDD2.t4 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0.9375 ps=4.25 w=3.75 l=0.16
X9 B.t5 B.t3 B.t4 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0 ps=0 w=3.75 l=0.16
X10 VTAIL.t5 VN.t4 VDD2.t3 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0.9375 ps=4.25 w=3.75 l=0.16
X11 VDD2.t2 VN.t5 VTAIL.t2 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=1.78125 ps=8.45 w=3.75 l=0.16
X12 VTAIL.t11 VP.t3 VDD1.t4 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0.9375 ps=4.25 w=3.75 l=0.16
X13 B.t2 B.t0 B.t1 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0 ps=0 w=3.75 l=0.16
X14 VTAIL.t4 VN.t6 VDD2.t1 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X15 VTAIL.t12 VP.t4 VDD1.t3 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
X16 VDD1.t2 VP.t5 VTAIL.t8 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=1.78125 ps=8.45 w=3.75 l=0.16
X17 VTAIL.t13 VP.t6 VDD1.t1 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=1.78125 pd=8.45 as=0.9375 ps=4.25 w=3.75 l=0.16
X18 VDD1.t0 VP.t7 VTAIL.t9 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=1.78125 ps=8.45 w=3.75 l=0.16
X19 VTAIL.t3 VN.t7 VDD2.t0 w_n1630_n1718# sky130_fd_pr__pfet_01v8 ad=0.9375 pd=4.25 as=0.9375 ps=4.25 w=3.75 l=0.16
R0 VP.n17 VP.t5 797.217
R1 VP.n11 VP.t3 797.217
R2 VP.n4 VP.t6 797.217
R3 VP.n9 VP.t7 797.217
R4 VP.n16 VP.t1 762.163
R5 VP.n1 VP.t0 762.163
R6 VP.n3 VP.t2 762.163
R7 VP.n8 VP.t4 762.163
R8 VP.n5 VP.n4 161.489
R9 VP.n18 VP.n17 161.3
R10 VP.n6 VP.n5 161.3
R11 VP.n7 VP.n2 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n15 VP.n0 161.3
R14 VP.n14 VP.n13 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n15 VP.n14 73.0308
R17 VP.n7 VP.n6 73.0308
R18 VP.n11 VP.n1 61.346
R19 VP.n17 VP.n16 61.346
R20 VP.n4 VP.n3 61.346
R21 VP.n9 VP.n8 61.346
R22 VP.n12 VP.n10 34.0687
R23 VP.n14 VP.n1 11.6853
R24 VP.n16 VP.n15 11.6853
R25 VP.n6 VP.n3 11.6853
R26 VP.n8 VP.n7 11.6853
R27 VP.n5 VP.n2 0.189894
R28 VP.n10 VP.n2 0.189894
R29 VP.n13 VP.n12 0.189894
R30 VP.n13 VP.n0 0.189894
R31 VP.n18 VP.n0 0.189894
R32 VP VP.n18 0.0516364
R33 VTAIL.n11 VTAIL.t13 108.278
R34 VTAIL.n10 VTAIL.t1 108.278
R35 VTAIL.n7 VTAIL.t5 108.278
R36 VTAIL.n15 VTAIL.t2 108.278
R37 VTAIL.n2 VTAIL.t6 108.278
R38 VTAIL.n3 VTAIL.t8 108.278
R39 VTAIL.n6 VTAIL.t11 108.278
R40 VTAIL.n14 VTAIL.t9 108.278
R41 VTAIL.n13 VTAIL.n12 95.1441
R42 VTAIL.n9 VTAIL.n8 95.1441
R43 VTAIL.n1 VTAIL.n0 95.1439
R44 VTAIL.n5 VTAIL.n4 95.1439
R45 VTAIL.n15 VTAIL.n14 16.1686
R46 VTAIL.n7 VTAIL.n6 16.1686
R47 VTAIL.n0 VTAIL.t0 13.1338
R48 VTAIL.n0 VTAIL.t3 13.1338
R49 VTAIL.n4 VTAIL.t10 13.1338
R50 VTAIL.n4 VTAIL.t14 13.1338
R51 VTAIL.n12 VTAIL.t15 13.1338
R52 VTAIL.n12 VTAIL.t12 13.1338
R53 VTAIL.n8 VTAIL.t7 13.1338
R54 VTAIL.n8 VTAIL.t4 13.1338
R55 VTAIL.n9 VTAIL.n7 0.569465
R56 VTAIL.n10 VTAIL.n9 0.569465
R57 VTAIL.n13 VTAIL.n11 0.569465
R58 VTAIL.n14 VTAIL.n13 0.569465
R59 VTAIL.n6 VTAIL.n5 0.569465
R60 VTAIL.n5 VTAIL.n3 0.569465
R61 VTAIL.n2 VTAIL.n1 0.569465
R62 VTAIL VTAIL.n15 0.511276
R63 VTAIL.n11 VTAIL.n10 0.470328
R64 VTAIL.n3 VTAIL.n2 0.470328
R65 VTAIL VTAIL.n1 0.0586897
R66 VDD1 VDD1.n0 112.165
R67 VDD1.n3 VDD1.n2 112.052
R68 VDD1.n3 VDD1.n1 112.052
R69 VDD1.n5 VDD1.n4 111.823
R70 VDD1.n5 VDD1.n3 30.0914
R71 VDD1.n4 VDD1.t3 13.1338
R72 VDD1.n4 VDD1.t0 13.1338
R73 VDD1.n0 VDD1.t1 13.1338
R74 VDD1.n0 VDD1.t5 13.1338
R75 VDD1.n2 VDD1.t6 13.1338
R76 VDD1.n2 VDD1.t2 13.1338
R77 VDD1.n1 VDD1.t4 13.1338
R78 VDD1.n1 VDD1.t7 13.1338
R79 VDD1 VDD1.n5 0.226793
R80 B.n65 B.t3 816.256
R81 B.n73 B.t0 816.256
R82 B.n20 B.t9 816.256
R83 B.n28 B.t6 816.256
R84 B.n241 B.n240 585
R85 B.n242 B.n37 585
R86 B.n244 B.n243 585
R87 B.n245 B.n36 585
R88 B.n247 B.n246 585
R89 B.n248 B.n35 585
R90 B.n250 B.n249 585
R91 B.n251 B.n34 585
R92 B.n253 B.n252 585
R93 B.n254 B.n33 585
R94 B.n256 B.n255 585
R95 B.n257 B.n32 585
R96 B.n259 B.n258 585
R97 B.n260 B.n31 585
R98 B.n262 B.n261 585
R99 B.n263 B.n27 585
R100 B.n265 B.n264 585
R101 B.n266 B.n26 585
R102 B.n268 B.n267 585
R103 B.n269 B.n25 585
R104 B.n271 B.n270 585
R105 B.n272 B.n24 585
R106 B.n274 B.n273 585
R107 B.n275 B.n23 585
R108 B.n277 B.n276 585
R109 B.n278 B.n22 585
R110 B.n280 B.n279 585
R111 B.n282 B.n19 585
R112 B.n284 B.n283 585
R113 B.n285 B.n18 585
R114 B.n287 B.n286 585
R115 B.n288 B.n17 585
R116 B.n290 B.n289 585
R117 B.n291 B.n16 585
R118 B.n293 B.n292 585
R119 B.n294 B.n15 585
R120 B.n296 B.n295 585
R121 B.n297 B.n14 585
R122 B.n299 B.n298 585
R123 B.n300 B.n13 585
R124 B.n302 B.n301 585
R125 B.n303 B.n12 585
R126 B.n305 B.n304 585
R127 B.n306 B.n11 585
R128 B.n239 B.n38 585
R129 B.n238 B.n237 585
R130 B.n236 B.n39 585
R131 B.n235 B.n234 585
R132 B.n233 B.n40 585
R133 B.n232 B.n231 585
R134 B.n230 B.n41 585
R135 B.n229 B.n228 585
R136 B.n227 B.n42 585
R137 B.n226 B.n225 585
R138 B.n224 B.n43 585
R139 B.n223 B.n222 585
R140 B.n221 B.n44 585
R141 B.n220 B.n219 585
R142 B.n218 B.n45 585
R143 B.n217 B.n216 585
R144 B.n215 B.n46 585
R145 B.n214 B.n213 585
R146 B.n212 B.n47 585
R147 B.n211 B.n210 585
R148 B.n209 B.n48 585
R149 B.n208 B.n207 585
R150 B.n206 B.n49 585
R151 B.n205 B.n204 585
R152 B.n203 B.n50 585
R153 B.n202 B.n201 585
R154 B.n200 B.n51 585
R155 B.n199 B.n198 585
R156 B.n197 B.n52 585
R157 B.n196 B.n195 585
R158 B.n194 B.n53 585
R159 B.n193 B.n192 585
R160 B.n191 B.n54 585
R161 B.n190 B.n189 585
R162 B.n188 B.n55 585
R163 B.n187 B.n186 585
R164 B.n185 B.n56 585
R165 B.n118 B.n117 585
R166 B.n119 B.n82 585
R167 B.n121 B.n120 585
R168 B.n122 B.n81 585
R169 B.n124 B.n123 585
R170 B.n125 B.n80 585
R171 B.n127 B.n126 585
R172 B.n128 B.n79 585
R173 B.n130 B.n129 585
R174 B.n131 B.n78 585
R175 B.n133 B.n132 585
R176 B.n134 B.n77 585
R177 B.n136 B.n135 585
R178 B.n137 B.n76 585
R179 B.n139 B.n138 585
R180 B.n140 B.n75 585
R181 B.n142 B.n141 585
R182 B.n144 B.n72 585
R183 B.n146 B.n145 585
R184 B.n147 B.n71 585
R185 B.n149 B.n148 585
R186 B.n150 B.n70 585
R187 B.n152 B.n151 585
R188 B.n153 B.n69 585
R189 B.n155 B.n154 585
R190 B.n156 B.n68 585
R191 B.n158 B.n157 585
R192 B.n160 B.n159 585
R193 B.n161 B.n64 585
R194 B.n163 B.n162 585
R195 B.n164 B.n63 585
R196 B.n166 B.n165 585
R197 B.n167 B.n62 585
R198 B.n169 B.n168 585
R199 B.n170 B.n61 585
R200 B.n172 B.n171 585
R201 B.n173 B.n60 585
R202 B.n175 B.n174 585
R203 B.n176 B.n59 585
R204 B.n178 B.n177 585
R205 B.n179 B.n58 585
R206 B.n181 B.n180 585
R207 B.n182 B.n57 585
R208 B.n184 B.n183 585
R209 B.n116 B.n83 585
R210 B.n115 B.n114 585
R211 B.n113 B.n84 585
R212 B.n112 B.n111 585
R213 B.n110 B.n85 585
R214 B.n109 B.n108 585
R215 B.n107 B.n86 585
R216 B.n106 B.n105 585
R217 B.n104 B.n87 585
R218 B.n103 B.n102 585
R219 B.n101 B.n88 585
R220 B.n100 B.n99 585
R221 B.n98 B.n89 585
R222 B.n97 B.n96 585
R223 B.n95 B.n90 585
R224 B.n94 B.n93 585
R225 B.n92 B.n91 585
R226 B.n2 B.n0 585
R227 B.n333 B.n1 585
R228 B.n332 B.n331 585
R229 B.n330 B.n3 585
R230 B.n329 B.n328 585
R231 B.n327 B.n4 585
R232 B.n326 B.n325 585
R233 B.n324 B.n5 585
R234 B.n323 B.n322 585
R235 B.n321 B.n6 585
R236 B.n320 B.n319 585
R237 B.n318 B.n7 585
R238 B.n317 B.n316 585
R239 B.n315 B.n8 585
R240 B.n314 B.n313 585
R241 B.n312 B.n9 585
R242 B.n311 B.n310 585
R243 B.n309 B.n10 585
R244 B.n308 B.n307 585
R245 B.n335 B.n334 585
R246 B.n117 B.n116 492.5
R247 B.n308 B.n11 492.5
R248 B.n183 B.n56 492.5
R249 B.n241 B.n38 492.5
R250 B.n116 B.n115 163.367
R251 B.n115 B.n84 163.367
R252 B.n111 B.n84 163.367
R253 B.n111 B.n110 163.367
R254 B.n110 B.n109 163.367
R255 B.n109 B.n86 163.367
R256 B.n105 B.n86 163.367
R257 B.n105 B.n104 163.367
R258 B.n104 B.n103 163.367
R259 B.n103 B.n88 163.367
R260 B.n99 B.n88 163.367
R261 B.n99 B.n98 163.367
R262 B.n98 B.n97 163.367
R263 B.n97 B.n90 163.367
R264 B.n93 B.n90 163.367
R265 B.n93 B.n92 163.367
R266 B.n92 B.n2 163.367
R267 B.n334 B.n2 163.367
R268 B.n334 B.n333 163.367
R269 B.n333 B.n332 163.367
R270 B.n332 B.n3 163.367
R271 B.n328 B.n3 163.367
R272 B.n328 B.n327 163.367
R273 B.n327 B.n326 163.367
R274 B.n326 B.n5 163.367
R275 B.n322 B.n5 163.367
R276 B.n322 B.n321 163.367
R277 B.n321 B.n320 163.367
R278 B.n320 B.n7 163.367
R279 B.n316 B.n7 163.367
R280 B.n316 B.n315 163.367
R281 B.n315 B.n314 163.367
R282 B.n314 B.n9 163.367
R283 B.n310 B.n9 163.367
R284 B.n310 B.n309 163.367
R285 B.n309 B.n308 163.367
R286 B.n117 B.n82 163.367
R287 B.n121 B.n82 163.367
R288 B.n122 B.n121 163.367
R289 B.n123 B.n122 163.367
R290 B.n123 B.n80 163.367
R291 B.n127 B.n80 163.367
R292 B.n128 B.n127 163.367
R293 B.n129 B.n128 163.367
R294 B.n129 B.n78 163.367
R295 B.n133 B.n78 163.367
R296 B.n134 B.n133 163.367
R297 B.n135 B.n134 163.367
R298 B.n135 B.n76 163.367
R299 B.n139 B.n76 163.367
R300 B.n140 B.n139 163.367
R301 B.n141 B.n140 163.367
R302 B.n141 B.n72 163.367
R303 B.n146 B.n72 163.367
R304 B.n147 B.n146 163.367
R305 B.n148 B.n147 163.367
R306 B.n148 B.n70 163.367
R307 B.n152 B.n70 163.367
R308 B.n153 B.n152 163.367
R309 B.n154 B.n153 163.367
R310 B.n154 B.n68 163.367
R311 B.n158 B.n68 163.367
R312 B.n159 B.n158 163.367
R313 B.n159 B.n64 163.367
R314 B.n163 B.n64 163.367
R315 B.n164 B.n163 163.367
R316 B.n165 B.n164 163.367
R317 B.n165 B.n62 163.367
R318 B.n169 B.n62 163.367
R319 B.n170 B.n169 163.367
R320 B.n171 B.n170 163.367
R321 B.n171 B.n60 163.367
R322 B.n175 B.n60 163.367
R323 B.n176 B.n175 163.367
R324 B.n177 B.n176 163.367
R325 B.n177 B.n58 163.367
R326 B.n181 B.n58 163.367
R327 B.n182 B.n181 163.367
R328 B.n183 B.n182 163.367
R329 B.n187 B.n56 163.367
R330 B.n188 B.n187 163.367
R331 B.n189 B.n188 163.367
R332 B.n189 B.n54 163.367
R333 B.n193 B.n54 163.367
R334 B.n194 B.n193 163.367
R335 B.n195 B.n194 163.367
R336 B.n195 B.n52 163.367
R337 B.n199 B.n52 163.367
R338 B.n200 B.n199 163.367
R339 B.n201 B.n200 163.367
R340 B.n201 B.n50 163.367
R341 B.n205 B.n50 163.367
R342 B.n206 B.n205 163.367
R343 B.n207 B.n206 163.367
R344 B.n207 B.n48 163.367
R345 B.n211 B.n48 163.367
R346 B.n212 B.n211 163.367
R347 B.n213 B.n212 163.367
R348 B.n213 B.n46 163.367
R349 B.n217 B.n46 163.367
R350 B.n218 B.n217 163.367
R351 B.n219 B.n218 163.367
R352 B.n219 B.n44 163.367
R353 B.n223 B.n44 163.367
R354 B.n224 B.n223 163.367
R355 B.n225 B.n224 163.367
R356 B.n225 B.n42 163.367
R357 B.n229 B.n42 163.367
R358 B.n230 B.n229 163.367
R359 B.n231 B.n230 163.367
R360 B.n231 B.n40 163.367
R361 B.n235 B.n40 163.367
R362 B.n236 B.n235 163.367
R363 B.n237 B.n236 163.367
R364 B.n237 B.n38 163.367
R365 B.n304 B.n11 163.367
R366 B.n304 B.n303 163.367
R367 B.n303 B.n302 163.367
R368 B.n302 B.n13 163.367
R369 B.n298 B.n13 163.367
R370 B.n298 B.n297 163.367
R371 B.n297 B.n296 163.367
R372 B.n296 B.n15 163.367
R373 B.n292 B.n15 163.367
R374 B.n292 B.n291 163.367
R375 B.n291 B.n290 163.367
R376 B.n290 B.n17 163.367
R377 B.n286 B.n17 163.367
R378 B.n286 B.n285 163.367
R379 B.n285 B.n284 163.367
R380 B.n284 B.n19 163.367
R381 B.n279 B.n19 163.367
R382 B.n279 B.n278 163.367
R383 B.n278 B.n277 163.367
R384 B.n277 B.n23 163.367
R385 B.n273 B.n23 163.367
R386 B.n273 B.n272 163.367
R387 B.n272 B.n271 163.367
R388 B.n271 B.n25 163.367
R389 B.n267 B.n25 163.367
R390 B.n267 B.n266 163.367
R391 B.n266 B.n265 163.367
R392 B.n265 B.n27 163.367
R393 B.n261 B.n27 163.367
R394 B.n261 B.n260 163.367
R395 B.n260 B.n259 163.367
R396 B.n259 B.n32 163.367
R397 B.n255 B.n32 163.367
R398 B.n255 B.n254 163.367
R399 B.n254 B.n253 163.367
R400 B.n253 B.n34 163.367
R401 B.n249 B.n34 163.367
R402 B.n249 B.n248 163.367
R403 B.n248 B.n247 163.367
R404 B.n247 B.n36 163.367
R405 B.n243 B.n36 163.367
R406 B.n243 B.n242 163.367
R407 B.n242 B.n241 163.367
R408 B.n65 B.t5 139.734
R409 B.n28 B.t7 139.734
R410 B.n73 B.t2 139.731
R411 B.n20 B.t10 139.731
R412 B.n66 B.t4 126.934
R413 B.n29 B.t8 126.934
R414 B.n74 B.t1 126.931
R415 B.n21 B.t11 126.931
R416 B.n67 B.n66 59.5399
R417 B.n143 B.n74 59.5399
R418 B.n281 B.n21 59.5399
R419 B.n30 B.n29 59.5399
R420 B.n307 B.n306 32.0005
R421 B.n240 B.n239 32.0005
R422 B.n185 B.n184 32.0005
R423 B.n118 B.n83 32.0005
R424 B B.n335 18.0485
R425 B.n66 B.n65 12.8005
R426 B.n74 B.n73 12.8005
R427 B.n21 B.n20 12.8005
R428 B.n29 B.n28 12.8005
R429 B.n306 B.n305 10.6151
R430 B.n305 B.n12 10.6151
R431 B.n301 B.n12 10.6151
R432 B.n301 B.n300 10.6151
R433 B.n300 B.n299 10.6151
R434 B.n299 B.n14 10.6151
R435 B.n295 B.n14 10.6151
R436 B.n295 B.n294 10.6151
R437 B.n294 B.n293 10.6151
R438 B.n293 B.n16 10.6151
R439 B.n289 B.n16 10.6151
R440 B.n289 B.n288 10.6151
R441 B.n288 B.n287 10.6151
R442 B.n287 B.n18 10.6151
R443 B.n283 B.n18 10.6151
R444 B.n283 B.n282 10.6151
R445 B.n280 B.n22 10.6151
R446 B.n276 B.n22 10.6151
R447 B.n276 B.n275 10.6151
R448 B.n275 B.n274 10.6151
R449 B.n274 B.n24 10.6151
R450 B.n270 B.n24 10.6151
R451 B.n270 B.n269 10.6151
R452 B.n269 B.n268 10.6151
R453 B.n268 B.n26 10.6151
R454 B.n264 B.n263 10.6151
R455 B.n263 B.n262 10.6151
R456 B.n262 B.n31 10.6151
R457 B.n258 B.n31 10.6151
R458 B.n258 B.n257 10.6151
R459 B.n257 B.n256 10.6151
R460 B.n256 B.n33 10.6151
R461 B.n252 B.n33 10.6151
R462 B.n252 B.n251 10.6151
R463 B.n251 B.n250 10.6151
R464 B.n250 B.n35 10.6151
R465 B.n246 B.n35 10.6151
R466 B.n246 B.n245 10.6151
R467 B.n245 B.n244 10.6151
R468 B.n244 B.n37 10.6151
R469 B.n240 B.n37 10.6151
R470 B.n186 B.n185 10.6151
R471 B.n186 B.n55 10.6151
R472 B.n190 B.n55 10.6151
R473 B.n191 B.n190 10.6151
R474 B.n192 B.n191 10.6151
R475 B.n192 B.n53 10.6151
R476 B.n196 B.n53 10.6151
R477 B.n197 B.n196 10.6151
R478 B.n198 B.n197 10.6151
R479 B.n198 B.n51 10.6151
R480 B.n202 B.n51 10.6151
R481 B.n203 B.n202 10.6151
R482 B.n204 B.n203 10.6151
R483 B.n204 B.n49 10.6151
R484 B.n208 B.n49 10.6151
R485 B.n209 B.n208 10.6151
R486 B.n210 B.n209 10.6151
R487 B.n210 B.n47 10.6151
R488 B.n214 B.n47 10.6151
R489 B.n215 B.n214 10.6151
R490 B.n216 B.n215 10.6151
R491 B.n216 B.n45 10.6151
R492 B.n220 B.n45 10.6151
R493 B.n221 B.n220 10.6151
R494 B.n222 B.n221 10.6151
R495 B.n222 B.n43 10.6151
R496 B.n226 B.n43 10.6151
R497 B.n227 B.n226 10.6151
R498 B.n228 B.n227 10.6151
R499 B.n228 B.n41 10.6151
R500 B.n232 B.n41 10.6151
R501 B.n233 B.n232 10.6151
R502 B.n234 B.n233 10.6151
R503 B.n234 B.n39 10.6151
R504 B.n238 B.n39 10.6151
R505 B.n239 B.n238 10.6151
R506 B.n119 B.n118 10.6151
R507 B.n120 B.n119 10.6151
R508 B.n120 B.n81 10.6151
R509 B.n124 B.n81 10.6151
R510 B.n125 B.n124 10.6151
R511 B.n126 B.n125 10.6151
R512 B.n126 B.n79 10.6151
R513 B.n130 B.n79 10.6151
R514 B.n131 B.n130 10.6151
R515 B.n132 B.n131 10.6151
R516 B.n132 B.n77 10.6151
R517 B.n136 B.n77 10.6151
R518 B.n137 B.n136 10.6151
R519 B.n138 B.n137 10.6151
R520 B.n138 B.n75 10.6151
R521 B.n142 B.n75 10.6151
R522 B.n145 B.n144 10.6151
R523 B.n145 B.n71 10.6151
R524 B.n149 B.n71 10.6151
R525 B.n150 B.n149 10.6151
R526 B.n151 B.n150 10.6151
R527 B.n151 B.n69 10.6151
R528 B.n155 B.n69 10.6151
R529 B.n156 B.n155 10.6151
R530 B.n157 B.n156 10.6151
R531 B.n161 B.n160 10.6151
R532 B.n162 B.n161 10.6151
R533 B.n162 B.n63 10.6151
R534 B.n166 B.n63 10.6151
R535 B.n167 B.n166 10.6151
R536 B.n168 B.n167 10.6151
R537 B.n168 B.n61 10.6151
R538 B.n172 B.n61 10.6151
R539 B.n173 B.n172 10.6151
R540 B.n174 B.n173 10.6151
R541 B.n174 B.n59 10.6151
R542 B.n178 B.n59 10.6151
R543 B.n179 B.n178 10.6151
R544 B.n180 B.n179 10.6151
R545 B.n180 B.n57 10.6151
R546 B.n184 B.n57 10.6151
R547 B.n114 B.n83 10.6151
R548 B.n114 B.n113 10.6151
R549 B.n113 B.n112 10.6151
R550 B.n112 B.n85 10.6151
R551 B.n108 B.n85 10.6151
R552 B.n108 B.n107 10.6151
R553 B.n107 B.n106 10.6151
R554 B.n106 B.n87 10.6151
R555 B.n102 B.n87 10.6151
R556 B.n102 B.n101 10.6151
R557 B.n101 B.n100 10.6151
R558 B.n100 B.n89 10.6151
R559 B.n96 B.n89 10.6151
R560 B.n96 B.n95 10.6151
R561 B.n95 B.n94 10.6151
R562 B.n94 B.n91 10.6151
R563 B.n91 B.n0 10.6151
R564 B.n331 B.n1 10.6151
R565 B.n331 B.n330 10.6151
R566 B.n330 B.n329 10.6151
R567 B.n329 B.n4 10.6151
R568 B.n325 B.n4 10.6151
R569 B.n325 B.n324 10.6151
R570 B.n324 B.n323 10.6151
R571 B.n323 B.n6 10.6151
R572 B.n319 B.n6 10.6151
R573 B.n319 B.n318 10.6151
R574 B.n318 B.n317 10.6151
R575 B.n317 B.n8 10.6151
R576 B.n313 B.n8 10.6151
R577 B.n313 B.n312 10.6151
R578 B.n312 B.n311 10.6151
R579 B.n311 B.n10 10.6151
R580 B.n307 B.n10 10.6151
R581 B.n282 B.n281 9.36635
R582 B.n264 B.n30 9.36635
R583 B.n143 B.n142 9.36635
R584 B.n160 B.n67 9.36635
R585 B.n335 B.n0 2.81026
R586 B.n335 B.n1 2.81026
R587 B.n281 B.n280 1.24928
R588 B.n30 B.n26 1.24928
R589 B.n144 B.n143 1.24928
R590 B.n157 B.n67 1.24928
R591 VN.n7 VN.t5 797.217
R592 VN.n2 VN.t3 797.217
R593 VN.n16 VN.t4 797.217
R594 VN.n11 VN.t2 797.217
R595 VN.n6 VN.t7 762.163
R596 VN.n1 VN.t1 762.163
R597 VN.n15 VN.t0 762.163
R598 VN.n10 VN.t6 762.163
R599 VN.n12 VN.n11 161.489
R600 VN.n3 VN.n2 161.489
R601 VN.n8 VN.n7 161.3
R602 VN.n17 VN.n16 161.3
R603 VN.n14 VN.n9 161.3
R604 VN.n13 VN.n12 161.3
R605 VN.n5 VN.n0 161.3
R606 VN.n4 VN.n3 161.3
R607 VN.n5 VN.n4 73.0308
R608 VN.n14 VN.n13 73.0308
R609 VN.n2 VN.n1 61.346
R610 VN.n7 VN.n6 61.346
R611 VN.n16 VN.n15 61.346
R612 VN.n11 VN.n10 61.346
R613 VN VN.n17 34.4494
R614 VN.n4 VN.n1 11.6853
R615 VN.n6 VN.n5 11.6853
R616 VN.n15 VN.n14 11.6853
R617 VN.n13 VN.n10 11.6853
R618 VN.n17 VN.n9 0.189894
R619 VN.n12 VN.n9 0.189894
R620 VN.n3 VN.n0 0.189894
R621 VN.n8 VN.n0 0.189894
R622 VN VN.n8 0.0516364
R623 VDD2.n2 VDD2.n1 112.052
R624 VDD2.n2 VDD2.n0 112.052
R625 VDD2 VDD2.n5 112.049
R626 VDD2.n4 VDD2.n3 111.823
R627 VDD2.n4 VDD2.n2 29.5084
R628 VDD2.n5 VDD2.t1 13.1338
R629 VDD2.n5 VDD2.t5 13.1338
R630 VDD2.n3 VDD2.t3 13.1338
R631 VDD2.n3 VDD2.t7 13.1338
R632 VDD2.n1 VDD2.t0 13.1338
R633 VDD2.n1 VDD2.t2 13.1338
R634 VDD2.n0 VDD2.t4 13.1338
R635 VDD2.n0 VDD2.t6 13.1338
R636 VDD2 VDD2.n4 0.343172
C0 VN VTAIL 0.840228f
C1 VP VDD2 0.282351f
C2 B VDD1 0.738726f
C3 VDD2 VTAIL 6.44985f
C4 B w_n1630_n1718# 4.32422f
C5 VDD1 w_n1630_n1718# 0.928957f
C6 B VP 0.90732f
C7 VN VDD2 0.943401f
C8 VDD1 VP 1.07375f
C9 B VTAIL 1.42492f
C10 w_n1630_n1718# VP 2.65176f
C11 VDD1 VTAIL 6.41065f
C12 w_n1630_n1718# VTAIL 2.14637f
C13 B VN 0.576203f
C14 VDD1 VN 0.151549f
C15 VP VTAIL 0.854334f
C16 VN w_n1630_n1718# 2.44805f
C17 B VDD2 0.764041f
C18 VDD1 VDD2 0.644877f
C19 VN VP 3.35296f
C20 w_n1630_n1718# VDD2 0.948138f
C21 VDD2 VSUBS 0.833231f
C22 VDD1 VSUBS 1.051144f
C23 VTAIL VSUBS 0.353832f
C24 VN VSUBS 3.23069f
C25 VP VSUBS 0.721994f
C26 B VSUBS 1.619872f
C27 w_n1630_n1718# VSUBS 35.3058f
C28 VDD2.t4 VSUBS 0.106372f
C29 VDD2.t6 VSUBS 0.106372f
C30 VDD2.n0 VSUBS 0.474482f
C31 VDD2.t0 VSUBS 0.106372f
C32 VDD2.t2 VSUBS 0.106372f
C33 VDD2.n1 VSUBS 0.474482f
C34 VDD2.n2 VSUBS 1.65779f
C35 VDD2.t3 VSUBS 0.106372f
C36 VDD2.t7 VSUBS 0.106372f
C37 VDD2.n3 VSUBS 0.473666f
C38 VDD2.n4 VSUBS 1.5543f
C39 VDD2.t1 VSUBS 0.106372f
C40 VDD2.t5 VSUBS 0.106372f
C41 VDD2.n5 VSUBS 0.474466f
C42 VN.n0 VSUBS 0.064083f
C43 VN.t7 VSUBS 0.110724f
C44 VN.t1 VSUBS 0.110724f
C45 VN.n1 VSUBS 0.068221f
C46 VN.t3 VSUBS 0.11355f
C47 VN.n2 VSUBS 0.089106f
C48 VN.n3 VSUBS 0.133617f
C49 VN.n4 VSUBS 0.024419f
C50 VN.n5 VSUBS 0.024419f
C51 VN.n6 VSUBS 0.068221f
C52 VN.t5 VSUBS 0.11355f
C53 VN.n7 VSUBS 0.089024f
C54 VN.n8 VSUBS 0.049662f
C55 VN.n9 VSUBS 0.064083f
C56 VN.t4 VSUBS 0.11355f
C57 VN.t0 VSUBS 0.110724f
C58 VN.t6 VSUBS 0.110724f
C59 VN.n10 VSUBS 0.068221f
C60 VN.t2 VSUBS 0.11355f
C61 VN.n11 VSUBS 0.089106f
C62 VN.n12 VSUBS 0.133617f
C63 VN.n13 VSUBS 0.024419f
C64 VN.n14 VSUBS 0.024419f
C65 VN.n15 VSUBS 0.068221f
C66 VN.n16 VSUBS 0.089024f
C67 VN.n17 VSUBS 1.85417f
C68 B.n0 VSUBS 0.004792f
C69 B.n1 VSUBS 0.004792f
C70 B.n2 VSUBS 0.007578f
C71 B.n3 VSUBS 0.007578f
C72 B.n4 VSUBS 0.007578f
C73 B.n5 VSUBS 0.007578f
C74 B.n6 VSUBS 0.007578f
C75 B.n7 VSUBS 0.007578f
C76 B.n8 VSUBS 0.007578f
C77 B.n9 VSUBS 0.007578f
C78 B.n10 VSUBS 0.007578f
C79 B.n11 VSUBS 0.017687f
C80 B.n12 VSUBS 0.007578f
C81 B.n13 VSUBS 0.007578f
C82 B.n14 VSUBS 0.007578f
C83 B.n15 VSUBS 0.007578f
C84 B.n16 VSUBS 0.007578f
C85 B.n17 VSUBS 0.007578f
C86 B.n18 VSUBS 0.007578f
C87 B.n19 VSUBS 0.007578f
C88 B.t11 VSUBS 0.118235f
C89 B.t10 VSUBS 0.123391f
C90 B.t9 VSUBS 0.026517f
C91 B.n20 VSUBS 0.06907f
C92 B.n21 VSUBS 0.067093f
C93 B.n22 VSUBS 0.007578f
C94 B.n23 VSUBS 0.007578f
C95 B.n24 VSUBS 0.007578f
C96 B.n25 VSUBS 0.007578f
C97 B.n26 VSUBS 0.004235f
C98 B.n27 VSUBS 0.007578f
C99 B.t8 VSUBS 0.118235f
C100 B.t7 VSUBS 0.123391f
C101 B.t6 VSUBS 0.026517f
C102 B.n28 VSUBS 0.06907f
C103 B.n29 VSUBS 0.067092f
C104 B.n30 VSUBS 0.017558f
C105 B.n31 VSUBS 0.007578f
C106 B.n32 VSUBS 0.007578f
C107 B.n33 VSUBS 0.007578f
C108 B.n34 VSUBS 0.007578f
C109 B.n35 VSUBS 0.007578f
C110 B.n36 VSUBS 0.007578f
C111 B.n37 VSUBS 0.007578f
C112 B.n38 VSUBS 0.017308f
C113 B.n39 VSUBS 0.007578f
C114 B.n40 VSUBS 0.007578f
C115 B.n41 VSUBS 0.007578f
C116 B.n42 VSUBS 0.007578f
C117 B.n43 VSUBS 0.007578f
C118 B.n44 VSUBS 0.007578f
C119 B.n45 VSUBS 0.007578f
C120 B.n46 VSUBS 0.007578f
C121 B.n47 VSUBS 0.007578f
C122 B.n48 VSUBS 0.007578f
C123 B.n49 VSUBS 0.007578f
C124 B.n50 VSUBS 0.007578f
C125 B.n51 VSUBS 0.007578f
C126 B.n52 VSUBS 0.007578f
C127 B.n53 VSUBS 0.007578f
C128 B.n54 VSUBS 0.007578f
C129 B.n55 VSUBS 0.007578f
C130 B.n56 VSUBS 0.017308f
C131 B.n57 VSUBS 0.007578f
C132 B.n58 VSUBS 0.007578f
C133 B.n59 VSUBS 0.007578f
C134 B.n60 VSUBS 0.007578f
C135 B.n61 VSUBS 0.007578f
C136 B.n62 VSUBS 0.007578f
C137 B.n63 VSUBS 0.007578f
C138 B.n64 VSUBS 0.007578f
C139 B.t4 VSUBS 0.118235f
C140 B.t5 VSUBS 0.123391f
C141 B.t3 VSUBS 0.026517f
C142 B.n65 VSUBS 0.06907f
C143 B.n66 VSUBS 0.067092f
C144 B.n67 VSUBS 0.017558f
C145 B.n68 VSUBS 0.007578f
C146 B.n69 VSUBS 0.007578f
C147 B.n70 VSUBS 0.007578f
C148 B.n71 VSUBS 0.007578f
C149 B.n72 VSUBS 0.007578f
C150 B.t1 VSUBS 0.118235f
C151 B.t2 VSUBS 0.123391f
C152 B.t0 VSUBS 0.026517f
C153 B.n73 VSUBS 0.06907f
C154 B.n74 VSUBS 0.067093f
C155 B.n75 VSUBS 0.007578f
C156 B.n76 VSUBS 0.007578f
C157 B.n77 VSUBS 0.007578f
C158 B.n78 VSUBS 0.007578f
C159 B.n79 VSUBS 0.007578f
C160 B.n80 VSUBS 0.007578f
C161 B.n81 VSUBS 0.007578f
C162 B.n82 VSUBS 0.007578f
C163 B.n83 VSUBS 0.017308f
C164 B.n84 VSUBS 0.007578f
C165 B.n85 VSUBS 0.007578f
C166 B.n86 VSUBS 0.007578f
C167 B.n87 VSUBS 0.007578f
C168 B.n88 VSUBS 0.007578f
C169 B.n89 VSUBS 0.007578f
C170 B.n90 VSUBS 0.007578f
C171 B.n91 VSUBS 0.007578f
C172 B.n92 VSUBS 0.007578f
C173 B.n93 VSUBS 0.007578f
C174 B.n94 VSUBS 0.007578f
C175 B.n95 VSUBS 0.007578f
C176 B.n96 VSUBS 0.007578f
C177 B.n97 VSUBS 0.007578f
C178 B.n98 VSUBS 0.007578f
C179 B.n99 VSUBS 0.007578f
C180 B.n100 VSUBS 0.007578f
C181 B.n101 VSUBS 0.007578f
C182 B.n102 VSUBS 0.007578f
C183 B.n103 VSUBS 0.007578f
C184 B.n104 VSUBS 0.007578f
C185 B.n105 VSUBS 0.007578f
C186 B.n106 VSUBS 0.007578f
C187 B.n107 VSUBS 0.007578f
C188 B.n108 VSUBS 0.007578f
C189 B.n109 VSUBS 0.007578f
C190 B.n110 VSUBS 0.007578f
C191 B.n111 VSUBS 0.007578f
C192 B.n112 VSUBS 0.007578f
C193 B.n113 VSUBS 0.007578f
C194 B.n114 VSUBS 0.007578f
C195 B.n115 VSUBS 0.007578f
C196 B.n116 VSUBS 0.017308f
C197 B.n117 VSUBS 0.017687f
C198 B.n118 VSUBS 0.017687f
C199 B.n119 VSUBS 0.007578f
C200 B.n120 VSUBS 0.007578f
C201 B.n121 VSUBS 0.007578f
C202 B.n122 VSUBS 0.007578f
C203 B.n123 VSUBS 0.007578f
C204 B.n124 VSUBS 0.007578f
C205 B.n125 VSUBS 0.007578f
C206 B.n126 VSUBS 0.007578f
C207 B.n127 VSUBS 0.007578f
C208 B.n128 VSUBS 0.007578f
C209 B.n129 VSUBS 0.007578f
C210 B.n130 VSUBS 0.007578f
C211 B.n131 VSUBS 0.007578f
C212 B.n132 VSUBS 0.007578f
C213 B.n133 VSUBS 0.007578f
C214 B.n134 VSUBS 0.007578f
C215 B.n135 VSUBS 0.007578f
C216 B.n136 VSUBS 0.007578f
C217 B.n137 VSUBS 0.007578f
C218 B.n138 VSUBS 0.007578f
C219 B.n139 VSUBS 0.007578f
C220 B.n140 VSUBS 0.007578f
C221 B.n141 VSUBS 0.007578f
C222 B.n142 VSUBS 0.007133f
C223 B.n143 VSUBS 0.017558f
C224 B.n144 VSUBS 0.004235f
C225 B.n145 VSUBS 0.007578f
C226 B.n146 VSUBS 0.007578f
C227 B.n147 VSUBS 0.007578f
C228 B.n148 VSUBS 0.007578f
C229 B.n149 VSUBS 0.007578f
C230 B.n150 VSUBS 0.007578f
C231 B.n151 VSUBS 0.007578f
C232 B.n152 VSUBS 0.007578f
C233 B.n153 VSUBS 0.007578f
C234 B.n154 VSUBS 0.007578f
C235 B.n155 VSUBS 0.007578f
C236 B.n156 VSUBS 0.007578f
C237 B.n157 VSUBS 0.004235f
C238 B.n158 VSUBS 0.007578f
C239 B.n159 VSUBS 0.007578f
C240 B.n160 VSUBS 0.007133f
C241 B.n161 VSUBS 0.007578f
C242 B.n162 VSUBS 0.007578f
C243 B.n163 VSUBS 0.007578f
C244 B.n164 VSUBS 0.007578f
C245 B.n165 VSUBS 0.007578f
C246 B.n166 VSUBS 0.007578f
C247 B.n167 VSUBS 0.007578f
C248 B.n168 VSUBS 0.007578f
C249 B.n169 VSUBS 0.007578f
C250 B.n170 VSUBS 0.007578f
C251 B.n171 VSUBS 0.007578f
C252 B.n172 VSUBS 0.007578f
C253 B.n173 VSUBS 0.007578f
C254 B.n174 VSUBS 0.007578f
C255 B.n175 VSUBS 0.007578f
C256 B.n176 VSUBS 0.007578f
C257 B.n177 VSUBS 0.007578f
C258 B.n178 VSUBS 0.007578f
C259 B.n179 VSUBS 0.007578f
C260 B.n180 VSUBS 0.007578f
C261 B.n181 VSUBS 0.007578f
C262 B.n182 VSUBS 0.007578f
C263 B.n183 VSUBS 0.017687f
C264 B.n184 VSUBS 0.017687f
C265 B.n185 VSUBS 0.017308f
C266 B.n186 VSUBS 0.007578f
C267 B.n187 VSUBS 0.007578f
C268 B.n188 VSUBS 0.007578f
C269 B.n189 VSUBS 0.007578f
C270 B.n190 VSUBS 0.007578f
C271 B.n191 VSUBS 0.007578f
C272 B.n192 VSUBS 0.007578f
C273 B.n193 VSUBS 0.007578f
C274 B.n194 VSUBS 0.007578f
C275 B.n195 VSUBS 0.007578f
C276 B.n196 VSUBS 0.007578f
C277 B.n197 VSUBS 0.007578f
C278 B.n198 VSUBS 0.007578f
C279 B.n199 VSUBS 0.007578f
C280 B.n200 VSUBS 0.007578f
C281 B.n201 VSUBS 0.007578f
C282 B.n202 VSUBS 0.007578f
C283 B.n203 VSUBS 0.007578f
C284 B.n204 VSUBS 0.007578f
C285 B.n205 VSUBS 0.007578f
C286 B.n206 VSUBS 0.007578f
C287 B.n207 VSUBS 0.007578f
C288 B.n208 VSUBS 0.007578f
C289 B.n209 VSUBS 0.007578f
C290 B.n210 VSUBS 0.007578f
C291 B.n211 VSUBS 0.007578f
C292 B.n212 VSUBS 0.007578f
C293 B.n213 VSUBS 0.007578f
C294 B.n214 VSUBS 0.007578f
C295 B.n215 VSUBS 0.007578f
C296 B.n216 VSUBS 0.007578f
C297 B.n217 VSUBS 0.007578f
C298 B.n218 VSUBS 0.007578f
C299 B.n219 VSUBS 0.007578f
C300 B.n220 VSUBS 0.007578f
C301 B.n221 VSUBS 0.007578f
C302 B.n222 VSUBS 0.007578f
C303 B.n223 VSUBS 0.007578f
C304 B.n224 VSUBS 0.007578f
C305 B.n225 VSUBS 0.007578f
C306 B.n226 VSUBS 0.007578f
C307 B.n227 VSUBS 0.007578f
C308 B.n228 VSUBS 0.007578f
C309 B.n229 VSUBS 0.007578f
C310 B.n230 VSUBS 0.007578f
C311 B.n231 VSUBS 0.007578f
C312 B.n232 VSUBS 0.007578f
C313 B.n233 VSUBS 0.007578f
C314 B.n234 VSUBS 0.007578f
C315 B.n235 VSUBS 0.007578f
C316 B.n236 VSUBS 0.007578f
C317 B.n237 VSUBS 0.007578f
C318 B.n238 VSUBS 0.007578f
C319 B.n239 VSUBS 0.018222f
C320 B.n240 VSUBS 0.016773f
C321 B.n241 VSUBS 0.017687f
C322 B.n242 VSUBS 0.007578f
C323 B.n243 VSUBS 0.007578f
C324 B.n244 VSUBS 0.007578f
C325 B.n245 VSUBS 0.007578f
C326 B.n246 VSUBS 0.007578f
C327 B.n247 VSUBS 0.007578f
C328 B.n248 VSUBS 0.007578f
C329 B.n249 VSUBS 0.007578f
C330 B.n250 VSUBS 0.007578f
C331 B.n251 VSUBS 0.007578f
C332 B.n252 VSUBS 0.007578f
C333 B.n253 VSUBS 0.007578f
C334 B.n254 VSUBS 0.007578f
C335 B.n255 VSUBS 0.007578f
C336 B.n256 VSUBS 0.007578f
C337 B.n257 VSUBS 0.007578f
C338 B.n258 VSUBS 0.007578f
C339 B.n259 VSUBS 0.007578f
C340 B.n260 VSUBS 0.007578f
C341 B.n261 VSUBS 0.007578f
C342 B.n262 VSUBS 0.007578f
C343 B.n263 VSUBS 0.007578f
C344 B.n264 VSUBS 0.007133f
C345 B.n265 VSUBS 0.007578f
C346 B.n266 VSUBS 0.007578f
C347 B.n267 VSUBS 0.007578f
C348 B.n268 VSUBS 0.007578f
C349 B.n269 VSUBS 0.007578f
C350 B.n270 VSUBS 0.007578f
C351 B.n271 VSUBS 0.007578f
C352 B.n272 VSUBS 0.007578f
C353 B.n273 VSUBS 0.007578f
C354 B.n274 VSUBS 0.007578f
C355 B.n275 VSUBS 0.007578f
C356 B.n276 VSUBS 0.007578f
C357 B.n277 VSUBS 0.007578f
C358 B.n278 VSUBS 0.007578f
C359 B.n279 VSUBS 0.007578f
C360 B.n280 VSUBS 0.004235f
C361 B.n281 VSUBS 0.017558f
C362 B.n282 VSUBS 0.007133f
C363 B.n283 VSUBS 0.007578f
C364 B.n284 VSUBS 0.007578f
C365 B.n285 VSUBS 0.007578f
C366 B.n286 VSUBS 0.007578f
C367 B.n287 VSUBS 0.007578f
C368 B.n288 VSUBS 0.007578f
C369 B.n289 VSUBS 0.007578f
C370 B.n290 VSUBS 0.007578f
C371 B.n291 VSUBS 0.007578f
C372 B.n292 VSUBS 0.007578f
C373 B.n293 VSUBS 0.007578f
C374 B.n294 VSUBS 0.007578f
C375 B.n295 VSUBS 0.007578f
C376 B.n296 VSUBS 0.007578f
C377 B.n297 VSUBS 0.007578f
C378 B.n298 VSUBS 0.007578f
C379 B.n299 VSUBS 0.007578f
C380 B.n300 VSUBS 0.007578f
C381 B.n301 VSUBS 0.007578f
C382 B.n302 VSUBS 0.007578f
C383 B.n303 VSUBS 0.007578f
C384 B.n304 VSUBS 0.007578f
C385 B.n305 VSUBS 0.007578f
C386 B.n306 VSUBS 0.017687f
C387 B.n307 VSUBS 0.017308f
C388 B.n308 VSUBS 0.017308f
C389 B.n309 VSUBS 0.007578f
C390 B.n310 VSUBS 0.007578f
C391 B.n311 VSUBS 0.007578f
C392 B.n312 VSUBS 0.007578f
C393 B.n313 VSUBS 0.007578f
C394 B.n314 VSUBS 0.007578f
C395 B.n315 VSUBS 0.007578f
C396 B.n316 VSUBS 0.007578f
C397 B.n317 VSUBS 0.007578f
C398 B.n318 VSUBS 0.007578f
C399 B.n319 VSUBS 0.007578f
C400 B.n320 VSUBS 0.007578f
C401 B.n321 VSUBS 0.007578f
C402 B.n322 VSUBS 0.007578f
C403 B.n323 VSUBS 0.007578f
C404 B.n324 VSUBS 0.007578f
C405 B.n325 VSUBS 0.007578f
C406 B.n326 VSUBS 0.007578f
C407 B.n327 VSUBS 0.007578f
C408 B.n328 VSUBS 0.007578f
C409 B.n329 VSUBS 0.007578f
C410 B.n330 VSUBS 0.007578f
C411 B.n331 VSUBS 0.007578f
C412 B.n332 VSUBS 0.007578f
C413 B.n333 VSUBS 0.007578f
C414 B.n334 VSUBS 0.007578f
C415 B.n335 VSUBS 0.01716f
C416 VDD1.t1 VSUBS 0.104937f
C417 VDD1.t5 VSUBS 0.104937f
C418 VDD1.n0 VSUBS 0.468501f
C419 VDD1.t4 VSUBS 0.104937f
C420 VDD1.t7 VSUBS 0.104937f
C421 VDD1.n1 VSUBS 0.468082f
C422 VDD1.t6 VSUBS 0.104937f
C423 VDD1.t2 VSUBS 0.104937f
C424 VDD1.n2 VSUBS 0.468082f
C425 VDD1.n3 VSUBS 1.68582f
C426 VDD1.t3 VSUBS 0.104937f
C427 VDD1.t0 VSUBS 0.104937f
C428 VDD1.n4 VSUBS 0.467275f
C429 VDD1.n5 VSUBS 1.56049f
C430 VTAIL.t0 VSUBS 0.10644f
C431 VTAIL.t3 VSUBS 0.10644f
C432 VTAIL.n0 VSUBS 0.417406f
C433 VTAIL.n1 VSUBS 0.399425f
C434 VTAIL.t6 VSUBS 0.548041f
C435 VTAIL.n2 VSUBS 0.491826f
C436 VTAIL.t8 VSUBS 0.548041f
C437 VTAIL.n3 VSUBS 0.491826f
C438 VTAIL.t10 VSUBS 0.10644f
C439 VTAIL.t14 VSUBS 0.10644f
C440 VTAIL.n4 VSUBS 0.417406f
C441 VTAIL.n5 VSUBS 0.438442f
C442 VTAIL.t11 VSUBS 0.548041f
C443 VTAIL.n6 VSUBS 1.06836f
C444 VTAIL.t5 VSUBS 0.548043f
C445 VTAIL.n7 VSUBS 1.06836f
C446 VTAIL.t7 VSUBS 0.10644f
C447 VTAIL.t4 VSUBS 0.10644f
C448 VTAIL.n8 VSUBS 0.417409f
C449 VTAIL.n9 VSUBS 0.438439f
C450 VTAIL.t1 VSUBS 0.548043f
C451 VTAIL.n10 VSUBS 0.491824f
C452 VTAIL.t13 VSUBS 0.548043f
C453 VTAIL.n11 VSUBS 0.491824f
C454 VTAIL.t15 VSUBS 0.10644f
C455 VTAIL.t12 VSUBS 0.10644f
C456 VTAIL.n12 VSUBS 0.417409f
C457 VTAIL.n13 VSUBS 0.438439f
C458 VTAIL.t9 VSUBS 0.548041f
C459 VTAIL.n14 VSUBS 1.06836f
C460 VTAIL.t2 VSUBS 0.548041f
C461 VTAIL.n15 VSUBS 1.06392f
C462 VP.n0 VSUBS 0.068461f
C463 VP.t1 VSUBS 0.118289f
C464 VP.t0 VSUBS 0.118289f
C465 VP.n1 VSUBS 0.072882f
C466 VP.n2 VSUBS 0.068461f
C467 VP.t4 VSUBS 0.118289f
C468 VP.t2 VSUBS 0.118289f
C469 VP.n3 VSUBS 0.072882f
C470 VP.t6 VSUBS 0.121308f
C471 VP.n4 VSUBS 0.095193f
C472 VP.n5 VSUBS 0.142745f
C473 VP.n6 VSUBS 0.026088f
C474 VP.n7 VSUBS 0.026088f
C475 VP.n8 VSUBS 0.072882f
C476 VP.t7 VSUBS 0.121308f
C477 VP.n9 VSUBS 0.095106f
C478 VP.n10 VSUBS 1.93525f
C479 VP.t3 VSUBS 0.121308f
C480 VP.n11 VSUBS 0.095106f
C481 VP.n12 VSUBS 2.00748f
C482 VP.n13 VSUBS 0.068461f
C483 VP.n14 VSUBS 0.026088f
C484 VP.n15 VSUBS 0.026088f
C485 VP.n16 VSUBS 0.072882f
C486 VP.t5 VSUBS 0.121308f
C487 VP.n17 VSUBS 0.095106f
C488 VP.n18 VSUBS 0.053055f
.ends

