* NGSPICE file created from diff_pair_sample_1483.ext - technology: sky130A

.subckt diff_pair_sample_1483 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=2.2902 pd=14.21 as=5.4132 ps=28.54 w=13.88 l=1.96
X1 B.t11 B.t9 B.t10 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=0 ps=0 w=13.88 l=1.96
X2 B.t8 B.t6 B.t7 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=0 ps=0 w=13.88 l=1.96
X3 VTAIL.t5 VN.t1 VDD2.t2 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=2.2902 ps=14.21 w=13.88 l=1.96
X4 B.t5 B.t3 B.t4 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=0 ps=0 w=13.88 l=1.96
X5 VDD2.t1 VN.t2 VTAIL.t4 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=2.2902 pd=14.21 as=5.4132 ps=28.54 w=13.88 l=1.96
X6 VTAIL.t7 VN.t3 VDD2.t0 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=2.2902 ps=14.21 w=13.88 l=1.96
X7 VDD1.t3 VP.t0 VTAIL.t2 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=2.2902 pd=14.21 as=5.4132 ps=28.54 w=13.88 l=1.96
X8 B.t2 B.t0 B.t1 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=0 ps=0 w=13.88 l=1.96
X9 VTAIL.t3 VP.t1 VDD1.t2 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=2.2902 ps=14.21 w=13.88 l=1.96
X10 VDD1.t1 VP.t2 VTAIL.t0 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=2.2902 pd=14.21 as=5.4132 ps=28.54 w=13.88 l=1.96
X11 VTAIL.t1 VP.t3 VDD1.t0 w_n2344_n3744# sky130_fd_pr__pfet_01v8 ad=5.4132 pd=28.54 as=2.2902 ps=14.21 w=13.88 l=1.96
R0 VN.n0 VN.t1 205.95
R1 VN.n1 VN.t2 205.95
R2 VN.n0 VN.t0 205.424
R3 VN.n1 VN.t3 205.424
R4 VN VN.n1 53.4356
R5 VN VN.n0 7.44692
R6 VTAIL.n6 VTAIL.t2 56.8345
R7 VTAIL.n5 VTAIL.t3 56.8344
R8 VTAIL.n4 VTAIL.t4 56.8344
R9 VTAIL.n3 VTAIL.t7 56.8344
R10 VTAIL.n7 VTAIL.t6 56.8343
R11 VTAIL.n0 VTAIL.t5 56.8343
R12 VTAIL.n1 VTAIL.t0 56.8343
R13 VTAIL.n2 VTAIL.t1 56.8343
R14 VTAIL.n7 VTAIL.n6 26.3065
R15 VTAIL.n3 VTAIL.n2 26.3065
R16 VTAIL.n4 VTAIL.n3 1.97464
R17 VTAIL.n6 VTAIL.n5 1.97464
R18 VTAIL.n2 VTAIL.n1 1.97464
R19 VTAIL VTAIL.n0 1.04576
R20 VTAIL VTAIL.n7 0.929379
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 112.775
R24 VDD2.n2 VDD2.n1 71.1714
R25 VDD2.n1 VDD2.t0 2.34236
R26 VDD2.n1 VDD2.t1 2.34236
R27 VDD2.n0 VDD2.t2 2.34236
R28 VDD2.n0 VDD2.t3 2.34236
R29 VDD2 VDD2.n2 0.0586897
R30 B.n369 B.n102 585
R31 B.n368 B.n367 585
R32 B.n366 B.n103 585
R33 B.n365 B.n364 585
R34 B.n363 B.n104 585
R35 B.n362 B.n361 585
R36 B.n360 B.n105 585
R37 B.n359 B.n358 585
R38 B.n357 B.n106 585
R39 B.n356 B.n355 585
R40 B.n354 B.n107 585
R41 B.n353 B.n352 585
R42 B.n351 B.n108 585
R43 B.n350 B.n349 585
R44 B.n348 B.n109 585
R45 B.n347 B.n346 585
R46 B.n345 B.n110 585
R47 B.n344 B.n343 585
R48 B.n342 B.n111 585
R49 B.n341 B.n340 585
R50 B.n339 B.n112 585
R51 B.n338 B.n337 585
R52 B.n336 B.n113 585
R53 B.n335 B.n334 585
R54 B.n333 B.n114 585
R55 B.n332 B.n331 585
R56 B.n330 B.n115 585
R57 B.n329 B.n328 585
R58 B.n327 B.n116 585
R59 B.n326 B.n325 585
R60 B.n324 B.n117 585
R61 B.n323 B.n322 585
R62 B.n321 B.n118 585
R63 B.n320 B.n319 585
R64 B.n318 B.n119 585
R65 B.n317 B.n316 585
R66 B.n315 B.n120 585
R67 B.n314 B.n313 585
R68 B.n312 B.n121 585
R69 B.n311 B.n310 585
R70 B.n309 B.n122 585
R71 B.n308 B.n307 585
R72 B.n306 B.n123 585
R73 B.n305 B.n304 585
R74 B.n303 B.n124 585
R75 B.n302 B.n301 585
R76 B.n300 B.n125 585
R77 B.n299 B.n298 585
R78 B.n294 B.n126 585
R79 B.n293 B.n292 585
R80 B.n291 B.n127 585
R81 B.n290 B.n289 585
R82 B.n288 B.n128 585
R83 B.n287 B.n286 585
R84 B.n285 B.n129 585
R85 B.n284 B.n283 585
R86 B.n282 B.n130 585
R87 B.n280 B.n279 585
R88 B.n278 B.n133 585
R89 B.n277 B.n276 585
R90 B.n275 B.n134 585
R91 B.n274 B.n273 585
R92 B.n272 B.n135 585
R93 B.n271 B.n270 585
R94 B.n269 B.n136 585
R95 B.n268 B.n267 585
R96 B.n266 B.n137 585
R97 B.n265 B.n264 585
R98 B.n263 B.n138 585
R99 B.n262 B.n261 585
R100 B.n260 B.n139 585
R101 B.n259 B.n258 585
R102 B.n257 B.n140 585
R103 B.n256 B.n255 585
R104 B.n254 B.n141 585
R105 B.n253 B.n252 585
R106 B.n251 B.n142 585
R107 B.n250 B.n249 585
R108 B.n248 B.n143 585
R109 B.n247 B.n246 585
R110 B.n245 B.n144 585
R111 B.n244 B.n243 585
R112 B.n242 B.n145 585
R113 B.n241 B.n240 585
R114 B.n239 B.n146 585
R115 B.n238 B.n237 585
R116 B.n236 B.n147 585
R117 B.n235 B.n234 585
R118 B.n233 B.n148 585
R119 B.n232 B.n231 585
R120 B.n230 B.n149 585
R121 B.n229 B.n228 585
R122 B.n227 B.n150 585
R123 B.n226 B.n225 585
R124 B.n224 B.n151 585
R125 B.n223 B.n222 585
R126 B.n221 B.n152 585
R127 B.n220 B.n219 585
R128 B.n218 B.n153 585
R129 B.n217 B.n216 585
R130 B.n215 B.n154 585
R131 B.n214 B.n213 585
R132 B.n212 B.n155 585
R133 B.n211 B.n210 585
R134 B.n371 B.n370 585
R135 B.n372 B.n101 585
R136 B.n374 B.n373 585
R137 B.n375 B.n100 585
R138 B.n377 B.n376 585
R139 B.n378 B.n99 585
R140 B.n380 B.n379 585
R141 B.n381 B.n98 585
R142 B.n383 B.n382 585
R143 B.n384 B.n97 585
R144 B.n386 B.n385 585
R145 B.n387 B.n96 585
R146 B.n389 B.n388 585
R147 B.n390 B.n95 585
R148 B.n392 B.n391 585
R149 B.n393 B.n94 585
R150 B.n395 B.n394 585
R151 B.n396 B.n93 585
R152 B.n398 B.n397 585
R153 B.n399 B.n92 585
R154 B.n401 B.n400 585
R155 B.n402 B.n91 585
R156 B.n404 B.n403 585
R157 B.n405 B.n90 585
R158 B.n407 B.n406 585
R159 B.n408 B.n89 585
R160 B.n410 B.n409 585
R161 B.n411 B.n88 585
R162 B.n413 B.n412 585
R163 B.n414 B.n87 585
R164 B.n416 B.n415 585
R165 B.n417 B.n86 585
R166 B.n419 B.n418 585
R167 B.n420 B.n85 585
R168 B.n422 B.n421 585
R169 B.n423 B.n84 585
R170 B.n425 B.n424 585
R171 B.n426 B.n83 585
R172 B.n428 B.n427 585
R173 B.n429 B.n82 585
R174 B.n431 B.n430 585
R175 B.n432 B.n81 585
R176 B.n434 B.n433 585
R177 B.n435 B.n80 585
R178 B.n437 B.n436 585
R179 B.n438 B.n79 585
R180 B.n440 B.n439 585
R181 B.n441 B.n78 585
R182 B.n443 B.n442 585
R183 B.n444 B.n77 585
R184 B.n446 B.n445 585
R185 B.n447 B.n76 585
R186 B.n449 B.n448 585
R187 B.n450 B.n75 585
R188 B.n452 B.n451 585
R189 B.n453 B.n74 585
R190 B.n455 B.n454 585
R191 B.n456 B.n73 585
R192 B.n613 B.n16 585
R193 B.n612 B.n611 585
R194 B.n610 B.n17 585
R195 B.n609 B.n608 585
R196 B.n607 B.n18 585
R197 B.n606 B.n605 585
R198 B.n604 B.n19 585
R199 B.n603 B.n602 585
R200 B.n601 B.n20 585
R201 B.n600 B.n599 585
R202 B.n598 B.n21 585
R203 B.n597 B.n596 585
R204 B.n595 B.n22 585
R205 B.n594 B.n593 585
R206 B.n592 B.n23 585
R207 B.n591 B.n590 585
R208 B.n589 B.n24 585
R209 B.n588 B.n587 585
R210 B.n586 B.n25 585
R211 B.n585 B.n584 585
R212 B.n583 B.n26 585
R213 B.n582 B.n581 585
R214 B.n580 B.n27 585
R215 B.n579 B.n578 585
R216 B.n577 B.n28 585
R217 B.n576 B.n575 585
R218 B.n574 B.n29 585
R219 B.n573 B.n572 585
R220 B.n571 B.n30 585
R221 B.n570 B.n569 585
R222 B.n568 B.n31 585
R223 B.n567 B.n566 585
R224 B.n565 B.n32 585
R225 B.n564 B.n563 585
R226 B.n562 B.n33 585
R227 B.n561 B.n560 585
R228 B.n559 B.n34 585
R229 B.n558 B.n557 585
R230 B.n556 B.n35 585
R231 B.n555 B.n554 585
R232 B.n553 B.n36 585
R233 B.n552 B.n551 585
R234 B.n550 B.n37 585
R235 B.n549 B.n548 585
R236 B.n547 B.n38 585
R237 B.n546 B.n545 585
R238 B.n544 B.n39 585
R239 B.n542 B.n541 585
R240 B.n540 B.n42 585
R241 B.n539 B.n538 585
R242 B.n537 B.n43 585
R243 B.n536 B.n535 585
R244 B.n534 B.n44 585
R245 B.n533 B.n532 585
R246 B.n531 B.n45 585
R247 B.n530 B.n529 585
R248 B.n528 B.n46 585
R249 B.n527 B.n526 585
R250 B.n525 B.n47 585
R251 B.n524 B.n523 585
R252 B.n522 B.n51 585
R253 B.n521 B.n520 585
R254 B.n519 B.n52 585
R255 B.n518 B.n517 585
R256 B.n516 B.n53 585
R257 B.n515 B.n514 585
R258 B.n513 B.n54 585
R259 B.n512 B.n511 585
R260 B.n510 B.n55 585
R261 B.n509 B.n508 585
R262 B.n507 B.n56 585
R263 B.n506 B.n505 585
R264 B.n504 B.n57 585
R265 B.n503 B.n502 585
R266 B.n501 B.n58 585
R267 B.n500 B.n499 585
R268 B.n498 B.n59 585
R269 B.n497 B.n496 585
R270 B.n495 B.n60 585
R271 B.n494 B.n493 585
R272 B.n492 B.n61 585
R273 B.n491 B.n490 585
R274 B.n489 B.n62 585
R275 B.n488 B.n487 585
R276 B.n486 B.n63 585
R277 B.n485 B.n484 585
R278 B.n483 B.n64 585
R279 B.n482 B.n481 585
R280 B.n480 B.n65 585
R281 B.n479 B.n478 585
R282 B.n477 B.n66 585
R283 B.n476 B.n475 585
R284 B.n474 B.n67 585
R285 B.n473 B.n472 585
R286 B.n471 B.n68 585
R287 B.n470 B.n469 585
R288 B.n468 B.n69 585
R289 B.n467 B.n466 585
R290 B.n465 B.n70 585
R291 B.n464 B.n463 585
R292 B.n462 B.n71 585
R293 B.n461 B.n460 585
R294 B.n459 B.n72 585
R295 B.n458 B.n457 585
R296 B.n615 B.n614 585
R297 B.n616 B.n15 585
R298 B.n618 B.n617 585
R299 B.n619 B.n14 585
R300 B.n621 B.n620 585
R301 B.n622 B.n13 585
R302 B.n624 B.n623 585
R303 B.n625 B.n12 585
R304 B.n627 B.n626 585
R305 B.n628 B.n11 585
R306 B.n630 B.n629 585
R307 B.n631 B.n10 585
R308 B.n633 B.n632 585
R309 B.n634 B.n9 585
R310 B.n636 B.n635 585
R311 B.n637 B.n8 585
R312 B.n639 B.n638 585
R313 B.n640 B.n7 585
R314 B.n642 B.n641 585
R315 B.n643 B.n6 585
R316 B.n645 B.n644 585
R317 B.n646 B.n5 585
R318 B.n648 B.n647 585
R319 B.n649 B.n4 585
R320 B.n651 B.n650 585
R321 B.n652 B.n3 585
R322 B.n654 B.n653 585
R323 B.n655 B.n0 585
R324 B.n2 B.n1 585
R325 B.n170 B.n169 585
R326 B.n172 B.n171 585
R327 B.n173 B.n168 585
R328 B.n175 B.n174 585
R329 B.n176 B.n167 585
R330 B.n178 B.n177 585
R331 B.n179 B.n166 585
R332 B.n181 B.n180 585
R333 B.n182 B.n165 585
R334 B.n184 B.n183 585
R335 B.n185 B.n164 585
R336 B.n187 B.n186 585
R337 B.n188 B.n163 585
R338 B.n190 B.n189 585
R339 B.n191 B.n162 585
R340 B.n193 B.n192 585
R341 B.n194 B.n161 585
R342 B.n196 B.n195 585
R343 B.n197 B.n160 585
R344 B.n199 B.n198 585
R345 B.n200 B.n159 585
R346 B.n202 B.n201 585
R347 B.n203 B.n158 585
R348 B.n205 B.n204 585
R349 B.n206 B.n157 585
R350 B.n208 B.n207 585
R351 B.n209 B.n156 585
R352 B.n211 B.n156 458.866
R353 B.n371 B.n102 458.866
R354 B.n457 B.n456 458.866
R355 B.n614 B.n613 458.866
R356 B.n131 B.t6 377.49
R357 B.n295 B.t3 377.49
R358 B.n48 B.t0 377.49
R359 B.n40 B.t9 377.49
R360 B.n657 B.n656 256.663
R361 B.n656 B.n655 235.042
R362 B.n656 B.n2 235.042
R363 B.n212 B.n211 163.367
R364 B.n213 B.n212 163.367
R365 B.n213 B.n154 163.367
R366 B.n217 B.n154 163.367
R367 B.n218 B.n217 163.367
R368 B.n219 B.n218 163.367
R369 B.n219 B.n152 163.367
R370 B.n223 B.n152 163.367
R371 B.n224 B.n223 163.367
R372 B.n225 B.n224 163.367
R373 B.n225 B.n150 163.367
R374 B.n229 B.n150 163.367
R375 B.n230 B.n229 163.367
R376 B.n231 B.n230 163.367
R377 B.n231 B.n148 163.367
R378 B.n235 B.n148 163.367
R379 B.n236 B.n235 163.367
R380 B.n237 B.n236 163.367
R381 B.n237 B.n146 163.367
R382 B.n241 B.n146 163.367
R383 B.n242 B.n241 163.367
R384 B.n243 B.n242 163.367
R385 B.n243 B.n144 163.367
R386 B.n247 B.n144 163.367
R387 B.n248 B.n247 163.367
R388 B.n249 B.n248 163.367
R389 B.n249 B.n142 163.367
R390 B.n253 B.n142 163.367
R391 B.n254 B.n253 163.367
R392 B.n255 B.n254 163.367
R393 B.n255 B.n140 163.367
R394 B.n259 B.n140 163.367
R395 B.n260 B.n259 163.367
R396 B.n261 B.n260 163.367
R397 B.n261 B.n138 163.367
R398 B.n265 B.n138 163.367
R399 B.n266 B.n265 163.367
R400 B.n267 B.n266 163.367
R401 B.n267 B.n136 163.367
R402 B.n271 B.n136 163.367
R403 B.n272 B.n271 163.367
R404 B.n273 B.n272 163.367
R405 B.n273 B.n134 163.367
R406 B.n277 B.n134 163.367
R407 B.n278 B.n277 163.367
R408 B.n279 B.n278 163.367
R409 B.n279 B.n130 163.367
R410 B.n284 B.n130 163.367
R411 B.n285 B.n284 163.367
R412 B.n286 B.n285 163.367
R413 B.n286 B.n128 163.367
R414 B.n290 B.n128 163.367
R415 B.n291 B.n290 163.367
R416 B.n292 B.n291 163.367
R417 B.n292 B.n126 163.367
R418 B.n299 B.n126 163.367
R419 B.n300 B.n299 163.367
R420 B.n301 B.n300 163.367
R421 B.n301 B.n124 163.367
R422 B.n305 B.n124 163.367
R423 B.n306 B.n305 163.367
R424 B.n307 B.n306 163.367
R425 B.n307 B.n122 163.367
R426 B.n311 B.n122 163.367
R427 B.n312 B.n311 163.367
R428 B.n313 B.n312 163.367
R429 B.n313 B.n120 163.367
R430 B.n317 B.n120 163.367
R431 B.n318 B.n317 163.367
R432 B.n319 B.n318 163.367
R433 B.n319 B.n118 163.367
R434 B.n323 B.n118 163.367
R435 B.n324 B.n323 163.367
R436 B.n325 B.n324 163.367
R437 B.n325 B.n116 163.367
R438 B.n329 B.n116 163.367
R439 B.n330 B.n329 163.367
R440 B.n331 B.n330 163.367
R441 B.n331 B.n114 163.367
R442 B.n335 B.n114 163.367
R443 B.n336 B.n335 163.367
R444 B.n337 B.n336 163.367
R445 B.n337 B.n112 163.367
R446 B.n341 B.n112 163.367
R447 B.n342 B.n341 163.367
R448 B.n343 B.n342 163.367
R449 B.n343 B.n110 163.367
R450 B.n347 B.n110 163.367
R451 B.n348 B.n347 163.367
R452 B.n349 B.n348 163.367
R453 B.n349 B.n108 163.367
R454 B.n353 B.n108 163.367
R455 B.n354 B.n353 163.367
R456 B.n355 B.n354 163.367
R457 B.n355 B.n106 163.367
R458 B.n359 B.n106 163.367
R459 B.n360 B.n359 163.367
R460 B.n361 B.n360 163.367
R461 B.n361 B.n104 163.367
R462 B.n365 B.n104 163.367
R463 B.n366 B.n365 163.367
R464 B.n367 B.n366 163.367
R465 B.n367 B.n102 163.367
R466 B.n456 B.n455 163.367
R467 B.n455 B.n74 163.367
R468 B.n451 B.n74 163.367
R469 B.n451 B.n450 163.367
R470 B.n450 B.n449 163.367
R471 B.n449 B.n76 163.367
R472 B.n445 B.n76 163.367
R473 B.n445 B.n444 163.367
R474 B.n444 B.n443 163.367
R475 B.n443 B.n78 163.367
R476 B.n439 B.n78 163.367
R477 B.n439 B.n438 163.367
R478 B.n438 B.n437 163.367
R479 B.n437 B.n80 163.367
R480 B.n433 B.n80 163.367
R481 B.n433 B.n432 163.367
R482 B.n432 B.n431 163.367
R483 B.n431 B.n82 163.367
R484 B.n427 B.n82 163.367
R485 B.n427 B.n426 163.367
R486 B.n426 B.n425 163.367
R487 B.n425 B.n84 163.367
R488 B.n421 B.n84 163.367
R489 B.n421 B.n420 163.367
R490 B.n420 B.n419 163.367
R491 B.n419 B.n86 163.367
R492 B.n415 B.n86 163.367
R493 B.n415 B.n414 163.367
R494 B.n414 B.n413 163.367
R495 B.n413 B.n88 163.367
R496 B.n409 B.n88 163.367
R497 B.n409 B.n408 163.367
R498 B.n408 B.n407 163.367
R499 B.n407 B.n90 163.367
R500 B.n403 B.n90 163.367
R501 B.n403 B.n402 163.367
R502 B.n402 B.n401 163.367
R503 B.n401 B.n92 163.367
R504 B.n397 B.n92 163.367
R505 B.n397 B.n396 163.367
R506 B.n396 B.n395 163.367
R507 B.n395 B.n94 163.367
R508 B.n391 B.n94 163.367
R509 B.n391 B.n390 163.367
R510 B.n390 B.n389 163.367
R511 B.n389 B.n96 163.367
R512 B.n385 B.n96 163.367
R513 B.n385 B.n384 163.367
R514 B.n384 B.n383 163.367
R515 B.n383 B.n98 163.367
R516 B.n379 B.n98 163.367
R517 B.n379 B.n378 163.367
R518 B.n378 B.n377 163.367
R519 B.n377 B.n100 163.367
R520 B.n373 B.n100 163.367
R521 B.n373 B.n372 163.367
R522 B.n372 B.n371 163.367
R523 B.n613 B.n612 163.367
R524 B.n612 B.n17 163.367
R525 B.n608 B.n17 163.367
R526 B.n608 B.n607 163.367
R527 B.n607 B.n606 163.367
R528 B.n606 B.n19 163.367
R529 B.n602 B.n19 163.367
R530 B.n602 B.n601 163.367
R531 B.n601 B.n600 163.367
R532 B.n600 B.n21 163.367
R533 B.n596 B.n21 163.367
R534 B.n596 B.n595 163.367
R535 B.n595 B.n594 163.367
R536 B.n594 B.n23 163.367
R537 B.n590 B.n23 163.367
R538 B.n590 B.n589 163.367
R539 B.n589 B.n588 163.367
R540 B.n588 B.n25 163.367
R541 B.n584 B.n25 163.367
R542 B.n584 B.n583 163.367
R543 B.n583 B.n582 163.367
R544 B.n582 B.n27 163.367
R545 B.n578 B.n27 163.367
R546 B.n578 B.n577 163.367
R547 B.n577 B.n576 163.367
R548 B.n576 B.n29 163.367
R549 B.n572 B.n29 163.367
R550 B.n572 B.n571 163.367
R551 B.n571 B.n570 163.367
R552 B.n570 B.n31 163.367
R553 B.n566 B.n31 163.367
R554 B.n566 B.n565 163.367
R555 B.n565 B.n564 163.367
R556 B.n564 B.n33 163.367
R557 B.n560 B.n33 163.367
R558 B.n560 B.n559 163.367
R559 B.n559 B.n558 163.367
R560 B.n558 B.n35 163.367
R561 B.n554 B.n35 163.367
R562 B.n554 B.n553 163.367
R563 B.n553 B.n552 163.367
R564 B.n552 B.n37 163.367
R565 B.n548 B.n37 163.367
R566 B.n548 B.n547 163.367
R567 B.n547 B.n546 163.367
R568 B.n546 B.n39 163.367
R569 B.n541 B.n39 163.367
R570 B.n541 B.n540 163.367
R571 B.n540 B.n539 163.367
R572 B.n539 B.n43 163.367
R573 B.n535 B.n43 163.367
R574 B.n535 B.n534 163.367
R575 B.n534 B.n533 163.367
R576 B.n533 B.n45 163.367
R577 B.n529 B.n45 163.367
R578 B.n529 B.n528 163.367
R579 B.n528 B.n527 163.367
R580 B.n527 B.n47 163.367
R581 B.n523 B.n47 163.367
R582 B.n523 B.n522 163.367
R583 B.n522 B.n521 163.367
R584 B.n521 B.n52 163.367
R585 B.n517 B.n52 163.367
R586 B.n517 B.n516 163.367
R587 B.n516 B.n515 163.367
R588 B.n515 B.n54 163.367
R589 B.n511 B.n54 163.367
R590 B.n511 B.n510 163.367
R591 B.n510 B.n509 163.367
R592 B.n509 B.n56 163.367
R593 B.n505 B.n56 163.367
R594 B.n505 B.n504 163.367
R595 B.n504 B.n503 163.367
R596 B.n503 B.n58 163.367
R597 B.n499 B.n58 163.367
R598 B.n499 B.n498 163.367
R599 B.n498 B.n497 163.367
R600 B.n497 B.n60 163.367
R601 B.n493 B.n60 163.367
R602 B.n493 B.n492 163.367
R603 B.n492 B.n491 163.367
R604 B.n491 B.n62 163.367
R605 B.n487 B.n62 163.367
R606 B.n487 B.n486 163.367
R607 B.n486 B.n485 163.367
R608 B.n485 B.n64 163.367
R609 B.n481 B.n64 163.367
R610 B.n481 B.n480 163.367
R611 B.n480 B.n479 163.367
R612 B.n479 B.n66 163.367
R613 B.n475 B.n66 163.367
R614 B.n475 B.n474 163.367
R615 B.n474 B.n473 163.367
R616 B.n473 B.n68 163.367
R617 B.n469 B.n68 163.367
R618 B.n469 B.n468 163.367
R619 B.n468 B.n467 163.367
R620 B.n467 B.n70 163.367
R621 B.n463 B.n70 163.367
R622 B.n463 B.n462 163.367
R623 B.n462 B.n461 163.367
R624 B.n461 B.n72 163.367
R625 B.n457 B.n72 163.367
R626 B.n614 B.n15 163.367
R627 B.n618 B.n15 163.367
R628 B.n619 B.n618 163.367
R629 B.n620 B.n619 163.367
R630 B.n620 B.n13 163.367
R631 B.n624 B.n13 163.367
R632 B.n625 B.n624 163.367
R633 B.n626 B.n625 163.367
R634 B.n626 B.n11 163.367
R635 B.n630 B.n11 163.367
R636 B.n631 B.n630 163.367
R637 B.n632 B.n631 163.367
R638 B.n632 B.n9 163.367
R639 B.n636 B.n9 163.367
R640 B.n637 B.n636 163.367
R641 B.n638 B.n637 163.367
R642 B.n638 B.n7 163.367
R643 B.n642 B.n7 163.367
R644 B.n643 B.n642 163.367
R645 B.n644 B.n643 163.367
R646 B.n644 B.n5 163.367
R647 B.n648 B.n5 163.367
R648 B.n649 B.n648 163.367
R649 B.n650 B.n649 163.367
R650 B.n650 B.n3 163.367
R651 B.n654 B.n3 163.367
R652 B.n655 B.n654 163.367
R653 B.n170 B.n2 163.367
R654 B.n171 B.n170 163.367
R655 B.n171 B.n168 163.367
R656 B.n175 B.n168 163.367
R657 B.n176 B.n175 163.367
R658 B.n177 B.n176 163.367
R659 B.n177 B.n166 163.367
R660 B.n181 B.n166 163.367
R661 B.n182 B.n181 163.367
R662 B.n183 B.n182 163.367
R663 B.n183 B.n164 163.367
R664 B.n187 B.n164 163.367
R665 B.n188 B.n187 163.367
R666 B.n189 B.n188 163.367
R667 B.n189 B.n162 163.367
R668 B.n193 B.n162 163.367
R669 B.n194 B.n193 163.367
R670 B.n195 B.n194 163.367
R671 B.n195 B.n160 163.367
R672 B.n199 B.n160 163.367
R673 B.n200 B.n199 163.367
R674 B.n201 B.n200 163.367
R675 B.n201 B.n158 163.367
R676 B.n205 B.n158 163.367
R677 B.n206 B.n205 163.367
R678 B.n207 B.n206 163.367
R679 B.n207 B.n156 163.367
R680 B.n295 B.t4 156.577
R681 B.n48 B.t2 156.577
R682 B.n131 B.t7 156.56
R683 B.n40 B.t11 156.56
R684 B.n296 B.t5 112.165
R685 B.n49 B.t1 112.165
R686 B.n132 B.t8 112.148
R687 B.n41 B.t10 112.148
R688 B.n281 B.n132 59.5399
R689 B.n297 B.n296 59.5399
R690 B.n50 B.n49 59.5399
R691 B.n543 B.n41 59.5399
R692 B.n132 B.n131 44.4126
R693 B.n296 B.n295 44.4126
R694 B.n49 B.n48 44.4126
R695 B.n41 B.n40 44.4126
R696 B.n615 B.n16 29.8151
R697 B.n458 B.n73 29.8151
R698 B.n210 B.n209 29.8151
R699 B.n370 B.n369 29.8151
R700 B B.n657 18.0485
R701 B.n616 B.n615 10.6151
R702 B.n617 B.n616 10.6151
R703 B.n617 B.n14 10.6151
R704 B.n621 B.n14 10.6151
R705 B.n622 B.n621 10.6151
R706 B.n623 B.n622 10.6151
R707 B.n623 B.n12 10.6151
R708 B.n627 B.n12 10.6151
R709 B.n628 B.n627 10.6151
R710 B.n629 B.n628 10.6151
R711 B.n629 B.n10 10.6151
R712 B.n633 B.n10 10.6151
R713 B.n634 B.n633 10.6151
R714 B.n635 B.n634 10.6151
R715 B.n635 B.n8 10.6151
R716 B.n639 B.n8 10.6151
R717 B.n640 B.n639 10.6151
R718 B.n641 B.n640 10.6151
R719 B.n641 B.n6 10.6151
R720 B.n645 B.n6 10.6151
R721 B.n646 B.n645 10.6151
R722 B.n647 B.n646 10.6151
R723 B.n647 B.n4 10.6151
R724 B.n651 B.n4 10.6151
R725 B.n652 B.n651 10.6151
R726 B.n653 B.n652 10.6151
R727 B.n653 B.n0 10.6151
R728 B.n611 B.n16 10.6151
R729 B.n611 B.n610 10.6151
R730 B.n610 B.n609 10.6151
R731 B.n609 B.n18 10.6151
R732 B.n605 B.n18 10.6151
R733 B.n605 B.n604 10.6151
R734 B.n604 B.n603 10.6151
R735 B.n603 B.n20 10.6151
R736 B.n599 B.n20 10.6151
R737 B.n599 B.n598 10.6151
R738 B.n598 B.n597 10.6151
R739 B.n597 B.n22 10.6151
R740 B.n593 B.n22 10.6151
R741 B.n593 B.n592 10.6151
R742 B.n592 B.n591 10.6151
R743 B.n591 B.n24 10.6151
R744 B.n587 B.n24 10.6151
R745 B.n587 B.n586 10.6151
R746 B.n586 B.n585 10.6151
R747 B.n585 B.n26 10.6151
R748 B.n581 B.n26 10.6151
R749 B.n581 B.n580 10.6151
R750 B.n580 B.n579 10.6151
R751 B.n579 B.n28 10.6151
R752 B.n575 B.n28 10.6151
R753 B.n575 B.n574 10.6151
R754 B.n574 B.n573 10.6151
R755 B.n573 B.n30 10.6151
R756 B.n569 B.n30 10.6151
R757 B.n569 B.n568 10.6151
R758 B.n568 B.n567 10.6151
R759 B.n567 B.n32 10.6151
R760 B.n563 B.n32 10.6151
R761 B.n563 B.n562 10.6151
R762 B.n562 B.n561 10.6151
R763 B.n561 B.n34 10.6151
R764 B.n557 B.n34 10.6151
R765 B.n557 B.n556 10.6151
R766 B.n556 B.n555 10.6151
R767 B.n555 B.n36 10.6151
R768 B.n551 B.n36 10.6151
R769 B.n551 B.n550 10.6151
R770 B.n550 B.n549 10.6151
R771 B.n549 B.n38 10.6151
R772 B.n545 B.n38 10.6151
R773 B.n545 B.n544 10.6151
R774 B.n542 B.n42 10.6151
R775 B.n538 B.n42 10.6151
R776 B.n538 B.n537 10.6151
R777 B.n537 B.n536 10.6151
R778 B.n536 B.n44 10.6151
R779 B.n532 B.n44 10.6151
R780 B.n532 B.n531 10.6151
R781 B.n531 B.n530 10.6151
R782 B.n530 B.n46 10.6151
R783 B.n526 B.n525 10.6151
R784 B.n525 B.n524 10.6151
R785 B.n524 B.n51 10.6151
R786 B.n520 B.n51 10.6151
R787 B.n520 B.n519 10.6151
R788 B.n519 B.n518 10.6151
R789 B.n518 B.n53 10.6151
R790 B.n514 B.n53 10.6151
R791 B.n514 B.n513 10.6151
R792 B.n513 B.n512 10.6151
R793 B.n512 B.n55 10.6151
R794 B.n508 B.n55 10.6151
R795 B.n508 B.n507 10.6151
R796 B.n507 B.n506 10.6151
R797 B.n506 B.n57 10.6151
R798 B.n502 B.n57 10.6151
R799 B.n502 B.n501 10.6151
R800 B.n501 B.n500 10.6151
R801 B.n500 B.n59 10.6151
R802 B.n496 B.n59 10.6151
R803 B.n496 B.n495 10.6151
R804 B.n495 B.n494 10.6151
R805 B.n494 B.n61 10.6151
R806 B.n490 B.n61 10.6151
R807 B.n490 B.n489 10.6151
R808 B.n489 B.n488 10.6151
R809 B.n488 B.n63 10.6151
R810 B.n484 B.n63 10.6151
R811 B.n484 B.n483 10.6151
R812 B.n483 B.n482 10.6151
R813 B.n482 B.n65 10.6151
R814 B.n478 B.n65 10.6151
R815 B.n478 B.n477 10.6151
R816 B.n477 B.n476 10.6151
R817 B.n476 B.n67 10.6151
R818 B.n472 B.n67 10.6151
R819 B.n472 B.n471 10.6151
R820 B.n471 B.n470 10.6151
R821 B.n470 B.n69 10.6151
R822 B.n466 B.n69 10.6151
R823 B.n466 B.n465 10.6151
R824 B.n465 B.n464 10.6151
R825 B.n464 B.n71 10.6151
R826 B.n460 B.n71 10.6151
R827 B.n460 B.n459 10.6151
R828 B.n459 B.n458 10.6151
R829 B.n454 B.n73 10.6151
R830 B.n454 B.n453 10.6151
R831 B.n453 B.n452 10.6151
R832 B.n452 B.n75 10.6151
R833 B.n448 B.n75 10.6151
R834 B.n448 B.n447 10.6151
R835 B.n447 B.n446 10.6151
R836 B.n446 B.n77 10.6151
R837 B.n442 B.n77 10.6151
R838 B.n442 B.n441 10.6151
R839 B.n441 B.n440 10.6151
R840 B.n440 B.n79 10.6151
R841 B.n436 B.n79 10.6151
R842 B.n436 B.n435 10.6151
R843 B.n435 B.n434 10.6151
R844 B.n434 B.n81 10.6151
R845 B.n430 B.n81 10.6151
R846 B.n430 B.n429 10.6151
R847 B.n429 B.n428 10.6151
R848 B.n428 B.n83 10.6151
R849 B.n424 B.n83 10.6151
R850 B.n424 B.n423 10.6151
R851 B.n423 B.n422 10.6151
R852 B.n422 B.n85 10.6151
R853 B.n418 B.n85 10.6151
R854 B.n418 B.n417 10.6151
R855 B.n417 B.n416 10.6151
R856 B.n416 B.n87 10.6151
R857 B.n412 B.n87 10.6151
R858 B.n412 B.n411 10.6151
R859 B.n411 B.n410 10.6151
R860 B.n410 B.n89 10.6151
R861 B.n406 B.n89 10.6151
R862 B.n406 B.n405 10.6151
R863 B.n405 B.n404 10.6151
R864 B.n404 B.n91 10.6151
R865 B.n400 B.n91 10.6151
R866 B.n400 B.n399 10.6151
R867 B.n399 B.n398 10.6151
R868 B.n398 B.n93 10.6151
R869 B.n394 B.n93 10.6151
R870 B.n394 B.n393 10.6151
R871 B.n393 B.n392 10.6151
R872 B.n392 B.n95 10.6151
R873 B.n388 B.n95 10.6151
R874 B.n388 B.n387 10.6151
R875 B.n387 B.n386 10.6151
R876 B.n386 B.n97 10.6151
R877 B.n382 B.n97 10.6151
R878 B.n382 B.n381 10.6151
R879 B.n381 B.n380 10.6151
R880 B.n380 B.n99 10.6151
R881 B.n376 B.n99 10.6151
R882 B.n376 B.n375 10.6151
R883 B.n375 B.n374 10.6151
R884 B.n374 B.n101 10.6151
R885 B.n370 B.n101 10.6151
R886 B.n169 B.n1 10.6151
R887 B.n172 B.n169 10.6151
R888 B.n173 B.n172 10.6151
R889 B.n174 B.n173 10.6151
R890 B.n174 B.n167 10.6151
R891 B.n178 B.n167 10.6151
R892 B.n179 B.n178 10.6151
R893 B.n180 B.n179 10.6151
R894 B.n180 B.n165 10.6151
R895 B.n184 B.n165 10.6151
R896 B.n185 B.n184 10.6151
R897 B.n186 B.n185 10.6151
R898 B.n186 B.n163 10.6151
R899 B.n190 B.n163 10.6151
R900 B.n191 B.n190 10.6151
R901 B.n192 B.n191 10.6151
R902 B.n192 B.n161 10.6151
R903 B.n196 B.n161 10.6151
R904 B.n197 B.n196 10.6151
R905 B.n198 B.n197 10.6151
R906 B.n198 B.n159 10.6151
R907 B.n202 B.n159 10.6151
R908 B.n203 B.n202 10.6151
R909 B.n204 B.n203 10.6151
R910 B.n204 B.n157 10.6151
R911 B.n208 B.n157 10.6151
R912 B.n209 B.n208 10.6151
R913 B.n210 B.n155 10.6151
R914 B.n214 B.n155 10.6151
R915 B.n215 B.n214 10.6151
R916 B.n216 B.n215 10.6151
R917 B.n216 B.n153 10.6151
R918 B.n220 B.n153 10.6151
R919 B.n221 B.n220 10.6151
R920 B.n222 B.n221 10.6151
R921 B.n222 B.n151 10.6151
R922 B.n226 B.n151 10.6151
R923 B.n227 B.n226 10.6151
R924 B.n228 B.n227 10.6151
R925 B.n228 B.n149 10.6151
R926 B.n232 B.n149 10.6151
R927 B.n233 B.n232 10.6151
R928 B.n234 B.n233 10.6151
R929 B.n234 B.n147 10.6151
R930 B.n238 B.n147 10.6151
R931 B.n239 B.n238 10.6151
R932 B.n240 B.n239 10.6151
R933 B.n240 B.n145 10.6151
R934 B.n244 B.n145 10.6151
R935 B.n245 B.n244 10.6151
R936 B.n246 B.n245 10.6151
R937 B.n246 B.n143 10.6151
R938 B.n250 B.n143 10.6151
R939 B.n251 B.n250 10.6151
R940 B.n252 B.n251 10.6151
R941 B.n252 B.n141 10.6151
R942 B.n256 B.n141 10.6151
R943 B.n257 B.n256 10.6151
R944 B.n258 B.n257 10.6151
R945 B.n258 B.n139 10.6151
R946 B.n262 B.n139 10.6151
R947 B.n263 B.n262 10.6151
R948 B.n264 B.n263 10.6151
R949 B.n264 B.n137 10.6151
R950 B.n268 B.n137 10.6151
R951 B.n269 B.n268 10.6151
R952 B.n270 B.n269 10.6151
R953 B.n270 B.n135 10.6151
R954 B.n274 B.n135 10.6151
R955 B.n275 B.n274 10.6151
R956 B.n276 B.n275 10.6151
R957 B.n276 B.n133 10.6151
R958 B.n280 B.n133 10.6151
R959 B.n283 B.n282 10.6151
R960 B.n283 B.n129 10.6151
R961 B.n287 B.n129 10.6151
R962 B.n288 B.n287 10.6151
R963 B.n289 B.n288 10.6151
R964 B.n289 B.n127 10.6151
R965 B.n293 B.n127 10.6151
R966 B.n294 B.n293 10.6151
R967 B.n298 B.n294 10.6151
R968 B.n302 B.n125 10.6151
R969 B.n303 B.n302 10.6151
R970 B.n304 B.n303 10.6151
R971 B.n304 B.n123 10.6151
R972 B.n308 B.n123 10.6151
R973 B.n309 B.n308 10.6151
R974 B.n310 B.n309 10.6151
R975 B.n310 B.n121 10.6151
R976 B.n314 B.n121 10.6151
R977 B.n315 B.n314 10.6151
R978 B.n316 B.n315 10.6151
R979 B.n316 B.n119 10.6151
R980 B.n320 B.n119 10.6151
R981 B.n321 B.n320 10.6151
R982 B.n322 B.n321 10.6151
R983 B.n322 B.n117 10.6151
R984 B.n326 B.n117 10.6151
R985 B.n327 B.n326 10.6151
R986 B.n328 B.n327 10.6151
R987 B.n328 B.n115 10.6151
R988 B.n332 B.n115 10.6151
R989 B.n333 B.n332 10.6151
R990 B.n334 B.n333 10.6151
R991 B.n334 B.n113 10.6151
R992 B.n338 B.n113 10.6151
R993 B.n339 B.n338 10.6151
R994 B.n340 B.n339 10.6151
R995 B.n340 B.n111 10.6151
R996 B.n344 B.n111 10.6151
R997 B.n345 B.n344 10.6151
R998 B.n346 B.n345 10.6151
R999 B.n346 B.n109 10.6151
R1000 B.n350 B.n109 10.6151
R1001 B.n351 B.n350 10.6151
R1002 B.n352 B.n351 10.6151
R1003 B.n352 B.n107 10.6151
R1004 B.n356 B.n107 10.6151
R1005 B.n357 B.n356 10.6151
R1006 B.n358 B.n357 10.6151
R1007 B.n358 B.n105 10.6151
R1008 B.n362 B.n105 10.6151
R1009 B.n363 B.n362 10.6151
R1010 B.n364 B.n363 10.6151
R1011 B.n364 B.n103 10.6151
R1012 B.n368 B.n103 10.6151
R1013 B.n369 B.n368 10.6151
R1014 B.n544 B.n543 9.36635
R1015 B.n526 B.n50 9.36635
R1016 B.n281 B.n280 9.36635
R1017 B.n297 B.n125 9.36635
R1018 B.n657 B.n0 8.11757
R1019 B.n657 B.n1 8.11757
R1020 B.n543 B.n542 1.24928
R1021 B.n50 B.n46 1.24928
R1022 B.n282 B.n281 1.24928
R1023 B.n298 B.n297 1.24928
R1024 VP.n2 VP.t1 205.95
R1025 VP.n2 VP.t0 205.424
R1026 VP.n4 VP.t3 170.667
R1027 VP.n11 VP.t2 170.667
R1028 VP.n10 VP.n0 161.3
R1029 VP.n9 VP.n8 161.3
R1030 VP.n7 VP.n1 161.3
R1031 VP.n6 VP.n5 161.3
R1032 VP.n4 VP.n3 91.3749
R1033 VP.n12 VP.n11 91.3749
R1034 VP.n9 VP.n1 56.4773
R1035 VP.n3 VP.n2 53.1567
R1036 VP.n5 VP.n1 24.3439
R1037 VP.n10 VP.n9 24.3439
R1038 VP.n5 VP.n4 19.2318
R1039 VP.n11 VP.n10 19.2318
R1040 VP.n6 VP.n3 0.278398
R1041 VP.n12 VP.n0 0.278398
R1042 VP.n7 VP.n6 0.189894
R1043 VP.n8 VP.n7 0.189894
R1044 VP.n8 VP.n0 0.189894
R1045 VP VP.n12 0.153422
R1046 VDD1 VDD1.n1 113.299
R1047 VDD1 VDD1.n0 71.2296
R1048 VDD1.n0 VDD1.t2 2.34236
R1049 VDD1.n0 VDD1.t3 2.34236
R1050 VDD1.n1 VDD1.t0 2.34236
R1051 VDD1.n1 VDD1.t1 2.34236
C0 VP B 1.5005f
C1 VDD1 w_n2344_n3744# 1.38099f
C2 VTAIL w_n2344_n3744# 4.40615f
C3 VTAIL VDD1 5.8879f
C4 VN w_n2344_n3744# 3.89591f
C5 VN VDD1 0.148213f
C6 VN VTAIL 4.88364f
C7 VDD2 w_n2344_n3744# 1.42279f
C8 VDD2 VDD1 0.873787f
C9 VTAIL VDD2 5.93781f
C10 B w_n2344_n3744# 8.98545f
C11 VN VDD2 5.13527f
C12 VP w_n2344_n3744# 4.19562f
C13 B VDD1 1.20045f
C14 B VTAIL 5.22508f
C15 VP VDD1 5.33985f
C16 VP VTAIL 4.89775f
C17 VN B 1.00612f
C18 VN VP 6.084f
C19 B VDD2 1.24212f
C20 VP VDD2 0.353373f
C21 VDD2 VSUBS 0.88644f
C22 VDD1 VSUBS 5.6207f
C23 VTAIL VSUBS 1.228374f
C24 VN VSUBS 5.2816f
C25 VP VSUBS 2.025104f
C26 B VSUBS 3.878968f
C27 w_n2344_n3744# VSUBS 0.107758p
C28 VDD1.t2 VSUBS 0.292517f
C29 VDD1.t3 VSUBS 0.292517f
C30 VDD1.n0 VSUBS 2.33335f
C31 VDD1.t0 VSUBS 0.292517f
C32 VDD1.t1 VSUBS 0.292517f
C33 VDD1.n1 VSUBS 3.1127f
C34 VP.n0 VSUBS 0.050136f
C35 VP.t2 VSUBS 2.82945f
C36 VP.n1 VSUBS 0.055752f
C37 VP.t0 VSUBS 3.03179f
C38 VP.t1 VSUBS 3.03487f
C39 VP.n2 VSUBS 3.88072f
C40 VP.n3 VSUBS 2.15928f
C41 VP.t3 VSUBS 2.82945f
C42 VP.n4 VSUBS 1.11538f
C43 VP.n5 VSUBS 0.06384f
C44 VP.n6 VSUBS 0.050136f
C45 VP.n7 VSUBS 0.038025f
C46 VP.n8 VSUBS 0.038025f
C47 VP.n9 VSUBS 0.055752f
C48 VP.n10 VSUBS 0.06384f
C49 VP.n11 VSUBS 1.11538f
C50 VP.n12 VSUBS 0.046411f
C51 B.n0 VSUBS 0.006056f
C52 B.n1 VSUBS 0.006056f
C53 B.n2 VSUBS 0.008957f
C54 B.n3 VSUBS 0.006864f
C55 B.n4 VSUBS 0.006864f
C56 B.n5 VSUBS 0.006864f
C57 B.n6 VSUBS 0.006864f
C58 B.n7 VSUBS 0.006864f
C59 B.n8 VSUBS 0.006864f
C60 B.n9 VSUBS 0.006864f
C61 B.n10 VSUBS 0.006864f
C62 B.n11 VSUBS 0.006864f
C63 B.n12 VSUBS 0.006864f
C64 B.n13 VSUBS 0.006864f
C65 B.n14 VSUBS 0.006864f
C66 B.n15 VSUBS 0.006864f
C67 B.n16 VSUBS 0.015476f
C68 B.n17 VSUBS 0.006864f
C69 B.n18 VSUBS 0.006864f
C70 B.n19 VSUBS 0.006864f
C71 B.n20 VSUBS 0.006864f
C72 B.n21 VSUBS 0.006864f
C73 B.n22 VSUBS 0.006864f
C74 B.n23 VSUBS 0.006864f
C75 B.n24 VSUBS 0.006864f
C76 B.n25 VSUBS 0.006864f
C77 B.n26 VSUBS 0.006864f
C78 B.n27 VSUBS 0.006864f
C79 B.n28 VSUBS 0.006864f
C80 B.n29 VSUBS 0.006864f
C81 B.n30 VSUBS 0.006864f
C82 B.n31 VSUBS 0.006864f
C83 B.n32 VSUBS 0.006864f
C84 B.n33 VSUBS 0.006864f
C85 B.n34 VSUBS 0.006864f
C86 B.n35 VSUBS 0.006864f
C87 B.n36 VSUBS 0.006864f
C88 B.n37 VSUBS 0.006864f
C89 B.n38 VSUBS 0.006864f
C90 B.n39 VSUBS 0.006864f
C91 B.t10 VSUBS 0.449985f
C92 B.t11 VSUBS 0.466471f
C93 B.t9 VSUBS 1.1791f
C94 B.n40 VSUBS 0.225972f
C95 B.n41 VSUBS 0.067904f
C96 B.n42 VSUBS 0.006864f
C97 B.n43 VSUBS 0.006864f
C98 B.n44 VSUBS 0.006864f
C99 B.n45 VSUBS 0.006864f
C100 B.n46 VSUBS 0.003836f
C101 B.n47 VSUBS 0.006864f
C102 B.t1 VSUBS 0.449974f
C103 B.t2 VSUBS 0.466461f
C104 B.t0 VSUBS 1.1791f
C105 B.n48 VSUBS 0.225982f
C106 B.n49 VSUBS 0.067915f
C107 B.n50 VSUBS 0.015902f
C108 B.n51 VSUBS 0.006864f
C109 B.n52 VSUBS 0.006864f
C110 B.n53 VSUBS 0.006864f
C111 B.n54 VSUBS 0.006864f
C112 B.n55 VSUBS 0.006864f
C113 B.n56 VSUBS 0.006864f
C114 B.n57 VSUBS 0.006864f
C115 B.n58 VSUBS 0.006864f
C116 B.n59 VSUBS 0.006864f
C117 B.n60 VSUBS 0.006864f
C118 B.n61 VSUBS 0.006864f
C119 B.n62 VSUBS 0.006864f
C120 B.n63 VSUBS 0.006864f
C121 B.n64 VSUBS 0.006864f
C122 B.n65 VSUBS 0.006864f
C123 B.n66 VSUBS 0.006864f
C124 B.n67 VSUBS 0.006864f
C125 B.n68 VSUBS 0.006864f
C126 B.n69 VSUBS 0.006864f
C127 B.n70 VSUBS 0.006864f
C128 B.n71 VSUBS 0.006864f
C129 B.n72 VSUBS 0.006864f
C130 B.n73 VSUBS 0.014805f
C131 B.n74 VSUBS 0.006864f
C132 B.n75 VSUBS 0.006864f
C133 B.n76 VSUBS 0.006864f
C134 B.n77 VSUBS 0.006864f
C135 B.n78 VSUBS 0.006864f
C136 B.n79 VSUBS 0.006864f
C137 B.n80 VSUBS 0.006864f
C138 B.n81 VSUBS 0.006864f
C139 B.n82 VSUBS 0.006864f
C140 B.n83 VSUBS 0.006864f
C141 B.n84 VSUBS 0.006864f
C142 B.n85 VSUBS 0.006864f
C143 B.n86 VSUBS 0.006864f
C144 B.n87 VSUBS 0.006864f
C145 B.n88 VSUBS 0.006864f
C146 B.n89 VSUBS 0.006864f
C147 B.n90 VSUBS 0.006864f
C148 B.n91 VSUBS 0.006864f
C149 B.n92 VSUBS 0.006864f
C150 B.n93 VSUBS 0.006864f
C151 B.n94 VSUBS 0.006864f
C152 B.n95 VSUBS 0.006864f
C153 B.n96 VSUBS 0.006864f
C154 B.n97 VSUBS 0.006864f
C155 B.n98 VSUBS 0.006864f
C156 B.n99 VSUBS 0.006864f
C157 B.n100 VSUBS 0.006864f
C158 B.n101 VSUBS 0.006864f
C159 B.n102 VSUBS 0.015476f
C160 B.n103 VSUBS 0.006864f
C161 B.n104 VSUBS 0.006864f
C162 B.n105 VSUBS 0.006864f
C163 B.n106 VSUBS 0.006864f
C164 B.n107 VSUBS 0.006864f
C165 B.n108 VSUBS 0.006864f
C166 B.n109 VSUBS 0.006864f
C167 B.n110 VSUBS 0.006864f
C168 B.n111 VSUBS 0.006864f
C169 B.n112 VSUBS 0.006864f
C170 B.n113 VSUBS 0.006864f
C171 B.n114 VSUBS 0.006864f
C172 B.n115 VSUBS 0.006864f
C173 B.n116 VSUBS 0.006864f
C174 B.n117 VSUBS 0.006864f
C175 B.n118 VSUBS 0.006864f
C176 B.n119 VSUBS 0.006864f
C177 B.n120 VSUBS 0.006864f
C178 B.n121 VSUBS 0.006864f
C179 B.n122 VSUBS 0.006864f
C180 B.n123 VSUBS 0.006864f
C181 B.n124 VSUBS 0.006864f
C182 B.n125 VSUBS 0.00646f
C183 B.n126 VSUBS 0.006864f
C184 B.n127 VSUBS 0.006864f
C185 B.n128 VSUBS 0.006864f
C186 B.n129 VSUBS 0.006864f
C187 B.n130 VSUBS 0.006864f
C188 B.t8 VSUBS 0.449985f
C189 B.t7 VSUBS 0.466471f
C190 B.t6 VSUBS 1.1791f
C191 B.n131 VSUBS 0.225972f
C192 B.n132 VSUBS 0.067904f
C193 B.n133 VSUBS 0.006864f
C194 B.n134 VSUBS 0.006864f
C195 B.n135 VSUBS 0.006864f
C196 B.n136 VSUBS 0.006864f
C197 B.n137 VSUBS 0.006864f
C198 B.n138 VSUBS 0.006864f
C199 B.n139 VSUBS 0.006864f
C200 B.n140 VSUBS 0.006864f
C201 B.n141 VSUBS 0.006864f
C202 B.n142 VSUBS 0.006864f
C203 B.n143 VSUBS 0.006864f
C204 B.n144 VSUBS 0.006864f
C205 B.n145 VSUBS 0.006864f
C206 B.n146 VSUBS 0.006864f
C207 B.n147 VSUBS 0.006864f
C208 B.n148 VSUBS 0.006864f
C209 B.n149 VSUBS 0.006864f
C210 B.n150 VSUBS 0.006864f
C211 B.n151 VSUBS 0.006864f
C212 B.n152 VSUBS 0.006864f
C213 B.n153 VSUBS 0.006864f
C214 B.n154 VSUBS 0.006864f
C215 B.n155 VSUBS 0.006864f
C216 B.n156 VSUBS 0.014805f
C217 B.n157 VSUBS 0.006864f
C218 B.n158 VSUBS 0.006864f
C219 B.n159 VSUBS 0.006864f
C220 B.n160 VSUBS 0.006864f
C221 B.n161 VSUBS 0.006864f
C222 B.n162 VSUBS 0.006864f
C223 B.n163 VSUBS 0.006864f
C224 B.n164 VSUBS 0.006864f
C225 B.n165 VSUBS 0.006864f
C226 B.n166 VSUBS 0.006864f
C227 B.n167 VSUBS 0.006864f
C228 B.n168 VSUBS 0.006864f
C229 B.n169 VSUBS 0.006864f
C230 B.n170 VSUBS 0.006864f
C231 B.n171 VSUBS 0.006864f
C232 B.n172 VSUBS 0.006864f
C233 B.n173 VSUBS 0.006864f
C234 B.n174 VSUBS 0.006864f
C235 B.n175 VSUBS 0.006864f
C236 B.n176 VSUBS 0.006864f
C237 B.n177 VSUBS 0.006864f
C238 B.n178 VSUBS 0.006864f
C239 B.n179 VSUBS 0.006864f
C240 B.n180 VSUBS 0.006864f
C241 B.n181 VSUBS 0.006864f
C242 B.n182 VSUBS 0.006864f
C243 B.n183 VSUBS 0.006864f
C244 B.n184 VSUBS 0.006864f
C245 B.n185 VSUBS 0.006864f
C246 B.n186 VSUBS 0.006864f
C247 B.n187 VSUBS 0.006864f
C248 B.n188 VSUBS 0.006864f
C249 B.n189 VSUBS 0.006864f
C250 B.n190 VSUBS 0.006864f
C251 B.n191 VSUBS 0.006864f
C252 B.n192 VSUBS 0.006864f
C253 B.n193 VSUBS 0.006864f
C254 B.n194 VSUBS 0.006864f
C255 B.n195 VSUBS 0.006864f
C256 B.n196 VSUBS 0.006864f
C257 B.n197 VSUBS 0.006864f
C258 B.n198 VSUBS 0.006864f
C259 B.n199 VSUBS 0.006864f
C260 B.n200 VSUBS 0.006864f
C261 B.n201 VSUBS 0.006864f
C262 B.n202 VSUBS 0.006864f
C263 B.n203 VSUBS 0.006864f
C264 B.n204 VSUBS 0.006864f
C265 B.n205 VSUBS 0.006864f
C266 B.n206 VSUBS 0.006864f
C267 B.n207 VSUBS 0.006864f
C268 B.n208 VSUBS 0.006864f
C269 B.n209 VSUBS 0.014805f
C270 B.n210 VSUBS 0.015476f
C271 B.n211 VSUBS 0.015476f
C272 B.n212 VSUBS 0.006864f
C273 B.n213 VSUBS 0.006864f
C274 B.n214 VSUBS 0.006864f
C275 B.n215 VSUBS 0.006864f
C276 B.n216 VSUBS 0.006864f
C277 B.n217 VSUBS 0.006864f
C278 B.n218 VSUBS 0.006864f
C279 B.n219 VSUBS 0.006864f
C280 B.n220 VSUBS 0.006864f
C281 B.n221 VSUBS 0.006864f
C282 B.n222 VSUBS 0.006864f
C283 B.n223 VSUBS 0.006864f
C284 B.n224 VSUBS 0.006864f
C285 B.n225 VSUBS 0.006864f
C286 B.n226 VSUBS 0.006864f
C287 B.n227 VSUBS 0.006864f
C288 B.n228 VSUBS 0.006864f
C289 B.n229 VSUBS 0.006864f
C290 B.n230 VSUBS 0.006864f
C291 B.n231 VSUBS 0.006864f
C292 B.n232 VSUBS 0.006864f
C293 B.n233 VSUBS 0.006864f
C294 B.n234 VSUBS 0.006864f
C295 B.n235 VSUBS 0.006864f
C296 B.n236 VSUBS 0.006864f
C297 B.n237 VSUBS 0.006864f
C298 B.n238 VSUBS 0.006864f
C299 B.n239 VSUBS 0.006864f
C300 B.n240 VSUBS 0.006864f
C301 B.n241 VSUBS 0.006864f
C302 B.n242 VSUBS 0.006864f
C303 B.n243 VSUBS 0.006864f
C304 B.n244 VSUBS 0.006864f
C305 B.n245 VSUBS 0.006864f
C306 B.n246 VSUBS 0.006864f
C307 B.n247 VSUBS 0.006864f
C308 B.n248 VSUBS 0.006864f
C309 B.n249 VSUBS 0.006864f
C310 B.n250 VSUBS 0.006864f
C311 B.n251 VSUBS 0.006864f
C312 B.n252 VSUBS 0.006864f
C313 B.n253 VSUBS 0.006864f
C314 B.n254 VSUBS 0.006864f
C315 B.n255 VSUBS 0.006864f
C316 B.n256 VSUBS 0.006864f
C317 B.n257 VSUBS 0.006864f
C318 B.n258 VSUBS 0.006864f
C319 B.n259 VSUBS 0.006864f
C320 B.n260 VSUBS 0.006864f
C321 B.n261 VSUBS 0.006864f
C322 B.n262 VSUBS 0.006864f
C323 B.n263 VSUBS 0.006864f
C324 B.n264 VSUBS 0.006864f
C325 B.n265 VSUBS 0.006864f
C326 B.n266 VSUBS 0.006864f
C327 B.n267 VSUBS 0.006864f
C328 B.n268 VSUBS 0.006864f
C329 B.n269 VSUBS 0.006864f
C330 B.n270 VSUBS 0.006864f
C331 B.n271 VSUBS 0.006864f
C332 B.n272 VSUBS 0.006864f
C333 B.n273 VSUBS 0.006864f
C334 B.n274 VSUBS 0.006864f
C335 B.n275 VSUBS 0.006864f
C336 B.n276 VSUBS 0.006864f
C337 B.n277 VSUBS 0.006864f
C338 B.n278 VSUBS 0.006864f
C339 B.n279 VSUBS 0.006864f
C340 B.n280 VSUBS 0.00646f
C341 B.n281 VSUBS 0.015902f
C342 B.n282 VSUBS 0.003836f
C343 B.n283 VSUBS 0.006864f
C344 B.n284 VSUBS 0.006864f
C345 B.n285 VSUBS 0.006864f
C346 B.n286 VSUBS 0.006864f
C347 B.n287 VSUBS 0.006864f
C348 B.n288 VSUBS 0.006864f
C349 B.n289 VSUBS 0.006864f
C350 B.n290 VSUBS 0.006864f
C351 B.n291 VSUBS 0.006864f
C352 B.n292 VSUBS 0.006864f
C353 B.n293 VSUBS 0.006864f
C354 B.n294 VSUBS 0.006864f
C355 B.t5 VSUBS 0.449974f
C356 B.t4 VSUBS 0.466461f
C357 B.t3 VSUBS 1.1791f
C358 B.n295 VSUBS 0.225982f
C359 B.n296 VSUBS 0.067915f
C360 B.n297 VSUBS 0.015902f
C361 B.n298 VSUBS 0.003836f
C362 B.n299 VSUBS 0.006864f
C363 B.n300 VSUBS 0.006864f
C364 B.n301 VSUBS 0.006864f
C365 B.n302 VSUBS 0.006864f
C366 B.n303 VSUBS 0.006864f
C367 B.n304 VSUBS 0.006864f
C368 B.n305 VSUBS 0.006864f
C369 B.n306 VSUBS 0.006864f
C370 B.n307 VSUBS 0.006864f
C371 B.n308 VSUBS 0.006864f
C372 B.n309 VSUBS 0.006864f
C373 B.n310 VSUBS 0.006864f
C374 B.n311 VSUBS 0.006864f
C375 B.n312 VSUBS 0.006864f
C376 B.n313 VSUBS 0.006864f
C377 B.n314 VSUBS 0.006864f
C378 B.n315 VSUBS 0.006864f
C379 B.n316 VSUBS 0.006864f
C380 B.n317 VSUBS 0.006864f
C381 B.n318 VSUBS 0.006864f
C382 B.n319 VSUBS 0.006864f
C383 B.n320 VSUBS 0.006864f
C384 B.n321 VSUBS 0.006864f
C385 B.n322 VSUBS 0.006864f
C386 B.n323 VSUBS 0.006864f
C387 B.n324 VSUBS 0.006864f
C388 B.n325 VSUBS 0.006864f
C389 B.n326 VSUBS 0.006864f
C390 B.n327 VSUBS 0.006864f
C391 B.n328 VSUBS 0.006864f
C392 B.n329 VSUBS 0.006864f
C393 B.n330 VSUBS 0.006864f
C394 B.n331 VSUBS 0.006864f
C395 B.n332 VSUBS 0.006864f
C396 B.n333 VSUBS 0.006864f
C397 B.n334 VSUBS 0.006864f
C398 B.n335 VSUBS 0.006864f
C399 B.n336 VSUBS 0.006864f
C400 B.n337 VSUBS 0.006864f
C401 B.n338 VSUBS 0.006864f
C402 B.n339 VSUBS 0.006864f
C403 B.n340 VSUBS 0.006864f
C404 B.n341 VSUBS 0.006864f
C405 B.n342 VSUBS 0.006864f
C406 B.n343 VSUBS 0.006864f
C407 B.n344 VSUBS 0.006864f
C408 B.n345 VSUBS 0.006864f
C409 B.n346 VSUBS 0.006864f
C410 B.n347 VSUBS 0.006864f
C411 B.n348 VSUBS 0.006864f
C412 B.n349 VSUBS 0.006864f
C413 B.n350 VSUBS 0.006864f
C414 B.n351 VSUBS 0.006864f
C415 B.n352 VSUBS 0.006864f
C416 B.n353 VSUBS 0.006864f
C417 B.n354 VSUBS 0.006864f
C418 B.n355 VSUBS 0.006864f
C419 B.n356 VSUBS 0.006864f
C420 B.n357 VSUBS 0.006864f
C421 B.n358 VSUBS 0.006864f
C422 B.n359 VSUBS 0.006864f
C423 B.n360 VSUBS 0.006864f
C424 B.n361 VSUBS 0.006864f
C425 B.n362 VSUBS 0.006864f
C426 B.n363 VSUBS 0.006864f
C427 B.n364 VSUBS 0.006864f
C428 B.n365 VSUBS 0.006864f
C429 B.n366 VSUBS 0.006864f
C430 B.n367 VSUBS 0.006864f
C431 B.n368 VSUBS 0.006864f
C432 B.n369 VSUBS 0.014588f
C433 B.n370 VSUBS 0.015693f
C434 B.n371 VSUBS 0.014805f
C435 B.n372 VSUBS 0.006864f
C436 B.n373 VSUBS 0.006864f
C437 B.n374 VSUBS 0.006864f
C438 B.n375 VSUBS 0.006864f
C439 B.n376 VSUBS 0.006864f
C440 B.n377 VSUBS 0.006864f
C441 B.n378 VSUBS 0.006864f
C442 B.n379 VSUBS 0.006864f
C443 B.n380 VSUBS 0.006864f
C444 B.n381 VSUBS 0.006864f
C445 B.n382 VSUBS 0.006864f
C446 B.n383 VSUBS 0.006864f
C447 B.n384 VSUBS 0.006864f
C448 B.n385 VSUBS 0.006864f
C449 B.n386 VSUBS 0.006864f
C450 B.n387 VSUBS 0.006864f
C451 B.n388 VSUBS 0.006864f
C452 B.n389 VSUBS 0.006864f
C453 B.n390 VSUBS 0.006864f
C454 B.n391 VSUBS 0.006864f
C455 B.n392 VSUBS 0.006864f
C456 B.n393 VSUBS 0.006864f
C457 B.n394 VSUBS 0.006864f
C458 B.n395 VSUBS 0.006864f
C459 B.n396 VSUBS 0.006864f
C460 B.n397 VSUBS 0.006864f
C461 B.n398 VSUBS 0.006864f
C462 B.n399 VSUBS 0.006864f
C463 B.n400 VSUBS 0.006864f
C464 B.n401 VSUBS 0.006864f
C465 B.n402 VSUBS 0.006864f
C466 B.n403 VSUBS 0.006864f
C467 B.n404 VSUBS 0.006864f
C468 B.n405 VSUBS 0.006864f
C469 B.n406 VSUBS 0.006864f
C470 B.n407 VSUBS 0.006864f
C471 B.n408 VSUBS 0.006864f
C472 B.n409 VSUBS 0.006864f
C473 B.n410 VSUBS 0.006864f
C474 B.n411 VSUBS 0.006864f
C475 B.n412 VSUBS 0.006864f
C476 B.n413 VSUBS 0.006864f
C477 B.n414 VSUBS 0.006864f
C478 B.n415 VSUBS 0.006864f
C479 B.n416 VSUBS 0.006864f
C480 B.n417 VSUBS 0.006864f
C481 B.n418 VSUBS 0.006864f
C482 B.n419 VSUBS 0.006864f
C483 B.n420 VSUBS 0.006864f
C484 B.n421 VSUBS 0.006864f
C485 B.n422 VSUBS 0.006864f
C486 B.n423 VSUBS 0.006864f
C487 B.n424 VSUBS 0.006864f
C488 B.n425 VSUBS 0.006864f
C489 B.n426 VSUBS 0.006864f
C490 B.n427 VSUBS 0.006864f
C491 B.n428 VSUBS 0.006864f
C492 B.n429 VSUBS 0.006864f
C493 B.n430 VSUBS 0.006864f
C494 B.n431 VSUBS 0.006864f
C495 B.n432 VSUBS 0.006864f
C496 B.n433 VSUBS 0.006864f
C497 B.n434 VSUBS 0.006864f
C498 B.n435 VSUBS 0.006864f
C499 B.n436 VSUBS 0.006864f
C500 B.n437 VSUBS 0.006864f
C501 B.n438 VSUBS 0.006864f
C502 B.n439 VSUBS 0.006864f
C503 B.n440 VSUBS 0.006864f
C504 B.n441 VSUBS 0.006864f
C505 B.n442 VSUBS 0.006864f
C506 B.n443 VSUBS 0.006864f
C507 B.n444 VSUBS 0.006864f
C508 B.n445 VSUBS 0.006864f
C509 B.n446 VSUBS 0.006864f
C510 B.n447 VSUBS 0.006864f
C511 B.n448 VSUBS 0.006864f
C512 B.n449 VSUBS 0.006864f
C513 B.n450 VSUBS 0.006864f
C514 B.n451 VSUBS 0.006864f
C515 B.n452 VSUBS 0.006864f
C516 B.n453 VSUBS 0.006864f
C517 B.n454 VSUBS 0.006864f
C518 B.n455 VSUBS 0.006864f
C519 B.n456 VSUBS 0.014805f
C520 B.n457 VSUBS 0.015476f
C521 B.n458 VSUBS 0.015476f
C522 B.n459 VSUBS 0.006864f
C523 B.n460 VSUBS 0.006864f
C524 B.n461 VSUBS 0.006864f
C525 B.n462 VSUBS 0.006864f
C526 B.n463 VSUBS 0.006864f
C527 B.n464 VSUBS 0.006864f
C528 B.n465 VSUBS 0.006864f
C529 B.n466 VSUBS 0.006864f
C530 B.n467 VSUBS 0.006864f
C531 B.n468 VSUBS 0.006864f
C532 B.n469 VSUBS 0.006864f
C533 B.n470 VSUBS 0.006864f
C534 B.n471 VSUBS 0.006864f
C535 B.n472 VSUBS 0.006864f
C536 B.n473 VSUBS 0.006864f
C537 B.n474 VSUBS 0.006864f
C538 B.n475 VSUBS 0.006864f
C539 B.n476 VSUBS 0.006864f
C540 B.n477 VSUBS 0.006864f
C541 B.n478 VSUBS 0.006864f
C542 B.n479 VSUBS 0.006864f
C543 B.n480 VSUBS 0.006864f
C544 B.n481 VSUBS 0.006864f
C545 B.n482 VSUBS 0.006864f
C546 B.n483 VSUBS 0.006864f
C547 B.n484 VSUBS 0.006864f
C548 B.n485 VSUBS 0.006864f
C549 B.n486 VSUBS 0.006864f
C550 B.n487 VSUBS 0.006864f
C551 B.n488 VSUBS 0.006864f
C552 B.n489 VSUBS 0.006864f
C553 B.n490 VSUBS 0.006864f
C554 B.n491 VSUBS 0.006864f
C555 B.n492 VSUBS 0.006864f
C556 B.n493 VSUBS 0.006864f
C557 B.n494 VSUBS 0.006864f
C558 B.n495 VSUBS 0.006864f
C559 B.n496 VSUBS 0.006864f
C560 B.n497 VSUBS 0.006864f
C561 B.n498 VSUBS 0.006864f
C562 B.n499 VSUBS 0.006864f
C563 B.n500 VSUBS 0.006864f
C564 B.n501 VSUBS 0.006864f
C565 B.n502 VSUBS 0.006864f
C566 B.n503 VSUBS 0.006864f
C567 B.n504 VSUBS 0.006864f
C568 B.n505 VSUBS 0.006864f
C569 B.n506 VSUBS 0.006864f
C570 B.n507 VSUBS 0.006864f
C571 B.n508 VSUBS 0.006864f
C572 B.n509 VSUBS 0.006864f
C573 B.n510 VSUBS 0.006864f
C574 B.n511 VSUBS 0.006864f
C575 B.n512 VSUBS 0.006864f
C576 B.n513 VSUBS 0.006864f
C577 B.n514 VSUBS 0.006864f
C578 B.n515 VSUBS 0.006864f
C579 B.n516 VSUBS 0.006864f
C580 B.n517 VSUBS 0.006864f
C581 B.n518 VSUBS 0.006864f
C582 B.n519 VSUBS 0.006864f
C583 B.n520 VSUBS 0.006864f
C584 B.n521 VSUBS 0.006864f
C585 B.n522 VSUBS 0.006864f
C586 B.n523 VSUBS 0.006864f
C587 B.n524 VSUBS 0.006864f
C588 B.n525 VSUBS 0.006864f
C589 B.n526 VSUBS 0.00646f
C590 B.n527 VSUBS 0.006864f
C591 B.n528 VSUBS 0.006864f
C592 B.n529 VSUBS 0.006864f
C593 B.n530 VSUBS 0.006864f
C594 B.n531 VSUBS 0.006864f
C595 B.n532 VSUBS 0.006864f
C596 B.n533 VSUBS 0.006864f
C597 B.n534 VSUBS 0.006864f
C598 B.n535 VSUBS 0.006864f
C599 B.n536 VSUBS 0.006864f
C600 B.n537 VSUBS 0.006864f
C601 B.n538 VSUBS 0.006864f
C602 B.n539 VSUBS 0.006864f
C603 B.n540 VSUBS 0.006864f
C604 B.n541 VSUBS 0.006864f
C605 B.n542 VSUBS 0.003836f
C606 B.n543 VSUBS 0.015902f
C607 B.n544 VSUBS 0.00646f
C608 B.n545 VSUBS 0.006864f
C609 B.n546 VSUBS 0.006864f
C610 B.n547 VSUBS 0.006864f
C611 B.n548 VSUBS 0.006864f
C612 B.n549 VSUBS 0.006864f
C613 B.n550 VSUBS 0.006864f
C614 B.n551 VSUBS 0.006864f
C615 B.n552 VSUBS 0.006864f
C616 B.n553 VSUBS 0.006864f
C617 B.n554 VSUBS 0.006864f
C618 B.n555 VSUBS 0.006864f
C619 B.n556 VSUBS 0.006864f
C620 B.n557 VSUBS 0.006864f
C621 B.n558 VSUBS 0.006864f
C622 B.n559 VSUBS 0.006864f
C623 B.n560 VSUBS 0.006864f
C624 B.n561 VSUBS 0.006864f
C625 B.n562 VSUBS 0.006864f
C626 B.n563 VSUBS 0.006864f
C627 B.n564 VSUBS 0.006864f
C628 B.n565 VSUBS 0.006864f
C629 B.n566 VSUBS 0.006864f
C630 B.n567 VSUBS 0.006864f
C631 B.n568 VSUBS 0.006864f
C632 B.n569 VSUBS 0.006864f
C633 B.n570 VSUBS 0.006864f
C634 B.n571 VSUBS 0.006864f
C635 B.n572 VSUBS 0.006864f
C636 B.n573 VSUBS 0.006864f
C637 B.n574 VSUBS 0.006864f
C638 B.n575 VSUBS 0.006864f
C639 B.n576 VSUBS 0.006864f
C640 B.n577 VSUBS 0.006864f
C641 B.n578 VSUBS 0.006864f
C642 B.n579 VSUBS 0.006864f
C643 B.n580 VSUBS 0.006864f
C644 B.n581 VSUBS 0.006864f
C645 B.n582 VSUBS 0.006864f
C646 B.n583 VSUBS 0.006864f
C647 B.n584 VSUBS 0.006864f
C648 B.n585 VSUBS 0.006864f
C649 B.n586 VSUBS 0.006864f
C650 B.n587 VSUBS 0.006864f
C651 B.n588 VSUBS 0.006864f
C652 B.n589 VSUBS 0.006864f
C653 B.n590 VSUBS 0.006864f
C654 B.n591 VSUBS 0.006864f
C655 B.n592 VSUBS 0.006864f
C656 B.n593 VSUBS 0.006864f
C657 B.n594 VSUBS 0.006864f
C658 B.n595 VSUBS 0.006864f
C659 B.n596 VSUBS 0.006864f
C660 B.n597 VSUBS 0.006864f
C661 B.n598 VSUBS 0.006864f
C662 B.n599 VSUBS 0.006864f
C663 B.n600 VSUBS 0.006864f
C664 B.n601 VSUBS 0.006864f
C665 B.n602 VSUBS 0.006864f
C666 B.n603 VSUBS 0.006864f
C667 B.n604 VSUBS 0.006864f
C668 B.n605 VSUBS 0.006864f
C669 B.n606 VSUBS 0.006864f
C670 B.n607 VSUBS 0.006864f
C671 B.n608 VSUBS 0.006864f
C672 B.n609 VSUBS 0.006864f
C673 B.n610 VSUBS 0.006864f
C674 B.n611 VSUBS 0.006864f
C675 B.n612 VSUBS 0.006864f
C676 B.n613 VSUBS 0.015476f
C677 B.n614 VSUBS 0.014805f
C678 B.n615 VSUBS 0.014805f
C679 B.n616 VSUBS 0.006864f
C680 B.n617 VSUBS 0.006864f
C681 B.n618 VSUBS 0.006864f
C682 B.n619 VSUBS 0.006864f
C683 B.n620 VSUBS 0.006864f
C684 B.n621 VSUBS 0.006864f
C685 B.n622 VSUBS 0.006864f
C686 B.n623 VSUBS 0.006864f
C687 B.n624 VSUBS 0.006864f
C688 B.n625 VSUBS 0.006864f
C689 B.n626 VSUBS 0.006864f
C690 B.n627 VSUBS 0.006864f
C691 B.n628 VSUBS 0.006864f
C692 B.n629 VSUBS 0.006864f
C693 B.n630 VSUBS 0.006864f
C694 B.n631 VSUBS 0.006864f
C695 B.n632 VSUBS 0.006864f
C696 B.n633 VSUBS 0.006864f
C697 B.n634 VSUBS 0.006864f
C698 B.n635 VSUBS 0.006864f
C699 B.n636 VSUBS 0.006864f
C700 B.n637 VSUBS 0.006864f
C701 B.n638 VSUBS 0.006864f
C702 B.n639 VSUBS 0.006864f
C703 B.n640 VSUBS 0.006864f
C704 B.n641 VSUBS 0.006864f
C705 B.n642 VSUBS 0.006864f
C706 B.n643 VSUBS 0.006864f
C707 B.n644 VSUBS 0.006864f
C708 B.n645 VSUBS 0.006864f
C709 B.n646 VSUBS 0.006864f
C710 B.n647 VSUBS 0.006864f
C711 B.n648 VSUBS 0.006864f
C712 B.n649 VSUBS 0.006864f
C713 B.n650 VSUBS 0.006864f
C714 B.n651 VSUBS 0.006864f
C715 B.n652 VSUBS 0.006864f
C716 B.n653 VSUBS 0.006864f
C717 B.n654 VSUBS 0.006864f
C718 B.n655 VSUBS 0.008957f
C719 B.n656 VSUBS 0.009541f
C720 B.n657 VSUBS 0.018973f
C721 VDD2.t2 VSUBS 0.289843f
C722 VDD2.t3 VSUBS 0.289843f
C723 VDD2.n0 VSUBS 3.05873f
C724 VDD2.t0 VSUBS 0.289843f
C725 VDD2.t1 VSUBS 0.289843f
C726 VDD2.n1 VSUBS 2.31145f
C727 VDD2.n2 VSUBS 4.29667f
C728 VTAIL.t5 VSUBS 2.43647f
C729 VTAIL.n0 VSUBS 0.748902f
C730 VTAIL.t0 VSUBS 2.43647f
C731 VTAIL.n1 VSUBS 0.816834f
C732 VTAIL.t1 VSUBS 2.43647f
C733 VTAIL.n2 VSUBS 2.11022f
C734 VTAIL.t7 VSUBS 2.43649f
C735 VTAIL.n3 VSUBS 2.11021f
C736 VTAIL.t4 VSUBS 2.43649f
C737 VTAIL.n4 VSUBS 0.816817f
C738 VTAIL.t3 VSUBS 2.43649f
C739 VTAIL.n5 VSUBS 0.816817f
C740 VTAIL.t2 VSUBS 2.43648f
C741 VTAIL.n6 VSUBS 2.11021f
C742 VTAIL.t6 VSUBS 2.43647f
C743 VTAIL.n7 VSUBS 2.03378f
C744 VN.t1 VSUBS 2.95315f
C745 VN.t0 VSUBS 2.95015f
C746 VN.n0 VSUBS 2.02144f
C747 VN.t2 VSUBS 2.95315f
C748 VN.t3 VSUBS 2.95015f
C749 VN.n1 VSUBS 3.7951f
.ends

