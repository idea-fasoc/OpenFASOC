* NGSPICE file created from diff_pair_sample_1317.ext - technology: sky130A

.subckt diff_pair_sample_1317 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=0 ps=0 w=11.94 l=2.53
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=4.6566 ps=24.66 w=11.94 l=2.53
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=4.6566 ps=24.66 w=11.94 l=2.53
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=4.6566 ps=24.66 w=11.94 l=2.53
X4 B.t8 B.t6 B.t7 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=0 ps=0 w=11.94 l=2.53
X5 B.t5 B.t3 B.t4 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=0 ps=0 w=11.94 l=2.53
X6 B.t2 B.t0 B.t1 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=0 ps=0 w=11.94 l=2.53
X7 VDD1.t0 VP.t1 VTAIL.t2 w_n2114_n3356# sky130_fd_pr__pfet_01v8 ad=4.6566 pd=24.66 as=4.6566 ps=24.66 w=11.94 l=2.53
R0 B.n406 B.n405 585
R1 B.n407 B.n64 585
R2 B.n409 B.n408 585
R3 B.n410 B.n63 585
R4 B.n412 B.n411 585
R5 B.n413 B.n62 585
R6 B.n415 B.n414 585
R7 B.n416 B.n61 585
R8 B.n418 B.n417 585
R9 B.n419 B.n60 585
R10 B.n421 B.n420 585
R11 B.n422 B.n59 585
R12 B.n424 B.n423 585
R13 B.n425 B.n58 585
R14 B.n427 B.n426 585
R15 B.n428 B.n57 585
R16 B.n430 B.n429 585
R17 B.n431 B.n56 585
R18 B.n433 B.n432 585
R19 B.n434 B.n55 585
R20 B.n436 B.n435 585
R21 B.n437 B.n54 585
R22 B.n439 B.n438 585
R23 B.n440 B.n53 585
R24 B.n442 B.n441 585
R25 B.n443 B.n52 585
R26 B.n445 B.n444 585
R27 B.n446 B.n51 585
R28 B.n448 B.n447 585
R29 B.n449 B.n50 585
R30 B.n451 B.n450 585
R31 B.n452 B.n49 585
R32 B.n454 B.n453 585
R33 B.n455 B.n48 585
R34 B.n457 B.n456 585
R35 B.n458 B.n47 585
R36 B.n460 B.n459 585
R37 B.n461 B.n46 585
R38 B.n463 B.n462 585
R39 B.n464 B.n45 585
R40 B.n466 B.n465 585
R41 B.n468 B.n467 585
R42 B.n469 B.n41 585
R43 B.n471 B.n470 585
R44 B.n472 B.n40 585
R45 B.n474 B.n473 585
R46 B.n475 B.n39 585
R47 B.n477 B.n476 585
R48 B.n478 B.n38 585
R49 B.n480 B.n479 585
R50 B.n481 B.n35 585
R51 B.n484 B.n483 585
R52 B.n485 B.n34 585
R53 B.n487 B.n486 585
R54 B.n488 B.n33 585
R55 B.n490 B.n489 585
R56 B.n491 B.n32 585
R57 B.n493 B.n492 585
R58 B.n494 B.n31 585
R59 B.n496 B.n495 585
R60 B.n497 B.n30 585
R61 B.n499 B.n498 585
R62 B.n500 B.n29 585
R63 B.n502 B.n501 585
R64 B.n503 B.n28 585
R65 B.n505 B.n504 585
R66 B.n506 B.n27 585
R67 B.n508 B.n507 585
R68 B.n509 B.n26 585
R69 B.n511 B.n510 585
R70 B.n512 B.n25 585
R71 B.n514 B.n513 585
R72 B.n515 B.n24 585
R73 B.n517 B.n516 585
R74 B.n518 B.n23 585
R75 B.n520 B.n519 585
R76 B.n521 B.n22 585
R77 B.n523 B.n522 585
R78 B.n524 B.n21 585
R79 B.n526 B.n525 585
R80 B.n527 B.n20 585
R81 B.n529 B.n528 585
R82 B.n530 B.n19 585
R83 B.n532 B.n531 585
R84 B.n533 B.n18 585
R85 B.n535 B.n534 585
R86 B.n536 B.n17 585
R87 B.n538 B.n537 585
R88 B.n539 B.n16 585
R89 B.n541 B.n540 585
R90 B.n542 B.n15 585
R91 B.n544 B.n543 585
R92 B.n404 B.n65 585
R93 B.n403 B.n402 585
R94 B.n401 B.n66 585
R95 B.n400 B.n399 585
R96 B.n398 B.n67 585
R97 B.n397 B.n396 585
R98 B.n395 B.n68 585
R99 B.n394 B.n393 585
R100 B.n392 B.n69 585
R101 B.n391 B.n390 585
R102 B.n389 B.n70 585
R103 B.n388 B.n387 585
R104 B.n386 B.n71 585
R105 B.n385 B.n384 585
R106 B.n383 B.n72 585
R107 B.n382 B.n381 585
R108 B.n380 B.n73 585
R109 B.n379 B.n378 585
R110 B.n377 B.n74 585
R111 B.n376 B.n375 585
R112 B.n374 B.n75 585
R113 B.n373 B.n372 585
R114 B.n371 B.n76 585
R115 B.n370 B.n369 585
R116 B.n368 B.n77 585
R117 B.n367 B.n366 585
R118 B.n365 B.n78 585
R119 B.n364 B.n363 585
R120 B.n362 B.n79 585
R121 B.n361 B.n360 585
R122 B.n359 B.n80 585
R123 B.n358 B.n357 585
R124 B.n356 B.n81 585
R125 B.n355 B.n354 585
R126 B.n353 B.n82 585
R127 B.n352 B.n351 585
R128 B.n350 B.n83 585
R129 B.n349 B.n348 585
R130 B.n347 B.n84 585
R131 B.n346 B.n345 585
R132 B.n344 B.n85 585
R133 B.n343 B.n342 585
R134 B.n341 B.n86 585
R135 B.n340 B.n339 585
R136 B.n338 B.n87 585
R137 B.n337 B.n336 585
R138 B.n335 B.n88 585
R139 B.n334 B.n333 585
R140 B.n332 B.n89 585
R141 B.n331 B.n330 585
R142 B.n329 B.n90 585
R143 B.n190 B.n189 585
R144 B.n191 B.n140 585
R145 B.n193 B.n192 585
R146 B.n194 B.n139 585
R147 B.n196 B.n195 585
R148 B.n197 B.n138 585
R149 B.n199 B.n198 585
R150 B.n200 B.n137 585
R151 B.n202 B.n201 585
R152 B.n203 B.n136 585
R153 B.n205 B.n204 585
R154 B.n206 B.n135 585
R155 B.n208 B.n207 585
R156 B.n209 B.n134 585
R157 B.n211 B.n210 585
R158 B.n212 B.n133 585
R159 B.n214 B.n213 585
R160 B.n215 B.n132 585
R161 B.n217 B.n216 585
R162 B.n218 B.n131 585
R163 B.n220 B.n219 585
R164 B.n221 B.n130 585
R165 B.n223 B.n222 585
R166 B.n224 B.n129 585
R167 B.n226 B.n225 585
R168 B.n227 B.n128 585
R169 B.n229 B.n228 585
R170 B.n230 B.n127 585
R171 B.n232 B.n231 585
R172 B.n233 B.n126 585
R173 B.n235 B.n234 585
R174 B.n236 B.n125 585
R175 B.n238 B.n237 585
R176 B.n239 B.n124 585
R177 B.n241 B.n240 585
R178 B.n242 B.n123 585
R179 B.n244 B.n243 585
R180 B.n245 B.n122 585
R181 B.n247 B.n246 585
R182 B.n248 B.n121 585
R183 B.n250 B.n249 585
R184 B.n252 B.n251 585
R185 B.n253 B.n117 585
R186 B.n255 B.n254 585
R187 B.n256 B.n116 585
R188 B.n258 B.n257 585
R189 B.n259 B.n115 585
R190 B.n261 B.n260 585
R191 B.n262 B.n114 585
R192 B.n264 B.n263 585
R193 B.n265 B.n111 585
R194 B.n268 B.n267 585
R195 B.n269 B.n110 585
R196 B.n271 B.n270 585
R197 B.n272 B.n109 585
R198 B.n274 B.n273 585
R199 B.n275 B.n108 585
R200 B.n277 B.n276 585
R201 B.n278 B.n107 585
R202 B.n280 B.n279 585
R203 B.n281 B.n106 585
R204 B.n283 B.n282 585
R205 B.n284 B.n105 585
R206 B.n286 B.n285 585
R207 B.n287 B.n104 585
R208 B.n289 B.n288 585
R209 B.n290 B.n103 585
R210 B.n292 B.n291 585
R211 B.n293 B.n102 585
R212 B.n295 B.n294 585
R213 B.n296 B.n101 585
R214 B.n298 B.n297 585
R215 B.n299 B.n100 585
R216 B.n301 B.n300 585
R217 B.n302 B.n99 585
R218 B.n304 B.n303 585
R219 B.n305 B.n98 585
R220 B.n307 B.n306 585
R221 B.n308 B.n97 585
R222 B.n310 B.n309 585
R223 B.n311 B.n96 585
R224 B.n313 B.n312 585
R225 B.n314 B.n95 585
R226 B.n316 B.n315 585
R227 B.n317 B.n94 585
R228 B.n319 B.n318 585
R229 B.n320 B.n93 585
R230 B.n322 B.n321 585
R231 B.n323 B.n92 585
R232 B.n325 B.n324 585
R233 B.n326 B.n91 585
R234 B.n328 B.n327 585
R235 B.n188 B.n141 585
R236 B.n187 B.n186 585
R237 B.n185 B.n142 585
R238 B.n184 B.n183 585
R239 B.n182 B.n143 585
R240 B.n181 B.n180 585
R241 B.n179 B.n144 585
R242 B.n178 B.n177 585
R243 B.n176 B.n145 585
R244 B.n175 B.n174 585
R245 B.n173 B.n146 585
R246 B.n172 B.n171 585
R247 B.n170 B.n147 585
R248 B.n169 B.n168 585
R249 B.n167 B.n148 585
R250 B.n166 B.n165 585
R251 B.n164 B.n149 585
R252 B.n163 B.n162 585
R253 B.n161 B.n150 585
R254 B.n160 B.n159 585
R255 B.n158 B.n151 585
R256 B.n157 B.n156 585
R257 B.n155 B.n152 585
R258 B.n154 B.n153 585
R259 B.n2 B.n0 585
R260 B.n581 B.n1 585
R261 B.n580 B.n579 585
R262 B.n578 B.n3 585
R263 B.n577 B.n576 585
R264 B.n575 B.n4 585
R265 B.n574 B.n573 585
R266 B.n572 B.n5 585
R267 B.n571 B.n570 585
R268 B.n569 B.n6 585
R269 B.n568 B.n567 585
R270 B.n566 B.n7 585
R271 B.n565 B.n564 585
R272 B.n563 B.n8 585
R273 B.n562 B.n561 585
R274 B.n560 B.n9 585
R275 B.n559 B.n558 585
R276 B.n557 B.n10 585
R277 B.n556 B.n555 585
R278 B.n554 B.n11 585
R279 B.n553 B.n552 585
R280 B.n551 B.n12 585
R281 B.n550 B.n549 585
R282 B.n548 B.n13 585
R283 B.n547 B.n546 585
R284 B.n545 B.n14 585
R285 B.n583 B.n582 585
R286 B.n190 B.n141 526.135
R287 B.n545 B.n544 526.135
R288 B.n329 B.n328 526.135
R289 B.n406 B.n65 526.135
R290 B.n112 B.t2 429.834
R291 B.n42 B.t4 429.834
R292 B.n118 B.t11 429.832
R293 B.n36 B.t7 429.832
R294 B.n113 B.t1 374.366
R295 B.n43 B.t5 374.366
R296 B.n119 B.t10 374.366
R297 B.n37 B.t8 374.366
R298 B.n112 B.t0 321.675
R299 B.n118 B.t9 321.675
R300 B.n36 B.t6 321.675
R301 B.n42 B.t3 321.675
R302 B.n186 B.n141 163.367
R303 B.n186 B.n185 163.367
R304 B.n185 B.n184 163.367
R305 B.n184 B.n143 163.367
R306 B.n180 B.n143 163.367
R307 B.n180 B.n179 163.367
R308 B.n179 B.n178 163.367
R309 B.n178 B.n145 163.367
R310 B.n174 B.n145 163.367
R311 B.n174 B.n173 163.367
R312 B.n173 B.n172 163.367
R313 B.n172 B.n147 163.367
R314 B.n168 B.n147 163.367
R315 B.n168 B.n167 163.367
R316 B.n167 B.n166 163.367
R317 B.n166 B.n149 163.367
R318 B.n162 B.n149 163.367
R319 B.n162 B.n161 163.367
R320 B.n161 B.n160 163.367
R321 B.n160 B.n151 163.367
R322 B.n156 B.n151 163.367
R323 B.n156 B.n155 163.367
R324 B.n155 B.n154 163.367
R325 B.n154 B.n2 163.367
R326 B.n582 B.n2 163.367
R327 B.n582 B.n581 163.367
R328 B.n581 B.n580 163.367
R329 B.n580 B.n3 163.367
R330 B.n576 B.n3 163.367
R331 B.n576 B.n575 163.367
R332 B.n575 B.n574 163.367
R333 B.n574 B.n5 163.367
R334 B.n570 B.n5 163.367
R335 B.n570 B.n569 163.367
R336 B.n569 B.n568 163.367
R337 B.n568 B.n7 163.367
R338 B.n564 B.n7 163.367
R339 B.n564 B.n563 163.367
R340 B.n563 B.n562 163.367
R341 B.n562 B.n9 163.367
R342 B.n558 B.n9 163.367
R343 B.n558 B.n557 163.367
R344 B.n557 B.n556 163.367
R345 B.n556 B.n11 163.367
R346 B.n552 B.n11 163.367
R347 B.n552 B.n551 163.367
R348 B.n551 B.n550 163.367
R349 B.n550 B.n13 163.367
R350 B.n546 B.n13 163.367
R351 B.n546 B.n545 163.367
R352 B.n191 B.n190 163.367
R353 B.n192 B.n191 163.367
R354 B.n192 B.n139 163.367
R355 B.n196 B.n139 163.367
R356 B.n197 B.n196 163.367
R357 B.n198 B.n197 163.367
R358 B.n198 B.n137 163.367
R359 B.n202 B.n137 163.367
R360 B.n203 B.n202 163.367
R361 B.n204 B.n203 163.367
R362 B.n204 B.n135 163.367
R363 B.n208 B.n135 163.367
R364 B.n209 B.n208 163.367
R365 B.n210 B.n209 163.367
R366 B.n210 B.n133 163.367
R367 B.n214 B.n133 163.367
R368 B.n215 B.n214 163.367
R369 B.n216 B.n215 163.367
R370 B.n216 B.n131 163.367
R371 B.n220 B.n131 163.367
R372 B.n221 B.n220 163.367
R373 B.n222 B.n221 163.367
R374 B.n222 B.n129 163.367
R375 B.n226 B.n129 163.367
R376 B.n227 B.n226 163.367
R377 B.n228 B.n227 163.367
R378 B.n228 B.n127 163.367
R379 B.n232 B.n127 163.367
R380 B.n233 B.n232 163.367
R381 B.n234 B.n233 163.367
R382 B.n234 B.n125 163.367
R383 B.n238 B.n125 163.367
R384 B.n239 B.n238 163.367
R385 B.n240 B.n239 163.367
R386 B.n240 B.n123 163.367
R387 B.n244 B.n123 163.367
R388 B.n245 B.n244 163.367
R389 B.n246 B.n245 163.367
R390 B.n246 B.n121 163.367
R391 B.n250 B.n121 163.367
R392 B.n251 B.n250 163.367
R393 B.n251 B.n117 163.367
R394 B.n255 B.n117 163.367
R395 B.n256 B.n255 163.367
R396 B.n257 B.n256 163.367
R397 B.n257 B.n115 163.367
R398 B.n261 B.n115 163.367
R399 B.n262 B.n261 163.367
R400 B.n263 B.n262 163.367
R401 B.n263 B.n111 163.367
R402 B.n268 B.n111 163.367
R403 B.n269 B.n268 163.367
R404 B.n270 B.n269 163.367
R405 B.n270 B.n109 163.367
R406 B.n274 B.n109 163.367
R407 B.n275 B.n274 163.367
R408 B.n276 B.n275 163.367
R409 B.n276 B.n107 163.367
R410 B.n280 B.n107 163.367
R411 B.n281 B.n280 163.367
R412 B.n282 B.n281 163.367
R413 B.n282 B.n105 163.367
R414 B.n286 B.n105 163.367
R415 B.n287 B.n286 163.367
R416 B.n288 B.n287 163.367
R417 B.n288 B.n103 163.367
R418 B.n292 B.n103 163.367
R419 B.n293 B.n292 163.367
R420 B.n294 B.n293 163.367
R421 B.n294 B.n101 163.367
R422 B.n298 B.n101 163.367
R423 B.n299 B.n298 163.367
R424 B.n300 B.n299 163.367
R425 B.n300 B.n99 163.367
R426 B.n304 B.n99 163.367
R427 B.n305 B.n304 163.367
R428 B.n306 B.n305 163.367
R429 B.n306 B.n97 163.367
R430 B.n310 B.n97 163.367
R431 B.n311 B.n310 163.367
R432 B.n312 B.n311 163.367
R433 B.n312 B.n95 163.367
R434 B.n316 B.n95 163.367
R435 B.n317 B.n316 163.367
R436 B.n318 B.n317 163.367
R437 B.n318 B.n93 163.367
R438 B.n322 B.n93 163.367
R439 B.n323 B.n322 163.367
R440 B.n324 B.n323 163.367
R441 B.n324 B.n91 163.367
R442 B.n328 B.n91 163.367
R443 B.n330 B.n329 163.367
R444 B.n330 B.n89 163.367
R445 B.n334 B.n89 163.367
R446 B.n335 B.n334 163.367
R447 B.n336 B.n335 163.367
R448 B.n336 B.n87 163.367
R449 B.n340 B.n87 163.367
R450 B.n341 B.n340 163.367
R451 B.n342 B.n341 163.367
R452 B.n342 B.n85 163.367
R453 B.n346 B.n85 163.367
R454 B.n347 B.n346 163.367
R455 B.n348 B.n347 163.367
R456 B.n348 B.n83 163.367
R457 B.n352 B.n83 163.367
R458 B.n353 B.n352 163.367
R459 B.n354 B.n353 163.367
R460 B.n354 B.n81 163.367
R461 B.n358 B.n81 163.367
R462 B.n359 B.n358 163.367
R463 B.n360 B.n359 163.367
R464 B.n360 B.n79 163.367
R465 B.n364 B.n79 163.367
R466 B.n365 B.n364 163.367
R467 B.n366 B.n365 163.367
R468 B.n366 B.n77 163.367
R469 B.n370 B.n77 163.367
R470 B.n371 B.n370 163.367
R471 B.n372 B.n371 163.367
R472 B.n372 B.n75 163.367
R473 B.n376 B.n75 163.367
R474 B.n377 B.n376 163.367
R475 B.n378 B.n377 163.367
R476 B.n378 B.n73 163.367
R477 B.n382 B.n73 163.367
R478 B.n383 B.n382 163.367
R479 B.n384 B.n383 163.367
R480 B.n384 B.n71 163.367
R481 B.n388 B.n71 163.367
R482 B.n389 B.n388 163.367
R483 B.n390 B.n389 163.367
R484 B.n390 B.n69 163.367
R485 B.n394 B.n69 163.367
R486 B.n395 B.n394 163.367
R487 B.n396 B.n395 163.367
R488 B.n396 B.n67 163.367
R489 B.n400 B.n67 163.367
R490 B.n401 B.n400 163.367
R491 B.n402 B.n401 163.367
R492 B.n402 B.n65 163.367
R493 B.n544 B.n15 163.367
R494 B.n540 B.n15 163.367
R495 B.n540 B.n539 163.367
R496 B.n539 B.n538 163.367
R497 B.n538 B.n17 163.367
R498 B.n534 B.n17 163.367
R499 B.n534 B.n533 163.367
R500 B.n533 B.n532 163.367
R501 B.n532 B.n19 163.367
R502 B.n528 B.n19 163.367
R503 B.n528 B.n527 163.367
R504 B.n527 B.n526 163.367
R505 B.n526 B.n21 163.367
R506 B.n522 B.n21 163.367
R507 B.n522 B.n521 163.367
R508 B.n521 B.n520 163.367
R509 B.n520 B.n23 163.367
R510 B.n516 B.n23 163.367
R511 B.n516 B.n515 163.367
R512 B.n515 B.n514 163.367
R513 B.n514 B.n25 163.367
R514 B.n510 B.n25 163.367
R515 B.n510 B.n509 163.367
R516 B.n509 B.n508 163.367
R517 B.n508 B.n27 163.367
R518 B.n504 B.n27 163.367
R519 B.n504 B.n503 163.367
R520 B.n503 B.n502 163.367
R521 B.n502 B.n29 163.367
R522 B.n498 B.n29 163.367
R523 B.n498 B.n497 163.367
R524 B.n497 B.n496 163.367
R525 B.n496 B.n31 163.367
R526 B.n492 B.n31 163.367
R527 B.n492 B.n491 163.367
R528 B.n491 B.n490 163.367
R529 B.n490 B.n33 163.367
R530 B.n486 B.n33 163.367
R531 B.n486 B.n485 163.367
R532 B.n485 B.n484 163.367
R533 B.n484 B.n35 163.367
R534 B.n479 B.n35 163.367
R535 B.n479 B.n478 163.367
R536 B.n478 B.n477 163.367
R537 B.n477 B.n39 163.367
R538 B.n473 B.n39 163.367
R539 B.n473 B.n472 163.367
R540 B.n472 B.n471 163.367
R541 B.n471 B.n41 163.367
R542 B.n467 B.n41 163.367
R543 B.n467 B.n466 163.367
R544 B.n466 B.n45 163.367
R545 B.n462 B.n45 163.367
R546 B.n462 B.n461 163.367
R547 B.n461 B.n460 163.367
R548 B.n460 B.n47 163.367
R549 B.n456 B.n47 163.367
R550 B.n456 B.n455 163.367
R551 B.n455 B.n454 163.367
R552 B.n454 B.n49 163.367
R553 B.n450 B.n49 163.367
R554 B.n450 B.n449 163.367
R555 B.n449 B.n448 163.367
R556 B.n448 B.n51 163.367
R557 B.n444 B.n51 163.367
R558 B.n444 B.n443 163.367
R559 B.n443 B.n442 163.367
R560 B.n442 B.n53 163.367
R561 B.n438 B.n53 163.367
R562 B.n438 B.n437 163.367
R563 B.n437 B.n436 163.367
R564 B.n436 B.n55 163.367
R565 B.n432 B.n55 163.367
R566 B.n432 B.n431 163.367
R567 B.n431 B.n430 163.367
R568 B.n430 B.n57 163.367
R569 B.n426 B.n57 163.367
R570 B.n426 B.n425 163.367
R571 B.n425 B.n424 163.367
R572 B.n424 B.n59 163.367
R573 B.n420 B.n59 163.367
R574 B.n420 B.n419 163.367
R575 B.n419 B.n418 163.367
R576 B.n418 B.n61 163.367
R577 B.n414 B.n61 163.367
R578 B.n414 B.n413 163.367
R579 B.n413 B.n412 163.367
R580 B.n412 B.n63 163.367
R581 B.n408 B.n63 163.367
R582 B.n408 B.n407 163.367
R583 B.n407 B.n406 163.367
R584 B.n266 B.n113 59.5399
R585 B.n120 B.n119 59.5399
R586 B.n482 B.n37 59.5399
R587 B.n44 B.n43 59.5399
R588 B.n113 B.n112 55.4672
R589 B.n119 B.n118 55.4672
R590 B.n37 B.n36 55.4672
R591 B.n43 B.n42 55.4672
R592 B.n543 B.n14 34.1859
R593 B.n405 B.n404 34.1859
R594 B.n327 B.n90 34.1859
R595 B.n189 B.n188 34.1859
R596 B B.n583 18.0485
R597 B.n543 B.n542 10.6151
R598 B.n542 B.n541 10.6151
R599 B.n541 B.n16 10.6151
R600 B.n537 B.n16 10.6151
R601 B.n537 B.n536 10.6151
R602 B.n536 B.n535 10.6151
R603 B.n535 B.n18 10.6151
R604 B.n531 B.n18 10.6151
R605 B.n531 B.n530 10.6151
R606 B.n530 B.n529 10.6151
R607 B.n529 B.n20 10.6151
R608 B.n525 B.n20 10.6151
R609 B.n525 B.n524 10.6151
R610 B.n524 B.n523 10.6151
R611 B.n523 B.n22 10.6151
R612 B.n519 B.n22 10.6151
R613 B.n519 B.n518 10.6151
R614 B.n518 B.n517 10.6151
R615 B.n517 B.n24 10.6151
R616 B.n513 B.n24 10.6151
R617 B.n513 B.n512 10.6151
R618 B.n512 B.n511 10.6151
R619 B.n511 B.n26 10.6151
R620 B.n507 B.n26 10.6151
R621 B.n507 B.n506 10.6151
R622 B.n506 B.n505 10.6151
R623 B.n505 B.n28 10.6151
R624 B.n501 B.n28 10.6151
R625 B.n501 B.n500 10.6151
R626 B.n500 B.n499 10.6151
R627 B.n499 B.n30 10.6151
R628 B.n495 B.n30 10.6151
R629 B.n495 B.n494 10.6151
R630 B.n494 B.n493 10.6151
R631 B.n493 B.n32 10.6151
R632 B.n489 B.n32 10.6151
R633 B.n489 B.n488 10.6151
R634 B.n488 B.n487 10.6151
R635 B.n487 B.n34 10.6151
R636 B.n483 B.n34 10.6151
R637 B.n481 B.n480 10.6151
R638 B.n480 B.n38 10.6151
R639 B.n476 B.n38 10.6151
R640 B.n476 B.n475 10.6151
R641 B.n475 B.n474 10.6151
R642 B.n474 B.n40 10.6151
R643 B.n470 B.n40 10.6151
R644 B.n470 B.n469 10.6151
R645 B.n469 B.n468 10.6151
R646 B.n465 B.n464 10.6151
R647 B.n464 B.n463 10.6151
R648 B.n463 B.n46 10.6151
R649 B.n459 B.n46 10.6151
R650 B.n459 B.n458 10.6151
R651 B.n458 B.n457 10.6151
R652 B.n457 B.n48 10.6151
R653 B.n453 B.n48 10.6151
R654 B.n453 B.n452 10.6151
R655 B.n452 B.n451 10.6151
R656 B.n451 B.n50 10.6151
R657 B.n447 B.n50 10.6151
R658 B.n447 B.n446 10.6151
R659 B.n446 B.n445 10.6151
R660 B.n445 B.n52 10.6151
R661 B.n441 B.n52 10.6151
R662 B.n441 B.n440 10.6151
R663 B.n440 B.n439 10.6151
R664 B.n439 B.n54 10.6151
R665 B.n435 B.n54 10.6151
R666 B.n435 B.n434 10.6151
R667 B.n434 B.n433 10.6151
R668 B.n433 B.n56 10.6151
R669 B.n429 B.n56 10.6151
R670 B.n429 B.n428 10.6151
R671 B.n428 B.n427 10.6151
R672 B.n427 B.n58 10.6151
R673 B.n423 B.n58 10.6151
R674 B.n423 B.n422 10.6151
R675 B.n422 B.n421 10.6151
R676 B.n421 B.n60 10.6151
R677 B.n417 B.n60 10.6151
R678 B.n417 B.n416 10.6151
R679 B.n416 B.n415 10.6151
R680 B.n415 B.n62 10.6151
R681 B.n411 B.n62 10.6151
R682 B.n411 B.n410 10.6151
R683 B.n410 B.n409 10.6151
R684 B.n409 B.n64 10.6151
R685 B.n405 B.n64 10.6151
R686 B.n331 B.n90 10.6151
R687 B.n332 B.n331 10.6151
R688 B.n333 B.n332 10.6151
R689 B.n333 B.n88 10.6151
R690 B.n337 B.n88 10.6151
R691 B.n338 B.n337 10.6151
R692 B.n339 B.n338 10.6151
R693 B.n339 B.n86 10.6151
R694 B.n343 B.n86 10.6151
R695 B.n344 B.n343 10.6151
R696 B.n345 B.n344 10.6151
R697 B.n345 B.n84 10.6151
R698 B.n349 B.n84 10.6151
R699 B.n350 B.n349 10.6151
R700 B.n351 B.n350 10.6151
R701 B.n351 B.n82 10.6151
R702 B.n355 B.n82 10.6151
R703 B.n356 B.n355 10.6151
R704 B.n357 B.n356 10.6151
R705 B.n357 B.n80 10.6151
R706 B.n361 B.n80 10.6151
R707 B.n362 B.n361 10.6151
R708 B.n363 B.n362 10.6151
R709 B.n363 B.n78 10.6151
R710 B.n367 B.n78 10.6151
R711 B.n368 B.n367 10.6151
R712 B.n369 B.n368 10.6151
R713 B.n369 B.n76 10.6151
R714 B.n373 B.n76 10.6151
R715 B.n374 B.n373 10.6151
R716 B.n375 B.n374 10.6151
R717 B.n375 B.n74 10.6151
R718 B.n379 B.n74 10.6151
R719 B.n380 B.n379 10.6151
R720 B.n381 B.n380 10.6151
R721 B.n381 B.n72 10.6151
R722 B.n385 B.n72 10.6151
R723 B.n386 B.n385 10.6151
R724 B.n387 B.n386 10.6151
R725 B.n387 B.n70 10.6151
R726 B.n391 B.n70 10.6151
R727 B.n392 B.n391 10.6151
R728 B.n393 B.n392 10.6151
R729 B.n393 B.n68 10.6151
R730 B.n397 B.n68 10.6151
R731 B.n398 B.n397 10.6151
R732 B.n399 B.n398 10.6151
R733 B.n399 B.n66 10.6151
R734 B.n403 B.n66 10.6151
R735 B.n404 B.n403 10.6151
R736 B.n189 B.n140 10.6151
R737 B.n193 B.n140 10.6151
R738 B.n194 B.n193 10.6151
R739 B.n195 B.n194 10.6151
R740 B.n195 B.n138 10.6151
R741 B.n199 B.n138 10.6151
R742 B.n200 B.n199 10.6151
R743 B.n201 B.n200 10.6151
R744 B.n201 B.n136 10.6151
R745 B.n205 B.n136 10.6151
R746 B.n206 B.n205 10.6151
R747 B.n207 B.n206 10.6151
R748 B.n207 B.n134 10.6151
R749 B.n211 B.n134 10.6151
R750 B.n212 B.n211 10.6151
R751 B.n213 B.n212 10.6151
R752 B.n213 B.n132 10.6151
R753 B.n217 B.n132 10.6151
R754 B.n218 B.n217 10.6151
R755 B.n219 B.n218 10.6151
R756 B.n219 B.n130 10.6151
R757 B.n223 B.n130 10.6151
R758 B.n224 B.n223 10.6151
R759 B.n225 B.n224 10.6151
R760 B.n225 B.n128 10.6151
R761 B.n229 B.n128 10.6151
R762 B.n230 B.n229 10.6151
R763 B.n231 B.n230 10.6151
R764 B.n231 B.n126 10.6151
R765 B.n235 B.n126 10.6151
R766 B.n236 B.n235 10.6151
R767 B.n237 B.n236 10.6151
R768 B.n237 B.n124 10.6151
R769 B.n241 B.n124 10.6151
R770 B.n242 B.n241 10.6151
R771 B.n243 B.n242 10.6151
R772 B.n243 B.n122 10.6151
R773 B.n247 B.n122 10.6151
R774 B.n248 B.n247 10.6151
R775 B.n249 B.n248 10.6151
R776 B.n253 B.n252 10.6151
R777 B.n254 B.n253 10.6151
R778 B.n254 B.n116 10.6151
R779 B.n258 B.n116 10.6151
R780 B.n259 B.n258 10.6151
R781 B.n260 B.n259 10.6151
R782 B.n260 B.n114 10.6151
R783 B.n264 B.n114 10.6151
R784 B.n265 B.n264 10.6151
R785 B.n267 B.n110 10.6151
R786 B.n271 B.n110 10.6151
R787 B.n272 B.n271 10.6151
R788 B.n273 B.n272 10.6151
R789 B.n273 B.n108 10.6151
R790 B.n277 B.n108 10.6151
R791 B.n278 B.n277 10.6151
R792 B.n279 B.n278 10.6151
R793 B.n279 B.n106 10.6151
R794 B.n283 B.n106 10.6151
R795 B.n284 B.n283 10.6151
R796 B.n285 B.n284 10.6151
R797 B.n285 B.n104 10.6151
R798 B.n289 B.n104 10.6151
R799 B.n290 B.n289 10.6151
R800 B.n291 B.n290 10.6151
R801 B.n291 B.n102 10.6151
R802 B.n295 B.n102 10.6151
R803 B.n296 B.n295 10.6151
R804 B.n297 B.n296 10.6151
R805 B.n297 B.n100 10.6151
R806 B.n301 B.n100 10.6151
R807 B.n302 B.n301 10.6151
R808 B.n303 B.n302 10.6151
R809 B.n303 B.n98 10.6151
R810 B.n307 B.n98 10.6151
R811 B.n308 B.n307 10.6151
R812 B.n309 B.n308 10.6151
R813 B.n309 B.n96 10.6151
R814 B.n313 B.n96 10.6151
R815 B.n314 B.n313 10.6151
R816 B.n315 B.n314 10.6151
R817 B.n315 B.n94 10.6151
R818 B.n319 B.n94 10.6151
R819 B.n320 B.n319 10.6151
R820 B.n321 B.n320 10.6151
R821 B.n321 B.n92 10.6151
R822 B.n325 B.n92 10.6151
R823 B.n326 B.n325 10.6151
R824 B.n327 B.n326 10.6151
R825 B.n188 B.n187 10.6151
R826 B.n187 B.n142 10.6151
R827 B.n183 B.n142 10.6151
R828 B.n183 B.n182 10.6151
R829 B.n182 B.n181 10.6151
R830 B.n181 B.n144 10.6151
R831 B.n177 B.n144 10.6151
R832 B.n177 B.n176 10.6151
R833 B.n176 B.n175 10.6151
R834 B.n175 B.n146 10.6151
R835 B.n171 B.n146 10.6151
R836 B.n171 B.n170 10.6151
R837 B.n170 B.n169 10.6151
R838 B.n169 B.n148 10.6151
R839 B.n165 B.n148 10.6151
R840 B.n165 B.n164 10.6151
R841 B.n164 B.n163 10.6151
R842 B.n163 B.n150 10.6151
R843 B.n159 B.n150 10.6151
R844 B.n159 B.n158 10.6151
R845 B.n158 B.n157 10.6151
R846 B.n157 B.n152 10.6151
R847 B.n153 B.n152 10.6151
R848 B.n153 B.n0 10.6151
R849 B.n579 B.n1 10.6151
R850 B.n579 B.n578 10.6151
R851 B.n578 B.n577 10.6151
R852 B.n577 B.n4 10.6151
R853 B.n573 B.n4 10.6151
R854 B.n573 B.n572 10.6151
R855 B.n572 B.n571 10.6151
R856 B.n571 B.n6 10.6151
R857 B.n567 B.n6 10.6151
R858 B.n567 B.n566 10.6151
R859 B.n566 B.n565 10.6151
R860 B.n565 B.n8 10.6151
R861 B.n561 B.n8 10.6151
R862 B.n561 B.n560 10.6151
R863 B.n560 B.n559 10.6151
R864 B.n559 B.n10 10.6151
R865 B.n555 B.n10 10.6151
R866 B.n555 B.n554 10.6151
R867 B.n554 B.n553 10.6151
R868 B.n553 B.n12 10.6151
R869 B.n549 B.n12 10.6151
R870 B.n549 B.n548 10.6151
R871 B.n548 B.n547 10.6151
R872 B.n547 B.n14 10.6151
R873 B.n483 B.n482 9.36635
R874 B.n465 B.n44 9.36635
R875 B.n249 B.n120 9.36635
R876 B.n267 B.n266 9.36635
R877 B.n583 B.n0 2.81026
R878 B.n583 B.n1 2.81026
R879 B.n482 B.n481 1.24928
R880 B.n468 B.n44 1.24928
R881 B.n252 B.n120 1.24928
R882 B.n266 B.n265 1.24928
R883 VP.n0 VP.t1 207.377
R884 VP.n0 VP.t0 162.952
R885 VP VP.n0 0.336784
R886 VTAIL.n262 VTAIL.n261 756.745
R887 VTAIL.n64 VTAIL.n63 756.745
R888 VTAIL.n196 VTAIL.n195 756.745
R889 VTAIL.n130 VTAIL.n129 756.745
R890 VTAIL.n221 VTAIL.n220 585
R891 VTAIL.n223 VTAIL.n222 585
R892 VTAIL.n216 VTAIL.n215 585
R893 VTAIL.n229 VTAIL.n228 585
R894 VTAIL.n231 VTAIL.n230 585
R895 VTAIL.n212 VTAIL.n211 585
R896 VTAIL.n237 VTAIL.n236 585
R897 VTAIL.n239 VTAIL.n238 585
R898 VTAIL.n208 VTAIL.n207 585
R899 VTAIL.n245 VTAIL.n244 585
R900 VTAIL.n247 VTAIL.n246 585
R901 VTAIL.n204 VTAIL.n203 585
R902 VTAIL.n253 VTAIL.n252 585
R903 VTAIL.n255 VTAIL.n254 585
R904 VTAIL.n200 VTAIL.n199 585
R905 VTAIL.n261 VTAIL.n260 585
R906 VTAIL.n23 VTAIL.n22 585
R907 VTAIL.n25 VTAIL.n24 585
R908 VTAIL.n18 VTAIL.n17 585
R909 VTAIL.n31 VTAIL.n30 585
R910 VTAIL.n33 VTAIL.n32 585
R911 VTAIL.n14 VTAIL.n13 585
R912 VTAIL.n39 VTAIL.n38 585
R913 VTAIL.n41 VTAIL.n40 585
R914 VTAIL.n10 VTAIL.n9 585
R915 VTAIL.n47 VTAIL.n46 585
R916 VTAIL.n49 VTAIL.n48 585
R917 VTAIL.n6 VTAIL.n5 585
R918 VTAIL.n55 VTAIL.n54 585
R919 VTAIL.n57 VTAIL.n56 585
R920 VTAIL.n2 VTAIL.n1 585
R921 VTAIL.n63 VTAIL.n62 585
R922 VTAIL.n195 VTAIL.n194 585
R923 VTAIL.n134 VTAIL.n133 585
R924 VTAIL.n189 VTAIL.n188 585
R925 VTAIL.n187 VTAIL.n186 585
R926 VTAIL.n138 VTAIL.n137 585
R927 VTAIL.n181 VTAIL.n180 585
R928 VTAIL.n179 VTAIL.n178 585
R929 VTAIL.n142 VTAIL.n141 585
R930 VTAIL.n173 VTAIL.n172 585
R931 VTAIL.n171 VTAIL.n170 585
R932 VTAIL.n146 VTAIL.n145 585
R933 VTAIL.n165 VTAIL.n164 585
R934 VTAIL.n163 VTAIL.n162 585
R935 VTAIL.n150 VTAIL.n149 585
R936 VTAIL.n157 VTAIL.n156 585
R937 VTAIL.n155 VTAIL.n154 585
R938 VTAIL.n129 VTAIL.n128 585
R939 VTAIL.n68 VTAIL.n67 585
R940 VTAIL.n123 VTAIL.n122 585
R941 VTAIL.n121 VTAIL.n120 585
R942 VTAIL.n72 VTAIL.n71 585
R943 VTAIL.n115 VTAIL.n114 585
R944 VTAIL.n113 VTAIL.n112 585
R945 VTAIL.n76 VTAIL.n75 585
R946 VTAIL.n107 VTAIL.n106 585
R947 VTAIL.n105 VTAIL.n104 585
R948 VTAIL.n80 VTAIL.n79 585
R949 VTAIL.n99 VTAIL.n98 585
R950 VTAIL.n97 VTAIL.n96 585
R951 VTAIL.n84 VTAIL.n83 585
R952 VTAIL.n91 VTAIL.n90 585
R953 VTAIL.n89 VTAIL.n88 585
R954 VTAIL.n153 VTAIL.t2 327.466
R955 VTAIL.n87 VTAIL.t1 327.466
R956 VTAIL.n219 VTAIL.t0 327.466
R957 VTAIL.n21 VTAIL.t3 327.466
R958 VTAIL.n222 VTAIL.n221 171.744
R959 VTAIL.n222 VTAIL.n215 171.744
R960 VTAIL.n229 VTAIL.n215 171.744
R961 VTAIL.n230 VTAIL.n229 171.744
R962 VTAIL.n230 VTAIL.n211 171.744
R963 VTAIL.n237 VTAIL.n211 171.744
R964 VTAIL.n238 VTAIL.n237 171.744
R965 VTAIL.n238 VTAIL.n207 171.744
R966 VTAIL.n245 VTAIL.n207 171.744
R967 VTAIL.n246 VTAIL.n245 171.744
R968 VTAIL.n246 VTAIL.n203 171.744
R969 VTAIL.n253 VTAIL.n203 171.744
R970 VTAIL.n254 VTAIL.n253 171.744
R971 VTAIL.n254 VTAIL.n199 171.744
R972 VTAIL.n261 VTAIL.n199 171.744
R973 VTAIL.n24 VTAIL.n23 171.744
R974 VTAIL.n24 VTAIL.n17 171.744
R975 VTAIL.n31 VTAIL.n17 171.744
R976 VTAIL.n32 VTAIL.n31 171.744
R977 VTAIL.n32 VTAIL.n13 171.744
R978 VTAIL.n39 VTAIL.n13 171.744
R979 VTAIL.n40 VTAIL.n39 171.744
R980 VTAIL.n40 VTAIL.n9 171.744
R981 VTAIL.n47 VTAIL.n9 171.744
R982 VTAIL.n48 VTAIL.n47 171.744
R983 VTAIL.n48 VTAIL.n5 171.744
R984 VTAIL.n55 VTAIL.n5 171.744
R985 VTAIL.n56 VTAIL.n55 171.744
R986 VTAIL.n56 VTAIL.n1 171.744
R987 VTAIL.n63 VTAIL.n1 171.744
R988 VTAIL.n195 VTAIL.n133 171.744
R989 VTAIL.n188 VTAIL.n133 171.744
R990 VTAIL.n188 VTAIL.n187 171.744
R991 VTAIL.n187 VTAIL.n137 171.744
R992 VTAIL.n180 VTAIL.n137 171.744
R993 VTAIL.n180 VTAIL.n179 171.744
R994 VTAIL.n179 VTAIL.n141 171.744
R995 VTAIL.n172 VTAIL.n141 171.744
R996 VTAIL.n172 VTAIL.n171 171.744
R997 VTAIL.n171 VTAIL.n145 171.744
R998 VTAIL.n164 VTAIL.n145 171.744
R999 VTAIL.n164 VTAIL.n163 171.744
R1000 VTAIL.n163 VTAIL.n149 171.744
R1001 VTAIL.n156 VTAIL.n149 171.744
R1002 VTAIL.n156 VTAIL.n155 171.744
R1003 VTAIL.n129 VTAIL.n67 171.744
R1004 VTAIL.n122 VTAIL.n67 171.744
R1005 VTAIL.n122 VTAIL.n121 171.744
R1006 VTAIL.n121 VTAIL.n71 171.744
R1007 VTAIL.n114 VTAIL.n71 171.744
R1008 VTAIL.n114 VTAIL.n113 171.744
R1009 VTAIL.n113 VTAIL.n75 171.744
R1010 VTAIL.n106 VTAIL.n75 171.744
R1011 VTAIL.n106 VTAIL.n105 171.744
R1012 VTAIL.n105 VTAIL.n79 171.744
R1013 VTAIL.n98 VTAIL.n79 171.744
R1014 VTAIL.n98 VTAIL.n97 171.744
R1015 VTAIL.n97 VTAIL.n83 171.744
R1016 VTAIL.n90 VTAIL.n83 171.744
R1017 VTAIL.n90 VTAIL.n89 171.744
R1018 VTAIL.n221 VTAIL.t0 85.8723
R1019 VTAIL.n23 VTAIL.t3 85.8723
R1020 VTAIL.n155 VTAIL.t2 85.8723
R1021 VTAIL.n89 VTAIL.t1 85.8723
R1022 VTAIL.n263 VTAIL.n262 34.5126
R1023 VTAIL.n65 VTAIL.n64 34.5126
R1024 VTAIL.n197 VTAIL.n196 34.5126
R1025 VTAIL.n131 VTAIL.n130 34.5126
R1026 VTAIL.n131 VTAIL.n65 27.591
R1027 VTAIL.n263 VTAIL.n197 25.1255
R1028 VTAIL.n220 VTAIL.n219 16.3895
R1029 VTAIL.n22 VTAIL.n21 16.3895
R1030 VTAIL.n154 VTAIL.n153 16.3895
R1031 VTAIL.n88 VTAIL.n87 16.3895
R1032 VTAIL.n223 VTAIL.n218 12.8005
R1033 VTAIL.n25 VTAIL.n20 12.8005
R1034 VTAIL.n157 VTAIL.n152 12.8005
R1035 VTAIL.n91 VTAIL.n86 12.8005
R1036 VTAIL.n224 VTAIL.n216 12.0247
R1037 VTAIL.n260 VTAIL.n198 12.0247
R1038 VTAIL.n26 VTAIL.n18 12.0247
R1039 VTAIL.n62 VTAIL.n0 12.0247
R1040 VTAIL.n194 VTAIL.n132 12.0247
R1041 VTAIL.n158 VTAIL.n150 12.0247
R1042 VTAIL.n128 VTAIL.n66 12.0247
R1043 VTAIL.n92 VTAIL.n84 12.0247
R1044 VTAIL.n228 VTAIL.n227 11.249
R1045 VTAIL.n259 VTAIL.n200 11.249
R1046 VTAIL.n30 VTAIL.n29 11.249
R1047 VTAIL.n61 VTAIL.n2 11.249
R1048 VTAIL.n193 VTAIL.n134 11.249
R1049 VTAIL.n162 VTAIL.n161 11.249
R1050 VTAIL.n127 VTAIL.n68 11.249
R1051 VTAIL.n96 VTAIL.n95 11.249
R1052 VTAIL.n231 VTAIL.n214 10.4732
R1053 VTAIL.n256 VTAIL.n255 10.4732
R1054 VTAIL.n33 VTAIL.n16 10.4732
R1055 VTAIL.n58 VTAIL.n57 10.4732
R1056 VTAIL.n190 VTAIL.n189 10.4732
R1057 VTAIL.n165 VTAIL.n148 10.4732
R1058 VTAIL.n124 VTAIL.n123 10.4732
R1059 VTAIL.n99 VTAIL.n82 10.4732
R1060 VTAIL.n232 VTAIL.n212 9.69747
R1061 VTAIL.n252 VTAIL.n202 9.69747
R1062 VTAIL.n34 VTAIL.n14 9.69747
R1063 VTAIL.n54 VTAIL.n4 9.69747
R1064 VTAIL.n186 VTAIL.n136 9.69747
R1065 VTAIL.n166 VTAIL.n146 9.69747
R1066 VTAIL.n120 VTAIL.n70 9.69747
R1067 VTAIL.n100 VTAIL.n80 9.69747
R1068 VTAIL.n258 VTAIL.n198 9.45567
R1069 VTAIL.n60 VTAIL.n0 9.45567
R1070 VTAIL.n192 VTAIL.n132 9.45567
R1071 VTAIL.n126 VTAIL.n66 9.45567
R1072 VTAIL.n243 VTAIL.n242 9.3005
R1073 VTAIL.n206 VTAIL.n205 9.3005
R1074 VTAIL.n249 VTAIL.n248 9.3005
R1075 VTAIL.n251 VTAIL.n250 9.3005
R1076 VTAIL.n202 VTAIL.n201 9.3005
R1077 VTAIL.n257 VTAIL.n256 9.3005
R1078 VTAIL.n259 VTAIL.n258 9.3005
R1079 VTAIL.n210 VTAIL.n209 9.3005
R1080 VTAIL.n235 VTAIL.n234 9.3005
R1081 VTAIL.n233 VTAIL.n232 9.3005
R1082 VTAIL.n214 VTAIL.n213 9.3005
R1083 VTAIL.n227 VTAIL.n226 9.3005
R1084 VTAIL.n225 VTAIL.n224 9.3005
R1085 VTAIL.n218 VTAIL.n217 9.3005
R1086 VTAIL.n241 VTAIL.n240 9.3005
R1087 VTAIL.n45 VTAIL.n44 9.3005
R1088 VTAIL.n8 VTAIL.n7 9.3005
R1089 VTAIL.n51 VTAIL.n50 9.3005
R1090 VTAIL.n53 VTAIL.n52 9.3005
R1091 VTAIL.n4 VTAIL.n3 9.3005
R1092 VTAIL.n59 VTAIL.n58 9.3005
R1093 VTAIL.n61 VTAIL.n60 9.3005
R1094 VTAIL.n12 VTAIL.n11 9.3005
R1095 VTAIL.n37 VTAIL.n36 9.3005
R1096 VTAIL.n35 VTAIL.n34 9.3005
R1097 VTAIL.n16 VTAIL.n15 9.3005
R1098 VTAIL.n29 VTAIL.n28 9.3005
R1099 VTAIL.n27 VTAIL.n26 9.3005
R1100 VTAIL.n20 VTAIL.n19 9.3005
R1101 VTAIL.n43 VTAIL.n42 9.3005
R1102 VTAIL.n193 VTAIL.n192 9.3005
R1103 VTAIL.n191 VTAIL.n190 9.3005
R1104 VTAIL.n136 VTAIL.n135 9.3005
R1105 VTAIL.n185 VTAIL.n184 9.3005
R1106 VTAIL.n183 VTAIL.n182 9.3005
R1107 VTAIL.n140 VTAIL.n139 9.3005
R1108 VTAIL.n177 VTAIL.n176 9.3005
R1109 VTAIL.n175 VTAIL.n174 9.3005
R1110 VTAIL.n144 VTAIL.n143 9.3005
R1111 VTAIL.n169 VTAIL.n168 9.3005
R1112 VTAIL.n167 VTAIL.n166 9.3005
R1113 VTAIL.n148 VTAIL.n147 9.3005
R1114 VTAIL.n161 VTAIL.n160 9.3005
R1115 VTAIL.n159 VTAIL.n158 9.3005
R1116 VTAIL.n152 VTAIL.n151 9.3005
R1117 VTAIL.n74 VTAIL.n73 9.3005
R1118 VTAIL.n117 VTAIL.n116 9.3005
R1119 VTAIL.n119 VTAIL.n118 9.3005
R1120 VTAIL.n70 VTAIL.n69 9.3005
R1121 VTAIL.n125 VTAIL.n124 9.3005
R1122 VTAIL.n127 VTAIL.n126 9.3005
R1123 VTAIL.n111 VTAIL.n110 9.3005
R1124 VTAIL.n109 VTAIL.n108 9.3005
R1125 VTAIL.n78 VTAIL.n77 9.3005
R1126 VTAIL.n103 VTAIL.n102 9.3005
R1127 VTAIL.n101 VTAIL.n100 9.3005
R1128 VTAIL.n82 VTAIL.n81 9.3005
R1129 VTAIL.n95 VTAIL.n94 9.3005
R1130 VTAIL.n93 VTAIL.n92 9.3005
R1131 VTAIL.n86 VTAIL.n85 9.3005
R1132 VTAIL.n236 VTAIL.n235 8.92171
R1133 VTAIL.n251 VTAIL.n204 8.92171
R1134 VTAIL.n38 VTAIL.n37 8.92171
R1135 VTAIL.n53 VTAIL.n6 8.92171
R1136 VTAIL.n185 VTAIL.n138 8.92171
R1137 VTAIL.n170 VTAIL.n169 8.92171
R1138 VTAIL.n119 VTAIL.n72 8.92171
R1139 VTAIL.n104 VTAIL.n103 8.92171
R1140 VTAIL.n239 VTAIL.n210 8.14595
R1141 VTAIL.n248 VTAIL.n247 8.14595
R1142 VTAIL.n41 VTAIL.n12 8.14595
R1143 VTAIL.n50 VTAIL.n49 8.14595
R1144 VTAIL.n182 VTAIL.n181 8.14595
R1145 VTAIL.n173 VTAIL.n144 8.14595
R1146 VTAIL.n116 VTAIL.n115 8.14595
R1147 VTAIL.n107 VTAIL.n78 8.14595
R1148 VTAIL.n240 VTAIL.n208 7.3702
R1149 VTAIL.n244 VTAIL.n206 7.3702
R1150 VTAIL.n42 VTAIL.n10 7.3702
R1151 VTAIL.n46 VTAIL.n8 7.3702
R1152 VTAIL.n178 VTAIL.n140 7.3702
R1153 VTAIL.n174 VTAIL.n142 7.3702
R1154 VTAIL.n112 VTAIL.n74 7.3702
R1155 VTAIL.n108 VTAIL.n76 7.3702
R1156 VTAIL.n243 VTAIL.n208 6.59444
R1157 VTAIL.n244 VTAIL.n243 6.59444
R1158 VTAIL.n45 VTAIL.n10 6.59444
R1159 VTAIL.n46 VTAIL.n45 6.59444
R1160 VTAIL.n178 VTAIL.n177 6.59444
R1161 VTAIL.n177 VTAIL.n142 6.59444
R1162 VTAIL.n112 VTAIL.n111 6.59444
R1163 VTAIL.n111 VTAIL.n76 6.59444
R1164 VTAIL.n240 VTAIL.n239 5.81868
R1165 VTAIL.n247 VTAIL.n206 5.81868
R1166 VTAIL.n42 VTAIL.n41 5.81868
R1167 VTAIL.n49 VTAIL.n8 5.81868
R1168 VTAIL.n181 VTAIL.n140 5.81868
R1169 VTAIL.n174 VTAIL.n173 5.81868
R1170 VTAIL.n115 VTAIL.n74 5.81868
R1171 VTAIL.n108 VTAIL.n107 5.81868
R1172 VTAIL.n236 VTAIL.n210 5.04292
R1173 VTAIL.n248 VTAIL.n204 5.04292
R1174 VTAIL.n38 VTAIL.n12 5.04292
R1175 VTAIL.n50 VTAIL.n6 5.04292
R1176 VTAIL.n182 VTAIL.n138 5.04292
R1177 VTAIL.n170 VTAIL.n144 5.04292
R1178 VTAIL.n116 VTAIL.n72 5.04292
R1179 VTAIL.n104 VTAIL.n78 5.04292
R1180 VTAIL.n235 VTAIL.n212 4.26717
R1181 VTAIL.n252 VTAIL.n251 4.26717
R1182 VTAIL.n37 VTAIL.n14 4.26717
R1183 VTAIL.n54 VTAIL.n53 4.26717
R1184 VTAIL.n186 VTAIL.n185 4.26717
R1185 VTAIL.n169 VTAIL.n146 4.26717
R1186 VTAIL.n120 VTAIL.n119 4.26717
R1187 VTAIL.n103 VTAIL.n80 4.26717
R1188 VTAIL.n153 VTAIL.n151 3.70982
R1189 VTAIL.n87 VTAIL.n85 3.70982
R1190 VTAIL.n219 VTAIL.n217 3.70982
R1191 VTAIL.n21 VTAIL.n19 3.70982
R1192 VTAIL.n232 VTAIL.n231 3.49141
R1193 VTAIL.n255 VTAIL.n202 3.49141
R1194 VTAIL.n34 VTAIL.n33 3.49141
R1195 VTAIL.n57 VTAIL.n4 3.49141
R1196 VTAIL.n189 VTAIL.n136 3.49141
R1197 VTAIL.n166 VTAIL.n165 3.49141
R1198 VTAIL.n123 VTAIL.n70 3.49141
R1199 VTAIL.n100 VTAIL.n99 3.49141
R1200 VTAIL.n228 VTAIL.n214 2.71565
R1201 VTAIL.n256 VTAIL.n200 2.71565
R1202 VTAIL.n30 VTAIL.n16 2.71565
R1203 VTAIL.n58 VTAIL.n2 2.71565
R1204 VTAIL.n190 VTAIL.n134 2.71565
R1205 VTAIL.n162 VTAIL.n148 2.71565
R1206 VTAIL.n124 VTAIL.n68 2.71565
R1207 VTAIL.n96 VTAIL.n82 2.71565
R1208 VTAIL.n227 VTAIL.n216 1.93989
R1209 VTAIL.n260 VTAIL.n259 1.93989
R1210 VTAIL.n29 VTAIL.n18 1.93989
R1211 VTAIL.n62 VTAIL.n61 1.93989
R1212 VTAIL.n194 VTAIL.n193 1.93989
R1213 VTAIL.n161 VTAIL.n150 1.93989
R1214 VTAIL.n128 VTAIL.n127 1.93989
R1215 VTAIL.n95 VTAIL.n84 1.93989
R1216 VTAIL.n197 VTAIL.n131 1.70309
R1217 VTAIL.n224 VTAIL.n223 1.16414
R1218 VTAIL.n262 VTAIL.n198 1.16414
R1219 VTAIL.n26 VTAIL.n25 1.16414
R1220 VTAIL.n64 VTAIL.n0 1.16414
R1221 VTAIL.n196 VTAIL.n132 1.16414
R1222 VTAIL.n158 VTAIL.n157 1.16414
R1223 VTAIL.n130 VTAIL.n66 1.16414
R1224 VTAIL.n92 VTAIL.n91 1.16414
R1225 VTAIL VTAIL.n65 1.1449
R1226 VTAIL VTAIL.n263 0.55869
R1227 VTAIL.n220 VTAIL.n218 0.388379
R1228 VTAIL.n22 VTAIL.n20 0.388379
R1229 VTAIL.n154 VTAIL.n152 0.388379
R1230 VTAIL.n88 VTAIL.n86 0.388379
R1231 VTAIL.n225 VTAIL.n217 0.155672
R1232 VTAIL.n226 VTAIL.n225 0.155672
R1233 VTAIL.n226 VTAIL.n213 0.155672
R1234 VTAIL.n233 VTAIL.n213 0.155672
R1235 VTAIL.n234 VTAIL.n233 0.155672
R1236 VTAIL.n234 VTAIL.n209 0.155672
R1237 VTAIL.n241 VTAIL.n209 0.155672
R1238 VTAIL.n242 VTAIL.n241 0.155672
R1239 VTAIL.n242 VTAIL.n205 0.155672
R1240 VTAIL.n249 VTAIL.n205 0.155672
R1241 VTAIL.n250 VTAIL.n249 0.155672
R1242 VTAIL.n250 VTAIL.n201 0.155672
R1243 VTAIL.n257 VTAIL.n201 0.155672
R1244 VTAIL.n258 VTAIL.n257 0.155672
R1245 VTAIL.n27 VTAIL.n19 0.155672
R1246 VTAIL.n28 VTAIL.n27 0.155672
R1247 VTAIL.n28 VTAIL.n15 0.155672
R1248 VTAIL.n35 VTAIL.n15 0.155672
R1249 VTAIL.n36 VTAIL.n35 0.155672
R1250 VTAIL.n36 VTAIL.n11 0.155672
R1251 VTAIL.n43 VTAIL.n11 0.155672
R1252 VTAIL.n44 VTAIL.n43 0.155672
R1253 VTAIL.n44 VTAIL.n7 0.155672
R1254 VTAIL.n51 VTAIL.n7 0.155672
R1255 VTAIL.n52 VTAIL.n51 0.155672
R1256 VTAIL.n52 VTAIL.n3 0.155672
R1257 VTAIL.n59 VTAIL.n3 0.155672
R1258 VTAIL.n60 VTAIL.n59 0.155672
R1259 VTAIL.n192 VTAIL.n191 0.155672
R1260 VTAIL.n191 VTAIL.n135 0.155672
R1261 VTAIL.n184 VTAIL.n135 0.155672
R1262 VTAIL.n184 VTAIL.n183 0.155672
R1263 VTAIL.n183 VTAIL.n139 0.155672
R1264 VTAIL.n176 VTAIL.n139 0.155672
R1265 VTAIL.n176 VTAIL.n175 0.155672
R1266 VTAIL.n175 VTAIL.n143 0.155672
R1267 VTAIL.n168 VTAIL.n143 0.155672
R1268 VTAIL.n168 VTAIL.n167 0.155672
R1269 VTAIL.n167 VTAIL.n147 0.155672
R1270 VTAIL.n160 VTAIL.n147 0.155672
R1271 VTAIL.n160 VTAIL.n159 0.155672
R1272 VTAIL.n159 VTAIL.n151 0.155672
R1273 VTAIL.n126 VTAIL.n125 0.155672
R1274 VTAIL.n125 VTAIL.n69 0.155672
R1275 VTAIL.n118 VTAIL.n69 0.155672
R1276 VTAIL.n118 VTAIL.n117 0.155672
R1277 VTAIL.n117 VTAIL.n73 0.155672
R1278 VTAIL.n110 VTAIL.n73 0.155672
R1279 VTAIL.n110 VTAIL.n109 0.155672
R1280 VTAIL.n109 VTAIL.n77 0.155672
R1281 VTAIL.n102 VTAIL.n77 0.155672
R1282 VTAIL.n102 VTAIL.n101 0.155672
R1283 VTAIL.n101 VTAIL.n81 0.155672
R1284 VTAIL.n94 VTAIL.n81 0.155672
R1285 VTAIL.n94 VTAIL.n93 0.155672
R1286 VTAIL.n93 VTAIL.n85 0.155672
R1287 VDD1.n64 VDD1.n63 756.745
R1288 VDD1.n129 VDD1.n128 756.745
R1289 VDD1.n63 VDD1.n62 585
R1290 VDD1.n2 VDD1.n1 585
R1291 VDD1.n57 VDD1.n56 585
R1292 VDD1.n55 VDD1.n54 585
R1293 VDD1.n6 VDD1.n5 585
R1294 VDD1.n49 VDD1.n48 585
R1295 VDD1.n47 VDD1.n46 585
R1296 VDD1.n10 VDD1.n9 585
R1297 VDD1.n41 VDD1.n40 585
R1298 VDD1.n39 VDD1.n38 585
R1299 VDD1.n14 VDD1.n13 585
R1300 VDD1.n33 VDD1.n32 585
R1301 VDD1.n31 VDD1.n30 585
R1302 VDD1.n18 VDD1.n17 585
R1303 VDD1.n25 VDD1.n24 585
R1304 VDD1.n23 VDD1.n22 585
R1305 VDD1.n88 VDD1.n87 585
R1306 VDD1.n90 VDD1.n89 585
R1307 VDD1.n83 VDD1.n82 585
R1308 VDD1.n96 VDD1.n95 585
R1309 VDD1.n98 VDD1.n97 585
R1310 VDD1.n79 VDD1.n78 585
R1311 VDD1.n104 VDD1.n103 585
R1312 VDD1.n106 VDD1.n105 585
R1313 VDD1.n75 VDD1.n74 585
R1314 VDD1.n112 VDD1.n111 585
R1315 VDD1.n114 VDD1.n113 585
R1316 VDD1.n71 VDD1.n70 585
R1317 VDD1.n120 VDD1.n119 585
R1318 VDD1.n122 VDD1.n121 585
R1319 VDD1.n67 VDD1.n66 585
R1320 VDD1.n128 VDD1.n127 585
R1321 VDD1.n21 VDD1.t0 327.466
R1322 VDD1.n86 VDD1.t1 327.466
R1323 VDD1.n63 VDD1.n1 171.744
R1324 VDD1.n56 VDD1.n1 171.744
R1325 VDD1.n56 VDD1.n55 171.744
R1326 VDD1.n55 VDD1.n5 171.744
R1327 VDD1.n48 VDD1.n5 171.744
R1328 VDD1.n48 VDD1.n47 171.744
R1329 VDD1.n47 VDD1.n9 171.744
R1330 VDD1.n40 VDD1.n9 171.744
R1331 VDD1.n40 VDD1.n39 171.744
R1332 VDD1.n39 VDD1.n13 171.744
R1333 VDD1.n32 VDD1.n13 171.744
R1334 VDD1.n32 VDD1.n31 171.744
R1335 VDD1.n31 VDD1.n17 171.744
R1336 VDD1.n24 VDD1.n17 171.744
R1337 VDD1.n24 VDD1.n23 171.744
R1338 VDD1.n89 VDD1.n88 171.744
R1339 VDD1.n89 VDD1.n82 171.744
R1340 VDD1.n96 VDD1.n82 171.744
R1341 VDD1.n97 VDD1.n96 171.744
R1342 VDD1.n97 VDD1.n78 171.744
R1343 VDD1.n104 VDD1.n78 171.744
R1344 VDD1.n105 VDD1.n104 171.744
R1345 VDD1.n105 VDD1.n74 171.744
R1346 VDD1.n112 VDD1.n74 171.744
R1347 VDD1.n113 VDD1.n112 171.744
R1348 VDD1.n113 VDD1.n70 171.744
R1349 VDD1.n120 VDD1.n70 171.744
R1350 VDD1.n121 VDD1.n120 171.744
R1351 VDD1.n121 VDD1.n66 171.744
R1352 VDD1.n128 VDD1.n66 171.744
R1353 VDD1 VDD1.n129 91.2162
R1354 VDD1.n23 VDD1.t0 85.8723
R1355 VDD1.n88 VDD1.t1 85.8723
R1356 VDD1 VDD1.n64 51.866
R1357 VDD1.n22 VDD1.n21 16.3895
R1358 VDD1.n87 VDD1.n86 16.3895
R1359 VDD1.n25 VDD1.n20 12.8005
R1360 VDD1.n90 VDD1.n85 12.8005
R1361 VDD1.n62 VDD1.n0 12.0247
R1362 VDD1.n26 VDD1.n18 12.0247
R1363 VDD1.n91 VDD1.n83 12.0247
R1364 VDD1.n127 VDD1.n65 12.0247
R1365 VDD1.n61 VDD1.n2 11.249
R1366 VDD1.n30 VDD1.n29 11.249
R1367 VDD1.n95 VDD1.n94 11.249
R1368 VDD1.n126 VDD1.n67 11.249
R1369 VDD1.n58 VDD1.n57 10.4732
R1370 VDD1.n33 VDD1.n16 10.4732
R1371 VDD1.n98 VDD1.n81 10.4732
R1372 VDD1.n123 VDD1.n122 10.4732
R1373 VDD1.n54 VDD1.n4 9.69747
R1374 VDD1.n34 VDD1.n14 9.69747
R1375 VDD1.n99 VDD1.n79 9.69747
R1376 VDD1.n119 VDD1.n69 9.69747
R1377 VDD1.n60 VDD1.n0 9.45567
R1378 VDD1.n125 VDD1.n65 9.45567
R1379 VDD1.n61 VDD1.n60 9.3005
R1380 VDD1.n59 VDD1.n58 9.3005
R1381 VDD1.n4 VDD1.n3 9.3005
R1382 VDD1.n53 VDD1.n52 9.3005
R1383 VDD1.n51 VDD1.n50 9.3005
R1384 VDD1.n8 VDD1.n7 9.3005
R1385 VDD1.n45 VDD1.n44 9.3005
R1386 VDD1.n43 VDD1.n42 9.3005
R1387 VDD1.n12 VDD1.n11 9.3005
R1388 VDD1.n37 VDD1.n36 9.3005
R1389 VDD1.n35 VDD1.n34 9.3005
R1390 VDD1.n16 VDD1.n15 9.3005
R1391 VDD1.n29 VDD1.n28 9.3005
R1392 VDD1.n27 VDD1.n26 9.3005
R1393 VDD1.n20 VDD1.n19 9.3005
R1394 VDD1.n110 VDD1.n109 9.3005
R1395 VDD1.n73 VDD1.n72 9.3005
R1396 VDD1.n116 VDD1.n115 9.3005
R1397 VDD1.n118 VDD1.n117 9.3005
R1398 VDD1.n69 VDD1.n68 9.3005
R1399 VDD1.n124 VDD1.n123 9.3005
R1400 VDD1.n126 VDD1.n125 9.3005
R1401 VDD1.n77 VDD1.n76 9.3005
R1402 VDD1.n102 VDD1.n101 9.3005
R1403 VDD1.n100 VDD1.n99 9.3005
R1404 VDD1.n81 VDD1.n80 9.3005
R1405 VDD1.n94 VDD1.n93 9.3005
R1406 VDD1.n92 VDD1.n91 9.3005
R1407 VDD1.n85 VDD1.n84 9.3005
R1408 VDD1.n108 VDD1.n107 9.3005
R1409 VDD1.n53 VDD1.n6 8.92171
R1410 VDD1.n38 VDD1.n37 8.92171
R1411 VDD1.n103 VDD1.n102 8.92171
R1412 VDD1.n118 VDD1.n71 8.92171
R1413 VDD1.n50 VDD1.n49 8.14595
R1414 VDD1.n41 VDD1.n12 8.14595
R1415 VDD1.n106 VDD1.n77 8.14595
R1416 VDD1.n115 VDD1.n114 8.14595
R1417 VDD1.n46 VDD1.n8 7.3702
R1418 VDD1.n42 VDD1.n10 7.3702
R1419 VDD1.n107 VDD1.n75 7.3702
R1420 VDD1.n111 VDD1.n73 7.3702
R1421 VDD1.n46 VDD1.n45 6.59444
R1422 VDD1.n45 VDD1.n10 6.59444
R1423 VDD1.n110 VDD1.n75 6.59444
R1424 VDD1.n111 VDD1.n110 6.59444
R1425 VDD1.n49 VDD1.n8 5.81868
R1426 VDD1.n42 VDD1.n41 5.81868
R1427 VDD1.n107 VDD1.n106 5.81868
R1428 VDD1.n114 VDD1.n73 5.81868
R1429 VDD1.n50 VDD1.n6 5.04292
R1430 VDD1.n38 VDD1.n12 5.04292
R1431 VDD1.n103 VDD1.n77 5.04292
R1432 VDD1.n115 VDD1.n71 5.04292
R1433 VDD1.n54 VDD1.n53 4.26717
R1434 VDD1.n37 VDD1.n14 4.26717
R1435 VDD1.n102 VDD1.n79 4.26717
R1436 VDD1.n119 VDD1.n118 4.26717
R1437 VDD1.n21 VDD1.n19 3.70982
R1438 VDD1.n86 VDD1.n84 3.70982
R1439 VDD1.n57 VDD1.n4 3.49141
R1440 VDD1.n34 VDD1.n33 3.49141
R1441 VDD1.n99 VDD1.n98 3.49141
R1442 VDD1.n122 VDD1.n69 3.49141
R1443 VDD1.n58 VDD1.n2 2.71565
R1444 VDD1.n30 VDD1.n16 2.71565
R1445 VDD1.n95 VDD1.n81 2.71565
R1446 VDD1.n123 VDD1.n67 2.71565
R1447 VDD1.n62 VDD1.n61 1.93989
R1448 VDD1.n29 VDD1.n18 1.93989
R1449 VDD1.n94 VDD1.n83 1.93989
R1450 VDD1.n127 VDD1.n126 1.93989
R1451 VDD1.n64 VDD1.n0 1.16414
R1452 VDD1.n26 VDD1.n25 1.16414
R1453 VDD1.n91 VDD1.n90 1.16414
R1454 VDD1.n129 VDD1.n65 1.16414
R1455 VDD1.n22 VDD1.n20 0.388379
R1456 VDD1.n87 VDD1.n85 0.388379
R1457 VDD1.n60 VDD1.n59 0.155672
R1458 VDD1.n59 VDD1.n3 0.155672
R1459 VDD1.n52 VDD1.n3 0.155672
R1460 VDD1.n52 VDD1.n51 0.155672
R1461 VDD1.n51 VDD1.n7 0.155672
R1462 VDD1.n44 VDD1.n7 0.155672
R1463 VDD1.n44 VDD1.n43 0.155672
R1464 VDD1.n43 VDD1.n11 0.155672
R1465 VDD1.n36 VDD1.n11 0.155672
R1466 VDD1.n36 VDD1.n35 0.155672
R1467 VDD1.n35 VDD1.n15 0.155672
R1468 VDD1.n28 VDD1.n15 0.155672
R1469 VDD1.n28 VDD1.n27 0.155672
R1470 VDD1.n27 VDD1.n19 0.155672
R1471 VDD1.n92 VDD1.n84 0.155672
R1472 VDD1.n93 VDD1.n92 0.155672
R1473 VDD1.n93 VDD1.n80 0.155672
R1474 VDD1.n100 VDD1.n80 0.155672
R1475 VDD1.n101 VDD1.n100 0.155672
R1476 VDD1.n101 VDD1.n76 0.155672
R1477 VDD1.n108 VDD1.n76 0.155672
R1478 VDD1.n109 VDD1.n108 0.155672
R1479 VDD1.n109 VDD1.n72 0.155672
R1480 VDD1.n116 VDD1.n72 0.155672
R1481 VDD1.n117 VDD1.n116 0.155672
R1482 VDD1.n117 VDD1.n68 0.155672
R1483 VDD1.n124 VDD1.n68 0.155672
R1484 VDD1.n125 VDD1.n124 0.155672
R1485 VN VN.t1 207.475
R1486 VN VN.t0 163.288
R1487 VDD2.n129 VDD2.n128 756.745
R1488 VDD2.n64 VDD2.n63 756.745
R1489 VDD2.n128 VDD2.n127 585
R1490 VDD2.n67 VDD2.n66 585
R1491 VDD2.n122 VDD2.n121 585
R1492 VDD2.n120 VDD2.n119 585
R1493 VDD2.n71 VDD2.n70 585
R1494 VDD2.n114 VDD2.n113 585
R1495 VDD2.n112 VDD2.n111 585
R1496 VDD2.n75 VDD2.n74 585
R1497 VDD2.n106 VDD2.n105 585
R1498 VDD2.n104 VDD2.n103 585
R1499 VDD2.n79 VDD2.n78 585
R1500 VDD2.n98 VDD2.n97 585
R1501 VDD2.n96 VDD2.n95 585
R1502 VDD2.n83 VDD2.n82 585
R1503 VDD2.n90 VDD2.n89 585
R1504 VDD2.n88 VDD2.n87 585
R1505 VDD2.n23 VDD2.n22 585
R1506 VDD2.n25 VDD2.n24 585
R1507 VDD2.n18 VDD2.n17 585
R1508 VDD2.n31 VDD2.n30 585
R1509 VDD2.n33 VDD2.n32 585
R1510 VDD2.n14 VDD2.n13 585
R1511 VDD2.n39 VDD2.n38 585
R1512 VDD2.n41 VDD2.n40 585
R1513 VDD2.n10 VDD2.n9 585
R1514 VDD2.n47 VDD2.n46 585
R1515 VDD2.n49 VDD2.n48 585
R1516 VDD2.n6 VDD2.n5 585
R1517 VDD2.n55 VDD2.n54 585
R1518 VDD2.n57 VDD2.n56 585
R1519 VDD2.n2 VDD2.n1 585
R1520 VDD2.n63 VDD2.n62 585
R1521 VDD2.n86 VDD2.t0 327.466
R1522 VDD2.n21 VDD2.t1 327.466
R1523 VDD2.n128 VDD2.n66 171.744
R1524 VDD2.n121 VDD2.n66 171.744
R1525 VDD2.n121 VDD2.n120 171.744
R1526 VDD2.n120 VDD2.n70 171.744
R1527 VDD2.n113 VDD2.n70 171.744
R1528 VDD2.n113 VDD2.n112 171.744
R1529 VDD2.n112 VDD2.n74 171.744
R1530 VDD2.n105 VDD2.n74 171.744
R1531 VDD2.n105 VDD2.n104 171.744
R1532 VDD2.n104 VDD2.n78 171.744
R1533 VDD2.n97 VDD2.n78 171.744
R1534 VDD2.n97 VDD2.n96 171.744
R1535 VDD2.n96 VDD2.n82 171.744
R1536 VDD2.n89 VDD2.n82 171.744
R1537 VDD2.n89 VDD2.n88 171.744
R1538 VDD2.n24 VDD2.n23 171.744
R1539 VDD2.n24 VDD2.n17 171.744
R1540 VDD2.n31 VDD2.n17 171.744
R1541 VDD2.n32 VDD2.n31 171.744
R1542 VDD2.n32 VDD2.n13 171.744
R1543 VDD2.n39 VDD2.n13 171.744
R1544 VDD2.n40 VDD2.n39 171.744
R1545 VDD2.n40 VDD2.n9 171.744
R1546 VDD2.n47 VDD2.n9 171.744
R1547 VDD2.n48 VDD2.n47 171.744
R1548 VDD2.n48 VDD2.n5 171.744
R1549 VDD2.n55 VDD2.n5 171.744
R1550 VDD2.n56 VDD2.n55 171.744
R1551 VDD2.n56 VDD2.n1 171.744
R1552 VDD2.n63 VDD2.n1 171.744
R1553 VDD2.n130 VDD2.n64 90.075
R1554 VDD2.n88 VDD2.t0 85.8723
R1555 VDD2.n23 VDD2.t1 85.8723
R1556 VDD2.n130 VDD2.n129 51.1914
R1557 VDD2.n87 VDD2.n86 16.3895
R1558 VDD2.n22 VDD2.n21 16.3895
R1559 VDD2.n90 VDD2.n85 12.8005
R1560 VDD2.n25 VDD2.n20 12.8005
R1561 VDD2.n127 VDD2.n65 12.0247
R1562 VDD2.n91 VDD2.n83 12.0247
R1563 VDD2.n26 VDD2.n18 12.0247
R1564 VDD2.n62 VDD2.n0 12.0247
R1565 VDD2.n126 VDD2.n67 11.249
R1566 VDD2.n95 VDD2.n94 11.249
R1567 VDD2.n30 VDD2.n29 11.249
R1568 VDD2.n61 VDD2.n2 11.249
R1569 VDD2.n123 VDD2.n122 10.4732
R1570 VDD2.n98 VDD2.n81 10.4732
R1571 VDD2.n33 VDD2.n16 10.4732
R1572 VDD2.n58 VDD2.n57 10.4732
R1573 VDD2.n119 VDD2.n69 9.69747
R1574 VDD2.n99 VDD2.n79 9.69747
R1575 VDD2.n34 VDD2.n14 9.69747
R1576 VDD2.n54 VDD2.n4 9.69747
R1577 VDD2.n125 VDD2.n65 9.45567
R1578 VDD2.n60 VDD2.n0 9.45567
R1579 VDD2.n126 VDD2.n125 9.3005
R1580 VDD2.n124 VDD2.n123 9.3005
R1581 VDD2.n69 VDD2.n68 9.3005
R1582 VDD2.n118 VDD2.n117 9.3005
R1583 VDD2.n116 VDD2.n115 9.3005
R1584 VDD2.n73 VDD2.n72 9.3005
R1585 VDD2.n110 VDD2.n109 9.3005
R1586 VDD2.n108 VDD2.n107 9.3005
R1587 VDD2.n77 VDD2.n76 9.3005
R1588 VDD2.n102 VDD2.n101 9.3005
R1589 VDD2.n100 VDD2.n99 9.3005
R1590 VDD2.n81 VDD2.n80 9.3005
R1591 VDD2.n94 VDD2.n93 9.3005
R1592 VDD2.n92 VDD2.n91 9.3005
R1593 VDD2.n85 VDD2.n84 9.3005
R1594 VDD2.n45 VDD2.n44 9.3005
R1595 VDD2.n8 VDD2.n7 9.3005
R1596 VDD2.n51 VDD2.n50 9.3005
R1597 VDD2.n53 VDD2.n52 9.3005
R1598 VDD2.n4 VDD2.n3 9.3005
R1599 VDD2.n59 VDD2.n58 9.3005
R1600 VDD2.n61 VDD2.n60 9.3005
R1601 VDD2.n12 VDD2.n11 9.3005
R1602 VDD2.n37 VDD2.n36 9.3005
R1603 VDD2.n35 VDD2.n34 9.3005
R1604 VDD2.n16 VDD2.n15 9.3005
R1605 VDD2.n29 VDD2.n28 9.3005
R1606 VDD2.n27 VDD2.n26 9.3005
R1607 VDD2.n20 VDD2.n19 9.3005
R1608 VDD2.n43 VDD2.n42 9.3005
R1609 VDD2.n118 VDD2.n71 8.92171
R1610 VDD2.n103 VDD2.n102 8.92171
R1611 VDD2.n38 VDD2.n37 8.92171
R1612 VDD2.n53 VDD2.n6 8.92171
R1613 VDD2.n115 VDD2.n114 8.14595
R1614 VDD2.n106 VDD2.n77 8.14595
R1615 VDD2.n41 VDD2.n12 8.14595
R1616 VDD2.n50 VDD2.n49 8.14595
R1617 VDD2.n111 VDD2.n73 7.3702
R1618 VDD2.n107 VDD2.n75 7.3702
R1619 VDD2.n42 VDD2.n10 7.3702
R1620 VDD2.n46 VDD2.n8 7.3702
R1621 VDD2.n111 VDD2.n110 6.59444
R1622 VDD2.n110 VDD2.n75 6.59444
R1623 VDD2.n45 VDD2.n10 6.59444
R1624 VDD2.n46 VDD2.n45 6.59444
R1625 VDD2.n114 VDD2.n73 5.81868
R1626 VDD2.n107 VDD2.n106 5.81868
R1627 VDD2.n42 VDD2.n41 5.81868
R1628 VDD2.n49 VDD2.n8 5.81868
R1629 VDD2.n115 VDD2.n71 5.04292
R1630 VDD2.n103 VDD2.n77 5.04292
R1631 VDD2.n38 VDD2.n12 5.04292
R1632 VDD2.n50 VDD2.n6 5.04292
R1633 VDD2.n119 VDD2.n118 4.26717
R1634 VDD2.n102 VDD2.n79 4.26717
R1635 VDD2.n37 VDD2.n14 4.26717
R1636 VDD2.n54 VDD2.n53 4.26717
R1637 VDD2.n86 VDD2.n84 3.70982
R1638 VDD2.n21 VDD2.n19 3.70982
R1639 VDD2.n122 VDD2.n69 3.49141
R1640 VDD2.n99 VDD2.n98 3.49141
R1641 VDD2.n34 VDD2.n33 3.49141
R1642 VDD2.n57 VDD2.n4 3.49141
R1643 VDD2.n123 VDD2.n67 2.71565
R1644 VDD2.n95 VDD2.n81 2.71565
R1645 VDD2.n30 VDD2.n16 2.71565
R1646 VDD2.n58 VDD2.n2 2.71565
R1647 VDD2.n127 VDD2.n126 1.93989
R1648 VDD2.n94 VDD2.n83 1.93989
R1649 VDD2.n29 VDD2.n18 1.93989
R1650 VDD2.n62 VDD2.n61 1.93989
R1651 VDD2.n129 VDD2.n65 1.16414
R1652 VDD2.n91 VDD2.n90 1.16414
R1653 VDD2.n26 VDD2.n25 1.16414
R1654 VDD2.n64 VDD2.n0 1.16414
R1655 VDD2 VDD2.n130 0.675069
R1656 VDD2.n87 VDD2.n85 0.388379
R1657 VDD2.n22 VDD2.n20 0.388379
R1658 VDD2.n125 VDD2.n124 0.155672
R1659 VDD2.n124 VDD2.n68 0.155672
R1660 VDD2.n117 VDD2.n68 0.155672
R1661 VDD2.n117 VDD2.n116 0.155672
R1662 VDD2.n116 VDD2.n72 0.155672
R1663 VDD2.n109 VDD2.n72 0.155672
R1664 VDD2.n109 VDD2.n108 0.155672
R1665 VDD2.n108 VDD2.n76 0.155672
R1666 VDD2.n101 VDD2.n76 0.155672
R1667 VDD2.n101 VDD2.n100 0.155672
R1668 VDD2.n100 VDD2.n80 0.155672
R1669 VDD2.n93 VDD2.n80 0.155672
R1670 VDD2.n93 VDD2.n92 0.155672
R1671 VDD2.n92 VDD2.n84 0.155672
R1672 VDD2.n27 VDD2.n19 0.155672
R1673 VDD2.n28 VDD2.n27 0.155672
R1674 VDD2.n28 VDD2.n15 0.155672
R1675 VDD2.n35 VDD2.n15 0.155672
R1676 VDD2.n36 VDD2.n35 0.155672
R1677 VDD2.n36 VDD2.n11 0.155672
R1678 VDD2.n43 VDD2.n11 0.155672
R1679 VDD2.n44 VDD2.n43 0.155672
R1680 VDD2.n44 VDD2.n7 0.155672
R1681 VDD2.n51 VDD2.n7 0.155672
R1682 VDD2.n52 VDD2.n51 0.155672
R1683 VDD2.n52 VDD2.n3 0.155672
R1684 VDD2.n59 VDD2.n3 0.155672
R1685 VDD2.n60 VDD2.n59 0.155672
C0 VTAIL VN 2.41784f
C1 VDD1 B 1.69117f
C2 VDD1 VDD2 0.666192f
C3 VN w_n2114_n3356# 2.90775f
C4 VTAIL VDD1 5.04146f
C5 VDD1 w_n2114_n3356# 1.76908f
C6 VP B 1.4833f
C7 VDD1 VN 0.148424f
C8 VP VDD2 0.330458f
C9 VDD2 B 1.72063f
C10 VTAIL VP 2.43213f
C11 VP w_n2114_n3356# 3.17688f
C12 VTAIL B 3.61584f
C13 VTAIL VDD2 5.09155f
C14 VN VP 5.40635f
C15 B w_n2114_n3356# 8.71675f
C16 VDD2 w_n2114_n3356# 1.79411f
C17 VN B 1.04111f
C18 VN VDD2 2.75542f
C19 VTAIL w_n2114_n3356# 2.74861f
C20 VDD1 VP 2.9349f
C21 VDD2 VSUBS 0.881743f
C22 VDD1 VSUBS 3.63861f
C23 VTAIL VSUBS 0.993464f
C24 VN VSUBS 7.79751f
C25 VP VSUBS 1.662941f
C26 B VSUBS 3.852406f
C27 w_n2114_n3356# VSUBS 87.341995f
C28 VDD2.n0 VSUBS 0.011486f
C29 VDD2.n1 VSUBS 0.025896f
C30 VDD2.n2 VSUBS 0.011601f
C31 VDD2.n3 VSUBS 0.020389f
C32 VDD2.n4 VSUBS 0.010956f
C33 VDD2.n5 VSUBS 0.025896f
C34 VDD2.n6 VSUBS 0.011601f
C35 VDD2.n7 VSUBS 0.020389f
C36 VDD2.n8 VSUBS 0.010956f
C37 VDD2.n9 VSUBS 0.025896f
C38 VDD2.n10 VSUBS 0.011601f
C39 VDD2.n11 VSUBS 0.020389f
C40 VDD2.n12 VSUBS 0.010956f
C41 VDD2.n13 VSUBS 0.025896f
C42 VDD2.n14 VSUBS 0.011601f
C43 VDD2.n15 VSUBS 0.020389f
C44 VDD2.n16 VSUBS 0.010956f
C45 VDD2.n17 VSUBS 0.025896f
C46 VDD2.n18 VSUBS 0.011601f
C47 VDD2.n19 VSUBS 1.01864f
C48 VDD2.n20 VSUBS 0.010956f
C49 VDD2.t1 VSUBS 0.055287f
C50 VDD2.n21 VSUBS 0.125325f
C51 VDD2.n22 VSUBS 0.016474f
C52 VDD2.n23 VSUBS 0.019422f
C53 VDD2.n24 VSUBS 0.025896f
C54 VDD2.n25 VSUBS 0.011601f
C55 VDD2.n26 VSUBS 0.010956f
C56 VDD2.n27 VSUBS 0.020389f
C57 VDD2.n28 VSUBS 0.020389f
C58 VDD2.n29 VSUBS 0.010956f
C59 VDD2.n30 VSUBS 0.011601f
C60 VDD2.n31 VSUBS 0.025896f
C61 VDD2.n32 VSUBS 0.025896f
C62 VDD2.n33 VSUBS 0.011601f
C63 VDD2.n34 VSUBS 0.010956f
C64 VDD2.n35 VSUBS 0.020389f
C65 VDD2.n36 VSUBS 0.020389f
C66 VDD2.n37 VSUBS 0.010956f
C67 VDD2.n38 VSUBS 0.011601f
C68 VDD2.n39 VSUBS 0.025896f
C69 VDD2.n40 VSUBS 0.025896f
C70 VDD2.n41 VSUBS 0.011601f
C71 VDD2.n42 VSUBS 0.010956f
C72 VDD2.n43 VSUBS 0.020389f
C73 VDD2.n44 VSUBS 0.020389f
C74 VDD2.n45 VSUBS 0.010956f
C75 VDD2.n46 VSUBS 0.011601f
C76 VDD2.n47 VSUBS 0.025896f
C77 VDD2.n48 VSUBS 0.025896f
C78 VDD2.n49 VSUBS 0.011601f
C79 VDD2.n50 VSUBS 0.010956f
C80 VDD2.n51 VSUBS 0.020389f
C81 VDD2.n52 VSUBS 0.020389f
C82 VDD2.n53 VSUBS 0.010956f
C83 VDD2.n54 VSUBS 0.011601f
C84 VDD2.n55 VSUBS 0.025896f
C85 VDD2.n56 VSUBS 0.025896f
C86 VDD2.n57 VSUBS 0.011601f
C87 VDD2.n58 VSUBS 0.010956f
C88 VDD2.n59 VSUBS 0.020389f
C89 VDD2.n60 VSUBS 0.052142f
C90 VDD2.n61 VSUBS 0.010956f
C91 VDD2.n62 VSUBS 0.011601f
C92 VDD2.n63 VSUBS 0.057103f
C93 VDD2.n64 VSUBS 0.58746f
C94 VDD2.n65 VSUBS 0.011486f
C95 VDD2.n66 VSUBS 0.025896f
C96 VDD2.n67 VSUBS 0.011601f
C97 VDD2.n68 VSUBS 0.020389f
C98 VDD2.n69 VSUBS 0.010956f
C99 VDD2.n70 VSUBS 0.025896f
C100 VDD2.n71 VSUBS 0.011601f
C101 VDD2.n72 VSUBS 0.020389f
C102 VDD2.n73 VSUBS 0.010956f
C103 VDD2.n74 VSUBS 0.025896f
C104 VDD2.n75 VSUBS 0.011601f
C105 VDD2.n76 VSUBS 0.020389f
C106 VDD2.n77 VSUBS 0.010956f
C107 VDD2.n78 VSUBS 0.025896f
C108 VDD2.n79 VSUBS 0.011601f
C109 VDD2.n80 VSUBS 0.020389f
C110 VDD2.n81 VSUBS 0.010956f
C111 VDD2.n82 VSUBS 0.025896f
C112 VDD2.n83 VSUBS 0.011601f
C113 VDD2.n84 VSUBS 1.01864f
C114 VDD2.n85 VSUBS 0.010956f
C115 VDD2.t0 VSUBS 0.055287f
C116 VDD2.n86 VSUBS 0.125325f
C117 VDD2.n87 VSUBS 0.016474f
C118 VDD2.n88 VSUBS 0.019422f
C119 VDD2.n89 VSUBS 0.025896f
C120 VDD2.n90 VSUBS 0.011601f
C121 VDD2.n91 VSUBS 0.010956f
C122 VDD2.n92 VSUBS 0.020389f
C123 VDD2.n93 VSUBS 0.020389f
C124 VDD2.n94 VSUBS 0.010956f
C125 VDD2.n95 VSUBS 0.011601f
C126 VDD2.n96 VSUBS 0.025896f
C127 VDD2.n97 VSUBS 0.025896f
C128 VDD2.n98 VSUBS 0.011601f
C129 VDD2.n99 VSUBS 0.010956f
C130 VDD2.n100 VSUBS 0.020389f
C131 VDD2.n101 VSUBS 0.020389f
C132 VDD2.n102 VSUBS 0.010956f
C133 VDD2.n103 VSUBS 0.011601f
C134 VDD2.n104 VSUBS 0.025896f
C135 VDD2.n105 VSUBS 0.025896f
C136 VDD2.n106 VSUBS 0.011601f
C137 VDD2.n107 VSUBS 0.010956f
C138 VDD2.n108 VSUBS 0.020389f
C139 VDD2.n109 VSUBS 0.020389f
C140 VDD2.n110 VSUBS 0.010956f
C141 VDD2.n111 VSUBS 0.011601f
C142 VDD2.n112 VSUBS 0.025896f
C143 VDD2.n113 VSUBS 0.025896f
C144 VDD2.n114 VSUBS 0.011601f
C145 VDD2.n115 VSUBS 0.010956f
C146 VDD2.n116 VSUBS 0.020389f
C147 VDD2.n117 VSUBS 0.020389f
C148 VDD2.n118 VSUBS 0.010956f
C149 VDD2.n119 VSUBS 0.011601f
C150 VDD2.n120 VSUBS 0.025896f
C151 VDD2.n121 VSUBS 0.025896f
C152 VDD2.n122 VSUBS 0.011601f
C153 VDD2.n123 VSUBS 0.010956f
C154 VDD2.n124 VSUBS 0.020389f
C155 VDD2.n125 VSUBS 0.052142f
C156 VDD2.n126 VSUBS 0.010956f
C157 VDD2.n127 VSUBS 0.011601f
C158 VDD2.n128 VSUBS 0.057103f
C159 VDD2.n129 VSUBS 0.052248f
C160 VDD2.n130 VSUBS 2.49075f
C161 VN.t0 VSUBS 3.7302f
C162 VN.t1 VSUBS 4.36985f
C163 VDD1.n0 VSUBS 0.011377f
C164 VDD1.n1 VSUBS 0.025652f
C165 VDD1.n2 VSUBS 0.011491f
C166 VDD1.n3 VSUBS 0.020197f
C167 VDD1.n4 VSUBS 0.010853f
C168 VDD1.n5 VSUBS 0.025652f
C169 VDD1.n6 VSUBS 0.011491f
C170 VDD1.n7 VSUBS 0.020197f
C171 VDD1.n8 VSUBS 0.010853f
C172 VDD1.n9 VSUBS 0.025652f
C173 VDD1.n10 VSUBS 0.011491f
C174 VDD1.n11 VSUBS 0.020197f
C175 VDD1.n12 VSUBS 0.010853f
C176 VDD1.n13 VSUBS 0.025652f
C177 VDD1.n14 VSUBS 0.011491f
C178 VDD1.n15 VSUBS 0.020197f
C179 VDD1.n16 VSUBS 0.010853f
C180 VDD1.n17 VSUBS 0.025652f
C181 VDD1.n18 VSUBS 0.011491f
C182 VDD1.n19 VSUBS 1.00902f
C183 VDD1.n20 VSUBS 0.010853f
C184 VDD1.t0 VSUBS 0.054765f
C185 VDD1.n21 VSUBS 0.124142f
C186 VDD1.n22 VSUBS 0.016319f
C187 VDD1.n23 VSUBS 0.019239f
C188 VDD1.n24 VSUBS 0.025652f
C189 VDD1.n25 VSUBS 0.011491f
C190 VDD1.n26 VSUBS 0.010853f
C191 VDD1.n27 VSUBS 0.020197f
C192 VDD1.n28 VSUBS 0.020197f
C193 VDD1.n29 VSUBS 0.010853f
C194 VDD1.n30 VSUBS 0.011491f
C195 VDD1.n31 VSUBS 0.025652f
C196 VDD1.n32 VSUBS 0.025652f
C197 VDD1.n33 VSUBS 0.011491f
C198 VDD1.n34 VSUBS 0.010853f
C199 VDD1.n35 VSUBS 0.020197f
C200 VDD1.n36 VSUBS 0.020197f
C201 VDD1.n37 VSUBS 0.010853f
C202 VDD1.n38 VSUBS 0.011491f
C203 VDD1.n39 VSUBS 0.025652f
C204 VDD1.n40 VSUBS 0.025652f
C205 VDD1.n41 VSUBS 0.011491f
C206 VDD1.n42 VSUBS 0.010853f
C207 VDD1.n43 VSUBS 0.020197f
C208 VDD1.n44 VSUBS 0.020197f
C209 VDD1.n45 VSUBS 0.010853f
C210 VDD1.n46 VSUBS 0.011491f
C211 VDD1.n47 VSUBS 0.025652f
C212 VDD1.n48 VSUBS 0.025652f
C213 VDD1.n49 VSUBS 0.011491f
C214 VDD1.n50 VSUBS 0.010853f
C215 VDD1.n51 VSUBS 0.020197f
C216 VDD1.n52 VSUBS 0.020197f
C217 VDD1.n53 VSUBS 0.010853f
C218 VDD1.n54 VSUBS 0.011491f
C219 VDD1.n55 VSUBS 0.025652f
C220 VDD1.n56 VSUBS 0.025652f
C221 VDD1.n57 VSUBS 0.011491f
C222 VDD1.n58 VSUBS 0.010853f
C223 VDD1.n59 VSUBS 0.020197f
C224 VDD1.n60 VSUBS 0.05165f
C225 VDD1.n61 VSUBS 0.010853f
C226 VDD1.n62 VSUBS 0.011491f
C227 VDD1.n63 VSUBS 0.056564f
C228 VDD1.n64 VSUBS 0.052856f
C229 VDD1.n65 VSUBS 0.011377f
C230 VDD1.n66 VSUBS 0.025652f
C231 VDD1.n67 VSUBS 0.011491f
C232 VDD1.n68 VSUBS 0.020197f
C233 VDD1.n69 VSUBS 0.010853f
C234 VDD1.n70 VSUBS 0.025652f
C235 VDD1.n71 VSUBS 0.011491f
C236 VDD1.n72 VSUBS 0.020197f
C237 VDD1.n73 VSUBS 0.010853f
C238 VDD1.n74 VSUBS 0.025652f
C239 VDD1.n75 VSUBS 0.011491f
C240 VDD1.n76 VSUBS 0.020197f
C241 VDD1.n77 VSUBS 0.010853f
C242 VDD1.n78 VSUBS 0.025652f
C243 VDD1.n79 VSUBS 0.011491f
C244 VDD1.n80 VSUBS 0.020197f
C245 VDD1.n81 VSUBS 0.010853f
C246 VDD1.n82 VSUBS 0.025652f
C247 VDD1.n83 VSUBS 0.011491f
C248 VDD1.n84 VSUBS 1.00902f
C249 VDD1.n85 VSUBS 0.010853f
C250 VDD1.t1 VSUBS 0.054765f
C251 VDD1.n86 VSUBS 0.124142f
C252 VDD1.n87 VSUBS 0.016319f
C253 VDD1.n88 VSUBS 0.019239f
C254 VDD1.n89 VSUBS 0.025652f
C255 VDD1.n90 VSUBS 0.011491f
C256 VDD1.n91 VSUBS 0.010853f
C257 VDD1.n92 VSUBS 0.020197f
C258 VDD1.n93 VSUBS 0.020197f
C259 VDD1.n94 VSUBS 0.010853f
C260 VDD1.n95 VSUBS 0.011491f
C261 VDD1.n96 VSUBS 0.025652f
C262 VDD1.n97 VSUBS 0.025652f
C263 VDD1.n98 VSUBS 0.011491f
C264 VDD1.n99 VSUBS 0.010853f
C265 VDD1.n100 VSUBS 0.020197f
C266 VDD1.n101 VSUBS 0.020197f
C267 VDD1.n102 VSUBS 0.010853f
C268 VDD1.n103 VSUBS 0.011491f
C269 VDD1.n104 VSUBS 0.025652f
C270 VDD1.n105 VSUBS 0.025652f
C271 VDD1.n106 VSUBS 0.011491f
C272 VDD1.n107 VSUBS 0.010853f
C273 VDD1.n108 VSUBS 0.020197f
C274 VDD1.n109 VSUBS 0.020197f
C275 VDD1.n110 VSUBS 0.010853f
C276 VDD1.n111 VSUBS 0.011491f
C277 VDD1.n112 VSUBS 0.025652f
C278 VDD1.n113 VSUBS 0.025652f
C279 VDD1.n114 VSUBS 0.011491f
C280 VDD1.n115 VSUBS 0.010853f
C281 VDD1.n116 VSUBS 0.020197f
C282 VDD1.n117 VSUBS 0.020197f
C283 VDD1.n118 VSUBS 0.010853f
C284 VDD1.n119 VSUBS 0.011491f
C285 VDD1.n120 VSUBS 0.025652f
C286 VDD1.n121 VSUBS 0.025652f
C287 VDD1.n122 VSUBS 0.011491f
C288 VDD1.n123 VSUBS 0.010853f
C289 VDD1.n124 VSUBS 0.020197f
C290 VDD1.n125 VSUBS 0.05165f
C291 VDD1.n126 VSUBS 0.010853f
C292 VDD1.n127 VSUBS 0.011491f
C293 VDD1.n128 VSUBS 0.056564f
C294 VDD1.n129 VSUBS 0.620199f
C295 VTAIL.n0 VSUBS 0.016509f
C296 VTAIL.n1 VSUBS 0.037222f
C297 VTAIL.n2 VSUBS 0.016674f
C298 VTAIL.n3 VSUBS 0.029306f
C299 VTAIL.n4 VSUBS 0.015748f
C300 VTAIL.n5 VSUBS 0.037222f
C301 VTAIL.n6 VSUBS 0.016674f
C302 VTAIL.n7 VSUBS 0.029306f
C303 VTAIL.n8 VSUBS 0.015748f
C304 VTAIL.n9 VSUBS 0.037222f
C305 VTAIL.n10 VSUBS 0.016674f
C306 VTAIL.n11 VSUBS 0.029306f
C307 VTAIL.n12 VSUBS 0.015748f
C308 VTAIL.n13 VSUBS 0.037222f
C309 VTAIL.n14 VSUBS 0.016674f
C310 VTAIL.n15 VSUBS 0.029306f
C311 VTAIL.n16 VSUBS 0.015748f
C312 VTAIL.n17 VSUBS 0.037222f
C313 VTAIL.n18 VSUBS 0.016674f
C314 VTAIL.n19 VSUBS 1.46413f
C315 VTAIL.n20 VSUBS 0.015748f
C316 VTAIL.t3 VSUBS 0.079466f
C317 VTAIL.n21 VSUBS 0.180136f
C318 VTAIL.n22 VSUBS 0.023679f
C319 VTAIL.n23 VSUBS 0.027916f
C320 VTAIL.n24 VSUBS 0.037222f
C321 VTAIL.n25 VSUBS 0.016674f
C322 VTAIL.n26 VSUBS 0.015748f
C323 VTAIL.n27 VSUBS 0.029306f
C324 VTAIL.n28 VSUBS 0.029306f
C325 VTAIL.n29 VSUBS 0.015748f
C326 VTAIL.n30 VSUBS 0.016674f
C327 VTAIL.n31 VSUBS 0.037222f
C328 VTAIL.n32 VSUBS 0.037222f
C329 VTAIL.n33 VSUBS 0.016674f
C330 VTAIL.n34 VSUBS 0.015748f
C331 VTAIL.n35 VSUBS 0.029306f
C332 VTAIL.n36 VSUBS 0.029306f
C333 VTAIL.n37 VSUBS 0.015748f
C334 VTAIL.n38 VSUBS 0.016674f
C335 VTAIL.n39 VSUBS 0.037222f
C336 VTAIL.n40 VSUBS 0.037222f
C337 VTAIL.n41 VSUBS 0.016674f
C338 VTAIL.n42 VSUBS 0.015748f
C339 VTAIL.n43 VSUBS 0.029306f
C340 VTAIL.n44 VSUBS 0.029306f
C341 VTAIL.n45 VSUBS 0.015748f
C342 VTAIL.n46 VSUBS 0.016674f
C343 VTAIL.n47 VSUBS 0.037222f
C344 VTAIL.n48 VSUBS 0.037222f
C345 VTAIL.n49 VSUBS 0.016674f
C346 VTAIL.n50 VSUBS 0.015748f
C347 VTAIL.n51 VSUBS 0.029306f
C348 VTAIL.n52 VSUBS 0.029306f
C349 VTAIL.n53 VSUBS 0.015748f
C350 VTAIL.n54 VSUBS 0.016674f
C351 VTAIL.n55 VSUBS 0.037222f
C352 VTAIL.n56 VSUBS 0.037222f
C353 VTAIL.n57 VSUBS 0.016674f
C354 VTAIL.n58 VSUBS 0.015748f
C355 VTAIL.n59 VSUBS 0.029306f
C356 VTAIL.n60 VSUBS 0.074946f
C357 VTAIL.n61 VSUBS 0.015748f
C358 VTAIL.n62 VSUBS 0.016674f
C359 VTAIL.n63 VSUBS 0.082076f
C360 VTAIL.n64 VSUBS 0.054898f
C361 VTAIL.n65 VSUBS 1.97152f
C362 VTAIL.n66 VSUBS 0.016509f
C363 VTAIL.n67 VSUBS 0.037222f
C364 VTAIL.n68 VSUBS 0.016674f
C365 VTAIL.n69 VSUBS 0.029306f
C366 VTAIL.n70 VSUBS 0.015748f
C367 VTAIL.n71 VSUBS 0.037222f
C368 VTAIL.n72 VSUBS 0.016674f
C369 VTAIL.n73 VSUBS 0.029306f
C370 VTAIL.n74 VSUBS 0.015748f
C371 VTAIL.n75 VSUBS 0.037222f
C372 VTAIL.n76 VSUBS 0.016674f
C373 VTAIL.n77 VSUBS 0.029306f
C374 VTAIL.n78 VSUBS 0.015748f
C375 VTAIL.n79 VSUBS 0.037222f
C376 VTAIL.n80 VSUBS 0.016674f
C377 VTAIL.n81 VSUBS 0.029306f
C378 VTAIL.n82 VSUBS 0.015748f
C379 VTAIL.n83 VSUBS 0.037222f
C380 VTAIL.n84 VSUBS 0.016674f
C381 VTAIL.n85 VSUBS 1.46413f
C382 VTAIL.n86 VSUBS 0.015748f
C383 VTAIL.t1 VSUBS 0.079466f
C384 VTAIL.n87 VSUBS 0.180136f
C385 VTAIL.n88 VSUBS 0.023679f
C386 VTAIL.n89 VSUBS 0.027916f
C387 VTAIL.n90 VSUBS 0.037222f
C388 VTAIL.n91 VSUBS 0.016674f
C389 VTAIL.n92 VSUBS 0.015748f
C390 VTAIL.n93 VSUBS 0.029306f
C391 VTAIL.n94 VSUBS 0.029306f
C392 VTAIL.n95 VSUBS 0.015748f
C393 VTAIL.n96 VSUBS 0.016674f
C394 VTAIL.n97 VSUBS 0.037222f
C395 VTAIL.n98 VSUBS 0.037222f
C396 VTAIL.n99 VSUBS 0.016674f
C397 VTAIL.n100 VSUBS 0.015748f
C398 VTAIL.n101 VSUBS 0.029306f
C399 VTAIL.n102 VSUBS 0.029306f
C400 VTAIL.n103 VSUBS 0.015748f
C401 VTAIL.n104 VSUBS 0.016674f
C402 VTAIL.n105 VSUBS 0.037222f
C403 VTAIL.n106 VSUBS 0.037222f
C404 VTAIL.n107 VSUBS 0.016674f
C405 VTAIL.n108 VSUBS 0.015748f
C406 VTAIL.n109 VSUBS 0.029306f
C407 VTAIL.n110 VSUBS 0.029306f
C408 VTAIL.n111 VSUBS 0.015748f
C409 VTAIL.n112 VSUBS 0.016674f
C410 VTAIL.n113 VSUBS 0.037222f
C411 VTAIL.n114 VSUBS 0.037222f
C412 VTAIL.n115 VSUBS 0.016674f
C413 VTAIL.n116 VSUBS 0.015748f
C414 VTAIL.n117 VSUBS 0.029306f
C415 VTAIL.n118 VSUBS 0.029306f
C416 VTAIL.n119 VSUBS 0.015748f
C417 VTAIL.n120 VSUBS 0.016674f
C418 VTAIL.n121 VSUBS 0.037222f
C419 VTAIL.n122 VSUBS 0.037222f
C420 VTAIL.n123 VSUBS 0.016674f
C421 VTAIL.n124 VSUBS 0.015748f
C422 VTAIL.n125 VSUBS 0.029306f
C423 VTAIL.n126 VSUBS 0.074946f
C424 VTAIL.n127 VSUBS 0.015748f
C425 VTAIL.n128 VSUBS 0.016674f
C426 VTAIL.n129 VSUBS 0.082076f
C427 VTAIL.n130 VSUBS 0.054898f
C428 VTAIL.n131 VSUBS 2.02423f
C429 VTAIL.n132 VSUBS 0.016509f
C430 VTAIL.n133 VSUBS 0.037222f
C431 VTAIL.n134 VSUBS 0.016674f
C432 VTAIL.n135 VSUBS 0.029306f
C433 VTAIL.n136 VSUBS 0.015748f
C434 VTAIL.n137 VSUBS 0.037222f
C435 VTAIL.n138 VSUBS 0.016674f
C436 VTAIL.n139 VSUBS 0.029306f
C437 VTAIL.n140 VSUBS 0.015748f
C438 VTAIL.n141 VSUBS 0.037222f
C439 VTAIL.n142 VSUBS 0.016674f
C440 VTAIL.n143 VSUBS 0.029306f
C441 VTAIL.n144 VSUBS 0.015748f
C442 VTAIL.n145 VSUBS 0.037222f
C443 VTAIL.n146 VSUBS 0.016674f
C444 VTAIL.n147 VSUBS 0.029306f
C445 VTAIL.n148 VSUBS 0.015748f
C446 VTAIL.n149 VSUBS 0.037222f
C447 VTAIL.n150 VSUBS 0.016674f
C448 VTAIL.n151 VSUBS 1.46413f
C449 VTAIL.n152 VSUBS 0.015748f
C450 VTAIL.t2 VSUBS 0.079466f
C451 VTAIL.n153 VSUBS 0.180136f
C452 VTAIL.n154 VSUBS 0.023679f
C453 VTAIL.n155 VSUBS 0.027916f
C454 VTAIL.n156 VSUBS 0.037222f
C455 VTAIL.n157 VSUBS 0.016674f
C456 VTAIL.n158 VSUBS 0.015748f
C457 VTAIL.n159 VSUBS 0.029306f
C458 VTAIL.n160 VSUBS 0.029306f
C459 VTAIL.n161 VSUBS 0.015748f
C460 VTAIL.n162 VSUBS 0.016674f
C461 VTAIL.n163 VSUBS 0.037222f
C462 VTAIL.n164 VSUBS 0.037222f
C463 VTAIL.n165 VSUBS 0.016674f
C464 VTAIL.n166 VSUBS 0.015748f
C465 VTAIL.n167 VSUBS 0.029306f
C466 VTAIL.n168 VSUBS 0.029306f
C467 VTAIL.n169 VSUBS 0.015748f
C468 VTAIL.n170 VSUBS 0.016674f
C469 VTAIL.n171 VSUBS 0.037222f
C470 VTAIL.n172 VSUBS 0.037222f
C471 VTAIL.n173 VSUBS 0.016674f
C472 VTAIL.n174 VSUBS 0.015748f
C473 VTAIL.n175 VSUBS 0.029306f
C474 VTAIL.n176 VSUBS 0.029306f
C475 VTAIL.n177 VSUBS 0.015748f
C476 VTAIL.n178 VSUBS 0.016674f
C477 VTAIL.n179 VSUBS 0.037222f
C478 VTAIL.n180 VSUBS 0.037222f
C479 VTAIL.n181 VSUBS 0.016674f
C480 VTAIL.n182 VSUBS 0.015748f
C481 VTAIL.n183 VSUBS 0.029306f
C482 VTAIL.n184 VSUBS 0.029306f
C483 VTAIL.n185 VSUBS 0.015748f
C484 VTAIL.n186 VSUBS 0.016674f
C485 VTAIL.n187 VSUBS 0.037222f
C486 VTAIL.n188 VSUBS 0.037222f
C487 VTAIL.n189 VSUBS 0.016674f
C488 VTAIL.n190 VSUBS 0.015748f
C489 VTAIL.n191 VSUBS 0.029306f
C490 VTAIL.n192 VSUBS 0.074946f
C491 VTAIL.n193 VSUBS 0.015748f
C492 VTAIL.n194 VSUBS 0.016674f
C493 VTAIL.n195 VSUBS 0.082076f
C494 VTAIL.n196 VSUBS 0.054898f
C495 VTAIL.n197 VSUBS 1.79141f
C496 VTAIL.n198 VSUBS 0.016509f
C497 VTAIL.n199 VSUBS 0.037222f
C498 VTAIL.n200 VSUBS 0.016674f
C499 VTAIL.n201 VSUBS 0.029306f
C500 VTAIL.n202 VSUBS 0.015748f
C501 VTAIL.n203 VSUBS 0.037222f
C502 VTAIL.n204 VSUBS 0.016674f
C503 VTAIL.n205 VSUBS 0.029306f
C504 VTAIL.n206 VSUBS 0.015748f
C505 VTAIL.n207 VSUBS 0.037222f
C506 VTAIL.n208 VSUBS 0.016674f
C507 VTAIL.n209 VSUBS 0.029306f
C508 VTAIL.n210 VSUBS 0.015748f
C509 VTAIL.n211 VSUBS 0.037222f
C510 VTAIL.n212 VSUBS 0.016674f
C511 VTAIL.n213 VSUBS 0.029306f
C512 VTAIL.n214 VSUBS 0.015748f
C513 VTAIL.n215 VSUBS 0.037222f
C514 VTAIL.n216 VSUBS 0.016674f
C515 VTAIL.n217 VSUBS 1.46413f
C516 VTAIL.n218 VSUBS 0.015748f
C517 VTAIL.t0 VSUBS 0.079466f
C518 VTAIL.n219 VSUBS 0.180136f
C519 VTAIL.n220 VSUBS 0.023679f
C520 VTAIL.n221 VSUBS 0.027916f
C521 VTAIL.n222 VSUBS 0.037222f
C522 VTAIL.n223 VSUBS 0.016674f
C523 VTAIL.n224 VSUBS 0.015748f
C524 VTAIL.n225 VSUBS 0.029306f
C525 VTAIL.n226 VSUBS 0.029306f
C526 VTAIL.n227 VSUBS 0.015748f
C527 VTAIL.n228 VSUBS 0.016674f
C528 VTAIL.n229 VSUBS 0.037222f
C529 VTAIL.n230 VSUBS 0.037222f
C530 VTAIL.n231 VSUBS 0.016674f
C531 VTAIL.n232 VSUBS 0.015748f
C532 VTAIL.n233 VSUBS 0.029306f
C533 VTAIL.n234 VSUBS 0.029306f
C534 VTAIL.n235 VSUBS 0.015748f
C535 VTAIL.n236 VSUBS 0.016674f
C536 VTAIL.n237 VSUBS 0.037222f
C537 VTAIL.n238 VSUBS 0.037222f
C538 VTAIL.n239 VSUBS 0.016674f
C539 VTAIL.n240 VSUBS 0.015748f
C540 VTAIL.n241 VSUBS 0.029306f
C541 VTAIL.n242 VSUBS 0.029306f
C542 VTAIL.n243 VSUBS 0.015748f
C543 VTAIL.n244 VSUBS 0.016674f
C544 VTAIL.n245 VSUBS 0.037222f
C545 VTAIL.n246 VSUBS 0.037222f
C546 VTAIL.n247 VSUBS 0.016674f
C547 VTAIL.n248 VSUBS 0.015748f
C548 VTAIL.n249 VSUBS 0.029306f
C549 VTAIL.n250 VSUBS 0.029306f
C550 VTAIL.n251 VSUBS 0.015748f
C551 VTAIL.n252 VSUBS 0.016674f
C552 VTAIL.n253 VSUBS 0.037222f
C553 VTAIL.n254 VSUBS 0.037222f
C554 VTAIL.n255 VSUBS 0.016674f
C555 VTAIL.n256 VSUBS 0.015748f
C556 VTAIL.n257 VSUBS 0.029306f
C557 VTAIL.n258 VSUBS 0.074946f
C558 VTAIL.n259 VSUBS 0.015748f
C559 VTAIL.n260 VSUBS 0.016674f
C560 VTAIL.n261 VSUBS 0.082076f
C561 VTAIL.n262 VSUBS 0.054898f
C562 VTAIL.n263 VSUBS 1.68335f
C563 VP.t1 VSUBS 4.51391f
C564 VP.t0 VSUBS 3.85433f
C565 VP.n0 VSUBS 5.43523f
C566 B.n0 VSUBS 0.003874f
C567 B.n1 VSUBS 0.003874f
C568 B.n2 VSUBS 0.006127f
C569 B.n3 VSUBS 0.006127f
C570 B.n4 VSUBS 0.006127f
C571 B.n5 VSUBS 0.006127f
C572 B.n6 VSUBS 0.006127f
C573 B.n7 VSUBS 0.006127f
C574 B.n8 VSUBS 0.006127f
C575 B.n9 VSUBS 0.006127f
C576 B.n10 VSUBS 0.006127f
C577 B.n11 VSUBS 0.006127f
C578 B.n12 VSUBS 0.006127f
C579 B.n13 VSUBS 0.006127f
C580 B.n14 VSUBS 0.014616f
C581 B.n15 VSUBS 0.006127f
C582 B.n16 VSUBS 0.006127f
C583 B.n17 VSUBS 0.006127f
C584 B.n18 VSUBS 0.006127f
C585 B.n19 VSUBS 0.006127f
C586 B.n20 VSUBS 0.006127f
C587 B.n21 VSUBS 0.006127f
C588 B.n22 VSUBS 0.006127f
C589 B.n23 VSUBS 0.006127f
C590 B.n24 VSUBS 0.006127f
C591 B.n25 VSUBS 0.006127f
C592 B.n26 VSUBS 0.006127f
C593 B.n27 VSUBS 0.006127f
C594 B.n28 VSUBS 0.006127f
C595 B.n29 VSUBS 0.006127f
C596 B.n30 VSUBS 0.006127f
C597 B.n31 VSUBS 0.006127f
C598 B.n32 VSUBS 0.006127f
C599 B.n33 VSUBS 0.006127f
C600 B.n34 VSUBS 0.006127f
C601 B.n35 VSUBS 0.006127f
C602 B.t8 VSUBS 0.183345f
C603 B.t7 VSUBS 0.210558f
C604 B.t6 VSUBS 1.20242f
C605 B.n36 VSUBS 0.334454f
C606 B.n37 VSUBS 0.21962f
C607 B.n38 VSUBS 0.006127f
C608 B.n39 VSUBS 0.006127f
C609 B.n40 VSUBS 0.006127f
C610 B.n41 VSUBS 0.006127f
C611 B.t5 VSUBS 0.183347f
C612 B.t4 VSUBS 0.21056f
C613 B.t3 VSUBS 1.20242f
C614 B.n42 VSUBS 0.334451f
C615 B.n43 VSUBS 0.219618f
C616 B.n44 VSUBS 0.014195f
C617 B.n45 VSUBS 0.006127f
C618 B.n46 VSUBS 0.006127f
C619 B.n47 VSUBS 0.006127f
C620 B.n48 VSUBS 0.006127f
C621 B.n49 VSUBS 0.006127f
C622 B.n50 VSUBS 0.006127f
C623 B.n51 VSUBS 0.006127f
C624 B.n52 VSUBS 0.006127f
C625 B.n53 VSUBS 0.006127f
C626 B.n54 VSUBS 0.006127f
C627 B.n55 VSUBS 0.006127f
C628 B.n56 VSUBS 0.006127f
C629 B.n57 VSUBS 0.006127f
C630 B.n58 VSUBS 0.006127f
C631 B.n59 VSUBS 0.006127f
C632 B.n60 VSUBS 0.006127f
C633 B.n61 VSUBS 0.006127f
C634 B.n62 VSUBS 0.006127f
C635 B.n63 VSUBS 0.006127f
C636 B.n64 VSUBS 0.006127f
C637 B.n65 VSUBS 0.014616f
C638 B.n66 VSUBS 0.006127f
C639 B.n67 VSUBS 0.006127f
C640 B.n68 VSUBS 0.006127f
C641 B.n69 VSUBS 0.006127f
C642 B.n70 VSUBS 0.006127f
C643 B.n71 VSUBS 0.006127f
C644 B.n72 VSUBS 0.006127f
C645 B.n73 VSUBS 0.006127f
C646 B.n74 VSUBS 0.006127f
C647 B.n75 VSUBS 0.006127f
C648 B.n76 VSUBS 0.006127f
C649 B.n77 VSUBS 0.006127f
C650 B.n78 VSUBS 0.006127f
C651 B.n79 VSUBS 0.006127f
C652 B.n80 VSUBS 0.006127f
C653 B.n81 VSUBS 0.006127f
C654 B.n82 VSUBS 0.006127f
C655 B.n83 VSUBS 0.006127f
C656 B.n84 VSUBS 0.006127f
C657 B.n85 VSUBS 0.006127f
C658 B.n86 VSUBS 0.006127f
C659 B.n87 VSUBS 0.006127f
C660 B.n88 VSUBS 0.006127f
C661 B.n89 VSUBS 0.006127f
C662 B.n90 VSUBS 0.014616f
C663 B.n91 VSUBS 0.006127f
C664 B.n92 VSUBS 0.006127f
C665 B.n93 VSUBS 0.006127f
C666 B.n94 VSUBS 0.006127f
C667 B.n95 VSUBS 0.006127f
C668 B.n96 VSUBS 0.006127f
C669 B.n97 VSUBS 0.006127f
C670 B.n98 VSUBS 0.006127f
C671 B.n99 VSUBS 0.006127f
C672 B.n100 VSUBS 0.006127f
C673 B.n101 VSUBS 0.006127f
C674 B.n102 VSUBS 0.006127f
C675 B.n103 VSUBS 0.006127f
C676 B.n104 VSUBS 0.006127f
C677 B.n105 VSUBS 0.006127f
C678 B.n106 VSUBS 0.006127f
C679 B.n107 VSUBS 0.006127f
C680 B.n108 VSUBS 0.006127f
C681 B.n109 VSUBS 0.006127f
C682 B.n110 VSUBS 0.006127f
C683 B.n111 VSUBS 0.006127f
C684 B.t1 VSUBS 0.183347f
C685 B.t2 VSUBS 0.21056f
C686 B.t0 VSUBS 1.20242f
C687 B.n112 VSUBS 0.334451f
C688 B.n113 VSUBS 0.219618f
C689 B.n114 VSUBS 0.006127f
C690 B.n115 VSUBS 0.006127f
C691 B.n116 VSUBS 0.006127f
C692 B.n117 VSUBS 0.006127f
C693 B.t10 VSUBS 0.183345f
C694 B.t11 VSUBS 0.210558f
C695 B.t9 VSUBS 1.20242f
C696 B.n118 VSUBS 0.334454f
C697 B.n119 VSUBS 0.21962f
C698 B.n120 VSUBS 0.014195f
C699 B.n121 VSUBS 0.006127f
C700 B.n122 VSUBS 0.006127f
C701 B.n123 VSUBS 0.006127f
C702 B.n124 VSUBS 0.006127f
C703 B.n125 VSUBS 0.006127f
C704 B.n126 VSUBS 0.006127f
C705 B.n127 VSUBS 0.006127f
C706 B.n128 VSUBS 0.006127f
C707 B.n129 VSUBS 0.006127f
C708 B.n130 VSUBS 0.006127f
C709 B.n131 VSUBS 0.006127f
C710 B.n132 VSUBS 0.006127f
C711 B.n133 VSUBS 0.006127f
C712 B.n134 VSUBS 0.006127f
C713 B.n135 VSUBS 0.006127f
C714 B.n136 VSUBS 0.006127f
C715 B.n137 VSUBS 0.006127f
C716 B.n138 VSUBS 0.006127f
C717 B.n139 VSUBS 0.006127f
C718 B.n140 VSUBS 0.006127f
C719 B.n141 VSUBS 0.014616f
C720 B.n142 VSUBS 0.006127f
C721 B.n143 VSUBS 0.006127f
C722 B.n144 VSUBS 0.006127f
C723 B.n145 VSUBS 0.006127f
C724 B.n146 VSUBS 0.006127f
C725 B.n147 VSUBS 0.006127f
C726 B.n148 VSUBS 0.006127f
C727 B.n149 VSUBS 0.006127f
C728 B.n150 VSUBS 0.006127f
C729 B.n151 VSUBS 0.006127f
C730 B.n152 VSUBS 0.006127f
C731 B.n153 VSUBS 0.006127f
C732 B.n154 VSUBS 0.006127f
C733 B.n155 VSUBS 0.006127f
C734 B.n156 VSUBS 0.006127f
C735 B.n157 VSUBS 0.006127f
C736 B.n158 VSUBS 0.006127f
C737 B.n159 VSUBS 0.006127f
C738 B.n160 VSUBS 0.006127f
C739 B.n161 VSUBS 0.006127f
C740 B.n162 VSUBS 0.006127f
C741 B.n163 VSUBS 0.006127f
C742 B.n164 VSUBS 0.006127f
C743 B.n165 VSUBS 0.006127f
C744 B.n166 VSUBS 0.006127f
C745 B.n167 VSUBS 0.006127f
C746 B.n168 VSUBS 0.006127f
C747 B.n169 VSUBS 0.006127f
C748 B.n170 VSUBS 0.006127f
C749 B.n171 VSUBS 0.006127f
C750 B.n172 VSUBS 0.006127f
C751 B.n173 VSUBS 0.006127f
C752 B.n174 VSUBS 0.006127f
C753 B.n175 VSUBS 0.006127f
C754 B.n176 VSUBS 0.006127f
C755 B.n177 VSUBS 0.006127f
C756 B.n178 VSUBS 0.006127f
C757 B.n179 VSUBS 0.006127f
C758 B.n180 VSUBS 0.006127f
C759 B.n181 VSUBS 0.006127f
C760 B.n182 VSUBS 0.006127f
C761 B.n183 VSUBS 0.006127f
C762 B.n184 VSUBS 0.006127f
C763 B.n185 VSUBS 0.006127f
C764 B.n186 VSUBS 0.006127f
C765 B.n187 VSUBS 0.006127f
C766 B.n188 VSUBS 0.014616f
C767 B.n189 VSUBS 0.014936f
C768 B.n190 VSUBS 0.014936f
C769 B.n191 VSUBS 0.006127f
C770 B.n192 VSUBS 0.006127f
C771 B.n193 VSUBS 0.006127f
C772 B.n194 VSUBS 0.006127f
C773 B.n195 VSUBS 0.006127f
C774 B.n196 VSUBS 0.006127f
C775 B.n197 VSUBS 0.006127f
C776 B.n198 VSUBS 0.006127f
C777 B.n199 VSUBS 0.006127f
C778 B.n200 VSUBS 0.006127f
C779 B.n201 VSUBS 0.006127f
C780 B.n202 VSUBS 0.006127f
C781 B.n203 VSUBS 0.006127f
C782 B.n204 VSUBS 0.006127f
C783 B.n205 VSUBS 0.006127f
C784 B.n206 VSUBS 0.006127f
C785 B.n207 VSUBS 0.006127f
C786 B.n208 VSUBS 0.006127f
C787 B.n209 VSUBS 0.006127f
C788 B.n210 VSUBS 0.006127f
C789 B.n211 VSUBS 0.006127f
C790 B.n212 VSUBS 0.006127f
C791 B.n213 VSUBS 0.006127f
C792 B.n214 VSUBS 0.006127f
C793 B.n215 VSUBS 0.006127f
C794 B.n216 VSUBS 0.006127f
C795 B.n217 VSUBS 0.006127f
C796 B.n218 VSUBS 0.006127f
C797 B.n219 VSUBS 0.006127f
C798 B.n220 VSUBS 0.006127f
C799 B.n221 VSUBS 0.006127f
C800 B.n222 VSUBS 0.006127f
C801 B.n223 VSUBS 0.006127f
C802 B.n224 VSUBS 0.006127f
C803 B.n225 VSUBS 0.006127f
C804 B.n226 VSUBS 0.006127f
C805 B.n227 VSUBS 0.006127f
C806 B.n228 VSUBS 0.006127f
C807 B.n229 VSUBS 0.006127f
C808 B.n230 VSUBS 0.006127f
C809 B.n231 VSUBS 0.006127f
C810 B.n232 VSUBS 0.006127f
C811 B.n233 VSUBS 0.006127f
C812 B.n234 VSUBS 0.006127f
C813 B.n235 VSUBS 0.006127f
C814 B.n236 VSUBS 0.006127f
C815 B.n237 VSUBS 0.006127f
C816 B.n238 VSUBS 0.006127f
C817 B.n239 VSUBS 0.006127f
C818 B.n240 VSUBS 0.006127f
C819 B.n241 VSUBS 0.006127f
C820 B.n242 VSUBS 0.006127f
C821 B.n243 VSUBS 0.006127f
C822 B.n244 VSUBS 0.006127f
C823 B.n245 VSUBS 0.006127f
C824 B.n246 VSUBS 0.006127f
C825 B.n247 VSUBS 0.006127f
C826 B.n248 VSUBS 0.006127f
C827 B.n249 VSUBS 0.005766f
C828 B.n250 VSUBS 0.006127f
C829 B.n251 VSUBS 0.006127f
C830 B.n252 VSUBS 0.003424f
C831 B.n253 VSUBS 0.006127f
C832 B.n254 VSUBS 0.006127f
C833 B.n255 VSUBS 0.006127f
C834 B.n256 VSUBS 0.006127f
C835 B.n257 VSUBS 0.006127f
C836 B.n258 VSUBS 0.006127f
C837 B.n259 VSUBS 0.006127f
C838 B.n260 VSUBS 0.006127f
C839 B.n261 VSUBS 0.006127f
C840 B.n262 VSUBS 0.006127f
C841 B.n263 VSUBS 0.006127f
C842 B.n264 VSUBS 0.006127f
C843 B.n265 VSUBS 0.003424f
C844 B.n266 VSUBS 0.014195f
C845 B.n267 VSUBS 0.005766f
C846 B.n268 VSUBS 0.006127f
C847 B.n269 VSUBS 0.006127f
C848 B.n270 VSUBS 0.006127f
C849 B.n271 VSUBS 0.006127f
C850 B.n272 VSUBS 0.006127f
C851 B.n273 VSUBS 0.006127f
C852 B.n274 VSUBS 0.006127f
C853 B.n275 VSUBS 0.006127f
C854 B.n276 VSUBS 0.006127f
C855 B.n277 VSUBS 0.006127f
C856 B.n278 VSUBS 0.006127f
C857 B.n279 VSUBS 0.006127f
C858 B.n280 VSUBS 0.006127f
C859 B.n281 VSUBS 0.006127f
C860 B.n282 VSUBS 0.006127f
C861 B.n283 VSUBS 0.006127f
C862 B.n284 VSUBS 0.006127f
C863 B.n285 VSUBS 0.006127f
C864 B.n286 VSUBS 0.006127f
C865 B.n287 VSUBS 0.006127f
C866 B.n288 VSUBS 0.006127f
C867 B.n289 VSUBS 0.006127f
C868 B.n290 VSUBS 0.006127f
C869 B.n291 VSUBS 0.006127f
C870 B.n292 VSUBS 0.006127f
C871 B.n293 VSUBS 0.006127f
C872 B.n294 VSUBS 0.006127f
C873 B.n295 VSUBS 0.006127f
C874 B.n296 VSUBS 0.006127f
C875 B.n297 VSUBS 0.006127f
C876 B.n298 VSUBS 0.006127f
C877 B.n299 VSUBS 0.006127f
C878 B.n300 VSUBS 0.006127f
C879 B.n301 VSUBS 0.006127f
C880 B.n302 VSUBS 0.006127f
C881 B.n303 VSUBS 0.006127f
C882 B.n304 VSUBS 0.006127f
C883 B.n305 VSUBS 0.006127f
C884 B.n306 VSUBS 0.006127f
C885 B.n307 VSUBS 0.006127f
C886 B.n308 VSUBS 0.006127f
C887 B.n309 VSUBS 0.006127f
C888 B.n310 VSUBS 0.006127f
C889 B.n311 VSUBS 0.006127f
C890 B.n312 VSUBS 0.006127f
C891 B.n313 VSUBS 0.006127f
C892 B.n314 VSUBS 0.006127f
C893 B.n315 VSUBS 0.006127f
C894 B.n316 VSUBS 0.006127f
C895 B.n317 VSUBS 0.006127f
C896 B.n318 VSUBS 0.006127f
C897 B.n319 VSUBS 0.006127f
C898 B.n320 VSUBS 0.006127f
C899 B.n321 VSUBS 0.006127f
C900 B.n322 VSUBS 0.006127f
C901 B.n323 VSUBS 0.006127f
C902 B.n324 VSUBS 0.006127f
C903 B.n325 VSUBS 0.006127f
C904 B.n326 VSUBS 0.006127f
C905 B.n327 VSUBS 0.014936f
C906 B.n328 VSUBS 0.014936f
C907 B.n329 VSUBS 0.014616f
C908 B.n330 VSUBS 0.006127f
C909 B.n331 VSUBS 0.006127f
C910 B.n332 VSUBS 0.006127f
C911 B.n333 VSUBS 0.006127f
C912 B.n334 VSUBS 0.006127f
C913 B.n335 VSUBS 0.006127f
C914 B.n336 VSUBS 0.006127f
C915 B.n337 VSUBS 0.006127f
C916 B.n338 VSUBS 0.006127f
C917 B.n339 VSUBS 0.006127f
C918 B.n340 VSUBS 0.006127f
C919 B.n341 VSUBS 0.006127f
C920 B.n342 VSUBS 0.006127f
C921 B.n343 VSUBS 0.006127f
C922 B.n344 VSUBS 0.006127f
C923 B.n345 VSUBS 0.006127f
C924 B.n346 VSUBS 0.006127f
C925 B.n347 VSUBS 0.006127f
C926 B.n348 VSUBS 0.006127f
C927 B.n349 VSUBS 0.006127f
C928 B.n350 VSUBS 0.006127f
C929 B.n351 VSUBS 0.006127f
C930 B.n352 VSUBS 0.006127f
C931 B.n353 VSUBS 0.006127f
C932 B.n354 VSUBS 0.006127f
C933 B.n355 VSUBS 0.006127f
C934 B.n356 VSUBS 0.006127f
C935 B.n357 VSUBS 0.006127f
C936 B.n358 VSUBS 0.006127f
C937 B.n359 VSUBS 0.006127f
C938 B.n360 VSUBS 0.006127f
C939 B.n361 VSUBS 0.006127f
C940 B.n362 VSUBS 0.006127f
C941 B.n363 VSUBS 0.006127f
C942 B.n364 VSUBS 0.006127f
C943 B.n365 VSUBS 0.006127f
C944 B.n366 VSUBS 0.006127f
C945 B.n367 VSUBS 0.006127f
C946 B.n368 VSUBS 0.006127f
C947 B.n369 VSUBS 0.006127f
C948 B.n370 VSUBS 0.006127f
C949 B.n371 VSUBS 0.006127f
C950 B.n372 VSUBS 0.006127f
C951 B.n373 VSUBS 0.006127f
C952 B.n374 VSUBS 0.006127f
C953 B.n375 VSUBS 0.006127f
C954 B.n376 VSUBS 0.006127f
C955 B.n377 VSUBS 0.006127f
C956 B.n378 VSUBS 0.006127f
C957 B.n379 VSUBS 0.006127f
C958 B.n380 VSUBS 0.006127f
C959 B.n381 VSUBS 0.006127f
C960 B.n382 VSUBS 0.006127f
C961 B.n383 VSUBS 0.006127f
C962 B.n384 VSUBS 0.006127f
C963 B.n385 VSUBS 0.006127f
C964 B.n386 VSUBS 0.006127f
C965 B.n387 VSUBS 0.006127f
C966 B.n388 VSUBS 0.006127f
C967 B.n389 VSUBS 0.006127f
C968 B.n390 VSUBS 0.006127f
C969 B.n391 VSUBS 0.006127f
C970 B.n392 VSUBS 0.006127f
C971 B.n393 VSUBS 0.006127f
C972 B.n394 VSUBS 0.006127f
C973 B.n395 VSUBS 0.006127f
C974 B.n396 VSUBS 0.006127f
C975 B.n397 VSUBS 0.006127f
C976 B.n398 VSUBS 0.006127f
C977 B.n399 VSUBS 0.006127f
C978 B.n400 VSUBS 0.006127f
C979 B.n401 VSUBS 0.006127f
C980 B.n402 VSUBS 0.006127f
C981 B.n403 VSUBS 0.006127f
C982 B.n404 VSUBS 0.015308f
C983 B.n405 VSUBS 0.014245f
C984 B.n406 VSUBS 0.014936f
C985 B.n407 VSUBS 0.006127f
C986 B.n408 VSUBS 0.006127f
C987 B.n409 VSUBS 0.006127f
C988 B.n410 VSUBS 0.006127f
C989 B.n411 VSUBS 0.006127f
C990 B.n412 VSUBS 0.006127f
C991 B.n413 VSUBS 0.006127f
C992 B.n414 VSUBS 0.006127f
C993 B.n415 VSUBS 0.006127f
C994 B.n416 VSUBS 0.006127f
C995 B.n417 VSUBS 0.006127f
C996 B.n418 VSUBS 0.006127f
C997 B.n419 VSUBS 0.006127f
C998 B.n420 VSUBS 0.006127f
C999 B.n421 VSUBS 0.006127f
C1000 B.n422 VSUBS 0.006127f
C1001 B.n423 VSUBS 0.006127f
C1002 B.n424 VSUBS 0.006127f
C1003 B.n425 VSUBS 0.006127f
C1004 B.n426 VSUBS 0.006127f
C1005 B.n427 VSUBS 0.006127f
C1006 B.n428 VSUBS 0.006127f
C1007 B.n429 VSUBS 0.006127f
C1008 B.n430 VSUBS 0.006127f
C1009 B.n431 VSUBS 0.006127f
C1010 B.n432 VSUBS 0.006127f
C1011 B.n433 VSUBS 0.006127f
C1012 B.n434 VSUBS 0.006127f
C1013 B.n435 VSUBS 0.006127f
C1014 B.n436 VSUBS 0.006127f
C1015 B.n437 VSUBS 0.006127f
C1016 B.n438 VSUBS 0.006127f
C1017 B.n439 VSUBS 0.006127f
C1018 B.n440 VSUBS 0.006127f
C1019 B.n441 VSUBS 0.006127f
C1020 B.n442 VSUBS 0.006127f
C1021 B.n443 VSUBS 0.006127f
C1022 B.n444 VSUBS 0.006127f
C1023 B.n445 VSUBS 0.006127f
C1024 B.n446 VSUBS 0.006127f
C1025 B.n447 VSUBS 0.006127f
C1026 B.n448 VSUBS 0.006127f
C1027 B.n449 VSUBS 0.006127f
C1028 B.n450 VSUBS 0.006127f
C1029 B.n451 VSUBS 0.006127f
C1030 B.n452 VSUBS 0.006127f
C1031 B.n453 VSUBS 0.006127f
C1032 B.n454 VSUBS 0.006127f
C1033 B.n455 VSUBS 0.006127f
C1034 B.n456 VSUBS 0.006127f
C1035 B.n457 VSUBS 0.006127f
C1036 B.n458 VSUBS 0.006127f
C1037 B.n459 VSUBS 0.006127f
C1038 B.n460 VSUBS 0.006127f
C1039 B.n461 VSUBS 0.006127f
C1040 B.n462 VSUBS 0.006127f
C1041 B.n463 VSUBS 0.006127f
C1042 B.n464 VSUBS 0.006127f
C1043 B.n465 VSUBS 0.005766f
C1044 B.n466 VSUBS 0.006127f
C1045 B.n467 VSUBS 0.006127f
C1046 B.n468 VSUBS 0.003424f
C1047 B.n469 VSUBS 0.006127f
C1048 B.n470 VSUBS 0.006127f
C1049 B.n471 VSUBS 0.006127f
C1050 B.n472 VSUBS 0.006127f
C1051 B.n473 VSUBS 0.006127f
C1052 B.n474 VSUBS 0.006127f
C1053 B.n475 VSUBS 0.006127f
C1054 B.n476 VSUBS 0.006127f
C1055 B.n477 VSUBS 0.006127f
C1056 B.n478 VSUBS 0.006127f
C1057 B.n479 VSUBS 0.006127f
C1058 B.n480 VSUBS 0.006127f
C1059 B.n481 VSUBS 0.003424f
C1060 B.n482 VSUBS 0.014195f
C1061 B.n483 VSUBS 0.005766f
C1062 B.n484 VSUBS 0.006127f
C1063 B.n485 VSUBS 0.006127f
C1064 B.n486 VSUBS 0.006127f
C1065 B.n487 VSUBS 0.006127f
C1066 B.n488 VSUBS 0.006127f
C1067 B.n489 VSUBS 0.006127f
C1068 B.n490 VSUBS 0.006127f
C1069 B.n491 VSUBS 0.006127f
C1070 B.n492 VSUBS 0.006127f
C1071 B.n493 VSUBS 0.006127f
C1072 B.n494 VSUBS 0.006127f
C1073 B.n495 VSUBS 0.006127f
C1074 B.n496 VSUBS 0.006127f
C1075 B.n497 VSUBS 0.006127f
C1076 B.n498 VSUBS 0.006127f
C1077 B.n499 VSUBS 0.006127f
C1078 B.n500 VSUBS 0.006127f
C1079 B.n501 VSUBS 0.006127f
C1080 B.n502 VSUBS 0.006127f
C1081 B.n503 VSUBS 0.006127f
C1082 B.n504 VSUBS 0.006127f
C1083 B.n505 VSUBS 0.006127f
C1084 B.n506 VSUBS 0.006127f
C1085 B.n507 VSUBS 0.006127f
C1086 B.n508 VSUBS 0.006127f
C1087 B.n509 VSUBS 0.006127f
C1088 B.n510 VSUBS 0.006127f
C1089 B.n511 VSUBS 0.006127f
C1090 B.n512 VSUBS 0.006127f
C1091 B.n513 VSUBS 0.006127f
C1092 B.n514 VSUBS 0.006127f
C1093 B.n515 VSUBS 0.006127f
C1094 B.n516 VSUBS 0.006127f
C1095 B.n517 VSUBS 0.006127f
C1096 B.n518 VSUBS 0.006127f
C1097 B.n519 VSUBS 0.006127f
C1098 B.n520 VSUBS 0.006127f
C1099 B.n521 VSUBS 0.006127f
C1100 B.n522 VSUBS 0.006127f
C1101 B.n523 VSUBS 0.006127f
C1102 B.n524 VSUBS 0.006127f
C1103 B.n525 VSUBS 0.006127f
C1104 B.n526 VSUBS 0.006127f
C1105 B.n527 VSUBS 0.006127f
C1106 B.n528 VSUBS 0.006127f
C1107 B.n529 VSUBS 0.006127f
C1108 B.n530 VSUBS 0.006127f
C1109 B.n531 VSUBS 0.006127f
C1110 B.n532 VSUBS 0.006127f
C1111 B.n533 VSUBS 0.006127f
C1112 B.n534 VSUBS 0.006127f
C1113 B.n535 VSUBS 0.006127f
C1114 B.n536 VSUBS 0.006127f
C1115 B.n537 VSUBS 0.006127f
C1116 B.n538 VSUBS 0.006127f
C1117 B.n539 VSUBS 0.006127f
C1118 B.n540 VSUBS 0.006127f
C1119 B.n541 VSUBS 0.006127f
C1120 B.n542 VSUBS 0.006127f
C1121 B.n543 VSUBS 0.014936f
C1122 B.n544 VSUBS 0.014936f
C1123 B.n545 VSUBS 0.014616f
C1124 B.n546 VSUBS 0.006127f
C1125 B.n547 VSUBS 0.006127f
C1126 B.n548 VSUBS 0.006127f
C1127 B.n549 VSUBS 0.006127f
C1128 B.n550 VSUBS 0.006127f
C1129 B.n551 VSUBS 0.006127f
C1130 B.n552 VSUBS 0.006127f
C1131 B.n553 VSUBS 0.006127f
C1132 B.n554 VSUBS 0.006127f
C1133 B.n555 VSUBS 0.006127f
C1134 B.n556 VSUBS 0.006127f
C1135 B.n557 VSUBS 0.006127f
C1136 B.n558 VSUBS 0.006127f
C1137 B.n559 VSUBS 0.006127f
C1138 B.n560 VSUBS 0.006127f
C1139 B.n561 VSUBS 0.006127f
C1140 B.n562 VSUBS 0.006127f
C1141 B.n563 VSUBS 0.006127f
C1142 B.n564 VSUBS 0.006127f
C1143 B.n565 VSUBS 0.006127f
C1144 B.n566 VSUBS 0.006127f
C1145 B.n567 VSUBS 0.006127f
C1146 B.n568 VSUBS 0.006127f
C1147 B.n569 VSUBS 0.006127f
C1148 B.n570 VSUBS 0.006127f
C1149 B.n571 VSUBS 0.006127f
C1150 B.n572 VSUBS 0.006127f
C1151 B.n573 VSUBS 0.006127f
C1152 B.n574 VSUBS 0.006127f
C1153 B.n575 VSUBS 0.006127f
C1154 B.n576 VSUBS 0.006127f
C1155 B.n577 VSUBS 0.006127f
C1156 B.n578 VSUBS 0.006127f
C1157 B.n579 VSUBS 0.006127f
C1158 B.n580 VSUBS 0.006127f
C1159 B.n581 VSUBS 0.006127f
C1160 B.n582 VSUBS 0.006127f
C1161 B.n583 VSUBS 0.013873f
.ends

