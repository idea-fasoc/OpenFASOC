* NGSPICE file created from diff_pair_sample_0988.ext - technology: sky130A

.subckt diff_pair_sample_0988 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.31
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.31
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.31
X3 VDD1.t4 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.31
X4 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.31
X5 VDD2.t4 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.31
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.31
X7 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.31
X8 VTAIL.t0 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.31
X9 VTAIL.t9 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.31
X10 VTAIL.t5 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=1.97835 ps=12.32 w=11.99 l=3.31
X11 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.31
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=0 ps=0 w=11.99 l=3.31
X13 VDD1.t1 VP.t4 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.31
X14 VDD1.t0 VP.t5 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=4.6761 pd=24.76 as=1.97835 ps=12.32 w=11.99 l=3.31
X15 VDD2.t0 VN.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.97835 pd=12.32 as=4.6761 ps=24.76 w=11.99 l=3.31
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t5 120.597
R22 VP.n8 VP.t4 87.2993
R23 VP.n4 VP.t2 87.2993
R24 VP.n0 VP.t1 87.2993
R25 VP.n9 VP.t0 87.2993
R26 VP.n13 VP.t3 87.2993
R27 VP.n27 VP.n8 70.9831
R28 VP.n50 VP.n0 70.9831
R29 VP.n26 VP.n9 70.9831
R30 VP.n14 VP.n13 62.0573
R31 VP.n27 VP.n26 51.6357
R32 VP.n31 VP.n6 47.2923
R33 VP.n46 VP.n2 47.2923
R34 VP.n22 VP.n11 47.2923
R35 VP.n35 VP.n6 33.6945
R36 VP.n42 VP.n2 33.6945
R37 VP.n18 VP.n11 33.6945
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 19.0848
R51 VP.n48 VP.n0 19.0848
R52 VP.n24 VP.n9 19.0848
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 3.94731
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n270 VTAIL.n269 289.615
R81 VTAIL.n66 VTAIL.n65 289.615
R82 VTAIL.n204 VTAIL.n203 289.615
R83 VTAIL.n136 VTAIL.n135 289.615
R84 VTAIL.n229 VTAIL.n228 185
R85 VTAIL.n231 VTAIL.n230 185
R86 VTAIL.n224 VTAIL.n223 185
R87 VTAIL.n237 VTAIL.n236 185
R88 VTAIL.n239 VTAIL.n238 185
R89 VTAIL.n220 VTAIL.n219 185
R90 VTAIL.n245 VTAIL.n244 185
R91 VTAIL.n247 VTAIL.n246 185
R92 VTAIL.n216 VTAIL.n215 185
R93 VTAIL.n253 VTAIL.n252 185
R94 VTAIL.n255 VTAIL.n254 185
R95 VTAIL.n212 VTAIL.n211 185
R96 VTAIL.n261 VTAIL.n260 185
R97 VTAIL.n263 VTAIL.n262 185
R98 VTAIL.n208 VTAIL.n207 185
R99 VTAIL.n269 VTAIL.n268 185
R100 VTAIL.n25 VTAIL.n24 185
R101 VTAIL.n27 VTAIL.n26 185
R102 VTAIL.n20 VTAIL.n19 185
R103 VTAIL.n33 VTAIL.n32 185
R104 VTAIL.n35 VTAIL.n34 185
R105 VTAIL.n16 VTAIL.n15 185
R106 VTAIL.n41 VTAIL.n40 185
R107 VTAIL.n43 VTAIL.n42 185
R108 VTAIL.n12 VTAIL.n11 185
R109 VTAIL.n49 VTAIL.n48 185
R110 VTAIL.n51 VTAIL.n50 185
R111 VTAIL.n8 VTAIL.n7 185
R112 VTAIL.n57 VTAIL.n56 185
R113 VTAIL.n59 VTAIL.n58 185
R114 VTAIL.n4 VTAIL.n3 185
R115 VTAIL.n65 VTAIL.n64 185
R116 VTAIL.n203 VTAIL.n202 185
R117 VTAIL.n142 VTAIL.n141 185
R118 VTAIL.n197 VTAIL.n196 185
R119 VTAIL.n195 VTAIL.n194 185
R120 VTAIL.n146 VTAIL.n145 185
R121 VTAIL.n189 VTAIL.n188 185
R122 VTAIL.n187 VTAIL.n186 185
R123 VTAIL.n150 VTAIL.n149 185
R124 VTAIL.n181 VTAIL.n180 185
R125 VTAIL.n179 VTAIL.n178 185
R126 VTAIL.n154 VTAIL.n153 185
R127 VTAIL.n173 VTAIL.n172 185
R128 VTAIL.n171 VTAIL.n170 185
R129 VTAIL.n158 VTAIL.n157 185
R130 VTAIL.n165 VTAIL.n164 185
R131 VTAIL.n163 VTAIL.n162 185
R132 VTAIL.n135 VTAIL.n134 185
R133 VTAIL.n74 VTAIL.n73 185
R134 VTAIL.n129 VTAIL.n128 185
R135 VTAIL.n127 VTAIL.n126 185
R136 VTAIL.n78 VTAIL.n77 185
R137 VTAIL.n121 VTAIL.n120 185
R138 VTAIL.n119 VTAIL.n118 185
R139 VTAIL.n82 VTAIL.n81 185
R140 VTAIL.n113 VTAIL.n112 185
R141 VTAIL.n111 VTAIL.n110 185
R142 VTAIL.n86 VTAIL.n85 185
R143 VTAIL.n105 VTAIL.n104 185
R144 VTAIL.n103 VTAIL.n102 185
R145 VTAIL.n90 VTAIL.n89 185
R146 VTAIL.n97 VTAIL.n96 185
R147 VTAIL.n95 VTAIL.n94 185
R148 VTAIL.n93 VTAIL.t3 147.659
R149 VTAIL.n227 VTAIL.t11 147.659
R150 VTAIL.n23 VTAIL.t6 147.659
R151 VTAIL.n161 VTAIL.t7 147.659
R152 VTAIL.n230 VTAIL.n229 104.615
R153 VTAIL.n230 VTAIL.n223 104.615
R154 VTAIL.n237 VTAIL.n223 104.615
R155 VTAIL.n238 VTAIL.n237 104.615
R156 VTAIL.n238 VTAIL.n219 104.615
R157 VTAIL.n245 VTAIL.n219 104.615
R158 VTAIL.n246 VTAIL.n245 104.615
R159 VTAIL.n246 VTAIL.n215 104.615
R160 VTAIL.n253 VTAIL.n215 104.615
R161 VTAIL.n254 VTAIL.n253 104.615
R162 VTAIL.n254 VTAIL.n211 104.615
R163 VTAIL.n261 VTAIL.n211 104.615
R164 VTAIL.n262 VTAIL.n261 104.615
R165 VTAIL.n262 VTAIL.n207 104.615
R166 VTAIL.n269 VTAIL.n207 104.615
R167 VTAIL.n26 VTAIL.n25 104.615
R168 VTAIL.n26 VTAIL.n19 104.615
R169 VTAIL.n33 VTAIL.n19 104.615
R170 VTAIL.n34 VTAIL.n33 104.615
R171 VTAIL.n34 VTAIL.n15 104.615
R172 VTAIL.n41 VTAIL.n15 104.615
R173 VTAIL.n42 VTAIL.n41 104.615
R174 VTAIL.n42 VTAIL.n11 104.615
R175 VTAIL.n49 VTAIL.n11 104.615
R176 VTAIL.n50 VTAIL.n49 104.615
R177 VTAIL.n50 VTAIL.n7 104.615
R178 VTAIL.n57 VTAIL.n7 104.615
R179 VTAIL.n58 VTAIL.n57 104.615
R180 VTAIL.n58 VTAIL.n3 104.615
R181 VTAIL.n65 VTAIL.n3 104.615
R182 VTAIL.n203 VTAIL.n141 104.615
R183 VTAIL.n196 VTAIL.n141 104.615
R184 VTAIL.n196 VTAIL.n195 104.615
R185 VTAIL.n195 VTAIL.n145 104.615
R186 VTAIL.n188 VTAIL.n145 104.615
R187 VTAIL.n188 VTAIL.n187 104.615
R188 VTAIL.n187 VTAIL.n149 104.615
R189 VTAIL.n180 VTAIL.n149 104.615
R190 VTAIL.n180 VTAIL.n179 104.615
R191 VTAIL.n179 VTAIL.n153 104.615
R192 VTAIL.n172 VTAIL.n153 104.615
R193 VTAIL.n172 VTAIL.n171 104.615
R194 VTAIL.n171 VTAIL.n157 104.615
R195 VTAIL.n164 VTAIL.n157 104.615
R196 VTAIL.n164 VTAIL.n163 104.615
R197 VTAIL.n135 VTAIL.n73 104.615
R198 VTAIL.n128 VTAIL.n73 104.615
R199 VTAIL.n128 VTAIL.n127 104.615
R200 VTAIL.n127 VTAIL.n77 104.615
R201 VTAIL.n120 VTAIL.n77 104.615
R202 VTAIL.n120 VTAIL.n119 104.615
R203 VTAIL.n119 VTAIL.n81 104.615
R204 VTAIL.n112 VTAIL.n81 104.615
R205 VTAIL.n112 VTAIL.n111 104.615
R206 VTAIL.n111 VTAIL.n85 104.615
R207 VTAIL.n104 VTAIL.n85 104.615
R208 VTAIL.n104 VTAIL.n103 104.615
R209 VTAIL.n103 VTAIL.n89 104.615
R210 VTAIL.n96 VTAIL.n89 104.615
R211 VTAIL.n96 VTAIL.n95 104.615
R212 VTAIL.n229 VTAIL.t11 52.3082
R213 VTAIL.n25 VTAIL.t6 52.3082
R214 VTAIL.n163 VTAIL.t7 52.3082
R215 VTAIL.n95 VTAIL.t3 52.3082
R216 VTAIL.n139 VTAIL.n138 49.0664
R217 VTAIL.n71 VTAIL.n70 49.0664
R218 VTAIL.n1 VTAIL.n0 49.0662
R219 VTAIL.n69 VTAIL.n68 49.0662
R220 VTAIL.n271 VTAIL.n270 35.4823
R221 VTAIL.n67 VTAIL.n66 35.4823
R222 VTAIL.n205 VTAIL.n204 35.4823
R223 VTAIL.n137 VTAIL.n136 35.4823
R224 VTAIL.n71 VTAIL.n69 28.9789
R225 VTAIL.n271 VTAIL.n205 25.841
R226 VTAIL.n228 VTAIL.n227 15.6677
R227 VTAIL.n24 VTAIL.n23 15.6677
R228 VTAIL.n162 VTAIL.n161 15.6677
R229 VTAIL.n94 VTAIL.n93 15.6677
R230 VTAIL.n231 VTAIL.n226 12.8005
R231 VTAIL.n27 VTAIL.n22 12.8005
R232 VTAIL.n165 VTAIL.n160 12.8005
R233 VTAIL.n97 VTAIL.n92 12.8005
R234 VTAIL.n232 VTAIL.n224 12.0247
R235 VTAIL.n268 VTAIL.n206 12.0247
R236 VTAIL.n28 VTAIL.n20 12.0247
R237 VTAIL.n64 VTAIL.n2 12.0247
R238 VTAIL.n202 VTAIL.n140 12.0247
R239 VTAIL.n166 VTAIL.n158 12.0247
R240 VTAIL.n134 VTAIL.n72 12.0247
R241 VTAIL.n98 VTAIL.n90 12.0247
R242 VTAIL.n236 VTAIL.n235 11.249
R243 VTAIL.n267 VTAIL.n208 11.249
R244 VTAIL.n32 VTAIL.n31 11.249
R245 VTAIL.n63 VTAIL.n4 11.249
R246 VTAIL.n201 VTAIL.n142 11.249
R247 VTAIL.n170 VTAIL.n169 11.249
R248 VTAIL.n133 VTAIL.n74 11.249
R249 VTAIL.n102 VTAIL.n101 11.249
R250 VTAIL.n239 VTAIL.n222 10.4732
R251 VTAIL.n264 VTAIL.n263 10.4732
R252 VTAIL.n35 VTAIL.n18 10.4732
R253 VTAIL.n60 VTAIL.n59 10.4732
R254 VTAIL.n198 VTAIL.n197 10.4732
R255 VTAIL.n173 VTAIL.n156 10.4732
R256 VTAIL.n130 VTAIL.n129 10.4732
R257 VTAIL.n105 VTAIL.n88 10.4732
R258 VTAIL.n240 VTAIL.n220 9.69747
R259 VTAIL.n260 VTAIL.n210 9.69747
R260 VTAIL.n36 VTAIL.n16 9.69747
R261 VTAIL.n56 VTAIL.n6 9.69747
R262 VTAIL.n194 VTAIL.n144 9.69747
R263 VTAIL.n174 VTAIL.n154 9.69747
R264 VTAIL.n126 VTAIL.n76 9.69747
R265 VTAIL.n106 VTAIL.n86 9.69747
R266 VTAIL.n266 VTAIL.n206 9.45567
R267 VTAIL.n62 VTAIL.n2 9.45567
R268 VTAIL.n200 VTAIL.n140 9.45567
R269 VTAIL.n132 VTAIL.n72 9.45567
R270 VTAIL.n251 VTAIL.n250 9.3005
R271 VTAIL.n214 VTAIL.n213 9.3005
R272 VTAIL.n257 VTAIL.n256 9.3005
R273 VTAIL.n259 VTAIL.n258 9.3005
R274 VTAIL.n210 VTAIL.n209 9.3005
R275 VTAIL.n265 VTAIL.n264 9.3005
R276 VTAIL.n267 VTAIL.n266 9.3005
R277 VTAIL.n218 VTAIL.n217 9.3005
R278 VTAIL.n243 VTAIL.n242 9.3005
R279 VTAIL.n241 VTAIL.n240 9.3005
R280 VTAIL.n222 VTAIL.n221 9.3005
R281 VTAIL.n235 VTAIL.n234 9.3005
R282 VTAIL.n233 VTAIL.n232 9.3005
R283 VTAIL.n226 VTAIL.n225 9.3005
R284 VTAIL.n249 VTAIL.n248 9.3005
R285 VTAIL.n47 VTAIL.n46 9.3005
R286 VTAIL.n10 VTAIL.n9 9.3005
R287 VTAIL.n53 VTAIL.n52 9.3005
R288 VTAIL.n55 VTAIL.n54 9.3005
R289 VTAIL.n6 VTAIL.n5 9.3005
R290 VTAIL.n61 VTAIL.n60 9.3005
R291 VTAIL.n63 VTAIL.n62 9.3005
R292 VTAIL.n14 VTAIL.n13 9.3005
R293 VTAIL.n39 VTAIL.n38 9.3005
R294 VTAIL.n37 VTAIL.n36 9.3005
R295 VTAIL.n18 VTAIL.n17 9.3005
R296 VTAIL.n31 VTAIL.n30 9.3005
R297 VTAIL.n29 VTAIL.n28 9.3005
R298 VTAIL.n22 VTAIL.n21 9.3005
R299 VTAIL.n45 VTAIL.n44 9.3005
R300 VTAIL.n201 VTAIL.n200 9.3005
R301 VTAIL.n199 VTAIL.n198 9.3005
R302 VTAIL.n144 VTAIL.n143 9.3005
R303 VTAIL.n193 VTAIL.n192 9.3005
R304 VTAIL.n191 VTAIL.n190 9.3005
R305 VTAIL.n148 VTAIL.n147 9.3005
R306 VTAIL.n185 VTAIL.n184 9.3005
R307 VTAIL.n183 VTAIL.n182 9.3005
R308 VTAIL.n152 VTAIL.n151 9.3005
R309 VTAIL.n177 VTAIL.n176 9.3005
R310 VTAIL.n175 VTAIL.n174 9.3005
R311 VTAIL.n156 VTAIL.n155 9.3005
R312 VTAIL.n169 VTAIL.n168 9.3005
R313 VTAIL.n167 VTAIL.n166 9.3005
R314 VTAIL.n160 VTAIL.n159 9.3005
R315 VTAIL.n80 VTAIL.n79 9.3005
R316 VTAIL.n123 VTAIL.n122 9.3005
R317 VTAIL.n125 VTAIL.n124 9.3005
R318 VTAIL.n76 VTAIL.n75 9.3005
R319 VTAIL.n131 VTAIL.n130 9.3005
R320 VTAIL.n133 VTAIL.n132 9.3005
R321 VTAIL.n117 VTAIL.n116 9.3005
R322 VTAIL.n115 VTAIL.n114 9.3005
R323 VTAIL.n84 VTAIL.n83 9.3005
R324 VTAIL.n109 VTAIL.n108 9.3005
R325 VTAIL.n107 VTAIL.n106 9.3005
R326 VTAIL.n88 VTAIL.n87 9.3005
R327 VTAIL.n101 VTAIL.n100 9.3005
R328 VTAIL.n99 VTAIL.n98 9.3005
R329 VTAIL.n92 VTAIL.n91 9.3005
R330 VTAIL.n244 VTAIL.n243 8.92171
R331 VTAIL.n259 VTAIL.n212 8.92171
R332 VTAIL.n40 VTAIL.n39 8.92171
R333 VTAIL.n55 VTAIL.n8 8.92171
R334 VTAIL.n193 VTAIL.n146 8.92171
R335 VTAIL.n178 VTAIL.n177 8.92171
R336 VTAIL.n125 VTAIL.n78 8.92171
R337 VTAIL.n110 VTAIL.n109 8.92171
R338 VTAIL.n247 VTAIL.n218 8.14595
R339 VTAIL.n256 VTAIL.n255 8.14595
R340 VTAIL.n43 VTAIL.n14 8.14595
R341 VTAIL.n52 VTAIL.n51 8.14595
R342 VTAIL.n190 VTAIL.n189 8.14595
R343 VTAIL.n181 VTAIL.n152 8.14595
R344 VTAIL.n122 VTAIL.n121 8.14595
R345 VTAIL.n113 VTAIL.n84 8.14595
R346 VTAIL.n248 VTAIL.n216 7.3702
R347 VTAIL.n252 VTAIL.n214 7.3702
R348 VTAIL.n44 VTAIL.n12 7.3702
R349 VTAIL.n48 VTAIL.n10 7.3702
R350 VTAIL.n186 VTAIL.n148 7.3702
R351 VTAIL.n182 VTAIL.n150 7.3702
R352 VTAIL.n118 VTAIL.n80 7.3702
R353 VTAIL.n114 VTAIL.n82 7.3702
R354 VTAIL.n251 VTAIL.n216 6.59444
R355 VTAIL.n252 VTAIL.n251 6.59444
R356 VTAIL.n47 VTAIL.n12 6.59444
R357 VTAIL.n48 VTAIL.n47 6.59444
R358 VTAIL.n186 VTAIL.n185 6.59444
R359 VTAIL.n185 VTAIL.n150 6.59444
R360 VTAIL.n118 VTAIL.n117 6.59444
R361 VTAIL.n117 VTAIL.n82 6.59444
R362 VTAIL.n248 VTAIL.n247 5.81868
R363 VTAIL.n255 VTAIL.n214 5.81868
R364 VTAIL.n44 VTAIL.n43 5.81868
R365 VTAIL.n51 VTAIL.n10 5.81868
R366 VTAIL.n189 VTAIL.n148 5.81868
R367 VTAIL.n182 VTAIL.n181 5.81868
R368 VTAIL.n121 VTAIL.n80 5.81868
R369 VTAIL.n114 VTAIL.n113 5.81868
R370 VTAIL.n244 VTAIL.n218 5.04292
R371 VTAIL.n256 VTAIL.n212 5.04292
R372 VTAIL.n40 VTAIL.n14 5.04292
R373 VTAIL.n52 VTAIL.n8 5.04292
R374 VTAIL.n190 VTAIL.n146 5.04292
R375 VTAIL.n178 VTAIL.n152 5.04292
R376 VTAIL.n122 VTAIL.n78 5.04292
R377 VTAIL.n110 VTAIL.n84 5.04292
R378 VTAIL.n93 VTAIL.n91 4.38563
R379 VTAIL.n227 VTAIL.n225 4.38563
R380 VTAIL.n23 VTAIL.n21 4.38563
R381 VTAIL.n161 VTAIL.n159 4.38563
R382 VTAIL.n243 VTAIL.n220 4.26717
R383 VTAIL.n260 VTAIL.n259 4.26717
R384 VTAIL.n39 VTAIL.n16 4.26717
R385 VTAIL.n56 VTAIL.n55 4.26717
R386 VTAIL.n194 VTAIL.n193 4.26717
R387 VTAIL.n177 VTAIL.n154 4.26717
R388 VTAIL.n126 VTAIL.n125 4.26717
R389 VTAIL.n109 VTAIL.n86 4.26717
R390 VTAIL.n240 VTAIL.n239 3.49141
R391 VTAIL.n263 VTAIL.n210 3.49141
R392 VTAIL.n36 VTAIL.n35 3.49141
R393 VTAIL.n59 VTAIL.n6 3.49141
R394 VTAIL.n197 VTAIL.n144 3.49141
R395 VTAIL.n174 VTAIL.n173 3.49141
R396 VTAIL.n129 VTAIL.n76 3.49141
R397 VTAIL.n106 VTAIL.n105 3.49141
R398 VTAIL.n137 VTAIL.n71 3.13843
R399 VTAIL.n205 VTAIL.n139 3.13843
R400 VTAIL.n69 VTAIL.n67 3.13843
R401 VTAIL.n236 VTAIL.n222 2.71565
R402 VTAIL.n264 VTAIL.n208 2.71565
R403 VTAIL.n32 VTAIL.n18 2.71565
R404 VTAIL.n60 VTAIL.n4 2.71565
R405 VTAIL.n198 VTAIL.n142 2.71565
R406 VTAIL.n170 VTAIL.n156 2.71565
R407 VTAIL.n130 VTAIL.n74 2.71565
R408 VTAIL.n102 VTAIL.n88 2.71565
R409 VTAIL VTAIL.n271 2.29576
R410 VTAIL.n139 VTAIL.n137 2.03929
R411 VTAIL.n67 VTAIL.n1 2.03929
R412 VTAIL.n235 VTAIL.n224 1.93989
R413 VTAIL.n268 VTAIL.n267 1.93989
R414 VTAIL.n31 VTAIL.n20 1.93989
R415 VTAIL.n64 VTAIL.n63 1.93989
R416 VTAIL.n202 VTAIL.n201 1.93989
R417 VTAIL.n169 VTAIL.n158 1.93989
R418 VTAIL.n134 VTAIL.n133 1.93989
R419 VTAIL.n101 VTAIL.n90 1.93989
R420 VTAIL.n0 VTAIL.t2 1.65188
R421 VTAIL.n0 VTAIL.t0 1.65188
R422 VTAIL.n68 VTAIL.t8 1.65188
R423 VTAIL.n68 VTAIL.t9 1.65188
R424 VTAIL.n138 VTAIL.t4 1.65188
R425 VTAIL.n138 VTAIL.t5 1.65188
R426 VTAIL.n70 VTAIL.t10 1.65188
R427 VTAIL.n70 VTAIL.t1 1.65188
R428 VTAIL.n232 VTAIL.n231 1.16414
R429 VTAIL.n270 VTAIL.n206 1.16414
R430 VTAIL.n28 VTAIL.n27 1.16414
R431 VTAIL.n66 VTAIL.n2 1.16414
R432 VTAIL.n204 VTAIL.n140 1.16414
R433 VTAIL.n166 VTAIL.n165 1.16414
R434 VTAIL.n136 VTAIL.n72 1.16414
R435 VTAIL.n98 VTAIL.n97 1.16414
R436 VTAIL VTAIL.n1 0.843172
R437 VTAIL.n228 VTAIL.n226 0.388379
R438 VTAIL.n24 VTAIL.n22 0.388379
R439 VTAIL.n162 VTAIL.n160 0.388379
R440 VTAIL.n94 VTAIL.n92 0.388379
R441 VTAIL.n233 VTAIL.n225 0.155672
R442 VTAIL.n234 VTAIL.n233 0.155672
R443 VTAIL.n234 VTAIL.n221 0.155672
R444 VTAIL.n241 VTAIL.n221 0.155672
R445 VTAIL.n242 VTAIL.n241 0.155672
R446 VTAIL.n242 VTAIL.n217 0.155672
R447 VTAIL.n249 VTAIL.n217 0.155672
R448 VTAIL.n250 VTAIL.n249 0.155672
R449 VTAIL.n250 VTAIL.n213 0.155672
R450 VTAIL.n257 VTAIL.n213 0.155672
R451 VTAIL.n258 VTAIL.n257 0.155672
R452 VTAIL.n258 VTAIL.n209 0.155672
R453 VTAIL.n265 VTAIL.n209 0.155672
R454 VTAIL.n266 VTAIL.n265 0.155672
R455 VTAIL.n29 VTAIL.n21 0.155672
R456 VTAIL.n30 VTAIL.n29 0.155672
R457 VTAIL.n30 VTAIL.n17 0.155672
R458 VTAIL.n37 VTAIL.n17 0.155672
R459 VTAIL.n38 VTAIL.n37 0.155672
R460 VTAIL.n38 VTAIL.n13 0.155672
R461 VTAIL.n45 VTAIL.n13 0.155672
R462 VTAIL.n46 VTAIL.n45 0.155672
R463 VTAIL.n46 VTAIL.n9 0.155672
R464 VTAIL.n53 VTAIL.n9 0.155672
R465 VTAIL.n54 VTAIL.n53 0.155672
R466 VTAIL.n54 VTAIL.n5 0.155672
R467 VTAIL.n61 VTAIL.n5 0.155672
R468 VTAIL.n62 VTAIL.n61 0.155672
R469 VTAIL.n200 VTAIL.n199 0.155672
R470 VTAIL.n199 VTAIL.n143 0.155672
R471 VTAIL.n192 VTAIL.n143 0.155672
R472 VTAIL.n192 VTAIL.n191 0.155672
R473 VTAIL.n191 VTAIL.n147 0.155672
R474 VTAIL.n184 VTAIL.n147 0.155672
R475 VTAIL.n184 VTAIL.n183 0.155672
R476 VTAIL.n183 VTAIL.n151 0.155672
R477 VTAIL.n176 VTAIL.n151 0.155672
R478 VTAIL.n176 VTAIL.n175 0.155672
R479 VTAIL.n175 VTAIL.n155 0.155672
R480 VTAIL.n168 VTAIL.n155 0.155672
R481 VTAIL.n168 VTAIL.n167 0.155672
R482 VTAIL.n167 VTAIL.n159 0.155672
R483 VTAIL.n132 VTAIL.n131 0.155672
R484 VTAIL.n131 VTAIL.n75 0.155672
R485 VTAIL.n124 VTAIL.n75 0.155672
R486 VTAIL.n124 VTAIL.n123 0.155672
R487 VTAIL.n123 VTAIL.n79 0.155672
R488 VTAIL.n116 VTAIL.n79 0.155672
R489 VTAIL.n116 VTAIL.n115 0.155672
R490 VTAIL.n115 VTAIL.n83 0.155672
R491 VTAIL.n108 VTAIL.n83 0.155672
R492 VTAIL.n108 VTAIL.n107 0.155672
R493 VTAIL.n107 VTAIL.n87 0.155672
R494 VTAIL.n100 VTAIL.n87 0.155672
R495 VTAIL.n100 VTAIL.n99 0.155672
R496 VTAIL.n99 VTAIL.n91 0.155672
R497 VDD1.n64 VDD1.n63 289.615
R498 VDD1.n129 VDD1.n128 289.615
R499 VDD1.n63 VDD1.n62 185
R500 VDD1.n2 VDD1.n1 185
R501 VDD1.n57 VDD1.n56 185
R502 VDD1.n55 VDD1.n54 185
R503 VDD1.n6 VDD1.n5 185
R504 VDD1.n49 VDD1.n48 185
R505 VDD1.n47 VDD1.n46 185
R506 VDD1.n10 VDD1.n9 185
R507 VDD1.n41 VDD1.n40 185
R508 VDD1.n39 VDD1.n38 185
R509 VDD1.n14 VDD1.n13 185
R510 VDD1.n33 VDD1.n32 185
R511 VDD1.n31 VDD1.n30 185
R512 VDD1.n18 VDD1.n17 185
R513 VDD1.n25 VDD1.n24 185
R514 VDD1.n23 VDD1.n22 185
R515 VDD1.n88 VDD1.n87 185
R516 VDD1.n90 VDD1.n89 185
R517 VDD1.n83 VDD1.n82 185
R518 VDD1.n96 VDD1.n95 185
R519 VDD1.n98 VDD1.n97 185
R520 VDD1.n79 VDD1.n78 185
R521 VDD1.n104 VDD1.n103 185
R522 VDD1.n106 VDD1.n105 185
R523 VDD1.n75 VDD1.n74 185
R524 VDD1.n112 VDD1.n111 185
R525 VDD1.n114 VDD1.n113 185
R526 VDD1.n71 VDD1.n70 185
R527 VDD1.n120 VDD1.n119 185
R528 VDD1.n122 VDD1.n121 185
R529 VDD1.n67 VDD1.n66 185
R530 VDD1.n128 VDD1.n127 185
R531 VDD1.n21 VDD1.t0 147.659
R532 VDD1.n86 VDD1.t1 147.659
R533 VDD1.n63 VDD1.n1 104.615
R534 VDD1.n56 VDD1.n1 104.615
R535 VDD1.n56 VDD1.n55 104.615
R536 VDD1.n55 VDD1.n5 104.615
R537 VDD1.n48 VDD1.n5 104.615
R538 VDD1.n48 VDD1.n47 104.615
R539 VDD1.n47 VDD1.n9 104.615
R540 VDD1.n40 VDD1.n9 104.615
R541 VDD1.n40 VDD1.n39 104.615
R542 VDD1.n39 VDD1.n13 104.615
R543 VDD1.n32 VDD1.n13 104.615
R544 VDD1.n32 VDD1.n31 104.615
R545 VDD1.n31 VDD1.n17 104.615
R546 VDD1.n24 VDD1.n17 104.615
R547 VDD1.n24 VDD1.n23 104.615
R548 VDD1.n89 VDD1.n88 104.615
R549 VDD1.n89 VDD1.n82 104.615
R550 VDD1.n96 VDD1.n82 104.615
R551 VDD1.n97 VDD1.n96 104.615
R552 VDD1.n97 VDD1.n78 104.615
R553 VDD1.n104 VDD1.n78 104.615
R554 VDD1.n105 VDD1.n104 104.615
R555 VDD1.n105 VDD1.n74 104.615
R556 VDD1.n112 VDD1.n74 104.615
R557 VDD1.n113 VDD1.n112 104.615
R558 VDD1.n113 VDD1.n70 104.615
R559 VDD1.n120 VDD1.n70 104.615
R560 VDD1.n121 VDD1.n120 104.615
R561 VDD1.n121 VDD1.n66 104.615
R562 VDD1.n128 VDD1.n66 104.615
R563 VDD1.n131 VDD1.n130 66.4742
R564 VDD1.n133 VDD1.n132 65.7442
R565 VDD1 VDD1.n64 54.5727
R566 VDD1.n131 VDD1.n129 54.4592
R567 VDD1.n23 VDD1.t0 52.3082
R568 VDD1.n88 VDD1.t1 52.3082
R569 VDD1.n133 VDD1.n131 46.4018
R570 VDD1.n22 VDD1.n21 15.6677
R571 VDD1.n87 VDD1.n86 15.6677
R572 VDD1.n25 VDD1.n20 12.8005
R573 VDD1.n90 VDD1.n85 12.8005
R574 VDD1.n62 VDD1.n0 12.0247
R575 VDD1.n26 VDD1.n18 12.0247
R576 VDD1.n91 VDD1.n83 12.0247
R577 VDD1.n127 VDD1.n65 12.0247
R578 VDD1.n61 VDD1.n2 11.249
R579 VDD1.n30 VDD1.n29 11.249
R580 VDD1.n95 VDD1.n94 11.249
R581 VDD1.n126 VDD1.n67 11.249
R582 VDD1.n58 VDD1.n57 10.4732
R583 VDD1.n33 VDD1.n16 10.4732
R584 VDD1.n98 VDD1.n81 10.4732
R585 VDD1.n123 VDD1.n122 10.4732
R586 VDD1.n54 VDD1.n4 9.69747
R587 VDD1.n34 VDD1.n14 9.69747
R588 VDD1.n99 VDD1.n79 9.69747
R589 VDD1.n119 VDD1.n69 9.69747
R590 VDD1.n60 VDD1.n0 9.45567
R591 VDD1.n125 VDD1.n65 9.45567
R592 VDD1.n8 VDD1.n7 9.3005
R593 VDD1.n51 VDD1.n50 9.3005
R594 VDD1.n53 VDD1.n52 9.3005
R595 VDD1.n4 VDD1.n3 9.3005
R596 VDD1.n59 VDD1.n58 9.3005
R597 VDD1.n61 VDD1.n60 9.3005
R598 VDD1.n45 VDD1.n44 9.3005
R599 VDD1.n43 VDD1.n42 9.3005
R600 VDD1.n12 VDD1.n11 9.3005
R601 VDD1.n37 VDD1.n36 9.3005
R602 VDD1.n35 VDD1.n34 9.3005
R603 VDD1.n16 VDD1.n15 9.3005
R604 VDD1.n29 VDD1.n28 9.3005
R605 VDD1.n27 VDD1.n26 9.3005
R606 VDD1.n20 VDD1.n19 9.3005
R607 VDD1.n110 VDD1.n109 9.3005
R608 VDD1.n73 VDD1.n72 9.3005
R609 VDD1.n116 VDD1.n115 9.3005
R610 VDD1.n118 VDD1.n117 9.3005
R611 VDD1.n69 VDD1.n68 9.3005
R612 VDD1.n124 VDD1.n123 9.3005
R613 VDD1.n126 VDD1.n125 9.3005
R614 VDD1.n77 VDD1.n76 9.3005
R615 VDD1.n102 VDD1.n101 9.3005
R616 VDD1.n100 VDD1.n99 9.3005
R617 VDD1.n81 VDD1.n80 9.3005
R618 VDD1.n94 VDD1.n93 9.3005
R619 VDD1.n92 VDD1.n91 9.3005
R620 VDD1.n85 VDD1.n84 9.3005
R621 VDD1.n108 VDD1.n107 9.3005
R622 VDD1.n53 VDD1.n6 8.92171
R623 VDD1.n38 VDD1.n37 8.92171
R624 VDD1.n103 VDD1.n102 8.92171
R625 VDD1.n118 VDD1.n71 8.92171
R626 VDD1.n50 VDD1.n49 8.14595
R627 VDD1.n41 VDD1.n12 8.14595
R628 VDD1.n106 VDD1.n77 8.14595
R629 VDD1.n115 VDD1.n114 8.14595
R630 VDD1.n46 VDD1.n8 7.3702
R631 VDD1.n42 VDD1.n10 7.3702
R632 VDD1.n107 VDD1.n75 7.3702
R633 VDD1.n111 VDD1.n73 7.3702
R634 VDD1.n46 VDD1.n45 6.59444
R635 VDD1.n45 VDD1.n10 6.59444
R636 VDD1.n110 VDD1.n75 6.59444
R637 VDD1.n111 VDD1.n110 6.59444
R638 VDD1.n49 VDD1.n8 5.81868
R639 VDD1.n42 VDD1.n41 5.81868
R640 VDD1.n107 VDD1.n106 5.81868
R641 VDD1.n114 VDD1.n73 5.81868
R642 VDD1.n50 VDD1.n6 5.04292
R643 VDD1.n38 VDD1.n12 5.04292
R644 VDD1.n103 VDD1.n77 5.04292
R645 VDD1.n115 VDD1.n71 5.04292
R646 VDD1.n21 VDD1.n19 4.38563
R647 VDD1.n86 VDD1.n84 4.38563
R648 VDD1.n54 VDD1.n53 4.26717
R649 VDD1.n37 VDD1.n14 4.26717
R650 VDD1.n102 VDD1.n79 4.26717
R651 VDD1.n119 VDD1.n118 4.26717
R652 VDD1.n57 VDD1.n4 3.49141
R653 VDD1.n34 VDD1.n33 3.49141
R654 VDD1.n99 VDD1.n98 3.49141
R655 VDD1.n122 VDD1.n69 3.49141
R656 VDD1.n58 VDD1.n2 2.71565
R657 VDD1.n30 VDD1.n16 2.71565
R658 VDD1.n95 VDD1.n81 2.71565
R659 VDD1.n123 VDD1.n67 2.71565
R660 VDD1.n62 VDD1.n61 1.93989
R661 VDD1.n29 VDD1.n18 1.93989
R662 VDD1.n94 VDD1.n83 1.93989
R663 VDD1.n127 VDD1.n126 1.93989
R664 VDD1.n132 VDD1.t2 1.65188
R665 VDD1.n132 VDD1.t5 1.65188
R666 VDD1.n130 VDD1.t3 1.65188
R667 VDD1.n130 VDD1.t4 1.65188
R668 VDD1.n64 VDD1.n0 1.16414
R669 VDD1.n26 VDD1.n25 1.16414
R670 VDD1.n91 VDD1.n90 1.16414
R671 VDD1.n129 VDD1.n65 1.16414
R672 VDD1 VDD1.n133 0.726793
R673 VDD1.n22 VDD1.n20 0.388379
R674 VDD1.n87 VDD1.n85 0.388379
R675 VDD1.n60 VDD1.n59 0.155672
R676 VDD1.n59 VDD1.n3 0.155672
R677 VDD1.n52 VDD1.n3 0.155672
R678 VDD1.n52 VDD1.n51 0.155672
R679 VDD1.n51 VDD1.n7 0.155672
R680 VDD1.n44 VDD1.n7 0.155672
R681 VDD1.n44 VDD1.n43 0.155672
R682 VDD1.n43 VDD1.n11 0.155672
R683 VDD1.n36 VDD1.n11 0.155672
R684 VDD1.n36 VDD1.n35 0.155672
R685 VDD1.n35 VDD1.n15 0.155672
R686 VDD1.n28 VDD1.n15 0.155672
R687 VDD1.n28 VDD1.n27 0.155672
R688 VDD1.n27 VDD1.n19 0.155672
R689 VDD1.n92 VDD1.n84 0.155672
R690 VDD1.n93 VDD1.n92 0.155672
R691 VDD1.n93 VDD1.n80 0.155672
R692 VDD1.n100 VDD1.n80 0.155672
R693 VDD1.n101 VDD1.n100 0.155672
R694 VDD1.n101 VDD1.n76 0.155672
R695 VDD1.n108 VDD1.n76 0.155672
R696 VDD1.n109 VDD1.n108 0.155672
R697 VDD1.n109 VDD1.n72 0.155672
R698 VDD1.n116 VDD1.n72 0.155672
R699 VDD1.n117 VDD1.n116 0.155672
R700 VDD1.n117 VDD1.n68 0.155672
R701 VDD1.n124 VDD1.n68 0.155672
R702 VDD1.n125 VDD1.n124 0.155672
R703 B.n884 B.n883 585
R704 B.n885 B.n884 585
R705 B.n327 B.n141 585
R706 B.n326 B.n325 585
R707 B.n324 B.n323 585
R708 B.n322 B.n321 585
R709 B.n320 B.n319 585
R710 B.n318 B.n317 585
R711 B.n316 B.n315 585
R712 B.n314 B.n313 585
R713 B.n312 B.n311 585
R714 B.n310 B.n309 585
R715 B.n308 B.n307 585
R716 B.n306 B.n305 585
R717 B.n304 B.n303 585
R718 B.n302 B.n301 585
R719 B.n300 B.n299 585
R720 B.n298 B.n297 585
R721 B.n296 B.n295 585
R722 B.n294 B.n293 585
R723 B.n292 B.n291 585
R724 B.n290 B.n289 585
R725 B.n288 B.n287 585
R726 B.n286 B.n285 585
R727 B.n284 B.n283 585
R728 B.n282 B.n281 585
R729 B.n280 B.n279 585
R730 B.n278 B.n277 585
R731 B.n276 B.n275 585
R732 B.n274 B.n273 585
R733 B.n272 B.n271 585
R734 B.n270 B.n269 585
R735 B.n268 B.n267 585
R736 B.n266 B.n265 585
R737 B.n264 B.n263 585
R738 B.n262 B.n261 585
R739 B.n260 B.n259 585
R740 B.n258 B.n257 585
R741 B.n256 B.n255 585
R742 B.n254 B.n253 585
R743 B.n252 B.n251 585
R744 B.n250 B.n249 585
R745 B.n248 B.n247 585
R746 B.n245 B.n244 585
R747 B.n243 B.n242 585
R748 B.n241 B.n240 585
R749 B.n239 B.n238 585
R750 B.n237 B.n236 585
R751 B.n235 B.n234 585
R752 B.n233 B.n232 585
R753 B.n231 B.n230 585
R754 B.n229 B.n228 585
R755 B.n227 B.n226 585
R756 B.n225 B.n224 585
R757 B.n223 B.n222 585
R758 B.n221 B.n220 585
R759 B.n219 B.n218 585
R760 B.n217 B.n216 585
R761 B.n215 B.n214 585
R762 B.n213 B.n212 585
R763 B.n211 B.n210 585
R764 B.n209 B.n208 585
R765 B.n207 B.n206 585
R766 B.n205 B.n204 585
R767 B.n203 B.n202 585
R768 B.n201 B.n200 585
R769 B.n199 B.n198 585
R770 B.n197 B.n196 585
R771 B.n195 B.n194 585
R772 B.n193 B.n192 585
R773 B.n191 B.n190 585
R774 B.n189 B.n188 585
R775 B.n187 B.n186 585
R776 B.n185 B.n184 585
R777 B.n183 B.n182 585
R778 B.n181 B.n180 585
R779 B.n179 B.n178 585
R780 B.n177 B.n176 585
R781 B.n175 B.n174 585
R782 B.n173 B.n172 585
R783 B.n171 B.n170 585
R784 B.n169 B.n168 585
R785 B.n167 B.n166 585
R786 B.n165 B.n164 585
R787 B.n163 B.n162 585
R788 B.n161 B.n160 585
R789 B.n159 B.n158 585
R790 B.n157 B.n156 585
R791 B.n155 B.n154 585
R792 B.n153 B.n152 585
R793 B.n151 B.n150 585
R794 B.n149 B.n148 585
R795 B.n95 B.n94 585
R796 B.n888 B.n887 585
R797 B.n882 B.n142 585
R798 B.n142 B.n92 585
R799 B.n881 B.n91 585
R800 B.n892 B.n91 585
R801 B.n880 B.n90 585
R802 B.n893 B.n90 585
R803 B.n879 B.n89 585
R804 B.n894 B.n89 585
R805 B.n878 B.n877 585
R806 B.n877 B.n85 585
R807 B.n876 B.n84 585
R808 B.n900 B.n84 585
R809 B.n875 B.n83 585
R810 B.n901 B.n83 585
R811 B.n874 B.n82 585
R812 B.n902 B.n82 585
R813 B.n873 B.n872 585
R814 B.n872 B.n81 585
R815 B.n871 B.n77 585
R816 B.n908 B.n77 585
R817 B.n870 B.n76 585
R818 B.n909 B.n76 585
R819 B.n869 B.n75 585
R820 B.n910 B.n75 585
R821 B.n868 B.n867 585
R822 B.n867 B.n71 585
R823 B.n866 B.n70 585
R824 B.n916 B.n70 585
R825 B.n865 B.n69 585
R826 B.n917 B.n69 585
R827 B.n864 B.n68 585
R828 B.n918 B.n68 585
R829 B.n863 B.n862 585
R830 B.n862 B.n64 585
R831 B.n861 B.n63 585
R832 B.n924 B.n63 585
R833 B.n860 B.n62 585
R834 B.n925 B.n62 585
R835 B.n859 B.n61 585
R836 B.n926 B.n61 585
R837 B.n858 B.n857 585
R838 B.n857 B.n57 585
R839 B.n856 B.n56 585
R840 B.n932 B.n56 585
R841 B.n855 B.n55 585
R842 B.n933 B.n55 585
R843 B.n854 B.n54 585
R844 B.n934 B.n54 585
R845 B.n853 B.n852 585
R846 B.n852 B.n50 585
R847 B.n851 B.n49 585
R848 B.n940 B.n49 585
R849 B.n850 B.n48 585
R850 B.n941 B.n48 585
R851 B.n849 B.n47 585
R852 B.n942 B.n47 585
R853 B.n848 B.n847 585
R854 B.n847 B.n43 585
R855 B.n846 B.n42 585
R856 B.n948 B.n42 585
R857 B.n845 B.n41 585
R858 B.n949 B.n41 585
R859 B.n844 B.n40 585
R860 B.n950 B.n40 585
R861 B.n843 B.n842 585
R862 B.n842 B.n36 585
R863 B.n841 B.n35 585
R864 B.n956 B.n35 585
R865 B.n840 B.n34 585
R866 B.n957 B.n34 585
R867 B.n839 B.n33 585
R868 B.n958 B.n33 585
R869 B.n838 B.n837 585
R870 B.n837 B.n29 585
R871 B.n836 B.n28 585
R872 B.n964 B.n28 585
R873 B.n835 B.n27 585
R874 B.n965 B.n27 585
R875 B.n834 B.n26 585
R876 B.n966 B.n26 585
R877 B.n833 B.n832 585
R878 B.n832 B.n22 585
R879 B.n831 B.n21 585
R880 B.n972 B.n21 585
R881 B.n830 B.n20 585
R882 B.n973 B.n20 585
R883 B.n829 B.n19 585
R884 B.n974 B.n19 585
R885 B.n828 B.n827 585
R886 B.n827 B.n18 585
R887 B.n826 B.n14 585
R888 B.n980 B.n14 585
R889 B.n825 B.n13 585
R890 B.n981 B.n13 585
R891 B.n824 B.n12 585
R892 B.n982 B.n12 585
R893 B.n823 B.n822 585
R894 B.n822 B.n8 585
R895 B.n821 B.n7 585
R896 B.n988 B.n7 585
R897 B.n820 B.n6 585
R898 B.n989 B.n6 585
R899 B.n819 B.n5 585
R900 B.n990 B.n5 585
R901 B.n818 B.n817 585
R902 B.n817 B.n4 585
R903 B.n816 B.n328 585
R904 B.n816 B.n815 585
R905 B.n806 B.n329 585
R906 B.n330 B.n329 585
R907 B.n808 B.n807 585
R908 B.n809 B.n808 585
R909 B.n805 B.n335 585
R910 B.n335 B.n334 585
R911 B.n804 B.n803 585
R912 B.n803 B.n802 585
R913 B.n337 B.n336 585
R914 B.n795 B.n337 585
R915 B.n794 B.n793 585
R916 B.n796 B.n794 585
R917 B.n792 B.n342 585
R918 B.n342 B.n341 585
R919 B.n791 B.n790 585
R920 B.n790 B.n789 585
R921 B.n344 B.n343 585
R922 B.n345 B.n344 585
R923 B.n782 B.n781 585
R924 B.n783 B.n782 585
R925 B.n780 B.n350 585
R926 B.n350 B.n349 585
R927 B.n779 B.n778 585
R928 B.n778 B.n777 585
R929 B.n352 B.n351 585
R930 B.n353 B.n352 585
R931 B.n770 B.n769 585
R932 B.n771 B.n770 585
R933 B.n768 B.n358 585
R934 B.n358 B.n357 585
R935 B.n767 B.n766 585
R936 B.n766 B.n765 585
R937 B.n360 B.n359 585
R938 B.n361 B.n360 585
R939 B.n758 B.n757 585
R940 B.n759 B.n758 585
R941 B.n756 B.n366 585
R942 B.n366 B.n365 585
R943 B.n755 B.n754 585
R944 B.n754 B.n753 585
R945 B.n368 B.n367 585
R946 B.n369 B.n368 585
R947 B.n746 B.n745 585
R948 B.n747 B.n746 585
R949 B.n744 B.n374 585
R950 B.n374 B.n373 585
R951 B.n743 B.n742 585
R952 B.n742 B.n741 585
R953 B.n376 B.n375 585
R954 B.n377 B.n376 585
R955 B.n734 B.n733 585
R956 B.n735 B.n734 585
R957 B.n732 B.n381 585
R958 B.n385 B.n381 585
R959 B.n731 B.n730 585
R960 B.n730 B.n729 585
R961 B.n383 B.n382 585
R962 B.n384 B.n383 585
R963 B.n722 B.n721 585
R964 B.n723 B.n722 585
R965 B.n720 B.n390 585
R966 B.n390 B.n389 585
R967 B.n719 B.n718 585
R968 B.n718 B.n717 585
R969 B.n392 B.n391 585
R970 B.n393 B.n392 585
R971 B.n710 B.n709 585
R972 B.n711 B.n710 585
R973 B.n708 B.n398 585
R974 B.n398 B.n397 585
R975 B.n707 B.n706 585
R976 B.n706 B.n705 585
R977 B.n400 B.n399 585
R978 B.n401 B.n400 585
R979 B.n698 B.n697 585
R980 B.n699 B.n698 585
R981 B.n696 B.n406 585
R982 B.n406 B.n405 585
R983 B.n695 B.n694 585
R984 B.n694 B.n693 585
R985 B.n408 B.n407 585
R986 B.n686 B.n408 585
R987 B.n685 B.n684 585
R988 B.n687 B.n685 585
R989 B.n683 B.n413 585
R990 B.n413 B.n412 585
R991 B.n682 B.n681 585
R992 B.n681 B.n680 585
R993 B.n415 B.n414 585
R994 B.n416 B.n415 585
R995 B.n673 B.n672 585
R996 B.n674 B.n673 585
R997 B.n671 B.n421 585
R998 B.n421 B.n420 585
R999 B.n670 B.n669 585
R1000 B.n669 B.n668 585
R1001 B.n423 B.n422 585
R1002 B.n424 B.n423 585
R1003 B.n664 B.n663 585
R1004 B.n427 B.n426 585
R1005 B.n660 B.n659 585
R1006 B.n661 B.n660 585
R1007 B.n658 B.n473 585
R1008 B.n657 B.n656 585
R1009 B.n655 B.n654 585
R1010 B.n653 B.n652 585
R1011 B.n651 B.n650 585
R1012 B.n649 B.n648 585
R1013 B.n647 B.n646 585
R1014 B.n645 B.n644 585
R1015 B.n643 B.n642 585
R1016 B.n641 B.n640 585
R1017 B.n639 B.n638 585
R1018 B.n637 B.n636 585
R1019 B.n635 B.n634 585
R1020 B.n633 B.n632 585
R1021 B.n631 B.n630 585
R1022 B.n629 B.n628 585
R1023 B.n627 B.n626 585
R1024 B.n625 B.n624 585
R1025 B.n623 B.n622 585
R1026 B.n621 B.n620 585
R1027 B.n619 B.n618 585
R1028 B.n617 B.n616 585
R1029 B.n615 B.n614 585
R1030 B.n613 B.n612 585
R1031 B.n611 B.n610 585
R1032 B.n609 B.n608 585
R1033 B.n607 B.n606 585
R1034 B.n605 B.n604 585
R1035 B.n603 B.n602 585
R1036 B.n601 B.n600 585
R1037 B.n599 B.n598 585
R1038 B.n597 B.n596 585
R1039 B.n595 B.n594 585
R1040 B.n593 B.n592 585
R1041 B.n591 B.n590 585
R1042 B.n589 B.n588 585
R1043 B.n587 B.n586 585
R1044 B.n585 B.n584 585
R1045 B.n583 B.n582 585
R1046 B.n580 B.n579 585
R1047 B.n578 B.n577 585
R1048 B.n576 B.n575 585
R1049 B.n574 B.n573 585
R1050 B.n572 B.n571 585
R1051 B.n570 B.n569 585
R1052 B.n568 B.n567 585
R1053 B.n566 B.n565 585
R1054 B.n564 B.n563 585
R1055 B.n562 B.n561 585
R1056 B.n560 B.n559 585
R1057 B.n558 B.n557 585
R1058 B.n556 B.n555 585
R1059 B.n554 B.n553 585
R1060 B.n552 B.n551 585
R1061 B.n550 B.n549 585
R1062 B.n548 B.n547 585
R1063 B.n546 B.n545 585
R1064 B.n544 B.n543 585
R1065 B.n542 B.n541 585
R1066 B.n540 B.n539 585
R1067 B.n538 B.n537 585
R1068 B.n536 B.n535 585
R1069 B.n534 B.n533 585
R1070 B.n532 B.n531 585
R1071 B.n530 B.n529 585
R1072 B.n528 B.n527 585
R1073 B.n526 B.n525 585
R1074 B.n524 B.n523 585
R1075 B.n522 B.n521 585
R1076 B.n520 B.n519 585
R1077 B.n518 B.n517 585
R1078 B.n516 B.n515 585
R1079 B.n514 B.n513 585
R1080 B.n512 B.n511 585
R1081 B.n510 B.n509 585
R1082 B.n508 B.n507 585
R1083 B.n506 B.n505 585
R1084 B.n504 B.n503 585
R1085 B.n502 B.n501 585
R1086 B.n500 B.n499 585
R1087 B.n498 B.n497 585
R1088 B.n496 B.n495 585
R1089 B.n494 B.n493 585
R1090 B.n492 B.n491 585
R1091 B.n490 B.n489 585
R1092 B.n488 B.n487 585
R1093 B.n486 B.n485 585
R1094 B.n484 B.n483 585
R1095 B.n482 B.n481 585
R1096 B.n480 B.n479 585
R1097 B.n665 B.n425 585
R1098 B.n425 B.n424 585
R1099 B.n667 B.n666 585
R1100 B.n668 B.n667 585
R1101 B.n419 B.n418 585
R1102 B.n420 B.n419 585
R1103 B.n676 B.n675 585
R1104 B.n675 B.n674 585
R1105 B.n677 B.n417 585
R1106 B.n417 B.n416 585
R1107 B.n679 B.n678 585
R1108 B.n680 B.n679 585
R1109 B.n411 B.n410 585
R1110 B.n412 B.n411 585
R1111 B.n689 B.n688 585
R1112 B.n688 B.n687 585
R1113 B.n690 B.n409 585
R1114 B.n686 B.n409 585
R1115 B.n692 B.n691 585
R1116 B.n693 B.n692 585
R1117 B.n404 B.n403 585
R1118 B.n405 B.n404 585
R1119 B.n701 B.n700 585
R1120 B.n700 B.n699 585
R1121 B.n702 B.n402 585
R1122 B.n402 B.n401 585
R1123 B.n704 B.n703 585
R1124 B.n705 B.n704 585
R1125 B.n396 B.n395 585
R1126 B.n397 B.n396 585
R1127 B.n713 B.n712 585
R1128 B.n712 B.n711 585
R1129 B.n714 B.n394 585
R1130 B.n394 B.n393 585
R1131 B.n716 B.n715 585
R1132 B.n717 B.n716 585
R1133 B.n388 B.n387 585
R1134 B.n389 B.n388 585
R1135 B.n725 B.n724 585
R1136 B.n724 B.n723 585
R1137 B.n726 B.n386 585
R1138 B.n386 B.n384 585
R1139 B.n728 B.n727 585
R1140 B.n729 B.n728 585
R1141 B.n380 B.n379 585
R1142 B.n385 B.n380 585
R1143 B.n737 B.n736 585
R1144 B.n736 B.n735 585
R1145 B.n738 B.n378 585
R1146 B.n378 B.n377 585
R1147 B.n740 B.n739 585
R1148 B.n741 B.n740 585
R1149 B.n372 B.n371 585
R1150 B.n373 B.n372 585
R1151 B.n749 B.n748 585
R1152 B.n748 B.n747 585
R1153 B.n750 B.n370 585
R1154 B.n370 B.n369 585
R1155 B.n752 B.n751 585
R1156 B.n753 B.n752 585
R1157 B.n364 B.n363 585
R1158 B.n365 B.n364 585
R1159 B.n761 B.n760 585
R1160 B.n760 B.n759 585
R1161 B.n762 B.n362 585
R1162 B.n362 B.n361 585
R1163 B.n764 B.n763 585
R1164 B.n765 B.n764 585
R1165 B.n356 B.n355 585
R1166 B.n357 B.n356 585
R1167 B.n773 B.n772 585
R1168 B.n772 B.n771 585
R1169 B.n774 B.n354 585
R1170 B.n354 B.n353 585
R1171 B.n776 B.n775 585
R1172 B.n777 B.n776 585
R1173 B.n348 B.n347 585
R1174 B.n349 B.n348 585
R1175 B.n785 B.n784 585
R1176 B.n784 B.n783 585
R1177 B.n786 B.n346 585
R1178 B.n346 B.n345 585
R1179 B.n788 B.n787 585
R1180 B.n789 B.n788 585
R1181 B.n340 B.n339 585
R1182 B.n341 B.n340 585
R1183 B.n798 B.n797 585
R1184 B.n797 B.n796 585
R1185 B.n799 B.n338 585
R1186 B.n795 B.n338 585
R1187 B.n801 B.n800 585
R1188 B.n802 B.n801 585
R1189 B.n333 B.n332 585
R1190 B.n334 B.n333 585
R1191 B.n811 B.n810 585
R1192 B.n810 B.n809 585
R1193 B.n812 B.n331 585
R1194 B.n331 B.n330 585
R1195 B.n814 B.n813 585
R1196 B.n815 B.n814 585
R1197 B.n2 B.n0 585
R1198 B.n4 B.n2 585
R1199 B.n3 B.n1 585
R1200 B.n989 B.n3 585
R1201 B.n987 B.n986 585
R1202 B.n988 B.n987 585
R1203 B.n985 B.n9 585
R1204 B.n9 B.n8 585
R1205 B.n984 B.n983 585
R1206 B.n983 B.n982 585
R1207 B.n11 B.n10 585
R1208 B.n981 B.n11 585
R1209 B.n979 B.n978 585
R1210 B.n980 B.n979 585
R1211 B.n977 B.n15 585
R1212 B.n18 B.n15 585
R1213 B.n976 B.n975 585
R1214 B.n975 B.n974 585
R1215 B.n17 B.n16 585
R1216 B.n973 B.n17 585
R1217 B.n971 B.n970 585
R1218 B.n972 B.n971 585
R1219 B.n969 B.n23 585
R1220 B.n23 B.n22 585
R1221 B.n968 B.n967 585
R1222 B.n967 B.n966 585
R1223 B.n25 B.n24 585
R1224 B.n965 B.n25 585
R1225 B.n963 B.n962 585
R1226 B.n964 B.n963 585
R1227 B.n961 B.n30 585
R1228 B.n30 B.n29 585
R1229 B.n960 B.n959 585
R1230 B.n959 B.n958 585
R1231 B.n32 B.n31 585
R1232 B.n957 B.n32 585
R1233 B.n955 B.n954 585
R1234 B.n956 B.n955 585
R1235 B.n953 B.n37 585
R1236 B.n37 B.n36 585
R1237 B.n952 B.n951 585
R1238 B.n951 B.n950 585
R1239 B.n39 B.n38 585
R1240 B.n949 B.n39 585
R1241 B.n947 B.n946 585
R1242 B.n948 B.n947 585
R1243 B.n945 B.n44 585
R1244 B.n44 B.n43 585
R1245 B.n944 B.n943 585
R1246 B.n943 B.n942 585
R1247 B.n46 B.n45 585
R1248 B.n941 B.n46 585
R1249 B.n939 B.n938 585
R1250 B.n940 B.n939 585
R1251 B.n937 B.n51 585
R1252 B.n51 B.n50 585
R1253 B.n936 B.n935 585
R1254 B.n935 B.n934 585
R1255 B.n53 B.n52 585
R1256 B.n933 B.n53 585
R1257 B.n931 B.n930 585
R1258 B.n932 B.n931 585
R1259 B.n929 B.n58 585
R1260 B.n58 B.n57 585
R1261 B.n928 B.n927 585
R1262 B.n927 B.n926 585
R1263 B.n60 B.n59 585
R1264 B.n925 B.n60 585
R1265 B.n923 B.n922 585
R1266 B.n924 B.n923 585
R1267 B.n921 B.n65 585
R1268 B.n65 B.n64 585
R1269 B.n920 B.n919 585
R1270 B.n919 B.n918 585
R1271 B.n67 B.n66 585
R1272 B.n917 B.n67 585
R1273 B.n915 B.n914 585
R1274 B.n916 B.n915 585
R1275 B.n913 B.n72 585
R1276 B.n72 B.n71 585
R1277 B.n912 B.n911 585
R1278 B.n911 B.n910 585
R1279 B.n74 B.n73 585
R1280 B.n909 B.n74 585
R1281 B.n907 B.n906 585
R1282 B.n908 B.n907 585
R1283 B.n905 B.n78 585
R1284 B.n81 B.n78 585
R1285 B.n904 B.n903 585
R1286 B.n903 B.n902 585
R1287 B.n80 B.n79 585
R1288 B.n901 B.n80 585
R1289 B.n899 B.n898 585
R1290 B.n900 B.n899 585
R1291 B.n897 B.n86 585
R1292 B.n86 B.n85 585
R1293 B.n896 B.n895 585
R1294 B.n895 B.n894 585
R1295 B.n88 B.n87 585
R1296 B.n893 B.n88 585
R1297 B.n891 B.n890 585
R1298 B.n892 B.n891 585
R1299 B.n889 B.n93 585
R1300 B.n93 B.n92 585
R1301 B.n992 B.n991 585
R1302 B.n991 B.n990 585
R1303 B.n663 B.n425 468.476
R1304 B.n887 B.n93 468.476
R1305 B.n479 B.n423 468.476
R1306 B.n884 B.n142 468.476
R1307 B.n476 B.t19 352.409
R1308 B.n143 B.t15 352.409
R1309 B.n474 B.t9 352.409
R1310 B.n145 B.t12 352.409
R1311 B.n476 B.t17 296.214
R1312 B.n474 B.t6 296.214
R1313 B.n145 B.t10 296.214
R1314 B.n143 B.t14 296.214
R1315 B.n477 B.t18 281.815
R1316 B.n144 B.t16 281.815
R1317 B.n475 B.t8 281.815
R1318 B.n146 B.t13 281.815
R1319 B.n885 B.n140 256.663
R1320 B.n885 B.n139 256.663
R1321 B.n885 B.n138 256.663
R1322 B.n885 B.n137 256.663
R1323 B.n885 B.n136 256.663
R1324 B.n885 B.n135 256.663
R1325 B.n885 B.n134 256.663
R1326 B.n885 B.n133 256.663
R1327 B.n885 B.n132 256.663
R1328 B.n885 B.n131 256.663
R1329 B.n885 B.n130 256.663
R1330 B.n885 B.n129 256.663
R1331 B.n885 B.n128 256.663
R1332 B.n885 B.n127 256.663
R1333 B.n885 B.n126 256.663
R1334 B.n885 B.n125 256.663
R1335 B.n885 B.n124 256.663
R1336 B.n885 B.n123 256.663
R1337 B.n885 B.n122 256.663
R1338 B.n885 B.n121 256.663
R1339 B.n885 B.n120 256.663
R1340 B.n885 B.n119 256.663
R1341 B.n885 B.n118 256.663
R1342 B.n885 B.n117 256.663
R1343 B.n885 B.n116 256.663
R1344 B.n885 B.n115 256.663
R1345 B.n885 B.n114 256.663
R1346 B.n885 B.n113 256.663
R1347 B.n885 B.n112 256.663
R1348 B.n885 B.n111 256.663
R1349 B.n885 B.n110 256.663
R1350 B.n885 B.n109 256.663
R1351 B.n885 B.n108 256.663
R1352 B.n885 B.n107 256.663
R1353 B.n885 B.n106 256.663
R1354 B.n885 B.n105 256.663
R1355 B.n885 B.n104 256.663
R1356 B.n885 B.n103 256.663
R1357 B.n885 B.n102 256.663
R1358 B.n885 B.n101 256.663
R1359 B.n885 B.n100 256.663
R1360 B.n885 B.n99 256.663
R1361 B.n885 B.n98 256.663
R1362 B.n885 B.n97 256.663
R1363 B.n885 B.n96 256.663
R1364 B.n886 B.n885 256.663
R1365 B.n662 B.n661 256.663
R1366 B.n661 B.n428 256.663
R1367 B.n661 B.n429 256.663
R1368 B.n661 B.n430 256.663
R1369 B.n661 B.n431 256.663
R1370 B.n661 B.n432 256.663
R1371 B.n661 B.n433 256.663
R1372 B.n661 B.n434 256.663
R1373 B.n661 B.n435 256.663
R1374 B.n661 B.n436 256.663
R1375 B.n661 B.n437 256.663
R1376 B.n661 B.n438 256.663
R1377 B.n661 B.n439 256.663
R1378 B.n661 B.n440 256.663
R1379 B.n661 B.n441 256.663
R1380 B.n661 B.n442 256.663
R1381 B.n661 B.n443 256.663
R1382 B.n661 B.n444 256.663
R1383 B.n661 B.n445 256.663
R1384 B.n661 B.n446 256.663
R1385 B.n661 B.n447 256.663
R1386 B.n661 B.n448 256.663
R1387 B.n661 B.n449 256.663
R1388 B.n661 B.n450 256.663
R1389 B.n661 B.n451 256.663
R1390 B.n661 B.n452 256.663
R1391 B.n661 B.n453 256.663
R1392 B.n661 B.n454 256.663
R1393 B.n661 B.n455 256.663
R1394 B.n661 B.n456 256.663
R1395 B.n661 B.n457 256.663
R1396 B.n661 B.n458 256.663
R1397 B.n661 B.n459 256.663
R1398 B.n661 B.n460 256.663
R1399 B.n661 B.n461 256.663
R1400 B.n661 B.n462 256.663
R1401 B.n661 B.n463 256.663
R1402 B.n661 B.n464 256.663
R1403 B.n661 B.n465 256.663
R1404 B.n661 B.n466 256.663
R1405 B.n661 B.n467 256.663
R1406 B.n661 B.n468 256.663
R1407 B.n661 B.n469 256.663
R1408 B.n661 B.n470 256.663
R1409 B.n661 B.n471 256.663
R1410 B.n661 B.n472 256.663
R1411 B.n667 B.n425 163.367
R1412 B.n667 B.n419 163.367
R1413 B.n675 B.n419 163.367
R1414 B.n675 B.n417 163.367
R1415 B.n679 B.n417 163.367
R1416 B.n679 B.n411 163.367
R1417 B.n688 B.n411 163.367
R1418 B.n688 B.n409 163.367
R1419 B.n692 B.n409 163.367
R1420 B.n692 B.n404 163.367
R1421 B.n700 B.n404 163.367
R1422 B.n700 B.n402 163.367
R1423 B.n704 B.n402 163.367
R1424 B.n704 B.n396 163.367
R1425 B.n712 B.n396 163.367
R1426 B.n712 B.n394 163.367
R1427 B.n716 B.n394 163.367
R1428 B.n716 B.n388 163.367
R1429 B.n724 B.n388 163.367
R1430 B.n724 B.n386 163.367
R1431 B.n728 B.n386 163.367
R1432 B.n728 B.n380 163.367
R1433 B.n736 B.n380 163.367
R1434 B.n736 B.n378 163.367
R1435 B.n740 B.n378 163.367
R1436 B.n740 B.n372 163.367
R1437 B.n748 B.n372 163.367
R1438 B.n748 B.n370 163.367
R1439 B.n752 B.n370 163.367
R1440 B.n752 B.n364 163.367
R1441 B.n760 B.n364 163.367
R1442 B.n760 B.n362 163.367
R1443 B.n764 B.n362 163.367
R1444 B.n764 B.n356 163.367
R1445 B.n772 B.n356 163.367
R1446 B.n772 B.n354 163.367
R1447 B.n776 B.n354 163.367
R1448 B.n776 B.n348 163.367
R1449 B.n784 B.n348 163.367
R1450 B.n784 B.n346 163.367
R1451 B.n788 B.n346 163.367
R1452 B.n788 B.n340 163.367
R1453 B.n797 B.n340 163.367
R1454 B.n797 B.n338 163.367
R1455 B.n801 B.n338 163.367
R1456 B.n801 B.n333 163.367
R1457 B.n810 B.n333 163.367
R1458 B.n810 B.n331 163.367
R1459 B.n814 B.n331 163.367
R1460 B.n814 B.n2 163.367
R1461 B.n991 B.n2 163.367
R1462 B.n991 B.n3 163.367
R1463 B.n987 B.n3 163.367
R1464 B.n987 B.n9 163.367
R1465 B.n983 B.n9 163.367
R1466 B.n983 B.n11 163.367
R1467 B.n979 B.n11 163.367
R1468 B.n979 B.n15 163.367
R1469 B.n975 B.n15 163.367
R1470 B.n975 B.n17 163.367
R1471 B.n971 B.n17 163.367
R1472 B.n971 B.n23 163.367
R1473 B.n967 B.n23 163.367
R1474 B.n967 B.n25 163.367
R1475 B.n963 B.n25 163.367
R1476 B.n963 B.n30 163.367
R1477 B.n959 B.n30 163.367
R1478 B.n959 B.n32 163.367
R1479 B.n955 B.n32 163.367
R1480 B.n955 B.n37 163.367
R1481 B.n951 B.n37 163.367
R1482 B.n951 B.n39 163.367
R1483 B.n947 B.n39 163.367
R1484 B.n947 B.n44 163.367
R1485 B.n943 B.n44 163.367
R1486 B.n943 B.n46 163.367
R1487 B.n939 B.n46 163.367
R1488 B.n939 B.n51 163.367
R1489 B.n935 B.n51 163.367
R1490 B.n935 B.n53 163.367
R1491 B.n931 B.n53 163.367
R1492 B.n931 B.n58 163.367
R1493 B.n927 B.n58 163.367
R1494 B.n927 B.n60 163.367
R1495 B.n923 B.n60 163.367
R1496 B.n923 B.n65 163.367
R1497 B.n919 B.n65 163.367
R1498 B.n919 B.n67 163.367
R1499 B.n915 B.n67 163.367
R1500 B.n915 B.n72 163.367
R1501 B.n911 B.n72 163.367
R1502 B.n911 B.n74 163.367
R1503 B.n907 B.n74 163.367
R1504 B.n907 B.n78 163.367
R1505 B.n903 B.n78 163.367
R1506 B.n903 B.n80 163.367
R1507 B.n899 B.n80 163.367
R1508 B.n899 B.n86 163.367
R1509 B.n895 B.n86 163.367
R1510 B.n895 B.n88 163.367
R1511 B.n891 B.n88 163.367
R1512 B.n891 B.n93 163.367
R1513 B.n660 B.n427 163.367
R1514 B.n660 B.n473 163.367
R1515 B.n656 B.n655 163.367
R1516 B.n652 B.n651 163.367
R1517 B.n648 B.n647 163.367
R1518 B.n644 B.n643 163.367
R1519 B.n640 B.n639 163.367
R1520 B.n636 B.n635 163.367
R1521 B.n632 B.n631 163.367
R1522 B.n628 B.n627 163.367
R1523 B.n624 B.n623 163.367
R1524 B.n620 B.n619 163.367
R1525 B.n616 B.n615 163.367
R1526 B.n612 B.n611 163.367
R1527 B.n608 B.n607 163.367
R1528 B.n604 B.n603 163.367
R1529 B.n600 B.n599 163.367
R1530 B.n596 B.n595 163.367
R1531 B.n592 B.n591 163.367
R1532 B.n588 B.n587 163.367
R1533 B.n584 B.n583 163.367
R1534 B.n579 B.n578 163.367
R1535 B.n575 B.n574 163.367
R1536 B.n571 B.n570 163.367
R1537 B.n567 B.n566 163.367
R1538 B.n563 B.n562 163.367
R1539 B.n559 B.n558 163.367
R1540 B.n555 B.n554 163.367
R1541 B.n551 B.n550 163.367
R1542 B.n547 B.n546 163.367
R1543 B.n543 B.n542 163.367
R1544 B.n539 B.n538 163.367
R1545 B.n535 B.n534 163.367
R1546 B.n531 B.n530 163.367
R1547 B.n527 B.n526 163.367
R1548 B.n523 B.n522 163.367
R1549 B.n519 B.n518 163.367
R1550 B.n515 B.n514 163.367
R1551 B.n511 B.n510 163.367
R1552 B.n507 B.n506 163.367
R1553 B.n503 B.n502 163.367
R1554 B.n499 B.n498 163.367
R1555 B.n495 B.n494 163.367
R1556 B.n491 B.n490 163.367
R1557 B.n487 B.n486 163.367
R1558 B.n483 B.n482 163.367
R1559 B.n669 B.n423 163.367
R1560 B.n669 B.n421 163.367
R1561 B.n673 B.n421 163.367
R1562 B.n673 B.n415 163.367
R1563 B.n681 B.n415 163.367
R1564 B.n681 B.n413 163.367
R1565 B.n685 B.n413 163.367
R1566 B.n685 B.n408 163.367
R1567 B.n694 B.n408 163.367
R1568 B.n694 B.n406 163.367
R1569 B.n698 B.n406 163.367
R1570 B.n698 B.n400 163.367
R1571 B.n706 B.n400 163.367
R1572 B.n706 B.n398 163.367
R1573 B.n710 B.n398 163.367
R1574 B.n710 B.n392 163.367
R1575 B.n718 B.n392 163.367
R1576 B.n718 B.n390 163.367
R1577 B.n722 B.n390 163.367
R1578 B.n722 B.n383 163.367
R1579 B.n730 B.n383 163.367
R1580 B.n730 B.n381 163.367
R1581 B.n734 B.n381 163.367
R1582 B.n734 B.n376 163.367
R1583 B.n742 B.n376 163.367
R1584 B.n742 B.n374 163.367
R1585 B.n746 B.n374 163.367
R1586 B.n746 B.n368 163.367
R1587 B.n754 B.n368 163.367
R1588 B.n754 B.n366 163.367
R1589 B.n758 B.n366 163.367
R1590 B.n758 B.n360 163.367
R1591 B.n766 B.n360 163.367
R1592 B.n766 B.n358 163.367
R1593 B.n770 B.n358 163.367
R1594 B.n770 B.n352 163.367
R1595 B.n778 B.n352 163.367
R1596 B.n778 B.n350 163.367
R1597 B.n782 B.n350 163.367
R1598 B.n782 B.n344 163.367
R1599 B.n790 B.n344 163.367
R1600 B.n790 B.n342 163.367
R1601 B.n794 B.n342 163.367
R1602 B.n794 B.n337 163.367
R1603 B.n803 B.n337 163.367
R1604 B.n803 B.n335 163.367
R1605 B.n808 B.n335 163.367
R1606 B.n808 B.n329 163.367
R1607 B.n816 B.n329 163.367
R1608 B.n817 B.n816 163.367
R1609 B.n817 B.n5 163.367
R1610 B.n6 B.n5 163.367
R1611 B.n7 B.n6 163.367
R1612 B.n822 B.n7 163.367
R1613 B.n822 B.n12 163.367
R1614 B.n13 B.n12 163.367
R1615 B.n14 B.n13 163.367
R1616 B.n827 B.n14 163.367
R1617 B.n827 B.n19 163.367
R1618 B.n20 B.n19 163.367
R1619 B.n21 B.n20 163.367
R1620 B.n832 B.n21 163.367
R1621 B.n832 B.n26 163.367
R1622 B.n27 B.n26 163.367
R1623 B.n28 B.n27 163.367
R1624 B.n837 B.n28 163.367
R1625 B.n837 B.n33 163.367
R1626 B.n34 B.n33 163.367
R1627 B.n35 B.n34 163.367
R1628 B.n842 B.n35 163.367
R1629 B.n842 B.n40 163.367
R1630 B.n41 B.n40 163.367
R1631 B.n42 B.n41 163.367
R1632 B.n847 B.n42 163.367
R1633 B.n847 B.n47 163.367
R1634 B.n48 B.n47 163.367
R1635 B.n49 B.n48 163.367
R1636 B.n852 B.n49 163.367
R1637 B.n852 B.n54 163.367
R1638 B.n55 B.n54 163.367
R1639 B.n56 B.n55 163.367
R1640 B.n857 B.n56 163.367
R1641 B.n857 B.n61 163.367
R1642 B.n62 B.n61 163.367
R1643 B.n63 B.n62 163.367
R1644 B.n862 B.n63 163.367
R1645 B.n862 B.n68 163.367
R1646 B.n69 B.n68 163.367
R1647 B.n70 B.n69 163.367
R1648 B.n867 B.n70 163.367
R1649 B.n867 B.n75 163.367
R1650 B.n76 B.n75 163.367
R1651 B.n77 B.n76 163.367
R1652 B.n872 B.n77 163.367
R1653 B.n872 B.n82 163.367
R1654 B.n83 B.n82 163.367
R1655 B.n84 B.n83 163.367
R1656 B.n877 B.n84 163.367
R1657 B.n877 B.n89 163.367
R1658 B.n90 B.n89 163.367
R1659 B.n91 B.n90 163.367
R1660 B.n142 B.n91 163.367
R1661 B.n148 B.n95 163.367
R1662 B.n152 B.n151 163.367
R1663 B.n156 B.n155 163.367
R1664 B.n160 B.n159 163.367
R1665 B.n164 B.n163 163.367
R1666 B.n168 B.n167 163.367
R1667 B.n172 B.n171 163.367
R1668 B.n176 B.n175 163.367
R1669 B.n180 B.n179 163.367
R1670 B.n184 B.n183 163.367
R1671 B.n188 B.n187 163.367
R1672 B.n192 B.n191 163.367
R1673 B.n196 B.n195 163.367
R1674 B.n200 B.n199 163.367
R1675 B.n204 B.n203 163.367
R1676 B.n208 B.n207 163.367
R1677 B.n212 B.n211 163.367
R1678 B.n216 B.n215 163.367
R1679 B.n220 B.n219 163.367
R1680 B.n224 B.n223 163.367
R1681 B.n228 B.n227 163.367
R1682 B.n232 B.n231 163.367
R1683 B.n236 B.n235 163.367
R1684 B.n240 B.n239 163.367
R1685 B.n244 B.n243 163.367
R1686 B.n249 B.n248 163.367
R1687 B.n253 B.n252 163.367
R1688 B.n257 B.n256 163.367
R1689 B.n261 B.n260 163.367
R1690 B.n265 B.n264 163.367
R1691 B.n269 B.n268 163.367
R1692 B.n273 B.n272 163.367
R1693 B.n277 B.n276 163.367
R1694 B.n281 B.n280 163.367
R1695 B.n285 B.n284 163.367
R1696 B.n289 B.n288 163.367
R1697 B.n293 B.n292 163.367
R1698 B.n297 B.n296 163.367
R1699 B.n301 B.n300 163.367
R1700 B.n305 B.n304 163.367
R1701 B.n309 B.n308 163.367
R1702 B.n313 B.n312 163.367
R1703 B.n317 B.n316 163.367
R1704 B.n321 B.n320 163.367
R1705 B.n325 B.n324 163.367
R1706 B.n884 B.n141 163.367
R1707 B.n661 B.n424 75.8186
R1708 B.n885 B.n92 75.8186
R1709 B.n663 B.n662 71.676
R1710 B.n473 B.n428 71.676
R1711 B.n655 B.n429 71.676
R1712 B.n651 B.n430 71.676
R1713 B.n647 B.n431 71.676
R1714 B.n643 B.n432 71.676
R1715 B.n639 B.n433 71.676
R1716 B.n635 B.n434 71.676
R1717 B.n631 B.n435 71.676
R1718 B.n627 B.n436 71.676
R1719 B.n623 B.n437 71.676
R1720 B.n619 B.n438 71.676
R1721 B.n615 B.n439 71.676
R1722 B.n611 B.n440 71.676
R1723 B.n607 B.n441 71.676
R1724 B.n603 B.n442 71.676
R1725 B.n599 B.n443 71.676
R1726 B.n595 B.n444 71.676
R1727 B.n591 B.n445 71.676
R1728 B.n587 B.n446 71.676
R1729 B.n583 B.n447 71.676
R1730 B.n578 B.n448 71.676
R1731 B.n574 B.n449 71.676
R1732 B.n570 B.n450 71.676
R1733 B.n566 B.n451 71.676
R1734 B.n562 B.n452 71.676
R1735 B.n558 B.n453 71.676
R1736 B.n554 B.n454 71.676
R1737 B.n550 B.n455 71.676
R1738 B.n546 B.n456 71.676
R1739 B.n542 B.n457 71.676
R1740 B.n538 B.n458 71.676
R1741 B.n534 B.n459 71.676
R1742 B.n530 B.n460 71.676
R1743 B.n526 B.n461 71.676
R1744 B.n522 B.n462 71.676
R1745 B.n518 B.n463 71.676
R1746 B.n514 B.n464 71.676
R1747 B.n510 B.n465 71.676
R1748 B.n506 B.n466 71.676
R1749 B.n502 B.n467 71.676
R1750 B.n498 B.n468 71.676
R1751 B.n494 B.n469 71.676
R1752 B.n490 B.n470 71.676
R1753 B.n486 B.n471 71.676
R1754 B.n482 B.n472 71.676
R1755 B.n887 B.n886 71.676
R1756 B.n148 B.n96 71.676
R1757 B.n152 B.n97 71.676
R1758 B.n156 B.n98 71.676
R1759 B.n160 B.n99 71.676
R1760 B.n164 B.n100 71.676
R1761 B.n168 B.n101 71.676
R1762 B.n172 B.n102 71.676
R1763 B.n176 B.n103 71.676
R1764 B.n180 B.n104 71.676
R1765 B.n184 B.n105 71.676
R1766 B.n188 B.n106 71.676
R1767 B.n192 B.n107 71.676
R1768 B.n196 B.n108 71.676
R1769 B.n200 B.n109 71.676
R1770 B.n204 B.n110 71.676
R1771 B.n208 B.n111 71.676
R1772 B.n212 B.n112 71.676
R1773 B.n216 B.n113 71.676
R1774 B.n220 B.n114 71.676
R1775 B.n224 B.n115 71.676
R1776 B.n228 B.n116 71.676
R1777 B.n232 B.n117 71.676
R1778 B.n236 B.n118 71.676
R1779 B.n240 B.n119 71.676
R1780 B.n244 B.n120 71.676
R1781 B.n249 B.n121 71.676
R1782 B.n253 B.n122 71.676
R1783 B.n257 B.n123 71.676
R1784 B.n261 B.n124 71.676
R1785 B.n265 B.n125 71.676
R1786 B.n269 B.n126 71.676
R1787 B.n273 B.n127 71.676
R1788 B.n277 B.n128 71.676
R1789 B.n281 B.n129 71.676
R1790 B.n285 B.n130 71.676
R1791 B.n289 B.n131 71.676
R1792 B.n293 B.n132 71.676
R1793 B.n297 B.n133 71.676
R1794 B.n301 B.n134 71.676
R1795 B.n305 B.n135 71.676
R1796 B.n309 B.n136 71.676
R1797 B.n313 B.n137 71.676
R1798 B.n317 B.n138 71.676
R1799 B.n321 B.n139 71.676
R1800 B.n325 B.n140 71.676
R1801 B.n141 B.n140 71.676
R1802 B.n324 B.n139 71.676
R1803 B.n320 B.n138 71.676
R1804 B.n316 B.n137 71.676
R1805 B.n312 B.n136 71.676
R1806 B.n308 B.n135 71.676
R1807 B.n304 B.n134 71.676
R1808 B.n300 B.n133 71.676
R1809 B.n296 B.n132 71.676
R1810 B.n292 B.n131 71.676
R1811 B.n288 B.n130 71.676
R1812 B.n284 B.n129 71.676
R1813 B.n280 B.n128 71.676
R1814 B.n276 B.n127 71.676
R1815 B.n272 B.n126 71.676
R1816 B.n268 B.n125 71.676
R1817 B.n264 B.n124 71.676
R1818 B.n260 B.n123 71.676
R1819 B.n256 B.n122 71.676
R1820 B.n252 B.n121 71.676
R1821 B.n248 B.n120 71.676
R1822 B.n243 B.n119 71.676
R1823 B.n239 B.n118 71.676
R1824 B.n235 B.n117 71.676
R1825 B.n231 B.n116 71.676
R1826 B.n227 B.n115 71.676
R1827 B.n223 B.n114 71.676
R1828 B.n219 B.n113 71.676
R1829 B.n215 B.n112 71.676
R1830 B.n211 B.n111 71.676
R1831 B.n207 B.n110 71.676
R1832 B.n203 B.n109 71.676
R1833 B.n199 B.n108 71.676
R1834 B.n195 B.n107 71.676
R1835 B.n191 B.n106 71.676
R1836 B.n187 B.n105 71.676
R1837 B.n183 B.n104 71.676
R1838 B.n179 B.n103 71.676
R1839 B.n175 B.n102 71.676
R1840 B.n171 B.n101 71.676
R1841 B.n167 B.n100 71.676
R1842 B.n163 B.n99 71.676
R1843 B.n159 B.n98 71.676
R1844 B.n155 B.n97 71.676
R1845 B.n151 B.n96 71.676
R1846 B.n886 B.n95 71.676
R1847 B.n662 B.n427 71.676
R1848 B.n656 B.n428 71.676
R1849 B.n652 B.n429 71.676
R1850 B.n648 B.n430 71.676
R1851 B.n644 B.n431 71.676
R1852 B.n640 B.n432 71.676
R1853 B.n636 B.n433 71.676
R1854 B.n632 B.n434 71.676
R1855 B.n628 B.n435 71.676
R1856 B.n624 B.n436 71.676
R1857 B.n620 B.n437 71.676
R1858 B.n616 B.n438 71.676
R1859 B.n612 B.n439 71.676
R1860 B.n608 B.n440 71.676
R1861 B.n604 B.n441 71.676
R1862 B.n600 B.n442 71.676
R1863 B.n596 B.n443 71.676
R1864 B.n592 B.n444 71.676
R1865 B.n588 B.n445 71.676
R1866 B.n584 B.n446 71.676
R1867 B.n579 B.n447 71.676
R1868 B.n575 B.n448 71.676
R1869 B.n571 B.n449 71.676
R1870 B.n567 B.n450 71.676
R1871 B.n563 B.n451 71.676
R1872 B.n559 B.n452 71.676
R1873 B.n555 B.n453 71.676
R1874 B.n551 B.n454 71.676
R1875 B.n547 B.n455 71.676
R1876 B.n543 B.n456 71.676
R1877 B.n539 B.n457 71.676
R1878 B.n535 B.n458 71.676
R1879 B.n531 B.n459 71.676
R1880 B.n527 B.n460 71.676
R1881 B.n523 B.n461 71.676
R1882 B.n519 B.n462 71.676
R1883 B.n515 B.n463 71.676
R1884 B.n511 B.n464 71.676
R1885 B.n507 B.n465 71.676
R1886 B.n503 B.n466 71.676
R1887 B.n499 B.n467 71.676
R1888 B.n495 B.n468 71.676
R1889 B.n491 B.n469 71.676
R1890 B.n487 B.n470 71.676
R1891 B.n483 B.n471 71.676
R1892 B.n479 B.n472 71.676
R1893 B.n477 B.n476 70.5944
R1894 B.n475 B.n474 70.5944
R1895 B.n146 B.n145 70.5944
R1896 B.n144 B.n143 70.5944
R1897 B.n478 B.n477 59.5399
R1898 B.n581 B.n475 59.5399
R1899 B.n147 B.n146 59.5399
R1900 B.n246 B.n144 59.5399
R1901 B.n668 B.n424 43.3251
R1902 B.n668 B.n420 43.3251
R1903 B.n674 B.n420 43.3251
R1904 B.n674 B.n416 43.3251
R1905 B.n680 B.n416 43.3251
R1906 B.n680 B.n412 43.3251
R1907 B.n687 B.n412 43.3251
R1908 B.n687 B.n686 43.3251
R1909 B.n693 B.n405 43.3251
R1910 B.n699 B.n405 43.3251
R1911 B.n699 B.n401 43.3251
R1912 B.n705 B.n401 43.3251
R1913 B.n705 B.n397 43.3251
R1914 B.n711 B.n397 43.3251
R1915 B.n711 B.n393 43.3251
R1916 B.n717 B.n393 43.3251
R1917 B.n717 B.n389 43.3251
R1918 B.n723 B.n389 43.3251
R1919 B.n723 B.n384 43.3251
R1920 B.n729 B.n384 43.3251
R1921 B.n729 B.n385 43.3251
R1922 B.n735 B.n377 43.3251
R1923 B.n741 B.n377 43.3251
R1924 B.n741 B.n373 43.3251
R1925 B.n747 B.n373 43.3251
R1926 B.n747 B.n369 43.3251
R1927 B.n753 B.n369 43.3251
R1928 B.n753 B.n365 43.3251
R1929 B.n759 B.n365 43.3251
R1930 B.n759 B.n361 43.3251
R1931 B.n765 B.n361 43.3251
R1932 B.n771 B.n357 43.3251
R1933 B.n771 B.n353 43.3251
R1934 B.n777 B.n353 43.3251
R1935 B.n777 B.n349 43.3251
R1936 B.n783 B.n349 43.3251
R1937 B.n783 B.n345 43.3251
R1938 B.n789 B.n345 43.3251
R1939 B.n789 B.n341 43.3251
R1940 B.n796 B.n341 43.3251
R1941 B.n796 B.n795 43.3251
R1942 B.n802 B.n334 43.3251
R1943 B.n809 B.n334 43.3251
R1944 B.n809 B.n330 43.3251
R1945 B.n815 B.n330 43.3251
R1946 B.n815 B.n4 43.3251
R1947 B.n990 B.n4 43.3251
R1948 B.n990 B.n989 43.3251
R1949 B.n989 B.n988 43.3251
R1950 B.n988 B.n8 43.3251
R1951 B.n982 B.n8 43.3251
R1952 B.n982 B.n981 43.3251
R1953 B.n981 B.n980 43.3251
R1954 B.n974 B.n18 43.3251
R1955 B.n974 B.n973 43.3251
R1956 B.n973 B.n972 43.3251
R1957 B.n972 B.n22 43.3251
R1958 B.n966 B.n22 43.3251
R1959 B.n966 B.n965 43.3251
R1960 B.n965 B.n964 43.3251
R1961 B.n964 B.n29 43.3251
R1962 B.n958 B.n29 43.3251
R1963 B.n958 B.n957 43.3251
R1964 B.n956 B.n36 43.3251
R1965 B.n950 B.n36 43.3251
R1966 B.n950 B.n949 43.3251
R1967 B.n949 B.n948 43.3251
R1968 B.n948 B.n43 43.3251
R1969 B.n942 B.n43 43.3251
R1970 B.n942 B.n941 43.3251
R1971 B.n941 B.n940 43.3251
R1972 B.n940 B.n50 43.3251
R1973 B.n934 B.n50 43.3251
R1974 B.n933 B.n932 43.3251
R1975 B.n932 B.n57 43.3251
R1976 B.n926 B.n57 43.3251
R1977 B.n926 B.n925 43.3251
R1978 B.n925 B.n924 43.3251
R1979 B.n924 B.n64 43.3251
R1980 B.n918 B.n64 43.3251
R1981 B.n918 B.n917 43.3251
R1982 B.n917 B.n916 43.3251
R1983 B.n916 B.n71 43.3251
R1984 B.n910 B.n71 43.3251
R1985 B.n910 B.n909 43.3251
R1986 B.n909 B.n908 43.3251
R1987 B.n902 B.n81 43.3251
R1988 B.n902 B.n901 43.3251
R1989 B.n901 B.n900 43.3251
R1990 B.n900 B.n85 43.3251
R1991 B.n894 B.n85 43.3251
R1992 B.n894 B.n893 43.3251
R1993 B.n893 B.n892 43.3251
R1994 B.n892 B.n92 43.3251
R1995 B.n802 B.t3 41.4138
R1996 B.n980 B.t2 41.4138
R1997 B.n686 B.t7 31.2197
R1998 B.n81 B.t11 31.2197
R1999 B.n889 B.n888 30.4395
R2000 B.n883 B.n882 30.4395
R2001 B.n480 B.n422 30.4395
R2002 B.n665 B.n664 30.4395
R2003 B.t1 B.n357 28.6712
R2004 B.n957 B.t0 28.6712
R2005 B.n385 B.t4 27.397
R2006 B.t5 B.n933 27.397
R2007 B B.n992 18.0485
R2008 B.n735 B.t4 15.9287
R2009 B.n934 B.t5 15.9287
R2010 B.n765 B.t1 14.6544
R2011 B.t0 B.n956 14.6544
R2012 B.n693 B.t7 12.1059
R2013 B.n908 B.t11 12.1059
R2014 B.n888 B.n94 10.6151
R2015 B.n149 B.n94 10.6151
R2016 B.n150 B.n149 10.6151
R2017 B.n153 B.n150 10.6151
R2018 B.n154 B.n153 10.6151
R2019 B.n157 B.n154 10.6151
R2020 B.n158 B.n157 10.6151
R2021 B.n161 B.n158 10.6151
R2022 B.n162 B.n161 10.6151
R2023 B.n165 B.n162 10.6151
R2024 B.n166 B.n165 10.6151
R2025 B.n169 B.n166 10.6151
R2026 B.n170 B.n169 10.6151
R2027 B.n173 B.n170 10.6151
R2028 B.n174 B.n173 10.6151
R2029 B.n177 B.n174 10.6151
R2030 B.n178 B.n177 10.6151
R2031 B.n181 B.n178 10.6151
R2032 B.n182 B.n181 10.6151
R2033 B.n185 B.n182 10.6151
R2034 B.n186 B.n185 10.6151
R2035 B.n189 B.n186 10.6151
R2036 B.n190 B.n189 10.6151
R2037 B.n193 B.n190 10.6151
R2038 B.n194 B.n193 10.6151
R2039 B.n197 B.n194 10.6151
R2040 B.n198 B.n197 10.6151
R2041 B.n201 B.n198 10.6151
R2042 B.n202 B.n201 10.6151
R2043 B.n205 B.n202 10.6151
R2044 B.n206 B.n205 10.6151
R2045 B.n209 B.n206 10.6151
R2046 B.n210 B.n209 10.6151
R2047 B.n213 B.n210 10.6151
R2048 B.n214 B.n213 10.6151
R2049 B.n217 B.n214 10.6151
R2050 B.n218 B.n217 10.6151
R2051 B.n221 B.n218 10.6151
R2052 B.n222 B.n221 10.6151
R2053 B.n225 B.n222 10.6151
R2054 B.n226 B.n225 10.6151
R2055 B.n230 B.n229 10.6151
R2056 B.n233 B.n230 10.6151
R2057 B.n234 B.n233 10.6151
R2058 B.n237 B.n234 10.6151
R2059 B.n238 B.n237 10.6151
R2060 B.n241 B.n238 10.6151
R2061 B.n242 B.n241 10.6151
R2062 B.n245 B.n242 10.6151
R2063 B.n250 B.n247 10.6151
R2064 B.n251 B.n250 10.6151
R2065 B.n254 B.n251 10.6151
R2066 B.n255 B.n254 10.6151
R2067 B.n258 B.n255 10.6151
R2068 B.n259 B.n258 10.6151
R2069 B.n262 B.n259 10.6151
R2070 B.n263 B.n262 10.6151
R2071 B.n266 B.n263 10.6151
R2072 B.n267 B.n266 10.6151
R2073 B.n270 B.n267 10.6151
R2074 B.n271 B.n270 10.6151
R2075 B.n274 B.n271 10.6151
R2076 B.n275 B.n274 10.6151
R2077 B.n278 B.n275 10.6151
R2078 B.n279 B.n278 10.6151
R2079 B.n282 B.n279 10.6151
R2080 B.n283 B.n282 10.6151
R2081 B.n286 B.n283 10.6151
R2082 B.n287 B.n286 10.6151
R2083 B.n290 B.n287 10.6151
R2084 B.n291 B.n290 10.6151
R2085 B.n294 B.n291 10.6151
R2086 B.n295 B.n294 10.6151
R2087 B.n298 B.n295 10.6151
R2088 B.n299 B.n298 10.6151
R2089 B.n302 B.n299 10.6151
R2090 B.n303 B.n302 10.6151
R2091 B.n306 B.n303 10.6151
R2092 B.n307 B.n306 10.6151
R2093 B.n310 B.n307 10.6151
R2094 B.n311 B.n310 10.6151
R2095 B.n314 B.n311 10.6151
R2096 B.n315 B.n314 10.6151
R2097 B.n318 B.n315 10.6151
R2098 B.n319 B.n318 10.6151
R2099 B.n322 B.n319 10.6151
R2100 B.n323 B.n322 10.6151
R2101 B.n326 B.n323 10.6151
R2102 B.n327 B.n326 10.6151
R2103 B.n883 B.n327 10.6151
R2104 B.n670 B.n422 10.6151
R2105 B.n671 B.n670 10.6151
R2106 B.n672 B.n671 10.6151
R2107 B.n672 B.n414 10.6151
R2108 B.n682 B.n414 10.6151
R2109 B.n683 B.n682 10.6151
R2110 B.n684 B.n683 10.6151
R2111 B.n684 B.n407 10.6151
R2112 B.n695 B.n407 10.6151
R2113 B.n696 B.n695 10.6151
R2114 B.n697 B.n696 10.6151
R2115 B.n697 B.n399 10.6151
R2116 B.n707 B.n399 10.6151
R2117 B.n708 B.n707 10.6151
R2118 B.n709 B.n708 10.6151
R2119 B.n709 B.n391 10.6151
R2120 B.n719 B.n391 10.6151
R2121 B.n720 B.n719 10.6151
R2122 B.n721 B.n720 10.6151
R2123 B.n721 B.n382 10.6151
R2124 B.n731 B.n382 10.6151
R2125 B.n732 B.n731 10.6151
R2126 B.n733 B.n732 10.6151
R2127 B.n733 B.n375 10.6151
R2128 B.n743 B.n375 10.6151
R2129 B.n744 B.n743 10.6151
R2130 B.n745 B.n744 10.6151
R2131 B.n745 B.n367 10.6151
R2132 B.n755 B.n367 10.6151
R2133 B.n756 B.n755 10.6151
R2134 B.n757 B.n756 10.6151
R2135 B.n757 B.n359 10.6151
R2136 B.n767 B.n359 10.6151
R2137 B.n768 B.n767 10.6151
R2138 B.n769 B.n768 10.6151
R2139 B.n769 B.n351 10.6151
R2140 B.n779 B.n351 10.6151
R2141 B.n780 B.n779 10.6151
R2142 B.n781 B.n780 10.6151
R2143 B.n781 B.n343 10.6151
R2144 B.n791 B.n343 10.6151
R2145 B.n792 B.n791 10.6151
R2146 B.n793 B.n792 10.6151
R2147 B.n793 B.n336 10.6151
R2148 B.n804 B.n336 10.6151
R2149 B.n805 B.n804 10.6151
R2150 B.n807 B.n805 10.6151
R2151 B.n807 B.n806 10.6151
R2152 B.n806 B.n328 10.6151
R2153 B.n818 B.n328 10.6151
R2154 B.n819 B.n818 10.6151
R2155 B.n820 B.n819 10.6151
R2156 B.n821 B.n820 10.6151
R2157 B.n823 B.n821 10.6151
R2158 B.n824 B.n823 10.6151
R2159 B.n825 B.n824 10.6151
R2160 B.n826 B.n825 10.6151
R2161 B.n828 B.n826 10.6151
R2162 B.n829 B.n828 10.6151
R2163 B.n830 B.n829 10.6151
R2164 B.n831 B.n830 10.6151
R2165 B.n833 B.n831 10.6151
R2166 B.n834 B.n833 10.6151
R2167 B.n835 B.n834 10.6151
R2168 B.n836 B.n835 10.6151
R2169 B.n838 B.n836 10.6151
R2170 B.n839 B.n838 10.6151
R2171 B.n840 B.n839 10.6151
R2172 B.n841 B.n840 10.6151
R2173 B.n843 B.n841 10.6151
R2174 B.n844 B.n843 10.6151
R2175 B.n845 B.n844 10.6151
R2176 B.n846 B.n845 10.6151
R2177 B.n848 B.n846 10.6151
R2178 B.n849 B.n848 10.6151
R2179 B.n850 B.n849 10.6151
R2180 B.n851 B.n850 10.6151
R2181 B.n853 B.n851 10.6151
R2182 B.n854 B.n853 10.6151
R2183 B.n855 B.n854 10.6151
R2184 B.n856 B.n855 10.6151
R2185 B.n858 B.n856 10.6151
R2186 B.n859 B.n858 10.6151
R2187 B.n860 B.n859 10.6151
R2188 B.n861 B.n860 10.6151
R2189 B.n863 B.n861 10.6151
R2190 B.n864 B.n863 10.6151
R2191 B.n865 B.n864 10.6151
R2192 B.n866 B.n865 10.6151
R2193 B.n868 B.n866 10.6151
R2194 B.n869 B.n868 10.6151
R2195 B.n870 B.n869 10.6151
R2196 B.n871 B.n870 10.6151
R2197 B.n873 B.n871 10.6151
R2198 B.n874 B.n873 10.6151
R2199 B.n875 B.n874 10.6151
R2200 B.n876 B.n875 10.6151
R2201 B.n878 B.n876 10.6151
R2202 B.n879 B.n878 10.6151
R2203 B.n880 B.n879 10.6151
R2204 B.n881 B.n880 10.6151
R2205 B.n882 B.n881 10.6151
R2206 B.n664 B.n426 10.6151
R2207 B.n659 B.n426 10.6151
R2208 B.n659 B.n658 10.6151
R2209 B.n658 B.n657 10.6151
R2210 B.n657 B.n654 10.6151
R2211 B.n654 B.n653 10.6151
R2212 B.n653 B.n650 10.6151
R2213 B.n650 B.n649 10.6151
R2214 B.n649 B.n646 10.6151
R2215 B.n646 B.n645 10.6151
R2216 B.n645 B.n642 10.6151
R2217 B.n642 B.n641 10.6151
R2218 B.n641 B.n638 10.6151
R2219 B.n638 B.n637 10.6151
R2220 B.n637 B.n634 10.6151
R2221 B.n634 B.n633 10.6151
R2222 B.n633 B.n630 10.6151
R2223 B.n630 B.n629 10.6151
R2224 B.n629 B.n626 10.6151
R2225 B.n626 B.n625 10.6151
R2226 B.n625 B.n622 10.6151
R2227 B.n622 B.n621 10.6151
R2228 B.n621 B.n618 10.6151
R2229 B.n618 B.n617 10.6151
R2230 B.n617 B.n614 10.6151
R2231 B.n614 B.n613 10.6151
R2232 B.n613 B.n610 10.6151
R2233 B.n610 B.n609 10.6151
R2234 B.n609 B.n606 10.6151
R2235 B.n606 B.n605 10.6151
R2236 B.n605 B.n602 10.6151
R2237 B.n602 B.n601 10.6151
R2238 B.n601 B.n598 10.6151
R2239 B.n598 B.n597 10.6151
R2240 B.n597 B.n594 10.6151
R2241 B.n594 B.n593 10.6151
R2242 B.n593 B.n590 10.6151
R2243 B.n590 B.n589 10.6151
R2244 B.n589 B.n586 10.6151
R2245 B.n586 B.n585 10.6151
R2246 B.n585 B.n582 10.6151
R2247 B.n580 B.n577 10.6151
R2248 B.n577 B.n576 10.6151
R2249 B.n576 B.n573 10.6151
R2250 B.n573 B.n572 10.6151
R2251 B.n572 B.n569 10.6151
R2252 B.n569 B.n568 10.6151
R2253 B.n568 B.n565 10.6151
R2254 B.n565 B.n564 10.6151
R2255 B.n561 B.n560 10.6151
R2256 B.n560 B.n557 10.6151
R2257 B.n557 B.n556 10.6151
R2258 B.n556 B.n553 10.6151
R2259 B.n553 B.n552 10.6151
R2260 B.n552 B.n549 10.6151
R2261 B.n549 B.n548 10.6151
R2262 B.n548 B.n545 10.6151
R2263 B.n545 B.n544 10.6151
R2264 B.n544 B.n541 10.6151
R2265 B.n541 B.n540 10.6151
R2266 B.n540 B.n537 10.6151
R2267 B.n537 B.n536 10.6151
R2268 B.n536 B.n533 10.6151
R2269 B.n533 B.n532 10.6151
R2270 B.n532 B.n529 10.6151
R2271 B.n529 B.n528 10.6151
R2272 B.n528 B.n525 10.6151
R2273 B.n525 B.n524 10.6151
R2274 B.n524 B.n521 10.6151
R2275 B.n521 B.n520 10.6151
R2276 B.n520 B.n517 10.6151
R2277 B.n517 B.n516 10.6151
R2278 B.n516 B.n513 10.6151
R2279 B.n513 B.n512 10.6151
R2280 B.n512 B.n509 10.6151
R2281 B.n509 B.n508 10.6151
R2282 B.n508 B.n505 10.6151
R2283 B.n505 B.n504 10.6151
R2284 B.n504 B.n501 10.6151
R2285 B.n501 B.n500 10.6151
R2286 B.n500 B.n497 10.6151
R2287 B.n497 B.n496 10.6151
R2288 B.n496 B.n493 10.6151
R2289 B.n493 B.n492 10.6151
R2290 B.n492 B.n489 10.6151
R2291 B.n489 B.n488 10.6151
R2292 B.n488 B.n485 10.6151
R2293 B.n485 B.n484 10.6151
R2294 B.n484 B.n481 10.6151
R2295 B.n481 B.n480 10.6151
R2296 B.n666 B.n665 10.6151
R2297 B.n666 B.n418 10.6151
R2298 B.n676 B.n418 10.6151
R2299 B.n677 B.n676 10.6151
R2300 B.n678 B.n677 10.6151
R2301 B.n678 B.n410 10.6151
R2302 B.n689 B.n410 10.6151
R2303 B.n690 B.n689 10.6151
R2304 B.n691 B.n690 10.6151
R2305 B.n691 B.n403 10.6151
R2306 B.n701 B.n403 10.6151
R2307 B.n702 B.n701 10.6151
R2308 B.n703 B.n702 10.6151
R2309 B.n703 B.n395 10.6151
R2310 B.n713 B.n395 10.6151
R2311 B.n714 B.n713 10.6151
R2312 B.n715 B.n714 10.6151
R2313 B.n715 B.n387 10.6151
R2314 B.n725 B.n387 10.6151
R2315 B.n726 B.n725 10.6151
R2316 B.n727 B.n726 10.6151
R2317 B.n727 B.n379 10.6151
R2318 B.n737 B.n379 10.6151
R2319 B.n738 B.n737 10.6151
R2320 B.n739 B.n738 10.6151
R2321 B.n739 B.n371 10.6151
R2322 B.n749 B.n371 10.6151
R2323 B.n750 B.n749 10.6151
R2324 B.n751 B.n750 10.6151
R2325 B.n751 B.n363 10.6151
R2326 B.n761 B.n363 10.6151
R2327 B.n762 B.n761 10.6151
R2328 B.n763 B.n762 10.6151
R2329 B.n763 B.n355 10.6151
R2330 B.n773 B.n355 10.6151
R2331 B.n774 B.n773 10.6151
R2332 B.n775 B.n774 10.6151
R2333 B.n775 B.n347 10.6151
R2334 B.n785 B.n347 10.6151
R2335 B.n786 B.n785 10.6151
R2336 B.n787 B.n786 10.6151
R2337 B.n787 B.n339 10.6151
R2338 B.n798 B.n339 10.6151
R2339 B.n799 B.n798 10.6151
R2340 B.n800 B.n799 10.6151
R2341 B.n800 B.n332 10.6151
R2342 B.n811 B.n332 10.6151
R2343 B.n812 B.n811 10.6151
R2344 B.n813 B.n812 10.6151
R2345 B.n813 B.n0 10.6151
R2346 B.n986 B.n1 10.6151
R2347 B.n986 B.n985 10.6151
R2348 B.n985 B.n984 10.6151
R2349 B.n984 B.n10 10.6151
R2350 B.n978 B.n10 10.6151
R2351 B.n978 B.n977 10.6151
R2352 B.n977 B.n976 10.6151
R2353 B.n976 B.n16 10.6151
R2354 B.n970 B.n16 10.6151
R2355 B.n970 B.n969 10.6151
R2356 B.n969 B.n968 10.6151
R2357 B.n968 B.n24 10.6151
R2358 B.n962 B.n24 10.6151
R2359 B.n962 B.n961 10.6151
R2360 B.n961 B.n960 10.6151
R2361 B.n960 B.n31 10.6151
R2362 B.n954 B.n31 10.6151
R2363 B.n954 B.n953 10.6151
R2364 B.n953 B.n952 10.6151
R2365 B.n952 B.n38 10.6151
R2366 B.n946 B.n38 10.6151
R2367 B.n946 B.n945 10.6151
R2368 B.n945 B.n944 10.6151
R2369 B.n944 B.n45 10.6151
R2370 B.n938 B.n45 10.6151
R2371 B.n938 B.n937 10.6151
R2372 B.n937 B.n936 10.6151
R2373 B.n936 B.n52 10.6151
R2374 B.n930 B.n52 10.6151
R2375 B.n930 B.n929 10.6151
R2376 B.n929 B.n928 10.6151
R2377 B.n928 B.n59 10.6151
R2378 B.n922 B.n59 10.6151
R2379 B.n922 B.n921 10.6151
R2380 B.n921 B.n920 10.6151
R2381 B.n920 B.n66 10.6151
R2382 B.n914 B.n66 10.6151
R2383 B.n914 B.n913 10.6151
R2384 B.n913 B.n912 10.6151
R2385 B.n912 B.n73 10.6151
R2386 B.n906 B.n73 10.6151
R2387 B.n906 B.n905 10.6151
R2388 B.n905 B.n904 10.6151
R2389 B.n904 B.n79 10.6151
R2390 B.n898 B.n79 10.6151
R2391 B.n898 B.n897 10.6151
R2392 B.n897 B.n896 10.6151
R2393 B.n896 B.n87 10.6151
R2394 B.n890 B.n87 10.6151
R2395 B.n890 B.n889 10.6151
R2396 B.n229 B.n147 6.5566
R2397 B.n246 B.n245 6.5566
R2398 B.n581 B.n580 6.5566
R2399 B.n564 B.n478 6.5566
R2400 B.n226 B.n147 4.05904
R2401 B.n247 B.n246 4.05904
R2402 B.n582 B.n581 4.05904
R2403 B.n561 B.n478 4.05904
R2404 B.n992 B.n0 2.81026
R2405 B.n992 B.n1 2.81026
R2406 B.n795 B.t3 1.91188
R2407 B.n18 B.t2 1.91188
R2408 VN.n34 VN.n33 161.3
R2409 VN.n32 VN.n19 161.3
R2410 VN.n31 VN.n30 161.3
R2411 VN.n29 VN.n20 161.3
R2412 VN.n28 VN.n27 161.3
R2413 VN.n26 VN.n21 161.3
R2414 VN.n25 VN.n24 161.3
R2415 VN.n16 VN.n15 161.3
R2416 VN.n14 VN.n1 161.3
R2417 VN.n13 VN.n12 161.3
R2418 VN.n11 VN.n2 161.3
R2419 VN.n10 VN.n9 161.3
R2420 VN.n8 VN.n3 161.3
R2421 VN.n7 VN.n6 161.3
R2422 VN.n23 VN.t4 120.597
R2423 VN.n5 VN.t0 120.597
R2424 VN.n4 VN.t3 87.2993
R2425 VN.n0 VN.t5 87.2993
R2426 VN.n22 VN.t2 87.2993
R2427 VN.n18 VN.t1 87.2993
R2428 VN.n17 VN.n0 70.9831
R2429 VN.n35 VN.n18 70.9831
R2430 VN.n5 VN.n4 62.0573
R2431 VN.n23 VN.n22 62.0573
R2432 VN VN.n35 51.8011
R2433 VN.n13 VN.n2 47.2923
R2434 VN.n31 VN.n20 47.2923
R2435 VN.n9 VN.n2 33.6945
R2436 VN.n27 VN.n20 33.6945
R2437 VN.n8 VN.n7 24.4675
R2438 VN.n9 VN.n8 24.4675
R2439 VN.n14 VN.n13 24.4675
R2440 VN.n15 VN.n14 24.4675
R2441 VN.n27 VN.n26 24.4675
R2442 VN.n26 VN.n25 24.4675
R2443 VN.n33 VN.n32 24.4675
R2444 VN.n32 VN.n31 24.4675
R2445 VN.n15 VN.n0 19.0848
R2446 VN.n33 VN.n18 19.0848
R2447 VN.n7 VN.n4 12.234
R2448 VN.n25 VN.n22 12.234
R2449 VN.n24 VN.n23 3.94734
R2450 VN.n6 VN.n5 3.94734
R2451 VN.n35 VN.n34 0.354971
R2452 VN.n17 VN.n16 0.354971
R2453 VN VN.n17 0.26696
R2454 VN.n34 VN.n19 0.189894
R2455 VN.n30 VN.n19 0.189894
R2456 VN.n30 VN.n29 0.189894
R2457 VN.n29 VN.n28 0.189894
R2458 VN.n28 VN.n21 0.189894
R2459 VN.n24 VN.n21 0.189894
R2460 VN.n6 VN.n3 0.189894
R2461 VN.n10 VN.n3 0.189894
R2462 VN.n11 VN.n10 0.189894
R2463 VN.n12 VN.n11 0.189894
R2464 VN.n12 VN.n1 0.189894
R2465 VN.n16 VN.n1 0.189894
R2466 VDD2.n131 VDD2.n130 289.615
R2467 VDD2.n64 VDD2.n63 289.615
R2468 VDD2.n130 VDD2.n129 185
R2469 VDD2.n69 VDD2.n68 185
R2470 VDD2.n124 VDD2.n123 185
R2471 VDD2.n122 VDD2.n121 185
R2472 VDD2.n73 VDD2.n72 185
R2473 VDD2.n116 VDD2.n115 185
R2474 VDD2.n114 VDD2.n113 185
R2475 VDD2.n77 VDD2.n76 185
R2476 VDD2.n108 VDD2.n107 185
R2477 VDD2.n106 VDD2.n105 185
R2478 VDD2.n81 VDD2.n80 185
R2479 VDD2.n100 VDD2.n99 185
R2480 VDD2.n98 VDD2.n97 185
R2481 VDD2.n85 VDD2.n84 185
R2482 VDD2.n92 VDD2.n91 185
R2483 VDD2.n90 VDD2.n89 185
R2484 VDD2.n23 VDD2.n22 185
R2485 VDD2.n25 VDD2.n24 185
R2486 VDD2.n18 VDD2.n17 185
R2487 VDD2.n31 VDD2.n30 185
R2488 VDD2.n33 VDD2.n32 185
R2489 VDD2.n14 VDD2.n13 185
R2490 VDD2.n39 VDD2.n38 185
R2491 VDD2.n41 VDD2.n40 185
R2492 VDD2.n10 VDD2.n9 185
R2493 VDD2.n47 VDD2.n46 185
R2494 VDD2.n49 VDD2.n48 185
R2495 VDD2.n6 VDD2.n5 185
R2496 VDD2.n55 VDD2.n54 185
R2497 VDD2.n57 VDD2.n56 185
R2498 VDD2.n2 VDD2.n1 185
R2499 VDD2.n63 VDD2.n62 185
R2500 VDD2.n88 VDD2.t4 147.659
R2501 VDD2.n21 VDD2.t5 147.659
R2502 VDD2.n130 VDD2.n68 104.615
R2503 VDD2.n123 VDD2.n68 104.615
R2504 VDD2.n123 VDD2.n122 104.615
R2505 VDD2.n122 VDD2.n72 104.615
R2506 VDD2.n115 VDD2.n72 104.615
R2507 VDD2.n115 VDD2.n114 104.615
R2508 VDD2.n114 VDD2.n76 104.615
R2509 VDD2.n107 VDD2.n76 104.615
R2510 VDD2.n107 VDD2.n106 104.615
R2511 VDD2.n106 VDD2.n80 104.615
R2512 VDD2.n99 VDD2.n80 104.615
R2513 VDD2.n99 VDD2.n98 104.615
R2514 VDD2.n98 VDD2.n84 104.615
R2515 VDD2.n91 VDD2.n84 104.615
R2516 VDD2.n91 VDD2.n90 104.615
R2517 VDD2.n24 VDD2.n23 104.615
R2518 VDD2.n24 VDD2.n17 104.615
R2519 VDD2.n31 VDD2.n17 104.615
R2520 VDD2.n32 VDD2.n31 104.615
R2521 VDD2.n32 VDD2.n13 104.615
R2522 VDD2.n39 VDD2.n13 104.615
R2523 VDD2.n40 VDD2.n39 104.615
R2524 VDD2.n40 VDD2.n9 104.615
R2525 VDD2.n47 VDD2.n9 104.615
R2526 VDD2.n48 VDD2.n47 104.615
R2527 VDD2.n48 VDD2.n5 104.615
R2528 VDD2.n55 VDD2.n5 104.615
R2529 VDD2.n56 VDD2.n55 104.615
R2530 VDD2.n56 VDD2.n1 104.615
R2531 VDD2.n63 VDD2.n1 104.615
R2532 VDD2.n66 VDD2.n65 66.4742
R2533 VDD2 VDD2.n133 66.4705
R2534 VDD2.n66 VDD2.n64 54.4592
R2535 VDD2.n90 VDD2.t4 52.3082
R2536 VDD2.n23 VDD2.t5 52.3082
R2537 VDD2.n132 VDD2.n131 52.1611
R2538 VDD2.n132 VDD2.n66 44.2498
R2539 VDD2.n89 VDD2.n88 15.6677
R2540 VDD2.n22 VDD2.n21 15.6677
R2541 VDD2.n92 VDD2.n87 12.8005
R2542 VDD2.n25 VDD2.n20 12.8005
R2543 VDD2.n129 VDD2.n67 12.0247
R2544 VDD2.n93 VDD2.n85 12.0247
R2545 VDD2.n26 VDD2.n18 12.0247
R2546 VDD2.n62 VDD2.n0 12.0247
R2547 VDD2.n128 VDD2.n69 11.249
R2548 VDD2.n97 VDD2.n96 11.249
R2549 VDD2.n30 VDD2.n29 11.249
R2550 VDD2.n61 VDD2.n2 11.249
R2551 VDD2.n125 VDD2.n124 10.4732
R2552 VDD2.n100 VDD2.n83 10.4732
R2553 VDD2.n33 VDD2.n16 10.4732
R2554 VDD2.n58 VDD2.n57 10.4732
R2555 VDD2.n121 VDD2.n71 9.69747
R2556 VDD2.n101 VDD2.n81 9.69747
R2557 VDD2.n34 VDD2.n14 9.69747
R2558 VDD2.n54 VDD2.n4 9.69747
R2559 VDD2.n127 VDD2.n67 9.45567
R2560 VDD2.n60 VDD2.n0 9.45567
R2561 VDD2.n75 VDD2.n74 9.3005
R2562 VDD2.n118 VDD2.n117 9.3005
R2563 VDD2.n120 VDD2.n119 9.3005
R2564 VDD2.n71 VDD2.n70 9.3005
R2565 VDD2.n126 VDD2.n125 9.3005
R2566 VDD2.n128 VDD2.n127 9.3005
R2567 VDD2.n112 VDD2.n111 9.3005
R2568 VDD2.n110 VDD2.n109 9.3005
R2569 VDD2.n79 VDD2.n78 9.3005
R2570 VDD2.n104 VDD2.n103 9.3005
R2571 VDD2.n102 VDD2.n101 9.3005
R2572 VDD2.n83 VDD2.n82 9.3005
R2573 VDD2.n96 VDD2.n95 9.3005
R2574 VDD2.n94 VDD2.n93 9.3005
R2575 VDD2.n87 VDD2.n86 9.3005
R2576 VDD2.n45 VDD2.n44 9.3005
R2577 VDD2.n8 VDD2.n7 9.3005
R2578 VDD2.n51 VDD2.n50 9.3005
R2579 VDD2.n53 VDD2.n52 9.3005
R2580 VDD2.n4 VDD2.n3 9.3005
R2581 VDD2.n59 VDD2.n58 9.3005
R2582 VDD2.n61 VDD2.n60 9.3005
R2583 VDD2.n12 VDD2.n11 9.3005
R2584 VDD2.n37 VDD2.n36 9.3005
R2585 VDD2.n35 VDD2.n34 9.3005
R2586 VDD2.n16 VDD2.n15 9.3005
R2587 VDD2.n29 VDD2.n28 9.3005
R2588 VDD2.n27 VDD2.n26 9.3005
R2589 VDD2.n20 VDD2.n19 9.3005
R2590 VDD2.n43 VDD2.n42 9.3005
R2591 VDD2.n120 VDD2.n73 8.92171
R2592 VDD2.n105 VDD2.n104 8.92171
R2593 VDD2.n38 VDD2.n37 8.92171
R2594 VDD2.n53 VDD2.n6 8.92171
R2595 VDD2.n117 VDD2.n116 8.14595
R2596 VDD2.n108 VDD2.n79 8.14595
R2597 VDD2.n41 VDD2.n12 8.14595
R2598 VDD2.n50 VDD2.n49 8.14595
R2599 VDD2.n113 VDD2.n75 7.3702
R2600 VDD2.n109 VDD2.n77 7.3702
R2601 VDD2.n42 VDD2.n10 7.3702
R2602 VDD2.n46 VDD2.n8 7.3702
R2603 VDD2.n113 VDD2.n112 6.59444
R2604 VDD2.n112 VDD2.n77 6.59444
R2605 VDD2.n45 VDD2.n10 6.59444
R2606 VDD2.n46 VDD2.n45 6.59444
R2607 VDD2.n116 VDD2.n75 5.81868
R2608 VDD2.n109 VDD2.n108 5.81868
R2609 VDD2.n42 VDD2.n41 5.81868
R2610 VDD2.n49 VDD2.n8 5.81868
R2611 VDD2.n117 VDD2.n73 5.04292
R2612 VDD2.n105 VDD2.n79 5.04292
R2613 VDD2.n38 VDD2.n12 5.04292
R2614 VDD2.n50 VDD2.n6 5.04292
R2615 VDD2.n88 VDD2.n86 4.38563
R2616 VDD2.n21 VDD2.n19 4.38563
R2617 VDD2.n121 VDD2.n120 4.26717
R2618 VDD2.n104 VDD2.n81 4.26717
R2619 VDD2.n37 VDD2.n14 4.26717
R2620 VDD2.n54 VDD2.n53 4.26717
R2621 VDD2.n124 VDD2.n71 3.49141
R2622 VDD2.n101 VDD2.n100 3.49141
R2623 VDD2.n34 VDD2.n33 3.49141
R2624 VDD2.n57 VDD2.n4 3.49141
R2625 VDD2.n125 VDD2.n69 2.71565
R2626 VDD2.n97 VDD2.n83 2.71565
R2627 VDD2.n30 VDD2.n16 2.71565
R2628 VDD2.n58 VDD2.n2 2.71565
R2629 VDD2 VDD2.n132 2.41214
R2630 VDD2.n129 VDD2.n128 1.93989
R2631 VDD2.n96 VDD2.n85 1.93989
R2632 VDD2.n29 VDD2.n18 1.93989
R2633 VDD2.n62 VDD2.n61 1.93989
R2634 VDD2.n133 VDD2.t3 1.65188
R2635 VDD2.n133 VDD2.t1 1.65188
R2636 VDD2.n65 VDD2.t2 1.65188
R2637 VDD2.n65 VDD2.t0 1.65188
R2638 VDD2.n131 VDD2.n67 1.16414
R2639 VDD2.n93 VDD2.n92 1.16414
R2640 VDD2.n26 VDD2.n25 1.16414
R2641 VDD2.n64 VDD2.n0 1.16414
R2642 VDD2.n89 VDD2.n87 0.388379
R2643 VDD2.n22 VDD2.n20 0.388379
R2644 VDD2.n127 VDD2.n126 0.155672
R2645 VDD2.n126 VDD2.n70 0.155672
R2646 VDD2.n119 VDD2.n70 0.155672
R2647 VDD2.n119 VDD2.n118 0.155672
R2648 VDD2.n118 VDD2.n74 0.155672
R2649 VDD2.n111 VDD2.n74 0.155672
R2650 VDD2.n111 VDD2.n110 0.155672
R2651 VDD2.n110 VDD2.n78 0.155672
R2652 VDD2.n103 VDD2.n78 0.155672
R2653 VDD2.n103 VDD2.n102 0.155672
R2654 VDD2.n102 VDD2.n82 0.155672
R2655 VDD2.n95 VDD2.n82 0.155672
R2656 VDD2.n95 VDD2.n94 0.155672
R2657 VDD2.n94 VDD2.n86 0.155672
R2658 VDD2.n27 VDD2.n19 0.155672
R2659 VDD2.n28 VDD2.n27 0.155672
R2660 VDD2.n28 VDD2.n15 0.155672
R2661 VDD2.n35 VDD2.n15 0.155672
R2662 VDD2.n36 VDD2.n35 0.155672
R2663 VDD2.n36 VDD2.n11 0.155672
R2664 VDD2.n43 VDD2.n11 0.155672
R2665 VDD2.n44 VDD2.n43 0.155672
R2666 VDD2.n44 VDD2.n7 0.155672
R2667 VDD2.n51 VDD2.n7 0.155672
R2668 VDD2.n52 VDD2.n51 0.155672
R2669 VDD2.n52 VDD2.n3 0.155672
R2670 VDD2.n59 VDD2.n3 0.155672
R2671 VDD2.n60 VDD2.n59 0.155672
C0 VP VTAIL 7.34796f
C1 VP VDD2 0.518438f
C2 VP VDD1 7.36703f
C3 VTAIL VDD2 7.99395f
C4 VTAIL VDD1 7.93772f
C5 VDD1 VDD2 1.68334f
C6 VP VN 7.6127f
C7 VN VTAIL 7.333721f
C8 VN VDD2 7.00328f
C9 VN VDD1 0.151625f
C10 VDD2 B 6.515678f
C11 VDD1 B 6.688505f
C12 VTAIL B 8.266823f
C13 VN B 14.96641f
C14 VP B 13.663165f
C15 VDD2.n0 B 0.012057f
C16 VDD2.n1 B 0.027129f
C17 VDD2.n2 B 0.012153f
C18 VDD2.n3 B 0.02136f
C19 VDD2.n4 B 0.011478f
C20 VDD2.n5 B 0.027129f
C21 VDD2.n6 B 0.012153f
C22 VDD2.n7 B 0.02136f
C23 VDD2.n8 B 0.011478f
C24 VDD2.n9 B 0.027129f
C25 VDD2.n10 B 0.012153f
C26 VDD2.n11 B 0.02136f
C27 VDD2.n12 B 0.011478f
C28 VDD2.n13 B 0.027129f
C29 VDD2.n14 B 0.012153f
C30 VDD2.n15 B 0.02136f
C31 VDD2.n16 B 0.011478f
C32 VDD2.n17 B 0.027129f
C33 VDD2.n18 B 0.012153f
C34 VDD2.n19 B 1.09504f
C35 VDD2.n20 B 0.011478f
C36 VDD2.t5 B 0.044513f
C37 VDD2.n21 B 0.123193f
C38 VDD2.n22 B 0.016026f
C39 VDD2.n23 B 0.020347f
C40 VDD2.n24 B 0.027129f
C41 VDD2.n25 B 0.012153f
C42 VDD2.n26 B 0.011478f
C43 VDD2.n27 B 0.02136f
C44 VDD2.n28 B 0.02136f
C45 VDD2.n29 B 0.011478f
C46 VDD2.n30 B 0.012153f
C47 VDD2.n31 B 0.027129f
C48 VDD2.n32 B 0.027129f
C49 VDD2.n33 B 0.012153f
C50 VDD2.n34 B 0.011478f
C51 VDD2.n35 B 0.02136f
C52 VDD2.n36 B 0.02136f
C53 VDD2.n37 B 0.011478f
C54 VDD2.n38 B 0.012153f
C55 VDD2.n39 B 0.027129f
C56 VDD2.n40 B 0.027129f
C57 VDD2.n41 B 0.012153f
C58 VDD2.n42 B 0.011478f
C59 VDD2.n43 B 0.02136f
C60 VDD2.n44 B 0.02136f
C61 VDD2.n45 B 0.011478f
C62 VDD2.n46 B 0.012153f
C63 VDD2.n47 B 0.027129f
C64 VDD2.n48 B 0.027129f
C65 VDD2.n49 B 0.012153f
C66 VDD2.n50 B 0.011478f
C67 VDD2.n51 B 0.02136f
C68 VDD2.n52 B 0.02136f
C69 VDD2.n53 B 0.011478f
C70 VDD2.n54 B 0.012153f
C71 VDD2.n55 B 0.027129f
C72 VDD2.n56 B 0.027129f
C73 VDD2.n57 B 0.012153f
C74 VDD2.n58 B 0.011478f
C75 VDD2.n59 B 0.02136f
C76 VDD2.n60 B 0.056083f
C77 VDD2.n61 B 0.011478f
C78 VDD2.n62 B 0.012153f
C79 VDD2.n63 B 0.055417f
C80 VDD2.n64 B 0.070525f
C81 VDD2.t2 B 0.20238f
C82 VDD2.t0 B 0.20238f
C83 VDD2.n65 B 1.81729f
C84 VDD2.n66 B 2.54453f
C85 VDD2.n67 B 0.012057f
C86 VDD2.n68 B 0.027129f
C87 VDD2.n69 B 0.012153f
C88 VDD2.n70 B 0.02136f
C89 VDD2.n71 B 0.011478f
C90 VDD2.n72 B 0.027129f
C91 VDD2.n73 B 0.012153f
C92 VDD2.n74 B 0.02136f
C93 VDD2.n75 B 0.011478f
C94 VDD2.n76 B 0.027129f
C95 VDD2.n77 B 0.012153f
C96 VDD2.n78 B 0.02136f
C97 VDD2.n79 B 0.011478f
C98 VDD2.n80 B 0.027129f
C99 VDD2.n81 B 0.012153f
C100 VDD2.n82 B 0.02136f
C101 VDD2.n83 B 0.011478f
C102 VDD2.n84 B 0.027129f
C103 VDD2.n85 B 0.012153f
C104 VDD2.n86 B 1.09504f
C105 VDD2.n87 B 0.011478f
C106 VDD2.t4 B 0.044513f
C107 VDD2.n88 B 0.123193f
C108 VDD2.n89 B 0.016026f
C109 VDD2.n90 B 0.020347f
C110 VDD2.n91 B 0.027129f
C111 VDD2.n92 B 0.012153f
C112 VDD2.n93 B 0.011478f
C113 VDD2.n94 B 0.02136f
C114 VDD2.n95 B 0.02136f
C115 VDD2.n96 B 0.011478f
C116 VDD2.n97 B 0.012153f
C117 VDD2.n98 B 0.027129f
C118 VDD2.n99 B 0.027129f
C119 VDD2.n100 B 0.012153f
C120 VDD2.n101 B 0.011478f
C121 VDD2.n102 B 0.02136f
C122 VDD2.n103 B 0.02136f
C123 VDD2.n104 B 0.011478f
C124 VDD2.n105 B 0.012153f
C125 VDD2.n106 B 0.027129f
C126 VDD2.n107 B 0.027129f
C127 VDD2.n108 B 0.012153f
C128 VDD2.n109 B 0.011478f
C129 VDD2.n110 B 0.02136f
C130 VDD2.n111 B 0.02136f
C131 VDD2.n112 B 0.011478f
C132 VDD2.n113 B 0.012153f
C133 VDD2.n114 B 0.027129f
C134 VDD2.n115 B 0.027129f
C135 VDD2.n116 B 0.012153f
C136 VDD2.n117 B 0.011478f
C137 VDD2.n118 B 0.02136f
C138 VDD2.n119 B 0.02136f
C139 VDD2.n120 B 0.011478f
C140 VDD2.n121 B 0.012153f
C141 VDD2.n122 B 0.027129f
C142 VDD2.n123 B 0.027129f
C143 VDD2.n124 B 0.012153f
C144 VDD2.n125 B 0.011478f
C145 VDD2.n126 B 0.02136f
C146 VDD2.n127 B 0.056083f
C147 VDD2.n128 B 0.011478f
C148 VDD2.n129 B 0.012153f
C149 VDD2.n130 B 0.055417f
C150 VDD2.n131 B 0.061986f
C151 VDD2.n132 B 2.35634f
C152 VDD2.t3 B 0.20238f
C153 VDD2.t1 B 0.20238f
C154 VDD2.n133 B 1.81726f
C155 VN.t5 B 2.152f
C156 VN.n0 B 0.840642f
C157 VN.n1 B 0.019902f
C158 VN.n2 B 0.017378f
C159 VN.n3 B 0.019902f
C160 VN.t3 B 2.152f
C161 VN.n4 B 0.822621f
C162 VN.t0 B 2.40124f
C163 VN.n5 B 0.783407f
C164 VN.n6 B 0.232193f
C165 VN.n7 B 0.027936f
C166 VN.n8 B 0.037092f
C167 VN.n9 B 0.0402f
C168 VN.n10 B 0.019902f
C169 VN.n11 B 0.019902f
C170 VN.n12 B 0.019902f
C171 VN.n13 B 0.037621f
C172 VN.n14 B 0.037092f
C173 VN.n15 B 0.033064f
C174 VN.n16 B 0.032121f
C175 VN.n17 B 0.044349f
C176 VN.t1 B 2.152f
C177 VN.n18 B 0.840642f
C178 VN.n19 B 0.019902f
C179 VN.n20 B 0.017378f
C180 VN.n21 B 0.019902f
C181 VN.t2 B 2.152f
C182 VN.n22 B 0.822621f
C183 VN.t4 B 2.40124f
C184 VN.n23 B 0.783407f
C185 VN.n24 B 0.232193f
C186 VN.n25 B 0.027936f
C187 VN.n26 B 0.037092f
C188 VN.n27 B 0.0402f
C189 VN.n28 B 0.019902f
C190 VN.n29 B 0.019902f
C191 VN.n30 B 0.019902f
C192 VN.n31 B 0.037621f
C193 VN.n32 B 0.037092f
C194 VN.n33 B 0.033064f
C195 VN.n34 B 0.032121f
C196 VN.n35 B 1.19102f
C197 VDD1.n0 B 0.012234f
C198 VDD1.n1 B 0.027527f
C199 VDD1.n2 B 0.012331f
C200 VDD1.n3 B 0.021673f
C201 VDD1.n4 B 0.011646f
C202 VDD1.n5 B 0.027527f
C203 VDD1.n6 B 0.012331f
C204 VDD1.n7 B 0.021673f
C205 VDD1.n8 B 0.011646f
C206 VDD1.n9 B 0.027527f
C207 VDD1.n10 B 0.012331f
C208 VDD1.n11 B 0.021673f
C209 VDD1.n12 B 0.011646f
C210 VDD1.n13 B 0.027527f
C211 VDD1.n14 B 0.012331f
C212 VDD1.n15 B 0.021673f
C213 VDD1.n16 B 0.011646f
C214 VDD1.n17 B 0.027527f
C215 VDD1.n18 B 0.012331f
C216 VDD1.n19 B 1.11109f
C217 VDD1.n20 B 0.011646f
C218 VDD1.t0 B 0.045165f
C219 VDD1.n21 B 0.125f
C220 VDD1.n22 B 0.016261f
C221 VDD1.n23 B 0.020645f
C222 VDD1.n24 B 0.027527f
C223 VDD1.n25 B 0.012331f
C224 VDD1.n26 B 0.011646f
C225 VDD1.n27 B 0.021673f
C226 VDD1.n28 B 0.021673f
C227 VDD1.n29 B 0.011646f
C228 VDD1.n30 B 0.012331f
C229 VDD1.n31 B 0.027527f
C230 VDD1.n32 B 0.027527f
C231 VDD1.n33 B 0.012331f
C232 VDD1.n34 B 0.011646f
C233 VDD1.n35 B 0.021673f
C234 VDD1.n36 B 0.021673f
C235 VDD1.n37 B 0.011646f
C236 VDD1.n38 B 0.012331f
C237 VDD1.n39 B 0.027527f
C238 VDD1.n40 B 0.027527f
C239 VDD1.n41 B 0.012331f
C240 VDD1.n42 B 0.011646f
C241 VDD1.n43 B 0.021673f
C242 VDD1.n44 B 0.021673f
C243 VDD1.n45 B 0.011646f
C244 VDD1.n46 B 0.012331f
C245 VDD1.n47 B 0.027527f
C246 VDD1.n48 B 0.027527f
C247 VDD1.n49 B 0.012331f
C248 VDD1.n50 B 0.011646f
C249 VDD1.n51 B 0.021673f
C250 VDD1.n52 B 0.021673f
C251 VDD1.n53 B 0.011646f
C252 VDD1.n54 B 0.012331f
C253 VDD1.n55 B 0.027527f
C254 VDD1.n56 B 0.027527f
C255 VDD1.n57 B 0.012331f
C256 VDD1.n58 B 0.011646f
C257 VDD1.n59 B 0.021673f
C258 VDD1.n60 B 0.056906f
C259 VDD1.n61 B 0.011646f
C260 VDD1.n62 B 0.012331f
C261 VDD1.n63 B 0.05623f
C262 VDD1.n64 B 0.072309f
C263 VDD1.n65 B 0.012234f
C264 VDD1.n66 B 0.027527f
C265 VDD1.n67 B 0.012331f
C266 VDD1.n68 B 0.021673f
C267 VDD1.n69 B 0.011646f
C268 VDD1.n70 B 0.027527f
C269 VDD1.n71 B 0.012331f
C270 VDD1.n72 B 0.021673f
C271 VDD1.n73 B 0.011646f
C272 VDD1.n74 B 0.027527f
C273 VDD1.n75 B 0.012331f
C274 VDD1.n76 B 0.021673f
C275 VDD1.n77 B 0.011646f
C276 VDD1.n78 B 0.027527f
C277 VDD1.n79 B 0.012331f
C278 VDD1.n80 B 0.021673f
C279 VDD1.n81 B 0.011646f
C280 VDD1.n82 B 0.027527f
C281 VDD1.n83 B 0.012331f
C282 VDD1.n84 B 1.11109f
C283 VDD1.n85 B 0.011646f
C284 VDD1.t1 B 0.045165f
C285 VDD1.n86 B 0.125f
C286 VDD1.n87 B 0.016261f
C287 VDD1.n88 B 0.020645f
C288 VDD1.n89 B 0.027527f
C289 VDD1.n90 B 0.012331f
C290 VDD1.n91 B 0.011646f
C291 VDD1.n92 B 0.021673f
C292 VDD1.n93 B 0.021673f
C293 VDD1.n94 B 0.011646f
C294 VDD1.n95 B 0.012331f
C295 VDD1.n96 B 0.027527f
C296 VDD1.n97 B 0.027527f
C297 VDD1.n98 B 0.012331f
C298 VDD1.n99 B 0.011646f
C299 VDD1.n100 B 0.021673f
C300 VDD1.n101 B 0.021673f
C301 VDD1.n102 B 0.011646f
C302 VDD1.n103 B 0.012331f
C303 VDD1.n104 B 0.027527f
C304 VDD1.n105 B 0.027527f
C305 VDD1.n106 B 0.012331f
C306 VDD1.n107 B 0.011646f
C307 VDD1.n108 B 0.021673f
C308 VDD1.n109 B 0.021673f
C309 VDD1.n110 B 0.011646f
C310 VDD1.n111 B 0.012331f
C311 VDD1.n112 B 0.027527f
C312 VDD1.n113 B 0.027527f
C313 VDD1.n114 B 0.012331f
C314 VDD1.n115 B 0.011646f
C315 VDD1.n116 B 0.021673f
C316 VDD1.n117 B 0.021673f
C317 VDD1.n118 B 0.011646f
C318 VDD1.n119 B 0.012331f
C319 VDD1.n120 B 0.027527f
C320 VDD1.n121 B 0.027527f
C321 VDD1.n122 B 0.012331f
C322 VDD1.n123 B 0.011646f
C323 VDD1.n124 B 0.021673f
C324 VDD1.n125 B 0.056906f
C325 VDD1.n126 B 0.011646f
C326 VDD1.n127 B 0.012331f
C327 VDD1.n128 B 0.05623f
C328 VDD1.n129 B 0.07156f
C329 VDD1.t3 B 0.205348f
C330 VDD1.t4 B 0.205348f
C331 VDD1.n130 B 1.84394f
C332 VDD1.n131 B 2.70573f
C333 VDD1.t2 B 0.205348f
C334 VDD1.t5 B 0.205348f
C335 VDD1.n132 B 1.83901f
C336 VDD1.n133 B 2.58267f
C337 VTAIL.t2 B 0.228396f
C338 VTAIL.t0 B 0.228396f
C339 VTAIL.n0 B 1.98268f
C340 VTAIL.n1 B 0.442927f
C341 VTAIL.n2 B 0.013607f
C342 VTAIL.n3 B 0.030617f
C343 VTAIL.n4 B 0.013715f
C344 VTAIL.n5 B 0.024105f
C345 VTAIL.n6 B 0.012953f
C346 VTAIL.n7 B 0.030617f
C347 VTAIL.n8 B 0.013715f
C348 VTAIL.n9 B 0.024105f
C349 VTAIL.n10 B 0.012953f
C350 VTAIL.n11 B 0.030617f
C351 VTAIL.n12 B 0.013715f
C352 VTAIL.n13 B 0.024105f
C353 VTAIL.n14 B 0.012953f
C354 VTAIL.n15 B 0.030617f
C355 VTAIL.n16 B 0.013715f
C356 VTAIL.n17 B 0.024105f
C357 VTAIL.n18 B 0.012953f
C358 VTAIL.n19 B 0.030617f
C359 VTAIL.n20 B 0.013715f
C360 VTAIL.n21 B 1.2358f
C361 VTAIL.n22 B 0.012953f
C362 VTAIL.t6 B 0.050235f
C363 VTAIL.n23 B 0.13903f
C364 VTAIL.n24 B 0.018086f
C365 VTAIL.n25 B 0.022963f
C366 VTAIL.n26 B 0.030617f
C367 VTAIL.n27 B 0.013715f
C368 VTAIL.n28 B 0.012953f
C369 VTAIL.n29 B 0.024105f
C370 VTAIL.n30 B 0.024105f
C371 VTAIL.n31 B 0.012953f
C372 VTAIL.n32 B 0.013715f
C373 VTAIL.n33 B 0.030617f
C374 VTAIL.n34 B 0.030617f
C375 VTAIL.n35 B 0.013715f
C376 VTAIL.n36 B 0.012953f
C377 VTAIL.n37 B 0.024105f
C378 VTAIL.n38 B 0.024105f
C379 VTAIL.n39 B 0.012953f
C380 VTAIL.n40 B 0.013715f
C381 VTAIL.n41 B 0.030617f
C382 VTAIL.n42 B 0.030617f
C383 VTAIL.n43 B 0.013715f
C384 VTAIL.n44 B 0.012953f
C385 VTAIL.n45 B 0.024105f
C386 VTAIL.n46 B 0.024105f
C387 VTAIL.n47 B 0.012953f
C388 VTAIL.n48 B 0.013715f
C389 VTAIL.n49 B 0.030617f
C390 VTAIL.n50 B 0.030617f
C391 VTAIL.n51 B 0.013715f
C392 VTAIL.n52 B 0.012953f
C393 VTAIL.n53 B 0.024105f
C394 VTAIL.n54 B 0.024105f
C395 VTAIL.n55 B 0.012953f
C396 VTAIL.n56 B 0.013715f
C397 VTAIL.n57 B 0.030617f
C398 VTAIL.n58 B 0.030617f
C399 VTAIL.n59 B 0.013715f
C400 VTAIL.n60 B 0.012953f
C401 VTAIL.n61 B 0.024105f
C402 VTAIL.n62 B 0.063293f
C403 VTAIL.n63 B 0.012953f
C404 VTAIL.n64 B 0.013715f
C405 VTAIL.n65 B 0.062541f
C406 VTAIL.n66 B 0.05335f
C407 VTAIL.n67 B 0.425848f
C408 VTAIL.t8 B 0.228396f
C409 VTAIL.t9 B 0.228396f
C410 VTAIL.n68 B 1.98268f
C411 VTAIL.n69 B 2.08061f
C412 VTAIL.t10 B 0.228396f
C413 VTAIL.t1 B 0.228396f
C414 VTAIL.n70 B 1.98269f
C415 VTAIL.n71 B 2.0806f
C416 VTAIL.n72 B 0.013607f
C417 VTAIL.n73 B 0.030617f
C418 VTAIL.n74 B 0.013715f
C419 VTAIL.n75 B 0.024105f
C420 VTAIL.n76 B 0.012953f
C421 VTAIL.n77 B 0.030617f
C422 VTAIL.n78 B 0.013715f
C423 VTAIL.n79 B 0.024105f
C424 VTAIL.n80 B 0.012953f
C425 VTAIL.n81 B 0.030617f
C426 VTAIL.n82 B 0.013715f
C427 VTAIL.n83 B 0.024105f
C428 VTAIL.n84 B 0.012953f
C429 VTAIL.n85 B 0.030617f
C430 VTAIL.n86 B 0.013715f
C431 VTAIL.n87 B 0.024105f
C432 VTAIL.n88 B 0.012953f
C433 VTAIL.n89 B 0.030617f
C434 VTAIL.n90 B 0.013715f
C435 VTAIL.n91 B 1.2358f
C436 VTAIL.n92 B 0.012953f
C437 VTAIL.t3 B 0.050235f
C438 VTAIL.n93 B 0.13903f
C439 VTAIL.n94 B 0.018086f
C440 VTAIL.n95 B 0.022963f
C441 VTAIL.n96 B 0.030617f
C442 VTAIL.n97 B 0.013715f
C443 VTAIL.n98 B 0.012953f
C444 VTAIL.n99 B 0.024105f
C445 VTAIL.n100 B 0.024105f
C446 VTAIL.n101 B 0.012953f
C447 VTAIL.n102 B 0.013715f
C448 VTAIL.n103 B 0.030617f
C449 VTAIL.n104 B 0.030617f
C450 VTAIL.n105 B 0.013715f
C451 VTAIL.n106 B 0.012953f
C452 VTAIL.n107 B 0.024105f
C453 VTAIL.n108 B 0.024105f
C454 VTAIL.n109 B 0.012953f
C455 VTAIL.n110 B 0.013715f
C456 VTAIL.n111 B 0.030617f
C457 VTAIL.n112 B 0.030617f
C458 VTAIL.n113 B 0.013715f
C459 VTAIL.n114 B 0.012953f
C460 VTAIL.n115 B 0.024105f
C461 VTAIL.n116 B 0.024105f
C462 VTAIL.n117 B 0.012953f
C463 VTAIL.n118 B 0.013715f
C464 VTAIL.n119 B 0.030617f
C465 VTAIL.n120 B 0.030617f
C466 VTAIL.n121 B 0.013715f
C467 VTAIL.n122 B 0.012953f
C468 VTAIL.n123 B 0.024105f
C469 VTAIL.n124 B 0.024105f
C470 VTAIL.n125 B 0.012953f
C471 VTAIL.n126 B 0.013715f
C472 VTAIL.n127 B 0.030617f
C473 VTAIL.n128 B 0.030617f
C474 VTAIL.n129 B 0.013715f
C475 VTAIL.n130 B 0.012953f
C476 VTAIL.n131 B 0.024105f
C477 VTAIL.n132 B 0.063293f
C478 VTAIL.n133 B 0.012953f
C479 VTAIL.n134 B 0.013715f
C480 VTAIL.n135 B 0.062541f
C481 VTAIL.n136 B 0.05335f
C482 VTAIL.n137 B 0.425848f
C483 VTAIL.t4 B 0.228396f
C484 VTAIL.t5 B 0.228396f
C485 VTAIL.n138 B 1.98269f
C486 VTAIL.n139 B 0.621201f
C487 VTAIL.n140 B 0.013607f
C488 VTAIL.n141 B 0.030617f
C489 VTAIL.n142 B 0.013715f
C490 VTAIL.n143 B 0.024105f
C491 VTAIL.n144 B 0.012953f
C492 VTAIL.n145 B 0.030617f
C493 VTAIL.n146 B 0.013715f
C494 VTAIL.n147 B 0.024105f
C495 VTAIL.n148 B 0.012953f
C496 VTAIL.n149 B 0.030617f
C497 VTAIL.n150 B 0.013715f
C498 VTAIL.n151 B 0.024105f
C499 VTAIL.n152 B 0.012953f
C500 VTAIL.n153 B 0.030617f
C501 VTAIL.n154 B 0.013715f
C502 VTAIL.n155 B 0.024105f
C503 VTAIL.n156 B 0.012953f
C504 VTAIL.n157 B 0.030617f
C505 VTAIL.n158 B 0.013715f
C506 VTAIL.n159 B 1.2358f
C507 VTAIL.n160 B 0.012953f
C508 VTAIL.t7 B 0.050235f
C509 VTAIL.n161 B 0.13903f
C510 VTAIL.n162 B 0.018086f
C511 VTAIL.n163 B 0.022963f
C512 VTAIL.n164 B 0.030617f
C513 VTAIL.n165 B 0.013715f
C514 VTAIL.n166 B 0.012953f
C515 VTAIL.n167 B 0.024105f
C516 VTAIL.n168 B 0.024105f
C517 VTAIL.n169 B 0.012953f
C518 VTAIL.n170 B 0.013715f
C519 VTAIL.n171 B 0.030617f
C520 VTAIL.n172 B 0.030617f
C521 VTAIL.n173 B 0.013715f
C522 VTAIL.n174 B 0.012953f
C523 VTAIL.n175 B 0.024105f
C524 VTAIL.n176 B 0.024105f
C525 VTAIL.n177 B 0.012953f
C526 VTAIL.n178 B 0.013715f
C527 VTAIL.n179 B 0.030617f
C528 VTAIL.n180 B 0.030617f
C529 VTAIL.n181 B 0.013715f
C530 VTAIL.n182 B 0.012953f
C531 VTAIL.n183 B 0.024105f
C532 VTAIL.n184 B 0.024105f
C533 VTAIL.n185 B 0.012953f
C534 VTAIL.n186 B 0.013715f
C535 VTAIL.n187 B 0.030617f
C536 VTAIL.n188 B 0.030617f
C537 VTAIL.n189 B 0.013715f
C538 VTAIL.n190 B 0.012953f
C539 VTAIL.n191 B 0.024105f
C540 VTAIL.n192 B 0.024105f
C541 VTAIL.n193 B 0.012953f
C542 VTAIL.n194 B 0.013715f
C543 VTAIL.n195 B 0.030617f
C544 VTAIL.n196 B 0.030617f
C545 VTAIL.n197 B 0.013715f
C546 VTAIL.n198 B 0.012953f
C547 VTAIL.n199 B 0.024105f
C548 VTAIL.n200 B 0.063293f
C549 VTAIL.n201 B 0.012953f
C550 VTAIL.n202 B 0.013715f
C551 VTAIL.n203 B 0.062541f
C552 VTAIL.n204 B 0.05335f
C553 VTAIL.n205 B 1.64151f
C554 VTAIL.n206 B 0.013607f
C555 VTAIL.n207 B 0.030617f
C556 VTAIL.n208 B 0.013715f
C557 VTAIL.n209 B 0.024105f
C558 VTAIL.n210 B 0.012953f
C559 VTAIL.n211 B 0.030617f
C560 VTAIL.n212 B 0.013715f
C561 VTAIL.n213 B 0.024105f
C562 VTAIL.n214 B 0.012953f
C563 VTAIL.n215 B 0.030617f
C564 VTAIL.n216 B 0.013715f
C565 VTAIL.n217 B 0.024105f
C566 VTAIL.n218 B 0.012953f
C567 VTAIL.n219 B 0.030617f
C568 VTAIL.n220 B 0.013715f
C569 VTAIL.n221 B 0.024105f
C570 VTAIL.n222 B 0.012953f
C571 VTAIL.n223 B 0.030617f
C572 VTAIL.n224 B 0.013715f
C573 VTAIL.n225 B 1.2358f
C574 VTAIL.n226 B 0.012953f
C575 VTAIL.t11 B 0.050235f
C576 VTAIL.n227 B 0.13903f
C577 VTAIL.n228 B 0.018086f
C578 VTAIL.n229 B 0.022963f
C579 VTAIL.n230 B 0.030617f
C580 VTAIL.n231 B 0.013715f
C581 VTAIL.n232 B 0.012953f
C582 VTAIL.n233 B 0.024105f
C583 VTAIL.n234 B 0.024105f
C584 VTAIL.n235 B 0.012953f
C585 VTAIL.n236 B 0.013715f
C586 VTAIL.n237 B 0.030617f
C587 VTAIL.n238 B 0.030617f
C588 VTAIL.n239 B 0.013715f
C589 VTAIL.n240 B 0.012953f
C590 VTAIL.n241 B 0.024105f
C591 VTAIL.n242 B 0.024105f
C592 VTAIL.n243 B 0.012953f
C593 VTAIL.n244 B 0.013715f
C594 VTAIL.n245 B 0.030617f
C595 VTAIL.n246 B 0.030617f
C596 VTAIL.n247 B 0.013715f
C597 VTAIL.n248 B 0.012953f
C598 VTAIL.n249 B 0.024105f
C599 VTAIL.n250 B 0.024105f
C600 VTAIL.n251 B 0.012953f
C601 VTAIL.n252 B 0.013715f
C602 VTAIL.n253 B 0.030617f
C603 VTAIL.n254 B 0.030617f
C604 VTAIL.n255 B 0.013715f
C605 VTAIL.n256 B 0.012953f
C606 VTAIL.n257 B 0.024105f
C607 VTAIL.n258 B 0.024105f
C608 VTAIL.n259 B 0.012953f
C609 VTAIL.n260 B 0.013715f
C610 VTAIL.n261 B 0.030617f
C611 VTAIL.n262 B 0.030617f
C612 VTAIL.n263 B 0.013715f
C613 VTAIL.n264 B 0.012953f
C614 VTAIL.n265 B 0.024105f
C615 VTAIL.n266 B 0.063293f
C616 VTAIL.n267 B 0.012953f
C617 VTAIL.n268 B 0.013715f
C618 VTAIL.n269 B 0.062541f
C619 VTAIL.n270 B 0.05335f
C620 VTAIL.n271 B 1.57606f
C621 VP.t1 B 2.1941f
C622 VP.n0 B 0.857091f
C623 VP.n1 B 0.020291f
C624 VP.n2 B 0.017718f
C625 VP.n3 B 0.020291f
C626 VP.t2 B 2.1941f
C627 VP.n4 B 0.770953f
C628 VP.n5 B 0.020291f
C629 VP.n6 B 0.017718f
C630 VP.n7 B 0.020291f
C631 VP.t4 B 2.1941f
C632 VP.n8 B 0.857091f
C633 VP.t0 B 2.1941f
C634 VP.n9 B 0.857091f
C635 VP.n10 B 0.020291f
C636 VP.n11 B 0.017718f
C637 VP.n12 B 0.020291f
C638 VP.t3 B 2.1941f
C639 VP.n13 B 0.838718f
C640 VP.t5 B 2.44822f
C641 VP.n14 B 0.798737f
C642 VP.n15 B 0.236737f
C643 VP.n16 B 0.028483f
C644 VP.n17 B 0.037818f
C645 VP.n18 B 0.040987f
C646 VP.n19 B 0.020291f
C647 VP.n20 B 0.020291f
C648 VP.n21 B 0.020291f
C649 VP.n22 B 0.038357f
C650 VP.n23 B 0.037818f
C651 VP.n24 B 0.033711f
C652 VP.n25 B 0.03275f
C653 VP.n26 B 1.20612f
C654 VP.n27 B 1.22025f
C655 VP.n28 B 0.03275f
C656 VP.n29 B 0.033711f
C657 VP.n30 B 0.037818f
C658 VP.n31 B 0.038357f
C659 VP.n32 B 0.020291f
C660 VP.n33 B 0.020291f
C661 VP.n34 B 0.020291f
C662 VP.n35 B 0.040987f
C663 VP.n36 B 0.037818f
C664 VP.n37 B 0.028483f
C665 VP.n38 B 0.020291f
C666 VP.n39 B 0.020291f
C667 VP.n40 B 0.028483f
C668 VP.n41 B 0.037818f
C669 VP.n42 B 0.040987f
C670 VP.n43 B 0.020291f
C671 VP.n44 B 0.020291f
C672 VP.n45 B 0.020291f
C673 VP.n46 B 0.038357f
C674 VP.n47 B 0.037818f
C675 VP.n48 B 0.033711f
C676 VP.n49 B 0.03275f
C677 VP.n50 B 0.045217f
.ends

