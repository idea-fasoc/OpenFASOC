* NGSPICE file created from diff_pair_sample_1390.ext - technology: sky130A

.subckt diff_pair_sample_1390 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X1 VDD2.t8 VN.t1 VTAIL.t15 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X2 VTAIL.t5 VP.t0 VDD1.t9 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X3 VTAIL.t14 VN.t2 VDD2.t7 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X4 VTAIL.t13 VN.t3 VDD2.t6 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X5 VDD1.t8 VP.t1 VTAIL.t3 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X6 VDD2.t5 VN.t4 VTAIL.t10 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=1.0923 ps=6.95 w=6.62 l=3.28
X7 B.t11 B.t9 B.t10 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=0 ps=0 w=6.62 l=3.28
X8 VTAIL.t17 VP.t2 VDD1.t7 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X9 VDD1.t6 VP.t3 VTAIL.t18 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=1.0923 ps=6.95 w=6.62 l=3.28
X10 VTAIL.t11 VN.t5 VDD2.t4 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X11 VDD2.t3 VN.t6 VTAIL.t16 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=2.5818 ps=14.02 w=6.62 l=3.28
X12 VTAIL.t1 VP.t4 VDD1.t5 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X13 B.t8 B.t6 B.t7 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=0 ps=0 w=6.62 l=3.28
X14 VDD2.t2 VN.t7 VTAIL.t7 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=2.5818 ps=14.02 w=6.62 l=3.28
X15 VDD2.t1 VN.t8 VTAIL.t8 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=1.0923 ps=6.95 w=6.62 l=3.28
X16 VDD1.t4 VP.t5 VTAIL.t0 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=1.0923 ps=6.95 w=6.62 l=3.28
X17 VDD1.t3 VP.t6 VTAIL.t2 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X18 VTAIL.t19 VP.t7 VDD1.t2 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X19 VTAIL.t9 VN.t9 VDD2.t0 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=1.0923 ps=6.95 w=6.62 l=3.28
X20 VDD1.t1 VP.t8 VTAIL.t4 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=2.5818 ps=14.02 w=6.62 l=3.28
X21 B.t5 B.t3 B.t4 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=0 ps=0 w=6.62 l=3.28
X22 VDD1.t0 VP.t9 VTAIL.t6 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=1.0923 pd=6.95 as=2.5818 ps=14.02 w=6.62 l=3.28
X23 B.t2 B.t0 B.t1 w_n5302_n2292# sky130_fd_pr__pfet_01v8 ad=2.5818 pd=14.02 as=0 ps=0 w=6.62 l=3.28
R0 VN.n96 VN.n95 161.3
R1 VN.n94 VN.n50 161.3
R2 VN.n93 VN.n92 161.3
R3 VN.n91 VN.n51 161.3
R4 VN.n90 VN.n89 161.3
R5 VN.n88 VN.n52 161.3
R6 VN.n87 VN.n86 161.3
R7 VN.n85 VN.n84 161.3
R8 VN.n83 VN.n54 161.3
R9 VN.n82 VN.n81 161.3
R10 VN.n80 VN.n55 161.3
R11 VN.n79 VN.n78 161.3
R12 VN.n77 VN.n56 161.3
R13 VN.n76 VN.n75 161.3
R14 VN.n74 VN.n57 161.3
R15 VN.n73 VN.n72 161.3
R16 VN.n71 VN.n58 161.3
R17 VN.n70 VN.n69 161.3
R18 VN.n68 VN.n59 161.3
R19 VN.n67 VN.n66 161.3
R20 VN.n65 VN.n60 161.3
R21 VN.n64 VN.n63 161.3
R22 VN.n47 VN.n46 161.3
R23 VN.n45 VN.n1 161.3
R24 VN.n44 VN.n43 161.3
R25 VN.n42 VN.n2 161.3
R26 VN.n41 VN.n40 161.3
R27 VN.n39 VN.n3 161.3
R28 VN.n38 VN.n37 161.3
R29 VN.n36 VN.n35 161.3
R30 VN.n34 VN.n5 161.3
R31 VN.n33 VN.n32 161.3
R32 VN.n31 VN.n6 161.3
R33 VN.n30 VN.n29 161.3
R34 VN.n28 VN.n7 161.3
R35 VN.n27 VN.n26 161.3
R36 VN.n25 VN.n8 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n13 VN.t8 81.0196
R45 VN.n62 VN.t6 81.0196
R46 VN.n48 VN.n0 79.4252
R47 VN.n97 VN.n49 79.4252
R48 VN.n13 VN.n12 69.3368
R49 VN.n62 VN.n61 69.3368
R50 VN.n21 VN.n10 56.5617
R51 VN.n29 VN.n6 56.5617
R52 VN.n70 VN.n59 56.5617
R53 VN.n78 VN.n55 56.5617
R54 VN VN.n97 52.9489
R55 VN.n40 VN.n2 48.8116
R56 VN.n89 VN.n51 48.8116
R57 VN.n8 VN.t1 48.6414
R58 VN.n12 VN.t2 48.6414
R59 VN.n4 VN.t5 48.6414
R60 VN.n0 VN.t7 48.6414
R61 VN.n57 VN.t0 48.6414
R62 VN.n61 VN.t3 48.6414
R63 VN.n53 VN.t9 48.6414
R64 VN.n49 VN.t4 48.6414
R65 VN.n44 VN.n2 32.3425
R66 VN.n93 VN.n51 32.3425
R67 VN.n16 VN.n15 24.5923
R68 VN.n17 VN.n16 24.5923
R69 VN.n17 VN.n10 24.5923
R70 VN.n22 VN.n21 24.5923
R71 VN.n23 VN.n22 24.5923
R72 VN.n23 VN.n8 24.5923
R73 VN.n27 VN.n8 24.5923
R74 VN.n28 VN.n27 24.5923
R75 VN.n29 VN.n28 24.5923
R76 VN.n33 VN.n6 24.5923
R77 VN.n34 VN.n33 24.5923
R78 VN.n35 VN.n34 24.5923
R79 VN.n39 VN.n38 24.5923
R80 VN.n40 VN.n39 24.5923
R81 VN.n45 VN.n44 24.5923
R82 VN.n46 VN.n45 24.5923
R83 VN.n66 VN.n59 24.5923
R84 VN.n66 VN.n65 24.5923
R85 VN.n65 VN.n64 24.5923
R86 VN.n78 VN.n77 24.5923
R87 VN.n77 VN.n76 24.5923
R88 VN.n76 VN.n57 24.5923
R89 VN.n72 VN.n57 24.5923
R90 VN.n72 VN.n71 24.5923
R91 VN.n71 VN.n70 24.5923
R92 VN.n89 VN.n88 24.5923
R93 VN.n88 VN.n87 24.5923
R94 VN.n84 VN.n83 24.5923
R95 VN.n83 VN.n82 24.5923
R96 VN.n82 VN.n55 24.5923
R97 VN.n95 VN.n94 24.5923
R98 VN.n94 VN.n93 24.5923
R99 VN.n38 VN.n4 19.1821
R100 VN.n87 VN.n53 19.1821
R101 VN.n46 VN.n0 10.8209
R102 VN.n95 VN.n49 10.8209
R103 VN.n15 VN.n12 5.4107
R104 VN.n35 VN.n4 5.4107
R105 VN.n64 VN.n61 5.4107
R106 VN.n84 VN.n53 5.4107
R107 VN.n14 VN.n13 4.34643
R108 VN.n63 VN.n62 4.34643
R109 VN.n97 VN.n96 0.354861
R110 VN.n48 VN.n47 0.354861
R111 VN VN.n48 0.267071
R112 VN.n96 VN.n50 0.189894
R113 VN.n92 VN.n50 0.189894
R114 VN.n92 VN.n91 0.189894
R115 VN.n91 VN.n90 0.189894
R116 VN.n90 VN.n52 0.189894
R117 VN.n86 VN.n52 0.189894
R118 VN.n86 VN.n85 0.189894
R119 VN.n85 VN.n54 0.189894
R120 VN.n81 VN.n54 0.189894
R121 VN.n81 VN.n80 0.189894
R122 VN.n80 VN.n79 0.189894
R123 VN.n79 VN.n56 0.189894
R124 VN.n75 VN.n56 0.189894
R125 VN.n75 VN.n74 0.189894
R126 VN.n74 VN.n73 0.189894
R127 VN.n73 VN.n58 0.189894
R128 VN.n69 VN.n58 0.189894
R129 VN.n69 VN.n68 0.189894
R130 VN.n68 VN.n67 0.189894
R131 VN.n67 VN.n60 0.189894
R132 VN.n63 VN.n60 0.189894
R133 VN.n14 VN.n11 0.189894
R134 VN.n18 VN.n11 0.189894
R135 VN.n19 VN.n18 0.189894
R136 VN.n20 VN.n19 0.189894
R137 VN.n20 VN.n9 0.189894
R138 VN.n24 VN.n9 0.189894
R139 VN.n25 VN.n24 0.189894
R140 VN.n26 VN.n25 0.189894
R141 VN.n26 VN.n7 0.189894
R142 VN.n30 VN.n7 0.189894
R143 VN.n31 VN.n30 0.189894
R144 VN.n32 VN.n31 0.189894
R145 VN.n32 VN.n5 0.189894
R146 VN.n36 VN.n5 0.189894
R147 VN.n37 VN.n36 0.189894
R148 VN.n37 VN.n3 0.189894
R149 VN.n41 VN.n3 0.189894
R150 VN.n42 VN.n41 0.189894
R151 VN.n43 VN.n42 0.189894
R152 VN.n43 VN.n1 0.189894
R153 VN.n47 VN.n1 0.189894
R154 VTAIL.n152 VTAIL.n122 756.745
R155 VTAIL.n32 VTAIL.n2 756.745
R156 VTAIL.n116 VTAIL.n86 756.745
R157 VTAIL.n76 VTAIL.n46 756.745
R158 VTAIL.n135 VTAIL.n134 585
R159 VTAIL.n137 VTAIL.n136 585
R160 VTAIL.n130 VTAIL.n129 585
R161 VTAIL.n143 VTAIL.n142 585
R162 VTAIL.n145 VTAIL.n144 585
R163 VTAIL.n126 VTAIL.n125 585
R164 VTAIL.n151 VTAIL.n150 585
R165 VTAIL.n153 VTAIL.n152 585
R166 VTAIL.n15 VTAIL.n14 585
R167 VTAIL.n17 VTAIL.n16 585
R168 VTAIL.n10 VTAIL.n9 585
R169 VTAIL.n23 VTAIL.n22 585
R170 VTAIL.n25 VTAIL.n24 585
R171 VTAIL.n6 VTAIL.n5 585
R172 VTAIL.n31 VTAIL.n30 585
R173 VTAIL.n33 VTAIL.n32 585
R174 VTAIL.n117 VTAIL.n116 585
R175 VTAIL.n115 VTAIL.n114 585
R176 VTAIL.n90 VTAIL.n89 585
R177 VTAIL.n109 VTAIL.n108 585
R178 VTAIL.n107 VTAIL.n106 585
R179 VTAIL.n94 VTAIL.n93 585
R180 VTAIL.n101 VTAIL.n100 585
R181 VTAIL.n99 VTAIL.n98 585
R182 VTAIL.n77 VTAIL.n76 585
R183 VTAIL.n75 VTAIL.n74 585
R184 VTAIL.n50 VTAIL.n49 585
R185 VTAIL.n69 VTAIL.n68 585
R186 VTAIL.n67 VTAIL.n66 585
R187 VTAIL.n54 VTAIL.n53 585
R188 VTAIL.n61 VTAIL.n60 585
R189 VTAIL.n59 VTAIL.n58 585
R190 VTAIL.n133 VTAIL.t7 327.514
R191 VTAIL.n13 VTAIL.t4 327.514
R192 VTAIL.n97 VTAIL.t6 327.514
R193 VTAIL.n57 VTAIL.t16 327.514
R194 VTAIL.n136 VTAIL.n135 171.744
R195 VTAIL.n136 VTAIL.n129 171.744
R196 VTAIL.n143 VTAIL.n129 171.744
R197 VTAIL.n144 VTAIL.n143 171.744
R198 VTAIL.n144 VTAIL.n125 171.744
R199 VTAIL.n151 VTAIL.n125 171.744
R200 VTAIL.n152 VTAIL.n151 171.744
R201 VTAIL.n16 VTAIL.n15 171.744
R202 VTAIL.n16 VTAIL.n9 171.744
R203 VTAIL.n23 VTAIL.n9 171.744
R204 VTAIL.n24 VTAIL.n23 171.744
R205 VTAIL.n24 VTAIL.n5 171.744
R206 VTAIL.n31 VTAIL.n5 171.744
R207 VTAIL.n32 VTAIL.n31 171.744
R208 VTAIL.n116 VTAIL.n115 171.744
R209 VTAIL.n115 VTAIL.n89 171.744
R210 VTAIL.n108 VTAIL.n89 171.744
R211 VTAIL.n108 VTAIL.n107 171.744
R212 VTAIL.n107 VTAIL.n93 171.744
R213 VTAIL.n100 VTAIL.n93 171.744
R214 VTAIL.n100 VTAIL.n99 171.744
R215 VTAIL.n76 VTAIL.n75 171.744
R216 VTAIL.n75 VTAIL.n49 171.744
R217 VTAIL.n68 VTAIL.n49 171.744
R218 VTAIL.n68 VTAIL.n67 171.744
R219 VTAIL.n67 VTAIL.n53 171.744
R220 VTAIL.n60 VTAIL.n53 171.744
R221 VTAIL.n60 VTAIL.n59 171.744
R222 VTAIL.n135 VTAIL.t7 85.8723
R223 VTAIL.n15 VTAIL.t4 85.8723
R224 VTAIL.n99 VTAIL.t6 85.8723
R225 VTAIL.n59 VTAIL.t16 85.8723
R226 VTAIL.n85 VTAIL.n84 69.7808
R227 VTAIL.n83 VTAIL.n82 69.7808
R228 VTAIL.n45 VTAIL.n44 69.7808
R229 VTAIL.n43 VTAIL.n42 69.7808
R230 VTAIL.n159 VTAIL.n158 69.7806
R231 VTAIL.n1 VTAIL.n0 69.7806
R232 VTAIL.n39 VTAIL.n38 69.7806
R233 VTAIL.n41 VTAIL.n40 69.7806
R234 VTAIL.n157 VTAIL.n156 30.246
R235 VTAIL.n37 VTAIL.n36 30.246
R236 VTAIL.n121 VTAIL.n120 30.246
R237 VTAIL.n81 VTAIL.n80 30.246
R238 VTAIL.n43 VTAIL.n41 24.2979
R239 VTAIL.n157 VTAIL.n121 21.1858
R240 VTAIL.n134 VTAIL.n133 16.3884
R241 VTAIL.n14 VTAIL.n13 16.3884
R242 VTAIL.n98 VTAIL.n97 16.3884
R243 VTAIL.n58 VTAIL.n57 16.3884
R244 VTAIL.n137 VTAIL.n132 12.8005
R245 VTAIL.n17 VTAIL.n12 12.8005
R246 VTAIL.n101 VTAIL.n96 12.8005
R247 VTAIL.n61 VTAIL.n56 12.8005
R248 VTAIL.n138 VTAIL.n130 12.0247
R249 VTAIL.n18 VTAIL.n10 12.0247
R250 VTAIL.n102 VTAIL.n94 12.0247
R251 VTAIL.n62 VTAIL.n54 12.0247
R252 VTAIL.n142 VTAIL.n141 11.249
R253 VTAIL.n22 VTAIL.n21 11.249
R254 VTAIL.n106 VTAIL.n105 11.249
R255 VTAIL.n66 VTAIL.n65 11.249
R256 VTAIL.n145 VTAIL.n128 10.4732
R257 VTAIL.n25 VTAIL.n8 10.4732
R258 VTAIL.n109 VTAIL.n92 10.4732
R259 VTAIL.n69 VTAIL.n52 10.4732
R260 VTAIL.n146 VTAIL.n126 9.69747
R261 VTAIL.n26 VTAIL.n6 9.69747
R262 VTAIL.n110 VTAIL.n90 9.69747
R263 VTAIL.n70 VTAIL.n50 9.69747
R264 VTAIL.n156 VTAIL.n155 9.45567
R265 VTAIL.n36 VTAIL.n35 9.45567
R266 VTAIL.n120 VTAIL.n119 9.45567
R267 VTAIL.n80 VTAIL.n79 9.45567
R268 VTAIL.n124 VTAIL.n123 9.3005
R269 VTAIL.n149 VTAIL.n148 9.3005
R270 VTAIL.n147 VTAIL.n146 9.3005
R271 VTAIL.n128 VTAIL.n127 9.3005
R272 VTAIL.n141 VTAIL.n140 9.3005
R273 VTAIL.n139 VTAIL.n138 9.3005
R274 VTAIL.n132 VTAIL.n131 9.3005
R275 VTAIL.n155 VTAIL.n154 9.3005
R276 VTAIL.n4 VTAIL.n3 9.3005
R277 VTAIL.n29 VTAIL.n28 9.3005
R278 VTAIL.n27 VTAIL.n26 9.3005
R279 VTAIL.n8 VTAIL.n7 9.3005
R280 VTAIL.n21 VTAIL.n20 9.3005
R281 VTAIL.n19 VTAIL.n18 9.3005
R282 VTAIL.n12 VTAIL.n11 9.3005
R283 VTAIL.n35 VTAIL.n34 9.3005
R284 VTAIL.n119 VTAIL.n118 9.3005
R285 VTAIL.n88 VTAIL.n87 9.3005
R286 VTAIL.n113 VTAIL.n112 9.3005
R287 VTAIL.n111 VTAIL.n110 9.3005
R288 VTAIL.n92 VTAIL.n91 9.3005
R289 VTAIL.n105 VTAIL.n104 9.3005
R290 VTAIL.n103 VTAIL.n102 9.3005
R291 VTAIL.n96 VTAIL.n95 9.3005
R292 VTAIL.n79 VTAIL.n78 9.3005
R293 VTAIL.n48 VTAIL.n47 9.3005
R294 VTAIL.n73 VTAIL.n72 9.3005
R295 VTAIL.n71 VTAIL.n70 9.3005
R296 VTAIL.n52 VTAIL.n51 9.3005
R297 VTAIL.n65 VTAIL.n64 9.3005
R298 VTAIL.n63 VTAIL.n62 9.3005
R299 VTAIL.n56 VTAIL.n55 9.3005
R300 VTAIL.n150 VTAIL.n149 8.92171
R301 VTAIL.n30 VTAIL.n29 8.92171
R302 VTAIL.n114 VTAIL.n113 8.92171
R303 VTAIL.n74 VTAIL.n73 8.92171
R304 VTAIL.n153 VTAIL.n124 8.14595
R305 VTAIL.n33 VTAIL.n4 8.14595
R306 VTAIL.n117 VTAIL.n88 8.14595
R307 VTAIL.n77 VTAIL.n48 8.14595
R308 VTAIL.n154 VTAIL.n122 7.3702
R309 VTAIL.n34 VTAIL.n2 7.3702
R310 VTAIL.n118 VTAIL.n86 7.3702
R311 VTAIL.n78 VTAIL.n46 7.3702
R312 VTAIL.n156 VTAIL.n122 6.59444
R313 VTAIL.n36 VTAIL.n2 6.59444
R314 VTAIL.n120 VTAIL.n86 6.59444
R315 VTAIL.n80 VTAIL.n46 6.59444
R316 VTAIL.n154 VTAIL.n153 5.81868
R317 VTAIL.n34 VTAIL.n33 5.81868
R318 VTAIL.n118 VTAIL.n117 5.81868
R319 VTAIL.n78 VTAIL.n77 5.81868
R320 VTAIL.n150 VTAIL.n124 5.04292
R321 VTAIL.n30 VTAIL.n4 5.04292
R322 VTAIL.n114 VTAIL.n88 5.04292
R323 VTAIL.n74 VTAIL.n48 5.04292
R324 VTAIL.n158 VTAIL.t15 4.91062
R325 VTAIL.n158 VTAIL.t11 4.91062
R326 VTAIL.n0 VTAIL.t8 4.91062
R327 VTAIL.n0 VTAIL.t14 4.91062
R328 VTAIL.n38 VTAIL.t3 4.91062
R329 VTAIL.n38 VTAIL.t5 4.91062
R330 VTAIL.n40 VTAIL.t0 4.91062
R331 VTAIL.n40 VTAIL.t19 4.91062
R332 VTAIL.n84 VTAIL.t2 4.91062
R333 VTAIL.n84 VTAIL.t1 4.91062
R334 VTAIL.n82 VTAIL.t18 4.91062
R335 VTAIL.n82 VTAIL.t17 4.91062
R336 VTAIL.n44 VTAIL.t12 4.91062
R337 VTAIL.n44 VTAIL.t13 4.91062
R338 VTAIL.n42 VTAIL.t10 4.91062
R339 VTAIL.n42 VTAIL.t9 4.91062
R340 VTAIL.n149 VTAIL.n126 4.26717
R341 VTAIL.n29 VTAIL.n6 4.26717
R342 VTAIL.n113 VTAIL.n90 4.26717
R343 VTAIL.n73 VTAIL.n50 4.26717
R344 VTAIL.n133 VTAIL.n131 3.71088
R345 VTAIL.n13 VTAIL.n11 3.71088
R346 VTAIL.n97 VTAIL.n95 3.71088
R347 VTAIL.n57 VTAIL.n55 3.71088
R348 VTAIL.n146 VTAIL.n145 3.49141
R349 VTAIL.n26 VTAIL.n25 3.49141
R350 VTAIL.n110 VTAIL.n109 3.49141
R351 VTAIL.n70 VTAIL.n69 3.49141
R352 VTAIL.n45 VTAIL.n43 3.11257
R353 VTAIL.n81 VTAIL.n45 3.11257
R354 VTAIL.n85 VTAIL.n83 3.11257
R355 VTAIL.n121 VTAIL.n85 3.11257
R356 VTAIL.n41 VTAIL.n39 3.11257
R357 VTAIL.n39 VTAIL.n37 3.11257
R358 VTAIL.n159 VTAIL.n157 3.11257
R359 VTAIL.n142 VTAIL.n128 2.71565
R360 VTAIL.n22 VTAIL.n8 2.71565
R361 VTAIL.n106 VTAIL.n92 2.71565
R362 VTAIL.n66 VTAIL.n52 2.71565
R363 VTAIL VTAIL.n1 2.39274
R364 VTAIL.n83 VTAIL.n81 2.02636
R365 VTAIL.n37 VTAIL.n1 2.02636
R366 VTAIL.n141 VTAIL.n130 1.93989
R367 VTAIL.n21 VTAIL.n10 1.93989
R368 VTAIL.n105 VTAIL.n94 1.93989
R369 VTAIL.n65 VTAIL.n54 1.93989
R370 VTAIL.n138 VTAIL.n137 1.16414
R371 VTAIL.n18 VTAIL.n17 1.16414
R372 VTAIL.n102 VTAIL.n101 1.16414
R373 VTAIL.n62 VTAIL.n61 1.16414
R374 VTAIL VTAIL.n159 0.720328
R375 VTAIL.n134 VTAIL.n132 0.388379
R376 VTAIL.n14 VTAIL.n12 0.388379
R377 VTAIL.n98 VTAIL.n96 0.388379
R378 VTAIL.n58 VTAIL.n56 0.388379
R379 VTAIL.n139 VTAIL.n131 0.155672
R380 VTAIL.n140 VTAIL.n139 0.155672
R381 VTAIL.n140 VTAIL.n127 0.155672
R382 VTAIL.n147 VTAIL.n127 0.155672
R383 VTAIL.n148 VTAIL.n147 0.155672
R384 VTAIL.n148 VTAIL.n123 0.155672
R385 VTAIL.n155 VTAIL.n123 0.155672
R386 VTAIL.n19 VTAIL.n11 0.155672
R387 VTAIL.n20 VTAIL.n19 0.155672
R388 VTAIL.n20 VTAIL.n7 0.155672
R389 VTAIL.n27 VTAIL.n7 0.155672
R390 VTAIL.n28 VTAIL.n27 0.155672
R391 VTAIL.n28 VTAIL.n3 0.155672
R392 VTAIL.n35 VTAIL.n3 0.155672
R393 VTAIL.n119 VTAIL.n87 0.155672
R394 VTAIL.n112 VTAIL.n87 0.155672
R395 VTAIL.n112 VTAIL.n111 0.155672
R396 VTAIL.n111 VTAIL.n91 0.155672
R397 VTAIL.n104 VTAIL.n91 0.155672
R398 VTAIL.n104 VTAIL.n103 0.155672
R399 VTAIL.n103 VTAIL.n95 0.155672
R400 VTAIL.n79 VTAIL.n47 0.155672
R401 VTAIL.n72 VTAIL.n47 0.155672
R402 VTAIL.n72 VTAIL.n71 0.155672
R403 VTAIL.n71 VTAIL.n51 0.155672
R404 VTAIL.n64 VTAIL.n51 0.155672
R405 VTAIL.n64 VTAIL.n63 0.155672
R406 VTAIL.n63 VTAIL.n55 0.155672
R407 VDD2.n69 VDD2.n39 756.745
R408 VDD2.n30 VDD2.n0 756.745
R409 VDD2.n70 VDD2.n69 585
R410 VDD2.n68 VDD2.n67 585
R411 VDD2.n43 VDD2.n42 585
R412 VDD2.n62 VDD2.n61 585
R413 VDD2.n60 VDD2.n59 585
R414 VDD2.n47 VDD2.n46 585
R415 VDD2.n54 VDD2.n53 585
R416 VDD2.n52 VDD2.n51 585
R417 VDD2.n13 VDD2.n12 585
R418 VDD2.n15 VDD2.n14 585
R419 VDD2.n8 VDD2.n7 585
R420 VDD2.n21 VDD2.n20 585
R421 VDD2.n23 VDD2.n22 585
R422 VDD2.n4 VDD2.n3 585
R423 VDD2.n29 VDD2.n28 585
R424 VDD2.n31 VDD2.n30 585
R425 VDD2.n50 VDD2.t5 327.514
R426 VDD2.n11 VDD2.t1 327.514
R427 VDD2.n69 VDD2.n68 171.744
R428 VDD2.n68 VDD2.n42 171.744
R429 VDD2.n61 VDD2.n42 171.744
R430 VDD2.n61 VDD2.n60 171.744
R431 VDD2.n60 VDD2.n46 171.744
R432 VDD2.n53 VDD2.n46 171.744
R433 VDD2.n53 VDD2.n52 171.744
R434 VDD2.n14 VDD2.n13 171.744
R435 VDD2.n14 VDD2.n7 171.744
R436 VDD2.n21 VDD2.n7 171.744
R437 VDD2.n22 VDD2.n21 171.744
R438 VDD2.n22 VDD2.n3 171.744
R439 VDD2.n29 VDD2.n3 171.744
R440 VDD2.n30 VDD2.n29 171.744
R441 VDD2.n38 VDD2.n37 88.7381
R442 VDD2 VDD2.n77 88.7353
R443 VDD2.n76 VDD2.n75 86.4596
R444 VDD2.n36 VDD2.n35 86.4594
R445 VDD2.n52 VDD2.t5 85.8723
R446 VDD2.n13 VDD2.t1 85.8723
R447 VDD2.n36 VDD2.n34 50.0368
R448 VDD2.n74 VDD2.n73 46.9247
R449 VDD2.n74 VDD2.n38 44.2045
R450 VDD2.n12 VDD2.n11 16.3884
R451 VDD2.n51 VDD2.n50 16.3884
R452 VDD2.n54 VDD2.n49 12.8005
R453 VDD2.n15 VDD2.n10 12.8005
R454 VDD2.n55 VDD2.n47 12.0247
R455 VDD2.n16 VDD2.n8 12.0247
R456 VDD2.n59 VDD2.n58 11.249
R457 VDD2.n20 VDD2.n19 11.249
R458 VDD2.n62 VDD2.n45 10.4732
R459 VDD2.n23 VDD2.n6 10.4732
R460 VDD2.n63 VDD2.n43 9.69747
R461 VDD2.n24 VDD2.n4 9.69747
R462 VDD2.n73 VDD2.n72 9.45567
R463 VDD2.n34 VDD2.n33 9.45567
R464 VDD2.n72 VDD2.n71 9.3005
R465 VDD2.n41 VDD2.n40 9.3005
R466 VDD2.n66 VDD2.n65 9.3005
R467 VDD2.n64 VDD2.n63 9.3005
R468 VDD2.n45 VDD2.n44 9.3005
R469 VDD2.n58 VDD2.n57 9.3005
R470 VDD2.n56 VDD2.n55 9.3005
R471 VDD2.n49 VDD2.n48 9.3005
R472 VDD2.n2 VDD2.n1 9.3005
R473 VDD2.n27 VDD2.n26 9.3005
R474 VDD2.n25 VDD2.n24 9.3005
R475 VDD2.n6 VDD2.n5 9.3005
R476 VDD2.n19 VDD2.n18 9.3005
R477 VDD2.n17 VDD2.n16 9.3005
R478 VDD2.n10 VDD2.n9 9.3005
R479 VDD2.n33 VDD2.n32 9.3005
R480 VDD2.n67 VDD2.n66 8.92171
R481 VDD2.n28 VDD2.n27 8.92171
R482 VDD2.n70 VDD2.n41 8.14595
R483 VDD2.n31 VDD2.n2 8.14595
R484 VDD2.n71 VDD2.n39 7.3702
R485 VDD2.n32 VDD2.n0 7.3702
R486 VDD2.n73 VDD2.n39 6.59444
R487 VDD2.n34 VDD2.n0 6.59444
R488 VDD2.n71 VDD2.n70 5.81868
R489 VDD2.n32 VDD2.n31 5.81868
R490 VDD2.n67 VDD2.n41 5.04292
R491 VDD2.n28 VDD2.n2 5.04292
R492 VDD2.n77 VDD2.t6 4.91062
R493 VDD2.n77 VDD2.t3 4.91062
R494 VDD2.n75 VDD2.t0 4.91062
R495 VDD2.n75 VDD2.t9 4.91062
R496 VDD2.n37 VDD2.t4 4.91062
R497 VDD2.n37 VDD2.t2 4.91062
R498 VDD2.n35 VDD2.t7 4.91062
R499 VDD2.n35 VDD2.t8 4.91062
R500 VDD2.n66 VDD2.n43 4.26717
R501 VDD2.n27 VDD2.n4 4.26717
R502 VDD2.n50 VDD2.n48 3.71088
R503 VDD2.n11 VDD2.n9 3.71088
R504 VDD2.n63 VDD2.n62 3.49141
R505 VDD2.n24 VDD2.n23 3.49141
R506 VDD2.n76 VDD2.n74 3.11257
R507 VDD2.n59 VDD2.n45 2.71565
R508 VDD2.n20 VDD2.n6 2.71565
R509 VDD2.n58 VDD2.n47 1.93989
R510 VDD2.n19 VDD2.n8 1.93989
R511 VDD2.n55 VDD2.n54 1.16414
R512 VDD2.n16 VDD2.n15 1.16414
R513 VDD2 VDD2.n76 0.836707
R514 VDD2.n38 VDD2.n36 0.723171
R515 VDD2.n51 VDD2.n49 0.388379
R516 VDD2.n12 VDD2.n10 0.388379
R517 VDD2.n72 VDD2.n40 0.155672
R518 VDD2.n65 VDD2.n40 0.155672
R519 VDD2.n65 VDD2.n64 0.155672
R520 VDD2.n64 VDD2.n44 0.155672
R521 VDD2.n57 VDD2.n44 0.155672
R522 VDD2.n57 VDD2.n56 0.155672
R523 VDD2.n56 VDD2.n48 0.155672
R524 VDD2.n17 VDD2.n9 0.155672
R525 VDD2.n18 VDD2.n17 0.155672
R526 VDD2.n18 VDD2.n5 0.155672
R527 VDD2.n25 VDD2.n5 0.155672
R528 VDD2.n26 VDD2.n25 0.155672
R529 VDD2.n26 VDD2.n1 0.155672
R530 VDD2.n33 VDD2.n1 0.155672
R531 VP.n32 VP.n31 161.3
R532 VP.n33 VP.n28 161.3
R533 VP.n35 VP.n34 161.3
R534 VP.n36 VP.n27 161.3
R535 VP.n38 VP.n37 161.3
R536 VP.n39 VP.n26 161.3
R537 VP.n41 VP.n40 161.3
R538 VP.n42 VP.n25 161.3
R539 VP.n44 VP.n43 161.3
R540 VP.n45 VP.n24 161.3
R541 VP.n47 VP.n46 161.3
R542 VP.n48 VP.n23 161.3
R543 VP.n50 VP.n49 161.3
R544 VP.n51 VP.n22 161.3
R545 VP.n53 VP.n52 161.3
R546 VP.n55 VP.n54 161.3
R547 VP.n56 VP.n20 161.3
R548 VP.n58 VP.n57 161.3
R549 VP.n59 VP.n19 161.3
R550 VP.n61 VP.n60 161.3
R551 VP.n62 VP.n18 161.3
R552 VP.n64 VP.n63 161.3
R553 VP.n111 VP.n110 161.3
R554 VP.n109 VP.n1 161.3
R555 VP.n108 VP.n107 161.3
R556 VP.n106 VP.n2 161.3
R557 VP.n105 VP.n104 161.3
R558 VP.n103 VP.n3 161.3
R559 VP.n102 VP.n101 161.3
R560 VP.n100 VP.n99 161.3
R561 VP.n98 VP.n5 161.3
R562 VP.n97 VP.n96 161.3
R563 VP.n95 VP.n6 161.3
R564 VP.n94 VP.n93 161.3
R565 VP.n92 VP.n7 161.3
R566 VP.n91 VP.n90 161.3
R567 VP.n89 VP.n8 161.3
R568 VP.n88 VP.n87 161.3
R569 VP.n86 VP.n9 161.3
R570 VP.n85 VP.n84 161.3
R571 VP.n83 VP.n10 161.3
R572 VP.n82 VP.n81 161.3
R573 VP.n80 VP.n11 161.3
R574 VP.n79 VP.n78 161.3
R575 VP.n77 VP.n76 161.3
R576 VP.n75 VP.n13 161.3
R577 VP.n74 VP.n73 161.3
R578 VP.n72 VP.n14 161.3
R579 VP.n71 VP.n70 161.3
R580 VP.n69 VP.n15 161.3
R581 VP.n68 VP.n67 161.3
R582 VP.n30 VP.t3 81.0194
R583 VP.n66 VP.n16 79.4252
R584 VP.n112 VP.n0 79.4252
R585 VP.n65 VP.n17 79.4252
R586 VP.n30 VP.n29 69.3368
R587 VP.n85 VP.n10 56.5617
R588 VP.n93 VP.n6 56.5617
R589 VP.n46 VP.n23 56.5617
R590 VP.n38 VP.n27 56.5617
R591 VP.n66 VP.n65 52.7836
R592 VP.n74 VP.n14 48.8116
R593 VP.n104 VP.n2 48.8116
R594 VP.n57 VP.n19 48.8116
R595 VP.n8 VP.t1 48.6414
R596 VP.n16 VP.t5 48.6414
R597 VP.n12 VP.t7 48.6414
R598 VP.n4 VP.t0 48.6414
R599 VP.n0 VP.t8 48.6414
R600 VP.n25 VP.t6 48.6414
R601 VP.n17 VP.t9 48.6414
R602 VP.n21 VP.t4 48.6414
R603 VP.n29 VP.t2 48.6414
R604 VP.n70 VP.n14 32.3425
R605 VP.n108 VP.n2 32.3425
R606 VP.n61 VP.n19 32.3425
R607 VP.n69 VP.n68 24.5923
R608 VP.n70 VP.n69 24.5923
R609 VP.n75 VP.n74 24.5923
R610 VP.n76 VP.n75 24.5923
R611 VP.n80 VP.n79 24.5923
R612 VP.n81 VP.n80 24.5923
R613 VP.n81 VP.n10 24.5923
R614 VP.n86 VP.n85 24.5923
R615 VP.n87 VP.n86 24.5923
R616 VP.n87 VP.n8 24.5923
R617 VP.n91 VP.n8 24.5923
R618 VP.n92 VP.n91 24.5923
R619 VP.n93 VP.n92 24.5923
R620 VP.n97 VP.n6 24.5923
R621 VP.n98 VP.n97 24.5923
R622 VP.n99 VP.n98 24.5923
R623 VP.n103 VP.n102 24.5923
R624 VP.n104 VP.n103 24.5923
R625 VP.n109 VP.n108 24.5923
R626 VP.n110 VP.n109 24.5923
R627 VP.n62 VP.n61 24.5923
R628 VP.n63 VP.n62 24.5923
R629 VP.n50 VP.n23 24.5923
R630 VP.n51 VP.n50 24.5923
R631 VP.n52 VP.n51 24.5923
R632 VP.n56 VP.n55 24.5923
R633 VP.n57 VP.n56 24.5923
R634 VP.n39 VP.n38 24.5923
R635 VP.n40 VP.n39 24.5923
R636 VP.n40 VP.n25 24.5923
R637 VP.n44 VP.n25 24.5923
R638 VP.n45 VP.n44 24.5923
R639 VP.n46 VP.n45 24.5923
R640 VP.n33 VP.n32 24.5923
R641 VP.n34 VP.n33 24.5923
R642 VP.n34 VP.n27 24.5923
R643 VP.n76 VP.n12 19.1821
R644 VP.n102 VP.n4 19.1821
R645 VP.n55 VP.n21 19.1821
R646 VP.n68 VP.n16 10.8209
R647 VP.n110 VP.n0 10.8209
R648 VP.n63 VP.n17 10.8209
R649 VP.n79 VP.n12 5.4107
R650 VP.n99 VP.n4 5.4107
R651 VP.n52 VP.n21 5.4107
R652 VP.n32 VP.n29 5.4107
R653 VP.n31 VP.n30 4.34641
R654 VP.n65 VP.n64 0.354861
R655 VP.n67 VP.n66 0.354861
R656 VP.n112 VP.n111 0.354861
R657 VP VP.n112 0.267071
R658 VP.n31 VP.n28 0.189894
R659 VP.n35 VP.n28 0.189894
R660 VP.n36 VP.n35 0.189894
R661 VP.n37 VP.n36 0.189894
R662 VP.n37 VP.n26 0.189894
R663 VP.n41 VP.n26 0.189894
R664 VP.n42 VP.n41 0.189894
R665 VP.n43 VP.n42 0.189894
R666 VP.n43 VP.n24 0.189894
R667 VP.n47 VP.n24 0.189894
R668 VP.n48 VP.n47 0.189894
R669 VP.n49 VP.n48 0.189894
R670 VP.n49 VP.n22 0.189894
R671 VP.n53 VP.n22 0.189894
R672 VP.n54 VP.n53 0.189894
R673 VP.n54 VP.n20 0.189894
R674 VP.n58 VP.n20 0.189894
R675 VP.n59 VP.n58 0.189894
R676 VP.n60 VP.n59 0.189894
R677 VP.n60 VP.n18 0.189894
R678 VP.n64 VP.n18 0.189894
R679 VP.n67 VP.n15 0.189894
R680 VP.n71 VP.n15 0.189894
R681 VP.n72 VP.n71 0.189894
R682 VP.n73 VP.n72 0.189894
R683 VP.n73 VP.n13 0.189894
R684 VP.n77 VP.n13 0.189894
R685 VP.n78 VP.n77 0.189894
R686 VP.n78 VP.n11 0.189894
R687 VP.n82 VP.n11 0.189894
R688 VP.n83 VP.n82 0.189894
R689 VP.n84 VP.n83 0.189894
R690 VP.n84 VP.n9 0.189894
R691 VP.n88 VP.n9 0.189894
R692 VP.n89 VP.n88 0.189894
R693 VP.n90 VP.n89 0.189894
R694 VP.n90 VP.n7 0.189894
R695 VP.n94 VP.n7 0.189894
R696 VP.n95 VP.n94 0.189894
R697 VP.n96 VP.n95 0.189894
R698 VP.n96 VP.n5 0.189894
R699 VP.n100 VP.n5 0.189894
R700 VP.n101 VP.n100 0.189894
R701 VP.n101 VP.n3 0.189894
R702 VP.n105 VP.n3 0.189894
R703 VP.n106 VP.n105 0.189894
R704 VP.n107 VP.n106 0.189894
R705 VP.n107 VP.n1 0.189894
R706 VP.n111 VP.n1 0.189894
R707 VDD1.n30 VDD1.n0 756.745
R708 VDD1.n67 VDD1.n37 756.745
R709 VDD1.n31 VDD1.n30 585
R710 VDD1.n29 VDD1.n28 585
R711 VDD1.n4 VDD1.n3 585
R712 VDD1.n23 VDD1.n22 585
R713 VDD1.n21 VDD1.n20 585
R714 VDD1.n8 VDD1.n7 585
R715 VDD1.n15 VDD1.n14 585
R716 VDD1.n13 VDD1.n12 585
R717 VDD1.n50 VDD1.n49 585
R718 VDD1.n52 VDD1.n51 585
R719 VDD1.n45 VDD1.n44 585
R720 VDD1.n58 VDD1.n57 585
R721 VDD1.n60 VDD1.n59 585
R722 VDD1.n41 VDD1.n40 585
R723 VDD1.n66 VDD1.n65 585
R724 VDD1.n68 VDD1.n67 585
R725 VDD1.n11 VDD1.t6 327.514
R726 VDD1.n48 VDD1.t4 327.514
R727 VDD1.n30 VDD1.n29 171.744
R728 VDD1.n29 VDD1.n3 171.744
R729 VDD1.n22 VDD1.n3 171.744
R730 VDD1.n22 VDD1.n21 171.744
R731 VDD1.n21 VDD1.n7 171.744
R732 VDD1.n14 VDD1.n7 171.744
R733 VDD1.n14 VDD1.n13 171.744
R734 VDD1.n51 VDD1.n50 171.744
R735 VDD1.n51 VDD1.n44 171.744
R736 VDD1.n58 VDD1.n44 171.744
R737 VDD1.n59 VDD1.n58 171.744
R738 VDD1.n59 VDD1.n40 171.744
R739 VDD1.n66 VDD1.n40 171.744
R740 VDD1.n67 VDD1.n66 171.744
R741 VDD1.n75 VDD1.n74 88.7381
R742 VDD1.n36 VDD1.n35 86.4596
R743 VDD1.n77 VDD1.n76 86.4594
R744 VDD1.n73 VDD1.n72 86.4594
R745 VDD1.n13 VDD1.t6 85.8723
R746 VDD1.n50 VDD1.t4 85.8723
R747 VDD1.n36 VDD1.n34 50.0368
R748 VDD1.n73 VDD1.n71 50.0368
R749 VDD1.n77 VDD1.n75 46.3436
R750 VDD1.n49 VDD1.n48 16.3884
R751 VDD1.n12 VDD1.n11 16.3884
R752 VDD1.n15 VDD1.n10 12.8005
R753 VDD1.n52 VDD1.n47 12.8005
R754 VDD1.n16 VDD1.n8 12.0247
R755 VDD1.n53 VDD1.n45 12.0247
R756 VDD1.n20 VDD1.n19 11.249
R757 VDD1.n57 VDD1.n56 11.249
R758 VDD1.n23 VDD1.n6 10.4732
R759 VDD1.n60 VDD1.n43 10.4732
R760 VDD1.n24 VDD1.n4 9.69747
R761 VDD1.n61 VDD1.n41 9.69747
R762 VDD1.n34 VDD1.n33 9.45567
R763 VDD1.n71 VDD1.n70 9.45567
R764 VDD1.n33 VDD1.n32 9.3005
R765 VDD1.n2 VDD1.n1 9.3005
R766 VDD1.n27 VDD1.n26 9.3005
R767 VDD1.n25 VDD1.n24 9.3005
R768 VDD1.n6 VDD1.n5 9.3005
R769 VDD1.n19 VDD1.n18 9.3005
R770 VDD1.n17 VDD1.n16 9.3005
R771 VDD1.n10 VDD1.n9 9.3005
R772 VDD1.n39 VDD1.n38 9.3005
R773 VDD1.n64 VDD1.n63 9.3005
R774 VDD1.n62 VDD1.n61 9.3005
R775 VDD1.n43 VDD1.n42 9.3005
R776 VDD1.n56 VDD1.n55 9.3005
R777 VDD1.n54 VDD1.n53 9.3005
R778 VDD1.n47 VDD1.n46 9.3005
R779 VDD1.n70 VDD1.n69 9.3005
R780 VDD1.n28 VDD1.n27 8.92171
R781 VDD1.n65 VDD1.n64 8.92171
R782 VDD1.n31 VDD1.n2 8.14595
R783 VDD1.n68 VDD1.n39 8.14595
R784 VDD1.n32 VDD1.n0 7.3702
R785 VDD1.n69 VDD1.n37 7.3702
R786 VDD1.n34 VDD1.n0 6.59444
R787 VDD1.n71 VDD1.n37 6.59444
R788 VDD1.n32 VDD1.n31 5.81868
R789 VDD1.n69 VDD1.n68 5.81868
R790 VDD1.n28 VDD1.n2 5.04292
R791 VDD1.n65 VDD1.n39 5.04292
R792 VDD1.n76 VDD1.t5 4.91062
R793 VDD1.n76 VDD1.t0 4.91062
R794 VDD1.n35 VDD1.t7 4.91062
R795 VDD1.n35 VDD1.t3 4.91062
R796 VDD1.n74 VDD1.t9 4.91062
R797 VDD1.n74 VDD1.t1 4.91062
R798 VDD1.n72 VDD1.t2 4.91062
R799 VDD1.n72 VDD1.t8 4.91062
R800 VDD1.n27 VDD1.n4 4.26717
R801 VDD1.n64 VDD1.n41 4.26717
R802 VDD1.n11 VDD1.n9 3.71088
R803 VDD1.n48 VDD1.n46 3.71088
R804 VDD1.n24 VDD1.n23 3.49141
R805 VDD1.n61 VDD1.n60 3.49141
R806 VDD1.n20 VDD1.n6 2.71565
R807 VDD1.n57 VDD1.n43 2.71565
R808 VDD1 VDD1.n77 2.27636
R809 VDD1.n19 VDD1.n8 1.93989
R810 VDD1.n56 VDD1.n45 1.93989
R811 VDD1.n16 VDD1.n15 1.16414
R812 VDD1.n53 VDD1.n52 1.16414
R813 VDD1 VDD1.n36 0.836707
R814 VDD1.n75 VDD1.n73 0.723171
R815 VDD1.n12 VDD1.n10 0.388379
R816 VDD1.n49 VDD1.n47 0.388379
R817 VDD1.n33 VDD1.n1 0.155672
R818 VDD1.n26 VDD1.n1 0.155672
R819 VDD1.n26 VDD1.n25 0.155672
R820 VDD1.n25 VDD1.n5 0.155672
R821 VDD1.n18 VDD1.n5 0.155672
R822 VDD1.n18 VDD1.n17 0.155672
R823 VDD1.n17 VDD1.n9 0.155672
R824 VDD1.n54 VDD1.n46 0.155672
R825 VDD1.n55 VDD1.n54 0.155672
R826 VDD1.n55 VDD1.n42 0.155672
R827 VDD1.n62 VDD1.n42 0.155672
R828 VDD1.n63 VDD1.n62 0.155672
R829 VDD1.n63 VDD1.n38 0.155672
R830 VDD1.n70 VDD1.n38 0.155672
R831 B.n633 B.n72 585
R832 B.n635 B.n634 585
R833 B.n636 B.n71 585
R834 B.n638 B.n637 585
R835 B.n639 B.n70 585
R836 B.n641 B.n640 585
R837 B.n642 B.n69 585
R838 B.n644 B.n643 585
R839 B.n645 B.n68 585
R840 B.n647 B.n646 585
R841 B.n648 B.n67 585
R842 B.n650 B.n649 585
R843 B.n651 B.n66 585
R844 B.n653 B.n652 585
R845 B.n654 B.n65 585
R846 B.n656 B.n655 585
R847 B.n657 B.n64 585
R848 B.n659 B.n658 585
R849 B.n660 B.n63 585
R850 B.n662 B.n661 585
R851 B.n663 B.n62 585
R852 B.n665 B.n664 585
R853 B.n666 B.n61 585
R854 B.n668 B.n667 585
R855 B.n669 B.n60 585
R856 B.n671 B.n670 585
R857 B.n673 B.n57 585
R858 B.n675 B.n674 585
R859 B.n676 B.n56 585
R860 B.n678 B.n677 585
R861 B.n679 B.n55 585
R862 B.n681 B.n680 585
R863 B.n682 B.n54 585
R864 B.n684 B.n683 585
R865 B.n685 B.n51 585
R866 B.n688 B.n687 585
R867 B.n689 B.n50 585
R868 B.n691 B.n690 585
R869 B.n692 B.n49 585
R870 B.n694 B.n693 585
R871 B.n695 B.n48 585
R872 B.n697 B.n696 585
R873 B.n698 B.n47 585
R874 B.n700 B.n699 585
R875 B.n701 B.n46 585
R876 B.n703 B.n702 585
R877 B.n704 B.n45 585
R878 B.n706 B.n705 585
R879 B.n707 B.n44 585
R880 B.n709 B.n708 585
R881 B.n710 B.n43 585
R882 B.n712 B.n711 585
R883 B.n713 B.n42 585
R884 B.n715 B.n714 585
R885 B.n716 B.n41 585
R886 B.n718 B.n717 585
R887 B.n719 B.n40 585
R888 B.n721 B.n720 585
R889 B.n722 B.n39 585
R890 B.n724 B.n723 585
R891 B.n725 B.n38 585
R892 B.n632 B.n631 585
R893 B.n630 B.n73 585
R894 B.n629 B.n628 585
R895 B.n627 B.n74 585
R896 B.n626 B.n625 585
R897 B.n624 B.n75 585
R898 B.n623 B.n622 585
R899 B.n621 B.n76 585
R900 B.n620 B.n619 585
R901 B.n618 B.n77 585
R902 B.n617 B.n616 585
R903 B.n615 B.n78 585
R904 B.n614 B.n613 585
R905 B.n612 B.n79 585
R906 B.n611 B.n610 585
R907 B.n609 B.n80 585
R908 B.n608 B.n607 585
R909 B.n606 B.n81 585
R910 B.n605 B.n604 585
R911 B.n603 B.n82 585
R912 B.n602 B.n601 585
R913 B.n600 B.n83 585
R914 B.n599 B.n598 585
R915 B.n597 B.n84 585
R916 B.n596 B.n595 585
R917 B.n594 B.n85 585
R918 B.n593 B.n592 585
R919 B.n591 B.n86 585
R920 B.n590 B.n589 585
R921 B.n588 B.n87 585
R922 B.n587 B.n586 585
R923 B.n585 B.n88 585
R924 B.n584 B.n583 585
R925 B.n582 B.n89 585
R926 B.n581 B.n580 585
R927 B.n579 B.n90 585
R928 B.n578 B.n577 585
R929 B.n576 B.n91 585
R930 B.n575 B.n574 585
R931 B.n573 B.n92 585
R932 B.n572 B.n571 585
R933 B.n570 B.n93 585
R934 B.n569 B.n568 585
R935 B.n567 B.n94 585
R936 B.n566 B.n565 585
R937 B.n564 B.n95 585
R938 B.n563 B.n562 585
R939 B.n561 B.n96 585
R940 B.n560 B.n559 585
R941 B.n558 B.n97 585
R942 B.n557 B.n556 585
R943 B.n555 B.n98 585
R944 B.n554 B.n553 585
R945 B.n552 B.n99 585
R946 B.n551 B.n550 585
R947 B.n549 B.n100 585
R948 B.n548 B.n547 585
R949 B.n546 B.n101 585
R950 B.n545 B.n544 585
R951 B.n543 B.n102 585
R952 B.n542 B.n541 585
R953 B.n540 B.n103 585
R954 B.n539 B.n538 585
R955 B.n537 B.n104 585
R956 B.n536 B.n535 585
R957 B.n534 B.n105 585
R958 B.n533 B.n532 585
R959 B.n531 B.n106 585
R960 B.n530 B.n529 585
R961 B.n528 B.n107 585
R962 B.n527 B.n526 585
R963 B.n525 B.n108 585
R964 B.n524 B.n523 585
R965 B.n522 B.n109 585
R966 B.n521 B.n520 585
R967 B.n519 B.n110 585
R968 B.n518 B.n517 585
R969 B.n516 B.n111 585
R970 B.n515 B.n514 585
R971 B.n513 B.n112 585
R972 B.n512 B.n511 585
R973 B.n510 B.n113 585
R974 B.n509 B.n508 585
R975 B.n507 B.n114 585
R976 B.n506 B.n505 585
R977 B.n504 B.n115 585
R978 B.n503 B.n502 585
R979 B.n501 B.n116 585
R980 B.n500 B.n499 585
R981 B.n498 B.n117 585
R982 B.n497 B.n496 585
R983 B.n495 B.n118 585
R984 B.n494 B.n493 585
R985 B.n492 B.n119 585
R986 B.n491 B.n490 585
R987 B.n489 B.n120 585
R988 B.n488 B.n487 585
R989 B.n486 B.n121 585
R990 B.n485 B.n484 585
R991 B.n483 B.n122 585
R992 B.n482 B.n481 585
R993 B.n480 B.n123 585
R994 B.n479 B.n478 585
R995 B.n477 B.n124 585
R996 B.n476 B.n475 585
R997 B.n474 B.n125 585
R998 B.n473 B.n472 585
R999 B.n471 B.n126 585
R1000 B.n470 B.n469 585
R1001 B.n468 B.n127 585
R1002 B.n467 B.n466 585
R1003 B.n465 B.n128 585
R1004 B.n464 B.n463 585
R1005 B.n462 B.n129 585
R1006 B.n461 B.n460 585
R1007 B.n459 B.n130 585
R1008 B.n458 B.n457 585
R1009 B.n456 B.n131 585
R1010 B.n455 B.n454 585
R1011 B.n453 B.n132 585
R1012 B.n452 B.n451 585
R1013 B.n450 B.n133 585
R1014 B.n449 B.n448 585
R1015 B.n447 B.n134 585
R1016 B.n446 B.n445 585
R1017 B.n444 B.n135 585
R1018 B.n443 B.n442 585
R1019 B.n441 B.n136 585
R1020 B.n440 B.n439 585
R1021 B.n438 B.n137 585
R1022 B.n437 B.n436 585
R1023 B.n435 B.n138 585
R1024 B.n434 B.n433 585
R1025 B.n432 B.n139 585
R1026 B.n431 B.n430 585
R1027 B.n429 B.n140 585
R1028 B.n428 B.n427 585
R1029 B.n426 B.n141 585
R1030 B.n425 B.n424 585
R1031 B.n423 B.n142 585
R1032 B.n422 B.n421 585
R1033 B.n420 B.n143 585
R1034 B.n419 B.n418 585
R1035 B.n417 B.n144 585
R1036 B.n416 B.n415 585
R1037 B.n323 B.n322 585
R1038 B.n324 B.n179 585
R1039 B.n326 B.n325 585
R1040 B.n327 B.n178 585
R1041 B.n329 B.n328 585
R1042 B.n330 B.n177 585
R1043 B.n332 B.n331 585
R1044 B.n333 B.n176 585
R1045 B.n335 B.n334 585
R1046 B.n336 B.n175 585
R1047 B.n338 B.n337 585
R1048 B.n339 B.n174 585
R1049 B.n341 B.n340 585
R1050 B.n342 B.n173 585
R1051 B.n344 B.n343 585
R1052 B.n345 B.n172 585
R1053 B.n347 B.n346 585
R1054 B.n348 B.n171 585
R1055 B.n350 B.n349 585
R1056 B.n351 B.n170 585
R1057 B.n353 B.n352 585
R1058 B.n354 B.n169 585
R1059 B.n356 B.n355 585
R1060 B.n357 B.n168 585
R1061 B.n359 B.n358 585
R1062 B.n360 B.n165 585
R1063 B.n363 B.n362 585
R1064 B.n364 B.n164 585
R1065 B.n366 B.n365 585
R1066 B.n367 B.n163 585
R1067 B.n369 B.n368 585
R1068 B.n370 B.n162 585
R1069 B.n372 B.n371 585
R1070 B.n373 B.n161 585
R1071 B.n375 B.n374 585
R1072 B.n377 B.n376 585
R1073 B.n378 B.n157 585
R1074 B.n380 B.n379 585
R1075 B.n381 B.n156 585
R1076 B.n383 B.n382 585
R1077 B.n384 B.n155 585
R1078 B.n386 B.n385 585
R1079 B.n387 B.n154 585
R1080 B.n389 B.n388 585
R1081 B.n390 B.n153 585
R1082 B.n392 B.n391 585
R1083 B.n393 B.n152 585
R1084 B.n395 B.n394 585
R1085 B.n396 B.n151 585
R1086 B.n398 B.n397 585
R1087 B.n399 B.n150 585
R1088 B.n401 B.n400 585
R1089 B.n402 B.n149 585
R1090 B.n404 B.n403 585
R1091 B.n405 B.n148 585
R1092 B.n407 B.n406 585
R1093 B.n408 B.n147 585
R1094 B.n410 B.n409 585
R1095 B.n411 B.n146 585
R1096 B.n413 B.n412 585
R1097 B.n414 B.n145 585
R1098 B.n321 B.n180 585
R1099 B.n320 B.n319 585
R1100 B.n318 B.n181 585
R1101 B.n317 B.n316 585
R1102 B.n315 B.n182 585
R1103 B.n314 B.n313 585
R1104 B.n312 B.n183 585
R1105 B.n311 B.n310 585
R1106 B.n309 B.n184 585
R1107 B.n308 B.n307 585
R1108 B.n306 B.n185 585
R1109 B.n305 B.n304 585
R1110 B.n303 B.n186 585
R1111 B.n302 B.n301 585
R1112 B.n300 B.n187 585
R1113 B.n299 B.n298 585
R1114 B.n297 B.n188 585
R1115 B.n296 B.n295 585
R1116 B.n294 B.n189 585
R1117 B.n293 B.n292 585
R1118 B.n291 B.n190 585
R1119 B.n290 B.n289 585
R1120 B.n288 B.n191 585
R1121 B.n287 B.n286 585
R1122 B.n285 B.n192 585
R1123 B.n284 B.n283 585
R1124 B.n282 B.n193 585
R1125 B.n281 B.n280 585
R1126 B.n279 B.n194 585
R1127 B.n278 B.n277 585
R1128 B.n276 B.n195 585
R1129 B.n275 B.n274 585
R1130 B.n273 B.n196 585
R1131 B.n272 B.n271 585
R1132 B.n270 B.n197 585
R1133 B.n269 B.n268 585
R1134 B.n267 B.n198 585
R1135 B.n266 B.n265 585
R1136 B.n264 B.n199 585
R1137 B.n263 B.n262 585
R1138 B.n261 B.n200 585
R1139 B.n260 B.n259 585
R1140 B.n258 B.n201 585
R1141 B.n257 B.n256 585
R1142 B.n255 B.n202 585
R1143 B.n254 B.n253 585
R1144 B.n252 B.n203 585
R1145 B.n251 B.n250 585
R1146 B.n249 B.n204 585
R1147 B.n248 B.n247 585
R1148 B.n246 B.n205 585
R1149 B.n245 B.n244 585
R1150 B.n243 B.n206 585
R1151 B.n242 B.n241 585
R1152 B.n240 B.n207 585
R1153 B.n239 B.n238 585
R1154 B.n237 B.n208 585
R1155 B.n236 B.n235 585
R1156 B.n234 B.n209 585
R1157 B.n233 B.n232 585
R1158 B.n231 B.n210 585
R1159 B.n230 B.n229 585
R1160 B.n228 B.n211 585
R1161 B.n227 B.n226 585
R1162 B.n225 B.n212 585
R1163 B.n224 B.n223 585
R1164 B.n222 B.n213 585
R1165 B.n221 B.n220 585
R1166 B.n219 B.n214 585
R1167 B.n218 B.n217 585
R1168 B.n216 B.n215 585
R1169 B.n2 B.n0 585
R1170 B.n833 B.n1 585
R1171 B.n832 B.n831 585
R1172 B.n830 B.n3 585
R1173 B.n829 B.n828 585
R1174 B.n827 B.n4 585
R1175 B.n826 B.n825 585
R1176 B.n824 B.n5 585
R1177 B.n823 B.n822 585
R1178 B.n821 B.n6 585
R1179 B.n820 B.n819 585
R1180 B.n818 B.n7 585
R1181 B.n817 B.n816 585
R1182 B.n815 B.n8 585
R1183 B.n814 B.n813 585
R1184 B.n812 B.n9 585
R1185 B.n811 B.n810 585
R1186 B.n809 B.n10 585
R1187 B.n808 B.n807 585
R1188 B.n806 B.n11 585
R1189 B.n805 B.n804 585
R1190 B.n803 B.n12 585
R1191 B.n802 B.n801 585
R1192 B.n800 B.n13 585
R1193 B.n799 B.n798 585
R1194 B.n797 B.n14 585
R1195 B.n796 B.n795 585
R1196 B.n794 B.n15 585
R1197 B.n793 B.n792 585
R1198 B.n791 B.n16 585
R1199 B.n790 B.n789 585
R1200 B.n788 B.n17 585
R1201 B.n787 B.n786 585
R1202 B.n785 B.n18 585
R1203 B.n784 B.n783 585
R1204 B.n782 B.n19 585
R1205 B.n781 B.n780 585
R1206 B.n779 B.n20 585
R1207 B.n778 B.n777 585
R1208 B.n776 B.n21 585
R1209 B.n775 B.n774 585
R1210 B.n773 B.n22 585
R1211 B.n772 B.n771 585
R1212 B.n770 B.n23 585
R1213 B.n769 B.n768 585
R1214 B.n767 B.n24 585
R1215 B.n766 B.n765 585
R1216 B.n764 B.n25 585
R1217 B.n763 B.n762 585
R1218 B.n761 B.n26 585
R1219 B.n760 B.n759 585
R1220 B.n758 B.n27 585
R1221 B.n757 B.n756 585
R1222 B.n755 B.n28 585
R1223 B.n754 B.n753 585
R1224 B.n752 B.n29 585
R1225 B.n751 B.n750 585
R1226 B.n749 B.n30 585
R1227 B.n748 B.n747 585
R1228 B.n746 B.n31 585
R1229 B.n745 B.n744 585
R1230 B.n743 B.n32 585
R1231 B.n742 B.n741 585
R1232 B.n740 B.n33 585
R1233 B.n739 B.n738 585
R1234 B.n737 B.n34 585
R1235 B.n736 B.n735 585
R1236 B.n734 B.n35 585
R1237 B.n733 B.n732 585
R1238 B.n731 B.n36 585
R1239 B.n730 B.n729 585
R1240 B.n728 B.n37 585
R1241 B.n727 B.n726 585
R1242 B.n835 B.n834 585
R1243 B.n322 B.n321 482.89
R1244 B.n726 B.n725 482.89
R1245 B.n416 B.n145 482.89
R1246 B.n633 B.n632 482.89
R1247 B.n158 B.t5 349.036
R1248 B.n58 B.t1 349.036
R1249 B.n166 B.t8 349.034
R1250 B.n52 B.t10 349.034
R1251 B.n159 B.t4 279.022
R1252 B.n59 B.t2 279.022
R1253 B.n167 B.t7 279.022
R1254 B.n53 B.t11 279.022
R1255 B.n158 B.t3 257.526
R1256 B.n166 B.t6 257.526
R1257 B.n52 B.t9 257.526
R1258 B.n58 B.t0 257.526
R1259 B.n321 B.n320 163.367
R1260 B.n320 B.n181 163.367
R1261 B.n316 B.n181 163.367
R1262 B.n316 B.n315 163.367
R1263 B.n315 B.n314 163.367
R1264 B.n314 B.n183 163.367
R1265 B.n310 B.n183 163.367
R1266 B.n310 B.n309 163.367
R1267 B.n309 B.n308 163.367
R1268 B.n308 B.n185 163.367
R1269 B.n304 B.n185 163.367
R1270 B.n304 B.n303 163.367
R1271 B.n303 B.n302 163.367
R1272 B.n302 B.n187 163.367
R1273 B.n298 B.n187 163.367
R1274 B.n298 B.n297 163.367
R1275 B.n297 B.n296 163.367
R1276 B.n296 B.n189 163.367
R1277 B.n292 B.n189 163.367
R1278 B.n292 B.n291 163.367
R1279 B.n291 B.n290 163.367
R1280 B.n290 B.n191 163.367
R1281 B.n286 B.n191 163.367
R1282 B.n286 B.n285 163.367
R1283 B.n285 B.n284 163.367
R1284 B.n284 B.n193 163.367
R1285 B.n280 B.n193 163.367
R1286 B.n280 B.n279 163.367
R1287 B.n279 B.n278 163.367
R1288 B.n278 B.n195 163.367
R1289 B.n274 B.n195 163.367
R1290 B.n274 B.n273 163.367
R1291 B.n273 B.n272 163.367
R1292 B.n272 B.n197 163.367
R1293 B.n268 B.n197 163.367
R1294 B.n268 B.n267 163.367
R1295 B.n267 B.n266 163.367
R1296 B.n266 B.n199 163.367
R1297 B.n262 B.n199 163.367
R1298 B.n262 B.n261 163.367
R1299 B.n261 B.n260 163.367
R1300 B.n260 B.n201 163.367
R1301 B.n256 B.n201 163.367
R1302 B.n256 B.n255 163.367
R1303 B.n255 B.n254 163.367
R1304 B.n254 B.n203 163.367
R1305 B.n250 B.n203 163.367
R1306 B.n250 B.n249 163.367
R1307 B.n249 B.n248 163.367
R1308 B.n248 B.n205 163.367
R1309 B.n244 B.n205 163.367
R1310 B.n244 B.n243 163.367
R1311 B.n243 B.n242 163.367
R1312 B.n242 B.n207 163.367
R1313 B.n238 B.n207 163.367
R1314 B.n238 B.n237 163.367
R1315 B.n237 B.n236 163.367
R1316 B.n236 B.n209 163.367
R1317 B.n232 B.n209 163.367
R1318 B.n232 B.n231 163.367
R1319 B.n231 B.n230 163.367
R1320 B.n230 B.n211 163.367
R1321 B.n226 B.n211 163.367
R1322 B.n226 B.n225 163.367
R1323 B.n225 B.n224 163.367
R1324 B.n224 B.n213 163.367
R1325 B.n220 B.n213 163.367
R1326 B.n220 B.n219 163.367
R1327 B.n219 B.n218 163.367
R1328 B.n218 B.n215 163.367
R1329 B.n215 B.n2 163.367
R1330 B.n834 B.n2 163.367
R1331 B.n834 B.n833 163.367
R1332 B.n833 B.n832 163.367
R1333 B.n832 B.n3 163.367
R1334 B.n828 B.n3 163.367
R1335 B.n828 B.n827 163.367
R1336 B.n827 B.n826 163.367
R1337 B.n826 B.n5 163.367
R1338 B.n822 B.n5 163.367
R1339 B.n822 B.n821 163.367
R1340 B.n821 B.n820 163.367
R1341 B.n820 B.n7 163.367
R1342 B.n816 B.n7 163.367
R1343 B.n816 B.n815 163.367
R1344 B.n815 B.n814 163.367
R1345 B.n814 B.n9 163.367
R1346 B.n810 B.n9 163.367
R1347 B.n810 B.n809 163.367
R1348 B.n809 B.n808 163.367
R1349 B.n808 B.n11 163.367
R1350 B.n804 B.n11 163.367
R1351 B.n804 B.n803 163.367
R1352 B.n803 B.n802 163.367
R1353 B.n802 B.n13 163.367
R1354 B.n798 B.n13 163.367
R1355 B.n798 B.n797 163.367
R1356 B.n797 B.n796 163.367
R1357 B.n796 B.n15 163.367
R1358 B.n792 B.n15 163.367
R1359 B.n792 B.n791 163.367
R1360 B.n791 B.n790 163.367
R1361 B.n790 B.n17 163.367
R1362 B.n786 B.n17 163.367
R1363 B.n786 B.n785 163.367
R1364 B.n785 B.n784 163.367
R1365 B.n784 B.n19 163.367
R1366 B.n780 B.n19 163.367
R1367 B.n780 B.n779 163.367
R1368 B.n779 B.n778 163.367
R1369 B.n778 B.n21 163.367
R1370 B.n774 B.n21 163.367
R1371 B.n774 B.n773 163.367
R1372 B.n773 B.n772 163.367
R1373 B.n772 B.n23 163.367
R1374 B.n768 B.n23 163.367
R1375 B.n768 B.n767 163.367
R1376 B.n767 B.n766 163.367
R1377 B.n766 B.n25 163.367
R1378 B.n762 B.n25 163.367
R1379 B.n762 B.n761 163.367
R1380 B.n761 B.n760 163.367
R1381 B.n760 B.n27 163.367
R1382 B.n756 B.n27 163.367
R1383 B.n756 B.n755 163.367
R1384 B.n755 B.n754 163.367
R1385 B.n754 B.n29 163.367
R1386 B.n750 B.n29 163.367
R1387 B.n750 B.n749 163.367
R1388 B.n749 B.n748 163.367
R1389 B.n748 B.n31 163.367
R1390 B.n744 B.n31 163.367
R1391 B.n744 B.n743 163.367
R1392 B.n743 B.n742 163.367
R1393 B.n742 B.n33 163.367
R1394 B.n738 B.n33 163.367
R1395 B.n738 B.n737 163.367
R1396 B.n737 B.n736 163.367
R1397 B.n736 B.n35 163.367
R1398 B.n732 B.n35 163.367
R1399 B.n732 B.n731 163.367
R1400 B.n731 B.n730 163.367
R1401 B.n730 B.n37 163.367
R1402 B.n726 B.n37 163.367
R1403 B.n322 B.n179 163.367
R1404 B.n326 B.n179 163.367
R1405 B.n327 B.n326 163.367
R1406 B.n328 B.n327 163.367
R1407 B.n328 B.n177 163.367
R1408 B.n332 B.n177 163.367
R1409 B.n333 B.n332 163.367
R1410 B.n334 B.n333 163.367
R1411 B.n334 B.n175 163.367
R1412 B.n338 B.n175 163.367
R1413 B.n339 B.n338 163.367
R1414 B.n340 B.n339 163.367
R1415 B.n340 B.n173 163.367
R1416 B.n344 B.n173 163.367
R1417 B.n345 B.n344 163.367
R1418 B.n346 B.n345 163.367
R1419 B.n346 B.n171 163.367
R1420 B.n350 B.n171 163.367
R1421 B.n351 B.n350 163.367
R1422 B.n352 B.n351 163.367
R1423 B.n352 B.n169 163.367
R1424 B.n356 B.n169 163.367
R1425 B.n357 B.n356 163.367
R1426 B.n358 B.n357 163.367
R1427 B.n358 B.n165 163.367
R1428 B.n363 B.n165 163.367
R1429 B.n364 B.n363 163.367
R1430 B.n365 B.n364 163.367
R1431 B.n365 B.n163 163.367
R1432 B.n369 B.n163 163.367
R1433 B.n370 B.n369 163.367
R1434 B.n371 B.n370 163.367
R1435 B.n371 B.n161 163.367
R1436 B.n375 B.n161 163.367
R1437 B.n376 B.n375 163.367
R1438 B.n376 B.n157 163.367
R1439 B.n380 B.n157 163.367
R1440 B.n381 B.n380 163.367
R1441 B.n382 B.n381 163.367
R1442 B.n382 B.n155 163.367
R1443 B.n386 B.n155 163.367
R1444 B.n387 B.n386 163.367
R1445 B.n388 B.n387 163.367
R1446 B.n388 B.n153 163.367
R1447 B.n392 B.n153 163.367
R1448 B.n393 B.n392 163.367
R1449 B.n394 B.n393 163.367
R1450 B.n394 B.n151 163.367
R1451 B.n398 B.n151 163.367
R1452 B.n399 B.n398 163.367
R1453 B.n400 B.n399 163.367
R1454 B.n400 B.n149 163.367
R1455 B.n404 B.n149 163.367
R1456 B.n405 B.n404 163.367
R1457 B.n406 B.n405 163.367
R1458 B.n406 B.n147 163.367
R1459 B.n410 B.n147 163.367
R1460 B.n411 B.n410 163.367
R1461 B.n412 B.n411 163.367
R1462 B.n412 B.n145 163.367
R1463 B.n417 B.n416 163.367
R1464 B.n418 B.n417 163.367
R1465 B.n418 B.n143 163.367
R1466 B.n422 B.n143 163.367
R1467 B.n423 B.n422 163.367
R1468 B.n424 B.n423 163.367
R1469 B.n424 B.n141 163.367
R1470 B.n428 B.n141 163.367
R1471 B.n429 B.n428 163.367
R1472 B.n430 B.n429 163.367
R1473 B.n430 B.n139 163.367
R1474 B.n434 B.n139 163.367
R1475 B.n435 B.n434 163.367
R1476 B.n436 B.n435 163.367
R1477 B.n436 B.n137 163.367
R1478 B.n440 B.n137 163.367
R1479 B.n441 B.n440 163.367
R1480 B.n442 B.n441 163.367
R1481 B.n442 B.n135 163.367
R1482 B.n446 B.n135 163.367
R1483 B.n447 B.n446 163.367
R1484 B.n448 B.n447 163.367
R1485 B.n448 B.n133 163.367
R1486 B.n452 B.n133 163.367
R1487 B.n453 B.n452 163.367
R1488 B.n454 B.n453 163.367
R1489 B.n454 B.n131 163.367
R1490 B.n458 B.n131 163.367
R1491 B.n459 B.n458 163.367
R1492 B.n460 B.n459 163.367
R1493 B.n460 B.n129 163.367
R1494 B.n464 B.n129 163.367
R1495 B.n465 B.n464 163.367
R1496 B.n466 B.n465 163.367
R1497 B.n466 B.n127 163.367
R1498 B.n470 B.n127 163.367
R1499 B.n471 B.n470 163.367
R1500 B.n472 B.n471 163.367
R1501 B.n472 B.n125 163.367
R1502 B.n476 B.n125 163.367
R1503 B.n477 B.n476 163.367
R1504 B.n478 B.n477 163.367
R1505 B.n478 B.n123 163.367
R1506 B.n482 B.n123 163.367
R1507 B.n483 B.n482 163.367
R1508 B.n484 B.n483 163.367
R1509 B.n484 B.n121 163.367
R1510 B.n488 B.n121 163.367
R1511 B.n489 B.n488 163.367
R1512 B.n490 B.n489 163.367
R1513 B.n490 B.n119 163.367
R1514 B.n494 B.n119 163.367
R1515 B.n495 B.n494 163.367
R1516 B.n496 B.n495 163.367
R1517 B.n496 B.n117 163.367
R1518 B.n500 B.n117 163.367
R1519 B.n501 B.n500 163.367
R1520 B.n502 B.n501 163.367
R1521 B.n502 B.n115 163.367
R1522 B.n506 B.n115 163.367
R1523 B.n507 B.n506 163.367
R1524 B.n508 B.n507 163.367
R1525 B.n508 B.n113 163.367
R1526 B.n512 B.n113 163.367
R1527 B.n513 B.n512 163.367
R1528 B.n514 B.n513 163.367
R1529 B.n514 B.n111 163.367
R1530 B.n518 B.n111 163.367
R1531 B.n519 B.n518 163.367
R1532 B.n520 B.n519 163.367
R1533 B.n520 B.n109 163.367
R1534 B.n524 B.n109 163.367
R1535 B.n525 B.n524 163.367
R1536 B.n526 B.n525 163.367
R1537 B.n526 B.n107 163.367
R1538 B.n530 B.n107 163.367
R1539 B.n531 B.n530 163.367
R1540 B.n532 B.n531 163.367
R1541 B.n532 B.n105 163.367
R1542 B.n536 B.n105 163.367
R1543 B.n537 B.n536 163.367
R1544 B.n538 B.n537 163.367
R1545 B.n538 B.n103 163.367
R1546 B.n542 B.n103 163.367
R1547 B.n543 B.n542 163.367
R1548 B.n544 B.n543 163.367
R1549 B.n544 B.n101 163.367
R1550 B.n548 B.n101 163.367
R1551 B.n549 B.n548 163.367
R1552 B.n550 B.n549 163.367
R1553 B.n550 B.n99 163.367
R1554 B.n554 B.n99 163.367
R1555 B.n555 B.n554 163.367
R1556 B.n556 B.n555 163.367
R1557 B.n556 B.n97 163.367
R1558 B.n560 B.n97 163.367
R1559 B.n561 B.n560 163.367
R1560 B.n562 B.n561 163.367
R1561 B.n562 B.n95 163.367
R1562 B.n566 B.n95 163.367
R1563 B.n567 B.n566 163.367
R1564 B.n568 B.n567 163.367
R1565 B.n568 B.n93 163.367
R1566 B.n572 B.n93 163.367
R1567 B.n573 B.n572 163.367
R1568 B.n574 B.n573 163.367
R1569 B.n574 B.n91 163.367
R1570 B.n578 B.n91 163.367
R1571 B.n579 B.n578 163.367
R1572 B.n580 B.n579 163.367
R1573 B.n580 B.n89 163.367
R1574 B.n584 B.n89 163.367
R1575 B.n585 B.n584 163.367
R1576 B.n586 B.n585 163.367
R1577 B.n586 B.n87 163.367
R1578 B.n590 B.n87 163.367
R1579 B.n591 B.n590 163.367
R1580 B.n592 B.n591 163.367
R1581 B.n592 B.n85 163.367
R1582 B.n596 B.n85 163.367
R1583 B.n597 B.n596 163.367
R1584 B.n598 B.n597 163.367
R1585 B.n598 B.n83 163.367
R1586 B.n602 B.n83 163.367
R1587 B.n603 B.n602 163.367
R1588 B.n604 B.n603 163.367
R1589 B.n604 B.n81 163.367
R1590 B.n608 B.n81 163.367
R1591 B.n609 B.n608 163.367
R1592 B.n610 B.n609 163.367
R1593 B.n610 B.n79 163.367
R1594 B.n614 B.n79 163.367
R1595 B.n615 B.n614 163.367
R1596 B.n616 B.n615 163.367
R1597 B.n616 B.n77 163.367
R1598 B.n620 B.n77 163.367
R1599 B.n621 B.n620 163.367
R1600 B.n622 B.n621 163.367
R1601 B.n622 B.n75 163.367
R1602 B.n626 B.n75 163.367
R1603 B.n627 B.n626 163.367
R1604 B.n628 B.n627 163.367
R1605 B.n628 B.n73 163.367
R1606 B.n632 B.n73 163.367
R1607 B.n725 B.n724 163.367
R1608 B.n724 B.n39 163.367
R1609 B.n720 B.n39 163.367
R1610 B.n720 B.n719 163.367
R1611 B.n719 B.n718 163.367
R1612 B.n718 B.n41 163.367
R1613 B.n714 B.n41 163.367
R1614 B.n714 B.n713 163.367
R1615 B.n713 B.n712 163.367
R1616 B.n712 B.n43 163.367
R1617 B.n708 B.n43 163.367
R1618 B.n708 B.n707 163.367
R1619 B.n707 B.n706 163.367
R1620 B.n706 B.n45 163.367
R1621 B.n702 B.n45 163.367
R1622 B.n702 B.n701 163.367
R1623 B.n701 B.n700 163.367
R1624 B.n700 B.n47 163.367
R1625 B.n696 B.n47 163.367
R1626 B.n696 B.n695 163.367
R1627 B.n695 B.n694 163.367
R1628 B.n694 B.n49 163.367
R1629 B.n690 B.n49 163.367
R1630 B.n690 B.n689 163.367
R1631 B.n689 B.n688 163.367
R1632 B.n688 B.n51 163.367
R1633 B.n683 B.n51 163.367
R1634 B.n683 B.n682 163.367
R1635 B.n682 B.n681 163.367
R1636 B.n681 B.n55 163.367
R1637 B.n677 B.n55 163.367
R1638 B.n677 B.n676 163.367
R1639 B.n676 B.n675 163.367
R1640 B.n675 B.n57 163.367
R1641 B.n670 B.n57 163.367
R1642 B.n670 B.n669 163.367
R1643 B.n669 B.n668 163.367
R1644 B.n668 B.n61 163.367
R1645 B.n664 B.n61 163.367
R1646 B.n664 B.n663 163.367
R1647 B.n663 B.n662 163.367
R1648 B.n662 B.n63 163.367
R1649 B.n658 B.n63 163.367
R1650 B.n658 B.n657 163.367
R1651 B.n657 B.n656 163.367
R1652 B.n656 B.n65 163.367
R1653 B.n652 B.n65 163.367
R1654 B.n652 B.n651 163.367
R1655 B.n651 B.n650 163.367
R1656 B.n650 B.n67 163.367
R1657 B.n646 B.n67 163.367
R1658 B.n646 B.n645 163.367
R1659 B.n645 B.n644 163.367
R1660 B.n644 B.n69 163.367
R1661 B.n640 B.n69 163.367
R1662 B.n640 B.n639 163.367
R1663 B.n639 B.n638 163.367
R1664 B.n638 B.n71 163.367
R1665 B.n634 B.n71 163.367
R1666 B.n634 B.n633 163.367
R1667 B.n159 B.n158 70.0126
R1668 B.n167 B.n166 70.0126
R1669 B.n53 B.n52 70.0126
R1670 B.n59 B.n58 70.0126
R1671 B.n160 B.n159 59.5399
R1672 B.n361 B.n167 59.5399
R1673 B.n686 B.n53 59.5399
R1674 B.n672 B.n59 59.5399
R1675 B.n727 B.n38 31.3761
R1676 B.n631 B.n72 31.3761
R1677 B.n415 B.n414 31.3761
R1678 B.n323 B.n180 31.3761
R1679 B B.n835 18.0485
R1680 B.n723 B.n38 10.6151
R1681 B.n723 B.n722 10.6151
R1682 B.n722 B.n721 10.6151
R1683 B.n721 B.n40 10.6151
R1684 B.n717 B.n40 10.6151
R1685 B.n717 B.n716 10.6151
R1686 B.n716 B.n715 10.6151
R1687 B.n715 B.n42 10.6151
R1688 B.n711 B.n42 10.6151
R1689 B.n711 B.n710 10.6151
R1690 B.n710 B.n709 10.6151
R1691 B.n709 B.n44 10.6151
R1692 B.n705 B.n44 10.6151
R1693 B.n705 B.n704 10.6151
R1694 B.n704 B.n703 10.6151
R1695 B.n703 B.n46 10.6151
R1696 B.n699 B.n46 10.6151
R1697 B.n699 B.n698 10.6151
R1698 B.n698 B.n697 10.6151
R1699 B.n697 B.n48 10.6151
R1700 B.n693 B.n48 10.6151
R1701 B.n693 B.n692 10.6151
R1702 B.n692 B.n691 10.6151
R1703 B.n691 B.n50 10.6151
R1704 B.n687 B.n50 10.6151
R1705 B.n685 B.n684 10.6151
R1706 B.n684 B.n54 10.6151
R1707 B.n680 B.n54 10.6151
R1708 B.n680 B.n679 10.6151
R1709 B.n679 B.n678 10.6151
R1710 B.n678 B.n56 10.6151
R1711 B.n674 B.n56 10.6151
R1712 B.n674 B.n673 10.6151
R1713 B.n671 B.n60 10.6151
R1714 B.n667 B.n60 10.6151
R1715 B.n667 B.n666 10.6151
R1716 B.n666 B.n665 10.6151
R1717 B.n665 B.n62 10.6151
R1718 B.n661 B.n62 10.6151
R1719 B.n661 B.n660 10.6151
R1720 B.n660 B.n659 10.6151
R1721 B.n659 B.n64 10.6151
R1722 B.n655 B.n64 10.6151
R1723 B.n655 B.n654 10.6151
R1724 B.n654 B.n653 10.6151
R1725 B.n653 B.n66 10.6151
R1726 B.n649 B.n66 10.6151
R1727 B.n649 B.n648 10.6151
R1728 B.n648 B.n647 10.6151
R1729 B.n647 B.n68 10.6151
R1730 B.n643 B.n68 10.6151
R1731 B.n643 B.n642 10.6151
R1732 B.n642 B.n641 10.6151
R1733 B.n641 B.n70 10.6151
R1734 B.n637 B.n70 10.6151
R1735 B.n637 B.n636 10.6151
R1736 B.n636 B.n635 10.6151
R1737 B.n635 B.n72 10.6151
R1738 B.n415 B.n144 10.6151
R1739 B.n419 B.n144 10.6151
R1740 B.n420 B.n419 10.6151
R1741 B.n421 B.n420 10.6151
R1742 B.n421 B.n142 10.6151
R1743 B.n425 B.n142 10.6151
R1744 B.n426 B.n425 10.6151
R1745 B.n427 B.n426 10.6151
R1746 B.n427 B.n140 10.6151
R1747 B.n431 B.n140 10.6151
R1748 B.n432 B.n431 10.6151
R1749 B.n433 B.n432 10.6151
R1750 B.n433 B.n138 10.6151
R1751 B.n437 B.n138 10.6151
R1752 B.n438 B.n437 10.6151
R1753 B.n439 B.n438 10.6151
R1754 B.n439 B.n136 10.6151
R1755 B.n443 B.n136 10.6151
R1756 B.n444 B.n443 10.6151
R1757 B.n445 B.n444 10.6151
R1758 B.n445 B.n134 10.6151
R1759 B.n449 B.n134 10.6151
R1760 B.n450 B.n449 10.6151
R1761 B.n451 B.n450 10.6151
R1762 B.n451 B.n132 10.6151
R1763 B.n455 B.n132 10.6151
R1764 B.n456 B.n455 10.6151
R1765 B.n457 B.n456 10.6151
R1766 B.n457 B.n130 10.6151
R1767 B.n461 B.n130 10.6151
R1768 B.n462 B.n461 10.6151
R1769 B.n463 B.n462 10.6151
R1770 B.n463 B.n128 10.6151
R1771 B.n467 B.n128 10.6151
R1772 B.n468 B.n467 10.6151
R1773 B.n469 B.n468 10.6151
R1774 B.n469 B.n126 10.6151
R1775 B.n473 B.n126 10.6151
R1776 B.n474 B.n473 10.6151
R1777 B.n475 B.n474 10.6151
R1778 B.n475 B.n124 10.6151
R1779 B.n479 B.n124 10.6151
R1780 B.n480 B.n479 10.6151
R1781 B.n481 B.n480 10.6151
R1782 B.n481 B.n122 10.6151
R1783 B.n485 B.n122 10.6151
R1784 B.n486 B.n485 10.6151
R1785 B.n487 B.n486 10.6151
R1786 B.n487 B.n120 10.6151
R1787 B.n491 B.n120 10.6151
R1788 B.n492 B.n491 10.6151
R1789 B.n493 B.n492 10.6151
R1790 B.n493 B.n118 10.6151
R1791 B.n497 B.n118 10.6151
R1792 B.n498 B.n497 10.6151
R1793 B.n499 B.n498 10.6151
R1794 B.n499 B.n116 10.6151
R1795 B.n503 B.n116 10.6151
R1796 B.n504 B.n503 10.6151
R1797 B.n505 B.n504 10.6151
R1798 B.n505 B.n114 10.6151
R1799 B.n509 B.n114 10.6151
R1800 B.n510 B.n509 10.6151
R1801 B.n511 B.n510 10.6151
R1802 B.n511 B.n112 10.6151
R1803 B.n515 B.n112 10.6151
R1804 B.n516 B.n515 10.6151
R1805 B.n517 B.n516 10.6151
R1806 B.n517 B.n110 10.6151
R1807 B.n521 B.n110 10.6151
R1808 B.n522 B.n521 10.6151
R1809 B.n523 B.n522 10.6151
R1810 B.n523 B.n108 10.6151
R1811 B.n527 B.n108 10.6151
R1812 B.n528 B.n527 10.6151
R1813 B.n529 B.n528 10.6151
R1814 B.n529 B.n106 10.6151
R1815 B.n533 B.n106 10.6151
R1816 B.n534 B.n533 10.6151
R1817 B.n535 B.n534 10.6151
R1818 B.n535 B.n104 10.6151
R1819 B.n539 B.n104 10.6151
R1820 B.n540 B.n539 10.6151
R1821 B.n541 B.n540 10.6151
R1822 B.n541 B.n102 10.6151
R1823 B.n545 B.n102 10.6151
R1824 B.n546 B.n545 10.6151
R1825 B.n547 B.n546 10.6151
R1826 B.n547 B.n100 10.6151
R1827 B.n551 B.n100 10.6151
R1828 B.n552 B.n551 10.6151
R1829 B.n553 B.n552 10.6151
R1830 B.n553 B.n98 10.6151
R1831 B.n557 B.n98 10.6151
R1832 B.n558 B.n557 10.6151
R1833 B.n559 B.n558 10.6151
R1834 B.n559 B.n96 10.6151
R1835 B.n563 B.n96 10.6151
R1836 B.n564 B.n563 10.6151
R1837 B.n565 B.n564 10.6151
R1838 B.n565 B.n94 10.6151
R1839 B.n569 B.n94 10.6151
R1840 B.n570 B.n569 10.6151
R1841 B.n571 B.n570 10.6151
R1842 B.n571 B.n92 10.6151
R1843 B.n575 B.n92 10.6151
R1844 B.n576 B.n575 10.6151
R1845 B.n577 B.n576 10.6151
R1846 B.n577 B.n90 10.6151
R1847 B.n581 B.n90 10.6151
R1848 B.n582 B.n581 10.6151
R1849 B.n583 B.n582 10.6151
R1850 B.n583 B.n88 10.6151
R1851 B.n587 B.n88 10.6151
R1852 B.n588 B.n587 10.6151
R1853 B.n589 B.n588 10.6151
R1854 B.n589 B.n86 10.6151
R1855 B.n593 B.n86 10.6151
R1856 B.n594 B.n593 10.6151
R1857 B.n595 B.n594 10.6151
R1858 B.n595 B.n84 10.6151
R1859 B.n599 B.n84 10.6151
R1860 B.n600 B.n599 10.6151
R1861 B.n601 B.n600 10.6151
R1862 B.n601 B.n82 10.6151
R1863 B.n605 B.n82 10.6151
R1864 B.n606 B.n605 10.6151
R1865 B.n607 B.n606 10.6151
R1866 B.n607 B.n80 10.6151
R1867 B.n611 B.n80 10.6151
R1868 B.n612 B.n611 10.6151
R1869 B.n613 B.n612 10.6151
R1870 B.n613 B.n78 10.6151
R1871 B.n617 B.n78 10.6151
R1872 B.n618 B.n617 10.6151
R1873 B.n619 B.n618 10.6151
R1874 B.n619 B.n76 10.6151
R1875 B.n623 B.n76 10.6151
R1876 B.n624 B.n623 10.6151
R1877 B.n625 B.n624 10.6151
R1878 B.n625 B.n74 10.6151
R1879 B.n629 B.n74 10.6151
R1880 B.n630 B.n629 10.6151
R1881 B.n631 B.n630 10.6151
R1882 B.n324 B.n323 10.6151
R1883 B.n325 B.n324 10.6151
R1884 B.n325 B.n178 10.6151
R1885 B.n329 B.n178 10.6151
R1886 B.n330 B.n329 10.6151
R1887 B.n331 B.n330 10.6151
R1888 B.n331 B.n176 10.6151
R1889 B.n335 B.n176 10.6151
R1890 B.n336 B.n335 10.6151
R1891 B.n337 B.n336 10.6151
R1892 B.n337 B.n174 10.6151
R1893 B.n341 B.n174 10.6151
R1894 B.n342 B.n341 10.6151
R1895 B.n343 B.n342 10.6151
R1896 B.n343 B.n172 10.6151
R1897 B.n347 B.n172 10.6151
R1898 B.n348 B.n347 10.6151
R1899 B.n349 B.n348 10.6151
R1900 B.n349 B.n170 10.6151
R1901 B.n353 B.n170 10.6151
R1902 B.n354 B.n353 10.6151
R1903 B.n355 B.n354 10.6151
R1904 B.n355 B.n168 10.6151
R1905 B.n359 B.n168 10.6151
R1906 B.n360 B.n359 10.6151
R1907 B.n362 B.n164 10.6151
R1908 B.n366 B.n164 10.6151
R1909 B.n367 B.n366 10.6151
R1910 B.n368 B.n367 10.6151
R1911 B.n368 B.n162 10.6151
R1912 B.n372 B.n162 10.6151
R1913 B.n373 B.n372 10.6151
R1914 B.n374 B.n373 10.6151
R1915 B.n378 B.n377 10.6151
R1916 B.n379 B.n378 10.6151
R1917 B.n379 B.n156 10.6151
R1918 B.n383 B.n156 10.6151
R1919 B.n384 B.n383 10.6151
R1920 B.n385 B.n384 10.6151
R1921 B.n385 B.n154 10.6151
R1922 B.n389 B.n154 10.6151
R1923 B.n390 B.n389 10.6151
R1924 B.n391 B.n390 10.6151
R1925 B.n391 B.n152 10.6151
R1926 B.n395 B.n152 10.6151
R1927 B.n396 B.n395 10.6151
R1928 B.n397 B.n396 10.6151
R1929 B.n397 B.n150 10.6151
R1930 B.n401 B.n150 10.6151
R1931 B.n402 B.n401 10.6151
R1932 B.n403 B.n402 10.6151
R1933 B.n403 B.n148 10.6151
R1934 B.n407 B.n148 10.6151
R1935 B.n408 B.n407 10.6151
R1936 B.n409 B.n408 10.6151
R1937 B.n409 B.n146 10.6151
R1938 B.n413 B.n146 10.6151
R1939 B.n414 B.n413 10.6151
R1940 B.n319 B.n180 10.6151
R1941 B.n319 B.n318 10.6151
R1942 B.n318 B.n317 10.6151
R1943 B.n317 B.n182 10.6151
R1944 B.n313 B.n182 10.6151
R1945 B.n313 B.n312 10.6151
R1946 B.n312 B.n311 10.6151
R1947 B.n311 B.n184 10.6151
R1948 B.n307 B.n184 10.6151
R1949 B.n307 B.n306 10.6151
R1950 B.n306 B.n305 10.6151
R1951 B.n305 B.n186 10.6151
R1952 B.n301 B.n186 10.6151
R1953 B.n301 B.n300 10.6151
R1954 B.n300 B.n299 10.6151
R1955 B.n299 B.n188 10.6151
R1956 B.n295 B.n188 10.6151
R1957 B.n295 B.n294 10.6151
R1958 B.n294 B.n293 10.6151
R1959 B.n293 B.n190 10.6151
R1960 B.n289 B.n190 10.6151
R1961 B.n289 B.n288 10.6151
R1962 B.n288 B.n287 10.6151
R1963 B.n287 B.n192 10.6151
R1964 B.n283 B.n192 10.6151
R1965 B.n283 B.n282 10.6151
R1966 B.n282 B.n281 10.6151
R1967 B.n281 B.n194 10.6151
R1968 B.n277 B.n194 10.6151
R1969 B.n277 B.n276 10.6151
R1970 B.n276 B.n275 10.6151
R1971 B.n275 B.n196 10.6151
R1972 B.n271 B.n196 10.6151
R1973 B.n271 B.n270 10.6151
R1974 B.n270 B.n269 10.6151
R1975 B.n269 B.n198 10.6151
R1976 B.n265 B.n198 10.6151
R1977 B.n265 B.n264 10.6151
R1978 B.n264 B.n263 10.6151
R1979 B.n263 B.n200 10.6151
R1980 B.n259 B.n200 10.6151
R1981 B.n259 B.n258 10.6151
R1982 B.n258 B.n257 10.6151
R1983 B.n257 B.n202 10.6151
R1984 B.n253 B.n202 10.6151
R1985 B.n253 B.n252 10.6151
R1986 B.n252 B.n251 10.6151
R1987 B.n251 B.n204 10.6151
R1988 B.n247 B.n204 10.6151
R1989 B.n247 B.n246 10.6151
R1990 B.n246 B.n245 10.6151
R1991 B.n245 B.n206 10.6151
R1992 B.n241 B.n206 10.6151
R1993 B.n241 B.n240 10.6151
R1994 B.n240 B.n239 10.6151
R1995 B.n239 B.n208 10.6151
R1996 B.n235 B.n208 10.6151
R1997 B.n235 B.n234 10.6151
R1998 B.n234 B.n233 10.6151
R1999 B.n233 B.n210 10.6151
R2000 B.n229 B.n210 10.6151
R2001 B.n229 B.n228 10.6151
R2002 B.n228 B.n227 10.6151
R2003 B.n227 B.n212 10.6151
R2004 B.n223 B.n212 10.6151
R2005 B.n223 B.n222 10.6151
R2006 B.n222 B.n221 10.6151
R2007 B.n221 B.n214 10.6151
R2008 B.n217 B.n214 10.6151
R2009 B.n217 B.n216 10.6151
R2010 B.n216 B.n0 10.6151
R2011 B.n831 B.n1 10.6151
R2012 B.n831 B.n830 10.6151
R2013 B.n830 B.n829 10.6151
R2014 B.n829 B.n4 10.6151
R2015 B.n825 B.n4 10.6151
R2016 B.n825 B.n824 10.6151
R2017 B.n824 B.n823 10.6151
R2018 B.n823 B.n6 10.6151
R2019 B.n819 B.n6 10.6151
R2020 B.n819 B.n818 10.6151
R2021 B.n818 B.n817 10.6151
R2022 B.n817 B.n8 10.6151
R2023 B.n813 B.n8 10.6151
R2024 B.n813 B.n812 10.6151
R2025 B.n812 B.n811 10.6151
R2026 B.n811 B.n10 10.6151
R2027 B.n807 B.n10 10.6151
R2028 B.n807 B.n806 10.6151
R2029 B.n806 B.n805 10.6151
R2030 B.n805 B.n12 10.6151
R2031 B.n801 B.n12 10.6151
R2032 B.n801 B.n800 10.6151
R2033 B.n800 B.n799 10.6151
R2034 B.n799 B.n14 10.6151
R2035 B.n795 B.n14 10.6151
R2036 B.n795 B.n794 10.6151
R2037 B.n794 B.n793 10.6151
R2038 B.n793 B.n16 10.6151
R2039 B.n789 B.n16 10.6151
R2040 B.n789 B.n788 10.6151
R2041 B.n788 B.n787 10.6151
R2042 B.n787 B.n18 10.6151
R2043 B.n783 B.n18 10.6151
R2044 B.n783 B.n782 10.6151
R2045 B.n782 B.n781 10.6151
R2046 B.n781 B.n20 10.6151
R2047 B.n777 B.n20 10.6151
R2048 B.n777 B.n776 10.6151
R2049 B.n776 B.n775 10.6151
R2050 B.n775 B.n22 10.6151
R2051 B.n771 B.n22 10.6151
R2052 B.n771 B.n770 10.6151
R2053 B.n770 B.n769 10.6151
R2054 B.n769 B.n24 10.6151
R2055 B.n765 B.n24 10.6151
R2056 B.n765 B.n764 10.6151
R2057 B.n764 B.n763 10.6151
R2058 B.n763 B.n26 10.6151
R2059 B.n759 B.n26 10.6151
R2060 B.n759 B.n758 10.6151
R2061 B.n758 B.n757 10.6151
R2062 B.n757 B.n28 10.6151
R2063 B.n753 B.n28 10.6151
R2064 B.n753 B.n752 10.6151
R2065 B.n752 B.n751 10.6151
R2066 B.n751 B.n30 10.6151
R2067 B.n747 B.n30 10.6151
R2068 B.n747 B.n746 10.6151
R2069 B.n746 B.n745 10.6151
R2070 B.n745 B.n32 10.6151
R2071 B.n741 B.n32 10.6151
R2072 B.n741 B.n740 10.6151
R2073 B.n740 B.n739 10.6151
R2074 B.n739 B.n34 10.6151
R2075 B.n735 B.n34 10.6151
R2076 B.n735 B.n734 10.6151
R2077 B.n734 B.n733 10.6151
R2078 B.n733 B.n36 10.6151
R2079 B.n729 B.n36 10.6151
R2080 B.n729 B.n728 10.6151
R2081 B.n728 B.n727 10.6151
R2082 B.n686 B.n685 6.5566
R2083 B.n673 B.n672 6.5566
R2084 B.n362 B.n361 6.5566
R2085 B.n374 B.n160 6.5566
R2086 B.n687 B.n686 4.05904
R2087 B.n672 B.n671 4.05904
R2088 B.n361 B.n360 4.05904
R2089 B.n377 B.n160 4.05904
R2090 B.n835 B.n0 2.81026
R2091 B.n835 B.n1 2.81026
C0 VTAIL VN 7.80301f
C1 B VN 1.39504f
C2 VP VDD1 6.89078f
C3 VP w_n5302_n2292# 12.136401f
C4 VP VDD2 0.670335f
C5 w_n5302_n2292# VDD1 2.67765f
C6 VDD2 VDD1 2.61697f
C7 w_n5302_n2292# VDD2 2.85655f
C8 VP VN 8.40059f
C9 VDD1 VN 0.155268f
C10 w_n5302_n2292# VN 11.444f
C11 VDD2 VN 6.37884f
C12 VTAIL B 2.73571f
C13 VTAIL VP 7.8172f
C14 VTAIL VDD1 8.44554f
C15 VTAIL w_n5302_n2292# 2.57236f
C16 VTAIL VDD2 8.50264f
C17 VP B 2.56309f
C18 B VDD1 2.31459f
C19 B w_n5302_n2292# 10.1887f
C20 B VDD2 2.45899f
C21 VDD2 VSUBS 2.376669f
C22 VDD1 VSUBS 2.117297f
C23 VTAIL VSUBS 0.765429f
C24 VN VSUBS 8.54943f
C25 VP VSUBS 4.645096f
C26 B VSUBS 5.757561f
C27 w_n5302_n2292# VSUBS 0.151361p
C28 B.n0 VSUBS 0.007128f
C29 B.n1 VSUBS 0.007128f
C30 B.n2 VSUBS 0.011272f
C31 B.n3 VSUBS 0.011272f
C32 B.n4 VSUBS 0.011272f
C33 B.n5 VSUBS 0.011272f
C34 B.n6 VSUBS 0.011272f
C35 B.n7 VSUBS 0.011272f
C36 B.n8 VSUBS 0.011272f
C37 B.n9 VSUBS 0.011272f
C38 B.n10 VSUBS 0.011272f
C39 B.n11 VSUBS 0.011272f
C40 B.n12 VSUBS 0.011272f
C41 B.n13 VSUBS 0.011272f
C42 B.n14 VSUBS 0.011272f
C43 B.n15 VSUBS 0.011272f
C44 B.n16 VSUBS 0.011272f
C45 B.n17 VSUBS 0.011272f
C46 B.n18 VSUBS 0.011272f
C47 B.n19 VSUBS 0.011272f
C48 B.n20 VSUBS 0.011272f
C49 B.n21 VSUBS 0.011272f
C50 B.n22 VSUBS 0.011272f
C51 B.n23 VSUBS 0.011272f
C52 B.n24 VSUBS 0.011272f
C53 B.n25 VSUBS 0.011272f
C54 B.n26 VSUBS 0.011272f
C55 B.n27 VSUBS 0.011272f
C56 B.n28 VSUBS 0.011272f
C57 B.n29 VSUBS 0.011272f
C58 B.n30 VSUBS 0.011272f
C59 B.n31 VSUBS 0.011272f
C60 B.n32 VSUBS 0.011272f
C61 B.n33 VSUBS 0.011272f
C62 B.n34 VSUBS 0.011272f
C63 B.n35 VSUBS 0.011272f
C64 B.n36 VSUBS 0.011272f
C65 B.n37 VSUBS 0.011272f
C66 B.n38 VSUBS 0.026047f
C67 B.n39 VSUBS 0.011272f
C68 B.n40 VSUBS 0.011272f
C69 B.n41 VSUBS 0.011272f
C70 B.n42 VSUBS 0.011272f
C71 B.n43 VSUBS 0.011272f
C72 B.n44 VSUBS 0.011272f
C73 B.n45 VSUBS 0.011272f
C74 B.n46 VSUBS 0.011272f
C75 B.n47 VSUBS 0.011272f
C76 B.n48 VSUBS 0.011272f
C77 B.n49 VSUBS 0.011272f
C78 B.n50 VSUBS 0.011272f
C79 B.n51 VSUBS 0.011272f
C80 B.t11 VSUBS 0.161711f
C81 B.t10 VSUBS 0.213632f
C82 B.t9 VSUBS 1.66444f
C83 B.n52 VSUBS 0.355154f
C84 B.n53 VSUBS 0.274918f
C85 B.n54 VSUBS 0.011272f
C86 B.n55 VSUBS 0.011272f
C87 B.n56 VSUBS 0.011272f
C88 B.n57 VSUBS 0.011272f
C89 B.t2 VSUBS 0.161714f
C90 B.t1 VSUBS 0.213634f
C91 B.t0 VSUBS 1.66444f
C92 B.n58 VSUBS 0.355151f
C93 B.n59 VSUBS 0.274915f
C94 B.n60 VSUBS 0.011272f
C95 B.n61 VSUBS 0.011272f
C96 B.n62 VSUBS 0.011272f
C97 B.n63 VSUBS 0.011272f
C98 B.n64 VSUBS 0.011272f
C99 B.n65 VSUBS 0.011272f
C100 B.n66 VSUBS 0.011272f
C101 B.n67 VSUBS 0.011272f
C102 B.n68 VSUBS 0.011272f
C103 B.n69 VSUBS 0.011272f
C104 B.n70 VSUBS 0.011272f
C105 B.n71 VSUBS 0.011272f
C106 B.n72 VSUBS 0.024661f
C107 B.n73 VSUBS 0.011272f
C108 B.n74 VSUBS 0.011272f
C109 B.n75 VSUBS 0.011272f
C110 B.n76 VSUBS 0.011272f
C111 B.n77 VSUBS 0.011272f
C112 B.n78 VSUBS 0.011272f
C113 B.n79 VSUBS 0.011272f
C114 B.n80 VSUBS 0.011272f
C115 B.n81 VSUBS 0.011272f
C116 B.n82 VSUBS 0.011272f
C117 B.n83 VSUBS 0.011272f
C118 B.n84 VSUBS 0.011272f
C119 B.n85 VSUBS 0.011272f
C120 B.n86 VSUBS 0.011272f
C121 B.n87 VSUBS 0.011272f
C122 B.n88 VSUBS 0.011272f
C123 B.n89 VSUBS 0.011272f
C124 B.n90 VSUBS 0.011272f
C125 B.n91 VSUBS 0.011272f
C126 B.n92 VSUBS 0.011272f
C127 B.n93 VSUBS 0.011272f
C128 B.n94 VSUBS 0.011272f
C129 B.n95 VSUBS 0.011272f
C130 B.n96 VSUBS 0.011272f
C131 B.n97 VSUBS 0.011272f
C132 B.n98 VSUBS 0.011272f
C133 B.n99 VSUBS 0.011272f
C134 B.n100 VSUBS 0.011272f
C135 B.n101 VSUBS 0.011272f
C136 B.n102 VSUBS 0.011272f
C137 B.n103 VSUBS 0.011272f
C138 B.n104 VSUBS 0.011272f
C139 B.n105 VSUBS 0.011272f
C140 B.n106 VSUBS 0.011272f
C141 B.n107 VSUBS 0.011272f
C142 B.n108 VSUBS 0.011272f
C143 B.n109 VSUBS 0.011272f
C144 B.n110 VSUBS 0.011272f
C145 B.n111 VSUBS 0.011272f
C146 B.n112 VSUBS 0.011272f
C147 B.n113 VSUBS 0.011272f
C148 B.n114 VSUBS 0.011272f
C149 B.n115 VSUBS 0.011272f
C150 B.n116 VSUBS 0.011272f
C151 B.n117 VSUBS 0.011272f
C152 B.n118 VSUBS 0.011272f
C153 B.n119 VSUBS 0.011272f
C154 B.n120 VSUBS 0.011272f
C155 B.n121 VSUBS 0.011272f
C156 B.n122 VSUBS 0.011272f
C157 B.n123 VSUBS 0.011272f
C158 B.n124 VSUBS 0.011272f
C159 B.n125 VSUBS 0.011272f
C160 B.n126 VSUBS 0.011272f
C161 B.n127 VSUBS 0.011272f
C162 B.n128 VSUBS 0.011272f
C163 B.n129 VSUBS 0.011272f
C164 B.n130 VSUBS 0.011272f
C165 B.n131 VSUBS 0.011272f
C166 B.n132 VSUBS 0.011272f
C167 B.n133 VSUBS 0.011272f
C168 B.n134 VSUBS 0.011272f
C169 B.n135 VSUBS 0.011272f
C170 B.n136 VSUBS 0.011272f
C171 B.n137 VSUBS 0.011272f
C172 B.n138 VSUBS 0.011272f
C173 B.n139 VSUBS 0.011272f
C174 B.n140 VSUBS 0.011272f
C175 B.n141 VSUBS 0.011272f
C176 B.n142 VSUBS 0.011272f
C177 B.n143 VSUBS 0.011272f
C178 B.n144 VSUBS 0.011272f
C179 B.n145 VSUBS 0.026047f
C180 B.n146 VSUBS 0.011272f
C181 B.n147 VSUBS 0.011272f
C182 B.n148 VSUBS 0.011272f
C183 B.n149 VSUBS 0.011272f
C184 B.n150 VSUBS 0.011272f
C185 B.n151 VSUBS 0.011272f
C186 B.n152 VSUBS 0.011272f
C187 B.n153 VSUBS 0.011272f
C188 B.n154 VSUBS 0.011272f
C189 B.n155 VSUBS 0.011272f
C190 B.n156 VSUBS 0.011272f
C191 B.n157 VSUBS 0.011272f
C192 B.t4 VSUBS 0.161714f
C193 B.t5 VSUBS 0.213634f
C194 B.t3 VSUBS 1.66444f
C195 B.n158 VSUBS 0.355151f
C196 B.n159 VSUBS 0.274915f
C197 B.n160 VSUBS 0.026115f
C198 B.n161 VSUBS 0.011272f
C199 B.n162 VSUBS 0.011272f
C200 B.n163 VSUBS 0.011272f
C201 B.n164 VSUBS 0.011272f
C202 B.n165 VSUBS 0.011272f
C203 B.t7 VSUBS 0.161711f
C204 B.t8 VSUBS 0.213632f
C205 B.t6 VSUBS 1.66444f
C206 B.n166 VSUBS 0.355154f
C207 B.n167 VSUBS 0.274918f
C208 B.n168 VSUBS 0.011272f
C209 B.n169 VSUBS 0.011272f
C210 B.n170 VSUBS 0.011272f
C211 B.n171 VSUBS 0.011272f
C212 B.n172 VSUBS 0.011272f
C213 B.n173 VSUBS 0.011272f
C214 B.n174 VSUBS 0.011272f
C215 B.n175 VSUBS 0.011272f
C216 B.n176 VSUBS 0.011272f
C217 B.n177 VSUBS 0.011272f
C218 B.n178 VSUBS 0.011272f
C219 B.n179 VSUBS 0.011272f
C220 B.n180 VSUBS 0.025337f
C221 B.n181 VSUBS 0.011272f
C222 B.n182 VSUBS 0.011272f
C223 B.n183 VSUBS 0.011272f
C224 B.n184 VSUBS 0.011272f
C225 B.n185 VSUBS 0.011272f
C226 B.n186 VSUBS 0.011272f
C227 B.n187 VSUBS 0.011272f
C228 B.n188 VSUBS 0.011272f
C229 B.n189 VSUBS 0.011272f
C230 B.n190 VSUBS 0.011272f
C231 B.n191 VSUBS 0.011272f
C232 B.n192 VSUBS 0.011272f
C233 B.n193 VSUBS 0.011272f
C234 B.n194 VSUBS 0.011272f
C235 B.n195 VSUBS 0.011272f
C236 B.n196 VSUBS 0.011272f
C237 B.n197 VSUBS 0.011272f
C238 B.n198 VSUBS 0.011272f
C239 B.n199 VSUBS 0.011272f
C240 B.n200 VSUBS 0.011272f
C241 B.n201 VSUBS 0.011272f
C242 B.n202 VSUBS 0.011272f
C243 B.n203 VSUBS 0.011272f
C244 B.n204 VSUBS 0.011272f
C245 B.n205 VSUBS 0.011272f
C246 B.n206 VSUBS 0.011272f
C247 B.n207 VSUBS 0.011272f
C248 B.n208 VSUBS 0.011272f
C249 B.n209 VSUBS 0.011272f
C250 B.n210 VSUBS 0.011272f
C251 B.n211 VSUBS 0.011272f
C252 B.n212 VSUBS 0.011272f
C253 B.n213 VSUBS 0.011272f
C254 B.n214 VSUBS 0.011272f
C255 B.n215 VSUBS 0.011272f
C256 B.n216 VSUBS 0.011272f
C257 B.n217 VSUBS 0.011272f
C258 B.n218 VSUBS 0.011272f
C259 B.n219 VSUBS 0.011272f
C260 B.n220 VSUBS 0.011272f
C261 B.n221 VSUBS 0.011272f
C262 B.n222 VSUBS 0.011272f
C263 B.n223 VSUBS 0.011272f
C264 B.n224 VSUBS 0.011272f
C265 B.n225 VSUBS 0.011272f
C266 B.n226 VSUBS 0.011272f
C267 B.n227 VSUBS 0.011272f
C268 B.n228 VSUBS 0.011272f
C269 B.n229 VSUBS 0.011272f
C270 B.n230 VSUBS 0.011272f
C271 B.n231 VSUBS 0.011272f
C272 B.n232 VSUBS 0.011272f
C273 B.n233 VSUBS 0.011272f
C274 B.n234 VSUBS 0.011272f
C275 B.n235 VSUBS 0.011272f
C276 B.n236 VSUBS 0.011272f
C277 B.n237 VSUBS 0.011272f
C278 B.n238 VSUBS 0.011272f
C279 B.n239 VSUBS 0.011272f
C280 B.n240 VSUBS 0.011272f
C281 B.n241 VSUBS 0.011272f
C282 B.n242 VSUBS 0.011272f
C283 B.n243 VSUBS 0.011272f
C284 B.n244 VSUBS 0.011272f
C285 B.n245 VSUBS 0.011272f
C286 B.n246 VSUBS 0.011272f
C287 B.n247 VSUBS 0.011272f
C288 B.n248 VSUBS 0.011272f
C289 B.n249 VSUBS 0.011272f
C290 B.n250 VSUBS 0.011272f
C291 B.n251 VSUBS 0.011272f
C292 B.n252 VSUBS 0.011272f
C293 B.n253 VSUBS 0.011272f
C294 B.n254 VSUBS 0.011272f
C295 B.n255 VSUBS 0.011272f
C296 B.n256 VSUBS 0.011272f
C297 B.n257 VSUBS 0.011272f
C298 B.n258 VSUBS 0.011272f
C299 B.n259 VSUBS 0.011272f
C300 B.n260 VSUBS 0.011272f
C301 B.n261 VSUBS 0.011272f
C302 B.n262 VSUBS 0.011272f
C303 B.n263 VSUBS 0.011272f
C304 B.n264 VSUBS 0.011272f
C305 B.n265 VSUBS 0.011272f
C306 B.n266 VSUBS 0.011272f
C307 B.n267 VSUBS 0.011272f
C308 B.n268 VSUBS 0.011272f
C309 B.n269 VSUBS 0.011272f
C310 B.n270 VSUBS 0.011272f
C311 B.n271 VSUBS 0.011272f
C312 B.n272 VSUBS 0.011272f
C313 B.n273 VSUBS 0.011272f
C314 B.n274 VSUBS 0.011272f
C315 B.n275 VSUBS 0.011272f
C316 B.n276 VSUBS 0.011272f
C317 B.n277 VSUBS 0.011272f
C318 B.n278 VSUBS 0.011272f
C319 B.n279 VSUBS 0.011272f
C320 B.n280 VSUBS 0.011272f
C321 B.n281 VSUBS 0.011272f
C322 B.n282 VSUBS 0.011272f
C323 B.n283 VSUBS 0.011272f
C324 B.n284 VSUBS 0.011272f
C325 B.n285 VSUBS 0.011272f
C326 B.n286 VSUBS 0.011272f
C327 B.n287 VSUBS 0.011272f
C328 B.n288 VSUBS 0.011272f
C329 B.n289 VSUBS 0.011272f
C330 B.n290 VSUBS 0.011272f
C331 B.n291 VSUBS 0.011272f
C332 B.n292 VSUBS 0.011272f
C333 B.n293 VSUBS 0.011272f
C334 B.n294 VSUBS 0.011272f
C335 B.n295 VSUBS 0.011272f
C336 B.n296 VSUBS 0.011272f
C337 B.n297 VSUBS 0.011272f
C338 B.n298 VSUBS 0.011272f
C339 B.n299 VSUBS 0.011272f
C340 B.n300 VSUBS 0.011272f
C341 B.n301 VSUBS 0.011272f
C342 B.n302 VSUBS 0.011272f
C343 B.n303 VSUBS 0.011272f
C344 B.n304 VSUBS 0.011272f
C345 B.n305 VSUBS 0.011272f
C346 B.n306 VSUBS 0.011272f
C347 B.n307 VSUBS 0.011272f
C348 B.n308 VSUBS 0.011272f
C349 B.n309 VSUBS 0.011272f
C350 B.n310 VSUBS 0.011272f
C351 B.n311 VSUBS 0.011272f
C352 B.n312 VSUBS 0.011272f
C353 B.n313 VSUBS 0.011272f
C354 B.n314 VSUBS 0.011272f
C355 B.n315 VSUBS 0.011272f
C356 B.n316 VSUBS 0.011272f
C357 B.n317 VSUBS 0.011272f
C358 B.n318 VSUBS 0.011272f
C359 B.n319 VSUBS 0.011272f
C360 B.n320 VSUBS 0.011272f
C361 B.n321 VSUBS 0.025337f
C362 B.n322 VSUBS 0.026047f
C363 B.n323 VSUBS 0.026047f
C364 B.n324 VSUBS 0.011272f
C365 B.n325 VSUBS 0.011272f
C366 B.n326 VSUBS 0.011272f
C367 B.n327 VSUBS 0.011272f
C368 B.n328 VSUBS 0.011272f
C369 B.n329 VSUBS 0.011272f
C370 B.n330 VSUBS 0.011272f
C371 B.n331 VSUBS 0.011272f
C372 B.n332 VSUBS 0.011272f
C373 B.n333 VSUBS 0.011272f
C374 B.n334 VSUBS 0.011272f
C375 B.n335 VSUBS 0.011272f
C376 B.n336 VSUBS 0.011272f
C377 B.n337 VSUBS 0.011272f
C378 B.n338 VSUBS 0.011272f
C379 B.n339 VSUBS 0.011272f
C380 B.n340 VSUBS 0.011272f
C381 B.n341 VSUBS 0.011272f
C382 B.n342 VSUBS 0.011272f
C383 B.n343 VSUBS 0.011272f
C384 B.n344 VSUBS 0.011272f
C385 B.n345 VSUBS 0.011272f
C386 B.n346 VSUBS 0.011272f
C387 B.n347 VSUBS 0.011272f
C388 B.n348 VSUBS 0.011272f
C389 B.n349 VSUBS 0.011272f
C390 B.n350 VSUBS 0.011272f
C391 B.n351 VSUBS 0.011272f
C392 B.n352 VSUBS 0.011272f
C393 B.n353 VSUBS 0.011272f
C394 B.n354 VSUBS 0.011272f
C395 B.n355 VSUBS 0.011272f
C396 B.n356 VSUBS 0.011272f
C397 B.n357 VSUBS 0.011272f
C398 B.n358 VSUBS 0.011272f
C399 B.n359 VSUBS 0.011272f
C400 B.n360 VSUBS 0.007791f
C401 B.n361 VSUBS 0.026115f
C402 B.n362 VSUBS 0.009117f
C403 B.n363 VSUBS 0.011272f
C404 B.n364 VSUBS 0.011272f
C405 B.n365 VSUBS 0.011272f
C406 B.n366 VSUBS 0.011272f
C407 B.n367 VSUBS 0.011272f
C408 B.n368 VSUBS 0.011272f
C409 B.n369 VSUBS 0.011272f
C410 B.n370 VSUBS 0.011272f
C411 B.n371 VSUBS 0.011272f
C412 B.n372 VSUBS 0.011272f
C413 B.n373 VSUBS 0.011272f
C414 B.n374 VSUBS 0.009117f
C415 B.n375 VSUBS 0.011272f
C416 B.n376 VSUBS 0.011272f
C417 B.n377 VSUBS 0.007791f
C418 B.n378 VSUBS 0.011272f
C419 B.n379 VSUBS 0.011272f
C420 B.n380 VSUBS 0.011272f
C421 B.n381 VSUBS 0.011272f
C422 B.n382 VSUBS 0.011272f
C423 B.n383 VSUBS 0.011272f
C424 B.n384 VSUBS 0.011272f
C425 B.n385 VSUBS 0.011272f
C426 B.n386 VSUBS 0.011272f
C427 B.n387 VSUBS 0.011272f
C428 B.n388 VSUBS 0.011272f
C429 B.n389 VSUBS 0.011272f
C430 B.n390 VSUBS 0.011272f
C431 B.n391 VSUBS 0.011272f
C432 B.n392 VSUBS 0.011272f
C433 B.n393 VSUBS 0.011272f
C434 B.n394 VSUBS 0.011272f
C435 B.n395 VSUBS 0.011272f
C436 B.n396 VSUBS 0.011272f
C437 B.n397 VSUBS 0.011272f
C438 B.n398 VSUBS 0.011272f
C439 B.n399 VSUBS 0.011272f
C440 B.n400 VSUBS 0.011272f
C441 B.n401 VSUBS 0.011272f
C442 B.n402 VSUBS 0.011272f
C443 B.n403 VSUBS 0.011272f
C444 B.n404 VSUBS 0.011272f
C445 B.n405 VSUBS 0.011272f
C446 B.n406 VSUBS 0.011272f
C447 B.n407 VSUBS 0.011272f
C448 B.n408 VSUBS 0.011272f
C449 B.n409 VSUBS 0.011272f
C450 B.n410 VSUBS 0.011272f
C451 B.n411 VSUBS 0.011272f
C452 B.n412 VSUBS 0.011272f
C453 B.n413 VSUBS 0.011272f
C454 B.n414 VSUBS 0.026047f
C455 B.n415 VSUBS 0.025337f
C456 B.n416 VSUBS 0.025337f
C457 B.n417 VSUBS 0.011272f
C458 B.n418 VSUBS 0.011272f
C459 B.n419 VSUBS 0.011272f
C460 B.n420 VSUBS 0.011272f
C461 B.n421 VSUBS 0.011272f
C462 B.n422 VSUBS 0.011272f
C463 B.n423 VSUBS 0.011272f
C464 B.n424 VSUBS 0.011272f
C465 B.n425 VSUBS 0.011272f
C466 B.n426 VSUBS 0.011272f
C467 B.n427 VSUBS 0.011272f
C468 B.n428 VSUBS 0.011272f
C469 B.n429 VSUBS 0.011272f
C470 B.n430 VSUBS 0.011272f
C471 B.n431 VSUBS 0.011272f
C472 B.n432 VSUBS 0.011272f
C473 B.n433 VSUBS 0.011272f
C474 B.n434 VSUBS 0.011272f
C475 B.n435 VSUBS 0.011272f
C476 B.n436 VSUBS 0.011272f
C477 B.n437 VSUBS 0.011272f
C478 B.n438 VSUBS 0.011272f
C479 B.n439 VSUBS 0.011272f
C480 B.n440 VSUBS 0.011272f
C481 B.n441 VSUBS 0.011272f
C482 B.n442 VSUBS 0.011272f
C483 B.n443 VSUBS 0.011272f
C484 B.n444 VSUBS 0.011272f
C485 B.n445 VSUBS 0.011272f
C486 B.n446 VSUBS 0.011272f
C487 B.n447 VSUBS 0.011272f
C488 B.n448 VSUBS 0.011272f
C489 B.n449 VSUBS 0.011272f
C490 B.n450 VSUBS 0.011272f
C491 B.n451 VSUBS 0.011272f
C492 B.n452 VSUBS 0.011272f
C493 B.n453 VSUBS 0.011272f
C494 B.n454 VSUBS 0.011272f
C495 B.n455 VSUBS 0.011272f
C496 B.n456 VSUBS 0.011272f
C497 B.n457 VSUBS 0.011272f
C498 B.n458 VSUBS 0.011272f
C499 B.n459 VSUBS 0.011272f
C500 B.n460 VSUBS 0.011272f
C501 B.n461 VSUBS 0.011272f
C502 B.n462 VSUBS 0.011272f
C503 B.n463 VSUBS 0.011272f
C504 B.n464 VSUBS 0.011272f
C505 B.n465 VSUBS 0.011272f
C506 B.n466 VSUBS 0.011272f
C507 B.n467 VSUBS 0.011272f
C508 B.n468 VSUBS 0.011272f
C509 B.n469 VSUBS 0.011272f
C510 B.n470 VSUBS 0.011272f
C511 B.n471 VSUBS 0.011272f
C512 B.n472 VSUBS 0.011272f
C513 B.n473 VSUBS 0.011272f
C514 B.n474 VSUBS 0.011272f
C515 B.n475 VSUBS 0.011272f
C516 B.n476 VSUBS 0.011272f
C517 B.n477 VSUBS 0.011272f
C518 B.n478 VSUBS 0.011272f
C519 B.n479 VSUBS 0.011272f
C520 B.n480 VSUBS 0.011272f
C521 B.n481 VSUBS 0.011272f
C522 B.n482 VSUBS 0.011272f
C523 B.n483 VSUBS 0.011272f
C524 B.n484 VSUBS 0.011272f
C525 B.n485 VSUBS 0.011272f
C526 B.n486 VSUBS 0.011272f
C527 B.n487 VSUBS 0.011272f
C528 B.n488 VSUBS 0.011272f
C529 B.n489 VSUBS 0.011272f
C530 B.n490 VSUBS 0.011272f
C531 B.n491 VSUBS 0.011272f
C532 B.n492 VSUBS 0.011272f
C533 B.n493 VSUBS 0.011272f
C534 B.n494 VSUBS 0.011272f
C535 B.n495 VSUBS 0.011272f
C536 B.n496 VSUBS 0.011272f
C537 B.n497 VSUBS 0.011272f
C538 B.n498 VSUBS 0.011272f
C539 B.n499 VSUBS 0.011272f
C540 B.n500 VSUBS 0.011272f
C541 B.n501 VSUBS 0.011272f
C542 B.n502 VSUBS 0.011272f
C543 B.n503 VSUBS 0.011272f
C544 B.n504 VSUBS 0.011272f
C545 B.n505 VSUBS 0.011272f
C546 B.n506 VSUBS 0.011272f
C547 B.n507 VSUBS 0.011272f
C548 B.n508 VSUBS 0.011272f
C549 B.n509 VSUBS 0.011272f
C550 B.n510 VSUBS 0.011272f
C551 B.n511 VSUBS 0.011272f
C552 B.n512 VSUBS 0.011272f
C553 B.n513 VSUBS 0.011272f
C554 B.n514 VSUBS 0.011272f
C555 B.n515 VSUBS 0.011272f
C556 B.n516 VSUBS 0.011272f
C557 B.n517 VSUBS 0.011272f
C558 B.n518 VSUBS 0.011272f
C559 B.n519 VSUBS 0.011272f
C560 B.n520 VSUBS 0.011272f
C561 B.n521 VSUBS 0.011272f
C562 B.n522 VSUBS 0.011272f
C563 B.n523 VSUBS 0.011272f
C564 B.n524 VSUBS 0.011272f
C565 B.n525 VSUBS 0.011272f
C566 B.n526 VSUBS 0.011272f
C567 B.n527 VSUBS 0.011272f
C568 B.n528 VSUBS 0.011272f
C569 B.n529 VSUBS 0.011272f
C570 B.n530 VSUBS 0.011272f
C571 B.n531 VSUBS 0.011272f
C572 B.n532 VSUBS 0.011272f
C573 B.n533 VSUBS 0.011272f
C574 B.n534 VSUBS 0.011272f
C575 B.n535 VSUBS 0.011272f
C576 B.n536 VSUBS 0.011272f
C577 B.n537 VSUBS 0.011272f
C578 B.n538 VSUBS 0.011272f
C579 B.n539 VSUBS 0.011272f
C580 B.n540 VSUBS 0.011272f
C581 B.n541 VSUBS 0.011272f
C582 B.n542 VSUBS 0.011272f
C583 B.n543 VSUBS 0.011272f
C584 B.n544 VSUBS 0.011272f
C585 B.n545 VSUBS 0.011272f
C586 B.n546 VSUBS 0.011272f
C587 B.n547 VSUBS 0.011272f
C588 B.n548 VSUBS 0.011272f
C589 B.n549 VSUBS 0.011272f
C590 B.n550 VSUBS 0.011272f
C591 B.n551 VSUBS 0.011272f
C592 B.n552 VSUBS 0.011272f
C593 B.n553 VSUBS 0.011272f
C594 B.n554 VSUBS 0.011272f
C595 B.n555 VSUBS 0.011272f
C596 B.n556 VSUBS 0.011272f
C597 B.n557 VSUBS 0.011272f
C598 B.n558 VSUBS 0.011272f
C599 B.n559 VSUBS 0.011272f
C600 B.n560 VSUBS 0.011272f
C601 B.n561 VSUBS 0.011272f
C602 B.n562 VSUBS 0.011272f
C603 B.n563 VSUBS 0.011272f
C604 B.n564 VSUBS 0.011272f
C605 B.n565 VSUBS 0.011272f
C606 B.n566 VSUBS 0.011272f
C607 B.n567 VSUBS 0.011272f
C608 B.n568 VSUBS 0.011272f
C609 B.n569 VSUBS 0.011272f
C610 B.n570 VSUBS 0.011272f
C611 B.n571 VSUBS 0.011272f
C612 B.n572 VSUBS 0.011272f
C613 B.n573 VSUBS 0.011272f
C614 B.n574 VSUBS 0.011272f
C615 B.n575 VSUBS 0.011272f
C616 B.n576 VSUBS 0.011272f
C617 B.n577 VSUBS 0.011272f
C618 B.n578 VSUBS 0.011272f
C619 B.n579 VSUBS 0.011272f
C620 B.n580 VSUBS 0.011272f
C621 B.n581 VSUBS 0.011272f
C622 B.n582 VSUBS 0.011272f
C623 B.n583 VSUBS 0.011272f
C624 B.n584 VSUBS 0.011272f
C625 B.n585 VSUBS 0.011272f
C626 B.n586 VSUBS 0.011272f
C627 B.n587 VSUBS 0.011272f
C628 B.n588 VSUBS 0.011272f
C629 B.n589 VSUBS 0.011272f
C630 B.n590 VSUBS 0.011272f
C631 B.n591 VSUBS 0.011272f
C632 B.n592 VSUBS 0.011272f
C633 B.n593 VSUBS 0.011272f
C634 B.n594 VSUBS 0.011272f
C635 B.n595 VSUBS 0.011272f
C636 B.n596 VSUBS 0.011272f
C637 B.n597 VSUBS 0.011272f
C638 B.n598 VSUBS 0.011272f
C639 B.n599 VSUBS 0.011272f
C640 B.n600 VSUBS 0.011272f
C641 B.n601 VSUBS 0.011272f
C642 B.n602 VSUBS 0.011272f
C643 B.n603 VSUBS 0.011272f
C644 B.n604 VSUBS 0.011272f
C645 B.n605 VSUBS 0.011272f
C646 B.n606 VSUBS 0.011272f
C647 B.n607 VSUBS 0.011272f
C648 B.n608 VSUBS 0.011272f
C649 B.n609 VSUBS 0.011272f
C650 B.n610 VSUBS 0.011272f
C651 B.n611 VSUBS 0.011272f
C652 B.n612 VSUBS 0.011272f
C653 B.n613 VSUBS 0.011272f
C654 B.n614 VSUBS 0.011272f
C655 B.n615 VSUBS 0.011272f
C656 B.n616 VSUBS 0.011272f
C657 B.n617 VSUBS 0.011272f
C658 B.n618 VSUBS 0.011272f
C659 B.n619 VSUBS 0.011272f
C660 B.n620 VSUBS 0.011272f
C661 B.n621 VSUBS 0.011272f
C662 B.n622 VSUBS 0.011272f
C663 B.n623 VSUBS 0.011272f
C664 B.n624 VSUBS 0.011272f
C665 B.n625 VSUBS 0.011272f
C666 B.n626 VSUBS 0.011272f
C667 B.n627 VSUBS 0.011272f
C668 B.n628 VSUBS 0.011272f
C669 B.n629 VSUBS 0.011272f
C670 B.n630 VSUBS 0.011272f
C671 B.n631 VSUBS 0.026724f
C672 B.n632 VSUBS 0.025337f
C673 B.n633 VSUBS 0.026047f
C674 B.n634 VSUBS 0.011272f
C675 B.n635 VSUBS 0.011272f
C676 B.n636 VSUBS 0.011272f
C677 B.n637 VSUBS 0.011272f
C678 B.n638 VSUBS 0.011272f
C679 B.n639 VSUBS 0.011272f
C680 B.n640 VSUBS 0.011272f
C681 B.n641 VSUBS 0.011272f
C682 B.n642 VSUBS 0.011272f
C683 B.n643 VSUBS 0.011272f
C684 B.n644 VSUBS 0.011272f
C685 B.n645 VSUBS 0.011272f
C686 B.n646 VSUBS 0.011272f
C687 B.n647 VSUBS 0.011272f
C688 B.n648 VSUBS 0.011272f
C689 B.n649 VSUBS 0.011272f
C690 B.n650 VSUBS 0.011272f
C691 B.n651 VSUBS 0.011272f
C692 B.n652 VSUBS 0.011272f
C693 B.n653 VSUBS 0.011272f
C694 B.n654 VSUBS 0.011272f
C695 B.n655 VSUBS 0.011272f
C696 B.n656 VSUBS 0.011272f
C697 B.n657 VSUBS 0.011272f
C698 B.n658 VSUBS 0.011272f
C699 B.n659 VSUBS 0.011272f
C700 B.n660 VSUBS 0.011272f
C701 B.n661 VSUBS 0.011272f
C702 B.n662 VSUBS 0.011272f
C703 B.n663 VSUBS 0.011272f
C704 B.n664 VSUBS 0.011272f
C705 B.n665 VSUBS 0.011272f
C706 B.n666 VSUBS 0.011272f
C707 B.n667 VSUBS 0.011272f
C708 B.n668 VSUBS 0.011272f
C709 B.n669 VSUBS 0.011272f
C710 B.n670 VSUBS 0.011272f
C711 B.n671 VSUBS 0.007791f
C712 B.n672 VSUBS 0.026115f
C713 B.n673 VSUBS 0.009117f
C714 B.n674 VSUBS 0.011272f
C715 B.n675 VSUBS 0.011272f
C716 B.n676 VSUBS 0.011272f
C717 B.n677 VSUBS 0.011272f
C718 B.n678 VSUBS 0.011272f
C719 B.n679 VSUBS 0.011272f
C720 B.n680 VSUBS 0.011272f
C721 B.n681 VSUBS 0.011272f
C722 B.n682 VSUBS 0.011272f
C723 B.n683 VSUBS 0.011272f
C724 B.n684 VSUBS 0.011272f
C725 B.n685 VSUBS 0.009117f
C726 B.n686 VSUBS 0.026115f
C727 B.n687 VSUBS 0.007791f
C728 B.n688 VSUBS 0.011272f
C729 B.n689 VSUBS 0.011272f
C730 B.n690 VSUBS 0.011272f
C731 B.n691 VSUBS 0.011272f
C732 B.n692 VSUBS 0.011272f
C733 B.n693 VSUBS 0.011272f
C734 B.n694 VSUBS 0.011272f
C735 B.n695 VSUBS 0.011272f
C736 B.n696 VSUBS 0.011272f
C737 B.n697 VSUBS 0.011272f
C738 B.n698 VSUBS 0.011272f
C739 B.n699 VSUBS 0.011272f
C740 B.n700 VSUBS 0.011272f
C741 B.n701 VSUBS 0.011272f
C742 B.n702 VSUBS 0.011272f
C743 B.n703 VSUBS 0.011272f
C744 B.n704 VSUBS 0.011272f
C745 B.n705 VSUBS 0.011272f
C746 B.n706 VSUBS 0.011272f
C747 B.n707 VSUBS 0.011272f
C748 B.n708 VSUBS 0.011272f
C749 B.n709 VSUBS 0.011272f
C750 B.n710 VSUBS 0.011272f
C751 B.n711 VSUBS 0.011272f
C752 B.n712 VSUBS 0.011272f
C753 B.n713 VSUBS 0.011272f
C754 B.n714 VSUBS 0.011272f
C755 B.n715 VSUBS 0.011272f
C756 B.n716 VSUBS 0.011272f
C757 B.n717 VSUBS 0.011272f
C758 B.n718 VSUBS 0.011272f
C759 B.n719 VSUBS 0.011272f
C760 B.n720 VSUBS 0.011272f
C761 B.n721 VSUBS 0.011272f
C762 B.n722 VSUBS 0.011272f
C763 B.n723 VSUBS 0.011272f
C764 B.n724 VSUBS 0.011272f
C765 B.n725 VSUBS 0.026047f
C766 B.n726 VSUBS 0.025337f
C767 B.n727 VSUBS 0.025337f
C768 B.n728 VSUBS 0.011272f
C769 B.n729 VSUBS 0.011272f
C770 B.n730 VSUBS 0.011272f
C771 B.n731 VSUBS 0.011272f
C772 B.n732 VSUBS 0.011272f
C773 B.n733 VSUBS 0.011272f
C774 B.n734 VSUBS 0.011272f
C775 B.n735 VSUBS 0.011272f
C776 B.n736 VSUBS 0.011272f
C777 B.n737 VSUBS 0.011272f
C778 B.n738 VSUBS 0.011272f
C779 B.n739 VSUBS 0.011272f
C780 B.n740 VSUBS 0.011272f
C781 B.n741 VSUBS 0.011272f
C782 B.n742 VSUBS 0.011272f
C783 B.n743 VSUBS 0.011272f
C784 B.n744 VSUBS 0.011272f
C785 B.n745 VSUBS 0.011272f
C786 B.n746 VSUBS 0.011272f
C787 B.n747 VSUBS 0.011272f
C788 B.n748 VSUBS 0.011272f
C789 B.n749 VSUBS 0.011272f
C790 B.n750 VSUBS 0.011272f
C791 B.n751 VSUBS 0.011272f
C792 B.n752 VSUBS 0.011272f
C793 B.n753 VSUBS 0.011272f
C794 B.n754 VSUBS 0.011272f
C795 B.n755 VSUBS 0.011272f
C796 B.n756 VSUBS 0.011272f
C797 B.n757 VSUBS 0.011272f
C798 B.n758 VSUBS 0.011272f
C799 B.n759 VSUBS 0.011272f
C800 B.n760 VSUBS 0.011272f
C801 B.n761 VSUBS 0.011272f
C802 B.n762 VSUBS 0.011272f
C803 B.n763 VSUBS 0.011272f
C804 B.n764 VSUBS 0.011272f
C805 B.n765 VSUBS 0.011272f
C806 B.n766 VSUBS 0.011272f
C807 B.n767 VSUBS 0.011272f
C808 B.n768 VSUBS 0.011272f
C809 B.n769 VSUBS 0.011272f
C810 B.n770 VSUBS 0.011272f
C811 B.n771 VSUBS 0.011272f
C812 B.n772 VSUBS 0.011272f
C813 B.n773 VSUBS 0.011272f
C814 B.n774 VSUBS 0.011272f
C815 B.n775 VSUBS 0.011272f
C816 B.n776 VSUBS 0.011272f
C817 B.n777 VSUBS 0.011272f
C818 B.n778 VSUBS 0.011272f
C819 B.n779 VSUBS 0.011272f
C820 B.n780 VSUBS 0.011272f
C821 B.n781 VSUBS 0.011272f
C822 B.n782 VSUBS 0.011272f
C823 B.n783 VSUBS 0.011272f
C824 B.n784 VSUBS 0.011272f
C825 B.n785 VSUBS 0.011272f
C826 B.n786 VSUBS 0.011272f
C827 B.n787 VSUBS 0.011272f
C828 B.n788 VSUBS 0.011272f
C829 B.n789 VSUBS 0.011272f
C830 B.n790 VSUBS 0.011272f
C831 B.n791 VSUBS 0.011272f
C832 B.n792 VSUBS 0.011272f
C833 B.n793 VSUBS 0.011272f
C834 B.n794 VSUBS 0.011272f
C835 B.n795 VSUBS 0.011272f
C836 B.n796 VSUBS 0.011272f
C837 B.n797 VSUBS 0.011272f
C838 B.n798 VSUBS 0.011272f
C839 B.n799 VSUBS 0.011272f
C840 B.n800 VSUBS 0.011272f
C841 B.n801 VSUBS 0.011272f
C842 B.n802 VSUBS 0.011272f
C843 B.n803 VSUBS 0.011272f
C844 B.n804 VSUBS 0.011272f
C845 B.n805 VSUBS 0.011272f
C846 B.n806 VSUBS 0.011272f
C847 B.n807 VSUBS 0.011272f
C848 B.n808 VSUBS 0.011272f
C849 B.n809 VSUBS 0.011272f
C850 B.n810 VSUBS 0.011272f
C851 B.n811 VSUBS 0.011272f
C852 B.n812 VSUBS 0.011272f
C853 B.n813 VSUBS 0.011272f
C854 B.n814 VSUBS 0.011272f
C855 B.n815 VSUBS 0.011272f
C856 B.n816 VSUBS 0.011272f
C857 B.n817 VSUBS 0.011272f
C858 B.n818 VSUBS 0.011272f
C859 B.n819 VSUBS 0.011272f
C860 B.n820 VSUBS 0.011272f
C861 B.n821 VSUBS 0.011272f
C862 B.n822 VSUBS 0.011272f
C863 B.n823 VSUBS 0.011272f
C864 B.n824 VSUBS 0.011272f
C865 B.n825 VSUBS 0.011272f
C866 B.n826 VSUBS 0.011272f
C867 B.n827 VSUBS 0.011272f
C868 B.n828 VSUBS 0.011272f
C869 B.n829 VSUBS 0.011272f
C870 B.n830 VSUBS 0.011272f
C871 B.n831 VSUBS 0.011272f
C872 B.n832 VSUBS 0.011272f
C873 B.n833 VSUBS 0.011272f
C874 B.n834 VSUBS 0.011272f
C875 B.n835 VSUBS 0.025523f
C876 VDD1.n0 VSUBS 0.036587f
C877 VDD1.n1 VSUBS 0.03422f
C878 VDD1.n2 VSUBS 0.018388f
C879 VDD1.n3 VSUBS 0.043463f
C880 VDD1.n4 VSUBS 0.01947f
C881 VDD1.n5 VSUBS 0.03422f
C882 VDD1.n6 VSUBS 0.018388f
C883 VDD1.n7 VSUBS 0.043463f
C884 VDD1.n8 VSUBS 0.01947f
C885 VDD1.n9 VSUBS 0.882167f
C886 VDD1.n10 VSUBS 0.018388f
C887 VDD1.t6 VSUBS 0.092852f
C888 VDD1.n11 VSUBS 0.157136f
C889 VDD1.n12 VSUBS 0.027644f
C890 VDD1.n13 VSUBS 0.032597f
C891 VDD1.n14 VSUBS 0.043463f
C892 VDD1.n15 VSUBS 0.01947f
C893 VDD1.n16 VSUBS 0.018388f
C894 VDD1.n17 VSUBS 0.03422f
C895 VDD1.n18 VSUBS 0.03422f
C896 VDD1.n19 VSUBS 0.018388f
C897 VDD1.n20 VSUBS 0.01947f
C898 VDD1.n21 VSUBS 0.043463f
C899 VDD1.n22 VSUBS 0.043463f
C900 VDD1.n23 VSUBS 0.01947f
C901 VDD1.n24 VSUBS 0.018388f
C902 VDD1.n25 VSUBS 0.03422f
C903 VDD1.n26 VSUBS 0.03422f
C904 VDD1.n27 VSUBS 0.018388f
C905 VDD1.n28 VSUBS 0.01947f
C906 VDD1.n29 VSUBS 0.043463f
C907 VDD1.n30 VSUBS 0.101767f
C908 VDD1.n31 VSUBS 0.01947f
C909 VDD1.n32 VSUBS 0.018388f
C910 VDD1.n33 VSUBS 0.074422f
C911 VDD1.n34 VSUBS 0.099819f
C912 VDD1.t7 VSUBS 0.179014f
C913 VDD1.t3 VSUBS 0.179014f
C914 VDD1.n35 VSUBS 1.21314f
C915 VDD1.n36 VSUBS 1.39373f
C916 VDD1.n37 VSUBS 0.036587f
C917 VDD1.n38 VSUBS 0.03422f
C918 VDD1.n39 VSUBS 0.018388f
C919 VDD1.n40 VSUBS 0.043463f
C920 VDD1.n41 VSUBS 0.01947f
C921 VDD1.n42 VSUBS 0.03422f
C922 VDD1.n43 VSUBS 0.018388f
C923 VDD1.n44 VSUBS 0.043463f
C924 VDD1.n45 VSUBS 0.01947f
C925 VDD1.n46 VSUBS 0.882167f
C926 VDD1.n47 VSUBS 0.018388f
C927 VDD1.t4 VSUBS 0.092852f
C928 VDD1.n48 VSUBS 0.157136f
C929 VDD1.n49 VSUBS 0.027644f
C930 VDD1.n50 VSUBS 0.032597f
C931 VDD1.n51 VSUBS 0.043463f
C932 VDD1.n52 VSUBS 0.01947f
C933 VDD1.n53 VSUBS 0.018388f
C934 VDD1.n54 VSUBS 0.03422f
C935 VDD1.n55 VSUBS 0.03422f
C936 VDD1.n56 VSUBS 0.018388f
C937 VDD1.n57 VSUBS 0.01947f
C938 VDD1.n58 VSUBS 0.043463f
C939 VDD1.n59 VSUBS 0.043463f
C940 VDD1.n60 VSUBS 0.01947f
C941 VDD1.n61 VSUBS 0.018388f
C942 VDD1.n62 VSUBS 0.03422f
C943 VDD1.n63 VSUBS 0.03422f
C944 VDD1.n64 VSUBS 0.018388f
C945 VDD1.n65 VSUBS 0.01947f
C946 VDD1.n66 VSUBS 0.043463f
C947 VDD1.n67 VSUBS 0.101767f
C948 VDD1.n68 VSUBS 0.01947f
C949 VDD1.n69 VSUBS 0.018388f
C950 VDD1.n70 VSUBS 0.074422f
C951 VDD1.n71 VSUBS 0.099819f
C952 VDD1.t2 VSUBS 0.179014f
C953 VDD1.t8 VSUBS 0.179014f
C954 VDD1.n72 VSUBS 1.21313f
C955 VDD1.n73 VSUBS 1.38231f
C956 VDD1.t9 VSUBS 0.179014f
C957 VDD1.t1 VSUBS 0.179014f
C958 VDD1.n74 VSUBS 1.24358f
C959 VDD1.n75 VSUBS 4.49598f
C960 VDD1.t5 VSUBS 0.179014f
C961 VDD1.t0 VSUBS 0.179014f
C962 VDD1.n76 VSUBS 1.21313f
C963 VDD1.n77 VSUBS 4.46079f
C964 VP.t8 VSUBS 2.00198f
C965 VP.n0 VSUBS 0.860976f
C966 VP.n1 VSUBS 0.034644f
C967 VP.n2 VSUBS 0.031309f
C968 VP.n3 VSUBS 0.034644f
C969 VP.t0 VSUBS 2.00198f
C970 VP.n4 VSUBS 0.734425f
C971 VP.n5 VSUBS 0.034644f
C972 VP.n6 VSUBS 0.045088f
C973 VP.n7 VSUBS 0.034644f
C974 VP.t1 VSUBS 2.00198f
C975 VP.n8 VSUBS 0.766954f
C976 VP.n9 VSUBS 0.034644f
C977 VP.n10 VSUBS 0.045088f
C978 VP.n11 VSUBS 0.034644f
C979 VP.t7 VSUBS 2.00198f
C980 VP.n12 VSUBS 0.734425f
C981 VP.n13 VSUBS 0.034644f
C982 VP.n14 VSUBS 0.031309f
C983 VP.n15 VSUBS 0.034644f
C984 VP.t5 VSUBS 2.00198f
C985 VP.n16 VSUBS 0.860976f
C986 VP.t9 VSUBS 2.00198f
C987 VP.n17 VSUBS 0.860976f
C988 VP.n18 VSUBS 0.034644f
C989 VP.n19 VSUBS 0.031309f
C990 VP.n20 VSUBS 0.034644f
C991 VP.t4 VSUBS 2.00198f
C992 VP.n21 VSUBS 0.734425f
C993 VP.n22 VSUBS 0.034644f
C994 VP.n23 VSUBS 0.045088f
C995 VP.n24 VSUBS 0.034644f
C996 VP.t6 VSUBS 2.00198f
C997 VP.n25 VSUBS 0.766954f
C998 VP.n26 VSUBS 0.034644f
C999 VP.n27 VSUBS 0.045088f
C1000 VP.n28 VSUBS 0.034644f
C1001 VP.t2 VSUBS 2.00198f
C1002 VP.n29 VSUBS 0.841302f
C1003 VP.t3 VSUBS 2.39159f
C1004 VP.n30 VSUBS 0.805537f
C1005 VP.n31 VSUBS 0.408113f
C1006 VP.n32 VSUBS 0.039506f
C1007 VP.n33 VSUBS 0.064244f
C1008 VP.n34 VSUBS 0.064244f
C1009 VP.n35 VSUBS 0.034644f
C1010 VP.n36 VSUBS 0.034644f
C1011 VP.n37 VSUBS 0.034644f
C1012 VP.n38 VSUBS 0.055632f
C1013 VP.n39 VSUBS 0.064244f
C1014 VP.n40 VSUBS 0.064244f
C1015 VP.n41 VSUBS 0.034644f
C1016 VP.n42 VSUBS 0.034644f
C1017 VP.n43 VSUBS 0.034644f
C1018 VP.n44 VSUBS 0.064244f
C1019 VP.n45 VSUBS 0.064244f
C1020 VP.n46 VSUBS 0.055632f
C1021 VP.n47 VSUBS 0.034644f
C1022 VP.n48 VSUBS 0.034644f
C1023 VP.n49 VSUBS 0.034644f
C1024 VP.n50 VSUBS 0.064244f
C1025 VP.n51 VSUBS 0.064244f
C1026 VP.n52 VSUBS 0.039506f
C1027 VP.n53 VSUBS 0.034644f
C1028 VP.n54 VSUBS 0.034644f
C1029 VP.n55 VSUBS 0.057266f
C1030 VP.n56 VSUBS 0.064244f
C1031 VP.n57 VSUBS 0.064244f
C1032 VP.n58 VSUBS 0.034644f
C1033 VP.n59 VSUBS 0.034644f
C1034 VP.n60 VSUBS 0.034644f
C1035 VP.n61 VSUBS 0.069412f
C1036 VP.n62 VSUBS 0.064244f
C1037 VP.n63 VSUBS 0.046483f
C1038 VP.n64 VSUBS 0.055905f
C1039 VP.n65 VSUBS 2.13097f
C1040 VP.n66 VSUBS 2.15463f
C1041 VP.n67 VSUBS 0.055905f
C1042 VP.n68 VSUBS 0.046483f
C1043 VP.n69 VSUBS 0.064244f
C1044 VP.n70 VSUBS 0.069412f
C1045 VP.n71 VSUBS 0.034644f
C1046 VP.n72 VSUBS 0.034644f
C1047 VP.n73 VSUBS 0.034644f
C1048 VP.n74 VSUBS 0.064244f
C1049 VP.n75 VSUBS 0.064244f
C1050 VP.n76 VSUBS 0.057266f
C1051 VP.n77 VSUBS 0.034644f
C1052 VP.n78 VSUBS 0.034644f
C1053 VP.n79 VSUBS 0.039506f
C1054 VP.n80 VSUBS 0.064244f
C1055 VP.n81 VSUBS 0.064244f
C1056 VP.n82 VSUBS 0.034644f
C1057 VP.n83 VSUBS 0.034644f
C1058 VP.n84 VSUBS 0.034644f
C1059 VP.n85 VSUBS 0.055632f
C1060 VP.n86 VSUBS 0.064244f
C1061 VP.n87 VSUBS 0.064244f
C1062 VP.n88 VSUBS 0.034644f
C1063 VP.n89 VSUBS 0.034644f
C1064 VP.n90 VSUBS 0.034644f
C1065 VP.n91 VSUBS 0.064244f
C1066 VP.n92 VSUBS 0.064244f
C1067 VP.n93 VSUBS 0.055632f
C1068 VP.n94 VSUBS 0.034644f
C1069 VP.n95 VSUBS 0.034644f
C1070 VP.n96 VSUBS 0.034644f
C1071 VP.n97 VSUBS 0.064244f
C1072 VP.n98 VSUBS 0.064244f
C1073 VP.n99 VSUBS 0.039506f
C1074 VP.n100 VSUBS 0.034644f
C1075 VP.n101 VSUBS 0.034644f
C1076 VP.n102 VSUBS 0.057266f
C1077 VP.n103 VSUBS 0.064244f
C1078 VP.n104 VSUBS 0.064244f
C1079 VP.n105 VSUBS 0.034644f
C1080 VP.n106 VSUBS 0.034644f
C1081 VP.n107 VSUBS 0.034644f
C1082 VP.n108 VSUBS 0.069412f
C1083 VP.n109 VSUBS 0.064244f
C1084 VP.n110 VSUBS 0.046483f
C1085 VP.n111 VSUBS 0.055905f
C1086 VP.n112 VSUBS 0.088453f
C1087 VDD2.n0 VSUBS 0.03679f
C1088 VDD2.n1 VSUBS 0.03441f
C1089 VDD2.n2 VSUBS 0.01849f
C1090 VDD2.n3 VSUBS 0.043704f
C1091 VDD2.n4 VSUBS 0.019578f
C1092 VDD2.n5 VSUBS 0.03441f
C1093 VDD2.n6 VSUBS 0.01849f
C1094 VDD2.n7 VSUBS 0.043704f
C1095 VDD2.n8 VSUBS 0.019578f
C1096 VDD2.n9 VSUBS 0.887062f
C1097 VDD2.n10 VSUBS 0.01849f
C1098 VDD2.t1 VSUBS 0.093368f
C1099 VDD2.n11 VSUBS 0.158008f
C1100 VDD2.n12 VSUBS 0.027797f
C1101 VDD2.n13 VSUBS 0.032778f
C1102 VDD2.n14 VSUBS 0.043704f
C1103 VDD2.n15 VSUBS 0.019578f
C1104 VDD2.n16 VSUBS 0.01849f
C1105 VDD2.n17 VSUBS 0.03441f
C1106 VDD2.n18 VSUBS 0.03441f
C1107 VDD2.n19 VSUBS 0.01849f
C1108 VDD2.n20 VSUBS 0.019578f
C1109 VDD2.n21 VSUBS 0.043704f
C1110 VDD2.n22 VSUBS 0.043704f
C1111 VDD2.n23 VSUBS 0.019578f
C1112 VDD2.n24 VSUBS 0.01849f
C1113 VDD2.n25 VSUBS 0.03441f
C1114 VDD2.n26 VSUBS 0.03441f
C1115 VDD2.n27 VSUBS 0.01849f
C1116 VDD2.n28 VSUBS 0.019578f
C1117 VDD2.n29 VSUBS 0.043704f
C1118 VDD2.n30 VSUBS 0.102332f
C1119 VDD2.n31 VSUBS 0.019578f
C1120 VDD2.n32 VSUBS 0.01849f
C1121 VDD2.n33 VSUBS 0.074835f
C1122 VDD2.n34 VSUBS 0.100373f
C1123 VDD2.t7 VSUBS 0.180008f
C1124 VDD2.t8 VSUBS 0.180008f
C1125 VDD2.n35 VSUBS 1.21986f
C1126 VDD2.n36 VSUBS 1.38998f
C1127 VDD2.t4 VSUBS 0.180008f
C1128 VDD2.t2 VSUBS 0.180008f
C1129 VDD2.n37 VSUBS 1.25048f
C1130 VDD2.n38 VSUBS 4.32971f
C1131 VDD2.n39 VSUBS 0.03679f
C1132 VDD2.n40 VSUBS 0.03441f
C1133 VDD2.n41 VSUBS 0.01849f
C1134 VDD2.n42 VSUBS 0.043704f
C1135 VDD2.n43 VSUBS 0.019578f
C1136 VDD2.n44 VSUBS 0.03441f
C1137 VDD2.n45 VSUBS 0.01849f
C1138 VDD2.n46 VSUBS 0.043704f
C1139 VDD2.n47 VSUBS 0.019578f
C1140 VDD2.n48 VSUBS 0.887062f
C1141 VDD2.n49 VSUBS 0.01849f
C1142 VDD2.t5 VSUBS 0.093368f
C1143 VDD2.n50 VSUBS 0.158008f
C1144 VDD2.n51 VSUBS 0.027797f
C1145 VDD2.n52 VSUBS 0.032778f
C1146 VDD2.n53 VSUBS 0.043704f
C1147 VDD2.n54 VSUBS 0.019578f
C1148 VDD2.n55 VSUBS 0.01849f
C1149 VDD2.n56 VSUBS 0.03441f
C1150 VDD2.n57 VSUBS 0.03441f
C1151 VDD2.n58 VSUBS 0.01849f
C1152 VDD2.n59 VSUBS 0.019578f
C1153 VDD2.n60 VSUBS 0.043704f
C1154 VDD2.n61 VSUBS 0.043704f
C1155 VDD2.n62 VSUBS 0.019578f
C1156 VDD2.n63 VSUBS 0.01849f
C1157 VDD2.n64 VSUBS 0.03441f
C1158 VDD2.n65 VSUBS 0.03441f
C1159 VDD2.n66 VSUBS 0.01849f
C1160 VDD2.n67 VSUBS 0.019578f
C1161 VDD2.n68 VSUBS 0.043704f
C1162 VDD2.n69 VSUBS 0.102332f
C1163 VDD2.n70 VSUBS 0.019578f
C1164 VDD2.n71 VSUBS 0.01849f
C1165 VDD2.n72 VSUBS 0.074835f
C1166 VDD2.n73 VSUBS 0.074958f
C1167 VDD2.n74 VSUBS 3.76656f
C1168 VDD2.t0 VSUBS 0.180008f
C1169 VDD2.t9 VSUBS 0.180008f
C1170 VDD2.n75 VSUBS 1.21987f
C1171 VDD2.n76 VSUBS 1.01826f
C1172 VDD2.t6 VSUBS 0.180008f
C1173 VDD2.t3 VSUBS 0.180008f
C1174 VDD2.n77 VSUBS 1.25043f
C1175 VTAIL.t8 VSUBS 0.175472f
C1176 VTAIL.t14 VSUBS 0.175472f
C1177 VTAIL.n0 VSUBS 1.05539f
C1178 VTAIL.n1 VSUBS 1.13152f
C1179 VTAIL.n2 VSUBS 0.035863f
C1180 VTAIL.n3 VSUBS 0.033542f
C1181 VTAIL.n4 VSUBS 0.018024f
C1182 VTAIL.n5 VSUBS 0.042603f
C1183 VTAIL.n6 VSUBS 0.019085f
C1184 VTAIL.n7 VSUBS 0.033542f
C1185 VTAIL.n8 VSUBS 0.018024f
C1186 VTAIL.n9 VSUBS 0.042603f
C1187 VTAIL.n10 VSUBS 0.019085f
C1188 VTAIL.n11 VSUBS 0.864708f
C1189 VTAIL.n12 VSUBS 0.018024f
C1190 VTAIL.t4 VSUBS 0.091015f
C1191 VTAIL.n13 VSUBS 0.154026f
C1192 VTAIL.n14 VSUBS 0.027097f
C1193 VTAIL.n15 VSUBS 0.031952f
C1194 VTAIL.n16 VSUBS 0.042603f
C1195 VTAIL.n17 VSUBS 0.019085f
C1196 VTAIL.n18 VSUBS 0.018024f
C1197 VTAIL.n19 VSUBS 0.033542f
C1198 VTAIL.n20 VSUBS 0.033542f
C1199 VTAIL.n21 VSUBS 0.018024f
C1200 VTAIL.n22 VSUBS 0.019085f
C1201 VTAIL.n23 VSUBS 0.042603f
C1202 VTAIL.n24 VSUBS 0.042603f
C1203 VTAIL.n25 VSUBS 0.019085f
C1204 VTAIL.n26 VSUBS 0.018024f
C1205 VTAIL.n27 VSUBS 0.033542f
C1206 VTAIL.n28 VSUBS 0.033542f
C1207 VTAIL.n29 VSUBS 0.018024f
C1208 VTAIL.n30 VSUBS 0.019085f
C1209 VTAIL.n31 VSUBS 0.042603f
C1210 VTAIL.n32 VSUBS 0.099753f
C1211 VTAIL.n33 VSUBS 0.019085f
C1212 VTAIL.n34 VSUBS 0.018024f
C1213 VTAIL.n35 VSUBS 0.07295f
C1214 VTAIL.n36 VSUBS 0.04987f
C1215 VTAIL.n37 VSUBS 0.58138f
C1216 VTAIL.t3 VSUBS 0.175472f
C1217 VTAIL.t5 VSUBS 0.175472f
C1218 VTAIL.n38 VSUBS 1.05539f
C1219 VTAIL.n39 VSUBS 1.32672f
C1220 VTAIL.t0 VSUBS 0.175472f
C1221 VTAIL.t19 VSUBS 0.175472f
C1222 VTAIL.n40 VSUBS 1.05539f
C1223 VTAIL.n41 VSUBS 2.73552f
C1224 VTAIL.t10 VSUBS 0.175472f
C1225 VTAIL.t9 VSUBS 0.175472f
C1226 VTAIL.n42 VSUBS 1.0554f
C1227 VTAIL.n43 VSUBS 2.73551f
C1228 VTAIL.t12 VSUBS 0.175472f
C1229 VTAIL.t13 VSUBS 0.175472f
C1230 VTAIL.n44 VSUBS 1.0554f
C1231 VTAIL.n45 VSUBS 1.32671f
C1232 VTAIL.n46 VSUBS 0.035863f
C1233 VTAIL.n47 VSUBS 0.033542f
C1234 VTAIL.n48 VSUBS 0.018024f
C1235 VTAIL.n49 VSUBS 0.042603f
C1236 VTAIL.n50 VSUBS 0.019085f
C1237 VTAIL.n51 VSUBS 0.033542f
C1238 VTAIL.n52 VSUBS 0.018024f
C1239 VTAIL.n53 VSUBS 0.042603f
C1240 VTAIL.n54 VSUBS 0.019085f
C1241 VTAIL.n55 VSUBS 0.864708f
C1242 VTAIL.n56 VSUBS 0.018024f
C1243 VTAIL.t16 VSUBS 0.091015f
C1244 VTAIL.n57 VSUBS 0.154026f
C1245 VTAIL.n58 VSUBS 0.027097f
C1246 VTAIL.n59 VSUBS 0.031952f
C1247 VTAIL.n60 VSUBS 0.042603f
C1248 VTAIL.n61 VSUBS 0.019085f
C1249 VTAIL.n62 VSUBS 0.018024f
C1250 VTAIL.n63 VSUBS 0.033542f
C1251 VTAIL.n64 VSUBS 0.033542f
C1252 VTAIL.n65 VSUBS 0.018024f
C1253 VTAIL.n66 VSUBS 0.019085f
C1254 VTAIL.n67 VSUBS 0.042603f
C1255 VTAIL.n68 VSUBS 0.042603f
C1256 VTAIL.n69 VSUBS 0.019085f
C1257 VTAIL.n70 VSUBS 0.018024f
C1258 VTAIL.n71 VSUBS 0.033542f
C1259 VTAIL.n72 VSUBS 0.033542f
C1260 VTAIL.n73 VSUBS 0.018024f
C1261 VTAIL.n74 VSUBS 0.019085f
C1262 VTAIL.n75 VSUBS 0.042603f
C1263 VTAIL.n76 VSUBS 0.099753f
C1264 VTAIL.n77 VSUBS 0.019085f
C1265 VTAIL.n78 VSUBS 0.018024f
C1266 VTAIL.n79 VSUBS 0.07295f
C1267 VTAIL.n80 VSUBS 0.04987f
C1268 VTAIL.n81 VSUBS 0.58138f
C1269 VTAIL.t18 VSUBS 0.175472f
C1270 VTAIL.t17 VSUBS 0.175472f
C1271 VTAIL.n82 VSUBS 1.0554f
C1272 VTAIL.n83 VSUBS 1.20931f
C1273 VTAIL.t2 VSUBS 0.175472f
C1274 VTAIL.t1 VSUBS 0.175472f
C1275 VTAIL.n84 VSUBS 1.0554f
C1276 VTAIL.n85 VSUBS 1.32671f
C1277 VTAIL.n86 VSUBS 0.035863f
C1278 VTAIL.n87 VSUBS 0.033542f
C1279 VTAIL.n88 VSUBS 0.018024f
C1280 VTAIL.n89 VSUBS 0.042603f
C1281 VTAIL.n90 VSUBS 0.019085f
C1282 VTAIL.n91 VSUBS 0.033542f
C1283 VTAIL.n92 VSUBS 0.018024f
C1284 VTAIL.n93 VSUBS 0.042603f
C1285 VTAIL.n94 VSUBS 0.019085f
C1286 VTAIL.n95 VSUBS 0.864708f
C1287 VTAIL.n96 VSUBS 0.018024f
C1288 VTAIL.t6 VSUBS 0.091015f
C1289 VTAIL.n97 VSUBS 0.154026f
C1290 VTAIL.n98 VSUBS 0.027097f
C1291 VTAIL.n99 VSUBS 0.031952f
C1292 VTAIL.n100 VSUBS 0.042603f
C1293 VTAIL.n101 VSUBS 0.019085f
C1294 VTAIL.n102 VSUBS 0.018024f
C1295 VTAIL.n103 VSUBS 0.033542f
C1296 VTAIL.n104 VSUBS 0.033542f
C1297 VTAIL.n105 VSUBS 0.018024f
C1298 VTAIL.n106 VSUBS 0.019085f
C1299 VTAIL.n107 VSUBS 0.042603f
C1300 VTAIL.n108 VSUBS 0.042603f
C1301 VTAIL.n109 VSUBS 0.019085f
C1302 VTAIL.n110 VSUBS 0.018024f
C1303 VTAIL.n111 VSUBS 0.033542f
C1304 VTAIL.n112 VSUBS 0.033542f
C1305 VTAIL.n113 VSUBS 0.018024f
C1306 VTAIL.n114 VSUBS 0.019085f
C1307 VTAIL.n115 VSUBS 0.042603f
C1308 VTAIL.n116 VSUBS 0.099753f
C1309 VTAIL.n117 VSUBS 0.019085f
C1310 VTAIL.n118 VSUBS 0.018024f
C1311 VTAIL.n119 VSUBS 0.07295f
C1312 VTAIL.n120 VSUBS 0.04987f
C1313 VTAIL.n121 VSUBS 1.77122f
C1314 VTAIL.n122 VSUBS 0.035863f
C1315 VTAIL.n123 VSUBS 0.033542f
C1316 VTAIL.n124 VSUBS 0.018024f
C1317 VTAIL.n125 VSUBS 0.042603f
C1318 VTAIL.n126 VSUBS 0.019085f
C1319 VTAIL.n127 VSUBS 0.033542f
C1320 VTAIL.n128 VSUBS 0.018024f
C1321 VTAIL.n129 VSUBS 0.042603f
C1322 VTAIL.n130 VSUBS 0.019085f
C1323 VTAIL.n131 VSUBS 0.864708f
C1324 VTAIL.n132 VSUBS 0.018024f
C1325 VTAIL.t7 VSUBS 0.091015f
C1326 VTAIL.n133 VSUBS 0.154026f
C1327 VTAIL.n134 VSUBS 0.027097f
C1328 VTAIL.n135 VSUBS 0.031952f
C1329 VTAIL.n136 VSUBS 0.042603f
C1330 VTAIL.n137 VSUBS 0.019085f
C1331 VTAIL.n138 VSUBS 0.018024f
C1332 VTAIL.n139 VSUBS 0.033542f
C1333 VTAIL.n140 VSUBS 0.033542f
C1334 VTAIL.n141 VSUBS 0.018024f
C1335 VTAIL.n142 VSUBS 0.019085f
C1336 VTAIL.n143 VSUBS 0.042603f
C1337 VTAIL.n144 VSUBS 0.042603f
C1338 VTAIL.n145 VSUBS 0.019085f
C1339 VTAIL.n146 VSUBS 0.018024f
C1340 VTAIL.n147 VSUBS 0.033542f
C1341 VTAIL.n148 VSUBS 0.033542f
C1342 VTAIL.n149 VSUBS 0.018024f
C1343 VTAIL.n150 VSUBS 0.019085f
C1344 VTAIL.n151 VSUBS 0.042603f
C1345 VTAIL.n152 VSUBS 0.099753f
C1346 VTAIL.n153 VSUBS 0.019085f
C1347 VTAIL.n154 VSUBS 0.018024f
C1348 VTAIL.n155 VSUBS 0.07295f
C1349 VTAIL.n156 VSUBS 0.04987f
C1350 VTAIL.n157 VSUBS 1.77122f
C1351 VTAIL.t15 VSUBS 0.175472f
C1352 VTAIL.t11 VSUBS 0.175472f
C1353 VTAIL.n158 VSUBS 1.05539f
C1354 VTAIL.n159 VSUBS 1.06816f
C1355 VN.t7 VSUBS 1.79841f
C1356 VN.n0 VSUBS 0.773426f
C1357 VN.n1 VSUBS 0.031121f
C1358 VN.n2 VSUBS 0.028125f
C1359 VN.n3 VSUBS 0.031121f
C1360 VN.t5 VSUBS 1.79841f
C1361 VN.n4 VSUBS 0.659744f
C1362 VN.n5 VSUBS 0.031121f
C1363 VN.n6 VSUBS 0.040503f
C1364 VN.n7 VSUBS 0.031121f
C1365 VN.t1 VSUBS 1.79841f
C1366 VN.n8 VSUBS 0.688965f
C1367 VN.n9 VSUBS 0.031121f
C1368 VN.n10 VSUBS 0.040503f
C1369 VN.n11 VSUBS 0.031121f
C1370 VN.t2 VSUBS 1.79841f
C1371 VN.n12 VSUBS 0.755753f
C1372 VN.t8 VSUBS 2.1484f
C1373 VN.n13 VSUBS 0.723624f
C1374 VN.n14 VSUBS 0.366613f
C1375 VN.n15 VSUBS 0.035488f
C1376 VN.n16 VSUBS 0.057711f
C1377 VN.n17 VSUBS 0.057711f
C1378 VN.n18 VSUBS 0.031121f
C1379 VN.n19 VSUBS 0.031121f
C1380 VN.n20 VSUBS 0.031121f
C1381 VN.n21 VSUBS 0.049975f
C1382 VN.n22 VSUBS 0.057711f
C1383 VN.n23 VSUBS 0.057711f
C1384 VN.n24 VSUBS 0.031121f
C1385 VN.n25 VSUBS 0.031121f
C1386 VN.n26 VSUBS 0.031121f
C1387 VN.n27 VSUBS 0.057711f
C1388 VN.n28 VSUBS 0.057711f
C1389 VN.n29 VSUBS 0.049975f
C1390 VN.n30 VSUBS 0.031121f
C1391 VN.n31 VSUBS 0.031121f
C1392 VN.n32 VSUBS 0.031121f
C1393 VN.n33 VSUBS 0.057711f
C1394 VN.n34 VSUBS 0.057711f
C1395 VN.n35 VSUBS 0.035488f
C1396 VN.n36 VSUBS 0.031121f
C1397 VN.n37 VSUBS 0.031121f
C1398 VN.n38 VSUBS 0.051443f
C1399 VN.n39 VSUBS 0.057711f
C1400 VN.n40 VSUBS 0.057711f
C1401 VN.n41 VSUBS 0.031121f
C1402 VN.n42 VSUBS 0.031121f
C1403 VN.n43 VSUBS 0.031121f
C1404 VN.n44 VSUBS 0.062353f
C1405 VN.n45 VSUBS 0.057711f
C1406 VN.n46 VSUBS 0.041756f
C1407 VN.n47 VSUBS 0.050221f
C1408 VN.n48 VSUBS 0.079458f
C1409 VN.t4 VSUBS 1.79841f
C1410 VN.n49 VSUBS 0.773426f
C1411 VN.n50 VSUBS 0.031121f
C1412 VN.n51 VSUBS 0.028125f
C1413 VN.n52 VSUBS 0.031121f
C1414 VN.t9 VSUBS 1.79841f
C1415 VN.n53 VSUBS 0.659744f
C1416 VN.n54 VSUBS 0.031121f
C1417 VN.n55 VSUBS 0.040503f
C1418 VN.n56 VSUBS 0.031121f
C1419 VN.t0 VSUBS 1.79841f
C1420 VN.n57 VSUBS 0.688965f
C1421 VN.n58 VSUBS 0.031121f
C1422 VN.n59 VSUBS 0.040503f
C1423 VN.n60 VSUBS 0.031121f
C1424 VN.t3 VSUBS 1.79841f
C1425 VN.n61 VSUBS 0.755753f
C1426 VN.t6 VSUBS 2.1484f
C1427 VN.n62 VSUBS 0.723624f
C1428 VN.n63 VSUBS 0.366613f
C1429 VN.n64 VSUBS 0.035488f
C1430 VN.n65 VSUBS 0.057711f
C1431 VN.n66 VSUBS 0.057711f
C1432 VN.n67 VSUBS 0.031121f
C1433 VN.n68 VSUBS 0.031121f
C1434 VN.n69 VSUBS 0.031121f
C1435 VN.n70 VSUBS 0.049975f
C1436 VN.n71 VSUBS 0.057711f
C1437 VN.n72 VSUBS 0.057711f
C1438 VN.n73 VSUBS 0.031121f
C1439 VN.n74 VSUBS 0.031121f
C1440 VN.n75 VSUBS 0.031121f
C1441 VN.n76 VSUBS 0.057711f
C1442 VN.n77 VSUBS 0.057711f
C1443 VN.n78 VSUBS 0.049975f
C1444 VN.n79 VSUBS 0.031121f
C1445 VN.n80 VSUBS 0.031121f
C1446 VN.n81 VSUBS 0.031121f
C1447 VN.n82 VSUBS 0.057711f
C1448 VN.n83 VSUBS 0.057711f
C1449 VN.n84 VSUBS 0.035488f
C1450 VN.n85 VSUBS 0.031121f
C1451 VN.n86 VSUBS 0.031121f
C1452 VN.n87 VSUBS 0.051443f
C1453 VN.n88 VSUBS 0.057711f
C1454 VN.n89 VSUBS 0.057711f
C1455 VN.n90 VSUBS 0.031121f
C1456 VN.n91 VSUBS 0.031121f
C1457 VN.n92 VSUBS 0.031121f
C1458 VN.n93 VSUBS 0.062353f
C1459 VN.n94 VSUBS 0.057711f
C1460 VN.n95 VSUBS 0.041756f
C1461 VN.n96 VSUBS 0.050221f
C1462 VN.n97 VSUBS 1.92678f
.ends

