* NGSPICE file created from diff_pair_sample_0065.ext - technology: sky130A

.subckt diff_pair_sample_0065 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X1 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X2 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=3.84
X3 VDD1.t1 VP.t1 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=3.84
X4 VDD1.t0 VP.t2 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=3.84
X5 VDD1.t6 VP.t3 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=3.84
X6 VTAIL.t19 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X7 VDD2.t6 VN.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=3.84
X8 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=3.84
X9 VTAIL.t2 VN.t4 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X10 VDD1.t5 VP.t4 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X11 VTAIL.t7 VN.t5 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X12 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=3.84
X13 VTAIL.t13 VP.t5 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X14 VDD2.t3 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X15 VDD1.t7 VP.t6 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=3.84
X16 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=3.84
X17 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=3.84
X18 VDD1.t4 VP.t7 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X19 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=3.84
X20 VTAIL.t10 VP.t8 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X21 VTAIL.t6 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X22 VTAIL.t9 VP.t9 VDD1.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=3.84
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=3.84
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n31 VP.t6 104.216
R60 VP.n75 VP.n74 85.5092
R61 VP.n130 VP.n0 85.5092
R62 VP.n73 VP.n18 85.5092
R63 VP.n75 VP.t2 71.0453
R64 VP.n89 VP.t9 71.0453
R65 VP.n102 VP.t7 71.0453
R66 VP.n115 VP.t5 71.0453
R67 VP.n0 VP.t1 71.0453
R68 VP.n18 VP.t3 71.0453
R69 VP.n58 VP.t8 71.0453
R70 VP.n45 VP.t4 71.0453
R71 VP.n32 VP.t0 71.0453
R72 VP.n74 VP.n73 59.4271
R73 VP.n96 VP.n95 56.4773
R74 VP.n109 VP.n108 56.4773
R75 VP.n52 VP.n51 56.4773
R76 VP.n39 VP.n38 56.4773
R77 VP.n32 VP.n31 54.3527
R78 VP.n82 VP.n81 40.8975
R79 VP.n122 VP.n2 40.8975
R80 VP.n65 VP.n20 40.8975
R81 VP.n83 VP.n82 39.9237
R82 VP.n122 VP.n121 39.9237
R83 VP.n65 VP.n64 39.9237
R84 VP.n77 VP.n76 24.3439
R85 VP.n77 VP.n16 24.3439
R86 VP.n81 VP.n16 24.3439
R87 VP.n83 VP.n14 24.3439
R88 VP.n87 VP.n14 24.3439
R89 VP.n88 VP.n87 24.3439
R90 VP.n90 VP.n12 24.3439
R91 VP.n94 VP.n12 24.3439
R92 VP.n95 VP.n94 24.3439
R93 VP.n96 VP.n10 24.3439
R94 VP.n100 VP.n10 24.3439
R95 VP.n101 VP.n100 24.3439
R96 VP.n103 VP.n8 24.3439
R97 VP.n107 VP.n8 24.3439
R98 VP.n108 VP.n107 24.3439
R99 VP.n109 VP.n6 24.3439
R100 VP.n113 VP.n6 24.3439
R101 VP.n114 VP.n113 24.3439
R102 VP.n116 VP.n4 24.3439
R103 VP.n120 VP.n4 24.3439
R104 VP.n121 VP.n120 24.3439
R105 VP.n126 VP.n2 24.3439
R106 VP.n127 VP.n126 24.3439
R107 VP.n128 VP.n127 24.3439
R108 VP.n69 VP.n20 24.3439
R109 VP.n70 VP.n69 24.3439
R110 VP.n71 VP.n70 24.3439
R111 VP.n52 VP.n24 24.3439
R112 VP.n56 VP.n24 24.3439
R113 VP.n57 VP.n56 24.3439
R114 VP.n59 VP.n22 24.3439
R115 VP.n63 VP.n22 24.3439
R116 VP.n64 VP.n63 24.3439
R117 VP.n39 VP.n28 24.3439
R118 VP.n43 VP.n28 24.3439
R119 VP.n44 VP.n43 24.3439
R120 VP.n46 VP.n26 24.3439
R121 VP.n50 VP.n26 24.3439
R122 VP.n51 VP.n50 24.3439
R123 VP.n33 VP.n30 24.3439
R124 VP.n37 VP.n30 24.3439
R125 VP.n38 VP.n37 24.3439
R126 VP.n90 VP.n89 20.449
R127 VP.n115 VP.n114 20.449
R128 VP.n58 VP.n57 20.449
R129 VP.n33 VP.n32 20.449
R130 VP.n102 VP.n101 12.1722
R131 VP.n103 VP.n102 12.1722
R132 VP.n45 VP.n44 12.1722
R133 VP.n46 VP.n45 12.1722
R134 VP.n76 VP.n75 4.38232
R135 VP.n128 VP.n0 4.38232
R136 VP.n71 VP.n18 4.38232
R137 VP.n89 VP.n88 3.89545
R138 VP.n116 VP.n115 3.89545
R139 VP.n59 VP.n58 3.89545
R140 VP.n34 VP.n31 2.44071
R141 VP.n73 VP.n72 0.355081
R142 VP.n74 VP.n17 0.355081
R143 VP.n130 VP.n129 0.355081
R144 VP VP.n130 0.26685
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VDD1.n56 VDD1.n0 289.615
R203 VDD1.n119 VDD1.n63 289.615
R204 VDD1.n57 VDD1.n56 185
R205 VDD1.n55 VDD1.n54 185
R206 VDD1.n4 VDD1.n3 185
R207 VDD1.n49 VDD1.n48 185
R208 VDD1.n47 VDD1.n46 185
R209 VDD1.n8 VDD1.n7 185
R210 VDD1.n12 VDD1.n10 185
R211 VDD1.n41 VDD1.n40 185
R212 VDD1.n39 VDD1.n38 185
R213 VDD1.n14 VDD1.n13 185
R214 VDD1.n33 VDD1.n32 185
R215 VDD1.n31 VDD1.n30 185
R216 VDD1.n18 VDD1.n17 185
R217 VDD1.n25 VDD1.n24 185
R218 VDD1.n23 VDD1.n22 185
R219 VDD1.n84 VDD1.n83 185
R220 VDD1.n86 VDD1.n85 185
R221 VDD1.n79 VDD1.n78 185
R222 VDD1.n92 VDD1.n91 185
R223 VDD1.n94 VDD1.n93 185
R224 VDD1.n75 VDD1.n74 185
R225 VDD1.n101 VDD1.n100 185
R226 VDD1.n102 VDD1.n73 185
R227 VDD1.n104 VDD1.n103 185
R228 VDD1.n71 VDD1.n70 185
R229 VDD1.n110 VDD1.n109 185
R230 VDD1.n112 VDD1.n111 185
R231 VDD1.n67 VDD1.n66 185
R232 VDD1.n118 VDD1.n117 185
R233 VDD1.n120 VDD1.n119 185
R234 VDD1.n21 VDD1.t7 149.524
R235 VDD1.n82 VDD1.t0 149.524
R236 VDD1.n56 VDD1.n55 104.615
R237 VDD1.n55 VDD1.n3 104.615
R238 VDD1.n48 VDD1.n3 104.615
R239 VDD1.n48 VDD1.n47 104.615
R240 VDD1.n47 VDD1.n7 104.615
R241 VDD1.n12 VDD1.n7 104.615
R242 VDD1.n40 VDD1.n12 104.615
R243 VDD1.n40 VDD1.n39 104.615
R244 VDD1.n39 VDD1.n13 104.615
R245 VDD1.n32 VDD1.n13 104.615
R246 VDD1.n32 VDD1.n31 104.615
R247 VDD1.n31 VDD1.n17 104.615
R248 VDD1.n24 VDD1.n17 104.615
R249 VDD1.n24 VDD1.n23 104.615
R250 VDD1.n85 VDD1.n84 104.615
R251 VDD1.n85 VDD1.n78 104.615
R252 VDD1.n92 VDD1.n78 104.615
R253 VDD1.n93 VDD1.n92 104.615
R254 VDD1.n93 VDD1.n74 104.615
R255 VDD1.n101 VDD1.n74 104.615
R256 VDD1.n102 VDD1.n101 104.615
R257 VDD1.n103 VDD1.n102 104.615
R258 VDD1.n103 VDD1.n70 104.615
R259 VDD1.n110 VDD1.n70 104.615
R260 VDD1.n111 VDD1.n110 104.615
R261 VDD1.n111 VDD1.n66 104.615
R262 VDD1.n118 VDD1.n66 104.615
R263 VDD1.n119 VDD1.n118 104.615
R264 VDD1.n127 VDD1.n126 63.179
R265 VDD1.n62 VDD1.n61 60.5384
R266 VDD1.n129 VDD1.n128 60.5382
R267 VDD1.n125 VDD1.n124 60.5382
R268 VDD1.n129 VDD1.n127 52.9298
R269 VDD1.n23 VDD1.t7 52.3082
R270 VDD1.n84 VDD1.t0 52.3082
R271 VDD1.n62 VDD1.n60 50.9074
R272 VDD1.n125 VDD1.n123 50.9074
R273 VDD1.n10 VDD1.n8 13.1884
R274 VDD1.n104 VDD1.n71 13.1884
R275 VDD1.n46 VDD1.n45 12.8005
R276 VDD1.n42 VDD1.n41 12.8005
R277 VDD1.n105 VDD1.n73 12.8005
R278 VDD1.n109 VDD1.n108 12.8005
R279 VDD1.n49 VDD1.n6 12.0247
R280 VDD1.n38 VDD1.n11 12.0247
R281 VDD1.n100 VDD1.n99 12.0247
R282 VDD1.n112 VDD1.n69 12.0247
R283 VDD1.n50 VDD1.n4 11.249
R284 VDD1.n37 VDD1.n14 11.249
R285 VDD1.n98 VDD1.n75 11.249
R286 VDD1.n113 VDD1.n67 11.249
R287 VDD1.n54 VDD1.n53 10.4732
R288 VDD1.n34 VDD1.n33 10.4732
R289 VDD1.n95 VDD1.n94 10.4732
R290 VDD1.n117 VDD1.n116 10.4732
R291 VDD1.n22 VDD1.n21 10.2747
R292 VDD1.n83 VDD1.n82 10.2747
R293 VDD1.n57 VDD1.n2 9.69747
R294 VDD1.n30 VDD1.n16 9.69747
R295 VDD1.n91 VDD1.n77 9.69747
R296 VDD1.n120 VDD1.n65 9.69747
R297 VDD1.n60 VDD1.n59 9.45567
R298 VDD1.n123 VDD1.n122 9.45567
R299 VDD1.n20 VDD1.n19 9.3005
R300 VDD1.n27 VDD1.n26 9.3005
R301 VDD1.n29 VDD1.n28 9.3005
R302 VDD1.n16 VDD1.n15 9.3005
R303 VDD1.n35 VDD1.n34 9.3005
R304 VDD1.n37 VDD1.n36 9.3005
R305 VDD1.n11 VDD1.n9 9.3005
R306 VDD1.n43 VDD1.n42 9.3005
R307 VDD1.n59 VDD1.n58 9.3005
R308 VDD1.n2 VDD1.n1 9.3005
R309 VDD1.n53 VDD1.n52 9.3005
R310 VDD1.n51 VDD1.n50 9.3005
R311 VDD1.n6 VDD1.n5 9.3005
R312 VDD1.n45 VDD1.n44 9.3005
R313 VDD1.n122 VDD1.n121 9.3005
R314 VDD1.n65 VDD1.n64 9.3005
R315 VDD1.n116 VDD1.n115 9.3005
R316 VDD1.n114 VDD1.n113 9.3005
R317 VDD1.n69 VDD1.n68 9.3005
R318 VDD1.n108 VDD1.n107 9.3005
R319 VDD1.n81 VDD1.n80 9.3005
R320 VDD1.n88 VDD1.n87 9.3005
R321 VDD1.n90 VDD1.n89 9.3005
R322 VDD1.n77 VDD1.n76 9.3005
R323 VDD1.n96 VDD1.n95 9.3005
R324 VDD1.n98 VDD1.n97 9.3005
R325 VDD1.n99 VDD1.n72 9.3005
R326 VDD1.n106 VDD1.n105 9.3005
R327 VDD1.n58 VDD1.n0 8.92171
R328 VDD1.n29 VDD1.n18 8.92171
R329 VDD1.n90 VDD1.n79 8.92171
R330 VDD1.n121 VDD1.n63 8.92171
R331 VDD1.n26 VDD1.n25 8.14595
R332 VDD1.n87 VDD1.n86 8.14595
R333 VDD1.n22 VDD1.n20 7.3702
R334 VDD1.n83 VDD1.n81 7.3702
R335 VDD1.n25 VDD1.n20 5.81868
R336 VDD1.n86 VDD1.n81 5.81868
R337 VDD1.n60 VDD1.n0 5.04292
R338 VDD1.n26 VDD1.n18 5.04292
R339 VDD1.n87 VDD1.n79 5.04292
R340 VDD1.n123 VDD1.n63 5.04292
R341 VDD1.n58 VDD1.n57 4.26717
R342 VDD1.n30 VDD1.n29 4.26717
R343 VDD1.n91 VDD1.n90 4.26717
R344 VDD1.n121 VDD1.n120 4.26717
R345 VDD1.n54 VDD1.n2 3.49141
R346 VDD1.n33 VDD1.n16 3.49141
R347 VDD1.n94 VDD1.n77 3.49141
R348 VDD1.n117 VDD1.n65 3.49141
R349 VDD1.n21 VDD1.n19 2.84303
R350 VDD1.n82 VDD1.n80 2.84303
R351 VDD1.n53 VDD1.n4 2.71565
R352 VDD1.n34 VDD1.n14 2.71565
R353 VDD1.n95 VDD1.n75 2.71565
R354 VDD1.n116 VDD1.n67 2.71565
R355 VDD1 VDD1.n129 2.63843
R356 VDD1.n50 VDD1.n49 1.93989
R357 VDD1.n38 VDD1.n37 1.93989
R358 VDD1.n100 VDD1.n98 1.93989
R359 VDD1.n113 VDD1.n112 1.93989
R360 VDD1.n128 VDD1.t3 1.74962
R361 VDD1.n128 VDD1.t6 1.74962
R362 VDD1.n61 VDD1.t2 1.74962
R363 VDD1.n61 VDD1.t5 1.74962
R364 VDD1.n126 VDD1.t8 1.74962
R365 VDD1.n126 VDD1.t1 1.74962
R366 VDD1.n124 VDD1.t9 1.74962
R367 VDD1.n124 VDD1.t4 1.74962
R368 VDD1.n46 VDD1.n6 1.16414
R369 VDD1.n41 VDD1.n11 1.16414
R370 VDD1.n99 VDD1.n73 1.16414
R371 VDD1.n109 VDD1.n69 1.16414
R372 VDD1 VDD1.n62 0.957397
R373 VDD1.n127 VDD1.n125 0.843861
R374 VDD1.n45 VDD1.n8 0.388379
R375 VDD1.n42 VDD1.n10 0.388379
R376 VDD1.n105 VDD1.n104 0.388379
R377 VDD1.n108 VDD1.n71 0.388379
R378 VDD1.n59 VDD1.n1 0.155672
R379 VDD1.n52 VDD1.n1 0.155672
R380 VDD1.n52 VDD1.n51 0.155672
R381 VDD1.n51 VDD1.n5 0.155672
R382 VDD1.n44 VDD1.n5 0.155672
R383 VDD1.n44 VDD1.n43 0.155672
R384 VDD1.n43 VDD1.n9 0.155672
R385 VDD1.n36 VDD1.n9 0.155672
R386 VDD1.n36 VDD1.n35 0.155672
R387 VDD1.n35 VDD1.n15 0.155672
R388 VDD1.n28 VDD1.n15 0.155672
R389 VDD1.n28 VDD1.n27 0.155672
R390 VDD1.n27 VDD1.n19 0.155672
R391 VDD1.n88 VDD1.n80 0.155672
R392 VDD1.n89 VDD1.n88 0.155672
R393 VDD1.n89 VDD1.n76 0.155672
R394 VDD1.n96 VDD1.n76 0.155672
R395 VDD1.n97 VDD1.n96 0.155672
R396 VDD1.n97 VDD1.n72 0.155672
R397 VDD1.n106 VDD1.n72 0.155672
R398 VDD1.n107 VDD1.n106 0.155672
R399 VDD1.n107 VDD1.n68 0.155672
R400 VDD1.n114 VDD1.n68 0.155672
R401 VDD1.n115 VDD1.n114 0.155672
R402 VDD1.n115 VDD1.n64 0.155672
R403 VDD1.n122 VDD1.n64 0.155672
R404 VTAIL.n256 VTAIL.n200 289.615
R405 VTAIL.n58 VTAIL.n2 289.615
R406 VTAIL.n194 VTAIL.n138 289.615
R407 VTAIL.n128 VTAIL.n72 289.615
R408 VTAIL.n221 VTAIL.n220 185
R409 VTAIL.n223 VTAIL.n222 185
R410 VTAIL.n216 VTAIL.n215 185
R411 VTAIL.n229 VTAIL.n228 185
R412 VTAIL.n231 VTAIL.n230 185
R413 VTAIL.n212 VTAIL.n211 185
R414 VTAIL.n238 VTAIL.n237 185
R415 VTAIL.n239 VTAIL.n210 185
R416 VTAIL.n241 VTAIL.n240 185
R417 VTAIL.n208 VTAIL.n207 185
R418 VTAIL.n247 VTAIL.n246 185
R419 VTAIL.n249 VTAIL.n248 185
R420 VTAIL.n204 VTAIL.n203 185
R421 VTAIL.n255 VTAIL.n254 185
R422 VTAIL.n257 VTAIL.n256 185
R423 VTAIL.n23 VTAIL.n22 185
R424 VTAIL.n25 VTAIL.n24 185
R425 VTAIL.n18 VTAIL.n17 185
R426 VTAIL.n31 VTAIL.n30 185
R427 VTAIL.n33 VTAIL.n32 185
R428 VTAIL.n14 VTAIL.n13 185
R429 VTAIL.n40 VTAIL.n39 185
R430 VTAIL.n41 VTAIL.n12 185
R431 VTAIL.n43 VTAIL.n42 185
R432 VTAIL.n10 VTAIL.n9 185
R433 VTAIL.n49 VTAIL.n48 185
R434 VTAIL.n51 VTAIL.n50 185
R435 VTAIL.n6 VTAIL.n5 185
R436 VTAIL.n57 VTAIL.n56 185
R437 VTAIL.n59 VTAIL.n58 185
R438 VTAIL.n195 VTAIL.n194 185
R439 VTAIL.n193 VTAIL.n192 185
R440 VTAIL.n142 VTAIL.n141 185
R441 VTAIL.n187 VTAIL.n186 185
R442 VTAIL.n185 VTAIL.n184 185
R443 VTAIL.n146 VTAIL.n145 185
R444 VTAIL.n150 VTAIL.n148 185
R445 VTAIL.n179 VTAIL.n178 185
R446 VTAIL.n177 VTAIL.n176 185
R447 VTAIL.n152 VTAIL.n151 185
R448 VTAIL.n171 VTAIL.n170 185
R449 VTAIL.n169 VTAIL.n168 185
R450 VTAIL.n156 VTAIL.n155 185
R451 VTAIL.n163 VTAIL.n162 185
R452 VTAIL.n161 VTAIL.n160 185
R453 VTAIL.n129 VTAIL.n128 185
R454 VTAIL.n127 VTAIL.n126 185
R455 VTAIL.n76 VTAIL.n75 185
R456 VTAIL.n121 VTAIL.n120 185
R457 VTAIL.n119 VTAIL.n118 185
R458 VTAIL.n80 VTAIL.n79 185
R459 VTAIL.n84 VTAIL.n82 185
R460 VTAIL.n113 VTAIL.n112 185
R461 VTAIL.n111 VTAIL.n110 185
R462 VTAIL.n86 VTAIL.n85 185
R463 VTAIL.n105 VTAIL.n104 185
R464 VTAIL.n103 VTAIL.n102 185
R465 VTAIL.n90 VTAIL.n89 185
R466 VTAIL.n97 VTAIL.n96 185
R467 VTAIL.n95 VTAIL.n94 185
R468 VTAIL.n219 VTAIL.t5 149.524
R469 VTAIL.n21 VTAIL.t17 149.524
R470 VTAIL.n159 VTAIL.t15 149.524
R471 VTAIL.n93 VTAIL.t3 149.524
R472 VTAIL.n222 VTAIL.n221 104.615
R473 VTAIL.n222 VTAIL.n215 104.615
R474 VTAIL.n229 VTAIL.n215 104.615
R475 VTAIL.n230 VTAIL.n229 104.615
R476 VTAIL.n230 VTAIL.n211 104.615
R477 VTAIL.n238 VTAIL.n211 104.615
R478 VTAIL.n239 VTAIL.n238 104.615
R479 VTAIL.n240 VTAIL.n239 104.615
R480 VTAIL.n240 VTAIL.n207 104.615
R481 VTAIL.n247 VTAIL.n207 104.615
R482 VTAIL.n248 VTAIL.n247 104.615
R483 VTAIL.n248 VTAIL.n203 104.615
R484 VTAIL.n255 VTAIL.n203 104.615
R485 VTAIL.n256 VTAIL.n255 104.615
R486 VTAIL.n24 VTAIL.n23 104.615
R487 VTAIL.n24 VTAIL.n17 104.615
R488 VTAIL.n31 VTAIL.n17 104.615
R489 VTAIL.n32 VTAIL.n31 104.615
R490 VTAIL.n32 VTAIL.n13 104.615
R491 VTAIL.n40 VTAIL.n13 104.615
R492 VTAIL.n41 VTAIL.n40 104.615
R493 VTAIL.n42 VTAIL.n41 104.615
R494 VTAIL.n42 VTAIL.n9 104.615
R495 VTAIL.n49 VTAIL.n9 104.615
R496 VTAIL.n50 VTAIL.n49 104.615
R497 VTAIL.n50 VTAIL.n5 104.615
R498 VTAIL.n57 VTAIL.n5 104.615
R499 VTAIL.n58 VTAIL.n57 104.615
R500 VTAIL.n194 VTAIL.n193 104.615
R501 VTAIL.n193 VTAIL.n141 104.615
R502 VTAIL.n186 VTAIL.n141 104.615
R503 VTAIL.n186 VTAIL.n185 104.615
R504 VTAIL.n185 VTAIL.n145 104.615
R505 VTAIL.n150 VTAIL.n145 104.615
R506 VTAIL.n178 VTAIL.n150 104.615
R507 VTAIL.n178 VTAIL.n177 104.615
R508 VTAIL.n177 VTAIL.n151 104.615
R509 VTAIL.n170 VTAIL.n151 104.615
R510 VTAIL.n170 VTAIL.n169 104.615
R511 VTAIL.n169 VTAIL.n155 104.615
R512 VTAIL.n162 VTAIL.n155 104.615
R513 VTAIL.n162 VTAIL.n161 104.615
R514 VTAIL.n128 VTAIL.n127 104.615
R515 VTAIL.n127 VTAIL.n75 104.615
R516 VTAIL.n120 VTAIL.n75 104.615
R517 VTAIL.n120 VTAIL.n119 104.615
R518 VTAIL.n119 VTAIL.n79 104.615
R519 VTAIL.n84 VTAIL.n79 104.615
R520 VTAIL.n112 VTAIL.n84 104.615
R521 VTAIL.n112 VTAIL.n111 104.615
R522 VTAIL.n111 VTAIL.n85 104.615
R523 VTAIL.n104 VTAIL.n85 104.615
R524 VTAIL.n104 VTAIL.n103 104.615
R525 VTAIL.n103 VTAIL.n89 104.615
R526 VTAIL.n96 VTAIL.n89 104.615
R527 VTAIL.n96 VTAIL.n95 104.615
R528 VTAIL.n221 VTAIL.t5 52.3082
R529 VTAIL.n23 VTAIL.t17 52.3082
R530 VTAIL.n161 VTAIL.t15 52.3082
R531 VTAIL.n95 VTAIL.t3 52.3082
R532 VTAIL.n137 VTAIL.n136 43.8596
R533 VTAIL.n135 VTAIL.n134 43.8596
R534 VTAIL.n71 VTAIL.n70 43.8596
R535 VTAIL.n69 VTAIL.n68 43.8596
R536 VTAIL.n263 VTAIL.n262 43.8594
R537 VTAIL.n1 VTAIL.n0 43.8594
R538 VTAIL.n65 VTAIL.n64 43.8594
R539 VTAIL.n67 VTAIL.n66 43.8594
R540 VTAIL.n261 VTAIL.n260 30.6338
R541 VTAIL.n63 VTAIL.n62 30.6338
R542 VTAIL.n199 VTAIL.n198 30.6338
R543 VTAIL.n133 VTAIL.n132 30.6338
R544 VTAIL.n69 VTAIL.n67 29.3152
R545 VTAIL.n261 VTAIL.n199 25.7203
R546 VTAIL.n241 VTAIL.n208 13.1884
R547 VTAIL.n43 VTAIL.n10 13.1884
R548 VTAIL.n148 VTAIL.n146 13.1884
R549 VTAIL.n82 VTAIL.n80 13.1884
R550 VTAIL.n242 VTAIL.n210 12.8005
R551 VTAIL.n246 VTAIL.n245 12.8005
R552 VTAIL.n44 VTAIL.n12 12.8005
R553 VTAIL.n48 VTAIL.n47 12.8005
R554 VTAIL.n184 VTAIL.n183 12.8005
R555 VTAIL.n180 VTAIL.n179 12.8005
R556 VTAIL.n118 VTAIL.n117 12.8005
R557 VTAIL.n114 VTAIL.n113 12.8005
R558 VTAIL.n237 VTAIL.n236 12.0247
R559 VTAIL.n249 VTAIL.n206 12.0247
R560 VTAIL.n39 VTAIL.n38 12.0247
R561 VTAIL.n51 VTAIL.n8 12.0247
R562 VTAIL.n187 VTAIL.n144 12.0247
R563 VTAIL.n176 VTAIL.n149 12.0247
R564 VTAIL.n121 VTAIL.n78 12.0247
R565 VTAIL.n110 VTAIL.n83 12.0247
R566 VTAIL.n235 VTAIL.n212 11.249
R567 VTAIL.n250 VTAIL.n204 11.249
R568 VTAIL.n37 VTAIL.n14 11.249
R569 VTAIL.n52 VTAIL.n6 11.249
R570 VTAIL.n188 VTAIL.n142 11.249
R571 VTAIL.n175 VTAIL.n152 11.249
R572 VTAIL.n122 VTAIL.n76 11.249
R573 VTAIL.n109 VTAIL.n86 11.249
R574 VTAIL.n232 VTAIL.n231 10.4732
R575 VTAIL.n254 VTAIL.n253 10.4732
R576 VTAIL.n34 VTAIL.n33 10.4732
R577 VTAIL.n56 VTAIL.n55 10.4732
R578 VTAIL.n192 VTAIL.n191 10.4732
R579 VTAIL.n172 VTAIL.n171 10.4732
R580 VTAIL.n126 VTAIL.n125 10.4732
R581 VTAIL.n106 VTAIL.n105 10.4732
R582 VTAIL.n220 VTAIL.n219 10.2747
R583 VTAIL.n22 VTAIL.n21 10.2747
R584 VTAIL.n160 VTAIL.n159 10.2747
R585 VTAIL.n94 VTAIL.n93 10.2747
R586 VTAIL.n228 VTAIL.n214 9.69747
R587 VTAIL.n257 VTAIL.n202 9.69747
R588 VTAIL.n30 VTAIL.n16 9.69747
R589 VTAIL.n59 VTAIL.n4 9.69747
R590 VTAIL.n195 VTAIL.n140 9.69747
R591 VTAIL.n168 VTAIL.n154 9.69747
R592 VTAIL.n129 VTAIL.n74 9.69747
R593 VTAIL.n102 VTAIL.n88 9.69747
R594 VTAIL.n260 VTAIL.n259 9.45567
R595 VTAIL.n62 VTAIL.n61 9.45567
R596 VTAIL.n198 VTAIL.n197 9.45567
R597 VTAIL.n132 VTAIL.n131 9.45567
R598 VTAIL.n259 VTAIL.n258 9.3005
R599 VTAIL.n202 VTAIL.n201 9.3005
R600 VTAIL.n253 VTAIL.n252 9.3005
R601 VTAIL.n251 VTAIL.n250 9.3005
R602 VTAIL.n206 VTAIL.n205 9.3005
R603 VTAIL.n245 VTAIL.n244 9.3005
R604 VTAIL.n218 VTAIL.n217 9.3005
R605 VTAIL.n225 VTAIL.n224 9.3005
R606 VTAIL.n227 VTAIL.n226 9.3005
R607 VTAIL.n214 VTAIL.n213 9.3005
R608 VTAIL.n233 VTAIL.n232 9.3005
R609 VTAIL.n235 VTAIL.n234 9.3005
R610 VTAIL.n236 VTAIL.n209 9.3005
R611 VTAIL.n243 VTAIL.n242 9.3005
R612 VTAIL.n61 VTAIL.n60 9.3005
R613 VTAIL.n4 VTAIL.n3 9.3005
R614 VTAIL.n55 VTAIL.n54 9.3005
R615 VTAIL.n53 VTAIL.n52 9.3005
R616 VTAIL.n8 VTAIL.n7 9.3005
R617 VTAIL.n47 VTAIL.n46 9.3005
R618 VTAIL.n20 VTAIL.n19 9.3005
R619 VTAIL.n27 VTAIL.n26 9.3005
R620 VTAIL.n29 VTAIL.n28 9.3005
R621 VTAIL.n16 VTAIL.n15 9.3005
R622 VTAIL.n35 VTAIL.n34 9.3005
R623 VTAIL.n37 VTAIL.n36 9.3005
R624 VTAIL.n38 VTAIL.n11 9.3005
R625 VTAIL.n45 VTAIL.n44 9.3005
R626 VTAIL.n158 VTAIL.n157 9.3005
R627 VTAIL.n165 VTAIL.n164 9.3005
R628 VTAIL.n167 VTAIL.n166 9.3005
R629 VTAIL.n154 VTAIL.n153 9.3005
R630 VTAIL.n173 VTAIL.n172 9.3005
R631 VTAIL.n175 VTAIL.n174 9.3005
R632 VTAIL.n149 VTAIL.n147 9.3005
R633 VTAIL.n181 VTAIL.n180 9.3005
R634 VTAIL.n197 VTAIL.n196 9.3005
R635 VTAIL.n140 VTAIL.n139 9.3005
R636 VTAIL.n191 VTAIL.n190 9.3005
R637 VTAIL.n189 VTAIL.n188 9.3005
R638 VTAIL.n144 VTAIL.n143 9.3005
R639 VTAIL.n183 VTAIL.n182 9.3005
R640 VTAIL.n92 VTAIL.n91 9.3005
R641 VTAIL.n99 VTAIL.n98 9.3005
R642 VTAIL.n101 VTAIL.n100 9.3005
R643 VTAIL.n88 VTAIL.n87 9.3005
R644 VTAIL.n107 VTAIL.n106 9.3005
R645 VTAIL.n109 VTAIL.n108 9.3005
R646 VTAIL.n83 VTAIL.n81 9.3005
R647 VTAIL.n115 VTAIL.n114 9.3005
R648 VTAIL.n131 VTAIL.n130 9.3005
R649 VTAIL.n74 VTAIL.n73 9.3005
R650 VTAIL.n125 VTAIL.n124 9.3005
R651 VTAIL.n123 VTAIL.n122 9.3005
R652 VTAIL.n78 VTAIL.n77 9.3005
R653 VTAIL.n117 VTAIL.n116 9.3005
R654 VTAIL.n227 VTAIL.n216 8.92171
R655 VTAIL.n258 VTAIL.n200 8.92171
R656 VTAIL.n29 VTAIL.n18 8.92171
R657 VTAIL.n60 VTAIL.n2 8.92171
R658 VTAIL.n196 VTAIL.n138 8.92171
R659 VTAIL.n167 VTAIL.n156 8.92171
R660 VTAIL.n130 VTAIL.n72 8.92171
R661 VTAIL.n101 VTAIL.n90 8.92171
R662 VTAIL.n224 VTAIL.n223 8.14595
R663 VTAIL.n26 VTAIL.n25 8.14595
R664 VTAIL.n164 VTAIL.n163 8.14595
R665 VTAIL.n98 VTAIL.n97 8.14595
R666 VTAIL.n220 VTAIL.n218 7.3702
R667 VTAIL.n22 VTAIL.n20 7.3702
R668 VTAIL.n160 VTAIL.n158 7.3702
R669 VTAIL.n94 VTAIL.n92 7.3702
R670 VTAIL.n223 VTAIL.n218 5.81868
R671 VTAIL.n25 VTAIL.n20 5.81868
R672 VTAIL.n163 VTAIL.n158 5.81868
R673 VTAIL.n97 VTAIL.n92 5.81868
R674 VTAIL.n224 VTAIL.n216 5.04292
R675 VTAIL.n260 VTAIL.n200 5.04292
R676 VTAIL.n26 VTAIL.n18 5.04292
R677 VTAIL.n62 VTAIL.n2 5.04292
R678 VTAIL.n198 VTAIL.n138 5.04292
R679 VTAIL.n164 VTAIL.n156 5.04292
R680 VTAIL.n132 VTAIL.n72 5.04292
R681 VTAIL.n98 VTAIL.n90 5.04292
R682 VTAIL.n228 VTAIL.n227 4.26717
R683 VTAIL.n258 VTAIL.n257 4.26717
R684 VTAIL.n30 VTAIL.n29 4.26717
R685 VTAIL.n60 VTAIL.n59 4.26717
R686 VTAIL.n196 VTAIL.n195 4.26717
R687 VTAIL.n168 VTAIL.n167 4.26717
R688 VTAIL.n130 VTAIL.n129 4.26717
R689 VTAIL.n102 VTAIL.n101 4.26717
R690 VTAIL.n71 VTAIL.n69 3.59533
R691 VTAIL.n133 VTAIL.n71 3.59533
R692 VTAIL.n137 VTAIL.n135 3.59533
R693 VTAIL.n199 VTAIL.n137 3.59533
R694 VTAIL.n67 VTAIL.n65 3.59533
R695 VTAIL.n65 VTAIL.n63 3.59533
R696 VTAIL.n263 VTAIL.n261 3.59533
R697 VTAIL.n231 VTAIL.n214 3.49141
R698 VTAIL.n254 VTAIL.n202 3.49141
R699 VTAIL.n33 VTAIL.n16 3.49141
R700 VTAIL.n56 VTAIL.n4 3.49141
R701 VTAIL.n192 VTAIL.n140 3.49141
R702 VTAIL.n171 VTAIL.n154 3.49141
R703 VTAIL.n126 VTAIL.n74 3.49141
R704 VTAIL.n105 VTAIL.n88 3.49141
R705 VTAIL.n219 VTAIL.n217 2.84303
R706 VTAIL.n21 VTAIL.n19 2.84303
R707 VTAIL.n159 VTAIL.n157 2.84303
R708 VTAIL.n93 VTAIL.n91 2.84303
R709 VTAIL VTAIL.n1 2.75481
R710 VTAIL.n232 VTAIL.n212 2.71565
R711 VTAIL.n253 VTAIL.n204 2.71565
R712 VTAIL.n34 VTAIL.n14 2.71565
R713 VTAIL.n55 VTAIL.n6 2.71565
R714 VTAIL.n191 VTAIL.n142 2.71565
R715 VTAIL.n172 VTAIL.n152 2.71565
R716 VTAIL.n125 VTAIL.n76 2.71565
R717 VTAIL.n106 VTAIL.n86 2.71565
R718 VTAIL.n135 VTAIL.n133 2.26774
R719 VTAIL.n63 VTAIL.n1 2.26774
R720 VTAIL.n237 VTAIL.n235 1.93989
R721 VTAIL.n250 VTAIL.n249 1.93989
R722 VTAIL.n39 VTAIL.n37 1.93989
R723 VTAIL.n52 VTAIL.n51 1.93989
R724 VTAIL.n188 VTAIL.n187 1.93989
R725 VTAIL.n176 VTAIL.n175 1.93989
R726 VTAIL.n122 VTAIL.n121 1.93989
R727 VTAIL.n110 VTAIL.n109 1.93989
R728 VTAIL.n262 VTAIL.t4 1.74962
R729 VTAIL.n262 VTAIL.t6 1.74962
R730 VTAIL.n0 VTAIL.t8 1.74962
R731 VTAIL.n0 VTAIL.t2 1.74962
R732 VTAIL.n64 VTAIL.t11 1.74962
R733 VTAIL.n64 VTAIL.t13 1.74962
R734 VTAIL.n66 VTAIL.t16 1.74962
R735 VTAIL.n66 VTAIL.t9 1.74962
R736 VTAIL.n136 VTAIL.t14 1.74962
R737 VTAIL.n136 VTAIL.t10 1.74962
R738 VTAIL.n134 VTAIL.t12 1.74962
R739 VTAIL.n134 VTAIL.t18 1.74962
R740 VTAIL.n70 VTAIL.t0 1.74962
R741 VTAIL.n70 VTAIL.t19 1.74962
R742 VTAIL.n68 VTAIL.t1 1.74962
R743 VTAIL.n68 VTAIL.t7 1.74962
R744 VTAIL.n236 VTAIL.n210 1.16414
R745 VTAIL.n246 VTAIL.n206 1.16414
R746 VTAIL.n38 VTAIL.n12 1.16414
R747 VTAIL.n48 VTAIL.n8 1.16414
R748 VTAIL.n184 VTAIL.n144 1.16414
R749 VTAIL.n179 VTAIL.n149 1.16414
R750 VTAIL.n118 VTAIL.n78 1.16414
R751 VTAIL.n113 VTAIL.n83 1.16414
R752 VTAIL VTAIL.n263 0.841017
R753 VTAIL.n242 VTAIL.n241 0.388379
R754 VTAIL.n245 VTAIL.n208 0.388379
R755 VTAIL.n44 VTAIL.n43 0.388379
R756 VTAIL.n47 VTAIL.n10 0.388379
R757 VTAIL.n183 VTAIL.n146 0.388379
R758 VTAIL.n180 VTAIL.n148 0.388379
R759 VTAIL.n117 VTAIL.n80 0.388379
R760 VTAIL.n114 VTAIL.n82 0.388379
R761 VTAIL.n225 VTAIL.n217 0.155672
R762 VTAIL.n226 VTAIL.n225 0.155672
R763 VTAIL.n226 VTAIL.n213 0.155672
R764 VTAIL.n233 VTAIL.n213 0.155672
R765 VTAIL.n234 VTAIL.n233 0.155672
R766 VTAIL.n234 VTAIL.n209 0.155672
R767 VTAIL.n243 VTAIL.n209 0.155672
R768 VTAIL.n244 VTAIL.n243 0.155672
R769 VTAIL.n244 VTAIL.n205 0.155672
R770 VTAIL.n251 VTAIL.n205 0.155672
R771 VTAIL.n252 VTAIL.n251 0.155672
R772 VTAIL.n252 VTAIL.n201 0.155672
R773 VTAIL.n259 VTAIL.n201 0.155672
R774 VTAIL.n27 VTAIL.n19 0.155672
R775 VTAIL.n28 VTAIL.n27 0.155672
R776 VTAIL.n28 VTAIL.n15 0.155672
R777 VTAIL.n35 VTAIL.n15 0.155672
R778 VTAIL.n36 VTAIL.n35 0.155672
R779 VTAIL.n36 VTAIL.n11 0.155672
R780 VTAIL.n45 VTAIL.n11 0.155672
R781 VTAIL.n46 VTAIL.n45 0.155672
R782 VTAIL.n46 VTAIL.n7 0.155672
R783 VTAIL.n53 VTAIL.n7 0.155672
R784 VTAIL.n54 VTAIL.n53 0.155672
R785 VTAIL.n54 VTAIL.n3 0.155672
R786 VTAIL.n61 VTAIL.n3 0.155672
R787 VTAIL.n197 VTAIL.n139 0.155672
R788 VTAIL.n190 VTAIL.n139 0.155672
R789 VTAIL.n190 VTAIL.n189 0.155672
R790 VTAIL.n189 VTAIL.n143 0.155672
R791 VTAIL.n182 VTAIL.n143 0.155672
R792 VTAIL.n182 VTAIL.n181 0.155672
R793 VTAIL.n181 VTAIL.n147 0.155672
R794 VTAIL.n174 VTAIL.n147 0.155672
R795 VTAIL.n174 VTAIL.n173 0.155672
R796 VTAIL.n173 VTAIL.n153 0.155672
R797 VTAIL.n166 VTAIL.n153 0.155672
R798 VTAIL.n166 VTAIL.n165 0.155672
R799 VTAIL.n165 VTAIL.n157 0.155672
R800 VTAIL.n131 VTAIL.n73 0.155672
R801 VTAIL.n124 VTAIL.n73 0.155672
R802 VTAIL.n124 VTAIL.n123 0.155672
R803 VTAIL.n123 VTAIL.n77 0.155672
R804 VTAIL.n116 VTAIL.n77 0.155672
R805 VTAIL.n116 VTAIL.n115 0.155672
R806 VTAIL.n115 VTAIL.n81 0.155672
R807 VTAIL.n108 VTAIL.n81 0.155672
R808 VTAIL.n108 VTAIL.n107 0.155672
R809 VTAIL.n107 VTAIL.n87 0.155672
R810 VTAIL.n100 VTAIL.n87 0.155672
R811 VTAIL.n100 VTAIL.n99 0.155672
R812 VTAIL.n99 VTAIL.n91 0.155672
R813 B.n1110 B.n1109 585
R814 B.n1111 B.n1110 585
R815 B.n373 B.n192 585
R816 B.n372 B.n371 585
R817 B.n370 B.n369 585
R818 B.n368 B.n367 585
R819 B.n366 B.n365 585
R820 B.n364 B.n363 585
R821 B.n362 B.n361 585
R822 B.n360 B.n359 585
R823 B.n358 B.n357 585
R824 B.n356 B.n355 585
R825 B.n354 B.n353 585
R826 B.n352 B.n351 585
R827 B.n350 B.n349 585
R828 B.n348 B.n347 585
R829 B.n346 B.n345 585
R830 B.n344 B.n343 585
R831 B.n342 B.n341 585
R832 B.n340 B.n339 585
R833 B.n338 B.n337 585
R834 B.n336 B.n335 585
R835 B.n334 B.n333 585
R836 B.n332 B.n331 585
R837 B.n330 B.n329 585
R838 B.n328 B.n327 585
R839 B.n326 B.n325 585
R840 B.n324 B.n323 585
R841 B.n322 B.n321 585
R842 B.n320 B.n319 585
R843 B.n318 B.n317 585
R844 B.n316 B.n315 585
R845 B.n314 B.n313 585
R846 B.n312 B.n311 585
R847 B.n310 B.n309 585
R848 B.n308 B.n307 585
R849 B.n306 B.n305 585
R850 B.n304 B.n303 585
R851 B.n302 B.n301 585
R852 B.n300 B.n299 585
R853 B.n298 B.n297 585
R854 B.n295 B.n294 585
R855 B.n293 B.n292 585
R856 B.n291 B.n290 585
R857 B.n289 B.n288 585
R858 B.n287 B.n286 585
R859 B.n285 B.n284 585
R860 B.n283 B.n282 585
R861 B.n281 B.n280 585
R862 B.n279 B.n278 585
R863 B.n277 B.n276 585
R864 B.n275 B.n274 585
R865 B.n273 B.n272 585
R866 B.n271 B.n270 585
R867 B.n269 B.n268 585
R868 B.n267 B.n266 585
R869 B.n265 B.n264 585
R870 B.n263 B.n262 585
R871 B.n261 B.n260 585
R872 B.n259 B.n258 585
R873 B.n257 B.n256 585
R874 B.n255 B.n254 585
R875 B.n253 B.n252 585
R876 B.n251 B.n250 585
R877 B.n249 B.n248 585
R878 B.n247 B.n246 585
R879 B.n245 B.n244 585
R880 B.n243 B.n242 585
R881 B.n241 B.n240 585
R882 B.n239 B.n238 585
R883 B.n237 B.n236 585
R884 B.n235 B.n234 585
R885 B.n233 B.n232 585
R886 B.n231 B.n230 585
R887 B.n229 B.n228 585
R888 B.n227 B.n226 585
R889 B.n225 B.n224 585
R890 B.n223 B.n222 585
R891 B.n221 B.n220 585
R892 B.n219 B.n218 585
R893 B.n217 B.n216 585
R894 B.n215 B.n214 585
R895 B.n213 B.n212 585
R896 B.n211 B.n210 585
R897 B.n209 B.n208 585
R898 B.n207 B.n206 585
R899 B.n205 B.n204 585
R900 B.n203 B.n202 585
R901 B.n201 B.n200 585
R902 B.n199 B.n198 585
R903 B.n1108 B.n147 585
R904 B.n1112 B.n147 585
R905 B.n1107 B.n146 585
R906 B.n1113 B.n146 585
R907 B.n1106 B.n1105 585
R908 B.n1105 B.n142 585
R909 B.n1104 B.n141 585
R910 B.n1119 B.n141 585
R911 B.n1103 B.n140 585
R912 B.n1120 B.n140 585
R913 B.n1102 B.n139 585
R914 B.n1121 B.n139 585
R915 B.n1101 B.n1100 585
R916 B.n1100 B.n135 585
R917 B.n1099 B.n134 585
R918 B.n1127 B.n134 585
R919 B.n1098 B.n133 585
R920 B.n1128 B.n133 585
R921 B.n1097 B.n132 585
R922 B.n1129 B.n132 585
R923 B.n1096 B.n1095 585
R924 B.n1095 B.n128 585
R925 B.n1094 B.n127 585
R926 B.n1135 B.n127 585
R927 B.n1093 B.n126 585
R928 B.n1136 B.n126 585
R929 B.n1092 B.n125 585
R930 B.n1137 B.n125 585
R931 B.n1091 B.n1090 585
R932 B.n1090 B.n121 585
R933 B.n1089 B.n120 585
R934 B.n1143 B.n120 585
R935 B.n1088 B.n119 585
R936 B.n1144 B.n119 585
R937 B.n1087 B.n118 585
R938 B.n1145 B.n118 585
R939 B.n1086 B.n1085 585
R940 B.n1085 B.n114 585
R941 B.n1084 B.n113 585
R942 B.n1151 B.n113 585
R943 B.n1083 B.n112 585
R944 B.n1152 B.n112 585
R945 B.n1082 B.n111 585
R946 B.n1153 B.n111 585
R947 B.n1081 B.n1080 585
R948 B.n1080 B.n107 585
R949 B.n1079 B.n106 585
R950 B.n1159 B.n106 585
R951 B.n1078 B.n105 585
R952 B.n1160 B.n105 585
R953 B.n1077 B.n104 585
R954 B.n1161 B.n104 585
R955 B.n1076 B.n1075 585
R956 B.n1075 B.n100 585
R957 B.n1074 B.n99 585
R958 B.n1167 B.n99 585
R959 B.n1073 B.n98 585
R960 B.n1168 B.n98 585
R961 B.n1072 B.n97 585
R962 B.n1169 B.n97 585
R963 B.n1071 B.n1070 585
R964 B.n1070 B.n93 585
R965 B.n1069 B.n92 585
R966 B.n1175 B.n92 585
R967 B.n1068 B.n91 585
R968 B.n1176 B.n91 585
R969 B.n1067 B.n90 585
R970 B.n1177 B.n90 585
R971 B.n1066 B.n1065 585
R972 B.n1065 B.n86 585
R973 B.n1064 B.n85 585
R974 B.n1183 B.n85 585
R975 B.n1063 B.n84 585
R976 B.n1184 B.n84 585
R977 B.n1062 B.n83 585
R978 B.n1185 B.n83 585
R979 B.n1061 B.n1060 585
R980 B.n1060 B.n79 585
R981 B.n1059 B.n78 585
R982 B.n1191 B.n78 585
R983 B.n1058 B.n77 585
R984 B.n1192 B.n77 585
R985 B.n1057 B.n76 585
R986 B.n1193 B.n76 585
R987 B.n1056 B.n1055 585
R988 B.n1055 B.n72 585
R989 B.n1054 B.n71 585
R990 B.n1199 B.n71 585
R991 B.n1053 B.n70 585
R992 B.n1200 B.n70 585
R993 B.n1052 B.n69 585
R994 B.n1201 B.n69 585
R995 B.n1051 B.n1050 585
R996 B.n1050 B.n65 585
R997 B.n1049 B.n64 585
R998 B.n1207 B.n64 585
R999 B.n1048 B.n63 585
R1000 B.n1208 B.n63 585
R1001 B.n1047 B.n62 585
R1002 B.n1209 B.n62 585
R1003 B.n1046 B.n1045 585
R1004 B.n1045 B.n58 585
R1005 B.n1044 B.n57 585
R1006 B.n1215 B.n57 585
R1007 B.n1043 B.n56 585
R1008 B.n1216 B.n56 585
R1009 B.n1042 B.n55 585
R1010 B.n1217 B.n55 585
R1011 B.n1041 B.n1040 585
R1012 B.n1040 B.n51 585
R1013 B.n1039 B.n50 585
R1014 B.n1223 B.n50 585
R1015 B.n1038 B.n49 585
R1016 B.n1224 B.n49 585
R1017 B.n1037 B.n48 585
R1018 B.n1225 B.n48 585
R1019 B.n1036 B.n1035 585
R1020 B.n1035 B.n44 585
R1021 B.n1034 B.n43 585
R1022 B.n1231 B.n43 585
R1023 B.n1033 B.n42 585
R1024 B.n1232 B.n42 585
R1025 B.n1032 B.n41 585
R1026 B.n1233 B.n41 585
R1027 B.n1031 B.n1030 585
R1028 B.n1030 B.n37 585
R1029 B.n1029 B.n36 585
R1030 B.n1239 B.n36 585
R1031 B.n1028 B.n35 585
R1032 B.n1240 B.n35 585
R1033 B.n1027 B.n34 585
R1034 B.n1241 B.n34 585
R1035 B.n1026 B.n1025 585
R1036 B.n1025 B.n30 585
R1037 B.n1024 B.n29 585
R1038 B.n1247 B.n29 585
R1039 B.n1023 B.n28 585
R1040 B.n1248 B.n28 585
R1041 B.n1022 B.n27 585
R1042 B.n1249 B.n27 585
R1043 B.n1021 B.n1020 585
R1044 B.n1020 B.n23 585
R1045 B.n1019 B.n22 585
R1046 B.n1255 B.n22 585
R1047 B.n1018 B.n21 585
R1048 B.n1256 B.n21 585
R1049 B.n1017 B.n20 585
R1050 B.n1257 B.n20 585
R1051 B.n1016 B.n1015 585
R1052 B.n1015 B.n16 585
R1053 B.n1014 B.n15 585
R1054 B.n1263 B.n15 585
R1055 B.n1013 B.n14 585
R1056 B.n1264 B.n14 585
R1057 B.n1012 B.n13 585
R1058 B.n1265 B.n13 585
R1059 B.n1011 B.n1010 585
R1060 B.n1010 B.n12 585
R1061 B.n1009 B.n1008 585
R1062 B.n1009 B.n8 585
R1063 B.n1007 B.n7 585
R1064 B.n1272 B.n7 585
R1065 B.n1006 B.n6 585
R1066 B.n1273 B.n6 585
R1067 B.n1005 B.n5 585
R1068 B.n1274 B.n5 585
R1069 B.n1004 B.n1003 585
R1070 B.n1003 B.n4 585
R1071 B.n1002 B.n374 585
R1072 B.n1002 B.n1001 585
R1073 B.n992 B.n375 585
R1074 B.n376 B.n375 585
R1075 B.n994 B.n993 585
R1076 B.n995 B.n994 585
R1077 B.n991 B.n381 585
R1078 B.n381 B.n380 585
R1079 B.n990 B.n989 585
R1080 B.n989 B.n988 585
R1081 B.n383 B.n382 585
R1082 B.n384 B.n383 585
R1083 B.n981 B.n980 585
R1084 B.n982 B.n981 585
R1085 B.n979 B.n389 585
R1086 B.n389 B.n388 585
R1087 B.n978 B.n977 585
R1088 B.n977 B.n976 585
R1089 B.n391 B.n390 585
R1090 B.n392 B.n391 585
R1091 B.n969 B.n968 585
R1092 B.n970 B.n969 585
R1093 B.n967 B.n397 585
R1094 B.n397 B.n396 585
R1095 B.n966 B.n965 585
R1096 B.n965 B.n964 585
R1097 B.n399 B.n398 585
R1098 B.n400 B.n399 585
R1099 B.n957 B.n956 585
R1100 B.n958 B.n957 585
R1101 B.n955 B.n405 585
R1102 B.n405 B.n404 585
R1103 B.n954 B.n953 585
R1104 B.n953 B.n952 585
R1105 B.n407 B.n406 585
R1106 B.n408 B.n407 585
R1107 B.n945 B.n944 585
R1108 B.n946 B.n945 585
R1109 B.n943 B.n413 585
R1110 B.n413 B.n412 585
R1111 B.n942 B.n941 585
R1112 B.n941 B.n940 585
R1113 B.n415 B.n414 585
R1114 B.n416 B.n415 585
R1115 B.n933 B.n932 585
R1116 B.n934 B.n933 585
R1117 B.n931 B.n421 585
R1118 B.n421 B.n420 585
R1119 B.n930 B.n929 585
R1120 B.n929 B.n928 585
R1121 B.n423 B.n422 585
R1122 B.n424 B.n423 585
R1123 B.n921 B.n920 585
R1124 B.n922 B.n921 585
R1125 B.n919 B.n429 585
R1126 B.n429 B.n428 585
R1127 B.n918 B.n917 585
R1128 B.n917 B.n916 585
R1129 B.n431 B.n430 585
R1130 B.n432 B.n431 585
R1131 B.n909 B.n908 585
R1132 B.n910 B.n909 585
R1133 B.n907 B.n437 585
R1134 B.n437 B.n436 585
R1135 B.n906 B.n905 585
R1136 B.n905 B.n904 585
R1137 B.n439 B.n438 585
R1138 B.n440 B.n439 585
R1139 B.n897 B.n896 585
R1140 B.n898 B.n897 585
R1141 B.n895 B.n445 585
R1142 B.n445 B.n444 585
R1143 B.n894 B.n893 585
R1144 B.n893 B.n892 585
R1145 B.n447 B.n446 585
R1146 B.n448 B.n447 585
R1147 B.n885 B.n884 585
R1148 B.n886 B.n885 585
R1149 B.n883 B.n453 585
R1150 B.n453 B.n452 585
R1151 B.n882 B.n881 585
R1152 B.n881 B.n880 585
R1153 B.n455 B.n454 585
R1154 B.n456 B.n455 585
R1155 B.n873 B.n872 585
R1156 B.n874 B.n873 585
R1157 B.n871 B.n460 585
R1158 B.n464 B.n460 585
R1159 B.n870 B.n869 585
R1160 B.n869 B.n868 585
R1161 B.n462 B.n461 585
R1162 B.n463 B.n462 585
R1163 B.n861 B.n860 585
R1164 B.n862 B.n861 585
R1165 B.n859 B.n469 585
R1166 B.n469 B.n468 585
R1167 B.n858 B.n857 585
R1168 B.n857 B.n856 585
R1169 B.n471 B.n470 585
R1170 B.n472 B.n471 585
R1171 B.n849 B.n848 585
R1172 B.n850 B.n849 585
R1173 B.n847 B.n477 585
R1174 B.n477 B.n476 585
R1175 B.n846 B.n845 585
R1176 B.n845 B.n844 585
R1177 B.n479 B.n478 585
R1178 B.n480 B.n479 585
R1179 B.n837 B.n836 585
R1180 B.n838 B.n837 585
R1181 B.n835 B.n484 585
R1182 B.n488 B.n484 585
R1183 B.n834 B.n833 585
R1184 B.n833 B.n832 585
R1185 B.n486 B.n485 585
R1186 B.n487 B.n486 585
R1187 B.n825 B.n824 585
R1188 B.n826 B.n825 585
R1189 B.n823 B.n493 585
R1190 B.n493 B.n492 585
R1191 B.n822 B.n821 585
R1192 B.n821 B.n820 585
R1193 B.n495 B.n494 585
R1194 B.n496 B.n495 585
R1195 B.n813 B.n812 585
R1196 B.n814 B.n813 585
R1197 B.n811 B.n501 585
R1198 B.n501 B.n500 585
R1199 B.n810 B.n809 585
R1200 B.n809 B.n808 585
R1201 B.n503 B.n502 585
R1202 B.n504 B.n503 585
R1203 B.n801 B.n800 585
R1204 B.n802 B.n801 585
R1205 B.n799 B.n509 585
R1206 B.n509 B.n508 585
R1207 B.n798 B.n797 585
R1208 B.n797 B.n796 585
R1209 B.n511 B.n510 585
R1210 B.n512 B.n511 585
R1211 B.n789 B.n788 585
R1212 B.n790 B.n789 585
R1213 B.n787 B.n517 585
R1214 B.n517 B.n516 585
R1215 B.n786 B.n785 585
R1216 B.n785 B.n784 585
R1217 B.n519 B.n518 585
R1218 B.n520 B.n519 585
R1219 B.n777 B.n776 585
R1220 B.n778 B.n777 585
R1221 B.n775 B.n525 585
R1222 B.n525 B.n524 585
R1223 B.n774 B.n773 585
R1224 B.n773 B.n772 585
R1225 B.n527 B.n526 585
R1226 B.n528 B.n527 585
R1227 B.n765 B.n764 585
R1228 B.n766 B.n765 585
R1229 B.n763 B.n533 585
R1230 B.n533 B.n532 585
R1231 B.n757 B.n756 585
R1232 B.n755 B.n579 585
R1233 B.n754 B.n578 585
R1234 B.n759 B.n578 585
R1235 B.n753 B.n752 585
R1236 B.n751 B.n750 585
R1237 B.n749 B.n748 585
R1238 B.n747 B.n746 585
R1239 B.n745 B.n744 585
R1240 B.n743 B.n742 585
R1241 B.n741 B.n740 585
R1242 B.n739 B.n738 585
R1243 B.n737 B.n736 585
R1244 B.n735 B.n734 585
R1245 B.n733 B.n732 585
R1246 B.n731 B.n730 585
R1247 B.n729 B.n728 585
R1248 B.n727 B.n726 585
R1249 B.n725 B.n724 585
R1250 B.n723 B.n722 585
R1251 B.n721 B.n720 585
R1252 B.n719 B.n718 585
R1253 B.n717 B.n716 585
R1254 B.n715 B.n714 585
R1255 B.n713 B.n712 585
R1256 B.n711 B.n710 585
R1257 B.n709 B.n708 585
R1258 B.n707 B.n706 585
R1259 B.n705 B.n704 585
R1260 B.n703 B.n702 585
R1261 B.n701 B.n700 585
R1262 B.n699 B.n698 585
R1263 B.n697 B.n696 585
R1264 B.n695 B.n694 585
R1265 B.n693 B.n692 585
R1266 B.n691 B.n690 585
R1267 B.n689 B.n688 585
R1268 B.n687 B.n686 585
R1269 B.n685 B.n684 585
R1270 B.n683 B.n682 585
R1271 B.n681 B.n680 585
R1272 B.n678 B.n677 585
R1273 B.n676 B.n675 585
R1274 B.n674 B.n673 585
R1275 B.n672 B.n671 585
R1276 B.n670 B.n669 585
R1277 B.n668 B.n667 585
R1278 B.n666 B.n665 585
R1279 B.n664 B.n663 585
R1280 B.n662 B.n661 585
R1281 B.n660 B.n659 585
R1282 B.n658 B.n657 585
R1283 B.n656 B.n655 585
R1284 B.n654 B.n653 585
R1285 B.n652 B.n651 585
R1286 B.n650 B.n649 585
R1287 B.n648 B.n647 585
R1288 B.n646 B.n645 585
R1289 B.n644 B.n643 585
R1290 B.n642 B.n641 585
R1291 B.n640 B.n639 585
R1292 B.n638 B.n637 585
R1293 B.n636 B.n635 585
R1294 B.n634 B.n633 585
R1295 B.n632 B.n631 585
R1296 B.n630 B.n629 585
R1297 B.n628 B.n627 585
R1298 B.n626 B.n625 585
R1299 B.n624 B.n623 585
R1300 B.n622 B.n621 585
R1301 B.n620 B.n619 585
R1302 B.n618 B.n617 585
R1303 B.n616 B.n615 585
R1304 B.n614 B.n613 585
R1305 B.n612 B.n611 585
R1306 B.n610 B.n609 585
R1307 B.n608 B.n607 585
R1308 B.n606 B.n605 585
R1309 B.n604 B.n603 585
R1310 B.n602 B.n601 585
R1311 B.n600 B.n599 585
R1312 B.n598 B.n597 585
R1313 B.n596 B.n595 585
R1314 B.n594 B.n593 585
R1315 B.n592 B.n591 585
R1316 B.n590 B.n589 585
R1317 B.n588 B.n587 585
R1318 B.n586 B.n585 585
R1319 B.n535 B.n534 585
R1320 B.n762 B.n761 585
R1321 B.n531 B.n530 585
R1322 B.n532 B.n531 585
R1323 B.n768 B.n767 585
R1324 B.n767 B.n766 585
R1325 B.n769 B.n529 585
R1326 B.n529 B.n528 585
R1327 B.n771 B.n770 585
R1328 B.n772 B.n771 585
R1329 B.n523 B.n522 585
R1330 B.n524 B.n523 585
R1331 B.n780 B.n779 585
R1332 B.n779 B.n778 585
R1333 B.n781 B.n521 585
R1334 B.n521 B.n520 585
R1335 B.n783 B.n782 585
R1336 B.n784 B.n783 585
R1337 B.n515 B.n514 585
R1338 B.n516 B.n515 585
R1339 B.n792 B.n791 585
R1340 B.n791 B.n790 585
R1341 B.n793 B.n513 585
R1342 B.n513 B.n512 585
R1343 B.n795 B.n794 585
R1344 B.n796 B.n795 585
R1345 B.n507 B.n506 585
R1346 B.n508 B.n507 585
R1347 B.n804 B.n803 585
R1348 B.n803 B.n802 585
R1349 B.n805 B.n505 585
R1350 B.n505 B.n504 585
R1351 B.n807 B.n806 585
R1352 B.n808 B.n807 585
R1353 B.n499 B.n498 585
R1354 B.n500 B.n499 585
R1355 B.n816 B.n815 585
R1356 B.n815 B.n814 585
R1357 B.n817 B.n497 585
R1358 B.n497 B.n496 585
R1359 B.n819 B.n818 585
R1360 B.n820 B.n819 585
R1361 B.n491 B.n490 585
R1362 B.n492 B.n491 585
R1363 B.n828 B.n827 585
R1364 B.n827 B.n826 585
R1365 B.n829 B.n489 585
R1366 B.n489 B.n487 585
R1367 B.n831 B.n830 585
R1368 B.n832 B.n831 585
R1369 B.n483 B.n482 585
R1370 B.n488 B.n483 585
R1371 B.n840 B.n839 585
R1372 B.n839 B.n838 585
R1373 B.n841 B.n481 585
R1374 B.n481 B.n480 585
R1375 B.n843 B.n842 585
R1376 B.n844 B.n843 585
R1377 B.n475 B.n474 585
R1378 B.n476 B.n475 585
R1379 B.n852 B.n851 585
R1380 B.n851 B.n850 585
R1381 B.n853 B.n473 585
R1382 B.n473 B.n472 585
R1383 B.n855 B.n854 585
R1384 B.n856 B.n855 585
R1385 B.n467 B.n466 585
R1386 B.n468 B.n467 585
R1387 B.n864 B.n863 585
R1388 B.n863 B.n862 585
R1389 B.n865 B.n465 585
R1390 B.n465 B.n463 585
R1391 B.n867 B.n866 585
R1392 B.n868 B.n867 585
R1393 B.n459 B.n458 585
R1394 B.n464 B.n459 585
R1395 B.n876 B.n875 585
R1396 B.n875 B.n874 585
R1397 B.n877 B.n457 585
R1398 B.n457 B.n456 585
R1399 B.n879 B.n878 585
R1400 B.n880 B.n879 585
R1401 B.n451 B.n450 585
R1402 B.n452 B.n451 585
R1403 B.n888 B.n887 585
R1404 B.n887 B.n886 585
R1405 B.n889 B.n449 585
R1406 B.n449 B.n448 585
R1407 B.n891 B.n890 585
R1408 B.n892 B.n891 585
R1409 B.n443 B.n442 585
R1410 B.n444 B.n443 585
R1411 B.n900 B.n899 585
R1412 B.n899 B.n898 585
R1413 B.n901 B.n441 585
R1414 B.n441 B.n440 585
R1415 B.n903 B.n902 585
R1416 B.n904 B.n903 585
R1417 B.n435 B.n434 585
R1418 B.n436 B.n435 585
R1419 B.n912 B.n911 585
R1420 B.n911 B.n910 585
R1421 B.n913 B.n433 585
R1422 B.n433 B.n432 585
R1423 B.n915 B.n914 585
R1424 B.n916 B.n915 585
R1425 B.n427 B.n426 585
R1426 B.n428 B.n427 585
R1427 B.n924 B.n923 585
R1428 B.n923 B.n922 585
R1429 B.n925 B.n425 585
R1430 B.n425 B.n424 585
R1431 B.n927 B.n926 585
R1432 B.n928 B.n927 585
R1433 B.n419 B.n418 585
R1434 B.n420 B.n419 585
R1435 B.n936 B.n935 585
R1436 B.n935 B.n934 585
R1437 B.n937 B.n417 585
R1438 B.n417 B.n416 585
R1439 B.n939 B.n938 585
R1440 B.n940 B.n939 585
R1441 B.n411 B.n410 585
R1442 B.n412 B.n411 585
R1443 B.n948 B.n947 585
R1444 B.n947 B.n946 585
R1445 B.n949 B.n409 585
R1446 B.n409 B.n408 585
R1447 B.n951 B.n950 585
R1448 B.n952 B.n951 585
R1449 B.n403 B.n402 585
R1450 B.n404 B.n403 585
R1451 B.n960 B.n959 585
R1452 B.n959 B.n958 585
R1453 B.n961 B.n401 585
R1454 B.n401 B.n400 585
R1455 B.n963 B.n962 585
R1456 B.n964 B.n963 585
R1457 B.n395 B.n394 585
R1458 B.n396 B.n395 585
R1459 B.n972 B.n971 585
R1460 B.n971 B.n970 585
R1461 B.n973 B.n393 585
R1462 B.n393 B.n392 585
R1463 B.n975 B.n974 585
R1464 B.n976 B.n975 585
R1465 B.n387 B.n386 585
R1466 B.n388 B.n387 585
R1467 B.n984 B.n983 585
R1468 B.n983 B.n982 585
R1469 B.n985 B.n385 585
R1470 B.n385 B.n384 585
R1471 B.n987 B.n986 585
R1472 B.n988 B.n987 585
R1473 B.n379 B.n378 585
R1474 B.n380 B.n379 585
R1475 B.n997 B.n996 585
R1476 B.n996 B.n995 585
R1477 B.n998 B.n377 585
R1478 B.n377 B.n376 585
R1479 B.n1000 B.n999 585
R1480 B.n1001 B.n1000 585
R1481 B.n3 B.n0 585
R1482 B.n4 B.n3 585
R1483 B.n1271 B.n1 585
R1484 B.n1272 B.n1271 585
R1485 B.n1270 B.n1269 585
R1486 B.n1270 B.n8 585
R1487 B.n1268 B.n9 585
R1488 B.n12 B.n9 585
R1489 B.n1267 B.n1266 585
R1490 B.n1266 B.n1265 585
R1491 B.n11 B.n10 585
R1492 B.n1264 B.n11 585
R1493 B.n1262 B.n1261 585
R1494 B.n1263 B.n1262 585
R1495 B.n1260 B.n17 585
R1496 B.n17 B.n16 585
R1497 B.n1259 B.n1258 585
R1498 B.n1258 B.n1257 585
R1499 B.n19 B.n18 585
R1500 B.n1256 B.n19 585
R1501 B.n1254 B.n1253 585
R1502 B.n1255 B.n1254 585
R1503 B.n1252 B.n24 585
R1504 B.n24 B.n23 585
R1505 B.n1251 B.n1250 585
R1506 B.n1250 B.n1249 585
R1507 B.n26 B.n25 585
R1508 B.n1248 B.n26 585
R1509 B.n1246 B.n1245 585
R1510 B.n1247 B.n1246 585
R1511 B.n1244 B.n31 585
R1512 B.n31 B.n30 585
R1513 B.n1243 B.n1242 585
R1514 B.n1242 B.n1241 585
R1515 B.n33 B.n32 585
R1516 B.n1240 B.n33 585
R1517 B.n1238 B.n1237 585
R1518 B.n1239 B.n1238 585
R1519 B.n1236 B.n38 585
R1520 B.n38 B.n37 585
R1521 B.n1235 B.n1234 585
R1522 B.n1234 B.n1233 585
R1523 B.n40 B.n39 585
R1524 B.n1232 B.n40 585
R1525 B.n1230 B.n1229 585
R1526 B.n1231 B.n1230 585
R1527 B.n1228 B.n45 585
R1528 B.n45 B.n44 585
R1529 B.n1227 B.n1226 585
R1530 B.n1226 B.n1225 585
R1531 B.n47 B.n46 585
R1532 B.n1224 B.n47 585
R1533 B.n1222 B.n1221 585
R1534 B.n1223 B.n1222 585
R1535 B.n1220 B.n52 585
R1536 B.n52 B.n51 585
R1537 B.n1219 B.n1218 585
R1538 B.n1218 B.n1217 585
R1539 B.n54 B.n53 585
R1540 B.n1216 B.n54 585
R1541 B.n1214 B.n1213 585
R1542 B.n1215 B.n1214 585
R1543 B.n1212 B.n59 585
R1544 B.n59 B.n58 585
R1545 B.n1211 B.n1210 585
R1546 B.n1210 B.n1209 585
R1547 B.n61 B.n60 585
R1548 B.n1208 B.n61 585
R1549 B.n1206 B.n1205 585
R1550 B.n1207 B.n1206 585
R1551 B.n1204 B.n66 585
R1552 B.n66 B.n65 585
R1553 B.n1203 B.n1202 585
R1554 B.n1202 B.n1201 585
R1555 B.n68 B.n67 585
R1556 B.n1200 B.n68 585
R1557 B.n1198 B.n1197 585
R1558 B.n1199 B.n1198 585
R1559 B.n1196 B.n73 585
R1560 B.n73 B.n72 585
R1561 B.n1195 B.n1194 585
R1562 B.n1194 B.n1193 585
R1563 B.n75 B.n74 585
R1564 B.n1192 B.n75 585
R1565 B.n1190 B.n1189 585
R1566 B.n1191 B.n1190 585
R1567 B.n1188 B.n80 585
R1568 B.n80 B.n79 585
R1569 B.n1187 B.n1186 585
R1570 B.n1186 B.n1185 585
R1571 B.n82 B.n81 585
R1572 B.n1184 B.n82 585
R1573 B.n1182 B.n1181 585
R1574 B.n1183 B.n1182 585
R1575 B.n1180 B.n87 585
R1576 B.n87 B.n86 585
R1577 B.n1179 B.n1178 585
R1578 B.n1178 B.n1177 585
R1579 B.n89 B.n88 585
R1580 B.n1176 B.n89 585
R1581 B.n1174 B.n1173 585
R1582 B.n1175 B.n1174 585
R1583 B.n1172 B.n94 585
R1584 B.n94 B.n93 585
R1585 B.n1171 B.n1170 585
R1586 B.n1170 B.n1169 585
R1587 B.n96 B.n95 585
R1588 B.n1168 B.n96 585
R1589 B.n1166 B.n1165 585
R1590 B.n1167 B.n1166 585
R1591 B.n1164 B.n101 585
R1592 B.n101 B.n100 585
R1593 B.n1163 B.n1162 585
R1594 B.n1162 B.n1161 585
R1595 B.n103 B.n102 585
R1596 B.n1160 B.n103 585
R1597 B.n1158 B.n1157 585
R1598 B.n1159 B.n1158 585
R1599 B.n1156 B.n108 585
R1600 B.n108 B.n107 585
R1601 B.n1155 B.n1154 585
R1602 B.n1154 B.n1153 585
R1603 B.n110 B.n109 585
R1604 B.n1152 B.n110 585
R1605 B.n1150 B.n1149 585
R1606 B.n1151 B.n1150 585
R1607 B.n1148 B.n115 585
R1608 B.n115 B.n114 585
R1609 B.n1147 B.n1146 585
R1610 B.n1146 B.n1145 585
R1611 B.n117 B.n116 585
R1612 B.n1144 B.n117 585
R1613 B.n1142 B.n1141 585
R1614 B.n1143 B.n1142 585
R1615 B.n1140 B.n122 585
R1616 B.n122 B.n121 585
R1617 B.n1139 B.n1138 585
R1618 B.n1138 B.n1137 585
R1619 B.n124 B.n123 585
R1620 B.n1136 B.n124 585
R1621 B.n1134 B.n1133 585
R1622 B.n1135 B.n1134 585
R1623 B.n1132 B.n129 585
R1624 B.n129 B.n128 585
R1625 B.n1131 B.n1130 585
R1626 B.n1130 B.n1129 585
R1627 B.n131 B.n130 585
R1628 B.n1128 B.n131 585
R1629 B.n1126 B.n1125 585
R1630 B.n1127 B.n1126 585
R1631 B.n1124 B.n136 585
R1632 B.n136 B.n135 585
R1633 B.n1123 B.n1122 585
R1634 B.n1122 B.n1121 585
R1635 B.n138 B.n137 585
R1636 B.n1120 B.n138 585
R1637 B.n1118 B.n1117 585
R1638 B.n1119 B.n1118 585
R1639 B.n1116 B.n143 585
R1640 B.n143 B.n142 585
R1641 B.n1115 B.n1114 585
R1642 B.n1114 B.n1113 585
R1643 B.n145 B.n144 585
R1644 B.n1112 B.n145 585
R1645 B.n1275 B.n1274 585
R1646 B.n1273 B.n2 585
R1647 B.n198 B.n145 516.524
R1648 B.n1110 B.n147 516.524
R1649 B.n761 B.n533 516.524
R1650 B.n757 B.n531 516.524
R1651 B.n193 B.t22 351.168
R1652 B.n582 B.t20 351.168
R1653 B.n195 B.t12 351.168
R1654 B.n580 B.t17 351.168
R1655 B.n195 B.t10 280.42
R1656 B.n193 B.t21 280.42
R1657 B.n582 B.t18 280.42
R1658 B.n580 B.t14 280.42
R1659 B.n194 B.t23 270.296
R1660 B.n583 B.t19 270.296
R1661 B.n196 B.t13 270.296
R1662 B.n581 B.t16 270.296
R1663 B.n1111 B.n191 256.663
R1664 B.n1111 B.n190 256.663
R1665 B.n1111 B.n189 256.663
R1666 B.n1111 B.n188 256.663
R1667 B.n1111 B.n187 256.663
R1668 B.n1111 B.n186 256.663
R1669 B.n1111 B.n185 256.663
R1670 B.n1111 B.n184 256.663
R1671 B.n1111 B.n183 256.663
R1672 B.n1111 B.n182 256.663
R1673 B.n1111 B.n181 256.663
R1674 B.n1111 B.n180 256.663
R1675 B.n1111 B.n179 256.663
R1676 B.n1111 B.n178 256.663
R1677 B.n1111 B.n177 256.663
R1678 B.n1111 B.n176 256.663
R1679 B.n1111 B.n175 256.663
R1680 B.n1111 B.n174 256.663
R1681 B.n1111 B.n173 256.663
R1682 B.n1111 B.n172 256.663
R1683 B.n1111 B.n171 256.663
R1684 B.n1111 B.n170 256.663
R1685 B.n1111 B.n169 256.663
R1686 B.n1111 B.n168 256.663
R1687 B.n1111 B.n167 256.663
R1688 B.n1111 B.n166 256.663
R1689 B.n1111 B.n165 256.663
R1690 B.n1111 B.n164 256.663
R1691 B.n1111 B.n163 256.663
R1692 B.n1111 B.n162 256.663
R1693 B.n1111 B.n161 256.663
R1694 B.n1111 B.n160 256.663
R1695 B.n1111 B.n159 256.663
R1696 B.n1111 B.n158 256.663
R1697 B.n1111 B.n157 256.663
R1698 B.n1111 B.n156 256.663
R1699 B.n1111 B.n155 256.663
R1700 B.n1111 B.n154 256.663
R1701 B.n1111 B.n153 256.663
R1702 B.n1111 B.n152 256.663
R1703 B.n1111 B.n151 256.663
R1704 B.n1111 B.n150 256.663
R1705 B.n1111 B.n149 256.663
R1706 B.n1111 B.n148 256.663
R1707 B.n759 B.n758 256.663
R1708 B.n759 B.n536 256.663
R1709 B.n759 B.n537 256.663
R1710 B.n759 B.n538 256.663
R1711 B.n759 B.n539 256.663
R1712 B.n759 B.n540 256.663
R1713 B.n759 B.n541 256.663
R1714 B.n759 B.n542 256.663
R1715 B.n759 B.n543 256.663
R1716 B.n759 B.n544 256.663
R1717 B.n759 B.n545 256.663
R1718 B.n759 B.n546 256.663
R1719 B.n759 B.n547 256.663
R1720 B.n759 B.n548 256.663
R1721 B.n759 B.n549 256.663
R1722 B.n759 B.n550 256.663
R1723 B.n759 B.n551 256.663
R1724 B.n759 B.n552 256.663
R1725 B.n759 B.n553 256.663
R1726 B.n759 B.n554 256.663
R1727 B.n759 B.n555 256.663
R1728 B.n759 B.n556 256.663
R1729 B.n759 B.n557 256.663
R1730 B.n759 B.n558 256.663
R1731 B.n759 B.n559 256.663
R1732 B.n759 B.n560 256.663
R1733 B.n759 B.n561 256.663
R1734 B.n759 B.n562 256.663
R1735 B.n759 B.n563 256.663
R1736 B.n759 B.n564 256.663
R1737 B.n759 B.n565 256.663
R1738 B.n759 B.n566 256.663
R1739 B.n759 B.n567 256.663
R1740 B.n759 B.n568 256.663
R1741 B.n759 B.n569 256.663
R1742 B.n759 B.n570 256.663
R1743 B.n759 B.n571 256.663
R1744 B.n759 B.n572 256.663
R1745 B.n759 B.n573 256.663
R1746 B.n759 B.n574 256.663
R1747 B.n759 B.n575 256.663
R1748 B.n759 B.n576 256.663
R1749 B.n759 B.n577 256.663
R1750 B.n760 B.n759 256.663
R1751 B.n1277 B.n1276 256.663
R1752 B.n202 B.n201 163.367
R1753 B.n206 B.n205 163.367
R1754 B.n210 B.n209 163.367
R1755 B.n214 B.n213 163.367
R1756 B.n218 B.n217 163.367
R1757 B.n222 B.n221 163.367
R1758 B.n226 B.n225 163.367
R1759 B.n230 B.n229 163.367
R1760 B.n234 B.n233 163.367
R1761 B.n238 B.n237 163.367
R1762 B.n242 B.n241 163.367
R1763 B.n246 B.n245 163.367
R1764 B.n250 B.n249 163.367
R1765 B.n254 B.n253 163.367
R1766 B.n258 B.n257 163.367
R1767 B.n262 B.n261 163.367
R1768 B.n266 B.n265 163.367
R1769 B.n270 B.n269 163.367
R1770 B.n274 B.n273 163.367
R1771 B.n278 B.n277 163.367
R1772 B.n282 B.n281 163.367
R1773 B.n286 B.n285 163.367
R1774 B.n290 B.n289 163.367
R1775 B.n294 B.n293 163.367
R1776 B.n299 B.n298 163.367
R1777 B.n303 B.n302 163.367
R1778 B.n307 B.n306 163.367
R1779 B.n311 B.n310 163.367
R1780 B.n315 B.n314 163.367
R1781 B.n319 B.n318 163.367
R1782 B.n323 B.n322 163.367
R1783 B.n327 B.n326 163.367
R1784 B.n331 B.n330 163.367
R1785 B.n335 B.n334 163.367
R1786 B.n339 B.n338 163.367
R1787 B.n343 B.n342 163.367
R1788 B.n347 B.n346 163.367
R1789 B.n351 B.n350 163.367
R1790 B.n355 B.n354 163.367
R1791 B.n359 B.n358 163.367
R1792 B.n363 B.n362 163.367
R1793 B.n367 B.n366 163.367
R1794 B.n371 B.n370 163.367
R1795 B.n1110 B.n192 163.367
R1796 B.n765 B.n533 163.367
R1797 B.n765 B.n527 163.367
R1798 B.n773 B.n527 163.367
R1799 B.n773 B.n525 163.367
R1800 B.n777 B.n525 163.367
R1801 B.n777 B.n519 163.367
R1802 B.n785 B.n519 163.367
R1803 B.n785 B.n517 163.367
R1804 B.n789 B.n517 163.367
R1805 B.n789 B.n511 163.367
R1806 B.n797 B.n511 163.367
R1807 B.n797 B.n509 163.367
R1808 B.n801 B.n509 163.367
R1809 B.n801 B.n503 163.367
R1810 B.n809 B.n503 163.367
R1811 B.n809 B.n501 163.367
R1812 B.n813 B.n501 163.367
R1813 B.n813 B.n495 163.367
R1814 B.n821 B.n495 163.367
R1815 B.n821 B.n493 163.367
R1816 B.n825 B.n493 163.367
R1817 B.n825 B.n486 163.367
R1818 B.n833 B.n486 163.367
R1819 B.n833 B.n484 163.367
R1820 B.n837 B.n484 163.367
R1821 B.n837 B.n479 163.367
R1822 B.n845 B.n479 163.367
R1823 B.n845 B.n477 163.367
R1824 B.n849 B.n477 163.367
R1825 B.n849 B.n471 163.367
R1826 B.n857 B.n471 163.367
R1827 B.n857 B.n469 163.367
R1828 B.n861 B.n469 163.367
R1829 B.n861 B.n462 163.367
R1830 B.n869 B.n462 163.367
R1831 B.n869 B.n460 163.367
R1832 B.n873 B.n460 163.367
R1833 B.n873 B.n455 163.367
R1834 B.n881 B.n455 163.367
R1835 B.n881 B.n453 163.367
R1836 B.n885 B.n453 163.367
R1837 B.n885 B.n447 163.367
R1838 B.n893 B.n447 163.367
R1839 B.n893 B.n445 163.367
R1840 B.n897 B.n445 163.367
R1841 B.n897 B.n439 163.367
R1842 B.n905 B.n439 163.367
R1843 B.n905 B.n437 163.367
R1844 B.n909 B.n437 163.367
R1845 B.n909 B.n431 163.367
R1846 B.n917 B.n431 163.367
R1847 B.n917 B.n429 163.367
R1848 B.n921 B.n429 163.367
R1849 B.n921 B.n423 163.367
R1850 B.n929 B.n423 163.367
R1851 B.n929 B.n421 163.367
R1852 B.n933 B.n421 163.367
R1853 B.n933 B.n415 163.367
R1854 B.n941 B.n415 163.367
R1855 B.n941 B.n413 163.367
R1856 B.n945 B.n413 163.367
R1857 B.n945 B.n407 163.367
R1858 B.n953 B.n407 163.367
R1859 B.n953 B.n405 163.367
R1860 B.n957 B.n405 163.367
R1861 B.n957 B.n399 163.367
R1862 B.n965 B.n399 163.367
R1863 B.n965 B.n397 163.367
R1864 B.n969 B.n397 163.367
R1865 B.n969 B.n391 163.367
R1866 B.n977 B.n391 163.367
R1867 B.n977 B.n389 163.367
R1868 B.n981 B.n389 163.367
R1869 B.n981 B.n383 163.367
R1870 B.n989 B.n383 163.367
R1871 B.n989 B.n381 163.367
R1872 B.n994 B.n381 163.367
R1873 B.n994 B.n375 163.367
R1874 B.n1002 B.n375 163.367
R1875 B.n1003 B.n1002 163.367
R1876 B.n1003 B.n5 163.367
R1877 B.n6 B.n5 163.367
R1878 B.n7 B.n6 163.367
R1879 B.n1009 B.n7 163.367
R1880 B.n1010 B.n1009 163.367
R1881 B.n1010 B.n13 163.367
R1882 B.n14 B.n13 163.367
R1883 B.n15 B.n14 163.367
R1884 B.n1015 B.n15 163.367
R1885 B.n1015 B.n20 163.367
R1886 B.n21 B.n20 163.367
R1887 B.n22 B.n21 163.367
R1888 B.n1020 B.n22 163.367
R1889 B.n1020 B.n27 163.367
R1890 B.n28 B.n27 163.367
R1891 B.n29 B.n28 163.367
R1892 B.n1025 B.n29 163.367
R1893 B.n1025 B.n34 163.367
R1894 B.n35 B.n34 163.367
R1895 B.n36 B.n35 163.367
R1896 B.n1030 B.n36 163.367
R1897 B.n1030 B.n41 163.367
R1898 B.n42 B.n41 163.367
R1899 B.n43 B.n42 163.367
R1900 B.n1035 B.n43 163.367
R1901 B.n1035 B.n48 163.367
R1902 B.n49 B.n48 163.367
R1903 B.n50 B.n49 163.367
R1904 B.n1040 B.n50 163.367
R1905 B.n1040 B.n55 163.367
R1906 B.n56 B.n55 163.367
R1907 B.n57 B.n56 163.367
R1908 B.n1045 B.n57 163.367
R1909 B.n1045 B.n62 163.367
R1910 B.n63 B.n62 163.367
R1911 B.n64 B.n63 163.367
R1912 B.n1050 B.n64 163.367
R1913 B.n1050 B.n69 163.367
R1914 B.n70 B.n69 163.367
R1915 B.n71 B.n70 163.367
R1916 B.n1055 B.n71 163.367
R1917 B.n1055 B.n76 163.367
R1918 B.n77 B.n76 163.367
R1919 B.n78 B.n77 163.367
R1920 B.n1060 B.n78 163.367
R1921 B.n1060 B.n83 163.367
R1922 B.n84 B.n83 163.367
R1923 B.n85 B.n84 163.367
R1924 B.n1065 B.n85 163.367
R1925 B.n1065 B.n90 163.367
R1926 B.n91 B.n90 163.367
R1927 B.n92 B.n91 163.367
R1928 B.n1070 B.n92 163.367
R1929 B.n1070 B.n97 163.367
R1930 B.n98 B.n97 163.367
R1931 B.n99 B.n98 163.367
R1932 B.n1075 B.n99 163.367
R1933 B.n1075 B.n104 163.367
R1934 B.n105 B.n104 163.367
R1935 B.n106 B.n105 163.367
R1936 B.n1080 B.n106 163.367
R1937 B.n1080 B.n111 163.367
R1938 B.n112 B.n111 163.367
R1939 B.n113 B.n112 163.367
R1940 B.n1085 B.n113 163.367
R1941 B.n1085 B.n118 163.367
R1942 B.n119 B.n118 163.367
R1943 B.n120 B.n119 163.367
R1944 B.n1090 B.n120 163.367
R1945 B.n1090 B.n125 163.367
R1946 B.n126 B.n125 163.367
R1947 B.n127 B.n126 163.367
R1948 B.n1095 B.n127 163.367
R1949 B.n1095 B.n132 163.367
R1950 B.n133 B.n132 163.367
R1951 B.n134 B.n133 163.367
R1952 B.n1100 B.n134 163.367
R1953 B.n1100 B.n139 163.367
R1954 B.n140 B.n139 163.367
R1955 B.n141 B.n140 163.367
R1956 B.n1105 B.n141 163.367
R1957 B.n1105 B.n146 163.367
R1958 B.n147 B.n146 163.367
R1959 B.n579 B.n578 163.367
R1960 B.n752 B.n578 163.367
R1961 B.n750 B.n749 163.367
R1962 B.n746 B.n745 163.367
R1963 B.n742 B.n741 163.367
R1964 B.n738 B.n737 163.367
R1965 B.n734 B.n733 163.367
R1966 B.n730 B.n729 163.367
R1967 B.n726 B.n725 163.367
R1968 B.n722 B.n721 163.367
R1969 B.n718 B.n717 163.367
R1970 B.n714 B.n713 163.367
R1971 B.n710 B.n709 163.367
R1972 B.n706 B.n705 163.367
R1973 B.n702 B.n701 163.367
R1974 B.n698 B.n697 163.367
R1975 B.n694 B.n693 163.367
R1976 B.n690 B.n689 163.367
R1977 B.n686 B.n685 163.367
R1978 B.n682 B.n681 163.367
R1979 B.n677 B.n676 163.367
R1980 B.n673 B.n672 163.367
R1981 B.n669 B.n668 163.367
R1982 B.n665 B.n664 163.367
R1983 B.n661 B.n660 163.367
R1984 B.n657 B.n656 163.367
R1985 B.n653 B.n652 163.367
R1986 B.n649 B.n648 163.367
R1987 B.n645 B.n644 163.367
R1988 B.n641 B.n640 163.367
R1989 B.n637 B.n636 163.367
R1990 B.n633 B.n632 163.367
R1991 B.n629 B.n628 163.367
R1992 B.n625 B.n624 163.367
R1993 B.n621 B.n620 163.367
R1994 B.n617 B.n616 163.367
R1995 B.n613 B.n612 163.367
R1996 B.n609 B.n608 163.367
R1997 B.n605 B.n604 163.367
R1998 B.n601 B.n600 163.367
R1999 B.n597 B.n596 163.367
R2000 B.n593 B.n592 163.367
R2001 B.n589 B.n588 163.367
R2002 B.n585 B.n535 163.367
R2003 B.n767 B.n531 163.367
R2004 B.n767 B.n529 163.367
R2005 B.n771 B.n529 163.367
R2006 B.n771 B.n523 163.367
R2007 B.n779 B.n523 163.367
R2008 B.n779 B.n521 163.367
R2009 B.n783 B.n521 163.367
R2010 B.n783 B.n515 163.367
R2011 B.n791 B.n515 163.367
R2012 B.n791 B.n513 163.367
R2013 B.n795 B.n513 163.367
R2014 B.n795 B.n507 163.367
R2015 B.n803 B.n507 163.367
R2016 B.n803 B.n505 163.367
R2017 B.n807 B.n505 163.367
R2018 B.n807 B.n499 163.367
R2019 B.n815 B.n499 163.367
R2020 B.n815 B.n497 163.367
R2021 B.n819 B.n497 163.367
R2022 B.n819 B.n491 163.367
R2023 B.n827 B.n491 163.367
R2024 B.n827 B.n489 163.367
R2025 B.n831 B.n489 163.367
R2026 B.n831 B.n483 163.367
R2027 B.n839 B.n483 163.367
R2028 B.n839 B.n481 163.367
R2029 B.n843 B.n481 163.367
R2030 B.n843 B.n475 163.367
R2031 B.n851 B.n475 163.367
R2032 B.n851 B.n473 163.367
R2033 B.n855 B.n473 163.367
R2034 B.n855 B.n467 163.367
R2035 B.n863 B.n467 163.367
R2036 B.n863 B.n465 163.367
R2037 B.n867 B.n465 163.367
R2038 B.n867 B.n459 163.367
R2039 B.n875 B.n459 163.367
R2040 B.n875 B.n457 163.367
R2041 B.n879 B.n457 163.367
R2042 B.n879 B.n451 163.367
R2043 B.n887 B.n451 163.367
R2044 B.n887 B.n449 163.367
R2045 B.n891 B.n449 163.367
R2046 B.n891 B.n443 163.367
R2047 B.n899 B.n443 163.367
R2048 B.n899 B.n441 163.367
R2049 B.n903 B.n441 163.367
R2050 B.n903 B.n435 163.367
R2051 B.n911 B.n435 163.367
R2052 B.n911 B.n433 163.367
R2053 B.n915 B.n433 163.367
R2054 B.n915 B.n427 163.367
R2055 B.n923 B.n427 163.367
R2056 B.n923 B.n425 163.367
R2057 B.n927 B.n425 163.367
R2058 B.n927 B.n419 163.367
R2059 B.n935 B.n419 163.367
R2060 B.n935 B.n417 163.367
R2061 B.n939 B.n417 163.367
R2062 B.n939 B.n411 163.367
R2063 B.n947 B.n411 163.367
R2064 B.n947 B.n409 163.367
R2065 B.n951 B.n409 163.367
R2066 B.n951 B.n403 163.367
R2067 B.n959 B.n403 163.367
R2068 B.n959 B.n401 163.367
R2069 B.n963 B.n401 163.367
R2070 B.n963 B.n395 163.367
R2071 B.n971 B.n395 163.367
R2072 B.n971 B.n393 163.367
R2073 B.n975 B.n393 163.367
R2074 B.n975 B.n387 163.367
R2075 B.n983 B.n387 163.367
R2076 B.n983 B.n385 163.367
R2077 B.n987 B.n385 163.367
R2078 B.n987 B.n379 163.367
R2079 B.n996 B.n379 163.367
R2080 B.n996 B.n377 163.367
R2081 B.n1000 B.n377 163.367
R2082 B.n1000 B.n3 163.367
R2083 B.n1275 B.n3 163.367
R2084 B.n1271 B.n2 163.367
R2085 B.n1271 B.n1270 163.367
R2086 B.n1270 B.n9 163.367
R2087 B.n1266 B.n9 163.367
R2088 B.n1266 B.n11 163.367
R2089 B.n1262 B.n11 163.367
R2090 B.n1262 B.n17 163.367
R2091 B.n1258 B.n17 163.367
R2092 B.n1258 B.n19 163.367
R2093 B.n1254 B.n19 163.367
R2094 B.n1254 B.n24 163.367
R2095 B.n1250 B.n24 163.367
R2096 B.n1250 B.n26 163.367
R2097 B.n1246 B.n26 163.367
R2098 B.n1246 B.n31 163.367
R2099 B.n1242 B.n31 163.367
R2100 B.n1242 B.n33 163.367
R2101 B.n1238 B.n33 163.367
R2102 B.n1238 B.n38 163.367
R2103 B.n1234 B.n38 163.367
R2104 B.n1234 B.n40 163.367
R2105 B.n1230 B.n40 163.367
R2106 B.n1230 B.n45 163.367
R2107 B.n1226 B.n45 163.367
R2108 B.n1226 B.n47 163.367
R2109 B.n1222 B.n47 163.367
R2110 B.n1222 B.n52 163.367
R2111 B.n1218 B.n52 163.367
R2112 B.n1218 B.n54 163.367
R2113 B.n1214 B.n54 163.367
R2114 B.n1214 B.n59 163.367
R2115 B.n1210 B.n59 163.367
R2116 B.n1210 B.n61 163.367
R2117 B.n1206 B.n61 163.367
R2118 B.n1206 B.n66 163.367
R2119 B.n1202 B.n66 163.367
R2120 B.n1202 B.n68 163.367
R2121 B.n1198 B.n68 163.367
R2122 B.n1198 B.n73 163.367
R2123 B.n1194 B.n73 163.367
R2124 B.n1194 B.n75 163.367
R2125 B.n1190 B.n75 163.367
R2126 B.n1190 B.n80 163.367
R2127 B.n1186 B.n80 163.367
R2128 B.n1186 B.n82 163.367
R2129 B.n1182 B.n82 163.367
R2130 B.n1182 B.n87 163.367
R2131 B.n1178 B.n87 163.367
R2132 B.n1178 B.n89 163.367
R2133 B.n1174 B.n89 163.367
R2134 B.n1174 B.n94 163.367
R2135 B.n1170 B.n94 163.367
R2136 B.n1170 B.n96 163.367
R2137 B.n1166 B.n96 163.367
R2138 B.n1166 B.n101 163.367
R2139 B.n1162 B.n101 163.367
R2140 B.n1162 B.n103 163.367
R2141 B.n1158 B.n103 163.367
R2142 B.n1158 B.n108 163.367
R2143 B.n1154 B.n108 163.367
R2144 B.n1154 B.n110 163.367
R2145 B.n1150 B.n110 163.367
R2146 B.n1150 B.n115 163.367
R2147 B.n1146 B.n115 163.367
R2148 B.n1146 B.n117 163.367
R2149 B.n1142 B.n117 163.367
R2150 B.n1142 B.n122 163.367
R2151 B.n1138 B.n122 163.367
R2152 B.n1138 B.n124 163.367
R2153 B.n1134 B.n124 163.367
R2154 B.n1134 B.n129 163.367
R2155 B.n1130 B.n129 163.367
R2156 B.n1130 B.n131 163.367
R2157 B.n1126 B.n131 163.367
R2158 B.n1126 B.n136 163.367
R2159 B.n1122 B.n136 163.367
R2160 B.n1122 B.n138 163.367
R2161 B.n1118 B.n138 163.367
R2162 B.n1118 B.n143 163.367
R2163 B.n1114 B.n143 163.367
R2164 B.n1114 B.n145 163.367
R2165 B.n759 B.n532 90.811
R2166 B.n1112 B.n1111 90.811
R2167 B.n196 B.n195 80.8732
R2168 B.n194 B.n193 80.8732
R2169 B.n583 B.n582 80.8732
R2170 B.n581 B.n580 80.8732
R2171 B.n198 B.n148 71.676
R2172 B.n202 B.n149 71.676
R2173 B.n206 B.n150 71.676
R2174 B.n210 B.n151 71.676
R2175 B.n214 B.n152 71.676
R2176 B.n218 B.n153 71.676
R2177 B.n222 B.n154 71.676
R2178 B.n226 B.n155 71.676
R2179 B.n230 B.n156 71.676
R2180 B.n234 B.n157 71.676
R2181 B.n238 B.n158 71.676
R2182 B.n242 B.n159 71.676
R2183 B.n246 B.n160 71.676
R2184 B.n250 B.n161 71.676
R2185 B.n254 B.n162 71.676
R2186 B.n258 B.n163 71.676
R2187 B.n262 B.n164 71.676
R2188 B.n266 B.n165 71.676
R2189 B.n270 B.n166 71.676
R2190 B.n274 B.n167 71.676
R2191 B.n278 B.n168 71.676
R2192 B.n282 B.n169 71.676
R2193 B.n286 B.n170 71.676
R2194 B.n290 B.n171 71.676
R2195 B.n294 B.n172 71.676
R2196 B.n299 B.n173 71.676
R2197 B.n303 B.n174 71.676
R2198 B.n307 B.n175 71.676
R2199 B.n311 B.n176 71.676
R2200 B.n315 B.n177 71.676
R2201 B.n319 B.n178 71.676
R2202 B.n323 B.n179 71.676
R2203 B.n327 B.n180 71.676
R2204 B.n331 B.n181 71.676
R2205 B.n335 B.n182 71.676
R2206 B.n339 B.n183 71.676
R2207 B.n343 B.n184 71.676
R2208 B.n347 B.n185 71.676
R2209 B.n351 B.n186 71.676
R2210 B.n355 B.n187 71.676
R2211 B.n359 B.n188 71.676
R2212 B.n363 B.n189 71.676
R2213 B.n367 B.n190 71.676
R2214 B.n371 B.n191 71.676
R2215 B.n192 B.n191 71.676
R2216 B.n370 B.n190 71.676
R2217 B.n366 B.n189 71.676
R2218 B.n362 B.n188 71.676
R2219 B.n358 B.n187 71.676
R2220 B.n354 B.n186 71.676
R2221 B.n350 B.n185 71.676
R2222 B.n346 B.n184 71.676
R2223 B.n342 B.n183 71.676
R2224 B.n338 B.n182 71.676
R2225 B.n334 B.n181 71.676
R2226 B.n330 B.n180 71.676
R2227 B.n326 B.n179 71.676
R2228 B.n322 B.n178 71.676
R2229 B.n318 B.n177 71.676
R2230 B.n314 B.n176 71.676
R2231 B.n310 B.n175 71.676
R2232 B.n306 B.n174 71.676
R2233 B.n302 B.n173 71.676
R2234 B.n298 B.n172 71.676
R2235 B.n293 B.n171 71.676
R2236 B.n289 B.n170 71.676
R2237 B.n285 B.n169 71.676
R2238 B.n281 B.n168 71.676
R2239 B.n277 B.n167 71.676
R2240 B.n273 B.n166 71.676
R2241 B.n269 B.n165 71.676
R2242 B.n265 B.n164 71.676
R2243 B.n261 B.n163 71.676
R2244 B.n257 B.n162 71.676
R2245 B.n253 B.n161 71.676
R2246 B.n249 B.n160 71.676
R2247 B.n245 B.n159 71.676
R2248 B.n241 B.n158 71.676
R2249 B.n237 B.n157 71.676
R2250 B.n233 B.n156 71.676
R2251 B.n229 B.n155 71.676
R2252 B.n225 B.n154 71.676
R2253 B.n221 B.n153 71.676
R2254 B.n217 B.n152 71.676
R2255 B.n213 B.n151 71.676
R2256 B.n209 B.n150 71.676
R2257 B.n205 B.n149 71.676
R2258 B.n201 B.n148 71.676
R2259 B.n758 B.n757 71.676
R2260 B.n752 B.n536 71.676
R2261 B.n749 B.n537 71.676
R2262 B.n745 B.n538 71.676
R2263 B.n741 B.n539 71.676
R2264 B.n737 B.n540 71.676
R2265 B.n733 B.n541 71.676
R2266 B.n729 B.n542 71.676
R2267 B.n725 B.n543 71.676
R2268 B.n721 B.n544 71.676
R2269 B.n717 B.n545 71.676
R2270 B.n713 B.n546 71.676
R2271 B.n709 B.n547 71.676
R2272 B.n705 B.n548 71.676
R2273 B.n701 B.n549 71.676
R2274 B.n697 B.n550 71.676
R2275 B.n693 B.n551 71.676
R2276 B.n689 B.n552 71.676
R2277 B.n685 B.n553 71.676
R2278 B.n681 B.n554 71.676
R2279 B.n676 B.n555 71.676
R2280 B.n672 B.n556 71.676
R2281 B.n668 B.n557 71.676
R2282 B.n664 B.n558 71.676
R2283 B.n660 B.n559 71.676
R2284 B.n656 B.n560 71.676
R2285 B.n652 B.n561 71.676
R2286 B.n648 B.n562 71.676
R2287 B.n644 B.n563 71.676
R2288 B.n640 B.n564 71.676
R2289 B.n636 B.n565 71.676
R2290 B.n632 B.n566 71.676
R2291 B.n628 B.n567 71.676
R2292 B.n624 B.n568 71.676
R2293 B.n620 B.n569 71.676
R2294 B.n616 B.n570 71.676
R2295 B.n612 B.n571 71.676
R2296 B.n608 B.n572 71.676
R2297 B.n604 B.n573 71.676
R2298 B.n600 B.n574 71.676
R2299 B.n596 B.n575 71.676
R2300 B.n592 B.n576 71.676
R2301 B.n588 B.n577 71.676
R2302 B.n760 B.n535 71.676
R2303 B.n758 B.n579 71.676
R2304 B.n750 B.n536 71.676
R2305 B.n746 B.n537 71.676
R2306 B.n742 B.n538 71.676
R2307 B.n738 B.n539 71.676
R2308 B.n734 B.n540 71.676
R2309 B.n730 B.n541 71.676
R2310 B.n726 B.n542 71.676
R2311 B.n722 B.n543 71.676
R2312 B.n718 B.n544 71.676
R2313 B.n714 B.n545 71.676
R2314 B.n710 B.n546 71.676
R2315 B.n706 B.n547 71.676
R2316 B.n702 B.n548 71.676
R2317 B.n698 B.n549 71.676
R2318 B.n694 B.n550 71.676
R2319 B.n690 B.n551 71.676
R2320 B.n686 B.n552 71.676
R2321 B.n682 B.n553 71.676
R2322 B.n677 B.n554 71.676
R2323 B.n673 B.n555 71.676
R2324 B.n669 B.n556 71.676
R2325 B.n665 B.n557 71.676
R2326 B.n661 B.n558 71.676
R2327 B.n657 B.n559 71.676
R2328 B.n653 B.n560 71.676
R2329 B.n649 B.n561 71.676
R2330 B.n645 B.n562 71.676
R2331 B.n641 B.n563 71.676
R2332 B.n637 B.n564 71.676
R2333 B.n633 B.n565 71.676
R2334 B.n629 B.n566 71.676
R2335 B.n625 B.n567 71.676
R2336 B.n621 B.n568 71.676
R2337 B.n617 B.n569 71.676
R2338 B.n613 B.n570 71.676
R2339 B.n609 B.n571 71.676
R2340 B.n605 B.n572 71.676
R2341 B.n601 B.n573 71.676
R2342 B.n597 B.n574 71.676
R2343 B.n593 B.n575 71.676
R2344 B.n589 B.n576 71.676
R2345 B.n585 B.n577 71.676
R2346 B.n761 B.n760 71.676
R2347 B.n1276 B.n1275 71.676
R2348 B.n1276 B.n2 71.676
R2349 B.n197 B.n196 59.5399
R2350 B.n296 B.n194 59.5399
R2351 B.n584 B.n583 59.5399
R2352 B.n679 B.n581 59.5399
R2353 B.n766 B.n532 45.0743
R2354 B.n766 B.n528 45.0743
R2355 B.n772 B.n528 45.0743
R2356 B.n772 B.n524 45.0743
R2357 B.n778 B.n524 45.0743
R2358 B.n778 B.n520 45.0743
R2359 B.n784 B.n520 45.0743
R2360 B.n784 B.n516 45.0743
R2361 B.n790 B.n516 45.0743
R2362 B.n796 B.n512 45.0743
R2363 B.n796 B.n508 45.0743
R2364 B.n802 B.n508 45.0743
R2365 B.n802 B.n504 45.0743
R2366 B.n808 B.n504 45.0743
R2367 B.n808 B.n500 45.0743
R2368 B.n814 B.n500 45.0743
R2369 B.n814 B.n496 45.0743
R2370 B.n820 B.n496 45.0743
R2371 B.n820 B.n492 45.0743
R2372 B.n826 B.n492 45.0743
R2373 B.n826 B.n487 45.0743
R2374 B.n832 B.n487 45.0743
R2375 B.n832 B.n488 45.0743
R2376 B.n838 B.n480 45.0743
R2377 B.n844 B.n480 45.0743
R2378 B.n844 B.n476 45.0743
R2379 B.n850 B.n476 45.0743
R2380 B.n850 B.n472 45.0743
R2381 B.n856 B.n472 45.0743
R2382 B.n856 B.n468 45.0743
R2383 B.n862 B.n468 45.0743
R2384 B.n862 B.n463 45.0743
R2385 B.n868 B.n463 45.0743
R2386 B.n868 B.n464 45.0743
R2387 B.n874 B.n456 45.0743
R2388 B.n880 B.n456 45.0743
R2389 B.n880 B.n452 45.0743
R2390 B.n886 B.n452 45.0743
R2391 B.n886 B.n448 45.0743
R2392 B.n892 B.n448 45.0743
R2393 B.n892 B.n444 45.0743
R2394 B.n898 B.n444 45.0743
R2395 B.n898 B.n440 45.0743
R2396 B.n904 B.n440 45.0743
R2397 B.n904 B.n436 45.0743
R2398 B.n910 B.n436 45.0743
R2399 B.n916 B.n432 45.0743
R2400 B.n916 B.n428 45.0743
R2401 B.n922 B.n428 45.0743
R2402 B.n922 B.n424 45.0743
R2403 B.n928 B.n424 45.0743
R2404 B.n928 B.n420 45.0743
R2405 B.n934 B.n420 45.0743
R2406 B.n934 B.n416 45.0743
R2407 B.n940 B.n416 45.0743
R2408 B.n940 B.n412 45.0743
R2409 B.n946 B.n412 45.0743
R2410 B.n952 B.n408 45.0743
R2411 B.n952 B.n404 45.0743
R2412 B.n958 B.n404 45.0743
R2413 B.n958 B.n400 45.0743
R2414 B.n964 B.n400 45.0743
R2415 B.n964 B.n396 45.0743
R2416 B.n970 B.n396 45.0743
R2417 B.n970 B.n392 45.0743
R2418 B.n976 B.n392 45.0743
R2419 B.n976 B.n388 45.0743
R2420 B.n982 B.n388 45.0743
R2421 B.n988 B.n384 45.0743
R2422 B.n988 B.n380 45.0743
R2423 B.n995 B.n380 45.0743
R2424 B.n995 B.n376 45.0743
R2425 B.n1001 B.n376 45.0743
R2426 B.n1001 B.n4 45.0743
R2427 B.n1274 B.n4 45.0743
R2428 B.n1274 B.n1273 45.0743
R2429 B.n1273 B.n1272 45.0743
R2430 B.n1272 B.n8 45.0743
R2431 B.n12 B.n8 45.0743
R2432 B.n1265 B.n12 45.0743
R2433 B.n1265 B.n1264 45.0743
R2434 B.n1264 B.n1263 45.0743
R2435 B.n1263 B.n16 45.0743
R2436 B.n1257 B.n1256 45.0743
R2437 B.n1256 B.n1255 45.0743
R2438 B.n1255 B.n23 45.0743
R2439 B.n1249 B.n23 45.0743
R2440 B.n1249 B.n1248 45.0743
R2441 B.n1248 B.n1247 45.0743
R2442 B.n1247 B.n30 45.0743
R2443 B.n1241 B.n30 45.0743
R2444 B.n1241 B.n1240 45.0743
R2445 B.n1240 B.n1239 45.0743
R2446 B.n1239 B.n37 45.0743
R2447 B.n1233 B.n1232 45.0743
R2448 B.n1232 B.n1231 45.0743
R2449 B.n1231 B.n44 45.0743
R2450 B.n1225 B.n44 45.0743
R2451 B.n1225 B.n1224 45.0743
R2452 B.n1224 B.n1223 45.0743
R2453 B.n1223 B.n51 45.0743
R2454 B.n1217 B.n51 45.0743
R2455 B.n1217 B.n1216 45.0743
R2456 B.n1216 B.n1215 45.0743
R2457 B.n1215 B.n58 45.0743
R2458 B.n1209 B.n1208 45.0743
R2459 B.n1208 B.n1207 45.0743
R2460 B.n1207 B.n65 45.0743
R2461 B.n1201 B.n65 45.0743
R2462 B.n1201 B.n1200 45.0743
R2463 B.n1200 B.n1199 45.0743
R2464 B.n1199 B.n72 45.0743
R2465 B.n1193 B.n72 45.0743
R2466 B.n1193 B.n1192 45.0743
R2467 B.n1192 B.n1191 45.0743
R2468 B.n1191 B.n79 45.0743
R2469 B.n1185 B.n79 45.0743
R2470 B.n1184 B.n1183 45.0743
R2471 B.n1183 B.n86 45.0743
R2472 B.n1177 B.n86 45.0743
R2473 B.n1177 B.n1176 45.0743
R2474 B.n1176 B.n1175 45.0743
R2475 B.n1175 B.n93 45.0743
R2476 B.n1169 B.n93 45.0743
R2477 B.n1169 B.n1168 45.0743
R2478 B.n1168 B.n1167 45.0743
R2479 B.n1167 B.n100 45.0743
R2480 B.n1161 B.n100 45.0743
R2481 B.n1160 B.n1159 45.0743
R2482 B.n1159 B.n107 45.0743
R2483 B.n1153 B.n107 45.0743
R2484 B.n1153 B.n1152 45.0743
R2485 B.n1152 B.n1151 45.0743
R2486 B.n1151 B.n114 45.0743
R2487 B.n1145 B.n114 45.0743
R2488 B.n1145 B.n1144 45.0743
R2489 B.n1144 B.n1143 45.0743
R2490 B.n1143 B.n121 45.0743
R2491 B.n1137 B.n121 45.0743
R2492 B.n1137 B.n1136 45.0743
R2493 B.n1136 B.n1135 45.0743
R2494 B.n1135 B.n128 45.0743
R2495 B.n1129 B.n1128 45.0743
R2496 B.n1128 B.n1127 45.0743
R2497 B.n1127 B.n135 45.0743
R2498 B.n1121 B.n135 45.0743
R2499 B.n1121 B.n1120 45.0743
R2500 B.n1120 B.n1119 45.0743
R2501 B.n1119 B.n142 45.0743
R2502 B.n1113 B.n142 45.0743
R2503 B.n1113 B.n1112 45.0743
R2504 B.n464 B.t7 43.7486
R2505 B.t6 B.n1184 43.7486
R2506 B.t15 B.n512 34.4687
R2507 B.t0 B.n432 34.4687
R2508 B.n982 B.t3 34.4687
R2509 B.n1257 B.t8 34.4687
R2510 B.t4 B.n58 34.4687
R2511 B.t11 B.n128 34.4687
R2512 B.n756 B.n530 33.5615
R2513 B.n763 B.n762 33.5615
R2514 B.n1109 B.n1108 33.5615
R2515 B.n199 B.n144 33.5615
R2516 B.n488 B.t1 31.8173
R2517 B.t5 B.n1160 31.8173
R2518 B.n946 B.t9 22.5374
R2519 B.t9 B.n408 22.5374
R2520 B.t2 B.n37 22.5374
R2521 B.n1233 B.t2 22.5374
R2522 B B.n1277 18.0485
R2523 B.n838 B.t1 13.2575
R2524 B.n1161 B.t5 13.2575
R2525 B.n768 B.n530 10.6151
R2526 B.n769 B.n768 10.6151
R2527 B.n770 B.n769 10.6151
R2528 B.n770 B.n522 10.6151
R2529 B.n780 B.n522 10.6151
R2530 B.n781 B.n780 10.6151
R2531 B.n782 B.n781 10.6151
R2532 B.n782 B.n514 10.6151
R2533 B.n792 B.n514 10.6151
R2534 B.n793 B.n792 10.6151
R2535 B.n794 B.n793 10.6151
R2536 B.n794 B.n506 10.6151
R2537 B.n804 B.n506 10.6151
R2538 B.n805 B.n804 10.6151
R2539 B.n806 B.n805 10.6151
R2540 B.n806 B.n498 10.6151
R2541 B.n816 B.n498 10.6151
R2542 B.n817 B.n816 10.6151
R2543 B.n818 B.n817 10.6151
R2544 B.n818 B.n490 10.6151
R2545 B.n828 B.n490 10.6151
R2546 B.n829 B.n828 10.6151
R2547 B.n830 B.n829 10.6151
R2548 B.n830 B.n482 10.6151
R2549 B.n840 B.n482 10.6151
R2550 B.n841 B.n840 10.6151
R2551 B.n842 B.n841 10.6151
R2552 B.n842 B.n474 10.6151
R2553 B.n852 B.n474 10.6151
R2554 B.n853 B.n852 10.6151
R2555 B.n854 B.n853 10.6151
R2556 B.n854 B.n466 10.6151
R2557 B.n864 B.n466 10.6151
R2558 B.n865 B.n864 10.6151
R2559 B.n866 B.n865 10.6151
R2560 B.n866 B.n458 10.6151
R2561 B.n876 B.n458 10.6151
R2562 B.n877 B.n876 10.6151
R2563 B.n878 B.n877 10.6151
R2564 B.n878 B.n450 10.6151
R2565 B.n888 B.n450 10.6151
R2566 B.n889 B.n888 10.6151
R2567 B.n890 B.n889 10.6151
R2568 B.n890 B.n442 10.6151
R2569 B.n900 B.n442 10.6151
R2570 B.n901 B.n900 10.6151
R2571 B.n902 B.n901 10.6151
R2572 B.n902 B.n434 10.6151
R2573 B.n912 B.n434 10.6151
R2574 B.n913 B.n912 10.6151
R2575 B.n914 B.n913 10.6151
R2576 B.n914 B.n426 10.6151
R2577 B.n924 B.n426 10.6151
R2578 B.n925 B.n924 10.6151
R2579 B.n926 B.n925 10.6151
R2580 B.n926 B.n418 10.6151
R2581 B.n936 B.n418 10.6151
R2582 B.n937 B.n936 10.6151
R2583 B.n938 B.n937 10.6151
R2584 B.n938 B.n410 10.6151
R2585 B.n948 B.n410 10.6151
R2586 B.n949 B.n948 10.6151
R2587 B.n950 B.n949 10.6151
R2588 B.n950 B.n402 10.6151
R2589 B.n960 B.n402 10.6151
R2590 B.n961 B.n960 10.6151
R2591 B.n962 B.n961 10.6151
R2592 B.n962 B.n394 10.6151
R2593 B.n972 B.n394 10.6151
R2594 B.n973 B.n972 10.6151
R2595 B.n974 B.n973 10.6151
R2596 B.n974 B.n386 10.6151
R2597 B.n984 B.n386 10.6151
R2598 B.n985 B.n984 10.6151
R2599 B.n986 B.n985 10.6151
R2600 B.n986 B.n378 10.6151
R2601 B.n997 B.n378 10.6151
R2602 B.n998 B.n997 10.6151
R2603 B.n999 B.n998 10.6151
R2604 B.n999 B.n0 10.6151
R2605 B.n756 B.n755 10.6151
R2606 B.n755 B.n754 10.6151
R2607 B.n754 B.n753 10.6151
R2608 B.n753 B.n751 10.6151
R2609 B.n751 B.n748 10.6151
R2610 B.n748 B.n747 10.6151
R2611 B.n747 B.n744 10.6151
R2612 B.n744 B.n743 10.6151
R2613 B.n743 B.n740 10.6151
R2614 B.n740 B.n739 10.6151
R2615 B.n739 B.n736 10.6151
R2616 B.n736 B.n735 10.6151
R2617 B.n735 B.n732 10.6151
R2618 B.n732 B.n731 10.6151
R2619 B.n731 B.n728 10.6151
R2620 B.n728 B.n727 10.6151
R2621 B.n727 B.n724 10.6151
R2622 B.n724 B.n723 10.6151
R2623 B.n723 B.n720 10.6151
R2624 B.n720 B.n719 10.6151
R2625 B.n719 B.n716 10.6151
R2626 B.n716 B.n715 10.6151
R2627 B.n715 B.n712 10.6151
R2628 B.n712 B.n711 10.6151
R2629 B.n711 B.n708 10.6151
R2630 B.n708 B.n707 10.6151
R2631 B.n707 B.n704 10.6151
R2632 B.n704 B.n703 10.6151
R2633 B.n703 B.n700 10.6151
R2634 B.n700 B.n699 10.6151
R2635 B.n699 B.n696 10.6151
R2636 B.n696 B.n695 10.6151
R2637 B.n695 B.n692 10.6151
R2638 B.n692 B.n691 10.6151
R2639 B.n691 B.n688 10.6151
R2640 B.n688 B.n687 10.6151
R2641 B.n687 B.n684 10.6151
R2642 B.n684 B.n683 10.6151
R2643 B.n683 B.n680 10.6151
R2644 B.n678 B.n675 10.6151
R2645 B.n675 B.n674 10.6151
R2646 B.n674 B.n671 10.6151
R2647 B.n671 B.n670 10.6151
R2648 B.n670 B.n667 10.6151
R2649 B.n667 B.n666 10.6151
R2650 B.n666 B.n663 10.6151
R2651 B.n663 B.n662 10.6151
R2652 B.n659 B.n658 10.6151
R2653 B.n658 B.n655 10.6151
R2654 B.n655 B.n654 10.6151
R2655 B.n654 B.n651 10.6151
R2656 B.n651 B.n650 10.6151
R2657 B.n650 B.n647 10.6151
R2658 B.n647 B.n646 10.6151
R2659 B.n646 B.n643 10.6151
R2660 B.n643 B.n642 10.6151
R2661 B.n642 B.n639 10.6151
R2662 B.n639 B.n638 10.6151
R2663 B.n638 B.n635 10.6151
R2664 B.n635 B.n634 10.6151
R2665 B.n634 B.n631 10.6151
R2666 B.n631 B.n630 10.6151
R2667 B.n630 B.n627 10.6151
R2668 B.n627 B.n626 10.6151
R2669 B.n626 B.n623 10.6151
R2670 B.n623 B.n622 10.6151
R2671 B.n622 B.n619 10.6151
R2672 B.n619 B.n618 10.6151
R2673 B.n618 B.n615 10.6151
R2674 B.n615 B.n614 10.6151
R2675 B.n614 B.n611 10.6151
R2676 B.n611 B.n610 10.6151
R2677 B.n610 B.n607 10.6151
R2678 B.n607 B.n606 10.6151
R2679 B.n606 B.n603 10.6151
R2680 B.n603 B.n602 10.6151
R2681 B.n602 B.n599 10.6151
R2682 B.n599 B.n598 10.6151
R2683 B.n598 B.n595 10.6151
R2684 B.n595 B.n594 10.6151
R2685 B.n594 B.n591 10.6151
R2686 B.n591 B.n590 10.6151
R2687 B.n590 B.n587 10.6151
R2688 B.n587 B.n586 10.6151
R2689 B.n586 B.n534 10.6151
R2690 B.n762 B.n534 10.6151
R2691 B.n764 B.n763 10.6151
R2692 B.n764 B.n526 10.6151
R2693 B.n774 B.n526 10.6151
R2694 B.n775 B.n774 10.6151
R2695 B.n776 B.n775 10.6151
R2696 B.n776 B.n518 10.6151
R2697 B.n786 B.n518 10.6151
R2698 B.n787 B.n786 10.6151
R2699 B.n788 B.n787 10.6151
R2700 B.n788 B.n510 10.6151
R2701 B.n798 B.n510 10.6151
R2702 B.n799 B.n798 10.6151
R2703 B.n800 B.n799 10.6151
R2704 B.n800 B.n502 10.6151
R2705 B.n810 B.n502 10.6151
R2706 B.n811 B.n810 10.6151
R2707 B.n812 B.n811 10.6151
R2708 B.n812 B.n494 10.6151
R2709 B.n822 B.n494 10.6151
R2710 B.n823 B.n822 10.6151
R2711 B.n824 B.n823 10.6151
R2712 B.n824 B.n485 10.6151
R2713 B.n834 B.n485 10.6151
R2714 B.n835 B.n834 10.6151
R2715 B.n836 B.n835 10.6151
R2716 B.n836 B.n478 10.6151
R2717 B.n846 B.n478 10.6151
R2718 B.n847 B.n846 10.6151
R2719 B.n848 B.n847 10.6151
R2720 B.n848 B.n470 10.6151
R2721 B.n858 B.n470 10.6151
R2722 B.n859 B.n858 10.6151
R2723 B.n860 B.n859 10.6151
R2724 B.n860 B.n461 10.6151
R2725 B.n870 B.n461 10.6151
R2726 B.n871 B.n870 10.6151
R2727 B.n872 B.n871 10.6151
R2728 B.n872 B.n454 10.6151
R2729 B.n882 B.n454 10.6151
R2730 B.n883 B.n882 10.6151
R2731 B.n884 B.n883 10.6151
R2732 B.n884 B.n446 10.6151
R2733 B.n894 B.n446 10.6151
R2734 B.n895 B.n894 10.6151
R2735 B.n896 B.n895 10.6151
R2736 B.n896 B.n438 10.6151
R2737 B.n906 B.n438 10.6151
R2738 B.n907 B.n906 10.6151
R2739 B.n908 B.n907 10.6151
R2740 B.n908 B.n430 10.6151
R2741 B.n918 B.n430 10.6151
R2742 B.n919 B.n918 10.6151
R2743 B.n920 B.n919 10.6151
R2744 B.n920 B.n422 10.6151
R2745 B.n930 B.n422 10.6151
R2746 B.n931 B.n930 10.6151
R2747 B.n932 B.n931 10.6151
R2748 B.n932 B.n414 10.6151
R2749 B.n942 B.n414 10.6151
R2750 B.n943 B.n942 10.6151
R2751 B.n944 B.n943 10.6151
R2752 B.n944 B.n406 10.6151
R2753 B.n954 B.n406 10.6151
R2754 B.n955 B.n954 10.6151
R2755 B.n956 B.n955 10.6151
R2756 B.n956 B.n398 10.6151
R2757 B.n966 B.n398 10.6151
R2758 B.n967 B.n966 10.6151
R2759 B.n968 B.n967 10.6151
R2760 B.n968 B.n390 10.6151
R2761 B.n978 B.n390 10.6151
R2762 B.n979 B.n978 10.6151
R2763 B.n980 B.n979 10.6151
R2764 B.n980 B.n382 10.6151
R2765 B.n990 B.n382 10.6151
R2766 B.n991 B.n990 10.6151
R2767 B.n993 B.n991 10.6151
R2768 B.n993 B.n992 10.6151
R2769 B.n992 B.n374 10.6151
R2770 B.n1004 B.n374 10.6151
R2771 B.n1005 B.n1004 10.6151
R2772 B.n1006 B.n1005 10.6151
R2773 B.n1007 B.n1006 10.6151
R2774 B.n1008 B.n1007 10.6151
R2775 B.n1011 B.n1008 10.6151
R2776 B.n1012 B.n1011 10.6151
R2777 B.n1013 B.n1012 10.6151
R2778 B.n1014 B.n1013 10.6151
R2779 B.n1016 B.n1014 10.6151
R2780 B.n1017 B.n1016 10.6151
R2781 B.n1018 B.n1017 10.6151
R2782 B.n1019 B.n1018 10.6151
R2783 B.n1021 B.n1019 10.6151
R2784 B.n1022 B.n1021 10.6151
R2785 B.n1023 B.n1022 10.6151
R2786 B.n1024 B.n1023 10.6151
R2787 B.n1026 B.n1024 10.6151
R2788 B.n1027 B.n1026 10.6151
R2789 B.n1028 B.n1027 10.6151
R2790 B.n1029 B.n1028 10.6151
R2791 B.n1031 B.n1029 10.6151
R2792 B.n1032 B.n1031 10.6151
R2793 B.n1033 B.n1032 10.6151
R2794 B.n1034 B.n1033 10.6151
R2795 B.n1036 B.n1034 10.6151
R2796 B.n1037 B.n1036 10.6151
R2797 B.n1038 B.n1037 10.6151
R2798 B.n1039 B.n1038 10.6151
R2799 B.n1041 B.n1039 10.6151
R2800 B.n1042 B.n1041 10.6151
R2801 B.n1043 B.n1042 10.6151
R2802 B.n1044 B.n1043 10.6151
R2803 B.n1046 B.n1044 10.6151
R2804 B.n1047 B.n1046 10.6151
R2805 B.n1048 B.n1047 10.6151
R2806 B.n1049 B.n1048 10.6151
R2807 B.n1051 B.n1049 10.6151
R2808 B.n1052 B.n1051 10.6151
R2809 B.n1053 B.n1052 10.6151
R2810 B.n1054 B.n1053 10.6151
R2811 B.n1056 B.n1054 10.6151
R2812 B.n1057 B.n1056 10.6151
R2813 B.n1058 B.n1057 10.6151
R2814 B.n1059 B.n1058 10.6151
R2815 B.n1061 B.n1059 10.6151
R2816 B.n1062 B.n1061 10.6151
R2817 B.n1063 B.n1062 10.6151
R2818 B.n1064 B.n1063 10.6151
R2819 B.n1066 B.n1064 10.6151
R2820 B.n1067 B.n1066 10.6151
R2821 B.n1068 B.n1067 10.6151
R2822 B.n1069 B.n1068 10.6151
R2823 B.n1071 B.n1069 10.6151
R2824 B.n1072 B.n1071 10.6151
R2825 B.n1073 B.n1072 10.6151
R2826 B.n1074 B.n1073 10.6151
R2827 B.n1076 B.n1074 10.6151
R2828 B.n1077 B.n1076 10.6151
R2829 B.n1078 B.n1077 10.6151
R2830 B.n1079 B.n1078 10.6151
R2831 B.n1081 B.n1079 10.6151
R2832 B.n1082 B.n1081 10.6151
R2833 B.n1083 B.n1082 10.6151
R2834 B.n1084 B.n1083 10.6151
R2835 B.n1086 B.n1084 10.6151
R2836 B.n1087 B.n1086 10.6151
R2837 B.n1088 B.n1087 10.6151
R2838 B.n1089 B.n1088 10.6151
R2839 B.n1091 B.n1089 10.6151
R2840 B.n1092 B.n1091 10.6151
R2841 B.n1093 B.n1092 10.6151
R2842 B.n1094 B.n1093 10.6151
R2843 B.n1096 B.n1094 10.6151
R2844 B.n1097 B.n1096 10.6151
R2845 B.n1098 B.n1097 10.6151
R2846 B.n1099 B.n1098 10.6151
R2847 B.n1101 B.n1099 10.6151
R2848 B.n1102 B.n1101 10.6151
R2849 B.n1103 B.n1102 10.6151
R2850 B.n1104 B.n1103 10.6151
R2851 B.n1106 B.n1104 10.6151
R2852 B.n1107 B.n1106 10.6151
R2853 B.n1108 B.n1107 10.6151
R2854 B.n1269 B.n1 10.6151
R2855 B.n1269 B.n1268 10.6151
R2856 B.n1268 B.n1267 10.6151
R2857 B.n1267 B.n10 10.6151
R2858 B.n1261 B.n10 10.6151
R2859 B.n1261 B.n1260 10.6151
R2860 B.n1260 B.n1259 10.6151
R2861 B.n1259 B.n18 10.6151
R2862 B.n1253 B.n18 10.6151
R2863 B.n1253 B.n1252 10.6151
R2864 B.n1252 B.n1251 10.6151
R2865 B.n1251 B.n25 10.6151
R2866 B.n1245 B.n25 10.6151
R2867 B.n1245 B.n1244 10.6151
R2868 B.n1244 B.n1243 10.6151
R2869 B.n1243 B.n32 10.6151
R2870 B.n1237 B.n32 10.6151
R2871 B.n1237 B.n1236 10.6151
R2872 B.n1236 B.n1235 10.6151
R2873 B.n1235 B.n39 10.6151
R2874 B.n1229 B.n39 10.6151
R2875 B.n1229 B.n1228 10.6151
R2876 B.n1228 B.n1227 10.6151
R2877 B.n1227 B.n46 10.6151
R2878 B.n1221 B.n46 10.6151
R2879 B.n1221 B.n1220 10.6151
R2880 B.n1220 B.n1219 10.6151
R2881 B.n1219 B.n53 10.6151
R2882 B.n1213 B.n53 10.6151
R2883 B.n1213 B.n1212 10.6151
R2884 B.n1212 B.n1211 10.6151
R2885 B.n1211 B.n60 10.6151
R2886 B.n1205 B.n60 10.6151
R2887 B.n1205 B.n1204 10.6151
R2888 B.n1204 B.n1203 10.6151
R2889 B.n1203 B.n67 10.6151
R2890 B.n1197 B.n67 10.6151
R2891 B.n1197 B.n1196 10.6151
R2892 B.n1196 B.n1195 10.6151
R2893 B.n1195 B.n74 10.6151
R2894 B.n1189 B.n74 10.6151
R2895 B.n1189 B.n1188 10.6151
R2896 B.n1188 B.n1187 10.6151
R2897 B.n1187 B.n81 10.6151
R2898 B.n1181 B.n81 10.6151
R2899 B.n1181 B.n1180 10.6151
R2900 B.n1180 B.n1179 10.6151
R2901 B.n1179 B.n88 10.6151
R2902 B.n1173 B.n88 10.6151
R2903 B.n1173 B.n1172 10.6151
R2904 B.n1172 B.n1171 10.6151
R2905 B.n1171 B.n95 10.6151
R2906 B.n1165 B.n95 10.6151
R2907 B.n1165 B.n1164 10.6151
R2908 B.n1164 B.n1163 10.6151
R2909 B.n1163 B.n102 10.6151
R2910 B.n1157 B.n102 10.6151
R2911 B.n1157 B.n1156 10.6151
R2912 B.n1156 B.n1155 10.6151
R2913 B.n1155 B.n109 10.6151
R2914 B.n1149 B.n109 10.6151
R2915 B.n1149 B.n1148 10.6151
R2916 B.n1148 B.n1147 10.6151
R2917 B.n1147 B.n116 10.6151
R2918 B.n1141 B.n116 10.6151
R2919 B.n1141 B.n1140 10.6151
R2920 B.n1140 B.n1139 10.6151
R2921 B.n1139 B.n123 10.6151
R2922 B.n1133 B.n123 10.6151
R2923 B.n1133 B.n1132 10.6151
R2924 B.n1132 B.n1131 10.6151
R2925 B.n1131 B.n130 10.6151
R2926 B.n1125 B.n130 10.6151
R2927 B.n1125 B.n1124 10.6151
R2928 B.n1124 B.n1123 10.6151
R2929 B.n1123 B.n137 10.6151
R2930 B.n1117 B.n137 10.6151
R2931 B.n1117 B.n1116 10.6151
R2932 B.n1116 B.n1115 10.6151
R2933 B.n1115 B.n144 10.6151
R2934 B.n200 B.n199 10.6151
R2935 B.n203 B.n200 10.6151
R2936 B.n204 B.n203 10.6151
R2937 B.n207 B.n204 10.6151
R2938 B.n208 B.n207 10.6151
R2939 B.n211 B.n208 10.6151
R2940 B.n212 B.n211 10.6151
R2941 B.n215 B.n212 10.6151
R2942 B.n216 B.n215 10.6151
R2943 B.n219 B.n216 10.6151
R2944 B.n220 B.n219 10.6151
R2945 B.n223 B.n220 10.6151
R2946 B.n224 B.n223 10.6151
R2947 B.n227 B.n224 10.6151
R2948 B.n228 B.n227 10.6151
R2949 B.n231 B.n228 10.6151
R2950 B.n232 B.n231 10.6151
R2951 B.n235 B.n232 10.6151
R2952 B.n236 B.n235 10.6151
R2953 B.n239 B.n236 10.6151
R2954 B.n240 B.n239 10.6151
R2955 B.n243 B.n240 10.6151
R2956 B.n244 B.n243 10.6151
R2957 B.n247 B.n244 10.6151
R2958 B.n248 B.n247 10.6151
R2959 B.n251 B.n248 10.6151
R2960 B.n252 B.n251 10.6151
R2961 B.n255 B.n252 10.6151
R2962 B.n256 B.n255 10.6151
R2963 B.n259 B.n256 10.6151
R2964 B.n260 B.n259 10.6151
R2965 B.n263 B.n260 10.6151
R2966 B.n264 B.n263 10.6151
R2967 B.n267 B.n264 10.6151
R2968 B.n268 B.n267 10.6151
R2969 B.n271 B.n268 10.6151
R2970 B.n272 B.n271 10.6151
R2971 B.n275 B.n272 10.6151
R2972 B.n276 B.n275 10.6151
R2973 B.n280 B.n279 10.6151
R2974 B.n283 B.n280 10.6151
R2975 B.n284 B.n283 10.6151
R2976 B.n287 B.n284 10.6151
R2977 B.n288 B.n287 10.6151
R2978 B.n291 B.n288 10.6151
R2979 B.n292 B.n291 10.6151
R2980 B.n295 B.n292 10.6151
R2981 B.n300 B.n297 10.6151
R2982 B.n301 B.n300 10.6151
R2983 B.n304 B.n301 10.6151
R2984 B.n305 B.n304 10.6151
R2985 B.n308 B.n305 10.6151
R2986 B.n309 B.n308 10.6151
R2987 B.n312 B.n309 10.6151
R2988 B.n313 B.n312 10.6151
R2989 B.n316 B.n313 10.6151
R2990 B.n317 B.n316 10.6151
R2991 B.n320 B.n317 10.6151
R2992 B.n321 B.n320 10.6151
R2993 B.n324 B.n321 10.6151
R2994 B.n325 B.n324 10.6151
R2995 B.n328 B.n325 10.6151
R2996 B.n329 B.n328 10.6151
R2997 B.n332 B.n329 10.6151
R2998 B.n333 B.n332 10.6151
R2999 B.n336 B.n333 10.6151
R3000 B.n337 B.n336 10.6151
R3001 B.n340 B.n337 10.6151
R3002 B.n341 B.n340 10.6151
R3003 B.n344 B.n341 10.6151
R3004 B.n345 B.n344 10.6151
R3005 B.n348 B.n345 10.6151
R3006 B.n349 B.n348 10.6151
R3007 B.n352 B.n349 10.6151
R3008 B.n353 B.n352 10.6151
R3009 B.n356 B.n353 10.6151
R3010 B.n357 B.n356 10.6151
R3011 B.n360 B.n357 10.6151
R3012 B.n361 B.n360 10.6151
R3013 B.n364 B.n361 10.6151
R3014 B.n365 B.n364 10.6151
R3015 B.n368 B.n365 10.6151
R3016 B.n369 B.n368 10.6151
R3017 B.n372 B.n369 10.6151
R3018 B.n373 B.n372 10.6151
R3019 B.n1109 B.n373 10.6151
R3020 B.n790 B.t15 10.6061
R3021 B.n910 B.t0 10.6061
R3022 B.t3 B.n384 10.6061
R3023 B.t8 B.n16 10.6061
R3024 B.n1209 B.t4 10.6061
R3025 B.n1129 B.t11 10.6061
R3026 B.n1277 B.n0 8.11757
R3027 B.n1277 B.n1 8.11757
R3028 B.n679 B.n678 6.5566
R3029 B.n662 B.n584 6.5566
R3030 B.n279 B.n197 6.5566
R3031 B.n296 B.n295 6.5566
R3032 B.n680 B.n679 4.05904
R3033 B.n659 B.n584 4.05904
R3034 B.n276 B.n197 4.05904
R3035 B.n297 B.n296 4.05904
R3036 B.n874 B.t7 1.3262
R3037 B.n1185 B.t6 1.3262
R3038 VN.n110 VN.n109 161.3
R3039 VN.n108 VN.n57 161.3
R3040 VN.n107 VN.n106 161.3
R3041 VN.n105 VN.n58 161.3
R3042 VN.n104 VN.n103 161.3
R3043 VN.n102 VN.n59 161.3
R3044 VN.n101 VN.n100 161.3
R3045 VN.n99 VN.n60 161.3
R3046 VN.n98 VN.n97 161.3
R3047 VN.n95 VN.n61 161.3
R3048 VN.n94 VN.n93 161.3
R3049 VN.n92 VN.n62 161.3
R3050 VN.n91 VN.n90 161.3
R3051 VN.n89 VN.n63 161.3
R3052 VN.n88 VN.n87 161.3
R3053 VN.n86 VN.n64 161.3
R3054 VN.n85 VN.n84 161.3
R3055 VN.n82 VN.n65 161.3
R3056 VN.n81 VN.n80 161.3
R3057 VN.n79 VN.n66 161.3
R3058 VN.n78 VN.n77 161.3
R3059 VN.n76 VN.n67 161.3
R3060 VN.n75 VN.n74 161.3
R3061 VN.n73 VN.n68 161.3
R3062 VN.n72 VN.n71 161.3
R3063 VN.n54 VN.n53 161.3
R3064 VN.n52 VN.n1 161.3
R3065 VN.n51 VN.n50 161.3
R3066 VN.n49 VN.n2 161.3
R3067 VN.n48 VN.n47 161.3
R3068 VN.n46 VN.n3 161.3
R3069 VN.n45 VN.n44 161.3
R3070 VN.n43 VN.n4 161.3
R3071 VN.n42 VN.n41 161.3
R3072 VN.n39 VN.n5 161.3
R3073 VN.n38 VN.n37 161.3
R3074 VN.n36 VN.n6 161.3
R3075 VN.n35 VN.n34 161.3
R3076 VN.n33 VN.n7 161.3
R3077 VN.n32 VN.n31 161.3
R3078 VN.n30 VN.n8 161.3
R3079 VN.n29 VN.n28 161.3
R3080 VN.n26 VN.n9 161.3
R3081 VN.n25 VN.n24 161.3
R3082 VN.n23 VN.n10 161.3
R3083 VN.n22 VN.n21 161.3
R3084 VN.n20 VN.n11 161.3
R3085 VN.n19 VN.n18 161.3
R3086 VN.n17 VN.n12 161.3
R3087 VN.n16 VN.n15 161.3
R3088 VN.n69 VN.t7 104.216
R3089 VN.n13 VN.t3 104.216
R3090 VN.n55 VN.n0 85.5092
R3091 VN.n111 VN.n56 85.5092
R3092 VN.n14 VN.t4 71.0453
R3093 VN.n27 VN.t6 71.0453
R3094 VN.n40 VN.t9 71.0453
R3095 VN.n0 VN.t1 71.0453
R3096 VN.n70 VN.t2 71.0453
R3097 VN.n83 VN.t0 71.0453
R3098 VN.n96 VN.t5 71.0453
R3099 VN.n56 VN.t8 71.0453
R3100 VN VN.n111 59.5926
R3101 VN.n21 VN.n20 56.4773
R3102 VN.n34 VN.n33 56.4773
R3103 VN.n77 VN.n76 56.4773
R3104 VN.n90 VN.n89 56.4773
R3105 VN.n70 VN.n69 54.3527
R3106 VN.n14 VN.n13 54.3527
R3107 VN.n47 VN.n2 40.8975
R3108 VN.n103 VN.n58 40.8975
R3109 VN.n47 VN.n46 39.9237
R3110 VN.n103 VN.n102 39.9237
R3111 VN.n15 VN.n12 24.3439
R3112 VN.n19 VN.n12 24.3439
R3113 VN.n20 VN.n19 24.3439
R3114 VN.n21 VN.n10 24.3439
R3115 VN.n25 VN.n10 24.3439
R3116 VN.n26 VN.n25 24.3439
R3117 VN.n28 VN.n8 24.3439
R3118 VN.n32 VN.n8 24.3439
R3119 VN.n33 VN.n32 24.3439
R3120 VN.n34 VN.n6 24.3439
R3121 VN.n38 VN.n6 24.3439
R3122 VN.n39 VN.n38 24.3439
R3123 VN.n41 VN.n4 24.3439
R3124 VN.n45 VN.n4 24.3439
R3125 VN.n46 VN.n45 24.3439
R3126 VN.n51 VN.n2 24.3439
R3127 VN.n52 VN.n51 24.3439
R3128 VN.n53 VN.n52 24.3439
R3129 VN.n76 VN.n75 24.3439
R3130 VN.n75 VN.n68 24.3439
R3131 VN.n71 VN.n68 24.3439
R3132 VN.n89 VN.n88 24.3439
R3133 VN.n88 VN.n64 24.3439
R3134 VN.n84 VN.n64 24.3439
R3135 VN.n82 VN.n81 24.3439
R3136 VN.n81 VN.n66 24.3439
R3137 VN.n77 VN.n66 24.3439
R3138 VN.n102 VN.n101 24.3439
R3139 VN.n101 VN.n60 24.3439
R3140 VN.n97 VN.n60 24.3439
R3141 VN.n95 VN.n94 24.3439
R3142 VN.n94 VN.n62 24.3439
R3143 VN.n90 VN.n62 24.3439
R3144 VN.n109 VN.n108 24.3439
R3145 VN.n108 VN.n107 24.3439
R3146 VN.n107 VN.n58 24.3439
R3147 VN.n15 VN.n14 20.449
R3148 VN.n40 VN.n39 20.449
R3149 VN.n71 VN.n70 20.449
R3150 VN.n96 VN.n95 20.449
R3151 VN.n27 VN.n26 12.1722
R3152 VN.n28 VN.n27 12.1722
R3153 VN.n84 VN.n83 12.1722
R3154 VN.n83 VN.n82 12.1722
R3155 VN.n53 VN.n0 4.38232
R3156 VN.n109 VN.n56 4.38232
R3157 VN.n41 VN.n40 3.89545
R3158 VN.n97 VN.n96 3.89545
R3159 VN.n72 VN.n69 2.44072
R3160 VN.n16 VN.n13 2.44072
R3161 VN.n111 VN.n110 0.355081
R3162 VN.n55 VN.n54 0.355081
R3163 VN VN.n55 0.26685
R3164 VN.n110 VN.n57 0.189894
R3165 VN.n106 VN.n57 0.189894
R3166 VN.n106 VN.n105 0.189894
R3167 VN.n105 VN.n104 0.189894
R3168 VN.n104 VN.n59 0.189894
R3169 VN.n100 VN.n59 0.189894
R3170 VN.n100 VN.n99 0.189894
R3171 VN.n99 VN.n98 0.189894
R3172 VN.n98 VN.n61 0.189894
R3173 VN.n93 VN.n61 0.189894
R3174 VN.n93 VN.n92 0.189894
R3175 VN.n92 VN.n91 0.189894
R3176 VN.n91 VN.n63 0.189894
R3177 VN.n87 VN.n63 0.189894
R3178 VN.n87 VN.n86 0.189894
R3179 VN.n86 VN.n85 0.189894
R3180 VN.n85 VN.n65 0.189894
R3181 VN.n80 VN.n65 0.189894
R3182 VN.n80 VN.n79 0.189894
R3183 VN.n79 VN.n78 0.189894
R3184 VN.n78 VN.n67 0.189894
R3185 VN.n74 VN.n67 0.189894
R3186 VN.n74 VN.n73 0.189894
R3187 VN.n73 VN.n72 0.189894
R3188 VN.n17 VN.n16 0.189894
R3189 VN.n18 VN.n17 0.189894
R3190 VN.n18 VN.n11 0.189894
R3191 VN.n22 VN.n11 0.189894
R3192 VN.n23 VN.n22 0.189894
R3193 VN.n24 VN.n23 0.189894
R3194 VN.n24 VN.n9 0.189894
R3195 VN.n29 VN.n9 0.189894
R3196 VN.n30 VN.n29 0.189894
R3197 VN.n31 VN.n30 0.189894
R3198 VN.n31 VN.n7 0.189894
R3199 VN.n35 VN.n7 0.189894
R3200 VN.n36 VN.n35 0.189894
R3201 VN.n37 VN.n36 0.189894
R3202 VN.n37 VN.n5 0.189894
R3203 VN.n42 VN.n5 0.189894
R3204 VN.n43 VN.n42 0.189894
R3205 VN.n44 VN.n43 0.189894
R3206 VN.n44 VN.n3 0.189894
R3207 VN.n48 VN.n3 0.189894
R3208 VN.n49 VN.n48 0.189894
R3209 VN.n50 VN.n49 0.189894
R3210 VN.n50 VN.n1 0.189894
R3211 VN.n54 VN.n1 0.189894
R3212 VDD2.n121 VDD2.n65 289.615
R3213 VDD2.n56 VDD2.n0 289.615
R3214 VDD2.n122 VDD2.n121 185
R3215 VDD2.n120 VDD2.n119 185
R3216 VDD2.n69 VDD2.n68 185
R3217 VDD2.n114 VDD2.n113 185
R3218 VDD2.n112 VDD2.n111 185
R3219 VDD2.n73 VDD2.n72 185
R3220 VDD2.n77 VDD2.n75 185
R3221 VDD2.n106 VDD2.n105 185
R3222 VDD2.n104 VDD2.n103 185
R3223 VDD2.n79 VDD2.n78 185
R3224 VDD2.n98 VDD2.n97 185
R3225 VDD2.n96 VDD2.n95 185
R3226 VDD2.n83 VDD2.n82 185
R3227 VDD2.n90 VDD2.n89 185
R3228 VDD2.n88 VDD2.n87 185
R3229 VDD2.n21 VDD2.n20 185
R3230 VDD2.n23 VDD2.n22 185
R3231 VDD2.n16 VDD2.n15 185
R3232 VDD2.n29 VDD2.n28 185
R3233 VDD2.n31 VDD2.n30 185
R3234 VDD2.n12 VDD2.n11 185
R3235 VDD2.n38 VDD2.n37 185
R3236 VDD2.n39 VDD2.n10 185
R3237 VDD2.n41 VDD2.n40 185
R3238 VDD2.n8 VDD2.n7 185
R3239 VDD2.n47 VDD2.n46 185
R3240 VDD2.n49 VDD2.n48 185
R3241 VDD2.n4 VDD2.n3 185
R3242 VDD2.n55 VDD2.n54 185
R3243 VDD2.n57 VDD2.n56 185
R3244 VDD2.n86 VDD2.t1 149.524
R3245 VDD2.n19 VDD2.t6 149.524
R3246 VDD2.n121 VDD2.n120 104.615
R3247 VDD2.n120 VDD2.n68 104.615
R3248 VDD2.n113 VDD2.n68 104.615
R3249 VDD2.n113 VDD2.n112 104.615
R3250 VDD2.n112 VDD2.n72 104.615
R3251 VDD2.n77 VDD2.n72 104.615
R3252 VDD2.n105 VDD2.n77 104.615
R3253 VDD2.n105 VDD2.n104 104.615
R3254 VDD2.n104 VDD2.n78 104.615
R3255 VDD2.n97 VDD2.n78 104.615
R3256 VDD2.n97 VDD2.n96 104.615
R3257 VDD2.n96 VDD2.n82 104.615
R3258 VDD2.n89 VDD2.n82 104.615
R3259 VDD2.n89 VDD2.n88 104.615
R3260 VDD2.n22 VDD2.n21 104.615
R3261 VDD2.n22 VDD2.n15 104.615
R3262 VDD2.n29 VDD2.n15 104.615
R3263 VDD2.n30 VDD2.n29 104.615
R3264 VDD2.n30 VDD2.n11 104.615
R3265 VDD2.n38 VDD2.n11 104.615
R3266 VDD2.n39 VDD2.n38 104.615
R3267 VDD2.n40 VDD2.n39 104.615
R3268 VDD2.n40 VDD2.n7 104.615
R3269 VDD2.n47 VDD2.n7 104.615
R3270 VDD2.n48 VDD2.n47 104.615
R3271 VDD2.n48 VDD2.n3 104.615
R3272 VDD2.n55 VDD2.n3 104.615
R3273 VDD2.n56 VDD2.n55 104.615
R3274 VDD2.n64 VDD2.n63 63.179
R3275 VDD2 VDD2.n129 63.1761
R3276 VDD2.n128 VDD2.n127 60.5384
R3277 VDD2.n62 VDD2.n61 60.5382
R3278 VDD2.n88 VDD2.t1 52.3082
R3279 VDD2.n21 VDD2.t6 52.3082
R3280 VDD2.n62 VDD2.n60 50.9074
R3281 VDD2.n126 VDD2.n64 50.5493
R3282 VDD2.n126 VDD2.n125 47.3126
R3283 VDD2.n75 VDD2.n73 13.1884
R3284 VDD2.n41 VDD2.n8 13.1884
R3285 VDD2.n111 VDD2.n110 12.8005
R3286 VDD2.n107 VDD2.n106 12.8005
R3287 VDD2.n42 VDD2.n10 12.8005
R3288 VDD2.n46 VDD2.n45 12.8005
R3289 VDD2.n114 VDD2.n71 12.0247
R3290 VDD2.n103 VDD2.n76 12.0247
R3291 VDD2.n37 VDD2.n36 12.0247
R3292 VDD2.n49 VDD2.n6 12.0247
R3293 VDD2.n115 VDD2.n69 11.249
R3294 VDD2.n102 VDD2.n79 11.249
R3295 VDD2.n35 VDD2.n12 11.249
R3296 VDD2.n50 VDD2.n4 11.249
R3297 VDD2.n119 VDD2.n118 10.4732
R3298 VDD2.n99 VDD2.n98 10.4732
R3299 VDD2.n32 VDD2.n31 10.4732
R3300 VDD2.n54 VDD2.n53 10.4732
R3301 VDD2.n87 VDD2.n86 10.2747
R3302 VDD2.n20 VDD2.n19 10.2747
R3303 VDD2.n122 VDD2.n67 9.69747
R3304 VDD2.n95 VDD2.n81 9.69747
R3305 VDD2.n28 VDD2.n14 9.69747
R3306 VDD2.n57 VDD2.n2 9.69747
R3307 VDD2.n125 VDD2.n124 9.45567
R3308 VDD2.n60 VDD2.n59 9.45567
R3309 VDD2.n85 VDD2.n84 9.3005
R3310 VDD2.n92 VDD2.n91 9.3005
R3311 VDD2.n94 VDD2.n93 9.3005
R3312 VDD2.n81 VDD2.n80 9.3005
R3313 VDD2.n100 VDD2.n99 9.3005
R3314 VDD2.n102 VDD2.n101 9.3005
R3315 VDD2.n76 VDD2.n74 9.3005
R3316 VDD2.n108 VDD2.n107 9.3005
R3317 VDD2.n124 VDD2.n123 9.3005
R3318 VDD2.n67 VDD2.n66 9.3005
R3319 VDD2.n118 VDD2.n117 9.3005
R3320 VDD2.n116 VDD2.n115 9.3005
R3321 VDD2.n71 VDD2.n70 9.3005
R3322 VDD2.n110 VDD2.n109 9.3005
R3323 VDD2.n59 VDD2.n58 9.3005
R3324 VDD2.n2 VDD2.n1 9.3005
R3325 VDD2.n53 VDD2.n52 9.3005
R3326 VDD2.n51 VDD2.n50 9.3005
R3327 VDD2.n6 VDD2.n5 9.3005
R3328 VDD2.n45 VDD2.n44 9.3005
R3329 VDD2.n18 VDD2.n17 9.3005
R3330 VDD2.n25 VDD2.n24 9.3005
R3331 VDD2.n27 VDD2.n26 9.3005
R3332 VDD2.n14 VDD2.n13 9.3005
R3333 VDD2.n33 VDD2.n32 9.3005
R3334 VDD2.n35 VDD2.n34 9.3005
R3335 VDD2.n36 VDD2.n9 9.3005
R3336 VDD2.n43 VDD2.n42 9.3005
R3337 VDD2.n123 VDD2.n65 8.92171
R3338 VDD2.n94 VDD2.n83 8.92171
R3339 VDD2.n27 VDD2.n16 8.92171
R3340 VDD2.n58 VDD2.n0 8.92171
R3341 VDD2.n91 VDD2.n90 8.14595
R3342 VDD2.n24 VDD2.n23 8.14595
R3343 VDD2.n87 VDD2.n85 7.3702
R3344 VDD2.n20 VDD2.n18 7.3702
R3345 VDD2.n90 VDD2.n85 5.81868
R3346 VDD2.n23 VDD2.n18 5.81868
R3347 VDD2.n125 VDD2.n65 5.04292
R3348 VDD2.n91 VDD2.n83 5.04292
R3349 VDD2.n24 VDD2.n16 5.04292
R3350 VDD2.n60 VDD2.n0 5.04292
R3351 VDD2.n123 VDD2.n122 4.26717
R3352 VDD2.n95 VDD2.n94 4.26717
R3353 VDD2.n28 VDD2.n27 4.26717
R3354 VDD2.n58 VDD2.n57 4.26717
R3355 VDD2.n128 VDD2.n126 3.59533
R3356 VDD2.n119 VDD2.n67 3.49141
R3357 VDD2.n98 VDD2.n81 3.49141
R3358 VDD2.n31 VDD2.n14 3.49141
R3359 VDD2.n54 VDD2.n2 3.49141
R3360 VDD2.n86 VDD2.n84 2.84303
R3361 VDD2.n19 VDD2.n17 2.84303
R3362 VDD2.n118 VDD2.n69 2.71565
R3363 VDD2.n99 VDD2.n79 2.71565
R3364 VDD2.n32 VDD2.n12 2.71565
R3365 VDD2.n53 VDD2.n4 2.71565
R3366 VDD2.n115 VDD2.n114 1.93989
R3367 VDD2.n103 VDD2.n102 1.93989
R3368 VDD2.n37 VDD2.n35 1.93989
R3369 VDD2.n50 VDD2.n49 1.93989
R3370 VDD2.n129 VDD2.t7 1.74962
R3371 VDD2.n129 VDD2.t2 1.74962
R3372 VDD2.n127 VDD2.t4 1.74962
R3373 VDD2.n127 VDD2.t9 1.74962
R3374 VDD2.n63 VDD2.t0 1.74962
R3375 VDD2.n63 VDD2.t8 1.74962
R3376 VDD2.n61 VDD2.t5 1.74962
R3377 VDD2.n61 VDD2.t3 1.74962
R3378 VDD2.n111 VDD2.n71 1.16414
R3379 VDD2.n106 VDD2.n76 1.16414
R3380 VDD2.n36 VDD2.n10 1.16414
R3381 VDD2.n46 VDD2.n6 1.16414
R3382 VDD2 VDD2.n128 0.957397
R3383 VDD2.n64 VDD2.n62 0.843861
R3384 VDD2.n110 VDD2.n73 0.388379
R3385 VDD2.n107 VDD2.n75 0.388379
R3386 VDD2.n42 VDD2.n41 0.388379
R3387 VDD2.n45 VDD2.n8 0.388379
R3388 VDD2.n124 VDD2.n66 0.155672
R3389 VDD2.n117 VDD2.n66 0.155672
R3390 VDD2.n117 VDD2.n116 0.155672
R3391 VDD2.n116 VDD2.n70 0.155672
R3392 VDD2.n109 VDD2.n70 0.155672
R3393 VDD2.n109 VDD2.n108 0.155672
R3394 VDD2.n108 VDD2.n74 0.155672
R3395 VDD2.n101 VDD2.n74 0.155672
R3396 VDD2.n101 VDD2.n100 0.155672
R3397 VDD2.n100 VDD2.n80 0.155672
R3398 VDD2.n93 VDD2.n80 0.155672
R3399 VDD2.n93 VDD2.n92 0.155672
R3400 VDD2.n92 VDD2.n84 0.155672
R3401 VDD2.n25 VDD2.n17 0.155672
R3402 VDD2.n26 VDD2.n25 0.155672
R3403 VDD2.n26 VDD2.n13 0.155672
R3404 VDD2.n33 VDD2.n13 0.155672
R3405 VDD2.n34 VDD2.n33 0.155672
R3406 VDD2.n34 VDD2.n9 0.155672
R3407 VDD2.n43 VDD2.n9 0.155672
R3408 VDD2.n44 VDD2.n43 0.155672
R3409 VDD2.n44 VDD2.n5 0.155672
R3410 VDD2.n51 VDD2.n5 0.155672
R3411 VDD2.n52 VDD2.n51 0.155672
R3412 VDD2.n52 VDD2.n1 0.155672
R3413 VDD2.n59 VDD2.n1 0.155672
C0 VDD2 VTAIL 10.8394f
C1 VTAIL VDD1 10.779099f
C2 VDD2 VDD1 2.98143f
C3 VP VTAIL 11.9982f
C4 VP VDD2 0.740775f
C5 VP VDD1 11.3592f
C6 VN VTAIL 11.9834f
C7 VN VDD2 10.7775f
C8 VN VDD1 0.155742f
C9 VP VN 10.1092f
C10 VDD2 B 8.552464f
C11 VDD1 B 8.520507f
C12 VTAIL B 8.857284f
C13 VN B 24.029488f
C14 VP B 22.619402f
C15 VDD2.n0 B 0.033117f
C16 VDD2.n1 B 0.025001f
C17 VDD2.n2 B 0.013434f
C18 VDD2.n3 B 0.031754f
C19 VDD2.n4 B 0.014225f
C20 VDD2.n5 B 0.025001f
C21 VDD2.n6 B 0.013434f
C22 VDD2.n7 B 0.031754f
C23 VDD2.n8 B 0.01383f
C24 VDD2.n9 B 0.025001f
C25 VDD2.n10 B 0.014225f
C26 VDD2.n11 B 0.031754f
C27 VDD2.n12 B 0.014225f
C28 VDD2.n13 B 0.025001f
C29 VDD2.n14 B 0.013434f
C30 VDD2.n15 B 0.031754f
C31 VDD2.n16 B 0.014225f
C32 VDD2.n17 B 1.18563f
C33 VDD2.n18 B 0.013434f
C34 VDD2.t6 B 0.053539f
C35 VDD2.n19 B 0.173726f
C36 VDD2.n20 B 0.022448f
C37 VDD2.n21 B 0.023815f
C38 VDD2.n22 B 0.031754f
C39 VDD2.n23 B 0.014225f
C40 VDD2.n24 B 0.013434f
C41 VDD2.n25 B 0.025001f
C42 VDD2.n26 B 0.025001f
C43 VDD2.n27 B 0.013434f
C44 VDD2.n28 B 0.014225f
C45 VDD2.n29 B 0.031754f
C46 VDD2.n30 B 0.031754f
C47 VDD2.n31 B 0.014225f
C48 VDD2.n32 B 0.013434f
C49 VDD2.n33 B 0.025001f
C50 VDD2.n34 B 0.025001f
C51 VDD2.n35 B 0.013434f
C52 VDD2.n36 B 0.013434f
C53 VDD2.n37 B 0.014225f
C54 VDD2.n38 B 0.031754f
C55 VDD2.n39 B 0.031754f
C56 VDD2.n40 B 0.031754f
C57 VDD2.n41 B 0.01383f
C58 VDD2.n42 B 0.013434f
C59 VDD2.n43 B 0.025001f
C60 VDD2.n44 B 0.025001f
C61 VDD2.n45 B 0.013434f
C62 VDD2.n46 B 0.014225f
C63 VDD2.n47 B 0.031754f
C64 VDD2.n48 B 0.031754f
C65 VDD2.n49 B 0.014225f
C66 VDD2.n50 B 0.013434f
C67 VDD2.n51 B 0.025001f
C68 VDD2.n52 B 0.025001f
C69 VDD2.n53 B 0.013434f
C70 VDD2.n54 B 0.014225f
C71 VDD2.n55 B 0.031754f
C72 VDD2.n56 B 0.065162f
C73 VDD2.n57 B 0.014225f
C74 VDD2.n58 B 0.013434f
C75 VDD2.n59 B 0.055056f
C76 VDD2.n60 B 0.077032f
C77 VDD2.t5 B 0.223642f
C78 VDD2.t3 B 0.223642f
C79 VDD2.n61 B 1.98381f
C80 VDD2.n62 B 0.878446f
C81 VDD2.t0 B 0.223642f
C82 VDD2.t8 B 0.223642f
C83 VDD2.n63 B 2.01392f
C84 VDD2.n64 B 3.50863f
C85 VDD2.n65 B 0.033117f
C86 VDD2.n66 B 0.025001f
C87 VDD2.n67 B 0.013434f
C88 VDD2.n68 B 0.031754f
C89 VDD2.n69 B 0.014225f
C90 VDD2.n70 B 0.025001f
C91 VDD2.n71 B 0.013434f
C92 VDD2.n72 B 0.031754f
C93 VDD2.n73 B 0.01383f
C94 VDD2.n74 B 0.025001f
C95 VDD2.n75 B 0.01383f
C96 VDD2.n76 B 0.013434f
C97 VDD2.n77 B 0.031754f
C98 VDD2.n78 B 0.031754f
C99 VDD2.n79 B 0.014225f
C100 VDD2.n80 B 0.025001f
C101 VDD2.n81 B 0.013434f
C102 VDD2.n82 B 0.031754f
C103 VDD2.n83 B 0.014225f
C104 VDD2.n84 B 1.18563f
C105 VDD2.n85 B 0.013434f
C106 VDD2.t1 B 0.053539f
C107 VDD2.n86 B 0.173726f
C108 VDD2.n87 B 0.022448f
C109 VDD2.n88 B 0.023815f
C110 VDD2.n89 B 0.031754f
C111 VDD2.n90 B 0.014225f
C112 VDD2.n91 B 0.013434f
C113 VDD2.n92 B 0.025001f
C114 VDD2.n93 B 0.025001f
C115 VDD2.n94 B 0.013434f
C116 VDD2.n95 B 0.014225f
C117 VDD2.n96 B 0.031754f
C118 VDD2.n97 B 0.031754f
C119 VDD2.n98 B 0.014225f
C120 VDD2.n99 B 0.013434f
C121 VDD2.n100 B 0.025001f
C122 VDD2.n101 B 0.025001f
C123 VDD2.n102 B 0.013434f
C124 VDD2.n103 B 0.014225f
C125 VDD2.n104 B 0.031754f
C126 VDD2.n105 B 0.031754f
C127 VDD2.n106 B 0.014225f
C128 VDD2.n107 B 0.013434f
C129 VDD2.n108 B 0.025001f
C130 VDD2.n109 B 0.025001f
C131 VDD2.n110 B 0.013434f
C132 VDD2.n111 B 0.014225f
C133 VDD2.n112 B 0.031754f
C134 VDD2.n113 B 0.031754f
C135 VDD2.n114 B 0.014225f
C136 VDD2.n115 B 0.013434f
C137 VDD2.n116 B 0.025001f
C138 VDD2.n117 B 0.025001f
C139 VDD2.n118 B 0.013434f
C140 VDD2.n119 B 0.014225f
C141 VDD2.n120 B 0.031754f
C142 VDD2.n121 B 0.065162f
C143 VDD2.n122 B 0.014225f
C144 VDD2.n123 B 0.013434f
C145 VDD2.n124 B 0.055056f
C146 VDD2.n125 B 0.053293f
C147 VDD2.n126 B 3.3206f
C148 VDD2.t4 B 0.223642f
C149 VDD2.t9 B 0.223642f
C150 VDD2.n127 B 1.98382f
C151 VDD2.n128 B 0.574466f
C152 VDD2.t7 B 0.223642f
C153 VDD2.t2 B 0.223642f
C154 VDD2.n129 B 2.01387f
C155 VN.t1 B 1.99034f
C156 VN.n0 B 0.764808f
C157 VN.n1 B 0.016834f
C158 VN.n2 B 0.033548f
C159 VN.n3 B 0.016834f
C160 VN.n4 B 0.031532f
C161 VN.n5 B 0.016834f
C162 VN.t9 B 1.99034f
C163 VN.n6 B 0.031532f
C164 VN.n7 B 0.016834f
C165 VN.n8 B 0.031532f
C166 VN.n9 B 0.016834f
C167 VN.t6 B 1.99034f
C168 VN.n10 B 0.031532f
C169 VN.n11 B 0.016834f
C170 VN.n12 B 0.031532f
C171 VN.t3 B 2.25625f
C172 VN.n13 B 0.725988f
C173 VN.t4 B 1.99034f
C174 VN.n14 B 0.765975f
C175 VN.n15 B 0.029041f
C176 VN.n16 B 0.216889f
C177 VN.n17 B 0.016834f
C178 VN.n18 B 0.016834f
C179 VN.n19 B 0.031532f
C180 VN.n20 B 0.020666f
C181 VN.n21 B 0.028697f
C182 VN.n22 B 0.016834f
C183 VN.n23 B 0.016834f
C184 VN.n24 B 0.016834f
C185 VN.n25 B 0.031532f
C186 VN.n26 B 0.023748f
C187 VN.n27 B 0.699145f
C188 VN.n28 B 0.023748f
C189 VN.n29 B 0.016834f
C190 VN.n30 B 0.016834f
C191 VN.n31 B 0.016834f
C192 VN.n32 B 0.031532f
C193 VN.n33 B 0.028697f
C194 VN.n34 B 0.020666f
C195 VN.n35 B 0.016834f
C196 VN.n36 B 0.016834f
C197 VN.n37 B 0.016834f
C198 VN.n38 B 0.031532f
C199 VN.n39 B 0.029041f
C200 VN.n40 B 0.699145f
C201 VN.n41 B 0.018454f
C202 VN.n42 B 0.016834f
C203 VN.n43 B 0.016834f
C204 VN.n44 B 0.016834f
C205 VN.n45 B 0.031532f
C206 VN.n46 B 0.033719f
C207 VN.n47 B 0.013628f
C208 VN.n48 B 0.016834f
C209 VN.n49 B 0.016834f
C210 VN.n50 B 0.016834f
C211 VN.n51 B 0.031532f
C212 VN.n52 B 0.031532f
C213 VN.n53 B 0.018766f
C214 VN.n54 B 0.027174f
C215 VN.n55 B 0.05137f
C216 VN.t8 B 1.99034f
C217 VN.n56 B 0.764808f
C218 VN.n57 B 0.016834f
C219 VN.n58 B 0.033548f
C220 VN.n59 B 0.016834f
C221 VN.n60 B 0.031532f
C222 VN.n61 B 0.016834f
C223 VN.t5 B 1.99034f
C224 VN.n62 B 0.031532f
C225 VN.n63 B 0.016834f
C226 VN.n64 B 0.031532f
C227 VN.n65 B 0.016834f
C228 VN.t0 B 1.99034f
C229 VN.n66 B 0.031532f
C230 VN.n67 B 0.016834f
C231 VN.n68 B 0.031532f
C232 VN.t7 B 2.25625f
C233 VN.n69 B 0.725988f
C234 VN.t2 B 1.99034f
C235 VN.n70 B 0.765975f
C236 VN.n71 B 0.029041f
C237 VN.n72 B 0.216889f
C238 VN.n73 B 0.016834f
C239 VN.n74 B 0.016834f
C240 VN.n75 B 0.031532f
C241 VN.n76 B 0.020666f
C242 VN.n77 B 0.028697f
C243 VN.n78 B 0.016834f
C244 VN.n79 B 0.016834f
C245 VN.n80 B 0.016834f
C246 VN.n81 B 0.031532f
C247 VN.n82 B 0.023748f
C248 VN.n83 B 0.699145f
C249 VN.n84 B 0.023748f
C250 VN.n85 B 0.016834f
C251 VN.n86 B 0.016834f
C252 VN.n87 B 0.016834f
C253 VN.n88 B 0.031532f
C254 VN.n89 B 0.028697f
C255 VN.n90 B 0.020666f
C256 VN.n91 B 0.016834f
C257 VN.n92 B 0.016834f
C258 VN.n93 B 0.016834f
C259 VN.n94 B 0.031532f
C260 VN.n95 B 0.029041f
C261 VN.n96 B 0.699145f
C262 VN.n97 B 0.018454f
C263 VN.n98 B 0.016834f
C264 VN.n99 B 0.016834f
C265 VN.n100 B 0.016834f
C266 VN.n101 B 0.031532f
C267 VN.n102 B 0.033719f
C268 VN.n103 B 0.013628f
C269 VN.n104 B 0.016834f
C270 VN.n105 B 0.016834f
C271 VN.n106 B 0.016834f
C272 VN.n107 B 0.031532f
C273 VN.n108 B 0.031532f
C274 VN.n109 B 0.018766f
C275 VN.n110 B 0.027174f
C276 VN.n111 B 1.23486f
C277 VTAIL.t8 B 0.234363f
C278 VTAIL.t2 B 0.234363f
C279 VTAIL.n0 B 1.99799f
C280 VTAIL.n1 B 0.686977f
C281 VTAIL.n2 B 0.034704f
C282 VTAIL.n3 B 0.026199f
C283 VTAIL.n4 B 0.014078f
C284 VTAIL.n5 B 0.033276f
C285 VTAIL.n6 B 0.014906f
C286 VTAIL.n7 B 0.026199f
C287 VTAIL.n8 B 0.014078f
C288 VTAIL.n9 B 0.033276f
C289 VTAIL.n10 B 0.014492f
C290 VTAIL.n11 B 0.026199f
C291 VTAIL.n12 B 0.014906f
C292 VTAIL.n13 B 0.033276f
C293 VTAIL.n14 B 0.014906f
C294 VTAIL.n15 B 0.026199f
C295 VTAIL.n16 B 0.014078f
C296 VTAIL.n17 B 0.033276f
C297 VTAIL.n18 B 0.014906f
C298 VTAIL.n19 B 1.24247f
C299 VTAIL.n20 B 0.014078f
C300 VTAIL.t17 B 0.056105f
C301 VTAIL.n21 B 0.182054f
C302 VTAIL.n22 B 0.023524f
C303 VTAIL.n23 B 0.024957f
C304 VTAIL.n24 B 0.033276f
C305 VTAIL.n25 B 0.014906f
C306 VTAIL.n26 B 0.014078f
C307 VTAIL.n27 B 0.026199f
C308 VTAIL.n28 B 0.026199f
C309 VTAIL.n29 B 0.014078f
C310 VTAIL.n30 B 0.014906f
C311 VTAIL.n31 B 0.033276f
C312 VTAIL.n32 B 0.033276f
C313 VTAIL.n33 B 0.014906f
C314 VTAIL.n34 B 0.014078f
C315 VTAIL.n35 B 0.026199f
C316 VTAIL.n36 B 0.026199f
C317 VTAIL.n37 B 0.014078f
C318 VTAIL.n38 B 0.014078f
C319 VTAIL.n39 B 0.014906f
C320 VTAIL.n40 B 0.033276f
C321 VTAIL.n41 B 0.033276f
C322 VTAIL.n42 B 0.033276f
C323 VTAIL.n43 B 0.014492f
C324 VTAIL.n44 B 0.014078f
C325 VTAIL.n45 B 0.026199f
C326 VTAIL.n46 B 0.026199f
C327 VTAIL.n47 B 0.014078f
C328 VTAIL.n48 B 0.014906f
C329 VTAIL.n49 B 0.033276f
C330 VTAIL.n50 B 0.033276f
C331 VTAIL.n51 B 0.014906f
C332 VTAIL.n52 B 0.014078f
C333 VTAIL.n53 B 0.026199f
C334 VTAIL.n54 B 0.026199f
C335 VTAIL.n55 B 0.014078f
C336 VTAIL.n56 B 0.014906f
C337 VTAIL.n57 B 0.033276f
C338 VTAIL.n58 B 0.068286f
C339 VTAIL.n59 B 0.014906f
C340 VTAIL.n60 B 0.014078f
C341 VTAIL.n61 B 0.057695f
C342 VTAIL.n62 B 0.037733f
C343 VTAIL.n63 B 0.515637f
C344 VTAIL.t11 B 0.234363f
C345 VTAIL.t13 B 0.234363f
C346 VTAIL.n64 B 1.99799f
C347 VTAIL.n65 B 0.870008f
C348 VTAIL.t16 B 0.234363f
C349 VTAIL.t9 B 0.234363f
C350 VTAIL.n66 B 1.99799f
C351 VTAIL.n67 B 2.35319f
C352 VTAIL.t1 B 0.234363f
C353 VTAIL.t7 B 0.234363f
C354 VTAIL.n68 B 1.99801f
C355 VTAIL.n69 B 2.35318f
C356 VTAIL.t0 B 0.234363f
C357 VTAIL.t19 B 0.234363f
C358 VTAIL.n70 B 1.99801f
C359 VTAIL.n71 B 0.869996f
C360 VTAIL.n72 B 0.034704f
C361 VTAIL.n73 B 0.026199f
C362 VTAIL.n74 B 0.014078f
C363 VTAIL.n75 B 0.033276f
C364 VTAIL.n76 B 0.014906f
C365 VTAIL.n77 B 0.026199f
C366 VTAIL.n78 B 0.014078f
C367 VTAIL.n79 B 0.033276f
C368 VTAIL.n80 B 0.014492f
C369 VTAIL.n81 B 0.026199f
C370 VTAIL.n82 B 0.014492f
C371 VTAIL.n83 B 0.014078f
C372 VTAIL.n84 B 0.033276f
C373 VTAIL.n85 B 0.033276f
C374 VTAIL.n86 B 0.014906f
C375 VTAIL.n87 B 0.026199f
C376 VTAIL.n88 B 0.014078f
C377 VTAIL.n89 B 0.033276f
C378 VTAIL.n90 B 0.014906f
C379 VTAIL.n91 B 1.24247f
C380 VTAIL.n92 B 0.014078f
C381 VTAIL.t3 B 0.056105f
C382 VTAIL.n93 B 0.182054f
C383 VTAIL.n94 B 0.023524f
C384 VTAIL.n95 B 0.024957f
C385 VTAIL.n96 B 0.033276f
C386 VTAIL.n97 B 0.014906f
C387 VTAIL.n98 B 0.014078f
C388 VTAIL.n99 B 0.026199f
C389 VTAIL.n100 B 0.026199f
C390 VTAIL.n101 B 0.014078f
C391 VTAIL.n102 B 0.014906f
C392 VTAIL.n103 B 0.033276f
C393 VTAIL.n104 B 0.033276f
C394 VTAIL.n105 B 0.014906f
C395 VTAIL.n106 B 0.014078f
C396 VTAIL.n107 B 0.026199f
C397 VTAIL.n108 B 0.026199f
C398 VTAIL.n109 B 0.014078f
C399 VTAIL.n110 B 0.014906f
C400 VTAIL.n111 B 0.033276f
C401 VTAIL.n112 B 0.033276f
C402 VTAIL.n113 B 0.014906f
C403 VTAIL.n114 B 0.014078f
C404 VTAIL.n115 B 0.026199f
C405 VTAIL.n116 B 0.026199f
C406 VTAIL.n117 B 0.014078f
C407 VTAIL.n118 B 0.014906f
C408 VTAIL.n119 B 0.033276f
C409 VTAIL.n120 B 0.033276f
C410 VTAIL.n121 B 0.014906f
C411 VTAIL.n122 B 0.014078f
C412 VTAIL.n123 B 0.026199f
C413 VTAIL.n124 B 0.026199f
C414 VTAIL.n125 B 0.014078f
C415 VTAIL.n126 B 0.014906f
C416 VTAIL.n127 B 0.033276f
C417 VTAIL.n128 B 0.068286f
C418 VTAIL.n129 B 0.014906f
C419 VTAIL.n130 B 0.014078f
C420 VTAIL.n131 B 0.057695f
C421 VTAIL.n132 B 0.037733f
C422 VTAIL.n133 B 0.515637f
C423 VTAIL.t12 B 0.234363f
C424 VTAIL.t18 B 0.234363f
C425 VTAIL.n134 B 1.99801f
C426 VTAIL.n135 B 0.757921f
C427 VTAIL.t14 B 0.234363f
C428 VTAIL.t10 B 0.234363f
C429 VTAIL.n136 B 1.99801f
C430 VTAIL.n137 B 0.869996f
C431 VTAIL.n138 B 0.034704f
C432 VTAIL.n139 B 0.026199f
C433 VTAIL.n140 B 0.014078f
C434 VTAIL.n141 B 0.033276f
C435 VTAIL.n142 B 0.014906f
C436 VTAIL.n143 B 0.026199f
C437 VTAIL.n144 B 0.014078f
C438 VTAIL.n145 B 0.033276f
C439 VTAIL.n146 B 0.014492f
C440 VTAIL.n147 B 0.026199f
C441 VTAIL.n148 B 0.014492f
C442 VTAIL.n149 B 0.014078f
C443 VTAIL.n150 B 0.033276f
C444 VTAIL.n151 B 0.033276f
C445 VTAIL.n152 B 0.014906f
C446 VTAIL.n153 B 0.026199f
C447 VTAIL.n154 B 0.014078f
C448 VTAIL.n155 B 0.033276f
C449 VTAIL.n156 B 0.014906f
C450 VTAIL.n157 B 1.24247f
C451 VTAIL.n158 B 0.014078f
C452 VTAIL.t15 B 0.056105f
C453 VTAIL.n159 B 0.182054f
C454 VTAIL.n160 B 0.023524f
C455 VTAIL.n161 B 0.024957f
C456 VTAIL.n162 B 0.033276f
C457 VTAIL.n163 B 0.014906f
C458 VTAIL.n164 B 0.014078f
C459 VTAIL.n165 B 0.026199f
C460 VTAIL.n166 B 0.026199f
C461 VTAIL.n167 B 0.014078f
C462 VTAIL.n168 B 0.014906f
C463 VTAIL.n169 B 0.033276f
C464 VTAIL.n170 B 0.033276f
C465 VTAIL.n171 B 0.014906f
C466 VTAIL.n172 B 0.014078f
C467 VTAIL.n173 B 0.026199f
C468 VTAIL.n174 B 0.026199f
C469 VTAIL.n175 B 0.014078f
C470 VTAIL.n176 B 0.014906f
C471 VTAIL.n177 B 0.033276f
C472 VTAIL.n178 B 0.033276f
C473 VTAIL.n179 B 0.014906f
C474 VTAIL.n180 B 0.014078f
C475 VTAIL.n181 B 0.026199f
C476 VTAIL.n182 B 0.026199f
C477 VTAIL.n183 B 0.014078f
C478 VTAIL.n184 B 0.014906f
C479 VTAIL.n185 B 0.033276f
C480 VTAIL.n186 B 0.033276f
C481 VTAIL.n187 B 0.014906f
C482 VTAIL.n188 B 0.014078f
C483 VTAIL.n189 B 0.026199f
C484 VTAIL.n190 B 0.026199f
C485 VTAIL.n191 B 0.014078f
C486 VTAIL.n192 B 0.014906f
C487 VTAIL.n193 B 0.033276f
C488 VTAIL.n194 B 0.068286f
C489 VTAIL.n195 B 0.014906f
C490 VTAIL.n196 B 0.014078f
C491 VTAIL.n197 B 0.057695f
C492 VTAIL.n198 B 0.037733f
C493 VTAIL.n199 B 1.80742f
C494 VTAIL.n200 B 0.034704f
C495 VTAIL.n201 B 0.026199f
C496 VTAIL.n202 B 0.014078f
C497 VTAIL.n203 B 0.033276f
C498 VTAIL.n204 B 0.014906f
C499 VTAIL.n205 B 0.026199f
C500 VTAIL.n206 B 0.014078f
C501 VTAIL.n207 B 0.033276f
C502 VTAIL.n208 B 0.014492f
C503 VTAIL.n209 B 0.026199f
C504 VTAIL.n210 B 0.014906f
C505 VTAIL.n211 B 0.033276f
C506 VTAIL.n212 B 0.014906f
C507 VTAIL.n213 B 0.026199f
C508 VTAIL.n214 B 0.014078f
C509 VTAIL.n215 B 0.033276f
C510 VTAIL.n216 B 0.014906f
C511 VTAIL.n217 B 1.24247f
C512 VTAIL.n218 B 0.014078f
C513 VTAIL.t5 B 0.056105f
C514 VTAIL.n219 B 0.182054f
C515 VTAIL.n220 B 0.023524f
C516 VTAIL.n221 B 0.024957f
C517 VTAIL.n222 B 0.033276f
C518 VTAIL.n223 B 0.014906f
C519 VTAIL.n224 B 0.014078f
C520 VTAIL.n225 B 0.026199f
C521 VTAIL.n226 B 0.026199f
C522 VTAIL.n227 B 0.014078f
C523 VTAIL.n228 B 0.014906f
C524 VTAIL.n229 B 0.033276f
C525 VTAIL.n230 B 0.033276f
C526 VTAIL.n231 B 0.014906f
C527 VTAIL.n232 B 0.014078f
C528 VTAIL.n233 B 0.026199f
C529 VTAIL.n234 B 0.026199f
C530 VTAIL.n235 B 0.014078f
C531 VTAIL.n236 B 0.014078f
C532 VTAIL.n237 B 0.014906f
C533 VTAIL.n238 B 0.033276f
C534 VTAIL.n239 B 0.033276f
C535 VTAIL.n240 B 0.033276f
C536 VTAIL.n241 B 0.014492f
C537 VTAIL.n242 B 0.014078f
C538 VTAIL.n243 B 0.026199f
C539 VTAIL.n244 B 0.026199f
C540 VTAIL.n245 B 0.014078f
C541 VTAIL.n246 B 0.014906f
C542 VTAIL.n247 B 0.033276f
C543 VTAIL.n248 B 0.033276f
C544 VTAIL.n249 B 0.014906f
C545 VTAIL.n250 B 0.014078f
C546 VTAIL.n251 B 0.026199f
C547 VTAIL.n252 B 0.026199f
C548 VTAIL.n253 B 0.014078f
C549 VTAIL.n254 B 0.014906f
C550 VTAIL.n255 B 0.033276f
C551 VTAIL.n256 B 0.068286f
C552 VTAIL.n257 B 0.014906f
C553 VTAIL.n258 B 0.014078f
C554 VTAIL.n259 B 0.057695f
C555 VTAIL.n260 B 0.037733f
C556 VTAIL.n261 B 1.80742f
C557 VTAIL.t4 B 0.234363f
C558 VTAIL.t6 B 0.234363f
C559 VTAIL.n262 B 1.99799f
C560 VTAIL.n263 B 0.637489f
C561 VDD1.n0 B 0.033798f
C562 VDD1.n1 B 0.025515f
C563 VDD1.n2 B 0.01371f
C564 VDD1.n3 B 0.032407f
C565 VDD1.n4 B 0.014517f
C566 VDD1.n5 B 0.025515f
C567 VDD1.n6 B 0.01371f
C568 VDD1.n7 B 0.032407f
C569 VDD1.n8 B 0.014114f
C570 VDD1.n9 B 0.025515f
C571 VDD1.n10 B 0.014114f
C572 VDD1.n11 B 0.01371f
C573 VDD1.n12 B 0.032407f
C574 VDD1.n13 B 0.032407f
C575 VDD1.n14 B 0.014517f
C576 VDD1.n15 B 0.025515f
C577 VDD1.n16 B 0.01371f
C578 VDD1.n17 B 0.032407f
C579 VDD1.n18 B 0.014517f
C580 VDD1.n19 B 1.21001f
C581 VDD1.n20 B 0.01371f
C582 VDD1.t7 B 0.05464f
C583 VDD1.n21 B 0.177298f
C584 VDD1.n22 B 0.022909f
C585 VDD1.n23 B 0.024305f
C586 VDD1.n24 B 0.032407f
C587 VDD1.n25 B 0.014517f
C588 VDD1.n26 B 0.01371f
C589 VDD1.n27 B 0.025515f
C590 VDD1.n28 B 0.025515f
C591 VDD1.n29 B 0.01371f
C592 VDD1.n30 B 0.014517f
C593 VDD1.n31 B 0.032407f
C594 VDD1.n32 B 0.032407f
C595 VDD1.n33 B 0.014517f
C596 VDD1.n34 B 0.01371f
C597 VDD1.n35 B 0.025515f
C598 VDD1.n36 B 0.025515f
C599 VDD1.n37 B 0.01371f
C600 VDD1.n38 B 0.014517f
C601 VDD1.n39 B 0.032407f
C602 VDD1.n40 B 0.032407f
C603 VDD1.n41 B 0.014517f
C604 VDD1.n42 B 0.01371f
C605 VDD1.n43 B 0.025515f
C606 VDD1.n44 B 0.025515f
C607 VDD1.n45 B 0.01371f
C608 VDD1.n46 B 0.014517f
C609 VDD1.n47 B 0.032407f
C610 VDD1.n48 B 0.032407f
C611 VDD1.n49 B 0.014517f
C612 VDD1.n50 B 0.01371f
C613 VDD1.n51 B 0.025515f
C614 VDD1.n52 B 0.025515f
C615 VDD1.n53 B 0.01371f
C616 VDD1.n54 B 0.014517f
C617 VDD1.n55 B 0.032407f
C618 VDD1.n56 B 0.066502f
C619 VDD1.n57 B 0.014517f
C620 VDD1.n58 B 0.01371f
C621 VDD1.n59 B 0.056188f
C622 VDD1.n60 B 0.078615f
C623 VDD1.t2 B 0.22824f
C624 VDD1.t5 B 0.22824f
C625 VDD1.n61 B 2.02461f
C626 VDD1.n62 B 0.905131f
C627 VDD1.n63 B 0.033798f
C628 VDD1.n64 B 0.025515f
C629 VDD1.n65 B 0.01371f
C630 VDD1.n66 B 0.032407f
C631 VDD1.n67 B 0.014517f
C632 VDD1.n68 B 0.025515f
C633 VDD1.n69 B 0.01371f
C634 VDD1.n70 B 0.032407f
C635 VDD1.n71 B 0.014114f
C636 VDD1.n72 B 0.025515f
C637 VDD1.n73 B 0.014517f
C638 VDD1.n74 B 0.032407f
C639 VDD1.n75 B 0.014517f
C640 VDD1.n76 B 0.025515f
C641 VDD1.n77 B 0.01371f
C642 VDD1.n78 B 0.032407f
C643 VDD1.n79 B 0.014517f
C644 VDD1.n80 B 1.21001f
C645 VDD1.n81 B 0.01371f
C646 VDD1.t0 B 0.05464f
C647 VDD1.n82 B 0.177298f
C648 VDD1.n83 B 0.022909f
C649 VDD1.n84 B 0.024305f
C650 VDD1.n85 B 0.032407f
C651 VDD1.n86 B 0.014517f
C652 VDD1.n87 B 0.01371f
C653 VDD1.n88 B 0.025515f
C654 VDD1.n89 B 0.025515f
C655 VDD1.n90 B 0.01371f
C656 VDD1.n91 B 0.014517f
C657 VDD1.n92 B 0.032407f
C658 VDD1.n93 B 0.032407f
C659 VDD1.n94 B 0.014517f
C660 VDD1.n95 B 0.01371f
C661 VDD1.n96 B 0.025515f
C662 VDD1.n97 B 0.025515f
C663 VDD1.n98 B 0.01371f
C664 VDD1.n99 B 0.01371f
C665 VDD1.n100 B 0.014517f
C666 VDD1.n101 B 0.032407f
C667 VDD1.n102 B 0.032407f
C668 VDD1.n103 B 0.032407f
C669 VDD1.n104 B 0.014114f
C670 VDD1.n105 B 0.01371f
C671 VDD1.n106 B 0.025515f
C672 VDD1.n107 B 0.025515f
C673 VDD1.n108 B 0.01371f
C674 VDD1.n109 B 0.014517f
C675 VDD1.n110 B 0.032407f
C676 VDD1.n111 B 0.032407f
C677 VDD1.n112 B 0.014517f
C678 VDD1.n113 B 0.01371f
C679 VDD1.n114 B 0.025515f
C680 VDD1.n115 B 0.025515f
C681 VDD1.n116 B 0.01371f
C682 VDD1.n117 B 0.014517f
C683 VDD1.n118 B 0.032407f
C684 VDD1.n119 B 0.066502f
C685 VDD1.n120 B 0.014517f
C686 VDD1.n121 B 0.01371f
C687 VDD1.n122 B 0.056188f
C688 VDD1.n123 B 0.078615f
C689 VDD1.t9 B 0.22824f
C690 VDD1.t4 B 0.22824f
C691 VDD1.n124 B 2.0246f
C692 VDD1.n125 B 0.896507f
C693 VDD1.t8 B 0.22824f
C694 VDD1.t1 B 0.22824f
C695 VDD1.n126 B 2.05533f
C696 VDD1.n127 B 3.74281f
C697 VDD1.t3 B 0.22824f
C698 VDD1.t6 B 0.22824f
C699 VDD1.n128 B 2.0246f
C700 VDD1.n129 B 3.71275f
C701 VP.t1 B 2.0281f
C702 VP.n0 B 0.779317f
C703 VP.n1 B 0.017153f
C704 VP.n2 B 0.034185f
C705 VP.n3 B 0.017153f
C706 VP.n4 B 0.03213f
C707 VP.n5 B 0.017153f
C708 VP.t5 B 2.0281f
C709 VP.n6 B 0.03213f
C710 VP.n7 B 0.017153f
C711 VP.n8 B 0.03213f
C712 VP.n9 B 0.017153f
C713 VP.t7 B 2.0281f
C714 VP.n10 B 0.03213f
C715 VP.n11 B 0.017153f
C716 VP.n12 B 0.03213f
C717 VP.n13 B 0.017153f
C718 VP.t9 B 2.0281f
C719 VP.n14 B 0.03213f
C720 VP.n15 B 0.017153f
C721 VP.n16 B 0.03213f
C722 VP.n17 B 0.02769f
C723 VP.t2 B 2.0281f
C724 VP.t3 B 2.0281f
C725 VP.n18 B 0.779317f
C726 VP.n19 B 0.017153f
C727 VP.n20 B 0.034185f
C728 VP.n21 B 0.017153f
C729 VP.n22 B 0.03213f
C730 VP.n23 B 0.017153f
C731 VP.t8 B 2.0281f
C732 VP.n24 B 0.03213f
C733 VP.n25 B 0.017153f
C734 VP.n26 B 0.03213f
C735 VP.n27 B 0.017153f
C736 VP.t4 B 2.0281f
C737 VP.n28 B 0.03213f
C738 VP.n29 B 0.017153f
C739 VP.n30 B 0.03213f
C740 VP.t6 B 2.29905f
C741 VP.n31 B 0.739761f
C742 VP.t0 B 2.0281f
C743 VP.n32 B 0.780506f
C744 VP.n33 B 0.029592f
C745 VP.n34 B 0.221004f
C746 VP.n35 B 0.017153f
C747 VP.n36 B 0.017153f
C748 VP.n37 B 0.03213f
C749 VP.n38 B 0.021058f
C750 VP.n39 B 0.029242f
C751 VP.n40 B 0.017153f
C752 VP.n41 B 0.017153f
C753 VP.n42 B 0.017153f
C754 VP.n43 B 0.03213f
C755 VP.n44 B 0.024198f
C756 VP.n45 B 0.712408f
C757 VP.n46 B 0.024198f
C758 VP.n47 B 0.017153f
C759 VP.n48 B 0.017153f
C760 VP.n49 B 0.017153f
C761 VP.n50 B 0.03213f
C762 VP.n51 B 0.029242f
C763 VP.n52 B 0.021058f
C764 VP.n53 B 0.017153f
C765 VP.n54 B 0.017153f
C766 VP.n55 B 0.017153f
C767 VP.n56 B 0.03213f
C768 VP.n57 B 0.029592f
C769 VP.n58 B 0.712408f
C770 VP.n59 B 0.018804f
C771 VP.n60 B 0.017153f
C772 VP.n61 B 0.017153f
C773 VP.n62 B 0.017153f
C774 VP.n63 B 0.03213f
C775 VP.n64 B 0.034359f
C776 VP.n65 B 0.013886f
C777 VP.n66 B 0.017153f
C778 VP.n67 B 0.017153f
C779 VP.n68 B 0.017153f
C780 VP.n69 B 0.03213f
C781 VP.n70 B 0.03213f
C782 VP.n71 B 0.019122f
C783 VP.n72 B 0.02769f
C784 VP.n73 B 1.25166f
C785 VP.n74 B 1.262f
C786 VP.n75 B 0.779317f
C787 VP.n76 B 0.019122f
C788 VP.n77 B 0.03213f
C789 VP.n78 B 0.017153f
C790 VP.n79 B 0.017153f
C791 VP.n80 B 0.017153f
C792 VP.n81 B 0.034185f
C793 VP.n82 B 0.013886f
C794 VP.n83 B 0.034359f
C795 VP.n84 B 0.017153f
C796 VP.n85 B 0.017153f
C797 VP.n86 B 0.017153f
C798 VP.n87 B 0.03213f
C799 VP.n88 B 0.018804f
C800 VP.n89 B 0.712408f
C801 VP.n90 B 0.029592f
C802 VP.n91 B 0.017153f
C803 VP.n92 B 0.017153f
C804 VP.n93 B 0.017153f
C805 VP.n94 B 0.03213f
C806 VP.n95 B 0.021058f
C807 VP.n96 B 0.029242f
C808 VP.n97 B 0.017153f
C809 VP.n98 B 0.017153f
C810 VP.n99 B 0.017153f
C811 VP.n100 B 0.03213f
C812 VP.n101 B 0.024198f
C813 VP.n102 B 0.712408f
C814 VP.n103 B 0.024198f
C815 VP.n104 B 0.017153f
C816 VP.n105 B 0.017153f
C817 VP.n106 B 0.017153f
C818 VP.n107 B 0.03213f
C819 VP.n108 B 0.029242f
C820 VP.n109 B 0.021058f
C821 VP.n110 B 0.017153f
C822 VP.n111 B 0.017153f
C823 VP.n112 B 0.017153f
C824 VP.n113 B 0.03213f
C825 VP.n114 B 0.029592f
C826 VP.n115 B 0.712408f
C827 VP.n116 B 0.018804f
C828 VP.n117 B 0.017153f
C829 VP.n118 B 0.017153f
C830 VP.n119 B 0.017153f
C831 VP.n120 B 0.03213f
C832 VP.n121 B 0.034359f
C833 VP.n122 B 0.013886f
C834 VP.n123 B 0.017153f
C835 VP.n124 B 0.017153f
C836 VP.n125 B 0.017153f
C837 VP.n126 B 0.03213f
C838 VP.n127 B 0.03213f
C839 VP.n128 B 0.019122f
C840 VP.n129 B 0.02769f
C841 VP.n130 B 0.052344f
.ends

