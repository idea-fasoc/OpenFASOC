* NGSPICE file created from diff_pair_sample_0858.ext - technology: sky130A

.subckt diff_pair_sample_0858 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=2.19945 ps=13.66 w=13.33 l=4
X1 B.t11 B.t9 B.t10 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=0 ps=0 w=13.33 l=4
X2 VDD1.t5 VP.t0 VTAIL.t0 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=5.1987 ps=27.44 w=13.33 l=4
X3 VTAIL.t3 VP.t1 VDD1.t4 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=2.19945 ps=13.66 w=13.33 l=4
X4 VTAIL.t11 VN.t1 VDD2.t4 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=2.19945 ps=13.66 w=13.33 l=4
X5 VDD1.t3 VP.t2 VTAIL.t4 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=2.19945 ps=13.66 w=13.33 l=4
X6 VDD1.t2 VP.t3 VTAIL.t5 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=5.1987 ps=27.44 w=13.33 l=4
X7 VDD2.t3 VN.t2 VTAIL.t8 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=5.1987 ps=27.44 w=13.33 l=4
X8 B.t8 B.t6 B.t7 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=0 ps=0 w=13.33 l=4
X9 VTAIL.t2 VP.t4 VDD1.t1 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=2.19945 ps=13.66 w=13.33 l=4
X10 B.t5 B.t3 B.t4 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=0 ps=0 w=13.33 l=4
X11 B.t2 B.t0 B.t1 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=0 ps=0 w=13.33 l=4
X12 VDD1.t0 VP.t5 VTAIL.t1 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=2.19945 ps=13.66 w=13.33 l=4
X13 VTAIL.t6 VN.t3 VDD2.t2 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=2.19945 ps=13.66 w=13.33 l=4
X14 VDD2.t1 VN.t4 VTAIL.t10 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=2.19945 pd=13.66 as=5.1987 ps=27.44 w=13.33 l=4
X15 VDD2.t0 VN.t5 VTAIL.t7 w_n4434_n3634# sky130_fd_pr__pfet_01v8 ad=5.1987 pd=27.44 as=2.19945 ps=13.66 w=13.33 l=4
R0 VN.n37 VN.n20 161.3
R1 VN.n36 VN.n35 161.3
R2 VN.n34 VN.n21 161.3
R3 VN.n33 VN.n32 161.3
R4 VN.n31 VN.n22 161.3
R5 VN.n30 VN.n29 161.3
R6 VN.n28 VN.n23 161.3
R7 VN.n27 VN.n26 161.3
R8 VN.n17 VN.n0 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n1 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n11 VN.n2 161.3
R13 VN.n10 VN.n9 161.3
R14 VN.n8 VN.n3 161.3
R15 VN.n7 VN.n6 161.3
R16 VN.n4 VN.t5 113.513
R17 VN.n24 VN.t2 113.513
R18 VN.n5 VN.t1 80.3137
R19 VN.n18 VN.t4 80.3137
R20 VN.n25 VN.t3 80.3137
R21 VN.n38 VN.t0 80.3137
R22 VN.n19 VN.n18 66.0336
R23 VN.n39 VN.n38 66.0336
R24 VN.n12 VN.n11 56.5193
R25 VN.n32 VN.n31 56.5193
R26 VN VN.n39 55.3943
R27 VN.n25 VN.n24 50.5569
R28 VN.n5 VN.n4 50.5569
R29 VN.n6 VN.n5 24.4675
R30 VN.n6 VN.n3 24.4675
R31 VN.n10 VN.n3 24.4675
R32 VN.n11 VN.n10 24.4675
R33 VN.n12 VN.n1 24.4675
R34 VN.n16 VN.n1 24.4675
R35 VN.n17 VN.n16 24.4675
R36 VN.n31 VN.n30 24.4675
R37 VN.n30 VN.n23 24.4675
R38 VN.n26 VN.n23 24.4675
R39 VN.n26 VN.n25 24.4675
R40 VN.n37 VN.n36 24.4675
R41 VN.n36 VN.n21 24.4675
R42 VN.n32 VN.n21 24.4675
R43 VN.n18 VN.n17 16.1487
R44 VN.n38 VN.n37 16.1487
R45 VN.n7 VN.n4 2.09747
R46 VN.n27 VN.n24 2.09747
R47 VN.n39 VN.n20 0.417535
R48 VN.n19 VN.n0 0.417535
R49 VN VN.n19 0.394291
R50 VN.n35 VN.n20 0.189894
R51 VN.n35 VN.n34 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n22 0.189894
R54 VN.n29 VN.n22 0.189894
R55 VN.n29 VN.n28 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n9 VN.n8 0.189894
R59 VN.n9 VN.n2 0.189894
R60 VN.n13 VN.n2 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n15 VN.n14 0.189894
R63 VN.n15 VN.n0 0.189894
R64 VTAIL.n249 VTAIL.n248 585
R65 VTAIL.n251 VTAIL.n250 585
R66 VTAIL.n244 VTAIL.n243 585
R67 VTAIL.n257 VTAIL.n256 585
R68 VTAIL.n259 VTAIL.n258 585
R69 VTAIL.n240 VTAIL.n239 585
R70 VTAIL.n265 VTAIL.n264 585
R71 VTAIL.n267 VTAIL.n266 585
R72 VTAIL.n236 VTAIL.n235 585
R73 VTAIL.n273 VTAIL.n272 585
R74 VTAIL.n275 VTAIL.n274 585
R75 VTAIL.n232 VTAIL.n231 585
R76 VTAIL.n281 VTAIL.n280 585
R77 VTAIL.n283 VTAIL.n282 585
R78 VTAIL.n228 VTAIL.n227 585
R79 VTAIL.n289 VTAIL.n288 585
R80 VTAIL.n291 VTAIL.n290 585
R81 VTAIL.n27 VTAIL.n26 585
R82 VTAIL.n29 VTAIL.n28 585
R83 VTAIL.n22 VTAIL.n21 585
R84 VTAIL.n35 VTAIL.n34 585
R85 VTAIL.n37 VTAIL.n36 585
R86 VTAIL.n18 VTAIL.n17 585
R87 VTAIL.n43 VTAIL.n42 585
R88 VTAIL.n45 VTAIL.n44 585
R89 VTAIL.n14 VTAIL.n13 585
R90 VTAIL.n51 VTAIL.n50 585
R91 VTAIL.n53 VTAIL.n52 585
R92 VTAIL.n10 VTAIL.n9 585
R93 VTAIL.n59 VTAIL.n58 585
R94 VTAIL.n61 VTAIL.n60 585
R95 VTAIL.n6 VTAIL.n5 585
R96 VTAIL.n67 VTAIL.n66 585
R97 VTAIL.n69 VTAIL.n68 585
R98 VTAIL.n219 VTAIL.n218 585
R99 VTAIL.n217 VTAIL.n216 585
R100 VTAIL.n156 VTAIL.n155 585
R101 VTAIL.n211 VTAIL.n210 585
R102 VTAIL.n209 VTAIL.n208 585
R103 VTAIL.n160 VTAIL.n159 585
R104 VTAIL.n203 VTAIL.n202 585
R105 VTAIL.n201 VTAIL.n200 585
R106 VTAIL.n164 VTAIL.n163 585
R107 VTAIL.n195 VTAIL.n194 585
R108 VTAIL.n193 VTAIL.n192 585
R109 VTAIL.n168 VTAIL.n167 585
R110 VTAIL.n187 VTAIL.n186 585
R111 VTAIL.n185 VTAIL.n184 585
R112 VTAIL.n172 VTAIL.n171 585
R113 VTAIL.n179 VTAIL.n178 585
R114 VTAIL.n177 VTAIL.n176 585
R115 VTAIL.n145 VTAIL.n144 585
R116 VTAIL.n143 VTAIL.n142 585
R117 VTAIL.n82 VTAIL.n81 585
R118 VTAIL.n137 VTAIL.n136 585
R119 VTAIL.n135 VTAIL.n134 585
R120 VTAIL.n86 VTAIL.n85 585
R121 VTAIL.n129 VTAIL.n128 585
R122 VTAIL.n127 VTAIL.n126 585
R123 VTAIL.n90 VTAIL.n89 585
R124 VTAIL.n121 VTAIL.n120 585
R125 VTAIL.n119 VTAIL.n118 585
R126 VTAIL.n94 VTAIL.n93 585
R127 VTAIL.n113 VTAIL.n112 585
R128 VTAIL.n111 VTAIL.n110 585
R129 VTAIL.n98 VTAIL.n97 585
R130 VTAIL.n105 VTAIL.n104 585
R131 VTAIL.n103 VTAIL.n102 585
R132 VTAIL.n290 VTAIL.n224 498.474
R133 VTAIL.n68 VTAIL.n2 498.474
R134 VTAIL.n218 VTAIL.n152 498.474
R135 VTAIL.n144 VTAIL.n78 498.474
R136 VTAIL.n247 VTAIL.t10 327.466
R137 VTAIL.n25 VTAIL.t5 327.466
R138 VTAIL.n175 VTAIL.t0 327.466
R139 VTAIL.n101 VTAIL.t8 327.466
R140 VTAIL.n250 VTAIL.n249 171.744
R141 VTAIL.n250 VTAIL.n243 171.744
R142 VTAIL.n257 VTAIL.n243 171.744
R143 VTAIL.n258 VTAIL.n257 171.744
R144 VTAIL.n258 VTAIL.n239 171.744
R145 VTAIL.n265 VTAIL.n239 171.744
R146 VTAIL.n266 VTAIL.n265 171.744
R147 VTAIL.n266 VTAIL.n235 171.744
R148 VTAIL.n273 VTAIL.n235 171.744
R149 VTAIL.n274 VTAIL.n273 171.744
R150 VTAIL.n274 VTAIL.n231 171.744
R151 VTAIL.n281 VTAIL.n231 171.744
R152 VTAIL.n282 VTAIL.n281 171.744
R153 VTAIL.n282 VTAIL.n227 171.744
R154 VTAIL.n289 VTAIL.n227 171.744
R155 VTAIL.n290 VTAIL.n289 171.744
R156 VTAIL.n28 VTAIL.n27 171.744
R157 VTAIL.n28 VTAIL.n21 171.744
R158 VTAIL.n35 VTAIL.n21 171.744
R159 VTAIL.n36 VTAIL.n35 171.744
R160 VTAIL.n36 VTAIL.n17 171.744
R161 VTAIL.n43 VTAIL.n17 171.744
R162 VTAIL.n44 VTAIL.n43 171.744
R163 VTAIL.n44 VTAIL.n13 171.744
R164 VTAIL.n51 VTAIL.n13 171.744
R165 VTAIL.n52 VTAIL.n51 171.744
R166 VTAIL.n52 VTAIL.n9 171.744
R167 VTAIL.n59 VTAIL.n9 171.744
R168 VTAIL.n60 VTAIL.n59 171.744
R169 VTAIL.n60 VTAIL.n5 171.744
R170 VTAIL.n67 VTAIL.n5 171.744
R171 VTAIL.n68 VTAIL.n67 171.744
R172 VTAIL.n218 VTAIL.n217 171.744
R173 VTAIL.n217 VTAIL.n155 171.744
R174 VTAIL.n210 VTAIL.n155 171.744
R175 VTAIL.n210 VTAIL.n209 171.744
R176 VTAIL.n209 VTAIL.n159 171.744
R177 VTAIL.n202 VTAIL.n159 171.744
R178 VTAIL.n202 VTAIL.n201 171.744
R179 VTAIL.n201 VTAIL.n163 171.744
R180 VTAIL.n194 VTAIL.n163 171.744
R181 VTAIL.n194 VTAIL.n193 171.744
R182 VTAIL.n193 VTAIL.n167 171.744
R183 VTAIL.n186 VTAIL.n167 171.744
R184 VTAIL.n186 VTAIL.n185 171.744
R185 VTAIL.n185 VTAIL.n171 171.744
R186 VTAIL.n178 VTAIL.n171 171.744
R187 VTAIL.n178 VTAIL.n177 171.744
R188 VTAIL.n144 VTAIL.n143 171.744
R189 VTAIL.n143 VTAIL.n81 171.744
R190 VTAIL.n136 VTAIL.n81 171.744
R191 VTAIL.n136 VTAIL.n135 171.744
R192 VTAIL.n135 VTAIL.n85 171.744
R193 VTAIL.n128 VTAIL.n85 171.744
R194 VTAIL.n128 VTAIL.n127 171.744
R195 VTAIL.n127 VTAIL.n89 171.744
R196 VTAIL.n120 VTAIL.n89 171.744
R197 VTAIL.n120 VTAIL.n119 171.744
R198 VTAIL.n119 VTAIL.n93 171.744
R199 VTAIL.n112 VTAIL.n93 171.744
R200 VTAIL.n112 VTAIL.n111 171.744
R201 VTAIL.n111 VTAIL.n97 171.744
R202 VTAIL.n104 VTAIL.n97 171.744
R203 VTAIL.n104 VTAIL.n103 171.744
R204 VTAIL.n249 VTAIL.t10 85.8723
R205 VTAIL.n27 VTAIL.t5 85.8723
R206 VTAIL.n177 VTAIL.t0 85.8723
R207 VTAIL.n103 VTAIL.t8 85.8723
R208 VTAIL.n151 VTAIL.n150 57.809
R209 VTAIL.n77 VTAIL.n76 57.809
R210 VTAIL.n1 VTAIL.n0 57.8088
R211 VTAIL.n75 VTAIL.n74 57.8088
R212 VTAIL.n295 VTAIL.n294 34.7066
R213 VTAIL.n73 VTAIL.n72 34.7066
R214 VTAIL.n223 VTAIL.n222 34.7066
R215 VTAIL.n149 VTAIL.n148 34.7066
R216 VTAIL.n77 VTAIL.n75 31.3238
R217 VTAIL.n295 VTAIL.n223 27.591
R218 VTAIL.n248 VTAIL.n247 16.3895
R219 VTAIL.n26 VTAIL.n25 16.3895
R220 VTAIL.n176 VTAIL.n175 16.3895
R221 VTAIL.n102 VTAIL.n101 16.3895
R222 VTAIL.n251 VTAIL.n246 12.8005
R223 VTAIL.n292 VTAIL.n291 12.8005
R224 VTAIL.n29 VTAIL.n24 12.8005
R225 VTAIL.n70 VTAIL.n69 12.8005
R226 VTAIL.n220 VTAIL.n219 12.8005
R227 VTAIL.n179 VTAIL.n174 12.8005
R228 VTAIL.n146 VTAIL.n145 12.8005
R229 VTAIL.n105 VTAIL.n100 12.8005
R230 VTAIL.n252 VTAIL.n244 12.0247
R231 VTAIL.n288 VTAIL.n226 12.0247
R232 VTAIL.n30 VTAIL.n22 12.0247
R233 VTAIL.n66 VTAIL.n4 12.0247
R234 VTAIL.n216 VTAIL.n154 12.0247
R235 VTAIL.n180 VTAIL.n172 12.0247
R236 VTAIL.n142 VTAIL.n80 12.0247
R237 VTAIL.n106 VTAIL.n98 12.0247
R238 VTAIL.n256 VTAIL.n255 11.249
R239 VTAIL.n287 VTAIL.n228 11.249
R240 VTAIL.n34 VTAIL.n33 11.249
R241 VTAIL.n65 VTAIL.n6 11.249
R242 VTAIL.n215 VTAIL.n156 11.249
R243 VTAIL.n184 VTAIL.n183 11.249
R244 VTAIL.n141 VTAIL.n82 11.249
R245 VTAIL.n110 VTAIL.n109 11.249
R246 VTAIL.n259 VTAIL.n242 10.4732
R247 VTAIL.n284 VTAIL.n283 10.4732
R248 VTAIL.n37 VTAIL.n20 10.4732
R249 VTAIL.n62 VTAIL.n61 10.4732
R250 VTAIL.n212 VTAIL.n211 10.4732
R251 VTAIL.n187 VTAIL.n170 10.4732
R252 VTAIL.n138 VTAIL.n137 10.4732
R253 VTAIL.n113 VTAIL.n96 10.4732
R254 VTAIL.n260 VTAIL.n240 9.69747
R255 VTAIL.n280 VTAIL.n230 9.69747
R256 VTAIL.n38 VTAIL.n18 9.69747
R257 VTAIL.n58 VTAIL.n8 9.69747
R258 VTAIL.n208 VTAIL.n158 9.69747
R259 VTAIL.n188 VTAIL.n168 9.69747
R260 VTAIL.n134 VTAIL.n84 9.69747
R261 VTAIL.n114 VTAIL.n94 9.69747
R262 VTAIL.n294 VTAIL.n293 9.45567
R263 VTAIL.n72 VTAIL.n71 9.45567
R264 VTAIL.n222 VTAIL.n221 9.45567
R265 VTAIL.n148 VTAIL.n147 9.45567
R266 VTAIL.n269 VTAIL.n268 9.3005
R267 VTAIL.n238 VTAIL.n237 9.3005
R268 VTAIL.n263 VTAIL.n262 9.3005
R269 VTAIL.n261 VTAIL.n260 9.3005
R270 VTAIL.n242 VTAIL.n241 9.3005
R271 VTAIL.n255 VTAIL.n254 9.3005
R272 VTAIL.n253 VTAIL.n252 9.3005
R273 VTAIL.n246 VTAIL.n245 9.3005
R274 VTAIL.n271 VTAIL.n270 9.3005
R275 VTAIL.n234 VTAIL.n233 9.3005
R276 VTAIL.n277 VTAIL.n276 9.3005
R277 VTAIL.n279 VTAIL.n278 9.3005
R278 VTAIL.n230 VTAIL.n229 9.3005
R279 VTAIL.n285 VTAIL.n284 9.3005
R280 VTAIL.n287 VTAIL.n286 9.3005
R281 VTAIL.n226 VTAIL.n225 9.3005
R282 VTAIL.n293 VTAIL.n292 9.3005
R283 VTAIL.n47 VTAIL.n46 9.3005
R284 VTAIL.n16 VTAIL.n15 9.3005
R285 VTAIL.n41 VTAIL.n40 9.3005
R286 VTAIL.n39 VTAIL.n38 9.3005
R287 VTAIL.n20 VTAIL.n19 9.3005
R288 VTAIL.n33 VTAIL.n32 9.3005
R289 VTAIL.n31 VTAIL.n30 9.3005
R290 VTAIL.n24 VTAIL.n23 9.3005
R291 VTAIL.n49 VTAIL.n48 9.3005
R292 VTAIL.n12 VTAIL.n11 9.3005
R293 VTAIL.n55 VTAIL.n54 9.3005
R294 VTAIL.n57 VTAIL.n56 9.3005
R295 VTAIL.n8 VTAIL.n7 9.3005
R296 VTAIL.n63 VTAIL.n62 9.3005
R297 VTAIL.n65 VTAIL.n64 9.3005
R298 VTAIL.n4 VTAIL.n3 9.3005
R299 VTAIL.n71 VTAIL.n70 9.3005
R300 VTAIL.n162 VTAIL.n161 9.3005
R301 VTAIL.n205 VTAIL.n204 9.3005
R302 VTAIL.n207 VTAIL.n206 9.3005
R303 VTAIL.n158 VTAIL.n157 9.3005
R304 VTAIL.n213 VTAIL.n212 9.3005
R305 VTAIL.n215 VTAIL.n214 9.3005
R306 VTAIL.n154 VTAIL.n153 9.3005
R307 VTAIL.n221 VTAIL.n220 9.3005
R308 VTAIL.n199 VTAIL.n198 9.3005
R309 VTAIL.n197 VTAIL.n196 9.3005
R310 VTAIL.n166 VTAIL.n165 9.3005
R311 VTAIL.n191 VTAIL.n190 9.3005
R312 VTAIL.n189 VTAIL.n188 9.3005
R313 VTAIL.n170 VTAIL.n169 9.3005
R314 VTAIL.n183 VTAIL.n182 9.3005
R315 VTAIL.n181 VTAIL.n180 9.3005
R316 VTAIL.n174 VTAIL.n173 9.3005
R317 VTAIL.n88 VTAIL.n87 9.3005
R318 VTAIL.n131 VTAIL.n130 9.3005
R319 VTAIL.n133 VTAIL.n132 9.3005
R320 VTAIL.n84 VTAIL.n83 9.3005
R321 VTAIL.n139 VTAIL.n138 9.3005
R322 VTAIL.n141 VTAIL.n140 9.3005
R323 VTAIL.n80 VTAIL.n79 9.3005
R324 VTAIL.n147 VTAIL.n146 9.3005
R325 VTAIL.n125 VTAIL.n124 9.3005
R326 VTAIL.n123 VTAIL.n122 9.3005
R327 VTAIL.n92 VTAIL.n91 9.3005
R328 VTAIL.n117 VTAIL.n116 9.3005
R329 VTAIL.n115 VTAIL.n114 9.3005
R330 VTAIL.n96 VTAIL.n95 9.3005
R331 VTAIL.n109 VTAIL.n108 9.3005
R332 VTAIL.n107 VTAIL.n106 9.3005
R333 VTAIL.n100 VTAIL.n99 9.3005
R334 VTAIL.n264 VTAIL.n263 8.92171
R335 VTAIL.n279 VTAIL.n232 8.92171
R336 VTAIL.n42 VTAIL.n41 8.92171
R337 VTAIL.n57 VTAIL.n10 8.92171
R338 VTAIL.n207 VTAIL.n160 8.92171
R339 VTAIL.n192 VTAIL.n191 8.92171
R340 VTAIL.n133 VTAIL.n86 8.92171
R341 VTAIL.n118 VTAIL.n117 8.92171
R342 VTAIL.n267 VTAIL.n238 8.14595
R343 VTAIL.n276 VTAIL.n275 8.14595
R344 VTAIL.n45 VTAIL.n16 8.14595
R345 VTAIL.n54 VTAIL.n53 8.14595
R346 VTAIL.n204 VTAIL.n203 8.14595
R347 VTAIL.n195 VTAIL.n166 8.14595
R348 VTAIL.n130 VTAIL.n129 8.14595
R349 VTAIL.n121 VTAIL.n92 8.14595
R350 VTAIL.n294 VTAIL.n224 7.75445
R351 VTAIL.n72 VTAIL.n2 7.75445
R352 VTAIL.n222 VTAIL.n152 7.75445
R353 VTAIL.n148 VTAIL.n78 7.75445
R354 VTAIL.n268 VTAIL.n236 7.3702
R355 VTAIL.n272 VTAIL.n234 7.3702
R356 VTAIL.n46 VTAIL.n14 7.3702
R357 VTAIL.n50 VTAIL.n12 7.3702
R358 VTAIL.n200 VTAIL.n162 7.3702
R359 VTAIL.n196 VTAIL.n164 7.3702
R360 VTAIL.n126 VTAIL.n88 7.3702
R361 VTAIL.n122 VTAIL.n90 7.3702
R362 VTAIL.n271 VTAIL.n236 6.59444
R363 VTAIL.n272 VTAIL.n271 6.59444
R364 VTAIL.n49 VTAIL.n14 6.59444
R365 VTAIL.n50 VTAIL.n49 6.59444
R366 VTAIL.n200 VTAIL.n199 6.59444
R367 VTAIL.n199 VTAIL.n164 6.59444
R368 VTAIL.n126 VTAIL.n125 6.59444
R369 VTAIL.n125 VTAIL.n90 6.59444
R370 VTAIL.n292 VTAIL.n224 6.08283
R371 VTAIL.n70 VTAIL.n2 6.08283
R372 VTAIL.n220 VTAIL.n152 6.08283
R373 VTAIL.n146 VTAIL.n78 6.08283
R374 VTAIL.n268 VTAIL.n267 5.81868
R375 VTAIL.n275 VTAIL.n234 5.81868
R376 VTAIL.n46 VTAIL.n45 5.81868
R377 VTAIL.n53 VTAIL.n12 5.81868
R378 VTAIL.n203 VTAIL.n162 5.81868
R379 VTAIL.n196 VTAIL.n195 5.81868
R380 VTAIL.n129 VTAIL.n88 5.81868
R381 VTAIL.n122 VTAIL.n121 5.81868
R382 VTAIL.n264 VTAIL.n238 5.04292
R383 VTAIL.n276 VTAIL.n232 5.04292
R384 VTAIL.n42 VTAIL.n16 5.04292
R385 VTAIL.n54 VTAIL.n10 5.04292
R386 VTAIL.n204 VTAIL.n160 5.04292
R387 VTAIL.n192 VTAIL.n166 5.04292
R388 VTAIL.n130 VTAIL.n86 5.04292
R389 VTAIL.n118 VTAIL.n92 5.04292
R390 VTAIL.n263 VTAIL.n240 4.26717
R391 VTAIL.n280 VTAIL.n279 4.26717
R392 VTAIL.n41 VTAIL.n18 4.26717
R393 VTAIL.n58 VTAIL.n57 4.26717
R394 VTAIL.n208 VTAIL.n207 4.26717
R395 VTAIL.n191 VTAIL.n168 4.26717
R396 VTAIL.n134 VTAIL.n133 4.26717
R397 VTAIL.n117 VTAIL.n94 4.26717
R398 VTAIL.n149 VTAIL.n77 3.73326
R399 VTAIL.n223 VTAIL.n151 3.73326
R400 VTAIL.n75 VTAIL.n73 3.73326
R401 VTAIL.n247 VTAIL.n245 3.70982
R402 VTAIL.n25 VTAIL.n23 3.70982
R403 VTAIL.n175 VTAIL.n173 3.70982
R404 VTAIL.n101 VTAIL.n99 3.70982
R405 VTAIL.n260 VTAIL.n259 3.49141
R406 VTAIL.n283 VTAIL.n230 3.49141
R407 VTAIL.n38 VTAIL.n37 3.49141
R408 VTAIL.n61 VTAIL.n8 3.49141
R409 VTAIL.n211 VTAIL.n158 3.49141
R410 VTAIL.n188 VTAIL.n187 3.49141
R411 VTAIL.n137 VTAIL.n84 3.49141
R412 VTAIL.n114 VTAIL.n113 3.49141
R413 VTAIL VTAIL.n295 2.74188
R414 VTAIL.n256 VTAIL.n242 2.71565
R415 VTAIL.n284 VTAIL.n228 2.71565
R416 VTAIL.n34 VTAIL.n20 2.71565
R417 VTAIL.n62 VTAIL.n6 2.71565
R418 VTAIL.n212 VTAIL.n156 2.71565
R419 VTAIL.n184 VTAIL.n170 2.71565
R420 VTAIL.n138 VTAIL.n82 2.71565
R421 VTAIL.n110 VTAIL.n96 2.71565
R422 VTAIL.n0 VTAIL.t7 2.43898
R423 VTAIL.n0 VTAIL.t11 2.43898
R424 VTAIL.n74 VTAIL.t4 2.43898
R425 VTAIL.n74 VTAIL.t2 2.43898
R426 VTAIL.n150 VTAIL.t1 2.43898
R427 VTAIL.n150 VTAIL.t3 2.43898
R428 VTAIL.n76 VTAIL.t9 2.43898
R429 VTAIL.n76 VTAIL.t6 2.43898
R430 VTAIL.n151 VTAIL.n149 2.33671
R431 VTAIL.n73 VTAIL.n1 2.33671
R432 VTAIL.n255 VTAIL.n244 1.93989
R433 VTAIL.n288 VTAIL.n287 1.93989
R434 VTAIL.n33 VTAIL.n22 1.93989
R435 VTAIL.n66 VTAIL.n65 1.93989
R436 VTAIL.n216 VTAIL.n215 1.93989
R437 VTAIL.n183 VTAIL.n172 1.93989
R438 VTAIL.n142 VTAIL.n141 1.93989
R439 VTAIL.n109 VTAIL.n98 1.93989
R440 VTAIL.n252 VTAIL.n251 1.16414
R441 VTAIL.n291 VTAIL.n226 1.16414
R442 VTAIL.n30 VTAIL.n29 1.16414
R443 VTAIL.n69 VTAIL.n4 1.16414
R444 VTAIL.n219 VTAIL.n154 1.16414
R445 VTAIL.n180 VTAIL.n179 1.16414
R446 VTAIL.n145 VTAIL.n80 1.16414
R447 VTAIL.n106 VTAIL.n105 1.16414
R448 VTAIL VTAIL.n1 0.991879
R449 VTAIL.n248 VTAIL.n246 0.388379
R450 VTAIL.n26 VTAIL.n24 0.388379
R451 VTAIL.n176 VTAIL.n174 0.388379
R452 VTAIL.n102 VTAIL.n100 0.388379
R453 VTAIL.n253 VTAIL.n245 0.155672
R454 VTAIL.n254 VTAIL.n253 0.155672
R455 VTAIL.n254 VTAIL.n241 0.155672
R456 VTAIL.n261 VTAIL.n241 0.155672
R457 VTAIL.n262 VTAIL.n261 0.155672
R458 VTAIL.n262 VTAIL.n237 0.155672
R459 VTAIL.n269 VTAIL.n237 0.155672
R460 VTAIL.n270 VTAIL.n269 0.155672
R461 VTAIL.n270 VTAIL.n233 0.155672
R462 VTAIL.n277 VTAIL.n233 0.155672
R463 VTAIL.n278 VTAIL.n277 0.155672
R464 VTAIL.n278 VTAIL.n229 0.155672
R465 VTAIL.n285 VTAIL.n229 0.155672
R466 VTAIL.n286 VTAIL.n285 0.155672
R467 VTAIL.n286 VTAIL.n225 0.155672
R468 VTAIL.n293 VTAIL.n225 0.155672
R469 VTAIL.n31 VTAIL.n23 0.155672
R470 VTAIL.n32 VTAIL.n31 0.155672
R471 VTAIL.n32 VTAIL.n19 0.155672
R472 VTAIL.n39 VTAIL.n19 0.155672
R473 VTAIL.n40 VTAIL.n39 0.155672
R474 VTAIL.n40 VTAIL.n15 0.155672
R475 VTAIL.n47 VTAIL.n15 0.155672
R476 VTAIL.n48 VTAIL.n47 0.155672
R477 VTAIL.n48 VTAIL.n11 0.155672
R478 VTAIL.n55 VTAIL.n11 0.155672
R479 VTAIL.n56 VTAIL.n55 0.155672
R480 VTAIL.n56 VTAIL.n7 0.155672
R481 VTAIL.n63 VTAIL.n7 0.155672
R482 VTAIL.n64 VTAIL.n63 0.155672
R483 VTAIL.n64 VTAIL.n3 0.155672
R484 VTAIL.n71 VTAIL.n3 0.155672
R485 VTAIL.n221 VTAIL.n153 0.155672
R486 VTAIL.n214 VTAIL.n153 0.155672
R487 VTAIL.n214 VTAIL.n213 0.155672
R488 VTAIL.n213 VTAIL.n157 0.155672
R489 VTAIL.n206 VTAIL.n157 0.155672
R490 VTAIL.n206 VTAIL.n205 0.155672
R491 VTAIL.n205 VTAIL.n161 0.155672
R492 VTAIL.n198 VTAIL.n161 0.155672
R493 VTAIL.n198 VTAIL.n197 0.155672
R494 VTAIL.n197 VTAIL.n165 0.155672
R495 VTAIL.n190 VTAIL.n165 0.155672
R496 VTAIL.n190 VTAIL.n189 0.155672
R497 VTAIL.n189 VTAIL.n169 0.155672
R498 VTAIL.n182 VTAIL.n169 0.155672
R499 VTAIL.n182 VTAIL.n181 0.155672
R500 VTAIL.n181 VTAIL.n173 0.155672
R501 VTAIL.n147 VTAIL.n79 0.155672
R502 VTAIL.n140 VTAIL.n79 0.155672
R503 VTAIL.n140 VTAIL.n139 0.155672
R504 VTAIL.n139 VTAIL.n83 0.155672
R505 VTAIL.n132 VTAIL.n83 0.155672
R506 VTAIL.n132 VTAIL.n131 0.155672
R507 VTAIL.n131 VTAIL.n87 0.155672
R508 VTAIL.n124 VTAIL.n87 0.155672
R509 VTAIL.n124 VTAIL.n123 0.155672
R510 VTAIL.n123 VTAIL.n91 0.155672
R511 VTAIL.n116 VTAIL.n91 0.155672
R512 VTAIL.n116 VTAIL.n115 0.155672
R513 VTAIL.n115 VTAIL.n95 0.155672
R514 VTAIL.n108 VTAIL.n95 0.155672
R515 VTAIL.n108 VTAIL.n107 0.155672
R516 VTAIL.n107 VTAIL.n99 0.155672
R517 VDD2.n140 VDD2.n139 585
R518 VDD2.n138 VDD2.n137 585
R519 VDD2.n77 VDD2.n76 585
R520 VDD2.n132 VDD2.n131 585
R521 VDD2.n130 VDD2.n129 585
R522 VDD2.n81 VDD2.n80 585
R523 VDD2.n124 VDD2.n123 585
R524 VDD2.n122 VDD2.n121 585
R525 VDD2.n85 VDD2.n84 585
R526 VDD2.n116 VDD2.n115 585
R527 VDD2.n114 VDD2.n113 585
R528 VDD2.n89 VDD2.n88 585
R529 VDD2.n108 VDD2.n107 585
R530 VDD2.n106 VDD2.n105 585
R531 VDD2.n93 VDD2.n92 585
R532 VDD2.n100 VDD2.n99 585
R533 VDD2.n98 VDD2.n97 585
R534 VDD2.n25 VDD2.n24 585
R535 VDD2.n27 VDD2.n26 585
R536 VDD2.n20 VDD2.n19 585
R537 VDD2.n33 VDD2.n32 585
R538 VDD2.n35 VDD2.n34 585
R539 VDD2.n16 VDD2.n15 585
R540 VDD2.n41 VDD2.n40 585
R541 VDD2.n43 VDD2.n42 585
R542 VDD2.n12 VDD2.n11 585
R543 VDD2.n49 VDD2.n48 585
R544 VDD2.n51 VDD2.n50 585
R545 VDD2.n8 VDD2.n7 585
R546 VDD2.n57 VDD2.n56 585
R547 VDD2.n59 VDD2.n58 585
R548 VDD2.n4 VDD2.n3 585
R549 VDD2.n65 VDD2.n64 585
R550 VDD2.n67 VDD2.n66 585
R551 VDD2.n139 VDD2.n73 498.474
R552 VDD2.n66 VDD2.n0 498.474
R553 VDD2.n96 VDD2.t5 327.466
R554 VDD2.n23 VDD2.t0 327.466
R555 VDD2.n139 VDD2.n138 171.744
R556 VDD2.n138 VDD2.n76 171.744
R557 VDD2.n131 VDD2.n76 171.744
R558 VDD2.n131 VDD2.n130 171.744
R559 VDD2.n130 VDD2.n80 171.744
R560 VDD2.n123 VDD2.n80 171.744
R561 VDD2.n123 VDD2.n122 171.744
R562 VDD2.n122 VDD2.n84 171.744
R563 VDD2.n115 VDD2.n84 171.744
R564 VDD2.n115 VDD2.n114 171.744
R565 VDD2.n114 VDD2.n88 171.744
R566 VDD2.n107 VDD2.n88 171.744
R567 VDD2.n107 VDD2.n106 171.744
R568 VDD2.n106 VDD2.n92 171.744
R569 VDD2.n99 VDD2.n92 171.744
R570 VDD2.n99 VDD2.n98 171.744
R571 VDD2.n26 VDD2.n25 171.744
R572 VDD2.n26 VDD2.n19 171.744
R573 VDD2.n33 VDD2.n19 171.744
R574 VDD2.n34 VDD2.n33 171.744
R575 VDD2.n34 VDD2.n15 171.744
R576 VDD2.n41 VDD2.n15 171.744
R577 VDD2.n42 VDD2.n41 171.744
R578 VDD2.n42 VDD2.n11 171.744
R579 VDD2.n49 VDD2.n11 171.744
R580 VDD2.n50 VDD2.n49 171.744
R581 VDD2.n50 VDD2.n7 171.744
R582 VDD2.n57 VDD2.n7 171.744
R583 VDD2.n58 VDD2.n57 171.744
R584 VDD2.n58 VDD2.n3 171.744
R585 VDD2.n65 VDD2.n3 171.744
R586 VDD2.n66 VDD2.n65 171.744
R587 VDD2.n98 VDD2.t5 85.8723
R588 VDD2.n25 VDD2.t0 85.8723
R589 VDD2.n72 VDD2.n71 75.3655
R590 VDD2 VDD2.n145 75.3626
R591 VDD2.n72 VDD2.n70 54.1296
R592 VDD2.n144 VDD2.n143 51.3853
R593 VDD2.n144 VDD2.n72 47.3381
R594 VDD2.n97 VDD2.n96 16.3895
R595 VDD2.n24 VDD2.n23 16.3895
R596 VDD2.n141 VDD2.n140 12.8005
R597 VDD2.n100 VDD2.n95 12.8005
R598 VDD2.n27 VDD2.n22 12.8005
R599 VDD2.n68 VDD2.n67 12.8005
R600 VDD2.n137 VDD2.n75 12.0247
R601 VDD2.n101 VDD2.n93 12.0247
R602 VDD2.n28 VDD2.n20 12.0247
R603 VDD2.n64 VDD2.n2 12.0247
R604 VDD2.n136 VDD2.n77 11.249
R605 VDD2.n105 VDD2.n104 11.249
R606 VDD2.n32 VDD2.n31 11.249
R607 VDD2.n63 VDD2.n4 11.249
R608 VDD2.n133 VDD2.n132 10.4732
R609 VDD2.n108 VDD2.n91 10.4732
R610 VDD2.n35 VDD2.n18 10.4732
R611 VDD2.n60 VDD2.n59 10.4732
R612 VDD2.n129 VDD2.n79 9.69747
R613 VDD2.n109 VDD2.n89 9.69747
R614 VDD2.n36 VDD2.n16 9.69747
R615 VDD2.n56 VDD2.n6 9.69747
R616 VDD2.n143 VDD2.n142 9.45567
R617 VDD2.n70 VDD2.n69 9.45567
R618 VDD2.n83 VDD2.n82 9.3005
R619 VDD2.n126 VDD2.n125 9.3005
R620 VDD2.n128 VDD2.n127 9.3005
R621 VDD2.n79 VDD2.n78 9.3005
R622 VDD2.n134 VDD2.n133 9.3005
R623 VDD2.n136 VDD2.n135 9.3005
R624 VDD2.n75 VDD2.n74 9.3005
R625 VDD2.n142 VDD2.n141 9.3005
R626 VDD2.n120 VDD2.n119 9.3005
R627 VDD2.n118 VDD2.n117 9.3005
R628 VDD2.n87 VDD2.n86 9.3005
R629 VDD2.n112 VDD2.n111 9.3005
R630 VDD2.n110 VDD2.n109 9.3005
R631 VDD2.n91 VDD2.n90 9.3005
R632 VDD2.n104 VDD2.n103 9.3005
R633 VDD2.n102 VDD2.n101 9.3005
R634 VDD2.n95 VDD2.n94 9.3005
R635 VDD2.n45 VDD2.n44 9.3005
R636 VDD2.n14 VDD2.n13 9.3005
R637 VDD2.n39 VDD2.n38 9.3005
R638 VDD2.n37 VDD2.n36 9.3005
R639 VDD2.n18 VDD2.n17 9.3005
R640 VDD2.n31 VDD2.n30 9.3005
R641 VDD2.n29 VDD2.n28 9.3005
R642 VDD2.n22 VDD2.n21 9.3005
R643 VDD2.n47 VDD2.n46 9.3005
R644 VDD2.n10 VDD2.n9 9.3005
R645 VDD2.n53 VDD2.n52 9.3005
R646 VDD2.n55 VDD2.n54 9.3005
R647 VDD2.n6 VDD2.n5 9.3005
R648 VDD2.n61 VDD2.n60 9.3005
R649 VDD2.n63 VDD2.n62 9.3005
R650 VDD2.n2 VDD2.n1 9.3005
R651 VDD2.n69 VDD2.n68 9.3005
R652 VDD2.n128 VDD2.n81 8.92171
R653 VDD2.n113 VDD2.n112 8.92171
R654 VDD2.n40 VDD2.n39 8.92171
R655 VDD2.n55 VDD2.n8 8.92171
R656 VDD2.n125 VDD2.n124 8.14595
R657 VDD2.n116 VDD2.n87 8.14595
R658 VDD2.n43 VDD2.n14 8.14595
R659 VDD2.n52 VDD2.n51 8.14595
R660 VDD2.n143 VDD2.n73 7.75445
R661 VDD2.n70 VDD2.n0 7.75445
R662 VDD2.n121 VDD2.n83 7.3702
R663 VDD2.n117 VDD2.n85 7.3702
R664 VDD2.n44 VDD2.n12 7.3702
R665 VDD2.n48 VDD2.n10 7.3702
R666 VDD2.n121 VDD2.n120 6.59444
R667 VDD2.n120 VDD2.n85 6.59444
R668 VDD2.n47 VDD2.n12 6.59444
R669 VDD2.n48 VDD2.n47 6.59444
R670 VDD2.n141 VDD2.n73 6.08283
R671 VDD2.n68 VDD2.n0 6.08283
R672 VDD2.n124 VDD2.n83 5.81868
R673 VDD2.n117 VDD2.n116 5.81868
R674 VDD2.n44 VDD2.n43 5.81868
R675 VDD2.n51 VDD2.n10 5.81868
R676 VDD2.n125 VDD2.n81 5.04292
R677 VDD2.n113 VDD2.n87 5.04292
R678 VDD2.n40 VDD2.n14 5.04292
R679 VDD2.n52 VDD2.n8 5.04292
R680 VDD2.n129 VDD2.n128 4.26717
R681 VDD2.n112 VDD2.n89 4.26717
R682 VDD2.n39 VDD2.n16 4.26717
R683 VDD2.n56 VDD2.n55 4.26717
R684 VDD2.n96 VDD2.n94 3.70982
R685 VDD2.n23 VDD2.n21 3.70982
R686 VDD2.n132 VDD2.n79 3.49141
R687 VDD2.n109 VDD2.n108 3.49141
R688 VDD2.n36 VDD2.n35 3.49141
R689 VDD2.n59 VDD2.n6 3.49141
R690 VDD2 VDD2.n144 2.85826
R691 VDD2.n133 VDD2.n77 2.71565
R692 VDD2.n105 VDD2.n91 2.71565
R693 VDD2.n32 VDD2.n18 2.71565
R694 VDD2.n60 VDD2.n4 2.71565
R695 VDD2.n145 VDD2.t2 2.43898
R696 VDD2.n145 VDD2.t3 2.43898
R697 VDD2.n71 VDD2.t4 2.43898
R698 VDD2.n71 VDD2.t1 2.43898
R699 VDD2.n137 VDD2.n136 1.93989
R700 VDD2.n104 VDD2.n93 1.93989
R701 VDD2.n31 VDD2.n20 1.93989
R702 VDD2.n64 VDD2.n63 1.93989
R703 VDD2.n140 VDD2.n75 1.16414
R704 VDD2.n101 VDD2.n100 1.16414
R705 VDD2.n28 VDD2.n27 1.16414
R706 VDD2.n67 VDD2.n2 1.16414
R707 VDD2.n97 VDD2.n95 0.388379
R708 VDD2.n24 VDD2.n22 0.388379
R709 VDD2.n142 VDD2.n74 0.155672
R710 VDD2.n135 VDD2.n74 0.155672
R711 VDD2.n135 VDD2.n134 0.155672
R712 VDD2.n134 VDD2.n78 0.155672
R713 VDD2.n127 VDD2.n78 0.155672
R714 VDD2.n127 VDD2.n126 0.155672
R715 VDD2.n126 VDD2.n82 0.155672
R716 VDD2.n119 VDD2.n82 0.155672
R717 VDD2.n119 VDD2.n118 0.155672
R718 VDD2.n118 VDD2.n86 0.155672
R719 VDD2.n111 VDD2.n86 0.155672
R720 VDD2.n111 VDD2.n110 0.155672
R721 VDD2.n110 VDD2.n90 0.155672
R722 VDD2.n103 VDD2.n90 0.155672
R723 VDD2.n103 VDD2.n102 0.155672
R724 VDD2.n102 VDD2.n94 0.155672
R725 VDD2.n29 VDD2.n21 0.155672
R726 VDD2.n30 VDD2.n29 0.155672
R727 VDD2.n30 VDD2.n17 0.155672
R728 VDD2.n37 VDD2.n17 0.155672
R729 VDD2.n38 VDD2.n37 0.155672
R730 VDD2.n38 VDD2.n13 0.155672
R731 VDD2.n45 VDD2.n13 0.155672
R732 VDD2.n46 VDD2.n45 0.155672
R733 VDD2.n46 VDD2.n9 0.155672
R734 VDD2.n53 VDD2.n9 0.155672
R735 VDD2.n54 VDD2.n53 0.155672
R736 VDD2.n54 VDD2.n5 0.155672
R737 VDD2.n61 VDD2.n5 0.155672
R738 VDD2.n62 VDD2.n61 0.155672
R739 VDD2.n62 VDD2.n1 0.155672
R740 VDD2.n69 VDD2.n1 0.155672
R741 B.n650 B.n649 585
R742 B.n651 B.n86 585
R743 B.n653 B.n652 585
R744 B.n654 B.n85 585
R745 B.n656 B.n655 585
R746 B.n657 B.n84 585
R747 B.n659 B.n658 585
R748 B.n660 B.n83 585
R749 B.n662 B.n661 585
R750 B.n663 B.n82 585
R751 B.n665 B.n664 585
R752 B.n666 B.n81 585
R753 B.n668 B.n667 585
R754 B.n669 B.n80 585
R755 B.n671 B.n670 585
R756 B.n672 B.n79 585
R757 B.n674 B.n673 585
R758 B.n675 B.n78 585
R759 B.n677 B.n676 585
R760 B.n678 B.n77 585
R761 B.n680 B.n679 585
R762 B.n681 B.n76 585
R763 B.n683 B.n682 585
R764 B.n684 B.n75 585
R765 B.n686 B.n685 585
R766 B.n687 B.n74 585
R767 B.n689 B.n688 585
R768 B.n690 B.n73 585
R769 B.n692 B.n691 585
R770 B.n693 B.n72 585
R771 B.n695 B.n694 585
R772 B.n696 B.n71 585
R773 B.n698 B.n697 585
R774 B.n699 B.n70 585
R775 B.n701 B.n700 585
R776 B.n702 B.n69 585
R777 B.n704 B.n703 585
R778 B.n705 B.n68 585
R779 B.n707 B.n706 585
R780 B.n708 B.n67 585
R781 B.n710 B.n709 585
R782 B.n711 B.n66 585
R783 B.n713 B.n712 585
R784 B.n714 B.n65 585
R785 B.n716 B.n715 585
R786 B.n717 B.n62 585
R787 B.n720 B.n719 585
R788 B.n721 B.n61 585
R789 B.n723 B.n722 585
R790 B.n724 B.n60 585
R791 B.n726 B.n725 585
R792 B.n727 B.n59 585
R793 B.n729 B.n728 585
R794 B.n730 B.n55 585
R795 B.n732 B.n731 585
R796 B.n733 B.n54 585
R797 B.n735 B.n734 585
R798 B.n736 B.n53 585
R799 B.n738 B.n737 585
R800 B.n739 B.n52 585
R801 B.n741 B.n740 585
R802 B.n742 B.n51 585
R803 B.n744 B.n743 585
R804 B.n745 B.n50 585
R805 B.n747 B.n746 585
R806 B.n748 B.n49 585
R807 B.n750 B.n749 585
R808 B.n751 B.n48 585
R809 B.n753 B.n752 585
R810 B.n754 B.n47 585
R811 B.n756 B.n755 585
R812 B.n757 B.n46 585
R813 B.n759 B.n758 585
R814 B.n760 B.n45 585
R815 B.n762 B.n761 585
R816 B.n763 B.n44 585
R817 B.n765 B.n764 585
R818 B.n766 B.n43 585
R819 B.n768 B.n767 585
R820 B.n769 B.n42 585
R821 B.n771 B.n770 585
R822 B.n772 B.n41 585
R823 B.n774 B.n773 585
R824 B.n775 B.n40 585
R825 B.n777 B.n776 585
R826 B.n778 B.n39 585
R827 B.n780 B.n779 585
R828 B.n781 B.n38 585
R829 B.n783 B.n782 585
R830 B.n784 B.n37 585
R831 B.n786 B.n785 585
R832 B.n787 B.n36 585
R833 B.n789 B.n788 585
R834 B.n790 B.n35 585
R835 B.n792 B.n791 585
R836 B.n793 B.n34 585
R837 B.n795 B.n794 585
R838 B.n796 B.n33 585
R839 B.n798 B.n797 585
R840 B.n799 B.n32 585
R841 B.n801 B.n800 585
R842 B.n648 B.n87 585
R843 B.n647 B.n646 585
R844 B.n645 B.n88 585
R845 B.n644 B.n643 585
R846 B.n642 B.n89 585
R847 B.n641 B.n640 585
R848 B.n639 B.n90 585
R849 B.n638 B.n637 585
R850 B.n636 B.n91 585
R851 B.n635 B.n634 585
R852 B.n633 B.n92 585
R853 B.n632 B.n631 585
R854 B.n630 B.n93 585
R855 B.n629 B.n628 585
R856 B.n627 B.n94 585
R857 B.n626 B.n625 585
R858 B.n624 B.n95 585
R859 B.n623 B.n622 585
R860 B.n621 B.n96 585
R861 B.n620 B.n619 585
R862 B.n618 B.n97 585
R863 B.n617 B.n616 585
R864 B.n615 B.n98 585
R865 B.n614 B.n613 585
R866 B.n612 B.n99 585
R867 B.n611 B.n610 585
R868 B.n609 B.n100 585
R869 B.n608 B.n607 585
R870 B.n606 B.n101 585
R871 B.n605 B.n604 585
R872 B.n603 B.n102 585
R873 B.n602 B.n601 585
R874 B.n600 B.n103 585
R875 B.n599 B.n598 585
R876 B.n597 B.n104 585
R877 B.n596 B.n595 585
R878 B.n594 B.n105 585
R879 B.n593 B.n592 585
R880 B.n591 B.n106 585
R881 B.n590 B.n589 585
R882 B.n588 B.n107 585
R883 B.n587 B.n586 585
R884 B.n585 B.n108 585
R885 B.n584 B.n583 585
R886 B.n582 B.n109 585
R887 B.n581 B.n580 585
R888 B.n579 B.n110 585
R889 B.n578 B.n577 585
R890 B.n576 B.n111 585
R891 B.n575 B.n574 585
R892 B.n573 B.n112 585
R893 B.n572 B.n571 585
R894 B.n570 B.n113 585
R895 B.n569 B.n568 585
R896 B.n567 B.n114 585
R897 B.n566 B.n565 585
R898 B.n564 B.n115 585
R899 B.n563 B.n562 585
R900 B.n561 B.n116 585
R901 B.n560 B.n559 585
R902 B.n558 B.n117 585
R903 B.n557 B.n556 585
R904 B.n555 B.n118 585
R905 B.n554 B.n553 585
R906 B.n552 B.n119 585
R907 B.n551 B.n550 585
R908 B.n549 B.n120 585
R909 B.n548 B.n547 585
R910 B.n546 B.n121 585
R911 B.n545 B.n544 585
R912 B.n543 B.n122 585
R913 B.n542 B.n541 585
R914 B.n540 B.n123 585
R915 B.n539 B.n538 585
R916 B.n537 B.n124 585
R917 B.n536 B.n535 585
R918 B.n534 B.n125 585
R919 B.n533 B.n532 585
R920 B.n531 B.n126 585
R921 B.n530 B.n529 585
R922 B.n528 B.n127 585
R923 B.n527 B.n526 585
R924 B.n525 B.n128 585
R925 B.n524 B.n523 585
R926 B.n522 B.n129 585
R927 B.n521 B.n520 585
R928 B.n519 B.n130 585
R929 B.n518 B.n517 585
R930 B.n516 B.n131 585
R931 B.n515 B.n514 585
R932 B.n513 B.n132 585
R933 B.n512 B.n511 585
R934 B.n510 B.n133 585
R935 B.n509 B.n508 585
R936 B.n507 B.n134 585
R937 B.n506 B.n505 585
R938 B.n504 B.n135 585
R939 B.n503 B.n502 585
R940 B.n501 B.n136 585
R941 B.n500 B.n499 585
R942 B.n498 B.n137 585
R943 B.n497 B.n496 585
R944 B.n495 B.n138 585
R945 B.n494 B.n493 585
R946 B.n492 B.n139 585
R947 B.n491 B.n490 585
R948 B.n489 B.n140 585
R949 B.n488 B.n487 585
R950 B.n486 B.n141 585
R951 B.n485 B.n484 585
R952 B.n483 B.n142 585
R953 B.n482 B.n481 585
R954 B.n480 B.n143 585
R955 B.n479 B.n478 585
R956 B.n477 B.n144 585
R957 B.n476 B.n475 585
R958 B.n474 B.n145 585
R959 B.n473 B.n472 585
R960 B.n471 B.n146 585
R961 B.n316 B.n315 585
R962 B.n317 B.n198 585
R963 B.n319 B.n318 585
R964 B.n320 B.n197 585
R965 B.n322 B.n321 585
R966 B.n323 B.n196 585
R967 B.n325 B.n324 585
R968 B.n326 B.n195 585
R969 B.n328 B.n327 585
R970 B.n329 B.n194 585
R971 B.n331 B.n330 585
R972 B.n332 B.n193 585
R973 B.n334 B.n333 585
R974 B.n335 B.n192 585
R975 B.n337 B.n336 585
R976 B.n338 B.n191 585
R977 B.n340 B.n339 585
R978 B.n341 B.n190 585
R979 B.n343 B.n342 585
R980 B.n344 B.n189 585
R981 B.n346 B.n345 585
R982 B.n347 B.n188 585
R983 B.n349 B.n348 585
R984 B.n350 B.n187 585
R985 B.n352 B.n351 585
R986 B.n353 B.n186 585
R987 B.n355 B.n354 585
R988 B.n356 B.n185 585
R989 B.n358 B.n357 585
R990 B.n359 B.n184 585
R991 B.n361 B.n360 585
R992 B.n362 B.n183 585
R993 B.n364 B.n363 585
R994 B.n365 B.n182 585
R995 B.n367 B.n366 585
R996 B.n368 B.n181 585
R997 B.n370 B.n369 585
R998 B.n371 B.n180 585
R999 B.n373 B.n372 585
R1000 B.n374 B.n179 585
R1001 B.n376 B.n375 585
R1002 B.n377 B.n178 585
R1003 B.n379 B.n378 585
R1004 B.n380 B.n177 585
R1005 B.n382 B.n381 585
R1006 B.n383 B.n174 585
R1007 B.n386 B.n385 585
R1008 B.n387 B.n173 585
R1009 B.n389 B.n388 585
R1010 B.n390 B.n172 585
R1011 B.n392 B.n391 585
R1012 B.n393 B.n171 585
R1013 B.n395 B.n394 585
R1014 B.n396 B.n170 585
R1015 B.n401 B.n400 585
R1016 B.n402 B.n169 585
R1017 B.n404 B.n403 585
R1018 B.n405 B.n168 585
R1019 B.n407 B.n406 585
R1020 B.n408 B.n167 585
R1021 B.n410 B.n409 585
R1022 B.n411 B.n166 585
R1023 B.n413 B.n412 585
R1024 B.n414 B.n165 585
R1025 B.n416 B.n415 585
R1026 B.n417 B.n164 585
R1027 B.n419 B.n418 585
R1028 B.n420 B.n163 585
R1029 B.n422 B.n421 585
R1030 B.n423 B.n162 585
R1031 B.n425 B.n424 585
R1032 B.n426 B.n161 585
R1033 B.n428 B.n427 585
R1034 B.n429 B.n160 585
R1035 B.n431 B.n430 585
R1036 B.n432 B.n159 585
R1037 B.n434 B.n433 585
R1038 B.n435 B.n158 585
R1039 B.n437 B.n436 585
R1040 B.n438 B.n157 585
R1041 B.n440 B.n439 585
R1042 B.n441 B.n156 585
R1043 B.n443 B.n442 585
R1044 B.n444 B.n155 585
R1045 B.n446 B.n445 585
R1046 B.n447 B.n154 585
R1047 B.n449 B.n448 585
R1048 B.n450 B.n153 585
R1049 B.n452 B.n451 585
R1050 B.n453 B.n152 585
R1051 B.n455 B.n454 585
R1052 B.n456 B.n151 585
R1053 B.n458 B.n457 585
R1054 B.n459 B.n150 585
R1055 B.n461 B.n460 585
R1056 B.n462 B.n149 585
R1057 B.n464 B.n463 585
R1058 B.n465 B.n148 585
R1059 B.n467 B.n466 585
R1060 B.n468 B.n147 585
R1061 B.n470 B.n469 585
R1062 B.n314 B.n199 585
R1063 B.n313 B.n312 585
R1064 B.n311 B.n200 585
R1065 B.n310 B.n309 585
R1066 B.n308 B.n201 585
R1067 B.n307 B.n306 585
R1068 B.n305 B.n202 585
R1069 B.n304 B.n303 585
R1070 B.n302 B.n203 585
R1071 B.n301 B.n300 585
R1072 B.n299 B.n204 585
R1073 B.n298 B.n297 585
R1074 B.n296 B.n205 585
R1075 B.n295 B.n294 585
R1076 B.n293 B.n206 585
R1077 B.n292 B.n291 585
R1078 B.n290 B.n207 585
R1079 B.n289 B.n288 585
R1080 B.n287 B.n208 585
R1081 B.n286 B.n285 585
R1082 B.n284 B.n209 585
R1083 B.n283 B.n282 585
R1084 B.n281 B.n210 585
R1085 B.n280 B.n279 585
R1086 B.n278 B.n211 585
R1087 B.n277 B.n276 585
R1088 B.n275 B.n212 585
R1089 B.n274 B.n273 585
R1090 B.n272 B.n213 585
R1091 B.n271 B.n270 585
R1092 B.n269 B.n214 585
R1093 B.n268 B.n267 585
R1094 B.n266 B.n215 585
R1095 B.n265 B.n264 585
R1096 B.n263 B.n216 585
R1097 B.n262 B.n261 585
R1098 B.n260 B.n217 585
R1099 B.n259 B.n258 585
R1100 B.n257 B.n218 585
R1101 B.n256 B.n255 585
R1102 B.n254 B.n219 585
R1103 B.n253 B.n252 585
R1104 B.n251 B.n220 585
R1105 B.n250 B.n249 585
R1106 B.n248 B.n221 585
R1107 B.n247 B.n246 585
R1108 B.n245 B.n222 585
R1109 B.n244 B.n243 585
R1110 B.n242 B.n223 585
R1111 B.n241 B.n240 585
R1112 B.n239 B.n224 585
R1113 B.n238 B.n237 585
R1114 B.n236 B.n225 585
R1115 B.n235 B.n234 585
R1116 B.n233 B.n226 585
R1117 B.n232 B.n231 585
R1118 B.n230 B.n227 585
R1119 B.n229 B.n228 585
R1120 B.n2 B.n0 585
R1121 B.n889 B.n1 585
R1122 B.n888 B.n887 585
R1123 B.n886 B.n3 585
R1124 B.n885 B.n884 585
R1125 B.n883 B.n4 585
R1126 B.n882 B.n881 585
R1127 B.n880 B.n5 585
R1128 B.n879 B.n878 585
R1129 B.n877 B.n6 585
R1130 B.n876 B.n875 585
R1131 B.n874 B.n7 585
R1132 B.n873 B.n872 585
R1133 B.n871 B.n8 585
R1134 B.n870 B.n869 585
R1135 B.n868 B.n9 585
R1136 B.n867 B.n866 585
R1137 B.n865 B.n10 585
R1138 B.n864 B.n863 585
R1139 B.n862 B.n11 585
R1140 B.n861 B.n860 585
R1141 B.n859 B.n12 585
R1142 B.n858 B.n857 585
R1143 B.n856 B.n13 585
R1144 B.n855 B.n854 585
R1145 B.n853 B.n14 585
R1146 B.n852 B.n851 585
R1147 B.n850 B.n15 585
R1148 B.n849 B.n848 585
R1149 B.n847 B.n16 585
R1150 B.n846 B.n845 585
R1151 B.n844 B.n17 585
R1152 B.n843 B.n842 585
R1153 B.n841 B.n18 585
R1154 B.n840 B.n839 585
R1155 B.n838 B.n19 585
R1156 B.n837 B.n836 585
R1157 B.n835 B.n20 585
R1158 B.n834 B.n833 585
R1159 B.n832 B.n21 585
R1160 B.n831 B.n830 585
R1161 B.n829 B.n22 585
R1162 B.n828 B.n827 585
R1163 B.n826 B.n23 585
R1164 B.n825 B.n824 585
R1165 B.n823 B.n24 585
R1166 B.n822 B.n821 585
R1167 B.n820 B.n25 585
R1168 B.n819 B.n818 585
R1169 B.n817 B.n26 585
R1170 B.n816 B.n815 585
R1171 B.n814 B.n27 585
R1172 B.n813 B.n812 585
R1173 B.n811 B.n28 585
R1174 B.n810 B.n809 585
R1175 B.n808 B.n29 585
R1176 B.n807 B.n806 585
R1177 B.n805 B.n30 585
R1178 B.n804 B.n803 585
R1179 B.n802 B.n31 585
R1180 B.n891 B.n890 585
R1181 B.n397 B.t8 483.418
R1182 B.n63 B.t10 483.418
R1183 B.n175 B.t5 483.418
R1184 B.n56 B.t1 483.418
R1185 B.n315 B.n314 478.086
R1186 B.n800 B.n31 478.086
R1187 B.n469 B.n146 478.086
R1188 B.n649 B.n648 478.086
R1189 B.n398 B.t7 399.442
R1190 B.n64 B.t11 399.442
R1191 B.n176 B.t4 399.442
R1192 B.n57 B.t2 399.442
R1193 B.n397 B.t6 289.805
R1194 B.n175 B.t3 289.805
R1195 B.n56 B.t0 289.805
R1196 B.n63 B.t9 289.805
R1197 B.n314 B.n313 163.367
R1198 B.n313 B.n200 163.367
R1199 B.n309 B.n200 163.367
R1200 B.n309 B.n308 163.367
R1201 B.n308 B.n307 163.367
R1202 B.n307 B.n202 163.367
R1203 B.n303 B.n202 163.367
R1204 B.n303 B.n302 163.367
R1205 B.n302 B.n301 163.367
R1206 B.n301 B.n204 163.367
R1207 B.n297 B.n204 163.367
R1208 B.n297 B.n296 163.367
R1209 B.n296 B.n295 163.367
R1210 B.n295 B.n206 163.367
R1211 B.n291 B.n206 163.367
R1212 B.n291 B.n290 163.367
R1213 B.n290 B.n289 163.367
R1214 B.n289 B.n208 163.367
R1215 B.n285 B.n208 163.367
R1216 B.n285 B.n284 163.367
R1217 B.n284 B.n283 163.367
R1218 B.n283 B.n210 163.367
R1219 B.n279 B.n210 163.367
R1220 B.n279 B.n278 163.367
R1221 B.n278 B.n277 163.367
R1222 B.n277 B.n212 163.367
R1223 B.n273 B.n212 163.367
R1224 B.n273 B.n272 163.367
R1225 B.n272 B.n271 163.367
R1226 B.n271 B.n214 163.367
R1227 B.n267 B.n214 163.367
R1228 B.n267 B.n266 163.367
R1229 B.n266 B.n265 163.367
R1230 B.n265 B.n216 163.367
R1231 B.n261 B.n216 163.367
R1232 B.n261 B.n260 163.367
R1233 B.n260 B.n259 163.367
R1234 B.n259 B.n218 163.367
R1235 B.n255 B.n218 163.367
R1236 B.n255 B.n254 163.367
R1237 B.n254 B.n253 163.367
R1238 B.n253 B.n220 163.367
R1239 B.n249 B.n220 163.367
R1240 B.n249 B.n248 163.367
R1241 B.n248 B.n247 163.367
R1242 B.n247 B.n222 163.367
R1243 B.n243 B.n222 163.367
R1244 B.n243 B.n242 163.367
R1245 B.n242 B.n241 163.367
R1246 B.n241 B.n224 163.367
R1247 B.n237 B.n224 163.367
R1248 B.n237 B.n236 163.367
R1249 B.n236 B.n235 163.367
R1250 B.n235 B.n226 163.367
R1251 B.n231 B.n226 163.367
R1252 B.n231 B.n230 163.367
R1253 B.n230 B.n229 163.367
R1254 B.n229 B.n2 163.367
R1255 B.n890 B.n2 163.367
R1256 B.n890 B.n889 163.367
R1257 B.n889 B.n888 163.367
R1258 B.n888 B.n3 163.367
R1259 B.n884 B.n3 163.367
R1260 B.n884 B.n883 163.367
R1261 B.n883 B.n882 163.367
R1262 B.n882 B.n5 163.367
R1263 B.n878 B.n5 163.367
R1264 B.n878 B.n877 163.367
R1265 B.n877 B.n876 163.367
R1266 B.n876 B.n7 163.367
R1267 B.n872 B.n7 163.367
R1268 B.n872 B.n871 163.367
R1269 B.n871 B.n870 163.367
R1270 B.n870 B.n9 163.367
R1271 B.n866 B.n9 163.367
R1272 B.n866 B.n865 163.367
R1273 B.n865 B.n864 163.367
R1274 B.n864 B.n11 163.367
R1275 B.n860 B.n11 163.367
R1276 B.n860 B.n859 163.367
R1277 B.n859 B.n858 163.367
R1278 B.n858 B.n13 163.367
R1279 B.n854 B.n13 163.367
R1280 B.n854 B.n853 163.367
R1281 B.n853 B.n852 163.367
R1282 B.n852 B.n15 163.367
R1283 B.n848 B.n15 163.367
R1284 B.n848 B.n847 163.367
R1285 B.n847 B.n846 163.367
R1286 B.n846 B.n17 163.367
R1287 B.n842 B.n17 163.367
R1288 B.n842 B.n841 163.367
R1289 B.n841 B.n840 163.367
R1290 B.n840 B.n19 163.367
R1291 B.n836 B.n19 163.367
R1292 B.n836 B.n835 163.367
R1293 B.n835 B.n834 163.367
R1294 B.n834 B.n21 163.367
R1295 B.n830 B.n21 163.367
R1296 B.n830 B.n829 163.367
R1297 B.n829 B.n828 163.367
R1298 B.n828 B.n23 163.367
R1299 B.n824 B.n23 163.367
R1300 B.n824 B.n823 163.367
R1301 B.n823 B.n822 163.367
R1302 B.n822 B.n25 163.367
R1303 B.n818 B.n25 163.367
R1304 B.n818 B.n817 163.367
R1305 B.n817 B.n816 163.367
R1306 B.n816 B.n27 163.367
R1307 B.n812 B.n27 163.367
R1308 B.n812 B.n811 163.367
R1309 B.n811 B.n810 163.367
R1310 B.n810 B.n29 163.367
R1311 B.n806 B.n29 163.367
R1312 B.n806 B.n805 163.367
R1313 B.n805 B.n804 163.367
R1314 B.n804 B.n31 163.367
R1315 B.n315 B.n198 163.367
R1316 B.n319 B.n198 163.367
R1317 B.n320 B.n319 163.367
R1318 B.n321 B.n320 163.367
R1319 B.n321 B.n196 163.367
R1320 B.n325 B.n196 163.367
R1321 B.n326 B.n325 163.367
R1322 B.n327 B.n326 163.367
R1323 B.n327 B.n194 163.367
R1324 B.n331 B.n194 163.367
R1325 B.n332 B.n331 163.367
R1326 B.n333 B.n332 163.367
R1327 B.n333 B.n192 163.367
R1328 B.n337 B.n192 163.367
R1329 B.n338 B.n337 163.367
R1330 B.n339 B.n338 163.367
R1331 B.n339 B.n190 163.367
R1332 B.n343 B.n190 163.367
R1333 B.n344 B.n343 163.367
R1334 B.n345 B.n344 163.367
R1335 B.n345 B.n188 163.367
R1336 B.n349 B.n188 163.367
R1337 B.n350 B.n349 163.367
R1338 B.n351 B.n350 163.367
R1339 B.n351 B.n186 163.367
R1340 B.n355 B.n186 163.367
R1341 B.n356 B.n355 163.367
R1342 B.n357 B.n356 163.367
R1343 B.n357 B.n184 163.367
R1344 B.n361 B.n184 163.367
R1345 B.n362 B.n361 163.367
R1346 B.n363 B.n362 163.367
R1347 B.n363 B.n182 163.367
R1348 B.n367 B.n182 163.367
R1349 B.n368 B.n367 163.367
R1350 B.n369 B.n368 163.367
R1351 B.n369 B.n180 163.367
R1352 B.n373 B.n180 163.367
R1353 B.n374 B.n373 163.367
R1354 B.n375 B.n374 163.367
R1355 B.n375 B.n178 163.367
R1356 B.n379 B.n178 163.367
R1357 B.n380 B.n379 163.367
R1358 B.n381 B.n380 163.367
R1359 B.n381 B.n174 163.367
R1360 B.n386 B.n174 163.367
R1361 B.n387 B.n386 163.367
R1362 B.n388 B.n387 163.367
R1363 B.n388 B.n172 163.367
R1364 B.n392 B.n172 163.367
R1365 B.n393 B.n392 163.367
R1366 B.n394 B.n393 163.367
R1367 B.n394 B.n170 163.367
R1368 B.n401 B.n170 163.367
R1369 B.n402 B.n401 163.367
R1370 B.n403 B.n402 163.367
R1371 B.n403 B.n168 163.367
R1372 B.n407 B.n168 163.367
R1373 B.n408 B.n407 163.367
R1374 B.n409 B.n408 163.367
R1375 B.n409 B.n166 163.367
R1376 B.n413 B.n166 163.367
R1377 B.n414 B.n413 163.367
R1378 B.n415 B.n414 163.367
R1379 B.n415 B.n164 163.367
R1380 B.n419 B.n164 163.367
R1381 B.n420 B.n419 163.367
R1382 B.n421 B.n420 163.367
R1383 B.n421 B.n162 163.367
R1384 B.n425 B.n162 163.367
R1385 B.n426 B.n425 163.367
R1386 B.n427 B.n426 163.367
R1387 B.n427 B.n160 163.367
R1388 B.n431 B.n160 163.367
R1389 B.n432 B.n431 163.367
R1390 B.n433 B.n432 163.367
R1391 B.n433 B.n158 163.367
R1392 B.n437 B.n158 163.367
R1393 B.n438 B.n437 163.367
R1394 B.n439 B.n438 163.367
R1395 B.n439 B.n156 163.367
R1396 B.n443 B.n156 163.367
R1397 B.n444 B.n443 163.367
R1398 B.n445 B.n444 163.367
R1399 B.n445 B.n154 163.367
R1400 B.n449 B.n154 163.367
R1401 B.n450 B.n449 163.367
R1402 B.n451 B.n450 163.367
R1403 B.n451 B.n152 163.367
R1404 B.n455 B.n152 163.367
R1405 B.n456 B.n455 163.367
R1406 B.n457 B.n456 163.367
R1407 B.n457 B.n150 163.367
R1408 B.n461 B.n150 163.367
R1409 B.n462 B.n461 163.367
R1410 B.n463 B.n462 163.367
R1411 B.n463 B.n148 163.367
R1412 B.n467 B.n148 163.367
R1413 B.n468 B.n467 163.367
R1414 B.n469 B.n468 163.367
R1415 B.n473 B.n146 163.367
R1416 B.n474 B.n473 163.367
R1417 B.n475 B.n474 163.367
R1418 B.n475 B.n144 163.367
R1419 B.n479 B.n144 163.367
R1420 B.n480 B.n479 163.367
R1421 B.n481 B.n480 163.367
R1422 B.n481 B.n142 163.367
R1423 B.n485 B.n142 163.367
R1424 B.n486 B.n485 163.367
R1425 B.n487 B.n486 163.367
R1426 B.n487 B.n140 163.367
R1427 B.n491 B.n140 163.367
R1428 B.n492 B.n491 163.367
R1429 B.n493 B.n492 163.367
R1430 B.n493 B.n138 163.367
R1431 B.n497 B.n138 163.367
R1432 B.n498 B.n497 163.367
R1433 B.n499 B.n498 163.367
R1434 B.n499 B.n136 163.367
R1435 B.n503 B.n136 163.367
R1436 B.n504 B.n503 163.367
R1437 B.n505 B.n504 163.367
R1438 B.n505 B.n134 163.367
R1439 B.n509 B.n134 163.367
R1440 B.n510 B.n509 163.367
R1441 B.n511 B.n510 163.367
R1442 B.n511 B.n132 163.367
R1443 B.n515 B.n132 163.367
R1444 B.n516 B.n515 163.367
R1445 B.n517 B.n516 163.367
R1446 B.n517 B.n130 163.367
R1447 B.n521 B.n130 163.367
R1448 B.n522 B.n521 163.367
R1449 B.n523 B.n522 163.367
R1450 B.n523 B.n128 163.367
R1451 B.n527 B.n128 163.367
R1452 B.n528 B.n527 163.367
R1453 B.n529 B.n528 163.367
R1454 B.n529 B.n126 163.367
R1455 B.n533 B.n126 163.367
R1456 B.n534 B.n533 163.367
R1457 B.n535 B.n534 163.367
R1458 B.n535 B.n124 163.367
R1459 B.n539 B.n124 163.367
R1460 B.n540 B.n539 163.367
R1461 B.n541 B.n540 163.367
R1462 B.n541 B.n122 163.367
R1463 B.n545 B.n122 163.367
R1464 B.n546 B.n545 163.367
R1465 B.n547 B.n546 163.367
R1466 B.n547 B.n120 163.367
R1467 B.n551 B.n120 163.367
R1468 B.n552 B.n551 163.367
R1469 B.n553 B.n552 163.367
R1470 B.n553 B.n118 163.367
R1471 B.n557 B.n118 163.367
R1472 B.n558 B.n557 163.367
R1473 B.n559 B.n558 163.367
R1474 B.n559 B.n116 163.367
R1475 B.n563 B.n116 163.367
R1476 B.n564 B.n563 163.367
R1477 B.n565 B.n564 163.367
R1478 B.n565 B.n114 163.367
R1479 B.n569 B.n114 163.367
R1480 B.n570 B.n569 163.367
R1481 B.n571 B.n570 163.367
R1482 B.n571 B.n112 163.367
R1483 B.n575 B.n112 163.367
R1484 B.n576 B.n575 163.367
R1485 B.n577 B.n576 163.367
R1486 B.n577 B.n110 163.367
R1487 B.n581 B.n110 163.367
R1488 B.n582 B.n581 163.367
R1489 B.n583 B.n582 163.367
R1490 B.n583 B.n108 163.367
R1491 B.n587 B.n108 163.367
R1492 B.n588 B.n587 163.367
R1493 B.n589 B.n588 163.367
R1494 B.n589 B.n106 163.367
R1495 B.n593 B.n106 163.367
R1496 B.n594 B.n593 163.367
R1497 B.n595 B.n594 163.367
R1498 B.n595 B.n104 163.367
R1499 B.n599 B.n104 163.367
R1500 B.n600 B.n599 163.367
R1501 B.n601 B.n600 163.367
R1502 B.n601 B.n102 163.367
R1503 B.n605 B.n102 163.367
R1504 B.n606 B.n605 163.367
R1505 B.n607 B.n606 163.367
R1506 B.n607 B.n100 163.367
R1507 B.n611 B.n100 163.367
R1508 B.n612 B.n611 163.367
R1509 B.n613 B.n612 163.367
R1510 B.n613 B.n98 163.367
R1511 B.n617 B.n98 163.367
R1512 B.n618 B.n617 163.367
R1513 B.n619 B.n618 163.367
R1514 B.n619 B.n96 163.367
R1515 B.n623 B.n96 163.367
R1516 B.n624 B.n623 163.367
R1517 B.n625 B.n624 163.367
R1518 B.n625 B.n94 163.367
R1519 B.n629 B.n94 163.367
R1520 B.n630 B.n629 163.367
R1521 B.n631 B.n630 163.367
R1522 B.n631 B.n92 163.367
R1523 B.n635 B.n92 163.367
R1524 B.n636 B.n635 163.367
R1525 B.n637 B.n636 163.367
R1526 B.n637 B.n90 163.367
R1527 B.n641 B.n90 163.367
R1528 B.n642 B.n641 163.367
R1529 B.n643 B.n642 163.367
R1530 B.n643 B.n88 163.367
R1531 B.n647 B.n88 163.367
R1532 B.n648 B.n647 163.367
R1533 B.n800 B.n799 163.367
R1534 B.n799 B.n798 163.367
R1535 B.n798 B.n33 163.367
R1536 B.n794 B.n33 163.367
R1537 B.n794 B.n793 163.367
R1538 B.n793 B.n792 163.367
R1539 B.n792 B.n35 163.367
R1540 B.n788 B.n35 163.367
R1541 B.n788 B.n787 163.367
R1542 B.n787 B.n786 163.367
R1543 B.n786 B.n37 163.367
R1544 B.n782 B.n37 163.367
R1545 B.n782 B.n781 163.367
R1546 B.n781 B.n780 163.367
R1547 B.n780 B.n39 163.367
R1548 B.n776 B.n39 163.367
R1549 B.n776 B.n775 163.367
R1550 B.n775 B.n774 163.367
R1551 B.n774 B.n41 163.367
R1552 B.n770 B.n41 163.367
R1553 B.n770 B.n769 163.367
R1554 B.n769 B.n768 163.367
R1555 B.n768 B.n43 163.367
R1556 B.n764 B.n43 163.367
R1557 B.n764 B.n763 163.367
R1558 B.n763 B.n762 163.367
R1559 B.n762 B.n45 163.367
R1560 B.n758 B.n45 163.367
R1561 B.n758 B.n757 163.367
R1562 B.n757 B.n756 163.367
R1563 B.n756 B.n47 163.367
R1564 B.n752 B.n47 163.367
R1565 B.n752 B.n751 163.367
R1566 B.n751 B.n750 163.367
R1567 B.n750 B.n49 163.367
R1568 B.n746 B.n49 163.367
R1569 B.n746 B.n745 163.367
R1570 B.n745 B.n744 163.367
R1571 B.n744 B.n51 163.367
R1572 B.n740 B.n51 163.367
R1573 B.n740 B.n739 163.367
R1574 B.n739 B.n738 163.367
R1575 B.n738 B.n53 163.367
R1576 B.n734 B.n53 163.367
R1577 B.n734 B.n733 163.367
R1578 B.n733 B.n732 163.367
R1579 B.n732 B.n55 163.367
R1580 B.n728 B.n55 163.367
R1581 B.n728 B.n727 163.367
R1582 B.n727 B.n726 163.367
R1583 B.n726 B.n60 163.367
R1584 B.n722 B.n60 163.367
R1585 B.n722 B.n721 163.367
R1586 B.n721 B.n720 163.367
R1587 B.n720 B.n62 163.367
R1588 B.n715 B.n62 163.367
R1589 B.n715 B.n714 163.367
R1590 B.n714 B.n713 163.367
R1591 B.n713 B.n66 163.367
R1592 B.n709 B.n66 163.367
R1593 B.n709 B.n708 163.367
R1594 B.n708 B.n707 163.367
R1595 B.n707 B.n68 163.367
R1596 B.n703 B.n68 163.367
R1597 B.n703 B.n702 163.367
R1598 B.n702 B.n701 163.367
R1599 B.n701 B.n70 163.367
R1600 B.n697 B.n70 163.367
R1601 B.n697 B.n696 163.367
R1602 B.n696 B.n695 163.367
R1603 B.n695 B.n72 163.367
R1604 B.n691 B.n72 163.367
R1605 B.n691 B.n690 163.367
R1606 B.n690 B.n689 163.367
R1607 B.n689 B.n74 163.367
R1608 B.n685 B.n74 163.367
R1609 B.n685 B.n684 163.367
R1610 B.n684 B.n683 163.367
R1611 B.n683 B.n76 163.367
R1612 B.n679 B.n76 163.367
R1613 B.n679 B.n678 163.367
R1614 B.n678 B.n677 163.367
R1615 B.n677 B.n78 163.367
R1616 B.n673 B.n78 163.367
R1617 B.n673 B.n672 163.367
R1618 B.n672 B.n671 163.367
R1619 B.n671 B.n80 163.367
R1620 B.n667 B.n80 163.367
R1621 B.n667 B.n666 163.367
R1622 B.n666 B.n665 163.367
R1623 B.n665 B.n82 163.367
R1624 B.n661 B.n82 163.367
R1625 B.n661 B.n660 163.367
R1626 B.n660 B.n659 163.367
R1627 B.n659 B.n84 163.367
R1628 B.n655 B.n84 163.367
R1629 B.n655 B.n654 163.367
R1630 B.n654 B.n653 163.367
R1631 B.n653 B.n86 163.367
R1632 B.n649 B.n86 163.367
R1633 B.n398 B.n397 83.9763
R1634 B.n176 B.n175 83.9763
R1635 B.n57 B.n56 83.9763
R1636 B.n64 B.n63 83.9763
R1637 B.n399 B.n398 59.5399
R1638 B.n384 B.n176 59.5399
R1639 B.n58 B.n57 59.5399
R1640 B.n718 B.n64 59.5399
R1641 B.n802 B.n801 31.0639
R1642 B.n650 B.n87 31.0639
R1643 B.n471 B.n470 31.0639
R1644 B.n316 B.n199 31.0639
R1645 B B.n891 18.0485
R1646 B.n801 B.n32 10.6151
R1647 B.n797 B.n32 10.6151
R1648 B.n797 B.n796 10.6151
R1649 B.n796 B.n795 10.6151
R1650 B.n795 B.n34 10.6151
R1651 B.n791 B.n34 10.6151
R1652 B.n791 B.n790 10.6151
R1653 B.n790 B.n789 10.6151
R1654 B.n789 B.n36 10.6151
R1655 B.n785 B.n36 10.6151
R1656 B.n785 B.n784 10.6151
R1657 B.n784 B.n783 10.6151
R1658 B.n783 B.n38 10.6151
R1659 B.n779 B.n38 10.6151
R1660 B.n779 B.n778 10.6151
R1661 B.n778 B.n777 10.6151
R1662 B.n777 B.n40 10.6151
R1663 B.n773 B.n40 10.6151
R1664 B.n773 B.n772 10.6151
R1665 B.n772 B.n771 10.6151
R1666 B.n771 B.n42 10.6151
R1667 B.n767 B.n42 10.6151
R1668 B.n767 B.n766 10.6151
R1669 B.n766 B.n765 10.6151
R1670 B.n765 B.n44 10.6151
R1671 B.n761 B.n44 10.6151
R1672 B.n761 B.n760 10.6151
R1673 B.n760 B.n759 10.6151
R1674 B.n759 B.n46 10.6151
R1675 B.n755 B.n46 10.6151
R1676 B.n755 B.n754 10.6151
R1677 B.n754 B.n753 10.6151
R1678 B.n753 B.n48 10.6151
R1679 B.n749 B.n48 10.6151
R1680 B.n749 B.n748 10.6151
R1681 B.n748 B.n747 10.6151
R1682 B.n747 B.n50 10.6151
R1683 B.n743 B.n50 10.6151
R1684 B.n743 B.n742 10.6151
R1685 B.n742 B.n741 10.6151
R1686 B.n741 B.n52 10.6151
R1687 B.n737 B.n52 10.6151
R1688 B.n737 B.n736 10.6151
R1689 B.n736 B.n735 10.6151
R1690 B.n735 B.n54 10.6151
R1691 B.n731 B.n730 10.6151
R1692 B.n730 B.n729 10.6151
R1693 B.n729 B.n59 10.6151
R1694 B.n725 B.n59 10.6151
R1695 B.n725 B.n724 10.6151
R1696 B.n724 B.n723 10.6151
R1697 B.n723 B.n61 10.6151
R1698 B.n719 B.n61 10.6151
R1699 B.n717 B.n716 10.6151
R1700 B.n716 B.n65 10.6151
R1701 B.n712 B.n65 10.6151
R1702 B.n712 B.n711 10.6151
R1703 B.n711 B.n710 10.6151
R1704 B.n710 B.n67 10.6151
R1705 B.n706 B.n67 10.6151
R1706 B.n706 B.n705 10.6151
R1707 B.n705 B.n704 10.6151
R1708 B.n704 B.n69 10.6151
R1709 B.n700 B.n69 10.6151
R1710 B.n700 B.n699 10.6151
R1711 B.n699 B.n698 10.6151
R1712 B.n698 B.n71 10.6151
R1713 B.n694 B.n71 10.6151
R1714 B.n694 B.n693 10.6151
R1715 B.n693 B.n692 10.6151
R1716 B.n692 B.n73 10.6151
R1717 B.n688 B.n73 10.6151
R1718 B.n688 B.n687 10.6151
R1719 B.n687 B.n686 10.6151
R1720 B.n686 B.n75 10.6151
R1721 B.n682 B.n75 10.6151
R1722 B.n682 B.n681 10.6151
R1723 B.n681 B.n680 10.6151
R1724 B.n680 B.n77 10.6151
R1725 B.n676 B.n77 10.6151
R1726 B.n676 B.n675 10.6151
R1727 B.n675 B.n674 10.6151
R1728 B.n674 B.n79 10.6151
R1729 B.n670 B.n79 10.6151
R1730 B.n670 B.n669 10.6151
R1731 B.n669 B.n668 10.6151
R1732 B.n668 B.n81 10.6151
R1733 B.n664 B.n81 10.6151
R1734 B.n664 B.n663 10.6151
R1735 B.n663 B.n662 10.6151
R1736 B.n662 B.n83 10.6151
R1737 B.n658 B.n83 10.6151
R1738 B.n658 B.n657 10.6151
R1739 B.n657 B.n656 10.6151
R1740 B.n656 B.n85 10.6151
R1741 B.n652 B.n85 10.6151
R1742 B.n652 B.n651 10.6151
R1743 B.n651 B.n650 10.6151
R1744 B.n472 B.n471 10.6151
R1745 B.n472 B.n145 10.6151
R1746 B.n476 B.n145 10.6151
R1747 B.n477 B.n476 10.6151
R1748 B.n478 B.n477 10.6151
R1749 B.n478 B.n143 10.6151
R1750 B.n482 B.n143 10.6151
R1751 B.n483 B.n482 10.6151
R1752 B.n484 B.n483 10.6151
R1753 B.n484 B.n141 10.6151
R1754 B.n488 B.n141 10.6151
R1755 B.n489 B.n488 10.6151
R1756 B.n490 B.n489 10.6151
R1757 B.n490 B.n139 10.6151
R1758 B.n494 B.n139 10.6151
R1759 B.n495 B.n494 10.6151
R1760 B.n496 B.n495 10.6151
R1761 B.n496 B.n137 10.6151
R1762 B.n500 B.n137 10.6151
R1763 B.n501 B.n500 10.6151
R1764 B.n502 B.n501 10.6151
R1765 B.n502 B.n135 10.6151
R1766 B.n506 B.n135 10.6151
R1767 B.n507 B.n506 10.6151
R1768 B.n508 B.n507 10.6151
R1769 B.n508 B.n133 10.6151
R1770 B.n512 B.n133 10.6151
R1771 B.n513 B.n512 10.6151
R1772 B.n514 B.n513 10.6151
R1773 B.n514 B.n131 10.6151
R1774 B.n518 B.n131 10.6151
R1775 B.n519 B.n518 10.6151
R1776 B.n520 B.n519 10.6151
R1777 B.n520 B.n129 10.6151
R1778 B.n524 B.n129 10.6151
R1779 B.n525 B.n524 10.6151
R1780 B.n526 B.n525 10.6151
R1781 B.n526 B.n127 10.6151
R1782 B.n530 B.n127 10.6151
R1783 B.n531 B.n530 10.6151
R1784 B.n532 B.n531 10.6151
R1785 B.n532 B.n125 10.6151
R1786 B.n536 B.n125 10.6151
R1787 B.n537 B.n536 10.6151
R1788 B.n538 B.n537 10.6151
R1789 B.n538 B.n123 10.6151
R1790 B.n542 B.n123 10.6151
R1791 B.n543 B.n542 10.6151
R1792 B.n544 B.n543 10.6151
R1793 B.n544 B.n121 10.6151
R1794 B.n548 B.n121 10.6151
R1795 B.n549 B.n548 10.6151
R1796 B.n550 B.n549 10.6151
R1797 B.n550 B.n119 10.6151
R1798 B.n554 B.n119 10.6151
R1799 B.n555 B.n554 10.6151
R1800 B.n556 B.n555 10.6151
R1801 B.n556 B.n117 10.6151
R1802 B.n560 B.n117 10.6151
R1803 B.n561 B.n560 10.6151
R1804 B.n562 B.n561 10.6151
R1805 B.n562 B.n115 10.6151
R1806 B.n566 B.n115 10.6151
R1807 B.n567 B.n566 10.6151
R1808 B.n568 B.n567 10.6151
R1809 B.n568 B.n113 10.6151
R1810 B.n572 B.n113 10.6151
R1811 B.n573 B.n572 10.6151
R1812 B.n574 B.n573 10.6151
R1813 B.n574 B.n111 10.6151
R1814 B.n578 B.n111 10.6151
R1815 B.n579 B.n578 10.6151
R1816 B.n580 B.n579 10.6151
R1817 B.n580 B.n109 10.6151
R1818 B.n584 B.n109 10.6151
R1819 B.n585 B.n584 10.6151
R1820 B.n586 B.n585 10.6151
R1821 B.n586 B.n107 10.6151
R1822 B.n590 B.n107 10.6151
R1823 B.n591 B.n590 10.6151
R1824 B.n592 B.n591 10.6151
R1825 B.n592 B.n105 10.6151
R1826 B.n596 B.n105 10.6151
R1827 B.n597 B.n596 10.6151
R1828 B.n598 B.n597 10.6151
R1829 B.n598 B.n103 10.6151
R1830 B.n602 B.n103 10.6151
R1831 B.n603 B.n602 10.6151
R1832 B.n604 B.n603 10.6151
R1833 B.n604 B.n101 10.6151
R1834 B.n608 B.n101 10.6151
R1835 B.n609 B.n608 10.6151
R1836 B.n610 B.n609 10.6151
R1837 B.n610 B.n99 10.6151
R1838 B.n614 B.n99 10.6151
R1839 B.n615 B.n614 10.6151
R1840 B.n616 B.n615 10.6151
R1841 B.n616 B.n97 10.6151
R1842 B.n620 B.n97 10.6151
R1843 B.n621 B.n620 10.6151
R1844 B.n622 B.n621 10.6151
R1845 B.n622 B.n95 10.6151
R1846 B.n626 B.n95 10.6151
R1847 B.n627 B.n626 10.6151
R1848 B.n628 B.n627 10.6151
R1849 B.n628 B.n93 10.6151
R1850 B.n632 B.n93 10.6151
R1851 B.n633 B.n632 10.6151
R1852 B.n634 B.n633 10.6151
R1853 B.n634 B.n91 10.6151
R1854 B.n638 B.n91 10.6151
R1855 B.n639 B.n638 10.6151
R1856 B.n640 B.n639 10.6151
R1857 B.n640 B.n89 10.6151
R1858 B.n644 B.n89 10.6151
R1859 B.n645 B.n644 10.6151
R1860 B.n646 B.n645 10.6151
R1861 B.n646 B.n87 10.6151
R1862 B.n317 B.n316 10.6151
R1863 B.n318 B.n317 10.6151
R1864 B.n318 B.n197 10.6151
R1865 B.n322 B.n197 10.6151
R1866 B.n323 B.n322 10.6151
R1867 B.n324 B.n323 10.6151
R1868 B.n324 B.n195 10.6151
R1869 B.n328 B.n195 10.6151
R1870 B.n329 B.n328 10.6151
R1871 B.n330 B.n329 10.6151
R1872 B.n330 B.n193 10.6151
R1873 B.n334 B.n193 10.6151
R1874 B.n335 B.n334 10.6151
R1875 B.n336 B.n335 10.6151
R1876 B.n336 B.n191 10.6151
R1877 B.n340 B.n191 10.6151
R1878 B.n341 B.n340 10.6151
R1879 B.n342 B.n341 10.6151
R1880 B.n342 B.n189 10.6151
R1881 B.n346 B.n189 10.6151
R1882 B.n347 B.n346 10.6151
R1883 B.n348 B.n347 10.6151
R1884 B.n348 B.n187 10.6151
R1885 B.n352 B.n187 10.6151
R1886 B.n353 B.n352 10.6151
R1887 B.n354 B.n353 10.6151
R1888 B.n354 B.n185 10.6151
R1889 B.n358 B.n185 10.6151
R1890 B.n359 B.n358 10.6151
R1891 B.n360 B.n359 10.6151
R1892 B.n360 B.n183 10.6151
R1893 B.n364 B.n183 10.6151
R1894 B.n365 B.n364 10.6151
R1895 B.n366 B.n365 10.6151
R1896 B.n366 B.n181 10.6151
R1897 B.n370 B.n181 10.6151
R1898 B.n371 B.n370 10.6151
R1899 B.n372 B.n371 10.6151
R1900 B.n372 B.n179 10.6151
R1901 B.n376 B.n179 10.6151
R1902 B.n377 B.n376 10.6151
R1903 B.n378 B.n377 10.6151
R1904 B.n378 B.n177 10.6151
R1905 B.n382 B.n177 10.6151
R1906 B.n383 B.n382 10.6151
R1907 B.n385 B.n173 10.6151
R1908 B.n389 B.n173 10.6151
R1909 B.n390 B.n389 10.6151
R1910 B.n391 B.n390 10.6151
R1911 B.n391 B.n171 10.6151
R1912 B.n395 B.n171 10.6151
R1913 B.n396 B.n395 10.6151
R1914 B.n400 B.n396 10.6151
R1915 B.n404 B.n169 10.6151
R1916 B.n405 B.n404 10.6151
R1917 B.n406 B.n405 10.6151
R1918 B.n406 B.n167 10.6151
R1919 B.n410 B.n167 10.6151
R1920 B.n411 B.n410 10.6151
R1921 B.n412 B.n411 10.6151
R1922 B.n412 B.n165 10.6151
R1923 B.n416 B.n165 10.6151
R1924 B.n417 B.n416 10.6151
R1925 B.n418 B.n417 10.6151
R1926 B.n418 B.n163 10.6151
R1927 B.n422 B.n163 10.6151
R1928 B.n423 B.n422 10.6151
R1929 B.n424 B.n423 10.6151
R1930 B.n424 B.n161 10.6151
R1931 B.n428 B.n161 10.6151
R1932 B.n429 B.n428 10.6151
R1933 B.n430 B.n429 10.6151
R1934 B.n430 B.n159 10.6151
R1935 B.n434 B.n159 10.6151
R1936 B.n435 B.n434 10.6151
R1937 B.n436 B.n435 10.6151
R1938 B.n436 B.n157 10.6151
R1939 B.n440 B.n157 10.6151
R1940 B.n441 B.n440 10.6151
R1941 B.n442 B.n441 10.6151
R1942 B.n442 B.n155 10.6151
R1943 B.n446 B.n155 10.6151
R1944 B.n447 B.n446 10.6151
R1945 B.n448 B.n447 10.6151
R1946 B.n448 B.n153 10.6151
R1947 B.n452 B.n153 10.6151
R1948 B.n453 B.n452 10.6151
R1949 B.n454 B.n453 10.6151
R1950 B.n454 B.n151 10.6151
R1951 B.n458 B.n151 10.6151
R1952 B.n459 B.n458 10.6151
R1953 B.n460 B.n459 10.6151
R1954 B.n460 B.n149 10.6151
R1955 B.n464 B.n149 10.6151
R1956 B.n465 B.n464 10.6151
R1957 B.n466 B.n465 10.6151
R1958 B.n466 B.n147 10.6151
R1959 B.n470 B.n147 10.6151
R1960 B.n312 B.n199 10.6151
R1961 B.n312 B.n311 10.6151
R1962 B.n311 B.n310 10.6151
R1963 B.n310 B.n201 10.6151
R1964 B.n306 B.n201 10.6151
R1965 B.n306 B.n305 10.6151
R1966 B.n305 B.n304 10.6151
R1967 B.n304 B.n203 10.6151
R1968 B.n300 B.n203 10.6151
R1969 B.n300 B.n299 10.6151
R1970 B.n299 B.n298 10.6151
R1971 B.n298 B.n205 10.6151
R1972 B.n294 B.n205 10.6151
R1973 B.n294 B.n293 10.6151
R1974 B.n293 B.n292 10.6151
R1975 B.n292 B.n207 10.6151
R1976 B.n288 B.n207 10.6151
R1977 B.n288 B.n287 10.6151
R1978 B.n287 B.n286 10.6151
R1979 B.n286 B.n209 10.6151
R1980 B.n282 B.n209 10.6151
R1981 B.n282 B.n281 10.6151
R1982 B.n281 B.n280 10.6151
R1983 B.n280 B.n211 10.6151
R1984 B.n276 B.n211 10.6151
R1985 B.n276 B.n275 10.6151
R1986 B.n275 B.n274 10.6151
R1987 B.n274 B.n213 10.6151
R1988 B.n270 B.n213 10.6151
R1989 B.n270 B.n269 10.6151
R1990 B.n269 B.n268 10.6151
R1991 B.n268 B.n215 10.6151
R1992 B.n264 B.n215 10.6151
R1993 B.n264 B.n263 10.6151
R1994 B.n263 B.n262 10.6151
R1995 B.n262 B.n217 10.6151
R1996 B.n258 B.n217 10.6151
R1997 B.n258 B.n257 10.6151
R1998 B.n257 B.n256 10.6151
R1999 B.n256 B.n219 10.6151
R2000 B.n252 B.n219 10.6151
R2001 B.n252 B.n251 10.6151
R2002 B.n251 B.n250 10.6151
R2003 B.n250 B.n221 10.6151
R2004 B.n246 B.n221 10.6151
R2005 B.n246 B.n245 10.6151
R2006 B.n245 B.n244 10.6151
R2007 B.n244 B.n223 10.6151
R2008 B.n240 B.n223 10.6151
R2009 B.n240 B.n239 10.6151
R2010 B.n239 B.n238 10.6151
R2011 B.n238 B.n225 10.6151
R2012 B.n234 B.n225 10.6151
R2013 B.n234 B.n233 10.6151
R2014 B.n233 B.n232 10.6151
R2015 B.n232 B.n227 10.6151
R2016 B.n228 B.n227 10.6151
R2017 B.n228 B.n0 10.6151
R2018 B.n887 B.n1 10.6151
R2019 B.n887 B.n886 10.6151
R2020 B.n886 B.n885 10.6151
R2021 B.n885 B.n4 10.6151
R2022 B.n881 B.n4 10.6151
R2023 B.n881 B.n880 10.6151
R2024 B.n880 B.n879 10.6151
R2025 B.n879 B.n6 10.6151
R2026 B.n875 B.n6 10.6151
R2027 B.n875 B.n874 10.6151
R2028 B.n874 B.n873 10.6151
R2029 B.n873 B.n8 10.6151
R2030 B.n869 B.n8 10.6151
R2031 B.n869 B.n868 10.6151
R2032 B.n868 B.n867 10.6151
R2033 B.n867 B.n10 10.6151
R2034 B.n863 B.n10 10.6151
R2035 B.n863 B.n862 10.6151
R2036 B.n862 B.n861 10.6151
R2037 B.n861 B.n12 10.6151
R2038 B.n857 B.n12 10.6151
R2039 B.n857 B.n856 10.6151
R2040 B.n856 B.n855 10.6151
R2041 B.n855 B.n14 10.6151
R2042 B.n851 B.n14 10.6151
R2043 B.n851 B.n850 10.6151
R2044 B.n850 B.n849 10.6151
R2045 B.n849 B.n16 10.6151
R2046 B.n845 B.n16 10.6151
R2047 B.n845 B.n844 10.6151
R2048 B.n844 B.n843 10.6151
R2049 B.n843 B.n18 10.6151
R2050 B.n839 B.n18 10.6151
R2051 B.n839 B.n838 10.6151
R2052 B.n838 B.n837 10.6151
R2053 B.n837 B.n20 10.6151
R2054 B.n833 B.n20 10.6151
R2055 B.n833 B.n832 10.6151
R2056 B.n832 B.n831 10.6151
R2057 B.n831 B.n22 10.6151
R2058 B.n827 B.n22 10.6151
R2059 B.n827 B.n826 10.6151
R2060 B.n826 B.n825 10.6151
R2061 B.n825 B.n24 10.6151
R2062 B.n821 B.n24 10.6151
R2063 B.n821 B.n820 10.6151
R2064 B.n820 B.n819 10.6151
R2065 B.n819 B.n26 10.6151
R2066 B.n815 B.n26 10.6151
R2067 B.n815 B.n814 10.6151
R2068 B.n814 B.n813 10.6151
R2069 B.n813 B.n28 10.6151
R2070 B.n809 B.n28 10.6151
R2071 B.n809 B.n808 10.6151
R2072 B.n808 B.n807 10.6151
R2073 B.n807 B.n30 10.6151
R2074 B.n803 B.n30 10.6151
R2075 B.n803 B.n802 10.6151
R2076 B.n731 B.n58 6.5566
R2077 B.n719 B.n718 6.5566
R2078 B.n385 B.n384 6.5566
R2079 B.n400 B.n399 6.5566
R2080 B.n58 B.n54 4.05904
R2081 B.n718 B.n717 4.05904
R2082 B.n384 B.n383 4.05904
R2083 B.n399 B.n169 4.05904
R2084 B.n891 B.n0 2.81026
R2085 B.n891 B.n1 2.81026
R2086 VP.n16 VP.n15 161.3
R2087 VP.n17 VP.n12 161.3
R2088 VP.n19 VP.n18 161.3
R2089 VP.n20 VP.n11 161.3
R2090 VP.n22 VP.n21 161.3
R2091 VP.n23 VP.n10 161.3
R2092 VP.n25 VP.n24 161.3
R2093 VP.n26 VP.n9 161.3
R2094 VP.n55 VP.n0 161.3
R2095 VP.n54 VP.n53 161.3
R2096 VP.n52 VP.n1 161.3
R2097 VP.n51 VP.n50 161.3
R2098 VP.n49 VP.n2 161.3
R2099 VP.n48 VP.n47 161.3
R2100 VP.n46 VP.n3 161.3
R2101 VP.n45 VP.n44 161.3
R2102 VP.n43 VP.n4 161.3
R2103 VP.n42 VP.n41 161.3
R2104 VP.n40 VP.n5 161.3
R2105 VP.n39 VP.n38 161.3
R2106 VP.n37 VP.n6 161.3
R2107 VP.n36 VP.n35 161.3
R2108 VP.n34 VP.n7 161.3
R2109 VP.n33 VP.n32 161.3
R2110 VP.n31 VP.n8 161.3
R2111 VP.n13 VP.t5 113.513
R2112 VP.n43 VP.t4 80.3137
R2113 VP.n30 VP.t2 80.3137
R2114 VP.n56 VP.t3 80.3137
R2115 VP.n27 VP.t0 80.3137
R2116 VP.n14 VP.t1 80.3137
R2117 VP.n30 VP.n29 66.0336
R2118 VP.n57 VP.n56 66.0336
R2119 VP.n28 VP.n27 66.0336
R2120 VP.n37 VP.n36 56.5193
R2121 VP.n50 VP.n49 56.5193
R2122 VP.n21 VP.n20 56.5193
R2123 VP.n29 VP.n28 55.3563
R2124 VP.n14 VP.n13 50.5569
R2125 VP.n32 VP.n31 24.4675
R2126 VP.n32 VP.n7 24.4675
R2127 VP.n36 VP.n7 24.4675
R2128 VP.n38 VP.n37 24.4675
R2129 VP.n38 VP.n5 24.4675
R2130 VP.n42 VP.n5 24.4675
R2131 VP.n43 VP.n42 24.4675
R2132 VP.n44 VP.n43 24.4675
R2133 VP.n44 VP.n3 24.4675
R2134 VP.n48 VP.n3 24.4675
R2135 VP.n49 VP.n48 24.4675
R2136 VP.n50 VP.n1 24.4675
R2137 VP.n54 VP.n1 24.4675
R2138 VP.n55 VP.n54 24.4675
R2139 VP.n21 VP.n10 24.4675
R2140 VP.n25 VP.n10 24.4675
R2141 VP.n26 VP.n25 24.4675
R2142 VP.n15 VP.n14 24.4675
R2143 VP.n15 VP.n12 24.4675
R2144 VP.n19 VP.n12 24.4675
R2145 VP.n20 VP.n19 24.4675
R2146 VP.n31 VP.n30 16.1487
R2147 VP.n56 VP.n55 16.1487
R2148 VP.n27 VP.n26 16.1487
R2149 VP.n16 VP.n13 2.09745
R2150 VP.n28 VP.n9 0.417535
R2151 VP.n29 VP.n8 0.417535
R2152 VP.n57 VP.n0 0.417535
R2153 VP VP.n57 0.394291
R2154 VP.n17 VP.n16 0.189894
R2155 VP.n18 VP.n17 0.189894
R2156 VP.n18 VP.n11 0.189894
R2157 VP.n22 VP.n11 0.189894
R2158 VP.n23 VP.n22 0.189894
R2159 VP.n24 VP.n23 0.189894
R2160 VP.n24 VP.n9 0.189894
R2161 VP.n33 VP.n8 0.189894
R2162 VP.n34 VP.n33 0.189894
R2163 VP.n35 VP.n34 0.189894
R2164 VP.n35 VP.n6 0.189894
R2165 VP.n39 VP.n6 0.189894
R2166 VP.n40 VP.n39 0.189894
R2167 VP.n41 VP.n40 0.189894
R2168 VP.n41 VP.n4 0.189894
R2169 VP.n45 VP.n4 0.189894
R2170 VP.n46 VP.n45 0.189894
R2171 VP.n47 VP.n46 0.189894
R2172 VP.n47 VP.n2 0.189894
R2173 VP.n51 VP.n2 0.189894
R2174 VP.n52 VP.n51 0.189894
R2175 VP.n53 VP.n52 0.189894
R2176 VP.n53 VP.n0 0.189894
R2177 VDD1.n67 VDD1.n66 585
R2178 VDD1.n65 VDD1.n64 585
R2179 VDD1.n4 VDD1.n3 585
R2180 VDD1.n59 VDD1.n58 585
R2181 VDD1.n57 VDD1.n56 585
R2182 VDD1.n8 VDD1.n7 585
R2183 VDD1.n51 VDD1.n50 585
R2184 VDD1.n49 VDD1.n48 585
R2185 VDD1.n12 VDD1.n11 585
R2186 VDD1.n43 VDD1.n42 585
R2187 VDD1.n41 VDD1.n40 585
R2188 VDD1.n16 VDD1.n15 585
R2189 VDD1.n35 VDD1.n34 585
R2190 VDD1.n33 VDD1.n32 585
R2191 VDD1.n20 VDD1.n19 585
R2192 VDD1.n27 VDD1.n26 585
R2193 VDD1.n25 VDD1.n24 585
R2194 VDD1.n96 VDD1.n95 585
R2195 VDD1.n98 VDD1.n97 585
R2196 VDD1.n91 VDD1.n90 585
R2197 VDD1.n104 VDD1.n103 585
R2198 VDD1.n106 VDD1.n105 585
R2199 VDD1.n87 VDD1.n86 585
R2200 VDD1.n112 VDD1.n111 585
R2201 VDD1.n114 VDD1.n113 585
R2202 VDD1.n83 VDD1.n82 585
R2203 VDD1.n120 VDD1.n119 585
R2204 VDD1.n122 VDD1.n121 585
R2205 VDD1.n79 VDD1.n78 585
R2206 VDD1.n128 VDD1.n127 585
R2207 VDD1.n130 VDD1.n129 585
R2208 VDD1.n75 VDD1.n74 585
R2209 VDD1.n136 VDD1.n135 585
R2210 VDD1.n138 VDD1.n137 585
R2211 VDD1.n66 VDD1.n0 498.474
R2212 VDD1.n137 VDD1.n71 498.474
R2213 VDD1.n23 VDD1.t0 327.466
R2214 VDD1.n94 VDD1.t3 327.466
R2215 VDD1.n66 VDD1.n65 171.744
R2216 VDD1.n65 VDD1.n3 171.744
R2217 VDD1.n58 VDD1.n3 171.744
R2218 VDD1.n58 VDD1.n57 171.744
R2219 VDD1.n57 VDD1.n7 171.744
R2220 VDD1.n50 VDD1.n7 171.744
R2221 VDD1.n50 VDD1.n49 171.744
R2222 VDD1.n49 VDD1.n11 171.744
R2223 VDD1.n42 VDD1.n11 171.744
R2224 VDD1.n42 VDD1.n41 171.744
R2225 VDD1.n41 VDD1.n15 171.744
R2226 VDD1.n34 VDD1.n15 171.744
R2227 VDD1.n34 VDD1.n33 171.744
R2228 VDD1.n33 VDD1.n19 171.744
R2229 VDD1.n26 VDD1.n19 171.744
R2230 VDD1.n26 VDD1.n25 171.744
R2231 VDD1.n97 VDD1.n96 171.744
R2232 VDD1.n97 VDD1.n90 171.744
R2233 VDD1.n104 VDD1.n90 171.744
R2234 VDD1.n105 VDD1.n104 171.744
R2235 VDD1.n105 VDD1.n86 171.744
R2236 VDD1.n112 VDD1.n86 171.744
R2237 VDD1.n113 VDD1.n112 171.744
R2238 VDD1.n113 VDD1.n82 171.744
R2239 VDD1.n120 VDD1.n82 171.744
R2240 VDD1.n121 VDD1.n120 171.744
R2241 VDD1.n121 VDD1.n78 171.744
R2242 VDD1.n128 VDD1.n78 171.744
R2243 VDD1.n129 VDD1.n128 171.744
R2244 VDD1.n129 VDD1.n74 171.744
R2245 VDD1.n136 VDD1.n74 171.744
R2246 VDD1.n137 VDD1.n136 171.744
R2247 VDD1.n25 VDD1.t0 85.8723
R2248 VDD1.n96 VDD1.t3 85.8723
R2249 VDD1.n143 VDD1.n142 75.3655
R2250 VDD1.n145 VDD1.n144 74.4876
R2251 VDD1 VDD1.n70 54.2431
R2252 VDD1.n143 VDD1.n141 54.1296
R2253 VDD1.n145 VDD1.n143 49.7875
R2254 VDD1.n24 VDD1.n23 16.3895
R2255 VDD1.n95 VDD1.n94 16.3895
R2256 VDD1.n68 VDD1.n67 12.8005
R2257 VDD1.n27 VDD1.n22 12.8005
R2258 VDD1.n98 VDD1.n93 12.8005
R2259 VDD1.n139 VDD1.n138 12.8005
R2260 VDD1.n64 VDD1.n2 12.0247
R2261 VDD1.n28 VDD1.n20 12.0247
R2262 VDD1.n99 VDD1.n91 12.0247
R2263 VDD1.n135 VDD1.n73 12.0247
R2264 VDD1.n63 VDD1.n4 11.249
R2265 VDD1.n32 VDD1.n31 11.249
R2266 VDD1.n103 VDD1.n102 11.249
R2267 VDD1.n134 VDD1.n75 11.249
R2268 VDD1.n60 VDD1.n59 10.4732
R2269 VDD1.n35 VDD1.n18 10.4732
R2270 VDD1.n106 VDD1.n89 10.4732
R2271 VDD1.n131 VDD1.n130 10.4732
R2272 VDD1.n56 VDD1.n6 9.69747
R2273 VDD1.n36 VDD1.n16 9.69747
R2274 VDD1.n107 VDD1.n87 9.69747
R2275 VDD1.n127 VDD1.n77 9.69747
R2276 VDD1.n70 VDD1.n69 9.45567
R2277 VDD1.n141 VDD1.n140 9.45567
R2278 VDD1.n10 VDD1.n9 9.3005
R2279 VDD1.n53 VDD1.n52 9.3005
R2280 VDD1.n55 VDD1.n54 9.3005
R2281 VDD1.n6 VDD1.n5 9.3005
R2282 VDD1.n61 VDD1.n60 9.3005
R2283 VDD1.n63 VDD1.n62 9.3005
R2284 VDD1.n2 VDD1.n1 9.3005
R2285 VDD1.n69 VDD1.n68 9.3005
R2286 VDD1.n47 VDD1.n46 9.3005
R2287 VDD1.n45 VDD1.n44 9.3005
R2288 VDD1.n14 VDD1.n13 9.3005
R2289 VDD1.n39 VDD1.n38 9.3005
R2290 VDD1.n37 VDD1.n36 9.3005
R2291 VDD1.n18 VDD1.n17 9.3005
R2292 VDD1.n31 VDD1.n30 9.3005
R2293 VDD1.n29 VDD1.n28 9.3005
R2294 VDD1.n22 VDD1.n21 9.3005
R2295 VDD1.n116 VDD1.n115 9.3005
R2296 VDD1.n85 VDD1.n84 9.3005
R2297 VDD1.n110 VDD1.n109 9.3005
R2298 VDD1.n108 VDD1.n107 9.3005
R2299 VDD1.n89 VDD1.n88 9.3005
R2300 VDD1.n102 VDD1.n101 9.3005
R2301 VDD1.n100 VDD1.n99 9.3005
R2302 VDD1.n93 VDD1.n92 9.3005
R2303 VDD1.n118 VDD1.n117 9.3005
R2304 VDD1.n81 VDD1.n80 9.3005
R2305 VDD1.n124 VDD1.n123 9.3005
R2306 VDD1.n126 VDD1.n125 9.3005
R2307 VDD1.n77 VDD1.n76 9.3005
R2308 VDD1.n132 VDD1.n131 9.3005
R2309 VDD1.n134 VDD1.n133 9.3005
R2310 VDD1.n73 VDD1.n72 9.3005
R2311 VDD1.n140 VDD1.n139 9.3005
R2312 VDD1.n55 VDD1.n8 8.92171
R2313 VDD1.n40 VDD1.n39 8.92171
R2314 VDD1.n111 VDD1.n110 8.92171
R2315 VDD1.n126 VDD1.n79 8.92171
R2316 VDD1.n52 VDD1.n51 8.14595
R2317 VDD1.n43 VDD1.n14 8.14595
R2318 VDD1.n114 VDD1.n85 8.14595
R2319 VDD1.n123 VDD1.n122 8.14595
R2320 VDD1.n70 VDD1.n0 7.75445
R2321 VDD1.n141 VDD1.n71 7.75445
R2322 VDD1.n48 VDD1.n10 7.3702
R2323 VDD1.n44 VDD1.n12 7.3702
R2324 VDD1.n115 VDD1.n83 7.3702
R2325 VDD1.n119 VDD1.n81 7.3702
R2326 VDD1.n48 VDD1.n47 6.59444
R2327 VDD1.n47 VDD1.n12 6.59444
R2328 VDD1.n118 VDD1.n83 6.59444
R2329 VDD1.n119 VDD1.n118 6.59444
R2330 VDD1.n68 VDD1.n0 6.08283
R2331 VDD1.n139 VDD1.n71 6.08283
R2332 VDD1.n51 VDD1.n10 5.81868
R2333 VDD1.n44 VDD1.n43 5.81868
R2334 VDD1.n115 VDD1.n114 5.81868
R2335 VDD1.n122 VDD1.n81 5.81868
R2336 VDD1.n52 VDD1.n8 5.04292
R2337 VDD1.n40 VDD1.n14 5.04292
R2338 VDD1.n111 VDD1.n85 5.04292
R2339 VDD1.n123 VDD1.n79 5.04292
R2340 VDD1.n56 VDD1.n55 4.26717
R2341 VDD1.n39 VDD1.n16 4.26717
R2342 VDD1.n110 VDD1.n87 4.26717
R2343 VDD1.n127 VDD1.n126 4.26717
R2344 VDD1.n23 VDD1.n21 3.70982
R2345 VDD1.n94 VDD1.n92 3.70982
R2346 VDD1.n59 VDD1.n6 3.49141
R2347 VDD1.n36 VDD1.n35 3.49141
R2348 VDD1.n107 VDD1.n106 3.49141
R2349 VDD1.n130 VDD1.n77 3.49141
R2350 VDD1.n60 VDD1.n4 2.71565
R2351 VDD1.n32 VDD1.n18 2.71565
R2352 VDD1.n103 VDD1.n89 2.71565
R2353 VDD1.n131 VDD1.n75 2.71565
R2354 VDD1.n144 VDD1.t4 2.43898
R2355 VDD1.n144 VDD1.t5 2.43898
R2356 VDD1.n142 VDD1.t1 2.43898
R2357 VDD1.n142 VDD1.t2 2.43898
R2358 VDD1.n64 VDD1.n63 1.93989
R2359 VDD1.n31 VDD1.n20 1.93989
R2360 VDD1.n102 VDD1.n91 1.93989
R2361 VDD1.n135 VDD1.n134 1.93989
R2362 VDD1.n67 VDD1.n2 1.16414
R2363 VDD1.n28 VDD1.n27 1.16414
R2364 VDD1.n99 VDD1.n98 1.16414
R2365 VDD1.n138 VDD1.n73 1.16414
R2366 VDD1 VDD1.n145 0.8755
R2367 VDD1.n24 VDD1.n22 0.388379
R2368 VDD1.n95 VDD1.n93 0.388379
R2369 VDD1.n69 VDD1.n1 0.155672
R2370 VDD1.n62 VDD1.n1 0.155672
R2371 VDD1.n62 VDD1.n61 0.155672
R2372 VDD1.n61 VDD1.n5 0.155672
R2373 VDD1.n54 VDD1.n5 0.155672
R2374 VDD1.n54 VDD1.n53 0.155672
R2375 VDD1.n53 VDD1.n9 0.155672
R2376 VDD1.n46 VDD1.n9 0.155672
R2377 VDD1.n46 VDD1.n45 0.155672
R2378 VDD1.n45 VDD1.n13 0.155672
R2379 VDD1.n38 VDD1.n13 0.155672
R2380 VDD1.n38 VDD1.n37 0.155672
R2381 VDD1.n37 VDD1.n17 0.155672
R2382 VDD1.n30 VDD1.n17 0.155672
R2383 VDD1.n30 VDD1.n29 0.155672
R2384 VDD1.n29 VDD1.n21 0.155672
R2385 VDD1.n100 VDD1.n92 0.155672
R2386 VDD1.n101 VDD1.n100 0.155672
R2387 VDD1.n101 VDD1.n88 0.155672
R2388 VDD1.n108 VDD1.n88 0.155672
R2389 VDD1.n109 VDD1.n108 0.155672
R2390 VDD1.n109 VDD1.n84 0.155672
R2391 VDD1.n116 VDD1.n84 0.155672
R2392 VDD1.n117 VDD1.n116 0.155672
R2393 VDD1.n117 VDD1.n80 0.155672
R2394 VDD1.n124 VDD1.n80 0.155672
R2395 VDD1.n125 VDD1.n124 0.155672
R2396 VDD1.n125 VDD1.n76 0.155672
R2397 VDD1.n132 VDD1.n76 0.155672
R2398 VDD1.n133 VDD1.n132 0.155672
R2399 VDD1.n133 VDD1.n72 0.155672
R2400 VDD1.n140 VDD1.n72 0.155672
C0 VP VN 8.5389f
C1 VTAIL VDD2 8.742129f
C2 VN VDD1 0.152746f
C3 B VP 2.44891f
C4 VN VDD2 7.94563f
C5 w_n4434_n3634# VTAIL 3.27735f
C6 B VDD1 2.56335f
C7 VP VDD1 8.36691f
C8 B VDD2 2.67102f
C9 w_n4434_n3634# VN 8.77271f
C10 VP VDD2 0.576502f
C11 VDD1 VDD2 1.95416f
C12 w_n4434_n3634# B 11.9825f
C13 w_n4434_n3634# VP 9.34986f
C14 w_n4434_n3634# VDD1 2.71903f
C15 w_n4434_n3634# VDD2 2.84887f
C16 VN VTAIL 8.378441f
C17 B VTAIL 4.52341f
C18 VP VTAIL 8.39339f
C19 B VN 1.47824f
C20 VTAIL VDD1 8.68103f
C21 VDD2 VSUBS 2.30035f
C22 VDD1 VSUBS 2.36324f
C23 VTAIL VSUBS 1.506865f
C24 VN VSUBS 7.28388f
C25 VP VSUBS 4.084047f
C26 B VSUBS 6.131589f
C27 w_n4434_n3634# VSUBS 0.197987p
C28 VDD1.n0 VSUBS 0.030313f
C29 VDD1.n1 VSUBS 0.028438f
C30 VDD1.n2 VSUBS 0.015282f
C31 VDD1.n3 VSUBS 0.03612f
C32 VDD1.n4 VSUBS 0.016181f
C33 VDD1.n5 VSUBS 0.028438f
C34 VDD1.n6 VSUBS 0.015282f
C35 VDD1.n7 VSUBS 0.03612f
C36 VDD1.n8 VSUBS 0.016181f
C37 VDD1.n9 VSUBS 0.028438f
C38 VDD1.n10 VSUBS 0.015282f
C39 VDD1.n11 VSUBS 0.03612f
C40 VDD1.n12 VSUBS 0.016181f
C41 VDD1.n13 VSUBS 0.028438f
C42 VDD1.n14 VSUBS 0.015282f
C43 VDD1.n15 VSUBS 0.03612f
C44 VDD1.n16 VSUBS 0.016181f
C45 VDD1.n17 VSUBS 0.028438f
C46 VDD1.n18 VSUBS 0.015282f
C47 VDD1.n19 VSUBS 0.03612f
C48 VDD1.n20 VSUBS 0.016181f
C49 VDD1.n21 VSUBS 1.60025f
C50 VDD1.n22 VSUBS 0.015282f
C51 VDD1.t0 VSUBS 0.077209f
C52 VDD1.n23 VSUBS 0.186459f
C53 VDD1.n24 VSUBS 0.022978f
C54 VDD1.n25 VSUBS 0.02709f
C55 VDD1.n26 VSUBS 0.03612f
C56 VDD1.n27 VSUBS 0.016181f
C57 VDD1.n28 VSUBS 0.015282f
C58 VDD1.n29 VSUBS 0.028438f
C59 VDD1.n30 VSUBS 0.028438f
C60 VDD1.n31 VSUBS 0.015282f
C61 VDD1.n32 VSUBS 0.016181f
C62 VDD1.n33 VSUBS 0.03612f
C63 VDD1.n34 VSUBS 0.03612f
C64 VDD1.n35 VSUBS 0.016181f
C65 VDD1.n36 VSUBS 0.015282f
C66 VDD1.n37 VSUBS 0.028438f
C67 VDD1.n38 VSUBS 0.028438f
C68 VDD1.n39 VSUBS 0.015282f
C69 VDD1.n40 VSUBS 0.016181f
C70 VDD1.n41 VSUBS 0.03612f
C71 VDD1.n42 VSUBS 0.03612f
C72 VDD1.n43 VSUBS 0.016181f
C73 VDD1.n44 VSUBS 0.015282f
C74 VDD1.n45 VSUBS 0.028438f
C75 VDD1.n46 VSUBS 0.028438f
C76 VDD1.n47 VSUBS 0.015282f
C77 VDD1.n48 VSUBS 0.016181f
C78 VDD1.n49 VSUBS 0.03612f
C79 VDD1.n50 VSUBS 0.03612f
C80 VDD1.n51 VSUBS 0.016181f
C81 VDD1.n52 VSUBS 0.015282f
C82 VDD1.n53 VSUBS 0.028438f
C83 VDD1.n54 VSUBS 0.028438f
C84 VDD1.n55 VSUBS 0.015282f
C85 VDD1.n56 VSUBS 0.016181f
C86 VDD1.n57 VSUBS 0.03612f
C87 VDD1.n58 VSUBS 0.03612f
C88 VDD1.n59 VSUBS 0.016181f
C89 VDD1.n60 VSUBS 0.015282f
C90 VDD1.n61 VSUBS 0.028438f
C91 VDD1.n62 VSUBS 0.028438f
C92 VDD1.n63 VSUBS 0.015282f
C93 VDD1.n64 VSUBS 0.016181f
C94 VDD1.n65 VSUBS 0.03612f
C95 VDD1.n66 VSUBS 0.089133f
C96 VDD1.n67 VSUBS 0.016181f
C97 VDD1.n68 VSUBS 0.030009f
C98 VDD1.n69 VSUBS 0.070784f
C99 VDD1.n70 VSUBS 0.104392f
C100 VDD1.n71 VSUBS 0.030313f
C101 VDD1.n72 VSUBS 0.028438f
C102 VDD1.n73 VSUBS 0.015282f
C103 VDD1.n74 VSUBS 0.03612f
C104 VDD1.n75 VSUBS 0.016181f
C105 VDD1.n76 VSUBS 0.028438f
C106 VDD1.n77 VSUBS 0.015282f
C107 VDD1.n78 VSUBS 0.03612f
C108 VDD1.n79 VSUBS 0.016181f
C109 VDD1.n80 VSUBS 0.028438f
C110 VDD1.n81 VSUBS 0.015282f
C111 VDD1.n82 VSUBS 0.03612f
C112 VDD1.n83 VSUBS 0.016181f
C113 VDD1.n84 VSUBS 0.028438f
C114 VDD1.n85 VSUBS 0.015282f
C115 VDD1.n86 VSUBS 0.03612f
C116 VDD1.n87 VSUBS 0.016181f
C117 VDD1.n88 VSUBS 0.028438f
C118 VDD1.n89 VSUBS 0.015282f
C119 VDD1.n90 VSUBS 0.03612f
C120 VDD1.n91 VSUBS 0.016181f
C121 VDD1.n92 VSUBS 1.60025f
C122 VDD1.n93 VSUBS 0.015282f
C123 VDD1.t3 VSUBS 0.077209f
C124 VDD1.n94 VSUBS 0.186459f
C125 VDD1.n95 VSUBS 0.022978f
C126 VDD1.n96 VSUBS 0.02709f
C127 VDD1.n97 VSUBS 0.03612f
C128 VDD1.n98 VSUBS 0.016181f
C129 VDD1.n99 VSUBS 0.015282f
C130 VDD1.n100 VSUBS 0.028438f
C131 VDD1.n101 VSUBS 0.028438f
C132 VDD1.n102 VSUBS 0.015282f
C133 VDD1.n103 VSUBS 0.016181f
C134 VDD1.n104 VSUBS 0.03612f
C135 VDD1.n105 VSUBS 0.03612f
C136 VDD1.n106 VSUBS 0.016181f
C137 VDD1.n107 VSUBS 0.015282f
C138 VDD1.n108 VSUBS 0.028438f
C139 VDD1.n109 VSUBS 0.028438f
C140 VDD1.n110 VSUBS 0.015282f
C141 VDD1.n111 VSUBS 0.016181f
C142 VDD1.n112 VSUBS 0.03612f
C143 VDD1.n113 VSUBS 0.03612f
C144 VDD1.n114 VSUBS 0.016181f
C145 VDD1.n115 VSUBS 0.015282f
C146 VDD1.n116 VSUBS 0.028438f
C147 VDD1.n117 VSUBS 0.028438f
C148 VDD1.n118 VSUBS 0.015282f
C149 VDD1.n119 VSUBS 0.016181f
C150 VDD1.n120 VSUBS 0.03612f
C151 VDD1.n121 VSUBS 0.03612f
C152 VDD1.n122 VSUBS 0.016181f
C153 VDD1.n123 VSUBS 0.015282f
C154 VDD1.n124 VSUBS 0.028438f
C155 VDD1.n125 VSUBS 0.028438f
C156 VDD1.n126 VSUBS 0.015282f
C157 VDD1.n127 VSUBS 0.016181f
C158 VDD1.n128 VSUBS 0.03612f
C159 VDD1.n129 VSUBS 0.03612f
C160 VDD1.n130 VSUBS 0.016181f
C161 VDD1.n131 VSUBS 0.015282f
C162 VDD1.n132 VSUBS 0.028438f
C163 VDD1.n133 VSUBS 0.028438f
C164 VDD1.n134 VSUBS 0.015282f
C165 VDD1.n135 VSUBS 0.016181f
C166 VDD1.n136 VSUBS 0.03612f
C167 VDD1.n137 VSUBS 0.089133f
C168 VDD1.n138 VSUBS 0.016181f
C169 VDD1.n139 VSUBS 0.030009f
C170 VDD1.n140 VSUBS 0.070784f
C171 VDD1.n141 VSUBS 0.103242f
C172 VDD1.t1 VSUBS 0.299564f
C173 VDD1.t2 VSUBS 0.299564f
C174 VDD1.n142 VSUBS 2.41065f
C175 VDD1.n143 VSUBS 4.30238f
C176 VDD1.t4 VSUBS 0.299564f
C177 VDD1.t5 VSUBS 0.299564f
C178 VDD1.n144 VSUBS 2.39949f
C179 VDD1.n145 VSUBS 4.02488f
C180 VP.n0 VSUBS 0.048432f
C181 VP.t3 VSUBS 3.75129f
C182 VP.n1 VSUBS 0.047988f
C183 VP.n2 VSUBS 0.025748f
C184 VP.n3 VSUBS 0.047988f
C185 VP.n4 VSUBS 0.025748f
C186 VP.t4 VSUBS 3.75129f
C187 VP.n5 VSUBS 0.047988f
C188 VP.n6 VSUBS 0.025748f
C189 VP.n7 VSUBS 0.047988f
C190 VP.n8 VSUBS 0.048432f
C191 VP.t2 VSUBS 3.75129f
C192 VP.n9 VSUBS 0.048432f
C193 VP.t0 VSUBS 3.75129f
C194 VP.n10 VSUBS 0.047988f
C195 VP.n11 VSUBS 0.025748f
C196 VP.n12 VSUBS 0.047988f
C197 VP.t5 VSUBS 4.19369f
C198 VP.n13 VSUBS 1.33983f
C199 VP.t1 VSUBS 3.75129f
C200 VP.n14 VSUBS 1.41395f
C201 VP.n15 VSUBS 0.047988f
C202 VP.n16 VSUBS 0.342474f
C203 VP.n17 VSUBS 0.025748f
C204 VP.n18 VSUBS 0.025748f
C205 VP.n19 VSUBS 0.047988f
C206 VP.n20 VSUBS 0.031492f
C207 VP.n21 VSUBS 0.043689f
C208 VP.n22 VSUBS 0.025748f
C209 VP.n23 VSUBS 0.025748f
C210 VP.n24 VSUBS 0.025748f
C211 VP.n25 VSUBS 0.047988f
C212 VP.n26 VSUBS 0.039933f
C213 VP.n27 VSUBS 1.41275f
C214 VP.n28 VSUBS 1.72841f
C215 VP.n29 VSUBS 1.74513f
C216 VP.n30 VSUBS 1.41275f
C217 VP.n31 VSUBS 0.039933f
C218 VP.n32 VSUBS 0.047988f
C219 VP.n33 VSUBS 0.025748f
C220 VP.n34 VSUBS 0.025748f
C221 VP.n35 VSUBS 0.025748f
C222 VP.n36 VSUBS 0.043689f
C223 VP.n37 VSUBS 0.031492f
C224 VP.n38 VSUBS 0.047988f
C225 VP.n39 VSUBS 0.025748f
C226 VP.n40 VSUBS 0.025748f
C227 VP.n41 VSUBS 0.025748f
C228 VP.n42 VSUBS 0.047988f
C229 VP.n43 VSUBS 1.33049f
C230 VP.n44 VSUBS 0.047988f
C231 VP.n45 VSUBS 0.025748f
C232 VP.n46 VSUBS 0.025748f
C233 VP.n47 VSUBS 0.025748f
C234 VP.n48 VSUBS 0.047988f
C235 VP.n49 VSUBS 0.031492f
C236 VP.n50 VSUBS 0.043689f
C237 VP.n51 VSUBS 0.025748f
C238 VP.n52 VSUBS 0.025748f
C239 VP.n53 VSUBS 0.025748f
C240 VP.n54 VSUBS 0.047988f
C241 VP.n55 VSUBS 0.039933f
C242 VP.n56 VSUBS 1.41275f
C243 VP.n57 VSUBS 0.087724f
C244 B.n0 VSUBS 0.005021f
C245 B.n1 VSUBS 0.005021f
C246 B.n2 VSUBS 0.00794f
C247 B.n3 VSUBS 0.00794f
C248 B.n4 VSUBS 0.00794f
C249 B.n5 VSUBS 0.00794f
C250 B.n6 VSUBS 0.00794f
C251 B.n7 VSUBS 0.00794f
C252 B.n8 VSUBS 0.00794f
C253 B.n9 VSUBS 0.00794f
C254 B.n10 VSUBS 0.00794f
C255 B.n11 VSUBS 0.00794f
C256 B.n12 VSUBS 0.00794f
C257 B.n13 VSUBS 0.00794f
C258 B.n14 VSUBS 0.00794f
C259 B.n15 VSUBS 0.00794f
C260 B.n16 VSUBS 0.00794f
C261 B.n17 VSUBS 0.00794f
C262 B.n18 VSUBS 0.00794f
C263 B.n19 VSUBS 0.00794f
C264 B.n20 VSUBS 0.00794f
C265 B.n21 VSUBS 0.00794f
C266 B.n22 VSUBS 0.00794f
C267 B.n23 VSUBS 0.00794f
C268 B.n24 VSUBS 0.00794f
C269 B.n25 VSUBS 0.00794f
C270 B.n26 VSUBS 0.00794f
C271 B.n27 VSUBS 0.00794f
C272 B.n28 VSUBS 0.00794f
C273 B.n29 VSUBS 0.00794f
C274 B.n30 VSUBS 0.00794f
C275 B.n31 VSUBS 0.017321f
C276 B.n32 VSUBS 0.00794f
C277 B.n33 VSUBS 0.00794f
C278 B.n34 VSUBS 0.00794f
C279 B.n35 VSUBS 0.00794f
C280 B.n36 VSUBS 0.00794f
C281 B.n37 VSUBS 0.00794f
C282 B.n38 VSUBS 0.00794f
C283 B.n39 VSUBS 0.00794f
C284 B.n40 VSUBS 0.00794f
C285 B.n41 VSUBS 0.00794f
C286 B.n42 VSUBS 0.00794f
C287 B.n43 VSUBS 0.00794f
C288 B.n44 VSUBS 0.00794f
C289 B.n45 VSUBS 0.00794f
C290 B.n46 VSUBS 0.00794f
C291 B.n47 VSUBS 0.00794f
C292 B.n48 VSUBS 0.00794f
C293 B.n49 VSUBS 0.00794f
C294 B.n50 VSUBS 0.00794f
C295 B.n51 VSUBS 0.00794f
C296 B.n52 VSUBS 0.00794f
C297 B.n53 VSUBS 0.00794f
C298 B.n54 VSUBS 0.005488f
C299 B.n55 VSUBS 0.00794f
C300 B.t2 VSUBS 0.273201f
C301 B.t1 VSUBS 0.325597f
C302 B.t0 VSUBS 2.81335f
C303 B.n56 VSUBS 0.519891f
C304 B.n57 VSUBS 0.312953f
C305 B.n58 VSUBS 0.018397f
C306 B.n59 VSUBS 0.00794f
C307 B.n60 VSUBS 0.00794f
C308 B.n61 VSUBS 0.00794f
C309 B.n62 VSUBS 0.00794f
C310 B.t11 VSUBS 0.273204f
C311 B.t10 VSUBS 0.3256f
C312 B.t9 VSUBS 2.81335f
C313 B.n63 VSUBS 0.519888f
C314 B.n64 VSUBS 0.312949f
C315 B.n65 VSUBS 0.00794f
C316 B.n66 VSUBS 0.00794f
C317 B.n67 VSUBS 0.00794f
C318 B.n68 VSUBS 0.00794f
C319 B.n69 VSUBS 0.00794f
C320 B.n70 VSUBS 0.00794f
C321 B.n71 VSUBS 0.00794f
C322 B.n72 VSUBS 0.00794f
C323 B.n73 VSUBS 0.00794f
C324 B.n74 VSUBS 0.00794f
C325 B.n75 VSUBS 0.00794f
C326 B.n76 VSUBS 0.00794f
C327 B.n77 VSUBS 0.00794f
C328 B.n78 VSUBS 0.00794f
C329 B.n79 VSUBS 0.00794f
C330 B.n80 VSUBS 0.00794f
C331 B.n81 VSUBS 0.00794f
C332 B.n82 VSUBS 0.00794f
C333 B.n83 VSUBS 0.00794f
C334 B.n84 VSUBS 0.00794f
C335 B.n85 VSUBS 0.00794f
C336 B.n86 VSUBS 0.00794f
C337 B.n87 VSUBS 0.018307f
C338 B.n88 VSUBS 0.00794f
C339 B.n89 VSUBS 0.00794f
C340 B.n90 VSUBS 0.00794f
C341 B.n91 VSUBS 0.00794f
C342 B.n92 VSUBS 0.00794f
C343 B.n93 VSUBS 0.00794f
C344 B.n94 VSUBS 0.00794f
C345 B.n95 VSUBS 0.00794f
C346 B.n96 VSUBS 0.00794f
C347 B.n97 VSUBS 0.00794f
C348 B.n98 VSUBS 0.00794f
C349 B.n99 VSUBS 0.00794f
C350 B.n100 VSUBS 0.00794f
C351 B.n101 VSUBS 0.00794f
C352 B.n102 VSUBS 0.00794f
C353 B.n103 VSUBS 0.00794f
C354 B.n104 VSUBS 0.00794f
C355 B.n105 VSUBS 0.00794f
C356 B.n106 VSUBS 0.00794f
C357 B.n107 VSUBS 0.00794f
C358 B.n108 VSUBS 0.00794f
C359 B.n109 VSUBS 0.00794f
C360 B.n110 VSUBS 0.00794f
C361 B.n111 VSUBS 0.00794f
C362 B.n112 VSUBS 0.00794f
C363 B.n113 VSUBS 0.00794f
C364 B.n114 VSUBS 0.00794f
C365 B.n115 VSUBS 0.00794f
C366 B.n116 VSUBS 0.00794f
C367 B.n117 VSUBS 0.00794f
C368 B.n118 VSUBS 0.00794f
C369 B.n119 VSUBS 0.00794f
C370 B.n120 VSUBS 0.00794f
C371 B.n121 VSUBS 0.00794f
C372 B.n122 VSUBS 0.00794f
C373 B.n123 VSUBS 0.00794f
C374 B.n124 VSUBS 0.00794f
C375 B.n125 VSUBS 0.00794f
C376 B.n126 VSUBS 0.00794f
C377 B.n127 VSUBS 0.00794f
C378 B.n128 VSUBS 0.00794f
C379 B.n129 VSUBS 0.00794f
C380 B.n130 VSUBS 0.00794f
C381 B.n131 VSUBS 0.00794f
C382 B.n132 VSUBS 0.00794f
C383 B.n133 VSUBS 0.00794f
C384 B.n134 VSUBS 0.00794f
C385 B.n135 VSUBS 0.00794f
C386 B.n136 VSUBS 0.00794f
C387 B.n137 VSUBS 0.00794f
C388 B.n138 VSUBS 0.00794f
C389 B.n139 VSUBS 0.00794f
C390 B.n140 VSUBS 0.00794f
C391 B.n141 VSUBS 0.00794f
C392 B.n142 VSUBS 0.00794f
C393 B.n143 VSUBS 0.00794f
C394 B.n144 VSUBS 0.00794f
C395 B.n145 VSUBS 0.00794f
C396 B.n146 VSUBS 0.017321f
C397 B.n147 VSUBS 0.00794f
C398 B.n148 VSUBS 0.00794f
C399 B.n149 VSUBS 0.00794f
C400 B.n150 VSUBS 0.00794f
C401 B.n151 VSUBS 0.00794f
C402 B.n152 VSUBS 0.00794f
C403 B.n153 VSUBS 0.00794f
C404 B.n154 VSUBS 0.00794f
C405 B.n155 VSUBS 0.00794f
C406 B.n156 VSUBS 0.00794f
C407 B.n157 VSUBS 0.00794f
C408 B.n158 VSUBS 0.00794f
C409 B.n159 VSUBS 0.00794f
C410 B.n160 VSUBS 0.00794f
C411 B.n161 VSUBS 0.00794f
C412 B.n162 VSUBS 0.00794f
C413 B.n163 VSUBS 0.00794f
C414 B.n164 VSUBS 0.00794f
C415 B.n165 VSUBS 0.00794f
C416 B.n166 VSUBS 0.00794f
C417 B.n167 VSUBS 0.00794f
C418 B.n168 VSUBS 0.00794f
C419 B.n169 VSUBS 0.005488f
C420 B.n170 VSUBS 0.00794f
C421 B.n171 VSUBS 0.00794f
C422 B.n172 VSUBS 0.00794f
C423 B.n173 VSUBS 0.00794f
C424 B.n174 VSUBS 0.00794f
C425 B.t4 VSUBS 0.273201f
C426 B.t5 VSUBS 0.325597f
C427 B.t3 VSUBS 2.81335f
C428 B.n175 VSUBS 0.519891f
C429 B.n176 VSUBS 0.312953f
C430 B.n177 VSUBS 0.00794f
C431 B.n178 VSUBS 0.00794f
C432 B.n179 VSUBS 0.00794f
C433 B.n180 VSUBS 0.00794f
C434 B.n181 VSUBS 0.00794f
C435 B.n182 VSUBS 0.00794f
C436 B.n183 VSUBS 0.00794f
C437 B.n184 VSUBS 0.00794f
C438 B.n185 VSUBS 0.00794f
C439 B.n186 VSUBS 0.00794f
C440 B.n187 VSUBS 0.00794f
C441 B.n188 VSUBS 0.00794f
C442 B.n189 VSUBS 0.00794f
C443 B.n190 VSUBS 0.00794f
C444 B.n191 VSUBS 0.00794f
C445 B.n192 VSUBS 0.00794f
C446 B.n193 VSUBS 0.00794f
C447 B.n194 VSUBS 0.00794f
C448 B.n195 VSUBS 0.00794f
C449 B.n196 VSUBS 0.00794f
C450 B.n197 VSUBS 0.00794f
C451 B.n198 VSUBS 0.00794f
C452 B.n199 VSUBS 0.017321f
C453 B.n200 VSUBS 0.00794f
C454 B.n201 VSUBS 0.00794f
C455 B.n202 VSUBS 0.00794f
C456 B.n203 VSUBS 0.00794f
C457 B.n204 VSUBS 0.00794f
C458 B.n205 VSUBS 0.00794f
C459 B.n206 VSUBS 0.00794f
C460 B.n207 VSUBS 0.00794f
C461 B.n208 VSUBS 0.00794f
C462 B.n209 VSUBS 0.00794f
C463 B.n210 VSUBS 0.00794f
C464 B.n211 VSUBS 0.00794f
C465 B.n212 VSUBS 0.00794f
C466 B.n213 VSUBS 0.00794f
C467 B.n214 VSUBS 0.00794f
C468 B.n215 VSUBS 0.00794f
C469 B.n216 VSUBS 0.00794f
C470 B.n217 VSUBS 0.00794f
C471 B.n218 VSUBS 0.00794f
C472 B.n219 VSUBS 0.00794f
C473 B.n220 VSUBS 0.00794f
C474 B.n221 VSUBS 0.00794f
C475 B.n222 VSUBS 0.00794f
C476 B.n223 VSUBS 0.00794f
C477 B.n224 VSUBS 0.00794f
C478 B.n225 VSUBS 0.00794f
C479 B.n226 VSUBS 0.00794f
C480 B.n227 VSUBS 0.00794f
C481 B.n228 VSUBS 0.00794f
C482 B.n229 VSUBS 0.00794f
C483 B.n230 VSUBS 0.00794f
C484 B.n231 VSUBS 0.00794f
C485 B.n232 VSUBS 0.00794f
C486 B.n233 VSUBS 0.00794f
C487 B.n234 VSUBS 0.00794f
C488 B.n235 VSUBS 0.00794f
C489 B.n236 VSUBS 0.00794f
C490 B.n237 VSUBS 0.00794f
C491 B.n238 VSUBS 0.00794f
C492 B.n239 VSUBS 0.00794f
C493 B.n240 VSUBS 0.00794f
C494 B.n241 VSUBS 0.00794f
C495 B.n242 VSUBS 0.00794f
C496 B.n243 VSUBS 0.00794f
C497 B.n244 VSUBS 0.00794f
C498 B.n245 VSUBS 0.00794f
C499 B.n246 VSUBS 0.00794f
C500 B.n247 VSUBS 0.00794f
C501 B.n248 VSUBS 0.00794f
C502 B.n249 VSUBS 0.00794f
C503 B.n250 VSUBS 0.00794f
C504 B.n251 VSUBS 0.00794f
C505 B.n252 VSUBS 0.00794f
C506 B.n253 VSUBS 0.00794f
C507 B.n254 VSUBS 0.00794f
C508 B.n255 VSUBS 0.00794f
C509 B.n256 VSUBS 0.00794f
C510 B.n257 VSUBS 0.00794f
C511 B.n258 VSUBS 0.00794f
C512 B.n259 VSUBS 0.00794f
C513 B.n260 VSUBS 0.00794f
C514 B.n261 VSUBS 0.00794f
C515 B.n262 VSUBS 0.00794f
C516 B.n263 VSUBS 0.00794f
C517 B.n264 VSUBS 0.00794f
C518 B.n265 VSUBS 0.00794f
C519 B.n266 VSUBS 0.00794f
C520 B.n267 VSUBS 0.00794f
C521 B.n268 VSUBS 0.00794f
C522 B.n269 VSUBS 0.00794f
C523 B.n270 VSUBS 0.00794f
C524 B.n271 VSUBS 0.00794f
C525 B.n272 VSUBS 0.00794f
C526 B.n273 VSUBS 0.00794f
C527 B.n274 VSUBS 0.00794f
C528 B.n275 VSUBS 0.00794f
C529 B.n276 VSUBS 0.00794f
C530 B.n277 VSUBS 0.00794f
C531 B.n278 VSUBS 0.00794f
C532 B.n279 VSUBS 0.00794f
C533 B.n280 VSUBS 0.00794f
C534 B.n281 VSUBS 0.00794f
C535 B.n282 VSUBS 0.00794f
C536 B.n283 VSUBS 0.00794f
C537 B.n284 VSUBS 0.00794f
C538 B.n285 VSUBS 0.00794f
C539 B.n286 VSUBS 0.00794f
C540 B.n287 VSUBS 0.00794f
C541 B.n288 VSUBS 0.00794f
C542 B.n289 VSUBS 0.00794f
C543 B.n290 VSUBS 0.00794f
C544 B.n291 VSUBS 0.00794f
C545 B.n292 VSUBS 0.00794f
C546 B.n293 VSUBS 0.00794f
C547 B.n294 VSUBS 0.00794f
C548 B.n295 VSUBS 0.00794f
C549 B.n296 VSUBS 0.00794f
C550 B.n297 VSUBS 0.00794f
C551 B.n298 VSUBS 0.00794f
C552 B.n299 VSUBS 0.00794f
C553 B.n300 VSUBS 0.00794f
C554 B.n301 VSUBS 0.00794f
C555 B.n302 VSUBS 0.00794f
C556 B.n303 VSUBS 0.00794f
C557 B.n304 VSUBS 0.00794f
C558 B.n305 VSUBS 0.00794f
C559 B.n306 VSUBS 0.00794f
C560 B.n307 VSUBS 0.00794f
C561 B.n308 VSUBS 0.00794f
C562 B.n309 VSUBS 0.00794f
C563 B.n310 VSUBS 0.00794f
C564 B.n311 VSUBS 0.00794f
C565 B.n312 VSUBS 0.00794f
C566 B.n313 VSUBS 0.00794f
C567 B.n314 VSUBS 0.017321f
C568 B.n315 VSUBS 0.018644f
C569 B.n316 VSUBS 0.018644f
C570 B.n317 VSUBS 0.00794f
C571 B.n318 VSUBS 0.00794f
C572 B.n319 VSUBS 0.00794f
C573 B.n320 VSUBS 0.00794f
C574 B.n321 VSUBS 0.00794f
C575 B.n322 VSUBS 0.00794f
C576 B.n323 VSUBS 0.00794f
C577 B.n324 VSUBS 0.00794f
C578 B.n325 VSUBS 0.00794f
C579 B.n326 VSUBS 0.00794f
C580 B.n327 VSUBS 0.00794f
C581 B.n328 VSUBS 0.00794f
C582 B.n329 VSUBS 0.00794f
C583 B.n330 VSUBS 0.00794f
C584 B.n331 VSUBS 0.00794f
C585 B.n332 VSUBS 0.00794f
C586 B.n333 VSUBS 0.00794f
C587 B.n334 VSUBS 0.00794f
C588 B.n335 VSUBS 0.00794f
C589 B.n336 VSUBS 0.00794f
C590 B.n337 VSUBS 0.00794f
C591 B.n338 VSUBS 0.00794f
C592 B.n339 VSUBS 0.00794f
C593 B.n340 VSUBS 0.00794f
C594 B.n341 VSUBS 0.00794f
C595 B.n342 VSUBS 0.00794f
C596 B.n343 VSUBS 0.00794f
C597 B.n344 VSUBS 0.00794f
C598 B.n345 VSUBS 0.00794f
C599 B.n346 VSUBS 0.00794f
C600 B.n347 VSUBS 0.00794f
C601 B.n348 VSUBS 0.00794f
C602 B.n349 VSUBS 0.00794f
C603 B.n350 VSUBS 0.00794f
C604 B.n351 VSUBS 0.00794f
C605 B.n352 VSUBS 0.00794f
C606 B.n353 VSUBS 0.00794f
C607 B.n354 VSUBS 0.00794f
C608 B.n355 VSUBS 0.00794f
C609 B.n356 VSUBS 0.00794f
C610 B.n357 VSUBS 0.00794f
C611 B.n358 VSUBS 0.00794f
C612 B.n359 VSUBS 0.00794f
C613 B.n360 VSUBS 0.00794f
C614 B.n361 VSUBS 0.00794f
C615 B.n362 VSUBS 0.00794f
C616 B.n363 VSUBS 0.00794f
C617 B.n364 VSUBS 0.00794f
C618 B.n365 VSUBS 0.00794f
C619 B.n366 VSUBS 0.00794f
C620 B.n367 VSUBS 0.00794f
C621 B.n368 VSUBS 0.00794f
C622 B.n369 VSUBS 0.00794f
C623 B.n370 VSUBS 0.00794f
C624 B.n371 VSUBS 0.00794f
C625 B.n372 VSUBS 0.00794f
C626 B.n373 VSUBS 0.00794f
C627 B.n374 VSUBS 0.00794f
C628 B.n375 VSUBS 0.00794f
C629 B.n376 VSUBS 0.00794f
C630 B.n377 VSUBS 0.00794f
C631 B.n378 VSUBS 0.00794f
C632 B.n379 VSUBS 0.00794f
C633 B.n380 VSUBS 0.00794f
C634 B.n381 VSUBS 0.00794f
C635 B.n382 VSUBS 0.00794f
C636 B.n383 VSUBS 0.005488f
C637 B.n384 VSUBS 0.018397f
C638 B.n385 VSUBS 0.006422f
C639 B.n386 VSUBS 0.00794f
C640 B.n387 VSUBS 0.00794f
C641 B.n388 VSUBS 0.00794f
C642 B.n389 VSUBS 0.00794f
C643 B.n390 VSUBS 0.00794f
C644 B.n391 VSUBS 0.00794f
C645 B.n392 VSUBS 0.00794f
C646 B.n393 VSUBS 0.00794f
C647 B.n394 VSUBS 0.00794f
C648 B.n395 VSUBS 0.00794f
C649 B.n396 VSUBS 0.00794f
C650 B.t7 VSUBS 0.273204f
C651 B.t8 VSUBS 0.3256f
C652 B.t6 VSUBS 2.81335f
C653 B.n397 VSUBS 0.519888f
C654 B.n398 VSUBS 0.312949f
C655 B.n399 VSUBS 0.018397f
C656 B.n400 VSUBS 0.006422f
C657 B.n401 VSUBS 0.00794f
C658 B.n402 VSUBS 0.00794f
C659 B.n403 VSUBS 0.00794f
C660 B.n404 VSUBS 0.00794f
C661 B.n405 VSUBS 0.00794f
C662 B.n406 VSUBS 0.00794f
C663 B.n407 VSUBS 0.00794f
C664 B.n408 VSUBS 0.00794f
C665 B.n409 VSUBS 0.00794f
C666 B.n410 VSUBS 0.00794f
C667 B.n411 VSUBS 0.00794f
C668 B.n412 VSUBS 0.00794f
C669 B.n413 VSUBS 0.00794f
C670 B.n414 VSUBS 0.00794f
C671 B.n415 VSUBS 0.00794f
C672 B.n416 VSUBS 0.00794f
C673 B.n417 VSUBS 0.00794f
C674 B.n418 VSUBS 0.00794f
C675 B.n419 VSUBS 0.00794f
C676 B.n420 VSUBS 0.00794f
C677 B.n421 VSUBS 0.00794f
C678 B.n422 VSUBS 0.00794f
C679 B.n423 VSUBS 0.00794f
C680 B.n424 VSUBS 0.00794f
C681 B.n425 VSUBS 0.00794f
C682 B.n426 VSUBS 0.00794f
C683 B.n427 VSUBS 0.00794f
C684 B.n428 VSUBS 0.00794f
C685 B.n429 VSUBS 0.00794f
C686 B.n430 VSUBS 0.00794f
C687 B.n431 VSUBS 0.00794f
C688 B.n432 VSUBS 0.00794f
C689 B.n433 VSUBS 0.00794f
C690 B.n434 VSUBS 0.00794f
C691 B.n435 VSUBS 0.00794f
C692 B.n436 VSUBS 0.00794f
C693 B.n437 VSUBS 0.00794f
C694 B.n438 VSUBS 0.00794f
C695 B.n439 VSUBS 0.00794f
C696 B.n440 VSUBS 0.00794f
C697 B.n441 VSUBS 0.00794f
C698 B.n442 VSUBS 0.00794f
C699 B.n443 VSUBS 0.00794f
C700 B.n444 VSUBS 0.00794f
C701 B.n445 VSUBS 0.00794f
C702 B.n446 VSUBS 0.00794f
C703 B.n447 VSUBS 0.00794f
C704 B.n448 VSUBS 0.00794f
C705 B.n449 VSUBS 0.00794f
C706 B.n450 VSUBS 0.00794f
C707 B.n451 VSUBS 0.00794f
C708 B.n452 VSUBS 0.00794f
C709 B.n453 VSUBS 0.00794f
C710 B.n454 VSUBS 0.00794f
C711 B.n455 VSUBS 0.00794f
C712 B.n456 VSUBS 0.00794f
C713 B.n457 VSUBS 0.00794f
C714 B.n458 VSUBS 0.00794f
C715 B.n459 VSUBS 0.00794f
C716 B.n460 VSUBS 0.00794f
C717 B.n461 VSUBS 0.00794f
C718 B.n462 VSUBS 0.00794f
C719 B.n463 VSUBS 0.00794f
C720 B.n464 VSUBS 0.00794f
C721 B.n465 VSUBS 0.00794f
C722 B.n466 VSUBS 0.00794f
C723 B.n467 VSUBS 0.00794f
C724 B.n468 VSUBS 0.00794f
C725 B.n469 VSUBS 0.018644f
C726 B.n470 VSUBS 0.018644f
C727 B.n471 VSUBS 0.017321f
C728 B.n472 VSUBS 0.00794f
C729 B.n473 VSUBS 0.00794f
C730 B.n474 VSUBS 0.00794f
C731 B.n475 VSUBS 0.00794f
C732 B.n476 VSUBS 0.00794f
C733 B.n477 VSUBS 0.00794f
C734 B.n478 VSUBS 0.00794f
C735 B.n479 VSUBS 0.00794f
C736 B.n480 VSUBS 0.00794f
C737 B.n481 VSUBS 0.00794f
C738 B.n482 VSUBS 0.00794f
C739 B.n483 VSUBS 0.00794f
C740 B.n484 VSUBS 0.00794f
C741 B.n485 VSUBS 0.00794f
C742 B.n486 VSUBS 0.00794f
C743 B.n487 VSUBS 0.00794f
C744 B.n488 VSUBS 0.00794f
C745 B.n489 VSUBS 0.00794f
C746 B.n490 VSUBS 0.00794f
C747 B.n491 VSUBS 0.00794f
C748 B.n492 VSUBS 0.00794f
C749 B.n493 VSUBS 0.00794f
C750 B.n494 VSUBS 0.00794f
C751 B.n495 VSUBS 0.00794f
C752 B.n496 VSUBS 0.00794f
C753 B.n497 VSUBS 0.00794f
C754 B.n498 VSUBS 0.00794f
C755 B.n499 VSUBS 0.00794f
C756 B.n500 VSUBS 0.00794f
C757 B.n501 VSUBS 0.00794f
C758 B.n502 VSUBS 0.00794f
C759 B.n503 VSUBS 0.00794f
C760 B.n504 VSUBS 0.00794f
C761 B.n505 VSUBS 0.00794f
C762 B.n506 VSUBS 0.00794f
C763 B.n507 VSUBS 0.00794f
C764 B.n508 VSUBS 0.00794f
C765 B.n509 VSUBS 0.00794f
C766 B.n510 VSUBS 0.00794f
C767 B.n511 VSUBS 0.00794f
C768 B.n512 VSUBS 0.00794f
C769 B.n513 VSUBS 0.00794f
C770 B.n514 VSUBS 0.00794f
C771 B.n515 VSUBS 0.00794f
C772 B.n516 VSUBS 0.00794f
C773 B.n517 VSUBS 0.00794f
C774 B.n518 VSUBS 0.00794f
C775 B.n519 VSUBS 0.00794f
C776 B.n520 VSUBS 0.00794f
C777 B.n521 VSUBS 0.00794f
C778 B.n522 VSUBS 0.00794f
C779 B.n523 VSUBS 0.00794f
C780 B.n524 VSUBS 0.00794f
C781 B.n525 VSUBS 0.00794f
C782 B.n526 VSUBS 0.00794f
C783 B.n527 VSUBS 0.00794f
C784 B.n528 VSUBS 0.00794f
C785 B.n529 VSUBS 0.00794f
C786 B.n530 VSUBS 0.00794f
C787 B.n531 VSUBS 0.00794f
C788 B.n532 VSUBS 0.00794f
C789 B.n533 VSUBS 0.00794f
C790 B.n534 VSUBS 0.00794f
C791 B.n535 VSUBS 0.00794f
C792 B.n536 VSUBS 0.00794f
C793 B.n537 VSUBS 0.00794f
C794 B.n538 VSUBS 0.00794f
C795 B.n539 VSUBS 0.00794f
C796 B.n540 VSUBS 0.00794f
C797 B.n541 VSUBS 0.00794f
C798 B.n542 VSUBS 0.00794f
C799 B.n543 VSUBS 0.00794f
C800 B.n544 VSUBS 0.00794f
C801 B.n545 VSUBS 0.00794f
C802 B.n546 VSUBS 0.00794f
C803 B.n547 VSUBS 0.00794f
C804 B.n548 VSUBS 0.00794f
C805 B.n549 VSUBS 0.00794f
C806 B.n550 VSUBS 0.00794f
C807 B.n551 VSUBS 0.00794f
C808 B.n552 VSUBS 0.00794f
C809 B.n553 VSUBS 0.00794f
C810 B.n554 VSUBS 0.00794f
C811 B.n555 VSUBS 0.00794f
C812 B.n556 VSUBS 0.00794f
C813 B.n557 VSUBS 0.00794f
C814 B.n558 VSUBS 0.00794f
C815 B.n559 VSUBS 0.00794f
C816 B.n560 VSUBS 0.00794f
C817 B.n561 VSUBS 0.00794f
C818 B.n562 VSUBS 0.00794f
C819 B.n563 VSUBS 0.00794f
C820 B.n564 VSUBS 0.00794f
C821 B.n565 VSUBS 0.00794f
C822 B.n566 VSUBS 0.00794f
C823 B.n567 VSUBS 0.00794f
C824 B.n568 VSUBS 0.00794f
C825 B.n569 VSUBS 0.00794f
C826 B.n570 VSUBS 0.00794f
C827 B.n571 VSUBS 0.00794f
C828 B.n572 VSUBS 0.00794f
C829 B.n573 VSUBS 0.00794f
C830 B.n574 VSUBS 0.00794f
C831 B.n575 VSUBS 0.00794f
C832 B.n576 VSUBS 0.00794f
C833 B.n577 VSUBS 0.00794f
C834 B.n578 VSUBS 0.00794f
C835 B.n579 VSUBS 0.00794f
C836 B.n580 VSUBS 0.00794f
C837 B.n581 VSUBS 0.00794f
C838 B.n582 VSUBS 0.00794f
C839 B.n583 VSUBS 0.00794f
C840 B.n584 VSUBS 0.00794f
C841 B.n585 VSUBS 0.00794f
C842 B.n586 VSUBS 0.00794f
C843 B.n587 VSUBS 0.00794f
C844 B.n588 VSUBS 0.00794f
C845 B.n589 VSUBS 0.00794f
C846 B.n590 VSUBS 0.00794f
C847 B.n591 VSUBS 0.00794f
C848 B.n592 VSUBS 0.00794f
C849 B.n593 VSUBS 0.00794f
C850 B.n594 VSUBS 0.00794f
C851 B.n595 VSUBS 0.00794f
C852 B.n596 VSUBS 0.00794f
C853 B.n597 VSUBS 0.00794f
C854 B.n598 VSUBS 0.00794f
C855 B.n599 VSUBS 0.00794f
C856 B.n600 VSUBS 0.00794f
C857 B.n601 VSUBS 0.00794f
C858 B.n602 VSUBS 0.00794f
C859 B.n603 VSUBS 0.00794f
C860 B.n604 VSUBS 0.00794f
C861 B.n605 VSUBS 0.00794f
C862 B.n606 VSUBS 0.00794f
C863 B.n607 VSUBS 0.00794f
C864 B.n608 VSUBS 0.00794f
C865 B.n609 VSUBS 0.00794f
C866 B.n610 VSUBS 0.00794f
C867 B.n611 VSUBS 0.00794f
C868 B.n612 VSUBS 0.00794f
C869 B.n613 VSUBS 0.00794f
C870 B.n614 VSUBS 0.00794f
C871 B.n615 VSUBS 0.00794f
C872 B.n616 VSUBS 0.00794f
C873 B.n617 VSUBS 0.00794f
C874 B.n618 VSUBS 0.00794f
C875 B.n619 VSUBS 0.00794f
C876 B.n620 VSUBS 0.00794f
C877 B.n621 VSUBS 0.00794f
C878 B.n622 VSUBS 0.00794f
C879 B.n623 VSUBS 0.00794f
C880 B.n624 VSUBS 0.00794f
C881 B.n625 VSUBS 0.00794f
C882 B.n626 VSUBS 0.00794f
C883 B.n627 VSUBS 0.00794f
C884 B.n628 VSUBS 0.00794f
C885 B.n629 VSUBS 0.00794f
C886 B.n630 VSUBS 0.00794f
C887 B.n631 VSUBS 0.00794f
C888 B.n632 VSUBS 0.00794f
C889 B.n633 VSUBS 0.00794f
C890 B.n634 VSUBS 0.00794f
C891 B.n635 VSUBS 0.00794f
C892 B.n636 VSUBS 0.00794f
C893 B.n637 VSUBS 0.00794f
C894 B.n638 VSUBS 0.00794f
C895 B.n639 VSUBS 0.00794f
C896 B.n640 VSUBS 0.00794f
C897 B.n641 VSUBS 0.00794f
C898 B.n642 VSUBS 0.00794f
C899 B.n643 VSUBS 0.00794f
C900 B.n644 VSUBS 0.00794f
C901 B.n645 VSUBS 0.00794f
C902 B.n646 VSUBS 0.00794f
C903 B.n647 VSUBS 0.00794f
C904 B.n648 VSUBS 0.017321f
C905 B.n649 VSUBS 0.018644f
C906 B.n650 VSUBS 0.017657f
C907 B.n651 VSUBS 0.00794f
C908 B.n652 VSUBS 0.00794f
C909 B.n653 VSUBS 0.00794f
C910 B.n654 VSUBS 0.00794f
C911 B.n655 VSUBS 0.00794f
C912 B.n656 VSUBS 0.00794f
C913 B.n657 VSUBS 0.00794f
C914 B.n658 VSUBS 0.00794f
C915 B.n659 VSUBS 0.00794f
C916 B.n660 VSUBS 0.00794f
C917 B.n661 VSUBS 0.00794f
C918 B.n662 VSUBS 0.00794f
C919 B.n663 VSUBS 0.00794f
C920 B.n664 VSUBS 0.00794f
C921 B.n665 VSUBS 0.00794f
C922 B.n666 VSUBS 0.00794f
C923 B.n667 VSUBS 0.00794f
C924 B.n668 VSUBS 0.00794f
C925 B.n669 VSUBS 0.00794f
C926 B.n670 VSUBS 0.00794f
C927 B.n671 VSUBS 0.00794f
C928 B.n672 VSUBS 0.00794f
C929 B.n673 VSUBS 0.00794f
C930 B.n674 VSUBS 0.00794f
C931 B.n675 VSUBS 0.00794f
C932 B.n676 VSUBS 0.00794f
C933 B.n677 VSUBS 0.00794f
C934 B.n678 VSUBS 0.00794f
C935 B.n679 VSUBS 0.00794f
C936 B.n680 VSUBS 0.00794f
C937 B.n681 VSUBS 0.00794f
C938 B.n682 VSUBS 0.00794f
C939 B.n683 VSUBS 0.00794f
C940 B.n684 VSUBS 0.00794f
C941 B.n685 VSUBS 0.00794f
C942 B.n686 VSUBS 0.00794f
C943 B.n687 VSUBS 0.00794f
C944 B.n688 VSUBS 0.00794f
C945 B.n689 VSUBS 0.00794f
C946 B.n690 VSUBS 0.00794f
C947 B.n691 VSUBS 0.00794f
C948 B.n692 VSUBS 0.00794f
C949 B.n693 VSUBS 0.00794f
C950 B.n694 VSUBS 0.00794f
C951 B.n695 VSUBS 0.00794f
C952 B.n696 VSUBS 0.00794f
C953 B.n697 VSUBS 0.00794f
C954 B.n698 VSUBS 0.00794f
C955 B.n699 VSUBS 0.00794f
C956 B.n700 VSUBS 0.00794f
C957 B.n701 VSUBS 0.00794f
C958 B.n702 VSUBS 0.00794f
C959 B.n703 VSUBS 0.00794f
C960 B.n704 VSUBS 0.00794f
C961 B.n705 VSUBS 0.00794f
C962 B.n706 VSUBS 0.00794f
C963 B.n707 VSUBS 0.00794f
C964 B.n708 VSUBS 0.00794f
C965 B.n709 VSUBS 0.00794f
C966 B.n710 VSUBS 0.00794f
C967 B.n711 VSUBS 0.00794f
C968 B.n712 VSUBS 0.00794f
C969 B.n713 VSUBS 0.00794f
C970 B.n714 VSUBS 0.00794f
C971 B.n715 VSUBS 0.00794f
C972 B.n716 VSUBS 0.00794f
C973 B.n717 VSUBS 0.005488f
C974 B.n718 VSUBS 0.018397f
C975 B.n719 VSUBS 0.006422f
C976 B.n720 VSUBS 0.00794f
C977 B.n721 VSUBS 0.00794f
C978 B.n722 VSUBS 0.00794f
C979 B.n723 VSUBS 0.00794f
C980 B.n724 VSUBS 0.00794f
C981 B.n725 VSUBS 0.00794f
C982 B.n726 VSUBS 0.00794f
C983 B.n727 VSUBS 0.00794f
C984 B.n728 VSUBS 0.00794f
C985 B.n729 VSUBS 0.00794f
C986 B.n730 VSUBS 0.00794f
C987 B.n731 VSUBS 0.006422f
C988 B.n732 VSUBS 0.00794f
C989 B.n733 VSUBS 0.00794f
C990 B.n734 VSUBS 0.00794f
C991 B.n735 VSUBS 0.00794f
C992 B.n736 VSUBS 0.00794f
C993 B.n737 VSUBS 0.00794f
C994 B.n738 VSUBS 0.00794f
C995 B.n739 VSUBS 0.00794f
C996 B.n740 VSUBS 0.00794f
C997 B.n741 VSUBS 0.00794f
C998 B.n742 VSUBS 0.00794f
C999 B.n743 VSUBS 0.00794f
C1000 B.n744 VSUBS 0.00794f
C1001 B.n745 VSUBS 0.00794f
C1002 B.n746 VSUBS 0.00794f
C1003 B.n747 VSUBS 0.00794f
C1004 B.n748 VSUBS 0.00794f
C1005 B.n749 VSUBS 0.00794f
C1006 B.n750 VSUBS 0.00794f
C1007 B.n751 VSUBS 0.00794f
C1008 B.n752 VSUBS 0.00794f
C1009 B.n753 VSUBS 0.00794f
C1010 B.n754 VSUBS 0.00794f
C1011 B.n755 VSUBS 0.00794f
C1012 B.n756 VSUBS 0.00794f
C1013 B.n757 VSUBS 0.00794f
C1014 B.n758 VSUBS 0.00794f
C1015 B.n759 VSUBS 0.00794f
C1016 B.n760 VSUBS 0.00794f
C1017 B.n761 VSUBS 0.00794f
C1018 B.n762 VSUBS 0.00794f
C1019 B.n763 VSUBS 0.00794f
C1020 B.n764 VSUBS 0.00794f
C1021 B.n765 VSUBS 0.00794f
C1022 B.n766 VSUBS 0.00794f
C1023 B.n767 VSUBS 0.00794f
C1024 B.n768 VSUBS 0.00794f
C1025 B.n769 VSUBS 0.00794f
C1026 B.n770 VSUBS 0.00794f
C1027 B.n771 VSUBS 0.00794f
C1028 B.n772 VSUBS 0.00794f
C1029 B.n773 VSUBS 0.00794f
C1030 B.n774 VSUBS 0.00794f
C1031 B.n775 VSUBS 0.00794f
C1032 B.n776 VSUBS 0.00794f
C1033 B.n777 VSUBS 0.00794f
C1034 B.n778 VSUBS 0.00794f
C1035 B.n779 VSUBS 0.00794f
C1036 B.n780 VSUBS 0.00794f
C1037 B.n781 VSUBS 0.00794f
C1038 B.n782 VSUBS 0.00794f
C1039 B.n783 VSUBS 0.00794f
C1040 B.n784 VSUBS 0.00794f
C1041 B.n785 VSUBS 0.00794f
C1042 B.n786 VSUBS 0.00794f
C1043 B.n787 VSUBS 0.00794f
C1044 B.n788 VSUBS 0.00794f
C1045 B.n789 VSUBS 0.00794f
C1046 B.n790 VSUBS 0.00794f
C1047 B.n791 VSUBS 0.00794f
C1048 B.n792 VSUBS 0.00794f
C1049 B.n793 VSUBS 0.00794f
C1050 B.n794 VSUBS 0.00794f
C1051 B.n795 VSUBS 0.00794f
C1052 B.n796 VSUBS 0.00794f
C1053 B.n797 VSUBS 0.00794f
C1054 B.n798 VSUBS 0.00794f
C1055 B.n799 VSUBS 0.00794f
C1056 B.n800 VSUBS 0.018644f
C1057 B.n801 VSUBS 0.018644f
C1058 B.n802 VSUBS 0.017321f
C1059 B.n803 VSUBS 0.00794f
C1060 B.n804 VSUBS 0.00794f
C1061 B.n805 VSUBS 0.00794f
C1062 B.n806 VSUBS 0.00794f
C1063 B.n807 VSUBS 0.00794f
C1064 B.n808 VSUBS 0.00794f
C1065 B.n809 VSUBS 0.00794f
C1066 B.n810 VSUBS 0.00794f
C1067 B.n811 VSUBS 0.00794f
C1068 B.n812 VSUBS 0.00794f
C1069 B.n813 VSUBS 0.00794f
C1070 B.n814 VSUBS 0.00794f
C1071 B.n815 VSUBS 0.00794f
C1072 B.n816 VSUBS 0.00794f
C1073 B.n817 VSUBS 0.00794f
C1074 B.n818 VSUBS 0.00794f
C1075 B.n819 VSUBS 0.00794f
C1076 B.n820 VSUBS 0.00794f
C1077 B.n821 VSUBS 0.00794f
C1078 B.n822 VSUBS 0.00794f
C1079 B.n823 VSUBS 0.00794f
C1080 B.n824 VSUBS 0.00794f
C1081 B.n825 VSUBS 0.00794f
C1082 B.n826 VSUBS 0.00794f
C1083 B.n827 VSUBS 0.00794f
C1084 B.n828 VSUBS 0.00794f
C1085 B.n829 VSUBS 0.00794f
C1086 B.n830 VSUBS 0.00794f
C1087 B.n831 VSUBS 0.00794f
C1088 B.n832 VSUBS 0.00794f
C1089 B.n833 VSUBS 0.00794f
C1090 B.n834 VSUBS 0.00794f
C1091 B.n835 VSUBS 0.00794f
C1092 B.n836 VSUBS 0.00794f
C1093 B.n837 VSUBS 0.00794f
C1094 B.n838 VSUBS 0.00794f
C1095 B.n839 VSUBS 0.00794f
C1096 B.n840 VSUBS 0.00794f
C1097 B.n841 VSUBS 0.00794f
C1098 B.n842 VSUBS 0.00794f
C1099 B.n843 VSUBS 0.00794f
C1100 B.n844 VSUBS 0.00794f
C1101 B.n845 VSUBS 0.00794f
C1102 B.n846 VSUBS 0.00794f
C1103 B.n847 VSUBS 0.00794f
C1104 B.n848 VSUBS 0.00794f
C1105 B.n849 VSUBS 0.00794f
C1106 B.n850 VSUBS 0.00794f
C1107 B.n851 VSUBS 0.00794f
C1108 B.n852 VSUBS 0.00794f
C1109 B.n853 VSUBS 0.00794f
C1110 B.n854 VSUBS 0.00794f
C1111 B.n855 VSUBS 0.00794f
C1112 B.n856 VSUBS 0.00794f
C1113 B.n857 VSUBS 0.00794f
C1114 B.n858 VSUBS 0.00794f
C1115 B.n859 VSUBS 0.00794f
C1116 B.n860 VSUBS 0.00794f
C1117 B.n861 VSUBS 0.00794f
C1118 B.n862 VSUBS 0.00794f
C1119 B.n863 VSUBS 0.00794f
C1120 B.n864 VSUBS 0.00794f
C1121 B.n865 VSUBS 0.00794f
C1122 B.n866 VSUBS 0.00794f
C1123 B.n867 VSUBS 0.00794f
C1124 B.n868 VSUBS 0.00794f
C1125 B.n869 VSUBS 0.00794f
C1126 B.n870 VSUBS 0.00794f
C1127 B.n871 VSUBS 0.00794f
C1128 B.n872 VSUBS 0.00794f
C1129 B.n873 VSUBS 0.00794f
C1130 B.n874 VSUBS 0.00794f
C1131 B.n875 VSUBS 0.00794f
C1132 B.n876 VSUBS 0.00794f
C1133 B.n877 VSUBS 0.00794f
C1134 B.n878 VSUBS 0.00794f
C1135 B.n879 VSUBS 0.00794f
C1136 B.n880 VSUBS 0.00794f
C1137 B.n881 VSUBS 0.00794f
C1138 B.n882 VSUBS 0.00794f
C1139 B.n883 VSUBS 0.00794f
C1140 B.n884 VSUBS 0.00794f
C1141 B.n885 VSUBS 0.00794f
C1142 B.n886 VSUBS 0.00794f
C1143 B.n887 VSUBS 0.00794f
C1144 B.n888 VSUBS 0.00794f
C1145 B.n889 VSUBS 0.00794f
C1146 B.n890 VSUBS 0.00794f
C1147 B.n891 VSUBS 0.01798f
C1148 VDD2.n0 VSUBS 0.030048f
C1149 VDD2.n1 VSUBS 0.02819f
C1150 VDD2.n2 VSUBS 0.015148f
C1151 VDD2.n3 VSUBS 0.035804f
C1152 VDD2.n4 VSUBS 0.016039f
C1153 VDD2.n5 VSUBS 0.02819f
C1154 VDD2.n6 VSUBS 0.015148f
C1155 VDD2.n7 VSUBS 0.035804f
C1156 VDD2.n8 VSUBS 0.016039f
C1157 VDD2.n9 VSUBS 0.02819f
C1158 VDD2.n10 VSUBS 0.015148f
C1159 VDD2.n11 VSUBS 0.035804f
C1160 VDD2.n12 VSUBS 0.016039f
C1161 VDD2.n13 VSUBS 0.02819f
C1162 VDD2.n14 VSUBS 0.015148f
C1163 VDD2.n15 VSUBS 0.035804f
C1164 VDD2.n16 VSUBS 0.016039f
C1165 VDD2.n17 VSUBS 0.02819f
C1166 VDD2.n18 VSUBS 0.015148f
C1167 VDD2.n19 VSUBS 0.035804f
C1168 VDD2.n20 VSUBS 0.016039f
C1169 VDD2.n21 VSUBS 1.58625f
C1170 VDD2.n22 VSUBS 0.015148f
C1171 VDD2.t0 VSUBS 0.076534f
C1172 VDD2.n23 VSUBS 0.184828f
C1173 VDD2.n24 VSUBS 0.022777f
C1174 VDD2.n25 VSUBS 0.026853f
C1175 VDD2.n26 VSUBS 0.035804f
C1176 VDD2.n27 VSUBS 0.016039f
C1177 VDD2.n28 VSUBS 0.015148f
C1178 VDD2.n29 VSUBS 0.02819f
C1179 VDD2.n30 VSUBS 0.02819f
C1180 VDD2.n31 VSUBS 0.015148f
C1181 VDD2.n32 VSUBS 0.016039f
C1182 VDD2.n33 VSUBS 0.035804f
C1183 VDD2.n34 VSUBS 0.035804f
C1184 VDD2.n35 VSUBS 0.016039f
C1185 VDD2.n36 VSUBS 0.015148f
C1186 VDD2.n37 VSUBS 0.02819f
C1187 VDD2.n38 VSUBS 0.02819f
C1188 VDD2.n39 VSUBS 0.015148f
C1189 VDD2.n40 VSUBS 0.016039f
C1190 VDD2.n41 VSUBS 0.035804f
C1191 VDD2.n42 VSUBS 0.035804f
C1192 VDD2.n43 VSUBS 0.016039f
C1193 VDD2.n44 VSUBS 0.015148f
C1194 VDD2.n45 VSUBS 0.02819f
C1195 VDD2.n46 VSUBS 0.02819f
C1196 VDD2.n47 VSUBS 0.015148f
C1197 VDD2.n48 VSUBS 0.016039f
C1198 VDD2.n49 VSUBS 0.035804f
C1199 VDD2.n50 VSUBS 0.035804f
C1200 VDD2.n51 VSUBS 0.016039f
C1201 VDD2.n52 VSUBS 0.015148f
C1202 VDD2.n53 VSUBS 0.02819f
C1203 VDD2.n54 VSUBS 0.02819f
C1204 VDD2.n55 VSUBS 0.015148f
C1205 VDD2.n56 VSUBS 0.016039f
C1206 VDD2.n57 VSUBS 0.035804f
C1207 VDD2.n58 VSUBS 0.035804f
C1208 VDD2.n59 VSUBS 0.016039f
C1209 VDD2.n60 VSUBS 0.015148f
C1210 VDD2.n61 VSUBS 0.02819f
C1211 VDD2.n62 VSUBS 0.02819f
C1212 VDD2.n63 VSUBS 0.015148f
C1213 VDD2.n64 VSUBS 0.016039f
C1214 VDD2.n65 VSUBS 0.035804f
C1215 VDD2.n66 VSUBS 0.088353f
C1216 VDD2.n67 VSUBS 0.016039f
C1217 VDD2.n68 VSUBS 0.029747f
C1218 VDD2.n69 VSUBS 0.070165f
C1219 VDD2.n70 VSUBS 0.102339f
C1220 VDD2.t4 VSUBS 0.296944f
C1221 VDD2.t1 VSUBS 0.296944f
C1222 VDD2.n71 VSUBS 2.38957f
C1223 VDD2.n72 VSUBS 4.08105f
C1224 VDD2.n73 VSUBS 0.030048f
C1225 VDD2.n74 VSUBS 0.02819f
C1226 VDD2.n75 VSUBS 0.015148f
C1227 VDD2.n76 VSUBS 0.035804f
C1228 VDD2.n77 VSUBS 0.016039f
C1229 VDD2.n78 VSUBS 0.02819f
C1230 VDD2.n79 VSUBS 0.015148f
C1231 VDD2.n80 VSUBS 0.035804f
C1232 VDD2.n81 VSUBS 0.016039f
C1233 VDD2.n82 VSUBS 0.02819f
C1234 VDD2.n83 VSUBS 0.015148f
C1235 VDD2.n84 VSUBS 0.035804f
C1236 VDD2.n85 VSUBS 0.016039f
C1237 VDD2.n86 VSUBS 0.02819f
C1238 VDD2.n87 VSUBS 0.015148f
C1239 VDD2.n88 VSUBS 0.035804f
C1240 VDD2.n89 VSUBS 0.016039f
C1241 VDD2.n90 VSUBS 0.02819f
C1242 VDD2.n91 VSUBS 0.015148f
C1243 VDD2.n92 VSUBS 0.035804f
C1244 VDD2.n93 VSUBS 0.016039f
C1245 VDD2.n94 VSUBS 1.58625f
C1246 VDD2.n95 VSUBS 0.015148f
C1247 VDD2.t5 VSUBS 0.076534f
C1248 VDD2.n96 VSUBS 0.184828f
C1249 VDD2.n97 VSUBS 0.022777f
C1250 VDD2.n98 VSUBS 0.026853f
C1251 VDD2.n99 VSUBS 0.035804f
C1252 VDD2.n100 VSUBS 0.016039f
C1253 VDD2.n101 VSUBS 0.015148f
C1254 VDD2.n102 VSUBS 0.02819f
C1255 VDD2.n103 VSUBS 0.02819f
C1256 VDD2.n104 VSUBS 0.015148f
C1257 VDD2.n105 VSUBS 0.016039f
C1258 VDD2.n106 VSUBS 0.035804f
C1259 VDD2.n107 VSUBS 0.035804f
C1260 VDD2.n108 VSUBS 0.016039f
C1261 VDD2.n109 VSUBS 0.015148f
C1262 VDD2.n110 VSUBS 0.02819f
C1263 VDD2.n111 VSUBS 0.02819f
C1264 VDD2.n112 VSUBS 0.015148f
C1265 VDD2.n113 VSUBS 0.016039f
C1266 VDD2.n114 VSUBS 0.035804f
C1267 VDD2.n115 VSUBS 0.035804f
C1268 VDD2.n116 VSUBS 0.016039f
C1269 VDD2.n117 VSUBS 0.015148f
C1270 VDD2.n118 VSUBS 0.02819f
C1271 VDD2.n119 VSUBS 0.02819f
C1272 VDD2.n120 VSUBS 0.015148f
C1273 VDD2.n121 VSUBS 0.016039f
C1274 VDD2.n122 VSUBS 0.035804f
C1275 VDD2.n123 VSUBS 0.035804f
C1276 VDD2.n124 VSUBS 0.016039f
C1277 VDD2.n125 VSUBS 0.015148f
C1278 VDD2.n126 VSUBS 0.02819f
C1279 VDD2.n127 VSUBS 0.02819f
C1280 VDD2.n128 VSUBS 0.015148f
C1281 VDD2.n129 VSUBS 0.016039f
C1282 VDD2.n130 VSUBS 0.035804f
C1283 VDD2.n131 VSUBS 0.035804f
C1284 VDD2.n132 VSUBS 0.016039f
C1285 VDD2.n133 VSUBS 0.015148f
C1286 VDD2.n134 VSUBS 0.02819f
C1287 VDD2.n135 VSUBS 0.02819f
C1288 VDD2.n136 VSUBS 0.015148f
C1289 VDD2.n137 VSUBS 0.016039f
C1290 VDD2.n138 VSUBS 0.035804f
C1291 VDD2.n139 VSUBS 0.088353f
C1292 VDD2.n140 VSUBS 0.016039f
C1293 VDD2.n141 VSUBS 0.029747f
C1294 VDD2.n142 VSUBS 0.070165f
C1295 VDD2.n143 VSUBS 0.086792f
C1296 VDD2.n144 VSUBS 3.43742f
C1297 VDD2.t2 VSUBS 0.296944f
C1298 VDD2.t3 VSUBS 0.296944f
C1299 VDD2.n145 VSUBS 2.38952f
C1300 VTAIL.t7 VSUBS 0.313448f
C1301 VTAIL.t11 VSUBS 0.313448f
C1302 VTAIL.n0 VSUBS 2.35437f
C1303 VTAIL.n1 VSUBS 0.982466f
C1304 VTAIL.n2 VSUBS 0.031718f
C1305 VTAIL.n3 VSUBS 0.029756f
C1306 VTAIL.n4 VSUBS 0.01599f
C1307 VTAIL.n5 VSUBS 0.037794f
C1308 VTAIL.n6 VSUBS 0.01693f
C1309 VTAIL.n7 VSUBS 0.029756f
C1310 VTAIL.n8 VSUBS 0.01599f
C1311 VTAIL.n9 VSUBS 0.037794f
C1312 VTAIL.n10 VSUBS 0.01693f
C1313 VTAIL.n11 VSUBS 0.029756f
C1314 VTAIL.n12 VSUBS 0.01599f
C1315 VTAIL.n13 VSUBS 0.037794f
C1316 VTAIL.n14 VSUBS 0.01693f
C1317 VTAIL.n15 VSUBS 0.029756f
C1318 VTAIL.n16 VSUBS 0.01599f
C1319 VTAIL.n17 VSUBS 0.037794f
C1320 VTAIL.n18 VSUBS 0.01693f
C1321 VTAIL.n19 VSUBS 0.029756f
C1322 VTAIL.n20 VSUBS 0.01599f
C1323 VTAIL.n21 VSUBS 0.037794f
C1324 VTAIL.n22 VSUBS 0.01693f
C1325 VTAIL.n23 VSUBS 1.67442f
C1326 VTAIL.n24 VSUBS 0.01599f
C1327 VTAIL.t5 VSUBS 0.080788f
C1328 VTAIL.n25 VSUBS 0.195101f
C1329 VTAIL.n26 VSUBS 0.024043f
C1330 VTAIL.n27 VSUBS 0.028346f
C1331 VTAIL.n28 VSUBS 0.037794f
C1332 VTAIL.n29 VSUBS 0.01693f
C1333 VTAIL.n30 VSUBS 0.01599f
C1334 VTAIL.n31 VSUBS 0.029756f
C1335 VTAIL.n32 VSUBS 0.029756f
C1336 VTAIL.n33 VSUBS 0.01599f
C1337 VTAIL.n34 VSUBS 0.01693f
C1338 VTAIL.n35 VSUBS 0.037794f
C1339 VTAIL.n36 VSUBS 0.037794f
C1340 VTAIL.n37 VSUBS 0.01693f
C1341 VTAIL.n38 VSUBS 0.01599f
C1342 VTAIL.n39 VSUBS 0.029756f
C1343 VTAIL.n40 VSUBS 0.029756f
C1344 VTAIL.n41 VSUBS 0.01599f
C1345 VTAIL.n42 VSUBS 0.01693f
C1346 VTAIL.n43 VSUBS 0.037794f
C1347 VTAIL.n44 VSUBS 0.037794f
C1348 VTAIL.n45 VSUBS 0.01693f
C1349 VTAIL.n46 VSUBS 0.01599f
C1350 VTAIL.n47 VSUBS 0.029756f
C1351 VTAIL.n48 VSUBS 0.029756f
C1352 VTAIL.n49 VSUBS 0.01599f
C1353 VTAIL.n50 VSUBS 0.01693f
C1354 VTAIL.n51 VSUBS 0.037794f
C1355 VTAIL.n52 VSUBS 0.037794f
C1356 VTAIL.n53 VSUBS 0.01693f
C1357 VTAIL.n54 VSUBS 0.01599f
C1358 VTAIL.n55 VSUBS 0.029756f
C1359 VTAIL.n56 VSUBS 0.029756f
C1360 VTAIL.n57 VSUBS 0.01599f
C1361 VTAIL.n58 VSUBS 0.01693f
C1362 VTAIL.n59 VSUBS 0.037794f
C1363 VTAIL.n60 VSUBS 0.037794f
C1364 VTAIL.n61 VSUBS 0.01693f
C1365 VTAIL.n62 VSUBS 0.01599f
C1366 VTAIL.n63 VSUBS 0.029756f
C1367 VTAIL.n64 VSUBS 0.029756f
C1368 VTAIL.n65 VSUBS 0.01599f
C1369 VTAIL.n66 VSUBS 0.01693f
C1370 VTAIL.n67 VSUBS 0.037794f
C1371 VTAIL.n68 VSUBS 0.093264f
C1372 VTAIL.n69 VSUBS 0.01693f
C1373 VTAIL.n70 VSUBS 0.0314f
C1374 VTAIL.n71 VSUBS 0.074065f
C1375 VTAIL.n72 VSUBS 0.071108f
C1376 VTAIL.n73 VSUBS 0.610307f
C1377 VTAIL.t4 VSUBS 0.313448f
C1378 VTAIL.t2 VSUBS 0.313448f
C1379 VTAIL.n74 VSUBS 2.35437f
C1380 VTAIL.n75 VSUBS 3.24315f
C1381 VTAIL.t9 VSUBS 0.313448f
C1382 VTAIL.t6 VSUBS 0.313448f
C1383 VTAIL.n76 VSUBS 2.35438f
C1384 VTAIL.n77 VSUBS 3.24313f
C1385 VTAIL.n78 VSUBS 0.031718f
C1386 VTAIL.n79 VSUBS 0.029756f
C1387 VTAIL.n80 VSUBS 0.01599f
C1388 VTAIL.n81 VSUBS 0.037794f
C1389 VTAIL.n82 VSUBS 0.01693f
C1390 VTAIL.n83 VSUBS 0.029756f
C1391 VTAIL.n84 VSUBS 0.01599f
C1392 VTAIL.n85 VSUBS 0.037794f
C1393 VTAIL.n86 VSUBS 0.01693f
C1394 VTAIL.n87 VSUBS 0.029756f
C1395 VTAIL.n88 VSUBS 0.01599f
C1396 VTAIL.n89 VSUBS 0.037794f
C1397 VTAIL.n90 VSUBS 0.01693f
C1398 VTAIL.n91 VSUBS 0.029756f
C1399 VTAIL.n92 VSUBS 0.01599f
C1400 VTAIL.n93 VSUBS 0.037794f
C1401 VTAIL.n94 VSUBS 0.01693f
C1402 VTAIL.n95 VSUBS 0.029756f
C1403 VTAIL.n96 VSUBS 0.01599f
C1404 VTAIL.n97 VSUBS 0.037794f
C1405 VTAIL.n98 VSUBS 0.01693f
C1406 VTAIL.n99 VSUBS 1.67442f
C1407 VTAIL.n100 VSUBS 0.01599f
C1408 VTAIL.t8 VSUBS 0.080787f
C1409 VTAIL.n101 VSUBS 0.195101f
C1410 VTAIL.n102 VSUBS 0.024043f
C1411 VTAIL.n103 VSUBS 0.028346f
C1412 VTAIL.n104 VSUBS 0.037794f
C1413 VTAIL.n105 VSUBS 0.01693f
C1414 VTAIL.n106 VSUBS 0.01599f
C1415 VTAIL.n107 VSUBS 0.029756f
C1416 VTAIL.n108 VSUBS 0.029756f
C1417 VTAIL.n109 VSUBS 0.01599f
C1418 VTAIL.n110 VSUBS 0.01693f
C1419 VTAIL.n111 VSUBS 0.037794f
C1420 VTAIL.n112 VSUBS 0.037794f
C1421 VTAIL.n113 VSUBS 0.01693f
C1422 VTAIL.n114 VSUBS 0.01599f
C1423 VTAIL.n115 VSUBS 0.029756f
C1424 VTAIL.n116 VSUBS 0.029756f
C1425 VTAIL.n117 VSUBS 0.01599f
C1426 VTAIL.n118 VSUBS 0.01693f
C1427 VTAIL.n119 VSUBS 0.037794f
C1428 VTAIL.n120 VSUBS 0.037794f
C1429 VTAIL.n121 VSUBS 0.01693f
C1430 VTAIL.n122 VSUBS 0.01599f
C1431 VTAIL.n123 VSUBS 0.029756f
C1432 VTAIL.n124 VSUBS 0.029756f
C1433 VTAIL.n125 VSUBS 0.01599f
C1434 VTAIL.n126 VSUBS 0.01693f
C1435 VTAIL.n127 VSUBS 0.037794f
C1436 VTAIL.n128 VSUBS 0.037794f
C1437 VTAIL.n129 VSUBS 0.01693f
C1438 VTAIL.n130 VSUBS 0.01599f
C1439 VTAIL.n131 VSUBS 0.029756f
C1440 VTAIL.n132 VSUBS 0.029756f
C1441 VTAIL.n133 VSUBS 0.01599f
C1442 VTAIL.n134 VSUBS 0.01693f
C1443 VTAIL.n135 VSUBS 0.037794f
C1444 VTAIL.n136 VSUBS 0.037794f
C1445 VTAIL.n137 VSUBS 0.01693f
C1446 VTAIL.n138 VSUBS 0.01599f
C1447 VTAIL.n139 VSUBS 0.029756f
C1448 VTAIL.n140 VSUBS 0.029756f
C1449 VTAIL.n141 VSUBS 0.01599f
C1450 VTAIL.n142 VSUBS 0.01693f
C1451 VTAIL.n143 VSUBS 0.037794f
C1452 VTAIL.n144 VSUBS 0.093264f
C1453 VTAIL.n145 VSUBS 0.01693f
C1454 VTAIL.n146 VSUBS 0.0314f
C1455 VTAIL.n147 VSUBS 0.074065f
C1456 VTAIL.n148 VSUBS 0.071108f
C1457 VTAIL.n149 VSUBS 0.610307f
C1458 VTAIL.t1 VSUBS 0.313448f
C1459 VTAIL.t3 VSUBS 0.313448f
C1460 VTAIL.n150 VSUBS 2.35438f
C1461 VTAIL.n151 VSUBS 1.2453f
C1462 VTAIL.n152 VSUBS 0.031718f
C1463 VTAIL.n153 VSUBS 0.029756f
C1464 VTAIL.n154 VSUBS 0.01599f
C1465 VTAIL.n155 VSUBS 0.037794f
C1466 VTAIL.n156 VSUBS 0.01693f
C1467 VTAIL.n157 VSUBS 0.029756f
C1468 VTAIL.n158 VSUBS 0.01599f
C1469 VTAIL.n159 VSUBS 0.037794f
C1470 VTAIL.n160 VSUBS 0.01693f
C1471 VTAIL.n161 VSUBS 0.029756f
C1472 VTAIL.n162 VSUBS 0.01599f
C1473 VTAIL.n163 VSUBS 0.037794f
C1474 VTAIL.n164 VSUBS 0.01693f
C1475 VTAIL.n165 VSUBS 0.029756f
C1476 VTAIL.n166 VSUBS 0.01599f
C1477 VTAIL.n167 VSUBS 0.037794f
C1478 VTAIL.n168 VSUBS 0.01693f
C1479 VTAIL.n169 VSUBS 0.029756f
C1480 VTAIL.n170 VSUBS 0.01599f
C1481 VTAIL.n171 VSUBS 0.037794f
C1482 VTAIL.n172 VSUBS 0.01693f
C1483 VTAIL.n173 VSUBS 1.67442f
C1484 VTAIL.n174 VSUBS 0.01599f
C1485 VTAIL.t0 VSUBS 0.080787f
C1486 VTAIL.n175 VSUBS 0.195101f
C1487 VTAIL.n176 VSUBS 0.024043f
C1488 VTAIL.n177 VSUBS 0.028346f
C1489 VTAIL.n178 VSUBS 0.037794f
C1490 VTAIL.n179 VSUBS 0.01693f
C1491 VTAIL.n180 VSUBS 0.01599f
C1492 VTAIL.n181 VSUBS 0.029756f
C1493 VTAIL.n182 VSUBS 0.029756f
C1494 VTAIL.n183 VSUBS 0.01599f
C1495 VTAIL.n184 VSUBS 0.01693f
C1496 VTAIL.n185 VSUBS 0.037794f
C1497 VTAIL.n186 VSUBS 0.037794f
C1498 VTAIL.n187 VSUBS 0.01693f
C1499 VTAIL.n188 VSUBS 0.01599f
C1500 VTAIL.n189 VSUBS 0.029756f
C1501 VTAIL.n190 VSUBS 0.029756f
C1502 VTAIL.n191 VSUBS 0.01599f
C1503 VTAIL.n192 VSUBS 0.01693f
C1504 VTAIL.n193 VSUBS 0.037794f
C1505 VTAIL.n194 VSUBS 0.037794f
C1506 VTAIL.n195 VSUBS 0.01693f
C1507 VTAIL.n196 VSUBS 0.01599f
C1508 VTAIL.n197 VSUBS 0.029756f
C1509 VTAIL.n198 VSUBS 0.029756f
C1510 VTAIL.n199 VSUBS 0.01599f
C1511 VTAIL.n200 VSUBS 0.01693f
C1512 VTAIL.n201 VSUBS 0.037794f
C1513 VTAIL.n202 VSUBS 0.037794f
C1514 VTAIL.n203 VSUBS 0.01693f
C1515 VTAIL.n204 VSUBS 0.01599f
C1516 VTAIL.n205 VSUBS 0.029756f
C1517 VTAIL.n206 VSUBS 0.029756f
C1518 VTAIL.n207 VSUBS 0.01599f
C1519 VTAIL.n208 VSUBS 0.01693f
C1520 VTAIL.n209 VSUBS 0.037794f
C1521 VTAIL.n210 VSUBS 0.037794f
C1522 VTAIL.n211 VSUBS 0.01693f
C1523 VTAIL.n212 VSUBS 0.01599f
C1524 VTAIL.n213 VSUBS 0.029756f
C1525 VTAIL.n214 VSUBS 0.029756f
C1526 VTAIL.n215 VSUBS 0.01599f
C1527 VTAIL.n216 VSUBS 0.01693f
C1528 VTAIL.n217 VSUBS 0.037794f
C1529 VTAIL.n218 VSUBS 0.093264f
C1530 VTAIL.n219 VSUBS 0.01693f
C1531 VTAIL.n220 VSUBS 0.0314f
C1532 VTAIL.n221 VSUBS 0.074065f
C1533 VTAIL.n222 VSUBS 0.071108f
C1534 VTAIL.n223 VSUBS 2.25024f
C1535 VTAIL.n224 VSUBS 0.031718f
C1536 VTAIL.n225 VSUBS 0.029756f
C1537 VTAIL.n226 VSUBS 0.01599f
C1538 VTAIL.n227 VSUBS 0.037794f
C1539 VTAIL.n228 VSUBS 0.01693f
C1540 VTAIL.n229 VSUBS 0.029756f
C1541 VTAIL.n230 VSUBS 0.01599f
C1542 VTAIL.n231 VSUBS 0.037794f
C1543 VTAIL.n232 VSUBS 0.01693f
C1544 VTAIL.n233 VSUBS 0.029756f
C1545 VTAIL.n234 VSUBS 0.01599f
C1546 VTAIL.n235 VSUBS 0.037794f
C1547 VTAIL.n236 VSUBS 0.01693f
C1548 VTAIL.n237 VSUBS 0.029756f
C1549 VTAIL.n238 VSUBS 0.01599f
C1550 VTAIL.n239 VSUBS 0.037794f
C1551 VTAIL.n240 VSUBS 0.01693f
C1552 VTAIL.n241 VSUBS 0.029756f
C1553 VTAIL.n242 VSUBS 0.01599f
C1554 VTAIL.n243 VSUBS 0.037794f
C1555 VTAIL.n244 VSUBS 0.01693f
C1556 VTAIL.n245 VSUBS 1.67442f
C1557 VTAIL.n246 VSUBS 0.01599f
C1558 VTAIL.t10 VSUBS 0.080788f
C1559 VTAIL.n247 VSUBS 0.195101f
C1560 VTAIL.n248 VSUBS 0.024043f
C1561 VTAIL.n249 VSUBS 0.028346f
C1562 VTAIL.n250 VSUBS 0.037794f
C1563 VTAIL.n251 VSUBS 0.01693f
C1564 VTAIL.n252 VSUBS 0.01599f
C1565 VTAIL.n253 VSUBS 0.029756f
C1566 VTAIL.n254 VSUBS 0.029756f
C1567 VTAIL.n255 VSUBS 0.01599f
C1568 VTAIL.n256 VSUBS 0.01693f
C1569 VTAIL.n257 VSUBS 0.037794f
C1570 VTAIL.n258 VSUBS 0.037794f
C1571 VTAIL.n259 VSUBS 0.01693f
C1572 VTAIL.n260 VSUBS 0.01599f
C1573 VTAIL.n261 VSUBS 0.029756f
C1574 VTAIL.n262 VSUBS 0.029756f
C1575 VTAIL.n263 VSUBS 0.01599f
C1576 VTAIL.n264 VSUBS 0.01693f
C1577 VTAIL.n265 VSUBS 0.037794f
C1578 VTAIL.n266 VSUBS 0.037794f
C1579 VTAIL.n267 VSUBS 0.01693f
C1580 VTAIL.n268 VSUBS 0.01599f
C1581 VTAIL.n269 VSUBS 0.029756f
C1582 VTAIL.n270 VSUBS 0.029756f
C1583 VTAIL.n271 VSUBS 0.01599f
C1584 VTAIL.n272 VSUBS 0.01693f
C1585 VTAIL.n273 VSUBS 0.037794f
C1586 VTAIL.n274 VSUBS 0.037794f
C1587 VTAIL.n275 VSUBS 0.01693f
C1588 VTAIL.n276 VSUBS 0.01599f
C1589 VTAIL.n277 VSUBS 0.029756f
C1590 VTAIL.n278 VSUBS 0.029756f
C1591 VTAIL.n279 VSUBS 0.01599f
C1592 VTAIL.n280 VSUBS 0.01693f
C1593 VTAIL.n281 VSUBS 0.037794f
C1594 VTAIL.n282 VSUBS 0.037794f
C1595 VTAIL.n283 VSUBS 0.01693f
C1596 VTAIL.n284 VSUBS 0.01599f
C1597 VTAIL.n285 VSUBS 0.029756f
C1598 VTAIL.n286 VSUBS 0.029756f
C1599 VTAIL.n287 VSUBS 0.01599f
C1600 VTAIL.n288 VSUBS 0.01693f
C1601 VTAIL.n289 VSUBS 0.037794f
C1602 VTAIL.n290 VSUBS 0.093264f
C1603 VTAIL.n291 VSUBS 0.01693f
C1604 VTAIL.n292 VSUBS 0.0314f
C1605 VTAIL.n293 VSUBS 0.074065f
C1606 VTAIL.n294 VSUBS 0.071108f
C1607 VTAIL.n295 VSUBS 2.15518f
C1608 VN.n0 VSUBS 0.043939f
C1609 VN.t4 VSUBS 3.40324f
C1610 VN.n1 VSUBS 0.043536f
C1611 VN.n2 VSUBS 0.023359f
C1612 VN.n3 VSUBS 0.043536f
C1613 VN.t5 VSUBS 3.8046f
C1614 VN.n4 VSUBS 1.21552f
C1615 VN.t1 VSUBS 3.40324f
C1616 VN.n5 VSUBS 1.28276f
C1617 VN.n6 VSUBS 0.043536f
C1618 VN.n7 VSUBS 0.310699f
C1619 VN.n8 VSUBS 0.023359f
C1620 VN.n9 VSUBS 0.023359f
C1621 VN.n10 VSUBS 0.043536f
C1622 VN.n11 VSUBS 0.02857f
C1623 VN.n12 VSUBS 0.039635f
C1624 VN.n13 VSUBS 0.023359f
C1625 VN.n14 VSUBS 0.023359f
C1626 VN.n15 VSUBS 0.023359f
C1627 VN.n16 VSUBS 0.043536f
C1628 VN.n17 VSUBS 0.036228f
C1629 VN.n18 VSUBS 1.28167f
C1630 VN.n19 VSUBS 0.079585f
C1631 VN.n20 VSUBS 0.043939f
C1632 VN.t0 VSUBS 3.40324f
C1633 VN.n21 VSUBS 0.043536f
C1634 VN.n22 VSUBS 0.023359f
C1635 VN.n23 VSUBS 0.043536f
C1636 VN.t2 VSUBS 3.8046f
C1637 VN.n24 VSUBS 1.21552f
C1638 VN.t3 VSUBS 3.40324f
C1639 VN.n25 VSUBS 1.28276f
C1640 VN.n26 VSUBS 0.043536f
C1641 VN.n27 VSUBS 0.310699f
C1642 VN.n28 VSUBS 0.023359f
C1643 VN.n29 VSUBS 0.023359f
C1644 VN.n30 VSUBS 0.043536f
C1645 VN.n31 VSUBS 0.02857f
C1646 VN.n32 VSUBS 0.039635f
C1647 VN.n33 VSUBS 0.023359f
C1648 VN.n34 VSUBS 0.023359f
C1649 VN.n35 VSUBS 0.023359f
C1650 VN.n36 VSUBS 0.043536f
C1651 VN.n37 VSUBS 0.036228f
C1652 VN.n38 VSUBS 1.28167f
C1653 VN.n39 VSUBS 1.57372f
.ends

