* NGSPICE file created from diff_pair_sample_1693.ext - technology: sky130A

.subckt diff_pair_sample_1693 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=3.23235 ps=19.92 w=19.59 l=3.18
X1 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=3.23235 ps=19.92 w=19.59 l=3.18
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=0 ps=0 w=19.59 l=3.18
X3 VDD1.t4 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=3.23235 ps=19.92 w=19.59 l=3.18
X4 VDD1.t3 VP.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=7.6401 ps=39.96 w=19.59 l=3.18
X5 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=7.6401 ps=39.96 w=19.59 l=3.18
X6 VTAIL.t9 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=3.23235 ps=19.92 w=19.59 l=3.18
X7 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=3.23235 ps=19.92 w=19.59 l=3.18
X8 VTAIL.t8 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=3.23235 ps=19.92 w=19.59 l=3.18
X9 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=7.6401 ps=39.96 w=19.59 l=3.18
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=0 ps=0 w=19.59 l=3.18
X11 VTAIL.t0 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=3.23235 ps=19.92 w=19.59 l=3.18
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=0 ps=0 w=19.59 l=3.18
X13 VDD1.t0 VP.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=7.6401 ps=39.96 w=19.59 l=3.18
X14 VTAIL.t5 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.23235 pd=19.92 as=3.23235 ps=19.92 w=19.59 l=3.18
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6401 pd=39.96 as=0 ps=0 w=19.59 l=3.18
R0 VP.n14 VP.t0 181.172
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n12 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n11 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n10 161.3
R7 VP.n25 VP.n24 161.3
R8 VP.n49 VP.n48 161.3
R9 VP.n47 VP.n1 161.3
R10 VP.n46 VP.n45 161.3
R11 VP.n44 VP.n2 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n41 VP.n3 161.3
R14 VP.n40 VP.n39 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n8 VP.t1 148.465
R23 VP.n4 VP.t4 148.465
R24 VP.n0 VP.t5 148.465
R25 VP.n9 VP.t2 148.465
R26 VP.n13 VP.t3 148.465
R27 VP.n27 VP.n8 77.3446
R28 VP.n50 VP.n0 77.3446
R29 VP.n26 VP.n9 77.3446
R30 VP.n14 VP.n13 62.0352
R31 VP.n27 VP.n26 56.7531
R32 VP.n31 VP.n6 40.979
R33 VP.n46 VP.n2 40.979
R34 VP.n22 VP.n11 40.979
R35 VP.n35 VP.n6 40.0078
R36 VP.n42 VP.n2 40.0078
R37 VP.n18 VP.n11 40.0078
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 12.7233
R51 VP.n48 VP.n0 12.7233
R52 VP.n24 VP.n9 12.7233
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 4.25366
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n442 VTAIL.n338 289.615
R81 VTAIL.n106 VTAIL.n2 289.615
R82 VTAIL.n332 VTAIL.n228 289.615
R83 VTAIL.n220 VTAIL.n116 289.615
R84 VTAIL.n375 VTAIL.n374 185
R85 VTAIL.n377 VTAIL.n376 185
R86 VTAIL.n370 VTAIL.n369 185
R87 VTAIL.n383 VTAIL.n382 185
R88 VTAIL.n385 VTAIL.n384 185
R89 VTAIL.n366 VTAIL.n365 185
R90 VTAIL.n391 VTAIL.n390 185
R91 VTAIL.n393 VTAIL.n392 185
R92 VTAIL.n362 VTAIL.n361 185
R93 VTAIL.n399 VTAIL.n398 185
R94 VTAIL.n401 VTAIL.n400 185
R95 VTAIL.n358 VTAIL.n357 185
R96 VTAIL.n407 VTAIL.n406 185
R97 VTAIL.n409 VTAIL.n408 185
R98 VTAIL.n354 VTAIL.n353 185
R99 VTAIL.n416 VTAIL.n415 185
R100 VTAIL.n417 VTAIL.n352 185
R101 VTAIL.n419 VTAIL.n418 185
R102 VTAIL.n350 VTAIL.n349 185
R103 VTAIL.n425 VTAIL.n424 185
R104 VTAIL.n427 VTAIL.n426 185
R105 VTAIL.n346 VTAIL.n345 185
R106 VTAIL.n433 VTAIL.n432 185
R107 VTAIL.n435 VTAIL.n434 185
R108 VTAIL.n342 VTAIL.n341 185
R109 VTAIL.n441 VTAIL.n440 185
R110 VTAIL.n443 VTAIL.n442 185
R111 VTAIL.n39 VTAIL.n38 185
R112 VTAIL.n41 VTAIL.n40 185
R113 VTAIL.n34 VTAIL.n33 185
R114 VTAIL.n47 VTAIL.n46 185
R115 VTAIL.n49 VTAIL.n48 185
R116 VTAIL.n30 VTAIL.n29 185
R117 VTAIL.n55 VTAIL.n54 185
R118 VTAIL.n57 VTAIL.n56 185
R119 VTAIL.n26 VTAIL.n25 185
R120 VTAIL.n63 VTAIL.n62 185
R121 VTAIL.n65 VTAIL.n64 185
R122 VTAIL.n22 VTAIL.n21 185
R123 VTAIL.n71 VTAIL.n70 185
R124 VTAIL.n73 VTAIL.n72 185
R125 VTAIL.n18 VTAIL.n17 185
R126 VTAIL.n80 VTAIL.n79 185
R127 VTAIL.n81 VTAIL.n16 185
R128 VTAIL.n83 VTAIL.n82 185
R129 VTAIL.n14 VTAIL.n13 185
R130 VTAIL.n89 VTAIL.n88 185
R131 VTAIL.n91 VTAIL.n90 185
R132 VTAIL.n10 VTAIL.n9 185
R133 VTAIL.n97 VTAIL.n96 185
R134 VTAIL.n99 VTAIL.n98 185
R135 VTAIL.n6 VTAIL.n5 185
R136 VTAIL.n105 VTAIL.n104 185
R137 VTAIL.n107 VTAIL.n106 185
R138 VTAIL.n333 VTAIL.n332 185
R139 VTAIL.n331 VTAIL.n330 185
R140 VTAIL.n232 VTAIL.n231 185
R141 VTAIL.n325 VTAIL.n324 185
R142 VTAIL.n323 VTAIL.n322 185
R143 VTAIL.n236 VTAIL.n235 185
R144 VTAIL.n317 VTAIL.n316 185
R145 VTAIL.n315 VTAIL.n314 185
R146 VTAIL.n240 VTAIL.n239 185
R147 VTAIL.n244 VTAIL.n242 185
R148 VTAIL.n309 VTAIL.n308 185
R149 VTAIL.n307 VTAIL.n306 185
R150 VTAIL.n246 VTAIL.n245 185
R151 VTAIL.n301 VTAIL.n300 185
R152 VTAIL.n299 VTAIL.n298 185
R153 VTAIL.n250 VTAIL.n249 185
R154 VTAIL.n293 VTAIL.n292 185
R155 VTAIL.n291 VTAIL.n290 185
R156 VTAIL.n254 VTAIL.n253 185
R157 VTAIL.n285 VTAIL.n284 185
R158 VTAIL.n283 VTAIL.n282 185
R159 VTAIL.n258 VTAIL.n257 185
R160 VTAIL.n277 VTAIL.n276 185
R161 VTAIL.n275 VTAIL.n274 185
R162 VTAIL.n262 VTAIL.n261 185
R163 VTAIL.n269 VTAIL.n268 185
R164 VTAIL.n267 VTAIL.n266 185
R165 VTAIL.n221 VTAIL.n220 185
R166 VTAIL.n219 VTAIL.n218 185
R167 VTAIL.n120 VTAIL.n119 185
R168 VTAIL.n213 VTAIL.n212 185
R169 VTAIL.n211 VTAIL.n210 185
R170 VTAIL.n124 VTAIL.n123 185
R171 VTAIL.n205 VTAIL.n204 185
R172 VTAIL.n203 VTAIL.n202 185
R173 VTAIL.n128 VTAIL.n127 185
R174 VTAIL.n132 VTAIL.n130 185
R175 VTAIL.n197 VTAIL.n196 185
R176 VTAIL.n195 VTAIL.n194 185
R177 VTAIL.n134 VTAIL.n133 185
R178 VTAIL.n189 VTAIL.n188 185
R179 VTAIL.n187 VTAIL.n186 185
R180 VTAIL.n138 VTAIL.n137 185
R181 VTAIL.n181 VTAIL.n180 185
R182 VTAIL.n179 VTAIL.n178 185
R183 VTAIL.n142 VTAIL.n141 185
R184 VTAIL.n173 VTAIL.n172 185
R185 VTAIL.n171 VTAIL.n170 185
R186 VTAIL.n146 VTAIL.n145 185
R187 VTAIL.n165 VTAIL.n164 185
R188 VTAIL.n163 VTAIL.n162 185
R189 VTAIL.n150 VTAIL.n149 185
R190 VTAIL.n157 VTAIL.n156 185
R191 VTAIL.n155 VTAIL.n154 185
R192 VTAIL.n373 VTAIL.t3 147.659
R193 VTAIL.n37 VTAIL.t10 147.659
R194 VTAIL.n265 VTAIL.t11 147.659
R195 VTAIL.n153 VTAIL.t2 147.659
R196 VTAIL.n376 VTAIL.n375 104.615
R197 VTAIL.n376 VTAIL.n369 104.615
R198 VTAIL.n383 VTAIL.n369 104.615
R199 VTAIL.n384 VTAIL.n383 104.615
R200 VTAIL.n384 VTAIL.n365 104.615
R201 VTAIL.n391 VTAIL.n365 104.615
R202 VTAIL.n392 VTAIL.n391 104.615
R203 VTAIL.n392 VTAIL.n361 104.615
R204 VTAIL.n399 VTAIL.n361 104.615
R205 VTAIL.n400 VTAIL.n399 104.615
R206 VTAIL.n400 VTAIL.n357 104.615
R207 VTAIL.n407 VTAIL.n357 104.615
R208 VTAIL.n408 VTAIL.n407 104.615
R209 VTAIL.n408 VTAIL.n353 104.615
R210 VTAIL.n416 VTAIL.n353 104.615
R211 VTAIL.n417 VTAIL.n416 104.615
R212 VTAIL.n418 VTAIL.n417 104.615
R213 VTAIL.n418 VTAIL.n349 104.615
R214 VTAIL.n425 VTAIL.n349 104.615
R215 VTAIL.n426 VTAIL.n425 104.615
R216 VTAIL.n426 VTAIL.n345 104.615
R217 VTAIL.n433 VTAIL.n345 104.615
R218 VTAIL.n434 VTAIL.n433 104.615
R219 VTAIL.n434 VTAIL.n341 104.615
R220 VTAIL.n441 VTAIL.n341 104.615
R221 VTAIL.n442 VTAIL.n441 104.615
R222 VTAIL.n40 VTAIL.n39 104.615
R223 VTAIL.n40 VTAIL.n33 104.615
R224 VTAIL.n47 VTAIL.n33 104.615
R225 VTAIL.n48 VTAIL.n47 104.615
R226 VTAIL.n48 VTAIL.n29 104.615
R227 VTAIL.n55 VTAIL.n29 104.615
R228 VTAIL.n56 VTAIL.n55 104.615
R229 VTAIL.n56 VTAIL.n25 104.615
R230 VTAIL.n63 VTAIL.n25 104.615
R231 VTAIL.n64 VTAIL.n63 104.615
R232 VTAIL.n64 VTAIL.n21 104.615
R233 VTAIL.n71 VTAIL.n21 104.615
R234 VTAIL.n72 VTAIL.n71 104.615
R235 VTAIL.n72 VTAIL.n17 104.615
R236 VTAIL.n80 VTAIL.n17 104.615
R237 VTAIL.n81 VTAIL.n80 104.615
R238 VTAIL.n82 VTAIL.n81 104.615
R239 VTAIL.n82 VTAIL.n13 104.615
R240 VTAIL.n89 VTAIL.n13 104.615
R241 VTAIL.n90 VTAIL.n89 104.615
R242 VTAIL.n90 VTAIL.n9 104.615
R243 VTAIL.n97 VTAIL.n9 104.615
R244 VTAIL.n98 VTAIL.n97 104.615
R245 VTAIL.n98 VTAIL.n5 104.615
R246 VTAIL.n105 VTAIL.n5 104.615
R247 VTAIL.n106 VTAIL.n105 104.615
R248 VTAIL.n332 VTAIL.n331 104.615
R249 VTAIL.n331 VTAIL.n231 104.615
R250 VTAIL.n324 VTAIL.n231 104.615
R251 VTAIL.n324 VTAIL.n323 104.615
R252 VTAIL.n323 VTAIL.n235 104.615
R253 VTAIL.n316 VTAIL.n235 104.615
R254 VTAIL.n316 VTAIL.n315 104.615
R255 VTAIL.n315 VTAIL.n239 104.615
R256 VTAIL.n244 VTAIL.n239 104.615
R257 VTAIL.n308 VTAIL.n244 104.615
R258 VTAIL.n308 VTAIL.n307 104.615
R259 VTAIL.n307 VTAIL.n245 104.615
R260 VTAIL.n300 VTAIL.n245 104.615
R261 VTAIL.n300 VTAIL.n299 104.615
R262 VTAIL.n299 VTAIL.n249 104.615
R263 VTAIL.n292 VTAIL.n249 104.615
R264 VTAIL.n292 VTAIL.n291 104.615
R265 VTAIL.n291 VTAIL.n253 104.615
R266 VTAIL.n284 VTAIL.n253 104.615
R267 VTAIL.n284 VTAIL.n283 104.615
R268 VTAIL.n283 VTAIL.n257 104.615
R269 VTAIL.n276 VTAIL.n257 104.615
R270 VTAIL.n276 VTAIL.n275 104.615
R271 VTAIL.n275 VTAIL.n261 104.615
R272 VTAIL.n268 VTAIL.n261 104.615
R273 VTAIL.n268 VTAIL.n267 104.615
R274 VTAIL.n220 VTAIL.n219 104.615
R275 VTAIL.n219 VTAIL.n119 104.615
R276 VTAIL.n212 VTAIL.n119 104.615
R277 VTAIL.n212 VTAIL.n211 104.615
R278 VTAIL.n211 VTAIL.n123 104.615
R279 VTAIL.n204 VTAIL.n123 104.615
R280 VTAIL.n204 VTAIL.n203 104.615
R281 VTAIL.n203 VTAIL.n127 104.615
R282 VTAIL.n132 VTAIL.n127 104.615
R283 VTAIL.n196 VTAIL.n132 104.615
R284 VTAIL.n196 VTAIL.n195 104.615
R285 VTAIL.n195 VTAIL.n133 104.615
R286 VTAIL.n188 VTAIL.n133 104.615
R287 VTAIL.n188 VTAIL.n187 104.615
R288 VTAIL.n187 VTAIL.n137 104.615
R289 VTAIL.n180 VTAIL.n137 104.615
R290 VTAIL.n180 VTAIL.n179 104.615
R291 VTAIL.n179 VTAIL.n141 104.615
R292 VTAIL.n172 VTAIL.n141 104.615
R293 VTAIL.n172 VTAIL.n171 104.615
R294 VTAIL.n171 VTAIL.n145 104.615
R295 VTAIL.n164 VTAIL.n145 104.615
R296 VTAIL.n164 VTAIL.n163 104.615
R297 VTAIL.n163 VTAIL.n149 104.615
R298 VTAIL.n156 VTAIL.n149 104.615
R299 VTAIL.n156 VTAIL.n155 104.615
R300 VTAIL.n375 VTAIL.t3 52.3082
R301 VTAIL.n39 VTAIL.t10 52.3082
R302 VTAIL.n267 VTAIL.t11 52.3082
R303 VTAIL.n155 VTAIL.t2 52.3082
R304 VTAIL.n227 VTAIL.n226 42.1779
R305 VTAIL.n115 VTAIL.n114 42.1779
R306 VTAIL.n1 VTAIL.n0 42.1777
R307 VTAIL.n113 VTAIL.n112 42.1777
R308 VTAIL.n115 VTAIL.n113 35.3065
R309 VTAIL.n447 VTAIL.n337 32.2807
R310 VTAIL.n447 VTAIL.n446 30.4399
R311 VTAIL.n111 VTAIL.n110 30.4399
R312 VTAIL.n337 VTAIL.n336 30.4399
R313 VTAIL.n225 VTAIL.n224 30.4399
R314 VTAIL.n374 VTAIL.n373 15.6677
R315 VTAIL.n38 VTAIL.n37 15.6677
R316 VTAIL.n266 VTAIL.n265 15.6677
R317 VTAIL.n154 VTAIL.n153 15.6677
R318 VTAIL.n419 VTAIL.n350 13.1884
R319 VTAIL.n83 VTAIL.n14 13.1884
R320 VTAIL.n242 VTAIL.n240 13.1884
R321 VTAIL.n130 VTAIL.n128 13.1884
R322 VTAIL.n377 VTAIL.n372 12.8005
R323 VTAIL.n420 VTAIL.n352 12.8005
R324 VTAIL.n424 VTAIL.n423 12.8005
R325 VTAIL.n41 VTAIL.n36 12.8005
R326 VTAIL.n84 VTAIL.n16 12.8005
R327 VTAIL.n88 VTAIL.n87 12.8005
R328 VTAIL.n314 VTAIL.n313 12.8005
R329 VTAIL.n310 VTAIL.n309 12.8005
R330 VTAIL.n269 VTAIL.n264 12.8005
R331 VTAIL.n202 VTAIL.n201 12.8005
R332 VTAIL.n198 VTAIL.n197 12.8005
R333 VTAIL.n157 VTAIL.n152 12.8005
R334 VTAIL.n378 VTAIL.n370 12.0247
R335 VTAIL.n415 VTAIL.n414 12.0247
R336 VTAIL.n427 VTAIL.n348 12.0247
R337 VTAIL.n42 VTAIL.n34 12.0247
R338 VTAIL.n79 VTAIL.n78 12.0247
R339 VTAIL.n91 VTAIL.n12 12.0247
R340 VTAIL.n317 VTAIL.n238 12.0247
R341 VTAIL.n306 VTAIL.n243 12.0247
R342 VTAIL.n270 VTAIL.n262 12.0247
R343 VTAIL.n205 VTAIL.n126 12.0247
R344 VTAIL.n194 VTAIL.n131 12.0247
R345 VTAIL.n158 VTAIL.n150 12.0247
R346 VTAIL.n382 VTAIL.n381 11.249
R347 VTAIL.n413 VTAIL.n354 11.249
R348 VTAIL.n428 VTAIL.n346 11.249
R349 VTAIL.n46 VTAIL.n45 11.249
R350 VTAIL.n77 VTAIL.n18 11.249
R351 VTAIL.n92 VTAIL.n10 11.249
R352 VTAIL.n318 VTAIL.n236 11.249
R353 VTAIL.n305 VTAIL.n246 11.249
R354 VTAIL.n274 VTAIL.n273 11.249
R355 VTAIL.n206 VTAIL.n124 11.249
R356 VTAIL.n193 VTAIL.n134 11.249
R357 VTAIL.n162 VTAIL.n161 11.249
R358 VTAIL.n385 VTAIL.n368 10.4732
R359 VTAIL.n410 VTAIL.n409 10.4732
R360 VTAIL.n432 VTAIL.n431 10.4732
R361 VTAIL.n49 VTAIL.n32 10.4732
R362 VTAIL.n74 VTAIL.n73 10.4732
R363 VTAIL.n96 VTAIL.n95 10.4732
R364 VTAIL.n322 VTAIL.n321 10.4732
R365 VTAIL.n302 VTAIL.n301 10.4732
R366 VTAIL.n277 VTAIL.n260 10.4732
R367 VTAIL.n210 VTAIL.n209 10.4732
R368 VTAIL.n190 VTAIL.n189 10.4732
R369 VTAIL.n165 VTAIL.n148 10.4732
R370 VTAIL.n386 VTAIL.n366 9.69747
R371 VTAIL.n406 VTAIL.n356 9.69747
R372 VTAIL.n435 VTAIL.n344 9.69747
R373 VTAIL.n50 VTAIL.n30 9.69747
R374 VTAIL.n70 VTAIL.n20 9.69747
R375 VTAIL.n99 VTAIL.n8 9.69747
R376 VTAIL.n325 VTAIL.n234 9.69747
R377 VTAIL.n298 VTAIL.n248 9.69747
R378 VTAIL.n278 VTAIL.n258 9.69747
R379 VTAIL.n213 VTAIL.n122 9.69747
R380 VTAIL.n186 VTAIL.n136 9.69747
R381 VTAIL.n166 VTAIL.n146 9.69747
R382 VTAIL.n446 VTAIL.n445 9.45567
R383 VTAIL.n110 VTAIL.n109 9.45567
R384 VTAIL.n336 VTAIL.n335 9.45567
R385 VTAIL.n224 VTAIL.n223 9.45567
R386 VTAIL.n445 VTAIL.n444 9.3005
R387 VTAIL.n439 VTAIL.n438 9.3005
R388 VTAIL.n437 VTAIL.n436 9.3005
R389 VTAIL.n344 VTAIL.n343 9.3005
R390 VTAIL.n431 VTAIL.n430 9.3005
R391 VTAIL.n429 VTAIL.n428 9.3005
R392 VTAIL.n348 VTAIL.n347 9.3005
R393 VTAIL.n423 VTAIL.n422 9.3005
R394 VTAIL.n395 VTAIL.n394 9.3005
R395 VTAIL.n364 VTAIL.n363 9.3005
R396 VTAIL.n389 VTAIL.n388 9.3005
R397 VTAIL.n387 VTAIL.n386 9.3005
R398 VTAIL.n368 VTAIL.n367 9.3005
R399 VTAIL.n381 VTAIL.n380 9.3005
R400 VTAIL.n379 VTAIL.n378 9.3005
R401 VTAIL.n372 VTAIL.n371 9.3005
R402 VTAIL.n397 VTAIL.n396 9.3005
R403 VTAIL.n360 VTAIL.n359 9.3005
R404 VTAIL.n403 VTAIL.n402 9.3005
R405 VTAIL.n405 VTAIL.n404 9.3005
R406 VTAIL.n356 VTAIL.n355 9.3005
R407 VTAIL.n411 VTAIL.n410 9.3005
R408 VTAIL.n413 VTAIL.n412 9.3005
R409 VTAIL.n414 VTAIL.n351 9.3005
R410 VTAIL.n421 VTAIL.n420 9.3005
R411 VTAIL.n340 VTAIL.n339 9.3005
R412 VTAIL.n109 VTAIL.n108 9.3005
R413 VTAIL.n103 VTAIL.n102 9.3005
R414 VTAIL.n101 VTAIL.n100 9.3005
R415 VTAIL.n8 VTAIL.n7 9.3005
R416 VTAIL.n95 VTAIL.n94 9.3005
R417 VTAIL.n93 VTAIL.n92 9.3005
R418 VTAIL.n12 VTAIL.n11 9.3005
R419 VTAIL.n87 VTAIL.n86 9.3005
R420 VTAIL.n59 VTAIL.n58 9.3005
R421 VTAIL.n28 VTAIL.n27 9.3005
R422 VTAIL.n53 VTAIL.n52 9.3005
R423 VTAIL.n51 VTAIL.n50 9.3005
R424 VTAIL.n32 VTAIL.n31 9.3005
R425 VTAIL.n45 VTAIL.n44 9.3005
R426 VTAIL.n43 VTAIL.n42 9.3005
R427 VTAIL.n36 VTAIL.n35 9.3005
R428 VTAIL.n61 VTAIL.n60 9.3005
R429 VTAIL.n24 VTAIL.n23 9.3005
R430 VTAIL.n67 VTAIL.n66 9.3005
R431 VTAIL.n69 VTAIL.n68 9.3005
R432 VTAIL.n20 VTAIL.n19 9.3005
R433 VTAIL.n75 VTAIL.n74 9.3005
R434 VTAIL.n77 VTAIL.n76 9.3005
R435 VTAIL.n78 VTAIL.n15 9.3005
R436 VTAIL.n85 VTAIL.n84 9.3005
R437 VTAIL.n4 VTAIL.n3 9.3005
R438 VTAIL.n252 VTAIL.n251 9.3005
R439 VTAIL.n295 VTAIL.n294 9.3005
R440 VTAIL.n297 VTAIL.n296 9.3005
R441 VTAIL.n248 VTAIL.n247 9.3005
R442 VTAIL.n303 VTAIL.n302 9.3005
R443 VTAIL.n305 VTAIL.n304 9.3005
R444 VTAIL.n243 VTAIL.n241 9.3005
R445 VTAIL.n311 VTAIL.n310 9.3005
R446 VTAIL.n335 VTAIL.n334 9.3005
R447 VTAIL.n230 VTAIL.n229 9.3005
R448 VTAIL.n329 VTAIL.n328 9.3005
R449 VTAIL.n327 VTAIL.n326 9.3005
R450 VTAIL.n234 VTAIL.n233 9.3005
R451 VTAIL.n321 VTAIL.n320 9.3005
R452 VTAIL.n319 VTAIL.n318 9.3005
R453 VTAIL.n238 VTAIL.n237 9.3005
R454 VTAIL.n313 VTAIL.n312 9.3005
R455 VTAIL.n289 VTAIL.n288 9.3005
R456 VTAIL.n287 VTAIL.n286 9.3005
R457 VTAIL.n256 VTAIL.n255 9.3005
R458 VTAIL.n281 VTAIL.n280 9.3005
R459 VTAIL.n279 VTAIL.n278 9.3005
R460 VTAIL.n260 VTAIL.n259 9.3005
R461 VTAIL.n273 VTAIL.n272 9.3005
R462 VTAIL.n271 VTAIL.n270 9.3005
R463 VTAIL.n264 VTAIL.n263 9.3005
R464 VTAIL.n140 VTAIL.n139 9.3005
R465 VTAIL.n183 VTAIL.n182 9.3005
R466 VTAIL.n185 VTAIL.n184 9.3005
R467 VTAIL.n136 VTAIL.n135 9.3005
R468 VTAIL.n191 VTAIL.n190 9.3005
R469 VTAIL.n193 VTAIL.n192 9.3005
R470 VTAIL.n131 VTAIL.n129 9.3005
R471 VTAIL.n199 VTAIL.n198 9.3005
R472 VTAIL.n223 VTAIL.n222 9.3005
R473 VTAIL.n118 VTAIL.n117 9.3005
R474 VTAIL.n217 VTAIL.n216 9.3005
R475 VTAIL.n215 VTAIL.n214 9.3005
R476 VTAIL.n122 VTAIL.n121 9.3005
R477 VTAIL.n209 VTAIL.n208 9.3005
R478 VTAIL.n207 VTAIL.n206 9.3005
R479 VTAIL.n126 VTAIL.n125 9.3005
R480 VTAIL.n201 VTAIL.n200 9.3005
R481 VTAIL.n177 VTAIL.n176 9.3005
R482 VTAIL.n175 VTAIL.n174 9.3005
R483 VTAIL.n144 VTAIL.n143 9.3005
R484 VTAIL.n169 VTAIL.n168 9.3005
R485 VTAIL.n167 VTAIL.n166 9.3005
R486 VTAIL.n148 VTAIL.n147 9.3005
R487 VTAIL.n161 VTAIL.n160 9.3005
R488 VTAIL.n159 VTAIL.n158 9.3005
R489 VTAIL.n152 VTAIL.n151 9.3005
R490 VTAIL.n390 VTAIL.n389 8.92171
R491 VTAIL.n405 VTAIL.n358 8.92171
R492 VTAIL.n436 VTAIL.n342 8.92171
R493 VTAIL.n54 VTAIL.n53 8.92171
R494 VTAIL.n69 VTAIL.n22 8.92171
R495 VTAIL.n100 VTAIL.n6 8.92171
R496 VTAIL.n326 VTAIL.n232 8.92171
R497 VTAIL.n297 VTAIL.n250 8.92171
R498 VTAIL.n282 VTAIL.n281 8.92171
R499 VTAIL.n214 VTAIL.n120 8.92171
R500 VTAIL.n185 VTAIL.n138 8.92171
R501 VTAIL.n170 VTAIL.n169 8.92171
R502 VTAIL.n393 VTAIL.n364 8.14595
R503 VTAIL.n402 VTAIL.n401 8.14595
R504 VTAIL.n440 VTAIL.n439 8.14595
R505 VTAIL.n57 VTAIL.n28 8.14595
R506 VTAIL.n66 VTAIL.n65 8.14595
R507 VTAIL.n104 VTAIL.n103 8.14595
R508 VTAIL.n330 VTAIL.n329 8.14595
R509 VTAIL.n294 VTAIL.n293 8.14595
R510 VTAIL.n285 VTAIL.n256 8.14595
R511 VTAIL.n218 VTAIL.n217 8.14595
R512 VTAIL.n182 VTAIL.n181 8.14595
R513 VTAIL.n173 VTAIL.n144 8.14595
R514 VTAIL.n394 VTAIL.n362 7.3702
R515 VTAIL.n398 VTAIL.n360 7.3702
R516 VTAIL.n443 VTAIL.n340 7.3702
R517 VTAIL.n446 VTAIL.n338 7.3702
R518 VTAIL.n58 VTAIL.n26 7.3702
R519 VTAIL.n62 VTAIL.n24 7.3702
R520 VTAIL.n107 VTAIL.n4 7.3702
R521 VTAIL.n110 VTAIL.n2 7.3702
R522 VTAIL.n336 VTAIL.n228 7.3702
R523 VTAIL.n333 VTAIL.n230 7.3702
R524 VTAIL.n290 VTAIL.n252 7.3702
R525 VTAIL.n286 VTAIL.n254 7.3702
R526 VTAIL.n224 VTAIL.n116 7.3702
R527 VTAIL.n221 VTAIL.n118 7.3702
R528 VTAIL.n178 VTAIL.n140 7.3702
R529 VTAIL.n174 VTAIL.n142 7.3702
R530 VTAIL.n397 VTAIL.n362 6.59444
R531 VTAIL.n398 VTAIL.n397 6.59444
R532 VTAIL.n444 VTAIL.n443 6.59444
R533 VTAIL.n444 VTAIL.n338 6.59444
R534 VTAIL.n61 VTAIL.n26 6.59444
R535 VTAIL.n62 VTAIL.n61 6.59444
R536 VTAIL.n108 VTAIL.n107 6.59444
R537 VTAIL.n108 VTAIL.n2 6.59444
R538 VTAIL.n334 VTAIL.n228 6.59444
R539 VTAIL.n334 VTAIL.n333 6.59444
R540 VTAIL.n290 VTAIL.n289 6.59444
R541 VTAIL.n289 VTAIL.n254 6.59444
R542 VTAIL.n222 VTAIL.n116 6.59444
R543 VTAIL.n222 VTAIL.n221 6.59444
R544 VTAIL.n178 VTAIL.n177 6.59444
R545 VTAIL.n177 VTAIL.n142 6.59444
R546 VTAIL.n394 VTAIL.n393 5.81868
R547 VTAIL.n401 VTAIL.n360 5.81868
R548 VTAIL.n440 VTAIL.n340 5.81868
R549 VTAIL.n58 VTAIL.n57 5.81868
R550 VTAIL.n65 VTAIL.n24 5.81868
R551 VTAIL.n104 VTAIL.n4 5.81868
R552 VTAIL.n330 VTAIL.n230 5.81868
R553 VTAIL.n293 VTAIL.n252 5.81868
R554 VTAIL.n286 VTAIL.n285 5.81868
R555 VTAIL.n218 VTAIL.n118 5.81868
R556 VTAIL.n181 VTAIL.n140 5.81868
R557 VTAIL.n174 VTAIL.n173 5.81868
R558 VTAIL.n390 VTAIL.n364 5.04292
R559 VTAIL.n402 VTAIL.n358 5.04292
R560 VTAIL.n439 VTAIL.n342 5.04292
R561 VTAIL.n54 VTAIL.n28 5.04292
R562 VTAIL.n66 VTAIL.n22 5.04292
R563 VTAIL.n103 VTAIL.n6 5.04292
R564 VTAIL.n329 VTAIL.n232 5.04292
R565 VTAIL.n294 VTAIL.n250 5.04292
R566 VTAIL.n282 VTAIL.n256 5.04292
R567 VTAIL.n217 VTAIL.n120 5.04292
R568 VTAIL.n182 VTAIL.n138 5.04292
R569 VTAIL.n170 VTAIL.n144 5.04292
R570 VTAIL.n373 VTAIL.n371 4.38563
R571 VTAIL.n37 VTAIL.n35 4.38563
R572 VTAIL.n265 VTAIL.n263 4.38563
R573 VTAIL.n153 VTAIL.n151 4.38563
R574 VTAIL.n389 VTAIL.n366 4.26717
R575 VTAIL.n406 VTAIL.n405 4.26717
R576 VTAIL.n436 VTAIL.n435 4.26717
R577 VTAIL.n53 VTAIL.n30 4.26717
R578 VTAIL.n70 VTAIL.n69 4.26717
R579 VTAIL.n100 VTAIL.n99 4.26717
R580 VTAIL.n326 VTAIL.n325 4.26717
R581 VTAIL.n298 VTAIL.n297 4.26717
R582 VTAIL.n281 VTAIL.n258 4.26717
R583 VTAIL.n214 VTAIL.n213 4.26717
R584 VTAIL.n186 VTAIL.n185 4.26717
R585 VTAIL.n169 VTAIL.n146 4.26717
R586 VTAIL.n386 VTAIL.n385 3.49141
R587 VTAIL.n409 VTAIL.n356 3.49141
R588 VTAIL.n432 VTAIL.n344 3.49141
R589 VTAIL.n50 VTAIL.n49 3.49141
R590 VTAIL.n73 VTAIL.n20 3.49141
R591 VTAIL.n96 VTAIL.n8 3.49141
R592 VTAIL.n322 VTAIL.n234 3.49141
R593 VTAIL.n301 VTAIL.n248 3.49141
R594 VTAIL.n278 VTAIL.n277 3.49141
R595 VTAIL.n210 VTAIL.n122 3.49141
R596 VTAIL.n189 VTAIL.n136 3.49141
R597 VTAIL.n166 VTAIL.n165 3.49141
R598 VTAIL.n225 VTAIL.n115 3.02636
R599 VTAIL.n337 VTAIL.n227 3.02636
R600 VTAIL.n113 VTAIL.n111 3.02636
R601 VTAIL.n382 VTAIL.n368 2.71565
R602 VTAIL.n410 VTAIL.n354 2.71565
R603 VTAIL.n431 VTAIL.n346 2.71565
R604 VTAIL.n46 VTAIL.n32 2.71565
R605 VTAIL.n74 VTAIL.n18 2.71565
R606 VTAIL.n95 VTAIL.n10 2.71565
R607 VTAIL.n321 VTAIL.n236 2.71565
R608 VTAIL.n302 VTAIL.n246 2.71565
R609 VTAIL.n274 VTAIL.n260 2.71565
R610 VTAIL.n209 VTAIL.n124 2.71565
R611 VTAIL.n190 VTAIL.n134 2.71565
R612 VTAIL.n162 VTAIL.n148 2.71565
R613 VTAIL VTAIL.n447 2.21171
R614 VTAIL.n227 VTAIL.n225 1.98326
R615 VTAIL.n111 VTAIL.n1 1.98326
R616 VTAIL.n381 VTAIL.n370 1.93989
R617 VTAIL.n415 VTAIL.n413 1.93989
R618 VTAIL.n428 VTAIL.n427 1.93989
R619 VTAIL.n45 VTAIL.n34 1.93989
R620 VTAIL.n79 VTAIL.n77 1.93989
R621 VTAIL.n92 VTAIL.n91 1.93989
R622 VTAIL.n318 VTAIL.n317 1.93989
R623 VTAIL.n306 VTAIL.n305 1.93989
R624 VTAIL.n273 VTAIL.n262 1.93989
R625 VTAIL.n206 VTAIL.n205 1.93989
R626 VTAIL.n194 VTAIL.n193 1.93989
R627 VTAIL.n161 VTAIL.n150 1.93989
R628 VTAIL.n378 VTAIL.n377 1.16414
R629 VTAIL.n414 VTAIL.n352 1.16414
R630 VTAIL.n424 VTAIL.n348 1.16414
R631 VTAIL.n42 VTAIL.n41 1.16414
R632 VTAIL.n78 VTAIL.n16 1.16414
R633 VTAIL.n88 VTAIL.n12 1.16414
R634 VTAIL.n314 VTAIL.n238 1.16414
R635 VTAIL.n309 VTAIL.n243 1.16414
R636 VTAIL.n270 VTAIL.n269 1.16414
R637 VTAIL.n202 VTAIL.n126 1.16414
R638 VTAIL.n197 VTAIL.n131 1.16414
R639 VTAIL.n158 VTAIL.n157 1.16414
R640 VTAIL.n0 VTAIL.t4 1.01122
R641 VTAIL.n0 VTAIL.t0 1.01122
R642 VTAIL.n112 VTAIL.t6 1.01122
R643 VTAIL.n112 VTAIL.t8 1.01122
R644 VTAIL.n226 VTAIL.t7 1.01122
R645 VTAIL.n226 VTAIL.t9 1.01122
R646 VTAIL.n114 VTAIL.t1 1.01122
R647 VTAIL.n114 VTAIL.t5 1.01122
R648 VTAIL VTAIL.n1 0.815155
R649 VTAIL.n374 VTAIL.n372 0.388379
R650 VTAIL.n420 VTAIL.n419 0.388379
R651 VTAIL.n423 VTAIL.n350 0.388379
R652 VTAIL.n38 VTAIL.n36 0.388379
R653 VTAIL.n84 VTAIL.n83 0.388379
R654 VTAIL.n87 VTAIL.n14 0.388379
R655 VTAIL.n313 VTAIL.n240 0.388379
R656 VTAIL.n310 VTAIL.n242 0.388379
R657 VTAIL.n266 VTAIL.n264 0.388379
R658 VTAIL.n201 VTAIL.n128 0.388379
R659 VTAIL.n198 VTAIL.n130 0.388379
R660 VTAIL.n154 VTAIL.n152 0.388379
R661 VTAIL.n379 VTAIL.n371 0.155672
R662 VTAIL.n380 VTAIL.n379 0.155672
R663 VTAIL.n380 VTAIL.n367 0.155672
R664 VTAIL.n387 VTAIL.n367 0.155672
R665 VTAIL.n388 VTAIL.n387 0.155672
R666 VTAIL.n388 VTAIL.n363 0.155672
R667 VTAIL.n395 VTAIL.n363 0.155672
R668 VTAIL.n396 VTAIL.n395 0.155672
R669 VTAIL.n396 VTAIL.n359 0.155672
R670 VTAIL.n403 VTAIL.n359 0.155672
R671 VTAIL.n404 VTAIL.n403 0.155672
R672 VTAIL.n404 VTAIL.n355 0.155672
R673 VTAIL.n411 VTAIL.n355 0.155672
R674 VTAIL.n412 VTAIL.n411 0.155672
R675 VTAIL.n412 VTAIL.n351 0.155672
R676 VTAIL.n421 VTAIL.n351 0.155672
R677 VTAIL.n422 VTAIL.n421 0.155672
R678 VTAIL.n422 VTAIL.n347 0.155672
R679 VTAIL.n429 VTAIL.n347 0.155672
R680 VTAIL.n430 VTAIL.n429 0.155672
R681 VTAIL.n430 VTAIL.n343 0.155672
R682 VTAIL.n437 VTAIL.n343 0.155672
R683 VTAIL.n438 VTAIL.n437 0.155672
R684 VTAIL.n438 VTAIL.n339 0.155672
R685 VTAIL.n445 VTAIL.n339 0.155672
R686 VTAIL.n43 VTAIL.n35 0.155672
R687 VTAIL.n44 VTAIL.n43 0.155672
R688 VTAIL.n44 VTAIL.n31 0.155672
R689 VTAIL.n51 VTAIL.n31 0.155672
R690 VTAIL.n52 VTAIL.n51 0.155672
R691 VTAIL.n52 VTAIL.n27 0.155672
R692 VTAIL.n59 VTAIL.n27 0.155672
R693 VTAIL.n60 VTAIL.n59 0.155672
R694 VTAIL.n60 VTAIL.n23 0.155672
R695 VTAIL.n67 VTAIL.n23 0.155672
R696 VTAIL.n68 VTAIL.n67 0.155672
R697 VTAIL.n68 VTAIL.n19 0.155672
R698 VTAIL.n75 VTAIL.n19 0.155672
R699 VTAIL.n76 VTAIL.n75 0.155672
R700 VTAIL.n76 VTAIL.n15 0.155672
R701 VTAIL.n85 VTAIL.n15 0.155672
R702 VTAIL.n86 VTAIL.n85 0.155672
R703 VTAIL.n86 VTAIL.n11 0.155672
R704 VTAIL.n93 VTAIL.n11 0.155672
R705 VTAIL.n94 VTAIL.n93 0.155672
R706 VTAIL.n94 VTAIL.n7 0.155672
R707 VTAIL.n101 VTAIL.n7 0.155672
R708 VTAIL.n102 VTAIL.n101 0.155672
R709 VTAIL.n102 VTAIL.n3 0.155672
R710 VTAIL.n109 VTAIL.n3 0.155672
R711 VTAIL.n335 VTAIL.n229 0.155672
R712 VTAIL.n328 VTAIL.n229 0.155672
R713 VTAIL.n328 VTAIL.n327 0.155672
R714 VTAIL.n327 VTAIL.n233 0.155672
R715 VTAIL.n320 VTAIL.n233 0.155672
R716 VTAIL.n320 VTAIL.n319 0.155672
R717 VTAIL.n319 VTAIL.n237 0.155672
R718 VTAIL.n312 VTAIL.n237 0.155672
R719 VTAIL.n312 VTAIL.n311 0.155672
R720 VTAIL.n311 VTAIL.n241 0.155672
R721 VTAIL.n304 VTAIL.n241 0.155672
R722 VTAIL.n304 VTAIL.n303 0.155672
R723 VTAIL.n303 VTAIL.n247 0.155672
R724 VTAIL.n296 VTAIL.n247 0.155672
R725 VTAIL.n296 VTAIL.n295 0.155672
R726 VTAIL.n295 VTAIL.n251 0.155672
R727 VTAIL.n288 VTAIL.n251 0.155672
R728 VTAIL.n288 VTAIL.n287 0.155672
R729 VTAIL.n287 VTAIL.n255 0.155672
R730 VTAIL.n280 VTAIL.n255 0.155672
R731 VTAIL.n280 VTAIL.n279 0.155672
R732 VTAIL.n279 VTAIL.n259 0.155672
R733 VTAIL.n272 VTAIL.n259 0.155672
R734 VTAIL.n272 VTAIL.n271 0.155672
R735 VTAIL.n271 VTAIL.n263 0.155672
R736 VTAIL.n223 VTAIL.n117 0.155672
R737 VTAIL.n216 VTAIL.n117 0.155672
R738 VTAIL.n216 VTAIL.n215 0.155672
R739 VTAIL.n215 VTAIL.n121 0.155672
R740 VTAIL.n208 VTAIL.n121 0.155672
R741 VTAIL.n208 VTAIL.n207 0.155672
R742 VTAIL.n207 VTAIL.n125 0.155672
R743 VTAIL.n200 VTAIL.n125 0.155672
R744 VTAIL.n200 VTAIL.n199 0.155672
R745 VTAIL.n199 VTAIL.n129 0.155672
R746 VTAIL.n192 VTAIL.n129 0.155672
R747 VTAIL.n192 VTAIL.n191 0.155672
R748 VTAIL.n191 VTAIL.n135 0.155672
R749 VTAIL.n184 VTAIL.n135 0.155672
R750 VTAIL.n184 VTAIL.n183 0.155672
R751 VTAIL.n183 VTAIL.n139 0.155672
R752 VTAIL.n176 VTAIL.n139 0.155672
R753 VTAIL.n176 VTAIL.n175 0.155672
R754 VTAIL.n175 VTAIL.n143 0.155672
R755 VTAIL.n168 VTAIL.n143 0.155672
R756 VTAIL.n168 VTAIL.n167 0.155672
R757 VTAIL.n167 VTAIL.n147 0.155672
R758 VTAIL.n160 VTAIL.n147 0.155672
R759 VTAIL.n160 VTAIL.n159 0.155672
R760 VTAIL.n159 VTAIL.n151 0.155672
R761 VDD1.n104 VDD1.n0 289.615
R762 VDD1.n213 VDD1.n109 289.615
R763 VDD1.n105 VDD1.n104 185
R764 VDD1.n103 VDD1.n102 185
R765 VDD1.n4 VDD1.n3 185
R766 VDD1.n97 VDD1.n96 185
R767 VDD1.n95 VDD1.n94 185
R768 VDD1.n8 VDD1.n7 185
R769 VDD1.n89 VDD1.n88 185
R770 VDD1.n87 VDD1.n86 185
R771 VDD1.n12 VDD1.n11 185
R772 VDD1.n16 VDD1.n14 185
R773 VDD1.n81 VDD1.n80 185
R774 VDD1.n79 VDD1.n78 185
R775 VDD1.n18 VDD1.n17 185
R776 VDD1.n73 VDD1.n72 185
R777 VDD1.n71 VDD1.n70 185
R778 VDD1.n22 VDD1.n21 185
R779 VDD1.n65 VDD1.n64 185
R780 VDD1.n63 VDD1.n62 185
R781 VDD1.n26 VDD1.n25 185
R782 VDD1.n57 VDD1.n56 185
R783 VDD1.n55 VDD1.n54 185
R784 VDD1.n30 VDD1.n29 185
R785 VDD1.n49 VDD1.n48 185
R786 VDD1.n47 VDD1.n46 185
R787 VDD1.n34 VDD1.n33 185
R788 VDD1.n41 VDD1.n40 185
R789 VDD1.n39 VDD1.n38 185
R790 VDD1.n146 VDD1.n145 185
R791 VDD1.n148 VDD1.n147 185
R792 VDD1.n141 VDD1.n140 185
R793 VDD1.n154 VDD1.n153 185
R794 VDD1.n156 VDD1.n155 185
R795 VDD1.n137 VDD1.n136 185
R796 VDD1.n162 VDD1.n161 185
R797 VDD1.n164 VDD1.n163 185
R798 VDD1.n133 VDD1.n132 185
R799 VDD1.n170 VDD1.n169 185
R800 VDD1.n172 VDD1.n171 185
R801 VDD1.n129 VDD1.n128 185
R802 VDD1.n178 VDD1.n177 185
R803 VDD1.n180 VDD1.n179 185
R804 VDD1.n125 VDD1.n124 185
R805 VDD1.n187 VDD1.n186 185
R806 VDD1.n188 VDD1.n123 185
R807 VDD1.n190 VDD1.n189 185
R808 VDD1.n121 VDD1.n120 185
R809 VDD1.n196 VDD1.n195 185
R810 VDD1.n198 VDD1.n197 185
R811 VDD1.n117 VDD1.n116 185
R812 VDD1.n204 VDD1.n203 185
R813 VDD1.n206 VDD1.n205 185
R814 VDD1.n113 VDD1.n112 185
R815 VDD1.n212 VDD1.n211 185
R816 VDD1.n214 VDD1.n213 185
R817 VDD1.n37 VDD1.t5 147.659
R818 VDD1.n144 VDD1.t4 147.659
R819 VDD1.n104 VDD1.n103 104.615
R820 VDD1.n103 VDD1.n3 104.615
R821 VDD1.n96 VDD1.n3 104.615
R822 VDD1.n96 VDD1.n95 104.615
R823 VDD1.n95 VDD1.n7 104.615
R824 VDD1.n88 VDD1.n7 104.615
R825 VDD1.n88 VDD1.n87 104.615
R826 VDD1.n87 VDD1.n11 104.615
R827 VDD1.n16 VDD1.n11 104.615
R828 VDD1.n80 VDD1.n16 104.615
R829 VDD1.n80 VDD1.n79 104.615
R830 VDD1.n79 VDD1.n17 104.615
R831 VDD1.n72 VDD1.n17 104.615
R832 VDD1.n72 VDD1.n71 104.615
R833 VDD1.n71 VDD1.n21 104.615
R834 VDD1.n64 VDD1.n21 104.615
R835 VDD1.n64 VDD1.n63 104.615
R836 VDD1.n63 VDD1.n25 104.615
R837 VDD1.n56 VDD1.n25 104.615
R838 VDD1.n56 VDD1.n55 104.615
R839 VDD1.n55 VDD1.n29 104.615
R840 VDD1.n48 VDD1.n29 104.615
R841 VDD1.n48 VDD1.n47 104.615
R842 VDD1.n47 VDD1.n33 104.615
R843 VDD1.n40 VDD1.n33 104.615
R844 VDD1.n40 VDD1.n39 104.615
R845 VDD1.n147 VDD1.n146 104.615
R846 VDD1.n147 VDD1.n140 104.615
R847 VDD1.n154 VDD1.n140 104.615
R848 VDD1.n155 VDD1.n154 104.615
R849 VDD1.n155 VDD1.n136 104.615
R850 VDD1.n162 VDD1.n136 104.615
R851 VDD1.n163 VDD1.n162 104.615
R852 VDD1.n163 VDD1.n132 104.615
R853 VDD1.n170 VDD1.n132 104.615
R854 VDD1.n171 VDD1.n170 104.615
R855 VDD1.n171 VDD1.n128 104.615
R856 VDD1.n178 VDD1.n128 104.615
R857 VDD1.n179 VDD1.n178 104.615
R858 VDD1.n179 VDD1.n124 104.615
R859 VDD1.n187 VDD1.n124 104.615
R860 VDD1.n188 VDD1.n187 104.615
R861 VDD1.n189 VDD1.n188 104.615
R862 VDD1.n189 VDD1.n120 104.615
R863 VDD1.n196 VDD1.n120 104.615
R864 VDD1.n197 VDD1.n196 104.615
R865 VDD1.n197 VDD1.n116 104.615
R866 VDD1.n204 VDD1.n116 104.615
R867 VDD1.n205 VDD1.n204 104.615
R868 VDD1.n205 VDD1.n112 104.615
R869 VDD1.n212 VDD1.n112 104.615
R870 VDD1.n213 VDD1.n212 104.615
R871 VDD1.n219 VDD1.n218 59.5576
R872 VDD1.n221 VDD1.n220 58.8565
R873 VDD1.n221 VDD1.n219 52.5332
R874 VDD1.n39 VDD1.t5 52.3082
R875 VDD1.n146 VDD1.t4 52.3082
R876 VDD1 VDD1.n108 49.4463
R877 VDD1.n219 VDD1.n217 49.3327
R878 VDD1.n38 VDD1.n37 15.6677
R879 VDD1.n145 VDD1.n144 15.6677
R880 VDD1.n14 VDD1.n12 13.1884
R881 VDD1.n190 VDD1.n121 13.1884
R882 VDD1.n86 VDD1.n85 12.8005
R883 VDD1.n82 VDD1.n81 12.8005
R884 VDD1.n41 VDD1.n36 12.8005
R885 VDD1.n148 VDD1.n143 12.8005
R886 VDD1.n191 VDD1.n123 12.8005
R887 VDD1.n195 VDD1.n194 12.8005
R888 VDD1.n89 VDD1.n10 12.0247
R889 VDD1.n78 VDD1.n15 12.0247
R890 VDD1.n42 VDD1.n34 12.0247
R891 VDD1.n149 VDD1.n141 12.0247
R892 VDD1.n186 VDD1.n185 12.0247
R893 VDD1.n198 VDD1.n119 12.0247
R894 VDD1.n90 VDD1.n8 11.249
R895 VDD1.n77 VDD1.n18 11.249
R896 VDD1.n46 VDD1.n45 11.249
R897 VDD1.n153 VDD1.n152 11.249
R898 VDD1.n184 VDD1.n125 11.249
R899 VDD1.n199 VDD1.n117 11.249
R900 VDD1.n94 VDD1.n93 10.4732
R901 VDD1.n74 VDD1.n73 10.4732
R902 VDD1.n49 VDD1.n32 10.4732
R903 VDD1.n156 VDD1.n139 10.4732
R904 VDD1.n181 VDD1.n180 10.4732
R905 VDD1.n203 VDD1.n202 10.4732
R906 VDD1.n97 VDD1.n6 9.69747
R907 VDD1.n70 VDD1.n20 9.69747
R908 VDD1.n50 VDD1.n30 9.69747
R909 VDD1.n157 VDD1.n137 9.69747
R910 VDD1.n177 VDD1.n127 9.69747
R911 VDD1.n206 VDD1.n115 9.69747
R912 VDD1.n108 VDD1.n107 9.45567
R913 VDD1.n217 VDD1.n216 9.45567
R914 VDD1.n24 VDD1.n23 9.3005
R915 VDD1.n67 VDD1.n66 9.3005
R916 VDD1.n69 VDD1.n68 9.3005
R917 VDD1.n20 VDD1.n19 9.3005
R918 VDD1.n75 VDD1.n74 9.3005
R919 VDD1.n77 VDD1.n76 9.3005
R920 VDD1.n15 VDD1.n13 9.3005
R921 VDD1.n83 VDD1.n82 9.3005
R922 VDD1.n107 VDD1.n106 9.3005
R923 VDD1.n2 VDD1.n1 9.3005
R924 VDD1.n101 VDD1.n100 9.3005
R925 VDD1.n99 VDD1.n98 9.3005
R926 VDD1.n6 VDD1.n5 9.3005
R927 VDD1.n93 VDD1.n92 9.3005
R928 VDD1.n91 VDD1.n90 9.3005
R929 VDD1.n10 VDD1.n9 9.3005
R930 VDD1.n85 VDD1.n84 9.3005
R931 VDD1.n61 VDD1.n60 9.3005
R932 VDD1.n59 VDD1.n58 9.3005
R933 VDD1.n28 VDD1.n27 9.3005
R934 VDD1.n53 VDD1.n52 9.3005
R935 VDD1.n51 VDD1.n50 9.3005
R936 VDD1.n32 VDD1.n31 9.3005
R937 VDD1.n45 VDD1.n44 9.3005
R938 VDD1.n43 VDD1.n42 9.3005
R939 VDD1.n36 VDD1.n35 9.3005
R940 VDD1.n216 VDD1.n215 9.3005
R941 VDD1.n210 VDD1.n209 9.3005
R942 VDD1.n208 VDD1.n207 9.3005
R943 VDD1.n115 VDD1.n114 9.3005
R944 VDD1.n202 VDD1.n201 9.3005
R945 VDD1.n200 VDD1.n199 9.3005
R946 VDD1.n119 VDD1.n118 9.3005
R947 VDD1.n194 VDD1.n193 9.3005
R948 VDD1.n166 VDD1.n165 9.3005
R949 VDD1.n135 VDD1.n134 9.3005
R950 VDD1.n160 VDD1.n159 9.3005
R951 VDD1.n158 VDD1.n157 9.3005
R952 VDD1.n139 VDD1.n138 9.3005
R953 VDD1.n152 VDD1.n151 9.3005
R954 VDD1.n150 VDD1.n149 9.3005
R955 VDD1.n143 VDD1.n142 9.3005
R956 VDD1.n168 VDD1.n167 9.3005
R957 VDD1.n131 VDD1.n130 9.3005
R958 VDD1.n174 VDD1.n173 9.3005
R959 VDD1.n176 VDD1.n175 9.3005
R960 VDD1.n127 VDD1.n126 9.3005
R961 VDD1.n182 VDD1.n181 9.3005
R962 VDD1.n184 VDD1.n183 9.3005
R963 VDD1.n185 VDD1.n122 9.3005
R964 VDD1.n192 VDD1.n191 9.3005
R965 VDD1.n111 VDD1.n110 9.3005
R966 VDD1.n98 VDD1.n4 8.92171
R967 VDD1.n69 VDD1.n22 8.92171
R968 VDD1.n54 VDD1.n53 8.92171
R969 VDD1.n161 VDD1.n160 8.92171
R970 VDD1.n176 VDD1.n129 8.92171
R971 VDD1.n207 VDD1.n113 8.92171
R972 VDD1.n102 VDD1.n101 8.14595
R973 VDD1.n66 VDD1.n65 8.14595
R974 VDD1.n57 VDD1.n28 8.14595
R975 VDD1.n164 VDD1.n135 8.14595
R976 VDD1.n173 VDD1.n172 8.14595
R977 VDD1.n211 VDD1.n210 8.14595
R978 VDD1.n108 VDD1.n0 7.3702
R979 VDD1.n105 VDD1.n2 7.3702
R980 VDD1.n62 VDD1.n24 7.3702
R981 VDD1.n58 VDD1.n26 7.3702
R982 VDD1.n165 VDD1.n133 7.3702
R983 VDD1.n169 VDD1.n131 7.3702
R984 VDD1.n214 VDD1.n111 7.3702
R985 VDD1.n217 VDD1.n109 7.3702
R986 VDD1.n106 VDD1.n0 6.59444
R987 VDD1.n106 VDD1.n105 6.59444
R988 VDD1.n62 VDD1.n61 6.59444
R989 VDD1.n61 VDD1.n26 6.59444
R990 VDD1.n168 VDD1.n133 6.59444
R991 VDD1.n169 VDD1.n168 6.59444
R992 VDD1.n215 VDD1.n214 6.59444
R993 VDD1.n215 VDD1.n109 6.59444
R994 VDD1.n102 VDD1.n2 5.81868
R995 VDD1.n65 VDD1.n24 5.81868
R996 VDD1.n58 VDD1.n57 5.81868
R997 VDD1.n165 VDD1.n164 5.81868
R998 VDD1.n172 VDD1.n131 5.81868
R999 VDD1.n211 VDD1.n111 5.81868
R1000 VDD1.n101 VDD1.n4 5.04292
R1001 VDD1.n66 VDD1.n22 5.04292
R1002 VDD1.n54 VDD1.n28 5.04292
R1003 VDD1.n161 VDD1.n135 5.04292
R1004 VDD1.n173 VDD1.n129 5.04292
R1005 VDD1.n210 VDD1.n113 5.04292
R1006 VDD1.n37 VDD1.n35 4.38563
R1007 VDD1.n144 VDD1.n142 4.38563
R1008 VDD1.n98 VDD1.n97 4.26717
R1009 VDD1.n70 VDD1.n69 4.26717
R1010 VDD1.n53 VDD1.n30 4.26717
R1011 VDD1.n160 VDD1.n137 4.26717
R1012 VDD1.n177 VDD1.n176 4.26717
R1013 VDD1.n207 VDD1.n206 4.26717
R1014 VDD1.n94 VDD1.n6 3.49141
R1015 VDD1.n73 VDD1.n20 3.49141
R1016 VDD1.n50 VDD1.n49 3.49141
R1017 VDD1.n157 VDD1.n156 3.49141
R1018 VDD1.n180 VDD1.n127 3.49141
R1019 VDD1.n203 VDD1.n115 3.49141
R1020 VDD1.n93 VDD1.n8 2.71565
R1021 VDD1.n74 VDD1.n18 2.71565
R1022 VDD1.n46 VDD1.n32 2.71565
R1023 VDD1.n153 VDD1.n139 2.71565
R1024 VDD1.n181 VDD1.n125 2.71565
R1025 VDD1.n202 VDD1.n117 2.71565
R1026 VDD1.n90 VDD1.n89 1.93989
R1027 VDD1.n78 VDD1.n77 1.93989
R1028 VDD1.n45 VDD1.n34 1.93989
R1029 VDD1.n152 VDD1.n141 1.93989
R1030 VDD1.n186 VDD1.n184 1.93989
R1031 VDD1.n199 VDD1.n198 1.93989
R1032 VDD1.n86 VDD1.n10 1.16414
R1033 VDD1.n81 VDD1.n15 1.16414
R1034 VDD1.n42 VDD1.n41 1.16414
R1035 VDD1.n149 VDD1.n148 1.16414
R1036 VDD1.n185 VDD1.n123 1.16414
R1037 VDD1.n195 VDD1.n119 1.16414
R1038 VDD1.n220 VDD1.t2 1.01122
R1039 VDD1.n220 VDD1.t3 1.01122
R1040 VDD1.n218 VDD1.t1 1.01122
R1041 VDD1.n218 VDD1.t0 1.01122
R1042 VDD1 VDD1.n221 0.698776
R1043 VDD1.n85 VDD1.n12 0.388379
R1044 VDD1.n82 VDD1.n14 0.388379
R1045 VDD1.n38 VDD1.n36 0.388379
R1046 VDD1.n145 VDD1.n143 0.388379
R1047 VDD1.n191 VDD1.n190 0.388379
R1048 VDD1.n194 VDD1.n121 0.388379
R1049 VDD1.n107 VDD1.n1 0.155672
R1050 VDD1.n100 VDD1.n1 0.155672
R1051 VDD1.n100 VDD1.n99 0.155672
R1052 VDD1.n99 VDD1.n5 0.155672
R1053 VDD1.n92 VDD1.n5 0.155672
R1054 VDD1.n92 VDD1.n91 0.155672
R1055 VDD1.n91 VDD1.n9 0.155672
R1056 VDD1.n84 VDD1.n9 0.155672
R1057 VDD1.n84 VDD1.n83 0.155672
R1058 VDD1.n83 VDD1.n13 0.155672
R1059 VDD1.n76 VDD1.n13 0.155672
R1060 VDD1.n76 VDD1.n75 0.155672
R1061 VDD1.n75 VDD1.n19 0.155672
R1062 VDD1.n68 VDD1.n19 0.155672
R1063 VDD1.n68 VDD1.n67 0.155672
R1064 VDD1.n67 VDD1.n23 0.155672
R1065 VDD1.n60 VDD1.n23 0.155672
R1066 VDD1.n60 VDD1.n59 0.155672
R1067 VDD1.n59 VDD1.n27 0.155672
R1068 VDD1.n52 VDD1.n27 0.155672
R1069 VDD1.n52 VDD1.n51 0.155672
R1070 VDD1.n51 VDD1.n31 0.155672
R1071 VDD1.n44 VDD1.n31 0.155672
R1072 VDD1.n44 VDD1.n43 0.155672
R1073 VDD1.n43 VDD1.n35 0.155672
R1074 VDD1.n150 VDD1.n142 0.155672
R1075 VDD1.n151 VDD1.n150 0.155672
R1076 VDD1.n151 VDD1.n138 0.155672
R1077 VDD1.n158 VDD1.n138 0.155672
R1078 VDD1.n159 VDD1.n158 0.155672
R1079 VDD1.n159 VDD1.n134 0.155672
R1080 VDD1.n166 VDD1.n134 0.155672
R1081 VDD1.n167 VDD1.n166 0.155672
R1082 VDD1.n167 VDD1.n130 0.155672
R1083 VDD1.n174 VDD1.n130 0.155672
R1084 VDD1.n175 VDD1.n174 0.155672
R1085 VDD1.n175 VDD1.n126 0.155672
R1086 VDD1.n182 VDD1.n126 0.155672
R1087 VDD1.n183 VDD1.n182 0.155672
R1088 VDD1.n183 VDD1.n122 0.155672
R1089 VDD1.n192 VDD1.n122 0.155672
R1090 VDD1.n193 VDD1.n192 0.155672
R1091 VDD1.n193 VDD1.n118 0.155672
R1092 VDD1.n200 VDD1.n118 0.155672
R1093 VDD1.n201 VDD1.n200 0.155672
R1094 VDD1.n201 VDD1.n114 0.155672
R1095 VDD1.n208 VDD1.n114 0.155672
R1096 VDD1.n209 VDD1.n208 0.155672
R1097 VDD1.n209 VDD1.n110 0.155672
R1098 VDD1.n216 VDD1.n110 0.155672
R1099 B.n1094 B.n1093 585
R1100 B.n1095 B.n1094 585
R1101 B.n437 B.n160 585
R1102 B.n436 B.n435 585
R1103 B.n434 B.n433 585
R1104 B.n432 B.n431 585
R1105 B.n430 B.n429 585
R1106 B.n428 B.n427 585
R1107 B.n426 B.n425 585
R1108 B.n424 B.n423 585
R1109 B.n422 B.n421 585
R1110 B.n420 B.n419 585
R1111 B.n418 B.n417 585
R1112 B.n416 B.n415 585
R1113 B.n414 B.n413 585
R1114 B.n412 B.n411 585
R1115 B.n410 B.n409 585
R1116 B.n408 B.n407 585
R1117 B.n406 B.n405 585
R1118 B.n404 B.n403 585
R1119 B.n402 B.n401 585
R1120 B.n400 B.n399 585
R1121 B.n398 B.n397 585
R1122 B.n396 B.n395 585
R1123 B.n394 B.n393 585
R1124 B.n392 B.n391 585
R1125 B.n390 B.n389 585
R1126 B.n388 B.n387 585
R1127 B.n386 B.n385 585
R1128 B.n384 B.n383 585
R1129 B.n382 B.n381 585
R1130 B.n380 B.n379 585
R1131 B.n378 B.n377 585
R1132 B.n376 B.n375 585
R1133 B.n374 B.n373 585
R1134 B.n372 B.n371 585
R1135 B.n370 B.n369 585
R1136 B.n368 B.n367 585
R1137 B.n366 B.n365 585
R1138 B.n364 B.n363 585
R1139 B.n362 B.n361 585
R1140 B.n360 B.n359 585
R1141 B.n358 B.n357 585
R1142 B.n356 B.n355 585
R1143 B.n354 B.n353 585
R1144 B.n352 B.n351 585
R1145 B.n350 B.n349 585
R1146 B.n348 B.n347 585
R1147 B.n346 B.n345 585
R1148 B.n344 B.n343 585
R1149 B.n342 B.n341 585
R1150 B.n340 B.n339 585
R1151 B.n338 B.n337 585
R1152 B.n336 B.n335 585
R1153 B.n334 B.n333 585
R1154 B.n332 B.n331 585
R1155 B.n330 B.n329 585
R1156 B.n328 B.n327 585
R1157 B.n326 B.n325 585
R1158 B.n324 B.n323 585
R1159 B.n322 B.n321 585
R1160 B.n320 B.n319 585
R1161 B.n318 B.n317 585
R1162 B.n316 B.n315 585
R1163 B.n314 B.n313 585
R1164 B.n311 B.n310 585
R1165 B.n309 B.n308 585
R1166 B.n307 B.n306 585
R1167 B.n305 B.n304 585
R1168 B.n303 B.n302 585
R1169 B.n301 B.n300 585
R1170 B.n299 B.n298 585
R1171 B.n297 B.n296 585
R1172 B.n295 B.n294 585
R1173 B.n293 B.n292 585
R1174 B.n291 B.n290 585
R1175 B.n289 B.n288 585
R1176 B.n287 B.n286 585
R1177 B.n285 B.n284 585
R1178 B.n283 B.n282 585
R1179 B.n281 B.n280 585
R1180 B.n279 B.n278 585
R1181 B.n277 B.n276 585
R1182 B.n275 B.n274 585
R1183 B.n273 B.n272 585
R1184 B.n271 B.n270 585
R1185 B.n269 B.n268 585
R1186 B.n267 B.n266 585
R1187 B.n265 B.n264 585
R1188 B.n263 B.n262 585
R1189 B.n261 B.n260 585
R1190 B.n259 B.n258 585
R1191 B.n257 B.n256 585
R1192 B.n255 B.n254 585
R1193 B.n253 B.n252 585
R1194 B.n251 B.n250 585
R1195 B.n249 B.n248 585
R1196 B.n247 B.n246 585
R1197 B.n245 B.n244 585
R1198 B.n243 B.n242 585
R1199 B.n241 B.n240 585
R1200 B.n239 B.n238 585
R1201 B.n237 B.n236 585
R1202 B.n235 B.n234 585
R1203 B.n233 B.n232 585
R1204 B.n231 B.n230 585
R1205 B.n229 B.n228 585
R1206 B.n227 B.n226 585
R1207 B.n225 B.n224 585
R1208 B.n223 B.n222 585
R1209 B.n221 B.n220 585
R1210 B.n219 B.n218 585
R1211 B.n217 B.n216 585
R1212 B.n215 B.n214 585
R1213 B.n213 B.n212 585
R1214 B.n211 B.n210 585
R1215 B.n209 B.n208 585
R1216 B.n207 B.n206 585
R1217 B.n205 B.n204 585
R1218 B.n203 B.n202 585
R1219 B.n201 B.n200 585
R1220 B.n199 B.n198 585
R1221 B.n197 B.n196 585
R1222 B.n195 B.n194 585
R1223 B.n193 B.n192 585
R1224 B.n191 B.n190 585
R1225 B.n189 B.n188 585
R1226 B.n187 B.n186 585
R1227 B.n185 B.n184 585
R1228 B.n183 B.n182 585
R1229 B.n181 B.n180 585
R1230 B.n179 B.n178 585
R1231 B.n177 B.n176 585
R1232 B.n175 B.n174 585
R1233 B.n173 B.n172 585
R1234 B.n171 B.n170 585
R1235 B.n169 B.n168 585
R1236 B.n167 B.n166 585
R1237 B.n1092 B.n91 585
R1238 B.n1096 B.n91 585
R1239 B.n1091 B.n90 585
R1240 B.n1097 B.n90 585
R1241 B.n1090 B.n1089 585
R1242 B.n1089 B.n86 585
R1243 B.n1088 B.n85 585
R1244 B.n1103 B.n85 585
R1245 B.n1087 B.n84 585
R1246 B.n1104 B.n84 585
R1247 B.n1086 B.n83 585
R1248 B.n1105 B.n83 585
R1249 B.n1085 B.n1084 585
R1250 B.n1084 B.n79 585
R1251 B.n1083 B.n78 585
R1252 B.n1111 B.n78 585
R1253 B.n1082 B.n77 585
R1254 B.n1112 B.n77 585
R1255 B.n1081 B.n76 585
R1256 B.n1113 B.n76 585
R1257 B.n1080 B.n1079 585
R1258 B.n1079 B.n72 585
R1259 B.n1078 B.n71 585
R1260 B.n1119 B.n71 585
R1261 B.n1077 B.n70 585
R1262 B.n1120 B.n70 585
R1263 B.n1076 B.n69 585
R1264 B.n1121 B.n69 585
R1265 B.n1075 B.n1074 585
R1266 B.n1074 B.n65 585
R1267 B.n1073 B.n64 585
R1268 B.n1127 B.n64 585
R1269 B.n1072 B.n63 585
R1270 B.n1128 B.n63 585
R1271 B.n1071 B.n62 585
R1272 B.n1129 B.n62 585
R1273 B.n1070 B.n1069 585
R1274 B.n1069 B.n58 585
R1275 B.n1068 B.n57 585
R1276 B.n1135 B.n57 585
R1277 B.n1067 B.n56 585
R1278 B.n1136 B.n56 585
R1279 B.n1066 B.n55 585
R1280 B.n1137 B.n55 585
R1281 B.n1065 B.n1064 585
R1282 B.n1064 B.n54 585
R1283 B.n1063 B.n50 585
R1284 B.n1143 B.n50 585
R1285 B.n1062 B.n49 585
R1286 B.n1144 B.n49 585
R1287 B.n1061 B.n48 585
R1288 B.n1145 B.n48 585
R1289 B.n1060 B.n1059 585
R1290 B.n1059 B.n44 585
R1291 B.n1058 B.n43 585
R1292 B.n1151 B.n43 585
R1293 B.n1057 B.n42 585
R1294 B.n1152 B.n42 585
R1295 B.n1056 B.n41 585
R1296 B.n1153 B.n41 585
R1297 B.n1055 B.n1054 585
R1298 B.n1054 B.n37 585
R1299 B.n1053 B.n36 585
R1300 B.n1159 B.n36 585
R1301 B.n1052 B.n35 585
R1302 B.n1160 B.n35 585
R1303 B.n1051 B.n34 585
R1304 B.n1161 B.n34 585
R1305 B.n1050 B.n1049 585
R1306 B.n1049 B.n30 585
R1307 B.n1048 B.n29 585
R1308 B.n1167 B.n29 585
R1309 B.n1047 B.n28 585
R1310 B.n1168 B.n28 585
R1311 B.n1046 B.n27 585
R1312 B.n1169 B.n27 585
R1313 B.n1045 B.n1044 585
R1314 B.n1044 B.n23 585
R1315 B.n1043 B.n22 585
R1316 B.n1175 B.n22 585
R1317 B.n1042 B.n21 585
R1318 B.n1176 B.n21 585
R1319 B.n1041 B.n20 585
R1320 B.n1177 B.n20 585
R1321 B.n1040 B.n1039 585
R1322 B.n1039 B.n19 585
R1323 B.n1038 B.n15 585
R1324 B.n1183 B.n15 585
R1325 B.n1037 B.n14 585
R1326 B.n1184 B.n14 585
R1327 B.n1036 B.n13 585
R1328 B.n1185 B.n13 585
R1329 B.n1035 B.n1034 585
R1330 B.n1034 B.n12 585
R1331 B.n1033 B.n1032 585
R1332 B.n1033 B.n8 585
R1333 B.n1031 B.n7 585
R1334 B.n1192 B.n7 585
R1335 B.n1030 B.n6 585
R1336 B.n1193 B.n6 585
R1337 B.n1029 B.n5 585
R1338 B.n1194 B.n5 585
R1339 B.n1028 B.n1027 585
R1340 B.n1027 B.n4 585
R1341 B.n1026 B.n438 585
R1342 B.n1026 B.n1025 585
R1343 B.n1016 B.n439 585
R1344 B.n440 B.n439 585
R1345 B.n1018 B.n1017 585
R1346 B.n1019 B.n1018 585
R1347 B.n1015 B.n445 585
R1348 B.n445 B.n444 585
R1349 B.n1014 B.n1013 585
R1350 B.n1013 B.n1012 585
R1351 B.n447 B.n446 585
R1352 B.n1005 B.n447 585
R1353 B.n1004 B.n1003 585
R1354 B.n1006 B.n1004 585
R1355 B.n1002 B.n452 585
R1356 B.n452 B.n451 585
R1357 B.n1001 B.n1000 585
R1358 B.n1000 B.n999 585
R1359 B.n454 B.n453 585
R1360 B.n455 B.n454 585
R1361 B.n992 B.n991 585
R1362 B.n993 B.n992 585
R1363 B.n990 B.n460 585
R1364 B.n460 B.n459 585
R1365 B.n989 B.n988 585
R1366 B.n988 B.n987 585
R1367 B.n462 B.n461 585
R1368 B.n463 B.n462 585
R1369 B.n980 B.n979 585
R1370 B.n981 B.n980 585
R1371 B.n978 B.n467 585
R1372 B.n471 B.n467 585
R1373 B.n977 B.n976 585
R1374 B.n976 B.n975 585
R1375 B.n469 B.n468 585
R1376 B.n470 B.n469 585
R1377 B.n968 B.n967 585
R1378 B.n969 B.n968 585
R1379 B.n966 B.n476 585
R1380 B.n476 B.n475 585
R1381 B.n965 B.n964 585
R1382 B.n964 B.n963 585
R1383 B.n478 B.n477 585
R1384 B.n479 B.n478 585
R1385 B.n956 B.n955 585
R1386 B.n957 B.n956 585
R1387 B.n954 B.n484 585
R1388 B.n484 B.n483 585
R1389 B.n953 B.n952 585
R1390 B.n952 B.n951 585
R1391 B.n486 B.n485 585
R1392 B.n944 B.n486 585
R1393 B.n943 B.n942 585
R1394 B.n945 B.n943 585
R1395 B.n941 B.n491 585
R1396 B.n491 B.n490 585
R1397 B.n940 B.n939 585
R1398 B.n939 B.n938 585
R1399 B.n493 B.n492 585
R1400 B.n494 B.n493 585
R1401 B.n931 B.n930 585
R1402 B.n932 B.n931 585
R1403 B.n929 B.n499 585
R1404 B.n499 B.n498 585
R1405 B.n928 B.n927 585
R1406 B.n927 B.n926 585
R1407 B.n501 B.n500 585
R1408 B.n502 B.n501 585
R1409 B.n919 B.n918 585
R1410 B.n920 B.n919 585
R1411 B.n917 B.n507 585
R1412 B.n507 B.n506 585
R1413 B.n916 B.n915 585
R1414 B.n915 B.n914 585
R1415 B.n509 B.n508 585
R1416 B.n510 B.n509 585
R1417 B.n907 B.n906 585
R1418 B.n908 B.n907 585
R1419 B.n905 B.n514 585
R1420 B.n518 B.n514 585
R1421 B.n904 B.n903 585
R1422 B.n903 B.n902 585
R1423 B.n516 B.n515 585
R1424 B.n517 B.n516 585
R1425 B.n895 B.n894 585
R1426 B.n896 B.n895 585
R1427 B.n893 B.n523 585
R1428 B.n523 B.n522 585
R1429 B.n892 B.n891 585
R1430 B.n891 B.n890 585
R1431 B.n525 B.n524 585
R1432 B.n526 B.n525 585
R1433 B.n883 B.n882 585
R1434 B.n884 B.n883 585
R1435 B.n881 B.n531 585
R1436 B.n531 B.n530 585
R1437 B.n875 B.n874 585
R1438 B.n873 B.n601 585
R1439 B.n872 B.n600 585
R1440 B.n877 B.n600 585
R1441 B.n871 B.n870 585
R1442 B.n869 B.n868 585
R1443 B.n867 B.n866 585
R1444 B.n865 B.n864 585
R1445 B.n863 B.n862 585
R1446 B.n861 B.n860 585
R1447 B.n859 B.n858 585
R1448 B.n857 B.n856 585
R1449 B.n855 B.n854 585
R1450 B.n853 B.n852 585
R1451 B.n851 B.n850 585
R1452 B.n849 B.n848 585
R1453 B.n847 B.n846 585
R1454 B.n845 B.n844 585
R1455 B.n843 B.n842 585
R1456 B.n841 B.n840 585
R1457 B.n839 B.n838 585
R1458 B.n837 B.n836 585
R1459 B.n835 B.n834 585
R1460 B.n833 B.n832 585
R1461 B.n831 B.n830 585
R1462 B.n829 B.n828 585
R1463 B.n827 B.n826 585
R1464 B.n825 B.n824 585
R1465 B.n823 B.n822 585
R1466 B.n821 B.n820 585
R1467 B.n819 B.n818 585
R1468 B.n817 B.n816 585
R1469 B.n815 B.n814 585
R1470 B.n813 B.n812 585
R1471 B.n811 B.n810 585
R1472 B.n809 B.n808 585
R1473 B.n807 B.n806 585
R1474 B.n805 B.n804 585
R1475 B.n803 B.n802 585
R1476 B.n801 B.n800 585
R1477 B.n799 B.n798 585
R1478 B.n797 B.n796 585
R1479 B.n795 B.n794 585
R1480 B.n793 B.n792 585
R1481 B.n791 B.n790 585
R1482 B.n789 B.n788 585
R1483 B.n787 B.n786 585
R1484 B.n785 B.n784 585
R1485 B.n783 B.n782 585
R1486 B.n781 B.n780 585
R1487 B.n779 B.n778 585
R1488 B.n777 B.n776 585
R1489 B.n775 B.n774 585
R1490 B.n773 B.n772 585
R1491 B.n771 B.n770 585
R1492 B.n769 B.n768 585
R1493 B.n767 B.n766 585
R1494 B.n765 B.n764 585
R1495 B.n763 B.n762 585
R1496 B.n761 B.n760 585
R1497 B.n759 B.n758 585
R1498 B.n757 B.n756 585
R1499 B.n755 B.n754 585
R1500 B.n753 B.n752 585
R1501 B.n751 B.n750 585
R1502 B.n748 B.n747 585
R1503 B.n746 B.n745 585
R1504 B.n744 B.n743 585
R1505 B.n742 B.n741 585
R1506 B.n740 B.n739 585
R1507 B.n738 B.n737 585
R1508 B.n736 B.n735 585
R1509 B.n734 B.n733 585
R1510 B.n732 B.n731 585
R1511 B.n730 B.n729 585
R1512 B.n728 B.n727 585
R1513 B.n726 B.n725 585
R1514 B.n724 B.n723 585
R1515 B.n722 B.n721 585
R1516 B.n720 B.n719 585
R1517 B.n718 B.n717 585
R1518 B.n716 B.n715 585
R1519 B.n714 B.n713 585
R1520 B.n712 B.n711 585
R1521 B.n710 B.n709 585
R1522 B.n708 B.n707 585
R1523 B.n706 B.n705 585
R1524 B.n704 B.n703 585
R1525 B.n702 B.n701 585
R1526 B.n700 B.n699 585
R1527 B.n698 B.n697 585
R1528 B.n696 B.n695 585
R1529 B.n694 B.n693 585
R1530 B.n692 B.n691 585
R1531 B.n690 B.n689 585
R1532 B.n688 B.n687 585
R1533 B.n686 B.n685 585
R1534 B.n684 B.n683 585
R1535 B.n682 B.n681 585
R1536 B.n680 B.n679 585
R1537 B.n678 B.n677 585
R1538 B.n676 B.n675 585
R1539 B.n674 B.n673 585
R1540 B.n672 B.n671 585
R1541 B.n670 B.n669 585
R1542 B.n668 B.n667 585
R1543 B.n666 B.n665 585
R1544 B.n664 B.n663 585
R1545 B.n662 B.n661 585
R1546 B.n660 B.n659 585
R1547 B.n658 B.n657 585
R1548 B.n656 B.n655 585
R1549 B.n654 B.n653 585
R1550 B.n652 B.n651 585
R1551 B.n650 B.n649 585
R1552 B.n648 B.n647 585
R1553 B.n646 B.n645 585
R1554 B.n644 B.n643 585
R1555 B.n642 B.n641 585
R1556 B.n640 B.n639 585
R1557 B.n638 B.n637 585
R1558 B.n636 B.n635 585
R1559 B.n634 B.n633 585
R1560 B.n632 B.n631 585
R1561 B.n630 B.n629 585
R1562 B.n628 B.n627 585
R1563 B.n626 B.n625 585
R1564 B.n624 B.n623 585
R1565 B.n622 B.n621 585
R1566 B.n620 B.n619 585
R1567 B.n618 B.n617 585
R1568 B.n616 B.n615 585
R1569 B.n614 B.n613 585
R1570 B.n612 B.n611 585
R1571 B.n610 B.n609 585
R1572 B.n608 B.n607 585
R1573 B.n533 B.n532 585
R1574 B.n880 B.n879 585
R1575 B.n529 B.n528 585
R1576 B.n530 B.n529 585
R1577 B.n886 B.n885 585
R1578 B.n885 B.n884 585
R1579 B.n887 B.n527 585
R1580 B.n527 B.n526 585
R1581 B.n889 B.n888 585
R1582 B.n890 B.n889 585
R1583 B.n521 B.n520 585
R1584 B.n522 B.n521 585
R1585 B.n898 B.n897 585
R1586 B.n897 B.n896 585
R1587 B.n899 B.n519 585
R1588 B.n519 B.n517 585
R1589 B.n901 B.n900 585
R1590 B.n902 B.n901 585
R1591 B.n513 B.n512 585
R1592 B.n518 B.n513 585
R1593 B.n910 B.n909 585
R1594 B.n909 B.n908 585
R1595 B.n911 B.n511 585
R1596 B.n511 B.n510 585
R1597 B.n913 B.n912 585
R1598 B.n914 B.n913 585
R1599 B.n505 B.n504 585
R1600 B.n506 B.n505 585
R1601 B.n922 B.n921 585
R1602 B.n921 B.n920 585
R1603 B.n923 B.n503 585
R1604 B.n503 B.n502 585
R1605 B.n925 B.n924 585
R1606 B.n926 B.n925 585
R1607 B.n497 B.n496 585
R1608 B.n498 B.n497 585
R1609 B.n934 B.n933 585
R1610 B.n933 B.n932 585
R1611 B.n935 B.n495 585
R1612 B.n495 B.n494 585
R1613 B.n937 B.n936 585
R1614 B.n938 B.n937 585
R1615 B.n489 B.n488 585
R1616 B.n490 B.n489 585
R1617 B.n947 B.n946 585
R1618 B.n946 B.n945 585
R1619 B.n948 B.n487 585
R1620 B.n944 B.n487 585
R1621 B.n950 B.n949 585
R1622 B.n951 B.n950 585
R1623 B.n482 B.n481 585
R1624 B.n483 B.n482 585
R1625 B.n959 B.n958 585
R1626 B.n958 B.n957 585
R1627 B.n960 B.n480 585
R1628 B.n480 B.n479 585
R1629 B.n962 B.n961 585
R1630 B.n963 B.n962 585
R1631 B.n474 B.n473 585
R1632 B.n475 B.n474 585
R1633 B.n971 B.n970 585
R1634 B.n970 B.n969 585
R1635 B.n972 B.n472 585
R1636 B.n472 B.n470 585
R1637 B.n974 B.n973 585
R1638 B.n975 B.n974 585
R1639 B.n466 B.n465 585
R1640 B.n471 B.n466 585
R1641 B.n983 B.n982 585
R1642 B.n982 B.n981 585
R1643 B.n984 B.n464 585
R1644 B.n464 B.n463 585
R1645 B.n986 B.n985 585
R1646 B.n987 B.n986 585
R1647 B.n458 B.n457 585
R1648 B.n459 B.n458 585
R1649 B.n995 B.n994 585
R1650 B.n994 B.n993 585
R1651 B.n996 B.n456 585
R1652 B.n456 B.n455 585
R1653 B.n998 B.n997 585
R1654 B.n999 B.n998 585
R1655 B.n450 B.n449 585
R1656 B.n451 B.n450 585
R1657 B.n1008 B.n1007 585
R1658 B.n1007 B.n1006 585
R1659 B.n1009 B.n448 585
R1660 B.n1005 B.n448 585
R1661 B.n1011 B.n1010 585
R1662 B.n1012 B.n1011 585
R1663 B.n443 B.n442 585
R1664 B.n444 B.n443 585
R1665 B.n1021 B.n1020 585
R1666 B.n1020 B.n1019 585
R1667 B.n1022 B.n441 585
R1668 B.n441 B.n440 585
R1669 B.n1024 B.n1023 585
R1670 B.n1025 B.n1024 585
R1671 B.n3 B.n0 585
R1672 B.n4 B.n3 585
R1673 B.n1191 B.n1 585
R1674 B.n1192 B.n1191 585
R1675 B.n1190 B.n1189 585
R1676 B.n1190 B.n8 585
R1677 B.n1188 B.n9 585
R1678 B.n12 B.n9 585
R1679 B.n1187 B.n1186 585
R1680 B.n1186 B.n1185 585
R1681 B.n11 B.n10 585
R1682 B.n1184 B.n11 585
R1683 B.n1182 B.n1181 585
R1684 B.n1183 B.n1182 585
R1685 B.n1180 B.n16 585
R1686 B.n19 B.n16 585
R1687 B.n1179 B.n1178 585
R1688 B.n1178 B.n1177 585
R1689 B.n18 B.n17 585
R1690 B.n1176 B.n18 585
R1691 B.n1174 B.n1173 585
R1692 B.n1175 B.n1174 585
R1693 B.n1172 B.n24 585
R1694 B.n24 B.n23 585
R1695 B.n1171 B.n1170 585
R1696 B.n1170 B.n1169 585
R1697 B.n26 B.n25 585
R1698 B.n1168 B.n26 585
R1699 B.n1166 B.n1165 585
R1700 B.n1167 B.n1166 585
R1701 B.n1164 B.n31 585
R1702 B.n31 B.n30 585
R1703 B.n1163 B.n1162 585
R1704 B.n1162 B.n1161 585
R1705 B.n33 B.n32 585
R1706 B.n1160 B.n33 585
R1707 B.n1158 B.n1157 585
R1708 B.n1159 B.n1158 585
R1709 B.n1156 B.n38 585
R1710 B.n38 B.n37 585
R1711 B.n1155 B.n1154 585
R1712 B.n1154 B.n1153 585
R1713 B.n40 B.n39 585
R1714 B.n1152 B.n40 585
R1715 B.n1150 B.n1149 585
R1716 B.n1151 B.n1150 585
R1717 B.n1148 B.n45 585
R1718 B.n45 B.n44 585
R1719 B.n1147 B.n1146 585
R1720 B.n1146 B.n1145 585
R1721 B.n47 B.n46 585
R1722 B.n1144 B.n47 585
R1723 B.n1142 B.n1141 585
R1724 B.n1143 B.n1142 585
R1725 B.n1140 B.n51 585
R1726 B.n54 B.n51 585
R1727 B.n1139 B.n1138 585
R1728 B.n1138 B.n1137 585
R1729 B.n53 B.n52 585
R1730 B.n1136 B.n53 585
R1731 B.n1134 B.n1133 585
R1732 B.n1135 B.n1134 585
R1733 B.n1132 B.n59 585
R1734 B.n59 B.n58 585
R1735 B.n1131 B.n1130 585
R1736 B.n1130 B.n1129 585
R1737 B.n61 B.n60 585
R1738 B.n1128 B.n61 585
R1739 B.n1126 B.n1125 585
R1740 B.n1127 B.n1126 585
R1741 B.n1124 B.n66 585
R1742 B.n66 B.n65 585
R1743 B.n1123 B.n1122 585
R1744 B.n1122 B.n1121 585
R1745 B.n68 B.n67 585
R1746 B.n1120 B.n68 585
R1747 B.n1118 B.n1117 585
R1748 B.n1119 B.n1118 585
R1749 B.n1116 B.n73 585
R1750 B.n73 B.n72 585
R1751 B.n1115 B.n1114 585
R1752 B.n1114 B.n1113 585
R1753 B.n75 B.n74 585
R1754 B.n1112 B.n75 585
R1755 B.n1110 B.n1109 585
R1756 B.n1111 B.n1110 585
R1757 B.n1108 B.n80 585
R1758 B.n80 B.n79 585
R1759 B.n1107 B.n1106 585
R1760 B.n1106 B.n1105 585
R1761 B.n82 B.n81 585
R1762 B.n1104 B.n82 585
R1763 B.n1102 B.n1101 585
R1764 B.n1103 B.n1102 585
R1765 B.n1100 B.n87 585
R1766 B.n87 B.n86 585
R1767 B.n1099 B.n1098 585
R1768 B.n1098 B.n1097 585
R1769 B.n89 B.n88 585
R1770 B.n1096 B.n89 585
R1771 B.n1195 B.n1194 585
R1772 B.n1193 B.n2 585
R1773 B.n166 B.n89 521.33
R1774 B.n1094 B.n91 521.33
R1775 B.n879 B.n531 521.33
R1776 B.n875 B.n529 521.33
R1777 B.n161 B.t18 481.05
R1778 B.n604 B.t16 481.05
R1779 B.n163 B.t8 481.05
R1780 B.n602 B.t13 481.05
R1781 B.n162 B.t19 412.978
R1782 B.n605 B.t15 412.978
R1783 B.n164 B.t9 412.978
R1784 B.n603 B.t12 412.978
R1785 B.n163 B.t6 357.247
R1786 B.n161 B.t17 357.247
R1787 B.n604 B.t14 357.247
R1788 B.n602 B.t10 357.247
R1789 B.n1095 B.n159 256.663
R1790 B.n1095 B.n158 256.663
R1791 B.n1095 B.n157 256.663
R1792 B.n1095 B.n156 256.663
R1793 B.n1095 B.n155 256.663
R1794 B.n1095 B.n154 256.663
R1795 B.n1095 B.n153 256.663
R1796 B.n1095 B.n152 256.663
R1797 B.n1095 B.n151 256.663
R1798 B.n1095 B.n150 256.663
R1799 B.n1095 B.n149 256.663
R1800 B.n1095 B.n148 256.663
R1801 B.n1095 B.n147 256.663
R1802 B.n1095 B.n146 256.663
R1803 B.n1095 B.n145 256.663
R1804 B.n1095 B.n144 256.663
R1805 B.n1095 B.n143 256.663
R1806 B.n1095 B.n142 256.663
R1807 B.n1095 B.n141 256.663
R1808 B.n1095 B.n140 256.663
R1809 B.n1095 B.n139 256.663
R1810 B.n1095 B.n138 256.663
R1811 B.n1095 B.n137 256.663
R1812 B.n1095 B.n136 256.663
R1813 B.n1095 B.n135 256.663
R1814 B.n1095 B.n134 256.663
R1815 B.n1095 B.n133 256.663
R1816 B.n1095 B.n132 256.663
R1817 B.n1095 B.n131 256.663
R1818 B.n1095 B.n130 256.663
R1819 B.n1095 B.n129 256.663
R1820 B.n1095 B.n128 256.663
R1821 B.n1095 B.n127 256.663
R1822 B.n1095 B.n126 256.663
R1823 B.n1095 B.n125 256.663
R1824 B.n1095 B.n124 256.663
R1825 B.n1095 B.n123 256.663
R1826 B.n1095 B.n122 256.663
R1827 B.n1095 B.n121 256.663
R1828 B.n1095 B.n120 256.663
R1829 B.n1095 B.n119 256.663
R1830 B.n1095 B.n118 256.663
R1831 B.n1095 B.n117 256.663
R1832 B.n1095 B.n116 256.663
R1833 B.n1095 B.n115 256.663
R1834 B.n1095 B.n114 256.663
R1835 B.n1095 B.n113 256.663
R1836 B.n1095 B.n112 256.663
R1837 B.n1095 B.n111 256.663
R1838 B.n1095 B.n110 256.663
R1839 B.n1095 B.n109 256.663
R1840 B.n1095 B.n108 256.663
R1841 B.n1095 B.n107 256.663
R1842 B.n1095 B.n106 256.663
R1843 B.n1095 B.n105 256.663
R1844 B.n1095 B.n104 256.663
R1845 B.n1095 B.n103 256.663
R1846 B.n1095 B.n102 256.663
R1847 B.n1095 B.n101 256.663
R1848 B.n1095 B.n100 256.663
R1849 B.n1095 B.n99 256.663
R1850 B.n1095 B.n98 256.663
R1851 B.n1095 B.n97 256.663
R1852 B.n1095 B.n96 256.663
R1853 B.n1095 B.n95 256.663
R1854 B.n1095 B.n94 256.663
R1855 B.n1095 B.n93 256.663
R1856 B.n1095 B.n92 256.663
R1857 B.n877 B.n876 256.663
R1858 B.n877 B.n534 256.663
R1859 B.n877 B.n535 256.663
R1860 B.n877 B.n536 256.663
R1861 B.n877 B.n537 256.663
R1862 B.n877 B.n538 256.663
R1863 B.n877 B.n539 256.663
R1864 B.n877 B.n540 256.663
R1865 B.n877 B.n541 256.663
R1866 B.n877 B.n542 256.663
R1867 B.n877 B.n543 256.663
R1868 B.n877 B.n544 256.663
R1869 B.n877 B.n545 256.663
R1870 B.n877 B.n546 256.663
R1871 B.n877 B.n547 256.663
R1872 B.n877 B.n548 256.663
R1873 B.n877 B.n549 256.663
R1874 B.n877 B.n550 256.663
R1875 B.n877 B.n551 256.663
R1876 B.n877 B.n552 256.663
R1877 B.n877 B.n553 256.663
R1878 B.n877 B.n554 256.663
R1879 B.n877 B.n555 256.663
R1880 B.n877 B.n556 256.663
R1881 B.n877 B.n557 256.663
R1882 B.n877 B.n558 256.663
R1883 B.n877 B.n559 256.663
R1884 B.n877 B.n560 256.663
R1885 B.n877 B.n561 256.663
R1886 B.n877 B.n562 256.663
R1887 B.n877 B.n563 256.663
R1888 B.n877 B.n564 256.663
R1889 B.n877 B.n565 256.663
R1890 B.n877 B.n566 256.663
R1891 B.n877 B.n567 256.663
R1892 B.n877 B.n568 256.663
R1893 B.n877 B.n569 256.663
R1894 B.n877 B.n570 256.663
R1895 B.n877 B.n571 256.663
R1896 B.n877 B.n572 256.663
R1897 B.n877 B.n573 256.663
R1898 B.n877 B.n574 256.663
R1899 B.n877 B.n575 256.663
R1900 B.n877 B.n576 256.663
R1901 B.n877 B.n577 256.663
R1902 B.n877 B.n578 256.663
R1903 B.n877 B.n579 256.663
R1904 B.n877 B.n580 256.663
R1905 B.n877 B.n581 256.663
R1906 B.n877 B.n582 256.663
R1907 B.n877 B.n583 256.663
R1908 B.n877 B.n584 256.663
R1909 B.n877 B.n585 256.663
R1910 B.n877 B.n586 256.663
R1911 B.n877 B.n587 256.663
R1912 B.n877 B.n588 256.663
R1913 B.n877 B.n589 256.663
R1914 B.n877 B.n590 256.663
R1915 B.n877 B.n591 256.663
R1916 B.n877 B.n592 256.663
R1917 B.n877 B.n593 256.663
R1918 B.n877 B.n594 256.663
R1919 B.n877 B.n595 256.663
R1920 B.n877 B.n596 256.663
R1921 B.n877 B.n597 256.663
R1922 B.n877 B.n598 256.663
R1923 B.n877 B.n599 256.663
R1924 B.n878 B.n877 256.663
R1925 B.n1197 B.n1196 256.663
R1926 B.n170 B.n169 163.367
R1927 B.n174 B.n173 163.367
R1928 B.n178 B.n177 163.367
R1929 B.n182 B.n181 163.367
R1930 B.n186 B.n185 163.367
R1931 B.n190 B.n189 163.367
R1932 B.n194 B.n193 163.367
R1933 B.n198 B.n197 163.367
R1934 B.n202 B.n201 163.367
R1935 B.n206 B.n205 163.367
R1936 B.n210 B.n209 163.367
R1937 B.n214 B.n213 163.367
R1938 B.n218 B.n217 163.367
R1939 B.n222 B.n221 163.367
R1940 B.n226 B.n225 163.367
R1941 B.n230 B.n229 163.367
R1942 B.n234 B.n233 163.367
R1943 B.n238 B.n237 163.367
R1944 B.n242 B.n241 163.367
R1945 B.n246 B.n245 163.367
R1946 B.n250 B.n249 163.367
R1947 B.n254 B.n253 163.367
R1948 B.n258 B.n257 163.367
R1949 B.n262 B.n261 163.367
R1950 B.n266 B.n265 163.367
R1951 B.n270 B.n269 163.367
R1952 B.n274 B.n273 163.367
R1953 B.n278 B.n277 163.367
R1954 B.n282 B.n281 163.367
R1955 B.n286 B.n285 163.367
R1956 B.n290 B.n289 163.367
R1957 B.n294 B.n293 163.367
R1958 B.n298 B.n297 163.367
R1959 B.n302 B.n301 163.367
R1960 B.n306 B.n305 163.367
R1961 B.n310 B.n309 163.367
R1962 B.n315 B.n314 163.367
R1963 B.n319 B.n318 163.367
R1964 B.n323 B.n322 163.367
R1965 B.n327 B.n326 163.367
R1966 B.n331 B.n330 163.367
R1967 B.n335 B.n334 163.367
R1968 B.n339 B.n338 163.367
R1969 B.n343 B.n342 163.367
R1970 B.n347 B.n346 163.367
R1971 B.n351 B.n350 163.367
R1972 B.n355 B.n354 163.367
R1973 B.n359 B.n358 163.367
R1974 B.n363 B.n362 163.367
R1975 B.n367 B.n366 163.367
R1976 B.n371 B.n370 163.367
R1977 B.n375 B.n374 163.367
R1978 B.n379 B.n378 163.367
R1979 B.n383 B.n382 163.367
R1980 B.n387 B.n386 163.367
R1981 B.n391 B.n390 163.367
R1982 B.n395 B.n394 163.367
R1983 B.n399 B.n398 163.367
R1984 B.n403 B.n402 163.367
R1985 B.n407 B.n406 163.367
R1986 B.n411 B.n410 163.367
R1987 B.n415 B.n414 163.367
R1988 B.n419 B.n418 163.367
R1989 B.n423 B.n422 163.367
R1990 B.n427 B.n426 163.367
R1991 B.n431 B.n430 163.367
R1992 B.n435 B.n434 163.367
R1993 B.n1094 B.n160 163.367
R1994 B.n883 B.n531 163.367
R1995 B.n883 B.n525 163.367
R1996 B.n891 B.n525 163.367
R1997 B.n891 B.n523 163.367
R1998 B.n895 B.n523 163.367
R1999 B.n895 B.n516 163.367
R2000 B.n903 B.n516 163.367
R2001 B.n903 B.n514 163.367
R2002 B.n907 B.n514 163.367
R2003 B.n907 B.n509 163.367
R2004 B.n915 B.n509 163.367
R2005 B.n915 B.n507 163.367
R2006 B.n919 B.n507 163.367
R2007 B.n919 B.n501 163.367
R2008 B.n927 B.n501 163.367
R2009 B.n927 B.n499 163.367
R2010 B.n931 B.n499 163.367
R2011 B.n931 B.n493 163.367
R2012 B.n939 B.n493 163.367
R2013 B.n939 B.n491 163.367
R2014 B.n943 B.n491 163.367
R2015 B.n943 B.n486 163.367
R2016 B.n952 B.n486 163.367
R2017 B.n952 B.n484 163.367
R2018 B.n956 B.n484 163.367
R2019 B.n956 B.n478 163.367
R2020 B.n964 B.n478 163.367
R2021 B.n964 B.n476 163.367
R2022 B.n968 B.n476 163.367
R2023 B.n968 B.n469 163.367
R2024 B.n976 B.n469 163.367
R2025 B.n976 B.n467 163.367
R2026 B.n980 B.n467 163.367
R2027 B.n980 B.n462 163.367
R2028 B.n988 B.n462 163.367
R2029 B.n988 B.n460 163.367
R2030 B.n992 B.n460 163.367
R2031 B.n992 B.n454 163.367
R2032 B.n1000 B.n454 163.367
R2033 B.n1000 B.n452 163.367
R2034 B.n1004 B.n452 163.367
R2035 B.n1004 B.n447 163.367
R2036 B.n1013 B.n447 163.367
R2037 B.n1013 B.n445 163.367
R2038 B.n1018 B.n445 163.367
R2039 B.n1018 B.n439 163.367
R2040 B.n1026 B.n439 163.367
R2041 B.n1027 B.n1026 163.367
R2042 B.n1027 B.n5 163.367
R2043 B.n6 B.n5 163.367
R2044 B.n7 B.n6 163.367
R2045 B.n1033 B.n7 163.367
R2046 B.n1034 B.n1033 163.367
R2047 B.n1034 B.n13 163.367
R2048 B.n14 B.n13 163.367
R2049 B.n15 B.n14 163.367
R2050 B.n1039 B.n15 163.367
R2051 B.n1039 B.n20 163.367
R2052 B.n21 B.n20 163.367
R2053 B.n22 B.n21 163.367
R2054 B.n1044 B.n22 163.367
R2055 B.n1044 B.n27 163.367
R2056 B.n28 B.n27 163.367
R2057 B.n29 B.n28 163.367
R2058 B.n1049 B.n29 163.367
R2059 B.n1049 B.n34 163.367
R2060 B.n35 B.n34 163.367
R2061 B.n36 B.n35 163.367
R2062 B.n1054 B.n36 163.367
R2063 B.n1054 B.n41 163.367
R2064 B.n42 B.n41 163.367
R2065 B.n43 B.n42 163.367
R2066 B.n1059 B.n43 163.367
R2067 B.n1059 B.n48 163.367
R2068 B.n49 B.n48 163.367
R2069 B.n50 B.n49 163.367
R2070 B.n1064 B.n50 163.367
R2071 B.n1064 B.n55 163.367
R2072 B.n56 B.n55 163.367
R2073 B.n57 B.n56 163.367
R2074 B.n1069 B.n57 163.367
R2075 B.n1069 B.n62 163.367
R2076 B.n63 B.n62 163.367
R2077 B.n64 B.n63 163.367
R2078 B.n1074 B.n64 163.367
R2079 B.n1074 B.n69 163.367
R2080 B.n70 B.n69 163.367
R2081 B.n71 B.n70 163.367
R2082 B.n1079 B.n71 163.367
R2083 B.n1079 B.n76 163.367
R2084 B.n77 B.n76 163.367
R2085 B.n78 B.n77 163.367
R2086 B.n1084 B.n78 163.367
R2087 B.n1084 B.n83 163.367
R2088 B.n84 B.n83 163.367
R2089 B.n85 B.n84 163.367
R2090 B.n1089 B.n85 163.367
R2091 B.n1089 B.n90 163.367
R2092 B.n91 B.n90 163.367
R2093 B.n601 B.n600 163.367
R2094 B.n870 B.n600 163.367
R2095 B.n868 B.n867 163.367
R2096 B.n864 B.n863 163.367
R2097 B.n860 B.n859 163.367
R2098 B.n856 B.n855 163.367
R2099 B.n852 B.n851 163.367
R2100 B.n848 B.n847 163.367
R2101 B.n844 B.n843 163.367
R2102 B.n840 B.n839 163.367
R2103 B.n836 B.n835 163.367
R2104 B.n832 B.n831 163.367
R2105 B.n828 B.n827 163.367
R2106 B.n824 B.n823 163.367
R2107 B.n820 B.n819 163.367
R2108 B.n816 B.n815 163.367
R2109 B.n812 B.n811 163.367
R2110 B.n808 B.n807 163.367
R2111 B.n804 B.n803 163.367
R2112 B.n800 B.n799 163.367
R2113 B.n796 B.n795 163.367
R2114 B.n792 B.n791 163.367
R2115 B.n788 B.n787 163.367
R2116 B.n784 B.n783 163.367
R2117 B.n780 B.n779 163.367
R2118 B.n776 B.n775 163.367
R2119 B.n772 B.n771 163.367
R2120 B.n768 B.n767 163.367
R2121 B.n764 B.n763 163.367
R2122 B.n760 B.n759 163.367
R2123 B.n756 B.n755 163.367
R2124 B.n752 B.n751 163.367
R2125 B.n747 B.n746 163.367
R2126 B.n743 B.n742 163.367
R2127 B.n739 B.n738 163.367
R2128 B.n735 B.n734 163.367
R2129 B.n731 B.n730 163.367
R2130 B.n727 B.n726 163.367
R2131 B.n723 B.n722 163.367
R2132 B.n719 B.n718 163.367
R2133 B.n715 B.n714 163.367
R2134 B.n711 B.n710 163.367
R2135 B.n707 B.n706 163.367
R2136 B.n703 B.n702 163.367
R2137 B.n699 B.n698 163.367
R2138 B.n695 B.n694 163.367
R2139 B.n691 B.n690 163.367
R2140 B.n687 B.n686 163.367
R2141 B.n683 B.n682 163.367
R2142 B.n679 B.n678 163.367
R2143 B.n675 B.n674 163.367
R2144 B.n671 B.n670 163.367
R2145 B.n667 B.n666 163.367
R2146 B.n663 B.n662 163.367
R2147 B.n659 B.n658 163.367
R2148 B.n655 B.n654 163.367
R2149 B.n651 B.n650 163.367
R2150 B.n647 B.n646 163.367
R2151 B.n643 B.n642 163.367
R2152 B.n639 B.n638 163.367
R2153 B.n635 B.n634 163.367
R2154 B.n631 B.n630 163.367
R2155 B.n627 B.n626 163.367
R2156 B.n623 B.n622 163.367
R2157 B.n619 B.n618 163.367
R2158 B.n615 B.n614 163.367
R2159 B.n611 B.n610 163.367
R2160 B.n607 B.n533 163.367
R2161 B.n885 B.n529 163.367
R2162 B.n885 B.n527 163.367
R2163 B.n889 B.n527 163.367
R2164 B.n889 B.n521 163.367
R2165 B.n897 B.n521 163.367
R2166 B.n897 B.n519 163.367
R2167 B.n901 B.n519 163.367
R2168 B.n901 B.n513 163.367
R2169 B.n909 B.n513 163.367
R2170 B.n909 B.n511 163.367
R2171 B.n913 B.n511 163.367
R2172 B.n913 B.n505 163.367
R2173 B.n921 B.n505 163.367
R2174 B.n921 B.n503 163.367
R2175 B.n925 B.n503 163.367
R2176 B.n925 B.n497 163.367
R2177 B.n933 B.n497 163.367
R2178 B.n933 B.n495 163.367
R2179 B.n937 B.n495 163.367
R2180 B.n937 B.n489 163.367
R2181 B.n946 B.n489 163.367
R2182 B.n946 B.n487 163.367
R2183 B.n950 B.n487 163.367
R2184 B.n950 B.n482 163.367
R2185 B.n958 B.n482 163.367
R2186 B.n958 B.n480 163.367
R2187 B.n962 B.n480 163.367
R2188 B.n962 B.n474 163.367
R2189 B.n970 B.n474 163.367
R2190 B.n970 B.n472 163.367
R2191 B.n974 B.n472 163.367
R2192 B.n974 B.n466 163.367
R2193 B.n982 B.n466 163.367
R2194 B.n982 B.n464 163.367
R2195 B.n986 B.n464 163.367
R2196 B.n986 B.n458 163.367
R2197 B.n994 B.n458 163.367
R2198 B.n994 B.n456 163.367
R2199 B.n998 B.n456 163.367
R2200 B.n998 B.n450 163.367
R2201 B.n1007 B.n450 163.367
R2202 B.n1007 B.n448 163.367
R2203 B.n1011 B.n448 163.367
R2204 B.n1011 B.n443 163.367
R2205 B.n1020 B.n443 163.367
R2206 B.n1020 B.n441 163.367
R2207 B.n1024 B.n441 163.367
R2208 B.n1024 B.n3 163.367
R2209 B.n1195 B.n3 163.367
R2210 B.n1191 B.n2 163.367
R2211 B.n1191 B.n1190 163.367
R2212 B.n1190 B.n9 163.367
R2213 B.n1186 B.n9 163.367
R2214 B.n1186 B.n11 163.367
R2215 B.n1182 B.n11 163.367
R2216 B.n1182 B.n16 163.367
R2217 B.n1178 B.n16 163.367
R2218 B.n1178 B.n18 163.367
R2219 B.n1174 B.n18 163.367
R2220 B.n1174 B.n24 163.367
R2221 B.n1170 B.n24 163.367
R2222 B.n1170 B.n26 163.367
R2223 B.n1166 B.n26 163.367
R2224 B.n1166 B.n31 163.367
R2225 B.n1162 B.n31 163.367
R2226 B.n1162 B.n33 163.367
R2227 B.n1158 B.n33 163.367
R2228 B.n1158 B.n38 163.367
R2229 B.n1154 B.n38 163.367
R2230 B.n1154 B.n40 163.367
R2231 B.n1150 B.n40 163.367
R2232 B.n1150 B.n45 163.367
R2233 B.n1146 B.n45 163.367
R2234 B.n1146 B.n47 163.367
R2235 B.n1142 B.n47 163.367
R2236 B.n1142 B.n51 163.367
R2237 B.n1138 B.n51 163.367
R2238 B.n1138 B.n53 163.367
R2239 B.n1134 B.n53 163.367
R2240 B.n1134 B.n59 163.367
R2241 B.n1130 B.n59 163.367
R2242 B.n1130 B.n61 163.367
R2243 B.n1126 B.n61 163.367
R2244 B.n1126 B.n66 163.367
R2245 B.n1122 B.n66 163.367
R2246 B.n1122 B.n68 163.367
R2247 B.n1118 B.n68 163.367
R2248 B.n1118 B.n73 163.367
R2249 B.n1114 B.n73 163.367
R2250 B.n1114 B.n75 163.367
R2251 B.n1110 B.n75 163.367
R2252 B.n1110 B.n80 163.367
R2253 B.n1106 B.n80 163.367
R2254 B.n1106 B.n82 163.367
R2255 B.n1102 B.n82 163.367
R2256 B.n1102 B.n87 163.367
R2257 B.n1098 B.n87 163.367
R2258 B.n1098 B.n89 163.367
R2259 B.n166 B.n92 71.676
R2260 B.n170 B.n93 71.676
R2261 B.n174 B.n94 71.676
R2262 B.n178 B.n95 71.676
R2263 B.n182 B.n96 71.676
R2264 B.n186 B.n97 71.676
R2265 B.n190 B.n98 71.676
R2266 B.n194 B.n99 71.676
R2267 B.n198 B.n100 71.676
R2268 B.n202 B.n101 71.676
R2269 B.n206 B.n102 71.676
R2270 B.n210 B.n103 71.676
R2271 B.n214 B.n104 71.676
R2272 B.n218 B.n105 71.676
R2273 B.n222 B.n106 71.676
R2274 B.n226 B.n107 71.676
R2275 B.n230 B.n108 71.676
R2276 B.n234 B.n109 71.676
R2277 B.n238 B.n110 71.676
R2278 B.n242 B.n111 71.676
R2279 B.n246 B.n112 71.676
R2280 B.n250 B.n113 71.676
R2281 B.n254 B.n114 71.676
R2282 B.n258 B.n115 71.676
R2283 B.n262 B.n116 71.676
R2284 B.n266 B.n117 71.676
R2285 B.n270 B.n118 71.676
R2286 B.n274 B.n119 71.676
R2287 B.n278 B.n120 71.676
R2288 B.n282 B.n121 71.676
R2289 B.n286 B.n122 71.676
R2290 B.n290 B.n123 71.676
R2291 B.n294 B.n124 71.676
R2292 B.n298 B.n125 71.676
R2293 B.n302 B.n126 71.676
R2294 B.n306 B.n127 71.676
R2295 B.n310 B.n128 71.676
R2296 B.n315 B.n129 71.676
R2297 B.n319 B.n130 71.676
R2298 B.n323 B.n131 71.676
R2299 B.n327 B.n132 71.676
R2300 B.n331 B.n133 71.676
R2301 B.n335 B.n134 71.676
R2302 B.n339 B.n135 71.676
R2303 B.n343 B.n136 71.676
R2304 B.n347 B.n137 71.676
R2305 B.n351 B.n138 71.676
R2306 B.n355 B.n139 71.676
R2307 B.n359 B.n140 71.676
R2308 B.n363 B.n141 71.676
R2309 B.n367 B.n142 71.676
R2310 B.n371 B.n143 71.676
R2311 B.n375 B.n144 71.676
R2312 B.n379 B.n145 71.676
R2313 B.n383 B.n146 71.676
R2314 B.n387 B.n147 71.676
R2315 B.n391 B.n148 71.676
R2316 B.n395 B.n149 71.676
R2317 B.n399 B.n150 71.676
R2318 B.n403 B.n151 71.676
R2319 B.n407 B.n152 71.676
R2320 B.n411 B.n153 71.676
R2321 B.n415 B.n154 71.676
R2322 B.n419 B.n155 71.676
R2323 B.n423 B.n156 71.676
R2324 B.n427 B.n157 71.676
R2325 B.n431 B.n158 71.676
R2326 B.n435 B.n159 71.676
R2327 B.n160 B.n159 71.676
R2328 B.n434 B.n158 71.676
R2329 B.n430 B.n157 71.676
R2330 B.n426 B.n156 71.676
R2331 B.n422 B.n155 71.676
R2332 B.n418 B.n154 71.676
R2333 B.n414 B.n153 71.676
R2334 B.n410 B.n152 71.676
R2335 B.n406 B.n151 71.676
R2336 B.n402 B.n150 71.676
R2337 B.n398 B.n149 71.676
R2338 B.n394 B.n148 71.676
R2339 B.n390 B.n147 71.676
R2340 B.n386 B.n146 71.676
R2341 B.n382 B.n145 71.676
R2342 B.n378 B.n144 71.676
R2343 B.n374 B.n143 71.676
R2344 B.n370 B.n142 71.676
R2345 B.n366 B.n141 71.676
R2346 B.n362 B.n140 71.676
R2347 B.n358 B.n139 71.676
R2348 B.n354 B.n138 71.676
R2349 B.n350 B.n137 71.676
R2350 B.n346 B.n136 71.676
R2351 B.n342 B.n135 71.676
R2352 B.n338 B.n134 71.676
R2353 B.n334 B.n133 71.676
R2354 B.n330 B.n132 71.676
R2355 B.n326 B.n131 71.676
R2356 B.n322 B.n130 71.676
R2357 B.n318 B.n129 71.676
R2358 B.n314 B.n128 71.676
R2359 B.n309 B.n127 71.676
R2360 B.n305 B.n126 71.676
R2361 B.n301 B.n125 71.676
R2362 B.n297 B.n124 71.676
R2363 B.n293 B.n123 71.676
R2364 B.n289 B.n122 71.676
R2365 B.n285 B.n121 71.676
R2366 B.n281 B.n120 71.676
R2367 B.n277 B.n119 71.676
R2368 B.n273 B.n118 71.676
R2369 B.n269 B.n117 71.676
R2370 B.n265 B.n116 71.676
R2371 B.n261 B.n115 71.676
R2372 B.n257 B.n114 71.676
R2373 B.n253 B.n113 71.676
R2374 B.n249 B.n112 71.676
R2375 B.n245 B.n111 71.676
R2376 B.n241 B.n110 71.676
R2377 B.n237 B.n109 71.676
R2378 B.n233 B.n108 71.676
R2379 B.n229 B.n107 71.676
R2380 B.n225 B.n106 71.676
R2381 B.n221 B.n105 71.676
R2382 B.n217 B.n104 71.676
R2383 B.n213 B.n103 71.676
R2384 B.n209 B.n102 71.676
R2385 B.n205 B.n101 71.676
R2386 B.n201 B.n100 71.676
R2387 B.n197 B.n99 71.676
R2388 B.n193 B.n98 71.676
R2389 B.n189 B.n97 71.676
R2390 B.n185 B.n96 71.676
R2391 B.n181 B.n95 71.676
R2392 B.n177 B.n94 71.676
R2393 B.n173 B.n93 71.676
R2394 B.n169 B.n92 71.676
R2395 B.n876 B.n875 71.676
R2396 B.n870 B.n534 71.676
R2397 B.n867 B.n535 71.676
R2398 B.n863 B.n536 71.676
R2399 B.n859 B.n537 71.676
R2400 B.n855 B.n538 71.676
R2401 B.n851 B.n539 71.676
R2402 B.n847 B.n540 71.676
R2403 B.n843 B.n541 71.676
R2404 B.n839 B.n542 71.676
R2405 B.n835 B.n543 71.676
R2406 B.n831 B.n544 71.676
R2407 B.n827 B.n545 71.676
R2408 B.n823 B.n546 71.676
R2409 B.n819 B.n547 71.676
R2410 B.n815 B.n548 71.676
R2411 B.n811 B.n549 71.676
R2412 B.n807 B.n550 71.676
R2413 B.n803 B.n551 71.676
R2414 B.n799 B.n552 71.676
R2415 B.n795 B.n553 71.676
R2416 B.n791 B.n554 71.676
R2417 B.n787 B.n555 71.676
R2418 B.n783 B.n556 71.676
R2419 B.n779 B.n557 71.676
R2420 B.n775 B.n558 71.676
R2421 B.n771 B.n559 71.676
R2422 B.n767 B.n560 71.676
R2423 B.n763 B.n561 71.676
R2424 B.n759 B.n562 71.676
R2425 B.n755 B.n563 71.676
R2426 B.n751 B.n564 71.676
R2427 B.n746 B.n565 71.676
R2428 B.n742 B.n566 71.676
R2429 B.n738 B.n567 71.676
R2430 B.n734 B.n568 71.676
R2431 B.n730 B.n569 71.676
R2432 B.n726 B.n570 71.676
R2433 B.n722 B.n571 71.676
R2434 B.n718 B.n572 71.676
R2435 B.n714 B.n573 71.676
R2436 B.n710 B.n574 71.676
R2437 B.n706 B.n575 71.676
R2438 B.n702 B.n576 71.676
R2439 B.n698 B.n577 71.676
R2440 B.n694 B.n578 71.676
R2441 B.n690 B.n579 71.676
R2442 B.n686 B.n580 71.676
R2443 B.n682 B.n581 71.676
R2444 B.n678 B.n582 71.676
R2445 B.n674 B.n583 71.676
R2446 B.n670 B.n584 71.676
R2447 B.n666 B.n585 71.676
R2448 B.n662 B.n586 71.676
R2449 B.n658 B.n587 71.676
R2450 B.n654 B.n588 71.676
R2451 B.n650 B.n589 71.676
R2452 B.n646 B.n590 71.676
R2453 B.n642 B.n591 71.676
R2454 B.n638 B.n592 71.676
R2455 B.n634 B.n593 71.676
R2456 B.n630 B.n594 71.676
R2457 B.n626 B.n595 71.676
R2458 B.n622 B.n596 71.676
R2459 B.n618 B.n597 71.676
R2460 B.n614 B.n598 71.676
R2461 B.n610 B.n599 71.676
R2462 B.n878 B.n533 71.676
R2463 B.n876 B.n601 71.676
R2464 B.n868 B.n534 71.676
R2465 B.n864 B.n535 71.676
R2466 B.n860 B.n536 71.676
R2467 B.n856 B.n537 71.676
R2468 B.n852 B.n538 71.676
R2469 B.n848 B.n539 71.676
R2470 B.n844 B.n540 71.676
R2471 B.n840 B.n541 71.676
R2472 B.n836 B.n542 71.676
R2473 B.n832 B.n543 71.676
R2474 B.n828 B.n544 71.676
R2475 B.n824 B.n545 71.676
R2476 B.n820 B.n546 71.676
R2477 B.n816 B.n547 71.676
R2478 B.n812 B.n548 71.676
R2479 B.n808 B.n549 71.676
R2480 B.n804 B.n550 71.676
R2481 B.n800 B.n551 71.676
R2482 B.n796 B.n552 71.676
R2483 B.n792 B.n553 71.676
R2484 B.n788 B.n554 71.676
R2485 B.n784 B.n555 71.676
R2486 B.n780 B.n556 71.676
R2487 B.n776 B.n557 71.676
R2488 B.n772 B.n558 71.676
R2489 B.n768 B.n559 71.676
R2490 B.n764 B.n560 71.676
R2491 B.n760 B.n561 71.676
R2492 B.n756 B.n562 71.676
R2493 B.n752 B.n563 71.676
R2494 B.n747 B.n564 71.676
R2495 B.n743 B.n565 71.676
R2496 B.n739 B.n566 71.676
R2497 B.n735 B.n567 71.676
R2498 B.n731 B.n568 71.676
R2499 B.n727 B.n569 71.676
R2500 B.n723 B.n570 71.676
R2501 B.n719 B.n571 71.676
R2502 B.n715 B.n572 71.676
R2503 B.n711 B.n573 71.676
R2504 B.n707 B.n574 71.676
R2505 B.n703 B.n575 71.676
R2506 B.n699 B.n576 71.676
R2507 B.n695 B.n577 71.676
R2508 B.n691 B.n578 71.676
R2509 B.n687 B.n579 71.676
R2510 B.n683 B.n580 71.676
R2511 B.n679 B.n581 71.676
R2512 B.n675 B.n582 71.676
R2513 B.n671 B.n583 71.676
R2514 B.n667 B.n584 71.676
R2515 B.n663 B.n585 71.676
R2516 B.n659 B.n586 71.676
R2517 B.n655 B.n587 71.676
R2518 B.n651 B.n588 71.676
R2519 B.n647 B.n589 71.676
R2520 B.n643 B.n590 71.676
R2521 B.n639 B.n591 71.676
R2522 B.n635 B.n592 71.676
R2523 B.n631 B.n593 71.676
R2524 B.n627 B.n594 71.676
R2525 B.n623 B.n595 71.676
R2526 B.n619 B.n596 71.676
R2527 B.n615 B.n597 71.676
R2528 B.n611 B.n598 71.676
R2529 B.n607 B.n599 71.676
R2530 B.n879 B.n878 71.676
R2531 B.n1196 B.n1195 71.676
R2532 B.n1196 B.n2 71.676
R2533 B.n164 B.n163 68.0732
R2534 B.n162 B.n161 68.0732
R2535 B.n605 B.n604 68.0732
R2536 B.n603 B.n602 68.0732
R2537 B.n165 B.n164 59.5399
R2538 B.n312 B.n162 59.5399
R2539 B.n606 B.n605 59.5399
R2540 B.n749 B.n603 59.5399
R2541 B.n877 B.n530 51.76
R2542 B.n1096 B.n1095 51.76
R2543 B.n874 B.n528 33.8737
R2544 B.n881 B.n880 33.8737
R2545 B.n1093 B.n1092 33.8737
R2546 B.n167 B.n88 33.8737
R2547 B.n884 B.n530 30.0829
R2548 B.n884 B.n526 30.0829
R2549 B.n890 B.n526 30.0829
R2550 B.n890 B.n522 30.0829
R2551 B.n896 B.n522 30.0829
R2552 B.n896 B.n517 30.0829
R2553 B.n902 B.n517 30.0829
R2554 B.n902 B.n518 30.0829
R2555 B.n908 B.n510 30.0829
R2556 B.n914 B.n510 30.0829
R2557 B.n914 B.n506 30.0829
R2558 B.n920 B.n506 30.0829
R2559 B.n920 B.n502 30.0829
R2560 B.n926 B.n502 30.0829
R2561 B.n926 B.n498 30.0829
R2562 B.n932 B.n498 30.0829
R2563 B.n932 B.n494 30.0829
R2564 B.n938 B.n494 30.0829
R2565 B.n938 B.n490 30.0829
R2566 B.n945 B.n490 30.0829
R2567 B.n945 B.n944 30.0829
R2568 B.n951 B.n483 30.0829
R2569 B.n957 B.n483 30.0829
R2570 B.n957 B.n479 30.0829
R2571 B.n963 B.n479 30.0829
R2572 B.n963 B.n475 30.0829
R2573 B.n969 B.n475 30.0829
R2574 B.n969 B.n470 30.0829
R2575 B.n975 B.n470 30.0829
R2576 B.n975 B.n471 30.0829
R2577 B.n981 B.n463 30.0829
R2578 B.n987 B.n463 30.0829
R2579 B.n987 B.n459 30.0829
R2580 B.n993 B.n459 30.0829
R2581 B.n993 B.n455 30.0829
R2582 B.n999 B.n455 30.0829
R2583 B.n999 B.n451 30.0829
R2584 B.n1006 B.n451 30.0829
R2585 B.n1006 B.n1005 30.0829
R2586 B.n1012 B.n444 30.0829
R2587 B.n1019 B.n444 30.0829
R2588 B.n1019 B.n440 30.0829
R2589 B.n1025 B.n440 30.0829
R2590 B.n1025 B.n4 30.0829
R2591 B.n1194 B.n4 30.0829
R2592 B.n1194 B.n1193 30.0829
R2593 B.n1193 B.n1192 30.0829
R2594 B.n1192 B.n8 30.0829
R2595 B.n12 B.n8 30.0829
R2596 B.n1185 B.n12 30.0829
R2597 B.n1185 B.n1184 30.0829
R2598 B.n1184 B.n1183 30.0829
R2599 B.n1177 B.n19 30.0829
R2600 B.n1177 B.n1176 30.0829
R2601 B.n1176 B.n1175 30.0829
R2602 B.n1175 B.n23 30.0829
R2603 B.n1169 B.n23 30.0829
R2604 B.n1169 B.n1168 30.0829
R2605 B.n1168 B.n1167 30.0829
R2606 B.n1167 B.n30 30.0829
R2607 B.n1161 B.n30 30.0829
R2608 B.n1160 B.n1159 30.0829
R2609 B.n1159 B.n37 30.0829
R2610 B.n1153 B.n37 30.0829
R2611 B.n1153 B.n1152 30.0829
R2612 B.n1152 B.n1151 30.0829
R2613 B.n1151 B.n44 30.0829
R2614 B.n1145 B.n44 30.0829
R2615 B.n1145 B.n1144 30.0829
R2616 B.n1144 B.n1143 30.0829
R2617 B.n1137 B.n54 30.0829
R2618 B.n1137 B.n1136 30.0829
R2619 B.n1136 B.n1135 30.0829
R2620 B.n1135 B.n58 30.0829
R2621 B.n1129 B.n58 30.0829
R2622 B.n1129 B.n1128 30.0829
R2623 B.n1128 B.n1127 30.0829
R2624 B.n1127 B.n65 30.0829
R2625 B.n1121 B.n65 30.0829
R2626 B.n1121 B.n1120 30.0829
R2627 B.n1120 B.n1119 30.0829
R2628 B.n1119 B.n72 30.0829
R2629 B.n1113 B.n72 30.0829
R2630 B.n1112 B.n1111 30.0829
R2631 B.n1111 B.n79 30.0829
R2632 B.n1105 B.n79 30.0829
R2633 B.n1105 B.n1104 30.0829
R2634 B.n1104 B.n1103 30.0829
R2635 B.n1103 B.n86 30.0829
R2636 B.n1097 B.n86 30.0829
R2637 B.n1097 B.n1096 30.0829
R2638 B.n951 B.t1 27.4286
R2639 B.n1143 B.t3 27.4286
R2640 B.n1005 B.t2 22.1199
R2641 B.n19 B.t4 22.1199
R2642 B B.n1197 18.0485
R2643 B.n981 B.t5 17.6961
R2644 B.n1161 B.t0 17.6961
R2645 B.n518 B.t11 16.8113
R2646 B.t7 B.n1112 16.8113
R2647 B.n908 B.t11 13.2722
R2648 B.n1113 B.t7 13.2722
R2649 B.n471 B.t5 12.3874
R2650 B.t0 B.n1160 12.3874
R2651 B.n886 B.n528 10.6151
R2652 B.n887 B.n886 10.6151
R2653 B.n888 B.n887 10.6151
R2654 B.n888 B.n520 10.6151
R2655 B.n898 B.n520 10.6151
R2656 B.n899 B.n898 10.6151
R2657 B.n900 B.n899 10.6151
R2658 B.n900 B.n512 10.6151
R2659 B.n910 B.n512 10.6151
R2660 B.n911 B.n910 10.6151
R2661 B.n912 B.n911 10.6151
R2662 B.n912 B.n504 10.6151
R2663 B.n922 B.n504 10.6151
R2664 B.n923 B.n922 10.6151
R2665 B.n924 B.n923 10.6151
R2666 B.n924 B.n496 10.6151
R2667 B.n934 B.n496 10.6151
R2668 B.n935 B.n934 10.6151
R2669 B.n936 B.n935 10.6151
R2670 B.n936 B.n488 10.6151
R2671 B.n947 B.n488 10.6151
R2672 B.n948 B.n947 10.6151
R2673 B.n949 B.n948 10.6151
R2674 B.n949 B.n481 10.6151
R2675 B.n959 B.n481 10.6151
R2676 B.n960 B.n959 10.6151
R2677 B.n961 B.n960 10.6151
R2678 B.n961 B.n473 10.6151
R2679 B.n971 B.n473 10.6151
R2680 B.n972 B.n971 10.6151
R2681 B.n973 B.n972 10.6151
R2682 B.n973 B.n465 10.6151
R2683 B.n983 B.n465 10.6151
R2684 B.n984 B.n983 10.6151
R2685 B.n985 B.n984 10.6151
R2686 B.n985 B.n457 10.6151
R2687 B.n995 B.n457 10.6151
R2688 B.n996 B.n995 10.6151
R2689 B.n997 B.n996 10.6151
R2690 B.n997 B.n449 10.6151
R2691 B.n1008 B.n449 10.6151
R2692 B.n1009 B.n1008 10.6151
R2693 B.n1010 B.n1009 10.6151
R2694 B.n1010 B.n442 10.6151
R2695 B.n1021 B.n442 10.6151
R2696 B.n1022 B.n1021 10.6151
R2697 B.n1023 B.n1022 10.6151
R2698 B.n1023 B.n0 10.6151
R2699 B.n874 B.n873 10.6151
R2700 B.n873 B.n872 10.6151
R2701 B.n872 B.n871 10.6151
R2702 B.n871 B.n869 10.6151
R2703 B.n869 B.n866 10.6151
R2704 B.n866 B.n865 10.6151
R2705 B.n865 B.n862 10.6151
R2706 B.n862 B.n861 10.6151
R2707 B.n861 B.n858 10.6151
R2708 B.n858 B.n857 10.6151
R2709 B.n857 B.n854 10.6151
R2710 B.n854 B.n853 10.6151
R2711 B.n853 B.n850 10.6151
R2712 B.n850 B.n849 10.6151
R2713 B.n849 B.n846 10.6151
R2714 B.n846 B.n845 10.6151
R2715 B.n845 B.n842 10.6151
R2716 B.n842 B.n841 10.6151
R2717 B.n841 B.n838 10.6151
R2718 B.n838 B.n837 10.6151
R2719 B.n837 B.n834 10.6151
R2720 B.n834 B.n833 10.6151
R2721 B.n833 B.n830 10.6151
R2722 B.n830 B.n829 10.6151
R2723 B.n829 B.n826 10.6151
R2724 B.n826 B.n825 10.6151
R2725 B.n825 B.n822 10.6151
R2726 B.n822 B.n821 10.6151
R2727 B.n821 B.n818 10.6151
R2728 B.n818 B.n817 10.6151
R2729 B.n817 B.n814 10.6151
R2730 B.n814 B.n813 10.6151
R2731 B.n813 B.n810 10.6151
R2732 B.n810 B.n809 10.6151
R2733 B.n809 B.n806 10.6151
R2734 B.n806 B.n805 10.6151
R2735 B.n805 B.n802 10.6151
R2736 B.n802 B.n801 10.6151
R2737 B.n801 B.n798 10.6151
R2738 B.n798 B.n797 10.6151
R2739 B.n797 B.n794 10.6151
R2740 B.n794 B.n793 10.6151
R2741 B.n793 B.n790 10.6151
R2742 B.n790 B.n789 10.6151
R2743 B.n789 B.n786 10.6151
R2744 B.n786 B.n785 10.6151
R2745 B.n785 B.n782 10.6151
R2746 B.n782 B.n781 10.6151
R2747 B.n781 B.n778 10.6151
R2748 B.n778 B.n777 10.6151
R2749 B.n777 B.n774 10.6151
R2750 B.n774 B.n773 10.6151
R2751 B.n773 B.n770 10.6151
R2752 B.n770 B.n769 10.6151
R2753 B.n769 B.n766 10.6151
R2754 B.n766 B.n765 10.6151
R2755 B.n765 B.n762 10.6151
R2756 B.n762 B.n761 10.6151
R2757 B.n761 B.n758 10.6151
R2758 B.n758 B.n757 10.6151
R2759 B.n757 B.n754 10.6151
R2760 B.n754 B.n753 10.6151
R2761 B.n753 B.n750 10.6151
R2762 B.n748 B.n745 10.6151
R2763 B.n745 B.n744 10.6151
R2764 B.n744 B.n741 10.6151
R2765 B.n741 B.n740 10.6151
R2766 B.n740 B.n737 10.6151
R2767 B.n737 B.n736 10.6151
R2768 B.n736 B.n733 10.6151
R2769 B.n733 B.n732 10.6151
R2770 B.n729 B.n728 10.6151
R2771 B.n728 B.n725 10.6151
R2772 B.n725 B.n724 10.6151
R2773 B.n724 B.n721 10.6151
R2774 B.n721 B.n720 10.6151
R2775 B.n720 B.n717 10.6151
R2776 B.n717 B.n716 10.6151
R2777 B.n716 B.n713 10.6151
R2778 B.n713 B.n712 10.6151
R2779 B.n712 B.n709 10.6151
R2780 B.n709 B.n708 10.6151
R2781 B.n708 B.n705 10.6151
R2782 B.n705 B.n704 10.6151
R2783 B.n704 B.n701 10.6151
R2784 B.n701 B.n700 10.6151
R2785 B.n700 B.n697 10.6151
R2786 B.n697 B.n696 10.6151
R2787 B.n696 B.n693 10.6151
R2788 B.n693 B.n692 10.6151
R2789 B.n692 B.n689 10.6151
R2790 B.n689 B.n688 10.6151
R2791 B.n688 B.n685 10.6151
R2792 B.n685 B.n684 10.6151
R2793 B.n684 B.n681 10.6151
R2794 B.n681 B.n680 10.6151
R2795 B.n680 B.n677 10.6151
R2796 B.n677 B.n676 10.6151
R2797 B.n676 B.n673 10.6151
R2798 B.n673 B.n672 10.6151
R2799 B.n672 B.n669 10.6151
R2800 B.n669 B.n668 10.6151
R2801 B.n668 B.n665 10.6151
R2802 B.n665 B.n664 10.6151
R2803 B.n664 B.n661 10.6151
R2804 B.n661 B.n660 10.6151
R2805 B.n660 B.n657 10.6151
R2806 B.n657 B.n656 10.6151
R2807 B.n656 B.n653 10.6151
R2808 B.n653 B.n652 10.6151
R2809 B.n652 B.n649 10.6151
R2810 B.n649 B.n648 10.6151
R2811 B.n648 B.n645 10.6151
R2812 B.n645 B.n644 10.6151
R2813 B.n644 B.n641 10.6151
R2814 B.n641 B.n640 10.6151
R2815 B.n640 B.n637 10.6151
R2816 B.n637 B.n636 10.6151
R2817 B.n636 B.n633 10.6151
R2818 B.n633 B.n632 10.6151
R2819 B.n632 B.n629 10.6151
R2820 B.n629 B.n628 10.6151
R2821 B.n628 B.n625 10.6151
R2822 B.n625 B.n624 10.6151
R2823 B.n624 B.n621 10.6151
R2824 B.n621 B.n620 10.6151
R2825 B.n620 B.n617 10.6151
R2826 B.n617 B.n616 10.6151
R2827 B.n616 B.n613 10.6151
R2828 B.n613 B.n612 10.6151
R2829 B.n612 B.n609 10.6151
R2830 B.n609 B.n608 10.6151
R2831 B.n608 B.n532 10.6151
R2832 B.n880 B.n532 10.6151
R2833 B.n882 B.n881 10.6151
R2834 B.n882 B.n524 10.6151
R2835 B.n892 B.n524 10.6151
R2836 B.n893 B.n892 10.6151
R2837 B.n894 B.n893 10.6151
R2838 B.n894 B.n515 10.6151
R2839 B.n904 B.n515 10.6151
R2840 B.n905 B.n904 10.6151
R2841 B.n906 B.n905 10.6151
R2842 B.n906 B.n508 10.6151
R2843 B.n916 B.n508 10.6151
R2844 B.n917 B.n916 10.6151
R2845 B.n918 B.n917 10.6151
R2846 B.n918 B.n500 10.6151
R2847 B.n928 B.n500 10.6151
R2848 B.n929 B.n928 10.6151
R2849 B.n930 B.n929 10.6151
R2850 B.n930 B.n492 10.6151
R2851 B.n940 B.n492 10.6151
R2852 B.n941 B.n940 10.6151
R2853 B.n942 B.n941 10.6151
R2854 B.n942 B.n485 10.6151
R2855 B.n953 B.n485 10.6151
R2856 B.n954 B.n953 10.6151
R2857 B.n955 B.n954 10.6151
R2858 B.n955 B.n477 10.6151
R2859 B.n965 B.n477 10.6151
R2860 B.n966 B.n965 10.6151
R2861 B.n967 B.n966 10.6151
R2862 B.n967 B.n468 10.6151
R2863 B.n977 B.n468 10.6151
R2864 B.n978 B.n977 10.6151
R2865 B.n979 B.n978 10.6151
R2866 B.n979 B.n461 10.6151
R2867 B.n989 B.n461 10.6151
R2868 B.n990 B.n989 10.6151
R2869 B.n991 B.n990 10.6151
R2870 B.n991 B.n453 10.6151
R2871 B.n1001 B.n453 10.6151
R2872 B.n1002 B.n1001 10.6151
R2873 B.n1003 B.n1002 10.6151
R2874 B.n1003 B.n446 10.6151
R2875 B.n1014 B.n446 10.6151
R2876 B.n1015 B.n1014 10.6151
R2877 B.n1017 B.n1015 10.6151
R2878 B.n1017 B.n1016 10.6151
R2879 B.n1016 B.n438 10.6151
R2880 B.n1028 B.n438 10.6151
R2881 B.n1029 B.n1028 10.6151
R2882 B.n1030 B.n1029 10.6151
R2883 B.n1031 B.n1030 10.6151
R2884 B.n1032 B.n1031 10.6151
R2885 B.n1035 B.n1032 10.6151
R2886 B.n1036 B.n1035 10.6151
R2887 B.n1037 B.n1036 10.6151
R2888 B.n1038 B.n1037 10.6151
R2889 B.n1040 B.n1038 10.6151
R2890 B.n1041 B.n1040 10.6151
R2891 B.n1042 B.n1041 10.6151
R2892 B.n1043 B.n1042 10.6151
R2893 B.n1045 B.n1043 10.6151
R2894 B.n1046 B.n1045 10.6151
R2895 B.n1047 B.n1046 10.6151
R2896 B.n1048 B.n1047 10.6151
R2897 B.n1050 B.n1048 10.6151
R2898 B.n1051 B.n1050 10.6151
R2899 B.n1052 B.n1051 10.6151
R2900 B.n1053 B.n1052 10.6151
R2901 B.n1055 B.n1053 10.6151
R2902 B.n1056 B.n1055 10.6151
R2903 B.n1057 B.n1056 10.6151
R2904 B.n1058 B.n1057 10.6151
R2905 B.n1060 B.n1058 10.6151
R2906 B.n1061 B.n1060 10.6151
R2907 B.n1062 B.n1061 10.6151
R2908 B.n1063 B.n1062 10.6151
R2909 B.n1065 B.n1063 10.6151
R2910 B.n1066 B.n1065 10.6151
R2911 B.n1067 B.n1066 10.6151
R2912 B.n1068 B.n1067 10.6151
R2913 B.n1070 B.n1068 10.6151
R2914 B.n1071 B.n1070 10.6151
R2915 B.n1072 B.n1071 10.6151
R2916 B.n1073 B.n1072 10.6151
R2917 B.n1075 B.n1073 10.6151
R2918 B.n1076 B.n1075 10.6151
R2919 B.n1077 B.n1076 10.6151
R2920 B.n1078 B.n1077 10.6151
R2921 B.n1080 B.n1078 10.6151
R2922 B.n1081 B.n1080 10.6151
R2923 B.n1082 B.n1081 10.6151
R2924 B.n1083 B.n1082 10.6151
R2925 B.n1085 B.n1083 10.6151
R2926 B.n1086 B.n1085 10.6151
R2927 B.n1087 B.n1086 10.6151
R2928 B.n1088 B.n1087 10.6151
R2929 B.n1090 B.n1088 10.6151
R2930 B.n1091 B.n1090 10.6151
R2931 B.n1092 B.n1091 10.6151
R2932 B.n1189 B.n1 10.6151
R2933 B.n1189 B.n1188 10.6151
R2934 B.n1188 B.n1187 10.6151
R2935 B.n1187 B.n10 10.6151
R2936 B.n1181 B.n10 10.6151
R2937 B.n1181 B.n1180 10.6151
R2938 B.n1180 B.n1179 10.6151
R2939 B.n1179 B.n17 10.6151
R2940 B.n1173 B.n17 10.6151
R2941 B.n1173 B.n1172 10.6151
R2942 B.n1172 B.n1171 10.6151
R2943 B.n1171 B.n25 10.6151
R2944 B.n1165 B.n25 10.6151
R2945 B.n1165 B.n1164 10.6151
R2946 B.n1164 B.n1163 10.6151
R2947 B.n1163 B.n32 10.6151
R2948 B.n1157 B.n32 10.6151
R2949 B.n1157 B.n1156 10.6151
R2950 B.n1156 B.n1155 10.6151
R2951 B.n1155 B.n39 10.6151
R2952 B.n1149 B.n39 10.6151
R2953 B.n1149 B.n1148 10.6151
R2954 B.n1148 B.n1147 10.6151
R2955 B.n1147 B.n46 10.6151
R2956 B.n1141 B.n46 10.6151
R2957 B.n1141 B.n1140 10.6151
R2958 B.n1140 B.n1139 10.6151
R2959 B.n1139 B.n52 10.6151
R2960 B.n1133 B.n52 10.6151
R2961 B.n1133 B.n1132 10.6151
R2962 B.n1132 B.n1131 10.6151
R2963 B.n1131 B.n60 10.6151
R2964 B.n1125 B.n60 10.6151
R2965 B.n1125 B.n1124 10.6151
R2966 B.n1124 B.n1123 10.6151
R2967 B.n1123 B.n67 10.6151
R2968 B.n1117 B.n67 10.6151
R2969 B.n1117 B.n1116 10.6151
R2970 B.n1116 B.n1115 10.6151
R2971 B.n1115 B.n74 10.6151
R2972 B.n1109 B.n74 10.6151
R2973 B.n1109 B.n1108 10.6151
R2974 B.n1108 B.n1107 10.6151
R2975 B.n1107 B.n81 10.6151
R2976 B.n1101 B.n81 10.6151
R2977 B.n1101 B.n1100 10.6151
R2978 B.n1100 B.n1099 10.6151
R2979 B.n1099 B.n88 10.6151
R2980 B.n168 B.n167 10.6151
R2981 B.n171 B.n168 10.6151
R2982 B.n172 B.n171 10.6151
R2983 B.n175 B.n172 10.6151
R2984 B.n176 B.n175 10.6151
R2985 B.n179 B.n176 10.6151
R2986 B.n180 B.n179 10.6151
R2987 B.n183 B.n180 10.6151
R2988 B.n184 B.n183 10.6151
R2989 B.n187 B.n184 10.6151
R2990 B.n188 B.n187 10.6151
R2991 B.n191 B.n188 10.6151
R2992 B.n192 B.n191 10.6151
R2993 B.n195 B.n192 10.6151
R2994 B.n196 B.n195 10.6151
R2995 B.n199 B.n196 10.6151
R2996 B.n200 B.n199 10.6151
R2997 B.n203 B.n200 10.6151
R2998 B.n204 B.n203 10.6151
R2999 B.n207 B.n204 10.6151
R3000 B.n208 B.n207 10.6151
R3001 B.n211 B.n208 10.6151
R3002 B.n212 B.n211 10.6151
R3003 B.n215 B.n212 10.6151
R3004 B.n216 B.n215 10.6151
R3005 B.n219 B.n216 10.6151
R3006 B.n220 B.n219 10.6151
R3007 B.n223 B.n220 10.6151
R3008 B.n224 B.n223 10.6151
R3009 B.n227 B.n224 10.6151
R3010 B.n228 B.n227 10.6151
R3011 B.n231 B.n228 10.6151
R3012 B.n232 B.n231 10.6151
R3013 B.n235 B.n232 10.6151
R3014 B.n236 B.n235 10.6151
R3015 B.n239 B.n236 10.6151
R3016 B.n240 B.n239 10.6151
R3017 B.n243 B.n240 10.6151
R3018 B.n244 B.n243 10.6151
R3019 B.n247 B.n244 10.6151
R3020 B.n248 B.n247 10.6151
R3021 B.n251 B.n248 10.6151
R3022 B.n252 B.n251 10.6151
R3023 B.n255 B.n252 10.6151
R3024 B.n256 B.n255 10.6151
R3025 B.n259 B.n256 10.6151
R3026 B.n260 B.n259 10.6151
R3027 B.n263 B.n260 10.6151
R3028 B.n264 B.n263 10.6151
R3029 B.n267 B.n264 10.6151
R3030 B.n268 B.n267 10.6151
R3031 B.n271 B.n268 10.6151
R3032 B.n272 B.n271 10.6151
R3033 B.n275 B.n272 10.6151
R3034 B.n276 B.n275 10.6151
R3035 B.n279 B.n276 10.6151
R3036 B.n280 B.n279 10.6151
R3037 B.n283 B.n280 10.6151
R3038 B.n284 B.n283 10.6151
R3039 B.n287 B.n284 10.6151
R3040 B.n288 B.n287 10.6151
R3041 B.n291 B.n288 10.6151
R3042 B.n292 B.n291 10.6151
R3043 B.n296 B.n295 10.6151
R3044 B.n299 B.n296 10.6151
R3045 B.n300 B.n299 10.6151
R3046 B.n303 B.n300 10.6151
R3047 B.n304 B.n303 10.6151
R3048 B.n307 B.n304 10.6151
R3049 B.n308 B.n307 10.6151
R3050 B.n311 B.n308 10.6151
R3051 B.n316 B.n313 10.6151
R3052 B.n317 B.n316 10.6151
R3053 B.n320 B.n317 10.6151
R3054 B.n321 B.n320 10.6151
R3055 B.n324 B.n321 10.6151
R3056 B.n325 B.n324 10.6151
R3057 B.n328 B.n325 10.6151
R3058 B.n329 B.n328 10.6151
R3059 B.n332 B.n329 10.6151
R3060 B.n333 B.n332 10.6151
R3061 B.n336 B.n333 10.6151
R3062 B.n337 B.n336 10.6151
R3063 B.n340 B.n337 10.6151
R3064 B.n341 B.n340 10.6151
R3065 B.n344 B.n341 10.6151
R3066 B.n345 B.n344 10.6151
R3067 B.n348 B.n345 10.6151
R3068 B.n349 B.n348 10.6151
R3069 B.n352 B.n349 10.6151
R3070 B.n353 B.n352 10.6151
R3071 B.n356 B.n353 10.6151
R3072 B.n357 B.n356 10.6151
R3073 B.n360 B.n357 10.6151
R3074 B.n361 B.n360 10.6151
R3075 B.n364 B.n361 10.6151
R3076 B.n365 B.n364 10.6151
R3077 B.n368 B.n365 10.6151
R3078 B.n369 B.n368 10.6151
R3079 B.n372 B.n369 10.6151
R3080 B.n373 B.n372 10.6151
R3081 B.n376 B.n373 10.6151
R3082 B.n377 B.n376 10.6151
R3083 B.n380 B.n377 10.6151
R3084 B.n381 B.n380 10.6151
R3085 B.n384 B.n381 10.6151
R3086 B.n385 B.n384 10.6151
R3087 B.n388 B.n385 10.6151
R3088 B.n389 B.n388 10.6151
R3089 B.n392 B.n389 10.6151
R3090 B.n393 B.n392 10.6151
R3091 B.n396 B.n393 10.6151
R3092 B.n397 B.n396 10.6151
R3093 B.n400 B.n397 10.6151
R3094 B.n401 B.n400 10.6151
R3095 B.n404 B.n401 10.6151
R3096 B.n405 B.n404 10.6151
R3097 B.n408 B.n405 10.6151
R3098 B.n409 B.n408 10.6151
R3099 B.n412 B.n409 10.6151
R3100 B.n413 B.n412 10.6151
R3101 B.n416 B.n413 10.6151
R3102 B.n417 B.n416 10.6151
R3103 B.n420 B.n417 10.6151
R3104 B.n421 B.n420 10.6151
R3105 B.n424 B.n421 10.6151
R3106 B.n425 B.n424 10.6151
R3107 B.n428 B.n425 10.6151
R3108 B.n429 B.n428 10.6151
R3109 B.n432 B.n429 10.6151
R3110 B.n433 B.n432 10.6151
R3111 B.n436 B.n433 10.6151
R3112 B.n437 B.n436 10.6151
R3113 B.n1093 B.n437 10.6151
R3114 B.n1197 B.n0 8.11757
R3115 B.n1197 B.n1 8.11757
R3116 B.n1012 B.t2 7.9635
R3117 B.n1183 B.t4 7.9635
R3118 B.n749 B.n748 6.5566
R3119 B.n732 B.n606 6.5566
R3120 B.n295 B.n165 6.5566
R3121 B.n312 B.n311 6.5566
R3122 B.n750 B.n749 4.05904
R3123 B.n729 B.n606 4.05904
R3124 B.n292 B.n165 4.05904
R3125 B.n313 B.n312 4.05904
R3126 B.n944 B.t1 2.65483
R3127 B.n54 B.t3 2.65483
R3128 VN.n23 VN.t3 181.173
R3129 VN.n5 VN.t0 181.173
R3130 VN.n34 VN.n33 161.3
R3131 VN.n32 VN.n19 161.3
R3132 VN.n31 VN.n30 161.3
R3133 VN.n29 VN.n20 161.3
R3134 VN.n28 VN.n27 161.3
R3135 VN.n26 VN.n21 161.3
R3136 VN.n25 VN.n24 161.3
R3137 VN.n16 VN.n15 161.3
R3138 VN.n14 VN.n1 161.3
R3139 VN.n13 VN.n12 161.3
R3140 VN.n11 VN.n2 161.3
R3141 VN.n10 VN.n9 161.3
R3142 VN.n8 VN.n3 161.3
R3143 VN.n7 VN.n6 161.3
R3144 VN.n4 VN.t4 148.465
R3145 VN.n0 VN.t1 148.465
R3146 VN.n22 VN.t5 148.465
R3147 VN.n18 VN.t2 148.465
R3148 VN.n17 VN.n0 77.3446
R3149 VN.n35 VN.n18 77.3446
R3150 VN.n5 VN.n4 62.0351
R3151 VN.n23 VN.n22 62.0351
R3152 VN VN.n35 56.9185
R3153 VN.n13 VN.n2 40.979
R3154 VN.n31 VN.n20 40.979
R3155 VN.n9 VN.n2 40.0078
R3156 VN.n27 VN.n20 40.0078
R3157 VN.n8 VN.n7 24.4675
R3158 VN.n9 VN.n8 24.4675
R3159 VN.n14 VN.n13 24.4675
R3160 VN.n15 VN.n14 24.4675
R3161 VN.n27 VN.n26 24.4675
R3162 VN.n26 VN.n25 24.4675
R3163 VN.n33 VN.n32 24.4675
R3164 VN.n32 VN.n31 24.4675
R3165 VN.n15 VN.n0 12.7233
R3166 VN.n33 VN.n18 12.7233
R3167 VN.n7 VN.n4 12.234
R3168 VN.n25 VN.n22 12.234
R3169 VN.n24 VN.n23 4.25368
R3170 VN.n6 VN.n5 4.25368
R3171 VN.n35 VN.n34 0.354971
R3172 VN.n17 VN.n16 0.354971
R3173 VN VN.n17 0.26696
R3174 VN.n34 VN.n19 0.189894
R3175 VN.n30 VN.n19 0.189894
R3176 VN.n30 VN.n29 0.189894
R3177 VN.n29 VN.n28 0.189894
R3178 VN.n28 VN.n21 0.189894
R3179 VN.n24 VN.n21 0.189894
R3180 VN.n6 VN.n3 0.189894
R3181 VN.n10 VN.n3 0.189894
R3182 VN.n11 VN.n10 0.189894
R3183 VN.n12 VN.n11 0.189894
R3184 VN.n12 VN.n1 0.189894
R3185 VN.n16 VN.n1 0.189894
R3186 VDD2.n215 VDD2.n111 289.615
R3187 VDD2.n104 VDD2.n0 289.615
R3188 VDD2.n216 VDD2.n215 185
R3189 VDD2.n214 VDD2.n213 185
R3190 VDD2.n115 VDD2.n114 185
R3191 VDD2.n208 VDD2.n207 185
R3192 VDD2.n206 VDD2.n205 185
R3193 VDD2.n119 VDD2.n118 185
R3194 VDD2.n200 VDD2.n199 185
R3195 VDD2.n198 VDD2.n197 185
R3196 VDD2.n123 VDD2.n122 185
R3197 VDD2.n127 VDD2.n125 185
R3198 VDD2.n192 VDD2.n191 185
R3199 VDD2.n190 VDD2.n189 185
R3200 VDD2.n129 VDD2.n128 185
R3201 VDD2.n184 VDD2.n183 185
R3202 VDD2.n182 VDD2.n181 185
R3203 VDD2.n133 VDD2.n132 185
R3204 VDD2.n176 VDD2.n175 185
R3205 VDD2.n174 VDD2.n173 185
R3206 VDD2.n137 VDD2.n136 185
R3207 VDD2.n168 VDD2.n167 185
R3208 VDD2.n166 VDD2.n165 185
R3209 VDD2.n141 VDD2.n140 185
R3210 VDD2.n160 VDD2.n159 185
R3211 VDD2.n158 VDD2.n157 185
R3212 VDD2.n145 VDD2.n144 185
R3213 VDD2.n152 VDD2.n151 185
R3214 VDD2.n150 VDD2.n149 185
R3215 VDD2.n37 VDD2.n36 185
R3216 VDD2.n39 VDD2.n38 185
R3217 VDD2.n32 VDD2.n31 185
R3218 VDD2.n45 VDD2.n44 185
R3219 VDD2.n47 VDD2.n46 185
R3220 VDD2.n28 VDD2.n27 185
R3221 VDD2.n53 VDD2.n52 185
R3222 VDD2.n55 VDD2.n54 185
R3223 VDD2.n24 VDD2.n23 185
R3224 VDD2.n61 VDD2.n60 185
R3225 VDD2.n63 VDD2.n62 185
R3226 VDD2.n20 VDD2.n19 185
R3227 VDD2.n69 VDD2.n68 185
R3228 VDD2.n71 VDD2.n70 185
R3229 VDD2.n16 VDD2.n15 185
R3230 VDD2.n78 VDD2.n77 185
R3231 VDD2.n79 VDD2.n14 185
R3232 VDD2.n81 VDD2.n80 185
R3233 VDD2.n12 VDD2.n11 185
R3234 VDD2.n87 VDD2.n86 185
R3235 VDD2.n89 VDD2.n88 185
R3236 VDD2.n8 VDD2.n7 185
R3237 VDD2.n95 VDD2.n94 185
R3238 VDD2.n97 VDD2.n96 185
R3239 VDD2.n4 VDD2.n3 185
R3240 VDD2.n103 VDD2.n102 185
R3241 VDD2.n105 VDD2.n104 185
R3242 VDD2.n148 VDD2.t3 147.659
R3243 VDD2.n35 VDD2.t5 147.659
R3244 VDD2.n215 VDD2.n214 104.615
R3245 VDD2.n214 VDD2.n114 104.615
R3246 VDD2.n207 VDD2.n114 104.615
R3247 VDD2.n207 VDD2.n206 104.615
R3248 VDD2.n206 VDD2.n118 104.615
R3249 VDD2.n199 VDD2.n118 104.615
R3250 VDD2.n199 VDD2.n198 104.615
R3251 VDD2.n198 VDD2.n122 104.615
R3252 VDD2.n127 VDD2.n122 104.615
R3253 VDD2.n191 VDD2.n127 104.615
R3254 VDD2.n191 VDD2.n190 104.615
R3255 VDD2.n190 VDD2.n128 104.615
R3256 VDD2.n183 VDD2.n128 104.615
R3257 VDD2.n183 VDD2.n182 104.615
R3258 VDD2.n182 VDD2.n132 104.615
R3259 VDD2.n175 VDD2.n132 104.615
R3260 VDD2.n175 VDD2.n174 104.615
R3261 VDD2.n174 VDD2.n136 104.615
R3262 VDD2.n167 VDD2.n136 104.615
R3263 VDD2.n167 VDD2.n166 104.615
R3264 VDD2.n166 VDD2.n140 104.615
R3265 VDD2.n159 VDD2.n140 104.615
R3266 VDD2.n159 VDD2.n158 104.615
R3267 VDD2.n158 VDD2.n144 104.615
R3268 VDD2.n151 VDD2.n144 104.615
R3269 VDD2.n151 VDD2.n150 104.615
R3270 VDD2.n38 VDD2.n37 104.615
R3271 VDD2.n38 VDD2.n31 104.615
R3272 VDD2.n45 VDD2.n31 104.615
R3273 VDD2.n46 VDD2.n45 104.615
R3274 VDD2.n46 VDD2.n27 104.615
R3275 VDD2.n53 VDD2.n27 104.615
R3276 VDD2.n54 VDD2.n53 104.615
R3277 VDD2.n54 VDD2.n23 104.615
R3278 VDD2.n61 VDD2.n23 104.615
R3279 VDD2.n62 VDD2.n61 104.615
R3280 VDD2.n62 VDD2.n19 104.615
R3281 VDD2.n69 VDD2.n19 104.615
R3282 VDD2.n70 VDD2.n69 104.615
R3283 VDD2.n70 VDD2.n15 104.615
R3284 VDD2.n78 VDD2.n15 104.615
R3285 VDD2.n79 VDD2.n78 104.615
R3286 VDD2.n80 VDD2.n79 104.615
R3287 VDD2.n80 VDD2.n11 104.615
R3288 VDD2.n87 VDD2.n11 104.615
R3289 VDD2.n88 VDD2.n87 104.615
R3290 VDD2.n88 VDD2.n7 104.615
R3291 VDD2.n95 VDD2.n7 104.615
R3292 VDD2.n96 VDD2.n95 104.615
R3293 VDD2.n96 VDD2.n3 104.615
R3294 VDD2.n103 VDD2.n3 104.615
R3295 VDD2.n104 VDD2.n103 104.615
R3296 VDD2.n110 VDD2.n109 59.5576
R3297 VDD2 VDD2.n221 59.5548
R3298 VDD2.n150 VDD2.t3 52.3082
R3299 VDD2.n37 VDD2.t5 52.3082
R3300 VDD2.n220 VDD2.n110 50.4373
R3301 VDD2.n110 VDD2.n108 49.3327
R3302 VDD2.n220 VDD2.n219 47.1187
R3303 VDD2.n149 VDD2.n148 15.6677
R3304 VDD2.n36 VDD2.n35 15.6677
R3305 VDD2.n125 VDD2.n123 13.1884
R3306 VDD2.n81 VDD2.n12 13.1884
R3307 VDD2.n197 VDD2.n196 12.8005
R3308 VDD2.n193 VDD2.n192 12.8005
R3309 VDD2.n152 VDD2.n147 12.8005
R3310 VDD2.n39 VDD2.n34 12.8005
R3311 VDD2.n82 VDD2.n14 12.8005
R3312 VDD2.n86 VDD2.n85 12.8005
R3313 VDD2.n200 VDD2.n121 12.0247
R3314 VDD2.n189 VDD2.n126 12.0247
R3315 VDD2.n153 VDD2.n145 12.0247
R3316 VDD2.n40 VDD2.n32 12.0247
R3317 VDD2.n77 VDD2.n76 12.0247
R3318 VDD2.n89 VDD2.n10 12.0247
R3319 VDD2.n201 VDD2.n119 11.249
R3320 VDD2.n188 VDD2.n129 11.249
R3321 VDD2.n157 VDD2.n156 11.249
R3322 VDD2.n44 VDD2.n43 11.249
R3323 VDD2.n75 VDD2.n16 11.249
R3324 VDD2.n90 VDD2.n8 11.249
R3325 VDD2.n205 VDD2.n204 10.4732
R3326 VDD2.n185 VDD2.n184 10.4732
R3327 VDD2.n160 VDD2.n143 10.4732
R3328 VDD2.n47 VDD2.n30 10.4732
R3329 VDD2.n72 VDD2.n71 10.4732
R3330 VDD2.n94 VDD2.n93 10.4732
R3331 VDD2.n208 VDD2.n117 9.69747
R3332 VDD2.n181 VDD2.n131 9.69747
R3333 VDD2.n161 VDD2.n141 9.69747
R3334 VDD2.n48 VDD2.n28 9.69747
R3335 VDD2.n68 VDD2.n18 9.69747
R3336 VDD2.n97 VDD2.n6 9.69747
R3337 VDD2.n219 VDD2.n218 9.45567
R3338 VDD2.n108 VDD2.n107 9.45567
R3339 VDD2.n135 VDD2.n134 9.3005
R3340 VDD2.n178 VDD2.n177 9.3005
R3341 VDD2.n180 VDD2.n179 9.3005
R3342 VDD2.n131 VDD2.n130 9.3005
R3343 VDD2.n186 VDD2.n185 9.3005
R3344 VDD2.n188 VDD2.n187 9.3005
R3345 VDD2.n126 VDD2.n124 9.3005
R3346 VDD2.n194 VDD2.n193 9.3005
R3347 VDD2.n218 VDD2.n217 9.3005
R3348 VDD2.n113 VDD2.n112 9.3005
R3349 VDD2.n212 VDD2.n211 9.3005
R3350 VDD2.n210 VDD2.n209 9.3005
R3351 VDD2.n117 VDD2.n116 9.3005
R3352 VDD2.n204 VDD2.n203 9.3005
R3353 VDD2.n202 VDD2.n201 9.3005
R3354 VDD2.n121 VDD2.n120 9.3005
R3355 VDD2.n196 VDD2.n195 9.3005
R3356 VDD2.n172 VDD2.n171 9.3005
R3357 VDD2.n170 VDD2.n169 9.3005
R3358 VDD2.n139 VDD2.n138 9.3005
R3359 VDD2.n164 VDD2.n163 9.3005
R3360 VDD2.n162 VDD2.n161 9.3005
R3361 VDD2.n143 VDD2.n142 9.3005
R3362 VDD2.n156 VDD2.n155 9.3005
R3363 VDD2.n154 VDD2.n153 9.3005
R3364 VDD2.n147 VDD2.n146 9.3005
R3365 VDD2.n107 VDD2.n106 9.3005
R3366 VDD2.n101 VDD2.n100 9.3005
R3367 VDD2.n99 VDD2.n98 9.3005
R3368 VDD2.n6 VDD2.n5 9.3005
R3369 VDD2.n93 VDD2.n92 9.3005
R3370 VDD2.n91 VDD2.n90 9.3005
R3371 VDD2.n10 VDD2.n9 9.3005
R3372 VDD2.n85 VDD2.n84 9.3005
R3373 VDD2.n57 VDD2.n56 9.3005
R3374 VDD2.n26 VDD2.n25 9.3005
R3375 VDD2.n51 VDD2.n50 9.3005
R3376 VDD2.n49 VDD2.n48 9.3005
R3377 VDD2.n30 VDD2.n29 9.3005
R3378 VDD2.n43 VDD2.n42 9.3005
R3379 VDD2.n41 VDD2.n40 9.3005
R3380 VDD2.n34 VDD2.n33 9.3005
R3381 VDD2.n59 VDD2.n58 9.3005
R3382 VDD2.n22 VDD2.n21 9.3005
R3383 VDD2.n65 VDD2.n64 9.3005
R3384 VDD2.n67 VDD2.n66 9.3005
R3385 VDD2.n18 VDD2.n17 9.3005
R3386 VDD2.n73 VDD2.n72 9.3005
R3387 VDD2.n75 VDD2.n74 9.3005
R3388 VDD2.n76 VDD2.n13 9.3005
R3389 VDD2.n83 VDD2.n82 9.3005
R3390 VDD2.n2 VDD2.n1 9.3005
R3391 VDD2.n209 VDD2.n115 8.92171
R3392 VDD2.n180 VDD2.n133 8.92171
R3393 VDD2.n165 VDD2.n164 8.92171
R3394 VDD2.n52 VDD2.n51 8.92171
R3395 VDD2.n67 VDD2.n20 8.92171
R3396 VDD2.n98 VDD2.n4 8.92171
R3397 VDD2.n213 VDD2.n212 8.14595
R3398 VDD2.n177 VDD2.n176 8.14595
R3399 VDD2.n168 VDD2.n139 8.14595
R3400 VDD2.n55 VDD2.n26 8.14595
R3401 VDD2.n64 VDD2.n63 8.14595
R3402 VDD2.n102 VDD2.n101 8.14595
R3403 VDD2.n219 VDD2.n111 7.3702
R3404 VDD2.n216 VDD2.n113 7.3702
R3405 VDD2.n173 VDD2.n135 7.3702
R3406 VDD2.n169 VDD2.n137 7.3702
R3407 VDD2.n56 VDD2.n24 7.3702
R3408 VDD2.n60 VDD2.n22 7.3702
R3409 VDD2.n105 VDD2.n2 7.3702
R3410 VDD2.n108 VDD2.n0 7.3702
R3411 VDD2.n217 VDD2.n111 6.59444
R3412 VDD2.n217 VDD2.n216 6.59444
R3413 VDD2.n173 VDD2.n172 6.59444
R3414 VDD2.n172 VDD2.n137 6.59444
R3415 VDD2.n59 VDD2.n24 6.59444
R3416 VDD2.n60 VDD2.n59 6.59444
R3417 VDD2.n106 VDD2.n105 6.59444
R3418 VDD2.n106 VDD2.n0 6.59444
R3419 VDD2.n213 VDD2.n113 5.81868
R3420 VDD2.n176 VDD2.n135 5.81868
R3421 VDD2.n169 VDD2.n168 5.81868
R3422 VDD2.n56 VDD2.n55 5.81868
R3423 VDD2.n63 VDD2.n22 5.81868
R3424 VDD2.n102 VDD2.n2 5.81868
R3425 VDD2.n212 VDD2.n115 5.04292
R3426 VDD2.n177 VDD2.n133 5.04292
R3427 VDD2.n165 VDD2.n139 5.04292
R3428 VDD2.n52 VDD2.n26 5.04292
R3429 VDD2.n64 VDD2.n20 5.04292
R3430 VDD2.n101 VDD2.n4 5.04292
R3431 VDD2.n148 VDD2.n146 4.38563
R3432 VDD2.n35 VDD2.n33 4.38563
R3433 VDD2.n209 VDD2.n208 4.26717
R3434 VDD2.n181 VDD2.n180 4.26717
R3435 VDD2.n164 VDD2.n141 4.26717
R3436 VDD2.n51 VDD2.n28 4.26717
R3437 VDD2.n68 VDD2.n67 4.26717
R3438 VDD2.n98 VDD2.n97 4.26717
R3439 VDD2.n205 VDD2.n117 3.49141
R3440 VDD2.n184 VDD2.n131 3.49141
R3441 VDD2.n161 VDD2.n160 3.49141
R3442 VDD2.n48 VDD2.n47 3.49141
R3443 VDD2.n71 VDD2.n18 3.49141
R3444 VDD2.n94 VDD2.n6 3.49141
R3445 VDD2.n204 VDD2.n119 2.71565
R3446 VDD2.n185 VDD2.n129 2.71565
R3447 VDD2.n157 VDD2.n143 2.71565
R3448 VDD2.n44 VDD2.n30 2.71565
R3449 VDD2.n72 VDD2.n16 2.71565
R3450 VDD2.n93 VDD2.n8 2.71565
R3451 VDD2 VDD2.n220 2.32809
R3452 VDD2.n201 VDD2.n200 1.93989
R3453 VDD2.n189 VDD2.n188 1.93989
R3454 VDD2.n156 VDD2.n145 1.93989
R3455 VDD2.n43 VDD2.n32 1.93989
R3456 VDD2.n77 VDD2.n75 1.93989
R3457 VDD2.n90 VDD2.n89 1.93989
R3458 VDD2.n197 VDD2.n121 1.16414
R3459 VDD2.n192 VDD2.n126 1.16414
R3460 VDD2.n153 VDD2.n152 1.16414
R3461 VDD2.n40 VDD2.n39 1.16414
R3462 VDD2.n76 VDD2.n14 1.16414
R3463 VDD2.n86 VDD2.n10 1.16414
R3464 VDD2.n221 VDD2.t0 1.01122
R3465 VDD2.n221 VDD2.t2 1.01122
R3466 VDD2.n109 VDD2.t1 1.01122
R3467 VDD2.n109 VDD2.t4 1.01122
R3468 VDD2.n196 VDD2.n123 0.388379
R3469 VDD2.n193 VDD2.n125 0.388379
R3470 VDD2.n149 VDD2.n147 0.388379
R3471 VDD2.n36 VDD2.n34 0.388379
R3472 VDD2.n82 VDD2.n81 0.388379
R3473 VDD2.n85 VDD2.n12 0.388379
R3474 VDD2.n218 VDD2.n112 0.155672
R3475 VDD2.n211 VDD2.n112 0.155672
R3476 VDD2.n211 VDD2.n210 0.155672
R3477 VDD2.n210 VDD2.n116 0.155672
R3478 VDD2.n203 VDD2.n116 0.155672
R3479 VDD2.n203 VDD2.n202 0.155672
R3480 VDD2.n202 VDD2.n120 0.155672
R3481 VDD2.n195 VDD2.n120 0.155672
R3482 VDD2.n195 VDD2.n194 0.155672
R3483 VDD2.n194 VDD2.n124 0.155672
R3484 VDD2.n187 VDD2.n124 0.155672
R3485 VDD2.n187 VDD2.n186 0.155672
R3486 VDD2.n186 VDD2.n130 0.155672
R3487 VDD2.n179 VDD2.n130 0.155672
R3488 VDD2.n179 VDD2.n178 0.155672
R3489 VDD2.n178 VDD2.n134 0.155672
R3490 VDD2.n171 VDD2.n134 0.155672
R3491 VDD2.n171 VDD2.n170 0.155672
R3492 VDD2.n170 VDD2.n138 0.155672
R3493 VDD2.n163 VDD2.n138 0.155672
R3494 VDD2.n163 VDD2.n162 0.155672
R3495 VDD2.n162 VDD2.n142 0.155672
R3496 VDD2.n155 VDD2.n142 0.155672
R3497 VDD2.n155 VDD2.n154 0.155672
R3498 VDD2.n154 VDD2.n146 0.155672
R3499 VDD2.n41 VDD2.n33 0.155672
R3500 VDD2.n42 VDD2.n41 0.155672
R3501 VDD2.n42 VDD2.n29 0.155672
R3502 VDD2.n49 VDD2.n29 0.155672
R3503 VDD2.n50 VDD2.n49 0.155672
R3504 VDD2.n50 VDD2.n25 0.155672
R3505 VDD2.n57 VDD2.n25 0.155672
R3506 VDD2.n58 VDD2.n57 0.155672
R3507 VDD2.n58 VDD2.n21 0.155672
R3508 VDD2.n65 VDD2.n21 0.155672
R3509 VDD2.n66 VDD2.n65 0.155672
R3510 VDD2.n66 VDD2.n17 0.155672
R3511 VDD2.n73 VDD2.n17 0.155672
R3512 VDD2.n74 VDD2.n73 0.155672
R3513 VDD2.n74 VDD2.n13 0.155672
R3514 VDD2.n83 VDD2.n13 0.155672
R3515 VDD2.n84 VDD2.n83 0.155672
R3516 VDD2.n84 VDD2.n9 0.155672
R3517 VDD2.n91 VDD2.n9 0.155672
R3518 VDD2.n92 VDD2.n91 0.155672
R3519 VDD2.n92 VDD2.n5 0.155672
R3520 VDD2.n99 VDD2.n5 0.155672
R3521 VDD2.n100 VDD2.n99 0.155672
R3522 VDD2.n100 VDD2.n1 0.155672
R3523 VDD2.n107 VDD2.n1 0.155672
C0 VN VTAIL 11.074f
C1 VN VDD1 0.15133f
C2 VTAIL VDD1 10.449901f
C3 VN VDD2 11.1254f
C4 VN VP 8.900161f
C5 VTAIL VDD2 10.5037f
C6 VTAIL VP 11.088401f
C7 VDD1 VDD2 1.6325f
C8 VDD1 VP 11.4777f
C9 VDD2 VP 0.50781f
C10 VDD2 B 7.775245f
C11 VDD1 B 7.925521f
C12 VTAIL B 11.268877f
C13 VN B 15.220701f
C14 VP B 13.797174f
C15 VDD2.n0 B 0.029469f
C16 VDD2.n1 B 0.021066f
C17 VDD2.n2 B 0.01132f
C18 VDD2.n3 B 0.026757f
C19 VDD2.n4 B 0.011986f
C20 VDD2.n5 B 0.021066f
C21 VDD2.n6 B 0.01132f
C22 VDD2.n7 B 0.026757f
C23 VDD2.n8 B 0.011986f
C24 VDD2.n9 B 0.021066f
C25 VDD2.n10 B 0.01132f
C26 VDD2.n11 B 0.026757f
C27 VDD2.n12 B 0.011653f
C28 VDD2.n13 B 0.021066f
C29 VDD2.n14 B 0.011986f
C30 VDD2.n15 B 0.026757f
C31 VDD2.n16 B 0.011986f
C32 VDD2.n17 B 0.021066f
C33 VDD2.n18 B 0.01132f
C34 VDD2.n19 B 0.026757f
C35 VDD2.n20 B 0.011986f
C36 VDD2.n21 B 0.021066f
C37 VDD2.n22 B 0.01132f
C38 VDD2.n23 B 0.026757f
C39 VDD2.n24 B 0.011986f
C40 VDD2.n25 B 0.021066f
C41 VDD2.n26 B 0.01132f
C42 VDD2.n27 B 0.026757f
C43 VDD2.n28 B 0.011986f
C44 VDD2.n29 B 0.021066f
C45 VDD2.n30 B 0.01132f
C46 VDD2.n31 B 0.026757f
C47 VDD2.n32 B 0.011986f
C48 VDD2.n33 B 1.81376f
C49 VDD2.n34 B 0.01132f
C50 VDD2.t5 B 0.04445f
C51 VDD2.n35 B 0.161643f
C52 VDD2.n36 B 0.015806f
C53 VDD2.n37 B 0.020068f
C54 VDD2.n38 B 0.026757f
C55 VDD2.n39 B 0.011986f
C56 VDD2.n40 B 0.01132f
C57 VDD2.n41 B 0.021066f
C58 VDD2.n42 B 0.021066f
C59 VDD2.n43 B 0.01132f
C60 VDD2.n44 B 0.011986f
C61 VDD2.n45 B 0.026757f
C62 VDD2.n46 B 0.026757f
C63 VDD2.n47 B 0.011986f
C64 VDD2.n48 B 0.01132f
C65 VDD2.n49 B 0.021066f
C66 VDD2.n50 B 0.021066f
C67 VDD2.n51 B 0.01132f
C68 VDD2.n52 B 0.011986f
C69 VDD2.n53 B 0.026757f
C70 VDD2.n54 B 0.026757f
C71 VDD2.n55 B 0.011986f
C72 VDD2.n56 B 0.01132f
C73 VDD2.n57 B 0.021066f
C74 VDD2.n58 B 0.021066f
C75 VDD2.n59 B 0.01132f
C76 VDD2.n60 B 0.011986f
C77 VDD2.n61 B 0.026757f
C78 VDD2.n62 B 0.026757f
C79 VDD2.n63 B 0.011986f
C80 VDD2.n64 B 0.01132f
C81 VDD2.n65 B 0.021066f
C82 VDD2.n66 B 0.021066f
C83 VDD2.n67 B 0.01132f
C84 VDD2.n68 B 0.011986f
C85 VDD2.n69 B 0.026757f
C86 VDD2.n70 B 0.026757f
C87 VDD2.n71 B 0.011986f
C88 VDD2.n72 B 0.01132f
C89 VDD2.n73 B 0.021066f
C90 VDD2.n74 B 0.021066f
C91 VDD2.n75 B 0.01132f
C92 VDD2.n76 B 0.01132f
C93 VDD2.n77 B 0.011986f
C94 VDD2.n78 B 0.026757f
C95 VDD2.n79 B 0.026757f
C96 VDD2.n80 B 0.026757f
C97 VDD2.n81 B 0.011653f
C98 VDD2.n82 B 0.01132f
C99 VDD2.n83 B 0.021066f
C100 VDD2.n84 B 0.021066f
C101 VDD2.n85 B 0.01132f
C102 VDD2.n86 B 0.011986f
C103 VDD2.n87 B 0.026757f
C104 VDD2.n88 B 0.026757f
C105 VDD2.n89 B 0.011986f
C106 VDD2.n90 B 0.01132f
C107 VDD2.n91 B 0.021066f
C108 VDD2.n92 B 0.021066f
C109 VDD2.n93 B 0.01132f
C110 VDD2.n94 B 0.011986f
C111 VDD2.n95 B 0.026757f
C112 VDD2.n96 B 0.026757f
C113 VDD2.n97 B 0.011986f
C114 VDD2.n98 B 0.01132f
C115 VDD2.n99 B 0.021066f
C116 VDD2.n100 B 0.021066f
C117 VDD2.n101 B 0.01132f
C118 VDD2.n102 B 0.011986f
C119 VDD2.n103 B 0.026757f
C120 VDD2.n104 B 0.057673f
C121 VDD2.n105 B 0.011986f
C122 VDD2.n106 B 0.01132f
C123 VDD2.n107 B 0.046104f
C124 VDD2.n108 B 0.055239f
C125 VDD2.t1 B 0.326121f
C126 VDD2.t4 B 0.326121f
C127 VDD2.n109 B 2.98323f
C128 VDD2.n110 B 2.87274f
C129 VDD2.n111 B 0.029469f
C130 VDD2.n112 B 0.021066f
C131 VDD2.n113 B 0.01132f
C132 VDD2.n114 B 0.026757f
C133 VDD2.n115 B 0.011986f
C134 VDD2.n116 B 0.021066f
C135 VDD2.n117 B 0.01132f
C136 VDD2.n118 B 0.026757f
C137 VDD2.n119 B 0.011986f
C138 VDD2.n120 B 0.021066f
C139 VDD2.n121 B 0.01132f
C140 VDD2.n122 B 0.026757f
C141 VDD2.n123 B 0.011653f
C142 VDD2.n124 B 0.021066f
C143 VDD2.n125 B 0.011653f
C144 VDD2.n126 B 0.01132f
C145 VDD2.n127 B 0.026757f
C146 VDD2.n128 B 0.026757f
C147 VDD2.n129 B 0.011986f
C148 VDD2.n130 B 0.021066f
C149 VDD2.n131 B 0.01132f
C150 VDD2.n132 B 0.026757f
C151 VDD2.n133 B 0.011986f
C152 VDD2.n134 B 0.021066f
C153 VDD2.n135 B 0.01132f
C154 VDD2.n136 B 0.026757f
C155 VDD2.n137 B 0.011986f
C156 VDD2.n138 B 0.021066f
C157 VDD2.n139 B 0.01132f
C158 VDD2.n140 B 0.026757f
C159 VDD2.n141 B 0.011986f
C160 VDD2.n142 B 0.021066f
C161 VDD2.n143 B 0.01132f
C162 VDD2.n144 B 0.026757f
C163 VDD2.n145 B 0.011986f
C164 VDD2.n146 B 1.81376f
C165 VDD2.n147 B 0.01132f
C166 VDD2.t3 B 0.04445f
C167 VDD2.n148 B 0.161643f
C168 VDD2.n149 B 0.015806f
C169 VDD2.n150 B 0.020068f
C170 VDD2.n151 B 0.026757f
C171 VDD2.n152 B 0.011986f
C172 VDD2.n153 B 0.01132f
C173 VDD2.n154 B 0.021066f
C174 VDD2.n155 B 0.021066f
C175 VDD2.n156 B 0.01132f
C176 VDD2.n157 B 0.011986f
C177 VDD2.n158 B 0.026757f
C178 VDD2.n159 B 0.026757f
C179 VDD2.n160 B 0.011986f
C180 VDD2.n161 B 0.01132f
C181 VDD2.n162 B 0.021066f
C182 VDD2.n163 B 0.021066f
C183 VDD2.n164 B 0.01132f
C184 VDD2.n165 B 0.011986f
C185 VDD2.n166 B 0.026757f
C186 VDD2.n167 B 0.026757f
C187 VDD2.n168 B 0.011986f
C188 VDD2.n169 B 0.01132f
C189 VDD2.n170 B 0.021066f
C190 VDD2.n171 B 0.021066f
C191 VDD2.n172 B 0.01132f
C192 VDD2.n173 B 0.011986f
C193 VDD2.n174 B 0.026757f
C194 VDD2.n175 B 0.026757f
C195 VDD2.n176 B 0.011986f
C196 VDD2.n177 B 0.01132f
C197 VDD2.n178 B 0.021066f
C198 VDD2.n179 B 0.021066f
C199 VDD2.n180 B 0.01132f
C200 VDD2.n181 B 0.011986f
C201 VDD2.n182 B 0.026757f
C202 VDD2.n183 B 0.026757f
C203 VDD2.n184 B 0.011986f
C204 VDD2.n185 B 0.01132f
C205 VDD2.n186 B 0.021066f
C206 VDD2.n187 B 0.021066f
C207 VDD2.n188 B 0.01132f
C208 VDD2.n189 B 0.011986f
C209 VDD2.n190 B 0.026757f
C210 VDD2.n191 B 0.026757f
C211 VDD2.n192 B 0.011986f
C212 VDD2.n193 B 0.01132f
C213 VDD2.n194 B 0.021066f
C214 VDD2.n195 B 0.021066f
C215 VDD2.n196 B 0.01132f
C216 VDD2.n197 B 0.011986f
C217 VDD2.n198 B 0.026757f
C218 VDD2.n199 B 0.026757f
C219 VDD2.n200 B 0.011986f
C220 VDD2.n201 B 0.01132f
C221 VDD2.n202 B 0.021066f
C222 VDD2.n203 B 0.021066f
C223 VDD2.n204 B 0.01132f
C224 VDD2.n205 B 0.011986f
C225 VDD2.n206 B 0.026757f
C226 VDD2.n207 B 0.026757f
C227 VDD2.n208 B 0.011986f
C228 VDD2.n209 B 0.01132f
C229 VDD2.n210 B 0.021066f
C230 VDD2.n211 B 0.021066f
C231 VDD2.n212 B 0.01132f
C232 VDD2.n213 B 0.011986f
C233 VDD2.n214 B 0.026757f
C234 VDD2.n215 B 0.057673f
C235 VDD2.n216 B 0.011986f
C236 VDD2.n217 B 0.01132f
C237 VDD2.n218 B 0.046104f
C238 VDD2.n219 B 0.04673f
C239 VDD2.n220 B 2.77664f
C240 VDD2.t0 B 0.326121f
C241 VDD2.t2 B 0.326121f
C242 VDD2.n221 B 2.9832f
C243 VN.t1 B 3.29186f
C244 VN.n0 B 1.20465f
C245 VN.n1 B 0.019182f
C246 VN.n2 B 0.015514f
C247 VN.n3 B 0.019182f
C248 VN.t4 B 3.29186f
C249 VN.n4 B 1.19688f
C250 VN.t0 B 3.52056f
C251 VN.n5 B 1.1551f
C252 VN.n6 B 0.223139f
C253 VN.n7 B 0.026925f
C254 VN.n8 B 0.03575f
C255 VN.n9 B 0.038218f
C256 VN.n10 B 0.019182f
C257 VN.n11 B 0.019182f
C258 VN.n12 B 0.019182f
C259 VN.n13 B 0.038026f
C260 VN.n14 B 0.03575f
C261 VN.n15 B 0.027278f
C262 VN.n16 B 0.030959f
C263 VN.n17 B 0.04686f
C264 VN.t2 B 3.29186f
C265 VN.n18 B 1.20465f
C266 VN.n19 B 0.019182f
C267 VN.n20 B 0.015514f
C268 VN.n21 B 0.019182f
C269 VN.t5 B 3.29186f
C270 VN.n22 B 1.19688f
C271 VN.t3 B 3.52056f
C272 VN.n23 B 1.1551f
C273 VN.n24 B 0.223139f
C274 VN.n25 B 0.026925f
C275 VN.n26 B 0.03575f
C276 VN.n27 B 0.038218f
C277 VN.n28 B 0.019182f
C278 VN.n29 B 0.019182f
C279 VN.n30 B 0.019182f
C280 VN.n31 B 0.038026f
C281 VN.n32 B 0.03575f
C282 VN.n33 B 0.027278f
C283 VN.n34 B 0.030959f
C284 VN.n35 B 1.30961f
C285 VDD1.n0 B 0.029771f
C286 VDD1.n1 B 0.021282f
C287 VDD1.n2 B 0.011436f
C288 VDD1.n3 B 0.027031f
C289 VDD1.n4 B 0.012109f
C290 VDD1.n5 B 0.021282f
C291 VDD1.n6 B 0.011436f
C292 VDD1.n7 B 0.027031f
C293 VDD1.n8 B 0.012109f
C294 VDD1.n9 B 0.021282f
C295 VDD1.n10 B 0.011436f
C296 VDD1.n11 B 0.027031f
C297 VDD1.n12 B 0.011773f
C298 VDD1.n13 B 0.021282f
C299 VDD1.n14 B 0.011773f
C300 VDD1.n15 B 0.011436f
C301 VDD1.n16 B 0.027031f
C302 VDD1.n17 B 0.027031f
C303 VDD1.n18 B 0.012109f
C304 VDD1.n19 B 0.021282f
C305 VDD1.n20 B 0.011436f
C306 VDD1.n21 B 0.027031f
C307 VDD1.n22 B 0.012109f
C308 VDD1.n23 B 0.021282f
C309 VDD1.n24 B 0.011436f
C310 VDD1.n25 B 0.027031f
C311 VDD1.n26 B 0.012109f
C312 VDD1.n27 B 0.021282f
C313 VDD1.n28 B 0.011436f
C314 VDD1.n29 B 0.027031f
C315 VDD1.n30 B 0.012109f
C316 VDD1.n31 B 0.021282f
C317 VDD1.n32 B 0.011436f
C318 VDD1.n33 B 0.027031f
C319 VDD1.n34 B 0.012109f
C320 VDD1.n35 B 1.83235f
C321 VDD1.n36 B 0.011436f
C322 VDD1.t5 B 0.044906f
C323 VDD1.n37 B 0.1633f
C324 VDD1.n38 B 0.015968f
C325 VDD1.n39 B 0.020273f
C326 VDD1.n40 B 0.027031f
C327 VDD1.n41 B 0.012109f
C328 VDD1.n42 B 0.011436f
C329 VDD1.n43 B 0.021282f
C330 VDD1.n44 B 0.021282f
C331 VDD1.n45 B 0.011436f
C332 VDD1.n46 B 0.012109f
C333 VDD1.n47 B 0.027031f
C334 VDD1.n48 B 0.027031f
C335 VDD1.n49 B 0.012109f
C336 VDD1.n50 B 0.011436f
C337 VDD1.n51 B 0.021282f
C338 VDD1.n52 B 0.021282f
C339 VDD1.n53 B 0.011436f
C340 VDD1.n54 B 0.012109f
C341 VDD1.n55 B 0.027031f
C342 VDD1.n56 B 0.027031f
C343 VDD1.n57 B 0.012109f
C344 VDD1.n58 B 0.011436f
C345 VDD1.n59 B 0.021282f
C346 VDD1.n60 B 0.021282f
C347 VDD1.n61 B 0.011436f
C348 VDD1.n62 B 0.012109f
C349 VDD1.n63 B 0.027031f
C350 VDD1.n64 B 0.027031f
C351 VDD1.n65 B 0.012109f
C352 VDD1.n66 B 0.011436f
C353 VDD1.n67 B 0.021282f
C354 VDD1.n68 B 0.021282f
C355 VDD1.n69 B 0.011436f
C356 VDD1.n70 B 0.012109f
C357 VDD1.n71 B 0.027031f
C358 VDD1.n72 B 0.027031f
C359 VDD1.n73 B 0.012109f
C360 VDD1.n74 B 0.011436f
C361 VDD1.n75 B 0.021282f
C362 VDD1.n76 B 0.021282f
C363 VDD1.n77 B 0.011436f
C364 VDD1.n78 B 0.012109f
C365 VDD1.n79 B 0.027031f
C366 VDD1.n80 B 0.027031f
C367 VDD1.n81 B 0.012109f
C368 VDD1.n82 B 0.011436f
C369 VDD1.n83 B 0.021282f
C370 VDD1.n84 B 0.021282f
C371 VDD1.n85 B 0.011436f
C372 VDD1.n86 B 0.012109f
C373 VDD1.n87 B 0.027031f
C374 VDD1.n88 B 0.027031f
C375 VDD1.n89 B 0.012109f
C376 VDD1.n90 B 0.011436f
C377 VDD1.n91 B 0.021282f
C378 VDD1.n92 B 0.021282f
C379 VDD1.n93 B 0.011436f
C380 VDD1.n94 B 0.012109f
C381 VDD1.n95 B 0.027031f
C382 VDD1.n96 B 0.027031f
C383 VDD1.n97 B 0.012109f
C384 VDD1.n98 B 0.011436f
C385 VDD1.n99 B 0.021282f
C386 VDD1.n100 B 0.021282f
C387 VDD1.n101 B 0.011436f
C388 VDD1.n102 B 0.012109f
C389 VDD1.n103 B 0.027031f
C390 VDD1.n104 B 0.058264f
C391 VDD1.n105 B 0.012109f
C392 VDD1.n106 B 0.011436f
C393 VDD1.n107 B 0.046576f
C394 VDD1.n108 B 0.056582f
C395 VDD1.n109 B 0.029771f
C396 VDD1.n110 B 0.021282f
C397 VDD1.n111 B 0.011436f
C398 VDD1.n112 B 0.027031f
C399 VDD1.n113 B 0.012109f
C400 VDD1.n114 B 0.021282f
C401 VDD1.n115 B 0.011436f
C402 VDD1.n116 B 0.027031f
C403 VDD1.n117 B 0.012109f
C404 VDD1.n118 B 0.021282f
C405 VDD1.n119 B 0.011436f
C406 VDD1.n120 B 0.027031f
C407 VDD1.n121 B 0.011773f
C408 VDD1.n122 B 0.021282f
C409 VDD1.n123 B 0.012109f
C410 VDD1.n124 B 0.027031f
C411 VDD1.n125 B 0.012109f
C412 VDD1.n126 B 0.021282f
C413 VDD1.n127 B 0.011436f
C414 VDD1.n128 B 0.027031f
C415 VDD1.n129 B 0.012109f
C416 VDD1.n130 B 0.021282f
C417 VDD1.n131 B 0.011436f
C418 VDD1.n132 B 0.027031f
C419 VDD1.n133 B 0.012109f
C420 VDD1.n134 B 0.021282f
C421 VDD1.n135 B 0.011436f
C422 VDD1.n136 B 0.027031f
C423 VDD1.n137 B 0.012109f
C424 VDD1.n138 B 0.021282f
C425 VDD1.n139 B 0.011436f
C426 VDD1.n140 B 0.027031f
C427 VDD1.n141 B 0.012109f
C428 VDD1.n142 B 1.83235f
C429 VDD1.n143 B 0.011436f
C430 VDD1.t4 B 0.044906f
C431 VDD1.n144 B 0.1633f
C432 VDD1.n145 B 0.015968f
C433 VDD1.n146 B 0.020273f
C434 VDD1.n147 B 0.027031f
C435 VDD1.n148 B 0.012109f
C436 VDD1.n149 B 0.011436f
C437 VDD1.n150 B 0.021282f
C438 VDD1.n151 B 0.021282f
C439 VDD1.n152 B 0.011436f
C440 VDD1.n153 B 0.012109f
C441 VDD1.n154 B 0.027031f
C442 VDD1.n155 B 0.027031f
C443 VDD1.n156 B 0.012109f
C444 VDD1.n157 B 0.011436f
C445 VDD1.n158 B 0.021282f
C446 VDD1.n159 B 0.021282f
C447 VDD1.n160 B 0.011436f
C448 VDD1.n161 B 0.012109f
C449 VDD1.n162 B 0.027031f
C450 VDD1.n163 B 0.027031f
C451 VDD1.n164 B 0.012109f
C452 VDD1.n165 B 0.011436f
C453 VDD1.n166 B 0.021282f
C454 VDD1.n167 B 0.021282f
C455 VDD1.n168 B 0.011436f
C456 VDD1.n169 B 0.012109f
C457 VDD1.n170 B 0.027031f
C458 VDD1.n171 B 0.027031f
C459 VDD1.n172 B 0.012109f
C460 VDD1.n173 B 0.011436f
C461 VDD1.n174 B 0.021282f
C462 VDD1.n175 B 0.021282f
C463 VDD1.n176 B 0.011436f
C464 VDD1.n177 B 0.012109f
C465 VDD1.n178 B 0.027031f
C466 VDD1.n179 B 0.027031f
C467 VDD1.n180 B 0.012109f
C468 VDD1.n181 B 0.011436f
C469 VDD1.n182 B 0.021282f
C470 VDD1.n183 B 0.021282f
C471 VDD1.n184 B 0.011436f
C472 VDD1.n185 B 0.011436f
C473 VDD1.n186 B 0.012109f
C474 VDD1.n187 B 0.027031f
C475 VDD1.n188 B 0.027031f
C476 VDD1.n189 B 0.027031f
C477 VDD1.n190 B 0.011773f
C478 VDD1.n191 B 0.011436f
C479 VDD1.n192 B 0.021282f
C480 VDD1.n193 B 0.021282f
C481 VDD1.n194 B 0.011436f
C482 VDD1.n195 B 0.012109f
C483 VDD1.n196 B 0.027031f
C484 VDD1.n197 B 0.027031f
C485 VDD1.n198 B 0.012109f
C486 VDD1.n199 B 0.011436f
C487 VDD1.n200 B 0.021282f
C488 VDD1.n201 B 0.021282f
C489 VDD1.n202 B 0.011436f
C490 VDD1.n203 B 0.012109f
C491 VDD1.n204 B 0.027031f
C492 VDD1.n205 B 0.027031f
C493 VDD1.n206 B 0.012109f
C494 VDD1.n207 B 0.011436f
C495 VDD1.n208 B 0.021282f
C496 VDD1.n209 B 0.021282f
C497 VDD1.n210 B 0.011436f
C498 VDD1.n211 B 0.012109f
C499 VDD1.n212 B 0.027031f
C500 VDD1.n213 B 0.058264f
C501 VDD1.n214 B 0.012109f
C502 VDD1.n215 B 0.011436f
C503 VDD1.n216 B 0.046576f
C504 VDD1.n217 B 0.055806f
C505 VDD1.t1 B 0.329463f
C506 VDD1.t0 B 0.329463f
C507 VDD1.n218 B 3.01381f
C508 VDD1.n219 B 3.02552f
C509 VDD1.t2 B 0.329463f
C510 VDD1.t3 B 0.329463f
C511 VDD1.n220 B 3.00856f
C512 VDD1.n221 B 3.00571f
C513 VTAIL.t4 B 0.348475f
C514 VTAIL.t0 B 0.348475f
C515 VTAIL.n0 B 3.10838f
C516 VTAIL.n1 B 0.437006f
C517 VTAIL.n2 B 0.031489f
C518 VTAIL.n3 B 0.02251f
C519 VTAIL.n4 B 0.012096f
C520 VTAIL.n5 B 0.028591f
C521 VTAIL.n6 B 0.012808f
C522 VTAIL.n7 B 0.02251f
C523 VTAIL.n8 B 0.012096f
C524 VTAIL.n9 B 0.028591f
C525 VTAIL.n10 B 0.012808f
C526 VTAIL.n11 B 0.02251f
C527 VTAIL.n12 B 0.012096f
C528 VTAIL.n13 B 0.028591f
C529 VTAIL.n14 B 0.012452f
C530 VTAIL.n15 B 0.02251f
C531 VTAIL.n16 B 0.012808f
C532 VTAIL.n17 B 0.028591f
C533 VTAIL.n18 B 0.012808f
C534 VTAIL.n19 B 0.02251f
C535 VTAIL.n20 B 0.012096f
C536 VTAIL.n21 B 0.028591f
C537 VTAIL.n22 B 0.012808f
C538 VTAIL.n23 B 0.02251f
C539 VTAIL.n24 B 0.012096f
C540 VTAIL.n25 B 0.028591f
C541 VTAIL.n26 B 0.012808f
C542 VTAIL.n27 B 0.02251f
C543 VTAIL.n28 B 0.012096f
C544 VTAIL.n29 B 0.028591f
C545 VTAIL.n30 B 0.012808f
C546 VTAIL.n31 B 0.02251f
C547 VTAIL.n32 B 0.012096f
C548 VTAIL.n33 B 0.028591f
C549 VTAIL.n34 B 0.012808f
C550 VTAIL.n35 B 1.93809f
C551 VTAIL.n36 B 0.012096f
C552 VTAIL.t10 B 0.047497f
C553 VTAIL.n37 B 0.172723f
C554 VTAIL.n38 B 0.016889f
C555 VTAIL.n39 B 0.021443f
C556 VTAIL.n40 B 0.028591f
C557 VTAIL.n41 B 0.012808f
C558 VTAIL.n42 B 0.012096f
C559 VTAIL.n43 B 0.02251f
C560 VTAIL.n44 B 0.02251f
C561 VTAIL.n45 B 0.012096f
C562 VTAIL.n46 B 0.012808f
C563 VTAIL.n47 B 0.028591f
C564 VTAIL.n48 B 0.028591f
C565 VTAIL.n49 B 0.012808f
C566 VTAIL.n50 B 0.012096f
C567 VTAIL.n51 B 0.02251f
C568 VTAIL.n52 B 0.02251f
C569 VTAIL.n53 B 0.012096f
C570 VTAIL.n54 B 0.012808f
C571 VTAIL.n55 B 0.028591f
C572 VTAIL.n56 B 0.028591f
C573 VTAIL.n57 B 0.012808f
C574 VTAIL.n58 B 0.012096f
C575 VTAIL.n59 B 0.02251f
C576 VTAIL.n60 B 0.02251f
C577 VTAIL.n61 B 0.012096f
C578 VTAIL.n62 B 0.012808f
C579 VTAIL.n63 B 0.028591f
C580 VTAIL.n64 B 0.028591f
C581 VTAIL.n65 B 0.012808f
C582 VTAIL.n66 B 0.012096f
C583 VTAIL.n67 B 0.02251f
C584 VTAIL.n68 B 0.02251f
C585 VTAIL.n69 B 0.012096f
C586 VTAIL.n70 B 0.012808f
C587 VTAIL.n71 B 0.028591f
C588 VTAIL.n72 B 0.028591f
C589 VTAIL.n73 B 0.012808f
C590 VTAIL.n74 B 0.012096f
C591 VTAIL.n75 B 0.02251f
C592 VTAIL.n76 B 0.02251f
C593 VTAIL.n77 B 0.012096f
C594 VTAIL.n78 B 0.012096f
C595 VTAIL.n79 B 0.012808f
C596 VTAIL.n80 B 0.028591f
C597 VTAIL.n81 B 0.028591f
C598 VTAIL.n82 B 0.028591f
C599 VTAIL.n83 B 0.012452f
C600 VTAIL.n84 B 0.012096f
C601 VTAIL.n85 B 0.02251f
C602 VTAIL.n86 B 0.02251f
C603 VTAIL.n87 B 0.012096f
C604 VTAIL.n88 B 0.012808f
C605 VTAIL.n89 B 0.028591f
C606 VTAIL.n90 B 0.028591f
C607 VTAIL.n91 B 0.012808f
C608 VTAIL.n92 B 0.012096f
C609 VTAIL.n93 B 0.02251f
C610 VTAIL.n94 B 0.02251f
C611 VTAIL.n95 B 0.012096f
C612 VTAIL.n96 B 0.012808f
C613 VTAIL.n97 B 0.028591f
C614 VTAIL.n98 B 0.028591f
C615 VTAIL.n99 B 0.012808f
C616 VTAIL.n100 B 0.012096f
C617 VTAIL.n101 B 0.02251f
C618 VTAIL.n102 B 0.02251f
C619 VTAIL.n103 B 0.012096f
C620 VTAIL.n104 B 0.012808f
C621 VTAIL.n105 B 0.028591f
C622 VTAIL.n106 B 0.061626f
C623 VTAIL.n107 B 0.012808f
C624 VTAIL.n108 B 0.012096f
C625 VTAIL.n109 B 0.049264f
C626 VTAIL.n110 B 0.034367f
C627 VTAIL.n111 B 0.380959f
C628 VTAIL.t6 B 0.348475f
C629 VTAIL.t8 B 0.348475f
C630 VTAIL.n112 B 3.10838f
C631 VTAIL.n113 B 2.42325f
C632 VTAIL.t1 B 0.348475f
C633 VTAIL.t5 B 0.348475f
C634 VTAIL.n114 B 3.10839f
C635 VTAIL.n115 B 2.42324f
C636 VTAIL.n116 B 0.031489f
C637 VTAIL.n117 B 0.02251f
C638 VTAIL.n118 B 0.012096f
C639 VTAIL.n119 B 0.028591f
C640 VTAIL.n120 B 0.012808f
C641 VTAIL.n121 B 0.02251f
C642 VTAIL.n122 B 0.012096f
C643 VTAIL.n123 B 0.028591f
C644 VTAIL.n124 B 0.012808f
C645 VTAIL.n125 B 0.02251f
C646 VTAIL.n126 B 0.012096f
C647 VTAIL.n127 B 0.028591f
C648 VTAIL.n128 B 0.012452f
C649 VTAIL.n129 B 0.02251f
C650 VTAIL.n130 B 0.012452f
C651 VTAIL.n131 B 0.012096f
C652 VTAIL.n132 B 0.028591f
C653 VTAIL.n133 B 0.028591f
C654 VTAIL.n134 B 0.012808f
C655 VTAIL.n135 B 0.02251f
C656 VTAIL.n136 B 0.012096f
C657 VTAIL.n137 B 0.028591f
C658 VTAIL.n138 B 0.012808f
C659 VTAIL.n139 B 0.02251f
C660 VTAIL.n140 B 0.012096f
C661 VTAIL.n141 B 0.028591f
C662 VTAIL.n142 B 0.012808f
C663 VTAIL.n143 B 0.02251f
C664 VTAIL.n144 B 0.012096f
C665 VTAIL.n145 B 0.028591f
C666 VTAIL.n146 B 0.012808f
C667 VTAIL.n147 B 0.02251f
C668 VTAIL.n148 B 0.012096f
C669 VTAIL.n149 B 0.028591f
C670 VTAIL.n150 B 0.012808f
C671 VTAIL.n151 B 1.93809f
C672 VTAIL.n152 B 0.012096f
C673 VTAIL.t2 B 0.047497f
C674 VTAIL.n153 B 0.172723f
C675 VTAIL.n154 B 0.016889f
C676 VTAIL.n155 B 0.021443f
C677 VTAIL.n156 B 0.028591f
C678 VTAIL.n157 B 0.012808f
C679 VTAIL.n158 B 0.012096f
C680 VTAIL.n159 B 0.02251f
C681 VTAIL.n160 B 0.02251f
C682 VTAIL.n161 B 0.012096f
C683 VTAIL.n162 B 0.012808f
C684 VTAIL.n163 B 0.028591f
C685 VTAIL.n164 B 0.028591f
C686 VTAIL.n165 B 0.012808f
C687 VTAIL.n166 B 0.012096f
C688 VTAIL.n167 B 0.02251f
C689 VTAIL.n168 B 0.02251f
C690 VTAIL.n169 B 0.012096f
C691 VTAIL.n170 B 0.012808f
C692 VTAIL.n171 B 0.028591f
C693 VTAIL.n172 B 0.028591f
C694 VTAIL.n173 B 0.012808f
C695 VTAIL.n174 B 0.012096f
C696 VTAIL.n175 B 0.02251f
C697 VTAIL.n176 B 0.02251f
C698 VTAIL.n177 B 0.012096f
C699 VTAIL.n178 B 0.012808f
C700 VTAIL.n179 B 0.028591f
C701 VTAIL.n180 B 0.028591f
C702 VTAIL.n181 B 0.012808f
C703 VTAIL.n182 B 0.012096f
C704 VTAIL.n183 B 0.02251f
C705 VTAIL.n184 B 0.02251f
C706 VTAIL.n185 B 0.012096f
C707 VTAIL.n186 B 0.012808f
C708 VTAIL.n187 B 0.028591f
C709 VTAIL.n188 B 0.028591f
C710 VTAIL.n189 B 0.012808f
C711 VTAIL.n190 B 0.012096f
C712 VTAIL.n191 B 0.02251f
C713 VTAIL.n192 B 0.02251f
C714 VTAIL.n193 B 0.012096f
C715 VTAIL.n194 B 0.012808f
C716 VTAIL.n195 B 0.028591f
C717 VTAIL.n196 B 0.028591f
C718 VTAIL.n197 B 0.012808f
C719 VTAIL.n198 B 0.012096f
C720 VTAIL.n199 B 0.02251f
C721 VTAIL.n200 B 0.02251f
C722 VTAIL.n201 B 0.012096f
C723 VTAIL.n202 B 0.012808f
C724 VTAIL.n203 B 0.028591f
C725 VTAIL.n204 B 0.028591f
C726 VTAIL.n205 B 0.012808f
C727 VTAIL.n206 B 0.012096f
C728 VTAIL.n207 B 0.02251f
C729 VTAIL.n208 B 0.02251f
C730 VTAIL.n209 B 0.012096f
C731 VTAIL.n210 B 0.012808f
C732 VTAIL.n211 B 0.028591f
C733 VTAIL.n212 B 0.028591f
C734 VTAIL.n213 B 0.012808f
C735 VTAIL.n214 B 0.012096f
C736 VTAIL.n215 B 0.02251f
C737 VTAIL.n216 B 0.02251f
C738 VTAIL.n217 B 0.012096f
C739 VTAIL.n218 B 0.012808f
C740 VTAIL.n219 B 0.028591f
C741 VTAIL.n220 B 0.061626f
C742 VTAIL.n221 B 0.012808f
C743 VTAIL.n222 B 0.012096f
C744 VTAIL.n223 B 0.049264f
C745 VTAIL.n224 B 0.034367f
C746 VTAIL.n225 B 0.380959f
C747 VTAIL.t7 B 0.348475f
C748 VTAIL.t9 B 0.348475f
C749 VTAIL.n226 B 3.10839f
C750 VTAIL.n227 B 0.597379f
C751 VTAIL.n228 B 0.031489f
C752 VTAIL.n229 B 0.02251f
C753 VTAIL.n230 B 0.012096f
C754 VTAIL.n231 B 0.028591f
C755 VTAIL.n232 B 0.012808f
C756 VTAIL.n233 B 0.02251f
C757 VTAIL.n234 B 0.012096f
C758 VTAIL.n235 B 0.028591f
C759 VTAIL.n236 B 0.012808f
C760 VTAIL.n237 B 0.02251f
C761 VTAIL.n238 B 0.012096f
C762 VTAIL.n239 B 0.028591f
C763 VTAIL.n240 B 0.012452f
C764 VTAIL.n241 B 0.02251f
C765 VTAIL.n242 B 0.012452f
C766 VTAIL.n243 B 0.012096f
C767 VTAIL.n244 B 0.028591f
C768 VTAIL.n245 B 0.028591f
C769 VTAIL.n246 B 0.012808f
C770 VTAIL.n247 B 0.02251f
C771 VTAIL.n248 B 0.012096f
C772 VTAIL.n249 B 0.028591f
C773 VTAIL.n250 B 0.012808f
C774 VTAIL.n251 B 0.02251f
C775 VTAIL.n252 B 0.012096f
C776 VTAIL.n253 B 0.028591f
C777 VTAIL.n254 B 0.012808f
C778 VTAIL.n255 B 0.02251f
C779 VTAIL.n256 B 0.012096f
C780 VTAIL.n257 B 0.028591f
C781 VTAIL.n258 B 0.012808f
C782 VTAIL.n259 B 0.02251f
C783 VTAIL.n260 B 0.012096f
C784 VTAIL.n261 B 0.028591f
C785 VTAIL.n262 B 0.012808f
C786 VTAIL.n263 B 1.93809f
C787 VTAIL.n264 B 0.012096f
C788 VTAIL.t11 B 0.047497f
C789 VTAIL.n265 B 0.172723f
C790 VTAIL.n266 B 0.016889f
C791 VTAIL.n267 B 0.021443f
C792 VTAIL.n268 B 0.028591f
C793 VTAIL.n269 B 0.012808f
C794 VTAIL.n270 B 0.012096f
C795 VTAIL.n271 B 0.02251f
C796 VTAIL.n272 B 0.02251f
C797 VTAIL.n273 B 0.012096f
C798 VTAIL.n274 B 0.012808f
C799 VTAIL.n275 B 0.028591f
C800 VTAIL.n276 B 0.028591f
C801 VTAIL.n277 B 0.012808f
C802 VTAIL.n278 B 0.012096f
C803 VTAIL.n279 B 0.02251f
C804 VTAIL.n280 B 0.02251f
C805 VTAIL.n281 B 0.012096f
C806 VTAIL.n282 B 0.012808f
C807 VTAIL.n283 B 0.028591f
C808 VTAIL.n284 B 0.028591f
C809 VTAIL.n285 B 0.012808f
C810 VTAIL.n286 B 0.012096f
C811 VTAIL.n287 B 0.02251f
C812 VTAIL.n288 B 0.02251f
C813 VTAIL.n289 B 0.012096f
C814 VTAIL.n290 B 0.012808f
C815 VTAIL.n291 B 0.028591f
C816 VTAIL.n292 B 0.028591f
C817 VTAIL.n293 B 0.012808f
C818 VTAIL.n294 B 0.012096f
C819 VTAIL.n295 B 0.02251f
C820 VTAIL.n296 B 0.02251f
C821 VTAIL.n297 B 0.012096f
C822 VTAIL.n298 B 0.012808f
C823 VTAIL.n299 B 0.028591f
C824 VTAIL.n300 B 0.028591f
C825 VTAIL.n301 B 0.012808f
C826 VTAIL.n302 B 0.012096f
C827 VTAIL.n303 B 0.02251f
C828 VTAIL.n304 B 0.02251f
C829 VTAIL.n305 B 0.012096f
C830 VTAIL.n306 B 0.012808f
C831 VTAIL.n307 B 0.028591f
C832 VTAIL.n308 B 0.028591f
C833 VTAIL.n309 B 0.012808f
C834 VTAIL.n310 B 0.012096f
C835 VTAIL.n311 B 0.02251f
C836 VTAIL.n312 B 0.02251f
C837 VTAIL.n313 B 0.012096f
C838 VTAIL.n314 B 0.012808f
C839 VTAIL.n315 B 0.028591f
C840 VTAIL.n316 B 0.028591f
C841 VTAIL.n317 B 0.012808f
C842 VTAIL.n318 B 0.012096f
C843 VTAIL.n319 B 0.02251f
C844 VTAIL.n320 B 0.02251f
C845 VTAIL.n321 B 0.012096f
C846 VTAIL.n322 B 0.012808f
C847 VTAIL.n323 B 0.028591f
C848 VTAIL.n324 B 0.028591f
C849 VTAIL.n325 B 0.012808f
C850 VTAIL.n326 B 0.012096f
C851 VTAIL.n327 B 0.02251f
C852 VTAIL.n328 B 0.02251f
C853 VTAIL.n329 B 0.012096f
C854 VTAIL.n330 B 0.012808f
C855 VTAIL.n331 B 0.028591f
C856 VTAIL.n332 B 0.061626f
C857 VTAIL.n333 B 0.012808f
C858 VTAIL.n334 B 0.012096f
C859 VTAIL.n335 B 0.049264f
C860 VTAIL.n336 B 0.034367f
C861 VTAIL.n337 B 1.98734f
C862 VTAIL.n338 B 0.031489f
C863 VTAIL.n339 B 0.02251f
C864 VTAIL.n340 B 0.012096f
C865 VTAIL.n341 B 0.028591f
C866 VTAIL.n342 B 0.012808f
C867 VTAIL.n343 B 0.02251f
C868 VTAIL.n344 B 0.012096f
C869 VTAIL.n345 B 0.028591f
C870 VTAIL.n346 B 0.012808f
C871 VTAIL.n347 B 0.02251f
C872 VTAIL.n348 B 0.012096f
C873 VTAIL.n349 B 0.028591f
C874 VTAIL.n350 B 0.012452f
C875 VTAIL.n351 B 0.02251f
C876 VTAIL.n352 B 0.012808f
C877 VTAIL.n353 B 0.028591f
C878 VTAIL.n354 B 0.012808f
C879 VTAIL.n355 B 0.02251f
C880 VTAIL.n356 B 0.012096f
C881 VTAIL.n357 B 0.028591f
C882 VTAIL.n358 B 0.012808f
C883 VTAIL.n359 B 0.02251f
C884 VTAIL.n360 B 0.012096f
C885 VTAIL.n361 B 0.028591f
C886 VTAIL.n362 B 0.012808f
C887 VTAIL.n363 B 0.02251f
C888 VTAIL.n364 B 0.012096f
C889 VTAIL.n365 B 0.028591f
C890 VTAIL.n366 B 0.012808f
C891 VTAIL.n367 B 0.02251f
C892 VTAIL.n368 B 0.012096f
C893 VTAIL.n369 B 0.028591f
C894 VTAIL.n370 B 0.012808f
C895 VTAIL.n371 B 1.93809f
C896 VTAIL.n372 B 0.012096f
C897 VTAIL.t3 B 0.047497f
C898 VTAIL.n373 B 0.172723f
C899 VTAIL.n374 B 0.016889f
C900 VTAIL.n375 B 0.021443f
C901 VTAIL.n376 B 0.028591f
C902 VTAIL.n377 B 0.012808f
C903 VTAIL.n378 B 0.012096f
C904 VTAIL.n379 B 0.02251f
C905 VTAIL.n380 B 0.02251f
C906 VTAIL.n381 B 0.012096f
C907 VTAIL.n382 B 0.012808f
C908 VTAIL.n383 B 0.028591f
C909 VTAIL.n384 B 0.028591f
C910 VTAIL.n385 B 0.012808f
C911 VTAIL.n386 B 0.012096f
C912 VTAIL.n387 B 0.02251f
C913 VTAIL.n388 B 0.02251f
C914 VTAIL.n389 B 0.012096f
C915 VTAIL.n390 B 0.012808f
C916 VTAIL.n391 B 0.028591f
C917 VTAIL.n392 B 0.028591f
C918 VTAIL.n393 B 0.012808f
C919 VTAIL.n394 B 0.012096f
C920 VTAIL.n395 B 0.02251f
C921 VTAIL.n396 B 0.02251f
C922 VTAIL.n397 B 0.012096f
C923 VTAIL.n398 B 0.012808f
C924 VTAIL.n399 B 0.028591f
C925 VTAIL.n400 B 0.028591f
C926 VTAIL.n401 B 0.012808f
C927 VTAIL.n402 B 0.012096f
C928 VTAIL.n403 B 0.02251f
C929 VTAIL.n404 B 0.02251f
C930 VTAIL.n405 B 0.012096f
C931 VTAIL.n406 B 0.012808f
C932 VTAIL.n407 B 0.028591f
C933 VTAIL.n408 B 0.028591f
C934 VTAIL.n409 B 0.012808f
C935 VTAIL.n410 B 0.012096f
C936 VTAIL.n411 B 0.02251f
C937 VTAIL.n412 B 0.02251f
C938 VTAIL.n413 B 0.012096f
C939 VTAIL.n414 B 0.012096f
C940 VTAIL.n415 B 0.012808f
C941 VTAIL.n416 B 0.028591f
C942 VTAIL.n417 B 0.028591f
C943 VTAIL.n418 B 0.028591f
C944 VTAIL.n419 B 0.012452f
C945 VTAIL.n420 B 0.012096f
C946 VTAIL.n421 B 0.02251f
C947 VTAIL.n422 B 0.02251f
C948 VTAIL.n423 B 0.012096f
C949 VTAIL.n424 B 0.012808f
C950 VTAIL.n425 B 0.028591f
C951 VTAIL.n426 B 0.028591f
C952 VTAIL.n427 B 0.012808f
C953 VTAIL.n428 B 0.012096f
C954 VTAIL.n429 B 0.02251f
C955 VTAIL.n430 B 0.02251f
C956 VTAIL.n431 B 0.012096f
C957 VTAIL.n432 B 0.012808f
C958 VTAIL.n433 B 0.028591f
C959 VTAIL.n434 B 0.028591f
C960 VTAIL.n435 B 0.012808f
C961 VTAIL.n436 B 0.012096f
C962 VTAIL.n437 B 0.02251f
C963 VTAIL.n438 B 0.02251f
C964 VTAIL.n439 B 0.012096f
C965 VTAIL.n440 B 0.012808f
C966 VTAIL.n441 B 0.028591f
C967 VTAIL.n442 B 0.061626f
C968 VTAIL.n443 B 0.012808f
C969 VTAIL.n444 B 0.012096f
C970 VTAIL.n445 B 0.049264f
C971 VTAIL.n446 B 0.034367f
C972 VTAIL.n447 B 1.92825f
C973 VP.t5 B 3.33709f
C974 VP.n0 B 1.22121f
C975 VP.n1 B 0.019445f
C976 VP.n2 B 0.015727f
C977 VP.n3 B 0.019445f
C978 VP.t4 B 3.33709f
C979 VP.n4 B 1.14951f
C980 VP.n5 B 0.019445f
C981 VP.n6 B 0.015727f
C982 VP.n7 B 0.019445f
C983 VP.t1 B 3.33709f
C984 VP.n8 B 1.22121f
C985 VP.t2 B 3.33709f
C986 VP.n9 B 1.22121f
C987 VP.n10 B 0.019445f
C988 VP.n11 B 0.015727f
C989 VP.n12 B 0.019445f
C990 VP.t3 B 3.33709f
C991 VP.n13 B 1.21332f
C992 VP.t0 B 3.56894f
C993 VP.n14 B 1.17097f
C994 VP.n15 B 0.226206f
C995 VP.n16 B 0.027295f
C996 VP.n17 B 0.036242f
C997 VP.n18 B 0.038743f
C998 VP.n19 B 0.019445f
C999 VP.n20 B 0.019445f
C1000 VP.n21 B 0.019445f
C1001 VP.n22 B 0.038548f
C1002 VP.n23 B 0.036242f
C1003 VP.n24 B 0.027653f
C1004 VP.n25 B 0.031385f
C1005 VP.n26 B 1.31997f
C1006 VP.n27 B 1.33228f
C1007 VP.n28 B 0.031385f
C1008 VP.n29 B 0.027653f
C1009 VP.n30 B 0.036242f
C1010 VP.n31 B 0.038548f
C1011 VP.n32 B 0.019445f
C1012 VP.n33 B 0.019445f
C1013 VP.n34 B 0.019445f
C1014 VP.n35 B 0.038743f
C1015 VP.n36 B 0.036242f
C1016 VP.n37 B 0.027295f
C1017 VP.n38 B 0.019445f
C1018 VP.n39 B 0.019445f
C1019 VP.n40 B 0.027295f
C1020 VP.n41 B 0.036242f
C1021 VP.n42 B 0.038743f
C1022 VP.n43 B 0.019445f
C1023 VP.n44 B 0.019445f
C1024 VP.n45 B 0.019445f
C1025 VP.n46 B 0.038548f
C1026 VP.n47 B 0.036242f
C1027 VP.n48 B 0.027653f
C1028 VP.n49 B 0.031385f
C1029 VP.n50 B 0.047504f
.ends

