* NGSPICE file created from diff_pair_sample_1619.ext - technology: sky130A

.subckt diff_pair_sample_1619 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t19 B.t5 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X1 VDD2.t9 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X2 VTAIL.t3 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X3 VTAIL.t6 VN.t2 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X4 VDD1.t8 VP.t1 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=3.3423 ps=17.92 w=8.57 l=2.14
X5 VDD2.t6 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=1.41405 ps=8.9 w=8.57 l=2.14
X6 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=0 ps=0 w=8.57 l=2.14
X7 VDD1.t7 VP.t2 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=1.41405 ps=8.9 w=8.57 l=2.14
X8 VTAIL.t16 VP.t3 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X9 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=0 ps=0 w=8.57 l=2.14
X10 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=1.41405 ps=8.9 w=8.57 l=2.14
X11 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=0 ps=0 w=8.57 l=2.14
X12 VTAIL.t8 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=0 ps=0 w=8.57 l=2.14
X14 VTAIL.t0 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X15 VTAIL.t18 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X16 VTAIL.t17 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X17 VDD2.t2 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X18 VDD2.t1 VN.t8 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=3.3423 ps=17.92 w=8.57 l=2.14
X19 VDD1.t3 VP.t6 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=3.3423 ps=17.92 w=8.57 l=2.14
X20 VTAIL.t14 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X21 VDD1.t1 VP.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=1.41405 ps=8.9 w=8.57 l=2.14
X22 VDD2.t0 VN.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.41405 pd=8.9 as=3.3423 ps=17.92 w=8.57 l=2.14
X23 VDD1.t0 VP.t9 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3423 pd=17.92 as=1.41405 ps=8.9 w=8.57 l=2.14
R0 VP.n20 VP.n19 161.3
R1 VP.n21 VP.n16 161.3
R2 VP.n23 VP.n22 161.3
R3 VP.n24 VP.n15 161.3
R4 VP.n26 VP.n25 161.3
R5 VP.n27 VP.n14 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n13 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n34 VP.n12 161.3
R10 VP.n36 VP.n35 161.3
R11 VP.n37 VP.n11 161.3
R12 VP.n39 VP.n38 161.3
R13 VP.n40 VP.n10 161.3
R14 VP.n74 VP.n0 161.3
R15 VP.n73 VP.n72 161.3
R16 VP.n71 VP.n1 161.3
R17 VP.n70 VP.n69 161.3
R18 VP.n68 VP.n2 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n3 161.3
R21 VP.n63 VP.n62 161.3
R22 VP.n61 VP.n4 161.3
R23 VP.n60 VP.n59 161.3
R24 VP.n58 VP.n5 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n6 161.3
R27 VP.n54 VP.n53 161.3
R28 VP.n52 VP.n51 161.3
R29 VP.n50 VP.n8 161.3
R30 VP.n49 VP.n48 161.3
R31 VP.n47 VP.n9 161.3
R32 VP.n46 VP.n45 161.3
R33 VP.n18 VP.t2 130.905
R34 VP.n60 VP.t8 96.5131
R35 VP.n44 VP.t9 96.5131
R36 VP.n7 VP.t4 96.5131
R37 VP.n67 VP.t7 96.5131
R38 VP.n75 VP.t1 96.5131
R39 VP.n26 VP.t0 96.5131
R40 VP.n41 VP.t6 96.5131
R41 VP.n33 VP.t3 96.5131
R42 VP.n17 VP.t5 96.5131
R43 VP.n44 VP.n43 89.2255
R44 VP.n76 VP.n75 89.2255
R45 VP.n42 VP.n41 89.2255
R46 VP.n49 VP.n9 56.5193
R47 VP.n56 VP.n55 56.5193
R48 VP.n62 VP.n3 56.5193
R49 VP.n73 VP.n1 56.5193
R50 VP.n39 VP.n11 56.5193
R51 VP.n28 VP.n13 56.5193
R52 VP.n22 VP.n21 56.5193
R53 VP.n43 VP.n42 48.1019
R54 VP.n18 VP.n17 47.6808
R55 VP.n45 VP.n9 24.4675
R56 VP.n50 VP.n49 24.4675
R57 VP.n51 VP.n50 24.4675
R58 VP.n55 VP.n54 24.4675
R59 VP.n56 VP.n5 24.4675
R60 VP.n60 VP.n5 24.4675
R61 VP.n61 VP.n60 24.4675
R62 VP.n62 VP.n61 24.4675
R63 VP.n66 VP.n3 24.4675
R64 VP.n69 VP.n68 24.4675
R65 VP.n69 VP.n1 24.4675
R66 VP.n74 VP.n73 24.4675
R67 VP.n40 VP.n39 24.4675
R68 VP.n32 VP.n13 24.4675
R69 VP.n35 VP.n34 24.4675
R70 VP.n35 VP.n11 24.4675
R71 VP.n22 VP.n15 24.4675
R72 VP.n26 VP.n15 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 22.9995
R77 VP.n67 VP.n66 22.9995
R78 VP.n33 VP.n32 22.9995
R79 VP.n20 VP.n17 22.9995
R80 VP.n45 VP.n44 21.5315
R81 VP.n75 VP.n74 21.5315
R82 VP.n41 VP.n40 21.5315
R83 VP.n19 VP.n18 8.82758
R84 VP.n51 VP.n7 1.46852
R85 VP.n68 VP.n67 1.46852
R86 VP.n34 VP.n33 1.46852
R87 VP.n42 VP.n10 0.278367
R88 VP.n46 VP.n43 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153454
R122 VTAIL.n192 VTAIL.n152 289.615
R123 VTAIL.n42 VTAIL.n2 289.615
R124 VTAIL.n146 VTAIL.n106 289.615
R125 VTAIL.n96 VTAIL.n56 289.615
R126 VTAIL.n167 VTAIL.n166 185
R127 VTAIL.n164 VTAIL.n163 185
R128 VTAIL.n173 VTAIL.n172 185
R129 VTAIL.n175 VTAIL.n174 185
R130 VTAIL.n160 VTAIL.n159 185
R131 VTAIL.n181 VTAIL.n180 185
R132 VTAIL.n184 VTAIL.n183 185
R133 VTAIL.n182 VTAIL.n156 185
R134 VTAIL.n189 VTAIL.n155 185
R135 VTAIL.n191 VTAIL.n190 185
R136 VTAIL.n193 VTAIL.n192 185
R137 VTAIL.n17 VTAIL.n16 185
R138 VTAIL.n14 VTAIL.n13 185
R139 VTAIL.n23 VTAIL.n22 185
R140 VTAIL.n25 VTAIL.n24 185
R141 VTAIL.n10 VTAIL.n9 185
R142 VTAIL.n31 VTAIL.n30 185
R143 VTAIL.n34 VTAIL.n33 185
R144 VTAIL.n32 VTAIL.n6 185
R145 VTAIL.n39 VTAIL.n5 185
R146 VTAIL.n41 VTAIL.n40 185
R147 VTAIL.n43 VTAIL.n42 185
R148 VTAIL.n147 VTAIL.n146 185
R149 VTAIL.n145 VTAIL.n144 185
R150 VTAIL.n143 VTAIL.n109 185
R151 VTAIL.n113 VTAIL.n110 185
R152 VTAIL.n138 VTAIL.n137 185
R153 VTAIL.n136 VTAIL.n135 185
R154 VTAIL.n115 VTAIL.n114 185
R155 VTAIL.n130 VTAIL.n129 185
R156 VTAIL.n128 VTAIL.n127 185
R157 VTAIL.n119 VTAIL.n118 185
R158 VTAIL.n122 VTAIL.n121 185
R159 VTAIL.n97 VTAIL.n96 185
R160 VTAIL.n95 VTAIL.n94 185
R161 VTAIL.n93 VTAIL.n59 185
R162 VTAIL.n63 VTAIL.n60 185
R163 VTAIL.n88 VTAIL.n87 185
R164 VTAIL.n86 VTAIL.n85 185
R165 VTAIL.n65 VTAIL.n64 185
R166 VTAIL.n80 VTAIL.n79 185
R167 VTAIL.n78 VTAIL.n77 185
R168 VTAIL.n69 VTAIL.n68 185
R169 VTAIL.n72 VTAIL.n71 185
R170 VTAIL.t7 VTAIL.n165 149.524
R171 VTAIL.t12 VTAIL.n15 149.524
R172 VTAIL.t13 VTAIL.n120 149.524
R173 VTAIL.t9 VTAIL.n70 149.524
R174 VTAIL.n166 VTAIL.n163 104.615
R175 VTAIL.n173 VTAIL.n163 104.615
R176 VTAIL.n174 VTAIL.n173 104.615
R177 VTAIL.n174 VTAIL.n159 104.615
R178 VTAIL.n181 VTAIL.n159 104.615
R179 VTAIL.n183 VTAIL.n181 104.615
R180 VTAIL.n183 VTAIL.n182 104.615
R181 VTAIL.n182 VTAIL.n155 104.615
R182 VTAIL.n191 VTAIL.n155 104.615
R183 VTAIL.n192 VTAIL.n191 104.615
R184 VTAIL.n16 VTAIL.n13 104.615
R185 VTAIL.n23 VTAIL.n13 104.615
R186 VTAIL.n24 VTAIL.n23 104.615
R187 VTAIL.n24 VTAIL.n9 104.615
R188 VTAIL.n31 VTAIL.n9 104.615
R189 VTAIL.n33 VTAIL.n31 104.615
R190 VTAIL.n33 VTAIL.n32 104.615
R191 VTAIL.n32 VTAIL.n5 104.615
R192 VTAIL.n41 VTAIL.n5 104.615
R193 VTAIL.n42 VTAIL.n41 104.615
R194 VTAIL.n146 VTAIL.n145 104.615
R195 VTAIL.n145 VTAIL.n109 104.615
R196 VTAIL.n113 VTAIL.n109 104.615
R197 VTAIL.n137 VTAIL.n113 104.615
R198 VTAIL.n137 VTAIL.n136 104.615
R199 VTAIL.n136 VTAIL.n114 104.615
R200 VTAIL.n129 VTAIL.n114 104.615
R201 VTAIL.n129 VTAIL.n128 104.615
R202 VTAIL.n128 VTAIL.n118 104.615
R203 VTAIL.n121 VTAIL.n118 104.615
R204 VTAIL.n96 VTAIL.n95 104.615
R205 VTAIL.n95 VTAIL.n59 104.615
R206 VTAIL.n63 VTAIL.n59 104.615
R207 VTAIL.n87 VTAIL.n63 104.615
R208 VTAIL.n87 VTAIL.n86 104.615
R209 VTAIL.n86 VTAIL.n64 104.615
R210 VTAIL.n79 VTAIL.n64 104.615
R211 VTAIL.n79 VTAIL.n78 104.615
R212 VTAIL.n78 VTAIL.n68 104.615
R213 VTAIL.n71 VTAIL.n68 104.615
R214 VTAIL.n166 VTAIL.t7 52.3082
R215 VTAIL.n16 VTAIL.t12 52.3082
R216 VTAIL.n121 VTAIL.t13 52.3082
R217 VTAIL.n71 VTAIL.t9 52.3082
R218 VTAIL.n105 VTAIL.n104 47.7321
R219 VTAIL.n103 VTAIL.n102 47.7321
R220 VTAIL.n55 VTAIL.n54 47.7321
R221 VTAIL.n53 VTAIL.n52 47.7321
R222 VTAIL.n199 VTAIL.n198 47.7319
R223 VTAIL.n1 VTAIL.n0 47.7319
R224 VTAIL.n49 VTAIL.n48 47.7319
R225 VTAIL.n51 VTAIL.n50 47.7319
R226 VTAIL.n197 VTAIL.n196 33.155
R227 VTAIL.n47 VTAIL.n46 33.155
R228 VTAIL.n151 VTAIL.n150 33.155
R229 VTAIL.n101 VTAIL.n100 33.155
R230 VTAIL.n53 VTAIL.n51 24.0134
R231 VTAIL.n197 VTAIL.n151 21.8841
R232 VTAIL.n190 VTAIL.n189 13.1884
R233 VTAIL.n40 VTAIL.n39 13.1884
R234 VTAIL.n144 VTAIL.n143 13.1884
R235 VTAIL.n94 VTAIL.n93 13.1884
R236 VTAIL.n188 VTAIL.n156 12.8005
R237 VTAIL.n193 VTAIL.n154 12.8005
R238 VTAIL.n38 VTAIL.n6 12.8005
R239 VTAIL.n43 VTAIL.n4 12.8005
R240 VTAIL.n147 VTAIL.n108 12.8005
R241 VTAIL.n142 VTAIL.n110 12.8005
R242 VTAIL.n97 VTAIL.n58 12.8005
R243 VTAIL.n92 VTAIL.n60 12.8005
R244 VTAIL.n185 VTAIL.n184 12.0247
R245 VTAIL.n194 VTAIL.n152 12.0247
R246 VTAIL.n35 VTAIL.n34 12.0247
R247 VTAIL.n44 VTAIL.n2 12.0247
R248 VTAIL.n148 VTAIL.n106 12.0247
R249 VTAIL.n139 VTAIL.n138 12.0247
R250 VTAIL.n98 VTAIL.n56 12.0247
R251 VTAIL.n89 VTAIL.n88 12.0247
R252 VTAIL.n180 VTAIL.n158 11.249
R253 VTAIL.n30 VTAIL.n8 11.249
R254 VTAIL.n135 VTAIL.n112 11.249
R255 VTAIL.n85 VTAIL.n62 11.249
R256 VTAIL.n179 VTAIL.n160 10.4732
R257 VTAIL.n29 VTAIL.n10 10.4732
R258 VTAIL.n134 VTAIL.n115 10.4732
R259 VTAIL.n84 VTAIL.n65 10.4732
R260 VTAIL.n167 VTAIL.n165 10.2747
R261 VTAIL.n17 VTAIL.n15 10.2747
R262 VTAIL.n122 VTAIL.n120 10.2747
R263 VTAIL.n72 VTAIL.n70 10.2747
R264 VTAIL.n176 VTAIL.n175 9.69747
R265 VTAIL.n26 VTAIL.n25 9.69747
R266 VTAIL.n131 VTAIL.n130 9.69747
R267 VTAIL.n81 VTAIL.n80 9.69747
R268 VTAIL.n196 VTAIL.n195 9.45567
R269 VTAIL.n46 VTAIL.n45 9.45567
R270 VTAIL.n150 VTAIL.n149 9.45567
R271 VTAIL.n100 VTAIL.n99 9.45567
R272 VTAIL.n195 VTAIL.n194 9.3005
R273 VTAIL.n154 VTAIL.n153 9.3005
R274 VTAIL.n169 VTAIL.n168 9.3005
R275 VTAIL.n171 VTAIL.n170 9.3005
R276 VTAIL.n162 VTAIL.n161 9.3005
R277 VTAIL.n177 VTAIL.n176 9.3005
R278 VTAIL.n179 VTAIL.n178 9.3005
R279 VTAIL.n158 VTAIL.n157 9.3005
R280 VTAIL.n186 VTAIL.n185 9.3005
R281 VTAIL.n188 VTAIL.n187 9.3005
R282 VTAIL.n45 VTAIL.n44 9.3005
R283 VTAIL.n4 VTAIL.n3 9.3005
R284 VTAIL.n19 VTAIL.n18 9.3005
R285 VTAIL.n21 VTAIL.n20 9.3005
R286 VTAIL.n12 VTAIL.n11 9.3005
R287 VTAIL.n27 VTAIL.n26 9.3005
R288 VTAIL.n29 VTAIL.n28 9.3005
R289 VTAIL.n8 VTAIL.n7 9.3005
R290 VTAIL.n36 VTAIL.n35 9.3005
R291 VTAIL.n38 VTAIL.n37 9.3005
R292 VTAIL.n124 VTAIL.n123 9.3005
R293 VTAIL.n126 VTAIL.n125 9.3005
R294 VTAIL.n117 VTAIL.n116 9.3005
R295 VTAIL.n132 VTAIL.n131 9.3005
R296 VTAIL.n134 VTAIL.n133 9.3005
R297 VTAIL.n112 VTAIL.n111 9.3005
R298 VTAIL.n140 VTAIL.n139 9.3005
R299 VTAIL.n142 VTAIL.n141 9.3005
R300 VTAIL.n149 VTAIL.n148 9.3005
R301 VTAIL.n108 VTAIL.n107 9.3005
R302 VTAIL.n74 VTAIL.n73 9.3005
R303 VTAIL.n76 VTAIL.n75 9.3005
R304 VTAIL.n67 VTAIL.n66 9.3005
R305 VTAIL.n82 VTAIL.n81 9.3005
R306 VTAIL.n84 VTAIL.n83 9.3005
R307 VTAIL.n62 VTAIL.n61 9.3005
R308 VTAIL.n90 VTAIL.n89 9.3005
R309 VTAIL.n92 VTAIL.n91 9.3005
R310 VTAIL.n99 VTAIL.n98 9.3005
R311 VTAIL.n58 VTAIL.n57 9.3005
R312 VTAIL.n172 VTAIL.n162 8.92171
R313 VTAIL.n22 VTAIL.n12 8.92171
R314 VTAIL.n127 VTAIL.n117 8.92171
R315 VTAIL.n77 VTAIL.n67 8.92171
R316 VTAIL.n171 VTAIL.n164 8.14595
R317 VTAIL.n21 VTAIL.n14 8.14595
R318 VTAIL.n126 VTAIL.n119 8.14595
R319 VTAIL.n76 VTAIL.n69 8.14595
R320 VTAIL.n168 VTAIL.n167 7.3702
R321 VTAIL.n18 VTAIL.n17 7.3702
R322 VTAIL.n123 VTAIL.n122 7.3702
R323 VTAIL.n73 VTAIL.n72 7.3702
R324 VTAIL.n168 VTAIL.n164 5.81868
R325 VTAIL.n18 VTAIL.n14 5.81868
R326 VTAIL.n123 VTAIL.n119 5.81868
R327 VTAIL.n73 VTAIL.n69 5.81868
R328 VTAIL.n172 VTAIL.n171 5.04292
R329 VTAIL.n22 VTAIL.n21 5.04292
R330 VTAIL.n127 VTAIL.n126 5.04292
R331 VTAIL.n77 VTAIL.n76 5.04292
R332 VTAIL.n175 VTAIL.n162 4.26717
R333 VTAIL.n25 VTAIL.n12 4.26717
R334 VTAIL.n130 VTAIL.n117 4.26717
R335 VTAIL.n80 VTAIL.n67 4.26717
R336 VTAIL.n176 VTAIL.n160 3.49141
R337 VTAIL.n26 VTAIL.n10 3.49141
R338 VTAIL.n131 VTAIL.n115 3.49141
R339 VTAIL.n81 VTAIL.n65 3.49141
R340 VTAIL.n169 VTAIL.n165 2.84303
R341 VTAIL.n19 VTAIL.n15 2.84303
R342 VTAIL.n124 VTAIL.n120 2.84303
R343 VTAIL.n74 VTAIL.n70 2.84303
R344 VTAIL.n180 VTAIL.n179 2.71565
R345 VTAIL.n30 VTAIL.n29 2.71565
R346 VTAIL.n135 VTAIL.n134 2.71565
R347 VTAIL.n85 VTAIL.n84 2.71565
R348 VTAIL.n198 VTAIL.t5 2.31088
R349 VTAIL.n198 VTAIL.t8 2.31088
R350 VTAIL.n0 VTAIL.t2 2.31088
R351 VTAIL.n0 VTAIL.t0 2.31088
R352 VTAIL.n48 VTAIL.t11 2.31088
R353 VTAIL.n48 VTAIL.t14 2.31088
R354 VTAIL.n50 VTAIL.t15 2.31088
R355 VTAIL.n50 VTAIL.t18 2.31088
R356 VTAIL.n104 VTAIL.t19 2.31088
R357 VTAIL.n104 VTAIL.t16 2.31088
R358 VTAIL.n102 VTAIL.t10 2.31088
R359 VTAIL.n102 VTAIL.t17 2.31088
R360 VTAIL.n54 VTAIL.t4 2.31088
R361 VTAIL.n54 VTAIL.t3 2.31088
R362 VTAIL.n52 VTAIL.t1 2.31088
R363 VTAIL.n52 VTAIL.t6 2.31088
R364 VTAIL.n55 VTAIL.n53 2.12981
R365 VTAIL.n101 VTAIL.n55 2.12981
R366 VTAIL.n105 VTAIL.n103 2.12981
R367 VTAIL.n151 VTAIL.n105 2.12981
R368 VTAIL.n51 VTAIL.n49 2.12981
R369 VTAIL.n49 VTAIL.n47 2.12981
R370 VTAIL.n199 VTAIL.n197 2.12981
R371 VTAIL.n184 VTAIL.n158 1.93989
R372 VTAIL.n196 VTAIL.n152 1.93989
R373 VTAIL.n34 VTAIL.n8 1.93989
R374 VTAIL.n46 VTAIL.n2 1.93989
R375 VTAIL.n150 VTAIL.n106 1.93989
R376 VTAIL.n138 VTAIL.n112 1.93989
R377 VTAIL.n100 VTAIL.n56 1.93989
R378 VTAIL.n88 VTAIL.n62 1.93989
R379 VTAIL VTAIL.n1 1.65567
R380 VTAIL.n103 VTAIL.n101 1.53498
R381 VTAIL.n47 VTAIL.n1 1.53498
R382 VTAIL.n185 VTAIL.n156 1.16414
R383 VTAIL.n194 VTAIL.n193 1.16414
R384 VTAIL.n35 VTAIL.n6 1.16414
R385 VTAIL.n44 VTAIL.n43 1.16414
R386 VTAIL.n148 VTAIL.n147 1.16414
R387 VTAIL.n139 VTAIL.n110 1.16414
R388 VTAIL.n98 VTAIL.n97 1.16414
R389 VTAIL.n89 VTAIL.n60 1.16414
R390 VTAIL VTAIL.n199 0.474638
R391 VTAIL.n189 VTAIL.n188 0.388379
R392 VTAIL.n190 VTAIL.n154 0.388379
R393 VTAIL.n39 VTAIL.n38 0.388379
R394 VTAIL.n40 VTAIL.n4 0.388379
R395 VTAIL.n144 VTAIL.n108 0.388379
R396 VTAIL.n143 VTAIL.n142 0.388379
R397 VTAIL.n94 VTAIL.n58 0.388379
R398 VTAIL.n93 VTAIL.n92 0.388379
R399 VTAIL.n170 VTAIL.n169 0.155672
R400 VTAIL.n170 VTAIL.n161 0.155672
R401 VTAIL.n177 VTAIL.n161 0.155672
R402 VTAIL.n178 VTAIL.n177 0.155672
R403 VTAIL.n178 VTAIL.n157 0.155672
R404 VTAIL.n186 VTAIL.n157 0.155672
R405 VTAIL.n187 VTAIL.n186 0.155672
R406 VTAIL.n187 VTAIL.n153 0.155672
R407 VTAIL.n195 VTAIL.n153 0.155672
R408 VTAIL.n20 VTAIL.n19 0.155672
R409 VTAIL.n20 VTAIL.n11 0.155672
R410 VTAIL.n27 VTAIL.n11 0.155672
R411 VTAIL.n28 VTAIL.n27 0.155672
R412 VTAIL.n28 VTAIL.n7 0.155672
R413 VTAIL.n36 VTAIL.n7 0.155672
R414 VTAIL.n37 VTAIL.n36 0.155672
R415 VTAIL.n37 VTAIL.n3 0.155672
R416 VTAIL.n45 VTAIL.n3 0.155672
R417 VTAIL.n149 VTAIL.n107 0.155672
R418 VTAIL.n141 VTAIL.n107 0.155672
R419 VTAIL.n141 VTAIL.n140 0.155672
R420 VTAIL.n140 VTAIL.n111 0.155672
R421 VTAIL.n133 VTAIL.n111 0.155672
R422 VTAIL.n133 VTAIL.n132 0.155672
R423 VTAIL.n132 VTAIL.n116 0.155672
R424 VTAIL.n125 VTAIL.n116 0.155672
R425 VTAIL.n125 VTAIL.n124 0.155672
R426 VTAIL.n99 VTAIL.n57 0.155672
R427 VTAIL.n91 VTAIL.n57 0.155672
R428 VTAIL.n91 VTAIL.n90 0.155672
R429 VTAIL.n90 VTAIL.n61 0.155672
R430 VTAIL.n83 VTAIL.n61 0.155672
R431 VTAIL.n83 VTAIL.n82 0.155672
R432 VTAIL.n82 VTAIL.n66 0.155672
R433 VTAIL.n75 VTAIL.n66 0.155672
R434 VTAIL.n75 VTAIL.n74 0.155672
R435 VDD1.n40 VDD1.n0 289.615
R436 VDD1.n87 VDD1.n47 289.615
R437 VDD1.n41 VDD1.n40 185
R438 VDD1.n39 VDD1.n38 185
R439 VDD1.n37 VDD1.n3 185
R440 VDD1.n7 VDD1.n4 185
R441 VDD1.n32 VDD1.n31 185
R442 VDD1.n30 VDD1.n29 185
R443 VDD1.n9 VDD1.n8 185
R444 VDD1.n24 VDD1.n23 185
R445 VDD1.n22 VDD1.n21 185
R446 VDD1.n13 VDD1.n12 185
R447 VDD1.n16 VDD1.n15 185
R448 VDD1.n62 VDD1.n61 185
R449 VDD1.n59 VDD1.n58 185
R450 VDD1.n68 VDD1.n67 185
R451 VDD1.n70 VDD1.n69 185
R452 VDD1.n55 VDD1.n54 185
R453 VDD1.n76 VDD1.n75 185
R454 VDD1.n79 VDD1.n78 185
R455 VDD1.n77 VDD1.n51 185
R456 VDD1.n84 VDD1.n50 185
R457 VDD1.n86 VDD1.n85 185
R458 VDD1.n88 VDD1.n87 185
R459 VDD1.t7 VDD1.n14 149.524
R460 VDD1.t0 VDD1.n60 149.524
R461 VDD1.n40 VDD1.n39 104.615
R462 VDD1.n39 VDD1.n3 104.615
R463 VDD1.n7 VDD1.n3 104.615
R464 VDD1.n31 VDD1.n7 104.615
R465 VDD1.n31 VDD1.n30 104.615
R466 VDD1.n30 VDD1.n8 104.615
R467 VDD1.n23 VDD1.n8 104.615
R468 VDD1.n23 VDD1.n22 104.615
R469 VDD1.n22 VDD1.n12 104.615
R470 VDD1.n15 VDD1.n12 104.615
R471 VDD1.n61 VDD1.n58 104.615
R472 VDD1.n68 VDD1.n58 104.615
R473 VDD1.n69 VDD1.n68 104.615
R474 VDD1.n69 VDD1.n54 104.615
R475 VDD1.n76 VDD1.n54 104.615
R476 VDD1.n78 VDD1.n76 104.615
R477 VDD1.n78 VDD1.n77 104.615
R478 VDD1.n77 VDD1.n50 104.615
R479 VDD1.n86 VDD1.n50 104.615
R480 VDD1.n87 VDD1.n86 104.615
R481 VDD1.n95 VDD1.n94 65.9523
R482 VDD1.n46 VDD1.n45 64.4109
R483 VDD1.n97 VDD1.n96 64.4107
R484 VDD1.n93 VDD1.n92 64.4107
R485 VDD1.n15 VDD1.t7 52.3082
R486 VDD1.n61 VDD1.t0 52.3082
R487 VDD1.n46 VDD1.n44 51.9631
R488 VDD1.n93 VDD1.n91 51.9631
R489 VDD1.n97 VDD1.n95 42.8651
R490 VDD1.n38 VDD1.n37 13.1884
R491 VDD1.n85 VDD1.n84 13.1884
R492 VDD1.n41 VDD1.n2 12.8005
R493 VDD1.n36 VDD1.n4 12.8005
R494 VDD1.n83 VDD1.n51 12.8005
R495 VDD1.n88 VDD1.n49 12.8005
R496 VDD1.n42 VDD1.n0 12.0247
R497 VDD1.n33 VDD1.n32 12.0247
R498 VDD1.n80 VDD1.n79 12.0247
R499 VDD1.n89 VDD1.n47 12.0247
R500 VDD1.n29 VDD1.n6 11.249
R501 VDD1.n75 VDD1.n53 11.249
R502 VDD1.n28 VDD1.n9 10.4732
R503 VDD1.n74 VDD1.n55 10.4732
R504 VDD1.n16 VDD1.n14 10.2747
R505 VDD1.n62 VDD1.n60 10.2747
R506 VDD1.n25 VDD1.n24 9.69747
R507 VDD1.n71 VDD1.n70 9.69747
R508 VDD1.n44 VDD1.n43 9.45567
R509 VDD1.n91 VDD1.n90 9.45567
R510 VDD1.n18 VDD1.n17 9.3005
R511 VDD1.n20 VDD1.n19 9.3005
R512 VDD1.n11 VDD1.n10 9.3005
R513 VDD1.n26 VDD1.n25 9.3005
R514 VDD1.n28 VDD1.n27 9.3005
R515 VDD1.n6 VDD1.n5 9.3005
R516 VDD1.n34 VDD1.n33 9.3005
R517 VDD1.n36 VDD1.n35 9.3005
R518 VDD1.n43 VDD1.n42 9.3005
R519 VDD1.n2 VDD1.n1 9.3005
R520 VDD1.n90 VDD1.n89 9.3005
R521 VDD1.n49 VDD1.n48 9.3005
R522 VDD1.n64 VDD1.n63 9.3005
R523 VDD1.n66 VDD1.n65 9.3005
R524 VDD1.n57 VDD1.n56 9.3005
R525 VDD1.n72 VDD1.n71 9.3005
R526 VDD1.n74 VDD1.n73 9.3005
R527 VDD1.n53 VDD1.n52 9.3005
R528 VDD1.n81 VDD1.n80 9.3005
R529 VDD1.n83 VDD1.n82 9.3005
R530 VDD1.n21 VDD1.n11 8.92171
R531 VDD1.n67 VDD1.n57 8.92171
R532 VDD1.n20 VDD1.n13 8.14595
R533 VDD1.n66 VDD1.n59 8.14595
R534 VDD1.n17 VDD1.n16 7.3702
R535 VDD1.n63 VDD1.n62 7.3702
R536 VDD1.n17 VDD1.n13 5.81868
R537 VDD1.n63 VDD1.n59 5.81868
R538 VDD1.n21 VDD1.n20 5.04292
R539 VDD1.n67 VDD1.n66 5.04292
R540 VDD1.n24 VDD1.n11 4.26717
R541 VDD1.n70 VDD1.n57 4.26717
R542 VDD1.n25 VDD1.n9 3.49141
R543 VDD1.n71 VDD1.n55 3.49141
R544 VDD1.n64 VDD1.n60 2.84303
R545 VDD1.n18 VDD1.n14 2.84303
R546 VDD1.n29 VDD1.n28 2.71565
R547 VDD1.n75 VDD1.n74 2.71565
R548 VDD1.n96 VDD1.t6 2.31088
R549 VDD1.n96 VDD1.t3 2.31088
R550 VDD1.n45 VDD1.t4 2.31088
R551 VDD1.n45 VDD1.t9 2.31088
R552 VDD1.n94 VDD1.t2 2.31088
R553 VDD1.n94 VDD1.t8 2.31088
R554 VDD1.n92 VDD1.t5 2.31088
R555 VDD1.n92 VDD1.t1 2.31088
R556 VDD1.n44 VDD1.n0 1.93989
R557 VDD1.n32 VDD1.n6 1.93989
R558 VDD1.n79 VDD1.n53 1.93989
R559 VDD1.n91 VDD1.n47 1.93989
R560 VDD1 VDD1.n97 1.53929
R561 VDD1.n42 VDD1.n41 1.16414
R562 VDD1.n33 VDD1.n4 1.16414
R563 VDD1.n80 VDD1.n51 1.16414
R564 VDD1.n89 VDD1.n88 1.16414
R565 VDD1 VDD1.n46 0.591017
R566 VDD1.n95 VDD1.n93 0.477482
R567 VDD1.n38 VDD1.n2 0.388379
R568 VDD1.n37 VDD1.n36 0.388379
R569 VDD1.n84 VDD1.n83 0.388379
R570 VDD1.n85 VDD1.n49 0.388379
R571 VDD1.n43 VDD1.n1 0.155672
R572 VDD1.n35 VDD1.n1 0.155672
R573 VDD1.n35 VDD1.n34 0.155672
R574 VDD1.n34 VDD1.n5 0.155672
R575 VDD1.n27 VDD1.n5 0.155672
R576 VDD1.n27 VDD1.n26 0.155672
R577 VDD1.n26 VDD1.n10 0.155672
R578 VDD1.n19 VDD1.n10 0.155672
R579 VDD1.n19 VDD1.n18 0.155672
R580 VDD1.n65 VDD1.n64 0.155672
R581 VDD1.n65 VDD1.n56 0.155672
R582 VDD1.n72 VDD1.n56 0.155672
R583 VDD1.n73 VDD1.n72 0.155672
R584 VDD1.n73 VDD1.n52 0.155672
R585 VDD1.n81 VDD1.n52 0.155672
R586 VDD1.n82 VDD1.n81 0.155672
R587 VDD1.n82 VDD1.n48 0.155672
R588 VDD1.n90 VDD1.n48 0.155672
R589 B.n786 B.n785 585
R590 B.n787 B.n786 585
R591 B.n278 B.n132 585
R592 B.n277 B.n276 585
R593 B.n275 B.n274 585
R594 B.n273 B.n272 585
R595 B.n271 B.n270 585
R596 B.n269 B.n268 585
R597 B.n267 B.n266 585
R598 B.n265 B.n264 585
R599 B.n263 B.n262 585
R600 B.n261 B.n260 585
R601 B.n259 B.n258 585
R602 B.n257 B.n256 585
R603 B.n255 B.n254 585
R604 B.n253 B.n252 585
R605 B.n251 B.n250 585
R606 B.n249 B.n248 585
R607 B.n247 B.n246 585
R608 B.n245 B.n244 585
R609 B.n243 B.n242 585
R610 B.n241 B.n240 585
R611 B.n239 B.n238 585
R612 B.n237 B.n236 585
R613 B.n235 B.n234 585
R614 B.n233 B.n232 585
R615 B.n231 B.n230 585
R616 B.n229 B.n228 585
R617 B.n227 B.n226 585
R618 B.n225 B.n224 585
R619 B.n223 B.n222 585
R620 B.n221 B.n220 585
R621 B.n219 B.n218 585
R622 B.n216 B.n215 585
R623 B.n214 B.n213 585
R624 B.n212 B.n211 585
R625 B.n210 B.n209 585
R626 B.n208 B.n207 585
R627 B.n206 B.n205 585
R628 B.n204 B.n203 585
R629 B.n202 B.n201 585
R630 B.n200 B.n199 585
R631 B.n198 B.n197 585
R632 B.n196 B.n195 585
R633 B.n194 B.n193 585
R634 B.n192 B.n191 585
R635 B.n190 B.n189 585
R636 B.n188 B.n187 585
R637 B.n186 B.n185 585
R638 B.n184 B.n183 585
R639 B.n182 B.n181 585
R640 B.n180 B.n179 585
R641 B.n178 B.n177 585
R642 B.n176 B.n175 585
R643 B.n174 B.n173 585
R644 B.n172 B.n171 585
R645 B.n170 B.n169 585
R646 B.n168 B.n167 585
R647 B.n166 B.n165 585
R648 B.n164 B.n163 585
R649 B.n162 B.n161 585
R650 B.n160 B.n159 585
R651 B.n158 B.n157 585
R652 B.n156 B.n155 585
R653 B.n154 B.n153 585
R654 B.n152 B.n151 585
R655 B.n150 B.n149 585
R656 B.n148 B.n147 585
R657 B.n146 B.n145 585
R658 B.n144 B.n143 585
R659 B.n142 B.n141 585
R660 B.n140 B.n139 585
R661 B.n96 B.n95 585
R662 B.n790 B.n789 585
R663 B.n784 B.n133 585
R664 B.n133 B.n93 585
R665 B.n783 B.n92 585
R666 B.n794 B.n92 585
R667 B.n782 B.n91 585
R668 B.n795 B.n91 585
R669 B.n781 B.n90 585
R670 B.n796 B.n90 585
R671 B.n780 B.n779 585
R672 B.n779 B.n86 585
R673 B.n778 B.n85 585
R674 B.n802 B.n85 585
R675 B.n777 B.n84 585
R676 B.n803 B.n84 585
R677 B.n776 B.n83 585
R678 B.n804 B.n83 585
R679 B.n775 B.n774 585
R680 B.n774 B.n79 585
R681 B.n773 B.n78 585
R682 B.n810 B.n78 585
R683 B.n772 B.n77 585
R684 B.n811 B.n77 585
R685 B.n771 B.n76 585
R686 B.n812 B.n76 585
R687 B.n770 B.n769 585
R688 B.n769 B.n72 585
R689 B.n768 B.n71 585
R690 B.n818 B.n71 585
R691 B.n767 B.n70 585
R692 B.n819 B.n70 585
R693 B.n766 B.n69 585
R694 B.n820 B.n69 585
R695 B.n765 B.n764 585
R696 B.n764 B.n65 585
R697 B.n763 B.n64 585
R698 B.n826 B.n64 585
R699 B.n762 B.n63 585
R700 B.n827 B.n63 585
R701 B.n761 B.n62 585
R702 B.n828 B.n62 585
R703 B.n760 B.n759 585
R704 B.n759 B.n58 585
R705 B.n758 B.n57 585
R706 B.n834 B.n57 585
R707 B.n757 B.n56 585
R708 B.n835 B.n56 585
R709 B.n756 B.n55 585
R710 B.n836 B.n55 585
R711 B.n755 B.n754 585
R712 B.n754 B.n54 585
R713 B.n753 B.n50 585
R714 B.n842 B.n50 585
R715 B.n752 B.n49 585
R716 B.n843 B.n49 585
R717 B.n751 B.n48 585
R718 B.n844 B.n48 585
R719 B.n750 B.n749 585
R720 B.n749 B.n44 585
R721 B.n748 B.n43 585
R722 B.n850 B.n43 585
R723 B.n747 B.n42 585
R724 B.n851 B.n42 585
R725 B.n746 B.n41 585
R726 B.n852 B.n41 585
R727 B.n745 B.n744 585
R728 B.n744 B.n37 585
R729 B.n743 B.n36 585
R730 B.n858 B.n36 585
R731 B.n742 B.n35 585
R732 B.n859 B.n35 585
R733 B.n741 B.n34 585
R734 B.n860 B.n34 585
R735 B.n740 B.n739 585
R736 B.n739 B.n30 585
R737 B.n738 B.n29 585
R738 B.n866 B.n29 585
R739 B.n737 B.n28 585
R740 B.n867 B.n28 585
R741 B.n736 B.n27 585
R742 B.t0 B.n27 585
R743 B.n735 B.n734 585
R744 B.n734 B.n23 585
R745 B.n733 B.n22 585
R746 B.n873 B.n22 585
R747 B.n732 B.n21 585
R748 B.n874 B.n21 585
R749 B.n731 B.n20 585
R750 B.n875 B.n20 585
R751 B.n730 B.n729 585
R752 B.n729 B.n16 585
R753 B.n728 B.n15 585
R754 B.n881 B.n15 585
R755 B.n727 B.n14 585
R756 B.n882 B.n14 585
R757 B.n726 B.n13 585
R758 B.n883 B.n13 585
R759 B.n725 B.n724 585
R760 B.n724 B.n12 585
R761 B.n723 B.n722 585
R762 B.n723 B.n8 585
R763 B.n721 B.n7 585
R764 B.n890 B.n7 585
R765 B.n720 B.n6 585
R766 B.n891 B.n6 585
R767 B.n719 B.n5 585
R768 B.n892 B.n5 585
R769 B.n718 B.n717 585
R770 B.n717 B.n4 585
R771 B.n716 B.n279 585
R772 B.n716 B.n715 585
R773 B.n706 B.n280 585
R774 B.n281 B.n280 585
R775 B.n708 B.n707 585
R776 B.n709 B.n708 585
R777 B.n705 B.n285 585
R778 B.n289 B.n285 585
R779 B.n704 B.n703 585
R780 B.n703 B.n702 585
R781 B.n287 B.n286 585
R782 B.n288 B.n287 585
R783 B.n695 B.n694 585
R784 B.n696 B.n695 585
R785 B.n693 B.n294 585
R786 B.n294 B.n293 585
R787 B.n692 B.n691 585
R788 B.n691 B.n690 585
R789 B.n296 B.n295 585
R790 B.n297 B.n296 585
R791 B.n684 B.n683 585
R792 B.t3 B.n684 585
R793 B.n682 B.n302 585
R794 B.n302 B.n301 585
R795 B.n681 B.n680 585
R796 B.n680 B.n679 585
R797 B.n304 B.n303 585
R798 B.n305 B.n304 585
R799 B.n672 B.n671 585
R800 B.n673 B.n672 585
R801 B.n670 B.n310 585
R802 B.n310 B.n309 585
R803 B.n669 B.n668 585
R804 B.n668 B.n667 585
R805 B.n312 B.n311 585
R806 B.n313 B.n312 585
R807 B.n660 B.n659 585
R808 B.n661 B.n660 585
R809 B.n658 B.n318 585
R810 B.n318 B.n317 585
R811 B.n657 B.n656 585
R812 B.n656 B.n655 585
R813 B.n320 B.n319 585
R814 B.n321 B.n320 585
R815 B.n648 B.n647 585
R816 B.n649 B.n648 585
R817 B.n646 B.n326 585
R818 B.n326 B.n325 585
R819 B.n645 B.n644 585
R820 B.n644 B.n643 585
R821 B.n328 B.n327 585
R822 B.n636 B.n328 585
R823 B.n635 B.n634 585
R824 B.n637 B.n635 585
R825 B.n633 B.n333 585
R826 B.n333 B.n332 585
R827 B.n632 B.n631 585
R828 B.n631 B.n630 585
R829 B.n335 B.n334 585
R830 B.n336 B.n335 585
R831 B.n623 B.n622 585
R832 B.n624 B.n623 585
R833 B.n621 B.n341 585
R834 B.n341 B.n340 585
R835 B.n620 B.n619 585
R836 B.n619 B.n618 585
R837 B.n343 B.n342 585
R838 B.n344 B.n343 585
R839 B.n611 B.n610 585
R840 B.n612 B.n611 585
R841 B.n609 B.n349 585
R842 B.n349 B.n348 585
R843 B.n608 B.n607 585
R844 B.n607 B.n606 585
R845 B.n351 B.n350 585
R846 B.n352 B.n351 585
R847 B.n599 B.n598 585
R848 B.n600 B.n599 585
R849 B.n597 B.n357 585
R850 B.n357 B.n356 585
R851 B.n596 B.n595 585
R852 B.n595 B.n594 585
R853 B.n359 B.n358 585
R854 B.n360 B.n359 585
R855 B.n587 B.n586 585
R856 B.n588 B.n587 585
R857 B.n585 B.n364 585
R858 B.n368 B.n364 585
R859 B.n584 B.n583 585
R860 B.n583 B.n582 585
R861 B.n366 B.n365 585
R862 B.n367 B.n366 585
R863 B.n575 B.n574 585
R864 B.n576 B.n575 585
R865 B.n573 B.n373 585
R866 B.n373 B.n372 585
R867 B.n572 B.n571 585
R868 B.n571 B.n570 585
R869 B.n375 B.n374 585
R870 B.n376 B.n375 585
R871 B.n566 B.n565 585
R872 B.n379 B.n378 585
R873 B.n562 B.n561 585
R874 B.n563 B.n562 585
R875 B.n560 B.n415 585
R876 B.n559 B.n558 585
R877 B.n557 B.n556 585
R878 B.n555 B.n554 585
R879 B.n553 B.n552 585
R880 B.n551 B.n550 585
R881 B.n549 B.n548 585
R882 B.n547 B.n546 585
R883 B.n545 B.n544 585
R884 B.n543 B.n542 585
R885 B.n541 B.n540 585
R886 B.n539 B.n538 585
R887 B.n537 B.n536 585
R888 B.n535 B.n534 585
R889 B.n533 B.n532 585
R890 B.n531 B.n530 585
R891 B.n529 B.n528 585
R892 B.n527 B.n526 585
R893 B.n525 B.n524 585
R894 B.n523 B.n522 585
R895 B.n521 B.n520 585
R896 B.n519 B.n518 585
R897 B.n517 B.n516 585
R898 B.n515 B.n514 585
R899 B.n513 B.n512 585
R900 B.n511 B.n510 585
R901 B.n509 B.n508 585
R902 B.n507 B.n506 585
R903 B.n505 B.n504 585
R904 B.n502 B.n501 585
R905 B.n500 B.n499 585
R906 B.n498 B.n497 585
R907 B.n496 B.n495 585
R908 B.n494 B.n493 585
R909 B.n492 B.n491 585
R910 B.n490 B.n489 585
R911 B.n488 B.n487 585
R912 B.n486 B.n485 585
R913 B.n484 B.n483 585
R914 B.n482 B.n481 585
R915 B.n480 B.n479 585
R916 B.n478 B.n477 585
R917 B.n476 B.n475 585
R918 B.n474 B.n473 585
R919 B.n472 B.n471 585
R920 B.n470 B.n469 585
R921 B.n468 B.n467 585
R922 B.n466 B.n465 585
R923 B.n464 B.n463 585
R924 B.n462 B.n461 585
R925 B.n460 B.n459 585
R926 B.n458 B.n457 585
R927 B.n456 B.n455 585
R928 B.n454 B.n453 585
R929 B.n452 B.n451 585
R930 B.n450 B.n449 585
R931 B.n448 B.n447 585
R932 B.n446 B.n445 585
R933 B.n444 B.n443 585
R934 B.n442 B.n441 585
R935 B.n440 B.n439 585
R936 B.n438 B.n437 585
R937 B.n436 B.n435 585
R938 B.n434 B.n433 585
R939 B.n432 B.n431 585
R940 B.n430 B.n429 585
R941 B.n428 B.n427 585
R942 B.n426 B.n425 585
R943 B.n424 B.n423 585
R944 B.n422 B.n421 585
R945 B.n567 B.n377 585
R946 B.n377 B.n376 585
R947 B.n569 B.n568 585
R948 B.n570 B.n569 585
R949 B.n371 B.n370 585
R950 B.n372 B.n371 585
R951 B.n578 B.n577 585
R952 B.n577 B.n576 585
R953 B.n579 B.n369 585
R954 B.n369 B.n367 585
R955 B.n581 B.n580 585
R956 B.n582 B.n581 585
R957 B.n363 B.n362 585
R958 B.n368 B.n363 585
R959 B.n590 B.n589 585
R960 B.n589 B.n588 585
R961 B.n591 B.n361 585
R962 B.n361 B.n360 585
R963 B.n593 B.n592 585
R964 B.n594 B.n593 585
R965 B.n355 B.n354 585
R966 B.n356 B.n355 585
R967 B.n602 B.n601 585
R968 B.n601 B.n600 585
R969 B.n603 B.n353 585
R970 B.n353 B.n352 585
R971 B.n605 B.n604 585
R972 B.n606 B.n605 585
R973 B.n347 B.n346 585
R974 B.n348 B.n347 585
R975 B.n614 B.n613 585
R976 B.n613 B.n612 585
R977 B.n615 B.n345 585
R978 B.n345 B.n344 585
R979 B.n617 B.n616 585
R980 B.n618 B.n617 585
R981 B.n339 B.n338 585
R982 B.n340 B.n339 585
R983 B.n626 B.n625 585
R984 B.n625 B.n624 585
R985 B.n627 B.n337 585
R986 B.n337 B.n336 585
R987 B.n629 B.n628 585
R988 B.n630 B.n629 585
R989 B.n331 B.n330 585
R990 B.n332 B.n331 585
R991 B.n639 B.n638 585
R992 B.n638 B.n637 585
R993 B.n640 B.n329 585
R994 B.n636 B.n329 585
R995 B.n642 B.n641 585
R996 B.n643 B.n642 585
R997 B.n324 B.n323 585
R998 B.n325 B.n324 585
R999 B.n651 B.n650 585
R1000 B.n650 B.n649 585
R1001 B.n652 B.n322 585
R1002 B.n322 B.n321 585
R1003 B.n654 B.n653 585
R1004 B.n655 B.n654 585
R1005 B.n316 B.n315 585
R1006 B.n317 B.n316 585
R1007 B.n663 B.n662 585
R1008 B.n662 B.n661 585
R1009 B.n664 B.n314 585
R1010 B.n314 B.n313 585
R1011 B.n666 B.n665 585
R1012 B.n667 B.n666 585
R1013 B.n308 B.n307 585
R1014 B.n309 B.n308 585
R1015 B.n675 B.n674 585
R1016 B.n674 B.n673 585
R1017 B.n676 B.n306 585
R1018 B.n306 B.n305 585
R1019 B.n678 B.n677 585
R1020 B.n679 B.n678 585
R1021 B.n300 B.n299 585
R1022 B.n301 B.n300 585
R1023 B.n686 B.n685 585
R1024 B.n685 B.t3 585
R1025 B.n687 B.n298 585
R1026 B.n298 B.n297 585
R1027 B.n689 B.n688 585
R1028 B.n690 B.n689 585
R1029 B.n292 B.n291 585
R1030 B.n293 B.n292 585
R1031 B.n698 B.n697 585
R1032 B.n697 B.n696 585
R1033 B.n699 B.n290 585
R1034 B.n290 B.n288 585
R1035 B.n701 B.n700 585
R1036 B.n702 B.n701 585
R1037 B.n284 B.n283 585
R1038 B.n289 B.n284 585
R1039 B.n711 B.n710 585
R1040 B.n710 B.n709 585
R1041 B.n712 B.n282 585
R1042 B.n282 B.n281 585
R1043 B.n714 B.n713 585
R1044 B.n715 B.n714 585
R1045 B.n3 B.n0 585
R1046 B.n4 B.n3 585
R1047 B.n889 B.n1 585
R1048 B.n890 B.n889 585
R1049 B.n888 B.n887 585
R1050 B.n888 B.n8 585
R1051 B.n886 B.n9 585
R1052 B.n12 B.n9 585
R1053 B.n885 B.n884 585
R1054 B.n884 B.n883 585
R1055 B.n11 B.n10 585
R1056 B.n882 B.n11 585
R1057 B.n880 B.n879 585
R1058 B.n881 B.n880 585
R1059 B.n878 B.n17 585
R1060 B.n17 B.n16 585
R1061 B.n877 B.n876 585
R1062 B.n876 B.n875 585
R1063 B.n19 B.n18 585
R1064 B.n874 B.n19 585
R1065 B.n872 B.n871 585
R1066 B.n873 B.n872 585
R1067 B.n870 B.n24 585
R1068 B.n24 B.n23 585
R1069 B.n869 B.n868 585
R1070 B.n868 B.t0 585
R1071 B.n26 B.n25 585
R1072 B.n867 B.n26 585
R1073 B.n865 B.n864 585
R1074 B.n866 B.n865 585
R1075 B.n863 B.n31 585
R1076 B.n31 B.n30 585
R1077 B.n862 B.n861 585
R1078 B.n861 B.n860 585
R1079 B.n33 B.n32 585
R1080 B.n859 B.n33 585
R1081 B.n857 B.n856 585
R1082 B.n858 B.n857 585
R1083 B.n855 B.n38 585
R1084 B.n38 B.n37 585
R1085 B.n854 B.n853 585
R1086 B.n853 B.n852 585
R1087 B.n40 B.n39 585
R1088 B.n851 B.n40 585
R1089 B.n849 B.n848 585
R1090 B.n850 B.n849 585
R1091 B.n847 B.n45 585
R1092 B.n45 B.n44 585
R1093 B.n846 B.n845 585
R1094 B.n845 B.n844 585
R1095 B.n47 B.n46 585
R1096 B.n843 B.n47 585
R1097 B.n841 B.n840 585
R1098 B.n842 B.n841 585
R1099 B.n839 B.n51 585
R1100 B.n54 B.n51 585
R1101 B.n838 B.n837 585
R1102 B.n837 B.n836 585
R1103 B.n53 B.n52 585
R1104 B.n835 B.n53 585
R1105 B.n833 B.n832 585
R1106 B.n834 B.n833 585
R1107 B.n831 B.n59 585
R1108 B.n59 B.n58 585
R1109 B.n830 B.n829 585
R1110 B.n829 B.n828 585
R1111 B.n61 B.n60 585
R1112 B.n827 B.n61 585
R1113 B.n825 B.n824 585
R1114 B.n826 B.n825 585
R1115 B.n823 B.n66 585
R1116 B.n66 B.n65 585
R1117 B.n822 B.n821 585
R1118 B.n821 B.n820 585
R1119 B.n68 B.n67 585
R1120 B.n819 B.n68 585
R1121 B.n817 B.n816 585
R1122 B.n818 B.n817 585
R1123 B.n815 B.n73 585
R1124 B.n73 B.n72 585
R1125 B.n814 B.n813 585
R1126 B.n813 B.n812 585
R1127 B.n75 B.n74 585
R1128 B.n811 B.n75 585
R1129 B.n809 B.n808 585
R1130 B.n810 B.n809 585
R1131 B.n807 B.n80 585
R1132 B.n80 B.n79 585
R1133 B.n806 B.n805 585
R1134 B.n805 B.n804 585
R1135 B.n82 B.n81 585
R1136 B.n803 B.n82 585
R1137 B.n801 B.n800 585
R1138 B.n802 B.n801 585
R1139 B.n799 B.n87 585
R1140 B.n87 B.n86 585
R1141 B.n798 B.n797 585
R1142 B.n797 B.n796 585
R1143 B.n89 B.n88 585
R1144 B.n795 B.n89 585
R1145 B.n793 B.n792 585
R1146 B.n794 B.n793 585
R1147 B.n791 B.n94 585
R1148 B.n94 B.n93 585
R1149 B.n893 B.n892 585
R1150 B.n891 B.n2 585
R1151 B.n789 B.n94 502.111
R1152 B.n786 B.n133 502.111
R1153 B.n421 B.n375 502.111
R1154 B.n565 B.n377 502.111
R1155 B.n136 B.t10 303.741
R1156 B.n134 B.t14 303.741
R1157 B.n418 B.t21 303.741
R1158 B.n416 B.t17 303.741
R1159 B.n134 B.t15 270.769
R1160 B.n418 B.t23 270.769
R1161 B.n136 B.t12 270.769
R1162 B.n416 B.t20 270.769
R1163 B.n787 B.n131 256.663
R1164 B.n787 B.n130 256.663
R1165 B.n787 B.n129 256.663
R1166 B.n787 B.n128 256.663
R1167 B.n787 B.n127 256.663
R1168 B.n787 B.n126 256.663
R1169 B.n787 B.n125 256.663
R1170 B.n787 B.n124 256.663
R1171 B.n787 B.n123 256.663
R1172 B.n787 B.n122 256.663
R1173 B.n787 B.n121 256.663
R1174 B.n787 B.n120 256.663
R1175 B.n787 B.n119 256.663
R1176 B.n787 B.n118 256.663
R1177 B.n787 B.n117 256.663
R1178 B.n787 B.n116 256.663
R1179 B.n787 B.n115 256.663
R1180 B.n787 B.n114 256.663
R1181 B.n787 B.n113 256.663
R1182 B.n787 B.n112 256.663
R1183 B.n787 B.n111 256.663
R1184 B.n787 B.n110 256.663
R1185 B.n787 B.n109 256.663
R1186 B.n787 B.n108 256.663
R1187 B.n787 B.n107 256.663
R1188 B.n787 B.n106 256.663
R1189 B.n787 B.n105 256.663
R1190 B.n787 B.n104 256.663
R1191 B.n787 B.n103 256.663
R1192 B.n787 B.n102 256.663
R1193 B.n787 B.n101 256.663
R1194 B.n787 B.n100 256.663
R1195 B.n787 B.n99 256.663
R1196 B.n787 B.n98 256.663
R1197 B.n787 B.n97 256.663
R1198 B.n788 B.n787 256.663
R1199 B.n564 B.n563 256.663
R1200 B.n563 B.n380 256.663
R1201 B.n563 B.n381 256.663
R1202 B.n563 B.n382 256.663
R1203 B.n563 B.n383 256.663
R1204 B.n563 B.n384 256.663
R1205 B.n563 B.n385 256.663
R1206 B.n563 B.n386 256.663
R1207 B.n563 B.n387 256.663
R1208 B.n563 B.n388 256.663
R1209 B.n563 B.n389 256.663
R1210 B.n563 B.n390 256.663
R1211 B.n563 B.n391 256.663
R1212 B.n563 B.n392 256.663
R1213 B.n563 B.n393 256.663
R1214 B.n563 B.n394 256.663
R1215 B.n563 B.n395 256.663
R1216 B.n563 B.n396 256.663
R1217 B.n563 B.n397 256.663
R1218 B.n563 B.n398 256.663
R1219 B.n563 B.n399 256.663
R1220 B.n563 B.n400 256.663
R1221 B.n563 B.n401 256.663
R1222 B.n563 B.n402 256.663
R1223 B.n563 B.n403 256.663
R1224 B.n563 B.n404 256.663
R1225 B.n563 B.n405 256.663
R1226 B.n563 B.n406 256.663
R1227 B.n563 B.n407 256.663
R1228 B.n563 B.n408 256.663
R1229 B.n563 B.n409 256.663
R1230 B.n563 B.n410 256.663
R1231 B.n563 B.n411 256.663
R1232 B.n563 B.n412 256.663
R1233 B.n563 B.n413 256.663
R1234 B.n563 B.n414 256.663
R1235 B.n895 B.n894 256.663
R1236 B.n135 B.t16 222.867
R1237 B.n419 B.t22 222.867
R1238 B.n137 B.t13 222.867
R1239 B.n417 B.t19 222.867
R1240 B.n139 B.n96 163.367
R1241 B.n143 B.n142 163.367
R1242 B.n147 B.n146 163.367
R1243 B.n151 B.n150 163.367
R1244 B.n155 B.n154 163.367
R1245 B.n159 B.n158 163.367
R1246 B.n163 B.n162 163.367
R1247 B.n167 B.n166 163.367
R1248 B.n171 B.n170 163.367
R1249 B.n175 B.n174 163.367
R1250 B.n179 B.n178 163.367
R1251 B.n183 B.n182 163.367
R1252 B.n187 B.n186 163.367
R1253 B.n191 B.n190 163.367
R1254 B.n195 B.n194 163.367
R1255 B.n199 B.n198 163.367
R1256 B.n203 B.n202 163.367
R1257 B.n207 B.n206 163.367
R1258 B.n211 B.n210 163.367
R1259 B.n215 B.n214 163.367
R1260 B.n220 B.n219 163.367
R1261 B.n224 B.n223 163.367
R1262 B.n228 B.n227 163.367
R1263 B.n232 B.n231 163.367
R1264 B.n236 B.n235 163.367
R1265 B.n240 B.n239 163.367
R1266 B.n244 B.n243 163.367
R1267 B.n248 B.n247 163.367
R1268 B.n252 B.n251 163.367
R1269 B.n256 B.n255 163.367
R1270 B.n260 B.n259 163.367
R1271 B.n264 B.n263 163.367
R1272 B.n268 B.n267 163.367
R1273 B.n272 B.n271 163.367
R1274 B.n276 B.n275 163.367
R1275 B.n786 B.n132 163.367
R1276 B.n571 B.n375 163.367
R1277 B.n571 B.n373 163.367
R1278 B.n575 B.n373 163.367
R1279 B.n575 B.n366 163.367
R1280 B.n583 B.n366 163.367
R1281 B.n583 B.n364 163.367
R1282 B.n587 B.n364 163.367
R1283 B.n587 B.n359 163.367
R1284 B.n595 B.n359 163.367
R1285 B.n595 B.n357 163.367
R1286 B.n599 B.n357 163.367
R1287 B.n599 B.n351 163.367
R1288 B.n607 B.n351 163.367
R1289 B.n607 B.n349 163.367
R1290 B.n611 B.n349 163.367
R1291 B.n611 B.n343 163.367
R1292 B.n619 B.n343 163.367
R1293 B.n619 B.n341 163.367
R1294 B.n623 B.n341 163.367
R1295 B.n623 B.n335 163.367
R1296 B.n631 B.n335 163.367
R1297 B.n631 B.n333 163.367
R1298 B.n635 B.n333 163.367
R1299 B.n635 B.n328 163.367
R1300 B.n644 B.n328 163.367
R1301 B.n644 B.n326 163.367
R1302 B.n648 B.n326 163.367
R1303 B.n648 B.n320 163.367
R1304 B.n656 B.n320 163.367
R1305 B.n656 B.n318 163.367
R1306 B.n660 B.n318 163.367
R1307 B.n660 B.n312 163.367
R1308 B.n668 B.n312 163.367
R1309 B.n668 B.n310 163.367
R1310 B.n672 B.n310 163.367
R1311 B.n672 B.n304 163.367
R1312 B.n680 B.n304 163.367
R1313 B.n680 B.n302 163.367
R1314 B.n684 B.n302 163.367
R1315 B.n684 B.n296 163.367
R1316 B.n691 B.n296 163.367
R1317 B.n691 B.n294 163.367
R1318 B.n695 B.n294 163.367
R1319 B.n695 B.n287 163.367
R1320 B.n703 B.n287 163.367
R1321 B.n703 B.n285 163.367
R1322 B.n708 B.n285 163.367
R1323 B.n708 B.n280 163.367
R1324 B.n716 B.n280 163.367
R1325 B.n717 B.n716 163.367
R1326 B.n717 B.n5 163.367
R1327 B.n6 B.n5 163.367
R1328 B.n7 B.n6 163.367
R1329 B.n723 B.n7 163.367
R1330 B.n724 B.n723 163.367
R1331 B.n724 B.n13 163.367
R1332 B.n14 B.n13 163.367
R1333 B.n15 B.n14 163.367
R1334 B.n729 B.n15 163.367
R1335 B.n729 B.n20 163.367
R1336 B.n21 B.n20 163.367
R1337 B.n22 B.n21 163.367
R1338 B.n734 B.n22 163.367
R1339 B.n734 B.n27 163.367
R1340 B.n28 B.n27 163.367
R1341 B.n29 B.n28 163.367
R1342 B.n739 B.n29 163.367
R1343 B.n739 B.n34 163.367
R1344 B.n35 B.n34 163.367
R1345 B.n36 B.n35 163.367
R1346 B.n744 B.n36 163.367
R1347 B.n744 B.n41 163.367
R1348 B.n42 B.n41 163.367
R1349 B.n43 B.n42 163.367
R1350 B.n749 B.n43 163.367
R1351 B.n749 B.n48 163.367
R1352 B.n49 B.n48 163.367
R1353 B.n50 B.n49 163.367
R1354 B.n754 B.n50 163.367
R1355 B.n754 B.n55 163.367
R1356 B.n56 B.n55 163.367
R1357 B.n57 B.n56 163.367
R1358 B.n759 B.n57 163.367
R1359 B.n759 B.n62 163.367
R1360 B.n63 B.n62 163.367
R1361 B.n64 B.n63 163.367
R1362 B.n764 B.n64 163.367
R1363 B.n764 B.n69 163.367
R1364 B.n70 B.n69 163.367
R1365 B.n71 B.n70 163.367
R1366 B.n769 B.n71 163.367
R1367 B.n769 B.n76 163.367
R1368 B.n77 B.n76 163.367
R1369 B.n78 B.n77 163.367
R1370 B.n774 B.n78 163.367
R1371 B.n774 B.n83 163.367
R1372 B.n84 B.n83 163.367
R1373 B.n85 B.n84 163.367
R1374 B.n779 B.n85 163.367
R1375 B.n779 B.n90 163.367
R1376 B.n91 B.n90 163.367
R1377 B.n92 B.n91 163.367
R1378 B.n133 B.n92 163.367
R1379 B.n562 B.n379 163.367
R1380 B.n562 B.n415 163.367
R1381 B.n558 B.n557 163.367
R1382 B.n554 B.n553 163.367
R1383 B.n550 B.n549 163.367
R1384 B.n546 B.n545 163.367
R1385 B.n542 B.n541 163.367
R1386 B.n538 B.n537 163.367
R1387 B.n534 B.n533 163.367
R1388 B.n530 B.n529 163.367
R1389 B.n526 B.n525 163.367
R1390 B.n522 B.n521 163.367
R1391 B.n518 B.n517 163.367
R1392 B.n514 B.n513 163.367
R1393 B.n510 B.n509 163.367
R1394 B.n506 B.n505 163.367
R1395 B.n501 B.n500 163.367
R1396 B.n497 B.n496 163.367
R1397 B.n493 B.n492 163.367
R1398 B.n489 B.n488 163.367
R1399 B.n485 B.n484 163.367
R1400 B.n481 B.n480 163.367
R1401 B.n477 B.n476 163.367
R1402 B.n473 B.n472 163.367
R1403 B.n469 B.n468 163.367
R1404 B.n465 B.n464 163.367
R1405 B.n461 B.n460 163.367
R1406 B.n457 B.n456 163.367
R1407 B.n453 B.n452 163.367
R1408 B.n449 B.n448 163.367
R1409 B.n445 B.n444 163.367
R1410 B.n441 B.n440 163.367
R1411 B.n437 B.n436 163.367
R1412 B.n433 B.n432 163.367
R1413 B.n429 B.n428 163.367
R1414 B.n425 B.n424 163.367
R1415 B.n569 B.n377 163.367
R1416 B.n569 B.n371 163.367
R1417 B.n577 B.n371 163.367
R1418 B.n577 B.n369 163.367
R1419 B.n581 B.n369 163.367
R1420 B.n581 B.n363 163.367
R1421 B.n589 B.n363 163.367
R1422 B.n589 B.n361 163.367
R1423 B.n593 B.n361 163.367
R1424 B.n593 B.n355 163.367
R1425 B.n601 B.n355 163.367
R1426 B.n601 B.n353 163.367
R1427 B.n605 B.n353 163.367
R1428 B.n605 B.n347 163.367
R1429 B.n613 B.n347 163.367
R1430 B.n613 B.n345 163.367
R1431 B.n617 B.n345 163.367
R1432 B.n617 B.n339 163.367
R1433 B.n625 B.n339 163.367
R1434 B.n625 B.n337 163.367
R1435 B.n629 B.n337 163.367
R1436 B.n629 B.n331 163.367
R1437 B.n638 B.n331 163.367
R1438 B.n638 B.n329 163.367
R1439 B.n642 B.n329 163.367
R1440 B.n642 B.n324 163.367
R1441 B.n650 B.n324 163.367
R1442 B.n650 B.n322 163.367
R1443 B.n654 B.n322 163.367
R1444 B.n654 B.n316 163.367
R1445 B.n662 B.n316 163.367
R1446 B.n662 B.n314 163.367
R1447 B.n666 B.n314 163.367
R1448 B.n666 B.n308 163.367
R1449 B.n674 B.n308 163.367
R1450 B.n674 B.n306 163.367
R1451 B.n678 B.n306 163.367
R1452 B.n678 B.n300 163.367
R1453 B.n685 B.n300 163.367
R1454 B.n685 B.n298 163.367
R1455 B.n689 B.n298 163.367
R1456 B.n689 B.n292 163.367
R1457 B.n697 B.n292 163.367
R1458 B.n697 B.n290 163.367
R1459 B.n701 B.n290 163.367
R1460 B.n701 B.n284 163.367
R1461 B.n710 B.n284 163.367
R1462 B.n710 B.n282 163.367
R1463 B.n714 B.n282 163.367
R1464 B.n714 B.n3 163.367
R1465 B.n893 B.n3 163.367
R1466 B.n889 B.n2 163.367
R1467 B.n889 B.n888 163.367
R1468 B.n888 B.n9 163.367
R1469 B.n884 B.n9 163.367
R1470 B.n884 B.n11 163.367
R1471 B.n880 B.n11 163.367
R1472 B.n880 B.n17 163.367
R1473 B.n876 B.n17 163.367
R1474 B.n876 B.n19 163.367
R1475 B.n872 B.n19 163.367
R1476 B.n872 B.n24 163.367
R1477 B.n868 B.n24 163.367
R1478 B.n868 B.n26 163.367
R1479 B.n865 B.n26 163.367
R1480 B.n865 B.n31 163.367
R1481 B.n861 B.n31 163.367
R1482 B.n861 B.n33 163.367
R1483 B.n857 B.n33 163.367
R1484 B.n857 B.n38 163.367
R1485 B.n853 B.n38 163.367
R1486 B.n853 B.n40 163.367
R1487 B.n849 B.n40 163.367
R1488 B.n849 B.n45 163.367
R1489 B.n845 B.n45 163.367
R1490 B.n845 B.n47 163.367
R1491 B.n841 B.n47 163.367
R1492 B.n841 B.n51 163.367
R1493 B.n837 B.n51 163.367
R1494 B.n837 B.n53 163.367
R1495 B.n833 B.n53 163.367
R1496 B.n833 B.n59 163.367
R1497 B.n829 B.n59 163.367
R1498 B.n829 B.n61 163.367
R1499 B.n825 B.n61 163.367
R1500 B.n825 B.n66 163.367
R1501 B.n821 B.n66 163.367
R1502 B.n821 B.n68 163.367
R1503 B.n817 B.n68 163.367
R1504 B.n817 B.n73 163.367
R1505 B.n813 B.n73 163.367
R1506 B.n813 B.n75 163.367
R1507 B.n809 B.n75 163.367
R1508 B.n809 B.n80 163.367
R1509 B.n805 B.n80 163.367
R1510 B.n805 B.n82 163.367
R1511 B.n801 B.n82 163.367
R1512 B.n801 B.n87 163.367
R1513 B.n797 B.n87 163.367
R1514 B.n797 B.n89 163.367
R1515 B.n793 B.n89 163.367
R1516 B.n793 B.n94 163.367
R1517 B.n563 B.n376 108.849
R1518 B.n787 B.n93 108.849
R1519 B.n789 B.n788 71.676
R1520 B.n139 B.n97 71.676
R1521 B.n143 B.n98 71.676
R1522 B.n147 B.n99 71.676
R1523 B.n151 B.n100 71.676
R1524 B.n155 B.n101 71.676
R1525 B.n159 B.n102 71.676
R1526 B.n163 B.n103 71.676
R1527 B.n167 B.n104 71.676
R1528 B.n171 B.n105 71.676
R1529 B.n175 B.n106 71.676
R1530 B.n179 B.n107 71.676
R1531 B.n183 B.n108 71.676
R1532 B.n187 B.n109 71.676
R1533 B.n191 B.n110 71.676
R1534 B.n195 B.n111 71.676
R1535 B.n199 B.n112 71.676
R1536 B.n203 B.n113 71.676
R1537 B.n207 B.n114 71.676
R1538 B.n211 B.n115 71.676
R1539 B.n215 B.n116 71.676
R1540 B.n220 B.n117 71.676
R1541 B.n224 B.n118 71.676
R1542 B.n228 B.n119 71.676
R1543 B.n232 B.n120 71.676
R1544 B.n236 B.n121 71.676
R1545 B.n240 B.n122 71.676
R1546 B.n244 B.n123 71.676
R1547 B.n248 B.n124 71.676
R1548 B.n252 B.n125 71.676
R1549 B.n256 B.n126 71.676
R1550 B.n260 B.n127 71.676
R1551 B.n264 B.n128 71.676
R1552 B.n268 B.n129 71.676
R1553 B.n272 B.n130 71.676
R1554 B.n276 B.n131 71.676
R1555 B.n132 B.n131 71.676
R1556 B.n275 B.n130 71.676
R1557 B.n271 B.n129 71.676
R1558 B.n267 B.n128 71.676
R1559 B.n263 B.n127 71.676
R1560 B.n259 B.n126 71.676
R1561 B.n255 B.n125 71.676
R1562 B.n251 B.n124 71.676
R1563 B.n247 B.n123 71.676
R1564 B.n243 B.n122 71.676
R1565 B.n239 B.n121 71.676
R1566 B.n235 B.n120 71.676
R1567 B.n231 B.n119 71.676
R1568 B.n227 B.n118 71.676
R1569 B.n223 B.n117 71.676
R1570 B.n219 B.n116 71.676
R1571 B.n214 B.n115 71.676
R1572 B.n210 B.n114 71.676
R1573 B.n206 B.n113 71.676
R1574 B.n202 B.n112 71.676
R1575 B.n198 B.n111 71.676
R1576 B.n194 B.n110 71.676
R1577 B.n190 B.n109 71.676
R1578 B.n186 B.n108 71.676
R1579 B.n182 B.n107 71.676
R1580 B.n178 B.n106 71.676
R1581 B.n174 B.n105 71.676
R1582 B.n170 B.n104 71.676
R1583 B.n166 B.n103 71.676
R1584 B.n162 B.n102 71.676
R1585 B.n158 B.n101 71.676
R1586 B.n154 B.n100 71.676
R1587 B.n150 B.n99 71.676
R1588 B.n146 B.n98 71.676
R1589 B.n142 B.n97 71.676
R1590 B.n788 B.n96 71.676
R1591 B.n565 B.n564 71.676
R1592 B.n415 B.n380 71.676
R1593 B.n557 B.n381 71.676
R1594 B.n553 B.n382 71.676
R1595 B.n549 B.n383 71.676
R1596 B.n545 B.n384 71.676
R1597 B.n541 B.n385 71.676
R1598 B.n537 B.n386 71.676
R1599 B.n533 B.n387 71.676
R1600 B.n529 B.n388 71.676
R1601 B.n525 B.n389 71.676
R1602 B.n521 B.n390 71.676
R1603 B.n517 B.n391 71.676
R1604 B.n513 B.n392 71.676
R1605 B.n509 B.n393 71.676
R1606 B.n505 B.n394 71.676
R1607 B.n500 B.n395 71.676
R1608 B.n496 B.n396 71.676
R1609 B.n492 B.n397 71.676
R1610 B.n488 B.n398 71.676
R1611 B.n484 B.n399 71.676
R1612 B.n480 B.n400 71.676
R1613 B.n476 B.n401 71.676
R1614 B.n472 B.n402 71.676
R1615 B.n468 B.n403 71.676
R1616 B.n464 B.n404 71.676
R1617 B.n460 B.n405 71.676
R1618 B.n456 B.n406 71.676
R1619 B.n452 B.n407 71.676
R1620 B.n448 B.n408 71.676
R1621 B.n444 B.n409 71.676
R1622 B.n440 B.n410 71.676
R1623 B.n436 B.n411 71.676
R1624 B.n432 B.n412 71.676
R1625 B.n428 B.n413 71.676
R1626 B.n424 B.n414 71.676
R1627 B.n564 B.n379 71.676
R1628 B.n558 B.n380 71.676
R1629 B.n554 B.n381 71.676
R1630 B.n550 B.n382 71.676
R1631 B.n546 B.n383 71.676
R1632 B.n542 B.n384 71.676
R1633 B.n538 B.n385 71.676
R1634 B.n534 B.n386 71.676
R1635 B.n530 B.n387 71.676
R1636 B.n526 B.n388 71.676
R1637 B.n522 B.n389 71.676
R1638 B.n518 B.n390 71.676
R1639 B.n514 B.n391 71.676
R1640 B.n510 B.n392 71.676
R1641 B.n506 B.n393 71.676
R1642 B.n501 B.n394 71.676
R1643 B.n497 B.n395 71.676
R1644 B.n493 B.n396 71.676
R1645 B.n489 B.n397 71.676
R1646 B.n485 B.n398 71.676
R1647 B.n481 B.n399 71.676
R1648 B.n477 B.n400 71.676
R1649 B.n473 B.n401 71.676
R1650 B.n469 B.n402 71.676
R1651 B.n465 B.n403 71.676
R1652 B.n461 B.n404 71.676
R1653 B.n457 B.n405 71.676
R1654 B.n453 B.n406 71.676
R1655 B.n449 B.n407 71.676
R1656 B.n445 B.n408 71.676
R1657 B.n441 B.n409 71.676
R1658 B.n437 B.n410 71.676
R1659 B.n433 B.n411 71.676
R1660 B.n429 B.n412 71.676
R1661 B.n425 B.n413 71.676
R1662 B.n421 B.n414 71.676
R1663 B.n894 B.n893 71.676
R1664 B.n894 B.n2 71.676
R1665 B.n138 B.n137 59.5399
R1666 B.n217 B.n135 59.5399
R1667 B.n420 B.n419 59.5399
R1668 B.n503 B.n417 59.5399
R1669 B.n570 B.n376 54.0272
R1670 B.n570 B.n372 54.0272
R1671 B.n576 B.n372 54.0272
R1672 B.n576 B.n367 54.0272
R1673 B.n582 B.n367 54.0272
R1674 B.n582 B.n368 54.0272
R1675 B.n588 B.n360 54.0272
R1676 B.n594 B.n360 54.0272
R1677 B.n594 B.n356 54.0272
R1678 B.n600 B.n356 54.0272
R1679 B.n600 B.n352 54.0272
R1680 B.n606 B.n352 54.0272
R1681 B.n606 B.n348 54.0272
R1682 B.n612 B.n348 54.0272
R1683 B.n612 B.n344 54.0272
R1684 B.n618 B.n344 54.0272
R1685 B.n624 B.n340 54.0272
R1686 B.n624 B.n336 54.0272
R1687 B.n630 B.n336 54.0272
R1688 B.n630 B.n332 54.0272
R1689 B.n637 B.n332 54.0272
R1690 B.n637 B.n636 54.0272
R1691 B.n643 B.n325 54.0272
R1692 B.n649 B.n325 54.0272
R1693 B.n649 B.n321 54.0272
R1694 B.n655 B.n321 54.0272
R1695 B.n655 B.n317 54.0272
R1696 B.n661 B.n317 54.0272
R1697 B.n667 B.n313 54.0272
R1698 B.n667 B.n309 54.0272
R1699 B.n673 B.n309 54.0272
R1700 B.n673 B.n305 54.0272
R1701 B.n679 B.n305 54.0272
R1702 B.n679 B.n301 54.0272
R1703 B.t3 B.n301 54.0272
R1704 B.t3 B.n297 54.0272
R1705 B.n690 B.n297 54.0272
R1706 B.n690 B.n293 54.0272
R1707 B.n696 B.n293 54.0272
R1708 B.n696 B.n288 54.0272
R1709 B.n702 B.n288 54.0272
R1710 B.n702 B.n289 54.0272
R1711 B.n709 B.n281 54.0272
R1712 B.n715 B.n281 54.0272
R1713 B.n715 B.n4 54.0272
R1714 B.n892 B.n4 54.0272
R1715 B.n892 B.n891 54.0272
R1716 B.n891 B.n890 54.0272
R1717 B.n890 B.n8 54.0272
R1718 B.n12 B.n8 54.0272
R1719 B.n883 B.n12 54.0272
R1720 B.n882 B.n881 54.0272
R1721 B.n881 B.n16 54.0272
R1722 B.n875 B.n16 54.0272
R1723 B.n875 B.n874 54.0272
R1724 B.n874 B.n873 54.0272
R1725 B.n873 B.n23 54.0272
R1726 B.t0 B.n23 54.0272
R1727 B.t0 B.n867 54.0272
R1728 B.n867 B.n866 54.0272
R1729 B.n866 B.n30 54.0272
R1730 B.n860 B.n30 54.0272
R1731 B.n860 B.n859 54.0272
R1732 B.n859 B.n858 54.0272
R1733 B.n858 B.n37 54.0272
R1734 B.n852 B.n851 54.0272
R1735 B.n851 B.n850 54.0272
R1736 B.n850 B.n44 54.0272
R1737 B.n844 B.n44 54.0272
R1738 B.n844 B.n843 54.0272
R1739 B.n843 B.n842 54.0272
R1740 B.n836 B.n54 54.0272
R1741 B.n836 B.n835 54.0272
R1742 B.n835 B.n834 54.0272
R1743 B.n834 B.n58 54.0272
R1744 B.n828 B.n58 54.0272
R1745 B.n828 B.n827 54.0272
R1746 B.n826 B.n65 54.0272
R1747 B.n820 B.n65 54.0272
R1748 B.n820 B.n819 54.0272
R1749 B.n819 B.n818 54.0272
R1750 B.n818 B.n72 54.0272
R1751 B.n812 B.n72 54.0272
R1752 B.n812 B.n811 54.0272
R1753 B.n811 B.n810 54.0272
R1754 B.n810 B.n79 54.0272
R1755 B.n804 B.n79 54.0272
R1756 B.n803 B.n802 54.0272
R1757 B.n802 B.n86 54.0272
R1758 B.n796 B.n86 54.0272
R1759 B.n796 B.n795 54.0272
R1760 B.n795 B.n794 54.0272
R1761 B.n794 B.n93 54.0272
R1762 B.n137 B.n136 47.9035
R1763 B.n135 B.n134 47.9035
R1764 B.n419 B.n418 47.9035
R1765 B.n417 B.n416 47.9035
R1766 B.t1 B.n340 42.9041
R1767 B.n827 B.t7 42.9041
R1768 B.n368 B.t18 39.726
R1769 B.n661 B.t4 39.726
R1770 B.n709 B.t9 39.726
R1771 B.n883 B.t2 39.726
R1772 B.n852 B.t5 39.726
R1773 B.t11 B.n803 39.726
R1774 B.n567 B.n566 32.6249
R1775 B.n422 B.n374 32.6249
R1776 B.n785 B.n784 32.6249
R1777 B.n791 B.n790 32.6249
R1778 B.n643 B.t6 28.6029
R1779 B.n842 B.t8 28.6029
R1780 B.n636 B.t6 25.4248
R1781 B.n54 B.t8 25.4248
R1782 B B.n895 18.0485
R1783 B.n588 B.t18 14.3017
R1784 B.t4 B.n313 14.3017
R1785 B.n289 B.t9 14.3017
R1786 B.t2 B.n882 14.3017
R1787 B.t5 B.n37 14.3017
R1788 B.n804 B.t11 14.3017
R1789 B.n618 B.t1 11.1236
R1790 B.t7 B.n826 11.1236
R1791 B.n568 B.n567 10.6151
R1792 B.n568 B.n370 10.6151
R1793 B.n578 B.n370 10.6151
R1794 B.n579 B.n578 10.6151
R1795 B.n580 B.n579 10.6151
R1796 B.n580 B.n362 10.6151
R1797 B.n590 B.n362 10.6151
R1798 B.n591 B.n590 10.6151
R1799 B.n592 B.n591 10.6151
R1800 B.n592 B.n354 10.6151
R1801 B.n602 B.n354 10.6151
R1802 B.n603 B.n602 10.6151
R1803 B.n604 B.n603 10.6151
R1804 B.n604 B.n346 10.6151
R1805 B.n614 B.n346 10.6151
R1806 B.n615 B.n614 10.6151
R1807 B.n616 B.n615 10.6151
R1808 B.n616 B.n338 10.6151
R1809 B.n626 B.n338 10.6151
R1810 B.n627 B.n626 10.6151
R1811 B.n628 B.n627 10.6151
R1812 B.n628 B.n330 10.6151
R1813 B.n639 B.n330 10.6151
R1814 B.n640 B.n639 10.6151
R1815 B.n641 B.n640 10.6151
R1816 B.n641 B.n323 10.6151
R1817 B.n651 B.n323 10.6151
R1818 B.n652 B.n651 10.6151
R1819 B.n653 B.n652 10.6151
R1820 B.n653 B.n315 10.6151
R1821 B.n663 B.n315 10.6151
R1822 B.n664 B.n663 10.6151
R1823 B.n665 B.n664 10.6151
R1824 B.n665 B.n307 10.6151
R1825 B.n675 B.n307 10.6151
R1826 B.n676 B.n675 10.6151
R1827 B.n677 B.n676 10.6151
R1828 B.n677 B.n299 10.6151
R1829 B.n686 B.n299 10.6151
R1830 B.n687 B.n686 10.6151
R1831 B.n688 B.n687 10.6151
R1832 B.n688 B.n291 10.6151
R1833 B.n698 B.n291 10.6151
R1834 B.n699 B.n698 10.6151
R1835 B.n700 B.n699 10.6151
R1836 B.n700 B.n283 10.6151
R1837 B.n711 B.n283 10.6151
R1838 B.n712 B.n711 10.6151
R1839 B.n713 B.n712 10.6151
R1840 B.n713 B.n0 10.6151
R1841 B.n566 B.n378 10.6151
R1842 B.n561 B.n378 10.6151
R1843 B.n561 B.n560 10.6151
R1844 B.n560 B.n559 10.6151
R1845 B.n559 B.n556 10.6151
R1846 B.n556 B.n555 10.6151
R1847 B.n555 B.n552 10.6151
R1848 B.n552 B.n551 10.6151
R1849 B.n551 B.n548 10.6151
R1850 B.n548 B.n547 10.6151
R1851 B.n547 B.n544 10.6151
R1852 B.n544 B.n543 10.6151
R1853 B.n543 B.n540 10.6151
R1854 B.n540 B.n539 10.6151
R1855 B.n539 B.n536 10.6151
R1856 B.n536 B.n535 10.6151
R1857 B.n535 B.n532 10.6151
R1858 B.n532 B.n531 10.6151
R1859 B.n531 B.n528 10.6151
R1860 B.n528 B.n527 10.6151
R1861 B.n527 B.n524 10.6151
R1862 B.n524 B.n523 10.6151
R1863 B.n523 B.n520 10.6151
R1864 B.n520 B.n519 10.6151
R1865 B.n519 B.n516 10.6151
R1866 B.n516 B.n515 10.6151
R1867 B.n515 B.n512 10.6151
R1868 B.n512 B.n511 10.6151
R1869 B.n511 B.n508 10.6151
R1870 B.n508 B.n507 10.6151
R1871 B.n507 B.n504 10.6151
R1872 B.n502 B.n499 10.6151
R1873 B.n499 B.n498 10.6151
R1874 B.n498 B.n495 10.6151
R1875 B.n495 B.n494 10.6151
R1876 B.n494 B.n491 10.6151
R1877 B.n491 B.n490 10.6151
R1878 B.n490 B.n487 10.6151
R1879 B.n487 B.n486 10.6151
R1880 B.n483 B.n482 10.6151
R1881 B.n482 B.n479 10.6151
R1882 B.n479 B.n478 10.6151
R1883 B.n478 B.n475 10.6151
R1884 B.n475 B.n474 10.6151
R1885 B.n474 B.n471 10.6151
R1886 B.n471 B.n470 10.6151
R1887 B.n470 B.n467 10.6151
R1888 B.n467 B.n466 10.6151
R1889 B.n466 B.n463 10.6151
R1890 B.n463 B.n462 10.6151
R1891 B.n462 B.n459 10.6151
R1892 B.n459 B.n458 10.6151
R1893 B.n458 B.n455 10.6151
R1894 B.n455 B.n454 10.6151
R1895 B.n454 B.n451 10.6151
R1896 B.n451 B.n450 10.6151
R1897 B.n450 B.n447 10.6151
R1898 B.n447 B.n446 10.6151
R1899 B.n446 B.n443 10.6151
R1900 B.n443 B.n442 10.6151
R1901 B.n442 B.n439 10.6151
R1902 B.n439 B.n438 10.6151
R1903 B.n438 B.n435 10.6151
R1904 B.n435 B.n434 10.6151
R1905 B.n434 B.n431 10.6151
R1906 B.n431 B.n430 10.6151
R1907 B.n430 B.n427 10.6151
R1908 B.n427 B.n426 10.6151
R1909 B.n426 B.n423 10.6151
R1910 B.n423 B.n422 10.6151
R1911 B.n572 B.n374 10.6151
R1912 B.n573 B.n572 10.6151
R1913 B.n574 B.n573 10.6151
R1914 B.n574 B.n365 10.6151
R1915 B.n584 B.n365 10.6151
R1916 B.n585 B.n584 10.6151
R1917 B.n586 B.n585 10.6151
R1918 B.n586 B.n358 10.6151
R1919 B.n596 B.n358 10.6151
R1920 B.n597 B.n596 10.6151
R1921 B.n598 B.n597 10.6151
R1922 B.n598 B.n350 10.6151
R1923 B.n608 B.n350 10.6151
R1924 B.n609 B.n608 10.6151
R1925 B.n610 B.n609 10.6151
R1926 B.n610 B.n342 10.6151
R1927 B.n620 B.n342 10.6151
R1928 B.n621 B.n620 10.6151
R1929 B.n622 B.n621 10.6151
R1930 B.n622 B.n334 10.6151
R1931 B.n632 B.n334 10.6151
R1932 B.n633 B.n632 10.6151
R1933 B.n634 B.n633 10.6151
R1934 B.n634 B.n327 10.6151
R1935 B.n645 B.n327 10.6151
R1936 B.n646 B.n645 10.6151
R1937 B.n647 B.n646 10.6151
R1938 B.n647 B.n319 10.6151
R1939 B.n657 B.n319 10.6151
R1940 B.n658 B.n657 10.6151
R1941 B.n659 B.n658 10.6151
R1942 B.n659 B.n311 10.6151
R1943 B.n669 B.n311 10.6151
R1944 B.n670 B.n669 10.6151
R1945 B.n671 B.n670 10.6151
R1946 B.n671 B.n303 10.6151
R1947 B.n681 B.n303 10.6151
R1948 B.n682 B.n681 10.6151
R1949 B.n683 B.n682 10.6151
R1950 B.n683 B.n295 10.6151
R1951 B.n692 B.n295 10.6151
R1952 B.n693 B.n692 10.6151
R1953 B.n694 B.n693 10.6151
R1954 B.n694 B.n286 10.6151
R1955 B.n704 B.n286 10.6151
R1956 B.n705 B.n704 10.6151
R1957 B.n707 B.n705 10.6151
R1958 B.n707 B.n706 10.6151
R1959 B.n706 B.n279 10.6151
R1960 B.n718 B.n279 10.6151
R1961 B.n719 B.n718 10.6151
R1962 B.n720 B.n719 10.6151
R1963 B.n721 B.n720 10.6151
R1964 B.n722 B.n721 10.6151
R1965 B.n725 B.n722 10.6151
R1966 B.n726 B.n725 10.6151
R1967 B.n727 B.n726 10.6151
R1968 B.n728 B.n727 10.6151
R1969 B.n730 B.n728 10.6151
R1970 B.n731 B.n730 10.6151
R1971 B.n732 B.n731 10.6151
R1972 B.n733 B.n732 10.6151
R1973 B.n735 B.n733 10.6151
R1974 B.n736 B.n735 10.6151
R1975 B.n737 B.n736 10.6151
R1976 B.n738 B.n737 10.6151
R1977 B.n740 B.n738 10.6151
R1978 B.n741 B.n740 10.6151
R1979 B.n742 B.n741 10.6151
R1980 B.n743 B.n742 10.6151
R1981 B.n745 B.n743 10.6151
R1982 B.n746 B.n745 10.6151
R1983 B.n747 B.n746 10.6151
R1984 B.n748 B.n747 10.6151
R1985 B.n750 B.n748 10.6151
R1986 B.n751 B.n750 10.6151
R1987 B.n752 B.n751 10.6151
R1988 B.n753 B.n752 10.6151
R1989 B.n755 B.n753 10.6151
R1990 B.n756 B.n755 10.6151
R1991 B.n757 B.n756 10.6151
R1992 B.n758 B.n757 10.6151
R1993 B.n760 B.n758 10.6151
R1994 B.n761 B.n760 10.6151
R1995 B.n762 B.n761 10.6151
R1996 B.n763 B.n762 10.6151
R1997 B.n765 B.n763 10.6151
R1998 B.n766 B.n765 10.6151
R1999 B.n767 B.n766 10.6151
R2000 B.n768 B.n767 10.6151
R2001 B.n770 B.n768 10.6151
R2002 B.n771 B.n770 10.6151
R2003 B.n772 B.n771 10.6151
R2004 B.n773 B.n772 10.6151
R2005 B.n775 B.n773 10.6151
R2006 B.n776 B.n775 10.6151
R2007 B.n777 B.n776 10.6151
R2008 B.n778 B.n777 10.6151
R2009 B.n780 B.n778 10.6151
R2010 B.n781 B.n780 10.6151
R2011 B.n782 B.n781 10.6151
R2012 B.n783 B.n782 10.6151
R2013 B.n784 B.n783 10.6151
R2014 B.n887 B.n1 10.6151
R2015 B.n887 B.n886 10.6151
R2016 B.n886 B.n885 10.6151
R2017 B.n885 B.n10 10.6151
R2018 B.n879 B.n10 10.6151
R2019 B.n879 B.n878 10.6151
R2020 B.n878 B.n877 10.6151
R2021 B.n877 B.n18 10.6151
R2022 B.n871 B.n18 10.6151
R2023 B.n871 B.n870 10.6151
R2024 B.n870 B.n869 10.6151
R2025 B.n869 B.n25 10.6151
R2026 B.n864 B.n25 10.6151
R2027 B.n864 B.n863 10.6151
R2028 B.n863 B.n862 10.6151
R2029 B.n862 B.n32 10.6151
R2030 B.n856 B.n32 10.6151
R2031 B.n856 B.n855 10.6151
R2032 B.n855 B.n854 10.6151
R2033 B.n854 B.n39 10.6151
R2034 B.n848 B.n39 10.6151
R2035 B.n848 B.n847 10.6151
R2036 B.n847 B.n846 10.6151
R2037 B.n846 B.n46 10.6151
R2038 B.n840 B.n46 10.6151
R2039 B.n840 B.n839 10.6151
R2040 B.n839 B.n838 10.6151
R2041 B.n838 B.n52 10.6151
R2042 B.n832 B.n52 10.6151
R2043 B.n832 B.n831 10.6151
R2044 B.n831 B.n830 10.6151
R2045 B.n830 B.n60 10.6151
R2046 B.n824 B.n60 10.6151
R2047 B.n824 B.n823 10.6151
R2048 B.n823 B.n822 10.6151
R2049 B.n822 B.n67 10.6151
R2050 B.n816 B.n67 10.6151
R2051 B.n816 B.n815 10.6151
R2052 B.n815 B.n814 10.6151
R2053 B.n814 B.n74 10.6151
R2054 B.n808 B.n74 10.6151
R2055 B.n808 B.n807 10.6151
R2056 B.n807 B.n806 10.6151
R2057 B.n806 B.n81 10.6151
R2058 B.n800 B.n81 10.6151
R2059 B.n800 B.n799 10.6151
R2060 B.n799 B.n798 10.6151
R2061 B.n798 B.n88 10.6151
R2062 B.n792 B.n88 10.6151
R2063 B.n792 B.n791 10.6151
R2064 B.n790 B.n95 10.6151
R2065 B.n140 B.n95 10.6151
R2066 B.n141 B.n140 10.6151
R2067 B.n144 B.n141 10.6151
R2068 B.n145 B.n144 10.6151
R2069 B.n148 B.n145 10.6151
R2070 B.n149 B.n148 10.6151
R2071 B.n152 B.n149 10.6151
R2072 B.n153 B.n152 10.6151
R2073 B.n156 B.n153 10.6151
R2074 B.n157 B.n156 10.6151
R2075 B.n160 B.n157 10.6151
R2076 B.n161 B.n160 10.6151
R2077 B.n164 B.n161 10.6151
R2078 B.n165 B.n164 10.6151
R2079 B.n168 B.n165 10.6151
R2080 B.n169 B.n168 10.6151
R2081 B.n172 B.n169 10.6151
R2082 B.n173 B.n172 10.6151
R2083 B.n176 B.n173 10.6151
R2084 B.n177 B.n176 10.6151
R2085 B.n180 B.n177 10.6151
R2086 B.n181 B.n180 10.6151
R2087 B.n184 B.n181 10.6151
R2088 B.n185 B.n184 10.6151
R2089 B.n188 B.n185 10.6151
R2090 B.n189 B.n188 10.6151
R2091 B.n192 B.n189 10.6151
R2092 B.n193 B.n192 10.6151
R2093 B.n196 B.n193 10.6151
R2094 B.n197 B.n196 10.6151
R2095 B.n201 B.n200 10.6151
R2096 B.n204 B.n201 10.6151
R2097 B.n205 B.n204 10.6151
R2098 B.n208 B.n205 10.6151
R2099 B.n209 B.n208 10.6151
R2100 B.n212 B.n209 10.6151
R2101 B.n213 B.n212 10.6151
R2102 B.n216 B.n213 10.6151
R2103 B.n221 B.n218 10.6151
R2104 B.n222 B.n221 10.6151
R2105 B.n225 B.n222 10.6151
R2106 B.n226 B.n225 10.6151
R2107 B.n229 B.n226 10.6151
R2108 B.n230 B.n229 10.6151
R2109 B.n233 B.n230 10.6151
R2110 B.n234 B.n233 10.6151
R2111 B.n237 B.n234 10.6151
R2112 B.n238 B.n237 10.6151
R2113 B.n241 B.n238 10.6151
R2114 B.n242 B.n241 10.6151
R2115 B.n245 B.n242 10.6151
R2116 B.n246 B.n245 10.6151
R2117 B.n249 B.n246 10.6151
R2118 B.n250 B.n249 10.6151
R2119 B.n253 B.n250 10.6151
R2120 B.n254 B.n253 10.6151
R2121 B.n257 B.n254 10.6151
R2122 B.n258 B.n257 10.6151
R2123 B.n261 B.n258 10.6151
R2124 B.n262 B.n261 10.6151
R2125 B.n265 B.n262 10.6151
R2126 B.n266 B.n265 10.6151
R2127 B.n269 B.n266 10.6151
R2128 B.n270 B.n269 10.6151
R2129 B.n273 B.n270 10.6151
R2130 B.n274 B.n273 10.6151
R2131 B.n277 B.n274 10.6151
R2132 B.n278 B.n277 10.6151
R2133 B.n785 B.n278 10.6151
R2134 B.n895 B.n0 8.11757
R2135 B.n895 B.n1 8.11757
R2136 B.n503 B.n502 6.5566
R2137 B.n486 B.n420 6.5566
R2138 B.n200 B.n138 6.5566
R2139 B.n217 B.n216 6.5566
R2140 B.n504 B.n503 4.05904
R2141 B.n483 B.n420 4.05904
R2142 B.n197 B.n138 4.05904
R2143 B.n218 B.n217 4.05904
R2144 VN.n63 VN.n33 161.3
R2145 VN.n62 VN.n61 161.3
R2146 VN.n60 VN.n34 161.3
R2147 VN.n59 VN.n58 161.3
R2148 VN.n57 VN.n35 161.3
R2149 VN.n55 VN.n54 161.3
R2150 VN.n53 VN.n36 161.3
R2151 VN.n52 VN.n51 161.3
R2152 VN.n50 VN.n37 161.3
R2153 VN.n49 VN.n48 161.3
R2154 VN.n47 VN.n38 161.3
R2155 VN.n46 VN.n45 161.3
R2156 VN.n44 VN.n39 161.3
R2157 VN.n43 VN.n42 161.3
R2158 VN.n30 VN.n0 161.3
R2159 VN.n29 VN.n28 161.3
R2160 VN.n27 VN.n1 161.3
R2161 VN.n26 VN.n25 161.3
R2162 VN.n24 VN.n2 161.3
R2163 VN.n22 VN.n21 161.3
R2164 VN.n20 VN.n3 161.3
R2165 VN.n19 VN.n18 161.3
R2166 VN.n17 VN.n4 161.3
R2167 VN.n16 VN.n15 161.3
R2168 VN.n14 VN.n5 161.3
R2169 VN.n13 VN.n12 161.3
R2170 VN.n11 VN.n6 161.3
R2171 VN.n10 VN.n9 161.3
R2172 VN.n8 VN.t3 130.905
R2173 VN.n41 VN.t8 130.905
R2174 VN.n16 VN.t0 96.5131
R2175 VN.n7 VN.t6 96.5131
R2176 VN.n23 VN.t5 96.5131
R2177 VN.n31 VN.t9 96.5131
R2178 VN.n49 VN.t7 96.5131
R2179 VN.n40 VN.t1 96.5131
R2180 VN.n56 VN.t2 96.5131
R2181 VN.n64 VN.t4 96.5131
R2182 VN.n32 VN.n31 89.2255
R2183 VN.n65 VN.n64 89.2255
R2184 VN.n12 VN.n11 56.5193
R2185 VN.n18 VN.n3 56.5193
R2186 VN.n29 VN.n1 56.5193
R2187 VN.n45 VN.n44 56.5193
R2188 VN.n51 VN.n36 56.5193
R2189 VN.n62 VN.n34 56.5193
R2190 VN VN.n65 48.3807
R2191 VN.n8 VN.n7 47.6808
R2192 VN.n41 VN.n40 47.6808
R2193 VN.n11 VN.n10 24.4675
R2194 VN.n12 VN.n5 24.4675
R2195 VN.n16 VN.n5 24.4675
R2196 VN.n17 VN.n16 24.4675
R2197 VN.n18 VN.n17 24.4675
R2198 VN.n22 VN.n3 24.4675
R2199 VN.n25 VN.n24 24.4675
R2200 VN.n25 VN.n1 24.4675
R2201 VN.n30 VN.n29 24.4675
R2202 VN.n44 VN.n43 24.4675
R2203 VN.n51 VN.n50 24.4675
R2204 VN.n50 VN.n49 24.4675
R2205 VN.n49 VN.n38 24.4675
R2206 VN.n45 VN.n38 24.4675
R2207 VN.n58 VN.n34 24.4675
R2208 VN.n58 VN.n57 24.4675
R2209 VN.n55 VN.n36 24.4675
R2210 VN.n63 VN.n62 24.4675
R2211 VN.n10 VN.n7 22.9995
R2212 VN.n23 VN.n22 22.9995
R2213 VN.n43 VN.n40 22.9995
R2214 VN.n56 VN.n55 22.9995
R2215 VN.n31 VN.n30 21.5315
R2216 VN.n64 VN.n63 21.5315
R2217 VN.n42 VN.n41 8.82758
R2218 VN.n9 VN.n8 8.82758
R2219 VN.n24 VN.n23 1.46852
R2220 VN.n57 VN.n56 1.46852
R2221 VN.n65 VN.n33 0.278367
R2222 VN.n32 VN.n0 0.278367
R2223 VN.n61 VN.n33 0.189894
R2224 VN.n61 VN.n60 0.189894
R2225 VN.n60 VN.n59 0.189894
R2226 VN.n59 VN.n35 0.189894
R2227 VN.n54 VN.n35 0.189894
R2228 VN.n54 VN.n53 0.189894
R2229 VN.n53 VN.n52 0.189894
R2230 VN.n52 VN.n37 0.189894
R2231 VN.n48 VN.n37 0.189894
R2232 VN.n48 VN.n47 0.189894
R2233 VN.n47 VN.n46 0.189894
R2234 VN.n46 VN.n39 0.189894
R2235 VN.n42 VN.n39 0.189894
R2236 VN.n9 VN.n6 0.189894
R2237 VN.n13 VN.n6 0.189894
R2238 VN.n14 VN.n13 0.189894
R2239 VN.n15 VN.n14 0.189894
R2240 VN.n15 VN.n4 0.189894
R2241 VN.n19 VN.n4 0.189894
R2242 VN.n20 VN.n19 0.189894
R2243 VN.n21 VN.n20 0.189894
R2244 VN.n21 VN.n2 0.189894
R2245 VN.n26 VN.n2 0.189894
R2246 VN.n27 VN.n26 0.189894
R2247 VN.n28 VN.n27 0.189894
R2248 VN.n28 VN.n0 0.189894
R2249 VN VN.n32 0.153454
R2250 VDD2.n89 VDD2.n49 289.615
R2251 VDD2.n40 VDD2.n0 289.615
R2252 VDD2.n90 VDD2.n89 185
R2253 VDD2.n88 VDD2.n87 185
R2254 VDD2.n86 VDD2.n52 185
R2255 VDD2.n56 VDD2.n53 185
R2256 VDD2.n81 VDD2.n80 185
R2257 VDD2.n79 VDD2.n78 185
R2258 VDD2.n58 VDD2.n57 185
R2259 VDD2.n73 VDD2.n72 185
R2260 VDD2.n71 VDD2.n70 185
R2261 VDD2.n62 VDD2.n61 185
R2262 VDD2.n65 VDD2.n64 185
R2263 VDD2.n15 VDD2.n14 185
R2264 VDD2.n12 VDD2.n11 185
R2265 VDD2.n21 VDD2.n20 185
R2266 VDD2.n23 VDD2.n22 185
R2267 VDD2.n8 VDD2.n7 185
R2268 VDD2.n29 VDD2.n28 185
R2269 VDD2.n32 VDD2.n31 185
R2270 VDD2.n30 VDD2.n4 185
R2271 VDD2.n37 VDD2.n3 185
R2272 VDD2.n39 VDD2.n38 185
R2273 VDD2.n41 VDD2.n40 185
R2274 VDD2.t5 VDD2.n63 149.524
R2275 VDD2.t6 VDD2.n13 149.524
R2276 VDD2.n89 VDD2.n88 104.615
R2277 VDD2.n88 VDD2.n52 104.615
R2278 VDD2.n56 VDD2.n52 104.615
R2279 VDD2.n80 VDD2.n56 104.615
R2280 VDD2.n80 VDD2.n79 104.615
R2281 VDD2.n79 VDD2.n57 104.615
R2282 VDD2.n72 VDD2.n57 104.615
R2283 VDD2.n72 VDD2.n71 104.615
R2284 VDD2.n71 VDD2.n61 104.615
R2285 VDD2.n64 VDD2.n61 104.615
R2286 VDD2.n14 VDD2.n11 104.615
R2287 VDD2.n21 VDD2.n11 104.615
R2288 VDD2.n22 VDD2.n21 104.615
R2289 VDD2.n22 VDD2.n7 104.615
R2290 VDD2.n29 VDD2.n7 104.615
R2291 VDD2.n31 VDD2.n29 104.615
R2292 VDD2.n31 VDD2.n30 104.615
R2293 VDD2.n30 VDD2.n3 104.615
R2294 VDD2.n39 VDD2.n3 104.615
R2295 VDD2.n40 VDD2.n39 104.615
R2296 VDD2.n48 VDD2.n47 65.9523
R2297 VDD2 VDD2.n97 65.9495
R2298 VDD2.n96 VDD2.n95 64.4109
R2299 VDD2.n46 VDD2.n45 64.4107
R2300 VDD2.n64 VDD2.t5 52.3082
R2301 VDD2.n14 VDD2.t6 52.3082
R2302 VDD2.n46 VDD2.n44 51.9631
R2303 VDD2.n94 VDD2.n93 49.8338
R2304 VDD2.n94 VDD2.n48 41.2174
R2305 VDD2.n87 VDD2.n86 13.1884
R2306 VDD2.n38 VDD2.n37 13.1884
R2307 VDD2.n90 VDD2.n51 12.8005
R2308 VDD2.n85 VDD2.n53 12.8005
R2309 VDD2.n36 VDD2.n4 12.8005
R2310 VDD2.n41 VDD2.n2 12.8005
R2311 VDD2.n91 VDD2.n49 12.0247
R2312 VDD2.n82 VDD2.n81 12.0247
R2313 VDD2.n33 VDD2.n32 12.0247
R2314 VDD2.n42 VDD2.n0 12.0247
R2315 VDD2.n78 VDD2.n55 11.249
R2316 VDD2.n28 VDD2.n6 11.249
R2317 VDD2.n77 VDD2.n58 10.4732
R2318 VDD2.n27 VDD2.n8 10.4732
R2319 VDD2.n65 VDD2.n63 10.2747
R2320 VDD2.n15 VDD2.n13 10.2747
R2321 VDD2.n74 VDD2.n73 9.69747
R2322 VDD2.n24 VDD2.n23 9.69747
R2323 VDD2.n93 VDD2.n92 9.45567
R2324 VDD2.n44 VDD2.n43 9.45567
R2325 VDD2.n67 VDD2.n66 9.3005
R2326 VDD2.n69 VDD2.n68 9.3005
R2327 VDD2.n60 VDD2.n59 9.3005
R2328 VDD2.n75 VDD2.n74 9.3005
R2329 VDD2.n77 VDD2.n76 9.3005
R2330 VDD2.n55 VDD2.n54 9.3005
R2331 VDD2.n83 VDD2.n82 9.3005
R2332 VDD2.n85 VDD2.n84 9.3005
R2333 VDD2.n92 VDD2.n91 9.3005
R2334 VDD2.n51 VDD2.n50 9.3005
R2335 VDD2.n43 VDD2.n42 9.3005
R2336 VDD2.n2 VDD2.n1 9.3005
R2337 VDD2.n17 VDD2.n16 9.3005
R2338 VDD2.n19 VDD2.n18 9.3005
R2339 VDD2.n10 VDD2.n9 9.3005
R2340 VDD2.n25 VDD2.n24 9.3005
R2341 VDD2.n27 VDD2.n26 9.3005
R2342 VDD2.n6 VDD2.n5 9.3005
R2343 VDD2.n34 VDD2.n33 9.3005
R2344 VDD2.n36 VDD2.n35 9.3005
R2345 VDD2.n70 VDD2.n60 8.92171
R2346 VDD2.n20 VDD2.n10 8.92171
R2347 VDD2.n69 VDD2.n62 8.14595
R2348 VDD2.n19 VDD2.n12 8.14595
R2349 VDD2.n66 VDD2.n65 7.3702
R2350 VDD2.n16 VDD2.n15 7.3702
R2351 VDD2.n66 VDD2.n62 5.81868
R2352 VDD2.n16 VDD2.n12 5.81868
R2353 VDD2.n70 VDD2.n69 5.04292
R2354 VDD2.n20 VDD2.n19 5.04292
R2355 VDD2.n73 VDD2.n60 4.26717
R2356 VDD2.n23 VDD2.n10 4.26717
R2357 VDD2.n74 VDD2.n58 3.49141
R2358 VDD2.n24 VDD2.n8 3.49141
R2359 VDD2.n17 VDD2.n13 2.84303
R2360 VDD2.n67 VDD2.n63 2.84303
R2361 VDD2.n78 VDD2.n77 2.71565
R2362 VDD2.n28 VDD2.n27 2.71565
R2363 VDD2.n97 VDD2.t8 2.31088
R2364 VDD2.n97 VDD2.t1 2.31088
R2365 VDD2.n95 VDD2.t7 2.31088
R2366 VDD2.n95 VDD2.t2 2.31088
R2367 VDD2.n47 VDD2.t4 2.31088
R2368 VDD2.n47 VDD2.t0 2.31088
R2369 VDD2.n45 VDD2.t3 2.31088
R2370 VDD2.n45 VDD2.t9 2.31088
R2371 VDD2.n96 VDD2.n94 2.12981
R2372 VDD2.n93 VDD2.n49 1.93989
R2373 VDD2.n81 VDD2.n55 1.93989
R2374 VDD2.n32 VDD2.n6 1.93989
R2375 VDD2.n44 VDD2.n0 1.93989
R2376 VDD2.n91 VDD2.n90 1.16414
R2377 VDD2.n82 VDD2.n53 1.16414
R2378 VDD2.n33 VDD2.n4 1.16414
R2379 VDD2.n42 VDD2.n41 1.16414
R2380 VDD2 VDD2.n96 0.591017
R2381 VDD2.n48 VDD2.n46 0.477482
R2382 VDD2.n87 VDD2.n51 0.388379
R2383 VDD2.n86 VDD2.n85 0.388379
R2384 VDD2.n37 VDD2.n36 0.388379
R2385 VDD2.n38 VDD2.n2 0.388379
R2386 VDD2.n92 VDD2.n50 0.155672
R2387 VDD2.n84 VDD2.n50 0.155672
R2388 VDD2.n84 VDD2.n83 0.155672
R2389 VDD2.n83 VDD2.n54 0.155672
R2390 VDD2.n76 VDD2.n54 0.155672
R2391 VDD2.n76 VDD2.n75 0.155672
R2392 VDD2.n75 VDD2.n59 0.155672
R2393 VDD2.n68 VDD2.n59 0.155672
R2394 VDD2.n68 VDD2.n67 0.155672
R2395 VDD2.n18 VDD2.n17 0.155672
R2396 VDD2.n18 VDD2.n9 0.155672
R2397 VDD2.n25 VDD2.n9 0.155672
R2398 VDD2.n26 VDD2.n25 0.155672
R2399 VDD2.n26 VDD2.n5 0.155672
R2400 VDD2.n34 VDD2.n5 0.155672
R2401 VDD2.n35 VDD2.n34 0.155672
R2402 VDD2.n35 VDD2.n1 0.155672
R2403 VDD2.n43 VDD2.n1 0.155672
C0 VTAIL VDD1 8.64974f
C1 VN VP 7.08344f
C2 VDD1 VP 7.80726f
C3 VTAIL VP 8.049589f
C4 VN VDD2 7.43816f
C5 VDD1 VDD2 1.87569f
C6 VTAIL VDD2 8.697989f
C7 VN VDD1 0.15246f
C8 VDD2 VP 0.524758f
C9 VN VTAIL 8.03533f
C10 VDD2 B 6.032603f
C11 VDD1 B 6.029297f
C12 VTAIL B 6.506651f
C13 VN B 15.678321f
C14 VP B 14.215964f
C15 VDD2.n0 B 0.029034f
C16 VDD2.n1 B 0.022259f
C17 VDD2.n2 B 0.011961f
C18 VDD2.n3 B 0.028271f
C19 VDD2.n4 B 0.012665f
C20 VDD2.n5 B 0.022259f
C21 VDD2.n6 B 0.011961f
C22 VDD2.n7 B 0.028271f
C23 VDD2.n8 B 0.012665f
C24 VDD2.n9 B 0.022259f
C25 VDD2.n10 B 0.011961f
C26 VDD2.n11 B 0.028271f
C27 VDD2.n12 B 0.012665f
C28 VDD2.n13 B 0.131185f
C29 VDD2.t6 B 0.047344f
C30 VDD2.n14 B 0.021204f
C31 VDD2.n15 B 0.019986f
C32 VDD2.n16 B 0.011961f
C33 VDD2.n17 B 0.783323f
C34 VDD2.n18 B 0.022259f
C35 VDD2.n19 B 0.011961f
C36 VDD2.n20 B 0.012665f
C37 VDD2.n21 B 0.028271f
C38 VDD2.n22 B 0.028271f
C39 VDD2.n23 B 0.012665f
C40 VDD2.n24 B 0.011961f
C41 VDD2.n25 B 0.022259f
C42 VDD2.n26 B 0.022259f
C43 VDD2.n27 B 0.011961f
C44 VDD2.n28 B 0.012665f
C45 VDD2.n29 B 0.028271f
C46 VDD2.n30 B 0.028271f
C47 VDD2.n31 B 0.028271f
C48 VDD2.n32 B 0.012665f
C49 VDD2.n33 B 0.011961f
C50 VDD2.n34 B 0.022259f
C51 VDD2.n35 B 0.022259f
C52 VDD2.n36 B 0.011961f
C53 VDD2.n37 B 0.012313f
C54 VDD2.n38 B 0.012313f
C55 VDD2.n39 B 0.028271f
C56 VDD2.n40 B 0.057219f
C57 VDD2.n41 B 0.012665f
C58 VDD2.n42 B 0.011961f
C59 VDD2.n43 B 0.052971f
C60 VDD2.n44 B 0.055061f
C61 VDD2.t3 B 0.150744f
C62 VDD2.t9 B 0.150744f
C63 VDD2.n45 B 1.31262f
C64 VDD2.n46 B 0.554794f
C65 VDD2.t4 B 0.150744f
C66 VDD2.t0 B 0.150744f
C67 VDD2.n47 B 1.32316f
C68 VDD2.n48 B 2.18156f
C69 VDD2.n49 B 0.029034f
C70 VDD2.n50 B 0.022259f
C71 VDD2.n51 B 0.011961f
C72 VDD2.n52 B 0.028271f
C73 VDD2.n53 B 0.012665f
C74 VDD2.n54 B 0.022259f
C75 VDD2.n55 B 0.011961f
C76 VDD2.n56 B 0.028271f
C77 VDD2.n57 B 0.028271f
C78 VDD2.n58 B 0.012665f
C79 VDD2.n59 B 0.022259f
C80 VDD2.n60 B 0.011961f
C81 VDD2.n61 B 0.028271f
C82 VDD2.n62 B 0.012665f
C83 VDD2.n63 B 0.131185f
C84 VDD2.t5 B 0.047344f
C85 VDD2.n64 B 0.021204f
C86 VDD2.n65 B 0.019986f
C87 VDD2.n66 B 0.011961f
C88 VDD2.n67 B 0.783323f
C89 VDD2.n68 B 0.022259f
C90 VDD2.n69 B 0.011961f
C91 VDD2.n70 B 0.012665f
C92 VDD2.n71 B 0.028271f
C93 VDD2.n72 B 0.028271f
C94 VDD2.n73 B 0.012665f
C95 VDD2.n74 B 0.011961f
C96 VDD2.n75 B 0.022259f
C97 VDD2.n76 B 0.022259f
C98 VDD2.n77 B 0.011961f
C99 VDD2.n78 B 0.012665f
C100 VDD2.n79 B 0.028271f
C101 VDD2.n80 B 0.028271f
C102 VDD2.n81 B 0.012665f
C103 VDD2.n82 B 0.011961f
C104 VDD2.n83 B 0.022259f
C105 VDD2.n84 B 0.022259f
C106 VDD2.n85 B 0.011961f
C107 VDD2.n86 B 0.012313f
C108 VDD2.n87 B 0.012313f
C109 VDD2.n88 B 0.028271f
C110 VDD2.n89 B 0.057219f
C111 VDD2.n90 B 0.012665f
C112 VDD2.n91 B 0.011961f
C113 VDD2.n92 B 0.052971f
C114 VDD2.n93 B 0.047011f
C115 VDD2.n94 B 2.17735f
C116 VDD2.t7 B 0.150744f
C117 VDD2.t2 B 0.150744f
C118 VDD2.n95 B 1.31262f
C119 VDD2.n96 B 0.373446f
C120 VDD2.t8 B 0.150744f
C121 VDD2.t1 B 0.150744f
C122 VDD2.n97 B 1.32313f
C123 VN.n0 B 0.033068f
C124 VN.t9 B 1.23899f
C125 VN.n1 B 0.033472f
C126 VN.n2 B 0.025082f
C127 VN.t5 B 1.23899f
C128 VN.n3 B 0.037666f
C129 VN.n4 B 0.025082f
C130 VN.t0 B 1.23899f
C131 VN.n5 B 0.046747f
C132 VN.n6 B 0.025082f
C133 VN.t6 B 1.23899f
C134 VN.n7 B 0.527173f
C135 VN.t3 B 1.39445f
C136 VN.n8 B 0.506015f
C137 VN.n9 B 0.21183f
C138 VN.n10 B 0.045362f
C139 VN.n11 B 0.037666f
C140 VN.n12 B 0.035569f
C141 VN.n13 B 0.025082f
C142 VN.n14 B 0.025082f
C143 VN.n15 B 0.025082f
C144 VN.n16 B 0.476459f
C145 VN.n17 B 0.046747f
C146 VN.n18 B 0.035569f
C147 VN.n19 B 0.025082f
C148 VN.n20 B 0.025082f
C149 VN.n21 B 0.025082f
C150 VN.n22 B 0.045362f
C151 VN.n23 B 0.452791f
C152 VN.n24 B 0.025052f
C153 VN.n25 B 0.046747f
C154 VN.n26 B 0.025082f
C155 VN.n27 B 0.025082f
C156 VN.n28 B 0.025082f
C157 VN.n29 B 0.039763f
C158 VN.n30 B 0.043977f
C159 VN.n31 B 0.537768f
C160 VN.n32 B 0.029601f
C161 VN.n33 B 0.033068f
C162 VN.t4 B 1.23899f
C163 VN.n34 B 0.033472f
C164 VN.n35 B 0.025082f
C165 VN.t2 B 1.23899f
C166 VN.n36 B 0.037666f
C167 VN.n37 B 0.025082f
C168 VN.t7 B 1.23899f
C169 VN.n38 B 0.046747f
C170 VN.n39 B 0.025082f
C171 VN.t1 B 1.23899f
C172 VN.n40 B 0.527173f
C173 VN.t8 B 1.39445f
C174 VN.n41 B 0.506015f
C175 VN.n42 B 0.21183f
C176 VN.n43 B 0.045362f
C177 VN.n44 B 0.037666f
C178 VN.n45 B 0.035569f
C179 VN.n46 B 0.025082f
C180 VN.n47 B 0.025082f
C181 VN.n48 B 0.025082f
C182 VN.n49 B 0.476459f
C183 VN.n50 B 0.046747f
C184 VN.n51 B 0.035569f
C185 VN.n52 B 0.025082f
C186 VN.n53 B 0.025082f
C187 VN.n54 B 0.025082f
C188 VN.n55 B 0.045362f
C189 VN.n56 B 0.452791f
C190 VN.n57 B 0.025052f
C191 VN.n58 B 0.046747f
C192 VN.n59 B 0.025082f
C193 VN.n60 B 0.025082f
C194 VN.n61 B 0.025082f
C195 VN.n62 B 0.039763f
C196 VN.n63 B 0.043977f
C197 VN.n64 B 0.537768f
C198 VN.n65 B 1.32034f
C199 VDD1.n0 B 0.029425f
C200 VDD1.n1 B 0.022559f
C201 VDD1.n2 B 0.012122f
C202 VDD1.n3 B 0.028652f
C203 VDD1.n4 B 0.012835f
C204 VDD1.n5 B 0.022559f
C205 VDD1.n6 B 0.012122f
C206 VDD1.n7 B 0.028652f
C207 VDD1.n8 B 0.028652f
C208 VDD1.n9 B 0.012835f
C209 VDD1.n10 B 0.022559f
C210 VDD1.n11 B 0.012122f
C211 VDD1.n12 B 0.028652f
C212 VDD1.n13 B 0.012835f
C213 VDD1.n14 B 0.13295f
C214 VDD1.t7 B 0.047981f
C215 VDD1.n15 B 0.021489f
C216 VDD1.n16 B 0.020255f
C217 VDD1.n17 B 0.012122f
C218 VDD1.n18 B 0.793866f
C219 VDD1.n19 B 0.022559f
C220 VDD1.n20 B 0.012122f
C221 VDD1.n21 B 0.012835f
C222 VDD1.n22 B 0.028652f
C223 VDD1.n23 B 0.028652f
C224 VDD1.n24 B 0.012835f
C225 VDD1.n25 B 0.012122f
C226 VDD1.n26 B 0.022559f
C227 VDD1.n27 B 0.022559f
C228 VDD1.n28 B 0.012122f
C229 VDD1.n29 B 0.012835f
C230 VDD1.n30 B 0.028652f
C231 VDD1.n31 B 0.028652f
C232 VDD1.n32 B 0.012835f
C233 VDD1.n33 B 0.012122f
C234 VDD1.n34 B 0.022559f
C235 VDD1.n35 B 0.022559f
C236 VDD1.n36 B 0.012122f
C237 VDD1.n37 B 0.012478f
C238 VDD1.n38 B 0.012478f
C239 VDD1.n39 B 0.028652f
C240 VDD1.n40 B 0.057989f
C241 VDD1.n41 B 0.012835f
C242 VDD1.n42 B 0.012122f
C243 VDD1.n43 B 0.053684f
C244 VDD1.n44 B 0.055802f
C245 VDD1.t4 B 0.152773f
C246 VDD1.t9 B 0.152773f
C247 VDD1.n45 B 1.33029f
C248 VDD1.n46 B 0.569411f
C249 VDD1.n47 B 0.029425f
C250 VDD1.n48 B 0.022559f
C251 VDD1.n49 B 0.012122f
C252 VDD1.n50 B 0.028652f
C253 VDD1.n51 B 0.012835f
C254 VDD1.n52 B 0.022559f
C255 VDD1.n53 B 0.012122f
C256 VDD1.n54 B 0.028652f
C257 VDD1.n55 B 0.012835f
C258 VDD1.n56 B 0.022559f
C259 VDD1.n57 B 0.012122f
C260 VDD1.n58 B 0.028652f
C261 VDD1.n59 B 0.012835f
C262 VDD1.n60 B 0.13295f
C263 VDD1.t0 B 0.047981f
C264 VDD1.n61 B 0.021489f
C265 VDD1.n62 B 0.020255f
C266 VDD1.n63 B 0.012122f
C267 VDD1.n64 B 0.793866f
C268 VDD1.n65 B 0.022559f
C269 VDD1.n66 B 0.012122f
C270 VDD1.n67 B 0.012835f
C271 VDD1.n68 B 0.028652f
C272 VDD1.n69 B 0.028652f
C273 VDD1.n70 B 0.012835f
C274 VDD1.n71 B 0.012122f
C275 VDD1.n72 B 0.022559f
C276 VDD1.n73 B 0.022559f
C277 VDD1.n74 B 0.012122f
C278 VDD1.n75 B 0.012835f
C279 VDD1.n76 B 0.028652f
C280 VDD1.n77 B 0.028652f
C281 VDD1.n78 B 0.028652f
C282 VDD1.n79 B 0.012835f
C283 VDD1.n80 B 0.012122f
C284 VDD1.n81 B 0.022559f
C285 VDD1.n82 B 0.022559f
C286 VDD1.n83 B 0.012122f
C287 VDD1.n84 B 0.012478f
C288 VDD1.n85 B 0.012478f
C289 VDD1.n86 B 0.028652f
C290 VDD1.n87 B 0.057989f
C291 VDD1.n88 B 0.012835f
C292 VDD1.n89 B 0.012122f
C293 VDD1.n90 B 0.053684f
C294 VDD1.n91 B 0.055802f
C295 VDD1.t5 B 0.152773f
C296 VDD1.t1 B 0.152773f
C297 VDD1.n92 B 1.33028f
C298 VDD1.n93 B 0.562261f
C299 VDD1.t2 B 0.152773f
C300 VDD1.t8 B 0.152773f
C301 VDD1.n94 B 1.34096f
C302 VDD1.n95 B 2.31063f
C303 VDD1.t6 B 0.152773f
C304 VDD1.t3 B 0.152773f
C305 VDD1.n96 B 1.33028f
C306 VDD1.n97 B 2.44766f
C307 VTAIL.t2 B 0.174818f
C308 VTAIL.t0 B 0.174818f
C309 VTAIL.n0 B 1.45167f
C310 VTAIL.n1 B 0.507652f
C311 VTAIL.n2 B 0.033671f
C312 VTAIL.n3 B 0.025814f
C313 VTAIL.n4 B 0.013871f
C314 VTAIL.n5 B 0.032786f
C315 VTAIL.n6 B 0.014687f
C316 VTAIL.n7 B 0.025814f
C317 VTAIL.n8 B 0.013871f
C318 VTAIL.n9 B 0.032786f
C319 VTAIL.n10 B 0.014687f
C320 VTAIL.n11 B 0.025814f
C321 VTAIL.n12 B 0.013871f
C322 VTAIL.n13 B 0.032786f
C323 VTAIL.n14 B 0.014687f
C324 VTAIL.n15 B 0.152135f
C325 VTAIL.t12 B 0.054905f
C326 VTAIL.n16 B 0.02459f
C327 VTAIL.n17 B 0.023177f
C328 VTAIL.n18 B 0.013871f
C329 VTAIL.n19 B 0.908419f
C330 VTAIL.n20 B 0.025814f
C331 VTAIL.n21 B 0.013871f
C332 VTAIL.n22 B 0.014687f
C333 VTAIL.n23 B 0.032786f
C334 VTAIL.n24 B 0.032786f
C335 VTAIL.n25 B 0.014687f
C336 VTAIL.n26 B 0.013871f
C337 VTAIL.n27 B 0.025814f
C338 VTAIL.n28 B 0.025814f
C339 VTAIL.n29 B 0.013871f
C340 VTAIL.n30 B 0.014687f
C341 VTAIL.n31 B 0.032786f
C342 VTAIL.n32 B 0.032786f
C343 VTAIL.n33 B 0.032786f
C344 VTAIL.n34 B 0.014687f
C345 VTAIL.n35 B 0.013871f
C346 VTAIL.n36 B 0.025814f
C347 VTAIL.n37 B 0.025814f
C348 VTAIL.n38 B 0.013871f
C349 VTAIL.n39 B 0.014279f
C350 VTAIL.n40 B 0.014279f
C351 VTAIL.n41 B 0.032786f
C352 VTAIL.n42 B 0.066357f
C353 VTAIL.n43 B 0.014687f
C354 VTAIL.n44 B 0.013871f
C355 VTAIL.n45 B 0.061431f
C356 VTAIL.n46 B 0.036708f
C357 VTAIL.n47 B 0.327788f
C358 VTAIL.t11 B 0.174818f
C359 VTAIL.t14 B 0.174818f
C360 VTAIL.n48 B 1.45167f
C361 VTAIL.n49 B 0.596566f
C362 VTAIL.t15 B 0.174818f
C363 VTAIL.t18 B 0.174818f
C364 VTAIL.n50 B 1.45167f
C365 VTAIL.n51 B 1.73884f
C366 VTAIL.t1 B 0.174818f
C367 VTAIL.t6 B 0.174818f
C368 VTAIL.n52 B 1.45168f
C369 VTAIL.n53 B 1.73883f
C370 VTAIL.t4 B 0.174818f
C371 VTAIL.t3 B 0.174818f
C372 VTAIL.n54 B 1.45168f
C373 VTAIL.n55 B 0.596557f
C374 VTAIL.n56 B 0.033671f
C375 VTAIL.n57 B 0.025814f
C376 VTAIL.n58 B 0.013871f
C377 VTAIL.n59 B 0.032786f
C378 VTAIL.n60 B 0.014687f
C379 VTAIL.n61 B 0.025814f
C380 VTAIL.n62 B 0.013871f
C381 VTAIL.n63 B 0.032786f
C382 VTAIL.n64 B 0.032786f
C383 VTAIL.n65 B 0.014687f
C384 VTAIL.n66 B 0.025814f
C385 VTAIL.n67 B 0.013871f
C386 VTAIL.n68 B 0.032786f
C387 VTAIL.n69 B 0.014687f
C388 VTAIL.n70 B 0.152135f
C389 VTAIL.t9 B 0.054905f
C390 VTAIL.n71 B 0.02459f
C391 VTAIL.n72 B 0.023177f
C392 VTAIL.n73 B 0.013871f
C393 VTAIL.n74 B 0.908419f
C394 VTAIL.n75 B 0.025814f
C395 VTAIL.n76 B 0.013871f
C396 VTAIL.n77 B 0.014687f
C397 VTAIL.n78 B 0.032786f
C398 VTAIL.n79 B 0.032786f
C399 VTAIL.n80 B 0.014687f
C400 VTAIL.n81 B 0.013871f
C401 VTAIL.n82 B 0.025814f
C402 VTAIL.n83 B 0.025814f
C403 VTAIL.n84 B 0.013871f
C404 VTAIL.n85 B 0.014687f
C405 VTAIL.n86 B 0.032786f
C406 VTAIL.n87 B 0.032786f
C407 VTAIL.n88 B 0.014687f
C408 VTAIL.n89 B 0.013871f
C409 VTAIL.n90 B 0.025814f
C410 VTAIL.n91 B 0.025814f
C411 VTAIL.n92 B 0.013871f
C412 VTAIL.n93 B 0.014279f
C413 VTAIL.n94 B 0.014279f
C414 VTAIL.n95 B 0.032786f
C415 VTAIL.n96 B 0.066357f
C416 VTAIL.n97 B 0.014687f
C417 VTAIL.n98 B 0.013871f
C418 VTAIL.n99 B 0.061431f
C419 VTAIL.n100 B 0.036708f
C420 VTAIL.n101 B 0.327788f
C421 VTAIL.t10 B 0.174818f
C422 VTAIL.t17 B 0.174818f
C423 VTAIL.n102 B 1.45168f
C424 VTAIL.n103 B 0.547081f
C425 VTAIL.t19 B 0.174818f
C426 VTAIL.t16 B 0.174818f
C427 VTAIL.n104 B 1.45168f
C428 VTAIL.n105 B 0.596557f
C429 VTAIL.n106 B 0.033671f
C430 VTAIL.n107 B 0.025814f
C431 VTAIL.n108 B 0.013871f
C432 VTAIL.n109 B 0.032786f
C433 VTAIL.n110 B 0.014687f
C434 VTAIL.n111 B 0.025814f
C435 VTAIL.n112 B 0.013871f
C436 VTAIL.n113 B 0.032786f
C437 VTAIL.n114 B 0.032786f
C438 VTAIL.n115 B 0.014687f
C439 VTAIL.n116 B 0.025814f
C440 VTAIL.n117 B 0.013871f
C441 VTAIL.n118 B 0.032786f
C442 VTAIL.n119 B 0.014687f
C443 VTAIL.n120 B 0.152135f
C444 VTAIL.t13 B 0.054905f
C445 VTAIL.n121 B 0.02459f
C446 VTAIL.n122 B 0.023177f
C447 VTAIL.n123 B 0.013871f
C448 VTAIL.n124 B 0.908419f
C449 VTAIL.n125 B 0.025814f
C450 VTAIL.n126 B 0.013871f
C451 VTAIL.n127 B 0.014687f
C452 VTAIL.n128 B 0.032786f
C453 VTAIL.n129 B 0.032786f
C454 VTAIL.n130 B 0.014687f
C455 VTAIL.n131 B 0.013871f
C456 VTAIL.n132 B 0.025814f
C457 VTAIL.n133 B 0.025814f
C458 VTAIL.n134 B 0.013871f
C459 VTAIL.n135 B 0.014687f
C460 VTAIL.n136 B 0.032786f
C461 VTAIL.n137 B 0.032786f
C462 VTAIL.n138 B 0.014687f
C463 VTAIL.n139 B 0.013871f
C464 VTAIL.n140 B 0.025814f
C465 VTAIL.n141 B 0.025814f
C466 VTAIL.n142 B 0.013871f
C467 VTAIL.n143 B 0.014279f
C468 VTAIL.n144 B 0.014279f
C469 VTAIL.n145 B 0.032786f
C470 VTAIL.n146 B 0.066357f
C471 VTAIL.n147 B 0.014687f
C472 VTAIL.n148 B 0.013871f
C473 VTAIL.n149 B 0.061431f
C474 VTAIL.n150 B 0.036708f
C475 VTAIL.n151 B 1.34243f
C476 VTAIL.n152 B 0.033671f
C477 VTAIL.n153 B 0.025814f
C478 VTAIL.n154 B 0.013871f
C479 VTAIL.n155 B 0.032786f
C480 VTAIL.n156 B 0.014687f
C481 VTAIL.n157 B 0.025814f
C482 VTAIL.n158 B 0.013871f
C483 VTAIL.n159 B 0.032786f
C484 VTAIL.n160 B 0.014687f
C485 VTAIL.n161 B 0.025814f
C486 VTAIL.n162 B 0.013871f
C487 VTAIL.n163 B 0.032786f
C488 VTAIL.n164 B 0.014687f
C489 VTAIL.n165 B 0.152135f
C490 VTAIL.t7 B 0.054905f
C491 VTAIL.n166 B 0.02459f
C492 VTAIL.n167 B 0.023177f
C493 VTAIL.n168 B 0.013871f
C494 VTAIL.n169 B 0.908419f
C495 VTAIL.n170 B 0.025814f
C496 VTAIL.n171 B 0.013871f
C497 VTAIL.n172 B 0.014687f
C498 VTAIL.n173 B 0.032786f
C499 VTAIL.n174 B 0.032786f
C500 VTAIL.n175 B 0.014687f
C501 VTAIL.n176 B 0.013871f
C502 VTAIL.n177 B 0.025814f
C503 VTAIL.n178 B 0.025814f
C504 VTAIL.n179 B 0.013871f
C505 VTAIL.n180 B 0.014687f
C506 VTAIL.n181 B 0.032786f
C507 VTAIL.n182 B 0.032786f
C508 VTAIL.n183 B 0.032786f
C509 VTAIL.n184 B 0.014687f
C510 VTAIL.n185 B 0.013871f
C511 VTAIL.n186 B 0.025814f
C512 VTAIL.n187 B 0.025814f
C513 VTAIL.n188 B 0.013871f
C514 VTAIL.n189 B 0.014279f
C515 VTAIL.n190 B 0.014279f
C516 VTAIL.n191 B 0.032786f
C517 VTAIL.n192 B 0.066357f
C518 VTAIL.n193 B 0.014687f
C519 VTAIL.n194 B 0.013871f
C520 VTAIL.n195 B 0.061431f
C521 VTAIL.n196 B 0.036708f
C522 VTAIL.n197 B 1.34243f
C523 VTAIL.t5 B 0.174818f
C524 VTAIL.t8 B 0.174818f
C525 VTAIL.n198 B 1.45167f
C526 VTAIL.n199 B 0.458893f
C527 VP.n0 B 0.033709f
C528 VP.t1 B 1.263f
C529 VP.n1 B 0.034121f
C530 VP.n2 B 0.025568f
C531 VP.t7 B 1.263f
C532 VP.n3 B 0.038396f
C533 VP.n4 B 0.025568f
C534 VP.t8 B 1.263f
C535 VP.n5 B 0.047652f
C536 VP.n6 B 0.025568f
C537 VP.t4 B 1.263f
C538 VP.n7 B 0.461564f
C539 VP.n8 B 0.025568f
C540 VP.n9 B 0.040533f
C541 VP.n10 B 0.033709f
C542 VP.t6 B 1.263f
C543 VP.n11 B 0.034121f
C544 VP.n12 B 0.025568f
C545 VP.t3 B 1.263f
C546 VP.n13 B 0.038396f
C547 VP.n14 B 0.025568f
C548 VP.t0 B 1.263f
C549 VP.n15 B 0.047652f
C550 VP.n16 B 0.025568f
C551 VP.t5 B 1.263f
C552 VP.n17 B 0.537387f
C553 VP.t2 B 1.42147f
C554 VP.n18 B 0.515819f
C555 VP.n19 B 0.215934f
C556 VP.n20 B 0.046241f
C557 VP.n21 B 0.038396f
C558 VP.n22 B 0.036258f
C559 VP.n23 B 0.025568f
C560 VP.n24 B 0.025568f
C561 VP.n25 B 0.025568f
C562 VP.n26 B 0.48569f
C563 VP.n27 B 0.047652f
C564 VP.n28 B 0.036258f
C565 VP.n29 B 0.025568f
C566 VP.n30 B 0.025568f
C567 VP.n31 B 0.025568f
C568 VP.n32 B 0.046241f
C569 VP.n33 B 0.461564f
C570 VP.n34 B 0.025538f
C571 VP.n35 B 0.047652f
C572 VP.n36 B 0.025568f
C573 VP.n37 B 0.025568f
C574 VP.n38 B 0.025568f
C575 VP.n39 B 0.040533f
C576 VP.n40 B 0.044829f
C577 VP.n41 B 0.548187f
C578 VP.n42 B 1.33209f
C579 VP.n43 B 1.3512f
C580 VP.t9 B 1.263f
C581 VP.n44 B 0.548187f
C582 VP.n45 B 0.044829f
C583 VP.n46 B 0.033709f
C584 VP.n47 B 0.025568f
C585 VP.n48 B 0.025568f
C586 VP.n49 B 0.034121f
C587 VP.n50 B 0.047652f
C588 VP.n51 B 0.025538f
C589 VP.n52 B 0.025568f
C590 VP.n53 B 0.025568f
C591 VP.n54 B 0.046241f
C592 VP.n55 B 0.038396f
C593 VP.n56 B 0.036258f
C594 VP.n57 B 0.025568f
C595 VP.n58 B 0.025568f
C596 VP.n59 B 0.025568f
C597 VP.n60 B 0.48569f
C598 VP.n61 B 0.047652f
C599 VP.n62 B 0.036258f
C600 VP.n63 B 0.025568f
C601 VP.n64 B 0.025568f
C602 VP.n65 B 0.025568f
C603 VP.n66 B 0.046241f
C604 VP.n67 B 0.461564f
C605 VP.n68 B 0.025538f
C606 VP.n69 B 0.047652f
C607 VP.n70 B 0.025568f
C608 VP.n71 B 0.025568f
C609 VP.n72 B 0.025568f
C610 VP.n73 B 0.040533f
C611 VP.n74 B 0.044829f
C612 VP.n75 B 0.548187f
C613 VP.n76 B 0.030175f
.ends

