* NGSPICE file created from diff_pair_sample_1419.ext - technology: sky130A

.subckt diff_pair_sample_1419 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=6.7821 ps=35.56 w=17.39 l=2.94
X1 VTAIL.t1 VN.t0 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X2 VTAIL.t0 VN.t1 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X3 VTAIL.t13 VP.t1 VDD1.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X4 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X5 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=0 ps=0 w=17.39 l=2.94
X6 VTAIL.t19 VN.t3 VDD2.t6 B.t23 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X7 VDD2.t5 VN.t4 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=2.86935 ps=17.72 w=17.39 l=2.94
X8 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X9 VDD2.t3 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=6.7821 ps=35.56 w=17.39 l=2.94
X10 VTAIL.t17 VP.t2 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X11 VDD1.t6 VP.t3 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=6.7821 ps=35.56 w=17.39 l=2.94
X12 VDD1.t5 VP.t4 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X13 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=2.86935 ps=17.72 w=17.39 l=2.94
X14 VTAIL.t16 VP.t5 VDD1.t4 B.t23 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X15 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=0 ps=0 w=17.39 l=2.94
X16 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=6.7821 ps=35.56 w=17.39 l=2.94
X17 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=0 ps=0 w=17.39 l=2.94
X18 VDD1.t3 VP.t6 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=2.86935 ps=17.72 w=17.39 l=2.94
X19 VTAIL.t18 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X20 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=0 ps=0 w=17.39 l=2.94
X21 VDD1.t1 VP.t8 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7821 pd=35.56 as=2.86935 ps=17.72 w=17.39 l=2.94
X22 VDD1.t0 VP.t9 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
X23 VTAIL.t2 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.86935 pd=17.72 as=2.86935 ps=17.72 w=17.39 l=2.94
R0 VP.n24 VP.t6 175.234
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n23 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n22 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n34 VP.n21 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n20 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n19 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n18 161.3
R13 VP.n46 VP.n45 161.3
R14 VP.n47 VP.n17 161.3
R15 VP.n49 VP.n48 161.3
R16 VP.n50 VP.n16 161.3
R17 VP.n52 VP.n51 161.3
R18 VP.n53 VP.n15 161.3
R19 VP.n55 VP.n54 161.3
R20 VP.n56 VP.n14 161.3
R21 VP.n102 VP.n0 161.3
R22 VP.n101 VP.n100 161.3
R23 VP.n99 VP.n1 161.3
R24 VP.n98 VP.n97 161.3
R25 VP.n96 VP.n2 161.3
R26 VP.n95 VP.n94 161.3
R27 VP.n93 VP.n3 161.3
R28 VP.n92 VP.n91 161.3
R29 VP.n89 VP.n4 161.3
R30 VP.n88 VP.n87 161.3
R31 VP.n86 VP.n5 161.3
R32 VP.n85 VP.n84 161.3
R33 VP.n83 VP.n6 161.3
R34 VP.n82 VP.n81 161.3
R35 VP.n80 VP.n7 161.3
R36 VP.n79 VP.n78 161.3
R37 VP.n77 VP.n8 161.3
R38 VP.n76 VP.n75 161.3
R39 VP.n74 VP.n9 161.3
R40 VP.n73 VP.n72 161.3
R41 VP.n70 VP.n10 161.3
R42 VP.n69 VP.n68 161.3
R43 VP.n67 VP.n11 161.3
R44 VP.n66 VP.n65 161.3
R45 VP.n64 VP.n12 161.3
R46 VP.n63 VP.n62 161.3
R47 VP.n61 VP.n13 161.3
R48 VP.n82 VP.t4 142.552
R49 VP.n59 VP.t8 142.552
R50 VP.n71 VP.t7 142.552
R51 VP.n90 VP.t5 142.552
R52 VP.n103 VP.t3 142.552
R53 VP.n36 VP.t9 142.552
R54 VP.n57 VP.t0 142.552
R55 VP.n44 VP.t2 142.552
R56 VP.n25 VP.t1 142.552
R57 VP.n60 VP.n59 108.799
R58 VP.n104 VP.n103 108.799
R59 VP.n58 VP.n57 108.799
R60 VP.n25 VP.n24 60.6237
R61 VP.n60 VP.n58 59.0261
R62 VP.n77 VP.n76 53.6055
R63 VP.n88 VP.n5 53.6055
R64 VP.n42 VP.n19 53.6055
R65 VP.n31 VP.n30 53.6055
R66 VP.n65 VP.n11 49.7204
R67 VP.n97 VP.n96 49.7204
R68 VP.n51 VP.n50 49.7204
R69 VP.n65 VP.n64 31.2664
R70 VP.n97 VP.n1 31.2664
R71 VP.n51 VP.n15 31.2664
R72 VP.n78 VP.n77 27.3813
R73 VP.n84 VP.n5 27.3813
R74 VP.n38 VP.n19 27.3813
R75 VP.n32 VP.n31 27.3813
R76 VP.n63 VP.n13 24.4675
R77 VP.n64 VP.n63 24.4675
R78 VP.n69 VP.n11 24.4675
R79 VP.n70 VP.n69 24.4675
R80 VP.n72 VP.n9 24.4675
R81 VP.n76 VP.n9 24.4675
R82 VP.n78 VP.n7 24.4675
R83 VP.n82 VP.n7 24.4675
R84 VP.n83 VP.n82 24.4675
R85 VP.n84 VP.n83 24.4675
R86 VP.n89 VP.n88 24.4675
R87 VP.n91 VP.n89 24.4675
R88 VP.n95 VP.n3 24.4675
R89 VP.n96 VP.n95 24.4675
R90 VP.n101 VP.n1 24.4675
R91 VP.n102 VP.n101 24.4675
R92 VP.n55 VP.n15 24.4675
R93 VP.n56 VP.n55 24.4675
R94 VP.n43 VP.n42 24.4675
R95 VP.n45 VP.n43 24.4675
R96 VP.n49 VP.n17 24.4675
R97 VP.n50 VP.n49 24.4675
R98 VP.n32 VP.n21 24.4675
R99 VP.n36 VP.n21 24.4675
R100 VP.n37 VP.n36 24.4675
R101 VP.n38 VP.n37 24.4675
R102 VP.n26 VP.n23 24.4675
R103 VP.n30 VP.n23 24.4675
R104 VP.n72 VP.n71 13.2127
R105 VP.n91 VP.n90 13.2127
R106 VP.n45 VP.n44 13.2127
R107 VP.n26 VP.n25 13.2127
R108 VP.n71 VP.n70 11.2553
R109 VP.n90 VP.n3 11.2553
R110 VP.n44 VP.n17 11.2553
R111 VP.n27 VP.n24 5.12434
R112 VP.n59 VP.n13 1.95786
R113 VP.n103 VP.n102 1.95786
R114 VP.n57 VP.n56 1.95786
R115 VP.n58 VP.n14 0.278367
R116 VP.n61 VP.n60 0.278367
R117 VP.n104 VP.n0 0.278367
R118 VP.n28 VP.n27 0.189894
R119 VP.n29 VP.n28 0.189894
R120 VP.n29 VP.n22 0.189894
R121 VP.n33 VP.n22 0.189894
R122 VP.n34 VP.n33 0.189894
R123 VP.n35 VP.n34 0.189894
R124 VP.n35 VP.n20 0.189894
R125 VP.n39 VP.n20 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n18 0.189894
R129 VP.n46 VP.n18 0.189894
R130 VP.n47 VP.n46 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n16 0.189894
R133 VP.n52 VP.n16 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n14 0.189894
R137 VP.n62 VP.n61 0.189894
R138 VP.n62 VP.n12 0.189894
R139 VP.n66 VP.n12 0.189894
R140 VP.n67 VP.n66 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n68 VP.n10 0.189894
R143 VP.n73 VP.n10 0.189894
R144 VP.n74 VP.n73 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n75 VP.n8 0.189894
R147 VP.n79 VP.n8 0.189894
R148 VP.n80 VP.n79 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n81 VP.n6 0.189894
R151 VP.n85 VP.n6 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n87 VP.n4 0.189894
R155 VP.n92 VP.n4 0.189894
R156 VP.n93 VP.n92 0.189894
R157 VP.n94 VP.n93 0.189894
R158 VP.n94 VP.n2 0.189894
R159 VP.n98 VP.n2 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n100 VP.n99 0.189894
R162 VP.n100 VP.n0 0.189894
R163 VP VP.n104 0.153454
R164 VTAIL.n396 VTAIL.n395 289.615
R165 VTAIL.n96 VTAIL.n95 289.615
R166 VTAIL.n300 VTAIL.n299 289.615
R167 VTAIL.n200 VTAIL.n199 289.615
R168 VTAIL.n332 VTAIL.n331 185
R169 VTAIL.n337 VTAIL.n336 185
R170 VTAIL.n339 VTAIL.n338 185
R171 VTAIL.n328 VTAIL.n327 185
R172 VTAIL.n345 VTAIL.n344 185
R173 VTAIL.n347 VTAIL.n346 185
R174 VTAIL.n324 VTAIL.n323 185
R175 VTAIL.n354 VTAIL.n353 185
R176 VTAIL.n355 VTAIL.n322 185
R177 VTAIL.n357 VTAIL.n356 185
R178 VTAIL.n320 VTAIL.n319 185
R179 VTAIL.n363 VTAIL.n362 185
R180 VTAIL.n365 VTAIL.n364 185
R181 VTAIL.n316 VTAIL.n315 185
R182 VTAIL.n371 VTAIL.n370 185
R183 VTAIL.n373 VTAIL.n372 185
R184 VTAIL.n312 VTAIL.n311 185
R185 VTAIL.n379 VTAIL.n378 185
R186 VTAIL.n381 VTAIL.n380 185
R187 VTAIL.n308 VTAIL.n307 185
R188 VTAIL.n387 VTAIL.n386 185
R189 VTAIL.n389 VTAIL.n388 185
R190 VTAIL.n304 VTAIL.n303 185
R191 VTAIL.n395 VTAIL.n394 185
R192 VTAIL.n32 VTAIL.n31 185
R193 VTAIL.n37 VTAIL.n36 185
R194 VTAIL.n39 VTAIL.n38 185
R195 VTAIL.n28 VTAIL.n27 185
R196 VTAIL.n45 VTAIL.n44 185
R197 VTAIL.n47 VTAIL.n46 185
R198 VTAIL.n24 VTAIL.n23 185
R199 VTAIL.n54 VTAIL.n53 185
R200 VTAIL.n55 VTAIL.n22 185
R201 VTAIL.n57 VTAIL.n56 185
R202 VTAIL.n20 VTAIL.n19 185
R203 VTAIL.n63 VTAIL.n62 185
R204 VTAIL.n65 VTAIL.n64 185
R205 VTAIL.n16 VTAIL.n15 185
R206 VTAIL.n71 VTAIL.n70 185
R207 VTAIL.n73 VTAIL.n72 185
R208 VTAIL.n12 VTAIL.n11 185
R209 VTAIL.n79 VTAIL.n78 185
R210 VTAIL.n81 VTAIL.n80 185
R211 VTAIL.n8 VTAIL.n7 185
R212 VTAIL.n87 VTAIL.n86 185
R213 VTAIL.n89 VTAIL.n88 185
R214 VTAIL.n4 VTAIL.n3 185
R215 VTAIL.n95 VTAIL.n94 185
R216 VTAIL.n299 VTAIL.n298 185
R217 VTAIL.n208 VTAIL.n207 185
R218 VTAIL.n293 VTAIL.n292 185
R219 VTAIL.n291 VTAIL.n290 185
R220 VTAIL.n212 VTAIL.n211 185
R221 VTAIL.n285 VTAIL.n284 185
R222 VTAIL.n283 VTAIL.n282 185
R223 VTAIL.n216 VTAIL.n215 185
R224 VTAIL.n277 VTAIL.n276 185
R225 VTAIL.n275 VTAIL.n274 185
R226 VTAIL.n220 VTAIL.n219 185
R227 VTAIL.n269 VTAIL.n268 185
R228 VTAIL.n267 VTAIL.n266 185
R229 VTAIL.n224 VTAIL.n223 185
R230 VTAIL.n261 VTAIL.n260 185
R231 VTAIL.n259 VTAIL.n226 185
R232 VTAIL.n258 VTAIL.n257 185
R233 VTAIL.n229 VTAIL.n227 185
R234 VTAIL.n252 VTAIL.n251 185
R235 VTAIL.n250 VTAIL.n249 185
R236 VTAIL.n233 VTAIL.n232 185
R237 VTAIL.n244 VTAIL.n243 185
R238 VTAIL.n242 VTAIL.n241 185
R239 VTAIL.n237 VTAIL.n236 185
R240 VTAIL.n199 VTAIL.n198 185
R241 VTAIL.n108 VTAIL.n107 185
R242 VTAIL.n193 VTAIL.n192 185
R243 VTAIL.n191 VTAIL.n190 185
R244 VTAIL.n112 VTAIL.n111 185
R245 VTAIL.n185 VTAIL.n184 185
R246 VTAIL.n183 VTAIL.n182 185
R247 VTAIL.n116 VTAIL.n115 185
R248 VTAIL.n177 VTAIL.n176 185
R249 VTAIL.n175 VTAIL.n174 185
R250 VTAIL.n120 VTAIL.n119 185
R251 VTAIL.n169 VTAIL.n168 185
R252 VTAIL.n167 VTAIL.n166 185
R253 VTAIL.n124 VTAIL.n123 185
R254 VTAIL.n161 VTAIL.n160 185
R255 VTAIL.n159 VTAIL.n126 185
R256 VTAIL.n158 VTAIL.n157 185
R257 VTAIL.n129 VTAIL.n127 185
R258 VTAIL.n152 VTAIL.n151 185
R259 VTAIL.n150 VTAIL.n149 185
R260 VTAIL.n133 VTAIL.n132 185
R261 VTAIL.n144 VTAIL.n143 185
R262 VTAIL.n142 VTAIL.n141 185
R263 VTAIL.n137 VTAIL.n136 185
R264 VTAIL.n333 VTAIL.t5 149.524
R265 VTAIL.n33 VTAIL.t10 149.524
R266 VTAIL.n238 VTAIL.t15 149.524
R267 VTAIL.n138 VTAIL.t3 149.524
R268 VTAIL.n337 VTAIL.n331 104.615
R269 VTAIL.n338 VTAIL.n337 104.615
R270 VTAIL.n338 VTAIL.n327 104.615
R271 VTAIL.n345 VTAIL.n327 104.615
R272 VTAIL.n346 VTAIL.n345 104.615
R273 VTAIL.n346 VTAIL.n323 104.615
R274 VTAIL.n354 VTAIL.n323 104.615
R275 VTAIL.n355 VTAIL.n354 104.615
R276 VTAIL.n356 VTAIL.n355 104.615
R277 VTAIL.n356 VTAIL.n319 104.615
R278 VTAIL.n363 VTAIL.n319 104.615
R279 VTAIL.n364 VTAIL.n363 104.615
R280 VTAIL.n364 VTAIL.n315 104.615
R281 VTAIL.n371 VTAIL.n315 104.615
R282 VTAIL.n372 VTAIL.n371 104.615
R283 VTAIL.n372 VTAIL.n311 104.615
R284 VTAIL.n379 VTAIL.n311 104.615
R285 VTAIL.n380 VTAIL.n379 104.615
R286 VTAIL.n380 VTAIL.n307 104.615
R287 VTAIL.n387 VTAIL.n307 104.615
R288 VTAIL.n388 VTAIL.n387 104.615
R289 VTAIL.n388 VTAIL.n303 104.615
R290 VTAIL.n395 VTAIL.n303 104.615
R291 VTAIL.n37 VTAIL.n31 104.615
R292 VTAIL.n38 VTAIL.n37 104.615
R293 VTAIL.n38 VTAIL.n27 104.615
R294 VTAIL.n45 VTAIL.n27 104.615
R295 VTAIL.n46 VTAIL.n45 104.615
R296 VTAIL.n46 VTAIL.n23 104.615
R297 VTAIL.n54 VTAIL.n23 104.615
R298 VTAIL.n55 VTAIL.n54 104.615
R299 VTAIL.n56 VTAIL.n55 104.615
R300 VTAIL.n56 VTAIL.n19 104.615
R301 VTAIL.n63 VTAIL.n19 104.615
R302 VTAIL.n64 VTAIL.n63 104.615
R303 VTAIL.n64 VTAIL.n15 104.615
R304 VTAIL.n71 VTAIL.n15 104.615
R305 VTAIL.n72 VTAIL.n71 104.615
R306 VTAIL.n72 VTAIL.n11 104.615
R307 VTAIL.n79 VTAIL.n11 104.615
R308 VTAIL.n80 VTAIL.n79 104.615
R309 VTAIL.n80 VTAIL.n7 104.615
R310 VTAIL.n87 VTAIL.n7 104.615
R311 VTAIL.n88 VTAIL.n87 104.615
R312 VTAIL.n88 VTAIL.n3 104.615
R313 VTAIL.n95 VTAIL.n3 104.615
R314 VTAIL.n299 VTAIL.n207 104.615
R315 VTAIL.n292 VTAIL.n207 104.615
R316 VTAIL.n292 VTAIL.n291 104.615
R317 VTAIL.n291 VTAIL.n211 104.615
R318 VTAIL.n284 VTAIL.n211 104.615
R319 VTAIL.n284 VTAIL.n283 104.615
R320 VTAIL.n283 VTAIL.n215 104.615
R321 VTAIL.n276 VTAIL.n215 104.615
R322 VTAIL.n276 VTAIL.n275 104.615
R323 VTAIL.n275 VTAIL.n219 104.615
R324 VTAIL.n268 VTAIL.n219 104.615
R325 VTAIL.n268 VTAIL.n267 104.615
R326 VTAIL.n267 VTAIL.n223 104.615
R327 VTAIL.n260 VTAIL.n223 104.615
R328 VTAIL.n260 VTAIL.n259 104.615
R329 VTAIL.n259 VTAIL.n258 104.615
R330 VTAIL.n258 VTAIL.n227 104.615
R331 VTAIL.n251 VTAIL.n227 104.615
R332 VTAIL.n251 VTAIL.n250 104.615
R333 VTAIL.n250 VTAIL.n232 104.615
R334 VTAIL.n243 VTAIL.n232 104.615
R335 VTAIL.n243 VTAIL.n242 104.615
R336 VTAIL.n242 VTAIL.n236 104.615
R337 VTAIL.n199 VTAIL.n107 104.615
R338 VTAIL.n192 VTAIL.n107 104.615
R339 VTAIL.n192 VTAIL.n191 104.615
R340 VTAIL.n191 VTAIL.n111 104.615
R341 VTAIL.n184 VTAIL.n111 104.615
R342 VTAIL.n184 VTAIL.n183 104.615
R343 VTAIL.n183 VTAIL.n115 104.615
R344 VTAIL.n176 VTAIL.n115 104.615
R345 VTAIL.n176 VTAIL.n175 104.615
R346 VTAIL.n175 VTAIL.n119 104.615
R347 VTAIL.n168 VTAIL.n119 104.615
R348 VTAIL.n168 VTAIL.n167 104.615
R349 VTAIL.n167 VTAIL.n123 104.615
R350 VTAIL.n160 VTAIL.n123 104.615
R351 VTAIL.n160 VTAIL.n159 104.615
R352 VTAIL.n159 VTAIL.n158 104.615
R353 VTAIL.n158 VTAIL.n127 104.615
R354 VTAIL.n151 VTAIL.n127 104.615
R355 VTAIL.n151 VTAIL.n150 104.615
R356 VTAIL.n150 VTAIL.n132 104.615
R357 VTAIL.n143 VTAIL.n132 104.615
R358 VTAIL.n143 VTAIL.n142 104.615
R359 VTAIL.n142 VTAIL.n136 104.615
R360 VTAIL.t5 VTAIL.n331 52.3082
R361 VTAIL.t10 VTAIL.n31 52.3082
R362 VTAIL.t15 VTAIL.n236 52.3082
R363 VTAIL.t3 VTAIL.n136 52.3082
R364 VTAIL.n205 VTAIL.n204 47.8278
R365 VTAIL.n203 VTAIL.n202 47.8278
R366 VTAIL.n105 VTAIL.n104 47.8278
R367 VTAIL.n103 VTAIL.n102 47.8278
R368 VTAIL.n399 VTAIL.n398 47.8268
R369 VTAIL.n1 VTAIL.n0 47.8268
R370 VTAIL.n99 VTAIL.n98 47.8268
R371 VTAIL.n101 VTAIL.n100 47.8268
R372 VTAIL.n397 VTAIL.n396 34.7066
R373 VTAIL.n97 VTAIL.n96 34.7066
R374 VTAIL.n301 VTAIL.n300 34.7066
R375 VTAIL.n201 VTAIL.n200 34.7066
R376 VTAIL.n103 VTAIL.n101 32.9962
R377 VTAIL.n397 VTAIL.n301 30.1772
R378 VTAIL.n357 VTAIL.n322 13.1884
R379 VTAIL.n57 VTAIL.n22 13.1884
R380 VTAIL.n261 VTAIL.n226 13.1884
R381 VTAIL.n161 VTAIL.n126 13.1884
R382 VTAIL.n353 VTAIL.n352 12.8005
R383 VTAIL.n358 VTAIL.n320 12.8005
R384 VTAIL.n53 VTAIL.n52 12.8005
R385 VTAIL.n58 VTAIL.n20 12.8005
R386 VTAIL.n262 VTAIL.n224 12.8005
R387 VTAIL.n257 VTAIL.n228 12.8005
R388 VTAIL.n162 VTAIL.n124 12.8005
R389 VTAIL.n157 VTAIL.n128 12.8005
R390 VTAIL.n351 VTAIL.n324 12.0247
R391 VTAIL.n362 VTAIL.n361 12.0247
R392 VTAIL.n51 VTAIL.n24 12.0247
R393 VTAIL.n62 VTAIL.n61 12.0247
R394 VTAIL.n266 VTAIL.n265 12.0247
R395 VTAIL.n256 VTAIL.n229 12.0247
R396 VTAIL.n166 VTAIL.n165 12.0247
R397 VTAIL.n156 VTAIL.n129 12.0247
R398 VTAIL.n348 VTAIL.n347 11.249
R399 VTAIL.n365 VTAIL.n318 11.249
R400 VTAIL.n394 VTAIL.n302 11.249
R401 VTAIL.n48 VTAIL.n47 11.249
R402 VTAIL.n65 VTAIL.n18 11.249
R403 VTAIL.n94 VTAIL.n2 11.249
R404 VTAIL.n298 VTAIL.n206 11.249
R405 VTAIL.n269 VTAIL.n222 11.249
R406 VTAIL.n253 VTAIL.n252 11.249
R407 VTAIL.n198 VTAIL.n106 11.249
R408 VTAIL.n169 VTAIL.n122 11.249
R409 VTAIL.n153 VTAIL.n152 11.249
R410 VTAIL.n344 VTAIL.n326 10.4732
R411 VTAIL.n366 VTAIL.n316 10.4732
R412 VTAIL.n393 VTAIL.n304 10.4732
R413 VTAIL.n44 VTAIL.n26 10.4732
R414 VTAIL.n66 VTAIL.n16 10.4732
R415 VTAIL.n93 VTAIL.n4 10.4732
R416 VTAIL.n297 VTAIL.n208 10.4732
R417 VTAIL.n270 VTAIL.n220 10.4732
R418 VTAIL.n249 VTAIL.n231 10.4732
R419 VTAIL.n197 VTAIL.n108 10.4732
R420 VTAIL.n170 VTAIL.n120 10.4732
R421 VTAIL.n149 VTAIL.n131 10.4732
R422 VTAIL.n333 VTAIL.n332 10.2747
R423 VTAIL.n33 VTAIL.n32 10.2747
R424 VTAIL.n238 VTAIL.n237 10.2747
R425 VTAIL.n138 VTAIL.n137 10.2747
R426 VTAIL.n343 VTAIL.n328 9.69747
R427 VTAIL.n370 VTAIL.n369 9.69747
R428 VTAIL.n390 VTAIL.n389 9.69747
R429 VTAIL.n43 VTAIL.n28 9.69747
R430 VTAIL.n70 VTAIL.n69 9.69747
R431 VTAIL.n90 VTAIL.n89 9.69747
R432 VTAIL.n294 VTAIL.n293 9.69747
R433 VTAIL.n274 VTAIL.n273 9.69747
R434 VTAIL.n248 VTAIL.n233 9.69747
R435 VTAIL.n194 VTAIL.n193 9.69747
R436 VTAIL.n174 VTAIL.n173 9.69747
R437 VTAIL.n148 VTAIL.n133 9.69747
R438 VTAIL.n392 VTAIL.n302 9.45567
R439 VTAIL.n92 VTAIL.n2 9.45567
R440 VTAIL.n296 VTAIL.n206 9.45567
R441 VTAIL.n196 VTAIL.n106 9.45567
R442 VTAIL.n310 VTAIL.n309 9.3005
R443 VTAIL.n383 VTAIL.n382 9.3005
R444 VTAIL.n385 VTAIL.n384 9.3005
R445 VTAIL.n306 VTAIL.n305 9.3005
R446 VTAIL.n391 VTAIL.n390 9.3005
R447 VTAIL.n393 VTAIL.n392 9.3005
R448 VTAIL.n375 VTAIL.n374 9.3005
R449 VTAIL.n314 VTAIL.n313 9.3005
R450 VTAIL.n369 VTAIL.n368 9.3005
R451 VTAIL.n367 VTAIL.n366 9.3005
R452 VTAIL.n318 VTAIL.n317 9.3005
R453 VTAIL.n361 VTAIL.n360 9.3005
R454 VTAIL.n359 VTAIL.n358 9.3005
R455 VTAIL.n335 VTAIL.n334 9.3005
R456 VTAIL.n330 VTAIL.n329 9.3005
R457 VTAIL.n341 VTAIL.n340 9.3005
R458 VTAIL.n343 VTAIL.n342 9.3005
R459 VTAIL.n326 VTAIL.n325 9.3005
R460 VTAIL.n349 VTAIL.n348 9.3005
R461 VTAIL.n351 VTAIL.n350 9.3005
R462 VTAIL.n352 VTAIL.n321 9.3005
R463 VTAIL.n377 VTAIL.n376 9.3005
R464 VTAIL.n10 VTAIL.n9 9.3005
R465 VTAIL.n83 VTAIL.n82 9.3005
R466 VTAIL.n85 VTAIL.n84 9.3005
R467 VTAIL.n6 VTAIL.n5 9.3005
R468 VTAIL.n91 VTAIL.n90 9.3005
R469 VTAIL.n93 VTAIL.n92 9.3005
R470 VTAIL.n75 VTAIL.n74 9.3005
R471 VTAIL.n14 VTAIL.n13 9.3005
R472 VTAIL.n69 VTAIL.n68 9.3005
R473 VTAIL.n67 VTAIL.n66 9.3005
R474 VTAIL.n18 VTAIL.n17 9.3005
R475 VTAIL.n61 VTAIL.n60 9.3005
R476 VTAIL.n59 VTAIL.n58 9.3005
R477 VTAIL.n35 VTAIL.n34 9.3005
R478 VTAIL.n30 VTAIL.n29 9.3005
R479 VTAIL.n41 VTAIL.n40 9.3005
R480 VTAIL.n43 VTAIL.n42 9.3005
R481 VTAIL.n26 VTAIL.n25 9.3005
R482 VTAIL.n49 VTAIL.n48 9.3005
R483 VTAIL.n51 VTAIL.n50 9.3005
R484 VTAIL.n52 VTAIL.n21 9.3005
R485 VTAIL.n77 VTAIL.n76 9.3005
R486 VTAIL.n297 VTAIL.n296 9.3005
R487 VTAIL.n295 VTAIL.n294 9.3005
R488 VTAIL.n210 VTAIL.n209 9.3005
R489 VTAIL.n289 VTAIL.n288 9.3005
R490 VTAIL.n287 VTAIL.n286 9.3005
R491 VTAIL.n214 VTAIL.n213 9.3005
R492 VTAIL.n281 VTAIL.n280 9.3005
R493 VTAIL.n279 VTAIL.n278 9.3005
R494 VTAIL.n218 VTAIL.n217 9.3005
R495 VTAIL.n273 VTAIL.n272 9.3005
R496 VTAIL.n271 VTAIL.n270 9.3005
R497 VTAIL.n222 VTAIL.n221 9.3005
R498 VTAIL.n265 VTAIL.n264 9.3005
R499 VTAIL.n263 VTAIL.n262 9.3005
R500 VTAIL.n228 VTAIL.n225 9.3005
R501 VTAIL.n256 VTAIL.n255 9.3005
R502 VTAIL.n254 VTAIL.n253 9.3005
R503 VTAIL.n231 VTAIL.n230 9.3005
R504 VTAIL.n248 VTAIL.n247 9.3005
R505 VTAIL.n246 VTAIL.n245 9.3005
R506 VTAIL.n235 VTAIL.n234 9.3005
R507 VTAIL.n240 VTAIL.n239 9.3005
R508 VTAIL.n140 VTAIL.n139 9.3005
R509 VTAIL.n135 VTAIL.n134 9.3005
R510 VTAIL.n146 VTAIL.n145 9.3005
R511 VTAIL.n148 VTAIL.n147 9.3005
R512 VTAIL.n131 VTAIL.n130 9.3005
R513 VTAIL.n154 VTAIL.n153 9.3005
R514 VTAIL.n156 VTAIL.n155 9.3005
R515 VTAIL.n128 VTAIL.n125 9.3005
R516 VTAIL.n187 VTAIL.n186 9.3005
R517 VTAIL.n189 VTAIL.n188 9.3005
R518 VTAIL.n110 VTAIL.n109 9.3005
R519 VTAIL.n195 VTAIL.n194 9.3005
R520 VTAIL.n197 VTAIL.n196 9.3005
R521 VTAIL.n114 VTAIL.n113 9.3005
R522 VTAIL.n181 VTAIL.n180 9.3005
R523 VTAIL.n179 VTAIL.n178 9.3005
R524 VTAIL.n118 VTAIL.n117 9.3005
R525 VTAIL.n173 VTAIL.n172 9.3005
R526 VTAIL.n171 VTAIL.n170 9.3005
R527 VTAIL.n122 VTAIL.n121 9.3005
R528 VTAIL.n165 VTAIL.n164 9.3005
R529 VTAIL.n163 VTAIL.n162 9.3005
R530 VTAIL.n340 VTAIL.n339 8.92171
R531 VTAIL.n373 VTAIL.n314 8.92171
R532 VTAIL.n386 VTAIL.n306 8.92171
R533 VTAIL.n40 VTAIL.n39 8.92171
R534 VTAIL.n73 VTAIL.n14 8.92171
R535 VTAIL.n86 VTAIL.n6 8.92171
R536 VTAIL.n290 VTAIL.n210 8.92171
R537 VTAIL.n277 VTAIL.n218 8.92171
R538 VTAIL.n245 VTAIL.n244 8.92171
R539 VTAIL.n190 VTAIL.n110 8.92171
R540 VTAIL.n177 VTAIL.n118 8.92171
R541 VTAIL.n145 VTAIL.n144 8.92171
R542 VTAIL.n336 VTAIL.n330 8.14595
R543 VTAIL.n374 VTAIL.n312 8.14595
R544 VTAIL.n385 VTAIL.n308 8.14595
R545 VTAIL.n36 VTAIL.n30 8.14595
R546 VTAIL.n74 VTAIL.n12 8.14595
R547 VTAIL.n85 VTAIL.n8 8.14595
R548 VTAIL.n289 VTAIL.n212 8.14595
R549 VTAIL.n278 VTAIL.n216 8.14595
R550 VTAIL.n241 VTAIL.n235 8.14595
R551 VTAIL.n189 VTAIL.n112 8.14595
R552 VTAIL.n178 VTAIL.n116 8.14595
R553 VTAIL.n141 VTAIL.n135 8.14595
R554 VTAIL.n335 VTAIL.n332 7.3702
R555 VTAIL.n378 VTAIL.n377 7.3702
R556 VTAIL.n382 VTAIL.n381 7.3702
R557 VTAIL.n35 VTAIL.n32 7.3702
R558 VTAIL.n78 VTAIL.n77 7.3702
R559 VTAIL.n82 VTAIL.n81 7.3702
R560 VTAIL.n286 VTAIL.n285 7.3702
R561 VTAIL.n282 VTAIL.n281 7.3702
R562 VTAIL.n240 VTAIL.n237 7.3702
R563 VTAIL.n186 VTAIL.n185 7.3702
R564 VTAIL.n182 VTAIL.n181 7.3702
R565 VTAIL.n140 VTAIL.n137 7.3702
R566 VTAIL.n378 VTAIL.n310 6.59444
R567 VTAIL.n381 VTAIL.n310 6.59444
R568 VTAIL.n78 VTAIL.n10 6.59444
R569 VTAIL.n81 VTAIL.n10 6.59444
R570 VTAIL.n285 VTAIL.n214 6.59444
R571 VTAIL.n282 VTAIL.n214 6.59444
R572 VTAIL.n185 VTAIL.n114 6.59444
R573 VTAIL.n182 VTAIL.n114 6.59444
R574 VTAIL.n336 VTAIL.n335 5.81868
R575 VTAIL.n377 VTAIL.n312 5.81868
R576 VTAIL.n382 VTAIL.n308 5.81868
R577 VTAIL.n36 VTAIL.n35 5.81868
R578 VTAIL.n77 VTAIL.n12 5.81868
R579 VTAIL.n82 VTAIL.n8 5.81868
R580 VTAIL.n286 VTAIL.n212 5.81868
R581 VTAIL.n281 VTAIL.n216 5.81868
R582 VTAIL.n241 VTAIL.n240 5.81868
R583 VTAIL.n186 VTAIL.n112 5.81868
R584 VTAIL.n181 VTAIL.n116 5.81868
R585 VTAIL.n141 VTAIL.n140 5.81868
R586 VTAIL.n339 VTAIL.n330 5.04292
R587 VTAIL.n374 VTAIL.n373 5.04292
R588 VTAIL.n386 VTAIL.n385 5.04292
R589 VTAIL.n39 VTAIL.n30 5.04292
R590 VTAIL.n74 VTAIL.n73 5.04292
R591 VTAIL.n86 VTAIL.n85 5.04292
R592 VTAIL.n290 VTAIL.n289 5.04292
R593 VTAIL.n278 VTAIL.n277 5.04292
R594 VTAIL.n244 VTAIL.n235 5.04292
R595 VTAIL.n190 VTAIL.n189 5.04292
R596 VTAIL.n178 VTAIL.n177 5.04292
R597 VTAIL.n144 VTAIL.n135 5.04292
R598 VTAIL.n340 VTAIL.n328 4.26717
R599 VTAIL.n370 VTAIL.n314 4.26717
R600 VTAIL.n389 VTAIL.n306 4.26717
R601 VTAIL.n40 VTAIL.n28 4.26717
R602 VTAIL.n70 VTAIL.n14 4.26717
R603 VTAIL.n89 VTAIL.n6 4.26717
R604 VTAIL.n293 VTAIL.n210 4.26717
R605 VTAIL.n274 VTAIL.n218 4.26717
R606 VTAIL.n245 VTAIL.n233 4.26717
R607 VTAIL.n193 VTAIL.n110 4.26717
R608 VTAIL.n174 VTAIL.n118 4.26717
R609 VTAIL.n145 VTAIL.n133 4.26717
R610 VTAIL.n344 VTAIL.n343 3.49141
R611 VTAIL.n369 VTAIL.n316 3.49141
R612 VTAIL.n390 VTAIL.n304 3.49141
R613 VTAIL.n44 VTAIL.n43 3.49141
R614 VTAIL.n69 VTAIL.n16 3.49141
R615 VTAIL.n90 VTAIL.n4 3.49141
R616 VTAIL.n294 VTAIL.n208 3.49141
R617 VTAIL.n273 VTAIL.n220 3.49141
R618 VTAIL.n249 VTAIL.n248 3.49141
R619 VTAIL.n194 VTAIL.n108 3.49141
R620 VTAIL.n173 VTAIL.n120 3.49141
R621 VTAIL.n149 VTAIL.n148 3.49141
R622 VTAIL.n334 VTAIL.n333 2.84303
R623 VTAIL.n34 VTAIL.n33 2.84303
R624 VTAIL.n239 VTAIL.n238 2.84303
R625 VTAIL.n139 VTAIL.n138 2.84303
R626 VTAIL.n105 VTAIL.n103 2.81947
R627 VTAIL.n201 VTAIL.n105 2.81947
R628 VTAIL.n205 VTAIL.n203 2.81947
R629 VTAIL.n301 VTAIL.n205 2.81947
R630 VTAIL.n101 VTAIL.n99 2.81947
R631 VTAIL.n99 VTAIL.n97 2.81947
R632 VTAIL.n399 VTAIL.n397 2.81947
R633 VTAIL.n347 VTAIL.n326 2.71565
R634 VTAIL.n366 VTAIL.n365 2.71565
R635 VTAIL.n394 VTAIL.n393 2.71565
R636 VTAIL.n47 VTAIL.n26 2.71565
R637 VTAIL.n66 VTAIL.n65 2.71565
R638 VTAIL.n94 VTAIL.n93 2.71565
R639 VTAIL.n298 VTAIL.n297 2.71565
R640 VTAIL.n270 VTAIL.n269 2.71565
R641 VTAIL.n252 VTAIL.n231 2.71565
R642 VTAIL.n198 VTAIL.n197 2.71565
R643 VTAIL.n170 VTAIL.n169 2.71565
R644 VTAIL.n152 VTAIL.n131 2.71565
R645 VTAIL VTAIL.n1 2.17291
R646 VTAIL.n348 VTAIL.n324 1.93989
R647 VTAIL.n362 VTAIL.n318 1.93989
R648 VTAIL.n396 VTAIL.n302 1.93989
R649 VTAIL.n48 VTAIL.n24 1.93989
R650 VTAIL.n62 VTAIL.n18 1.93989
R651 VTAIL.n96 VTAIL.n2 1.93989
R652 VTAIL.n300 VTAIL.n206 1.93989
R653 VTAIL.n266 VTAIL.n222 1.93989
R654 VTAIL.n253 VTAIL.n229 1.93989
R655 VTAIL.n200 VTAIL.n106 1.93989
R656 VTAIL.n166 VTAIL.n122 1.93989
R657 VTAIL.n153 VTAIL.n129 1.93989
R658 VTAIL.n203 VTAIL.n201 1.87981
R659 VTAIL.n97 VTAIL.n1 1.87981
R660 VTAIL.n353 VTAIL.n351 1.16414
R661 VTAIL.n361 VTAIL.n320 1.16414
R662 VTAIL.n53 VTAIL.n51 1.16414
R663 VTAIL.n61 VTAIL.n20 1.16414
R664 VTAIL.n265 VTAIL.n224 1.16414
R665 VTAIL.n257 VTAIL.n256 1.16414
R666 VTAIL.n165 VTAIL.n124 1.16414
R667 VTAIL.n157 VTAIL.n156 1.16414
R668 VTAIL.n398 VTAIL.t6 1.13909
R669 VTAIL.n398 VTAIL.t0 1.13909
R670 VTAIL.n0 VTAIL.t8 1.13909
R671 VTAIL.n0 VTAIL.t1 1.13909
R672 VTAIL.n98 VTAIL.t9 1.13909
R673 VTAIL.n98 VTAIL.t16 1.13909
R674 VTAIL.n100 VTAIL.t12 1.13909
R675 VTAIL.n100 VTAIL.t18 1.13909
R676 VTAIL.n204 VTAIL.t11 1.13909
R677 VTAIL.n204 VTAIL.t17 1.13909
R678 VTAIL.n202 VTAIL.t14 1.13909
R679 VTAIL.n202 VTAIL.t13 1.13909
R680 VTAIL.n104 VTAIL.t4 1.13909
R681 VTAIL.n104 VTAIL.t19 1.13909
R682 VTAIL.n102 VTAIL.t7 1.13909
R683 VTAIL.n102 VTAIL.t2 1.13909
R684 VTAIL VTAIL.n399 0.647052
R685 VTAIL.n352 VTAIL.n322 0.388379
R686 VTAIL.n358 VTAIL.n357 0.388379
R687 VTAIL.n52 VTAIL.n22 0.388379
R688 VTAIL.n58 VTAIL.n57 0.388379
R689 VTAIL.n262 VTAIL.n261 0.388379
R690 VTAIL.n228 VTAIL.n226 0.388379
R691 VTAIL.n162 VTAIL.n161 0.388379
R692 VTAIL.n128 VTAIL.n126 0.388379
R693 VTAIL.n334 VTAIL.n329 0.155672
R694 VTAIL.n341 VTAIL.n329 0.155672
R695 VTAIL.n342 VTAIL.n341 0.155672
R696 VTAIL.n342 VTAIL.n325 0.155672
R697 VTAIL.n349 VTAIL.n325 0.155672
R698 VTAIL.n350 VTAIL.n349 0.155672
R699 VTAIL.n350 VTAIL.n321 0.155672
R700 VTAIL.n359 VTAIL.n321 0.155672
R701 VTAIL.n360 VTAIL.n359 0.155672
R702 VTAIL.n360 VTAIL.n317 0.155672
R703 VTAIL.n367 VTAIL.n317 0.155672
R704 VTAIL.n368 VTAIL.n367 0.155672
R705 VTAIL.n368 VTAIL.n313 0.155672
R706 VTAIL.n375 VTAIL.n313 0.155672
R707 VTAIL.n376 VTAIL.n375 0.155672
R708 VTAIL.n376 VTAIL.n309 0.155672
R709 VTAIL.n383 VTAIL.n309 0.155672
R710 VTAIL.n384 VTAIL.n383 0.155672
R711 VTAIL.n384 VTAIL.n305 0.155672
R712 VTAIL.n391 VTAIL.n305 0.155672
R713 VTAIL.n392 VTAIL.n391 0.155672
R714 VTAIL.n34 VTAIL.n29 0.155672
R715 VTAIL.n41 VTAIL.n29 0.155672
R716 VTAIL.n42 VTAIL.n41 0.155672
R717 VTAIL.n42 VTAIL.n25 0.155672
R718 VTAIL.n49 VTAIL.n25 0.155672
R719 VTAIL.n50 VTAIL.n49 0.155672
R720 VTAIL.n50 VTAIL.n21 0.155672
R721 VTAIL.n59 VTAIL.n21 0.155672
R722 VTAIL.n60 VTAIL.n59 0.155672
R723 VTAIL.n60 VTAIL.n17 0.155672
R724 VTAIL.n67 VTAIL.n17 0.155672
R725 VTAIL.n68 VTAIL.n67 0.155672
R726 VTAIL.n68 VTAIL.n13 0.155672
R727 VTAIL.n75 VTAIL.n13 0.155672
R728 VTAIL.n76 VTAIL.n75 0.155672
R729 VTAIL.n76 VTAIL.n9 0.155672
R730 VTAIL.n83 VTAIL.n9 0.155672
R731 VTAIL.n84 VTAIL.n83 0.155672
R732 VTAIL.n84 VTAIL.n5 0.155672
R733 VTAIL.n91 VTAIL.n5 0.155672
R734 VTAIL.n92 VTAIL.n91 0.155672
R735 VTAIL.n296 VTAIL.n295 0.155672
R736 VTAIL.n295 VTAIL.n209 0.155672
R737 VTAIL.n288 VTAIL.n209 0.155672
R738 VTAIL.n288 VTAIL.n287 0.155672
R739 VTAIL.n287 VTAIL.n213 0.155672
R740 VTAIL.n280 VTAIL.n213 0.155672
R741 VTAIL.n280 VTAIL.n279 0.155672
R742 VTAIL.n279 VTAIL.n217 0.155672
R743 VTAIL.n272 VTAIL.n217 0.155672
R744 VTAIL.n272 VTAIL.n271 0.155672
R745 VTAIL.n271 VTAIL.n221 0.155672
R746 VTAIL.n264 VTAIL.n221 0.155672
R747 VTAIL.n264 VTAIL.n263 0.155672
R748 VTAIL.n263 VTAIL.n225 0.155672
R749 VTAIL.n255 VTAIL.n225 0.155672
R750 VTAIL.n255 VTAIL.n254 0.155672
R751 VTAIL.n254 VTAIL.n230 0.155672
R752 VTAIL.n247 VTAIL.n230 0.155672
R753 VTAIL.n247 VTAIL.n246 0.155672
R754 VTAIL.n246 VTAIL.n234 0.155672
R755 VTAIL.n239 VTAIL.n234 0.155672
R756 VTAIL.n196 VTAIL.n195 0.155672
R757 VTAIL.n195 VTAIL.n109 0.155672
R758 VTAIL.n188 VTAIL.n109 0.155672
R759 VTAIL.n188 VTAIL.n187 0.155672
R760 VTAIL.n187 VTAIL.n113 0.155672
R761 VTAIL.n180 VTAIL.n113 0.155672
R762 VTAIL.n180 VTAIL.n179 0.155672
R763 VTAIL.n179 VTAIL.n117 0.155672
R764 VTAIL.n172 VTAIL.n117 0.155672
R765 VTAIL.n172 VTAIL.n171 0.155672
R766 VTAIL.n171 VTAIL.n121 0.155672
R767 VTAIL.n164 VTAIL.n121 0.155672
R768 VTAIL.n164 VTAIL.n163 0.155672
R769 VTAIL.n163 VTAIL.n125 0.155672
R770 VTAIL.n155 VTAIL.n125 0.155672
R771 VTAIL.n155 VTAIL.n154 0.155672
R772 VTAIL.n154 VTAIL.n130 0.155672
R773 VTAIL.n147 VTAIL.n130 0.155672
R774 VTAIL.n147 VTAIL.n146 0.155672
R775 VTAIL.n146 VTAIL.n134 0.155672
R776 VTAIL.n139 VTAIL.n134 0.155672
R777 VDD1.n94 VDD1.n93 289.615
R778 VDD1.n191 VDD1.n190 289.615
R779 VDD1.n93 VDD1.n92 185
R780 VDD1.n2 VDD1.n1 185
R781 VDD1.n87 VDD1.n86 185
R782 VDD1.n85 VDD1.n84 185
R783 VDD1.n6 VDD1.n5 185
R784 VDD1.n79 VDD1.n78 185
R785 VDD1.n77 VDD1.n76 185
R786 VDD1.n10 VDD1.n9 185
R787 VDD1.n71 VDD1.n70 185
R788 VDD1.n69 VDD1.n68 185
R789 VDD1.n14 VDD1.n13 185
R790 VDD1.n63 VDD1.n62 185
R791 VDD1.n61 VDD1.n60 185
R792 VDD1.n18 VDD1.n17 185
R793 VDD1.n55 VDD1.n54 185
R794 VDD1.n53 VDD1.n20 185
R795 VDD1.n52 VDD1.n51 185
R796 VDD1.n23 VDD1.n21 185
R797 VDD1.n46 VDD1.n45 185
R798 VDD1.n44 VDD1.n43 185
R799 VDD1.n27 VDD1.n26 185
R800 VDD1.n38 VDD1.n37 185
R801 VDD1.n36 VDD1.n35 185
R802 VDD1.n31 VDD1.n30 185
R803 VDD1.n127 VDD1.n126 185
R804 VDD1.n132 VDD1.n131 185
R805 VDD1.n134 VDD1.n133 185
R806 VDD1.n123 VDD1.n122 185
R807 VDD1.n140 VDD1.n139 185
R808 VDD1.n142 VDD1.n141 185
R809 VDD1.n119 VDD1.n118 185
R810 VDD1.n149 VDD1.n148 185
R811 VDD1.n150 VDD1.n117 185
R812 VDD1.n152 VDD1.n151 185
R813 VDD1.n115 VDD1.n114 185
R814 VDD1.n158 VDD1.n157 185
R815 VDD1.n160 VDD1.n159 185
R816 VDD1.n111 VDD1.n110 185
R817 VDD1.n166 VDD1.n165 185
R818 VDD1.n168 VDD1.n167 185
R819 VDD1.n107 VDD1.n106 185
R820 VDD1.n174 VDD1.n173 185
R821 VDD1.n176 VDD1.n175 185
R822 VDD1.n103 VDD1.n102 185
R823 VDD1.n182 VDD1.n181 185
R824 VDD1.n184 VDD1.n183 185
R825 VDD1.n99 VDD1.n98 185
R826 VDD1.n190 VDD1.n189 185
R827 VDD1.n32 VDD1.t3 149.524
R828 VDD1.n128 VDD1.t1 149.524
R829 VDD1.n93 VDD1.n1 104.615
R830 VDD1.n86 VDD1.n1 104.615
R831 VDD1.n86 VDD1.n85 104.615
R832 VDD1.n85 VDD1.n5 104.615
R833 VDD1.n78 VDD1.n5 104.615
R834 VDD1.n78 VDD1.n77 104.615
R835 VDD1.n77 VDD1.n9 104.615
R836 VDD1.n70 VDD1.n9 104.615
R837 VDD1.n70 VDD1.n69 104.615
R838 VDD1.n69 VDD1.n13 104.615
R839 VDD1.n62 VDD1.n13 104.615
R840 VDD1.n62 VDD1.n61 104.615
R841 VDD1.n61 VDD1.n17 104.615
R842 VDD1.n54 VDD1.n17 104.615
R843 VDD1.n54 VDD1.n53 104.615
R844 VDD1.n53 VDD1.n52 104.615
R845 VDD1.n52 VDD1.n21 104.615
R846 VDD1.n45 VDD1.n21 104.615
R847 VDD1.n45 VDD1.n44 104.615
R848 VDD1.n44 VDD1.n26 104.615
R849 VDD1.n37 VDD1.n26 104.615
R850 VDD1.n37 VDD1.n36 104.615
R851 VDD1.n36 VDD1.n30 104.615
R852 VDD1.n132 VDD1.n126 104.615
R853 VDD1.n133 VDD1.n132 104.615
R854 VDD1.n133 VDD1.n122 104.615
R855 VDD1.n140 VDD1.n122 104.615
R856 VDD1.n141 VDD1.n140 104.615
R857 VDD1.n141 VDD1.n118 104.615
R858 VDD1.n149 VDD1.n118 104.615
R859 VDD1.n150 VDD1.n149 104.615
R860 VDD1.n151 VDD1.n150 104.615
R861 VDD1.n151 VDD1.n114 104.615
R862 VDD1.n158 VDD1.n114 104.615
R863 VDD1.n159 VDD1.n158 104.615
R864 VDD1.n159 VDD1.n110 104.615
R865 VDD1.n166 VDD1.n110 104.615
R866 VDD1.n167 VDD1.n166 104.615
R867 VDD1.n167 VDD1.n106 104.615
R868 VDD1.n174 VDD1.n106 104.615
R869 VDD1.n175 VDD1.n174 104.615
R870 VDD1.n175 VDD1.n102 104.615
R871 VDD1.n182 VDD1.n102 104.615
R872 VDD1.n183 VDD1.n182 104.615
R873 VDD1.n183 VDD1.n98 104.615
R874 VDD1.n190 VDD1.n98 104.615
R875 VDD1.n195 VDD1.n194 66.5645
R876 VDD1.n96 VDD1.n95 64.5066
R877 VDD1.n193 VDD1.n192 64.5056
R878 VDD1.n197 VDD1.n196 64.5054
R879 VDD1.n96 VDD1.n94 54.2043
R880 VDD1.n193 VDD1.n191 54.2043
R881 VDD1.n197 VDD1.n195 54.0893
R882 VDD1.t3 VDD1.n30 52.3082
R883 VDD1.t1 VDD1.n126 52.3082
R884 VDD1.n55 VDD1.n20 13.1884
R885 VDD1.n152 VDD1.n117 13.1884
R886 VDD1.n56 VDD1.n18 12.8005
R887 VDD1.n51 VDD1.n22 12.8005
R888 VDD1.n148 VDD1.n147 12.8005
R889 VDD1.n153 VDD1.n115 12.8005
R890 VDD1.n60 VDD1.n59 12.0247
R891 VDD1.n50 VDD1.n23 12.0247
R892 VDD1.n146 VDD1.n119 12.0247
R893 VDD1.n157 VDD1.n156 12.0247
R894 VDD1.n92 VDD1.n0 11.249
R895 VDD1.n63 VDD1.n16 11.249
R896 VDD1.n47 VDD1.n46 11.249
R897 VDD1.n143 VDD1.n142 11.249
R898 VDD1.n160 VDD1.n113 11.249
R899 VDD1.n189 VDD1.n97 11.249
R900 VDD1.n91 VDD1.n2 10.4732
R901 VDD1.n64 VDD1.n14 10.4732
R902 VDD1.n43 VDD1.n25 10.4732
R903 VDD1.n139 VDD1.n121 10.4732
R904 VDD1.n161 VDD1.n111 10.4732
R905 VDD1.n188 VDD1.n99 10.4732
R906 VDD1.n32 VDD1.n31 10.2747
R907 VDD1.n128 VDD1.n127 10.2747
R908 VDD1.n88 VDD1.n87 9.69747
R909 VDD1.n68 VDD1.n67 9.69747
R910 VDD1.n42 VDD1.n27 9.69747
R911 VDD1.n138 VDD1.n123 9.69747
R912 VDD1.n165 VDD1.n164 9.69747
R913 VDD1.n185 VDD1.n184 9.69747
R914 VDD1.n90 VDD1.n0 9.45567
R915 VDD1.n187 VDD1.n97 9.45567
R916 VDD1.n34 VDD1.n33 9.3005
R917 VDD1.n29 VDD1.n28 9.3005
R918 VDD1.n40 VDD1.n39 9.3005
R919 VDD1.n42 VDD1.n41 9.3005
R920 VDD1.n25 VDD1.n24 9.3005
R921 VDD1.n48 VDD1.n47 9.3005
R922 VDD1.n50 VDD1.n49 9.3005
R923 VDD1.n22 VDD1.n19 9.3005
R924 VDD1.n81 VDD1.n80 9.3005
R925 VDD1.n83 VDD1.n82 9.3005
R926 VDD1.n4 VDD1.n3 9.3005
R927 VDD1.n89 VDD1.n88 9.3005
R928 VDD1.n91 VDD1.n90 9.3005
R929 VDD1.n8 VDD1.n7 9.3005
R930 VDD1.n75 VDD1.n74 9.3005
R931 VDD1.n73 VDD1.n72 9.3005
R932 VDD1.n12 VDD1.n11 9.3005
R933 VDD1.n67 VDD1.n66 9.3005
R934 VDD1.n65 VDD1.n64 9.3005
R935 VDD1.n16 VDD1.n15 9.3005
R936 VDD1.n59 VDD1.n58 9.3005
R937 VDD1.n57 VDD1.n56 9.3005
R938 VDD1.n105 VDD1.n104 9.3005
R939 VDD1.n178 VDD1.n177 9.3005
R940 VDD1.n180 VDD1.n179 9.3005
R941 VDD1.n101 VDD1.n100 9.3005
R942 VDD1.n186 VDD1.n185 9.3005
R943 VDD1.n188 VDD1.n187 9.3005
R944 VDD1.n170 VDD1.n169 9.3005
R945 VDD1.n109 VDD1.n108 9.3005
R946 VDD1.n164 VDD1.n163 9.3005
R947 VDD1.n162 VDD1.n161 9.3005
R948 VDD1.n113 VDD1.n112 9.3005
R949 VDD1.n156 VDD1.n155 9.3005
R950 VDD1.n154 VDD1.n153 9.3005
R951 VDD1.n130 VDD1.n129 9.3005
R952 VDD1.n125 VDD1.n124 9.3005
R953 VDD1.n136 VDD1.n135 9.3005
R954 VDD1.n138 VDD1.n137 9.3005
R955 VDD1.n121 VDD1.n120 9.3005
R956 VDD1.n144 VDD1.n143 9.3005
R957 VDD1.n146 VDD1.n145 9.3005
R958 VDD1.n147 VDD1.n116 9.3005
R959 VDD1.n172 VDD1.n171 9.3005
R960 VDD1.n84 VDD1.n4 8.92171
R961 VDD1.n71 VDD1.n12 8.92171
R962 VDD1.n39 VDD1.n38 8.92171
R963 VDD1.n135 VDD1.n134 8.92171
R964 VDD1.n168 VDD1.n109 8.92171
R965 VDD1.n181 VDD1.n101 8.92171
R966 VDD1.n83 VDD1.n6 8.14595
R967 VDD1.n72 VDD1.n10 8.14595
R968 VDD1.n35 VDD1.n29 8.14595
R969 VDD1.n131 VDD1.n125 8.14595
R970 VDD1.n169 VDD1.n107 8.14595
R971 VDD1.n180 VDD1.n103 8.14595
R972 VDD1.n80 VDD1.n79 7.3702
R973 VDD1.n76 VDD1.n75 7.3702
R974 VDD1.n34 VDD1.n31 7.3702
R975 VDD1.n130 VDD1.n127 7.3702
R976 VDD1.n173 VDD1.n172 7.3702
R977 VDD1.n177 VDD1.n176 7.3702
R978 VDD1.n79 VDD1.n8 6.59444
R979 VDD1.n76 VDD1.n8 6.59444
R980 VDD1.n173 VDD1.n105 6.59444
R981 VDD1.n176 VDD1.n105 6.59444
R982 VDD1.n80 VDD1.n6 5.81868
R983 VDD1.n75 VDD1.n10 5.81868
R984 VDD1.n35 VDD1.n34 5.81868
R985 VDD1.n131 VDD1.n130 5.81868
R986 VDD1.n172 VDD1.n107 5.81868
R987 VDD1.n177 VDD1.n103 5.81868
R988 VDD1.n84 VDD1.n83 5.04292
R989 VDD1.n72 VDD1.n71 5.04292
R990 VDD1.n38 VDD1.n29 5.04292
R991 VDD1.n134 VDD1.n125 5.04292
R992 VDD1.n169 VDD1.n168 5.04292
R993 VDD1.n181 VDD1.n180 5.04292
R994 VDD1.n87 VDD1.n4 4.26717
R995 VDD1.n68 VDD1.n12 4.26717
R996 VDD1.n39 VDD1.n27 4.26717
R997 VDD1.n135 VDD1.n123 4.26717
R998 VDD1.n165 VDD1.n109 4.26717
R999 VDD1.n184 VDD1.n101 4.26717
R1000 VDD1.n88 VDD1.n2 3.49141
R1001 VDD1.n67 VDD1.n14 3.49141
R1002 VDD1.n43 VDD1.n42 3.49141
R1003 VDD1.n139 VDD1.n138 3.49141
R1004 VDD1.n164 VDD1.n111 3.49141
R1005 VDD1.n185 VDD1.n99 3.49141
R1006 VDD1.n129 VDD1.n128 2.84303
R1007 VDD1.n33 VDD1.n32 2.84303
R1008 VDD1.n92 VDD1.n91 2.71565
R1009 VDD1.n64 VDD1.n63 2.71565
R1010 VDD1.n46 VDD1.n25 2.71565
R1011 VDD1.n142 VDD1.n121 2.71565
R1012 VDD1.n161 VDD1.n160 2.71565
R1013 VDD1.n189 VDD1.n188 2.71565
R1014 VDD1 VDD1.n197 2.05653
R1015 VDD1.n94 VDD1.n0 1.93989
R1016 VDD1.n60 VDD1.n16 1.93989
R1017 VDD1.n47 VDD1.n23 1.93989
R1018 VDD1.n143 VDD1.n119 1.93989
R1019 VDD1.n157 VDD1.n113 1.93989
R1020 VDD1.n191 VDD1.n97 1.93989
R1021 VDD1.n59 VDD1.n18 1.16414
R1022 VDD1.n51 VDD1.n50 1.16414
R1023 VDD1.n148 VDD1.n146 1.16414
R1024 VDD1.n156 VDD1.n115 1.16414
R1025 VDD1.n196 VDD1.t7 1.13909
R1026 VDD1.n196 VDD1.t9 1.13909
R1027 VDD1.n95 VDD1.t8 1.13909
R1028 VDD1.n95 VDD1.t0 1.13909
R1029 VDD1.n194 VDD1.t4 1.13909
R1030 VDD1.n194 VDD1.t6 1.13909
R1031 VDD1.n192 VDD1.t2 1.13909
R1032 VDD1.n192 VDD1.t5 1.13909
R1033 VDD1 VDD1.n96 0.763431
R1034 VDD1.n195 VDD1.n193 0.649895
R1035 VDD1.n56 VDD1.n55 0.388379
R1036 VDD1.n22 VDD1.n20 0.388379
R1037 VDD1.n147 VDD1.n117 0.388379
R1038 VDD1.n153 VDD1.n152 0.388379
R1039 VDD1.n90 VDD1.n89 0.155672
R1040 VDD1.n89 VDD1.n3 0.155672
R1041 VDD1.n82 VDD1.n3 0.155672
R1042 VDD1.n82 VDD1.n81 0.155672
R1043 VDD1.n81 VDD1.n7 0.155672
R1044 VDD1.n74 VDD1.n7 0.155672
R1045 VDD1.n74 VDD1.n73 0.155672
R1046 VDD1.n73 VDD1.n11 0.155672
R1047 VDD1.n66 VDD1.n11 0.155672
R1048 VDD1.n66 VDD1.n65 0.155672
R1049 VDD1.n65 VDD1.n15 0.155672
R1050 VDD1.n58 VDD1.n15 0.155672
R1051 VDD1.n58 VDD1.n57 0.155672
R1052 VDD1.n57 VDD1.n19 0.155672
R1053 VDD1.n49 VDD1.n19 0.155672
R1054 VDD1.n49 VDD1.n48 0.155672
R1055 VDD1.n48 VDD1.n24 0.155672
R1056 VDD1.n41 VDD1.n24 0.155672
R1057 VDD1.n41 VDD1.n40 0.155672
R1058 VDD1.n40 VDD1.n28 0.155672
R1059 VDD1.n33 VDD1.n28 0.155672
R1060 VDD1.n129 VDD1.n124 0.155672
R1061 VDD1.n136 VDD1.n124 0.155672
R1062 VDD1.n137 VDD1.n136 0.155672
R1063 VDD1.n137 VDD1.n120 0.155672
R1064 VDD1.n144 VDD1.n120 0.155672
R1065 VDD1.n145 VDD1.n144 0.155672
R1066 VDD1.n145 VDD1.n116 0.155672
R1067 VDD1.n154 VDD1.n116 0.155672
R1068 VDD1.n155 VDD1.n154 0.155672
R1069 VDD1.n155 VDD1.n112 0.155672
R1070 VDD1.n162 VDD1.n112 0.155672
R1071 VDD1.n163 VDD1.n162 0.155672
R1072 VDD1.n163 VDD1.n108 0.155672
R1073 VDD1.n170 VDD1.n108 0.155672
R1074 VDD1.n171 VDD1.n170 0.155672
R1075 VDD1.n171 VDD1.n104 0.155672
R1076 VDD1.n178 VDD1.n104 0.155672
R1077 VDD1.n179 VDD1.n178 0.155672
R1078 VDD1.n179 VDD1.n100 0.155672
R1079 VDD1.n186 VDD1.n100 0.155672
R1080 VDD1.n187 VDD1.n186 0.155672
R1081 B.n918 B.n917 585
R1082 B.n918 B.n120 585
R1083 B.n921 B.n920 585
R1084 B.n922 B.n187 585
R1085 B.n924 B.n923 585
R1086 B.n926 B.n186 585
R1087 B.n929 B.n928 585
R1088 B.n930 B.n185 585
R1089 B.n932 B.n931 585
R1090 B.n934 B.n184 585
R1091 B.n937 B.n936 585
R1092 B.n938 B.n183 585
R1093 B.n940 B.n939 585
R1094 B.n942 B.n182 585
R1095 B.n945 B.n944 585
R1096 B.n946 B.n181 585
R1097 B.n948 B.n947 585
R1098 B.n950 B.n180 585
R1099 B.n953 B.n952 585
R1100 B.n954 B.n179 585
R1101 B.n956 B.n955 585
R1102 B.n958 B.n178 585
R1103 B.n961 B.n960 585
R1104 B.n962 B.n177 585
R1105 B.n964 B.n963 585
R1106 B.n966 B.n176 585
R1107 B.n969 B.n968 585
R1108 B.n970 B.n175 585
R1109 B.n972 B.n971 585
R1110 B.n974 B.n174 585
R1111 B.n977 B.n976 585
R1112 B.n978 B.n173 585
R1113 B.n980 B.n979 585
R1114 B.n982 B.n172 585
R1115 B.n985 B.n984 585
R1116 B.n986 B.n171 585
R1117 B.n988 B.n987 585
R1118 B.n990 B.n170 585
R1119 B.n993 B.n992 585
R1120 B.n994 B.n169 585
R1121 B.n996 B.n995 585
R1122 B.n998 B.n168 585
R1123 B.n1001 B.n1000 585
R1124 B.n1002 B.n167 585
R1125 B.n1004 B.n1003 585
R1126 B.n1006 B.n166 585
R1127 B.n1009 B.n1008 585
R1128 B.n1010 B.n165 585
R1129 B.n1012 B.n1011 585
R1130 B.n1014 B.n164 585
R1131 B.n1017 B.n1016 585
R1132 B.n1018 B.n163 585
R1133 B.n1020 B.n1019 585
R1134 B.n1022 B.n162 585
R1135 B.n1025 B.n1024 585
R1136 B.n1026 B.n161 585
R1137 B.n1028 B.n1027 585
R1138 B.n1030 B.n160 585
R1139 B.n1033 B.n1032 585
R1140 B.n1035 B.n157 585
R1141 B.n1037 B.n1036 585
R1142 B.n1039 B.n156 585
R1143 B.n1042 B.n1041 585
R1144 B.n1043 B.n155 585
R1145 B.n1045 B.n1044 585
R1146 B.n1047 B.n154 585
R1147 B.n1049 B.n1048 585
R1148 B.n1051 B.n1050 585
R1149 B.n1054 B.n1053 585
R1150 B.n1055 B.n149 585
R1151 B.n1057 B.n1056 585
R1152 B.n1059 B.n148 585
R1153 B.n1062 B.n1061 585
R1154 B.n1063 B.n147 585
R1155 B.n1065 B.n1064 585
R1156 B.n1067 B.n146 585
R1157 B.n1070 B.n1069 585
R1158 B.n1071 B.n145 585
R1159 B.n1073 B.n1072 585
R1160 B.n1075 B.n144 585
R1161 B.n1078 B.n1077 585
R1162 B.n1079 B.n143 585
R1163 B.n1081 B.n1080 585
R1164 B.n1083 B.n142 585
R1165 B.n1086 B.n1085 585
R1166 B.n1087 B.n141 585
R1167 B.n1089 B.n1088 585
R1168 B.n1091 B.n140 585
R1169 B.n1094 B.n1093 585
R1170 B.n1095 B.n139 585
R1171 B.n1097 B.n1096 585
R1172 B.n1099 B.n138 585
R1173 B.n1102 B.n1101 585
R1174 B.n1103 B.n137 585
R1175 B.n1105 B.n1104 585
R1176 B.n1107 B.n136 585
R1177 B.n1110 B.n1109 585
R1178 B.n1111 B.n135 585
R1179 B.n1113 B.n1112 585
R1180 B.n1115 B.n134 585
R1181 B.n1118 B.n1117 585
R1182 B.n1119 B.n133 585
R1183 B.n1121 B.n1120 585
R1184 B.n1123 B.n132 585
R1185 B.n1126 B.n1125 585
R1186 B.n1127 B.n131 585
R1187 B.n1129 B.n1128 585
R1188 B.n1131 B.n130 585
R1189 B.n1134 B.n1133 585
R1190 B.n1135 B.n129 585
R1191 B.n1137 B.n1136 585
R1192 B.n1139 B.n128 585
R1193 B.n1142 B.n1141 585
R1194 B.n1143 B.n127 585
R1195 B.n1145 B.n1144 585
R1196 B.n1147 B.n126 585
R1197 B.n1150 B.n1149 585
R1198 B.n1151 B.n125 585
R1199 B.n1153 B.n1152 585
R1200 B.n1155 B.n124 585
R1201 B.n1158 B.n1157 585
R1202 B.n1159 B.n123 585
R1203 B.n1161 B.n1160 585
R1204 B.n1163 B.n122 585
R1205 B.n1166 B.n1165 585
R1206 B.n1167 B.n121 585
R1207 B.n916 B.n119 585
R1208 B.n1170 B.n119 585
R1209 B.n915 B.n118 585
R1210 B.n1171 B.n118 585
R1211 B.n914 B.n117 585
R1212 B.n1172 B.n117 585
R1213 B.n913 B.n912 585
R1214 B.n912 B.n113 585
R1215 B.n911 B.n112 585
R1216 B.n1178 B.n112 585
R1217 B.n910 B.n111 585
R1218 B.n1179 B.n111 585
R1219 B.n909 B.n110 585
R1220 B.n1180 B.n110 585
R1221 B.n908 B.n907 585
R1222 B.n907 B.n106 585
R1223 B.n906 B.n105 585
R1224 B.n1186 B.n105 585
R1225 B.n905 B.n104 585
R1226 B.n1187 B.n104 585
R1227 B.n904 B.n103 585
R1228 B.n1188 B.n103 585
R1229 B.n903 B.n902 585
R1230 B.n902 B.n99 585
R1231 B.n901 B.n98 585
R1232 B.n1194 B.n98 585
R1233 B.n900 B.n97 585
R1234 B.n1195 B.n97 585
R1235 B.n899 B.n96 585
R1236 B.n1196 B.n96 585
R1237 B.n898 B.n897 585
R1238 B.n897 B.n92 585
R1239 B.n896 B.n91 585
R1240 B.n1202 B.n91 585
R1241 B.n895 B.n90 585
R1242 B.n1203 B.n90 585
R1243 B.n894 B.n89 585
R1244 B.n1204 B.n89 585
R1245 B.n893 B.n892 585
R1246 B.n892 B.n85 585
R1247 B.n891 B.n84 585
R1248 B.n1210 B.n84 585
R1249 B.n890 B.n83 585
R1250 B.n1211 B.n83 585
R1251 B.n889 B.n82 585
R1252 B.n1212 B.n82 585
R1253 B.n888 B.n887 585
R1254 B.n887 B.n78 585
R1255 B.n886 B.n77 585
R1256 B.n1218 B.n77 585
R1257 B.n885 B.n76 585
R1258 B.n1219 B.n76 585
R1259 B.n884 B.n75 585
R1260 B.n1220 B.n75 585
R1261 B.n883 B.n882 585
R1262 B.n882 B.n71 585
R1263 B.n881 B.n70 585
R1264 B.n1226 B.n70 585
R1265 B.n880 B.n69 585
R1266 B.n1227 B.n69 585
R1267 B.n879 B.n68 585
R1268 B.n1228 B.n68 585
R1269 B.n878 B.n877 585
R1270 B.n877 B.n64 585
R1271 B.n876 B.n63 585
R1272 B.n1234 B.n63 585
R1273 B.n875 B.n62 585
R1274 B.n1235 B.n62 585
R1275 B.n874 B.n61 585
R1276 B.n1236 B.n61 585
R1277 B.n873 B.n872 585
R1278 B.n872 B.n57 585
R1279 B.n871 B.n56 585
R1280 B.n1242 B.n56 585
R1281 B.n870 B.n55 585
R1282 B.n1243 B.n55 585
R1283 B.n869 B.n54 585
R1284 B.n1244 B.n54 585
R1285 B.n868 B.n867 585
R1286 B.n867 B.n50 585
R1287 B.n866 B.n49 585
R1288 B.n1250 B.n49 585
R1289 B.n865 B.n48 585
R1290 B.n1251 B.n48 585
R1291 B.n864 B.n47 585
R1292 B.n1252 B.n47 585
R1293 B.n863 B.n862 585
R1294 B.n862 B.n43 585
R1295 B.n861 B.n42 585
R1296 B.n1258 B.n42 585
R1297 B.n860 B.n41 585
R1298 B.n1259 B.n41 585
R1299 B.n859 B.n40 585
R1300 B.n1260 B.n40 585
R1301 B.n858 B.n857 585
R1302 B.n857 B.n36 585
R1303 B.n856 B.n35 585
R1304 B.n1266 B.n35 585
R1305 B.n855 B.n34 585
R1306 B.n1267 B.n34 585
R1307 B.n854 B.n33 585
R1308 B.n1268 B.n33 585
R1309 B.n853 B.n852 585
R1310 B.n852 B.n29 585
R1311 B.n851 B.n28 585
R1312 B.n1274 B.n28 585
R1313 B.n850 B.n27 585
R1314 B.n1275 B.n27 585
R1315 B.n849 B.n26 585
R1316 B.n1276 B.n26 585
R1317 B.n848 B.n847 585
R1318 B.n847 B.n22 585
R1319 B.n846 B.n21 585
R1320 B.n1282 B.n21 585
R1321 B.n845 B.n20 585
R1322 B.n1283 B.n20 585
R1323 B.n844 B.n19 585
R1324 B.n1284 B.n19 585
R1325 B.n843 B.n842 585
R1326 B.n842 B.n18 585
R1327 B.n841 B.n14 585
R1328 B.n1290 B.n14 585
R1329 B.n840 B.n13 585
R1330 B.n1291 B.n13 585
R1331 B.n839 B.n12 585
R1332 B.n1292 B.n12 585
R1333 B.n838 B.n837 585
R1334 B.n837 B.n8 585
R1335 B.n836 B.n7 585
R1336 B.n1298 B.n7 585
R1337 B.n835 B.n6 585
R1338 B.n1299 B.n6 585
R1339 B.n834 B.n5 585
R1340 B.n1300 B.n5 585
R1341 B.n833 B.n832 585
R1342 B.n832 B.n4 585
R1343 B.n831 B.n188 585
R1344 B.n831 B.n830 585
R1345 B.n821 B.n189 585
R1346 B.n190 B.n189 585
R1347 B.n823 B.n822 585
R1348 B.n824 B.n823 585
R1349 B.n820 B.n195 585
R1350 B.n195 B.n194 585
R1351 B.n819 B.n818 585
R1352 B.n818 B.n817 585
R1353 B.n197 B.n196 585
R1354 B.n810 B.n197 585
R1355 B.n809 B.n808 585
R1356 B.n811 B.n809 585
R1357 B.n807 B.n202 585
R1358 B.n202 B.n201 585
R1359 B.n806 B.n805 585
R1360 B.n805 B.n804 585
R1361 B.n204 B.n203 585
R1362 B.n205 B.n204 585
R1363 B.n797 B.n796 585
R1364 B.n798 B.n797 585
R1365 B.n795 B.n210 585
R1366 B.n210 B.n209 585
R1367 B.n794 B.n793 585
R1368 B.n793 B.n792 585
R1369 B.n212 B.n211 585
R1370 B.n213 B.n212 585
R1371 B.n785 B.n784 585
R1372 B.n786 B.n785 585
R1373 B.n783 B.n217 585
R1374 B.n221 B.n217 585
R1375 B.n782 B.n781 585
R1376 B.n781 B.n780 585
R1377 B.n219 B.n218 585
R1378 B.n220 B.n219 585
R1379 B.n773 B.n772 585
R1380 B.n774 B.n773 585
R1381 B.n771 B.n226 585
R1382 B.n226 B.n225 585
R1383 B.n770 B.n769 585
R1384 B.n769 B.n768 585
R1385 B.n228 B.n227 585
R1386 B.n229 B.n228 585
R1387 B.n761 B.n760 585
R1388 B.n762 B.n761 585
R1389 B.n759 B.n234 585
R1390 B.n234 B.n233 585
R1391 B.n758 B.n757 585
R1392 B.n757 B.n756 585
R1393 B.n236 B.n235 585
R1394 B.n237 B.n236 585
R1395 B.n749 B.n748 585
R1396 B.n750 B.n749 585
R1397 B.n747 B.n242 585
R1398 B.n242 B.n241 585
R1399 B.n746 B.n745 585
R1400 B.n745 B.n744 585
R1401 B.n244 B.n243 585
R1402 B.n245 B.n244 585
R1403 B.n737 B.n736 585
R1404 B.n738 B.n737 585
R1405 B.n735 B.n250 585
R1406 B.n250 B.n249 585
R1407 B.n734 B.n733 585
R1408 B.n733 B.n732 585
R1409 B.n252 B.n251 585
R1410 B.n253 B.n252 585
R1411 B.n725 B.n724 585
R1412 B.n726 B.n725 585
R1413 B.n723 B.n258 585
R1414 B.n258 B.n257 585
R1415 B.n722 B.n721 585
R1416 B.n721 B.n720 585
R1417 B.n260 B.n259 585
R1418 B.n261 B.n260 585
R1419 B.n713 B.n712 585
R1420 B.n714 B.n713 585
R1421 B.n711 B.n266 585
R1422 B.n266 B.n265 585
R1423 B.n710 B.n709 585
R1424 B.n709 B.n708 585
R1425 B.n268 B.n267 585
R1426 B.n269 B.n268 585
R1427 B.n701 B.n700 585
R1428 B.n702 B.n701 585
R1429 B.n699 B.n273 585
R1430 B.n277 B.n273 585
R1431 B.n698 B.n697 585
R1432 B.n697 B.n696 585
R1433 B.n275 B.n274 585
R1434 B.n276 B.n275 585
R1435 B.n689 B.n688 585
R1436 B.n690 B.n689 585
R1437 B.n687 B.n282 585
R1438 B.n282 B.n281 585
R1439 B.n686 B.n685 585
R1440 B.n685 B.n684 585
R1441 B.n284 B.n283 585
R1442 B.n285 B.n284 585
R1443 B.n677 B.n676 585
R1444 B.n678 B.n677 585
R1445 B.n675 B.n290 585
R1446 B.n290 B.n289 585
R1447 B.n674 B.n673 585
R1448 B.n673 B.n672 585
R1449 B.n292 B.n291 585
R1450 B.n293 B.n292 585
R1451 B.n665 B.n664 585
R1452 B.n666 B.n665 585
R1453 B.n663 B.n298 585
R1454 B.n298 B.n297 585
R1455 B.n662 B.n661 585
R1456 B.n661 B.n660 585
R1457 B.n300 B.n299 585
R1458 B.n301 B.n300 585
R1459 B.n653 B.n652 585
R1460 B.n654 B.n653 585
R1461 B.n651 B.n306 585
R1462 B.n306 B.n305 585
R1463 B.n650 B.n649 585
R1464 B.n649 B.n648 585
R1465 B.n308 B.n307 585
R1466 B.n309 B.n308 585
R1467 B.n641 B.n640 585
R1468 B.n642 B.n641 585
R1469 B.n639 B.n314 585
R1470 B.n314 B.n313 585
R1471 B.n638 B.n637 585
R1472 B.n637 B.n636 585
R1473 B.n633 B.n318 585
R1474 B.n632 B.n631 585
R1475 B.n629 B.n319 585
R1476 B.n629 B.n317 585
R1477 B.n628 B.n627 585
R1478 B.n626 B.n625 585
R1479 B.n624 B.n321 585
R1480 B.n622 B.n621 585
R1481 B.n620 B.n322 585
R1482 B.n619 B.n618 585
R1483 B.n616 B.n323 585
R1484 B.n614 B.n613 585
R1485 B.n612 B.n324 585
R1486 B.n611 B.n610 585
R1487 B.n608 B.n325 585
R1488 B.n606 B.n605 585
R1489 B.n604 B.n326 585
R1490 B.n603 B.n602 585
R1491 B.n600 B.n327 585
R1492 B.n598 B.n597 585
R1493 B.n596 B.n328 585
R1494 B.n595 B.n594 585
R1495 B.n592 B.n329 585
R1496 B.n590 B.n589 585
R1497 B.n588 B.n330 585
R1498 B.n587 B.n586 585
R1499 B.n584 B.n331 585
R1500 B.n582 B.n581 585
R1501 B.n580 B.n332 585
R1502 B.n579 B.n578 585
R1503 B.n576 B.n333 585
R1504 B.n574 B.n573 585
R1505 B.n572 B.n334 585
R1506 B.n571 B.n570 585
R1507 B.n568 B.n335 585
R1508 B.n566 B.n565 585
R1509 B.n564 B.n336 585
R1510 B.n563 B.n562 585
R1511 B.n560 B.n337 585
R1512 B.n558 B.n557 585
R1513 B.n556 B.n338 585
R1514 B.n555 B.n554 585
R1515 B.n552 B.n339 585
R1516 B.n550 B.n549 585
R1517 B.n548 B.n340 585
R1518 B.n547 B.n546 585
R1519 B.n544 B.n341 585
R1520 B.n542 B.n541 585
R1521 B.n540 B.n342 585
R1522 B.n539 B.n538 585
R1523 B.n536 B.n343 585
R1524 B.n534 B.n533 585
R1525 B.n532 B.n344 585
R1526 B.n531 B.n530 585
R1527 B.n528 B.n345 585
R1528 B.n526 B.n525 585
R1529 B.n524 B.n346 585
R1530 B.n523 B.n522 585
R1531 B.n520 B.n347 585
R1532 B.n518 B.n517 585
R1533 B.n516 B.n348 585
R1534 B.n515 B.n514 585
R1535 B.n512 B.n352 585
R1536 B.n510 B.n509 585
R1537 B.n508 B.n353 585
R1538 B.n507 B.n506 585
R1539 B.n504 B.n354 585
R1540 B.n502 B.n501 585
R1541 B.n499 B.n355 585
R1542 B.n498 B.n497 585
R1543 B.n495 B.n358 585
R1544 B.n493 B.n492 585
R1545 B.n491 B.n359 585
R1546 B.n490 B.n489 585
R1547 B.n487 B.n360 585
R1548 B.n485 B.n484 585
R1549 B.n483 B.n361 585
R1550 B.n482 B.n481 585
R1551 B.n479 B.n362 585
R1552 B.n477 B.n476 585
R1553 B.n475 B.n363 585
R1554 B.n474 B.n473 585
R1555 B.n471 B.n364 585
R1556 B.n469 B.n468 585
R1557 B.n467 B.n365 585
R1558 B.n466 B.n465 585
R1559 B.n463 B.n366 585
R1560 B.n461 B.n460 585
R1561 B.n459 B.n367 585
R1562 B.n458 B.n457 585
R1563 B.n455 B.n368 585
R1564 B.n453 B.n452 585
R1565 B.n451 B.n369 585
R1566 B.n450 B.n449 585
R1567 B.n447 B.n370 585
R1568 B.n445 B.n444 585
R1569 B.n443 B.n371 585
R1570 B.n442 B.n441 585
R1571 B.n439 B.n372 585
R1572 B.n437 B.n436 585
R1573 B.n435 B.n373 585
R1574 B.n434 B.n433 585
R1575 B.n431 B.n374 585
R1576 B.n429 B.n428 585
R1577 B.n427 B.n375 585
R1578 B.n426 B.n425 585
R1579 B.n423 B.n376 585
R1580 B.n421 B.n420 585
R1581 B.n419 B.n377 585
R1582 B.n418 B.n417 585
R1583 B.n415 B.n378 585
R1584 B.n413 B.n412 585
R1585 B.n411 B.n379 585
R1586 B.n410 B.n409 585
R1587 B.n407 B.n380 585
R1588 B.n405 B.n404 585
R1589 B.n403 B.n381 585
R1590 B.n402 B.n401 585
R1591 B.n399 B.n382 585
R1592 B.n397 B.n396 585
R1593 B.n395 B.n383 585
R1594 B.n394 B.n393 585
R1595 B.n391 B.n384 585
R1596 B.n389 B.n388 585
R1597 B.n387 B.n386 585
R1598 B.n316 B.n315 585
R1599 B.n635 B.n634 585
R1600 B.n636 B.n635 585
R1601 B.n312 B.n311 585
R1602 B.n313 B.n312 585
R1603 B.n644 B.n643 585
R1604 B.n643 B.n642 585
R1605 B.n645 B.n310 585
R1606 B.n310 B.n309 585
R1607 B.n647 B.n646 585
R1608 B.n648 B.n647 585
R1609 B.n304 B.n303 585
R1610 B.n305 B.n304 585
R1611 B.n656 B.n655 585
R1612 B.n655 B.n654 585
R1613 B.n657 B.n302 585
R1614 B.n302 B.n301 585
R1615 B.n659 B.n658 585
R1616 B.n660 B.n659 585
R1617 B.n296 B.n295 585
R1618 B.n297 B.n296 585
R1619 B.n668 B.n667 585
R1620 B.n667 B.n666 585
R1621 B.n669 B.n294 585
R1622 B.n294 B.n293 585
R1623 B.n671 B.n670 585
R1624 B.n672 B.n671 585
R1625 B.n288 B.n287 585
R1626 B.n289 B.n288 585
R1627 B.n680 B.n679 585
R1628 B.n679 B.n678 585
R1629 B.n681 B.n286 585
R1630 B.n286 B.n285 585
R1631 B.n683 B.n682 585
R1632 B.n684 B.n683 585
R1633 B.n280 B.n279 585
R1634 B.n281 B.n280 585
R1635 B.n692 B.n691 585
R1636 B.n691 B.n690 585
R1637 B.n693 B.n278 585
R1638 B.n278 B.n276 585
R1639 B.n695 B.n694 585
R1640 B.n696 B.n695 585
R1641 B.n272 B.n271 585
R1642 B.n277 B.n272 585
R1643 B.n704 B.n703 585
R1644 B.n703 B.n702 585
R1645 B.n705 B.n270 585
R1646 B.n270 B.n269 585
R1647 B.n707 B.n706 585
R1648 B.n708 B.n707 585
R1649 B.n264 B.n263 585
R1650 B.n265 B.n264 585
R1651 B.n716 B.n715 585
R1652 B.n715 B.n714 585
R1653 B.n717 B.n262 585
R1654 B.n262 B.n261 585
R1655 B.n719 B.n718 585
R1656 B.n720 B.n719 585
R1657 B.n256 B.n255 585
R1658 B.n257 B.n256 585
R1659 B.n728 B.n727 585
R1660 B.n727 B.n726 585
R1661 B.n729 B.n254 585
R1662 B.n254 B.n253 585
R1663 B.n731 B.n730 585
R1664 B.n732 B.n731 585
R1665 B.n248 B.n247 585
R1666 B.n249 B.n248 585
R1667 B.n740 B.n739 585
R1668 B.n739 B.n738 585
R1669 B.n741 B.n246 585
R1670 B.n246 B.n245 585
R1671 B.n743 B.n742 585
R1672 B.n744 B.n743 585
R1673 B.n240 B.n239 585
R1674 B.n241 B.n240 585
R1675 B.n752 B.n751 585
R1676 B.n751 B.n750 585
R1677 B.n753 B.n238 585
R1678 B.n238 B.n237 585
R1679 B.n755 B.n754 585
R1680 B.n756 B.n755 585
R1681 B.n232 B.n231 585
R1682 B.n233 B.n232 585
R1683 B.n764 B.n763 585
R1684 B.n763 B.n762 585
R1685 B.n765 B.n230 585
R1686 B.n230 B.n229 585
R1687 B.n767 B.n766 585
R1688 B.n768 B.n767 585
R1689 B.n224 B.n223 585
R1690 B.n225 B.n224 585
R1691 B.n776 B.n775 585
R1692 B.n775 B.n774 585
R1693 B.n777 B.n222 585
R1694 B.n222 B.n220 585
R1695 B.n779 B.n778 585
R1696 B.n780 B.n779 585
R1697 B.n216 B.n215 585
R1698 B.n221 B.n216 585
R1699 B.n788 B.n787 585
R1700 B.n787 B.n786 585
R1701 B.n789 B.n214 585
R1702 B.n214 B.n213 585
R1703 B.n791 B.n790 585
R1704 B.n792 B.n791 585
R1705 B.n208 B.n207 585
R1706 B.n209 B.n208 585
R1707 B.n800 B.n799 585
R1708 B.n799 B.n798 585
R1709 B.n801 B.n206 585
R1710 B.n206 B.n205 585
R1711 B.n803 B.n802 585
R1712 B.n804 B.n803 585
R1713 B.n200 B.n199 585
R1714 B.n201 B.n200 585
R1715 B.n813 B.n812 585
R1716 B.n812 B.n811 585
R1717 B.n814 B.n198 585
R1718 B.n810 B.n198 585
R1719 B.n816 B.n815 585
R1720 B.n817 B.n816 585
R1721 B.n193 B.n192 585
R1722 B.n194 B.n193 585
R1723 B.n826 B.n825 585
R1724 B.n825 B.n824 585
R1725 B.n827 B.n191 585
R1726 B.n191 B.n190 585
R1727 B.n829 B.n828 585
R1728 B.n830 B.n829 585
R1729 B.n2 B.n0 585
R1730 B.n4 B.n2 585
R1731 B.n3 B.n1 585
R1732 B.n1299 B.n3 585
R1733 B.n1297 B.n1296 585
R1734 B.n1298 B.n1297 585
R1735 B.n1295 B.n9 585
R1736 B.n9 B.n8 585
R1737 B.n1294 B.n1293 585
R1738 B.n1293 B.n1292 585
R1739 B.n11 B.n10 585
R1740 B.n1291 B.n11 585
R1741 B.n1289 B.n1288 585
R1742 B.n1290 B.n1289 585
R1743 B.n1287 B.n15 585
R1744 B.n18 B.n15 585
R1745 B.n1286 B.n1285 585
R1746 B.n1285 B.n1284 585
R1747 B.n17 B.n16 585
R1748 B.n1283 B.n17 585
R1749 B.n1281 B.n1280 585
R1750 B.n1282 B.n1281 585
R1751 B.n1279 B.n23 585
R1752 B.n23 B.n22 585
R1753 B.n1278 B.n1277 585
R1754 B.n1277 B.n1276 585
R1755 B.n25 B.n24 585
R1756 B.n1275 B.n25 585
R1757 B.n1273 B.n1272 585
R1758 B.n1274 B.n1273 585
R1759 B.n1271 B.n30 585
R1760 B.n30 B.n29 585
R1761 B.n1270 B.n1269 585
R1762 B.n1269 B.n1268 585
R1763 B.n32 B.n31 585
R1764 B.n1267 B.n32 585
R1765 B.n1265 B.n1264 585
R1766 B.n1266 B.n1265 585
R1767 B.n1263 B.n37 585
R1768 B.n37 B.n36 585
R1769 B.n1262 B.n1261 585
R1770 B.n1261 B.n1260 585
R1771 B.n39 B.n38 585
R1772 B.n1259 B.n39 585
R1773 B.n1257 B.n1256 585
R1774 B.n1258 B.n1257 585
R1775 B.n1255 B.n44 585
R1776 B.n44 B.n43 585
R1777 B.n1254 B.n1253 585
R1778 B.n1253 B.n1252 585
R1779 B.n46 B.n45 585
R1780 B.n1251 B.n46 585
R1781 B.n1249 B.n1248 585
R1782 B.n1250 B.n1249 585
R1783 B.n1247 B.n51 585
R1784 B.n51 B.n50 585
R1785 B.n1246 B.n1245 585
R1786 B.n1245 B.n1244 585
R1787 B.n53 B.n52 585
R1788 B.n1243 B.n53 585
R1789 B.n1241 B.n1240 585
R1790 B.n1242 B.n1241 585
R1791 B.n1239 B.n58 585
R1792 B.n58 B.n57 585
R1793 B.n1238 B.n1237 585
R1794 B.n1237 B.n1236 585
R1795 B.n60 B.n59 585
R1796 B.n1235 B.n60 585
R1797 B.n1233 B.n1232 585
R1798 B.n1234 B.n1233 585
R1799 B.n1231 B.n65 585
R1800 B.n65 B.n64 585
R1801 B.n1230 B.n1229 585
R1802 B.n1229 B.n1228 585
R1803 B.n67 B.n66 585
R1804 B.n1227 B.n67 585
R1805 B.n1225 B.n1224 585
R1806 B.n1226 B.n1225 585
R1807 B.n1223 B.n72 585
R1808 B.n72 B.n71 585
R1809 B.n1222 B.n1221 585
R1810 B.n1221 B.n1220 585
R1811 B.n74 B.n73 585
R1812 B.n1219 B.n74 585
R1813 B.n1217 B.n1216 585
R1814 B.n1218 B.n1217 585
R1815 B.n1215 B.n79 585
R1816 B.n79 B.n78 585
R1817 B.n1214 B.n1213 585
R1818 B.n1213 B.n1212 585
R1819 B.n81 B.n80 585
R1820 B.n1211 B.n81 585
R1821 B.n1209 B.n1208 585
R1822 B.n1210 B.n1209 585
R1823 B.n1207 B.n86 585
R1824 B.n86 B.n85 585
R1825 B.n1206 B.n1205 585
R1826 B.n1205 B.n1204 585
R1827 B.n88 B.n87 585
R1828 B.n1203 B.n88 585
R1829 B.n1201 B.n1200 585
R1830 B.n1202 B.n1201 585
R1831 B.n1199 B.n93 585
R1832 B.n93 B.n92 585
R1833 B.n1198 B.n1197 585
R1834 B.n1197 B.n1196 585
R1835 B.n95 B.n94 585
R1836 B.n1195 B.n95 585
R1837 B.n1193 B.n1192 585
R1838 B.n1194 B.n1193 585
R1839 B.n1191 B.n100 585
R1840 B.n100 B.n99 585
R1841 B.n1190 B.n1189 585
R1842 B.n1189 B.n1188 585
R1843 B.n102 B.n101 585
R1844 B.n1187 B.n102 585
R1845 B.n1185 B.n1184 585
R1846 B.n1186 B.n1185 585
R1847 B.n1183 B.n107 585
R1848 B.n107 B.n106 585
R1849 B.n1182 B.n1181 585
R1850 B.n1181 B.n1180 585
R1851 B.n109 B.n108 585
R1852 B.n1179 B.n109 585
R1853 B.n1177 B.n1176 585
R1854 B.n1178 B.n1177 585
R1855 B.n1175 B.n114 585
R1856 B.n114 B.n113 585
R1857 B.n1174 B.n1173 585
R1858 B.n1173 B.n1172 585
R1859 B.n116 B.n115 585
R1860 B.n1171 B.n116 585
R1861 B.n1169 B.n1168 585
R1862 B.n1170 B.n1169 585
R1863 B.n1302 B.n1301 585
R1864 B.n1301 B.n1300 585
R1865 B.n356 B.t12 438.156
R1866 B.n158 B.t18 438.156
R1867 B.n349 B.t15 438.156
R1868 B.n150 B.t21 438.156
R1869 B.n635 B.n318 430.038
R1870 B.n1169 B.n121 430.038
R1871 B.n637 B.n316 430.038
R1872 B.n918 B.n119 430.038
R1873 B.n357 B.t11 374.738
R1874 B.n159 B.t19 374.738
R1875 B.n350 B.t14 374.738
R1876 B.n151 B.t22 374.738
R1877 B.n356 B.t9 351.06
R1878 B.n349 B.t13 351.06
R1879 B.n150 B.t20 351.06
R1880 B.n158 B.t16 351.06
R1881 B.n919 B.n120 256.663
R1882 B.n925 B.n120 256.663
R1883 B.n927 B.n120 256.663
R1884 B.n933 B.n120 256.663
R1885 B.n935 B.n120 256.663
R1886 B.n941 B.n120 256.663
R1887 B.n943 B.n120 256.663
R1888 B.n949 B.n120 256.663
R1889 B.n951 B.n120 256.663
R1890 B.n957 B.n120 256.663
R1891 B.n959 B.n120 256.663
R1892 B.n965 B.n120 256.663
R1893 B.n967 B.n120 256.663
R1894 B.n973 B.n120 256.663
R1895 B.n975 B.n120 256.663
R1896 B.n981 B.n120 256.663
R1897 B.n983 B.n120 256.663
R1898 B.n989 B.n120 256.663
R1899 B.n991 B.n120 256.663
R1900 B.n997 B.n120 256.663
R1901 B.n999 B.n120 256.663
R1902 B.n1005 B.n120 256.663
R1903 B.n1007 B.n120 256.663
R1904 B.n1013 B.n120 256.663
R1905 B.n1015 B.n120 256.663
R1906 B.n1021 B.n120 256.663
R1907 B.n1023 B.n120 256.663
R1908 B.n1029 B.n120 256.663
R1909 B.n1031 B.n120 256.663
R1910 B.n1038 B.n120 256.663
R1911 B.n1040 B.n120 256.663
R1912 B.n1046 B.n120 256.663
R1913 B.n153 B.n120 256.663
R1914 B.n1052 B.n120 256.663
R1915 B.n1058 B.n120 256.663
R1916 B.n1060 B.n120 256.663
R1917 B.n1066 B.n120 256.663
R1918 B.n1068 B.n120 256.663
R1919 B.n1074 B.n120 256.663
R1920 B.n1076 B.n120 256.663
R1921 B.n1082 B.n120 256.663
R1922 B.n1084 B.n120 256.663
R1923 B.n1090 B.n120 256.663
R1924 B.n1092 B.n120 256.663
R1925 B.n1098 B.n120 256.663
R1926 B.n1100 B.n120 256.663
R1927 B.n1106 B.n120 256.663
R1928 B.n1108 B.n120 256.663
R1929 B.n1114 B.n120 256.663
R1930 B.n1116 B.n120 256.663
R1931 B.n1122 B.n120 256.663
R1932 B.n1124 B.n120 256.663
R1933 B.n1130 B.n120 256.663
R1934 B.n1132 B.n120 256.663
R1935 B.n1138 B.n120 256.663
R1936 B.n1140 B.n120 256.663
R1937 B.n1146 B.n120 256.663
R1938 B.n1148 B.n120 256.663
R1939 B.n1154 B.n120 256.663
R1940 B.n1156 B.n120 256.663
R1941 B.n1162 B.n120 256.663
R1942 B.n1164 B.n120 256.663
R1943 B.n630 B.n317 256.663
R1944 B.n320 B.n317 256.663
R1945 B.n623 B.n317 256.663
R1946 B.n617 B.n317 256.663
R1947 B.n615 B.n317 256.663
R1948 B.n609 B.n317 256.663
R1949 B.n607 B.n317 256.663
R1950 B.n601 B.n317 256.663
R1951 B.n599 B.n317 256.663
R1952 B.n593 B.n317 256.663
R1953 B.n591 B.n317 256.663
R1954 B.n585 B.n317 256.663
R1955 B.n583 B.n317 256.663
R1956 B.n577 B.n317 256.663
R1957 B.n575 B.n317 256.663
R1958 B.n569 B.n317 256.663
R1959 B.n567 B.n317 256.663
R1960 B.n561 B.n317 256.663
R1961 B.n559 B.n317 256.663
R1962 B.n553 B.n317 256.663
R1963 B.n551 B.n317 256.663
R1964 B.n545 B.n317 256.663
R1965 B.n543 B.n317 256.663
R1966 B.n537 B.n317 256.663
R1967 B.n535 B.n317 256.663
R1968 B.n529 B.n317 256.663
R1969 B.n527 B.n317 256.663
R1970 B.n521 B.n317 256.663
R1971 B.n519 B.n317 256.663
R1972 B.n513 B.n317 256.663
R1973 B.n511 B.n317 256.663
R1974 B.n505 B.n317 256.663
R1975 B.n503 B.n317 256.663
R1976 B.n496 B.n317 256.663
R1977 B.n494 B.n317 256.663
R1978 B.n488 B.n317 256.663
R1979 B.n486 B.n317 256.663
R1980 B.n480 B.n317 256.663
R1981 B.n478 B.n317 256.663
R1982 B.n472 B.n317 256.663
R1983 B.n470 B.n317 256.663
R1984 B.n464 B.n317 256.663
R1985 B.n462 B.n317 256.663
R1986 B.n456 B.n317 256.663
R1987 B.n454 B.n317 256.663
R1988 B.n448 B.n317 256.663
R1989 B.n446 B.n317 256.663
R1990 B.n440 B.n317 256.663
R1991 B.n438 B.n317 256.663
R1992 B.n432 B.n317 256.663
R1993 B.n430 B.n317 256.663
R1994 B.n424 B.n317 256.663
R1995 B.n422 B.n317 256.663
R1996 B.n416 B.n317 256.663
R1997 B.n414 B.n317 256.663
R1998 B.n408 B.n317 256.663
R1999 B.n406 B.n317 256.663
R2000 B.n400 B.n317 256.663
R2001 B.n398 B.n317 256.663
R2002 B.n392 B.n317 256.663
R2003 B.n390 B.n317 256.663
R2004 B.n385 B.n317 256.663
R2005 B.n635 B.n312 163.367
R2006 B.n643 B.n312 163.367
R2007 B.n643 B.n310 163.367
R2008 B.n647 B.n310 163.367
R2009 B.n647 B.n304 163.367
R2010 B.n655 B.n304 163.367
R2011 B.n655 B.n302 163.367
R2012 B.n659 B.n302 163.367
R2013 B.n659 B.n296 163.367
R2014 B.n667 B.n296 163.367
R2015 B.n667 B.n294 163.367
R2016 B.n671 B.n294 163.367
R2017 B.n671 B.n288 163.367
R2018 B.n679 B.n288 163.367
R2019 B.n679 B.n286 163.367
R2020 B.n683 B.n286 163.367
R2021 B.n683 B.n280 163.367
R2022 B.n691 B.n280 163.367
R2023 B.n691 B.n278 163.367
R2024 B.n695 B.n278 163.367
R2025 B.n695 B.n272 163.367
R2026 B.n703 B.n272 163.367
R2027 B.n703 B.n270 163.367
R2028 B.n707 B.n270 163.367
R2029 B.n707 B.n264 163.367
R2030 B.n715 B.n264 163.367
R2031 B.n715 B.n262 163.367
R2032 B.n719 B.n262 163.367
R2033 B.n719 B.n256 163.367
R2034 B.n727 B.n256 163.367
R2035 B.n727 B.n254 163.367
R2036 B.n731 B.n254 163.367
R2037 B.n731 B.n248 163.367
R2038 B.n739 B.n248 163.367
R2039 B.n739 B.n246 163.367
R2040 B.n743 B.n246 163.367
R2041 B.n743 B.n240 163.367
R2042 B.n751 B.n240 163.367
R2043 B.n751 B.n238 163.367
R2044 B.n755 B.n238 163.367
R2045 B.n755 B.n232 163.367
R2046 B.n763 B.n232 163.367
R2047 B.n763 B.n230 163.367
R2048 B.n767 B.n230 163.367
R2049 B.n767 B.n224 163.367
R2050 B.n775 B.n224 163.367
R2051 B.n775 B.n222 163.367
R2052 B.n779 B.n222 163.367
R2053 B.n779 B.n216 163.367
R2054 B.n787 B.n216 163.367
R2055 B.n787 B.n214 163.367
R2056 B.n791 B.n214 163.367
R2057 B.n791 B.n208 163.367
R2058 B.n799 B.n208 163.367
R2059 B.n799 B.n206 163.367
R2060 B.n803 B.n206 163.367
R2061 B.n803 B.n200 163.367
R2062 B.n812 B.n200 163.367
R2063 B.n812 B.n198 163.367
R2064 B.n816 B.n198 163.367
R2065 B.n816 B.n193 163.367
R2066 B.n825 B.n193 163.367
R2067 B.n825 B.n191 163.367
R2068 B.n829 B.n191 163.367
R2069 B.n829 B.n2 163.367
R2070 B.n1301 B.n2 163.367
R2071 B.n1301 B.n3 163.367
R2072 B.n1297 B.n3 163.367
R2073 B.n1297 B.n9 163.367
R2074 B.n1293 B.n9 163.367
R2075 B.n1293 B.n11 163.367
R2076 B.n1289 B.n11 163.367
R2077 B.n1289 B.n15 163.367
R2078 B.n1285 B.n15 163.367
R2079 B.n1285 B.n17 163.367
R2080 B.n1281 B.n17 163.367
R2081 B.n1281 B.n23 163.367
R2082 B.n1277 B.n23 163.367
R2083 B.n1277 B.n25 163.367
R2084 B.n1273 B.n25 163.367
R2085 B.n1273 B.n30 163.367
R2086 B.n1269 B.n30 163.367
R2087 B.n1269 B.n32 163.367
R2088 B.n1265 B.n32 163.367
R2089 B.n1265 B.n37 163.367
R2090 B.n1261 B.n37 163.367
R2091 B.n1261 B.n39 163.367
R2092 B.n1257 B.n39 163.367
R2093 B.n1257 B.n44 163.367
R2094 B.n1253 B.n44 163.367
R2095 B.n1253 B.n46 163.367
R2096 B.n1249 B.n46 163.367
R2097 B.n1249 B.n51 163.367
R2098 B.n1245 B.n51 163.367
R2099 B.n1245 B.n53 163.367
R2100 B.n1241 B.n53 163.367
R2101 B.n1241 B.n58 163.367
R2102 B.n1237 B.n58 163.367
R2103 B.n1237 B.n60 163.367
R2104 B.n1233 B.n60 163.367
R2105 B.n1233 B.n65 163.367
R2106 B.n1229 B.n65 163.367
R2107 B.n1229 B.n67 163.367
R2108 B.n1225 B.n67 163.367
R2109 B.n1225 B.n72 163.367
R2110 B.n1221 B.n72 163.367
R2111 B.n1221 B.n74 163.367
R2112 B.n1217 B.n74 163.367
R2113 B.n1217 B.n79 163.367
R2114 B.n1213 B.n79 163.367
R2115 B.n1213 B.n81 163.367
R2116 B.n1209 B.n81 163.367
R2117 B.n1209 B.n86 163.367
R2118 B.n1205 B.n86 163.367
R2119 B.n1205 B.n88 163.367
R2120 B.n1201 B.n88 163.367
R2121 B.n1201 B.n93 163.367
R2122 B.n1197 B.n93 163.367
R2123 B.n1197 B.n95 163.367
R2124 B.n1193 B.n95 163.367
R2125 B.n1193 B.n100 163.367
R2126 B.n1189 B.n100 163.367
R2127 B.n1189 B.n102 163.367
R2128 B.n1185 B.n102 163.367
R2129 B.n1185 B.n107 163.367
R2130 B.n1181 B.n107 163.367
R2131 B.n1181 B.n109 163.367
R2132 B.n1177 B.n109 163.367
R2133 B.n1177 B.n114 163.367
R2134 B.n1173 B.n114 163.367
R2135 B.n1173 B.n116 163.367
R2136 B.n1169 B.n116 163.367
R2137 B.n631 B.n629 163.367
R2138 B.n629 B.n628 163.367
R2139 B.n625 B.n624 163.367
R2140 B.n622 B.n322 163.367
R2141 B.n618 B.n616 163.367
R2142 B.n614 B.n324 163.367
R2143 B.n610 B.n608 163.367
R2144 B.n606 B.n326 163.367
R2145 B.n602 B.n600 163.367
R2146 B.n598 B.n328 163.367
R2147 B.n594 B.n592 163.367
R2148 B.n590 B.n330 163.367
R2149 B.n586 B.n584 163.367
R2150 B.n582 B.n332 163.367
R2151 B.n578 B.n576 163.367
R2152 B.n574 B.n334 163.367
R2153 B.n570 B.n568 163.367
R2154 B.n566 B.n336 163.367
R2155 B.n562 B.n560 163.367
R2156 B.n558 B.n338 163.367
R2157 B.n554 B.n552 163.367
R2158 B.n550 B.n340 163.367
R2159 B.n546 B.n544 163.367
R2160 B.n542 B.n342 163.367
R2161 B.n538 B.n536 163.367
R2162 B.n534 B.n344 163.367
R2163 B.n530 B.n528 163.367
R2164 B.n526 B.n346 163.367
R2165 B.n522 B.n520 163.367
R2166 B.n518 B.n348 163.367
R2167 B.n514 B.n512 163.367
R2168 B.n510 B.n353 163.367
R2169 B.n506 B.n504 163.367
R2170 B.n502 B.n355 163.367
R2171 B.n497 B.n495 163.367
R2172 B.n493 B.n359 163.367
R2173 B.n489 B.n487 163.367
R2174 B.n485 B.n361 163.367
R2175 B.n481 B.n479 163.367
R2176 B.n477 B.n363 163.367
R2177 B.n473 B.n471 163.367
R2178 B.n469 B.n365 163.367
R2179 B.n465 B.n463 163.367
R2180 B.n461 B.n367 163.367
R2181 B.n457 B.n455 163.367
R2182 B.n453 B.n369 163.367
R2183 B.n449 B.n447 163.367
R2184 B.n445 B.n371 163.367
R2185 B.n441 B.n439 163.367
R2186 B.n437 B.n373 163.367
R2187 B.n433 B.n431 163.367
R2188 B.n429 B.n375 163.367
R2189 B.n425 B.n423 163.367
R2190 B.n421 B.n377 163.367
R2191 B.n417 B.n415 163.367
R2192 B.n413 B.n379 163.367
R2193 B.n409 B.n407 163.367
R2194 B.n405 B.n381 163.367
R2195 B.n401 B.n399 163.367
R2196 B.n397 B.n383 163.367
R2197 B.n393 B.n391 163.367
R2198 B.n389 B.n386 163.367
R2199 B.n637 B.n314 163.367
R2200 B.n641 B.n314 163.367
R2201 B.n641 B.n308 163.367
R2202 B.n649 B.n308 163.367
R2203 B.n649 B.n306 163.367
R2204 B.n653 B.n306 163.367
R2205 B.n653 B.n300 163.367
R2206 B.n661 B.n300 163.367
R2207 B.n661 B.n298 163.367
R2208 B.n665 B.n298 163.367
R2209 B.n665 B.n292 163.367
R2210 B.n673 B.n292 163.367
R2211 B.n673 B.n290 163.367
R2212 B.n677 B.n290 163.367
R2213 B.n677 B.n284 163.367
R2214 B.n685 B.n284 163.367
R2215 B.n685 B.n282 163.367
R2216 B.n689 B.n282 163.367
R2217 B.n689 B.n275 163.367
R2218 B.n697 B.n275 163.367
R2219 B.n697 B.n273 163.367
R2220 B.n701 B.n273 163.367
R2221 B.n701 B.n268 163.367
R2222 B.n709 B.n268 163.367
R2223 B.n709 B.n266 163.367
R2224 B.n713 B.n266 163.367
R2225 B.n713 B.n260 163.367
R2226 B.n721 B.n260 163.367
R2227 B.n721 B.n258 163.367
R2228 B.n725 B.n258 163.367
R2229 B.n725 B.n252 163.367
R2230 B.n733 B.n252 163.367
R2231 B.n733 B.n250 163.367
R2232 B.n737 B.n250 163.367
R2233 B.n737 B.n244 163.367
R2234 B.n745 B.n244 163.367
R2235 B.n745 B.n242 163.367
R2236 B.n749 B.n242 163.367
R2237 B.n749 B.n236 163.367
R2238 B.n757 B.n236 163.367
R2239 B.n757 B.n234 163.367
R2240 B.n761 B.n234 163.367
R2241 B.n761 B.n228 163.367
R2242 B.n769 B.n228 163.367
R2243 B.n769 B.n226 163.367
R2244 B.n773 B.n226 163.367
R2245 B.n773 B.n219 163.367
R2246 B.n781 B.n219 163.367
R2247 B.n781 B.n217 163.367
R2248 B.n785 B.n217 163.367
R2249 B.n785 B.n212 163.367
R2250 B.n793 B.n212 163.367
R2251 B.n793 B.n210 163.367
R2252 B.n797 B.n210 163.367
R2253 B.n797 B.n204 163.367
R2254 B.n805 B.n204 163.367
R2255 B.n805 B.n202 163.367
R2256 B.n809 B.n202 163.367
R2257 B.n809 B.n197 163.367
R2258 B.n818 B.n197 163.367
R2259 B.n818 B.n195 163.367
R2260 B.n823 B.n195 163.367
R2261 B.n823 B.n189 163.367
R2262 B.n831 B.n189 163.367
R2263 B.n832 B.n831 163.367
R2264 B.n832 B.n5 163.367
R2265 B.n6 B.n5 163.367
R2266 B.n7 B.n6 163.367
R2267 B.n837 B.n7 163.367
R2268 B.n837 B.n12 163.367
R2269 B.n13 B.n12 163.367
R2270 B.n14 B.n13 163.367
R2271 B.n842 B.n14 163.367
R2272 B.n842 B.n19 163.367
R2273 B.n20 B.n19 163.367
R2274 B.n21 B.n20 163.367
R2275 B.n847 B.n21 163.367
R2276 B.n847 B.n26 163.367
R2277 B.n27 B.n26 163.367
R2278 B.n28 B.n27 163.367
R2279 B.n852 B.n28 163.367
R2280 B.n852 B.n33 163.367
R2281 B.n34 B.n33 163.367
R2282 B.n35 B.n34 163.367
R2283 B.n857 B.n35 163.367
R2284 B.n857 B.n40 163.367
R2285 B.n41 B.n40 163.367
R2286 B.n42 B.n41 163.367
R2287 B.n862 B.n42 163.367
R2288 B.n862 B.n47 163.367
R2289 B.n48 B.n47 163.367
R2290 B.n49 B.n48 163.367
R2291 B.n867 B.n49 163.367
R2292 B.n867 B.n54 163.367
R2293 B.n55 B.n54 163.367
R2294 B.n56 B.n55 163.367
R2295 B.n872 B.n56 163.367
R2296 B.n872 B.n61 163.367
R2297 B.n62 B.n61 163.367
R2298 B.n63 B.n62 163.367
R2299 B.n877 B.n63 163.367
R2300 B.n877 B.n68 163.367
R2301 B.n69 B.n68 163.367
R2302 B.n70 B.n69 163.367
R2303 B.n882 B.n70 163.367
R2304 B.n882 B.n75 163.367
R2305 B.n76 B.n75 163.367
R2306 B.n77 B.n76 163.367
R2307 B.n887 B.n77 163.367
R2308 B.n887 B.n82 163.367
R2309 B.n83 B.n82 163.367
R2310 B.n84 B.n83 163.367
R2311 B.n892 B.n84 163.367
R2312 B.n892 B.n89 163.367
R2313 B.n90 B.n89 163.367
R2314 B.n91 B.n90 163.367
R2315 B.n897 B.n91 163.367
R2316 B.n897 B.n96 163.367
R2317 B.n97 B.n96 163.367
R2318 B.n98 B.n97 163.367
R2319 B.n902 B.n98 163.367
R2320 B.n902 B.n103 163.367
R2321 B.n104 B.n103 163.367
R2322 B.n105 B.n104 163.367
R2323 B.n907 B.n105 163.367
R2324 B.n907 B.n110 163.367
R2325 B.n111 B.n110 163.367
R2326 B.n112 B.n111 163.367
R2327 B.n912 B.n112 163.367
R2328 B.n912 B.n117 163.367
R2329 B.n118 B.n117 163.367
R2330 B.n119 B.n118 163.367
R2331 B.n1165 B.n1163 163.367
R2332 B.n1161 B.n123 163.367
R2333 B.n1157 B.n1155 163.367
R2334 B.n1153 B.n125 163.367
R2335 B.n1149 B.n1147 163.367
R2336 B.n1145 B.n127 163.367
R2337 B.n1141 B.n1139 163.367
R2338 B.n1137 B.n129 163.367
R2339 B.n1133 B.n1131 163.367
R2340 B.n1129 B.n131 163.367
R2341 B.n1125 B.n1123 163.367
R2342 B.n1121 B.n133 163.367
R2343 B.n1117 B.n1115 163.367
R2344 B.n1113 B.n135 163.367
R2345 B.n1109 B.n1107 163.367
R2346 B.n1105 B.n137 163.367
R2347 B.n1101 B.n1099 163.367
R2348 B.n1097 B.n139 163.367
R2349 B.n1093 B.n1091 163.367
R2350 B.n1089 B.n141 163.367
R2351 B.n1085 B.n1083 163.367
R2352 B.n1081 B.n143 163.367
R2353 B.n1077 B.n1075 163.367
R2354 B.n1073 B.n145 163.367
R2355 B.n1069 B.n1067 163.367
R2356 B.n1065 B.n147 163.367
R2357 B.n1061 B.n1059 163.367
R2358 B.n1057 B.n149 163.367
R2359 B.n1053 B.n1051 163.367
R2360 B.n1048 B.n1047 163.367
R2361 B.n1045 B.n155 163.367
R2362 B.n1041 B.n1039 163.367
R2363 B.n1037 B.n157 163.367
R2364 B.n1032 B.n1030 163.367
R2365 B.n1028 B.n161 163.367
R2366 B.n1024 B.n1022 163.367
R2367 B.n1020 B.n163 163.367
R2368 B.n1016 B.n1014 163.367
R2369 B.n1012 B.n165 163.367
R2370 B.n1008 B.n1006 163.367
R2371 B.n1004 B.n167 163.367
R2372 B.n1000 B.n998 163.367
R2373 B.n996 B.n169 163.367
R2374 B.n992 B.n990 163.367
R2375 B.n988 B.n171 163.367
R2376 B.n984 B.n982 163.367
R2377 B.n980 B.n173 163.367
R2378 B.n976 B.n974 163.367
R2379 B.n972 B.n175 163.367
R2380 B.n968 B.n966 163.367
R2381 B.n964 B.n177 163.367
R2382 B.n960 B.n958 163.367
R2383 B.n956 B.n179 163.367
R2384 B.n952 B.n950 163.367
R2385 B.n948 B.n181 163.367
R2386 B.n944 B.n942 163.367
R2387 B.n940 B.n183 163.367
R2388 B.n936 B.n934 163.367
R2389 B.n932 B.n185 163.367
R2390 B.n928 B.n926 163.367
R2391 B.n924 B.n187 163.367
R2392 B.n920 B.n918 163.367
R2393 B.n630 B.n318 71.676
R2394 B.n628 B.n320 71.676
R2395 B.n624 B.n623 71.676
R2396 B.n617 B.n322 71.676
R2397 B.n616 B.n615 71.676
R2398 B.n609 B.n324 71.676
R2399 B.n608 B.n607 71.676
R2400 B.n601 B.n326 71.676
R2401 B.n600 B.n599 71.676
R2402 B.n593 B.n328 71.676
R2403 B.n592 B.n591 71.676
R2404 B.n585 B.n330 71.676
R2405 B.n584 B.n583 71.676
R2406 B.n577 B.n332 71.676
R2407 B.n576 B.n575 71.676
R2408 B.n569 B.n334 71.676
R2409 B.n568 B.n567 71.676
R2410 B.n561 B.n336 71.676
R2411 B.n560 B.n559 71.676
R2412 B.n553 B.n338 71.676
R2413 B.n552 B.n551 71.676
R2414 B.n545 B.n340 71.676
R2415 B.n544 B.n543 71.676
R2416 B.n537 B.n342 71.676
R2417 B.n536 B.n535 71.676
R2418 B.n529 B.n344 71.676
R2419 B.n528 B.n527 71.676
R2420 B.n521 B.n346 71.676
R2421 B.n520 B.n519 71.676
R2422 B.n513 B.n348 71.676
R2423 B.n512 B.n511 71.676
R2424 B.n505 B.n353 71.676
R2425 B.n504 B.n503 71.676
R2426 B.n496 B.n355 71.676
R2427 B.n495 B.n494 71.676
R2428 B.n488 B.n359 71.676
R2429 B.n487 B.n486 71.676
R2430 B.n480 B.n361 71.676
R2431 B.n479 B.n478 71.676
R2432 B.n472 B.n363 71.676
R2433 B.n471 B.n470 71.676
R2434 B.n464 B.n365 71.676
R2435 B.n463 B.n462 71.676
R2436 B.n456 B.n367 71.676
R2437 B.n455 B.n454 71.676
R2438 B.n448 B.n369 71.676
R2439 B.n447 B.n446 71.676
R2440 B.n440 B.n371 71.676
R2441 B.n439 B.n438 71.676
R2442 B.n432 B.n373 71.676
R2443 B.n431 B.n430 71.676
R2444 B.n424 B.n375 71.676
R2445 B.n423 B.n422 71.676
R2446 B.n416 B.n377 71.676
R2447 B.n415 B.n414 71.676
R2448 B.n408 B.n379 71.676
R2449 B.n407 B.n406 71.676
R2450 B.n400 B.n381 71.676
R2451 B.n399 B.n398 71.676
R2452 B.n392 B.n383 71.676
R2453 B.n391 B.n390 71.676
R2454 B.n386 B.n385 71.676
R2455 B.n1164 B.n121 71.676
R2456 B.n1163 B.n1162 71.676
R2457 B.n1156 B.n123 71.676
R2458 B.n1155 B.n1154 71.676
R2459 B.n1148 B.n125 71.676
R2460 B.n1147 B.n1146 71.676
R2461 B.n1140 B.n127 71.676
R2462 B.n1139 B.n1138 71.676
R2463 B.n1132 B.n129 71.676
R2464 B.n1131 B.n1130 71.676
R2465 B.n1124 B.n131 71.676
R2466 B.n1123 B.n1122 71.676
R2467 B.n1116 B.n133 71.676
R2468 B.n1115 B.n1114 71.676
R2469 B.n1108 B.n135 71.676
R2470 B.n1107 B.n1106 71.676
R2471 B.n1100 B.n137 71.676
R2472 B.n1099 B.n1098 71.676
R2473 B.n1092 B.n139 71.676
R2474 B.n1091 B.n1090 71.676
R2475 B.n1084 B.n141 71.676
R2476 B.n1083 B.n1082 71.676
R2477 B.n1076 B.n143 71.676
R2478 B.n1075 B.n1074 71.676
R2479 B.n1068 B.n145 71.676
R2480 B.n1067 B.n1066 71.676
R2481 B.n1060 B.n147 71.676
R2482 B.n1059 B.n1058 71.676
R2483 B.n1052 B.n149 71.676
R2484 B.n1051 B.n153 71.676
R2485 B.n1047 B.n1046 71.676
R2486 B.n1040 B.n155 71.676
R2487 B.n1039 B.n1038 71.676
R2488 B.n1031 B.n157 71.676
R2489 B.n1030 B.n1029 71.676
R2490 B.n1023 B.n161 71.676
R2491 B.n1022 B.n1021 71.676
R2492 B.n1015 B.n163 71.676
R2493 B.n1014 B.n1013 71.676
R2494 B.n1007 B.n165 71.676
R2495 B.n1006 B.n1005 71.676
R2496 B.n999 B.n167 71.676
R2497 B.n998 B.n997 71.676
R2498 B.n991 B.n169 71.676
R2499 B.n990 B.n989 71.676
R2500 B.n983 B.n171 71.676
R2501 B.n982 B.n981 71.676
R2502 B.n975 B.n173 71.676
R2503 B.n974 B.n973 71.676
R2504 B.n967 B.n175 71.676
R2505 B.n966 B.n965 71.676
R2506 B.n959 B.n177 71.676
R2507 B.n958 B.n957 71.676
R2508 B.n951 B.n179 71.676
R2509 B.n950 B.n949 71.676
R2510 B.n943 B.n181 71.676
R2511 B.n942 B.n941 71.676
R2512 B.n935 B.n183 71.676
R2513 B.n934 B.n933 71.676
R2514 B.n927 B.n185 71.676
R2515 B.n926 B.n925 71.676
R2516 B.n919 B.n187 71.676
R2517 B.n920 B.n919 71.676
R2518 B.n925 B.n924 71.676
R2519 B.n928 B.n927 71.676
R2520 B.n933 B.n932 71.676
R2521 B.n936 B.n935 71.676
R2522 B.n941 B.n940 71.676
R2523 B.n944 B.n943 71.676
R2524 B.n949 B.n948 71.676
R2525 B.n952 B.n951 71.676
R2526 B.n957 B.n956 71.676
R2527 B.n960 B.n959 71.676
R2528 B.n965 B.n964 71.676
R2529 B.n968 B.n967 71.676
R2530 B.n973 B.n972 71.676
R2531 B.n976 B.n975 71.676
R2532 B.n981 B.n980 71.676
R2533 B.n984 B.n983 71.676
R2534 B.n989 B.n988 71.676
R2535 B.n992 B.n991 71.676
R2536 B.n997 B.n996 71.676
R2537 B.n1000 B.n999 71.676
R2538 B.n1005 B.n1004 71.676
R2539 B.n1008 B.n1007 71.676
R2540 B.n1013 B.n1012 71.676
R2541 B.n1016 B.n1015 71.676
R2542 B.n1021 B.n1020 71.676
R2543 B.n1024 B.n1023 71.676
R2544 B.n1029 B.n1028 71.676
R2545 B.n1032 B.n1031 71.676
R2546 B.n1038 B.n1037 71.676
R2547 B.n1041 B.n1040 71.676
R2548 B.n1046 B.n1045 71.676
R2549 B.n1048 B.n153 71.676
R2550 B.n1053 B.n1052 71.676
R2551 B.n1058 B.n1057 71.676
R2552 B.n1061 B.n1060 71.676
R2553 B.n1066 B.n1065 71.676
R2554 B.n1069 B.n1068 71.676
R2555 B.n1074 B.n1073 71.676
R2556 B.n1077 B.n1076 71.676
R2557 B.n1082 B.n1081 71.676
R2558 B.n1085 B.n1084 71.676
R2559 B.n1090 B.n1089 71.676
R2560 B.n1093 B.n1092 71.676
R2561 B.n1098 B.n1097 71.676
R2562 B.n1101 B.n1100 71.676
R2563 B.n1106 B.n1105 71.676
R2564 B.n1109 B.n1108 71.676
R2565 B.n1114 B.n1113 71.676
R2566 B.n1117 B.n1116 71.676
R2567 B.n1122 B.n1121 71.676
R2568 B.n1125 B.n1124 71.676
R2569 B.n1130 B.n1129 71.676
R2570 B.n1133 B.n1132 71.676
R2571 B.n1138 B.n1137 71.676
R2572 B.n1141 B.n1140 71.676
R2573 B.n1146 B.n1145 71.676
R2574 B.n1149 B.n1148 71.676
R2575 B.n1154 B.n1153 71.676
R2576 B.n1157 B.n1156 71.676
R2577 B.n1162 B.n1161 71.676
R2578 B.n1165 B.n1164 71.676
R2579 B.n631 B.n630 71.676
R2580 B.n625 B.n320 71.676
R2581 B.n623 B.n622 71.676
R2582 B.n618 B.n617 71.676
R2583 B.n615 B.n614 71.676
R2584 B.n610 B.n609 71.676
R2585 B.n607 B.n606 71.676
R2586 B.n602 B.n601 71.676
R2587 B.n599 B.n598 71.676
R2588 B.n594 B.n593 71.676
R2589 B.n591 B.n590 71.676
R2590 B.n586 B.n585 71.676
R2591 B.n583 B.n582 71.676
R2592 B.n578 B.n577 71.676
R2593 B.n575 B.n574 71.676
R2594 B.n570 B.n569 71.676
R2595 B.n567 B.n566 71.676
R2596 B.n562 B.n561 71.676
R2597 B.n559 B.n558 71.676
R2598 B.n554 B.n553 71.676
R2599 B.n551 B.n550 71.676
R2600 B.n546 B.n545 71.676
R2601 B.n543 B.n542 71.676
R2602 B.n538 B.n537 71.676
R2603 B.n535 B.n534 71.676
R2604 B.n530 B.n529 71.676
R2605 B.n527 B.n526 71.676
R2606 B.n522 B.n521 71.676
R2607 B.n519 B.n518 71.676
R2608 B.n514 B.n513 71.676
R2609 B.n511 B.n510 71.676
R2610 B.n506 B.n505 71.676
R2611 B.n503 B.n502 71.676
R2612 B.n497 B.n496 71.676
R2613 B.n494 B.n493 71.676
R2614 B.n489 B.n488 71.676
R2615 B.n486 B.n485 71.676
R2616 B.n481 B.n480 71.676
R2617 B.n478 B.n477 71.676
R2618 B.n473 B.n472 71.676
R2619 B.n470 B.n469 71.676
R2620 B.n465 B.n464 71.676
R2621 B.n462 B.n461 71.676
R2622 B.n457 B.n456 71.676
R2623 B.n454 B.n453 71.676
R2624 B.n449 B.n448 71.676
R2625 B.n446 B.n445 71.676
R2626 B.n441 B.n440 71.676
R2627 B.n438 B.n437 71.676
R2628 B.n433 B.n432 71.676
R2629 B.n430 B.n429 71.676
R2630 B.n425 B.n424 71.676
R2631 B.n422 B.n421 71.676
R2632 B.n417 B.n416 71.676
R2633 B.n414 B.n413 71.676
R2634 B.n409 B.n408 71.676
R2635 B.n406 B.n405 71.676
R2636 B.n401 B.n400 71.676
R2637 B.n398 B.n397 71.676
R2638 B.n393 B.n392 71.676
R2639 B.n390 B.n389 71.676
R2640 B.n385 B.n316 71.676
R2641 B.n357 B.n356 63.4187
R2642 B.n350 B.n349 63.4187
R2643 B.n151 B.n150 63.4187
R2644 B.n159 B.n158 63.4187
R2645 B.n500 B.n357 59.5399
R2646 B.n351 B.n350 59.5399
R2647 B.n152 B.n151 59.5399
R2648 B.n1034 B.n159 59.5399
R2649 B.n636 B.n317 53.8721
R2650 B.n1170 B.n120 53.8721
R2651 B.n636 B.n313 33.0029
R2652 B.n642 B.n313 33.0029
R2653 B.n642 B.n309 33.0029
R2654 B.n648 B.n309 33.0029
R2655 B.n648 B.n305 33.0029
R2656 B.n654 B.n305 33.0029
R2657 B.n654 B.n301 33.0029
R2658 B.n660 B.n301 33.0029
R2659 B.n666 B.n297 33.0029
R2660 B.n666 B.n293 33.0029
R2661 B.n672 B.n293 33.0029
R2662 B.n672 B.n289 33.0029
R2663 B.n678 B.n289 33.0029
R2664 B.n678 B.n285 33.0029
R2665 B.n684 B.n285 33.0029
R2666 B.n684 B.n281 33.0029
R2667 B.n690 B.n281 33.0029
R2668 B.n690 B.n276 33.0029
R2669 B.n696 B.n276 33.0029
R2670 B.n696 B.n277 33.0029
R2671 B.n702 B.n269 33.0029
R2672 B.n708 B.n269 33.0029
R2673 B.n708 B.n265 33.0029
R2674 B.n714 B.n265 33.0029
R2675 B.n714 B.n261 33.0029
R2676 B.n720 B.n261 33.0029
R2677 B.n720 B.n257 33.0029
R2678 B.n726 B.n257 33.0029
R2679 B.n732 B.n253 33.0029
R2680 B.n732 B.n249 33.0029
R2681 B.n738 B.n249 33.0029
R2682 B.n738 B.n245 33.0029
R2683 B.n744 B.n245 33.0029
R2684 B.n744 B.n241 33.0029
R2685 B.n750 B.n241 33.0029
R2686 B.n750 B.n237 33.0029
R2687 B.n756 B.n237 33.0029
R2688 B.n762 B.n233 33.0029
R2689 B.n762 B.n229 33.0029
R2690 B.n768 B.n229 33.0029
R2691 B.n768 B.n225 33.0029
R2692 B.n774 B.n225 33.0029
R2693 B.n774 B.n220 33.0029
R2694 B.n780 B.n220 33.0029
R2695 B.n780 B.n221 33.0029
R2696 B.n786 B.n213 33.0029
R2697 B.n792 B.n213 33.0029
R2698 B.n792 B.n209 33.0029
R2699 B.n798 B.n209 33.0029
R2700 B.n798 B.n205 33.0029
R2701 B.n804 B.n205 33.0029
R2702 B.n804 B.n201 33.0029
R2703 B.n811 B.n201 33.0029
R2704 B.n811 B.n810 33.0029
R2705 B.n817 B.n194 33.0029
R2706 B.n824 B.n194 33.0029
R2707 B.n824 B.n190 33.0029
R2708 B.n830 B.n190 33.0029
R2709 B.n830 B.n4 33.0029
R2710 B.n1300 B.n4 33.0029
R2711 B.n1300 B.n1299 33.0029
R2712 B.n1299 B.n1298 33.0029
R2713 B.n1298 B.n8 33.0029
R2714 B.n1292 B.n8 33.0029
R2715 B.n1292 B.n1291 33.0029
R2716 B.n1291 B.n1290 33.0029
R2717 B.n1284 B.n18 33.0029
R2718 B.n1284 B.n1283 33.0029
R2719 B.n1283 B.n1282 33.0029
R2720 B.n1282 B.n22 33.0029
R2721 B.n1276 B.n22 33.0029
R2722 B.n1276 B.n1275 33.0029
R2723 B.n1275 B.n1274 33.0029
R2724 B.n1274 B.n29 33.0029
R2725 B.n1268 B.n29 33.0029
R2726 B.n1267 B.n1266 33.0029
R2727 B.n1266 B.n36 33.0029
R2728 B.n1260 B.n36 33.0029
R2729 B.n1260 B.n1259 33.0029
R2730 B.n1259 B.n1258 33.0029
R2731 B.n1258 B.n43 33.0029
R2732 B.n1252 B.n43 33.0029
R2733 B.n1252 B.n1251 33.0029
R2734 B.n1250 B.n50 33.0029
R2735 B.n1244 B.n50 33.0029
R2736 B.n1244 B.n1243 33.0029
R2737 B.n1243 B.n1242 33.0029
R2738 B.n1242 B.n57 33.0029
R2739 B.n1236 B.n57 33.0029
R2740 B.n1236 B.n1235 33.0029
R2741 B.n1235 B.n1234 33.0029
R2742 B.n1234 B.n64 33.0029
R2743 B.n1228 B.n1227 33.0029
R2744 B.n1227 B.n1226 33.0029
R2745 B.n1226 B.n71 33.0029
R2746 B.n1220 B.n71 33.0029
R2747 B.n1220 B.n1219 33.0029
R2748 B.n1219 B.n1218 33.0029
R2749 B.n1218 B.n78 33.0029
R2750 B.n1212 B.n78 33.0029
R2751 B.n1211 B.n1210 33.0029
R2752 B.n1210 B.n85 33.0029
R2753 B.n1204 B.n85 33.0029
R2754 B.n1204 B.n1203 33.0029
R2755 B.n1203 B.n1202 33.0029
R2756 B.n1202 B.n92 33.0029
R2757 B.n1196 B.n92 33.0029
R2758 B.n1196 B.n1195 33.0029
R2759 B.n1195 B.n1194 33.0029
R2760 B.n1194 B.n99 33.0029
R2761 B.n1188 B.n99 33.0029
R2762 B.n1188 B.n1187 33.0029
R2763 B.n1186 B.n106 33.0029
R2764 B.n1180 B.n106 33.0029
R2765 B.n1180 B.n1179 33.0029
R2766 B.n1179 B.n1178 33.0029
R2767 B.n1178 B.n113 33.0029
R2768 B.n1172 B.n113 33.0029
R2769 B.n1172 B.n1171 33.0029
R2770 B.n1171 B.n1170 33.0029
R2771 B.n221 B.t23 32.0323
R2772 B.t1 B.n1267 32.0323
R2773 B.n702 B.t7 29.1203
R2774 B.n1212 B.t5 29.1203
R2775 B.n1168 B.n1167 27.942
R2776 B.n917 B.n916 27.942
R2777 B.n638 B.n315 27.942
R2778 B.n634 B.n633 27.942
R2779 B.n726 B.t2 24.267
R2780 B.n1228 B.t0 24.267
R2781 B.t10 B.n297 23.2963
R2782 B.n1187 B.t17 23.2963
R2783 B.t4 B.n233 21.355
R2784 B.n1251 B.t6 21.355
R2785 B.n810 B.t3 19.4137
R2786 B.n18 B.t8 19.4137
R2787 B B.n1302 18.0485
R2788 B.n817 B.t3 13.5897
R2789 B.n1290 B.t8 13.5897
R2790 B.n756 B.t4 11.6484
R2791 B.t6 B.n1250 11.6484
R2792 B.n1167 B.n1166 10.6151
R2793 B.n1166 B.n122 10.6151
R2794 B.n1160 B.n122 10.6151
R2795 B.n1160 B.n1159 10.6151
R2796 B.n1159 B.n1158 10.6151
R2797 B.n1158 B.n124 10.6151
R2798 B.n1152 B.n124 10.6151
R2799 B.n1152 B.n1151 10.6151
R2800 B.n1151 B.n1150 10.6151
R2801 B.n1150 B.n126 10.6151
R2802 B.n1144 B.n126 10.6151
R2803 B.n1144 B.n1143 10.6151
R2804 B.n1143 B.n1142 10.6151
R2805 B.n1142 B.n128 10.6151
R2806 B.n1136 B.n128 10.6151
R2807 B.n1136 B.n1135 10.6151
R2808 B.n1135 B.n1134 10.6151
R2809 B.n1134 B.n130 10.6151
R2810 B.n1128 B.n130 10.6151
R2811 B.n1128 B.n1127 10.6151
R2812 B.n1127 B.n1126 10.6151
R2813 B.n1126 B.n132 10.6151
R2814 B.n1120 B.n132 10.6151
R2815 B.n1120 B.n1119 10.6151
R2816 B.n1119 B.n1118 10.6151
R2817 B.n1118 B.n134 10.6151
R2818 B.n1112 B.n134 10.6151
R2819 B.n1112 B.n1111 10.6151
R2820 B.n1111 B.n1110 10.6151
R2821 B.n1110 B.n136 10.6151
R2822 B.n1104 B.n136 10.6151
R2823 B.n1104 B.n1103 10.6151
R2824 B.n1103 B.n1102 10.6151
R2825 B.n1102 B.n138 10.6151
R2826 B.n1096 B.n138 10.6151
R2827 B.n1096 B.n1095 10.6151
R2828 B.n1095 B.n1094 10.6151
R2829 B.n1094 B.n140 10.6151
R2830 B.n1088 B.n140 10.6151
R2831 B.n1088 B.n1087 10.6151
R2832 B.n1087 B.n1086 10.6151
R2833 B.n1086 B.n142 10.6151
R2834 B.n1080 B.n142 10.6151
R2835 B.n1080 B.n1079 10.6151
R2836 B.n1079 B.n1078 10.6151
R2837 B.n1078 B.n144 10.6151
R2838 B.n1072 B.n144 10.6151
R2839 B.n1072 B.n1071 10.6151
R2840 B.n1071 B.n1070 10.6151
R2841 B.n1070 B.n146 10.6151
R2842 B.n1064 B.n146 10.6151
R2843 B.n1064 B.n1063 10.6151
R2844 B.n1063 B.n1062 10.6151
R2845 B.n1062 B.n148 10.6151
R2846 B.n1056 B.n148 10.6151
R2847 B.n1056 B.n1055 10.6151
R2848 B.n1055 B.n1054 10.6151
R2849 B.n1050 B.n1049 10.6151
R2850 B.n1049 B.n154 10.6151
R2851 B.n1044 B.n154 10.6151
R2852 B.n1044 B.n1043 10.6151
R2853 B.n1043 B.n1042 10.6151
R2854 B.n1042 B.n156 10.6151
R2855 B.n1036 B.n156 10.6151
R2856 B.n1036 B.n1035 10.6151
R2857 B.n1033 B.n160 10.6151
R2858 B.n1027 B.n160 10.6151
R2859 B.n1027 B.n1026 10.6151
R2860 B.n1026 B.n1025 10.6151
R2861 B.n1025 B.n162 10.6151
R2862 B.n1019 B.n162 10.6151
R2863 B.n1019 B.n1018 10.6151
R2864 B.n1018 B.n1017 10.6151
R2865 B.n1017 B.n164 10.6151
R2866 B.n1011 B.n164 10.6151
R2867 B.n1011 B.n1010 10.6151
R2868 B.n1010 B.n1009 10.6151
R2869 B.n1009 B.n166 10.6151
R2870 B.n1003 B.n166 10.6151
R2871 B.n1003 B.n1002 10.6151
R2872 B.n1002 B.n1001 10.6151
R2873 B.n1001 B.n168 10.6151
R2874 B.n995 B.n168 10.6151
R2875 B.n995 B.n994 10.6151
R2876 B.n994 B.n993 10.6151
R2877 B.n993 B.n170 10.6151
R2878 B.n987 B.n170 10.6151
R2879 B.n987 B.n986 10.6151
R2880 B.n986 B.n985 10.6151
R2881 B.n985 B.n172 10.6151
R2882 B.n979 B.n172 10.6151
R2883 B.n979 B.n978 10.6151
R2884 B.n978 B.n977 10.6151
R2885 B.n977 B.n174 10.6151
R2886 B.n971 B.n174 10.6151
R2887 B.n971 B.n970 10.6151
R2888 B.n970 B.n969 10.6151
R2889 B.n969 B.n176 10.6151
R2890 B.n963 B.n176 10.6151
R2891 B.n963 B.n962 10.6151
R2892 B.n962 B.n961 10.6151
R2893 B.n961 B.n178 10.6151
R2894 B.n955 B.n178 10.6151
R2895 B.n955 B.n954 10.6151
R2896 B.n954 B.n953 10.6151
R2897 B.n953 B.n180 10.6151
R2898 B.n947 B.n180 10.6151
R2899 B.n947 B.n946 10.6151
R2900 B.n946 B.n945 10.6151
R2901 B.n945 B.n182 10.6151
R2902 B.n939 B.n182 10.6151
R2903 B.n939 B.n938 10.6151
R2904 B.n938 B.n937 10.6151
R2905 B.n937 B.n184 10.6151
R2906 B.n931 B.n184 10.6151
R2907 B.n931 B.n930 10.6151
R2908 B.n930 B.n929 10.6151
R2909 B.n929 B.n186 10.6151
R2910 B.n923 B.n186 10.6151
R2911 B.n923 B.n922 10.6151
R2912 B.n922 B.n921 10.6151
R2913 B.n921 B.n917 10.6151
R2914 B.n639 B.n638 10.6151
R2915 B.n640 B.n639 10.6151
R2916 B.n640 B.n307 10.6151
R2917 B.n650 B.n307 10.6151
R2918 B.n651 B.n650 10.6151
R2919 B.n652 B.n651 10.6151
R2920 B.n652 B.n299 10.6151
R2921 B.n662 B.n299 10.6151
R2922 B.n663 B.n662 10.6151
R2923 B.n664 B.n663 10.6151
R2924 B.n664 B.n291 10.6151
R2925 B.n674 B.n291 10.6151
R2926 B.n675 B.n674 10.6151
R2927 B.n676 B.n675 10.6151
R2928 B.n676 B.n283 10.6151
R2929 B.n686 B.n283 10.6151
R2930 B.n687 B.n686 10.6151
R2931 B.n688 B.n687 10.6151
R2932 B.n688 B.n274 10.6151
R2933 B.n698 B.n274 10.6151
R2934 B.n699 B.n698 10.6151
R2935 B.n700 B.n699 10.6151
R2936 B.n700 B.n267 10.6151
R2937 B.n710 B.n267 10.6151
R2938 B.n711 B.n710 10.6151
R2939 B.n712 B.n711 10.6151
R2940 B.n712 B.n259 10.6151
R2941 B.n722 B.n259 10.6151
R2942 B.n723 B.n722 10.6151
R2943 B.n724 B.n723 10.6151
R2944 B.n724 B.n251 10.6151
R2945 B.n734 B.n251 10.6151
R2946 B.n735 B.n734 10.6151
R2947 B.n736 B.n735 10.6151
R2948 B.n736 B.n243 10.6151
R2949 B.n746 B.n243 10.6151
R2950 B.n747 B.n746 10.6151
R2951 B.n748 B.n747 10.6151
R2952 B.n748 B.n235 10.6151
R2953 B.n758 B.n235 10.6151
R2954 B.n759 B.n758 10.6151
R2955 B.n760 B.n759 10.6151
R2956 B.n760 B.n227 10.6151
R2957 B.n770 B.n227 10.6151
R2958 B.n771 B.n770 10.6151
R2959 B.n772 B.n771 10.6151
R2960 B.n772 B.n218 10.6151
R2961 B.n782 B.n218 10.6151
R2962 B.n783 B.n782 10.6151
R2963 B.n784 B.n783 10.6151
R2964 B.n784 B.n211 10.6151
R2965 B.n794 B.n211 10.6151
R2966 B.n795 B.n794 10.6151
R2967 B.n796 B.n795 10.6151
R2968 B.n796 B.n203 10.6151
R2969 B.n806 B.n203 10.6151
R2970 B.n807 B.n806 10.6151
R2971 B.n808 B.n807 10.6151
R2972 B.n808 B.n196 10.6151
R2973 B.n819 B.n196 10.6151
R2974 B.n820 B.n819 10.6151
R2975 B.n822 B.n820 10.6151
R2976 B.n822 B.n821 10.6151
R2977 B.n821 B.n188 10.6151
R2978 B.n833 B.n188 10.6151
R2979 B.n834 B.n833 10.6151
R2980 B.n835 B.n834 10.6151
R2981 B.n836 B.n835 10.6151
R2982 B.n838 B.n836 10.6151
R2983 B.n839 B.n838 10.6151
R2984 B.n840 B.n839 10.6151
R2985 B.n841 B.n840 10.6151
R2986 B.n843 B.n841 10.6151
R2987 B.n844 B.n843 10.6151
R2988 B.n845 B.n844 10.6151
R2989 B.n846 B.n845 10.6151
R2990 B.n848 B.n846 10.6151
R2991 B.n849 B.n848 10.6151
R2992 B.n850 B.n849 10.6151
R2993 B.n851 B.n850 10.6151
R2994 B.n853 B.n851 10.6151
R2995 B.n854 B.n853 10.6151
R2996 B.n855 B.n854 10.6151
R2997 B.n856 B.n855 10.6151
R2998 B.n858 B.n856 10.6151
R2999 B.n859 B.n858 10.6151
R3000 B.n860 B.n859 10.6151
R3001 B.n861 B.n860 10.6151
R3002 B.n863 B.n861 10.6151
R3003 B.n864 B.n863 10.6151
R3004 B.n865 B.n864 10.6151
R3005 B.n866 B.n865 10.6151
R3006 B.n868 B.n866 10.6151
R3007 B.n869 B.n868 10.6151
R3008 B.n870 B.n869 10.6151
R3009 B.n871 B.n870 10.6151
R3010 B.n873 B.n871 10.6151
R3011 B.n874 B.n873 10.6151
R3012 B.n875 B.n874 10.6151
R3013 B.n876 B.n875 10.6151
R3014 B.n878 B.n876 10.6151
R3015 B.n879 B.n878 10.6151
R3016 B.n880 B.n879 10.6151
R3017 B.n881 B.n880 10.6151
R3018 B.n883 B.n881 10.6151
R3019 B.n884 B.n883 10.6151
R3020 B.n885 B.n884 10.6151
R3021 B.n886 B.n885 10.6151
R3022 B.n888 B.n886 10.6151
R3023 B.n889 B.n888 10.6151
R3024 B.n890 B.n889 10.6151
R3025 B.n891 B.n890 10.6151
R3026 B.n893 B.n891 10.6151
R3027 B.n894 B.n893 10.6151
R3028 B.n895 B.n894 10.6151
R3029 B.n896 B.n895 10.6151
R3030 B.n898 B.n896 10.6151
R3031 B.n899 B.n898 10.6151
R3032 B.n900 B.n899 10.6151
R3033 B.n901 B.n900 10.6151
R3034 B.n903 B.n901 10.6151
R3035 B.n904 B.n903 10.6151
R3036 B.n905 B.n904 10.6151
R3037 B.n906 B.n905 10.6151
R3038 B.n908 B.n906 10.6151
R3039 B.n909 B.n908 10.6151
R3040 B.n910 B.n909 10.6151
R3041 B.n911 B.n910 10.6151
R3042 B.n913 B.n911 10.6151
R3043 B.n914 B.n913 10.6151
R3044 B.n915 B.n914 10.6151
R3045 B.n916 B.n915 10.6151
R3046 B.n633 B.n632 10.6151
R3047 B.n632 B.n319 10.6151
R3048 B.n627 B.n319 10.6151
R3049 B.n627 B.n626 10.6151
R3050 B.n626 B.n321 10.6151
R3051 B.n621 B.n321 10.6151
R3052 B.n621 B.n620 10.6151
R3053 B.n620 B.n619 10.6151
R3054 B.n619 B.n323 10.6151
R3055 B.n613 B.n323 10.6151
R3056 B.n613 B.n612 10.6151
R3057 B.n612 B.n611 10.6151
R3058 B.n611 B.n325 10.6151
R3059 B.n605 B.n325 10.6151
R3060 B.n605 B.n604 10.6151
R3061 B.n604 B.n603 10.6151
R3062 B.n603 B.n327 10.6151
R3063 B.n597 B.n327 10.6151
R3064 B.n597 B.n596 10.6151
R3065 B.n596 B.n595 10.6151
R3066 B.n595 B.n329 10.6151
R3067 B.n589 B.n329 10.6151
R3068 B.n589 B.n588 10.6151
R3069 B.n588 B.n587 10.6151
R3070 B.n587 B.n331 10.6151
R3071 B.n581 B.n331 10.6151
R3072 B.n581 B.n580 10.6151
R3073 B.n580 B.n579 10.6151
R3074 B.n579 B.n333 10.6151
R3075 B.n573 B.n333 10.6151
R3076 B.n573 B.n572 10.6151
R3077 B.n572 B.n571 10.6151
R3078 B.n571 B.n335 10.6151
R3079 B.n565 B.n335 10.6151
R3080 B.n565 B.n564 10.6151
R3081 B.n564 B.n563 10.6151
R3082 B.n563 B.n337 10.6151
R3083 B.n557 B.n337 10.6151
R3084 B.n557 B.n556 10.6151
R3085 B.n556 B.n555 10.6151
R3086 B.n555 B.n339 10.6151
R3087 B.n549 B.n339 10.6151
R3088 B.n549 B.n548 10.6151
R3089 B.n548 B.n547 10.6151
R3090 B.n547 B.n341 10.6151
R3091 B.n541 B.n341 10.6151
R3092 B.n541 B.n540 10.6151
R3093 B.n540 B.n539 10.6151
R3094 B.n539 B.n343 10.6151
R3095 B.n533 B.n343 10.6151
R3096 B.n533 B.n532 10.6151
R3097 B.n532 B.n531 10.6151
R3098 B.n531 B.n345 10.6151
R3099 B.n525 B.n345 10.6151
R3100 B.n525 B.n524 10.6151
R3101 B.n524 B.n523 10.6151
R3102 B.n523 B.n347 10.6151
R3103 B.n517 B.n516 10.6151
R3104 B.n516 B.n515 10.6151
R3105 B.n515 B.n352 10.6151
R3106 B.n509 B.n352 10.6151
R3107 B.n509 B.n508 10.6151
R3108 B.n508 B.n507 10.6151
R3109 B.n507 B.n354 10.6151
R3110 B.n501 B.n354 10.6151
R3111 B.n499 B.n498 10.6151
R3112 B.n498 B.n358 10.6151
R3113 B.n492 B.n358 10.6151
R3114 B.n492 B.n491 10.6151
R3115 B.n491 B.n490 10.6151
R3116 B.n490 B.n360 10.6151
R3117 B.n484 B.n360 10.6151
R3118 B.n484 B.n483 10.6151
R3119 B.n483 B.n482 10.6151
R3120 B.n482 B.n362 10.6151
R3121 B.n476 B.n362 10.6151
R3122 B.n476 B.n475 10.6151
R3123 B.n475 B.n474 10.6151
R3124 B.n474 B.n364 10.6151
R3125 B.n468 B.n364 10.6151
R3126 B.n468 B.n467 10.6151
R3127 B.n467 B.n466 10.6151
R3128 B.n466 B.n366 10.6151
R3129 B.n460 B.n366 10.6151
R3130 B.n460 B.n459 10.6151
R3131 B.n459 B.n458 10.6151
R3132 B.n458 B.n368 10.6151
R3133 B.n452 B.n368 10.6151
R3134 B.n452 B.n451 10.6151
R3135 B.n451 B.n450 10.6151
R3136 B.n450 B.n370 10.6151
R3137 B.n444 B.n370 10.6151
R3138 B.n444 B.n443 10.6151
R3139 B.n443 B.n442 10.6151
R3140 B.n442 B.n372 10.6151
R3141 B.n436 B.n372 10.6151
R3142 B.n436 B.n435 10.6151
R3143 B.n435 B.n434 10.6151
R3144 B.n434 B.n374 10.6151
R3145 B.n428 B.n374 10.6151
R3146 B.n428 B.n427 10.6151
R3147 B.n427 B.n426 10.6151
R3148 B.n426 B.n376 10.6151
R3149 B.n420 B.n376 10.6151
R3150 B.n420 B.n419 10.6151
R3151 B.n419 B.n418 10.6151
R3152 B.n418 B.n378 10.6151
R3153 B.n412 B.n378 10.6151
R3154 B.n412 B.n411 10.6151
R3155 B.n411 B.n410 10.6151
R3156 B.n410 B.n380 10.6151
R3157 B.n404 B.n380 10.6151
R3158 B.n404 B.n403 10.6151
R3159 B.n403 B.n402 10.6151
R3160 B.n402 B.n382 10.6151
R3161 B.n396 B.n382 10.6151
R3162 B.n396 B.n395 10.6151
R3163 B.n395 B.n394 10.6151
R3164 B.n394 B.n384 10.6151
R3165 B.n388 B.n384 10.6151
R3166 B.n388 B.n387 10.6151
R3167 B.n387 B.n315 10.6151
R3168 B.n634 B.n311 10.6151
R3169 B.n644 B.n311 10.6151
R3170 B.n645 B.n644 10.6151
R3171 B.n646 B.n645 10.6151
R3172 B.n646 B.n303 10.6151
R3173 B.n656 B.n303 10.6151
R3174 B.n657 B.n656 10.6151
R3175 B.n658 B.n657 10.6151
R3176 B.n658 B.n295 10.6151
R3177 B.n668 B.n295 10.6151
R3178 B.n669 B.n668 10.6151
R3179 B.n670 B.n669 10.6151
R3180 B.n670 B.n287 10.6151
R3181 B.n680 B.n287 10.6151
R3182 B.n681 B.n680 10.6151
R3183 B.n682 B.n681 10.6151
R3184 B.n682 B.n279 10.6151
R3185 B.n692 B.n279 10.6151
R3186 B.n693 B.n692 10.6151
R3187 B.n694 B.n693 10.6151
R3188 B.n694 B.n271 10.6151
R3189 B.n704 B.n271 10.6151
R3190 B.n705 B.n704 10.6151
R3191 B.n706 B.n705 10.6151
R3192 B.n706 B.n263 10.6151
R3193 B.n716 B.n263 10.6151
R3194 B.n717 B.n716 10.6151
R3195 B.n718 B.n717 10.6151
R3196 B.n718 B.n255 10.6151
R3197 B.n728 B.n255 10.6151
R3198 B.n729 B.n728 10.6151
R3199 B.n730 B.n729 10.6151
R3200 B.n730 B.n247 10.6151
R3201 B.n740 B.n247 10.6151
R3202 B.n741 B.n740 10.6151
R3203 B.n742 B.n741 10.6151
R3204 B.n742 B.n239 10.6151
R3205 B.n752 B.n239 10.6151
R3206 B.n753 B.n752 10.6151
R3207 B.n754 B.n753 10.6151
R3208 B.n754 B.n231 10.6151
R3209 B.n764 B.n231 10.6151
R3210 B.n765 B.n764 10.6151
R3211 B.n766 B.n765 10.6151
R3212 B.n766 B.n223 10.6151
R3213 B.n776 B.n223 10.6151
R3214 B.n777 B.n776 10.6151
R3215 B.n778 B.n777 10.6151
R3216 B.n778 B.n215 10.6151
R3217 B.n788 B.n215 10.6151
R3218 B.n789 B.n788 10.6151
R3219 B.n790 B.n789 10.6151
R3220 B.n790 B.n207 10.6151
R3221 B.n800 B.n207 10.6151
R3222 B.n801 B.n800 10.6151
R3223 B.n802 B.n801 10.6151
R3224 B.n802 B.n199 10.6151
R3225 B.n813 B.n199 10.6151
R3226 B.n814 B.n813 10.6151
R3227 B.n815 B.n814 10.6151
R3228 B.n815 B.n192 10.6151
R3229 B.n826 B.n192 10.6151
R3230 B.n827 B.n826 10.6151
R3231 B.n828 B.n827 10.6151
R3232 B.n828 B.n0 10.6151
R3233 B.n1296 B.n1 10.6151
R3234 B.n1296 B.n1295 10.6151
R3235 B.n1295 B.n1294 10.6151
R3236 B.n1294 B.n10 10.6151
R3237 B.n1288 B.n10 10.6151
R3238 B.n1288 B.n1287 10.6151
R3239 B.n1287 B.n1286 10.6151
R3240 B.n1286 B.n16 10.6151
R3241 B.n1280 B.n16 10.6151
R3242 B.n1280 B.n1279 10.6151
R3243 B.n1279 B.n1278 10.6151
R3244 B.n1278 B.n24 10.6151
R3245 B.n1272 B.n24 10.6151
R3246 B.n1272 B.n1271 10.6151
R3247 B.n1271 B.n1270 10.6151
R3248 B.n1270 B.n31 10.6151
R3249 B.n1264 B.n31 10.6151
R3250 B.n1264 B.n1263 10.6151
R3251 B.n1263 B.n1262 10.6151
R3252 B.n1262 B.n38 10.6151
R3253 B.n1256 B.n38 10.6151
R3254 B.n1256 B.n1255 10.6151
R3255 B.n1255 B.n1254 10.6151
R3256 B.n1254 B.n45 10.6151
R3257 B.n1248 B.n45 10.6151
R3258 B.n1248 B.n1247 10.6151
R3259 B.n1247 B.n1246 10.6151
R3260 B.n1246 B.n52 10.6151
R3261 B.n1240 B.n52 10.6151
R3262 B.n1240 B.n1239 10.6151
R3263 B.n1239 B.n1238 10.6151
R3264 B.n1238 B.n59 10.6151
R3265 B.n1232 B.n59 10.6151
R3266 B.n1232 B.n1231 10.6151
R3267 B.n1231 B.n1230 10.6151
R3268 B.n1230 B.n66 10.6151
R3269 B.n1224 B.n66 10.6151
R3270 B.n1224 B.n1223 10.6151
R3271 B.n1223 B.n1222 10.6151
R3272 B.n1222 B.n73 10.6151
R3273 B.n1216 B.n73 10.6151
R3274 B.n1216 B.n1215 10.6151
R3275 B.n1215 B.n1214 10.6151
R3276 B.n1214 B.n80 10.6151
R3277 B.n1208 B.n80 10.6151
R3278 B.n1208 B.n1207 10.6151
R3279 B.n1207 B.n1206 10.6151
R3280 B.n1206 B.n87 10.6151
R3281 B.n1200 B.n87 10.6151
R3282 B.n1200 B.n1199 10.6151
R3283 B.n1199 B.n1198 10.6151
R3284 B.n1198 B.n94 10.6151
R3285 B.n1192 B.n94 10.6151
R3286 B.n1192 B.n1191 10.6151
R3287 B.n1191 B.n1190 10.6151
R3288 B.n1190 B.n101 10.6151
R3289 B.n1184 B.n101 10.6151
R3290 B.n1184 B.n1183 10.6151
R3291 B.n1183 B.n1182 10.6151
R3292 B.n1182 B.n108 10.6151
R3293 B.n1176 B.n108 10.6151
R3294 B.n1176 B.n1175 10.6151
R3295 B.n1175 B.n1174 10.6151
R3296 B.n1174 B.n115 10.6151
R3297 B.n1168 B.n115 10.6151
R3298 B.n660 B.t10 9.7071
R3299 B.t17 B.n1186 9.7071
R3300 B.t2 B.n253 8.73644
R3301 B.t0 B.n64 8.73644
R3302 B.n1050 B.n152 6.5566
R3303 B.n1035 B.n1034 6.5566
R3304 B.n517 B.n351 6.5566
R3305 B.n501 B.n500 6.5566
R3306 B.n1054 B.n152 4.05904
R3307 B.n1034 B.n1033 4.05904
R3308 B.n351 B.n347 4.05904
R3309 B.n500 B.n499 4.05904
R3310 B.n277 B.t7 3.88314
R3311 B.t5 B.n1211 3.88314
R3312 B.n1302 B.n0 2.81026
R3313 B.n1302 B.n1 2.81026
R3314 B.n786 B.t23 0.97116
R3315 B.n1268 B.t1 0.97116
R3316 VN.n10 VN.t4 175.234
R3317 VN.n56 VN.t8 175.234
R3318 VN.n87 VN.n45 161.3
R3319 VN.n86 VN.n85 161.3
R3320 VN.n84 VN.n46 161.3
R3321 VN.n83 VN.n82 161.3
R3322 VN.n81 VN.n47 161.3
R3323 VN.n80 VN.n79 161.3
R3324 VN.n78 VN.n48 161.3
R3325 VN.n77 VN.n76 161.3
R3326 VN.n75 VN.n49 161.3
R3327 VN.n74 VN.n73 161.3
R3328 VN.n72 VN.n51 161.3
R3329 VN.n71 VN.n70 161.3
R3330 VN.n69 VN.n52 161.3
R3331 VN.n68 VN.n67 161.3
R3332 VN.n66 VN.n53 161.3
R3333 VN.n65 VN.n64 161.3
R3334 VN.n63 VN.n54 161.3
R3335 VN.n62 VN.n61 161.3
R3336 VN.n60 VN.n55 161.3
R3337 VN.n59 VN.n58 161.3
R3338 VN.n42 VN.n0 161.3
R3339 VN.n41 VN.n40 161.3
R3340 VN.n39 VN.n1 161.3
R3341 VN.n38 VN.n37 161.3
R3342 VN.n36 VN.n2 161.3
R3343 VN.n35 VN.n34 161.3
R3344 VN.n33 VN.n3 161.3
R3345 VN.n32 VN.n31 161.3
R3346 VN.n29 VN.n4 161.3
R3347 VN.n28 VN.n27 161.3
R3348 VN.n26 VN.n5 161.3
R3349 VN.n25 VN.n24 161.3
R3350 VN.n23 VN.n6 161.3
R3351 VN.n22 VN.n21 161.3
R3352 VN.n20 VN.n7 161.3
R3353 VN.n19 VN.n18 161.3
R3354 VN.n17 VN.n8 161.3
R3355 VN.n16 VN.n15 161.3
R3356 VN.n14 VN.n9 161.3
R3357 VN.n13 VN.n12 161.3
R3358 VN.n22 VN.t5 142.552
R3359 VN.n11 VN.t0 142.552
R3360 VN.n30 VN.t1 142.552
R3361 VN.n43 VN.t6 142.552
R3362 VN.n68 VN.t2 142.552
R3363 VN.n57 VN.t3 142.552
R3364 VN.n50 VN.t9 142.552
R3365 VN.n88 VN.t7 142.552
R3366 VN.n44 VN.n43 108.799
R3367 VN.n89 VN.n88 108.799
R3368 VN.n11 VN.n10 60.6237
R3369 VN.n57 VN.n56 60.6237
R3370 VN VN.n89 59.305
R3371 VN.n17 VN.n16 53.6055
R3372 VN.n28 VN.n5 53.6055
R3373 VN.n63 VN.n62 53.6055
R3374 VN.n74 VN.n51 53.6055
R3375 VN.n37 VN.n36 49.7204
R3376 VN.n82 VN.n81 49.7204
R3377 VN.n37 VN.n1 31.2664
R3378 VN.n82 VN.n46 31.2664
R3379 VN.n18 VN.n17 27.3813
R3380 VN.n24 VN.n5 27.3813
R3381 VN.n64 VN.n63 27.3813
R3382 VN.n70 VN.n51 27.3813
R3383 VN.n12 VN.n9 24.4675
R3384 VN.n16 VN.n9 24.4675
R3385 VN.n18 VN.n7 24.4675
R3386 VN.n22 VN.n7 24.4675
R3387 VN.n23 VN.n22 24.4675
R3388 VN.n24 VN.n23 24.4675
R3389 VN.n29 VN.n28 24.4675
R3390 VN.n31 VN.n29 24.4675
R3391 VN.n35 VN.n3 24.4675
R3392 VN.n36 VN.n35 24.4675
R3393 VN.n41 VN.n1 24.4675
R3394 VN.n42 VN.n41 24.4675
R3395 VN.n62 VN.n55 24.4675
R3396 VN.n58 VN.n55 24.4675
R3397 VN.n70 VN.n69 24.4675
R3398 VN.n69 VN.n68 24.4675
R3399 VN.n68 VN.n53 24.4675
R3400 VN.n64 VN.n53 24.4675
R3401 VN.n81 VN.n80 24.4675
R3402 VN.n80 VN.n48 24.4675
R3403 VN.n76 VN.n75 24.4675
R3404 VN.n75 VN.n74 24.4675
R3405 VN.n87 VN.n86 24.4675
R3406 VN.n86 VN.n46 24.4675
R3407 VN.n12 VN.n11 13.2127
R3408 VN.n31 VN.n30 13.2127
R3409 VN.n58 VN.n57 13.2127
R3410 VN.n76 VN.n50 13.2127
R3411 VN.n30 VN.n3 11.2553
R3412 VN.n50 VN.n48 11.2553
R3413 VN.n59 VN.n56 5.12434
R3414 VN.n13 VN.n10 5.12434
R3415 VN.n43 VN.n42 1.95786
R3416 VN.n88 VN.n87 1.95786
R3417 VN.n89 VN.n45 0.278367
R3418 VN.n44 VN.n0 0.278367
R3419 VN.n85 VN.n45 0.189894
R3420 VN.n85 VN.n84 0.189894
R3421 VN.n84 VN.n83 0.189894
R3422 VN.n83 VN.n47 0.189894
R3423 VN.n79 VN.n47 0.189894
R3424 VN.n79 VN.n78 0.189894
R3425 VN.n78 VN.n77 0.189894
R3426 VN.n77 VN.n49 0.189894
R3427 VN.n73 VN.n49 0.189894
R3428 VN.n73 VN.n72 0.189894
R3429 VN.n72 VN.n71 0.189894
R3430 VN.n71 VN.n52 0.189894
R3431 VN.n67 VN.n52 0.189894
R3432 VN.n67 VN.n66 0.189894
R3433 VN.n66 VN.n65 0.189894
R3434 VN.n65 VN.n54 0.189894
R3435 VN.n61 VN.n54 0.189894
R3436 VN.n61 VN.n60 0.189894
R3437 VN.n60 VN.n59 0.189894
R3438 VN.n14 VN.n13 0.189894
R3439 VN.n15 VN.n14 0.189894
R3440 VN.n15 VN.n8 0.189894
R3441 VN.n19 VN.n8 0.189894
R3442 VN.n20 VN.n19 0.189894
R3443 VN.n21 VN.n20 0.189894
R3444 VN.n21 VN.n6 0.189894
R3445 VN.n25 VN.n6 0.189894
R3446 VN.n26 VN.n25 0.189894
R3447 VN.n27 VN.n26 0.189894
R3448 VN.n27 VN.n4 0.189894
R3449 VN.n32 VN.n4 0.189894
R3450 VN.n33 VN.n32 0.189894
R3451 VN.n34 VN.n33 0.189894
R3452 VN.n34 VN.n2 0.189894
R3453 VN.n38 VN.n2 0.189894
R3454 VN.n39 VN.n38 0.189894
R3455 VN.n40 VN.n39 0.189894
R3456 VN.n40 VN.n0 0.189894
R3457 VN VN.n44 0.153454
R3458 VDD2.n193 VDD2.n192 289.615
R3459 VDD2.n94 VDD2.n93 289.615
R3460 VDD2.n192 VDD2.n191 185
R3461 VDD2.n101 VDD2.n100 185
R3462 VDD2.n186 VDD2.n185 185
R3463 VDD2.n184 VDD2.n183 185
R3464 VDD2.n105 VDD2.n104 185
R3465 VDD2.n178 VDD2.n177 185
R3466 VDD2.n176 VDD2.n175 185
R3467 VDD2.n109 VDD2.n108 185
R3468 VDD2.n170 VDD2.n169 185
R3469 VDD2.n168 VDD2.n167 185
R3470 VDD2.n113 VDD2.n112 185
R3471 VDD2.n162 VDD2.n161 185
R3472 VDD2.n160 VDD2.n159 185
R3473 VDD2.n117 VDD2.n116 185
R3474 VDD2.n154 VDD2.n153 185
R3475 VDD2.n152 VDD2.n119 185
R3476 VDD2.n151 VDD2.n150 185
R3477 VDD2.n122 VDD2.n120 185
R3478 VDD2.n145 VDD2.n144 185
R3479 VDD2.n143 VDD2.n142 185
R3480 VDD2.n126 VDD2.n125 185
R3481 VDD2.n137 VDD2.n136 185
R3482 VDD2.n135 VDD2.n134 185
R3483 VDD2.n130 VDD2.n129 185
R3484 VDD2.n30 VDD2.n29 185
R3485 VDD2.n35 VDD2.n34 185
R3486 VDD2.n37 VDD2.n36 185
R3487 VDD2.n26 VDD2.n25 185
R3488 VDD2.n43 VDD2.n42 185
R3489 VDD2.n45 VDD2.n44 185
R3490 VDD2.n22 VDD2.n21 185
R3491 VDD2.n52 VDD2.n51 185
R3492 VDD2.n53 VDD2.n20 185
R3493 VDD2.n55 VDD2.n54 185
R3494 VDD2.n18 VDD2.n17 185
R3495 VDD2.n61 VDD2.n60 185
R3496 VDD2.n63 VDD2.n62 185
R3497 VDD2.n14 VDD2.n13 185
R3498 VDD2.n69 VDD2.n68 185
R3499 VDD2.n71 VDD2.n70 185
R3500 VDD2.n10 VDD2.n9 185
R3501 VDD2.n77 VDD2.n76 185
R3502 VDD2.n79 VDD2.n78 185
R3503 VDD2.n6 VDD2.n5 185
R3504 VDD2.n85 VDD2.n84 185
R3505 VDD2.n87 VDD2.n86 185
R3506 VDD2.n2 VDD2.n1 185
R3507 VDD2.n93 VDD2.n92 185
R3508 VDD2.n131 VDD2.t2 149.524
R3509 VDD2.n31 VDD2.t5 149.524
R3510 VDD2.n192 VDD2.n100 104.615
R3511 VDD2.n185 VDD2.n100 104.615
R3512 VDD2.n185 VDD2.n184 104.615
R3513 VDD2.n184 VDD2.n104 104.615
R3514 VDD2.n177 VDD2.n104 104.615
R3515 VDD2.n177 VDD2.n176 104.615
R3516 VDD2.n176 VDD2.n108 104.615
R3517 VDD2.n169 VDD2.n108 104.615
R3518 VDD2.n169 VDD2.n168 104.615
R3519 VDD2.n168 VDD2.n112 104.615
R3520 VDD2.n161 VDD2.n112 104.615
R3521 VDD2.n161 VDD2.n160 104.615
R3522 VDD2.n160 VDD2.n116 104.615
R3523 VDD2.n153 VDD2.n116 104.615
R3524 VDD2.n153 VDD2.n152 104.615
R3525 VDD2.n152 VDD2.n151 104.615
R3526 VDD2.n151 VDD2.n120 104.615
R3527 VDD2.n144 VDD2.n120 104.615
R3528 VDD2.n144 VDD2.n143 104.615
R3529 VDD2.n143 VDD2.n125 104.615
R3530 VDD2.n136 VDD2.n125 104.615
R3531 VDD2.n136 VDD2.n135 104.615
R3532 VDD2.n135 VDD2.n129 104.615
R3533 VDD2.n35 VDD2.n29 104.615
R3534 VDD2.n36 VDD2.n35 104.615
R3535 VDD2.n36 VDD2.n25 104.615
R3536 VDD2.n43 VDD2.n25 104.615
R3537 VDD2.n44 VDD2.n43 104.615
R3538 VDD2.n44 VDD2.n21 104.615
R3539 VDD2.n52 VDD2.n21 104.615
R3540 VDD2.n53 VDD2.n52 104.615
R3541 VDD2.n54 VDD2.n53 104.615
R3542 VDD2.n54 VDD2.n17 104.615
R3543 VDD2.n61 VDD2.n17 104.615
R3544 VDD2.n62 VDD2.n61 104.615
R3545 VDD2.n62 VDD2.n13 104.615
R3546 VDD2.n69 VDD2.n13 104.615
R3547 VDD2.n70 VDD2.n69 104.615
R3548 VDD2.n70 VDD2.n9 104.615
R3549 VDD2.n77 VDD2.n9 104.615
R3550 VDD2.n78 VDD2.n77 104.615
R3551 VDD2.n78 VDD2.n5 104.615
R3552 VDD2.n85 VDD2.n5 104.615
R3553 VDD2.n86 VDD2.n85 104.615
R3554 VDD2.n86 VDD2.n1 104.615
R3555 VDD2.n93 VDD2.n1 104.615
R3556 VDD2.n98 VDD2.n97 66.5645
R3557 VDD2 VDD2.n197 66.5615
R3558 VDD2.n196 VDD2.n195 64.5066
R3559 VDD2.n96 VDD2.n95 64.5056
R3560 VDD2.n96 VDD2.n94 54.2043
R3561 VDD2.t2 VDD2.n129 52.3082
R3562 VDD2.t5 VDD2.n29 52.3082
R3563 VDD2.n194 VDD2.n98 52.0968
R3564 VDD2.n194 VDD2.n193 51.3853
R3565 VDD2.n154 VDD2.n119 13.1884
R3566 VDD2.n55 VDD2.n20 13.1884
R3567 VDD2.n155 VDD2.n117 12.8005
R3568 VDD2.n150 VDD2.n121 12.8005
R3569 VDD2.n51 VDD2.n50 12.8005
R3570 VDD2.n56 VDD2.n18 12.8005
R3571 VDD2.n159 VDD2.n158 12.0247
R3572 VDD2.n149 VDD2.n122 12.0247
R3573 VDD2.n49 VDD2.n22 12.0247
R3574 VDD2.n60 VDD2.n59 12.0247
R3575 VDD2.n191 VDD2.n99 11.249
R3576 VDD2.n162 VDD2.n115 11.249
R3577 VDD2.n146 VDD2.n145 11.249
R3578 VDD2.n46 VDD2.n45 11.249
R3579 VDD2.n63 VDD2.n16 11.249
R3580 VDD2.n92 VDD2.n0 11.249
R3581 VDD2.n190 VDD2.n101 10.4732
R3582 VDD2.n163 VDD2.n113 10.4732
R3583 VDD2.n142 VDD2.n124 10.4732
R3584 VDD2.n42 VDD2.n24 10.4732
R3585 VDD2.n64 VDD2.n14 10.4732
R3586 VDD2.n91 VDD2.n2 10.4732
R3587 VDD2.n131 VDD2.n130 10.2747
R3588 VDD2.n31 VDD2.n30 10.2747
R3589 VDD2.n187 VDD2.n186 9.69747
R3590 VDD2.n167 VDD2.n166 9.69747
R3591 VDD2.n141 VDD2.n126 9.69747
R3592 VDD2.n41 VDD2.n26 9.69747
R3593 VDD2.n68 VDD2.n67 9.69747
R3594 VDD2.n88 VDD2.n87 9.69747
R3595 VDD2.n189 VDD2.n99 9.45567
R3596 VDD2.n90 VDD2.n0 9.45567
R3597 VDD2.n133 VDD2.n132 9.3005
R3598 VDD2.n128 VDD2.n127 9.3005
R3599 VDD2.n139 VDD2.n138 9.3005
R3600 VDD2.n141 VDD2.n140 9.3005
R3601 VDD2.n124 VDD2.n123 9.3005
R3602 VDD2.n147 VDD2.n146 9.3005
R3603 VDD2.n149 VDD2.n148 9.3005
R3604 VDD2.n121 VDD2.n118 9.3005
R3605 VDD2.n180 VDD2.n179 9.3005
R3606 VDD2.n182 VDD2.n181 9.3005
R3607 VDD2.n103 VDD2.n102 9.3005
R3608 VDD2.n188 VDD2.n187 9.3005
R3609 VDD2.n190 VDD2.n189 9.3005
R3610 VDD2.n107 VDD2.n106 9.3005
R3611 VDD2.n174 VDD2.n173 9.3005
R3612 VDD2.n172 VDD2.n171 9.3005
R3613 VDD2.n111 VDD2.n110 9.3005
R3614 VDD2.n166 VDD2.n165 9.3005
R3615 VDD2.n164 VDD2.n163 9.3005
R3616 VDD2.n115 VDD2.n114 9.3005
R3617 VDD2.n158 VDD2.n157 9.3005
R3618 VDD2.n156 VDD2.n155 9.3005
R3619 VDD2.n8 VDD2.n7 9.3005
R3620 VDD2.n81 VDD2.n80 9.3005
R3621 VDD2.n83 VDD2.n82 9.3005
R3622 VDD2.n4 VDD2.n3 9.3005
R3623 VDD2.n89 VDD2.n88 9.3005
R3624 VDD2.n91 VDD2.n90 9.3005
R3625 VDD2.n73 VDD2.n72 9.3005
R3626 VDD2.n12 VDD2.n11 9.3005
R3627 VDD2.n67 VDD2.n66 9.3005
R3628 VDD2.n65 VDD2.n64 9.3005
R3629 VDD2.n16 VDD2.n15 9.3005
R3630 VDD2.n59 VDD2.n58 9.3005
R3631 VDD2.n57 VDD2.n56 9.3005
R3632 VDD2.n33 VDD2.n32 9.3005
R3633 VDD2.n28 VDD2.n27 9.3005
R3634 VDD2.n39 VDD2.n38 9.3005
R3635 VDD2.n41 VDD2.n40 9.3005
R3636 VDD2.n24 VDD2.n23 9.3005
R3637 VDD2.n47 VDD2.n46 9.3005
R3638 VDD2.n49 VDD2.n48 9.3005
R3639 VDD2.n50 VDD2.n19 9.3005
R3640 VDD2.n75 VDD2.n74 9.3005
R3641 VDD2.n183 VDD2.n103 8.92171
R3642 VDD2.n170 VDD2.n111 8.92171
R3643 VDD2.n138 VDD2.n137 8.92171
R3644 VDD2.n38 VDD2.n37 8.92171
R3645 VDD2.n71 VDD2.n12 8.92171
R3646 VDD2.n84 VDD2.n4 8.92171
R3647 VDD2.n182 VDD2.n105 8.14595
R3648 VDD2.n171 VDD2.n109 8.14595
R3649 VDD2.n134 VDD2.n128 8.14595
R3650 VDD2.n34 VDD2.n28 8.14595
R3651 VDD2.n72 VDD2.n10 8.14595
R3652 VDD2.n83 VDD2.n6 8.14595
R3653 VDD2.n179 VDD2.n178 7.3702
R3654 VDD2.n175 VDD2.n174 7.3702
R3655 VDD2.n133 VDD2.n130 7.3702
R3656 VDD2.n33 VDD2.n30 7.3702
R3657 VDD2.n76 VDD2.n75 7.3702
R3658 VDD2.n80 VDD2.n79 7.3702
R3659 VDD2.n178 VDD2.n107 6.59444
R3660 VDD2.n175 VDD2.n107 6.59444
R3661 VDD2.n76 VDD2.n8 6.59444
R3662 VDD2.n79 VDD2.n8 6.59444
R3663 VDD2.n179 VDD2.n105 5.81868
R3664 VDD2.n174 VDD2.n109 5.81868
R3665 VDD2.n134 VDD2.n133 5.81868
R3666 VDD2.n34 VDD2.n33 5.81868
R3667 VDD2.n75 VDD2.n10 5.81868
R3668 VDD2.n80 VDD2.n6 5.81868
R3669 VDD2.n183 VDD2.n182 5.04292
R3670 VDD2.n171 VDD2.n170 5.04292
R3671 VDD2.n137 VDD2.n128 5.04292
R3672 VDD2.n37 VDD2.n28 5.04292
R3673 VDD2.n72 VDD2.n71 5.04292
R3674 VDD2.n84 VDD2.n83 5.04292
R3675 VDD2.n186 VDD2.n103 4.26717
R3676 VDD2.n167 VDD2.n111 4.26717
R3677 VDD2.n138 VDD2.n126 4.26717
R3678 VDD2.n38 VDD2.n26 4.26717
R3679 VDD2.n68 VDD2.n12 4.26717
R3680 VDD2.n87 VDD2.n4 4.26717
R3681 VDD2.n187 VDD2.n101 3.49141
R3682 VDD2.n166 VDD2.n113 3.49141
R3683 VDD2.n142 VDD2.n141 3.49141
R3684 VDD2.n42 VDD2.n41 3.49141
R3685 VDD2.n67 VDD2.n14 3.49141
R3686 VDD2.n88 VDD2.n2 3.49141
R3687 VDD2.n32 VDD2.n31 2.84303
R3688 VDD2.n132 VDD2.n131 2.84303
R3689 VDD2.n196 VDD2.n194 2.81947
R3690 VDD2.n191 VDD2.n190 2.71565
R3691 VDD2.n163 VDD2.n162 2.71565
R3692 VDD2.n145 VDD2.n124 2.71565
R3693 VDD2.n45 VDD2.n24 2.71565
R3694 VDD2.n64 VDD2.n63 2.71565
R3695 VDD2.n92 VDD2.n91 2.71565
R3696 VDD2.n193 VDD2.n99 1.93989
R3697 VDD2.n159 VDD2.n115 1.93989
R3698 VDD2.n146 VDD2.n122 1.93989
R3699 VDD2.n46 VDD2.n22 1.93989
R3700 VDD2.n60 VDD2.n16 1.93989
R3701 VDD2.n94 VDD2.n0 1.93989
R3702 VDD2.n158 VDD2.n117 1.16414
R3703 VDD2.n150 VDD2.n149 1.16414
R3704 VDD2.n51 VDD2.n49 1.16414
R3705 VDD2.n59 VDD2.n18 1.16414
R3706 VDD2.n197 VDD2.t6 1.13909
R3707 VDD2.n197 VDD2.t1 1.13909
R3708 VDD2.n195 VDD2.t0 1.13909
R3709 VDD2.n195 VDD2.t7 1.13909
R3710 VDD2.n97 VDD2.t8 1.13909
R3711 VDD2.n97 VDD2.t3 1.13909
R3712 VDD2.n95 VDD2.t9 1.13909
R3713 VDD2.n95 VDD2.t4 1.13909
R3714 VDD2 VDD2.n196 0.763431
R3715 VDD2.n98 VDD2.n96 0.649895
R3716 VDD2.n155 VDD2.n154 0.388379
R3717 VDD2.n121 VDD2.n119 0.388379
R3718 VDD2.n50 VDD2.n20 0.388379
R3719 VDD2.n56 VDD2.n55 0.388379
R3720 VDD2.n189 VDD2.n188 0.155672
R3721 VDD2.n188 VDD2.n102 0.155672
R3722 VDD2.n181 VDD2.n102 0.155672
R3723 VDD2.n181 VDD2.n180 0.155672
R3724 VDD2.n180 VDD2.n106 0.155672
R3725 VDD2.n173 VDD2.n106 0.155672
R3726 VDD2.n173 VDD2.n172 0.155672
R3727 VDD2.n172 VDD2.n110 0.155672
R3728 VDD2.n165 VDD2.n110 0.155672
R3729 VDD2.n165 VDD2.n164 0.155672
R3730 VDD2.n164 VDD2.n114 0.155672
R3731 VDD2.n157 VDD2.n114 0.155672
R3732 VDD2.n157 VDD2.n156 0.155672
R3733 VDD2.n156 VDD2.n118 0.155672
R3734 VDD2.n148 VDD2.n118 0.155672
R3735 VDD2.n148 VDD2.n147 0.155672
R3736 VDD2.n147 VDD2.n123 0.155672
R3737 VDD2.n140 VDD2.n123 0.155672
R3738 VDD2.n140 VDD2.n139 0.155672
R3739 VDD2.n139 VDD2.n127 0.155672
R3740 VDD2.n132 VDD2.n127 0.155672
R3741 VDD2.n32 VDD2.n27 0.155672
R3742 VDD2.n39 VDD2.n27 0.155672
R3743 VDD2.n40 VDD2.n39 0.155672
R3744 VDD2.n40 VDD2.n23 0.155672
R3745 VDD2.n47 VDD2.n23 0.155672
R3746 VDD2.n48 VDD2.n47 0.155672
R3747 VDD2.n48 VDD2.n19 0.155672
R3748 VDD2.n57 VDD2.n19 0.155672
R3749 VDD2.n58 VDD2.n57 0.155672
R3750 VDD2.n58 VDD2.n15 0.155672
R3751 VDD2.n65 VDD2.n15 0.155672
R3752 VDD2.n66 VDD2.n65 0.155672
R3753 VDD2.n66 VDD2.n11 0.155672
R3754 VDD2.n73 VDD2.n11 0.155672
R3755 VDD2.n74 VDD2.n73 0.155672
R3756 VDD2.n74 VDD2.n7 0.155672
R3757 VDD2.n81 VDD2.n7 0.155672
R3758 VDD2.n82 VDD2.n81 0.155672
R3759 VDD2.n82 VDD2.n3 0.155672
R3760 VDD2.n89 VDD2.n3 0.155672
R3761 VDD2.n90 VDD2.n89 0.155672
C0 VDD2 VTAIL 12.8925f
C1 VDD2 VDD1 2.39616f
C2 VP VDD2 0.627314f
C3 VTAIL VDD1 12.839999f
C4 VN VDD2 15.5879f
C5 VP VTAIL 16.1481f
C6 VP VDD1 16.0564f
C7 VN VTAIL 16.133799f
C8 VN VDD1 0.154108f
C9 VP VN 9.896719f
C10 VDD2 B 8.537965f
C11 VDD1 B 8.528261f
C12 VTAIL B 10.643201f
C13 VN B 20.18013f
C14 VP B 18.665607f
C15 VDD2.n0 B 0.013342f
C16 VDD2.n1 B 0.03002f
C17 VDD2.n2 B 0.013448f
C18 VDD2.n3 B 0.023636f
C19 VDD2.n4 B 0.012701f
C20 VDD2.n5 B 0.03002f
C21 VDD2.n6 B 0.013448f
C22 VDD2.n7 B 0.023636f
C23 VDD2.n8 B 0.012701f
C24 VDD2.n9 B 0.03002f
C25 VDD2.n10 B 0.013448f
C26 VDD2.n11 B 0.023636f
C27 VDD2.n12 B 0.012701f
C28 VDD2.n13 B 0.03002f
C29 VDD2.n14 B 0.013448f
C30 VDD2.n15 B 0.023636f
C31 VDD2.n16 B 0.012701f
C32 VDD2.n17 B 0.03002f
C33 VDD2.n18 B 0.013448f
C34 VDD2.n19 B 0.023636f
C35 VDD2.n20 B 0.013075f
C36 VDD2.n21 B 0.03002f
C37 VDD2.n22 B 0.013448f
C38 VDD2.n23 B 0.023636f
C39 VDD2.n24 B 0.012701f
C40 VDD2.n25 B 0.03002f
C41 VDD2.n26 B 0.013448f
C42 VDD2.n27 B 0.023636f
C43 VDD2.n28 B 0.012701f
C44 VDD2.n29 B 0.022515f
C45 VDD2.n30 B 0.021222f
C46 VDD2.t5 B 0.051389f
C47 VDD2.n31 B 0.219323f
C48 VDD2.n32 B 1.75905f
C49 VDD2.n33 B 0.012701f
C50 VDD2.n34 B 0.013448f
C51 VDD2.n35 B 0.03002f
C52 VDD2.n36 B 0.03002f
C53 VDD2.n37 B 0.013448f
C54 VDD2.n38 B 0.012701f
C55 VDD2.n39 B 0.023636f
C56 VDD2.n40 B 0.023636f
C57 VDD2.n41 B 0.012701f
C58 VDD2.n42 B 0.013448f
C59 VDD2.n43 B 0.03002f
C60 VDD2.n44 B 0.03002f
C61 VDD2.n45 B 0.013448f
C62 VDD2.n46 B 0.012701f
C63 VDD2.n47 B 0.023636f
C64 VDD2.n48 B 0.023636f
C65 VDD2.n49 B 0.012701f
C66 VDD2.n50 B 0.012701f
C67 VDD2.n51 B 0.013448f
C68 VDD2.n52 B 0.03002f
C69 VDD2.n53 B 0.03002f
C70 VDD2.n54 B 0.03002f
C71 VDD2.n55 B 0.013075f
C72 VDD2.n56 B 0.012701f
C73 VDD2.n57 B 0.023636f
C74 VDD2.n58 B 0.023636f
C75 VDD2.n59 B 0.012701f
C76 VDD2.n60 B 0.013448f
C77 VDD2.n61 B 0.03002f
C78 VDD2.n62 B 0.03002f
C79 VDD2.n63 B 0.013448f
C80 VDD2.n64 B 0.012701f
C81 VDD2.n65 B 0.023636f
C82 VDD2.n66 B 0.023636f
C83 VDD2.n67 B 0.012701f
C84 VDD2.n68 B 0.013448f
C85 VDD2.n69 B 0.03002f
C86 VDD2.n70 B 0.03002f
C87 VDD2.n71 B 0.013448f
C88 VDD2.n72 B 0.012701f
C89 VDD2.n73 B 0.023636f
C90 VDD2.n74 B 0.023636f
C91 VDD2.n75 B 0.012701f
C92 VDD2.n76 B 0.013448f
C93 VDD2.n77 B 0.03002f
C94 VDD2.n78 B 0.03002f
C95 VDD2.n79 B 0.013448f
C96 VDD2.n80 B 0.012701f
C97 VDD2.n81 B 0.023636f
C98 VDD2.n82 B 0.023636f
C99 VDD2.n83 B 0.012701f
C100 VDD2.n84 B 0.013448f
C101 VDD2.n85 B 0.03002f
C102 VDD2.n86 B 0.03002f
C103 VDD2.n87 B 0.013448f
C104 VDD2.n88 B 0.012701f
C105 VDD2.n89 B 0.023636f
C106 VDD2.n90 B 0.06206f
C107 VDD2.n91 B 0.012701f
C108 VDD2.n92 B 0.013448f
C109 VDD2.n93 B 0.060195f
C110 VDD2.n94 B 0.081605f
C111 VDD2.t9 B 0.324809f
C112 VDD2.t4 B 0.324809f
C113 VDD2.n95 B 2.96524f
C114 VDD2.n96 B 0.699459f
C115 VDD2.t8 B 0.324809f
C116 VDD2.t3 B 0.324809f
C117 VDD2.n97 B 2.98277f
C118 VDD2.n98 B 3.22576f
C119 VDD2.n99 B 0.013342f
C120 VDD2.n100 B 0.03002f
C121 VDD2.n101 B 0.013448f
C122 VDD2.n102 B 0.023636f
C123 VDD2.n103 B 0.012701f
C124 VDD2.n104 B 0.03002f
C125 VDD2.n105 B 0.013448f
C126 VDD2.n106 B 0.023636f
C127 VDD2.n107 B 0.012701f
C128 VDD2.n108 B 0.03002f
C129 VDD2.n109 B 0.013448f
C130 VDD2.n110 B 0.023636f
C131 VDD2.n111 B 0.012701f
C132 VDD2.n112 B 0.03002f
C133 VDD2.n113 B 0.013448f
C134 VDD2.n114 B 0.023636f
C135 VDD2.n115 B 0.012701f
C136 VDD2.n116 B 0.03002f
C137 VDD2.n117 B 0.013448f
C138 VDD2.n118 B 0.023636f
C139 VDD2.n119 B 0.013075f
C140 VDD2.n120 B 0.03002f
C141 VDD2.n121 B 0.012701f
C142 VDD2.n122 B 0.013448f
C143 VDD2.n123 B 0.023636f
C144 VDD2.n124 B 0.012701f
C145 VDD2.n125 B 0.03002f
C146 VDD2.n126 B 0.013448f
C147 VDD2.n127 B 0.023636f
C148 VDD2.n128 B 0.012701f
C149 VDD2.n129 B 0.022515f
C150 VDD2.n130 B 0.021222f
C151 VDD2.t2 B 0.051389f
C152 VDD2.n131 B 0.219324f
C153 VDD2.n132 B 1.75905f
C154 VDD2.n133 B 0.012701f
C155 VDD2.n134 B 0.013448f
C156 VDD2.n135 B 0.03002f
C157 VDD2.n136 B 0.03002f
C158 VDD2.n137 B 0.013448f
C159 VDD2.n138 B 0.012701f
C160 VDD2.n139 B 0.023636f
C161 VDD2.n140 B 0.023636f
C162 VDD2.n141 B 0.012701f
C163 VDD2.n142 B 0.013448f
C164 VDD2.n143 B 0.03002f
C165 VDD2.n144 B 0.03002f
C166 VDD2.n145 B 0.013448f
C167 VDD2.n146 B 0.012701f
C168 VDD2.n147 B 0.023636f
C169 VDD2.n148 B 0.023636f
C170 VDD2.n149 B 0.012701f
C171 VDD2.n150 B 0.013448f
C172 VDD2.n151 B 0.03002f
C173 VDD2.n152 B 0.03002f
C174 VDD2.n153 B 0.03002f
C175 VDD2.n154 B 0.013075f
C176 VDD2.n155 B 0.012701f
C177 VDD2.n156 B 0.023636f
C178 VDD2.n157 B 0.023636f
C179 VDD2.n158 B 0.012701f
C180 VDD2.n159 B 0.013448f
C181 VDD2.n160 B 0.03002f
C182 VDD2.n161 B 0.03002f
C183 VDD2.n162 B 0.013448f
C184 VDD2.n163 B 0.012701f
C185 VDD2.n164 B 0.023636f
C186 VDD2.n165 B 0.023636f
C187 VDD2.n166 B 0.012701f
C188 VDD2.n167 B 0.013448f
C189 VDD2.n168 B 0.03002f
C190 VDD2.n169 B 0.03002f
C191 VDD2.n170 B 0.013448f
C192 VDD2.n171 B 0.012701f
C193 VDD2.n172 B 0.023636f
C194 VDD2.n173 B 0.023636f
C195 VDD2.n174 B 0.012701f
C196 VDD2.n175 B 0.013448f
C197 VDD2.n176 B 0.03002f
C198 VDD2.n177 B 0.03002f
C199 VDD2.n178 B 0.013448f
C200 VDD2.n179 B 0.012701f
C201 VDD2.n180 B 0.023636f
C202 VDD2.n181 B 0.023636f
C203 VDD2.n182 B 0.012701f
C204 VDD2.n183 B 0.013448f
C205 VDD2.n184 B 0.03002f
C206 VDD2.n185 B 0.03002f
C207 VDD2.n186 B 0.013448f
C208 VDD2.n187 B 0.012701f
C209 VDD2.n188 B 0.023636f
C210 VDD2.n189 B 0.06206f
C211 VDD2.n190 B 0.012701f
C212 VDD2.n191 B 0.013448f
C213 VDD2.n192 B 0.060195f
C214 VDD2.n193 B 0.067947f
C215 VDD2.n194 B 3.24846f
C216 VDD2.t0 B 0.324809f
C217 VDD2.t7 B 0.324809f
C218 VDD2.n195 B 2.96523f
C219 VDD2.n196 B 0.458317f
C220 VDD2.t6 B 0.324809f
C221 VDD2.t1 B 0.324809f
C222 VDD2.n197 B 2.98272f
C223 VN.n0 B 0.024974f
C224 VN.t6 B 2.66211f
C225 VN.n1 B 0.038034f
C226 VN.n2 B 0.018943f
C227 VN.n3 B 0.025892f
C228 VN.n4 B 0.018943f
C229 VN.n5 B 0.020268f
C230 VN.n6 B 0.018943f
C231 VN.t5 B 2.66211f
C232 VN.n7 B 0.035305f
C233 VN.n8 B 0.018943f
C234 VN.n9 B 0.035305f
C235 VN.t4 B 2.85834f
C236 VN.n10 B 0.953105f
C237 VN.t0 B 2.66211f
C238 VN.n11 B 0.982398f
C239 VN.n12 B 0.027287f
C240 VN.n13 B 0.20179f
C241 VN.n14 B 0.018943f
C242 VN.n15 B 0.018943f
C243 VN.n16 B 0.03341f
C244 VN.n17 B 0.020268f
C245 VN.n18 B 0.036937f
C246 VN.n19 B 0.018943f
C247 VN.n20 B 0.018943f
C248 VN.n21 B 0.018943f
C249 VN.n22 B 0.940018f
C250 VN.n23 B 0.035305f
C251 VN.n24 B 0.036937f
C252 VN.n25 B 0.018943f
C253 VN.n26 B 0.018943f
C254 VN.n27 B 0.018943f
C255 VN.n28 B 0.03341f
C256 VN.n29 B 0.035305f
C257 VN.t1 B 2.66211f
C258 VN.n30 B 0.922143f
C259 VN.n31 B 0.027287f
C260 VN.n32 B 0.018943f
C261 VN.n33 B 0.018943f
C262 VN.n34 B 0.018943f
C263 VN.n35 B 0.035305f
C264 VN.n36 B 0.034951f
C265 VN.n37 B 0.01763f
C266 VN.n38 B 0.018943f
C267 VN.n39 B 0.018943f
C268 VN.n40 B 0.018943f
C269 VN.n41 B 0.035305f
C270 VN.n42 B 0.019269f
C271 VN.n43 B 0.985833f
C272 VN.n44 B 0.036787f
C273 VN.n45 B 0.024974f
C274 VN.t7 B 2.66211f
C275 VN.n46 B 0.038034f
C276 VN.n47 B 0.018943f
C277 VN.n48 B 0.025892f
C278 VN.n49 B 0.018943f
C279 VN.t9 B 2.66211f
C280 VN.n50 B 0.922143f
C281 VN.n51 B 0.020268f
C282 VN.n52 B 0.018943f
C283 VN.t2 B 2.66211f
C284 VN.n53 B 0.035305f
C285 VN.n54 B 0.018943f
C286 VN.n55 B 0.035305f
C287 VN.t8 B 2.85834f
C288 VN.n56 B 0.953105f
C289 VN.t3 B 2.66211f
C290 VN.n57 B 0.982398f
C291 VN.n58 B 0.027287f
C292 VN.n59 B 0.20179f
C293 VN.n60 B 0.018943f
C294 VN.n61 B 0.018943f
C295 VN.n62 B 0.03341f
C296 VN.n63 B 0.020268f
C297 VN.n64 B 0.036937f
C298 VN.n65 B 0.018943f
C299 VN.n66 B 0.018943f
C300 VN.n67 B 0.018943f
C301 VN.n68 B 0.940018f
C302 VN.n69 B 0.035305f
C303 VN.n70 B 0.036937f
C304 VN.n71 B 0.018943f
C305 VN.n72 B 0.018943f
C306 VN.n73 B 0.018943f
C307 VN.n74 B 0.03341f
C308 VN.n75 B 0.035305f
C309 VN.n76 B 0.027287f
C310 VN.n77 B 0.018943f
C311 VN.n78 B 0.018943f
C312 VN.n79 B 0.018943f
C313 VN.n80 B 0.035305f
C314 VN.n81 B 0.034951f
C315 VN.n82 B 0.01763f
C316 VN.n83 B 0.018943f
C317 VN.n84 B 0.018943f
C318 VN.n85 B 0.018943f
C319 VN.n86 B 0.035305f
C320 VN.n87 B 0.019269f
C321 VN.n88 B 0.985833f
C322 VN.n89 B 1.34942f
C323 VDD1.n0 B 0.013477f
C324 VDD1.n1 B 0.030323f
C325 VDD1.n2 B 0.013584f
C326 VDD1.n3 B 0.023875f
C327 VDD1.n4 B 0.012829f
C328 VDD1.n5 B 0.030323f
C329 VDD1.n6 B 0.013584f
C330 VDD1.n7 B 0.023875f
C331 VDD1.n8 B 0.012829f
C332 VDD1.n9 B 0.030323f
C333 VDD1.n10 B 0.013584f
C334 VDD1.n11 B 0.023875f
C335 VDD1.n12 B 0.012829f
C336 VDD1.n13 B 0.030323f
C337 VDD1.n14 B 0.013584f
C338 VDD1.n15 B 0.023875f
C339 VDD1.n16 B 0.012829f
C340 VDD1.n17 B 0.030323f
C341 VDD1.n18 B 0.013584f
C342 VDD1.n19 B 0.023875f
C343 VDD1.n20 B 0.013207f
C344 VDD1.n21 B 0.030323f
C345 VDD1.n22 B 0.012829f
C346 VDD1.n23 B 0.013584f
C347 VDD1.n24 B 0.023875f
C348 VDD1.n25 B 0.012829f
C349 VDD1.n26 B 0.030323f
C350 VDD1.n27 B 0.013584f
C351 VDD1.n28 B 0.023875f
C352 VDD1.n29 B 0.012829f
C353 VDD1.n30 B 0.022743f
C354 VDD1.n31 B 0.021436f
C355 VDD1.t3 B 0.051907f
C356 VDD1.n32 B 0.221537f
C357 VDD1.n33 B 1.7768f
C358 VDD1.n34 B 0.012829f
C359 VDD1.n35 B 0.013584f
C360 VDD1.n36 B 0.030323f
C361 VDD1.n37 B 0.030323f
C362 VDD1.n38 B 0.013584f
C363 VDD1.n39 B 0.012829f
C364 VDD1.n40 B 0.023875f
C365 VDD1.n41 B 0.023875f
C366 VDD1.n42 B 0.012829f
C367 VDD1.n43 B 0.013584f
C368 VDD1.n44 B 0.030323f
C369 VDD1.n45 B 0.030323f
C370 VDD1.n46 B 0.013584f
C371 VDD1.n47 B 0.012829f
C372 VDD1.n48 B 0.023875f
C373 VDD1.n49 B 0.023875f
C374 VDD1.n50 B 0.012829f
C375 VDD1.n51 B 0.013584f
C376 VDD1.n52 B 0.030323f
C377 VDD1.n53 B 0.030323f
C378 VDD1.n54 B 0.030323f
C379 VDD1.n55 B 0.013207f
C380 VDD1.n56 B 0.012829f
C381 VDD1.n57 B 0.023875f
C382 VDD1.n58 B 0.023875f
C383 VDD1.n59 B 0.012829f
C384 VDD1.n60 B 0.013584f
C385 VDD1.n61 B 0.030323f
C386 VDD1.n62 B 0.030323f
C387 VDD1.n63 B 0.013584f
C388 VDD1.n64 B 0.012829f
C389 VDD1.n65 B 0.023875f
C390 VDD1.n66 B 0.023875f
C391 VDD1.n67 B 0.012829f
C392 VDD1.n68 B 0.013584f
C393 VDD1.n69 B 0.030323f
C394 VDD1.n70 B 0.030323f
C395 VDD1.n71 B 0.013584f
C396 VDD1.n72 B 0.012829f
C397 VDD1.n73 B 0.023875f
C398 VDD1.n74 B 0.023875f
C399 VDD1.n75 B 0.012829f
C400 VDD1.n76 B 0.013584f
C401 VDD1.n77 B 0.030323f
C402 VDD1.n78 B 0.030323f
C403 VDD1.n79 B 0.013584f
C404 VDD1.n80 B 0.012829f
C405 VDD1.n81 B 0.023875f
C406 VDD1.n82 B 0.023875f
C407 VDD1.n83 B 0.012829f
C408 VDD1.n84 B 0.013584f
C409 VDD1.n85 B 0.030323f
C410 VDD1.n86 B 0.030323f
C411 VDD1.n87 B 0.013584f
C412 VDD1.n88 B 0.012829f
C413 VDD1.n89 B 0.023875f
C414 VDD1.n90 B 0.062686f
C415 VDD1.n91 B 0.012829f
C416 VDD1.n92 B 0.013584f
C417 VDD1.n93 B 0.060803f
C418 VDD1.n94 B 0.082428f
C419 VDD1.t8 B 0.328087f
C420 VDD1.t0 B 0.328087f
C421 VDD1.n95 B 2.99515f
C422 VDD1.n96 B 0.714407f
C423 VDD1.n97 B 0.013477f
C424 VDD1.n98 B 0.030323f
C425 VDD1.n99 B 0.013584f
C426 VDD1.n100 B 0.023875f
C427 VDD1.n101 B 0.012829f
C428 VDD1.n102 B 0.030323f
C429 VDD1.n103 B 0.013584f
C430 VDD1.n104 B 0.023875f
C431 VDD1.n105 B 0.012829f
C432 VDD1.n106 B 0.030323f
C433 VDD1.n107 B 0.013584f
C434 VDD1.n108 B 0.023875f
C435 VDD1.n109 B 0.012829f
C436 VDD1.n110 B 0.030323f
C437 VDD1.n111 B 0.013584f
C438 VDD1.n112 B 0.023875f
C439 VDD1.n113 B 0.012829f
C440 VDD1.n114 B 0.030323f
C441 VDD1.n115 B 0.013584f
C442 VDD1.n116 B 0.023875f
C443 VDD1.n117 B 0.013207f
C444 VDD1.n118 B 0.030323f
C445 VDD1.n119 B 0.013584f
C446 VDD1.n120 B 0.023875f
C447 VDD1.n121 B 0.012829f
C448 VDD1.n122 B 0.030323f
C449 VDD1.n123 B 0.013584f
C450 VDD1.n124 B 0.023875f
C451 VDD1.n125 B 0.012829f
C452 VDD1.n126 B 0.022743f
C453 VDD1.n127 B 0.021436f
C454 VDD1.t1 B 0.051907f
C455 VDD1.n128 B 0.221537f
C456 VDD1.n129 B 1.7768f
C457 VDD1.n130 B 0.012829f
C458 VDD1.n131 B 0.013584f
C459 VDD1.n132 B 0.030323f
C460 VDD1.n133 B 0.030323f
C461 VDD1.n134 B 0.013584f
C462 VDD1.n135 B 0.012829f
C463 VDD1.n136 B 0.023875f
C464 VDD1.n137 B 0.023875f
C465 VDD1.n138 B 0.012829f
C466 VDD1.n139 B 0.013584f
C467 VDD1.n140 B 0.030323f
C468 VDD1.n141 B 0.030323f
C469 VDD1.n142 B 0.013584f
C470 VDD1.n143 B 0.012829f
C471 VDD1.n144 B 0.023875f
C472 VDD1.n145 B 0.023875f
C473 VDD1.n146 B 0.012829f
C474 VDD1.n147 B 0.012829f
C475 VDD1.n148 B 0.013584f
C476 VDD1.n149 B 0.030323f
C477 VDD1.n150 B 0.030323f
C478 VDD1.n151 B 0.030323f
C479 VDD1.n152 B 0.013207f
C480 VDD1.n153 B 0.012829f
C481 VDD1.n154 B 0.023875f
C482 VDD1.n155 B 0.023875f
C483 VDD1.n156 B 0.012829f
C484 VDD1.n157 B 0.013584f
C485 VDD1.n158 B 0.030323f
C486 VDD1.n159 B 0.030323f
C487 VDD1.n160 B 0.013584f
C488 VDD1.n161 B 0.012829f
C489 VDD1.n162 B 0.023875f
C490 VDD1.n163 B 0.023875f
C491 VDD1.n164 B 0.012829f
C492 VDD1.n165 B 0.013584f
C493 VDD1.n166 B 0.030323f
C494 VDD1.n167 B 0.030323f
C495 VDD1.n168 B 0.013584f
C496 VDD1.n169 B 0.012829f
C497 VDD1.n170 B 0.023875f
C498 VDD1.n171 B 0.023875f
C499 VDD1.n172 B 0.012829f
C500 VDD1.n173 B 0.013584f
C501 VDD1.n174 B 0.030323f
C502 VDD1.n175 B 0.030323f
C503 VDD1.n176 B 0.013584f
C504 VDD1.n177 B 0.012829f
C505 VDD1.n178 B 0.023875f
C506 VDD1.n179 B 0.023875f
C507 VDD1.n180 B 0.012829f
C508 VDD1.n181 B 0.013584f
C509 VDD1.n182 B 0.030323f
C510 VDD1.n183 B 0.030323f
C511 VDD1.n184 B 0.013584f
C512 VDD1.n185 B 0.012829f
C513 VDD1.n186 B 0.023875f
C514 VDD1.n187 B 0.062686f
C515 VDD1.n188 B 0.012829f
C516 VDD1.n189 B 0.013584f
C517 VDD1.n190 B 0.060803f
C518 VDD1.n191 B 0.082428f
C519 VDD1.t2 B 0.328087f
C520 VDD1.t5 B 0.328087f
C521 VDD1.n192 B 2.99516f
C522 VDD1.n193 B 0.706518f
C523 VDD1.t4 B 0.328087f
C524 VDD1.t6 B 0.328087f
C525 VDD1.n194 B 3.01287f
C526 VDD1.n195 B 3.38985f
C527 VDD1.t7 B 0.328087f
C528 VDD1.t9 B 0.328087f
C529 VDD1.n196 B 2.99515f
C530 VDD1.n197 B 3.54466f
C531 VTAIL.t8 B 0.328148f
C532 VTAIL.t1 B 0.328148f
C533 VTAIL.n0 B 2.93195f
C534 VTAIL.n1 B 0.530488f
C535 VTAIL.n2 B 0.013479f
C536 VTAIL.n3 B 0.030329f
C537 VTAIL.n4 B 0.013586f
C538 VTAIL.n5 B 0.023879f
C539 VTAIL.n6 B 0.012832f
C540 VTAIL.n7 B 0.030329f
C541 VTAIL.n8 B 0.013586f
C542 VTAIL.n9 B 0.023879f
C543 VTAIL.n10 B 0.012832f
C544 VTAIL.n11 B 0.030329f
C545 VTAIL.n12 B 0.013586f
C546 VTAIL.n13 B 0.023879f
C547 VTAIL.n14 B 0.012832f
C548 VTAIL.n15 B 0.030329f
C549 VTAIL.n16 B 0.013586f
C550 VTAIL.n17 B 0.023879f
C551 VTAIL.n18 B 0.012832f
C552 VTAIL.n19 B 0.030329f
C553 VTAIL.n20 B 0.013586f
C554 VTAIL.n21 B 0.023879f
C555 VTAIL.n22 B 0.013209f
C556 VTAIL.n23 B 0.030329f
C557 VTAIL.n24 B 0.013586f
C558 VTAIL.n25 B 0.023879f
C559 VTAIL.n26 B 0.012832f
C560 VTAIL.n27 B 0.030329f
C561 VTAIL.n28 B 0.013586f
C562 VTAIL.n29 B 0.023879f
C563 VTAIL.n30 B 0.012832f
C564 VTAIL.n31 B 0.022747f
C565 VTAIL.n32 B 0.02144f
C566 VTAIL.t10 B 0.051917f
C567 VTAIL.n33 B 0.221578f
C568 VTAIL.n34 B 1.77713f
C569 VTAIL.n35 B 0.012832f
C570 VTAIL.n36 B 0.013586f
C571 VTAIL.n37 B 0.030329f
C572 VTAIL.n38 B 0.030329f
C573 VTAIL.n39 B 0.013586f
C574 VTAIL.n40 B 0.012832f
C575 VTAIL.n41 B 0.023879f
C576 VTAIL.n42 B 0.023879f
C577 VTAIL.n43 B 0.012832f
C578 VTAIL.n44 B 0.013586f
C579 VTAIL.n45 B 0.030329f
C580 VTAIL.n46 B 0.030329f
C581 VTAIL.n47 B 0.013586f
C582 VTAIL.n48 B 0.012832f
C583 VTAIL.n49 B 0.023879f
C584 VTAIL.n50 B 0.023879f
C585 VTAIL.n51 B 0.012832f
C586 VTAIL.n52 B 0.012832f
C587 VTAIL.n53 B 0.013586f
C588 VTAIL.n54 B 0.030329f
C589 VTAIL.n55 B 0.030329f
C590 VTAIL.n56 B 0.030329f
C591 VTAIL.n57 B 0.013209f
C592 VTAIL.n58 B 0.012832f
C593 VTAIL.n59 B 0.023879f
C594 VTAIL.n60 B 0.023879f
C595 VTAIL.n61 B 0.012832f
C596 VTAIL.n62 B 0.013586f
C597 VTAIL.n63 B 0.030329f
C598 VTAIL.n64 B 0.030329f
C599 VTAIL.n65 B 0.013586f
C600 VTAIL.n66 B 0.012832f
C601 VTAIL.n67 B 0.023879f
C602 VTAIL.n68 B 0.023879f
C603 VTAIL.n69 B 0.012832f
C604 VTAIL.n70 B 0.013586f
C605 VTAIL.n71 B 0.030329f
C606 VTAIL.n72 B 0.030329f
C607 VTAIL.n73 B 0.013586f
C608 VTAIL.n74 B 0.012832f
C609 VTAIL.n75 B 0.023879f
C610 VTAIL.n76 B 0.023879f
C611 VTAIL.n77 B 0.012832f
C612 VTAIL.n78 B 0.013586f
C613 VTAIL.n79 B 0.030329f
C614 VTAIL.n80 B 0.030329f
C615 VTAIL.n81 B 0.013586f
C616 VTAIL.n82 B 0.012832f
C617 VTAIL.n83 B 0.023879f
C618 VTAIL.n84 B 0.023879f
C619 VTAIL.n85 B 0.012832f
C620 VTAIL.n86 B 0.013586f
C621 VTAIL.n87 B 0.030329f
C622 VTAIL.n88 B 0.030329f
C623 VTAIL.n89 B 0.013586f
C624 VTAIL.n90 B 0.012832f
C625 VTAIL.n91 B 0.023879f
C626 VTAIL.n92 B 0.062698f
C627 VTAIL.n93 B 0.012832f
C628 VTAIL.n94 B 0.013586f
C629 VTAIL.n95 B 0.060814f
C630 VTAIL.n96 B 0.052189f
C631 VTAIL.n97 B 0.384294f
C632 VTAIL.t9 B 0.328148f
C633 VTAIL.t16 B 0.328148f
C634 VTAIL.n98 B 2.93195f
C635 VTAIL.n99 B 0.652537f
C636 VTAIL.t12 B 0.328148f
C637 VTAIL.t18 B 0.328148f
C638 VTAIL.n100 B 2.93195f
C639 VTAIL.n101 B 2.3473f
C640 VTAIL.t7 B 0.328148f
C641 VTAIL.t2 B 0.328148f
C642 VTAIL.n102 B 2.93194f
C643 VTAIL.n103 B 2.3473f
C644 VTAIL.t4 B 0.328148f
C645 VTAIL.t19 B 0.328148f
C646 VTAIL.n104 B 2.93194f
C647 VTAIL.n105 B 0.652546f
C648 VTAIL.n106 B 0.013479f
C649 VTAIL.n107 B 0.030329f
C650 VTAIL.n108 B 0.013586f
C651 VTAIL.n109 B 0.023879f
C652 VTAIL.n110 B 0.012832f
C653 VTAIL.n111 B 0.030329f
C654 VTAIL.n112 B 0.013586f
C655 VTAIL.n113 B 0.023879f
C656 VTAIL.n114 B 0.012832f
C657 VTAIL.n115 B 0.030329f
C658 VTAIL.n116 B 0.013586f
C659 VTAIL.n117 B 0.023879f
C660 VTAIL.n118 B 0.012832f
C661 VTAIL.n119 B 0.030329f
C662 VTAIL.n120 B 0.013586f
C663 VTAIL.n121 B 0.023879f
C664 VTAIL.n122 B 0.012832f
C665 VTAIL.n123 B 0.030329f
C666 VTAIL.n124 B 0.013586f
C667 VTAIL.n125 B 0.023879f
C668 VTAIL.n126 B 0.013209f
C669 VTAIL.n127 B 0.030329f
C670 VTAIL.n128 B 0.012832f
C671 VTAIL.n129 B 0.013586f
C672 VTAIL.n130 B 0.023879f
C673 VTAIL.n131 B 0.012832f
C674 VTAIL.n132 B 0.030329f
C675 VTAIL.n133 B 0.013586f
C676 VTAIL.n134 B 0.023879f
C677 VTAIL.n135 B 0.012832f
C678 VTAIL.n136 B 0.022747f
C679 VTAIL.n137 B 0.02144f
C680 VTAIL.t3 B 0.051917f
C681 VTAIL.n138 B 0.221578f
C682 VTAIL.n139 B 1.77713f
C683 VTAIL.n140 B 0.012832f
C684 VTAIL.n141 B 0.013586f
C685 VTAIL.n142 B 0.030329f
C686 VTAIL.n143 B 0.030329f
C687 VTAIL.n144 B 0.013586f
C688 VTAIL.n145 B 0.012832f
C689 VTAIL.n146 B 0.023879f
C690 VTAIL.n147 B 0.023879f
C691 VTAIL.n148 B 0.012832f
C692 VTAIL.n149 B 0.013586f
C693 VTAIL.n150 B 0.030329f
C694 VTAIL.n151 B 0.030329f
C695 VTAIL.n152 B 0.013586f
C696 VTAIL.n153 B 0.012832f
C697 VTAIL.n154 B 0.023879f
C698 VTAIL.n155 B 0.023879f
C699 VTAIL.n156 B 0.012832f
C700 VTAIL.n157 B 0.013586f
C701 VTAIL.n158 B 0.030329f
C702 VTAIL.n159 B 0.030329f
C703 VTAIL.n160 B 0.030329f
C704 VTAIL.n161 B 0.013209f
C705 VTAIL.n162 B 0.012832f
C706 VTAIL.n163 B 0.023879f
C707 VTAIL.n164 B 0.023879f
C708 VTAIL.n165 B 0.012832f
C709 VTAIL.n166 B 0.013586f
C710 VTAIL.n167 B 0.030329f
C711 VTAIL.n168 B 0.030329f
C712 VTAIL.n169 B 0.013586f
C713 VTAIL.n170 B 0.012832f
C714 VTAIL.n171 B 0.023879f
C715 VTAIL.n172 B 0.023879f
C716 VTAIL.n173 B 0.012832f
C717 VTAIL.n174 B 0.013586f
C718 VTAIL.n175 B 0.030329f
C719 VTAIL.n176 B 0.030329f
C720 VTAIL.n177 B 0.013586f
C721 VTAIL.n178 B 0.012832f
C722 VTAIL.n179 B 0.023879f
C723 VTAIL.n180 B 0.023879f
C724 VTAIL.n181 B 0.012832f
C725 VTAIL.n182 B 0.013586f
C726 VTAIL.n183 B 0.030329f
C727 VTAIL.n184 B 0.030329f
C728 VTAIL.n185 B 0.013586f
C729 VTAIL.n186 B 0.012832f
C730 VTAIL.n187 B 0.023879f
C731 VTAIL.n188 B 0.023879f
C732 VTAIL.n189 B 0.012832f
C733 VTAIL.n190 B 0.013586f
C734 VTAIL.n191 B 0.030329f
C735 VTAIL.n192 B 0.030329f
C736 VTAIL.n193 B 0.013586f
C737 VTAIL.n194 B 0.012832f
C738 VTAIL.n195 B 0.023879f
C739 VTAIL.n196 B 0.062698f
C740 VTAIL.n197 B 0.012832f
C741 VTAIL.n198 B 0.013586f
C742 VTAIL.n199 B 0.060814f
C743 VTAIL.n200 B 0.052189f
C744 VTAIL.n201 B 0.384294f
C745 VTAIL.t14 B 0.328148f
C746 VTAIL.t13 B 0.328148f
C747 VTAIL.n202 B 2.93194f
C748 VTAIL.n203 B 0.580245f
C749 VTAIL.t11 B 0.328148f
C750 VTAIL.t17 B 0.328148f
C751 VTAIL.n204 B 2.93194f
C752 VTAIL.n205 B 0.652546f
C753 VTAIL.n206 B 0.013479f
C754 VTAIL.n207 B 0.030329f
C755 VTAIL.n208 B 0.013586f
C756 VTAIL.n209 B 0.023879f
C757 VTAIL.n210 B 0.012832f
C758 VTAIL.n211 B 0.030329f
C759 VTAIL.n212 B 0.013586f
C760 VTAIL.n213 B 0.023879f
C761 VTAIL.n214 B 0.012832f
C762 VTAIL.n215 B 0.030329f
C763 VTAIL.n216 B 0.013586f
C764 VTAIL.n217 B 0.023879f
C765 VTAIL.n218 B 0.012832f
C766 VTAIL.n219 B 0.030329f
C767 VTAIL.n220 B 0.013586f
C768 VTAIL.n221 B 0.023879f
C769 VTAIL.n222 B 0.012832f
C770 VTAIL.n223 B 0.030329f
C771 VTAIL.n224 B 0.013586f
C772 VTAIL.n225 B 0.023879f
C773 VTAIL.n226 B 0.013209f
C774 VTAIL.n227 B 0.030329f
C775 VTAIL.n228 B 0.012832f
C776 VTAIL.n229 B 0.013586f
C777 VTAIL.n230 B 0.023879f
C778 VTAIL.n231 B 0.012832f
C779 VTAIL.n232 B 0.030329f
C780 VTAIL.n233 B 0.013586f
C781 VTAIL.n234 B 0.023879f
C782 VTAIL.n235 B 0.012832f
C783 VTAIL.n236 B 0.022747f
C784 VTAIL.n237 B 0.02144f
C785 VTAIL.t15 B 0.051917f
C786 VTAIL.n238 B 0.221578f
C787 VTAIL.n239 B 1.77713f
C788 VTAIL.n240 B 0.012832f
C789 VTAIL.n241 B 0.013586f
C790 VTAIL.n242 B 0.030329f
C791 VTAIL.n243 B 0.030329f
C792 VTAIL.n244 B 0.013586f
C793 VTAIL.n245 B 0.012832f
C794 VTAIL.n246 B 0.023879f
C795 VTAIL.n247 B 0.023879f
C796 VTAIL.n248 B 0.012832f
C797 VTAIL.n249 B 0.013586f
C798 VTAIL.n250 B 0.030329f
C799 VTAIL.n251 B 0.030329f
C800 VTAIL.n252 B 0.013586f
C801 VTAIL.n253 B 0.012832f
C802 VTAIL.n254 B 0.023879f
C803 VTAIL.n255 B 0.023879f
C804 VTAIL.n256 B 0.012832f
C805 VTAIL.n257 B 0.013586f
C806 VTAIL.n258 B 0.030329f
C807 VTAIL.n259 B 0.030329f
C808 VTAIL.n260 B 0.030329f
C809 VTAIL.n261 B 0.013209f
C810 VTAIL.n262 B 0.012832f
C811 VTAIL.n263 B 0.023879f
C812 VTAIL.n264 B 0.023879f
C813 VTAIL.n265 B 0.012832f
C814 VTAIL.n266 B 0.013586f
C815 VTAIL.n267 B 0.030329f
C816 VTAIL.n268 B 0.030329f
C817 VTAIL.n269 B 0.013586f
C818 VTAIL.n270 B 0.012832f
C819 VTAIL.n271 B 0.023879f
C820 VTAIL.n272 B 0.023879f
C821 VTAIL.n273 B 0.012832f
C822 VTAIL.n274 B 0.013586f
C823 VTAIL.n275 B 0.030329f
C824 VTAIL.n276 B 0.030329f
C825 VTAIL.n277 B 0.013586f
C826 VTAIL.n278 B 0.012832f
C827 VTAIL.n279 B 0.023879f
C828 VTAIL.n280 B 0.023879f
C829 VTAIL.n281 B 0.012832f
C830 VTAIL.n282 B 0.013586f
C831 VTAIL.n283 B 0.030329f
C832 VTAIL.n284 B 0.030329f
C833 VTAIL.n285 B 0.013586f
C834 VTAIL.n286 B 0.012832f
C835 VTAIL.n287 B 0.023879f
C836 VTAIL.n288 B 0.023879f
C837 VTAIL.n289 B 0.012832f
C838 VTAIL.n290 B 0.013586f
C839 VTAIL.n291 B 0.030329f
C840 VTAIL.n292 B 0.030329f
C841 VTAIL.n293 B 0.013586f
C842 VTAIL.n294 B 0.012832f
C843 VTAIL.n295 B 0.023879f
C844 VTAIL.n296 B 0.062698f
C845 VTAIL.n297 B 0.012832f
C846 VTAIL.n298 B 0.013586f
C847 VTAIL.n299 B 0.060814f
C848 VTAIL.n300 B 0.052189f
C849 VTAIL.n301 B 1.93445f
C850 VTAIL.n302 B 0.013479f
C851 VTAIL.n303 B 0.030329f
C852 VTAIL.n304 B 0.013586f
C853 VTAIL.n305 B 0.023879f
C854 VTAIL.n306 B 0.012832f
C855 VTAIL.n307 B 0.030329f
C856 VTAIL.n308 B 0.013586f
C857 VTAIL.n309 B 0.023879f
C858 VTAIL.n310 B 0.012832f
C859 VTAIL.n311 B 0.030329f
C860 VTAIL.n312 B 0.013586f
C861 VTAIL.n313 B 0.023879f
C862 VTAIL.n314 B 0.012832f
C863 VTAIL.n315 B 0.030329f
C864 VTAIL.n316 B 0.013586f
C865 VTAIL.n317 B 0.023879f
C866 VTAIL.n318 B 0.012832f
C867 VTAIL.n319 B 0.030329f
C868 VTAIL.n320 B 0.013586f
C869 VTAIL.n321 B 0.023879f
C870 VTAIL.n322 B 0.013209f
C871 VTAIL.n323 B 0.030329f
C872 VTAIL.n324 B 0.013586f
C873 VTAIL.n325 B 0.023879f
C874 VTAIL.n326 B 0.012832f
C875 VTAIL.n327 B 0.030329f
C876 VTAIL.n328 B 0.013586f
C877 VTAIL.n329 B 0.023879f
C878 VTAIL.n330 B 0.012832f
C879 VTAIL.n331 B 0.022747f
C880 VTAIL.n332 B 0.02144f
C881 VTAIL.t5 B 0.051917f
C882 VTAIL.n333 B 0.221578f
C883 VTAIL.n334 B 1.77713f
C884 VTAIL.n335 B 0.012832f
C885 VTAIL.n336 B 0.013586f
C886 VTAIL.n337 B 0.030329f
C887 VTAIL.n338 B 0.030329f
C888 VTAIL.n339 B 0.013586f
C889 VTAIL.n340 B 0.012832f
C890 VTAIL.n341 B 0.023879f
C891 VTAIL.n342 B 0.023879f
C892 VTAIL.n343 B 0.012832f
C893 VTAIL.n344 B 0.013586f
C894 VTAIL.n345 B 0.030329f
C895 VTAIL.n346 B 0.030329f
C896 VTAIL.n347 B 0.013586f
C897 VTAIL.n348 B 0.012832f
C898 VTAIL.n349 B 0.023879f
C899 VTAIL.n350 B 0.023879f
C900 VTAIL.n351 B 0.012832f
C901 VTAIL.n352 B 0.012832f
C902 VTAIL.n353 B 0.013586f
C903 VTAIL.n354 B 0.030329f
C904 VTAIL.n355 B 0.030329f
C905 VTAIL.n356 B 0.030329f
C906 VTAIL.n357 B 0.013209f
C907 VTAIL.n358 B 0.012832f
C908 VTAIL.n359 B 0.023879f
C909 VTAIL.n360 B 0.023879f
C910 VTAIL.n361 B 0.012832f
C911 VTAIL.n362 B 0.013586f
C912 VTAIL.n363 B 0.030329f
C913 VTAIL.n364 B 0.030329f
C914 VTAIL.n365 B 0.013586f
C915 VTAIL.n366 B 0.012832f
C916 VTAIL.n367 B 0.023879f
C917 VTAIL.n368 B 0.023879f
C918 VTAIL.n369 B 0.012832f
C919 VTAIL.n370 B 0.013586f
C920 VTAIL.n371 B 0.030329f
C921 VTAIL.n372 B 0.030329f
C922 VTAIL.n373 B 0.013586f
C923 VTAIL.n374 B 0.012832f
C924 VTAIL.n375 B 0.023879f
C925 VTAIL.n376 B 0.023879f
C926 VTAIL.n377 B 0.012832f
C927 VTAIL.n378 B 0.013586f
C928 VTAIL.n379 B 0.030329f
C929 VTAIL.n380 B 0.030329f
C930 VTAIL.n381 B 0.013586f
C931 VTAIL.n382 B 0.012832f
C932 VTAIL.n383 B 0.023879f
C933 VTAIL.n384 B 0.023879f
C934 VTAIL.n385 B 0.012832f
C935 VTAIL.n386 B 0.013586f
C936 VTAIL.n387 B 0.030329f
C937 VTAIL.n388 B 0.030329f
C938 VTAIL.n389 B 0.013586f
C939 VTAIL.n390 B 0.012832f
C940 VTAIL.n391 B 0.023879f
C941 VTAIL.n392 B 0.062698f
C942 VTAIL.n393 B 0.012832f
C943 VTAIL.n394 B 0.013586f
C944 VTAIL.n395 B 0.060814f
C945 VTAIL.n396 B 0.052189f
C946 VTAIL.n397 B 1.93445f
C947 VTAIL.t6 B 0.328148f
C948 VTAIL.t0 B 0.328148f
C949 VTAIL.n398 B 2.93195f
C950 VTAIL.n399 B 0.485384f
C951 VP.n0 B 0.025291f
C952 VP.t3 B 2.69584f
C953 VP.n1 B 0.038515f
C954 VP.n2 B 0.019183f
C955 VP.n3 B 0.02622f
C956 VP.n4 B 0.019183f
C957 VP.n5 B 0.020524f
C958 VP.n6 B 0.019183f
C959 VP.t4 B 2.69584f
C960 VP.n7 B 0.035752f
C961 VP.n8 B 0.019183f
C962 VP.n9 B 0.035752f
C963 VP.n10 B 0.019183f
C964 VP.t7 B 2.69584f
C965 VP.n11 B 0.035393f
C966 VP.n12 B 0.019183f
C967 VP.n13 B 0.019513f
C968 VP.n14 B 0.025291f
C969 VP.t0 B 2.69584f
C970 VP.n15 B 0.038515f
C971 VP.n16 B 0.019183f
C972 VP.n17 B 0.02622f
C973 VP.n18 B 0.019183f
C974 VP.n19 B 0.020524f
C975 VP.n20 B 0.019183f
C976 VP.t9 B 2.69584f
C977 VP.n21 B 0.035752f
C978 VP.n22 B 0.019183f
C979 VP.n23 B 0.035752f
C980 VP.t6 B 2.89454f
C981 VP.n24 B 0.965178f
C982 VP.t1 B 2.69584f
C983 VP.n25 B 0.994842f
C984 VP.n26 B 0.027632f
C985 VP.n27 B 0.204347f
C986 VP.n28 B 0.019183f
C987 VP.n29 B 0.019183f
C988 VP.n30 B 0.033833f
C989 VP.n31 B 0.020524f
C990 VP.n32 B 0.037405f
C991 VP.n33 B 0.019183f
C992 VP.n34 B 0.019183f
C993 VP.n35 B 0.019183f
C994 VP.n36 B 0.951925f
C995 VP.n37 B 0.035752f
C996 VP.n38 B 0.037405f
C997 VP.n39 B 0.019183f
C998 VP.n40 B 0.019183f
C999 VP.n41 B 0.019183f
C1000 VP.n42 B 0.033833f
C1001 VP.n43 B 0.035752f
C1002 VP.t2 B 2.69584f
C1003 VP.n44 B 0.933824f
C1004 VP.n45 B 0.027632f
C1005 VP.n46 B 0.019183f
C1006 VP.n47 B 0.019183f
C1007 VP.n48 B 0.019183f
C1008 VP.n49 B 0.035752f
C1009 VP.n50 B 0.035393f
C1010 VP.n51 B 0.017854f
C1011 VP.n52 B 0.019183f
C1012 VP.n53 B 0.019183f
C1013 VP.n54 B 0.019183f
C1014 VP.n55 B 0.035752f
C1015 VP.n56 B 0.019513f
C1016 VP.n57 B 0.998321f
C1017 VP.n58 B 1.35645f
C1018 VP.t8 B 2.69584f
C1019 VP.n59 B 0.998321f
C1020 VP.n60 B 1.36814f
C1021 VP.n61 B 0.025291f
C1022 VP.n62 B 0.019183f
C1023 VP.n63 B 0.035752f
C1024 VP.n64 B 0.038515f
C1025 VP.n65 B 0.017854f
C1026 VP.n66 B 0.019183f
C1027 VP.n67 B 0.019183f
C1028 VP.n68 B 0.019183f
C1029 VP.n69 B 0.035752f
C1030 VP.n70 B 0.02622f
C1031 VP.n71 B 0.933824f
C1032 VP.n72 B 0.027632f
C1033 VP.n73 B 0.019183f
C1034 VP.n74 B 0.019183f
C1035 VP.n75 B 0.019183f
C1036 VP.n76 B 0.033833f
C1037 VP.n77 B 0.020524f
C1038 VP.n78 B 0.037405f
C1039 VP.n79 B 0.019183f
C1040 VP.n80 B 0.019183f
C1041 VP.n81 B 0.019183f
C1042 VP.n82 B 0.951925f
C1043 VP.n83 B 0.035752f
C1044 VP.n84 B 0.037405f
C1045 VP.n85 B 0.019183f
C1046 VP.n86 B 0.019183f
C1047 VP.n87 B 0.019183f
C1048 VP.n88 B 0.033833f
C1049 VP.n89 B 0.035752f
C1050 VP.t5 B 2.69584f
C1051 VP.n90 B 0.933824f
C1052 VP.n91 B 0.027632f
C1053 VP.n92 B 0.019183f
C1054 VP.n93 B 0.019183f
C1055 VP.n94 B 0.019183f
C1056 VP.n95 B 0.035752f
C1057 VP.n96 B 0.035393f
C1058 VP.n97 B 0.017854f
C1059 VP.n98 B 0.019183f
C1060 VP.n99 B 0.019183f
C1061 VP.n100 B 0.019183f
C1062 VP.n101 B 0.035752f
C1063 VP.n102 B 0.019513f
C1064 VP.n103 B 0.998321f
C1065 VP.n104 B 0.037253f
.ends

