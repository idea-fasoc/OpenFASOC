* NGSPICE file created from diff_pair_sample_0990.ext - technology: sky130A

.subckt diff_pair_sample_0990 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X1 VDD1.t4 VP.t1 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X2 VTAIL.t13 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X3 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=1.17315 ps=7.44 w=7.11 l=1.52
X4 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=0 ps=0 w=7.11 l=1.52
X6 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=2.7729 ps=15 w=7.11 l=1.52
X7 VTAIL.t12 VP.t3 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=1.17315 ps=7.44 w=7.11 l=1.52
X8 VTAIL.t11 VP.t4 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=1.17315 ps=7.44 w=7.11 l=1.52
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=0 ps=0 w=7.11 l=1.52
X10 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X11 VTAIL.t1 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=1.17315 ps=7.44 w=7.11 l=1.52
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=0 ps=0 w=7.11 l=1.52
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7729 pd=15 as=0 ps=0 w=7.11 l=1.52
X14 VDD2.t2 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=2.7729 ps=15 w=7.11 l=1.52
X15 VDD1.t5 VP.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=2.7729 ps=15 w=7.11 l=1.52
X16 VDD1.t1 VP.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=2.7729 ps=15 w=7.11 l=1.52
X17 VDD1.t2 VP.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X18 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
X19 VDD2.t0 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.17315 pd=7.44 as=1.17315 ps=7.44 w=7.11 l=1.52
R0 VP.n26 VP.n25 172.31
R1 VP.n46 VP.n45 172.31
R2 VP.n24 VP.n23 172.31
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n44 VP.n0 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n1 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n37 VP.n2 161.3
R15 VP.n36 VP.n35 161.3
R16 VP.n34 VP.n3 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n30 VP.n4 161.3
R19 VP.n29 VP.n28 161.3
R20 VP.n27 VP.n5 161.3
R21 VP.n11 VP.t4 148.417
R22 VP.n25 VP.t3 112.731
R23 VP.n31 VP.t1 112.731
R24 VP.n38 VP.t0 112.731
R25 VP.n45 VP.t6 112.731
R26 VP.n23 VP.t5 112.731
R27 VP.n16 VP.t2 112.731
R28 VP.n10 VP.t7 112.731
R29 VP.n30 VP.n29 55.0624
R30 VP.n43 VP.n1 55.0624
R31 VP.n21 VP.n7 55.0624
R32 VP.n11 VP.n10 45.8064
R33 VP.n26 VP.n24 42.1217
R34 VP.n36 VP.n3 40.4934
R35 VP.n37 VP.n36 40.4934
R36 VP.n15 VP.n14 40.4934
R37 VP.n14 VP.n9 40.4934
R38 VP.n29 VP.n5 25.9244
R39 VP.n44 VP.n43 25.9244
R40 VP.n22 VP.n21 25.9244
R41 VP.n32 VP.n30 24.4675
R42 VP.n39 VP.n1 24.4675
R43 VP.n17 VP.n7 24.4675
R44 VP.n31 VP.n3 20.7975
R45 VP.n38 VP.n37 20.7975
R46 VP.n16 VP.n15 20.7975
R47 VP.n10 VP.n9 20.7975
R48 VP.n12 VP.n11 17.4308
R49 VP.n25 VP.n5 13.4574
R50 VP.n45 VP.n44 13.4574
R51 VP.n23 VP.n22 13.4574
R52 VP.n32 VP.n31 3.67055
R53 VP.n39 VP.n38 3.67055
R54 VP.n17 VP.n16 3.67055
R55 VP.n13 VP.n12 0.189894
R56 VP.n13 VP.n8 0.189894
R57 VP.n18 VP.n8 0.189894
R58 VP.n19 VP.n18 0.189894
R59 VP.n20 VP.n19 0.189894
R60 VP.n20 VP.n6 0.189894
R61 VP.n24 VP.n6 0.189894
R62 VP.n27 VP.n26 0.189894
R63 VP.n28 VP.n27 0.189894
R64 VP.n28 VP.n4 0.189894
R65 VP.n33 VP.n4 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n35 VP.n34 0.189894
R68 VP.n35 VP.n2 0.189894
R69 VP.n40 VP.n2 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n42 VP.n41 0.189894
R72 VP.n42 VP.n0 0.189894
R73 VP.n46 VP.n0 0.189894
R74 VP VP.n46 0.0516364
R75 VDD1 VDD1.n0 67.0487
R76 VDD1.n3 VDD1.n2 66.9351
R77 VDD1.n3 VDD1.n1 66.9351
R78 VDD1.n5 VDD1.n4 66.1929
R79 VDD1.n5 VDD1.n3 37.6043
R80 VDD1.n4 VDD1.t3 2.78531
R81 VDD1.n4 VDD1.t5 2.78531
R82 VDD1.n0 VDD1.t6 2.78531
R83 VDD1.n0 VDD1.t2 2.78531
R84 VDD1.n2 VDD1.t0 2.78531
R85 VDD1.n2 VDD1.t1 2.78531
R86 VDD1.n1 VDD1.t7 2.78531
R87 VDD1.n1 VDD1.t4 2.78531
R88 VDD1 VDD1.n5 0.739724
R89 VTAIL.n11 VTAIL.t11 52.2991
R90 VTAIL.n10 VTAIL.t2 52.2991
R91 VTAIL.n7 VTAIL.t3 52.2991
R92 VTAIL.n15 VTAIL.t7 52.2989
R93 VTAIL.n2 VTAIL.t1 52.2989
R94 VTAIL.n3 VTAIL.t9 52.2989
R95 VTAIL.n6 VTAIL.t12 52.2989
R96 VTAIL.n14 VTAIL.t10 52.2989
R97 VTAIL.n13 VTAIL.n12 49.5143
R98 VTAIL.n9 VTAIL.n8 49.5143
R99 VTAIL.n1 VTAIL.n0 49.5142
R100 VTAIL.n5 VTAIL.n4 49.5142
R101 VTAIL.n15 VTAIL.n14 20.091
R102 VTAIL.n7 VTAIL.n6 20.091
R103 VTAIL.n0 VTAIL.t6 2.78531
R104 VTAIL.n0 VTAIL.t4 2.78531
R105 VTAIL.n4 VTAIL.t14 2.78531
R106 VTAIL.n4 VTAIL.t15 2.78531
R107 VTAIL.n12 VTAIL.t8 2.78531
R108 VTAIL.n12 VTAIL.t13 2.78531
R109 VTAIL.n8 VTAIL.t0 2.78531
R110 VTAIL.n8 VTAIL.t5 2.78531
R111 VTAIL.n9 VTAIL.n7 1.59533
R112 VTAIL.n10 VTAIL.n9 1.59533
R113 VTAIL.n13 VTAIL.n11 1.59533
R114 VTAIL.n14 VTAIL.n13 1.59533
R115 VTAIL.n6 VTAIL.n5 1.59533
R116 VTAIL.n5 VTAIL.n3 1.59533
R117 VTAIL.n2 VTAIL.n1 1.59533
R118 VTAIL VTAIL.n15 1.53714
R119 VTAIL.n11 VTAIL.n10 0.470328
R120 VTAIL.n3 VTAIL.n2 0.470328
R121 VTAIL VTAIL.n1 0.0586897
R122 B.n613 B.n612 585
R123 B.n226 B.n98 585
R124 B.n225 B.n224 585
R125 B.n223 B.n222 585
R126 B.n221 B.n220 585
R127 B.n219 B.n218 585
R128 B.n217 B.n216 585
R129 B.n215 B.n214 585
R130 B.n213 B.n212 585
R131 B.n211 B.n210 585
R132 B.n209 B.n208 585
R133 B.n207 B.n206 585
R134 B.n205 B.n204 585
R135 B.n203 B.n202 585
R136 B.n201 B.n200 585
R137 B.n199 B.n198 585
R138 B.n197 B.n196 585
R139 B.n195 B.n194 585
R140 B.n193 B.n192 585
R141 B.n191 B.n190 585
R142 B.n189 B.n188 585
R143 B.n187 B.n186 585
R144 B.n185 B.n184 585
R145 B.n183 B.n182 585
R146 B.n181 B.n180 585
R147 B.n179 B.n178 585
R148 B.n177 B.n176 585
R149 B.n174 B.n173 585
R150 B.n172 B.n171 585
R151 B.n170 B.n169 585
R152 B.n168 B.n167 585
R153 B.n166 B.n165 585
R154 B.n164 B.n163 585
R155 B.n162 B.n161 585
R156 B.n160 B.n159 585
R157 B.n158 B.n157 585
R158 B.n156 B.n155 585
R159 B.n153 B.n152 585
R160 B.n151 B.n150 585
R161 B.n149 B.n148 585
R162 B.n147 B.n146 585
R163 B.n145 B.n144 585
R164 B.n143 B.n142 585
R165 B.n141 B.n140 585
R166 B.n139 B.n138 585
R167 B.n137 B.n136 585
R168 B.n135 B.n134 585
R169 B.n133 B.n132 585
R170 B.n131 B.n130 585
R171 B.n129 B.n128 585
R172 B.n127 B.n126 585
R173 B.n125 B.n124 585
R174 B.n123 B.n122 585
R175 B.n121 B.n120 585
R176 B.n119 B.n118 585
R177 B.n117 B.n116 585
R178 B.n115 B.n114 585
R179 B.n113 B.n112 585
R180 B.n111 B.n110 585
R181 B.n109 B.n108 585
R182 B.n107 B.n106 585
R183 B.n105 B.n104 585
R184 B.n67 B.n66 585
R185 B.n618 B.n617 585
R186 B.n611 B.n99 585
R187 B.n99 B.n64 585
R188 B.n610 B.n63 585
R189 B.n622 B.n63 585
R190 B.n609 B.n62 585
R191 B.n623 B.n62 585
R192 B.n608 B.n61 585
R193 B.n624 B.n61 585
R194 B.n607 B.n606 585
R195 B.n606 B.n57 585
R196 B.n605 B.n56 585
R197 B.n630 B.n56 585
R198 B.n604 B.n55 585
R199 B.n631 B.n55 585
R200 B.n603 B.n54 585
R201 B.n632 B.n54 585
R202 B.n602 B.n601 585
R203 B.n601 B.n50 585
R204 B.n600 B.n49 585
R205 B.n638 B.n49 585
R206 B.n599 B.n48 585
R207 B.n639 B.n48 585
R208 B.n598 B.n47 585
R209 B.n640 B.n47 585
R210 B.n597 B.n596 585
R211 B.n596 B.n43 585
R212 B.n595 B.n42 585
R213 B.n646 B.n42 585
R214 B.n594 B.n41 585
R215 B.n647 B.n41 585
R216 B.n593 B.n40 585
R217 B.n648 B.n40 585
R218 B.n592 B.n591 585
R219 B.n591 B.n36 585
R220 B.n590 B.n35 585
R221 B.n654 B.n35 585
R222 B.n589 B.n34 585
R223 B.n655 B.n34 585
R224 B.n588 B.n33 585
R225 B.n656 B.n33 585
R226 B.n587 B.n586 585
R227 B.n586 B.n32 585
R228 B.n585 B.n28 585
R229 B.n662 B.n28 585
R230 B.n584 B.n27 585
R231 B.n663 B.n27 585
R232 B.n583 B.n26 585
R233 B.n664 B.n26 585
R234 B.n582 B.n581 585
R235 B.n581 B.n22 585
R236 B.n580 B.n21 585
R237 B.n670 B.n21 585
R238 B.n579 B.n20 585
R239 B.n671 B.n20 585
R240 B.n578 B.n19 585
R241 B.n672 B.n19 585
R242 B.n577 B.n576 585
R243 B.n576 B.n15 585
R244 B.n575 B.n14 585
R245 B.n678 B.n14 585
R246 B.n574 B.n13 585
R247 B.n679 B.n13 585
R248 B.n573 B.n12 585
R249 B.n680 B.n12 585
R250 B.n572 B.n571 585
R251 B.n571 B.n570 585
R252 B.n569 B.n568 585
R253 B.n569 B.n8 585
R254 B.n567 B.n7 585
R255 B.n687 B.n7 585
R256 B.n566 B.n6 585
R257 B.n688 B.n6 585
R258 B.n565 B.n5 585
R259 B.n689 B.n5 585
R260 B.n564 B.n563 585
R261 B.n563 B.n4 585
R262 B.n562 B.n227 585
R263 B.n562 B.n561 585
R264 B.n552 B.n228 585
R265 B.n229 B.n228 585
R266 B.n554 B.n553 585
R267 B.n555 B.n554 585
R268 B.n551 B.n234 585
R269 B.n234 B.n233 585
R270 B.n550 B.n549 585
R271 B.n549 B.n548 585
R272 B.n236 B.n235 585
R273 B.n237 B.n236 585
R274 B.n541 B.n540 585
R275 B.n542 B.n541 585
R276 B.n539 B.n242 585
R277 B.n242 B.n241 585
R278 B.n538 B.n537 585
R279 B.n537 B.n536 585
R280 B.n244 B.n243 585
R281 B.n245 B.n244 585
R282 B.n529 B.n528 585
R283 B.n530 B.n529 585
R284 B.n527 B.n250 585
R285 B.n250 B.n249 585
R286 B.n526 B.n525 585
R287 B.n525 B.n524 585
R288 B.n252 B.n251 585
R289 B.n517 B.n252 585
R290 B.n516 B.n515 585
R291 B.n518 B.n516 585
R292 B.n514 B.n257 585
R293 B.n257 B.n256 585
R294 B.n513 B.n512 585
R295 B.n512 B.n511 585
R296 B.n259 B.n258 585
R297 B.n260 B.n259 585
R298 B.n504 B.n503 585
R299 B.n505 B.n504 585
R300 B.n502 B.n264 585
R301 B.n268 B.n264 585
R302 B.n501 B.n500 585
R303 B.n500 B.n499 585
R304 B.n266 B.n265 585
R305 B.n267 B.n266 585
R306 B.n492 B.n491 585
R307 B.n493 B.n492 585
R308 B.n490 B.n273 585
R309 B.n273 B.n272 585
R310 B.n489 B.n488 585
R311 B.n488 B.n487 585
R312 B.n275 B.n274 585
R313 B.n276 B.n275 585
R314 B.n480 B.n479 585
R315 B.n481 B.n480 585
R316 B.n478 B.n280 585
R317 B.n284 B.n280 585
R318 B.n477 B.n476 585
R319 B.n476 B.n475 585
R320 B.n282 B.n281 585
R321 B.n283 B.n282 585
R322 B.n468 B.n467 585
R323 B.n469 B.n468 585
R324 B.n466 B.n289 585
R325 B.n289 B.n288 585
R326 B.n465 B.n464 585
R327 B.n464 B.n463 585
R328 B.n291 B.n290 585
R329 B.n292 B.n291 585
R330 B.n459 B.n458 585
R331 B.n295 B.n294 585
R332 B.n455 B.n454 585
R333 B.n456 B.n455 585
R334 B.n453 B.n327 585
R335 B.n452 B.n451 585
R336 B.n450 B.n449 585
R337 B.n448 B.n447 585
R338 B.n446 B.n445 585
R339 B.n444 B.n443 585
R340 B.n442 B.n441 585
R341 B.n440 B.n439 585
R342 B.n438 B.n437 585
R343 B.n436 B.n435 585
R344 B.n434 B.n433 585
R345 B.n432 B.n431 585
R346 B.n430 B.n429 585
R347 B.n428 B.n427 585
R348 B.n426 B.n425 585
R349 B.n424 B.n423 585
R350 B.n422 B.n421 585
R351 B.n420 B.n419 585
R352 B.n418 B.n417 585
R353 B.n416 B.n415 585
R354 B.n414 B.n413 585
R355 B.n412 B.n411 585
R356 B.n410 B.n409 585
R357 B.n408 B.n407 585
R358 B.n406 B.n405 585
R359 B.n404 B.n403 585
R360 B.n402 B.n401 585
R361 B.n400 B.n399 585
R362 B.n398 B.n397 585
R363 B.n396 B.n395 585
R364 B.n394 B.n393 585
R365 B.n392 B.n391 585
R366 B.n390 B.n389 585
R367 B.n388 B.n387 585
R368 B.n386 B.n385 585
R369 B.n384 B.n383 585
R370 B.n382 B.n381 585
R371 B.n380 B.n379 585
R372 B.n378 B.n377 585
R373 B.n376 B.n375 585
R374 B.n374 B.n373 585
R375 B.n372 B.n371 585
R376 B.n370 B.n369 585
R377 B.n368 B.n367 585
R378 B.n366 B.n365 585
R379 B.n364 B.n363 585
R380 B.n362 B.n361 585
R381 B.n360 B.n359 585
R382 B.n358 B.n357 585
R383 B.n356 B.n355 585
R384 B.n354 B.n353 585
R385 B.n352 B.n351 585
R386 B.n350 B.n349 585
R387 B.n348 B.n347 585
R388 B.n346 B.n345 585
R389 B.n344 B.n343 585
R390 B.n342 B.n341 585
R391 B.n340 B.n339 585
R392 B.n338 B.n337 585
R393 B.n336 B.n335 585
R394 B.n334 B.n326 585
R395 B.n456 B.n326 585
R396 B.n460 B.n293 585
R397 B.n293 B.n292 585
R398 B.n462 B.n461 585
R399 B.n463 B.n462 585
R400 B.n287 B.n286 585
R401 B.n288 B.n287 585
R402 B.n471 B.n470 585
R403 B.n470 B.n469 585
R404 B.n472 B.n285 585
R405 B.n285 B.n283 585
R406 B.n474 B.n473 585
R407 B.n475 B.n474 585
R408 B.n279 B.n278 585
R409 B.n284 B.n279 585
R410 B.n483 B.n482 585
R411 B.n482 B.n481 585
R412 B.n484 B.n277 585
R413 B.n277 B.n276 585
R414 B.n486 B.n485 585
R415 B.n487 B.n486 585
R416 B.n271 B.n270 585
R417 B.n272 B.n271 585
R418 B.n495 B.n494 585
R419 B.n494 B.n493 585
R420 B.n496 B.n269 585
R421 B.n269 B.n267 585
R422 B.n498 B.n497 585
R423 B.n499 B.n498 585
R424 B.n263 B.n262 585
R425 B.n268 B.n263 585
R426 B.n507 B.n506 585
R427 B.n506 B.n505 585
R428 B.n508 B.n261 585
R429 B.n261 B.n260 585
R430 B.n510 B.n509 585
R431 B.n511 B.n510 585
R432 B.n255 B.n254 585
R433 B.n256 B.n255 585
R434 B.n520 B.n519 585
R435 B.n519 B.n518 585
R436 B.n521 B.n253 585
R437 B.n517 B.n253 585
R438 B.n523 B.n522 585
R439 B.n524 B.n523 585
R440 B.n248 B.n247 585
R441 B.n249 B.n248 585
R442 B.n532 B.n531 585
R443 B.n531 B.n530 585
R444 B.n533 B.n246 585
R445 B.n246 B.n245 585
R446 B.n535 B.n534 585
R447 B.n536 B.n535 585
R448 B.n240 B.n239 585
R449 B.n241 B.n240 585
R450 B.n544 B.n543 585
R451 B.n543 B.n542 585
R452 B.n545 B.n238 585
R453 B.n238 B.n237 585
R454 B.n547 B.n546 585
R455 B.n548 B.n547 585
R456 B.n232 B.n231 585
R457 B.n233 B.n232 585
R458 B.n557 B.n556 585
R459 B.n556 B.n555 585
R460 B.n558 B.n230 585
R461 B.n230 B.n229 585
R462 B.n560 B.n559 585
R463 B.n561 B.n560 585
R464 B.n3 B.n0 585
R465 B.n4 B.n3 585
R466 B.n686 B.n1 585
R467 B.n687 B.n686 585
R468 B.n685 B.n684 585
R469 B.n685 B.n8 585
R470 B.n683 B.n9 585
R471 B.n570 B.n9 585
R472 B.n682 B.n681 585
R473 B.n681 B.n680 585
R474 B.n11 B.n10 585
R475 B.n679 B.n11 585
R476 B.n677 B.n676 585
R477 B.n678 B.n677 585
R478 B.n675 B.n16 585
R479 B.n16 B.n15 585
R480 B.n674 B.n673 585
R481 B.n673 B.n672 585
R482 B.n18 B.n17 585
R483 B.n671 B.n18 585
R484 B.n669 B.n668 585
R485 B.n670 B.n669 585
R486 B.n667 B.n23 585
R487 B.n23 B.n22 585
R488 B.n666 B.n665 585
R489 B.n665 B.n664 585
R490 B.n25 B.n24 585
R491 B.n663 B.n25 585
R492 B.n661 B.n660 585
R493 B.n662 B.n661 585
R494 B.n659 B.n29 585
R495 B.n32 B.n29 585
R496 B.n658 B.n657 585
R497 B.n657 B.n656 585
R498 B.n31 B.n30 585
R499 B.n655 B.n31 585
R500 B.n653 B.n652 585
R501 B.n654 B.n653 585
R502 B.n651 B.n37 585
R503 B.n37 B.n36 585
R504 B.n650 B.n649 585
R505 B.n649 B.n648 585
R506 B.n39 B.n38 585
R507 B.n647 B.n39 585
R508 B.n645 B.n644 585
R509 B.n646 B.n645 585
R510 B.n643 B.n44 585
R511 B.n44 B.n43 585
R512 B.n642 B.n641 585
R513 B.n641 B.n640 585
R514 B.n46 B.n45 585
R515 B.n639 B.n46 585
R516 B.n637 B.n636 585
R517 B.n638 B.n637 585
R518 B.n635 B.n51 585
R519 B.n51 B.n50 585
R520 B.n634 B.n633 585
R521 B.n633 B.n632 585
R522 B.n53 B.n52 585
R523 B.n631 B.n53 585
R524 B.n629 B.n628 585
R525 B.n630 B.n629 585
R526 B.n627 B.n58 585
R527 B.n58 B.n57 585
R528 B.n626 B.n625 585
R529 B.n625 B.n624 585
R530 B.n60 B.n59 585
R531 B.n623 B.n60 585
R532 B.n621 B.n620 585
R533 B.n622 B.n621 585
R534 B.n619 B.n65 585
R535 B.n65 B.n64 585
R536 B.n690 B.n689 585
R537 B.n688 B.n2 585
R538 B.n617 B.n65 473.281
R539 B.n613 B.n99 473.281
R540 B.n326 B.n291 473.281
R541 B.n458 B.n293 473.281
R542 B.n102 B.t12 318.245
R543 B.n100 B.t16 318.245
R544 B.n331 B.t8 318.245
R545 B.n328 B.t19 318.245
R546 B.n615 B.n614 256.663
R547 B.n615 B.n97 256.663
R548 B.n615 B.n96 256.663
R549 B.n615 B.n95 256.663
R550 B.n615 B.n94 256.663
R551 B.n615 B.n93 256.663
R552 B.n615 B.n92 256.663
R553 B.n615 B.n91 256.663
R554 B.n615 B.n90 256.663
R555 B.n615 B.n89 256.663
R556 B.n615 B.n88 256.663
R557 B.n615 B.n87 256.663
R558 B.n615 B.n86 256.663
R559 B.n615 B.n85 256.663
R560 B.n615 B.n84 256.663
R561 B.n615 B.n83 256.663
R562 B.n615 B.n82 256.663
R563 B.n615 B.n81 256.663
R564 B.n615 B.n80 256.663
R565 B.n615 B.n79 256.663
R566 B.n615 B.n78 256.663
R567 B.n615 B.n77 256.663
R568 B.n615 B.n76 256.663
R569 B.n615 B.n75 256.663
R570 B.n615 B.n74 256.663
R571 B.n615 B.n73 256.663
R572 B.n615 B.n72 256.663
R573 B.n615 B.n71 256.663
R574 B.n615 B.n70 256.663
R575 B.n615 B.n69 256.663
R576 B.n615 B.n68 256.663
R577 B.n616 B.n615 256.663
R578 B.n457 B.n456 256.663
R579 B.n456 B.n296 256.663
R580 B.n456 B.n297 256.663
R581 B.n456 B.n298 256.663
R582 B.n456 B.n299 256.663
R583 B.n456 B.n300 256.663
R584 B.n456 B.n301 256.663
R585 B.n456 B.n302 256.663
R586 B.n456 B.n303 256.663
R587 B.n456 B.n304 256.663
R588 B.n456 B.n305 256.663
R589 B.n456 B.n306 256.663
R590 B.n456 B.n307 256.663
R591 B.n456 B.n308 256.663
R592 B.n456 B.n309 256.663
R593 B.n456 B.n310 256.663
R594 B.n456 B.n311 256.663
R595 B.n456 B.n312 256.663
R596 B.n456 B.n313 256.663
R597 B.n456 B.n314 256.663
R598 B.n456 B.n315 256.663
R599 B.n456 B.n316 256.663
R600 B.n456 B.n317 256.663
R601 B.n456 B.n318 256.663
R602 B.n456 B.n319 256.663
R603 B.n456 B.n320 256.663
R604 B.n456 B.n321 256.663
R605 B.n456 B.n322 256.663
R606 B.n456 B.n323 256.663
R607 B.n456 B.n324 256.663
R608 B.n456 B.n325 256.663
R609 B.n692 B.n691 256.663
R610 B.n104 B.n67 163.367
R611 B.n108 B.n107 163.367
R612 B.n112 B.n111 163.367
R613 B.n116 B.n115 163.367
R614 B.n120 B.n119 163.367
R615 B.n124 B.n123 163.367
R616 B.n128 B.n127 163.367
R617 B.n132 B.n131 163.367
R618 B.n136 B.n135 163.367
R619 B.n140 B.n139 163.367
R620 B.n144 B.n143 163.367
R621 B.n148 B.n147 163.367
R622 B.n152 B.n151 163.367
R623 B.n157 B.n156 163.367
R624 B.n161 B.n160 163.367
R625 B.n165 B.n164 163.367
R626 B.n169 B.n168 163.367
R627 B.n173 B.n172 163.367
R628 B.n178 B.n177 163.367
R629 B.n182 B.n181 163.367
R630 B.n186 B.n185 163.367
R631 B.n190 B.n189 163.367
R632 B.n194 B.n193 163.367
R633 B.n198 B.n197 163.367
R634 B.n202 B.n201 163.367
R635 B.n206 B.n205 163.367
R636 B.n210 B.n209 163.367
R637 B.n214 B.n213 163.367
R638 B.n218 B.n217 163.367
R639 B.n222 B.n221 163.367
R640 B.n224 B.n98 163.367
R641 B.n464 B.n291 163.367
R642 B.n464 B.n289 163.367
R643 B.n468 B.n289 163.367
R644 B.n468 B.n282 163.367
R645 B.n476 B.n282 163.367
R646 B.n476 B.n280 163.367
R647 B.n480 B.n280 163.367
R648 B.n480 B.n275 163.367
R649 B.n488 B.n275 163.367
R650 B.n488 B.n273 163.367
R651 B.n492 B.n273 163.367
R652 B.n492 B.n266 163.367
R653 B.n500 B.n266 163.367
R654 B.n500 B.n264 163.367
R655 B.n504 B.n264 163.367
R656 B.n504 B.n259 163.367
R657 B.n512 B.n259 163.367
R658 B.n512 B.n257 163.367
R659 B.n516 B.n257 163.367
R660 B.n516 B.n252 163.367
R661 B.n525 B.n252 163.367
R662 B.n525 B.n250 163.367
R663 B.n529 B.n250 163.367
R664 B.n529 B.n244 163.367
R665 B.n537 B.n244 163.367
R666 B.n537 B.n242 163.367
R667 B.n541 B.n242 163.367
R668 B.n541 B.n236 163.367
R669 B.n549 B.n236 163.367
R670 B.n549 B.n234 163.367
R671 B.n554 B.n234 163.367
R672 B.n554 B.n228 163.367
R673 B.n562 B.n228 163.367
R674 B.n563 B.n562 163.367
R675 B.n563 B.n5 163.367
R676 B.n6 B.n5 163.367
R677 B.n7 B.n6 163.367
R678 B.n569 B.n7 163.367
R679 B.n571 B.n569 163.367
R680 B.n571 B.n12 163.367
R681 B.n13 B.n12 163.367
R682 B.n14 B.n13 163.367
R683 B.n576 B.n14 163.367
R684 B.n576 B.n19 163.367
R685 B.n20 B.n19 163.367
R686 B.n21 B.n20 163.367
R687 B.n581 B.n21 163.367
R688 B.n581 B.n26 163.367
R689 B.n27 B.n26 163.367
R690 B.n28 B.n27 163.367
R691 B.n586 B.n28 163.367
R692 B.n586 B.n33 163.367
R693 B.n34 B.n33 163.367
R694 B.n35 B.n34 163.367
R695 B.n591 B.n35 163.367
R696 B.n591 B.n40 163.367
R697 B.n41 B.n40 163.367
R698 B.n42 B.n41 163.367
R699 B.n596 B.n42 163.367
R700 B.n596 B.n47 163.367
R701 B.n48 B.n47 163.367
R702 B.n49 B.n48 163.367
R703 B.n601 B.n49 163.367
R704 B.n601 B.n54 163.367
R705 B.n55 B.n54 163.367
R706 B.n56 B.n55 163.367
R707 B.n606 B.n56 163.367
R708 B.n606 B.n61 163.367
R709 B.n62 B.n61 163.367
R710 B.n63 B.n62 163.367
R711 B.n99 B.n63 163.367
R712 B.n455 B.n295 163.367
R713 B.n455 B.n327 163.367
R714 B.n451 B.n450 163.367
R715 B.n447 B.n446 163.367
R716 B.n443 B.n442 163.367
R717 B.n439 B.n438 163.367
R718 B.n435 B.n434 163.367
R719 B.n431 B.n430 163.367
R720 B.n427 B.n426 163.367
R721 B.n423 B.n422 163.367
R722 B.n419 B.n418 163.367
R723 B.n415 B.n414 163.367
R724 B.n411 B.n410 163.367
R725 B.n407 B.n406 163.367
R726 B.n403 B.n402 163.367
R727 B.n399 B.n398 163.367
R728 B.n395 B.n394 163.367
R729 B.n391 B.n390 163.367
R730 B.n387 B.n386 163.367
R731 B.n383 B.n382 163.367
R732 B.n379 B.n378 163.367
R733 B.n375 B.n374 163.367
R734 B.n371 B.n370 163.367
R735 B.n367 B.n366 163.367
R736 B.n363 B.n362 163.367
R737 B.n359 B.n358 163.367
R738 B.n355 B.n354 163.367
R739 B.n351 B.n350 163.367
R740 B.n347 B.n346 163.367
R741 B.n343 B.n342 163.367
R742 B.n339 B.n338 163.367
R743 B.n335 B.n326 163.367
R744 B.n462 B.n293 163.367
R745 B.n462 B.n287 163.367
R746 B.n470 B.n287 163.367
R747 B.n470 B.n285 163.367
R748 B.n474 B.n285 163.367
R749 B.n474 B.n279 163.367
R750 B.n482 B.n279 163.367
R751 B.n482 B.n277 163.367
R752 B.n486 B.n277 163.367
R753 B.n486 B.n271 163.367
R754 B.n494 B.n271 163.367
R755 B.n494 B.n269 163.367
R756 B.n498 B.n269 163.367
R757 B.n498 B.n263 163.367
R758 B.n506 B.n263 163.367
R759 B.n506 B.n261 163.367
R760 B.n510 B.n261 163.367
R761 B.n510 B.n255 163.367
R762 B.n519 B.n255 163.367
R763 B.n519 B.n253 163.367
R764 B.n523 B.n253 163.367
R765 B.n523 B.n248 163.367
R766 B.n531 B.n248 163.367
R767 B.n531 B.n246 163.367
R768 B.n535 B.n246 163.367
R769 B.n535 B.n240 163.367
R770 B.n543 B.n240 163.367
R771 B.n543 B.n238 163.367
R772 B.n547 B.n238 163.367
R773 B.n547 B.n232 163.367
R774 B.n556 B.n232 163.367
R775 B.n556 B.n230 163.367
R776 B.n560 B.n230 163.367
R777 B.n560 B.n3 163.367
R778 B.n690 B.n3 163.367
R779 B.n686 B.n2 163.367
R780 B.n686 B.n685 163.367
R781 B.n685 B.n9 163.367
R782 B.n681 B.n9 163.367
R783 B.n681 B.n11 163.367
R784 B.n677 B.n11 163.367
R785 B.n677 B.n16 163.367
R786 B.n673 B.n16 163.367
R787 B.n673 B.n18 163.367
R788 B.n669 B.n18 163.367
R789 B.n669 B.n23 163.367
R790 B.n665 B.n23 163.367
R791 B.n665 B.n25 163.367
R792 B.n661 B.n25 163.367
R793 B.n661 B.n29 163.367
R794 B.n657 B.n29 163.367
R795 B.n657 B.n31 163.367
R796 B.n653 B.n31 163.367
R797 B.n653 B.n37 163.367
R798 B.n649 B.n37 163.367
R799 B.n649 B.n39 163.367
R800 B.n645 B.n39 163.367
R801 B.n645 B.n44 163.367
R802 B.n641 B.n44 163.367
R803 B.n641 B.n46 163.367
R804 B.n637 B.n46 163.367
R805 B.n637 B.n51 163.367
R806 B.n633 B.n51 163.367
R807 B.n633 B.n53 163.367
R808 B.n629 B.n53 163.367
R809 B.n629 B.n58 163.367
R810 B.n625 B.n58 163.367
R811 B.n625 B.n60 163.367
R812 B.n621 B.n60 163.367
R813 B.n621 B.n65 163.367
R814 B.n100 B.t17 110.812
R815 B.n331 B.t11 110.812
R816 B.n102 B.t14 110.805
R817 B.n328 B.t21 110.805
R818 B.n456 B.n292 98.5875
R819 B.n615 B.n64 98.5875
R820 B.n101 B.t18 74.9334
R821 B.n332 B.t10 74.9334
R822 B.n103 B.t15 74.9256
R823 B.n329 B.t20 74.9256
R824 B.n617 B.n616 71.676
R825 B.n104 B.n68 71.676
R826 B.n108 B.n69 71.676
R827 B.n112 B.n70 71.676
R828 B.n116 B.n71 71.676
R829 B.n120 B.n72 71.676
R830 B.n124 B.n73 71.676
R831 B.n128 B.n74 71.676
R832 B.n132 B.n75 71.676
R833 B.n136 B.n76 71.676
R834 B.n140 B.n77 71.676
R835 B.n144 B.n78 71.676
R836 B.n148 B.n79 71.676
R837 B.n152 B.n80 71.676
R838 B.n157 B.n81 71.676
R839 B.n161 B.n82 71.676
R840 B.n165 B.n83 71.676
R841 B.n169 B.n84 71.676
R842 B.n173 B.n85 71.676
R843 B.n178 B.n86 71.676
R844 B.n182 B.n87 71.676
R845 B.n186 B.n88 71.676
R846 B.n190 B.n89 71.676
R847 B.n194 B.n90 71.676
R848 B.n198 B.n91 71.676
R849 B.n202 B.n92 71.676
R850 B.n206 B.n93 71.676
R851 B.n210 B.n94 71.676
R852 B.n214 B.n95 71.676
R853 B.n218 B.n96 71.676
R854 B.n222 B.n97 71.676
R855 B.n614 B.n98 71.676
R856 B.n614 B.n613 71.676
R857 B.n224 B.n97 71.676
R858 B.n221 B.n96 71.676
R859 B.n217 B.n95 71.676
R860 B.n213 B.n94 71.676
R861 B.n209 B.n93 71.676
R862 B.n205 B.n92 71.676
R863 B.n201 B.n91 71.676
R864 B.n197 B.n90 71.676
R865 B.n193 B.n89 71.676
R866 B.n189 B.n88 71.676
R867 B.n185 B.n87 71.676
R868 B.n181 B.n86 71.676
R869 B.n177 B.n85 71.676
R870 B.n172 B.n84 71.676
R871 B.n168 B.n83 71.676
R872 B.n164 B.n82 71.676
R873 B.n160 B.n81 71.676
R874 B.n156 B.n80 71.676
R875 B.n151 B.n79 71.676
R876 B.n147 B.n78 71.676
R877 B.n143 B.n77 71.676
R878 B.n139 B.n76 71.676
R879 B.n135 B.n75 71.676
R880 B.n131 B.n74 71.676
R881 B.n127 B.n73 71.676
R882 B.n123 B.n72 71.676
R883 B.n119 B.n71 71.676
R884 B.n115 B.n70 71.676
R885 B.n111 B.n69 71.676
R886 B.n107 B.n68 71.676
R887 B.n616 B.n67 71.676
R888 B.n458 B.n457 71.676
R889 B.n327 B.n296 71.676
R890 B.n450 B.n297 71.676
R891 B.n446 B.n298 71.676
R892 B.n442 B.n299 71.676
R893 B.n438 B.n300 71.676
R894 B.n434 B.n301 71.676
R895 B.n430 B.n302 71.676
R896 B.n426 B.n303 71.676
R897 B.n422 B.n304 71.676
R898 B.n418 B.n305 71.676
R899 B.n414 B.n306 71.676
R900 B.n410 B.n307 71.676
R901 B.n406 B.n308 71.676
R902 B.n402 B.n309 71.676
R903 B.n398 B.n310 71.676
R904 B.n394 B.n311 71.676
R905 B.n390 B.n312 71.676
R906 B.n386 B.n313 71.676
R907 B.n382 B.n314 71.676
R908 B.n378 B.n315 71.676
R909 B.n374 B.n316 71.676
R910 B.n370 B.n317 71.676
R911 B.n366 B.n318 71.676
R912 B.n362 B.n319 71.676
R913 B.n358 B.n320 71.676
R914 B.n354 B.n321 71.676
R915 B.n350 B.n322 71.676
R916 B.n346 B.n323 71.676
R917 B.n342 B.n324 71.676
R918 B.n338 B.n325 71.676
R919 B.n457 B.n295 71.676
R920 B.n451 B.n296 71.676
R921 B.n447 B.n297 71.676
R922 B.n443 B.n298 71.676
R923 B.n439 B.n299 71.676
R924 B.n435 B.n300 71.676
R925 B.n431 B.n301 71.676
R926 B.n427 B.n302 71.676
R927 B.n423 B.n303 71.676
R928 B.n419 B.n304 71.676
R929 B.n415 B.n305 71.676
R930 B.n411 B.n306 71.676
R931 B.n407 B.n307 71.676
R932 B.n403 B.n308 71.676
R933 B.n399 B.n309 71.676
R934 B.n395 B.n310 71.676
R935 B.n391 B.n311 71.676
R936 B.n387 B.n312 71.676
R937 B.n383 B.n313 71.676
R938 B.n379 B.n314 71.676
R939 B.n375 B.n315 71.676
R940 B.n371 B.n316 71.676
R941 B.n367 B.n317 71.676
R942 B.n363 B.n318 71.676
R943 B.n359 B.n319 71.676
R944 B.n355 B.n320 71.676
R945 B.n351 B.n321 71.676
R946 B.n347 B.n322 71.676
R947 B.n343 B.n323 71.676
R948 B.n339 B.n324 71.676
R949 B.n335 B.n325 71.676
R950 B.n691 B.n690 71.676
R951 B.n691 B.n2 71.676
R952 B.n463 B.n292 60.3961
R953 B.n463 B.n288 60.3961
R954 B.n469 B.n288 60.3961
R955 B.n469 B.n283 60.3961
R956 B.n475 B.n283 60.3961
R957 B.n475 B.n284 60.3961
R958 B.n481 B.n276 60.3961
R959 B.n487 B.n276 60.3961
R960 B.n487 B.n272 60.3961
R961 B.n493 B.n272 60.3961
R962 B.n493 B.n267 60.3961
R963 B.n499 B.n267 60.3961
R964 B.n499 B.n268 60.3961
R965 B.n505 B.n260 60.3961
R966 B.n511 B.n260 60.3961
R967 B.n511 B.n256 60.3961
R968 B.n518 B.n256 60.3961
R969 B.n518 B.n517 60.3961
R970 B.n524 B.n249 60.3961
R971 B.n530 B.n249 60.3961
R972 B.n530 B.n245 60.3961
R973 B.n536 B.n245 60.3961
R974 B.n542 B.n241 60.3961
R975 B.n542 B.n237 60.3961
R976 B.n548 B.n237 60.3961
R977 B.n548 B.n233 60.3961
R978 B.n555 B.n233 60.3961
R979 B.n561 B.n229 60.3961
R980 B.n561 B.n4 60.3961
R981 B.n689 B.n4 60.3961
R982 B.n689 B.n688 60.3961
R983 B.n688 B.n687 60.3961
R984 B.n687 B.n8 60.3961
R985 B.n570 B.n8 60.3961
R986 B.n680 B.n679 60.3961
R987 B.n679 B.n678 60.3961
R988 B.n678 B.n15 60.3961
R989 B.n672 B.n15 60.3961
R990 B.n672 B.n671 60.3961
R991 B.n670 B.n22 60.3961
R992 B.n664 B.n22 60.3961
R993 B.n664 B.n663 60.3961
R994 B.n663 B.n662 60.3961
R995 B.n656 B.n32 60.3961
R996 B.n656 B.n655 60.3961
R997 B.n655 B.n654 60.3961
R998 B.n654 B.n36 60.3961
R999 B.n648 B.n36 60.3961
R1000 B.n647 B.n646 60.3961
R1001 B.n646 B.n43 60.3961
R1002 B.n640 B.n43 60.3961
R1003 B.n640 B.n639 60.3961
R1004 B.n639 B.n638 60.3961
R1005 B.n638 B.n50 60.3961
R1006 B.n632 B.n50 60.3961
R1007 B.n631 B.n630 60.3961
R1008 B.n630 B.n57 60.3961
R1009 B.n624 B.n57 60.3961
R1010 B.n624 B.n623 60.3961
R1011 B.n623 B.n622 60.3961
R1012 B.n622 B.n64 60.3961
R1013 B.n154 B.n103 59.5399
R1014 B.n175 B.n101 59.5399
R1015 B.n333 B.n332 59.5399
R1016 B.n330 B.n329 59.5399
R1017 B.n268 B.t3 51.5144
R1018 B.t7 B.n647 51.5144
R1019 B.t2 B.n229 49.7381
R1020 B.n570 B.t1 49.7381
R1021 B.n481 B.t9 47.9617
R1022 B.n632 B.t13 47.9617
R1023 B.n536 B.t5 44.4091
R1024 B.t6 B.n670 44.4091
R1025 B.n524 B.t0 42.6327
R1026 B.n662 B.t4 42.6327
R1027 B.n103 B.n102 35.8793
R1028 B.n101 B.n100 35.8793
R1029 B.n332 B.n331 35.8793
R1030 B.n329 B.n328 35.8793
R1031 B.n460 B.n459 30.7517
R1032 B.n334 B.n290 30.7517
R1033 B.n619 B.n618 30.7517
R1034 B.n612 B.n611 30.7517
R1035 B B.n692 18.0485
R1036 B.n517 B.t0 17.7639
R1037 B.n32 B.t4 17.7639
R1038 B.t5 B.n241 15.9876
R1039 B.n671 B.t6 15.9876
R1040 B.n284 B.t9 12.4349
R1041 B.t13 B.n631 12.4349
R1042 B.n555 B.t2 10.6586
R1043 B.n680 B.t1 10.6586
R1044 B.n461 B.n460 10.6151
R1045 B.n461 B.n286 10.6151
R1046 B.n471 B.n286 10.6151
R1047 B.n472 B.n471 10.6151
R1048 B.n473 B.n472 10.6151
R1049 B.n473 B.n278 10.6151
R1050 B.n483 B.n278 10.6151
R1051 B.n484 B.n483 10.6151
R1052 B.n485 B.n484 10.6151
R1053 B.n485 B.n270 10.6151
R1054 B.n495 B.n270 10.6151
R1055 B.n496 B.n495 10.6151
R1056 B.n497 B.n496 10.6151
R1057 B.n497 B.n262 10.6151
R1058 B.n507 B.n262 10.6151
R1059 B.n508 B.n507 10.6151
R1060 B.n509 B.n508 10.6151
R1061 B.n509 B.n254 10.6151
R1062 B.n520 B.n254 10.6151
R1063 B.n521 B.n520 10.6151
R1064 B.n522 B.n521 10.6151
R1065 B.n522 B.n247 10.6151
R1066 B.n532 B.n247 10.6151
R1067 B.n533 B.n532 10.6151
R1068 B.n534 B.n533 10.6151
R1069 B.n534 B.n239 10.6151
R1070 B.n544 B.n239 10.6151
R1071 B.n545 B.n544 10.6151
R1072 B.n546 B.n545 10.6151
R1073 B.n546 B.n231 10.6151
R1074 B.n557 B.n231 10.6151
R1075 B.n558 B.n557 10.6151
R1076 B.n559 B.n558 10.6151
R1077 B.n559 B.n0 10.6151
R1078 B.n459 B.n294 10.6151
R1079 B.n454 B.n294 10.6151
R1080 B.n454 B.n453 10.6151
R1081 B.n453 B.n452 10.6151
R1082 B.n452 B.n449 10.6151
R1083 B.n449 B.n448 10.6151
R1084 B.n448 B.n445 10.6151
R1085 B.n445 B.n444 10.6151
R1086 B.n444 B.n441 10.6151
R1087 B.n441 B.n440 10.6151
R1088 B.n440 B.n437 10.6151
R1089 B.n437 B.n436 10.6151
R1090 B.n436 B.n433 10.6151
R1091 B.n433 B.n432 10.6151
R1092 B.n432 B.n429 10.6151
R1093 B.n429 B.n428 10.6151
R1094 B.n428 B.n425 10.6151
R1095 B.n425 B.n424 10.6151
R1096 B.n424 B.n421 10.6151
R1097 B.n421 B.n420 10.6151
R1098 B.n420 B.n417 10.6151
R1099 B.n417 B.n416 10.6151
R1100 B.n416 B.n413 10.6151
R1101 B.n413 B.n412 10.6151
R1102 B.n412 B.n409 10.6151
R1103 B.n409 B.n408 10.6151
R1104 B.n405 B.n404 10.6151
R1105 B.n404 B.n401 10.6151
R1106 B.n401 B.n400 10.6151
R1107 B.n400 B.n397 10.6151
R1108 B.n397 B.n396 10.6151
R1109 B.n396 B.n393 10.6151
R1110 B.n393 B.n392 10.6151
R1111 B.n392 B.n389 10.6151
R1112 B.n389 B.n388 10.6151
R1113 B.n385 B.n384 10.6151
R1114 B.n384 B.n381 10.6151
R1115 B.n381 B.n380 10.6151
R1116 B.n380 B.n377 10.6151
R1117 B.n377 B.n376 10.6151
R1118 B.n376 B.n373 10.6151
R1119 B.n373 B.n372 10.6151
R1120 B.n372 B.n369 10.6151
R1121 B.n369 B.n368 10.6151
R1122 B.n368 B.n365 10.6151
R1123 B.n365 B.n364 10.6151
R1124 B.n364 B.n361 10.6151
R1125 B.n361 B.n360 10.6151
R1126 B.n360 B.n357 10.6151
R1127 B.n357 B.n356 10.6151
R1128 B.n356 B.n353 10.6151
R1129 B.n353 B.n352 10.6151
R1130 B.n352 B.n349 10.6151
R1131 B.n349 B.n348 10.6151
R1132 B.n348 B.n345 10.6151
R1133 B.n345 B.n344 10.6151
R1134 B.n344 B.n341 10.6151
R1135 B.n341 B.n340 10.6151
R1136 B.n340 B.n337 10.6151
R1137 B.n337 B.n336 10.6151
R1138 B.n336 B.n334 10.6151
R1139 B.n465 B.n290 10.6151
R1140 B.n466 B.n465 10.6151
R1141 B.n467 B.n466 10.6151
R1142 B.n467 B.n281 10.6151
R1143 B.n477 B.n281 10.6151
R1144 B.n478 B.n477 10.6151
R1145 B.n479 B.n478 10.6151
R1146 B.n479 B.n274 10.6151
R1147 B.n489 B.n274 10.6151
R1148 B.n490 B.n489 10.6151
R1149 B.n491 B.n490 10.6151
R1150 B.n491 B.n265 10.6151
R1151 B.n501 B.n265 10.6151
R1152 B.n502 B.n501 10.6151
R1153 B.n503 B.n502 10.6151
R1154 B.n503 B.n258 10.6151
R1155 B.n513 B.n258 10.6151
R1156 B.n514 B.n513 10.6151
R1157 B.n515 B.n514 10.6151
R1158 B.n515 B.n251 10.6151
R1159 B.n526 B.n251 10.6151
R1160 B.n527 B.n526 10.6151
R1161 B.n528 B.n527 10.6151
R1162 B.n528 B.n243 10.6151
R1163 B.n538 B.n243 10.6151
R1164 B.n539 B.n538 10.6151
R1165 B.n540 B.n539 10.6151
R1166 B.n540 B.n235 10.6151
R1167 B.n550 B.n235 10.6151
R1168 B.n551 B.n550 10.6151
R1169 B.n553 B.n551 10.6151
R1170 B.n553 B.n552 10.6151
R1171 B.n552 B.n227 10.6151
R1172 B.n564 B.n227 10.6151
R1173 B.n565 B.n564 10.6151
R1174 B.n566 B.n565 10.6151
R1175 B.n567 B.n566 10.6151
R1176 B.n568 B.n567 10.6151
R1177 B.n572 B.n568 10.6151
R1178 B.n573 B.n572 10.6151
R1179 B.n574 B.n573 10.6151
R1180 B.n575 B.n574 10.6151
R1181 B.n577 B.n575 10.6151
R1182 B.n578 B.n577 10.6151
R1183 B.n579 B.n578 10.6151
R1184 B.n580 B.n579 10.6151
R1185 B.n582 B.n580 10.6151
R1186 B.n583 B.n582 10.6151
R1187 B.n584 B.n583 10.6151
R1188 B.n585 B.n584 10.6151
R1189 B.n587 B.n585 10.6151
R1190 B.n588 B.n587 10.6151
R1191 B.n589 B.n588 10.6151
R1192 B.n590 B.n589 10.6151
R1193 B.n592 B.n590 10.6151
R1194 B.n593 B.n592 10.6151
R1195 B.n594 B.n593 10.6151
R1196 B.n595 B.n594 10.6151
R1197 B.n597 B.n595 10.6151
R1198 B.n598 B.n597 10.6151
R1199 B.n599 B.n598 10.6151
R1200 B.n600 B.n599 10.6151
R1201 B.n602 B.n600 10.6151
R1202 B.n603 B.n602 10.6151
R1203 B.n604 B.n603 10.6151
R1204 B.n605 B.n604 10.6151
R1205 B.n607 B.n605 10.6151
R1206 B.n608 B.n607 10.6151
R1207 B.n609 B.n608 10.6151
R1208 B.n610 B.n609 10.6151
R1209 B.n611 B.n610 10.6151
R1210 B.n684 B.n1 10.6151
R1211 B.n684 B.n683 10.6151
R1212 B.n683 B.n682 10.6151
R1213 B.n682 B.n10 10.6151
R1214 B.n676 B.n10 10.6151
R1215 B.n676 B.n675 10.6151
R1216 B.n675 B.n674 10.6151
R1217 B.n674 B.n17 10.6151
R1218 B.n668 B.n17 10.6151
R1219 B.n668 B.n667 10.6151
R1220 B.n667 B.n666 10.6151
R1221 B.n666 B.n24 10.6151
R1222 B.n660 B.n24 10.6151
R1223 B.n660 B.n659 10.6151
R1224 B.n659 B.n658 10.6151
R1225 B.n658 B.n30 10.6151
R1226 B.n652 B.n30 10.6151
R1227 B.n652 B.n651 10.6151
R1228 B.n651 B.n650 10.6151
R1229 B.n650 B.n38 10.6151
R1230 B.n644 B.n38 10.6151
R1231 B.n644 B.n643 10.6151
R1232 B.n643 B.n642 10.6151
R1233 B.n642 B.n45 10.6151
R1234 B.n636 B.n45 10.6151
R1235 B.n636 B.n635 10.6151
R1236 B.n635 B.n634 10.6151
R1237 B.n634 B.n52 10.6151
R1238 B.n628 B.n52 10.6151
R1239 B.n628 B.n627 10.6151
R1240 B.n627 B.n626 10.6151
R1241 B.n626 B.n59 10.6151
R1242 B.n620 B.n59 10.6151
R1243 B.n620 B.n619 10.6151
R1244 B.n618 B.n66 10.6151
R1245 B.n105 B.n66 10.6151
R1246 B.n106 B.n105 10.6151
R1247 B.n109 B.n106 10.6151
R1248 B.n110 B.n109 10.6151
R1249 B.n113 B.n110 10.6151
R1250 B.n114 B.n113 10.6151
R1251 B.n117 B.n114 10.6151
R1252 B.n118 B.n117 10.6151
R1253 B.n121 B.n118 10.6151
R1254 B.n122 B.n121 10.6151
R1255 B.n125 B.n122 10.6151
R1256 B.n126 B.n125 10.6151
R1257 B.n129 B.n126 10.6151
R1258 B.n130 B.n129 10.6151
R1259 B.n133 B.n130 10.6151
R1260 B.n134 B.n133 10.6151
R1261 B.n137 B.n134 10.6151
R1262 B.n138 B.n137 10.6151
R1263 B.n141 B.n138 10.6151
R1264 B.n142 B.n141 10.6151
R1265 B.n145 B.n142 10.6151
R1266 B.n146 B.n145 10.6151
R1267 B.n149 B.n146 10.6151
R1268 B.n150 B.n149 10.6151
R1269 B.n153 B.n150 10.6151
R1270 B.n158 B.n155 10.6151
R1271 B.n159 B.n158 10.6151
R1272 B.n162 B.n159 10.6151
R1273 B.n163 B.n162 10.6151
R1274 B.n166 B.n163 10.6151
R1275 B.n167 B.n166 10.6151
R1276 B.n170 B.n167 10.6151
R1277 B.n171 B.n170 10.6151
R1278 B.n174 B.n171 10.6151
R1279 B.n179 B.n176 10.6151
R1280 B.n180 B.n179 10.6151
R1281 B.n183 B.n180 10.6151
R1282 B.n184 B.n183 10.6151
R1283 B.n187 B.n184 10.6151
R1284 B.n188 B.n187 10.6151
R1285 B.n191 B.n188 10.6151
R1286 B.n192 B.n191 10.6151
R1287 B.n195 B.n192 10.6151
R1288 B.n196 B.n195 10.6151
R1289 B.n199 B.n196 10.6151
R1290 B.n200 B.n199 10.6151
R1291 B.n203 B.n200 10.6151
R1292 B.n204 B.n203 10.6151
R1293 B.n207 B.n204 10.6151
R1294 B.n208 B.n207 10.6151
R1295 B.n211 B.n208 10.6151
R1296 B.n212 B.n211 10.6151
R1297 B.n215 B.n212 10.6151
R1298 B.n216 B.n215 10.6151
R1299 B.n219 B.n216 10.6151
R1300 B.n220 B.n219 10.6151
R1301 B.n223 B.n220 10.6151
R1302 B.n225 B.n223 10.6151
R1303 B.n226 B.n225 10.6151
R1304 B.n612 B.n226 10.6151
R1305 B.n408 B.n330 9.36635
R1306 B.n385 B.n333 9.36635
R1307 B.n154 B.n153 9.36635
R1308 B.n176 B.n175 9.36635
R1309 B.n505 B.t3 8.88221
R1310 B.n648 B.t7 8.88221
R1311 B.n692 B.n0 8.11757
R1312 B.n692 B.n1 8.11757
R1313 B.n405 B.n330 1.24928
R1314 B.n388 B.n333 1.24928
R1315 B.n155 B.n154 1.24928
R1316 B.n175 B.n174 1.24928
R1317 VN.n18 VN.n17 172.31
R1318 VN.n37 VN.n36 172.31
R1319 VN.n35 VN.n19 161.3
R1320 VN.n34 VN.n33 161.3
R1321 VN.n32 VN.n20 161.3
R1322 VN.n31 VN.n30 161.3
R1323 VN.n28 VN.n21 161.3
R1324 VN.n27 VN.n26 161.3
R1325 VN.n25 VN.n22 161.3
R1326 VN.n16 VN.n0 161.3
R1327 VN.n15 VN.n14 161.3
R1328 VN.n13 VN.n1 161.3
R1329 VN.n12 VN.n11 161.3
R1330 VN.n9 VN.n2 161.3
R1331 VN.n8 VN.n7 161.3
R1332 VN.n6 VN.n3 161.3
R1333 VN.n5 VN.t4 148.417
R1334 VN.n24 VN.t5 148.417
R1335 VN.n4 VN.t7 112.731
R1336 VN.n10 VN.t6 112.731
R1337 VN.n17 VN.t2 112.731
R1338 VN.n23 VN.t1 112.731
R1339 VN.n29 VN.t3 112.731
R1340 VN.n36 VN.t0 112.731
R1341 VN.n15 VN.n1 55.0624
R1342 VN.n34 VN.n20 55.0624
R1343 VN.n5 VN.n4 45.8064
R1344 VN.n24 VN.n23 45.8064
R1345 VN VN.n37 42.5024
R1346 VN.n8 VN.n3 40.4934
R1347 VN.n9 VN.n8 40.4934
R1348 VN.n27 VN.n22 40.4934
R1349 VN.n28 VN.n27 40.4934
R1350 VN.n16 VN.n15 25.9244
R1351 VN.n35 VN.n34 25.9244
R1352 VN.n11 VN.n1 24.4675
R1353 VN.n30 VN.n20 24.4675
R1354 VN.n4 VN.n3 20.7975
R1355 VN.n10 VN.n9 20.7975
R1356 VN.n23 VN.n22 20.7975
R1357 VN.n29 VN.n28 20.7975
R1358 VN.n25 VN.n24 17.4308
R1359 VN.n6 VN.n5 17.4308
R1360 VN.n17 VN.n16 13.4574
R1361 VN.n36 VN.n35 13.4574
R1362 VN.n11 VN.n10 3.67055
R1363 VN.n30 VN.n29 3.67055
R1364 VN.n37 VN.n19 0.189894
R1365 VN.n33 VN.n19 0.189894
R1366 VN.n33 VN.n32 0.189894
R1367 VN.n32 VN.n31 0.189894
R1368 VN.n31 VN.n21 0.189894
R1369 VN.n26 VN.n21 0.189894
R1370 VN.n26 VN.n25 0.189894
R1371 VN.n7 VN.n6 0.189894
R1372 VN.n7 VN.n2 0.189894
R1373 VN.n12 VN.n2 0.189894
R1374 VN.n13 VN.n12 0.189894
R1375 VN.n14 VN.n13 0.189894
R1376 VN.n14 VN.n0 0.189894
R1377 VN.n18 VN.n0 0.189894
R1378 VN VN.n18 0.0516364
R1379 VDD2.n2 VDD2.n1 66.9351
R1380 VDD2.n2 VDD2.n0 66.9351
R1381 VDD2 VDD2.n5 66.9321
R1382 VDD2.n4 VDD2.n3 66.1931
R1383 VDD2.n4 VDD2.n2 37.0213
R1384 VDD2.n5 VDD2.t6 2.78531
R1385 VDD2.n5 VDD2.t2 2.78531
R1386 VDD2.n3 VDD2.t7 2.78531
R1387 VDD2.n3 VDD2.t4 2.78531
R1388 VDD2.n1 VDD2.t1 2.78531
R1389 VDD2.n1 VDD2.t5 2.78531
R1390 VDD2.n0 VDD2.t3 2.78531
R1391 VDD2.n0 VDD2.t0 2.78531
R1392 VDD2 VDD2.n4 0.856103
C0 VDD1 VP 4.92039f
C1 VN VDD2 4.66627f
C2 VTAIL VDD1 6.20166f
C3 VP VDD2 0.404746f
C4 VN VP 5.43324f
C5 VTAIL VDD2 6.24883f
C6 VTAIL VN 5.02448f
C7 VTAIL VP 5.03859f
C8 VDD1 VDD2 1.23071f
C9 VDD1 VN 0.149774f
C10 VDD2 B 3.914333f
C11 VDD1 B 4.236868f
C12 VTAIL B 6.565649f
C13 VN B 10.868641f
C14 VP B 9.383996f
C15 VDD2.t3 B 0.139322f
C16 VDD2.t0 B 0.139322f
C17 VDD2.n0 B 1.18916f
C18 VDD2.t1 B 0.139322f
C19 VDD2.t5 B 0.139322f
C20 VDD2.n1 B 1.18916f
C21 VDD2.n2 B 2.33373f
C22 VDD2.t7 B 0.139322f
C23 VDD2.t4 B 0.139322f
C24 VDD2.n3 B 1.18471f
C25 VDD2.n4 B 2.17599f
C26 VDD2.t6 B 0.139322f
C27 VDD2.t2 B 0.139322f
C28 VDD2.n5 B 1.18913f
C29 VN.n0 B 0.032167f
C30 VN.t2 B 0.928574f
C31 VN.n1 B 0.055673f
C32 VN.n2 B 0.032167f
C33 VN.t6 B 0.928574f
C34 VN.n3 B 0.059491f
C35 VN.t4 B 1.04464f
C36 VN.t7 B 0.928574f
C37 VN.n4 B 0.425638f
C38 VN.n5 B 0.418387f
C39 VN.n6 B 0.205657f
C40 VN.n7 B 0.032167f
C41 VN.n8 B 0.026004f
C42 VN.n9 B 0.059491f
C43 VN.n10 B 0.354345f
C44 VN.n11 B 0.034792f
C45 VN.n12 B 0.032167f
C46 VN.n13 B 0.032167f
C47 VN.n14 B 0.032167f
C48 VN.n15 B 0.036682f
C49 VN.n16 B 0.048193f
C50 VN.n17 B 0.426812f
C51 VN.n18 B 0.029875f
C52 VN.n19 B 0.032167f
C53 VN.t0 B 0.928574f
C54 VN.n20 B 0.055673f
C55 VN.n21 B 0.032167f
C56 VN.t3 B 0.928574f
C57 VN.n22 B 0.059491f
C58 VN.t5 B 1.04464f
C59 VN.t1 B 0.928574f
C60 VN.n23 B 0.425638f
C61 VN.n24 B 0.418387f
C62 VN.n25 B 0.205657f
C63 VN.n26 B 0.032167f
C64 VN.n27 B 0.026004f
C65 VN.n28 B 0.059491f
C66 VN.n29 B 0.354345f
C67 VN.n30 B 0.034792f
C68 VN.n31 B 0.032167f
C69 VN.n32 B 0.032167f
C70 VN.n33 B 0.032167f
C71 VN.n34 B 0.036682f
C72 VN.n35 B 0.048193f
C73 VN.n36 B 0.426812f
C74 VN.n37 B 1.36024f
C75 VTAIL.t6 B 0.118123f
C76 VTAIL.t4 B 0.118123f
C77 VTAIL.n0 B 0.947516f
C78 VTAIL.n1 B 0.31334f
C79 VTAIL.t1 B 1.20835f
C80 VTAIL.n2 B 0.402547f
C81 VTAIL.t9 B 1.20835f
C82 VTAIL.n3 B 0.402547f
C83 VTAIL.t14 B 0.118123f
C84 VTAIL.t15 B 0.118123f
C85 VTAIL.n4 B 0.947516f
C86 VTAIL.n5 B 0.417437f
C87 VTAIL.t12 B 1.20835f
C88 VTAIL.n6 B 1.17956f
C89 VTAIL.t3 B 1.20835f
C90 VTAIL.n7 B 1.17955f
C91 VTAIL.t0 B 0.118123f
C92 VTAIL.t5 B 0.118123f
C93 VTAIL.n8 B 0.947517f
C94 VTAIL.n9 B 0.417435f
C95 VTAIL.t2 B 1.20835f
C96 VTAIL.n10 B 0.402542f
C97 VTAIL.t11 B 1.20835f
C98 VTAIL.n11 B 0.402542f
C99 VTAIL.t8 B 0.118123f
C100 VTAIL.t13 B 0.118123f
C101 VTAIL.n12 B 0.947517f
C102 VTAIL.n13 B 0.417435f
C103 VTAIL.t10 B 1.20835f
C104 VTAIL.n14 B 1.17956f
C105 VTAIL.t7 B 1.20835f
C106 VTAIL.n15 B 1.17562f
C107 VDD1.t6 B 0.140696f
C108 VDD1.t2 B 0.140696f
C109 VDD1.n0 B 1.20168f
C110 VDD1.t7 B 0.140696f
C111 VDD1.t4 B 0.140696f
C112 VDD1.n1 B 1.20089f
C113 VDD1.t0 B 0.140696f
C114 VDD1.t1 B 0.140696f
C115 VDD1.n2 B 1.20089f
C116 VDD1.n3 B 2.40976f
C117 VDD1.t3 B 0.140696f
C118 VDD1.t5 B 0.140696f
C119 VDD1.n4 B 1.19639f
C120 VDD1.n5 B 2.22755f
C121 VP.n0 B 0.032691f
C122 VP.t6 B 0.943699f
C123 VP.n1 B 0.05658f
C124 VP.n2 B 0.032691f
C125 VP.t0 B 0.943699f
C126 VP.n3 B 0.06046f
C127 VP.n4 B 0.032691f
C128 VP.n5 B 0.048978f
C129 VP.n6 B 0.032691f
C130 VP.t5 B 0.943699f
C131 VP.n7 B 0.05658f
C132 VP.n8 B 0.032691f
C133 VP.t2 B 0.943699f
C134 VP.n9 B 0.06046f
C135 VP.t4 B 1.06166f
C136 VP.t7 B 0.943699f
C137 VP.n10 B 0.432571f
C138 VP.n11 B 0.425202f
C139 VP.n12 B 0.209007f
C140 VP.n13 B 0.032691f
C141 VP.n14 B 0.026428f
C142 VP.n15 B 0.06046f
C143 VP.n16 B 0.360117f
C144 VP.n17 B 0.035358f
C145 VP.n18 B 0.032691f
C146 VP.n19 B 0.032691f
C147 VP.n20 B 0.032691f
C148 VP.n21 B 0.03728f
C149 VP.n22 B 0.048978f
C150 VP.n23 B 0.433764f
C151 VP.n24 B 1.36094f
C152 VP.t3 B 0.943699f
C153 VP.n25 B 0.433764f
C154 VP.n26 B 1.38884f
C155 VP.n27 B 0.032691f
C156 VP.n28 B 0.032691f
C157 VP.n29 B 0.03728f
C158 VP.n30 B 0.05658f
C159 VP.t1 B 0.943699f
C160 VP.n31 B 0.360117f
C161 VP.n32 B 0.035358f
C162 VP.n33 B 0.032691f
C163 VP.n34 B 0.032691f
C164 VP.n35 B 0.032691f
C165 VP.n36 B 0.026428f
C166 VP.n37 B 0.06046f
C167 VP.n38 B 0.360117f
C168 VP.n39 B 0.035358f
C169 VP.n40 B 0.032691f
C170 VP.n41 B 0.032691f
C171 VP.n42 B 0.032691f
C172 VP.n43 B 0.03728f
C173 VP.n44 B 0.048978f
C174 VP.n45 B 0.433764f
C175 VP.n46 B 0.030362f
.ends

