* NGSPICE file created from diff_pair_sample_0417.ext - technology: sky130A

.subckt diff_pair_sample_0417 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X1 VTAIL.t14 VN.t1 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0.71115 ps=4.64 w=4.31 l=0.39
X2 VTAIL.t1 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X3 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0 ps=0 w=4.31 l=0.39
X4 VDD2.t0 VN.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X5 VDD1.t6 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=1.6809 ps=9.4 w=4.31 l=0.39
X6 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X7 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0.71115 ps=4.64 w=4.31 l=0.39
X8 VTAIL.t12 VN.t3 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X9 VDD2.t2 VN.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=1.6809 ps=9.4 w=4.31 l=0.39
X10 VDD2.t3 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X11 VTAIL.t2 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0.71115 ps=4.64 w=4.31 l=0.39
X12 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0 ps=0 w=4.31 l=0.39
X13 VDD1.t2 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=1.6809 ps=9.4 w=4.31 l=0.39
X14 VDD1.t1 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X15 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0 ps=0 w=4.31 l=0.39
X16 VTAIL.t9 VN.t6 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0.71115 ps=4.64 w=4.31 l=0.39
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6809 pd=9.4 as=0 ps=0 w=4.31 l=0.39
X18 VDD1.t0 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=0.71115 ps=4.64 w=4.31 l=0.39
X19 VDD2.t6 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.71115 pd=4.64 as=1.6809 ps=9.4 w=4.31 l=0.39
R0 VN.n1 VN.t6 400.493
R1 VN.n7 VN.t4 400.493
R2 VN.n4 VN.t7 387.399
R3 VN.n10 VN.t1 387.399
R4 VN.n2 VN.t2 367.68
R5 VN.n3 VN.t3 367.68
R6 VN.n8 VN.t0 367.68
R7 VN.n9 VN.t5 367.68
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 161.3
R11 VN.n3 VN.n0 161.3
R12 VN.n7 VN.n6 74.3446
R13 VN.n1 VN.n0 74.3446
R14 VN.n3 VN.n2 48.2005
R15 VN.n9 VN.n8 48.2005
R16 VN VN.n11 35.2372
R17 VN.n4 VN.n3 28.4823
R18 VN.n10 VN.n9 28.4823
R19 VN.n8 VN.n7 13.0795
R20 VN.n2 VN.n1 13.0795
R21 VN.n11 VN.n6 0.189894
R22 VN.n5 VN.n0 0.189894
R23 VN VN.n5 0.0516364
R24 VDD2.n2 VDD2.n1 74.3065
R25 VDD2.n2 VDD2.n0 74.3065
R26 VDD2 VDD2.n5 74.3038
R27 VDD2.n4 VDD2.n3 74.0518
R28 VDD2.n4 VDD2.n2 30.2239
R29 VDD2.n5 VDD2.t4 4.59447
R30 VDD2.n5 VDD2.t2 4.59447
R31 VDD2.n3 VDD2.t1 4.59447
R32 VDD2.n3 VDD2.t3 4.59447
R33 VDD2.n1 VDD2.t5 4.59447
R34 VDD2.n1 VDD2.t6 4.59447
R35 VDD2.n0 VDD2.t7 4.59447
R36 VDD2.n0 VDD2.t0 4.59447
R37 VDD2 VDD2.n4 0.369034
R38 VTAIL.n11 VTAIL.t7 61.967
R39 VTAIL.n10 VTAIL.t11 61.967
R40 VTAIL.n7 VTAIL.t14 61.967
R41 VTAIL.n14 VTAIL.t6 61.9667
R42 VTAIL.n15 VTAIL.t8 61.9667
R43 VTAIL.n2 VTAIL.t9 61.9667
R44 VTAIL.n3 VTAIL.t0 61.9667
R45 VTAIL.n6 VTAIL.t2 61.9667
R46 VTAIL.n13 VTAIL.n12 57.373
R47 VTAIL.n9 VTAIL.n8 57.373
R48 VTAIL.n1 VTAIL.n0 57.3728
R49 VTAIL.n5 VTAIL.n4 57.3728
R50 VTAIL.n15 VTAIL.n14 16.7031
R51 VTAIL.n7 VTAIL.n6 16.7031
R52 VTAIL.n0 VTAIL.t13 4.59447
R53 VTAIL.n0 VTAIL.t12 4.59447
R54 VTAIL.n4 VTAIL.t5 4.59447
R55 VTAIL.n4 VTAIL.t1 4.59447
R56 VTAIL.n12 VTAIL.t3 4.59447
R57 VTAIL.n12 VTAIL.t4 4.59447
R58 VTAIL.n8 VTAIL.t10 4.59447
R59 VTAIL.n8 VTAIL.t15 4.59447
R60 VTAIL.n9 VTAIL.n7 0.62119
R61 VTAIL.n10 VTAIL.n9 0.62119
R62 VTAIL.n13 VTAIL.n11 0.62119
R63 VTAIL.n14 VTAIL.n13 0.62119
R64 VTAIL.n6 VTAIL.n5 0.62119
R65 VTAIL.n5 VTAIL.n3 0.62119
R66 VTAIL.n2 VTAIL.n1 0.62119
R67 VTAIL VTAIL.n15 0.563
R68 VTAIL.n11 VTAIL.n10 0.470328
R69 VTAIL.n3 VTAIL.n2 0.470328
R70 VTAIL VTAIL.n1 0.0586897
R71 B.n306 B.n305 585
R72 B.n308 B.n66 585
R73 B.n311 B.n310 585
R74 B.n312 B.n65 585
R75 B.n314 B.n313 585
R76 B.n316 B.n64 585
R77 B.n319 B.n318 585
R78 B.n320 B.n63 585
R79 B.n322 B.n321 585
R80 B.n324 B.n62 585
R81 B.n327 B.n326 585
R82 B.n328 B.n61 585
R83 B.n330 B.n329 585
R84 B.n332 B.n60 585
R85 B.n335 B.n334 585
R86 B.n336 B.n59 585
R87 B.n338 B.n337 585
R88 B.n340 B.n58 585
R89 B.n343 B.n342 585
R90 B.n345 B.n55 585
R91 B.n347 B.n346 585
R92 B.n349 B.n54 585
R93 B.n352 B.n351 585
R94 B.n353 B.n53 585
R95 B.n355 B.n354 585
R96 B.n357 B.n52 585
R97 B.n360 B.n359 585
R98 B.n361 B.n48 585
R99 B.n363 B.n362 585
R100 B.n365 B.n47 585
R101 B.n368 B.n367 585
R102 B.n369 B.n46 585
R103 B.n371 B.n370 585
R104 B.n373 B.n45 585
R105 B.n376 B.n375 585
R106 B.n377 B.n44 585
R107 B.n379 B.n378 585
R108 B.n381 B.n43 585
R109 B.n384 B.n383 585
R110 B.n385 B.n42 585
R111 B.n387 B.n386 585
R112 B.n389 B.n41 585
R113 B.n392 B.n391 585
R114 B.n393 B.n40 585
R115 B.n395 B.n394 585
R116 B.n397 B.n39 585
R117 B.n400 B.n399 585
R118 B.n401 B.n38 585
R119 B.n304 B.n36 585
R120 B.n404 B.n36 585
R121 B.n303 B.n35 585
R122 B.n405 B.n35 585
R123 B.n302 B.n34 585
R124 B.n406 B.n34 585
R125 B.n301 B.n300 585
R126 B.n300 B.n30 585
R127 B.n299 B.n29 585
R128 B.n412 B.n29 585
R129 B.n298 B.n28 585
R130 B.n413 B.n28 585
R131 B.n297 B.n27 585
R132 B.n414 B.n27 585
R133 B.n296 B.n295 585
R134 B.n295 B.n23 585
R135 B.n294 B.n22 585
R136 B.n420 B.n22 585
R137 B.n293 B.n21 585
R138 B.n421 B.n21 585
R139 B.n292 B.n20 585
R140 B.n422 B.n20 585
R141 B.n291 B.n290 585
R142 B.n290 B.n19 585
R143 B.n289 B.n15 585
R144 B.n428 B.n15 585
R145 B.n288 B.n14 585
R146 B.n429 B.n14 585
R147 B.n287 B.n13 585
R148 B.n430 B.n13 585
R149 B.n286 B.n285 585
R150 B.n285 B.n12 585
R151 B.n284 B.n283 585
R152 B.n284 B.n8 585
R153 B.n282 B.n7 585
R154 B.n437 B.n7 585
R155 B.n281 B.n6 585
R156 B.n438 B.n6 585
R157 B.n280 B.n5 585
R158 B.n439 B.n5 585
R159 B.n279 B.n278 585
R160 B.n278 B.n4 585
R161 B.n277 B.n67 585
R162 B.n277 B.n276 585
R163 B.n266 B.n68 585
R164 B.n269 B.n68 585
R165 B.n268 B.n267 585
R166 B.n270 B.n268 585
R167 B.n265 B.n72 585
R168 B.n75 B.n72 585
R169 B.n264 B.n263 585
R170 B.n263 B.n262 585
R171 B.n74 B.n73 585
R172 B.n255 B.n74 585
R173 B.n254 B.n253 585
R174 B.n256 B.n254 585
R175 B.n252 B.n79 585
R176 B.n83 B.n79 585
R177 B.n251 B.n250 585
R178 B.n250 B.n249 585
R179 B.n81 B.n80 585
R180 B.n82 B.n81 585
R181 B.n242 B.n241 585
R182 B.n243 B.n242 585
R183 B.n240 B.n88 585
R184 B.n88 B.n87 585
R185 B.n239 B.n238 585
R186 B.n238 B.n237 585
R187 B.n90 B.n89 585
R188 B.n91 B.n90 585
R189 B.n230 B.n229 585
R190 B.n231 B.n230 585
R191 B.n228 B.n96 585
R192 B.n96 B.n95 585
R193 B.n227 B.n226 585
R194 B.n226 B.n225 585
R195 B.n222 B.n100 585
R196 B.n221 B.n220 585
R197 B.n218 B.n101 585
R198 B.n218 B.n99 585
R199 B.n217 B.n216 585
R200 B.n215 B.n214 585
R201 B.n213 B.n103 585
R202 B.n211 B.n210 585
R203 B.n209 B.n104 585
R204 B.n208 B.n207 585
R205 B.n205 B.n105 585
R206 B.n203 B.n202 585
R207 B.n201 B.n106 585
R208 B.n200 B.n199 585
R209 B.n197 B.n107 585
R210 B.n195 B.n194 585
R211 B.n193 B.n108 585
R212 B.n192 B.n191 585
R213 B.n189 B.n109 585
R214 B.n187 B.n186 585
R215 B.n184 B.n110 585
R216 B.n183 B.n182 585
R217 B.n180 B.n113 585
R218 B.n178 B.n177 585
R219 B.n176 B.n114 585
R220 B.n175 B.n174 585
R221 B.n172 B.n115 585
R222 B.n170 B.n169 585
R223 B.n168 B.n116 585
R224 B.n167 B.n166 585
R225 B.n164 B.n163 585
R226 B.n162 B.n161 585
R227 B.n160 B.n121 585
R228 B.n158 B.n157 585
R229 B.n156 B.n122 585
R230 B.n155 B.n154 585
R231 B.n152 B.n123 585
R232 B.n150 B.n149 585
R233 B.n148 B.n124 585
R234 B.n147 B.n146 585
R235 B.n144 B.n125 585
R236 B.n142 B.n141 585
R237 B.n140 B.n126 585
R238 B.n139 B.n138 585
R239 B.n136 B.n127 585
R240 B.n134 B.n133 585
R241 B.n132 B.n128 585
R242 B.n131 B.n130 585
R243 B.n98 B.n97 585
R244 B.n99 B.n98 585
R245 B.n224 B.n223 585
R246 B.n225 B.n224 585
R247 B.n94 B.n93 585
R248 B.n95 B.n94 585
R249 B.n233 B.n232 585
R250 B.n232 B.n231 585
R251 B.n234 B.n92 585
R252 B.n92 B.n91 585
R253 B.n236 B.n235 585
R254 B.n237 B.n236 585
R255 B.n86 B.n85 585
R256 B.n87 B.n86 585
R257 B.n245 B.n244 585
R258 B.n244 B.n243 585
R259 B.n246 B.n84 585
R260 B.n84 B.n82 585
R261 B.n248 B.n247 585
R262 B.n249 B.n248 585
R263 B.n78 B.n77 585
R264 B.n83 B.n78 585
R265 B.n258 B.n257 585
R266 B.n257 B.n256 585
R267 B.n259 B.n76 585
R268 B.n255 B.n76 585
R269 B.n261 B.n260 585
R270 B.n262 B.n261 585
R271 B.n71 B.n70 585
R272 B.n75 B.n71 585
R273 B.n272 B.n271 585
R274 B.n271 B.n270 585
R275 B.n273 B.n69 585
R276 B.n269 B.n69 585
R277 B.n275 B.n274 585
R278 B.n276 B.n275 585
R279 B.n3 B.n0 585
R280 B.n4 B.n3 585
R281 B.n436 B.n1 585
R282 B.n437 B.n436 585
R283 B.n435 B.n434 585
R284 B.n435 B.n8 585
R285 B.n433 B.n9 585
R286 B.n12 B.n9 585
R287 B.n432 B.n431 585
R288 B.n431 B.n430 585
R289 B.n11 B.n10 585
R290 B.n429 B.n11 585
R291 B.n427 B.n426 585
R292 B.n428 B.n427 585
R293 B.n425 B.n16 585
R294 B.n19 B.n16 585
R295 B.n424 B.n423 585
R296 B.n423 B.n422 585
R297 B.n18 B.n17 585
R298 B.n421 B.n18 585
R299 B.n419 B.n418 585
R300 B.n420 B.n419 585
R301 B.n417 B.n24 585
R302 B.n24 B.n23 585
R303 B.n416 B.n415 585
R304 B.n415 B.n414 585
R305 B.n26 B.n25 585
R306 B.n413 B.n26 585
R307 B.n411 B.n410 585
R308 B.n412 B.n411 585
R309 B.n409 B.n31 585
R310 B.n31 B.n30 585
R311 B.n408 B.n407 585
R312 B.n407 B.n406 585
R313 B.n33 B.n32 585
R314 B.n405 B.n33 585
R315 B.n403 B.n402 585
R316 B.n404 B.n403 585
R317 B.n440 B.n439 585
R318 B.n438 B.n2 585
R319 B.n403 B.n38 497.305
R320 B.n306 B.n36 497.305
R321 B.n226 B.n98 497.305
R322 B.n224 B.n100 497.305
R323 B.n49 B.t12 476.142
R324 B.n56 B.t8 476.142
R325 B.n117 B.t15 476.142
R326 B.n111 B.t19 476.142
R327 B.n307 B.n37 256.663
R328 B.n309 B.n37 256.663
R329 B.n315 B.n37 256.663
R330 B.n317 B.n37 256.663
R331 B.n323 B.n37 256.663
R332 B.n325 B.n37 256.663
R333 B.n331 B.n37 256.663
R334 B.n333 B.n37 256.663
R335 B.n339 B.n37 256.663
R336 B.n341 B.n37 256.663
R337 B.n348 B.n37 256.663
R338 B.n350 B.n37 256.663
R339 B.n356 B.n37 256.663
R340 B.n358 B.n37 256.663
R341 B.n364 B.n37 256.663
R342 B.n366 B.n37 256.663
R343 B.n372 B.n37 256.663
R344 B.n374 B.n37 256.663
R345 B.n380 B.n37 256.663
R346 B.n382 B.n37 256.663
R347 B.n388 B.n37 256.663
R348 B.n390 B.n37 256.663
R349 B.n396 B.n37 256.663
R350 B.n398 B.n37 256.663
R351 B.n219 B.n99 256.663
R352 B.n102 B.n99 256.663
R353 B.n212 B.n99 256.663
R354 B.n206 B.n99 256.663
R355 B.n204 B.n99 256.663
R356 B.n198 B.n99 256.663
R357 B.n196 B.n99 256.663
R358 B.n190 B.n99 256.663
R359 B.n188 B.n99 256.663
R360 B.n181 B.n99 256.663
R361 B.n179 B.n99 256.663
R362 B.n173 B.n99 256.663
R363 B.n171 B.n99 256.663
R364 B.n165 B.n99 256.663
R365 B.n120 B.n99 256.663
R366 B.n159 B.n99 256.663
R367 B.n153 B.n99 256.663
R368 B.n151 B.n99 256.663
R369 B.n145 B.n99 256.663
R370 B.n143 B.n99 256.663
R371 B.n137 B.n99 256.663
R372 B.n135 B.n99 256.663
R373 B.n129 B.n99 256.663
R374 B.n442 B.n441 256.663
R375 B.n399 B.n397 163.367
R376 B.n395 B.n40 163.367
R377 B.n391 B.n389 163.367
R378 B.n387 B.n42 163.367
R379 B.n383 B.n381 163.367
R380 B.n379 B.n44 163.367
R381 B.n375 B.n373 163.367
R382 B.n371 B.n46 163.367
R383 B.n367 B.n365 163.367
R384 B.n363 B.n48 163.367
R385 B.n359 B.n357 163.367
R386 B.n355 B.n53 163.367
R387 B.n351 B.n349 163.367
R388 B.n347 B.n55 163.367
R389 B.n342 B.n340 163.367
R390 B.n338 B.n59 163.367
R391 B.n334 B.n332 163.367
R392 B.n330 B.n61 163.367
R393 B.n326 B.n324 163.367
R394 B.n322 B.n63 163.367
R395 B.n318 B.n316 163.367
R396 B.n314 B.n65 163.367
R397 B.n310 B.n308 163.367
R398 B.n226 B.n96 163.367
R399 B.n230 B.n96 163.367
R400 B.n230 B.n90 163.367
R401 B.n238 B.n90 163.367
R402 B.n238 B.n88 163.367
R403 B.n242 B.n88 163.367
R404 B.n242 B.n81 163.367
R405 B.n250 B.n81 163.367
R406 B.n250 B.n79 163.367
R407 B.n254 B.n79 163.367
R408 B.n254 B.n74 163.367
R409 B.n263 B.n74 163.367
R410 B.n263 B.n72 163.367
R411 B.n268 B.n72 163.367
R412 B.n268 B.n68 163.367
R413 B.n277 B.n68 163.367
R414 B.n278 B.n277 163.367
R415 B.n278 B.n5 163.367
R416 B.n6 B.n5 163.367
R417 B.n7 B.n6 163.367
R418 B.n284 B.n7 163.367
R419 B.n285 B.n284 163.367
R420 B.n285 B.n13 163.367
R421 B.n14 B.n13 163.367
R422 B.n15 B.n14 163.367
R423 B.n290 B.n15 163.367
R424 B.n290 B.n20 163.367
R425 B.n21 B.n20 163.367
R426 B.n22 B.n21 163.367
R427 B.n295 B.n22 163.367
R428 B.n295 B.n27 163.367
R429 B.n28 B.n27 163.367
R430 B.n29 B.n28 163.367
R431 B.n300 B.n29 163.367
R432 B.n300 B.n34 163.367
R433 B.n35 B.n34 163.367
R434 B.n36 B.n35 163.367
R435 B.n220 B.n218 163.367
R436 B.n218 B.n217 163.367
R437 B.n214 B.n213 163.367
R438 B.n211 B.n104 163.367
R439 B.n207 B.n205 163.367
R440 B.n203 B.n106 163.367
R441 B.n199 B.n197 163.367
R442 B.n195 B.n108 163.367
R443 B.n191 B.n189 163.367
R444 B.n187 B.n110 163.367
R445 B.n182 B.n180 163.367
R446 B.n178 B.n114 163.367
R447 B.n174 B.n172 163.367
R448 B.n170 B.n116 163.367
R449 B.n166 B.n164 163.367
R450 B.n161 B.n160 163.367
R451 B.n158 B.n122 163.367
R452 B.n154 B.n152 163.367
R453 B.n150 B.n124 163.367
R454 B.n146 B.n144 163.367
R455 B.n142 B.n126 163.367
R456 B.n138 B.n136 163.367
R457 B.n134 B.n128 163.367
R458 B.n130 B.n98 163.367
R459 B.n224 B.n94 163.367
R460 B.n232 B.n94 163.367
R461 B.n232 B.n92 163.367
R462 B.n236 B.n92 163.367
R463 B.n236 B.n86 163.367
R464 B.n244 B.n86 163.367
R465 B.n244 B.n84 163.367
R466 B.n248 B.n84 163.367
R467 B.n248 B.n78 163.367
R468 B.n257 B.n78 163.367
R469 B.n257 B.n76 163.367
R470 B.n261 B.n76 163.367
R471 B.n261 B.n71 163.367
R472 B.n271 B.n71 163.367
R473 B.n271 B.n69 163.367
R474 B.n275 B.n69 163.367
R475 B.n275 B.n3 163.367
R476 B.n440 B.n3 163.367
R477 B.n436 B.n2 163.367
R478 B.n436 B.n435 163.367
R479 B.n435 B.n9 163.367
R480 B.n431 B.n9 163.367
R481 B.n431 B.n11 163.367
R482 B.n427 B.n11 163.367
R483 B.n427 B.n16 163.367
R484 B.n423 B.n16 163.367
R485 B.n423 B.n18 163.367
R486 B.n419 B.n18 163.367
R487 B.n419 B.n24 163.367
R488 B.n415 B.n24 163.367
R489 B.n415 B.n26 163.367
R490 B.n411 B.n26 163.367
R491 B.n411 B.n31 163.367
R492 B.n407 B.n31 163.367
R493 B.n407 B.n33 163.367
R494 B.n403 B.n33 163.367
R495 B.n225 B.n99 157.226
R496 B.n404 B.n37 157.226
R497 B.n56 B.t10 89.4327
R498 B.n117 B.t18 89.4327
R499 B.n49 B.t13 89.4289
R500 B.n111 B.t21 89.4289
R501 B.n225 B.n95 78.0391
R502 B.n231 B.n95 78.0391
R503 B.n231 B.n91 78.0391
R504 B.n237 B.n91 78.0391
R505 B.n243 B.n87 78.0391
R506 B.n243 B.n82 78.0391
R507 B.n249 B.n82 78.0391
R508 B.n249 B.n83 78.0391
R509 B.n256 B.n255 78.0391
R510 B.n262 B.n75 78.0391
R511 B.n270 B.n269 78.0391
R512 B.n276 B.n4 78.0391
R513 B.n439 B.n4 78.0391
R514 B.n439 B.n438 78.0391
R515 B.n438 B.n437 78.0391
R516 B.n437 B.n8 78.0391
R517 B.n430 B.n12 78.0391
R518 B.n429 B.n428 78.0391
R519 B.n422 B.n19 78.0391
R520 B.n421 B.n420 78.0391
R521 B.n420 B.n23 78.0391
R522 B.n414 B.n23 78.0391
R523 B.n414 B.n413 78.0391
R524 B.n412 B.n30 78.0391
R525 B.n406 B.n30 78.0391
R526 B.n406 B.n405 78.0391
R527 B.n405 B.n404 78.0391
R528 B.n57 B.t11 75.4691
R529 B.n118 B.t17 75.4691
R530 B.n50 B.t14 75.4652
R531 B.n112 B.t20 75.4652
R532 B.n398 B.n38 71.676
R533 B.n397 B.n396 71.676
R534 B.n390 B.n40 71.676
R535 B.n389 B.n388 71.676
R536 B.n382 B.n42 71.676
R537 B.n381 B.n380 71.676
R538 B.n374 B.n44 71.676
R539 B.n373 B.n372 71.676
R540 B.n366 B.n46 71.676
R541 B.n365 B.n364 71.676
R542 B.n358 B.n48 71.676
R543 B.n357 B.n356 71.676
R544 B.n350 B.n53 71.676
R545 B.n349 B.n348 71.676
R546 B.n341 B.n55 71.676
R547 B.n340 B.n339 71.676
R548 B.n333 B.n59 71.676
R549 B.n332 B.n331 71.676
R550 B.n325 B.n61 71.676
R551 B.n324 B.n323 71.676
R552 B.n317 B.n63 71.676
R553 B.n316 B.n315 71.676
R554 B.n309 B.n65 71.676
R555 B.n308 B.n307 71.676
R556 B.n307 B.n306 71.676
R557 B.n310 B.n309 71.676
R558 B.n315 B.n314 71.676
R559 B.n318 B.n317 71.676
R560 B.n323 B.n322 71.676
R561 B.n326 B.n325 71.676
R562 B.n331 B.n330 71.676
R563 B.n334 B.n333 71.676
R564 B.n339 B.n338 71.676
R565 B.n342 B.n341 71.676
R566 B.n348 B.n347 71.676
R567 B.n351 B.n350 71.676
R568 B.n356 B.n355 71.676
R569 B.n359 B.n358 71.676
R570 B.n364 B.n363 71.676
R571 B.n367 B.n366 71.676
R572 B.n372 B.n371 71.676
R573 B.n375 B.n374 71.676
R574 B.n380 B.n379 71.676
R575 B.n383 B.n382 71.676
R576 B.n388 B.n387 71.676
R577 B.n391 B.n390 71.676
R578 B.n396 B.n395 71.676
R579 B.n399 B.n398 71.676
R580 B.n219 B.n100 71.676
R581 B.n217 B.n102 71.676
R582 B.n213 B.n212 71.676
R583 B.n206 B.n104 71.676
R584 B.n205 B.n204 71.676
R585 B.n198 B.n106 71.676
R586 B.n197 B.n196 71.676
R587 B.n190 B.n108 71.676
R588 B.n189 B.n188 71.676
R589 B.n181 B.n110 71.676
R590 B.n180 B.n179 71.676
R591 B.n173 B.n114 71.676
R592 B.n172 B.n171 71.676
R593 B.n165 B.n116 71.676
R594 B.n164 B.n120 71.676
R595 B.n160 B.n159 71.676
R596 B.n153 B.n122 71.676
R597 B.n152 B.n151 71.676
R598 B.n145 B.n124 71.676
R599 B.n144 B.n143 71.676
R600 B.n137 B.n126 71.676
R601 B.n136 B.n135 71.676
R602 B.n129 B.n128 71.676
R603 B.n220 B.n219 71.676
R604 B.n214 B.n102 71.676
R605 B.n212 B.n211 71.676
R606 B.n207 B.n206 71.676
R607 B.n204 B.n203 71.676
R608 B.n199 B.n198 71.676
R609 B.n196 B.n195 71.676
R610 B.n191 B.n190 71.676
R611 B.n188 B.n187 71.676
R612 B.n182 B.n181 71.676
R613 B.n179 B.n178 71.676
R614 B.n174 B.n173 71.676
R615 B.n171 B.n170 71.676
R616 B.n166 B.n165 71.676
R617 B.n161 B.n120 71.676
R618 B.n159 B.n158 71.676
R619 B.n154 B.n153 71.676
R620 B.n151 B.n150 71.676
R621 B.n146 B.n145 71.676
R622 B.n143 B.n142 71.676
R623 B.n138 B.n137 71.676
R624 B.n135 B.n134 71.676
R625 B.n130 B.n129 71.676
R626 B.n441 B.n440 71.676
R627 B.n441 B.n2 71.676
R628 B.t16 B.n87 65.4152
R629 B.n269 B.t0 65.4152
R630 B.n12 B.t7 65.4152
R631 B.n413 B.t9 65.4152
R632 B.n51 B.n50 59.5399
R633 B.n344 B.n57 59.5399
R634 B.n119 B.n118 59.5399
R635 B.n185 B.n112 59.5399
R636 B.n75 B.t1 56.2342
R637 B.t3 B.n429 56.2342
R638 B.n255 B.t5 47.0532
R639 B.n19 B.t4 47.0532
R640 B.n256 B.t2 40.1674
R641 B.n422 B.t6 40.1674
R642 B.n83 B.t2 37.8722
R643 B.t6 B.n421 37.8722
R644 B.n223 B.n222 32.3127
R645 B.n227 B.n97 32.3127
R646 B.n305 B.n304 32.3127
R647 B.n402 B.n401 32.3127
R648 B.n262 B.t5 30.9864
R649 B.n428 B.t4 30.9864
R650 B.n270 B.t1 21.8054
R651 B.n430 B.t3 21.8054
R652 B B.n442 18.0485
R653 B.n50 B.n49 13.9641
R654 B.n57 B.n56 13.9641
R655 B.n118 B.n117 13.9641
R656 B.n112 B.n111 13.9641
R657 B.n237 B.t16 12.6244
R658 B.n276 B.t0 12.6244
R659 B.t7 B.n8 12.6244
R660 B.t9 B.n412 12.6244
R661 B.n223 B.n93 10.6151
R662 B.n233 B.n93 10.6151
R663 B.n234 B.n233 10.6151
R664 B.n235 B.n234 10.6151
R665 B.n235 B.n85 10.6151
R666 B.n245 B.n85 10.6151
R667 B.n246 B.n245 10.6151
R668 B.n247 B.n246 10.6151
R669 B.n247 B.n77 10.6151
R670 B.n258 B.n77 10.6151
R671 B.n259 B.n258 10.6151
R672 B.n260 B.n259 10.6151
R673 B.n260 B.n70 10.6151
R674 B.n272 B.n70 10.6151
R675 B.n273 B.n272 10.6151
R676 B.n274 B.n273 10.6151
R677 B.n274 B.n0 10.6151
R678 B.n222 B.n221 10.6151
R679 B.n221 B.n101 10.6151
R680 B.n216 B.n101 10.6151
R681 B.n216 B.n215 10.6151
R682 B.n215 B.n103 10.6151
R683 B.n210 B.n103 10.6151
R684 B.n210 B.n209 10.6151
R685 B.n209 B.n208 10.6151
R686 B.n208 B.n105 10.6151
R687 B.n202 B.n105 10.6151
R688 B.n202 B.n201 10.6151
R689 B.n201 B.n200 10.6151
R690 B.n200 B.n107 10.6151
R691 B.n194 B.n107 10.6151
R692 B.n194 B.n193 10.6151
R693 B.n193 B.n192 10.6151
R694 B.n192 B.n109 10.6151
R695 B.n186 B.n109 10.6151
R696 B.n184 B.n183 10.6151
R697 B.n183 B.n113 10.6151
R698 B.n177 B.n113 10.6151
R699 B.n177 B.n176 10.6151
R700 B.n176 B.n175 10.6151
R701 B.n175 B.n115 10.6151
R702 B.n169 B.n115 10.6151
R703 B.n169 B.n168 10.6151
R704 B.n168 B.n167 10.6151
R705 B.n163 B.n162 10.6151
R706 B.n162 B.n121 10.6151
R707 B.n157 B.n121 10.6151
R708 B.n157 B.n156 10.6151
R709 B.n156 B.n155 10.6151
R710 B.n155 B.n123 10.6151
R711 B.n149 B.n123 10.6151
R712 B.n149 B.n148 10.6151
R713 B.n148 B.n147 10.6151
R714 B.n147 B.n125 10.6151
R715 B.n141 B.n125 10.6151
R716 B.n141 B.n140 10.6151
R717 B.n140 B.n139 10.6151
R718 B.n139 B.n127 10.6151
R719 B.n133 B.n127 10.6151
R720 B.n133 B.n132 10.6151
R721 B.n132 B.n131 10.6151
R722 B.n131 B.n97 10.6151
R723 B.n228 B.n227 10.6151
R724 B.n229 B.n228 10.6151
R725 B.n229 B.n89 10.6151
R726 B.n239 B.n89 10.6151
R727 B.n240 B.n239 10.6151
R728 B.n241 B.n240 10.6151
R729 B.n241 B.n80 10.6151
R730 B.n251 B.n80 10.6151
R731 B.n252 B.n251 10.6151
R732 B.n253 B.n252 10.6151
R733 B.n253 B.n73 10.6151
R734 B.n264 B.n73 10.6151
R735 B.n265 B.n264 10.6151
R736 B.n267 B.n265 10.6151
R737 B.n267 B.n266 10.6151
R738 B.n266 B.n67 10.6151
R739 B.n279 B.n67 10.6151
R740 B.n280 B.n279 10.6151
R741 B.n281 B.n280 10.6151
R742 B.n282 B.n281 10.6151
R743 B.n283 B.n282 10.6151
R744 B.n286 B.n283 10.6151
R745 B.n287 B.n286 10.6151
R746 B.n288 B.n287 10.6151
R747 B.n289 B.n288 10.6151
R748 B.n291 B.n289 10.6151
R749 B.n292 B.n291 10.6151
R750 B.n293 B.n292 10.6151
R751 B.n294 B.n293 10.6151
R752 B.n296 B.n294 10.6151
R753 B.n297 B.n296 10.6151
R754 B.n298 B.n297 10.6151
R755 B.n299 B.n298 10.6151
R756 B.n301 B.n299 10.6151
R757 B.n302 B.n301 10.6151
R758 B.n303 B.n302 10.6151
R759 B.n304 B.n303 10.6151
R760 B.n434 B.n1 10.6151
R761 B.n434 B.n433 10.6151
R762 B.n433 B.n432 10.6151
R763 B.n432 B.n10 10.6151
R764 B.n426 B.n10 10.6151
R765 B.n426 B.n425 10.6151
R766 B.n425 B.n424 10.6151
R767 B.n424 B.n17 10.6151
R768 B.n418 B.n17 10.6151
R769 B.n418 B.n417 10.6151
R770 B.n417 B.n416 10.6151
R771 B.n416 B.n25 10.6151
R772 B.n410 B.n25 10.6151
R773 B.n410 B.n409 10.6151
R774 B.n409 B.n408 10.6151
R775 B.n408 B.n32 10.6151
R776 B.n402 B.n32 10.6151
R777 B.n401 B.n400 10.6151
R778 B.n400 B.n39 10.6151
R779 B.n394 B.n39 10.6151
R780 B.n394 B.n393 10.6151
R781 B.n393 B.n392 10.6151
R782 B.n392 B.n41 10.6151
R783 B.n386 B.n41 10.6151
R784 B.n386 B.n385 10.6151
R785 B.n385 B.n384 10.6151
R786 B.n384 B.n43 10.6151
R787 B.n378 B.n43 10.6151
R788 B.n378 B.n377 10.6151
R789 B.n377 B.n376 10.6151
R790 B.n376 B.n45 10.6151
R791 B.n370 B.n45 10.6151
R792 B.n370 B.n369 10.6151
R793 B.n369 B.n368 10.6151
R794 B.n368 B.n47 10.6151
R795 B.n362 B.n361 10.6151
R796 B.n361 B.n360 10.6151
R797 B.n360 B.n52 10.6151
R798 B.n354 B.n52 10.6151
R799 B.n354 B.n353 10.6151
R800 B.n353 B.n352 10.6151
R801 B.n352 B.n54 10.6151
R802 B.n346 B.n54 10.6151
R803 B.n346 B.n345 10.6151
R804 B.n343 B.n58 10.6151
R805 B.n337 B.n58 10.6151
R806 B.n337 B.n336 10.6151
R807 B.n336 B.n335 10.6151
R808 B.n335 B.n60 10.6151
R809 B.n329 B.n60 10.6151
R810 B.n329 B.n328 10.6151
R811 B.n328 B.n327 10.6151
R812 B.n327 B.n62 10.6151
R813 B.n321 B.n62 10.6151
R814 B.n321 B.n320 10.6151
R815 B.n320 B.n319 10.6151
R816 B.n319 B.n64 10.6151
R817 B.n313 B.n64 10.6151
R818 B.n313 B.n312 10.6151
R819 B.n312 B.n311 10.6151
R820 B.n311 B.n66 10.6151
R821 B.n305 B.n66 10.6151
R822 B.n186 B.n185 9.36635
R823 B.n163 B.n119 9.36635
R824 B.n51 B.n47 9.36635
R825 B.n344 B.n343 9.36635
R826 B.n442 B.n0 8.11757
R827 B.n442 B.n1 8.11757
R828 B.n185 B.n184 1.24928
R829 B.n167 B.n119 1.24928
R830 B.n362 B.n51 1.24928
R831 B.n345 B.n344 1.24928
R832 VP.n3 VP.t3 400.493
R833 VP.n12 VP.t1 387.399
R834 VP.n1 VP.t4 387.399
R835 VP.n6 VP.t5 387.399
R836 VP.n10 VP.t7 367.68
R837 VP.n11 VP.t0 367.68
R838 VP.n5 VP.t2 367.68
R839 VP.n4 VP.t6 367.68
R840 VP.n13 VP.n12 161.3
R841 VP.n5 VP.n2 161.3
R842 VP.n7 VP.n6 161.3
R843 VP.n11 VP.n0 161.3
R844 VP.n10 VP.n9 161.3
R845 VP.n8 VP.n1 161.3
R846 VP.n3 VP.n2 74.3446
R847 VP.n11 VP.n10 48.2005
R848 VP.n5 VP.n4 48.2005
R849 VP.n8 VP.n7 34.8566
R850 VP.n10 VP.n1 28.4823
R851 VP.n12 VP.n11 28.4823
R852 VP.n6 VP.n5 28.4823
R853 VP.n4 VP.n3 13.0795
R854 VP.n7 VP.n2 0.189894
R855 VP.n9 VP.n8 0.189894
R856 VP.n9 VP.n0 0.189894
R857 VP.n13 VP.n0 0.189894
R858 VP VP.n13 0.0516364
R859 VDD1 VDD1.n0 74.4203
R860 VDD1.n3 VDD1.n2 74.3065
R861 VDD1.n3 VDD1.n1 74.3065
R862 VDD1.n5 VDD1.n4 74.0516
R863 VDD1.n5 VDD1.n3 30.8069
R864 VDD1.n4 VDD1.t5 4.59447
R865 VDD1.n4 VDD1.t2 4.59447
R866 VDD1.n0 VDD1.t4 4.59447
R867 VDD1.n0 VDD1.t1 4.59447
R868 VDD1.n2 VDD1.t7 4.59447
R869 VDD1.n2 VDD1.t6 4.59447
R870 VDD1.n1 VDD1.t3 4.59447
R871 VDD1.n1 VDD1.t0 4.59447
R872 VDD1 VDD1.n5 0.252655
C0 VP VDD2 0.288475f
C1 VP VDD1 1.78966f
C2 VDD2 VDD1 0.671967f
C3 VP VTAIL 1.64743f
C4 VP VN 3.53774f
C5 VDD2 VTAIL 6.44378f
C6 VDD2 VN 1.65316f
C7 VDD1 VTAIL 6.40418f
C8 VDD1 VN 0.151395f
C9 VN VTAIL 1.63332f
C10 VDD2 B 2.495482f
C11 VDD1 B 2.692564f
C12 VTAIL B 4.230626f
C13 VN B 5.713959f
C14 VP B 4.783612f
C15 VDD1.t4 B 0.0791f
C16 VDD1.t1 B 0.0791f
C17 VDD1.n0 B 0.630776f
C18 VDD1.t3 B 0.0791f
C19 VDD1.t0 B 0.0791f
C20 VDD1.n1 B 0.630348f
C21 VDD1.t7 B 0.0791f
C22 VDD1.t6 B 0.0791f
C23 VDD1.n2 B 0.630348f
C24 VDD1.n3 B 1.46018f
C25 VDD1.t5 B 0.0791f
C26 VDD1.t2 B 0.0791f
C27 VDD1.n4 B 0.629458f
C28 VDD1.n5 B 1.4753f
C29 VP.n0 B 0.027284f
C30 VP.t4 B 0.138349f
C31 VP.n1 B 0.070707f
C32 VP.n2 B 0.0909f
C33 VP.t2 B 0.134889f
C34 VP.t6 B 0.134889f
C35 VP.t3 B 0.140662f
C36 VP.n3 B 0.0686f
C37 VP.n4 B 0.075177f
C38 VP.n5 B 0.075177f
C39 VP.t5 B 0.138349f
C40 VP.n6 B 0.070707f
C41 VP.n7 B 0.80658f
C42 VP.n8 B 0.834718f
C43 VP.n9 B 0.027284f
C44 VP.t7 B 0.134889f
C45 VP.n10 B 0.075177f
C46 VP.t0 B 0.134889f
C47 VP.n11 B 0.075177f
C48 VP.t1 B 0.138349f
C49 VP.n12 B 0.070707f
C50 VP.n13 B 0.021144f
C51 VTAIL.t13 B 0.066767f
C52 VTAIL.t12 B 0.066767f
C53 VTAIL.n0 B 0.487671f
C54 VTAIL.n1 B 0.213742f
C55 VTAIL.t9 B 0.625058f
C56 VTAIL.n2 B 0.284448f
C57 VTAIL.t0 B 0.625058f
C58 VTAIL.n3 B 0.284448f
C59 VTAIL.t5 B 0.066767f
C60 VTAIL.t1 B 0.066767f
C61 VTAIL.n4 B 0.487671f
C62 VTAIL.n5 B 0.249273f
C63 VTAIL.t2 B 0.625058f
C64 VTAIL.n6 B 0.794959f
C65 VTAIL.t14 B 0.62506f
C66 VTAIL.n7 B 0.794957f
C67 VTAIL.t10 B 0.066767f
C68 VTAIL.t15 B 0.066767f
C69 VTAIL.n8 B 0.487673f
C70 VTAIL.n9 B 0.249271f
C71 VTAIL.t11 B 0.62506f
C72 VTAIL.n10 B 0.284445f
C73 VTAIL.t7 B 0.62506f
C74 VTAIL.n11 B 0.284445f
C75 VTAIL.t3 B 0.066767f
C76 VTAIL.t4 B 0.066767f
C77 VTAIL.n12 B 0.487673f
C78 VTAIL.n13 B 0.249271f
C79 VTAIL.t6 B 0.625058f
C80 VTAIL.n14 B 0.794959f
C81 VTAIL.t8 B 0.625058f
C82 VTAIL.n15 B 0.791284f
C83 VDD2.t7 B 0.080174f
C84 VDD2.t0 B 0.080174f
C85 VDD2.n0 B 0.638912f
C86 VDD2.t5 B 0.080174f
C87 VDD2.t6 B 0.080174f
C88 VDD2.n1 B 0.638912f
C89 VDD2.n2 B 1.4293f
C90 VDD2.t1 B 0.080174f
C91 VDD2.t3 B 0.080174f
C92 VDD2.n3 B 0.638012f
C93 VDD2.n4 B 1.46794f
C94 VDD2.t4 B 0.080174f
C95 VDD2.t2 B 0.080174f
C96 VDD2.n5 B 0.638893f
C97 VN.n0 B 0.089915f
C98 VN.t6 B 0.139138f
C99 VN.n1 B 0.067856f
C100 VN.t2 B 0.133427f
C101 VN.n2 B 0.074362f
C102 VN.t3 B 0.133427f
C103 VN.n3 B 0.074362f
C104 VN.t7 B 0.13685f
C105 VN.n4 B 0.069941f
C106 VN.n5 B 0.020915f
C107 VN.n6 B 0.089915f
C108 VN.t1 B 0.13685f
C109 VN.t0 B 0.133427f
C110 VN.t4 B 0.139138f
C111 VN.n7 B 0.067856f
C112 VN.n8 B 0.074362f
C113 VN.t5 B 0.133427f
C114 VN.n9 B 0.074362f
C115 VN.n10 B 0.069941f
C116 VN.n11 B 0.815782f
.ends

