* NGSPICE file created from diff_pair_sample_0287.ext - technology: sky130A

.subckt diff_pair_sample_0287 VTAIL VN VP B VDD2 VDD1
X0 B.t16 B.t14 B.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=0 ps=0 w=10.85 l=2.6
X1 VDD1.t3 VP.t0 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.79025 pd=11.18 as=4.2315 ps=22.48 w=10.85 l=2.6
X2 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=0 ps=0 w=10.85 l=2.6
X3 VDD1.t2 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.79025 pd=11.18 as=4.2315 ps=22.48 w=10.85 l=2.6
X4 VTAIL.t0 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=1.79025 ps=11.18 w=10.85 l=2.6
X5 VTAIL.t4 VP.t2 VDD1.t1 B.t17 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=1.79025 ps=11.18 w=10.85 l=2.6
X6 VTAIL.t3 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=1.79025 ps=11.18 w=10.85 l=2.6
X7 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=0 ps=0 w=10.85 l=2.6
X8 VDD2.t2 VN.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.79025 pd=11.18 as=4.2315 ps=22.48 w=10.85 l=2.6
X9 VTAIL.t7 VN.t2 VDD2.t1 B.t17 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=1.79025 ps=11.18 w=10.85 l=2.6
X10 B.t6 B.t3 B.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2315 pd=22.48 as=0 ps=0 w=10.85 l=2.6
X11 VDD2.t0 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.79025 pd=11.18 as=4.2315 ps=22.48 w=10.85 l=2.6
R0 B.n547 B.n546 585
R1 B.n548 B.n113 585
R2 B.n550 B.n549 585
R3 B.n552 B.n112 585
R4 B.n555 B.n554 585
R5 B.n556 B.n111 585
R6 B.n558 B.n557 585
R7 B.n560 B.n110 585
R8 B.n563 B.n562 585
R9 B.n564 B.n109 585
R10 B.n566 B.n565 585
R11 B.n568 B.n108 585
R12 B.n571 B.n570 585
R13 B.n572 B.n107 585
R14 B.n574 B.n573 585
R15 B.n576 B.n106 585
R16 B.n579 B.n578 585
R17 B.n580 B.n105 585
R18 B.n582 B.n581 585
R19 B.n584 B.n104 585
R20 B.n587 B.n586 585
R21 B.n588 B.n103 585
R22 B.n590 B.n589 585
R23 B.n592 B.n102 585
R24 B.n595 B.n594 585
R25 B.n596 B.n101 585
R26 B.n598 B.n597 585
R27 B.n600 B.n100 585
R28 B.n603 B.n602 585
R29 B.n604 B.n99 585
R30 B.n606 B.n605 585
R31 B.n608 B.n98 585
R32 B.n611 B.n610 585
R33 B.n612 B.n97 585
R34 B.n614 B.n613 585
R35 B.n616 B.n96 585
R36 B.n618 B.n617 585
R37 B.n620 B.n619 585
R38 B.n623 B.n622 585
R39 B.n624 B.n91 585
R40 B.n626 B.n625 585
R41 B.n628 B.n90 585
R42 B.n631 B.n630 585
R43 B.n632 B.n89 585
R44 B.n634 B.n633 585
R45 B.n636 B.n88 585
R46 B.n638 B.n637 585
R47 B.n640 B.n639 585
R48 B.n643 B.n642 585
R49 B.n644 B.n83 585
R50 B.n646 B.n645 585
R51 B.n648 B.n82 585
R52 B.n651 B.n650 585
R53 B.n652 B.n81 585
R54 B.n654 B.n653 585
R55 B.n656 B.n80 585
R56 B.n659 B.n658 585
R57 B.n660 B.n79 585
R58 B.n662 B.n661 585
R59 B.n664 B.n78 585
R60 B.n667 B.n666 585
R61 B.n668 B.n77 585
R62 B.n670 B.n669 585
R63 B.n672 B.n76 585
R64 B.n675 B.n674 585
R65 B.n676 B.n75 585
R66 B.n678 B.n677 585
R67 B.n680 B.n74 585
R68 B.n683 B.n682 585
R69 B.n684 B.n73 585
R70 B.n686 B.n685 585
R71 B.n688 B.n72 585
R72 B.n691 B.n690 585
R73 B.n692 B.n71 585
R74 B.n694 B.n693 585
R75 B.n696 B.n70 585
R76 B.n699 B.n698 585
R77 B.n700 B.n69 585
R78 B.n702 B.n701 585
R79 B.n704 B.n68 585
R80 B.n707 B.n706 585
R81 B.n708 B.n67 585
R82 B.n710 B.n709 585
R83 B.n712 B.n66 585
R84 B.n715 B.n714 585
R85 B.n716 B.n65 585
R86 B.n544 B.n63 585
R87 B.n719 B.n63 585
R88 B.n543 B.n62 585
R89 B.n720 B.n62 585
R90 B.n542 B.n61 585
R91 B.n721 B.n61 585
R92 B.n541 B.n540 585
R93 B.n540 B.n57 585
R94 B.n539 B.n56 585
R95 B.n727 B.n56 585
R96 B.n538 B.n55 585
R97 B.n728 B.n55 585
R98 B.n537 B.n54 585
R99 B.n729 B.n54 585
R100 B.n536 B.n535 585
R101 B.n535 B.n53 585
R102 B.n534 B.n49 585
R103 B.n735 B.n49 585
R104 B.n533 B.n48 585
R105 B.n736 B.n48 585
R106 B.n532 B.n47 585
R107 B.n737 B.n47 585
R108 B.n531 B.n530 585
R109 B.n530 B.n43 585
R110 B.n529 B.n42 585
R111 B.n743 B.n42 585
R112 B.n528 B.n41 585
R113 B.n744 B.n41 585
R114 B.n527 B.n40 585
R115 B.n745 B.n40 585
R116 B.n526 B.n525 585
R117 B.n525 B.n36 585
R118 B.n524 B.n35 585
R119 B.n751 B.n35 585
R120 B.n523 B.n34 585
R121 B.n752 B.n34 585
R122 B.n522 B.n33 585
R123 B.n753 B.n33 585
R124 B.n521 B.n520 585
R125 B.n520 B.n32 585
R126 B.n519 B.n28 585
R127 B.n759 B.n28 585
R128 B.n518 B.n27 585
R129 B.n760 B.n27 585
R130 B.n517 B.n26 585
R131 B.n761 B.n26 585
R132 B.n516 B.n515 585
R133 B.n515 B.n22 585
R134 B.n514 B.n21 585
R135 B.n767 B.n21 585
R136 B.n513 B.n20 585
R137 B.n768 B.n20 585
R138 B.n512 B.n19 585
R139 B.n769 B.n19 585
R140 B.n511 B.n510 585
R141 B.n510 B.n15 585
R142 B.n509 B.n14 585
R143 B.n775 B.n14 585
R144 B.n508 B.n13 585
R145 B.n776 B.n13 585
R146 B.n507 B.n12 585
R147 B.n777 B.n12 585
R148 B.n506 B.n505 585
R149 B.n505 B.n8 585
R150 B.n504 B.n7 585
R151 B.n783 B.n7 585
R152 B.n503 B.n6 585
R153 B.n784 B.n6 585
R154 B.n502 B.n5 585
R155 B.n785 B.n5 585
R156 B.n501 B.n500 585
R157 B.n500 B.n4 585
R158 B.n499 B.n114 585
R159 B.n499 B.n498 585
R160 B.n489 B.n115 585
R161 B.n116 B.n115 585
R162 B.n491 B.n490 585
R163 B.n492 B.n491 585
R164 B.n488 B.n121 585
R165 B.n121 B.n120 585
R166 B.n487 B.n486 585
R167 B.n486 B.n485 585
R168 B.n123 B.n122 585
R169 B.n124 B.n123 585
R170 B.n478 B.n477 585
R171 B.n479 B.n478 585
R172 B.n476 B.n129 585
R173 B.n129 B.n128 585
R174 B.n475 B.n474 585
R175 B.n474 B.n473 585
R176 B.n131 B.n130 585
R177 B.n132 B.n131 585
R178 B.n466 B.n465 585
R179 B.n467 B.n466 585
R180 B.n464 B.n137 585
R181 B.n137 B.n136 585
R182 B.n463 B.n462 585
R183 B.n462 B.n461 585
R184 B.n139 B.n138 585
R185 B.n454 B.n139 585
R186 B.n453 B.n452 585
R187 B.n455 B.n453 585
R188 B.n451 B.n144 585
R189 B.n144 B.n143 585
R190 B.n450 B.n449 585
R191 B.n449 B.n448 585
R192 B.n146 B.n145 585
R193 B.n147 B.n146 585
R194 B.n441 B.n440 585
R195 B.n442 B.n441 585
R196 B.n439 B.n152 585
R197 B.n152 B.n151 585
R198 B.n438 B.n437 585
R199 B.n437 B.n436 585
R200 B.n154 B.n153 585
R201 B.n155 B.n154 585
R202 B.n429 B.n428 585
R203 B.n430 B.n429 585
R204 B.n427 B.n160 585
R205 B.n160 B.n159 585
R206 B.n426 B.n425 585
R207 B.n425 B.n424 585
R208 B.n162 B.n161 585
R209 B.n417 B.n162 585
R210 B.n416 B.n415 585
R211 B.n418 B.n416 585
R212 B.n414 B.n167 585
R213 B.n167 B.n166 585
R214 B.n413 B.n412 585
R215 B.n412 B.n411 585
R216 B.n169 B.n168 585
R217 B.n170 B.n169 585
R218 B.n404 B.n403 585
R219 B.n405 B.n404 585
R220 B.n402 B.n175 585
R221 B.n175 B.n174 585
R222 B.n401 B.n400 585
R223 B.n400 B.n399 585
R224 B.n396 B.n179 585
R225 B.n395 B.n394 585
R226 B.n392 B.n180 585
R227 B.n392 B.n178 585
R228 B.n391 B.n390 585
R229 B.n389 B.n388 585
R230 B.n387 B.n182 585
R231 B.n385 B.n384 585
R232 B.n383 B.n183 585
R233 B.n382 B.n381 585
R234 B.n379 B.n184 585
R235 B.n377 B.n376 585
R236 B.n375 B.n185 585
R237 B.n374 B.n373 585
R238 B.n371 B.n186 585
R239 B.n369 B.n368 585
R240 B.n367 B.n187 585
R241 B.n366 B.n365 585
R242 B.n363 B.n188 585
R243 B.n361 B.n360 585
R244 B.n359 B.n189 585
R245 B.n358 B.n357 585
R246 B.n355 B.n190 585
R247 B.n353 B.n352 585
R248 B.n351 B.n191 585
R249 B.n350 B.n349 585
R250 B.n347 B.n192 585
R251 B.n345 B.n344 585
R252 B.n343 B.n193 585
R253 B.n342 B.n341 585
R254 B.n339 B.n194 585
R255 B.n337 B.n336 585
R256 B.n335 B.n195 585
R257 B.n334 B.n333 585
R258 B.n331 B.n196 585
R259 B.n329 B.n328 585
R260 B.n327 B.n197 585
R261 B.n326 B.n325 585
R262 B.n323 B.n198 585
R263 B.n321 B.n320 585
R264 B.n319 B.n199 585
R265 B.n318 B.n317 585
R266 B.n315 B.n203 585
R267 B.n313 B.n312 585
R268 B.n311 B.n204 585
R269 B.n310 B.n309 585
R270 B.n307 B.n205 585
R271 B.n305 B.n304 585
R272 B.n303 B.n206 585
R273 B.n301 B.n300 585
R274 B.n298 B.n209 585
R275 B.n296 B.n295 585
R276 B.n294 B.n210 585
R277 B.n293 B.n292 585
R278 B.n290 B.n211 585
R279 B.n288 B.n287 585
R280 B.n286 B.n212 585
R281 B.n285 B.n284 585
R282 B.n282 B.n213 585
R283 B.n280 B.n279 585
R284 B.n278 B.n214 585
R285 B.n277 B.n276 585
R286 B.n274 B.n215 585
R287 B.n272 B.n271 585
R288 B.n270 B.n216 585
R289 B.n269 B.n268 585
R290 B.n266 B.n217 585
R291 B.n264 B.n263 585
R292 B.n262 B.n218 585
R293 B.n261 B.n260 585
R294 B.n258 B.n219 585
R295 B.n256 B.n255 585
R296 B.n254 B.n220 585
R297 B.n253 B.n252 585
R298 B.n250 B.n221 585
R299 B.n248 B.n247 585
R300 B.n246 B.n222 585
R301 B.n245 B.n244 585
R302 B.n242 B.n223 585
R303 B.n240 B.n239 585
R304 B.n238 B.n224 585
R305 B.n237 B.n236 585
R306 B.n234 B.n225 585
R307 B.n232 B.n231 585
R308 B.n230 B.n226 585
R309 B.n229 B.n228 585
R310 B.n177 B.n176 585
R311 B.n178 B.n177 585
R312 B.n398 B.n397 585
R313 B.n399 B.n398 585
R314 B.n173 B.n172 585
R315 B.n174 B.n173 585
R316 B.n407 B.n406 585
R317 B.n406 B.n405 585
R318 B.n408 B.n171 585
R319 B.n171 B.n170 585
R320 B.n410 B.n409 585
R321 B.n411 B.n410 585
R322 B.n165 B.n164 585
R323 B.n166 B.n165 585
R324 B.n420 B.n419 585
R325 B.n419 B.n418 585
R326 B.n421 B.n163 585
R327 B.n417 B.n163 585
R328 B.n423 B.n422 585
R329 B.n424 B.n423 585
R330 B.n158 B.n157 585
R331 B.n159 B.n158 585
R332 B.n432 B.n431 585
R333 B.n431 B.n430 585
R334 B.n433 B.n156 585
R335 B.n156 B.n155 585
R336 B.n435 B.n434 585
R337 B.n436 B.n435 585
R338 B.n150 B.n149 585
R339 B.n151 B.n150 585
R340 B.n444 B.n443 585
R341 B.n443 B.n442 585
R342 B.n445 B.n148 585
R343 B.n148 B.n147 585
R344 B.n447 B.n446 585
R345 B.n448 B.n447 585
R346 B.n142 B.n141 585
R347 B.n143 B.n142 585
R348 B.n457 B.n456 585
R349 B.n456 B.n455 585
R350 B.n458 B.n140 585
R351 B.n454 B.n140 585
R352 B.n460 B.n459 585
R353 B.n461 B.n460 585
R354 B.n135 B.n134 585
R355 B.n136 B.n135 585
R356 B.n469 B.n468 585
R357 B.n468 B.n467 585
R358 B.n470 B.n133 585
R359 B.n133 B.n132 585
R360 B.n472 B.n471 585
R361 B.n473 B.n472 585
R362 B.n127 B.n126 585
R363 B.n128 B.n127 585
R364 B.n481 B.n480 585
R365 B.n480 B.n479 585
R366 B.n482 B.n125 585
R367 B.n125 B.n124 585
R368 B.n484 B.n483 585
R369 B.n485 B.n484 585
R370 B.n119 B.n118 585
R371 B.n120 B.n119 585
R372 B.n494 B.n493 585
R373 B.n493 B.n492 585
R374 B.n495 B.n117 585
R375 B.n117 B.n116 585
R376 B.n497 B.n496 585
R377 B.n498 B.n497 585
R378 B.n2 B.n0 585
R379 B.n4 B.n2 585
R380 B.n3 B.n1 585
R381 B.n784 B.n3 585
R382 B.n782 B.n781 585
R383 B.n783 B.n782 585
R384 B.n780 B.n9 585
R385 B.n9 B.n8 585
R386 B.n779 B.n778 585
R387 B.n778 B.n777 585
R388 B.n11 B.n10 585
R389 B.n776 B.n11 585
R390 B.n774 B.n773 585
R391 B.n775 B.n774 585
R392 B.n772 B.n16 585
R393 B.n16 B.n15 585
R394 B.n771 B.n770 585
R395 B.n770 B.n769 585
R396 B.n18 B.n17 585
R397 B.n768 B.n18 585
R398 B.n766 B.n765 585
R399 B.n767 B.n766 585
R400 B.n764 B.n23 585
R401 B.n23 B.n22 585
R402 B.n763 B.n762 585
R403 B.n762 B.n761 585
R404 B.n25 B.n24 585
R405 B.n760 B.n25 585
R406 B.n758 B.n757 585
R407 B.n759 B.n758 585
R408 B.n756 B.n29 585
R409 B.n32 B.n29 585
R410 B.n755 B.n754 585
R411 B.n754 B.n753 585
R412 B.n31 B.n30 585
R413 B.n752 B.n31 585
R414 B.n750 B.n749 585
R415 B.n751 B.n750 585
R416 B.n748 B.n37 585
R417 B.n37 B.n36 585
R418 B.n747 B.n746 585
R419 B.n746 B.n745 585
R420 B.n39 B.n38 585
R421 B.n744 B.n39 585
R422 B.n742 B.n741 585
R423 B.n743 B.n742 585
R424 B.n740 B.n44 585
R425 B.n44 B.n43 585
R426 B.n739 B.n738 585
R427 B.n738 B.n737 585
R428 B.n46 B.n45 585
R429 B.n736 B.n46 585
R430 B.n734 B.n733 585
R431 B.n735 B.n734 585
R432 B.n732 B.n50 585
R433 B.n53 B.n50 585
R434 B.n731 B.n730 585
R435 B.n730 B.n729 585
R436 B.n52 B.n51 585
R437 B.n728 B.n52 585
R438 B.n726 B.n725 585
R439 B.n727 B.n726 585
R440 B.n724 B.n58 585
R441 B.n58 B.n57 585
R442 B.n723 B.n722 585
R443 B.n722 B.n721 585
R444 B.n60 B.n59 585
R445 B.n720 B.n60 585
R446 B.n718 B.n717 585
R447 B.n719 B.n718 585
R448 B.n787 B.n786 585
R449 B.n786 B.n785 585
R450 B.n398 B.n179 497.305
R451 B.n718 B.n65 497.305
R452 B.n400 B.n177 497.305
R453 B.n546 B.n63 497.305
R454 B.n207 B.t16 319.481
R455 B.n92 B.t9 319.481
R456 B.n200 B.t6 319.481
R457 B.n84 B.t12 319.481
R458 B.n207 B.t14 308.618
R459 B.n200 B.t3 308.618
R460 B.n84 B.t11 308.618
R461 B.n92 B.t7 308.618
R462 B.n208 B.t15 262.656
R463 B.n93 B.t10 262.656
R464 B.n201 B.t5 262.656
R465 B.n85 B.t13 262.656
R466 B.n545 B.n64 256.663
R467 B.n551 B.n64 256.663
R468 B.n553 B.n64 256.663
R469 B.n559 B.n64 256.663
R470 B.n561 B.n64 256.663
R471 B.n567 B.n64 256.663
R472 B.n569 B.n64 256.663
R473 B.n575 B.n64 256.663
R474 B.n577 B.n64 256.663
R475 B.n583 B.n64 256.663
R476 B.n585 B.n64 256.663
R477 B.n591 B.n64 256.663
R478 B.n593 B.n64 256.663
R479 B.n599 B.n64 256.663
R480 B.n601 B.n64 256.663
R481 B.n607 B.n64 256.663
R482 B.n609 B.n64 256.663
R483 B.n615 B.n64 256.663
R484 B.n95 B.n64 256.663
R485 B.n621 B.n64 256.663
R486 B.n627 B.n64 256.663
R487 B.n629 B.n64 256.663
R488 B.n635 B.n64 256.663
R489 B.n87 B.n64 256.663
R490 B.n641 B.n64 256.663
R491 B.n647 B.n64 256.663
R492 B.n649 B.n64 256.663
R493 B.n655 B.n64 256.663
R494 B.n657 B.n64 256.663
R495 B.n663 B.n64 256.663
R496 B.n665 B.n64 256.663
R497 B.n671 B.n64 256.663
R498 B.n673 B.n64 256.663
R499 B.n679 B.n64 256.663
R500 B.n681 B.n64 256.663
R501 B.n687 B.n64 256.663
R502 B.n689 B.n64 256.663
R503 B.n695 B.n64 256.663
R504 B.n697 B.n64 256.663
R505 B.n703 B.n64 256.663
R506 B.n705 B.n64 256.663
R507 B.n711 B.n64 256.663
R508 B.n713 B.n64 256.663
R509 B.n393 B.n178 256.663
R510 B.n181 B.n178 256.663
R511 B.n386 B.n178 256.663
R512 B.n380 B.n178 256.663
R513 B.n378 B.n178 256.663
R514 B.n372 B.n178 256.663
R515 B.n370 B.n178 256.663
R516 B.n364 B.n178 256.663
R517 B.n362 B.n178 256.663
R518 B.n356 B.n178 256.663
R519 B.n354 B.n178 256.663
R520 B.n348 B.n178 256.663
R521 B.n346 B.n178 256.663
R522 B.n340 B.n178 256.663
R523 B.n338 B.n178 256.663
R524 B.n332 B.n178 256.663
R525 B.n330 B.n178 256.663
R526 B.n324 B.n178 256.663
R527 B.n322 B.n178 256.663
R528 B.n316 B.n178 256.663
R529 B.n314 B.n178 256.663
R530 B.n308 B.n178 256.663
R531 B.n306 B.n178 256.663
R532 B.n299 B.n178 256.663
R533 B.n297 B.n178 256.663
R534 B.n291 B.n178 256.663
R535 B.n289 B.n178 256.663
R536 B.n283 B.n178 256.663
R537 B.n281 B.n178 256.663
R538 B.n275 B.n178 256.663
R539 B.n273 B.n178 256.663
R540 B.n267 B.n178 256.663
R541 B.n265 B.n178 256.663
R542 B.n259 B.n178 256.663
R543 B.n257 B.n178 256.663
R544 B.n251 B.n178 256.663
R545 B.n249 B.n178 256.663
R546 B.n243 B.n178 256.663
R547 B.n241 B.n178 256.663
R548 B.n235 B.n178 256.663
R549 B.n233 B.n178 256.663
R550 B.n227 B.n178 256.663
R551 B.n398 B.n173 163.367
R552 B.n406 B.n173 163.367
R553 B.n406 B.n171 163.367
R554 B.n410 B.n171 163.367
R555 B.n410 B.n165 163.367
R556 B.n419 B.n165 163.367
R557 B.n419 B.n163 163.367
R558 B.n423 B.n163 163.367
R559 B.n423 B.n158 163.367
R560 B.n431 B.n158 163.367
R561 B.n431 B.n156 163.367
R562 B.n435 B.n156 163.367
R563 B.n435 B.n150 163.367
R564 B.n443 B.n150 163.367
R565 B.n443 B.n148 163.367
R566 B.n447 B.n148 163.367
R567 B.n447 B.n142 163.367
R568 B.n456 B.n142 163.367
R569 B.n456 B.n140 163.367
R570 B.n460 B.n140 163.367
R571 B.n460 B.n135 163.367
R572 B.n468 B.n135 163.367
R573 B.n468 B.n133 163.367
R574 B.n472 B.n133 163.367
R575 B.n472 B.n127 163.367
R576 B.n480 B.n127 163.367
R577 B.n480 B.n125 163.367
R578 B.n484 B.n125 163.367
R579 B.n484 B.n119 163.367
R580 B.n493 B.n119 163.367
R581 B.n493 B.n117 163.367
R582 B.n497 B.n117 163.367
R583 B.n497 B.n2 163.367
R584 B.n786 B.n2 163.367
R585 B.n786 B.n3 163.367
R586 B.n782 B.n3 163.367
R587 B.n782 B.n9 163.367
R588 B.n778 B.n9 163.367
R589 B.n778 B.n11 163.367
R590 B.n774 B.n11 163.367
R591 B.n774 B.n16 163.367
R592 B.n770 B.n16 163.367
R593 B.n770 B.n18 163.367
R594 B.n766 B.n18 163.367
R595 B.n766 B.n23 163.367
R596 B.n762 B.n23 163.367
R597 B.n762 B.n25 163.367
R598 B.n758 B.n25 163.367
R599 B.n758 B.n29 163.367
R600 B.n754 B.n29 163.367
R601 B.n754 B.n31 163.367
R602 B.n750 B.n31 163.367
R603 B.n750 B.n37 163.367
R604 B.n746 B.n37 163.367
R605 B.n746 B.n39 163.367
R606 B.n742 B.n39 163.367
R607 B.n742 B.n44 163.367
R608 B.n738 B.n44 163.367
R609 B.n738 B.n46 163.367
R610 B.n734 B.n46 163.367
R611 B.n734 B.n50 163.367
R612 B.n730 B.n50 163.367
R613 B.n730 B.n52 163.367
R614 B.n726 B.n52 163.367
R615 B.n726 B.n58 163.367
R616 B.n722 B.n58 163.367
R617 B.n722 B.n60 163.367
R618 B.n718 B.n60 163.367
R619 B.n394 B.n392 163.367
R620 B.n392 B.n391 163.367
R621 B.n388 B.n387 163.367
R622 B.n385 B.n183 163.367
R623 B.n381 B.n379 163.367
R624 B.n377 B.n185 163.367
R625 B.n373 B.n371 163.367
R626 B.n369 B.n187 163.367
R627 B.n365 B.n363 163.367
R628 B.n361 B.n189 163.367
R629 B.n357 B.n355 163.367
R630 B.n353 B.n191 163.367
R631 B.n349 B.n347 163.367
R632 B.n345 B.n193 163.367
R633 B.n341 B.n339 163.367
R634 B.n337 B.n195 163.367
R635 B.n333 B.n331 163.367
R636 B.n329 B.n197 163.367
R637 B.n325 B.n323 163.367
R638 B.n321 B.n199 163.367
R639 B.n317 B.n315 163.367
R640 B.n313 B.n204 163.367
R641 B.n309 B.n307 163.367
R642 B.n305 B.n206 163.367
R643 B.n300 B.n298 163.367
R644 B.n296 B.n210 163.367
R645 B.n292 B.n290 163.367
R646 B.n288 B.n212 163.367
R647 B.n284 B.n282 163.367
R648 B.n280 B.n214 163.367
R649 B.n276 B.n274 163.367
R650 B.n272 B.n216 163.367
R651 B.n268 B.n266 163.367
R652 B.n264 B.n218 163.367
R653 B.n260 B.n258 163.367
R654 B.n256 B.n220 163.367
R655 B.n252 B.n250 163.367
R656 B.n248 B.n222 163.367
R657 B.n244 B.n242 163.367
R658 B.n240 B.n224 163.367
R659 B.n236 B.n234 163.367
R660 B.n232 B.n226 163.367
R661 B.n228 B.n177 163.367
R662 B.n400 B.n175 163.367
R663 B.n404 B.n175 163.367
R664 B.n404 B.n169 163.367
R665 B.n412 B.n169 163.367
R666 B.n412 B.n167 163.367
R667 B.n416 B.n167 163.367
R668 B.n416 B.n162 163.367
R669 B.n425 B.n162 163.367
R670 B.n425 B.n160 163.367
R671 B.n429 B.n160 163.367
R672 B.n429 B.n154 163.367
R673 B.n437 B.n154 163.367
R674 B.n437 B.n152 163.367
R675 B.n441 B.n152 163.367
R676 B.n441 B.n146 163.367
R677 B.n449 B.n146 163.367
R678 B.n449 B.n144 163.367
R679 B.n453 B.n144 163.367
R680 B.n453 B.n139 163.367
R681 B.n462 B.n139 163.367
R682 B.n462 B.n137 163.367
R683 B.n466 B.n137 163.367
R684 B.n466 B.n131 163.367
R685 B.n474 B.n131 163.367
R686 B.n474 B.n129 163.367
R687 B.n478 B.n129 163.367
R688 B.n478 B.n123 163.367
R689 B.n486 B.n123 163.367
R690 B.n486 B.n121 163.367
R691 B.n491 B.n121 163.367
R692 B.n491 B.n115 163.367
R693 B.n499 B.n115 163.367
R694 B.n500 B.n499 163.367
R695 B.n500 B.n5 163.367
R696 B.n6 B.n5 163.367
R697 B.n7 B.n6 163.367
R698 B.n505 B.n7 163.367
R699 B.n505 B.n12 163.367
R700 B.n13 B.n12 163.367
R701 B.n14 B.n13 163.367
R702 B.n510 B.n14 163.367
R703 B.n510 B.n19 163.367
R704 B.n20 B.n19 163.367
R705 B.n21 B.n20 163.367
R706 B.n515 B.n21 163.367
R707 B.n515 B.n26 163.367
R708 B.n27 B.n26 163.367
R709 B.n28 B.n27 163.367
R710 B.n520 B.n28 163.367
R711 B.n520 B.n33 163.367
R712 B.n34 B.n33 163.367
R713 B.n35 B.n34 163.367
R714 B.n525 B.n35 163.367
R715 B.n525 B.n40 163.367
R716 B.n41 B.n40 163.367
R717 B.n42 B.n41 163.367
R718 B.n530 B.n42 163.367
R719 B.n530 B.n47 163.367
R720 B.n48 B.n47 163.367
R721 B.n49 B.n48 163.367
R722 B.n535 B.n49 163.367
R723 B.n535 B.n54 163.367
R724 B.n55 B.n54 163.367
R725 B.n56 B.n55 163.367
R726 B.n540 B.n56 163.367
R727 B.n540 B.n61 163.367
R728 B.n62 B.n61 163.367
R729 B.n63 B.n62 163.367
R730 B.n714 B.n712 163.367
R731 B.n710 B.n67 163.367
R732 B.n706 B.n704 163.367
R733 B.n702 B.n69 163.367
R734 B.n698 B.n696 163.367
R735 B.n694 B.n71 163.367
R736 B.n690 B.n688 163.367
R737 B.n686 B.n73 163.367
R738 B.n682 B.n680 163.367
R739 B.n678 B.n75 163.367
R740 B.n674 B.n672 163.367
R741 B.n670 B.n77 163.367
R742 B.n666 B.n664 163.367
R743 B.n662 B.n79 163.367
R744 B.n658 B.n656 163.367
R745 B.n654 B.n81 163.367
R746 B.n650 B.n648 163.367
R747 B.n646 B.n83 163.367
R748 B.n642 B.n640 163.367
R749 B.n637 B.n636 163.367
R750 B.n634 B.n89 163.367
R751 B.n630 B.n628 163.367
R752 B.n626 B.n91 163.367
R753 B.n622 B.n620 163.367
R754 B.n617 B.n616 163.367
R755 B.n614 B.n97 163.367
R756 B.n610 B.n608 163.367
R757 B.n606 B.n99 163.367
R758 B.n602 B.n600 163.367
R759 B.n598 B.n101 163.367
R760 B.n594 B.n592 163.367
R761 B.n590 B.n103 163.367
R762 B.n586 B.n584 163.367
R763 B.n582 B.n105 163.367
R764 B.n578 B.n576 163.367
R765 B.n574 B.n107 163.367
R766 B.n570 B.n568 163.367
R767 B.n566 B.n109 163.367
R768 B.n562 B.n560 163.367
R769 B.n558 B.n111 163.367
R770 B.n554 B.n552 163.367
R771 B.n550 B.n113 163.367
R772 B.n399 B.n178 82.5431
R773 B.n719 B.n64 82.5431
R774 B.n393 B.n179 71.676
R775 B.n391 B.n181 71.676
R776 B.n387 B.n386 71.676
R777 B.n380 B.n183 71.676
R778 B.n379 B.n378 71.676
R779 B.n372 B.n185 71.676
R780 B.n371 B.n370 71.676
R781 B.n364 B.n187 71.676
R782 B.n363 B.n362 71.676
R783 B.n356 B.n189 71.676
R784 B.n355 B.n354 71.676
R785 B.n348 B.n191 71.676
R786 B.n347 B.n346 71.676
R787 B.n340 B.n193 71.676
R788 B.n339 B.n338 71.676
R789 B.n332 B.n195 71.676
R790 B.n331 B.n330 71.676
R791 B.n324 B.n197 71.676
R792 B.n323 B.n322 71.676
R793 B.n316 B.n199 71.676
R794 B.n315 B.n314 71.676
R795 B.n308 B.n204 71.676
R796 B.n307 B.n306 71.676
R797 B.n299 B.n206 71.676
R798 B.n298 B.n297 71.676
R799 B.n291 B.n210 71.676
R800 B.n290 B.n289 71.676
R801 B.n283 B.n212 71.676
R802 B.n282 B.n281 71.676
R803 B.n275 B.n214 71.676
R804 B.n274 B.n273 71.676
R805 B.n267 B.n216 71.676
R806 B.n266 B.n265 71.676
R807 B.n259 B.n218 71.676
R808 B.n258 B.n257 71.676
R809 B.n251 B.n220 71.676
R810 B.n250 B.n249 71.676
R811 B.n243 B.n222 71.676
R812 B.n242 B.n241 71.676
R813 B.n235 B.n224 71.676
R814 B.n234 B.n233 71.676
R815 B.n227 B.n226 71.676
R816 B.n713 B.n65 71.676
R817 B.n712 B.n711 71.676
R818 B.n705 B.n67 71.676
R819 B.n704 B.n703 71.676
R820 B.n697 B.n69 71.676
R821 B.n696 B.n695 71.676
R822 B.n689 B.n71 71.676
R823 B.n688 B.n687 71.676
R824 B.n681 B.n73 71.676
R825 B.n680 B.n679 71.676
R826 B.n673 B.n75 71.676
R827 B.n672 B.n671 71.676
R828 B.n665 B.n77 71.676
R829 B.n664 B.n663 71.676
R830 B.n657 B.n79 71.676
R831 B.n656 B.n655 71.676
R832 B.n649 B.n81 71.676
R833 B.n648 B.n647 71.676
R834 B.n641 B.n83 71.676
R835 B.n640 B.n87 71.676
R836 B.n636 B.n635 71.676
R837 B.n629 B.n89 71.676
R838 B.n628 B.n627 71.676
R839 B.n621 B.n91 71.676
R840 B.n620 B.n95 71.676
R841 B.n616 B.n615 71.676
R842 B.n609 B.n97 71.676
R843 B.n608 B.n607 71.676
R844 B.n601 B.n99 71.676
R845 B.n600 B.n599 71.676
R846 B.n593 B.n101 71.676
R847 B.n592 B.n591 71.676
R848 B.n585 B.n103 71.676
R849 B.n584 B.n583 71.676
R850 B.n577 B.n105 71.676
R851 B.n576 B.n575 71.676
R852 B.n569 B.n107 71.676
R853 B.n568 B.n567 71.676
R854 B.n561 B.n109 71.676
R855 B.n560 B.n559 71.676
R856 B.n553 B.n111 71.676
R857 B.n552 B.n551 71.676
R858 B.n545 B.n113 71.676
R859 B.n546 B.n545 71.676
R860 B.n551 B.n550 71.676
R861 B.n554 B.n553 71.676
R862 B.n559 B.n558 71.676
R863 B.n562 B.n561 71.676
R864 B.n567 B.n566 71.676
R865 B.n570 B.n569 71.676
R866 B.n575 B.n574 71.676
R867 B.n578 B.n577 71.676
R868 B.n583 B.n582 71.676
R869 B.n586 B.n585 71.676
R870 B.n591 B.n590 71.676
R871 B.n594 B.n593 71.676
R872 B.n599 B.n598 71.676
R873 B.n602 B.n601 71.676
R874 B.n607 B.n606 71.676
R875 B.n610 B.n609 71.676
R876 B.n615 B.n614 71.676
R877 B.n617 B.n95 71.676
R878 B.n622 B.n621 71.676
R879 B.n627 B.n626 71.676
R880 B.n630 B.n629 71.676
R881 B.n635 B.n634 71.676
R882 B.n637 B.n87 71.676
R883 B.n642 B.n641 71.676
R884 B.n647 B.n646 71.676
R885 B.n650 B.n649 71.676
R886 B.n655 B.n654 71.676
R887 B.n658 B.n657 71.676
R888 B.n663 B.n662 71.676
R889 B.n666 B.n665 71.676
R890 B.n671 B.n670 71.676
R891 B.n674 B.n673 71.676
R892 B.n679 B.n678 71.676
R893 B.n682 B.n681 71.676
R894 B.n687 B.n686 71.676
R895 B.n690 B.n689 71.676
R896 B.n695 B.n694 71.676
R897 B.n698 B.n697 71.676
R898 B.n703 B.n702 71.676
R899 B.n706 B.n705 71.676
R900 B.n711 B.n710 71.676
R901 B.n714 B.n713 71.676
R902 B.n394 B.n393 71.676
R903 B.n388 B.n181 71.676
R904 B.n386 B.n385 71.676
R905 B.n381 B.n380 71.676
R906 B.n378 B.n377 71.676
R907 B.n373 B.n372 71.676
R908 B.n370 B.n369 71.676
R909 B.n365 B.n364 71.676
R910 B.n362 B.n361 71.676
R911 B.n357 B.n356 71.676
R912 B.n354 B.n353 71.676
R913 B.n349 B.n348 71.676
R914 B.n346 B.n345 71.676
R915 B.n341 B.n340 71.676
R916 B.n338 B.n337 71.676
R917 B.n333 B.n332 71.676
R918 B.n330 B.n329 71.676
R919 B.n325 B.n324 71.676
R920 B.n322 B.n321 71.676
R921 B.n317 B.n316 71.676
R922 B.n314 B.n313 71.676
R923 B.n309 B.n308 71.676
R924 B.n306 B.n305 71.676
R925 B.n300 B.n299 71.676
R926 B.n297 B.n296 71.676
R927 B.n292 B.n291 71.676
R928 B.n289 B.n288 71.676
R929 B.n284 B.n283 71.676
R930 B.n281 B.n280 71.676
R931 B.n276 B.n275 71.676
R932 B.n273 B.n272 71.676
R933 B.n268 B.n267 71.676
R934 B.n265 B.n264 71.676
R935 B.n260 B.n259 71.676
R936 B.n257 B.n256 71.676
R937 B.n252 B.n251 71.676
R938 B.n249 B.n248 71.676
R939 B.n244 B.n243 71.676
R940 B.n241 B.n240 71.676
R941 B.n236 B.n235 71.676
R942 B.n233 B.n232 71.676
R943 B.n228 B.n227 71.676
R944 B.n302 B.n208 59.5399
R945 B.n202 B.n201 59.5399
R946 B.n86 B.n85 59.5399
R947 B.n94 B.n93 59.5399
R948 B.n208 B.n207 56.8247
R949 B.n201 B.n200 56.8247
R950 B.n85 B.n84 56.8247
R951 B.n93 B.n92 56.8247
R952 B.n399 B.n174 46.3881
R953 B.n405 B.n174 46.3881
R954 B.n405 B.n170 46.3881
R955 B.n411 B.n170 46.3881
R956 B.n411 B.n166 46.3881
R957 B.n418 B.n166 46.3881
R958 B.n418 B.n417 46.3881
R959 B.n424 B.n159 46.3881
R960 B.n430 B.n159 46.3881
R961 B.n430 B.n155 46.3881
R962 B.n436 B.n155 46.3881
R963 B.n436 B.n151 46.3881
R964 B.n442 B.n151 46.3881
R965 B.n442 B.n147 46.3881
R966 B.n448 B.n147 46.3881
R967 B.n448 B.n143 46.3881
R968 B.n455 B.n143 46.3881
R969 B.n455 B.n454 46.3881
R970 B.n461 B.n136 46.3881
R971 B.n467 B.n136 46.3881
R972 B.n467 B.n132 46.3881
R973 B.n473 B.n132 46.3881
R974 B.n473 B.n128 46.3881
R975 B.n479 B.n128 46.3881
R976 B.n479 B.n124 46.3881
R977 B.n485 B.n124 46.3881
R978 B.n492 B.n120 46.3881
R979 B.n492 B.n116 46.3881
R980 B.n498 B.n116 46.3881
R981 B.n498 B.n4 46.3881
R982 B.n785 B.n4 46.3881
R983 B.n785 B.n784 46.3881
R984 B.n784 B.n783 46.3881
R985 B.n783 B.n8 46.3881
R986 B.n777 B.n8 46.3881
R987 B.n777 B.n776 46.3881
R988 B.n775 B.n15 46.3881
R989 B.n769 B.n15 46.3881
R990 B.n769 B.n768 46.3881
R991 B.n768 B.n767 46.3881
R992 B.n767 B.n22 46.3881
R993 B.n761 B.n22 46.3881
R994 B.n761 B.n760 46.3881
R995 B.n760 B.n759 46.3881
R996 B.n753 B.n32 46.3881
R997 B.n753 B.n752 46.3881
R998 B.n752 B.n751 46.3881
R999 B.n751 B.n36 46.3881
R1000 B.n745 B.n36 46.3881
R1001 B.n745 B.n744 46.3881
R1002 B.n744 B.n743 46.3881
R1003 B.n743 B.n43 46.3881
R1004 B.n737 B.n43 46.3881
R1005 B.n737 B.n736 46.3881
R1006 B.n736 B.n735 46.3881
R1007 B.n729 B.n53 46.3881
R1008 B.n729 B.n728 46.3881
R1009 B.n728 B.n727 46.3881
R1010 B.n727 B.n57 46.3881
R1011 B.n721 B.n57 46.3881
R1012 B.n721 B.n720 46.3881
R1013 B.n720 B.n719 46.3881
R1014 B.t0 B.n120 42.2951
R1015 B.n776 B.t17 42.2951
R1016 B.n717 B.n716 32.3127
R1017 B.n547 B.n544 32.3127
R1018 B.n401 B.n176 32.3127
R1019 B.n397 B.n396 32.3127
R1020 B.n417 B.t4 30.016
R1021 B.n53 B.t8 30.016
R1022 B.n461 B.t1 24.5586
R1023 B.n759 B.t2 24.5586
R1024 B.n454 B.t1 21.83
R1025 B.n32 B.t2 21.83
R1026 B B.n787 18.0485
R1027 B.n424 B.t4 16.3726
R1028 B.n735 B.t8 16.3726
R1029 B.n716 B.n715 10.6151
R1030 B.n715 B.n66 10.6151
R1031 B.n709 B.n66 10.6151
R1032 B.n709 B.n708 10.6151
R1033 B.n708 B.n707 10.6151
R1034 B.n707 B.n68 10.6151
R1035 B.n701 B.n68 10.6151
R1036 B.n701 B.n700 10.6151
R1037 B.n700 B.n699 10.6151
R1038 B.n699 B.n70 10.6151
R1039 B.n693 B.n70 10.6151
R1040 B.n693 B.n692 10.6151
R1041 B.n692 B.n691 10.6151
R1042 B.n691 B.n72 10.6151
R1043 B.n685 B.n72 10.6151
R1044 B.n685 B.n684 10.6151
R1045 B.n684 B.n683 10.6151
R1046 B.n683 B.n74 10.6151
R1047 B.n677 B.n74 10.6151
R1048 B.n677 B.n676 10.6151
R1049 B.n676 B.n675 10.6151
R1050 B.n675 B.n76 10.6151
R1051 B.n669 B.n76 10.6151
R1052 B.n669 B.n668 10.6151
R1053 B.n668 B.n667 10.6151
R1054 B.n667 B.n78 10.6151
R1055 B.n661 B.n78 10.6151
R1056 B.n661 B.n660 10.6151
R1057 B.n660 B.n659 10.6151
R1058 B.n659 B.n80 10.6151
R1059 B.n653 B.n80 10.6151
R1060 B.n653 B.n652 10.6151
R1061 B.n652 B.n651 10.6151
R1062 B.n651 B.n82 10.6151
R1063 B.n645 B.n82 10.6151
R1064 B.n645 B.n644 10.6151
R1065 B.n644 B.n643 10.6151
R1066 B.n639 B.n638 10.6151
R1067 B.n638 B.n88 10.6151
R1068 B.n633 B.n88 10.6151
R1069 B.n633 B.n632 10.6151
R1070 B.n632 B.n631 10.6151
R1071 B.n631 B.n90 10.6151
R1072 B.n625 B.n90 10.6151
R1073 B.n625 B.n624 10.6151
R1074 B.n624 B.n623 10.6151
R1075 B.n619 B.n618 10.6151
R1076 B.n618 B.n96 10.6151
R1077 B.n613 B.n96 10.6151
R1078 B.n613 B.n612 10.6151
R1079 B.n612 B.n611 10.6151
R1080 B.n611 B.n98 10.6151
R1081 B.n605 B.n98 10.6151
R1082 B.n605 B.n604 10.6151
R1083 B.n604 B.n603 10.6151
R1084 B.n603 B.n100 10.6151
R1085 B.n597 B.n100 10.6151
R1086 B.n597 B.n596 10.6151
R1087 B.n596 B.n595 10.6151
R1088 B.n595 B.n102 10.6151
R1089 B.n589 B.n102 10.6151
R1090 B.n589 B.n588 10.6151
R1091 B.n588 B.n587 10.6151
R1092 B.n587 B.n104 10.6151
R1093 B.n581 B.n104 10.6151
R1094 B.n581 B.n580 10.6151
R1095 B.n580 B.n579 10.6151
R1096 B.n579 B.n106 10.6151
R1097 B.n573 B.n106 10.6151
R1098 B.n573 B.n572 10.6151
R1099 B.n572 B.n571 10.6151
R1100 B.n571 B.n108 10.6151
R1101 B.n565 B.n108 10.6151
R1102 B.n565 B.n564 10.6151
R1103 B.n564 B.n563 10.6151
R1104 B.n563 B.n110 10.6151
R1105 B.n557 B.n110 10.6151
R1106 B.n557 B.n556 10.6151
R1107 B.n556 B.n555 10.6151
R1108 B.n555 B.n112 10.6151
R1109 B.n549 B.n112 10.6151
R1110 B.n549 B.n548 10.6151
R1111 B.n548 B.n547 10.6151
R1112 B.n402 B.n401 10.6151
R1113 B.n403 B.n402 10.6151
R1114 B.n403 B.n168 10.6151
R1115 B.n413 B.n168 10.6151
R1116 B.n414 B.n413 10.6151
R1117 B.n415 B.n414 10.6151
R1118 B.n415 B.n161 10.6151
R1119 B.n426 B.n161 10.6151
R1120 B.n427 B.n426 10.6151
R1121 B.n428 B.n427 10.6151
R1122 B.n428 B.n153 10.6151
R1123 B.n438 B.n153 10.6151
R1124 B.n439 B.n438 10.6151
R1125 B.n440 B.n439 10.6151
R1126 B.n440 B.n145 10.6151
R1127 B.n450 B.n145 10.6151
R1128 B.n451 B.n450 10.6151
R1129 B.n452 B.n451 10.6151
R1130 B.n452 B.n138 10.6151
R1131 B.n463 B.n138 10.6151
R1132 B.n464 B.n463 10.6151
R1133 B.n465 B.n464 10.6151
R1134 B.n465 B.n130 10.6151
R1135 B.n475 B.n130 10.6151
R1136 B.n476 B.n475 10.6151
R1137 B.n477 B.n476 10.6151
R1138 B.n477 B.n122 10.6151
R1139 B.n487 B.n122 10.6151
R1140 B.n488 B.n487 10.6151
R1141 B.n490 B.n488 10.6151
R1142 B.n490 B.n489 10.6151
R1143 B.n489 B.n114 10.6151
R1144 B.n501 B.n114 10.6151
R1145 B.n502 B.n501 10.6151
R1146 B.n503 B.n502 10.6151
R1147 B.n504 B.n503 10.6151
R1148 B.n506 B.n504 10.6151
R1149 B.n507 B.n506 10.6151
R1150 B.n508 B.n507 10.6151
R1151 B.n509 B.n508 10.6151
R1152 B.n511 B.n509 10.6151
R1153 B.n512 B.n511 10.6151
R1154 B.n513 B.n512 10.6151
R1155 B.n514 B.n513 10.6151
R1156 B.n516 B.n514 10.6151
R1157 B.n517 B.n516 10.6151
R1158 B.n518 B.n517 10.6151
R1159 B.n519 B.n518 10.6151
R1160 B.n521 B.n519 10.6151
R1161 B.n522 B.n521 10.6151
R1162 B.n523 B.n522 10.6151
R1163 B.n524 B.n523 10.6151
R1164 B.n526 B.n524 10.6151
R1165 B.n527 B.n526 10.6151
R1166 B.n528 B.n527 10.6151
R1167 B.n529 B.n528 10.6151
R1168 B.n531 B.n529 10.6151
R1169 B.n532 B.n531 10.6151
R1170 B.n533 B.n532 10.6151
R1171 B.n534 B.n533 10.6151
R1172 B.n536 B.n534 10.6151
R1173 B.n537 B.n536 10.6151
R1174 B.n538 B.n537 10.6151
R1175 B.n539 B.n538 10.6151
R1176 B.n541 B.n539 10.6151
R1177 B.n542 B.n541 10.6151
R1178 B.n543 B.n542 10.6151
R1179 B.n544 B.n543 10.6151
R1180 B.n396 B.n395 10.6151
R1181 B.n395 B.n180 10.6151
R1182 B.n390 B.n180 10.6151
R1183 B.n390 B.n389 10.6151
R1184 B.n389 B.n182 10.6151
R1185 B.n384 B.n182 10.6151
R1186 B.n384 B.n383 10.6151
R1187 B.n383 B.n382 10.6151
R1188 B.n382 B.n184 10.6151
R1189 B.n376 B.n184 10.6151
R1190 B.n376 B.n375 10.6151
R1191 B.n375 B.n374 10.6151
R1192 B.n374 B.n186 10.6151
R1193 B.n368 B.n186 10.6151
R1194 B.n368 B.n367 10.6151
R1195 B.n367 B.n366 10.6151
R1196 B.n366 B.n188 10.6151
R1197 B.n360 B.n188 10.6151
R1198 B.n360 B.n359 10.6151
R1199 B.n359 B.n358 10.6151
R1200 B.n358 B.n190 10.6151
R1201 B.n352 B.n190 10.6151
R1202 B.n352 B.n351 10.6151
R1203 B.n351 B.n350 10.6151
R1204 B.n350 B.n192 10.6151
R1205 B.n344 B.n192 10.6151
R1206 B.n344 B.n343 10.6151
R1207 B.n343 B.n342 10.6151
R1208 B.n342 B.n194 10.6151
R1209 B.n336 B.n194 10.6151
R1210 B.n336 B.n335 10.6151
R1211 B.n335 B.n334 10.6151
R1212 B.n334 B.n196 10.6151
R1213 B.n328 B.n196 10.6151
R1214 B.n328 B.n327 10.6151
R1215 B.n327 B.n326 10.6151
R1216 B.n326 B.n198 10.6151
R1217 B.n320 B.n319 10.6151
R1218 B.n319 B.n318 10.6151
R1219 B.n318 B.n203 10.6151
R1220 B.n312 B.n203 10.6151
R1221 B.n312 B.n311 10.6151
R1222 B.n311 B.n310 10.6151
R1223 B.n310 B.n205 10.6151
R1224 B.n304 B.n205 10.6151
R1225 B.n304 B.n303 10.6151
R1226 B.n301 B.n209 10.6151
R1227 B.n295 B.n209 10.6151
R1228 B.n295 B.n294 10.6151
R1229 B.n294 B.n293 10.6151
R1230 B.n293 B.n211 10.6151
R1231 B.n287 B.n211 10.6151
R1232 B.n287 B.n286 10.6151
R1233 B.n286 B.n285 10.6151
R1234 B.n285 B.n213 10.6151
R1235 B.n279 B.n213 10.6151
R1236 B.n279 B.n278 10.6151
R1237 B.n278 B.n277 10.6151
R1238 B.n277 B.n215 10.6151
R1239 B.n271 B.n215 10.6151
R1240 B.n271 B.n270 10.6151
R1241 B.n270 B.n269 10.6151
R1242 B.n269 B.n217 10.6151
R1243 B.n263 B.n217 10.6151
R1244 B.n263 B.n262 10.6151
R1245 B.n262 B.n261 10.6151
R1246 B.n261 B.n219 10.6151
R1247 B.n255 B.n219 10.6151
R1248 B.n255 B.n254 10.6151
R1249 B.n254 B.n253 10.6151
R1250 B.n253 B.n221 10.6151
R1251 B.n247 B.n221 10.6151
R1252 B.n247 B.n246 10.6151
R1253 B.n246 B.n245 10.6151
R1254 B.n245 B.n223 10.6151
R1255 B.n239 B.n223 10.6151
R1256 B.n239 B.n238 10.6151
R1257 B.n238 B.n237 10.6151
R1258 B.n237 B.n225 10.6151
R1259 B.n231 B.n225 10.6151
R1260 B.n231 B.n230 10.6151
R1261 B.n230 B.n229 10.6151
R1262 B.n229 B.n176 10.6151
R1263 B.n397 B.n172 10.6151
R1264 B.n407 B.n172 10.6151
R1265 B.n408 B.n407 10.6151
R1266 B.n409 B.n408 10.6151
R1267 B.n409 B.n164 10.6151
R1268 B.n420 B.n164 10.6151
R1269 B.n421 B.n420 10.6151
R1270 B.n422 B.n421 10.6151
R1271 B.n422 B.n157 10.6151
R1272 B.n432 B.n157 10.6151
R1273 B.n433 B.n432 10.6151
R1274 B.n434 B.n433 10.6151
R1275 B.n434 B.n149 10.6151
R1276 B.n444 B.n149 10.6151
R1277 B.n445 B.n444 10.6151
R1278 B.n446 B.n445 10.6151
R1279 B.n446 B.n141 10.6151
R1280 B.n457 B.n141 10.6151
R1281 B.n458 B.n457 10.6151
R1282 B.n459 B.n458 10.6151
R1283 B.n459 B.n134 10.6151
R1284 B.n469 B.n134 10.6151
R1285 B.n470 B.n469 10.6151
R1286 B.n471 B.n470 10.6151
R1287 B.n471 B.n126 10.6151
R1288 B.n481 B.n126 10.6151
R1289 B.n482 B.n481 10.6151
R1290 B.n483 B.n482 10.6151
R1291 B.n483 B.n118 10.6151
R1292 B.n494 B.n118 10.6151
R1293 B.n495 B.n494 10.6151
R1294 B.n496 B.n495 10.6151
R1295 B.n496 B.n0 10.6151
R1296 B.n781 B.n1 10.6151
R1297 B.n781 B.n780 10.6151
R1298 B.n780 B.n779 10.6151
R1299 B.n779 B.n10 10.6151
R1300 B.n773 B.n10 10.6151
R1301 B.n773 B.n772 10.6151
R1302 B.n772 B.n771 10.6151
R1303 B.n771 B.n17 10.6151
R1304 B.n765 B.n17 10.6151
R1305 B.n765 B.n764 10.6151
R1306 B.n764 B.n763 10.6151
R1307 B.n763 B.n24 10.6151
R1308 B.n757 B.n24 10.6151
R1309 B.n757 B.n756 10.6151
R1310 B.n756 B.n755 10.6151
R1311 B.n755 B.n30 10.6151
R1312 B.n749 B.n30 10.6151
R1313 B.n749 B.n748 10.6151
R1314 B.n748 B.n747 10.6151
R1315 B.n747 B.n38 10.6151
R1316 B.n741 B.n38 10.6151
R1317 B.n741 B.n740 10.6151
R1318 B.n740 B.n739 10.6151
R1319 B.n739 B.n45 10.6151
R1320 B.n733 B.n45 10.6151
R1321 B.n733 B.n732 10.6151
R1322 B.n732 B.n731 10.6151
R1323 B.n731 B.n51 10.6151
R1324 B.n725 B.n51 10.6151
R1325 B.n725 B.n724 10.6151
R1326 B.n724 B.n723 10.6151
R1327 B.n723 B.n59 10.6151
R1328 B.n717 B.n59 10.6151
R1329 B.n643 B.n86 9.36635
R1330 B.n619 B.n94 9.36635
R1331 B.n202 B.n198 9.36635
R1332 B.n302 B.n301 9.36635
R1333 B.n485 B.t0 4.09352
R1334 B.t17 B.n775 4.09352
R1335 B.n787 B.n0 2.81026
R1336 B.n787 B.n1 2.81026
R1337 B.n639 B.n86 1.24928
R1338 B.n623 B.n94 1.24928
R1339 B.n320 B.n202 1.24928
R1340 B.n303 B.n302 1.24928
R1341 VP.n14 VP.n0 161.3
R1342 VP.n13 VP.n12 161.3
R1343 VP.n11 VP.n1 161.3
R1344 VP.n10 VP.n9 161.3
R1345 VP.n8 VP.n2 161.3
R1346 VP.n7 VP.n6 161.3
R1347 VP.n4 VP.t2 136.763
R1348 VP.n4 VP.t0 135.988
R1349 VP.n3 VP.t3 100.572
R1350 VP.n15 VP.t1 100.572
R1351 VP.n5 VP.n3 100.236
R1352 VP.n16 VP.n15 100.236
R1353 VP.n9 VP.n1 56.5193
R1354 VP.n5 VP.n4 49.7913
R1355 VP.n8 VP.n7 24.4675
R1356 VP.n9 VP.n8 24.4675
R1357 VP.n13 VP.n1 24.4675
R1358 VP.n14 VP.n13 24.4675
R1359 VP.n7 VP.n3 10.5213
R1360 VP.n15 VP.n14 10.5213
R1361 VP.n6 VP.n5 0.278367
R1362 VP.n16 VP.n0 0.278367
R1363 VP.n6 VP.n2 0.189894
R1364 VP.n10 VP.n2 0.189894
R1365 VP.n11 VP.n10 0.189894
R1366 VP.n12 VP.n11 0.189894
R1367 VP.n12 VP.n0 0.189894
R1368 VP VP.n16 0.153454
R1369 VTAIL.n458 VTAIL.n406 289.615
R1370 VTAIL.n52 VTAIL.n0 289.615
R1371 VTAIL.n110 VTAIL.n58 289.615
R1372 VTAIL.n168 VTAIL.n116 289.615
R1373 VTAIL.n400 VTAIL.n348 289.615
R1374 VTAIL.n342 VTAIL.n290 289.615
R1375 VTAIL.n284 VTAIL.n232 289.615
R1376 VTAIL.n226 VTAIL.n174 289.615
R1377 VTAIL.n425 VTAIL.n424 185
R1378 VTAIL.n422 VTAIL.n421 185
R1379 VTAIL.n431 VTAIL.n430 185
R1380 VTAIL.n433 VTAIL.n432 185
R1381 VTAIL.n418 VTAIL.n417 185
R1382 VTAIL.n439 VTAIL.n438 185
R1383 VTAIL.n442 VTAIL.n441 185
R1384 VTAIL.n440 VTAIL.n414 185
R1385 VTAIL.n447 VTAIL.n413 185
R1386 VTAIL.n449 VTAIL.n448 185
R1387 VTAIL.n451 VTAIL.n450 185
R1388 VTAIL.n410 VTAIL.n409 185
R1389 VTAIL.n457 VTAIL.n456 185
R1390 VTAIL.n459 VTAIL.n458 185
R1391 VTAIL.n19 VTAIL.n18 185
R1392 VTAIL.n16 VTAIL.n15 185
R1393 VTAIL.n25 VTAIL.n24 185
R1394 VTAIL.n27 VTAIL.n26 185
R1395 VTAIL.n12 VTAIL.n11 185
R1396 VTAIL.n33 VTAIL.n32 185
R1397 VTAIL.n36 VTAIL.n35 185
R1398 VTAIL.n34 VTAIL.n8 185
R1399 VTAIL.n41 VTAIL.n7 185
R1400 VTAIL.n43 VTAIL.n42 185
R1401 VTAIL.n45 VTAIL.n44 185
R1402 VTAIL.n4 VTAIL.n3 185
R1403 VTAIL.n51 VTAIL.n50 185
R1404 VTAIL.n53 VTAIL.n52 185
R1405 VTAIL.n77 VTAIL.n76 185
R1406 VTAIL.n74 VTAIL.n73 185
R1407 VTAIL.n83 VTAIL.n82 185
R1408 VTAIL.n85 VTAIL.n84 185
R1409 VTAIL.n70 VTAIL.n69 185
R1410 VTAIL.n91 VTAIL.n90 185
R1411 VTAIL.n94 VTAIL.n93 185
R1412 VTAIL.n92 VTAIL.n66 185
R1413 VTAIL.n99 VTAIL.n65 185
R1414 VTAIL.n101 VTAIL.n100 185
R1415 VTAIL.n103 VTAIL.n102 185
R1416 VTAIL.n62 VTAIL.n61 185
R1417 VTAIL.n109 VTAIL.n108 185
R1418 VTAIL.n111 VTAIL.n110 185
R1419 VTAIL.n135 VTAIL.n134 185
R1420 VTAIL.n132 VTAIL.n131 185
R1421 VTAIL.n141 VTAIL.n140 185
R1422 VTAIL.n143 VTAIL.n142 185
R1423 VTAIL.n128 VTAIL.n127 185
R1424 VTAIL.n149 VTAIL.n148 185
R1425 VTAIL.n152 VTAIL.n151 185
R1426 VTAIL.n150 VTAIL.n124 185
R1427 VTAIL.n157 VTAIL.n123 185
R1428 VTAIL.n159 VTAIL.n158 185
R1429 VTAIL.n161 VTAIL.n160 185
R1430 VTAIL.n120 VTAIL.n119 185
R1431 VTAIL.n167 VTAIL.n166 185
R1432 VTAIL.n169 VTAIL.n168 185
R1433 VTAIL.n401 VTAIL.n400 185
R1434 VTAIL.n399 VTAIL.n398 185
R1435 VTAIL.n352 VTAIL.n351 185
R1436 VTAIL.n393 VTAIL.n392 185
R1437 VTAIL.n391 VTAIL.n390 185
R1438 VTAIL.n389 VTAIL.n355 185
R1439 VTAIL.n359 VTAIL.n356 185
R1440 VTAIL.n384 VTAIL.n383 185
R1441 VTAIL.n382 VTAIL.n381 185
R1442 VTAIL.n361 VTAIL.n360 185
R1443 VTAIL.n376 VTAIL.n375 185
R1444 VTAIL.n374 VTAIL.n373 185
R1445 VTAIL.n365 VTAIL.n364 185
R1446 VTAIL.n368 VTAIL.n367 185
R1447 VTAIL.n343 VTAIL.n342 185
R1448 VTAIL.n341 VTAIL.n340 185
R1449 VTAIL.n294 VTAIL.n293 185
R1450 VTAIL.n335 VTAIL.n334 185
R1451 VTAIL.n333 VTAIL.n332 185
R1452 VTAIL.n331 VTAIL.n297 185
R1453 VTAIL.n301 VTAIL.n298 185
R1454 VTAIL.n326 VTAIL.n325 185
R1455 VTAIL.n324 VTAIL.n323 185
R1456 VTAIL.n303 VTAIL.n302 185
R1457 VTAIL.n318 VTAIL.n317 185
R1458 VTAIL.n316 VTAIL.n315 185
R1459 VTAIL.n307 VTAIL.n306 185
R1460 VTAIL.n310 VTAIL.n309 185
R1461 VTAIL.n285 VTAIL.n284 185
R1462 VTAIL.n283 VTAIL.n282 185
R1463 VTAIL.n236 VTAIL.n235 185
R1464 VTAIL.n277 VTAIL.n276 185
R1465 VTAIL.n275 VTAIL.n274 185
R1466 VTAIL.n273 VTAIL.n239 185
R1467 VTAIL.n243 VTAIL.n240 185
R1468 VTAIL.n268 VTAIL.n267 185
R1469 VTAIL.n266 VTAIL.n265 185
R1470 VTAIL.n245 VTAIL.n244 185
R1471 VTAIL.n260 VTAIL.n259 185
R1472 VTAIL.n258 VTAIL.n257 185
R1473 VTAIL.n249 VTAIL.n248 185
R1474 VTAIL.n252 VTAIL.n251 185
R1475 VTAIL.n227 VTAIL.n226 185
R1476 VTAIL.n225 VTAIL.n224 185
R1477 VTAIL.n178 VTAIL.n177 185
R1478 VTAIL.n219 VTAIL.n218 185
R1479 VTAIL.n217 VTAIL.n216 185
R1480 VTAIL.n215 VTAIL.n181 185
R1481 VTAIL.n185 VTAIL.n182 185
R1482 VTAIL.n210 VTAIL.n209 185
R1483 VTAIL.n208 VTAIL.n207 185
R1484 VTAIL.n187 VTAIL.n186 185
R1485 VTAIL.n202 VTAIL.n201 185
R1486 VTAIL.n200 VTAIL.n199 185
R1487 VTAIL.n191 VTAIL.n190 185
R1488 VTAIL.n194 VTAIL.n193 185
R1489 VTAIL.t6 VTAIL.n423 149.524
R1490 VTAIL.t7 VTAIL.n17 149.524
R1491 VTAIL.t2 VTAIL.n75 149.524
R1492 VTAIL.t3 VTAIL.n133 149.524
R1493 VTAIL.t1 VTAIL.n366 149.524
R1494 VTAIL.t4 VTAIL.n308 149.524
R1495 VTAIL.t5 VTAIL.n250 149.524
R1496 VTAIL.t0 VTAIL.n192 149.524
R1497 VTAIL.n424 VTAIL.n421 104.615
R1498 VTAIL.n431 VTAIL.n421 104.615
R1499 VTAIL.n432 VTAIL.n431 104.615
R1500 VTAIL.n432 VTAIL.n417 104.615
R1501 VTAIL.n439 VTAIL.n417 104.615
R1502 VTAIL.n441 VTAIL.n439 104.615
R1503 VTAIL.n441 VTAIL.n440 104.615
R1504 VTAIL.n440 VTAIL.n413 104.615
R1505 VTAIL.n449 VTAIL.n413 104.615
R1506 VTAIL.n450 VTAIL.n449 104.615
R1507 VTAIL.n450 VTAIL.n409 104.615
R1508 VTAIL.n457 VTAIL.n409 104.615
R1509 VTAIL.n458 VTAIL.n457 104.615
R1510 VTAIL.n18 VTAIL.n15 104.615
R1511 VTAIL.n25 VTAIL.n15 104.615
R1512 VTAIL.n26 VTAIL.n25 104.615
R1513 VTAIL.n26 VTAIL.n11 104.615
R1514 VTAIL.n33 VTAIL.n11 104.615
R1515 VTAIL.n35 VTAIL.n33 104.615
R1516 VTAIL.n35 VTAIL.n34 104.615
R1517 VTAIL.n34 VTAIL.n7 104.615
R1518 VTAIL.n43 VTAIL.n7 104.615
R1519 VTAIL.n44 VTAIL.n43 104.615
R1520 VTAIL.n44 VTAIL.n3 104.615
R1521 VTAIL.n51 VTAIL.n3 104.615
R1522 VTAIL.n52 VTAIL.n51 104.615
R1523 VTAIL.n76 VTAIL.n73 104.615
R1524 VTAIL.n83 VTAIL.n73 104.615
R1525 VTAIL.n84 VTAIL.n83 104.615
R1526 VTAIL.n84 VTAIL.n69 104.615
R1527 VTAIL.n91 VTAIL.n69 104.615
R1528 VTAIL.n93 VTAIL.n91 104.615
R1529 VTAIL.n93 VTAIL.n92 104.615
R1530 VTAIL.n92 VTAIL.n65 104.615
R1531 VTAIL.n101 VTAIL.n65 104.615
R1532 VTAIL.n102 VTAIL.n101 104.615
R1533 VTAIL.n102 VTAIL.n61 104.615
R1534 VTAIL.n109 VTAIL.n61 104.615
R1535 VTAIL.n110 VTAIL.n109 104.615
R1536 VTAIL.n134 VTAIL.n131 104.615
R1537 VTAIL.n141 VTAIL.n131 104.615
R1538 VTAIL.n142 VTAIL.n141 104.615
R1539 VTAIL.n142 VTAIL.n127 104.615
R1540 VTAIL.n149 VTAIL.n127 104.615
R1541 VTAIL.n151 VTAIL.n149 104.615
R1542 VTAIL.n151 VTAIL.n150 104.615
R1543 VTAIL.n150 VTAIL.n123 104.615
R1544 VTAIL.n159 VTAIL.n123 104.615
R1545 VTAIL.n160 VTAIL.n159 104.615
R1546 VTAIL.n160 VTAIL.n119 104.615
R1547 VTAIL.n167 VTAIL.n119 104.615
R1548 VTAIL.n168 VTAIL.n167 104.615
R1549 VTAIL.n400 VTAIL.n399 104.615
R1550 VTAIL.n399 VTAIL.n351 104.615
R1551 VTAIL.n392 VTAIL.n351 104.615
R1552 VTAIL.n392 VTAIL.n391 104.615
R1553 VTAIL.n391 VTAIL.n355 104.615
R1554 VTAIL.n359 VTAIL.n355 104.615
R1555 VTAIL.n383 VTAIL.n359 104.615
R1556 VTAIL.n383 VTAIL.n382 104.615
R1557 VTAIL.n382 VTAIL.n360 104.615
R1558 VTAIL.n375 VTAIL.n360 104.615
R1559 VTAIL.n375 VTAIL.n374 104.615
R1560 VTAIL.n374 VTAIL.n364 104.615
R1561 VTAIL.n367 VTAIL.n364 104.615
R1562 VTAIL.n342 VTAIL.n341 104.615
R1563 VTAIL.n341 VTAIL.n293 104.615
R1564 VTAIL.n334 VTAIL.n293 104.615
R1565 VTAIL.n334 VTAIL.n333 104.615
R1566 VTAIL.n333 VTAIL.n297 104.615
R1567 VTAIL.n301 VTAIL.n297 104.615
R1568 VTAIL.n325 VTAIL.n301 104.615
R1569 VTAIL.n325 VTAIL.n324 104.615
R1570 VTAIL.n324 VTAIL.n302 104.615
R1571 VTAIL.n317 VTAIL.n302 104.615
R1572 VTAIL.n317 VTAIL.n316 104.615
R1573 VTAIL.n316 VTAIL.n306 104.615
R1574 VTAIL.n309 VTAIL.n306 104.615
R1575 VTAIL.n284 VTAIL.n283 104.615
R1576 VTAIL.n283 VTAIL.n235 104.615
R1577 VTAIL.n276 VTAIL.n235 104.615
R1578 VTAIL.n276 VTAIL.n275 104.615
R1579 VTAIL.n275 VTAIL.n239 104.615
R1580 VTAIL.n243 VTAIL.n239 104.615
R1581 VTAIL.n267 VTAIL.n243 104.615
R1582 VTAIL.n267 VTAIL.n266 104.615
R1583 VTAIL.n266 VTAIL.n244 104.615
R1584 VTAIL.n259 VTAIL.n244 104.615
R1585 VTAIL.n259 VTAIL.n258 104.615
R1586 VTAIL.n258 VTAIL.n248 104.615
R1587 VTAIL.n251 VTAIL.n248 104.615
R1588 VTAIL.n226 VTAIL.n225 104.615
R1589 VTAIL.n225 VTAIL.n177 104.615
R1590 VTAIL.n218 VTAIL.n177 104.615
R1591 VTAIL.n218 VTAIL.n217 104.615
R1592 VTAIL.n217 VTAIL.n181 104.615
R1593 VTAIL.n185 VTAIL.n181 104.615
R1594 VTAIL.n209 VTAIL.n185 104.615
R1595 VTAIL.n209 VTAIL.n208 104.615
R1596 VTAIL.n208 VTAIL.n186 104.615
R1597 VTAIL.n201 VTAIL.n186 104.615
R1598 VTAIL.n201 VTAIL.n200 104.615
R1599 VTAIL.n200 VTAIL.n190 104.615
R1600 VTAIL.n193 VTAIL.n190 104.615
R1601 VTAIL.n424 VTAIL.t6 52.3082
R1602 VTAIL.n18 VTAIL.t7 52.3082
R1603 VTAIL.n76 VTAIL.t2 52.3082
R1604 VTAIL.n134 VTAIL.t3 52.3082
R1605 VTAIL.n367 VTAIL.t1 52.3082
R1606 VTAIL.n309 VTAIL.t4 52.3082
R1607 VTAIL.n251 VTAIL.t5 52.3082
R1608 VTAIL.n193 VTAIL.t0 52.3082
R1609 VTAIL.n463 VTAIL.n462 35.4823
R1610 VTAIL.n57 VTAIL.n56 35.4823
R1611 VTAIL.n115 VTAIL.n114 35.4823
R1612 VTAIL.n173 VTAIL.n172 35.4823
R1613 VTAIL.n405 VTAIL.n404 35.4823
R1614 VTAIL.n347 VTAIL.n346 35.4823
R1615 VTAIL.n289 VTAIL.n288 35.4823
R1616 VTAIL.n231 VTAIL.n230 35.4823
R1617 VTAIL.n463 VTAIL.n405 24.2462
R1618 VTAIL.n231 VTAIL.n173 24.2462
R1619 VTAIL.n448 VTAIL.n447 13.1884
R1620 VTAIL.n42 VTAIL.n41 13.1884
R1621 VTAIL.n100 VTAIL.n99 13.1884
R1622 VTAIL.n158 VTAIL.n157 13.1884
R1623 VTAIL.n390 VTAIL.n389 13.1884
R1624 VTAIL.n332 VTAIL.n331 13.1884
R1625 VTAIL.n274 VTAIL.n273 13.1884
R1626 VTAIL.n216 VTAIL.n215 13.1884
R1627 VTAIL.n446 VTAIL.n414 12.8005
R1628 VTAIL.n451 VTAIL.n412 12.8005
R1629 VTAIL.n40 VTAIL.n8 12.8005
R1630 VTAIL.n45 VTAIL.n6 12.8005
R1631 VTAIL.n98 VTAIL.n66 12.8005
R1632 VTAIL.n103 VTAIL.n64 12.8005
R1633 VTAIL.n156 VTAIL.n124 12.8005
R1634 VTAIL.n161 VTAIL.n122 12.8005
R1635 VTAIL.n393 VTAIL.n354 12.8005
R1636 VTAIL.n388 VTAIL.n356 12.8005
R1637 VTAIL.n335 VTAIL.n296 12.8005
R1638 VTAIL.n330 VTAIL.n298 12.8005
R1639 VTAIL.n277 VTAIL.n238 12.8005
R1640 VTAIL.n272 VTAIL.n240 12.8005
R1641 VTAIL.n219 VTAIL.n180 12.8005
R1642 VTAIL.n214 VTAIL.n182 12.8005
R1643 VTAIL.n443 VTAIL.n442 12.0247
R1644 VTAIL.n452 VTAIL.n410 12.0247
R1645 VTAIL.n37 VTAIL.n36 12.0247
R1646 VTAIL.n46 VTAIL.n4 12.0247
R1647 VTAIL.n95 VTAIL.n94 12.0247
R1648 VTAIL.n104 VTAIL.n62 12.0247
R1649 VTAIL.n153 VTAIL.n152 12.0247
R1650 VTAIL.n162 VTAIL.n120 12.0247
R1651 VTAIL.n394 VTAIL.n352 12.0247
R1652 VTAIL.n385 VTAIL.n384 12.0247
R1653 VTAIL.n336 VTAIL.n294 12.0247
R1654 VTAIL.n327 VTAIL.n326 12.0247
R1655 VTAIL.n278 VTAIL.n236 12.0247
R1656 VTAIL.n269 VTAIL.n268 12.0247
R1657 VTAIL.n220 VTAIL.n178 12.0247
R1658 VTAIL.n211 VTAIL.n210 12.0247
R1659 VTAIL.n438 VTAIL.n416 11.249
R1660 VTAIL.n456 VTAIL.n455 11.249
R1661 VTAIL.n32 VTAIL.n10 11.249
R1662 VTAIL.n50 VTAIL.n49 11.249
R1663 VTAIL.n90 VTAIL.n68 11.249
R1664 VTAIL.n108 VTAIL.n107 11.249
R1665 VTAIL.n148 VTAIL.n126 11.249
R1666 VTAIL.n166 VTAIL.n165 11.249
R1667 VTAIL.n398 VTAIL.n397 11.249
R1668 VTAIL.n381 VTAIL.n358 11.249
R1669 VTAIL.n340 VTAIL.n339 11.249
R1670 VTAIL.n323 VTAIL.n300 11.249
R1671 VTAIL.n282 VTAIL.n281 11.249
R1672 VTAIL.n265 VTAIL.n242 11.249
R1673 VTAIL.n224 VTAIL.n223 11.249
R1674 VTAIL.n207 VTAIL.n184 11.249
R1675 VTAIL.n437 VTAIL.n418 10.4732
R1676 VTAIL.n459 VTAIL.n408 10.4732
R1677 VTAIL.n31 VTAIL.n12 10.4732
R1678 VTAIL.n53 VTAIL.n2 10.4732
R1679 VTAIL.n89 VTAIL.n70 10.4732
R1680 VTAIL.n111 VTAIL.n60 10.4732
R1681 VTAIL.n147 VTAIL.n128 10.4732
R1682 VTAIL.n169 VTAIL.n118 10.4732
R1683 VTAIL.n401 VTAIL.n350 10.4732
R1684 VTAIL.n380 VTAIL.n361 10.4732
R1685 VTAIL.n343 VTAIL.n292 10.4732
R1686 VTAIL.n322 VTAIL.n303 10.4732
R1687 VTAIL.n285 VTAIL.n234 10.4732
R1688 VTAIL.n264 VTAIL.n245 10.4732
R1689 VTAIL.n227 VTAIL.n176 10.4732
R1690 VTAIL.n206 VTAIL.n187 10.4732
R1691 VTAIL.n425 VTAIL.n423 10.2747
R1692 VTAIL.n19 VTAIL.n17 10.2747
R1693 VTAIL.n77 VTAIL.n75 10.2747
R1694 VTAIL.n135 VTAIL.n133 10.2747
R1695 VTAIL.n368 VTAIL.n366 10.2747
R1696 VTAIL.n310 VTAIL.n308 10.2747
R1697 VTAIL.n252 VTAIL.n250 10.2747
R1698 VTAIL.n194 VTAIL.n192 10.2747
R1699 VTAIL.n434 VTAIL.n433 9.69747
R1700 VTAIL.n460 VTAIL.n406 9.69747
R1701 VTAIL.n28 VTAIL.n27 9.69747
R1702 VTAIL.n54 VTAIL.n0 9.69747
R1703 VTAIL.n86 VTAIL.n85 9.69747
R1704 VTAIL.n112 VTAIL.n58 9.69747
R1705 VTAIL.n144 VTAIL.n143 9.69747
R1706 VTAIL.n170 VTAIL.n116 9.69747
R1707 VTAIL.n402 VTAIL.n348 9.69747
R1708 VTAIL.n377 VTAIL.n376 9.69747
R1709 VTAIL.n344 VTAIL.n290 9.69747
R1710 VTAIL.n319 VTAIL.n318 9.69747
R1711 VTAIL.n286 VTAIL.n232 9.69747
R1712 VTAIL.n261 VTAIL.n260 9.69747
R1713 VTAIL.n228 VTAIL.n174 9.69747
R1714 VTAIL.n203 VTAIL.n202 9.69747
R1715 VTAIL.n462 VTAIL.n461 9.45567
R1716 VTAIL.n56 VTAIL.n55 9.45567
R1717 VTAIL.n114 VTAIL.n113 9.45567
R1718 VTAIL.n172 VTAIL.n171 9.45567
R1719 VTAIL.n404 VTAIL.n403 9.45567
R1720 VTAIL.n346 VTAIL.n345 9.45567
R1721 VTAIL.n288 VTAIL.n287 9.45567
R1722 VTAIL.n230 VTAIL.n229 9.45567
R1723 VTAIL.n461 VTAIL.n460 9.3005
R1724 VTAIL.n408 VTAIL.n407 9.3005
R1725 VTAIL.n455 VTAIL.n454 9.3005
R1726 VTAIL.n453 VTAIL.n452 9.3005
R1727 VTAIL.n412 VTAIL.n411 9.3005
R1728 VTAIL.n427 VTAIL.n426 9.3005
R1729 VTAIL.n429 VTAIL.n428 9.3005
R1730 VTAIL.n420 VTAIL.n419 9.3005
R1731 VTAIL.n435 VTAIL.n434 9.3005
R1732 VTAIL.n437 VTAIL.n436 9.3005
R1733 VTAIL.n416 VTAIL.n415 9.3005
R1734 VTAIL.n444 VTAIL.n443 9.3005
R1735 VTAIL.n446 VTAIL.n445 9.3005
R1736 VTAIL.n55 VTAIL.n54 9.3005
R1737 VTAIL.n2 VTAIL.n1 9.3005
R1738 VTAIL.n49 VTAIL.n48 9.3005
R1739 VTAIL.n47 VTAIL.n46 9.3005
R1740 VTAIL.n6 VTAIL.n5 9.3005
R1741 VTAIL.n21 VTAIL.n20 9.3005
R1742 VTAIL.n23 VTAIL.n22 9.3005
R1743 VTAIL.n14 VTAIL.n13 9.3005
R1744 VTAIL.n29 VTAIL.n28 9.3005
R1745 VTAIL.n31 VTAIL.n30 9.3005
R1746 VTAIL.n10 VTAIL.n9 9.3005
R1747 VTAIL.n38 VTAIL.n37 9.3005
R1748 VTAIL.n40 VTAIL.n39 9.3005
R1749 VTAIL.n113 VTAIL.n112 9.3005
R1750 VTAIL.n60 VTAIL.n59 9.3005
R1751 VTAIL.n107 VTAIL.n106 9.3005
R1752 VTAIL.n105 VTAIL.n104 9.3005
R1753 VTAIL.n64 VTAIL.n63 9.3005
R1754 VTAIL.n79 VTAIL.n78 9.3005
R1755 VTAIL.n81 VTAIL.n80 9.3005
R1756 VTAIL.n72 VTAIL.n71 9.3005
R1757 VTAIL.n87 VTAIL.n86 9.3005
R1758 VTAIL.n89 VTAIL.n88 9.3005
R1759 VTAIL.n68 VTAIL.n67 9.3005
R1760 VTAIL.n96 VTAIL.n95 9.3005
R1761 VTAIL.n98 VTAIL.n97 9.3005
R1762 VTAIL.n171 VTAIL.n170 9.3005
R1763 VTAIL.n118 VTAIL.n117 9.3005
R1764 VTAIL.n165 VTAIL.n164 9.3005
R1765 VTAIL.n163 VTAIL.n162 9.3005
R1766 VTAIL.n122 VTAIL.n121 9.3005
R1767 VTAIL.n137 VTAIL.n136 9.3005
R1768 VTAIL.n139 VTAIL.n138 9.3005
R1769 VTAIL.n130 VTAIL.n129 9.3005
R1770 VTAIL.n145 VTAIL.n144 9.3005
R1771 VTAIL.n147 VTAIL.n146 9.3005
R1772 VTAIL.n126 VTAIL.n125 9.3005
R1773 VTAIL.n154 VTAIL.n153 9.3005
R1774 VTAIL.n156 VTAIL.n155 9.3005
R1775 VTAIL.n370 VTAIL.n369 9.3005
R1776 VTAIL.n372 VTAIL.n371 9.3005
R1777 VTAIL.n363 VTAIL.n362 9.3005
R1778 VTAIL.n378 VTAIL.n377 9.3005
R1779 VTAIL.n380 VTAIL.n379 9.3005
R1780 VTAIL.n358 VTAIL.n357 9.3005
R1781 VTAIL.n386 VTAIL.n385 9.3005
R1782 VTAIL.n388 VTAIL.n387 9.3005
R1783 VTAIL.n403 VTAIL.n402 9.3005
R1784 VTAIL.n350 VTAIL.n349 9.3005
R1785 VTAIL.n397 VTAIL.n396 9.3005
R1786 VTAIL.n395 VTAIL.n394 9.3005
R1787 VTAIL.n354 VTAIL.n353 9.3005
R1788 VTAIL.n312 VTAIL.n311 9.3005
R1789 VTAIL.n314 VTAIL.n313 9.3005
R1790 VTAIL.n305 VTAIL.n304 9.3005
R1791 VTAIL.n320 VTAIL.n319 9.3005
R1792 VTAIL.n322 VTAIL.n321 9.3005
R1793 VTAIL.n300 VTAIL.n299 9.3005
R1794 VTAIL.n328 VTAIL.n327 9.3005
R1795 VTAIL.n330 VTAIL.n329 9.3005
R1796 VTAIL.n345 VTAIL.n344 9.3005
R1797 VTAIL.n292 VTAIL.n291 9.3005
R1798 VTAIL.n339 VTAIL.n338 9.3005
R1799 VTAIL.n337 VTAIL.n336 9.3005
R1800 VTAIL.n296 VTAIL.n295 9.3005
R1801 VTAIL.n254 VTAIL.n253 9.3005
R1802 VTAIL.n256 VTAIL.n255 9.3005
R1803 VTAIL.n247 VTAIL.n246 9.3005
R1804 VTAIL.n262 VTAIL.n261 9.3005
R1805 VTAIL.n264 VTAIL.n263 9.3005
R1806 VTAIL.n242 VTAIL.n241 9.3005
R1807 VTAIL.n270 VTAIL.n269 9.3005
R1808 VTAIL.n272 VTAIL.n271 9.3005
R1809 VTAIL.n287 VTAIL.n286 9.3005
R1810 VTAIL.n234 VTAIL.n233 9.3005
R1811 VTAIL.n281 VTAIL.n280 9.3005
R1812 VTAIL.n279 VTAIL.n278 9.3005
R1813 VTAIL.n238 VTAIL.n237 9.3005
R1814 VTAIL.n196 VTAIL.n195 9.3005
R1815 VTAIL.n198 VTAIL.n197 9.3005
R1816 VTAIL.n189 VTAIL.n188 9.3005
R1817 VTAIL.n204 VTAIL.n203 9.3005
R1818 VTAIL.n206 VTAIL.n205 9.3005
R1819 VTAIL.n184 VTAIL.n183 9.3005
R1820 VTAIL.n212 VTAIL.n211 9.3005
R1821 VTAIL.n214 VTAIL.n213 9.3005
R1822 VTAIL.n229 VTAIL.n228 9.3005
R1823 VTAIL.n176 VTAIL.n175 9.3005
R1824 VTAIL.n223 VTAIL.n222 9.3005
R1825 VTAIL.n221 VTAIL.n220 9.3005
R1826 VTAIL.n180 VTAIL.n179 9.3005
R1827 VTAIL.n430 VTAIL.n420 8.92171
R1828 VTAIL.n24 VTAIL.n14 8.92171
R1829 VTAIL.n82 VTAIL.n72 8.92171
R1830 VTAIL.n140 VTAIL.n130 8.92171
R1831 VTAIL.n373 VTAIL.n363 8.92171
R1832 VTAIL.n315 VTAIL.n305 8.92171
R1833 VTAIL.n257 VTAIL.n247 8.92171
R1834 VTAIL.n199 VTAIL.n189 8.92171
R1835 VTAIL.n429 VTAIL.n422 8.14595
R1836 VTAIL.n23 VTAIL.n16 8.14595
R1837 VTAIL.n81 VTAIL.n74 8.14595
R1838 VTAIL.n139 VTAIL.n132 8.14595
R1839 VTAIL.n372 VTAIL.n365 8.14595
R1840 VTAIL.n314 VTAIL.n307 8.14595
R1841 VTAIL.n256 VTAIL.n249 8.14595
R1842 VTAIL.n198 VTAIL.n191 8.14595
R1843 VTAIL.n426 VTAIL.n425 7.3702
R1844 VTAIL.n20 VTAIL.n19 7.3702
R1845 VTAIL.n78 VTAIL.n77 7.3702
R1846 VTAIL.n136 VTAIL.n135 7.3702
R1847 VTAIL.n369 VTAIL.n368 7.3702
R1848 VTAIL.n311 VTAIL.n310 7.3702
R1849 VTAIL.n253 VTAIL.n252 7.3702
R1850 VTAIL.n195 VTAIL.n194 7.3702
R1851 VTAIL.n426 VTAIL.n422 5.81868
R1852 VTAIL.n20 VTAIL.n16 5.81868
R1853 VTAIL.n78 VTAIL.n74 5.81868
R1854 VTAIL.n136 VTAIL.n132 5.81868
R1855 VTAIL.n369 VTAIL.n365 5.81868
R1856 VTAIL.n311 VTAIL.n307 5.81868
R1857 VTAIL.n253 VTAIL.n249 5.81868
R1858 VTAIL.n195 VTAIL.n191 5.81868
R1859 VTAIL.n430 VTAIL.n429 5.04292
R1860 VTAIL.n24 VTAIL.n23 5.04292
R1861 VTAIL.n82 VTAIL.n81 5.04292
R1862 VTAIL.n140 VTAIL.n139 5.04292
R1863 VTAIL.n373 VTAIL.n372 5.04292
R1864 VTAIL.n315 VTAIL.n314 5.04292
R1865 VTAIL.n257 VTAIL.n256 5.04292
R1866 VTAIL.n199 VTAIL.n198 5.04292
R1867 VTAIL.n433 VTAIL.n420 4.26717
R1868 VTAIL.n462 VTAIL.n406 4.26717
R1869 VTAIL.n27 VTAIL.n14 4.26717
R1870 VTAIL.n56 VTAIL.n0 4.26717
R1871 VTAIL.n85 VTAIL.n72 4.26717
R1872 VTAIL.n114 VTAIL.n58 4.26717
R1873 VTAIL.n143 VTAIL.n130 4.26717
R1874 VTAIL.n172 VTAIL.n116 4.26717
R1875 VTAIL.n404 VTAIL.n348 4.26717
R1876 VTAIL.n376 VTAIL.n363 4.26717
R1877 VTAIL.n346 VTAIL.n290 4.26717
R1878 VTAIL.n318 VTAIL.n305 4.26717
R1879 VTAIL.n288 VTAIL.n232 4.26717
R1880 VTAIL.n260 VTAIL.n247 4.26717
R1881 VTAIL.n230 VTAIL.n174 4.26717
R1882 VTAIL.n202 VTAIL.n189 4.26717
R1883 VTAIL.n434 VTAIL.n418 3.49141
R1884 VTAIL.n460 VTAIL.n459 3.49141
R1885 VTAIL.n28 VTAIL.n12 3.49141
R1886 VTAIL.n54 VTAIL.n53 3.49141
R1887 VTAIL.n86 VTAIL.n70 3.49141
R1888 VTAIL.n112 VTAIL.n111 3.49141
R1889 VTAIL.n144 VTAIL.n128 3.49141
R1890 VTAIL.n170 VTAIL.n169 3.49141
R1891 VTAIL.n402 VTAIL.n401 3.49141
R1892 VTAIL.n377 VTAIL.n361 3.49141
R1893 VTAIL.n344 VTAIL.n343 3.49141
R1894 VTAIL.n319 VTAIL.n303 3.49141
R1895 VTAIL.n286 VTAIL.n285 3.49141
R1896 VTAIL.n261 VTAIL.n245 3.49141
R1897 VTAIL.n228 VTAIL.n227 3.49141
R1898 VTAIL.n203 VTAIL.n187 3.49141
R1899 VTAIL.n427 VTAIL.n423 2.84303
R1900 VTAIL.n21 VTAIL.n17 2.84303
R1901 VTAIL.n79 VTAIL.n75 2.84303
R1902 VTAIL.n137 VTAIL.n133 2.84303
R1903 VTAIL.n370 VTAIL.n366 2.84303
R1904 VTAIL.n312 VTAIL.n308 2.84303
R1905 VTAIL.n254 VTAIL.n250 2.84303
R1906 VTAIL.n196 VTAIL.n192 2.84303
R1907 VTAIL.n438 VTAIL.n437 2.71565
R1908 VTAIL.n456 VTAIL.n408 2.71565
R1909 VTAIL.n32 VTAIL.n31 2.71565
R1910 VTAIL.n50 VTAIL.n2 2.71565
R1911 VTAIL.n90 VTAIL.n89 2.71565
R1912 VTAIL.n108 VTAIL.n60 2.71565
R1913 VTAIL.n148 VTAIL.n147 2.71565
R1914 VTAIL.n166 VTAIL.n118 2.71565
R1915 VTAIL.n398 VTAIL.n350 2.71565
R1916 VTAIL.n381 VTAIL.n380 2.71565
R1917 VTAIL.n340 VTAIL.n292 2.71565
R1918 VTAIL.n323 VTAIL.n322 2.71565
R1919 VTAIL.n282 VTAIL.n234 2.71565
R1920 VTAIL.n265 VTAIL.n264 2.71565
R1921 VTAIL.n224 VTAIL.n176 2.71565
R1922 VTAIL.n207 VTAIL.n206 2.71565
R1923 VTAIL.n289 VTAIL.n231 2.52636
R1924 VTAIL.n405 VTAIL.n347 2.52636
R1925 VTAIL.n173 VTAIL.n115 2.52636
R1926 VTAIL.n442 VTAIL.n416 1.93989
R1927 VTAIL.n455 VTAIL.n410 1.93989
R1928 VTAIL.n36 VTAIL.n10 1.93989
R1929 VTAIL.n49 VTAIL.n4 1.93989
R1930 VTAIL.n94 VTAIL.n68 1.93989
R1931 VTAIL.n107 VTAIL.n62 1.93989
R1932 VTAIL.n152 VTAIL.n126 1.93989
R1933 VTAIL.n165 VTAIL.n120 1.93989
R1934 VTAIL.n397 VTAIL.n352 1.93989
R1935 VTAIL.n384 VTAIL.n358 1.93989
R1936 VTAIL.n339 VTAIL.n294 1.93989
R1937 VTAIL.n326 VTAIL.n300 1.93989
R1938 VTAIL.n281 VTAIL.n236 1.93989
R1939 VTAIL.n268 VTAIL.n242 1.93989
R1940 VTAIL.n223 VTAIL.n178 1.93989
R1941 VTAIL.n210 VTAIL.n184 1.93989
R1942 VTAIL VTAIL.n57 1.32162
R1943 VTAIL VTAIL.n463 1.20524
R1944 VTAIL.n443 VTAIL.n414 1.16414
R1945 VTAIL.n452 VTAIL.n451 1.16414
R1946 VTAIL.n37 VTAIL.n8 1.16414
R1947 VTAIL.n46 VTAIL.n45 1.16414
R1948 VTAIL.n95 VTAIL.n66 1.16414
R1949 VTAIL.n104 VTAIL.n103 1.16414
R1950 VTAIL.n153 VTAIL.n124 1.16414
R1951 VTAIL.n162 VTAIL.n161 1.16414
R1952 VTAIL.n394 VTAIL.n393 1.16414
R1953 VTAIL.n385 VTAIL.n356 1.16414
R1954 VTAIL.n336 VTAIL.n335 1.16414
R1955 VTAIL.n327 VTAIL.n298 1.16414
R1956 VTAIL.n278 VTAIL.n277 1.16414
R1957 VTAIL.n269 VTAIL.n240 1.16414
R1958 VTAIL.n220 VTAIL.n219 1.16414
R1959 VTAIL.n211 VTAIL.n182 1.16414
R1960 VTAIL.n347 VTAIL.n289 0.470328
R1961 VTAIL.n115 VTAIL.n57 0.470328
R1962 VTAIL.n447 VTAIL.n446 0.388379
R1963 VTAIL.n448 VTAIL.n412 0.388379
R1964 VTAIL.n41 VTAIL.n40 0.388379
R1965 VTAIL.n42 VTAIL.n6 0.388379
R1966 VTAIL.n99 VTAIL.n98 0.388379
R1967 VTAIL.n100 VTAIL.n64 0.388379
R1968 VTAIL.n157 VTAIL.n156 0.388379
R1969 VTAIL.n158 VTAIL.n122 0.388379
R1970 VTAIL.n390 VTAIL.n354 0.388379
R1971 VTAIL.n389 VTAIL.n388 0.388379
R1972 VTAIL.n332 VTAIL.n296 0.388379
R1973 VTAIL.n331 VTAIL.n330 0.388379
R1974 VTAIL.n274 VTAIL.n238 0.388379
R1975 VTAIL.n273 VTAIL.n272 0.388379
R1976 VTAIL.n216 VTAIL.n180 0.388379
R1977 VTAIL.n215 VTAIL.n214 0.388379
R1978 VTAIL.n428 VTAIL.n427 0.155672
R1979 VTAIL.n428 VTAIL.n419 0.155672
R1980 VTAIL.n435 VTAIL.n419 0.155672
R1981 VTAIL.n436 VTAIL.n435 0.155672
R1982 VTAIL.n436 VTAIL.n415 0.155672
R1983 VTAIL.n444 VTAIL.n415 0.155672
R1984 VTAIL.n445 VTAIL.n444 0.155672
R1985 VTAIL.n445 VTAIL.n411 0.155672
R1986 VTAIL.n453 VTAIL.n411 0.155672
R1987 VTAIL.n454 VTAIL.n453 0.155672
R1988 VTAIL.n454 VTAIL.n407 0.155672
R1989 VTAIL.n461 VTAIL.n407 0.155672
R1990 VTAIL.n22 VTAIL.n21 0.155672
R1991 VTAIL.n22 VTAIL.n13 0.155672
R1992 VTAIL.n29 VTAIL.n13 0.155672
R1993 VTAIL.n30 VTAIL.n29 0.155672
R1994 VTAIL.n30 VTAIL.n9 0.155672
R1995 VTAIL.n38 VTAIL.n9 0.155672
R1996 VTAIL.n39 VTAIL.n38 0.155672
R1997 VTAIL.n39 VTAIL.n5 0.155672
R1998 VTAIL.n47 VTAIL.n5 0.155672
R1999 VTAIL.n48 VTAIL.n47 0.155672
R2000 VTAIL.n48 VTAIL.n1 0.155672
R2001 VTAIL.n55 VTAIL.n1 0.155672
R2002 VTAIL.n80 VTAIL.n79 0.155672
R2003 VTAIL.n80 VTAIL.n71 0.155672
R2004 VTAIL.n87 VTAIL.n71 0.155672
R2005 VTAIL.n88 VTAIL.n87 0.155672
R2006 VTAIL.n88 VTAIL.n67 0.155672
R2007 VTAIL.n96 VTAIL.n67 0.155672
R2008 VTAIL.n97 VTAIL.n96 0.155672
R2009 VTAIL.n97 VTAIL.n63 0.155672
R2010 VTAIL.n105 VTAIL.n63 0.155672
R2011 VTAIL.n106 VTAIL.n105 0.155672
R2012 VTAIL.n106 VTAIL.n59 0.155672
R2013 VTAIL.n113 VTAIL.n59 0.155672
R2014 VTAIL.n138 VTAIL.n137 0.155672
R2015 VTAIL.n138 VTAIL.n129 0.155672
R2016 VTAIL.n145 VTAIL.n129 0.155672
R2017 VTAIL.n146 VTAIL.n145 0.155672
R2018 VTAIL.n146 VTAIL.n125 0.155672
R2019 VTAIL.n154 VTAIL.n125 0.155672
R2020 VTAIL.n155 VTAIL.n154 0.155672
R2021 VTAIL.n155 VTAIL.n121 0.155672
R2022 VTAIL.n163 VTAIL.n121 0.155672
R2023 VTAIL.n164 VTAIL.n163 0.155672
R2024 VTAIL.n164 VTAIL.n117 0.155672
R2025 VTAIL.n171 VTAIL.n117 0.155672
R2026 VTAIL.n403 VTAIL.n349 0.155672
R2027 VTAIL.n396 VTAIL.n349 0.155672
R2028 VTAIL.n396 VTAIL.n395 0.155672
R2029 VTAIL.n395 VTAIL.n353 0.155672
R2030 VTAIL.n387 VTAIL.n353 0.155672
R2031 VTAIL.n387 VTAIL.n386 0.155672
R2032 VTAIL.n386 VTAIL.n357 0.155672
R2033 VTAIL.n379 VTAIL.n357 0.155672
R2034 VTAIL.n379 VTAIL.n378 0.155672
R2035 VTAIL.n378 VTAIL.n362 0.155672
R2036 VTAIL.n371 VTAIL.n362 0.155672
R2037 VTAIL.n371 VTAIL.n370 0.155672
R2038 VTAIL.n345 VTAIL.n291 0.155672
R2039 VTAIL.n338 VTAIL.n291 0.155672
R2040 VTAIL.n338 VTAIL.n337 0.155672
R2041 VTAIL.n337 VTAIL.n295 0.155672
R2042 VTAIL.n329 VTAIL.n295 0.155672
R2043 VTAIL.n329 VTAIL.n328 0.155672
R2044 VTAIL.n328 VTAIL.n299 0.155672
R2045 VTAIL.n321 VTAIL.n299 0.155672
R2046 VTAIL.n321 VTAIL.n320 0.155672
R2047 VTAIL.n320 VTAIL.n304 0.155672
R2048 VTAIL.n313 VTAIL.n304 0.155672
R2049 VTAIL.n313 VTAIL.n312 0.155672
R2050 VTAIL.n287 VTAIL.n233 0.155672
R2051 VTAIL.n280 VTAIL.n233 0.155672
R2052 VTAIL.n280 VTAIL.n279 0.155672
R2053 VTAIL.n279 VTAIL.n237 0.155672
R2054 VTAIL.n271 VTAIL.n237 0.155672
R2055 VTAIL.n271 VTAIL.n270 0.155672
R2056 VTAIL.n270 VTAIL.n241 0.155672
R2057 VTAIL.n263 VTAIL.n241 0.155672
R2058 VTAIL.n263 VTAIL.n262 0.155672
R2059 VTAIL.n262 VTAIL.n246 0.155672
R2060 VTAIL.n255 VTAIL.n246 0.155672
R2061 VTAIL.n255 VTAIL.n254 0.155672
R2062 VTAIL.n229 VTAIL.n175 0.155672
R2063 VTAIL.n222 VTAIL.n175 0.155672
R2064 VTAIL.n222 VTAIL.n221 0.155672
R2065 VTAIL.n221 VTAIL.n179 0.155672
R2066 VTAIL.n213 VTAIL.n179 0.155672
R2067 VTAIL.n213 VTAIL.n212 0.155672
R2068 VTAIL.n212 VTAIL.n183 0.155672
R2069 VTAIL.n205 VTAIL.n183 0.155672
R2070 VTAIL.n205 VTAIL.n204 0.155672
R2071 VTAIL.n204 VTAIL.n188 0.155672
R2072 VTAIL.n197 VTAIL.n188 0.155672
R2073 VTAIL.n197 VTAIL.n196 0.155672
R2074 VDD1 VDD1.n1 106.808
R2075 VDD1 VDD1.n0 65.6953
R2076 VDD1.n0 VDD1.t1 1.82538
R2077 VDD1.n0 VDD1.t3 1.82538
R2078 VDD1.n1 VDD1.t0 1.82538
R2079 VDD1.n1 VDD1.t2 1.82538
R2080 VN.n0 VN.t2 136.763
R2081 VN.n1 VN.t1 136.763
R2082 VN.n0 VN.t3 135.988
R2083 VN.n1 VN.t0 135.988
R2084 VN VN.n1 50.0702
R2085 VN VN.n0 4.33156
R2086 VDD2.n2 VDD2.n0 106.282
R2087 VDD2.n2 VDD2.n1 65.6371
R2088 VDD2.n1 VDD2.t3 1.82538
R2089 VDD2.n1 VDD2.t2 1.82538
R2090 VDD2.n0 VDD2.t1 1.82538
R2091 VDD2.n0 VDD2.t0 1.82538
R2092 VDD2 VDD2.n2 0.0586897
C0 VP VTAIL 4.29903f
C1 VP VDD2 0.394441f
C2 VTAIL VDD1 5.13382f
C3 VDD1 VDD2 1.0204f
C4 VTAIL VDD2 5.18803f
C5 VP VN 5.97629f
C6 VDD1 VN 0.149135f
C7 VTAIL VN 4.28493f
C8 VDD2 VN 4.32171f
C9 VP VDD1 4.56628f
C10 VDD2 B 3.690534f
C11 VDD1 B 7.73228f
C12 VTAIL B 9.38606f
C13 VN B 10.592231f
C14 VP B 8.851472f
C15 VDD2.t1 B 0.230627f
C16 VDD2.t0 B 0.230627f
C17 VDD2.n0 B 2.65552f
C18 VDD2.t3 B 0.230627f
C19 VDD2.t2 B 0.230627f
C20 VDD2.n1 B 2.04505f
C21 VDD2.n2 B 3.65221f
C22 VN.t2 B 2.20701f
C23 VN.t3 B 2.20221f
C24 VN.n0 B 1.39349f
C25 VN.t1 B 2.20701f
C26 VN.t0 B 2.20221f
C27 VN.n1 B 2.75201f
C28 VDD1.t1 B 0.233045f
C29 VDD1.t3 B 0.233045f
C30 VDD1.n0 B 2.06689f
C31 VDD1.t0 B 0.233045f
C32 VDD1.t2 B 0.233045f
C33 VDD1.n1 B 2.70915f
C34 VTAIL.n0 B 0.024572f
C35 VTAIL.n1 B 0.016758f
C36 VTAIL.n2 B 0.009005f
C37 VTAIL.n3 B 0.021284f
C38 VTAIL.n4 B 0.009535f
C39 VTAIL.n5 B 0.016758f
C40 VTAIL.n6 B 0.009005f
C41 VTAIL.n7 B 0.021284f
C42 VTAIL.n8 B 0.009535f
C43 VTAIL.n9 B 0.016758f
C44 VTAIL.n10 B 0.009005f
C45 VTAIL.n11 B 0.021284f
C46 VTAIL.n12 B 0.009535f
C47 VTAIL.n13 B 0.016758f
C48 VTAIL.n14 B 0.009005f
C49 VTAIL.n15 B 0.021284f
C50 VTAIL.n16 B 0.009535f
C51 VTAIL.n17 B 0.113425f
C52 VTAIL.t7 B 0.035845f
C53 VTAIL.n18 B 0.015963f
C54 VTAIL.n19 B 0.015046f
C55 VTAIL.n20 B 0.009005f
C56 VTAIL.n21 B 0.759686f
C57 VTAIL.n22 B 0.016758f
C58 VTAIL.n23 B 0.009005f
C59 VTAIL.n24 B 0.009535f
C60 VTAIL.n25 B 0.021284f
C61 VTAIL.n26 B 0.021284f
C62 VTAIL.n27 B 0.009535f
C63 VTAIL.n28 B 0.009005f
C64 VTAIL.n29 B 0.016758f
C65 VTAIL.n30 B 0.016758f
C66 VTAIL.n31 B 0.009005f
C67 VTAIL.n32 B 0.009535f
C68 VTAIL.n33 B 0.021284f
C69 VTAIL.n34 B 0.021284f
C70 VTAIL.n35 B 0.021284f
C71 VTAIL.n36 B 0.009535f
C72 VTAIL.n37 B 0.009005f
C73 VTAIL.n38 B 0.016758f
C74 VTAIL.n39 B 0.016758f
C75 VTAIL.n40 B 0.009005f
C76 VTAIL.n41 B 0.00927f
C77 VTAIL.n42 B 0.00927f
C78 VTAIL.n43 B 0.021284f
C79 VTAIL.n44 B 0.021284f
C80 VTAIL.n45 B 0.009535f
C81 VTAIL.n46 B 0.009005f
C82 VTAIL.n47 B 0.016758f
C83 VTAIL.n48 B 0.016758f
C84 VTAIL.n49 B 0.009005f
C85 VTAIL.n50 B 0.009535f
C86 VTAIL.n51 B 0.021284f
C87 VTAIL.n52 B 0.047877f
C88 VTAIL.n53 B 0.009535f
C89 VTAIL.n54 B 0.009005f
C90 VTAIL.n55 B 0.042627f
C91 VTAIL.n56 B 0.027088f
C92 VTAIL.n57 B 0.113221f
C93 VTAIL.n58 B 0.024572f
C94 VTAIL.n59 B 0.016758f
C95 VTAIL.n60 B 0.009005f
C96 VTAIL.n61 B 0.021284f
C97 VTAIL.n62 B 0.009535f
C98 VTAIL.n63 B 0.016758f
C99 VTAIL.n64 B 0.009005f
C100 VTAIL.n65 B 0.021284f
C101 VTAIL.n66 B 0.009535f
C102 VTAIL.n67 B 0.016758f
C103 VTAIL.n68 B 0.009005f
C104 VTAIL.n69 B 0.021284f
C105 VTAIL.n70 B 0.009535f
C106 VTAIL.n71 B 0.016758f
C107 VTAIL.n72 B 0.009005f
C108 VTAIL.n73 B 0.021284f
C109 VTAIL.n74 B 0.009535f
C110 VTAIL.n75 B 0.113425f
C111 VTAIL.t2 B 0.035845f
C112 VTAIL.n76 B 0.015963f
C113 VTAIL.n77 B 0.015046f
C114 VTAIL.n78 B 0.009005f
C115 VTAIL.n79 B 0.759686f
C116 VTAIL.n80 B 0.016758f
C117 VTAIL.n81 B 0.009005f
C118 VTAIL.n82 B 0.009535f
C119 VTAIL.n83 B 0.021284f
C120 VTAIL.n84 B 0.021284f
C121 VTAIL.n85 B 0.009535f
C122 VTAIL.n86 B 0.009005f
C123 VTAIL.n87 B 0.016758f
C124 VTAIL.n88 B 0.016758f
C125 VTAIL.n89 B 0.009005f
C126 VTAIL.n90 B 0.009535f
C127 VTAIL.n91 B 0.021284f
C128 VTAIL.n92 B 0.021284f
C129 VTAIL.n93 B 0.021284f
C130 VTAIL.n94 B 0.009535f
C131 VTAIL.n95 B 0.009005f
C132 VTAIL.n96 B 0.016758f
C133 VTAIL.n97 B 0.016758f
C134 VTAIL.n98 B 0.009005f
C135 VTAIL.n99 B 0.00927f
C136 VTAIL.n100 B 0.00927f
C137 VTAIL.n101 B 0.021284f
C138 VTAIL.n102 B 0.021284f
C139 VTAIL.n103 B 0.009535f
C140 VTAIL.n104 B 0.009005f
C141 VTAIL.n105 B 0.016758f
C142 VTAIL.n106 B 0.016758f
C143 VTAIL.n107 B 0.009005f
C144 VTAIL.n108 B 0.009535f
C145 VTAIL.n109 B 0.021284f
C146 VTAIL.n110 B 0.047877f
C147 VTAIL.n111 B 0.009535f
C148 VTAIL.n112 B 0.009005f
C149 VTAIL.n113 B 0.042627f
C150 VTAIL.n114 B 0.027088f
C151 VTAIL.n115 B 0.178274f
C152 VTAIL.n116 B 0.024572f
C153 VTAIL.n117 B 0.016758f
C154 VTAIL.n118 B 0.009005f
C155 VTAIL.n119 B 0.021284f
C156 VTAIL.n120 B 0.009535f
C157 VTAIL.n121 B 0.016758f
C158 VTAIL.n122 B 0.009005f
C159 VTAIL.n123 B 0.021284f
C160 VTAIL.n124 B 0.009535f
C161 VTAIL.n125 B 0.016758f
C162 VTAIL.n126 B 0.009005f
C163 VTAIL.n127 B 0.021284f
C164 VTAIL.n128 B 0.009535f
C165 VTAIL.n129 B 0.016758f
C166 VTAIL.n130 B 0.009005f
C167 VTAIL.n131 B 0.021284f
C168 VTAIL.n132 B 0.009535f
C169 VTAIL.n133 B 0.113425f
C170 VTAIL.t3 B 0.035845f
C171 VTAIL.n134 B 0.015963f
C172 VTAIL.n135 B 0.015046f
C173 VTAIL.n136 B 0.009005f
C174 VTAIL.n137 B 0.759686f
C175 VTAIL.n138 B 0.016758f
C176 VTAIL.n139 B 0.009005f
C177 VTAIL.n140 B 0.009535f
C178 VTAIL.n141 B 0.021284f
C179 VTAIL.n142 B 0.021284f
C180 VTAIL.n143 B 0.009535f
C181 VTAIL.n144 B 0.009005f
C182 VTAIL.n145 B 0.016758f
C183 VTAIL.n146 B 0.016758f
C184 VTAIL.n147 B 0.009005f
C185 VTAIL.n148 B 0.009535f
C186 VTAIL.n149 B 0.021284f
C187 VTAIL.n150 B 0.021284f
C188 VTAIL.n151 B 0.021284f
C189 VTAIL.n152 B 0.009535f
C190 VTAIL.n153 B 0.009005f
C191 VTAIL.n154 B 0.016758f
C192 VTAIL.n155 B 0.016758f
C193 VTAIL.n156 B 0.009005f
C194 VTAIL.n157 B 0.00927f
C195 VTAIL.n158 B 0.00927f
C196 VTAIL.n159 B 0.021284f
C197 VTAIL.n160 B 0.021284f
C198 VTAIL.n161 B 0.009535f
C199 VTAIL.n162 B 0.009005f
C200 VTAIL.n163 B 0.016758f
C201 VTAIL.n164 B 0.016758f
C202 VTAIL.n165 B 0.009005f
C203 VTAIL.n166 B 0.009535f
C204 VTAIL.n167 B 0.021284f
C205 VTAIL.n168 B 0.047877f
C206 VTAIL.n169 B 0.009535f
C207 VTAIL.n170 B 0.009005f
C208 VTAIL.n171 B 0.042627f
C209 VTAIL.n172 B 0.027088f
C210 VTAIL.n173 B 1.02199f
C211 VTAIL.n174 B 0.024572f
C212 VTAIL.n175 B 0.016758f
C213 VTAIL.n176 B 0.009005f
C214 VTAIL.n177 B 0.021284f
C215 VTAIL.n178 B 0.009535f
C216 VTAIL.n179 B 0.016758f
C217 VTAIL.n180 B 0.009005f
C218 VTAIL.n181 B 0.021284f
C219 VTAIL.n182 B 0.009535f
C220 VTAIL.n183 B 0.016758f
C221 VTAIL.n184 B 0.009005f
C222 VTAIL.n185 B 0.021284f
C223 VTAIL.n186 B 0.021284f
C224 VTAIL.n187 B 0.009535f
C225 VTAIL.n188 B 0.016758f
C226 VTAIL.n189 B 0.009005f
C227 VTAIL.n190 B 0.021284f
C228 VTAIL.n191 B 0.009535f
C229 VTAIL.n192 B 0.113425f
C230 VTAIL.t0 B 0.035845f
C231 VTAIL.n193 B 0.015963f
C232 VTAIL.n194 B 0.015046f
C233 VTAIL.n195 B 0.009005f
C234 VTAIL.n196 B 0.759686f
C235 VTAIL.n197 B 0.016758f
C236 VTAIL.n198 B 0.009005f
C237 VTAIL.n199 B 0.009535f
C238 VTAIL.n200 B 0.021284f
C239 VTAIL.n201 B 0.021284f
C240 VTAIL.n202 B 0.009535f
C241 VTAIL.n203 B 0.009005f
C242 VTAIL.n204 B 0.016758f
C243 VTAIL.n205 B 0.016758f
C244 VTAIL.n206 B 0.009005f
C245 VTAIL.n207 B 0.009535f
C246 VTAIL.n208 B 0.021284f
C247 VTAIL.n209 B 0.021284f
C248 VTAIL.n210 B 0.009535f
C249 VTAIL.n211 B 0.009005f
C250 VTAIL.n212 B 0.016758f
C251 VTAIL.n213 B 0.016758f
C252 VTAIL.n214 B 0.009005f
C253 VTAIL.n215 B 0.00927f
C254 VTAIL.n216 B 0.00927f
C255 VTAIL.n217 B 0.021284f
C256 VTAIL.n218 B 0.021284f
C257 VTAIL.n219 B 0.009535f
C258 VTAIL.n220 B 0.009005f
C259 VTAIL.n221 B 0.016758f
C260 VTAIL.n222 B 0.016758f
C261 VTAIL.n223 B 0.009005f
C262 VTAIL.n224 B 0.009535f
C263 VTAIL.n225 B 0.021284f
C264 VTAIL.n226 B 0.047877f
C265 VTAIL.n227 B 0.009535f
C266 VTAIL.n228 B 0.009005f
C267 VTAIL.n229 B 0.042627f
C268 VTAIL.n230 B 0.027088f
C269 VTAIL.n231 B 1.02199f
C270 VTAIL.n232 B 0.024572f
C271 VTAIL.n233 B 0.016758f
C272 VTAIL.n234 B 0.009005f
C273 VTAIL.n235 B 0.021284f
C274 VTAIL.n236 B 0.009535f
C275 VTAIL.n237 B 0.016758f
C276 VTAIL.n238 B 0.009005f
C277 VTAIL.n239 B 0.021284f
C278 VTAIL.n240 B 0.009535f
C279 VTAIL.n241 B 0.016758f
C280 VTAIL.n242 B 0.009005f
C281 VTAIL.n243 B 0.021284f
C282 VTAIL.n244 B 0.021284f
C283 VTAIL.n245 B 0.009535f
C284 VTAIL.n246 B 0.016758f
C285 VTAIL.n247 B 0.009005f
C286 VTAIL.n248 B 0.021284f
C287 VTAIL.n249 B 0.009535f
C288 VTAIL.n250 B 0.113425f
C289 VTAIL.t5 B 0.035845f
C290 VTAIL.n251 B 0.015963f
C291 VTAIL.n252 B 0.015046f
C292 VTAIL.n253 B 0.009005f
C293 VTAIL.n254 B 0.759686f
C294 VTAIL.n255 B 0.016758f
C295 VTAIL.n256 B 0.009005f
C296 VTAIL.n257 B 0.009535f
C297 VTAIL.n258 B 0.021284f
C298 VTAIL.n259 B 0.021284f
C299 VTAIL.n260 B 0.009535f
C300 VTAIL.n261 B 0.009005f
C301 VTAIL.n262 B 0.016758f
C302 VTAIL.n263 B 0.016758f
C303 VTAIL.n264 B 0.009005f
C304 VTAIL.n265 B 0.009535f
C305 VTAIL.n266 B 0.021284f
C306 VTAIL.n267 B 0.021284f
C307 VTAIL.n268 B 0.009535f
C308 VTAIL.n269 B 0.009005f
C309 VTAIL.n270 B 0.016758f
C310 VTAIL.n271 B 0.016758f
C311 VTAIL.n272 B 0.009005f
C312 VTAIL.n273 B 0.00927f
C313 VTAIL.n274 B 0.00927f
C314 VTAIL.n275 B 0.021284f
C315 VTAIL.n276 B 0.021284f
C316 VTAIL.n277 B 0.009535f
C317 VTAIL.n278 B 0.009005f
C318 VTAIL.n279 B 0.016758f
C319 VTAIL.n280 B 0.016758f
C320 VTAIL.n281 B 0.009005f
C321 VTAIL.n282 B 0.009535f
C322 VTAIL.n283 B 0.021284f
C323 VTAIL.n284 B 0.047877f
C324 VTAIL.n285 B 0.009535f
C325 VTAIL.n286 B 0.009005f
C326 VTAIL.n287 B 0.042627f
C327 VTAIL.n288 B 0.027088f
C328 VTAIL.n289 B 0.178274f
C329 VTAIL.n290 B 0.024572f
C330 VTAIL.n291 B 0.016758f
C331 VTAIL.n292 B 0.009005f
C332 VTAIL.n293 B 0.021284f
C333 VTAIL.n294 B 0.009535f
C334 VTAIL.n295 B 0.016758f
C335 VTAIL.n296 B 0.009005f
C336 VTAIL.n297 B 0.021284f
C337 VTAIL.n298 B 0.009535f
C338 VTAIL.n299 B 0.016758f
C339 VTAIL.n300 B 0.009005f
C340 VTAIL.n301 B 0.021284f
C341 VTAIL.n302 B 0.021284f
C342 VTAIL.n303 B 0.009535f
C343 VTAIL.n304 B 0.016758f
C344 VTAIL.n305 B 0.009005f
C345 VTAIL.n306 B 0.021284f
C346 VTAIL.n307 B 0.009535f
C347 VTAIL.n308 B 0.113425f
C348 VTAIL.t4 B 0.035845f
C349 VTAIL.n309 B 0.015963f
C350 VTAIL.n310 B 0.015046f
C351 VTAIL.n311 B 0.009005f
C352 VTAIL.n312 B 0.759686f
C353 VTAIL.n313 B 0.016758f
C354 VTAIL.n314 B 0.009005f
C355 VTAIL.n315 B 0.009535f
C356 VTAIL.n316 B 0.021284f
C357 VTAIL.n317 B 0.021284f
C358 VTAIL.n318 B 0.009535f
C359 VTAIL.n319 B 0.009005f
C360 VTAIL.n320 B 0.016758f
C361 VTAIL.n321 B 0.016758f
C362 VTAIL.n322 B 0.009005f
C363 VTAIL.n323 B 0.009535f
C364 VTAIL.n324 B 0.021284f
C365 VTAIL.n325 B 0.021284f
C366 VTAIL.n326 B 0.009535f
C367 VTAIL.n327 B 0.009005f
C368 VTAIL.n328 B 0.016758f
C369 VTAIL.n329 B 0.016758f
C370 VTAIL.n330 B 0.009005f
C371 VTAIL.n331 B 0.00927f
C372 VTAIL.n332 B 0.00927f
C373 VTAIL.n333 B 0.021284f
C374 VTAIL.n334 B 0.021284f
C375 VTAIL.n335 B 0.009535f
C376 VTAIL.n336 B 0.009005f
C377 VTAIL.n337 B 0.016758f
C378 VTAIL.n338 B 0.016758f
C379 VTAIL.n339 B 0.009005f
C380 VTAIL.n340 B 0.009535f
C381 VTAIL.n341 B 0.021284f
C382 VTAIL.n342 B 0.047877f
C383 VTAIL.n343 B 0.009535f
C384 VTAIL.n344 B 0.009005f
C385 VTAIL.n345 B 0.042627f
C386 VTAIL.n346 B 0.027088f
C387 VTAIL.n347 B 0.178274f
C388 VTAIL.n348 B 0.024572f
C389 VTAIL.n349 B 0.016758f
C390 VTAIL.n350 B 0.009005f
C391 VTAIL.n351 B 0.021284f
C392 VTAIL.n352 B 0.009535f
C393 VTAIL.n353 B 0.016758f
C394 VTAIL.n354 B 0.009005f
C395 VTAIL.n355 B 0.021284f
C396 VTAIL.n356 B 0.009535f
C397 VTAIL.n357 B 0.016758f
C398 VTAIL.n358 B 0.009005f
C399 VTAIL.n359 B 0.021284f
C400 VTAIL.n360 B 0.021284f
C401 VTAIL.n361 B 0.009535f
C402 VTAIL.n362 B 0.016758f
C403 VTAIL.n363 B 0.009005f
C404 VTAIL.n364 B 0.021284f
C405 VTAIL.n365 B 0.009535f
C406 VTAIL.n366 B 0.113425f
C407 VTAIL.t1 B 0.035845f
C408 VTAIL.n367 B 0.015963f
C409 VTAIL.n368 B 0.015046f
C410 VTAIL.n369 B 0.009005f
C411 VTAIL.n370 B 0.759686f
C412 VTAIL.n371 B 0.016758f
C413 VTAIL.n372 B 0.009005f
C414 VTAIL.n373 B 0.009535f
C415 VTAIL.n374 B 0.021284f
C416 VTAIL.n375 B 0.021284f
C417 VTAIL.n376 B 0.009535f
C418 VTAIL.n377 B 0.009005f
C419 VTAIL.n378 B 0.016758f
C420 VTAIL.n379 B 0.016758f
C421 VTAIL.n380 B 0.009005f
C422 VTAIL.n381 B 0.009535f
C423 VTAIL.n382 B 0.021284f
C424 VTAIL.n383 B 0.021284f
C425 VTAIL.n384 B 0.009535f
C426 VTAIL.n385 B 0.009005f
C427 VTAIL.n386 B 0.016758f
C428 VTAIL.n387 B 0.016758f
C429 VTAIL.n388 B 0.009005f
C430 VTAIL.n389 B 0.00927f
C431 VTAIL.n390 B 0.00927f
C432 VTAIL.n391 B 0.021284f
C433 VTAIL.n392 B 0.021284f
C434 VTAIL.n393 B 0.009535f
C435 VTAIL.n394 B 0.009005f
C436 VTAIL.n395 B 0.016758f
C437 VTAIL.n396 B 0.016758f
C438 VTAIL.n397 B 0.009005f
C439 VTAIL.n398 B 0.009535f
C440 VTAIL.n399 B 0.021284f
C441 VTAIL.n400 B 0.047877f
C442 VTAIL.n401 B 0.009535f
C443 VTAIL.n402 B 0.009005f
C444 VTAIL.n403 B 0.042627f
C445 VTAIL.n404 B 0.027088f
C446 VTAIL.n405 B 1.02199f
C447 VTAIL.n406 B 0.024572f
C448 VTAIL.n407 B 0.016758f
C449 VTAIL.n408 B 0.009005f
C450 VTAIL.n409 B 0.021284f
C451 VTAIL.n410 B 0.009535f
C452 VTAIL.n411 B 0.016758f
C453 VTAIL.n412 B 0.009005f
C454 VTAIL.n413 B 0.021284f
C455 VTAIL.n414 B 0.009535f
C456 VTAIL.n415 B 0.016758f
C457 VTAIL.n416 B 0.009005f
C458 VTAIL.n417 B 0.021284f
C459 VTAIL.n418 B 0.009535f
C460 VTAIL.n419 B 0.016758f
C461 VTAIL.n420 B 0.009005f
C462 VTAIL.n421 B 0.021284f
C463 VTAIL.n422 B 0.009535f
C464 VTAIL.n423 B 0.113425f
C465 VTAIL.t6 B 0.035845f
C466 VTAIL.n424 B 0.015963f
C467 VTAIL.n425 B 0.015046f
C468 VTAIL.n426 B 0.009005f
C469 VTAIL.n427 B 0.759686f
C470 VTAIL.n428 B 0.016758f
C471 VTAIL.n429 B 0.009005f
C472 VTAIL.n430 B 0.009535f
C473 VTAIL.n431 B 0.021284f
C474 VTAIL.n432 B 0.021284f
C475 VTAIL.n433 B 0.009535f
C476 VTAIL.n434 B 0.009005f
C477 VTAIL.n435 B 0.016758f
C478 VTAIL.n436 B 0.016758f
C479 VTAIL.n437 B 0.009005f
C480 VTAIL.n438 B 0.009535f
C481 VTAIL.n439 B 0.021284f
C482 VTAIL.n440 B 0.021284f
C483 VTAIL.n441 B 0.021284f
C484 VTAIL.n442 B 0.009535f
C485 VTAIL.n443 B 0.009005f
C486 VTAIL.n444 B 0.016758f
C487 VTAIL.n445 B 0.016758f
C488 VTAIL.n446 B 0.009005f
C489 VTAIL.n447 B 0.00927f
C490 VTAIL.n448 B 0.00927f
C491 VTAIL.n449 B 0.021284f
C492 VTAIL.n450 B 0.021284f
C493 VTAIL.n451 B 0.009535f
C494 VTAIL.n452 B 0.009005f
C495 VTAIL.n453 B 0.016758f
C496 VTAIL.n454 B 0.016758f
C497 VTAIL.n455 B 0.009005f
C498 VTAIL.n456 B 0.009535f
C499 VTAIL.n457 B 0.021284f
C500 VTAIL.n458 B 0.047877f
C501 VTAIL.n459 B 0.009535f
C502 VTAIL.n460 B 0.009005f
C503 VTAIL.n461 B 0.042627f
C504 VTAIL.n462 B 0.027088f
C505 VTAIL.n463 B 0.950657f
C506 VP.n0 B 0.03479f
C507 VP.t1 B 2.02209f
C508 VP.n1 B 0.038522f
C509 VP.n2 B 0.026388f
C510 VP.t3 B 2.02209f
C511 VP.n3 B 0.809022f
C512 VP.t0 B 2.25306f
C513 VP.t2 B 2.25796f
C514 VP.n4 B 2.80165f
C515 VP.n5 B 1.42659f
C516 VP.n6 B 0.03479f
C517 VP.n7 B 0.03534f
C518 VP.n8 B 0.049181f
C519 VP.n9 B 0.038522f
C520 VP.n10 B 0.026388f
C521 VP.n11 B 0.026388f
C522 VP.n12 B 0.026388f
C523 VP.n13 B 0.049181f
C524 VP.n14 B 0.03534f
C525 VP.n15 B 0.809022f
C526 VP.n16 B 0.042563f
.ends

