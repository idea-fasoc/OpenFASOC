* NGSPICE file created from diff_pair_sample_1584.ext - technology: sky130A

.subckt diff_pair_sample_1584 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t8 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X1 VDD2.t9 VN.t0 VTAIL.t1 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X2 VDD1.t6 VP.t1 VTAIL.t10 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X3 VTAIL.t0 VN.t1 VDD2.t8 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X4 VTAIL.t9 VP.t2 VDD1.t1 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X5 VDD1.t9 VP.t3 VTAIL.t8 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=0.37
X6 VDD2.t7 VN.t2 VTAIL.t16 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=0.37
X7 VDD1.t7 VP.t4 VTAIL.t7 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=0.37
X8 VDD2.t6 VN.t3 VTAIL.t12 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X9 VDD1.t2 VP.t5 VTAIL.t6 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=0.37
X10 VTAIL.t18 VN.t4 VDD2.t5 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X11 VDD2.t4 VN.t5 VTAIL.t15 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=0.37
X12 VDD2.t3 VN.t6 VTAIL.t14 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=0.37
X13 VDD2.t2 VN.t7 VTAIL.t13 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=0.37
X14 VTAIL.t19 VN.t8 VDD2.t1 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X15 VTAIL.t17 VN.t9 VDD2.t0 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X16 VTAIL.t5 VP.t6 VDD1.t4 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X17 VTAIL.t4 VP.t7 VDD1.t5 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X18 B.t11 B.t9 B.t10 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=0.37
X19 VDD1.t3 VP.t8 VTAIL.t3 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=0.37
X20 B.t8 B.t6 B.t7 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=0.37
X21 VDD1.t0 VP.t9 VTAIL.t2 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=0.37
X22 B.t5 B.t3 B.t4 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=0.37
X23 B.t2 B.t0 B.t1 w_n1810_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=0.37
R0 VP.n5 VP.t5 385.087
R1 VP.n15 VP.t3 364.106
R2 VP.n16 VP.t0 364.106
R3 VP.n1 VP.t1 364.106
R4 VP.n21 VP.t7 364.106
R5 VP.n22 VP.t9 364.106
R6 VP.n12 VP.t4 364.106
R7 VP.n11 VP.t6 364.106
R8 VP.n4 VP.t8 364.106
R9 VP.n6 VP.t2 364.106
R10 VP.n23 VP.n22 161.3
R11 VP.n8 VP.n7 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n11 VP.n3 161.3
R14 VP.n13 VP.n12 161.3
R15 VP.n21 VP.n0 161.3
R16 VP.n20 VP.n19 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n2 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n8 VP.n5 70.4033
R21 VP.n16 VP.n15 48.2005
R22 VP.n22 VP.n21 48.2005
R23 VP.n12 VP.n11 48.2005
R24 VP.n17 VP.n16 38.7066
R25 VP.n21 VP.n20 38.7066
R26 VP.n11 VP.n10 38.7066
R27 VP.n7 VP.n6 38.7066
R28 VP.n14 VP.n13 34.8793
R29 VP.n6 VP.n5 20.9576
R30 VP.n17 VP.n1 9.49444
R31 VP.n20 VP.n1 9.49444
R32 VP.n10 VP.n4 9.49444
R33 VP.n7 VP.n4 9.49444
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n3 0.189894
R36 VP.n13 VP.n3 0.189894
R37 VP.n14 VP.n2 0.189894
R38 VP.n18 VP.n2 0.189894
R39 VP.n19 VP.n18 0.189894
R40 VP.n19 VP.n0 0.189894
R41 VP.n23 VP.n0 0.189894
R42 VP VP.n23 0.0516364
R43 VDD1.n14 VDD1.n0 756.745
R44 VDD1.n35 VDD1.n21 756.745
R45 VDD1.n15 VDD1.n14 585
R46 VDD1.n13 VDD1.n12 585
R47 VDD1.n4 VDD1.n3 585
R48 VDD1.n7 VDD1.n6 585
R49 VDD1.n28 VDD1.n27 585
R50 VDD1.n25 VDD1.n24 585
R51 VDD1.n34 VDD1.n33 585
R52 VDD1.n36 VDD1.n35 585
R53 VDD1.t2 VDD1.n5 330.707
R54 VDD1.t9 VDD1.n26 330.707
R55 VDD1.n14 VDD1.n13 171.744
R56 VDD1.n13 VDD1.n3 171.744
R57 VDD1.n6 VDD1.n3 171.744
R58 VDD1.n27 VDD1.n24 171.744
R59 VDD1.n34 VDD1.n24 171.744
R60 VDD1.n35 VDD1.n34 171.744
R61 VDD1.n43 VDD1.n42 116.099
R62 VDD1.n20 VDD1.n19 115.701
R63 VDD1.n45 VDD1.n44 115.701
R64 VDD1.n41 VDD1.n40 115.701
R65 VDD1.n6 VDD1.t2 85.8723
R66 VDD1.n27 VDD1.t9 85.8723
R67 VDD1.n20 VDD1.n18 51.6009
R68 VDD1.n41 VDD1.n39 51.6009
R69 VDD1.n45 VDD1.n43 30.8716
R70 VDD1.n7 VDD1.n5 16.3201
R71 VDD1.n28 VDD1.n26 16.3201
R72 VDD1.n8 VDD1.n4 12.8005
R73 VDD1.n29 VDD1.n25 12.8005
R74 VDD1.n12 VDD1.n11 12.0247
R75 VDD1.n33 VDD1.n32 12.0247
R76 VDD1.n15 VDD1.n2 11.249
R77 VDD1.n36 VDD1.n23 11.249
R78 VDD1.n16 VDD1.n0 10.4732
R79 VDD1.n37 VDD1.n21 10.4732
R80 VDD1.n18 VDD1.n17 9.45567
R81 VDD1.n39 VDD1.n38 9.45567
R82 VDD1.n17 VDD1.n16 9.3005
R83 VDD1.n2 VDD1.n1 9.3005
R84 VDD1.n11 VDD1.n10 9.3005
R85 VDD1.n9 VDD1.n8 9.3005
R86 VDD1.n38 VDD1.n37 9.3005
R87 VDD1.n23 VDD1.n22 9.3005
R88 VDD1.n32 VDD1.n31 9.3005
R89 VDD1.n30 VDD1.n29 9.3005
R90 VDD1.n44 VDD1.t4 8.22961
R91 VDD1.n44 VDD1.t7 8.22961
R92 VDD1.n19 VDD1.t1 8.22961
R93 VDD1.n19 VDD1.t3 8.22961
R94 VDD1.n42 VDD1.t5 8.22961
R95 VDD1.n42 VDD1.t0 8.22961
R96 VDD1.n40 VDD1.t8 8.22961
R97 VDD1.n40 VDD1.t6 8.22961
R98 VDD1.n9 VDD1.n5 3.78097
R99 VDD1.n30 VDD1.n26 3.78097
R100 VDD1.n18 VDD1.n0 3.49141
R101 VDD1.n39 VDD1.n21 3.49141
R102 VDD1.n16 VDD1.n15 2.71565
R103 VDD1.n37 VDD1.n36 2.71565
R104 VDD1.n12 VDD1.n2 1.93989
R105 VDD1.n33 VDD1.n23 1.93989
R106 VDD1.n11 VDD1.n4 1.16414
R107 VDD1.n32 VDD1.n25 1.16414
R108 VDD1 VDD1.n45 0.394897
R109 VDD1.n8 VDD1.n7 0.388379
R110 VDD1.n29 VDD1.n28 0.388379
R111 VDD1 VDD1.n20 0.209552
R112 VDD1.n17 VDD1.n1 0.155672
R113 VDD1.n10 VDD1.n1 0.155672
R114 VDD1.n10 VDD1.n9 0.155672
R115 VDD1.n31 VDD1.n30 0.155672
R116 VDD1.n31 VDD1.n22 0.155672
R117 VDD1.n38 VDD1.n22 0.155672
R118 VDD1.n43 VDD1.n41 0.096016
R119 VTAIL.n88 VTAIL.n74 756.745
R120 VTAIL.n16 VTAIL.n2 756.745
R121 VTAIL.n68 VTAIL.n54 756.745
R122 VTAIL.n44 VTAIL.n30 756.745
R123 VTAIL.n81 VTAIL.n80 585
R124 VTAIL.n78 VTAIL.n77 585
R125 VTAIL.n87 VTAIL.n86 585
R126 VTAIL.n89 VTAIL.n88 585
R127 VTAIL.n9 VTAIL.n8 585
R128 VTAIL.n6 VTAIL.n5 585
R129 VTAIL.n15 VTAIL.n14 585
R130 VTAIL.n17 VTAIL.n16 585
R131 VTAIL.n69 VTAIL.n68 585
R132 VTAIL.n67 VTAIL.n66 585
R133 VTAIL.n58 VTAIL.n57 585
R134 VTAIL.n61 VTAIL.n60 585
R135 VTAIL.n45 VTAIL.n44 585
R136 VTAIL.n43 VTAIL.n42 585
R137 VTAIL.n34 VTAIL.n33 585
R138 VTAIL.n37 VTAIL.n36 585
R139 VTAIL.t13 VTAIL.n79 330.707
R140 VTAIL.t2 VTAIL.n7 330.707
R141 VTAIL.t7 VTAIL.n59 330.707
R142 VTAIL.t16 VTAIL.n35 330.707
R143 VTAIL.n80 VTAIL.n77 171.744
R144 VTAIL.n87 VTAIL.n77 171.744
R145 VTAIL.n88 VTAIL.n87 171.744
R146 VTAIL.n8 VTAIL.n5 171.744
R147 VTAIL.n15 VTAIL.n5 171.744
R148 VTAIL.n16 VTAIL.n15 171.744
R149 VTAIL.n68 VTAIL.n67 171.744
R150 VTAIL.n67 VTAIL.n57 171.744
R151 VTAIL.n60 VTAIL.n57 171.744
R152 VTAIL.n44 VTAIL.n43 171.744
R153 VTAIL.n43 VTAIL.n33 171.744
R154 VTAIL.n36 VTAIL.n33 171.744
R155 VTAIL.n53 VTAIL.n52 99.0229
R156 VTAIL.n51 VTAIL.n50 99.0229
R157 VTAIL.n29 VTAIL.n28 99.0229
R158 VTAIL.n27 VTAIL.n26 99.0229
R159 VTAIL.n95 VTAIL.n94 99.0227
R160 VTAIL.n1 VTAIL.n0 99.0227
R161 VTAIL.n23 VTAIL.n22 99.0227
R162 VTAIL.n25 VTAIL.n24 99.0227
R163 VTAIL.n80 VTAIL.t13 85.8723
R164 VTAIL.n8 VTAIL.t2 85.8723
R165 VTAIL.n60 VTAIL.t7 85.8723
R166 VTAIL.n36 VTAIL.t16 85.8723
R167 VTAIL.n93 VTAIL.n92 34.3187
R168 VTAIL.n21 VTAIL.n20 34.3187
R169 VTAIL.n73 VTAIL.n72 34.3187
R170 VTAIL.n49 VTAIL.n48 34.3187
R171 VTAIL.n27 VTAIL.n25 16.9789
R172 VTAIL.n93 VTAIL.n73 16.3755
R173 VTAIL.n81 VTAIL.n79 16.3201
R174 VTAIL.n9 VTAIL.n7 16.3201
R175 VTAIL.n61 VTAIL.n59 16.3201
R176 VTAIL.n37 VTAIL.n35 16.3201
R177 VTAIL.n82 VTAIL.n78 12.8005
R178 VTAIL.n10 VTAIL.n6 12.8005
R179 VTAIL.n62 VTAIL.n58 12.8005
R180 VTAIL.n38 VTAIL.n34 12.8005
R181 VTAIL.n86 VTAIL.n85 12.0247
R182 VTAIL.n14 VTAIL.n13 12.0247
R183 VTAIL.n66 VTAIL.n65 12.0247
R184 VTAIL.n42 VTAIL.n41 12.0247
R185 VTAIL.n89 VTAIL.n76 11.249
R186 VTAIL.n17 VTAIL.n4 11.249
R187 VTAIL.n69 VTAIL.n56 11.249
R188 VTAIL.n45 VTAIL.n32 11.249
R189 VTAIL.n90 VTAIL.n74 10.4732
R190 VTAIL.n18 VTAIL.n2 10.4732
R191 VTAIL.n70 VTAIL.n54 10.4732
R192 VTAIL.n46 VTAIL.n30 10.4732
R193 VTAIL.n92 VTAIL.n91 9.45567
R194 VTAIL.n20 VTAIL.n19 9.45567
R195 VTAIL.n72 VTAIL.n71 9.45567
R196 VTAIL.n48 VTAIL.n47 9.45567
R197 VTAIL.n91 VTAIL.n90 9.3005
R198 VTAIL.n76 VTAIL.n75 9.3005
R199 VTAIL.n85 VTAIL.n84 9.3005
R200 VTAIL.n83 VTAIL.n82 9.3005
R201 VTAIL.n19 VTAIL.n18 9.3005
R202 VTAIL.n4 VTAIL.n3 9.3005
R203 VTAIL.n13 VTAIL.n12 9.3005
R204 VTAIL.n11 VTAIL.n10 9.3005
R205 VTAIL.n71 VTAIL.n70 9.3005
R206 VTAIL.n56 VTAIL.n55 9.3005
R207 VTAIL.n65 VTAIL.n64 9.3005
R208 VTAIL.n63 VTAIL.n62 9.3005
R209 VTAIL.n47 VTAIL.n46 9.3005
R210 VTAIL.n32 VTAIL.n31 9.3005
R211 VTAIL.n41 VTAIL.n40 9.3005
R212 VTAIL.n39 VTAIL.n38 9.3005
R213 VTAIL.n94 VTAIL.t12 8.22961
R214 VTAIL.n94 VTAIL.t17 8.22961
R215 VTAIL.n0 VTAIL.t15 8.22961
R216 VTAIL.n0 VTAIL.t18 8.22961
R217 VTAIL.n22 VTAIL.t10 8.22961
R218 VTAIL.n22 VTAIL.t4 8.22961
R219 VTAIL.n24 VTAIL.t8 8.22961
R220 VTAIL.n24 VTAIL.t11 8.22961
R221 VTAIL.n52 VTAIL.t3 8.22961
R222 VTAIL.n52 VTAIL.t5 8.22961
R223 VTAIL.n50 VTAIL.t6 8.22961
R224 VTAIL.n50 VTAIL.t9 8.22961
R225 VTAIL.n28 VTAIL.t1 8.22961
R226 VTAIL.n28 VTAIL.t0 8.22961
R227 VTAIL.n26 VTAIL.t14 8.22961
R228 VTAIL.n26 VTAIL.t19 8.22961
R229 VTAIL.n83 VTAIL.n79 3.78097
R230 VTAIL.n11 VTAIL.n7 3.78097
R231 VTAIL.n63 VTAIL.n59 3.78097
R232 VTAIL.n39 VTAIL.n35 3.78097
R233 VTAIL.n92 VTAIL.n74 3.49141
R234 VTAIL.n20 VTAIL.n2 3.49141
R235 VTAIL.n72 VTAIL.n54 3.49141
R236 VTAIL.n48 VTAIL.n30 3.49141
R237 VTAIL.n90 VTAIL.n89 2.71565
R238 VTAIL.n18 VTAIL.n17 2.71565
R239 VTAIL.n70 VTAIL.n69 2.71565
R240 VTAIL.n46 VTAIL.n45 2.71565
R241 VTAIL.n86 VTAIL.n76 1.93989
R242 VTAIL.n14 VTAIL.n4 1.93989
R243 VTAIL.n66 VTAIL.n56 1.93989
R244 VTAIL.n42 VTAIL.n32 1.93989
R245 VTAIL.n85 VTAIL.n78 1.16414
R246 VTAIL.n13 VTAIL.n6 1.16414
R247 VTAIL.n65 VTAIL.n58 1.16414
R248 VTAIL.n41 VTAIL.n34 1.16414
R249 VTAIL.n51 VTAIL.n49 0.772052
R250 VTAIL.n21 VTAIL.n1 0.772052
R251 VTAIL.n29 VTAIL.n27 0.603948
R252 VTAIL.n49 VTAIL.n29 0.603948
R253 VTAIL.n53 VTAIL.n51 0.603948
R254 VTAIL.n73 VTAIL.n53 0.603948
R255 VTAIL.n25 VTAIL.n23 0.603948
R256 VTAIL.n23 VTAIL.n21 0.603948
R257 VTAIL.n95 VTAIL.n93 0.603948
R258 VTAIL VTAIL.n1 0.511276
R259 VTAIL.n82 VTAIL.n81 0.388379
R260 VTAIL.n10 VTAIL.n9 0.388379
R261 VTAIL.n62 VTAIL.n61 0.388379
R262 VTAIL.n38 VTAIL.n37 0.388379
R263 VTAIL.n84 VTAIL.n83 0.155672
R264 VTAIL.n84 VTAIL.n75 0.155672
R265 VTAIL.n91 VTAIL.n75 0.155672
R266 VTAIL.n12 VTAIL.n11 0.155672
R267 VTAIL.n12 VTAIL.n3 0.155672
R268 VTAIL.n19 VTAIL.n3 0.155672
R269 VTAIL.n71 VTAIL.n55 0.155672
R270 VTAIL.n64 VTAIL.n55 0.155672
R271 VTAIL.n64 VTAIL.n63 0.155672
R272 VTAIL.n47 VTAIL.n31 0.155672
R273 VTAIL.n40 VTAIL.n31 0.155672
R274 VTAIL.n40 VTAIL.n39 0.155672
R275 VTAIL VTAIL.n95 0.0931724
R276 VN.n2 VN.t5 385.087
R277 VN.n13 VN.t2 385.087
R278 VN.n3 VN.t4 364.106
R279 VN.n1 VN.t3 364.106
R280 VN.n8 VN.t9 364.106
R281 VN.n9 VN.t7 364.106
R282 VN.n14 VN.t1 364.106
R283 VN.n12 VN.t0 364.106
R284 VN.n19 VN.t8 364.106
R285 VN.n20 VN.t6 364.106
R286 VN.n10 VN.n9 161.3
R287 VN.n21 VN.n20 161.3
R288 VN.n19 VN.n11 161.3
R289 VN.n18 VN.n17 161.3
R290 VN.n16 VN.n15 161.3
R291 VN.n8 VN.n0 161.3
R292 VN.n7 VN.n6 161.3
R293 VN.n5 VN.n4 161.3
R294 VN.n16 VN.n13 70.4033
R295 VN.n5 VN.n2 70.4033
R296 VN.n9 VN.n8 48.2005
R297 VN.n20 VN.n19 48.2005
R298 VN.n4 VN.n3 38.7066
R299 VN.n8 VN.n7 38.7066
R300 VN.n15 VN.n14 38.7066
R301 VN.n19 VN.n18 38.7066
R302 VN VN.n21 35.26
R303 VN.n14 VN.n13 20.9576
R304 VN.n3 VN.n2 20.9576
R305 VN.n4 VN.n1 9.49444
R306 VN.n7 VN.n1 9.49444
R307 VN.n15 VN.n12 9.49444
R308 VN.n18 VN.n12 9.49444
R309 VN.n21 VN.n11 0.189894
R310 VN.n17 VN.n11 0.189894
R311 VN.n17 VN.n16 0.189894
R312 VN.n6 VN.n5 0.189894
R313 VN.n6 VN.n0 0.189894
R314 VN.n10 VN.n0 0.189894
R315 VN VN.n10 0.0516364
R316 VDD2.n37 VDD2.n23 756.745
R317 VDD2.n14 VDD2.n0 756.745
R318 VDD2.n38 VDD2.n37 585
R319 VDD2.n36 VDD2.n35 585
R320 VDD2.n27 VDD2.n26 585
R321 VDD2.n30 VDD2.n29 585
R322 VDD2.n7 VDD2.n6 585
R323 VDD2.n4 VDD2.n3 585
R324 VDD2.n13 VDD2.n12 585
R325 VDD2.n15 VDD2.n14 585
R326 VDD2.t3 VDD2.n28 330.707
R327 VDD2.t4 VDD2.n5 330.707
R328 VDD2.n37 VDD2.n36 171.744
R329 VDD2.n36 VDD2.n26 171.744
R330 VDD2.n29 VDD2.n26 171.744
R331 VDD2.n6 VDD2.n3 171.744
R332 VDD2.n13 VDD2.n3 171.744
R333 VDD2.n14 VDD2.n13 171.744
R334 VDD2.n22 VDD2.n21 116.099
R335 VDD2 VDD2.n45 116.096
R336 VDD2.n44 VDD2.n43 115.701
R337 VDD2.n20 VDD2.n19 115.701
R338 VDD2.n29 VDD2.t3 85.8723
R339 VDD2.n6 VDD2.t4 85.8723
R340 VDD2.n20 VDD2.n18 51.6009
R341 VDD2.n42 VDD2.n41 50.9975
R342 VDD2.n42 VDD2.n22 29.9868
R343 VDD2.n30 VDD2.n28 16.3201
R344 VDD2.n7 VDD2.n5 16.3201
R345 VDD2.n31 VDD2.n27 12.8005
R346 VDD2.n8 VDD2.n4 12.8005
R347 VDD2.n35 VDD2.n34 12.0247
R348 VDD2.n12 VDD2.n11 12.0247
R349 VDD2.n38 VDD2.n25 11.249
R350 VDD2.n15 VDD2.n2 11.249
R351 VDD2.n39 VDD2.n23 10.4732
R352 VDD2.n16 VDD2.n0 10.4732
R353 VDD2.n41 VDD2.n40 9.45567
R354 VDD2.n18 VDD2.n17 9.45567
R355 VDD2.n40 VDD2.n39 9.3005
R356 VDD2.n25 VDD2.n24 9.3005
R357 VDD2.n34 VDD2.n33 9.3005
R358 VDD2.n32 VDD2.n31 9.3005
R359 VDD2.n17 VDD2.n16 9.3005
R360 VDD2.n2 VDD2.n1 9.3005
R361 VDD2.n11 VDD2.n10 9.3005
R362 VDD2.n9 VDD2.n8 9.3005
R363 VDD2.n45 VDD2.t8 8.22961
R364 VDD2.n45 VDD2.t7 8.22961
R365 VDD2.n43 VDD2.t1 8.22961
R366 VDD2.n43 VDD2.t9 8.22961
R367 VDD2.n21 VDD2.t0 8.22961
R368 VDD2.n21 VDD2.t2 8.22961
R369 VDD2.n19 VDD2.t5 8.22961
R370 VDD2.n19 VDD2.t6 8.22961
R371 VDD2.n32 VDD2.n28 3.78097
R372 VDD2.n9 VDD2.n5 3.78097
R373 VDD2.n41 VDD2.n23 3.49141
R374 VDD2.n18 VDD2.n0 3.49141
R375 VDD2.n39 VDD2.n38 2.71565
R376 VDD2.n16 VDD2.n15 2.71565
R377 VDD2.n35 VDD2.n25 1.93989
R378 VDD2.n12 VDD2.n2 1.93989
R379 VDD2.n34 VDD2.n27 1.16414
R380 VDD2.n11 VDD2.n4 1.16414
R381 VDD2.n44 VDD2.n42 0.603948
R382 VDD2.n31 VDD2.n30 0.388379
R383 VDD2.n8 VDD2.n7 0.388379
R384 VDD2 VDD2.n44 0.209552
R385 VDD2.n40 VDD2.n24 0.155672
R386 VDD2.n33 VDD2.n24 0.155672
R387 VDD2.n33 VDD2.n32 0.155672
R388 VDD2.n10 VDD2.n9 0.155672
R389 VDD2.n10 VDD2.n1 0.155672
R390 VDD2.n17 VDD2.n1 0.155672
R391 VDD2.n22 VDD2.n20 0.096016
R392 B.n193 B.n192 585
R393 B.n191 B.n60 585
R394 B.n190 B.n189 585
R395 B.n188 B.n61 585
R396 B.n187 B.n186 585
R397 B.n185 B.n62 585
R398 B.n184 B.n183 585
R399 B.n182 B.n63 585
R400 B.n181 B.n180 585
R401 B.n179 B.n64 585
R402 B.n178 B.n177 585
R403 B.n176 B.n65 585
R404 B.n175 B.n174 585
R405 B.n173 B.n66 585
R406 B.n172 B.n171 585
R407 B.n170 B.n67 585
R408 B.n169 B.n168 585
R409 B.n167 B.n68 585
R410 B.n166 B.n165 585
R411 B.n161 B.n69 585
R412 B.n160 B.n159 585
R413 B.n158 B.n70 585
R414 B.n157 B.n156 585
R415 B.n155 B.n71 585
R416 B.n154 B.n153 585
R417 B.n152 B.n72 585
R418 B.n151 B.n150 585
R419 B.n148 B.n73 585
R420 B.n147 B.n146 585
R421 B.n145 B.n76 585
R422 B.n144 B.n143 585
R423 B.n142 B.n77 585
R424 B.n141 B.n140 585
R425 B.n139 B.n78 585
R426 B.n138 B.n137 585
R427 B.n136 B.n79 585
R428 B.n135 B.n134 585
R429 B.n133 B.n80 585
R430 B.n132 B.n131 585
R431 B.n130 B.n81 585
R432 B.n129 B.n128 585
R433 B.n127 B.n82 585
R434 B.n126 B.n125 585
R435 B.n124 B.n83 585
R436 B.n123 B.n122 585
R437 B.n194 B.n59 585
R438 B.n196 B.n195 585
R439 B.n197 B.n58 585
R440 B.n199 B.n198 585
R441 B.n200 B.n57 585
R442 B.n202 B.n201 585
R443 B.n203 B.n56 585
R444 B.n205 B.n204 585
R445 B.n206 B.n55 585
R446 B.n208 B.n207 585
R447 B.n209 B.n54 585
R448 B.n211 B.n210 585
R449 B.n212 B.n53 585
R450 B.n214 B.n213 585
R451 B.n215 B.n52 585
R452 B.n217 B.n216 585
R453 B.n218 B.n51 585
R454 B.n220 B.n219 585
R455 B.n221 B.n50 585
R456 B.n223 B.n222 585
R457 B.n224 B.n49 585
R458 B.n226 B.n225 585
R459 B.n227 B.n48 585
R460 B.n229 B.n228 585
R461 B.n230 B.n47 585
R462 B.n232 B.n231 585
R463 B.n233 B.n46 585
R464 B.n235 B.n234 585
R465 B.n236 B.n45 585
R466 B.n238 B.n237 585
R467 B.n239 B.n44 585
R468 B.n241 B.n240 585
R469 B.n242 B.n43 585
R470 B.n244 B.n243 585
R471 B.n245 B.n42 585
R472 B.n247 B.n246 585
R473 B.n248 B.n41 585
R474 B.n250 B.n249 585
R475 B.n251 B.n40 585
R476 B.n253 B.n252 585
R477 B.n254 B.n39 585
R478 B.n256 B.n255 585
R479 B.n325 B.n12 585
R480 B.n324 B.n323 585
R481 B.n322 B.n13 585
R482 B.n321 B.n320 585
R483 B.n319 B.n14 585
R484 B.n318 B.n317 585
R485 B.n316 B.n15 585
R486 B.n315 B.n314 585
R487 B.n313 B.n16 585
R488 B.n312 B.n311 585
R489 B.n310 B.n17 585
R490 B.n309 B.n308 585
R491 B.n307 B.n18 585
R492 B.n306 B.n305 585
R493 B.n304 B.n19 585
R494 B.n303 B.n302 585
R495 B.n301 B.n20 585
R496 B.n300 B.n299 585
R497 B.n297 B.n21 585
R498 B.n296 B.n295 585
R499 B.n294 B.n24 585
R500 B.n293 B.n292 585
R501 B.n291 B.n25 585
R502 B.n290 B.n289 585
R503 B.n288 B.n26 585
R504 B.n287 B.n286 585
R505 B.n285 B.n27 585
R506 B.n283 B.n282 585
R507 B.n281 B.n30 585
R508 B.n280 B.n279 585
R509 B.n278 B.n31 585
R510 B.n277 B.n276 585
R511 B.n275 B.n32 585
R512 B.n274 B.n273 585
R513 B.n272 B.n33 585
R514 B.n271 B.n270 585
R515 B.n269 B.n34 585
R516 B.n268 B.n267 585
R517 B.n266 B.n35 585
R518 B.n265 B.n264 585
R519 B.n263 B.n36 585
R520 B.n262 B.n261 585
R521 B.n260 B.n37 585
R522 B.n259 B.n258 585
R523 B.n257 B.n38 585
R524 B.n327 B.n326 585
R525 B.n328 B.n11 585
R526 B.n330 B.n329 585
R527 B.n331 B.n10 585
R528 B.n333 B.n332 585
R529 B.n334 B.n9 585
R530 B.n336 B.n335 585
R531 B.n337 B.n8 585
R532 B.n339 B.n338 585
R533 B.n340 B.n7 585
R534 B.n342 B.n341 585
R535 B.n343 B.n6 585
R536 B.n345 B.n344 585
R537 B.n346 B.n5 585
R538 B.n348 B.n347 585
R539 B.n349 B.n4 585
R540 B.n351 B.n350 585
R541 B.n352 B.n3 585
R542 B.n354 B.n353 585
R543 B.n355 B.n0 585
R544 B.n2 B.n1 585
R545 B.n94 B.n93 585
R546 B.n96 B.n95 585
R547 B.n97 B.n92 585
R548 B.n99 B.n98 585
R549 B.n100 B.n91 585
R550 B.n102 B.n101 585
R551 B.n103 B.n90 585
R552 B.n105 B.n104 585
R553 B.n106 B.n89 585
R554 B.n108 B.n107 585
R555 B.n109 B.n88 585
R556 B.n111 B.n110 585
R557 B.n112 B.n87 585
R558 B.n114 B.n113 585
R559 B.n115 B.n86 585
R560 B.n117 B.n116 585
R561 B.n118 B.n85 585
R562 B.n120 B.n119 585
R563 B.n121 B.n84 585
R564 B.n122 B.n121 530.939
R565 B.n192 B.n59 530.939
R566 B.n257 B.n256 530.939
R567 B.n326 B.n325 530.939
R568 B.n74 B.t9 467.925
R569 B.n162 B.t6 467.925
R570 B.n28 B.t0 467.925
R571 B.n22 B.t3 467.925
R572 B.n357 B.n356 256.663
R573 B.n162 B.t7 248.236
R574 B.n28 B.t2 248.236
R575 B.n74 B.t10 248.236
R576 B.n22 B.t5 248.236
R577 B.n356 B.n355 235.042
R578 B.n356 B.n2 235.042
R579 B.n163 B.t8 234.66
R580 B.n29 B.t1 234.66
R581 B.n75 B.t11 234.66
R582 B.n23 B.t4 234.66
R583 B.n122 B.n83 163.367
R584 B.n126 B.n83 163.367
R585 B.n127 B.n126 163.367
R586 B.n128 B.n127 163.367
R587 B.n128 B.n81 163.367
R588 B.n132 B.n81 163.367
R589 B.n133 B.n132 163.367
R590 B.n134 B.n133 163.367
R591 B.n134 B.n79 163.367
R592 B.n138 B.n79 163.367
R593 B.n139 B.n138 163.367
R594 B.n140 B.n139 163.367
R595 B.n140 B.n77 163.367
R596 B.n144 B.n77 163.367
R597 B.n145 B.n144 163.367
R598 B.n146 B.n145 163.367
R599 B.n146 B.n73 163.367
R600 B.n151 B.n73 163.367
R601 B.n152 B.n151 163.367
R602 B.n153 B.n152 163.367
R603 B.n153 B.n71 163.367
R604 B.n157 B.n71 163.367
R605 B.n158 B.n157 163.367
R606 B.n159 B.n158 163.367
R607 B.n159 B.n69 163.367
R608 B.n166 B.n69 163.367
R609 B.n167 B.n166 163.367
R610 B.n168 B.n167 163.367
R611 B.n168 B.n67 163.367
R612 B.n172 B.n67 163.367
R613 B.n173 B.n172 163.367
R614 B.n174 B.n173 163.367
R615 B.n174 B.n65 163.367
R616 B.n178 B.n65 163.367
R617 B.n179 B.n178 163.367
R618 B.n180 B.n179 163.367
R619 B.n180 B.n63 163.367
R620 B.n184 B.n63 163.367
R621 B.n185 B.n184 163.367
R622 B.n186 B.n185 163.367
R623 B.n186 B.n61 163.367
R624 B.n190 B.n61 163.367
R625 B.n191 B.n190 163.367
R626 B.n192 B.n191 163.367
R627 B.n256 B.n39 163.367
R628 B.n252 B.n39 163.367
R629 B.n252 B.n251 163.367
R630 B.n251 B.n250 163.367
R631 B.n250 B.n41 163.367
R632 B.n246 B.n41 163.367
R633 B.n246 B.n245 163.367
R634 B.n245 B.n244 163.367
R635 B.n244 B.n43 163.367
R636 B.n240 B.n43 163.367
R637 B.n240 B.n239 163.367
R638 B.n239 B.n238 163.367
R639 B.n238 B.n45 163.367
R640 B.n234 B.n45 163.367
R641 B.n234 B.n233 163.367
R642 B.n233 B.n232 163.367
R643 B.n232 B.n47 163.367
R644 B.n228 B.n47 163.367
R645 B.n228 B.n227 163.367
R646 B.n227 B.n226 163.367
R647 B.n226 B.n49 163.367
R648 B.n222 B.n49 163.367
R649 B.n222 B.n221 163.367
R650 B.n221 B.n220 163.367
R651 B.n220 B.n51 163.367
R652 B.n216 B.n51 163.367
R653 B.n216 B.n215 163.367
R654 B.n215 B.n214 163.367
R655 B.n214 B.n53 163.367
R656 B.n210 B.n53 163.367
R657 B.n210 B.n209 163.367
R658 B.n209 B.n208 163.367
R659 B.n208 B.n55 163.367
R660 B.n204 B.n55 163.367
R661 B.n204 B.n203 163.367
R662 B.n203 B.n202 163.367
R663 B.n202 B.n57 163.367
R664 B.n198 B.n57 163.367
R665 B.n198 B.n197 163.367
R666 B.n197 B.n196 163.367
R667 B.n196 B.n59 163.367
R668 B.n325 B.n324 163.367
R669 B.n324 B.n13 163.367
R670 B.n320 B.n13 163.367
R671 B.n320 B.n319 163.367
R672 B.n319 B.n318 163.367
R673 B.n318 B.n15 163.367
R674 B.n314 B.n15 163.367
R675 B.n314 B.n313 163.367
R676 B.n313 B.n312 163.367
R677 B.n312 B.n17 163.367
R678 B.n308 B.n17 163.367
R679 B.n308 B.n307 163.367
R680 B.n307 B.n306 163.367
R681 B.n306 B.n19 163.367
R682 B.n302 B.n19 163.367
R683 B.n302 B.n301 163.367
R684 B.n301 B.n300 163.367
R685 B.n300 B.n21 163.367
R686 B.n295 B.n21 163.367
R687 B.n295 B.n294 163.367
R688 B.n294 B.n293 163.367
R689 B.n293 B.n25 163.367
R690 B.n289 B.n25 163.367
R691 B.n289 B.n288 163.367
R692 B.n288 B.n287 163.367
R693 B.n287 B.n27 163.367
R694 B.n282 B.n27 163.367
R695 B.n282 B.n281 163.367
R696 B.n281 B.n280 163.367
R697 B.n280 B.n31 163.367
R698 B.n276 B.n31 163.367
R699 B.n276 B.n275 163.367
R700 B.n275 B.n274 163.367
R701 B.n274 B.n33 163.367
R702 B.n270 B.n33 163.367
R703 B.n270 B.n269 163.367
R704 B.n269 B.n268 163.367
R705 B.n268 B.n35 163.367
R706 B.n264 B.n35 163.367
R707 B.n264 B.n263 163.367
R708 B.n263 B.n262 163.367
R709 B.n262 B.n37 163.367
R710 B.n258 B.n37 163.367
R711 B.n258 B.n257 163.367
R712 B.n326 B.n11 163.367
R713 B.n330 B.n11 163.367
R714 B.n331 B.n330 163.367
R715 B.n332 B.n331 163.367
R716 B.n332 B.n9 163.367
R717 B.n336 B.n9 163.367
R718 B.n337 B.n336 163.367
R719 B.n338 B.n337 163.367
R720 B.n338 B.n7 163.367
R721 B.n342 B.n7 163.367
R722 B.n343 B.n342 163.367
R723 B.n344 B.n343 163.367
R724 B.n344 B.n5 163.367
R725 B.n348 B.n5 163.367
R726 B.n349 B.n348 163.367
R727 B.n350 B.n349 163.367
R728 B.n350 B.n3 163.367
R729 B.n354 B.n3 163.367
R730 B.n355 B.n354 163.367
R731 B.n93 B.n2 163.367
R732 B.n96 B.n93 163.367
R733 B.n97 B.n96 163.367
R734 B.n98 B.n97 163.367
R735 B.n98 B.n91 163.367
R736 B.n102 B.n91 163.367
R737 B.n103 B.n102 163.367
R738 B.n104 B.n103 163.367
R739 B.n104 B.n89 163.367
R740 B.n108 B.n89 163.367
R741 B.n109 B.n108 163.367
R742 B.n110 B.n109 163.367
R743 B.n110 B.n87 163.367
R744 B.n114 B.n87 163.367
R745 B.n115 B.n114 163.367
R746 B.n116 B.n115 163.367
R747 B.n116 B.n85 163.367
R748 B.n120 B.n85 163.367
R749 B.n121 B.n120 163.367
R750 B.n149 B.n75 59.5399
R751 B.n164 B.n163 59.5399
R752 B.n284 B.n29 59.5399
R753 B.n298 B.n23 59.5399
R754 B.n327 B.n12 34.4981
R755 B.n255 B.n38 34.4981
R756 B.n194 B.n193 34.4981
R757 B.n123 B.n84 34.4981
R758 B B.n357 18.0485
R759 B.n75 B.n74 13.5763
R760 B.n163 B.n162 13.5763
R761 B.n29 B.n28 13.5763
R762 B.n23 B.n22 13.5763
R763 B.n328 B.n327 10.6151
R764 B.n329 B.n328 10.6151
R765 B.n329 B.n10 10.6151
R766 B.n333 B.n10 10.6151
R767 B.n334 B.n333 10.6151
R768 B.n335 B.n334 10.6151
R769 B.n335 B.n8 10.6151
R770 B.n339 B.n8 10.6151
R771 B.n340 B.n339 10.6151
R772 B.n341 B.n340 10.6151
R773 B.n341 B.n6 10.6151
R774 B.n345 B.n6 10.6151
R775 B.n346 B.n345 10.6151
R776 B.n347 B.n346 10.6151
R777 B.n347 B.n4 10.6151
R778 B.n351 B.n4 10.6151
R779 B.n352 B.n351 10.6151
R780 B.n353 B.n352 10.6151
R781 B.n353 B.n0 10.6151
R782 B.n323 B.n12 10.6151
R783 B.n323 B.n322 10.6151
R784 B.n322 B.n321 10.6151
R785 B.n321 B.n14 10.6151
R786 B.n317 B.n14 10.6151
R787 B.n317 B.n316 10.6151
R788 B.n316 B.n315 10.6151
R789 B.n315 B.n16 10.6151
R790 B.n311 B.n16 10.6151
R791 B.n311 B.n310 10.6151
R792 B.n310 B.n309 10.6151
R793 B.n309 B.n18 10.6151
R794 B.n305 B.n18 10.6151
R795 B.n305 B.n304 10.6151
R796 B.n304 B.n303 10.6151
R797 B.n303 B.n20 10.6151
R798 B.n299 B.n20 10.6151
R799 B.n297 B.n296 10.6151
R800 B.n296 B.n24 10.6151
R801 B.n292 B.n24 10.6151
R802 B.n292 B.n291 10.6151
R803 B.n291 B.n290 10.6151
R804 B.n290 B.n26 10.6151
R805 B.n286 B.n26 10.6151
R806 B.n286 B.n285 10.6151
R807 B.n283 B.n30 10.6151
R808 B.n279 B.n30 10.6151
R809 B.n279 B.n278 10.6151
R810 B.n278 B.n277 10.6151
R811 B.n277 B.n32 10.6151
R812 B.n273 B.n32 10.6151
R813 B.n273 B.n272 10.6151
R814 B.n272 B.n271 10.6151
R815 B.n271 B.n34 10.6151
R816 B.n267 B.n34 10.6151
R817 B.n267 B.n266 10.6151
R818 B.n266 B.n265 10.6151
R819 B.n265 B.n36 10.6151
R820 B.n261 B.n36 10.6151
R821 B.n261 B.n260 10.6151
R822 B.n260 B.n259 10.6151
R823 B.n259 B.n38 10.6151
R824 B.n255 B.n254 10.6151
R825 B.n254 B.n253 10.6151
R826 B.n253 B.n40 10.6151
R827 B.n249 B.n40 10.6151
R828 B.n249 B.n248 10.6151
R829 B.n248 B.n247 10.6151
R830 B.n247 B.n42 10.6151
R831 B.n243 B.n42 10.6151
R832 B.n243 B.n242 10.6151
R833 B.n242 B.n241 10.6151
R834 B.n241 B.n44 10.6151
R835 B.n237 B.n44 10.6151
R836 B.n237 B.n236 10.6151
R837 B.n236 B.n235 10.6151
R838 B.n235 B.n46 10.6151
R839 B.n231 B.n46 10.6151
R840 B.n231 B.n230 10.6151
R841 B.n230 B.n229 10.6151
R842 B.n229 B.n48 10.6151
R843 B.n225 B.n48 10.6151
R844 B.n225 B.n224 10.6151
R845 B.n224 B.n223 10.6151
R846 B.n223 B.n50 10.6151
R847 B.n219 B.n50 10.6151
R848 B.n219 B.n218 10.6151
R849 B.n218 B.n217 10.6151
R850 B.n217 B.n52 10.6151
R851 B.n213 B.n52 10.6151
R852 B.n213 B.n212 10.6151
R853 B.n212 B.n211 10.6151
R854 B.n211 B.n54 10.6151
R855 B.n207 B.n54 10.6151
R856 B.n207 B.n206 10.6151
R857 B.n206 B.n205 10.6151
R858 B.n205 B.n56 10.6151
R859 B.n201 B.n56 10.6151
R860 B.n201 B.n200 10.6151
R861 B.n200 B.n199 10.6151
R862 B.n199 B.n58 10.6151
R863 B.n195 B.n58 10.6151
R864 B.n195 B.n194 10.6151
R865 B.n94 B.n1 10.6151
R866 B.n95 B.n94 10.6151
R867 B.n95 B.n92 10.6151
R868 B.n99 B.n92 10.6151
R869 B.n100 B.n99 10.6151
R870 B.n101 B.n100 10.6151
R871 B.n101 B.n90 10.6151
R872 B.n105 B.n90 10.6151
R873 B.n106 B.n105 10.6151
R874 B.n107 B.n106 10.6151
R875 B.n107 B.n88 10.6151
R876 B.n111 B.n88 10.6151
R877 B.n112 B.n111 10.6151
R878 B.n113 B.n112 10.6151
R879 B.n113 B.n86 10.6151
R880 B.n117 B.n86 10.6151
R881 B.n118 B.n117 10.6151
R882 B.n119 B.n118 10.6151
R883 B.n119 B.n84 10.6151
R884 B.n124 B.n123 10.6151
R885 B.n125 B.n124 10.6151
R886 B.n125 B.n82 10.6151
R887 B.n129 B.n82 10.6151
R888 B.n130 B.n129 10.6151
R889 B.n131 B.n130 10.6151
R890 B.n131 B.n80 10.6151
R891 B.n135 B.n80 10.6151
R892 B.n136 B.n135 10.6151
R893 B.n137 B.n136 10.6151
R894 B.n137 B.n78 10.6151
R895 B.n141 B.n78 10.6151
R896 B.n142 B.n141 10.6151
R897 B.n143 B.n142 10.6151
R898 B.n143 B.n76 10.6151
R899 B.n147 B.n76 10.6151
R900 B.n148 B.n147 10.6151
R901 B.n150 B.n72 10.6151
R902 B.n154 B.n72 10.6151
R903 B.n155 B.n154 10.6151
R904 B.n156 B.n155 10.6151
R905 B.n156 B.n70 10.6151
R906 B.n160 B.n70 10.6151
R907 B.n161 B.n160 10.6151
R908 B.n165 B.n161 10.6151
R909 B.n169 B.n68 10.6151
R910 B.n170 B.n169 10.6151
R911 B.n171 B.n170 10.6151
R912 B.n171 B.n66 10.6151
R913 B.n175 B.n66 10.6151
R914 B.n176 B.n175 10.6151
R915 B.n177 B.n176 10.6151
R916 B.n177 B.n64 10.6151
R917 B.n181 B.n64 10.6151
R918 B.n182 B.n181 10.6151
R919 B.n183 B.n182 10.6151
R920 B.n183 B.n62 10.6151
R921 B.n187 B.n62 10.6151
R922 B.n188 B.n187 10.6151
R923 B.n189 B.n188 10.6151
R924 B.n189 B.n60 10.6151
R925 B.n193 B.n60 10.6151
R926 B.n357 B.n0 8.11757
R927 B.n357 B.n1 8.11757
R928 B.n298 B.n297 6.5566
R929 B.n285 B.n284 6.5566
R930 B.n150 B.n149 6.5566
R931 B.n165 B.n164 6.5566
R932 B.n299 B.n298 4.05904
R933 B.n284 B.n283 4.05904
R934 B.n149 B.n148 4.05904
R935 B.n164 B.n68 4.05904
C0 VN B 0.620706f
C1 VTAIL VP 1.83097f
C2 VDD1 VDD2 0.765806f
C3 VTAIL VN 1.81666f
C4 B w_n1810_n1758# 4.54014f
C5 VN VP 3.62877f
C6 VTAIL w_n1810_n1758# 1.71585f
C7 VDD2 B 1.01848f
C8 VDD1 B 0.986775f
C9 w_n1810_n1758# VP 3.26548f
C10 VN w_n1810_n1758# 3.03766f
C11 VTAIL VDD2 7.74377f
C12 VTAIL VDD1 7.70779f
C13 VDD2 VP 0.302975f
C14 VDD1 VP 1.91869f
C15 VN VDD2 1.77059f
C16 VN VDD1 0.152613f
C17 VTAIL B 1.15246f
C18 B VP 0.99289f
C19 VDD2 w_n1810_n1758# 1.31153f
C20 VDD1 w_n1810_n1758# 1.28424f
C21 VDD2 VSUBS 0.889577f
C22 VDD1 VSUBS 0.762555f
C23 VTAIL VSUBS 0.317774f
C24 VN VSUBS 3.15238f
C25 VP VSUBS 1.004208f
C26 B VSUBS 1.830802f
C27 w_n1810_n1758# VSUBS 40.0734f
C28 B.n0 VSUBS 0.006527f
C29 B.n1 VSUBS 0.006527f
C30 B.n2 VSUBS 0.009653f
C31 B.n3 VSUBS 0.007397f
C32 B.n4 VSUBS 0.007397f
C33 B.n5 VSUBS 0.007397f
C34 B.n6 VSUBS 0.007397f
C35 B.n7 VSUBS 0.007397f
C36 B.n8 VSUBS 0.007397f
C37 B.n9 VSUBS 0.007397f
C38 B.n10 VSUBS 0.007397f
C39 B.n11 VSUBS 0.007397f
C40 B.n12 VSUBS 0.018161f
C41 B.n13 VSUBS 0.007397f
C42 B.n14 VSUBS 0.007397f
C43 B.n15 VSUBS 0.007397f
C44 B.n16 VSUBS 0.007397f
C45 B.n17 VSUBS 0.007397f
C46 B.n18 VSUBS 0.007397f
C47 B.n19 VSUBS 0.007397f
C48 B.n20 VSUBS 0.007397f
C49 B.n21 VSUBS 0.007397f
C50 B.t4 VSUBS 0.060458f
C51 B.t5 VSUBS 0.06597f
C52 B.t3 VSUBS 0.065974f
C53 B.n22 VSUBS 0.118759f
C54 B.n23 VSUBS 0.111335f
C55 B.n24 VSUBS 0.007397f
C56 B.n25 VSUBS 0.007397f
C57 B.n26 VSUBS 0.007397f
C58 B.n27 VSUBS 0.007397f
C59 B.t1 VSUBS 0.060459f
C60 B.t2 VSUBS 0.065971f
C61 B.t0 VSUBS 0.065974f
C62 B.n28 VSUBS 0.118758f
C63 B.n29 VSUBS 0.111334f
C64 B.n30 VSUBS 0.007397f
C65 B.n31 VSUBS 0.007397f
C66 B.n32 VSUBS 0.007397f
C67 B.n33 VSUBS 0.007397f
C68 B.n34 VSUBS 0.007397f
C69 B.n35 VSUBS 0.007397f
C70 B.n36 VSUBS 0.007397f
C71 B.n37 VSUBS 0.007397f
C72 B.n38 VSUBS 0.018161f
C73 B.n39 VSUBS 0.007397f
C74 B.n40 VSUBS 0.007397f
C75 B.n41 VSUBS 0.007397f
C76 B.n42 VSUBS 0.007397f
C77 B.n43 VSUBS 0.007397f
C78 B.n44 VSUBS 0.007397f
C79 B.n45 VSUBS 0.007397f
C80 B.n46 VSUBS 0.007397f
C81 B.n47 VSUBS 0.007397f
C82 B.n48 VSUBS 0.007397f
C83 B.n49 VSUBS 0.007397f
C84 B.n50 VSUBS 0.007397f
C85 B.n51 VSUBS 0.007397f
C86 B.n52 VSUBS 0.007397f
C87 B.n53 VSUBS 0.007397f
C88 B.n54 VSUBS 0.007397f
C89 B.n55 VSUBS 0.007397f
C90 B.n56 VSUBS 0.007397f
C91 B.n57 VSUBS 0.007397f
C92 B.n58 VSUBS 0.007397f
C93 B.n59 VSUBS 0.017737f
C94 B.n60 VSUBS 0.007397f
C95 B.n61 VSUBS 0.007397f
C96 B.n62 VSUBS 0.007397f
C97 B.n63 VSUBS 0.007397f
C98 B.n64 VSUBS 0.007397f
C99 B.n65 VSUBS 0.007397f
C100 B.n66 VSUBS 0.007397f
C101 B.n67 VSUBS 0.007397f
C102 B.n68 VSUBS 0.005113f
C103 B.n69 VSUBS 0.007397f
C104 B.n70 VSUBS 0.007397f
C105 B.n71 VSUBS 0.007397f
C106 B.n72 VSUBS 0.007397f
C107 B.n73 VSUBS 0.007397f
C108 B.t11 VSUBS 0.060458f
C109 B.t10 VSUBS 0.06597f
C110 B.t9 VSUBS 0.065974f
C111 B.n74 VSUBS 0.118759f
C112 B.n75 VSUBS 0.111335f
C113 B.n76 VSUBS 0.007397f
C114 B.n77 VSUBS 0.007397f
C115 B.n78 VSUBS 0.007397f
C116 B.n79 VSUBS 0.007397f
C117 B.n80 VSUBS 0.007397f
C118 B.n81 VSUBS 0.007397f
C119 B.n82 VSUBS 0.007397f
C120 B.n83 VSUBS 0.007397f
C121 B.n84 VSUBS 0.017737f
C122 B.n85 VSUBS 0.007397f
C123 B.n86 VSUBS 0.007397f
C124 B.n87 VSUBS 0.007397f
C125 B.n88 VSUBS 0.007397f
C126 B.n89 VSUBS 0.007397f
C127 B.n90 VSUBS 0.007397f
C128 B.n91 VSUBS 0.007397f
C129 B.n92 VSUBS 0.007397f
C130 B.n93 VSUBS 0.007397f
C131 B.n94 VSUBS 0.007397f
C132 B.n95 VSUBS 0.007397f
C133 B.n96 VSUBS 0.007397f
C134 B.n97 VSUBS 0.007397f
C135 B.n98 VSUBS 0.007397f
C136 B.n99 VSUBS 0.007397f
C137 B.n100 VSUBS 0.007397f
C138 B.n101 VSUBS 0.007397f
C139 B.n102 VSUBS 0.007397f
C140 B.n103 VSUBS 0.007397f
C141 B.n104 VSUBS 0.007397f
C142 B.n105 VSUBS 0.007397f
C143 B.n106 VSUBS 0.007397f
C144 B.n107 VSUBS 0.007397f
C145 B.n108 VSUBS 0.007397f
C146 B.n109 VSUBS 0.007397f
C147 B.n110 VSUBS 0.007397f
C148 B.n111 VSUBS 0.007397f
C149 B.n112 VSUBS 0.007397f
C150 B.n113 VSUBS 0.007397f
C151 B.n114 VSUBS 0.007397f
C152 B.n115 VSUBS 0.007397f
C153 B.n116 VSUBS 0.007397f
C154 B.n117 VSUBS 0.007397f
C155 B.n118 VSUBS 0.007397f
C156 B.n119 VSUBS 0.007397f
C157 B.n120 VSUBS 0.007397f
C158 B.n121 VSUBS 0.017737f
C159 B.n122 VSUBS 0.018161f
C160 B.n123 VSUBS 0.018161f
C161 B.n124 VSUBS 0.007397f
C162 B.n125 VSUBS 0.007397f
C163 B.n126 VSUBS 0.007397f
C164 B.n127 VSUBS 0.007397f
C165 B.n128 VSUBS 0.007397f
C166 B.n129 VSUBS 0.007397f
C167 B.n130 VSUBS 0.007397f
C168 B.n131 VSUBS 0.007397f
C169 B.n132 VSUBS 0.007397f
C170 B.n133 VSUBS 0.007397f
C171 B.n134 VSUBS 0.007397f
C172 B.n135 VSUBS 0.007397f
C173 B.n136 VSUBS 0.007397f
C174 B.n137 VSUBS 0.007397f
C175 B.n138 VSUBS 0.007397f
C176 B.n139 VSUBS 0.007397f
C177 B.n140 VSUBS 0.007397f
C178 B.n141 VSUBS 0.007397f
C179 B.n142 VSUBS 0.007397f
C180 B.n143 VSUBS 0.007397f
C181 B.n144 VSUBS 0.007397f
C182 B.n145 VSUBS 0.007397f
C183 B.n146 VSUBS 0.007397f
C184 B.n147 VSUBS 0.007397f
C185 B.n148 VSUBS 0.005113f
C186 B.n149 VSUBS 0.017138f
C187 B.n150 VSUBS 0.005983f
C188 B.n151 VSUBS 0.007397f
C189 B.n152 VSUBS 0.007397f
C190 B.n153 VSUBS 0.007397f
C191 B.n154 VSUBS 0.007397f
C192 B.n155 VSUBS 0.007397f
C193 B.n156 VSUBS 0.007397f
C194 B.n157 VSUBS 0.007397f
C195 B.n158 VSUBS 0.007397f
C196 B.n159 VSUBS 0.007397f
C197 B.n160 VSUBS 0.007397f
C198 B.n161 VSUBS 0.007397f
C199 B.t8 VSUBS 0.060459f
C200 B.t7 VSUBS 0.065971f
C201 B.t6 VSUBS 0.065974f
C202 B.n162 VSUBS 0.118758f
C203 B.n163 VSUBS 0.111334f
C204 B.n164 VSUBS 0.017138f
C205 B.n165 VSUBS 0.005983f
C206 B.n166 VSUBS 0.007397f
C207 B.n167 VSUBS 0.007397f
C208 B.n168 VSUBS 0.007397f
C209 B.n169 VSUBS 0.007397f
C210 B.n170 VSUBS 0.007397f
C211 B.n171 VSUBS 0.007397f
C212 B.n172 VSUBS 0.007397f
C213 B.n173 VSUBS 0.007397f
C214 B.n174 VSUBS 0.007397f
C215 B.n175 VSUBS 0.007397f
C216 B.n176 VSUBS 0.007397f
C217 B.n177 VSUBS 0.007397f
C218 B.n178 VSUBS 0.007397f
C219 B.n179 VSUBS 0.007397f
C220 B.n180 VSUBS 0.007397f
C221 B.n181 VSUBS 0.007397f
C222 B.n182 VSUBS 0.007397f
C223 B.n183 VSUBS 0.007397f
C224 B.n184 VSUBS 0.007397f
C225 B.n185 VSUBS 0.007397f
C226 B.n186 VSUBS 0.007397f
C227 B.n187 VSUBS 0.007397f
C228 B.n188 VSUBS 0.007397f
C229 B.n189 VSUBS 0.007397f
C230 B.n190 VSUBS 0.007397f
C231 B.n191 VSUBS 0.007397f
C232 B.n192 VSUBS 0.018161f
C233 B.n193 VSUBS 0.017333f
C234 B.n194 VSUBS 0.018564f
C235 B.n195 VSUBS 0.007397f
C236 B.n196 VSUBS 0.007397f
C237 B.n197 VSUBS 0.007397f
C238 B.n198 VSUBS 0.007397f
C239 B.n199 VSUBS 0.007397f
C240 B.n200 VSUBS 0.007397f
C241 B.n201 VSUBS 0.007397f
C242 B.n202 VSUBS 0.007397f
C243 B.n203 VSUBS 0.007397f
C244 B.n204 VSUBS 0.007397f
C245 B.n205 VSUBS 0.007397f
C246 B.n206 VSUBS 0.007397f
C247 B.n207 VSUBS 0.007397f
C248 B.n208 VSUBS 0.007397f
C249 B.n209 VSUBS 0.007397f
C250 B.n210 VSUBS 0.007397f
C251 B.n211 VSUBS 0.007397f
C252 B.n212 VSUBS 0.007397f
C253 B.n213 VSUBS 0.007397f
C254 B.n214 VSUBS 0.007397f
C255 B.n215 VSUBS 0.007397f
C256 B.n216 VSUBS 0.007397f
C257 B.n217 VSUBS 0.007397f
C258 B.n218 VSUBS 0.007397f
C259 B.n219 VSUBS 0.007397f
C260 B.n220 VSUBS 0.007397f
C261 B.n221 VSUBS 0.007397f
C262 B.n222 VSUBS 0.007397f
C263 B.n223 VSUBS 0.007397f
C264 B.n224 VSUBS 0.007397f
C265 B.n225 VSUBS 0.007397f
C266 B.n226 VSUBS 0.007397f
C267 B.n227 VSUBS 0.007397f
C268 B.n228 VSUBS 0.007397f
C269 B.n229 VSUBS 0.007397f
C270 B.n230 VSUBS 0.007397f
C271 B.n231 VSUBS 0.007397f
C272 B.n232 VSUBS 0.007397f
C273 B.n233 VSUBS 0.007397f
C274 B.n234 VSUBS 0.007397f
C275 B.n235 VSUBS 0.007397f
C276 B.n236 VSUBS 0.007397f
C277 B.n237 VSUBS 0.007397f
C278 B.n238 VSUBS 0.007397f
C279 B.n239 VSUBS 0.007397f
C280 B.n240 VSUBS 0.007397f
C281 B.n241 VSUBS 0.007397f
C282 B.n242 VSUBS 0.007397f
C283 B.n243 VSUBS 0.007397f
C284 B.n244 VSUBS 0.007397f
C285 B.n245 VSUBS 0.007397f
C286 B.n246 VSUBS 0.007397f
C287 B.n247 VSUBS 0.007397f
C288 B.n248 VSUBS 0.007397f
C289 B.n249 VSUBS 0.007397f
C290 B.n250 VSUBS 0.007397f
C291 B.n251 VSUBS 0.007397f
C292 B.n252 VSUBS 0.007397f
C293 B.n253 VSUBS 0.007397f
C294 B.n254 VSUBS 0.007397f
C295 B.n255 VSUBS 0.017737f
C296 B.n256 VSUBS 0.017737f
C297 B.n257 VSUBS 0.018161f
C298 B.n258 VSUBS 0.007397f
C299 B.n259 VSUBS 0.007397f
C300 B.n260 VSUBS 0.007397f
C301 B.n261 VSUBS 0.007397f
C302 B.n262 VSUBS 0.007397f
C303 B.n263 VSUBS 0.007397f
C304 B.n264 VSUBS 0.007397f
C305 B.n265 VSUBS 0.007397f
C306 B.n266 VSUBS 0.007397f
C307 B.n267 VSUBS 0.007397f
C308 B.n268 VSUBS 0.007397f
C309 B.n269 VSUBS 0.007397f
C310 B.n270 VSUBS 0.007397f
C311 B.n271 VSUBS 0.007397f
C312 B.n272 VSUBS 0.007397f
C313 B.n273 VSUBS 0.007397f
C314 B.n274 VSUBS 0.007397f
C315 B.n275 VSUBS 0.007397f
C316 B.n276 VSUBS 0.007397f
C317 B.n277 VSUBS 0.007397f
C318 B.n278 VSUBS 0.007397f
C319 B.n279 VSUBS 0.007397f
C320 B.n280 VSUBS 0.007397f
C321 B.n281 VSUBS 0.007397f
C322 B.n282 VSUBS 0.007397f
C323 B.n283 VSUBS 0.005113f
C324 B.n284 VSUBS 0.017138f
C325 B.n285 VSUBS 0.005983f
C326 B.n286 VSUBS 0.007397f
C327 B.n287 VSUBS 0.007397f
C328 B.n288 VSUBS 0.007397f
C329 B.n289 VSUBS 0.007397f
C330 B.n290 VSUBS 0.007397f
C331 B.n291 VSUBS 0.007397f
C332 B.n292 VSUBS 0.007397f
C333 B.n293 VSUBS 0.007397f
C334 B.n294 VSUBS 0.007397f
C335 B.n295 VSUBS 0.007397f
C336 B.n296 VSUBS 0.007397f
C337 B.n297 VSUBS 0.005983f
C338 B.n298 VSUBS 0.017138f
C339 B.n299 VSUBS 0.005113f
C340 B.n300 VSUBS 0.007397f
C341 B.n301 VSUBS 0.007397f
C342 B.n302 VSUBS 0.007397f
C343 B.n303 VSUBS 0.007397f
C344 B.n304 VSUBS 0.007397f
C345 B.n305 VSUBS 0.007397f
C346 B.n306 VSUBS 0.007397f
C347 B.n307 VSUBS 0.007397f
C348 B.n308 VSUBS 0.007397f
C349 B.n309 VSUBS 0.007397f
C350 B.n310 VSUBS 0.007397f
C351 B.n311 VSUBS 0.007397f
C352 B.n312 VSUBS 0.007397f
C353 B.n313 VSUBS 0.007397f
C354 B.n314 VSUBS 0.007397f
C355 B.n315 VSUBS 0.007397f
C356 B.n316 VSUBS 0.007397f
C357 B.n317 VSUBS 0.007397f
C358 B.n318 VSUBS 0.007397f
C359 B.n319 VSUBS 0.007397f
C360 B.n320 VSUBS 0.007397f
C361 B.n321 VSUBS 0.007397f
C362 B.n322 VSUBS 0.007397f
C363 B.n323 VSUBS 0.007397f
C364 B.n324 VSUBS 0.007397f
C365 B.n325 VSUBS 0.018161f
C366 B.n326 VSUBS 0.017737f
C367 B.n327 VSUBS 0.017737f
C368 B.n328 VSUBS 0.007397f
C369 B.n329 VSUBS 0.007397f
C370 B.n330 VSUBS 0.007397f
C371 B.n331 VSUBS 0.007397f
C372 B.n332 VSUBS 0.007397f
C373 B.n333 VSUBS 0.007397f
C374 B.n334 VSUBS 0.007397f
C375 B.n335 VSUBS 0.007397f
C376 B.n336 VSUBS 0.007397f
C377 B.n337 VSUBS 0.007397f
C378 B.n338 VSUBS 0.007397f
C379 B.n339 VSUBS 0.007397f
C380 B.n340 VSUBS 0.007397f
C381 B.n341 VSUBS 0.007397f
C382 B.n342 VSUBS 0.007397f
C383 B.n343 VSUBS 0.007397f
C384 B.n344 VSUBS 0.007397f
C385 B.n345 VSUBS 0.007397f
C386 B.n346 VSUBS 0.007397f
C387 B.n347 VSUBS 0.007397f
C388 B.n348 VSUBS 0.007397f
C389 B.n349 VSUBS 0.007397f
C390 B.n350 VSUBS 0.007397f
C391 B.n351 VSUBS 0.007397f
C392 B.n352 VSUBS 0.007397f
C393 B.n353 VSUBS 0.007397f
C394 B.n354 VSUBS 0.007397f
C395 B.n355 VSUBS 0.009653f
C396 B.n356 VSUBS 0.010283f
C397 B.n357 VSUBS 0.020448f
C398 VDD2.n0 VSUBS 0.024392f
C399 VDD2.n1 VSUBS 0.02237f
C400 VDD2.n2 VSUBS 0.012021f
C401 VDD2.n3 VSUBS 0.028413f
C402 VDD2.n4 VSUBS 0.012728f
C403 VDD2.n5 VSUBS 0.086761f
C404 VDD2.t4 VSUBS 0.062868f
C405 VDD2.n6 VSUBS 0.021309f
C406 VDD2.n7 VSUBS 0.017871f
C407 VDD2.n8 VSUBS 0.012021f
C408 VDD2.n9 VSUBS 0.301769f
C409 VDD2.n10 VSUBS 0.02237f
C410 VDD2.n11 VSUBS 0.012021f
C411 VDD2.n12 VSUBS 0.012728f
C412 VDD2.n13 VSUBS 0.028413f
C413 VDD2.n14 VSUBS 0.068142f
C414 VDD2.n15 VSUBS 0.012728f
C415 VDD2.n16 VSUBS 0.012021f
C416 VDD2.n17 VSUBS 0.055069f
C417 VDD2.n18 VSUBS 0.050796f
C418 VDD2.t5 VSUBS 0.069826f
C419 VDD2.t6 VSUBS 0.069826f
C420 VDD2.n19 VSUBS 0.4065f
C421 VDD2.n20 VSUBS 0.458105f
C422 VDD2.t0 VSUBS 0.069826f
C423 VDD2.t2 VSUBS 0.069826f
C424 VDD2.n21 VSUBS 0.407859f
C425 VDD2.n22 VSUBS 1.25251f
C426 VDD2.n23 VSUBS 0.024392f
C427 VDD2.n24 VSUBS 0.02237f
C428 VDD2.n25 VSUBS 0.012021f
C429 VDD2.n26 VSUBS 0.028413f
C430 VDD2.n27 VSUBS 0.012728f
C431 VDD2.n28 VSUBS 0.086761f
C432 VDD2.t3 VSUBS 0.062868f
C433 VDD2.n29 VSUBS 0.021309f
C434 VDD2.n30 VSUBS 0.017871f
C435 VDD2.n31 VSUBS 0.012021f
C436 VDD2.n32 VSUBS 0.301769f
C437 VDD2.n33 VSUBS 0.02237f
C438 VDD2.n34 VSUBS 0.012021f
C439 VDD2.n35 VSUBS 0.012728f
C440 VDD2.n36 VSUBS 0.028413f
C441 VDD2.n37 VSUBS 0.068142f
C442 VDD2.n38 VSUBS 0.012728f
C443 VDD2.n39 VSUBS 0.012021f
C444 VDD2.n40 VSUBS 0.055069f
C445 VDD2.n41 VSUBS 0.049761f
C446 VDD2.n42 VSUBS 1.23817f
C447 VDD2.t1 VSUBS 0.069826f
C448 VDD2.t9 VSUBS 0.069826f
C449 VDD2.n43 VSUBS 0.406502f
C450 VDD2.n44 VSUBS 0.373394f
C451 VDD2.t8 VSUBS 0.069826f
C452 VDD2.t7 VSUBS 0.069826f
C453 VDD2.n45 VSUBS 0.407845f
C454 VN.n0 VSUBS 0.047091f
C455 VN.t3 VSUBS 0.203293f
C456 VN.n1 VSUBS 0.105502f
C457 VN.t5 VSUBS 0.209421f
C458 VN.n2 VSUBS 0.106613f
C459 VN.t4 VSUBS 0.203293f
C460 VN.n3 VSUBS 0.120108f
C461 VN.n4 VSUBS 0.010686f
C462 VN.n5 VSUBS 0.145881f
C463 VN.n6 VSUBS 0.047091f
C464 VN.n7 VSUBS 0.010686f
C465 VN.t9 VSUBS 0.203293f
C466 VN.n8 VSUBS 0.120108f
C467 VN.t7 VSUBS 0.203293f
C468 VN.n9 VSUBS 0.112414f
C469 VN.n10 VSUBS 0.036494f
C470 VN.n11 VSUBS 0.047091f
C471 VN.t0 VSUBS 0.203293f
C472 VN.n12 VSUBS 0.105502f
C473 VN.t2 VSUBS 0.209421f
C474 VN.n13 VSUBS 0.106613f
C475 VN.t1 VSUBS 0.203293f
C476 VN.n14 VSUBS 0.120108f
C477 VN.n15 VSUBS 0.010686f
C478 VN.n16 VSUBS 0.145881f
C479 VN.n17 VSUBS 0.047091f
C480 VN.n18 VSUBS 0.010686f
C481 VN.t8 VSUBS 0.203293f
C482 VN.n19 VSUBS 0.120108f
C483 VN.t6 VSUBS 0.203293f
C484 VN.n20 VSUBS 0.112414f
C485 VN.n21 VSUBS 1.42517f
C486 VTAIL.t15 VSUBS 0.079379f
C487 VTAIL.t18 VSUBS 0.079379f
C488 VTAIL.n0 VSUBS 0.402644f
C489 VTAIL.n1 VSUBS 0.487879f
C490 VTAIL.n2 VSUBS 0.027728f
C491 VTAIL.n3 VSUBS 0.025431f
C492 VTAIL.n4 VSUBS 0.013665f
C493 VTAIL.n5 VSUBS 0.0323f
C494 VTAIL.n6 VSUBS 0.014469f
C495 VTAIL.n7 VSUBS 0.098631f
C496 VTAIL.t2 VSUBS 0.071468f
C497 VTAIL.n8 VSUBS 0.024225f
C498 VTAIL.n9 VSUBS 0.020316f
C499 VTAIL.n10 VSUBS 0.013665f
C500 VTAIL.n11 VSUBS 0.343052f
C501 VTAIL.n12 VSUBS 0.025431f
C502 VTAIL.n13 VSUBS 0.013665f
C503 VTAIL.n14 VSUBS 0.014469f
C504 VTAIL.n15 VSUBS 0.0323f
C505 VTAIL.n16 VSUBS 0.077464f
C506 VTAIL.n17 VSUBS 0.014469f
C507 VTAIL.n18 VSUBS 0.013665f
C508 VTAIL.n19 VSUBS 0.062603f
C509 VTAIL.n20 VSUBS 0.039038f
C510 VTAIL.n21 VSUBS 0.136551f
C511 VTAIL.t10 VSUBS 0.079379f
C512 VTAIL.t4 VSUBS 0.079379f
C513 VTAIL.n22 VSUBS 0.402644f
C514 VTAIL.n23 VSUBS 0.481698f
C515 VTAIL.t8 VSUBS 0.079379f
C516 VTAIL.t11 VSUBS 0.079379f
C517 VTAIL.n24 VSUBS 0.402644f
C518 VTAIL.n25 VSUBS 1.15562f
C519 VTAIL.t14 VSUBS 0.079379f
C520 VTAIL.t19 VSUBS 0.079379f
C521 VTAIL.n26 VSUBS 0.402646f
C522 VTAIL.n27 VSUBS 1.15562f
C523 VTAIL.t1 VSUBS 0.079379f
C524 VTAIL.t0 VSUBS 0.079379f
C525 VTAIL.n28 VSUBS 0.402646f
C526 VTAIL.n29 VSUBS 0.481696f
C527 VTAIL.n30 VSUBS 0.027728f
C528 VTAIL.n31 VSUBS 0.025431f
C529 VTAIL.n32 VSUBS 0.013665f
C530 VTAIL.n33 VSUBS 0.0323f
C531 VTAIL.n34 VSUBS 0.014469f
C532 VTAIL.n35 VSUBS 0.098631f
C533 VTAIL.t16 VSUBS 0.071468f
C534 VTAIL.n36 VSUBS 0.024225f
C535 VTAIL.n37 VSUBS 0.020316f
C536 VTAIL.n38 VSUBS 0.013665f
C537 VTAIL.n39 VSUBS 0.343052f
C538 VTAIL.n40 VSUBS 0.025431f
C539 VTAIL.n41 VSUBS 0.013665f
C540 VTAIL.n42 VSUBS 0.014469f
C541 VTAIL.n43 VSUBS 0.0323f
C542 VTAIL.n44 VSUBS 0.077464f
C543 VTAIL.n45 VSUBS 0.014469f
C544 VTAIL.n46 VSUBS 0.013665f
C545 VTAIL.n47 VSUBS 0.062603f
C546 VTAIL.n48 VSUBS 0.039038f
C547 VTAIL.n49 VSUBS 0.136551f
C548 VTAIL.t6 VSUBS 0.079379f
C549 VTAIL.t9 VSUBS 0.079379f
C550 VTAIL.n50 VSUBS 0.402646f
C551 VTAIL.n51 VSUBS 0.495471f
C552 VTAIL.t3 VSUBS 0.079379f
C553 VTAIL.t5 VSUBS 0.079379f
C554 VTAIL.n52 VSUBS 0.402646f
C555 VTAIL.n53 VSUBS 0.481696f
C556 VTAIL.n54 VSUBS 0.027728f
C557 VTAIL.n55 VSUBS 0.025431f
C558 VTAIL.n56 VSUBS 0.013665f
C559 VTAIL.n57 VSUBS 0.0323f
C560 VTAIL.n58 VSUBS 0.014469f
C561 VTAIL.n59 VSUBS 0.098631f
C562 VTAIL.t7 VSUBS 0.071468f
C563 VTAIL.n60 VSUBS 0.024225f
C564 VTAIL.n61 VSUBS 0.020316f
C565 VTAIL.n62 VSUBS 0.013665f
C566 VTAIL.n63 VSUBS 0.343052f
C567 VTAIL.n64 VSUBS 0.025431f
C568 VTAIL.n65 VSUBS 0.013665f
C569 VTAIL.n66 VSUBS 0.014469f
C570 VTAIL.n67 VSUBS 0.0323f
C571 VTAIL.n68 VSUBS 0.077464f
C572 VTAIL.n69 VSUBS 0.014469f
C573 VTAIL.n70 VSUBS 0.013665f
C574 VTAIL.n71 VSUBS 0.062603f
C575 VTAIL.n72 VSUBS 0.039038f
C576 VTAIL.n73 VSUBS 0.747247f
C577 VTAIL.n74 VSUBS 0.027728f
C578 VTAIL.n75 VSUBS 0.025431f
C579 VTAIL.n76 VSUBS 0.013665f
C580 VTAIL.n77 VSUBS 0.0323f
C581 VTAIL.n78 VSUBS 0.014469f
C582 VTAIL.n79 VSUBS 0.098631f
C583 VTAIL.t13 VSUBS 0.071468f
C584 VTAIL.n80 VSUBS 0.024225f
C585 VTAIL.n81 VSUBS 0.020316f
C586 VTAIL.n82 VSUBS 0.013665f
C587 VTAIL.n83 VSUBS 0.343052f
C588 VTAIL.n84 VSUBS 0.025431f
C589 VTAIL.n85 VSUBS 0.013665f
C590 VTAIL.n86 VSUBS 0.014469f
C591 VTAIL.n87 VSUBS 0.0323f
C592 VTAIL.n88 VSUBS 0.077464f
C593 VTAIL.n89 VSUBS 0.014469f
C594 VTAIL.n90 VSUBS 0.013665f
C595 VTAIL.n91 VSUBS 0.062603f
C596 VTAIL.n92 VSUBS 0.039038f
C597 VTAIL.n93 VSUBS 0.747247f
C598 VTAIL.t12 VSUBS 0.079379f
C599 VTAIL.t17 VSUBS 0.079379f
C600 VTAIL.n94 VSUBS 0.402644f
C601 VTAIL.n95 VSUBS 0.439844f
C602 VDD1.n0 VSUBS 0.024133f
C603 VDD1.n1 VSUBS 0.022133f
C604 VDD1.n2 VSUBS 0.011893f
C605 VDD1.n3 VSUBS 0.028111f
C606 VDD1.n4 VSUBS 0.012593f
C607 VDD1.n5 VSUBS 0.08584f
C608 VDD1.t2 VSUBS 0.0622f
C609 VDD1.n6 VSUBS 0.021083f
C610 VDD1.n7 VSUBS 0.017681f
C611 VDD1.n8 VSUBS 0.011893f
C612 VDD1.n9 VSUBS 0.298565f
C613 VDD1.n10 VSUBS 0.022133f
C614 VDD1.n11 VSUBS 0.011893f
C615 VDD1.n12 VSUBS 0.012593f
C616 VDD1.n13 VSUBS 0.028111f
C617 VDD1.n14 VSUBS 0.067419f
C618 VDD1.n15 VSUBS 0.012593f
C619 VDD1.n16 VSUBS 0.011893f
C620 VDD1.n17 VSUBS 0.054484f
C621 VDD1.n18 VSUBS 0.050257f
C622 VDD1.t1 VSUBS 0.069085f
C623 VDD1.t3 VSUBS 0.069085f
C624 VDD1.n19 VSUBS 0.402186f
C625 VDD1.n20 VSUBS 0.455964f
C626 VDD1.n21 VSUBS 0.024133f
C627 VDD1.n22 VSUBS 0.022133f
C628 VDD1.n23 VSUBS 0.011893f
C629 VDD1.n24 VSUBS 0.028111f
C630 VDD1.n25 VSUBS 0.012593f
C631 VDD1.n26 VSUBS 0.08584f
C632 VDD1.t9 VSUBS 0.0622f
C633 VDD1.n27 VSUBS 0.021083f
C634 VDD1.n28 VSUBS 0.017681f
C635 VDD1.n29 VSUBS 0.011893f
C636 VDD1.n30 VSUBS 0.298565f
C637 VDD1.n31 VSUBS 0.022133f
C638 VDD1.n32 VSUBS 0.011893f
C639 VDD1.n33 VSUBS 0.012593f
C640 VDD1.n34 VSUBS 0.028111f
C641 VDD1.n35 VSUBS 0.067419f
C642 VDD1.n36 VSUBS 0.012593f
C643 VDD1.n37 VSUBS 0.011893f
C644 VDD1.n38 VSUBS 0.054484f
C645 VDD1.n39 VSUBS 0.050257f
C646 VDD1.t8 VSUBS 0.069085f
C647 VDD1.t6 VSUBS 0.069085f
C648 VDD1.n40 VSUBS 0.402185f
C649 VDD1.n41 VSUBS 0.453241f
C650 VDD1.t5 VSUBS 0.069085f
C651 VDD1.t0 VSUBS 0.069085f
C652 VDD1.n42 VSUBS 0.403529f
C653 VDD1.n43 VSUBS 1.29838f
C654 VDD1.t4 VSUBS 0.069085f
C655 VDD1.t7 VSUBS 0.069085f
C656 VDD1.n44 VSUBS 0.402185f
C657 VDD1.n45 VSUBS 1.55161f
C658 VP.n0 VSUBS 0.04973f
C659 VP.t1 VSUBS 0.214687f
C660 VP.n1 VSUBS 0.111415f
C661 VP.n2 VSUBS 0.04973f
C662 VP.n3 VSUBS 0.04973f
C663 VP.t4 VSUBS 0.214687f
C664 VP.t6 VSUBS 0.214687f
C665 VP.t8 VSUBS 0.214687f
C666 VP.n4 VSUBS 0.111415f
C667 VP.t5 VSUBS 0.221158f
C668 VP.n5 VSUBS 0.112588f
C669 VP.t2 VSUBS 0.214687f
C670 VP.n6 VSUBS 0.126839f
C671 VP.n7 VSUBS 0.011285f
C672 VP.n8 VSUBS 0.154057f
C673 VP.n9 VSUBS 0.04973f
C674 VP.n10 VSUBS 0.011285f
C675 VP.n11 VSUBS 0.126839f
C676 VP.n12 VSUBS 0.118714f
C677 VP.n13 VSUBS 1.47199f
C678 VP.n14 VSUBS 1.52324f
C679 VP.t3 VSUBS 0.214687f
C680 VP.n15 VSUBS 0.118714f
C681 VP.t0 VSUBS 0.214687f
C682 VP.n16 VSUBS 0.126839f
C683 VP.n17 VSUBS 0.011285f
C684 VP.n18 VSUBS 0.04973f
C685 VP.n19 VSUBS 0.04973f
C686 VP.n20 VSUBS 0.011285f
C687 VP.t7 VSUBS 0.214687f
C688 VP.n21 VSUBS 0.126839f
C689 VP.t9 VSUBS 0.214687f
C690 VP.n22 VSUBS 0.118714f
C691 VP.n23 VSUBS 0.038539f
.ends

