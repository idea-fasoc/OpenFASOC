* NGSPICE file created from diff_pair_sample_0138.ext - technology: sky130A

.subckt diff_pair_sample_0138 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=0 ps=0 w=17.09 l=2.74
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=6.6651 ps=34.96 w=17.09 l=2.74
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=6.6651 ps=34.96 w=17.09 l=2.74
X3 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=6.6651 ps=34.96 w=17.09 l=2.74
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=0 ps=0 w=17.09 l=2.74
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=0 ps=0 w=17.09 l=2.74
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=6.6651 ps=34.96 w=17.09 l=2.74
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6651 pd=34.96 as=0 ps=0 w=17.09 l=2.74
R0 B.n592 B.n117 585
R1 B.n117 B.n50 585
R2 B.n594 B.n593 585
R3 B.n596 B.n116 585
R4 B.n599 B.n598 585
R5 B.n600 B.n115 585
R6 B.n602 B.n601 585
R7 B.n604 B.n114 585
R8 B.n607 B.n606 585
R9 B.n608 B.n113 585
R10 B.n610 B.n609 585
R11 B.n612 B.n112 585
R12 B.n615 B.n614 585
R13 B.n616 B.n111 585
R14 B.n618 B.n617 585
R15 B.n620 B.n110 585
R16 B.n623 B.n622 585
R17 B.n624 B.n109 585
R18 B.n626 B.n625 585
R19 B.n628 B.n108 585
R20 B.n631 B.n630 585
R21 B.n632 B.n107 585
R22 B.n634 B.n633 585
R23 B.n636 B.n106 585
R24 B.n639 B.n638 585
R25 B.n640 B.n105 585
R26 B.n642 B.n641 585
R27 B.n644 B.n104 585
R28 B.n647 B.n646 585
R29 B.n648 B.n103 585
R30 B.n650 B.n649 585
R31 B.n652 B.n102 585
R32 B.n655 B.n654 585
R33 B.n656 B.n101 585
R34 B.n658 B.n657 585
R35 B.n660 B.n100 585
R36 B.n663 B.n662 585
R37 B.n664 B.n99 585
R38 B.n666 B.n665 585
R39 B.n668 B.n98 585
R40 B.n671 B.n670 585
R41 B.n672 B.n97 585
R42 B.n674 B.n673 585
R43 B.n676 B.n96 585
R44 B.n679 B.n678 585
R45 B.n680 B.n95 585
R46 B.n682 B.n681 585
R47 B.n684 B.n94 585
R48 B.n687 B.n686 585
R49 B.n688 B.n93 585
R50 B.n690 B.n689 585
R51 B.n692 B.n92 585
R52 B.n695 B.n694 585
R53 B.n696 B.n91 585
R54 B.n698 B.n697 585
R55 B.n700 B.n90 585
R56 B.n702 B.n701 585
R57 B.n704 B.n703 585
R58 B.n707 B.n706 585
R59 B.n708 B.n85 585
R60 B.n710 B.n709 585
R61 B.n712 B.n84 585
R62 B.n715 B.n714 585
R63 B.n716 B.n83 585
R64 B.n718 B.n717 585
R65 B.n720 B.n82 585
R66 B.n723 B.n722 585
R67 B.n725 B.n79 585
R68 B.n727 B.n726 585
R69 B.n729 B.n78 585
R70 B.n732 B.n731 585
R71 B.n733 B.n77 585
R72 B.n735 B.n734 585
R73 B.n737 B.n76 585
R74 B.n740 B.n739 585
R75 B.n741 B.n75 585
R76 B.n743 B.n742 585
R77 B.n745 B.n74 585
R78 B.n748 B.n747 585
R79 B.n749 B.n73 585
R80 B.n751 B.n750 585
R81 B.n753 B.n72 585
R82 B.n756 B.n755 585
R83 B.n757 B.n71 585
R84 B.n759 B.n758 585
R85 B.n761 B.n70 585
R86 B.n764 B.n763 585
R87 B.n765 B.n69 585
R88 B.n767 B.n766 585
R89 B.n769 B.n68 585
R90 B.n772 B.n771 585
R91 B.n773 B.n67 585
R92 B.n775 B.n774 585
R93 B.n777 B.n66 585
R94 B.n780 B.n779 585
R95 B.n781 B.n65 585
R96 B.n783 B.n782 585
R97 B.n785 B.n64 585
R98 B.n788 B.n787 585
R99 B.n789 B.n63 585
R100 B.n791 B.n790 585
R101 B.n793 B.n62 585
R102 B.n796 B.n795 585
R103 B.n797 B.n61 585
R104 B.n799 B.n798 585
R105 B.n801 B.n60 585
R106 B.n804 B.n803 585
R107 B.n805 B.n59 585
R108 B.n807 B.n806 585
R109 B.n809 B.n58 585
R110 B.n812 B.n811 585
R111 B.n813 B.n57 585
R112 B.n815 B.n814 585
R113 B.n817 B.n56 585
R114 B.n820 B.n819 585
R115 B.n821 B.n55 585
R116 B.n823 B.n822 585
R117 B.n825 B.n54 585
R118 B.n828 B.n827 585
R119 B.n829 B.n53 585
R120 B.n831 B.n830 585
R121 B.n833 B.n52 585
R122 B.n836 B.n835 585
R123 B.n837 B.n51 585
R124 B.n591 B.n49 585
R125 B.n840 B.n49 585
R126 B.n590 B.n48 585
R127 B.n841 B.n48 585
R128 B.n589 B.n47 585
R129 B.n842 B.n47 585
R130 B.n588 B.n587 585
R131 B.n587 B.n43 585
R132 B.n586 B.n42 585
R133 B.n848 B.n42 585
R134 B.n585 B.n41 585
R135 B.n849 B.n41 585
R136 B.n584 B.n40 585
R137 B.n850 B.n40 585
R138 B.n583 B.n582 585
R139 B.n582 B.n39 585
R140 B.n581 B.n35 585
R141 B.n856 B.n35 585
R142 B.n580 B.n34 585
R143 B.n857 B.n34 585
R144 B.n579 B.n33 585
R145 B.n858 B.n33 585
R146 B.n578 B.n577 585
R147 B.n577 B.n29 585
R148 B.n576 B.n28 585
R149 B.n864 B.n28 585
R150 B.n575 B.n27 585
R151 B.n865 B.n27 585
R152 B.n574 B.n26 585
R153 B.n866 B.n26 585
R154 B.n573 B.n572 585
R155 B.n572 B.n22 585
R156 B.n571 B.n21 585
R157 B.n872 B.n21 585
R158 B.n570 B.n20 585
R159 B.n873 B.n20 585
R160 B.n569 B.n19 585
R161 B.n874 B.n19 585
R162 B.n568 B.n567 585
R163 B.n567 B.n18 585
R164 B.n566 B.n14 585
R165 B.n880 B.n14 585
R166 B.n565 B.n13 585
R167 B.n881 B.n13 585
R168 B.n564 B.n12 585
R169 B.n882 B.n12 585
R170 B.n563 B.n562 585
R171 B.n562 B.n8 585
R172 B.n561 B.n7 585
R173 B.n888 B.n7 585
R174 B.n560 B.n6 585
R175 B.n889 B.n6 585
R176 B.n559 B.n5 585
R177 B.n890 B.n5 585
R178 B.n558 B.n557 585
R179 B.n557 B.n4 585
R180 B.n556 B.n118 585
R181 B.n556 B.n555 585
R182 B.n546 B.n119 585
R183 B.n120 B.n119 585
R184 B.n548 B.n547 585
R185 B.n549 B.n548 585
R186 B.n545 B.n125 585
R187 B.n125 B.n124 585
R188 B.n544 B.n543 585
R189 B.n543 B.n542 585
R190 B.n127 B.n126 585
R191 B.n535 B.n127 585
R192 B.n534 B.n533 585
R193 B.n536 B.n534 585
R194 B.n532 B.n132 585
R195 B.n132 B.n131 585
R196 B.n531 B.n530 585
R197 B.n530 B.n529 585
R198 B.n134 B.n133 585
R199 B.n135 B.n134 585
R200 B.n522 B.n521 585
R201 B.n523 B.n522 585
R202 B.n520 B.n140 585
R203 B.n140 B.n139 585
R204 B.n519 B.n518 585
R205 B.n518 B.n517 585
R206 B.n142 B.n141 585
R207 B.n143 B.n142 585
R208 B.n510 B.n509 585
R209 B.n511 B.n510 585
R210 B.n508 B.n148 585
R211 B.n148 B.n147 585
R212 B.n507 B.n506 585
R213 B.n506 B.n505 585
R214 B.n150 B.n149 585
R215 B.n498 B.n150 585
R216 B.n497 B.n496 585
R217 B.n499 B.n497 585
R218 B.n495 B.n155 585
R219 B.n155 B.n154 585
R220 B.n494 B.n493 585
R221 B.n493 B.n492 585
R222 B.n157 B.n156 585
R223 B.n158 B.n157 585
R224 B.n485 B.n484 585
R225 B.n486 B.n485 585
R226 B.n483 B.n163 585
R227 B.n163 B.n162 585
R228 B.n482 B.n481 585
R229 B.n481 B.n480 585
R230 B.n477 B.n167 585
R231 B.n476 B.n475 585
R232 B.n473 B.n168 585
R233 B.n473 B.n166 585
R234 B.n472 B.n471 585
R235 B.n470 B.n469 585
R236 B.n468 B.n170 585
R237 B.n466 B.n465 585
R238 B.n464 B.n171 585
R239 B.n463 B.n462 585
R240 B.n460 B.n172 585
R241 B.n458 B.n457 585
R242 B.n456 B.n173 585
R243 B.n455 B.n454 585
R244 B.n452 B.n174 585
R245 B.n450 B.n449 585
R246 B.n448 B.n175 585
R247 B.n447 B.n446 585
R248 B.n444 B.n176 585
R249 B.n442 B.n441 585
R250 B.n440 B.n177 585
R251 B.n439 B.n438 585
R252 B.n436 B.n178 585
R253 B.n434 B.n433 585
R254 B.n432 B.n179 585
R255 B.n431 B.n430 585
R256 B.n428 B.n180 585
R257 B.n426 B.n425 585
R258 B.n424 B.n181 585
R259 B.n423 B.n422 585
R260 B.n420 B.n182 585
R261 B.n418 B.n417 585
R262 B.n416 B.n183 585
R263 B.n415 B.n414 585
R264 B.n412 B.n184 585
R265 B.n410 B.n409 585
R266 B.n408 B.n185 585
R267 B.n407 B.n406 585
R268 B.n404 B.n186 585
R269 B.n402 B.n401 585
R270 B.n400 B.n187 585
R271 B.n399 B.n398 585
R272 B.n396 B.n188 585
R273 B.n394 B.n393 585
R274 B.n392 B.n189 585
R275 B.n391 B.n390 585
R276 B.n388 B.n190 585
R277 B.n386 B.n385 585
R278 B.n384 B.n191 585
R279 B.n383 B.n382 585
R280 B.n380 B.n192 585
R281 B.n378 B.n377 585
R282 B.n376 B.n193 585
R283 B.n375 B.n374 585
R284 B.n372 B.n194 585
R285 B.n370 B.n369 585
R286 B.n368 B.n195 585
R287 B.n367 B.n366 585
R288 B.n364 B.n363 585
R289 B.n362 B.n361 585
R290 B.n360 B.n200 585
R291 B.n358 B.n357 585
R292 B.n356 B.n201 585
R293 B.n355 B.n354 585
R294 B.n352 B.n202 585
R295 B.n350 B.n349 585
R296 B.n348 B.n203 585
R297 B.n346 B.n345 585
R298 B.n343 B.n206 585
R299 B.n341 B.n340 585
R300 B.n339 B.n207 585
R301 B.n338 B.n337 585
R302 B.n335 B.n208 585
R303 B.n333 B.n332 585
R304 B.n331 B.n209 585
R305 B.n330 B.n329 585
R306 B.n327 B.n210 585
R307 B.n325 B.n324 585
R308 B.n323 B.n211 585
R309 B.n322 B.n321 585
R310 B.n319 B.n212 585
R311 B.n317 B.n316 585
R312 B.n315 B.n213 585
R313 B.n314 B.n313 585
R314 B.n311 B.n214 585
R315 B.n309 B.n308 585
R316 B.n307 B.n215 585
R317 B.n306 B.n305 585
R318 B.n303 B.n216 585
R319 B.n301 B.n300 585
R320 B.n299 B.n217 585
R321 B.n298 B.n297 585
R322 B.n295 B.n218 585
R323 B.n293 B.n292 585
R324 B.n291 B.n219 585
R325 B.n290 B.n289 585
R326 B.n287 B.n220 585
R327 B.n285 B.n284 585
R328 B.n283 B.n221 585
R329 B.n282 B.n281 585
R330 B.n279 B.n222 585
R331 B.n277 B.n276 585
R332 B.n275 B.n223 585
R333 B.n274 B.n273 585
R334 B.n271 B.n224 585
R335 B.n269 B.n268 585
R336 B.n267 B.n225 585
R337 B.n266 B.n265 585
R338 B.n263 B.n226 585
R339 B.n261 B.n260 585
R340 B.n259 B.n227 585
R341 B.n258 B.n257 585
R342 B.n255 B.n228 585
R343 B.n253 B.n252 585
R344 B.n251 B.n229 585
R345 B.n250 B.n249 585
R346 B.n247 B.n230 585
R347 B.n245 B.n244 585
R348 B.n243 B.n231 585
R349 B.n242 B.n241 585
R350 B.n239 B.n232 585
R351 B.n237 B.n236 585
R352 B.n235 B.n234 585
R353 B.n165 B.n164 585
R354 B.n479 B.n478 585
R355 B.n480 B.n479 585
R356 B.n161 B.n160 585
R357 B.n162 B.n161 585
R358 B.n488 B.n487 585
R359 B.n487 B.n486 585
R360 B.n489 B.n159 585
R361 B.n159 B.n158 585
R362 B.n491 B.n490 585
R363 B.n492 B.n491 585
R364 B.n153 B.n152 585
R365 B.n154 B.n153 585
R366 B.n501 B.n500 585
R367 B.n500 B.n499 585
R368 B.n502 B.n151 585
R369 B.n498 B.n151 585
R370 B.n504 B.n503 585
R371 B.n505 B.n504 585
R372 B.n146 B.n145 585
R373 B.n147 B.n146 585
R374 B.n513 B.n512 585
R375 B.n512 B.n511 585
R376 B.n514 B.n144 585
R377 B.n144 B.n143 585
R378 B.n516 B.n515 585
R379 B.n517 B.n516 585
R380 B.n138 B.n137 585
R381 B.n139 B.n138 585
R382 B.n525 B.n524 585
R383 B.n524 B.n523 585
R384 B.n526 B.n136 585
R385 B.n136 B.n135 585
R386 B.n528 B.n527 585
R387 B.n529 B.n528 585
R388 B.n130 B.n129 585
R389 B.n131 B.n130 585
R390 B.n538 B.n537 585
R391 B.n537 B.n536 585
R392 B.n539 B.n128 585
R393 B.n535 B.n128 585
R394 B.n541 B.n540 585
R395 B.n542 B.n541 585
R396 B.n123 B.n122 585
R397 B.n124 B.n123 585
R398 B.n551 B.n550 585
R399 B.n550 B.n549 585
R400 B.n552 B.n121 585
R401 B.n121 B.n120 585
R402 B.n554 B.n553 585
R403 B.n555 B.n554 585
R404 B.n2 B.n0 585
R405 B.n4 B.n2 585
R406 B.n3 B.n1 585
R407 B.n889 B.n3 585
R408 B.n887 B.n886 585
R409 B.n888 B.n887 585
R410 B.n885 B.n9 585
R411 B.n9 B.n8 585
R412 B.n884 B.n883 585
R413 B.n883 B.n882 585
R414 B.n11 B.n10 585
R415 B.n881 B.n11 585
R416 B.n879 B.n878 585
R417 B.n880 B.n879 585
R418 B.n877 B.n15 585
R419 B.n18 B.n15 585
R420 B.n876 B.n875 585
R421 B.n875 B.n874 585
R422 B.n17 B.n16 585
R423 B.n873 B.n17 585
R424 B.n871 B.n870 585
R425 B.n872 B.n871 585
R426 B.n869 B.n23 585
R427 B.n23 B.n22 585
R428 B.n868 B.n867 585
R429 B.n867 B.n866 585
R430 B.n25 B.n24 585
R431 B.n865 B.n25 585
R432 B.n863 B.n862 585
R433 B.n864 B.n863 585
R434 B.n861 B.n30 585
R435 B.n30 B.n29 585
R436 B.n860 B.n859 585
R437 B.n859 B.n858 585
R438 B.n32 B.n31 585
R439 B.n857 B.n32 585
R440 B.n855 B.n854 585
R441 B.n856 B.n855 585
R442 B.n853 B.n36 585
R443 B.n39 B.n36 585
R444 B.n852 B.n851 585
R445 B.n851 B.n850 585
R446 B.n38 B.n37 585
R447 B.n849 B.n38 585
R448 B.n847 B.n846 585
R449 B.n848 B.n847 585
R450 B.n845 B.n44 585
R451 B.n44 B.n43 585
R452 B.n844 B.n843 585
R453 B.n843 B.n842 585
R454 B.n46 B.n45 585
R455 B.n841 B.n46 585
R456 B.n839 B.n838 585
R457 B.n840 B.n839 585
R458 B.n892 B.n891 585
R459 B.n891 B.n890 585
R460 B.n479 B.n167 506.916
R461 B.n839 B.n51 506.916
R462 B.n481 B.n165 506.916
R463 B.n117 B.n49 506.916
R464 B.n204 B.t13 358.567
R465 B.n196 B.t2 358.567
R466 B.n80 B.t10 358.567
R467 B.n86 B.t6 358.567
R468 B.n595 B.n50 256.663
R469 B.n597 B.n50 256.663
R470 B.n603 B.n50 256.663
R471 B.n605 B.n50 256.663
R472 B.n611 B.n50 256.663
R473 B.n613 B.n50 256.663
R474 B.n619 B.n50 256.663
R475 B.n621 B.n50 256.663
R476 B.n627 B.n50 256.663
R477 B.n629 B.n50 256.663
R478 B.n635 B.n50 256.663
R479 B.n637 B.n50 256.663
R480 B.n643 B.n50 256.663
R481 B.n645 B.n50 256.663
R482 B.n651 B.n50 256.663
R483 B.n653 B.n50 256.663
R484 B.n659 B.n50 256.663
R485 B.n661 B.n50 256.663
R486 B.n667 B.n50 256.663
R487 B.n669 B.n50 256.663
R488 B.n675 B.n50 256.663
R489 B.n677 B.n50 256.663
R490 B.n683 B.n50 256.663
R491 B.n685 B.n50 256.663
R492 B.n691 B.n50 256.663
R493 B.n693 B.n50 256.663
R494 B.n699 B.n50 256.663
R495 B.n89 B.n50 256.663
R496 B.n705 B.n50 256.663
R497 B.n711 B.n50 256.663
R498 B.n713 B.n50 256.663
R499 B.n719 B.n50 256.663
R500 B.n721 B.n50 256.663
R501 B.n728 B.n50 256.663
R502 B.n730 B.n50 256.663
R503 B.n736 B.n50 256.663
R504 B.n738 B.n50 256.663
R505 B.n744 B.n50 256.663
R506 B.n746 B.n50 256.663
R507 B.n752 B.n50 256.663
R508 B.n754 B.n50 256.663
R509 B.n760 B.n50 256.663
R510 B.n762 B.n50 256.663
R511 B.n768 B.n50 256.663
R512 B.n770 B.n50 256.663
R513 B.n776 B.n50 256.663
R514 B.n778 B.n50 256.663
R515 B.n784 B.n50 256.663
R516 B.n786 B.n50 256.663
R517 B.n792 B.n50 256.663
R518 B.n794 B.n50 256.663
R519 B.n800 B.n50 256.663
R520 B.n802 B.n50 256.663
R521 B.n808 B.n50 256.663
R522 B.n810 B.n50 256.663
R523 B.n816 B.n50 256.663
R524 B.n818 B.n50 256.663
R525 B.n824 B.n50 256.663
R526 B.n826 B.n50 256.663
R527 B.n832 B.n50 256.663
R528 B.n834 B.n50 256.663
R529 B.n474 B.n166 256.663
R530 B.n169 B.n166 256.663
R531 B.n467 B.n166 256.663
R532 B.n461 B.n166 256.663
R533 B.n459 B.n166 256.663
R534 B.n453 B.n166 256.663
R535 B.n451 B.n166 256.663
R536 B.n445 B.n166 256.663
R537 B.n443 B.n166 256.663
R538 B.n437 B.n166 256.663
R539 B.n435 B.n166 256.663
R540 B.n429 B.n166 256.663
R541 B.n427 B.n166 256.663
R542 B.n421 B.n166 256.663
R543 B.n419 B.n166 256.663
R544 B.n413 B.n166 256.663
R545 B.n411 B.n166 256.663
R546 B.n405 B.n166 256.663
R547 B.n403 B.n166 256.663
R548 B.n397 B.n166 256.663
R549 B.n395 B.n166 256.663
R550 B.n389 B.n166 256.663
R551 B.n387 B.n166 256.663
R552 B.n381 B.n166 256.663
R553 B.n379 B.n166 256.663
R554 B.n373 B.n166 256.663
R555 B.n371 B.n166 256.663
R556 B.n365 B.n166 256.663
R557 B.n199 B.n166 256.663
R558 B.n359 B.n166 256.663
R559 B.n353 B.n166 256.663
R560 B.n351 B.n166 256.663
R561 B.n344 B.n166 256.663
R562 B.n342 B.n166 256.663
R563 B.n336 B.n166 256.663
R564 B.n334 B.n166 256.663
R565 B.n328 B.n166 256.663
R566 B.n326 B.n166 256.663
R567 B.n320 B.n166 256.663
R568 B.n318 B.n166 256.663
R569 B.n312 B.n166 256.663
R570 B.n310 B.n166 256.663
R571 B.n304 B.n166 256.663
R572 B.n302 B.n166 256.663
R573 B.n296 B.n166 256.663
R574 B.n294 B.n166 256.663
R575 B.n288 B.n166 256.663
R576 B.n286 B.n166 256.663
R577 B.n280 B.n166 256.663
R578 B.n278 B.n166 256.663
R579 B.n272 B.n166 256.663
R580 B.n270 B.n166 256.663
R581 B.n264 B.n166 256.663
R582 B.n262 B.n166 256.663
R583 B.n256 B.n166 256.663
R584 B.n254 B.n166 256.663
R585 B.n248 B.n166 256.663
R586 B.n246 B.n166 256.663
R587 B.n240 B.n166 256.663
R588 B.n238 B.n166 256.663
R589 B.n233 B.n166 256.663
R590 B.n479 B.n161 163.367
R591 B.n487 B.n161 163.367
R592 B.n487 B.n159 163.367
R593 B.n491 B.n159 163.367
R594 B.n491 B.n153 163.367
R595 B.n500 B.n153 163.367
R596 B.n500 B.n151 163.367
R597 B.n504 B.n151 163.367
R598 B.n504 B.n146 163.367
R599 B.n512 B.n146 163.367
R600 B.n512 B.n144 163.367
R601 B.n516 B.n144 163.367
R602 B.n516 B.n138 163.367
R603 B.n524 B.n138 163.367
R604 B.n524 B.n136 163.367
R605 B.n528 B.n136 163.367
R606 B.n528 B.n130 163.367
R607 B.n537 B.n130 163.367
R608 B.n537 B.n128 163.367
R609 B.n541 B.n128 163.367
R610 B.n541 B.n123 163.367
R611 B.n550 B.n123 163.367
R612 B.n550 B.n121 163.367
R613 B.n554 B.n121 163.367
R614 B.n554 B.n2 163.367
R615 B.n891 B.n2 163.367
R616 B.n891 B.n3 163.367
R617 B.n887 B.n3 163.367
R618 B.n887 B.n9 163.367
R619 B.n883 B.n9 163.367
R620 B.n883 B.n11 163.367
R621 B.n879 B.n11 163.367
R622 B.n879 B.n15 163.367
R623 B.n875 B.n15 163.367
R624 B.n875 B.n17 163.367
R625 B.n871 B.n17 163.367
R626 B.n871 B.n23 163.367
R627 B.n867 B.n23 163.367
R628 B.n867 B.n25 163.367
R629 B.n863 B.n25 163.367
R630 B.n863 B.n30 163.367
R631 B.n859 B.n30 163.367
R632 B.n859 B.n32 163.367
R633 B.n855 B.n32 163.367
R634 B.n855 B.n36 163.367
R635 B.n851 B.n36 163.367
R636 B.n851 B.n38 163.367
R637 B.n847 B.n38 163.367
R638 B.n847 B.n44 163.367
R639 B.n843 B.n44 163.367
R640 B.n843 B.n46 163.367
R641 B.n839 B.n46 163.367
R642 B.n475 B.n473 163.367
R643 B.n473 B.n472 163.367
R644 B.n469 B.n468 163.367
R645 B.n466 B.n171 163.367
R646 B.n462 B.n460 163.367
R647 B.n458 B.n173 163.367
R648 B.n454 B.n452 163.367
R649 B.n450 B.n175 163.367
R650 B.n446 B.n444 163.367
R651 B.n442 B.n177 163.367
R652 B.n438 B.n436 163.367
R653 B.n434 B.n179 163.367
R654 B.n430 B.n428 163.367
R655 B.n426 B.n181 163.367
R656 B.n422 B.n420 163.367
R657 B.n418 B.n183 163.367
R658 B.n414 B.n412 163.367
R659 B.n410 B.n185 163.367
R660 B.n406 B.n404 163.367
R661 B.n402 B.n187 163.367
R662 B.n398 B.n396 163.367
R663 B.n394 B.n189 163.367
R664 B.n390 B.n388 163.367
R665 B.n386 B.n191 163.367
R666 B.n382 B.n380 163.367
R667 B.n378 B.n193 163.367
R668 B.n374 B.n372 163.367
R669 B.n370 B.n195 163.367
R670 B.n366 B.n364 163.367
R671 B.n361 B.n360 163.367
R672 B.n358 B.n201 163.367
R673 B.n354 B.n352 163.367
R674 B.n350 B.n203 163.367
R675 B.n345 B.n343 163.367
R676 B.n341 B.n207 163.367
R677 B.n337 B.n335 163.367
R678 B.n333 B.n209 163.367
R679 B.n329 B.n327 163.367
R680 B.n325 B.n211 163.367
R681 B.n321 B.n319 163.367
R682 B.n317 B.n213 163.367
R683 B.n313 B.n311 163.367
R684 B.n309 B.n215 163.367
R685 B.n305 B.n303 163.367
R686 B.n301 B.n217 163.367
R687 B.n297 B.n295 163.367
R688 B.n293 B.n219 163.367
R689 B.n289 B.n287 163.367
R690 B.n285 B.n221 163.367
R691 B.n281 B.n279 163.367
R692 B.n277 B.n223 163.367
R693 B.n273 B.n271 163.367
R694 B.n269 B.n225 163.367
R695 B.n265 B.n263 163.367
R696 B.n261 B.n227 163.367
R697 B.n257 B.n255 163.367
R698 B.n253 B.n229 163.367
R699 B.n249 B.n247 163.367
R700 B.n245 B.n231 163.367
R701 B.n241 B.n239 163.367
R702 B.n237 B.n234 163.367
R703 B.n481 B.n163 163.367
R704 B.n485 B.n163 163.367
R705 B.n485 B.n157 163.367
R706 B.n493 B.n157 163.367
R707 B.n493 B.n155 163.367
R708 B.n497 B.n155 163.367
R709 B.n497 B.n150 163.367
R710 B.n506 B.n150 163.367
R711 B.n506 B.n148 163.367
R712 B.n510 B.n148 163.367
R713 B.n510 B.n142 163.367
R714 B.n518 B.n142 163.367
R715 B.n518 B.n140 163.367
R716 B.n522 B.n140 163.367
R717 B.n522 B.n134 163.367
R718 B.n530 B.n134 163.367
R719 B.n530 B.n132 163.367
R720 B.n534 B.n132 163.367
R721 B.n534 B.n127 163.367
R722 B.n543 B.n127 163.367
R723 B.n543 B.n125 163.367
R724 B.n548 B.n125 163.367
R725 B.n548 B.n119 163.367
R726 B.n556 B.n119 163.367
R727 B.n557 B.n556 163.367
R728 B.n557 B.n5 163.367
R729 B.n6 B.n5 163.367
R730 B.n7 B.n6 163.367
R731 B.n562 B.n7 163.367
R732 B.n562 B.n12 163.367
R733 B.n13 B.n12 163.367
R734 B.n14 B.n13 163.367
R735 B.n567 B.n14 163.367
R736 B.n567 B.n19 163.367
R737 B.n20 B.n19 163.367
R738 B.n21 B.n20 163.367
R739 B.n572 B.n21 163.367
R740 B.n572 B.n26 163.367
R741 B.n27 B.n26 163.367
R742 B.n28 B.n27 163.367
R743 B.n577 B.n28 163.367
R744 B.n577 B.n33 163.367
R745 B.n34 B.n33 163.367
R746 B.n35 B.n34 163.367
R747 B.n582 B.n35 163.367
R748 B.n582 B.n40 163.367
R749 B.n41 B.n40 163.367
R750 B.n42 B.n41 163.367
R751 B.n587 B.n42 163.367
R752 B.n587 B.n47 163.367
R753 B.n48 B.n47 163.367
R754 B.n49 B.n48 163.367
R755 B.n835 B.n833 163.367
R756 B.n831 B.n53 163.367
R757 B.n827 B.n825 163.367
R758 B.n823 B.n55 163.367
R759 B.n819 B.n817 163.367
R760 B.n815 B.n57 163.367
R761 B.n811 B.n809 163.367
R762 B.n807 B.n59 163.367
R763 B.n803 B.n801 163.367
R764 B.n799 B.n61 163.367
R765 B.n795 B.n793 163.367
R766 B.n791 B.n63 163.367
R767 B.n787 B.n785 163.367
R768 B.n783 B.n65 163.367
R769 B.n779 B.n777 163.367
R770 B.n775 B.n67 163.367
R771 B.n771 B.n769 163.367
R772 B.n767 B.n69 163.367
R773 B.n763 B.n761 163.367
R774 B.n759 B.n71 163.367
R775 B.n755 B.n753 163.367
R776 B.n751 B.n73 163.367
R777 B.n747 B.n745 163.367
R778 B.n743 B.n75 163.367
R779 B.n739 B.n737 163.367
R780 B.n735 B.n77 163.367
R781 B.n731 B.n729 163.367
R782 B.n727 B.n79 163.367
R783 B.n722 B.n720 163.367
R784 B.n718 B.n83 163.367
R785 B.n714 B.n712 163.367
R786 B.n710 B.n85 163.367
R787 B.n706 B.n704 163.367
R788 B.n701 B.n700 163.367
R789 B.n698 B.n91 163.367
R790 B.n694 B.n692 163.367
R791 B.n690 B.n93 163.367
R792 B.n686 B.n684 163.367
R793 B.n682 B.n95 163.367
R794 B.n678 B.n676 163.367
R795 B.n674 B.n97 163.367
R796 B.n670 B.n668 163.367
R797 B.n666 B.n99 163.367
R798 B.n662 B.n660 163.367
R799 B.n658 B.n101 163.367
R800 B.n654 B.n652 163.367
R801 B.n650 B.n103 163.367
R802 B.n646 B.n644 163.367
R803 B.n642 B.n105 163.367
R804 B.n638 B.n636 163.367
R805 B.n634 B.n107 163.367
R806 B.n630 B.n628 163.367
R807 B.n626 B.n109 163.367
R808 B.n622 B.n620 163.367
R809 B.n618 B.n111 163.367
R810 B.n614 B.n612 163.367
R811 B.n610 B.n113 163.367
R812 B.n606 B.n604 163.367
R813 B.n602 B.n115 163.367
R814 B.n598 B.n596 163.367
R815 B.n594 B.n117 163.367
R816 B.n204 B.t15 128.59
R817 B.n86 B.t8 128.59
R818 B.n196 B.t5 128.569
R819 B.n80 B.t11 128.569
R820 B.n474 B.n167 71.676
R821 B.n472 B.n169 71.676
R822 B.n468 B.n467 71.676
R823 B.n461 B.n171 71.676
R824 B.n460 B.n459 71.676
R825 B.n453 B.n173 71.676
R826 B.n452 B.n451 71.676
R827 B.n445 B.n175 71.676
R828 B.n444 B.n443 71.676
R829 B.n437 B.n177 71.676
R830 B.n436 B.n435 71.676
R831 B.n429 B.n179 71.676
R832 B.n428 B.n427 71.676
R833 B.n421 B.n181 71.676
R834 B.n420 B.n419 71.676
R835 B.n413 B.n183 71.676
R836 B.n412 B.n411 71.676
R837 B.n405 B.n185 71.676
R838 B.n404 B.n403 71.676
R839 B.n397 B.n187 71.676
R840 B.n396 B.n395 71.676
R841 B.n389 B.n189 71.676
R842 B.n388 B.n387 71.676
R843 B.n381 B.n191 71.676
R844 B.n380 B.n379 71.676
R845 B.n373 B.n193 71.676
R846 B.n372 B.n371 71.676
R847 B.n365 B.n195 71.676
R848 B.n364 B.n199 71.676
R849 B.n360 B.n359 71.676
R850 B.n353 B.n201 71.676
R851 B.n352 B.n351 71.676
R852 B.n344 B.n203 71.676
R853 B.n343 B.n342 71.676
R854 B.n336 B.n207 71.676
R855 B.n335 B.n334 71.676
R856 B.n328 B.n209 71.676
R857 B.n327 B.n326 71.676
R858 B.n320 B.n211 71.676
R859 B.n319 B.n318 71.676
R860 B.n312 B.n213 71.676
R861 B.n311 B.n310 71.676
R862 B.n304 B.n215 71.676
R863 B.n303 B.n302 71.676
R864 B.n296 B.n217 71.676
R865 B.n295 B.n294 71.676
R866 B.n288 B.n219 71.676
R867 B.n287 B.n286 71.676
R868 B.n280 B.n221 71.676
R869 B.n279 B.n278 71.676
R870 B.n272 B.n223 71.676
R871 B.n271 B.n270 71.676
R872 B.n264 B.n225 71.676
R873 B.n263 B.n262 71.676
R874 B.n256 B.n227 71.676
R875 B.n255 B.n254 71.676
R876 B.n248 B.n229 71.676
R877 B.n247 B.n246 71.676
R878 B.n240 B.n231 71.676
R879 B.n239 B.n238 71.676
R880 B.n234 B.n233 71.676
R881 B.n834 B.n51 71.676
R882 B.n833 B.n832 71.676
R883 B.n826 B.n53 71.676
R884 B.n825 B.n824 71.676
R885 B.n818 B.n55 71.676
R886 B.n817 B.n816 71.676
R887 B.n810 B.n57 71.676
R888 B.n809 B.n808 71.676
R889 B.n802 B.n59 71.676
R890 B.n801 B.n800 71.676
R891 B.n794 B.n61 71.676
R892 B.n793 B.n792 71.676
R893 B.n786 B.n63 71.676
R894 B.n785 B.n784 71.676
R895 B.n778 B.n65 71.676
R896 B.n777 B.n776 71.676
R897 B.n770 B.n67 71.676
R898 B.n769 B.n768 71.676
R899 B.n762 B.n69 71.676
R900 B.n761 B.n760 71.676
R901 B.n754 B.n71 71.676
R902 B.n753 B.n752 71.676
R903 B.n746 B.n73 71.676
R904 B.n745 B.n744 71.676
R905 B.n738 B.n75 71.676
R906 B.n737 B.n736 71.676
R907 B.n730 B.n77 71.676
R908 B.n729 B.n728 71.676
R909 B.n721 B.n79 71.676
R910 B.n720 B.n719 71.676
R911 B.n713 B.n83 71.676
R912 B.n712 B.n711 71.676
R913 B.n705 B.n85 71.676
R914 B.n704 B.n89 71.676
R915 B.n700 B.n699 71.676
R916 B.n693 B.n91 71.676
R917 B.n692 B.n691 71.676
R918 B.n685 B.n93 71.676
R919 B.n684 B.n683 71.676
R920 B.n677 B.n95 71.676
R921 B.n676 B.n675 71.676
R922 B.n669 B.n97 71.676
R923 B.n668 B.n667 71.676
R924 B.n661 B.n99 71.676
R925 B.n660 B.n659 71.676
R926 B.n653 B.n101 71.676
R927 B.n652 B.n651 71.676
R928 B.n645 B.n103 71.676
R929 B.n644 B.n643 71.676
R930 B.n637 B.n105 71.676
R931 B.n636 B.n635 71.676
R932 B.n629 B.n107 71.676
R933 B.n628 B.n627 71.676
R934 B.n621 B.n109 71.676
R935 B.n620 B.n619 71.676
R936 B.n613 B.n111 71.676
R937 B.n612 B.n611 71.676
R938 B.n605 B.n113 71.676
R939 B.n604 B.n603 71.676
R940 B.n597 B.n115 71.676
R941 B.n596 B.n595 71.676
R942 B.n595 B.n594 71.676
R943 B.n598 B.n597 71.676
R944 B.n603 B.n602 71.676
R945 B.n606 B.n605 71.676
R946 B.n611 B.n610 71.676
R947 B.n614 B.n613 71.676
R948 B.n619 B.n618 71.676
R949 B.n622 B.n621 71.676
R950 B.n627 B.n626 71.676
R951 B.n630 B.n629 71.676
R952 B.n635 B.n634 71.676
R953 B.n638 B.n637 71.676
R954 B.n643 B.n642 71.676
R955 B.n646 B.n645 71.676
R956 B.n651 B.n650 71.676
R957 B.n654 B.n653 71.676
R958 B.n659 B.n658 71.676
R959 B.n662 B.n661 71.676
R960 B.n667 B.n666 71.676
R961 B.n670 B.n669 71.676
R962 B.n675 B.n674 71.676
R963 B.n678 B.n677 71.676
R964 B.n683 B.n682 71.676
R965 B.n686 B.n685 71.676
R966 B.n691 B.n690 71.676
R967 B.n694 B.n693 71.676
R968 B.n699 B.n698 71.676
R969 B.n701 B.n89 71.676
R970 B.n706 B.n705 71.676
R971 B.n711 B.n710 71.676
R972 B.n714 B.n713 71.676
R973 B.n719 B.n718 71.676
R974 B.n722 B.n721 71.676
R975 B.n728 B.n727 71.676
R976 B.n731 B.n730 71.676
R977 B.n736 B.n735 71.676
R978 B.n739 B.n738 71.676
R979 B.n744 B.n743 71.676
R980 B.n747 B.n746 71.676
R981 B.n752 B.n751 71.676
R982 B.n755 B.n754 71.676
R983 B.n760 B.n759 71.676
R984 B.n763 B.n762 71.676
R985 B.n768 B.n767 71.676
R986 B.n771 B.n770 71.676
R987 B.n776 B.n775 71.676
R988 B.n779 B.n778 71.676
R989 B.n784 B.n783 71.676
R990 B.n787 B.n786 71.676
R991 B.n792 B.n791 71.676
R992 B.n795 B.n794 71.676
R993 B.n800 B.n799 71.676
R994 B.n803 B.n802 71.676
R995 B.n808 B.n807 71.676
R996 B.n811 B.n810 71.676
R997 B.n816 B.n815 71.676
R998 B.n819 B.n818 71.676
R999 B.n824 B.n823 71.676
R1000 B.n827 B.n826 71.676
R1001 B.n832 B.n831 71.676
R1002 B.n835 B.n834 71.676
R1003 B.n475 B.n474 71.676
R1004 B.n469 B.n169 71.676
R1005 B.n467 B.n466 71.676
R1006 B.n462 B.n461 71.676
R1007 B.n459 B.n458 71.676
R1008 B.n454 B.n453 71.676
R1009 B.n451 B.n450 71.676
R1010 B.n446 B.n445 71.676
R1011 B.n443 B.n442 71.676
R1012 B.n438 B.n437 71.676
R1013 B.n435 B.n434 71.676
R1014 B.n430 B.n429 71.676
R1015 B.n427 B.n426 71.676
R1016 B.n422 B.n421 71.676
R1017 B.n419 B.n418 71.676
R1018 B.n414 B.n413 71.676
R1019 B.n411 B.n410 71.676
R1020 B.n406 B.n405 71.676
R1021 B.n403 B.n402 71.676
R1022 B.n398 B.n397 71.676
R1023 B.n395 B.n394 71.676
R1024 B.n390 B.n389 71.676
R1025 B.n387 B.n386 71.676
R1026 B.n382 B.n381 71.676
R1027 B.n379 B.n378 71.676
R1028 B.n374 B.n373 71.676
R1029 B.n371 B.n370 71.676
R1030 B.n366 B.n365 71.676
R1031 B.n361 B.n199 71.676
R1032 B.n359 B.n358 71.676
R1033 B.n354 B.n353 71.676
R1034 B.n351 B.n350 71.676
R1035 B.n345 B.n344 71.676
R1036 B.n342 B.n341 71.676
R1037 B.n337 B.n336 71.676
R1038 B.n334 B.n333 71.676
R1039 B.n329 B.n328 71.676
R1040 B.n326 B.n325 71.676
R1041 B.n321 B.n320 71.676
R1042 B.n318 B.n317 71.676
R1043 B.n313 B.n312 71.676
R1044 B.n310 B.n309 71.676
R1045 B.n305 B.n304 71.676
R1046 B.n302 B.n301 71.676
R1047 B.n297 B.n296 71.676
R1048 B.n294 B.n293 71.676
R1049 B.n289 B.n288 71.676
R1050 B.n286 B.n285 71.676
R1051 B.n281 B.n280 71.676
R1052 B.n278 B.n277 71.676
R1053 B.n273 B.n272 71.676
R1054 B.n270 B.n269 71.676
R1055 B.n265 B.n264 71.676
R1056 B.n262 B.n261 71.676
R1057 B.n257 B.n256 71.676
R1058 B.n254 B.n253 71.676
R1059 B.n249 B.n248 71.676
R1060 B.n246 B.n245 71.676
R1061 B.n241 B.n240 71.676
R1062 B.n238 B.n237 71.676
R1063 B.n233 B.n165 71.676
R1064 B.n205 B.t14 69.0514
R1065 B.n87 B.t9 69.0514
R1066 B.n197 B.t4 69.0287
R1067 B.n81 B.t12 69.0287
R1068 B.n480 B.n166 66.3989
R1069 B.n840 B.n50 66.3989
R1070 B.n347 B.n205 59.5399
R1071 B.n205 B.n204 59.5399
R1072 B.n198 B.n197 59.5399
R1073 B.n197 B.n196 59.5399
R1074 B.n81 B.n80 59.5399
R1075 B.n724 B.n81 59.5399
R1076 B.n87 B.n86 59.5399
R1077 B.n88 B.n87 59.5399
R1078 B.n480 B.n162 33.4456
R1079 B.n486 B.n162 33.4456
R1080 B.n486 B.n158 33.4456
R1081 B.n492 B.n158 33.4456
R1082 B.n492 B.n154 33.4456
R1083 B.n499 B.n154 33.4456
R1084 B.n499 B.n498 33.4456
R1085 B.n505 B.n147 33.4456
R1086 B.n511 B.n147 33.4456
R1087 B.n511 B.n143 33.4456
R1088 B.n517 B.n143 33.4456
R1089 B.n517 B.n139 33.4456
R1090 B.n523 B.n139 33.4456
R1091 B.n523 B.n135 33.4456
R1092 B.n529 B.n135 33.4456
R1093 B.n529 B.n131 33.4456
R1094 B.n536 B.n131 33.4456
R1095 B.n536 B.n535 33.4456
R1096 B.n542 B.n124 33.4456
R1097 B.n549 B.n124 33.4456
R1098 B.n549 B.n120 33.4456
R1099 B.n555 B.n120 33.4456
R1100 B.n555 B.n4 33.4456
R1101 B.n890 B.n4 33.4456
R1102 B.n890 B.n889 33.4456
R1103 B.n889 B.n888 33.4456
R1104 B.n888 B.n8 33.4456
R1105 B.n882 B.n8 33.4456
R1106 B.n882 B.n881 33.4456
R1107 B.n881 B.n880 33.4456
R1108 B.n874 B.n18 33.4456
R1109 B.n874 B.n873 33.4456
R1110 B.n873 B.n872 33.4456
R1111 B.n872 B.n22 33.4456
R1112 B.n866 B.n22 33.4456
R1113 B.n866 B.n865 33.4456
R1114 B.n865 B.n864 33.4456
R1115 B.n864 B.n29 33.4456
R1116 B.n858 B.n29 33.4456
R1117 B.n858 B.n857 33.4456
R1118 B.n857 B.n856 33.4456
R1119 B.n850 B.n39 33.4456
R1120 B.n850 B.n849 33.4456
R1121 B.n849 B.n848 33.4456
R1122 B.n848 B.n43 33.4456
R1123 B.n842 B.n43 33.4456
R1124 B.n842 B.n841 33.4456
R1125 B.n841 B.n840 33.4456
R1126 B.n838 B.n837 32.9371
R1127 B.n592 B.n591 32.9371
R1128 B.n482 B.n164 32.9371
R1129 B.n478 B.n477 32.9371
R1130 B.n535 B.t0 29.5109
R1131 B.n18 B.t1 29.5109
R1132 B.n498 B.t3 21.6415
R1133 B.n39 B.t7 21.6415
R1134 B B.n892 18.0485
R1135 B.n505 B.t3 11.8047
R1136 B.n856 B.t7 11.8047
R1137 B.n837 B.n836 10.6151
R1138 B.n836 B.n52 10.6151
R1139 B.n830 B.n52 10.6151
R1140 B.n830 B.n829 10.6151
R1141 B.n829 B.n828 10.6151
R1142 B.n828 B.n54 10.6151
R1143 B.n822 B.n54 10.6151
R1144 B.n822 B.n821 10.6151
R1145 B.n821 B.n820 10.6151
R1146 B.n820 B.n56 10.6151
R1147 B.n814 B.n56 10.6151
R1148 B.n814 B.n813 10.6151
R1149 B.n813 B.n812 10.6151
R1150 B.n812 B.n58 10.6151
R1151 B.n806 B.n58 10.6151
R1152 B.n806 B.n805 10.6151
R1153 B.n805 B.n804 10.6151
R1154 B.n804 B.n60 10.6151
R1155 B.n798 B.n60 10.6151
R1156 B.n798 B.n797 10.6151
R1157 B.n797 B.n796 10.6151
R1158 B.n796 B.n62 10.6151
R1159 B.n790 B.n62 10.6151
R1160 B.n790 B.n789 10.6151
R1161 B.n789 B.n788 10.6151
R1162 B.n788 B.n64 10.6151
R1163 B.n782 B.n64 10.6151
R1164 B.n782 B.n781 10.6151
R1165 B.n781 B.n780 10.6151
R1166 B.n780 B.n66 10.6151
R1167 B.n774 B.n66 10.6151
R1168 B.n774 B.n773 10.6151
R1169 B.n773 B.n772 10.6151
R1170 B.n772 B.n68 10.6151
R1171 B.n766 B.n68 10.6151
R1172 B.n766 B.n765 10.6151
R1173 B.n765 B.n764 10.6151
R1174 B.n764 B.n70 10.6151
R1175 B.n758 B.n70 10.6151
R1176 B.n758 B.n757 10.6151
R1177 B.n757 B.n756 10.6151
R1178 B.n756 B.n72 10.6151
R1179 B.n750 B.n72 10.6151
R1180 B.n750 B.n749 10.6151
R1181 B.n749 B.n748 10.6151
R1182 B.n748 B.n74 10.6151
R1183 B.n742 B.n74 10.6151
R1184 B.n742 B.n741 10.6151
R1185 B.n741 B.n740 10.6151
R1186 B.n740 B.n76 10.6151
R1187 B.n734 B.n76 10.6151
R1188 B.n734 B.n733 10.6151
R1189 B.n733 B.n732 10.6151
R1190 B.n732 B.n78 10.6151
R1191 B.n726 B.n78 10.6151
R1192 B.n726 B.n725 10.6151
R1193 B.n723 B.n82 10.6151
R1194 B.n717 B.n82 10.6151
R1195 B.n717 B.n716 10.6151
R1196 B.n716 B.n715 10.6151
R1197 B.n715 B.n84 10.6151
R1198 B.n709 B.n84 10.6151
R1199 B.n709 B.n708 10.6151
R1200 B.n708 B.n707 10.6151
R1201 B.n703 B.n702 10.6151
R1202 B.n702 B.n90 10.6151
R1203 B.n697 B.n90 10.6151
R1204 B.n697 B.n696 10.6151
R1205 B.n696 B.n695 10.6151
R1206 B.n695 B.n92 10.6151
R1207 B.n689 B.n92 10.6151
R1208 B.n689 B.n688 10.6151
R1209 B.n688 B.n687 10.6151
R1210 B.n687 B.n94 10.6151
R1211 B.n681 B.n94 10.6151
R1212 B.n681 B.n680 10.6151
R1213 B.n680 B.n679 10.6151
R1214 B.n679 B.n96 10.6151
R1215 B.n673 B.n96 10.6151
R1216 B.n673 B.n672 10.6151
R1217 B.n672 B.n671 10.6151
R1218 B.n671 B.n98 10.6151
R1219 B.n665 B.n98 10.6151
R1220 B.n665 B.n664 10.6151
R1221 B.n664 B.n663 10.6151
R1222 B.n663 B.n100 10.6151
R1223 B.n657 B.n100 10.6151
R1224 B.n657 B.n656 10.6151
R1225 B.n656 B.n655 10.6151
R1226 B.n655 B.n102 10.6151
R1227 B.n649 B.n102 10.6151
R1228 B.n649 B.n648 10.6151
R1229 B.n648 B.n647 10.6151
R1230 B.n647 B.n104 10.6151
R1231 B.n641 B.n104 10.6151
R1232 B.n641 B.n640 10.6151
R1233 B.n640 B.n639 10.6151
R1234 B.n639 B.n106 10.6151
R1235 B.n633 B.n106 10.6151
R1236 B.n633 B.n632 10.6151
R1237 B.n632 B.n631 10.6151
R1238 B.n631 B.n108 10.6151
R1239 B.n625 B.n108 10.6151
R1240 B.n625 B.n624 10.6151
R1241 B.n624 B.n623 10.6151
R1242 B.n623 B.n110 10.6151
R1243 B.n617 B.n110 10.6151
R1244 B.n617 B.n616 10.6151
R1245 B.n616 B.n615 10.6151
R1246 B.n615 B.n112 10.6151
R1247 B.n609 B.n112 10.6151
R1248 B.n609 B.n608 10.6151
R1249 B.n608 B.n607 10.6151
R1250 B.n607 B.n114 10.6151
R1251 B.n601 B.n114 10.6151
R1252 B.n601 B.n600 10.6151
R1253 B.n600 B.n599 10.6151
R1254 B.n599 B.n116 10.6151
R1255 B.n593 B.n116 10.6151
R1256 B.n593 B.n592 10.6151
R1257 B.n483 B.n482 10.6151
R1258 B.n484 B.n483 10.6151
R1259 B.n484 B.n156 10.6151
R1260 B.n494 B.n156 10.6151
R1261 B.n495 B.n494 10.6151
R1262 B.n496 B.n495 10.6151
R1263 B.n496 B.n149 10.6151
R1264 B.n507 B.n149 10.6151
R1265 B.n508 B.n507 10.6151
R1266 B.n509 B.n508 10.6151
R1267 B.n509 B.n141 10.6151
R1268 B.n519 B.n141 10.6151
R1269 B.n520 B.n519 10.6151
R1270 B.n521 B.n520 10.6151
R1271 B.n521 B.n133 10.6151
R1272 B.n531 B.n133 10.6151
R1273 B.n532 B.n531 10.6151
R1274 B.n533 B.n532 10.6151
R1275 B.n533 B.n126 10.6151
R1276 B.n544 B.n126 10.6151
R1277 B.n545 B.n544 10.6151
R1278 B.n547 B.n545 10.6151
R1279 B.n547 B.n546 10.6151
R1280 B.n546 B.n118 10.6151
R1281 B.n558 B.n118 10.6151
R1282 B.n559 B.n558 10.6151
R1283 B.n560 B.n559 10.6151
R1284 B.n561 B.n560 10.6151
R1285 B.n563 B.n561 10.6151
R1286 B.n564 B.n563 10.6151
R1287 B.n565 B.n564 10.6151
R1288 B.n566 B.n565 10.6151
R1289 B.n568 B.n566 10.6151
R1290 B.n569 B.n568 10.6151
R1291 B.n570 B.n569 10.6151
R1292 B.n571 B.n570 10.6151
R1293 B.n573 B.n571 10.6151
R1294 B.n574 B.n573 10.6151
R1295 B.n575 B.n574 10.6151
R1296 B.n576 B.n575 10.6151
R1297 B.n578 B.n576 10.6151
R1298 B.n579 B.n578 10.6151
R1299 B.n580 B.n579 10.6151
R1300 B.n581 B.n580 10.6151
R1301 B.n583 B.n581 10.6151
R1302 B.n584 B.n583 10.6151
R1303 B.n585 B.n584 10.6151
R1304 B.n586 B.n585 10.6151
R1305 B.n588 B.n586 10.6151
R1306 B.n589 B.n588 10.6151
R1307 B.n590 B.n589 10.6151
R1308 B.n591 B.n590 10.6151
R1309 B.n477 B.n476 10.6151
R1310 B.n476 B.n168 10.6151
R1311 B.n471 B.n168 10.6151
R1312 B.n471 B.n470 10.6151
R1313 B.n470 B.n170 10.6151
R1314 B.n465 B.n170 10.6151
R1315 B.n465 B.n464 10.6151
R1316 B.n464 B.n463 10.6151
R1317 B.n463 B.n172 10.6151
R1318 B.n457 B.n172 10.6151
R1319 B.n457 B.n456 10.6151
R1320 B.n456 B.n455 10.6151
R1321 B.n455 B.n174 10.6151
R1322 B.n449 B.n174 10.6151
R1323 B.n449 B.n448 10.6151
R1324 B.n448 B.n447 10.6151
R1325 B.n447 B.n176 10.6151
R1326 B.n441 B.n176 10.6151
R1327 B.n441 B.n440 10.6151
R1328 B.n440 B.n439 10.6151
R1329 B.n439 B.n178 10.6151
R1330 B.n433 B.n178 10.6151
R1331 B.n433 B.n432 10.6151
R1332 B.n432 B.n431 10.6151
R1333 B.n431 B.n180 10.6151
R1334 B.n425 B.n180 10.6151
R1335 B.n425 B.n424 10.6151
R1336 B.n424 B.n423 10.6151
R1337 B.n423 B.n182 10.6151
R1338 B.n417 B.n182 10.6151
R1339 B.n417 B.n416 10.6151
R1340 B.n416 B.n415 10.6151
R1341 B.n415 B.n184 10.6151
R1342 B.n409 B.n184 10.6151
R1343 B.n409 B.n408 10.6151
R1344 B.n408 B.n407 10.6151
R1345 B.n407 B.n186 10.6151
R1346 B.n401 B.n186 10.6151
R1347 B.n401 B.n400 10.6151
R1348 B.n400 B.n399 10.6151
R1349 B.n399 B.n188 10.6151
R1350 B.n393 B.n188 10.6151
R1351 B.n393 B.n392 10.6151
R1352 B.n392 B.n391 10.6151
R1353 B.n391 B.n190 10.6151
R1354 B.n385 B.n190 10.6151
R1355 B.n385 B.n384 10.6151
R1356 B.n384 B.n383 10.6151
R1357 B.n383 B.n192 10.6151
R1358 B.n377 B.n192 10.6151
R1359 B.n377 B.n376 10.6151
R1360 B.n376 B.n375 10.6151
R1361 B.n375 B.n194 10.6151
R1362 B.n369 B.n194 10.6151
R1363 B.n369 B.n368 10.6151
R1364 B.n368 B.n367 10.6151
R1365 B.n363 B.n362 10.6151
R1366 B.n362 B.n200 10.6151
R1367 B.n357 B.n200 10.6151
R1368 B.n357 B.n356 10.6151
R1369 B.n356 B.n355 10.6151
R1370 B.n355 B.n202 10.6151
R1371 B.n349 B.n202 10.6151
R1372 B.n349 B.n348 10.6151
R1373 B.n346 B.n206 10.6151
R1374 B.n340 B.n206 10.6151
R1375 B.n340 B.n339 10.6151
R1376 B.n339 B.n338 10.6151
R1377 B.n338 B.n208 10.6151
R1378 B.n332 B.n208 10.6151
R1379 B.n332 B.n331 10.6151
R1380 B.n331 B.n330 10.6151
R1381 B.n330 B.n210 10.6151
R1382 B.n324 B.n210 10.6151
R1383 B.n324 B.n323 10.6151
R1384 B.n323 B.n322 10.6151
R1385 B.n322 B.n212 10.6151
R1386 B.n316 B.n212 10.6151
R1387 B.n316 B.n315 10.6151
R1388 B.n315 B.n314 10.6151
R1389 B.n314 B.n214 10.6151
R1390 B.n308 B.n214 10.6151
R1391 B.n308 B.n307 10.6151
R1392 B.n307 B.n306 10.6151
R1393 B.n306 B.n216 10.6151
R1394 B.n300 B.n216 10.6151
R1395 B.n300 B.n299 10.6151
R1396 B.n299 B.n298 10.6151
R1397 B.n298 B.n218 10.6151
R1398 B.n292 B.n218 10.6151
R1399 B.n292 B.n291 10.6151
R1400 B.n291 B.n290 10.6151
R1401 B.n290 B.n220 10.6151
R1402 B.n284 B.n220 10.6151
R1403 B.n284 B.n283 10.6151
R1404 B.n283 B.n282 10.6151
R1405 B.n282 B.n222 10.6151
R1406 B.n276 B.n222 10.6151
R1407 B.n276 B.n275 10.6151
R1408 B.n275 B.n274 10.6151
R1409 B.n274 B.n224 10.6151
R1410 B.n268 B.n224 10.6151
R1411 B.n268 B.n267 10.6151
R1412 B.n267 B.n266 10.6151
R1413 B.n266 B.n226 10.6151
R1414 B.n260 B.n226 10.6151
R1415 B.n260 B.n259 10.6151
R1416 B.n259 B.n258 10.6151
R1417 B.n258 B.n228 10.6151
R1418 B.n252 B.n228 10.6151
R1419 B.n252 B.n251 10.6151
R1420 B.n251 B.n250 10.6151
R1421 B.n250 B.n230 10.6151
R1422 B.n244 B.n230 10.6151
R1423 B.n244 B.n243 10.6151
R1424 B.n243 B.n242 10.6151
R1425 B.n242 B.n232 10.6151
R1426 B.n236 B.n232 10.6151
R1427 B.n236 B.n235 10.6151
R1428 B.n235 B.n164 10.6151
R1429 B.n478 B.n160 10.6151
R1430 B.n488 B.n160 10.6151
R1431 B.n489 B.n488 10.6151
R1432 B.n490 B.n489 10.6151
R1433 B.n490 B.n152 10.6151
R1434 B.n501 B.n152 10.6151
R1435 B.n502 B.n501 10.6151
R1436 B.n503 B.n502 10.6151
R1437 B.n503 B.n145 10.6151
R1438 B.n513 B.n145 10.6151
R1439 B.n514 B.n513 10.6151
R1440 B.n515 B.n514 10.6151
R1441 B.n515 B.n137 10.6151
R1442 B.n525 B.n137 10.6151
R1443 B.n526 B.n525 10.6151
R1444 B.n527 B.n526 10.6151
R1445 B.n527 B.n129 10.6151
R1446 B.n538 B.n129 10.6151
R1447 B.n539 B.n538 10.6151
R1448 B.n540 B.n539 10.6151
R1449 B.n540 B.n122 10.6151
R1450 B.n551 B.n122 10.6151
R1451 B.n552 B.n551 10.6151
R1452 B.n553 B.n552 10.6151
R1453 B.n553 B.n0 10.6151
R1454 B.n886 B.n1 10.6151
R1455 B.n886 B.n885 10.6151
R1456 B.n885 B.n884 10.6151
R1457 B.n884 B.n10 10.6151
R1458 B.n878 B.n10 10.6151
R1459 B.n878 B.n877 10.6151
R1460 B.n877 B.n876 10.6151
R1461 B.n876 B.n16 10.6151
R1462 B.n870 B.n16 10.6151
R1463 B.n870 B.n869 10.6151
R1464 B.n869 B.n868 10.6151
R1465 B.n868 B.n24 10.6151
R1466 B.n862 B.n24 10.6151
R1467 B.n862 B.n861 10.6151
R1468 B.n861 B.n860 10.6151
R1469 B.n860 B.n31 10.6151
R1470 B.n854 B.n31 10.6151
R1471 B.n854 B.n853 10.6151
R1472 B.n853 B.n852 10.6151
R1473 B.n852 B.n37 10.6151
R1474 B.n846 B.n37 10.6151
R1475 B.n846 B.n845 10.6151
R1476 B.n845 B.n844 10.6151
R1477 B.n844 B.n45 10.6151
R1478 B.n838 B.n45 10.6151
R1479 B.n724 B.n723 6.5566
R1480 B.n707 B.n88 6.5566
R1481 B.n363 B.n198 6.5566
R1482 B.n348 B.n347 6.5566
R1483 B.n725 B.n724 4.05904
R1484 B.n703 B.n88 4.05904
R1485 B.n367 B.n198 4.05904
R1486 B.n347 B.n346 4.05904
R1487 B.n542 B.t0 3.93522
R1488 B.n880 B.t1 3.93522
R1489 B.n892 B.n0 2.81026
R1490 B.n892 B.n1 2.81026
R1491 VP.n0 VP.t1 240.298
R1492 VP.n0 VP.t0 191.413
R1493 VP VP.n0 0.431811
R1494 VTAIL.n1 VTAIL.t0 43.8242
R1495 VTAIL.n3 VTAIL.t1 43.8241
R1496 VTAIL.n0 VTAIL.t3 43.8241
R1497 VTAIL.n2 VTAIL.t2 43.8241
R1498 VTAIL.n1 VTAIL.n0 32.3927
R1499 VTAIL.n3 VTAIL.n2 29.7462
R1500 VTAIL.n2 VTAIL.n1 1.7936
R1501 VTAIL VTAIL.n0 1.19016
R1502 VTAIL VTAIL.n3 0.603948
R1503 VDD1 VDD1.t1 105.374
R1504 VDD1 VDD1.t0 61.2227
R1505 VN VN.t0 240.299
R1506 VN VN.t1 191.845
R1507 VDD2.n0 VDD2.t0 104.189
R1508 VDD2.n0 VDD2.t1 60.5029
R1509 VDD2 VDD2.n0 0.720328
C0 VDD2 VP 0.339334f
C1 VDD2 VTAIL 6.47053f
C2 VTAIL VP 3.34754f
C3 VDD2 VN 3.88473f
C4 VN VP 6.46655f
C5 VDD2 VDD1 0.692077f
C6 VDD1 VP 4.07256f
C7 VN VTAIL 3.33319f
C8 VTAIL VDD1 6.41995f
C9 VN VDD1 0.148186f
C10 VDD2 B 5.392844f
C11 VDD1 B 8.90967f
C12 VTAIL B 9.47753f
C13 VN B 12.08363f
C14 VP B 6.923559f
C15 VDD2.t0 B 3.8514f
C16 VDD2.t1 B 3.14455f
C17 VDD2.n0 B 3.2714f
C18 VN.t1 B 4.00609f
C19 VN.t0 B 4.5774f
C20 VDD1.t0 B 3.15561f
C21 VDD1.t1 B 3.90202f
C22 VTAIL.t3 B 3.02143f
C23 VTAIL.n0 B 1.89951f
C24 VTAIL.t0 B 3.02144f
C25 VTAIL.n1 B 1.938f
C26 VTAIL.t2 B 3.02142f
C27 VTAIL.n2 B 1.76913f
C28 VTAIL.t1 B 3.02143f
C29 VTAIL.n3 B 1.69321f
C30 VP.t0 B 4.07358f
C31 VP.t1 B 4.65656f
C32 VP.n0 B 5.09096f
.ends

