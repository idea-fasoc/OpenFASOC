* NGSPICE file created from diff_pair_sample_0513.ext - technology: sky130A

.subckt diff_pair_sample_0513 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X1 VTAIL.t18 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X2 VDD1.t9 VP.t0 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X3 VDD2.t7 VN.t2 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=1.2243 ps=7.75 w=7.42 l=2.37
X4 VDD1.t8 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=2.8938 ps=15.62 w=7.42 l=2.37
X5 VDD2.t6 VN.t3 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X6 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=0 ps=0 w=7.42 l=2.37
X7 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X8 VTAIL.t15 VN.t4 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X9 VTAIL.t0 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X10 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=0 ps=0 w=7.42 l=2.37
X11 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=1.2243 ps=7.75 w=7.42 l=2.37
X12 VDD1.t4 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=1.2243 ps=7.75 w=7.42 l=2.37
X13 VDD2.t9 VN.t5 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=2.8938 ps=15.62 w=7.42 l=2.37
X14 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=0 ps=0 w=7.42 l=2.37
X15 VDD2.t2 VN.t6 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=2.8938 ps=15.62 w=7.42 l=2.37
X16 VTAIL.t8 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X17 VTAIL.t12 VN.t7 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X18 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=2.8938 ps=15.62 w=7.42 l=2.37
X19 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X20 VDD2.t4 VN.t8 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=1.2243 ps=7.75 w=7.42 l=2.37
X21 VTAIL.t6 VP.t9 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X22 VDD2.t5 VN.t9 VTAIL.t10 B.t23 sky130_fd_pr__nfet_01v8 ad=1.2243 pd=7.75 as=1.2243 ps=7.75 w=7.42 l=2.37
X23 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.8938 pd=15.62 as=0 ps=0 w=7.42 l=2.37
R0 VN.n73 VN.n38 161.3
R1 VN.n72 VN.n71 161.3
R2 VN.n70 VN.n39 161.3
R3 VN.n69 VN.n68 161.3
R4 VN.n67 VN.n40 161.3
R5 VN.n66 VN.n65 161.3
R6 VN.n64 VN.n63 161.3
R7 VN.n62 VN.n42 161.3
R8 VN.n61 VN.n60 161.3
R9 VN.n59 VN.n43 161.3
R10 VN.n58 VN.n57 161.3
R11 VN.n55 VN.n44 161.3
R12 VN.n54 VN.n53 161.3
R13 VN.n52 VN.n45 161.3
R14 VN.n51 VN.n50 161.3
R15 VN.n49 VN.n46 161.3
R16 VN.n35 VN.n0 161.3
R17 VN.n34 VN.n33 161.3
R18 VN.n32 VN.n1 161.3
R19 VN.n31 VN.n30 161.3
R20 VN.n29 VN.n2 161.3
R21 VN.n28 VN.n27 161.3
R22 VN.n26 VN.n25 161.3
R23 VN.n24 VN.n4 161.3
R24 VN.n23 VN.n22 161.3
R25 VN.n21 VN.n5 161.3
R26 VN.n20 VN.n19 161.3
R27 VN.n17 VN.n6 161.3
R28 VN.n16 VN.n15 161.3
R29 VN.n14 VN.n7 161.3
R30 VN.n13 VN.n12 161.3
R31 VN.n11 VN.n8 161.3
R32 VN.n9 VN.t2 108.352
R33 VN.n47 VN.t5 108.352
R34 VN.n37 VN.n36 103.531
R35 VN.n75 VN.n74 103.531
R36 VN.n10 VN.t7 75.4528
R37 VN.n18 VN.t3 75.4528
R38 VN.n3 VN.t1 75.4528
R39 VN.n36 VN.t6 75.4528
R40 VN.n48 VN.t0 75.4528
R41 VN.n56 VN.t9 75.4528
R42 VN.n41 VN.t4 75.4528
R43 VN.n74 VN.t8 75.4528
R44 VN.n30 VN.n1 56.5617
R45 VN.n68 VN.n39 56.5617
R46 VN.n10 VN.n9 50.3824
R47 VN.n48 VN.n47 50.3824
R48 VN.n12 VN.n7 50.2647
R49 VN.n24 VN.n23 50.2647
R50 VN.n50 VN.n45 50.2647
R51 VN.n62 VN.n61 50.2647
R52 VN VN.n75 48.5967
R53 VN.n16 VN.n7 30.8893
R54 VN.n23 VN.n5 30.8893
R55 VN.n54 VN.n45 30.8893
R56 VN.n61 VN.n43 30.8893
R57 VN.n12 VN.n11 24.5923
R58 VN.n17 VN.n16 24.5923
R59 VN.n19 VN.n5 24.5923
R60 VN.n25 VN.n24 24.5923
R61 VN.n29 VN.n28 24.5923
R62 VN.n30 VN.n29 24.5923
R63 VN.n34 VN.n1 24.5923
R64 VN.n35 VN.n34 24.5923
R65 VN.n50 VN.n49 24.5923
R66 VN.n57 VN.n43 24.5923
R67 VN.n55 VN.n54 24.5923
R68 VN.n68 VN.n67 24.5923
R69 VN.n67 VN.n66 24.5923
R70 VN.n63 VN.n62 24.5923
R71 VN.n73 VN.n72 24.5923
R72 VN.n72 VN.n39 24.5923
R73 VN.n11 VN.n10 22.1332
R74 VN.n25 VN.n3 22.1332
R75 VN.n49 VN.n48 22.1332
R76 VN.n63 VN.n41 22.1332
R77 VN.n18 VN.n17 12.2964
R78 VN.n19 VN.n18 12.2964
R79 VN.n57 VN.n56 12.2964
R80 VN.n56 VN.n55 12.2964
R81 VN.n36 VN.n35 7.37805
R82 VN.n74 VN.n73 7.37805
R83 VN.n47 VN.n46 6.9978
R84 VN.n9 VN.n8 6.9978
R85 VN.n28 VN.n3 2.45968
R86 VN.n66 VN.n41 2.45968
R87 VN.n75 VN.n38 0.278335
R88 VN.n37 VN.n0 0.278335
R89 VN.n71 VN.n38 0.189894
R90 VN.n71 VN.n70 0.189894
R91 VN.n70 VN.n69 0.189894
R92 VN.n69 VN.n40 0.189894
R93 VN.n65 VN.n40 0.189894
R94 VN.n65 VN.n64 0.189894
R95 VN.n64 VN.n42 0.189894
R96 VN.n60 VN.n42 0.189894
R97 VN.n60 VN.n59 0.189894
R98 VN.n59 VN.n58 0.189894
R99 VN.n58 VN.n44 0.189894
R100 VN.n53 VN.n44 0.189894
R101 VN.n53 VN.n52 0.189894
R102 VN.n52 VN.n51 0.189894
R103 VN.n51 VN.n46 0.189894
R104 VN.n13 VN.n8 0.189894
R105 VN.n14 VN.n13 0.189894
R106 VN.n15 VN.n14 0.189894
R107 VN.n15 VN.n6 0.189894
R108 VN.n20 VN.n6 0.189894
R109 VN.n21 VN.n20 0.189894
R110 VN.n22 VN.n21 0.189894
R111 VN.n22 VN.n4 0.189894
R112 VN.n26 VN.n4 0.189894
R113 VN.n27 VN.n26 0.189894
R114 VN.n27 VN.n2 0.189894
R115 VN.n31 VN.n2 0.189894
R116 VN.n32 VN.n31 0.189894
R117 VN.n33 VN.n32 0.189894
R118 VN.n33 VN.n0 0.189894
R119 VN VN.n37 0.153485
R120 VDD2.n77 VDD2.n43 289.615
R121 VDD2.n34 VDD2.n0 289.615
R122 VDD2.n78 VDD2.n77 185
R123 VDD2.n76 VDD2.n75 185
R124 VDD2.n47 VDD2.n46 185
R125 VDD2.n70 VDD2.n69 185
R126 VDD2.n68 VDD2.n67 185
R127 VDD2.n51 VDD2.n50 185
R128 VDD2.n62 VDD2.n61 185
R129 VDD2.n60 VDD2.n59 185
R130 VDD2.n55 VDD2.n54 185
R131 VDD2.n12 VDD2.n11 185
R132 VDD2.n17 VDD2.n16 185
R133 VDD2.n19 VDD2.n18 185
R134 VDD2.n8 VDD2.n7 185
R135 VDD2.n25 VDD2.n24 185
R136 VDD2.n27 VDD2.n26 185
R137 VDD2.n4 VDD2.n3 185
R138 VDD2.n33 VDD2.n32 185
R139 VDD2.n35 VDD2.n34 185
R140 VDD2.n56 VDD2.t4 147.659
R141 VDD2.n13 VDD2.t7 147.659
R142 VDD2.n77 VDD2.n76 104.615
R143 VDD2.n76 VDD2.n46 104.615
R144 VDD2.n69 VDD2.n46 104.615
R145 VDD2.n69 VDD2.n68 104.615
R146 VDD2.n68 VDD2.n50 104.615
R147 VDD2.n61 VDD2.n50 104.615
R148 VDD2.n61 VDD2.n60 104.615
R149 VDD2.n60 VDD2.n54 104.615
R150 VDD2.n17 VDD2.n11 104.615
R151 VDD2.n18 VDD2.n17 104.615
R152 VDD2.n18 VDD2.n7 104.615
R153 VDD2.n25 VDD2.n7 104.615
R154 VDD2.n26 VDD2.n25 104.615
R155 VDD2.n26 VDD2.n3 104.615
R156 VDD2.n33 VDD2.n3 104.615
R157 VDD2.n34 VDD2.n33 104.615
R158 VDD2.n42 VDD2.n41 66.5028
R159 VDD2 VDD2.n85 66.5
R160 VDD2.n84 VDD2.n83 64.8126
R161 VDD2.n40 VDD2.n39 64.8125
R162 VDD2.t4 VDD2.n54 52.3082
R163 VDD2.t7 VDD2.n11 52.3082
R164 VDD2.n40 VDD2.n38 50.8038
R165 VDD2.n82 VDD2.n81 48.4763
R166 VDD2.n82 VDD2.n42 41.1679
R167 VDD2.n56 VDD2.n55 15.6677
R168 VDD2.n13 VDD2.n12 15.6677
R169 VDD2.n59 VDD2.n58 12.8005
R170 VDD2.n16 VDD2.n15 12.8005
R171 VDD2.n62 VDD2.n53 12.0247
R172 VDD2.n19 VDD2.n10 12.0247
R173 VDD2.n63 VDD2.n51 11.249
R174 VDD2.n20 VDD2.n8 11.249
R175 VDD2.n67 VDD2.n66 10.4732
R176 VDD2.n24 VDD2.n23 10.4732
R177 VDD2.n70 VDD2.n49 9.69747
R178 VDD2.n27 VDD2.n6 9.69747
R179 VDD2.n81 VDD2.n80 9.45567
R180 VDD2.n38 VDD2.n37 9.45567
R181 VDD2.n80 VDD2.n79 9.3005
R182 VDD2.n45 VDD2.n44 9.3005
R183 VDD2.n74 VDD2.n73 9.3005
R184 VDD2.n72 VDD2.n71 9.3005
R185 VDD2.n49 VDD2.n48 9.3005
R186 VDD2.n66 VDD2.n65 9.3005
R187 VDD2.n64 VDD2.n63 9.3005
R188 VDD2.n53 VDD2.n52 9.3005
R189 VDD2.n58 VDD2.n57 9.3005
R190 VDD2.n37 VDD2.n36 9.3005
R191 VDD2.n31 VDD2.n30 9.3005
R192 VDD2.n29 VDD2.n28 9.3005
R193 VDD2.n6 VDD2.n5 9.3005
R194 VDD2.n23 VDD2.n22 9.3005
R195 VDD2.n21 VDD2.n20 9.3005
R196 VDD2.n10 VDD2.n9 9.3005
R197 VDD2.n15 VDD2.n14 9.3005
R198 VDD2.n2 VDD2.n1 9.3005
R199 VDD2.n71 VDD2.n47 8.92171
R200 VDD2.n28 VDD2.n4 8.92171
R201 VDD2.n75 VDD2.n74 8.14595
R202 VDD2.n32 VDD2.n31 8.14595
R203 VDD2.n81 VDD2.n43 7.3702
R204 VDD2.n78 VDD2.n45 7.3702
R205 VDD2.n35 VDD2.n2 7.3702
R206 VDD2.n38 VDD2.n0 7.3702
R207 VDD2.n79 VDD2.n43 6.59444
R208 VDD2.n79 VDD2.n78 6.59444
R209 VDD2.n36 VDD2.n35 6.59444
R210 VDD2.n36 VDD2.n0 6.59444
R211 VDD2.n75 VDD2.n45 5.81868
R212 VDD2.n32 VDD2.n2 5.81868
R213 VDD2.n74 VDD2.n47 5.04292
R214 VDD2.n31 VDD2.n4 5.04292
R215 VDD2.n57 VDD2.n56 4.38565
R216 VDD2.n14 VDD2.n13 4.38565
R217 VDD2.n71 VDD2.n70 4.26717
R218 VDD2.n28 VDD2.n27 4.26717
R219 VDD2.n67 VDD2.n49 3.49141
R220 VDD2.n24 VDD2.n6 3.49141
R221 VDD2.n66 VDD2.n51 2.71565
R222 VDD2.n23 VDD2.n8 2.71565
R223 VDD2.n85 VDD2.t1 2.66896
R224 VDD2.n85 VDD2.t9 2.66896
R225 VDD2.n83 VDD2.t0 2.66896
R226 VDD2.n83 VDD2.t5 2.66896
R227 VDD2.n41 VDD2.t8 2.66896
R228 VDD2.n41 VDD2.t2 2.66896
R229 VDD2.n39 VDD2.t3 2.66896
R230 VDD2.n39 VDD2.t6 2.66896
R231 VDD2.n84 VDD2.n82 2.32809
R232 VDD2.n63 VDD2.n62 1.93989
R233 VDD2.n20 VDD2.n19 1.93989
R234 VDD2.n59 VDD2.n53 1.16414
R235 VDD2.n16 VDD2.n10 1.16414
R236 VDD2 VDD2.n84 0.640586
R237 VDD2.n42 VDD2.n40 0.527051
R238 VDD2.n58 VDD2.n55 0.388379
R239 VDD2.n15 VDD2.n12 0.388379
R240 VDD2.n80 VDD2.n44 0.155672
R241 VDD2.n73 VDD2.n44 0.155672
R242 VDD2.n73 VDD2.n72 0.155672
R243 VDD2.n72 VDD2.n48 0.155672
R244 VDD2.n65 VDD2.n48 0.155672
R245 VDD2.n65 VDD2.n64 0.155672
R246 VDD2.n64 VDD2.n52 0.155672
R247 VDD2.n57 VDD2.n52 0.155672
R248 VDD2.n14 VDD2.n9 0.155672
R249 VDD2.n21 VDD2.n9 0.155672
R250 VDD2.n22 VDD2.n21 0.155672
R251 VDD2.n22 VDD2.n5 0.155672
R252 VDD2.n29 VDD2.n5 0.155672
R253 VDD2.n30 VDD2.n29 0.155672
R254 VDD2.n30 VDD2.n1 0.155672
R255 VDD2.n37 VDD2.n1 0.155672
R256 VTAIL.n168 VTAIL.n134 289.615
R257 VTAIL.n36 VTAIL.n2 289.615
R258 VTAIL.n128 VTAIL.n94 289.615
R259 VTAIL.n84 VTAIL.n50 289.615
R260 VTAIL.n146 VTAIL.n145 185
R261 VTAIL.n151 VTAIL.n150 185
R262 VTAIL.n153 VTAIL.n152 185
R263 VTAIL.n142 VTAIL.n141 185
R264 VTAIL.n159 VTAIL.n158 185
R265 VTAIL.n161 VTAIL.n160 185
R266 VTAIL.n138 VTAIL.n137 185
R267 VTAIL.n167 VTAIL.n166 185
R268 VTAIL.n169 VTAIL.n168 185
R269 VTAIL.n14 VTAIL.n13 185
R270 VTAIL.n19 VTAIL.n18 185
R271 VTAIL.n21 VTAIL.n20 185
R272 VTAIL.n10 VTAIL.n9 185
R273 VTAIL.n27 VTAIL.n26 185
R274 VTAIL.n29 VTAIL.n28 185
R275 VTAIL.n6 VTAIL.n5 185
R276 VTAIL.n35 VTAIL.n34 185
R277 VTAIL.n37 VTAIL.n36 185
R278 VTAIL.n129 VTAIL.n128 185
R279 VTAIL.n127 VTAIL.n126 185
R280 VTAIL.n98 VTAIL.n97 185
R281 VTAIL.n121 VTAIL.n120 185
R282 VTAIL.n119 VTAIL.n118 185
R283 VTAIL.n102 VTAIL.n101 185
R284 VTAIL.n113 VTAIL.n112 185
R285 VTAIL.n111 VTAIL.n110 185
R286 VTAIL.n106 VTAIL.n105 185
R287 VTAIL.n85 VTAIL.n84 185
R288 VTAIL.n83 VTAIL.n82 185
R289 VTAIL.n54 VTAIL.n53 185
R290 VTAIL.n77 VTAIL.n76 185
R291 VTAIL.n75 VTAIL.n74 185
R292 VTAIL.n58 VTAIL.n57 185
R293 VTAIL.n69 VTAIL.n68 185
R294 VTAIL.n67 VTAIL.n66 185
R295 VTAIL.n62 VTAIL.n61 185
R296 VTAIL.n147 VTAIL.t13 147.659
R297 VTAIL.n15 VTAIL.t7 147.659
R298 VTAIL.n107 VTAIL.t3 147.659
R299 VTAIL.n63 VTAIL.t14 147.659
R300 VTAIL.n151 VTAIL.n145 104.615
R301 VTAIL.n152 VTAIL.n151 104.615
R302 VTAIL.n152 VTAIL.n141 104.615
R303 VTAIL.n159 VTAIL.n141 104.615
R304 VTAIL.n160 VTAIL.n159 104.615
R305 VTAIL.n160 VTAIL.n137 104.615
R306 VTAIL.n167 VTAIL.n137 104.615
R307 VTAIL.n168 VTAIL.n167 104.615
R308 VTAIL.n19 VTAIL.n13 104.615
R309 VTAIL.n20 VTAIL.n19 104.615
R310 VTAIL.n20 VTAIL.n9 104.615
R311 VTAIL.n27 VTAIL.n9 104.615
R312 VTAIL.n28 VTAIL.n27 104.615
R313 VTAIL.n28 VTAIL.n5 104.615
R314 VTAIL.n35 VTAIL.n5 104.615
R315 VTAIL.n36 VTAIL.n35 104.615
R316 VTAIL.n128 VTAIL.n127 104.615
R317 VTAIL.n127 VTAIL.n97 104.615
R318 VTAIL.n120 VTAIL.n97 104.615
R319 VTAIL.n120 VTAIL.n119 104.615
R320 VTAIL.n119 VTAIL.n101 104.615
R321 VTAIL.n112 VTAIL.n101 104.615
R322 VTAIL.n112 VTAIL.n111 104.615
R323 VTAIL.n111 VTAIL.n105 104.615
R324 VTAIL.n84 VTAIL.n83 104.615
R325 VTAIL.n83 VTAIL.n53 104.615
R326 VTAIL.n76 VTAIL.n53 104.615
R327 VTAIL.n76 VTAIL.n75 104.615
R328 VTAIL.n75 VTAIL.n57 104.615
R329 VTAIL.n68 VTAIL.n57 104.615
R330 VTAIL.n68 VTAIL.n67 104.615
R331 VTAIL.n67 VTAIL.n61 104.615
R332 VTAIL.t13 VTAIL.n145 52.3082
R333 VTAIL.t7 VTAIL.n13 52.3082
R334 VTAIL.t3 VTAIL.n105 52.3082
R335 VTAIL.t14 VTAIL.n61 52.3082
R336 VTAIL.n93 VTAIL.n92 48.1338
R337 VTAIL.n91 VTAIL.n90 48.1338
R338 VTAIL.n49 VTAIL.n48 48.1338
R339 VTAIL.n47 VTAIL.n46 48.1338
R340 VTAIL.n175 VTAIL.n174 48.1337
R341 VTAIL.n1 VTAIL.n0 48.1337
R342 VTAIL.n43 VTAIL.n42 48.1337
R343 VTAIL.n45 VTAIL.n44 48.1337
R344 VTAIL.n173 VTAIL.n172 31.7975
R345 VTAIL.n41 VTAIL.n40 31.7975
R346 VTAIL.n133 VTAIL.n132 31.7975
R347 VTAIL.n89 VTAIL.n88 31.7975
R348 VTAIL.n47 VTAIL.n45 23.4186
R349 VTAIL.n173 VTAIL.n133 21.091
R350 VTAIL.n147 VTAIL.n146 15.6677
R351 VTAIL.n15 VTAIL.n14 15.6677
R352 VTAIL.n107 VTAIL.n106 15.6677
R353 VTAIL.n63 VTAIL.n62 15.6677
R354 VTAIL.n150 VTAIL.n149 12.8005
R355 VTAIL.n18 VTAIL.n17 12.8005
R356 VTAIL.n110 VTAIL.n109 12.8005
R357 VTAIL.n66 VTAIL.n65 12.8005
R358 VTAIL.n153 VTAIL.n144 12.0247
R359 VTAIL.n21 VTAIL.n12 12.0247
R360 VTAIL.n113 VTAIL.n104 12.0247
R361 VTAIL.n69 VTAIL.n60 12.0247
R362 VTAIL.n154 VTAIL.n142 11.249
R363 VTAIL.n22 VTAIL.n10 11.249
R364 VTAIL.n114 VTAIL.n102 11.249
R365 VTAIL.n70 VTAIL.n58 11.249
R366 VTAIL.n158 VTAIL.n157 10.4732
R367 VTAIL.n26 VTAIL.n25 10.4732
R368 VTAIL.n118 VTAIL.n117 10.4732
R369 VTAIL.n74 VTAIL.n73 10.4732
R370 VTAIL.n161 VTAIL.n140 9.69747
R371 VTAIL.n29 VTAIL.n8 9.69747
R372 VTAIL.n121 VTAIL.n100 9.69747
R373 VTAIL.n77 VTAIL.n56 9.69747
R374 VTAIL.n172 VTAIL.n171 9.45567
R375 VTAIL.n40 VTAIL.n39 9.45567
R376 VTAIL.n132 VTAIL.n131 9.45567
R377 VTAIL.n88 VTAIL.n87 9.45567
R378 VTAIL.n171 VTAIL.n170 9.3005
R379 VTAIL.n165 VTAIL.n164 9.3005
R380 VTAIL.n163 VTAIL.n162 9.3005
R381 VTAIL.n140 VTAIL.n139 9.3005
R382 VTAIL.n157 VTAIL.n156 9.3005
R383 VTAIL.n155 VTAIL.n154 9.3005
R384 VTAIL.n144 VTAIL.n143 9.3005
R385 VTAIL.n149 VTAIL.n148 9.3005
R386 VTAIL.n136 VTAIL.n135 9.3005
R387 VTAIL.n39 VTAIL.n38 9.3005
R388 VTAIL.n33 VTAIL.n32 9.3005
R389 VTAIL.n31 VTAIL.n30 9.3005
R390 VTAIL.n8 VTAIL.n7 9.3005
R391 VTAIL.n25 VTAIL.n24 9.3005
R392 VTAIL.n23 VTAIL.n22 9.3005
R393 VTAIL.n12 VTAIL.n11 9.3005
R394 VTAIL.n17 VTAIL.n16 9.3005
R395 VTAIL.n4 VTAIL.n3 9.3005
R396 VTAIL.n131 VTAIL.n130 9.3005
R397 VTAIL.n96 VTAIL.n95 9.3005
R398 VTAIL.n125 VTAIL.n124 9.3005
R399 VTAIL.n123 VTAIL.n122 9.3005
R400 VTAIL.n100 VTAIL.n99 9.3005
R401 VTAIL.n117 VTAIL.n116 9.3005
R402 VTAIL.n115 VTAIL.n114 9.3005
R403 VTAIL.n104 VTAIL.n103 9.3005
R404 VTAIL.n109 VTAIL.n108 9.3005
R405 VTAIL.n87 VTAIL.n86 9.3005
R406 VTAIL.n52 VTAIL.n51 9.3005
R407 VTAIL.n81 VTAIL.n80 9.3005
R408 VTAIL.n79 VTAIL.n78 9.3005
R409 VTAIL.n56 VTAIL.n55 9.3005
R410 VTAIL.n73 VTAIL.n72 9.3005
R411 VTAIL.n71 VTAIL.n70 9.3005
R412 VTAIL.n60 VTAIL.n59 9.3005
R413 VTAIL.n65 VTAIL.n64 9.3005
R414 VTAIL.n162 VTAIL.n138 8.92171
R415 VTAIL.n30 VTAIL.n6 8.92171
R416 VTAIL.n122 VTAIL.n98 8.92171
R417 VTAIL.n78 VTAIL.n54 8.92171
R418 VTAIL.n166 VTAIL.n165 8.14595
R419 VTAIL.n34 VTAIL.n33 8.14595
R420 VTAIL.n126 VTAIL.n125 8.14595
R421 VTAIL.n82 VTAIL.n81 8.14595
R422 VTAIL.n169 VTAIL.n136 7.3702
R423 VTAIL.n172 VTAIL.n134 7.3702
R424 VTAIL.n37 VTAIL.n4 7.3702
R425 VTAIL.n40 VTAIL.n2 7.3702
R426 VTAIL.n132 VTAIL.n94 7.3702
R427 VTAIL.n129 VTAIL.n96 7.3702
R428 VTAIL.n88 VTAIL.n50 7.3702
R429 VTAIL.n85 VTAIL.n52 7.3702
R430 VTAIL.n170 VTAIL.n169 6.59444
R431 VTAIL.n170 VTAIL.n134 6.59444
R432 VTAIL.n38 VTAIL.n37 6.59444
R433 VTAIL.n38 VTAIL.n2 6.59444
R434 VTAIL.n130 VTAIL.n94 6.59444
R435 VTAIL.n130 VTAIL.n129 6.59444
R436 VTAIL.n86 VTAIL.n50 6.59444
R437 VTAIL.n86 VTAIL.n85 6.59444
R438 VTAIL.n166 VTAIL.n136 5.81868
R439 VTAIL.n34 VTAIL.n4 5.81868
R440 VTAIL.n126 VTAIL.n96 5.81868
R441 VTAIL.n82 VTAIL.n52 5.81868
R442 VTAIL.n165 VTAIL.n138 5.04292
R443 VTAIL.n33 VTAIL.n6 5.04292
R444 VTAIL.n125 VTAIL.n98 5.04292
R445 VTAIL.n81 VTAIL.n54 5.04292
R446 VTAIL.n108 VTAIL.n107 4.38565
R447 VTAIL.n64 VTAIL.n63 4.38565
R448 VTAIL.n148 VTAIL.n147 4.38565
R449 VTAIL.n16 VTAIL.n15 4.38565
R450 VTAIL.n162 VTAIL.n161 4.26717
R451 VTAIL.n30 VTAIL.n29 4.26717
R452 VTAIL.n122 VTAIL.n121 4.26717
R453 VTAIL.n78 VTAIL.n77 4.26717
R454 VTAIL.n158 VTAIL.n140 3.49141
R455 VTAIL.n26 VTAIL.n8 3.49141
R456 VTAIL.n118 VTAIL.n100 3.49141
R457 VTAIL.n74 VTAIL.n56 3.49141
R458 VTAIL.n157 VTAIL.n142 2.71565
R459 VTAIL.n25 VTAIL.n10 2.71565
R460 VTAIL.n117 VTAIL.n102 2.71565
R461 VTAIL.n73 VTAIL.n58 2.71565
R462 VTAIL.n174 VTAIL.t16 2.66896
R463 VTAIL.n174 VTAIL.t18 2.66896
R464 VTAIL.n0 VTAIL.t17 2.66896
R465 VTAIL.n0 VTAIL.t12 2.66896
R466 VTAIL.n42 VTAIL.t9 2.66896
R467 VTAIL.n42 VTAIL.t0 2.66896
R468 VTAIL.n44 VTAIL.t5 2.66896
R469 VTAIL.n44 VTAIL.t8 2.66896
R470 VTAIL.n92 VTAIL.t2 2.66896
R471 VTAIL.n92 VTAIL.t1 2.66896
R472 VTAIL.n90 VTAIL.t4 2.66896
R473 VTAIL.n90 VTAIL.t6 2.66896
R474 VTAIL.n48 VTAIL.t10 2.66896
R475 VTAIL.n48 VTAIL.t19 2.66896
R476 VTAIL.n46 VTAIL.t11 2.66896
R477 VTAIL.n46 VTAIL.t15 2.66896
R478 VTAIL.n49 VTAIL.n47 2.32809
R479 VTAIL.n89 VTAIL.n49 2.32809
R480 VTAIL.n93 VTAIL.n91 2.32809
R481 VTAIL.n133 VTAIL.n93 2.32809
R482 VTAIL.n45 VTAIL.n43 2.32809
R483 VTAIL.n43 VTAIL.n41 2.32809
R484 VTAIL.n175 VTAIL.n173 2.32809
R485 VTAIL.n154 VTAIL.n153 1.93989
R486 VTAIL.n22 VTAIL.n21 1.93989
R487 VTAIL.n114 VTAIL.n113 1.93989
R488 VTAIL.n70 VTAIL.n69 1.93989
R489 VTAIL VTAIL.n1 1.80438
R490 VTAIL.n91 VTAIL.n89 1.63412
R491 VTAIL.n41 VTAIL.n1 1.63412
R492 VTAIL.n150 VTAIL.n144 1.16414
R493 VTAIL.n18 VTAIL.n12 1.16414
R494 VTAIL.n110 VTAIL.n104 1.16414
R495 VTAIL.n66 VTAIL.n60 1.16414
R496 VTAIL VTAIL.n175 0.524207
R497 VTAIL.n149 VTAIL.n146 0.388379
R498 VTAIL.n17 VTAIL.n14 0.388379
R499 VTAIL.n109 VTAIL.n106 0.388379
R500 VTAIL.n65 VTAIL.n62 0.388379
R501 VTAIL.n148 VTAIL.n143 0.155672
R502 VTAIL.n155 VTAIL.n143 0.155672
R503 VTAIL.n156 VTAIL.n155 0.155672
R504 VTAIL.n156 VTAIL.n139 0.155672
R505 VTAIL.n163 VTAIL.n139 0.155672
R506 VTAIL.n164 VTAIL.n163 0.155672
R507 VTAIL.n164 VTAIL.n135 0.155672
R508 VTAIL.n171 VTAIL.n135 0.155672
R509 VTAIL.n16 VTAIL.n11 0.155672
R510 VTAIL.n23 VTAIL.n11 0.155672
R511 VTAIL.n24 VTAIL.n23 0.155672
R512 VTAIL.n24 VTAIL.n7 0.155672
R513 VTAIL.n31 VTAIL.n7 0.155672
R514 VTAIL.n32 VTAIL.n31 0.155672
R515 VTAIL.n32 VTAIL.n3 0.155672
R516 VTAIL.n39 VTAIL.n3 0.155672
R517 VTAIL.n131 VTAIL.n95 0.155672
R518 VTAIL.n124 VTAIL.n95 0.155672
R519 VTAIL.n124 VTAIL.n123 0.155672
R520 VTAIL.n123 VTAIL.n99 0.155672
R521 VTAIL.n116 VTAIL.n99 0.155672
R522 VTAIL.n116 VTAIL.n115 0.155672
R523 VTAIL.n115 VTAIL.n103 0.155672
R524 VTAIL.n108 VTAIL.n103 0.155672
R525 VTAIL.n87 VTAIL.n51 0.155672
R526 VTAIL.n80 VTAIL.n51 0.155672
R527 VTAIL.n80 VTAIL.n79 0.155672
R528 VTAIL.n79 VTAIL.n55 0.155672
R529 VTAIL.n72 VTAIL.n55 0.155672
R530 VTAIL.n72 VTAIL.n71 0.155672
R531 VTAIL.n71 VTAIL.n59 0.155672
R532 VTAIL.n64 VTAIL.n59 0.155672
R533 B.n783 B.n782 585
R534 B.n267 B.n135 585
R535 B.n266 B.n265 585
R536 B.n264 B.n263 585
R537 B.n262 B.n261 585
R538 B.n260 B.n259 585
R539 B.n258 B.n257 585
R540 B.n256 B.n255 585
R541 B.n254 B.n253 585
R542 B.n252 B.n251 585
R543 B.n250 B.n249 585
R544 B.n248 B.n247 585
R545 B.n246 B.n245 585
R546 B.n244 B.n243 585
R547 B.n242 B.n241 585
R548 B.n240 B.n239 585
R549 B.n238 B.n237 585
R550 B.n236 B.n235 585
R551 B.n234 B.n233 585
R552 B.n232 B.n231 585
R553 B.n230 B.n229 585
R554 B.n228 B.n227 585
R555 B.n226 B.n225 585
R556 B.n224 B.n223 585
R557 B.n222 B.n221 585
R558 B.n220 B.n219 585
R559 B.n218 B.n217 585
R560 B.n216 B.n215 585
R561 B.n214 B.n213 585
R562 B.n212 B.n211 585
R563 B.n210 B.n209 585
R564 B.n208 B.n207 585
R565 B.n206 B.n205 585
R566 B.n204 B.n203 585
R567 B.n202 B.n201 585
R568 B.n200 B.n199 585
R569 B.n198 B.n197 585
R570 B.n196 B.n195 585
R571 B.n194 B.n193 585
R572 B.n192 B.n191 585
R573 B.n190 B.n189 585
R574 B.n188 B.n187 585
R575 B.n186 B.n185 585
R576 B.n184 B.n183 585
R577 B.n182 B.n181 585
R578 B.n180 B.n179 585
R579 B.n178 B.n177 585
R580 B.n176 B.n175 585
R581 B.n174 B.n173 585
R582 B.n172 B.n171 585
R583 B.n170 B.n169 585
R584 B.n168 B.n167 585
R585 B.n166 B.n165 585
R586 B.n164 B.n163 585
R587 B.n162 B.n161 585
R588 B.n160 B.n159 585
R589 B.n158 B.n157 585
R590 B.n156 B.n155 585
R591 B.n154 B.n153 585
R592 B.n152 B.n151 585
R593 B.n150 B.n149 585
R594 B.n148 B.n147 585
R595 B.n146 B.n145 585
R596 B.n144 B.n143 585
R597 B.n103 B.n102 585
R598 B.n788 B.n787 585
R599 B.n781 B.n136 585
R600 B.n136 B.n100 585
R601 B.n780 B.n99 585
R602 B.n792 B.n99 585
R603 B.n779 B.n98 585
R604 B.n793 B.n98 585
R605 B.n778 B.n97 585
R606 B.n794 B.n97 585
R607 B.n777 B.n776 585
R608 B.n776 B.n93 585
R609 B.n775 B.n92 585
R610 B.n800 B.n92 585
R611 B.n774 B.n91 585
R612 B.n801 B.n91 585
R613 B.n773 B.n90 585
R614 B.n802 B.n90 585
R615 B.n772 B.n771 585
R616 B.n771 B.n86 585
R617 B.n770 B.n85 585
R618 B.n808 B.n85 585
R619 B.n769 B.n84 585
R620 B.n809 B.n84 585
R621 B.n768 B.n83 585
R622 B.n810 B.n83 585
R623 B.n767 B.n766 585
R624 B.n766 B.n79 585
R625 B.n765 B.n78 585
R626 B.n816 B.n78 585
R627 B.n764 B.n77 585
R628 B.n817 B.n77 585
R629 B.n763 B.n76 585
R630 B.n818 B.n76 585
R631 B.n762 B.n761 585
R632 B.n761 B.n72 585
R633 B.n760 B.n71 585
R634 B.n824 B.n71 585
R635 B.n759 B.n70 585
R636 B.n825 B.n70 585
R637 B.n758 B.n69 585
R638 B.n826 B.n69 585
R639 B.n757 B.n756 585
R640 B.n756 B.n65 585
R641 B.n755 B.n64 585
R642 B.n832 B.n64 585
R643 B.n754 B.n63 585
R644 B.n833 B.n63 585
R645 B.n753 B.n62 585
R646 B.n834 B.n62 585
R647 B.n752 B.n751 585
R648 B.n751 B.n58 585
R649 B.n750 B.n57 585
R650 B.n840 B.n57 585
R651 B.n749 B.n56 585
R652 B.n841 B.n56 585
R653 B.n748 B.n55 585
R654 B.n842 B.n55 585
R655 B.n747 B.n746 585
R656 B.n746 B.n51 585
R657 B.n745 B.n50 585
R658 B.n848 B.n50 585
R659 B.n744 B.n49 585
R660 B.n849 B.n49 585
R661 B.n743 B.n48 585
R662 B.n850 B.n48 585
R663 B.n742 B.n741 585
R664 B.n741 B.n44 585
R665 B.n740 B.n43 585
R666 B.n856 B.n43 585
R667 B.n739 B.n42 585
R668 B.n857 B.n42 585
R669 B.n738 B.n41 585
R670 B.n858 B.n41 585
R671 B.n737 B.n736 585
R672 B.n736 B.n37 585
R673 B.n735 B.n36 585
R674 B.n864 B.n36 585
R675 B.n734 B.n35 585
R676 B.n865 B.n35 585
R677 B.n733 B.n34 585
R678 B.n866 B.n34 585
R679 B.n732 B.n731 585
R680 B.n731 B.n30 585
R681 B.n730 B.n29 585
R682 B.n872 B.n29 585
R683 B.n729 B.n28 585
R684 B.n873 B.n28 585
R685 B.n728 B.n27 585
R686 B.n874 B.n27 585
R687 B.n727 B.n726 585
R688 B.n726 B.n23 585
R689 B.n725 B.n22 585
R690 B.n880 B.n22 585
R691 B.n724 B.n21 585
R692 B.n881 B.n21 585
R693 B.n723 B.n20 585
R694 B.n882 B.n20 585
R695 B.n722 B.n721 585
R696 B.n721 B.n16 585
R697 B.n720 B.n15 585
R698 B.n888 B.n15 585
R699 B.n719 B.n14 585
R700 B.n889 B.n14 585
R701 B.n718 B.n13 585
R702 B.n890 B.n13 585
R703 B.n717 B.n716 585
R704 B.n716 B.n12 585
R705 B.n715 B.n714 585
R706 B.n715 B.n8 585
R707 B.n713 B.n7 585
R708 B.n897 B.n7 585
R709 B.n712 B.n6 585
R710 B.n898 B.n6 585
R711 B.n711 B.n5 585
R712 B.n899 B.n5 585
R713 B.n710 B.n709 585
R714 B.n709 B.n4 585
R715 B.n708 B.n268 585
R716 B.n708 B.n707 585
R717 B.n698 B.n269 585
R718 B.n270 B.n269 585
R719 B.n700 B.n699 585
R720 B.n701 B.n700 585
R721 B.n697 B.n275 585
R722 B.n275 B.n274 585
R723 B.n696 B.n695 585
R724 B.n695 B.n694 585
R725 B.n277 B.n276 585
R726 B.n278 B.n277 585
R727 B.n687 B.n686 585
R728 B.n688 B.n687 585
R729 B.n685 B.n283 585
R730 B.n283 B.n282 585
R731 B.n684 B.n683 585
R732 B.n683 B.n682 585
R733 B.n285 B.n284 585
R734 B.n286 B.n285 585
R735 B.n675 B.n674 585
R736 B.n676 B.n675 585
R737 B.n673 B.n291 585
R738 B.n291 B.n290 585
R739 B.n672 B.n671 585
R740 B.n671 B.n670 585
R741 B.n293 B.n292 585
R742 B.n294 B.n293 585
R743 B.n663 B.n662 585
R744 B.n664 B.n663 585
R745 B.n661 B.n299 585
R746 B.n299 B.n298 585
R747 B.n660 B.n659 585
R748 B.n659 B.n658 585
R749 B.n301 B.n300 585
R750 B.n302 B.n301 585
R751 B.n651 B.n650 585
R752 B.n652 B.n651 585
R753 B.n649 B.n306 585
R754 B.n310 B.n306 585
R755 B.n648 B.n647 585
R756 B.n647 B.n646 585
R757 B.n308 B.n307 585
R758 B.n309 B.n308 585
R759 B.n639 B.n638 585
R760 B.n640 B.n639 585
R761 B.n637 B.n315 585
R762 B.n315 B.n314 585
R763 B.n636 B.n635 585
R764 B.n635 B.n634 585
R765 B.n317 B.n316 585
R766 B.n318 B.n317 585
R767 B.n627 B.n626 585
R768 B.n628 B.n627 585
R769 B.n625 B.n322 585
R770 B.n326 B.n322 585
R771 B.n624 B.n623 585
R772 B.n623 B.n622 585
R773 B.n324 B.n323 585
R774 B.n325 B.n324 585
R775 B.n615 B.n614 585
R776 B.n616 B.n615 585
R777 B.n613 B.n331 585
R778 B.n331 B.n330 585
R779 B.n612 B.n611 585
R780 B.n611 B.n610 585
R781 B.n333 B.n332 585
R782 B.n334 B.n333 585
R783 B.n603 B.n602 585
R784 B.n604 B.n603 585
R785 B.n601 B.n338 585
R786 B.n342 B.n338 585
R787 B.n600 B.n599 585
R788 B.n599 B.n598 585
R789 B.n340 B.n339 585
R790 B.n341 B.n340 585
R791 B.n591 B.n590 585
R792 B.n592 B.n591 585
R793 B.n589 B.n347 585
R794 B.n347 B.n346 585
R795 B.n588 B.n587 585
R796 B.n587 B.n586 585
R797 B.n349 B.n348 585
R798 B.n350 B.n349 585
R799 B.n579 B.n578 585
R800 B.n580 B.n579 585
R801 B.n577 B.n355 585
R802 B.n355 B.n354 585
R803 B.n576 B.n575 585
R804 B.n575 B.n574 585
R805 B.n357 B.n356 585
R806 B.n358 B.n357 585
R807 B.n567 B.n566 585
R808 B.n568 B.n567 585
R809 B.n565 B.n363 585
R810 B.n363 B.n362 585
R811 B.n564 B.n563 585
R812 B.n563 B.n562 585
R813 B.n365 B.n364 585
R814 B.n366 B.n365 585
R815 B.n555 B.n554 585
R816 B.n556 B.n555 585
R817 B.n553 B.n371 585
R818 B.n371 B.n370 585
R819 B.n552 B.n551 585
R820 B.n551 B.n550 585
R821 B.n373 B.n372 585
R822 B.n374 B.n373 585
R823 B.n546 B.n545 585
R824 B.n377 B.n376 585
R825 B.n542 B.n541 585
R826 B.n543 B.n542 585
R827 B.n540 B.n410 585
R828 B.n539 B.n538 585
R829 B.n537 B.n536 585
R830 B.n535 B.n534 585
R831 B.n533 B.n532 585
R832 B.n531 B.n530 585
R833 B.n529 B.n528 585
R834 B.n527 B.n526 585
R835 B.n525 B.n524 585
R836 B.n523 B.n522 585
R837 B.n521 B.n520 585
R838 B.n519 B.n518 585
R839 B.n517 B.n516 585
R840 B.n515 B.n514 585
R841 B.n513 B.n512 585
R842 B.n511 B.n510 585
R843 B.n509 B.n508 585
R844 B.n507 B.n506 585
R845 B.n505 B.n504 585
R846 B.n503 B.n502 585
R847 B.n501 B.n500 585
R848 B.n499 B.n498 585
R849 B.n497 B.n496 585
R850 B.n495 B.n494 585
R851 B.n493 B.n492 585
R852 B.n490 B.n489 585
R853 B.n488 B.n487 585
R854 B.n486 B.n485 585
R855 B.n484 B.n483 585
R856 B.n482 B.n481 585
R857 B.n480 B.n479 585
R858 B.n478 B.n477 585
R859 B.n476 B.n475 585
R860 B.n474 B.n473 585
R861 B.n472 B.n471 585
R862 B.n469 B.n468 585
R863 B.n467 B.n466 585
R864 B.n465 B.n464 585
R865 B.n463 B.n462 585
R866 B.n461 B.n460 585
R867 B.n459 B.n458 585
R868 B.n457 B.n456 585
R869 B.n455 B.n454 585
R870 B.n453 B.n452 585
R871 B.n451 B.n450 585
R872 B.n449 B.n448 585
R873 B.n447 B.n446 585
R874 B.n445 B.n444 585
R875 B.n443 B.n442 585
R876 B.n441 B.n440 585
R877 B.n439 B.n438 585
R878 B.n437 B.n436 585
R879 B.n435 B.n434 585
R880 B.n433 B.n432 585
R881 B.n431 B.n430 585
R882 B.n429 B.n428 585
R883 B.n427 B.n426 585
R884 B.n425 B.n424 585
R885 B.n423 B.n422 585
R886 B.n421 B.n420 585
R887 B.n419 B.n418 585
R888 B.n417 B.n416 585
R889 B.n415 B.n409 585
R890 B.n543 B.n409 585
R891 B.n547 B.n375 585
R892 B.n375 B.n374 585
R893 B.n549 B.n548 585
R894 B.n550 B.n549 585
R895 B.n369 B.n368 585
R896 B.n370 B.n369 585
R897 B.n558 B.n557 585
R898 B.n557 B.n556 585
R899 B.n559 B.n367 585
R900 B.n367 B.n366 585
R901 B.n561 B.n560 585
R902 B.n562 B.n561 585
R903 B.n361 B.n360 585
R904 B.n362 B.n361 585
R905 B.n570 B.n569 585
R906 B.n569 B.n568 585
R907 B.n571 B.n359 585
R908 B.n359 B.n358 585
R909 B.n573 B.n572 585
R910 B.n574 B.n573 585
R911 B.n353 B.n352 585
R912 B.n354 B.n353 585
R913 B.n582 B.n581 585
R914 B.n581 B.n580 585
R915 B.n583 B.n351 585
R916 B.n351 B.n350 585
R917 B.n585 B.n584 585
R918 B.n586 B.n585 585
R919 B.n345 B.n344 585
R920 B.n346 B.n345 585
R921 B.n594 B.n593 585
R922 B.n593 B.n592 585
R923 B.n595 B.n343 585
R924 B.n343 B.n341 585
R925 B.n597 B.n596 585
R926 B.n598 B.n597 585
R927 B.n337 B.n336 585
R928 B.n342 B.n337 585
R929 B.n606 B.n605 585
R930 B.n605 B.n604 585
R931 B.n607 B.n335 585
R932 B.n335 B.n334 585
R933 B.n609 B.n608 585
R934 B.n610 B.n609 585
R935 B.n329 B.n328 585
R936 B.n330 B.n329 585
R937 B.n618 B.n617 585
R938 B.n617 B.n616 585
R939 B.n619 B.n327 585
R940 B.n327 B.n325 585
R941 B.n621 B.n620 585
R942 B.n622 B.n621 585
R943 B.n321 B.n320 585
R944 B.n326 B.n321 585
R945 B.n630 B.n629 585
R946 B.n629 B.n628 585
R947 B.n631 B.n319 585
R948 B.n319 B.n318 585
R949 B.n633 B.n632 585
R950 B.n634 B.n633 585
R951 B.n313 B.n312 585
R952 B.n314 B.n313 585
R953 B.n642 B.n641 585
R954 B.n641 B.n640 585
R955 B.n643 B.n311 585
R956 B.n311 B.n309 585
R957 B.n645 B.n644 585
R958 B.n646 B.n645 585
R959 B.n305 B.n304 585
R960 B.n310 B.n305 585
R961 B.n654 B.n653 585
R962 B.n653 B.n652 585
R963 B.n655 B.n303 585
R964 B.n303 B.n302 585
R965 B.n657 B.n656 585
R966 B.n658 B.n657 585
R967 B.n297 B.n296 585
R968 B.n298 B.n297 585
R969 B.n666 B.n665 585
R970 B.n665 B.n664 585
R971 B.n667 B.n295 585
R972 B.n295 B.n294 585
R973 B.n669 B.n668 585
R974 B.n670 B.n669 585
R975 B.n289 B.n288 585
R976 B.n290 B.n289 585
R977 B.n678 B.n677 585
R978 B.n677 B.n676 585
R979 B.n679 B.n287 585
R980 B.n287 B.n286 585
R981 B.n681 B.n680 585
R982 B.n682 B.n681 585
R983 B.n281 B.n280 585
R984 B.n282 B.n281 585
R985 B.n690 B.n689 585
R986 B.n689 B.n688 585
R987 B.n691 B.n279 585
R988 B.n279 B.n278 585
R989 B.n693 B.n692 585
R990 B.n694 B.n693 585
R991 B.n273 B.n272 585
R992 B.n274 B.n273 585
R993 B.n703 B.n702 585
R994 B.n702 B.n701 585
R995 B.n704 B.n271 585
R996 B.n271 B.n270 585
R997 B.n706 B.n705 585
R998 B.n707 B.n706 585
R999 B.n3 B.n0 585
R1000 B.n4 B.n3 585
R1001 B.n896 B.n1 585
R1002 B.n897 B.n896 585
R1003 B.n895 B.n894 585
R1004 B.n895 B.n8 585
R1005 B.n893 B.n9 585
R1006 B.n12 B.n9 585
R1007 B.n892 B.n891 585
R1008 B.n891 B.n890 585
R1009 B.n11 B.n10 585
R1010 B.n889 B.n11 585
R1011 B.n887 B.n886 585
R1012 B.n888 B.n887 585
R1013 B.n885 B.n17 585
R1014 B.n17 B.n16 585
R1015 B.n884 B.n883 585
R1016 B.n883 B.n882 585
R1017 B.n19 B.n18 585
R1018 B.n881 B.n19 585
R1019 B.n879 B.n878 585
R1020 B.n880 B.n879 585
R1021 B.n877 B.n24 585
R1022 B.n24 B.n23 585
R1023 B.n876 B.n875 585
R1024 B.n875 B.n874 585
R1025 B.n26 B.n25 585
R1026 B.n873 B.n26 585
R1027 B.n871 B.n870 585
R1028 B.n872 B.n871 585
R1029 B.n869 B.n31 585
R1030 B.n31 B.n30 585
R1031 B.n868 B.n867 585
R1032 B.n867 B.n866 585
R1033 B.n33 B.n32 585
R1034 B.n865 B.n33 585
R1035 B.n863 B.n862 585
R1036 B.n864 B.n863 585
R1037 B.n861 B.n38 585
R1038 B.n38 B.n37 585
R1039 B.n860 B.n859 585
R1040 B.n859 B.n858 585
R1041 B.n40 B.n39 585
R1042 B.n857 B.n40 585
R1043 B.n855 B.n854 585
R1044 B.n856 B.n855 585
R1045 B.n853 B.n45 585
R1046 B.n45 B.n44 585
R1047 B.n852 B.n851 585
R1048 B.n851 B.n850 585
R1049 B.n47 B.n46 585
R1050 B.n849 B.n47 585
R1051 B.n847 B.n846 585
R1052 B.n848 B.n847 585
R1053 B.n845 B.n52 585
R1054 B.n52 B.n51 585
R1055 B.n844 B.n843 585
R1056 B.n843 B.n842 585
R1057 B.n54 B.n53 585
R1058 B.n841 B.n54 585
R1059 B.n839 B.n838 585
R1060 B.n840 B.n839 585
R1061 B.n837 B.n59 585
R1062 B.n59 B.n58 585
R1063 B.n836 B.n835 585
R1064 B.n835 B.n834 585
R1065 B.n61 B.n60 585
R1066 B.n833 B.n61 585
R1067 B.n831 B.n830 585
R1068 B.n832 B.n831 585
R1069 B.n829 B.n66 585
R1070 B.n66 B.n65 585
R1071 B.n828 B.n827 585
R1072 B.n827 B.n826 585
R1073 B.n68 B.n67 585
R1074 B.n825 B.n68 585
R1075 B.n823 B.n822 585
R1076 B.n824 B.n823 585
R1077 B.n821 B.n73 585
R1078 B.n73 B.n72 585
R1079 B.n820 B.n819 585
R1080 B.n819 B.n818 585
R1081 B.n75 B.n74 585
R1082 B.n817 B.n75 585
R1083 B.n815 B.n814 585
R1084 B.n816 B.n815 585
R1085 B.n813 B.n80 585
R1086 B.n80 B.n79 585
R1087 B.n812 B.n811 585
R1088 B.n811 B.n810 585
R1089 B.n82 B.n81 585
R1090 B.n809 B.n82 585
R1091 B.n807 B.n806 585
R1092 B.n808 B.n807 585
R1093 B.n805 B.n87 585
R1094 B.n87 B.n86 585
R1095 B.n804 B.n803 585
R1096 B.n803 B.n802 585
R1097 B.n89 B.n88 585
R1098 B.n801 B.n89 585
R1099 B.n799 B.n798 585
R1100 B.n800 B.n799 585
R1101 B.n797 B.n94 585
R1102 B.n94 B.n93 585
R1103 B.n796 B.n795 585
R1104 B.n795 B.n794 585
R1105 B.n96 B.n95 585
R1106 B.n793 B.n96 585
R1107 B.n791 B.n790 585
R1108 B.n792 B.n791 585
R1109 B.n789 B.n101 585
R1110 B.n101 B.n100 585
R1111 B.n900 B.n899 585
R1112 B.n898 B.n2 585
R1113 B.n787 B.n101 530.939
R1114 B.n783 B.n136 530.939
R1115 B.n409 B.n373 530.939
R1116 B.n545 B.n375 530.939
R1117 B.n140 B.t20 283.123
R1118 B.n137 B.t16 283.123
R1119 B.n413 B.t9 283.123
R1120 B.n411 B.t13 283.123
R1121 B.n785 B.n784 256.663
R1122 B.n785 B.n134 256.663
R1123 B.n785 B.n133 256.663
R1124 B.n785 B.n132 256.663
R1125 B.n785 B.n131 256.663
R1126 B.n785 B.n130 256.663
R1127 B.n785 B.n129 256.663
R1128 B.n785 B.n128 256.663
R1129 B.n785 B.n127 256.663
R1130 B.n785 B.n126 256.663
R1131 B.n785 B.n125 256.663
R1132 B.n785 B.n124 256.663
R1133 B.n785 B.n123 256.663
R1134 B.n785 B.n122 256.663
R1135 B.n785 B.n121 256.663
R1136 B.n785 B.n120 256.663
R1137 B.n785 B.n119 256.663
R1138 B.n785 B.n118 256.663
R1139 B.n785 B.n117 256.663
R1140 B.n785 B.n116 256.663
R1141 B.n785 B.n115 256.663
R1142 B.n785 B.n114 256.663
R1143 B.n785 B.n113 256.663
R1144 B.n785 B.n112 256.663
R1145 B.n785 B.n111 256.663
R1146 B.n785 B.n110 256.663
R1147 B.n785 B.n109 256.663
R1148 B.n785 B.n108 256.663
R1149 B.n785 B.n107 256.663
R1150 B.n785 B.n106 256.663
R1151 B.n785 B.n105 256.663
R1152 B.n785 B.n104 256.663
R1153 B.n786 B.n785 256.663
R1154 B.n544 B.n543 256.663
R1155 B.n543 B.n378 256.663
R1156 B.n543 B.n379 256.663
R1157 B.n543 B.n380 256.663
R1158 B.n543 B.n381 256.663
R1159 B.n543 B.n382 256.663
R1160 B.n543 B.n383 256.663
R1161 B.n543 B.n384 256.663
R1162 B.n543 B.n385 256.663
R1163 B.n543 B.n386 256.663
R1164 B.n543 B.n387 256.663
R1165 B.n543 B.n388 256.663
R1166 B.n543 B.n389 256.663
R1167 B.n543 B.n390 256.663
R1168 B.n543 B.n391 256.663
R1169 B.n543 B.n392 256.663
R1170 B.n543 B.n393 256.663
R1171 B.n543 B.n394 256.663
R1172 B.n543 B.n395 256.663
R1173 B.n543 B.n396 256.663
R1174 B.n543 B.n397 256.663
R1175 B.n543 B.n398 256.663
R1176 B.n543 B.n399 256.663
R1177 B.n543 B.n400 256.663
R1178 B.n543 B.n401 256.663
R1179 B.n543 B.n402 256.663
R1180 B.n543 B.n403 256.663
R1181 B.n543 B.n404 256.663
R1182 B.n543 B.n405 256.663
R1183 B.n543 B.n406 256.663
R1184 B.n543 B.n407 256.663
R1185 B.n543 B.n408 256.663
R1186 B.n902 B.n901 256.663
R1187 B.n137 B.t18 255.888
R1188 B.n413 B.t12 255.888
R1189 B.n140 B.t21 255.888
R1190 B.n411 B.t15 255.888
R1191 B.n138 B.t19 203.525
R1192 B.n414 B.t11 203.525
R1193 B.n141 B.t22 203.525
R1194 B.n412 B.t14 203.525
R1195 B.n143 B.n103 163.367
R1196 B.n147 B.n146 163.367
R1197 B.n151 B.n150 163.367
R1198 B.n155 B.n154 163.367
R1199 B.n159 B.n158 163.367
R1200 B.n163 B.n162 163.367
R1201 B.n167 B.n166 163.367
R1202 B.n171 B.n170 163.367
R1203 B.n175 B.n174 163.367
R1204 B.n179 B.n178 163.367
R1205 B.n183 B.n182 163.367
R1206 B.n187 B.n186 163.367
R1207 B.n191 B.n190 163.367
R1208 B.n195 B.n194 163.367
R1209 B.n199 B.n198 163.367
R1210 B.n203 B.n202 163.367
R1211 B.n207 B.n206 163.367
R1212 B.n211 B.n210 163.367
R1213 B.n215 B.n214 163.367
R1214 B.n219 B.n218 163.367
R1215 B.n223 B.n222 163.367
R1216 B.n227 B.n226 163.367
R1217 B.n231 B.n230 163.367
R1218 B.n235 B.n234 163.367
R1219 B.n239 B.n238 163.367
R1220 B.n243 B.n242 163.367
R1221 B.n247 B.n246 163.367
R1222 B.n251 B.n250 163.367
R1223 B.n255 B.n254 163.367
R1224 B.n259 B.n258 163.367
R1225 B.n263 B.n262 163.367
R1226 B.n265 B.n135 163.367
R1227 B.n551 B.n373 163.367
R1228 B.n551 B.n371 163.367
R1229 B.n555 B.n371 163.367
R1230 B.n555 B.n365 163.367
R1231 B.n563 B.n365 163.367
R1232 B.n563 B.n363 163.367
R1233 B.n567 B.n363 163.367
R1234 B.n567 B.n357 163.367
R1235 B.n575 B.n357 163.367
R1236 B.n575 B.n355 163.367
R1237 B.n579 B.n355 163.367
R1238 B.n579 B.n349 163.367
R1239 B.n587 B.n349 163.367
R1240 B.n587 B.n347 163.367
R1241 B.n591 B.n347 163.367
R1242 B.n591 B.n340 163.367
R1243 B.n599 B.n340 163.367
R1244 B.n599 B.n338 163.367
R1245 B.n603 B.n338 163.367
R1246 B.n603 B.n333 163.367
R1247 B.n611 B.n333 163.367
R1248 B.n611 B.n331 163.367
R1249 B.n615 B.n331 163.367
R1250 B.n615 B.n324 163.367
R1251 B.n623 B.n324 163.367
R1252 B.n623 B.n322 163.367
R1253 B.n627 B.n322 163.367
R1254 B.n627 B.n317 163.367
R1255 B.n635 B.n317 163.367
R1256 B.n635 B.n315 163.367
R1257 B.n639 B.n315 163.367
R1258 B.n639 B.n308 163.367
R1259 B.n647 B.n308 163.367
R1260 B.n647 B.n306 163.367
R1261 B.n651 B.n306 163.367
R1262 B.n651 B.n301 163.367
R1263 B.n659 B.n301 163.367
R1264 B.n659 B.n299 163.367
R1265 B.n663 B.n299 163.367
R1266 B.n663 B.n293 163.367
R1267 B.n671 B.n293 163.367
R1268 B.n671 B.n291 163.367
R1269 B.n675 B.n291 163.367
R1270 B.n675 B.n285 163.367
R1271 B.n683 B.n285 163.367
R1272 B.n683 B.n283 163.367
R1273 B.n687 B.n283 163.367
R1274 B.n687 B.n277 163.367
R1275 B.n695 B.n277 163.367
R1276 B.n695 B.n275 163.367
R1277 B.n700 B.n275 163.367
R1278 B.n700 B.n269 163.367
R1279 B.n708 B.n269 163.367
R1280 B.n709 B.n708 163.367
R1281 B.n709 B.n5 163.367
R1282 B.n6 B.n5 163.367
R1283 B.n7 B.n6 163.367
R1284 B.n715 B.n7 163.367
R1285 B.n716 B.n715 163.367
R1286 B.n716 B.n13 163.367
R1287 B.n14 B.n13 163.367
R1288 B.n15 B.n14 163.367
R1289 B.n721 B.n15 163.367
R1290 B.n721 B.n20 163.367
R1291 B.n21 B.n20 163.367
R1292 B.n22 B.n21 163.367
R1293 B.n726 B.n22 163.367
R1294 B.n726 B.n27 163.367
R1295 B.n28 B.n27 163.367
R1296 B.n29 B.n28 163.367
R1297 B.n731 B.n29 163.367
R1298 B.n731 B.n34 163.367
R1299 B.n35 B.n34 163.367
R1300 B.n36 B.n35 163.367
R1301 B.n736 B.n36 163.367
R1302 B.n736 B.n41 163.367
R1303 B.n42 B.n41 163.367
R1304 B.n43 B.n42 163.367
R1305 B.n741 B.n43 163.367
R1306 B.n741 B.n48 163.367
R1307 B.n49 B.n48 163.367
R1308 B.n50 B.n49 163.367
R1309 B.n746 B.n50 163.367
R1310 B.n746 B.n55 163.367
R1311 B.n56 B.n55 163.367
R1312 B.n57 B.n56 163.367
R1313 B.n751 B.n57 163.367
R1314 B.n751 B.n62 163.367
R1315 B.n63 B.n62 163.367
R1316 B.n64 B.n63 163.367
R1317 B.n756 B.n64 163.367
R1318 B.n756 B.n69 163.367
R1319 B.n70 B.n69 163.367
R1320 B.n71 B.n70 163.367
R1321 B.n761 B.n71 163.367
R1322 B.n761 B.n76 163.367
R1323 B.n77 B.n76 163.367
R1324 B.n78 B.n77 163.367
R1325 B.n766 B.n78 163.367
R1326 B.n766 B.n83 163.367
R1327 B.n84 B.n83 163.367
R1328 B.n85 B.n84 163.367
R1329 B.n771 B.n85 163.367
R1330 B.n771 B.n90 163.367
R1331 B.n91 B.n90 163.367
R1332 B.n92 B.n91 163.367
R1333 B.n776 B.n92 163.367
R1334 B.n776 B.n97 163.367
R1335 B.n98 B.n97 163.367
R1336 B.n99 B.n98 163.367
R1337 B.n136 B.n99 163.367
R1338 B.n542 B.n377 163.367
R1339 B.n542 B.n410 163.367
R1340 B.n538 B.n537 163.367
R1341 B.n534 B.n533 163.367
R1342 B.n530 B.n529 163.367
R1343 B.n526 B.n525 163.367
R1344 B.n522 B.n521 163.367
R1345 B.n518 B.n517 163.367
R1346 B.n514 B.n513 163.367
R1347 B.n510 B.n509 163.367
R1348 B.n506 B.n505 163.367
R1349 B.n502 B.n501 163.367
R1350 B.n498 B.n497 163.367
R1351 B.n494 B.n493 163.367
R1352 B.n489 B.n488 163.367
R1353 B.n485 B.n484 163.367
R1354 B.n481 B.n480 163.367
R1355 B.n477 B.n476 163.367
R1356 B.n473 B.n472 163.367
R1357 B.n468 B.n467 163.367
R1358 B.n464 B.n463 163.367
R1359 B.n460 B.n459 163.367
R1360 B.n456 B.n455 163.367
R1361 B.n452 B.n451 163.367
R1362 B.n448 B.n447 163.367
R1363 B.n444 B.n443 163.367
R1364 B.n440 B.n439 163.367
R1365 B.n436 B.n435 163.367
R1366 B.n432 B.n431 163.367
R1367 B.n428 B.n427 163.367
R1368 B.n424 B.n423 163.367
R1369 B.n420 B.n419 163.367
R1370 B.n416 B.n409 163.367
R1371 B.n549 B.n375 163.367
R1372 B.n549 B.n369 163.367
R1373 B.n557 B.n369 163.367
R1374 B.n557 B.n367 163.367
R1375 B.n561 B.n367 163.367
R1376 B.n561 B.n361 163.367
R1377 B.n569 B.n361 163.367
R1378 B.n569 B.n359 163.367
R1379 B.n573 B.n359 163.367
R1380 B.n573 B.n353 163.367
R1381 B.n581 B.n353 163.367
R1382 B.n581 B.n351 163.367
R1383 B.n585 B.n351 163.367
R1384 B.n585 B.n345 163.367
R1385 B.n593 B.n345 163.367
R1386 B.n593 B.n343 163.367
R1387 B.n597 B.n343 163.367
R1388 B.n597 B.n337 163.367
R1389 B.n605 B.n337 163.367
R1390 B.n605 B.n335 163.367
R1391 B.n609 B.n335 163.367
R1392 B.n609 B.n329 163.367
R1393 B.n617 B.n329 163.367
R1394 B.n617 B.n327 163.367
R1395 B.n621 B.n327 163.367
R1396 B.n621 B.n321 163.367
R1397 B.n629 B.n321 163.367
R1398 B.n629 B.n319 163.367
R1399 B.n633 B.n319 163.367
R1400 B.n633 B.n313 163.367
R1401 B.n641 B.n313 163.367
R1402 B.n641 B.n311 163.367
R1403 B.n645 B.n311 163.367
R1404 B.n645 B.n305 163.367
R1405 B.n653 B.n305 163.367
R1406 B.n653 B.n303 163.367
R1407 B.n657 B.n303 163.367
R1408 B.n657 B.n297 163.367
R1409 B.n665 B.n297 163.367
R1410 B.n665 B.n295 163.367
R1411 B.n669 B.n295 163.367
R1412 B.n669 B.n289 163.367
R1413 B.n677 B.n289 163.367
R1414 B.n677 B.n287 163.367
R1415 B.n681 B.n287 163.367
R1416 B.n681 B.n281 163.367
R1417 B.n689 B.n281 163.367
R1418 B.n689 B.n279 163.367
R1419 B.n693 B.n279 163.367
R1420 B.n693 B.n273 163.367
R1421 B.n702 B.n273 163.367
R1422 B.n702 B.n271 163.367
R1423 B.n706 B.n271 163.367
R1424 B.n706 B.n3 163.367
R1425 B.n900 B.n3 163.367
R1426 B.n896 B.n2 163.367
R1427 B.n896 B.n895 163.367
R1428 B.n895 B.n9 163.367
R1429 B.n891 B.n9 163.367
R1430 B.n891 B.n11 163.367
R1431 B.n887 B.n11 163.367
R1432 B.n887 B.n17 163.367
R1433 B.n883 B.n17 163.367
R1434 B.n883 B.n19 163.367
R1435 B.n879 B.n19 163.367
R1436 B.n879 B.n24 163.367
R1437 B.n875 B.n24 163.367
R1438 B.n875 B.n26 163.367
R1439 B.n871 B.n26 163.367
R1440 B.n871 B.n31 163.367
R1441 B.n867 B.n31 163.367
R1442 B.n867 B.n33 163.367
R1443 B.n863 B.n33 163.367
R1444 B.n863 B.n38 163.367
R1445 B.n859 B.n38 163.367
R1446 B.n859 B.n40 163.367
R1447 B.n855 B.n40 163.367
R1448 B.n855 B.n45 163.367
R1449 B.n851 B.n45 163.367
R1450 B.n851 B.n47 163.367
R1451 B.n847 B.n47 163.367
R1452 B.n847 B.n52 163.367
R1453 B.n843 B.n52 163.367
R1454 B.n843 B.n54 163.367
R1455 B.n839 B.n54 163.367
R1456 B.n839 B.n59 163.367
R1457 B.n835 B.n59 163.367
R1458 B.n835 B.n61 163.367
R1459 B.n831 B.n61 163.367
R1460 B.n831 B.n66 163.367
R1461 B.n827 B.n66 163.367
R1462 B.n827 B.n68 163.367
R1463 B.n823 B.n68 163.367
R1464 B.n823 B.n73 163.367
R1465 B.n819 B.n73 163.367
R1466 B.n819 B.n75 163.367
R1467 B.n815 B.n75 163.367
R1468 B.n815 B.n80 163.367
R1469 B.n811 B.n80 163.367
R1470 B.n811 B.n82 163.367
R1471 B.n807 B.n82 163.367
R1472 B.n807 B.n87 163.367
R1473 B.n803 B.n87 163.367
R1474 B.n803 B.n89 163.367
R1475 B.n799 B.n89 163.367
R1476 B.n799 B.n94 163.367
R1477 B.n795 B.n94 163.367
R1478 B.n795 B.n96 163.367
R1479 B.n791 B.n96 163.367
R1480 B.n791 B.n101 163.367
R1481 B.n543 B.n374 122.174
R1482 B.n785 B.n100 122.174
R1483 B.n787 B.n786 71.676
R1484 B.n143 B.n104 71.676
R1485 B.n147 B.n105 71.676
R1486 B.n151 B.n106 71.676
R1487 B.n155 B.n107 71.676
R1488 B.n159 B.n108 71.676
R1489 B.n163 B.n109 71.676
R1490 B.n167 B.n110 71.676
R1491 B.n171 B.n111 71.676
R1492 B.n175 B.n112 71.676
R1493 B.n179 B.n113 71.676
R1494 B.n183 B.n114 71.676
R1495 B.n187 B.n115 71.676
R1496 B.n191 B.n116 71.676
R1497 B.n195 B.n117 71.676
R1498 B.n199 B.n118 71.676
R1499 B.n203 B.n119 71.676
R1500 B.n207 B.n120 71.676
R1501 B.n211 B.n121 71.676
R1502 B.n215 B.n122 71.676
R1503 B.n219 B.n123 71.676
R1504 B.n223 B.n124 71.676
R1505 B.n227 B.n125 71.676
R1506 B.n231 B.n126 71.676
R1507 B.n235 B.n127 71.676
R1508 B.n239 B.n128 71.676
R1509 B.n243 B.n129 71.676
R1510 B.n247 B.n130 71.676
R1511 B.n251 B.n131 71.676
R1512 B.n255 B.n132 71.676
R1513 B.n259 B.n133 71.676
R1514 B.n263 B.n134 71.676
R1515 B.n784 B.n135 71.676
R1516 B.n784 B.n783 71.676
R1517 B.n265 B.n134 71.676
R1518 B.n262 B.n133 71.676
R1519 B.n258 B.n132 71.676
R1520 B.n254 B.n131 71.676
R1521 B.n250 B.n130 71.676
R1522 B.n246 B.n129 71.676
R1523 B.n242 B.n128 71.676
R1524 B.n238 B.n127 71.676
R1525 B.n234 B.n126 71.676
R1526 B.n230 B.n125 71.676
R1527 B.n226 B.n124 71.676
R1528 B.n222 B.n123 71.676
R1529 B.n218 B.n122 71.676
R1530 B.n214 B.n121 71.676
R1531 B.n210 B.n120 71.676
R1532 B.n206 B.n119 71.676
R1533 B.n202 B.n118 71.676
R1534 B.n198 B.n117 71.676
R1535 B.n194 B.n116 71.676
R1536 B.n190 B.n115 71.676
R1537 B.n186 B.n114 71.676
R1538 B.n182 B.n113 71.676
R1539 B.n178 B.n112 71.676
R1540 B.n174 B.n111 71.676
R1541 B.n170 B.n110 71.676
R1542 B.n166 B.n109 71.676
R1543 B.n162 B.n108 71.676
R1544 B.n158 B.n107 71.676
R1545 B.n154 B.n106 71.676
R1546 B.n150 B.n105 71.676
R1547 B.n146 B.n104 71.676
R1548 B.n786 B.n103 71.676
R1549 B.n545 B.n544 71.676
R1550 B.n410 B.n378 71.676
R1551 B.n537 B.n379 71.676
R1552 B.n533 B.n380 71.676
R1553 B.n529 B.n381 71.676
R1554 B.n525 B.n382 71.676
R1555 B.n521 B.n383 71.676
R1556 B.n517 B.n384 71.676
R1557 B.n513 B.n385 71.676
R1558 B.n509 B.n386 71.676
R1559 B.n505 B.n387 71.676
R1560 B.n501 B.n388 71.676
R1561 B.n497 B.n389 71.676
R1562 B.n493 B.n390 71.676
R1563 B.n488 B.n391 71.676
R1564 B.n484 B.n392 71.676
R1565 B.n480 B.n393 71.676
R1566 B.n476 B.n394 71.676
R1567 B.n472 B.n395 71.676
R1568 B.n467 B.n396 71.676
R1569 B.n463 B.n397 71.676
R1570 B.n459 B.n398 71.676
R1571 B.n455 B.n399 71.676
R1572 B.n451 B.n400 71.676
R1573 B.n447 B.n401 71.676
R1574 B.n443 B.n402 71.676
R1575 B.n439 B.n403 71.676
R1576 B.n435 B.n404 71.676
R1577 B.n431 B.n405 71.676
R1578 B.n427 B.n406 71.676
R1579 B.n423 B.n407 71.676
R1580 B.n419 B.n408 71.676
R1581 B.n544 B.n377 71.676
R1582 B.n538 B.n378 71.676
R1583 B.n534 B.n379 71.676
R1584 B.n530 B.n380 71.676
R1585 B.n526 B.n381 71.676
R1586 B.n522 B.n382 71.676
R1587 B.n518 B.n383 71.676
R1588 B.n514 B.n384 71.676
R1589 B.n510 B.n385 71.676
R1590 B.n506 B.n386 71.676
R1591 B.n502 B.n387 71.676
R1592 B.n498 B.n388 71.676
R1593 B.n494 B.n389 71.676
R1594 B.n489 B.n390 71.676
R1595 B.n485 B.n391 71.676
R1596 B.n481 B.n392 71.676
R1597 B.n477 B.n393 71.676
R1598 B.n473 B.n394 71.676
R1599 B.n468 B.n395 71.676
R1600 B.n464 B.n396 71.676
R1601 B.n460 B.n397 71.676
R1602 B.n456 B.n398 71.676
R1603 B.n452 B.n399 71.676
R1604 B.n448 B.n400 71.676
R1605 B.n444 B.n401 71.676
R1606 B.n440 B.n402 71.676
R1607 B.n436 B.n403 71.676
R1608 B.n432 B.n404 71.676
R1609 B.n428 B.n405 71.676
R1610 B.n424 B.n406 71.676
R1611 B.n420 B.n407 71.676
R1612 B.n416 B.n408 71.676
R1613 B.n901 B.n900 71.676
R1614 B.n901 B.n2 71.676
R1615 B.n142 B.n141 59.5399
R1616 B.n139 B.n138 59.5399
R1617 B.n470 B.n414 59.5399
R1618 B.n491 B.n412 59.5399
R1619 B.n550 B.n374 58.9213
R1620 B.n550 B.n370 58.9213
R1621 B.n556 B.n370 58.9213
R1622 B.n556 B.n366 58.9213
R1623 B.n562 B.n366 58.9213
R1624 B.n562 B.n362 58.9213
R1625 B.n568 B.n362 58.9213
R1626 B.n574 B.n358 58.9213
R1627 B.n574 B.n354 58.9213
R1628 B.n580 B.n354 58.9213
R1629 B.n580 B.n350 58.9213
R1630 B.n586 B.n350 58.9213
R1631 B.n586 B.n346 58.9213
R1632 B.n592 B.n346 58.9213
R1633 B.n592 B.n341 58.9213
R1634 B.n598 B.n341 58.9213
R1635 B.n598 B.n342 58.9213
R1636 B.n604 B.n334 58.9213
R1637 B.n610 B.n334 58.9213
R1638 B.n610 B.n330 58.9213
R1639 B.n616 B.n330 58.9213
R1640 B.n616 B.n325 58.9213
R1641 B.n622 B.n325 58.9213
R1642 B.n622 B.n326 58.9213
R1643 B.n628 B.n318 58.9213
R1644 B.n634 B.n318 58.9213
R1645 B.n634 B.n314 58.9213
R1646 B.n640 B.n314 58.9213
R1647 B.n640 B.n309 58.9213
R1648 B.n646 B.n309 58.9213
R1649 B.n646 B.n310 58.9213
R1650 B.n652 B.n302 58.9213
R1651 B.n658 B.n302 58.9213
R1652 B.n658 B.n298 58.9213
R1653 B.n664 B.n298 58.9213
R1654 B.n664 B.n294 58.9213
R1655 B.n670 B.n294 58.9213
R1656 B.n676 B.n290 58.9213
R1657 B.n676 B.n286 58.9213
R1658 B.n682 B.n286 58.9213
R1659 B.n682 B.n282 58.9213
R1660 B.n688 B.n282 58.9213
R1661 B.n688 B.n278 58.9213
R1662 B.n694 B.n278 58.9213
R1663 B.n701 B.n274 58.9213
R1664 B.n701 B.n270 58.9213
R1665 B.n707 B.n270 58.9213
R1666 B.n707 B.n4 58.9213
R1667 B.n899 B.n4 58.9213
R1668 B.n899 B.n898 58.9213
R1669 B.n898 B.n897 58.9213
R1670 B.n897 B.n8 58.9213
R1671 B.n12 B.n8 58.9213
R1672 B.n890 B.n12 58.9213
R1673 B.n890 B.n889 58.9213
R1674 B.n888 B.n16 58.9213
R1675 B.n882 B.n16 58.9213
R1676 B.n882 B.n881 58.9213
R1677 B.n881 B.n880 58.9213
R1678 B.n880 B.n23 58.9213
R1679 B.n874 B.n23 58.9213
R1680 B.n874 B.n873 58.9213
R1681 B.n872 B.n30 58.9213
R1682 B.n866 B.n30 58.9213
R1683 B.n866 B.n865 58.9213
R1684 B.n865 B.n864 58.9213
R1685 B.n864 B.n37 58.9213
R1686 B.n858 B.n37 58.9213
R1687 B.n857 B.n856 58.9213
R1688 B.n856 B.n44 58.9213
R1689 B.n850 B.n44 58.9213
R1690 B.n850 B.n849 58.9213
R1691 B.n849 B.n848 58.9213
R1692 B.n848 B.n51 58.9213
R1693 B.n842 B.n51 58.9213
R1694 B.n841 B.n840 58.9213
R1695 B.n840 B.n58 58.9213
R1696 B.n834 B.n58 58.9213
R1697 B.n834 B.n833 58.9213
R1698 B.n833 B.n832 58.9213
R1699 B.n832 B.n65 58.9213
R1700 B.n826 B.n65 58.9213
R1701 B.n825 B.n824 58.9213
R1702 B.n824 B.n72 58.9213
R1703 B.n818 B.n72 58.9213
R1704 B.n818 B.n817 58.9213
R1705 B.n817 B.n816 58.9213
R1706 B.n816 B.n79 58.9213
R1707 B.n810 B.n79 58.9213
R1708 B.n810 B.n809 58.9213
R1709 B.n809 B.n808 58.9213
R1710 B.n808 B.n86 58.9213
R1711 B.n802 B.n801 58.9213
R1712 B.n801 B.n800 58.9213
R1713 B.n800 B.n93 58.9213
R1714 B.n794 B.n93 58.9213
R1715 B.n794 B.n793 58.9213
R1716 B.n793 B.n792 58.9213
R1717 B.n792 B.n100 58.9213
R1718 B.t10 B.n358 58.0549
R1719 B.n670 B.t0 58.0549
R1720 B.t6 B.n872 58.0549
R1721 B.t17 B.n86 58.0549
R1722 B.n652 B.t23 56.3219
R1723 B.n858 B.t2 56.3219
R1724 B.n694 B.t7 54.5889
R1725 B.t4 B.n888 54.5889
R1726 B.n628 B.t8 52.856
R1727 B.n842 B.t1 52.856
R1728 B.n141 B.n140 52.3641
R1729 B.n138 B.n137 52.3641
R1730 B.n414 B.n413 52.3641
R1731 B.n412 B.n411 52.3641
R1732 B.n604 B.t5 49.39
R1733 B.n826 B.t3 49.39
R1734 B.n547 B.n546 34.4981
R1735 B.n415 B.n372 34.4981
R1736 B.n782 B.n781 34.4981
R1737 B.n789 B.n788 34.4981
R1738 B B.n902 18.0485
R1739 B.n548 B.n547 10.6151
R1740 B.n548 B.n368 10.6151
R1741 B.n558 B.n368 10.6151
R1742 B.n559 B.n558 10.6151
R1743 B.n560 B.n559 10.6151
R1744 B.n560 B.n360 10.6151
R1745 B.n570 B.n360 10.6151
R1746 B.n571 B.n570 10.6151
R1747 B.n572 B.n571 10.6151
R1748 B.n572 B.n352 10.6151
R1749 B.n582 B.n352 10.6151
R1750 B.n583 B.n582 10.6151
R1751 B.n584 B.n583 10.6151
R1752 B.n584 B.n344 10.6151
R1753 B.n594 B.n344 10.6151
R1754 B.n595 B.n594 10.6151
R1755 B.n596 B.n595 10.6151
R1756 B.n596 B.n336 10.6151
R1757 B.n606 B.n336 10.6151
R1758 B.n607 B.n606 10.6151
R1759 B.n608 B.n607 10.6151
R1760 B.n608 B.n328 10.6151
R1761 B.n618 B.n328 10.6151
R1762 B.n619 B.n618 10.6151
R1763 B.n620 B.n619 10.6151
R1764 B.n620 B.n320 10.6151
R1765 B.n630 B.n320 10.6151
R1766 B.n631 B.n630 10.6151
R1767 B.n632 B.n631 10.6151
R1768 B.n632 B.n312 10.6151
R1769 B.n642 B.n312 10.6151
R1770 B.n643 B.n642 10.6151
R1771 B.n644 B.n643 10.6151
R1772 B.n644 B.n304 10.6151
R1773 B.n654 B.n304 10.6151
R1774 B.n655 B.n654 10.6151
R1775 B.n656 B.n655 10.6151
R1776 B.n656 B.n296 10.6151
R1777 B.n666 B.n296 10.6151
R1778 B.n667 B.n666 10.6151
R1779 B.n668 B.n667 10.6151
R1780 B.n668 B.n288 10.6151
R1781 B.n678 B.n288 10.6151
R1782 B.n679 B.n678 10.6151
R1783 B.n680 B.n679 10.6151
R1784 B.n680 B.n280 10.6151
R1785 B.n690 B.n280 10.6151
R1786 B.n691 B.n690 10.6151
R1787 B.n692 B.n691 10.6151
R1788 B.n692 B.n272 10.6151
R1789 B.n703 B.n272 10.6151
R1790 B.n704 B.n703 10.6151
R1791 B.n705 B.n704 10.6151
R1792 B.n705 B.n0 10.6151
R1793 B.n546 B.n376 10.6151
R1794 B.n541 B.n376 10.6151
R1795 B.n541 B.n540 10.6151
R1796 B.n540 B.n539 10.6151
R1797 B.n539 B.n536 10.6151
R1798 B.n536 B.n535 10.6151
R1799 B.n535 B.n532 10.6151
R1800 B.n532 B.n531 10.6151
R1801 B.n531 B.n528 10.6151
R1802 B.n528 B.n527 10.6151
R1803 B.n527 B.n524 10.6151
R1804 B.n524 B.n523 10.6151
R1805 B.n523 B.n520 10.6151
R1806 B.n520 B.n519 10.6151
R1807 B.n519 B.n516 10.6151
R1808 B.n516 B.n515 10.6151
R1809 B.n515 B.n512 10.6151
R1810 B.n512 B.n511 10.6151
R1811 B.n511 B.n508 10.6151
R1812 B.n508 B.n507 10.6151
R1813 B.n507 B.n504 10.6151
R1814 B.n504 B.n503 10.6151
R1815 B.n503 B.n500 10.6151
R1816 B.n500 B.n499 10.6151
R1817 B.n499 B.n496 10.6151
R1818 B.n496 B.n495 10.6151
R1819 B.n495 B.n492 10.6151
R1820 B.n490 B.n487 10.6151
R1821 B.n487 B.n486 10.6151
R1822 B.n486 B.n483 10.6151
R1823 B.n483 B.n482 10.6151
R1824 B.n482 B.n479 10.6151
R1825 B.n479 B.n478 10.6151
R1826 B.n478 B.n475 10.6151
R1827 B.n475 B.n474 10.6151
R1828 B.n474 B.n471 10.6151
R1829 B.n469 B.n466 10.6151
R1830 B.n466 B.n465 10.6151
R1831 B.n465 B.n462 10.6151
R1832 B.n462 B.n461 10.6151
R1833 B.n461 B.n458 10.6151
R1834 B.n458 B.n457 10.6151
R1835 B.n457 B.n454 10.6151
R1836 B.n454 B.n453 10.6151
R1837 B.n453 B.n450 10.6151
R1838 B.n450 B.n449 10.6151
R1839 B.n449 B.n446 10.6151
R1840 B.n446 B.n445 10.6151
R1841 B.n445 B.n442 10.6151
R1842 B.n442 B.n441 10.6151
R1843 B.n441 B.n438 10.6151
R1844 B.n438 B.n437 10.6151
R1845 B.n437 B.n434 10.6151
R1846 B.n434 B.n433 10.6151
R1847 B.n433 B.n430 10.6151
R1848 B.n430 B.n429 10.6151
R1849 B.n429 B.n426 10.6151
R1850 B.n426 B.n425 10.6151
R1851 B.n425 B.n422 10.6151
R1852 B.n422 B.n421 10.6151
R1853 B.n421 B.n418 10.6151
R1854 B.n418 B.n417 10.6151
R1855 B.n417 B.n415 10.6151
R1856 B.n552 B.n372 10.6151
R1857 B.n553 B.n552 10.6151
R1858 B.n554 B.n553 10.6151
R1859 B.n554 B.n364 10.6151
R1860 B.n564 B.n364 10.6151
R1861 B.n565 B.n564 10.6151
R1862 B.n566 B.n565 10.6151
R1863 B.n566 B.n356 10.6151
R1864 B.n576 B.n356 10.6151
R1865 B.n577 B.n576 10.6151
R1866 B.n578 B.n577 10.6151
R1867 B.n578 B.n348 10.6151
R1868 B.n588 B.n348 10.6151
R1869 B.n589 B.n588 10.6151
R1870 B.n590 B.n589 10.6151
R1871 B.n590 B.n339 10.6151
R1872 B.n600 B.n339 10.6151
R1873 B.n601 B.n600 10.6151
R1874 B.n602 B.n601 10.6151
R1875 B.n602 B.n332 10.6151
R1876 B.n612 B.n332 10.6151
R1877 B.n613 B.n612 10.6151
R1878 B.n614 B.n613 10.6151
R1879 B.n614 B.n323 10.6151
R1880 B.n624 B.n323 10.6151
R1881 B.n625 B.n624 10.6151
R1882 B.n626 B.n625 10.6151
R1883 B.n626 B.n316 10.6151
R1884 B.n636 B.n316 10.6151
R1885 B.n637 B.n636 10.6151
R1886 B.n638 B.n637 10.6151
R1887 B.n638 B.n307 10.6151
R1888 B.n648 B.n307 10.6151
R1889 B.n649 B.n648 10.6151
R1890 B.n650 B.n649 10.6151
R1891 B.n650 B.n300 10.6151
R1892 B.n660 B.n300 10.6151
R1893 B.n661 B.n660 10.6151
R1894 B.n662 B.n661 10.6151
R1895 B.n662 B.n292 10.6151
R1896 B.n672 B.n292 10.6151
R1897 B.n673 B.n672 10.6151
R1898 B.n674 B.n673 10.6151
R1899 B.n674 B.n284 10.6151
R1900 B.n684 B.n284 10.6151
R1901 B.n685 B.n684 10.6151
R1902 B.n686 B.n685 10.6151
R1903 B.n686 B.n276 10.6151
R1904 B.n696 B.n276 10.6151
R1905 B.n697 B.n696 10.6151
R1906 B.n699 B.n697 10.6151
R1907 B.n699 B.n698 10.6151
R1908 B.n698 B.n268 10.6151
R1909 B.n710 B.n268 10.6151
R1910 B.n711 B.n710 10.6151
R1911 B.n712 B.n711 10.6151
R1912 B.n713 B.n712 10.6151
R1913 B.n714 B.n713 10.6151
R1914 B.n717 B.n714 10.6151
R1915 B.n718 B.n717 10.6151
R1916 B.n719 B.n718 10.6151
R1917 B.n720 B.n719 10.6151
R1918 B.n722 B.n720 10.6151
R1919 B.n723 B.n722 10.6151
R1920 B.n724 B.n723 10.6151
R1921 B.n725 B.n724 10.6151
R1922 B.n727 B.n725 10.6151
R1923 B.n728 B.n727 10.6151
R1924 B.n729 B.n728 10.6151
R1925 B.n730 B.n729 10.6151
R1926 B.n732 B.n730 10.6151
R1927 B.n733 B.n732 10.6151
R1928 B.n734 B.n733 10.6151
R1929 B.n735 B.n734 10.6151
R1930 B.n737 B.n735 10.6151
R1931 B.n738 B.n737 10.6151
R1932 B.n739 B.n738 10.6151
R1933 B.n740 B.n739 10.6151
R1934 B.n742 B.n740 10.6151
R1935 B.n743 B.n742 10.6151
R1936 B.n744 B.n743 10.6151
R1937 B.n745 B.n744 10.6151
R1938 B.n747 B.n745 10.6151
R1939 B.n748 B.n747 10.6151
R1940 B.n749 B.n748 10.6151
R1941 B.n750 B.n749 10.6151
R1942 B.n752 B.n750 10.6151
R1943 B.n753 B.n752 10.6151
R1944 B.n754 B.n753 10.6151
R1945 B.n755 B.n754 10.6151
R1946 B.n757 B.n755 10.6151
R1947 B.n758 B.n757 10.6151
R1948 B.n759 B.n758 10.6151
R1949 B.n760 B.n759 10.6151
R1950 B.n762 B.n760 10.6151
R1951 B.n763 B.n762 10.6151
R1952 B.n764 B.n763 10.6151
R1953 B.n765 B.n764 10.6151
R1954 B.n767 B.n765 10.6151
R1955 B.n768 B.n767 10.6151
R1956 B.n769 B.n768 10.6151
R1957 B.n770 B.n769 10.6151
R1958 B.n772 B.n770 10.6151
R1959 B.n773 B.n772 10.6151
R1960 B.n774 B.n773 10.6151
R1961 B.n775 B.n774 10.6151
R1962 B.n777 B.n775 10.6151
R1963 B.n778 B.n777 10.6151
R1964 B.n779 B.n778 10.6151
R1965 B.n780 B.n779 10.6151
R1966 B.n781 B.n780 10.6151
R1967 B.n894 B.n1 10.6151
R1968 B.n894 B.n893 10.6151
R1969 B.n893 B.n892 10.6151
R1970 B.n892 B.n10 10.6151
R1971 B.n886 B.n10 10.6151
R1972 B.n886 B.n885 10.6151
R1973 B.n885 B.n884 10.6151
R1974 B.n884 B.n18 10.6151
R1975 B.n878 B.n18 10.6151
R1976 B.n878 B.n877 10.6151
R1977 B.n877 B.n876 10.6151
R1978 B.n876 B.n25 10.6151
R1979 B.n870 B.n25 10.6151
R1980 B.n870 B.n869 10.6151
R1981 B.n869 B.n868 10.6151
R1982 B.n868 B.n32 10.6151
R1983 B.n862 B.n32 10.6151
R1984 B.n862 B.n861 10.6151
R1985 B.n861 B.n860 10.6151
R1986 B.n860 B.n39 10.6151
R1987 B.n854 B.n39 10.6151
R1988 B.n854 B.n853 10.6151
R1989 B.n853 B.n852 10.6151
R1990 B.n852 B.n46 10.6151
R1991 B.n846 B.n46 10.6151
R1992 B.n846 B.n845 10.6151
R1993 B.n845 B.n844 10.6151
R1994 B.n844 B.n53 10.6151
R1995 B.n838 B.n53 10.6151
R1996 B.n838 B.n837 10.6151
R1997 B.n837 B.n836 10.6151
R1998 B.n836 B.n60 10.6151
R1999 B.n830 B.n60 10.6151
R2000 B.n830 B.n829 10.6151
R2001 B.n829 B.n828 10.6151
R2002 B.n828 B.n67 10.6151
R2003 B.n822 B.n67 10.6151
R2004 B.n822 B.n821 10.6151
R2005 B.n821 B.n820 10.6151
R2006 B.n820 B.n74 10.6151
R2007 B.n814 B.n74 10.6151
R2008 B.n814 B.n813 10.6151
R2009 B.n813 B.n812 10.6151
R2010 B.n812 B.n81 10.6151
R2011 B.n806 B.n81 10.6151
R2012 B.n806 B.n805 10.6151
R2013 B.n805 B.n804 10.6151
R2014 B.n804 B.n88 10.6151
R2015 B.n798 B.n88 10.6151
R2016 B.n798 B.n797 10.6151
R2017 B.n797 B.n796 10.6151
R2018 B.n796 B.n95 10.6151
R2019 B.n790 B.n95 10.6151
R2020 B.n790 B.n789 10.6151
R2021 B.n788 B.n102 10.6151
R2022 B.n144 B.n102 10.6151
R2023 B.n145 B.n144 10.6151
R2024 B.n148 B.n145 10.6151
R2025 B.n149 B.n148 10.6151
R2026 B.n152 B.n149 10.6151
R2027 B.n153 B.n152 10.6151
R2028 B.n156 B.n153 10.6151
R2029 B.n157 B.n156 10.6151
R2030 B.n160 B.n157 10.6151
R2031 B.n161 B.n160 10.6151
R2032 B.n164 B.n161 10.6151
R2033 B.n165 B.n164 10.6151
R2034 B.n168 B.n165 10.6151
R2035 B.n169 B.n168 10.6151
R2036 B.n172 B.n169 10.6151
R2037 B.n173 B.n172 10.6151
R2038 B.n176 B.n173 10.6151
R2039 B.n177 B.n176 10.6151
R2040 B.n180 B.n177 10.6151
R2041 B.n181 B.n180 10.6151
R2042 B.n184 B.n181 10.6151
R2043 B.n185 B.n184 10.6151
R2044 B.n188 B.n185 10.6151
R2045 B.n189 B.n188 10.6151
R2046 B.n192 B.n189 10.6151
R2047 B.n193 B.n192 10.6151
R2048 B.n197 B.n196 10.6151
R2049 B.n200 B.n197 10.6151
R2050 B.n201 B.n200 10.6151
R2051 B.n204 B.n201 10.6151
R2052 B.n205 B.n204 10.6151
R2053 B.n208 B.n205 10.6151
R2054 B.n209 B.n208 10.6151
R2055 B.n212 B.n209 10.6151
R2056 B.n213 B.n212 10.6151
R2057 B.n217 B.n216 10.6151
R2058 B.n220 B.n217 10.6151
R2059 B.n221 B.n220 10.6151
R2060 B.n224 B.n221 10.6151
R2061 B.n225 B.n224 10.6151
R2062 B.n228 B.n225 10.6151
R2063 B.n229 B.n228 10.6151
R2064 B.n232 B.n229 10.6151
R2065 B.n233 B.n232 10.6151
R2066 B.n236 B.n233 10.6151
R2067 B.n237 B.n236 10.6151
R2068 B.n240 B.n237 10.6151
R2069 B.n241 B.n240 10.6151
R2070 B.n244 B.n241 10.6151
R2071 B.n245 B.n244 10.6151
R2072 B.n248 B.n245 10.6151
R2073 B.n249 B.n248 10.6151
R2074 B.n252 B.n249 10.6151
R2075 B.n253 B.n252 10.6151
R2076 B.n256 B.n253 10.6151
R2077 B.n257 B.n256 10.6151
R2078 B.n260 B.n257 10.6151
R2079 B.n261 B.n260 10.6151
R2080 B.n264 B.n261 10.6151
R2081 B.n266 B.n264 10.6151
R2082 B.n267 B.n266 10.6151
R2083 B.n782 B.n267 10.6151
R2084 B.n342 B.t5 9.53181
R2085 B.t3 B.n825 9.53181
R2086 B.n492 B.n491 9.36635
R2087 B.n470 B.n469 9.36635
R2088 B.n193 B.n142 9.36635
R2089 B.n216 B.n139 9.36635
R2090 B.n902 B.n0 8.11757
R2091 B.n902 B.n1 8.11757
R2092 B.n326 B.t8 6.06588
R2093 B.t1 B.n841 6.06588
R2094 B.t7 B.n274 4.33291
R2095 B.n889 B.t4 4.33291
R2096 B.n310 B.t23 2.59995
R2097 B.t2 B.n857 2.59995
R2098 B.n491 B.n490 1.24928
R2099 B.n471 B.n470 1.24928
R2100 B.n196 B.n142 1.24928
R2101 B.n213 B.n139 1.24928
R2102 B.n568 B.t10 0.866983
R2103 B.t0 B.n290 0.866983
R2104 B.n873 B.t6 0.866983
R2105 B.n802 B.t17 0.866983
R2106 VP.n23 VP.n20 161.3
R2107 VP.n25 VP.n24 161.3
R2108 VP.n26 VP.n19 161.3
R2109 VP.n28 VP.n27 161.3
R2110 VP.n29 VP.n18 161.3
R2111 VP.n32 VP.n31 161.3
R2112 VP.n33 VP.n17 161.3
R2113 VP.n35 VP.n34 161.3
R2114 VP.n36 VP.n16 161.3
R2115 VP.n38 VP.n37 161.3
R2116 VP.n40 VP.n39 161.3
R2117 VP.n41 VP.n14 161.3
R2118 VP.n43 VP.n42 161.3
R2119 VP.n44 VP.n13 161.3
R2120 VP.n46 VP.n45 161.3
R2121 VP.n47 VP.n12 161.3
R2122 VP.n86 VP.n0 161.3
R2123 VP.n85 VP.n84 161.3
R2124 VP.n83 VP.n1 161.3
R2125 VP.n82 VP.n81 161.3
R2126 VP.n80 VP.n2 161.3
R2127 VP.n79 VP.n78 161.3
R2128 VP.n77 VP.n76 161.3
R2129 VP.n75 VP.n4 161.3
R2130 VP.n74 VP.n73 161.3
R2131 VP.n72 VP.n5 161.3
R2132 VP.n71 VP.n70 161.3
R2133 VP.n68 VP.n6 161.3
R2134 VP.n67 VP.n66 161.3
R2135 VP.n65 VP.n7 161.3
R2136 VP.n64 VP.n63 161.3
R2137 VP.n62 VP.n8 161.3
R2138 VP.n60 VP.n59 161.3
R2139 VP.n58 VP.n9 161.3
R2140 VP.n57 VP.n56 161.3
R2141 VP.n55 VP.n10 161.3
R2142 VP.n54 VP.n53 161.3
R2143 VP.n52 VP.n11 161.3
R2144 VP.n21 VP.t4 108.352
R2145 VP.n51 VP.n50 103.531
R2146 VP.n88 VP.n87 103.531
R2147 VP.n49 VP.n48 103.531
R2148 VP.n50 VP.t5 75.4528
R2149 VP.n61 VP.t6 75.4528
R2150 VP.n69 VP.t0 75.4528
R2151 VP.n3 VP.t3 75.4528
R2152 VP.n87 VP.t7 75.4528
R2153 VP.n48 VP.t1 75.4528
R2154 VP.n15 VP.t8 75.4528
R2155 VP.n30 VP.t2 75.4528
R2156 VP.n22 VP.t9 75.4528
R2157 VP.n56 VP.n55 56.5617
R2158 VP.n81 VP.n1 56.5617
R2159 VP.n42 VP.n13 56.5617
R2160 VP.n22 VP.n21 50.3824
R2161 VP.n63 VP.n7 50.2647
R2162 VP.n75 VP.n74 50.2647
R2163 VP.n36 VP.n35 50.2647
R2164 VP.n24 VP.n19 50.2647
R2165 VP.n51 VP.n49 48.3178
R2166 VP.n67 VP.n7 30.8893
R2167 VP.n74 VP.n5 30.8893
R2168 VP.n35 VP.n17 30.8893
R2169 VP.n28 VP.n19 30.8893
R2170 VP.n54 VP.n11 24.5923
R2171 VP.n55 VP.n54 24.5923
R2172 VP.n56 VP.n9 24.5923
R2173 VP.n60 VP.n9 24.5923
R2174 VP.n63 VP.n62 24.5923
R2175 VP.n68 VP.n67 24.5923
R2176 VP.n70 VP.n5 24.5923
R2177 VP.n76 VP.n75 24.5923
R2178 VP.n80 VP.n79 24.5923
R2179 VP.n81 VP.n80 24.5923
R2180 VP.n85 VP.n1 24.5923
R2181 VP.n86 VP.n85 24.5923
R2182 VP.n46 VP.n13 24.5923
R2183 VP.n47 VP.n46 24.5923
R2184 VP.n37 VP.n36 24.5923
R2185 VP.n41 VP.n40 24.5923
R2186 VP.n42 VP.n41 24.5923
R2187 VP.n29 VP.n28 24.5923
R2188 VP.n31 VP.n17 24.5923
R2189 VP.n24 VP.n23 24.5923
R2190 VP.n62 VP.n61 22.1332
R2191 VP.n76 VP.n3 22.1332
R2192 VP.n37 VP.n15 22.1332
R2193 VP.n23 VP.n22 22.1332
R2194 VP.n69 VP.n68 12.2964
R2195 VP.n70 VP.n69 12.2964
R2196 VP.n30 VP.n29 12.2964
R2197 VP.n31 VP.n30 12.2964
R2198 VP.n50 VP.n11 7.37805
R2199 VP.n87 VP.n86 7.37805
R2200 VP.n48 VP.n47 7.37805
R2201 VP.n21 VP.n20 6.9978
R2202 VP.n61 VP.n60 2.45968
R2203 VP.n79 VP.n3 2.45968
R2204 VP.n40 VP.n15 2.45968
R2205 VP.n49 VP.n12 0.278335
R2206 VP.n52 VP.n51 0.278335
R2207 VP.n88 VP.n0 0.278335
R2208 VP.n25 VP.n20 0.189894
R2209 VP.n26 VP.n25 0.189894
R2210 VP.n27 VP.n26 0.189894
R2211 VP.n27 VP.n18 0.189894
R2212 VP.n32 VP.n18 0.189894
R2213 VP.n33 VP.n32 0.189894
R2214 VP.n34 VP.n33 0.189894
R2215 VP.n34 VP.n16 0.189894
R2216 VP.n38 VP.n16 0.189894
R2217 VP.n39 VP.n38 0.189894
R2218 VP.n39 VP.n14 0.189894
R2219 VP.n43 VP.n14 0.189894
R2220 VP.n44 VP.n43 0.189894
R2221 VP.n45 VP.n44 0.189894
R2222 VP.n45 VP.n12 0.189894
R2223 VP.n53 VP.n52 0.189894
R2224 VP.n53 VP.n10 0.189894
R2225 VP.n57 VP.n10 0.189894
R2226 VP.n58 VP.n57 0.189894
R2227 VP.n59 VP.n58 0.189894
R2228 VP.n59 VP.n8 0.189894
R2229 VP.n64 VP.n8 0.189894
R2230 VP.n65 VP.n64 0.189894
R2231 VP.n66 VP.n65 0.189894
R2232 VP.n66 VP.n6 0.189894
R2233 VP.n71 VP.n6 0.189894
R2234 VP.n72 VP.n71 0.189894
R2235 VP.n73 VP.n72 0.189894
R2236 VP.n73 VP.n4 0.189894
R2237 VP.n77 VP.n4 0.189894
R2238 VP.n78 VP.n77 0.189894
R2239 VP.n78 VP.n2 0.189894
R2240 VP.n82 VP.n2 0.189894
R2241 VP.n83 VP.n82 0.189894
R2242 VP.n84 VP.n83 0.189894
R2243 VP.n84 VP.n0 0.189894
R2244 VP VP.n88 0.153485
R2245 VDD1.n34 VDD1.n0 289.615
R2246 VDD1.n75 VDD1.n41 289.615
R2247 VDD1.n35 VDD1.n34 185
R2248 VDD1.n33 VDD1.n32 185
R2249 VDD1.n4 VDD1.n3 185
R2250 VDD1.n27 VDD1.n26 185
R2251 VDD1.n25 VDD1.n24 185
R2252 VDD1.n8 VDD1.n7 185
R2253 VDD1.n19 VDD1.n18 185
R2254 VDD1.n17 VDD1.n16 185
R2255 VDD1.n12 VDD1.n11 185
R2256 VDD1.n53 VDD1.n52 185
R2257 VDD1.n58 VDD1.n57 185
R2258 VDD1.n60 VDD1.n59 185
R2259 VDD1.n49 VDD1.n48 185
R2260 VDD1.n66 VDD1.n65 185
R2261 VDD1.n68 VDD1.n67 185
R2262 VDD1.n45 VDD1.n44 185
R2263 VDD1.n74 VDD1.n73 185
R2264 VDD1.n76 VDD1.n75 185
R2265 VDD1.n13 VDD1.t5 147.659
R2266 VDD1.n54 VDD1.t4 147.659
R2267 VDD1.n34 VDD1.n33 104.615
R2268 VDD1.n33 VDD1.n3 104.615
R2269 VDD1.n26 VDD1.n3 104.615
R2270 VDD1.n26 VDD1.n25 104.615
R2271 VDD1.n25 VDD1.n7 104.615
R2272 VDD1.n18 VDD1.n7 104.615
R2273 VDD1.n18 VDD1.n17 104.615
R2274 VDD1.n17 VDD1.n11 104.615
R2275 VDD1.n58 VDD1.n52 104.615
R2276 VDD1.n59 VDD1.n58 104.615
R2277 VDD1.n59 VDD1.n48 104.615
R2278 VDD1.n66 VDD1.n48 104.615
R2279 VDD1.n67 VDD1.n66 104.615
R2280 VDD1.n67 VDD1.n44 104.615
R2281 VDD1.n74 VDD1.n44 104.615
R2282 VDD1.n75 VDD1.n74 104.615
R2283 VDD1.n83 VDD1.n82 66.5028
R2284 VDD1.n40 VDD1.n39 64.8126
R2285 VDD1.n85 VDD1.n84 64.8125
R2286 VDD1.n81 VDD1.n80 64.8125
R2287 VDD1.t5 VDD1.n11 52.3082
R2288 VDD1.t4 VDD1.n52 52.3082
R2289 VDD1.n40 VDD1.n38 50.8038
R2290 VDD1.n81 VDD1.n79 50.8038
R2291 VDD1.n85 VDD1.n83 42.9147
R2292 VDD1.n13 VDD1.n12 15.6677
R2293 VDD1.n54 VDD1.n53 15.6677
R2294 VDD1.n16 VDD1.n15 12.8005
R2295 VDD1.n57 VDD1.n56 12.8005
R2296 VDD1.n19 VDD1.n10 12.0247
R2297 VDD1.n60 VDD1.n51 12.0247
R2298 VDD1.n20 VDD1.n8 11.249
R2299 VDD1.n61 VDD1.n49 11.249
R2300 VDD1.n24 VDD1.n23 10.4732
R2301 VDD1.n65 VDD1.n64 10.4732
R2302 VDD1.n27 VDD1.n6 9.69747
R2303 VDD1.n68 VDD1.n47 9.69747
R2304 VDD1.n38 VDD1.n37 9.45567
R2305 VDD1.n79 VDD1.n78 9.45567
R2306 VDD1.n37 VDD1.n36 9.3005
R2307 VDD1.n2 VDD1.n1 9.3005
R2308 VDD1.n31 VDD1.n30 9.3005
R2309 VDD1.n29 VDD1.n28 9.3005
R2310 VDD1.n6 VDD1.n5 9.3005
R2311 VDD1.n23 VDD1.n22 9.3005
R2312 VDD1.n21 VDD1.n20 9.3005
R2313 VDD1.n10 VDD1.n9 9.3005
R2314 VDD1.n15 VDD1.n14 9.3005
R2315 VDD1.n78 VDD1.n77 9.3005
R2316 VDD1.n72 VDD1.n71 9.3005
R2317 VDD1.n70 VDD1.n69 9.3005
R2318 VDD1.n47 VDD1.n46 9.3005
R2319 VDD1.n64 VDD1.n63 9.3005
R2320 VDD1.n62 VDD1.n61 9.3005
R2321 VDD1.n51 VDD1.n50 9.3005
R2322 VDD1.n56 VDD1.n55 9.3005
R2323 VDD1.n43 VDD1.n42 9.3005
R2324 VDD1.n28 VDD1.n4 8.92171
R2325 VDD1.n69 VDD1.n45 8.92171
R2326 VDD1.n32 VDD1.n31 8.14595
R2327 VDD1.n73 VDD1.n72 8.14595
R2328 VDD1.n38 VDD1.n0 7.3702
R2329 VDD1.n35 VDD1.n2 7.3702
R2330 VDD1.n76 VDD1.n43 7.3702
R2331 VDD1.n79 VDD1.n41 7.3702
R2332 VDD1.n36 VDD1.n0 6.59444
R2333 VDD1.n36 VDD1.n35 6.59444
R2334 VDD1.n77 VDD1.n76 6.59444
R2335 VDD1.n77 VDD1.n41 6.59444
R2336 VDD1.n32 VDD1.n2 5.81868
R2337 VDD1.n73 VDD1.n43 5.81868
R2338 VDD1.n31 VDD1.n4 5.04292
R2339 VDD1.n72 VDD1.n45 5.04292
R2340 VDD1.n14 VDD1.n13 4.38565
R2341 VDD1.n55 VDD1.n54 4.38565
R2342 VDD1.n28 VDD1.n27 4.26717
R2343 VDD1.n69 VDD1.n68 4.26717
R2344 VDD1.n24 VDD1.n6 3.49141
R2345 VDD1.n65 VDD1.n47 3.49141
R2346 VDD1.n23 VDD1.n8 2.71565
R2347 VDD1.n64 VDD1.n49 2.71565
R2348 VDD1.n84 VDD1.t1 2.66896
R2349 VDD1.n84 VDD1.t8 2.66896
R2350 VDD1.n39 VDD1.t0 2.66896
R2351 VDD1.n39 VDD1.t7 2.66896
R2352 VDD1.n82 VDD1.t6 2.66896
R2353 VDD1.n82 VDD1.t2 2.66896
R2354 VDD1.n80 VDD1.t3 2.66896
R2355 VDD1.n80 VDD1.t9 2.66896
R2356 VDD1.n20 VDD1.n19 1.93989
R2357 VDD1.n61 VDD1.n60 1.93989
R2358 VDD1 VDD1.n85 1.688
R2359 VDD1.n16 VDD1.n10 1.16414
R2360 VDD1.n57 VDD1.n51 1.16414
R2361 VDD1 VDD1.n40 0.640586
R2362 VDD1.n83 VDD1.n81 0.527051
R2363 VDD1.n15 VDD1.n12 0.388379
R2364 VDD1.n56 VDD1.n53 0.388379
R2365 VDD1.n37 VDD1.n1 0.155672
R2366 VDD1.n30 VDD1.n1 0.155672
R2367 VDD1.n30 VDD1.n29 0.155672
R2368 VDD1.n29 VDD1.n5 0.155672
R2369 VDD1.n22 VDD1.n5 0.155672
R2370 VDD1.n22 VDD1.n21 0.155672
R2371 VDD1.n21 VDD1.n9 0.155672
R2372 VDD1.n14 VDD1.n9 0.155672
R2373 VDD1.n55 VDD1.n50 0.155672
R2374 VDD1.n62 VDD1.n50 0.155672
R2375 VDD1.n63 VDD1.n62 0.155672
R2376 VDD1.n63 VDD1.n46 0.155672
R2377 VDD1.n70 VDD1.n46 0.155672
R2378 VDD1.n71 VDD1.n70 0.155672
R2379 VDD1.n71 VDD1.n42 0.155672
R2380 VDD1.n78 VDD1.n42 0.155672
C0 VDD1 VP 7.05947f
C1 VN VTAIL 7.40723f
C2 VDD2 VP 0.554219f
C3 VTAIL VP 7.42146f
C4 VN VP 7.209f
C5 VDD1 VDD2 2.02438f
C6 VTAIL VDD1 8.15632f
C7 VTAIL VDD2 8.20662f
C8 VN VDD1 0.153198f
C9 VN VDD2 6.66145f
C10 VDD2 B 6.181821f
C11 VDD1 B 6.113869f
C12 VTAIL B 6.225391f
C13 VN B 16.688778f
C14 VP B 15.250366f
C15 VDD1.n0 B 0.037397f
C16 VDD1.n1 B 0.025861f
C17 VDD1.n2 B 0.013897f
C18 VDD1.n3 B 0.032847f
C19 VDD1.n4 B 0.014714f
C20 VDD1.n5 B 0.025861f
C21 VDD1.n6 B 0.013897f
C22 VDD1.n7 B 0.032847f
C23 VDD1.n8 B 0.014714f
C24 VDD1.n9 B 0.025861f
C25 VDD1.n10 B 0.013897f
C26 VDD1.n11 B 0.024635f
C27 VDD1.n12 B 0.019404f
C28 VDD1.t5 B 0.053535f
C29 VDD1.n13 B 0.119622f
C30 VDD1.n14 B 0.784021f
C31 VDD1.n15 B 0.013897f
C32 VDD1.n16 B 0.014714f
C33 VDD1.n17 B 0.032847f
C34 VDD1.n18 B 0.032847f
C35 VDD1.n19 B 0.014714f
C36 VDD1.n20 B 0.013897f
C37 VDD1.n21 B 0.025861f
C38 VDD1.n22 B 0.025861f
C39 VDD1.n23 B 0.013897f
C40 VDD1.n24 B 0.014714f
C41 VDD1.n25 B 0.032847f
C42 VDD1.n26 B 0.032847f
C43 VDD1.n27 B 0.014714f
C44 VDD1.n28 B 0.013897f
C45 VDD1.n29 B 0.025861f
C46 VDD1.n30 B 0.025861f
C47 VDD1.n31 B 0.013897f
C48 VDD1.n32 B 0.014714f
C49 VDD1.n33 B 0.032847f
C50 VDD1.n34 B 0.072959f
C51 VDD1.n35 B 0.014714f
C52 VDD1.n36 B 0.013897f
C53 VDD1.n37 B 0.05907f
C54 VDD1.n38 B 0.070003f
C55 VDD1.t0 B 0.151637f
C56 VDD1.t7 B 0.151637f
C57 VDD1.n39 B 1.29448f
C58 VDD1.n40 B 0.693679f
C59 VDD1.n41 B 0.037397f
C60 VDD1.n42 B 0.025861f
C61 VDD1.n43 B 0.013897f
C62 VDD1.n44 B 0.032847f
C63 VDD1.n45 B 0.014714f
C64 VDD1.n46 B 0.025861f
C65 VDD1.n47 B 0.013897f
C66 VDD1.n48 B 0.032847f
C67 VDD1.n49 B 0.014714f
C68 VDD1.n50 B 0.025861f
C69 VDD1.n51 B 0.013897f
C70 VDD1.n52 B 0.024635f
C71 VDD1.n53 B 0.019404f
C72 VDD1.t4 B 0.053535f
C73 VDD1.n54 B 0.119622f
C74 VDD1.n55 B 0.784021f
C75 VDD1.n56 B 0.013897f
C76 VDD1.n57 B 0.014714f
C77 VDD1.n58 B 0.032847f
C78 VDD1.n59 B 0.032847f
C79 VDD1.n60 B 0.014714f
C80 VDD1.n61 B 0.013897f
C81 VDD1.n62 B 0.025861f
C82 VDD1.n63 B 0.025861f
C83 VDD1.n64 B 0.013897f
C84 VDD1.n65 B 0.014714f
C85 VDD1.n66 B 0.032847f
C86 VDD1.n67 B 0.032847f
C87 VDD1.n68 B 0.014714f
C88 VDD1.n69 B 0.013897f
C89 VDD1.n70 B 0.025861f
C90 VDD1.n71 B 0.025861f
C91 VDD1.n72 B 0.013897f
C92 VDD1.n73 B 0.014714f
C93 VDD1.n74 B 0.032847f
C94 VDD1.n75 B 0.072959f
C95 VDD1.n76 B 0.014714f
C96 VDD1.n77 B 0.013897f
C97 VDD1.n78 B 0.05907f
C98 VDD1.n79 B 0.070003f
C99 VDD1.t3 B 0.151637f
C100 VDD1.t9 B 0.151637f
C101 VDD1.n80 B 1.29447f
C102 VDD1.n81 B 0.685363f
C103 VDD1.t6 B 0.151637f
C104 VDD1.t2 B 0.151637f
C105 VDD1.n82 B 1.3087f
C106 VDD1.n83 B 2.71326f
C107 VDD1.t1 B 0.151637f
C108 VDD1.t8 B 0.151637f
C109 VDD1.n84 B 1.29447f
C110 VDD1.n85 B 2.81975f
C111 VP.n0 B 0.032518f
C112 VP.t7 B 1.161f
C113 VP.n1 B 0.032444f
C114 VP.n2 B 0.024666f
C115 VP.t3 B 1.161f
C116 VP.n3 B 0.427786f
C117 VP.n4 B 0.024666f
C118 VP.n5 B 0.049148f
C119 VP.n6 B 0.024666f
C120 VP.t0 B 1.161f
C121 VP.n7 B 0.023257f
C122 VP.n8 B 0.024666f
C123 VP.t6 B 1.161f
C124 VP.n9 B 0.045741f
C125 VP.n10 B 0.024666f
C126 VP.n11 B 0.029934f
C127 VP.n12 B 0.032518f
C128 VP.t1 B 1.161f
C129 VP.n13 B 0.032444f
C130 VP.n14 B 0.024666f
C131 VP.t8 B 1.161f
C132 VP.n15 B 0.427786f
C133 VP.n16 B 0.024666f
C134 VP.n17 B 0.049148f
C135 VP.n18 B 0.024666f
C136 VP.t2 B 1.161f
C137 VP.n19 B 0.023257f
C138 VP.n20 B 0.232379f
C139 VP.t9 B 1.161f
C140 VP.t4 B 1.33375f
C141 VP.n21 B 0.481009f
C142 VP.n22 B 0.50495f
C143 VP.n23 B 0.043483f
C144 VP.n24 B 0.045049f
C145 VP.n25 B 0.024666f
C146 VP.n26 B 0.024666f
C147 VP.n27 B 0.024666f
C148 VP.n28 B 0.049148f
C149 VP.n29 B 0.034451f
C150 VP.n30 B 0.427786f
C151 VP.n31 B 0.034451f
C152 VP.n32 B 0.024666f
C153 VP.n33 B 0.024666f
C154 VP.n34 B 0.024666f
C155 VP.n35 B 0.023257f
C156 VP.n36 B 0.045049f
C157 VP.n37 B 0.043483f
C158 VP.n38 B 0.024666f
C159 VP.n39 B 0.024666f
C160 VP.n40 B 0.025418f
C161 VP.n41 B 0.045741f
C162 VP.n42 B 0.039268f
C163 VP.n43 B 0.024666f
C164 VP.n44 B 0.024666f
C165 VP.n45 B 0.024666f
C166 VP.n46 B 0.045741f
C167 VP.n47 B 0.029934f
C168 VP.n48 B 0.498918f
C169 VP.n49 B 1.30304f
C170 VP.t5 B 1.161f
C171 VP.n50 B 0.498918f
C172 VP.n51 B 1.32144f
C173 VP.n52 B 0.032518f
C174 VP.n53 B 0.024666f
C175 VP.n54 B 0.045741f
C176 VP.n55 B 0.032444f
C177 VP.n56 B 0.039268f
C178 VP.n57 B 0.024666f
C179 VP.n58 B 0.024666f
C180 VP.n59 B 0.024666f
C181 VP.n60 B 0.025418f
C182 VP.n61 B 0.427786f
C183 VP.n62 B 0.043483f
C184 VP.n63 B 0.045049f
C185 VP.n64 B 0.024666f
C186 VP.n65 B 0.024666f
C187 VP.n66 B 0.024666f
C188 VP.n67 B 0.049148f
C189 VP.n68 B 0.034451f
C190 VP.n69 B 0.427786f
C191 VP.n70 B 0.034451f
C192 VP.n71 B 0.024666f
C193 VP.n72 B 0.024666f
C194 VP.n73 B 0.024666f
C195 VP.n74 B 0.023257f
C196 VP.n75 B 0.045049f
C197 VP.n76 B 0.043483f
C198 VP.n77 B 0.024666f
C199 VP.n78 B 0.024666f
C200 VP.n79 B 0.025418f
C201 VP.n80 B 0.045741f
C202 VP.n81 B 0.039268f
C203 VP.n82 B 0.024666f
C204 VP.n83 B 0.024666f
C205 VP.n84 B 0.024666f
C206 VP.n85 B 0.045741f
C207 VP.n86 B 0.029934f
C208 VP.n87 B 0.498918f
C209 VP.n88 B 0.039752f
C210 VTAIL.t17 B 0.157119f
C211 VTAIL.t12 B 0.157119f
C212 VTAIL.n0 B 1.26614f
C213 VTAIL.n1 B 0.557444f
C214 VTAIL.n2 B 0.038749f
C215 VTAIL.n3 B 0.026796f
C216 VTAIL.n4 B 0.014399f
C217 VTAIL.n5 B 0.034034f
C218 VTAIL.n6 B 0.015246f
C219 VTAIL.n7 B 0.026796f
C220 VTAIL.n8 B 0.014399f
C221 VTAIL.n9 B 0.034034f
C222 VTAIL.n10 B 0.015246f
C223 VTAIL.n11 B 0.026796f
C224 VTAIL.n12 B 0.014399f
C225 VTAIL.n13 B 0.025526f
C226 VTAIL.n14 B 0.020105f
C227 VTAIL.t7 B 0.055471f
C228 VTAIL.n15 B 0.123947f
C229 VTAIL.n16 B 0.812366f
C230 VTAIL.n17 B 0.014399f
C231 VTAIL.n18 B 0.015246f
C232 VTAIL.n19 B 0.034034f
C233 VTAIL.n20 B 0.034034f
C234 VTAIL.n21 B 0.015246f
C235 VTAIL.n22 B 0.014399f
C236 VTAIL.n23 B 0.026796f
C237 VTAIL.n24 B 0.026796f
C238 VTAIL.n25 B 0.014399f
C239 VTAIL.n26 B 0.015246f
C240 VTAIL.n27 B 0.034034f
C241 VTAIL.n28 B 0.034034f
C242 VTAIL.n29 B 0.015246f
C243 VTAIL.n30 B 0.014399f
C244 VTAIL.n31 B 0.026796f
C245 VTAIL.n32 B 0.026796f
C246 VTAIL.n33 B 0.014399f
C247 VTAIL.n34 B 0.015246f
C248 VTAIL.n35 B 0.034034f
C249 VTAIL.n36 B 0.075596f
C250 VTAIL.n37 B 0.015246f
C251 VTAIL.n38 B 0.014399f
C252 VTAIL.n39 B 0.061206f
C253 VTAIL.n40 B 0.042474f
C254 VTAIL.n41 B 0.364496f
C255 VTAIL.t9 B 0.157119f
C256 VTAIL.t0 B 0.157119f
C257 VTAIL.n42 B 1.26614f
C258 VTAIL.n43 B 0.662582f
C259 VTAIL.t5 B 0.157119f
C260 VTAIL.t8 B 0.157119f
C261 VTAIL.n44 B 1.26614f
C262 VTAIL.n45 B 1.77984f
C263 VTAIL.t11 B 0.157119f
C264 VTAIL.t15 B 0.157119f
C265 VTAIL.n46 B 1.26615f
C266 VTAIL.n47 B 1.77984f
C267 VTAIL.t10 B 0.157119f
C268 VTAIL.t19 B 0.157119f
C269 VTAIL.n48 B 1.26615f
C270 VTAIL.n49 B 0.662573f
C271 VTAIL.n50 B 0.038749f
C272 VTAIL.n51 B 0.026796f
C273 VTAIL.n52 B 0.014399f
C274 VTAIL.n53 B 0.034034f
C275 VTAIL.n54 B 0.015246f
C276 VTAIL.n55 B 0.026796f
C277 VTAIL.n56 B 0.014399f
C278 VTAIL.n57 B 0.034034f
C279 VTAIL.n58 B 0.015246f
C280 VTAIL.n59 B 0.026796f
C281 VTAIL.n60 B 0.014399f
C282 VTAIL.n61 B 0.025526f
C283 VTAIL.n62 B 0.020105f
C284 VTAIL.t14 B 0.055471f
C285 VTAIL.n63 B 0.123947f
C286 VTAIL.n64 B 0.812366f
C287 VTAIL.n65 B 0.014399f
C288 VTAIL.n66 B 0.015246f
C289 VTAIL.n67 B 0.034034f
C290 VTAIL.n68 B 0.034034f
C291 VTAIL.n69 B 0.015246f
C292 VTAIL.n70 B 0.014399f
C293 VTAIL.n71 B 0.026796f
C294 VTAIL.n72 B 0.026796f
C295 VTAIL.n73 B 0.014399f
C296 VTAIL.n74 B 0.015246f
C297 VTAIL.n75 B 0.034034f
C298 VTAIL.n76 B 0.034034f
C299 VTAIL.n77 B 0.015246f
C300 VTAIL.n78 B 0.014399f
C301 VTAIL.n79 B 0.026796f
C302 VTAIL.n80 B 0.026796f
C303 VTAIL.n81 B 0.014399f
C304 VTAIL.n82 B 0.015246f
C305 VTAIL.n83 B 0.034034f
C306 VTAIL.n84 B 0.075596f
C307 VTAIL.n85 B 0.015246f
C308 VTAIL.n86 B 0.014399f
C309 VTAIL.n87 B 0.061206f
C310 VTAIL.n88 B 0.042474f
C311 VTAIL.n89 B 0.364496f
C312 VTAIL.t4 B 0.157119f
C313 VTAIL.t6 B 0.157119f
C314 VTAIL.n90 B 1.26615f
C315 VTAIL.n91 B 0.602654f
C316 VTAIL.t2 B 0.157119f
C317 VTAIL.t1 B 0.157119f
C318 VTAIL.n92 B 1.26615f
C319 VTAIL.n93 B 0.662573f
C320 VTAIL.n94 B 0.038749f
C321 VTAIL.n95 B 0.026796f
C322 VTAIL.n96 B 0.014399f
C323 VTAIL.n97 B 0.034034f
C324 VTAIL.n98 B 0.015246f
C325 VTAIL.n99 B 0.026796f
C326 VTAIL.n100 B 0.014399f
C327 VTAIL.n101 B 0.034034f
C328 VTAIL.n102 B 0.015246f
C329 VTAIL.n103 B 0.026796f
C330 VTAIL.n104 B 0.014399f
C331 VTAIL.n105 B 0.025526f
C332 VTAIL.n106 B 0.020105f
C333 VTAIL.t3 B 0.055471f
C334 VTAIL.n107 B 0.123947f
C335 VTAIL.n108 B 0.812366f
C336 VTAIL.n109 B 0.014399f
C337 VTAIL.n110 B 0.015246f
C338 VTAIL.n111 B 0.034034f
C339 VTAIL.n112 B 0.034034f
C340 VTAIL.n113 B 0.015246f
C341 VTAIL.n114 B 0.014399f
C342 VTAIL.n115 B 0.026796f
C343 VTAIL.n116 B 0.026796f
C344 VTAIL.n117 B 0.014399f
C345 VTAIL.n118 B 0.015246f
C346 VTAIL.n119 B 0.034034f
C347 VTAIL.n120 B 0.034034f
C348 VTAIL.n121 B 0.015246f
C349 VTAIL.n122 B 0.014399f
C350 VTAIL.n123 B 0.026796f
C351 VTAIL.n124 B 0.026796f
C352 VTAIL.n125 B 0.014399f
C353 VTAIL.n126 B 0.015246f
C354 VTAIL.n127 B 0.034034f
C355 VTAIL.n128 B 0.075596f
C356 VTAIL.n129 B 0.015246f
C357 VTAIL.n130 B 0.014399f
C358 VTAIL.n131 B 0.061206f
C359 VTAIL.n132 B 0.042474f
C360 VTAIL.n133 B 1.34071f
C361 VTAIL.n134 B 0.038749f
C362 VTAIL.n135 B 0.026796f
C363 VTAIL.n136 B 0.014399f
C364 VTAIL.n137 B 0.034034f
C365 VTAIL.n138 B 0.015246f
C366 VTAIL.n139 B 0.026796f
C367 VTAIL.n140 B 0.014399f
C368 VTAIL.n141 B 0.034034f
C369 VTAIL.n142 B 0.015246f
C370 VTAIL.n143 B 0.026796f
C371 VTAIL.n144 B 0.014399f
C372 VTAIL.n145 B 0.025526f
C373 VTAIL.n146 B 0.020105f
C374 VTAIL.t13 B 0.055471f
C375 VTAIL.n147 B 0.123947f
C376 VTAIL.n148 B 0.812366f
C377 VTAIL.n149 B 0.014399f
C378 VTAIL.n150 B 0.015246f
C379 VTAIL.n151 B 0.034034f
C380 VTAIL.n152 B 0.034034f
C381 VTAIL.n153 B 0.015246f
C382 VTAIL.n154 B 0.014399f
C383 VTAIL.n155 B 0.026796f
C384 VTAIL.n156 B 0.026796f
C385 VTAIL.n157 B 0.014399f
C386 VTAIL.n158 B 0.015246f
C387 VTAIL.n159 B 0.034034f
C388 VTAIL.n160 B 0.034034f
C389 VTAIL.n161 B 0.015246f
C390 VTAIL.n162 B 0.014399f
C391 VTAIL.n163 B 0.026796f
C392 VTAIL.n164 B 0.026796f
C393 VTAIL.n165 B 0.014399f
C394 VTAIL.n166 B 0.015246f
C395 VTAIL.n167 B 0.034034f
C396 VTAIL.n168 B 0.075596f
C397 VTAIL.n169 B 0.015246f
C398 VTAIL.n170 B 0.014399f
C399 VTAIL.n171 B 0.061206f
C400 VTAIL.n172 B 0.042474f
C401 VTAIL.n173 B 1.34071f
C402 VTAIL.t16 B 0.157119f
C403 VTAIL.t18 B 0.157119f
C404 VTAIL.n174 B 1.26614f
C405 VTAIL.n175 B 0.506829f
C406 VDD2.n0 B 0.036735f
C407 VDD2.n1 B 0.025403f
C408 VDD2.n2 B 0.013651f
C409 VDD2.n3 B 0.032265f
C410 VDD2.n4 B 0.014454f
C411 VDD2.n5 B 0.025403f
C412 VDD2.n6 B 0.013651f
C413 VDD2.n7 B 0.032265f
C414 VDD2.n8 B 0.014454f
C415 VDD2.n9 B 0.025403f
C416 VDD2.n10 B 0.013651f
C417 VDD2.n11 B 0.024199f
C418 VDD2.n12 B 0.01906f
C419 VDD2.t7 B 0.052588f
C420 VDD2.n13 B 0.117505f
C421 VDD2.n14 B 0.770146f
C422 VDD2.n15 B 0.013651f
C423 VDD2.n16 B 0.014454f
C424 VDD2.n17 B 0.032265f
C425 VDD2.n18 B 0.032265f
C426 VDD2.n19 B 0.014454f
C427 VDD2.n20 B 0.013651f
C428 VDD2.n21 B 0.025403f
C429 VDD2.n22 B 0.025403f
C430 VDD2.n23 B 0.013651f
C431 VDD2.n24 B 0.014454f
C432 VDD2.n25 B 0.032265f
C433 VDD2.n26 B 0.032265f
C434 VDD2.n27 B 0.014454f
C435 VDD2.n28 B 0.013651f
C436 VDD2.n29 B 0.025403f
C437 VDD2.n30 B 0.025403f
C438 VDD2.n31 B 0.013651f
C439 VDD2.n32 B 0.014454f
C440 VDD2.n33 B 0.032265f
C441 VDD2.n34 B 0.071668f
C442 VDD2.n35 B 0.014454f
C443 VDD2.n36 B 0.013651f
C444 VDD2.n37 B 0.058025f
C445 VDD2.n38 B 0.068764f
C446 VDD2.t3 B 0.148954f
C447 VDD2.t6 B 0.148954f
C448 VDD2.n39 B 1.27156f
C449 VDD2.n40 B 0.673233f
C450 VDD2.t8 B 0.148954f
C451 VDD2.t2 B 0.148954f
C452 VDD2.n41 B 1.28554f
C453 VDD2.n42 B 2.54788f
C454 VDD2.n43 B 0.036735f
C455 VDD2.n44 B 0.025403f
C456 VDD2.n45 B 0.013651f
C457 VDD2.n46 B 0.032265f
C458 VDD2.n47 B 0.014454f
C459 VDD2.n48 B 0.025403f
C460 VDD2.n49 B 0.013651f
C461 VDD2.n50 B 0.032265f
C462 VDD2.n51 B 0.014454f
C463 VDD2.n52 B 0.025403f
C464 VDD2.n53 B 0.013651f
C465 VDD2.n54 B 0.024199f
C466 VDD2.n55 B 0.01906f
C467 VDD2.t4 B 0.052588f
C468 VDD2.n56 B 0.117505f
C469 VDD2.n57 B 0.770146f
C470 VDD2.n58 B 0.013651f
C471 VDD2.n59 B 0.014454f
C472 VDD2.n60 B 0.032265f
C473 VDD2.n61 B 0.032265f
C474 VDD2.n62 B 0.014454f
C475 VDD2.n63 B 0.013651f
C476 VDD2.n64 B 0.025403f
C477 VDD2.n65 B 0.025403f
C478 VDD2.n66 B 0.013651f
C479 VDD2.n67 B 0.014454f
C480 VDD2.n68 B 0.032265f
C481 VDD2.n69 B 0.032265f
C482 VDD2.n70 B 0.014454f
C483 VDD2.n71 B 0.013651f
C484 VDD2.n72 B 0.025403f
C485 VDD2.n73 B 0.025403f
C486 VDD2.n74 B 0.013651f
C487 VDD2.n75 B 0.014454f
C488 VDD2.n76 B 0.032265f
C489 VDD2.n77 B 0.071668f
C490 VDD2.n78 B 0.014454f
C491 VDD2.n79 B 0.013651f
C492 VDD2.n80 B 0.058025f
C493 VDD2.n81 B 0.057812f
C494 VDD2.n82 B 2.48314f
C495 VDD2.t0 B 0.148954f
C496 VDD2.t5 B 0.148954f
C497 VDD2.n83 B 1.27157f
C498 VDD2.n84 B 0.453309f
C499 VDD2.t1 B 0.148954f
C500 VDD2.t9 B 0.148954f
C501 VDD2.n85 B 1.2855f
C502 VN.n0 B 0.031868f
C503 VN.t6 B 1.13778f
C504 VN.n1 B 0.031795f
C505 VN.n2 B 0.024173f
C506 VN.t1 B 1.13778f
C507 VN.n3 B 0.41923f
C508 VN.n4 B 0.024173f
C509 VN.n5 B 0.048165f
C510 VN.n6 B 0.024173f
C511 VN.t3 B 1.13778f
C512 VN.n7 B 0.022791f
C513 VN.n8 B 0.227732f
C514 VN.t7 B 1.13778f
C515 VN.t2 B 1.30708f
C516 VN.n9 B 0.471389f
C517 VN.n10 B 0.494851f
C518 VN.n11 B 0.042613f
C519 VN.n12 B 0.044148f
C520 VN.n13 B 0.024173f
C521 VN.n14 B 0.024173f
C522 VN.n15 B 0.024173f
C523 VN.n16 B 0.048165f
C524 VN.n17 B 0.033762f
C525 VN.n18 B 0.41923f
C526 VN.n19 B 0.033762f
C527 VN.n20 B 0.024173f
C528 VN.n21 B 0.024173f
C529 VN.n22 B 0.024173f
C530 VN.n23 B 0.022791f
C531 VN.n24 B 0.044148f
C532 VN.n25 B 0.042613f
C533 VN.n26 B 0.024173f
C534 VN.n27 B 0.024173f
C535 VN.n28 B 0.02491f
C536 VN.n29 B 0.044826f
C537 VN.n30 B 0.038483f
C538 VN.n31 B 0.024173f
C539 VN.n32 B 0.024173f
C540 VN.n33 B 0.024173f
C541 VN.n34 B 0.044826f
C542 VN.n35 B 0.029336f
C543 VN.n36 B 0.48894f
C544 VN.n37 B 0.038957f
C545 VN.n38 B 0.031868f
C546 VN.t8 B 1.13778f
C547 VN.n39 B 0.031795f
C548 VN.n40 B 0.024173f
C549 VN.t4 B 1.13778f
C550 VN.n41 B 0.41923f
C551 VN.n42 B 0.024173f
C552 VN.n43 B 0.048165f
C553 VN.n44 B 0.024173f
C554 VN.t9 B 1.13778f
C555 VN.n45 B 0.022791f
C556 VN.n46 B 0.227732f
C557 VN.t0 B 1.13778f
C558 VN.t5 B 1.30708f
C559 VN.n47 B 0.471389f
C560 VN.n48 B 0.494851f
C561 VN.n49 B 0.042613f
C562 VN.n50 B 0.044148f
C563 VN.n51 B 0.024173f
C564 VN.n52 B 0.024173f
C565 VN.n53 B 0.024173f
C566 VN.n54 B 0.048165f
C567 VN.n55 B 0.033762f
C568 VN.n56 B 0.41923f
C569 VN.n57 B 0.033762f
C570 VN.n58 B 0.024173f
C571 VN.n59 B 0.024173f
C572 VN.n60 B 0.024173f
C573 VN.n61 B 0.022791f
C574 VN.n62 B 0.044148f
C575 VN.n63 B 0.042613f
C576 VN.n64 B 0.024173f
C577 VN.n65 B 0.024173f
C578 VN.n66 B 0.02491f
C579 VN.n67 B 0.044826f
C580 VN.n68 B 0.038483f
C581 VN.n69 B 0.024173f
C582 VN.n70 B 0.024173f
C583 VN.n71 B 0.024173f
C584 VN.n72 B 0.044826f
C585 VN.n73 B 0.029336f
C586 VN.n74 B 0.48894f
C587 VN.n75 B 1.29004f
.ends

