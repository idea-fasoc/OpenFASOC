* NGSPICE file created from diff_pair_sample_0625.ext - technology: sky130A

.subckt diff_pair_sample_0625 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=0.46
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.46
X2 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.46
X3 VTAIL.t9 VP.t1 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X4 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X5 VDD2.t6 VN.t1 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X6 VTAIL.t1 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=0.46
X7 VDD1.t2 VP.t2 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X8 VDD2.t4 VN.t3 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=0.46
X9 VDD1.t7 VP.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X10 VTAIL.t11 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X11 VTAIL.t6 VP.t4 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X12 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=0.46
X13 VDD1.t0 VP.t5 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=0.46
X14 VTAIL.t4 VP.t6 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0.5478 ps=3.65 w=3.32 l=0.46
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.46
X16 VDD2.t1 VN.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=0.5478 ps=3.65 w=3.32 l=0.46
X17 VDD2.t0 VN.t7 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=0.46
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.46
X19 VDD1.t1 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5478 pd=3.65 as=1.2948 ps=7.42 w=3.32 l=0.46
R0 VP.n4 VP.t6 280.32
R1 VP.n10 VP.t0 259.337
R2 VP.n1 VP.t3 259.337
R3 VP.n15 VP.t1 259.337
R4 VP.n16 VP.t7 259.337
R5 VP.n8 VP.t5 259.337
R6 VP.n7 VP.t4 259.337
R7 VP.n3 VP.t2 259.337
R8 VP.n17 VP.n16 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n7 VP.n2 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n15 VP.n0 161.3
R13 VP.n14 VP.n13 161.3
R14 VP.n12 VP.n1 161.3
R15 VP.n11 VP.n10 161.3
R16 VP.n5 VP.n4 70.4033
R17 VP.n10 VP.n1 48.2005
R18 VP.n16 VP.n15 48.2005
R19 VP.n8 VP.n7 48.2005
R20 VP.n11 VP.n9 34.3414
R21 VP.n14 VP.n1 24.1005
R22 VP.n15 VP.n14 24.1005
R23 VP.n6 VP.n3 24.1005
R24 VP.n7 VP.n6 24.1005
R25 VP.n4 VP.n3 20.9576
R26 VP.n5 VP.n2 0.189894
R27 VP.n9 VP.n2 0.189894
R28 VP.n12 VP.n11 0.189894
R29 VP.n13 VP.n12 0.189894
R30 VP.n13 VP.n0 0.189894
R31 VP.n17 VP.n0 0.189894
R32 VP VP.n17 0.0516364
R33 VDD1 VDD1.n0 82.0267
R34 VDD1.n3 VDD1.n2 81.913
R35 VDD1.n3 VDD1.n1 81.913
R36 VDD1.n5 VDD1.n4 81.6279
R37 VDD1.n5 VDD1.n3 30.225
R38 VDD1.n4 VDD1.t4 5.96436
R39 VDD1.n4 VDD1.t0 5.96436
R40 VDD1.n0 VDD1.t5 5.96436
R41 VDD1.n0 VDD1.t2 5.96436
R42 VDD1.n2 VDD1.t3 5.96436
R43 VDD1.n2 VDD1.t1 5.96436
R44 VDD1.n1 VDD1.t6 5.96436
R45 VDD1.n1 VDD1.t7 5.96436
R46 VDD1 VDD1.n5 0.282828
R47 VTAIL.n130 VTAIL.n120 289.615
R48 VTAIL.n12 VTAIL.n2 289.615
R49 VTAIL.n28 VTAIL.n18 289.615
R50 VTAIL.n46 VTAIL.n36 289.615
R51 VTAIL.n114 VTAIL.n104 289.615
R52 VTAIL.n96 VTAIL.n86 289.615
R53 VTAIL.n80 VTAIL.n70 289.615
R54 VTAIL.n62 VTAIL.n52 289.615
R55 VTAIL.n124 VTAIL.n123 185
R56 VTAIL.n129 VTAIL.n128 185
R57 VTAIL.n131 VTAIL.n130 185
R58 VTAIL.n6 VTAIL.n5 185
R59 VTAIL.n11 VTAIL.n10 185
R60 VTAIL.n13 VTAIL.n12 185
R61 VTAIL.n22 VTAIL.n21 185
R62 VTAIL.n27 VTAIL.n26 185
R63 VTAIL.n29 VTAIL.n28 185
R64 VTAIL.n40 VTAIL.n39 185
R65 VTAIL.n45 VTAIL.n44 185
R66 VTAIL.n47 VTAIL.n46 185
R67 VTAIL.n115 VTAIL.n114 185
R68 VTAIL.n113 VTAIL.n112 185
R69 VTAIL.n108 VTAIL.n107 185
R70 VTAIL.n97 VTAIL.n96 185
R71 VTAIL.n95 VTAIL.n94 185
R72 VTAIL.n90 VTAIL.n89 185
R73 VTAIL.n81 VTAIL.n80 185
R74 VTAIL.n79 VTAIL.n78 185
R75 VTAIL.n74 VTAIL.n73 185
R76 VTAIL.n63 VTAIL.n62 185
R77 VTAIL.n61 VTAIL.n60 185
R78 VTAIL.n56 VTAIL.n55 185
R79 VTAIL.n125 VTAIL.t14 148.606
R80 VTAIL.n7 VTAIL.t0 148.606
R81 VTAIL.n23 VTAIL.t3 148.606
R82 VTAIL.n41 VTAIL.t10 148.606
R83 VTAIL.n109 VTAIL.t5 148.606
R84 VTAIL.n91 VTAIL.t4 148.606
R85 VTAIL.n75 VTAIL.t15 148.606
R86 VTAIL.n57 VTAIL.t1 148.606
R87 VTAIL.n129 VTAIL.n123 104.615
R88 VTAIL.n130 VTAIL.n129 104.615
R89 VTAIL.n11 VTAIL.n5 104.615
R90 VTAIL.n12 VTAIL.n11 104.615
R91 VTAIL.n27 VTAIL.n21 104.615
R92 VTAIL.n28 VTAIL.n27 104.615
R93 VTAIL.n45 VTAIL.n39 104.615
R94 VTAIL.n46 VTAIL.n45 104.615
R95 VTAIL.n114 VTAIL.n113 104.615
R96 VTAIL.n113 VTAIL.n107 104.615
R97 VTAIL.n96 VTAIL.n95 104.615
R98 VTAIL.n95 VTAIL.n89 104.615
R99 VTAIL.n80 VTAIL.n79 104.615
R100 VTAIL.n79 VTAIL.n73 104.615
R101 VTAIL.n62 VTAIL.n61 104.615
R102 VTAIL.n61 VTAIL.n55 104.615
R103 VTAIL.n103 VTAIL.n102 64.9492
R104 VTAIL.n69 VTAIL.n68 64.9492
R105 VTAIL.n1 VTAIL.n0 64.9491
R106 VTAIL.n35 VTAIL.n34 64.9491
R107 VTAIL.t14 VTAIL.n123 52.3082
R108 VTAIL.t0 VTAIL.n5 52.3082
R109 VTAIL.t3 VTAIL.n21 52.3082
R110 VTAIL.t10 VTAIL.n39 52.3082
R111 VTAIL.t5 VTAIL.n107 52.3082
R112 VTAIL.t4 VTAIL.n89 52.3082
R113 VTAIL.t15 VTAIL.n73 52.3082
R114 VTAIL.t1 VTAIL.n55 52.3082
R115 VTAIL.n135 VTAIL.n134 36.0641
R116 VTAIL.n17 VTAIL.n16 36.0641
R117 VTAIL.n33 VTAIL.n32 36.0641
R118 VTAIL.n51 VTAIL.n50 36.0641
R119 VTAIL.n119 VTAIL.n118 36.0641
R120 VTAIL.n101 VTAIL.n100 36.0641
R121 VTAIL.n85 VTAIL.n84 36.0641
R122 VTAIL.n67 VTAIL.n66 36.0641
R123 VTAIL.n135 VTAIL.n119 15.91
R124 VTAIL.n67 VTAIL.n51 15.91
R125 VTAIL.n125 VTAIL.n124 15.5966
R126 VTAIL.n7 VTAIL.n6 15.5966
R127 VTAIL.n23 VTAIL.n22 15.5966
R128 VTAIL.n41 VTAIL.n40 15.5966
R129 VTAIL.n109 VTAIL.n108 15.5966
R130 VTAIL.n91 VTAIL.n90 15.5966
R131 VTAIL.n75 VTAIL.n74 15.5966
R132 VTAIL.n57 VTAIL.n56 15.5966
R133 VTAIL.n128 VTAIL.n127 12.8005
R134 VTAIL.n10 VTAIL.n9 12.8005
R135 VTAIL.n26 VTAIL.n25 12.8005
R136 VTAIL.n44 VTAIL.n43 12.8005
R137 VTAIL.n112 VTAIL.n111 12.8005
R138 VTAIL.n94 VTAIL.n93 12.8005
R139 VTAIL.n78 VTAIL.n77 12.8005
R140 VTAIL.n60 VTAIL.n59 12.8005
R141 VTAIL.n131 VTAIL.n122 12.0247
R142 VTAIL.n13 VTAIL.n4 12.0247
R143 VTAIL.n29 VTAIL.n20 12.0247
R144 VTAIL.n47 VTAIL.n38 12.0247
R145 VTAIL.n115 VTAIL.n106 12.0247
R146 VTAIL.n97 VTAIL.n88 12.0247
R147 VTAIL.n81 VTAIL.n72 12.0247
R148 VTAIL.n63 VTAIL.n54 12.0247
R149 VTAIL.n132 VTAIL.n120 11.249
R150 VTAIL.n14 VTAIL.n2 11.249
R151 VTAIL.n30 VTAIL.n18 11.249
R152 VTAIL.n48 VTAIL.n36 11.249
R153 VTAIL.n116 VTAIL.n104 11.249
R154 VTAIL.n98 VTAIL.n86 11.249
R155 VTAIL.n82 VTAIL.n70 11.249
R156 VTAIL.n64 VTAIL.n52 11.249
R157 VTAIL.n134 VTAIL.n133 9.45567
R158 VTAIL.n16 VTAIL.n15 9.45567
R159 VTAIL.n32 VTAIL.n31 9.45567
R160 VTAIL.n50 VTAIL.n49 9.45567
R161 VTAIL.n118 VTAIL.n117 9.45567
R162 VTAIL.n100 VTAIL.n99 9.45567
R163 VTAIL.n84 VTAIL.n83 9.45567
R164 VTAIL.n66 VTAIL.n65 9.45567
R165 VTAIL.n133 VTAIL.n132 9.3005
R166 VTAIL.n122 VTAIL.n121 9.3005
R167 VTAIL.n127 VTAIL.n126 9.3005
R168 VTAIL.n15 VTAIL.n14 9.3005
R169 VTAIL.n4 VTAIL.n3 9.3005
R170 VTAIL.n9 VTAIL.n8 9.3005
R171 VTAIL.n31 VTAIL.n30 9.3005
R172 VTAIL.n20 VTAIL.n19 9.3005
R173 VTAIL.n25 VTAIL.n24 9.3005
R174 VTAIL.n49 VTAIL.n48 9.3005
R175 VTAIL.n38 VTAIL.n37 9.3005
R176 VTAIL.n43 VTAIL.n42 9.3005
R177 VTAIL.n117 VTAIL.n116 9.3005
R178 VTAIL.n106 VTAIL.n105 9.3005
R179 VTAIL.n111 VTAIL.n110 9.3005
R180 VTAIL.n99 VTAIL.n98 9.3005
R181 VTAIL.n88 VTAIL.n87 9.3005
R182 VTAIL.n93 VTAIL.n92 9.3005
R183 VTAIL.n83 VTAIL.n82 9.3005
R184 VTAIL.n72 VTAIL.n71 9.3005
R185 VTAIL.n77 VTAIL.n76 9.3005
R186 VTAIL.n65 VTAIL.n64 9.3005
R187 VTAIL.n54 VTAIL.n53 9.3005
R188 VTAIL.n59 VTAIL.n58 9.3005
R189 VTAIL.n0 VTAIL.t13 5.96436
R190 VTAIL.n0 VTAIL.t2 5.96436
R191 VTAIL.n34 VTAIL.t7 5.96436
R192 VTAIL.n34 VTAIL.t9 5.96436
R193 VTAIL.n102 VTAIL.t8 5.96436
R194 VTAIL.n102 VTAIL.t6 5.96436
R195 VTAIL.n68 VTAIL.t12 5.96436
R196 VTAIL.n68 VTAIL.t11 5.96436
R197 VTAIL.n126 VTAIL.n125 4.46457
R198 VTAIL.n8 VTAIL.n7 4.46457
R199 VTAIL.n24 VTAIL.n23 4.46457
R200 VTAIL.n42 VTAIL.n41 4.46457
R201 VTAIL.n110 VTAIL.n109 4.46457
R202 VTAIL.n92 VTAIL.n91 4.46457
R203 VTAIL.n76 VTAIL.n75 4.46457
R204 VTAIL.n58 VTAIL.n57 4.46457
R205 VTAIL.n134 VTAIL.n120 2.71565
R206 VTAIL.n16 VTAIL.n2 2.71565
R207 VTAIL.n32 VTAIL.n18 2.71565
R208 VTAIL.n50 VTAIL.n36 2.71565
R209 VTAIL.n118 VTAIL.n104 2.71565
R210 VTAIL.n100 VTAIL.n86 2.71565
R211 VTAIL.n84 VTAIL.n70 2.71565
R212 VTAIL.n66 VTAIL.n52 2.71565
R213 VTAIL.n132 VTAIL.n131 1.93989
R214 VTAIL.n14 VTAIL.n13 1.93989
R215 VTAIL.n30 VTAIL.n29 1.93989
R216 VTAIL.n48 VTAIL.n47 1.93989
R217 VTAIL.n116 VTAIL.n115 1.93989
R218 VTAIL.n98 VTAIL.n97 1.93989
R219 VTAIL.n82 VTAIL.n81 1.93989
R220 VTAIL.n64 VTAIL.n63 1.93989
R221 VTAIL.n128 VTAIL.n122 1.16414
R222 VTAIL.n10 VTAIL.n4 1.16414
R223 VTAIL.n26 VTAIL.n20 1.16414
R224 VTAIL.n44 VTAIL.n38 1.16414
R225 VTAIL.n112 VTAIL.n106 1.16414
R226 VTAIL.n94 VTAIL.n88 1.16414
R227 VTAIL.n78 VTAIL.n72 1.16414
R228 VTAIL.n60 VTAIL.n54 1.16414
R229 VTAIL.n69 VTAIL.n67 0.681535
R230 VTAIL.n85 VTAIL.n69 0.681535
R231 VTAIL.n103 VTAIL.n101 0.681535
R232 VTAIL.n119 VTAIL.n103 0.681535
R233 VTAIL.n51 VTAIL.n35 0.681535
R234 VTAIL.n35 VTAIL.n33 0.681535
R235 VTAIL.n17 VTAIL.n1 0.681535
R236 VTAIL VTAIL.n135 0.623345
R237 VTAIL.n101 VTAIL.n85 0.470328
R238 VTAIL.n33 VTAIL.n17 0.470328
R239 VTAIL.n127 VTAIL.n124 0.388379
R240 VTAIL.n9 VTAIL.n6 0.388379
R241 VTAIL.n25 VTAIL.n22 0.388379
R242 VTAIL.n43 VTAIL.n40 0.388379
R243 VTAIL.n111 VTAIL.n108 0.388379
R244 VTAIL.n93 VTAIL.n90 0.388379
R245 VTAIL.n77 VTAIL.n74 0.388379
R246 VTAIL.n59 VTAIL.n56 0.388379
R247 VTAIL.n126 VTAIL.n121 0.155672
R248 VTAIL.n133 VTAIL.n121 0.155672
R249 VTAIL.n8 VTAIL.n3 0.155672
R250 VTAIL.n15 VTAIL.n3 0.155672
R251 VTAIL.n24 VTAIL.n19 0.155672
R252 VTAIL.n31 VTAIL.n19 0.155672
R253 VTAIL.n42 VTAIL.n37 0.155672
R254 VTAIL.n49 VTAIL.n37 0.155672
R255 VTAIL.n117 VTAIL.n105 0.155672
R256 VTAIL.n110 VTAIL.n105 0.155672
R257 VTAIL.n99 VTAIL.n87 0.155672
R258 VTAIL.n92 VTAIL.n87 0.155672
R259 VTAIL.n83 VTAIL.n71 0.155672
R260 VTAIL.n76 VTAIL.n71 0.155672
R261 VTAIL.n65 VTAIL.n53 0.155672
R262 VTAIL.n58 VTAIL.n53 0.155672
R263 VTAIL VTAIL.n1 0.0586897
R264 B.n375 B.n374 585
R265 B.n144 B.n60 585
R266 B.n143 B.n142 585
R267 B.n141 B.n140 585
R268 B.n139 B.n138 585
R269 B.n137 B.n136 585
R270 B.n135 B.n134 585
R271 B.n133 B.n132 585
R272 B.n131 B.n130 585
R273 B.n129 B.n128 585
R274 B.n127 B.n126 585
R275 B.n125 B.n124 585
R276 B.n123 B.n122 585
R277 B.n121 B.n120 585
R278 B.n119 B.n118 585
R279 B.n117 B.n116 585
R280 B.n115 B.n114 585
R281 B.n113 B.n112 585
R282 B.n111 B.n110 585
R283 B.n109 B.n108 585
R284 B.n107 B.n106 585
R285 B.n105 B.n104 585
R286 B.n103 B.n102 585
R287 B.n101 B.n100 585
R288 B.n99 B.n98 585
R289 B.n97 B.n96 585
R290 B.n95 B.n94 585
R291 B.n93 B.n92 585
R292 B.n91 B.n90 585
R293 B.n89 B.n88 585
R294 B.n87 B.n86 585
R295 B.n85 B.n84 585
R296 B.n83 B.n82 585
R297 B.n81 B.n80 585
R298 B.n79 B.n78 585
R299 B.n77 B.n76 585
R300 B.n75 B.n74 585
R301 B.n73 B.n72 585
R302 B.n71 B.n70 585
R303 B.n69 B.n68 585
R304 B.n40 B.n39 585
R305 B.n380 B.n379 585
R306 B.n373 B.n61 585
R307 B.n61 B.n37 585
R308 B.n372 B.n36 585
R309 B.n384 B.n36 585
R310 B.n371 B.n35 585
R311 B.n385 B.n35 585
R312 B.n370 B.n34 585
R313 B.n386 B.n34 585
R314 B.n369 B.n368 585
R315 B.n368 B.n33 585
R316 B.n367 B.n29 585
R317 B.n392 B.n29 585
R318 B.n366 B.n28 585
R319 B.n393 B.n28 585
R320 B.n365 B.n27 585
R321 B.n394 B.n27 585
R322 B.n364 B.n363 585
R323 B.n363 B.n23 585
R324 B.n362 B.n22 585
R325 B.n400 B.n22 585
R326 B.n361 B.n21 585
R327 B.n401 B.n21 585
R328 B.n360 B.n20 585
R329 B.n402 B.n20 585
R330 B.n359 B.n358 585
R331 B.n358 B.n19 585
R332 B.n357 B.n15 585
R333 B.n408 B.n15 585
R334 B.n356 B.n14 585
R335 B.n409 B.n14 585
R336 B.n355 B.n13 585
R337 B.n410 B.n13 585
R338 B.n354 B.n353 585
R339 B.n353 B.n12 585
R340 B.n352 B.n351 585
R341 B.n352 B.n8 585
R342 B.n350 B.n7 585
R343 B.n417 B.n7 585
R344 B.n349 B.n6 585
R345 B.n418 B.n6 585
R346 B.n348 B.n5 585
R347 B.n419 B.n5 585
R348 B.n347 B.n346 585
R349 B.n346 B.n4 585
R350 B.n345 B.n145 585
R351 B.n345 B.n344 585
R352 B.n334 B.n146 585
R353 B.n337 B.n146 585
R354 B.n336 B.n335 585
R355 B.n338 B.n336 585
R356 B.n333 B.n150 585
R357 B.n153 B.n150 585
R358 B.n332 B.n331 585
R359 B.n331 B.n330 585
R360 B.n152 B.n151 585
R361 B.n323 B.n152 585
R362 B.n322 B.n321 585
R363 B.n324 B.n322 585
R364 B.n320 B.n158 585
R365 B.n158 B.n157 585
R366 B.n319 B.n318 585
R367 B.n318 B.n317 585
R368 B.n160 B.n159 585
R369 B.n161 B.n160 585
R370 B.n310 B.n309 585
R371 B.n311 B.n310 585
R372 B.n308 B.n166 585
R373 B.n166 B.n165 585
R374 B.n307 B.n306 585
R375 B.n306 B.n305 585
R376 B.n168 B.n167 585
R377 B.n298 B.n168 585
R378 B.n297 B.n296 585
R379 B.n299 B.n297 585
R380 B.n295 B.n173 585
R381 B.n173 B.n172 585
R382 B.n294 B.n293 585
R383 B.n293 B.n292 585
R384 B.n175 B.n174 585
R385 B.n176 B.n175 585
R386 B.n288 B.n287 585
R387 B.n179 B.n178 585
R388 B.n284 B.n283 585
R389 B.n285 B.n284 585
R390 B.n282 B.n200 585
R391 B.n281 B.n280 585
R392 B.n279 B.n278 585
R393 B.n277 B.n276 585
R394 B.n275 B.n274 585
R395 B.n273 B.n272 585
R396 B.n271 B.n270 585
R397 B.n269 B.n268 585
R398 B.n267 B.n266 585
R399 B.n265 B.n264 585
R400 B.n263 B.n262 585
R401 B.n261 B.n260 585
R402 B.n259 B.n258 585
R403 B.n256 B.n255 585
R404 B.n254 B.n253 585
R405 B.n252 B.n251 585
R406 B.n250 B.n249 585
R407 B.n248 B.n247 585
R408 B.n246 B.n245 585
R409 B.n244 B.n243 585
R410 B.n242 B.n241 585
R411 B.n240 B.n239 585
R412 B.n238 B.n237 585
R413 B.n235 B.n234 585
R414 B.n233 B.n232 585
R415 B.n231 B.n230 585
R416 B.n229 B.n228 585
R417 B.n227 B.n226 585
R418 B.n225 B.n224 585
R419 B.n223 B.n222 585
R420 B.n221 B.n220 585
R421 B.n219 B.n218 585
R422 B.n217 B.n216 585
R423 B.n215 B.n214 585
R424 B.n213 B.n212 585
R425 B.n211 B.n210 585
R426 B.n209 B.n208 585
R427 B.n207 B.n206 585
R428 B.n205 B.n199 585
R429 B.n285 B.n199 585
R430 B.n289 B.n177 585
R431 B.n177 B.n176 585
R432 B.n291 B.n290 585
R433 B.n292 B.n291 585
R434 B.n171 B.n170 585
R435 B.n172 B.n171 585
R436 B.n301 B.n300 585
R437 B.n300 B.n299 585
R438 B.n302 B.n169 585
R439 B.n298 B.n169 585
R440 B.n304 B.n303 585
R441 B.n305 B.n304 585
R442 B.n164 B.n163 585
R443 B.n165 B.n164 585
R444 B.n313 B.n312 585
R445 B.n312 B.n311 585
R446 B.n314 B.n162 585
R447 B.n162 B.n161 585
R448 B.n316 B.n315 585
R449 B.n317 B.n316 585
R450 B.n156 B.n155 585
R451 B.n157 B.n156 585
R452 B.n326 B.n325 585
R453 B.n325 B.n324 585
R454 B.n327 B.n154 585
R455 B.n323 B.n154 585
R456 B.n329 B.n328 585
R457 B.n330 B.n329 585
R458 B.n149 B.n148 585
R459 B.n153 B.n149 585
R460 B.n340 B.n339 585
R461 B.n339 B.n338 585
R462 B.n341 B.n147 585
R463 B.n337 B.n147 585
R464 B.n343 B.n342 585
R465 B.n344 B.n343 585
R466 B.n3 B.n0 585
R467 B.n4 B.n3 585
R468 B.n416 B.n1 585
R469 B.n417 B.n416 585
R470 B.n415 B.n414 585
R471 B.n415 B.n8 585
R472 B.n413 B.n9 585
R473 B.n12 B.n9 585
R474 B.n412 B.n411 585
R475 B.n411 B.n410 585
R476 B.n11 B.n10 585
R477 B.n409 B.n11 585
R478 B.n407 B.n406 585
R479 B.n408 B.n407 585
R480 B.n405 B.n16 585
R481 B.n19 B.n16 585
R482 B.n404 B.n403 585
R483 B.n403 B.n402 585
R484 B.n18 B.n17 585
R485 B.n401 B.n18 585
R486 B.n399 B.n398 585
R487 B.n400 B.n399 585
R488 B.n397 B.n24 585
R489 B.n24 B.n23 585
R490 B.n396 B.n395 585
R491 B.n395 B.n394 585
R492 B.n26 B.n25 585
R493 B.n393 B.n26 585
R494 B.n391 B.n390 585
R495 B.n392 B.n391 585
R496 B.n389 B.n30 585
R497 B.n33 B.n30 585
R498 B.n388 B.n387 585
R499 B.n387 B.n386 585
R500 B.n32 B.n31 585
R501 B.n385 B.n32 585
R502 B.n383 B.n382 585
R503 B.n384 B.n383 585
R504 B.n381 B.n38 585
R505 B.n38 B.n37 585
R506 B.n420 B.n419 585
R507 B.n418 B.n2 585
R508 B.n379 B.n38 516.524
R509 B.n375 B.n61 516.524
R510 B.n199 B.n175 516.524
R511 B.n287 B.n177 516.524
R512 B.n65 B.t16 381.396
R513 B.n62 B.t12 381.396
R514 B.n203 B.t19 381.396
R515 B.n201 B.t8 381.396
R516 B.n377 B.n376 256.663
R517 B.n377 B.n59 256.663
R518 B.n377 B.n58 256.663
R519 B.n377 B.n57 256.663
R520 B.n377 B.n56 256.663
R521 B.n377 B.n55 256.663
R522 B.n377 B.n54 256.663
R523 B.n377 B.n53 256.663
R524 B.n377 B.n52 256.663
R525 B.n377 B.n51 256.663
R526 B.n377 B.n50 256.663
R527 B.n377 B.n49 256.663
R528 B.n377 B.n48 256.663
R529 B.n377 B.n47 256.663
R530 B.n377 B.n46 256.663
R531 B.n377 B.n45 256.663
R532 B.n377 B.n44 256.663
R533 B.n377 B.n43 256.663
R534 B.n377 B.n42 256.663
R535 B.n377 B.n41 256.663
R536 B.n378 B.n377 256.663
R537 B.n286 B.n285 256.663
R538 B.n285 B.n180 256.663
R539 B.n285 B.n181 256.663
R540 B.n285 B.n182 256.663
R541 B.n285 B.n183 256.663
R542 B.n285 B.n184 256.663
R543 B.n285 B.n185 256.663
R544 B.n285 B.n186 256.663
R545 B.n285 B.n187 256.663
R546 B.n285 B.n188 256.663
R547 B.n285 B.n189 256.663
R548 B.n285 B.n190 256.663
R549 B.n285 B.n191 256.663
R550 B.n285 B.n192 256.663
R551 B.n285 B.n193 256.663
R552 B.n285 B.n194 256.663
R553 B.n285 B.n195 256.663
R554 B.n285 B.n196 256.663
R555 B.n285 B.n197 256.663
R556 B.n285 B.n198 256.663
R557 B.n422 B.n421 256.663
R558 B.n285 B.n176 177.894
R559 B.n377 B.n37 177.894
R560 B.n68 B.n40 163.367
R561 B.n72 B.n71 163.367
R562 B.n76 B.n75 163.367
R563 B.n80 B.n79 163.367
R564 B.n84 B.n83 163.367
R565 B.n88 B.n87 163.367
R566 B.n92 B.n91 163.367
R567 B.n96 B.n95 163.367
R568 B.n100 B.n99 163.367
R569 B.n104 B.n103 163.367
R570 B.n108 B.n107 163.367
R571 B.n112 B.n111 163.367
R572 B.n116 B.n115 163.367
R573 B.n120 B.n119 163.367
R574 B.n124 B.n123 163.367
R575 B.n128 B.n127 163.367
R576 B.n132 B.n131 163.367
R577 B.n136 B.n135 163.367
R578 B.n140 B.n139 163.367
R579 B.n142 B.n60 163.367
R580 B.n293 B.n175 163.367
R581 B.n293 B.n173 163.367
R582 B.n297 B.n173 163.367
R583 B.n297 B.n168 163.367
R584 B.n306 B.n168 163.367
R585 B.n306 B.n166 163.367
R586 B.n310 B.n166 163.367
R587 B.n310 B.n160 163.367
R588 B.n318 B.n160 163.367
R589 B.n318 B.n158 163.367
R590 B.n322 B.n158 163.367
R591 B.n322 B.n152 163.367
R592 B.n331 B.n152 163.367
R593 B.n331 B.n150 163.367
R594 B.n336 B.n150 163.367
R595 B.n336 B.n146 163.367
R596 B.n345 B.n146 163.367
R597 B.n346 B.n345 163.367
R598 B.n346 B.n5 163.367
R599 B.n6 B.n5 163.367
R600 B.n7 B.n6 163.367
R601 B.n352 B.n7 163.367
R602 B.n353 B.n352 163.367
R603 B.n353 B.n13 163.367
R604 B.n14 B.n13 163.367
R605 B.n15 B.n14 163.367
R606 B.n358 B.n15 163.367
R607 B.n358 B.n20 163.367
R608 B.n21 B.n20 163.367
R609 B.n22 B.n21 163.367
R610 B.n363 B.n22 163.367
R611 B.n363 B.n27 163.367
R612 B.n28 B.n27 163.367
R613 B.n29 B.n28 163.367
R614 B.n368 B.n29 163.367
R615 B.n368 B.n34 163.367
R616 B.n35 B.n34 163.367
R617 B.n36 B.n35 163.367
R618 B.n61 B.n36 163.367
R619 B.n284 B.n179 163.367
R620 B.n284 B.n200 163.367
R621 B.n280 B.n279 163.367
R622 B.n276 B.n275 163.367
R623 B.n272 B.n271 163.367
R624 B.n268 B.n267 163.367
R625 B.n264 B.n263 163.367
R626 B.n260 B.n259 163.367
R627 B.n255 B.n254 163.367
R628 B.n251 B.n250 163.367
R629 B.n247 B.n246 163.367
R630 B.n243 B.n242 163.367
R631 B.n239 B.n238 163.367
R632 B.n234 B.n233 163.367
R633 B.n230 B.n229 163.367
R634 B.n226 B.n225 163.367
R635 B.n222 B.n221 163.367
R636 B.n218 B.n217 163.367
R637 B.n214 B.n213 163.367
R638 B.n210 B.n209 163.367
R639 B.n206 B.n199 163.367
R640 B.n291 B.n177 163.367
R641 B.n291 B.n171 163.367
R642 B.n300 B.n171 163.367
R643 B.n300 B.n169 163.367
R644 B.n304 B.n169 163.367
R645 B.n304 B.n164 163.367
R646 B.n312 B.n164 163.367
R647 B.n312 B.n162 163.367
R648 B.n316 B.n162 163.367
R649 B.n316 B.n156 163.367
R650 B.n325 B.n156 163.367
R651 B.n325 B.n154 163.367
R652 B.n329 B.n154 163.367
R653 B.n329 B.n149 163.367
R654 B.n339 B.n149 163.367
R655 B.n339 B.n147 163.367
R656 B.n343 B.n147 163.367
R657 B.n343 B.n3 163.367
R658 B.n420 B.n3 163.367
R659 B.n416 B.n2 163.367
R660 B.n416 B.n415 163.367
R661 B.n415 B.n9 163.367
R662 B.n411 B.n9 163.367
R663 B.n411 B.n11 163.367
R664 B.n407 B.n11 163.367
R665 B.n407 B.n16 163.367
R666 B.n403 B.n16 163.367
R667 B.n403 B.n18 163.367
R668 B.n399 B.n18 163.367
R669 B.n399 B.n24 163.367
R670 B.n395 B.n24 163.367
R671 B.n395 B.n26 163.367
R672 B.n391 B.n26 163.367
R673 B.n391 B.n30 163.367
R674 B.n387 B.n30 163.367
R675 B.n387 B.n32 163.367
R676 B.n383 B.n32 163.367
R677 B.n383 B.n38 163.367
R678 B.n62 B.t14 149.827
R679 B.n203 B.t21 149.827
R680 B.n65 B.t17 149.827
R681 B.n201 B.t11 149.827
R682 B.n63 B.t15 134.506
R683 B.n204 B.t20 134.506
R684 B.n66 B.t18 134.506
R685 B.n202 B.t10 134.506
R686 B.n292 B.n176 87.0278
R687 B.n292 B.n172 87.0278
R688 B.n299 B.n172 87.0278
R689 B.n299 B.n298 87.0278
R690 B.n305 B.n165 87.0278
R691 B.n311 B.n165 87.0278
R692 B.n311 B.n161 87.0278
R693 B.n317 B.n161 87.0278
R694 B.n324 B.n157 87.0278
R695 B.n324 B.n323 87.0278
R696 B.n330 B.n153 87.0278
R697 B.n338 B.n337 87.0278
R698 B.n344 B.n4 87.0278
R699 B.n419 B.n4 87.0278
R700 B.n419 B.n418 87.0278
R701 B.n418 B.n417 87.0278
R702 B.n417 B.n8 87.0278
R703 B.n410 B.n12 87.0278
R704 B.n409 B.n408 87.0278
R705 B.n402 B.n19 87.0278
R706 B.n402 B.n401 87.0278
R707 B.n400 B.n23 87.0278
R708 B.n394 B.n23 87.0278
R709 B.n394 B.n393 87.0278
R710 B.n393 B.n392 87.0278
R711 B.n386 B.n33 87.0278
R712 B.n386 B.n385 87.0278
R713 B.n385 B.n384 87.0278
R714 B.n384 B.n37 87.0278
R715 B.n330 B.t5 79.349
R716 B.n408 B.t2 79.349
R717 B.n379 B.n378 71.676
R718 B.n68 B.n41 71.676
R719 B.n72 B.n42 71.676
R720 B.n76 B.n43 71.676
R721 B.n80 B.n44 71.676
R722 B.n84 B.n45 71.676
R723 B.n88 B.n46 71.676
R724 B.n92 B.n47 71.676
R725 B.n96 B.n48 71.676
R726 B.n100 B.n49 71.676
R727 B.n104 B.n50 71.676
R728 B.n108 B.n51 71.676
R729 B.n112 B.n52 71.676
R730 B.n116 B.n53 71.676
R731 B.n120 B.n54 71.676
R732 B.n124 B.n55 71.676
R733 B.n128 B.n56 71.676
R734 B.n132 B.n57 71.676
R735 B.n136 B.n58 71.676
R736 B.n140 B.n59 71.676
R737 B.n376 B.n60 71.676
R738 B.n376 B.n375 71.676
R739 B.n142 B.n59 71.676
R740 B.n139 B.n58 71.676
R741 B.n135 B.n57 71.676
R742 B.n131 B.n56 71.676
R743 B.n127 B.n55 71.676
R744 B.n123 B.n54 71.676
R745 B.n119 B.n53 71.676
R746 B.n115 B.n52 71.676
R747 B.n111 B.n51 71.676
R748 B.n107 B.n50 71.676
R749 B.n103 B.n49 71.676
R750 B.n99 B.n48 71.676
R751 B.n95 B.n47 71.676
R752 B.n91 B.n46 71.676
R753 B.n87 B.n45 71.676
R754 B.n83 B.n44 71.676
R755 B.n79 B.n43 71.676
R756 B.n75 B.n42 71.676
R757 B.n71 B.n41 71.676
R758 B.n378 B.n40 71.676
R759 B.n287 B.n286 71.676
R760 B.n200 B.n180 71.676
R761 B.n279 B.n181 71.676
R762 B.n275 B.n182 71.676
R763 B.n271 B.n183 71.676
R764 B.n267 B.n184 71.676
R765 B.n263 B.n185 71.676
R766 B.n259 B.n186 71.676
R767 B.n254 B.n187 71.676
R768 B.n250 B.n188 71.676
R769 B.n246 B.n189 71.676
R770 B.n242 B.n190 71.676
R771 B.n238 B.n191 71.676
R772 B.n233 B.n192 71.676
R773 B.n229 B.n193 71.676
R774 B.n225 B.n194 71.676
R775 B.n221 B.n195 71.676
R776 B.n217 B.n196 71.676
R777 B.n213 B.n197 71.676
R778 B.n209 B.n198 71.676
R779 B.n286 B.n179 71.676
R780 B.n280 B.n180 71.676
R781 B.n276 B.n181 71.676
R782 B.n272 B.n182 71.676
R783 B.n268 B.n183 71.676
R784 B.n264 B.n184 71.676
R785 B.n260 B.n185 71.676
R786 B.n255 B.n186 71.676
R787 B.n251 B.n187 71.676
R788 B.n247 B.n188 71.676
R789 B.n243 B.n189 71.676
R790 B.n239 B.n190 71.676
R791 B.n234 B.n191 71.676
R792 B.n230 B.n192 71.676
R793 B.n226 B.n193 71.676
R794 B.n222 B.n194 71.676
R795 B.n218 B.n195 71.676
R796 B.n214 B.n196 71.676
R797 B.n210 B.n197 71.676
R798 B.n206 B.n198 71.676
R799 B.n421 B.n420 71.676
R800 B.n421 B.n2 71.676
R801 B.n305 B.t9 66.5508
R802 B.n317 B.t1 66.5508
R803 B.t4 B.n400 66.5508
R804 B.n392 B.t13 66.5508
R805 B.n337 B.t3 63.9912
R806 B.n12 B.t0 63.9912
R807 B.n67 B.n66 59.5399
R808 B.n64 B.n63 59.5399
R809 B.n236 B.n204 59.5399
R810 B.n257 B.n202 59.5399
R811 B.n338 B.t7 51.1931
R812 B.n410 B.t6 51.1931
R813 B.n153 B.t7 35.8353
R814 B.t6 B.n409 35.8353
R815 B.n289 B.n288 33.5615
R816 B.n205 B.n174 33.5615
R817 B.n374 B.n373 33.5615
R818 B.n381 B.n380 33.5615
R819 B.n344 B.t3 23.0371
R820 B.t0 B.n8 23.0371
R821 B.n298 B.t9 20.4775
R822 B.t1 B.n157 20.4775
R823 B.n401 B.t4 20.4775
R824 B.n33 B.t13 20.4775
R825 B B.n422 18.0485
R826 B.n66 B.n65 15.3217
R827 B.n63 B.n62 15.3217
R828 B.n204 B.n203 15.3217
R829 B.n202 B.n201 15.3217
R830 B.n290 B.n289 10.6151
R831 B.n290 B.n170 10.6151
R832 B.n301 B.n170 10.6151
R833 B.n302 B.n301 10.6151
R834 B.n303 B.n302 10.6151
R835 B.n303 B.n163 10.6151
R836 B.n313 B.n163 10.6151
R837 B.n314 B.n313 10.6151
R838 B.n315 B.n314 10.6151
R839 B.n315 B.n155 10.6151
R840 B.n326 B.n155 10.6151
R841 B.n327 B.n326 10.6151
R842 B.n328 B.n327 10.6151
R843 B.n328 B.n148 10.6151
R844 B.n340 B.n148 10.6151
R845 B.n341 B.n340 10.6151
R846 B.n342 B.n341 10.6151
R847 B.n342 B.n0 10.6151
R848 B.n288 B.n178 10.6151
R849 B.n283 B.n178 10.6151
R850 B.n283 B.n282 10.6151
R851 B.n282 B.n281 10.6151
R852 B.n281 B.n278 10.6151
R853 B.n278 B.n277 10.6151
R854 B.n277 B.n274 10.6151
R855 B.n274 B.n273 10.6151
R856 B.n273 B.n270 10.6151
R857 B.n270 B.n269 10.6151
R858 B.n269 B.n266 10.6151
R859 B.n266 B.n265 10.6151
R860 B.n265 B.n262 10.6151
R861 B.n262 B.n261 10.6151
R862 B.n261 B.n258 10.6151
R863 B.n256 B.n253 10.6151
R864 B.n253 B.n252 10.6151
R865 B.n252 B.n249 10.6151
R866 B.n249 B.n248 10.6151
R867 B.n248 B.n245 10.6151
R868 B.n245 B.n244 10.6151
R869 B.n244 B.n241 10.6151
R870 B.n241 B.n240 10.6151
R871 B.n240 B.n237 10.6151
R872 B.n235 B.n232 10.6151
R873 B.n232 B.n231 10.6151
R874 B.n231 B.n228 10.6151
R875 B.n228 B.n227 10.6151
R876 B.n227 B.n224 10.6151
R877 B.n224 B.n223 10.6151
R878 B.n223 B.n220 10.6151
R879 B.n220 B.n219 10.6151
R880 B.n219 B.n216 10.6151
R881 B.n216 B.n215 10.6151
R882 B.n215 B.n212 10.6151
R883 B.n212 B.n211 10.6151
R884 B.n211 B.n208 10.6151
R885 B.n208 B.n207 10.6151
R886 B.n207 B.n205 10.6151
R887 B.n294 B.n174 10.6151
R888 B.n295 B.n294 10.6151
R889 B.n296 B.n295 10.6151
R890 B.n296 B.n167 10.6151
R891 B.n307 B.n167 10.6151
R892 B.n308 B.n307 10.6151
R893 B.n309 B.n308 10.6151
R894 B.n309 B.n159 10.6151
R895 B.n319 B.n159 10.6151
R896 B.n320 B.n319 10.6151
R897 B.n321 B.n320 10.6151
R898 B.n321 B.n151 10.6151
R899 B.n332 B.n151 10.6151
R900 B.n333 B.n332 10.6151
R901 B.n335 B.n333 10.6151
R902 B.n335 B.n334 10.6151
R903 B.n334 B.n145 10.6151
R904 B.n347 B.n145 10.6151
R905 B.n348 B.n347 10.6151
R906 B.n349 B.n348 10.6151
R907 B.n350 B.n349 10.6151
R908 B.n351 B.n350 10.6151
R909 B.n354 B.n351 10.6151
R910 B.n355 B.n354 10.6151
R911 B.n356 B.n355 10.6151
R912 B.n357 B.n356 10.6151
R913 B.n359 B.n357 10.6151
R914 B.n360 B.n359 10.6151
R915 B.n361 B.n360 10.6151
R916 B.n362 B.n361 10.6151
R917 B.n364 B.n362 10.6151
R918 B.n365 B.n364 10.6151
R919 B.n366 B.n365 10.6151
R920 B.n367 B.n366 10.6151
R921 B.n369 B.n367 10.6151
R922 B.n370 B.n369 10.6151
R923 B.n371 B.n370 10.6151
R924 B.n372 B.n371 10.6151
R925 B.n373 B.n372 10.6151
R926 B.n414 B.n1 10.6151
R927 B.n414 B.n413 10.6151
R928 B.n413 B.n412 10.6151
R929 B.n412 B.n10 10.6151
R930 B.n406 B.n10 10.6151
R931 B.n406 B.n405 10.6151
R932 B.n405 B.n404 10.6151
R933 B.n404 B.n17 10.6151
R934 B.n398 B.n17 10.6151
R935 B.n398 B.n397 10.6151
R936 B.n397 B.n396 10.6151
R937 B.n396 B.n25 10.6151
R938 B.n390 B.n25 10.6151
R939 B.n390 B.n389 10.6151
R940 B.n389 B.n388 10.6151
R941 B.n388 B.n31 10.6151
R942 B.n382 B.n31 10.6151
R943 B.n382 B.n381 10.6151
R944 B.n380 B.n39 10.6151
R945 B.n69 B.n39 10.6151
R946 B.n70 B.n69 10.6151
R947 B.n73 B.n70 10.6151
R948 B.n74 B.n73 10.6151
R949 B.n77 B.n74 10.6151
R950 B.n78 B.n77 10.6151
R951 B.n81 B.n78 10.6151
R952 B.n82 B.n81 10.6151
R953 B.n85 B.n82 10.6151
R954 B.n86 B.n85 10.6151
R955 B.n89 B.n86 10.6151
R956 B.n90 B.n89 10.6151
R957 B.n93 B.n90 10.6151
R958 B.n94 B.n93 10.6151
R959 B.n98 B.n97 10.6151
R960 B.n101 B.n98 10.6151
R961 B.n102 B.n101 10.6151
R962 B.n105 B.n102 10.6151
R963 B.n106 B.n105 10.6151
R964 B.n109 B.n106 10.6151
R965 B.n110 B.n109 10.6151
R966 B.n113 B.n110 10.6151
R967 B.n114 B.n113 10.6151
R968 B.n118 B.n117 10.6151
R969 B.n121 B.n118 10.6151
R970 B.n122 B.n121 10.6151
R971 B.n125 B.n122 10.6151
R972 B.n126 B.n125 10.6151
R973 B.n129 B.n126 10.6151
R974 B.n130 B.n129 10.6151
R975 B.n133 B.n130 10.6151
R976 B.n134 B.n133 10.6151
R977 B.n137 B.n134 10.6151
R978 B.n138 B.n137 10.6151
R979 B.n141 B.n138 10.6151
R980 B.n143 B.n141 10.6151
R981 B.n144 B.n143 10.6151
R982 B.n374 B.n144 10.6151
R983 B.n258 B.n257 9.36635
R984 B.n236 B.n235 9.36635
R985 B.n94 B.n67 9.36635
R986 B.n117 B.n64 9.36635
R987 B.n422 B.n0 8.11757
R988 B.n422 B.n1 8.11757
R989 B.n323 B.t5 7.67938
R990 B.n19 B.t2 7.67938
R991 B.n257 B.n256 1.24928
R992 B.n237 B.n236 1.24928
R993 B.n97 B.n67 1.24928
R994 B.n114 B.n64 1.24928
R995 VN.n2 VN.t5 280.32
R996 VN.n10 VN.t3 280.32
R997 VN.n1 VN.t6 259.337
R998 VN.n5 VN.t0 259.337
R999 VN.n6 VN.t7 259.337
R1000 VN.n9 VN.t4 259.337
R1001 VN.n13 VN.t1 259.337
R1002 VN.n14 VN.t2 259.337
R1003 VN.n7 VN.n6 161.3
R1004 VN.n15 VN.n14 161.3
R1005 VN.n13 VN.n8 161.3
R1006 VN.n12 VN.n11 161.3
R1007 VN.n5 VN.n0 161.3
R1008 VN.n4 VN.n3 161.3
R1009 VN.n11 VN.n10 70.4033
R1010 VN.n3 VN.n2 70.4033
R1011 VN.n6 VN.n5 48.2005
R1012 VN.n14 VN.n13 48.2005
R1013 VN VN.n15 34.7221
R1014 VN.n4 VN.n1 24.1005
R1015 VN.n5 VN.n4 24.1005
R1016 VN.n13 VN.n12 24.1005
R1017 VN.n12 VN.n9 24.1005
R1018 VN.n10 VN.n9 20.9576
R1019 VN.n2 VN.n1 20.9576
R1020 VN.n15 VN.n8 0.189894
R1021 VN.n11 VN.n8 0.189894
R1022 VN.n3 VN.n0 0.189894
R1023 VN.n7 VN.n0 0.189894
R1024 VN VN.n7 0.0516364
R1025 VDD2.n2 VDD2.n1 81.913
R1026 VDD2.n2 VDD2.n0 81.913
R1027 VDD2 VDD2.n5 81.9102
R1028 VDD2.n4 VDD2.n3 81.628
R1029 VDD2.n4 VDD2.n2 29.642
R1030 VDD2.n5 VDD2.t3 5.96436
R1031 VDD2.n5 VDD2.t4 5.96436
R1032 VDD2.n3 VDD2.t5 5.96436
R1033 VDD2.n3 VDD2.t6 5.96436
R1034 VDD2.n1 VDD2.t7 5.96436
R1035 VDD2.n1 VDD2.t0 5.96436
R1036 VDD2.n0 VDD2.t2 5.96436
R1037 VDD2.n0 VDD2.t1 5.96436
R1038 VDD2 VDD2.n4 0.399207
C0 VP VDD2 0.297488f
C1 VN VP 3.44175f
C2 VN VDD2 1.46589f
C3 VTAIL VP 1.56471f
C4 VDD1 VP 1.60967f
C5 VTAIL VDD2 5.13771f
C6 VDD1 VDD2 0.709053f
C7 VN VTAIL 1.5506f
C8 VDD1 VN 0.152957f
C9 VDD1 VTAIL 5.09764f
C10 VDD2 B 2.472439f
C11 VDD1 B 2.675775f
C12 VTAIL B 3.709781f
C13 VN B 5.890039f
C14 VP B 4.980482f
C15 VDD2.t2 B 0.057313f
C16 VDD2.t1 B 0.057313f
C17 VDD2.n0 B 0.43412f
C18 VDD2.t7 B 0.057313f
C19 VDD2.t0 B 0.057313f
C20 VDD2.n1 B 0.43412f
C21 VDD2.n2 B 1.30539f
C22 VDD2.t5 B 0.057313f
C23 VDD2.t6 B 0.057313f
C24 VDD2.n3 B 0.433265f
C25 VDD2.n4 B 1.30911f
C26 VDD2.t3 B 0.057313f
C27 VDD2.t4 B 0.057313f
C28 VDD2.n5 B 0.434105f
C29 VN.n0 B 0.026844f
C30 VN.t6 B 0.122158f
C31 VN.n1 B 0.073535f
C32 VN.t5 B 0.12746f
C33 VN.n2 B 0.065698f
C34 VN.n3 B 0.085797f
C35 VN.n4 B 0.006091f
C36 VN.t0 B 0.122158f
C37 VN.n5 B 0.073535f
C38 VN.t7 B 0.122158f
C39 VN.n6 B 0.070804f
C40 VN.n7 B 0.020803f
C41 VN.n8 B 0.026844f
C42 VN.t4 B 0.122158f
C43 VN.n9 B 0.073535f
C44 VN.t3 B 0.12746f
C45 VN.n10 B 0.065698f
C46 VN.n11 B 0.085797f
C47 VN.n12 B 0.006091f
C48 VN.t1 B 0.122158f
C49 VN.n13 B 0.073535f
C50 VN.t2 B 0.122158f
C51 VN.n14 B 0.070804f
C52 VN.n15 B 0.788675f
C53 VTAIL.t13 B 0.050189f
C54 VTAIL.t2 B 0.050189f
C55 VTAIL.n0 B 0.342639f
C56 VTAIL.n1 B 0.203166f
C57 VTAIL.n2 B 0.027406f
C58 VTAIL.n3 B 0.01913f
C59 VTAIL.n4 B 0.01028f
C60 VTAIL.n5 B 0.018223f
C61 VTAIL.n6 B 0.014168f
C62 VTAIL.t0 B 0.041441f
C63 VTAIL.n7 B 0.072243f
C64 VTAIL.n8 B 0.215156f
C65 VTAIL.n9 B 0.01028f
C66 VTAIL.n10 B 0.010885f
C67 VTAIL.n11 B 0.024298f
C68 VTAIL.n12 B 0.053513f
C69 VTAIL.n13 B 0.010885f
C70 VTAIL.n14 B 0.01028f
C71 VTAIL.n15 B 0.049445f
C72 VTAIL.n16 B 0.030189f
C73 VTAIL.n17 B 0.090238f
C74 VTAIL.n18 B 0.027406f
C75 VTAIL.n19 B 0.01913f
C76 VTAIL.n20 B 0.01028f
C77 VTAIL.n21 B 0.018223f
C78 VTAIL.n22 B 0.014168f
C79 VTAIL.t3 B 0.041441f
C80 VTAIL.n23 B 0.072243f
C81 VTAIL.n24 B 0.215156f
C82 VTAIL.n25 B 0.01028f
C83 VTAIL.n26 B 0.010885f
C84 VTAIL.n27 B 0.024298f
C85 VTAIL.n28 B 0.053513f
C86 VTAIL.n29 B 0.010885f
C87 VTAIL.n30 B 0.01028f
C88 VTAIL.n31 B 0.049445f
C89 VTAIL.n32 B 0.030189f
C90 VTAIL.n33 B 0.090238f
C91 VTAIL.t7 B 0.050189f
C92 VTAIL.t9 B 0.050189f
C93 VTAIL.n34 B 0.342639f
C94 VTAIL.n35 B 0.241559f
C95 VTAIL.n36 B 0.027406f
C96 VTAIL.n37 B 0.01913f
C97 VTAIL.n38 B 0.01028f
C98 VTAIL.n39 B 0.018223f
C99 VTAIL.n40 B 0.014168f
C100 VTAIL.t10 B 0.041441f
C101 VTAIL.n41 B 0.072243f
C102 VTAIL.n42 B 0.215156f
C103 VTAIL.n43 B 0.01028f
C104 VTAIL.n44 B 0.010885f
C105 VTAIL.n45 B 0.024298f
C106 VTAIL.n46 B 0.053513f
C107 VTAIL.n47 B 0.010885f
C108 VTAIL.n48 B 0.01028f
C109 VTAIL.n49 B 0.049445f
C110 VTAIL.n50 B 0.030189f
C111 VTAIL.n51 B 0.539543f
C112 VTAIL.n52 B 0.027406f
C113 VTAIL.n53 B 0.01913f
C114 VTAIL.n54 B 0.01028f
C115 VTAIL.n55 B 0.018223f
C116 VTAIL.n56 B 0.014168f
C117 VTAIL.t1 B 0.041441f
C118 VTAIL.n57 B 0.072243f
C119 VTAIL.n58 B 0.215156f
C120 VTAIL.n59 B 0.01028f
C121 VTAIL.n60 B 0.010885f
C122 VTAIL.n61 B 0.024298f
C123 VTAIL.n62 B 0.053513f
C124 VTAIL.n63 B 0.010885f
C125 VTAIL.n64 B 0.01028f
C126 VTAIL.n65 B 0.049445f
C127 VTAIL.n66 B 0.030189f
C128 VTAIL.n67 B 0.539543f
C129 VTAIL.t12 B 0.050189f
C130 VTAIL.t11 B 0.050189f
C131 VTAIL.n68 B 0.342641f
C132 VTAIL.n69 B 0.241557f
C133 VTAIL.n70 B 0.027406f
C134 VTAIL.n71 B 0.01913f
C135 VTAIL.n72 B 0.01028f
C136 VTAIL.n73 B 0.018223f
C137 VTAIL.n74 B 0.014168f
C138 VTAIL.t15 B 0.041441f
C139 VTAIL.n75 B 0.072243f
C140 VTAIL.n76 B 0.215156f
C141 VTAIL.n77 B 0.01028f
C142 VTAIL.n78 B 0.010885f
C143 VTAIL.n79 B 0.024298f
C144 VTAIL.n80 B 0.053513f
C145 VTAIL.n81 B 0.010885f
C146 VTAIL.n82 B 0.01028f
C147 VTAIL.n83 B 0.049445f
C148 VTAIL.n84 B 0.030189f
C149 VTAIL.n85 B 0.090238f
C150 VTAIL.n86 B 0.027406f
C151 VTAIL.n87 B 0.01913f
C152 VTAIL.n88 B 0.01028f
C153 VTAIL.n89 B 0.018223f
C154 VTAIL.n90 B 0.014168f
C155 VTAIL.t4 B 0.041441f
C156 VTAIL.n91 B 0.072243f
C157 VTAIL.n92 B 0.215156f
C158 VTAIL.n93 B 0.01028f
C159 VTAIL.n94 B 0.010885f
C160 VTAIL.n95 B 0.024298f
C161 VTAIL.n96 B 0.053513f
C162 VTAIL.n97 B 0.010885f
C163 VTAIL.n98 B 0.01028f
C164 VTAIL.n99 B 0.049445f
C165 VTAIL.n100 B 0.030189f
C166 VTAIL.n101 B 0.090238f
C167 VTAIL.t8 B 0.050189f
C168 VTAIL.t6 B 0.050189f
C169 VTAIL.n102 B 0.342641f
C170 VTAIL.n103 B 0.241557f
C171 VTAIL.n104 B 0.027406f
C172 VTAIL.n105 B 0.01913f
C173 VTAIL.n106 B 0.01028f
C174 VTAIL.n107 B 0.018223f
C175 VTAIL.n108 B 0.014168f
C176 VTAIL.t5 B 0.041441f
C177 VTAIL.n109 B 0.072243f
C178 VTAIL.n110 B 0.215156f
C179 VTAIL.n111 B 0.01028f
C180 VTAIL.n112 B 0.010885f
C181 VTAIL.n113 B 0.024298f
C182 VTAIL.n114 B 0.053513f
C183 VTAIL.n115 B 0.010885f
C184 VTAIL.n116 B 0.01028f
C185 VTAIL.n117 B 0.049445f
C186 VTAIL.n118 B 0.030189f
C187 VTAIL.n119 B 0.539543f
C188 VTAIL.n120 B 0.027406f
C189 VTAIL.n121 B 0.01913f
C190 VTAIL.n122 B 0.01028f
C191 VTAIL.n123 B 0.018223f
C192 VTAIL.n124 B 0.014168f
C193 VTAIL.t14 B 0.041441f
C194 VTAIL.n125 B 0.072243f
C195 VTAIL.n126 B 0.215156f
C196 VTAIL.n127 B 0.01028f
C197 VTAIL.n128 B 0.010885f
C198 VTAIL.n129 B 0.024298f
C199 VTAIL.n130 B 0.053513f
C200 VTAIL.n131 B 0.010885f
C201 VTAIL.n132 B 0.01028f
C202 VTAIL.n133 B 0.049445f
C203 VTAIL.n134 B 0.030189f
C204 VTAIL.n135 B 0.535956f
C205 VDD1.t5 B 0.056421f
C206 VDD1.t2 B 0.056421f
C207 VDD1.n0 B 0.427725f
C208 VDD1.t6 B 0.056421f
C209 VDD1.t7 B 0.056421f
C210 VDD1.n1 B 0.427359f
C211 VDD1.t3 B 0.056421f
C212 VDD1.t1 B 0.056421f
C213 VDD1.n2 B 0.427359f
C214 VDD1.n3 B 1.33133f
C215 VDD1.t4 B 0.056421f
C216 VDD1.t0 B 0.056421f
C217 VDD1.n4 B 0.426515f
C218 VDD1.n5 B 1.31382f
C219 VP.n0 B 0.027145f
C220 VP.t3 B 0.123529f
C221 VP.n1 B 0.07436f
C222 VP.n2 B 0.027145f
C223 VP.t5 B 0.123529f
C224 VP.t4 B 0.123529f
C225 VP.t2 B 0.123529f
C226 VP.n3 B 0.07436f
C227 VP.t6 B 0.128891f
C228 VP.n4 B 0.066436f
C229 VP.n5 B 0.08676f
C230 VP.n6 B 0.00616f
C231 VP.n7 B 0.07436f
C232 VP.n8 B 0.071599f
C233 VP.n9 B 0.779457f
C234 VP.t0 B 0.123529f
C235 VP.n10 B 0.071599f
C236 VP.n11 B 0.807953f
C237 VP.n12 B 0.027145f
C238 VP.n13 B 0.027145f
C239 VP.n14 B 0.00616f
C240 VP.t1 B 0.123529f
C241 VP.n15 B 0.07436f
C242 VP.t7 B 0.123529f
C243 VP.n16 B 0.071599f
C244 VP.n17 B 0.021037f
.ends

