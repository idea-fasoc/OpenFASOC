* NGSPICE file created from diff_pair_sample_1319.ext - technology: sky130A

.subckt diff_pair_sample_1319 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=1.1427 ps=6.64 w=2.93 l=2.06
X1 B.t11 B.t9 B.t10 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=0 ps=0 w=2.93 l=2.06
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=1.1427 ps=6.64 w=2.93 l=2.06
X3 B.t8 B.t6 B.t7 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=0 ps=0 w=2.93 l=2.06
X4 VDD2.t1 VN.t0 VTAIL.t0 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=1.1427 ps=6.64 w=2.93 l=2.06
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=1.1427 ps=6.64 w=2.93 l=2.06
X6 B.t5 B.t3 B.t4 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=0 ps=0 w=2.93 l=2.06
X7 B.t2 B.t0 B.t1 w_n1926_n1554# sky130_fd_pr__pfet_01v8 ad=1.1427 pd=6.64 as=0 ps=0 w=2.93 l=2.06
R0 VP.n0 VP.t1 129.493
R1 VP.n0 VP.t0 93.1394
R2 VP VP.n0 0.241678
R3 VTAIL.n1 VTAIL.t0 135.782
R4 VTAIL.n3 VTAIL.t1 135.781
R5 VTAIL.n0 VTAIL.t3 135.781
R6 VTAIL.n2 VTAIL.t2 135.781
R7 VTAIL.n1 VTAIL.n0 19.0134
R8 VTAIL.n3 VTAIL.n2 16.9531
R9 VTAIL.n2 VTAIL.n1 1.5005
R10 VTAIL VTAIL.n0 1.0436
R11 VTAIL VTAIL.n3 0.457397
R12 VDD1 VDD1.t1 183.806
R13 VDD1 VDD1.t0 153.035
R14 B.n254 B.n37 585
R15 B.n256 B.n255 585
R16 B.n257 B.n36 585
R17 B.n259 B.n258 585
R18 B.n260 B.n35 585
R19 B.n262 B.n261 585
R20 B.n263 B.n34 585
R21 B.n265 B.n264 585
R22 B.n266 B.n33 585
R23 B.n268 B.n267 585
R24 B.n269 B.n32 585
R25 B.n271 B.n270 585
R26 B.n272 B.n31 585
R27 B.n274 B.n273 585
R28 B.n275 B.n28 585
R29 B.n278 B.n277 585
R30 B.n279 B.n27 585
R31 B.n281 B.n280 585
R32 B.n282 B.n26 585
R33 B.n284 B.n283 585
R34 B.n285 B.n25 585
R35 B.n287 B.n286 585
R36 B.n288 B.n21 585
R37 B.n290 B.n289 585
R38 B.n291 B.n20 585
R39 B.n293 B.n292 585
R40 B.n294 B.n19 585
R41 B.n296 B.n295 585
R42 B.n297 B.n18 585
R43 B.n299 B.n298 585
R44 B.n300 B.n17 585
R45 B.n302 B.n301 585
R46 B.n303 B.n16 585
R47 B.n305 B.n304 585
R48 B.n306 B.n15 585
R49 B.n308 B.n307 585
R50 B.n309 B.n14 585
R51 B.n311 B.n310 585
R52 B.n312 B.n13 585
R53 B.n253 B.n252 585
R54 B.n251 B.n38 585
R55 B.n250 B.n249 585
R56 B.n248 B.n39 585
R57 B.n247 B.n246 585
R58 B.n245 B.n40 585
R59 B.n244 B.n243 585
R60 B.n242 B.n41 585
R61 B.n241 B.n240 585
R62 B.n239 B.n42 585
R63 B.n238 B.n237 585
R64 B.n236 B.n43 585
R65 B.n235 B.n234 585
R66 B.n233 B.n44 585
R67 B.n232 B.n231 585
R68 B.n230 B.n45 585
R69 B.n229 B.n228 585
R70 B.n227 B.n46 585
R71 B.n226 B.n225 585
R72 B.n224 B.n47 585
R73 B.n223 B.n222 585
R74 B.n221 B.n48 585
R75 B.n220 B.n219 585
R76 B.n218 B.n49 585
R77 B.n217 B.n216 585
R78 B.n215 B.n50 585
R79 B.n214 B.n213 585
R80 B.n212 B.n51 585
R81 B.n211 B.n210 585
R82 B.n209 B.n52 585
R83 B.n208 B.n207 585
R84 B.n206 B.n53 585
R85 B.n205 B.n204 585
R86 B.n203 B.n54 585
R87 B.n202 B.n201 585
R88 B.n200 B.n55 585
R89 B.n199 B.n198 585
R90 B.n197 B.n56 585
R91 B.n196 B.n195 585
R92 B.n194 B.n57 585
R93 B.n193 B.n192 585
R94 B.n191 B.n58 585
R95 B.n190 B.n189 585
R96 B.n188 B.n59 585
R97 B.n187 B.n186 585
R98 B.n124 B.n81 585
R99 B.n126 B.n125 585
R100 B.n127 B.n80 585
R101 B.n129 B.n128 585
R102 B.n130 B.n79 585
R103 B.n132 B.n131 585
R104 B.n133 B.n78 585
R105 B.n135 B.n134 585
R106 B.n136 B.n77 585
R107 B.n138 B.n137 585
R108 B.n139 B.n76 585
R109 B.n141 B.n140 585
R110 B.n142 B.n75 585
R111 B.n144 B.n143 585
R112 B.n145 B.n72 585
R113 B.n148 B.n147 585
R114 B.n149 B.n71 585
R115 B.n151 B.n150 585
R116 B.n152 B.n70 585
R117 B.n154 B.n153 585
R118 B.n155 B.n69 585
R119 B.n157 B.n156 585
R120 B.n158 B.n68 585
R121 B.n163 B.n162 585
R122 B.n164 B.n67 585
R123 B.n166 B.n165 585
R124 B.n167 B.n66 585
R125 B.n169 B.n168 585
R126 B.n170 B.n65 585
R127 B.n172 B.n171 585
R128 B.n173 B.n64 585
R129 B.n175 B.n174 585
R130 B.n176 B.n63 585
R131 B.n178 B.n177 585
R132 B.n179 B.n62 585
R133 B.n181 B.n180 585
R134 B.n182 B.n61 585
R135 B.n184 B.n183 585
R136 B.n185 B.n60 585
R137 B.n123 B.n122 585
R138 B.n121 B.n82 585
R139 B.n120 B.n119 585
R140 B.n118 B.n83 585
R141 B.n117 B.n116 585
R142 B.n115 B.n84 585
R143 B.n114 B.n113 585
R144 B.n112 B.n85 585
R145 B.n111 B.n110 585
R146 B.n109 B.n86 585
R147 B.n108 B.n107 585
R148 B.n106 B.n87 585
R149 B.n105 B.n104 585
R150 B.n103 B.n88 585
R151 B.n102 B.n101 585
R152 B.n100 B.n89 585
R153 B.n99 B.n98 585
R154 B.n97 B.n90 585
R155 B.n96 B.n95 585
R156 B.n94 B.n91 585
R157 B.n93 B.n92 585
R158 B.n2 B.n0 585
R159 B.n345 B.n1 585
R160 B.n344 B.n343 585
R161 B.n342 B.n3 585
R162 B.n341 B.n340 585
R163 B.n339 B.n4 585
R164 B.n338 B.n337 585
R165 B.n336 B.n5 585
R166 B.n335 B.n334 585
R167 B.n333 B.n6 585
R168 B.n332 B.n331 585
R169 B.n330 B.n7 585
R170 B.n329 B.n328 585
R171 B.n327 B.n8 585
R172 B.n326 B.n325 585
R173 B.n324 B.n9 585
R174 B.n323 B.n322 585
R175 B.n321 B.n10 585
R176 B.n320 B.n319 585
R177 B.n318 B.n11 585
R178 B.n317 B.n316 585
R179 B.n315 B.n12 585
R180 B.n314 B.n313 585
R181 B.n347 B.n346 585
R182 B.n124 B.n123 564.573
R183 B.n314 B.n13 564.573
R184 B.n187 B.n60 564.573
R185 B.n254 B.n253 564.573
R186 B.n159 B.t9 241.333
R187 B.n73 B.t0 241.333
R188 B.n22 B.t6 241.333
R189 B.n29 B.t3 241.333
R190 B.n159 B.t11 190.476
R191 B.n29 B.t4 190.476
R192 B.n73 B.t2 190.475
R193 B.n22 B.t7 190.475
R194 B.n123 B.n82 163.367
R195 B.n119 B.n82 163.367
R196 B.n119 B.n118 163.367
R197 B.n118 B.n117 163.367
R198 B.n117 B.n84 163.367
R199 B.n113 B.n84 163.367
R200 B.n113 B.n112 163.367
R201 B.n112 B.n111 163.367
R202 B.n111 B.n86 163.367
R203 B.n107 B.n86 163.367
R204 B.n107 B.n106 163.367
R205 B.n106 B.n105 163.367
R206 B.n105 B.n88 163.367
R207 B.n101 B.n88 163.367
R208 B.n101 B.n100 163.367
R209 B.n100 B.n99 163.367
R210 B.n99 B.n90 163.367
R211 B.n95 B.n90 163.367
R212 B.n95 B.n94 163.367
R213 B.n94 B.n93 163.367
R214 B.n93 B.n2 163.367
R215 B.n346 B.n2 163.367
R216 B.n346 B.n345 163.367
R217 B.n345 B.n344 163.367
R218 B.n344 B.n3 163.367
R219 B.n340 B.n3 163.367
R220 B.n340 B.n339 163.367
R221 B.n339 B.n338 163.367
R222 B.n338 B.n5 163.367
R223 B.n334 B.n5 163.367
R224 B.n334 B.n333 163.367
R225 B.n333 B.n332 163.367
R226 B.n332 B.n7 163.367
R227 B.n328 B.n7 163.367
R228 B.n328 B.n327 163.367
R229 B.n327 B.n326 163.367
R230 B.n326 B.n9 163.367
R231 B.n322 B.n9 163.367
R232 B.n322 B.n321 163.367
R233 B.n321 B.n320 163.367
R234 B.n320 B.n11 163.367
R235 B.n316 B.n11 163.367
R236 B.n316 B.n315 163.367
R237 B.n315 B.n314 163.367
R238 B.n125 B.n124 163.367
R239 B.n125 B.n80 163.367
R240 B.n129 B.n80 163.367
R241 B.n130 B.n129 163.367
R242 B.n131 B.n130 163.367
R243 B.n131 B.n78 163.367
R244 B.n135 B.n78 163.367
R245 B.n136 B.n135 163.367
R246 B.n137 B.n136 163.367
R247 B.n137 B.n76 163.367
R248 B.n141 B.n76 163.367
R249 B.n142 B.n141 163.367
R250 B.n143 B.n142 163.367
R251 B.n143 B.n72 163.367
R252 B.n148 B.n72 163.367
R253 B.n149 B.n148 163.367
R254 B.n150 B.n149 163.367
R255 B.n150 B.n70 163.367
R256 B.n154 B.n70 163.367
R257 B.n155 B.n154 163.367
R258 B.n156 B.n155 163.367
R259 B.n156 B.n68 163.367
R260 B.n163 B.n68 163.367
R261 B.n164 B.n163 163.367
R262 B.n165 B.n164 163.367
R263 B.n165 B.n66 163.367
R264 B.n169 B.n66 163.367
R265 B.n170 B.n169 163.367
R266 B.n171 B.n170 163.367
R267 B.n171 B.n64 163.367
R268 B.n175 B.n64 163.367
R269 B.n176 B.n175 163.367
R270 B.n177 B.n176 163.367
R271 B.n177 B.n62 163.367
R272 B.n181 B.n62 163.367
R273 B.n182 B.n181 163.367
R274 B.n183 B.n182 163.367
R275 B.n183 B.n60 163.367
R276 B.n188 B.n187 163.367
R277 B.n189 B.n188 163.367
R278 B.n189 B.n58 163.367
R279 B.n193 B.n58 163.367
R280 B.n194 B.n193 163.367
R281 B.n195 B.n194 163.367
R282 B.n195 B.n56 163.367
R283 B.n199 B.n56 163.367
R284 B.n200 B.n199 163.367
R285 B.n201 B.n200 163.367
R286 B.n201 B.n54 163.367
R287 B.n205 B.n54 163.367
R288 B.n206 B.n205 163.367
R289 B.n207 B.n206 163.367
R290 B.n207 B.n52 163.367
R291 B.n211 B.n52 163.367
R292 B.n212 B.n211 163.367
R293 B.n213 B.n212 163.367
R294 B.n213 B.n50 163.367
R295 B.n217 B.n50 163.367
R296 B.n218 B.n217 163.367
R297 B.n219 B.n218 163.367
R298 B.n219 B.n48 163.367
R299 B.n223 B.n48 163.367
R300 B.n224 B.n223 163.367
R301 B.n225 B.n224 163.367
R302 B.n225 B.n46 163.367
R303 B.n229 B.n46 163.367
R304 B.n230 B.n229 163.367
R305 B.n231 B.n230 163.367
R306 B.n231 B.n44 163.367
R307 B.n235 B.n44 163.367
R308 B.n236 B.n235 163.367
R309 B.n237 B.n236 163.367
R310 B.n237 B.n42 163.367
R311 B.n241 B.n42 163.367
R312 B.n242 B.n241 163.367
R313 B.n243 B.n242 163.367
R314 B.n243 B.n40 163.367
R315 B.n247 B.n40 163.367
R316 B.n248 B.n247 163.367
R317 B.n249 B.n248 163.367
R318 B.n249 B.n38 163.367
R319 B.n253 B.n38 163.367
R320 B.n310 B.n13 163.367
R321 B.n310 B.n309 163.367
R322 B.n309 B.n308 163.367
R323 B.n308 B.n15 163.367
R324 B.n304 B.n15 163.367
R325 B.n304 B.n303 163.367
R326 B.n303 B.n302 163.367
R327 B.n302 B.n17 163.367
R328 B.n298 B.n17 163.367
R329 B.n298 B.n297 163.367
R330 B.n297 B.n296 163.367
R331 B.n296 B.n19 163.367
R332 B.n292 B.n19 163.367
R333 B.n292 B.n291 163.367
R334 B.n291 B.n290 163.367
R335 B.n290 B.n21 163.367
R336 B.n286 B.n21 163.367
R337 B.n286 B.n285 163.367
R338 B.n285 B.n284 163.367
R339 B.n284 B.n26 163.367
R340 B.n280 B.n26 163.367
R341 B.n280 B.n279 163.367
R342 B.n279 B.n278 163.367
R343 B.n278 B.n28 163.367
R344 B.n273 B.n28 163.367
R345 B.n273 B.n272 163.367
R346 B.n272 B.n271 163.367
R347 B.n271 B.n32 163.367
R348 B.n267 B.n32 163.367
R349 B.n267 B.n266 163.367
R350 B.n266 B.n265 163.367
R351 B.n265 B.n34 163.367
R352 B.n261 B.n34 163.367
R353 B.n261 B.n260 163.367
R354 B.n260 B.n259 163.367
R355 B.n259 B.n36 163.367
R356 B.n255 B.n36 163.367
R357 B.n255 B.n254 163.367
R358 B.n160 B.t10 144.125
R359 B.n30 B.t5 144.125
R360 B.n74 B.t1 144.123
R361 B.n23 B.t8 144.123
R362 B.n161 B.n160 59.5399
R363 B.n146 B.n74 59.5399
R364 B.n24 B.n23 59.5399
R365 B.n276 B.n30 59.5399
R366 B.n160 B.n159 46.352
R367 B.n74 B.n73 46.352
R368 B.n23 B.n22 46.352
R369 B.n30 B.n29 46.352
R370 B.n313 B.n312 36.6834
R371 B.n252 B.n37 36.6834
R372 B.n186 B.n185 36.6834
R373 B.n122 B.n81 36.6834
R374 B B.n347 18.0485
R375 B.n312 B.n311 10.6151
R376 B.n311 B.n14 10.6151
R377 B.n307 B.n14 10.6151
R378 B.n307 B.n306 10.6151
R379 B.n306 B.n305 10.6151
R380 B.n305 B.n16 10.6151
R381 B.n301 B.n16 10.6151
R382 B.n301 B.n300 10.6151
R383 B.n300 B.n299 10.6151
R384 B.n299 B.n18 10.6151
R385 B.n295 B.n18 10.6151
R386 B.n295 B.n294 10.6151
R387 B.n294 B.n293 10.6151
R388 B.n293 B.n20 10.6151
R389 B.n289 B.n288 10.6151
R390 B.n288 B.n287 10.6151
R391 B.n287 B.n25 10.6151
R392 B.n283 B.n25 10.6151
R393 B.n283 B.n282 10.6151
R394 B.n282 B.n281 10.6151
R395 B.n281 B.n27 10.6151
R396 B.n277 B.n27 10.6151
R397 B.n275 B.n274 10.6151
R398 B.n274 B.n31 10.6151
R399 B.n270 B.n31 10.6151
R400 B.n270 B.n269 10.6151
R401 B.n269 B.n268 10.6151
R402 B.n268 B.n33 10.6151
R403 B.n264 B.n33 10.6151
R404 B.n264 B.n263 10.6151
R405 B.n263 B.n262 10.6151
R406 B.n262 B.n35 10.6151
R407 B.n258 B.n35 10.6151
R408 B.n258 B.n257 10.6151
R409 B.n257 B.n256 10.6151
R410 B.n256 B.n37 10.6151
R411 B.n186 B.n59 10.6151
R412 B.n190 B.n59 10.6151
R413 B.n191 B.n190 10.6151
R414 B.n192 B.n191 10.6151
R415 B.n192 B.n57 10.6151
R416 B.n196 B.n57 10.6151
R417 B.n197 B.n196 10.6151
R418 B.n198 B.n197 10.6151
R419 B.n198 B.n55 10.6151
R420 B.n202 B.n55 10.6151
R421 B.n203 B.n202 10.6151
R422 B.n204 B.n203 10.6151
R423 B.n204 B.n53 10.6151
R424 B.n208 B.n53 10.6151
R425 B.n209 B.n208 10.6151
R426 B.n210 B.n209 10.6151
R427 B.n210 B.n51 10.6151
R428 B.n214 B.n51 10.6151
R429 B.n215 B.n214 10.6151
R430 B.n216 B.n215 10.6151
R431 B.n216 B.n49 10.6151
R432 B.n220 B.n49 10.6151
R433 B.n221 B.n220 10.6151
R434 B.n222 B.n221 10.6151
R435 B.n222 B.n47 10.6151
R436 B.n226 B.n47 10.6151
R437 B.n227 B.n226 10.6151
R438 B.n228 B.n227 10.6151
R439 B.n228 B.n45 10.6151
R440 B.n232 B.n45 10.6151
R441 B.n233 B.n232 10.6151
R442 B.n234 B.n233 10.6151
R443 B.n234 B.n43 10.6151
R444 B.n238 B.n43 10.6151
R445 B.n239 B.n238 10.6151
R446 B.n240 B.n239 10.6151
R447 B.n240 B.n41 10.6151
R448 B.n244 B.n41 10.6151
R449 B.n245 B.n244 10.6151
R450 B.n246 B.n245 10.6151
R451 B.n246 B.n39 10.6151
R452 B.n250 B.n39 10.6151
R453 B.n251 B.n250 10.6151
R454 B.n252 B.n251 10.6151
R455 B.n126 B.n81 10.6151
R456 B.n127 B.n126 10.6151
R457 B.n128 B.n127 10.6151
R458 B.n128 B.n79 10.6151
R459 B.n132 B.n79 10.6151
R460 B.n133 B.n132 10.6151
R461 B.n134 B.n133 10.6151
R462 B.n134 B.n77 10.6151
R463 B.n138 B.n77 10.6151
R464 B.n139 B.n138 10.6151
R465 B.n140 B.n139 10.6151
R466 B.n140 B.n75 10.6151
R467 B.n144 B.n75 10.6151
R468 B.n145 B.n144 10.6151
R469 B.n147 B.n71 10.6151
R470 B.n151 B.n71 10.6151
R471 B.n152 B.n151 10.6151
R472 B.n153 B.n152 10.6151
R473 B.n153 B.n69 10.6151
R474 B.n157 B.n69 10.6151
R475 B.n158 B.n157 10.6151
R476 B.n162 B.n158 10.6151
R477 B.n166 B.n67 10.6151
R478 B.n167 B.n166 10.6151
R479 B.n168 B.n167 10.6151
R480 B.n168 B.n65 10.6151
R481 B.n172 B.n65 10.6151
R482 B.n173 B.n172 10.6151
R483 B.n174 B.n173 10.6151
R484 B.n174 B.n63 10.6151
R485 B.n178 B.n63 10.6151
R486 B.n179 B.n178 10.6151
R487 B.n180 B.n179 10.6151
R488 B.n180 B.n61 10.6151
R489 B.n184 B.n61 10.6151
R490 B.n185 B.n184 10.6151
R491 B.n122 B.n121 10.6151
R492 B.n121 B.n120 10.6151
R493 B.n120 B.n83 10.6151
R494 B.n116 B.n83 10.6151
R495 B.n116 B.n115 10.6151
R496 B.n115 B.n114 10.6151
R497 B.n114 B.n85 10.6151
R498 B.n110 B.n85 10.6151
R499 B.n110 B.n109 10.6151
R500 B.n109 B.n108 10.6151
R501 B.n108 B.n87 10.6151
R502 B.n104 B.n87 10.6151
R503 B.n104 B.n103 10.6151
R504 B.n103 B.n102 10.6151
R505 B.n102 B.n89 10.6151
R506 B.n98 B.n89 10.6151
R507 B.n98 B.n97 10.6151
R508 B.n97 B.n96 10.6151
R509 B.n96 B.n91 10.6151
R510 B.n92 B.n91 10.6151
R511 B.n92 B.n0 10.6151
R512 B.n343 B.n1 10.6151
R513 B.n343 B.n342 10.6151
R514 B.n342 B.n341 10.6151
R515 B.n341 B.n4 10.6151
R516 B.n337 B.n4 10.6151
R517 B.n337 B.n336 10.6151
R518 B.n336 B.n335 10.6151
R519 B.n335 B.n6 10.6151
R520 B.n331 B.n6 10.6151
R521 B.n331 B.n330 10.6151
R522 B.n330 B.n329 10.6151
R523 B.n329 B.n8 10.6151
R524 B.n325 B.n8 10.6151
R525 B.n325 B.n324 10.6151
R526 B.n324 B.n323 10.6151
R527 B.n323 B.n10 10.6151
R528 B.n319 B.n10 10.6151
R529 B.n319 B.n318 10.6151
R530 B.n318 B.n317 10.6151
R531 B.n317 B.n12 10.6151
R532 B.n313 B.n12 10.6151
R533 B.n289 B.n24 6.5566
R534 B.n277 B.n276 6.5566
R535 B.n147 B.n146 6.5566
R536 B.n162 B.n161 6.5566
R537 B.n24 B.n20 4.05904
R538 B.n276 B.n275 4.05904
R539 B.n146 B.n145 4.05904
R540 B.n161 B.n67 4.05904
R541 B.n347 B.n0 2.81026
R542 B.n347 B.n1 2.81026
R543 VN VN.t0 129.684
R544 VN VN.t1 93.3806
R545 VDD2.n0 VDD2.t0 182.767
R546 VDD2.n0 VDD2.t1 152.46
R547 VDD2 VDD2.n0 0.573776
C0 VDD2 VTAIL 2.56186f
C1 w_n1926_n1554# B 5.694991f
C2 VN B 0.833939f
C3 VDD2 B 0.949859f
C4 VP w_n1926_n1554# 2.65971f
C5 VTAIL VDD1 2.51295f
C6 VP VN 3.52586f
C7 VDD2 VP 0.315241f
C8 VDD1 B 0.924377f
C9 VDD1 VP 1.0033f
C10 VN w_n1926_n1554# 2.41799f
C11 VDD2 w_n1926_n1554# 1.09857f
C12 VTAIL B 1.42871f
C13 VDD2 VN 0.8426f
C14 VTAIL VP 0.999601f
C15 VDD1 w_n1926_n1554# 1.07968f
C16 VDD1 VN 0.15304f
C17 VDD2 VDD1 0.609067f
C18 VP B 1.23276f
C19 VTAIL w_n1926_n1554# 1.42152f
C20 VTAIL VN 0.985437f
C21 VDD2 VSUBS 0.52864f
C22 VDD1 VSUBS 2.501195f
C23 VTAIL VSUBS 0.378839f
C24 VN VSUBS 5.00419f
C25 VP VSUBS 1.080126f
C26 B VSUBS 2.58901f
C27 w_n1926_n1554# VSUBS 37.9268f
C28 VDD2.t0 VSUBS 0.42024f
C29 VDD2.t1 VSUBS 0.283974f
C30 VDD2.n0 VSUBS 1.80987f
C31 VN.t1 VSUBS 1.06974f
C32 VN.t0 VSUBS 1.58962f
C33 B.n0 VSUBS 0.005126f
C34 B.n1 VSUBS 0.005126f
C35 B.n2 VSUBS 0.008107f
C36 B.n3 VSUBS 0.008107f
C37 B.n4 VSUBS 0.008107f
C38 B.n5 VSUBS 0.008107f
C39 B.n6 VSUBS 0.008107f
C40 B.n7 VSUBS 0.008107f
C41 B.n8 VSUBS 0.008107f
C42 B.n9 VSUBS 0.008107f
C43 B.n10 VSUBS 0.008107f
C44 B.n11 VSUBS 0.008107f
C45 B.n12 VSUBS 0.008107f
C46 B.n13 VSUBS 0.020869f
C47 B.n14 VSUBS 0.008107f
C48 B.n15 VSUBS 0.008107f
C49 B.n16 VSUBS 0.008107f
C50 B.n17 VSUBS 0.008107f
C51 B.n18 VSUBS 0.008107f
C52 B.n19 VSUBS 0.008107f
C53 B.n20 VSUBS 0.005603f
C54 B.n21 VSUBS 0.008107f
C55 B.t8 VSUBS 0.08103f
C56 B.t7 VSUBS 0.095895f
C57 B.t6 VSUBS 0.33783f
C58 B.n22 VSUBS 0.088668f
C59 B.n23 VSUBS 0.072647f
C60 B.n24 VSUBS 0.018783f
C61 B.n25 VSUBS 0.008107f
C62 B.n26 VSUBS 0.008107f
C63 B.n27 VSUBS 0.008107f
C64 B.n28 VSUBS 0.008107f
C65 B.t5 VSUBS 0.08103f
C66 B.t4 VSUBS 0.095895f
C67 B.t3 VSUBS 0.33783f
C68 B.n29 VSUBS 0.088668f
C69 B.n30 VSUBS 0.072647f
C70 B.n31 VSUBS 0.008107f
C71 B.n32 VSUBS 0.008107f
C72 B.n33 VSUBS 0.008107f
C73 B.n34 VSUBS 0.008107f
C74 B.n35 VSUBS 0.008107f
C75 B.n36 VSUBS 0.008107f
C76 B.n37 VSUBS 0.020017f
C77 B.n38 VSUBS 0.008107f
C78 B.n39 VSUBS 0.008107f
C79 B.n40 VSUBS 0.008107f
C80 B.n41 VSUBS 0.008107f
C81 B.n42 VSUBS 0.008107f
C82 B.n43 VSUBS 0.008107f
C83 B.n44 VSUBS 0.008107f
C84 B.n45 VSUBS 0.008107f
C85 B.n46 VSUBS 0.008107f
C86 B.n47 VSUBS 0.008107f
C87 B.n48 VSUBS 0.008107f
C88 B.n49 VSUBS 0.008107f
C89 B.n50 VSUBS 0.008107f
C90 B.n51 VSUBS 0.008107f
C91 B.n52 VSUBS 0.008107f
C92 B.n53 VSUBS 0.008107f
C93 B.n54 VSUBS 0.008107f
C94 B.n55 VSUBS 0.008107f
C95 B.n56 VSUBS 0.008107f
C96 B.n57 VSUBS 0.008107f
C97 B.n58 VSUBS 0.008107f
C98 B.n59 VSUBS 0.008107f
C99 B.n60 VSUBS 0.020869f
C100 B.n61 VSUBS 0.008107f
C101 B.n62 VSUBS 0.008107f
C102 B.n63 VSUBS 0.008107f
C103 B.n64 VSUBS 0.008107f
C104 B.n65 VSUBS 0.008107f
C105 B.n66 VSUBS 0.008107f
C106 B.n67 VSUBS 0.005603f
C107 B.n68 VSUBS 0.008107f
C108 B.n69 VSUBS 0.008107f
C109 B.n70 VSUBS 0.008107f
C110 B.n71 VSUBS 0.008107f
C111 B.n72 VSUBS 0.008107f
C112 B.t1 VSUBS 0.08103f
C113 B.t2 VSUBS 0.095895f
C114 B.t0 VSUBS 0.33783f
C115 B.n73 VSUBS 0.088668f
C116 B.n74 VSUBS 0.072647f
C117 B.n75 VSUBS 0.008107f
C118 B.n76 VSUBS 0.008107f
C119 B.n77 VSUBS 0.008107f
C120 B.n78 VSUBS 0.008107f
C121 B.n79 VSUBS 0.008107f
C122 B.n80 VSUBS 0.008107f
C123 B.n81 VSUBS 0.020869f
C124 B.n82 VSUBS 0.008107f
C125 B.n83 VSUBS 0.008107f
C126 B.n84 VSUBS 0.008107f
C127 B.n85 VSUBS 0.008107f
C128 B.n86 VSUBS 0.008107f
C129 B.n87 VSUBS 0.008107f
C130 B.n88 VSUBS 0.008107f
C131 B.n89 VSUBS 0.008107f
C132 B.n90 VSUBS 0.008107f
C133 B.n91 VSUBS 0.008107f
C134 B.n92 VSUBS 0.008107f
C135 B.n93 VSUBS 0.008107f
C136 B.n94 VSUBS 0.008107f
C137 B.n95 VSUBS 0.008107f
C138 B.n96 VSUBS 0.008107f
C139 B.n97 VSUBS 0.008107f
C140 B.n98 VSUBS 0.008107f
C141 B.n99 VSUBS 0.008107f
C142 B.n100 VSUBS 0.008107f
C143 B.n101 VSUBS 0.008107f
C144 B.n102 VSUBS 0.008107f
C145 B.n103 VSUBS 0.008107f
C146 B.n104 VSUBS 0.008107f
C147 B.n105 VSUBS 0.008107f
C148 B.n106 VSUBS 0.008107f
C149 B.n107 VSUBS 0.008107f
C150 B.n108 VSUBS 0.008107f
C151 B.n109 VSUBS 0.008107f
C152 B.n110 VSUBS 0.008107f
C153 B.n111 VSUBS 0.008107f
C154 B.n112 VSUBS 0.008107f
C155 B.n113 VSUBS 0.008107f
C156 B.n114 VSUBS 0.008107f
C157 B.n115 VSUBS 0.008107f
C158 B.n116 VSUBS 0.008107f
C159 B.n117 VSUBS 0.008107f
C160 B.n118 VSUBS 0.008107f
C161 B.n119 VSUBS 0.008107f
C162 B.n120 VSUBS 0.008107f
C163 B.n121 VSUBS 0.008107f
C164 B.n122 VSUBS 0.020141f
C165 B.n123 VSUBS 0.020141f
C166 B.n124 VSUBS 0.020869f
C167 B.n125 VSUBS 0.008107f
C168 B.n126 VSUBS 0.008107f
C169 B.n127 VSUBS 0.008107f
C170 B.n128 VSUBS 0.008107f
C171 B.n129 VSUBS 0.008107f
C172 B.n130 VSUBS 0.008107f
C173 B.n131 VSUBS 0.008107f
C174 B.n132 VSUBS 0.008107f
C175 B.n133 VSUBS 0.008107f
C176 B.n134 VSUBS 0.008107f
C177 B.n135 VSUBS 0.008107f
C178 B.n136 VSUBS 0.008107f
C179 B.n137 VSUBS 0.008107f
C180 B.n138 VSUBS 0.008107f
C181 B.n139 VSUBS 0.008107f
C182 B.n140 VSUBS 0.008107f
C183 B.n141 VSUBS 0.008107f
C184 B.n142 VSUBS 0.008107f
C185 B.n143 VSUBS 0.008107f
C186 B.n144 VSUBS 0.008107f
C187 B.n145 VSUBS 0.005603f
C188 B.n146 VSUBS 0.018783f
C189 B.n147 VSUBS 0.006557f
C190 B.n148 VSUBS 0.008107f
C191 B.n149 VSUBS 0.008107f
C192 B.n150 VSUBS 0.008107f
C193 B.n151 VSUBS 0.008107f
C194 B.n152 VSUBS 0.008107f
C195 B.n153 VSUBS 0.008107f
C196 B.n154 VSUBS 0.008107f
C197 B.n155 VSUBS 0.008107f
C198 B.n156 VSUBS 0.008107f
C199 B.n157 VSUBS 0.008107f
C200 B.n158 VSUBS 0.008107f
C201 B.t10 VSUBS 0.08103f
C202 B.t11 VSUBS 0.095895f
C203 B.t9 VSUBS 0.33783f
C204 B.n159 VSUBS 0.088668f
C205 B.n160 VSUBS 0.072647f
C206 B.n161 VSUBS 0.018783f
C207 B.n162 VSUBS 0.006557f
C208 B.n163 VSUBS 0.008107f
C209 B.n164 VSUBS 0.008107f
C210 B.n165 VSUBS 0.008107f
C211 B.n166 VSUBS 0.008107f
C212 B.n167 VSUBS 0.008107f
C213 B.n168 VSUBS 0.008107f
C214 B.n169 VSUBS 0.008107f
C215 B.n170 VSUBS 0.008107f
C216 B.n171 VSUBS 0.008107f
C217 B.n172 VSUBS 0.008107f
C218 B.n173 VSUBS 0.008107f
C219 B.n174 VSUBS 0.008107f
C220 B.n175 VSUBS 0.008107f
C221 B.n176 VSUBS 0.008107f
C222 B.n177 VSUBS 0.008107f
C223 B.n178 VSUBS 0.008107f
C224 B.n179 VSUBS 0.008107f
C225 B.n180 VSUBS 0.008107f
C226 B.n181 VSUBS 0.008107f
C227 B.n182 VSUBS 0.008107f
C228 B.n183 VSUBS 0.008107f
C229 B.n184 VSUBS 0.008107f
C230 B.n185 VSUBS 0.020869f
C231 B.n186 VSUBS 0.020141f
C232 B.n187 VSUBS 0.020141f
C233 B.n188 VSUBS 0.008107f
C234 B.n189 VSUBS 0.008107f
C235 B.n190 VSUBS 0.008107f
C236 B.n191 VSUBS 0.008107f
C237 B.n192 VSUBS 0.008107f
C238 B.n193 VSUBS 0.008107f
C239 B.n194 VSUBS 0.008107f
C240 B.n195 VSUBS 0.008107f
C241 B.n196 VSUBS 0.008107f
C242 B.n197 VSUBS 0.008107f
C243 B.n198 VSUBS 0.008107f
C244 B.n199 VSUBS 0.008107f
C245 B.n200 VSUBS 0.008107f
C246 B.n201 VSUBS 0.008107f
C247 B.n202 VSUBS 0.008107f
C248 B.n203 VSUBS 0.008107f
C249 B.n204 VSUBS 0.008107f
C250 B.n205 VSUBS 0.008107f
C251 B.n206 VSUBS 0.008107f
C252 B.n207 VSUBS 0.008107f
C253 B.n208 VSUBS 0.008107f
C254 B.n209 VSUBS 0.008107f
C255 B.n210 VSUBS 0.008107f
C256 B.n211 VSUBS 0.008107f
C257 B.n212 VSUBS 0.008107f
C258 B.n213 VSUBS 0.008107f
C259 B.n214 VSUBS 0.008107f
C260 B.n215 VSUBS 0.008107f
C261 B.n216 VSUBS 0.008107f
C262 B.n217 VSUBS 0.008107f
C263 B.n218 VSUBS 0.008107f
C264 B.n219 VSUBS 0.008107f
C265 B.n220 VSUBS 0.008107f
C266 B.n221 VSUBS 0.008107f
C267 B.n222 VSUBS 0.008107f
C268 B.n223 VSUBS 0.008107f
C269 B.n224 VSUBS 0.008107f
C270 B.n225 VSUBS 0.008107f
C271 B.n226 VSUBS 0.008107f
C272 B.n227 VSUBS 0.008107f
C273 B.n228 VSUBS 0.008107f
C274 B.n229 VSUBS 0.008107f
C275 B.n230 VSUBS 0.008107f
C276 B.n231 VSUBS 0.008107f
C277 B.n232 VSUBS 0.008107f
C278 B.n233 VSUBS 0.008107f
C279 B.n234 VSUBS 0.008107f
C280 B.n235 VSUBS 0.008107f
C281 B.n236 VSUBS 0.008107f
C282 B.n237 VSUBS 0.008107f
C283 B.n238 VSUBS 0.008107f
C284 B.n239 VSUBS 0.008107f
C285 B.n240 VSUBS 0.008107f
C286 B.n241 VSUBS 0.008107f
C287 B.n242 VSUBS 0.008107f
C288 B.n243 VSUBS 0.008107f
C289 B.n244 VSUBS 0.008107f
C290 B.n245 VSUBS 0.008107f
C291 B.n246 VSUBS 0.008107f
C292 B.n247 VSUBS 0.008107f
C293 B.n248 VSUBS 0.008107f
C294 B.n249 VSUBS 0.008107f
C295 B.n250 VSUBS 0.008107f
C296 B.n251 VSUBS 0.008107f
C297 B.n252 VSUBS 0.020994f
C298 B.n253 VSUBS 0.020141f
C299 B.n254 VSUBS 0.020869f
C300 B.n255 VSUBS 0.008107f
C301 B.n256 VSUBS 0.008107f
C302 B.n257 VSUBS 0.008107f
C303 B.n258 VSUBS 0.008107f
C304 B.n259 VSUBS 0.008107f
C305 B.n260 VSUBS 0.008107f
C306 B.n261 VSUBS 0.008107f
C307 B.n262 VSUBS 0.008107f
C308 B.n263 VSUBS 0.008107f
C309 B.n264 VSUBS 0.008107f
C310 B.n265 VSUBS 0.008107f
C311 B.n266 VSUBS 0.008107f
C312 B.n267 VSUBS 0.008107f
C313 B.n268 VSUBS 0.008107f
C314 B.n269 VSUBS 0.008107f
C315 B.n270 VSUBS 0.008107f
C316 B.n271 VSUBS 0.008107f
C317 B.n272 VSUBS 0.008107f
C318 B.n273 VSUBS 0.008107f
C319 B.n274 VSUBS 0.008107f
C320 B.n275 VSUBS 0.005603f
C321 B.n276 VSUBS 0.018783f
C322 B.n277 VSUBS 0.006557f
C323 B.n278 VSUBS 0.008107f
C324 B.n279 VSUBS 0.008107f
C325 B.n280 VSUBS 0.008107f
C326 B.n281 VSUBS 0.008107f
C327 B.n282 VSUBS 0.008107f
C328 B.n283 VSUBS 0.008107f
C329 B.n284 VSUBS 0.008107f
C330 B.n285 VSUBS 0.008107f
C331 B.n286 VSUBS 0.008107f
C332 B.n287 VSUBS 0.008107f
C333 B.n288 VSUBS 0.008107f
C334 B.n289 VSUBS 0.006557f
C335 B.n290 VSUBS 0.008107f
C336 B.n291 VSUBS 0.008107f
C337 B.n292 VSUBS 0.008107f
C338 B.n293 VSUBS 0.008107f
C339 B.n294 VSUBS 0.008107f
C340 B.n295 VSUBS 0.008107f
C341 B.n296 VSUBS 0.008107f
C342 B.n297 VSUBS 0.008107f
C343 B.n298 VSUBS 0.008107f
C344 B.n299 VSUBS 0.008107f
C345 B.n300 VSUBS 0.008107f
C346 B.n301 VSUBS 0.008107f
C347 B.n302 VSUBS 0.008107f
C348 B.n303 VSUBS 0.008107f
C349 B.n304 VSUBS 0.008107f
C350 B.n305 VSUBS 0.008107f
C351 B.n306 VSUBS 0.008107f
C352 B.n307 VSUBS 0.008107f
C353 B.n308 VSUBS 0.008107f
C354 B.n309 VSUBS 0.008107f
C355 B.n310 VSUBS 0.008107f
C356 B.n311 VSUBS 0.008107f
C357 B.n312 VSUBS 0.020869f
C358 B.n313 VSUBS 0.020141f
C359 B.n314 VSUBS 0.020141f
C360 B.n315 VSUBS 0.008107f
C361 B.n316 VSUBS 0.008107f
C362 B.n317 VSUBS 0.008107f
C363 B.n318 VSUBS 0.008107f
C364 B.n319 VSUBS 0.008107f
C365 B.n320 VSUBS 0.008107f
C366 B.n321 VSUBS 0.008107f
C367 B.n322 VSUBS 0.008107f
C368 B.n323 VSUBS 0.008107f
C369 B.n324 VSUBS 0.008107f
C370 B.n325 VSUBS 0.008107f
C371 B.n326 VSUBS 0.008107f
C372 B.n327 VSUBS 0.008107f
C373 B.n328 VSUBS 0.008107f
C374 B.n329 VSUBS 0.008107f
C375 B.n330 VSUBS 0.008107f
C376 B.n331 VSUBS 0.008107f
C377 B.n332 VSUBS 0.008107f
C378 B.n333 VSUBS 0.008107f
C379 B.n334 VSUBS 0.008107f
C380 B.n335 VSUBS 0.008107f
C381 B.n336 VSUBS 0.008107f
C382 B.n337 VSUBS 0.008107f
C383 B.n338 VSUBS 0.008107f
C384 B.n339 VSUBS 0.008107f
C385 B.n340 VSUBS 0.008107f
C386 B.n341 VSUBS 0.008107f
C387 B.n342 VSUBS 0.008107f
C388 B.n343 VSUBS 0.008107f
C389 B.n344 VSUBS 0.008107f
C390 B.n345 VSUBS 0.008107f
C391 B.n346 VSUBS 0.008107f
C392 B.n347 VSUBS 0.018357f
C393 VDD1.t0 VSUBS 0.267713f
C394 VDD1.t1 VSUBS 0.406236f
C395 VTAIL.t3 VSUBS 0.299373f
C396 VTAIL.n0 VSUBS 1.01129f
C397 VTAIL.t0 VSUBS 0.299374f
C398 VTAIL.n1 VSUBS 1.03971f
C399 VTAIL.t2 VSUBS 0.299373f
C400 VTAIL.n2 VSUBS 0.911545f
C401 VTAIL.t1 VSUBS 0.299373f
C402 VTAIL.n3 VSUBS 0.846659f
C403 VP.t1 VSUBS 1.68038f
C404 VP.t0 VSUBS 1.13583f
C405 VP.n0 VSUBS 3.29791f
.ends

