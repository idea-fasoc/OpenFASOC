* NGSPICE file created from diff_pair_sample_0541.ext - technology: sky130A

.subckt diff_pair_sample_0541 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=0 ps=0 w=17.45 l=1.69
X1 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=0 ps=0 w=17.45 l=1.69
X2 VTAIL.t15 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X3 VTAIL.t2 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X4 VTAIL.t14 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=2.87925 ps=17.78 w=17.45 l=1.69
X5 VTAIL.t6 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=2.87925 ps=17.78 w=17.45 l=1.69
X6 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=0 ps=0 w=17.45 l=1.69
X7 VTAIL.t7 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X8 VTAIL.t13 VN.t2 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X9 VDD1.t4 VP.t3 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X10 VDD2.t1 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=6.8055 ps=35.68 w=17.45 l=1.69
X11 VDD2.t3 VN.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X12 VDD2.t0 VN.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=6.8055 ps=35.68 w=17.45 l=1.69
X13 VDD1.t3 VP.t4 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=6.8055 ps=35.68 w=17.45 l=1.69
X14 VTAIL.t1 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=2.87925 ps=17.78 w=17.45 l=1.69
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=0 ps=0 w=17.45 l=1.69
X16 VTAIL.t9 VN.t6 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=6.8055 pd=35.68 as=2.87925 ps=17.78 w=17.45 l=1.69
X17 VDD1.t1 VP.t6 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
X18 VDD1.t0 VP.t7 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=6.8055 ps=35.68 w=17.45 l=1.69
X19 VDD2.t4 VN.t7 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.87925 pd=17.78 as=2.87925 ps=17.78 w=17.45 l=1.69
R0 B.n694 B.n693 585
R1 B.n694 B.n71 585
R2 B.n697 B.n696 585
R3 B.n698 B.n138 585
R4 B.n700 B.n699 585
R5 B.n702 B.n137 585
R6 B.n705 B.n704 585
R7 B.n706 B.n136 585
R8 B.n708 B.n707 585
R9 B.n710 B.n135 585
R10 B.n713 B.n712 585
R11 B.n714 B.n134 585
R12 B.n716 B.n715 585
R13 B.n718 B.n133 585
R14 B.n721 B.n720 585
R15 B.n722 B.n132 585
R16 B.n724 B.n723 585
R17 B.n726 B.n131 585
R18 B.n729 B.n728 585
R19 B.n730 B.n130 585
R20 B.n732 B.n731 585
R21 B.n734 B.n129 585
R22 B.n737 B.n736 585
R23 B.n738 B.n128 585
R24 B.n740 B.n739 585
R25 B.n742 B.n127 585
R26 B.n745 B.n744 585
R27 B.n746 B.n126 585
R28 B.n748 B.n747 585
R29 B.n750 B.n125 585
R30 B.n753 B.n752 585
R31 B.n754 B.n124 585
R32 B.n756 B.n755 585
R33 B.n758 B.n123 585
R34 B.n761 B.n760 585
R35 B.n762 B.n122 585
R36 B.n764 B.n763 585
R37 B.n766 B.n121 585
R38 B.n769 B.n768 585
R39 B.n770 B.n120 585
R40 B.n772 B.n771 585
R41 B.n774 B.n119 585
R42 B.n777 B.n776 585
R43 B.n778 B.n118 585
R44 B.n780 B.n779 585
R45 B.n782 B.n117 585
R46 B.n785 B.n784 585
R47 B.n786 B.n116 585
R48 B.n788 B.n787 585
R49 B.n790 B.n115 585
R50 B.n793 B.n792 585
R51 B.n794 B.n114 585
R52 B.n796 B.n795 585
R53 B.n798 B.n113 585
R54 B.n801 B.n800 585
R55 B.n802 B.n112 585
R56 B.n804 B.n803 585
R57 B.n806 B.n111 585
R58 B.n809 B.n808 585
R59 B.n811 B.n108 585
R60 B.n813 B.n812 585
R61 B.n815 B.n107 585
R62 B.n818 B.n817 585
R63 B.n819 B.n106 585
R64 B.n821 B.n820 585
R65 B.n823 B.n105 585
R66 B.n825 B.n824 585
R67 B.n827 B.n826 585
R68 B.n830 B.n829 585
R69 B.n831 B.n100 585
R70 B.n833 B.n832 585
R71 B.n835 B.n99 585
R72 B.n838 B.n837 585
R73 B.n839 B.n98 585
R74 B.n841 B.n840 585
R75 B.n843 B.n97 585
R76 B.n846 B.n845 585
R77 B.n847 B.n96 585
R78 B.n849 B.n848 585
R79 B.n851 B.n95 585
R80 B.n854 B.n853 585
R81 B.n855 B.n94 585
R82 B.n857 B.n856 585
R83 B.n859 B.n93 585
R84 B.n862 B.n861 585
R85 B.n863 B.n92 585
R86 B.n865 B.n864 585
R87 B.n867 B.n91 585
R88 B.n870 B.n869 585
R89 B.n871 B.n90 585
R90 B.n873 B.n872 585
R91 B.n875 B.n89 585
R92 B.n878 B.n877 585
R93 B.n879 B.n88 585
R94 B.n881 B.n880 585
R95 B.n883 B.n87 585
R96 B.n886 B.n885 585
R97 B.n887 B.n86 585
R98 B.n889 B.n888 585
R99 B.n891 B.n85 585
R100 B.n894 B.n893 585
R101 B.n895 B.n84 585
R102 B.n897 B.n896 585
R103 B.n899 B.n83 585
R104 B.n902 B.n901 585
R105 B.n903 B.n82 585
R106 B.n905 B.n904 585
R107 B.n907 B.n81 585
R108 B.n910 B.n909 585
R109 B.n911 B.n80 585
R110 B.n913 B.n912 585
R111 B.n915 B.n79 585
R112 B.n918 B.n917 585
R113 B.n919 B.n78 585
R114 B.n921 B.n920 585
R115 B.n923 B.n77 585
R116 B.n926 B.n925 585
R117 B.n927 B.n76 585
R118 B.n929 B.n928 585
R119 B.n931 B.n75 585
R120 B.n934 B.n933 585
R121 B.n935 B.n74 585
R122 B.n937 B.n936 585
R123 B.n939 B.n73 585
R124 B.n942 B.n941 585
R125 B.n943 B.n72 585
R126 B.n692 B.n70 585
R127 B.n946 B.n70 585
R128 B.n691 B.n69 585
R129 B.n947 B.n69 585
R130 B.n690 B.n68 585
R131 B.n948 B.n68 585
R132 B.n689 B.n688 585
R133 B.n688 B.n64 585
R134 B.n687 B.n63 585
R135 B.n954 B.n63 585
R136 B.n686 B.n62 585
R137 B.n955 B.n62 585
R138 B.n685 B.n61 585
R139 B.n956 B.n61 585
R140 B.n684 B.n683 585
R141 B.n683 B.n57 585
R142 B.n682 B.n56 585
R143 B.n962 B.n56 585
R144 B.n681 B.n55 585
R145 B.n963 B.n55 585
R146 B.n680 B.n54 585
R147 B.n964 B.n54 585
R148 B.n679 B.n678 585
R149 B.n678 B.n50 585
R150 B.n677 B.n49 585
R151 B.n970 B.n49 585
R152 B.n676 B.n48 585
R153 B.n971 B.n48 585
R154 B.n675 B.n47 585
R155 B.n972 B.n47 585
R156 B.n674 B.n673 585
R157 B.n673 B.n46 585
R158 B.n672 B.n42 585
R159 B.n978 B.n42 585
R160 B.n671 B.n41 585
R161 B.n979 B.n41 585
R162 B.n670 B.n40 585
R163 B.n980 B.n40 585
R164 B.n669 B.n668 585
R165 B.n668 B.n36 585
R166 B.n667 B.n35 585
R167 B.n986 B.n35 585
R168 B.n666 B.n34 585
R169 B.n987 B.n34 585
R170 B.n665 B.n33 585
R171 B.n988 B.n33 585
R172 B.n664 B.n663 585
R173 B.n663 B.n29 585
R174 B.n662 B.n28 585
R175 B.n994 B.n28 585
R176 B.n661 B.n27 585
R177 B.n995 B.n27 585
R178 B.n660 B.n26 585
R179 B.n996 B.n26 585
R180 B.n659 B.n658 585
R181 B.n658 B.n25 585
R182 B.n657 B.n21 585
R183 B.n1002 B.n21 585
R184 B.n656 B.n20 585
R185 B.n1003 B.n20 585
R186 B.n655 B.n19 585
R187 B.n1004 B.n19 585
R188 B.n654 B.n653 585
R189 B.n653 B.n15 585
R190 B.n652 B.n14 585
R191 B.n1010 B.n14 585
R192 B.n651 B.n13 585
R193 B.n1011 B.n13 585
R194 B.n650 B.n12 585
R195 B.n1012 B.n12 585
R196 B.n649 B.n648 585
R197 B.n648 B.n8 585
R198 B.n647 B.n7 585
R199 B.n1018 B.n7 585
R200 B.n646 B.n6 585
R201 B.n1019 B.n6 585
R202 B.n645 B.n5 585
R203 B.n1020 B.n5 585
R204 B.n644 B.n643 585
R205 B.n643 B.n4 585
R206 B.n642 B.n139 585
R207 B.n642 B.n641 585
R208 B.n632 B.n140 585
R209 B.n141 B.n140 585
R210 B.n634 B.n633 585
R211 B.n635 B.n634 585
R212 B.n631 B.n145 585
R213 B.n149 B.n145 585
R214 B.n630 B.n629 585
R215 B.n629 B.n628 585
R216 B.n147 B.n146 585
R217 B.n148 B.n147 585
R218 B.n621 B.n620 585
R219 B.n622 B.n621 585
R220 B.n619 B.n154 585
R221 B.n154 B.n153 585
R222 B.n618 B.n617 585
R223 B.n617 B.n616 585
R224 B.n156 B.n155 585
R225 B.n609 B.n156 585
R226 B.n608 B.n607 585
R227 B.n610 B.n608 585
R228 B.n606 B.n161 585
R229 B.n161 B.n160 585
R230 B.n605 B.n604 585
R231 B.n604 B.n603 585
R232 B.n163 B.n162 585
R233 B.n164 B.n163 585
R234 B.n596 B.n595 585
R235 B.n597 B.n596 585
R236 B.n594 B.n168 585
R237 B.n172 B.n168 585
R238 B.n593 B.n592 585
R239 B.n592 B.n591 585
R240 B.n170 B.n169 585
R241 B.n171 B.n170 585
R242 B.n584 B.n583 585
R243 B.n585 B.n584 585
R244 B.n582 B.n177 585
R245 B.n177 B.n176 585
R246 B.n581 B.n580 585
R247 B.n580 B.n579 585
R248 B.n179 B.n178 585
R249 B.n572 B.n179 585
R250 B.n571 B.n570 585
R251 B.n573 B.n571 585
R252 B.n569 B.n184 585
R253 B.n184 B.n183 585
R254 B.n568 B.n567 585
R255 B.n567 B.n566 585
R256 B.n186 B.n185 585
R257 B.n187 B.n186 585
R258 B.n559 B.n558 585
R259 B.n560 B.n559 585
R260 B.n557 B.n192 585
R261 B.n192 B.n191 585
R262 B.n556 B.n555 585
R263 B.n555 B.n554 585
R264 B.n194 B.n193 585
R265 B.n195 B.n194 585
R266 B.n547 B.n546 585
R267 B.n548 B.n547 585
R268 B.n545 B.n200 585
R269 B.n200 B.n199 585
R270 B.n544 B.n543 585
R271 B.n543 B.n542 585
R272 B.n202 B.n201 585
R273 B.n203 B.n202 585
R274 B.n535 B.n534 585
R275 B.n536 B.n535 585
R276 B.n533 B.n208 585
R277 B.n208 B.n207 585
R278 B.n532 B.n531 585
R279 B.n531 B.n530 585
R280 B.n527 B.n212 585
R281 B.n526 B.n525 585
R282 B.n523 B.n213 585
R283 B.n523 B.n211 585
R284 B.n522 B.n521 585
R285 B.n520 B.n519 585
R286 B.n518 B.n215 585
R287 B.n516 B.n515 585
R288 B.n514 B.n216 585
R289 B.n513 B.n512 585
R290 B.n510 B.n217 585
R291 B.n508 B.n507 585
R292 B.n506 B.n218 585
R293 B.n505 B.n504 585
R294 B.n502 B.n219 585
R295 B.n500 B.n499 585
R296 B.n498 B.n220 585
R297 B.n497 B.n496 585
R298 B.n494 B.n221 585
R299 B.n492 B.n491 585
R300 B.n490 B.n222 585
R301 B.n489 B.n488 585
R302 B.n486 B.n223 585
R303 B.n484 B.n483 585
R304 B.n482 B.n224 585
R305 B.n481 B.n480 585
R306 B.n478 B.n225 585
R307 B.n476 B.n475 585
R308 B.n474 B.n226 585
R309 B.n473 B.n472 585
R310 B.n470 B.n227 585
R311 B.n468 B.n467 585
R312 B.n466 B.n228 585
R313 B.n465 B.n464 585
R314 B.n462 B.n229 585
R315 B.n460 B.n459 585
R316 B.n458 B.n230 585
R317 B.n457 B.n456 585
R318 B.n454 B.n231 585
R319 B.n452 B.n451 585
R320 B.n450 B.n232 585
R321 B.n449 B.n448 585
R322 B.n446 B.n233 585
R323 B.n444 B.n443 585
R324 B.n442 B.n234 585
R325 B.n441 B.n440 585
R326 B.n438 B.n235 585
R327 B.n436 B.n435 585
R328 B.n434 B.n236 585
R329 B.n433 B.n432 585
R330 B.n430 B.n237 585
R331 B.n428 B.n427 585
R332 B.n426 B.n238 585
R333 B.n425 B.n424 585
R334 B.n422 B.n239 585
R335 B.n420 B.n419 585
R336 B.n418 B.n240 585
R337 B.n417 B.n416 585
R338 B.n414 B.n241 585
R339 B.n412 B.n411 585
R340 B.n410 B.n242 585
R341 B.n409 B.n408 585
R342 B.n406 B.n246 585
R343 B.n404 B.n403 585
R344 B.n402 B.n247 585
R345 B.n401 B.n400 585
R346 B.n398 B.n248 585
R347 B.n396 B.n395 585
R348 B.n393 B.n249 585
R349 B.n392 B.n391 585
R350 B.n389 B.n252 585
R351 B.n387 B.n386 585
R352 B.n385 B.n253 585
R353 B.n384 B.n383 585
R354 B.n381 B.n254 585
R355 B.n379 B.n378 585
R356 B.n377 B.n255 585
R357 B.n376 B.n375 585
R358 B.n373 B.n256 585
R359 B.n371 B.n370 585
R360 B.n369 B.n257 585
R361 B.n368 B.n367 585
R362 B.n365 B.n258 585
R363 B.n363 B.n362 585
R364 B.n361 B.n259 585
R365 B.n360 B.n359 585
R366 B.n357 B.n260 585
R367 B.n355 B.n354 585
R368 B.n353 B.n261 585
R369 B.n352 B.n351 585
R370 B.n349 B.n262 585
R371 B.n347 B.n346 585
R372 B.n345 B.n263 585
R373 B.n344 B.n343 585
R374 B.n341 B.n264 585
R375 B.n339 B.n338 585
R376 B.n337 B.n265 585
R377 B.n336 B.n335 585
R378 B.n333 B.n266 585
R379 B.n331 B.n330 585
R380 B.n329 B.n267 585
R381 B.n328 B.n327 585
R382 B.n325 B.n268 585
R383 B.n323 B.n322 585
R384 B.n321 B.n269 585
R385 B.n320 B.n319 585
R386 B.n317 B.n270 585
R387 B.n315 B.n314 585
R388 B.n313 B.n271 585
R389 B.n312 B.n311 585
R390 B.n309 B.n272 585
R391 B.n307 B.n306 585
R392 B.n305 B.n273 585
R393 B.n304 B.n303 585
R394 B.n301 B.n274 585
R395 B.n299 B.n298 585
R396 B.n297 B.n275 585
R397 B.n296 B.n295 585
R398 B.n293 B.n276 585
R399 B.n291 B.n290 585
R400 B.n289 B.n277 585
R401 B.n288 B.n287 585
R402 B.n285 B.n278 585
R403 B.n283 B.n282 585
R404 B.n281 B.n280 585
R405 B.n210 B.n209 585
R406 B.n529 B.n528 585
R407 B.n530 B.n529 585
R408 B.n206 B.n205 585
R409 B.n207 B.n206 585
R410 B.n538 B.n537 585
R411 B.n537 B.n536 585
R412 B.n539 B.n204 585
R413 B.n204 B.n203 585
R414 B.n541 B.n540 585
R415 B.n542 B.n541 585
R416 B.n198 B.n197 585
R417 B.n199 B.n198 585
R418 B.n550 B.n549 585
R419 B.n549 B.n548 585
R420 B.n551 B.n196 585
R421 B.n196 B.n195 585
R422 B.n553 B.n552 585
R423 B.n554 B.n553 585
R424 B.n190 B.n189 585
R425 B.n191 B.n190 585
R426 B.n562 B.n561 585
R427 B.n561 B.n560 585
R428 B.n563 B.n188 585
R429 B.n188 B.n187 585
R430 B.n565 B.n564 585
R431 B.n566 B.n565 585
R432 B.n182 B.n181 585
R433 B.n183 B.n182 585
R434 B.n575 B.n574 585
R435 B.n574 B.n573 585
R436 B.n576 B.n180 585
R437 B.n572 B.n180 585
R438 B.n578 B.n577 585
R439 B.n579 B.n578 585
R440 B.n175 B.n174 585
R441 B.n176 B.n175 585
R442 B.n587 B.n586 585
R443 B.n586 B.n585 585
R444 B.n588 B.n173 585
R445 B.n173 B.n171 585
R446 B.n590 B.n589 585
R447 B.n591 B.n590 585
R448 B.n167 B.n166 585
R449 B.n172 B.n167 585
R450 B.n599 B.n598 585
R451 B.n598 B.n597 585
R452 B.n600 B.n165 585
R453 B.n165 B.n164 585
R454 B.n602 B.n601 585
R455 B.n603 B.n602 585
R456 B.n159 B.n158 585
R457 B.n160 B.n159 585
R458 B.n612 B.n611 585
R459 B.n611 B.n610 585
R460 B.n613 B.n157 585
R461 B.n609 B.n157 585
R462 B.n615 B.n614 585
R463 B.n616 B.n615 585
R464 B.n152 B.n151 585
R465 B.n153 B.n152 585
R466 B.n624 B.n623 585
R467 B.n623 B.n622 585
R468 B.n625 B.n150 585
R469 B.n150 B.n148 585
R470 B.n627 B.n626 585
R471 B.n628 B.n627 585
R472 B.n144 B.n143 585
R473 B.n149 B.n144 585
R474 B.n637 B.n636 585
R475 B.n636 B.n635 585
R476 B.n638 B.n142 585
R477 B.n142 B.n141 585
R478 B.n640 B.n639 585
R479 B.n641 B.n640 585
R480 B.n2 B.n0 585
R481 B.n4 B.n2 585
R482 B.n3 B.n1 585
R483 B.n1019 B.n3 585
R484 B.n1017 B.n1016 585
R485 B.n1018 B.n1017 585
R486 B.n1015 B.n9 585
R487 B.n9 B.n8 585
R488 B.n1014 B.n1013 585
R489 B.n1013 B.n1012 585
R490 B.n11 B.n10 585
R491 B.n1011 B.n11 585
R492 B.n1009 B.n1008 585
R493 B.n1010 B.n1009 585
R494 B.n1007 B.n16 585
R495 B.n16 B.n15 585
R496 B.n1006 B.n1005 585
R497 B.n1005 B.n1004 585
R498 B.n18 B.n17 585
R499 B.n1003 B.n18 585
R500 B.n1001 B.n1000 585
R501 B.n1002 B.n1001 585
R502 B.n999 B.n22 585
R503 B.n25 B.n22 585
R504 B.n998 B.n997 585
R505 B.n997 B.n996 585
R506 B.n24 B.n23 585
R507 B.n995 B.n24 585
R508 B.n993 B.n992 585
R509 B.n994 B.n993 585
R510 B.n991 B.n30 585
R511 B.n30 B.n29 585
R512 B.n990 B.n989 585
R513 B.n989 B.n988 585
R514 B.n32 B.n31 585
R515 B.n987 B.n32 585
R516 B.n985 B.n984 585
R517 B.n986 B.n985 585
R518 B.n983 B.n37 585
R519 B.n37 B.n36 585
R520 B.n982 B.n981 585
R521 B.n981 B.n980 585
R522 B.n39 B.n38 585
R523 B.n979 B.n39 585
R524 B.n977 B.n976 585
R525 B.n978 B.n977 585
R526 B.n975 B.n43 585
R527 B.n46 B.n43 585
R528 B.n974 B.n973 585
R529 B.n973 B.n972 585
R530 B.n45 B.n44 585
R531 B.n971 B.n45 585
R532 B.n969 B.n968 585
R533 B.n970 B.n969 585
R534 B.n967 B.n51 585
R535 B.n51 B.n50 585
R536 B.n966 B.n965 585
R537 B.n965 B.n964 585
R538 B.n53 B.n52 585
R539 B.n963 B.n53 585
R540 B.n961 B.n960 585
R541 B.n962 B.n961 585
R542 B.n959 B.n58 585
R543 B.n58 B.n57 585
R544 B.n958 B.n957 585
R545 B.n957 B.n956 585
R546 B.n60 B.n59 585
R547 B.n955 B.n60 585
R548 B.n953 B.n952 585
R549 B.n954 B.n953 585
R550 B.n951 B.n65 585
R551 B.n65 B.n64 585
R552 B.n950 B.n949 585
R553 B.n949 B.n948 585
R554 B.n67 B.n66 585
R555 B.n947 B.n67 585
R556 B.n945 B.n944 585
R557 B.n946 B.n945 585
R558 B.n1022 B.n1021 585
R559 B.n1021 B.n1020 585
R560 B.n529 B.n212 458.866
R561 B.n945 B.n72 458.866
R562 B.n531 B.n210 458.866
R563 B.n694 B.n70 458.866
R564 B.n250 B.t19 454.928
R565 B.n243 B.t12 454.928
R566 B.n101 B.t8 454.928
R567 B.n109 B.t16 454.928
R568 B.n250 B.t21 415.077
R569 B.n109 B.t17 415.077
R570 B.n243 B.t15 415.077
R571 B.n101 B.t10 415.077
R572 B.n251 B.t20 375.901
R573 B.n110 B.t18 375.901
R574 B.n244 B.t14 375.901
R575 B.n102 B.t11 375.901
R576 B.n695 B.n71 256.663
R577 B.n701 B.n71 256.663
R578 B.n703 B.n71 256.663
R579 B.n709 B.n71 256.663
R580 B.n711 B.n71 256.663
R581 B.n717 B.n71 256.663
R582 B.n719 B.n71 256.663
R583 B.n725 B.n71 256.663
R584 B.n727 B.n71 256.663
R585 B.n733 B.n71 256.663
R586 B.n735 B.n71 256.663
R587 B.n741 B.n71 256.663
R588 B.n743 B.n71 256.663
R589 B.n749 B.n71 256.663
R590 B.n751 B.n71 256.663
R591 B.n757 B.n71 256.663
R592 B.n759 B.n71 256.663
R593 B.n765 B.n71 256.663
R594 B.n767 B.n71 256.663
R595 B.n773 B.n71 256.663
R596 B.n775 B.n71 256.663
R597 B.n781 B.n71 256.663
R598 B.n783 B.n71 256.663
R599 B.n789 B.n71 256.663
R600 B.n791 B.n71 256.663
R601 B.n797 B.n71 256.663
R602 B.n799 B.n71 256.663
R603 B.n805 B.n71 256.663
R604 B.n807 B.n71 256.663
R605 B.n814 B.n71 256.663
R606 B.n816 B.n71 256.663
R607 B.n822 B.n71 256.663
R608 B.n104 B.n71 256.663
R609 B.n828 B.n71 256.663
R610 B.n834 B.n71 256.663
R611 B.n836 B.n71 256.663
R612 B.n842 B.n71 256.663
R613 B.n844 B.n71 256.663
R614 B.n850 B.n71 256.663
R615 B.n852 B.n71 256.663
R616 B.n858 B.n71 256.663
R617 B.n860 B.n71 256.663
R618 B.n866 B.n71 256.663
R619 B.n868 B.n71 256.663
R620 B.n874 B.n71 256.663
R621 B.n876 B.n71 256.663
R622 B.n882 B.n71 256.663
R623 B.n884 B.n71 256.663
R624 B.n890 B.n71 256.663
R625 B.n892 B.n71 256.663
R626 B.n898 B.n71 256.663
R627 B.n900 B.n71 256.663
R628 B.n906 B.n71 256.663
R629 B.n908 B.n71 256.663
R630 B.n914 B.n71 256.663
R631 B.n916 B.n71 256.663
R632 B.n922 B.n71 256.663
R633 B.n924 B.n71 256.663
R634 B.n930 B.n71 256.663
R635 B.n932 B.n71 256.663
R636 B.n938 B.n71 256.663
R637 B.n940 B.n71 256.663
R638 B.n524 B.n211 256.663
R639 B.n214 B.n211 256.663
R640 B.n517 B.n211 256.663
R641 B.n511 B.n211 256.663
R642 B.n509 B.n211 256.663
R643 B.n503 B.n211 256.663
R644 B.n501 B.n211 256.663
R645 B.n495 B.n211 256.663
R646 B.n493 B.n211 256.663
R647 B.n487 B.n211 256.663
R648 B.n485 B.n211 256.663
R649 B.n479 B.n211 256.663
R650 B.n477 B.n211 256.663
R651 B.n471 B.n211 256.663
R652 B.n469 B.n211 256.663
R653 B.n463 B.n211 256.663
R654 B.n461 B.n211 256.663
R655 B.n455 B.n211 256.663
R656 B.n453 B.n211 256.663
R657 B.n447 B.n211 256.663
R658 B.n445 B.n211 256.663
R659 B.n439 B.n211 256.663
R660 B.n437 B.n211 256.663
R661 B.n431 B.n211 256.663
R662 B.n429 B.n211 256.663
R663 B.n423 B.n211 256.663
R664 B.n421 B.n211 256.663
R665 B.n415 B.n211 256.663
R666 B.n413 B.n211 256.663
R667 B.n407 B.n211 256.663
R668 B.n405 B.n211 256.663
R669 B.n399 B.n211 256.663
R670 B.n397 B.n211 256.663
R671 B.n390 B.n211 256.663
R672 B.n388 B.n211 256.663
R673 B.n382 B.n211 256.663
R674 B.n380 B.n211 256.663
R675 B.n374 B.n211 256.663
R676 B.n372 B.n211 256.663
R677 B.n366 B.n211 256.663
R678 B.n364 B.n211 256.663
R679 B.n358 B.n211 256.663
R680 B.n356 B.n211 256.663
R681 B.n350 B.n211 256.663
R682 B.n348 B.n211 256.663
R683 B.n342 B.n211 256.663
R684 B.n340 B.n211 256.663
R685 B.n334 B.n211 256.663
R686 B.n332 B.n211 256.663
R687 B.n326 B.n211 256.663
R688 B.n324 B.n211 256.663
R689 B.n318 B.n211 256.663
R690 B.n316 B.n211 256.663
R691 B.n310 B.n211 256.663
R692 B.n308 B.n211 256.663
R693 B.n302 B.n211 256.663
R694 B.n300 B.n211 256.663
R695 B.n294 B.n211 256.663
R696 B.n292 B.n211 256.663
R697 B.n286 B.n211 256.663
R698 B.n284 B.n211 256.663
R699 B.n279 B.n211 256.663
R700 B.n529 B.n206 163.367
R701 B.n537 B.n206 163.367
R702 B.n537 B.n204 163.367
R703 B.n541 B.n204 163.367
R704 B.n541 B.n198 163.367
R705 B.n549 B.n198 163.367
R706 B.n549 B.n196 163.367
R707 B.n553 B.n196 163.367
R708 B.n553 B.n190 163.367
R709 B.n561 B.n190 163.367
R710 B.n561 B.n188 163.367
R711 B.n565 B.n188 163.367
R712 B.n565 B.n182 163.367
R713 B.n574 B.n182 163.367
R714 B.n574 B.n180 163.367
R715 B.n578 B.n180 163.367
R716 B.n578 B.n175 163.367
R717 B.n586 B.n175 163.367
R718 B.n586 B.n173 163.367
R719 B.n590 B.n173 163.367
R720 B.n590 B.n167 163.367
R721 B.n598 B.n167 163.367
R722 B.n598 B.n165 163.367
R723 B.n602 B.n165 163.367
R724 B.n602 B.n159 163.367
R725 B.n611 B.n159 163.367
R726 B.n611 B.n157 163.367
R727 B.n615 B.n157 163.367
R728 B.n615 B.n152 163.367
R729 B.n623 B.n152 163.367
R730 B.n623 B.n150 163.367
R731 B.n627 B.n150 163.367
R732 B.n627 B.n144 163.367
R733 B.n636 B.n144 163.367
R734 B.n636 B.n142 163.367
R735 B.n640 B.n142 163.367
R736 B.n640 B.n2 163.367
R737 B.n1021 B.n2 163.367
R738 B.n1021 B.n3 163.367
R739 B.n1017 B.n3 163.367
R740 B.n1017 B.n9 163.367
R741 B.n1013 B.n9 163.367
R742 B.n1013 B.n11 163.367
R743 B.n1009 B.n11 163.367
R744 B.n1009 B.n16 163.367
R745 B.n1005 B.n16 163.367
R746 B.n1005 B.n18 163.367
R747 B.n1001 B.n18 163.367
R748 B.n1001 B.n22 163.367
R749 B.n997 B.n22 163.367
R750 B.n997 B.n24 163.367
R751 B.n993 B.n24 163.367
R752 B.n993 B.n30 163.367
R753 B.n989 B.n30 163.367
R754 B.n989 B.n32 163.367
R755 B.n985 B.n32 163.367
R756 B.n985 B.n37 163.367
R757 B.n981 B.n37 163.367
R758 B.n981 B.n39 163.367
R759 B.n977 B.n39 163.367
R760 B.n977 B.n43 163.367
R761 B.n973 B.n43 163.367
R762 B.n973 B.n45 163.367
R763 B.n969 B.n45 163.367
R764 B.n969 B.n51 163.367
R765 B.n965 B.n51 163.367
R766 B.n965 B.n53 163.367
R767 B.n961 B.n53 163.367
R768 B.n961 B.n58 163.367
R769 B.n957 B.n58 163.367
R770 B.n957 B.n60 163.367
R771 B.n953 B.n60 163.367
R772 B.n953 B.n65 163.367
R773 B.n949 B.n65 163.367
R774 B.n949 B.n67 163.367
R775 B.n945 B.n67 163.367
R776 B.n525 B.n523 163.367
R777 B.n523 B.n522 163.367
R778 B.n519 B.n518 163.367
R779 B.n516 B.n216 163.367
R780 B.n512 B.n510 163.367
R781 B.n508 B.n218 163.367
R782 B.n504 B.n502 163.367
R783 B.n500 B.n220 163.367
R784 B.n496 B.n494 163.367
R785 B.n492 B.n222 163.367
R786 B.n488 B.n486 163.367
R787 B.n484 B.n224 163.367
R788 B.n480 B.n478 163.367
R789 B.n476 B.n226 163.367
R790 B.n472 B.n470 163.367
R791 B.n468 B.n228 163.367
R792 B.n464 B.n462 163.367
R793 B.n460 B.n230 163.367
R794 B.n456 B.n454 163.367
R795 B.n452 B.n232 163.367
R796 B.n448 B.n446 163.367
R797 B.n444 B.n234 163.367
R798 B.n440 B.n438 163.367
R799 B.n436 B.n236 163.367
R800 B.n432 B.n430 163.367
R801 B.n428 B.n238 163.367
R802 B.n424 B.n422 163.367
R803 B.n420 B.n240 163.367
R804 B.n416 B.n414 163.367
R805 B.n412 B.n242 163.367
R806 B.n408 B.n406 163.367
R807 B.n404 B.n247 163.367
R808 B.n400 B.n398 163.367
R809 B.n396 B.n249 163.367
R810 B.n391 B.n389 163.367
R811 B.n387 B.n253 163.367
R812 B.n383 B.n381 163.367
R813 B.n379 B.n255 163.367
R814 B.n375 B.n373 163.367
R815 B.n371 B.n257 163.367
R816 B.n367 B.n365 163.367
R817 B.n363 B.n259 163.367
R818 B.n359 B.n357 163.367
R819 B.n355 B.n261 163.367
R820 B.n351 B.n349 163.367
R821 B.n347 B.n263 163.367
R822 B.n343 B.n341 163.367
R823 B.n339 B.n265 163.367
R824 B.n335 B.n333 163.367
R825 B.n331 B.n267 163.367
R826 B.n327 B.n325 163.367
R827 B.n323 B.n269 163.367
R828 B.n319 B.n317 163.367
R829 B.n315 B.n271 163.367
R830 B.n311 B.n309 163.367
R831 B.n307 B.n273 163.367
R832 B.n303 B.n301 163.367
R833 B.n299 B.n275 163.367
R834 B.n295 B.n293 163.367
R835 B.n291 B.n277 163.367
R836 B.n287 B.n285 163.367
R837 B.n283 B.n280 163.367
R838 B.n531 B.n208 163.367
R839 B.n535 B.n208 163.367
R840 B.n535 B.n202 163.367
R841 B.n543 B.n202 163.367
R842 B.n543 B.n200 163.367
R843 B.n547 B.n200 163.367
R844 B.n547 B.n194 163.367
R845 B.n555 B.n194 163.367
R846 B.n555 B.n192 163.367
R847 B.n559 B.n192 163.367
R848 B.n559 B.n186 163.367
R849 B.n567 B.n186 163.367
R850 B.n567 B.n184 163.367
R851 B.n571 B.n184 163.367
R852 B.n571 B.n179 163.367
R853 B.n580 B.n179 163.367
R854 B.n580 B.n177 163.367
R855 B.n584 B.n177 163.367
R856 B.n584 B.n170 163.367
R857 B.n592 B.n170 163.367
R858 B.n592 B.n168 163.367
R859 B.n596 B.n168 163.367
R860 B.n596 B.n163 163.367
R861 B.n604 B.n163 163.367
R862 B.n604 B.n161 163.367
R863 B.n608 B.n161 163.367
R864 B.n608 B.n156 163.367
R865 B.n617 B.n156 163.367
R866 B.n617 B.n154 163.367
R867 B.n621 B.n154 163.367
R868 B.n621 B.n147 163.367
R869 B.n629 B.n147 163.367
R870 B.n629 B.n145 163.367
R871 B.n634 B.n145 163.367
R872 B.n634 B.n140 163.367
R873 B.n642 B.n140 163.367
R874 B.n643 B.n642 163.367
R875 B.n643 B.n5 163.367
R876 B.n6 B.n5 163.367
R877 B.n7 B.n6 163.367
R878 B.n648 B.n7 163.367
R879 B.n648 B.n12 163.367
R880 B.n13 B.n12 163.367
R881 B.n14 B.n13 163.367
R882 B.n653 B.n14 163.367
R883 B.n653 B.n19 163.367
R884 B.n20 B.n19 163.367
R885 B.n21 B.n20 163.367
R886 B.n658 B.n21 163.367
R887 B.n658 B.n26 163.367
R888 B.n27 B.n26 163.367
R889 B.n28 B.n27 163.367
R890 B.n663 B.n28 163.367
R891 B.n663 B.n33 163.367
R892 B.n34 B.n33 163.367
R893 B.n35 B.n34 163.367
R894 B.n668 B.n35 163.367
R895 B.n668 B.n40 163.367
R896 B.n41 B.n40 163.367
R897 B.n42 B.n41 163.367
R898 B.n673 B.n42 163.367
R899 B.n673 B.n47 163.367
R900 B.n48 B.n47 163.367
R901 B.n49 B.n48 163.367
R902 B.n678 B.n49 163.367
R903 B.n678 B.n54 163.367
R904 B.n55 B.n54 163.367
R905 B.n56 B.n55 163.367
R906 B.n683 B.n56 163.367
R907 B.n683 B.n61 163.367
R908 B.n62 B.n61 163.367
R909 B.n63 B.n62 163.367
R910 B.n688 B.n63 163.367
R911 B.n688 B.n68 163.367
R912 B.n69 B.n68 163.367
R913 B.n70 B.n69 163.367
R914 B.n941 B.n939 163.367
R915 B.n937 B.n74 163.367
R916 B.n933 B.n931 163.367
R917 B.n929 B.n76 163.367
R918 B.n925 B.n923 163.367
R919 B.n921 B.n78 163.367
R920 B.n917 B.n915 163.367
R921 B.n913 B.n80 163.367
R922 B.n909 B.n907 163.367
R923 B.n905 B.n82 163.367
R924 B.n901 B.n899 163.367
R925 B.n897 B.n84 163.367
R926 B.n893 B.n891 163.367
R927 B.n889 B.n86 163.367
R928 B.n885 B.n883 163.367
R929 B.n881 B.n88 163.367
R930 B.n877 B.n875 163.367
R931 B.n873 B.n90 163.367
R932 B.n869 B.n867 163.367
R933 B.n865 B.n92 163.367
R934 B.n861 B.n859 163.367
R935 B.n857 B.n94 163.367
R936 B.n853 B.n851 163.367
R937 B.n849 B.n96 163.367
R938 B.n845 B.n843 163.367
R939 B.n841 B.n98 163.367
R940 B.n837 B.n835 163.367
R941 B.n833 B.n100 163.367
R942 B.n829 B.n827 163.367
R943 B.n824 B.n823 163.367
R944 B.n821 B.n106 163.367
R945 B.n817 B.n815 163.367
R946 B.n813 B.n108 163.367
R947 B.n808 B.n806 163.367
R948 B.n804 B.n112 163.367
R949 B.n800 B.n798 163.367
R950 B.n796 B.n114 163.367
R951 B.n792 B.n790 163.367
R952 B.n788 B.n116 163.367
R953 B.n784 B.n782 163.367
R954 B.n780 B.n118 163.367
R955 B.n776 B.n774 163.367
R956 B.n772 B.n120 163.367
R957 B.n768 B.n766 163.367
R958 B.n764 B.n122 163.367
R959 B.n760 B.n758 163.367
R960 B.n756 B.n124 163.367
R961 B.n752 B.n750 163.367
R962 B.n748 B.n126 163.367
R963 B.n744 B.n742 163.367
R964 B.n740 B.n128 163.367
R965 B.n736 B.n734 163.367
R966 B.n732 B.n130 163.367
R967 B.n728 B.n726 163.367
R968 B.n724 B.n132 163.367
R969 B.n720 B.n718 163.367
R970 B.n716 B.n134 163.367
R971 B.n712 B.n710 163.367
R972 B.n708 B.n136 163.367
R973 B.n704 B.n702 163.367
R974 B.n700 B.n138 163.367
R975 B.n696 B.n694 163.367
R976 B.n524 B.n212 71.676
R977 B.n522 B.n214 71.676
R978 B.n518 B.n517 71.676
R979 B.n511 B.n216 71.676
R980 B.n510 B.n509 71.676
R981 B.n503 B.n218 71.676
R982 B.n502 B.n501 71.676
R983 B.n495 B.n220 71.676
R984 B.n494 B.n493 71.676
R985 B.n487 B.n222 71.676
R986 B.n486 B.n485 71.676
R987 B.n479 B.n224 71.676
R988 B.n478 B.n477 71.676
R989 B.n471 B.n226 71.676
R990 B.n470 B.n469 71.676
R991 B.n463 B.n228 71.676
R992 B.n462 B.n461 71.676
R993 B.n455 B.n230 71.676
R994 B.n454 B.n453 71.676
R995 B.n447 B.n232 71.676
R996 B.n446 B.n445 71.676
R997 B.n439 B.n234 71.676
R998 B.n438 B.n437 71.676
R999 B.n431 B.n236 71.676
R1000 B.n430 B.n429 71.676
R1001 B.n423 B.n238 71.676
R1002 B.n422 B.n421 71.676
R1003 B.n415 B.n240 71.676
R1004 B.n414 B.n413 71.676
R1005 B.n407 B.n242 71.676
R1006 B.n406 B.n405 71.676
R1007 B.n399 B.n247 71.676
R1008 B.n398 B.n397 71.676
R1009 B.n390 B.n249 71.676
R1010 B.n389 B.n388 71.676
R1011 B.n382 B.n253 71.676
R1012 B.n381 B.n380 71.676
R1013 B.n374 B.n255 71.676
R1014 B.n373 B.n372 71.676
R1015 B.n366 B.n257 71.676
R1016 B.n365 B.n364 71.676
R1017 B.n358 B.n259 71.676
R1018 B.n357 B.n356 71.676
R1019 B.n350 B.n261 71.676
R1020 B.n349 B.n348 71.676
R1021 B.n342 B.n263 71.676
R1022 B.n341 B.n340 71.676
R1023 B.n334 B.n265 71.676
R1024 B.n333 B.n332 71.676
R1025 B.n326 B.n267 71.676
R1026 B.n325 B.n324 71.676
R1027 B.n318 B.n269 71.676
R1028 B.n317 B.n316 71.676
R1029 B.n310 B.n271 71.676
R1030 B.n309 B.n308 71.676
R1031 B.n302 B.n273 71.676
R1032 B.n301 B.n300 71.676
R1033 B.n294 B.n275 71.676
R1034 B.n293 B.n292 71.676
R1035 B.n286 B.n277 71.676
R1036 B.n285 B.n284 71.676
R1037 B.n280 B.n279 71.676
R1038 B.n940 B.n72 71.676
R1039 B.n939 B.n938 71.676
R1040 B.n932 B.n74 71.676
R1041 B.n931 B.n930 71.676
R1042 B.n924 B.n76 71.676
R1043 B.n923 B.n922 71.676
R1044 B.n916 B.n78 71.676
R1045 B.n915 B.n914 71.676
R1046 B.n908 B.n80 71.676
R1047 B.n907 B.n906 71.676
R1048 B.n900 B.n82 71.676
R1049 B.n899 B.n898 71.676
R1050 B.n892 B.n84 71.676
R1051 B.n891 B.n890 71.676
R1052 B.n884 B.n86 71.676
R1053 B.n883 B.n882 71.676
R1054 B.n876 B.n88 71.676
R1055 B.n875 B.n874 71.676
R1056 B.n868 B.n90 71.676
R1057 B.n867 B.n866 71.676
R1058 B.n860 B.n92 71.676
R1059 B.n859 B.n858 71.676
R1060 B.n852 B.n94 71.676
R1061 B.n851 B.n850 71.676
R1062 B.n844 B.n96 71.676
R1063 B.n843 B.n842 71.676
R1064 B.n836 B.n98 71.676
R1065 B.n835 B.n834 71.676
R1066 B.n828 B.n100 71.676
R1067 B.n827 B.n104 71.676
R1068 B.n823 B.n822 71.676
R1069 B.n816 B.n106 71.676
R1070 B.n815 B.n814 71.676
R1071 B.n807 B.n108 71.676
R1072 B.n806 B.n805 71.676
R1073 B.n799 B.n112 71.676
R1074 B.n798 B.n797 71.676
R1075 B.n791 B.n114 71.676
R1076 B.n790 B.n789 71.676
R1077 B.n783 B.n116 71.676
R1078 B.n782 B.n781 71.676
R1079 B.n775 B.n118 71.676
R1080 B.n774 B.n773 71.676
R1081 B.n767 B.n120 71.676
R1082 B.n766 B.n765 71.676
R1083 B.n759 B.n122 71.676
R1084 B.n758 B.n757 71.676
R1085 B.n751 B.n124 71.676
R1086 B.n750 B.n749 71.676
R1087 B.n743 B.n126 71.676
R1088 B.n742 B.n741 71.676
R1089 B.n735 B.n128 71.676
R1090 B.n734 B.n733 71.676
R1091 B.n727 B.n130 71.676
R1092 B.n726 B.n725 71.676
R1093 B.n719 B.n132 71.676
R1094 B.n718 B.n717 71.676
R1095 B.n711 B.n134 71.676
R1096 B.n710 B.n709 71.676
R1097 B.n703 B.n136 71.676
R1098 B.n702 B.n701 71.676
R1099 B.n695 B.n138 71.676
R1100 B.n696 B.n695 71.676
R1101 B.n701 B.n700 71.676
R1102 B.n704 B.n703 71.676
R1103 B.n709 B.n708 71.676
R1104 B.n712 B.n711 71.676
R1105 B.n717 B.n716 71.676
R1106 B.n720 B.n719 71.676
R1107 B.n725 B.n724 71.676
R1108 B.n728 B.n727 71.676
R1109 B.n733 B.n732 71.676
R1110 B.n736 B.n735 71.676
R1111 B.n741 B.n740 71.676
R1112 B.n744 B.n743 71.676
R1113 B.n749 B.n748 71.676
R1114 B.n752 B.n751 71.676
R1115 B.n757 B.n756 71.676
R1116 B.n760 B.n759 71.676
R1117 B.n765 B.n764 71.676
R1118 B.n768 B.n767 71.676
R1119 B.n773 B.n772 71.676
R1120 B.n776 B.n775 71.676
R1121 B.n781 B.n780 71.676
R1122 B.n784 B.n783 71.676
R1123 B.n789 B.n788 71.676
R1124 B.n792 B.n791 71.676
R1125 B.n797 B.n796 71.676
R1126 B.n800 B.n799 71.676
R1127 B.n805 B.n804 71.676
R1128 B.n808 B.n807 71.676
R1129 B.n814 B.n813 71.676
R1130 B.n817 B.n816 71.676
R1131 B.n822 B.n821 71.676
R1132 B.n824 B.n104 71.676
R1133 B.n829 B.n828 71.676
R1134 B.n834 B.n833 71.676
R1135 B.n837 B.n836 71.676
R1136 B.n842 B.n841 71.676
R1137 B.n845 B.n844 71.676
R1138 B.n850 B.n849 71.676
R1139 B.n853 B.n852 71.676
R1140 B.n858 B.n857 71.676
R1141 B.n861 B.n860 71.676
R1142 B.n866 B.n865 71.676
R1143 B.n869 B.n868 71.676
R1144 B.n874 B.n873 71.676
R1145 B.n877 B.n876 71.676
R1146 B.n882 B.n881 71.676
R1147 B.n885 B.n884 71.676
R1148 B.n890 B.n889 71.676
R1149 B.n893 B.n892 71.676
R1150 B.n898 B.n897 71.676
R1151 B.n901 B.n900 71.676
R1152 B.n906 B.n905 71.676
R1153 B.n909 B.n908 71.676
R1154 B.n914 B.n913 71.676
R1155 B.n917 B.n916 71.676
R1156 B.n922 B.n921 71.676
R1157 B.n925 B.n924 71.676
R1158 B.n930 B.n929 71.676
R1159 B.n933 B.n932 71.676
R1160 B.n938 B.n937 71.676
R1161 B.n941 B.n940 71.676
R1162 B.n525 B.n524 71.676
R1163 B.n519 B.n214 71.676
R1164 B.n517 B.n516 71.676
R1165 B.n512 B.n511 71.676
R1166 B.n509 B.n508 71.676
R1167 B.n504 B.n503 71.676
R1168 B.n501 B.n500 71.676
R1169 B.n496 B.n495 71.676
R1170 B.n493 B.n492 71.676
R1171 B.n488 B.n487 71.676
R1172 B.n485 B.n484 71.676
R1173 B.n480 B.n479 71.676
R1174 B.n477 B.n476 71.676
R1175 B.n472 B.n471 71.676
R1176 B.n469 B.n468 71.676
R1177 B.n464 B.n463 71.676
R1178 B.n461 B.n460 71.676
R1179 B.n456 B.n455 71.676
R1180 B.n453 B.n452 71.676
R1181 B.n448 B.n447 71.676
R1182 B.n445 B.n444 71.676
R1183 B.n440 B.n439 71.676
R1184 B.n437 B.n436 71.676
R1185 B.n432 B.n431 71.676
R1186 B.n429 B.n428 71.676
R1187 B.n424 B.n423 71.676
R1188 B.n421 B.n420 71.676
R1189 B.n416 B.n415 71.676
R1190 B.n413 B.n412 71.676
R1191 B.n408 B.n407 71.676
R1192 B.n405 B.n404 71.676
R1193 B.n400 B.n399 71.676
R1194 B.n397 B.n396 71.676
R1195 B.n391 B.n390 71.676
R1196 B.n388 B.n387 71.676
R1197 B.n383 B.n382 71.676
R1198 B.n380 B.n379 71.676
R1199 B.n375 B.n374 71.676
R1200 B.n372 B.n371 71.676
R1201 B.n367 B.n366 71.676
R1202 B.n364 B.n363 71.676
R1203 B.n359 B.n358 71.676
R1204 B.n356 B.n355 71.676
R1205 B.n351 B.n350 71.676
R1206 B.n348 B.n347 71.676
R1207 B.n343 B.n342 71.676
R1208 B.n340 B.n339 71.676
R1209 B.n335 B.n334 71.676
R1210 B.n332 B.n331 71.676
R1211 B.n327 B.n326 71.676
R1212 B.n324 B.n323 71.676
R1213 B.n319 B.n318 71.676
R1214 B.n316 B.n315 71.676
R1215 B.n311 B.n310 71.676
R1216 B.n308 B.n307 71.676
R1217 B.n303 B.n302 71.676
R1218 B.n300 B.n299 71.676
R1219 B.n295 B.n294 71.676
R1220 B.n292 B.n291 71.676
R1221 B.n287 B.n286 71.676
R1222 B.n284 B.n283 71.676
R1223 B.n279 B.n210 71.676
R1224 B.n394 B.n251 59.5399
R1225 B.n245 B.n244 59.5399
R1226 B.n103 B.n102 59.5399
R1227 B.n810 B.n110 59.5399
R1228 B.n530 B.n211 53.7299
R1229 B.n946 B.n71 53.7299
R1230 B.n251 B.n250 39.1763
R1231 B.n244 B.n243 39.1763
R1232 B.n102 B.n101 39.1763
R1233 B.n110 B.n109 39.1763
R1234 B.n530 B.n207 32.9158
R1235 B.n536 B.n207 32.9158
R1236 B.n536 B.n203 32.9158
R1237 B.n542 B.n203 32.9158
R1238 B.n542 B.n199 32.9158
R1239 B.n548 B.n199 32.9158
R1240 B.n554 B.n195 32.9158
R1241 B.n554 B.n191 32.9158
R1242 B.n560 B.n191 32.9158
R1243 B.n560 B.n187 32.9158
R1244 B.n566 B.n187 32.9158
R1245 B.n566 B.n183 32.9158
R1246 B.n573 B.n183 32.9158
R1247 B.n573 B.n572 32.9158
R1248 B.n579 B.n176 32.9158
R1249 B.n585 B.n176 32.9158
R1250 B.n585 B.n171 32.9158
R1251 B.n591 B.n171 32.9158
R1252 B.n591 B.n172 32.9158
R1253 B.n597 B.n164 32.9158
R1254 B.n603 B.n164 32.9158
R1255 B.n603 B.n160 32.9158
R1256 B.n610 B.n160 32.9158
R1257 B.n610 B.n609 32.9158
R1258 B.n616 B.n153 32.9158
R1259 B.n622 B.n153 32.9158
R1260 B.n622 B.n148 32.9158
R1261 B.n628 B.n148 32.9158
R1262 B.n628 B.n149 32.9158
R1263 B.n635 B.n141 32.9158
R1264 B.n641 B.n141 32.9158
R1265 B.n641 B.n4 32.9158
R1266 B.n1020 B.n4 32.9158
R1267 B.n1020 B.n1019 32.9158
R1268 B.n1019 B.n1018 32.9158
R1269 B.n1018 B.n8 32.9158
R1270 B.n1012 B.n8 32.9158
R1271 B.n1011 B.n1010 32.9158
R1272 B.n1010 B.n15 32.9158
R1273 B.n1004 B.n15 32.9158
R1274 B.n1004 B.n1003 32.9158
R1275 B.n1003 B.n1002 32.9158
R1276 B.n996 B.n25 32.9158
R1277 B.n996 B.n995 32.9158
R1278 B.n995 B.n994 32.9158
R1279 B.n994 B.n29 32.9158
R1280 B.n988 B.n29 32.9158
R1281 B.n987 B.n986 32.9158
R1282 B.n986 B.n36 32.9158
R1283 B.n980 B.n36 32.9158
R1284 B.n980 B.n979 32.9158
R1285 B.n979 B.n978 32.9158
R1286 B.n972 B.n46 32.9158
R1287 B.n972 B.n971 32.9158
R1288 B.n971 B.n970 32.9158
R1289 B.n970 B.n50 32.9158
R1290 B.n964 B.n50 32.9158
R1291 B.n964 B.n963 32.9158
R1292 B.n963 B.n962 32.9158
R1293 B.n962 B.n57 32.9158
R1294 B.n956 B.n955 32.9158
R1295 B.n955 B.n954 32.9158
R1296 B.n954 B.n64 32.9158
R1297 B.n948 B.n64 32.9158
R1298 B.n948 B.n947 32.9158
R1299 B.n947 B.n946 32.9158
R1300 B.n944 B.n943 29.8151
R1301 B.n532 B.n209 29.8151
R1302 B.n528 B.n527 29.8151
R1303 B.n693 B.n692 29.8151
R1304 B.n572 B.t4 19.8465
R1305 B.n46 B.t5 19.8465
R1306 B.n635 B.t3 18.8784
R1307 B.n1012 B.t6 18.8784
R1308 B B.n1022 18.0485
R1309 B.t13 B.n195 17.9103
R1310 B.n172 B.t7 17.9103
R1311 B.t1 B.n987 17.9103
R1312 B.t9 B.n57 17.9103
R1313 B.n616 B.t2 16.9422
R1314 B.n1002 B.t0 16.9422
R1315 B.n609 B.t2 15.9741
R1316 B.n25 B.t0 15.9741
R1317 B.n548 B.t13 15.006
R1318 B.n597 B.t7 15.006
R1319 B.n988 B.t1 15.006
R1320 B.n956 B.t9 15.006
R1321 B.n149 B.t3 14.0379
R1322 B.t6 B.n1011 14.0379
R1323 B.n579 B.t4 13.0698
R1324 B.n978 B.t5 13.0698
R1325 B.n943 B.n942 10.6151
R1326 B.n942 B.n73 10.6151
R1327 B.n936 B.n73 10.6151
R1328 B.n936 B.n935 10.6151
R1329 B.n935 B.n934 10.6151
R1330 B.n934 B.n75 10.6151
R1331 B.n928 B.n75 10.6151
R1332 B.n928 B.n927 10.6151
R1333 B.n927 B.n926 10.6151
R1334 B.n926 B.n77 10.6151
R1335 B.n920 B.n77 10.6151
R1336 B.n920 B.n919 10.6151
R1337 B.n919 B.n918 10.6151
R1338 B.n918 B.n79 10.6151
R1339 B.n912 B.n79 10.6151
R1340 B.n912 B.n911 10.6151
R1341 B.n911 B.n910 10.6151
R1342 B.n910 B.n81 10.6151
R1343 B.n904 B.n81 10.6151
R1344 B.n904 B.n903 10.6151
R1345 B.n903 B.n902 10.6151
R1346 B.n902 B.n83 10.6151
R1347 B.n896 B.n83 10.6151
R1348 B.n896 B.n895 10.6151
R1349 B.n895 B.n894 10.6151
R1350 B.n894 B.n85 10.6151
R1351 B.n888 B.n85 10.6151
R1352 B.n888 B.n887 10.6151
R1353 B.n887 B.n886 10.6151
R1354 B.n886 B.n87 10.6151
R1355 B.n880 B.n87 10.6151
R1356 B.n880 B.n879 10.6151
R1357 B.n879 B.n878 10.6151
R1358 B.n878 B.n89 10.6151
R1359 B.n872 B.n89 10.6151
R1360 B.n872 B.n871 10.6151
R1361 B.n871 B.n870 10.6151
R1362 B.n870 B.n91 10.6151
R1363 B.n864 B.n91 10.6151
R1364 B.n864 B.n863 10.6151
R1365 B.n863 B.n862 10.6151
R1366 B.n862 B.n93 10.6151
R1367 B.n856 B.n93 10.6151
R1368 B.n856 B.n855 10.6151
R1369 B.n855 B.n854 10.6151
R1370 B.n854 B.n95 10.6151
R1371 B.n848 B.n95 10.6151
R1372 B.n848 B.n847 10.6151
R1373 B.n847 B.n846 10.6151
R1374 B.n846 B.n97 10.6151
R1375 B.n840 B.n97 10.6151
R1376 B.n840 B.n839 10.6151
R1377 B.n839 B.n838 10.6151
R1378 B.n838 B.n99 10.6151
R1379 B.n832 B.n99 10.6151
R1380 B.n832 B.n831 10.6151
R1381 B.n831 B.n830 10.6151
R1382 B.n826 B.n825 10.6151
R1383 B.n825 B.n105 10.6151
R1384 B.n820 B.n105 10.6151
R1385 B.n820 B.n819 10.6151
R1386 B.n819 B.n818 10.6151
R1387 B.n818 B.n107 10.6151
R1388 B.n812 B.n107 10.6151
R1389 B.n812 B.n811 10.6151
R1390 B.n809 B.n111 10.6151
R1391 B.n803 B.n111 10.6151
R1392 B.n803 B.n802 10.6151
R1393 B.n802 B.n801 10.6151
R1394 B.n801 B.n113 10.6151
R1395 B.n795 B.n113 10.6151
R1396 B.n795 B.n794 10.6151
R1397 B.n794 B.n793 10.6151
R1398 B.n793 B.n115 10.6151
R1399 B.n787 B.n115 10.6151
R1400 B.n787 B.n786 10.6151
R1401 B.n786 B.n785 10.6151
R1402 B.n785 B.n117 10.6151
R1403 B.n779 B.n117 10.6151
R1404 B.n779 B.n778 10.6151
R1405 B.n778 B.n777 10.6151
R1406 B.n777 B.n119 10.6151
R1407 B.n771 B.n119 10.6151
R1408 B.n771 B.n770 10.6151
R1409 B.n770 B.n769 10.6151
R1410 B.n769 B.n121 10.6151
R1411 B.n763 B.n121 10.6151
R1412 B.n763 B.n762 10.6151
R1413 B.n762 B.n761 10.6151
R1414 B.n761 B.n123 10.6151
R1415 B.n755 B.n123 10.6151
R1416 B.n755 B.n754 10.6151
R1417 B.n754 B.n753 10.6151
R1418 B.n753 B.n125 10.6151
R1419 B.n747 B.n125 10.6151
R1420 B.n747 B.n746 10.6151
R1421 B.n746 B.n745 10.6151
R1422 B.n745 B.n127 10.6151
R1423 B.n739 B.n127 10.6151
R1424 B.n739 B.n738 10.6151
R1425 B.n738 B.n737 10.6151
R1426 B.n737 B.n129 10.6151
R1427 B.n731 B.n129 10.6151
R1428 B.n731 B.n730 10.6151
R1429 B.n730 B.n729 10.6151
R1430 B.n729 B.n131 10.6151
R1431 B.n723 B.n131 10.6151
R1432 B.n723 B.n722 10.6151
R1433 B.n722 B.n721 10.6151
R1434 B.n721 B.n133 10.6151
R1435 B.n715 B.n133 10.6151
R1436 B.n715 B.n714 10.6151
R1437 B.n714 B.n713 10.6151
R1438 B.n713 B.n135 10.6151
R1439 B.n707 B.n135 10.6151
R1440 B.n707 B.n706 10.6151
R1441 B.n706 B.n705 10.6151
R1442 B.n705 B.n137 10.6151
R1443 B.n699 B.n137 10.6151
R1444 B.n699 B.n698 10.6151
R1445 B.n698 B.n697 10.6151
R1446 B.n697 B.n693 10.6151
R1447 B.n533 B.n532 10.6151
R1448 B.n534 B.n533 10.6151
R1449 B.n534 B.n201 10.6151
R1450 B.n544 B.n201 10.6151
R1451 B.n545 B.n544 10.6151
R1452 B.n546 B.n545 10.6151
R1453 B.n546 B.n193 10.6151
R1454 B.n556 B.n193 10.6151
R1455 B.n557 B.n556 10.6151
R1456 B.n558 B.n557 10.6151
R1457 B.n558 B.n185 10.6151
R1458 B.n568 B.n185 10.6151
R1459 B.n569 B.n568 10.6151
R1460 B.n570 B.n569 10.6151
R1461 B.n570 B.n178 10.6151
R1462 B.n581 B.n178 10.6151
R1463 B.n582 B.n581 10.6151
R1464 B.n583 B.n582 10.6151
R1465 B.n583 B.n169 10.6151
R1466 B.n593 B.n169 10.6151
R1467 B.n594 B.n593 10.6151
R1468 B.n595 B.n594 10.6151
R1469 B.n595 B.n162 10.6151
R1470 B.n605 B.n162 10.6151
R1471 B.n606 B.n605 10.6151
R1472 B.n607 B.n606 10.6151
R1473 B.n607 B.n155 10.6151
R1474 B.n618 B.n155 10.6151
R1475 B.n619 B.n618 10.6151
R1476 B.n620 B.n619 10.6151
R1477 B.n620 B.n146 10.6151
R1478 B.n630 B.n146 10.6151
R1479 B.n631 B.n630 10.6151
R1480 B.n633 B.n631 10.6151
R1481 B.n633 B.n632 10.6151
R1482 B.n632 B.n139 10.6151
R1483 B.n644 B.n139 10.6151
R1484 B.n645 B.n644 10.6151
R1485 B.n646 B.n645 10.6151
R1486 B.n647 B.n646 10.6151
R1487 B.n649 B.n647 10.6151
R1488 B.n650 B.n649 10.6151
R1489 B.n651 B.n650 10.6151
R1490 B.n652 B.n651 10.6151
R1491 B.n654 B.n652 10.6151
R1492 B.n655 B.n654 10.6151
R1493 B.n656 B.n655 10.6151
R1494 B.n657 B.n656 10.6151
R1495 B.n659 B.n657 10.6151
R1496 B.n660 B.n659 10.6151
R1497 B.n661 B.n660 10.6151
R1498 B.n662 B.n661 10.6151
R1499 B.n664 B.n662 10.6151
R1500 B.n665 B.n664 10.6151
R1501 B.n666 B.n665 10.6151
R1502 B.n667 B.n666 10.6151
R1503 B.n669 B.n667 10.6151
R1504 B.n670 B.n669 10.6151
R1505 B.n671 B.n670 10.6151
R1506 B.n672 B.n671 10.6151
R1507 B.n674 B.n672 10.6151
R1508 B.n675 B.n674 10.6151
R1509 B.n676 B.n675 10.6151
R1510 B.n677 B.n676 10.6151
R1511 B.n679 B.n677 10.6151
R1512 B.n680 B.n679 10.6151
R1513 B.n681 B.n680 10.6151
R1514 B.n682 B.n681 10.6151
R1515 B.n684 B.n682 10.6151
R1516 B.n685 B.n684 10.6151
R1517 B.n686 B.n685 10.6151
R1518 B.n687 B.n686 10.6151
R1519 B.n689 B.n687 10.6151
R1520 B.n690 B.n689 10.6151
R1521 B.n691 B.n690 10.6151
R1522 B.n692 B.n691 10.6151
R1523 B.n527 B.n526 10.6151
R1524 B.n526 B.n213 10.6151
R1525 B.n521 B.n213 10.6151
R1526 B.n521 B.n520 10.6151
R1527 B.n520 B.n215 10.6151
R1528 B.n515 B.n215 10.6151
R1529 B.n515 B.n514 10.6151
R1530 B.n514 B.n513 10.6151
R1531 B.n513 B.n217 10.6151
R1532 B.n507 B.n217 10.6151
R1533 B.n507 B.n506 10.6151
R1534 B.n506 B.n505 10.6151
R1535 B.n505 B.n219 10.6151
R1536 B.n499 B.n219 10.6151
R1537 B.n499 B.n498 10.6151
R1538 B.n498 B.n497 10.6151
R1539 B.n497 B.n221 10.6151
R1540 B.n491 B.n221 10.6151
R1541 B.n491 B.n490 10.6151
R1542 B.n490 B.n489 10.6151
R1543 B.n489 B.n223 10.6151
R1544 B.n483 B.n223 10.6151
R1545 B.n483 B.n482 10.6151
R1546 B.n482 B.n481 10.6151
R1547 B.n481 B.n225 10.6151
R1548 B.n475 B.n225 10.6151
R1549 B.n475 B.n474 10.6151
R1550 B.n474 B.n473 10.6151
R1551 B.n473 B.n227 10.6151
R1552 B.n467 B.n227 10.6151
R1553 B.n467 B.n466 10.6151
R1554 B.n466 B.n465 10.6151
R1555 B.n465 B.n229 10.6151
R1556 B.n459 B.n229 10.6151
R1557 B.n459 B.n458 10.6151
R1558 B.n458 B.n457 10.6151
R1559 B.n457 B.n231 10.6151
R1560 B.n451 B.n231 10.6151
R1561 B.n451 B.n450 10.6151
R1562 B.n450 B.n449 10.6151
R1563 B.n449 B.n233 10.6151
R1564 B.n443 B.n233 10.6151
R1565 B.n443 B.n442 10.6151
R1566 B.n442 B.n441 10.6151
R1567 B.n441 B.n235 10.6151
R1568 B.n435 B.n235 10.6151
R1569 B.n435 B.n434 10.6151
R1570 B.n434 B.n433 10.6151
R1571 B.n433 B.n237 10.6151
R1572 B.n427 B.n237 10.6151
R1573 B.n427 B.n426 10.6151
R1574 B.n426 B.n425 10.6151
R1575 B.n425 B.n239 10.6151
R1576 B.n419 B.n239 10.6151
R1577 B.n419 B.n418 10.6151
R1578 B.n418 B.n417 10.6151
R1579 B.n417 B.n241 10.6151
R1580 B.n411 B.n410 10.6151
R1581 B.n410 B.n409 10.6151
R1582 B.n409 B.n246 10.6151
R1583 B.n403 B.n246 10.6151
R1584 B.n403 B.n402 10.6151
R1585 B.n402 B.n401 10.6151
R1586 B.n401 B.n248 10.6151
R1587 B.n395 B.n248 10.6151
R1588 B.n393 B.n392 10.6151
R1589 B.n392 B.n252 10.6151
R1590 B.n386 B.n252 10.6151
R1591 B.n386 B.n385 10.6151
R1592 B.n385 B.n384 10.6151
R1593 B.n384 B.n254 10.6151
R1594 B.n378 B.n254 10.6151
R1595 B.n378 B.n377 10.6151
R1596 B.n377 B.n376 10.6151
R1597 B.n376 B.n256 10.6151
R1598 B.n370 B.n256 10.6151
R1599 B.n370 B.n369 10.6151
R1600 B.n369 B.n368 10.6151
R1601 B.n368 B.n258 10.6151
R1602 B.n362 B.n258 10.6151
R1603 B.n362 B.n361 10.6151
R1604 B.n361 B.n360 10.6151
R1605 B.n360 B.n260 10.6151
R1606 B.n354 B.n260 10.6151
R1607 B.n354 B.n353 10.6151
R1608 B.n353 B.n352 10.6151
R1609 B.n352 B.n262 10.6151
R1610 B.n346 B.n262 10.6151
R1611 B.n346 B.n345 10.6151
R1612 B.n345 B.n344 10.6151
R1613 B.n344 B.n264 10.6151
R1614 B.n338 B.n264 10.6151
R1615 B.n338 B.n337 10.6151
R1616 B.n337 B.n336 10.6151
R1617 B.n336 B.n266 10.6151
R1618 B.n330 B.n266 10.6151
R1619 B.n330 B.n329 10.6151
R1620 B.n329 B.n328 10.6151
R1621 B.n328 B.n268 10.6151
R1622 B.n322 B.n268 10.6151
R1623 B.n322 B.n321 10.6151
R1624 B.n321 B.n320 10.6151
R1625 B.n320 B.n270 10.6151
R1626 B.n314 B.n270 10.6151
R1627 B.n314 B.n313 10.6151
R1628 B.n313 B.n312 10.6151
R1629 B.n312 B.n272 10.6151
R1630 B.n306 B.n272 10.6151
R1631 B.n306 B.n305 10.6151
R1632 B.n305 B.n304 10.6151
R1633 B.n304 B.n274 10.6151
R1634 B.n298 B.n274 10.6151
R1635 B.n298 B.n297 10.6151
R1636 B.n297 B.n296 10.6151
R1637 B.n296 B.n276 10.6151
R1638 B.n290 B.n276 10.6151
R1639 B.n290 B.n289 10.6151
R1640 B.n289 B.n288 10.6151
R1641 B.n288 B.n278 10.6151
R1642 B.n282 B.n278 10.6151
R1643 B.n282 B.n281 10.6151
R1644 B.n281 B.n209 10.6151
R1645 B.n528 B.n205 10.6151
R1646 B.n538 B.n205 10.6151
R1647 B.n539 B.n538 10.6151
R1648 B.n540 B.n539 10.6151
R1649 B.n540 B.n197 10.6151
R1650 B.n550 B.n197 10.6151
R1651 B.n551 B.n550 10.6151
R1652 B.n552 B.n551 10.6151
R1653 B.n552 B.n189 10.6151
R1654 B.n562 B.n189 10.6151
R1655 B.n563 B.n562 10.6151
R1656 B.n564 B.n563 10.6151
R1657 B.n564 B.n181 10.6151
R1658 B.n575 B.n181 10.6151
R1659 B.n576 B.n575 10.6151
R1660 B.n577 B.n576 10.6151
R1661 B.n577 B.n174 10.6151
R1662 B.n587 B.n174 10.6151
R1663 B.n588 B.n587 10.6151
R1664 B.n589 B.n588 10.6151
R1665 B.n589 B.n166 10.6151
R1666 B.n599 B.n166 10.6151
R1667 B.n600 B.n599 10.6151
R1668 B.n601 B.n600 10.6151
R1669 B.n601 B.n158 10.6151
R1670 B.n612 B.n158 10.6151
R1671 B.n613 B.n612 10.6151
R1672 B.n614 B.n613 10.6151
R1673 B.n614 B.n151 10.6151
R1674 B.n624 B.n151 10.6151
R1675 B.n625 B.n624 10.6151
R1676 B.n626 B.n625 10.6151
R1677 B.n626 B.n143 10.6151
R1678 B.n637 B.n143 10.6151
R1679 B.n638 B.n637 10.6151
R1680 B.n639 B.n638 10.6151
R1681 B.n639 B.n0 10.6151
R1682 B.n1016 B.n1 10.6151
R1683 B.n1016 B.n1015 10.6151
R1684 B.n1015 B.n1014 10.6151
R1685 B.n1014 B.n10 10.6151
R1686 B.n1008 B.n10 10.6151
R1687 B.n1008 B.n1007 10.6151
R1688 B.n1007 B.n1006 10.6151
R1689 B.n1006 B.n17 10.6151
R1690 B.n1000 B.n17 10.6151
R1691 B.n1000 B.n999 10.6151
R1692 B.n999 B.n998 10.6151
R1693 B.n998 B.n23 10.6151
R1694 B.n992 B.n23 10.6151
R1695 B.n992 B.n991 10.6151
R1696 B.n991 B.n990 10.6151
R1697 B.n990 B.n31 10.6151
R1698 B.n984 B.n31 10.6151
R1699 B.n984 B.n983 10.6151
R1700 B.n983 B.n982 10.6151
R1701 B.n982 B.n38 10.6151
R1702 B.n976 B.n38 10.6151
R1703 B.n976 B.n975 10.6151
R1704 B.n975 B.n974 10.6151
R1705 B.n974 B.n44 10.6151
R1706 B.n968 B.n44 10.6151
R1707 B.n968 B.n967 10.6151
R1708 B.n967 B.n966 10.6151
R1709 B.n966 B.n52 10.6151
R1710 B.n960 B.n52 10.6151
R1711 B.n960 B.n959 10.6151
R1712 B.n959 B.n958 10.6151
R1713 B.n958 B.n59 10.6151
R1714 B.n952 B.n59 10.6151
R1715 B.n952 B.n951 10.6151
R1716 B.n951 B.n950 10.6151
R1717 B.n950 B.n66 10.6151
R1718 B.n944 B.n66 10.6151
R1719 B.n826 B.n103 6.5566
R1720 B.n811 B.n810 6.5566
R1721 B.n411 B.n245 6.5566
R1722 B.n395 B.n394 6.5566
R1723 B.n830 B.n103 4.05904
R1724 B.n810 B.n809 4.05904
R1725 B.n245 B.n241 4.05904
R1726 B.n394 B.n393 4.05904
R1727 B.n1022 B.n0 2.81026
R1728 B.n1022 B.n1 2.81026
R1729 VN.n5 VN.t6 276.861
R1730 VN.n28 VN.t5 276.861
R1731 VN.n6 VN.t7 248.844
R1732 VN.n14 VN.t2 248.844
R1733 VN.n21 VN.t3 248.844
R1734 VN.n29 VN.t0 248.844
R1735 VN.n37 VN.t4 248.844
R1736 VN.n44 VN.t1 248.844
R1737 VN.n22 VN.n21 184.299
R1738 VN.n45 VN.n44 184.299
R1739 VN.n43 VN.n23 161.3
R1740 VN.n42 VN.n41 161.3
R1741 VN.n40 VN.n24 161.3
R1742 VN.n39 VN.n38 161.3
R1743 VN.n36 VN.n25 161.3
R1744 VN.n35 VN.n34 161.3
R1745 VN.n33 VN.n26 161.3
R1746 VN.n32 VN.n31 161.3
R1747 VN.n30 VN.n27 161.3
R1748 VN.n20 VN.n0 161.3
R1749 VN.n19 VN.n18 161.3
R1750 VN.n17 VN.n1 161.3
R1751 VN.n16 VN.n15 161.3
R1752 VN.n13 VN.n2 161.3
R1753 VN.n12 VN.n11 161.3
R1754 VN.n10 VN.n3 161.3
R1755 VN.n9 VN.n8 161.3
R1756 VN.n7 VN.n4 161.3
R1757 VN.n6 VN.n5 68.3373
R1758 VN.n29 VN.n28 68.3373
R1759 VN VN.n45 50.9872
R1760 VN.n19 VN.n1 42.4359
R1761 VN.n42 VN.n24 42.4359
R1762 VN.n8 VN.n3 40.4934
R1763 VN.n12 VN.n3 40.4934
R1764 VN.n31 VN.n26 40.4934
R1765 VN.n35 VN.n26 40.4934
R1766 VN.n15 VN.n1 38.5509
R1767 VN.n38 VN.n24 38.5509
R1768 VN.n8 VN.n7 24.4675
R1769 VN.n13 VN.n12 24.4675
R1770 VN.n20 VN.n19 24.4675
R1771 VN.n31 VN.n30 24.4675
R1772 VN.n36 VN.n35 24.4675
R1773 VN.n43 VN.n42 24.4675
R1774 VN.n15 VN.n14 23.9782
R1775 VN.n38 VN.n37 23.9782
R1776 VN.n28 VN.n27 18.9029
R1777 VN.n5 VN.n4 18.9029
R1778 VN.n21 VN.n20 1.46852
R1779 VN.n44 VN.n43 1.46852
R1780 VN.n7 VN.n6 0.48984
R1781 VN.n14 VN.n13 0.48984
R1782 VN.n30 VN.n29 0.48984
R1783 VN.n37 VN.n36 0.48984
R1784 VN.n45 VN.n23 0.189894
R1785 VN.n41 VN.n23 0.189894
R1786 VN.n41 VN.n40 0.189894
R1787 VN.n40 VN.n39 0.189894
R1788 VN.n39 VN.n25 0.189894
R1789 VN.n34 VN.n25 0.189894
R1790 VN.n34 VN.n33 0.189894
R1791 VN.n33 VN.n32 0.189894
R1792 VN.n32 VN.n27 0.189894
R1793 VN.n9 VN.n4 0.189894
R1794 VN.n10 VN.n9 0.189894
R1795 VN.n11 VN.n10 0.189894
R1796 VN.n11 VN.n2 0.189894
R1797 VN.n16 VN.n2 0.189894
R1798 VN.n17 VN.n16 0.189894
R1799 VN.n18 VN.n17 0.189894
R1800 VN.n18 VN.n0 0.189894
R1801 VN.n22 VN.n0 0.189894
R1802 VN VN.n22 0.0516364
R1803 VDD2.n2 VDD2.n1 60.1397
R1804 VDD2.n2 VDD2.n0 60.1397
R1805 VDD2 VDD2.n5 60.1369
R1806 VDD2.n4 VDD2.n3 59.3246
R1807 VDD2.n4 VDD2.n2 46.5946
R1808 VDD2.n5 VDD2.t7 1.13517
R1809 VDD2.n5 VDD2.t0 1.13517
R1810 VDD2.n3 VDD2.t6 1.13517
R1811 VDD2.n3 VDD2.t3 1.13517
R1812 VDD2.n1 VDD2.t2 1.13517
R1813 VDD2.n1 VDD2.t1 1.13517
R1814 VDD2.n0 VDD2.t5 1.13517
R1815 VDD2.n0 VDD2.t4 1.13517
R1816 VDD2 VDD2.n4 0.929379
R1817 VTAIL.n786 VTAIL.n694 289.615
R1818 VTAIL.n94 VTAIL.n2 289.615
R1819 VTAIL.n192 VTAIL.n100 289.615
R1820 VTAIL.n292 VTAIL.n200 289.615
R1821 VTAIL.n688 VTAIL.n596 289.615
R1822 VTAIL.n588 VTAIL.n496 289.615
R1823 VTAIL.n490 VTAIL.n398 289.615
R1824 VTAIL.n390 VTAIL.n298 289.615
R1825 VTAIL.n727 VTAIL.n726 185
R1826 VTAIL.n729 VTAIL.n728 185
R1827 VTAIL.n722 VTAIL.n721 185
R1828 VTAIL.n735 VTAIL.n734 185
R1829 VTAIL.n737 VTAIL.n736 185
R1830 VTAIL.n718 VTAIL.n717 185
R1831 VTAIL.n743 VTAIL.n742 185
R1832 VTAIL.n745 VTAIL.n744 185
R1833 VTAIL.n714 VTAIL.n713 185
R1834 VTAIL.n751 VTAIL.n750 185
R1835 VTAIL.n753 VTAIL.n752 185
R1836 VTAIL.n710 VTAIL.n709 185
R1837 VTAIL.n759 VTAIL.n758 185
R1838 VTAIL.n761 VTAIL.n760 185
R1839 VTAIL.n706 VTAIL.n705 185
R1840 VTAIL.n768 VTAIL.n767 185
R1841 VTAIL.n769 VTAIL.n704 185
R1842 VTAIL.n771 VTAIL.n770 185
R1843 VTAIL.n702 VTAIL.n701 185
R1844 VTAIL.n777 VTAIL.n776 185
R1845 VTAIL.n779 VTAIL.n778 185
R1846 VTAIL.n698 VTAIL.n697 185
R1847 VTAIL.n785 VTAIL.n784 185
R1848 VTAIL.n787 VTAIL.n786 185
R1849 VTAIL.n35 VTAIL.n34 185
R1850 VTAIL.n37 VTAIL.n36 185
R1851 VTAIL.n30 VTAIL.n29 185
R1852 VTAIL.n43 VTAIL.n42 185
R1853 VTAIL.n45 VTAIL.n44 185
R1854 VTAIL.n26 VTAIL.n25 185
R1855 VTAIL.n51 VTAIL.n50 185
R1856 VTAIL.n53 VTAIL.n52 185
R1857 VTAIL.n22 VTAIL.n21 185
R1858 VTAIL.n59 VTAIL.n58 185
R1859 VTAIL.n61 VTAIL.n60 185
R1860 VTAIL.n18 VTAIL.n17 185
R1861 VTAIL.n67 VTAIL.n66 185
R1862 VTAIL.n69 VTAIL.n68 185
R1863 VTAIL.n14 VTAIL.n13 185
R1864 VTAIL.n76 VTAIL.n75 185
R1865 VTAIL.n77 VTAIL.n12 185
R1866 VTAIL.n79 VTAIL.n78 185
R1867 VTAIL.n10 VTAIL.n9 185
R1868 VTAIL.n85 VTAIL.n84 185
R1869 VTAIL.n87 VTAIL.n86 185
R1870 VTAIL.n6 VTAIL.n5 185
R1871 VTAIL.n93 VTAIL.n92 185
R1872 VTAIL.n95 VTAIL.n94 185
R1873 VTAIL.n133 VTAIL.n132 185
R1874 VTAIL.n135 VTAIL.n134 185
R1875 VTAIL.n128 VTAIL.n127 185
R1876 VTAIL.n141 VTAIL.n140 185
R1877 VTAIL.n143 VTAIL.n142 185
R1878 VTAIL.n124 VTAIL.n123 185
R1879 VTAIL.n149 VTAIL.n148 185
R1880 VTAIL.n151 VTAIL.n150 185
R1881 VTAIL.n120 VTAIL.n119 185
R1882 VTAIL.n157 VTAIL.n156 185
R1883 VTAIL.n159 VTAIL.n158 185
R1884 VTAIL.n116 VTAIL.n115 185
R1885 VTAIL.n165 VTAIL.n164 185
R1886 VTAIL.n167 VTAIL.n166 185
R1887 VTAIL.n112 VTAIL.n111 185
R1888 VTAIL.n174 VTAIL.n173 185
R1889 VTAIL.n175 VTAIL.n110 185
R1890 VTAIL.n177 VTAIL.n176 185
R1891 VTAIL.n108 VTAIL.n107 185
R1892 VTAIL.n183 VTAIL.n182 185
R1893 VTAIL.n185 VTAIL.n184 185
R1894 VTAIL.n104 VTAIL.n103 185
R1895 VTAIL.n191 VTAIL.n190 185
R1896 VTAIL.n193 VTAIL.n192 185
R1897 VTAIL.n233 VTAIL.n232 185
R1898 VTAIL.n235 VTAIL.n234 185
R1899 VTAIL.n228 VTAIL.n227 185
R1900 VTAIL.n241 VTAIL.n240 185
R1901 VTAIL.n243 VTAIL.n242 185
R1902 VTAIL.n224 VTAIL.n223 185
R1903 VTAIL.n249 VTAIL.n248 185
R1904 VTAIL.n251 VTAIL.n250 185
R1905 VTAIL.n220 VTAIL.n219 185
R1906 VTAIL.n257 VTAIL.n256 185
R1907 VTAIL.n259 VTAIL.n258 185
R1908 VTAIL.n216 VTAIL.n215 185
R1909 VTAIL.n265 VTAIL.n264 185
R1910 VTAIL.n267 VTAIL.n266 185
R1911 VTAIL.n212 VTAIL.n211 185
R1912 VTAIL.n274 VTAIL.n273 185
R1913 VTAIL.n275 VTAIL.n210 185
R1914 VTAIL.n277 VTAIL.n276 185
R1915 VTAIL.n208 VTAIL.n207 185
R1916 VTAIL.n283 VTAIL.n282 185
R1917 VTAIL.n285 VTAIL.n284 185
R1918 VTAIL.n204 VTAIL.n203 185
R1919 VTAIL.n291 VTAIL.n290 185
R1920 VTAIL.n293 VTAIL.n292 185
R1921 VTAIL.n689 VTAIL.n688 185
R1922 VTAIL.n687 VTAIL.n686 185
R1923 VTAIL.n600 VTAIL.n599 185
R1924 VTAIL.n681 VTAIL.n680 185
R1925 VTAIL.n679 VTAIL.n678 185
R1926 VTAIL.n604 VTAIL.n603 185
R1927 VTAIL.n608 VTAIL.n606 185
R1928 VTAIL.n673 VTAIL.n672 185
R1929 VTAIL.n671 VTAIL.n670 185
R1930 VTAIL.n610 VTAIL.n609 185
R1931 VTAIL.n665 VTAIL.n664 185
R1932 VTAIL.n663 VTAIL.n662 185
R1933 VTAIL.n614 VTAIL.n613 185
R1934 VTAIL.n657 VTAIL.n656 185
R1935 VTAIL.n655 VTAIL.n654 185
R1936 VTAIL.n618 VTAIL.n617 185
R1937 VTAIL.n649 VTAIL.n648 185
R1938 VTAIL.n647 VTAIL.n646 185
R1939 VTAIL.n622 VTAIL.n621 185
R1940 VTAIL.n641 VTAIL.n640 185
R1941 VTAIL.n639 VTAIL.n638 185
R1942 VTAIL.n626 VTAIL.n625 185
R1943 VTAIL.n633 VTAIL.n632 185
R1944 VTAIL.n631 VTAIL.n630 185
R1945 VTAIL.n589 VTAIL.n588 185
R1946 VTAIL.n587 VTAIL.n586 185
R1947 VTAIL.n500 VTAIL.n499 185
R1948 VTAIL.n581 VTAIL.n580 185
R1949 VTAIL.n579 VTAIL.n578 185
R1950 VTAIL.n504 VTAIL.n503 185
R1951 VTAIL.n508 VTAIL.n506 185
R1952 VTAIL.n573 VTAIL.n572 185
R1953 VTAIL.n571 VTAIL.n570 185
R1954 VTAIL.n510 VTAIL.n509 185
R1955 VTAIL.n565 VTAIL.n564 185
R1956 VTAIL.n563 VTAIL.n562 185
R1957 VTAIL.n514 VTAIL.n513 185
R1958 VTAIL.n557 VTAIL.n556 185
R1959 VTAIL.n555 VTAIL.n554 185
R1960 VTAIL.n518 VTAIL.n517 185
R1961 VTAIL.n549 VTAIL.n548 185
R1962 VTAIL.n547 VTAIL.n546 185
R1963 VTAIL.n522 VTAIL.n521 185
R1964 VTAIL.n541 VTAIL.n540 185
R1965 VTAIL.n539 VTAIL.n538 185
R1966 VTAIL.n526 VTAIL.n525 185
R1967 VTAIL.n533 VTAIL.n532 185
R1968 VTAIL.n531 VTAIL.n530 185
R1969 VTAIL.n491 VTAIL.n490 185
R1970 VTAIL.n489 VTAIL.n488 185
R1971 VTAIL.n402 VTAIL.n401 185
R1972 VTAIL.n483 VTAIL.n482 185
R1973 VTAIL.n481 VTAIL.n480 185
R1974 VTAIL.n406 VTAIL.n405 185
R1975 VTAIL.n410 VTAIL.n408 185
R1976 VTAIL.n475 VTAIL.n474 185
R1977 VTAIL.n473 VTAIL.n472 185
R1978 VTAIL.n412 VTAIL.n411 185
R1979 VTAIL.n467 VTAIL.n466 185
R1980 VTAIL.n465 VTAIL.n464 185
R1981 VTAIL.n416 VTAIL.n415 185
R1982 VTAIL.n459 VTAIL.n458 185
R1983 VTAIL.n457 VTAIL.n456 185
R1984 VTAIL.n420 VTAIL.n419 185
R1985 VTAIL.n451 VTAIL.n450 185
R1986 VTAIL.n449 VTAIL.n448 185
R1987 VTAIL.n424 VTAIL.n423 185
R1988 VTAIL.n443 VTAIL.n442 185
R1989 VTAIL.n441 VTAIL.n440 185
R1990 VTAIL.n428 VTAIL.n427 185
R1991 VTAIL.n435 VTAIL.n434 185
R1992 VTAIL.n433 VTAIL.n432 185
R1993 VTAIL.n391 VTAIL.n390 185
R1994 VTAIL.n389 VTAIL.n388 185
R1995 VTAIL.n302 VTAIL.n301 185
R1996 VTAIL.n383 VTAIL.n382 185
R1997 VTAIL.n381 VTAIL.n380 185
R1998 VTAIL.n306 VTAIL.n305 185
R1999 VTAIL.n310 VTAIL.n308 185
R2000 VTAIL.n375 VTAIL.n374 185
R2001 VTAIL.n373 VTAIL.n372 185
R2002 VTAIL.n312 VTAIL.n311 185
R2003 VTAIL.n367 VTAIL.n366 185
R2004 VTAIL.n365 VTAIL.n364 185
R2005 VTAIL.n316 VTAIL.n315 185
R2006 VTAIL.n359 VTAIL.n358 185
R2007 VTAIL.n357 VTAIL.n356 185
R2008 VTAIL.n320 VTAIL.n319 185
R2009 VTAIL.n351 VTAIL.n350 185
R2010 VTAIL.n349 VTAIL.n348 185
R2011 VTAIL.n324 VTAIL.n323 185
R2012 VTAIL.n343 VTAIL.n342 185
R2013 VTAIL.n341 VTAIL.n340 185
R2014 VTAIL.n328 VTAIL.n327 185
R2015 VTAIL.n335 VTAIL.n334 185
R2016 VTAIL.n333 VTAIL.n332 185
R2017 VTAIL.n725 VTAIL.t12 147.659
R2018 VTAIL.n33 VTAIL.t9 147.659
R2019 VTAIL.n131 VTAIL.t0 147.659
R2020 VTAIL.n231 VTAIL.t1 147.659
R2021 VTAIL.n629 VTAIL.t3 147.659
R2022 VTAIL.n529 VTAIL.t6 147.659
R2023 VTAIL.n431 VTAIL.t10 147.659
R2024 VTAIL.n331 VTAIL.t14 147.659
R2025 VTAIL.n728 VTAIL.n727 104.615
R2026 VTAIL.n728 VTAIL.n721 104.615
R2027 VTAIL.n735 VTAIL.n721 104.615
R2028 VTAIL.n736 VTAIL.n735 104.615
R2029 VTAIL.n736 VTAIL.n717 104.615
R2030 VTAIL.n743 VTAIL.n717 104.615
R2031 VTAIL.n744 VTAIL.n743 104.615
R2032 VTAIL.n744 VTAIL.n713 104.615
R2033 VTAIL.n751 VTAIL.n713 104.615
R2034 VTAIL.n752 VTAIL.n751 104.615
R2035 VTAIL.n752 VTAIL.n709 104.615
R2036 VTAIL.n759 VTAIL.n709 104.615
R2037 VTAIL.n760 VTAIL.n759 104.615
R2038 VTAIL.n760 VTAIL.n705 104.615
R2039 VTAIL.n768 VTAIL.n705 104.615
R2040 VTAIL.n769 VTAIL.n768 104.615
R2041 VTAIL.n770 VTAIL.n769 104.615
R2042 VTAIL.n770 VTAIL.n701 104.615
R2043 VTAIL.n777 VTAIL.n701 104.615
R2044 VTAIL.n778 VTAIL.n777 104.615
R2045 VTAIL.n778 VTAIL.n697 104.615
R2046 VTAIL.n785 VTAIL.n697 104.615
R2047 VTAIL.n786 VTAIL.n785 104.615
R2048 VTAIL.n36 VTAIL.n35 104.615
R2049 VTAIL.n36 VTAIL.n29 104.615
R2050 VTAIL.n43 VTAIL.n29 104.615
R2051 VTAIL.n44 VTAIL.n43 104.615
R2052 VTAIL.n44 VTAIL.n25 104.615
R2053 VTAIL.n51 VTAIL.n25 104.615
R2054 VTAIL.n52 VTAIL.n51 104.615
R2055 VTAIL.n52 VTAIL.n21 104.615
R2056 VTAIL.n59 VTAIL.n21 104.615
R2057 VTAIL.n60 VTAIL.n59 104.615
R2058 VTAIL.n60 VTAIL.n17 104.615
R2059 VTAIL.n67 VTAIL.n17 104.615
R2060 VTAIL.n68 VTAIL.n67 104.615
R2061 VTAIL.n68 VTAIL.n13 104.615
R2062 VTAIL.n76 VTAIL.n13 104.615
R2063 VTAIL.n77 VTAIL.n76 104.615
R2064 VTAIL.n78 VTAIL.n77 104.615
R2065 VTAIL.n78 VTAIL.n9 104.615
R2066 VTAIL.n85 VTAIL.n9 104.615
R2067 VTAIL.n86 VTAIL.n85 104.615
R2068 VTAIL.n86 VTAIL.n5 104.615
R2069 VTAIL.n93 VTAIL.n5 104.615
R2070 VTAIL.n94 VTAIL.n93 104.615
R2071 VTAIL.n134 VTAIL.n133 104.615
R2072 VTAIL.n134 VTAIL.n127 104.615
R2073 VTAIL.n141 VTAIL.n127 104.615
R2074 VTAIL.n142 VTAIL.n141 104.615
R2075 VTAIL.n142 VTAIL.n123 104.615
R2076 VTAIL.n149 VTAIL.n123 104.615
R2077 VTAIL.n150 VTAIL.n149 104.615
R2078 VTAIL.n150 VTAIL.n119 104.615
R2079 VTAIL.n157 VTAIL.n119 104.615
R2080 VTAIL.n158 VTAIL.n157 104.615
R2081 VTAIL.n158 VTAIL.n115 104.615
R2082 VTAIL.n165 VTAIL.n115 104.615
R2083 VTAIL.n166 VTAIL.n165 104.615
R2084 VTAIL.n166 VTAIL.n111 104.615
R2085 VTAIL.n174 VTAIL.n111 104.615
R2086 VTAIL.n175 VTAIL.n174 104.615
R2087 VTAIL.n176 VTAIL.n175 104.615
R2088 VTAIL.n176 VTAIL.n107 104.615
R2089 VTAIL.n183 VTAIL.n107 104.615
R2090 VTAIL.n184 VTAIL.n183 104.615
R2091 VTAIL.n184 VTAIL.n103 104.615
R2092 VTAIL.n191 VTAIL.n103 104.615
R2093 VTAIL.n192 VTAIL.n191 104.615
R2094 VTAIL.n234 VTAIL.n233 104.615
R2095 VTAIL.n234 VTAIL.n227 104.615
R2096 VTAIL.n241 VTAIL.n227 104.615
R2097 VTAIL.n242 VTAIL.n241 104.615
R2098 VTAIL.n242 VTAIL.n223 104.615
R2099 VTAIL.n249 VTAIL.n223 104.615
R2100 VTAIL.n250 VTAIL.n249 104.615
R2101 VTAIL.n250 VTAIL.n219 104.615
R2102 VTAIL.n257 VTAIL.n219 104.615
R2103 VTAIL.n258 VTAIL.n257 104.615
R2104 VTAIL.n258 VTAIL.n215 104.615
R2105 VTAIL.n265 VTAIL.n215 104.615
R2106 VTAIL.n266 VTAIL.n265 104.615
R2107 VTAIL.n266 VTAIL.n211 104.615
R2108 VTAIL.n274 VTAIL.n211 104.615
R2109 VTAIL.n275 VTAIL.n274 104.615
R2110 VTAIL.n276 VTAIL.n275 104.615
R2111 VTAIL.n276 VTAIL.n207 104.615
R2112 VTAIL.n283 VTAIL.n207 104.615
R2113 VTAIL.n284 VTAIL.n283 104.615
R2114 VTAIL.n284 VTAIL.n203 104.615
R2115 VTAIL.n291 VTAIL.n203 104.615
R2116 VTAIL.n292 VTAIL.n291 104.615
R2117 VTAIL.n688 VTAIL.n687 104.615
R2118 VTAIL.n687 VTAIL.n599 104.615
R2119 VTAIL.n680 VTAIL.n599 104.615
R2120 VTAIL.n680 VTAIL.n679 104.615
R2121 VTAIL.n679 VTAIL.n603 104.615
R2122 VTAIL.n608 VTAIL.n603 104.615
R2123 VTAIL.n672 VTAIL.n608 104.615
R2124 VTAIL.n672 VTAIL.n671 104.615
R2125 VTAIL.n671 VTAIL.n609 104.615
R2126 VTAIL.n664 VTAIL.n609 104.615
R2127 VTAIL.n664 VTAIL.n663 104.615
R2128 VTAIL.n663 VTAIL.n613 104.615
R2129 VTAIL.n656 VTAIL.n613 104.615
R2130 VTAIL.n656 VTAIL.n655 104.615
R2131 VTAIL.n655 VTAIL.n617 104.615
R2132 VTAIL.n648 VTAIL.n617 104.615
R2133 VTAIL.n648 VTAIL.n647 104.615
R2134 VTAIL.n647 VTAIL.n621 104.615
R2135 VTAIL.n640 VTAIL.n621 104.615
R2136 VTAIL.n640 VTAIL.n639 104.615
R2137 VTAIL.n639 VTAIL.n625 104.615
R2138 VTAIL.n632 VTAIL.n625 104.615
R2139 VTAIL.n632 VTAIL.n631 104.615
R2140 VTAIL.n588 VTAIL.n587 104.615
R2141 VTAIL.n587 VTAIL.n499 104.615
R2142 VTAIL.n580 VTAIL.n499 104.615
R2143 VTAIL.n580 VTAIL.n579 104.615
R2144 VTAIL.n579 VTAIL.n503 104.615
R2145 VTAIL.n508 VTAIL.n503 104.615
R2146 VTAIL.n572 VTAIL.n508 104.615
R2147 VTAIL.n572 VTAIL.n571 104.615
R2148 VTAIL.n571 VTAIL.n509 104.615
R2149 VTAIL.n564 VTAIL.n509 104.615
R2150 VTAIL.n564 VTAIL.n563 104.615
R2151 VTAIL.n563 VTAIL.n513 104.615
R2152 VTAIL.n556 VTAIL.n513 104.615
R2153 VTAIL.n556 VTAIL.n555 104.615
R2154 VTAIL.n555 VTAIL.n517 104.615
R2155 VTAIL.n548 VTAIL.n517 104.615
R2156 VTAIL.n548 VTAIL.n547 104.615
R2157 VTAIL.n547 VTAIL.n521 104.615
R2158 VTAIL.n540 VTAIL.n521 104.615
R2159 VTAIL.n540 VTAIL.n539 104.615
R2160 VTAIL.n539 VTAIL.n525 104.615
R2161 VTAIL.n532 VTAIL.n525 104.615
R2162 VTAIL.n532 VTAIL.n531 104.615
R2163 VTAIL.n490 VTAIL.n489 104.615
R2164 VTAIL.n489 VTAIL.n401 104.615
R2165 VTAIL.n482 VTAIL.n401 104.615
R2166 VTAIL.n482 VTAIL.n481 104.615
R2167 VTAIL.n481 VTAIL.n405 104.615
R2168 VTAIL.n410 VTAIL.n405 104.615
R2169 VTAIL.n474 VTAIL.n410 104.615
R2170 VTAIL.n474 VTAIL.n473 104.615
R2171 VTAIL.n473 VTAIL.n411 104.615
R2172 VTAIL.n466 VTAIL.n411 104.615
R2173 VTAIL.n466 VTAIL.n465 104.615
R2174 VTAIL.n465 VTAIL.n415 104.615
R2175 VTAIL.n458 VTAIL.n415 104.615
R2176 VTAIL.n458 VTAIL.n457 104.615
R2177 VTAIL.n457 VTAIL.n419 104.615
R2178 VTAIL.n450 VTAIL.n419 104.615
R2179 VTAIL.n450 VTAIL.n449 104.615
R2180 VTAIL.n449 VTAIL.n423 104.615
R2181 VTAIL.n442 VTAIL.n423 104.615
R2182 VTAIL.n442 VTAIL.n441 104.615
R2183 VTAIL.n441 VTAIL.n427 104.615
R2184 VTAIL.n434 VTAIL.n427 104.615
R2185 VTAIL.n434 VTAIL.n433 104.615
R2186 VTAIL.n390 VTAIL.n389 104.615
R2187 VTAIL.n389 VTAIL.n301 104.615
R2188 VTAIL.n382 VTAIL.n301 104.615
R2189 VTAIL.n382 VTAIL.n381 104.615
R2190 VTAIL.n381 VTAIL.n305 104.615
R2191 VTAIL.n310 VTAIL.n305 104.615
R2192 VTAIL.n374 VTAIL.n310 104.615
R2193 VTAIL.n374 VTAIL.n373 104.615
R2194 VTAIL.n373 VTAIL.n311 104.615
R2195 VTAIL.n366 VTAIL.n311 104.615
R2196 VTAIL.n366 VTAIL.n365 104.615
R2197 VTAIL.n365 VTAIL.n315 104.615
R2198 VTAIL.n358 VTAIL.n315 104.615
R2199 VTAIL.n358 VTAIL.n357 104.615
R2200 VTAIL.n357 VTAIL.n319 104.615
R2201 VTAIL.n350 VTAIL.n319 104.615
R2202 VTAIL.n350 VTAIL.n349 104.615
R2203 VTAIL.n349 VTAIL.n323 104.615
R2204 VTAIL.n342 VTAIL.n323 104.615
R2205 VTAIL.n342 VTAIL.n341 104.615
R2206 VTAIL.n341 VTAIL.n327 104.615
R2207 VTAIL.n334 VTAIL.n327 104.615
R2208 VTAIL.n334 VTAIL.n333 104.615
R2209 VTAIL.n727 VTAIL.t12 52.3082
R2210 VTAIL.n35 VTAIL.t9 52.3082
R2211 VTAIL.n133 VTAIL.t0 52.3082
R2212 VTAIL.n233 VTAIL.t1 52.3082
R2213 VTAIL.n631 VTAIL.t3 52.3082
R2214 VTAIL.n531 VTAIL.t6 52.3082
R2215 VTAIL.n433 VTAIL.t10 52.3082
R2216 VTAIL.n333 VTAIL.t14 52.3082
R2217 VTAIL.n595 VTAIL.n594 42.6458
R2218 VTAIL.n397 VTAIL.n396 42.6458
R2219 VTAIL.n1 VTAIL.n0 42.6456
R2220 VTAIL.n199 VTAIL.n198 42.6456
R2221 VTAIL.n791 VTAIL.n790 30.8278
R2222 VTAIL.n99 VTAIL.n98 30.8278
R2223 VTAIL.n197 VTAIL.n196 30.8278
R2224 VTAIL.n297 VTAIL.n296 30.8278
R2225 VTAIL.n693 VTAIL.n692 30.8278
R2226 VTAIL.n593 VTAIL.n592 30.8278
R2227 VTAIL.n495 VTAIL.n494 30.8278
R2228 VTAIL.n395 VTAIL.n394 30.8278
R2229 VTAIL.n791 VTAIL.n693 29.1514
R2230 VTAIL.n395 VTAIL.n297 29.1514
R2231 VTAIL.n726 VTAIL.n725 15.6677
R2232 VTAIL.n34 VTAIL.n33 15.6677
R2233 VTAIL.n132 VTAIL.n131 15.6677
R2234 VTAIL.n232 VTAIL.n231 15.6677
R2235 VTAIL.n630 VTAIL.n629 15.6677
R2236 VTAIL.n530 VTAIL.n529 15.6677
R2237 VTAIL.n432 VTAIL.n431 15.6677
R2238 VTAIL.n332 VTAIL.n331 15.6677
R2239 VTAIL.n771 VTAIL.n702 13.1884
R2240 VTAIL.n79 VTAIL.n10 13.1884
R2241 VTAIL.n177 VTAIL.n108 13.1884
R2242 VTAIL.n277 VTAIL.n208 13.1884
R2243 VTAIL.n606 VTAIL.n604 13.1884
R2244 VTAIL.n506 VTAIL.n504 13.1884
R2245 VTAIL.n408 VTAIL.n406 13.1884
R2246 VTAIL.n308 VTAIL.n306 13.1884
R2247 VTAIL.n729 VTAIL.n724 12.8005
R2248 VTAIL.n772 VTAIL.n704 12.8005
R2249 VTAIL.n776 VTAIL.n775 12.8005
R2250 VTAIL.n37 VTAIL.n32 12.8005
R2251 VTAIL.n80 VTAIL.n12 12.8005
R2252 VTAIL.n84 VTAIL.n83 12.8005
R2253 VTAIL.n135 VTAIL.n130 12.8005
R2254 VTAIL.n178 VTAIL.n110 12.8005
R2255 VTAIL.n182 VTAIL.n181 12.8005
R2256 VTAIL.n235 VTAIL.n230 12.8005
R2257 VTAIL.n278 VTAIL.n210 12.8005
R2258 VTAIL.n282 VTAIL.n281 12.8005
R2259 VTAIL.n678 VTAIL.n677 12.8005
R2260 VTAIL.n674 VTAIL.n673 12.8005
R2261 VTAIL.n633 VTAIL.n628 12.8005
R2262 VTAIL.n578 VTAIL.n577 12.8005
R2263 VTAIL.n574 VTAIL.n573 12.8005
R2264 VTAIL.n533 VTAIL.n528 12.8005
R2265 VTAIL.n480 VTAIL.n479 12.8005
R2266 VTAIL.n476 VTAIL.n475 12.8005
R2267 VTAIL.n435 VTAIL.n430 12.8005
R2268 VTAIL.n380 VTAIL.n379 12.8005
R2269 VTAIL.n376 VTAIL.n375 12.8005
R2270 VTAIL.n335 VTAIL.n330 12.8005
R2271 VTAIL.n730 VTAIL.n722 12.0247
R2272 VTAIL.n767 VTAIL.n766 12.0247
R2273 VTAIL.n779 VTAIL.n700 12.0247
R2274 VTAIL.n38 VTAIL.n30 12.0247
R2275 VTAIL.n75 VTAIL.n74 12.0247
R2276 VTAIL.n87 VTAIL.n8 12.0247
R2277 VTAIL.n136 VTAIL.n128 12.0247
R2278 VTAIL.n173 VTAIL.n172 12.0247
R2279 VTAIL.n185 VTAIL.n106 12.0247
R2280 VTAIL.n236 VTAIL.n228 12.0247
R2281 VTAIL.n273 VTAIL.n272 12.0247
R2282 VTAIL.n285 VTAIL.n206 12.0247
R2283 VTAIL.n681 VTAIL.n602 12.0247
R2284 VTAIL.n670 VTAIL.n607 12.0247
R2285 VTAIL.n634 VTAIL.n626 12.0247
R2286 VTAIL.n581 VTAIL.n502 12.0247
R2287 VTAIL.n570 VTAIL.n507 12.0247
R2288 VTAIL.n534 VTAIL.n526 12.0247
R2289 VTAIL.n483 VTAIL.n404 12.0247
R2290 VTAIL.n472 VTAIL.n409 12.0247
R2291 VTAIL.n436 VTAIL.n428 12.0247
R2292 VTAIL.n383 VTAIL.n304 12.0247
R2293 VTAIL.n372 VTAIL.n309 12.0247
R2294 VTAIL.n336 VTAIL.n328 12.0247
R2295 VTAIL.n734 VTAIL.n733 11.249
R2296 VTAIL.n765 VTAIL.n706 11.249
R2297 VTAIL.n780 VTAIL.n698 11.249
R2298 VTAIL.n42 VTAIL.n41 11.249
R2299 VTAIL.n73 VTAIL.n14 11.249
R2300 VTAIL.n88 VTAIL.n6 11.249
R2301 VTAIL.n140 VTAIL.n139 11.249
R2302 VTAIL.n171 VTAIL.n112 11.249
R2303 VTAIL.n186 VTAIL.n104 11.249
R2304 VTAIL.n240 VTAIL.n239 11.249
R2305 VTAIL.n271 VTAIL.n212 11.249
R2306 VTAIL.n286 VTAIL.n204 11.249
R2307 VTAIL.n682 VTAIL.n600 11.249
R2308 VTAIL.n669 VTAIL.n610 11.249
R2309 VTAIL.n638 VTAIL.n637 11.249
R2310 VTAIL.n582 VTAIL.n500 11.249
R2311 VTAIL.n569 VTAIL.n510 11.249
R2312 VTAIL.n538 VTAIL.n537 11.249
R2313 VTAIL.n484 VTAIL.n402 11.249
R2314 VTAIL.n471 VTAIL.n412 11.249
R2315 VTAIL.n440 VTAIL.n439 11.249
R2316 VTAIL.n384 VTAIL.n302 11.249
R2317 VTAIL.n371 VTAIL.n312 11.249
R2318 VTAIL.n340 VTAIL.n339 11.249
R2319 VTAIL.n737 VTAIL.n720 10.4732
R2320 VTAIL.n762 VTAIL.n761 10.4732
R2321 VTAIL.n784 VTAIL.n783 10.4732
R2322 VTAIL.n45 VTAIL.n28 10.4732
R2323 VTAIL.n70 VTAIL.n69 10.4732
R2324 VTAIL.n92 VTAIL.n91 10.4732
R2325 VTAIL.n143 VTAIL.n126 10.4732
R2326 VTAIL.n168 VTAIL.n167 10.4732
R2327 VTAIL.n190 VTAIL.n189 10.4732
R2328 VTAIL.n243 VTAIL.n226 10.4732
R2329 VTAIL.n268 VTAIL.n267 10.4732
R2330 VTAIL.n290 VTAIL.n289 10.4732
R2331 VTAIL.n686 VTAIL.n685 10.4732
R2332 VTAIL.n666 VTAIL.n665 10.4732
R2333 VTAIL.n641 VTAIL.n624 10.4732
R2334 VTAIL.n586 VTAIL.n585 10.4732
R2335 VTAIL.n566 VTAIL.n565 10.4732
R2336 VTAIL.n541 VTAIL.n524 10.4732
R2337 VTAIL.n488 VTAIL.n487 10.4732
R2338 VTAIL.n468 VTAIL.n467 10.4732
R2339 VTAIL.n443 VTAIL.n426 10.4732
R2340 VTAIL.n388 VTAIL.n387 10.4732
R2341 VTAIL.n368 VTAIL.n367 10.4732
R2342 VTAIL.n343 VTAIL.n326 10.4732
R2343 VTAIL.n738 VTAIL.n718 9.69747
R2344 VTAIL.n758 VTAIL.n708 9.69747
R2345 VTAIL.n787 VTAIL.n696 9.69747
R2346 VTAIL.n46 VTAIL.n26 9.69747
R2347 VTAIL.n66 VTAIL.n16 9.69747
R2348 VTAIL.n95 VTAIL.n4 9.69747
R2349 VTAIL.n144 VTAIL.n124 9.69747
R2350 VTAIL.n164 VTAIL.n114 9.69747
R2351 VTAIL.n193 VTAIL.n102 9.69747
R2352 VTAIL.n244 VTAIL.n224 9.69747
R2353 VTAIL.n264 VTAIL.n214 9.69747
R2354 VTAIL.n293 VTAIL.n202 9.69747
R2355 VTAIL.n689 VTAIL.n598 9.69747
R2356 VTAIL.n662 VTAIL.n612 9.69747
R2357 VTAIL.n642 VTAIL.n622 9.69747
R2358 VTAIL.n589 VTAIL.n498 9.69747
R2359 VTAIL.n562 VTAIL.n512 9.69747
R2360 VTAIL.n542 VTAIL.n522 9.69747
R2361 VTAIL.n491 VTAIL.n400 9.69747
R2362 VTAIL.n464 VTAIL.n414 9.69747
R2363 VTAIL.n444 VTAIL.n424 9.69747
R2364 VTAIL.n391 VTAIL.n300 9.69747
R2365 VTAIL.n364 VTAIL.n314 9.69747
R2366 VTAIL.n344 VTAIL.n324 9.69747
R2367 VTAIL.n790 VTAIL.n789 9.45567
R2368 VTAIL.n98 VTAIL.n97 9.45567
R2369 VTAIL.n196 VTAIL.n195 9.45567
R2370 VTAIL.n296 VTAIL.n295 9.45567
R2371 VTAIL.n692 VTAIL.n691 9.45567
R2372 VTAIL.n592 VTAIL.n591 9.45567
R2373 VTAIL.n494 VTAIL.n493 9.45567
R2374 VTAIL.n394 VTAIL.n393 9.45567
R2375 VTAIL.n789 VTAIL.n788 9.3005
R2376 VTAIL.n696 VTAIL.n695 9.3005
R2377 VTAIL.n783 VTAIL.n782 9.3005
R2378 VTAIL.n781 VTAIL.n780 9.3005
R2379 VTAIL.n700 VTAIL.n699 9.3005
R2380 VTAIL.n775 VTAIL.n774 9.3005
R2381 VTAIL.n747 VTAIL.n746 9.3005
R2382 VTAIL.n716 VTAIL.n715 9.3005
R2383 VTAIL.n741 VTAIL.n740 9.3005
R2384 VTAIL.n739 VTAIL.n738 9.3005
R2385 VTAIL.n720 VTAIL.n719 9.3005
R2386 VTAIL.n733 VTAIL.n732 9.3005
R2387 VTAIL.n731 VTAIL.n730 9.3005
R2388 VTAIL.n724 VTAIL.n723 9.3005
R2389 VTAIL.n749 VTAIL.n748 9.3005
R2390 VTAIL.n712 VTAIL.n711 9.3005
R2391 VTAIL.n755 VTAIL.n754 9.3005
R2392 VTAIL.n757 VTAIL.n756 9.3005
R2393 VTAIL.n708 VTAIL.n707 9.3005
R2394 VTAIL.n763 VTAIL.n762 9.3005
R2395 VTAIL.n765 VTAIL.n764 9.3005
R2396 VTAIL.n766 VTAIL.n703 9.3005
R2397 VTAIL.n773 VTAIL.n772 9.3005
R2398 VTAIL.n97 VTAIL.n96 9.3005
R2399 VTAIL.n4 VTAIL.n3 9.3005
R2400 VTAIL.n91 VTAIL.n90 9.3005
R2401 VTAIL.n89 VTAIL.n88 9.3005
R2402 VTAIL.n8 VTAIL.n7 9.3005
R2403 VTAIL.n83 VTAIL.n82 9.3005
R2404 VTAIL.n55 VTAIL.n54 9.3005
R2405 VTAIL.n24 VTAIL.n23 9.3005
R2406 VTAIL.n49 VTAIL.n48 9.3005
R2407 VTAIL.n47 VTAIL.n46 9.3005
R2408 VTAIL.n28 VTAIL.n27 9.3005
R2409 VTAIL.n41 VTAIL.n40 9.3005
R2410 VTAIL.n39 VTAIL.n38 9.3005
R2411 VTAIL.n32 VTAIL.n31 9.3005
R2412 VTAIL.n57 VTAIL.n56 9.3005
R2413 VTAIL.n20 VTAIL.n19 9.3005
R2414 VTAIL.n63 VTAIL.n62 9.3005
R2415 VTAIL.n65 VTAIL.n64 9.3005
R2416 VTAIL.n16 VTAIL.n15 9.3005
R2417 VTAIL.n71 VTAIL.n70 9.3005
R2418 VTAIL.n73 VTAIL.n72 9.3005
R2419 VTAIL.n74 VTAIL.n11 9.3005
R2420 VTAIL.n81 VTAIL.n80 9.3005
R2421 VTAIL.n195 VTAIL.n194 9.3005
R2422 VTAIL.n102 VTAIL.n101 9.3005
R2423 VTAIL.n189 VTAIL.n188 9.3005
R2424 VTAIL.n187 VTAIL.n186 9.3005
R2425 VTAIL.n106 VTAIL.n105 9.3005
R2426 VTAIL.n181 VTAIL.n180 9.3005
R2427 VTAIL.n153 VTAIL.n152 9.3005
R2428 VTAIL.n122 VTAIL.n121 9.3005
R2429 VTAIL.n147 VTAIL.n146 9.3005
R2430 VTAIL.n145 VTAIL.n144 9.3005
R2431 VTAIL.n126 VTAIL.n125 9.3005
R2432 VTAIL.n139 VTAIL.n138 9.3005
R2433 VTAIL.n137 VTAIL.n136 9.3005
R2434 VTAIL.n130 VTAIL.n129 9.3005
R2435 VTAIL.n155 VTAIL.n154 9.3005
R2436 VTAIL.n118 VTAIL.n117 9.3005
R2437 VTAIL.n161 VTAIL.n160 9.3005
R2438 VTAIL.n163 VTAIL.n162 9.3005
R2439 VTAIL.n114 VTAIL.n113 9.3005
R2440 VTAIL.n169 VTAIL.n168 9.3005
R2441 VTAIL.n171 VTAIL.n170 9.3005
R2442 VTAIL.n172 VTAIL.n109 9.3005
R2443 VTAIL.n179 VTAIL.n178 9.3005
R2444 VTAIL.n295 VTAIL.n294 9.3005
R2445 VTAIL.n202 VTAIL.n201 9.3005
R2446 VTAIL.n289 VTAIL.n288 9.3005
R2447 VTAIL.n287 VTAIL.n286 9.3005
R2448 VTAIL.n206 VTAIL.n205 9.3005
R2449 VTAIL.n281 VTAIL.n280 9.3005
R2450 VTAIL.n253 VTAIL.n252 9.3005
R2451 VTAIL.n222 VTAIL.n221 9.3005
R2452 VTAIL.n247 VTAIL.n246 9.3005
R2453 VTAIL.n245 VTAIL.n244 9.3005
R2454 VTAIL.n226 VTAIL.n225 9.3005
R2455 VTAIL.n239 VTAIL.n238 9.3005
R2456 VTAIL.n237 VTAIL.n236 9.3005
R2457 VTAIL.n230 VTAIL.n229 9.3005
R2458 VTAIL.n255 VTAIL.n254 9.3005
R2459 VTAIL.n218 VTAIL.n217 9.3005
R2460 VTAIL.n261 VTAIL.n260 9.3005
R2461 VTAIL.n263 VTAIL.n262 9.3005
R2462 VTAIL.n214 VTAIL.n213 9.3005
R2463 VTAIL.n269 VTAIL.n268 9.3005
R2464 VTAIL.n271 VTAIL.n270 9.3005
R2465 VTAIL.n272 VTAIL.n209 9.3005
R2466 VTAIL.n279 VTAIL.n278 9.3005
R2467 VTAIL.n616 VTAIL.n615 9.3005
R2468 VTAIL.n659 VTAIL.n658 9.3005
R2469 VTAIL.n661 VTAIL.n660 9.3005
R2470 VTAIL.n612 VTAIL.n611 9.3005
R2471 VTAIL.n667 VTAIL.n666 9.3005
R2472 VTAIL.n669 VTAIL.n668 9.3005
R2473 VTAIL.n607 VTAIL.n605 9.3005
R2474 VTAIL.n675 VTAIL.n674 9.3005
R2475 VTAIL.n691 VTAIL.n690 9.3005
R2476 VTAIL.n598 VTAIL.n597 9.3005
R2477 VTAIL.n685 VTAIL.n684 9.3005
R2478 VTAIL.n683 VTAIL.n682 9.3005
R2479 VTAIL.n602 VTAIL.n601 9.3005
R2480 VTAIL.n677 VTAIL.n676 9.3005
R2481 VTAIL.n653 VTAIL.n652 9.3005
R2482 VTAIL.n651 VTAIL.n650 9.3005
R2483 VTAIL.n620 VTAIL.n619 9.3005
R2484 VTAIL.n645 VTAIL.n644 9.3005
R2485 VTAIL.n643 VTAIL.n642 9.3005
R2486 VTAIL.n624 VTAIL.n623 9.3005
R2487 VTAIL.n637 VTAIL.n636 9.3005
R2488 VTAIL.n635 VTAIL.n634 9.3005
R2489 VTAIL.n628 VTAIL.n627 9.3005
R2490 VTAIL.n516 VTAIL.n515 9.3005
R2491 VTAIL.n559 VTAIL.n558 9.3005
R2492 VTAIL.n561 VTAIL.n560 9.3005
R2493 VTAIL.n512 VTAIL.n511 9.3005
R2494 VTAIL.n567 VTAIL.n566 9.3005
R2495 VTAIL.n569 VTAIL.n568 9.3005
R2496 VTAIL.n507 VTAIL.n505 9.3005
R2497 VTAIL.n575 VTAIL.n574 9.3005
R2498 VTAIL.n591 VTAIL.n590 9.3005
R2499 VTAIL.n498 VTAIL.n497 9.3005
R2500 VTAIL.n585 VTAIL.n584 9.3005
R2501 VTAIL.n583 VTAIL.n582 9.3005
R2502 VTAIL.n502 VTAIL.n501 9.3005
R2503 VTAIL.n577 VTAIL.n576 9.3005
R2504 VTAIL.n553 VTAIL.n552 9.3005
R2505 VTAIL.n551 VTAIL.n550 9.3005
R2506 VTAIL.n520 VTAIL.n519 9.3005
R2507 VTAIL.n545 VTAIL.n544 9.3005
R2508 VTAIL.n543 VTAIL.n542 9.3005
R2509 VTAIL.n524 VTAIL.n523 9.3005
R2510 VTAIL.n537 VTAIL.n536 9.3005
R2511 VTAIL.n535 VTAIL.n534 9.3005
R2512 VTAIL.n528 VTAIL.n527 9.3005
R2513 VTAIL.n418 VTAIL.n417 9.3005
R2514 VTAIL.n461 VTAIL.n460 9.3005
R2515 VTAIL.n463 VTAIL.n462 9.3005
R2516 VTAIL.n414 VTAIL.n413 9.3005
R2517 VTAIL.n469 VTAIL.n468 9.3005
R2518 VTAIL.n471 VTAIL.n470 9.3005
R2519 VTAIL.n409 VTAIL.n407 9.3005
R2520 VTAIL.n477 VTAIL.n476 9.3005
R2521 VTAIL.n493 VTAIL.n492 9.3005
R2522 VTAIL.n400 VTAIL.n399 9.3005
R2523 VTAIL.n487 VTAIL.n486 9.3005
R2524 VTAIL.n485 VTAIL.n484 9.3005
R2525 VTAIL.n404 VTAIL.n403 9.3005
R2526 VTAIL.n479 VTAIL.n478 9.3005
R2527 VTAIL.n455 VTAIL.n454 9.3005
R2528 VTAIL.n453 VTAIL.n452 9.3005
R2529 VTAIL.n422 VTAIL.n421 9.3005
R2530 VTAIL.n447 VTAIL.n446 9.3005
R2531 VTAIL.n445 VTAIL.n444 9.3005
R2532 VTAIL.n426 VTAIL.n425 9.3005
R2533 VTAIL.n439 VTAIL.n438 9.3005
R2534 VTAIL.n437 VTAIL.n436 9.3005
R2535 VTAIL.n430 VTAIL.n429 9.3005
R2536 VTAIL.n318 VTAIL.n317 9.3005
R2537 VTAIL.n361 VTAIL.n360 9.3005
R2538 VTAIL.n363 VTAIL.n362 9.3005
R2539 VTAIL.n314 VTAIL.n313 9.3005
R2540 VTAIL.n369 VTAIL.n368 9.3005
R2541 VTAIL.n371 VTAIL.n370 9.3005
R2542 VTAIL.n309 VTAIL.n307 9.3005
R2543 VTAIL.n377 VTAIL.n376 9.3005
R2544 VTAIL.n393 VTAIL.n392 9.3005
R2545 VTAIL.n300 VTAIL.n299 9.3005
R2546 VTAIL.n387 VTAIL.n386 9.3005
R2547 VTAIL.n385 VTAIL.n384 9.3005
R2548 VTAIL.n304 VTAIL.n303 9.3005
R2549 VTAIL.n379 VTAIL.n378 9.3005
R2550 VTAIL.n355 VTAIL.n354 9.3005
R2551 VTAIL.n353 VTAIL.n352 9.3005
R2552 VTAIL.n322 VTAIL.n321 9.3005
R2553 VTAIL.n347 VTAIL.n346 9.3005
R2554 VTAIL.n345 VTAIL.n344 9.3005
R2555 VTAIL.n326 VTAIL.n325 9.3005
R2556 VTAIL.n339 VTAIL.n338 9.3005
R2557 VTAIL.n337 VTAIL.n336 9.3005
R2558 VTAIL.n330 VTAIL.n329 9.3005
R2559 VTAIL.n742 VTAIL.n741 8.92171
R2560 VTAIL.n757 VTAIL.n710 8.92171
R2561 VTAIL.n788 VTAIL.n694 8.92171
R2562 VTAIL.n50 VTAIL.n49 8.92171
R2563 VTAIL.n65 VTAIL.n18 8.92171
R2564 VTAIL.n96 VTAIL.n2 8.92171
R2565 VTAIL.n148 VTAIL.n147 8.92171
R2566 VTAIL.n163 VTAIL.n116 8.92171
R2567 VTAIL.n194 VTAIL.n100 8.92171
R2568 VTAIL.n248 VTAIL.n247 8.92171
R2569 VTAIL.n263 VTAIL.n216 8.92171
R2570 VTAIL.n294 VTAIL.n200 8.92171
R2571 VTAIL.n690 VTAIL.n596 8.92171
R2572 VTAIL.n661 VTAIL.n614 8.92171
R2573 VTAIL.n646 VTAIL.n645 8.92171
R2574 VTAIL.n590 VTAIL.n496 8.92171
R2575 VTAIL.n561 VTAIL.n514 8.92171
R2576 VTAIL.n546 VTAIL.n545 8.92171
R2577 VTAIL.n492 VTAIL.n398 8.92171
R2578 VTAIL.n463 VTAIL.n416 8.92171
R2579 VTAIL.n448 VTAIL.n447 8.92171
R2580 VTAIL.n392 VTAIL.n298 8.92171
R2581 VTAIL.n363 VTAIL.n316 8.92171
R2582 VTAIL.n348 VTAIL.n347 8.92171
R2583 VTAIL.n745 VTAIL.n716 8.14595
R2584 VTAIL.n754 VTAIL.n753 8.14595
R2585 VTAIL.n53 VTAIL.n24 8.14595
R2586 VTAIL.n62 VTAIL.n61 8.14595
R2587 VTAIL.n151 VTAIL.n122 8.14595
R2588 VTAIL.n160 VTAIL.n159 8.14595
R2589 VTAIL.n251 VTAIL.n222 8.14595
R2590 VTAIL.n260 VTAIL.n259 8.14595
R2591 VTAIL.n658 VTAIL.n657 8.14595
R2592 VTAIL.n649 VTAIL.n620 8.14595
R2593 VTAIL.n558 VTAIL.n557 8.14595
R2594 VTAIL.n549 VTAIL.n520 8.14595
R2595 VTAIL.n460 VTAIL.n459 8.14595
R2596 VTAIL.n451 VTAIL.n422 8.14595
R2597 VTAIL.n360 VTAIL.n359 8.14595
R2598 VTAIL.n351 VTAIL.n322 8.14595
R2599 VTAIL.n746 VTAIL.n714 7.3702
R2600 VTAIL.n750 VTAIL.n712 7.3702
R2601 VTAIL.n54 VTAIL.n22 7.3702
R2602 VTAIL.n58 VTAIL.n20 7.3702
R2603 VTAIL.n152 VTAIL.n120 7.3702
R2604 VTAIL.n156 VTAIL.n118 7.3702
R2605 VTAIL.n252 VTAIL.n220 7.3702
R2606 VTAIL.n256 VTAIL.n218 7.3702
R2607 VTAIL.n654 VTAIL.n616 7.3702
R2608 VTAIL.n650 VTAIL.n618 7.3702
R2609 VTAIL.n554 VTAIL.n516 7.3702
R2610 VTAIL.n550 VTAIL.n518 7.3702
R2611 VTAIL.n456 VTAIL.n418 7.3702
R2612 VTAIL.n452 VTAIL.n420 7.3702
R2613 VTAIL.n356 VTAIL.n318 7.3702
R2614 VTAIL.n352 VTAIL.n320 7.3702
R2615 VTAIL.n749 VTAIL.n714 6.59444
R2616 VTAIL.n750 VTAIL.n749 6.59444
R2617 VTAIL.n57 VTAIL.n22 6.59444
R2618 VTAIL.n58 VTAIL.n57 6.59444
R2619 VTAIL.n155 VTAIL.n120 6.59444
R2620 VTAIL.n156 VTAIL.n155 6.59444
R2621 VTAIL.n255 VTAIL.n220 6.59444
R2622 VTAIL.n256 VTAIL.n255 6.59444
R2623 VTAIL.n654 VTAIL.n653 6.59444
R2624 VTAIL.n653 VTAIL.n618 6.59444
R2625 VTAIL.n554 VTAIL.n553 6.59444
R2626 VTAIL.n553 VTAIL.n518 6.59444
R2627 VTAIL.n456 VTAIL.n455 6.59444
R2628 VTAIL.n455 VTAIL.n420 6.59444
R2629 VTAIL.n356 VTAIL.n355 6.59444
R2630 VTAIL.n355 VTAIL.n320 6.59444
R2631 VTAIL.n746 VTAIL.n745 5.81868
R2632 VTAIL.n753 VTAIL.n712 5.81868
R2633 VTAIL.n54 VTAIL.n53 5.81868
R2634 VTAIL.n61 VTAIL.n20 5.81868
R2635 VTAIL.n152 VTAIL.n151 5.81868
R2636 VTAIL.n159 VTAIL.n118 5.81868
R2637 VTAIL.n252 VTAIL.n251 5.81868
R2638 VTAIL.n259 VTAIL.n218 5.81868
R2639 VTAIL.n657 VTAIL.n616 5.81868
R2640 VTAIL.n650 VTAIL.n649 5.81868
R2641 VTAIL.n557 VTAIL.n516 5.81868
R2642 VTAIL.n550 VTAIL.n549 5.81868
R2643 VTAIL.n459 VTAIL.n418 5.81868
R2644 VTAIL.n452 VTAIL.n451 5.81868
R2645 VTAIL.n359 VTAIL.n318 5.81868
R2646 VTAIL.n352 VTAIL.n351 5.81868
R2647 VTAIL.n742 VTAIL.n716 5.04292
R2648 VTAIL.n754 VTAIL.n710 5.04292
R2649 VTAIL.n790 VTAIL.n694 5.04292
R2650 VTAIL.n50 VTAIL.n24 5.04292
R2651 VTAIL.n62 VTAIL.n18 5.04292
R2652 VTAIL.n98 VTAIL.n2 5.04292
R2653 VTAIL.n148 VTAIL.n122 5.04292
R2654 VTAIL.n160 VTAIL.n116 5.04292
R2655 VTAIL.n196 VTAIL.n100 5.04292
R2656 VTAIL.n248 VTAIL.n222 5.04292
R2657 VTAIL.n260 VTAIL.n216 5.04292
R2658 VTAIL.n296 VTAIL.n200 5.04292
R2659 VTAIL.n692 VTAIL.n596 5.04292
R2660 VTAIL.n658 VTAIL.n614 5.04292
R2661 VTAIL.n646 VTAIL.n620 5.04292
R2662 VTAIL.n592 VTAIL.n496 5.04292
R2663 VTAIL.n558 VTAIL.n514 5.04292
R2664 VTAIL.n546 VTAIL.n520 5.04292
R2665 VTAIL.n494 VTAIL.n398 5.04292
R2666 VTAIL.n460 VTAIL.n416 5.04292
R2667 VTAIL.n448 VTAIL.n422 5.04292
R2668 VTAIL.n394 VTAIL.n298 5.04292
R2669 VTAIL.n360 VTAIL.n316 5.04292
R2670 VTAIL.n348 VTAIL.n322 5.04292
R2671 VTAIL.n725 VTAIL.n723 4.38563
R2672 VTAIL.n33 VTAIL.n31 4.38563
R2673 VTAIL.n131 VTAIL.n129 4.38563
R2674 VTAIL.n231 VTAIL.n229 4.38563
R2675 VTAIL.n629 VTAIL.n627 4.38563
R2676 VTAIL.n529 VTAIL.n527 4.38563
R2677 VTAIL.n431 VTAIL.n429 4.38563
R2678 VTAIL.n331 VTAIL.n329 4.38563
R2679 VTAIL.n741 VTAIL.n718 4.26717
R2680 VTAIL.n758 VTAIL.n757 4.26717
R2681 VTAIL.n788 VTAIL.n787 4.26717
R2682 VTAIL.n49 VTAIL.n26 4.26717
R2683 VTAIL.n66 VTAIL.n65 4.26717
R2684 VTAIL.n96 VTAIL.n95 4.26717
R2685 VTAIL.n147 VTAIL.n124 4.26717
R2686 VTAIL.n164 VTAIL.n163 4.26717
R2687 VTAIL.n194 VTAIL.n193 4.26717
R2688 VTAIL.n247 VTAIL.n224 4.26717
R2689 VTAIL.n264 VTAIL.n263 4.26717
R2690 VTAIL.n294 VTAIL.n293 4.26717
R2691 VTAIL.n690 VTAIL.n689 4.26717
R2692 VTAIL.n662 VTAIL.n661 4.26717
R2693 VTAIL.n645 VTAIL.n622 4.26717
R2694 VTAIL.n590 VTAIL.n589 4.26717
R2695 VTAIL.n562 VTAIL.n561 4.26717
R2696 VTAIL.n545 VTAIL.n522 4.26717
R2697 VTAIL.n492 VTAIL.n491 4.26717
R2698 VTAIL.n464 VTAIL.n463 4.26717
R2699 VTAIL.n447 VTAIL.n424 4.26717
R2700 VTAIL.n392 VTAIL.n391 4.26717
R2701 VTAIL.n364 VTAIL.n363 4.26717
R2702 VTAIL.n347 VTAIL.n324 4.26717
R2703 VTAIL.n738 VTAIL.n737 3.49141
R2704 VTAIL.n761 VTAIL.n708 3.49141
R2705 VTAIL.n784 VTAIL.n696 3.49141
R2706 VTAIL.n46 VTAIL.n45 3.49141
R2707 VTAIL.n69 VTAIL.n16 3.49141
R2708 VTAIL.n92 VTAIL.n4 3.49141
R2709 VTAIL.n144 VTAIL.n143 3.49141
R2710 VTAIL.n167 VTAIL.n114 3.49141
R2711 VTAIL.n190 VTAIL.n102 3.49141
R2712 VTAIL.n244 VTAIL.n243 3.49141
R2713 VTAIL.n267 VTAIL.n214 3.49141
R2714 VTAIL.n290 VTAIL.n202 3.49141
R2715 VTAIL.n686 VTAIL.n598 3.49141
R2716 VTAIL.n665 VTAIL.n612 3.49141
R2717 VTAIL.n642 VTAIL.n641 3.49141
R2718 VTAIL.n586 VTAIL.n498 3.49141
R2719 VTAIL.n565 VTAIL.n512 3.49141
R2720 VTAIL.n542 VTAIL.n541 3.49141
R2721 VTAIL.n488 VTAIL.n400 3.49141
R2722 VTAIL.n467 VTAIL.n414 3.49141
R2723 VTAIL.n444 VTAIL.n443 3.49141
R2724 VTAIL.n388 VTAIL.n300 3.49141
R2725 VTAIL.n367 VTAIL.n314 3.49141
R2726 VTAIL.n344 VTAIL.n343 3.49141
R2727 VTAIL.n734 VTAIL.n720 2.71565
R2728 VTAIL.n762 VTAIL.n706 2.71565
R2729 VTAIL.n783 VTAIL.n698 2.71565
R2730 VTAIL.n42 VTAIL.n28 2.71565
R2731 VTAIL.n70 VTAIL.n14 2.71565
R2732 VTAIL.n91 VTAIL.n6 2.71565
R2733 VTAIL.n140 VTAIL.n126 2.71565
R2734 VTAIL.n168 VTAIL.n112 2.71565
R2735 VTAIL.n189 VTAIL.n104 2.71565
R2736 VTAIL.n240 VTAIL.n226 2.71565
R2737 VTAIL.n268 VTAIL.n212 2.71565
R2738 VTAIL.n289 VTAIL.n204 2.71565
R2739 VTAIL.n685 VTAIL.n600 2.71565
R2740 VTAIL.n666 VTAIL.n610 2.71565
R2741 VTAIL.n638 VTAIL.n624 2.71565
R2742 VTAIL.n585 VTAIL.n500 2.71565
R2743 VTAIL.n566 VTAIL.n510 2.71565
R2744 VTAIL.n538 VTAIL.n524 2.71565
R2745 VTAIL.n487 VTAIL.n402 2.71565
R2746 VTAIL.n468 VTAIL.n412 2.71565
R2747 VTAIL.n440 VTAIL.n426 2.71565
R2748 VTAIL.n387 VTAIL.n302 2.71565
R2749 VTAIL.n368 VTAIL.n312 2.71565
R2750 VTAIL.n340 VTAIL.n326 2.71565
R2751 VTAIL.n733 VTAIL.n722 1.93989
R2752 VTAIL.n767 VTAIL.n765 1.93989
R2753 VTAIL.n780 VTAIL.n779 1.93989
R2754 VTAIL.n41 VTAIL.n30 1.93989
R2755 VTAIL.n75 VTAIL.n73 1.93989
R2756 VTAIL.n88 VTAIL.n87 1.93989
R2757 VTAIL.n139 VTAIL.n128 1.93989
R2758 VTAIL.n173 VTAIL.n171 1.93989
R2759 VTAIL.n186 VTAIL.n185 1.93989
R2760 VTAIL.n239 VTAIL.n228 1.93989
R2761 VTAIL.n273 VTAIL.n271 1.93989
R2762 VTAIL.n286 VTAIL.n285 1.93989
R2763 VTAIL.n682 VTAIL.n681 1.93989
R2764 VTAIL.n670 VTAIL.n669 1.93989
R2765 VTAIL.n637 VTAIL.n626 1.93989
R2766 VTAIL.n582 VTAIL.n581 1.93989
R2767 VTAIL.n570 VTAIL.n569 1.93989
R2768 VTAIL.n537 VTAIL.n526 1.93989
R2769 VTAIL.n484 VTAIL.n483 1.93989
R2770 VTAIL.n472 VTAIL.n471 1.93989
R2771 VTAIL.n439 VTAIL.n428 1.93989
R2772 VTAIL.n384 VTAIL.n383 1.93989
R2773 VTAIL.n372 VTAIL.n371 1.93989
R2774 VTAIL.n339 VTAIL.n328 1.93989
R2775 VTAIL.n397 VTAIL.n395 1.74188
R2776 VTAIL.n495 VTAIL.n397 1.74188
R2777 VTAIL.n595 VTAIL.n593 1.74188
R2778 VTAIL.n693 VTAIL.n595 1.74188
R2779 VTAIL.n297 VTAIL.n199 1.74188
R2780 VTAIL.n199 VTAIL.n197 1.74188
R2781 VTAIL.n99 VTAIL.n1 1.74188
R2782 VTAIL VTAIL.n791 1.68369
R2783 VTAIL.n730 VTAIL.n729 1.16414
R2784 VTAIL.n766 VTAIL.n704 1.16414
R2785 VTAIL.n776 VTAIL.n700 1.16414
R2786 VTAIL.n38 VTAIL.n37 1.16414
R2787 VTAIL.n74 VTAIL.n12 1.16414
R2788 VTAIL.n84 VTAIL.n8 1.16414
R2789 VTAIL.n136 VTAIL.n135 1.16414
R2790 VTAIL.n172 VTAIL.n110 1.16414
R2791 VTAIL.n182 VTAIL.n106 1.16414
R2792 VTAIL.n236 VTAIL.n235 1.16414
R2793 VTAIL.n272 VTAIL.n210 1.16414
R2794 VTAIL.n282 VTAIL.n206 1.16414
R2795 VTAIL.n678 VTAIL.n602 1.16414
R2796 VTAIL.n673 VTAIL.n607 1.16414
R2797 VTAIL.n634 VTAIL.n633 1.16414
R2798 VTAIL.n578 VTAIL.n502 1.16414
R2799 VTAIL.n573 VTAIL.n507 1.16414
R2800 VTAIL.n534 VTAIL.n533 1.16414
R2801 VTAIL.n480 VTAIL.n404 1.16414
R2802 VTAIL.n475 VTAIL.n409 1.16414
R2803 VTAIL.n436 VTAIL.n435 1.16414
R2804 VTAIL.n380 VTAIL.n304 1.16414
R2805 VTAIL.n375 VTAIL.n309 1.16414
R2806 VTAIL.n336 VTAIL.n335 1.16414
R2807 VTAIL.n0 VTAIL.t8 1.13517
R2808 VTAIL.n0 VTAIL.t13 1.13517
R2809 VTAIL.n198 VTAIL.t4 1.13517
R2810 VTAIL.n198 VTAIL.t7 1.13517
R2811 VTAIL.n594 VTAIL.t5 1.13517
R2812 VTAIL.n594 VTAIL.t2 1.13517
R2813 VTAIL.n396 VTAIL.t11 1.13517
R2814 VTAIL.n396 VTAIL.t15 1.13517
R2815 VTAIL.n593 VTAIL.n495 0.470328
R2816 VTAIL.n197 VTAIL.n99 0.470328
R2817 VTAIL.n726 VTAIL.n724 0.388379
R2818 VTAIL.n772 VTAIL.n771 0.388379
R2819 VTAIL.n775 VTAIL.n702 0.388379
R2820 VTAIL.n34 VTAIL.n32 0.388379
R2821 VTAIL.n80 VTAIL.n79 0.388379
R2822 VTAIL.n83 VTAIL.n10 0.388379
R2823 VTAIL.n132 VTAIL.n130 0.388379
R2824 VTAIL.n178 VTAIL.n177 0.388379
R2825 VTAIL.n181 VTAIL.n108 0.388379
R2826 VTAIL.n232 VTAIL.n230 0.388379
R2827 VTAIL.n278 VTAIL.n277 0.388379
R2828 VTAIL.n281 VTAIL.n208 0.388379
R2829 VTAIL.n677 VTAIL.n604 0.388379
R2830 VTAIL.n674 VTAIL.n606 0.388379
R2831 VTAIL.n630 VTAIL.n628 0.388379
R2832 VTAIL.n577 VTAIL.n504 0.388379
R2833 VTAIL.n574 VTAIL.n506 0.388379
R2834 VTAIL.n530 VTAIL.n528 0.388379
R2835 VTAIL.n479 VTAIL.n406 0.388379
R2836 VTAIL.n476 VTAIL.n408 0.388379
R2837 VTAIL.n432 VTAIL.n430 0.388379
R2838 VTAIL.n379 VTAIL.n306 0.388379
R2839 VTAIL.n376 VTAIL.n308 0.388379
R2840 VTAIL.n332 VTAIL.n330 0.388379
R2841 VTAIL.n731 VTAIL.n723 0.155672
R2842 VTAIL.n732 VTAIL.n731 0.155672
R2843 VTAIL.n732 VTAIL.n719 0.155672
R2844 VTAIL.n739 VTAIL.n719 0.155672
R2845 VTAIL.n740 VTAIL.n739 0.155672
R2846 VTAIL.n740 VTAIL.n715 0.155672
R2847 VTAIL.n747 VTAIL.n715 0.155672
R2848 VTAIL.n748 VTAIL.n747 0.155672
R2849 VTAIL.n748 VTAIL.n711 0.155672
R2850 VTAIL.n755 VTAIL.n711 0.155672
R2851 VTAIL.n756 VTAIL.n755 0.155672
R2852 VTAIL.n756 VTAIL.n707 0.155672
R2853 VTAIL.n763 VTAIL.n707 0.155672
R2854 VTAIL.n764 VTAIL.n763 0.155672
R2855 VTAIL.n764 VTAIL.n703 0.155672
R2856 VTAIL.n773 VTAIL.n703 0.155672
R2857 VTAIL.n774 VTAIL.n773 0.155672
R2858 VTAIL.n774 VTAIL.n699 0.155672
R2859 VTAIL.n781 VTAIL.n699 0.155672
R2860 VTAIL.n782 VTAIL.n781 0.155672
R2861 VTAIL.n782 VTAIL.n695 0.155672
R2862 VTAIL.n789 VTAIL.n695 0.155672
R2863 VTAIL.n39 VTAIL.n31 0.155672
R2864 VTAIL.n40 VTAIL.n39 0.155672
R2865 VTAIL.n40 VTAIL.n27 0.155672
R2866 VTAIL.n47 VTAIL.n27 0.155672
R2867 VTAIL.n48 VTAIL.n47 0.155672
R2868 VTAIL.n48 VTAIL.n23 0.155672
R2869 VTAIL.n55 VTAIL.n23 0.155672
R2870 VTAIL.n56 VTAIL.n55 0.155672
R2871 VTAIL.n56 VTAIL.n19 0.155672
R2872 VTAIL.n63 VTAIL.n19 0.155672
R2873 VTAIL.n64 VTAIL.n63 0.155672
R2874 VTAIL.n64 VTAIL.n15 0.155672
R2875 VTAIL.n71 VTAIL.n15 0.155672
R2876 VTAIL.n72 VTAIL.n71 0.155672
R2877 VTAIL.n72 VTAIL.n11 0.155672
R2878 VTAIL.n81 VTAIL.n11 0.155672
R2879 VTAIL.n82 VTAIL.n81 0.155672
R2880 VTAIL.n82 VTAIL.n7 0.155672
R2881 VTAIL.n89 VTAIL.n7 0.155672
R2882 VTAIL.n90 VTAIL.n89 0.155672
R2883 VTAIL.n90 VTAIL.n3 0.155672
R2884 VTAIL.n97 VTAIL.n3 0.155672
R2885 VTAIL.n137 VTAIL.n129 0.155672
R2886 VTAIL.n138 VTAIL.n137 0.155672
R2887 VTAIL.n138 VTAIL.n125 0.155672
R2888 VTAIL.n145 VTAIL.n125 0.155672
R2889 VTAIL.n146 VTAIL.n145 0.155672
R2890 VTAIL.n146 VTAIL.n121 0.155672
R2891 VTAIL.n153 VTAIL.n121 0.155672
R2892 VTAIL.n154 VTAIL.n153 0.155672
R2893 VTAIL.n154 VTAIL.n117 0.155672
R2894 VTAIL.n161 VTAIL.n117 0.155672
R2895 VTAIL.n162 VTAIL.n161 0.155672
R2896 VTAIL.n162 VTAIL.n113 0.155672
R2897 VTAIL.n169 VTAIL.n113 0.155672
R2898 VTAIL.n170 VTAIL.n169 0.155672
R2899 VTAIL.n170 VTAIL.n109 0.155672
R2900 VTAIL.n179 VTAIL.n109 0.155672
R2901 VTAIL.n180 VTAIL.n179 0.155672
R2902 VTAIL.n180 VTAIL.n105 0.155672
R2903 VTAIL.n187 VTAIL.n105 0.155672
R2904 VTAIL.n188 VTAIL.n187 0.155672
R2905 VTAIL.n188 VTAIL.n101 0.155672
R2906 VTAIL.n195 VTAIL.n101 0.155672
R2907 VTAIL.n237 VTAIL.n229 0.155672
R2908 VTAIL.n238 VTAIL.n237 0.155672
R2909 VTAIL.n238 VTAIL.n225 0.155672
R2910 VTAIL.n245 VTAIL.n225 0.155672
R2911 VTAIL.n246 VTAIL.n245 0.155672
R2912 VTAIL.n246 VTAIL.n221 0.155672
R2913 VTAIL.n253 VTAIL.n221 0.155672
R2914 VTAIL.n254 VTAIL.n253 0.155672
R2915 VTAIL.n254 VTAIL.n217 0.155672
R2916 VTAIL.n261 VTAIL.n217 0.155672
R2917 VTAIL.n262 VTAIL.n261 0.155672
R2918 VTAIL.n262 VTAIL.n213 0.155672
R2919 VTAIL.n269 VTAIL.n213 0.155672
R2920 VTAIL.n270 VTAIL.n269 0.155672
R2921 VTAIL.n270 VTAIL.n209 0.155672
R2922 VTAIL.n279 VTAIL.n209 0.155672
R2923 VTAIL.n280 VTAIL.n279 0.155672
R2924 VTAIL.n280 VTAIL.n205 0.155672
R2925 VTAIL.n287 VTAIL.n205 0.155672
R2926 VTAIL.n288 VTAIL.n287 0.155672
R2927 VTAIL.n288 VTAIL.n201 0.155672
R2928 VTAIL.n295 VTAIL.n201 0.155672
R2929 VTAIL.n691 VTAIL.n597 0.155672
R2930 VTAIL.n684 VTAIL.n597 0.155672
R2931 VTAIL.n684 VTAIL.n683 0.155672
R2932 VTAIL.n683 VTAIL.n601 0.155672
R2933 VTAIL.n676 VTAIL.n601 0.155672
R2934 VTAIL.n676 VTAIL.n675 0.155672
R2935 VTAIL.n675 VTAIL.n605 0.155672
R2936 VTAIL.n668 VTAIL.n605 0.155672
R2937 VTAIL.n668 VTAIL.n667 0.155672
R2938 VTAIL.n667 VTAIL.n611 0.155672
R2939 VTAIL.n660 VTAIL.n611 0.155672
R2940 VTAIL.n660 VTAIL.n659 0.155672
R2941 VTAIL.n659 VTAIL.n615 0.155672
R2942 VTAIL.n652 VTAIL.n615 0.155672
R2943 VTAIL.n652 VTAIL.n651 0.155672
R2944 VTAIL.n651 VTAIL.n619 0.155672
R2945 VTAIL.n644 VTAIL.n619 0.155672
R2946 VTAIL.n644 VTAIL.n643 0.155672
R2947 VTAIL.n643 VTAIL.n623 0.155672
R2948 VTAIL.n636 VTAIL.n623 0.155672
R2949 VTAIL.n636 VTAIL.n635 0.155672
R2950 VTAIL.n635 VTAIL.n627 0.155672
R2951 VTAIL.n591 VTAIL.n497 0.155672
R2952 VTAIL.n584 VTAIL.n497 0.155672
R2953 VTAIL.n584 VTAIL.n583 0.155672
R2954 VTAIL.n583 VTAIL.n501 0.155672
R2955 VTAIL.n576 VTAIL.n501 0.155672
R2956 VTAIL.n576 VTAIL.n575 0.155672
R2957 VTAIL.n575 VTAIL.n505 0.155672
R2958 VTAIL.n568 VTAIL.n505 0.155672
R2959 VTAIL.n568 VTAIL.n567 0.155672
R2960 VTAIL.n567 VTAIL.n511 0.155672
R2961 VTAIL.n560 VTAIL.n511 0.155672
R2962 VTAIL.n560 VTAIL.n559 0.155672
R2963 VTAIL.n559 VTAIL.n515 0.155672
R2964 VTAIL.n552 VTAIL.n515 0.155672
R2965 VTAIL.n552 VTAIL.n551 0.155672
R2966 VTAIL.n551 VTAIL.n519 0.155672
R2967 VTAIL.n544 VTAIL.n519 0.155672
R2968 VTAIL.n544 VTAIL.n543 0.155672
R2969 VTAIL.n543 VTAIL.n523 0.155672
R2970 VTAIL.n536 VTAIL.n523 0.155672
R2971 VTAIL.n536 VTAIL.n535 0.155672
R2972 VTAIL.n535 VTAIL.n527 0.155672
R2973 VTAIL.n493 VTAIL.n399 0.155672
R2974 VTAIL.n486 VTAIL.n399 0.155672
R2975 VTAIL.n486 VTAIL.n485 0.155672
R2976 VTAIL.n485 VTAIL.n403 0.155672
R2977 VTAIL.n478 VTAIL.n403 0.155672
R2978 VTAIL.n478 VTAIL.n477 0.155672
R2979 VTAIL.n477 VTAIL.n407 0.155672
R2980 VTAIL.n470 VTAIL.n407 0.155672
R2981 VTAIL.n470 VTAIL.n469 0.155672
R2982 VTAIL.n469 VTAIL.n413 0.155672
R2983 VTAIL.n462 VTAIL.n413 0.155672
R2984 VTAIL.n462 VTAIL.n461 0.155672
R2985 VTAIL.n461 VTAIL.n417 0.155672
R2986 VTAIL.n454 VTAIL.n417 0.155672
R2987 VTAIL.n454 VTAIL.n453 0.155672
R2988 VTAIL.n453 VTAIL.n421 0.155672
R2989 VTAIL.n446 VTAIL.n421 0.155672
R2990 VTAIL.n446 VTAIL.n445 0.155672
R2991 VTAIL.n445 VTAIL.n425 0.155672
R2992 VTAIL.n438 VTAIL.n425 0.155672
R2993 VTAIL.n438 VTAIL.n437 0.155672
R2994 VTAIL.n437 VTAIL.n429 0.155672
R2995 VTAIL.n393 VTAIL.n299 0.155672
R2996 VTAIL.n386 VTAIL.n299 0.155672
R2997 VTAIL.n386 VTAIL.n385 0.155672
R2998 VTAIL.n385 VTAIL.n303 0.155672
R2999 VTAIL.n378 VTAIL.n303 0.155672
R3000 VTAIL.n378 VTAIL.n377 0.155672
R3001 VTAIL.n377 VTAIL.n307 0.155672
R3002 VTAIL.n370 VTAIL.n307 0.155672
R3003 VTAIL.n370 VTAIL.n369 0.155672
R3004 VTAIL.n369 VTAIL.n313 0.155672
R3005 VTAIL.n362 VTAIL.n313 0.155672
R3006 VTAIL.n362 VTAIL.n361 0.155672
R3007 VTAIL.n361 VTAIL.n317 0.155672
R3008 VTAIL.n354 VTAIL.n317 0.155672
R3009 VTAIL.n354 VTAIL.n353 0.155672
R3010 VTAIL.n353 VTAIL.n321 0.155672
R3011 VTAIL.n346 VTAIL.n321 0.155672
R3012 VTAIL.n346 VTAIL.n345 0.155672
R3013 VTAIL.n345 VTAIL.n325 0.155672
R3014 VTAIL.n338 VTAIL.n325 0.155672
R3015 VTAIL.n338 VTAIL.n337 0.155672
R3016 VTAIL.n337 VTAIL.n329 0.155672
R3017 VTAIL VTAIL.n1 0.0586897
R3018 VP.n12 VP.t1 276.861
R3019 VP.n31 VP.t5 248.844
R3020 VP.n38 VP.t3 248.844
R3021 VP.n46 VP.t2 248.844
R3022 VP.n53 VP.t7 248.844
R3023 VP.n28 VP.t4 248.844
R3024 VP.n21 VP.t0 248.844
R3025 VP.n13 VP.t6 248.844
R3026 VP.n31 VP.n30 184.299
R3027 VP.n54 VP.n53 184.299
R3028 VP.n29 VP.n28 184.299
R3029 VP.n14 VP.n11 161.3
R3030 VP.n16 VP.n15 161.3
R3031 VP.n17 VP.n10 161.3
R3032 VP.n19 VP.n18 161.3
R3033 VP.n20 VP.n9 161.3
R3034 VP.n23 VP.n22 161.3
R3035 VP.n24 VP.n8 161.3
R3036 VP.n26 VP.n25 161.3
R3037 VP.n27 VP.n7 161.3
R3038 VP.n52 VP.n0 161.3
R3039 VP.n51 VP.n50 161.3
R3040 VP.n49 VP.n1 161.3
R3041 VP.n48 VP.n47 161.3
R3042 VP.n45 VP.n2 161.3
R3043 VP.n44 VP.n43 161.3
R3044 VP.n42 VP.n3 161.3
R3045 VP.n41 VP.n40 161.3
R3046 VP.n39 VP.n4 161.3
R3047 VP.n37 VP.n36 161.3
R3048 VP.n35 VP.n5 161.3
R3049 VP.n34 VP.n33 161.3
R3050 VP.n32 VP.n6 161.3
R3051 VP.n13 VP.n12 68.3373
R3052 VP.n30 VP.n29 50.6066
R3053 VP.n33 VP.n5 42.4359
R3054 VP.n51 VP.n1 42.4359
R3055 VP.n26 VP.n8 42.4359
R3056 VP.n40 VP.n3 40.4934
R3057 VP.n44 VP.n3 40.4934
R3058 VP.n19 VP.n10 40.4934
R3059 VP.n15 VP.n10 40.4934
R3060 VP.n37 VP.n5 38.5509
R3061 VP.n47 VP.n1 38.5509
R3062 VP.n22 VP.n8 38.5509
R3063 VP.n33 VP.n32 24.4675
R3064 VP.n40 VP.n39 24.4675
R3065 VP.n45 VP.n44 24.4675
R3066 VP.n52 VP.n51 24.4675
R3067 VP.n27 VP.n26 24.4675
R3068 VP.n20 VP.n19 24.4675
R3069 VP.n15 VP.n14 24.4675
R3070 VP.n38 VP.n37 23.9782
R3071 VP.n47 VP.n46 23.9782
R3072 VP.n22 VP.n21 23.9782
R3073 VP.n12 VP.n11 18.9029
R3074 VP.n32 VP.n31 1.46852
R3075 VP.n53 VP.n52 1.46852
R3076 VP.n28 VP.n27 1.46852
R3077 VP.n39 VP.n38 0.48984
R3078 VP.n46 VP.n45 0.48984
R3079 VP.n21 VP.n20 0.48984
R3080 VP.n14 VP.n13 0.48984
R3081 VP.n16 VP.n11 0.189894
R3082 VP.n17 VP.n16 0.189894
R3083 VP.n18 VP.n17 0.189894
R3084 VP.n18 VP.n9 0.189894
R3085 VP.n23 VP.n9 0.189894
R3086 VP.n24 VP.n23 0.189894
R3087 VP.n25 VP.n24 0.189894
R3088 VP.n25 VP.n7 0.189894
R3089 VP.n29 VP.n7 0.189894
R3090 VP.n30 VP.n6 0.189894
R3091 VP.n34 VP.n6 0.189894
R3092 VP.n35 VP.n34 0.189894
R3093 VP.n36 VP.n35 0.189894
R3094 VP.n36 VP.n4 0.189894
R3095 VP.n41 VP.n4 0.189894
R3096 VP.n42 VP.n41 0.189894
R3097 VP.n43 VP.n42 0.189894
R3098 VP.n43 VP.n2 0.189894
R3099 VP.n48 VP.n2 0.189894
R3100 VP.n49 VP.n48 0.189894
R3101 VP.n50 VP.n49 0.189894
R3102 VP.n50 VP.n0 0.189894
R3103 VP.n54 VP.n0 0.189894
R3104 VP VP.n54 0.0516364
R3105 VDD1 VDD1.n0 60.2535
R3106 VDD1.n3 VDD1.n2 60.1397
R3107 VDD1.n3 VDD1.n1 60.1397
R3108 VDD1.n5 VDD1.n4 59.3244
R3109 VDD1.n5 VDD1.n3 47.1776
R3110 VDD1.n4 VDD1.t7 1.13517
R3111 VDD1.n4 VDD1.t3 1.13517
R3112 VDD1.n0 VDD1.t6 1.13517
R3113 VDD1.n0 VDD1.t1 1.13517
R3114 VDD1.n2 VDD1.t5 1.13517
R3115 VDD1.n2 VDD1.t0 1.13517
R3116 VDD1.n1 VDD1.t2 1.13517
R3117 VDD1.n1 VDD1.t4 1.13517
R3118 VDD1 VDD1.n5 0.813
C0 VN VDD2 11.2196f
C1 VTAIL VDD1 10.6233f
C2 VP VDD1 11.491401f
C3 VTAIL VDD2 10.671599f
C4 VP VDD2 0.422381f
C5 VN VTAIL 11.0915f
C6 VN VP 7.56139f
C7 VTAIL VP 11.105599f
C8 VDD1 VDD2 1.30082f
C9 VN VDD1 0.149627f
C10 VDD2 B 4.894075f
C11 VDD1 B 5.231587f
C12 VTAIL B 12.985244f
C13 VN B 12.5994f
C14 VP B 10.885587f
C15 VDD1.t6 B 0.344494f
C16 VDD1.t1 B 0.344494f
C17 VDD1.n0 B 3.13905f
C18 VDD1.t2 B 0.344494f
C19 VDD1.t4 B 0.344494f
C20 VDD1.n1 B 3.13812f
C21 VDD1.t5 B 0.344494f
C22 VDD1.t0 B 0.344494f
C23 VDD1.n2 B 3.13812f
C24 VDD1.n3 B 3.14756f
C25 VDD1.t7 B 0.344494f
C26 VDD1.t3 B 0.344494f
C27 VDD1.n4 B 3.13235f
C28 VDD1.n5 B 3.08123f
C29 VP.n0 B 0.028448f
C30 VP.t7 B 2.30624f
C31 VP.n1 B 0.023144f
C32 VP.n2 B 0.028448f
C33 VP.t2 B 2.30624f
C34 VP.n3 B 0.022998f
C35 VP.n4 B 0.028448f
C36 VP.t3 B 2.30624f
C37 VP.n5 B 0.023144f
C38 VP.n6 B 0.028448f
C39 VP.t5 B 2.30624f
C40 VP.n7 B 0.028448f
C41 VP.t4 B 2.30624f
C42 VP.n8 B 0.023144f
C43 VP.n9 B 0.028448f
C44 VP.t0 B 2.30624f
C45 VP.n10 B 0.022998f
C46 VP.n11 B 0.180261f
C47 VP.t6 B 2.30624f
C48 VP.t1 B 2.40024f
C49 VP.n12 B 0.890963f
C50 VP.n13 B 0.858149f
C51 VP.n14 B 0.027368f
C52 VP.n15 B 0.056541f
C53 VP.n16 B 0.028448f
C54 VP.n17 B 0.028448f
C55 VP.n18 B 0.028448f
C56 VP.n19 B 0.056541f
C57 VP.n20 B 0.027368f
C58 VP.n21 B 0.809894f
C59 VP.n22 B 0.056512f
C60 VP.n23 B 0.028448f
C61 VP.n24 B 0.028448f
C62 VP.n25 B 0.028448f
C63 VP.n26 B 0.0559f
C64 VP.n27 B 0.028415f
C65 VP.n28 B 0.866379f
C66 VP.n29 B 1.58291f
C67 VP.n30 B 1.60312f
C68 VP.n31 B 0.866379f
C69 VP.n32 B 0.028415f
C70 VP.n33 B 0.0559f
C71 VP.n34 B 0.028448f
C72 VP.n35 B 0.028448f
C73 VP.n36 B 0.028448f
C74 VP.n37 B 0.056512f
C75 VP.n38 B 0.809894f
C76 VP.n39 B 0.027368f
C77 VP.n40 B 0.056541f
C78 VP.n41 B 0.028448f
C79 VP.n42 B 0.028448f
C80 VP.n43 B 0.028448f
C81 VP.n44 B 0.056541f
C82 VP.n45 B 0.027368f
C83 VP.n46 B 0.809894f
C84 VP.n47 B 0.056512f
C85 VP.n48 B 0.028448f
C86 VP.n49 B 0.028448f
C87 VP.n50 B 0.028448f
C88 VP.n51 B 0.0559f
C89 VP.n52 B 0.028415f
C90 VP.n53 B 0.866379f
C91 VP.n54 B 0.0301f
C92 VTAIL.t8 B 0.253482f
C93 VTAIL.t13 B 0.253482f
C94 VTAIL.n0 B 2.246f
C95 VTAIL.n1 B 0.294298f
C96 VTAIL.n2 B 0.024474f
C97 VTAIL.n3 B 0.018382f
C98 VTAIL.n4 B 0.009878f
C99 VTAIL.n5 B 0.023348f
C100 VTAIL.n6 B 0.010459f
C101 VTAIL.n7 B 0.018382f
C102 VTAIL.n8 B 0.009878f
C103 VTAIL.n9 B 0.023348f
C104 VTAIL.n10 B 0.010168f
C105 VTAIL.n11 B 0.018382f
C106 VTAIL.n12 B 0.010459f
C107 VTAIL.n13 B 0.023348f
C108 VTAIL.n14 B 0.010459f
C109 VTAIL.n15 B 0.018382f
C110 VTAIL.n16 B 0.009878f
C111 VTAIL.n17 B 0.023348f
C112 VTAIL.n18 B 0.010459f
C113 VTAIL.n19 B 0.018382f
C114 VTAIL.n20 B 0.009878f
C115 VTAIL.n21 B 0.023348f
C116 VTAIL.n22 B 0.010459f
C117 VTAIL.n23 B 0.018382f
C118 VTAIL.n24 B 0.009878f
C119 VTAIL.n25 B 0.023348f
C120 VTAIL.n26 B 0.010459f
C121 VTAIL.n27 B 0.018382f
C122 VTAIL.n28 B 0.009878f
C123 VTAIL.n29 B 0.023348f
C124 VTAIL.n30 B 0.010459f
C125 VTAIL.n31 B 1.40238f
C126 VTAIL.n32 B 0.009878f
C127 VTAIL.t9 B 0.038652f
C128 VTAIL.n33 B 0.131184f
C129 VTAIL.n34 B 0.013792f
C130 VTAIL.n35 B 0.017511f
C131 VTAIL.n36 B 0.023348f
C132 VTAIL.n37 B 0.010459f
C133 VTAIL.n38 B 0.009878f
C134 VTAIL.n39 B 0.018382f
C135 VTAIL.n40 B 0.018382f
C136 VTAIL.n41 B 0.009878f
C137 VTAIL.n42 B 0.010459f
C138 VTAIL.n43 B 0.023348f
C139 VTAIL.n44 B 0.023348f
C140 VTAIL.n45 B 0.010459f
C141 VTAIL.n46 B 0.009878f
C142 VTAIL.n47 B 0.018382f
C143 VTAIL.n48 B 0.018382f
C144 VTAIL.n49 B 0.009878f
C145 VTAIL.n50 B 0.010459f
C146 VTAIL.n51 B 0.023348f
C147 VTAIL.n52 B 0.023348f
C148 VTAIL.n53 B 0.010459f
C149 VTAIL.n54 B 0.009878f
C150 VTAIL.n55 B 0.018382f
C151 VTAIL.n56 B 0.018382f
C152 VTAIL.n57 B 0.009878f
C153 VTAIL.n58 B 0.010459f
C154 VTAIL.n59 B 0.023348f
C155 VTAIL.n60 B 0.023348f
C156 VTAIL.n61 B 0.010459f
C157 VTAIL.n62 B 0.009878f
C158 VTAIL.n63 B 0.018382f
C159 VTAIL.n64 B 0.018382f
C160 VTAIL.n65 B 0.009878f
C161 VTAIL.n66 B 0.010459f
C162 VTAIL.n67 B 0.023348f
C163 VTAIL.n68 B 0.023348f
C164 VTAIL.n69 B 0.010459f
C165 VTAIL.n70 B 0.009878f
C166 VTAIL.n71 B 0.018382f
C167 VTAIL.n72 B 0.018382f
C168 VTAIL.n73 B 0.009878f
C169 VTAIL.n74 B 0.009878f
C170 VTAIL.n75 B 0.010459f
C171 VTAIL.n76 B 0.023348f
C172 VTAIL.n77 B 0.023348f
C173 VTAIL.n78 B 0.023348f
C174 VTAIL.n79 B 0.010168f
C175 VTAIL.n80 B 0.009878f
C176 VTAIL.n81 B 0.018382f
C177 VTAIL.n82 B 0.018382f
C178 VTAIL.n83 B 0.009878f
C179 VTAIL.n84 B 0.010459f
C180 VTAIL.n85 B 0.023348f
C181 VTAIL.n86 B 0.023348f
C182 VTAIL.n87 B 0.010459f
C183 VTAIL.n88 B 0.009878f
C184 VTAIL.n89 B 0.018382f
C185 VTAIL.n90 B 0.018382f
C186 VTAIL.n91 B 0.009878f
C187 VTAIL.n92 B 0.010459f
C188 VTAIL.n93 B 0.023348f
C189 VTAIL.n94 B 0.048131f
C190 VTAIL.n95 B 0.010459f
C191 VTAIL.n96 B 0.009878f
C192 VTAIL.n97 B 0.040732f
C193 VTAIL.n98 B 0.026628f
C194 VTAIL.n99 B 0.145682f
C195 VTAIL.n100 B 0.024474f
C196 VTAIL.n101 B 0.018382f
C197 VTAIL.n102 B 0.009878f
C198 VTAIL.n103 B 0.023348f
C199 VTAIL.n104 B 0.010459f
C200 VTAIL.n105 B 0.018382f
C201 VTAIL.n106 B 0.009878f
C202 VTAIL.n107 B 0.023348f
C203 VTAIL.n108 B 0.010168f
C204 VTAIL.n109 B 0.018382f
C205 VTAIL.n110 B 0.010459f
C206 VTAIL.n111 B 0.023348f
C207 VTAIL.n112 B 0.010459f
C208 VTAIL.n113 B 0.018382f
C209 VTAIL.n114 B 0.009878f
C210 VTAIL.n115 B 0.023348f
C211 VTAIL.n116 B 0.010459f
C212 VTAIL.n117 B 0.018382f
C213 VTAIL.n118 B 0.009878f
C214 VTAIL.n119 B 0.023348f
C215 VTAIL.n120 B 0.010459f
C216 VTAIL.n121 B 0.018382f
C217 VTAIL.n122 B 0.009878f
C218 VTAIL.n123 B 0.023348f
C219 VTAIL.n124 B 0.010459f
C220 VTAIL.n125 B 0.018382f
C221 VTAIL.n126 B 0.009878f
C222 VTAIL.n127 B 0.023348f
C223 VTAIL.n128 B 0.010459f
C224 VTAIL.n129 B 1.40238f
C225 VTAIL.n130 B 0.009878f
C226 VTAIL.t0 B 0.038652f
C227 VTAIL.n131 B 0.131184f
C228 VTAIL.n132 B 0.013792f
C229 VTAIL.n133 B 0.017511f
C230 VTAIL.n134 B 0.023348f
C231 VTAIL.n135 B 0.010459f
C232 VTAIL.n136 B 0.009878f
C233 VTAIL.n137 B 0.018382f
C234 VTAIL.n138 B 0.018382f
C235 VTAIL.n139 B 0.009878f
C236 VTAIL.n140 B 0.010459f
C237 VTAIL.n141 B 0.023348f
C238 VTAIL.n142 B 0.023348f
C239 VTAIL.n143 B 0.010459f
C240 VTAIL.n144 B 0.009878f
C241 VTAIL.n145 B 0.018382f
C242 VTAIL.n146 B 0.018382f
C243 VTAIL.n147 B 0.009878f
C244 VTAIL.n148 B 0.010459f
C245 VTAIL.n149 B 0.023348f
C246 VTAIL.n150 B 0.023348f
C247 VTAIL.n151 B 0.010459f
C248 VTAIL.n152 B 0.009878f
C249 VTAIL.n153 B 0.018382f
C250 VTAIL.n154 B 0.018382f
C251 VTAIL.n155 B 0.009878f
C252 VTAIL.n156 B 0.010459f
C253 VTAIL.n157 B 0.023348f
C254 VTAIL.n158 B 0.023348f
C255 VTAIL.n159 B 0.010459f
C256 VTAIL.n160 B 0.009878f
C257 VTAIL.n161 B 0.018382f
C258 VTAIL.n162 B 0.018382f
C259 VTAIL.n163 B 0.009878f
C260 VTAIL.n164 B 0.010459f
C261 VTAIL.n165 B 0.023348f
C262 VTAIL.n166 B 0.023348f
C263 VTAIL.n167 B 0.010459f
C264 VTAIL.n168 B 0.009878f
C265 VTAIL.n169 B 0.018382f
C266 VTAIL.n170 B 0.018382f
C267 VTAIL.n171 B 0.009878f
C268 VTAIL.n172 B 0.009878f
C269 VTAIL.n173 B 0.010459f
C270 VTAIL.n174 B 0.023348f
C271 VTAIL.n175 B 0.023348f
C272 VTAIL.n176 B 0.023348f
C273 VTAIL.n177 B 0.010168f
C274 VTAIL.n178 B 0.009878f
C275 VTAIL.n179 B 0.018382f
C276 VTAIL.n180 B 0.018382f
C277 VTAIL.n181 B 0.009878f
C278 VTAIL.n182 B 0.010459f
C279 VTAIL.n183 B 0.023348f
C280 VTAIL.n184 B 0.023348f
C281 VTAIL.n185 B 0.010459f
C282 VTAIL.n186 B 0.009878f
C283 VTAIL.n187 B 0.018382f
C284 VTAIL.n188 B 0.018382f
C285 VTAIL.n189 B 0.009878f
C286 VTAIL.n190 B 0.010459f
C287 VTAIL.n191 B 0.023348f
C288 VTAIL.n192 B 0.048131f
C289 VTAIL.n193 B 0.010459f
C290 VTAIL.n194 B 0.009878f
C291 VTAIL.n195 B 0.040732f
C292 VTAIL.n196 B 0.026628f
C293 VTAIL.n197 B 0.145682f
C294 VTAIL.t4 B 0.253482f
C295 VTAIL.t7 B 0.253482f
C296 VTAIL.n198 B 2.246f
C297 VTAIL.n199 B 0.393996f
C298 VTAIL.n200 B 0.024474f
C299 VTAIL.n201 B 0.018382f
C300 VTAIL.n202 B 0.009878f
C301 VTAIL.n203 B 0.023348f
C302 VTAIL.n204 B 0.010459f
C303 VTAIL.n205 B 0.018382f
C304 VTAIL.n206 B 0.009878f
C305 VTAIL.n207 B 0.023348f
C306 VTAIL.n208 B 0.010168f
C307 VTAIL.n209 B 0.018382f
C308 VTAIL.n210 B 0.010459f
C309 VTAIL.n211 B 0.023348f
C310 VTAIL.n212 B 0.010459f
C311 VTAIL.n213 B 0.018382f
C312 VTAIL.n214 B 0.009878f
C313 VTAIL.n215 B 0.023348f
C314 VTAIL.n216 B 0.010459f
C315 VTAIL.n217 B 0.018382f
C316 VTAIL.n218 B 0.009878f
C317 VTAIL.n219 B 0.023348f
C318 VTAIL.n220 B 0.010459f
C319 VTAIL.n221 B 0.018382f
C320 VTAIL.n222 B 0.009878f
C321 VTAIL.n223 B 0.023348f
C322 VTAIL.n224 B 0.010459f
C323 VTAIL.n225 B 0.018382f
C324 VTAIL.n226 B 0.009878f
C325 VTAIL.n227 B 0.023348f
C326 VTAIL.n228 B 0.010459f
C327 VTAIL.n229 B 1.40238f
C328 VTAIL.n230 B 0.009878f
C329 VTAIL.t1 B 0.038652f
C330 VTAIL.n231 B 0.131184f
C331 VTAIL.n232 B 0.013792f
C332 VTAIL.n233 B 0.017511f
C333 VTAIL.n234 B 0.023348f
C334 VTAIL.n235 B 0.010459f
C335 VTAIL.n236 B 0.009878f
C336 VTAIL.n237 B 0.018382f
C337 VTAIL.n238 B 0.018382f
C338 VTAIL.n239 B 0.009878f
C339 VTAIL.n240 B 0.010459f
C340 VTAIL.n241 B 0.023348f
C341 VTAIL.n242 B 0.023348f
C342 VTAIL.n243 B 0.010459f
C343 VTAIL.n244 B 0.009878f
C344 VTAIL.n245 B 0.018382f
C345 VTAIL.n246 B 0.018382f
C346 VTAIL.n247 B 0.009878f
C347 VTAIL.n248 B 0.010459f
C348 VTAIL.n249 B 0.023348f
C349 VTAIL.n250 B 0.023348f
C350 VTAIL.n251 B 0.010459f
C351 VTAIL.n252 B 0.009878f
C352 VTAIL.n253 B 0.018382f
C353 VTAIL.n254 B 0.018382f
C354 VTAIL.n255 B 0.009878f
C355 VTAIL.n256 B 0.010459f
C356 VTAIL.n257 B 0.023348f
C357 VTAIL.n258 B 0.023348f
C358 VTAIL.n259 B 0.010459f
C359 VTAIL.n260 B 0.009878f
C360 VTAIL.n261 B 0.018382f
C361 VTAIL.n262 B 0.018382f
C362 VTAIL.n263 B 0.009878f
C363 VTAIL.n264 B 0.010459f
C364 VTAIL.n265 B 0.023348f
C365 VTAIL.n266 B 0.023348f
C366 VTAIL.n267 B 0.010459f
C367 VTAIL.n268 B 0.009878f
C368 VTAIL.n269 B 0.018382f
C369 VTAIL.n270 B 0.018382f
C370 VTAIL.n271 B 0.009878f
C371 VTAIL.n272 B 0.009878f
C372 VTAIL.n273 B 0.010459f
C373 VTAIL.n274 B 0.023348f
C374 VTAIL.n275 B 0.023348f
C375 VTAIL.n276 B 0.023348f
C376 VTAIL.n277 B 0.010168f
C377 VTAIL.n278 B 0.009878f
C378 VTAIL.n279 B 0.018382f
C379 VTAIL.n280 B 0.018382f
C380 VTAIL.n281 B 0.009878f
C381 VTAIL.n282 B 0.010459f
C382 VTAIL.n283 B 0.023348f
C383 VTAIL.n284 B 0.023348f
C384 VTAIL.n285 B 0.010459f
C385 VTAIL.n286 B 0.009878f
C386 VTAIL.n287 B 0.018382f
C387 VTAIL.n288 B 0.018382f
C388 VTAIL.n289 B 0.009878f
C389 VTAIL.n290 B 0.010459f
C390 VTAIL.n291 B 0.023348f
C391 VTAIL.n292 B 0.048131f
C392 VTAIL.n293 B 0.010459f
C393 VTAIL.n294 B 0.009878f
C394 VTAIL.n295 B 0.040732f
C395 VTAIL.n296 B 0.026628f
C396 VTAIL.n297 B 1.36173f
C397 VTAIL.n298 B 0.024474f
C398 VTAIL.n299 B 0.018382f
C399 VTAIL.n300 B 0.009878f
C400 VTAIL.n301 B 0.023348f
C401 VTAIL.n302 B 0.010459f
C402 VTAIL.n303 B 0.018382f
C403 VTAIL.n304 B 0.009878f
C404 VTAIL.n305 B 0.023348f
C405 VTAIL.n306 B 0.010168f
C406 VTAIL.n307 B 0.018382f
C407 VTAIL.n308 B 0.010168f
C408 VTAIL.n309 B 0.009878f
C409 VTAIL.n310 B 0.023348f
C410 VTAIL.n311 B 0.023348f
C411 VTAIL.n312 B 0.010459f
C412 VTAIL.n313 B 0.018382f
C413 VTAIL.n314 B 0.009878f
C414 VTAIL.n315 B 0.023348f
C415 VTAIL.n316 B 0.010459f
C416 VTAIL.n317 B 0.018382f
C417 VTAIL.n318 B 0.009878f
C418 VTAIL.n319 B 0.023348f
C419 VTAIL.n320 B 0.010459f
C420 VTAIL.n321 B 0.018382f
C421 VTAIL.n322 B 0.009878f
C422 VTAIL.n323 B 0.023348f
C423 VTAIL.n324 B 0.010459f
C424 VTAIL.n325 B 0.018382f
C425 VTAIL.n326 B 0.009878f
C426 VTAIL.n327 B 0.023348f
C427 VTAIL.n328 B 0.010459f
C428 VTAIL.n329 B 1.40238f
C429 VTAIL.n330 B 0.009878f
C430 VTAIL.t14 B 0.038652f
C431 VTAIL.n331 B 0.131184f
C432 VTAIL.n332 B 0.013792f
C433 VTAIL.n333 B 0.017511f
C434 VTAIL.n334 B 0.023348f
C435 VTAIL.n335 B 0.010459f
C436 VTAIL.n336 B 0.009878f
C437 VTAIL.n337 B 0.018382f
C438 VTAIL.n338 B 0.018382f
C439 VTAIL.n339 B 0.009878f
C440 VTAIL.n340 B 0.010459f
C441 VTAIL.n341 B 0.023348f
C442 VTAIL.n342 B 0.023348f
C443 VTAIL.n343 B 0.010459f
C444 VTAIL.n344 B 0.009878f
C445 VTAIL.n345 B 0.018382f
C446 VTAIL.n346 B 0.018382f
C447 VTAIL.n347 B 0.009878f
C448 VTAIL.n348 B 0.010459f
C449 VTAIL.n349 B 0.023348f
C450 VTAIL.n350 B 0.023348f
C451 VTAIL.n351 B 0.010459f
C452 VTAIL.n352 B 0.009878f
C453 VTAIL.n353 B 0.018382f
C454 VTAIL.n354 B 0.018382f
C455 VTAIL.n355 B 0.009878f
C456 VTAIL.n356 B 0.010459f
C457 VTAIL.n357 B 0.023348f
C458 VTAIL.n358 B 0.023348f
C459 VTAIL.n359 B 0.010459f
C460 VTAIL.n360 B 0.009878f
C461 VTAIL.n361 B 0.018382f
C462 VTAIL.n362 B 0.018382f
C463 VTAIL.n363 B 0.009878f
C464 VTAIL.n364 B 0.010459f
C465 VTAIL.n365 B 0.023348f
C466 VTAIL.n366 B 0.023348f
C467 VTAIL.n367 B 0.010459f
C468 VTAIL.n368 B 0.009878f
C469 VTAIL.n369 B 0.018382f
C470 VTAIL.n370 B 0.018382f
C471 VTAIL.n371 B 0.009878f
C472 VTAIL.n372 B 0.010459f
C473 VTAIL.n373 B 0.023348f
C474 VTAIL.n374 B 0.023348f
C475 VTAIL.n375 B 0.010459f
C476 VTAIL.n376 B 0.009878f
C477 VTAIL.n377 B 0.018382f
C478 VTAIL.n378 B 0.018382f
C479 VTAIL.n379 B 0.009878f
C480 VTAIL.n380 B 0.010459f
C481 VTAIL.n381 B 0.023348f
C482 VTAIL.n382 B 0.023348f
C483 VTAIL.n383 B 0.010459f
C484 VTAIL.n384 B 0.009878f
C485 VTAIL.n385 B 0.018382f
C486 VTAIL.n386 B 0.018382f
C487 VTAIL.n387 B 0.009878f
C488 VTAIL.n388 B 0.010459f
C489 VTAIL.n389 B 0.023348f
C490 VTAIL.n390 B 0.048131f
C491 VTAIL.n391 B 0.010459f
C492 VTAIL.n392 B 0.009878f
C493 VTAIL.n393 B 0.040732f
C494 VTAIL.n394 B 0.026628f
C495 VTAIL.n395 B 1.36173f
C496 VTAIL.t11 B 0.253482f
C497 VTAIL.t15 B 0.253482f
C498 VTAIL.n396 B 2.24601f
C499 VTAIL.n397 B 0.393985f
C500 VTAIL.n398 B 0.024474f
C501 VTAIL.n399 B 0.018382f
C502 VTAIL.n400 B 0.009878f
C503 VTAIL.n401 B 0.023348f
C504 VTAIL.n402 B 0.010459f
C505 VTAIL.n403 B 0.018382f
C506 VTAIL.n404 B 0.009878f
C507 VTAIL.n405 B 0.023348f
C508 VTAIL.n406 B 0.010168f
C509 VTAIL.n407 B 0.018382f
C510 VTAIL.n408 B 0.010168f
C511 VTAIL.n409 B 0.009878f
C512 VTAIL.n410 B 0.023348f
C513 VTAIL.n411 B 0.023348f
C514 VTAIL.n412 B 0.010459f
C515 VTAIL.n413 B 0.018382f
C516 VTAIL.n414 B 0.009878f
C517 VTAIL.n415 B 0.023348f
C518 VTAIL.n416 B 0.010459f
C519 VTAIL.n417 B 0.018382f
C520 VTAIL.n418 B 0.009878f
C521 VTAIL.n419 B 0.023348f
C522 VTAIL.n420 B 0.010459f
C523 VTAIL.n421 B 0.018382f
C524 VTAIL.n422 B 0.009878f
C525 VTAIL.n423 B 0.023348f
C526 VTAIL.n424 B 0.010459f
C527 VTAIL.n425 B 0.018382f
C528 VTAIL.n426 B 0.009878f
C529 VTAIL.n427 B 0.023348f
C530 VTAIL.n428 B 0.010459f
C531 VTAIL.n429 B 1.40238f
C532 VTAIL.n430 B 0.009878f
C533 VTAIL.t10 B 0.038652f
C534 VTAIL.n431 B 0.131184f
C535 VTAIL.n432 B 0.013792f
C536 VTAIL.n433 B 0.017511f
C537 VTAIL.n434 B 0.023348f
C538 VTAIL.n435 B 0.010459f
C539 VTAIL.n436 B 0.009878f
C540 VTAIL.n437 B 0.018382f
C541 VTAIL.n438 B 0.018382f
C542 VTAIL.n439 B 0.009878f
C543 VTAIL.n440 B 0.010459f
C544 VTAIL.n441 B 0.023348f
C545 VTAIL.n442 B 0.023348f
C546 VTAIL.n443 B 0.010459f
C547 VTAIL.n444 B 0.009878f
C548 VTAIL.n445 B 0.018382f
C549 VTAIL.n446 B 0.018382f
C550 VTAIL.n447 B 0.009878f
C551 VTAIL.n448 B 0.010459f
C552 VTAIL.n449 B 0.023348f
C553 VTAIL.n450 B 0.023348f
C554 VTAIL.n451 B 0.010459f
C555 VTAIL.n452 B 0.009878f
C556 VTAIL.n453 B 0.018382f
C557 VTAIL.n454 B 0.018382f
C558 VTAIL.n455 B 0.009878f
C559 VTAIL.n456 B 0.010459f
C560 VTAIL.n457 B 0.023348f
C561 VTAIL.n458 B 0.023348f
C562 VTAIL.n459 B 0.010459f
C563 VTAIL.n460 B 0.009878f
C564 VTAIL.n461 B 0.018382f
C565 VTAIL.n462 B 0.018382f
C566 VTAIL.n463 B 0.009878f
C567 VTAIL.n464 B 0.010459f
C568 VTAIL.n465 B 0.023348f
C569 VTAIL.n466 B 0.023348f
C570 VTAIL.n467 B 0.010459f
C571 VTAIL.n468 B 0.009878f
C572 VTAIL.n469 B 0.018382f
C573 VTAIL.n470 B 0.018382f
C574 VTAIL.n471 B 0.009878f
C575 VTAIL.n472 B 0.010459f
C576 VTAIL.n473 B 0.023348f
C577 VTAIL.n474 B 0.023348f
C578 VTAIL.n475 B 0.010459f
C579 VTAIL.n476 B 0.009878f
C580 VTAIL.n477 B 0.018382f
C581 VTAIL.n478 B 0.018382f
C582 VTAIL.n479 B 0.009878f
C583 VTAIL.n480 B 0.010459f
C584 VTAIL.n481 B 0.023348f
C585 VTAIL.n482 B 0.023348f
C586 VTAIL.n483 B 0.010459f
C587 VTAIL.n484 B 0.009878f
C588 VTAIL.n485 B 0.018382f
C589 VTAIL.n486 B 0.018382f
C590 VTAIL.n487 B 0.009878f
C591 VTAIL.n488 B 0.010459f
C592 VTAIL.n489 B 0.023348f
C593 VTAIL.n490 B 0.048131f
C594 VTAIL.n491 B 0.010459f
C595 VTAIL.n492 B 0.009878f
C596 VTAIL.n493 B 0.040732f
C597 VTAIL.n494 B 0.026628f
C598 VTAIL.n495 B 0.145682f
C599 VTAIL.n496 B 0.024474f
C600 VTAIL.n497 B 0.018382f
C601 VTAIL.n498 B 0.009878f
C602 VTAIL.n499 B 0.023348f
C603 VTAIL.n500 B 0.010459f
C604 VTAIL.n501 B 0.018382f
C605 VTAIL.n502 B 0.009878f
C606 VTAIL.n503 B 0.023348f
C607 VTAIL.n504 B 0.010168f
C608 VTAIL.n505 B 0.018382f
C609 VTAIL.n506 B 0.010168f
C610 VTAIL.n507 B 0.009878f
C611 VTAIL.n508 B 0.023348f
C612 VTAIL.n509 B 0.023348f
C613 VTAIL.n510 B 0.010459f
C614 VTAIL.n511 B 0.018382f
C615 VTAIL.n512 B 0.009878f
C616 VTAIL.n513 B 0.023348f
C617 VTAIL.n514 B 0.010459f
C618 VTAIL.n515 B 0.018382f
C619 VTAIL.n516 B 0.009878f
C620 VTAIL.n517 B 0.023348f
C621 VTAIL.n518 B 0.010459f
C622 VTAIL.n519 B 0.018382f
C623 VTAIL.n520 B 0.009878f
C624 VTAIL.n521 B 0.023348f
C625 VTAIL.n522 B 0.010459f
C626 VTAIL.n523 B 0.018382f
C627 VTAIL.n524 B 0.009878f
C628 VTAIL.n525 B 0.023348f
C629 VTAIL.n526 B 0.010459f
C630 VTAIL.n527 B 1.40238f
C631 VTAIL.n528 B 0.009878f
C632 VTAIL.t6 B 0.038652f
C633 VTAIL.n529 B 0.131184f
C634 VTAIL.n530 B 0.013792f
C635 VTAIL.n531 B 0.017511f
C636 VTAIL.n532 B 0.023348f
C637 VTAIL.n533 B 0.010459f
C638 VTAIL.n534 B 0.009878f
C639 VTAIL.n535 B 0.018382f
C640 VTAIL.n536 B 0.018382f
C641 VTAIL.n537 B 0.009878f
C642 VTAIL.n538 B 0.010459f
C643 VTAIL.n539 B 0.023348f
C644 VTAIL.n540 B 0.023348f
C645 VTAIL.n541 B 0.010459f
C646 VTAIL.n542 B 0.009878f
C647 VTAIL.n543 B 0.018382f
C648 VTAIL.n544 B 0.018382f
C649 VTAIL.n545 B 0.009878f
C650 VTAIL.n546 B 0.010459f
C651 VTAIL.n547 B 0.023348f
C652 VTAIL.n548 B 0.023348f
C653 VTAIL.n549 B 0.010459f
C654 VTAIL.n550 B 0.009878f
C655 VTAIL.n551 B 0.018382f
C656 VTAIL.n552 B 0.018382f
C657 VTAIL.n553 B 0.009878f
C658 VTAIL.n554 B 0.010459f
C659 VTAIL.n555 B 0.023348f
C660 VTAIL.n556 B 0.023348f
C661 VTAIL.n557 B 0.010459f
C662 VTAIL.n558 B 0.009878f
C663 VTAIL.n559 B 0.018382f
C664 VTAIL.n560 B 0.018382f
C665 VTAIL.n561 B 0.009878f
C666 VTAIL.n562 B 0.010459f
C667 VTAIL.n563 B 0.023348f
C668 VTAIL.n564 B 0.023348f
C669 VTAIL.n565 B 0.010459f
C670 VTAIL.n566 B 0.009878f
C671 VTAIL.n567 B 0.018382f
C672 VTAIL.n568 B 0.018382f
C673 VTAIL.n569 B 0.009878f
C674 VTAIL.n570 B 0.010459f
C675 VTAIL.n571 B 0.023348f
C676 VTAIL.n572 B 0.023348f
C677 VTAIL.n573 B 0.010459f
C678 VTAIL.n574 B 0.009878f
C679 VTAIL.n575 B 0.018382f
C680 VTAIL.n576 B 0.018382f
C681 VTAIL.n577 B 0.009878f
C682 VTAIL.n578 B 0.010459f
C683 VTAIL.n579 B 0.023348f
C684 VTAIL.n580 B 0.023348f
C685 VTAIL.n581 B 0.010459f
C686 VTAIL.n582 B 0.009878f
C687 VTAIL.n583 B 0.018382f
C688 VTAIL.n584 B 0.018382f
C689 VTAIL.n585 B 0.009878f
C690 VTAIL.n586 B 0.010459f
C691 VTAIL.n587 B 0.023348f
C692 VTAIL.n588 B 0.048131f
C693 VTAIL.n589 B 0.010459f
C694 VTAIL.n590 B 0.009878f
C695 VTAIL.n591 B 0.040732f
C696 VTAIL.n592 B 0.026628f
C697 VTAIL.n593 B 0.145682f
C698 VTAIL.t5 B 0.253482f
C699 VTAIL.t2 B 0.253482f
C700 VTAIL.n594 B 2.24601f
C701 VTAIL.n595 B 0.393985f
C702 VTAIL.n596 B 0.024474f
C703 VTAIL.n597 B 0.018382f
C704 VTAIL.n598 B 0.009878f
C705 VTAIL.n599 B 0.023348f
C706 VTAIL.n600 B 0.010459f
C707 VTAIL.n601 B 0.018382f
C708 VTAIL.n602 B 0.009878f
C709 VTAIL.n603 B 0.023348f
C710 VTAIL.n604 B 0.010168f
C711 VTAIL.n605 B 0.018382f
C712 VTAIL.n606 B 0.010168f
C713 VTAIL.n607 B 0.009878f
C714 VTAIL.n608 B 0.023348f
C715 VTAIL.n609 B 0.023348f
C716 VTAIL.n610 B 0.010459f
C717 VTAIL.n611 B 0.018382f
C718 VTAIL.n612 B 0.009878f
C719 VTAIL.n613 B 0.023348f
C720 VTAIL.n614 B 0.010459f
C721 VTAIL.n615 B 0.018382f
C722 VTAIL.n616 B 0.009878f
C723 VTAIL.n617 B 0.023348f
C724 VTAIL.n618 B 0.010459f
C725 VTAIL.n619 B 0.018382f
C726 VTAIL.n620 B 0.009878f
C727 VTAIL.n621 B 0.023348f
C728 VTAIL.n622 B 0.010459f
C729 VTAIL.n623 B 0.018382f
C730 VTAIL.n624 B 0.009878f
C731 VTAIL.n625 B 0.023348f
C732 VTAIL.n626 B 0.010459f
C733 VTAIL.n627 B 1.40238f
C734 VTAIL.n628 B 0.009878f
C735 VTAIL.t3 B 0.038652f
C736 VTAIL.n629 B 0.131184f
C737 VTAIL.n630 B 0.013792f
C738 VTAIL.n631 B 0.017511f
C739 VTAIL.n632 B 0.023348f
C740 VTAIL.n633 B 0.010459f
C741 VTAIL.n634 B 0.009878f
C742 VTAIL.n635 B 0.018382f
C743 VTAIL.n636 B 0.018382f
C744 VTAIL.n637 B 0.009878f
C745 VTAIL.n638 B 0.010459f
C746 VTAIL.n639 B 0.023348f
C747 VTAIL.n640 B 0.023348f
C748 VTAIL.n641 B 0.010459f
C749 VTAIL.n642 B 0.009878f
C750 VTAIL.n643 B 0.018382f
C751 VTAIL.n644 B 0.018382f
C752 VTAIL.n645 B 0.009878f
C753 VTAIL.n646 B 0.010459f
C754 VTAIL.n647 B 0.023348f
C755 VTAIL.n648 B 0.023348f
C756 VTAIL.n649 B 0.010459f
C757 VTAIL.n650 B 0.009878f
C758 VTAIL.n651 B 0.018382f
C759 VTAIL.n652 B 0.018382f
C760 VTAIL.n653 B 0.009878f
C761 VTAIL.n654 B 0.010459f
C762 VTAIL.n655 B 0.023348f
C763 VTAIL.n656 B 0.023348f
C764 VTAIL.n657 B 0.010459f
C765 VTAIL.n658 B 0.009878f
C766 VTAIL.n659 B 0.018382f
C767 VTAIL.n660 B 0.018382f
C768 VTAIL.n661 B 0.009878f
C769 VTAIL.n662 B 0.010459f
C770 VTAIL.n663 B 0.023348f
C771 VTAIL.n664 B 0.023348f
C772 VTAIL.n665 B 0.010459f
C773 VTAIL.n666 B 0.009878f
C774 VTAIL.n667 B 0.018382f
C775 VTAIL.n668 B 0.018382f
C776 VTAIL.n669 B 0.009878f
C777 VTAIL.n670 B 0.010459f
C778 VTAIL.n671 B 0.023348f
C779 VTAIL.n672 B 0.023348f
C780 VTAIL.n673 B 0.010459f
C781 VTAIL.n674 B 0.009878f
C782 VTAIL.n675 B 0.018382f
C783 VTAIL.n676 B 0.018382f
C784 VTAIL.n677 B 0.009878f
C785 VTAIL.n678 B 0.010459f
C786 VTAIL.n679 B 0.023348f
C787 VTAIL.n680 B 0.023348f
C788 VTAIL.n681 B 0.010459f
C789 VTAIL.n682 B 0.009878f
C790 VTAIL.n683 B 0.018382f
C791 VTAIL.n684 B 0.018382f
C792 VTAIL.n685 B 0.009878f
C793 VTAIL.n686 B 0.010459f
C794 VTAIL.n687 B 0.023348f
C795 VTAIL.n688 B 0.048131f
C796 VTAIL.n689 B 0.010459f
C797 VTAIL.n690 B 0.009878f
C798 VTAIL.n691 B 0.040732f
C799 VTAIL.n692 B 0.026628f
C800 VTAIL.n693 B 1.36173f
C801 VTAIL.n694 B 0.024474f
C802 VTAIL.n695 B 0.018382f
C803 VTAIL.n696 B 0.009878f
C804 VTAIL.n697 B 0.023348f
C805 VTAIL.n698 B 0.010459f
C806 VTAIL.n699 B 0.018382f
C807 VTAIL.n700 B 0.009878f
C808 VTAIL.n701 B 0.023348f
C809 VTAIL.n702 B 0.010168f
C810 VTAIL.n703 B 0.018382f
C811 VTAIL.n704 B 0.010459f
C812 VTAIL.n705 B 0.023348f
C813 VTAIL.n706 B 0.010459f
C814 VTAIL.n707 B 0.018382f
C815 VTAIL.n708 B 0.009878f
C816 VTAIL.n709 B 0.023348f
C817 VTAIL.n710 B 0.010459f
C818 VTAIL.n711 B 0.018382f
C819 VTAIL.n712 B 0.009878f
C820 VTAIL.n713 B 0.023348f
C821 VTAIL.n714 B 0.010459f
C822 VTAIL.n715 B 0.018382f
C823 VTAIL.n716 B 0.009878f
C824 VTAIL.n717 B 0.023348f
C825 VTAIL.n718 B 0.010459f
C826 VTAIL.n719 B 0.018382f
C827 VTAIL.n720 B 0.009878f
C828 VTAIL.n721 B 0.023348f
C829 VTAIL.n722 B 0.010459f
C830 VTAIL.n723 B 1.40238f
C831 VTAIL.n724 B 0.009878f
C832 VTAIL.t12 B 0.038652f
C833 VTAIL.n725 B 0.131184f
C834 VTAIL.n726 B 0.013792f
C835 VTAIL.n727 B 0.017511f
C836 VTAIL.n728 B 0.023348f
C837 VTAIL.n729 B 0.010459f
C838 VTAIL.n730 B 0.009878f
C839 VTAIL.n731 B 0.018382f
C840 VTAIL.n732 B 0.018382f
C841 VTAIL.n733 B 0.009878f
C842 VTAIL.n734 B 0.010459f
C843 VTAIL.n735 B 0.023348f
C844 VTAIL.n736 B 0.023348f
C845 VTAIL.n737 B 0.010459f
C846 VTAIL.n738 B 0.009878f
C847 VTAIL.n739 B 0.018382f
C848 VTAIL.n740 B 0.018382f
C849 VTAIL.n741 B 0.009878f
C850 VTAIL.n742 B 0.010459f
C851 VTAIL.n743 B 0.023348f
C852 VTAIL.n744 B 0.023348f
C853 VTAIL.n745 B 0.010459f
C854 VTAIL.n746 B 0.009878f
C855 VTAIL.n747 B 0.018382f
C856 VTAIL.n748 B 0.018382f
C857 VTAIL.n749 B 0.009878f
C858 VTAIL.n750 B 0.010459f
C859 VTAIL.n751 B 0.023348f
C860 VTAIL.n752 B 0.023348f
C861 VTAIL.n753 B 0.010459f
C862 VTAIL.n754 B 0.009878f
C863 VTAIL.n755 B 0.018382f
C864 VTAIL.n756 B 0.018382f
C865 VTAIL.n757 B 0.009878f
C866 VTAIL.n758 B 0.010459f
C867 VTAIL.n759 B 0.023348f
C868 VTAIL.n760 B 0.023348f
C869 VTAIL.n761 B 0.010459f
C870 VTAIL.n762 B 0.009878f
C871 VTAIL.n763 B 0.018382f
C872 VTAIL.n764 B 0.018382f
C873 VTAIL.n765 B 0.009878f
C874 VTAIL.n766 B 0.009878f
C875 VTAIL.n767 B 0.010459f
C876 VTAIL.n768 B 0.023348f
C877 VTAIL.n769 B 0.023348f
C878 VTAIL.n770 B 0.023348f
C879 VTAIL.n771 B 0.010168f
C880 VTAIL.n772 B 0.009878f
C881 VTAIL.n773 B 0.018382f
C882 VTAIL.n774 B 0.018382f
C883 VTAIL.n775 B 0.009878f
C884 VTAIL.n776 B 0.010459f
C885 VTAIL.n777 B 0.023348f
C886 VTAIL.n778 B 0.023348f
C887 VTAIL.n779 B 0.010459f
C888 VTAIL.n780 B 0.009878f
C889 VTAIL.n781 B 0.018382f
C890 VTAIL.n782 B 0.018382f
C891 VTAIL.n783 B 0.009878f
C892 VTAIL.n784 B 0.010459f
C893 VTAIL.n785 B 0.023348f
C894 VTAIL.n786 B 0.048131f
C895 VTAIL.n787 B 0.010459f
C896 VTAIL.n788 B 0.009878f
C897 VTAIL.n789 B 0.040732f
C898 VTAIL.n790 B 0.026628f
C899 VTAIL.n791 B 1.35828f
C900 VDD2.t5 B 0.342807f
C901 VDD2.t4 B 0.342807f
C902 VDD2.n0 B 3.12276f
C903 VDD2.t2 B 0.342807f
C904 VDD2.t1 B 0.342807f
C905 VDD2.n1 B 3.12276f
C906 VDD2.n2 B 3.08009f
C907 VDD2.t6 B 0.342807f
C908 VDD2.t3 B 0.342807f
C909 VDD2.n3 B 3.11703f
C910 VDD2.n4 B 3.0357f
C911 VDD2.t7 B 0.342807f
C912 VDD2.t0 B 0.342807f
C913 VDD2.n5 B 3.12273f
C914 VN.n0 B 0.028129f
C915 VN.t3 B 2.28031f
C916 VN.n1 B 0.022884f
C917 VN.n2 B 0.028129f
C918 VN.t2 B 2.28031f
C919 VN.n3 B 0.022739f
C920 VN.n4 B 0.178235f
C921 VN.t7 B 2.28031f
C922 VN.t6 B 2.37325f
C923 VN.n5 B 0.880946f
C924 VN.n6 B 0.848501f
C925 VN.n7 B 0.02706f
C926 VN.n8 B 0.055905f
C927 VN.n9 B 0.028129f
C928 VN.n10 B 0.028129f
C929 VN.n11 B 0.028129f
C930 VN.n12 B 0.055905f
C931 VN.n13 B 0.02706f
C932 VN.n14 B 0.800789f
C933 VN.n15 B 0.055876f
C934 VN.n16 B 0.028129f
C935 VN.n17 B 0.028129f
C936 VN.n18 B 0.028129f
C937 VN.n19 B 0.055272f
C938 VN.n20 B 0.028095f
C939 VN.n21 B 0.856638f
C940 VN.n22 B 0.029762f
C941 VN.n23 B 0.028129f
C942 VN.t1 B 2.28031f
C943 VN.n24 B 0.022884f
C944 VN.n25 B 0.028129f
C945 VN.t4 B 2.28031f
C946 VN.n26 B 0.022739f
C947 VN.n27 B 0.178235f
C948 VN.t0 B 2.28031f
C949 VN.t5 B 2.37325f
C950 VN.n28 B 0.880946f
C951 VN.n29 B 0.848501f
C952 VN.n30 B 0.02706f
C953 VN.n31 B 0.055905f
C954 VN.n32 B 0.028129f
C955 VN.n33 B 0.028129f
C956 VN.n34 B 0.028129f
C957 VN.n35 B 0.055905f
C958 VN.n36 B 0.02706f
C959 VN.n37 B 0.800789f
C960 VN.n38 B 0.055876f
C961 VN.n39 B 0.028129f
C962 VN.n40 B 0.028129f
C963 VN.n41 B 0.028129f
C964 VN.n42 B 0.055272f
C965 VN.n43 B 0.028095f
C966 VN.n44 B 0.856638f
C967 VN.n45 B 1.58339f
.ends

