* NGSPICE file created from diff_pair_sample_0870.ext - technology: sky130A

.subckt diff_pair_sample_0870 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=6.474 ps=33.98 w=16.6 l=3.55
X1 VTAIL.t19 VN.t0 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X2 VDD1.t8 VP.t1 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=2.739 ps=16.93 w=16.6 l=3.55
X3 VDD2.t8 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X4 VDD1.t7 VP.t2 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=6.474 ps=33.98 w=16.6 l=3.55
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=0 ps=0 w=16.6 l=3.55
X6 VDD2.t7 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=6.474 ps=33.98 w=16.6 l=3.55
X7 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X8 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=0 ps=0 w=16.6 l=3.55
X9 VTAIL.t8 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X10 VTAIL.t15 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X11 VTAIL.t13 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X12 VTAIL.t10 VP.t5 VDD1.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X13 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=6.474 ps=33.98 w=16.6 l=3.55
X14 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=2.739 ps=16.93 w=16.6 l=3.55
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=0 ps=0 w=16.6 l=3.55
X16 VDD1.t3 VP.t6 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X17 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=2.739 ps=16.93 w=16.6 l=3.55
X18 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=0 ps=0 w=16.6 l=3.55
X20 VTAIL.t9 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X21 VDD1.t1 VP.t8 VTAIL.t18 B.t0 sky130_fd_pr__nfet_01v8 ad=6.474 pd=33.98 as=2.739 ps=16.93 w=16.6 l=3.55
X22 VTAIL.t3 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
X23 VDD1.t0 VP.t9 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=2.739 pd=16.93 as=2.739 ps=16.93 w=16.6 l=3.55
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n21 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n20 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n19 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n18 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n4 161.3
R31 VP.n105 VP.n104 161.3
R32 VP.n102 VP.n5 161.3
R33 VP.n101 VP.n100 161.3
R34 VP.n99 VP.n6 161.3
R35 VP.n98 VP.n97 161.3
R36 VP.n96 VP.n7 161.3
R37 VP.n95 VP.n94 161.3
R38 VP.n93 VP.n8 161.3
R39 VP.n92 VP.n91 161.3
R40 VP.n90 VP.n9 161.3
R41 VP.n89 VP.n88 161.3
R42 VP.n87 VP.n10 161.3
R43 VP.n86 VP.n85 161.3
R44 VP.n84 VP.n11 161.3
R45 VP.n83 VP.n82 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n79 VP.n13 161.3
R48 VP.n78 VP.n77 161.3
R49 VP.n76 VP.n14 161.3
R50 VP.n75 VP.n74 161.3
R51 VP.n73 VP.n15 161.3
R52 VP.n72 VP.n71 161.3
R53 VP.n70 VP.n16 161.3
R54 VP.n30 VP.t1 146.381
R55 VP.n8 VP.t9 112.694
R56 VP.n68 VP.t8 112.694
R57 VP.n12 VP.t7 112.694
R58 VP.n103 VP.t3 112.694
R59 VP.n0 VP.t2 112.694
R60 VP.n25 VP.t6 112.694
R61 VP.n17 VP.t0 112.694
R62 VP.n52 VP.t5 112.694
R63 VP.n29 VP.t4 112.694
R64 VP.n69 VP.n68 77.2324
R65 VP.n118 VP.n0 77.2324
R66 VP.n67 VP.n17 77.2324
R67 VP.n69 VP.n67 61.9082
R68 VP.n74 VP.n14 56.4773
R69 VP.n110 VP.n2 56.4773
R70 VP.n59 VP.n19 56.4773
R71 VP.n30 VP.n29 55.9619
R72 VP.n89 VP.n10 46.253
R73 VP.n97 VP.n6 46.253
R74 VP.n46 VP.n23 46.253
R75 VP.n38 VP.n27 46.253
R76 VP.n85 VP.n10 34.5682
R77 VP.n101 VP.n6 34.5682
R78 VP.n50 VP.n23 34.5682
R79 VP.n34 VP.n27 34.5682
R80 VP.n72 VP.n16 24.3439
R81 VP.n73 VP.n72 24.3439
R82 VP.n74 VP.n73 24.3439
R83 VP.n78 VP.n14 24.3439
R84 VP.n79 VP.n78 24.3439
R85 VP.n80 VP.n79 24.3439
R86 VP.n84 VP.n83 24.3439
R87 VP.n85 VP.n84 24.3439
R88 VP.n90 VP.n89 24.3439
R89 VP.n91 VP.n90 24.3439
R90 VP.n91 VP.n8 24.3439
R91 VP.n95 VP.n8 24.3439
R92 VP.n96 VP.n95 24.3439
R93 VP.n97 VP.n96 24.3439
R94 VP.n102 VP.n101 24.3439
R95 VP.n104 VP.n102 24.3439
R96 VP.n108 VP.n4 24.3439
R97 VP.n109 VP.n108 24.3439
R98 VP.n110 VP.n109 24.3439
R99 VP.n114 VP.n2 24.3439
R100 VP.n115 VP.n114 24.3439
R101 VP.n116 VP.n115 24.3439
R102 VP.n63 VP.n19 24.3439
R103 VP.n64 VP.n63 24.3439
R104 VP.n65 VP.n64 24.3439
R105 VP.n51 VP.n50 24.3439
R106 VP.n53 VP.n51 24.3439
R107 VP.n57 VP.n21 24.3439
R108 VP.n58 VP.n57 24.3439
R109 VP.n59 VP.n58 24.3439
R110 VP.n39 VP.n38 24.3439
R111 VP.n40 VP.n39 24.3439
R112 VP.n40 VP.n25 24.3439
R113 VP.n44 VP.n25 24.3439
R114 VP.n45 VP.n44 24.3439
R115 VP.n46 VP.n45 24.3439
R116 VP.n33 VP.n32 24.3439
R117 VP.n34 VP.n33 24.3439
R118 VP.n83 VP.n12 18.5015
R119 VP.n104 VP.n103 18.5015
R120 VP.n53 VP.n52 18.5015
R121 VP.n32 VP.n29 18.5015
R122 VP.n68 VP.n16 12.6591
R123 VP.n116 VP.n0 12.6591
R124 VP.n65 VP.n17 12.6591
R125 VP.n80 VP.n12 5.84292
R126 VP.n103 VP.n4 5.84292
R127 VP.n52 VP.n21 5.84292
R128 VP.n31 VP.n30 3.08091
R129 VP.n67 VP.n66 0.355081
R130 VP.n70 VP.n69 0.355081
R131 VP.n118 VP.n117 0.355081
R132 VP VP.n118 0.26685
R133 VP.n31 VP.n28 0.189894
R134 VP.n35 VP.n28 0.189894
R135 VP.n36 VP.n35 0.189894
R136 VP.n37 VP.n36 0.189894
R137 VP.n37 VP.n26 0.189894
R138 VP.n41 VP.n26 0.189894
R139 VP.n42 VP.n41 0.189894
R140 VP.n43 VP.n42 0.189894
R141 VP.n43 VP.n24 0.189894
R142 VP.n47 VP.n24 0.189894
R143 VP.n48 VP.n47 0.189894
R144 VP.n49 VP.n48 0.189894
R145 VP.n49 VP.n22 0.189894
R146 VP.n54 VP.n22 0.189894
R147 VP.n55 VP.n54 0.189894
R148 VP.n56 VP.n55 0.189894
R149 VP.n56 VP.n20 0.189894
R150 VP.n60 VP.n20 0.189894
R151 VP.n61 VP.n60 0.189894
R152 VP.n62 VP.n61 0.189894
R153 VP.n62 VP.n18 0.189894
R154 VP.n66 VP.n18 0.189894
R155 VP.n71 VP.n70 0.189894
R156 VP.n71 VP.n15 0.189894
R157 VP.n75 VP.n15 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n77 VP.n76 0.189894
R160 VP.n77 VP.n13 0.189894
R161 VP.n81 VP.n13 0.189894
R162 VP.n82 VP.n81 0.189894
R163 VP.n82 VP.n11 0.189894
R164 VP.n86 VP.n11 0.189894
R165 VP.n87 VP.n86 0.189894
R166 VP.n88 VP.n87 0.189894
R167 VP.n88 VP.n9 0.189894
R168 VP.n92 VP.n9 0.189894
R169 VP.n93 VP.n92 0.189894
R170 VP.n94 VP.n93 0.189894
R171 VP.n94 VP.n7 0.189894
R172 VP.n98 VP.n7 0.189894
R173 VP.n99 VP.n98 0.189894
R174 VP.n100 VP.n99 0.189894
R175 VP.n100 VP.n5 0.189894
R176 VP.n105 VP.n5 0.189894
R177 VP.n106 VP.n105 0.189894
R178 VP.n107 VP.n106 0.189894
R179 VP.n107 VP.n3 0.189894
R180 VP.n111 VP.n3 0.189894
R181 VP.n112 VP.n111 0.189894
R182 VP.n113 VP.n112 0.189894
R183 VP.n113 VP.n1 0.189894
R184 VP.n117 VP.n1 0.189894
R185 VTAIL.n11 VTAIL.t1 48.3667
R186 VTAIL.n17 VTAIL.t7 48.3664
R187 VTAIL.n2 VTAIL.t12 48.3664
R188 VTAIL.n16 VTAIL.t14 48.3664
R189 VTAIL.n15 VTAIL.n14 47.1739
R190 VTAIL.n13 VTAIL.n12 47.1739
R191 VTAIL.n10 VTAIL.n9 47.1739
R192 VTAIL.n8 VTAIL.n7 47.1739
R193 VTAIL.n19 VTAIL.n18 47.1736
R194 VTAIL.n1 VTAIL.n0 47.1736
R195 VTAIL.n4 VTAIL.n3 47.1736
R196 VTAIL.n6 VTAIL.n5 47.1736
R197 VTAIL.n8 VTAIL.n6 33.3669
R198 VTAIL.n17 VTAIL.n16 30.0221
R199 VTAIL.n10 VTAIL.n8 3.34533
R200 VTAIL.n11 VTAIL.n10 3.34533
R201 VTAIL.n15 VTAIL.n13 3.34533
R202 VTAIL.n16 VTAIL.n15 3.34533
R203 VTAIL.n6 VTAIL.n4 3.34533
R204 VTAIL.n4 VTAIL.n2 3.34533
R205 VTAIL.n19 VTAIL.n17 3.34533
R206 VTAIL VTAIL.n1 2.56731
R207 VTAIL.n13 VTAIL.n11 2.14274
R208 VTAIL.n2 VTAIL.n1 2.14274
R209 VTAIL.n18 VTAIL.t5 1.19327
R210 VTAIL.n18 VTAIL.t8 1.19327
R211 VTAIL.n0 VTAIL.t6 1.19327
R212 VTAIL.n0 VTAIL.t3 1.19327
R213 VTAIL.n3 VTAIL.t16 1.19327
R214 VTAIL.n3 VTAIL.t15 1.19327
R215 VTAIL.n5 VTAIL.t18 1.19327
R216 VTAIL.n5 VTAIL.t9 1.19327
R217 VTAIL.n14 VTAIL.t17 1.19327
R218 VTAIL.n14 VTAIL.t10 1.19327
R219 VTAIL.n12 VTAIL.t11 1.19327
R220 VTAIL.n12 VTAIL.t13 1.19327
R221 VTAIL.n9 VTAIL.t4 1.19327
R222 VTAIL.n9 VTAIL.t19 1.19327
R223 VTAIL.n7 VTAIL.t0 1.19327
R224 VTAIL.n7 VTAIL.t2 1.19327
R225 VTAIL VTAIL.n19 0.778517
R226 VDD1.n1 VDD1.t8 68.3903
R227 VDD1.n3 VDD1.t1 68.39
R228 VDD1.n5 VDD1.n4 66.3057
R229 VDD1.n1 VDD1.n0 63.8527
R230 VDD1.n7 VDD1.n6 63.8525
R231 VDD1.n3 VDD1.n2 63.8524
R232 VDD1.n7 VDD1.n5 56.169
R233 VDD1 VDD1.n7 2.45093
R234 VDD1.n6 VDD1.t4 1.19327
R235 VDD1.n6 VDD1.t9 1.19327
R236 VDD1.n0 VDD1.t5 1.19327
R237 VDD1.n0 VDD1.t3 1.19327
R238 VDD1.n4 VDD1.t6 1.19327
R239 VDD1.n4 VDD1.t7 1.19327
R240 VDD1.n2 VDD1.t2 1.19327
R241 VDD1.n2 VDD1.t0 1.19327
R242 VDD1 VDD1.n1 0.894897
R243 VDD1.n5 VDD1.n3 0.781361
R244 B.n1223 B.n1222 585
R245 B.n440 B.n199 585
R246 B.n439 B.n438 585
R247 B.n437 B.n436 585
R248 B.n435 B.n434 585
R249 B.n433 B.n432 585
R250 B.n431 B.n430 585
R251 B.n429 B.n428 585
R252 B.n427 B.n426 585
R253 B.n425 B.n424 585
R254 B.n423 B.n422 585
R255 B.n421 B.n420 585
R256 B.n419 B.n418 585
R257 B.n417 B.n416 585
R258 B.n415 B.n414 585
R259 B.n413 B.n412 585
R260 B.n411 B.n410 585
R261 B.n409 B.n408 585
R262 B.n407 B.n406 585
R263 B.n405 B.n404 585
R264 B.n403 B.n402 585
R265 B.n401 B.n400 585
R266 B.n399 B.n398 585
R267 B.n397 B.n396 585
R268 B.n395 B.n394 585
R269 B.n393 B.n392 585
R270 B.n391 B.n390 585
R271 B.n389 B.n388 585
R272 B.n387 B.n386 585
R273 B.n385 B.n384 585
R274 B.n383 B.n382 585
R275 B.n381 B.n380 585
R276 B.n379 B.n378 585
R277 B.n377 B.n376 585
R278 B.n375 B.n374 585
R279 B.n373 B.n372 585
R280 B.n371 B.n370 585
R281 B.n369 B.n368 585
R282 B.n367 B.n366 585
R283 B.n365 B.n364 585
R284 B.n363 B.n362 585
R285 B.n361 B.n360 585
R286 B.n359 B.n358 585
R287 B.n357 B.n356 585
R288 B.n355 B.n354 585
R289 B.n353 B.n352 585
R290 B.n351 B.n350 585
R291 B.n349 B.n348 585
R292 B.n347 B.n346 585
R293 B.n345 B.n344 585
R294 B.n343 B.n342 585
R295 B.n341 B.n340 585
R296 B.n339 B.n338 585
R297 B.n337 B.n336 585
R298 B.n335 B.n334 585
R299 B.n332 B.n331 585
R300 B.n330 B.n329 585
R301 B.n328 B.n327 585
R302 B.n326 B.n325 585
R303 B.n324 B.n323 585
R304 B.n322 B.n321 585
R305 B.n320 B.n319 585
R306 B.n318 B.n317 585
R307 B.n316 B.n315 585
R308 B.n314 B.n313 585
R309 B.n311 B.n310 585
R310 B.n309 B.n308 585
R311 B.n307 B.n306 585
R312 B.n305 B.n304 585
R313 B.n303 B.n302 585
R314 B.n301 B.n300 585
R315 B.n299 B.n298 585
R316 B.n297 B.n296 585
R317 B.n295 B.n294 585
R318 B.n293 B.n292 585
R319 B.n291 B.n290 585
R320 B.n289 B.n288 585
R321 B.n287 B.n286 585
R322 B.n285 B.n284 585
R323 B.n283 B.n282 585
R324 B.n281 B.n280 585
R325 B.n279 B.n278 585
R326 B.n277 B.n276 585
R327 B.n275 B.n274 585
R328 B.n273 B.n272 585
R329 B.n271 B.n270 585
R330 B.n269 B.n268 585
R331 B.n267 B.n266 585
R332 B.n265 B.n264 585
R333 B.n263 B.n262 585
R334 B.n261 B.n260 585
R335 B.n259 B.n258 585
R336 B.n257 B.n256 585
R337 B.n255 B.n254 585
R338 B.n253 B.n252 585
R339 B.n251 B.n250 585
R340 B.n249 B.n248 585
R341 B.n247 B.n246 585
R342 B.n245 B.n244 585
R343 B.n243 B.n242 585
R344 B.n241 B.n240 585
R345 B.n239 B.n238 585
R346 B.n237 B.n236 585
R347 B.n235 B.n234 585
R348 B.n233 B.n232 585
R349 B.n231 B.n230 585
R350 B.n229 B.n228 585
R351 B.n227 B.n226 585
R352 B.n225 B.n224 585
R353 B.n223 B.n222 585
R354 B.n221 B.n220 585
R355 B.n219 B.n218 585
R356 B.n217 B.n216 585
R357 B.n215 B.n214 585
R358 B.n213 B.n212 585
R359 B.n211 B.n210 585
R360 B.n209 B.n208 585
R361 B.n207 B.n206 585
R362 B.n205 B.n204 585
R363 B.n138 B.n137 585
R364 B.n1221 B.n139 585
R365 B.n1226 B.n139 585
R366 B.n1220 B.n1219 585
R367 B.n1219 B.n135 585
R368 B.n1218 B.n134 585
R369 B.n1232 B.n134 585
R370 B.n1217 B.n133 585
R371 B.n1233 B.n133 585
R372 B.n1216 B.n132 585
R373 B.n1234 B.n132 585
R374 B.n1215 B.n1214 585
R375 B.n1214 B.n128 585
R376 B.n1213 B.n127 585
R377 B.n1240 B.n127 585
R378 B.n1212 B.n126 585
R379 B.n1241 B.n126 585
R380 B.n1211 B.n125 585
R381 B.n1242 B.n125 585
R382 B.n1210 B.n1209 585
R383 B.n1209 B.n121 585
R384 B.n1208 B.n120 585
R385 B.n1248 B.n120 585
R386 B.n1207 B.n119 585
R387 B.n1249 B.n119 585
R388 B.n1206 B.n118 585
R389 B.n1250 B.n118 585
R390 B.n1205 B.n1204 585
R391 B.n1204 B.n114 585
R392 B.n1203 B.n113 585
R393 B.n1256 B.n113 585
R394 B.n1202 B.n112 585
R395 B.n1257 B.n112 585
R396 B.n1201 B.n111 585
R397 B.n1258 B.n111 585
R398 B.n1200 B.n1199 585
R399 B.n1199 B.n107 585
R400 B.n1198 B.n106 585
R401 B.n1264 B.n106 585
R402 B.n1197 B.n105 585
R403 B.n1265 B.n105 585
R404 B.n1196 B.n104 585
R405 B.n1266 B.n104 585
R406 B.n1195 B.n1194 585
R407 B.n1194 B.n100 585
R408 B.n1193 B.n99 585
R409 B.n1272 B.n99 585
R410 B.n1192 B.n98 585
R411 B.n1273 B.n98 585
R412 B.n1191 B.n97 585
R413 B.n1274 B.n97 585
R414 B.n1190 B.n1189 585
R415 B.n1189 B.n93 585
R416 B.n1188 B.n92 585
R417 B.n1280 B.n92 585
R418 B.n1187 B.n91 585
R419 B.n1281 B.n91 585
R420 B.n1186 B.n90 585
R421 B.n1282 B.n90 585
R422 B.n1185 B.n1184 585
R423 B.n1184 B.n86 585
R424 B.n1183 B.n85 585
R425 B.n1288 B.n85 585
R426 B.n1182 B.n84 585
R427 B.n1289 B.n84 585
R428 B.n1181 B.n83 585
R429 B.n1290 B.n83 585
R430 B.n1180 B.n1179 585
R431 B.n1179 B.n79 585
R432 B.n1178 B.n78 585
R433 B.n1296 B.n78 585
R434 B.n1177 B.n77 585
R435 B.n1297 B.n77 585
R436 B.n1176 B.n76 585
R437 B.n1298 B.n76 585
R438 B.n1175 B.n1174 585
R439 B.n1174 B.n72 585
R440 B.n1173 B.n71 585
R441 B.n1304 B.n71 585
R442 B.n1172 B.n70 585
R443 B.n1305 B.n70 585
R444 B.n1171 B.n69 585
R445 B.n1306 B.n69 585
R446 B.n1170 B.n1169 585
R447 B.n1169 B.n65 585
R448 B.n1168 B.n64 585
R449 B.n1312 B.n64 585
R450 B.n1167 B.n63 585
R451 B.n1313 B.n63 585
R452 B.n1166 B.n62 585
R453 B.n1314 B.n62 585
R454 B.n1165 B.n1164 585
R455 B.n1164 B.n58 585
R456 B.n1163 B.n57 585
R457 B.n1320 B.n57 585
R458 B.n1162 B.n56 585
R459 B.n1321 B.n56 585
R460 B.n1161 B.n55 585
R461 B.n1322 B.n55 585
R462 B.n1160 B.n1159 585
R463 B.n1159 B.n51 585
R464 B.n1158 B.n50 585
R465 B.n1328 B.n50 585
R466 B.n1157 B.n49 585
R467 B.n1329 B.n49 585
R468 B.n1156 B.n48 585
R469 B.n1330 B.n48 585
R470 B.n1155 B.n1154 585
R471 B.n1154 B.n44 585
R472 B.n1153 B.n43 585
R473 B.n1336 B.n43 585
R474 B.n1152 B.n42 585
R475 B.n1337 B.n42 585
R476 B.n1151 B.n41 585
R477 B.n1338 B.n41 585
R478 B.n1150 B.n1149 585
R479 B.n1149 B.n40 585
R480 B.n1148 B.n36 585
R481 B.n1344 B.n36 585
R482 B.n1147 B.n35 585
R483 B.n1345 B.n35 585
R484 B.n1146 B.n34 585
R485 B.n1346 B.n34 585
R486 B.n1145 B.n1144 585
R487 B.n1144 B.n30 585
R488 B.n1143 B.n29 585
R489 B.n1352 B.n29 585
R490 B.n1142 B.n28 585
R491 B.n1353 B.n28 585
R492 B.n1141 B.n27 585
R493 B.n1354 B.n27 585
R494 B.n1140 B.n1139 585
R495 B.n1139 B.n23 585
R496 B.n1138 B.n22 585
R497 B.n1360 B.n22 585
R498 B.n1137 B.n21 585
R499 B.n1361 B.n21 585
R500 B.n1136 B.n20 585
R501 B.n1362 B.n20 585
R502 B.n1135 B.n1134 585
R503 B.n1134 B.n19 585
R504 B.n1133 B.n15 585
R505 B.n1368 B.n15 585
R506 B.n1132 B.n14 585
R507 B.n1369 B.n14 585
R508 B.n1131 B.n13 585
R509 B.n1370 B.n13 585
R510 B.n1130 B.n1129 585
R511 B.n1129 B.n12 585
R512 B.n1128 B.n1127 585
R513 B.n1128 B.n8 585
R514 B.n1126 B.n7 585
R515 B.n1377 B.n7 585
R516 B.n1125 B.n6 585
R517 B.n1378 B.n6 585
R518 B.n1124 B.n5 585
R519 B.n1379 B.n5 585
R520 B.n1123 B.n1122 585
R521 B.n1122 B.n4 585
R522 B.n1121 B.n441 585
R523 B.n1121 B.n1120 585
R524 B.n1111 B.n442 585
R525 B.n443 B.n442 585
R526 B.n1113 B.n1112 585
R527 B.n1114 B.n1113 585
R528 B.n1110 B.n448 585
R529 B.n448 B.n447 585
R530 B.n1109 B.n1108 585
R531 B.n1108 B.n1107 585
R532 B.n450 B.n449 585
R533 B.n1100 B.n450 585
R534 B.n1099 B.n1098 585
R535 B.n1101 B.n1099 585
R536 B.n1097 B.n455 585
R537 B.n455 B.n454 585
R538 B.n1096 B.n1095 585
R539 B.n1095 B.n1094 585
R540 B.n457 B.n456 585
R541 B.n458 B.n457 585
R542 B.n1087 B.n1086 585
R543 B.n1088 B.n1087 585
R544 B.n1085 B.n463 585
R545 B.n463 B.n462 585
R546 B.n1084 B.n1083 585
R547 B.n1083 B.n1082 585
R548 B.n465 B.n464 585
R549 B.n466 B.n465 585
R550 B.n1075 B.n1074 585
R551 B.n1076 B.n1075 585
R552 B.n1073 B.n471 585
R553 B.n471 B.n470 585
R554 B.n1072 B.n1071 585
R555 B.n1071 B.n1070 585
R556 B.n473 B.n472 585
R557 B.n1063 B.n473 585
R558 B.n1062 B.n1061 585
R559 B.n1064 B.n1062 585
R560 B.n1060 B.n478 585
R561 B.n478 B.n477 585
R562 B.n1059 B.n1058 585
R563 B.n1058 B.n1057 585
R564 B.n480 B.n479 585
R565 B.n481 B.n480 585
R566 B.n1050 B.n1049 585
R567 B.n1051 B.n1050 585
R568 B.n1048 B.n486 585
R569 B.n486 B.n485 585
R570 B.n1047 B.n1046 585
R571 B.n1046 B.n1045 585
R572 B.n488 B.n487 585
R573 B.n489 B.n488 585
R574 B.n1038 B.n1037 585
R575 B.n1039 B.n1038 585
R576 B.n1036 B.n494 585
R577 B.n494 B.n493 585
R578 B.n1035 B.n1034 585
R579 B.n1034 B.n1033 585
R580 B.n496 B.n495 585
R581 B.n497 B.n496 585
R582 B.n1026 B.n1025 585
R583 B.n1027 B.n1026 585
R584 B.n1024 B.n502 585
R585 B.n502 B.n501 585
R586 B.n1023 B.n1022 585
R587 B.n1022 B.n1021 585
R588 B.n504 B.n503 585
R589 B.n505 B.n504 585
R590 B.n1014 B.n1013 585
R591 B.n1015 B.n1014 585
R592 B.n1012 B.n510 585
R593 B.n510 B.n509 585
R594 B.n1011 B.n1010 585
R595 B.n1010 B.n1009 585
R596 B.n512 B.n511 585
R597 B.n513 B.n512 585
R598 B.n1002 B.n1001 585
R599 B.n1003 B.n1002 585
R600 B.n1000 B.n518 585
R601 B.n518 B.n517 585
R602 B.n999 B.n998 585
R603 B.n998 B.n997 585
R604 B.n520 B.n519 585
R605 B.n521 B.n520 585
R606 B.n990 B.n989 585
R607 B.n991 B.n990 585
R608 B.n988 B.n526 585
R609 B.n526 B.n525 585
R610 B.n987 B.n986 585
R611 B.n986 B.n985 585
R612 B.n528 B.n527 585
R613 B.n529 B.n528 585
R614 B.n978 B.n977 585
R615 B.n979 B.n978 585
R616 B.n976 B.n534 585
R617 B.n534 B.n533 585
R618 B.n975 B.n974 585
R619 B.n974 B.n973 585
R620 B.n536 B.n535 585
R621 B.n537 B.n536 585
R622 B.n966 B.n965 585
R623 B.n967 B.n966 585
R624 B.n964 B.n541 585
R625 B.n545 B.n541 585
R626 B.n963 B.n962 585
R627 B.n962 B.n961 585
R628 B.n543 B.n542 585
R629 B.n544 B.n543 585
R630 B.n954 B.n953 585
R631 B.n955 B.n954 585
R632 B.n952 B.n550 585
R633 B.n550 B.n549 585
R634 B.n951 B.n950 585
R635 B.n950 B.n949 585
R636 B.n552 B.n551 585
R637 B.n553 B.n552 585
R638 B.n942 B.n941 585
R639 B.n943 B.n942 585
R640 B.n940 B.n558 585
R641 B.n558 B.n557 585
R642 B.n939 B.n938 585
R643 B.n938 B.n937 585
R644 B.n560 B.n559 585
R645 B.n561 B.n560 585
R646 B.n930 B.n929 585
R647 B.n931 B.n930 585
R648 B.n928 B.n566 585
R649 B.n566 B.n565 585
R650 B.n927 B.n926 585
R651 B.n926 B.n925 585
R652 B.n568 B.n567 585
R653 B.n569 B.n568 585
R654 B.n918 B.n917 585
R655 B.n919 B.n918 585
R656 B.n916 B.n574 585
R657 B.n574 B.n573 585
R658 B.n915 B.n914 585
R659 B.n914 B.n913 585
R660 B.n576 B.n575 585
R661 B.n577 B.n576 585
R662 B.n906 B.n905 585
R663 B.n907 B.n906 585
R664 B.n904 B.n582 585
R665 B.n582 B.n581 585
R666 B.n903 B.n902 585
R667 B.n902 B.n901 585
R668 B.n584 B.n583 585
R669 B.n585 B.n584 585
R670 B.n894 B.n893 585
R671 B.n895 B.n894 585
R672 B.n588 B.n587 585
R673 B.n657 B.n656 585
R674 B.n658 B.n654 585
R675 B.n654 B.n589 585
R676 B.n660 B.n659 585
R677 B.n662 B.n653 585
R678 B.n665 B.n664 585
R679 B.n666 B.n652 585
R680 B.n668 B.n667 585
R681 B.n670 B.n651 585
R682 B.n673 B.n672 585
R683 B.n674 B.n650 585
R684 B.n676 B.n675 585
R685 B.n678 B.n649 585
R686 B.n681 B.n680 585
R687 B.n682 B.n648 585
R688 B.n684 B.n683 585
R689 B.n686 B.n647 585
R690 B.n689 B.n688 585
R691 B.n690 B.n646 585
R692 B.n692 B.n691 585
R693 B.n694 B.n645 585
R694 B.n697 B.n696 585
R695 B.n698 B.n644 585
R696 B.n700 B.n699 585
R697 B.n702 B.n643 585
R698 B.n705 B.n704 585
R699 B.n706 B.n642 585
R700 B.n708 B.n707 585
R701 B.n710 B.n641 585
R702 B.n713 B.n712 585
R703 B.n714 B.n640 585
R704 B.n716 B.n715 585
R705 B.n718 B.n639 585
R706 B.n721 B.n720 585
R707 B.n722 B.n638 585
R708 B.n724 B.n723 585
R709 B.n726 B.n637 585
R710 B.n729 B.n728 585
R711 B.n730 B.n636 585
R712 B.n732 B.n731 585
R713 B.n734 B.n635 585
R714 B.n737 B.n736 585
R715 B.n738 B.n634 585
R716 B.n740 B.n739 585
R717 B.n742 B.n633 585
R718 B.n745 B.n744 585
R719 B.n746 B.n632 585
R720 B.n748 B.n747 585
R721 B.n750 B.n631 585
R722 B.n753 B.n752 585
R723 B.n754 B.n630 585
R724 B.n756 B.n755 585
R725 B.n758 B.n629 585
R726 B.n761 B.n760 585
R727 B.n762 B.n626 585
R728 B.n765 B.n764 585
R729 B.n767 B.n625 585
R730 B.n770 B.n769 585
R731 B.n771 B.n624 585
R732 B.n773 B.n772 585
R733 B.n775 B.n623 585
R734 B.n778 B.n777 585
R735 B.n779 B.n622 585
R736 B.n781 B.n780 585
R737 B.n783 B.n621 585
R738 B.n786 B.n785 585
R739 B.n787 B.n617 585
R740 B.n789 B.n788 585
R741 B.n791 B.n616 585
R742 B.n794 B.n793 585
R743 B.n795 B.n615 585
R744 B.n797 B.n796 585
R745 B.n799 B.n614 585
R746 B.n802 B.n801 585
R747 B.n803 B.n613 585
R748 B.n805 B.n804 585
R749 B.n807 B.n612 585
R750 B.n810 B.n809 585
R751 B.n811 B.n611 585
R752 B.n813 B.n812 585
R753 B.n815 B.n610 585
R754 B.n818 B.n817 585
R755 B.n819 B.n609 585
R756 B.n821 B.n820 585
R757 B.n823 B.n608 585
R758 B.n826 B.n825 585
R759 B.n827 B.n607 585
R760 B.n829 B.n828 585
R761 B.n831 B.n606 585
R762 B.n834 B.n833 585
R763 B.n835 B.n605 585
R764 B.n837 B.n836 585
R765 B.n839 B.n604 585
R766 B.n842 B.n841 585
R767 B.n843 B.n603 585
R768 B.n845 B.n844 585
R769 B.n847 B.n602 585
R770 B.n850 B.n849 585
R771 B.n851 B.n601 585
R772 B.n853 B.n852 585
R773 B.n855 B.n600 585
R774 B.n858 B.n857 585
R775 B.n859 B.n599 585
R776 B.n861 B.n860 585
R777 B.n863 B.n598 585
R778 B.n866 B.n865 585
R779 B.n867 B.n597 585
R780 B.n869 B.n868 585
R781 B.n871 B.n596 585
R782 B.n874 B.n873 585
R783 B.n875 B.n595 585
R784 B.n877 B.n876 585
R785 B.n879 B.n594 585
R786 B.n882 B.n881 585
R787 B.n883 B.n593 585
R788 B.n885 B.n884 585
R789 B.n887 B.n592 585
R790 B.n888 B.n591 585
R791 B.n891 B.n890 585
R792 B.n892 B.n590 585
R793 B.n590 B.n589 585
R794 B.n897 B.n896 585
R795 B.n896 B.n895 585
R796 B.n898 B.n586 585
R797 B.n586 B.n585 585
R798 B.n900 B.n899 585
R799 B.n901 B.n900 585
R800 B.n580 B.n579 585
R801 B.n581 B.n580 585
R802 B.n909 B.n908 585
R803 B.n908 B.n907 585
R804 B.n910 B.n578 585
R805 B.n578 B.n577 585
R806 B.n912 B.n911 585
R807 B.n913 B.n912 585
R808 B.n572 B.n571 585
R809 B.n573 B.n572 585
R810 B.n921 B.n920 585
R811 B.n920 B.n919 585
R812 B.n922 B.n570 585
R813 B.n570 B.n569 585
R814 B.n924 B.n923 585
R815 B.n925 B.n924 585
R816 B.n564 B.n563 585
R817 B.n565 B.n564 585
R818 B.n933 B.n932 585
R819 B.n932 B.n931 585
R820 B.n934 B.n562 585
R821 B.n562 B.n561 585
R822 B.n936 B.n935 585
R823 B.n937 B.n936 585
R824 B.n556 B.n555 585
R825 B.n557 B.n556 585
R826 B.n945 B.n944 585
R827 B.n944 B.n943 585
R828 B.n946 B.n554 585
R829 B.n554 B.n553 585
R830 B.n948 B.n947 585
R831 B.n949 B.n948 585
R832 B.n548 B.n547 585
R833 B.n549 B.n548 585
R834 B.n957 B.n956 585
R835 B.n956 B.n955 585
R836 B.n958 B.n546 585
R837 B.n546 B.n544 585
R838 B.n960 B.n959 585
R839 B.n961 B.n960 585
R840 B.n540 B.n539 585
R841 B.n545 B.n540 585
R842 B.n969 B.n968 585
R843 B.n968 B.n967 585
R844 B.n970 B.n538 585
R845 B.n538 B.n537 585
R846 B.n972 B.n971 585
R847 B.n973 B.n972 585
R848 B.n532 B.n531 585
R849 B.n533 B.n532 585
R850 B.n981 B.n980 585
R851 B.n980 B.n979 585
R852 B.n982 B.n530 585
R853 B.n530 B.n529 585
R854 B.n984 B.n983 585
R855 B.n985 B.n984 585
R856 B.n524 B.n523 585
R857 B.n525 B.n524 585
R858 B.n993 B.n992 585
R859 B.n992 B.n991 585
R860 B.n994 B.n522 585
R861 B.n522 B.n521 585
R862 B.n996 B.n995 585
R863 B.n997 B.n996 585
R864 B.n516 B.n515 585
R865 B.n517 B.n516 585
R866 B.n1005 B.n1004 585
R867 B.n1004 B.n1003 585
R868 B.n1006 B.n514 585
R869 B.n514 B.n513 585
R870 B.n1008 B.n1007 585
R871 B.n1009 B.n1008 585
R872 B.n508 B.n507 585
R873 B.n509 B.n508 585
R874 B.n1017 B.n1016 585
R875 B.n1016 B.n1015 585
R876 B.n1018 B.n506 585
R877 B.n506 B.n505 585
R878 B.n1020 B.n1019 585
R879 B.n1021 B.n1020 585
R880 B.n500 B.n499 585
R881 B.n501 B.n500 585
R882 B.n1029 B.n1028 585
R883 B.n1028 B.n1027 585
R884 B.n1030 B.n498 585
R885 B.n498 B.n497 585
R886 B.n1032 B.n1031 585
R887 B.n1033 B.n1032 585
R888 B.n492 B.n491 585
R889 B.n493 B.n492 585
R890 B.n1041 B.n1040 585
R891 B.n1040 B.n1039 585
R892 B.n1042 B.n490 585
R893 B.n490 B.n489 585
R894 B.n1044 B.n1043 585
R895 B.n1045 B.n1044 585
R896 B.n484 B.n483 585
R897 B.n485 B.n484 585
R898 B.n1053 B.n1052 585
R899 B.n1052 B.n1051 585
R900 B.n1054 B.n482 585
R901 B.n482 B.n481 585
R902 B.n1056 B.n1055 585
R903 B.n1057 B.n1056 585
R904 B.n476 B.n475 585
R905 B.n477 B.n476 585
R906 B.n1066 B.n1065 585
R907 B.n1065 B.n1064 585
R908 B.n1067 B.n474 585
R909 B.n1063 B.n474 585
R910 B.n1069 B.n1068 585
R911 B.n1070 B.n1069 585
R912 B.n469 B.n468 585
R913 B.n470 B.n469 585
R914 B.n1078 B.n1077 585
R915 B.n1077 B.n1076 585
R916 B.n1079 B.n467 585
R917 B.n467 B.n466 585
R918 B.n1081 B.n1080 585
R919 B.n1082 B.n1081 585
R920 B.n461 B.n460 585
R921 B.n462 B.n461 585
R922 B.n1090 B.n1089 585
R923 B.n1089 B.n1088 585
R924 B.n1091 B.n459 585
R925 B.n459 B.n458 585
R926 B.n1093 B.n1092 585
R927 B.n1094 B.n1093 585
R928 B.n453 B.n452 585
R929 B.n454 B.n453 585
R930 B.n1103 B.n1102 585
R931 B.n1102 B.n1101 585
R932 B.n1104 B.n451 585
R933 B.n1100 B.n451 585
R934 B.n1106 B.n1105 585
R935 B.n1107 B.n1106 585
R936 B.n446 B.n445 585
R937 B.n447 B.n446 585
R938 B.n1116 B.n1115 585
R939 B.n1115 B.n1114 585
R940 B.n1117 B.n444 585
R941 B.n444 B.n443 585
R942 B.n1119 B.n1118 585
R943 B.n1120 B.n1119 585
R944 B.n3 B.n0 585
R945 B.n4 B.n3 585
R946 B.n1376 B.n1 585
R947 B.n1377 B.n1376 585
R948 B.n1375 B.n1374 585
R949 B.n1375 B.n8 585
R950 B.n1373 B.n9 585
R951 B.n12 B.n9 585
R952 B.n1372 B.n1371 585
R953 B.n1371 B.n1370 585
R954 B.n11 B.n10 585
R955 B.n1369 B.n11 585
R956 B.n1367 B.n1366 585
R957 B.n1368 B.n1367 585
R958 B.n1365 B.n16 585
R959 B.n19 B.n16 585
R960 B.n1364 B.n1363 585
R961 B.n1363 B.n1362 585
R962 B.n18 B.n17 585
R963 B.n1361 B.n18 585
R964 B.n1359 B.n1358 585
R965 B.n1360 B.n1359 585
R966 B.n1357 B.n24 585
R967 B.n24 B.n23 585
R968 B.n1356 B.n1355 585
R969 B.n1355 B.n1354 585
R970 B.n26 B.n25 585
R971 B.n1353 B.n26 585
R972 B.n1351 B.n1350 585
R973 B.n1352 B.n1351 585
R974 B.n1349 B.n31 585
R975 B.n31 B.n30 585
R976 B.n1348 B.n1347 585
R977 B.n1347 B.n1346 585
R978 B.n33 B.n32 585
R979 B.n1345 B.n33 585
R980 B.n1343 B.n1342 585
R981 B.n1344 B.n1343 585
R982 B.n1341 B.n37 585
R983 B.n40 B.n37 585
R984 B.n1340 B.n1339 585
R985 B.n1339 B.n1338 585
R986 B.n39 B.n38 585
R987 B.n1337 B.n39 585
R988 B.n1335 B.n1334 585
R989 B.n1336 B.n1335 585
R990 B.n1333 B.n45 585
R991 B.n45 B.n44 585
R992 B.n1332 B.n1331 585
R993 B.n1331 B.n1330 585
R994 B.n47 B.n46 585
R995 B.n1329 B.n47 585
R996 B.n1327 B.n1326 585
R997 B.n1328 B.n1327 585
R998 B.n1325 B.n52 585
R999 B.n52 B.n51 585
R1000 B.n1324 B.n1323 585
R1001 B.n1323 B.n1322 585
R1002 B.n54 B.n53 585
R1003 B.n1321 B.n54 585
R1004 B.n1319 B.n1318 585
R1005 B.n1320 B.n1319 585
R1006 B.n1317 B.n59 585
R1007 B.n59 B.n58 585
R1008 B.n1316 B.n1315 585
R1009 B.n1315 B.n1314 585
R1010 B.n61 B.n60 585
R1011 B.n1313 B.n61 585
R1012 B.n1311 B.n1310 585
R1013 B.n1312 B.n1311 585
R1014 B.n1309 B.n66 585
R1015 B.n66 B.n65 585
R1016 B.n1308 B.n1307 585
R1017 B.n1307 B.n1306 585
R1018 B.n68 B.n67 585
R1019 B.n1305 B.n68 585
R1020 B.n1303 B.n1302 585
R1021 B.n1304 B.n1303 585
R1022 B.n1301 B.n73 585
R1023 B.n73 B.n72 585
R1024 B.n1300 B.n1299 585
R1025 B.n1299 B.n1298 585
R1026 B.n75 B.n74 585
R1027 B.n1297 B.n75 585
R1028 B.n1295 B.n1294 585
R1029 B.n1296 B.n1295 585
R1030 B.n1293 B.n80 585
R1031 B.n80 B.n79 585
R1032 B.n1292 B.n1291 585
R1033 B.n1291 B.n1290 585
R1034 B.n82 B.n81 585
R1035 B.n1289 B.n82 585
R1036 B.n1287 B.n1286 585
R1037 B.n1288 B.n1287 585
R1038 B.n1285 B.n87 585
R1039 B.n87 B.n86 585
R1040 B.n1284 B.n1283 585
R1041 B.n1283 B.n1282 585
R1042 B.n89 B.n88 585
R1043 B.n1281 B.n89 585
R1044 B.n1279 B.n1278 585
R1045 B.n1280 B.n1279 585
R1046 B.n1277 B.n94 585
R1047 B.n94 B.n93 585
R1048 B.n1276 B.n1275 585
R1049 B.n1275 B.n1274 585
R1050 B.n96 B.n95 585
R1051 B.n1273 B.n96 585
R1052 B.n1271 B.n1270 585
R1053 B.n1272 B.n1271 585
R1054 B.n1269 B.n101 585
R1055 B.n101 B.n100 585
R1056 B.n1268 B.n1267 585
R1057 B.n1267 B.n1266 585
R1058 B.n103 B.n102 585
R1059 B.n1265 B.n103 585
R1060 B.n1263 B.n1262 585
R1061 B.n1264 B.n1263 585
R1062 B.n1261 B.n108 585
R1063 B.n108 B.n107 585
R1064 B.n1260 B.n1259 585
R1065 B.n1259 B.n1258 585
R1066 B.n110 B.n109 585
R1067 B.n1257 B.n110 585
R1068 B.n1255 B.n1254 585
R1069 B.n1256 B.n1255 585
R1070 B.n1253 B.n115 585
R1071 B.n115 B.n114 585
R1072 B.n1252 B.n1251 585
R1073 B.n1251 B.n1250 585
R1074 B.n117 B.n116 585
R1075 B.n1249 B.n117 585
R1076 B.n1247 B.n1246 585
R1077 B.n1248 B.n1247 585
R1078 B.n1245 B.n122 585
R1079 B.n122 B.n121 585
R1080 B.n1244 B.n1243 585
R1081 B.n1243 B.n1242 585
R1082 B.n124 B.n123 585
R1083 B.n1241 B.n124 585
R1084 B.n1239 B.n1238 585
R1085 B.n1240 B.n1239 585
R1086 B.n1237 B.n129 585
R1087 B.n129 B.n128 585
R1088 B.n1236 B.n1235 585
R1089 B.n1235 B.n1234 585
R1090 B.n131 B.n130 585
R1091 B.n1233 B.n131 585
R1092 B.n1231 B.n1230 585
R1093 B.n1232 B.n1231 585
R1094 B.n1229 B.n136 585
R1095 B.n136 B.n135 585
R1096 B.n1228 B.n1227 585
R1097 B.n1227 B.n1226 585
R1098 B.n1380 B.n1379 585
R1099 B.n1378 B.n2 585
R1100 B.n1227 B.n138 502.111
R1101 B.n1223 B.n139 502.111
R1102 B.n894 B.n590 502.111
R1103 B.n896 B.n588 502.111
R1104 B.n202 B.t10 321.832
R1105 B.n200 B.t18 321.832
R1106 B.n618 B.t14 321.832
R1107 B.n627 B.t21 321.832
R1108 B.n1225 B.n1224 256.663
R1109 B.n1225 B.n198 256.663
R1110 B.n1225 B.n197 256.663
R1111 B.n1225 B.n196 256.663
R1112 B.n1225 B.n195 256.663
R1113 B.n1225 B.n194 256.663
R1114 B.n1225 B.n193 256.663
R1115 B.n1225 B.n192 256.663
R1116 B.n1225 B.n191 256.663
R1117 B.n1225 B.n190 256.663
R1118 B.n1225 B.n189 256.663
R1119 B.n1225 B.n188 256.663
R1120 B.n1225 B.n187 256.663
R1121 B.n1225 B.n186 256.663
R1122 B.n1225 B.n185 256.663
R1123 B.n1225 B.n184 256.663
R1124 B.n1225 B.n183 256.663
R1125 B.n1225 B.n182 256.663
R1126 B.n1225 B.n181 256.663
R1127 B.n1225 B.n180 256.663
R1128 B.n1225 B.n179 256.663
R1129 B.n1225 B.n178 256.663
R1130 B.n1225 B.n177 256.663
R1131 B.n1225 B.n176 256.663
R1132 B.n1225 B.n175 256.663
R1133 B.n1225 B.n174 256.663
R1134 B.n1225 B.n173 256.663
R1135 B.n1225 B.n172 256.663
R1136 B.n1225 B.n171 256.663
R1137 B.n1225 B.n170 256.663
R1138 B.n1225 B.n169 256.663
R1139 B.n1225 B.n168 256.663
R1140 B.n1225 B.n167 256.663
R1141 B.n1225 B.n166 256.663
R1142 B.n1225 B.n165 256.663
R1143 B.n1225 B.n164 256.663
R1144 B.n1225 B.n163 256.663
R1145 B.n1225 B.n162 256.663
R1146 B.n1225 B.n161 256.663
R1147 B.n1225 B.n160 256.663
R1148 B.n1225 B.n159 256.663
R1149 B.n1225 B.n158 256.663
R1150 B.n1225 B.n157 256.663
R1151 B.n1225 B.n156 256.663
R1152 B.n1225 B.n155 256.663
R1153 B.n1225 B.n154 256.663
R1154 B.n1225 B.n153 256.663
R1155 B.n1225 B.n152 256.663
R1156 B.n1225 B.n151 256.663
R1157 B.n1225 B.n150 256.663
R1158 B.n1225 B.n149 256.663
R1159 B.n1225 B.n148 256.663
R1160 B.n1225 B.n147 256.663
R1161 B.n1225 B.n146 256.663
R1162 B.n1225 B.n145 256.663
R1163 B.n1225 B.n144 256.663
R1164 B.n1225 B.n143 256.663
R1165 B.n1225 B.n142 256.663
R1166 B.n1225 B.n141 256.663
R1167 B.n1225 B.n140 256.663
R1168 B.n655 B.n589 256.663
R1169 B.n661 B.n589 256.663
R1170 B.n663 B.n589 256.663
R1171 B.n669 B.n589 256.663
R1172 B.n671 B.n589 256.663
R1173 B.n677 B.n589 256.663
R1174 B.n679 B.n589 256.663
R1175 B.n685 B.n589 256.663
R1176 B.n687 B.n589 256.663
R1177 B.n693 B.n589 256.663
R1178 B.n695 B.n589 256.663
R1179 B.n701 B.n589 256.663
R1180 B.n703 B.n589 256.663
R1181 B.n709 B.n589 256.663
R1182 B.n711 B.n589 256.663
R1183 B.n717 B.n589 256.663
R1184 B.n719 B.n589 256.663
R1185 B.n725 B.n589 256.663
R1186 B.n727 B.n589 256.663
R1187 B.n733 B.n589 256.663
R1188 B.n735 B.n589 256.663
R1189 B.n741 B.n589 256.663
R1190 B.n743 B.n589 256.663
R1191 B.n749 B.n589 256.663
R1192 B.n751 B.n589 256.663
R1193 B.n757 B.n589 256.663
R1194 B.n759 B.n589 256.663
R1195 B.n766 B.n589 256.663
R1196 B.n768 B.n589 256.663
R1197 B.n774 B.n589 256.663
R1198 B.n776 B.n589 256.663
R1199 B.n782 B.n589 256.663
R1200 B.n784 B.n589 256.663
R1201 B.n790 B.n589 256.663
R1202 B.n792 B.n589 256.663
R1203 B.n798 B.n589 256.663
R1204 B.n800 B.n589 256.663
R1205 B.n806 B.n589 256.663
R1206 B.n808 B.n589 256.663
R1207 B.n814 B.n589 256.663
R1208 B.n816 B.n589 256.663
R1209 B.n822 B.n589 256.663
R1210 B.n824 B.n589 256.663
R1211 B.n830 B.n589 256.663
R1212 B.n832 B.n589 256.663
R1213 B.n838 B.n589 256.663
R1214 B.n840 B.n589 256.663
R1215 B.n846 B.n589 256.663
R1216 B.n848 B.n589 256.663
R1217 B.n854 B.n589 256.663
R1218 B.n856 B.n589 256.663
R1219 B.n862 B.n589 256.663
R1220 B.n864 B.n589 256.663
R1221 B.n870 B.n589 256.663
R1222 B.n872 B.n589 256.663
R1223 B.n878 B.n589 256.663
R1224 B.n880 B.n589 256.663
R1225 B.n886 B.n589 256.663
R1226 B.n889 B.n589 256.663
R1227 B.n1382 B.n1381 256.663
R1228 B.n206 B.n205 163.367
R1229 B.n210 B.n209 163.367
R1230 B.n214 B.n213 163.367
R1231 B.n218 B.n217 163.367
R1232 B.n222 B.n221 163.367
R1233 B.n226 B.n225 163.367
R1234 B.n230 B.n229 163.367
R1235 B.n234 B.n233 163.367
R1236 B.n238 B.n237 163.367
R1237 B.n242 B.n241 163.367
R1238 B.n246 B.n245 163.367
R1239 B.n250 B.n249 163.367
R1240 B.n254 B.n253 163.367
R1241 B.n258 B.n257 163.367
R1242 B.n262 B.n261 163.367
R1243 B.n266 B.n265 163.367
R1244 B.n270 B.n269 163.367
R1245 B.n274 B.n273 163.367
R1246 B.n278 B.n277 163.367
R1247 B.n282 B.n281 163.367
R1248 B.n286 B.n285 163.367
R1249 B.n290 B.n289 163.367
R1250 B.n294 B.n293 163.367
R1251 B.n298 B.n297 163.367
R1252 B.n302 B.n301 163.367
R1253 B.n306 B.n305 163.367
R1254 B.n310 B.n309 163.367
R1255 B.n315 B.n314 163.367
R1256 B.n319 B.n318 163.367
R1257 B.n323 B.n322 163.367
R1258 B.n327 B.n326 163.367
R1259 B.n331 B.n330 163.367
R1260 B.n336 B.n335 163.367
R1261 B.n340 B.n339 163.367
R1262 B.n344 B.n343 163.367
R1263 B.n348 B.n347 163.367
R1264 B.n352 B.n351 163.367
R1265 B.n356 B.n355 163.367
R1266 B.n360 B.n359 163.367
R1267 B.n364 B.n363 163.367
R1268 B.n368 B.n367 163.367
R1269 B.n372 B.n371 163.367
R1270 B.n376 B.n375 163.367
R1271 B.n380 B.n379 163.367
R1272 B.n384 B.n383 163.367
R1273 B.n388 B.n387 163.367
R1274 B.n392 B.n391 163.367
R1275 B.n396 B.n395 163.367
R1276 B.n400 B.n399 163.367
R1277 B.n404 B.n403 163.367
R1278 B.n408 B.n407 163.367
R1279 B.n412 B.n411 163.367
R1280 B.n416 B.n415 163.367
R1281 B.n420 B.n419 163.367
R1282 B.n424 B.n423 163.367
R1283 B.n428 B.n427 163.367
R1284 B.n432 B.n431 163.367
R1285 B.n436 B.n435 163.367
R1286 B.n438 B.n199 163.367
R1287 B.n894 B.n584 163.367
R1288 B.n902 B.n584 163.367
R1289 B.n902 B.n582 163.367
R1290 B.n906 B.n582 163.367
R1291 B.n906 B.n576 163.367
R1292 B.n914 B.n576 163.367
R1293 B.n914 B.n574 163.367
R1294 B.n918 B.n574 163.367
R1295 B.n918 B.n568 163.367
R1296 B.n926 B.n568 163.367
R1297 B.n926 B.n566 163.367
R1298 B.n930 B.n566 163.367
R1299 B.n930 B.n560 163.367
R1300 B.n938 B.n560 163.367
R1301 B.n938 B.n558 163.367
R1302 B.n942 B.n558 163.367
R1303 B.n942 B.n552 163.367
R1304 B.n950 B.n552 163.367
R1305 B.n950 B.n550 163.367
R1306 B.n954 B.n550 163.367
R1307 B.n954 B.n543 163.367
R1308 B.n962 B.n543 163.367
R1309 B.n962 B.n541 163.367
R1310 B.n966 B.n541 163.367
R1311 B.n966 B.n536 163.367
R1312 B.n974 B.n536 163.367
R1313 B.n974 B.n534 163.367
R1314 B.n978 B.n534 163.367
R1315 B.n978 B.n528 163.367
R1316 B.n986 B.n528 163.367
R1317 B.n986 B.n526 163.367
R1318 B.n990 B.n526 163.367
R1319 B.n990 B.n520 163.367
R1320 B.n998 B.n520 163.367
R1321 B.n998 B.n518 163.367
R1322 B.n1002 B.n518 163.367
R1323 B.n1002 B.n512 163.367
R1324 B.n1010 B.n512 163.367
R1325 B.n1010 B.n510 163.367
R1326 B.n1014 B.n510 163.367
R1327 B.n1014 B.n504 163.367
R1328 B.n1022 B.n504 163.367
R1329 B.n1022 B.n502 163.367
R1330 B.n1026 B.n502 163.367
R1331 B.n1026 B.n496 163.367
R1332 B.n1034 B.n496 163.367
R1333 B.n1034 B.n494 163.367
R1334 B.n1038 B.n494 163.367
R1335 B.n1038 B.n488 163.367
R1336 B.n1046 B.n488 163.367
R1337 B.n1046 B.n486 163.367
R1338 B.n1050 B.n486 163.367
R1339 B.n1050 B.n480 163.367
R1340 B.n1058 B.n480 163.367
R1341 B.n1058 B.n478 163.367
R1342 B.n1062 B.n478 163.367
R1343 B.n1062 B.n473 163.367
R1344 B.n1071 B.n473 163.367
R1345 B.n1071 B.n471 163.367
R1346 B.n1075 B.n471 163.367
R1347 B.n1075 B.n465 163.367
R1348 B.n1083 B.n465 163.367
R1349 B.n1083 B.n463 163.367
R1350 B.n1087 B.n463 163.367
R1351 B.n1087 B.n457 163.367
R1352 B.n1095 B.n457 163.367
R1353 B.n1095 B.n455 163.367
R1354 B.n1099 B.n455 163.367
R1355 B.n1099 B.n450 163.367
R1356 B.n1108 B.n450 163.367
R1357 B.n1108 B.n448 163.367
R1358 B.n1113 B.n448 163.367
R1359 B.n1113 B.n442 163.367
R1360 B.n1121 B.n442 163.367
R1361 B.n1122 B.n1121 163.367
R1362 B.n1122 B.n5 163.367
R1363 B.n6 B.n5 163.367
R1364 B.n7 B.n6 163.367
R1365 B.n1128 B.n7 163.367
R1366 B.n1129 B.n1128 163.367
R1367 B.n1129 B.n13 163.367
R1368 B.n14 B.n13 163.367
R1369 B.n15 B.n14 163.367
R1370 B.n1134 B.n15 163.367
R1371 B.n1134 B.n20 163.367
R1372 B.n21 B.n20 163.367
R1373 B.n22 B.n21 163.367
R1374 B.n1139 B.n22 163.367
R1375 B.n1139 B.n27 163.367
R1376 B.n28 B.n27 163.367
R1377 B.n29 B.n28 163.367
R1378 B.n1144 B.n29 163.367
R1379 B.n1144 B.n34 163.367
R1380 B.n35 B.n34 163.367
R1381 B.n36 B.n35 163.367
R1382 B.n1149 B.n36 163.367
R1383 B.n1149 B.n41 163.367
R1384 B.n42 B.n41 163.367
R1385 B.n43 B.n42 163.367
R1386 B.n1154 B.n43 163.367
R1387 B.n1154 B.n48 163.367
R1388 B.n49 B.n48 163.367
R1389 B.n50 B.n49 163.367
R1390 B.n1159 B.n50 163.367
R1391 B.n1159 B.n55 163.367
R1392 B.n56 B.n55 163.367
R1393 B.n57 B.n56 163.367
R1394 B.n1164 B.n57 163.367
R1395 B.n1164 B.n62 163.367
R1396 B.n63 B.n62 163.367
R1397 B.n64 B.n63 163.367
R1398 B.n1169 B.n64 163.367
R1399 B.n1169 B.n69 163.367
R1400 B.n70 B.n69 163.367
R1401 B.n71 B.n70 163.367
R1402 B.n1174 B.n71 163.367
R1403 B.n1174 B.n76 163.367
R1404 B.n77 B.n76 163.367
R1405 B.n78 B.n77 163.367
R1406 B.n1179 B.n78 163.367
R1407 B.n1179 B.n83 163.367
R1408 B.n84 B.n83 163.367
R1409 B.n85 B.n84 163.367
R1410 B.n1184 B.n85 163.367
R1411 B.n1184 B.n90 163.367
R1412 B.n91 B.n90 163.367
R1413 B.n92 B.n91 163.367
R1414 B.n1189 B.n92 163.367
R1415 B.n1189 B.n97 163.367
R1416 B.n98 B.n97 163.367
R1417 B.n99 B.n98 163.367
R1418 B.n1194 B.n99 163.367
R1419 B.n1194 B.n104 163.367
R1420 B.n105 B.n104 163.367
R1421 B.n106 B.n105 163.367
R1422 B.n1199 B.n106 163.367
R1423 B.n1199 B.n111 163.367
R1424 B.n112 B.n111 163.367
R1425 B.n113 B.n112 163.367
R1426 B.n1204 B.n113 163.367
R1427 B.n1204 B.n118 163.367
R1428 B.n119 B.n118 163.367
R1429 B.n120 B.n119 163.367
R1430 B.n1209 B.n120 163.367
R1431 B.n1209 B.n125 163.367
R1432 B.n126 B.n125 163.367
R1433 B.n127 B.n126 163.367
R1434 B.n1214 B.n127 163.367
R1435 B.n1214 B.n132 163.367
R1436 B.n133 B.n132 163.367
R1437 B.n134 B.n133 163.367
R1438 B.n1219 B.n134 163.367
R1439 B.n1219 B.n139 163.367
R1440 B.n656 B.n654 163.367
R1441 B.n660 B.n654 163.367
R1442 B.n664 B.n662 163.367
R1443 B.n668 B.n652 163.367
R1444 B.n672 B.n670 163.367
R1445 B.n676 B.n650 163.367
R1446 B.n680 B.n678 163.367
R1447 B.n684 B.n648 163.367
R1448 B.n688 B.n686 163.367
R1449 B.n692 B.n646 163.367
R1450 B.n696 B.n694 163.367
R1451 B.n700 B.n644 163.367
R1452 B.n704 B.n702 163.367
R1453 B.n708 B.n642 163.367
R1454 B.n712 B.n710 163.367
R1455 B.n716 B.n640 163.367
R1456 B.n720 B.n718 163.367
R1457 B.n724 B.n638 163.367
R1458 B.n728 B.n726 163.367
R1459 B.n732 B.n636 163.367
R1460 B.n736 B.n734 163.367
R1461 B.n740 B.n634 163.367
R1462 B.n744 B.n742 163.367
R1463 B.n748 B.n632 163.367
R1464 B.n752 B.n750 163.367
R1465 B.n756 B.n630 163.367
R1466 B.n760 B.n758 163.367
R1467 B.n765 B.n626 163.367
R1468 B.n769 B.n767 163.367
R1469 B.n773 B.n624 163.367
R1470 B.n777 B.n775 163.367
R1471 B.n781 B.n622 163.367
R1472 B.n785 B.n783 163.367
R1473 B.n789 B.n617 163.367
R1474 B.n793 B.n791 163.367
R1475 B.n797 B.n615 163.367
R1476 B.n801 B.n799 163.367
R1477 B.n805 B.n613 163.367
R1478 B.n809 B.n807 163.367
R1479 B.n813 B.n611 163.367
R1480 B.n817 B.n815 163.367
R1481 B.n821 B.n609 163.367
R1482 B.n825 B.n823 163.367
R1483 B.n829 B.n607 163.367
R1484 B.n833 B.n831 163.367
R1485 B.n837 B.n605 163.367
R1486 B.n841 B.n839 163.367
R1487 B.n845 B.n603 163.367
R1488 B.n849 B.n847 163.367
R1489 B.n853 B.n601 163.367
R1490 B.n857 B.n855 163.367
R1491 B.n861 B.n599 163.367
R1492 B.n865 B.n863 163.367
R1493 B.n869 B.n597 163.367
R1494 B.n873 B.n871 163.367
R1495 B.n877 B.n595 163.367
R1496 B.n881 B.n879 163.367
R1497 B.n885 B.n593 163.367
R1498 B.n888 B.n887 163.367
R1499 B.n890 B.n590 163.367
R1500 B.n896 B.n586 163.367
R1501 B.n900 B.n586 163.367
R1502 B.n900 B.n580 163.367
R1503 B.n908 B.n580 163.367
R1504 B.n908 B.n578 163.367
R1505 B.n912 B.n578 163.367
R1506 B.n912 B.n572 163.367
R1507 B.n920 B.n572 163.367
R1508 B.n920 B.n570 163.367
R1509 B.n924 B.n570 163.367
R1510 B.n924 B.n564 163.367
R1511 B.n932 B.n564 163.367
R1512 B.n932 B.n562 163.367
R1513 B.n936 B.n562 163.367
R1514 B.n936 B.n556 163.367
R1515 B.n944 B.n556 163.367
R1516 B.n944 B.n554 163.367
R1517 B.n948 B.n554 163.367
R1518 B.n948 B.n548 163.367
R1519 B.n956 B.n548 163.367
R1520 B.n956 B.n546 163.367
R1521 B.n960 B.n546 163.367
R1522 B.n960 B.n540 163.367
R1523 B.n968 B.n540 163.367
R1524 B.n968 B.n538 163.367
R1525 B.n972 B.n538 163.367
R1526 B.n972 B.n532 163.367
R1527 B.n980 B.n532 163.367
R1528 B.n980 B.n530 163.367
R1529 B.n984 B.n530 163.367
R1530 B.n984 B.n524 163.367
R1531 B.n992 B.n524 163.367
R1532 B.n992 B.n522 163.367
R1533 B.n996 B.n522 163.367
R1534 B.n996 B.n516 163.367
R1535 B.n1004 B.n516 163.367
R1536 B.n1004 B.n514 163.367
R1537 B.n1008 B.n514 163.367
R1538 B.n1008 B.n508 163.367
R1539 B.n1016 B.n508 163.367
R1540 B.n1016 B.n506 163.367
R1541 B.n1020 B.n506 163.367
R1542 B.n1020 B.n500 163.367
R1543 B.n1028 B.n500 163.367
R1544 B.n1028 B.n498 163.367
R1545 B.n1032 B.n498 163.367
R1546 B.n1032 B.n492 163.367
R1547 B.n1040 B.n492 163.367
R1548 B.n1040 B.n490 163.367
R1549 B.n1044 B.n490 163.367
R1550 B.n1044 B.n484 163.367
R1551 B.n1052 B.n484 163.367
R1552 B.n1052 B.n482 163.367
R1553 B.n1056 B.n482 163.367
R1554 B.n1056 B.n476 163.367
R1555 B.n1065 B.n476 163.367
R1556 B.n1065 B.n474 163.367
R1557 B.n1069 B.n474 163.367
R1558 B.n1069 B.n469 163.367
R1559 B.n1077 B.n469 163.367
R1560 B.n1077 B.n467 163.367
R1561 B.n1081 B.n467 163.367
R1562 B.n1081 B.n461 163.367
R1563 B.n1089 B.n461 163.367
R1564 B.n1089 B.n459 163.367
R1565 B.n1093 B.n459 163.367
R1566 B.n1093 B.n453 163.367
R1567 B.n1102 B.n453 163.367
R1568 B.n1102 B.n451 163.367
R1569 B.n1106 B.n451 163.367
R1570 B.n1106 B.n446 163.367
R1571 B.n1115 B.n446 163.367
R1572 B.n1115 B.n444 163.367
R1573 B.n1119 B.n444 163.367
R1574 B.n1119 B.n3 163.367
R1575 B.n1380 B.n3 163.367
R1576 B.n1376 B.n2 163.367
R1577 B.n1376 B.n1375 163.367
R1578 B.n1375 B.n9 163.367
R1579 B.n1371 B.n9 163.367
R1580 B.n1371 B.n11 163.367
R1581 B.n1367 B.n11 163.367
R1582 B.n1367 B.n16 163.367
R1583 B.n1363 B.n16 163.367
R1584 B.n1363 B.n18 163.367
R1585 B.n1359 B.n18 163.367
R1586 B.n1359 B.n24 163.367
R1587 B.n1355 B.n24 163.367
R1588 B.n1355 B.n26 163.367
R1589 B.n1351 B.n26 163.367
R1590 B.n1351 B.n31 163.367
R1591 B.n1347 B.n31 163.367
R1592 B.n1347 B.n33 163.367
R1593 B.n1343 B.n33 163.367
R1594 B.n1343 B.n37 163.367
R1595 B.n1339 B.n37 163.367
R1596 B.n1339 B.n39 163.367
R1597 B.n1335 B.n39 163.367
R1598 B.n1335 B.n45 163.367
R1599 B.n1331 B.n45 163.367
R1600 B.n1331 B.n47 163.367
R1601 B.n1327 B.n47 163.367
R1602 B.n1327 B.n52 163.367
R1603 B.n1323 B.n52 163.367
R1604 B.n1323 B.n54 163.367
R1605 B.n1319 B.n54 163.367
R1606 B.n1319 B.n59 163.367
R1607 B.n1315 B.n59 163.367
R1608 B.n1315 B.n61 163.367
R1609 B.n1311 B.n61 163.367
R1610 B.n1311 B.n66 163.367
R1611 B.n1307 B.n66 163.367
R1612 B.n1307 B.n68 163.367
R1613 B.n1303 B.n68 163.367
R1614 B.n1303 B.n73 163.367
R1615 B.n1299 B.n73 163.367
R1616 B.n1299 B.n75 163.367
R1617 B.n1295 B.n75 163.367
R1618 B.n1295 B.n80 163.367
R1619 B.n1291 B.n80 163.367
R1620 B.n1291 B.n82 163.367
R1621 B.n1287 B.n82 163.367
R1622 B.n1287 B.n87 163.367
R1623 B.n1283 B.n87 163.367
R1624 B.n1283 B.n89 163.367
R1625 B.n1279 B.n89 163.367
R1626 B.n1279 B.n94 163.367
R1627 B.n1275 B.n94 163.367
R1628 B.n1275 B.n96 163.367
R1629 B.n1271 B.n96 163.367
R1630 B.n1271 B.n101 163.367
R1631 B.n1267 B.n101 163.367
R1632 B.n1267 B.n103 163.367
R1633 B.n1263 B.n103 163.367
R1634 B.n1263 B.n108 163.367
R1635 B.n1259 B.n108 163.367
R1636 B.n1259 B.n110 163.367
R1637 B.n1255 B.n110 163.367
R1638 B.n1255 B.n115 163.367
R1639 B.n1251 B.n115 163.367
R1640 B.n1251 B.n117 163.367
R1641 B.n1247 B.n117 163.367
R1642 B.n1247 B.n122 163.367
R1643 B.n1243 B.n122 163.367
R1644 B.n1243 B.n124 163.367
R1645 B.n1239 B.n124 163.367
R1646 B.n1239 B.n129 163.367
R1647 B.n1235 B.n129 163.367
R1648 B.n1235 B.n131 163.367
R1649 B.n1231 B.n131 163.367
R1650 B.n1231 B.n136 163.367
R1651 B.n1227 B.n136 163.367
R1652 B.n200 B.t19 148.018
R1653 B.n618 B.t17 148.018
R1654 B.n202 B.t12 147.996
R1655 B.n627 B.t23 147.996
R1656 B.n203 B.n202 75.249
R1657 B.n201 B.n200 75.249
R1658 B.n619 B.n618 75.249
R1659 B.n628 B.n627 75.249
R1660 B.n201 B.t20 72.7695
R1661 B.n619 B.t16 72.7695
R1662 B.n203 B.t13 72.7477
R1663 B.n628 B.t22 72.7477
R1664 B.n140 B.n138 71.676
R1665 B.n206 B.n141 71.676
R1666 B.n210 B.n142 71.676
R1667 B.n214 B.n143 71.676
R1668 B.n218 B.n144 71.676
R1669 B.n222 B.n145 71.676
R1670 B.n226 B.n146 71.676
R1671 B.n230 B.n147 71.676
R1672 B.n234 B.n148 71.676
R1673 B.n238 B.n149 71.676
R1674 B.n242 B.n150 71.676
R1675 B.n246 B.n151 71.676
R1676 B.n250 B.n152 71.676
R1677 B.n254 B.n153 71.676
R1678 B.n258 B.n154 71.676
R1679 B.n262 B.n155 71.676
R1680 B.n266 B.n156 71.676
R1681 B.n270 B.n157 71.676
R1682 B.n274 B.n158 71.676
R1683 B.n278 B.n159 71.676
R1684 B.n282 B.n160 71.676
R1685 B.n286 B.n161 71.676
R1686 B.n290 B.n162 71.676
R1687 B.n294 B.n163 71.676
R1688 B.n298 B.n164 71.676
R1689 B.n302 B.n165 71.676
R1690 B.n306 B.n166 71.676
R1691 B.n310 B.n167 71.676
R1692 B.n315 B.n168 71.676
R1693 B.n319 B.n169 71.676
R1694 B.n323 B.n170 71.676
R1695 B.n327 B.n171 71.676
R1696 B.n331 B.n172 71.676
R1697 B.n336 B.n173 71.676
R1698 B.n340 B.n174 71.676
R1699 B.n344 B.n175 71.676
R1700 B.n348 B.n176 71.676
R1701 B.n352 B.n177 71.676
R1702 B.n356 B.n178 71.676
R1703 B.n360 B.n179 71.676
R1704 B.n364 B.n180 71.676
R1705 B.n368 B.n181 71.676
R1706 B.n372 B.n182 71.676
R1707 B.n376 B.n183 71.676
R1708 B.n380 B.n184 71.676
R1709 B.n384 B.n185 71.676
R1710 B.n388 B.n186 71.676
R1711 B.n392 B.n187 71.676
R1712 B.n396 B.n188 71.676
R1713 B.n400 B.n189 71.676
R1714 B.n404 B.n190 71.676
R1715 B.n408 B.n191 71.676
R1716 B.n412 B.n192 71.676
R1717 B.n416 B.n193 71.676
R1718 B.n420 B.n194 71.676
R1719 B.n424 B.n195 71.676
R1720 B.n428 B.n196 71.676
R1721 B.n432 B.n197 71.676
R1722 B.n436 B.n198 71.676
R1723 B.n1224 B.n199 71.676
R1724 B.n1224 B.n1223 71.676
R1725 B.n438 B.n198 71.676
R1726 B.n435 B.n197 71.676
R1727 B.n431 B.n196 71.676
R1728 B.n427 B.n195 71.676
R1729 B.n423 B.n194 71.676
R1730 B.n419 B.n193 71.676
R1731 B.n415 B.n192 71.676
R1732 B.n411 B.n191 71.676
R1733 B.n407 B.n190 71.676
R1734 B.n403 B.n189 71.676
R1735 B.n399 B.n188 71.676
R1736 B.n395 B.n187 71.676
R1737 B.n391 B.n186 71.676
R1738 B.n387 B.n185 71.676
R1739 B.n383 B.n184 71.676
R1740 B.n379 B.n183 71.676
R1741 B.n375 B.n182 71.676
R1742 B.n371 B.n181 71.676
R1743 B.n367 B.n180 71.676
R1744 B.n363 B.n179 71.676
R1745 B.n359 B.n178 71.676
R1746 B.n355 B.n177 71.676
R1747 B.n351 B.n176 71.676
R1748 B.n347 B.n175 71.676
R1749 B.n343 B.n174 71.676
R1750 B.n339 B.n173 71.676
R1751 B.n335 B.n172 71.676
R1752 B.n330 B.n171 71.676
R1753 B.n326 B.n170 71.676
R1754 B.n322 B.n169 71.676
R1755 B.n318 B.n168 71.676
R1756 B.n314 B.n167 71.676
R1757 B.n309 B.n166 71.676
R1758 B.n305 B.n165 71.676
R1759 B.n301 B.n164 71.676
R1760 B.n297 B.n163 71.676
R1761 B.n293 B.n162 71.676
R1762 B.n289 B.n161 71.676
R1763 B.n285 B.n160 71.676
R1764 B.n281 B.n159 71.676
R1765 B.n277 B.n158 71.676
R1766 B.n273 B.n157 71.676
R1767 B.n269 B.n156 71.676
R1768 B.n265 B.n155 71.676
R1769 B.n261 B.n154 71.676
R1770 B.n257 B.n153 71.676
R1771 B.n253 B.n152 71.676
R1772 B.n249 B.n151 71.676
R1773 B.n245 B.n150 71.676
R1774 B.n241 B.n149 71.676
R1775 B.n237 B.n148 71.676
R1776 B.n233 B.n147 71.676
R1777 B.n229 B.n146 71.676
R1778 B.n225 B.n145 71.676
R1779 B.n221 B.n144 71.676
R1780 B.n217 B.n143 71.676
R1781 B.n213 B.n142 71.676
R1782 B.n209 B.n141 71.676
R1783 B.n205 B.n140 71.676
R1784 B.n655 B.n588 71.676
R1785 B.n661 B.n660 71.676
R1786 B.n664 B.n663 71.676
R1787 B.n669 B.n668 71.676
R1788 B.n672 B.n671 71.676
R1789 B.n677 B.n676 71.676
R1790 B.n680 B.n679 71.676
R1791 B.n685 B.n684 71.676
R1792 B.n688 B.n687 71.676
R1793 B.n693 B.n692 71.676
R1794 B.n696 B.n695 71.676
R1795 B.n701 B.n700 71.676
R1796 B.n704 B.n703 71.676
R1797 B.n709 B.n708 71.676
R1798 B.n712 B.n711 71.676
R1799 B.n717 B.n716 71.676
R1800 B.n720 B.n719 71.676
R1801 B.n725 B.n724 71.676
R1802 B.n728 B.n727 71.676
R1803 B.n733 B.n732 71.676
R1804 B.n736 B.n735 71.676
R1805 B.n741 B.n740 71.676
R1806 B.n744 B.n743 71.676
R1807 B.n749 B.n748 71.676
R1808 B.n752 B.n751 71.676
R1809 B.n757 B.n756 71.676
R1810 B.n760 B.n759 71.676
R1811 B.n766 B.n765 71.676
R1812 B.n769 B.n768 71.676
R1813 B.n774 B.n773 71.676
R1814 B.n777 B.n776 71.676
R1815 B.n782 B.n781 71.676
R1816 B.n785 B.n784 71.676
R1817 B.n790 B.n789 71.676
R1818 B.n793 B.n792 71.676
R1819 B.n798 B.n797 71.676
R1820 B.n801 B.n800 71.676
R1821 B.n806 B.n805 71.676
R1822 B.n809 B.n808 71.676
R1823 B.n814 B.n813 71.676
R1824 B.n817 B.n816 71.676
R1825 B.n822 B.n821 71.676
R1826 B.n825 B.n824 71.676
R1827 B.n830 B.n829 71.676
R1828 B.n833 B.n832 71.676
R1829 B.n838 B.n837 71.676
R1830 B.n841 B.n840 71.676
R1831 B.n846 B.n845 71.676
R1832 B.n849 B.n848 71.676
R1833 B.n854 B.n853 71.676
R1834 B.n857 B.n856 71.676
R1835 B.n862 B.n861 71.676
R1836 B.n865 B.n864 71.676
R1837 B.n870 B.n869 71.676
R1838 B.n873 B.n872 71.676
R1839 B.n878 B.n877 71.676
R1840 B.n881 B.n880 71.676
R1841 B.n886 B.n885 71.676
R1842 B.n889 B.n888 71.676
R1843 B.n656 B.n655 71.676
R1844 B.n662 B.n661 71.676
R1845 B.n663 B.n652 71.676
R1846 B.n670 B.n669 71.676
R1847 B.n671 B.n650 71.676
R1848 B.n678 B.n677 71.676
R1849 B.n679 B.n648 71.676
R1850 B.n686 B.n685 71.676
R1851 B.n687 B.n646 71.676
R1852 B.n694 B.n693 71.676
R1853 B.n695 B.n644 71.676
R1854 B.n702 B.n701 71.676
R1855 B.n703 B.n642 71.676
R1856 B.n710 B.n709 71.676
R1857 B.n711 B.n640 71.676
R1858 B.n718 B.n717 71.676
R1859 B.n719 B.n638 71.676
R1860 B.n726 B.n725 71.676
R1861 B.n727 B.n636 71.676
R1862 B.n734 B.n733 71.676
R1863 B.n735 B.n634 71.676
R1864 B.n742 B.n741 71.676
R1865 B.n743 B.n632 71.676
R1866 B.n750 B.n749 71.676
R1867 B.n751 B.n630 71.676
R1868 B.n758 B.n757 71.676
R1869 B.n759 B.n626 71.676
R1870 B.n767 B.n766 71.676
R1871 B.n768 B.n624 71.676
R1872 B.n775 B.n774 71.676
R1873 B.n776 B.n622 71.676
R1874 B.n783 B.n782 71.676
R1875 B.n784 B.n617 71.676
R1876 B.n791 B.n790 71.676
R1877 B.n792 B.n615 71.676
R1878 B.n799 B.n798 71.676
R1879 B.n800 B.n613 71.676
R1880 B.n807 B.n806 71.676
R1881 B.n808 B.n611 71.676
R1882 B.n815 B.n814 71.676
R1883 B.n816 B.n609 71.676
R1884 B.n823 B.n822 71.676
R1885 B.n824 B.n607 71.676
R1886 B.n831 B.n830 71.676
R1887 B.n832 B.n605 71.676
R1888 B.n839 B.n838 71.676
R1889 B.n840 B.n603 71.676
R1890 B.n847 B.n846 71.676
R1891 B.n848 B.n601 71.676
R1892 B.n855 B.n854 71.676
R1893 B.n856 B.n599 71.676
R1894 B.n863 B.n862 71.676
R1895 B.n864 B.n597 71.676
R1896 B.n871 B.n870 71.676
R1897 B.n872 B.n595 71.676
R1898 B.n879 B.n878 71.676
R1899 B.n880 B.n593 71.676
R1900 B.n887 B.n886 71.676
R1901 B.n890 B.n889 71.676
R1902 B.n1381 B.n1380 71.676
R1903 B.n1381 B.n2 71.676
R1904 B.n895 B.n589 64.8691
R1905 B.n1226 B.n1225 64.8691
R1906 B.n312 B.n203 59.5399
R1907 B.n333 B.n201 59.5399
R1908 B.n620 B.n619 59.5399
R1909 B.n763 B.n628 59.5399
R1910 B.n895 B.n585 34.1948
R1911 B.n901 B.n585 34.1948
R1912 B.n901 B.n581 34.1948
R1913 B.n907 B.n581 34.1948
R1914 B.n907 B.n577 34.1948
R1915 B.n913 B.n577 34.1948
R1916 B.n913 B.n573 34.1948
R1917 B.n919 B.n573 34.1948
R1918 B.n925 B.n569 34.1948
R1919 B.n925 B.n565 34.1948
R1920 B.n931 B.n565 34.1948
R1921 B.n931 B.n561 34.1948
R1922 B.n937 B.n561 34.1948
R1923 B.n937 B.n557 34.1948
R1924 B.n943 B.n557 34.1948
R1925 B.n943 B.n553 34.1948
R1926 B.n949 B.n553 34.1948
R1927 B.n949 B.n549 34.1948
R1928 B.n955 B.n549 34.1948
R1929 B.n955 B.n544 34.1948
R1930 B.n961 B.n544 34.1948
R1931 B.n961 B.n545 34.1948
R1932 B.n967 B.n537 34.1948
R1933 B.n973 B.n537 34.1948
R1934 B.n973 B.n533 34.1948
R1935 B.n979 B.n533 34.1948
R1936 B.n979 B.n529 34.1948
R1937 B.n985 B.n529 34.1948
R1938 B.n985 B.n525 34.1948
R1939 B.n991 B.n525 34.1948
R1940 B.n991 B.n521 34.1948
R1941 B.n997 B.n521 34.1948
R1942 B.n1003 B.n517 34.1948
R1943 B.n1003 B.n513 34.1948
R1944 B.n1009 B.n513 34.1948
R1945 B.n1009 B.n509 34.1948
R1946 B.n1015 B.n509 34.1948
R1947 B.n1015 B.n505 34.1948
R1948 B.n1021 B.n505 34.1948
R1949 B.n1021 B.n501 34.1948
R1950 B.n1027 B.n501 34.1948
R1951 B.n1027 B.n497 34.1948
R1952 B.n1033 B.n497 34.1948
R1953 B.n1039 B.n493 34.1948
R1954 B.n1039 B.n489 34.1948
R1955 B.n1045 B.n489 34.1948
R1956 B.n1045 B.n485 34.1948
R1957 B.n1051 B.n485 34.1948
R1958 B.n1051 B.n481 34.1948
R1959 B.n1057 B.n481 34.1948
R1960 B.n1057 B.n477 34.1948
R1961 B.n1064 B.n477 34.1948
R1962 B.n1064 B.n1063 34.1948
R1963 B.n1070 B.n470 34.1948
R1964 B.n1076 B.n470 34.1948
R1965 B.n1076 B.n466 34.1948
R1966 B.n1082 B.n466 34.1948
R1967 B.n1082 B.n462 34.1948
R1968 B.n1088 B.n462 34.1948
R1969 B.n1088 B.n458 34.1948
R1970 B.n1094 B.n458 34.1948
R1971 B.n1094 B.n454 34.1948
R1972 B.n1101 B.n454 34.1948
R1973 B.n1101 B.n1100 34.1948
R1974 B.n1107 B.n447 34.1948
R1975 B.n1114 B.n447 34.1948
R1976 B.n1114 B.n443 34.1948
R1977 B.n1120 B.n443 34.1948
R1978 B.n1120 B.n4 34.1948
R1979 B.n1379 B.n4 34.1948
R1980 B.n1379 B.n1378 34.1948
R1981 B.n1378 B.n1377 34.1948
R1982 B.n1377 B.n8 34.1948
R1983 B.n12 B.n8 34.1948
R1984 B.n1370 B.n12 34.1948
R1985 B.n1370 B.n1369 34.1948
R1986 B.n1369 B.n1368 34.1948
R1987 B.n1362 B.n19 34.1948
R1988 B.n1362 B.n1361 34.1948
R1989 B.n1361 B.n1360 34.1948
R1990 B.n1360 B.n23 34.1948
R1991 B.n1354 B.n23 34.1948
R1992 B.n1354 B.n1353 34.1948
R1993 B.n1353 B.n1352 34.1948
R1994 B.n1352 B.n30 34.1948
R1995 B.n1346 B.n30 34.1948
R1996 B.n1346 B.n1345 34.1948
R1997 B.n1345 B.n1344 34.1948
R1998 B.n1338 B.n40 34.1948
R1999 B.n1338 B.n1337 34.1948
R2000 B.n1337 B.n1336 34.1948
R2001 B.n1336 B.n44 34.1948
R2002 B.n1330 B.n44 34.1948
R2003 B.n1330 B.n1329 34.1948
R2004 B.n1329 B.n1328 34.1948
R2005 B.n1328 B.n51 34.1948
R2006 B.n1322 B.n51 34.1948
R2007 B.n1322 B.n1321 34.1948
R2008 B.n1320 B.n58 34.1948
R2009 B.n1314 B.n58 34.1948
R2010 B.n1314 B.n1313 34.1948
R2011 B.n1313 B.n1312 34.1948
R2012 B.n1312 B.n65 34.1948
R2013 B.n1306 B.n65 34.1948
R2014 B.n1306 B.n1305 34.1948
R2015 B.n1305 B.n1304 34.1948
R2016 B.n1304 B.n72 34.1948
R2017 B.n1298 B.n72 34.1948
R2018 B.n1298 B.n1297 34.1948
R2019 B.n1296 B.n79 34.1948
R2020 B.n1290 B.n79 34.1948
R2021 B.n1290 B.n1289 34.1948
R2022 B.n1289 B.n1288 34.1948
R2023 B.n1288 B.n86 34.1948
R2024 B.n1282 B.n86 34.1948
R2025 B.n1282 B.n1281 34.1948
R2026 B.n1281 B.n1280 34.1948
R2027 B.n1280 B.n93 34.1948
R2028 B.n1274 B.n93 34.1948
R2029 B.n1273 B.n1272 34.1948
R2030 B.n1272 B.n100 34.1948
R2031 B.n1266 B.n100 34.1948
R2032 B.n1266 B.n1265 34.1948
R2033 B.n1265 B.n1264 34.1948
R2034 B.n1264 B.n107 34.1948
R2035 B.n1258 B.n107 34.1948
R2036 B.n1258 B.n1257 34.1948
R2037 B.n1257 B.n1256 34.1948
R2038 B.n1256 B.n114 34.1948
R2039 B.n1250 B.n114 34.1948
R2040 B.n1250 B.n1249 34.1948
R2041 B.n1249 B.n1248 34.1948
R2042 B.n1248 B.n121 34.1948
R2043 B.n1242 B.n1241 34.1948
R2044 B.n1241 B.n1240 34.1948
R2045 B.n1240 B.n128 34.1948
R2046 B.n1234 B.n128 34.1948
R2047 B.n1234 B.n1233 34.1948
R2048 B.n1233 B.n1232 34.1948
R2049 B.n1232 B.n135 34.1948
R2050 B.n1226 B.n135 34.1948
R2051 B.n997 B.t2 32.6862
R2052 B.t8 B.n1296 32.6862
R2053 B.n897 B.n587 32.6249
R2054 B.n893 B.n892 32.6249
R2055 B.n1222 B.n1221 32.6249
R2056 B.n1228 B.n137 32.6249
R2057 B.n919 B.t15 31.6805
R2058 B.n1242 B.t11 31.6805
R2059 B.n1107 B.t1 27.6576
R2060 B.n1368 B.t6 27.6576
R2061 B.n1063 B.t9 26.6519
R2062 B.n40 B.t3 26.6519
R2063 B.t4 B.n493 21.6234
R2064 B.n1321 B.t5 21.6234
R2065 B.n545 B.t0 18.6062
R2066 B.t7 B.n1273 18.6062
R2067 B B.n1382 18.0485
R2068 B.n967 B.t0 15.5891
R2069 B.n1274 B.t7 15.5891
R2070 B.n1033 B.t4 12.5719
R2071 B.t5 B.n1320 12.5719
R2072 B.n898 B.n897 10.6151
R2073 B.n899 B.n898 10.6151
R2074 B.n899 B.n579 10.6151
R2075 B.n909 B.n579 10.6151
R2076 B.n910 B.n909 10.6151
R2077 B.n911 B.n910 10.6151
R2078 B.n911 B.n571 10.6151
R2079 B.n921 B.n571 10.6151
R2080 B.n922 B.n921 10.6151
R2081 B.n923 B.n922 10.6151
R2082 B.n923 B.n563 10.6151
R2083 B.n933 B.n563 10.6151
R2084 B.n934 B.n933 10.6151
R2085 B.n935 B.n934 10.6151
R2086 B.n935 B.n555 10.6151
R2087 B.n945 B.n555 10.6151
R2088 B.n946 B.n945 10.6151
R2089 B.n947 B.n946 10.6151
R2090 B.n947 B.n547 10.6151
R2091 B.n957 B.n547 10.6151
R2092 B.n958 B.n957 10.6151
R2093 B.n959 B.n958 10.6151
R2094 B.n959 B.n539 10.6151
R2095 B.n969 B.n539 10.6151
R2096 B.n970 B.n969 10.6151
R2097 B.n971 B.n970 10.6151
R2098 B.n971 B.n531 10.6151
R2099 B.n981 B.n531 10.6151
R2100 B.n982 B.n981 10.6151
R2101 B.n983 B.n982 10.6151
R2102 B.n983 B.n523 10.6151
R2103 B.n993 B.n523 10.6151
R2104 B.n994 B.n993 10.6151
R2105 B.n995 B.n994 10.6151
R2106 B.n995 B.n515 10.6151
R2107 B.n1005 B.n515 10.6151
R2108 B.n1006 B.n1005 10.6151
R2109 B.n1007 B.n1006 10.6151
R2110 B.n1007 B.n507 10.6151
R2111 B.n1017 B.n507 10.6151
R2112 B.n1018 B.n1017 10.6151
R2113 B.n1019 B.n1018 10.6151
R2114 B.n1019 B.n499 10.6151
R2115 B.n1029 B.n499 10.6151
R2116 B.n1030 B.n1029 10.6151
R2117 B.n1031 B.n1030 10.6151
R2118 B.n1031 B.n491 10.6151
R2119 B.n1041 B.n491 10.6151
R2120 B.n1042 B.n1041 10.6151
R2121 B.n1043 B.n1042 10.6151
R2122 B.n1043 B.n483 10.6151
R2123 B.n1053 B.n483 10.6151
R2124 B.n1054 B.n1053 10.6151
R2125 B.n1055 B.n1054 10.6151
R2126 B.n1055 B.n475 10.6151
R2127 B.n1066 B.n475 10.6151
R2128 B.n1067 B.n1066 10.6151
R2129 B.n1068 B.n1067 10.6151
R2130 B.n1068 B.n468 10.6151
R2131 B.n1078 B.n468 10.6151
R2132 B.n1079 B.n1078 10.6151
R2133 B.n1080 B.n1079 10.6151
R2134 B.n1080 B.n460 10.6151
R2135 B.n1090 B.n460 10.6151
R2136 B.n1091 B.n1090 10.6151
R2137 B.n1092 B.n1091 10.6151
R2138 B.n1092 B.n452 10.6151
R2139 B.n1103 B.n452 10.6151
R2140 B.n1104 B.n1103 10.6151
R2141 B.n1105 B.n1104 10.6151
R2142 B.n1105 B.n445 10.6151
R2143 B.n1116 B.n445 10.6151
R2144 B.n1117 B.n1116 10.6151
R2145 B.n1118 B.n1117 10.6151
R2146 B.n1118 B.n0 10.6151
R2147 B.n657 B.n587 10.6151
R2148 B.n658 B.n657 10.6151
R2149 B.n659 B.n658 10.6151
R2150 B.n659 B.n653 10.6151
R2151 B.n665 B.n653 10.6151
R2152 B.n666 B.n665 10.6151
R2153 B.n667 B.n666 10.6151
R2154 B.n667 B.n651 10.6151
R2155 B.n673 B.n651 10.6151
R2156 B.n674 B.n673 10.6151
R2157 B.n675 B.n674 10.6151
R2158 B.n675 B.n649 10.6151
R2159 B.n681 B.n649 10.6151
R2160 B.n682 B.n681 10.6151
R2161 B.n683 B.n682 10.6151
R2162 B.n683 B.n647 10.6151
R2163 B.n689 B.n647 10.6151
R2164 B.n690 B.n689 10.6151
R2165 B.n691 B.n690 10.6151
R2166 B.n691 B.n645 10.6151
R2167 B.n697 B.n645 10.6151
R2168 B.n698 B.n697 10.6151
R2169 B.n699 B.n698 10.6151
R2170 B.n699 B.n643 10.6151
R2171 B.n705 B.n643 10.6151
R2172 B.n706 B.n705 10.6151
R2173 B.n707 B.n706 10.6151
R2174 B.n707 B.n641 10.6151
R2175 B.n713 B.n641 10.6151
R2176 B.n714 B.n713 10.6151
R2177 B.n715 B.n714 10.6151
R2178 B.n715 B.n639 10.6151
R2179 B.n721 B.n639 10.6151
R2180 B.n722 B.n721 10.6151
R2181 B.n723 B.n722 10.6151
R2182 B.n723 B.n637 10.6151
R2183 B.n729 B.n637 10.6151
R2184 B.n730 B.n729 10.6151
R2185 B.n731 B.n730 10.6151
R2186 B.n731 B.n635 10.6151
R2187 B.n737 B.n635 10.6151
R2188 B.n738 B.n737 10.6151
R2189 B.n739 B.n738 10.6151
R2190 B.n739 B.n633 10.6151
R2191 B.n745 B.n633 10.6151
R2192 B.n746 B.n745 10.6151
R2193 B.n747 B.n746 10.6151
R2194 B.n747 B.n631 10.6151
R2195 B.n753 B.n631 10.6151
R2196 B.n754 B.n753 10.6151
R2197 B.n755 B.n754 10.6151
R2198 B.n755 B.n629 10.6151
R2199 B.n761 B.n629 10.6151
R2200 B.n762 B.n761 10.6151
R2201 B.n764 B.n625 10.6151
R2202 B.n770 B.n625 10.6151
R2203 B.n771 B.n770 10.6151
R2204 B.n772 B.n771 10.6151
R2205 B.n772 B.n623 10.6151
R2206 B.n778 B.n623 10.6151
R2207 B.n779 B.n778 10.6151
R2208 B.n780 B.n779 10.6151
R2209 B.n780 B.n621 10.6151
R2210 B.n787 B.n786 10.6151
R2211 B.n788 B.n787 10.6151
R2212 B.n788 B.n616 10.6151
R2213 B.n794 B.n616 10.6151
R2214 B.n795 B.n794 10.6151
R2215 B.n796 B.n795 10.6151
R2216 B.n796 B.n614 10.6151
R2217 B.n802 B.n614 10.6151
R2218 B.n803 B.n802 10.6151
R2219 B.n804 B.n803 10.6151
R2220 B.n804 B.n612 10.6151
R2221 B.n810 B.n612 10.6151
R2222 B.n811 B.n810 10.6151
R2223 B.n812 B.n811 10.6151
R2224 B.n812 B.n610 10.6151
R2225 B.n818 B.n610 10.6151
R2226 B.n819 B.n818 10.6151
R2227 B.n820 B.n819 10.6151
R2228 B.n820 B.n608 10.6151
R2229 B.n826 B.n608 10.6151
R2230 B.n827 B.n826 10.6151
R2231 B.n828 B.n827 10.6151
R2232 B.n828 B.n606 10.6151
R2233 B.n834 B.n606 10.6151
R2234 B.n835 B.n834 10.6151
R2235 B.n836 B.n835 10.6151
R2236 B.n836 B.n604 10.6151
R2237 B.n842 B.n604 10.6151
R2238 B.n843 B.n842 10.6151
R2239 B.n844 B.n843 10.6151
R2240 B.n844 B.n602 10.6151
R2241 B.n850 B.n602 10.6151
R2242 B.n851 B.n850 10.6151
R2243 B.n852 B.n851 10.6151
R2244 B.n852 B.n600 10.6151
R2245 B.n858 B.n600 10.6151
R2246 B.n859 B.n858 10.6151
R2247 B.n860 B.n859 10.6151
R2248 B.n860 B.n598 10.6151
R2249 B.n866 B.n598 10.6151
R2250 B.n867 B.n866 10.6151
R2251 B.n868 B.n867 10.6151
R2252 B.n868 B.n596 10.6151
R2253 B.n874 B.n596 10.6151
R2254 B.n875 B.n874 10.6151
R2255 B.n876 B.n875 10.6151
R2256 B.n876 B.n594 10.6151
R2257 B.n882 B.n594 10.6151
R2258 B.n883 B.n882 10.6151
R2259 B.n884 B.n883 10.6151
R2260 B.n884 B.n592 10.6151
R2261 B.n592 B.n591 10.6151
R2262 B.n891 B.n591 10.6151
R2263 B.n892 B.n891 10.6151
R2264 B.n893 B.n583 10.6151
R2265 B.n903 B.n583 10.6151
R2266 B.n904 B.n903 10.6151
R2267 B.n905 B.n904 10.6151
R2268 B.n905 B.n575 10.6151
R2269 B.n915 B.n575 10.6151
R2270 B.n916 B.n915 10.6151
R2271 B.n917 B.n916 10.6151
R2272 B.n917 B.n567 10.6151
R2273 B.n927 B.n567 10.6151
R2274 B.n928 B.n927 10.6151
R2275 B.n929 B.n928 10.6151
R2276 B.n929 B.n559 10.6151
R2277 B.n939 B.n559 10.6151
R2278 B.n940 B.n939 10.6151
R2279 B.n941 B.n940 10.6151
R2280 B.n941 B.n551 10.6151
R2281 B.n951 B.n551 10.6151
R2282 B.n952 B.n951 10.6151
R2283 B.n953 B.n952 10.6151
R2284 B.n953 B.n542 10.6151
R2285 B.n963 B.n542 10.6151
R2286 B.n964 B.n963 10.6151
R2287 B.n965 B.n964 10.6151
R2288 B.n965 B.n535 10.6151
R2289 B.n975 B.n535 10.6151
R2290 B.n976 B.n975 10.6151
R2291 B.n977 B.n976 10.6151
R2292 B.n977 B.n527 10.6151
R2293 B.n987 B.n527 10.6151
R2294 B.n988 B.n987 10.6151
R2295 B.n989 B.n988 10.6151
R2296 B.n989 B.n519 10.6151
R2297 B.n999 B.n519 10.6151
R2298 B.n1000 B.n999 10.6151
R2299 B.n1001 B.n1000 10.6151
R2300 B.n1001 B.n511 10.6151
R2301 B.n1011 B.n511 10.6151
R2302 B.n1012 B.n1011 10.6151
R2303 B.n1013 B.n1012 10.6151
R2304 B.n1013 B.n503 10.6151
R2305 B.n1023 B.n503 10.6151
R2306 B.n1024 B.n1023 10.6151
R2307 B.n1025 B.n1024 10.6151
R2308 B.n1025 B.n495 10.6151
R2309 B.n1035 B.n495 10.6151
R2310 B.n1036 B.n1035 10.6151
R2311 B.n1037 B.n1036 10.6151
R2312 B.n1037 B.n487 10.6151
R2313 B.n1047 B.n487 10.6151
R2314 B.n1048 B.n1047 10.6151
R2315 B.n1049 B.n1048 10.6151
R2316 B.n1049 B.n479 10.6151
R2317 B.n1059 B.n479 10.6151
R2318 B.n1060 B.n1059 10.6151
R2319 B.n1061 B.n1060 10.6151
R2320 B.n1061 B.n472 10.6151
R2321 B.n1072 B.n472 10.6151
R2322 B.n1073 B.n1072 10.6151
R2323 B.n1074 B.n1073 10.6151
R2324 B.n1074 B.n464 10.6151
R2325 B.n1084 B.n464 10.6151
R2326 B.n1085 B.n1084 10.6151
R2327 B.n1086 B.n1085 10.6151
R2328 B.n1086 B.n456 10.6151
R2329 B.n1096 B.n456 10.6151
R2330 B.n1097 B.n1096 10.6151
R2331 B.n1098 B.n1097 10.6151
R2332 B.n1098 B.n449 10.6151
R2333 B.n1109 B.n449 10.6151
R2334 B.n1110 B.n1109 10.6151
R2335 B.n1112 B.n1110 10.6151
R2336 B.n1112 B.n1111 10.6151
R2337 B.n1111 B.n441 10.6151
R2338 B.n1123 B.n441 10.6151
R2339 B.n1124 B.n1123 10.6151
R2340 B.n1125 B.n1124 10.6151
R2341 B.n1126 B.n1125 10.6151
R2342 B.n1127 B.n1126 10.6151
R2343 B.n1130 B.n1127 10.6151
R2344 B.n1131 B.n1130 10.6151
R2345 B.n1132 B.n1131 10.6151
R2346 B.n1133 B.n1132 10.6151
R2347 B.n1135 B.n1133 10.6151
R2348 B.n1136 B.n1135 10.6151
R2349 B.n1137 B.n1136 10.6151
R2350 B.n1138 B.n1137 10.6151
R2351 B.n1140 B.n1138 10.6151
R2352 B.n1141 B.n1140 10.6151
R2353 B.n1142 B.n1141 10.6151
R2354 B.n1143 B.n1142 10.6151
R2355 B.n1145 B.n1143 10.6151
R2356 B.n1146 B.n1145 10.6151
R2357 B.n1147 B.n1146 10.6151
R2358 B.n1148 B.n1147 10.6151
R2359 B.n1150 B.n1148 10.6151
R2360 B.n1151 B.n1150 10.6151
R2361 B.n1152 B.n1151 10.6151
R2362 B.n1153 B.n1152 10.6151
R2363 B.n1155 B.n1153 10.6151
R2364 B.n1156 B.n1155 10.6151
R2365 B.n1157 B.n1156 10.6151
R2366 B.n1158 B.n1157 10.6151
R2367 B.n1160 B.n1158 10.6151
R2368 B.n1161 B.n1160 10.6151
R2369 B.n1162 B.n1161 10.6151
R2370 B.n1163 B.n1162 10.6151
R2371 B.n1165 B.n1163 10.6151
R2372 B.n1166 B.n1165 10.6151
R2373 B.n1167 B.n1166 10.6151
R2374 B.n1168 B.n1167 10.6151
R2375 B.n1170 B.n1168 10.6151
R2376 B.n1171 B.n1170 10.6151
R2377 B.n1172 B.n1171 10.6151
R2378 B.n1173 B.n1172 10.6151
R2379 B.n1175 B.n1173 10.6151
R2380 B.n1176 B.n1175 10.6151
R2381 B.n1177 B.n1176 10.6151
R2382 B.n1178 B.n1177 10.6151
R2383 B.n1180 B.n1178 10.6151
R2384 B.n1181 B.n1180 10.6151
R2385 B.n1182 B.n1181 10.6151
R2386 B.n1183 B.n1182 10.6151
R2387 B.n1185 B.n1183 10.6151
R2388 B.n1186 B.n1185 10.6151
R2389 B.n1187 B.n1186 10.6151
R2390 B.n1188 B.n1187 10.6151
R2391 B.n1190 B.n1188 10.6151
R2392 B.n1191 B.n1190 10.6151
R2393 B.n1192 B.n1191 10.6151
R2394 B.n1193 B.n1192 10.6151
R2395 B.n1195 B.n1193 10.6151
R2396 B.n1196 B.n1195 10.6151
R2397 B.n1197 B.n1196 10.6151
R2398 B.n1198 B.n1197 10.6151
R2399 B.n1200 B.n1198 10.6151
R2400 B.n1201 B.n1200 10.6151
R2401 B.n1202 B.n1201 10.6151
R2402 B.n1203 B.n1202 10.6151
R2403 B.n1205 B.n1203 10.6151
R2404 B.n1206 B.n1205 10.6151
R2405 B.n1207 B.n1206 10.6151
R2406 B.n1208 B.n1207 10.6151
R2407 B.n1210 B.n1208 10.6151
R2408 B.n1211 B.n1210 10.6151
R2409 B.n1212 B.n1211 10.6151
R2410 B.n1213 B.n1212 10.6151
R2411 B.n1215 B.n1213 10.6151
R2412 B.n1216 B.n1215 10.6151
R2413 B.n1217 B.n1216 10.6151
R2414 B.n1218 B.n1217 10.6151
R2415 B.n1220 B.n1218 10.6151
R2416 B.n1221 B.n1220 10.6151
R2417 B.n1374 B.n1 10.6151
R2418 B.n1374 B.n1373 10.6151
R2419 B.n1373 B.n1372 10.6151
R2420 B.n1372 B.n10 10.6151
R2421 B.n1366 B.n10 10.6151
R2422 B.n1366 B.n1365 10.6151
R2423 B.n1365 B.n1364 10.6151
R2424 B.n1364 B.n17 10.6151
R2425 B.n1358 B.n17 10.6151
R2426 B.n1358 B.n1357 10.6151
R2427 B.n1357 B.n1356 10.6151
R2428 B.n1356 B.n25 10.6151
R2429 B.n1350 B.n25 10.6151
R2430 B.n1350 B.n1349 10.6151
R2431 B.n1349 B.n1348 10.6151
R2432 B.n1348 B.n32 10.6151
R2433 B.n1342 B.n32 10.6151
R2434 B.n1342 B.n1341 10.6151
R2435 B.n1341 B.n1340 10.6151
R2436 B.n1340 B.n38 10.6151
R2437 B.n1334 B.n38 10.6151
R2438 B.n1334 B.n1333 10.6151
R2439 B.n1333 B.n1332 10.6151
R2440 B.n1332 B.n46 10.6151
R2441 B.n1326 B.n46 10.6151
R2442 B.n1326 B.n1325 10.6151
R2443 B.n1325 B.n1324 10.6151
R2444 B.n1324 B.n53 10.6151
R2445 B.n1318 B.n53 10.6151
R2446 B.n1318 B.n1317 10.6151
R2447 B.n1317 B.n1316 10.6151
R2448 B.n1316 B.n60 10.6151
R2449 B.n1310 B.n60 10.6151
R2450 B.n1310 B.n1309 10.6151
R2451 B.n1309 B.n1308 10.6151
R2452 B.n1308 B.n67 10.6151
R2453 B.n1302 B.n67 10.6151
R2454 B.n1302 B.n1301 10.6151
R2455 B.n1301 B.n1300 10.6151
R2456 B.n1300 B.n74 10.6151
R2457 B.n1294 B.n74 10.6151
R2458 B.n1294 B.n1293 10.6151
R2459 B.n1293 B.n1292 10.6151
R2460 B.n1292 B.n81 10.6151
R2461 B.n1286 B.n81 10.6151
R2462 B.n1286 B.n1285 10.6151
R2463 B.n1285 B.n1284 10.6151
R2464 B.n1284 B.n88 10.6151
R2465 B.n1278 B.n88 10.6151
R2466 B.n1278 B.n1277 10.6151
R2467 B.n1277 B.n1276 10.6151
R2468 B.n1276 B.n95 10.6151
R2469 B.n1270 B.n95 10.6151
R2470 B.n1270 B.n1269 10.6151
R2471 B.n1269 B.n1268 10.6151
R2472 B.n1268 B.n102 10.6151
R2473 B.n1262 B.n102 10.6151
R2474 B.n1262 B.n1261 10.6151
R2475 B.n1261 B.n1260 10.6151
R2476 B.n1260 B.n109 10.6151
R2477 B.n1254 B.n109 10.6151
R2478 B.n1254 B.n1253 10.6151
R2479 B.n1253 B.n1252 10.6151
R2480 B.n1252 B.n116 10.6151
R2481 B.n1246 B.n116 10.6151
R2482 B.n1246 B.n1245 10.6151
R2483 B.n1245 B.n1244 10.6151
R2484 B.n1244 B.n123 10.6151
R2485 B.n1238 B.n123 10.6151
R2486 B.n1238 B.n1237 10.6151
R2487 B.n1237 B.n1236 10.6151
R2488 B.n1236 B.n130 10.6151
R2489 B.n1230 B.n130 10.6151
R2490 B.n1230 B.n1229 10.6151
R2491 B.n1229 B.n1228 10.6151
R2492 B.n204 B.n137 10.6151
R2493 B.n207 B.n204 10.6151
R2494 B.n208 B.n207 10.6151
R2495 B.n211 B.n208 10.6151
R2496 B.n212 B.n211 10.6151
R2497 B.n215 B.n212 10.6151
R2498 B.n216 B.n215 10.6151
R2499 B.n219 B.n216 10.6151
R2500 B.n220 B.n219 10.6151
R2501 B.n223 B.n220 10.6151
R2502 B.n224 B.n223 10.6151
R2503 B.n227 B.n224 10.6151
R2504 B.n228 B.n227 10.6151
R2505 B.n231 B.n228 10.6151
R2506 B.n232 B.n231 10.6151
R2507 B.n235 B.n232 10.6151
R2508 B.n236 B.n235 10.6151
R2509 B.n239 B.n236 10.6151
R2510 B.n240 B.n239 10.6151
R2511 B.n243 B.n240 10.6151
R2512 B.n244 B.n243 10.6151
R2513 B.n247 B.n244 10.6151
R2514 B.n248 B.n247 10.6151
R2515 B.n251 B.n248 10.6151
R2516 B.n252 B.n251 10.6151
R2517 B.n255 B.n252 10.6151
R2518 B.n256 B.n255 10.6151
R2519 B.n259 B.n256 10.6151
R2520 B.n260 B.n259 10.6151
R2521 B.n263 B.n260 10.6151
R2522 B.n264 B.n263 10.6151
R2523 B.n267 B.n264 10.6151
R2524 B.n268 B.n267 10.6151
R2525 B.n271 B.n268 10.6151
R2526 B.n272 B.n271 10.6151
R2527 B.n275 B.n272 10.6151
R2528 B.n276 B.n275 10.6151
R2529 B.n279 B.n276 10.6151
R2530 B.n280 B.n279 10.6151
R2531 B.n283 B.n280 10.6151
R2532 B.n284 B.n283 10.6151
R2533 B.n287 B.n284 10.6151
R2534 B.n288 B.n287 10.6151
R2535 B.n291 B.n288 10.6151
R2536 B.n292 B.n291 10.6151
R2537 B.n295 B.n292 10.6151
R2538 B.n296 B.n295 10.6151
R2539 B.n299 B.n296 10.6151
R2540 B.n300 B.n299 10.6151
R2541 B.n303 B.n300 10.6151
R2542 B.n304 B.n303 10.6151
R2543 B.n307 B.n304 10.6151
R2544 B.n308 B.n307 10.6151
R2545 B.n311 B.n308 10.6151
R2546 B.n316 B.n313 10.6151
R2547 B.n317 B.n316 10.6151
R2548 B.n320 B.n317 10.6151
R2549 B.n321 B.n320 10.6151
R2550 B.n324 B.n321 10.6151
R2551 B.n325 B.n324 10.6151
R2552 B.n328 B.n325 10.6151
R2553 B.n329 B.n328 10.6151
R2554 B.n332 B.n329 10.6151
R2555 B.n337 B.n334 10.6151
R2556 B.n338 B.n337 10.6151
R2557 B.n341 B.n338 10.6151
R2558 B.n342 B.n341 10.6151
R2559 B.n345 B.n342 10.6151
R2560 B.n346 B.n345 10.6151
R2561 B.n349 B.n346 10.6151
R2562 B.n350 B.n349 10.6151
R2563 B.n353 B.n350 10.6151
R2564 B.n354 B.n353 10.6151
R2565 B.n357 B.n354 10.6151
R2566 B.n358 B.n357 10.6151
R2567 B.n361 B.n358 10.6151
R2568 B.n362 B.n361 10.6151
R2569 B.n365 B.n362 10.6151
R2570 B.n366 B.n365 10.6151
R2571 B.n369 B.n366 10.6151
R2572 B.n370 B.n369 10.6151
R2573 B.n373 B.n370 10.6151
R2574 B.n374 B.n373 10.6151
R2575 B.n377 B.n374 10.6151
R2576 B.n378 B.n377 10.6151
R2577 B.n381 B.n378 10.6151
R2578 B.n382 B.n381 10.6151
R2579 B.n385 B.n382 10.6151
R2580 B.n386 B.n385 10.6151
R2581 B.n389 B.n386 10.6151
R2582 B.n390 B.n389 10.6151
R2583 B.n393 B.n390 10.6151
R2584 B.n394 B.n393 10.6151
R2585 B.n397 B.n394 10.6151
R2586 B.n398 B.n397 10.6151
R2587 B.n401 B.n398 10.6151
R2588 B.n402 B.n401 10.6151
R2589 B.n405 B.n402 10.6151
R2590 B.n406 B.n405 10.6151
R2591 B.n409 B.n406 10.6151
R2592 B.n410 B.n409 10.6151
R2593 B.n413 B.n410 10.6151
R2594 B.n414 B.n413 10.6151
R2595 B.n417 B.n414 10.6151
R2596 B.n418 B.n417 10.6151
R2597 B.n421 B.n418 10.6151
R2598 B.n422 B.n421 10.6151
R2599 B.n425 B.n422 10.6151
R2600 B.n426 B.n425 10.6151
R2601 B.n429 B.n426 10.6151
R2602 B.n430 B.n429 10.6151
R2603 B.n433 B.n430 10.6151
R2604 B.n434 B.n433 10.6151
R2605 B.n437 B.n434 10.6151
R2606 B.n439 B.n437 10.6151
R2607 B.n440 B.n439 10.6151
R2608 B.n1222 B.n440 10.6151
R2609 B.n763 B.n762 9.36635
R2610 B.n786 B.n620 9.36635
R2611 B.n312 B.n311 9.36635
R2612 B.n334 B.n333 9.36635
R2613 B.n1382 B.n0 8.11757
R2614 B.n1382 B.n1 8.11757
R2615 B.n1070 B.t9 7.54336
R2616 B.n1344 B.t3 7.54336
R2617 B.n1100 B.t1 6.53764
R2618 B.n19 B.t6 6.53764
R2619 B.t15 B.n569 2.51479
R2620 B.t11 B.n121 2.51479
R2621 B.t2 B.n517 1.50907
R2622 B.n1297 B.t8 1.50907
R2623 B.n764 B.n763 1.24928
R2624 B.n621 B.n620 1.24928
R2625 B.n313 B.n312 1.24928
R2626 B.n333 B.n332 1.24928
R2627 VN.n100 VN.n99 161.3
R2628 VN.n98 VN.n52 161.3
R2629 VN.n97 VN.n96 161.3
R2630 VN.n95 VN.n53 161.3
R2631 VN.n94 VN.n93 161.3
R2632 VN.n92 VN.n54 161.3
R2633 VN.n91 VN.n90 161.3
R2634 VN.n89 VN.n55 161.3
R2635 VN.n88 VN.n87 161.3
R2636 VN.n86 VN.n56 161.3
R2637 VN.n85 VN.n84 161.3
R2638 VN.n83 VN.n58 161.3
R2639 VN.n82 VN.n81 161.3
R2640 VN.n80 VN.n59 161.3
R2641 VN.n79 VN.n78 161.3
R2642 VN.n77 VN.n60 161.3
R2643 VN.n76 VN.n75 161.3
R2644 VN.n74 VN.n61 161.3
R2645 VN.n73 VN.n72 161.3
R2646 VN.n71 VN.n62 161.3
R2647 VN.n70 VN.n69 161.3
R2648 VN.n68 VN.n63 161.3
R2649 VN.n67 VN.n66 161.3
R2650 VN.n49 VN.n48 161.3
R2651 VN.n47 VN.n1 161.3
R2652 VN.n46 VN.n45 161.3
R2653 VN.n44 VN.n2 161.3
R2654 VN.n43 VN.n42 161.3
R2655 VN.n41 VN.n3 161.3
R2656 VN.n40 VN.n39 161.3
R2657 VN.n38 VN.n4 161.3
R2658 VN.n37 VN.n36 161.3
R2659 VN.n34 VN.n5 161.3
R2660 VN.n33 VN.n32 161.3
R2661 VN.n31 VN.n6 161.3
R2662 VN.n30 VN.n29 161.3
R2663 VN.n28 VN.n7 161.3
R2664 VN.n27 VN.n26 161.3
R2665 VN.n25 VN.n8 161.3
R2666 VN.n24 VN.n23 161.3
R2667 VN.n22 VN.n9 161.3
R2668 VN.n21 VN.n20 161.3
R2669 VN.n19 VN.n10 161.3
R2670 VN.n18 VN.n17 161.3
R2671 VN.n16 VN.n11 161.3
R2672 VN.n15 VN.n14 161.3
R2673 VN.n13 VN.t7 146.381
R2674 VN.n65 VN.t5 146.381
R2675 VN.n8 VN.t8 112.694
R2676 VN.n12 VN.t9 112.694
R2677 VN.n35 VN.t4 112.694
R2678 VN.n0 VN.t2 112.694
R2679 VN.n60 VN.t1 112.694
R2680 VN.n64 VN.t0 112.694
R2681 VN.n57 VN.t3 112.694
R2682 VN.n51 VN.t6 112.694
R2683 VN.n50 VN.n0 77.2324
R2684 VN.n101 VN.n51 77.2324
R2685 VN VN.n101 62.0737
R2686 VN.n42 VN.n2 56.4773
R2687 VN.n93 VN.n53 56.4773
R2688 VN.n13 VN.n12 55.9618
R2689 VN.n65 VN.n64 55.9618
R2690 VN.n21 VN.n10 46.253
R2691 VN.n29 VN.n6 46.253
R2692 VN.n73 VN.n62 46.253
R2693 VN.n81 VN.n58 46.253
R2694 VN.n17 VN.n10 34.5682
R2695 VN.n33 VN.n6 34.5682
R2696 VN.n69 VN.n62 34.5682
R2697 VN.n85 VN.n58 34.5682
R2698 VN.n16 VN.n15 24.3439
R2699 VN.n17 VN.n16 24.3439
R2700 VN.n22 VN.n21 24.3439
R2701 VN.n23 VN.n22 24.3439
R2702 VN.n23 VN.n8 24.3439
R2703 VN.n27 VN.n8 24.3439
R2704 VN.n28 VN.n27 24.3439
R2705 VN.n29 VN.n28 24.3439
R2706 VN.n34 VN.n33 24.3439
R2707 VN.n36 VN.n34 24.3439
R2708 VN.n40 VN.n4 24.3439
R2709 VN.n41 VN.n40 24.3439
R2710 VN.n42 VN.n41 24.3439
R2711 VN.n46 VN.n2 24.3439
R2712 VN.n47 VN.n46 24.3439
R2713 VN.n48 VN.n47 24.3439
R2714 VN.n69 VN.n68 24.3439
R2715 VN.n68 VN.n67 24.3439
R2716 VN.n81 VN.n80 24.3439
R2717 VN.n80 VN.n79 24.3439
R2718 VN.n79 VN.n60 24.3439
R2719 VN.n75 VN.n60 24.3439
R2720 VN.n75 VN.n74 24.3439
R2721 VN.n74 VN.n73 24.3439
R2722 VN.n93 VN.n92 24.3439
R2723 VN.n92 VN.n91 24.3439
R2724 VN.n91 VN.n55 24.3439
R2725 VN.n87 VN.n86 24.3439
R2726 VN.n86 VN.n85 24.3439
R2727 VN.n99 VN.n98 24.3439
R2728 VN.n98 VN.n97 24.3439
R2729 VN.n97 VN.n53 24.3439
R2730 VN.n15 VN.n12 18.5015
R2731 VN.n36 VN.n35 18.5015
R2732 VN.n67 VN.n64 18.5015
R2733 VN.n87 VN.n57 18.5015
R2734 VN.n48 VN.n0 12.6591
R2735 VN.n99 VN.n51 12.6591
R2736 VN.n35 VN.n4 5.84292
R2737 VN.n57 VN.n55 5.84292
R2738 VN.n14 VN.n13 3.08092
R2739 VN.n66 VN.n65 3.08092
R2740 VN.n101 VN.n100 0.355081
R2741 VN.n50 VN.n49 0.355081
R2742 VN VN.n50 0.26685
R2743 VN.n100 VN.n52 0.189894
R2744 VN.n96 VN.n52 0.189894
R2745 VN.n96 VN.n95 0.189894
R2746 VN.n95 VN.n94 0.189894
R2747 VN.n94 VN.n54 0.189894
R2748 VN.n90 VN.n54 0.189894
R2749 VN.n90 VN.n89 0.189894
R2750 VN.n89 VN.n88 0.189894
R2751 VN.n88 VN.n56 0.189894
R2752 VN.n84 VN.n56 0.189894
R2753 VN.n84 VN.n83 0.189894
R2754 VN.n83 VN.n82 0.189894
R2755 VN.n82 VN.n59 0.189894
R2756 VN.n78 VN.n59 0.189894
R2757 VN.n78 VN.n77 0.189894
R2758 VN.n77 VN.n76 0.189894
R2759 VN.n76 VN.n61 0.189894
R2760 VN.n72 VN.n61 0.189894
R2761 VN.n72 VN.n71 0.189894
R2762 VN.n71 VN.n70 0.189894
R2763 VN.n70 VN.n63 0.189894
R2764 VN.n66 VN.n63 0.189894
R2765 VN.n14 VN.n11 0.189894
R2766 VN.n18 VN.n11 0.189894
R2767 VN.n19 VN.n18 0.189894
R2768 VN.n20 VN.n19 0.189894
R2769 VN.n20 VN.n9 0.189894
R2770 VN.n24 VN.n9 0.189894
R2771 VN.n25 VN.n24 0.189894
R2772 VN.n26 VN.n25 0.189894
R2773 VN.n26 VN.n7 0.189894
R2774 VN.n30 VN.n7 0.189894
R2775 VN.n31 VN.n30 0.189894
R2776 VN.n32 VN.n31 0.189894
R2777 VN.n32 VN.n5 0.189894
R2778 VN.n37 VN.n5 0.189894
R2779 VN.n38 VN.n37 0.189894
R2780 VN.n39 VN.n38 0.189894
R2781 VN.n39 VN.n3 0.189894
R2782 VN.n43 VN.n3 0.189894
R2783 VN.n44 VN.n43 0.189894
R2784 VN.n45 VN.n44 0.189894
R2785 VN.n45 VN.n1 0.189894
R2786 VN.n49 VN.n1 0.189894
R2787 VDD2.n1 VDD2.t2 68.39
R2788 VDD2.n3 VDD2.n2 66.3057
R2789 VDD2 VDD2.n7 66.3029
R2790 VDD2.n4 VDD2.t3 65.0454
R2791 VDD2.n6 VDD2.n5 63.8527
R2792 VDD2.n1 VDD2.n0 63.8524
R2793 VDD2.n4 VDD2.n3 53.9136
R2794 VDD2.n6 VDD2.n4 3.34533
R2795 VDD2.n7 VDD2.t9 1.19327
R2796 VDD2.n7 VDD2.t4 1.19327
R2797 VDD2.n5 VDD2.t6 1.19327
R2798 VDD2.n5 VDD2.t8 1.19327
R2799 VDD2.n2 VDD2.t5 1.19327
R2800 VDD2.n2 VDD2.t7 1.19327
R2801 VDD2.n0 VDD2.t0 1.19327
R2802 VDD2.n0 VDD2.t1 1.19327
R2803 VDD2 VDD2.n6 0.894897
R2804 VDD2.n3 VDD2.n1 0.781361
C0 VP VDD2 0.704728f
C1 VTAIL VDD1 12.669701f
C2 VTAIL VDD2 12.727f
C3 VN VDD1 0.15518f
C4 VN VDD2 15.370099f
C5 VDD1 VDD2 2.79353f
C6 VP VTAIL 16.216f
C7 VP VN 10.657901f
C8 VN VTAIL 16.2017f
C9 VP VDD1 15.9151f
C10 VDD2 B 9.102519f
C11 VDD1 B 9.094422f
C12 VTAIL B 10.792514f
C13 VN B 23.03454f
C14 VP B 21.574484f
C15 VDD2.t2 B 3.67103f
C16 VDD2.t0 B 0.313746f
C17 VDD2.t1 B 0.313746f
C18 VDD2.n0 B 2.85198f
C19 VDD2.n1 B 1.01114f
C20 VDD2.t5 B 0.313746f
C21 VDD2.t7 B 0.313746f
C22 VDD2.n2 B 2.87606f
C23 VDD2.n3 B 3.52694f
C24 VDD2.t3 B 3.64541f
C25 VDD2.n4 B 3.67431f
C26 VDD2.t6 B 0.313746f
C27 VDD2.t8 B 0.313746f
C28 VDD2.n5 B 2.85198f
C29 VDD2.n6 B 0.52093f
C30 VDD2.t9 B 0.313746f
C31 VDD2.t4 B 0.313746f
C32 VDD2.n7 B 2.87601f
C33 VN.t2 B 2.70996f
C34 VN.n0 B 1.00606f
C35 VN.n1 B 0.016745f
C36 VN.n2 B 0.021262f
C37 VN.n3 B 0.016745f
C38 VN.n4 B 0.019596f
C39 VN.n5 B 0.016745f
C40 VN.n6 B 0.014347f
C41 VN.n7 B 0.016745f
C42 VN.t8 B 2.70996f
C43 VN.n8 B 0.953195f
C44 VN.n9 B 0.016745f
C45 VN.n10 B 0.014347f
C46 VN.n11 B 0.016745f
C47 VN.t9 B 2.70996f
C48 VN.n12 B 1.00012f
C49 VN.t7 B 2.95528f
C50 VN.n13 B 0.950672f
C51 VN.n14 B 0.20714f
C52 VN.n15 B 0.027649f
C53 VN.n16 B 0.031366f
C54 VN.n17 B 0.034022f
C55 VN.n18 B 0.016745f
C56 VN.n19 B 0.016745f
C57 VN.n20 B 0.016745f
C58 VN.n21 B 0.032099f
C59 VN.n22 B 0.031366f
C60 VN.n23 B 0.031366f
C61 VN.n24 B 0.016745f
C62 VN.n25 B 0.016745f
C63 VN.n26 B 0.016745f
C64 VN.n27 B 0.031366f
C65 VN.n28 B 0.031366f
C66 VN.n29 B 0.032099f
C67 VN.n30 B 0.016745f
C68 VN.n31 B 0.016745f
C69 VN.n32 B 0.016745f
C70 VN.n33 B 0.034022f
C71 VN.n34 B 0.031366f
C72 VN.t4 B 2.70996f
C73 VN.n35 B 0.937316f
C74 VN.n36 B 0.027649f
C75 VN.n37 B 0.016745f
C76 VN.n38 B 0.016745f
C77 VN.n39 B 0.016745f
C78 VN.n40 B 0.031366f
C79 VN.n41 B 0.031366f
C80 VN.n42 B 0.027841f
C81 VN.n43 B 0.016745f
C82 VN.n44 B 0.016745f
C83 VN.n45 B 0.016745f
C84 VN.n46 B 0.031366f
C85 VN.n47 B 0.031366f
C86 VN.n48 B 0.023932f
C87 VN.n49 B 0.027031f
C88 VN.n50 B 0.04367f
C89 VN.t6 B 2.70996f
C90 VN.n51 B 1.00606f
C91 VN.n52 B 0.016745f
C92 VN.n53 B 0.021262f
C93 VN.n54 B 0.016745f
C94 VN.n55 B 0.019596f
C95 VN.n56 B 0.016745f
C96 VN.t3 B 2.70996f
C97 VN.n57 B 0.937316f
C98 VN.n58 B 0.014347f
C99 VN.n59 B 0.016745f
C100 VN.t1 B 2.70996f
C101 VN.n60 B 0.953195f
C102 VN.n61 B 0.016745f
C103 VN.n62 B 0.014347f
C104 VN.n63 B 0.016745f
C105 VN.t0 B 2.70996f
C106 VN.n64 B 1.00012f
C107 VN.t5 B 2.95528f
C108 VN.n65 B 0.950672f
C109 VN.n66 B 0.20714f
C110 VN.n67 B 0.027649f
C111 VN.n68 B 0.031366f
C112 VN.n69 B 0.034022f
C113 VN.n70 B 0.016745f
C114 VN.n71 B 0.016745f
C115 VN.n72 B 0.016745f
C116 VN.n73 B 0.032099f
C117 VN.n74 B 0.031366f
C118 VN.n75 B 0.031366f
C119 VN.n76 B 0.016745f
C120 VN.n77 B 0.016745f
C121 VN.n78 B 0.016745f
C122 VN.n79 B 0.031366f
C123 VN.n80 B 0.031366f
C124 VN.n81 B 0.032099f
C125 VN.n82 B 0.016745f
C126 VN.n83 B 0.016745f
C127 VN.n84 B 0.016745f
C128 VN.n85 B 0.034022f
C129 VN.n86 B 0.031366f
C130 VN.n87 B 0.027649f
C131 VN.n88 B 0.016745f
C132 VN.n89 B 0.016745f
C133 VN.n90 B 0.016745f
C134 VN.n91 B 0.031366f
C135 VN.n92 B 0.031366f
C136 VN.n93 B 0.027841f
C137 VN.n94 B 0.016745f
C138 VN.n95 B 0.016745f
C139 VN.n96 B 0.016745f
C140 VN.n97 B 0.031366f
C141 VN.n98 B 0.031366f
C142 VN.n99 B 0.023932f
C143 VN.n100 B 0.027031f
C144 VN.n101 B 1.28896f
C145 VDD1.t8 B 3.7198f
C146 VDD1.t5 B 0.317914f
C147 VDD1.t3 B 0.317914f
C148 VDD1.n0 B 2.88987f
C149 VDD1.n1 B 1.03272f
C150 VDD1.t1 B 3.7198f
C151 VDD1.t2 B 0.317914f
C152 VDD1.t0 B 0.317914f
C153 VDD1.n2 B 2.88986f
C154 VDD1.n3 B 1.02458f
C155 VDD1.t6 B 0.317914f
C156 VDD1.t7 B 0.317914f
C157 VDD1.n4 B 2.91427f
C158 VDD1.n5 B 3.72349f
C159 VDD1.t4 B 0.317914f
C160 VDD1.t9 B 0.317914f
C161 VDD1.n6 B 2.88986f
C162 VDD1.n7 B 3.79124f
C163 VTAIL.t6 B 0.320118f
C164 VTAIL.t3 B 0.320118f
C165 VTAIL.n0 B 2.84148f
C166 VTAIL.n1 B 0.60371f
C167 VTAIL.t12 B 3.63081f
C168 VTAIL.n2 B 0.748599f
C169 VTAIL.t16 B 0.320118f
C170 VTAIL.t15 B 0.320118f
C171 VTAIL.n3 B 2.84148f
C172 VTAIL.n4 B 0.759451f
C173 VTAIL.t18 B 0.320118f
C174 VTAIL.t9 B 0.320118f
C175 VTAIL.n5 B 2.84148f
C176 VTAIL.n6 B 2.47922f
C177 VTAIL.t0 B 0.320118f
C178 VTAIL.t2 B 0.320118f
C179 VTAIL.n7 B 2.84148f
C180 VTAIL.n8 B 2.47922f
C181 VTAIL.t4 B 0.320118f
C182 VTAIL.t19 B 0.320118f
C183 VTAIL.n9 B 2.84148f
C184 VTAIL.n10 B 0.759448f
C185 VTAIL.t1 B 3.63082f
C186 VTAIL.n11 B 0.748595f
C187 VTAIL.t11 B 0.320118f
C188 VTAIL.t13 B 0.320118f
C189 VTAIL.n12 B 2.84148f
C190 VTAIL.n13 B 0.664885f
C191 VTAIL.t17 B 0.320118f
C192 VTAIL.t10 B 0.320118f
C193 VTAIL.n14 B 2.84148f
C194 VTAIL.n15 B 0.759448f
C195 VTAIL.t14 B 3.63081f
C196 VTAIL.n16 B 2.29992f
C197 VTAIL.t7 B 3.63081f
C198 VTAIL.n17 B 2.29992f
C199 VTAIL.t5 B 0.320118f
C200 VTAIL.t8 B 0.320118f
C201 VTAIL.n18 B 2.84148f
C202 VTAIL.n19 B 0.557615f
C203 VP.t2 B 2.74352f
C204 VP.n0 B 1.01851f
C205 VP.n1 B 0.016953f
C206 VP.n2 B 0.021525f
C207 VP.n3 B 0.016953f
C208 VP.n4 B 0.019839f
C209 VP.n5 B 0.016953f
C210 VP.n6 B 0.014525f
C211 VP.n7 B 0.016953f
C212 VP.t9 B 2.74352f
C213 VP.n8 B 0.964999f
C214 VP.n9 B 0.016953f
C215 VP.n10 B 0.014525f
C216 VP.n11 B 0.016953f
C217 VP.t7 B 2.74352f
C218 VP.n12 B 0.948923f
C219 VP.n13 B 0.016953f
C220 VP.n14 B 0.028186f
C221 VP.n15 B 0.016953f
C222 VP.n16 B 0.024229f
C223 VP.t0 B 2.74352f
C224 VP.n17 B 1.01851f
C225 VP.n18 B 0.016953f
C226 VP.n19 B 0.021525f
C227 VP.n20 B 0.016953f
C228 VP.n21 B 0.019839f
C229 VP.n22 B 0.016953f
C230 VP.n23 B 0.014525f
C231 VP.n24 B 0.016953f
C232 VP.t6 B 2.74352f
C233 VP.n25 B 0.964999f
C234 VP.n26 B 0.016953f
C235 VP.n27 B 0.014525f
C236 VP.n28 B 0.016953f
C237 VP.t4 B 2.74352f
C238 VP.n29 B 1.0125f
C239 VP.t1 B 2.99188f
C240 VP.n30 B 0.962445f
C241 VP.n31 B 0.209705f
C242 VP.n32 B 0.027991f
C243 VP.n33 B 0.031754f
C244 VP.n34 B 0.034444f
C245 VP.n35 B 0.016953f
C246 VP.n36 B 0.016953f
C247 VP.n37 B 0.016953f
C248 VP.n38 B 0.032497f
C249 VP.n39 B 0.031754f
C250 VP.n40 B 0.031754f
C251 VP.n41 B 0.016953f
C252 VP.n42 B 0.016953f
C253 VP.n43 B 0.016953f
C254 VP.n44 B 0.031754f
C255 VP.n45 B 0.031754f
C256 VP.n46 B 0.032497f
C257 VP.n47 B 0.016953f
C258 VP.n48 B 0.016953f
C259 VP.n49 B 0.016953f
C260 VP.n50 B 0.034444f
C261 VP.n51 B 0.031754f
C262 VP.t5 B 2.74352f
C263 VP.n52 B 0.948923f
C264 VP.n53 B 0.027991f
C265 VP.n54 B 0.016953f
C266 VP.n55 B 0.016953f
C267 VP.n56 B 0.016953f
C268 VP.n57 B 0.031754f
C269 VP.n58 B 0.031754f
C270 VP.n59 B 0.028186f
C271 VP.n60 B 0.016953f
C272 VP.n61 B 0.016953f
C273 VP.n62 B 0.016953f
C274 VP.n63 B 0.031754f
C275 VP.n64 B 0.031754f
C276 VP.n65 B 0.024229f
C277 VP.n66 B 0.027366f
C278 VP.n67 B 1.29845f
C279 VP.t8 B 2.74352f
C280 VP.n68 B 1.01851f
C281 VP.n69 B 1.30826f
C282 VP.n70 B 0.027366f
C283 VP.n71 B 0.016953f
C284 VP.n72 B 0.031754f
C285 VP.n73 B 0.031754f
C286 VP.n74 B 0.021525f
C287 VP.n75 B 0.016953f
C288 VP.n76 B 0.016953f
C289 VP.n77 B 0.016953f
C290 VP.n78 B 0.031754f
C291 VP.n79 B 0.031754f
C292 VP.n80 B 0.019839f
C293 VP.n81 B 0.016953f
C294 VP.n82 B 0.016953f
C295 VP.n83 B 0.027991f
C296 VP.n84 B 0.031754f
C297 VP.n85 B 0.034444f
C298 VP.n86 B 0.016953f
C299 VP.n87 B 0.016953f
C300 VP.n88 B 0.016953f
C301 VP.n89 B 0.032497f
C302 VP.n90 B 0.031754f
C303 VP.n91 B 0.031754f
C304 VP.n92 B 0.016953f
C305 VP.n93 B 0.016953f
C306 VP.n94 B 0.016953f
C307 VP.n95 B 0.031754f
C308 VP.n96 B 0.031754f
C309 VP.n97 B 0.032497f
C310 VP.n98 B 0.016953f
C311 VP.n99 B 0.016953f
C312 VP.n100 B 0.016953f
C313 VP.n101 B 0.034444f
C314 VP.n102 B 0.031754f
C315 VP.t3 B 2.74352f
C316 VP.n103 B 0.948923f
C317 VP.n104 B 0.027991f
C318 VP.n105 B 0.016953f
C319 VP.n106 B 0.016953f
C320 VP.n107 B 0.016953f
C321 VP.n108 B 0.031754f
C322 VP.n109 B 0.031754f
C323 VP.n110 B 0.028186f
C324 VP.n111 B 0.016953f
C325 VP.n112 B 0.016953f
C326 VP.n113 B 0.016953f
C327 VP.n114 B 0.031754f
C328 VP.n115 B 0.031754f
C329 VP.n116 B 0.024229f
C330 VP.n117 B 0.027366f
C331 VP.n118 B 0.044211f
.ends

