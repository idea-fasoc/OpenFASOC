* NGSPICE file created from diff_pair_sample_1023.ext - technology: sky130A

.subckt diff_pair_sample_1023 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=3.73
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=3.73
X2 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=3.73
X3 VDD1.t2 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=3.73
X4 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=3.73
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=3.73
X6 VTAIL.t6 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=3.73
X7 VDD2.t1 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=3.73
X8 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0032 pd=6.41 as=2.3712 ps=12.94 w=6.08 l=3.73
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=3.73
X10 VTAIL.t5 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=1.0032 ps=6.41 w=6.08 l=3.73
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3712 pd=12.94 as=0 ps=0 w=6.08 l=3.73
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n7 VP.n6 88.77
R10 VP.n22 VP.n0 88.77
R11 VP.n5 VP.t2 72.841
R12 VP.n5 VP.t0 71.5072
R13 VP.n6 VP.n5 47.1985
R14 VP.n14 VP.n13 40.577
R15 VP.n14 VP.n2 40.577
R16 VP.n7 VP.t3 39.2841
R17 VP.n0 VP.t1 39.2841
R18 VP.n8 VP.n4 24.5923
R19 VP.n12 VP.n4 24.5923
R20 VP.n13 VP.n12 24.5923
R21 VP.n18 VP.n2 24.5923
R22 VP.n19 VP.n18 24.5923
R23 VP.n20 VP.n19 24.5923
R24 VP.n8 VP.n7 1.47601
R25 VP.n20 VP.n0 1.47601
R26 VP.n9 VP.n6 0.354861
R27 VP.n22 VP.n21 0.354861
R28 VP VP.n22 0.267071
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VTAIL.n250 VTAIL.n224 289.615
R38 VTAIL.n26 VTAIL.n0 289.615
R39 VTAIL.n58 VTAIL.n32 289.615
R40 VTAIL.n90 VTAIL.n64 289.615
R41 VTAIL.n218 VTAIL.n192 289.615
R42 VTAIL.n186 VTAIL.n160 289.615
R43 VTAIL.n154 VTAIL.n128 289.615
R44 VTAIL.n122 VTAIL.n96 289.615
R45 VTAIL.n235 VTAIL.n234 185
R46 VTAIL.n232 VTAIL.n231 185
R47 VTAIL.n241 VTAIL.n240 185
R48 VTAIL.n243 VTAIL.n242 185
R49 VTAIL.n228 VTAIL.n227 185
R50 VTAIL.n249 VTAIL.n248 185
R51 VTAIL.n251 VTAIL.n250 185
R52 VTAIL.n11 VTAIL.n10 185
R53 VTAIL.n8 VTAIL.n7 185
R54 VTAIL.n17 VTAIL.n16 185
R55 VTAIL.n19 VTAIL.n18 185
R56 VTAIL.n4 VTAIL.n3 185
R57 VTAIL.n25 VTAIL.n24 185
R58 VTAIL.n27 VTAIL.n26 185
R59 VTAIL.n43 VTAIL.n42 185
R60 VTAIL.n40 VTAIL.n39 185
R61 VTAIL.n49 VTAIL.n48 185
R62 VTAIL.n51 VTAIL.n50 185
R63 VTAIL.n36 VTAIL.n35 185
R64 VTAIL.n57 VTAIL.n56 185
R65 VTAIL.n59 VTAIL.n58 185
R66 VTAIL.n75 VTAIL.n74 185
R67 VTAIL.n72 VTAIL.n71 185
R68 VTAIL.n81 VTAIL.n80 185
R69 VTAIL.n83 VTAIL.n82 185
R70 VTAIL.n68 VTAIL.n67 185
R71 VTAIL.n89 VTAIL.n88 185
R72 VTAIL.n91 VTAIL.n90 185
R73 VTAIL.n219 VTAIL.n218 185
R74 VTAIL.n217 VTAIL.n216 185
R75 VTAIL.n196 VTAIL.n195 185
R76 VTAIL.n211 VTAIL.n210 185
R77 VTAIL.n209 VTAIL.n208 185
R78 VTAIL.n200 VTAIL.n199 185
R79 VTAIL.n203 VTAIL.n202 185
R80 VTAIL.n187 VTAIL.n186 185
R81 VTAIL.n185 VTAIL.n184 185
R82 VTAIL.n164 VTAIL.n163 185
R83 VTAIL.n179 VTAIL.n178 185
R84 VTAIL.n177 VTAIL.n176 185
R85 VTAIL.n168 VTAIL.n167 185
R86 VTAIL.n171 VTAIL.n170 185
R87 VTAIL.n155 VTAIL.n154 185
R88 VTAIL.n153 VTAIL.n152 185
R89 VTAIL.n132 VTAIL.n131 185
R90 VTAIL.n147 VTAIL.n146 185
R91 VTAIL.n145 VTAIL.n144 185
R92 VTAIL.n136 VTAIL.n135 185
R93 VTAIL.n139 VTAIL.n138 185
R94 VTAIL.n123 VTAIL.n122 185
R95 VTAIL.n121 VTAIL.n120 185
R96 VTAIL.n100 VTAIL.n99 185
R97 VTAIL.n115 VTAIL.n114 185
R98 VTAIL.n113 VTAIL.n112 185
R99 VTAIL.n104 VTAIL.n103 185
R100 VTAIL.n107 VTAIL.n106 185
R101 VTAIL.t7 VTAIL.n233 147.661
R102 VTAIL.t0 VTAIL.n9 147.661
R103 VTAIL.t3 VTAIL.n41 147.661
R104 VTAIL.t5 VTAIL.n73 147.661
R105 VTAIL.t4 VTAIL.n201 147.661
R106 VTAIL.t6 VTAIL.n169 147.661
R107 VTAIL.t1 VTAIL.n137 147.661
R108 VTAIL.t2 VTAIL.n105 147.661
R109 VTAIL.n234 VTAIL.n231 104.615
R110 VTAIL.n241 VTAIL.n231 104.615
R111 VTAIL.n242 VTAIL.n241 104.615
R112 VTAIL.n242 VTAIL.n227 104.615
R113 VTAIL.n249 VTAIL.n227 104.615
R114 VTAIL.n250 VTAIL.n249 104.615
R115 VTAIL.n10 VTAIL.n7 104.615
R116 VTAIL.n17 VTAIL.n7 104.615
R117 VTAIL.n18 VTAIL.n17 104.615
R118 VTAIL.n18 VTAIL.n3 104.615
R119 VTAIL.n25 VTAIL.n3 104.615
R120 VTAIL.n26 VTAIL.n25 104.615
R121 VTAIL.n42 VTAIL.n39 104.615
R122 VTAIL.n49 VTAIL.n39 104.615
R123 VTAIL.n50 VTAIL.n49 104.615
R124 VTAIL.n50 VTAIL.n35 104.615
R125 VTAIL.n57 VTAIL.n35 104.615
R126 VTAIL.n58 VTAIL.n57 104.615
R127 VTAIL.n74 VTAIL.n71 104.615
R128 VTAIL.n81 VTAIL.n71 104.615
R129 VTAIL.n82 VTAIL.n81 104.615
R130 VTAIL.n82 VTAIL.n67 104.615
R131 VTAIL.n89 VTAIL.n67 104.615
R132 VTAIL.n90 VTAIL.n89 104.615
R133 VTAIL.n218 VTAIL.n217 104.615
R134 VTAIL.n217 VTAIL.n195 104.615
R135 VTAIL.n210 VTAIL.n195 104.615
R136 VTAIL.n210 VTAIL.n209 104.615
R137 VTAIL.n209 VTAIL.n199 104.615
R138 VTAIL.n202 VTAIL.n199 104.615
R139 VTAIL.n186 VTAIL.n185 104.615
R140 VTAIL.n185 VTAIL.n163 104.615
R141 VTAIL.n178 VTAIL.n163 104.615
R142 VTAIL.n178 VTAIL.n177 104.615
R143 VTAIL.n177 VTAIL.n167 104.615
R144 VTAIL.n170 VTAIL.n167 104.615
R145 VTAIL.n154 VTAIL.n153 104.615
R146 VTAIL.n153 VTAIL.n131 104.615
R147 VTAIL.n146 VTAIL.n131 104.615
R148 VTAIL.n146 VTAIL.n145 104.615
R149 VTAIL.n145 VTAIL.n135 104.615
R150 VTAIL.n138 VTAIL.n135 104.615
R151 VTAIL.n122 VTAIL.n121 104.615
R152 VTAIL.n121 VTAIL.n99 104.615
R153 VTAIL.n114 VTAIL.n99 104.615
R154 VTAIL.n114 VTAIL.n113 104.615
R155 VTAIL.n113 VTAIL.n103 104.615
R156 VTAIL.n106 VTAIL.n103 104.615
R157 VTAIL.n234 VTAIL.t7 52.3082
R158 VTAIL.n10 VTAIL.t0 52.3082
R159 VTAIL.n42 VTAIL.t3 52.3082
R160 VTAIL.n74 VTAIL.t5 52.3082
R161 VTAIL.n202 VTAIL.t4 52.3082
R162 VTAIL.n170 VTAIL.t6 52.3082
R163 VTAIL.n138 VTAIL.t1 52.3082
R164 VTAIL.n106 VTAIL.t2 52.3082
R165 VTAIL.n255 VTAIL.n254 33.7369
R166 VTAIL.n31 VTAIL.n30 33.7369
R167 VTAIL.n63 VTAIL.n62 33.7369
R168 VTAIL.n95 VTAIL.n94 33.7369
R169 VTAIL.n223 VTAIL.n222 33.7369
R170 VTAIL.n191 VTAIL.n190 33.7369
R171 VTAIL.n159 VTAIL.n158 33.7369
R172 VTAIL.n127 VTAIL.n126 33.7369
R173 VTAIL.n255 VTAIL.n223 21.1083
R174 VTAIL.n127 VTAIL.n95 21.1083
R175 VTAIL.n235 VTAIL.n233 15.6674
R176 VTAIL.n11 VTAIL.n9 15.6674
R177 VTAIL.n43 VTAIL.n41 15.6674
R178 VTAIL.n75 VTAIL.n73 15.6674
R179 VTAIL.n203 VTAIL.n201 15.6674
R180 VTAIL.n171 VTAIL.n169 15.6674
R181 VTAIL.n139 VTAIL.n137 15.6674
R182 VTAIL.n107 VTAIL.n105 15.6674
R183 VTAIL.n236 VTAIL.n232 12.8005
R184 VTAIL.n12 VTAIL.n8 12.8005
R185 VTAIL.n44 VTAIL.n40 12.8005
R186 VTAIL.n76 VTAIL.n72 12.8005
R187 VTAIL.n204 VTAIL.n200 12.8005
R188 VTAIL.n172 VTAIL.n168 12.8005
R189 VTAIL.n140 VTAIL.n136 12.8005
R190 VTAIL.n108 VTAIL.n104 12.8005
R191 VTAIL.n240 VTAIL.n239 12.0247
R192 VTAIL.n16 VTAIL.n15 12.0247
R193 VTAIL.n48 VTAIL.n47 12.0247
R194 VTAIL.n80 VTAIL.n79 12.0247
R195 VTAIL.n208 VTAIL.n207 12.0247
R196 VTAIL.n176 VTAIL.n175 12.0247
R197 VTAIL.n144 VTAIL.n143 12.0247
R198 VTAIL.n112 VTAIL.n111 12.0247
R199 VTAIL.n243 VTAIL.n230 11.249
R200 VTAIL.n19 VTAIL.n6 11.249
R201 VTAIL.n51 VTAIL.n38 11.249
R202 VTAIL.n83 VTAIL.n70 11.249
R203 VTAIL.n211 VTAIL.n198 11.249
R204 VTAIL.n179 VTAIL.n166 11.249
R205 VTAIL.n147 VTAIL.n134 11.249
R206 VTAIL.n115 VTAIL.n102 11.249
R207 VTAIL.n244 VTAIL.n228 10.4732
R208 VTAIL.n20 VTAIL.n4 10.4732
R209 VTAIL.n52 VTAIL.n36 10.4732
R210 VTAIL.n84 VTAIL.n68 10.4732
R211 VTAIL.n212 VTAIL.n196 10.4732
R212 VTAIL.n180 VTAIL.n164 10.4732
R213 VTAIL.n148 VTAIL.n132 10.4732
R214 VTAIL.n116 VTAIL.n100 10.4732
R215 VTAIL.n248 VTAIL.n247 9.69747
R216 VTAIL.n24 VTAIL.n23 9.69747
R217 VTAIL.n56 VTAIL.n55 9.69747
R218 VTAIL.n88 VTAIL.n87 9.69747
R219 VTAIL.n216 VTAIL.n215 9.69747
R220 VTAIL.n184 VTAIL.n183 9.69747
R221 VTAIL.n152 VTAIL.n151 9.69747
R222 VTAIL.n120 VTAIL.n119 9.69747
R223 VTAIL.n254 VTAIL.n253 9.45567
R224 VTAIL.n30 VTAIL.n29 9.45567
R225 VTAIL.n62 VTAIL.n61 9.45567
R226 VTAIL.n94 VTAIL.n93 9.45567
R227 VTAIL.n222 VTAIL.n221 9.45567
R228 VTAIL.n190 VTAIL.n189 9.45567
R229 VTAIL.n158 VTAIL.n157 9.45567
R230 VTAIL.n126 VTAIL.n125 9.45567
R231 VTAIL.n253 VTAIL.n252 9.3005
R232 VTAIL.n226 VTAIL.n225 9.3005
R233 VTAIL.n247 VTAIL.n246 9.3005
R234 VTAIL.n245 VTAIL.n244 9.3005
R235 VTAIL.n230 VTAIL.n229 9.3005
R236 VTAIL.n239 VTAIL.n238 9.3005
R237 VTAIL.n237 VTAIL.n236 9.3005
R238 VTAIL.n29 VTAIL.n28 9.3005
R239 VTAIL.n2 VTAIL.n1 9.3005
R240 VTAIL.n23 VTAIL.n22 9.3005
R241 VTAIL.n21 VTAIL.n20 9.3005
R242 VTAIL.n6 VTAIL.n5 9.3005
R243 VTAIL.n15 VTAIL.n14 9.3005
R244 VTAIL.n13 VTAIL.n12 9.3005
R245 VTAIL.n61 VTAIL.n60 9.3005
R246 VTAIL.n34 VTAIL.n33 9.3005
R247 VTAIL.n55 VTAIL.n54 9.3005
R248 VTAIL.n53 VTAIL.n52 9.3005
R249 VTAIL.n38 VTAIL.n37 9.3005
R250 VTAIL.n47 VTAIL.n46 9.3005
R251 VTAIL.n45 VTAIL.n44 9.3005
R252 VTAIL.n93 VTAIL.n92 9.3005
R253 VTAIL.n66 VTAIL.n65 9.3005
R254 VTAIL.n87 VTAIL.n86 9.3005
R255 VTAIL.n85 VTAIL.n84 9.3005
R256 VTAIL.n70 VTAIL.n69 9.3005
R257 VTAIL.n79 VTAIL.n78 9.3005
R258 VTAIL.n77 VTAIL.n76 9.3005
R259 VTAIL.n221 VTAIL.n220 9.3005
R260 VTAIL.n194 VTAIL.n193 9.3005
R261 VTAIL.n215 VTAIL.n214 9.3005
R262 VTAIL.n213 VTAIL.n212 9.3005
R263 VTAIL.n198 VTAIL.n197 9.3005
R264 VTAIL.n207 VTAIL.n206 9.3005
R265 VTAIL.n205 VTAIL.n204 9.3005
R266 VTAIL.n189 VTAIL.n188 9.3005
R267 VTAIL.n162 VTAIL.n161 9.3005
R268 VTAIL.n183 VTAIL.n182 9.3005
R269 VTAIL.n181 VTAIL.n180 9.3005
R270 VTAIL.n166 VTAIL.n165 9.3005
R271 VTAIL.n175 VTAIL.n174 9.3005
R272 VTAIL.n173 VTAIL.n172 9.3005
R273 VTAIL.n157 VTAIL.n156 9.3005
R274 VTAIL.n130 VTAIL.n129 9.3005
R275 VTAIL.n151 VTAIL.n150 9.3005
R276 VTAIL.n149 VTAIL.n148 9.3005
R277 VTAIL.n134 VTAIL.n133 9.3005
R278 VTAIL.n143 VTAIL.n142 9.3005
R279 VTAIL.n141 VTAIL.n140 9.3005
R280 VTAIL.n125 VTAIL.n124 9.3005
R281 VTAIL.n98 VTAIL.n97 9.3005
R282 VTAIL.n119 VTAIL.n118 9.3005
R283 VTAIL.n117 VTAIL.n116 9.3005
R284 VTAIL.n102 VTAIL.n101 9.3005
R285 VTAIL.n111 VTAIL.n110 9.3005
R286 VTAIL.n109 VTAIL.n108 9.3005
R287 VTAIL.n251 VTAIL.n226 8.92171
R288 VTAIL.n27 VTAIL.n2 8.92171
R289 VTAIL.n59 VTAIL.n34 8.92171
R290 VTAIL.n91 VTAIL.n66 8.92171
R291 VTAIL.n219 VTAIL.n194 8.92171
R292 VTAIL.n187 VTAIL.n162 8.92171
R293 VTAIL.n155 VTAIL.n130 8.92171
R294 VTAIL.n123 VTAIL.n98 8.92171
R295 VTAIL.n252 VTAIL.n224 8.14595
R296 VTAIL.n28 VTAIL.n0 8.14595
R297 VTAIL.n60 VTAIL.n32 8.14595
R298 VTAIL.n92 VTAIL.n64 8.14595
R299 VTAIL.n220 VTAIL.n192 8.14595
R300 VTAIL.n188 VTAIL.n160 8.14595
R301 VTAIL.n156 VTAIL.n128 8.14595
R302 VTAIL.n124 VTAIL.n96 8.14595
R303 VTAIL.n254 VTAIL.n224 5.81868
R304 VTAIL.n30 VTAIL.n0 5.81868
R305 VTAIL.n62 VTAIL.n32 5.81868
R306 VTAIL.n94 VTAIL.n64 5.81868
R307 VTAIL.n222 VTAIL.n192 5.81868
R308 VTAIL.n190 VTAIL.n160 5.81868
R309 VTAIL.n158 VTAIL.n128 5.81868
R310 VTAIL.n126 VTAIL.n96 5.81868
R311 VTAIL.n252 VTAIL.n251 5.04292
R312 VTAIL.n28 VTAIL.n27 5.04292
R313 VTAIL.n60 VTAIL.n59 5.04292
R314 VTAIL.n92 VTAIL.n91 5.04292
R315 VTAIL.n220 VTAIL.n219 5.04292
R316 VTAIL.n188 VTAIL.n187 5.04292
R317 VTAIL.n156 VTAIL.n155 5.04292
R318 VTAIL.n124 VTAIL.n123 5.04292
R319 VTAIL.n237 VTAIL.n233 4.38594
R320 VTAIL.n13 VTAIL.n9 4.38594
R321 VTAIL.n45 VTAIL.n41 4.38594
R322 VTAIL.n77 VTAIL.n73 4.38594
R323 VTAIL.n205 VTAIL.n201 4.38594
R324 VTAIL.n173 VTAIL.n169 4.38594
R325 VTAIL.n141 VTAIL.n137 4.38594
R326 VTAIL.n109 VTAIL.n105 4.38594
R327 VTAIL.n248 VTAIL.n226 4.26717
R328 VTAIL.n24 VTAIL.n2 4.26717
R329 VTAIL.n56 VTAIL.n34 4.26717
R330 VTAIL.n88 VTAIL.n66 4.26717
R331 VTAIL.n216 VTAIL.n194 4.26717
R332 VTAIL.n184 VTAIL.n162 4.26717
R333 VTAIL.n152 VTAIL.n130 4.26717
R334 VTAIL.n120 VTAIL.n98 4.26717
R335 VTAIL.n159 VTAIL.n127 3.5005
R336 VTAIL.n223 VTAIL.n191 3.5005
R337 VTAIL.n95 VTAIL.n63 3.5005
R338 VTAIL.n247 VTAIL.n228 3.49141
R339 VTAIL.n23 VTAIL.n4 3.49141
R340 VTAIL.n55 VTAIL.n36 3.49141
R341 VTAIL.n87 VTAIL.n68 3.49141
R342 VTAIL.n215 VTAIL.n196 3.49141
R343 VTAIL.n183 VTAIL.n164 3.49141
R344 VTAIL.n151 VTAIL.n132 3.49141
R345 VTAIL.n119 VTAIL.n100 3.49141
R346 VTAIL.n244 VTAIL.n243 2.71565
R347 VTAIL.n20 VTAIL.n19 2.71565
R348 VTAIL.n52 VTAIL.n51 2.71565
R349 VTAIL.n84 VTAIL.n83 2.71565
R350 VTAIL.n212 VTAIL.n211 2.71565
R351 VTAIL.n180 VTAIL.n179 2.71565
R352 VTAIL.n148 VTAIL.n147 2.71565
R353 VTAIL.n116 VTAIL.n115 2.71565
R354 VTAIL.n240 VTAIL.n230 1.93989
R355 VTAIL.n16 VTAIL.n6 1.93989
R356 VTAIL.n48 VTAIL.n38 1.93989
R357 VTAIL.n80 VTAIL.n70 1.93989
R358 VTAIL.n208 VTAIL.n198 1.93989
R359 VTAIL.n176 VTAIL.n166 1.93989
R360 VTAIL.n144 VTAIL.n134 1.93989
R361 VTAIL.n112 VTAIL.n102 1.93989
R362 VTAIL VTAIL.n31 1.80869
R363 VTAIL VTAIL.n255 1.69231
R364 VTAIL.n239 VTAIL.n232 1.16414
R365 VTAIL.n15 VTAIL.n8 1.16414
R366 VTAIL.n47 VTAIL.n40 1.16414
R367 VTAIL.n79 VTAIL.n72 1.16414
R368 VTAIL.n207 VTAIL.n200 1.16414
R369 VTAIL.n175 VTAIL.n168 1.16414
R370 VTAIL.n143 VTAIL.n136 1.16414
R371 VTAIL.n111 VTAIL.n104 1.16414
R372 VTAIL.n191 VTAIL.n159 0.470328
R373 VTAIL.n63 VTAIL.n31 0.470328
R374 VTAIL.n236 VTAIL.n235 0.388379
R375 VTAIL.n12 VTAIL.n11 0.388379
R376 VTAIL.n44 VTAIL.n43 0.388379
R377 VTAIL.n76 VTAIL.n75 0.388379
R378 VTAIL.n204 VTAIL.n203 0.388379
R379 VTAIL.n172 VTAIL.n171 0.388379
R380 VTAIL.n140 VTAIL.n139 0.388379
R381 VTAIL.n108 VTAIL.n107 0.388379
R382 VTAIL.n238 VTAIL.n237 0.155672
R383 VTAIL.n238 VTAIL.n229 0.155672
R384 VTAIL.n245 VTAIL.n229 0.155672
R385 VTAIL.n246 VTAIL.n245 0.155672
R386 VTAIL.n246 VTAIL.n225 0.155672
R387 VTAIL.n253 VTAIL.n225 0.155672
R388 VTAIL.n14 VTAIL.n13 0.155672
R389 VTAIL.n14 VTAIL.n5 0.155672
R390 VTAIL.n21 VTAIL.n5 0.155672
R391 VTAIL.n22 VTAIL.n21 0.155672
R392 VTAIL.n22 VTAIL.n1 0.155672
R393 VTAIL.n29 VTAIL.n1 0.155672
R394 VTAIL.n46 VTAIL.n45 0.155672
R395 VTAIL.n46 VTAIL.n37 0.155672
R396 VTAIL.n53 VTAIL.n37 0.155672
R397 VTAIL.n54 VTAIL.n53 0.155672
R398 VTAIL.n54 VTAIL.n33 0.155672
R399 VTAIL.n61 VTAIL.n33 0.155672
R400 VTAIL.n78 VTAIL.n77 0.155672
R401 VTAIL.n78 VTAIL.n69 0.155672
R402 VTAIL.n85 VTAIL.n69 0.155672
R403 VTAIL.n86 VTAIL.n85 0.155672
R404 VTAIL.n86 VTAIL.n65 0.155672
R405 VTAIL.n93 VTAIL.n65 0.155672
R406 VTAIL.n221 VTAIL.n193 0.155672
R407 VTAIL.n214 VTAIL.n193 0.155672
R408 VTAIL.n214 VTAIL.n213 0.155672
R409 VTAIL.n213 VTAIL.n197 0.155672
R410 VTAIL.n206 VTAIL.n197 0.155672
R411 VTAIL.n206 VTAIL.n205 0.155672
R412 VTAIL.n189 VTAIL.n161 0.155672
R413 VTAIL.n182 VTAIL.n161 0.155672
R414 VTAIL.n182 VTAIL.n181 0.155672
R415 VTAIL.n181 VTAIL.n165 0.155672
R416 VTAIL.n174 VTAIL.n165 0.155672
R417 VTAIL.n174 VTAIL.n173 0.155672
R418 VTAIL.n157 VTAIL.n129 0.155672
R419 VTAIL.n150 VTAIL.n129 0.155672
R420 VTAIL.n150 VTAIL.n149 0.155672
R421 VTAIL.n149 VTAIL.n133 0.155672
R422 VTAIL.n142 VTAIL.n133 0.155672
R423 VTAIL.n142 VTAIL.n141 0.155672
R424 VTAIL.n125 VTAIL.n97 0.155672
R425 VTAIL.n118 VTAIL.n97 0.155672
R426 VTAIL.n118 VTAIL.n117 0.155672
R427 VTAIL.n117 VTAIL.n101 0.155672
R428 VTAIL.n110 VTAIL.n101 0.155672
R429 VTAIL.n110 VTAIL.n109 0.155672
R430 VDD1 VDD1.n1 108.724
R431 VDD1 VDD1.n0 68.8004
R432 VDD1.n0 VDD1.t1 3.25708
R433 VDD1.n0 VDD1.t3 3.25708
R434 VDD1.n1 VDD1.t0 3.25708
R435 VDD1.n1 VDD1.t2 3.25708
R436 B.n654 B.n653 585
R437 B.n228 B.n111 585
R438 B.n227 B.n226 585
R439 B.n225 B.n224 585
R440 B.n223 B.n222 585
R441 B.n221 B.n220 585
R442 B.n219 B.n218 585
R443 B.n217 B.n216 585
R444 B.n215 B.n214 585
R445 B.n213 B.n212 585
R446 B.n211 B.n210 585
R447 B.n209 B.n208 585
R448 B.n207 B.n206 585
R449 B.n205 B.n204 585
R450 B.n203 B.n202 585
R451 B.n201 B.n200 585
R452 B.n199 B.n198 585
R453 B.n197 B.n196 585
R454 B.n195 B.n194 585
R455 B.n193 B.n192 585
R456 B.n191 B.n190 585
R457 B.n189 B.n188 585
R458 B.n187 B.n186 585
R459 B.n185 B.n184 585
R460 B.n183 B.n182 585
R461 B.n181 B.n180 585
R462 B.n179 B.n178 585
R463 B.n177 B.n176 585
R464 B.n175 B.n174 585
R465 B.n173 B.n172 585
R466 B.n171 B.n170 585
R467 B.n169 B.n168 585
R468 B.n167 B.n166 585
R469 B.n165 B.n164 585
R470 B.n163 B.n162 585
R471 B.n161 B.n160 585
R472 B.n159 B.n158 585
R473 B.n157 B.n156 585
R474 B.n155 B.n154 585
R475 B.n153 B.n152 585
R476 B.n151 B.n150 585
R477 B.n149 B.n148 585
R478 B.n147 B.n146 585
R479 B.n145 B.n144 585
R480 B.n143 B.n142 585
R481 B.n141 B.n140 585
R482 B.n139 B.n138 585
R483 B.n137 B.n136 585
R484 B.n135 B.n134 585
R485 B.n133 B.n132 585
R486 B.n131 B.n130 585
R487 B.n129 B.n128 585
R488 B.n127 B.n126 585
R489 B.n125 B.n124 585
R490 B.n123 B.n122 585
R491 B.n121 B.n120 585
R492 B.n119 B.n118 585
R493 B.n81 B.n80 585
R494 B.n652 B.n82 585
R495 B.n657 B.n82 585
R496 B.n651 B.n650 585
R497 B.n650 B.n78 585
R498 B.n649 B.n77 585
R499 B.n663 B.n77 585
R500 B.n648 B.n76 585
R501 B.n664 B.n76 585
R502 B.n647 B.n75 585
R503 B.n665 B.n75 585
R504 B.n646 B.n645 585
R505 B.n645 B.n71 585
R506 B.n644 B.n70 585
R507 B.n671 B.n70 585
R508 B.n643 B.n69 585
R509 B.n672 B.n69 585
R510 B.n642 B.n68 585
R511 B.n673 B.n68 585
R512 B.n641 B.n640 585
R513 B.n640 B.n67 585
R514 B.n639 B.n63 585
R515 B.n679 B.n63 585
R516 B.n638 B.n62 585
R517 B.n680 B.n62 585
R518 B.n637 B.n61 585
R519 B.n681 B.n61 585
R520 B.n636 B.n635 585
R521 B.n635 B.n57 585
R522 B.n634 B.n56 585
R523 B.n687 B.n56 585
R524 B.n633 B.n55 585
R525 B.n688 B.n55 585
R526 B.n632 B.n54 585
R527 B.n689 B.n54 585
R528 B.n631 B.n630 585
R529 B.n630 B.n50 585
R530 B.n629 B.n49 585
R531 B.n695 B.n49 585
R532 B.n628 B.n48 585
R533 B.n696 B.n48 585
R534 B.n627 B.n47 585
R535 B.n697 B.n47 585
R536 B.n626 B.n625 585
R537 B.n625 B.n43 585
R538 B.n624 B.n42 585
R539 B.n703 B.n42 585
R540 B.n623 B.n41 585
R541 B.n704 B.n41 585
R542 B.n622 B.n40 585
R543 B.n705 B.n40 585
R544 B.n621 B.n620 585
R545 B.n620 B.n36 585
R546 B.n619 B.n35 585
R547 B.n711 B.n35 585
R548 B.n618 B.n34 585
R549 B.n712 B.n34 585
R550 B.n617 B.n33 585
R551 B.n713 B.n33 585
R552 B.n616 B.n615 585
R553 B.n615 B.n29 585
R554 B.n614 B.n28 585
R555 B.n719 B.n28 585
R556 B.n613 B.n27 585
R557 B.n720 B.n27 585
R558 B.n612 B.n26 585
R559 B.n721 B.n26 585
R560 B.n611 B.n610 585
R561 B.n610 B.n22 585
R562 B.n609 B.n21 585
R563 B.n727 B.n21 585
R564 B.n608 B.n20 585
R565 B.n728 B.n20 585
R566 B.n607 B.n19 585
R567 B.n729 B.n19 585
R568 B.n606 B.n605 585
R569 B.n605 B.n15 585
R570 B.n604 B.n14 585
R571 B.n735 B.n14 585
R572 B.n603 B.n13 585
R573 B.n736 B.n13 585
R574 B.n602 B.n12 585
R575 B.n737 B.n12 585
R576 B.n601 B.n600 585
R577 B.n600 B.n8 585
R578 B.n599 B.n7 585
R579 B.n743 B.n7 585
R580 B.n598 B.n6 585
R581 B.n744 B.n6 585
R582 B.n597 B.n5 585
R583 B.n745 B.n5 585
R584 B.n596 B.n595 585
R585 B.n595 B.n4 585
R586 B.n594 B.n229 585
R587 B.n594 B.n593 585
R588 B.n584 B.n230 585
R589 B.n231 B.n230 585
R590 B.n586 B.n585 585
R591 B.n587 B.n586 585
R592 B.n583 B.n236 585
R593 B.n236 B.n235 585
R594 B.n582 B.n581 585
R595 B.n581 B.n580 585
R596 B.n238 B.n237 585
R597 B.n239 B.n238 585
R598 B.n573 B.n572 585
R599 B.n574 B.n573 585
R600 B.n571 B.n244 585
R601 B.n244 B.n243 585
R602 B.n570 B.n569 585
R603 B.n569 B.n568 585
R604 B.n246 B.n245 585
R605 B.n247 B.n246 585
R606 B.n561 B.n560 585
R607 B.n562 B.n561 585
R608 B.n559 B.n252 585
R609 B.n252 B.n251 585
R610 B.n558 B.n557 585
R611 B.n557 B.n556 585
R612 B.n254 B.n253 585
R613 B.n255 B.n254 585
R614 B.n549 B.n548 585
R615 B.n550 B.n549 585
R616 B.n547 B.n260 585
R617 B.n260 B.n259 585
R618 B.n546 B.n545 585
R619 B.n545 B.n544 585
R620 B.n262 B.n261 585
R621 B.n263 B.n262 585
R622 B.n537 B.n536 585
R623 B.n538 B.n537 585
R624 B.n535 B.n268 585
R625 B.n268 B.n267 585
R626 B.n534 B.n533 585
R627 B.n533 B.n532 585
R628 B.n270 B.n269 585
R629 B.n271 B.n270 585
R630 B.n525 B.n524 585
R631 B.n526 B.n525 585
R632 B.n523 B.n276 585
R633 B.n276 B.n275 585
R634 B.n522 B.n521 585
R635 B.n521 B.n520 585
R636 B.n278 B.n277 585
R637 B.n279 B.n278 585
R638 B.n513 B.n512 585
R639 B.n514 B.n513 585
R640 B.n511 B.n284 585
R641 B.n284 B.n283 585
R642 B.n510 B.n509 585
R643 B.n509 B.n508 585
R644 B.n286 B.n285 585
R645 B.n287 B.n286 585
R646 B.n501 B.n500 585
R647 B.n502 B.n501 585
R648 B.n499 B.n292 585
R649 B.n292 B.n291 585
R650 B.n498 B.n497 585
R651 B.n497 B.n496 585
R652 B.n294 B.n293 585
R653 B.n489 B.n294 585
R654 B.n488 B.n487 585
R655 B.n490 B.n488 585
R656 B.n486 B.n299 585
R657 B.n299 B.n298 585
R658 B.n485 B.n484 585
R659 B.n484 B.n483 585
R660 B.n301 B.n300 585
R661 B.n302 B.n301 585
R662 B.n476 B.n475 585
R663 B.n477 B.n476 585
R664 B.n474 B.n307 585
R665 B.n307 B.n306 585
R666 B.n473 B.n472 585
R667 B.n472 B.n471 585
R668 B.n309 B.n308 585
R669 B.n310 B.n309 585
R670 B.n464 B.n463 585
R671 B.n465 B.n464 585
R672 B.n313 B.n312 585
R673 B.n348 B.n346 585
R674 B.n349 B.n345 585
R675 B.n349 B.n314 585
R676 B.n352 B.n351 585
R677 B.n353 B.n344 585
R678 B.n355 B.n354 585
R679 B.n357 B.n343 585
R680 B.n360 B.n359 585
R681 B.n361 B.n342 585
R682 B.n363 B.n362 585
R683 B.n365 B.n341 585
R684 B.n368 B.n367 585
R685 B.n369 B.n340 585
R686 B.n371 B.n370 585
R687 B.n373 B.n339 585
R688 B.n376 B.n375 585
R689 B.n377 B.n338 585
R690 B.n379 B.n378 585
R691 B.n381 B.n337 585
R692 B.n384 B.n383 585
R693 B.n385 B.n336 585
R694 B.n387 B.n386 585
R695 B.n389 B.n335 585
R696 B.n392 B.n391 585
R697 B.n394 B.n332 585
R698 B.n396 B.n395 585
R699 B.n398 B.n331 585
R700 B.n401 B.n400 585
R701 B.n402 B.n330 585
R702 B.n404 B.n403 585
R703 B.n406 B.n329 585
R704 B.n409 B.n408 585
R705 B.n410 B.n328 585
R706 B.n415 B.n414 585
R707 B.n417 B.n327 585
R708 B.n420 B.n419 585
R709 B.n421 B.n326 585
R710 B.n423 B.n422 585
R711 B.n425 B.n325 585
R712 B.n428 B.n427 585
R713 B.n429 B.n324 585
R714 B.n431 B.n430 585
R715 B.n433 B.n323 585
R716 B.n436 B.n435 585
R717 B.n437 B.n322 585
R718 B.n439 B.n438 585
R719 B.n441 B.n321 585
R720 B.n444 B.n443 585
R721 B.n445 B.n320 585
R722 B.n447 B.n446 585
R723 B.n449 B.n319 585
R724 B.n452 B.n451 585
R725 B.n453 B.n318 585
R726 B.n455 B.n454 585
R727 B.n457 B.n317 585
R728 B.n458 B.n316 585
R729 B.n461 B.n460 585
R730 B.n462 B.n315 585
R731 B.n315 B.n314 585
R732 B.n467 B.n466 585
R733 B.n466 B.n465 585
R734 B.n468 B.n311 585
R735 B.n311 B.n310 585
R736 B.n470 B.n469 585
R737 B.n471 B.n470 585
R738 B.n305 B.n304 585
R739 B.n306 B.n305 585
R740 B.n479 B.n478 585
R741 B.n478 B.n477 585
R742 B.n480 B.n303 585
R743 B.n303 B.n302 585
R744 B.n482 B.n481 585
R745 B.n483 B.n482 585
R746 B.n297 B.n296 585
R747 B.n298 B.n297 585
R748 B.n492 B.n491 585
R749 B.n491 B.n490 585
R750 B.n493 B.n295 585
R751 B.n489 B.n295 585
R752 B.n495 B.n494 585
R753 B.n496 B.n495 585
R754 B.n290 B.n289 585
R755 B.n291 B.n290 585
R756 B.n504 B.n503 585
R757 B.n503 B.n502 585
R758 B.n505 B.n288 585
R759 B.n288 B.n287 585
R760 B.n507 B.n506 585
R761 B.n508 B.n507 585
R762 B.n282 B.n281 585
R763 B.n283 B.n282 585
R764 B.n516 B.n515 585
R765 B.n515 B.n514 585
R766 B.n517 B.n280 585
R767 B.n280 B.n279 585
R768 B.n519 B.n518 585
R769 B.n520 B.n519 585
R770 B.n274 B.n273 585
R771 B.n275 B.n274 585
R772 B.n528 B.n527 585
R773 B.n527 B.n526 585
R774 B.n529 B.n272 585
R775 B.n272 B.n271 585
R776 B.n531 B.n530 585
R777 B.n532 B.n531 585
R778 B.n266 B.n265 585
R779 B.n267 B.n266 585
R780 B.n540 B.n539 585
R781 B.n539 B.n538 585
R782 B.n541 B.n264 585
R783 B.n264 B.n263 585
R784 B.n543 B.n542 585
R785 B.n544 B.n543 585
R786 B.n258 B.n257 585
R787 B.n259 B.n258 585
R788 B.n552 B.n551 585
R789 B.n551 B.n550 585
R790 B.n553 B.n256 585
R791 B.n256 B.n255 585
R792 B.n555 B.n554 585
R793 B.n556 B.n555 585
R794 B.n250 B.n249 585
R795 B.n251 B.n250 585
R796 B.n564 B.n563 585
R797 B.n563 B.n562 585
R798 B.n565 B.n248 585
R799 B.n248 B.n247 585
R800 B.n567 B.n566 585
R801 B.n568 B.n567 585
R802 B.n242 B.n241 585
R803 B.n243 B.n242 585
R804 B.n576 B.n575 585
R805 B.n575 B.n574 585
R806 B.n577 B.n240 585
R807 B.n240 B.n239 585
R808 B.n579 B.n578 585
R809 B.n580 B.n579 585
R810 B.n234 B.n233 585
R811 B.n235 B.n234 585
R812 B.n589 B.n588 585
R813 B.n588 B.n587 585
R814 B.n590 B.n232 585
R815 B.n232 B.n231 585
R816 B.n592 B.n591 585
R817 B.n593 B.n592 585
R818 B.n2 B.n0 585
R819 B.n4 B.n2 585
R820 B.n3 B.n1 585
R821 B.n744 B.n3 585
R822 B.n742 B.n741 585
R823 B.n743 B.n742 585
R824 B.n740 B.n9 585
R825 B.n9 B.n8 585
R826 B.n739 B.n738 585
R827 B.n738 B.n737 585
R828 B.n11 B.n10 585
R829 B.n736 B.n11 585
R830 B.n734 B.n733 585
R831 B.n735 B.n734 585
R832 B.n732 B.n16 585
R833 B.n16 B.n15 585
R834 B.n731 B.n730 585
R835 B.n730 B.n729 585
R836 B.n18 B.n17 585
R837 B.n728 B.n18 585
R838 B.n726 B.n725 585
R839 B.n727 B.n726 585
R840 B.n724 B.n23 585
R841 B.n23 B.n22 585
R842 B.n723 B.n722 585
R843 B.n722 B.n721 585
R844 B.n25 B.n24 585
R845 B.n720 B.n25 585
R846 B.n718 B.n717 585
R847 B.n719 B.n718 585
R848 B.n716 B.n30 585
R849 B.n30 B.n29 585
R850 B.n715 B.n714 585
R851 B.n714 B.n713 585
R852 B.n32 B.n31 585
R853 B.n712 B.n32 585
R854 B.n710 B.n709 585
R855 B.n711 B.n710 585
R856 B.n708 B.n37 585
R857 B.n37 B.n36 585
R858 B.n707 B.n706 585
R859 B.n706 B.n705 585
R860 B.n39 B.n38 585
R861 B.n704 B.n39 585
R862 B.n702 B.n701 585
R863 B.n703 B.n702 585
R864 B.n700 B.n44 585
R865 B.n44 B.n43 585
R866 B.n699 B.n698 585
R867 B.n698 B.n697 585
R868 B.n46 B.n45 585
R869 B.n696 B.n46 585
R870 B.n694 B.n693 585
R871 B.n695 B.n694 585
R872 B.n692 B.n51 585
R873 B.n51 B.n50 585
R874 B.n691 B.n690 585
R875 B.n690 B.n689 585
R876 B.n53 B.n52 585
R877 B.n688 B.n53 585
R878 B.n686 B.n685 585
R879 B.n687 B.n686 585
R880 B.n684 B.n58 585
R881 B.n58 B.n57 585
R882 B.n683 B.n682 585
R883 B.n682 B.n681 585
R884 B.n60 B.n59 585
R885 B.n680 B.n60 585
R886 B.n678 B.n677 585
R887 B.n679 B.n678 585
R888 B.n676 B.n64 585
R889 B.n67 B.n64 585
R890 B.n675 B.n674 585
R891 B.n674 B.n673 585
R892 B.n66 B.n65 585
R893 B.n672 B.n66 585
R894 B.n670 B.n669 585
R895 B.n671 B.n670 585
R896 B.n668 B.n72 585
R897 B.n72 B.n71 585
R898 B.n667 B.n666 585
R899 B.n666 B.n665 585
R900 B.n74 B.n73 585
R901 B.n664 B.n74 585
R902 B.n662 B.n661 585
R903 B.n663 B.n662 585
R904 B.n660 B.n79 585
R905 B.n79 B.n78 585
R906 B.n659 B.n658 585
R907 B.n658 B.n657 585
R908 B.n747 B.n746 585
R909 B.n746 B.n745 585
R910 B.n466 B.n313 487.695
R911 B.n658 B.n81 487.695
R912 B.n464 B.n315 487.695
R913 B.n654 B.n82 487.695
R914 B.n411 B.t7 259.277
R915 B.n112 B.t16 259.277
R916 B.n333 B.t10 259.277
R917 B.n115 B.t13 259.277
R918 B.n656 B.n655 256.663
R919 B.n656 B.n110 256.663
R920 B.n656 B.n109 256.663
R921 B.n656 B.n108 256.663
R922 B.n656 B.n107 256.663
R923 B.n656 B.n106 256.663
R924 B.n656 B.n105 256.663
R925 B.n656 B.n104 256.663
R926 B.n656 B.n103 256.663
R927 B.n656 B.n102 256.663
R928 B.n656 B.n101 256.663
R929 B.n656 B.n100 256.663
R930 B.n656 B.n99 256.663
R931 B.n656 B.n98 256.663
R932 B.n656 B.n97 256.663
R933 B.n656 B.n96 256.663
R934 B.n656 B.n95 256.663
R935 B.n656 B.n94 256.663
R936 B.n656 B.n93 256.663
R937 B.n656 B.n92 256.663
R938 B.n656 B.n91 256.663
R939 B.n656 B.n90 256.663
R940 B.n656 B.n89 256.663
R941 B.n656 B.n88 256.663
R942 B.n656 B.n87 256.663
R943 B.n656 B.n86 256.663
R944 B.n656 B.n85 256.663
R945 B.n656 B.n84 256.663
R946 B.n656 B.n83 256.663
R947 B.n347 B.n314 256.663
R948 B.n350 B.n314 256.663
R949 B.n356 B.n314 256.663
R950 B.n358 B.n314 256.663
R951 B.n364 B.n314 256.663
R952 B.n366 B.n314 256.663
R953 B.n372 B.n314 256.663
R954 B.n374 B.n314 256.663
R955 B.n380 B.n314 256.663
R956 B.n382 B.n314 256.663
R957 B.n388 B.n314 256.663
R958 B.n390 B.n314 256.663
R959 B.n397 B.n314 256.663
R960 B.n399 B.n314 256.663
R961 B.n405 B.n314 256.663
R962 B.n407 B.n314 256.663
R963 B.n416 B.n314 256.663
R964 B.n418 B.n314 256.663
R965 B.n424 B.n314 256.663
R966 B.n426 B.n314 256.663
R967 B.n432 B.n314 256.663
R968 B.n434 B.n314 256.663
R969 B.n440 B.n314 256.663
R970 B.n442 B.n314 256.663
R971 B.n448 B.n314 256.663
R972 B.n450 B.n314 256.663
R973 B.n456 B.n314 256.663
R974 B.n459 B.n314 256.663
R975 B.n411 B.t4 248.572
R976 B.n333 B.t8 248.572
R977 B.n115 B.t11 248.572
R978 B.n112 B.t15 248.572
R979 B.n412 B.t6 180.538
R980 B.n113 B.t17 180.538
R981 B.n334 B.t9 180.538
R982 B.n116 B.t14 180.538
R983 B.n466 B.n311 163.367
R984 B.n470 B.n311 163.367
R985 B.n470 B.n305 163.367
R986 B.n478 B.n305 163.367
R987 B.n478 B.n303 163.367
R988 B.n482 B.n303 163.367
R989 B.n482 B.n297 163.367
R990 B.n491 B.n297 163.367
R991 B.n491 B.n295 163.367
R992 B.n495 B.n295 163.367
R993 B.n495 B.n290 163.367
R994 B.n503 B.n290 163.367
R995 B.n503 B.n288 163.367
R996 B.n507 B.n288 163.367
R997 B.n507 B.n282 163.367
R998 B.n515 B.n282 163.367
R999 B.n515 B.n280 163.367
R1000 B.n519 B.n280 163.367
R1001 B.n519 B.n274 163.367
R1002 B.n527 B.n274 163.367
R1003 B.n527 B.n272 163.367
R1004 B.n531 B.n272 163.367
R1005 B.n531 B.n266 163.367
R1006 B.n539 B.n266 163.367
R1007 B.n539 B.n264 163.367
R1008 B.n543 B.n264 163.367
R1009 B.n543 B.n258 163.367
R1010 B.n551 B.n258 163.367
R1011 B.n551 B.n256 163.367
R1012 B.n555 B.n256 163.367
R1013 B.n555 B.n250 163.367
R1014 B.n563 B.n250 163.367
R1015 B.n563 B.n248 163.367
R1016 B.n567 B.n248 163.367
R1017 B.n567 B.n242 163.367
R1018 B.n575 B.n242 163.367
R1019 B.n575 B.n240 163.367
R1020 B.n579 B.n240 163.367
R1021 B.n579 B.n234 163.367
R1022 B.n588 B.n234 163.367
R1023 B.n588 B.n232 163.367
R1024 B.n592 B.n232 163.367
R1025 B.n592 B.n2 163.367
R1026 B.n746 B.n2 163.367
R1027 B.n746 B.n3 163.367
R1028 B.n742 B.n3 163.367
R1029 B.n742 B.n9 163.367
R1030 B.n738 B.n9 163.367
R1031 B.n738 B.n11 163.367
R1032 B.n734 B.n11 163.367
R1033 B.n734 B.n16 163.367
R1034 B.n730 B.n16 163.367
R1035 B.n730 B.n18 163.367
R1036 B.n726 B.n18 163.367
R1037 B.n726 B.n23 163.367
R1038 B.n722 B.n23 163.367
R1039 B.n722 B.n25 163.367
R1040 B.n718 B.n25 163.367
R1041 B.n718 B.n30 163.367
R1042 B.n714 B.n30 163.367
R1043 B.n714 B.n32 163.367
R1044 B.n710 B.n32 163.367
R1045 B.n710 B.n37 163.367
R1046 B.n706 B.n37 163.367
R1047 B.n706 B.n39 163.367
R1048 B.n702 B.n39 163.367
R1049 B.n702 B.n44 163.367
R1050 B.n698 B.n44 163.367
R1051 B.n698 B.n46 163.367
R1052 B.n694 B.n46 163.367
R1053 B.n694 B.n51 163.367
R1054 B.n690 B.n51 163.367
R1055 B.n690 B.n53 163.367
R1056 B.n686 B.n53 163.367
R1057 B.n686 B.n58 163.367
R1058 B.n682 B.n58 163.367
R1059 B.n682 B.n60 163.367
R1060 B.n678 B.n60 163.367
R1061 B.n678 B.n64 163.367
R1062 B.n674 B.n64 163.367
R1063 B.n674 B.n66 163.367
R1064 B.n670 B.n66 163.367
R1065 B.n670 B.n72 163.367
R1066 B.n666 B.n72 163.367
R1067 B.n666 B.n74 163.367
R1068 B.n662 B.n74 163.367
R1069 B.n662 B.n79 163.367
R1070 B.n658 B.n79 163.367
R1071 B.n349 B.n348 163.367
R1072 B.n351 B.n349 163.367
R1073 B.n355 B.n344 163.367
R1074 B.n359 B.n357 163.367
R1075 B.n363 B.n342 163.367
R1076 B.n367 B.n365 163.367
R1077 B.n371 B.n340 163.367
R1078 B.n375 B.n373 163.367
R1079 B.n379 B.n338 163.367
R1080 B.n383 B.n381 163.367
R1081 B.n387 B.n336 163.367
R1082 B.n391 B.n389 163.367
R1083 B.n396 B.n332 163.367
R1084 B.n400 B.n398 163.367
R1085 B.n404 B.n330 163.367
R1086 B.n408 B.n406 163.367
R1087 B.n415 B.n328 163.367
R1088 B.n419 B.n417 163.367
R1089 B.n423 B.n326 163.367
R1090 B.n427 B.n425 163.367
R1091 B.n431 B.n324 163.367
R1092 B.n435 B.n433 163.367
R1093 B.n439 B.n322 163.367
R1094 B.n443 B.n441 163.367
R1095 B.n447 B.n320 163.367
R1096 B.n451 B.n449 163.367
R1097 B.n455 B.n318 163.367
R1098 B.n458 B.n457 163.367
R1099 B.n460 B.n315 163.367
R1100 B.n464 B.n309 163.367
R1101 B.n472 B.n309 163.367
R1102 B.n472 B.n307 163.367
R1103 B.n476 B.n307 163.367
R1104 B.n476 B.n301 163.367
R1105 B.n484 B.n301 163.367
R1106 B.n484 B.n299 163.367
R1107 B.n488 B.n299 163.367
R1108 B.n488 B.n294 163.367
R1109 B.n497 B.n294 163.367
R1110 B.n497 B.n292 163.367
R1111 B.n501 B.n292 163.367
R1112 B.n501 B.n286 163.367
R1113 B.n509 B.n286 163.367
R1114 B.n509 B.n284 163.367
R1115 B.n513 B.n284 163.367
R1116 B.n513 B.n278 163.367
R1117 B.n521 B.n278 163.367
R1118 B.n521 B.n276 163.367
R1119 B.n525 B.n276 163.367
R1120 B.n525 B.n270 163.367
R1121 B.n533 B.n270 163.367
R1122 B.n533 B.n268 163.367
R1123 B.n537 B.n268 163.367
R1124 B.n537 B.n262 163.367
R1125 B.n545 B.n262 163.367
R1126 B.n545 B.n260 163.367
R1127 B.n549 B.n260 163.367
R1128 B.n549 B.n254 163.367
R1129 B.n557 B.n254 163.367
R1130 B.n557 B.n252 163.367
R1131 B.n561 B.n252 163.367
R1132 B.n561 B.n246 163.367
R1133 B.n569 B.n246 163.367
R1134 B.n569 B.n244 163.367
R1135 B.n573 B.n244 163.367
R1136 B.n573 B.n238 163.367
R1137 B.n581 B.n238 163.367
R1138 B.n581 B.n236 163.367
R1139 B.n586 B.n236 163.367
R1140 B.n586 B.n230 163.367
R1141 B.n594 B.n230 163.367
R1142 B.n595 B.n594 163.367
R1143 B.n595 B.n5 163.367
R1144 B.n6 B.n5 163.367
R1145 B.n7 B.n6 163.367
R1146 B.n600 B.n7 163.367
R1147 B.n600 B.n12 163.367
R1148 B.n13 B.n12 163.367
R1149 B.n14 B.n13 163.367
R1150 B.n605 B.n14 163.367
R1151 B.n605 B.n19 163.367
R1152 B.n20 B.n19 163.367
R1153 B.n21 B.n20 163.367
R1154 B.n610 B.n21 163.367
R1155 B.n610 B.n26 163.367
R1156 B.n27 B.n26 163.367
R1157 B.n28 B.n27 163.367
R1158 B.n615 B.n28 163.367
R1159 B.n615 B.n33 163.367
R1160 B.n34 B.n33 163.367
R1161 B.n35 B.n34 163.367
R1162 B.n620 B.n35 163.367
R1163 B.n620 B.n40 163.367
R1164 B.n41 B.n40 163.367
R1165 B.n42 B.n41 163.367
R1166 B.n625 B.n42 163.367
R1167 B.n625 B.n47 163.367
R1168 B.n48 B.n47 163.367
R1169 B.n49 B.n48 163.367
R1170 B.n630 B.n49 163.367
R1171 B.n630 B.n54 163.367
R1172 B.n55 B.n54 163.367
R1173 B.n56 B.n55 163.367
R1174 B.n635 B.n56 163.367
R1175 B.n635 B.n61 163.367
R1176 B.n62 B.n61 163.367
R1177 B.n63 B.n62 163.367
R1178 B.n640 B.n63 163.367
R1179 B.n640 B.n68 163.367
R1180 B.n69 B.n68 163.367
R1181 B.n70 B.n69 163.367
R1182 B.n645 B.n70 163.367
R1183 B.n645 B.n75 163.367
R1184 B.n76 B.n75 163.367
R1185 B.n77 B.n76 163.367
R1186 B.n650 B.n77 163.367
R1187 B.n650 B.n82 163.367
R1188 B.n120 B.n119 163.367
R1189 B.n124 B.n123 163.367
R1190 B.n128 B.n127 163.367
R1191 B.n132 B.n131 163.367
R1192 B.n136 B.n135 163.367
R1193 B.n140 B.n139 163.367
R1194 B.n144 B.n143 163.367
R1195 B.n148 B.n147 163.367
R1196 B.n152 B.n151 163.367
R1197 B.n156 B.n155 163.367
R1198 B.n160 B.n159 163.367
R1199 B.n164 B.n163 163.367
R1200 B.n168 B.n167 163.367
R1201 B.n172 B.n171 163.367
R1202 B.n176 B.n175 163.367
R1203 B.n180 B.n179 163.367
R1204 B.n184 B.n183 163.367
R1205 B.n188 B.n187 163.367
R1206 B.n192 B.n191 163.367
R1207 B.n196 B.n195 163.367
R1208 B.n200 B.n199 163.367
R1209 B.n204 B.n203 163.367
R1210 B.n208 B.n207 163.367
R1211 B.n212 B.n211 163.367
R1212 B.n216 B.n215 163.367
R1213 B.n220 B.n219 163.367
R1214 B.n224 B.n223 163.367
R1215 B.n226 B.n111 163.367
R1216 B.n465 B.n314 115.281
R1217 B.n657 B.n656 115.281
R1218 B.n412 B.n411 78.7399
R1219 B.n334 B.n333 78.7399
R1220 B.n116 B.n115 78.7399
R1221 B.n113 B.n112 78.7399
R1222 B.n347 B.n313 71.676
R1223 B.n351 B.n350 71.676
R1224 B.n356 B.n355 71.676
R1225 B.n359 B.n358 71.676
R1226 B.n364 B.n363 71.676
R1227 B.n367 B.n366 71.676
R1228 B.n372 B.n371 71.676
R1229 B.n375 B.n374 71.676
R1230 B.n380 B.n379 71.676
R1231 B.n383 B.n382 71.676
R1232 B.n388 B.n387 71.676
R1233 B.n391 B.n390 71.676
R1234 B.n397 B.n396 71.676
R1235 B.n400 B.n399 71.676
R1236 B.n405 B.n404 71.676
R1237 B.n408 B.n407 71.676
R1238 B.n416 B.n415 71.676
R1239 B.n419 B.n418 71.676
R1240 B.n424 B.n423 71.676
R1241 B.n427 B.n426 71.676
R1242 B.n432 B.n431 71.676
R1243 B.n435 B.n434 71.676
R1244 B.n440 B.n439 71.676
R1245 B.n443 B.n442 71.676
R1246 B.n448 B.n447 71.676
R1247 B.n451 B.n450 71.676
R1248 B.n456 B.n455 71.676
R1249 B.n459 B.n458 71.676
R1250 B.n83 B.n81 71.676
R1251 B.n120 B.n84 71.676
R1252 B.n124 B.n85 71.676
R1253 B.n128 B.n86 71.676
R1254 B.n132 B.n87 71.676
R1255 B.n136 B.n88 71.676
R1256 B.n140 B.n89 71.676
R1257 B.n144 B.n90 71.676
R1258 B.n148 B.n91 71.676
R1259 B.n152 B.n92 71.676
R1260 B.n156 B.n93 71.676
R1261 B.n160 B.n94 71.676
R1262 B.n164 B.n95 71.676
R1263 B.n168 B.n96 71.676
R1264 B.n172 B.n97 71.676
R1265 B.n176 B.n98 71.676
R1266 B.n180 B.n99 71.676
R1267 B.n184 B.n100 71.676
R1268 B.n188 B.n101 71.676
R1269 B.n192 B.n102 71.676
R1270 B.n196 B.n103 71.676
R1271 B.n200 B.n104 71.676
R1272 B.n204 B.n105 71.676
R1273 B.n208 B.n106 71.676
R1274 B.n212 B.n107 71.676
R1275 B.n216 B.n108 71.676
R1276 B.n220 B.n109 71.676
R1277 B.n224 B.n110 71.676
R1278 B.n655 B.n111 71.676
R1279 B.n655 B.n654 71.676
R1280 B.n226 B.n110 71.676
R1281 B.n223 B.n109 71.676
R1282 B.n219 B.n108 71.676
R1283 B.n215 B.n107 71.676
R1284 B.n211 B.n106 71.676
R1285 B.n207 B.n105 71.676
R1286 B.n203 B.n104 71.676
R1287 B.n199 B.n103 71.676
R1288 B.n195 B.n102 71.676
R1289 B.n191 B.n101 71.676
R1290 B.n187 B.n100 71.676
R1291 B.n183 B.n99 71.676
R1292 B.n179 B.n98 71.676
R1293 B.n175 B.n97 71.676
R1294 B.n171 B.n96 71.676
R1295 B.n167 B.n95 71.676
R1296 B.n163 B.n94 71.676
R1297 B.n159 B.n93 71.676
R1298 B.n155 B.n92 71.676
R1299 B.n151 B.n91 71.676
R1300 B.n147 B.n90 71.676
R1301 B.n143 B.n89 71.676
R1302 B.n139 B.n88 71.676
R1303 B.n135 B.n87 71.676
R1304 B.n131 B.n86 71.676
R1305 B.n127 B.n85 71.676
R1306 B.n123 B.n84 71.676
R1307 B.n119 B.n83 71.676
R1308 B.n348 B.n347 71.676
R1309 B.n350 B.n344 71.676
R1310 B.n357 B.n356 71.676
R1311 B.n358 B.n342 71.676
R1312 B.n365 B.n364 71.676
R1313 B.n366 B.n340 71.676
R1314 B.n373 B.n372 71.676
R1315 B.n374 B.n338 71.676
R1316 B.n381 B.n380 71.676
R1317 B.n382 B.n336 71.676
R1318 B.n389 B.n388 71.676
R1319 B.n390 B.n332 71.676
R1320 B.n398 B.n397 71.676
R1321 B.n399 B.n330 71.676
R1322 B.n406 B.n405 71.676
R1323 B.n407 B.n328 71.676
R1324 B.n417 B.n416 71.676
R1325 B.n418 B.n326 71.676
R1326 B.n425 B.n424 71.676
R1327 B.n426 B.n324 71.676
R1328 B.n433 B.n432 71.676
R1329 B.n434 B.n322 71.676
R1330 B.n441 B.n440 71.676
R1331 B.n442 B.n320 71.676
R1332 B.n449 B.n448 71.676
R1333 B.n450 B.n318 71.676
R1334 B.n457 B.n456 71.676
R1335 B.n460 B.n459 71.676
R1336 B.n465 B.n310 65.8746
R1337 B.n471 B.n310 65.8746
R1338 B.n471 B.n306 65.8746
R1339 B.n477 B.n306 65.8746
R1340 B.n477 B.n302 65.8746
R1341 B.n483 B.n302 65.8746
R1342 B.n483 B.n298 65.8746
R1343 B.n490 B.n298 65.8746
R1344 B.n490 B.n489 65.8746
R1345 B.n496 B.n291 65.8746
R1346 B.n502 B.n291 65.8746
R1347 B.n502 B.n287 65.8746
R1348 B.n508 B.n287 65.8746
R1349 B.n508 B.n283 65.8746
R1350 B.n514 B.n283 65.8746
R1351 B.n514 B.n279 65.8746
R1352 B.n520 B.n279 65.8746
R1353 B.n520 B.n275 65.8746
R1354 B.n526 B.n275 65.8746
R1355 B.n526 B.n271 65.8746
R1356 B.n532 B.n271 65.8746
R1357 B.n532 B.n267 65.8746
R1358 B.n538 B.n267 65.8746
R1359 B.n544 B.n263 65.8746
R1360 B.n544 B.n259 65.8746
R1361 B.n550 B.n259 65.8746
R1362 B.n550 B.n255 65.8746
R1363 B.n556 B.n255 65.8746
R1364 B.n556 B.n251 65.8746
R1365 B.n562 B.n251 65.8746
R1366 B.n562 B.n247 65.8746
R1367 B.n568 B.n247 65.8746
R1368 B.n568 B.n243 65.8746
R1369 B.n574 B.n243 65.8746
R1370 B.n580 B.n239 65.8746
R1371 B.n580 B.n235 65.8746
R1372 B.n587 B.n235 65.8746
R1373 B.n587 B.n231 65.8746
R1374 B.n593 B.n231 65.8746
R1375 B.n593 B.n4 65.8746
R1376 B.n745 B.n4 65.8746
R1377 B.n745 B.n744 65.8746
R1378 B.n744 B.n743 65.8746
R1379 B.n743 B.n8 65.8746
R1380 B.n737 B.n8 65.8746
R1381 B.n737 B.n736 65.8746
R1382 B.n736 B.n735 65.8746
R1383 B.n735 B.n15 65.8746
R1384 B.n729 B.n728 65.8746
R1385 B.n728 B.n727 65.8746
R1386 B.n727 B.n22 65.8746
R1387 B.n721 B.n22 65.8746
R1388 B.n721 B.n720 65.8746
R1389 B.n720 B.n719 65.8746
R1390 B.n719 B.n29 65.8746
R1391 B.n713 B.n29 65.8746
R1392 B.n713 B.n712 65.8746
R1393 B.n712 B.n711 65.8746
R1394 B.n711 B.n36 65.8746
R1395 B.n705 B.n704 65.8746
R1396 B.n704 B.n703 65.8746
R1397 B.n703 B.n43 65.8746
R1398 B.n697 B.n43 65.8746
R1399 B.n697 B.n696 65.8746
R1400 B.n696 B.n695 65.8746
R1401 B.n695 B.n50 65.8746
R1402 B.n689 B.n50 65.8746
R1403 B.n689 B.n688 65.8746
R1404 B.n688 B.n687 65.8746
R1405 B.n687 B.n57 65.8746
R1406 B.n681 B.n57 65.8746
R1407 B.n681 B.n680 65.8746
R1408 B.n680 B.n679 65.8746
R1409 B.n673 B.n67 65.8746
R1410 B.n673 B.n672 65.8746
R1411 B.n672 B.n671 65.8746
R1412 B.n671 B.n71 65.8746
R1413 B.n665 B.n71 65.8746
R1414 B.n665 B.n664 65.8746
R1415 B.n664 B.n663 65.8746
R1416 B.n663 B.n78 65.8746
R1417 B.n657 B.n78 65.8746
R1418 B.n413 B.n412 59.5399
R1419 B.n393 B.n334 59.5399
R1420 B.n117 B.n116 59.5399
R1421 B.n114 B.n113 59.5399
R1422 B.n496 B.t5 43.5936
R1423 B.n679 B.t12 43.5936
R1424 B.t1 B.n239 37.7812
R1425 B.t0 B.n15 37.7812
R1426 B.t2 B.n263 33.9063
R1427 B.t3 B.n36 33.9063
R1428 B.n538 B.t2 31.9688
R1429 B.n705 B.t3 31.9688
R1430 B.n659 B.n80 31.6883
R1431 B.n653 B.n652 31.6883
R1432 B.n463 B.n462 31.6883
R1433 B.n467 B.n312 31.6883
R1434 B.n574 B.t1 28.0939
R1435 B.n729 B.t0 28.0939
R1436 B.n489 B.t5 22.2814
R1437 B.n67 B.t12 22.2814
R1438 B B.n747 18.0485
R1439 B.n118 B.n80 10.6151
R1440 B.n121 B.n118 10.6151
R1441 B.n122 B.n121 10.6151
R1442 B.n125 B.n122 10.6151
R1443 B.n126 B.n125 10.6151
R1444 B.n129 B.n126 10.6151
R1445 B.n130 B.n129 10.6151
R1446 B.n133 B.n130 10.6151
R1447 B.n134 B.n133 10.6151
R1448 B.n137 B.n134 10.6151
R1449 B.n138 B.n137 10.6151
R1450 B.n141 B.n138 10.6151
R1451 B.n142 B.n141 10.6151
R1452 B.n145 B.n142 10.6151
R1453 B.n146 B.n145 10.6151
R1454 B.n149 B.n146 10.6151
R1455 B.n150 B.n149 10.6151
R1456 B.n153 B.n150 10.6151
R1457 B.n154 B.n153 10.6151
R1458 B.n157 B.n154 10.6151
R1459 B.n158 B.n157 10.6151
R1460 B.n161 B.n158 10.6151
R1461 B.n162 B.n161 10.6151
R1462 B.n166 B.n165 10.6151
R1463 B.n169 B.n166 10.6151
R1464 B.n170 B.n169 10.6151
R1465 B.n173 B.n170 10.6151
R1466 B.n174 B.n173 10.6151
R1467 B.n177 B.n174 10.6151
R1468 B.n178 B.n177 10.6151
R1469 B.n181 B.n178 10.6151
R1470 B.n182 B.n181 10.6151
R1471 B.n186 B.n185 10.6151
R1472 B.n189 B.n186 10.6151
R1473 B.n190 B.n189 10.6151
R1474 B.n193 B.n190 10.6151
R1475 B.n194 B.n193 10.6151
R1476 B.n197 B.n194 10.6151
R1477 B.n198 B.n197 10.6151
R1478 B.n201 B.n198 10.6151
R1479 B.n202 B.n201 10.6151
R1480 B.n205 B.n202 10.6151
R1481 B.n206 B.n205 10.6151
R1482 B.n209 B.n206 10.6151
R1483 B.n210 B.n209 10.6151
R1484 B.n213 B.n210 10.6151
R1485 B.n214 B.n213 10.6151
R1486 B.n217 B.n214 10.6151
R1487 B.n218 B.n217 10.6151
R1488 B.n221 B.n218 10.6151
R1489 B.n222 B.n221 10.6151
R1490 B.n225 B.n222 10.6151
R1491 B.n227 B.n225 10.6151
R1492 B.n228 B.n227 10.6151
R1493 B.n653 B.n228 10.6151
R1494 B.n463 B.n308 10.6151
R1495 B.n473 B.n308 10.6151
R1496 B.n474 B.n473 10.6151
R1497 B.n475 B.n474 10.6151
R1498 B.n475 B.n300 10.6151
R1499 B.n485 B.n300 10.6151
R1500 B.n486 B.n485 10.6151
R1501 B.n487 B.n486 10.6151
R1502 B.n487 B.n293 10.6151
R1503 B.n498 B.n293 10.6151
R1504 B.n499 B.n498 10.6151
R1505 B.n500 B.n499 10.6151
R1506 B.n500 B.n285 10.6151
R1507 B.n510 B.n285 10.6151
R1508 B.n511 B.n510 10.6151
R1509 B.n512 B.n511 10.6151
R1510 B.n512 B.n277 10.6151
R1511 B.n522 B.n277 10.6151
R1512 B.n523 B.n522 10.6151
R1513 B.n524 B.n523 10.6151
R1514 B.n524 B.n269 10.6151
R1515 B.n534 B.n269 10.6151
R1516 B.n535 B.n534 10.6151
R1517 B.n536 B.n535 10.6151
R1518 B.n536 B.n261 10.6151
R1519 B.n546 B.n261 10.6151
R1520 B.n547 B.n546 10.6151
R1521 B.n548 B.n547 10.6151
R1522 B.n548 B.n253 10.6151
R1523 B.n558 B.n253 10.6151
R1524 B.n559 B.n558 10.6151
R1525 B.n560 B.n559 10.6151
R1526 B.n560 B.n245 10.6151
R1527 B.n570 B.n245 10.6151
R1528 B.n571 B.n570 10.6151
R1529 B.n572 B.n571 10.6151
R1530 B.n572 B.n237 10.6151
R1531 B.n582 B.n237 10.6151
R1532 B.n583 B.n582 10.6151
R1533 B.n585 B.n583 10.6151
R1534 B.n585 B.n584 10.6151
R1535 B.n584 B.n229 10.6151
R1536 B.n596 B.n229 10.6151
R1537 B.n597 B.n596 10.6151
R1538 B.n598 B.n597 10.6151
R1539 B.n599 B.n598 10.6151
R1540 B.n601 B.n599 10.6151
R1541 B.n602 B.n601 10.6151
R1542 B.n603 B.n602 10.6151
R1543 B.n604 B.n603 10.6151
R1544 B.n606 B.n604 10.6151
R1545 B.n607 B.n606 10.6151
R1546 B.n608 B.n607 10.6151
R1547 B.n609 B.n608 10.6151
R1548 B.n611 B.n609 10.6151
R1549 B.n612 B.n611 10.6151
R1550 B.n613 B.n612 10.6151
R1551 B.n614 B.n613 10.6151
R1552 B.n616 B.n614 10.6151
R1553 B.n617 B.n616 10.6151
R1554 B.n618 B.n617 10.6151
R1555 B.n619 B.n618 10.6151
R1556 B.n621 B.n619 10.6151
R1557 B.n622 B.n621 10.6151
R1558 B.n623 B.n622 10.6151
R1559 B.n624 B.n623 10.6151
R1560 B.n626 B.n624 10.6151
R1561 B.n627 B.n626 10.6151
R1562 B.n628 B.n627 10.6151
R1563 B.n629 B.n628 10.6151
R1564 B.n631 B.n629 10.6151
R1565 B.n632 B.n631 10.6151
R1566 B.n633 B.n632 10.6151
R1567 B.n634 B.n633 10.6151
R1568 B.n636 B.n634 10.6151
R1569 B.n637 B.n636 10.6151
R1570 B.n638 B.n637 10.6151
R1571 B.n639 B.n638 10.6151
R1572 B.n641 B.n639 10.6151
R1573 B.n642 B.n641 10.6151
R1574 B.n643 B.n642 10.6151
R1575 B.n644 B.n643 10.6151
R1576 B.n646 B.n644 10.6151
R1577 B.n647 B.n646 10.6151
R1578 B.n648 B.n647 10.6151
R1579 B.n649 B.n648 10.6151
R1580 B.n651 B.n649 10.6151
R1581 B.n652 B.n651 10.6151
R1582 B.n346 B.n312 10.6151
R1583 B.n346 B.n345 10.6151
R1584 B.n352 B.n345 10.6151
R1585 B.n353 B.n352 10.6151
R1586 B.n354 B.n353 10.6151
R1587 B.n354 B.n343 10.6151
R1588 B.n360 B.n343 10.6151
R1589 B.n361 B.n360 10.6151
R1590 B.n362 B.n361 10.6151
R1591 B.n362 B.n341 10.6151
R1592 B.n368 B.n341 10.6151
R1593 B.n369 B.n368 10.6151
R1594 B.n370 B.n369 10.6151
R1595 B.n370 B.n339 10.6151
R1596 B.n376 B.n339 10.6151
R1597 B.n377 B.n376 10.6151
R1598 B.n378 B.n377 10.6151
R1599 B.n378 B.n337 10.6151
R1600 B.n384 B.n337 10.6151
R1601 B.n385 B.n384 10.6151
R1602 B.n386 B.n385 10.6151
R1603 B.n386 B.n335 10.6151
R1604 B.n392 B.n335 10.6151
R1605 B.n395 B.n394 10.6151
R1606 B.n395 B.n331 10.6151
R1607 B.n401 B.n331 10.6151
R1608 B.n402 B.n401 10.6151
R1609 B.n403 B.n402 10.6151
R1610 B.n403 B.n329 10.6151
R1611 B.n409 B.n329 10.6151
R1612 B.n410 B.n409 10.6151
R1613 B.n414 B.n410 10.6151
R1614 B.n420 B.n327 10.6151
R1615 B.n421 B.n420 10.6151
R1616 B.n422 B.n421 10.6151
R1617 B.n422 B.n325 10.6151
R1618 B.n428 B.n325 10.6151
R1619 B.n429 B.n428 10.6151
R1620 B.n430 B.n429 10.6151
R1621 B.n430 B.n323 10.6151
R1622 B.n436 B.n323 10.6151
R1623 B.n437 B.n436 10.6151
R1624 B.n438 B.n437 10.6151
R1625 B.n438 B.n321 10.6151
R1626 B.n444 B.n321 10.6151
R1627 B.n445 B.n444 10.6151
R1628 B.n446 B.n445 10.6151
R1629 B.n446 B.n319 10.6151
R1630 B.n452 B.n319 10.6151
R1631 B.n453 B.n452 10.6151
R1632 B.n454 B.n453 10.6151
R1633 B.n454 B.n317 10.6151
R1634 B.n317 B.n316 10.6151
R1635 B.n461 B.n316 10.6151
R1636 B.n462 B.n461 10.6151
R1637 B.n468 B.n467 10.6151
R1638 B.n469 B.n468 10.6151
R1639 B.n469 B.n304 10.6151
R1640 B.n479 B.n304 10.6151
R1641 B.n480 B.n479 10.6151
R1642 B.n481 B.n480 10.6151
R1643 B.n481 B.n296 10.6151
R1644 B.n492 B.n296 10.6151
R1645 B.n493 B.n492 10.6151
R1646 B.n494 B.n493 10.6151
R1647 B.n494 B.n289 10.6151
R1648 B.n504 B.n289 10.6151
R1649 B.n505 B.n504 10.6151
R1650 B.n506 B.n505 10.6151
R1651 B.n506 B.n281 10.6151
R1652 B.n516 B.n281 10.6151
R1653 B.n517 B.n516 10.6151
R1654 B.n518 B.n517 10.6151
R1655 B.n518 B.n273 10.6151
R1656 B.n528 B.n273 10.6151
R1657 B.n529 B.n528 10.6151
R1658 B.n530 B.n529 10.6151
R1659 B.n530 B.n265 10.6151
R1660 B.n540 B.n265 10.6151
R1661 B.n541 B.n540 10.6151
R1662 B.n542 B.n541 10.6151
R1663 B.n542 B.n257 10.6151
R1664 B.n552 B.n257 10.6151
R1665 B.n553 B.n552 10.6151
R1666 B.n554 B.n553 10.6151
R1667 B.n554 B.n249 10.6151
R1668 B.n564 B.n249 10.6151
R1669 B.n565 B.n564 10.6151
R1670 B.n566 B.n565 10.6151
R1671 B.n566 B.n241 10.6151
R1672 B.n576 B.n241 10.6151
R1673 B.n577 B.n576 10.6151
R1674 B.n578 B.n577 10.6151
R1675 B.n578 B.n233 10.6151
R1676 B.n589 B.n233 10.6151
R1677 B.n590 B.n589 10.6151
R1678 B.n591 B.n590 10.6151
R1679 B.n591 B.n0 10.6151
R1680 B.n741 B.n1 10.6151
R1681 B.n741 B.n740 10.6151
R1682 B.n740 B.n739 10.6151
R1683 B.n739 B.n10 10.6151
R1684 B.n733 B.n10 10.6151
R1685 B.n733 B.n732 10.6151
R1686 B.n732 B.n731 10.6151
R1687 B.n731 B.n17 10.6151
R1688 B.n725 B.n17 10.6151
R1689 B.n725 B.n724 10.6151
R1690 B.n724 B.n723 10.6151
R1691 B.n723 B.n24 10.6151
R1692 B.n717 B.n24 10.6151
R1693 B.n717 B.n716 10.6151
R1694 B.n716 B.n715 10.6151
R1695 B.n715 B.n31 10.6151
R1696 B.n709 B.n31 10.6151
R1697 B.n709 B.n708 10.6151
R1698 B.n708 B.n707 10.6151
R1699 B.n707 B.n38 10.6151
R1700 B.n701 B.n38 10.6151
R1701 B.n701 B.n700 10.6151
R1702 B.n700 B.n699 10.6151
R1703 B.n699 B.n45 10.6151
R1704 B.n693 B.n45 10.6151
R1705 B.n693 B.n692 10.6151
R1706 B.n692 B.n691 10.6151
R1707 B.n691 B.n52 10.6151
R1708 B.n685 B.n52 10.6151
R1709 B.n685 B.n684 10.6151
R1710 B.n684 B.n683 10.6151
R1711 B.n683 B.n59 10.6151
R1712 B.n677 B.n59 10.6151
R1713 B.n677 B.n676 10.6151
R1714 B.n676 B.n675 10.6151
R1715 B.n675 B.n65 10.6151
R1716 B.n669 B.n65 10.6151
R1717 B.n669 B.n668 10.6151
R1718 B.n668 B.n667 10.6151
R1719 B.n667 B.n73 10.6151
R1720 B.n661 B.n73 10.6151
R1721 B.n661 B.n660 10.6151
R1722 B.n660 B.n659 10.6151
R1723 B.n162 B.n117 9.36635
R1724 B.n185 B.n114 9.36635
R1725 B.n393 B.n392 9.36635
R1726 B.n413 B.n327 9.36635
R1727 B.n747 B.n0 2.81026
R1728 B.n747 B.n1 2.81026
R1729 B.n165 B.n117 1.24928
R1730 B.n182 B.n114 1.24928
R1731 B.n394 B.n393 1.24928
R1732 B.n414 B.n413 1.24928
R1733 VN.n1 VN.t3 72.8411
R1734 VN.n0 VN.t0 72.8411
R1735 VN.n0 VN.t2 71.5072
R1736 VN.n1 VN.t1 71.5072
R1737 VN VN.n1 47.3638
R1738 VN VN.n0 1.90546
R1739 VDD2.n2 VDD2.n0 108.198
R1740 VDD2.n2 VDD2.n1 68.7422
R1741 VDD2.n1 VDD2.t2 3.25708
R1742 VDD2.n1 VDD2.t0 3.25708
R1743 VDD2.n0 VDD2.t3 3.25708
R1744 VDD2.n0 VDD2.t1 3.25708
R1745 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 4.48271f
C1 VDD2 VTAIL 4.54449f
C2 VP VN 5.90688f
C3 VP VDD1 3.0289f
C4 VDD2 VP 0.466397f
C5 VDD1 VN 0.150209f
C6 VDD2 VN 2.71374f
C7 VTAIL VP 3.23633f
C8 VDD2 VDD1 1.29942f
C9 VTAIL VN 3.22222f
C10 VDD2 B 3.949463f
C11 VDD1 B 8.024429f
C12 VTAIL B 6.766511f
C13 VN B 12.37859f
C14 VP B 10.774909f
C15 VDD2.t3 B 0.13536f
C16 VDD2.t1 B 0.13536f
C17 VDD2.n0 B 1.64812f
C18 VDD2.t2 B 0.13536f
C19 VDD2.t0 B 0.13536f
C20 VDD2.n1 B 1.13127f
C21 VDD2.n2 B 3.55537f
C22 VN.t2 B 1.71784f
C23 VN.t0 B 1.73046f
C24 VN.n0 B 1.02817f
C25 VN.t1 B 1.71784f
C26 VN.t3 B 1.73046f
C27 VN.n1 B 2.38555f
C28 VDD1.t1 B 0.138991f
C29 VDD1.t3 B 0.138991f
C30 VDD1.n0 B 1.16211f
C31 VDD1.t0 B 0.138991f
C32 VDD1.t2 B 0.138991f
C33 VDD1.n1 B 1.71798f
C34 VTAIL.n0 B 0.030239f
C35 VTAIL.n1 B 0.020718f
C36 VTAIL.n2 B 0.011133f
C37 VTAIL.n3 B 0.026314f
C38 VTAIL.n4 B 0.011788f
C39 VTAIL.n5 B 0.020718f
C40 VTAIL.n6 B 0.011133f
C41 VTAIL.n7 B 0.026314f
C42 VTAIL.n8 B 0.011788f
C43 VTAIL.n9 B 0.089117f
C44 VTAIL.t0 B 0.042915f
C45 VTAIL.n10 B 0.019736f
C46 VTAIL.n11 B 0.015543f
C47 VTAIL.n12 B 0.011133f
C48 VTAIL.n13 B 0.50049f
C49 VTAIL.n14 B 0.020718f
C50 VTAIL.n15 B 0.011133f
C51 VTAIL.n16 B 0.011788f
C52 VTAIL.n17 B 0.026314f
C53 VTAIL.n18 B 0.026314f
C54 VTAIL.n19 B 0.011788f
C55 VTAIL.n20 B 0.011133f
C56 VTAIL.n21 B 0.020718f
C57 VTAIL.n22 B 0.020718f
C58 VTAIL.n23 B 0.011133f
C59 VTAIL.n24 B 0.011788f
C60 VTAIL.n25 B 0.026314f
C61 VTAIL.n26 B 0.058943f
C62 VTAIL.n27 B 0.011788f
C63 VTAIL.n28 B 0.011133f
C64 VTAIL.n29 B 0.050152f
C65 VTAIL.n30 B 0.033252f
C66 VTAIL.n31 B 0.171048f
C67 VTAIL.n32 B 0.030239f
C68 VTAIL.n33 B 0.020718f
C69 VTAIL.n34 B 0.011133f
C70 VTAIL.n35 B 0.026314f
C71 VTAIL.n36 B 0.011788f
C72 VTAIL.n37 B 0.020718f
C73 VTAIL.n38 B 0.011133f
C74 VTAIL.n39 B 0.026314f
C75 VTAIL.n40 B 0.011788f
C76 VTAIL.n41 B 0.089117f
C77 VTAIL.t3 B 0.042915f
C78 VTAIL.n42 B 0.019736f
C79 VTAIL.n43 B 0.015543f
C80 VTAIL.n44 B 0.011133f
C81 VTAIL.n45 B 0.50049f
C82 VTAIL.n46 B 0.020718f
C83 VTAIL.n47 B 0.011133f
C84 VTAIL.n48 B 0.011788f
C85 VTAIL.n49 B 0.026314f
C86 VTAIL.n50 B 0.026314f
C87 VTAIL.n51 B 0.011788f
C88 VTAIL.n52 B 0.011133f
C89 VTAIL.n53 B 0.020718f
C90 VTAIL.n54 B 0.020718f
C91 VTAIL.n55 B 0.011133f
C92 VTAIL.n56 B 0.011788f
C93 VTAIL.n57 B 0.026314f
C94 VTAIL.n58 B 0.058943f
C95 VTAIL.n59 B 0.011788f
C96 VTAIL.n60 B 0.011133f
C97 VTAIL.n61 B 0.050152f
C98 VTAIL.n62 B 0.033252f
C99 VTAIL.n63 B 0.283989f
C100 VTAIL.n64 B 0.030239f
C101 VTAIL.n65 B 0.020718f
C102 VTAIL.n66 B 0.011133f
C103 VTAIL.n67 B 0.026314f
C104 VTAIL.n68 B 0.011788f
C105 VTAIL.n69 B 0.020718f
C106 VTAIL.n70 B 0.011133f
C107 VTAIL.n71 B 0.026314f
C108 VTAIL.n72 B 0.011788f
C109 VTAIL.n73 B 0.089117f
C110 VTAIL.t5 B 0.042915f
C111 VTAIL.n74 B 0.019736f
C112 VTAIL.n75 B 0.015543f
C113 VTAIL.n76 B 0.011133f
C114 VTAIL.n77 B 0.50049f
C115 VTAIL.n78 B 0.020718f
C116 VTAIL.n79 B 0.011133f
C117 VTAIL.n80 B 0.011788f
C118 VTAIL.n81 B 0.026314f
C119 VTAIL.n82 B 0.026314f
C120 VTAIL.n83 B 0.011788f
C121 VTAIL.n84 B 0.011133f
C122 VTAIL.n85 B 0.020718f
C123 VTAIL.n86 B 0.020718f
C124 VTAIL.n87 B 0.011133f
C125 VTAIL.n88 B 0.011788f
C126 VTAIL.n89 B 0.026314f
C127 VTAIL.n90 B 0.058943f
C128 VTAIL.n91 B 0.011788f
C129 VTAIL.n92 B 0.011133f
C130 VTAIL.n93 B 0.050152f
C131 VTAIL.n94 B 0.033252f
C132 VTAIL.n95 B 1.1176f
C133 VTAIL.n96 B 0.030239f
C134 VTAIL.n97 B 0.020718f
C135 VTAIL.n98 B 0.011133f
C136 VTAIL.n99 B 0.026314f
C137 VTAIL.n100 B 0.011788f
C138 VTAIL.n101 B 0.020718f
C139 VTAIL.n102 B 0.011133f
C140 VTAIL.n103 B 0.026314f
C141 VTAIL.n104 B 0.011788f
C142 VTAIL.n105 B 0.089117f
C143 VTAIL.t2 B 0.042915f
C144 VTAIL.n106 B 0.019736f
C145 VTAIL.n107 B 0.015543f
C146 VTAIL.n108 B 0.011133f
C147 VTAIL.n109 B 0.500491f
C148 VTAIL.n110 B 0.020718f
C149 VTAIL.n111 B 0.011133f
C150 VTAIL.n112 B 0.011788f
C151 VTAIL.n113 B 0.026314f
C152 VTAIL.n114 B 0.026314f
C153 VTAIL.n115 B 0.011788f
C154 VTAIL.n116 B 0.011133f
C155 VTAIL.n117 B 0.020718f
C156 VTAIL.n118 B 0.020718f
C157 VTAIL.n119 B 0.011133f
C158 VTAIL.n120 B 0.011788f
C159 VTAIL.n121 B 0.026314f
C160 VTAIL.n122 B 0.058943f
C161 VTAIL.n123 B 0.011788f
C162 VTAIL.n124 B 0.011133f
C163 VTAIL.n125 B 0.050152f
C164 VTAIL.n126 B 0.033252f
C165 VTAIL.n127 B 1.1176f
C166 VTAIL.n128 B 0.030239f
C167 VTAIL.n129 B 0.020718f
C168 VTAIL.n130 B 0.011133f
C169 VTAIL.n131 B 0.026314f
C170 VTAIL.n132 B 0.011788f
C171 VTAIL.n133 B 0.020718f
C172 VTAIL.n134 B 0.011133f
C173 VTAIL.n135 B 0.026314f
C174 VTAIL.n136 B 0.011788f
C175 VTAIL.n137 B 0.089117f
C176 VTAIL.t1 B 0.042915f
C177 VTAIL.n138 B 0.019736f
C178 VTAIL.n139 B 0.015543f
C179 VTAIL.n140 B 0.011133f
C180 VTAIL.n141 B 0.500491f
C181 VTAIL.n142 B 0.020718f
C182 VTAIL.n143 B 0.011133f
C183 VTAIL.n144 B 0.011788f
C184 VTAIL.n145 B 0.026314f
C185 VTAIL.n146 B 0.026314f
C186 VTAIL.n147 B 0.011788f
C187 VTAIL.n148 B 0.011133f
C188 VTAIL.n149 B 0.020718f
C189 VTAIL.n150 B 0.020718f
C190 VTAIL.n151 B 0.011133f
C191 VTAIL.n152 B 0.011788f
C192 VTAIL.n153 B 0.026314f
C193 VTAIL.n154 B 0.058943f
C194 VTAIL.n155 B 0.011788f
C195 VTAIL.n156 B 0.011133f
C196 VTAIL.n157 B 0.050152f
C197 VTAIL.n158 B 0.033252f
C198 VTAIL.n159 B 0.283989f
C199 VTAIL.n160 B 0.030239f
C200 VTAIL.n161 B 0.020718f
C201 VTAIL.n162 B 0.011133f
C202 VTAIL.n163 B 0.026314f
C203 VTAIL.n164 B 0.011788f
C204 VTAIL.n165 B 0.020718f
C205 VTAIL.n166 B 0.011133f
C206 VTAIL.n167 B 0.026314f
C207 VTAIL.n168 B 0.011788f
C208 VTAIL.n169 B 0.089117f
C209 VTAIL.t6 B 0.042915f
C210 VTAIL.n170 B 0.019736f
C211 VTAIL.n171 B 0.015543f
C212 VTAIL.n172 B 0.011133f
C213 VTAIL.n173 B 0.500491f
C214 VTAIL.n174 B 0.020718f
C215 VTAIL.n175 B 0.011133f
C216 VTAIL.n176 B 0.011788f
C217 VTAIL.n177 B 0.026314f
C218 VTAIL.n178 B 0.026314f
C219 VTAIL.n179 B 0.011788f
C220 VTAIL.n180 B 0.011133f
C221 VTAIL.n181 B 0.020718f
C222 VTAIL.n182 B 0.020718f
C223 VTAIL.n183 B 0.011133f
C224 VTAIL.n184 B 0.011788f
C225 VTAIL.n185 B 0.026314f
C226 VTAIL.n186 B 0.058943f
C227 VTAIL.n187 B 0.011788f
C228 VTAIL.n188 B 0.011133f
C229 VTAIL.n189 B 0.050152f
C230 VTAIL.n190 B 0.033252f
C231 VTAIL.n191 B 0.283989f
C232 VTAIL.n192 B 0.030239f
C233 VTAIL.n193 B 0.020718f
C234 VTAIL.n194 B 0.011133f
C235 VTAIL.n195 B 0.026314f
C236 VTAIL.n196 B 0.011788f
C237 VTAIL.n197 B 0.020718f
C238 VTAIL.n198 B 0.011133f
C239 VTAIL.n199 B 0.026314f
C240 VTAIL.n200 B 0.011788f
C241 VTAIL.n201 B 0.089117f
C242 VTAIL.t4 B 0.042915f
C243 VTAIL.n202 B 0.019736f
C244 VTAIL.n203 B 0.015543f
C245 VTAIL.n204 B 0.011133f
C246 VTAIL.n205 B 0.500491f
C247 VTAIL.n206 B 0.020718f
C248 VTAIL.n207 B 0.011133f
C249 VTAIL.n208 B 0.011788f
C250 VTAIL.n209 B 0.026314f
C251 VTAIL.n210 B 0.026314f
C252 VTAIL.n211 B 0.011788f
C253 VTAIL.n212 B 0.011133f
C254 VTAIL.n213 B 0.020718f
C255 VTAIL.n214 B 0.020718f
C256 VTAIL.n215 B 0.011133f
C257 VTAIL.n216 B 0.011788f
C258 VTAIL.n217 B 0.026314f
C259 VTAIL.n218 B 0.058943f
C260 VTAIL.n219 B 0.011788f
C261 VTAIL.n220 B 0.011133f
C262 VTAIL.n221 B 0.050152f
C263 VTAIL.n222 B 0.033252f
C264 VTAIL.n223 B 1.1176f
C265 VTAIL.n224 B 0.030239f
C266 VTAIL.n225 B 0.020718f
C267 VTAIL.n226 B 0.011133f
C268 VTAIL.n227 B 0.026314f
C269 VTAIL.n228 B 0.011788f
C270 VTAIL.n229 B 0.020718f
C271 VTAIL.n230 B 0.011133f
C272 VTAIL.n231 B 0.026314f
C273 VTAIL.n232 B 0.011788f
C274 VTAIL.n233 B 0.089117f
C275 VTAIL.t7 B 0.042915f
C276 VTAIL.n234 B 0.019736f
C277 VTAIL.n235 B 0.015543f
C278 VTAIL.n236 B 0.011133f
C279 VTAIL.n237 B 0.50049f
C280 VTAIL.n238 B 0.020718f
C281 VTAIL.n239 B 0.011133f
C282 VTAIL.n240 B 0.011788f
C283 VTAIL.n241 B 0.026314f
C284 VTAIL.n242 B 0.026314f
C285 VTAIL.n243 B 0.011788f
C286 VTAIL.n244 B 0.011133f
C287 VTAIL.n245 B 0.020718f
C288 VTAIL.n246 B 0.020718f
C289 VTAIL.n247 B 0.011133f
C290 VTAIL.n248 B 0.011788f
C291 VTAIL.n249 B 0.026314f
C292 VTAIL.n250 B 0.058943f
C293 VTAIL.n251 B 0.011788f
C294 VTAIL.n252 B 0.011133f
C295 VTAIL.n253 B 0.050152f
C296 VTAIL.n254 B 0.033252f
C297 VTAIL.n255 B 0.996893f
C298 VP.t1 B 1.44467f
C299 VP.n0 B 0.617835f
C300 VP.n1 B 0.024049f
C301 VP.n2 B 0.047546f
C302 VP.n3 B 0.024049f
C303 VP.n4 B 0.044597f
C304 VP.t2 B 1.77941f
C305 VP.t0 B 1.76644f
C306 VP.n5 B 2.44303f
C307 VP.n6 B 1.27884f
C308 VP.t3 B 1.44467f
C309 VP.n7 B 0.617835f
C310 VP.n8 B 0.023902f
C311 VP.n9 B 0.038809f
C312 VP.n10 B 0.024049f
C313 VP.n11 B 0.024049f
C314 VP.n12 B 0.044597f
C315 VP.n13 B 0.047546f
C316 VP.n14 B 0.019424f
C317 VP.n15 B 0.024049f
C318 VP.n16 B 0.024049f
C319 VP.n17 B 0.024049f
C320 VP.n18 B 0.044597f
C321 VP.n19 B 0.044597f
C322 VP.n20 B 0.023902f
C323 VP.n21 B 0.038809f
C324 VP.n22 B 0.07379f
.ends

