* NGSPICE file created from diff_pair_sample_1564.ext - technology: sky130A

.subckt diff_pair_sample_1564 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=0 ps=0 w=4.18 l=1.3
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=0 ps=0 w=4.18 l=1.3
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=1.6302 ps=9.14 w=4.18 l=1.3
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=1.6302 ps=9.14 w=4.18 l=1.3
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=0 ps=0 w=4.18 l=1.3
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=0 ps=0 w=4.18 l=1.3
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=1.6302 ps=9.14 w=4.18 l=1.3
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6302 pd=9.14 as=1.6302 ps=9.14 w=4.18 l=1.3
R0 B.n388 B.n387 585
R1 B.n389 B.n388 585
R2 B.n155 B.n58 585
R3 B.n154 B.n153 585
R4 B.n152 B.n151 585
R5 B.n150 B.n149 585
R6 B.n148 B.n147 585
R7 B.n146 B.n145 585
R8 B.n144 B.n143 585
R9 B.n142 B.n141 585
R10 B.n140 B.n139 585
R11 B.n138 B.n137 585
R12 B.n136 B.n135 585
R13 B.n134 B.n133 585
R14 B.n132 B.n131 585
R15 B.n130 B.n129 585
R16 B.n128 B.n127 585
R17 B.n126 B.n125 585
R18 B.n124 B.n123 585
R19 B.n122 B.n121 585
R20 B.n120 B.n119 585
R21 B.n118 B.n117 585
R22 B.n116 B.n115 585
R23 B.n114 B.n113 585
R24 B.n112 B.n111 585
R25 B.n110 B.n109 585
R26 B.n108 B.n107 585
R27 B.n106 B.n105 585
R28 B.n104 B.n103 585
R29 B.n101 B.n100 585
R30 B.n99 B.n98 585
R31 B.n97 B.n96 585
R32 B.n95 B.n94 585
R33 B.n93 B.n92 585
R34 B.n91 B.n90 585
R35 B.n89 B.n88 585
R36 B.n87 B.n86 585
R37 B.n85 B.n84 585
R38 B.n83 B.n82 585
R39 B.n81 B.n80 585
R40 B.n79 B.n78 585
R41 B.n77 B.n76 585
R42 B.n75 B.n74 585
R43 B.n73 B.n72 585
R44 B.n71 B.n70 585
R45 B.n69 B.n68 585
R46 B.n67 B.n66 585
R47 B.n65 B.n64 585
R48 B.n386 B.n34 585
R49 B.n390 B.n34 585
R50 B.n385 B.n33 585
R51 B.n391 B.n33 585
R52 B.n384 B.n383 585
R53 B.n383 B.n29 585
R54 B.n382 B.n28 585
R55 B.n397 B.n28 585
R56 B.n381 B.n27 585
R57 B.n398 B.n27 585
R58 B.n380 B.n26 585
R59 B.n399 B.n26 585
R60 B.n379 B.n378 585
R61 B.n378 B.n22 585
R62 B.n377 B.n21 585
R63 B.n405 B.n21 585
R64 B.n376 B.n20 585
R65 B.n406 B.n20 585
R66 B.n375 B.n19 585
R67 B.n407 B.n19 585
R68 B.n374 B.n373 585
R69 B.n373 B.n15 585
R70 B.n372 B.n14 585
R71 B.n413 B.n14 585
R72 B.n371 B.n13 585
R73 B.n414 B.n13 585
R74 B.n370 B.n12 585
R75 B.n415 B.n12 585
R76 B.n369 B.n368 585
R77 B.n368 B.n367 585
R78 B.n366 B.n365 585
R79 B.n366 B.n8 585
R80 B.n364 B.n7 585
R81 B.n422 B.n7 585
R82 B.n363 B.n6 585
R83 B.n423 B.n6 585
R84 B.n362 B.n5 585
R85 B.n424 B.n5 585
R86 B.n361 B.n360 585
R87 B.n360 B.n4 585
R88 B.n359 B.n156 585
R89 B.n359 B.n358 585
R90 B.n349 B.n157 585
R91 B.n158 B.n157 585
R92 B.n351 B.n350 585
R93 B.n352 B.n351 585
R94 B.n348 B.n163 585
R95 B.n163 B.n162 585
R96 B.n347 B.n346 585
R97 B.n346 B.n345 585
R98 B.n165 B.n164 585
R99 B.n166 B.n165 585
R100 B.n338 B.n337 585
R101 B.n339 B.n338 585
R102 B.n336 B.n171 585
R103 B.n171 B.n170 585
R104 B.n335 B.n334 585
R105 B.n334 B.n333 585
R106 B.n173 B.n172 585
R107 B.n174 B.n173 585
R108 B.n326 B.n325 585
R109 B.n327 B.n326 585
R110 B.n324 B.n179 585
R111 B.n179 B.n178 585
R112 B.n323 B.n322 585
R113 B.n322 B.n321 585
R114 B.n181 B.n180 585
R115 B.n182 B.n181 585
R116 B.n314 B.n313 585
R117 B.n315 B.n314 585
R118 B.n312 B.n187 585
R119 B.n187 B.n186 585
R120 B.n306 B.n305 585
R121 B.n304 B.n212 585
R122 B.n303 B.n211 585
R123 B.n308 B.n211 585
R124 B.n302 B.n301 585
R125 B.n300 B.n299 585
R126 B.n298 B.n297 585
R127 B.n296 B.n295 585
R128 B.n294 B.n293 585
R129 B.n292 B.n291 585
R130 B.n290 B.n289 585
R131 B.n288 B.n287 585
R132 B.n286 B.n285 585
R133 B.n284 B.n283 585
R134 B.n282 B.n281 585
R135 B.n280 B.n279 585
R136 B.n278 B.n277 585
R137 B.n276 B.n275 585
R138 B.n274 B.n273 585
R139 B.n272 B.n271 585
R140 B.n270 B.n269 585
R141 B.n268 B.n267 585
R142 B.n266 B.n265 585
R143 B.n264 B.n263 585
R144 B.n262 B.n261 585
R145 B.n260 B.n259 585
R146 B.n258 B.n257 585
R147 B.n256 B.n255 585
R148 B.n254 B.n253 585
R149 B.n251 B.n250 585
R150 B.n249 B.n248 585
R151 B.n247 B.n246 585
R152 B.n245 B.n244 585
R153 B.n243 B.n242 585
R154 B.n241 B.n240 585
R155 B.n239 B.n238 585
R156 B.n237 B.n236 585
R157 B.n235 B.n234 585
R158 B.n233 B.n232 585
R159 B.n231 B.n230 585
R160 B.n229 B.n228 585
R161 B.n227 B.n226 585
R162 B.n225 B.n224 585
R163 B.n223 B.n222 585
R164 B.n221 B.n220 585
R165 B.n219 B.n218 585
R166 B.n189 B.n188 585
R167 B.n311 B.n310 585
R168 B.n185 B.n184 585
R169 B.n186 B.n185 585
R170 B.n317 B.n316 585
R171 B.n316 B.n315 585
R172 B.n318 B.n183 585
R173 B.n183 B.n182 585
R174 B.n320 B.n319 585
R175 B.n321 B.n320 585
R176 B.n177 B.n176 585
R177 B.n178 B.n177 585
R178 B.n329 B.n328 585
R179 B.n328 B.n327 585
R180 B.n330 B.n175 585
R181 B.n175 B.n174 585
R182 B.n332 B.n331 585
R183 B.n333 B.n332 585
R184 B.n169 B.n168 585
R185 B.n170 B.n169 585
R186 B.n341 B.n340 585
R187 B.n340 B.n339 585
R188 B.n342 B.n167 585
R189 B.n167 B.n166 585
R190 B.n344 B.n343 585
R191 B.n345 B.n344 585
R192 B.n161 B.n160 585
R193 B.n162 B.n161 585
R194 B.n354 B.n353 585
R195 B.n353 B.n352 585
R196 B.n355 B.n159 585
R197 B.n159 B.n158 585
R198 B.n357 B.n356 585
R199 B.n358 B.n357 585
R200 B.n3 B.n0 585
R201 B.n4 B.n3 585
R202 B.n421 B.n1 585
R203 B.n422 B.n421 585
R204 B.n420 B.n419 585
R205 B.n420 B.n8 585
R206 B.n418 B.n9 585
R207 B.n367 B.n9 585
R208 B.n417 B.n416 585
R209 B.n416 B.n415 585
R210 B.n11 B.n10 585
R211 B.n414 B.n11 585
R212 B.n412 B.n411 585
R213 B.n413 B.n412 585
R214 B.n410 B.n16 585
R215 B.n16 B.n15 585
R216 B.n409 B.n408 585
R217 B.n408 B.n407 585
R218 B.n18 B.n17 585
R219 B.n406 B.n18 585
R220 B.n404 B.n403 585
R221 B.n405 B.n404 585
R222 B.n402 B.n23 585
R223 B.n23 B.n22 585
R224 B.n401 B.n400 585
R225 B.n400 B.n399 585
R226 B.n25 B.n24 585
R227 B.n398 B.n25 585
R228 B.n396 B.n395 585
R229 B.n397 B.n396 585
R230 B.n394 B.n30 585
R231 B.n30 B.n29 585
R232 B.n393 B.n392 585
R233 B.n392 B.n391 585
R234 B.n32 B.n31 585
R235 B.n390 B.n32 585
R236 B.n425 B.n424 585
R237 B.n423 B.n2 585
R238 B.n64 B.n32 516.524
R239 B.n388 B.n34 516.524
R240 B.n310 B.n187 516.524
R241 B.n306 B.n185 516.524
R242 B.n62 B.t6 282.099
R243 B.n59 B.t13 282.099
R244 B.n216 B.t10 282.099
R245 B.n213 B.t2 282.099
R246 B.n389 B.n57 256.663
R247 B.n389 B.n56 256.663
R248 B.n389 B.n55 256.663
R249 B.n389 B.n54 256.663
R250 B.n389 B.n53 256.663
R251 B.n389 B.n52 256.663
R252 B.n389 B.n51 256.663
R253 B.n389 B.n50 256.663
R254 B.n389 B.n49 256.663
R255 B.n389 B.n48 256.663
R256 B.n389 B.n47 256.663
R257 B.n389 B.n46 256.663
R258 B.n389 B.n45 256.663
R259 B.n389 B.n44 256.663
R260 B.n389 B.n43 256.663
R261 B.n389 B.n42 256.663
R262 B.n389 B.n41 256.663
R263 B.n389 B.n40 256.663
R264 B.n389 B.n39 256.663
R265 B.n389 B.n38 256.663
R266 B.n389 B.n37 256.663
R267 B.n389 B.n36 256.663
R268 B.n389 B.n35 256.663
R269 B.n308 B.n307 256.663
R270 B.n308 B.n190 256.663
R271 B.n308 B.n191 256.663
R272 B.n308 B.n192 256.663
R273 B.n308 B.n193 256.663
R274 B.n308 B.n194 256.663
R275 B.n308 B.n195 256.663
R276 B.n308 B.n196 256.663
R277 B.n308 B.n197 256.663
R278 B.n308 B.n198 256.663
R279 B.n308 B.n199 256.663
R280 B.n308 B.n200 256.663
R281 B.n308 B.n201 256.663
R282 B.n308 B.n202 256.663
R283 B.n308 B.n203 256.663
R284 B.n308 B.n204 256.663
R285 B.n308 B.n205 256.663
R286 B.n308 B.n206 256.663
R287 B.n308 B.n207 256.663
R288 B.n308 B.n208 256.663
R289 B.n308 B.n209 256.663
R290 B.n308 B.n210 256.663
R291 B.n309 B.n308 256.663
R292 B.n427 B.n426 256.663
R293 B.n68 B.n67 163.367
R294 B.n72 B.n71 163.367
R295 B.n76 B.n75 163.367
R296 B.n80 B.n79 163.367
R297 B.n84 B.n83 163.367
R298 B.n88 B.n87 163.367
R299 B.n92 B.n91 163.367
R300 B.n96 B.n95 163.367
R301 B.n100 B.n99 163.367
R302 B.n105 B.n104 163.367
R303 B.n109 B.n108 163.367
R304 B.n113 B.n112 163.367
R305 B.n117 B.n116 163.367
R306 B.n121 B.n120 163.367
R307 B.n125 B.n124 163.367
R308 B.n129 B.n128 163.367
R309 B.n133 B.n132 163.367
R310 B.n137 B.n136 163.367
R311 B.n141 B.n140 163.367
R312 B.n145 B.n144 163.367
R313 B.n149 B.n148 163.367
R314 B.n153 B.n152 163.367
R315 B.n388 B.n58 163.367
R316 B.n314 B.n187 163.367
R317 B.n314 B.n181 163.367
R318 B.n322 B.n181 163.367
R319 B.n322 B.n179 163.367
R320 B.n326 B.n179 163.367
R321 B.n326 B.n173 163.367
R322 B.n334 B.n173 163.367
R323 B.n334 B.n171 163.367
R324 B.n338 B.n171 163.367
R325 B.n338 B.n165 163.367
R326 B.n346 B.n165 163.367
R327 B.n346 B.n163 163.367
R328 B.n351 B.n163 163.367
R329 B.n351 B.n157 163.367
R330 B.n359 B.n157 163.367
R331 B.n360 B.n359 163.367
R332 B.n360 B.n5 163.367
R333 B.n6 B.n5 163.367
R334 B.n7 B.n6 163.367
R335 B.n366 B.n7 163.367
R336 B.n368 B.n366 163.367
R337 B.n368 B.n12 163.367
R338 B.n13 B.n12 163.367
R339 B.n14 B.n13 163.367
R340 B.n373 B.n14 163.367
R341 B.n373 B.n19 163.367
R342 B.n20 B.n19 163.367
R343 B.n21 B.n20 163.367
R344 B.n378 B.n21 163.367
R345 B.n378 B.n26 163.367
R346 B.n27 B.n26 163.367
R347 B.n28 B.n27 163.367
R348 B.n383 B.n28 163.367
R349 B.n383 B.n33 163.367
R350 B.n34 B.n33 163.367
R351 B.n212 B.n211 163.367
R352 B.n301 B.n211 163.367
R353 B.n299 B.n298 163.367
R354 B.n295 B.n294 163.367
R355 B.n291 B.n290 163.367
R356 B.n287 B.n286 163.367
R357 B.n283 B.n282 163.367
R358 B.n279 B.n278 163.367
R359 B.n275 B.n274 163.367
R360 B.n271 B.n270 163.367
R361 B.n267 B.n266 163.367
R362 B.n263 B.n262 163.367
R363 B.n259 B.n258 163.367
R364 B.n255 B.n254 163.367
R365 B.n250 B.n249 163.367
R366 B.n246 B.n245 163.367
R367 B.n242 B.n241 163.367
R368 B.n238 B.n237 163.367
R369 B.n234 B.n233 163.367
R370 B.n230 B.n229 163.367
R371 B.n226 B.n225 163.367
R372 B.n222 B.n221 163.367
R373 B.n218 B.n189 163.367
R374 B.n316 B.n185 163.367
R375 B.n316 B.n183 163.367
R376 B.n320 B.n183 163.367
R377 B.n320 B.n177 163.367
R378 B.n328 B.n177 163.367
R379 B.n328 B.n175 163.367
R380 B.n332 B.n175 163.367
R381 B.n332 B.n169 163.367
R382 B.n340 B.n169 163.367
R383 B.n340 B.n167 163.367
R384 B.n344 B.n167 163.367
R385 B.n344 B.n161 163.367
R386 B.n353 B.n161 163.367
R387 B.n353 B.n159 163.367
R388 B.n357 B.n159 163.367
R389 B.n357 B.n3 163.367
R390 B.n425 B.n3 163.367
R391 B.n421 B.n2 163.367
R392 B.n421 B.n420 163.367
R393 B.n420 B.n9 163.367
R394 B.n416 B.n9 163.367
R395 B.n416 B.n11 163.367
R396 B.n412 B.n11 163.367
R397 B.n412 B.n16 163.367
R398 B.n408 B.n16 163.367
R399 B.n408 B.n18 163.367
R400 B.n404 B.n18 163.367
R401 B.n404 B.n23 163.367
R402 B.n400 B.n23 163.367
R403 B.n400 B.n25 163.367
R404 B.n396 B.n25 163.367
R405 B.n396 B.n30 163.367
R406 B.n392 B.n30 163.367
R407 B.n392 B.n32 163.367
R408 B.n308 B.n186 159.387
R409 B.n390 B.n389 159.387
R410 B.n59 B.t14 104.703
R411 B.n216 B.t12 104.703
R412 B.n62 B.t8 104.7
R413 B.n213 B.t5 104.7
R414 B.n315 B.n186 79.1121
R415 B.n315 B.n182 79.1121
R416 B.n321 B.n182 79.1121
R417 B.n321 B.n178 79.1121
R418 B.n327 B.n178 79.1121
R419 B.n333 B.n174 79.1121
R420 B.n333 B.n170 79.1121
R421 B.n339 B.n170 79.1121
R422 B.n339 B.n166 79.1121
R423 B.n345 B.n166 79.1121
R424 B.n345 B.n162 79.1121
R425 B.n352 B.n162 79.1121
R426 B.n358 B.n158 79.1121
R427 B.n358 B.n4 79.1121
R428 B.n424 B.n4 79.1121
R429 B.n424 B.n423 79.1121
R430 B.n423 B.n422 79.1121
R431 B.n422 B.n8 79.1121
R432 B.n367 B.n8 79.1121
R433 B.n415 B.n414 79.1121
R434 B.n414 B.n413 79.1121
R435 B.n413 B.n15 79.1121
R436 B.n407 B.n15 79.1121
R437 B.n407 B.n406 79.1121
R438 B.n406 B.n405 79.1121
R439 B.n405 B.n22 79.1121
R440 B.n399 B.n398 79.1121
R441 B.n398 B.n397 79.1121
R442 B.n397 B.n29 79.1121
R443 B.n391 B.n29 79.1121
R444 B.n391 B.n390 79.1121
R445 B.n60 B.t15 73.0907
R446 B.n217 B.t11 73.0907
R447 B.n63 B.t9 73.0869
R448 B.n214 B.t4 73.0869
R449 B.n64 B.n35 71.676
R450 B.n68 B.n36 71.676
R451 B.n72 B.n37 71.676
R452 B.n76 B.n38 71.676
R453 B.n80 B.n39 71.676
R454 B.n84 B.n40 71.676
R455 B.n88 B.n41 71.676
R456 B.n92 B.n42 71.676
R457 B.n96 B.n43 71.676
R458 B.n100 B.n44 71.676
R459 B.n105 B.n45 71.676
R460 B.n109 B.n46 71.676
R461 B.n113 B.n47 71.676
R462 B.n117 B.n48 71.676
R463 B.n121 B.n49 71.676
R464 B.n125 B.n50 71.676
R465 B.n129 B.n51 71.676
R466 B.n133 B.n52 71.676
R467 B.n137 B.n53 71.676
R468 B.n141 B.n54 71.676
R469 B.n145 B.n55 71.676
R470 B.n149 B.n56 71.676
R471 B.n153 B.n57 71.676
R472 B.n58 B.n57 71.676
R473 B.n152 B.n56 71.676
R474 B.n148 B.n55 71.676
R475 B.n144 B.n54 71.676
R476 B.n140 B.n53 71.676
R477 B.n136 B.n52 71.676
R478 B.n132 B.n51 71.676
R479 B.n128 B.n50 71.676
R480 B.n124 B.n49 71.676
R481 B.n120 B.n48 71.676
R482 B.n116 B.n47 71.676
R483 B.n112 B.n46 71.676
R484 B.n108 B.n45 71.676
R485 B.n104 B.n44 71.676
R486 B.n99 B.n43 71.676
R487 B.n95 B.n42 71.676
R488 B.n91 B.n41 71.676
R489 B.n87 B.n40 71.676
R490 B.n83 B.n39 71.676
R491 B.n79 B.n38 71.676
R492 B.n75 B.n37 71.676
R493 B.n71 B.n36 71.676
R494 B.n67 B.n35 71.676
R495 B.n307 B.n306 71.676
R496 B.n301 B.n190 71.676
R497 B.n298 B.n191 71.676
R498 B.n294 B.n192 71.676
R499 B.n290 B.n193 71.676
R500 B.n286 B.n194 71.676
R501 B.n282 B.n195 71.676
R502 B.n278 B.n196 71.676
R503 B.n274 B.n197 71.676
R504 B.n270 B.n198 71.676
R505 B.n266 B.n199 71.676
R506 B.n262 B.n200 71.676
R507 B.n258 B.n201 71.676
R508 B.n254 B.n202 71.676
R509 B.n249 B.n203 71.676
R510 B.n245 B.n204 71.676
R511 B.n241 B.n205 71.676
R512 B.n237 B.n206 71.676
R513 B.n233 B.n207 71.676
R514 B.n229 B.n208 71.676
R515 B.n225 B.n209 71.676
R516 B.n221 B.n210 71.676
R517 B.n309 B.n189 71.676
R518 B.n307 B.n212 71.676
R519 B.n299 B.n190 71.676
R520 B.n295 B.n191 71.676
R521 B.n291 B.n192 71.676
R522 B.n287 B.n193 71.676
R523 B.n283 B.n194 71.676
R524 B.n279 B.n195 71.676
R525 B.n275 B.n196 71.676
R526 B.n271 B.n197 71.676
R527 B.n267 B.n198 71.676
R528 B.n263 B.n199 71.676
R529 B.n259 B.n200 71.676
R530 B.n255 B.n201 71.676
R531 B.n250 B.n202 71.676
R532 B.n246 B.n203 71.676
R533 B.n242 B.n204 71.676
R534 B.n238 B.n205 71.676
R535 B.n234 B.n206 71.676
R536 B.n230 B.n207 71.676
R537 B.n226 B.n208 71.676
R538 B.n222 B.n209 71.676
R539 B.n218 B.n210 71.676
R540 B.n310 B.n309 71.676
R541 B.n426 B.n425 71.676
R542 B.n426 B.n2 71.676
R543 B.n102 B.n63 59.5399
R544 B.n61 B.n60 59.5399
R545 B.n252 B.n217 59.5399
R546 B.n215 B.n214 59.5399
R547 B.n327 B.t3 39.5563
R548 B.t3 B.n174 39.5563
R549 B.n352 B.t1 39.5563
R550 B.t1 B.n158 39.5563
R551 B.n367 B.t0 39.5563
R552 B.n415 B.t0 39.5563
R553 B.t7 B.n22 39.5563
R554 B.n399 B.t7 39.5563
R555 B.n305 B.n184 33.5615
R556 B.n312 B.n311 33.5615
R557 B.n387 B.n386 33.5615
R558 B.n65 B.n31 33.5615
R559 B.n63 B.n62 31.6126
R560 B.n60 B.n59 31.6126
R561 B.n217 B.n216 31.6126
R562 B.n214 B.n213 31.6126
R563 B B.n427 18.0485
R564 B.n317 B.n184 10.6151
R565 B.n318 B.n317 10.6151
R566 B.n319 B.n318 10.6151
R567 B.n319 B.n176 10.6151
R568 B.n329 B.n176 10.6151
R569 B.n330 B.n329 10.6151
R570 B.n331 B.n330 10.6151
R571 B.n331 B.n168 10.6151
R572 B.n341 B.n168 10.6151
R573 B.n342 B.n341 10.6151
R574 B.n343 B.n342 10.6151
R575 B.n343 B.n160 10.6151
R576 B.n354 B.n160 10.6151
R577 B.n355 B.n354 10.6151
R578 B.n356 B.n355 10.6151
R579 B.n356 B.n0 10.6151
R580 B.n305 B.n304 10.6151
R581 B.n304 B.n303 10.6151
R582 B.n303 B.n302 10.6151
R583 B.n302 B.n300 10.6151
R584 B.n300 B.n297 10.6151
R585 B.n297 B.n296 10.6151
R586 B.n296 B.n293 10.6151
R587 B.n293 B.n292 10.6151
R588 B.n292 B.n289 10.6151
R589 B.n289 B.n288 10.6151
R590 B.n288 B.n285 10.6151
R591 B.n285 B.n284 10.6151
R592 B.n284 B.n281 10.6151
R593 B.n281 B.n280 10.6151
R594 B.n280 B.n277 10.6151
R595 B.n277 B.n276 10.6151
R596 B.n276 B.n273 10.6151
R597 B.n273 B.n272 10.6151
R598 B.n269 B.n268 10.6151
R599 B.n268 B.n265 10.6151
R600 B.n265 B.n264 10.6151
R601 B.n264 B.n261 10.6151
R602 B.n261 B.n260 10.6151
R603 B.n260 B.n257 10.6151
R604 B.n257 B.n256 10.6151
R605 B.n256 B.n253 10.6151
R606 B.n251 B.n248 10.6151
R607 B.n248 B.n247 10.6151
R608 B.n247 B.n244 10.6151
R609 B.n244 B.n243 10.6151
R610 B.n243 B.n240 10.6151
R611 B.n240 B.n239 10.6151
R612 B.n239 B.n236 10.6151
R613 B.n236 B.n235 10.6151
R614 B.n235 B.n232 10.6151
R615 B.n232 B.n231 10.6151
R616 B.n231 B.n228 10.6151
R617 B.n228 B.n227 10.6151
R618 B.n227 B.n224 10.6151
R619 B.n224 B.n223 10.6151
R620 B.n223 B.n220 10.6151
R621 B.n220 B.n219 10.6151
R622 B.n219 B.n188 10.6151
R623 B.n311 B.n188 10.6151
R624 B.n313 B.n312 10.6151
R625 B.n313 B.n180 10.6151
R626 B.n323 B.n180 10.6151
R627 B.n324 B.n323 10.6151
R628 B.n325 B.n324 10.6151
R629 B.n325 B.n172 10.6151
R630 B.n335 B.n172 10.6151
R631 B.n336 B.n335 10.6151
R632 B.n337 B.n336 10.6151
R633 B.n337 B.n164 10.6151
R634 B.n347 B.n164 10.6151
R635 B.n348 B.n347 10.6151
R636 B.n350 B.n348 10.6151
R637 B.n350 B.n349 10.6151
R638 B.n349 B.n156 10.6151
R639 B.n361 B.n156 10.6151
R640 B.n362 B.n361 10.6151
R641 B.n363 B.n362 10.6151
R642 B.n364 B.n363 10.6151
R643 B.n365 B.n364 10.6151
R644 B.n369 B.n365 10.6151
R645 B.n370 B.n369 10.6151
R646 B.n371 B.n370 10.6151
R647 B.n372 B.n371 10.6151
R648 B.n374 B.n372 10.6151
R649 B.n375 B.n374 10.6151
R650 B.n376 B.n375 10.6151
R651 B.n377 B.n376 10.6151
R652 B.n379 B.n377 10.6151
R653 B.n380 B.n379 10.6151
R654 B.n381 B.n380 10.6151
R655 B.n382 B.n381 10.6151
R656 B.n384 B.n382 10.6151
R657 B.n385 B.n384 10.6151
R658 B.n386 B.n385 10.6151
R659 B.n419 B.n1 10.6151
R660 B.n419 B.n418 10.6151
R661 B.n418 B.n417 10.6151
R662 B.n417 B.n10 10.6151
R663 B.n411 B.n10 10.6151
R664 B.n411 B.n410 10.6151
R665 B.n410 B.n409 10.6151
R666 B.n409 B.n17 10.6151
R667 B.n403 B.n17 10.6151
R668 B.n403 B.n402 10.6151
R669 B.n402 B.n401 10.6151
R670 B.n401 B.n24 10.6151
R671 B.n395 B.n24 10.6151
R672 B.n395 B.n394 10.6151
R673 B.n394 B.n393 10.6151
R674 B.n393 B.n31 10.6151
R675 B.n66 B.n65 10.6151
R676 B.n69 B.n66 10.6151
R677 B.n70 B.n69 10.6151
R678 B.n73 B.n70 10.6151
R679 B.n74 B.n73 10.6151
R680 B.n77 B.n74 10.6151
R681 B.n78 B.n77 10.6151
R682 B.n81 B.n78 10.6151
R683 B.n82 B.n81 10.6151
R684 B.n85 B.n82 10.6151
R685 B.n86 B.n85 10.6151
R686 B.n89 B.n86 10.6151
R687 B.n90 B.n89 10.6151
R688 B.n93 B.n90 10.6151
R689 B.n94 B.n93 10.6151
R690 B.n97 B.n94 10.6151
R691 B.n98 B.n97 10.6151
R692 B.n101 B.n98 10.6151
R693 B.n106 B.n103 10.6151
R694 B.n107 B.n106 10.6151
R695 B.n110 B.n107 10.6151
R696 B.n111 B.n110 10.6151
R697 B.n114 B.n111 10.6151
R698 B.n115 B.n114 10.6151
R699 B.n118 B.n115 10.6151
R700 B.n119 B.n118 10.6151
R701 B.n123 B.n122 10.6151
R702 B.n126 B.n123 10.6151
R703 B.n127 B.n126 10.6151
R704 B.n130 B.n127 10.6151
R705 B.n131 B.n130 10.6151
R706 B.n134 B.n131 10.6151
R707 B.n135 B.n134 10.6151
R708 B.n138 B.n135 10.6151
R709 B.n139 B.n138 10.6151
R710 B.n142 B.n139 10.6151
R711 B.n143 B.n142 10.6151
R712 B.n146 B.n143 10.6151
R713 B.n147 B.n146 10.6151
R714 B.n150 B.n147 10.6151
R715 B.n151 B.n150 10.6151
R716 B.n154 B.n151 10.6151
R717 B.n155 B.n154 10.6151
R718 B.n387 B.n155 10.6151
R719 B.n427 B.n0 8.11757
R720 B.n427 B.n1 8.11757
R721 B.n269 B.n215 6.5566
R722 B.n253 B.n252 6.5566
R723 B.n103 B.n102 6.5566
R724 B.n119 B.n61 6.5566
R725 B.n272 B.n215 4.05904
R726 B.n252 B.n251 4.05904
R727 B.n102 B.n101 4.05904
R728 B.n122 B.n61 4.05904
R729 VP.n0 VP.t0 223.597
R730 VP.n0 VP.t1 188.312
R731 VP VP.n0 0.146778
R732 VTAIL.n1 VTAIL.t1 59.5886
R733 VTAIL.n2 VTAIL.t3 59.5884
R734 VTAIL.n3 VTAIL.t0 59.5884
R735 VTAIL.n0 VTAIL.t2 59.5884
R736 VTAIL.n1 VTAIL.n0 18.7807
R737 VTAIL.n3 VTAIL.n2 17.3755
R738 VTAIL.n2 VTAIL.n1 1.17291
R739 VTAIL VTAIL.n0 0.87981
R740 VTAIL VTAIL.n3 0.293603
R741 VDD1 VDD1.t0 107.216
R742 VDD1 VDD1.t1 76.6767
R743 VN VN.t0 223.882
R744 VN VN.t1 188.458
R745 VDD2.n0 VDD2.t0 106.341
R746 VDD2.n0 VDD2.t1 76.2672
R747 VDD2 VDD2.n0 0.409983
C0 VP VTAIL 0.993336f
C1 VTAIL VN 0.979108f
C2 VP VDD2 0.2825f
C3 VDD2 VN 0.999261f
C4 VP VDD1 1.128f
C5 VN VDD1 0.152003f
C6 VDD2 VTAIL 2.76402f
C7 VTAIL VDD1 2.7211f
C8 VP VN 3.40117f
C9 VDD2 VDD1 0.522507f
C10 VDD2 B 2.53563f
C11 VDD1 B 4.14138f
C12 VTAIL B 3.472632f
C13 VN B 6.27446f
C14 VP B 4.128953f
C15 VDD2.t0 B 0.720529f
C16 VDD2.t1 B 0.519868f
C17 VDD2.n0 B 1.50306f
C18 VN.t1 B 0.585735f
C19 VN.t0 B 0.759609f
C20 VDD1.t1 B 0.492066f
C21 VDD1.t0 B 0.696058f
C22 VTAIL.t2 B 0.542248f
C23 VTAIL.n0 B 0.856195f
C24 VTAIL.t1 B 0.54225f
C25 VTAIL.n1 B 0.872974f
C26 VTAIL.t3 B 0.542248f
C27 VTAIL.n2 B 0.792529f
C28 VTAIL.t0 B 0.542248f
C29 VTAIL.n3 B 0.742187f
C30 VP.t0 B 0.765228f
C31 VP.t1 B 0.593004f
C32 VP.n0 B 2.01379f
.ends

