* NGSPICE file created from diff_pair_sample_0039.ext - technology: sky130A

.subckt diff_pair_sample_0039 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=3.1977 ps=19.71 w=19.38 l=1.56
X1 VDD1.t8 VP.t1 VTAIL.t13 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=7.5582 ps=39.54 w=19.38 l=1.56
X2 VTAIL.t15 VP.t2 VDD1.t7 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X3 VTAIL.t17 VP.t3 VDD1.t6 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X4 VDD2.t9 VN.t0 VTAIL.t8 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X5 VDD2.t8 VN.t1 VTAIL.t5 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=3.1977 ps=19.71 w=19.38 l=1.56
X6 VTAIL.t2 VN.t2 VDD2.t7 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X7 VDD2.t6 VN.t3 VTAIL.t9 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X8 B.t11 B.t9 B.t10 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=0 ps=0 w=19.38 l=1.56
X9 VTAIL.t7 VN.t4 VDD2.t5 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X10 VTAIL.t14 VP.t4 VDD1.t5 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X11 B.t8 B.t6 B.t7 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=0 ps=0 w=19.38 l=1.56
X12 VDD2.t4 VN.t5 VTAIL.t0 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=7.5582 ps=39.54 w=19.38 l=1.56
X13 VTAIL.t3 VN.t6 VDD2.t3 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X14 VDD1.t4 VP.t5 VTAIL.t18 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=7.5582 ps=39.54 w=19.38 l=1.56
X15 VDD1.t3 VP.t6 VTAIL.t12 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X16 VDD2.t2 VN.t7 VTAIL.t4 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=7.5582 ps=39.54 w=19.38 l=1.56
X17 VTAIL.t16 VP.t7 VDD1.t2 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X18 VDD1.t1 VP.t8 VTAIL.t19 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=3.1977 ps=19.71 w=19.38 l=1.56
X19 B.t5 B.t3 B.t4 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=0 ps=0 w=19.38 l=1.56
X20 VDD2.t1 VN.t8 VTAIL.t6 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=3.1977 ps=19.71 w=19.38 l=1.56
X21 VTAIL.t1 VN.t9 VDD2.t0 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X22 VDD1.t0 VP.t9 VTAIL.t11 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=3.1977 pd=19.71 as=3.1977 ps=19.71 w=19.38 l=1.56
X23 B.t2 B.t0 B.t1 w_n3238_n4844# sky130_fd_pr__pfet_01v8 ad=7.5582 pd=39.54 as=0 ps=0 w=19.38 l=1.56
R0 VP.n14 VP.t8 327.947
R1 VP.n39 VP.t0 299.397
R2 VP.n46 VP.t4 299.397
R3 VP.n53 VP.t9 299.397
R4 VP.n60 VP.t3 299.397
R5 VP.n67 VP.t5 299.397
R6 VP.n36 VP.t1 299.397
R7 VP.n29 VP.t2 299.397
R8 VP.n22 VP.t6 299.397
R9 VP.n15 VP.t7 299.397
R10 VP.n39 VP.n38 184.417
R11 VP.n68 VP.n67 184.417
R12 VP.n37 VP.n36 184.417
R13 VP.n17 VP.n16 161.3
R14 VP.n18 VP.n13 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n12 161.3
R17 VP.n24 VP.n23 161.3
R18 VP.n25 VP.n11 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n28 VP.n10 161.3
R21 VP.n31 VP.n30 161.3
R22 VP.n32 VP.n9 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n35 VP.n8 161.3
R25 VP.n66 VP.n0 161.3
R26 VP.n65 VP.n64 161.3
R27 VP.n63 VP.n1 161.3
R28 VP.n62 VP.n61 161.3
R29 VP.n59 VP.n2 161.3
R30 VP.n58 VP.n57 161.3
R31 VP.n56 VP.n3 161.3
R32 VP.n55 VP.n54 161.3
R33 VP.n52 VP.n4 161.3
R34 VP.n51 VP.n50 161.3
R35 VP.n49 VP.n5 161.3
R36 VP.n48 VP.n47 161.3
R37 VP.n45 VP.n6 161.3
R38 VP.n44 VP.n43 161.3
R39 VP.n42 VP.n7 161.3
R40 VP.n41 VP.n40 161.3
R41 VP.n15 VP.n14 60.7346
R42 VP.n51 VP.n5 56.5617
R43 VP.n58 VP.n3 56.5617
R44 VP.n27 VP.n11 56.5617
R45 VP.n20 VP.n13 56.5617
R46 VP.n38 VP.n37 52.8603
R47 VP.n44 VP.n7 48.8116
R48 VP.n65 VP.n1 48.8116
R49 VP.n34 VP.n9 48.8116
R50 VP.n45 VP.n44 32.3425
R51 VP.n61 VP.n1 32.3425
R52 VP.n30 VP.n9 32.3425
R53 VP.n40 VP.n7 24.5923
R54 VP.n47 VP.n5 24.5923
R55 VP.n52 VP.n51 24.5923
R56 VP.n54 VP.n3 24.5923
R57 VP.n59 VP.n58 24.5923
R58 VP.n66 VP.n65 24.5923
R59 VP.n35 VP.n34 24.5923
R60 VP.n28 VP.n27 24.5923
R61 VP.n21 VP.n20 24.5923
R62 VP.n23 VP.n11 24.5923
R63 VP.n16 VP.n13 24.5923
R64 VP.n17 VP.n14 18.7424
R65 VP.n46 VP.n45 17.7066
R66 VP.n61 VP.n60 17.7066
R67 VP.n30 VP.n29 17.7066
R68 VP.n53 VP.n52 12.2964
R69 VP.n54 VP.n53 12.2964
R70 VP.n22 VP.n21 12.2964
R71 VP.n23 VP.n22 12.2964
R72 VP.n47 VP.n46 6.88621
R73 VP.n60 VP.n59 6.88621
R74 VP.n29 VP.n28 6.88621
R75 VP.n16 VP.n15 6.88621
R76 VP.n40 VP.n39 1.47601
R77 VP.n67 VP.n66 1.47601
R78 VP.n36 VP.n35 1.47601
R79 VP.n18 VP.n17 0.189894
R80 VP.n19 VP.n18 0.189894
R81 VP.n19 VP.n12 0.189894
R82 VP.n24 VP.n12 0.189894
R83 VP.n25 VP.n24 0.189894
R84 VP.n26 VP.n25 0.189894
R85 VP.n26 VP.n10 0.189894
R86 VP.n31 VP.n10 0.189894
R87 VP.n32 VP.n31 0.189894
R88 VP.n33 VP.n32 0.189894
R89 VP.n33 VP.n8 0.189894
R90 VP.n37 VP.n8 0.189894
R91 VP.n41 VP.n38 0.189894
R92 VP.n42 VP.n41 0.189894
R93 VP.n43 VP.n42 0.189894
R94 VP.n43 VP.n6 0.189894
R95 VP.n48 VP.n6 0.189894
R96 VP.n49 VP.n48 0.189894
R97 VP.n50 VP.n49 0.189894
R98 VP.n50 VP.n4 0.189894
R99 VP.n55 VP.n4 0.189894
R100 VP.n56 VP.n55 0.189894
R101 VP.n57 VP.n56 0.189894
R102 VP.n57 VP.n2 0.189894
R103 VP.n62 VP.n2 0.189894
R104 VP.n63 VP.n62 0.189894
R105 VP.n64 VP.n63 0.189894
R106 VP.n64 VP.n0 0.189894
R107 VP.n68 VP.n0 0.189894
R108 VP VP.n68 0.0516364
R109 VTAIL.n11 VTAIL.t4 54.406
R110 VTAIL.n17 VTAIL.t0 54.4057
R111 VTAIL.n2 VTAIL.t18 54.4057
R112 VTAIL.n16 VTAIL.t13 54.4057
R113 VTAIL.n15 VTAIL.n14 52.7287
R114 VTAIL.n13 VTAIL.n12 52.7287
R115 VTAIL.n10 VTAIL.n9 52.7287
R116 VTAIL.n8 VTAIL.n7 52.7287
R117 VTAIL.n19 VTAIL.n18 52.7287
R118 VTAIL.n1 VTAIL.n0 52.7287
R119 VTAIL.n4 VTAIL.n3 52.7287
R120 VTAIL.n6 VTAIL.n5 52.7287
R121 VTAIL.n8 VTAIL.n6 32.3324
R122 VTAIL.n17 VTAIL.n16 30.7031
R123 VTAIL.n18 VTAIL.t9 1.67774
R124 VTAIL.n18 VTAIL.t1 1.67774
R125 VTAIL.n0 VTAIL.t6 1.67774
R126 VTAIL.n0 VTAIL.t7 1.67774
R127 VTAIL.n3 VTAIL.t11 1.67774
R128 VTAIL.n3 VTAIL.t17 1.67774
R129 VTAIL.n5 VTAIL.t10 1.67774
R130 VTAIL.n5 VTAIL.t14 1.67774
R131 VTAIL.n14 VTAIL.t12 1.67774
R132 VTAIL.n14 VTAIL.t15 1.67774
R133 VTAIL.n12 VTAIL.t19 1.67774
R134 VTAIL.n12 VTAIL.t16 1.67774
R135 VTAIL.n9 VTAIL.t8 1.67774
R136 VTAIL.n9 VTAIL.t3 1.67774
R137 VTAIL.n7 VTAIL.t5 1.67774
R138 VTAIL.n7 VTAIL.t2 1.67774
R139 VTAIL.n10 VTAIL.n8 1.62981
R140 VTAIL.n11 VTAIL.n10 1.62981
R141 VTAIL.n15 VTAIL.n13 1.62981
R142 VTAIL.n16 VTAIL.n15 1.62981
R143 VTAIL.n6 VTAIL.n4 1.62981
R144 VTAIL.n4 VTAIL.n2 1.62981
R145 VTAIL.n19 VTAIL.n17 1.62981
R146 VTAIL.n13 VTAIL.n11 1.28498
R147 VTAIL.n2 VTAIL.n1 1.28498
R148 VTAIL VTAIL.n1 1.28067
R149 VTAIL VTAIL.n19 0.349638
R150 VDD1.n1 VDD1.t1 72.7141
R151 VDD1.n3 VDD1.t9 72.7138
R152 VDD1.n5 VDD1.n4 70.5741
R153 VDD1.n1 VDD1.n0 69.4075
R154 VDD1.n3 VDD1.n2 69.4075
R155 VDD1.n7 VDD1.n6 69.4073
R156 VDD1.n7 VDD1.n5 49.5591
R157 VDD1.n6 VDD1.t7 1.67774
R158 VDD1.n6 VDD1.t8 1.67774
R159 VDD1.n0 VDD1.t2 1.67774
R160 VDD1.n0 VDD1.t3 1.67774
R161 VDD1.n4 VDD1.t6 1.67774
R162 VDD1.n4 VDD1.t4 1.67774
R163 VDD1.n2 VDD1.t5 1.67774
R164 VDD1.n2 VDD1.t0 1.67774
R165 VDD1 VDD1.n7 1.16429
R166 VDD1 VDD1.n1 0.466017
R167 VDD1.n5 VDD1.n3 0.352482
R168 VN.n6 VN.t8 327.947
R169 VN.n36 VN.t7 327.947
R170 VN.n7 VN.t4 299.397
R171 VN.n14 VN.t3 299.397
R172 VN.n21 VN.t9 299.397
R173 VN.n28 VN.t5 299.397
R174 VN.n37 VN.t6 299.397
R175 VN.n44 VN.t0 299.397
R176 VN.n51 VN.t2 299.397
R177 VN.n58 VN.t1 299.397
R178 VN.n29 VN.n28 184.417
R179 VN.n59 VN.n58 184.417
R180 VN.n57 VN.n30 161.3
R181 VN.n56 VN.n55 161.3
R182 VN.n54 VN.n31 161.3
R183 VN.n53 VN.n52 161.3
R184 VN.n50 VN.n32 161.3
R185 VN.n49 VN.n48 161.3
R186 VN.n47 VN.n33 161.3
R187 VN.n46 VN.n45 161.3
R188 VN.n43 VN.n34 161.3
R189 VN.n42 VN.n41 161.3
R190 VN.n40 VN.n35 161.3
R191 VN.n39 VN.n38 161.3
R192 VN.n27 VN.n0 161.3
R193 VN.n26 VN.n25 161.3
R194 VN.n24 VN.n1 161.3
R195 VN.n23 VN.n22 161.3
R196 VN.n20 VN.n2 161.3
R197 VN.n19 VN.n18 161.3
R198 VN.n17 VN.n3 161.3
R199 VN.n16 VN.n15 161.3
R200 VN.n13 VN.n4 161.3
R201 VN.n12 VN.n11 161.3
R202 VN.n10 VN.n5 161.3
R203 VN.n9 VN.n8 161.3
R204 VN.n7 VN.n6 60.7346
R205 VN.n37 VN.n36 60.7346
R206 VN.n12 VN.n5 56.5617
R207 VN.n19 VN.n3 56.5617
R208 VN.n42 VN.n35 56.5617
R209 VN.n49 VN.n33 56.5617
R210 VN VN.n59 53.241
R211 VN.n26 VN.n1 48.8116
R212 VN.n56 VN.n31 48.8116
R213 VN.n22 VN.n1 32.3425
R214 VN.n52 VN.n31 32.3425
R215 VN.n8 VN.n5 24.5923
R216 VN.n13 VN.n12 24.5923
R217 VN.n15 VN.n3 24.5923
R218 VN.n20 VN.n19 24.5923
R219 VN.n27 VN.n26 24.5923
R220 VN.n38 VN.n35 24.5923
R221 VN.n45 VN.n33 24.5923
R222 VN.n43 VN.n42 24.5923
R223 VN.n50 VN.n49 24.5923
R224 VN.n57 VN.n56 24.5923
R225 VN.n39 VN.n36 18.7424
R226 VN.n9 VN.n6 18.7424
R227 VN.n22 VN.n21 17.7066
R228 VN.n52 VN.n51 17.7066
R229 VN.n14 VN.n13 12.2964
R230 VN.n15 VN.n14 12.2964
R231 VN.n45 VN.n44 12.2964
R232 VN.n44 VN.n43 12.2964
R233 VN.n8 VN.n7 6.88621
R234 VN.n21 VN.n20 6.88621
R235 VN.n38 VN.n37 6.88621
R236 VN.n51 VN.n50 6.88621
R237 VN.n28 VN.n27 1.47601
R238 VN.n58 VN.n57 1.47601
R239 VN.n59 VN.n30 0.189894
R240 VN.n55 VN.n30 0.189894
R241 VN.n55 VN.n54 0.189894
R242 VN.n54 VN.n53 0.189894
R243 VN.n53 VN.n32 0.189894
R244 VN.n48 VN.n32 0.189894
R245 VN.n48 VN.n47 0.189894
R246 VN.n47 VN.n46 0.189894
R247 VN.n46 VN.n34 0.189894
R248 VN.n41 VN.n34 0.189894
R249 VN.n41 VN.n40 0.189894
R250 VN.n40 VN.n39 0.189894
R251 VN.n10 VN.n9 0.189894
R252 VN.n11 VN.n10 0.189894
R253 VN.n11 VN.n4 0.189894
R254 VN.n16 VN.n4 0.189894
R255 VN.n17 VN.n16 0.189894
R256 VN.n18 VN.n17 0.189894
R257 VN.n18 VN.n2 0.189894
R258 VN.n23 VN.n2 0.189894
R259 VN.n24 VN.n23 0.189894
R260 VN.n25 VN.n24 0.189894
R261 VN.n25 VN.n0 0.189894
R262 VN.n29 VN.n0 0.189894
R263 VN VN.n29 0.0516364
R264 VDD2.n1 VDD2.t1 72.7138
R265 VDD2.n4 VDD2.t8 71.0848
R266 VDD2.n3 VDD2.n2 70.5741
R267 VDD2 VDD2.n7 70.5711
R268 VDD2.n6 VDD2.n5 69.4075
R269 VDD2.n1 VDD2.n0 69.4075
R270 VDD2.n4 VDD2.n3 48.1614
R271 VDD2.n7 VDD2.t3 1.67774
R272 VDD2.n7 VDD2.t2 1.67774
R273 VDD2.n5 VDD2.t7 1.67774
R274 VDD2.n5 VDD2.t9 1.67774
R275 VDD2.n2 VDD2.t0 1.67774
R276 VDD2.n2 VDD2.t4 1.67774
R277 VDD2.n0 VDD2.t5 1.67774
R278 VDD2.n0 VDD2.t6 1.67774
R279 VDD2.n6 VDD2.n4 1.62981
R280 VDD2 VDD2.n6 0.466017
R281 VDD2.n3 VDD2.n1 0.352482
R282 B.n494 B.n137 585
R283 B.n493 B.n492 585
R284 B.n491 B.n138 585
R285 B.n490 B.n489 585
R286 B.n488 B.n139 585
R287 B.n487 B.n486 585
R288 B.n485 B.n140 585
R289 B.n484 B.n483 585
R290 B.n482 B.n141 585
R291 B.n481 B.n480 585
R292 B.n479 B.n142 585
R293 B.n478 B.n477 585
R294 B.n476 B.n143 585
R295 B.n475 B.n474 585
R296 B.n473 B.n144 585
R297 B.n472 B.n471 585
R298 B.n470 B.n145 585
R299 B.n469 B.n468 585
R300 B.n467 B.n146 585
R301 B.n466 B.n465 585
R302 B.n464 B.n147 585
R303 B.n463 B.n462 585
R304 B.n461 B.n148 585
R305 B.n460 B.n459 585
R306 B.n458 B.n149 585
R307 B.n457 B.n456 585
R308 B.n455 B.n150 585
R309 B.n454 B.n453 585
R310 B.n452 B.n151 585
R311 B.n451 B.n450 585
R312 B.n449 B.n152 585
R313 B.n448 B.n447 585
R314 B.n446 B.n153 585
R315 B.n445 B.n444 585
R316 B.n443 B.n154 585
R317 B.n442 B.n441 585
R318 B.n440 B.n155 585
R319 B.n439 B.n438 585
R320 B.n437 B.n156 585
R321 B.n436 B.n435 585
R322 B.n434 B.n157 585
R323 B.n433 B.n432 585
R324 B.n431 B.n158 585
R325 B.n430 B.n429 585
R326 B.n428 B.n159 585
R327 B.n427 B.n426 585
R328 B.n425 B.n160 585
R329 B.n424 B.n423 585
R330 B.n422 B.n161 585
R331 B.n421 B.n420 585
R332 B.n419 B.n162 585
R333 B.n418 B.n417 585
R334 B.n416 B.n163 585
R335 B.n415 B.n414 585
R336 B.n413 B.n164 585
R337 B.n412 B.n411 585
R338 B.n410 B.n165 585
R339 B.n409 B.n408 585
R340 B.n407 B.n166 585
R341 B.n406 B.n405 585
R342 B.n404 B.n167 585
R343 B.n403 B.n402 585
R344 B.n401 B.n168 585
R345 B.n400 B.n399 585
R346 B.n395 B.n169 585
R347 B.n394 B.n393 585
R348 B.n392 B.n170 585
R349 B.n391 B.n390 585
R350 B.n389 B.n171 585
R351 B.n388 B.n387 585
R352 B.n386 B.n172 585
R353 B.n385 B.n384 585
R354 B.n383 B.n173 585
R355 B.n381 B.n380 585
R356 B.n379 B.n176 585
R357 B.n378 B.n377 585
R358 B.n376 B.n177 585
R359 B.n375 B.n374 585
R360 B.n373 B.n178 585
R361 B.n372 B.n371 585
R362 B.n370 B.n179 585
R363 B.n369 B.n368 585
R364 B.n367 B.n180 585
R365 B.n366 B.n365 585
R366 B.n364 B.n181 585
R367 B.n363 B.n362 585
R368 B.n361 B.n182 585
R369 B.n360 B.n359 585
R370 B.n358 B.n183 585
R371 B.n357 B.n356 585
R372 B.n355 B.n184 585
R373 B.n354 B.n353 585
R374 B.n352 B.n185 585
R375 B.n351 B.n350 585
R376 B.n349 B.n186 585
R377 B.n348 B.n347 585
R378 B.n346 B.n187 585
R379 B.n345 B.n344 585
R380 B.n343 B.n188 585
R381 B.n342 B.n341 585
R382 B.n340 B.n189 585
R383 B.n339 B.n338 585
R384 B.n337 B.n190 585
R385 B.n336 B.n335 585
R386 B.n334 B.n191 585
R387 B.n333 B.n332 585
R388 B.n331 B.n192 585
R389 B.n330 B.n329 585
R390 B.n328 B.n193 585
R391 B.n327 B.n326 585
R392 B.n325 B.n194 585
R393 B.n324 B.n323 585
R394 B.n322 B.n195 585
R395 B.n321 B.n320 585
R396 B.n319 B.n196 585
R397 B.n318 B.n317 585
R398 B.n316 B.n197 585
R399 B.n315 B.n314 585
R400 B.n313 B.n198 585
R401 B.n312 B.n311 585
R402 B.n310 B.n199 585
R403 B.n309 B.n308 585
R404 B.n307 B.n200 585
R405 B.n306 B.n305 585
R406 B.n304 B.n201 585
R407 B.n303 B.n302 585
R408 B.n301 B.n202 585
R409 B.n300 B.n299 585
R410 B.n298 B.n203 585
R411 B.n297 B.n296 585
R412 B.n295 B.n204 585
R413 B.n294 B.n293 585
R414 B.n292 B.n205 585
R415 B.n291 B.n290 585
R416 B.n289 B.n206 585
R417 B.n288 B.n287 585
R418 B.n496 B.n495 585
R419 B.n497 B.n136 585
R420 B.n499 B.n498 585
R421 B.n500 B.n135 585
R422 B.n502 B.n501 585
R423 B.n503 B.n134 585
R424 B.n505 B.n504 585
R425 B.n506 B.n133 585
R426 B.n508 B.n507 585
R427 B.n509 B.n132 585
R428 B.n511 B.n510 585
R429 B.n512 B.n131 585
R430 B.n514 B.n513 585
R431 B.n515 B.n130 585
R432 B.n517 B.n516 585
R433 B.n518 B.n129 585
R434 B.n520 B.n519 585
R435 B.n521 B.n128 585
R436 B.n523 B.n522 585
R437 B.n524 B.n127 585
R438 B.n526 B.n525 585
R439 B.n527 B.n126 585
R440 B.n529 B.n528 585
R441 B.n530 B.n125 585
R442 B.n532 B.n531 585
R443 B.n533 B.n124 585
R444 B.n535 B.n534 585
R445 B.n536 B.n123 585
R446 B.n538 B.n537 585
R447 B.n539 B.n122 585
R448 B.n541 B.n540 585
R449 B.n542 B.n121 585
R450 B.n544 B.n543 585
R451 B.n545 B.n120 585
R452 B.n547 B.n546 585
R453 B.n548 B.n119 585
R454 B.n550 B.n549 585
R455 B.n551 B.n118 585
R456 B.n553 B.n552 585
R457 B.n554 B.n117 585
R458 B.n556 B.n555 585
R459 B.n557 B.n116 585
R460 B.n559 B.n558 585
R461 B.n560 B.n115 585
R462 B.n562 B.n561 585
R463 B.n563 B.n114 585
R464 B.n565 B.n564 585
R465 B.n566 B.n113 585
R466 B.n568 B.n567 585
R467 B.n569 B.n112 585
R468 B.n571 B.n570 585
R469 B.n572 B.n111 585
R470 B.n574 B.n573 585
R471 B.n575 B.n110 585
R472 B.n577 B.n576 585
R473 B.n578 B.n109 585
R474 B.n580 B.n579 585
R475 B.n581 B.n108 585
R476 B.n583 B.n582 585
R477 B.n584 B.n107 585
R478 B.n586 B.n585 585
R479 B.n587 B.n106 585
R480 B.n589 B.n588 585
R481 B.n590 B.n105 585
R482 B.n592 B.n591 585
R483 B.n593 B.n104 585
R484 B.n595 B.n594 585
R485 B.n596 B.n103 585
R486 B.n598 B.n597 585
R487 B.n599 B.n102 585
R488 B.n601 B.n600 585
R489 B.n602 B.n101 585
R490 B.n604 B.n603 585
R491 B.n605 B.n100 585
R492 B.n607 B.n606 585
R493 B.n608 B.n99 585
R494 B.n610 B.n609 585
R495 B.n611 B.n98 585
R496 B.n613 B.n612 585
R497 B.n614 B.n97 585
R498 B.n616 B.n615 585
R499 B.n617 B.n96 585
R500 B.n619 B.n618 585
R501 B.n620 B.n95 585
R502 B.n826 B.n825 585
R503 B.n824 B.n23 585
R504 B.n823 B.n822 585
R505 B.n821 B.n24 585
R506 B.n820 B.n819 585
R507 B.n818 B.n25 585
R508 B.n817 B.n816 585
R509 B.n815 B.n26 585
R510 B.n814 B.n813 585
R511 B.n812 B.n27 585
R512 B.n811 B.n810 585
R513 B.n809 B.n28 585
R514 B.n808 B.n807 585
R515 B.n806 B.n29 585
R516 B.n805 B.n804 585
R517 B.n803 B.n30 585
R518 B.n802 B.n801 585
R519 B.n800 B.n31 585
R520 B.n799 B.n798 585
R521 B.n797 B.n32 585
R522 B.n796 B.n795 585
R523 B.n794 B.n33 585
R524 B.n793 B.n792 585
R525 B.n791 B.n34 585
R526 B.n790 B.n789 585
R527 B.n788 B.n35 585
R528 B.n787 B.n786 585
R529 B.n785 B.n36 585
R530 B.n784 B.n783 585
R531 B.n782 B.n37 585
R532 B.n781 B.n780 585
R533 B.n779 B.n38 585
R534 B.n778 B.n777 585
R535 B.n776 B.n39 585
R536 B.n775 B.n774 585
R537 B.n773 B.n40 585
R538 B.n772 B.n771 585
R539 B.n770 B.n41 585
R540 B.n769 B.n768 585
R541 B.n767 B.n42 585
R542 B.n766 B.n765 585
R543 B.n764 B.n43 585
R544 B.n763 B.n762 585
R545 B.n761 B.n44 585
R546 B.n760 B.n759 585
R547 B.n758 B.n45 585
R548 B.n757 B.n756 585
R549 B.n755 B.n46 585
R550 B.n754 B.n753 585
R551 B.n752 B.n47 585
R552 B.n751 B.n750 585
R553 B.n749 B.n48 585
R554 B.n748 B.n747 585
R555 B.n746 B.n49 585
R556 B.n745 B.n744 585
R557 B.n743 B.n50 585
R558 B.n742 B.n741 585
R559 B.n740 B.n51 585
R560 B.n739 B.n738 585
R561 B.n737 B.n52 585
R562 B.n736 B.n735 585
R563 B.n734 B.n53 585
R564 B.n733 B.n732 585
R565 B.n731 B.n730 585
R566 B.n729 B.n57 585
R567 B.n728 B.n727 585
R568 B.n726 B.n58 585
R569 B.n725 B.n724 585
R570 B.n723 B.n59 585
R571 B.n722 B.n721 585
R572 B.n720 B.n60 585
R573 B.n719 B.n718 585
R574 B.n717 B.n61 585
R575 B.n715 B.n714 585
R576 B.n713 B.n64 585
R577 B.n712 B.n711 585
R578 B.n710 B.n65 585
R579 B.n709 B.n708 585
R580 B.n707 B.n66 585
R581 B.n706 B.n705 585
R582 B.n704 B.n67 585
R583 B.n703 B.n702 585
R584 B.n701 B.n68 585
R585 B.n700 B.n699 585
R586 B.n698 B.n69 585
R587 B.n697 B.n696 585
R588 B.n695 B.n70 585
R589 B.n694 B.n693 585
R590 B.n692 B.n71 585
R591 B.n691 B.n690 585
R592 B.n689 B.n72 585
R593 B.n688 B.n687 585
R594 B.n686 B.n73 585
R595 B.n685 B.n684 585
R596 B.n683 B.n74 585
R597 B.n682 B.n681 585
R598 B.n680 B.n75 585
R599 B.n679 B.n678 585
R600 B.n677 B.n76 585
R601 B.n676 B.n675 585
R602 B.n674 B.n77 585
R603 B.n673 B.n672 585
R604 B.n671 B.n78 585
R605 B.n670 B.n669 585
R606 B.n668 B.n79 585
R607 B.n667 B.n666 585
R608 B.n665 B.n80 585
R609 B.n664 B.n663 585
R610 B.n662 B.n81 585
R611 B.n661 B.n660 585
R612 B.n659 B.n82 585
R613 B.n658 B.n657 585
R614 B.n656 B.n83 585
R615 B.n655 B.n654 585
R616 B.n653 B.n84 585
R617 B.n652 B.n651 585
R618 B.n650 B.n85 585
R619 B.n649 B.n648 585
R620 B.n647 B.n86 585
R621 B.n646 B.n645 585
R622 B.n644 B.n87 585
R623 B.n643 B.n642 585
R624 B.n641 B.n88 585
R625 B.n640 B.n639 585
R626 B.n638 B.n89 585
R627 B.n637 B.n636 585
R628 B.n635 B.n90 585
R629 B.n634 B.n633 585
R630 B.n632 B.n91 585
R631 B.n631 B.n630 585
R632 B.n629 B.n92 585
R633 B.n628 B.n627 585
R634 B.n626 B.n93 585
R635 B.n625 B.n624 585
R636 B.n623 B.n94 585
R637 B.n622 B.n621 585
R638 B.n827 B.n22 585
R639 B.n829 B.n828 585
R640 B.n830 B.n21 585
R641 B.n832 B.n831 585
R642 B.n833 B.n20 585
R643 B.n835 B.n834 585
R644 B.n836 B.n19 585
R645 B.n838 B.n837 585
R646 B.n839 B.n18 585
R647 B.n841 B.n840 585
R648 B.n842 B.n17 585
R649 B.n844 B.n843 585
R650 B.n845 B.n16 585
R651 B.n847 B.n846 585
R652 B.n848 B.n15 585
R653 B.n850 B.n849 585
R654 B.n851 B.n14 585
R655 B.n853 B.n852 585
R656 B.n854 B.n13 585
R657 B.n856 B.n855 585
R658 B.n857 B.n12 585
R659 B.n859 B.n858 585
R660 B.n860 B.n11 585
R661 B.n862 B.n861 585
R662 B.n863 B.n10 585
R663 B.n865 B.n864 585
R664 B.n866 B.n9 585
R665 B.n868 B.n867 585
R666 B.n869 B.n8 585
R667 B.n871 B.n870 585
R668 B.n872 B.n7 585
R669 B.n874 B.n873 585
R670 B.n875 B.n6 585
R671 B.n877 B.n876 585
R672 B.n878 B.n5 585
R673 B.n880 B.n879 585
R674 B.n881 B.n4 585
R675 B.n883 B.n882 585
R676 B.n884 B.n3 585
R677 B.n886 B.n885 585
R678 B.n887 B.n0 585
R679 B.n2 B.n1 585
R680 B.n228 B.n227 585
R681 B.n229 B.n226 585
R682 B.n231 B.n230 585
R683 B.n232 B.n225 585
R684 B.n234 B.n233 585
R685 B.n235 B.n224 585
R686 B.n237 B.n236 585
R687 B.n238 B.n223 585
R688 B.n240 B.n239 585
R689 B.n241 B.n222 585
R690 B.n243 B.n242 585
R691 B.n244 B.n221 585
R692 B.n246 B.n245 585
R693 B.n247 B.n220 585
R694 B.n249 B.n248 585
R695 B.n250 B.n219 585
R696 B.n252 B.n251 585
R697 B.n253 B.n218 585
R698 B.n255 B.n254 585
R699 B.n256 B.n217 585
R700 B.n258 B.n257 585
R701 B.n259 B.n216 585
R702 B.n261 B.n260 585
R703 B.n262 B.n215 585
R704 B.n264 B.n263 585
R705 B.n265 B.n214 585
R706 B.n267 B.n266 585
R707 B.n268 B.n213 585
R708 B.n270 B.n269 585
R709 B.n271 B.n212 585
R710 B.n273 B.n272 585
R711 B.n274 B.n211 585
R712 B.n276 B.n275 585
R713 B.n277 B.n210 585
R714 B.n279 B.n278 585
R715 B.n280 B.n209 585
R716 B.n282 B.n281 585
R717 B.n283 B.n208 585
R718 B.n285 B.n284 585
R719 B.n286 B.n207 585
R720 B.n288 B.n207 511.721
R721 B.n496 B.n137 511.721
R722 B.n622 B.n95 511.721
R723 B.n827 B.n826 511.721
R724 B.n174 B.t9 505.053
R725 B.n396 B.t0 505.053
R726 B.n62 B.t3 505.053
R727 B.n54 B.t6 505.053
R728 B.n889 B.n888 256.663
R729 B.n888 B.n887 235.042
R730 B.n888 B.n2 235.042
R731 B.n289 B.n288 163.367
R732 B.n290 B.n289 163.367
R733 B.n290 B.n205 163.367
R734 B.n294 B.n205 163.367
R735 B.n295 B.n294 163.367
R736 B.n296 B.n295 163.367
R737 B.n296 B.n203 163.367
R738 B.n300 B.n203 163.367
R739 B.n301 B.n300 163.367
R740 B.n302 B.n301 163.367
R741 B.n302 B.n201 163.367
R742 B.n306 B.n201 163.367
R743 B.n307 B.n306 163.367
R744 B.n308 B.n307 163.367
R745 B.n308 B.n199 163.367
R746 B.n312 B.n199 163.367
R747 B.n313 B.n312 163.367
R748 B.n314 B.n313 163.367
R749 B.n314 B.n197 163.367
R750 B.n318 B.n197 163.367
R751 B.n319 B.n318 163.367
R752 B.n320 B.n319 163.367
R753 B.n320 B.n195 163.367
R754 B.n324 B.n195 163.367
R755 B.n325 B.n324 163.367
R756 B.n326 B.n325 163.367
R757 B.n326 B.n193 163.367
R758 B.n330 B.n193 163.367
R759 B.n331 B.n330 163.367
R760 B.n332 B.n331 163.367
R761 B.n332 B.n191 163.367
R762 B.n336 B.n191 163.367
R763 B.n337 B.n336 163.367
R764 B.n338 B.n337 163.367
R765 B.n338 B.n189 163.367
R766 B.n342 B.n189 163.367
R767 B.n343 B.n342 163.367
R768 B.n344 B.n343 163.367
R769 B.n344 B.n187 163.367
R770 B.n348 B.n187 163.367
R771 B.n349 B.n348 163.367
R772 B.n350 B.n349 163.367
R773 B.n350 B.n185 163.367
R774 B.n354 B.n185 163.367
R775 B.n355 B.n354 163.367
R776 B.n356 B.n355 163.367
R777 B.n356 B.n183 163.367
R778 B.n360 B.n183 163.367
R779 B.n361 B.n360 163.367
R780 B.n362 B.n361 163.367
R781 B.n362 B.n181 163.367
R782 B.n366 B.n181 163.367
R783 B.n367 B.n366 163.367
R784 B.n368 B.n367 163.367
R785 B.n368 B.n179 163.367
R786 B.n372 B.n179 163.367
R787 B.n373 B.n372 163.367
R788 B.n374 B.n373 163.367
R789 B.n374 B.n177 163.367
R790 B.n378 B.n177 163.367
R791 B.n379 B.n378 163.367
R792 B.n380 B.n379 163.367
R793 B.n380 B.n173 163.367
R794 B.n385 B.n173 163.367
R795 B.n386 B.n385 163.367
R796 B.n387 B.n386 163.367
R797 B.n387 B.n171 163.367
R798 B.n391 B.n171 163.367
R799 B.n392 B.n391 163.367
R800 B.n393 B.n392 163.367
R801 B.n393 B.n169 163.367
R802 B.n400 B.n169 163.367
R803 B.n401 B.n400 163.367
R804 B.n402 B.n401 163.367
R805 B.n402 B.n167 163.367
R806 B.n406 B.n167 163.367
R807 B.n407 B.n406 163.367
R808 B.n408 B.n407 163.367
R809 B.n408 B.n165 163.367
R810 B.n412 B.n165 163.367
R811 B.n413 B.n412 163.367
R812 B.n414 B.n413 163.367
R813 B.n414 B.n163 163.367
R814 B.n418 B.n163 163.367
R815 B.n419 B.n418 163.367
R816 B.n420 B.n419 163.367
R817 B.n420 B.n161 163.367
R818 B.n424 B.n161 163.367
R819 B.n425 B.n424 163.367
R820 B.n426 B.n425 163.367
R821 B.n426 B.n159 163.367
R822 B.n430 B.n159 163.367
R823 B.n431 B.n430 163.367
R824 B.n432 B.n431 163.367
R825 B.n432 B.n157 163.367
R826 B.n436 B.n157 163.367
R827 B.n437 B.n436 163.367
R828 B.n438 B.n437 163.367
R829 B.n438 B.n155 163.367
R830 B.n442 B.n155 163.367
R831 B.n443 B.n442 163.367
R832 B.n444 B.n443 163.367
R833 B.n444 B.n153 163.367
R834 B.n448 B.n153 163.367
R835 B.n449 B.n448 163.367
R836 B.n450 B.n449 163.367
R837 B.n450 B.n151 163.367
R838 B.n454 B.n151 163.367
R839 B.n455 B.n454 163.367
R840 B.n456 B.n455 163.367
R841 B.n456 B.n149 163.367
R842 B.n460 B.n149 163.367
R843 B.n461 B.n460 163.367
R844 B.n462 B.n461 163.367
R845 B.n462 B.n147 163.367
R846 B.n466 B.n147 163.367
R847 B.n467 B.n466 163.367
R848 B.n468 B.n467 163.367
R849 B.n468 B.n145 163.367
R850 B.n472 B.n145 163.367
R851 B.n473 B.n472 163.367
R852 B.n474 B.n473 163.367
R853 B.n474 B.n143 163.367
R854 B.n478 B.n143 163.367
R855 B.n479 B.n478 163.367
R856 B.n480 B.n479 163.367
R857 B.n480 B.n141 163.367
R858 B.n484 B.n141 163.367
R859 B.n485 B.n484 163.367
R860 B.n486 B.n485 163.367
R861 B.n486 B.n139 163.367
R862 B.n490 B.n139 163.367
R863 B.n491 B.n490 163.367
R864 B.n492 B.n491 163.367
R865 B.n492 B.n137 163.367
R866 B.n618 B.n95 163.367
R867 B.n618 B.n617 163.367
R868 B.n617 B.n616 163.367
R869 B.n616 B.n97 163.367
R870 B.n612 B.n97 163.367
R871 B.n612 B.n611 163.367
R872 B.n611 B.n610 163.367
R873 B.n610 B.n99 163.367
R874 B.n606 B.n99 163.367
R875 B.n606 B.n605 163.367
R876 B.n605 B.n604 163.367
R877 B.n604 B.n101 163.367
R878 B.n600 B.n101 163.367
R879 B.n600 B.n599 163.367
R880 B.n599 B.n598 163.367
R881 B.n598 B.n103 163.367
R882 B.n594 B.n103 163.367
R883 B.n594 B.n593 163.367
R884 B.n593 B.n592 163.367
R885 B.n592 B.n105 163.367
R886 B.n588 B.n105 163.367
R887 B.n588 B.n587 163.367
R888 B.n587 B.n586 163.367
R889 B.n586 B.n107 163.367
R890 B.n582 B.n107 163.367
R891 B.n582 B.n581 163.367
R892 B.n581 B.n580 163.367
R893 B.n580 B.n109 163.367
R894 B.n576 B.n109 163.367
R895 B.n576 B.n575 163.367
R896 B.n575 B.n574 163.367
R897 B.n574 B.n111 163.367
R898 B.n570 B.n111 163.367
R899 B.n570 B.n569 163.367
R900 B.n569 B.n568 163.367
R901 B.n568 B.n113 163.367
R902 B.n564 B.n113 163.367
R903 B.n564 B.n563 163.367
R904 B.n563 B.n562 163.367
R905 B.n562 B.n115 163.367
R906 B.n558 B.n115 163.367
R907 B.n558 B.n557 163.367
R908 B.n557 B.n556 163.367
R909 B.n556 B.n117 163.367
R910 B.n552 B.n117 163.367
R911 B.n552 B.n551 163.367
R912 B.n551 B.n550 163.367
R913 B.n550 B.n119 163.367
R914 B.n546 B.n119 163.367
R915 B.n546 B.n545 163.367
R916 B.n545 B.n544 163.367
R917 B.n544 B.n121 163.367
R918 B.n540 B.n121 163.367
R919 B.n540 B.n539 163.367
R920 B.n539 B.n538 163.367
R921 B.n538 B.n123 163.367
R922 B.n534 B.n123 163.367
R923 B.n534 B.n533 163.367
R924 B.n533 B.n532 163.367
R925 B.n532 B.n125 163.367
R926 B.n528 B.n125 163.367
R927 B.n528 B.n527 163.367
R928 B.n527 B.n526 163.367
R929 B.n526 B.n127 163.367
R930 B.n522 B.n127 163.367
R931 B.n522 B.n521 163.367
R932 B.n521 B.n520 163.367
R933 B.n520 B.n129 163.367
R934 B.n516 B.n129 163.367
R935 B.n516 B.n515 163.367
R936 B.n515 B.n514 163.367
R937 B.n514 B.n131 163.367
R938 B.n510 B.n131 163.367
R939 B.n510 B.n509 163.367
R940 B.n509 B.n508 163.367
R941 B.n508 B.n133 163.367
R942 B.n504 B.n133 163.367
R943 B.n504 B.n503 163.367
R944 B.n503 B.n502 163.367
R945 B.n502 B.n135 163.367
R946 B.n498 B.n135 163.367
R947 B.n498 B.n497 163.367
R948 B.n497 B.n496 163.367
R949 B.n826 B.n23 163.367
R950 B.n822 B.n23 163.367
R951 B.n822 B.n821 163.367
R952 B.n821 B.n820 163.367
R953 B.n820 B.n25 163.367
R954 B.n816 B.n25 163.367
R955 B.n816 B.n815 163.367
R956 B.n815 B.n814 163.367
R957 B.n814 B.n27 163.367
R958 B.n810 B.n27 163.367
R959 B.n810 B.n809 163.367
R960 B.n809 B.n808 163.367
R961 B.n808 B.n29 163.367
R962 B.n804 B.n29 163.367
R963 B.n804 B.n803 163.367
R964 B.n803 B.n802 163.367
R965 B.n802 B.n31 163.367
R966 B.n798 B.n31 163.367
R967 B.n798 B.n797 163.367
R968 B.n797 B.n796 163.367
R969 B.n796 B.n33 163.367
R970 B.n792 B.n33 163.367
R971 B.n792 B.n791 163.367
R972 B.n791 B.n790 163.367
R973 B.n790 B.n35 163.367
R974 B.n786 B.n35 163.367
R975 B.n786 B.n785 163.367
R976 B.n785 B.n784 163.367
R977 B.n784 B.n37 163.367
R978 B.n780 B.n37 163.367
R979 B.n780 B.n779 163.367
R980 B.n779 B.n778 163.367
R981 B.n778 B.n39 163.367
R982 B.n774 B.n39 163.367
R983 B.n774 B.n773 163.367
R984 B.n773 B.n772 163.367
R985 B.n772 B.n41 163.367
R986 B.n768 B.n41 163.367
R987 B.n768 B.n767 163.367
R988 B.n767 B.n766 163.367
R989 B.n766 B.n43 163.367
R990 B.n762 B.n43 163.367
R991 B.n762 B.n761 163.367
R992 B.n761 B.n760 163.367
R993 B.n760 B.n45 163.367
R994 B.n756 B.n45 163.367
R995 B.n756 B.n755 163.367
R996 B.n755 B.n754 163.367
R997 B.n754 B.n47 163.367
R998 B.n750 B.n47 163.367
R999 B.n750 B.n749 163.367
R1000 B.n749 B.n748 163.367
R1001 B.n748 B.n49 163.367
R1002 B.n744 B.n49 163.367
R1003 B.n744 B.n743 163.367
R1004 B.n743 B.n742 163.367
R1005 B.n742 B.n51 163.367
R1006 B.n738 B.n51 163.367
R1007 B.n738 B.n737 163.367
R1008 B.n737 B.n736 163.367
R1009 B.n736 B.n53 163.367
R1010 B.n732 B.n53 163.367
R1011 B.n732 B.n731 163.367
R1012 B.n731 B.n57 163.367
R1013 B.n727 B.n57 163.367
R1014 B.n727 B.n726 163.367
R1015 B.n726 B.n725 163.367
R1016 B.n725 B.n59 163.367
R1017 B.n721 B.n59 163.367
R1018 B.n721 B.n720 163.367
R1019 B.n720 B.n719 163.367
R1020 B.n719 B.n61 163.367
R1021 B.n714 B.n61 163.367
R1022 B.n714 B.n713 163.367
R1023 B.n713 B.n712 163.367
R1024 B.n712 B.n65 163.367
R1025 B.n708 B.n65 163.367
R1026 B.n708 B.n707 163.367
R1027 B.n707 B.n706 163.367
R1028 B.n706 B.n67 163.367
R1029 B.n702 B.n67 163.367
R1030 B.n702 B.n701 163.367
R1031 B.n701 B.n700 163.367
R1032 B.n700 B.n69 163.367
R1033 B.n696 B.n69 163.367
R1034 B.n696 B.n695 163.367
R1035 B.n695 B.n694 163.367
R1036 B.n694 B.n71 163.367
R1037 B.n690 B.n71 163.367
R1038 B.n690 B.n689 163.367
R1039 B.n689 B.n688 163.367
R1040 B.n688 B.n73 163.367
R1041 B.n684 B.n73 163.367
R1042 B.n684 B.n683 163.367
R1043 B.n683 B.n682 163.367
R1044 B.n682 B.n75 163.367
R1045 B.n678 B.n75 163.367
R1046 B.n678 B.n677 163.367
R1047 B.n677 B.n676 163.367
R1048 B.n676 B.n77 163.367
R1049 B.n672 B.n77 163.367
R1050 B.n672 B.n671 163.367
R1051 B.n671 B.n670 163.367
R1052 B.n670 B.n79 163.367
R1053 B.n666 B.n79 163.367
R1054 B.n666 B.n665 163.367
R1055 B.n665 B.n664 163.367
R1056 B.n664 B.n81 163.367
R1057 B.n660 B.n81 163.367
R1058 B.n660 B.n659 163.367
R1059 B.n659 B.n658 163.367
R1060 B.n658 B.n83 163.367
R1061 B.n654 B.n83 163.367
R1062 B.n654 B.n653 163.367
R1063 B.n653 B.n652 163.367
R1064 B.n652 B.n85 163.367
R1065 B.n648 B.n85 163.367
R1066 B.n648 B.n647 163.367
R1067 B.n647 B.n646 163.367
R1068 B.n646 B.n87 163.367
R1069 B.n642 B.n87 163.367
R1070 B.n642 B.n641 163.367
R1071 B.n641 B.n640 163.367
R1072 B.n640 B.n89 163.367
R1073 B.n636 B.n89 163.367
R1074 B.n636 B.n635 163.367
R1075 B.n635 B.n634 163.367
R1076 B.n634 B.n91 163.367
R1077 B.n630 B.n91 163.367
R1078 B.n630 B.n629 163.367
R1079 B.n629 B.n628 163.367
R1080 B.n628 B.n93 163.367
R1081 B.n624 B.n93 163.367
R1082 B.n624 B.n623 163.367
R1083 B.n623 B.n622 163.367
R1084 B.n828 B.n827 163.367
R1085 B.n828 B.n21 163.367
R1086 B.n832 B.n21 163.367
R1087 B.n833 B.n832 163.367
R1088 B.n834 B.n833 163.367
R1089 B.n834 B.n19 163.367
R1090 B.n838 B.n19 163.367
R1091 B.n839 B.n838 163.367
R1092 B.n840 B.n839 163.367
R1093 B.n840 B.n17 163.367
R1094 B.n844 B.n17 163.367
R1095 B.n845 B.n844 163.367
R1096 B.n846 B.n845 163.367
R1097 B.n846 B.n15 163.367
R1098 B.n850 B.n15 163.367
R1099 B.n851 B.n850 163.367
R1100 B.n852 B.n851 163.367
R1101 B.n852 B.n13 163.367
R1102 B.n856 B.n13 163.367
R1103 B.n857 B.n856 163.367
R1104 B.n858 B.n857 163.367
R1105 B.n858 B.n11 163.367
R1106 B.n862 B.n11 163.367
R1107 B.n863 B.n862 163.367
R1108 B.n864 B.n863 163.367
R1109 B.n864 B.n9 163.367
R1110 B.n868 B.n9 163.367
R1111 B.n869 B.n868 163.367
R1112 B.n870 B.n869 163.367
R1113 B.n870 B.n7 163.367
R1114 B.n874 B.n7 163.367
R1115 B.n875 B.n874 163.367
R1116 B.n876 B.n875 163.367
R1117 B.n876 B.n5 163.367
R1118 B.n880 B.n5 163.367
R1119 B.n881 B.n880 163.367
R1120 B.n882 B.n881 163.367
R1121 B.n882 B.n3 163.367
R1122 B.n886 B.n3 163.367
R1123 B.n887 B.n886 163.367
R1124 B.n228 B.n2 163.367
R1125 B.n229 B.n228 163.367
R1126 B.n230 B.n229 163.367
R1127 B.n230 B.n225 163.367
R1128 B.n234 B.n225 163.367
R1129 B.n235 B.n234 163.367
R1130 B.n236 B.n235 163.367
R1131 B.n236 B.n223 163.367
R1132 B.n240 B.n223 163.367
R1133 B.n241 B.n240 163.367
R1134 B.n242 B.n241 163.367
R1135 B.n242 B.n221 163.367
R1136 B.n246 B.n221 163.367
R1137 B.n247 B.n246 163.367
R1138 B.n248 B.n247 163.367
R1139 B.n248 B.n219 163.367
R1140 B.n252 B.n219 163.367
R1141 B.n253 B.n252 163.367
R1142 B.n254 B.n253 163.367
R1143 B.n254 B.n217 163.367
R1144 B.n258 B.n217 163.367
R1145 B.n259 B.n258 163.367
R1146 B.n260 B.n259 163.367
R1147 B.n260 B.n215 163.367
R1148 B.n264 B.n215 163.367
R1149 B.n265 B.n264 163.367
R1150 B.n266 B.n265 163.367
R1151 B.n266 B.n213 163.367
R1152 B.n270 B.n213 163.367
R1153 B.n271 B.n270 163.367
R1154 B.n272 B.n271 163.367
R1155 B.n272 B.n211 163.367
R1156 B.n276 B.n211 163.367
R1157 B.n277 B.n276 163.367
R1158 B.n278 B.n277 163.367
R1159 B.n278 B.n209 163.367
R1160 B.n282 B.n209 163.367
R1161 B.n283 B.n282 163.367
R1162 B.n284 B.n283 163.367
R1163 B.n284 B.n207 163.367
R1164 B.n396 B.t1 149.326
R1165 B.n62 B.t5 149.326
R1166 B.n174 B.t10 149.3
R1167 B.n54 B.t8 149.3
R1168 B.n397 B.t2 112.671
R1169 B.n63 B.t4 112.671
R1170 B.n175 B.t11 112.647
R1171 B.n55 B.t7 112.647
R1172 B.n382 B.n175 59.5399
R1173 B.n398 B.n397 59.5399
R1174 B.n716 B.n63 59.5399
R1175 B.n56 B.n55 59.5399
R1176 B.n175 B.n174 36.655
R1177 B.n397 B.n396 36.655
R1178 B.n63 B.n62 36.655
R1179 B.n55 B.n54 36.655
R1180 B.n825 B.n22 33.2493
R1181 B.n621 B.n620 33.2493
R1182 B.n495 B.n494 33.2493
R1183 B.n287 B.n286 33.2493
R1184 B B.n889 18.0485
R1185 B.n829 B.n22 10.6151
R1186 B.n830 B.n829 10.6151
R1187 B.n831 B.n830 10.6151
R1188 B.n831 B.n20 10.6151
R1189 B.n835 B.n20 10.6151
R1190 B.n836 B.n835 10.6151
R1191 B.n837 B.n836 10.6151
R1192 B.n837 B.n18 10.6151
R1193 B.n841 B.n18 10.6151
R1194 B.n842 B.n841 10.6151
R1195 B.n843 B.n842 10.6151
R1196 B.n843 B.n16 10.6151
R1197 B.n847 B.n16 10.6151
R1198 B.n848 B.n847 10.6151
R1199 B.n849 B.n848 10.6151
R1200 B.n849 B.n14 10.6151
R1201 B.n853 B.n14 10.6151
R1202 B.n854 B.n853 10.6151
R1203 B.n855 B.n854 10.6151
R1204 B.n855 B.n12 10.6151
R1205 B.n859 B.n12 10.6151
R1206 B.n860 B.n859 10.6151
R1207 B.n861 B.n860 10.6151
R1208 B.n861 B.n10 10.6151
R1209 B.n865 B.n10 10.6151
R1210 B.n866 B.n865 10.6151
R1211 B.n867 B.n866 10.6151
R1212 B.n867 B.n8 10.6151
R1213 B.n871 B.n8 10.6151
R1214 B.n872 B.n871 10.6151
R1215 B.n873 B.n872 10.6151
R1216 B.n873 B.n6 10.6151
R1217 B.n877 B.n6 10.6151
R1218 B.n878 B.n877 10.6151
R1219 B.n879 B.n878 10.6151
R1220 B.n879 B.n4 10.6151
R1221 B.n883 B.n4 10.6151
R1222 B.n884 B.n883 10.6151
R1223 B.n885 B.n884 10.6151
R1224 B.n885 B.n0 10.6151
R1225 B.n825 B.n824 10.6151
R1226 B.n824 B.n823 10.6151
R1227 B.n823 B.n24 10.6151
R1228 B.n819 B.n24 10.6151
R1229 B.n819 B.n818 10.6151
R1230 B.n818 B.n817 10.6151
R1231 B.n817 B.n26 10.6151
R1232 B.n813 B.n26 10.6151
R1233 B.n813 B.n812 10.6151
R1234 B.n812 B.n811 10.6151
R1235 B.n811 B.n28 10.6151
R1236 B.n807 B.n28 10.6151
R1237 B.n807 B.n806 10.6151
R1238 B.n806 B.n805 10.6151
R1239 B.n805 B.n30 10.6151
R1240 B.n801 B.n30 10.6151
R1241 B.n801 B.n800 10.6151
R1242 B.n800 B.n799 10.6151
R1243 B.n799 B.n32 10.6151
R1244 B.n795 B.n32 10.6151
R1245 B.n795 B.n794 10.6151
R1246 B.n794 B.n793 10.6151
R1247 B.n793 B.n34 10.6151
R1248 B.n789 B.n34 10.6151
R1249 B.n789 B.n788 10.6151
R1250 B.n788 B.n787 10.6151
R1251 B.n787 B.n36 10.6151
R1252 B.n783 B.n36 10.6151
R1253 B.n783 B.n782 10.6151
R1254 B.n782 B.n781 10.6151
R1255 B.n781 B.n38 10.6151
R1256 B.n777 B.n38 10.6151
R1257 B.n777 B.n776 10.6151
R1258 B.n776 B.n775 10.6151
R1259 B.n775 B.n40 10.6151
R1260 B.n771 B.n40 10.6151
R1261 B.n771 B.n770 10.6151
R1262 B.n770 B.n769 10.6151
R1263 B.n769 B.n42 10.6151
R1264 B.n765 B.n42 10.6151
R1265 B.n765 B.n764 10.6151
R1266 B.n764 B.n763 10.6151
R1267 B.n763 B.n44 10.6151
R1268 B.n759 B.n44 10.6151
R1269 B.n759 B.n758 10.6151
R1270 B.n758 B.n757 10.6151
R1271 B.n757 B.n46 10.6151
R1272 B.n753 B.n46 10.6151
R1273 B.n753 B.n752 10.6151
R1274 B.n752 B.n751 10.6151
R1275 B.n751 B.n48 10.6151
R1276 B.n747 B.n48 10.6151
R1277 B.n747 B.n746 10.6151
R1278 B.n746 B.n745 10.6151
R1279 B.n745 B.n50 10.6151
R1280 B.n741 B.n50 10.6151
R1281 B.n741 B.n740 10.6151
R1282 B.n740 B.n739 10.6151
R1283 B.n739 B.n52 10.6151
R1284 B.n735 B.n52 10.6151
R1285 B.n735 B.n734 10.6151
R1286 B.n734 B.n733 10.6151
R1287 B.n730 B.n729 10.6151
R1288 B.n729 B.n728 10.6151
R1289 B.n728 B.n58 10.6151
R1290 B.n724 B.n58 10.6151
R1291 B.n724 B.n723 10.6151
R1292 B.n723 B.n722 10.6151
R1293 B.n722 B.n60 10.6151
R1294 B.n718 B.n60 10.6151
R1295 B.n718 B.n717 10.6151
R1296 B.n715 B.n64 10.6151
R1297 B.n711 B.n64 10.6151
R1298 B.n711 B.n710 10.6151
R1299 B.n710 B.n709 10.6151
R1300 B.n709 B.n66 10.6151
R1301 B.n705 B.n66 10.6151
R1302 B.n705 B.n704 10.6151
R1303 B.n704 B.n703 10.6151
R1304 B.n703 B.n68 10.6151
R1305 B.n699 B.n68 10.6151
R1306 B.n699 B.n698 10.6151
R1307 B.n698 B.n697 10.6151
R1308 B.n697 B.n70 10.6151
R1309 B.n693 B.n70 10.6151
R1310 B.n693 B.n692 10.6151
R1311 B.n692 B.n691 10.6151
R1312 B.n691 B.n72 10.6151
R1313 B.n687 B.n72 10.6151
R1314 B.n687 B.n686 10.6151
R1315 B.n686 B.n685 10.6151
R1316 B.n685 B.n74 10.6151
R1317 B.n681 B.n74 10.6151
R1318 B.n681 B.n680 10.6151
R1319 B.n680 B.n679 10.6151
R1320 B.n679 B.n76 10.6151
R1321 B.n675 B.n76 10.6151
R1322 B.n675 B.n674 10.6151
R1323 B.n674 B.n673 10.6151
R1324 B.n673 B.n78 10.6151
R1325 B.n669 B.n78 10.6151
R1326 B.n669 B.n668 10.6151
R1327 B.n668 B.n667 10.6151
R1328 B.n667 B.n80 10.6151
R1329 B.n663 B.n80 10.6151
R1330 B.n663 B.n662 10.6151
R1331 B.n662 B.n661 10.6151
R1332 B.n661 B.n82 10.6151
R1333 B.n657 B.n82 10.6151
R1334 B.n657 B.n656 10.6151
R1335 B.n656 B.n655 10.6151
R1336 B.n655 B.n84 10.6151
R1337 B.n651 B.n84 10.6151
R1338 B.n651 B.n650 10.6151
R1339 B.n650 B.n649 10.6151
R1340 B.n649 B.n86 10.6151
R1341 B.n645 B.n86 10.6151
R1342 B.n645 B.n644 10.6151
R1343 B.n644 B.n643 10.6151
R1344 B.n643 B.n88 10.6151
R1345 B.n639 B.n88 10.6151
R1346 B.n639 B.n638 10.6151
R1347 B.n638 B.n637 10.6151
R1348 B.n637 B.n90 10.6151
R1349 B.n633 B.n90 10.6151
R1350 B.n633 B.n632 10.6151
R1351 B.n632 B.n631 10.6151
R1352 B.n631 B.n92 10.6151
R1353 B.n627 B.n92 10.6151
R1354 B.n627 B.n626 10.6151
R1355 B.n626 B.n625 10.6151
R1356 B.n625 B.n94 10.6151
R1357 B.n621 B.n94 10.6151
R1358 B.n620 B.n619 10.6151
R1359 B.n619 B.n96 10.6151
R1360 B.n615 B.n96 10.6151
R1361 B.n615 B.n614 10.6151
R1362 B.n614 B.n613 10.6151
R1363 B.n613 B.n98 10.6151
R1364 B.n609 B.n98 10.6151
R1365 B.n609 B.n608 10.6151
R1366 B.n608 B.n607 10.6151
R1367 B.n607 B.n100 10.6151
R1368 B.n603 B.n100 10.6151
R1369 B.n603 B.n602 10.6151
R1370 B.n602 B.n601 10.6151
R1371 B.n601 B.n102 10.6151
R1372 B.n597 B.n102 10.6151
R1373 B.n597 B.n596 10.6151
R1374 B.n596 B.n595 10.6151
R1375 B.n595 B.n104 10.6151
R1376 B.n591 B.n104 10.6151
R1377 B.n591 B.n590 10.6151
R1378 B.n590 B.n589 10.6151
R1379 B.n589 B.n106 10.6151
R1380 B.n585 B.n106 10.6151
R1381 B.n585 B.n584 10.6151
R1382 B.n584 B.n583 10.6151
R1383 B.n583 B.n108 10.6151
R1384 B.n579 B.n108 10.6151
R1385 B.n579 B.n578 10.6151
R1386 B.n578 B.n577 10.6151
R1387 B.n577 B.n110 10.6151
R1388 B.n573 B.n110 10.6151
R1389 B.n573 B.n572 10.6151
R1390 B.n572 B.n571 10.6151
R1391 B.n571 B.n112 10.6151
R1392 B.n567 B.n112 10.6151
R1393 B.n567 B.n566 10.6151
R1394 B.n566 B.n565 10.6151
R1395 B.n565 B.n114 10.6151
R1396 B.n561 B.n114 10.6151
R1397 B.n561 B.n560 10.6151
R1398 B.n560 B.n559 10.6151
R1399 B.n559 B.n116 10.6151
R1400 B.n555 B.n116 10.6151
R1401 B.n555 B.n554 10.6151
R1402 B.n554 B.n553 10.6151
R1403 B.n553 B.n118 10.6151
R1404 B.n549 B.n118 10.6151
R1405 B.n549 B.n548 10.6151
R1406 B.n548 B.n547 10.6151
R1407 B.n547 B.n120 10.6151
R1408 B.n543 B.n120 10.6151
R1409 B.n543 B.n542 10.6151
R1410 B.n542 B.n541 10.6151
R1411 B.n541 B.n122 10.6151
R1412 B.n537 B.n122 10.6151
R1413 B.n537 B.n536 10.6151
R1414 B.n536 B.n535 10.6151
R1415 B.n535 B.n124 10.6151
R1416 B.n531 B.n124 10.6151
R1417 B.n531 B.n530 10.6151
R1418 B.n530 B.n529 10.6151
R1419 B.n529 B.n126 10.6151
R1420 B.n525 B.n126 10.6151
R1421 B.n525 B.n524 10.6151
R1422 B.n524 B.n523 10.6151
R1423 B.n523 B.n128 10.6151
R1424 B.n519 B.n128 10.6151
R1425 B.n519 B.n518 10.6151
R1426 B.n518 B.n517 10.6151
R1427 B.n517 B.n130 10.6151
R1428 B.n513 B.n130 10.6151
R1429 B.n513 B.n512 10.6151
R1430 B.n512 B.n511 10.6151
R1431 B.n511 B.n132 10.6151
R1432 B.n507 B.n132 10.6151
R1433 B.n507 B.n506 10.6151
R1434 B.n506 B.n505 10.6151
R1435 B.n505 B.n134 10.6151
R1436 B.n501 B.n134 10.6151
R1437 B.n501 B.n500 10.6151
R1438 B.n500 B.n499 10.6151
R1439 B.n499 B.n136 10.6151
R1440 B.n495 B.n136 10.6151
R1441 B.n227 B.n1 10.6151
R1442 B.n227 B.n226 10.6151
R1443 B.n231 B.n226 10.6151
R1444 B.n232 B.n231 10.6151
R1445 B.n233 B.n232 10.6151
R1446 B.n233 B.n224 10.6151
R1447 B.n237 B.n224 10.6151
R1448 B.n238 B.n237 10.6151
R1449 B.n239 B.n238 10.6151
R1450 B.n239 B.n222 10.6151
R1451 B.n243 B.n222 10.6151
R1452 B.n244 B.n243 10.6151
R1453 B.n245 B.n244 10.6151
R1454 B.n245 B.n220 10.6151
R1455 B.n249 B.n220 10.6151
R1456 B.n250 B.n249 10.6151
R1457 B.n251 B.n250 10.6151
R1458 B.n251 B.n218 10.6151
R1459 B.n255 B.n218 10.6151
R1460 B.n256 B.n255 10.6151
R1461 B.n257 B.n256 10.6151
R1462 B.n257 B.n216 10.6151
R1463 B.n261 B.n216 10.6151
R1464 B.n262 B.n261 10.6151
R1465 B.n263 B.n262 10.6151
R1466 B.n263 B.n214 10.6151
R1467 B.n267 B.n214 10.6151
R1468 B.n268 B.n267 10.6151
R1469 B.n269 B.n268 10.6151
R1470 B.n269 B.n212 10.6151
R1471 B.n273 B.n212 10.6151
R1472 B.n274 B.n273 10.6151
R1473 B.n275 B.n274 10.6151
R1474 B.n275 B.n210 10.6151
R1475 B.n279 B.n210 10.6151
R1476 B.n280 B.n279 10.6151
R1477 B.n281 B.n280 10.6151
R1478 B.n281 B.n208 10.6151
R1479 B.n285 B.n208 10.6151
R1480 B.n286 B.n285 10.6151
R1481 B.n287 B.n206 10.6151
R1482 B.n291 B.n206 10.6151
R1483 B.n292 B.n291 10.6151
R1484 B.n293 B.n292 10.6151
R1485 B.n293 B.n204 10.6151
R1486 B.n297 B.n204 10.6151
R1487 B.n298 B.n297 10.6151
R1488 B.n299 B.n298 10.6151
R1489 B.n299 B.n202 10.6151
R1490 B.n303 B.n202 10.6151
R1491 B.n304 B.n303 10.6151
R1492 B.n305 B.n304 10.6151
R1493 B.n305 B.n200 10.6151
R1494 B.n309 B.n200 10.6151
R1495 B.n310 B.n309 10.6151
R1496 B.n311 B.n310 10.6151
R1497 B.n311 B.n198 10.6151
R1498 B.n315 B.n198 10.6151
R1499 B.n316 B.n315 10.6151
R1500 B.n317 B.n316 10.6151
R1501 B.n317 B.n196 10.6151
R1502 B.n321 B.n196 10.6151
R1503 B.n322 B.n321 10.6151
R1504 B.n323 B.n322 10.6151
R1505 B.n323 B.n194 10.6151
R1506 B.n327 B.n194 10.6151
R1507 B.n328 B.n327 10.6151
R1508 B.n329 B.n328 10.6151
R1509 B.n329 B.n192 10.6151
R1510 B.n333 B.n192 10.6151
R1511 B.n334 B.n333 10.6151
R1512 B.n335 B.n334 10.6151
R1513 B.n335 B.n190 10.6151
R1514 B.n339 B.n190 10.6151
R1515 B.n340 B.n339 10.6151
R1516 B.n341 B.n340 10.6151
R1517 B.n341 B.n188 10.6151
R1518 B.n345 B.n188 10.6151
R1519 B.n346 B.n345 10.6151
R1520 B.n347 B.n346 10.6151
R1521 B.n347 B.n186 10.6151
R1522 B.n351 B.n186 10.6151
R1523 B.n352 B.n351 10.6151
R1524 B.n353 B.n352 10.6151
R1525 B.n353 B.n184 10.6151
R1526 B.n357 B.n184 10.6151
R1527 B.n358 B.n357 10.6151
R1528 B.n359 B.n358 10.6151
R1529 B.n359 B.n182 10.6151
R1530 B.n363 B.n182 10.6151
R1531 B.n364 B.n363 10.6151
R1532 B.n365 B.n364 10.6151
R1533 B.n365 B.n180 10.6151
R1534 B.n369 B.n180 10.6151
R1535 B.n370 B.n369 10.6151
R1536 B.n371 B.n370 10.6151
R1537 B.n371 B.n178 10.6151
R1538 B.n375 B.n178 10.6151
R1539 B.n376 B.n375 10.6151
R1540 B.n377 B.n376 10.6151
R1541 B.n377 B.n176 10.6151
R1542 B.n381 B.n176 10.6151
R1543 B.n384 B.n383 10.6151
R1544 B.n384 B.n172 10.6151
R1545 B.n388 B.n172 10.6151
R1546 B.n389 B.n388 10.6151
R1547 B.n390 B.n389 10.6151
R1548 B.n390 B.n170 10.6151
R1549 B.n394 B.n170 10.6151
R1550 B.n395 B.n394 10.6151
R1551 B.n399 B.n395 10.6151
R1552 B.n403 B.n168 10.6151
R1553 B.n404 B.n403 10.6151
R1554 B.n405 B.n404 10.6151
R1555 B.n405 B.n166 10.6151
R1556 B.n409 B.n166 10.6151
R1557 B.n410 B.n409 10.6151
R1558 B.n411 B.n410 10.6151
R1559 B.n411 B.n164 10.6151
R1560 B.n415 B.n164 10.6151
R1561 B.n416 B.n415 10.6151
R1562 B.n417 B.n416 10.6151
R1563 B.n417 B.n162 10.6151
R1564 B.n421 B.n162 10.6151
R1565 B.n422 B.n421 10.6151
R1566 B.n423 B.n422 10.6151
R1567 B.n423 B.n160 10.6151
R1568 B.n427 B.n160 10.6151
R1569 B.n428 B.n427 10.6151
R1570 B.n429 B.n428 10.6151
R1571 B.n429 B.n158 10.6151
R1572 B.n433 B.n158 10.6151
R1573 B.n434 B.n433 10.6151
R1574 B.n435 B.n434 10.6151
R1575 B.n435 B.n156 10.6151
R1576 B.n439 B.n156 10.6151
R1577 B.n440 B.n439 10.6151
R1578 B.n441 B.n440 10.6151
R1579 B.n441 B.n154 10.6151
R1580 B.n445 B.n154 10.6151
R1581 B.n446 B.n445 10.6151
R1582 B.n447 B.n446 10.6151
R1583 B.n447 B.n152 10.6151
R1584 B.n451 B.n152 10.6151
R1585 B.n452 B.n451 10.6151
R1586 B.n453 B.n452 10.6151
R1587 B.n453 B.n150 10.6151
R1588 B.n457 B.n150 10.6151
R1589 B.n458 B.n457 10.6151
R1590 B.n459 B.n458 10.6151
R1591 B.n459 B.n148 10.6151
R1592 B.n463 B.n148 10.6151
R1593 B.n464 B.n463 10.6151
R1594 B.n465 B.n464 10.6151
R1595 B.n465 B.n146 10.6151
R1596 B.n469 B.n146 10.6151
R1597 B.n470 B.n469 10.6151
R1598 B.n471 B.n470 10.6151
R1599 B.n471 B.n144 10.6151
R1600 B.n475 B.n144 10.6151
R1601 B.n476 B.n475 10.6151
R1602 B.n477 B.n476 10.6151
R1603 B.n477 B.n142 10.6151
R1604 B.n481 B.n142 10.6151
R1605 B.n482 B.n481 10.6151
R1606 B.n483 B.n482 10.6151
R1607 B.n483 B.n140 10.6151
R1608 B.n487 B.n140 10.6151
R1609 B.n488 B.n487 10.6151
R1610 B.n489 B.n488 10.6151
R1611 B.n489 B.n138 10.6151
R1612 B.n493 B.n138 10.6151
R1613 B.n494 B.n493 10.6151
R1614 B.n733 B.n56 9.36635
R1615 B.n716 B.n715 9.36635
R1616 B.n382 B.n381 9.36635
R1617 B.n398 B.n168 9.36635
R1618 B.n889 B.n0 8.11757
R1619 B.n889 B.n1 8.11757
R1620 B.n730 B.n56 1.24928
R1621 B.n717 B.n716 1.24928
R1622 B.n383 B.n382 1.24928
R1623 B.n399 B.n398 1.24928
C0 VDD2 B 2.70726f
C1 VP VDD1 15.138599f
C2 VN VP 8.23139f
C3 VDD2 VDD1 1.49945f
C4 VN VDD2 14.8436f
C5 VTAIL w_n3238_n4844# 4.16276f
C6 VTAIL B 4.74989f
C7 B w_n3238_n4844# 10.8667f
C8 VP VDD2 0.452152f
C9 VTAIL VDD1 15.304999f
C10 VN VTAIL 14.750999f
C11 VDD1 w_n3238_n4844# 2.91729f
C12 VN w_n3238_n4844# 6.74932f
C13 B VDD1 2.62985f
C14 VN B 1.10827f
C15 VTAIL VP 14.7655f
C16 VP w_n3238_n4844# 7.16768f
C17 VTAIL VDD2 15.3448f
C18 VN VDD1 0.151306f
C19 VDD2 w_n3238_n4844# 3.00687f
C20 VP B 1.80603f
C21 VDD2 VSUBS 1.977315f
C22 VDD1 VSUBS 1.746972f
C23 VTAIL VSUBS 1.2917f
C24 VN VSUBS 6.42998f
C25 VP VSUBS 3.171281f
C26 B VSUBS 4.70025f
C27 w_n3238_n4844# VSUBS 0.191599p
C28 B.n0 VSUBS 0.007055f
C29 B.n1 VSUBS 0.007055f
C30 B.n2 VSUBS 0.010434f
C31 B.n3 VSUBS 0.007996f
C32 B.n4 VSUBS 0.007996f
C33 B.n5 VSUBS 0.007996f
C34 B.n6 VSUBS 0.007996f
C35 B.n7 VSUBS 0.007996f
C36 B.n8 VSUBS 0.007996f
C37 B.n9 VSUBS 0.007996f
C38 B.n10 VSUBS 0.007996f
C39 B.n11 VSUBS 0.007996f
C40 B.n12 VSUBS 0.007996f
C41 B.n13 VSUBS 0.007996f
C42 B.n14 VSUBS 0.007996f
C43 B.n15 VSUBS 0.007996f
C44 B.n16 VSUBS 0.007996f
C45 B.n17 VSUBS 0.007996f
C46 B.n18 VSUBS 0.007996f
C47 B.n19 VSUBS 0.007996f
C48 B.n20 VSUBS 0.007996f
C49 B.n21 VSUBS 0.007996f
C50 B.n22 VSUBS 0.018603f
C51 B.n23 VSUBS 0.007996f
C52 B.n24 VSUBS 0.007996f
C53 B.n25 VSUBS 0.007996f
C54 B.n26 VSUBS 0.007996f
C55 B.n27 VSUBS 0.007996f
C56 B.n28 VSUBS 0.007996f
C57 B.n29 VSUBS 0.007996f
C58 B.n30 VSUBS 0.007996f
C59 B.n31 VSUBS 0.007996f
C60 B.n32 VSUBS 0.007996f
C61 B.n33 VSUBS 0.007996f
C62 B.n34 VSUBS 0.007996f
C63 B.n35 VSUBS 0.007996f
C64 B.n36 VSUBS 0.007996f
C65 B.n37 VSUBS 0.007996f
C66 B.n38 VSUBS 0.007996f
C67 B.n39 VSUBS 0.007996f
C68 B.n40 VSUBS 0.007996f
C69 B.n41 VSUBS 0.007996f
C70 B.n42 VSUBS 0.007996f
C71 B.n43 VSUBS 0.007996f
C72 B.n44 VSUBS 0.007996f
C73 B.n45 VSUBS 0.007996f
C74 B.n46 VSUBS 0.007996f
C75 B.n47 VSUBS 0.007996f
C76 B.n48 VSUBS 0.007996f
C77 B.n49 VSUBS 0.007996f
C78 B.n50 VSUBS 0.007996f
C79 B.n51 VSUBS 0.007996f
C80 B.n52 VSUBS 0.007996f
C81 B.n53 VSUBS 0.007996f
C82 B.t7 VSUBS 0.751099f
C83 B.t8 VSUBS 0.767321f
C84 B.t6 VSUBS 1.46562f
C85 B.n54 VSUBS 0.342517f
C86 B.n55 VSUBS 0.077481f
C87 B.n56 VSUBS 0.018526f
C88 B.n57 VSUBS 0.007996f
C89 B.n58 VSUBS 0.007996f
C90 B.n59 VSUBS 0.007996f
C91 B.n60 VSUBS 0.007996f
C92 B.n61 VSUBS 0.007996f
C93 B.t4 VSUBS 0.751069f
C94 B.t5 VSUBS 0.767296f
C95 B.t3 VSUBS 1.46562f
C96 B.n62 VSUBS 0.342542f
C97 B.n63 VSUBS 0.07751f
C98 B.n64 VSUBS 0.007996f
C99 B.n65 VSUBS 0.007996f
C100 B.n66 VSUBS 0.007996f
C101 B.n67 VSUBS 0.007996f
C102 B.n68 VSUBS 0.007996f
C103 B.n69 VSUBS 0.007996f
C104 B.n70 VSUBS 0.007996f
C105 B.n71 VSUBS 0.007996f
C106 B.n72 VSUBS 0.007996f
C107 B.n73 VSUBS 0.007996f
C108 B.n74 VSUBS 0.007996f
C109 B.n75 VSUBS 0.007996f
C110 B.n76 VSUBS 0.007996f
C111 B.n77 VSUBS 0.007996f
C112 B.n78 VSUBS 0.007996f
C113 B.n79 VSUBS 0.007996f
C114 B.n80 VSUBS 0.007996f
C115 B.n81 VSUBS 0.007996f
C116 B.n82 VSUBS 0.007996f
C117 B.n83 VSUBS 0.007996f
C118 B.n84 VSUBS 0.007996f
C119 B.n85 VSUBS 0.007996f
C120 B.n86 VSUBS 0.007996f
C121 B.n87 VSUBS 0.007996f
C122 B.n88 VSUBS 0.007996f
C123 B.n89 VSUBS 0.007996f
C124 B.n90 VSUBS 0.007996f
C125 B.n91 VSUBS 0.007996f
C126 B.n92 VSUBS 0.007996f
C127 B.n93 VSUBS 0.007996f
C128 B.n94 VSUBS 0.007996f
C129 B.n95 VSUBS 0.018603f
C130 B.n96 VSUBS 0.007996f
C131 B.n97 VSUBS 0.007996f
C132 B.n98 VSUBS 0.007996f
C133 B.n99 VSUBS 0.007996f
C134 B.n100 VSUBS 0.007996f
C135 B.n101 VSUBS 0.007996f
C136 B.n102 VSUBS 0.007996f
C137 B.n103 VSUBS 0.007996f
C138 B.n104 VSUBS 0.007996f
C139 B.n105 VSUBS 0.007996f
C140 B.n106 VSUBS 0.007996f
C141 B.n107 VSUBS 0.007996f
C142 B.n108 VSUBS 0.007996f
C143 B.n109 VSUBS 0.007996f
C144 B.n110 VSUBS 0.007996f
C145 B.n111 VSUBS 0.007996f
C146 B.n112 VSUBS 0.007996f
C147 B.n113 VSUBS 0.007996f
C148 B.n114 VSUBS 0.007996f
C149 B.n115 VSUBS 0.007996f
C150 B.n116 VSUBS 0.007996f
C151 B.n117 VSUBS 0.007996f
C152 B.n118 VSUBS 0.007996f
C153 B.n119 VSUBS 0.007996f
C154 B.n120 VSUBS 0.007996f
C155 B.n121 VSUBS 0.007996f
C156 B.n122 VSUBS 0.007996f
C157 B.n123 VSUBS 0.007996f
C158 B.n124 VSUBS 0.007996f
C159 B.n125 VSUBS 0.007996f
C160 B.n126 VSUBS 0.007996f
C161 B.n127 VSUBS 0.007996f
C162 B.n128 VSUBS 0.007996f
C163 B.n129 VSUBS 0.007996f
C164 B.n130 VSUBS 0.007996f
C165 B.n131 VSUBS 0.007996f
C166 B.n132 VSUBS 0.007996f
C167 B.n133 VSUBS 0.007996f
C168 B.n134 VSUBS 0.007996f
C169 B.n135 VSUBS 0.007996f
C170 B.n136 VSUBS 0.007996f
C171 B.n137 VSUBS 0.01926f
C172 B.n138 VSUBS 0.007996f
C173 B.n139 VSUBS 0.007996f
C174 B.n140 VSUBS 0.007996f
C175 B.n141 VSUBS 0.007996f
C176 B.n142 VSUBS 0.007996f
C177 B.n143 VSUBS 0.007996f
C178 B.n144 VSUBS 0.007996f
C179 B.n145 VSUBS 0.007996f
C180 B.n146 VSUBS 0.007996f
C181 B.n147 VSUBS 0.007996f
C182 B.n148 VSUBS 0.007996f
C183 B.n149 VSUBS 0.007996f
C184 B.n150 VSUBS 0.007996f
C185 B.n151 VSUBS 0.007996f
C186 B.n152 VSUBS 0.007996f
C187 B.n153 VSUBS 0.007996f
C188 B.n154 VSUBS 0.007996f
C189 B.n155 VSUBS 0.007996f
C190 B.n156 VSUBS 0.007996f
C191 B.n157 VSUBS 0.007996f
C192 B.n158 VSUBS 0.007996f
C193 B.n159 VSUBS 0.007996f
C194 B.n160 VSUBS 0.007996f
C195 B.n161 VSUBS 0.007996f
C196 B.n162 VSUBS 0.007996f
C197 B.n163 VSUBS 0.007996f
C198 B.n164 VSUBS 0.007996f
C199 B.n165 VSUBS 0.007996f
C200 B.n166 VSUBS 0.007996f
C201 B.n167 VSUBS 0.007996f
C202 B.n168 VSUBS 0.007526f
C203 B.n169 VSUBS 0.007996f
C204 B.n170 VSUBS 0.007996f
C205 B.n171 VSUBS 0.007996f
C206 B.n172 VSUBS 0.007996f
C207 B.n173 VSUBS 0.007996f
C208 B.t11 VSUBS 0.751099f
C209 B.t10 VSUBS 0.767321f
C210 B.t9 VSUBS 1.46562f
C211 B.n174 VSUBS 0.342517f
C212 B.n175 VSUBS 0.077481f
C213 B.n176 VSUBS 0.007996f
C214 B.n177 VSUBS 0.007996f
C215 B.n178 VSUBS 0.007996f
C216 B.n179 VSUBS 0.007996f
C217 B.n180 VSUBS 0.007996f
C218 B.n181 VSUBS 0.007996f
C219 B.n182 VSUBS 0.007996f
C220 B.n183 VSUBS 0.007996f
C221 B.n184 VSUBS 0.007996f
C222 B.n185 VSUBS 0.007996f
C223 B.n186 VSUBS 0.007996f
C224 B.n187 VSUBS 0.007996f
C225 B.n188 VSUBS 0.007996f
C226 B.n189 VSUBS 0.007996f
C227 B.n190 VSUBS 0.007996f
C228 B.n191 VSUBS 0.007996f
C229 B.n192 VSUBS 0.007996f
C230 B.n193 VSUBS 0.007996f
C231 B.n194 VSUBS 0.007996f
C232 B.n195 VSUBS 0.007996f
C233 B.n196 VSUBS 0.007996f
C234 B.n197 VSUBS 0.007996f
C235 B.n198 VSUBS 0.007996f
C236 B.n199 VSUBS 0.007996f
C237 B.n200 VSUBS 0.007996f
C238 B.n201 VSUBS 0.007996f
C239 B.n202 VSUBS 0.007996f
C240 B.n203 VSUBS 0.007996f
C241 B.n204 VSUBS 0.007996f
C242 B.n205 VSUBS 0.007996f
C243 B.n206 VSUBS 0.007996f
C244 B.n207 VSUBS 0.018603f
C245 B.n208 VSUBS 0.007996f
C246 B.n209 VSUBS 0.007996f
C247 B.n210 VSUBS 0.007996f
C248 B.n211 VSUBS 0.007996f
C249 B.n212 VSUBS 0.007996f
C250 B.n213 VSUBS 0.007996f
C251 B.n214 VSUBS 0.007996f
C252 B.n215 VSUBS 0.007996f
C253 B.n216 VSUBS 0.007996f
C254 B.n217 VSUBS 0.007996f
C255 B.n218 VSUBS 0.007996f
C256 B.n219 VSUBS 0.007996f
C257 B.n220 VSUBS 0.007996f
C258 B.n221 VSUBS 0.007996f
C259 B.n222 VSUBS 0.007996f
C260 B.n223 VSUBS 0.007996f
C261 B.n224 VSUBS 0.007996f
C262 B.n225 VSUBS 0.007996f
C263 B.n226 VSUBS 0.007996f
C264 B.n227 VSUBS 0.007996f
C265 B.n228 VSUBS 0.007996f
C266 B.n229 VSUBS 0.007996f
C267 B.n230 VSUBS 0.007996f
C268 B.n231 VSUBS 0.007996f
C269 B.n232 VSUBS 0.007996f
C270 B.n233 VSUBS 0.007996f
C271 B.n234 VSUBS 0.007996f
C272 B.n235 VSUBS 0.007996f
C273 B.n236 VSUBS 0.007996f
C274 B.n237 VSUBS 0.007996f
C275 B.n238 VSUBS 0.007996f
C276 B.n239 VSUBS 0.007996f
C277 B.n240 VSUBS 0.007996f
C278 B.n241 VSUBS 0.007996f
C279 B.n242 VSUBS 0.007996f
C280 B.n243 VSUBS 0.007996f
C281 B.n244 VSUBS 0.007996f
C282 B.n245 VSUBS 0.007996f
C283 B.n246 VSUBS 0.007996f
C284 B.n247 VSUBS 0.007996f
C285 B.n248 VSUBS 0.007996f
C286 B.n249 VSUBS 0.007996f
C287 B.n250 VSUBS 0.007996f
C288 B.n251 VSUBS 0.007996f
C289 B.n252 VSUBS 0.007996f
C290 B.n253 VSUBS 0.007996f
C291 B.n254 VSUBS 0.007996f
C292 B.n255 VSUBS 0.007996f
C293 B.n256 VSUBS 0.007996f
C294 B.n257 VSUBS 0.007996f
C295 B.n258 VSUBS 0.007996f
C296 B.n259 VSUBS 0.007996f
C297 B.n260 VSUBS 0.007996f
C298 B.n261 VSUBS 0.007996f
C299 B.n262 VSUBS 0.007996f
C300 B.n263 VSUBS 0.007996f
C301 B.n264 VSUBS 0.007996f
C302 B.n265 VSUBS 0.007996f
C303 B.n266 VSUBS 0.007996f
C304 B.n267 VSUBS 0.007996f
C305 B.n268 VSUBS 0.007996f
C306 B.n269 VSUBS 0.007996f
C307 B.n270 VSUBS 0.007996f
C308 B.n271 VSUBS 0.007996f
C309 B.n272 VSUBS 0.007996f
C310 B.n273 VSUBS 0.007996f
C311 B.n274 VSUBS 0.007996f
C312 B.n275 VSUBS 0.007996f
C313 B.n276 VSUBS 0.007996f
C314 B.n277 VSUBS 0.007996f
C315 B.n278 VSUBS 0.007996f
C316 B.n279 VSUBS 0.007996f
C317 B.n280 VSUBS 0.007996f
C318 B.n281 VSUBS 0.007996f
C319 B.n282 VSUBS 0.007996f
C320 B.n283 VSUBS 0.007996f
C321 B.n284 VSUBS 0.007996f
C322 B.n285 VSUBS 0.007996f
C323 B.n286 VSUBS 0.018603f
C324 B.n287 VSUBS 0.01926f
C325 B.n288 VSUBS 0.01926f
C326 B.n289 VSUBS 0.007996f
C327 B.n290 VSUBS 0.007996f
C328 B.n291 VSUBS 0.007996f
C329 B.n292 VSUBS 0.007996f
C330 B.n293 VSUBS 0.007996f
C331 B.n294 VSUBS 0.007996f
C332 B.n295 VSUBS 0.007996f
C333 B.n296 VSUBS 0.007996f
C334 B.n297 VSUBS 0.007996f
C335 B.n298 VSUBS 0.007996f
C336 B.n299 VSUBS 0.007996f
C337 B.n300 VSUBS 0.007996f
C338 B.n301 VSUBS 0.007996f
C339 B.n302 VSUBS 0.007996f
C340 B.n303 VSUBS 0.007996f
C341 B.n304 VSUBS 0.007996f
C342 B.n305 VSUBS 0.007996f
C343 B.n306 VSUBS 0.007996f
C344 B.n307 VSUBS 0.007996f
C345 B.n308 VSUBS 0.007996f
C346 B.n309 VSUBS 0.007996f
C347 B.n310 VSUBS 0.007996f
C348 B.n311 VSUBS 0.007996f
C349 B.n312 VSUBS 0.007996f
C350 B.n313 VSUBS 0.007996f
C351 B.n314 VSUBS 0.007996f
C352 B.n315 VSUBS 0.007996f
C353 B.n316 VSUBS 0.007996f
C354 B.n317 VSUBS 0.007996f
C355 B.n318 VSUBS 0.007996f
C356 B.n319 VSUBS 0.007996f
C357 B.n320 VSUBS 0.007996f
C358 B.n321 VSUBS 0.007996f
C359 B.n322 VSUBS 0.007996f
C360 B.n323 VSUBS 0.007996f
C361 B.n324 VSUBS 0.007996f
C362 B.n325 VSUBS 0.007996f
C363 B.n326 VSUBS 0.007996f
C364 B.n327 VSUBS 0.007996f
C365 B.n328 VSUBS 0.007996f
C366 B.n329 VSUBS 0.007996f
C367 B.n330 VSUBS 0.007996f
C368 B.n331 VSUBS 0.007996f
C369 B.n332 VSUBS 0.007996f
C370 B.n333 VSUBS 0.007996f
C371 B.n334 VSUBS 0.007996f
C372 B.n335 VSUBS 0.007996f
C373 B.n336 VSUBS 0.007996f
C374 B.n337 VSUBS 0.007996f
C375 B.n338 VSUBS 0.007996f
C376 B.n339 VSUBS 0.007996f
C377 B.n340 VSUBS 0.007996f
C378 B.n341 VSUBS 0.007996f
C379 B.n342 VSUBS 0.007996f
C380 B.n343 VSUBS 0.007996f
C381 B.n344 VSUBS 0.007996f
C382 B.n345 VSUBS 0.007996f
C383 B.n346 VSUBS 0.007996f
C384 B.n347 VSUBS 0.007996f
C385 B.n348 VSUBS 0.007996f
C386 B.n349 VSUBS 0.007996f
C387 B.n350 VSUBS 0.007996f
C388 B.n351 VSUBS 0.007996f
C389 B.n352 VSUBS 0.007996f
C390 B.n353 VSUBS 0.007996f
C391 B.n354 VSUBS 0.007996f
C392 B.n355 VSUBS 0.007996f
C393 B.n356 VSUBS 0.007996f
C394 B.n357 VSUBS 0.007996f
C395 B.n358 VSUBS 0.007996f
C396 B.n359 VSUBS 0.007996f
C397 B.n360 VSUBS 0.007996f
C398 B.n361 VSUBS 0.007996f
C399 B.n362 VSUBS 0.007996f
C400 B.n363 VSUBS 0.007996f
C401 B.n364 VSUBS 0.007996f
C402 B.n365 VSUBS 0.007996f
C403 B.n366 VSUBS 0.007996f
C404 B.n367 VSUBS 0.007996f
C405 B.n368 VSUBS 0.007996f
C406 B.n369 VSUBS 0.007996f
C407 B.n370 VSUBS 0.007996f
C408 B.n371 VSUBS 0.007996f
C409 B.n372 VSUBS 0.007996f
C410 B.n373 VSUBS 0.007996f
C411 B.n374 VSUBS 0.007996f
C412 B.n375 VSUBS 0.007996f
C413 B.n376 VSUBS 0.007996f
C414 B.n377 VSUBS 0.007996f
C415 B.n378 VSUBS 0.007996f
C416 B.n379 VSUBS 0.007996f
C417 B.n380 VSUBS 0.007996f
C418 B.n381 VSUBS 0.007526f
C419 B.n382 VSUBS 0.018526f
C420 B.n383 VSUBS 0.004468f
C421 B.n384 VSUBS 0.007996f
C422 B.n385 VSUBS 0.007996f
C423 B.n386 VSUBS 0.007996f
C424 B.n387 VSUBS 0.007996f
C425 B.n388 VSUBS 0.007996f
C426 B.n389 VSUBS 0.007996f
C427 B.n390 VSUBS 0.007996f
C428 B.n391 VSUBS 0.007996f
C429 B.n392 VSUBS 0.007996f
C430 B.n393 VSUBS 0.007996f
C431 B.n394 VSUBS 0.007996f
C432 B.n395 VSUBS 0.007996f
C433 B.t2 VSUBS 0.751069f
C434 B.t1 VSUBS 0.767296f
C435 B.t0 VSUBS 1.46562f
C436 B.n396 VSUBS 0.342542f
C437 B.n397 VSUBS 0.07751f
C438 B.n398 VSUBS 0.018526f
C439 B.n399 VSUBS 0.004468f
C440 B.n400 VSUBS 0.007996f
C441 B.n401 VSUBS 0.007996f
C442 B.n402 VSUBS 0.007996f
C443 B.n403 VSUBS 0.007996f
C444 B.n404 VSUBS 0.007996f
C445 B.n405 VSUBS 0.007996f
C446 B.n406 VSUBS 0.007996f
C447 B.n407 VSUBS 0.007996f
C448 B.n408 VSUBS 0.007996f
C449 B.n409 VSUBS 0.007996f
C450 B.n410 VSUBS 0.007996f
C451 B.n411 VSUBS 0.007996f
C452 B.n412 VSUBS 0.007996f
C453 B.n413 VSUBS 0.007996f
C454 B.n414 VSUBS 0.007996f
C455 B.n415 VSUBS 0.007996f
C456 B.n416 VSUBS 0.007996f
C457 B.n417 VSUBS 0.007996f
C458 B.n418 VSUBS 0.007996f
C459 B.n419 VSUBS 0.007996f
C460 B.n420 VSUBS 0.007996f
C461 B.n421 VSUBS 0.007996f
C462 B.n422 VSUBS 0.007996f
C463 B.n423 VSUBS 0.007996f
C464 B.n424 VSUBS 0.007996f
C465 B.n425 VSUBS 0.007996f
C466 B.n426 VSUBS 0.007996f
C467 B.n427 VSUBS 0.007996f
C468 B.n428 VSUBS 0.007996f
C469 B.n429 VSUBS 0.007996f
C470 B.n430 VSUBS 0.007996f
C471 B.n431 VSUBS 0.007996f
C472 B.n432 VSUBS 0.007996f
C473 B.n433 VSUBS 0.007996f
C474 B.n434 VSUBS 0.007996f
C475 B.n435 VSUBS 0.007996f
C476 B.n436 VSUBS 0.007996f
C477 B.n437 VSUBS 0.007996f
C478 B.n438 VSUBS 0.007996f
C479 B.n439 VSUBS 0.007996f
C480 B.n440 VSUBS 0.007996f
C481 B.n441 VSUBS 0.007996f
C482 B.n442 VSUBS 0.007996f
C483 B.n443 VSUBS 0.007996f
C484 B.n444 VSUBS 0.007996f
C485 B.n445 VSUBS 0.007996f
C486 B.n446 VSUBS 0.007996f
C487 B.n447 VSUBS 0.007996f
C488 B.n448 VSUBS 0.007996f
C489 B.n449 VSUBS 0.007996f
C490 B.n450 VSUBS 0.007996f
C491 B.n451 VSUBS 0.007996f
C492 B.n452 VSUBS 0.007996f
C493 B.n453 VSUBS 0.007996f
C494 B.n454 VSUBS 0.007996f
C495 B.n455 VSUBS 0.007996f
C496 B.n456 VSUBS 0.007996f
C497 B.n457 VSUBS 0.007996f
C498 B.n458 VSUBS 0.007996f
C499 B.n459 VSUBS 0.007996f
C500 B.n460 VSUBS 0.007996f
C501 B.n461 VSUBS 0.007996f
C502 B.n462 VSUBS 0.007996f
C503 B.n463 VSUBS 0.007996f
C504 B.n464 VSUBS 0.007996f
C505 B.n465 VSUBS 0.007996f
C506 B.n466 VSUBS 0.007996f
C507 B.n467 VSUBS 0.007996f
C508 B.n468 VSUBS 0.007996f
C509 B.n469 VSUBS 0.007996f
C510 B.n470 VSUBS 0.007996f
C511 B.n471 VSUBS 0.007996f
C512 B.n472 VSUBS 0.007996f
C513 B.n473 VSUBS 0.007996f
C514 B.n474 VSUBS 0.007996f
C515 B.n475 VSUBS 0.007996f
C516 B.n476 VSUBS 0.007996f
C517 B.n477 VSUBS 0.007996f
C518 B.n478 VSUBS 0.007996f
C519 B.n479 VSUBS 0.007996f
C520 B.n480 VSUBS 0.007996f
C521 B.n481 VSUBS 0.007996f
C522 B.n482 VSUBS 0.007996f
C523 B.n483 VSUBS 0.007996f
C524 B.n484 VSUBS 0.007996f
C525 B.n485 VSUBS 0.007996f
C526 B.n486 VSUBS 0.007996f
C527 B.n487 VSUBS 0.007996f
C528 B.n488 VSUBS 0.007996f
C529 B.n489 VSUBS 0.007996f
C530 B.n490 VSUBS 0.007996f
C531 B.n491 VSUBS 0.007996f
C532 B.n492 VSUBS 0.007996f
C533 B.n493 VSUBS 0.007996f
C534 B.n494 VSUBS 0.018332f
C535 B.n495 VSUBS 0.019531f
C536 B.n496 VSUBS 0.018603f
C537 B.n497 VSUBS 0.007996f
C538 B.n498 VSUBS 0.007996f
C539 B.n499 VSUBS 0.007996f
C540 B.n500 VSUBS 0.007996f
C541 B.n501 VSUBS 0.007996f
C542 B.n502 VSUBS 0.007996f
C543 B.n503 VSUBS 0.007996f
C544 B.n504 VSUBS 0.007996f
C545 B.n505 VSUBS 0.007996f
C546 B.n506 VSUBS 0.007996f
C547 B.n507 VSUBS 0.007996f
C548 B.n508 VSUBS 0.007996f
C549 B.n509 VSUBS 0.007996f
C550 B.n510 VSUBS 0.007996f
C551 B.n511 VSUBS 0.007996f
C552 B.n512 VSUBS 0.007996f
C553 B.n513 VSUBS 0.007996f
C554 B.n514 VSUBS 0.007996f
C555 B.n515 VSUBS 0.007996f
C556 B.n516 VSUBS 0.007996f
C557 B.n517 VSUBS 0.007996f
C558 B.n518 VSUBS 0.007996f
C559 B.n519 VSUBS 0.007996f
C560 B.n520 VSUBS 0.007996f
C561 B.n521 VSUBS 0.007996f
C562 B.n522 VSUBS 0.007996f
C563 B.n523 VSUBS 0.007996f
C564 B.n524 VSUBS 0.007996f
C565 B.n525 VSUBS 0.007996f
C566 B.n526 VSUBS 0.007996f
C567 B.n527 VSUBS 0.007996f
C568 B.n528 VSUBS 0.007996f
C569 B.n529 VSUBS 0.007996f
C570 B.n530 VSUBS 0.007996f
C571 B.n531 VSUBS 0.007996f
C572 B.n532 VSUBS 0.007996f
C573 B.n533 VSUBS 0.007996f
C574 B.n534 VSUBS 0.007996f
C575 B.n535 VSUBS 0.007996f
C576 B.n536 VSUBS 0.007996f
C577 B.n537 VSUBS 0.007996f
C578 B.n538 VSUBS 0.007996f
C579 B.n539 VSUBS 0.007996f
C580 B.n540 VSUBS 0.007996f
C581 B.n541 VSUBS 0.007996f
C582 B.n542 VSUBS 0.007996f
C583 B.n543 VSUBS 0.007996f
C584 B.n544 VSUBS 0.007996f
C585 B.n545 VSUBS 0.007996f
C586 B.n546 VSUBS 0.007996f
C587 B.n547 VSUBS 0.007996f
C588 B.n548 VSUBS 0.007996f
C589 B.n549 VSUBS 0.007996f
C590 B.n550 VSUBS 0.007996f
C591 B.n551 VSUBS 0.007996f
C592 B.n552 VSUBS 0.007996f
C593 B.n553 VSUBS 0.007996f
C594 B.n554 VSUBS 0.007996f
C595 B.n555 VSUBS 0.007996f
C596 B.n556 VSUBS 0.007996f
C597 B.n557 VSUBS 0.007996f
C598 B.n558 VSUBS 0.007996f
C599 B.n559 VSUBS 0.007996f
C600 B.n560 VSUBS 0.007996f
C601 B.n561 VSUBS 0.007996f
C602 B.n562 VSUBS 0.007996f
C603 B.n563 VSUBS 0.007996f
C604 B.n564 VSUBS 0.007996f
C605 B.n565 VSUBS 0.007996f
C606 B.n566 VSUBS 0.007996f
C607 B.n567 VSUBS 0.007996f
C608 B.n568 VSUBS 0.007996f
C609 B.n569 VSUBS 0.007996f
C610 B.n570 VSUBS 0.007996f
C611 B.n571 VSUBS 0.007996f
C612 B.n572 VSUBS 0.007996f
C613 B.n573 VSUBS 0.007996f
C614 B.n574 VSUBS 0.007996f
C615 B.n575 VSUBS 0.007996f
C616 B.n576 VSUBS 0.007996f
C617 B.n577 VSUBS 0.007996f
C618 B.n578 VSUBS 0.007996f
C619 B.n579 VSUBS 0.007996f
C620 B.n580 VSUBS 0.007996f
C621 B.n581 VSUBS 0.007996f
C622 B.n582 VSUBS 0.007996f
C623 B.n583 VSUBS 0.007996f
C624 B.n584 VSUBS 0.007996f
C625 B.n585 VSUBS 0.007996f
C626 B.n586 VSUBS 0.007996f
C627 B.n587 VSUBS 0.007996f
C628 B.n588 VSUBS 0.007996f
C629 B.n589 VSUBS 0.007996f
C630 B.n590 VSUBS 0.007996f
C631 B.n591 VSUBS 0.007996f
C632 B.n592 VSUBS 0.007996f
C633 B.n593 VSUBS 0.007996f
C634 B.n594 VSUBS 0.007996f
C635 B.n595 VSUBS 0.007996f
C636 B.n596 VSUBS 0.007996f
C637 B.n597 VSUBS 0.007996f
C638 B.n598 VSUBS 0.007996f
C639 B.n599 VSUBS 0.007996f
C640 B.n600 VSUBS 0.007996f
C641 B.n601 VSUBS 0.007996f
C642 B.n602 VSUBS 0.007996f
C643 B.n603 VSUBS 0.007996f
C644 B.n604 VSUBS 0.007996f
C645 B.n605 VSUBS 0.007996f
C646 B.n606 VSUBS 0.007996f
C647 B.n607 VSUBS 0.007996f
C648 B.n608 VSUBS 0.007996f
C649 B.n609 VSUBS 0.007996f
C650 B.n610 VSUBS 0.007996f
C651 B.n611 VSUBS 0.007996f
C652 B.n612 VSUBS 0.007996f
C653 B.n613 VSUBS 0.007996f
C654 B.n614 VSUBS 0.007996f
C655 B.n615 VSUBS 0.007996f
C656 B.n616 VSUBS 0.007996f
C657 B.n617 VSUBS 0.007996f
C658 B.n618 VSUBS 0.007996f
C659 B.n619 VSUBS 0.007996f
C660 B.n620 VSUBS 0.018603f
C661 B.n621 VSUBS 0.01926f
C662 B.n622 VSUBS 0.01926f
C663 B.n623 VSUBS 0.007996f
C664 B.n624 VSUBS 0.007996f
C665 B.n625 VSUBS 0.007996f
C666 B.n626 VSUBS 0.007996f
C667 B.n627 VSUBS 0.007996f
C668 B.n628 VSUBS 0.007996f
C669 B.n629 VSUBS 0.007996f
C670 B.n630 VSUBS 0.007996f
C671 B.n631 VSUBS 0.007996f
C672 B.n632 VSUBS 0.007996f
C673 B.n633 VSUBS 0.007996f
C674 B.n634 VSUBS 0.007996f
C675 B.n635 VSUBS 0.007996f
C676 B.n636 VSUBS 0.007996f
C677 B.n637 VSUBS 0.007996f
C678 B.n638 VSUBS 0.007996f
C679 B.n639 VSUBS 0.007996f
C680 B.n640 VSUBS 0.007996f
C681 B.n641 VSUBS 0.007996f
C682 B.n642 VSUBS 0.007996f
C683 B.n643 VSUBS 0.007996f
C684 B.n644 VSUBS 0.007996f
C685 B.n645 VSUBS 0.007996f
C686 B.n646 VSUBS 0.007996f
C687 B.n647 VSUBS 0.007996f
C688 B.n648 VSUBS 0.007996f
C689 B.n649 VSUBS 0.007996f
C690 B.n650 VSUBS 0.007996f
C691 B.n651 VSUBS 0.007996f
C692 B.n652 VSUBS 0.007996f
C693 B.n653 VSUBS 0.007996f
C694 B.n654 VSUBS 0.007996f
C695 B.n655 VSUBS 0.007996f
C696 B.n656 VSUBS 0.007996f
C697 B.n657 VSUBS 0.007996f
C698 B.n658 VSUBS 0.007996f
C699 B.n659 VSUBS 0.007996f
C700 B.n660 VSUBS 0.007996f
C701 B.n661 VSUBS 0.007996f
C702 B.n662 VSUBS 0.007996f
C703 B.n663 VSUBS 0.007996f
C704 B.n664 VSUBS 0.007996f
C705 B.n665 VSUBS 0.007996f
C706 B.n666 VSUBS 0.007996f
C707 B.n667 VSUBS 0.007996f
C708 B.n668 VSUBS 0.007996f
C709 B.n669 VSUBS 0.007996f
C710 B.n670 VSUBS 0.007996f
C711 B.n671 VSUBS 0.007996f
C712 B.n672 VSUBS 0.007996f
C713 B.n673 VSUBS 0.007996f
C714 B.n674 VSUBS 0.007996f
C715 B.n675 VSUBS 0.007996f
C716 B.n676 VSUBS 0.007996f
C717 B.n677 VSUBS 0.007996f
C718 B.n678 VSUBS 0.007996f
C719 B.n679 VSUBS 0.007996f
C720 B.n680 VSUBS 0.007996f
C721 B.n681 VSUBS 0.007996f
C722 B.n682 VSUBS 0.007996f
C723 B.n683 VSUBS 0.007996f
C724 B.n684 VSUBS 0.007996f
C725 B.n685 VSUBS 0.007996f
C726 B.n686 VSUBS 0.007996f
C727 B.n687 VSUBS 0.007996f
C728 B.n688 VSUBS 0.007996f
C729 B.n689 VSUBS 0.007996f
C730 B.n690 VSUBS 0.007996f
C731 B.n691 VSUBS 0.007996f
C732 B.n692 VSUBS 0.007996f
C733 B.n693 VSUBS 0.007996f
C734 B.n694 VSUBS 0.007996f
C735 B.n695 VSUBS 0.007996f
C736 B.n696 VSUBS 0.007996f
C737 B.n697 VSUBS 0.007996f
C738 B.n698 VSUBS 0.007996f
C739 B.n699 VSUBS 0.007996f
C740 B.n700 VSUBS 0.007996f
C741 B.n701 VSUBS 0.007996f
C742 B.n702 VSUBS 0.007996f
C743 B.n703 VSUBS 0.007996f
C744 B.n704 VSUBS 0.007996f
C745 B.n705 VSUBS 0.007996f
C746 B.n706 VSUBS 0.007996f
C747 B.n707 VSUBS 0.007996f
C748 B.n708 VSUBS 0.007996f
C749 B.n709 VSUBS 0.007996f
C750 B.n710 VSUBS 0.007996f
C751 B.n711 VSUBS 0.007996f
C752 B.n712 VSUBS 0.007996f
C753 B.n713 VSUBS 0.007996f
C754 B.n714 VSUBS 0.007996f
C755 B.n715 VSUBS 0.007526f
C756 B.n716 VSUBS 0.018526f
C757 B.n717 VSUBS 0.004468f
C758 B.n718 VSUBS 0.007996f
C759 B.n719 VSUBS 0.007996f
C760 B.n720 VSUBS 0.007996f
C761 B.n721 VSUBS 0.007996f
C762 B.n722 VSUBS 0.007996f
C763 B.n723 VSUBS 0.007996f
C764 B.n724 VSUBS 0.007996f
C765 B.n725 VSUBS 0.007996f
C766 B.n726 VSUBS 0.007996f
C767 B.n727 VSUBS 0.007996f
C768 B.n728 VSUBS 0.007996f
C769 B.n729 VSUBS 0.007996f
C770 B.n730 VSUBS 0.004468f
C771 B.n731 VSUBS 0.007996f
C772 B.n732 VSUBS 0.007996f
C773 B.n733 VSUBS 0.007526f
C774 B.n734 VSUBS 0.007996f
C775 B.n735 VSUBS 0.007996f
C776 B.n736 VSUBS 0.007996f
C777 B.n737 VSUBS 0.007996f
C778 B.n738 VSUBS 0.007996f
C779 B.n739 VSUBS 0.007996f
C780 B.n740 VSUBS 0.007996f
C781 B.n741 VSUBS 0.007996f
C782 B.n742 VSUBS 0.007996f
C783 B.n743 VSUBS 0.007996f
C784 B.n744 VSUBS 0.007996f
C785 B.n745 VSUBS 0.007996f
C786 B.n746 VSUBS 0.007996f
C787 B.n747 VSUBS 0.007996f
C788 B.n748 VSUBS 0.007996f
C789 B.n749 VSUBS 0.007996f
C790 B.n750 VSUBS 0.007996f
C791 B.n751 VSUBS 0.007996f
C792 B.n752 VSUBS 0.007996f
C793 B.n753 VSUBS 0.007996f
C794 B.n754 VSUBS 0.007996f
C795 B.n755 VSUBS 0.007996f
C796 B.n756 VSUBS 0.007996f
C797 B.n757 VSUBS 0.007996f
C798 B.n758 VSUBS 0.007996f
C799 B.n759 VSUBS 0.007996f
C800 B.n760 VSUBS 0.007996f
C801 B.n761 VSUBS 0.007996f
C802 B.n762 VSUBS 0.007996f
C803 B.n763 VSUBS 0.007996f
C804 B.n764 VSUBS 0.007996f
C805 B.n765 VSUBS 0.007996f
C806 B.n766 VSUBS 0.007996f
C807 B.n767 VSUBS 0.007996f
C808 B.n768 VSUBS 0.007996f
C809 B.n769 VSUBS 0.007996f
C810 B.n770 VSUBS 0.007996f
C811 B.n771 VSUBS 0.007996f
C812 B.n772 VSUBS 0.007996f
C813 B.n773 VSUBS 0.007996f
C814 B.n774 VSUBS 0.007996f
C815 B.n775 VSUBS 0.007996f
C816 B.n776 VSUBS 0.007996f
C817 B.n777 VSUBS 0.007996f
C818 B.n778 VSUBS 0.007996f
C819 B.n779 VSUBS 0.007996f
C820 B.n780 VSUBS 0.007996f
C821 B.n781 VSUBS 0.007996f
C822 B.n782 VSUBS 0.007996f
C823 B.n783 VSUBS 0.007996f
C824 B.n784 VSUBS 0.007996f
C825 B.n785 VSUBS 0.007996f
C826 B.n786 VSUBS 0.007996f
C827 B.n787 VSUBS 0.007996f
C828 B.n788 VSUBS 0.007996f
C829 B.n789 VSUBS 0.007996f
C830 B.n790 VSUBS 0.007996f
C831 B.n791 VSUBS 0.007996f
C832 B.n792 VSUBS 0.007996f
C833 B.n793 VSUBS 0.007996f
C834 B.n794 VSUBS 0.007996f
C835 B.n795 VSUBS 0.007996f
C836 B.n796 VSUBS 0.007996f
C837 B.n797 VSUBS 0.007996f
C838 B.n798 VSUBS 0.007996f
C839 B.n799 VSUBS 0.007996f
C840 B.n800 VSUBS 0.007996f
C841 B.n801 VSUBS 0.007996f
C842 B.n802 VSUBS 0.007996f
C843 B.n803 VSUBS 0.007996f
C844 B.n804 VSUBS 0.007996f
C845 B.n805 VSUBS 0.007996f
C846 B.n806 VSUBS 0.007996f
C847 B.n807 VSUBS 0.007996f
C848 B.n808 VSUBS 0.007996f
C849 B.n809 VSUBS 0.007996f
C850 B.n810 VSUBS 0.007996f
C851 B.n811 VSUBS 0.007996f
C852 B.n812 VSUBS 0.007996f
C853 B.n813 VSUBS 0.007996f
C854 B.n814 VSUBS 0.007996f
C855 B.n815 VSUBS 0.007996f
C856 B.n816 VSUBS 0.007996f
C857 B.n817 VSUBS 0.007996f
C858 B.n818 VSUBS 0.007996f
C859 B.n819 VSUBS 0.007996f
C860 B.n820 VSUBS 0.007996f
C861 B.n821 VSUBS 0.007996f
C862 B.n822 VSUBS 0.007996f
C863 B.n823 VSUBS 0.007996f
C864 B.n824 VSUBS 0.007996f
C865 B.n825 VSUBS 0.01926f
C866 B.n826 VSUBS 0.01926f
C867 B.n827 VSUBS 0.018603f
C868 B.n828 VSUBS 0.007996f
C869 B.n829 VSUBS 0.007996f
C870 B.n830 VSUBS 0.007996f
C871 B.n831 VSUBS 0.007996f
C872 B.n832 VSUBS 0.007996f
C873 B.n833 VSUBS 0.007996f
C874 B.n834 VSUBS 0.007996f
C875 B.n835 VSUBS 0.007996f
C876 B.n836 VSUBS 0.007996f
C877 B.n837 VSUBS 0.007996f
C878 B.n838 VSUBS 0.007996f
C879 B.n839 VSUBS 0.007996f
C880 B.n840 VSUBS 0.007996f
C881 B.n841 VSUBS 0.007996f
C882 B.n842 VSUBS 0.007996f
C883 B.n843 VSUBS 0.007996f
C884 B.n844 VSUBS 0.007996f
C885 B.n845 VSUBS 0.007996f
C886 B.n846 VSUBS 0.007996f
C887 B.n847 VSUBS 0.007996f
C888 B.n848 VSUBS 0.007996f
C889 B.n849 VSUBS 0.007996f
C890 B.n850 VSUBS 0.007996f
C891 B.n851 VSUBS 0.007996f
C892 B.n852 VSUBS 0.007996f
C893 B.n853 VSUBS 0.007996f
C894 B.n854 VSUBS 0.007996f
C895 B.n855 VSUBS 0.007996f
C896 B.n856 VSUBS 0.007996f
C897 B.n857 VSUBS 0.007996f
C898 B.n858 VSUBS 0.007996f
C899 B.n859 VSUBS 0.007996f
C900 B.n860 VSUBS 0.007996f
C901 B.n861 VSUBS 0.007996f
C902 B.n862 VSUBS 0.007996f
C903 B.n863 VSUBS 0.007996f
C904 B.n864 VSUBS 0.007996f
C905 B.n865 VSUBS 0.007996f
C906 B.n866 VSUBS 0.007996f
C907 B.n867 VSUBS 0.007996f
C908 B.n868 VSUBS 0.007996f
C909 B.n869 VSUBS 0.007996f
C910 B.n870 VSUBS 0.007996f
C911 B.n871 VSUBS 0.007996f
C912 B.n872 VSUBS 0.007996f
C913 B.n873 VSUBS 0.007996f
C914 B.n874 VSUBS 0.007996f
C915 B.n875 VSUBS 0.007996f
C916 B.n876 VSUBS 0.007996f
C917 B.n877 VSUBS 0.007996f
C918 B.n878 VSUBS 0.007996f
C919 B.n879 VSUBS 0.007996f
C920 B.n880 VSUBS 0.007996f
C921 B.n881 VSUBS 0.007996f
C922 B.n882 VSUBS 0.007996f
C923 B.n883 VSUBS 0.007996f
C924 B.n884 VSUBS 0.007996f
C925 B.n885 VSUBS 0.007996f
C926 B.n886 VSUBS 0.007996f
C927 B.n887 VSUBS 0.010434f
C928 B.n888 VSUBS 0.011115f
C929 B.n889 VSUBS 0.022104f
C930 VDD2.t1 VSUBS 4.42097f
C931 VDD2.t5 VSUBS 0.404753f
C932 VDD2.t6 VSUBS 0.404753f
C933 VDD2.n0 VSUBS 3.39653f
C934 VDD2.n1 VSUBS 1.4433f
C935 VDD2.t0 VSUBS 0.404753f
C936 VDD2.t4 VSUBS 0.404753f
C937 VDD2.n2 VSUBS 3.40928f
C938 VDD2.n3 VSUBS 3.28165f
C939 VDD2.t8 VSUBS 4.40377f
C940 VDD2.n4 VSUBS 3.80376f
C941 VDD2.t7 VSUBS 0.404753f
C942 VDD2.t9 VSUBS 0.404753f
C943 VDD2.n5 VSUBS 3.39653f
C944 VDD2.n6 VSUBS 0.700395f
C945 VDD2.t3 VSUBS 0.404753f
C946 VDD2.t2 VSUBS 0.404753f
C947 VDD2.n7 VSUBS 3.40923f
C948 VN.n0 VSUBS 0.033442f
C949 VN.t5 VSUBS 2.7847f
C950 VN.n1 VSUBS 0.030222f
C951 VN.n2 VSUBS 0.033442f
C952 VN.t9 VSUBS 2.7847f
C953 VN.n3 VSUBS 0.043524f
C954 VN.n4 VSUBS 0.033442f
C955 VN.t3 VSUBS 2.7847f
C956 VN.n5 VSUBS 0.053702f
C957 VN.t8 VSUBS 2.88095f
C958 VN.n6 VSUBS 1.06668f
C959 VN.t4 VSUBS 2.7847f
C960 VN.n7 VSUBS 1.03355f
C961 VN.n8 VSUBS 0.039972f
C962 VN.n9 VSUBS 0.208268f
C963 VN.n10 VSUBS 0.033442f
C964 VN.n11 VSUBS 0.033442f
C965 VN.n12 VSUBS 0.043524f
C966 VN.n13 VSUBS 0.046708f
C967 VN.n14 VSUBS 0.975094f
C968 VN.n15 VSUBS 0.046708f
C969 VN.n16 VSUBS 0.033442f
C970 VN.n17 VSUBS 0.033442f
C971 VN.n18 VSUBS 0.033442f
C972 VN.n19 VSUBS 0.053702f
C973 VN.n20 VSUBS 0.039972f
C974 VN.n21 VSUBS 0.975094f
C975 VN.n22 VSUBS 0.058432f
C976 VN.n23 VSUBS 0.033442f
C977 VN.n24 VSUBS 0.033442f
C978 VN.n25 VSUBS 0.033442f
C979 VN.n26 VSUBS 0.062015f
C980 VN.n27 VSUBS 0.033237f
C981 VN.n28 VSUBS 1.03416f
C982 VN.n29 VSUBS 0.034381f
C983 VN.n30 VSUBS 0.033442f
C984 VN.t1 VSUBS 2.7847f
C985 VN.n31 VSUBS 0.030222f
C986 VN.n32 VSUBS 0.033442f
C987 VN.t2 VSUBS 2.7847f
C988 VN.n33 VSUBS 0.043524f
C989 VN.n34 VSUBS 0.033442f
C990 VN.t0 VSUBS 2.7847f
C991 VN.n35 VSUBS 0.053702f
C992 VN.t7 VSUBS 2.88095f
C993 VN.n36 VSUBS 1.06668f
C994 VN.t6 VSUBS 2.7847f
C995 VN.n37 VSUBS 1.03355f
C996 VN.n38 VSUBS 0.039972f
C997 VN.n39 VSUBS 0.208268f
C998 VN.n40 VSUBS 0.033442f
C999 VN.n41 VSUBS 0.033442f
C1000 VN.n42 VSUBS 0.043524f
C1001 VN.n43 VSUBS 0.046708f
C1002 VN.n44 VSUBS 0.975094f
C1003 VN.n45 VSUBS 0.046708f
C1004 VN.n46 VSUBS 0.033442f
C1005 VN.n47 VSUBS 0.033442f
C1006 VN.n48 VSUBS 0.033442f
C1007 VN.n49 VSUBS 0.053702f
C1008 VN.n50 VSUBS 0.039972f
C1009 VN.n51 VSUBS 0.975094f
C1010 VN.n52 VSUBS 0.058432f
C1011 VN.n53 VSUBS 0.033442f
C1012 VN.n54 VSUBS 0.033442f
C1013 VN.n55 VSUBS 0.033442f
C1014 VN.n56 VSUBS 0.062015f
C1015 VN.n57 VSUBS 0.033237f
C1016 VN.n58 VSUBS 1.03416f
C1017 VN.n59 VSUBS 2.0046f
C1018 VDD1.t1 VSUBS 4.42127f
C1019 VDD1.t2 VSUBS 0.404779f
C1020 VDD1.t3 VSUBS 0.404779f
C1021 VDD1.n0 VSUBS 3.39676f
C1022 VDD1.n1 VSUBS 1.45132f
C1023 VDD1.t9 VSUBS 4.421259f
C1024 VDD1.t5 VSUBS 0.404779f
C1025 VDD1.t0 VSUBS 0.404779f
C1026 VDD1.n2 VSUBS 3.39676f
C1027 VDD1.n3 VSUBS 1.44339f
C1028 VDD1.t6 VSUBS 0.404779f
C1029 VDD1.t4 VSUBS 0.404779f
C1030 VDD1.n4 VSUBS 3.40951f
C1031 VDD1.n5 VSUBS 3.38874f
C1032 VDD1.t7 VSUBS 0.404779f
C1033 VDD1.t8 VSUBS 0.404779f
C1034 VDD1.n6 VSUBS 3.39674f
C1035 VDD1.n7 VSUBS 3.79725f
C1036 VTAIL.t6 VSUBS 0.410696f
C1037 VTAIL.t7 VSUBS 0.410696f
C1038 VTAIL.n0 VSUBS 3.28048f
C1039 VTAIL.n1 VSUBS 0.880753f
C1040 VTAIL.t18 VSUBS 4.27755f
C1041 VTAIL.n2 VSUBS 1.03393f
C1042 VTAIL.t11 VSUBS 0.410696f
C1043 VTAIL.t17 VSUBS 0.410696f
C1044 VTAIL.n3 VSUBS 3.28048f
C1045 VTAIL.n4 VSUBS 0.940719f
C1046 VTAIL.t10 VSUBS 0.410696f
C1047 VTAIL.t14 VSUBS 0.410696f
C1048 VTAIL.n5 VSUBS 3.28048f
C1049 VTAIL.n6 VSUBS 2.88945f
C1050 VTAIL.t5 VSUBS 0.410696f
C1051 VTAIL.t2 VSUBS 0.410696f
C1052 VTAIL.n7 VSUBS 3.28048f
C1053 VTAIL.n8 VSUBS 2.88945f
C1054 VTAIL.t8 VSUBS 0.410696f
C1055 VTAIL.t3 VSUBS 0.410696f
C1056 VTAIL.n9 VSUBS 3.28048f
C1057 VTAIL.n10 VSUBS 0.94072f
C1058 VTAIL.t4 VSUBS 4.27756f
C1059 VTAIL.n11 VSUBS 1.03392f
C1060 VTAIL.t19 VSUBS 0.410696f
C1061 VTAIL.t16 VSUBS 0.410696f
C1062 VTAIL.n12 VSUBS 3.28048f
C1063 VTAIL.n13 VSUBS 0.910923f
C1064 VTAIL.t12 VSUBS 0.410696f
C1065 VTAIL.t15 VSUBS 0.410696f
C1066 VTAIL.n14 VSUBS 3.28048f
C1067 VTAIL.n15 VSUBS 0.94072f
C1068 VTAIL.t13 VSUBS 4.27755f
C1069 VTAIL.n16 VSUBS 2.87167f
C1070 VTAIL.t0 VSUBS 4.27755f
C1071 VTAIL.n17 VSUBS 2.87167f
C1072 VTAIL.t9 VSUBS 0.410696f
C1073 VTAIL.t1 VSUBS 0.410696f
C1074 VTAIL.n18 VSUBS 3.28048f
C1075 VTAIL.n19 VSUBS 0.830098f
C1076 VP.n0 VSUBS 0.034079f
C1077 VP.t5 VSUBS 2.83776f
C1078 VP.n1 VSUBS 0.030798f
C1079 VP.n2 VSUBS 0.034079f
C1080 VP.t3 VSUBS 2.83776f
C1081 VP.n3 VSUBS 0.044354f
C1082 VP.n4 VSUBS 0.034079f
C1083 VP.t9 VSUBS 2.83776f
C1084 VP.n5 VSUBS 0.054725f
C1085 VP.n6 VSUBS 0.034079f
C1086 VP.t4 VSUBS 2.83776f
C1087 VP.n7 VSUBS 0.063197f
C1088 VP.n8 VSUBS 0.034079f
C1089 VP.t1 VSUBS 2.83776f
C1090 VP.n9 VSUBS 0.030798f
C1091 VP.n10 VSUBS 0.034079f
C1092 VP.t2 VSUBS 2.83776f
C1093 VP.n11 VSUBS 0.044354f
C1094 VP.n12 VSUBS 0.034079f
C1095 VP.t6 VSUBS 2.83776f
C1096 VP.n13 VSUBS 0.054725f
C1097 VP.t8 VSUBS 2.93584f
C1098 VP.n14 VSUBS 1.087f
C1099 VP.t7 VSUBS 2.83776f
C1100 VP.n15 VSUBS 1.05324f
C1101 VP.n16 VSUBS 0.040734f
C1102 VP.n17 VSUBS 0.212237f
C1103 VP.n18 VSUBS 0.034079f
C1104 VP.n19 VSUBS 0.034079f
C1105 VP.n20 VSUBS 0.044354f
C1106 VP.n21 VSUBS 0.047598f
C1107 VP.n22 VSUBS 0.993673f
C1108 VP.n23 VSUBS 0.047598f
C1109 VP.n24 VSUBS 0.034079f
C1110 VP.n25 VSUBS 0.034079f
C1111 VP.n26 VSUBS 0.034079f
C1112 VP.n27 VSUBS 0.054725f
C1113 VP.n28 VSUBS 0.040734f
C1114 VP.n29 VSUBS 0.993673f
C1115 VP.n30 VSUBS 0.059545f
C1116 VP.n31 VSUBS 0.034079f
C1117 VP.n32 VSUBS 0.034079f
C1118 VP.n33 VSUBS 0.034079f
C1119 VP.n34 VSUBS 0.063197f
C1120 VP.n35 VSUBS 0.03387f
C1121 VP.n36 VSUBS 1.05386f
C1122 VP.n37 VSUBS 2.0207f
C1123 VP.n38 VSUBS 2.04394f
C1124 VP.t0 VSUBS 2.83776f
C1125 VP.n39 VSUBS 1.05386f
C1126 VP.n40 VSUBS 0.03387f
C1127 VP.n41 VSUBS 0.034079f
C1128 VP.n42 VSUBS 0.034079f
C1129 VP.n43 VSUBS 0.034079f
C1130 VP.n44 VSUBS 0.030798f
C1131 VP.n45 VSUBS 0.059545f
C1132 VP.n46 VSUBS 0.993673f
C1133 VP.n47 VSUBS 0.040734f
C1134 VP.n48 VSUBS 0.034079f
C1135 VP.n49 VSUBS 0.034079f
C1136 VP.n50 VSUBS 0.034079f
C1137 VP.n51 VSUBS 0.044354f
C1138 VP.n52 VSUBS 0.047598f
C1139 VP.n53 VSUBS 0.993673f
C1140 VP.n54 VSUBS 0.047598f
C1141 VP.n55 VSUBS 0.034079f
C1142 VP.n56 VSUBS 0.034079f
C1143 VP.n57 VSUBS 0.034079f
C1144 VP.n58 VSUBS 0.054725f
C1145 VP.n59 VSUBS 0.040734f
C1146 VP.n60 VSUBS 0.993673f
C1147 VP.n61 VSUBS 0.059545f
C1148 VP.n62 VSUBS 0.034079f
C1149 VP.n63 VSUBS 0.034079f
C1150 VP.n64 VSUBS 0.034079f
C1151 VP.n65 VSUBS 0.063197f
C1152 VP.n66 VSUBS 0.03387f
C1153 VP.n67 VSUBS 1.05386f
C1154 VP.n68 VSUBS 0.035036f
.ends

