* NGSPICE file created from diff_pair_sample_1208.ext - technology: sky130A

.subckt diff_pair_sample_1208 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X1 VDD1.t7 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=3.8844 ps=20.7 w=9.96 l=1.05
X2 VDD1.t6 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=3.8844 ps=20.7 w=9.96 l=1.05
X3 VTAIL.t14 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=1.6434 ps=10.29 w=9.96 l=1.05
X4 VDD2.t5 VN.t2 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X5 VTAIL.t3 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=1.6434 ps=10.29 w=9.96 l=1.05
X6 VDD2.t4 VN.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=3.8844 ps=20.7 w=9.96 l=1.05
X7 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X8 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=0 ps=0 w=9.96 l=1.05
X9 VTAIL.t11 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X10 VDD1.t3 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X11 VDD2.t7 VN.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X12 VDD2.t2 VN.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=3.8844 ps=20.7 w=9.96 l=1.05
X13 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=0 ps=0 w=9.96 l=1.05
X14 VTAIL.t2 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=1.6434 ps=10.29 w=9.96 l=1.05
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=0 ps=0 w=9.96 l=1.05
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=0 ps=0 w=9.96 l=1.05
X17 VTAIL.t5 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X18 VDD1.t0 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6434 pd=10.29 as=1.6434 ps=10.29 w=9.96 l=1.05
X19 VTAIL.t8 VN.t7 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8844 pd=20.7 as=1.6434 ps=10.29 w=9.96 l=1.05
R0 VN.n3 VN.t7 287.925
R1 VN.n16 VN.t6 287.925
R2 VN.n11 VN.t3 266.478
R3 VN.n24 VN.t1 266.478
R4 VN.n4 VN.t5 228.607
R5 VN.n1 VN.t0 228.607
R6 VN.n17 VN.t4 228.607
R7 VN.n14 VN.t2 228.607
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.4773
R19 VN.n19 VN.n18 56.4773
R20 VN.n11 VN.n10 43.0884
R21 VN.n24 VN.n23 43.0884
R22 VN VN.n25 42.4763
R23 VN.n4 VN.n3 35.3356
R24 VN.n17 VN.n16 35.3356
R25 VN.n16 VN.n15 28.7542
R26 VN.n3 VN.n2 28.7542
R27 VN.n10 VN.n9 27.752
R28 VN.n23 VN.n22 27.752
R29 VN.n5 VN.n4 21.4227
R30 VN.n6 VN.n1 21.4227
R31 VN.n18 VN.n17 21.4227
R32 VN.n19 VN.n14 21.4227
R33 VN.n9 VN.n1 2.92171
R34 VN.n22 VN.n14 2.92171
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 63.1796
R45 VDD2.n2 VDD2.n0 63.1796
R46 VDD2 VDD2.n5 63.1768
R47 VDD2.n4 VDD2.n3 62.6403
R48 VDD2.n4 VDD2.n2 37.6549
R49 VDD2.n5 VDD2.t1 1.98845
R50 VDD2.n5 VDD2.t2 1.98845
R51 VDD2.n3 VDD2.t6 1.98845
R52 VDD2.n3 VDD2.t5 1.98845
R53 VDD2.n1 VDD2.t0 1.98845
R54 VDD2.n1 VDD2.t4 1.98845
R55 VDD2.n0 VDD2.t3 1.98845
R56 VDD2.n0 VDD2.t7 1.98845
R57 VDD2 VDD2.n4 0.653517
R58 VTAIL.n434 VTAIL.n386 289.615
R59 VTAIL.n50 VTAIL.n2 289.615
R60 VTAIL.n104 VTAIL.n56 289.615
R61 VTAIL.n160 VTAIL.n112 289.615
R62 VTAIL.n380 VTAIL.n332 289.615
R63 VTAIL.n324 VTAIL.n276 289.615
R64 VTAIL.n270 VTAIL.n222 289.615
R65 VTAIL.n214 VTAIL.n166 289.615
R66 VTAIL.n402 VTAIL.n401 185
R67 VTAIL.n407 VTAIL.n406 185
R68 VTAIL.n409 VTAIL.n408 185
R69 VTAIL.n398 VTAIL.n397 185
R70 VTAIL.n415 VTAIL.n414 185
R71 VTAIL.n417 VTAIL.n416 185
R72 VTAIL.n394 VTAIL.n393 185
R73 VTAIL.n424 VTAIL.n423 185
R74 VTAIL.n425 VTAIL.n392 185
R75 VTAIL.n427 VTAIL.n426 185
R76 VTAIL.n390 VTAIL.n389 185
R77 VTAIL.n433 VTAIL.n432 185
R78 VTAIL.n435 VTAIL.n434 185
R79 VTAIL.n18 VTAIL.n17 185
R80 VTAIL.n23 VTAIL.n22 185
R81 VTAIL.n25 VTAIL.n24 185
R82 VTAIL.n14 VTAIL.n13 185
R83 VTAIL.n31 VTAIL.n30 185
R84 VTAIL.n33 VTAIL.n32 185
R85 VTAIL.n10 VTAIL.n9 185
R86 VTAIL.n40 VTAIL.n39 185
R87 VTAIL.n41 VTAIL.n8 185
R88 VTAIL.n43 VTAIL.n42 185
R89 VTAIL.n6 VTAIL.n5 185
R90 VTAIL.n49 VTAIL.n48 185
R91 VTAIL.n51 VTAIL.n50 185
R92 VTAIL.n72 VTAIL.n71 185
R93 VTAIL.n77 VTAIL.n76 185
R94 VTAIL.n79 VTAIL.n78 185
R95 VTAIL.n68 VTAIL.n67 185
R96 VTAIL.n85 VTAIL.n84 185
R97 VTAIL.n87 VTAIL.n86 185
R98 VTAIL.n64 VTAIL.n63 185
R99 VTAIL.n94 VTAIL.n93 185
R100 VTAIL.n95 VTAIL.n62 185
R101 VTAIL.n97 VTAIL.n96 185
R102 VTAIL.n60 VTAIL.n59 185
R103 VTAIL.n103 VTAIL.n102 185
R104 VTAIL.n105 VTAIL.n104 185
R105 VTAIL.n128 VTAIL.n127 185
R106 VTAIL.n133 VTAIL.n132 185
R107 VTAIL.n135 VTAIL.n134 185
R108 VTAIL.n124 VTAIL.n123 185
R109 VTAIL.n141 VTAIL.n140 185
R110 VTAIL.n143 VTAIL.n142 185
R111 VTAIL.n120 VTAIL.n119 185
R112 VTAIL.n150 VTAIL.n149 185
R113 VTAIL.n151 VTAIL.n118 185
R114 VTAIL.n153 VTAIL.n152 185
R115 VTAIL.n116 VTAIL.n115 185
R116 VTAIL.n159 VTAIL.n158 185
R117 VTAIL.n161 VTAIL.n160 185
R118 VTAIL.n381 VTAIL.n380 185
R119 VTAIL.n379 VTAIL.n378 185
R120 VTAIL.n336 VTAIL.n335 185
R121 VTAIL.n373 VTAIL.n372 185
R122 VTAIL.n371 VTAIL.n338 185
R123 VTAIL.n370 VTAIL.n369 185
R124 VTAIL.n341 VTAIL.n339 185
R125 VTAIL.n364 VTAIL.n363 185
R126 VTAIL.n362 VTAIL.n361 185
R127 VTAIL.n345 VTAIL.n344 185
R128 VTAIL.n356 VTAIL.n355 185
R129 VTAIL.n354 VTAIL.n353 185
R130 VTAIL.n349 VTAIL.n348 185
R131 VTAIL.n325 VTAIL.n324 185
R132 VTAIL.n323 VTAIL.n322 185
R133 VTAIL.n280 VTAIL.n279 185
R134 VTAIL.n317 VTAIL.n316 185
R135 VTAIL.n315 VTAIL.n282 185
R136 VTAIL.n314 VTAIL.n313 185
R137 VTAIL.n285 VTAIL.n283 185
R138 VTAIL.n308 VTAIL.n307 185
R139 VTAIL.n306 VTAIL.n305 185
R140 VTAIL.n289 VTAIL.n288 185
R141 VTAIL.n300 VTAIL.n299 185
R142 VTAIL.n298 VTAIL.n297 185
R143 VTAIL.n293 VTAIL.n292 185
R144 VTAIL.n271 VTAIL.n270 185
R145 VTAIL.n269 VTAIL.n268 185
R146 VTAIL.n226 VTAIL.n225 185
R147 VTAIL.n263 VTAIL.n262 185
R148 VTAIL.n261 VTAIL.n228 185
R149 VTAIL.n260 VTAIL.n259 185
R150 VTAIL.n231 VTAIL.n229 185
R151 VTAIL.n254 VTAIL.n253 185
R152 VTAIL.n252 VTAIL.n251 185
R153 VTAIL.n235 VTAIL.n234 185
R154 VTAIL.n246 VTAIL.n245 185
R155 VTAIL.n244 VTAIL.n243 185
R156 VTAIL.n239 VTAIL.n238 185
R157 VTAIL.n215 VTAIL.n214 185
R158 VTAIL.n213 VTAIL.n212 185
R159 VTAIL.n170 VTAIL.n169 185
R160 VTAIL.n207 VTAIL.n206 185
R161 VTAIL.n205 VTAIL.n172 185
R162 VTAIL.n204 VTAIL.n203 185
R163 VTAIL.n175 VTAIL.n173 185
R164 VTAIL.n198 VTAIL.n197 185
R165 VTAIL.n196 VTAIL.n195 185
R166 VTAIL.n179 VTAIL.n178 185
R167 VTAIL.n190 VTAIL.n189 185
R168 VTAIL.n188 VTAIL.n187 185
R169 VTAIL.n183 VTAIL.n182 185
R170 VTAIL.n403 VTAIL.t12 149.524
R171 VTAIL.n19 VTAIL.t8 149.524
R172 VTAIL.n73 VTAIL.t4 149.524
R173 VTAIL.n129 VTAIL.t3 149.524
R174 VTAIL.n350 VTAIL.t0 149.524
R175 VTAIL.n294 VTAIL.t2 149.524
R176 VTAIL.n240 VTAIL.t9 149.524
R177 VTAIL.n184 VTAIL.t14 149.524
R178 VTAIL.n407 VTAIL.n401 104.615
R179 VTAIL.n408 VTAIL.n407 104.615
R180 VTAIL.n408 VTAIL.n397 104.615
R181 VTAIL.n415 VTAIL.n397 104.615
R182 VTAIL.n416 VTAIL.n415 104.615
R183 VTAIL.n416 VTAIL.n393 104.615
R184 VTAIL.n424 VTAIL.n393 104.615
R185 VTAIL.n425 VTAIL.n424 104.615
R186 VTAIL.n426 VTAIL.n425 104.615
R187 VTAIL.n426 VTAIL.n389 104.615
R188 VTAIL.n433 VTAIL.n389 104.615
R189 VTAIL.n434 VTAIL.n433 104.615
R190 VTAIL.n23 VTAIL.n17 104.615
R191 VTAIL.n24 VTAIL.n23 104.615
R192 VTAIL.n24 VTAIL.n13 104.615
R193 VTAIL.n31 VTAIL.n13 104.615
R194 VTAIL.n32 VTAIL.n31 104.615
R195 VTAIL.n32 VTAIL.n9 104.615
R196 VTAIL.n40 VTAIL.n9 104.615
R197 VTAIL.n41 VTAIL.n40 104.615
R198 VTAIL.n42 VTAIL.n41 104.615
R199 VTAIL.n42 VTAIL.n5 104.615
R200 VTAIL.n49 VTAIL.n5 104.615
R201 VTAIL.n50 VTAIL.n49 104.615
R202 VTAIL.n77 VTAIL.n71 104.615
R203 VTAIL.n78 VTAIL.n77 104.615
R204 VTAIL.n78 VTAIL.n67 104.615
R205 VTAIL.n85 VTAIL.n67 104.615
R206 VTAIL.n86 VTAIL.n85 104.615
R207 VTAIL.n86 VTAIL.n63 104.615
R208 VTAIL.n94 VTAIL.n63 104.615
R209 VTAIL.n95 VTAIL.n94 104.615
R210 VTAIL.n96 VTAIL.n95 104.615
R211 VTAIL.n96 VTAIL.n59 104.615
R212 VTAIL.n103 VTAIL.n59 104.615
R213 VTAIL.n104 VTAIL.n103 104.615
R214 VTAIL.n133 VTAIL.n127 104.615
R215 VTAIL.n134 VTAIL.n133 104.615
R216 VTAIL.n134 VTAIL.n123 104.615
R217 VTAIL.n141 VTAIL.n123 104.615
R218 VTAIL.n142 VTAIL.n141 104.615
R219 VTAIL.n142 VTAIL.n119 104.615
R220 VTAIL.n150 VTAIL.n119 104.615
R221 VTAIL.n151 VTAIL.n150 104.615
R222 VTAIL.n152 VTAIL.n151 104.615
R223 VTAIL.n152 VTAIL.n115 104.615
R224 VTAIL.n159 VTAIL.n115 104.615
R225 VTAIL.n160 VTAIL.n159 104.615
R226 VTAIL.n380 VTAIL.n379 104.615
R227 VTAIL.n379 VTAIL.n335 104.615
R228 VTAIL.n372 VTAIL.n335 104.615
R229 VTAIL.n372 VTAIL.n371 104.615
R230 VTAIL.n371 VTAIL.n370 104.615
R231 VTAIL.n370 VTAIL.n339 104.615
R232 VTAIL.n363 VTAIL.n339 104.615
R233 VTAIL.n363 VTAIL.n362 104.615
R234 VTAIL.n362 VTAIL.n344 104.615
R235 VTAIL.n355 VTAIL.n344 104.615
R236 VTAIL.n355 VTAIL.n354 104.615
R237 VTAIL.n354 VTAIL.n348 104.615
R238 VTAIL.n324 VTAIL.n323 104.615
R239 VTAIL.n323 VTAIL.n279 104.615
R240 VTAIL.n316 VTAIL.n279 104.615
R241 VTAIL.n316 VTAIL.n315 104.615
R242 VTAIL.n315 VTAIL.n314 104.615
R243 VTAIL.n314 VTAIL.n283 104.615
R244 VTAIL.n307 VTAIL.n283 104.615
R245 VTAIL.n307 VTAIL.n306 104.615
R246 VTAIL.n306 VTAIL.n288 104.615
R247 VTAIL.n299 VTAIL.n288 104.615
R248 VTAIL.n299 VTAIL.n298 104.615
R249 VTAIL.n298 VTAIL.n292 104.615
R250 VTAIL.n270 VTAIL.n269 104.615
R251 VTAIL.n269 VTAIL.n225 104.615
R252 VTAIL.n262 VTAIL.n225 104.615
R253 VTAIL.n262 VTAIL.n261 104.615
R254 VTAIL.n261 VTAIL.n260 104.615
R255 VTAIL.n260 VTAIL.n229 104.615
R256 VTAIL.n253 VTAIL.n229 104.615
R257 VTAIL.n253 VTAIL.n252 104.615
R258 VTAIL.n252 VTAIL.n234 104.615
R259 VTAIL.n245 VTAIL.n234 104.615
R260 VTAIL.n245 VTAIL.n244 104.615
R261 VTAIL.n244 VTAIL.n238 104.615
R262 VTAIL.n214 VTAIL.n213 104.615
R263 VTAIL.n213 VTAIL.n169 104.615
R264 VTAIL.n206 VTAIL.n169 104.615
R265 VTAIL.n206 VTAIL.n205 104.615
R266 VTAIL.n205 VTAIL.n204 104.615
R267 VTAIL.n204 VTAIL.n173 104.615
R268 VTAIL.n197 VTAIL.n173 104.615
R269 VTAIL.n197 VTAIL.n196 104.615
R270 VTAIL.n196 VTAIL.n178 104.615
R271 VTAIL.n189 VTAIL.n178 104.615
R272 VTAIL.n189 VTAIL.n188 104.615
R273 VTAIL.n188 VTAIL.n182 104.615
R274 VTAIL.t12 VTAIL.n401 52.3082
R275 VTAIL.t8 VTAIL.n17 52.3082
R276 VTAIL.t4 VTAIL.n71 52.3082
R277 VTAIL.t3 VTAIL.n127 52.3082
R278 VTAIL.t0 VTAIL.n348 52.3082
R279 VTAIL.t2 VTAIL.n292 52.3082
R280 VTAIL.t9 VTAIL.n238 52.3082
R281 VTAIL.t14 VTAIL.n182 52.3082
R282 VTAIL.n331 VTAIL.n330 45.9615
R283 VTAIL.n221 VTAIL.n220 45.9615
R284 VTAIL.n1 VTAIL.n0 45.9614
R285 VTAIL.n111 VTAIL.n110 45.9614
R286 VTAIL.n439 VTAIL.n438 32.1853
R287 VTAIL.n55 VTAIL.n54 32.1853
R288 VTAIL.n109 VTAIL.n108 32.1853
R289 VTAIL.n165 VTAIL.n164 32.1853
R290 VTAIL.n385 VTAIL.n384 32.1853
R291 VTAIL.n329 VTAIL.n328 32.1853
R292 VTAIL.n275 VTAIL.n274 32.1853
R293 VTAIL.n219 VTAIL.n218 32.1853
R294 VTAIL.n439 VTAIL.n385 22.1427
R295 VTAIL.n219 VTAIL.n165 22.1427
R296 VTAIL.n427 VTAIL.n392 13.1884
R297 VTAIL.n43 VTAIL.n8 13.1884
R298 VTAIL.n97 VTAIL.n62 13.1884
R299 VTAIL.n153 VTAIL.n118 13.1884
R300 VTAIL.n373 VTAIL.n338 13.1884
R301 VTAIL.n317 VTAIL.n282 13.1884
R302 VTAIL.n263 VTAIL.n228 13.1884
R303 VTAIL.n207 VTAIL.n172 13.1884
R304 VTAIL.n423 VTAIL.n422 12.8005
R305 VTAIL.n428 VTAIL.n390 12.8005
R306 VTAIL.n39 VTAIL.n38 12.8005
R307 VTAIL.n44 VTAIL.n6 12.8005
R308 VTAIL.n93 VTAIL.n92 12.8005
R309 VTAIL.n98 VTAIL.n60 12.8005
R310 VTAIL.n149 VTAIL.n148 12.8005
R311 VTAIL.n154 VTAIL.n116 12.8005
R312 VTAIL.n374 VTAIL.n336 12.8005
R313 VTAIL.n369 VTAIL.n340 12.8005
R314 VTAIL.n318 VTAIL.n280 12.8005
R315 VTAIL.n313 VTAIL.n284 12.8005
R316 VTAIL.n264 VTAIL.n226 12.8005
R317 VTAIL.n259 VTAIL.n230 12.8005
R318 VTAIL.n208 VTAIL.n170 12.8005
R319 VTAIL.n203 VTAIL.n174 12.8005
R320 VTAIL.n421 VTAIL.n394 12.0247
R321 VTAIL.n432 VTAIL.n431 12.0247
R322 VTAIL.n37 VTAIL.n10 12.0247
R323 VTAIL.n48 VTAIL.n47 12.0247
R324 VTAIL.n91 VTAIL.n64 12.0247
R325 VTAIL.n102 VTAIL.n101 12.0247
R326 VTAIL.n147 VTAIL.n120 12.0247
R327 VTAIL.n158 VTAIL.n157 12.0247
R328 VTAIL.n378 VTAIL.n377 12.0247
R329 VTAIL.n368 VTAIL.n341 12.0247
R330 VTAIL.n322 VTAIL.n321 12.0247
R331 VTAIL.n312 VTAIL.n285 12.0247
R332 VTAIL.n268 VTAIL.n267 12.0247
R333 VTAIL.n258 VTAIL.n231 12.0247
R334 VTAIL.n212 VTAIL.n211 12.0247
R335 VTAIL.n202 VTAIL.n175 12.0247
R336 VTAIL.n418 VTAIL.n417 11.249
R337 VTAIL.n435 VTAIL.n388 11.249
R338 VTAIL.n34 VTAIL.n33 11.249
R339 VTAIL.n51 VTAIL.n4 11.249
R340 VTAIL.n88 VTAIL.n87 11.249
R341 VTAIL.n105 VTAIL.n58 11.249
R342 VTAIL.n144 VTAIL.n143 11.249
R343 VTAIL.n161 VTAIL.n114 11.249
R344 VTAIL.n381 VTAIL.n334 11.249
R345 VTAIL.n365 VTAIL.n364 11.249
R346 VTAIL.n325 VTAIL.n278 11.249
R347 VTAIL.n309 VTAIL.n308 11.249
R348 VTAIL.n271 VTAIL.n224 11.249
R349 VTAIL.n255 VTAIL.n254 11.249
R350 VTAIL.n215 VTAIL.n168 11.249
R351 VTAIL.n199 VTAIL.n198 11.249
R352 VTAIL.n414 VTAIL.n396 10.4732
R353 VTAIL.n436 VTAIL.n386 10.4732
R354 VTAIL.n30 VTAIL.n12 10.4732
R355 VTAIL.n52 VTAIL.n2 10.4732
R356 VTAIL.n84 VTAIL.n66 10.4732
R357 VTAIL.n106 VTAIL.n56 10.4732
R358 VTAIL.n140 VTAIL.n122 10.4732
R359 VTAIL.n162 VTAIL.n112 10.4732
R360 VTAIL.n382 VTAIL.n332 10.4732
R361 VTAIL.n361 VTAIL.n343 10.4732
R362 VTAIL.n326 VTAIL.n276 10.4732
R363 VTAIL.n305 VTAIL.n287 10.4732
R364 VTAIL.n272 VTAIL.n222 10.4732
R365 VTAIL.n251 VTAIL.n233 10.4732
R366 VTAIL.n216 VTAIL.n166 10.4732
R367 VTAIL.n195 VTAIL.n177 10.4732
R368 VTAIL.n403 VTAIL.n402 10.2747
R369 VTAIL.n19 VTAIL.n18 10.2747
R370 VTAIL.n73 VTAIL.n72 10.2747
R371 VTAIL.n129 VTAIL.n128 10.2747
R372 VTAIL.n350 VTAIL.n349 10.2747
R373 VTAIL.n294 VTAIL.n293 10.2747
R374 VTAIL.n240 VTAIL.n239 10.2747
R375 VTAIL.n184 VTAIL.n183 10.2747
R376 VTAIL.n413 VTAIL.n398 9.69747
R377 VTAIL.n29 VTAIL.n14 9.69747
R378 VTAIL.n83 VTAIL.n68 9.69747
R379 VTAIL.n139 VTAIL.n124 9.69747
R380 VTAIL.n360 VTAIL.n345 9.69747
R381 VTAIL.n304 VTAIL.n289 9.69747
R382 VTAIL.n250 VTAIL.n235 9.69747
R383 VTAIL.n194 VTAIL.n179 9.69747
R384 VTAIL.n438 VTAIL.n437 9.45567
R385 VTAIL.n54 VTAIL.n53 9.45567
R386 VTAIL.n108 VTAIL.n107 9.45567
R387 VTAIL.n164 VTAIL.n163 9.45567
R388 VTAIL.n384 VTAIL.n383 9.45567
R389 VTAIL.n328 VTAIL.n327 9.45567
R390 VTAIL.n274 VTAIL.n273 9.45567
R391 VTAIL.n218 VTAIL.n217 9.45567
R392 VTAIL.n437 VTAIL.n436 9.3005
R393 VTAIL.n388 VTAIL.n387 9.3005
R394 VTAIL.n431 VTAIL.n430 9.3005
R395 VTAIL.n429 VTAIL.n428 9.3005
R396 VTAIL.n405 VTAIL.n404 9.3005
R397 VTAIL.n400 VTAIL.n399 9.3005
R398 VTAIL.n411 VTAIL.n410 9.3005
R399 VTAIL.n413 VTAIL.n412 9.3005
R400 VTAIL.n396 VTAIL.n395 9.3005
R401 VTAIL.n419 VTAIL.n418 9.3005
R402 VTAIL.n421 VTAIL.n420 9.3005
R403 VTAIL.n422 VTAIL.n391 9.3005
R404 VTAIL.n53 VTAIL.n52 9.3005
R405 VTAIL.n4 VTAIL.n3 9.3005
R406 VTAIL.n47 VTAIL.n46 9.3005
R407 VTAIL.n45 VTAIL.n44 9.3005
R408 VTAIL.n21 VTAIL.n20 9.3005
R409 VTAIL.n16 VTAIL.n15 9.3005
R410 VTAIL.n27 VTAIL.n26 9.3005
R411 VTAIL.n29 VTAIL.n28 9.3005
R412 VTAIL.n12 VTAIL.n11 9.3005
R413 VTAIL.n35 VTAIL.n34 9.3005
R414 VTAIL.n37 VTAIL.n36 9.3005
R415 VTAIL.n38 VTAIL.n7 9.3005
R416 VTAIL.n107 VTAIL.n106 9.3005
R417 VTAIL.n58 VTAIL.n57 9.3005
R418 VTAIL.n101 VTAIL.n100 9.3005
R419 VTAIL.n99 VTAIL.n98 9.3005
R420 VTAIL.n75 VTAIL.n74 9.3005
R421 VTAIL.n70 VTAIL.n69 9.3005
R422 VTAIL.n81 VTAIL.n80 9.3005
R423 VTAIL.n83 VTAIL.n82 9.3005
R424 VTAIL.n66 VTAIL.n65 9.3005
R425 VTAIL.n89 VTAIL.n88 9.3005
R426 VTAIL.n91 VTAIL.n90 9.3005
R427 VTAIL.n92 VTAIL.n61 9.3005
R428 VTAIL.n163 VTAIL.n162 9.3005
R429 VTAIL.n114 VTAIL.n113 9.3005
R430 VTAIL.n157 VTAIL.n156 9.3005
R431 VTAIL.n155 VTAIL.n154 9.3005
R432 VTAIL.n131 VTAIL.n130 9.3005
R433 VTAIL.n126 VTAIL.n125 9.3005
R434 VTAIL.n137 VTAIL.n136 9.3005
R435 VTAIL.n139 VTAIL.n138 9.3005
R436 VTAIL.n122 VTAIL.n121 9.3005
R437 VTAIL.n145 VTAIL.n144 9.3005
R438 VTAIL.n147 VTAIL.n146 9.3005
R439 VTAIL.n148 VTAIL.n117 9.3005
R440 VTAIL.n352 VTAIL.n351 9.3005
R441 VTAIL.n347 VTAIL.n346 9.3005
R442 VTAIL.n358 VTAIL.n357 9.3005
R443 VTAIL.n360 VTAIL.n359 9.3005
R444 VTAIL.n343 VTAIL.n342 9.3005
R445 VTAIL.n366 VTAIL.n365 9.3005
R446 VTAIL.n368 VTAIL.n367 9.3005
R447 VTAIL.n340 VTAIL.n337 9.3005
R448 VTAIL.n383 VTAIL.n382 9.3005
R449 VTAIL.n334 VTAIL.n333 9.3005
R450 VTAIL.n377 VTAIL.n376 9.3005
R451 VTAIL.n375 VTAIL.n374 9.3005
R452 VTAIL.n296 VTAIL.n295 9.3005
R453 VTAIL.n291 VTAIL.n290 9.3005
R454 VTAIL.n302 VTAIL.n301 9.3005
R455 VTAIL.n304 VTAIL.n303 9.3005
R456 VTAIL.n287 VTAIL.n286 9.3005
R457 VTAIL.n310 VTAIL.n309 9.3005
R458 VTAIL.n312 VTAIL.n311 9.3005
R459 VTAIL.n284 VTAIL.n281 9.3005
R460 VTAIL.n327 VTAIL.n326 9.3005
R461 VTAIL.n278 VTAIL.n277 9.3005
R462 VTAIL.n321 VTAIL.n320 9.3005
R463 VTAIL.n319 VTAIL.n318 9.3005
R464 VTAIL.n242 VTAIL.n241 9.3005
R465 VTAIL.n237 VTAIL.n236 9.3005
R466 VTAIL.n248 VTAIL.n247 9.3005
R467 VTAIL.n250 VTAIL.n249 9.3005
R468 VTAIL.n233 VTAIL.n232 9.3005
R469 VTAIL.n256 VTAIL.n255 9.3005
R470 VTAIL.n258 VTAIL.n257 9.3005
R471 VTAIL.n230 VTAIL.n227 9.3005
R472 VTAIL.n273 VTAIL.n272 9.3005
R473 VTAIL.n224 VTAIL.n223 9.3005
R474 VTAIL.n267 VTAIL.n266 9.3005
R475 VTAIL.n265 VTAIL.n264 9.3005
R476 VTAIL.n186 VTAIL.n185 9.3005
R477 VTAIL.n181 VTAIL.n180 9.3005
R478 VTAIL.n192 VTAIL.n191 9.3005
R479 VTAIL.n194 VTAIL.n193 9.3005
R480 VTAIL.n177 VTAIL.n176 9.3005
R481 VTAIL.n200 VTAIL.n199 9.3005
R482 VTAIL.n202 VTAIL.n201 9.3005
R483 VTAIL.n174 VTAIL.n171 9.3005
R484 VTAIL.n217 VTAIL.n216 9.3005
R485 VTAIL.n168 VTAIL.n167 9.3005
R486 VTAIL.n211 VTAIL.n210 9.3005
R487 VTAIL.n209 VTAIL.n208 9.3005
R488 VTAIL.n410 VTAIL.n409 8.92171
R489 VTAIL.n26 VTAIL.n25 8.92171
R490 VTAIL.n80 VTAIL.n79 8.92171
R491 VTAIL.n136 VTAIL.n135 8.92171
R492 VTAIL.n357 VTAIL.n356 8.92171
R493 VTAIL.n301 VTAIL.n300 8.92171
R494 VTAIL.n247 VTAIL.n246 8.92171
R495 VTAIL.n191 VTAIL.n190 8.92171
R496 VTAIL.n406 VTAIL.n400 8.14595
R497 VTAIL.n22 VTAIL.n16 8.14595
R498 VTAIL.n76 VTAIL.n70 8.14595
R499 VTAIL.n132 VTAIL.n126 8.14595
R500 VTAIL.n353 VTAIL.n347 8.14595
R501 VTAIL.n297 VTAIL.n291 8.14595
R502 VTAIL.n243 VTAIL.n237 8.14595
R503 VTAIL.n187 VTAIL.n181 8.14595
R504 VTAIL.n405 VTAIL.n402 7.3702
R505 VTAIL.n21 VTAIL.n18 7.3702
R506 VTAIL.n75 VTAIL.n72 7.3702
R507 VTAIL.n131 VTAIL.n128 7.3702
R508 VTAIL.n352 VTAIL.n349 7.3702
R509 VTAIL.n296 VTAIL.n293 7.3702
R510 VTAIL.n242 VTAIL.n239 7.3702
R511 VTAIL.n186 VTAIL.n183 7.3702
R512 VTAIL.n406 VTAIL.n405 5.81868
R513 VTAIL.n22 VTAIL.n21 5.81868
R514 VTAIL.n76 VTAIL.n75 5.81868
R515 VTAIL.n132 VTAIL.n131 5.81868
R516 VTAIL.n353 VTAIL.n352 5.81868
R517 VTAIL.n297 VTAIL.n296 5.81868
R518 VTAIL.n243 VTAIL.n242 5.81868
R519 VTAIL.n187 VTAIL.n186 5.81868
R520 VTAIL.n409 VTAIL.n400 5.04292
R521 VTAIL.n25 VTAIL.n16 5.04292
R522 VTAIL.n79 VTAIL.n70 5.04292
R523 VTAIL.n135 VTAIL.n126 5.04292
R524 VTAIL.n356 VTAIL.n347 5.04292
R525 VTAIL.n300 VTAIL.n291 5.04292
R526 VTAIL.n246 VTAIL.n237 5.04292
R527 VTAIL.n190 VTAIL.n181 5.04292
R528 VTAIL.n410 VTAIL.n398 4.26717
R529 VTAIL.n26 VTAIL.n14 4.26717
R530 VTAIL.n80 VTAIL.n68 4.26717
R531 VTAIL.n136 VTAIL.n124 4.26717
R532 VTAIL.n357 VTAIL.n345 4.26717
R533 VTAIL.n301 VTAIL.n289 4.26717
R534 VTAIL.n247 VTAIL.n235 4.26717
R535 VTAIL.n191 VTAIL.n179 4.26717
R536 VTAIL.n414 VTAIL.n413 3.49141
R537 VTAIL.n438 VTAIL.n386 3.49141
R538 VTAIL.n30 VTAIL.n29 3.49141
R539 VTAIL.n54 VTAIL.n2 3.49141
R540 VTAIL.n84 VTAIL.n83 3.49141
R541 VTAIL.n108 VTAIL.n56 3.49141
R542 VTAIL.n140 VTAIL.n139 3.49141
R543 VTAIL.n164 VTAIL.n112 3.49141
R544 VTAIL.n384 VTAIL.n332 3.49141
R545 VTAIL.n361 VTAIL.n360 3.49141
R546 VTAIL.n328 VTAIL.n276 3.49141
R547 VTAIL.n305 VTAIL.n304 3.49141
R548 VTAIL.n274 VTAIL.n222 3.49141
R549 VTAIL.n251 VTAIL.n250 3.49141
R550 VTAIL.n218 VTAIL.n166 3.49141
R551 VTAIL.n195 VTAIL.n194 3.49141
R552 VTAIL.n404 VTAIL.n403 2.84303
R553 VTAIL.n20 VTAIL.n19 2.84303
R554 VTAIL.n74 VTAIL.n73 2.84303
R555 VTAIL.n130 VTAIL.n129 2.84303
R556 VTAIL.n351 VTAIL.n350 2.84303
R557 VTAIL.n295 VTAIL.n294 2.84303
R558 VTAIL.n241 VTAIL.n240 2.84303
R559 VTAIL.n185 VTAIL.n184 2.84303
R560 VTAIL.n417 VTAIL.n396 2.71565
R561 VTAIL.n436 VTAIL.n435 2.71565
R562 VTAIL.n33 VTAIL.n12 2.71565
R563 VTAIL.n52 VTAIL.n51 2.71565
R564 VTAIL.n87 VTAIL.n66 2.71565
R565 VTAIL.n106 VTAIL.n105 2.71565
R566 VTAIL.n143 VTAIL.n122 2.71565
R567 VTAIL.n162 VTAIL.n161 2.71565
R568 VTAIL.n382 VTAIL.n381 2.71565
R569 VTAIL.n364 VTAIL.n343 2.71565
R570 VTAIL.n326 VTAIL.n325 2.71565
R571 VTAIL.n308 VTAIL.n287 2.71565
R572 VTAIL.n272 VTAIL.n271 2.71565
R573 VTAIL.n254 VTAIL.n233 2.71565
R574 VTAIL.n216 VTAIL.n215 2.71565
R575 VTAIL.n198 VTAIL.n177 2.71565
R576 VTAIL.n0 VTAIL.t10 1.98845
R577 VTAIL.n0 VTAIL.t15 1.98845
R578 VTAIL.n110 VTAIL.t1 1.98845
R579 VTAIL.n110 VTAIL.t5 1.98845
R580 VTAIL.n330 VTAIL.t6 1.98845
R581 VTAIL.n330 VTAIL.t7 1.98845
R582 VTAIL.n220 VTAIL.t13 1.98845
R583 VTAIL.n220 VTAIL.t11 1.98845
R584 VTAIL.n418 VTAIL.n394 1.93989
R585 VTAIL.n432 VTAIL.n388 1.93989
R586 VTAIL.n34 VTAIL.n10 1.93989
R587 VTAIL.n48 VTAIL.n4 1.93989
R588 VTAIL.n88 VTAIL.n64 1.93989
R589 VTAIL.n102 VTAIL.n58 1.93989
R590 VTAIL.n144 VTAIL.n120 1.93989
R591 VTAIL.n158 VTAIL.n114 1.93989
R592 VTAIL.n378 VTAIL.n334 1.93989
R593 VTAIL.n365 VTAIL.n341 1.93989
R594 VTAIL.n322 VTAIL.n278 1.93989
R595 VTAIL.n309 VTAIL.n285 1.93989
R596 VTAIL.n268 VTAIL.n224 1.93989
R597 VTAIL.n255 VTAIL.n231 1.93989
R598 VTAIL.n212 VTAIL.n168 1.93989
R599 VTAIL.n199 VTAIL.n175 1.93989
R600 VTAIL.n221 VTAIL.n219 1.19016
R601 VTAIL.n275 VTAIL.n221 1.19016
R602 VTAIL.n331 VTAIL.n329 1.19016
R603 VTAIL.n385 VTAIL.n331 1.19016
R604 VTAIL.n165 VTAIL.n111 1.19016
R605 VTAIL.n111 VTAIL.n109 1.19016
R606 VTAIL.n55 VTAIL.n1 1.19016
R607 VTAIL.n423 VTAIL.n421 1.16414
R608 VTAIL.n431 VTAIL.n390 1.16414
R609 VTAIL.n39 VTAIL.n37 1.16414
R610 VTAIL.n47 VTAIL.n6 1.16414
R611 VTAIL.n93 VTAIL.n91 1.16414
R612 VTAIL.n101 VTAIL.n60 1.16414
R613 VTAIL.n149 VTAIL.n147 1.16414
R614 VTAIL.n157 VTAIL.n116 1.16414
R615 VTAIL.n377 VTAIL.n336 1.16414
R616 VTAIL.n369 VTAIL.n368 1.16414
R617 VTAIL.n321 VTAIL.n280 1.16414
R618 VTAIL.n313 VTAIL.n312 1.16414
R619 VTAIL.n267 VTAIL.n226 1.16414
R620 VTAIL.n259 VTAIL.n258 1.16414
R621 VTAIL.n211 VTAIL.n170 1.16414
R622 VTAIL.n203 VTAIL.n202 1.16414
R623 VTAIL VTAIL.n439 1.13197
R624 VTAIL.n329 VTAIL.n275 0.470328
R625 VTAIL.n109 VTAIL.n55 0.470328
R626 VTAIL.n422 VTAIL.n392 0.388379
R627 VTAIL.n428 VTAIL.n427 0.388379
R628 VTAIL.n38 VTAIL.n8 0.388379
R629 VTAIL.n44 VTAIL.n43 0.388379
R630 VTAIL.n92 VTAIL.n62 0.388379
R631 VTAIL.n98 VTAIL.n97 0.388379
R632 VTAIL.n148 VTAIL.n118 0.388379
R633 VTAIL.n154 VTAIL.n153 0.388379
R634 VTAIL.n374 VTAIL.n373 0.388379
R635 VTAIL.n340 VTAIL.n338 0.388379
R636 VTAIL.n318 VTAIL.n317 0.388379
R637 VTAIL.n284 VTAIL.n282 0.388379
R638 VTAIL.n264 VTAIL.n263 0.388379
R639 VTAIL.n230 VTAIL.n228 0.388379
R640 VTAIL.n208 VTAIL.n207 0.388379
R641 VTAIL.n174 VTAIL.n172 0.388379
R642 VTAIL.n404 VTAIL.n399 0.155672
R643 VTAIL.n411 VTAIL.n399 0.155672
R644 VTAIL.n412 VTAIL.n411 0.155672
R645 VTAIL.n412 VTAIL.n395 0.155672
R646 VTAIL.n419 VTAIL.n395 0.155672
R647 VTAIL.n420 VTAIL.n419 0.155672
R648 VTAIL.n420 VTAIL.n391 0.155672
R649 VTAIL.n429 VTAIL.n391 0.155672
R650 VTAIL.n430 VTAIL.n429 0.155672
R651 VTAIL.n430 VTAIL.n387 0.155672
R652 VTAIL.n437 VTAIL.n387 0.155672
R653 VTAIL.n20 VTAIL.n15 0.155672
R654 VTAIL.n27 VTAIL.n15 0.155672
R655 VTAIL.n28 VTAIL.n27 0.155672
R656 VTAIL.n28 VTAIL.n11 0.155672
R657 VTAIL.n35 VTAIL.n11 0.155672
R658 VTAIL.n36 VTAIL.n35 0.155672
R659 VTAIL.n36 VTAIL.n7 0.155672
R660 VTAIL.n45 VTAIL.n7 0.155672
R661 VTAIL.n46 VTAIL.n45 0.155672
R662 VTAIL.n46 VTAIL.n3 0.155672
R663 VTAIL.n53 VTAIL.n3 0.155672
R664 VTAIL.n74 VTAIL.n69 0.155672
R665 VTAIL.n81 VTAIL.n69 0.155672
R666 VTAIL.n82 VTAIL.n81 0.155672
R667 VTAIL.n82 VTAIL.n65 0.155672
R668 VTAIL.n89 VTAIL.n65 0.155672
R669 VTAIL.n90 VTAIL.n89 0.155672
R670 VTAIL.n90 VTAIL.n61 0.155672
R671 VTAIL.n99 VTAIL.n61 0.155672
R672 VTAIL.n100 VTAIL.n99 0.155672
R673 VTAIL.n100 VTAIL.n57 0.155672
R674 VTAIL.n107 VTAIL.n57 0.155672
R675 VTAIL.n130 VTAIL.n125 0.155672
R676 VTAIL.n137 VTAIL.n125 0.155672
R677 VTAIL.n138 VTAIL.n137 0.155672
R678 VTAIL.n138 VTAIL.n121 0.155672
R679 VTAIL.n145 VTAIL.n121 0.155672
R680 VTAIL.n146 VTAIL.n145 0.155672
R681 VTAIL.n146 VTAIL.n117 0.155672
R682 VTAIL.n155 VTAIL.n117 0.155672
R683 VTAIL.n156 VTAIL.n155 0.155672
R684 VTAIL.n156 VTAIL.n113 0.155672
R685 VTAIL.n163 VTAIL.n113 0.155672
R686 VTAIL.n383 VTAIL.n333 0.155672
R687 VTAIL.n376 VTAIL.n333 0.155672
R688 VTAIL.n376 VTAIL.n375 0.155672
R689 VTAIL.n375 VTAIL.n337 0.155672
R690 VTAIL.n367 VTAIL.n337 0.155672
R691 VTAIL.n367 VTAIL.n366 0.155672
R692 VTAIL.n366 VTAIL.n342 0.155672
R693 VTAIL.n359 VTAIL.n342 0.155672
R694 VTAIL.n359 VTAIL.n358 0.155672
R695 VTAIL.n358 VTAIL.n346 0.155672
R696 VTAIL.n351 VTAIL.n346 0.155672
R697 VTAIL.n327 VTAIL.n277 0.155672
R698 VTAIL.n320 VTAIL.n277 0.155672
R699 VTAIL.n320 VTAIL.n319 0.155672
R700 VTAIL.n319 VTAIL.n281 0.155672
R701 VTAIL.n311 VTAIL.n281 0.155672
R702 VTAIL.n311 VTAIL.n310 0.155672
R703 VTAIL.n310 VTAIL.n286 0.155672
R704 VTAIL.n303 VTAIL.n286 0.155672
R705 VTAIL.n303 VTAIL.n302 0.155672
R706 VTAIL.n302 VTAIL.n290 0.155672
R707 VTAIL.n295 VTAIL.n290 0.155672
R708 VTAIL.n273 VTAIL.n223 0.155672
R709 VTAIL.n266 VTAIL.n223 0.155672
R710 VTAIL.n266 VTAIL.n265 0.155672
R711 VTAIL.n265 VTAIL.n227 0.155672
R712 VTAIL.n257 VTAIL.n227 0.155672
R713 VTAIL.n257 VTAIL.n256 0.155672
R714 VTAIL.n256 VTAIL.n232 0.155672
R715 VTAIL.n249 VTAIL.n232 0.155672
R716 VTAIL.n249 VTAIL.n248 0.155672
R717 VTAIL.n248 VTAIL.n236 0.155672
R718 VTAIL.n241 VTAIL.n236 0.155672
R719 VTAIL.n217 VTAIL.n167 0.155672
R720 VTAIL.n210 VTAIL.n167 0.155672
R721 VTAIL.n210 VTAIL.n209 0.155672
R722 VTAIL.n209 VTAIL.n171 0.155672
R723 VTAIL.n201 VTAIL.n171 0.155672
R724 VTAIL.n201 VTAIL.n200 0.155672
R725 VTAIL.n200 VTAIL.n176 0.155672
R726 VTAIL.n193 VTAIL.n176 0.155672
R727 VTAIL.n193 VTAIL.n192 0.155672
R728 VTAIL.n192 VTAIL.n180 0.155672
R729 VTAIL.n185 VTAIL.n180 0.155672
R730 VTAIL VTAIL.n1 0.0586897
R731 B.n645 B.n644 585
R732 B.n646 B.n645 585
R733 B.n258 B.n95 585
R734 B.n257 B.n256 585
R735 B.n255 B.n254 585
R736 B.n253 B.n252 585
R737 B.n251 B.n250 585
R738 B.n249 B.n248 585
R739 B.n247 B.n246 585
R740 B.n245 B.n244 585
R741 B.n243 B.n242 585
R742 B.n241 B.n240 585
R743 B.n239 B.n238 585
R744 B.n237 B.n236 585
R745 B.n235 B.n234 585
R746 B.n233 B.n232 585
R747 B.n231 B.n230 585
R748 B.n229 B.n228 585
R749 B.n227 B.n226 585
R750 B.n225 B.n224 585
R751 B.n223 B.n222 585
R752 B.n221 B.n220 585
R753 B.n219 B.n218 585
R754 B.n217 B.n216 585
R755 B.n215 B.n214 585
R756 B.n213 B.n212 585
R757 B.n211 B.n210 585
R758 B.n209 B.n208 585
R759 B.n207 B.n206 585
R760 B.n205 B.n204 585
R761 B.n203 B.n202 585
R762 B.n201 B.n200 585
R763 B.n199 B.n198 585
R764 B.n197 B.n196 585
R765 B.n195 B.n194 585
R766 B.n193 B.n192 585
R767 B.n191 B.n190 585
R768 B.n188 B.n187 585
R769 B.n186 B.n185 585
R770 B.n184 B.n183 585
R771 B.n182 B.n181 585
R772 B.n180 B.n179 585
R773 B.n178 B.n177 585
R774 B.n176 B.n175 585
R775 B.n174 B.n173 585
R776 B.n172 B.n171 585
R777 B.n170 B.n169 585
R778 B.n168 B.n167 585
R779 B.n166 B.n165 585
R780 B.n164 B.n163 585
R781 B.n162 B.n161 585
R782 B.n160 B.n159 585
R783 B.n158 B.n157 585
R784 B.n156 B.n155 585
R785 B.n154 B.n153 585
R786 B.n152 B.n151 585
R787 B.n150 B.n149 585
R788 B.n148 B.n147 585
R789 B.n146 B.n145 585
R790 B.n144 B.n143 585
R791 B.n142 B.n141 585
R792 B.n140 B.n139 585
R793 B.n138 B.n137 585
R794 B.n136 B.n135 585
R795 B.n134 B.n133 585
R796 B.n132 B.n131 585
R797 B.n130 B.n129 585
R798 B.n128 B.n127 585
R799 B.n126 B.n125 585
R800 B.n124 B.n123 585
R801 B.n122 B.n121 585
R802 B.n120 B.n119 585
R803 B.n118 B.n117 585
R804 B.n116 B.n115 585
R805 B.n114 B.n113 585
R806 B.n112 B.n111 585
R807 B.n110 B.n109 585
R808 B.n108 B.n107 585
R809 B.n106 B.n105 585
R810 B.n104 B.n103 585
R811 B.n102 B.n101 585
R812 B.n53 B.n52 585
R813 B.n643 B.n54 585
R814 B.n647 B.n54 585
R815 B.n642 B.n641 585
R816 B.n641 B.n50 585
R817 B.n640 B.n49 585
R818 B.n653 B.n49 585
R819 B.n639 B.n48 585
R820 B.n654 B.n48 585
R821 B.n638 B.n47 585
R822 B.n655 B.n47 585
R823 B.n637 B.n636 585
R824 B.n636 B.n46 585
R825 B.n635 B.n42 585
R826 B.n661 B.n42 585
R827 B.n634 B.n41 585
R828 B.n662 B.n41 585
R829 B.n633 B.n40 585
R830 B.n663 B.n40 585
R831 B.n632 B.n631 585
R832 B.n631 B.n36 585
R833 B.n630 B.n35 585
R834 B.n669 B.n35 585
R835 B.n629 B.n34 585
R836 B.n670 B.n34 585
R837 B.n628 B.n33 585
R838 B.n671 B.n33 585
R839 B.n627 B.n626 585
R840 B.n626 B.n29 585
R841 B.n625 B.n28 585
R842 B.n677 B.n28 585
R843 B.n624 B.n27 585
R844 B.n678 B.n27 585
R845 B.n623 B.n26 585
R846 B.n679 B.n26 585
R847 B.n622 B.n621 585
R848 B.n621 B.n22 585
R849 B.n620 B.n21 585
R850 B.n685 B.n21 585
R851 B.n619 B.n20 585
R852 B.n686 B.n20 585
R853 B.n618 B.n19 585
R854 B.n687 B.n19 585
R855 B.n617 B.n616 585
R856 B.n616 B.n15 585
R857 B.n615 B.n14 585
R858 B.n693 B.n14 585
R859 B.n614 B.n13 585
R860 B.n694 B.n13 585
R861 B.n613 B.n12 585
R862 B.n695 B.n12 585
R863 B.n612 B.n611 585
R864 B.n611 B.n610 585
R865 B.n609 B.n608 585
R866 B.n609 B.n8 585
R867 B.n607 B.n7 585
R868 B.n702 B.n7 585
R869 B.n606 B.n6 585
R870 B.n703 B.n6 585
R871 B.n605 B.n5 585
R872 B.n704 B.n5 585
R873 B.n604 B.n603 585
R874 B.n603 B.n4 585
R875 B.n602 B.n259 585
R876 B.n602 B.n601 585
R877 B.n592 B.n260 585
R878 B.n261 B.n260 585
R879 B.n594 B.n593 585
R880 B.n595 B.n594 585
R881 B.n591 B.n266 585
R882 B.n266 B.n265 585
R883 B.n590 B.n589 585
R884 B.n589 B.n588 585
R885 B.n268 B.n267 585
R886 B.n269 B.n268 585
R887 B.n581 B.n580 585
R888 B.n582 B.n581 585
R889 B.n579 B.n274 585
R890 B.n274 B.n273 585
R891 B.n578 B.n577 585
R892 B.n577 B.n576 585
R893 B.n276 B.n275 585
R894 B.n277 B.n276 585
R895 B.n569 B.n568 585
R896 B.n570 B.n569 585
R897 B.n567 B.n282 585
R898 B.n282 B.n281 585
R899 B.n566 B.n565 585
R900 B.n565 B.n564 585
R901 B.n284 B.n283 585
R902 B.n285 B.n284 585
R903 B.n557 B.n556 585
R904 B.n558 B.n557 585
R905 B.n555 B.n290 585
R906 B.n290 B.n289 585
R907 B.n554 B.n553 585
R908 B.n553 B.n552 585
R909 B.n292 B.n291 585
R910 B.n293 B.n292 585
R911 B.n545 B.n544 585
R912 B.n546 B.n545 585
R913 B.n543 B.n298 585
R914 B.n298 B.n297 585
R915 B.n542 B.n541 585
R916 B.n541 B.n540 585
R917 B.n300 B.n299 585
R918 B.n533 B.n300 585
R919 B.n532 B.n531 585
R920 B.n534 B.n532 585
R921 B.n530 B.n305 585
R922 B.n305 B.n304 585
R923 B.n529 B.n528 585
R924 B.n528 B.n527 585
R925 B.n307 B.n306 585
R926 B.n308 B.n307 585
R927 B.n520 B.n519 585
R928 B.n521 B.n520 585
R929 B.n311 B.n310 585
R930 B.n359 B.n357 585
R931 B.n360 B.n356 585
R932 B.n360 B.n312 585
R933 B.n363 B.n362 585
R934 B.n364 B.n355 585
R935 B.n366 B.n365 585
R936 B.n368 B.n354 585
R937 B.n371 B.n370 585
R938 B.n372 B.n353 585
R939 B.n374 B.n373 585
R940 B.n376 B.n352 585
R941 B.n379 B.n378 585
R942 B.n380 B.n351 585
R943 B.n382 B.n381 585
R944 B.n384 B.n350 585
R945 B.n387 B.n386 585
R946 B.n388 B.n349 585
R947 B.n390 B.n389 585
R948 B.n392 B.n348 585
R949 B.n395 B.n394 585
R950 B.n396 B.n347 585
R951 B.n398 B.n397 585
R952 B.n400 B.n346 585
R953 B.n403 B.n402 585
R954 B.n404 B.n345 585
R955 B.n406 B.n405 585
R956 B.n408 B.n344 585
R957 B.n411 B.n410 585
R958 B.n412 B.n343 585
R959 B.n414 B.n413 585
R960 B.n416 B.n342 585
R961 B.n419 B.n418 585
R962 B.n420 B.n341 585
R963 B.n422 B.n421 585
R964 B.n424 B.n340 585
R965 B.n427 B.n426 585
R966 B.n429 B.n337 585
R967 B.n431 B.n430 585
R968 B.n433 B.n336 585
R969 B.n436 B.n435 585
R970 B.n437 B.n335 585
R971 B.n439 B.n438 585
R972 B.n441 B.n334 585
R973 B.n444 B.n443 585
R974 B.n445 B.n331 585
R975 B.n448 B.n447 585
R976 B.n450 B.n330 585
R977 B.n453 B.n452 585
R978 B.n454 B.n329 585
R979 B.n456 B.n455 585
R980 B.n458 B.n328 585
R981 B.n461 B.n460 585
R982 B.n462 B.n327 585
R983 B.n464 B.n463 585
R984 B.n466 B.n326 585
R985 B.n469 B.n468 585
R986 B.n470 B.n325 585
R987 B.n472 B.n471 585
R988 B.n474 B.n324 585
R989 B.n477 B.n476 585
R990 B.n478 B.n323 585
R991 B.n480 B.n479 585
R992 B.n482 B.n322 585
R993 B.n485 B.n484 585
R994 B.n486 B.n321 585
R995 B.n488 B.n487 585
R996 B.n490 B.n320 585
R997 B.n493 B.n492 585
R998 B.n494 B.n319 585
R999 B.n496 B.n495 585
R1000 B.n498 B.n318 585
R1001 B.n501 B.n500 585
R1002 B.n502 B.n317 585
R1003 B.n504 B.n503 585
R1004 B.n506 B.n316 585
R1005 B.n509 B.n508 585
R1006 B.n510 B.n315 585
R1007 B.n512 B.n511 585
R1008 B.n514 B.n314 585
R1009 B.n517 B.n516 585
R1010 B.n518 B.n313 585
R1011 B.n523 B.n522 585
R1012 B.n522 B.n521 585
R1013 B.n524 B.n309 585
R1014 B.n309 B.n308 585
R1015 B.n526 B.n525 585
R1016 B.n527 B.n526 585
R1017 B.n303 B.n302 585
R1018 B.n304 B.n303 585
R1019 B.n536 B.n535 585
R1020 B.n535 B.n534 585
R1021 B.n537 B.n301 585
R1022 B.n533 B.n301 585
R1023 B.n539 B.n538 585
R1024 B.n540 B.n539 585
R1025 B.n296 B.n295 585
R1026 B.n297 B.n296 585
R1027 B.n548 B.n547 585
R1028 B.n547 B.n546 585
R1029 B.n549 B.n294 585
R1030 B.n294 B.n293 585
R1031 B.n551 B.n550 585
R1032 B.n552 B.n551 585
R1033 B.n288 B.n287 585
R1034 B.n289 B.n288 585
R1035 B.n560 B.n559 585
R1036 B.n559 B.n558 585
R1037 B.n561 B.n286 585
R1038 B.n286 B.n285 585
R1039 B.n563 B.n562 585
R1040 B.n564 B.n563 585
R1041 B.n280 B.n279 585
R1042 B.n281 B.n280 585
R1043 B.n572 B.n571 585
R1044 B.n571 B.n570 585
R1045 B.n573 B.n278 585
R1046 B.n278 B.n277 585
R1047 B.n575 B.n574 585
R1048 B.n576 B.n575 585
R1049 B.n272 B.n271 585
R1050 B.n273 B.n272 585
R1051 B.n584 B.n583 585
R1052 B.n583 B.n582 585
R1053 B.n585 B.n270 585
R1054 B.n270 B.n269 585
R1055 B.n587 B.n586 585
R1056 B.n588 B.n587 585
R1057 B.n264 B.n263 585
R1058 B.n265 B.n264 585
R1059 B.n597 B.n596 585
R1060 B.n596 B.n595 585
R1061 B.n598 B.n262 585
R1062 B.n262 B.n261 585
R1063 B.n600 B.n599 585
R1064 B.n601 B.n600 585
R1065 B.n3 B.n0 585
R1066 B.n4 B.n3 585
R1067 B.n701 B.n1 585
R1068 B.n702 B.n701 585
R1069 B.n700 B.n699 585
R1070 B.n700 B.n8 585
R1071 B.n698 B.n9 585
R1072 B.n610 B.n9 585
R1073 B.n697 B.n696 585
R1074 B.n696 B.n695 585
R1075 B.n11 B.n10 585
R1076 B.n694 B.n11 585
R1077 B.n692 B.n691 585
R1078 B.n693 B.n692 585
R1079 B.n690 B.n16 585
R1080 B.n16 B.n15 585
R1081 B.n689 B.n688 585
R1082 B.n688 B.n687 585
R1083 B.n18 B.n17 585
R1084 B.n686 B.n18 585
R1085 B.n684 B.n683 585
R1086 B.n685 B.n684 585
R1087 B.n682 B.n23 585
R1088 B.n23 B.n22 585
R1089 B.n681 B.n680 585
R1090 B.n680 B.n679 585
R1091 B.n25 B.n24 585
R1092 B.n678 B.n25 585
R1093 B.n676 B.n675 585
R1094 B.n677 B.n676 585
R1095 B.n674 B.n30 585
R1096 B.n30 B.n29 585
R1097 B.n673 B.n672 585
R1098 B.n672 B.n671 585
R1099 B.n32 B.n31 585
R1100 B.n670 B.n32 585
R1101 B.n668 B.n667 585
R1102 B.n669 B.n668 585
R1103 B.n666 B.n37 585
R1104 B.n37 B.n36 585
R1105 B.n665 B.n664 585
R1106 B.n664 B.n663 585
R1107 B.n39 B.n38 585
R1108 B.n662 B.n39 585
R1109 B.n660 B.n659 585
R1110 B.n661 B.n660 585
R1111 B.n658 B.n43 585
R1112 B.n46 B.n43 585
R1113 B.n657 B.n656 585
R1114 B.n656 B.n655 585
R1115 B.n45 B.n44 585
R1116 B.n654 B.n45 585
R1117 B.n652 B.n651 585
R1118 B.n653 B.n652 585
R1119 B.n650 B.n51 585
R1120 B.n51 B.n50 585
R1121 B.n649 B.n648 585
R1122 B.n648 B.n647 585
R1123 B.n705 B.n704 585
R1124 B.n703 B.n2 585
R1125 B.n648 B.n53 468.476
R1126 B.n645 B.n54 468.476
R1127 B.n520 B.n313 468.476
R1128 B.n522 B.n311 468.476
R1129 B.n98 B.t19 431.861
R1130 B.n96 B.t8 431.861
R1131 B.n332 B.t16 431.861
R1132 B.n338 B.t12 431.861
R1133 B.n96 B.t10 273.635
R1134 B.n332 B.t18 273.635
R1135 B.n98 B.t20 273.635
R1136 B.n338 B.t15 273.635
R1137 B.n646 B.n94 256.663
R1138 B.n646 B.n93 256.663
R1139 B.n646 B.n92 256.663
R1140 B.n646 B.n91 256.663
R1141 B.n646 B.n90 256.663
R1142 B.n646 B.n89 256.663
R1143 B.n646 B.n88 256.663
R1144 B.n646 B.n87 256.663
R1145 B.n646 B.n86 256.663
R1146 B.n646 B.n85 256.663
R1147 B.n646 B.n84 256.663
R1148 B.n646 B.n83 256.663
R1149 B.n646 B.n82 256.663
R1150 B.n646 B.n81 256.663
R1151 B.n646 B.n80 256.663
R1152 B.n646 B.n79 256.663
R1153 B.n646 B.n78 256.663
R1154 B.n646 B.n77 256.663
R1155 B.n646 B.n76 256.663
R1156 B.n646 B.n75 256.663
R1157 B.n646 B.n74 256.663
R1158 B.n646 B.n73 256.663
R1159 B.n646 B.n72 256.663
R1160 B.n646 B.n71 256.663
R1161 B.n646 B.n70 256.663
R1162 B.n646 B.n69 256.663
R1163 B.n646 B.n68 256.663
R1164 B.n646 B.n67 256.663
R1165 B.n646 B.n66 256.663
R1166 B.n646 B.n65 256.663
R1167 B.n646 B.n64 256.663
R1168 B.n646 B.n63 256.663
R1169 B.n646 B.n62 256.663
R1170 B.n646 B.n61 256.663
R1171 B.n646 B.n60 256.663
R1172 B.n646 B.n59 256.663
R1173 B.n646 B.n58 256.663
R1174 B.n646 B.n57 256.663
R1175 B.n646 B.n56 256.663
R1176 B.n646 B.n55 256.663
R1177 B.n358 B.n312 256.663
R1178 B.n361 B.n312 256.663
R1179 B.n367 B.n312 256.663
R1180 B.n369 B.n312 256.663
R1181 B.n375 B.n312 256.663
R1182 B.n377 B.n312 256.663
R1183 B.n383 B.n312 256.663
R1184 B.n385 B.n312 256.663
R1185 B.n391 B.n312 256.663
R1186 B.n393 B.n312 256.663
R1187 B.n399 B.n312 256.663
R1188 B.n401 B.n312 256.663
R1189 B.n407 B.n312 256.663
R1190 B.n409 B.n312 256.663
R1191 B.n415 B.n312 256.663
R1192 B.n417 B.n312 256.663
R1193 B.n423 B.n312 256.663
R1194 B.n425 B.n312 256.663
R1195 B.n432 B.n312 256.663
R1196 B.n434 B.n312 256.663
R1197 B.n440 B.n312 256.663
R1198 B.n442 B.n312 256.663
R1199 B.n449 B.n312 256.663
R1200 B.n451 B.n312 256.663
R1201 B.n457 B.n312 256.663
R1202 B.n459 B.n312 256.663
R1203 B.n465 B.n312 256.663
R1204 B.n467 B.n312 256.663
R1205 B.n473 B.n312 256.663
R1206 B.n475 B.n312 256.663
R1207 B.n481 B.n312 256.663
R1208 B.n483 B.n312 256.663
R1209 B.n489 B.n312 256.663
R1210 B.n491 B.n312 256.663
R1211 B.n497 B.n312 256.663
R1212 B.n499 B.n312 256.663
R1213 B.n505 B.n312 256.663
R1214 B.n507 B.n312 256.663
R1215 B.n513 B.n312 256.663
R1216 B.n515 B.n312 256.663
R1217 B.n707 B.n706 256.663
R1218 B.n97 B.t11 246.871
R1219 B.n333 B.t17 246.871
R1220 B.n99 B.t21 246.871
R1221 B.n339 B.t14 246.871
R1222 B.n103 B.n102 163.367
R1223 B.n107 B.n106 163.367
R1224 B.n111 B.n110 163.367
R1225 B.n115 B.n114 163.367
R1226 B.n119 B.n118 163.367
R1227 B.n123 B.n122 163.367
R1228 B.n127 B.n126 163.367
R1229 B.n131 B.n130 163.367
R1230 B.n135 B.n134 163.367
R1231 B.n139 B.n138 163.367
R1232 B.n143 B.n142 163.367
R1233 B.n147 B.n146 163.367
R1234 B.n151 B.n150 163.367
R1235 B.n155 B.n154 163.367
R1236 B.n159 B.n158 163.367
R1237 B.n163 B.n162 163.367
R1238 B.n167 B.n166 163.367
R1239 B.n171 B.n170 163.367
R1240 B.n175 B.n174 163.367
R1241 B.n179 B.n178 163.367
R1242 B.n183 B.n182 163.367
R1243 B.n187 B.n186 163.367
R1244 B.n192 B.n191 163.367
R1245 B.n196 B.n195 163.367
R1246 B.n200 B.n199 163.367
R1247 B.n204 B.n203 163.367
R1248 B.n208 B.n207 163.367
R1249 B.n212 B.n211 163.367
R1250 B.n216 B.n215 163.367
R1251 B.n220 B.n219 163.367
R1252 B.n224 B.n223 163.367
R1253 B.n228 B.n227 163.367
R1254 B.n232 B.n231 163.367
R1255 B.n236 B.n235 163.367
R1256 B.n240 B.n239 163.367
R1257 B.n244 B.n243 163.367
R1258 B.n248 B.n247 163.367
R1259 B.n252 B.n251 163.367
R1260 B.n256 B.n255 163.367
R1261 B.n645 B.n95 163.367
R1262 B.n520 B.n307 163.367
R1263 B.n528 B.n307 163.367
R1264 B.n528 B.n305 163.367
R1265 B.n532 B.n305 163.367
R1266 B.n532 B.n300 163.367
R1267 B.n541 B.n300 163.367
R1268 B.n541 B.n298 163.367
R1269 B.n545 B.n298 163.367
R1270 B.n545 B.n292 163.367
R1271 B.n553 B.n292 163.367
R1272 B.n553 B.n290 163.367
R1273 B.n557 B.n290 163.367
R1274 B.n557 B.n284 163.367
R1275 B.n565 B.n284 163.367
R1276 B.n565 B.n282 163.367
R1277 B.n569 B.n282 163.367
R1278 B.n569 B.n276 163.367
R1279 B.n577 B.n276 163.367
R1280 B.n577 B.n274 163.367
R1281 B.n581 B.n274 163.367
R1282 B.n581 B.n268 163.367
R1283 B.n589 B.n268 163.367
R1284 B.n589 B.n266 163.367
R1285 B.n594 B.n266 163.367
R1286 B.n594 B.n260 163.367
R1287 B.n602 B.n260 163.367
R1288 B.n603 B.n602 163.367
R1289 B.n603 B.n5 163.367
R1290 B.n6 B.n5 163.367
R1291 B.n7 B.n6 163.367
R1292 B.n609 B.n7 163.367
R1293 B.n611 B.n609 163.367
R1294 B.n611 B.n12 163.367
R1295 B.n13 B.n12 163.367
R1296 B.n14 B.n13 163.367
R1297 B.n616 B.n14 163.367
R1298 B.n616 B.n19 163.367
R1299 B.n20 B.n19 163.367
R1300 B.n21 B.n20 163.367
R1301 B.n621 B.n21 163.367
R1302 B.n621 B.n26 163.367
R1303 B.n27 B.n26 163.367
R1304 B.n28 B.n27 163.367
R1305 B.n626 B.n28 163.367
R1306 B.n626 B.n33 163.367
R1307 B.n34 B.n33 163.367
R1308 B.n35 B.n34 163.367
R1309 B.n631 B.n35 163.367
R1310 B.n631 B.n40 163.367
R1311 B.n41 B.n40 163.367
R1312 B.n42 B.n41 163.367
R1313 B.n636 B.n42 163.367
R1314 B.n636 B.n47 163.367
R1315 B.n48 B.n47 163.367
R1316 B.n49 B.n48 163.367
R1317 B.n641 B.n49 163.367
R1318 B.n641 B.n54 163.367
R1319 B.n360 B.n359 163.367
R1320 B.n362 B.n360 163.367
R1321 B.n366 B.n355 163.367
R1322 B.n370 B.n368 163.367
R1323 B.n374 B.n353 163.367
R1324 B.n378 B.n376 163.367
R1325 B.n382 B.n351 163.367
R1326 B.n386 B.n384 163.367
R1327 B.n390 B.n349 163.367
R1328 B.n394 B.n392 163.367
R1329 B.n398 B.n347 163.367
R1330 B.n402 B.n400 163.367
R1331 B.n406 B.n345 163.367
R1332 B.n410 B.n408 163.367
R1333 B.n414 B.n343 163.367
R1334 B.n418 B.n416 163.367
R1335 B.n422 B.n341 163.367
R1336 B.n426 B.n424 163.367
R1337 B.n431 B.n337 163.367
R1338 B.n435 B.n433 163.367
R1339 B.n439 B.n335 163.367
R1340 B.n443 B.n441 163.367
R1341 B.n448 B.n331 163.367
R1342 B.n452 B.n450 163.367
R1343 B.n456 B.n329 163.367
R1344 B.n460 B.n458 163.367
R1345 B.n464 B.n327 163.367
R1346 B.n468 B.n466 163.367
R1347 B.n472 B.n325 163.367
R1348 B.n476 B.n474 163.367
R1349 B.n480 B.n323 163.367
R1350 B.n484 B.n482 163.367
R1351 B.n488 B.n321 163.367
R1352 B.n492 B.n490 163.367
R1353 B.n496 B.n319 163.367
R1354 B.n500 B.n498 163.367
R1355 B.n504 B.n317 163.367
R1356 B.n508 B.n506 163.367
R1357 B.n512 B.n315 163.367
R1358 B.n516 B.n514 163.367
R1359 B.n522 B.n309 163.367
R1360 B.n526 B.n309 163.367
R1361 B.n526 B.n303 163.367
R1362 B.n535 B.n303 163.367
R1363 B.n535 B.n301 163.367
R1364 B.n539 B.n301 163.367
R1365 B.n539 B.n296 163.367
R1366 B.n547 B.n296 163.367
R1367 B.n547 B.n294 163.367
R1368 B.n551 B.n294 163.367
R1369 B.n551 B.n288 163.367
R1370 B.n559 B.n288 163.367
R1371 B.n559 B.n286 163.367
R1372 B.n563 B.n286 163.367
R1373 B.n563 B.n280 163.367
R1374 B.n571 B.n280 163.367
R1375 B.n571 B.n278 163.367
R1376 B.n575 B.n278 163.367
R1377 B.n575 B.n272 163.367
R1378 B.n583 B.n272 163.367
R1379 B.n583 B.n270 163.367
R1380 B.n587 B.n270 163.367
R1381 B.n587 B.n264 163.367
R1382 B.n596 B.n264 163.367
R1383 B.n596 B.n262 163.367
R1384 B.n600 B.n262 163.367
R1385 B.n600 B.n3 163.367
R1386 B.n705 B.n3 163.367
R1387 B.n701 B.n2 163.367
R1388 B.n701 B.n700 163.367
R1389 B.n700 B.n9 163.367
R1390 B.n696 B.n9 163.367
R1391 B.n696 B.n11 163.367
R1392 B.n692 B.n11 163.367
R1393 B.n692 B.n16 163.367
R1394 B.n688 B.n16 163.367
R1395 B.n688 B.n18 163.367
R1396 B.n684 B.n18 163.367
R1397 B.n684 B.n23 163.367
R1398 B.n680 B.n23 163.367
R1399 B.n680 B.n25 163.367
R1400 B.n676 B.n25 163.367
R1401 B.n676 B.n30 163.367
R1402 B.n672 B.n30 163.367
R1403 B.n672 B.n32 163.367
R1404 B.n668 B.n32 163.367
R1405 B.n668 B.n37 163.367
R1406 B.n664 B.n37 163.367
R1407 B.n664 B.n39 163.367
R1408 B.n660 B.n39 163.367
R1409 B.n660 B.n43 163.367
R1410 B.n656 B.n43 163.367
R1411 B.n656 B.n45 163.367
R1412 B.n652 B.n45 163.367
R1413 B.n652 B.n51 163.367
R1414 B.n648 B.n51 163.367
R1415 B.n521 B.n312 84.477
R1416 B.n647 B.n646 84.477
R1417 B.n55 B.n53 71.676
R1418 B.n103 B.n56 71.676
R1419 B.n107 B.n57 71.676
R1420 B.n111 B.n58 71.676
R1421 B.n115 B.n59 71.676
R1422 B.n119 B.n60 71.676
R1423 B.n123 B.n61 71.676
R1424 B.n127 B.n62 71.676
R1425 B.n131 B.n63 71.676
R1426 B.n135 B.n64 71.676
R1427 B.n139 B.n65 71.676
R1428 B.n143 B.n66 71.676
R1429 B.n147 B.n67 71.676
R1430 B.n151 B.n68 71.676
R1431 B.n155 B.n69 71.676
R1432 B.n159 B.n70 71.676
R1433 B.n163 B.n71 71.676
R1434 B.n167 B.n72 71.676
R1435 B.n171 B.n73 71.676
R1436 B.n175 B.n74 71.676
R1437 B.n179 B.n75 71.676
R1438 B.n183 B.n76 71.676
R1439 B.n187 B.n77 71.676
R1440 B.n192 B.n78 71.676
R1441 B.n196 B.n79 71.676
R1442 B.n200 B.n80 71.676
R1443 B.n204 B.n81 71.676
R1444 B.n208 B.n82 71.676
R1445 B.n212 B.n83 71.676
R1446 B.n216 B.n84 71.676
R1447 B.n220 B.n85 71.676
R1448 B.n224 B.n86 71.676
R1449 B.n228 B.n87 71.676
R1450 B.n232 B.n88 71.676
R1451 B.n236 B.n89 71.676
R1452 B.n240 B.n90 71.676
R1453 B.n244 B.n91 71.676
R1454 B.n248 B.n92 71.676
R1455 B.n252 B.n93 71.676
R1456 B.n256 B.n94 71.676
R1457 B.n95 B.n94 71.676
R1458 B.n255 B.n93 71.676
R1459 B.n251 B.n92 71.676
R1460 B.n247 B.n91 71.676
R1461 B.n243 B.n90 71.676
R1462 B.n239 B.n89 71.676
R1463 B.n235 B.n88 71.676
R1464 B.n231 B.n87 71.676
R1465 B.n227 B.n86 71.676
R1466 B.n223 B.n85 71.676
R1467 B.n219 B.n84 71.676
R1468 B.n215 B.n83 71.676
R1469 B.n211 B.n82 71.676
R1470 B.n207 B.n81 71.676
R1471 B.n203 B.n80 71.676
R1472 B.n199 B.n79 71.676
R1473 B.n195 B.n78 71.676
R1474 B.n191 B.n77 71.676
R1475 B.n186 B.n76 71.676
R1476 B.n182 B.n75 71.676
R1477 B.n178 B.n74 71.676
R1478 B.n174 B.n73 71.676
R1479 B.n170 B.n72 71.676
R1480 B.n166 B.n71 71.676
R1481 B.n162 B.n70 71.676
R1482 B.n158 B.n69 71.676
R1483 B.n154 B.n68 71.676
R1484 B.n150 B.n67 71.676
R1485 B.n146 B.n66 71.676
R1486 B.n142 B.n65 71.676
R1487 B.n138 B.n64 71.676
R1488 B.n134 B.n63 71.676
R1489 B.n130 B.n62 71.676
R1490 B.n126 B.n61 71.676
R1491 B.n122 B.n60 71.676
R1492 B.n118 B.n59 71.676
R1493 B.n114 B.n58 71.676
R1494 B.n110 B.n57 71.676
R1495 B.n106 B.n56 71.676
R1496 B.n102 B.n55 71.676
R1497 B.n358 B.n311 71.676
R1498 B.n362 B.n361 71.676
R1499 B.n367 B.n366 71.676
R1500 B.n370 B.n369 71.676
R1501 B.n375 B.n374 71.676
R1502 B.n378 B.n377 71.676
R1503 B.n383 B.n382 71.676
R1504 B.n386 B.n385 71.676
R1505 B.n391 B.n390 71.676
R1506 B.n394 B.n393 71.676
R1507 B.n399 B.n398 71.676
R1508 B.n402 B.n401 71.676
R1509 B.n407 B.n406 71.676
R1510 B.n410 B.n409 71.676
R1511 B.n415 B.n414 71.676
R1512 B.n418 B.n417 71.676
R1513 B.n423 B.n422 71.676
R1514 B.n426 B.n425 71.676
R1515 B.n432 B.n431 71.676
R1516 B.n435 B.n434 71.676
R1517 B.n440 B.n439 71.676
R1518 B.n443 B.n442 71.676
R1519 B.n449 B.n448 71.676
R1520 B.n452 B.n451 71.676
R1521 B.n457 B.n456 71.676
R1522 B.n460 B.n459 71.676
R1523 B.n465 B.n464 71.676
R1524 B.n468 B.n467 71.676
R1525 B.n473 B.n472 71.676
R1526 B.n476 B.n475 71.676
R1527 B.n481 B.n480 71.676
R1528 B.n484 B.n483 71.676
R1529 B.n489 B.n488 71.676
R1530 B.n492 B.n491 71.676
R1531 B.n497 B.n496 71.676
R1532 B.n500 B.n499 71.676
R1533 B.n505 B.n504 71.676
R1534 B.n508 B.n507 71.676
R1535 B.n513 B.n512 71.676
R1536 B.n516 B.n515 71.676
R1537 B.n359 B.n358 71.676
R1538 B.n361 B.n355 71.676
R1539 B.n368 B.n367 71.676
R1540 B.n369 B.n353 71.676
R1541 B.n376 B.n375 71.676
R1542 B.n377 B.n351 71.676
R1543 B.n384 B.n383 71.676
R1544 B.n385 B.n349 71.676
R1545 B.n392 B.n391 71.676
R1546 B.n393 B.n347 71.676
R1547 B.n400 B.n399 71.676
R1548 B.n401 B.n345 71.676
R1549 B.n408 B.n407 71.676
R1550 B.n409 B.n343 71.676
R1551 B.n416 B.n415 71.676
R1552 B.n417 B.n341 71.676
R1553 B.n424 B.n423 71.676
R1554 B.n425 B.n337 71.676
R1555 B.n433 B.n432 71.676
R1556 B.n434 B.n335 71.676
R1557 B.n441 B.n440 71.676
R1558 B.n442 B.n331 71.676
R1559 B.n450 B.n449 71.676
R1560 B.n451 B.n329 71.676
R1561 B.n458 B.n457 71.676
R1562 B.n459 B.n327 71.676
R1563 B.n466 B.n465 71.676
R1564 B.n467 B.n325 71.676
R1565 B.n474 B.n473 71.676
R1566 B.n475 B.n323 71.676
R1567 B.n482 B.n481 71.676
R1568 B.n483 B.n321 71.676
R1569 B.n490 B.n489 71.676
R1570 B.n491 B.n319 71.676
R1571 B.n498 B.n497 71.676
R1572 B.n499 B.n317 71.676
R1573 B.n506 B.n505 71.676
R1574 B.n507 B.n315 71.676
R1575 B.n514 B.n513 71.676
R1576 B.n515 B.n313 71.676
R1577 B.n706 B.n705 71.676
R1578 B.n706 B.n2 71.676
R1579 B.n100 B.n99 59.5399
R1580 B.n189 B.n97 59.5399
R1581 B.n446 B.n333 59.5399
R1582 B.n428 B.n339 59.5399
R1583 B.n521 B.n308 49.098
R1584 B.n527 B.n308 49.098
R1585 B.n527 B.n304 49.098
R1586 B.n534 B.n304 49.098
R1587 B.n534 B.n533 49.098
R1588 B.n540 B.n297 49.098
R1589 B.n546 B.n297 49.098
R1590 B.n546 B.n293 49.098
R1591 B.n552 B.n293 49.098
R1592 B.n552 B.n289 49.098
R1593 B.n558 B.n289 49.098
R1594 B.n564 B.n285 49.098
R1595 B.n564 B.n281 49.098
R1596 B.n570 B.n281 49.098
R1597 B.n576 B.n277 49.098
R1598 B.n576 B.n273 49.098
R1599 B.n582 B.n273 49.098
R1600 B.n588 B.n269 49.098
R1601 B.n588 B.n265 49.098
R1602 B.n595 B.n265 49.098
R1603 B.n601 B.n261 49.098
R1604 B.n601 B.n4 49.098
R1605 B.n704 B.n4 49.098
R1606 B.n704 B.n703 49.098
R1607 B.n703 B.n702 49.098
R1608 B.n702 B.n8 49.098
R1609 B.n610 B.n8 49.098
R1610 B.n695 B.n694 49.098
R1611 B.n694 B.n693 49.098
R1612 B.n693 B.n15 49.098
R1613 B.n687 B.n686 49.098
R1614 B.n686 B.n685 49.098
R1615 B.n685 B.n22 49.098
R1616 B.n679 B.n678 49.098
R1617 B.n678 B.n677 49.098
R1618 B.n677 B.n29 49.098
R1619 B.n671 B.n670 49.098
R1620 B.n670 B.n669 49.098
R1621 B.n669 B.n36 49.098
R1622 B.n663 B.n36 49.098
R1623 B.n663 B.n662 49.098
R1624 B.n662 B.n661 49.098
R1625 B.n655 B.n46 49.098
R1626 B.n655 B.n654 49.098
R1627 B.n654 B.n653 49.098
R1628 B.n653 B.n50 49.098
R1629 B.n647 B.n50 49.098
R1630 B.n595 B.t4 42.5998
R1631 B.n695 B.t2 42.5998
R1632 B.n582 B.t5 39.7117
R1633 B.n687 B.t6 39.7117
R1634 B.n570 B.t1 36.8236
R1635 B.n679 B.t7 36.8236
R1636 B.n558 B.t3 33.9355
R1637 B.n671 B.t0 33.9355
R1638 B.n523 B.n310 30.4395
R1639 B.n519 B.n518 30.4395
R1640 B.n644 B.n643 30.4395
R1641 B.n649 B.n52 30.4395
R1642 B.n540 B.t13 28.1593
R1643 B.n661 B.t9 28.1593
R1644 B.n99 B.n98 26.7641
R1645 B.n97 B.n96 26.7641
R1646 B.n333 B.n332 26.7641
R1647 B.n339 B.n338 26.7641
R1648 B.n533 B.t13 20.9391
R1649 B.n46 B.t9 20.9391
R1650 B B.n707 18.0485
R1651 B.t3 B.n285 15.163
R1652 B.t0 B.n29 15.163
R1653 B.t1 B.n277 12.2749
R1654 B.t7 B.n22 12.2749
R1655 B.n524 B.n523 10.6151
R1656 B.n525 B.n524 10.6151
R1657 B.n525 B.n302 10.6151
R1658 B.n536 B.n302 10.6151
R1659 B.n537 B.n536 10.6151
R1660 B.n538 B.n537 10.6151
R1661 B.n538 B.n295 10.6151
R1662 B.n548 B.n295 10.6151
R1663 B.n549 B.n548 10.6151
R1664 B.n550 B.n549 10.6151
R1665 B.n550 B.n287 10.6151
R1666 B.n560 B.n287 10.6151
R1667 B.n561 B.n560 10.6151
R1668 B.n562 B.n561 10.6151
R1669 B.n562 B.n279 10.6151
R1670 B.n572 B.n279 10.6151
R1671 B.n573 B.n572 10.6151
R1672 B.n574 B.n573 10.6151
R1673 B.n574 B.n271 10.6151
R1674 B.n584 B.n271 10.6151
R1675 B.n585 B.n584 10.6151
R1676 B.n586 B.n585 10.6151
R1677 B.n586 B.n263 10.6151
R1678 B.n597 B.n263 10.6151
R1679 B.n598 B.n597 10.6151
R1680 B.n599 B.n598 10.6151
R1681 B.n599 B.n0 10.6151
R1682 B.n357 B.n310 10.6151
R1683 B.n357 B.n356 10.6151
R1684 B.n363 B.n356 10.6151
R1685 B.n364 B.n363 10.6151
R1686 B.n365 B.n364 10.6151
R1687 B.n365 B.n354 10.6151
R1688 B.n371 B.n354 10.6151
R1689 B.n372 B.n371 10.6151
R1690 B.n373 B.n372 10.6151
R1691 B.n373 B.n352 10.6151
R1692 B.n379 B.n352 10.6151
R1693 B.n380 B.n379 10.6151
R1694 B.n381 B.n380 10.6151
R1695 B.n381 B.n350 10.6151
R1696 B.n387 B.n350 10.6151
R1697 B.n388 B.n387 10.6151
R1698 B.n389 B.n388 10.6151
R1699 B.n389 B.n348 10.6151
R1700 B.n395 B.n348 10.6151
R1701 B.n396 B.n395 10.6151
R1702 B.n397 B.n396 10.6151
R1703 B.n397 B.n346 10.6151
R1704 B.n403 B.n346 10.6151
R1705 B.n404 B.n403 10.6151
R1706 B.n405 B.n404 10.6151
R1707 B.n405 B.n344 10.6151
R1708 B.n411 B.n344 10.6151
R1709 B.n412 B.n411 10.6151
R1710 B.n413 B.n412 10.6151
R1711 B.n413 B.n342 10.6151
R1712 B.n419 B.n342 10.6151
R1713 B.n420 B.n419 10.6151
R1714 B.n421 B.n420 10.6151
R1715 B.n421 B.n340 10.6151
R1716 B.n427 B.n340 10.6151
R1717 B.n430 B.n429 10.6151
R1718 B.n430 B.n336 10.6151
R1719 B.n436 B.n336 10.6151
R1720 B.n437 B.n436 10.6151
R1721 B.n438 B.n437 10.6151
R1722 B.n438 B.n334 10.6151
R1723 B.n444 B.n334 10.6151
R1724 B.n445 B.n444 10.6151
R1725 B.n447 B.n330 10.6151
R1726 B.n453 B.n330 10.6151
R1727 B.n454 B.n453 10.6151
R1728 B.n455 B.n454 10.6151
R1729 B.n455 B.n328 10.6151
R1730 B.n461 B.n328 10.6151
R1731 B.n462 B.n461 10.6151
R1732 B.n463 B.n462 10.6151
R1733 B.n463 B.n326 10.6151
R1734 B.n469 B.n326 10.6151
R1735 B.n470 B.n469 10.6151
R1736 B.n471 B.n470 10.6151
R1737 B.n471 B.n324 10.6151
R1738 B.n477 B.n324 10.6151
R1739 B.n478 B.n477 10.6151
R1740 B.n479 B.n478 10.6151
R1741 B.n479 B.n322 10.6151
R1742 B.n485 B.n322 10.6151
R1743 B.n486 B.n485 10.6151
R1744 B.n487 B.n486 10.6151
R1745 B.n487 B.n320 10.6151
R1746 B.n493 B.n320 10.6151
R1747 B.n494 B.n493 10.6151
R1748 B.n495 B.n494 10.6151
R1749 B.n495 B.n318 10.6151
R1750 B.n501 B.n318 10.6151
R1751 B.n502 B.n501 10.6151
R1752 B.n503 B.n502 10.6151
R1753 B.n503 B.n316 10.6151
R1754 B.n509 B.n316 10.6151
R1755 B.n510 B.n509 10.6151
R1756 B.n511 B.n510 10.6151
R1757 B.n511 B.n314 10.6151
R1758 B.n517 B.n314 10.6151
R1759 B.n518 B.n517 10.6151
R1760 B.n519 B.n306 10.6151
R1761 B.n529 B.n306 10.6151
R1762 B.n530 B.n529 10.6151
R1763 B.n531 B.n530 10.6151
R1764 B.n531 B.n299 10.6151
R1765 B.n542 B.n299 10.6151
R1766 B.n543 B.n542 10.6151
R1767 B.n544 B.n543 10.6151
R1768 B.n544 B.n291 10.6151
R1769 B.n554 B.n291 10.6151
R1770 B.n555 B.n554 10.6151
R1771 B.n556 B.n555 10.6151
R1772 B.n556 B.n283 10.6151
R1773 B.n566 B.n283 10.6151
R1774 B.n567 B.n566 10.6151
R1775 B.n568 B.n567 10.6151
R1776 B.n568 B.n275 10.6151
R1777 B.n578 B.n275 10.6151
R1778 B.n579 B.n578 10.6151
R1779 B.n580 B.n579 10.6151
R1780 B.n580 B.n267 10.6151
R1781 B.n590 B.n267 10.6151
R1782 B.n591 B.n590 10.6151
R1783 B.n593 B.n591 10.6151
R1784 B.n593 B.n592 10.6151
R1785 B.n592 B.n259 10.6151
R1786 B.n604 B.n259 10.6151
R1787 B.n605 B.n604 10.6151
R1788 B.n606 B.n605 10.6151
R1789 B.n607 B.n606 10.6151
R1790 B.n608 B.n607 10.6151
R1791 B.n612 B.n608 10.6151
R1792 B.n613 B.n612 10.6151
R1793 B.n614 B.n613 10.6151
R1794 B.n615 B.n614 10.6151
R1795 B.n617 B.n615 10.6151
R1796 B.n618 B.n617 10.6151
R1797 B.n619 B.n618 10.6151
R1798 B.n620 B.n619 10.6151
R1799 B.n622 B.n620 10.6151
R1800 B.n623 B.n622 10.6151
R1801 B.n624 B.n623 10.6151
R1802 B.n625 B.n624 10.6151
R1803 B.n627 B.n625 10.6151
R1804 B.n628 B.n627 10.6151
R1805 B.n629 B.n628 10.6151
R1806 B.n630 B.n629 10.6151
R1807 B.n632 B.n630 10.6151
R1808 B.n633 B.n632 10.6151
R1809 B.n634 B.n633 10.6151
R1810 B.n635 B.n634 10.6151
R1811 B.n637 B.n635 10.6151
R1812 B.n638 B.n637 10.6151
R1813 B.n639 B.n638 10.6151
R1814 B.n640 B.n639 10.6151
R1815 B.n642 B.n640 10.6151
R1816 B.n643 B.n642 10.6151
R1817 B.n699 B.n1 10.6151
R1818 B.n699 B.n698 10.6151
R1819 B.n698 B.n697 10.6151
R1820 B.n697 B.n10 10.6151
R1821 B.n691 B.n10 10.6151
R1822 B.n691 B.n690 10.6151
R1823 B.n690 B.n689 10.6151
R1824 B.n689 B.n17 10.6151
R1825 B.n683 B.n17 10.6151
R1826 B.n683 B.n682 10.6151
R1827 B.n682 B.n681 10.6151
R1828 B.n681 B.n24 10.6151
R1829 B.n675 B.n24 10.6151
R1830 B.n675 B.n674 10.6151
R1831 B.n674 B.n673 10.6151
R1832 B.n673 B.n31 10.6151
R1833 B.n667 B.n31 10.6151
R1834 B.n667 B.n666 10.6151
R1835 B.n666 B.n665 10.6151
R1836 B.n665 B.n38 10.6151
R1837 B.n659 B.n38 10.6151
R1838 B.n659 B.n658 10.6151
R1839 B.n658 B.n657 10.6151
R1840 B.n657 B.n44 10.6151
R1841 B.n651 B.n44 10.6151
R1842 B.n651 B.n650 10.6151
R1843 B.n650 B.n649 10.6151
R1844 B.n101 B.n52 10.6151
R1845 B.n104 B.n101 10.6151
R1846 B.n105 B.n104 10.6151
R1847 B.n108 B.n105 10.6151
R1848 B.n109 B.n108 10.6151
R1849 B.n112 B.n109 10.6151
R1850 B.n113 B.n112 10.6151
R1851 B.n116 B.n113 10.6151
R1852 B.n117 B.n116 10.6151
R1853 B.n120 B.n117 10.6151
R1854 B.n121 B.n120 10.6151
R1855 B.n124 B.n121 10.6151
R1856 B.n125 B.n124 10.6151
R1857 B.n128 B.n125 10.6151
R1858 B.n129 B.n128 10.6151
R1859 B.n132 B.n129 10.6151
R1860 B.n133 B.n132 10.6151
R1861 B.n136 B.n133 10.6151
R1862 B.n137 B.n136 10.6151
R1863 B.n140 B.n137 10.6151
R1864 B.n141 B.n140 10.6151
R1865 B.n144 B.n141 10.6151
R1866 B.n145 B.n144 10.6151
R1867 B.n148 B.n145 10.6151
R1868 B.n149 B.n148 10.6151
R1869 B.n152 B.n149 10.6151
R1870 B.n153 B.n152 10.6151
R1871 B.n156 B.n153 10.6151
R1872 B.n157 B.n156 10.6151
R1873 B.n160 B.n157 10.6151
R1874 B.n161 B.n160 10.6151
R1875 B.n164 B.n161 10.6151
R1876 B.n165 B.n164 10.6151
R1877 B.n168 B.n165 10.6151
R1878 B.n169 B.n168 10.6151
R1879 B.n173 B.n172 10.6151
R1880 B.n176 B.n173 10.6151
R1881 B.n177 B.n176 10.6151
R1882 B.n180 B.n177 10.6151
R1883 B.n181 B.n180 10.6151
R1884 B.n184 B.n181 10.6151
R1885 B.n185 B.n184 10.6151
R1886 B.n188 B.n185 10.6151
R1887 B.n193 B.n190 10.6151
R1888 B.n194 B.n193 10.6151
R1889 B.n197 B.n194 10.6151
R1890 B.n198 B.n197 10.6151
R1891 B.n201 B.n198 10.6151
R1892 B.n202 B.n201 10.6151
R1893 B.n205 B.n202 10.6151
R1894 B.n206 B.n205 10.6151
R1895 B.n209 B.n206 10.6151
R1896 B.n210 B.n209 10.6151
R1897 B.n213 B.n210 10.6151
R1898 B.n214 B.n213 10.6151
R1899 B.n217 B.n214 10.6151
R1900 B.n218 B.n217 10.6151
R1901 B.n221 B.n218 10.6151
R1902 B.n222 B.n221 10.6151
R1903 B.n225 B.n222 10.6151
R1904 B.n226 B.n225 10.6151
R1905 B.n229 B.n226 10.6151
R1906 B.n230 B.n229 10.6151
R1907 B.n233 B.n230 10.6151
R1908 B.n234 B.n233 10.6151
R1909 B.n237 B.n234 10.6151
R1910 B.n238 B.n237 10.6151
R1911 B.n241 B.n238 10.6151
R1912 B.n242 B.n241 10.6151
R1913 B.n245 B.n242 10.6151
R1914 B.n246 B.n245 10.6151
R1915 B.n249 B.n246 10.6151
R1916 B.n250 B.n249 10.6151
R1917 B.n253 B.n250 10.6151
R1918 B.n254 B.n253 10.6151
R1919 B.n257 B.n254 10.6151
R1920 B.n258 B.n257 10.6151
R1921 B.n644 B.n258 10.6151
R1922 B.t5 B.n269 9.38678
R1923 B.t6 B.n15 9.38678
R1924 B.n707 B.n0 8.11757
R1925 B.n707 B.n1 8.11757
R1926 B.n429 B.n428 6.5566
R1927 B.n446 B.n445 6.5566
R1928 B.n172 B.n100 6.5566
R1929 B.n189 B.n188 6.5566
R1930 B.t4 B.n261 6.49869
R1931 B.n610 B.t2 6.49869
R1932 B.n428 B.n427 4.05904
R1933 B.n447 B.n446 4.05904
R1934 B.n169 B.n100 4.05904
R1935 B.n190 B.n189 4.05904
R1936 VP.n7 VP.t5 287.925
R1937 VP.n17 VP.t2 266.478
R1938 VP.n29 VP.t0 266.478
R1939 VP.n15 VP.t1 266.478
R1940 VP.n22 VP.t7 228.607
R1941 VP.n1 VP.t6 228.607
R1942 VP.n5 VP.t3 228.607
R1943 VP.n8 VP.t4 228.607
R1944 VP.n9 VP.n6 161.3
R1945 VP.n11 VP.n10 161.3
R1946 VP.n13 VP.n12 161.3
R1947 VP.n14 VP.n4 161.3
R1948 VP.n28 VP.n0 161.3
R1949 VP.n27 VP.n26 161.3
R1950 VP.n25 VP.n24 161.3
R1951 VP.n23 VP.n2 161.3
R1952 VP.n21 VP.n20 161.3
R1953 VP.n19 VP.n3 161.3
R1954 VP.n16 VP.n15 80.6037
R1955 VP.n30 VP.n29 80.6037
R1956 VP.n18 VP.n17 80.6037
R1957 VP.n24 VP.n23 56.4773
R1958 VP.n10 VP.n9 56.4773
R1959 VP.n17 VP.n3 43.0884
R1960 VP.n29 VP.n28 43.0884
R1961 VP.n15 VP.n14 43.0884
R1962 VP.n18 VP.n16 42.1908
R1963 VP.n8 VP.n7 35.3356
R1964 VP.n7 VP.n6 28.7542
R1965 VP.n21 VP.n3 27.752
R1966 VP.n28 VP.n27 27.752
R1967 VP.n14 VP.n13 27.752
R1968 VP.n23 VP.n22 21.4227
R1969 VP.n24 VP.n1 21.4227
R1970 VP.n10 VP.n5 21.4227
R1971 VP.n9 VP.n8 21.4227
R1972 VP.n22 VP.n21 2.92171
R1973 VP.n27 VP.n1 2.92171
R1974 VP.n13 VP.n5 2.92171
R1975 VP.n16 VP.n4 0.285035
R1976 VP.n19 VP.n18 0.285035
R1977 VP.n30 VP.n0 0.285035
R1978 VP.n11 VP.n6 0.189894
R1979 VP.n12 VP.n11 0.189894
R1980 VP.n12 VP.n4 0.189894
R1981 VP.n20 VP.n19 0.189894
R1982 VP.n20 VP.n2 0.189894
R1983 VP.n25 VP.n2 0.189894
R1984 VP.n26 VP.n25 0.189894
R1985 VP.n26 VP.n0 0.189894
R1986 VP VP.n30 0.146778
R1987 VDD1 VDD1.n0 63.2933
R1988 VDD1.n3 VDD1.n2 63.1796
R1989 VDD1.n3 VDD1.n1 63.1796
R1990 VDD1.n5 VDD1.n4 62.6402
R1991 VDD1.n5 VDD1.n3 38.238
R1992 VDD1.n4 VDD1.t4 1.98845
R1993 VDD1.n4 VDD1.t6 1.98845
R1994 VDD1.n0 VDD1.t2 1.98845
R1995 VDD1.n0 VDD1.t3 1.98845
R1996 VDD1.n2 VDD1.t1 1.98845
R1997 VDD1.n2 VDD1.t7 1.98845
R1998 VDD1.n1 VDD1.t5 1.98845
R1999 VDD1.n1 VDD1.t0 1.98845
R2000 VDD1 VDD1.n5 0.537138
C0 VDD2 VDD1 1.00035f
C1 VN VTAIL 5.55449f
C2 VDD2 VN 5.58263f
C3 VDD1 VP 5.78783f
C4 VN VP 5.39585f
C5 VDD2 VTAIL 8.26759f
C6 VDD1 VN 0.148506f
C7 VP VTAIL 5.56859f
C8 VDD2 VP 0.354314f
C9 VDD1 VTAIL 8.22356f
C10 VDD2 B 3.669084f
C11 VDD1 B 3.93857f
C12 VTAIL B 8.105109f
C13 VN B 9.58845f
C14 VP B 7.888441f
C15 VDD1.t2 B 0.203322f
C16 VDD1.t3 B 0.203322f
C17 VDD1.n0 B 1.79361f
C18 VDD1.t5 B 0.203322f
C19 VDD1.t0 B 0.203322f
C20 VDD1.n1 B 1.79286f
C21 VDD1.t1 B 0.203322f
C22 VDD1.t7 B 0.203322f
C23 VDD1.n2 B 1.79286f
C24 VDD1.n3 B 2.37784f
C25 VDD1.t4 B 0.203322f
C26 VDD1.t6 B 0.203322f
C27 VDD1.n4 B 1.78974f
C28 VDD1.n5 B 2.35694f
C29 VP.n0 B 0.050902f
C30 VP.t6 B 1.0806f
C31 VP.n1 B 0.40795f
C32 VP.n2 B 0.038147f
C33 VP.t7 B 1.0806f
C34 VP.n3 B 0.036093f
C35 VP.n4 B 0.050902f
C36 VP.t1 B 1.14234f
C37 VP.t3 B 1.0806f
C38 VP.n5 B 0.40795f
C39 VP.n6 B 0.193444f
C40 VP.t4 B 1.0806f
C41 VP.t5 B 1.17783f
C42 VP.n7 B 0.458356f
C43 VP.n8 B 0.463913f
C44 VP.n9 B 0.051696f
C45 VP.n10 B 0.051696f
C46 VP.n11 B 0.038147f
C47 VP.n12 B 0.038147f
C48 VP.n13 B 0.044133f
C49 VP.n14 B 0.036093f
C50 VP.n15 B 0.467832f
C51 VP.n16 B 1.60012f
C52 VP.t2 B 1.14234f
C53 VP.n17 B 0.467832f
C54 VP.n18 B 1.63253f
C55 VP.n19 B 0.050902f
C56 VP.n20 B 0.038147f
C57 VP.n21 B 0.044133f
C58 VP.n22 B 0.40795f
C59 VP.n23 B 0.051696f
C60 VP.n24 B 0.051696f
C61 VP.n25 B 0.038147f
C62 VP.n26 B 0.038147f
C63 VP.n27 B 0.044133f
C64 VP.n28 B 0.036093f
C65 VP.t0 B 1.14234f
C66 VP.n29 B 0.467832f
C67 VP.n30 B 0.035726f
C68 VTAIL.t10 B 0.156249f
C69 VTAIL.t15 B 0.156249f
C70 VTAIL.n0 B 1.318f
C71 VTAIL.n1 B 0.272079f
C72 VTAIL.n2 B 0.026296f
C73 VTAIL.n3 B 0.019852f
C74 VTAIL.n4 B 0.010668f
C75 VTAIL.n5 B 0.025214f
C76 VTAIL.n6 B 0.011295f
C77 VTAIL.n7 B 0.019852f
C78 VTAIL.n8 B 0.010981f
C79 VTAIL.n9 B 0.025214f
C80 VTAIL.n10 B 0.011295f
C81 VTAIL.n11 B 0.019852f
C82 VTAIL.n12 B 0.010668f
C83 VTAIL.n13 B 0.025214f
C84 VTAIL.n14 B 0.011295f
C85 VTAIL.n15 B 0.019852f
C86 VTAIL.n16 B 0.010668f
C87 VTAIL.n17 B 0.018911f
C88 VTAIL.n18 B 0.017825f
C89 VTAIL.t8 B 0.042368f
C90 VTAIL.n19 B 0.127585f
C91 VTAIL.n20 B 0.821364f
C92 VTAIL.n21 B 0.010668f
C93 VTAIL.n22 B 0.011295f
C94 VTAIL.n23 B 0.025214f
C95 VTAIL.n24 B 0.025214f
C96 VTAIL.n25 B 0.011295f
C97 VTAIL.n26 B 0.010668f
C98 VTAIL.n27 B 0.019852f
C99 VTAIL.n28 B 0.019852f
C100 VTAIL.n29 B 0.010668f
C101 VTAIL.n30 B 0.011295f
C102 VTAIL.n31 B 0.025214f
C103 VTAIL.n32 B 0.025214f
C104 VTAIL.n33 B 0.011295f
C105 VTAIL.n34 B 0.010668f
C106 VTAIL.n35 B 0.019852f
C107 VTAIL.n36 B 0.019852f
C108 VTAIL.n37 B 0.010668f
C109 VTAIL.n38 B 0.010668f
C110 VTAIL.n39 B 0.011295f
C111 VTAIL.n40 B 0.025214f
C112 VTAIL.n41 B 0.025214f
C113 VTAIL.n42 B 0.025214f
C114 VTAIL.n43 B 0.010981f
C115 VTAIL.n44 B 0.010668f
C116 VTAIL.n45 B 0.019852f
C117 VTAIL.n46 B 0.019852f
C118 VTAIL.n47 B 0.010668f
C119 VTAIL.n48 B 0.011295f
C120 VTAIL.n49 B 0.025214f
C121 VTAIL.n50 B 0.051742f
C122 VTAIL.n51 B 0.011295f
C123 VTAIL.n52 B 0.010668f
C124 VTAIL.n53 B 0.045887f
C125 VTAIL.n54 B 0.02866f
C126 VTAIL.n55 B 0.123108f
C127 VTAIL.n56 B 0.026296f
C128 VTAIL.n57 B 0.019852f
C129 VTAIL.n58 B 0.010668f
C130 VTAIL.n59 B 0.025214f
C131 VTAIL.n60 B 0.011295f
C132 VTAIL.n61 B 0.019852f
C133 VTAIL.n62 B 0.010981f
C134 VTAIL.n63 B 0.025214f
C135 VTAIL.n64 B 0.011295f
C136 VTAIL.n65 B 0.019852f
C137 VTAIL.n66 B 0.010668f
C138 VTAIL.n67 B 0.025214f
C139 VTAIL.n68 B 0.011295f
C140 VTAIL.n69 B 0.019852f
C141 VTAIL.n70 B 0.010668f
C142 VTAIL.n71 B 0.018911f
C143 VTAIL.n72 B 0.017825f
C144 VTAIL.t4 B 0.042368f
C145 VTAIL.n73 B 0.127585f
C146 VTAIL.n74 B 0.821364f
C147 VTAIL.n75 B 0.010668f
C148 VTAIL.n76 B 0.011295f
C149 VTAIL.n77 B 0.025214f
C150 VTAIL.n78 B 0.025214f
C151 VTAIL.n79 B 0.011295f
C152 VTAIL.n80 B 0.010668f
C153 VTAIL.n81 B 0.019852f
C154 VTAIL.n82 B 0.019852f
C155 VTAIL.n83 B 0.010668f
C156 VTAIL.n84 B 0.011295f
C157 VTAIL.n85 B 0.025214f
C158 VTAIL.n86 B 0.025214f
C159 VTAIL.n87 B 0.011295f
C160 VTAIL.n88 B 0.010668f
C161 VTAIL.n89 B 0.019852f
C162 VTAIL.n90 B 0.019852f
C163 VTAIL.n91 B 0.010668f
C164 VTAIL.n92 B 0.010668f
C165 VTAIL.n93 B 0.011295f
C166 VTAIL.n94 B 0.025214f
C167 VTAIL.n95 B 0.025214f
C168 VTAIL.n96 B 0.025214f
C169 VTAIL.n97 B 0.010981f
C170 VTAIL.n98 B 0.010668f
C171 VTAIL.n99 B 0.019852f
C172 VTAIL.n100 B 0.019852f
C173 VTAIL.n101 B 0.010668f
C174 VTAIL.n102 B 0.011295f
C175 VTAIL.n103 B 0.025214f
C176 VTAIL.n104 B 0.051742f
C177 VTAIL.n105 B 0.011295f
C178 VTAIL.n106 B 0.010668f
C179 VTAIL.n107 B 0.045887f
C180 VTAIL.n108 B 0.02866f
C181 VTAIL.n109 B 0.123108f
C182 VTAIL.t1 B 0.156249f
C183 VTAIL.t5 B 0.156249f
C184 VTAIL.n110 B 1.318f
C185 VTAIL.n111 B 0.344456f
C186 VTAIL.n112 B 0.026296f
C187 VTAIL.n113 B 0.019852f
C188 VTAIL.n114 B 0.010668f
C189 VTAIL.n115 B 0.025214f
C190 VTAIL.n116 B 0.011295f
C191 VTAIL.n117 B 0.019852f
C192 VTAIL.n118 B 0.010981f
C193 VTAIL.n119 B 0.025214f
C194 VTAIL.n120 B 0.011295f
C195 VTAIL.n121 B 0.019852f
C196 VTAIL.n122 B 0.010668f
C197 VTAIL.n123 B 0.025214f
C198 VTAIL.n124 B 0.011295f
C199 VTAIL.n125 B 0.019852f
C200 VTAIL.n126 B 0.010668f
C201 VTAIL.n127 B 0.018911f
C202 VTAIL.n128 B 0.017825f
C203 VTAIL.t3 B 0.042368f
C204 VTAIL.n129 B 0.127585f
C205 VTAIL.n130 B 0.821364f
C206 VTAIL.n131 B 0.010668f
C207 VTAIL.n132 B 0.011295f
C208 VTAIL.n133 B 0.025214f
C209 VTAIL.n134 B 0.025214f
C210 VTAIL.n135 B 0.011295f
C211 VTAIL.n136 B 0.010668f
C212 VTAIL.n137 B 0.019852f
C213 VTAIL.n138 B 0.019852f
C214 VTAIL.n139 B 0.010668f
C215 VTAIL.n140 B 0.011295f
C216 VTAIL.n141 B 0.025214f
C217 VTAIL.n142 B 0.025214f
C218 VTAIL.n143 B 0.011295f
C219 VTAIL.n144 B 0.010668f
C220 VTAIL.n145 B 0.019852f
C221 VTAIL.n146 B 0.019852f
C222 VTAIL.n147 B 0.010668f
C223 VTAIL.n148 B 0.010668f
C224 VTAIL.n149 B 0.011295f
C225 VTAIL.n150 B 0.025214f
C226 VTAIL.n151 B 0.025214f
C227 VTAIL.n152 B 0.025214f
C228 VTAIL.n153 B 0.010981f
C229 VTAIL.n154 B 0.010668f
C230 VTAIL.n155 B 0.019852f
C231 VTAIL.n156 B 0.019852f
C232 VTAIL.n157 B 0.010668f
C233 VTAIL.n158 B 0.011295f
C234 VTAIL.n159 B 0.025214f
C235 VTAIL.n160 B 0.051742f
C236 VTAIL.n161 B 0.011295f
C237 VTAIL.n162 B 0.010668f
C238 VTAIL.n163 B 0.045887f
C239 VTAIL.n164 B 0.02866f
C240 VTAIL.n165 B 0.988057f
C241 VTAIL.n166 B 0.026296f
C242 VTAIL.n167 B 0.019852f
C243 VTAIL.n168 B 0.010668f
C244 VTAIL.n169 B 0.025214f
C245 VTAIL.n170 B 0.011295f
C246 VTAIL.n171 B 0.019852f
C247 VTAIL.n172 B 0.010981f
C248 VTAIL.n173 B 0.025214f
C249 VTAIL.n174 B 0.010668f
C250 VTAIL.n175 B 0.011295f
C251 VTAIL.n176 B 0.019852f
C252 VTAIL.n177 B 0.010668f
C253 VTAIL.n178 B 0.025214f
C254 VTAIL.n179 B 0.011295f
C255 VTAIL.n180 B 0.019852f
C256 VTAIL.n181 B 0.010668f
C257 VTAIL.n182 B 0.018911f
C258 VTAIL.n183 B 0.017825f
C259 VTAIL.t14 B 0.042368f
C260 VTAIL.n184 B 0.127585f
C261 VTAIL.n185 B 0.821364f
C262 VTAIL.n186 B 0.010668f
C263 VTAIL.n187 B 0.011295f
C264 VTAIL.n188 B 0.025214f
C265 VTAIL.n189 B 0.025214f
C266 VTAIL.n190 B 0.011295f
C267 VTAIL.n191 B 0.010668f
C268 VTAIL.n192 B 0.019852f
C269 VTAIL.n193 B 0.019852f
C270 VTAIL.n194 B 0.010668f
C271 VTAIL.n195 B 0.011295f
C272 VTAIL.n196 B 0.025214f
C273 VTAIL.n197 B 0.025214f
C274 VTAIL.n198 B 0.011295f
C275 VTAIL.n199 B 0.010668f
C276 VTAIL.n200 B 0.019852f
C277 VTAIL.n201 B 0.019852f
C278 VTAIL.n202 B 0.010668f
C279 VTAIL.n203 B 0.011295f
C280 VTAIL.n204 B 0.025214f
C281 VTAIL.n205 B 0.025214f
C282 VTAIL.n206 B 0.025214f
C283 VTAIL.n207 B 0.010981f
C284 VTAIL.n208 B 0.010668f
C285 VTAIL.n209 B 0.019852f
C286 VTAIL.n210 B 0.019852f
C287 VTAIL.n211 B 0.010668f
C288 VTAIL.n212 B 0.011295f
C289 VTAIL.n213 B 0.025214f
C290 VTAIL.n214 B 0.051742f
C291 VTAIL.n215 B 0.011295f
C292 VTAIL.n216 B 0.010668f
C293 VTAIL.n217 B 0.045887f
C294 VTAIL.n218 B 0.02866f
C295 VTAIL.n219 B 0.988057f
C296 VTAIL.t13 B 0.156249f
C297 VTAIL.t11 B 0.156249f
C298 VTAIL.n220 B 1.31801f
C299 VTAIL.n221 B 0.344448f
C300 VTAIL.n222 B 0.026296f
C301 VTAIL.n223 B 0.019852f
C302 VTAIL.n224 B 0.010668f
C303 VTAIL.n225 B 0.025214f
C304 VTAIL.n226 B 0.011295f
C305 VTAIL.n227 B 0.019852f
C306 VTAIL.n228 B 0.010981f
C307 VTAIL.n229 B 0.025214f
C308 VTAIL.n230 B 0.010668f
C309 VTAIL.n231 B 0.011295f
C310 VTAIL.n232 B 0.019852f
C311 VTAIL.n233 B 0.010668f
C312 VTAIL.n234 B 0.025214f
C313 VTAIL.n235 B 0.011295f
C314 VTAIL.n236 B 0.019852f
C315 VTAIL.n237 B 0.010668f
C316 VTAIL.n238 B 0.018911f
C317 VTAIL.n239 B 0.017825f
C318 VTAIL.t9 B 0.042368f
C319 VTAIL.n240 B 0.127585f
C320 VTAIL.n241 B 0.821364f
C321 VTAIL.n242 B 0.010668f
C322 VTAIL.n243 B 0.011295f
C323 VTAIL.n244 B 0.025214f
C324 VTAIL.n245 B 0.025214f
C325 VTAIL.n246 B 0.011295f
C326 VTAIL.n247 B 0.010668f
C327 VTAIL.n248 B 0.019852f
C328 VTAIL.n249 B 0.019852f
C329 VTAIL.n250 B 0.010668f
C330 VTAIL.n251 B 0.011295f
C331 VTAIL.n252 B 0.025214f
C332 VTAIL.n253 B 0.025214f
C333 VTAIL.n254 B 0.011295f
C334 VTAIL.n255 B 0.010668f
C335 VTAIL.n256 B 0.019852f
C336 VTAIL.n257 B 0.019852f
C337 VTAIL.n258 B 0.010668f
C338 VTAIL.n259 B 0.011295f
C339 VTAIL.n260 B 0.025214f
C340 VTAIL.n261 B 0.025214f
C341 VTAIL.n262 B 0.025214f
C342 VTAIL.n263 B 0.010981f
C343 VTAIL.n264 B 0.010668f
C344 VTAIL.n265 B 0.019852f
C345 VTAIL.n266 B 0.019852f
C346 VTAIL.n267 B 0.010668f
C347 VTAIL.n268 B 0.011295f
C348 VTAIL.n269 B 0.025214f
C349 VTAIL.n270 B 0.051742f
C350 VTAIL.n271 B 0.011295f
C351 VTAIL.n272 B 0.010668f
C352 VTAIL.n273 B 0.045887f
C353 VTAIL.n274 B 0.02866f
C354 VTAIL.n275 B 0.123108f
C355 VTAIL.n276 B 0.026296f
C356 VTAIL.n277 B 0.019852f
C357 VTAIL.n278 B 0.010668f
C358 VTAIL.n279 B 0.025214f
C359 VTAIL.n280 B 0.011295f
C360 VTAIL.n281 B 0.019852f
C361 VTAIL.n282 B 0.010981f
C362 VTAIL.n283 B 0.025214f
C363 VTAIL.n284 B 0.010668f
C364 VTAIL.n285 B 0.011295f
C365 VTAIL.n286 B 0.019852f
C366 VTAIL.n287 B 0.010668f
C367 VTAIL.n288 B 0.025214f
C368 VTAIL.n289 B 0.011295f
C369 VTAIL.n290 B 0.019852f
C370 VTAIL.n291 B 0.010668f
C371 VTAIL.n292 B 0.018911f
C372 VTAIL.n293 B 0.017825f
C373 VTAIL.t2 B 0.042368f
C374 VTAIL.n294 B 0.127585f
C375 VTAIL.n295 B 0.821364f
C376 VTAIL.n296 B 0.010668f
C377 VTAIL.n297 B 0.011295f
C378 VTAIL.n298 B 0.025214f
C379 VTAIL.n299 B 0.025214f
C380 VTAIL.n300 B 0.011295f
C381 VTAIL.n301 B 0.010668f
C382 VTAIL.n302 B 0.019852f
C383 VTAIL.n303 B 0.019852f
C384 VTAIL.n304 B 0.010668f
C385 VTAIL.n305 B 0.011295f
C386 VTAIL.n306 B 0.025214f
C387 VTAIL.n307 B 0.025214f
C388 VTAIL.n308 B 0.011295f
C389 VTAIL.n309 B 0.010668f
C390 VTAIL.n310 B 0.019852f
C391 VTAIL.n311 B 0.019852f
C392 VTAIL.n312 B 0.010668f
C393 VTAIL.n313 B 0.011295f
C394 VTAIL.n314 B 0.025214f
C395 VTAIL.n315 B 0.025214f
C396 VTAIL.n316 B 0.025214f
C397 VTAIL.n317 B 0.010981f
C398 VTAIL.n318 B 0.010668f
C399 VTAIL.n319 B 0.019852f
C400 VTAIL.n320 B 0.019852f
C401 VTAIL.n321 B 0.010668f
C402 VTAIL.n322 B 0.011295f
C403 VTAIL.n323 B 0.025214f
C404 VTAIL.n324 B 0.051742f
C405 VTAIL.n325 B 0.011295f
C406 VTAIL.n326 B 0.010668f
C407 VTAIL.n327 B 0.045887f
C408 VTAIL.n328 B 0.02866f
C409 VTAIL.n329 B 0.123108f
C410 VTAIL.t6 B 0.156249f
C411 VTAIL.t7 B 0.156249f
C412 VTAIL.n330 B 1.31801f
C413 VTAIL.n331 B 0.344448f
C414 VTAIL.n332 B 0.026296f
C415 VTAIL.n333 B 0.019852f
C416 VTAIL.n334 B 0.010668f
C417 VTAIL.n335 B 0.025214f
C418 VTAIL.n336 B 0.011295f
C419 VTAIL.n337 B 0.019852f
C420 VTAIL.n338 B 0.010981f
C421 VTAIL.n339 B 0.025214f
C422 VTAIL.n340 B 0.010668f
C423 VTAIL.n341 B 0.011295f
C424 VTAIL.n342 B 0.019852f
C425 VTAIL.n343 B 0.010668f
C426 VTAIL.n344 B 0.025214f
C427 VTAIL.n345 B 0.011295f
C428 VTAIL.n346 B 0.019852f
C429 VTAIL.n347 B 0.010668f
C430 VTAIL.n348 B 0.018911f
C431 VTAIL.n349 B 0.017825f
C432 VTAIL.t0 B 0.042368f
C433 VTAIL.n350 B 0.127585f
C434 VTAIL.n351 B 0.821364f
C435 VTAIL.n352 B 0.010668f
C436 VTAIL.n353 B 0.011295f
C437 VTAIL.n354 B 0.025214f
C438 VTAIL.n355 B 0.025214f
C439 VTAIL.n356 B 0.011295f
C440 VTAIL.n357 B 0.010668f
C441 VTAIL.n358 B 0.019852f
C442 VTAIL.n359 B 0.019852f
C443 VTAIL.n360 B 0.010668f
C444 VTAIL.n361 B 0.011295f
C445 VTAIL.n362 B 0.025214f
C446 VTAIL.n363 B 0.025214f
C447 VTAIL.n364 B 0.011295f
C448 VTAIL.n365 B 0.010668f
C449 VTAIL.n366 B 0.019852f
C450 VTAIL.n367 B 0.019852f
C451 VTAIL.n368 B 0.010668f
C452 VTAIL.n369 B 0.011295f
C453 VTAIL.n370 B 0.025214f
C454 VTAIL.n371 B 0.025214f
C455 VTAIL.n372 B 0.025214f
C456 VTAIL.n373 B 0.010981f
C457 VTAIL.n374 B 0.010668f
C458 VTAIL.n375 B 0.019852f
C459 VTAIL.n376 B 0.019852f
C460 VTAIL.n377 B 0.010668f
C461 VTAIL.n378 B 0.011295f
C462 VTAIL.n379 B 0.025214f
C463 VTAIL.n380 B 0.051742f
C464 VTAIL.n381 B 0.011295f
C465 VTAIL.n382 B 0.010668f
C466 VTAIL.n383 B 0.045887f
C467 VTAIL.n384 B 0.02866f
C468 VTAIL.n385 B 0.988057f
C469 VTAIL.n386 B 0.026296f
C470 VTAIL.n387 B 0.019852f
C471 VTAIL.n388 B 0.010668f
C472 VTAIL.n389 B 0.025214f
C473 VTAIL.n390 B 0.011295f
C474 VTAIL.n391 B 0.019852f
C475 VTAIL.n392 B 0.010981f
C476 VTAIL.n393 B 0.025214f
C477 VTAIL.n394 B 0.011295f
C478 VTAIL.n395 B 0.019852f
C479 VTAIL.n396 B 0.010668f
C480 VTAIL.n397 B 0.025214f
C481 VTAIL.n398 B 0.011295f
C482 VTAIL.n399 B 0.019852f
C483 VTAIL.n400 B 0.010668f
C484 VTAIL.n401 B 0.018911f
C485 VTAIL.n402 B 0.017825f
C486 VTAIL.t12 B 0.042368f
C487 VTAIL.n403 B 0.127585f
C488 VTAIL.n404 B 0.821364f
C489 VTAIL.n405 B 0.010668f
C490 VTAIL.n406 B 0.011295f
C491 VTAIL.n407 B 0.025214f
C492 VTAIL.n408 B 0.025214f
C493 VTAIL.n409 B 0.011295f
C494 VTAIL.n410 B 0.010668f
C495 VTAIL.n411 B 0.019852f
C496 VTAIL.n412 B 0.019852f
C497 VTAIL.n413 B 0.010668f
C498 VTAIL.n414 B 0.011295f
C499 VTAIL.n415 B 0.025214f
C500 VTAIL.n416 B 0.025214f
C501 VTAIL.n417 B 0.011295f
C502 VTAIL.n418 B 0.010668f
C503 VTAIL.n419 B 0.019852f
C504 VTAIL.n420 B 0.019852f
C505 VTAIL.n421 B 0.010668f
C506 VTAIL.n422 B 0.010668f
C507 VTAIL.n423 B 0.011295f
C508 VTAIL.n424 B 0.025214f
C509 VTAIL.n425 B 0.025214f
C510 VTAIL.n426 B 0.025214f
C511 VTAIL.n427 B 0.010981f
C512 VTAIL.n428 B 0.010668f
C513 VTAIL.n429 B 0.019852f
C514 VTAIL.n430 B 0.019852f
C515 VTAIL.n431 B 0.010668f
C516 VTAIL.n432 B 0.011295f
C517 VTAIL.n433 B 0.025214f
C518 VTAIL.n434 B 0.051742f
C519 VTAIL.n435 B 0.011295f
C520 VTAIL.n436 B 0.010668f
C521 VTAIL.n437 B 0.045887f
C522 VTAIL.n438 B 0.02866f
C523 VTAIL.n439 B 0.984335f
C524 VDD2.t3 B 0.203255f
C525 VDD2.t7 B 0.203255f
C526 VDD2.n0 B 1.79227f
C527 VDD2.t0 B 0.203255f
C528 VDD2.t4 B 0.203255f
C529 VDD2.n1 B 1.79227f
C530 VDD2.n2 B 2.32213f
C531 VDD2.t6 B 0.203255f
C532 VDD2.t5 B 0.203255f
C533 VDD2.n3 B 1.78915f
C534 VDD2.n4 B 2.32539f
C535 VDD2.t1 B 0.203255f
C536 VDD2.t2 B 0.203255f
C537 VDD2.n5 B 1.79224f
C538 VN.n0 B 0.050136f
C539 VN.t0 B 1.06434f
C540 VN.n1 B 0.401811f
C541 VN.n2 B 0.190533f
C542 VN.t5 B 1.06434f
C543 VN.t7 B 1.16011f
C544 VN.n3 B 0.451459f
C545 VN.n4 B 0.456932f
C546 VN.n5 B 0.050918f
C547 VN.n6 B 0.050918f
C548 VN.n7 B 0.037573f
C549 VN.n8 B 0.037573f
C550 VN.n9 B 0.043469f
C551 VN.n10 B 0.03555f
C552 VN.t3 B 1.12514f
C553 VN.n11 B 0.460792f
C554 VN.n12 B 0.035188f
C555 VN.n13 B 0.050136f
C556 VN.t2 B 1.06434f
C557 VN.n14 B 0.401811f
C558 VN.n15 B 0.190533f
C559 VN.t4 B 1.06434f
C560 VN.t6 B 1.16011f
C561 VN.n16 B 0.451459f
C562 VN.n17 B 0.456932f
C563 VN.n18 B 0.050918f
C564 VN.n19 B 0.050918f
C565 VN.n20 B 0.037573f
C566 VN.n21 B 0.037573f
C567 VN.n22 B 0.043469f
C568 VN.n23 B 0.03555f
C569 VN.t1 B 1.12514f
C570 VN.n24 B 0.460792f
C571 VN.n25 B 1.59711f
.ends

