* NGSPICE file created from diff_pair_sample_0197.ext - technology: sky130A

.subckt diff_pair_sample_0197 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=0 ps=0 w=16.68 l=0.95
X1 B.t8 B.t6 B.t7 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=0 ps=0 w=16.68 l=0.95
X2 VDD1.t3 VP.t0 VTAIL.t7 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=2.7522 pd=17.01 as=6.5052 ps=34.14 w=16.68 l=0.95
X3 VDD1.t2 VP.t1 VTAIL.t5 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=2.7522 pd=17.01 as=6.5052 ps=34.14 w=16.68 l=0.95
X4 VDD2.t3 VN.t0 VTAIL.t0 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=2.7522 pd=17.01 as=6.5052 ps=34.14 w=16.68 l=0.95
X5 VDD2.t2 VN.t1 VTAIL.t2 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=2.7522 pd=17.01 as=6.5052 ps=34.14 w=16.68 l=0.95
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=2.7522 ps=17.01 w=16.68 l=0.95
X7 B.t5 B.t3 B.t4 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=0 ps=0 w=16.68 l=0.95
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=2.7522 ps=17.01 w=16.68 l=0.95
X9 B.t2 B.t0 B.t1 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=0 ps=0 w=16.68 l=0.95
X10 VTAIL.t4 VP.t2 VDD1.t1 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=2.7522 ps=17.01 w=16.68 l=0.95
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n1738_n4304# sky130_fd_pr__pfet_01v8 ad=6.5052 pd=34.14 as=2.7522 ps=17.01 w=16.68 l=0.95
R0 B.n275 B.t9 625.721
R1 B.n124 B.t6 625.721
R2 B.n46 B.t0 625.721
R3 B.n40 B.t3 625.721
R4 B.n377 B.n96 585
R5 B.n376 B.n375 585
R6 B.n374 B.n97 585
R7 B.n373 B.n372 585
R8 B.n371 B.n98 585
R9 B.n370 B.n369 585
R10 B.n368 B.n99 585
R11 B.n367 B.n366 585
R12 B.n365 B.n100 585
R13 B.n364 B.n363 585
R14 B.n362 B.n101 585
R15 B.n361 B.n360 585
R16 B.n359 B.n102 585
R17 B.n358 B.n357 585
R18 B.n356 B.n103 585
R19 B.n355 B.n354 585
R20 B.n353 B.n104 585
R21 B.n352 B.n351 585
R22 B.n350 B.n105 585
R23 B.n349 B.n348 585
R24 B.n347 B.n106 585
R25 B.n346 B.n345 585
R26 B.n344 B.n107 585
R27 B.n343 B.n342 585
R28 B.n341 B.n108 585
R29 B.n340 B.n339 585
R30 B.n338 B.n109 585
R31 B.n337 B.n336 585
R32 B.n335 B.n110 585
R33 B.n334 B.n333 585
R34 B.n332 B.n111 585
R35 B.n331 B.n330 585
R36 B.n329 B.n112 585
R37 B.n328 B.n327 585
R38 B.n326 B.n113 585
R39 B.n325 B.n324 585
R40 B.n323 B.n114 585
R41 B.n322 B.n321 585
R42 B.n320 B.n115 585
R43 B.n319 B.n318 585
R44 B.n317 B.n116 585
R45 B.n316 B.n315 585
R46 B.n314 B.n117 585
R47 B.n313 B.n312 585
R48 B.n311 B.n118 585
R49 B.n310 B.n309 585
R50 B.n308 B.n119 585
R51 B.n307 B.n306 585
R52 B.n305 B.n120 585
R53 B.n304 B.n303 585
R54 B.n302 B.n121 585
R55 B.n301 B.n300 585
R56 B.n299 B.n122 585
R57 B.n298 B.n297 585
R58 B.n296 B.n123 585
R59 B.n294 B.n293 585
R60 B.n292 B.n126 585
R61 B.n291 B.n290 585
R62 B.n289 B.n127 585
R63 B.n288 B.n287 585
R64 B.n286 B.n128 585
R65 B.n285 B.n284 585
R66 B.n283 B.n129 585
R67 B.n282 B.n281 585
R68 B.n280 B.n130 585
R69 B.n279 B.n278 585
R70 B.n274 B.n131 585
R71 B.n273 B.n272 585
R72 B.n271 B.n132 585
R73 B.n270 B.n269 585
R74 B.n268 B.n133 585
R75 B.n267 B.n266 585
R76 B.n265 B.n134 585
R77 B.n264 B.n263 585
R78 B.n262 B.n135 585
R79 B.n261 B.n260 585
R80 B.n259 B.n136 585
R81 B.n258 B.n257 585
R82 B.n256 B.n137 585
R83 B.n255 B.n254 585
R84 B.n253 B.n138 585
R85 B.n252 B.n251 585
R86 B.n250 B.n139 585
R87 B.n249 B.n248 585
R88 B.n247 B.n140 585
R89 B.n246 B.n245 585
R90 B.n244 B.n141 585
R91 B.n243 B.n242 585
R92 B.n241 B.n142 585
R93 B.n240 B.n239 585
R94 B.n238 B.n143 585
R95 B.n237 B.n236 585
R96 B.n235 B.n144 585
R97 B.n234 B.n233 585
R98 B.n232 B.n145 585
R99 B.n231 B.n230 585
R100 B.n229 B.n146 585
R101 B.n228 B.n227 585
R102 B.n226 B.n147 585
R103 B.n225 B.n224 585
R104 B.n223 B.n148 585
R105 B.n222 B.n221 585
R106 B.n220 B.n149 585
R107 B.n219 B.n218 585
R108 B.n217 B.n150 585
R109 B.n216 B.n215 585
R110 B.n214 B.n151 585
R111 B.n213 B.n212 585
R112 B.n211 B.n152 585
R113 B.n210 B.n209 585
R114 B.n208 B.n153 585
R115 B.n207 B.n206 585
R116 B.n205 B.n154 585
R117 B.n204 B.n203 585
R118 B.n202 B.n155 585
R119 B.n201 B.n200 585
R120 B.n199 B.n156 585
R121 B.n198 B.n197 585
R122 B.n196 B.n157 585
R123 B.n195 B.n194 585
R124 B.n379 B.n378 585
R125 B.n380 B.n95 585
R126 B.n382 B.n381 585
R127 B.n383 B.n94 585
R128 B.n385 B.n384 585
R129 B.n386 B.n93 585
R130 B.n388 B.n387 585
R131 B.n389 B.n92 585
R132 B.n391 B.n390 585
R133 B.n392 B.n91 585
R134 B.n394 B.n393 585
R135 B.n395 B.n90 585
R136 B.n397 B.n396 585
R137 B.n398 B.n89 585
R138 B.n400 B.n399 585
R139 B.n401 B.n88 585
R140 B.n403 B.n402 585
R141 B.n404 B.n87 585
R142 B.n406 B.n405 585
R143 B.n407 B.n86 585
R144 B.n409 B.n408 585
R145 B.n410 B.n85 585
R146 B.n412 B.n411 585
R147 B.n413 B.n84 585
R148 B.n415 B.n414 585
R149 B.n416 B.n83 585
R150 B.n418 B.n417 585
R151 B.n419 B.n82 585
R152 B.n421 B.n420 585
R153 B.n422 B.n81 585
R154 B.n424 B.n423 585
R155 B.n425 B.n80 585
R156 B.n427 B.n426 585
R157 B.n428 B.n79 585
R158 B.n430 B.n429 585
R159 B.n431 B.n78 585
R160 B.n433 B.n432 585
R161 B.n434 B.n77 585
R162 B.n436 B.n435 585
R163 B.n437 B.n76 585
R164 B.n619 B.n618 585
R165 B.n617 B.n12 585
R166 B.n616 B.n615 585
R167 B.n614 B.n13 585
R168 B.n613 B.n612 585
R169 B.n611 B.n14 585
R170 B.n610 B.n609 585
R171 B.n608 B.n15 585
R172 B.n607 B.n606 585
R173 B.n605 B.n16 585
R174 B.n604 B.n603 585
R175 B.n602 B.n17 585
R176 B.n601 B.n600 585
R177 B.n599 B.n18 585
R178 B.n598 B.n597 585
R179 B.n596 B.n19 585
R180 B.n595 B.n594 585
R181 B.n593 B.n20 585
R182 B.n592 B.n591 585
R183 B.n590 B.n21 585
R184 B.n589 B.n588 585
R185 B.n587 B.n22 585
R186 B.n586 B.n585 585
R187 B.n584 B.n23 585
R188 B.n583 B.n582 585
R189 B.n581 B.n24 585
R190 B.n580 B.n579 585
R191 B.n578 B.n25 585
R192 B.n577 B.n576 585
R193 B.n575 B.n26 585
R194 B.n574 B.n573 585
R195 B.n572 B.n27 585
R196 B.n571 B.n570 585
R197 B.n569 B.n28 585
R198 B.n568 B.n567 585
R199 B.n566 B.n29 585
R200 B.n565 B.n564 585
R201 B.n563 B.n30 585
R202 B.n562 B.n561 585
R203 B.n560 B.n31 585
R204 B.n559 B.n558 585
R205 B.n557 B.n32 585
R206 B.n556 B.n555 585
R207 B.n554 B.n33 585
R208 B.n553 B.n552 585
R209 B.n551 B.n34 585
R210 B.n550 B.n549 585
R211 B.n548 B.n35 585
R212 B.n547 B.n546 585
R213 B.n545 B.n36 585
R214 B.n544 B.n543 585
R215 B.n542 B.n37 585
R216 B.n541 B.n540 585
R217 B.n539 B.n38 585
R218 B.n538 B.n537 585
R219 B.n535 B.n39 585
R220 B.n534 B.n533 585
R221 B.n532 B.n42 585
R222 B.n531 B.n530 585
R223 B.n529 B.n43 585
R224 B.n528 B.n527 585
R225 B.n526 B.n44 585
R226 B.n525 B.n524 585
R227 B.n523 B.n45 585
R228 B.n522 B.n521 585
R229 B.n520 B.n519 585
R230 B.n518 B.n49 585
R231 B.n517 B.n516 585
R232 B.n515 B.n50 585
R233 B.n514 B.n513 585
R234 B.n512 B.n51 585
R235 B.n511 B.n510 585
R236 B.n509 B.n52 585
R237 B.n508 B.n507 585
R238 B.n506 B.n53 585
R239 B.n505 B.n504 585
R240 B.n503 B.n54 585
R241 B.n502 B.n501 585
R242 B.n500 B.n55 585
R243 B.n499 B.n498 585
R244 B.n497 B.n56 585
R245 B.n496 B.n495 585
R246 B.n494 B.n57 585
R247 B.n493 B.n492 585
R248 B.n491 B.n58 585
R249 B.n490 B.n489 585
R250 B.n488 B.n59 585
R251 B.n487 B.n486 585
R252 B.n485 B.n60 585
R253 B.n484 B.n483 585
R254 B.n482 B.n61 585
R255 B.n481 B.n480 585
R256 B.n479 B.n62 585
R257 B.n478 B.n477 585
R258 B.n476 B.n63 585
R259 B.n475 B.n474 585
R260 B.n473 B.n64 585
R261 B.n472 B.n471 585
R262 B.n470 B.n65 585
R263 B.n469 B.n468 585
R264 B.n467 B.n66 585
R265 B.n466 B.n465 585
R266 B.n464 B.n67 585
R267 B.n463 B.n462 585
R268 B.n461 B.n68 585
R269 B.n460 B.n459 585
R270 B.n458 B.n69 585
R271 B.n457 B.n456 585
R272 B.n455 B.n70 585
R273 B.n454 B.n453 585
R274 B.n452 B.n71 585
R275 B.n451 B.n450 585
R276 B.n449 B.n72 585
R277 B.n448 B.n447 585
R278 B.n446 B.n73 585
R279 B.n445 B.n444 585
R280 B.n443 B.n74 585
R281 B.n442 B.n441 585
R282 B.n440 B.n75 585
R283 B.n439 B.n438 585
R284 B.n620 B.n11 585
R285 B.n622 B.n621 585
R286 B.n623 B.n10 585
R287 B.n625 B.n624 585
R288 B.n626 B.n9 585
R289 B.n628 B.n627 585
R290 B.n629 B.n8 585
R291 B.n631 B.n630 585
R292 B.n632 B.n7 585
R293 B.n634 B.n633 585
R294 B.n635 B.n6 585
R295 B.n637 B.n636 585
R296 B.n638 B.n5 585
R297 B.n640 B.n639 585
R298 B.n641 B.n4 585
R299 B.n643 B.n642 585
R300 B.n644 B.n3 585
R301 B.n646 B.n645 585
R302 B.n647 B.n0 585
R303 B.n2 B.n1 585
R304 B.n168 B.n167 585
R305 B.n169 B.n166 585
R306 B.n171 B.n170 585
R307 B.n172 B.n165 585
R308 B.n174 B.n173 585
R309 B.n175 B.n164 585
R310 B.n177 B.n176 585
R311 B.n178 B.n163 585
R312 B.n180 B.n179 585
R313 B.n181 B.n162 585
R314 B.n183 B.n182 585
R315 B.n184 B.n161 585
R316 B.n186 B.n185 585
R317 B.n187 B.n160 585
R318 B.n189 B.n188 585
R319 B.n190 B.n159 585
R320 B.n192 B.n191 585
R321 B.n193 B.n158 585
R322 B.n194 B.n193 511.721
R323 B.n378 B.n377 511.721
R324 B.n438 B.n437 511.721
R325 B.n618 B.n11 511.721
R326 B.n124 B.t7 484.538
R327 B.n46 B.t2 484.538
R328 B.n275 B.t10 484.538
R329 B.n40 B.t5 484.538
R330 B.n125 B.t8 459.714
R331 B.n47 B.t1 459.714
R332 B.n276 B.t11 459.714
R333 B.n41 B.t4 459.714
R334 B.n649 B.n648 256.663
R335 B.n648 B.n647 235.042
R336 B.n648 B.n2 235.042
R337 B.n194 B.n157 163.367
R338 B.n198 B.n157 163.367
R339 B.n199 B.n198 163.367
R340 B.n200 B.n199 163.367
R341 B.n200 B.n155 163.367
R342 B.n204 B.n155 163.367
R343 B.n205 B.n204 163.367
R344 B.n206 B.n205 163.367
R345 B.n206 B.n153 163.367
R346 B.n210 B.n153 163.367
R347 B.n211 B.n210 163.367
R348 B.n212 B.n211 163.367
R349 B.n212 B.n151 163.367
R350 B.n216 B.n151 163.367
R351 B.n217 B.n216 163.367
R352 B.n218 B.n217 163.367
R353 B.n218 B.n149 163.367
R354 B.n222 B.n149 163.367
R355 B.n223 B.n222 163.367
R356 B.n224 B.n223 163.367
R357 B.n224 B.n147 163.367
R358 B.n228 B.n147 163.367
R359 B.n229 B.n228 163.367
R360 B.n230 B.n229 163.367
R361 B.n230 B.n145 163.367
R362 B.n234 B.n145 163.367
R363 B.n235 B.n234 163.367
R364 B.n236 B.n235 163.367
R365 B.n236 B.n143 163.367
R366 B.n240 B.n143 163.367
R367 B.n241 B.n240 163.367
R368 B.n242 B.n241 163.367
R369 B.n242 B.n141 163.367
R370 B.n246 B.n141 163.367
R371 B.n247 B.n246 163.367
R372 B.n248 B.n247 163.367
R373 B.n248 B.n139 163.367
R374 B.n252 B.n139 163.367
R375 B.n253 B.n252 163.367
R376 B.n254 B.n253 163.367
R377 B.n254 B.n137 163.367
R378 B.n258 B.n137 163.367
R379 B.n259 B.n258 163.367
R380 B.n260 B.n259 163.367
R381 B.n260 B.n135 163.367
R382 B.n264 B.n135 163.367
R383 B.n265 B.n264 163.367
R384 B.n266 B.n265 163.367
R385 B.n266 B.n133 163.367
R386 B.n270 B.n133 163.367
R387 B.n271 B.n270 163.367
R388 B.n272 B.n271 163.367
R389 B.n272 B.n131 163.367
R390 B.n279 B.n131 163.367
R391 B.n280 B.n279 163.367
R392 B.n281 B.n280 163.367
R393 B.n281 B.n129 163.367
R394 B.n285 B.n129 163.367
R395 B.n286 B.n285 163.367
R396 B.n287 B.n286 163.367
R397 B.n287 B.n127 163.367
R398 B.n291 B.n127 163.367
R399 B.n292 B.n291 163.367
R400 B.n293 B.n292 163.367
R401 B.n293 B.n123 163.367
R402 B.n298 B.n123 163.367
R403 B.n299 B.n298 163.367
R404 B.n300 B.n299 163.367
R405 B.n300 B.n121 163.367
R406 B.n304 B.n121 163.367
R407 B.n305 B.n304 163.367
R408 B.n306 B.n305 163.367
R409 B.n306 B.n119 163.367
R410 B.n310 B.n119 163.367
R411 B.n311 B.n310 163.367
R412 B.n312 B.n311 163.367
R413 B.n312 B.n117 163.367
R414 B.n316 B.n117 163.367
R415 B.n317 B.n316 163.367
R416 B.n318 B.n317 163.367
R417 B.n318 B.n115 163.367
R418 B.n322 B.n115 163.367
R419 B.n323 B.n322 163.367
R420 B.n324 B.n323 163.367
R421 B.n324 B.n113 163.367
R422 B.n328 B.n113 163.367
R423 B.n329 B.n328 163.367
R424 B.n330 B.n329 163.367
R425 B.n330 B.n111 163.367
R426 B.n334 B.n111 163.367
R427 B.n335 B.n334 163.367
R428 B.n336 B.n335 163.367
R429 B.n336 B.n109 163.367
R430 B.n340 B.n109 163.367
R431 B.n341 B.n340 163.367
R432 B.n342 B.n341 163.367
R433 B.n342 B.n107 163.367
R434 B.n346 B.n107 163.367
R435 B.n347 B.n346 163.367
R436 B.n348 B.n347 163.367
R437 B.n348 B.n105 163.367
R438 B.n352 B.n105 163.367
R439 B.n353 B.n352 163.367
R440 B.n354 B.n353 163.367
R441 B.n354 B.n103 163.367
R442 B.n358 B.n103 163.367
R443 B.n359 B.n358 163.367
R444 B.n360 B.n359 163.367
R445 B.n360 B.n101 163.367
R446 B.n364 B.n101 163.367
R447 B.n365 B.n364 163.367
R448 B.n366 B.n365 163.367
R449 B.n366 B.n99 163.367
R450 B.n370 B.n99 163.367
R451 B.n371 B.n370 163.367
R452 B.n372 B.n371 163.367
R453 B.n372 B.n97 163.367
R454 B.n376 B.n97 163.367
R455 B.n377 B.n376 163.367
R456 B.n437 B.n436 163.367
R457 B.n436 B.n77 163.367
R458 B.n432 B.n77 163.367
R459 B.n432 B.n431 163.367
R460 B.n431 B.n430 163.367
R461 B.n430 B.n79 163.367
R462 B.n426 B.n79 163.367
R463 B.n426 B.n425 163.367
R464 B.n425 B.n424 163.367
R465 B.n424 B.n81 163.367
R466 B.n420 B.n81 163.367
R467 B.n420 B.n419 163.367
R468 B.n419 B.n418 163.367
R469 B.n418 B.n83 163.367
R470 B.n414 B.n83 163.367
R471 B.n414 B.n413 163.367
R472 B.n413 B.n412 163.367
R473 B.n412 B.n85 163.367
R474 B.n408 B.n85 163.367
R475 B.n408 B.n407 163.367
R476 B.n407 B.n406 163.367
R477 B.n406 B.n87 163.367
R478 B.n402 B.n87 163.367
R479 B.n402 B.n401 163.367
R480 B.n401 B.n400 163.367
R481 B.n400 B.n89 163.367
R482 B.n396 B.n89 163.367
R483 B.n396 B.n395 163.367
R484 B.n395 B.n394 163.367
R485 B.n394 B.n91 163.367
R486 B.n390 B.n91 163.367
R487 B.n390 B.n389 163.367
R488 B.n389 B.n388 163.367
R489 B.n388 B.n93 163.367
R490 B.n384 B.n93 163.367
R491 B.n384 B.n383 163.367
R492 B.n383 B.n382 163.367
R493 B.n382 B.n95 163.367
R494 B.n378 B.n95 163.367
R495 B.n618 B.n617 163.367
R496 B.n617 B.n616 163.367
R497 B.n616 B.n13 163.367
R498 B.n612 B.n13 163.367
R499 B.n612 B.n611 163.367
R500 B.n611 B.n610 163.367
R501 B.n610 B.n15 163.367
R502 B.n606 B.n15 163.367
R503 B.n606 B.n605 163.367
R504 B.n605 B.n604 163.367
R505 B.n604 B.n17 163.367
R506 B.n600 B.n17 163.367
R507 B.n600 B.n599 163.367
R508 B.n599 B.n598 163.367
R509 B.n598 B.n19 163.367
R510 B.n594 B.n19 163.367
R511 B.n594 B.n593 163.367
R512 B.n593 B.n592 163.367
R513 B.n592 B.n21 163.367
R514 B.n588 B.n21 163.367
R515 B.n588 B.n587 163.367
R516 B.n587 B.n586 163.367
R517 B.n586 B.n23 163.367
R518 B.n582 B.n23 163.367
R519 B.n582 B.n581 163.367
R520 B.n581 B.n580 163.367
R521 B.n580 B.n25 163.367
R522 B.n576 B.n25 163.367
R523 B.n576 B.n575 163.367
R524 B.n575 B.n574 163.367
R525 B.n574 B.n27 163.367
R526 B.n570 B.n27 163.367
R527 B.n570 B.n569 163.367
R528 B.n569 B.n568 163.367
R529 B.n568 B.n29 163.367
R530 B.n564 B.n29 163.367
R531 B.n564 B.n563 163.367
R532 B.n563 B.n562 163.367
R533 B.n562 B.n31 163.367
R534 B.n558 B.n31 163.367
R535 B.n558 B.n557 163.367
R536 B.n557 B.n556 163.367
R537 B.n556 B.n33 163.367
R538 B.n552 B.n33 163.367
R539 B.n552 B.n551 163.367
R540 B.n551 B.n550 163.367
R541 B.n550 B.n35 163.367
R542 B.n546 B.n35 163.367
R543 B.n546 B.n545 163.367
R544 B.n545 B.n544 163.367
R545 B.n544 B.n37 163.367
R546 B.n540 B.n37 163.367
R547 B.n540 B.n539 163.367
R548 B.n539 B.n538 163.367
R549 B.n538 B.n39 163.367
R550 B.n533 B.n39 163.367
R551 B.n533 B.n532 163.367
R552 B.n532 B.n531 163.367
R553 B.n531 B.n43 163.367
R554 B.n527 B.n43 163.367
R555 B.n527 B.n526 163.367
R556 B.n526 B.n525 163.367
R557 B.n525 B.n45 163.367
R558 B.n521 B.n45 163.367
R559 B.n521 B.n520 163.367
R560 B.n520 B.n49 163.367
R561 B.n516 B.n49 163.367
R562 B.n516 B.n515 163.367
R563 B.n515 B.n514 163.367
R564 B.n514 B.n51 163.367
R565 B.n510 B.n51 163.367
R566 B.n510 B.n509 163.367
R567 B.n509 B.n508 163.367
R568 B.n508 B.n53 163.367
R569 B.n504 B.n53 163.367
R570 B.n504 B.n503 163.367
R571 B.n503 B.n502 163.367
R572 B.n502 B.n55 163.367
R573 B.n498 B.n55 163.367
R574 B.n498 B.n497 163.367
R575 B.n497 B.n496 163.367
R576 B.n496 B.n57 163.367
R577 B.n492 B.n57 163.367
R578 B.n492 B.n491 163.367
R579 B.n491 B.n490 163.367
R580 B.n490 B.n59 163.367
R581 B.n486 B.n59 163.367
R582 B.n486 B.n485 163.367
R583 B.n485 B.n484 163.367
R584 B.n484 B.n61 163.367
R585 B.n480 B.n61 163.367
R586 B.n480 B.n479 163.367
R587 B.n479 B.n478 163.367
R588 B.n478 B.n63 163.367
R589 B.n474 B.n63 163.367
R590 B.n474 B.n473 163.367
R591 B.n473 B.n472 163.367
R592 B.n472 B.n65 163.367
R593 B.n468 B.n65 163.367
R594 B.n468 B.n467 163.367
R595 B.n467 B.n466 163.367
R596 B.n466 B.n67 163.367
R597 B.n462 B.n67 163.367
R598 B.n462 B.n461 163.367
R599 B.n461 B.n460 163.367
R600 B.n460 B.n69 163.367
R601 B.n456 B.n69 163.367
R602 B.n456 B.n455 163.367
R603 B.n455 B.n454 163.367
R604 B.n454 B.n71 163.367
R605 B.n450 B.n71 163.367
R606 B.n450 B.n449 163.367
R607 B.n449 B.n448 163.367
R608 B.n448 B.n73 163.367
R609 B.n444 B.n73 163.367
R610 B.n444 B.n443 163.367
R611 B.n443 B.n442 163.367
R612 B.n442 B.n75 163.367
R613 B.n438 B.n75 163.367
R614 B.n622 B.n11 163.367
R615 B.n623 B.n622 163.367
R616 B.n624 B.n623 163.367
R617 B.n624 B.n9 163.367
R618 B.n628 B.n9 163.367
R619 B.n629 B.n628 163.367
R620 B.n630 B.n629 163.367
R621 B.n630 B.n7 163.367
R622 B.n634 B.n7 163.367
R623 B.n635 B.n634 163.367
R624 B.n636 B.n635 163.367
R625 B.n636 B.n5 163.367
R626 B.n640 B.n5 163.367
R627 B.n641 B.n640 163.367
R628 B.n642 B.n641 163.367
R629 B.n642 B.n3 163.367
R630 B.n646 B.n3 163.367
R631 B.n647 B.n646 163.367
R632 B.n168 B.n2 163.367
R633 B.n169 B.n168 163.367
R634 B.n170 B.n169 163.367
R635 B.n170 B.n165 163.367
R636 B.n174 B.n165 163.367
R637 B.n175 B.n174 163.367
R638 B.n176 B.n175 163.367
R639 B.n176 B.n163 163.367
R640 B.n180 B.n163 163.367
R641 B.n181 B.n180 163.367
R642 B.n182 B.n181 163.367
R643 B.n182 B.n161 163.367
R644 B.n186 B.n161 163.367
R645 B.n187 B.n186 163.367
R646 B.n188 B.n187 163.367
R647 B.n188 B.n159 163.367
R648 B.n192 B.n159 163.367
R649 B.n193 B.n192 163.367
R650 B.n277 B.n276 59.5399
R651 B.n295 B.n125 59.5399
R652 B.n48 B.n47 59.5399
R653 B.n536 B.n41 59.5399
R654 B.n620 B.n619 33.2493
R655 B.n439 B.n76 33.2493
R656 B.n379 B.n96 33.2493
R657 B.n195 B.n158 33.2493
R658 B.n276 B.n275 24.8247
R659 B.n125 B.n124 24.8247
R660 B.n47 B.n46 24.8247
R661 B.n41 B.n40 24.8247
R662 B B.n649 18.0485
R663 B.n621 B.n620 10.6151
R664 B.n621 B.n10 10.6151
R665 B.n625 B.n10 10.6151
R666 B.n626 B.n625 10.6151
R667 B.n627 B.n626 10.6151
R668 B.n627 B.n8 10.6151
R669 B.n631 B.n8 10.6151
R670 B.n632 B.n631 10.6151
R671 B.n633 B.n632 10.6151
R672 B.n633 B.n6 10.6151
R673 B.n637 B.n6 10.6151
R674 B.n638 B.n637 10.6151
R675 B.n639 B.n638 10.6151
R676 B.n639 B.n4 10.6151
R677 B.n643 B.n4 10.6151
R678 B.n644 B.n643 10.6151
R679 B.n645 B.n644 10.6151
R680 B.n645 B.n0 10.6151
R681 B.n619 B.n12 10.6151
R682 B.n615 B.n12 10.6151
R683 B.n615 B.n614 10.6151
R684 B.n614 B.n613 10.6151
R685 B.n613 B.n14 10.6151
R686 B.n609 B.n14 10.6151
R687 B.n609 B.n608 10.6151
R688 B.n608 B.n607 10.6151
R689 B.n607 B.n16 10.6151
R690 B.n603 B.n16 10.6151
R691 B.n603 B.n602 10.6151
R692 B.n602 B.n601 10.6151
R693 B.n601 B.n18 10.6151
R694 B.n597 B.n18 10.6151
R695 B.n597 B.n596 10.6151
R696 B.n596 B.n595 10.6151
R697 B.n595 B.n20 10.6151
R698 B.n591 B.n20 10.6151
R699 B.n591 B.n590 10.6151
R700 B.n590 B.n589 10.6151
R701 B.n589 B.n22 10.6151
R702 B.n585 B.n22 10.6151
R703 B.n585 B.n584 10.6151
R704 B.n584 B.n583 10.6151
R705 B.n583 B.n24 10.6151
R706 B.n579 B.n24 10.6151
R707 B.n579 B.n578 10.6151
R708 B.n578 B.n577 10.6151
R709 B.n577 B.n26 10.6151
R710 B.n573 B.n26 10.6151
R711 B.n573 B.n572 10.6151
R712 B.n572 B.n571 10.6151
R713 B.n571 B.n28 10.6151
R714 B.n567 B.n28 10.6151
R715 B.n567 B.n566 10.6151
R716 B.n566 B.n565 10.6151
R717 B.n565 B.n30 10.6151
R718 B.n561 B.n30 10.6151
R719 B.n561 B.n560 10.6151
R720 B.n560 B.n559 10.6151
R721 B.n559 B.n32 10.6151
R722 B.n555 B.n32 10.6151
R723 B.n555 B.n554 10.6151
R724 B.n554 B.n553 10.6151
R725 B.n553 B.n34 10.6151
R726 B.n549 B.n34 10.6151
R727 B.n549 B.n548 10.6151
R728 B.n548 B.n547 10.6151
R729 B.n547 B.n36 10.6151
R730 B.n543 B.n36 10.6151
R731 B.n543 B.n542 10.6151
R732 B.n542 B.n541 10.6151
R733 B.n541 B.n38 10.6151
R734 B.n537 B.n38 10.6151
R735 B.n535 B.n534 10.6151
R736 B.n534 B.n42 10.6151
R737 B.n530 B.n42 10.6151
R738 B.n530 B.n529 10.6151
R739 B.n529 B.n528 10.6151
R740 B.n528 B.n44 10.6151
R741 B.n524 B.n44 10.6151
R742 B.n524 B.n523 10.6151
R743 B.n523 B.n522 10.6151
R744 B.n519 B.n518 10.6151
R745 B.n518 B.n517 10.6151
R746 B.n517 B.n50 10.6151
R747 B.n513 B.n50 10.6151
R748 B.n513 B.n512 10.6151
R749 B.n512 B.n511 10.6151
R750 B.n511 B.n52 10.6151
R751 B.n507 B.n52 10.6151
R752 B.n507 B.n506 10.6151
R753 B.n506 B.n505 10.6151
R754 B.n505 B.n54 10.6151
R755 B.n501 B.n54 10.6151
R756 B.n501 B.n500 10.6151
R757 B.n500 B.n499 10.6151
R758 B.n499 B.n56 10.6151
R759 B.n495 B.n56 10.6151
R760 B.n495 B.n494 10.6151
R761 B.n494 B.n493 10.6151
R762 B.n493 B.n58 10.6151
R763 B.n489 B.n58 10.6151
R764 B.n489 B.n488 10.6151
R765 B.n488 B.n487 10.6151
R766 B.n487 B.n60 10.6151
R767 B.n483 B.n60 10.6151
R768 B.n483 B.n482 10.6151
R769 B.n482 B.n481 10.6151
R770 B.n481 B.n62 10.6151
R771 B.n477 B.n62 10.6151
R772 B.n477 B.n476 10.6151
R773 B.n476 B.n475 10.6151
R774 B.n475 B.n64 10.6151
R775 B.n471 B.n64 10.6151
R776 B.n471 B.n470 10.6151
R777 B.n470 B.n469 10.6151
R778 B.n469 B.n66 10.6151
R779 B.n465 B.n66 10.6151
R780 B.n465 B.n464 10.6151
R781 B.n464 B.n463 10.6151
R782 B.n463 B.n68 10.6151
R783 B.n459 B.n68 10.6151
R784 B.n459 B.n458 10.6151
R785 B.n458 B.n457 10.6151
R786 B.n457 B.n70 10.6151
R787 B.n453 B.n70 10.6151
R788 B.n453 B.n452 10.6151
R789 B.n452 B.n451 10.6151
R790 B.n451 B.n72 10.6151
R791 B.n447 B.n72 10.6151
R792 B.n447 B.n446 10.6151
R793 B.n446 B.n445 10.6151
R794 B.n445 B.n74 10.6151
R795 B.n441 B.n74 10.6151
R796 B.n441 B.n440 10.6151
R797 B.n440 B.n439 10.6151
R798 B.n435 B.n76 10.6151
R799 B.n435 B.n434 10.6151
R800 B.n434 B.n433 10.6151
R801 B.n433 B.n78 10.6151
R802 B.n429 B.n78 10.6151
R803 B.n429 B.n428 10.6151
R804 B.n428 B.n427 10.6151
R805 B.n427 B.n80 10.6151
R806 B.n423 B.n80 10.6151
R807 B.n423 B.n422 10.6151
R808 B.n422 B.n421 10.6151
R809 B.n421 B.n82 10.6151
R810 B.n417 B.n82 10.6151
R811 B.n417 B.n416 10.6151
R812 B.n416 B.n415 10.6151
R813 B.n415 B.n84 10.6151
R814 B.n411 B.n84 10.6151
R815 B.n411 B.n410 10.6151
R816 B.n410 B.n409 10.6151
R817 B.n409 B.n86 10.6151
R818 B.n405 B.n86 10.6151
R819 B.n405 B.n404 10.6151
R820 B.n404 B.n403 10.6151
R821 B.n403 B.n88 10.6151
R822 B.n399 B.n88 10.6151
R823 B.n399 B.n398 10.6151
R824 B.n398 B.n397 10.6151
R825 B.n397 B.n90 10.6151
R826 B.n393 B.n90 10.6151
R827 B.n393 B.n392 10.6151
R828 B.n392 B.n391 10.6151
R829 B.n391 B.n92 10.6151
R830 B.n387 B.n92 10.6151
R831 B.n387 B.n386 10.6151
R832 B.n386 B.n385 10.6151
R833 B.n385 B.n94 10.6151
R834 B.n381 B.n94 10.6151
R835 B.n381 B.n380 10.6151
R836 B.n380 B.n379 10.6151
R837 B.n167 B.n1 10.6151
R838 B.n167 B.n166 10.6151
R839 B.n171 B.n166 10.6151
R840 B.n172 B.n171 10.6151
R841 B.n173 B.n172 10.6151
R842 B.n173 B.n164 10.6151
R843 B.n177 B.n164 10.6151
R844 B.n178 B.n177 10.6151
R845 B.n179 B.n178 10.6151
R846 B.n179 B.n162 10.6151
R847 B.n183 B.n162 10.6151
R848 B.n184 B.n183 10.6151
R849 B.n185 B.n184 10.6151
R850 B.n185 B.n160 10.6151
R851 B.n189 B.n160 10.6151
R852 B.n190 B.n189 10.6151
R853 B.n191 B.n190 10.6151
R854 B.n191 B.n158 10.6151
R855 B.n196 B.n195 10.6151
R856 B.n197 B.n196 10.6151
R857 B.n197 B.n156 10.6151
R858 B.n201 B.n156 10.6151
R859 B.n202 B.n201 10.6151
R860 B.n203 B.n202 10.6151
R861 B.n203 B.n154 10.6151
R862 B.n207 B.n154 10.6151
R863 B.n208 B.n207 10.6151
R864 B.n209 B.n208 10.6151
R865 B.n209 B.n152 10.6151
R866 B.n213 B.n152 10.6151
R867 B.n214 B.n213 10.6151
R868 B.n215 B.n214 10.6151
R869 B.n215 B.n150 10.6151
R870 B.n219 B.n150 10.6151
R871 B.n220 B.n219 10.6151
R872 B.n221 B.n220 10.6151
R873 B.n221 B.n148 10.6151
R874 B.n225 B.n148 10.6151
R875 B.n226 B.n225 10.6151
R876 B.n227 B.n226 10.6151
R877 B.n227 B.n146 10.6151
R878 B.n231 B.n146 10.6151
R879 B.n232 B.n231 10.6151
R880 B.n233 B.n232 10.6151
R881 B.n233 B.n144 10.6151
R882 B.n237 B.n144 10.6151
R883 B.n238 B.n237 10.6151
R884 B.n239 B.n238 10.6151
R885 B.n239 B.n142 10.6151
R886 B.n243 B.n142 10.6151
R887 B.n244 B.n243 10.6151
R888 B.n245 B.n244 10.6151
R889 B.n245 B.n140 10.6151
R890 B.n249 B.n140 10.6151
R891 B.n250 B.n249 10.6151
R892 B.n251 B.n250 10.6151
R893 B.n251 B.n138 10.6151
R894 B.n255 B.n138 10.6151
R895 B.n256 B.n255 10.6151
R896 B.n257 B.n256 10.6151
R897 B.n257 B.n136 10.6151
R898 B.n261 B.n136 10.6151
R899 B.n262 B.n261 10.6151
R900 B.n263 B.n262 10.6151
R901 B.n263 B.n134 10.6151
R902 B.n267 B.n134 10.6151
R903 B.n268 B.n267 10.6151
R904 B.n269 B.n268 10.6151
R905 B.n269 B.n132 10.6151
R906 B.n273 B.n132 10.6151
R907 B.n274 B.n273 10.6151
R908 B.n278 B.n274 10.6151
R909 B.n282 B.n130 10.6151
R910 B.n283 B.n282 10.6151
R911 B.n284 B.n283 10.6151
R912 B.n284 B.n128 10.6151
R913 B.n288 B.n128 10.6151
R914 B.n289 B.n288 10.6151
R915 B.n290 B.n289 10.6151
R916 B.n290 B.n126 10.6151
R917 B.n294 B.n126 10.6151
R918 B.n297 B.n296 10.6151
R919 B.n297 B.n122 10.6151
R920 B.n301 B.n122 10.6151
R921 B.n302 B.n301 10.6151
R922 B.n303 B.n302 10.6151
R923 B.n303 B.n120 10.6151
R924 B.n307 B.n120 10.6151
R925 B.n308 B.n307 10.6151
R926 B.n309 B.n308 10.6151
R927 B.n309 B.n118 10.6151
R928 B.n313 B.n118 10.6151
R929 B.n314 B.n313 10.6151
R930 B.n315 B.n314 10.6151
R931 B.n315 B.n116 10.6151
R932 B.n319 B.n116 10.6151
R933 B.n320 B.n319 10.6151
R934 B.n321 B.n320 10.6151
R935 B.n321 B.n114 10.6151
R936 B.n325 B.n114 10.6151
R937 B.n326 B.n325 10.6151
R938 B.n327 B.n326 10.6151
R939 B.n327 B.n112 10.6151
R940 B.n331 B.n112 10.6151
R941 B.n332 B.n331 10.6151
R942 B.n333 B.n332 10.6151
R943 B.n333 B.n110 10.6151
R944 B.n337 B.n110 10.6151
R945 B.n338 B.n337 10.6151
R946 B.n339 B.n338 10.6151
R947 B.n339 B.n108 10.6151
R948 B.n343 B.n108 10.6151
R949 B.n344 B.n343 10.6151
R950 B.n345 B.n344 10.6151
R951 B.n345 B.n106 10.6151
R952 B.n349 B.n106 10.6151
R953 B.n350 B.n349 10.6151
R954 B.n351 B.n350 10.6151
R955 B.n351 B.n104 10.6151
R956 B.n355 B.n104 10.6151
R957 B.n356 B.n355 10.6151
R958 B.n357 B.n356 10.6151
R959 B.n357 B.n102 10.6151
R960 B.n361 B.n102 10.6151
R961 B.n362 B.n361 10.6151
R962 B.n363 B.n362 10.6151
R963 B.n363 B.n100 10.6151
R964 B.n367 B.n100 10.6151
R965 B.n368 B.n367 10.6151
R966 B.n369 B.n368 10.6151
R967 B.n369 B.n98 10.6151
R968 B.n373 B.n98 10.6151
R969 B.n374 B.n373 10.6151
R970 B.n375 B.n374 10.6151
R971 B.n375 B.n96 10.6151
R972 B.n537 B.n536 9.36635
R973 B.n519 B.n48 9.36635
R974 B.n278 B.n277 9.36635
R975 B.n296 B.n295 9.36635
R976 B.n649 B.n0 8.11757
R977 B.n649 B.n1 8.11757
R978 B.n536 B.n535 1.24928
R979 B.n522 B.n48 1.24928
R980 B.n277 B.n130 1.24928
R981 B.n295 B.n294 1.24928
R982 VP.n0 VP.t3 483.103
R983 VP.n0 VP.t1 483.017
R984 VP.n2 VP.t2 464.497
R985 VP.n3 VP.t0 464.497
R986 VP.n4 VP.n3 80.6037
R987 VP.n2 VP.n1 80.6037
R988 VP.n1 VP.n0 76.0183
R989 VP.n3 VP.n2 48.2005
R990 VP.n4 VP.n1 0.380177
R991 VP VP.n4 0.146778
R992 VTAIL.n746 VTAIL.n658 756.745
R993 VTAIL.n88 VTAIL.n0 756.745
R994 VTAIL.n182 VTAIL.n94 756.745
R995 VTAIL.n276 VTAIL.n188 756.745
R996 VTAIL.n652 VTAIL.n564 756.745
R997 VTAIL.n558 VTAIL.n470 756.745
R998 VTAIL.n464 VTAIL.n376 756.745
R999 VTAIL.n370 VTAIL.n282 756.745
R1000 VTAIL.n689 VTAIL.n688 585
R1001 VTAIL.n686 VTAIL.n685 585
R1002 VTAIL.n695 VTAIL.n694 585
R1003 VTAIL.n697 VTAIL.n696 585
R1004 VTAIL.n682 VTAIL.n681 585
R1005 VTAIL.n703 VTAIL.n702 585
R1006 VTAIL.n705 VTAIL.n704 585
R1007 VTAIL.n678 VTAIL.n677 585
R1008 VTAIL.n711 VTAIL.n710 585
R1009 VTAIL.n713 VTAIL.n712 585
R1010 VTAIL.n674 VTAIL.n673 585
R1011 VTAIL.n719 VTAIL.n718 585
R1012 VTAIL.n721 VTAIL.n720 585
R1013 VTAIL.n670 VTAIL.n669 585
R1014 VTAIL.n727 VTAIL.n726 585
R1015 VTAIL.n730 VTAIL.n729 585
R1016 VTAIL.n728 VTAIL.n666 585
R1017 VTAIL.n735 VTAIL.n665 585
R1018 VTAIL.n737 VTAIL.n736 585
R1019 VTAIL.n739 VTAIL.n738 585
R1020 VTAIL.n662 VTAIL.n661 585
R1021 VTAIL.n745 VTAIL.n744 585
R1022 VTAIL.n747 VTAIL.n746 585
R1023 VTAIL.n31 VTAIL.n30 585
R1024 VTAIL.n28 VTAIL.n27 585
R1025 VTAIL.n37 VTAIL.n36 585
R1026 VTAIL.n39 VTAIL.n38 585
R1027 VTAIL.n24 VTAIL.n23 585
R1028 VTAIL.n45 VTAIL.n44 585
R1029 VTAIL.n47 VTAIL.n46 585
R1030 VTAIL.n20 VTAIL.n19 585
R1031 VTAIL.n53 VTAIL.n52 585
R1032 VTAIL.n55 VTAIL.n54 585
R1033 VTAIL.n16 VTAIL.n15 585
R1034 VTAIL.n61 VTAIL.n60 585
R1035 VTAIL.n63 VTAIL.n62 585
R1036 VTAIL.n12 VTAIL.n11 585
R1037 VTAIL.n69 VTAIL.n68 585
R1038 VTAIL.n72 VTAIL.n71 585
R1039 VTAIL.n70 VTAIL.n8 585
R1040 VTAIL.n77 VTAIL.n7 585
R1041 VTAIL.n79 VTAIL.n78 585
R1042 VTAIL.n81 VTAIL.n80 585
R1043 VTAIL.n4 VTAIL.n3 585
R1044 VTAIL.n87 VTAIL.n86 585
R1045 VTAIL.n89 VTAIL.n88 585
R1046 VTAIL.n125 VTAIL.n124 585
R1047 VTAIL.n122 VTAIL.n121 585
R1048 VTAIL.n131 VTAIL.n130 585
R1049 VTAIL.n133 VTAIL.n132 585
R1050 VTAIL.n118 VTAIL.n117 585
R1051 VTAIL.n139 VTAIL.n138 585
R1052 VTAIL.n141 VTAIL.n140 585
R1053 VTAIL.n114 VTAIL.n113 585
R1054 VTAIL.n147 VTAIL.n146 585
R1055 VTAIL.n149 VTAIL.n148 585
R1056 VTAIL.n110 VTAIL.n109 585
R1057 VTAIL.n155 VTAIL.n154 585
R1058 VTAIL.n157 VTAIL.n156 585
R1059 VTAIL.n106 VTAIL.n105 585
R1060 VTAIL.n163 VTAIL.n162 585
R1061 VTAIL.n166 VTAIL.n165 585
R1062 VTAIL.n164 VTAIL.n102 585
R1063 VTAIL.n171 VTAIL.n101 585
R1064 VTAIL.n173 VTAIL.n172 585
R1065 VTAIL.n175 VTAIL.n174 585
R1066 VTAIL.n98 VTAIL.n97 585
R1067 VTAIL.n181 VTAIL.n180 585
R1068 VTAIL.n183 VTAIL.n182 585
R1069 VTAIL.n219 VTAIL.n218 585
R1070 VTAIL.n216 VTAIL.n215 585
R1071 VTAIL.n225 VTAIL.n224 585
R1072 VTAIL.n227 VTAIL.n226 585
R1073 VTAIL.n212 VTAIL.n211 585
R1074 VTAIL.n233 VTAIL.n232 585
R1075 VTAIL.n235 VTAIL.n234 585
R1076 VTAIL.n208 VTAIL.n207 585
R1077 VTAIL.n241 VTAIL.n240 585
R1078 VTAIL.n243 VTAIL.n242 585
R1079 VTAIL.n204 VTAIL.n203 585
R1080 VTAIL.n249 VTAIL.n248 585
R1081 VTAIL.n251 VTAIL.n250 585
R1082 VTAIL.n200 VTAIL.n199 585
R1083 VTAIL.n257 VTAIL.n256 585
R1084 VTAIL.n260 VTAIL.n259 585
R1085 VTAIL.n258 VTAIL.n196 585
R1086 VTAIL.n265 VTAIL.n195 585
R1087 VTAIL.n267 VTAIL.n266 585
R1088 VTAIL.n269 VTAIL.n268 585
R1089 VTAIL.n192 VTAIL.n191 585
R1090 VTAIL.n275 VTAIL.n274 585
R1091 VTAIL.n277 VTAIL.n276 585
R1092 VTAIL.n653 VTAIL.n652 585
R1093 VTAIL.n651 VTAIL.n650 585
R1094 VTAIL.n568 VTAIL.n567 585
R1095 VTAIL.n645 VTAIL.n644 585
R1096 VTAIL.n643 VTAIL.n642 585
R1097 VTAIL.n641 VTAIL.n571 585
R1098 VTAIL.n575 VTAIL.n572 585
R1099 VTAIL.n636 VTAIL.n635 585
R1100 VTAIL.n634 VTAIL.n633 585
R1101 VTAIL.n577 VTAIL.n576 585
R1102 VTAIL.n628 VTAIL.n627 585
R1103 VTAIL.n626 VTAIL.n625 585
R1104 VTAIL.n581 VTAIL.n580 585
R1105 VTAIL.n620 VTAIL.n619 585
R1106 VTAIL.n618 VTAIL.n617 585
R1107 VTAIL.n585 VTAIL.n584 585
R1108 VTAIL.n612 VTAIL.n611 585
R1109 VTAIL.n610 VTAIL.n609 585
R1110 VTAIL.n589 VTAIL.n588 585
R1111 VTAIL.n604 VTAIL.n603 585
R1112 VTAIL.n602 VTAIL.n601 585
R1113 VTAIL.n593 VTAIL.n592 585
R1114 VTAIL.n596 VTAIL.n595 585
R1115 VTAIL.n559 VTAIL.n558 585
R1116 VTAIL.n557 VTAIL.n556 585
R1117 VTAIL.n474 VTAIL.n473 585
R1118 VTAIL.n551 VTAIL.n550 585
R1119 VTAIL.n549 VTAIL.n548 585
R1120 VTAIL.n547 VTAIL.n477 585
R1121 VTAIL.n481 VTAIL.n478 585
R1122 VTAIL.n542 VTAIL.n541 585
R1123 VTAIL.n540 VTAIL.n539 585
R1124 VTAIL.n483 VTAIL.n482 585
R1125 VTAIL.n534 VTAIL.n533 585
R1126 VTAIL.n532 VTAIL.n531 585
R1127 VTAIL.n487 VTAIL.n486 585
R1128 VTAIL.n526 VTAIL.n525 585
R1129 VTAIL.n524 VTAIL.n523 585
R1130 VTAIL.n491 VTAIL.n490 585
R1131 VTAIL.n518 VTAIL.n517 585
R1132 VTAIL.n516 VTAIL.n515 585
R1133 VTAIL.n495 VTAIL.n494 585
R1134 VTAIL.n510 VTAIL.n509 585
R1135 VTAIL.n508 VTAIL.n507 585
R1136 VTAIL.n499 VTAIL.n498 585
R1137 VTAIL.n502 VTAIL.n501 585
R1138 VTAIL.n465 VTAIL.n464 585
R1139 VTAIL.n463 VTAIL.n462 585
R1140 VTAIL.n380 VTAIL.n379 585
R1141 VTAIL.n457 VTAIL.n456 585
R1142 VTAIL.n455 VTAIL.n454 585
R1143 VTAIL.n453 VTAIL.n383 585
R1144 VTAIL.n387 VTAIL.n384 585
R1145 VTAIL.n448 VTAIL.n447 585
R1146 VTAIL.n446 VTAIL.n445 585
R1147 VTAIL.n389 VTAIL.n388 585
R1148 VTAIL.n440 VTAIL.n439 585
R1149 VTAIL.n438 VTAIL.n437 585
R1150 VTAIL.n393 VTAIL.n392 585
R1151 VTAIL.n432 VTAIL.n431 585
R1152 VTAIL.n430 VTAIL.n429 585
R1153 VTAIL.n397 VTAIL.n396 585
R1154 VTAIL.n424 VTAIL.n423 585
R1155 VTAIL.n422 VTAIL.n421 585
R1156 VTAIL.n401 VTAIL.n400 585
R1157 VTAIL.n416 VTAIL.n415 585
R1158 VTAIL.n414 VTAIL.n413 585
R1159 VTAIL.n405 VTAIL.n404 585
R1160 VTAIL.n408 VTAIL.n407 585
R1161 VTAIL.n371 VTAIL.n370 585
R1162 VTAIL.n369 VTAIL.n368 585
R1163 VTAIL.n286 VTAIL.n285 585
R1164 VTAIL.n363 VTAIL.n362 585
R1165 VTAIL.n361 VTAIL.n360 585
R1166 VTAIL.n359 VTAIL.n289 585
R1167 VTAIL.n293 VTAIL.n290 585
R1168 VTAIL.n354 VTAIL.n353 585
R1169 VTAIL.n352 VTAIL.n351 585
R1170 VTAIL.n295 VTAIL.n294 585
R1171 VTAIL.n346 VTAIL.n345 585
R1172 VTAIL.n344 VTAIL.n343 585
R1173 VTAIL.n299 VTAIL.n298 585
R1174 VTAIL.n338 VTAIL.n337 585
R1175 VTAIL.n336 VTAIL.n335 585
R1176 VTAIL.n303 VTAIL.n302 585
R1177 VTAIL.n330 VTAIL.n329 585
R1178 VTAIL.n328 VTAIL.n327 585
R1179 VTAIL.n307 VTAIL.n306 585
R1180 VTAIL.n322 VTAIL.n321 585
R1181 VTAIL.n320 VTAIL.n319 585
R1182 VTAIL.n311 VTAIL.n310 585
R1183 VTAIL.n314 VTAIL.n313 585
R1184 VTAIL.t5 VTAIL.n594 327.466
R1185 VTAIL.t6 VTAIL.n500 327.466
R1186 VTAIL.t2 VTAIL.n406 327.466
R1187 VTAIL.t3 VTAIL.n312 327.466
R1188 VTAIL.t0 VTAIL.n687 327.466
R1189 VTAIL.t1 VTAIL.n29 327.466
R1190 VTAIL.t7 VTAIL.n123 327.466
R1191 VTAIL.t4 VTAIL.n217 327.466
R1192 VTAIL.n688 VTAIL.n685 171.744
R1193 VTAIL.n695 VTAIL.n685 171.744
R1194 VTAIL.n696 VTAIL.n695 171.744
R1195 VTAIL.n696 VTAIL.n681 171.744
R1196 VTAIL.n703 VTAIL.n681 171.744
R1197 VTAIL.n704 VTAIL.n703 171.744
R1198 VTAIL.n704 VTAIL.n677 171.744
R1199 VTAIL.n711 VTAIL.n677 171.744
R1200 VTAIL.n712 VTAIL.n711 171.744
R1201 VTAIL.n712 VTAIL.n673 171.744
R1202 VTAIL.n719 VTAIL.n673 171.744
R1203 VTAIL.n720 VTAIL.n719 171.744
R1204 VTAIL.n720 VTAIL.n669 171.744
R1205 VTAIL.n727 VTAIL.n669 171.744
R1206 VTAIL.n729 VTAIL.n727 171.744
R1207 VTAIL.n729 VTAIL.n728 171.744
R1208 VTAIL.n728 VTAIL.n665 171.744
R1209 VTAIL.n737 VTAIL.n665 171.744
R1210 VTAIL.n738 VTAIL.n737 171.744
R1211 VTAIL.n738 VTAIL.n661 171.744
R1212 VTAIL.n745 VTAIL.n661 171.744
R1213 VTAIL.n746 VTAIL.n745 171.744
R1214 VTAIL.n30 VTAIL.n27 171.744
R1215 VTAIL.n37 VTAIL.n27 171.744
R1216 VTAIL.n38 VTAIL.n37 171.744
R1217 VTAIL.n38 VTAIL.n23 171.744
R1218 VTAIL.n45 VTAIL.n23 171.744
R1219 VTAIL.n46 VTAIL.n45 171.744
R1220 VTAIL.n46 VTAIL.n19 171.744
R1221 VTAIL.n53 VTAIL.n19 171.744
R1222 VTAIL.n54 VTAIL.n53 171.744
R1223 VTAIL.n54 VTAIL.n15 171.744
R1224 VTAIL.n61 VTAIL.n15 171.744
R1225 VTAIL.n62 VTAIL.n61 171.744
R1226 VTAIL.n62 VTAIL.n11 171.744
R1227 VTAIL.n69 VTAIL.n11 171.744
R1228 VTAIL.n71 VTAIL.n69 171.744
R1229 VTAIL.n71 VTAIL.n70 171.744
R1230 VTAIL.n70 VTAIL.n7 171.744
R1231 VTAIL.n79 VTAIL.n7 171.744
R1232 VTAIL.n80 VTAIL.n79 171.744
R1233 VTAIL.n80 VTAIL.n3 171.744
R1234 VTAIL.n87 VTAIL.n3 171.744
R1235 VTAIL.n88 VTAIL.n87 171.744
R1236 VTAIL.n124 VTAIL.n121 171.744
R1237 VTAIL.n131 VTAIL.n121 171.744
R1238 VTAIL.n132 VTAIL.n131 171.744
R1239 VTAIL.n132 VTAIL.n117 171.744
R1240 VTAIL.n139 VTAIL.n117 171.744
R1241 VTAIL.n140 VTAIL.n139 171.744
R1242 VTAIL.n140 VTAIL.n113 171.744
R1243 VTAIL.n147 VTAIL.n113 171.744
R1244 VTAIL.n148 VTAIL.n147 171.744
R1245 VTAIL.n148 VTAIL.n109 171.744
R1246 VTAIL.n155 VTAIL.n109 171.744
R1247 VTAIL.n156 VTAIL.n155 171.744
R1248 VTAIL.n156 VTAIL.n105 171.744
R1249 VTAIL.n163 VTAIL.n105 171.744
R1250 VTAIL.n165 VTAIL.n163 171.744
R1251 VTAIL.n165 VTAIL.n164 171.744
R1252 VTAIL.n164 VTAIL.n101 171.744
R1253 VTAIL.n173 VTAIL.n101 171.744
R1254 VTAIL.n174 VTAIL.n173 171.744
R1255 VTAIL.n174 VTAIL.n97 171.744
R1256 VTAIL.n181 VTAIL.n97 171.744
R1257 VTAIL.n182 VTAIL.n181 171.744
R1258 VTAIL.n218 VTAIL.n215 171.744
R1259 VTAIL.n225 VTAIL.n215 171.744
R1260 VTAIL.n226 VTAIL.n225 171.744
R1261 VTAIL.n226 VTAIL.n211 171.744
R1262 VTAIL.n233 VTAIL.n211 171.744
R1263 VTAIL.n234 VTAIL.n233 171.744
R1264 VTAIL.n234 VTAIL.n207 171.744
R1265 VTAIL.n241 VTAIL.n207 171.744
R1266 VTAIL.n242 VTAIL.n241 171.744
R1267 VTAIL.n242 VTAIL.n203 171.744
R1268 VTAIL.n249 VTAIL.n203 171.744
R1269 VTAIL.n250 VTAIL.n249 171.744
R1270 VTAIL.n250 VTAIL.n199 171.744
R1271 VTAIL.n257 VTAIL.n199 171.744
R1272 VTAIL.n259 VTAIL.n257 171.744
R1273 VTAIL.n259 VTAIL.n258 171.744
R1274 VTAIL.n258 VTAIL.n195 171.744
R1275 VTAIL.n267 VTAIL.n195 171.744
R1276 VTAIL.n268 VTAIL.n267 171.744
R1277 VTAIL.n268 VTAIL.n191 171.744
R1278 VTAIL.n275 VTAIL.n191 171.744
R1279 VTAIL.n276 VTAIL.n275 171.744
R1280 VTAIL.n652 VTAIL.n651 171.744
R1281 VTAIL.n651 VTAIL.n567 171.744
R1282 VTAIL.n644 VTAIL.n567 171.744
R1283 VTAIL.n644 VTAIL.n643 171.744
R1284 VTAIL.n643 VTAIL.n571 171.744
R1285 VTAIL.n575 VTAIL.n571 171.744
R1286 VTAIL.n635 VTAIL.n575 171.744
R1287 VTAIL.n635 VTAIL.n634 171.744
R1288 VTAIL.n634 VTAIL.n576 171.744
R1289 VTAIL.n627 VTAIL.n576 171.744
R1290 VTAIL.n627 VTAIL.n626 171.744
R1291 VTAIL.n626 VTAIL.n580 171.744
R1292 VTAIL.n619 VTAIL.n580 171.744
R1293 VTAIL.n619 VTAIL.n618 171.744
R1294 VTAIL.n618 VTAIL.n584 171.744
R1295 VTAIL.n611 VTAIL.n584 171.744
R1296 VTAIL.n611 VTAIL.n610 171.744
R1297 VTAIL.n610 VTAIL.n588 171.744
R1298 VTAIL.n603 VTAIL.n588 171.744
R1299 VTAIL.n603 VTAIL.n602 171.744
R1300 VTAIL.n602 VTAIL.n592 171.744
R1301 VTAIL.n595 VTAIL.n592 171.744
R1302 VTAIL.n558 VTAIL.n557 171.744
R1303 VTAIL.n557 VTAIL.n473 171.744
R1304 VTAIL.n550 VTAIL.n473 171.744
R1305 VTAIL.n550 VTAIL.n549 171.744
R1306 VTAIL.n549 VTAIL.n477 171.744
R1307 VTAIL.n481 VTAIL.n477 171.744
R1308 VTAIL.n541 VTAIL.n481 171.744
R1309 VTAIL.n541 VTAIL.n540 171.744
R1310 VTAIL.n540 VTAIL.n482 171.744
R1311 VTAIL.n533 VTAIL.n482 171.744
R1312 VTAIL.n533 VTAIL.n532 171.744
R1313 VTAIL.n532 VTAIL.n486 171.744
R1314 VTAIL.n525 VTAIL.n486 171.744
R1315 VTAIL.n525 VTAIL.n524 171.744
R1316 VTAIL.n524 VTAIL.n490 171.744
R1317 VTAIL.n517 VTAIL.n490 171.744
R1318 VTAIL.n517 VTAIL.n516 171.744
R1319 VTAIL.n516 VTAIL.n494 171.744
R1320 VTAIL.n509 VTAIL.n494 171.744
R1321 VTAIL.n509 VTAIL.n508 171.744
R1322 VTAIL.n508 VTAIL.n498 171.744
R1323 VTAIL.n501 VTAIL.n498 171.744
R1324 VTAIL.n464 VTAIL.n463 171.744
R1325 VTAIL.n463 VTAIL.n379 171.744
R1326 VTAIL.n456 VTAIL.n379 171.744
R1327 VTAIL.n456 VTAIL.n455 171.744
R1328 VTAIL.n455 VTAIL.n383 171.744
R1329 VTAIL.n387 VTAIL.n383 171.744
R1330 VTAIL.n447 VTAIL.n387 171.744
R1331 VTAIL.n447 VTAIL.n446 171.744
R1332 VTAIL.n446 VTAIL.n388 171.744
R1333 VTAIL.n439 VTAIL.n388 171.744
R1334 VTAIL.n439 VTAIL.n438 171.744
R1335 VTAIL.n438 VTAIL.n392 171.744
R1336 VTAIL.n431 VTAIL.n392 171.744
R1337 VTAIL.n431 VTAIL.n430 171.744
R1338 VTAIL.n430 VTAIL.n396 171.744
R1339 VTAIL.n423 VTAIL.n396 171.744
R1340 VTAIL.n423 VTAIL.n422 171.744
R1341 VTAIL.n422 VTAIL.n400 171.744
R1342 VTAIL.n415 VTAIL.n400 171.744
R1343 VTAIL.n415 VTAIL.n414 171.744
R1344 VTAIL.n414 VTAIL.n404 171.744
R1345 VTAIL.n407 VTAIL.n404 171.744
R1346 VTAIL.n370 VTAIL.n369 171.744
R1347 VTAIL.n369 VTAIL.n285 171.744
R1348 VTAIL.n362 VTAIL.n285 171.744
R1349 VTAIL.n362 VTAIL.n361 171.744
R1350 VTAIL.n361 VTAIL.n289 171.744
R1351 VTAIL.n293 VTAIL.n289 171.744
R1352 VTAIL.n353 VTAIL.n293 171.744
R1353 VTAIL.n353 VTAIL.n352 171.744
R1354 VTAIL.n352 VTAIL.n294 171.744
R1355 VTAIL.n345 VTAIL.n294 171.744
R1356 VTAIL.n345 VTAIL.n344 171.744
R1357 VTAIL.n344 VTAIL.n298 171.744
R1358 VTAIL.n337 VTAIL.n298 171.744
R1359 VTAIL.n337 VTAIL.n336 171.744
R1360 VTAIL.n336 VTAIL.n302 171.744
R1361 VTAIL.n329 VTAIL.n302 171.744
R1362 VTAIL.n329 VTAIL.n328 171.744
R1363 VTAIL.n328 VTAIL.n306 171.744
R1364 VTAIL.n321 VTAIL.n306 171.744
R1365 VTAIL.n321 VTAIL.n320 171.744
R1366 VTAIL.n320 VTAIL.n310 171.744
R1367 VTAIL.n313 VTAIL.n310 171.744
R1368 VTAIL.n688 VTAIL.t0 85.8723
R1369 VTAIL.n30 VTAIL.t1 85.8723
R1370 VTAIL.n124 VTAIL.t7 85.8723
R1371 VTAIL.n218 VTAIL.t4 85.8723
R1372 VTAIL.n595 VTAIL.t5 85.8723
R1373 VTAIL.n501 VTAIL.t6 85.8723
R1374 VTAIL.n407 VTAIL.t2 85.8723
R1375 VTAIL.n313 VTAIL.t3 85.8723
R1376 VTAIL.n751 VTAIL.n750 29.8581
R1377 VTAIL.n93 VTAIL.n92 29.8581
R1378 VTAIL.n187 VTAIL.n186 29.8581
R1379 VTAIL.n281 VTAIL.n280 29.8581
R1380 VTAIL.n657 VTAIL.n656 29.8581
R1381 VTAIL.n563 VTAIL.n562 29.8581
R1382 VTAIL.n469 VTAIL.n468 29.8581
R1383 VTAIL.n375 VTAIL.n374 29.8581
R1384 VTAIL.n751 VTAIL.n657 27.8496
R1385 VTAIL.n375 VTAIL.n281 27.8496
R1386 VTAIL.n689 VTAIL.n687 16.3895
R1387 VTAIL.n31 VTAIL.n29 16.3895
R1388 VTAIL.n125 VTAIL.n123 16.3895
R1389 VTAIL.n219 VTAIL.n217 16.3895
R1390 VTAIL.n596 VTAIL.n594 16.3895
R1391 VTAIL.n502 VTAIL.n500 16.3895
R1392 VTAIL.n408 VTAIL.n406 16.3895
R1393 VTAIL.n314 VTAIL.n312 16.3895
R1394 VTAIL.n736 VTAIL.n735 13.1884
R1395 VTAIL.n78 VTAIL.n77 13.1884
R1396 VTAIL.n172 VTAIL.n171 13.1884
R1397 VTAIL.n266 VTAIL.n265 13.1884
R1398 VTAIL.n642 VTAIL.n641 13.1884
R1399 VTAIL.n548 VTAIL.n547 13.1884
R1400 VTAIL.n454 VTAIL.n453 13.1884
R1401 VTAIL.n360 VTAIL.n359 13.1884
R1402 VTAIL.n690 VTAIL.n686 12.8005
R1403 VTAIL.n734 VTAIL.n666 12.8005
R1404 VTAIL.n739 VTAIL.n664 12.8005
R1405 VTAIL.n32 VTAIL.n28 12.8005
R1406 VTAIL.n76 VTAIL.n8 12.8005
R1407 VTAIL.n81 VTAIL.n6 12.8005
R1408 VTAIL.n126 VTAIL.n122 12.8005
R1409 VTAIL.n170 VTAIL.n102 12.8005
R1410 VTAIL.n175 VTAIL.n100 12.8005
R1411 VTAIL.n220 VTAIL.n216 12.8005
R1412 VTAIL.n264 VTAIL.n196 12.8005
R1413 VTAIL.n269 VTAIL.n194 12.8005
R1414 VTAIL.n645 VTAIL.n570 12.8005
R1415 VTAIL.n640 VTAIL.n572 12.8005
R1416 VTAIL.n597 VTAIL.n593 12.8005
R1417 VTAIL.n551 VTAIL.n476 12.8005
R1418 VTAIL.n546 VTAIL.n478 12.8005
R1419 VTAIL.n503 VTAIL.n499 12.8005
R1420 VTAIL.n457 VTAIL.n382 12.8005
R1421 VTAIL.n452 VTAIL.n384 12.8005
R1422 VTAIL.n409 VTAIL.n405 12.8005
R1423 VTAIL.n363 VTAIL.n288 12.8005
R1424 VTAIL.n358 VTAIL.n290 12.8005
R1425 VTAIL.n315 VTAIL.n311 12.8005
R1426 VTAIL.n694 VTAIL.n693 12.0247
R1427 VTAIL.n731 VTAIL.n730 12.0247
R1428 VTAIL.n740 VTAIL.n662 12.0247
R1429 VTAIL.n36 VTAIL.n35 12.0247
R1430 VTAIL.n73 VTAIL.n72 12.0247
R1431 VTAIL.n82 VTAIL.n4 12.0247
R1432 VTAIL.n130 VTAIL.n129 12.0247
R1433 VTAIL.n167 VTAIL.n166 12.0247
R1434 VTAIL.n176 VTAIL.n98 12.0247
R1435 VTAIL.n224 VTAIL.n223 12.0247
R1436 VTAIL.n261 VTAIL.n260 12.0247
R1437 VTAIL.n270 VTAIL.n192 12.0247
R1438 VTAIL.n646 VTAIL.n568 12.0247
R1439 VTAIL.n637 VTAIL.n636 12.0247
R1440 VTAIL.n601 VTAIL.n600 12.0247
R1441 VTAIL.n552 VTAIL.n474 12.0247
R1442 VTAIL.n543 VTAIL.n542 12.0247
R1443 VTAIL.n507 VTAIL.n506 12.0247
R1444 VTAIL.n458 VTAIL.n380 12.0247
R1445 VTAIL.n449 VTAIL.n448 12.0247
R1446 VTAIL.n413 VTAIL.n412 12.0247
R1447 VTAIL.n364 VTAIL.n286 12.0247
R1448 VTAIL.n355 VTAIL.n354 12.0247
R1449 VTAIL.n319 VTAIL.n318 12.0247
R1450 VTAIL.n697 VTAIL.n684 11.249
R1451 VTAIL.n726 VTAIL.n668 11.249
R1452 VTAIL.n744 VTAIL.n743 11.249
R1453 VTAIL.n39 VTAIL.n26 11.249
R1454 VTAIL.n68 VTAIL.n10 11.249
R1455 VTAIL.n86 VTAIL.n85 11.249
R1456 VTAIL.n133 VTAIL.n120 11.249
R1457 VTAIL.n162 VTAIL.n104 11.249
R1458 VTAIL.n180 VTAIL.n179 11.249
R1459 VTAIL.n227 VTAIL.n214 11.249
R1460 VTAIL.n256 VTAIL.n198 11.249
R1461 VTAIL.n274 VTAIL.n273 11.249
R1462 VTAIL.n650 VTAIL.n649 11.249
R1463 VTAIL.n633 VTAIL.n574 11.249
R1464 VTAIL.n604 VTAIL.n591 11.249
R1465 VTAIL.n556 VTAIL.n555 11.249
R1466 VTAIL.n539 VTAIL.n480 11.249
R1467 VTAIL.n510 VTAIL.n497 11.249
R1468 VTAIL.n462 VTAIL.n461 11.249
R1469 VTAIL.n445 VTAIL.n386 11.249
R1470 VTAIL.n416 VTAIL.n403 11.249
R1471 VTAIL.n368 VTAIL.n367 11.249
R1472 VTAIL.n351 VTAIL.n292 11.249
R1473 VTAIL.n322 VTAIL.n309 11.249
R1474 VTAIL.n698 VTAIL.n682 10.4732
R1475 VTAIL.n725 VTAIL.n670 10.4732
R1476 VTAIL.n747 VTAIL.n660 10.4732
R1477 VTAIL.n40 VTAIL.n24 10.4732
R1478 VTAIL.n67 VTAIL.n12 10.4732
R1479 VTAIL.n89 VTAIL.n2 10.4732
R1480 VTAIL.n134 VTAIL.n118 10.4732
R1481 VTAIL.n161 VTAIL.n106 10.4732
R1482 VTAIL.n183 VTAIL.n96 10.4732
R1483 VTAIL.n228 VTAIL.n212 10.4732
R1484 VTAIL.n255 VTAIL.n200 10.4732
R1485 VTAIL.n277 VTAIL.n190 10.4732
R1486 VTAIL.n653 VTAIL.n566 10.4732
R1487 VTAIL.n632 VTAIL.n577 10.4732
R1488 VTAIL.n605 VTAIL.n589 10.4732
R1489 VTAIL.n559 VTAIL.n472 10.4732
R1490 VTAIL.n538 VTAIL.n483 10.4732
R1491 VTAIL.n511 VTAIL.n495 10.4732
R1492 VTAIL.n465 VTAIL.n378 10.4732
R1493 VTAIL.n444 VTAIL.n389 10.4732
R1494 VTAIL.n417 VTAIL.n401 10.4732
R1495 VTAIL.n371 VTAIL.n284 10.4732
R1496 VTAIL.n350 VTAIL.n295 10.4732
R1497 VTAIL.n323 VTAIL.n307 10.4732
R1498 VTAIL.n702 VTAIL.n701 9.69747
R1499 VTAIL.n722 VTAIL.n721 9.69747
R1500 VTAIL.n748 VTAIL.n658 9.69747
R1501 VTAIL.n44 VTAIL.n43 9.69747
R1502 VTAIL.n64 VTAIL.n63 9.69747
R1503 VTAIL.n90 VTAIL.n0 9.69747
R1504 VTAIL.n138 VTAIL.n137 9.69747
R1505 VTAIL.n158 VTAIL.n157 9.69747
R1506 VTAIL.n184 VTAIL.n94 9.69747
R1507 VTAIL.n232 VTAIL.n231 9.69747
R1508 VTAIL.n252 VTAIL.n251 9.69747
R1509 VTAIL.n278 VTAIL.n188 9.69747
R1510 VTAIL.n654 VTAIL.n564 9.69747
R1511 VTAIL.n629 VTAIL.n628 9.69747
R1512 VTAIL.n609 VTAIL.n608 9.69747
R1513 VTAIL.n560 VTAIL.n470 9.69747
R1514 VTAIL.n535 VTAIL.n534 9.69747
R1515 VTAIL.n515 VTAIL.n514 9.69747
R1516 VTAIL.n466 VTAIL.n376 9.69747
R1517 VTAIL.n441 VTAIL.n440 9.69747
R1518 VTAIL.n421 VTAIL.n420 9.69747
R1519 VTAIL.n372 VTAIL.n282 9.69747
R1520 VTAIL.n347 VTAIL.n346 9.69747
R1521 VTAIL.n327 VTAIL.n326 9.69747
R1522 VTAIL.n750 VTAIL.n749 9.45567
R1523 VTAIL.n92 VTAIL.n91 9.45567
R1524 VTAIL.n186 VTAIL.n185 9.45567
R1525 VTAIL.n280 VTAIL.n279 9.45567
R1526 VTAIL.n656 VTAIL.n655 9.45567
R1527 VTAIL.n562 VTAIL.n561 9.45567
R1528 VTAIL.n468 VTAIL.n467 9.45567
R1529 VTAIL.n374 VTAIL.n373 9.45567
R1530 VTAIL.n749 VTAIL.n748 9.3005
R1531 VTAIL.n660 VTAIL.n659 9.3005
R1532 VTAIL.n743 VTAIL.n742 9.3005
R1533 VTAIL.n741 VTAIL.n740 9.3005
R1534 VTAIL.n664 VTAIL.n663 9.3005
R1535 VTAIL.n709 VTAIL.n708 9.3005
R1536 VTAIL.n707 VTAIL.n706 9.3005
R1537 VTAIL.n680 VTAIL.n679 9.3005
R1538 VTAIL.n701 VTAIL.n700 9.3005
R1539 VTAIL.n699 VTAIL.n698 9.3005
R1540 VTAIL.n684 VTAIL.n683 9.3005
R1541 VTAIL.n693 VTAIL.n692 9.3005
R1542 VTAIL.n691 VTAIL.n690 9.3005
R1543 VTAIL.n676 VTAIL.n675 9.3005
R1544 VTAIL.n715 VTAIL.n714 9.3005
R1545 VTAIL.n717 VTAIL.n716 9.3005
R1546 VTAIL.n672 VTAIL.n671 9.3005
R1547 VTAIL.n723 VTAIL.n722 9.3005
R1548 VTAIL.n725 VTAIL.n724 9.3005
R1549 VTAIL.n668 VTAIL.n667 9.3005
R1550 VTAIL.n732 VTAIL.n731 9.3005
R1551 VTAIL.n734 VTAIL.n733 9.3005
R1552 VTAIL.n91 VTAIL.n90 9.3005
R1553 VTAIL.n2 VTAIL.n1 9.3005
R1554 VTAIL.n85 VTAIL.n84 9.3005
R1555 VTAIL.n83 VTAIL.n82 9.3005
R1556 VTAIL.n6 VTAIL.n5 9.3005
R1557 VTAIL.n51 VTAIL.n50 9.3005
R1558 VTAIL.n49 VTAIL.n48 9.3005
R1559 VTAIL.n22 VTAIL.n21 9.3005
R1560 VTAIL.n43 VTAIL.n42 9.3005
R1561 VTAIL.n41 VTAIL.n40 9.3005
R1562 VTAIL.n26 VTAIL.n25 9.3005
R1563 VTAIL.n35 VTAIL.n34 9.3005
R1564 VTAIL.n33 VTAIL.n32 9.3005
R1565 VTAIL.n18 VTAIL.n17 9.3005
R1566 VTAIL.n57 VTAIL.n56 9.3005
R1567 VTAIL.n59 VTAIL.n58 9.3005
R1568 VTAIL.n14 VTAIL.n13 9.3005
R1569 VTAIL.n65 VTAIL.n64 9.3005
R1570 VTAIL.n67 VTAIL.n66 9.3005
R1571 VTAIL.n10 VTAIL.n9 9.3005
R1572 VTAIL.n74 VTAIL.n73 9.3005
R1573 VTAIL.n76 VTAIL.n75 9.3005
R1574 VTAIL.n185 VTAIL.n184 9.3005
R1575 VTAIL.n96 VTAIL.n95 9.3005
R1576 VTAIL.n179 VTAIL.n178 9.3005
R1577 VTAIL.n177 VTAIL.n176 9.3005
R1578 VTAIL.n100 VTAIL.n99 9.3005
R1579 VTAIL.n145 VTAIL.n144 9.3005
R1580 VTAIL.n143 VTAIL.n142 9.3005
R1581 VTAIL.n116 VTAIL.n115 9.3005
R1582 VTAIL.n137 VTAIL.n136 9.3005
R1583 VTAIL.n135 VTAIL.n134 9.3005
R1584 VTAIL.n120 VTAIL.n119 9.3005
R1585 VTAIL.n129 VTAIL.n128 9.3005
R1586 VTAIL.n127 VTAIL.n126 9.3005
R1587 VTAIL.n112 VTAIL.n111 9.3005
R1588 VTAIL.n151 VTAIL.n150 9.3005
R1589 VTAIL.n153 VTAIL.n152 9.3005
R1590 VTAIL.n108 VTAIL.n107 9.3005
R1591 VTAIL.n159 VTAIL.n158 9.3005
R1592 VTAIL.n161 VTAIL.n160 9.3005
R1593 VTAIL.n104 VTAIL.n103 9.3005
R1594 VTAIL.n168 VTAIL.n167 9.3005
R1595 VTAIL.n170 VTAIL.n169 9.3005
R1596 VTAIL.n279 VTAIL.n278 9.3005
R1597 VTAIL.n190 VTAIL.n189 9.3005
R1598 VTAIL.n273 VTAIL.n272 9.3005
R1599 VTAIL.n271 VTAIL.n270 9.3005
R1600 VTAIL.n194 VTAIL.n193 9.3005
R1601 VTAIL.n239 VTAIL.n238 9.3005
R1602 VTAIL.n237 VTAIL.n236 9.3005
R1603 VTAIL.n210 VTAIL.n209 9.3005
R1604 VTAIL.n231 VTAIL.n230 9.3005
R1605 VTAIL.n229 VTAIL.n228 9.3005
R1606 VTAIL.n214 VTAIL.n213 9.3005
R1607 VTAIL.n223 VTAIL.n222 9.3005
R1608 VTAIL.n221 VTAIL.n220 9.3005
R1609 VTAIL.n206 VTAIL.n205 9.3005
R1610 VTAIL.n245 VTAIL.n244 9.3005
R1611 VTAIL.n247 VTAIL.n246 9.3005
R1612 VTAIL.n202 VTAIL.n201 9.3005
R1613 VTAIL.n253 VTAIL.n252 9.3005
R1614 VTAIL.n255 VTAIL.n254 9.3005
R1615 VTAIL.n198 VTAIL.n197 9.3005
R1616 VTAIL.n262 VTAIL.n261 9.3005
R1617 VTAIL.n264 VTAIL.n263 9.3005
R1618 VTAIL.n622 VTAIL.n621 9.3005
R1619 VTAIL.n624 VTAIL.n623 9.3005
R1620 VTAIL.n579 VTAIL.n578 9.3005
R1621 VTAIL.n630 VTAIL.n629 9.3005
R1622 VTAIL.n632 VTAIL.n631 9.3005
R1623 VTAIL.n574 VTAIL.n573 9.3005
R1624 VTAIL.n638 VTAIL.n637 9.3005
R1625 VTAIL.n640 VTAIL.n639 9.3005
R1626 VTAIL.n655 VTAIL.n654 9.3005
R1627 VTAIL.n566 VTAIL.n565 9.3005
R1628 VTAIL.n649 VTAIL.n648 9.3005
R1629 VTAIL.n647 VTAIL.n646 9.3005
R1630 VTAIL.n570 VTAIL.n569 9.3005
R1631 VTAIL.n583 VTAIL.n582 9.3005
R1632 VTAIL.n616 VTAIL.n615 9.3005
R1633 VTAIL.n614 VTAIL.n613 9.3005
R1634 VTAIL.n587 VTAIL.n586 9.3005
R1635 VTAIL.n608 VTAIL.n607 9.3005
R1636 VTAIL.n606 VTAIL.n605 9.3005
R1637 VTAIL.n591 VTAIL.n590 9.3005
R1638 VTAIL.n600 VTAIL.n599 9.3005
R1639 VTAIL.n598 VTAIL.n597 9.3005
R1640 VTAIL.n528 VTAIL.n527 9.3005
R1641 VTAIL.n530 VTAIL.n529 9.3005
R1642 VTAIL.n485 VTAIL.n484 9.3005
R1643 VTAIL.n536 VTAIL.n535 9.3005
R1644 VTAIL.n538 VTAIL.n537 9.3005
R1645 VTAIL.n480 VTAIL.n479 9.3005
R1646 VTAIL.n544 VTAIL.n543 9.3005
R1647 VTAIL.n546 VTAIL.n545 9.3005
R1648 VTAIL.n561 VTAIL.n560 9.3005
R1649 VTAIL.n472 VTAIL.n471 9.3005
R1650 VTAIL.n555 VTAIL.n554 9.3005
R1651 VTAIL.n553 VTAIL.n552 9.3005
R1652 VTAIL.n476 VTAIL.n475 9.3005
R1653 VTAIL.n489 VTAIL.n488 9.3005
R1654 VTAIL.n522 VTAIL.n521 9.3005
R1655 VTAIL.n520 VTAIL.n519 9.3005
R1656 VTAIL.n493 VTAIL.n492 9.3005
R1657 VTAIL.n514 VTAIL.n513 9.3005
R1658 VTAIL.n512 VTAIL.n511 9.3005
R1659 VTAIL.n497 VTAIL.n496 9.3005
R1660 VTAIL.n506 VTAIL.n505 9.3005
R1661 VTAIL.n504 VTAIL.n503 9.3005
R1662 VTAIL.n434 VTAIL.n433 9.3005
R1663 VTAIL.n436 VTAIL.n435 9.3005
R1664 VTAIL.n391 VTAIL.n390 9.3005
R1665 VTAIL.n442 VTAIL.n441 9.3005
R1666 VTAIL.n444 VTAIL.n443 9.3005
R1667 VTAIL.n386 VTAIL.n385 9.3005
R1668 VTAIL.n450 VTAIL.n449 9.3005
R1669 VTAIL.n452 VTAIL.n451 9.3005
R1670 VTAIL.n467 VTAIL.n466 9.3005
R1671 VTAIL.n378 VTAIL.n377 9.3005
R1672 VTAIL.n461 VTAIL.n460 9.3005
R1673 VTAIL.n459 VTAIL.n458 9.3005
R1674 VTAIL.n382 VTAIL.n381 9.3005
R1675 VTAIL.n395 VTAIL.n394 9.3005
R1676 VTAIL.n428 VTAIL.n427 9.3005
R1677 VTAIL.n426 VTAIL.n425 9.3005
R1678 VTAIL.n399 VTAIL.n398 9.3005
R1679 VTAIL.n420 VTAIL.n419 9.3005
R1680 VTAIL.n418 VTAIL.n417 9.3005
R1681 VTAIL.n403 VTAIL.n402 9.3005
R1682 VTAIL.n412 VTAIL.n411 9.3005
R1683 VTAIL.n410 VTAIL.n409 9.3005
R1684 VTAIL.n340 VTAIL.n339 9.3005
R1685 VTAIL.n342 VTAIL.n341 9.3005
R1686 VTAIL.n297 VTAIL.n296 9.3005
R1687 VTAIL.n348 VTAIL.n347 9.3005
R1688 VTAIL.n350 VTAIL.n349 9.3005
R1689 VTAIL.n292 VTAIL.n291 9.3005
R1690 VTAIL.n356 VTAIL.n355 9.3005
R1691 VTAIL.n358 VTAIL.n357 9.3005
R1692 VTAIL.n373 VTAIL.n372 9.3005
R1693 VTAIL.n284 VTAIL.n283 9.3005
R1694 VTAIL.n367 VTAIL.n366 9.3005
R1695 VTAIL.n365 VTAIL.n364 9.3005
R1696 VTAIL.n288 VTAIL.n287 9.3005
R1697 VTAIL.n301 VTAIL.n300 9.3005
R1698 VTAIL.n334 VTAIL.n333 9.3005
R1699 VTAIL.n332 VTAIL.n331 9.3005
R1700 VTAIL.n305 VTAIL.n304 9.3005
R1701 VTAIL.n326 VTAIL.n325 9.3005
R1702 VTAIL.n324 VTAIL.n323 9.3005
R1703 VTAIL.n309 VTAIL.n308 9.3005
R1704 VTAIL.n318 VTAIL.n317 9.3005
R1705 VTAIL.n316 VTAIL.n315 9.3005
R1706 VTAIL.n705 VTAIL.n680 8.92171
R1707 VTAIL.n718 VTAIL.n672 8.92171
R1708 VTAIL.n47 VTAIL.n22 8.92171
R1709 VTAIL.n60 VTAIL.n14 8.92171
R1710 VTAIL.n141 VTAIL.n116 8.92171
R1711 VTAIL.n154 VTAIL.n108 8.92171
R1712 VTAIL.n235 VTAIL.n210 8.92171
R1713 VTAIL.n248 VTAIL.n202 8.92171
R1714 VTAIL.n625 VTAIL.n579 8.92171
R1715 VTAIL.n612 VTAIL.n587 8.92171
R1716 VTAIL.n531 VTAIL.n485 8.92171
R1717 VTAIL.n518 VTAIL.n493 8.92171
R1718 VTAIL.n437 VTAIL.n391 8.92171
R1719 VTAIL.n424 VTAIL.n399 8.92171
R1720 VTAIL.n343 VTAIL.n297 8.92171
R1721 VTAIL.n330 VTAIL.n305 8.92171
R1722 VTAIL.n706 VTAIL.n678 8.14595
R1723 VTAIL.n717 VTAIL.n674 8.14595
R1724 VTAIL.n48 VTAIL.n20 8.14595
R1725 VTAIL.n59 VTAIL.n16 8.14595
R1726 VTAIL.n142 VTAIL.n114 8.14595
R1727 VTAIL.n153 VTAIL.n110 8.14595
R1728 VTAIL.n236 VTAIL.n208 8.14595
R1729 VTAIL.n247 VTAIL.n204 8.14595
R1730 VTAIL.n624 VTAIL.n581 8.14595
R1731 VTAIL.n613 VTAIL.n585 8.14595
R1732 VTAIL.n530 VTAIL.n487 8.14595
R1733 VTAIL.n519 VTAIL.n491 8.14595
R1734 VTAIL.n436 VTAIL.n393 8.14595
R1735 VTAIL.n425 VTAIL.n397 8.14595
R1736 VTAIL.n342 VTAIL.n299 8.14595
R1737 VTAIL.n331 VTAIL.n303 8.14595
R1738 VTAIL.n710 VTAIL.n709 7.3702
R1739 VTAIL.n714 VTAIL.n713 7.3702
R1740 VTAIL.n52 VTAIL.n51 7.3702
R1741 VTAIL.n56 VTAIL.n55 7.3702
R1742 VTAIL.n146 VTAIL.n145 7.3702
R1743 VTAIL.n150 VTAIL.n149 7.3702
R1744 VTAIL.n240 VTAIL.n239 7.3702
R1745 VTAIL.n244 VTAIL.n243 7.3702
R1746 VTAIL.n621 VTAIL.n620 7.3702
R1747 VTAIL.n617 VTAIL.n616 7.3702
R1748 VTAIL.n527 VTAIL.n526 7.3702
R1749 VTAIL.n523 VTAIL.n522 7.3702
R1750 VTAIL.n433 VTAIL.n432 7.3702
R1751 VTAIL.n429 VTAIL.n428 7.3702
R1752 VTAIL.n339 VTAIL.n338 7.3702
R1753 VTAIL.n335 VTAIL.n334 7.3702
R1754 VTAIL.n710 VTAIL.n676 6.59444
R1755 VTAIL.n713 VTAIL.n676 6.59444
R1756 VTAIL.n52 VTAIL.n18 6.59444
R1757 VTAIL.n55 VTAIL.n18 6.59444
R1758 VTAIL.n146 VTAIL.n112 6.59444
R1759 VTAIL.n149 VTAIL.n112 6.59444
R1760 VTAIL.n240 VTAIL.n206 6.59444
R1761 VTAIL.n243 VTAIL.n206 6.59444
R1762 VTAIL.n620 VTAIL.n583 6.59444
R1763 VTAIL.n617 VTAIL.n583 6.59444
R1764 VTAIL.n526 VTAIL.n489 6.59444
R1765 VTAIL.n523 VTAIL.n489 6.59444
R1766 VTAIL.n432 VTAIL.n395 6.59444
R1767 VTAIL.n429 VTAIL.n395 6.59444
R1768 VTAIL.n338 VTAIL.n301 6.59444
R1769 VTAIL.n335 VTAIL.n301 6.59444
R1770 VTAIL.n709 VTAIL.n678 5.81868
R1771 VTAIL.n714 VTAIL.n674 5.81868
R1772 VTAIL.n51 VTAIL.n20 5.81868
R1773 VTAIL.n56 VTAIL.n16 5.81868
R1774 VTAIL.n145 VTAIL.n114 5.81868
R1775 VTAIL.n150 VTAIL.n110 5.81868
R1776 VTAIL.n239 VTAIL.n208 5.81868
R1777 VTAIL.n244 VTAIL.n204 5.81868
R1778 VTAIL.n621 VTAIL.n581 5.81868
R1779 VTAIL.n616 VTAIL.n585 5.81868
R1780 VTAIL.n527 VTAIL.n487 5.81868
R1781 VTAIL.n522 VTAIL.n491 5.81868
R1782 VTAIL.n433 VTAIL.n393 5.81868
R1783 VTAIL.n428 VTAIL.n397 5.81868
R1784 VTAIL.n339 VTAIL.n299 5.81868
R1785 VTAIL.n334 VTAIL.n303 5.81868
R1786 VTAIL.n706 VTAIL.n705 5.04292
R1787 VTAIL.n718 VTAIL.n717 5.04292
R1788 VTAIL.n48 VTAIL.n47 5.04292
R1789 VTAIL.n60 VTAIL.n59 5.04292
R1790 VTAIL.n142 VTAIL.n141 5.04292
R1791 VTAIL.n154 VTAIL.n153 5.04292
R1792 VTAIL.n236 VTAIL.n235 5.04292
R1793 VTAIL.n248 VTAIL.n247 5.04292
R1794 VTAIL.n625 VTAIL.n624 5.04292
R1795 VTAIL.n613 VTAIL.n612 5.04292
R1796 VTAIL.n531 VTAIL.n530 5.04292
R1797 VTAIL.n519 VTAIL.n518 5.04292
R1798 VTAIL.n437 VTAIL.n436 5.04292
R1799 VTAIL.n425 VTAIL.n424 5.04292
R1800 VTAIL.n343 VTAIL.n342 5.04292
R1801 VTAIL.n331 VTAIL.n330 5.04292
R1802 VTAIL.n702 VTAIL.n680 4.26717
R1803 VTAIL.n721 VTAIL.n672 4.26717
R1804 VTAIL.n750 VTAIL.n658 4.26717
R1805 VTAIL.n44 VTAIL.n22 4.26717
R1806 VTAIL.n63 VTAIL.n14 4.26717
R1807 VTAIL.n92 VTAIL.n0 4.26717
R1808 VTAIL.n138 VTAIL.n116 4.26717
R1809 VTAIL.n157 VTAIL.n108 4.26717
R1810 VTAIL.n186 VTAIL.n94 4.26717
R1811 VTAIL.n232 VTAIL.n210 4.26717
R1812 VTAIL.n251 VTAIL.n202 4.26717
R1813 VTAIL.n280 VTAIL.n188 4.26717
R1814 VTAIL.n656 VTAIL.n564 4.26717
R1815 VTAIL.n628 VTAIL.n579 4.26717
R1816 VTAIL.n609 VTAIL.n587 4.26717
R1817 VTAIL.n562 VTAIL.n470 4.26717
R1818 VTAIL.n534 VTAIL.n485 4.26717
R1819 VTAIL.n515 VTAIL.n493 4.26717
R1820 VTAIL.n468 VTAIL.n376 4.26717
R1821 VTAIL.n440 VTAIL.n391 4.26717
R1822 VTAIL.n421 VTAIL.n399 4.26717
R1823 VTAIL.n374 VTAIL.n282 4.26717
R1824 VTAIL.n346 VTAIL.n297 4.26717
R1825 VTAIL.n327 VTAIL.n305 4.26717
R1826 VTAIL.n691 VTAIL.n687 3.70982
R1827 VTAIL.n33 VTAIL.n29 3.70982
R1828 VTAIL.n127 VTAIL.n123 3.70982
R1829 VTAIL.n221 VTAIL.n217 3.70982
R1830 VTAIL.n598 VTAIL.n594 3.70982
R1831 VTAIL.n504 VTAIL.n500 3.70982
R1832 VTAIL.n410 VTAIL.n406 3.70982
R1833 VTAIL.n316 VTAIL.n312 3.70982
R1834 VTAIL.n701 VTAIL.n682 3.49141
R1835 VTAIL.n722 VTAIL.n670 3.49141
R1836 VTAIL.n748 VTAIL.n747 3.49141
R1837 VTAIL.n43 VTAIL.n24 3.49141
R1838 VTAIL.n64 VTAIL.n12 3.49141
R1839 VTAIL.n90 VTAIL.n89 3.49141
R1840 VTAIL.n137 VTAIL.n118 3.49141
R1841 VTAIL.n158 VTAIL.n106 3.49141
R1842 VTAIL.n184 VTAIL.n183 3.49141
R1843 VTAIL.n231 VTAIL.n212 3.49141
R1844 VTAIL.n252 VTAIL.n200 3.49141
R1845 VTAIL.n278 VTAIL.n277 3.49141
R1846 VTAIL.n654 VTAIL.n653 3.49141
R1847 VTAIL.n629 VTAIL.n577 3.49141
R1848 VTAIL.n608 VTAIL.n589 3.49141
R1849 VTAIL.n560 VTAIL.n559 3.49141
R1850 VTAIL.n535 VTAIL.n483 3.49141
R1851 VTAIL.n514 VTAIL.n495 3.49141
R1852 VTAIL.n466 VTAIL.n465 3.49141
R1853 VTAIL.n441 VTAIL.n389 3.49141
R1854 VTAIL.n420 VTAIL.n401 3.49141
R1855 VTAIL.n372 VTAIL.n371 3.49141
R1856 VTAIL.n347 VTAIL.n295 3.49141
R1857 VTAIL.n326 VTAIL.n307 3.49141
R1858 VTAIL.n698 VTAIL.n697 2.71565
R1859 VTAIL.n726 VTAIL.n725 2.71565
R1860 VTAIL.n744 VTAIL.n660 2.71565
R1861 VTAIL.n40 VTAIL.n39 2.71565
R1862 VTAIL.n68 VTAIL.n67 2.71565
R1863 VTAIL.n86 VTAIL.n2 2.71565
R1864 VTAIL.n134 VTAIL.n133 2.71565
R1865 VTAIL.n162 VTAIL.n161 2.71565
R1866 VTAIL.n180 VTAIL.n96 2.71565
R1867 VTAIL.n228 VTAIL.n227 2.71565
R1868 VTAIL.n256 VTAIL.n255 2.71565
R1869 VTAIL.n274 VTAIL.n190 2.71565
R1870 VTAIL.n650 VTAIL.n566 2.71565
R1871 VTAIL.n633 VTAIL.n632 2.71565
R1872 VTAIL.n605 VTAIL.n604 2.71565
R1873 VTAIL.n556 VTAIL.n472 2.71565
R1874 VTAIL.n539 VTAIL.n538 2.71565
R1875 VTAIL.n511 VTAIL.n510 2.71565
R1876 VTAIL.n462 VTAIL.n378 2.71565
R1877 VTAIL.n445 VTAIL.n444 2.71565
R1878 VTAIL.n417 VTAIL.n416 2.71565
R1879 VTAIL.n368 VTAIL.n284 2.71565
R1880 VTAIL.n351 VTAIL.n350 2.71565
R1881 VTAIL.n323 VTAIL.n322 2.71565
R1882 VTAIL.n694 VTAIL.n684 1.93989
R1883 VTAIL.n730 VTAIL.n668 1.93989
R1884 VTAIL.n743 VTAIL.n662 1.93989
R1885 VTAIL.n36 VTAIL.n26 1.93989
R1886 VTAIL.n72 VTAIL.n10 1.93989
R1887 VTAIL.n85 VTAIL.n4 1.93989
R1888 VTAIL.n130 VTAIL.n120 1.93989
R1889 VTAIL.n166 VTAIL.n104 1.93989
R1890 VTAIL.n179 VTAIL.n98 1.93989
R1891 VTAIL.n224 VTAIL.n214 1.93989
R1892 VTAIL.n260 VTAIL.n198 1.93989
R1893 VTAIL.n273 VTAIL.n192 1.93989
R1894 VTAIL.n649 VTAIL.n568 1.93989
R1895 VTAIL.n636 VTAIL.n574 1.93989
R1896 VTAIL.n601 VTAIL.n591 1.93989
R1897 VTAIL.n555 VTAIL.n474 1.93989
R1898 VTAIL.n542 VTAIL.n480 1.93989
R1899 VTAIL.n507 VTAIL.n497 1.93989
R1900 VTAIL.n461 VTAIL.n380 1.93989
R1901 VTAIL.n448 VTAIL.n386 1.93989
R1902 VTAIL.n413 VTAIL.n403 1.93989
R1903 VTAIL.n367 VTAIL.n286 1.93989
R1904 VTAIL.n354 VTAIL.n292 1.93989
R1905 VTAIL.n319 VTAIL.n309 1.93989
R1906 VTAIL.n693 VTAIL.n686 1.16414
R1907 VTAIL.n731 VTAIL.n666 1.16414
R1908 VTAIL.n740 VTAIL.n739 1.16414
R1909 VTAIL.n35 VTAIL.n28 1.16414
R1910 VTAIL.n73 VTAIL.n8 1.16414
R1911 VTAIL.n82 VTAIL.n81 1.16414
R1912 VTAIL.n129 VTAIL.n122 1.16414
R1913 VTAIL.n167 VTAIL.n102 1.16414
R1914 VTAIL.n176 VTAIL.n175 1.16414
R1915 VTAIL.n223 VTAIL.n216 1.16414
R1916 VTAIL.n261 VTAIL.n196 1.16414
R1917 VTAIL.n270 VTAIL.n269 1.16414
R1918 VTAIL.n646 VTAIL.n645 1.16414
R1919 VTAIL.n637 VTAIL.n572 1.16414
R1920 VTAIL.n600 VTAIL.n593 1.16414
R1921 VTAIL.n552 VTAIL.n551 1.16414
R1922 VTAIL.n543 VTAIL.n478 1.16414
R1923 VTAIL.n506 VTAIL.n499 1.16414
R1924 VTAIL.n458 VTAIL.n457 1.16414
R1925 VTAIL.n449 VTAIL.n384 1.16414
R1926 VTAIL.n412 VTAIL.n405 1.16414
R1927 VTAIL.n364 VTAIL.n363 1.16414
R1928 VTAIL.n355 VTAIL.n290 1.16414
R1929 VTAIL.n318 VTAIL.n311 1.16414
R1930 VTAIL.n469 VTAIL.n375 1.10395
R1931 VTAIL.n657 VTAIL.n563 1.10395
R1932 VTAIL.n281 VTAIL.n187 1.10395
R1933 VTAIL VTAIL.n93 0.610414
R1934 VTAIL VTAIL.n751 0.494034
R1935 VTAIL.n563 VTAIL.n469 0.470328
R1936 VTAIL.n187 VTAIL.n93 0.470328
R1937 VTAIL.n690 VTAIL.n689 0.388379
R1938 VTAIL.n735 VTAIL.n734 0.388379
R1939 VTAIL.n736 VTAIL.n664 0.388379
R1940 VTAIL.n32 VTAIL.n31 0.388379
R1941 VTAIL.n77 VTAIL.n76 0.388379
R1942 VTAIL.n78 VTAIL.n6 0.388379
R1943 VTAIL.n126 VTAIL.n125 0.388379
R1944 VTAIL.n171 VTAIL.n170 0.388379
R1945 VTAIL.n172 VTAIL.n100 0.388379
R1946 VTAIL.n220 VTAIL.n219 0.388379
R1947 VTAIL.n265 VTAIL.n264 0.388379
R1948 VTAIL.n266 VTAIL.n194 0.388379
R1949 VTAIL.n642 VTAIL.n570 0.388379
R1950 VTAIL.n641 VTAIL.n640 0.388379
R1951 VTAIL.n597 VTAIL.n596 0.388379
R1952 VTAIL.n548 VTAIL.n476 0.388379
R1953 VTAIL.n547 VTAIL.n546 0.388379
R1954 VTAIL.n503 VTAIL.n502 0.388379
R1955 VTAIL.n454 VTAIL.n382 0.388379
R1956 VTAIL.n453 VTAIL.n452 0.388379
R1957 VTAIL.n409 VTAIL.n408 0.388379
R1958 VTAIL.n360 VTAIL.n288 0.388379
R1959 VTAIL.n359 VTAIL.n358 0.388379
R1960 VTAIL.n315 VTAIL.n314 0.388379
R1961 VTAIL.n692 VTAIL.n691 0.155672
R1962 VTAIL.n692 VTAIL.n683 0.155672
R1963 VTAIL.n699 VTAIL.n683 0.155672
R1964 VTAIL.n700 VTAIL.n699 0.155672
R1965 VTAIL.n700 VTAIL.n679 0.155672
R1966 VTAIL.n707 VTAIL.n679 0.155672
R1967 VTAIL.n708 VTAIL.n707 0.155672
R1968 VTAIL.n708 VTAIL.n675 0.155672
R1969 VTAIL.n715 VTAIL.n675 0.155672
R1970 VTAIL.n716 VTAIL.n715 0.155672
R1971 VTAIL.n716 VTAIL.n671 0.155672
R1972 VTAIL.n723 VTAIL.n671 0.155672
R1973 VTAIL.n724 VTAIL.n723 0.155672
R1974 VTAIL.n724 VTAIL.n667 0.155672
R1975 VTAIL.n732 VTAIL.n667 0.155672
R1976 VTAIL.n733 VTAIL.n732 0.155672
R1977 VTAIL.n733 VTAIL.n663 0.155672
R1978 VTAIL.n741 VTAIL.n663 0.155672
R1979 VTAIL.n742 VTAIL.n741 0.155672
R1980 VTAIL.n742 VTAIL.n659 0.155672
R1981 VTAIL.n749 VTAIL.n659 0.155672
R1982 VTAIL.n34 VTAIL.n33 0.155672
R1983 VTAIL.n34 VTAIL.n25 0.155672
R1984 VTAIL.n41 VTAIL.n25 0.155672
R1985 VTAIL.n42 VTAIL.n41 0.155672
R1986 VTAIL.n42 VTAIL.n21 0.155672
R1987 VTAIL.n49 VTAIL.n21 0.155672
R1988 VTAIL.n50 VTAIL.n49 0.155672
R1989 VTAIL.n50 VTAIL.n17 0.155672
R1990 VTAIL.n57 VTAIL.n17 0.155672
R1991 VTAIL.n58 VTAIL.n57 0.155672
R1992 VTAIL.n58 VTAIL.n13 0.155672
R1993 VTAIL.n65 VTAIL.n13 0.155672
R1994 VTAIL.n66 VTAIL.n65 0.155672
R1995 VTAIL.n66 VTAIL.n9 0.155672
R1996 VTAIL.n74 VTAIL.n9 0.155672
R1997 VTAIL.n75 VTAIL.n74 0.155672
R1998 VTAIL.n75 VTAIL.n5 0.155672
R1999 VTAIL.n83 VTAIL.n5 0.155672
R2000 VTAIL.n84 VTAIL.n83 0.155672
R2001 VTAIL.n84 VTAIL.n1 0.155672
R2002 VTAIL.n91 VTAIL.n1 0.155672
R2003 VTAIL.n128 VTAIL.n127 0.155672
R2004 VTAIL.n128 VTAIL.n119 0.155672
R2005 VTAIL.n135 VTAIL.n119 0.155672
R2006 VTAIL.n136 VTAIL.n135 0.155672
R2007 VTAIL.n136 VTAIL.n115 0.155672
R2008 VTAIL.n143 VTAIL.n115 0.155672
R2009 VTAIL.n144 VTAIL.n143 0.155672
R2010 VTAIL.n144 VTAIL.n111 0.155672
R2011 VTAIL.n151 VTAIL.n111 0.155672
R2012 VTAIL.n152 VTAIL.n151 0.155672
R2013 VTAIL.n152 VTAIL.n107 0.155672
R2014 VTAIL.n159 VTAIL.n107 0.155672
R2015 VTAIL.n160 VTAIL.n159 0.155672
R2016 VTAIL.n160 VTAIL.n103 0.155672
R2017 VTAIL.n168 VTAIL.n103 0.155672
R2018 VTAIL.n169 VTAIL.n168 0.155672
R2019 VTAIL.n169 VTAIL.n99 0.155672
R2020 VTAIL.n177 VTAIL.n99 0.155672
R2021 VTAIL.n178 VTAIL.n177 0.155672
R2022 VTAIL.n178 VTAIL.n95 0.155672
R2023 VTAIL.n185 VTAIL.n95 0.155672
R2024 VTAIL.n222 VTAIL.n221 0.155672
R2025 VTAIL.n222 VTAIL.n213 0.155672
R2026 VTAIL.n229 VTAIL.n213 0.155672
R2027 VTAIL.n230 VTAIL.n229 0.155672
R2028 VTAIL.n230 VTAIL.n209 0.155672
R2029 VTAIL.n237 VTAIL.n209 0.155672
R2030 VTAIL.n238 VTAIL.n237 0.155672
R2031 VTAIL.n238 VTAIL.n205 0.155672
R2032 VTAIL.n245 VTAIL.n205 0.155672
R2033 VTAIL.n246 VTAIL.n245 0.155672
R2034 VTAIL.n246 VTAIL.n201 0.155672
R2035 VTAIL.n253 VTAIL.n201 0.155672
R2036 VTAIL.n254 VTAIL.n253 0.155672
R2037 VTAIL.n254 VTAIL.n197 0.155672
R2038 VTAIL.n262 VTAIL.n197 0.155672
R2039 VTAIL.n263 VTAIL.n262 0.155672
R2040 VTAIL.n263 VTAIL.n193 0.155672
R2041 VTAIL.n271 VTAIL.n193 0.155672
R2042 VTAIL.n272 VTAIL.n271 0.155672
R2043 VTAIL.n272 VTAIL.n189 0.155672
R2044 VTAIL.n279 VTAIL.n189 0.155672
R2045 VTAIL.n655 VTAIL.n565 0.155672
R2046 VTAIL.n648 VTAIL.n565 0.155672
R2047 VTAIL.n648 VTAIL.n647 0.155672
R2048 VTAIL.n647 VTAIL.n569 0.155672
R2049 VTAIL.n639 VTAIL.n569 0.155672
R2050 VTAIL.n639 VTAIL.n638 0.155672
R2051 VTAIL.n638 VTAIL.n573 0.155672
R2052 VTAIL.n631 VTAIL.n573 0.155672
R2053 VTAIL.n631 VTAIL.n630 0.155672
R2054 VTAIL.n630 VTAIL.n578 0.155672
R2055 VTAIL.n623 VTAIL.n578 0.155672
R2056 VTAIL.n623 VTAIL.n622 0.155672
R2057 VTAIL.n622 VTAIL.n582 0.155672
R2058 VTAIL.n615 VTAIL.n582 0.155672
R2059 VTAIL.n615 VTAIL.n614 0.155672
R2060 VTAIL.n614 VTAIL.n586 0.155672
R2061 VTAIL.n607 VTAIL.n586 0.155672
R2062 VTAIL.n607 VTAIL.n606 0.155672
R2063 VTAIL.n606 VTAIL.n590 0.155672
R2064 VTAIL.n599 VTAIL.n590 0.155672
R2065 VTAIL.n599 VTAIL.n598 0.155672
R2066 VTAIL.n561 VTAIL.n471 0.155672
R2067 VTAIL.n554 VTAIL.n471 0.155672
R2068 VTAIL.n554 VTAIL.n553 0.155672
R2069 VTAIL.n553 VTAIL.n475 0.155672
R2070 VTAIL.n545 VTAIL.n475 0.155672
R2071 VTAIL.n545 VTAIL.n544 0.155672
R2072 VTAIL.n544 VTAIL.n479 0.155672
R2073 VTAIL.n537 VTAIL.n479 0.155672
R2074 VTAIL.n537 VTAIL.n536 0.155672
R2075 VTAIL.n536 VTAIL.n484 0.155672
R2076 VTAIL.n529 VTAIL.n484 0.155672
R2077 VTAIL.n529 VTAIL.n528 0.155672
R2078 VTAIL.n528 VTAIL.n488 0.155672
R2079 VTAIL.n521 VTAIL.n488 0.155672
R2080 VTAIL.n521 VTAIL.n520 0.155672
R2081 VTAIL.n520 VTAIL.n492 0.155672
R2082 VTAIL.n513 VTAIL.n492 0.155672
R2083 VTAIL.n513 VTAIL.n512 0.155672
R2084 VTAIL.n512 VTAIL.n496 0.155672
R2085 VTAIL.n505 VTAIL.n496 0.155672
R2086 VTAIL.n505 VTAIL.n504 0.155672
R2087 VTAIL.n467 VTAIL.n377 0.155672
R2088 VTAIL.n460 VTAIL.n377 0.155672
R2089 VTAIL.n460 VTAIL.n459 0.155672
R2090 VTAIL.n459 VTAIL.n381 0.155672
R2091 VTAIL.n451 VTAIL.n381 0.155672
R2092 VTAIL.n451 VTAIL.n450 0.155672
R2093 VTAIL.n450 VTAIL.n385 0.155672
R2094 VTAIL.n443 VTAIL.n385 0.155672
R2095 VTAIL.n443 VTAIL.n442 0.155672
R2096 VTAIL.n442 VTAIL.n390 0.155672
R2097 VTAIL.n435 VTAIL.n390 0.155672
R2098 VTAIL.n435 VTAIL.n434 0.155672
R2099 VTAIL.n434 VTAIL.n394 0.155672
R2100 VTAIL.n427 VTAIL.n394 0.155672
R2101 VTAIL.n427 VTAIL.n426 0.155672
R2102 VTAIL.n426 VTAIL.n398 0.155672
R2103 VTAIL.n419 VTAIL.n398 0.155672
R2104 VTAIL.n419 VTAIL.n418 0.155672
R2105 VTAIL.n418 VTAIL.n402 0.155672
R2106 VTAIL.n411 VTAIL.n402 0.155672
R2107 VTAIL.n411 VTAIL.n410 0.155672
R2108 VTAIL.n373 VTAIL.n283 0.155672
R2109 VTAIL.n366 VTAIL.n283 0.155672
R2110 VTAIL.n366 VTAIL.n365 0.155672
R2111 VTAIL.n365 VTAIL.n287 0.155672
R2112 VTAIL.n357 VTAIL.n287 0.155672
R2113 VTAIL.n357 VTAIL.n356 0.155672
R2114 VTAIL.n356 VTAIL.n291 0.155672
R2115 VTAIL.n349 VTAIL.n291 0.155672
R2116 VTAIL.n349 VTAIL.n348 0.155672
R2117 VTAIL.n348 VTAIL.n296 0.155672
R2118 VTAIL.n341 VTAIL.n296 0.155672
R2119 VTAIL.n341 VTAIL.n340 0.155672
R2120 VTAIL.n340 VTAIL.n300 0.155672
R2121 VTAIL.n333 VTAIL.n300 0.155672
R2122 VTAIL.n333 VTAIL.n332 0.155672
R2123 VTAIL.n332 VTAIL.n304 0.155672
R2124 VTAIL.n325 VTAIL.n304 0.155672
R2125 VTAIL.n325 VTAIL.n324 0.155672
R2126 VTAIL.n324 VTAIL.n308 0.155672
R2127 VTAIL.n317 VTAIL.n308 0.155672
R2128 VTAIL.n317 VTAIL.n316 0.155672
R2129 VDD1 VDD1.n1 108.993
R2130 VDD1 VDD1.n0 67.1228
R2131 VDD1.n0 VDD1.t0 1.94924
R2132 VDD1.n0 VDD1.t2 1.94924
R2133 VDD1.n1 VDD1.t1 1.94924
R2134 VDD1.n1 VDD1.t3 1.94924
R2135 VN.n0 VN.t2 483.103
R2136 VN.n1 VN.t1 483.103
R2137 VN.n1 VN.t3 483.017
R2138 VN.n0 VN.t0 483.017
R2139 VN VN.n1 76.3039
R2140 VN VN.n0 31.2622
R2141 VDD2.n2 VDD2.n0 108.469
R2142 VDD2.n2 VDD2.n1 67.0646
R2143 VDD2.n1 VDD2.t0 1.94924
R2144 VDD2.n1 VDD2.t2 1.94924
R2145 VDD2.n0 VDD2.t1 1.94924
R2146 VDD2.n0 VDD2.t3 1.94924
R2147 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 4.35591f
C1 VTAIL w_n1738_n4304# 5.24016f
C2 VDD2 VDD1 0.626737f
C3 VN VDD1 0.147952f
C4 VDD2 VTAIL 7.95423f
C5 B VP 1.20828f
C6 w_n1738_n4304# B 8.52755f
C7 VTAIL VN 4.3418f
C8 VTAIL VDD1 7.91108f
C9 w_n1738_n4304# VP 2.94694f
C10 VDD2 B 1.12189f
C11 VN B 0.852115f
C12 VDD2 VP 0.289756f
C13 VDD2 w_n1738_n4304# 1.26682f
C14 B VDD1 1.09659f
C15 VN VP 5.86829f
C16 VN w_n1738_n4304# 2.72769f
C17 VDD1 VP 5.0153f
C18 w_n1738_n4304# VDD1 1.24716f
C19 VTAIL B 5.32227f
C20 VDD2 VN 4.87382f
C21 VDD2 VSUBS 0.822232f
C22 VDD1 VSUBS 5.633218f
C23 VTAIL VSUBS 1.139409f
C24 VN VSUBS 5.86609f
C25 VP VSUBS 1.616683f
C26 B VSUBS 3.240074f
C27 w_n1738_n4304# VSUBS 91.578705f
C28 VDD2.t1 VSUBS 0.362739f
C29 VDD2.t3 VSUBS 0.362739f
C30 VDD2.n0 VSUBS 3.83018f
C31 VDD2.t0 VSUBS 0.362739f
C32 VDD2.t2 VSUBS 0.362739f
C33 VDD2.n1 VSUBS 2.9724f
C34 VDD2.n2 VSUBS 4.54269f
C35 VN.t2 VSUBS 2.33279f
C36 VN.t0 VSUBS 2.33261f
C37 VN.n0 VSUBS 1.68128f
C38 VN.t1 VSUBS 2.33279f
C39 VN.t3 VSUBS 2.33261f
C40 VN.n1 VSUBS 3.17642f
C41 VDD1.t0 VSUBS 0.359903f
C42 VDD1.t2 VSUBS 0.359903f
C43 VDD1.n0 VSUBS 2.94974f
C44 VDD1.t1 VSUBS 0.359903f
C45 VDD1.t3 VSUBS 0.359903f
C46 VDD1.n1 VSUBS 3.8279f
C47 VTAIL.n0 VSUBS 0.022309f
C48 VTAIL.n1 VSUBS 0.022092f
C49 VTAIL.n2 VSUBS 0.011871f
C50 VTAIL.n3 VSUBS 0.028059f
C51 VTAIL.n4 VSUBS 0.01257f
C52 VTAIL.n5 VSUBS 0.022092f
C53 VTAIL.n6 VSUBS 0.011871f
C54 VTAIL.n7 VSUBS 0.028059f
C55 VTAIL.n8 VSUBS 0.01257f
C56 VTAIL.n9 VSUBS 0.022092f
C57 VTAIL.n10 VSUBS 0.011871f
C58 VTAIL.n11 VSUBS 0.028059f
C59 VTAIL.n12 VSUBS 0.01257f
C60 VTAIL.n13 VSUBS 0.022092f
C61 VTAIL.n14 VSUBS 0.011871f
C62 VTAIL.n15 VSUBS 0.028059f
C63 VTAIL.n16 VSUBS 0.01257f
C64 VTAIL.n17 VSUBS 0.022092f
C65 VTAIL.n18 VSUBS 0.011871f
C66 VTAIL.n19 VSUBS 0.028059f
C67 VTAIL.n20 VSUBS 0.01257f
C68 VTAIL.n21 VSUBS 0.022092f
C69 VTAIL.n22 VSUBS 0.011871f
C70 VTAIL.n23 VSUBS 0.028059f
C71 VTAIL.n24 VSUBS 0.01257f
C72 VTAIL.n25 VSUBS 0.022092f
C73 VTAIL.n26 VSUBS 0.011871f
C74 VTAIL.n27 VSUBS 0.028059f
C75 VTAIL.n28 VSUBS 0.01257f
C76 VTAIL.n29 VSUBS 0.166676f
C77 VTAIL.t1 VSUBS 0.060162f
C78 VTAIL.n30 VSUBS 0.021045f
C79 VTAIL.n31 VSUBS 0.01785f
C80 VTAIL.n32 VSUBS 0.011871f
C81 VTAIL.n33 VSUBS 1.5791f
C82 VTAIL.n34 VSUBS 0.022092f
C83 VTAIL.n35 VSUBS 0.011871f
C84 VTAIL.n36 VSUBS 0.01257f
C85 VTAIL.n37 VSUBS 0.028059f
C86 VTAIL.n38 VSUBS 0.028059f
C87 VTAIL.n39 VSUBS 0.01257f
C88 VTAIL.n40 VSUBS 0.011871f
C89 VTAIL.n41 VSUBS 0.022092f
C90 VTAIL.n42 VSUBS 0.022092f
C91 VTAIL.n43 VSUBS 0.011871f
C92 VTAIL.n44 VSUBS 0.01257f
C93 VTAIL.n45 VSUBS 0.028059f
C94 VTAIL.n46 VSUBS 0.028059f
C95 VTAIL.n47 VSUBS 0.01257f
C96 VTAIL.n48 VSUBS 0.011871f
C97 VTAIL.n49 VSUBS 0.022092f
C98 VTAIL.n50 VSUBS 0.022092f
C99 VTAIL.n51 VSUBS 0.011871f
C100 VTAIL.n52 VSUBS 0.01257f
C101 VTAIL.n53 VSUBS 0.028059f
C102 VTAIL.n54 VSUBS 0.028059f
C103 VTAIL.n55 VSUBS 0.01257f
C104 VTAIL.n56 VSUBS 0.011871f
C105 VTAIL.n57 VSUBS 0.022092f
C106 VTAIL.n58 VSUBS 0.022092f
C107 VTAIL.n59 VSUBS 0.011871f
C108 VTAIL.n60 VSUBS 0.01257f
C109 VTAIL.n61 VSUBS 0.028059f
C110 VTAIL.n62 VSUBS 0.028059f
C111 VTAIL.n63 VSUBS 0.01257f
C112 VTAIL.n64 VSUBS 0.011871f
C113 VTAIL.n65 VSUBS 0.022092f
C114 VTAIL.n66 VSUBS 0.022092f
C115 VTAIL.n67 VSUBS 0.011871f
C116 VTAIL.n68 VSUBS 0.01257f
C117 VTAIL.n69 VSUBS 0.028059f
C118 VTAIL.n70 VSUBS 0.028059f
C119 VTAIL.n71 VSUBS 0.028059f
C120 VTAIL.n72 VSUBS 0.01257f
C121 VTAIL.n73 VSUBS 0.011871f
C122 VTAIL.n74 VSUBS 0.022092f
C123 VTAIL.n75 VSUBS 0.022092f
C124 VTAIL.n76 VSUBS 0.011871f
C125 VTAIL.n77 VSUBS 0.01222f
C126 VTAIL.n78 VSUBS 0.01222f
C127 VTAIL.n79 VSUBS 0.028059f
C128 VTAIL.n80 VSUBS 0.028059f
C129 VTAIL.n81 VSUBS 0.01257f
C130 VTAIL.n82 VSUBS 0.011871f
C131 VTAIL.n83 VSUBS 0.022092f
C132 VTAIL.n84 VSUBS 0.022092f
C133 VTAIL.n85 VSUBS 0.011871f
C134 VTAIL.n86 VSUBS 0.01257f
C135 VTAIL.n87 VSUBS 0.028059f
C136 VTAIL.n88 VSUBS 0.061234f
C137 VTAIL.n89 VSUBS 0.01257f
C138 VTAIL.n90 VSUBS 0.011871f
C139 VTAIL.n91 VSUBS 0.047443f
C140 VTAIL.n92 VSUBS 0.030382f
C141 VTAIL.n93 VSUBS 0.09369f
C142 VTAIL.n94 VSUBS 0.022309f
C143 VTAIL.n95 VSUBS 0.022092f
C144 VTAIL.n96 VSUBS 0.011871f
C145 VTAIL.n97 VSUBS 0.028059f
C146 VTAIL.n98 VSUBS 0.01257f
C147 VTAIL.n99 VSUBS 0.022092f
C148 VTAIL.n100 VSUBS 0.011871f
C149 VTAIL.n101 VSUBS 0.028059f
C150 VTAIL.n102 VSUBS 0.01257f
C151 VTAIL.n103 VSUBS 0.022092f
C152 VTAIL.n104 VSUBS 0.011871f
C153 VTAIL.n105 VSUBS 0.028059f
C154 VTAIL.n106 VSUBS 0.01257f
C155 VTAIL.n107 VSUBS 0.022092f
C156 VTAIL.n108 VSUBS 0.011871f
C157 VTAIL.n109 VSUBS 0.028059f
C158 VTAIL.n110 VSUBS 0.01257f
C159 VTAIL.n111 VSUBS 0.022092f
C160 VTAIL.n112 VSUBS 0.011871f
C161 VTAIL.n113 VSUBS 0.028059f
C162 VTAIL.n114 VSUBS 0.01257f
C163 VTAIL.n115 VSUBS 0.022092f
C164 VTAIL.n116 VSUBS 0.011871f
C165 VTAIL.n117 VSUBS 0.028059f
C166 VTAIL.n118 VSUBS 0.01257f
C167 VTAIL.n119 VSUBS 0.022092f
C168 VTAIL.n120 VSUBS 0.011871f
C169 VTAIL.n121 VSUBS 0.028059f
C170 VTAIL.n122 VSUBS 0.01257f
C171 VTAIL.n123 VSUBS 0.166676f
C172 VTAIL.t7 VSUBS 0.060162f
C173 VTAIL.n124 VSUBS 0.021045f
C174 VTAIL.n125 VSUBS 0.01785f
C175 VTAIL.n126 VSUBS 0.011871f
C176 VTAIL.n127 VSUBS 1.5791f
C177 VTAIL.n128 VSUBS 0.022092f
C178 VTAIL.n129 VSUBS 0.011871f
C179 VTAIL.n130 VSUBS 0.01257f
C180 VTAIL.n131 VSUBS 0.028059f
C181 VTAIL.n132 VSUBS 0.028059f
C182 VTAIL.n133 VSUBS 0.01257f
C183 VTAIL.n134 VSUBS 0.011871f
C184 VTAIL.n135 VSUBS 0.022092f
C185 VTAIL.n136 VSUBS 0.022092f
C186 VTAIL.n137 VSUBS 0.011871f
C187 VTAIL.n138 VSUBS 0.01257f
C188 VTAIL.n139 VSUBS 0.028059f
C189 VTAIL.n140 VSUBS 0.028059f
C190 VTAIL.n141 VSUBS 0.01257f
C191 VTAIL.n142 VSUBS 0.011871f
C192 VTAIL.n143 VSUBS 0.022092f
C193 VTAIL.n144 VSUBS 0.022092f
C194 VTAIL.n145 VSUBS 0.011871f
C195 VTAIL.n146 VSUBS 0.01257f
C196 VTAIL.n147 VSUBS 0.028059f
C197 VTAIL.n148 VSUBS 0.028059f
C198 VTAIL.n149 VSUBS 0.01257f
C199 VTAIL.n150 VSUBS 0.011871f
C200 VTAIL.n151 VSUBS 0.022092f
C201 VTAIL.n152 VSUBS 0.022092f
C202 VTAIL.n153 VSUBS 0.011871f
C203 VTAIL.n154 VSUBS 0.01257f
C204 VTAIL.n155 VSUBS 0.028059f
C205 VTAIL.n156 VSUBS 0.028059f
C206 VTAIL.n157 VSUBS 0.01257f
C207 VTAIL.n158 VSUBS 0.011871f
C208 VTAIL.n159 VSUBS 0.022092f
C209 VTAIL.n160 VSUBS 0.022092f
C210 VTAIL.n161 VSUBS 0.011871f
C211 VTAIL.n162 VSUBS 0.01257f
C212 VTAIL.n163 VSUBS 0.028059f
C213 VTAIL.n164 VSUBS 0.028059f
C214 VTAIL.n165 VSUBS 0.028059f
C215 VTAIL.n166 VSUBS 0.01257f
C216 VTAIL.n167 VSUBS 0.011871f
C217 VTAIL.n168 VSUBS 0.022092f
C218 VTAIL.n169 VSUBS 0.022092f
C219 VTAIL.n170 VSUBS 0.011871f
C220 VTAIL.n171 VSUBS 0.01222f
C221 VTAIL.n172 VSUBS 0.01222f
C222 VTAIL.n173 VSUBS 0.028059f
C223 VTAIL.n174 VSUBS 0.028059f
C224 VTAIL.n175 VSUBS 0.01257f
C225 VTAIL.n176 VSUBS 0.011871f
C226 VTAIL.n177 VSUBS 0.022092f
C227 VTAIL.n178 VSUBS 0.022092f
C228 VTAIL.n179 VSUBS 0.011871f
C229 VTAIL.n180 VSUBS 0.01257f
C230 VTAIL.n181 VSUBS 0.028059f
C231 VTAIL.n182 VSUBS 0.061234f
C232 VTAIL.n183 VSUBS 0.01257f
C233 VTAIL.n184 VSUBS 0.011871f
C234 VTAIL.n185 VSUBS 0.047443f
C235 VTAIL.n186 VSUBS 0.030382f
C236 VTAIL.n187 VSUBS 0.128822f
C237 VTAIL.n188 VSUBS 0.022309f
C238 VTAIL.n189 VSUBS 0.022092f
C239 VTAIL.n190 VSUBS 0.011871f
C240 VTAIL.n191 VSUBS 0.028059f
C241 VTAIL.n192 VSUBS 0.01257f
C242 VTAIL.n193 VSUBS 0.022092f
C243 VTAIL.n194 VSUBS 0.011871f
C244 VTAIL.n195 VSUBS 0.028059f
C245 VTAIL.n196 VSUBS 0.01257f
C246 VTAIL.n197 VSUBS 0.022092f
C247 VTAIL.n198 VSUBS 0.011871f
C248 VTAIL.n199 VSUBS 0.028059f
C249 VTAIL.n200 VSUBS 0.01257f
C250 VTAIL.n201 VSUBS 0.022092f
C251 VTAIL.n202 VSUBS 0.011871f
C252 VTAIL.n203 VSUBS 0.028059f
C253 VTAIL.n204 VSUBS 0.01257f
C254 VTAIL.n205 VSUBS 0.022092f
C255 VTAIL.n206 VSUBS 0.011871f
C256 VTAIL.n207 VSUBS 0.028059f
C257 VTAIL.n208 VSUBS 0.01257f
C258 VTAIL.n209 VSUBS 0.022092f
C259 VTAIL.n210 VSUBS 0.011871f
C260 VTAIL.n211 VSUBS 0.028059f
C261 VTAIL.n212 VSUBS 0.01257f
C262 VTAIL.n213 VSUBS 0.022092f
C263 VTAIL.n214 VSUBS 0.011871f
C264 VTAIL.n215 VSUBS 0.028059f
C265 VTAIL.n216 VSUBS 0.01257f
C266 VTAIL.n217 VSUBS 0.166676f
C267 VTAIL.t4 VSUBS 0.060162f
C268 VTAIL.n218 VSUBS 0.021045f
C269 VTAIL.n219 VSUBS 0.01785f
C270 VTAIL.n220 VSUBS 0.011871f
C271 VTAIL.n221 VSUBS 1.5791f
C272 VTAIL.n222 VSUBS 0.022092f
C273 VTAIL.n223 VSUBS 0.011871f
C274 VTAIL.n224 VSUBS 0.01257f
C275 VTAIL.n225 VSUBS 0.028059f
C276 VTAIL.n226 VSUBS 0.028059f
C277 VTAIL.n227 VSUBS 0.01257f
C278 VTAIL.n228 VSUBS 0.011871f
C279 VTAIL.n229 VSUBS 0.022092f
C280 VTAIL.n230 VSUBS 0.022092f
C281 VTAIL.n231 VSUBS 0.011871f
C282 VTAIL.n232 VSUBS 0.01257f
C283 VTAIL.n233 VSUBS 0.028059f
C284 VTAIL.n234 VSUBS 0.028059f
C285 VTAIL.n235 VSUBS 0.01257f
C286 VTAIL.n236 VSUBS 0.011871f
C287 VTAIL.n237 VSUBS 0.022092f
C288 VTAIL.n238 VSUBS 0.022092f
C289 VTAIL.n239 VSUBS 0.011871f
C290 VTAIL.n240 VSUBS 0.01257f
C291 VTAIL.n241 VSUBS 0.028059f
C292 VTAIL.n242 VSUBS 0.028059f
C293 VTAIL.n243 VSUBS 0.01257f
C294 VTAIL.n244 VSUBS 0.011871f
C295 VTAIL.n245 VSUBS 0.022092f
C296 VTAIL.n246 VSUBS 0.022092f
C297 VTAIL.n247 VSUBS 0.011871f
C298 VTAIL.n248 VSUBS 0.01257f
C299 VTAIL.n249 VSUBS 0.028059f
C300 VTAIL.n250 VSUBS 0.028059f
C301 VTAIL.n251 VSUBS 0.01257f
C302 VTAIL.n252 VSUBS 0.011871f
C303 VTAIL.n253 VSUBS 0.022092f
C304 VTAIL.n254 VSUBS 0.022092f
C305 VTAIL.n255 VSUBS 0.011871f
C306 VTAIL.n256 VSUBS 0.01257f
C307 VTAIL.n257 VSUBS 0.028059f
C308 VTAIL.n258 VSUBS 0.028059f
C309 VTAIL.n259 VSUBS 0.028059f
C310 VTAIL.n260 VSUBS 0.01257f
C311 VTAIL.n261 VSUBS 0.011871f
C312 VTAIL.n262 VSUBS 0.022092f
C313 VTAIL.n263 VSUBS 0.022092f
C314 VTAIL.n264 VSUBS 0.011871f
C315 VTAIL.n265 VSUBS 0.01222f
C316 VTAIL.n266 VSUBS 0.01222f
C317 VTAIL.n267 VSUBS 0.028059f
C318 VTAIL.n268 VSUBS 0.028059f
C319 VTAIL.n269 VSUBS 0.01257f
C320 VTAIL.n270 VSUBS 0.011871f
C321 VTAIL.n271 VSUBS 0.022092f
C322 VTAIL.n272 VSUBS 0.022092f
C323 VTAIL.n273 VSUBS 0.011871f
C324 VTAIL.n274 VSUBS 0.01257f
C325 VTAIL.n275 VSUBS 0.028059f
C326 VTAIL.n276 VSUBS 0.061234f
C327 VTAIL.n277 VSUBS 0.01257f
C328 VTAIL.n278 VSUBS 0.011871f
C329 VTAIL.n279 VSUBS 0.047443f
C330 VTAIL.n280 VSUBS 0.030382f
C331 VTAIL.n281 VSUBS 1.49761f
C332 VTAIL.n282 VSUBS 0.022309f
C333 VTAIL.n283 VSUBS 0.022092f
C334 VTAIL.n284 VSUBS 0.011871f
C335 VTAIL.n285 VSUBS 0.028059f
C336 VTAIL.n286 VSUBS 0.01257f
C337 VTAIL.n287 VSUBS 0.022092f
C338 VTAIL.n288 VSUBS 0.011871f
C339 VTAIL.n289 VSUBS 0.028059f
C340 VTAIL.n290 VSUBS 0.01257f
C341 VTAIL.n291 VSUBS 0.022092f
C342 VTAIL.n292 VSUBS 0.011871f
C343 VTAIL.n293 VSUBS 0.028059f
C344 VTAIL.n294 VSUBS 0.028059f
C345 VTAIL.n295 VSUBS 0.01257f
C346 VTAIL.n296 VSUBS 0.022092f
C347 VTAIL.n297 VSUBS 0.011871f
C348 VTAIL.n298 VSUBS 0.028059f
C349 VTAIL.n299 VSUBS 0.01257f
C350 VTAIL.n300 VSUBS 0.022092f
C351 VTAIL.n301 VSUBS 0.011871f
C352 VTAIL.n302 VSUBS 0.028059f
C353 VTAIL.n303 VSUBS 0.01257f
C354 VTAIL.n304 VSUBS 0.022092f
C355 VTAIL.n305 VSUBS 0.011871f
C356 VTAIL.n306 VSUBS 0.028059f
C357 VTAIL.n307 VSUBS 0.01257f
C358 VTAIL.n308 VSUBS 0.022092f
C359 VTAIL.n309 VSUBS 0.011871f
C360 VTAIL.n310 VSUBS 0.028059f
C361 VTAIL.n311 VSUBS 0.01257f
C362 VTAIL.n312 VSUBS 0.166676f
C363 VTAIL.t3 VSUBS 0.060162f
C364 VTAIL.n313 VSUBS 0.021045f
C365 VTAIL.n314 VSUBS 0.01785f
C366 VTAIL.n315 VSUBS 0.011871f
C367 VTAIL.n316 VSUBS 1.5791f
C368 VTAIL.n317 VSUBS 0.022092f
C369 VTAIL.n318 VSUBS 0.011871f
C370 VTAIL.n319 VSUBS 0.01257f
C371 VTAIL.n320 VSUBS 0.028059f
C372 VTAIL.n321 VSUBS 0.028059f
C373 VTAIL.n322 VSUBS 0.01257f
C374 VTAIL.n323 VSUBS 0.011871f
C375 VTAIL.n324 VSUBS 0.022092f
C376 VTAIL.n325 VSUBS 0.022092f
C377 VTAIL.n326 VSUBS 0.011871f
C378 VTAIL.n327 VSUBS 0.01257f
C379 VTAIL.n328 VSUBS 0.028059f
C380 VTAIL.n329 VSUBS 0.028059f
C381 VTAIL.n330 VSUBS 0.01257f
C382 VTAIL.n331 VSUBS 0.011871f
C383 VTAIL.n332 VSUBS 0.022092f
C384 VTAIL.n333 VSUBS 0.022092f
C385 VTAIL.n334 VSUBS 0.011871f
C386 VTAIL.n335 VSUBS 0.01257f
C387 VTAIL.n336 VSUBS 0.028059f
C388 VTAIL.n337 VSUBS 0.028059f
C389 VTAIL.n338 VSUBS 0.01257f
C390 VTAIL.n339 VSUBS 0.011871f
C391 VTAIL.n340 VSUBS 0.022092f
C392 VTAIL.n341 VSUBS 0.022092f
C393 VTAIL.n342 VSUBS 0.011871f
C394 VTAIL.n343 VSUBS 0.01257f
C395 VTAIL.n344 VSUBS 0.028059f
C396 VTAIL.n345 VSUBS 0.028059f
C397 VTAIL.n346 VSUBS 0.01257f
C398 VTAIL.n347 VSUBS 0.011871f
C399 VTAIL.n348 VSUBS 0.022092f
C400 VTAIL.n349 VSUBS 0.022092f
C401 VTAIL.n350 VSUBS 0.011871f
C402 VTAIL.n351 VSUBS 0.01257f
C403 VTAIL.n352 VSUBS 0.028059f
C404 VTAIL.n353 VSUBS 0.028059f
C405 VTAIL.n354 VSUBS 0.01257f
C406 VTAIL.n355 VSUBS 0.011871f
C407 VTAIL.n356 VSUBS 0.022092f
C408 VTAIL.n357 VSUBS 0.022092f
C409 VTAIL.n358 VSUBS 0.011871f
C410 VTAIL.n359 VSUBS 0.01222f
C411 VTAIL.n360 VSUBS 0.01222f
C412 VTAIL.n361 VSUBS 0.028059f
C413 VTAIL.n362 VSUBS 0.028059f
C414 VTAIL.n363 VSUBS 0.01257f
C415 VTAIL.n364 VSUBS 0.011871f
C416 VTAIL.n365 VSUBS 0.022092f
C417 VTAIL.n366 VSUBS 0.022092f
C418 VTAIL.n367 VSUBS 0.011871f
C419 VTAIL.n368 VSUBS 0.01257f
C420 VTAIL.n369 VSUBS 0.028059f
C421 VTAIL.n370 VSUBS 0.061234f
C422 VTAIL.n371 VSUBS 0.01257f
C423 VTAIL.n372 VSUBS 0.011871f
C424 VTAIL.n373 VSUBS 0.047443f
C425 VTAIL.n374 VSUBS 0.030382f
C426 VTAIL.n375 VSUBS 1.49761f
C427 VTAIL.n376 VSUBS 0.022309f
C428 VTAIL.n377 VSUBS 0.022092f
C429 VTAIL.n378 VSUBS 0.011871f
C430 VTAIL.n379 VSUBS 0.028059f
C431 VTAIL.n380 VSUBS 0.01257f
C432 VTAIL.n381 VSUBS 0.022092f
C433 VTAIL.n382 VSUBS 0.011871f
C434 VTAIL.n383 VSUBS 0.028059f
C435 VTAIL.n384 VSUBS 0.01257f
C436 VTAIL.n385 VSUBS 0.022092f
C437 VTAIL.n386 VSUBS 0.011871f
C438 VTAIL.n387 VSUBS 0.028059f
C439 VTAIL.n388 VSUBS 0.028059f
C440 VTAIL.n389 VSUBS 0.01257f
C441 VTAIL.n390 VSUBS 0.022092f
C442 VTAIL.n391 VSUBS 0.011871f
C443 VTAIL.n392 VSUBS 0.028059f
C444 VTAIL.n393 VSUBS 0.01257f
C445 VTAIL.n394 VSUBS 0.022092f
C446 VTAIL.n395 VSUBS 0.011871f
C447 VTAIL.n396 VSUBS 0.028059f
C448 VTAIL.n397 VSUBS 0.01257f
C449 VTAIL.n398 VSUBS 0.022092f
C450 VTAIL.n399 VSUBS 0.011871f
C451 VTAIL.n400 VSUBS 0.028059f
C452 VTAIL.n401 VSUBS 0.01257f
C453 VTAIL.n402 VSUBS 0.022092f
C454 VTAIL.n403 VSUBS 0.011871f
C455 VTAIL.n404 VSUBS 0.028059f
C456 VTAIL.n405 VSUBS 0.01257f
C457 VTAIL.n406 VSUBS 0.166676f
C458 VTAIL.t2 VSUBS 0.060162f
C459 VTAIL.n407 VSUBS 0.021045f
C460 VTAIL.n408 VSUBS 0.01785f
C461 VTAIL.n409 VSUBS 0.011871f
C462 VTAIL.n410 VSUBS 1.5791f
C463 VTAIL.n411 VSUBS 0.022092f
C464 VTAIL.n412 VSUBS 0.011871f
C465 VTAIL.n413 VSUBS 0.01257f
C466 VTAIL.n414 VSUBS 0.028059f
C467 VTAIL.n415 VSUBS 0.028059f
C468 VTAIL.n416 VSUBS 0.01257f
C469 VTAIL.n417 VSUBS 0.011871f
C470 VTAIL.n418 VSUBS 0.022092f
C471 VTAIL.n419 VSUBS 0.022092f
C472 VTAIL.n420 VSUBS 0.011871f
C473 VTAIL.n421 VSUBS 0.01257f
C474 VTAIL.n422 VSUBS 0.028059f
C475 VTAIL.n423 VSUBS 0.028059f
C476 VTAIL.n424 VSUBS 0.01257f
C477 VTAIL.n425 VSUBS 0.011871f
C478 VTAIL.n426 VSUBS 0.022092f
C479 VTAIL.n427 VSUBS 0.022092f
C480 VTAIL.n428 VSUBS 0.011871f
C481 VTAIL.n429 VSUBS 0.01257f
C482 VTAIL.n430 VSUBS 0.028059f
C483 VTAIL.n431 VSUBS 0.028059f
C484 VTAIL.n432 VSUBS 0.01257f
C485 VTAIL.n433 VSUBS 0.011871f
C486 VTAIL.n434 VSUBS 0.022092f
C487 VTAIL.n435 VSUBS 0.022092f
C488 VTAIL.n436 VSUBS 0.011871f
C489 VTAIL.n437 VSUBS 0.01257f
C490 VTAIL.n438 VSUBS 0.028059f
C491 VTAIL.n439 VSUBS 0.028059f
C492 VTAIL.n440 VSUBS 0.01257f
C493 VTAIL.n441 VSUBS 0.011871f
C494 VTAIL.n442 VSUBS 0.022092f
C495 VTAIL.n443 VSUBS 0.022092f
C496 VTAIL.n444 VSUBS 0.011871f
C497 VTAIL.n445 VSUBS 0.01257f
C498 VTAIL.n446 VSUBS 0.028059f
C499 VTAIL.n447 VSUBS 0.028059f
C500 VTAIL.n448 VSUBS 0.01257f
C501 VTAIL.n449 VSUBS 0.011871f
C502 VTAIL.n450 VSUBS 0.022092f
C503 VTAIL.n451 VSUBS 0.022092f
C504 VTAIL.n452 VSUBS 0.011871f
C505 VTAIL.n453 VSUBS 0.01222f
C506 VTAIL.n454 VSUBS 0.01222f
C507 VTAIL.n455 VSUBS 0.028059f
C508 VTAIL.n456 VSUBS 0.028059f
C509 VTAIL.n457 VSUBS 0.01257f
C510 VTAIL.n458 VSUBS 0.011871f
C511 VTAIL.n459 VSUBS 0.022092f
C512 VTAIL.n460 VSUBS 0.022092f
C513 VTAIL.n461 VSUBS 0.011871f
C514 VTAIL.n462 VSUBS 0.01257f
C515 VTAIL.n463 VSUBS 0.028059f
C516 VTAIL.n464 VSUBS 0.061234f
C517 VTAIL.n465 VSUBS 0.01257f
C518 VTAIL.n466 VSUBS 0.011871f
C519 VTAIL.n467 VSUBS 0.047443f
C520 VTAIL.n468 VSUBS 0.030382f
C521 VTAIL.n469 VSUBS 0.128822f
C522 VTAIL.n470 VSUBS 0.022309f
C523 VTAIL.n471 VSUBS 0.022092f
C524 VTAIL.n472 VSUBS 0.011871f
C525 VTAIL.n473 VSUBS 0.028059f
C526 VTAIL.n474 VSUBS 0.01257f
C527 VTAIL.n475 VSUBS 0.022092f
C528 VTAIL.n476 VSUBS 0.011871f
C529 VTAIL.n477 VSUBS 0.028059f
C530 VTAIL.n478 VSUBS 0.01257f
C531 VTAIL.n479 VSUBS 0.022092f
C532 VTAIL.n480 VSUBS 0.011871f
C533 VTAIL.n481 VSUBS 0.028059f
C534 VTAIL.n482 VSUBS 0.028059f
C535 VTAIL.n483 VSUBS 0.01257f
C536 VTAIL.n484 VSUBS 0.022092f
C537 VTAIL.n485 VSUBS 0.011871f
C538 VTAIL.n486 VSUBS 0.028059f
C539 VTAIL.n487 VSUBS 0.01257f
C540 VTAIL.n488 VSUBS 0.022092f
C541 VTAIL.n489 VSUBS 0.011871f
C542 VTAIL.n490 VSUBS 0.028059f
C543 VTAIL.n491 VSUBS 0.01257f
C544 VTAIL.n492 VSUBS 0.022092f
C545 VTAIL.n493 VSUBS 0.011871f
C546 VTAIL.n494 VSUBS 0.028059f
C547 VTAIL.n495 VSUBS 0.01257f
C548 VTAIL.n496 VSUBS 0.022092f
C549 VTAIL.n497 VSUBS 0.011871f
C550 VTAIL.n498 VSUBS 0.028059f
C551 VTAIL.n499 VSUBS 0.01257f
C552 VTAIL.n500 VSUBS 0.166676f
C553 VTAIL.t6 VSUBS 0.060162f
C554 VTAIL.n501 VSUBS 0.021045f
C555 VTAIL.n502 VSUBS 0.01785f
C556 VTAIL.n503 VSUBS 0.011871f
C557 VTAIL.n504 VSUBS 1.5791f
C558 VTAIL.n505 VSUBS 0.022092f
C559 VTAIL.n506 VSUBS 0.011871f
C560 VTAIL.n507 VSUBS 0.01257f
C561 VTAIL.n508 VSUBS 0.028059f
C562 VTAIL.n509 VSUBS 0.028059f
C563 VTAIL.n510 VSUBS 0.01257f
C564 VTAIL.n511 VSUBS 0.011871f
C565 VTAIL.n512 VSUBS 0.022092f
C566 VTAIL.n513 VSUBS 0.022092f
C567 VTAIL.n514 VSUBS 0.011871f
C568 VTAIL.n515 VSUBS 0.01257f
C569 VTAIL.n516 VSUBS 0.028059f
C570 VTAIL.n517 VSUBS 0.028059f
C571 VTAIL.n518 VSUBS 0.01257f
C572 VTAIL.n519 VSUBS 0.011871f
C573 VTAIL.n520 VSUBS 0.022092f
C574 VTAIL.n521 VSUBS 0.022092f
C575 VTAIL.n522 VSUBS 0.011871f
C576 VTAIL.n523 VSUBS 0.01257f
C577 VTAIL.n524 VSUBS 0.028059f
C578 VTAIL.n525 VSUBS 0.028059f
C579 VTAIL.n526 VSUBS 0.01257f
C580 VTAIL.n527 VSUBS 0.011871f
C581 VTAIL.n528 VSUBS 0.022092f
C582 VTAIL.n529 VSUBS 0.022092f
C583 VTAIL.n530 VSUBS 0.011871f
C584 VTAIL.n531 VSUBS 0.01257f
C585 VTAIL.n532 VSUBS 0.028059f
C586 VTAIL.n533 VSUBS 0.028059f
C587 VTAIL.n534 VSUBS 0.01257f
C588 VTAIL.n535 VSUBS 0.011871f
C589 VTAIL.n536 VSUBS 0.022092f
C590 VTAIL.n537 VSUBS 0.022092f
C591 VTAIL.n538 VSUBS 0.011871f
C592 VTAIL.n539 VSUBS 0.01257f
C593 VTAIL.n540 VSUBS 0.028059f
C594 VTAIL.n541 VSUBS 0.028059f
C595 VTAIL.n542 VSUBS 0.01257f
C596 VTAIL.n543 VSUBS 0.011871f
C597 VTAIL.n544 VSUBS 0.022092f
C598 VTAIL.n545 VSUBS 0.022092f
C599 VTAIL.n546 VSUBS 0.011871f
C600 VTAIL.n547 VSUBS 0.01222f
C601 VTAIL.n548 VSUBS 0.01222f
C602 VTAIL.n549 VSUBS 0.028059f
C603 VTAIL.n550 VSUBS 0.028059f
C604 VTAIL.n551 VSUBS 0.01257f
C605 VTAIL.n552 VSUBS 0.011871f
C606 VTAIL.n553 VSUBS 0.022092f
C607 VTAIL.n554 VSUBS 0.022092f
C608 VTAIL.n555 VSUBS 0.011871f
C609 VTAIL.n556 VSUBS 0.01257f
C610 VTAIL.n557 VSUBS 0.028059f
C611 VTAIL.n558 VSUBS 0.061234f
C612 VTAIL.n559 VSUBS 0.01257f
C613 VTAIL.n560 VSUBS 0.011871f
C614 VTAIL.n561 VSUBS 0.047443f
C615 VTAIL.n562 VSUBS 0.030382f
C616 VTAIL.n563 VSUBS 0.128822f
C617 VTAIL.n564 VSUBS 0.022309f
C618 VTAIL.n565 VSUBS 0.022092f
C619 VTAIL.n566 VSUBS 0.011871f
C620 VTAIL.n567 VSUBS 0.028059f
C621 VTAIL.n568 VSUBS 0.01257f
C622 VTAIL.n569 VSUBS 0.022092f
C623 VTAIL.n570 VSUBS 0.011871f
C624 VTAIL.n571 VSUBS 0.028059f
C625 VTAIL.n572 VSUBS 0.01257f
C626 VTAIL.n573 VSUBS 0.022092f
C627 VTAIL.n574 VSUBS 0.011871f
C628 VTAIL.n575 VSUBS 0.028059f
C629 VTAIL.n576 VSUBS 0.028059f
C630 VTAIL.n577 VSUBS 0.01257f
C631 VTAIL.n578 VSUBS 0.022092f
C632 VTAIL.n579 VSUBS 0.011871f
C633 VTAIL.n580 VSUBS 0.028059f
C634 VTAIL.n581 VSUBS 0.01257f
C635 VTAIL.n582 VSUBS 0.022092f
C636 VTAIL.n583 VSUBS 0.011871f
C637 VTAIL.n584 VSUBS 0.028059f
C638 VTAIL.n585 VSUBS 0.01257f
C639 VTAIL.n586 VSUBS 0.022092f
C640 VTAIL.n587 VSUBS 0.011871f
C641 VTAIL.n588 VSUBS 0.028059f
C642 VTAIL.n589 VSUBS 0.01257f
C643 VTAIL.n590 VSUBS 0.022092f
C644 VTAIL.n591 VSUBS 0.011871f
C645 VTAIL.n592 VSUBS 0.028059f
C646 VTAIL.n593 VSUBS 0.01257f
C647 VTAIL.n594 VSUBS 0.166676f
C648 VTAIL.t5 VSUBS 0.060162f
C649 VTAIL.n595 VSUBS 0.021045f
C650 VTAIL.n596 VSUBS 0.01785f
C651 VTAIL.n597 VSUBS 0.011871f
C652 VTAIL.n598 VSUBS 1.5791f
C653 VTAIL.n599 VSUBS 0.022092f
C654 VTAIL.n600 VSUBS 0.011871f
C655 VTAIL.n601 VSUBS 0.01257f
C656 VTAIL.n602 VSUBS 0.028059f
C657 VTAIL.n603 VSUBS 0.028059f
C658 VTAIL.n604 VSUBS 0.01257f
C659 VTAIL.n605 VSUBS 0.011871f
C660 VTAIL.n606 VSUBS 0.022092f
C661 VTAIL.n607 VSUBS 0.022092f
C662 VTAIL.n608 VSUBS 0.011871f
C663 VTAIL.n609 VSUBS 0.01257f
C664 VTAIL.n610 VSUBS 0.028059f
C665 VTAIL.n611 VSUBS 0.028059f
C666 VTAIL.n612 VSUBS 0.01257f
C667 VTAIL.n613 VSUBS 0.011871f
C668 VTAIL.n614 VSUBS 0.022092f
C669 VTAIL.n615 VSUBS 0.022092f
C670 VTAIL.n616 VSUBS 0.011871f
C671 VTAIL.n617 VSUBS 0.01257f
C672 VTAIL.n618 VSUBS 0.028059f
C673 VTAIL.n619 VSUBS 0.028059f
C674 VTAIL.n620 VSUBS 0.01257f
C675 VTAIL.n621 VSUBS 0.011871f
C676 VTAIL.n622 VSUBS 0.022092f
C677 VTAIL.n623 VSUBS 0.022092f
C678 VTAIL.n624 VSUBS 0.011871f
C679 VTAIL.n625 VSUBS 0.01257f
C680 VTAIL.n626 VSUBS 0.028059f
C681 VTAIL.n627 VSUBS 0.028059f
C682 VTAIL.n628 VSUBS 0.01257f
C683 VTAIL.n629 VSUBS 0.011871f
C684 VTAIL.n630 VSUBS 0.022092f
C685 VTAIL.n631 VSUBS 0.022092f
C686 VTAIL.n632 VSUBS 0.011871f
C687 VTAIL.n633 VSUBS 0.01257f
C688 VTAIL.n634 VSUBS 0.028059f
C689 VTAIL.n635 VSUBS 0.028059f
C690 VTAIL.n636 VSUBS 0.01257f
C691 VTAIL.n637 VSUBS 0.011871f
C692 VTAIL.n638 VSUBS 0.022092f
C693 VTAIL.n639 VSUBS 0.022092f
C694 VTAIL.n640 VSUBS 0.011871f
C695 VTAIL.n641 VSUBS 0.01222f
C696 VTAIL.n642 VSUBS 0.01222f
C697 VTAIL.n643 VSUBS 0.028059f
C698 VTAIL.n644 VSUBS 0.028059f
C699 VTAIL.n645 VSUBS 0.01257f
C700 VTAIL.n646 VSUBS 0.011871f
C701 VTAIL.n647 VSUBS 0.022092f
C702 VTAIL.n648 VSUBS 0.022092f
C703 VTAIL.n649 VSUBS 0.011871f
C704 VTAIL.n650 VSUBS 0.01257f
C705 VTAIL.n651 VSUBS 0.028059f
C706 VTAIL.n652 VSUBS 0.061234f
C707 VTAIL.n653 VSUBS 0.01257f
C708 VTAIL.n654 VSUBS 0.011871f
C709 VTAIL.n655 VSUBS 0.047443f
C710 VTAIL.n656 VSUBS 0.030382f
C711 VTAIL.n657 VSUBS 1.49761f
C712 VTAIL.n658 VSUBS 0.022309f
C713 VTAIL.n659 VSUBS 0.022092f
C714 VTAIL.n660 VSUBS 0.011871f
C715 VTAIL.n661 VSUBS 0.028059f
C716 VTAIL.n662 VSUBS 0.01257f
C717 VTAIL.n663 VSUBS 0.022092f
C718 VTAIL.n664 VSUBS 0.011871f
C719 VTAIL.n665 VSUBS 0.028059f
C720 VTAIL.n666 VSUBS 0.01257f
C721 VTAIL.n667 VSUBS 0.022092f
C722 VTAIL.n668 VSUBS 0.011871f
C723 VTAIL.n669 VSUBS 0.028059f
C724 VTAIL.n670 VSUBS 0.01257f
C725 VTAIL.n671 VSUBS 0.022092f
C726 VTAIL.n672 VSUBS 0.011871f
C727 VTAIL.n673 VSUBS 0.028059f
C728 VTAIL.n674 VSUBS 0.01257f
C729 VTAIL.n675 VSUBS 0.022092f
C730 VTAIL.n676 VSUBS 0.011871f
C731 VTAIL.n677 VSUBS 0.028059f
C732 VTAIL.n678 VSUBS 0.01257f
C733 VTAIL.n679 VSUBS 0.022092f
C734 VTAIL.n680 VSUBS 0.011871f
C735 VTAIL.n681 VSUBS 0.028059f
C736 VTAIL.n682 VSUBS 0.01257f
C737 VTAIL.n683 VSUBS 0.022092f
C738 VTAIL.n684 VSUBS 0.011871f
C739 VTAIL.n685 VSUBS 0.028059f
C740 VTAIL.n686 VSUBS 0.01257f
C741 VTAIL.n687 VSUBS 0.166676f
C742 VTAIL.t0 VSUBS 0.060162f
C743 VTAIL.n688 VSUBS 0.021045f
C744 VTAIL.n689 VSUBS 0.01785f
C745 VTAIL.n690 VSUBS 0.011871f
C746 VTAIL.n691 VSUBS 1.5791f
C747 VTAIL.n692 VSUBS 0.022092f
C748 VTAIL.n693 VSUBS 0.011871f
C749 VTAIL.n694 VSUBS 0.01257f
C750 VTAIL.n695 VSUBS 0.028059f
C751 VTAIL.n696 VSUBS 0.028059f
C752 VTAIL.n697 VSUBS 0.01257f
C753 VTAIL.n698 VSUBS 0.011871f
C754 VTAIL.n699 VSUBS 0.022092f
C755 VTAIL.n700 VSUBS 0.022092f
C756 VTAIL.n701 VSUBS 0.011871f
C757 VTAIL.n702 VSUBS 0.01257f
C758 VTAIL.n703 VSUBS 0.028059f
C759 VTAIL.n704 VSUBS 0.028059f
C760 VTAIL.n705 VSUBS 0.01257f
C761 VTAIL.n706 VSUBS 0.011871f
C762 VTAIL.n707 VSUBS 0.022092f
C763 VTAIL.n708 VSUBS 0.022092f
C764 VTAIL.n709 VSUBS 0.011871f
C765 VTAIL.n710 VSUBS 0.01257f
C766 VTAIL.n711 VSUBS 0.028059f
C767 VTAIL.n712 VSUBS 0.028059f
C768 VTAIL.n713 VSUBS 0.01257f
C769 VTAIL.n714 VSUBS 0.011871f
C770 VTAIL.n715 VSUBS 0.022092f
C771 VTAIL.n716 VSUBS 0.022092f
C772 VTAIL.n717 VSUBS 0.011871f
C773 VTAIL.n718 VSUBS 0.01257f
C774 VTAIL.n719 VSUBS 0.028059f
C775 VTAIL.n720 VSUBS 0.028059f
C776 VTAIL.n721 VSUBS 0.01257f
C777 VTAIL.n722 VSUBS 0.011871f
C778 VTAIL.n723 VSUBS 0.022092f
C779 VTAIL.n724 VSUBS 0.022092f
C780 VTAIL.n725 VSUBS 0.011871f
C781 VTAIL.n726 VSUBS 0.01257f
C782 VTAIL.n727 VSUBS 0.028059f
C783 VTAIL.n728 VSUBS 0.028059f
C784 VTAIL.n729 VSUBS 0.028059f
C785 VTAIL.n730 VSUBS 0.01257f
C786 VTAIL.n731 VSUBS 0.011871f
C787 VTAIL.n732 VSUBS 0.022092f
C788 VTAIL.n733 VSUBS 0.022092f
C789 VTAIL.n734 VSUBS 0.011871f
C790 VTAIL.n735 VSUBS 0.01222f
C791 VTAIL.n736 VSUBS 0.01222f
C792 VTAIL.n737 VSUBS 0.028059f
C793 VTAIL.n738 VSUBS 0.028059f
C794 VTAIL.n739 VSUBS 0.01257f
C795 VTAIL.n740 VSUBS 0.011871f
C796 VTAIL.n741 VSUBS 0.022092f
C797 VTAIL.n742 VSUBS 0.022092f
C798 VTAIL.n743 VSUBS 0.011871f
C799 VTAIL.n744 VSUBS 0.01257f
C800 VTAIL.n745 VSUBS 0.028059f
C801 VTAIL.n746 VSUBS 0.061234f
C802 VTAIL.n747 VSUBS 0.01257f
C803 VTAIL.n748 VSUBS 0.011871f
C804 VTAIL.n749 VSUBS 0.047443f
C805 VTAIL.n750 VSUBS 0.030382f
C806 VTAIL.n751 VSUBS 1.45419f
C807 VP.t1 VSUBS 2.3947f
C808 VP.t3 VSUBS 2.39488f
C809 VP.n0 VSUBS 3.2398f
C810 VP.n1 VSUBS 3.54396f
C811 VP.t2 VSUBS 2.36032f
C812 VP.n2 VSUBS 0.896805f
C813 VP.t0 VSUBS 2.36032f
C814 VP.n3 VSUBS 0.896805f
C815 VP.n4 VSUBS 0.06671f
C816 B.n0 VSUBS 0.006605f
C817 B.n1 VSUBS 0.006605f
C818 B.n2 VSUBS 0.009768f
C819 B.n3 VSUBS 0.007485f
C820 B.n4 VSUBS 0.007485f
C821 B.n5 VSUBS 0.007485f
C822 B.n6 VSUBS 0.007485f
C823 B.n7 VSUBS 0.007485f
C824 B.n8 VSUBS 0.007485f
C825 B.n9 VSUBS 0.007485f
C826 B.n10 VSUBS 0.007485f
C827 B.n11 VSUBS 0.0175f
C828 B.n12 VSUBS 0.007485f
C829 B.n13 VSUBS 0.007485f
C830 B.n14 VSUBS 0.007485f
C831 B.n15 VSUBS 0.007485f
C832 B.n16 VSUBS 0.007485f
C833 B.n17 VSUBS 0.007485f
C834 B.n18 VSUBS 0.007485f
C835 B.n19 VSUBS 0.007485f
C836 B.n20 VSUBS 0.007485f
C837 B.n21 VSUBS 0.007485f
C838 B.n22 VSUBS 0.007485f
C839 B.n23 VSUBS 0.007485f
C840 B.n24 VSUBS 0.007485f
C841 B.n25 VSUBS 0.007485f
C842 B.n26 VSUBS 0.007485f
C843 B.n27 VSUBS 0.007485f
C844 B.n28 VSUBS 0.007485f
C845 B.n29 VSUBS 0.007485f
C846 B.n30 VSUBS 0.007485f
C847 B.n31 VSUBS 0.007485f
C848 B.n32 VSUBS 0.007485f
C849 B.n33 VSUBS 0.007485f
C850 B.n34 VSUBS 0.007485f
C851 B.n35 VSUBS 0.007485f
C852 B.n36 VSUBS 0.007485f
C853 B.n37 VSUBS 0.007485f
C854 B.n38 VSUBS 0.007485f
C855 B.n39 VSUBS 0.007485f
C856 B.t4 VSUBS 0.341241f
C857 B.t5 VSUBS 0.357464f
C858 B.t3 VSUBS 0.699755f
C859 B.n40 VSUBS 0.468704f
C860 B.n41 VSUBS 0.327316f
C861 B.n42 VSUBS 0.007485f
C862 B.n43 VSUBS 0.007485f
C863 B.n44 VSUBS 0.007485f
C864 B.n45 VSUBS 0.007485f
C865 B.t1 VSUBS 0.341245f
C866 B.t2 VSUBS 0.357467f
C867 B.t0 VSUBS 0.699755f
C868 B.n46 VSUBS 0.4687f
C869 B.n47 VSUBS 0.327312f
C870 B.n48 VSUBS 0.017342f
C871 B.n49 VSUBS 0.007485f
C872 B.n50 VSUBS 0.007485f
C873 B.n51 VSUBS 0.007485f
C874 B.n52 VSUBS 0.007485f
C875 B.n53 VSUBS 0.007485f
C876 B.n54 VSUBS 0.007485f
C877 B.n55 VSUBS 0.007485f
C878 B.n56 VSUBS 0.007485f
C879 B.n57 VSUBS 0.007485f
C880 B.n58 VSUBS 0.007485f
C881 B.n59 VSUBS 0.007485f
C882 B.n60 VSUBS 0.007485f
C883 B.n61 VSUBS 0.007485f
C884 B.n62 VSUBS 0.007485f
C885 B.n63 VSUBS 0.007485f
C886 B.n64 VSUBS 0.007485f
C887 B.n65 VSUBS 0.007485f
C888 B.n66 VSUBS 0.007485f
C889 B.n67 VSUBS 0.007485f
C890 B.n68 VSUBS 0.007485f
C891 B.n69 VSUBS 0.007485f
C892 B.n70 VSUBS 0.007485f
C893 B.n71 VSUBS 0.007485f
C894 B.n72 VSUBS 0.007485f
C895 B.n73 VSUBS 0.007485f
C896 B.n74 VSUBS 0.007485f
C897 B.n75 VSUBS 0.007485f
C898 B.n76 VSUBS 0.0175f
C899 B.n77 VSUBS 0.007485f
C900 B.n78 VSUBS 0.007485f
C901 B.n79 VSUBS 0.007485f
C902 B.n80 VSUBS 0.007485f
C903 B.n81 VSUBS 0.007485f
C904 B.n82 VSUBS 0.007485f
C905 B.n83 VSUBS 0.007485f
C906 B.n84 VSUBS 0.007485f
C907 B.n85 VSUBS 0.007485f
C908 B.n86 VSUBS 0.007485f
C909 B.n87 VSUBS 0.007485f
C910 B.n88 VSUBS 0.007485f
C911 B.n89 VSUBS 0.007485f
C912 B.n90 VSUBS 0.007485f
C913 B.n91 VSUBS 0.007485f
C914 B.n92 VSUBS 0.007485f
C915 B.n93 VSUBS 0.007485f
C916 B.n94 VSUBS 0.007485f
C917 B.n95 VSUBS 0.007485f
C918 B.n96 VSUBS 0.017076f
C919 B.n97 VSUBS 0.007485f
C920 B.n98 VSUBS 0.007485f
C921 B.n99 VSUBS 0.007485f
C922 B.n100 VSUBS 0.007485f
C923 B.n101 VSUBS 0.007485f
C924 B.n102 VSUBS 0.007485f
C925 B.n103 VSUBS 0.007485f
C926 B.n104 VSUBS 0.007485f
C927 B.n105 VSUBS 0.007485f
C928 B.n106 VSUBS 0.007485f
C929 B.n107 VSUBS 0.007485f
C930 B.n108 VSUBS 0.007485f
C931 B.n109 VSUBS 0.007485f
C932 B.n110 VSUBS 0.007485f
C933 B.n111 VSUBS 0.007485f
C934 B.n112 VSUBS 0.007485f
C935 B.n113 VSUBS 0.007485f
C936 B.n114 VSUBS 0.007485f
C937 B.n115 VSUBS 0.007485f
C938 B.n116 VSUBS 0.007485f
C939 B.n117 VSUBS 0.007485f
C940 B.n118 VSUBS 0.007485f
C941 B.n119 VSUBS 0.007485f
C942 B.n120 VSUBS 0.007485f
C943 B.n121 VSUBS 0.007485f
C944 B.n122 VSUBS 0.007485f
C945 B.n123 VSUBS 0.007485f
C946 B.t8 VSUBS 0.341245f
C947 B.t7 VSUBS 0.357467f
C948 B.t6 VSUBS 0.699755f
C949 B.n124 VSUBS 0.4687f
C950 B.n125 VSUBS 0.327312f
C951 B.n126 VSUBS 0.007485f
C952 B.n127 VSUBS 0.007485f
C953 B.n128 VSUBS 0.007485f
C954 B.n129 VSUBS 0.007485f
C955 B.n130 VSUBS 0.004183f
C956 B.n131 VSUBS 0.007485f
C957 B.n132 VSUBS 0.007485f
C958 B.n133 VSUBS 0.007485f
C959 B.n134 VSUBS 0.007485f
C960 B.n135 VSUBS 0.007485f
C961 B.n136 VSUBS 0.007485f
C962 B.n137 VSUBS 0.007485f
C963 B.n138 VSUBS 0.007485f
C964 B.n139 VSUBS 0.007485f
C965 B.n140 VSUBS 0.007485f
C966 B.n141 VSUBS 0.007485f
C967 B.n142 VSUBS 0.007485f
C968 B.n143 VSUBS 0.007485f
C969 B.n144 VSUBS 0.007485f
C970 B.n145 VSUBS 0.007485f
C971 B.n146 VSUBS 0.007485f
C972 B.n147 VSUBS 0.007485f
C973 B.n148 VSUBS 0.007485f
C974 B.n149 VSUBS 0.007485f
C975 B.n150 VSUBS 0.007485f
C976 B.n151 VSUBS 0.007485f
C977 B.n152 VSUBS 0.007485f
C978 B.n153 VSUBS 0.007485f
C979 B.n154 VSUBS 0.007485f
C980 B.n155 VSUBS 0.007485f
C981 B.n156 VSUBS 0.007485f
C982 B.n157 VSUBS 0.007485f
C983 B.n158 VSUBS 0.0175f
C984 B.n159 VSUBS 0.007485f
C985 B.n160 VSUBS 0.007485f
C986 B.n161 VSUBS 0.007485f
C987 B.n162 VSUBS 0.007485f
C988 B.n163 VSUBS 0.007485f
C989 B.n164 VSUBS 0.007485f
C990 B.n165 VSUBS 0.007485f
C991 B.n166 VSUBS 0.007485f
C992 B.n167 VSUBS 0.007485f
C993 B.n168 VSUBS 0.007485f
C994 B.n169 VSUBS 0.007485f
C995 B.n170 VSUBS 0.007485f
C996 B.n171 VSUBS 0.007485f
C997 B.n172 VSUBS 0.007485f
C998 B.n173 VSUBS 0.007485f
C999 B.n174 VSUBS 0.007485f
C1000 B.n175 VSUBS 0.007485f
C1001 B.n176 VSUBS 0.007485f
C1002 B.n177 VSUBS 0.007485f
C1003 B.n178 VSUBS 0.007485f
C1004 B.n179 VSUBS 0.007485f
C1005 B.n180 VSUBS 0.007485f
C1006 B.n181 VSUBS 0.007485f
C1007 B.n182 VSUBS 0.007485f
C1008 B.n183 VSUBS 0.007485f
C1009 B.n184 VSUBS 0.007485f
C1010 B.n185 VSUBS 0.007485f
C1011 B.n186 VSUBS 0.007485f
C1012 B.n187 VSUBS 0.007485f
C1013 B.n188 VSUBS 0.007485f
C1014 B.n189 VSUBS 0.007485f
C1015 B.n190 VSUBS 0.007485f
C1016 B.n191 VSUBS 0.007485f
C1017 B.n192 VSUBS 0.007485f
C1018 B.n193 VSUBS 0.0175f
C1019 B.n194 VSUBS 0.017945f
C1020 B.n195 VSUBS 0.017945f
C1021 B.n196 VSUBS 0.007485f
C1022 B.n197 VSUBS 0.007485f
C1023 B.n198 VSUBS 0.007485f
C1024 B.n199 VSUBS 0.007485f
C1025 B.n200 VSUBS 0.007485f
C1026 B.n201 VSUBS 0.007485f
C1027 B.n202 VSUBS 0.007485f
C1028 B.n203 VSUBS 0.007485f
C1029 B.n204 VSUBS 0.007485f
C1030 B.n205 VSUBS 0.007485f
C1031 B.n206 VSUBS 0.007485f
C1032 B.n207 VSUBS 0.007485f
C1033 B.n208 VSUBS 0.007485f
C1034 B.n209 VSUBS 0.007485f
C1035 B.n210 VSUBS 0.007485f
C1036 B.n211 VSUBS 0.007485f
C1037 B.n212 VSUBS 0.007485f
C1038 B.n213 VSUBS 0.007485f
C1039 B.n214 VSUBS 0.007485f
C1040 B.n215 VSUBS 0.007485f
C1041 B.n216 VSUBS 0.007485f
C1042 B.n217 VSUBS 0.007485f
C1043 B.n218 VSUBS 0.007485f
C1044 B.n219 VSUBS 0.007485f
C1045 B.n220 VSUBS 0.007485f
C1046 B.n221 VSUBS 0.007485f
C1047 B.n222 VSUBS 0.007485f
C1048 B.n223 VSUBS 0.007485f
C1049 B.n224 VSUBS 0.007485f
C1050 B.n225 VSUBS 0.007485f
C1051 B.n226 VSUBS 0.007485f
C1052 B.n227 VSUBS 0.007485f
C1053 B.n228 VSUBS 0.007485f
C1054 B.n229 VSUBS 0.007485f
C1055 B.n230 VSUBS 0.007485f
C1056 B.n231 VSUBS 0.007485f
C1057 B.n232 VSUBS 0.007485f
C1058 B.n233 VSUBS 0.007485f
C1059 B.n234 VSUBS 0.007485f
C1060 B.n235 VSUBS 0.007485f
C1061 B.n236 VSUBS 0.007485f
C1062 B.n237 VSUBS 0.007485f
C1063 B.n238 VSUBS 0.007485f
C1064 B.n239 VSUBS 0.007485f
C1065 B.n240 VSUBS 0.007485f
C1066 B.n241 VSUBS 0.007485f
C1067 B.n242 VSUBS 0.007485f
C1068 B.n243 VSUBS 0.007485f
C1069 B.n244 VSUBS 0.007485f
C1070 B.n245 VSUBS 0.007485f
C1071 B.n246 VSUBS 0.007485f
C1072 B.n247 VSUBS 0.007485f
C1073 B.n248 VSUBS 0.007485f
C1074 B.n249 VSUBS 0.007485f
C1075 B.n250 VSUBS 0.007485f
C1076 B.n251 VSUBS 0.007485f
C1077 B.n252 VSUBS 0.007485f
C1078 B.n253 VSUBS 0.007485f
C1079 B.n254 VSUBS 0.007485f
C1080 B.n255 VSUBS 0.007485f
C1081 B.n256 VSUBS 0.007485f
C1082 B.n257 VSUBS 0.007485f
C1083 B.n258 VSUBS 0.007485f
C1084 B.n259 VSUBS 0.007485f
C1085 B.n260 VSUBS 0.007485f
C1086 B.n261 VSUBS 0.007485f
C1087 B.n262 VSUBS 0.007485f
C1088 B.n263 VSUBS 0.007485f
C1089 B.n264 VSUBS 0.007485f
C1090 B.n265 VSUBS 0.007485f
C1091 B.n266 VSUBS 0.007485f
C1092 B.n267 VSUBS 0.007485f
C1093 B.n268 VSUBS 0.007485f
C1094 B.n269 VSUBS 0.007485f
C1095 B.n270 VSUBS 0.007485f
C1096 B.n271 VSUBS 0.007485f
C1097 B.n272 VSUBS 0.007485f
C1098 B.n273 VSUBS 0.007485f
C1099 B.n274 VSUBS 0.007485f
C1100 B.t11 VSUBS 0.341241f
C1101 B.t10 VSUBS 0.357464f
C1102 B.t9 VSUBS 0.699755f
C1103 B.n275 VSUBS 0.468704f
C1104 B.n276 VSUBS 0.327316f
C1105 B.n277 VSUBS 0.017342f
C1106 B.n278 VSUBS 0.007045f
C1107 B.n279 VSUBS 0.007485f
C1108 B.n280 VSUBS 0.007485f
C1109 B.n281 VSUBS 0.007485f
C1110 B.n282 VSUBS 0.007485f
C1111 B.n283 VSUBS 0.007485f
C1112 B.n284 VSUBS 0.007485f
C1113 B.n285 VSUBS 0.007485f
C1114 B.n286 VSUBS 0.007485f
C1115 B.n287 VSUBS 0.007485f
C1116 B.n288 VSUBS 0.007485f
C1117 B.n289 VSUBS 0.007485f
C1118 B.n290 VSUBS 0.007485f
C1119 B.n291 VSUBS 0.007485f
C1120 B.n292 VSUBS 0.007485f
C1121 B.n293 VSUBS 0.007485f
C1122 B.n294 VSUBS 0.004183f
C1123 B.n295 VSUBS 0.017342f
C1124 B.n296 VSUBS 0.007045f
C1125 B.n297 VSUBS 0.007485f
C1126 B.n298 VSUBS 0.007485f
C1127 B.n299 VSUBS 0.007485f
C1128 B.n300 VSUBS 0.007485f
C1129 B.n301 VSUBS 0.007485f
C1130 B.n302 VSUBS 0.007485f
C1131 B.n303 VSUBS 0.007485f
C1132 B.n304 VSUBS 0.007485f
C1133 B.n305 VSUBS 0.007485f
C1134 B.n306 VSUBS 0.007485f
C1135 B.n307 VSUBS 0.007485f
C1136 B.n308 VSUBS 0.007485f
C1137 B.n309 VSUBS 0.007485f
C1138 B.n310 VSUBS 0.007485f
C1139 B.n311 VSUBS 0.007485f
C1140 B.n312 VSUBS 0.007485f
C1141 B.n313 VSUBS 0.007485f
C1142 B.n314 VSUBS 0.007485f
C1143 B.n315 VSUBS 0.007485f
C1144 B.n316 VSUBS 0.007485f
C1145 B.n317 VSUBS 0.007485f
C1146 B.n318 VSUBS 0.007485f
C1147 B.n319 VSUBS 0.007485f
C1148 B.n320 VSUBS 0.007485f
C1149 B.n321 VSUBS 0.007485f
C1150 B.n322 VSUBS 0.007485f
C1151 B.n323 VSUBS 0.007485f
C1152 B.n324 VSUBS 0.007485f
C1153 B.n325 VSUBS 0.007485f
C1154 B.n326 VSUBS 0.007485f
C1155 B.n327 VSUBS 0.007485f
C1156 B.n328 VSUBS 0.007485f
C1157 B.n329 VSUBS 0.007485f
C1158 B.n330 VSUBS 0.007485f
C1159 B.n331 VSUBS 0.007485f
C1160 B.n332 VSUBS 0.007485f
C1161 B.n333 VSUBS 0.007485f
C1162 B.n334 VSUBS 0.007485f
C1163 B.n335 VSUBS 0.007485f
C1164 B.n336 VSUBS 0.007485f
C1165 B.n337 VSUBS 0.007485f
C1166 B.n338 VSUBS 0.007485f
C1167 B.n339 VSUBS 0.007485f
C1168 B.n340 VSUBS 0.007485f
C1169 B.n341 VSUBS 0.007485f
C1170 B.n342 VSUBS 0.007485f
C1171 B.n343 VSUBS 0.007485f
C1172 B.n344 VSUBS 0.007485f
C1173 B.n345 VSUBS 0.007485f
C1174 B.n346 VSUBS 0.007485f
C1175 B.n347 VSUBS 0.007485f
C1176 B.n348 VSUBS 0.007485f
C1177 B.n349 VSUBS 0.007485f
C1178 B.n350 VSUBS 0.007485f
C1179 B.n351 VSUBS 0.007485f
C1180 B.n352 VSUBS 0.007485f
C1181 B.n353 VSUBS 0.007485f
C1182 B.n354 VSUBS 0.007485f
C1183 B.n355 VSUBS 0.007485f
C1184 B.n356 VSUBS 0.007485f
C1185 B.n357 VSUBS 0.007485f
C1186 B.n358 VSUBS 0.007485f
C1187 B.n359 VSUBS 0.007485f
C1188 B.n360 VSUBS 0.007485f
C1189 B.n361 VSUBS 0.007485f
C1190 B.n362 VSUBS 0.007485f
C1191 B.n363 VSUBS 0.007485f
C1192 B.n364 VSUBS 0.007485f
C1193 B.n365 VSUBS 0.007485f
C1194 B.n366 VSUBS 0.007485f
C1195 B.n367 VSUBS 0.007485f
C1196 B.n368 VSUBS 0.007485f
C1197 B.n369 VSUBS 0.007485f
C1198 B.n370 VSUBS 0.007485f
C1199 B.n371 VSUBS 0.007485f
C1200 B.n372 VSUBS 0.007485f
C1201 B.n373 VSUBS 0.007485f
C1202 B.n374 VSUBS 0.007485f
C1203 B.n375 VSUBS 0.007485f
C1204 B.n376 VSUBS 0.007485f
C1205 B.n377 VSUBS 0.017945f
C1206 B.n378 VSUBS 0.0175f
C1207 B.n379 VSUBS 0.018368f
C1208 B.n380 VSUBS 0.007485f
C1209 B.n381 VSUBS 0.007485f
C1210 B.n382 VSUBS 0.007485f
C1211 B.n383 VSUBS 0.007485f
C1212 B.n384 VSUBS 0.007485f
C1213 B.n385 VSUBS 0.007485f
C1214 B.n386 VSUBS 0.007485f
C1215 B.n387 VSUBS 0.007485f
C1216 B.n388 VSUBS 0.007485f
C1217 B.n389 VSUBS 0.007485f
C1218 B.n390 VSUBS 0.007485f
C1219 B.n391 VSUBS 0.007485f
C1220 B.n392 VSUBS 0.007485f
C1221 B.n393 VSUBS 0.007485f
C1222 B.n394 VSUBS 0.007485f
C1223 B.n395 VSUBS 0.007485f
C1224 B.n396 VSUBS 0.007485f
C1225 B.n397 VSUBS 0.007485f
C1226 B.n398 VSUBS 0.007485f
C1227 B.n399 VSUBS 0.007485f
C1228 B.n400 VSUBS 0.007485f
C1229 B.n401 VSUBS 0.007485f
C1230 B.n402 VSUBS 0.007485f
C1231 B.n403 VSUBS 0.007485f
C1232 B.n404 VSUBS 0.007485f
C1233 B.n405 VSUBS 0.007485f
C1234 B.n406 VSUBS 0.007485f
C1235 B.n407 VSUBS 0.007485f
C1236 B.n408 VSUBS 0.007485f
C1237 B.n409 VSUBS 0.007485f
C1238 B.n410 VSUBS 0.007485f
C1239 B.n411 VSUBS 0.007485f
C1240 B.n412 VSUBS 0.007485f
C1241 B.n413 VSUBS 0.007485f
C1242 B.n414 VSUBS 0.007485f
C1243 B.n415 VSUBS 0.007485f
C1244 B.n416 VSUBS 0.007485f
C1245 B.n417 VSUBS 0.007485f
C1246 B.n418 VSUBS 0.007485f
C1247 B.n419 VSUBS 0.007485f
C1248 B.n420 VSUBS 0.007485f
C1249 B.n421 VSUBS 0.007485f
C1250 B.n422 VSUBS 0.007485f
C1251 B.n423 VSUBS 0.007485f
C1252 B.n424 VSUBS 0.007485f
C1253 B.n425 VSUBS 0.007485f
C1254 B.n426 VSUBS 0.007485f
C1255 B.n427 VSUBS 0.007485f
C1256 B.n428 VSUBS 0.007485f
C1257 B.n429 VSUBS 0.007485f
C1258 B.n430 VSUBS 0.007485f
C1259 B.n431 VSUBS 0.007485f
C1260 B.n432 VSUBS 0.007485f
C1261 B.n433 VSUBS 0.007485f
C1262 B.n434 VSUBS 0.007485f
C1263 B.n435 VSUBS 0.007485f
C1264 B.n436 VSUBS 0.007485f
C1265 B.n437 VSUBS 0.0175f
C1266 B.n438 VSUBS 0.017945f
C1267 B.n439 VSUBS 0.017945f
C1268 B.n440 VSUBS 0.007485f
C1269 B.n441 VSUBS 0.007485f
C1270 B.n442 VSUBS 0.007485f
C1271 B.n443 VSUBS 0.007485f
C1272 B.n444 VSUBS 0.007485f
C1273 B.n445 VSUBS 0.007485f
C1274 B.n446 VSUBS 0.007485f
C1275 B.n447 VSUBS 0.007485f
C1276 B.n448 VSUBS 0.007485f
C1277 B.n449 VSUBS 0.007485f
C1278 B.n450 VSUBS 0.007485f
C1279 B.n451 VSUBS 0.007485f
C1280 B.n452 VSUBS 0.007485f
C1281 B.n453 VSUBS 0.007485f
C1282 B.n454 VSUBS 0.007485f
C1283 B.n455 VSUBS 0.007485f
C1284 B.n456 VSUBS 0.007485f
C1285 B.n457 VSUBS 0.007485f
C1286 B.n458 VSUBS 0.007485f
C1287 B.n459 VSUBS 0.007485f
C1288 B.n460 VSUBS 0.007485f
C1289 B.n461 VSUBS 0.007485f
C1290 B.n462 VSUBS 0.007485f
C1291 B.n463 VSUBS 0.007485f
C1292 B.n464 VSUBS 0.007485f
C1293 B.n465 VSUBS 0.007485f
C1294 B.n466 VSUBS 0.007485f
C1295 B.n467 VSUBS 0.007485f
C1296 B.n468 VSUBS 0.007485f
C1297 B.n469 VSUBS 0.007485f
C1298 B.n470 VSUBS 0.007485f
C1299 B.n471 VSUBS 0.007485f
C1300 B.n472 VSUBS 0.007485f
C1301 B.n473 VSUBS 0.007485f
C1302 B.n474 VSUBS 0.007485f
C1303 B.n475 VSUBS 0.007485f
C1304 B.n476 VSUBS 0.007485f
C1305 B.n477 VSUBS 0.007485f
C1306 B.n478 VSUBS 0.007485f
C1307 B.n479 VSUBS 0.007485f
C1308 B.n480 VSUBS 0.007485f
C1309 B.n481 VSUBS 0.007485f
C1310 B.n482 VSUBS 0.007485f
C1311 B.n483 VSUBS 0.007485f
C1312 B.n484 VSUBS 0.007485f
C1313 B.n485 VSUBS 0.007485f
C1314 B.n486 VSUBS 0.007485f
C1315 B.n487 VSUBS 0.007485f
C1316 B.n488 VSUBS 0.007485f
C1317 B.n489 VSUBS 0.007485f
C1318 B.n490 VSUBS 0.007485f
C1319 B.n491 VSUBS 0.007485f
C1320 B.n492 VSUBS 0.007485f
C1321 B.n493 VSUBS 0.007485f
C1322 B.n494 VSUBS 0.007485f
C1323 B.n495 VSUBS 0.007485f
C1324 B.n496 VSUBS 0.007485f
C1325 B.n497 VSUBS 0.007485f
C1326 B.n498 VSUBS 0.007485f
C1327 B.n499 VSUBS 0.007485f
C1328 B.n500 VSUBS 0.007485f
C1329 B.n501 VSUBS 0.007485f
C1330 B.n502 VSUBS 0.007485f
C1331 B.n503 VSUBS 0.007485f
C1332 B.n504 VSUBS 0.007485f
C1333 B.n505 VSUBS 0.007485f
C1334 B.n506 VSUBS 0.007485f
C1335 B.n507 VSUBS 0.007485f
C1336 B.n508 VSUBS 0.007485f
C1337 B.n509 VSUBS 0.007485f
C1338 B.n510 VSUBS 0.007485f
C1339 B.n511 VSUBS 0.007485f
C1340 B.n512 VSUBS 0.007485f
C1341 B.n513 VSUBS 0.007485f
C1342 B.n514 VSUBS 0.007485f
C1343 B.n515 VSUBS 0.007485f
C1344 B.n516 VSUBS 0.007485f
C1345 B.n517 VSUBS 0.007485f
C1346 B.n518 VSUBS 0.007485f
C1347 B.n519 VSUBS 0.007045f
C1348 B.n520 VSUBS 0.007485f
C1349 B.n521 VSUBS 0.007485f
C1350 B.n522 VSUBS 0.004183f
C1351 B.n523 VSUBS 0.007485f
C1352 B.n524 VSUBS 0.007485f
C1353 B.n525 VSUBS 0.007485f
C1354 B.n526 VSUBS 0.007485f
C1355 B.n527 VSUBS 0.007485f
C1356 B.n528 VSUBS 0.007485f
C1357 B.n529 VSUBS 0.007485f
C1358 B.n530 VSUBS 0.007485f
C1359 B.n531 VSUBS 0.007485f
C1360 B.n532 VSUBS 0.007485f
C1361 B.n533 VSUBS 0.007485f
C1362 B.n534 VSUBS 0.007485f
C1363 B.n535 VSUBS 0.004183f
C1364 B.n536 VSUBS 0.017342f
C1365 B.n537 VSUBS 0.007045f
C1366 B.n538 VSUBS 0.007485f
C1367 B.n539 VSUBS 0.007485f
C1368 B.n540 VSUBS 0.007485f
C1369 B.n541 VSUBS 0.007485f
C1370 B.n542 VSUBS 0.007485f
C1371 B.n543 VSUBS 0.007485f
C1372 B.n544 VSUBS 0.007485f
C1373 B.n545 VSUBS 0.007485f
C1374 B.n546 VSUBS 0.007485f
C1375 B.n547 VSUBS 0.007485f
C1376 B.n548 VSUBS 0.007485f
C1377 B.n549 VSUBS 0.007485f
C1378 B.n550 VSUBS 0.007485f
C1379 B.n551 VSUBS 0.007485f
C1380 B.n552 VSUBS 0.007485f
C1381 B.n553 VSUBS 0.007485f
C1382 B.n554 VSUBS 0.007485f
C1383 B.n555 VSUBS 0.007485f
C1384 B.n556 VSUBS 0.007485f
C1385 B.n557 VSUBS 0.007485f
C1386 B.n558 VSUBS 0.007485f
C1387 B.n559 VSUBS 0.007485f
C1388 B.n560 VSUBS 0.007485f
C1389 B.n561 VSUBS 0.007485f
C1390 B.n562 VSUBS 0.007485f
C1391 B.n563 VSUBS 0.007485f
C1392 B.n564 VSUBS 0.007485f
C1393 B.n565 VSUBS 0.007485f
C1394 B.n566 VSUBS 0.007485f
C1395 B.n567 VSUBS 0.007485f
C1396 B.n568 VSUBS 0.007485f
C1397 B.n569 VSUBS 0.007485f
C1398 B.n570 VSUBS 0.007485f
C1399 B.n571 VSUBS 0.007485f
C1400 B.n572 VSUBS 0.007485f
C1401 B.n573 VSUBS 0.007485f
C1402 B.n574 VSUBS 0.007485f
C1403 B.n575 VSUBS 0.007485f
C1404 B.n576 VSUBS 0.007485f
C1405 B.n577 VSUBS 0.007485f
C1406 B.n578 VSUBS 0.007485f
C1407 B.n579 VSUBS 0.007485f
C1408 B.n580 VSUBS 0.007485f
C1409 B.n581 VSUBS 0.007485f
C1410 B.n582 VSUBS 0.007485f
C1411 B.n583 VSUBS 0.007485f
C1412 B.n584 VSUBS 0.007485f
C1413 B.n585 VSUBS 0.007485f
C1414 B.n586 VSUBS 0.007485f
C1415 B.n587 VSUBS 0.007485f
C1416 B.n588 VSUBS 0.007485f
C1417 B.n589 VSUBS 0.007485f
C1418 B.n590 VSUBS 0.007485f
C1419 B.n591 VSUBS 0.007485f
C1420 B.n592 VSUBS 0.007485f
C1421 B.n593 VSUBS 0.007485f
C1422 B.n594 VSUBS 0.007485f
C1423 B.n595 VSUBS 0.007485f
C1424 B.n596 VSUBS 0.007485f
C1425 B.n597 VSUBS 0.007485f
C1426 B.n598 VSUBS 0.007485f
C1427 B.n599 VSUBS 0.007485f
C1428 B.n600 VSUBS 0.007485f
C1429 B.n601 VSUBS 0.007485f
C1430 B.n602 VSUBS 0.007485f
C1431 B.n603 VSUBS 0.007485f
C1432 B.n604 VSUBS 0.007485f
C1433 B.n605 VSUBS 0.007485f
C1434 B.n606 VSUBS 0.007485f
C1435 B.n607 VSUBS 0.007485f
C1436 B.n608 VSUBS 0.007485f
C1437 B.n609 VSUBS 0.007485f
C1438 B.n610 VSUBS 0.007485f
C1439 B.n611 VSUBS 0.007485f
C1440 B.n612 VSUBS 0.007485f
C1441 B.n613 VSUBS 0.007485f
C1442 B.n614 VSUBS 0.007485f
C1443 B.n615 VSUBS 0.007485f
C1444 B.n616 VSUBS 0.007485f
C1445 B.n617 VSUBS 0.007485f
C1446 B.n618 VSUBS 0.017945f
C1447 B.n619 VSUBS 0.017945f
C1448 B.n620 VSUBS 0.0175f
C1449 B.n621 VSUBS 0.007485f
C1450 B.n622 VSUBS 0.007485f
C1451 B.n623 VSUBS 0.007485f
C1452 B.n624 VSUBS 0.007485f
C1453 B.n625 VSUBS 0.007485f
C1454 B.n626 VSUBS 0.007485f
C1455 B.n627 VSUBS 0.007485f
C1456 B.n628 VSUBS 0.007485f
C1457 B.n629 VSUBS 0.007485f
C1458 B.n630 VSUBS 0.007485f
C1459 B.n631 VSUBS 0.007485f
C1460 B.n632 VSUBS 0.007485f
C1461 B.n633 VSUBS 0.007485f
C1462 B.n634 VSUBS 0.007485f
C1463 B.n635 VSUBS 0.007485f
C1464 B.n636 VSUBS 0.007485f
C1465 B.n637 VSUBS 0.007485f
C1466 B.n638 VSUBS 0.007485f
C1467 B.n639 VSUBS 0.007485f
C1468 B.n640 VSUBS 0.007485f
C1469 B.n641 VSUBS 0.007485f
C1470 B.n642 VSUBS 0.007485f
C1471 B.n643 VSUBS 0.007485f
C1472 B.n644 VSUBS 0.007485f
C1473 B.n645 VSUBS 0.007485f
C1474 B.n646 VSUBS 0.007485f
C1475 B.n647 VSUBS 0.009768f
C1476 B.n648 VSUBS 0.010405f
C1477 B.n649 VSUBS 0.020691f
.ends

