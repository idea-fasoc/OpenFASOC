* NGSPICE file created from diff_pair_sample_0047.ext - technology: sky130A

.subckt diff_pair_sample_0047 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=1.16985 ps=7.42 w=7.09 l=3.1
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=3.1
X2 VTAIL.t2 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=1.16985 ps=7.42 w=7.09 l=3.1
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=3.1
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=3.1
X5 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.16985 pd=7.42 as=2.7651 ps=14.96 w=7.09 l=3.1
X6 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=1.16985 ps=7.42 w=7.09 l=3.1
X7 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.16985 pd=7.42 as=2.7651 ps=14.96 w=7.09 l=3.1
X8 VDD2.t2 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.16985 pd=7.42 as=2.7651 ps=14.96 w=7.09 l=3.1
X9 VTAIL.t5 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=1.16985 ps=7.42 w=7.09 l=3.1
X10 VDD2.t0 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.16985 pd=7.42 as=2.7651 ps=14.96 w=7.09 l=3.1
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=3.1
R0 VN.n1 VN.t1 89.6304
R1 VN.n0 VN.t2 89.6304
R2 VN.n0 VN.t3 88.6156
R3 VN.n1 VN.t0 88.6156
R4 VN VN.n1 47.236
R5 VN VN.n0 2.83069
R6 VDD2.n2 VDD2.n0 104.502
R7 VDD2.n2 VDD2.n1 65.805
R8 VDD2.n1 VDD2.t3 2.79317
R9 VDD2.n1 VDD2.t2 2.79317
R10 VDD2.n0 VDD2.t1 2.79317
R11 VDD2.n0 VDD2.t0 2.79317
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t2 51.9191
R14 VTAIL.n4 VTAIL.t6 51.9191
R15 VTAIL.n3 VTAIL.t7 51.9191
R16 VTAIL.n6 VTAIL.t0 51.9188
R17 VTAIL.n7 VTAIL.t4 51.9188
R18 VTAIL.n0 VTAIL.t5 51.9188
R19 VTAIL.n1 VTAIL.t3 51.9188
R20 VTAIL.n2 VTAIL.t1 51.9188
R21 VTAIL.n7 VTAIL.n6 21.4358
R22 VTAIL.n3 VTAIL.n2 21.4358
R23 VTAIL.n4 VTAIL.n3 2.9574
R24 VTAIL.n6 VTAIL.n5 2.9574
R25 VTAIL.n2 VTAIL.n1 2.9574
R26 VTAIL VTAIL.n0 1.53714
R27 VTAIL VTAIL.n7 1.42076
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n514 B.n513 585
R31 B.n516 B.n109 585
R32 B.n519 B.n518 585
R33 B.n520 B.n108 585
R34 B.n522 B.n521 585
R35 B.n524 B.n107 585
R36 B.n527 B.n526 585
R37 B.n528 B.n106 585
R38 B.n530 B.n529 585
R39 B.n532 B.n105 585
R40 B.n535 B.n534 585
R41 B.n536 B.n104 585
R42 B.n538 B.n537 585
R43 B.n540 B.n103 585
R44 B.n543 B.n542 585
R45 B.n544 B.n102 585
R46 B.n546 B.n545 585
R47 B.n548 B.n101 585
R48 B.n551 B.n550 585
R49 B.n552 B.n100 585
R50 B.n554 B.n553 585
R51 B.n556 B.n99 585
R52 B.n559 B.n558 585
R53 B.n560 B.n98 585
R54 B.n562 B.n561 585
R55 B.n564 B.n97 585
R56 B.n567 B.n566 585
R57 B.n569 B.n94 585
R58 B.n571 B.n570 585
R59 B.n573 B.n93 585
R60 B.n576 B.n575 585
R61 B.n577 B.n92 585
R62 B.n579 B.n578 585
R63 B.n581 B.n91 585
R64 B.n584 B.n583 585
R65 B.n585 B.n87 585
R66 B.n587 B.n586 585
R67 B.n589 B.n86 585
R68 B.n592 B.n591 585
R69 B.n593 B.n85 585
R70 B.n595 B.n594 585
R71 B.n597 B.n84 585
R72 B.n600 B.n599 585
R73 B.n601 B.n83 585
R74 B.n603 B.n602 585
R75 B.n605 B.n82 585
R76 B.n608 B.n607 585
R77 B.n609 B.n81 585
R78 B.n611 B.n610 585
R79 B.n613 B.n80 585
R80 B.n616 B.n615 585
R81 B.n617 B.n79 585
R82 B.n619 B.n618 585
R83 B.n621 B.n78 585
R84 B.n624 B.n623 585
R85 B.n625 B.n77 585
R86 B.n627 B.n626 585
R87 B.n629 B.n76 585
R88 B.n632 B.n631 585
R89 B.n633 B.n75 585
R90 B.n635 B.n634 585
R91 B.n637 B.n74 585
R92 B.n640 B.n639 585
R93 B.n641 B.n73 585
R94 B.n512 B.n71 585
R95 B.n644 B.n71 585
R96 B.n511 B.n70 585
R97 B.n645 B.n70 585
R98 B.n510 B.n69 585
R99 B.n646 B.n69 585
R100 B.n509 B.n508 585
R101 B.n508 B.n65 585
R102 B.n507 B.n64 585
R103 B.n652 B.n64 585
R104 B.n506 B.n63 585
R105 B.n653 B.n63 585
R106 B.n505 B.n62 585
R107 B.n654 B.n62 585
R108 B.n504 B.n503 585
R109 B.n503 B.n58 585
R110 B.n502 B.n57 585
R111 B.n660 B.n57 585
R112 B.n501 B.n56 585
R113 B.n661 B.n56 585
R114 B.n500 B.n55 585
R115 B.n662 B.n55 585
R116 B.n499 B.n498 585
R117 B.n498 B.n51 585
R118 B.n497 B.n50 585
R119 B.n668 B.n50 585
R120 B.n496 B.n49 585
R121 B.n669 B.n49 585
R122 B.n495 B.n48 585
R123 B.n670 B.n48 585
R124 B.n494 B.n493 585
R125 B.n493 B.n44 585
R126 B.n492 B.n43 585
R127 B.n676 B.n43 585
R128 B.n491 B.n42 585
R129 B.n677 B.n42 585
R130 B.n490 B.n41 585
R131 B.n678 B.n41 585
R132 B.n489 B.n488 585
R133 B.n488 B.n37 585
R134 B.n487 B.n36 585
R135 B.n684 B.n36 585
R136 B.n486 B.n35 585
R137 B.n685 B.n35 585
R138 B.n485 B.n34 585
R139 B.n686 B.n34 585
R140 B.n484 B.n483 585
R141 B.n483 B.n30 585
R142 B.n482 B.n29 585
R143 B.n692 B.n29 585
R144 B.n481 B.n28 585
R145 B.n693 B.n28 585
R146 B.n480 B.n27 585
R147 B.n694 B.n27 585
R148 B.n479 B.n478 585
R149 B.n478 B.n23 585
R150 B.n477 B.n22 585
R151 B.n700 B.n22 585
R152 B.n476 B.n21 585
R153 B.n701 B.n21 585
R154 B.n475 B.n20 585
R155 B.n702 B.n20 585
R156 B.n474 B.n473 585
R157 B.n473 B.n19 585
R158 B.n472 B.n15 585
R159 B.n708 B.n15 585
R160 B.n471 B.n14 585
R161 B.n709 B.n14 585
R162 B.n470 B.n13 585
R163 B.n710 B.n13 585
R164 B.n469 B.n468 585
R165 B.n468 B.n12 585
R166 B.n467 B.n466 585
R167 B.n467 B.n8 585
R168 B.n465 B.n7 585
R169 B.n717 B.n7 585
R170 B.n464 B.n6 585
R171 B.n718 B.n6 585
R172 B.n463 B.n5 585
R173 B.n719 B.n5 585
R174 B.n462 B.n461 585
R175 B.n461 B.n4 585
R176 B.n460 B.n110 585
R177 B.n460 B.n459 585
R178 B.n450 B.n111 585
R179 B.n112 B.n111 585
R180 B.n452 B.n451 585
R181 B.n453 B.n452 585
R182 B.n449 B.n117 585
R183 B.n117 B.n116 585
R184 B.n448 B.n447 585
R185 B.n447 B.n446 585
R186 B.n119 B.n118 585
R187 B.n439 B.n119 585
R188 B.n438 B.n437 585
R189 B.n440 B.n438 585
R190 B.n436 B.n124 585
R191 B.n124 B.n123 585
R192 B.n435 B.n434 585
R193 B.n434 B.n433 585
R194 B.n126 B.n125 585
R195 B.n127 B.n126 585
R196 B.n426 B.n425 585
R197 B.n427 B.n426 585
R198 B.n424 B.n132 585
R199 B.n132 B.n131 585
R200 B.n423 B.n422 585
R201 B.n422 B.n421 585
R202 B.n134 B.n133 585
R203 B.n135 B.n134 585
R204 B.n414 B.n413 585
R205 B.n415 B.n414 585
R206 B.n412 B.n139 585
R207 B.n143 B.n139 585
R208 B.n411 B.n410 585
R209 B.n410 B.n409 585
R210 B.n141 B.n140 585
R211 B.n142 B.n141 585
R212 B.n402 B.n401 585
R213 B.n403 B.n402 585
R214 B.n400 B.n148 585
R215 B.n148 B.n147 585
R216 B.n399 B.n398 585
R217 B.n398 B.n397 585
R218 B.n150 B.n149 585
R219 B.n151 B.n150 585
R220 B.n390 B.n389 585
R221 B.n391 B.n390 585
R222 B.n388 B.n156 585
R223 B.n156 B.n155 585
R224 B.n387 B.n386 585
R225 B.n386 B.n385 585
R226 B.n158 B.n157 585
R227 B.n159 B.n158 585
R228 B.n378 B.n377 585
R229 B.n379 B.n378 585
R230 B.n376 B.n164 585
R231 B.n164 B.n163 585
R232 B.n375 B.n374 585
R233 B.n374 B.n373 585
R234 B.n166 B.n165 585
R235 B.n167 B.n166 585
R236 B.n366 B.n365 585
R237 B.n367 B.n366 585
R238 B.n364 B.n172 585
R239 B.n172 B.n171 585
R240 B.n363 B.n362 585
R241 B.n362 B.n361 585
R242 B.n174 B.n173 585
R243 B.n175 B.n174 585
R244 B.n354 B.n353 585
R245 B.n355 B.n354 585
R246 B.n352 B.n180 585
R247 B.n180 B.n179 585
R248 B.n351 B.n350 585
R249 B.n350 B.n349 585
R250 B.n346 B.n184 585
R251 B.n345 B.n344 585
R252 B.n342 B.n185 585
R253 B.n342 B.n183 585
R254 B.n341 B.n340 585
R255 B.n339 B.n338 585
R256 B.n337 B.n187 585
R257 B.n335 B.n334 585
R258 B.n333 B.n188 585
R259 B.n332 B.n331 585
R260 B.n329 B.n189 585
R261 B.n327 B.n326 585
R262 B.n325 B.n190 585
R263 B.n324 B.n323 585
R264 B.n321 B.n191 585
R265 B.n319 B.n318 585
R266 B.n317 B.n192 585
R267 B.n316 B.n315 585
R268 B.n313 B.n193 585
R269 B.n311 B.n310 585
R270 B.n309 B.n194 585
R271 B.n308 B.n307 585
R272 B.n305 B.n195 585
R273 B.n303 B.n302 585
R274 B.n301 B.n196 585
R275 B.n300 B.n299 585
R276 B.n297 B.n197 585
R277 B.n295 B.n294 585
R278 B.n292 B.n198 585
R279 B.n291 B.n290 585
R280 B.n288 B.n201 585
R281 B.n286 B.n285 585
R282 B.n284 B.n202 585
R283 B.n283 B.n282 585
R284 B.n280 B.n203 585
R285 B.n278 B.n277 585
R286 B.n276 B.n204 585
R287 B.n275 B.n274 585
R288 B.n272 B.n271 585
R289 B.n270 B.n269 585
R290 B.n268 B.n209 585
R291 B.n266 B.n265 585
R292 B.n264 B.n210 585
R293 B.n263 B.n262 585
R294 B.n260 B.n211 585
R295 B.n258 B.n257 585
R296 B.n256 B.n212 585
R297 B.n255 B.n254 585
R298 B.n252 B.n213 585
R299 B.n250 B.n249 585
R300 B.n248 B.n214 585
R301 B.n247 B.n246 585
R302 B.n244 B.n215 585
R303 B.n242 B.n241 585
R304 B.n240 B.n216 585
R305 B.n239 B.n238 585
R306 B.n236 B.n217 585
R307 B.n234 B.n233 585
R308 B.n232 B.n218 585
R309 B.n231 B.n230 585
R310 B.n228 B.n219 585
R311 B.n226 B.n225 585
R312 B.n224 B.n220 585
R313 B.n223 B.n222 585
R314 B.n182 B.n181 585
R315 B.n183 B.n182 585
R316 B.n348 B.n347 585
R317 B.n349 B.n348 585
R318 B.n178 B.n177 585
R319 B.n179 B.n178 585
R320 B.n357 B.n356 585
R321 B.n356 B.n355 585
R322 B.n358 B.n176 585
R323 B.n176 B.n175 585
R324 B.n360 B.n359 585
R325 B.n361 B.n360 585
R326 B.n170 B.n169 585
R327 B.n171 B.n170 585
R328 B.n369 B.n368 585
R329 B.n368 B.n367 585
R330 B.n370 B.n168 585
R331 B.n168 B.n167 585
R332 B.n372 B.n371 585
R333 B.n373 B.n372 585
R334 B.n162 B.n161 585
R335 B.n163 B.n162 585
R336 B.n381 B.n380 585
R337 B.n380 B.n379 585
R338 B.n382 B.n160 585
R339 B.n160 B.n159 585
R340 B.n384 B.n383 585
R341 B.n385 B.n384 585
R342 B.n154 B.n153 585
R343 B.n155 B.n154 585
R344 B.n393 B.n392 585
R345 B.n392 B.n391 585
R346 B.n394 B.n152 585
R347 B.n152 B.n151 585
R348 B.n396 B.n395 585
R349 B.n397 B.n396 585
R350 B.n146 B.n145 585
R351 B.n147 B.n146 585
R352 B.n405 B.n404 585
R353 B.n404 B.n403 585
R354 B.n406 B.n144 585
R355 B.n144 B.n142 585
R356 B.n408 B.n407 585
R357 B.n409 B.n408 585
R358 B.n138 B.n137 585
R359 B.n143 B.n138 585
R360 B.n417 B.n416 585
R361 B.n416 B.n415 585
R362 B.n418 B.n136 585
R363 B.n136 B.n135 585
R364 B.n420 B.n419 585
R365 B.n421 B.n420 585
R366 B.n130 B.n129 585
R367 B.n131 B.n130 585
R368 B.n429 B.n428 585
R369 B.n428 B.n427 585
R370 B.n430 B.n128 585
R371 B.n128 B.n127 585
R372 B.n432 B.n431 585
R373 B.n433 B.n432 585
R374 B.n122 B.n121 585
R375 B.n123 B.n122 585
R376 B.n442 B.n441 585
R377 B.n441 B.n440 585
R378 B.n443 B.n120 585
R379 B.n439 B.n120 585
R380 B.n445 B.n444 585
R381 B.n446 B.n445 585
R382 B.n115 B.n114 585
R383 B.n116 B.n115 585
R384 B.n455 B.n454 585
R385 B.n454 B.n453 585
R386 B.n456 B.n113 585
R387 B.n113 B.n112 585
R388 B.n458 B.n457 585
R389 B.n459 B.n458 585
R390 B.n3 B.n0 585
R391 B.n4 B.n3 585
R392 B.n716 B.n1 585
R393 B.n717 B.n716 585
R394 B.n715 B.n714 585
R395 B.n715 B.n8 585
R396 B.n713 B.n9 585
R397 B.n12 B.n9 585
R398 B.n712 B.n711 585
R399 B.n711 B.n710 585
R400 B.n11 B.n10 585
R401 B.n709 B.n11 585
R402 B.n707 B.n706 585
R403 B.n708 B.n707 585
R404 B.n705 B.n16 585
R405 B.n19 B.n16 585
R406 B.n704 B.n703 585
R407 B.n703 B.n702 585
R408 B.n18 B.n17 585
R409 B.n701 B.n18 585
R410 B.n699 B.n698 585
R411 B.n700 B.n699 585
R412 B.n697 B.n24 585
R413 B.n24 B.n23 585
R414 B.n696 B.n695 585
R415 B.n695 B.n694 585
R416 B.n26 B.n25 585
R417 B.n693 B.n26 585
R418 B.n691 B.n690 585
R419 B.n692 B.n691 585
R420 B.n689 B.n31 585
R421 B.n31 B.n30 585
R422 B.n688 B.n687 585
R423 B.n687 B.n686 585
R424 B.n33 B.n32 585
R425 B.n685 B.n33 585
R426 B.n683 B.n682 585
R427 B.n684 B.n683 585
R428 B.n681 B.n38 585
R429 B.n38 B.n37 585
R430 B.n680 B.n679 585
R431 B.n679 B.n678 585
R432 B.n40 B.n39 585
R433 B.n677 B.n40 585
R434 B.n675 B.n674 585
R435 B.n676 B.n675 585
R436 B.n673 B.n45 585
R437 B.n45 B.n44 585
R438 B.n672 B.n671 585
R439 B.n671 B.n670 585
R440 B.n47 B.n46 585
R441 B.n669 B.n47 585
R442 B.n667 B.n666 585
R443 B.n668 B.n667 585
R444 B.n665 B.n52 585
R445 B.n52 B.n51 585
R446 B.n664 B.n663 585
R447 B.n663 B.n662 585
R448 B.n54 B.n53 585
R449 B.n661 B.n54 585
R450 B.n659 B.n658 585
R451 B.n660 B.n659 585
R452 B.n657 B.n59 585
R453 B.n59 B.n58 585
R454 B.n656 B.n655 585
R455 B.n655 B.n654 585
R456 B.n61 B.n60 585
R457 B.n653 B.n61 585
R458 B.n651 B.n650 585
R459 B.n652 B.n651 585
R460 B.n649 B.n66 585
R461 B.n66 B.n65 585
R462 B.n648 B.n647 585
R463 B.n647 B.n646 585
R464 B.n68 B.n67 585
R465 B.n645 B.n68 585
R466 B.n643 B.n642 585
R467 B.n644 B.n643 585
R468 B.n720 B.n719 585
R469 B.n718 B.n2 585
R470 B.n643 B.n73 473.281
R471 B.n514 B.n71 473.281
R472 B.n350 B.n182 473.281
R473 B.n348 B.n184 473.281
R474 B.n88 B.t8 263.813
R475 B.n95 B.t12 263.813
R476 B.n205 B.t4 263.813
R477 B.n199 B.t15 263.813
R478 B.n515 B.n72 256.663
R479 B.n517 B.n72 256.663
R480 B.n523 B.n72 256.663
R481 B.n525 B.n72 256.663
R482 B.n531 B.n72 256.663
R483 B.n533 B.n72 256.663
R484 B.n539 B.n72 256.663
R485 B.n541 B.n72 256.663
R486 B.n547 B.n72 256.663
R487 B.n549 B.n72 256.663
R488 B.n555 B.n72 256.663
R489 B.n557 B.n72 256.663
R490 B.n563 B.n72 256.663
R491 B.n565 B.n72 256.663
R492 B.n572 B.n72 256.663
R493 B.n574 B.n72 256.663
R494 B.n580 B.n72 256.663
R495 B.n582 B.n72 256.663
R496 B.n588 B.n72 256.663
R497 B.n590 B.n72 256.663
R498 B.n596 B.n72 256.663
R499 B.n598 B.n72 256.663
R500 B.n604 B.n72 256.663
R501 B.n606 B.n72 256.663
R502 B.n612 B.n72 256.663
R503 B.n614 B.n72 256.663
R504 B.n620 B.n72 256.663
R505 B.n622 B.n72 256.663
R506 B.n628 B.n72 256.663
R507 B.n630 B.n72 256.663
R508 B.n636 B.n72 256.663
R509 B.n638 B.n72 256.663
R510 B.n343 B.n183 256.663
R511 B.n186 B.n183 256.663
R512 B.n336 B.n183 256.663
R513 B.n330 B.n183 256.663
R514 B.n328 B.n183 256.663
R515 B.n322 B.n183 256.663
R516 B.n320 B.n183 256.663
R517 B.n314 B.n183 256.663
R518 B.n312 B.n183 256.663
R519 B.n306 B.n183 256.663
R520 B.n304 B.n183 256.663
R521 B.n298 B.n183 256.663
R522 B.n296 B.n183 256.663
R523 B.n289 B.n183 256.663
R524 B.n287 B.n183 256.663
R525 B.n281 B.n183 256.663
R526 B.n279 B.n183 256.663
R527 B.n273 B.n183 256.663
R528 B.n208 B.n183 256.663
R529 B.n267 B.n183 256.663
R530 B.n261 B.n183 256.663
R531 B.n259 B.n183 256.663
R532 B.n253 B.n183 256.663
R533 B.n251 B.n183 256.663
R534 B.n245 B.n183 256.663
R535 B.n243 B.n183 256.663
R536 B.n237 B.n183 256.663
R537 B.n235 B.n183 256.663
R538 B.n229 B.n183 256.663
R539 B.n227 B.n183 256.663
R540 B.n221 B.n183 256.663
R541 B.n722 B.n721 256.663
R542 B.n639 B.n637 163.367
R543 B.n635 B.n75 163.367
R544 B.n631 B.n629 163.367
R545 B.n627 B.n77 163.367
R546 B.n623 B.n621 163.367
R547 B.n619 B.n79 163.367
R548 B.n615 B.n613 163.367
R549 B.n611 B.n81 163.367
R550 B.n607 B.n605 163.367
R551 B.n603 B.n83 163.367
R552 B.n599 B.n597 163.367
R553 B.n595 B.n85 163.367
R554 B.n591 B.n589 163.367
R555 B.n587 B.n87 163.367
R556 B.n583 B.n581 163.367
R557 B.n579 B.n92 163.367
R558 B.n575 B.n573 163.367
R559 B.n571 B.n94 163.367
R560 B.n566 B.n564 163.367
R561 B.n562 B.n98 163.367
R562 B.n558 B.n556 163.367
R563 B.n554 B.n100 163.367
R564 B.n550 B.n548 163.367
R565 B.n546 B.n102 163.367
R566 B.n542 B.n540 163.367
R567 B.n538 B.n104 163.367
R568 B.n534 B.n532 163.367
R569 B.n530 B.n106 163.367
R570 B.n526 B.n524 163.367
R571 B.n522 B.n108 163.367
R572 B.n518 B.n516 163.367
R573 B.n350 B.n180 163.367
R574 B.n354 B.n180 163.367
R575 B.n354 B.n174 163.367
R576 B.n362 B.n174 163.367
R577 B.n362 B.n172 163.367
R578 B.n366 B.n172 163.367
R579 B.n366 B.n166 163.367
R580 B.n374 B.n166 163.367
R581 B.n374 B.n164 163.367
R582 B.n378 B.n164 163.367
R583 B.n378 B.n158 163.367
R584 B.n386 B.n158 163.367
R585 B.n386 B.n156 163.367
R586 B.n390 B.n156 163.367
R587 B.n390 B.n150 163.367
R588 B.n398 B.n150 163.367
R589 B.n398 B.n148 163.367
R590 B.n402 B.n148 163.367
R591 B.n402 B.n141 163.367
R592 B.n410 B.n141 163.367
R593 B.n410 B.n139 163.367
R594 B.n414 B.n139 163.367
R595 B.n414 B.n134 163.367
R596 B.n422 B.n134 163.367
R597 B.n422 B.n132 163.367
R598 B.n426 B.n132 163.367
R599 B.n426 B.n126 163.367
R600 B.n434 B.n126 163.367
R601 B.n434 B.n124 163.367
R602 B.n438 B.n124 163.367
R603 B.n438 B.n119 163.367
R604 B.n447 B.n119 163.367
R605 B.n447 B.n117 163.367
R606 B.n452 B.n117 163.367
R607 B.n452 B.n111 163.367
R608 B.n460 B.n111 163.367
R609 B.n461 B.n460 163.367
R610 B.n461 B.n5 163.367
R611 B.n6 B.n5 163.367
R612 B.n7 B.n6 163.367
R613 B.n467 B.n7 163.367
R614 B.n468 B.n467 163.367
R615 B.n468 B.n13 163.367
R616 B.n14 B.n13 163.367
R617 B.n15 B.n14 163.367
R618 B.n473 B.n15 163.367
R619 B.n473 B.n20 163.367
R620 B.n21 B.n20 163.367
R621 B.n22 B.n21 163.367
R622 B.n478 B.n22 163.367
R623 B.n478 B.n27 163.367
R624 B.n28 B.n27 163.367
R625 B.n29 B.n28 163.367
R626 B.n483 B.n29 163.367
R627 B.n483 B.n34 163.367
R628 B.n35 B.n34 163.367
R629 B.n36 B.n35 163.367
R630 B.n488 B.n36 163.367
R631 B.n488 B.n41 163.367
R632 B.n42 B.n41 163.367
R633 B.n43 B.n42 163.367
R634 B.n493 B.n43 163.367
R635 B.n493 B.n48 163.367
R636 B.n49 B.n48 163.367
R637 B.n50 B.n49 163.367
R638 B.n498 B.n50 163.367
R639 B.n498 B.n55 163.367
R640 B.n56 B.n55 163.367
R641 B.n57 B.n56 163.367
R642 B.n503 B.n57 163.367
R643 B.n503 B.n62 163.367
R644 B.n63 B.n62 163.367
R645 B.n64 B.n63 163.367
R646 B.n508 B.n64 163.367
R647 B.n508 B.n69 163.367
R648 B.n70 B.n69 163.367
R649 B.n71 B.n70 163.367
R650 B.n344 B.n342 163.367
R651 B.n342 B.n341 163.367
R652 B.n338 B.n337 163.367
R653 B.n335 B.n188 163.367
R654 B.n331 B.n329 163.367
R655 B.n327 B.n190 163.367
R656 B.n323 B.n321 163.367
R657 B.n319 B.n192 163.367
R658 B.n315 B.n313 163.367
R659 B.n311 B.n194 163.367
R660 B.n307 B.n305 163.367
R661 B.n303 B.n196 163.367
R662 B.n299 B.n297 163.367
R663 B.n295 B.n198 163.367
R664 B.n290 B.n288 163.367
R665 B.n286 B.n202 163.367
R666 B.n282 B.n280 163.367
R667 B.n278 B.n204 163.367
R668 B.n274 B.n272 163.367
R669 B.n269 B.n268 163.367
R670 B.n266 B.n210 163.367
R671 B.n262 B.n260 163.367
R672 B.n258 B.n212 163.367
R673 B.n254 B.n252 163.367
R674 B.n250 B.n214 163.367
R675 B.n246 B.n244 163.367
R676 B.n242 B.n216 163.367
R677 B.n238 B.n236 163.367
R678 B.n234 B.n218 163.367
R679 B.n230 B.n228 163.367
R680 B.n226 B.n220 163.367
R681 B.n222 B.n182 163.367
R682 B.n348 B.n178 163.367
R683 B.n356 B.n178 163.367
R684 B.n356 B.n176 163.367
R685 B.n360 B.n176 163.367
R686 B.n360 B.n170 163.367
R687 B.n368 B.n170 163.367
R688 B.n368 B.n168 163.367
R689 B.n372 B.n168 163.367
R690 B.n372 B.n162 163.367
R691 B.n380 B.n162 163.367
R692 B.n380 B.n160 163.367
R693 B.n384 B.n160 163.367
R694 B.n384 B.n154 163.367
R695 B.n392 B.n154 163.367
R696 B.n392 B.n152 163.367
R697 B.n396 B.n152 163.367
R698 B.n396 B.n146 163.367
R699 B.n404 B.n146 163.367
R700 B.n404 B.n144 163.367
R701 B.n408 B.n144 163.367
R702 B.n408 B.n138 163.367
R703 B.n416 B.n138 163.367
R704 B.n416 B.n136 163.367
R705 B.n420 B.n136 163.367
R706 B.n420 B.n130 163.367
R707 B.n428 B.n130 163.367
R708 B.n428 B.n128 163.367
R709 B.n432 B.n128 163.367
R710 B.n432 B.n122 163.367
R711 B.n441 B.n122 163.367
R712 B.n441 B.n120 163.367
R713 B.n445 B.n120 163.367
R714 B.n445 B.n115 163.367
R715 B.n454 B.n115 163.367
R716 B.n454 B.n113 163.367
R717 B.n458 B.n113 163.367
R718 B.n458 B.n3 163.367
R719 B.n720 B.n3 163.367
R720 B.n716 B.n2 163.367
R721 B.n716 B.n715 163.367
R722 B.n715 B.n9 163.367
R723 B.n711 B.n9 163.367
R724 B.n711 B.n11 163.367
R725 B.n707 B.n11 163.367
R726 B.n707 B.n16 163.367
R727 B.n703 B.n16 163.367
R728 B.n703 B.n18 163.367
R729 B.n699 B.n18 163.367
R730 B.n699 B.n24 163.367
R731 B.n695 B.n24 163.367
R732 B.n695 B.n26 163.367
R733 B.n691 B.n26 163.367
R734 B.n691 B.n31 163.367
R735 B.n687 B.n31 163.367
R736 B.n687 B.n33 163.367
R737 B.n683 B.n33 163.367
R738 B.n683 B.n38 163.367
R739 B.n679 B.n38 163.367
R740 B.n679 B.n40 163.367
R741 B.n675 B.n40 163.367
R742 B.n675 B.n45 163.367
R743 B.n671 B.n45 163.367
R744 B.n671 B.n47 163.367
R745 B.n667 B.n47 163.367
R746 B.n667 B.n52 163.367
R747 B.n663 B.n52 163.367
R748 B.n663 B.n54 163.367
R749 B.n659 B.n54 163.367
R750 B.n659 B.n59 163.367
R751 B.n655 B.n59 163.367
R752 B.n655 B.n61 163.367
R753 B.n651 B.n61 163.367
R754 B.n651 B.n66 163.367
R755 B.n647 B.n66 163.367
R756 B.n647 B.n68 163.367
R757 B.n643 B.n68 163.367
R758 B.n95 B.t13 141.075
R759 B.n205 B.t7 141.075
R760 B.n88 B.t10 141.066
R761 B.n199 B.t17 141.066
R762 B.n349 B.n183 102.305
R763 B.n644 B.n72 102.305
R764 B.n96 B.t14 74.5534
R765 B.n206 B.t6 74.5534
R766 B.n89 B.t11 74.5456
R767 B.n200 B.t16 74.5456
R768 B.n638 B.n73 71.676
R769 B.n637 B.n636 71.676
R770 B.n630 B.n75 71.676
R771 B.n629 B.n628 71.676
R772 B.n622 B.n77 71.676
R773 B.n621 B.n620 71.676
R774 B.n614 B.n79 71.676
R775 B.n613 B.n612 71.676
R776 B.n606 B.n81 71.676
R777 B.n605 B.n604 71.676
R778 B.n598 B.n83 71.676
R779 B.n597 B.n596 71.676
R780 B.n590 B.n85 71.676
R781 B.n589 B.n588 71.676
R782 B.n582 B.n87 71.676
R783 B.n581 B.n580 71.676
R784 B.n574 B.n92 71.676
R785 B.n573 B.n572 71.676
R786 B.n565 B.n94 71.676
R787 B.n564 B.n563 71.676
R788 B.n557 B.n98 71.676
R789 B.n556 B.n555 71.676
R790 B.n549 B.n100 71.676
R791 B.n548 B.n547 71.676
R792 B.n541 B.n102 71.676
R793 B.n540 B.n539 71.676
R794 B.n533 B.n104 71.676
R795 B.n532 B.n531 71.676
R796 B.n525 B.n106 71.676
R797 B.n524 B.n523 71.676
R798 B.n517 B.n108 71.676
R799 B.n516 B.n515 71.676
R800 B.n515 B.n514 71.676
R801 B.n518 B.n517 71.676
R802 B.n523 B.n522 71.676
R803 B.n526 B.n525 71.676
R804 B.n531 B.n530 71.676
R805 B.n534 B.n533 71.676
R806 B.n539 B.n538 71.676
R807 B.n542 B.n541 71.676
R808 B.n547 B.n546 71.676
R809 B.n550 B.n549 71.676
R810 B.n555 B.n554 71.676
R811 B.n558 B.n557 71.676
R812 B.n563 B.n562 71.676
R813 B.n566 B.n565 71.676
R814 B.n572 B.n571 71.676
R815 B.n575 B.n574 71.676
R816 B.n580 B.n579 71.676
R817 B.n583 B.n582 71.676
R818 B.n588 B.n587 71.676
R819 B.n591 B.n590 71.676
R820 B.n596 B.n595 71.676
R821 B.n599 B.n598 71.676
R822 B.n604 B.n603 71.676
R823 B.n607 B.n606 71.676
R824 B.n612 B.n611 71.676
R825 B.n615 B.n614 71.676
R826 B.n620 B.n619 71.676
R827 B.n623 B.n622 71.676
R828 B.n628 B.n627 71.676
R829 B.n631 B.n630 71.676
R830 B.n636 B.n635 71.676
R831 B.n639 B.n638 71.676
R832 B.n343 B.n184 71.676
R833 B.n341 B.n186 71.676
R834 B.n337 B.n336 71.676
R835 B.n330 B.n188 71.676
R836 B.n329 B.n328 71.676
R837 B.n322 B.n190 71.676
R838 B.n321 B.n320 71.676
R839 B.n314 B.n192 71.676
R840 B.n313 B.n312 71.676
R841 B.n306 B.n194 71.676
R842 B.n305 B.n304 71.676
R843 B.n298 B.n196 71.676
R844 B.n297 B.n296 71.676
R845 B.n289 B.n198 71.676
R846 B.n288 B.n287 71.676
R847 B.n281 B.n202 71.676
R848 B.n280 B.n279 71.676
R849 B.n273 B.n204 71.676
R850 B.n272 B.n208 71.676
R851 B.n268 B.n267 71.676
R852 B.n261 B.n210 71.676
R853 B.n260 B.n259 71.676
R854 B.n253 B.n212 71.676
R855 B.n252 B.n251 71.676
R856 B.n245 B.n214 71.676
R857 B.n244 B.n243 71.676
R858 B.n237 B.n216 71.676
R859 B.n236 B.n235 71.676
R860 B.n229 B.n218 71.676
R861 B.n228 B.n227 71.676
R862 B.n221 B.n220 71.676
R863 B.n344 B.n343 71.676
R864 B.n338 B.n186 71.676
R865 B.n336 B.n335 71.676
R866 B.n331 B.n330 71.676
R867 B.n328 B.n327 71.676
R868 B.n323 B.n322 71.676
R869 B.n320 B.n319 71.676
R870 B.n315 B.n314 71.676
R871 B.n312 B.n311 71.676
R872 B.n307 B.n306 71.676
R873 B.n304 B.n303 71.676
R874 B.n299 B.n298 71.676
R875 B.n296 B.n295 71.676
R876 B.n290 B.n289 71.676
R877 B.n287 B.n286 71.676
R878 B.n282 B.n281 71.676
R879 B.n279 B.n278 71.676
R880 B.n274 B.n273 71.676
R881 B.n269 B.n208 71.676
R882 B.n267 B.n266 71.676
R883 B.n262 B.n261 71.676
R884 B.n259 B.n258 71.676
R885 B.n254 B.n253 71.676
R886 B.n251 B.n250 71.676
R887 B.n246 B.n245 71.676
R888 B.n243 B.n242 71.676
R889 B.n238 B.n237 71.676
R890 B.n235 B.n234 71.676
R891 B.n230 B.n229 71.676
R892 B.n227 B.n226 71.676
R893 B.n222 B.n221 71.676
R894 B.n721 B.n720 71.676
R895 B.n721 B.n2 71.676
R896 B.n89 B.n88 66.5217
R897 B.n96 B.n95 66.5217
R898 B.n206 B.n205 66.5217
R899 B.n200 B.n199 66.5217
R900 B.n349 B.n179 60.4938
R901 B.n355 B.n179 60.4938
R902 B.n355 B.n175 60.4938
R903 B.n361 B.n175 60.4938
R904 B.n361 B.n171 60.4938
R905 B.n367 B.n171 60.4938
R906 B.n367 B.n167 60.4938
R907 B.n373 B.n167 60.4938
R908 B.n379 B.n163 60.4938
R909 B.n379 B.n159 60.4938
R910 B.n385 B.n159 60.4938
R911 B.n385 B.n155 60.4938
R912 B.n391 B.n155 60.4938
R913 B.n391 B.n151 60.4938
R914 B.n397 B.n151 60.4938
R915 B.n397 B.n147 60.4938
R916 B.n403 B.n147 60.4938
R917 B.n403 B.n142 60.4938
R918 B.n409 B.n142 60.4938
R919 B.n409 B.n143 60.4938
R920 B.n415 B.n135 60.4938
R921 B.n421 B.n135 60.4938
R922 B.n421 B.n131 60.4938
R923 B.n427 B.n131 60.4938
R924 B.n427 B.n127 60.4938
R925 B.n433 B.n127 60.4938
R926 B.n433 B.n123 60.4938
R927 B.n440 B.n123 60.4938
R928 B.n440 B.n439 60.4938
R929 B.n446 B.n116 60.4938
R930 B.n453 B.n116 60.4938
R931 B.n453 B.n112 60.4938
R932 B.n459 B.n112 60.4938
R933 B.n459 B.n4 60.4938
R934 B.n719 B.n4 60.4938
R935 B.n719 B.n718 60.4938
R936 B.n718 B.n717 60.4938
R937 B.n717 B.n8 60.4938
R938 B.n12 B.n8 60.4938
R939 B.n710 B.n12 60.4938
R940 B.n710 B.n709 60.4938
R941 B.n709 B.n708 60.4938
R942 B.n702 B.n19 60.4938
R943 B.n702 B.n701 60.4938
R944 B.n701 B.n700 60.4938
R945 B.n700 B.n23 60.4938
R946 B.n694 B.n23 60.4938
R947 B.n694 B.n693 60.4938
R948 B.n693 B.n692 60.4938
R949 B.n692 B.n30 60.4938
R950 B.n686 B.n30 60.4938
R951 B.n685 B.n684 60.4938
R952 B.n684 B.n37 60.4938
R953 B.n678 B.n37 60.4938
R954 B.n678 B.n677 60.4938
R955 B.n677 B.n676 60.4938
R956 B.n676 B.n44 60.4938
R957 B.n670 B.n44 60.4938
R958 B.n670 B.n669 60.4938
R959 B.n669 B.n668 60.4938
R960 B.n668 B.n51 60.4938
R961 B.n662 B.n51 60.4938
R962 B.n662 B.n661 60.4938
R963 B.n660 B.n58 60.4938
R964 B.n654 B.n58 60.4938
R965 B.n654 B.n653 60.4938
R966 B.n653 B.n652 60.4938
R967 B.n652 B.n65 60.4938
R968 B.n646 B.n65 60.4938
R969 B.n646 B.n645 60.4938
R970 B.n645 B.n644 60.4938
R971 B.n90 B.n89 59.5399
R972 B.n568 B.n96 59.5399
R973 B.n207 B.n206 59.5399
R974 B.n293 B.n200 59.5399
R975 B.n439 B.t3 51.5978
R976 B.n19 B.t2 51.5978
R977 B.n143 B.t1 46.2601
R978 B.t0 B.n685 46.2601
R979 B.t5 B.n163 32.0264
R980 B.n661 B.t9 32.0264
R981 B.n347 B.n346 30.7517
R982 B.n351 B.n181 30.7517
R983 B.n513 B.n512 30.7517
R984 B.n642 B.n641 30.7517
R985 B.n373 B.t5 28.4679
R986 B.t9 B.n660 28.4679
R987 B B.n722 18.0485
R988 B.n415 B.t1 14.2342
R989 B.n686 B.t0 14.2342
R990 B.n347 B.n177 10.6151
R991 B.n357 B.n177 10.6151
R992 B.n358 B.n357 10.6151
R993 B.n359 B.n358 10.6151
R994 B.n359 B.n169 10.6151
R995 B.n369 B.n169 10.6151
R996 B.n370 B.n369 10.6151
R997 B.n371 B.n370 10.6151
R998 B.n371 B.n161 10.6151
R999 B.n381 B.n161 10.6151
R1000 B.n382 B.n381 10.6151
R1001 B.n383 B.n382 10.6151
R1002 B.n383 B.n153 10.6151
R1003 B.n393 B.n153 10.6151
R1004 B.n394 B.n393 10.6151
R1005 B.n395 B.n394 10.6151
R1006 B.n395 B.n145 10.6151
R1007 B.n405 B.n145 10.6151
R1008 B.n406 B.n405 10.6151
R1009 B.n407 B.n406 10.6151
R1010 B.n407 B.n137 10.6151
R1011 B.n417 B.n137 10.6151
R1012 B.n418 B.n417 10.6151
R1013 B.n419 B.n418 10.6151
R1014 B.n419 B.n129 10.6151
R1015 B.n429 B.n129 10.6151
R1016 B.n430 B.n429 10.6151
R1017 B.n431 B.n430 10.6151
R1018 B.n431 B.n121 10.6151
R1019 B.n442 B.n121 10.6151
R1020 B.n443 B.n442 10.6151
R1021 B.n444 B.n443 10.6151
R1022 B.n444 B.n114 10.6151
R1023 B.n455 B.n114 10.6151
R1024 B.n456 B.n455 10.6151
R1025 B.n457 B.n456 10.6151
R1026 B.n457 B.n0 10.6151
R1027 B.n346 B.n345 10.6151
R1028 B.n345 B.n185 10.6151
R1029 B.n340 B.n185 10.6151
R1030 B.n340 B.n339 10.6151
R1031 B.n339 B.n187 10.6151
R1032 B.n334 B.n187 10.6151
R1033 B.n334 B.n333 10.6151
R1034 B.n333 B.n332 10.6151
R1035 B.n332 B.n189 10.6151
R1036 B.n326 B.n189 10.6151
R1037 B.n326 B.n325 10.6151
R1038 B.n325 B.n324 10.6151
R1039 B.n324 B.n191 10.6151
R1040 B.n318 B.n191 10.6151
R1041 B.n318 B.n317 10.6151
R1042 B.n317 B.n316 10.6151
R1043 B.n316 B.n193 10.6151
R1044 B.n310 B.n193 10.6151
R1045 B.n310 B.n309 10.6151
R1046 B.n309 B.n308 10.6151
R1047 B.n308 B.n195 10.6151
R1048 B.n302 B.n195 10.6151
R1049 B.n302 B.n301 10.6151
R1050 B.n301 B.n300 10.6151
R1051 B.n300 B.n197 10.6151
R1052 B.n294 B.n197 10.6151
R1053 B.n292 B.n291 10.6151
R1054 B.n291 B.n201 10.6151
R1055 B.n285 B.n201 10.6151
R1056 B.n285 B.n284 10.6151
R1057 B.n284 B.n283 10.6151
R1058 B.n283 B.n203 10.6151
R1059 B.n277 B.n203 10.6151
R1060 B.n277 B.n276 10.6151
R1061 B.n276 B.n275 10.6151
R1062 B.n271 B.n270 10.6151
R1063 B.n270 B.n209 10.6151
R1064 B.n265 B.n209 10.6151
R1065 B.n265 B.n264 10.6151
R1066 B.n264 B.n263 10.6151
R1067 B.n263 B.n211 10.6151
R1068 B.n257 B.n211 10.6151
R1069 B.n257 B.n256 10.6151
R1070 B.n256 B.n255 10.6151
R1071 B.n255 B.n213 10.6151
R1072 B.n249 B.n213 10.6151
R1073 B.n249 B.n248 10.6151
R1074 B.n248 B.n247 10.6151
R1075 B.n247 B.n215 10.6151
R1076 B.n241 B.n215 10.6151
R1077 B.n241 B.n240 10.6151
R1078 B.n240 B.n239 10.6151
R1079 B.n239 B.n217 10.6151
R1080 B.n233 B.n217 10.6151
R1081 B.n233 B.n232 10.6151
R1082 B.n232 B.n231 10.6151
R1083 B.n231 B.n219 10.6151
R1084 B.n225 B.n219 10.6151
R1085 B.n225 B.n224 10.6151
R1086 B.n224 B.n223 10.6151
R1087 B.n223 B.n181 10.6151
R1088 B.n352 B.n351 10.6151
R1089 B.n353 B.n352 10.6151
R1090 B.n353 B.n173 10.6151
R1091 B.n363 B.n173 10.6151
R1092 B.n364 B.n363 10.6151
R1093 B.n365 B.n364 10.6151
R1094 B.n365 B.n165 10.6151
R1095 B.n375 B.n165 10.6151
R1096 B.n376 B.n375 10.6151
R1097 B.n377 B.n376 10.6151
R1098 B.n377 B.n157 10.6151
R1099 B.n387 B.n157 10.6151
R1100 B.n388 B.n387 10.6151
R1101 B.n389 B.n388 10.6151
R1102 B.n389 B.n149 10.6151
R1103 B.n399 B.n149 10.6151
R1104 B.n400 B.n399 10.6151
R1105 B.n401 B.n400 10.6151
R1106 B.n401 B.n140 10.6151
R1107 B.n411 B.n140 10.6151
R1108 B.n412 B.n411 10.6151
R1109 B.n413 B.n412 10.6151
R1110 B.n413 B.n133 10.6151
R1111 B.n423 B.n133 10.6151
R1112 B.n424 B.n423 10.6151
R1113 B.n425 B.n424 10.6151
R1114 B.n425 B.n125 10.6151
R1115 B.n435 B.n125 10.6151
R1116 B.n436 B.n435 10.6151
R1117 B.n437 B.n436 10.6151
R1118 B.n437 B.n118 10.6151
R1119 B.n448 B.n118 10.6151
R1120 B.n449 B.n448 10.6151
R1121 B.n451 B.n449 10.6151
R1122 B.n451 B.n450 10.6151
R1123 B.n450 B.n110 10.6151
R1124 B.n462 B.n110 10.6151
R1125 B.n463 B.n462 10.6151
R1126 B.n464 B.n463 10.6151
R1127 B.n465 B.n464 10.6151
R1128 B.n466 B.n465 10.6151
R1129 B.n469 B.n466 10.6151
R1130 B.n470 B.n469 10.6151
R1131 B.n471 B.n470 10.6151
R1132 B.n472 B.n471 10.6151
R1133 B.n474 B.n472 10.6151
R1134 B.n475 B.n474 10.6151
R1135 B.n476 B.n475 10.6151
R1136 B.n477 B.n476 10.6151
R1137 B.n479 B.n477 10.6151
R1138 B.n480 B.n479 10.6151
R1139 B.n481 B.n480 10.6151
R1140 B.n482 B.n481 10.6151
R1141 B.n484 B.n482 10.6151
R1142 B.n485 B.n484 10.6151
R1143 B.n486 B.n485 10.6151
R1144 B.n487 B.n486 10.6151
R1145 B.n489 B.n487 10.6151
R1146 B.n490 B.n489 10.6151
R1147 B.n491 B.n490 10.6151
R1148 B.n492 B.n491 10.6151
R1149 B.n494 B.n492 10.6151
R1150 B.n495 B.n494 10.6151
R1151 B.n496 B.n495 10.6151
R1152 B.n497 B.n496 10.6151
R1153 B.n499 B.n497 10.6151
R1154 B.n500 B.n499 10.6151
R1155 B.n501 B.n500 10.6151
R1156 B.n502 B.n501 10.6151
R1157 B.n504 B.n502 10.6151
R1158 B.n505 B.n504 10.6151
R1159 B.n506 B.n505 10.6151
R1160 B.n507 B.n506 10.6151
R1161 B.n509 B.n507 10.6151
R1162 B.n510 B.n509 10.6151
R1163 B.n511 B.n510 10.6151
R1164 B.n512 B.n511 10.6151
R1165 B.n714 B.n1 10.6151
R1166 B.n714 B.n713 10.6151
R1167 B.n713 B.n712 10.6151
R1168 B.n712 B.n10 10.6151
R1169 B.n706 B.n10 10.6151
R1170 B.n706 B.n705 10.6151
R1171 B.n705 B.n704 10.6151
R1172 B.n704 B.n17 10.6151
R1173 B.n698 B.n17 10.6151
R1174 B.n698 B.n697 10.6151
R1175 B.n697 B.n696 10.6151
R1176 B.n696 B.n25 10.6151
R1177 B.n690 B.n25 10.6151
R1178 B.n690 B.n689 10.6151
R1179 B.n689 B.n688 10.6151
R1180 B.n688 B.n32 10.6151
R1181 B.n682 B.n32 10.6151
R1182 B.n682 B.n681 10.6151
R1183 B.n681 B.n680 10.6151
R1184 B.n680 B.n39 10.6151
R1185 B.n674 B.n39 10.6151
R1186 B.n674 B.n673 10.6151
R1187 B.n673 B.n672 10.6151
R1188 B.n672 B.n46 10.6151
R1189 B.n666 B.n46 10.6151
R1190 B.n666 B.n665 10.6151
R1191 B.n665 B.n664 10.6151
R1192 B.n664 B.n53 10.6151
R1193 B.n658 B.n53 10.6151
R1194 B.n658 B.n657 10.6151
R1195 B.n657 B.n656 10.6151
R1196 B.n656 B.n60 10.6151
R1197 B.n650 B.n60 10.6151
R1198 B.n650 B.n649 10.6151
R1199 B.n649 B.n648 10.6151
R1200 B.n648 B.n67 10.6151
R1201 B.n642 B.n67 10.6151
R1202 B.n641 B.n640 10.6151
R1203 B.n640 B.n74 10.6151
R1204 B.n634 B.n74 10.6151
R1205 B.n634 B.n633 10.6151
R1206 B.n633 B.n632 10.6151
R1207 B.n632 B.n76 10.6151
R1208 B.n626 B.n76 10.6151
R1209 B.n626 B.n625 10.6151
R1210 B.n625 B.n624 10.6151
R1211 B.n624 B.n78 10.6151
R1212 B.n618 B.n78 10.6151
R1213 B.n618 B.n617 10.6151
R1214 B.n617 B.n616 10.6151
R1215 B.n616 B.n80 10.6151
R1216 B.n610 B.n80 10.6151
R1217 B.n610 B.n609 10.6151
R1218 B.n609 B.n608 10.6151
R1219 B.n608 B.n82 10.6151
R1220 B.n602 B.n82 10.6151
R1221 B.n602 B.n601 10.6151
R1222 B.n601 B.n600 10.6151
R1223 B.n600 B.n84 10.6151
R1224 B.n594 B.n84 10.6151
R1225 B.n594 B.n593 10.6151
R1226 B.n593 B.n592 10.6151
R1227 B.n592 B.n86 10.6151
R1228 B.n586 B.n585 10.6151
R1229 B.n585 B.n584 10.6151
R1230 B.n584 B.n91 10.6151
R1231 B.n578 B.n91 10.6151
R1232 B.n578 B.n577 10.6151
R1233 B.n577 B.n576 10.6151
R1234 B.n576 B.n93 10.6151
R1235 B.n570 B.n93 10.6151
R1236 B.n570 B.n569 10.6151
R1237 B.n567 B.n97 10.6151
R1238 B.n561 B.n97 10.6151
R1239 B.n561 B.n560 10.6151
R1240 B.n560 B.n559 10.6151
R1241 B.n559 B.n99 10.6151
R1242 B.n553 B.n99 10.6151
R1243 B.n553 B.n552 10.6151
R1244 B.n552 B.n551 10.6151
R1245 B.n551 B.n101 10.6151
R1246 B.n545 B.n101 10.6151
R1247 B.n545 B.n544 10.6151
R1248 B.n544 B.n543 10.6151
R1249 B.n543 B.n103 10.6151
R1250 B.n537 B.n103 10.6151
R1251 B.n537 B.n536 10.6151
R1252 B.n536 B.n535 10.6151
R1253 B.n535 B.n105 10.6151
R1254 B.n529 B.n105 10.6151
R1255 B.n529 B.n528 10.6151
R1256 B.n528 B.n527 10.6151
R1257 B.n527 B.n107 10.6151
R1258 B.n521 B.n107 10.6151
R1259 B.n521 B.n520 10.6151
R1260 B.n520 B.n519 10.6151
R1261 B.n519 B.n109 10.6151
R1262 B.n513 B.n109 10.6151
R1263 B.n294 B.n293 9.36635
R1264 B.n271 B.n207 9.36635
R1265 B.n90 B.n86 9.36635
R1266 B.n568 B.n567 9.36635
R1267 B.n446 B.t3 8.89658
R1268 B.n708 B.t2 8.89658
R1269 B.n722 B.n0 8.11757
R1270 B.n722 B.n1 8.11757
R1271 B.n293 B.n292 1.24928
R1272 B.n275 B.n207 1.24928
R1273 B.n586 B.n90 1.24928
R1274 B.n569 B.n568 1.24928
R1275 VP.n15 VP.n14 161.3
R1276 VP.n13 VP.n1 161.3
R1277 VP.n12 VP.n11 161.3
R1278 VP.n10 VP.n2 161.3
R1279 VP.n9 VP.n8 161.3
R1280 VP.n7 VP.n3 161.3
R1281 VP.n4 VP.t0 89.6301
R1282 VP.n4 VP.t3 88.6156
R1283 VP.n6 VP.n5 67.3131
R1284 VP.n16 VP.n0 67.3131
R1285 VP.n12 VP.n2 56.5193
R1286 VP.n6 VP.t2 55.1195
R1287 VP.n0 VP.t1 55.1195
R1288 VP.n5 VP.n4 47.0706
R1289 VP.n8 VP.n7 24.4675
R1290 VP.n8 VP.n2 24.4675
R1291 VP.n13 VP.n12 24.4675
R1292 VP.n14 VP.n13 24.4675
R1293 VP.n7 VP.n6 22.7548
R1294 VP.n14 VP.n0 22.7548
R1295 VP.n5 VP.n3 0.354971
R1296 VP.n16 VP.n15 0.354971
R1297 VP VP.n16 0.26696
R1298 VP.n9 VP.n3 0.189894
R1299 VP.n10 VP.n9 0.189894
R1300 VP.n11 VP.n10 0.189894
R1301 VP.n11 VP.n1 0.189894
R1302 VP.n15 VP.n1 0.189894
R1303 VDD1 VDD1.n1 105.028
R1304 VDD1 VDD1.n0 65.8632
R1305 VDD1.n0 VDD1.t3 2.79317
R1306 VDD1.n0 VDD1.t0 2.79317
R1307 VDD1.n1 VDD1.t1 2.79317
R1308 VDD1.n1 VDD1.t2 2.79317
C0 VN VDD2 3.01725f
C1 VDD2 VTAIL 4.4803f
C2 VP VDD1 3.29305f
C3 VP VN 5.64059f
C4 VP VTAIL 3.36969f
C5 VDD1 VN 0.149595f
C6 VDD1 VTAIL 4.42274f
C7 VN VTAIL 3.35558f
C8 VP VDD2 0.426265f
C9 VDD1 VDD2 1.14914f
C10 VDD2 B 3.675934f
C11 VDD1 B 7.547071f
C12 VTAIL B 7.113105f
C13 VN B 11.170219f
C14 VP B 9.535129f
C15 VDD1.t3 B 0.157162f
C16 VDD1.t0 B 0.157162f
C17 VDD1.n0 B 1.33623f
C18 VDD1.t1 B 0.157162f
C19 VDD1.t2 B 0.157162f
C20 VDD1.n1 B 1.89534f
C21 VP.t1 B 1.51439f
C22 VP.n0 B 0.663576f
C23 VP.n1 B 0.025799f
C24 VP.n2 B 0.037662f
C25 VP.n3 B 0.041639f
C26 VP.t2 B 1.51439f
C27 VP.t0 B 1.80138f
C28 VP.t3 B 1.79327f
C29 VP.n4 B 2.4639f
C30 VP.n5 B 1.32753f
C31 VP.n6 B 0.663576f
C32 VP.n7 B 0.04642f
C33 VP.n8 B 0.048083f
C34 VP.n9 B 0.025799f
C35 VP.n10 B 0.025799f
C36 VP.n11 B 0.025799f
C37 VP.n12 B 0.037662f
C38 VP.n13 B 0.048083f
C39 VP.n14 B 0.04642f
C40 VP.n15 B 0.041639f
C41 VP.n16 B 0.050993f
C42 VTAIL.t5 B 1.10699f
C43 VTAIL.n0 B 0.367657f
C44 VTAIL.t3 B 1.10699f
C45 VTAIL.n1 B 0.456173f
C46 VTAIL.t1 B 1.10699f
C47 VTAIL.n2 B 1.25484f
C48 VTAIL.t7 B 1.107f
C49 VTAIL.n3 B 1.25483f
C50 VTAIL.t6 B 1.107f
C51 VTAIL.n4 B 0.456168f
C52 VTAIL.t2 B 1.107f
C53 VTAIL.n5 B 0.456168f
C54 VTAIL.t0 B 1.10699f
C55 VTAIL.n6 B 1.25484f
C56 VTAIL.t4 B 1.10699f
C57 VTAIL.n7 B 1.15907f
C58 VDD2.t1 B 0.155168f
C59 VDD2.t0 B 0.155168f
C60 VDD2.n0 B 1.84614f
C61 VDD2.t3 B 0.155168f
C62 VDD2.t2 B 0.155168f
C63 VDD2.n1 B 1.31883f
C64 VDD2.n2 B 3.44453f
C65 VN.t3 B 1.74439f
C66 VN.t2 B 1.75228f
C67 VN.n0 B 1.05714f
C68 VN.t1 B 1.75228f
C69 VN.t0 B 1.74439f
C70 VN.n1 B 2.40713f
.ends

