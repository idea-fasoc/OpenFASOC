* NGSPICE file created from diff_pair_sample_1678.ext - technology: sky130A

.subckt diff_pair_sample_1678 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=2.57
X1 VDD1.t7 VP.t0 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=2.57
X2 VDD1.t6 VP.t1 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X3 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X4 VTAIL.t10 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X5 VDD1.t4 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=2.57
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=2.57
X7 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X8 VTAIL.t15 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X9 VTAIL.t11 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=2.57
X10 VDD2.t4 VN.t3 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X11 VTAIL.t9 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=2.57
X12 VTAIL.t2 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=2.57
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=2.57
X14 VTAIL.t0 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=2.57
X15 VDD2.t1 VN.t6 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=2.57
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=2.57
X17 VTAIL.t13 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X18 VDD1.t0 VP.t7 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=1.66155 ps=10.4 w=10.07 l=2.57
X19 VDD2.t0 VN.t7 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=2.57
R0 B.n660 B.n138 585
R1 B.n138 B.n93 585
R2 B.n662 B.n661 585
R3 B.n664 B.n137 585
R4 B.n667 B.n666 585
R5 B.n668 B.n136 585
R6 B.n670 B.n669 585
R7 B.n672 B.n135 585
R8 B.n675 B.n674 585
R9 B.n676 B.n134 585
R10 B.n678 B.n677 585
R11 B.n680 B.n133 585
R12 B.n683 B.n682 585
R13 B.n684 B.n132 585
R14 B.n686 B.n685 585
R15 B.n688 B.n131 585
R16 B.n691 B.n690 585
R17 B.n692 B.n130 585
R18 B.n694 B.n693 585
R19 B.n696 B.n129 585
R20 B.n699 B.n698 585
R21 B.n700 B.n128 585
R22 B.n702 B.n701 585
R23 B.n704 B.n127 585
R24 B.n707 B.n706 585
R25 B.n708 B.n126 585
R26 B.n710 B.n709 585
R27 B.n712 B.n125 585
R28 B.n715 B.n714 585
R29 B.n716 B.n124 585
R30 B.n718 B.n717 585
R31 B.n720 B.n123 585
R32 B.n723 B.n722 585
R33 B.n724 B.n122 585
R34 B.n726 B.n725 585
R35 B.n728 B.n121 585
R36 B.n731 B.n730 585
R37 B.n733 B.n118 585
R38 B.n735 B.n734 585
R39 B.n737 B.n117 585
R40 B.n740 B.n739 585
R41 B.n741 B.n116 585
R42 B.n743 B.n742 585
R43 B.n745 B.n115 585
R44 B.n748 B.n747 585
R45 B.n749 B.n112 585
R46 B.n752 B.n751 585
R47 B.n754 B.n111 585
R48 B.n757 B.n756 585
R49 B.n758 B.n110 585
R50 B.n760 B.n759 585
R51 B.n762 B.n109 585
R52 B.n765 B.n764 585
R53 B.n766 B.n108 585
R54 B.n768 B.n767 585
R55 B.n770 B.n107 585
R56 B.n773 B.n772 585
R57 B.n774 B.n106 585
R58 B.n776 B.n775 585
R59 B.n778 B.n105 585
R60 B.n781 B.n780 585
R61 B.n782 B.n104 585
R62 B.n784 B.n783 585
R63 B.n786 B.n103 585
R64 B.n789 B.n788 585
R65 B.n790 B.n102 585
R66 B.n792 B.n791 585
R67 B.n794 B.n101 585
R68 B.n797 B.n796 585
R69 B.n798 B.n100 585
R70 B.n800 B.n799 585
R71 B.n802 B.n99 585
R72 B.n805 B.n804 585
R73 B.n806 B.n98 585
R74 B.n808 B.n807 585
R75 B.n810 B.n97 585
R76 B.n813 B.n812 585
R77 B.n814 B.n96 585
R78 B.n816 B.n815 585
R79 B.n818 B.n95 585
R80 B.n821 B.n820 585
R81 B.n822 B.n94 585
R82 B.n659 B.n92 585
R83 B.n825 B.n92 585
R84 B.n658 B.n91 585
R85 B.n826 B.n91 585
R86 B.n657 B.n90 585
R87 B.n827 B.n90 585
R88 B.n656 B.n655 585
R89 B.n655 B.n86 585
R90 B.n654 B.n85 585
R91 B.n833 B.n85 585
R92 B.n653 B.n84 585
R93 B.n834 B.n84 585
R94 B.n652 B.n83 585
R95 B.n835 B.n83 585
R96 B.n651 B.n650 585
R97 B.n650 B.n82 585
R98 B.n649 B.n78 585
R99 B.n841 B.n78 585
R100 B.n648 B.n77 585
R101 B.n842 B.n77 585
R102 B.n647 B.n76 585
R103 B.n843 B.n76 585
R104 B.n646 B.n645 585
R105 B.n645 B.n72 585
R106 B.n644 B.n71 585
R107 B.n849 B.n71 585
R108 B.n643 B.n70 585
R109 B.n850 B.n70 585
R110 B.n642 B.n69 585
R111 B.n851 B.n69 585
R112 B.n641 B.n640 585
R113 B.n640 B.n65 585
R114 B.n639 B.n64 585
R115 B.n857 B.n64 585
R116 B.n638 B.n63 585
R117 B.n858 B.n63 585
R118 B.n637 B.n62 585
R119 B.n859 B.n62 585
R120 B.n636 B.n635 585
R121 B.n635 B.n61 585
R122 B.n634 B.n57 585
R123 B.n865 B.n57 585
R124 B.n633 B.n56 585
R125 B.n866 B.n56 585
R126 B.n632 B.n55 585
R127 B.n867 B.n55 585
R128 B.n631 B.n630 585
R129 B.n630 B.n51 585
R130 B.n629 B.n50 585
R131 B.n873 B.n50 585
R132 B.n628 B.n49 585
R133 B.n874 B.n49 585
R134 B.n627 B.n48 585
R135 B.n875 B.n48 585
R136 B.n626 B.n625 585
R137 B.n625 B.n47 585
R138 B.n624 B.n43 585
R139 B.n881 B.n43 585
R140 B.n623 B.n42 585
R141 B.n882 B.n42 585
R142 B.n622 B.n41 585
R143 B.n883 B.n41 585
R144 B.n621 B.n620 585
R145 B.n620 B.n37 585
R146 B.n619 B.n36 585
R147 B.n889 B.n36 585
R148 B.n618 B.n35 585
R149 B.n890 B.n35 585
R150 B.n617 B.n34 585
R151 B.n891 B.n34 585
R152 B.n616 B.n615 585
R153 B.n615 B.n30 585
R154 B.n614 B.n29 585
R155 B.n897 B.n29 585
R156 B.n613 B.n28 585
R157 B.n898 B.n28 585
R158 B.n612 B.n27 585
R159 B.n899 B.n27 585
R160 B.n611 B.n610 585
R161 B.n610 B.n23 585
R162 B.n609 B.n22 585
R163 B.n905 B.n22 585
R164 B.n608 B.n21 585
R165 B.n906 B.n21 585
R166 B.n607 B.n20 585
R167 B.n907 B.n20 585
R168 B.n606 B.n605 585
R169 B.n605 B.n16 585
R170 B.n604 B.n15 585
R171 B.n913 B.n15 585
R172 B.n603 B.n14 585
R173 B.n914 B.n14 585
R174 B.n602 B.n13 585
R175 B.n915 B.n13 585
R176 B.n601 B.n600 585
R177 B.n600 B.n12 585
R178 B.n599 B.n598 585
R179 B.n599 B.n8 585
R180 B.n597 B.n7 585
R181 B.n922 B.n7 585
R182 B.n596 B.n6 585
R183 B.n923 B.n6 585
R184 B.n595 B.n5 585
R185 B.n924 B.n5 585
R186 B.n594 B.n593 585
R187 B.n593 B.n4 585
R188 B.n592 B.n139 585
R189 B.n592 B.n591 585
R190 B.n582 B.n140 585
R191 B.n141 B.n140 585
R192 B.n584 B.n583 585
R193 B.n585 B.n584 585
R194 B.n581 B.n146 585
R195 B.n146 B.n145 585
R196 B.n580 B.n579 585
R197 B.n579 B.n578 585
R198 B.n148 B.n147 585
R199 B.n149 B.n148 585
R200 B.n571 B.n570 585
R201 B.n572 B.n571 585
R202 B.n569 B.n154 585
R203 B.n154 B.n153 585
R204 B.n568 B.n567 585
R205 B.n567 B.n566 585
R206 B.n156 B.n155 585
R207 B.n157 B.n156 585
R208 B.n559 B.n558 585
R209 B.n560 B.n559 585
R210 B.n557 B.n162 585
R211 B.n162 B.n161 585
R212 B.n556 B.n555 585
R213 B.n555 B.n554 585
R214 B.n164 B.n163 585
R215 B.n165 B.n164 585
R216 B.n547 B.n546 585
R217 B.n548 B.n547 585
R218 B.n545 B.n170 585
R219 B.n170 B.n169 585
R220 B.n544 B.n543 585
R221 B.n543 B.n542 585
R222 B.n172 B.n171 585
R223 B.n173 B.n172 585
R224 B.n535 B.n534 585
R225 B.n536 B.n535 585
R226 B.n533 B.n178 585
R227 B.n178 B.n177 585
R228 B.n532 B.n531 585
R229 B.n531 B.n530 585
R230 B.n180 B.n179 585
R231 B.n523 B.n180 585
R232 B.n522 B.n521 585
R233 B.n524 B.n522 585
R234 B.n520 B.n185 585
R235 B.n185 B.n184 585
R236 B.n519 B.n518 585
R237 B.n518 B.n517 585
R238 B.n187 B.n186 585
R239 B.n188 B.n187 585
R240 B.n510 B.n509 585
R241 B.n511 B.n510 585
R242 B.n508 B.n193 585
R243 B.n193 B.n192 585
R244 B.n507 B.n506 585
R245 B.n506 B.n505 585
R246 B.n195 B.n194 585
R247 B.n498 B.n195 585
R248 B.n497 B.n496 585
R249 B.n499 B.n497 585
R250 B.n495 B.n200 585
R251 B.n200 B.n199 585
R252 B.n494 B.n493 585
R253 B.n493 B.n492 585
R254 B.n202 B.n201 585
R255 B.n203 B.n202 585
R256 B.n485 B.n484 585
R257 B.n486 B.n485 585
R258 B.n483 B.n208 585
R259 B.n208 B.n207 585
R260 B.n482 B.n481 585
R261 B.n481 B.n480 585
R262 B.n210 B.n209 585
R263 B.n211 B.n210 585
R264 B.n473 B.n472 585
R265 B.n474 B.n473 585
R266 B.n471 B.n216 585
R267 B.n216 B.n215 585
R268 B.n470 B.n469 585
R269 B.n469 B.n468 585
R270 B.n218 B.n217 585
R271 B.n461 B.n218 585
R272 B.n460 B.n459 585
R273 B.n462 B.n460 585
R274 B.n458 B.n223 585
R275 B.n223 B.n222 585
R276 B.n457 B.n456 585
R277 B.n456 B.n455 585
R278 B.n225 B.n224 585
R279 B.n226 B.n225 585
R280 B.n448 B.n447 585
R281 B.n449 B.n448 585
R282 B.n446 B.n231 585
R283 B.n231 B.n230 585
R284 B.n445 B.n444 585
R285 B.n444 B.n443 585
R286 B.n440 B.n235 585
R287 B.n439 B.n438 585
R288 B.n436 B.n236 585
R289 B.n436 B.n234 585
R290 B.n435 B.n434 585
R291 B.n433 B.n432 585
R292 B.n431 B.n238 585
R293 B.n429 B.n428 585
R294 B.n427 B.n239 585
R295 B.n426 B.n425 585
R296 B.n423 B.n240 585
R297 B.n421 B.n420 585
R298 B.n419 B.n241 585
R299 B.n418 B.n417 585
R300 B.n415 B.n242 585
R301 B.n413 B.n412 585
R302 B.n411 B.n243 585
R303 B.n410 B.n409 585
R304 B.n407 B.n244 585
R305 B.n405 B.n404 585
R306 B.n403 B.n245 585
R307 B.n402 B.n401 585
R308 B.n399 B.n246 585
R309 B.n397 B.n396 585
R310 B.n395 B.n247 585
R311 B.n394 B.n393 585
R312 B.n391 B.n248 585
R313 B.n389 B.n388 585
R314 B.n387 B.n249 585
R315 B.n386 B.n385 585
R316 B.n383 B.n250 585
R317 B.n381 B.n380 585
R318 B.n379 B.n251 585
R319 B.n378 B.n377 585
R320 B.n375 B.n252 585
R321 B.n373 B.n372 585
R322 B.n371 B.n253 585
R323 B.n369 B.n368 585
R324 B.n366 B.n256 585
R325 B.n364 B.n363 585
R326 B.n362 B.n257 585
R327 B.n361 B.n360 585
R328 B.n358 B.n258 585
R329 B.n356 B.n355 585
R330 B.n354 B.n259 585
R331 B.n353 B.n352 585
R332 B.n350 B.n349 585
R333 B.n348 B.n347 585
R334 B.n346 B.n264 585
R335 B.n344 B.n343 585
R336 B.n342 B.n265 585
R337 B.n341 B.n340 585
R338 B.n338 B.n266 585
R339 B.n336 B.n335 585
R340 B.n334 B.n267 585
R341 B.n333 B.n332 585
R342 B.n330 B.n268 585
R343 B.n328 B.n327 585
R344 B.n326 B.n269 585
R345 B.n325 B.n324 585
R346 B.n322 B.n270 585
R347 B.n320 B.n319 585
R348 B.n318 B.n271 585
R349 B.n317 B.n316 585
R350 B.n314 B.n272 585
R351 B.n312 B.n311 585
R352 B.n310 B.n273 585
R353 B.n309 B.n308 585
R354 B.n306 B.n274 585
R355 B.n304 B.n303 585
R356 B.n302 B.n275 585
R357 B.n301 B.n300 585
R358 B.n298 B.n276 585
R359 B.n296 B.n295 585
R360 B.n294 B.n277 585
R361 B.n293 B.n292 585
R362 B.n290 B.n278 585
R363 B.n288 B.n287 585
R364 B.n286 B.n279 585
R365 B.n285 B.n284 585
R366 B.n282 B.n280 585
R367 B.n233 B.n232 585
R368 B.n442 B.n441 585
R369 B.n443 B.n442 585
R370 B.n229 B.n228 585
R371 B.n230 B.n229 585
R372 B.n451 B.n450 585
R373 B.n450 B.n449 585
R374 B.n452 B.n227 585
R375 B.n227 B.n226 585
R376 B.n454 B.n453 585
R377 B.n455 B.n454 585
R378 B.n221 B.n220 585
R379 B.n222 B.n221 585
R380 B.n464 B.n463 585
R381 B.n463 B.n462 585
R382 B.n465 B.n219 585
R383 B.n461 B.n219 585
R384 B.n467 B.n466 585
R385 B.n468 B.n467 585
R386 B.n214 B.n213 585
R387 B.n215 B.n214 585
R388 B.n476 B.n475 585
R389 B.n475 B.n474 585
R390 B.n477 B.n212 585
R391 B.n212 B.n211 585
R392 B.n479 B.n478 585
R393 B.n480 B.n479 585
R394 B.n206 B.n205 585
R395 B.n207 B.n206 585
R396 B.n488 B.n487 585
R397 B.n487 B.n486 585
R398 B.n489 B.n204 585
R399 B.n204 B.n203 585
R400 B.n491 B.n490 585
R401 B.n492 B.n491 585
R402 B.n198 B.n197 585
R403 B.n199 B.n198 585
R404 B.n501 B.n500 585
R405 B.n500 B.n499 585
R406 B.n502 B.n196 585
R407 B.n498 B.n196 585
R408 B.n504 B.n503 585
R409 B.n505 B.n504 585
R410 B.n191 B.n190 585
R411 B.n192 B.n191 585
R412 B.n513 B.n512 585
R413 B.n512 B.n511 585
R414 B.n514 B.n189 585
R415 B.n189 B.n188 585
R416 B.n516 B.n515 585
R417 B.n517 B.n516 585
R418 B.n183 B.n182 585
R419 B.n184 B.n183 585
R420 B.n526 B.n525 585
R421 B.n525 B.n524 585
R422 B.n527 B.n181 585
R423 B.n523 B.n181 585
R424 B.n529 B.n528 585
R425 B.n530 B.n529 585
R426 B.n176 B.n175 585
R427 B.n177 B.n176 585
R428 B.n538 B.n537 585
R429 B.n537 B.n536 585
R430 B.n539 B.n174 585
R431 B.n174 B.n173 585
R432 B.n541 B.n540 585
R433 B.n542 B.n541 585
R434 B.n168 B.n167 585
R435 B.n169 B.n168 585
R436 B.n550 B.n549 585
R437 B.n549 B.n548 585
R438 B.n551 B.n166 585
R439 B.n166 B.n165 585
R440 B.n553 B.n552 585
R441 B.n554 B.n553 585
R442 B.n160 B.n159 585
R443 B.n161 B.n160 585
R444 B.n562 B.n561 585
R445 B.n561 B.n560 585
R446 B.n563 B.n158 585
R447 B.n158 B.n157 585
R448 B.n565 B.n564 585
R449 B.n566 B.n565 585
R450 B.n152 B.n151 585
R451 B.n153 B.n152 585
R452 B.n574 B.n573 585
R453 B.n573 B.n572 585
R454 B.n575 B.n150 585
R455 B.n150 B.n149 585
R456 B.n577 B.n576 585
R457 B.n578 B.n577 585
R458 B.n144 B.n143 585
R459 B.n145 B.n144 585
R460 B.n587 B.n586 585
R461 B.n586 B.n585 585
R462 B.n588 B.n142 585
R463 B.n142 B.n141 585
R464 B.n590 B.n589 585
R465 B.n591 B.n590 585
R466 B.n3 B.n0 585
R467 B.n4 B.n3 585
R468 B.n921 B.n1 585
R469 B.n922 B.n921 585
R470 B.n920 B.n919 585
R471 B.n920 B.n8 585
R472 B.n918 B.n9 585
R473 B.n12 B.n9 585
R474 B.n917 B.n916 585
R475 B.n916 B.n915 585
R476 B.n11 B.n10 585
R477 B.n914 B.n11 585
R478 B.n912 B.n911 585
R479 B.n913 B.n912 585
R480 B.n910 B.n17 585
R481 B.n17 B.n16 585
R482 B.n909 B.n908 585
R483 B.n908 B.n907 585
R484 B.n19 B.n18 585
R485 B.n906 B.n19 585
R486 B.n904 B.n903 585
R487 B.n905 B.n904 585
R488 B.n902 B.n24 585
R489 B.n24 B.n23 585
R490 B.n901 B.n900 585
R491 B.n900 B.n899 585
R492 B.n26 B.n25 585
R493 B.n898 B.n26 585
R494 B.n896 B.n895 585
R495 B.n897 B.n896 585
R496 B.n894 B.n31 585
R497 B.n31 B.n30 585
R498 B.n893 B.n892 585
R499 B.n892 B.n891 585
R500 B.n33 B.n32 585
R501 B.n890 B.n33 585
R502 B.n888 B.n887 585
R503 B.n889 B.n888 585
R504 B.n886 B.n38 585
R505 B.n38 B.n37 585
R506 B.n885 B.n884 585
R507 B.n884 B.n883 585
R508 B.n40 B.n39 585
R509 B.n882 B.n40 585
R510 B.n880 B.n879 585
R511 B.n881 B.n880 585
R512 B.n878 B.n44 585
R513 B.n47 B.n44 585
R514 B.n877 B.n876 585
R515 B.n876 B.n875 585
R516 B.n46 B.n45 585
R517 B.n874 B.n46 585
R518 B.n872 B.n871 585
R519 B.n873 B.n872 585
R520 B.n870 B.n52 585
R521 B.n52 B.n51 585
R522 B.n869 B.n868 585
R523 B.n868 B.n867 585
R524 B.n54 B.n53 585
R525 B.n866 B.n54 585
R526 B.n864 B.n863 585
R527 B.n865 B.n864 585
R528 B.n862 B.n58 585
R529 B.n61 B.n58 585
R530 B.n861 B.n860 585
R531 B.n860 B.n859 585
R532 B.n60 B.n59 585
R533 B.n858 B.n60 585
R534 B.n856 B.n855 585
R535 B.n857 B.n856 585
R536 B.n854 B.n66 585
R537 B.n66 B.n65 585
R538 B.n853 B.n852 585
R539 B.n852 B.n851 585
R540 B.n68 B.n67 585
R541 B.n850 B.n68 585
R542 B.n848 B.n847 585
R543 B.n849 B.n848 585
R544 B.n846 B.n73 585
R545 B.n73 B.n72 585
R546 B.n845 B.n844 585
R547 B.n844 B.n843 585
R548 B.n75 B.n74 585
R549 B.n842 B.n75 585
R550 B.n840 B.n839 585
R551 B.n841 B.n840 585
R552 B.n838 B.n79 585
R553 B.n82 B.n79 585
R554 B.n837 B.n836 585
R555 B.n836 B.n835 585
R556 B.n81 B.n80 585
R557 B.n834 B.n81 585
R558 B.n832 B.n831 585
R559 B.n833 B.n832 585
R560 B.n830 B.n87 585
R561 B.n87 B.n86 585
R562 B.n829 B.n828 585
R563 B.n828 B.n827 585
R564 B.n89 B.n88 585
R565 B.n826 B.n89 585
R566 B.n824 B.n823 585
R567 B.n825 B.n824 585
R568 B.n925 B.n924 585
R569 B.n923 B.n2 585
R570 B.n824 B.n94 578.989
R571 B.n138 B.n92 578.989
R572 B.n444 B.n233 578.989
R573 B.n442 B.n235 578.989
R574 B.n119 B.t10 305.248
R575 B.n260 B.t18 305.248
R576 B.n113 B.t20 305.248
R577 B.n254 B.t15 305.248
R578 B.n113 B.t19 302.433
R579 B.n119 B.t8 302.433
R580 B.n260 B.t16 302.433
R581 B.n254 B.t12 302.433
R582 B.n663 B.n93 256.663
R583 B.n665 B.n93 256.663
R584 B.n671 B.n93 256.663
R585 B.n673 B.n93 256.663
R586 B.n679 B.n93 256.663
R587 B.n681 B.n93 256.663
R588 B.n687 B.n93 256.663
R589 B.n689 B.n93 256.663
R590 B.n695 B.n93 256.663
R591 B.n697 B.n93 256.663
R592 B.n703 B.n93 256.663
R593 B.n705 B.n93 256.663
R594 B.n711 B.n93 256.663
R595 B.n713 B.n93 256.663
R596 B.n719 B.n93 256.663
R597 B.n721 B.n93 256.663
R598 B.n727 B.n93 256.663
R599 B.n729 B.n93 256.663
R600 B.n736 B.n93 256.663
R601 B.n738 B.n93 256.663
R602 B.n744 B.n93 256.663
R603 B.n746 B.n93 256.663
R604 B.n753 B.n93 256.663
R605 B.n755 B.n93 256.663
R606 B.n761 B.n93 256.663
R607 B.n763 B.n93 256.663
R608 B.n769 B.n93 256.663
R609 B.n771 B.n93 256.663
R610 B.n777 B.n93 256.663
R611 B.n779 B.n93 256.663
R612 B.n785 B.n93 256.663
R613 B.n787 B.n93 256.663
R614 B.n793 B.n93 256.663
R615 B.n795 B.n93 256.663
R616 B.n801 B.n93 256.663
R617 B.n803 B.n93 256.663
R618 B.n809 B.n93 256.663
R619 B.n811 B.n93 256.663
R620 B.n817 B.n93 256.663
R621 B.n819 B.n93 256.663
R622 B.n437 B.n234 256.663
R623 B.n237 B.n234 256.663
R624 B.n430 B.n234 256.663
R625 B.n424 B.n234 256.663
R626 B.n422 B.n234 256.663
R627 B.n416 B.n234 256.663
R628 B.n414 B.n234 256.663
R629 B.n408 B.n234 256.663
R630 B.n406 B.n234 256.663
R631 B.n400 B.n234 256.663
R632 B.n398 B.n234 256.663
R633 B.n392 B.n234 256.663
R634 B.n390 B.n234 256.663
R635 B.n384 B.n234 256.663
R636 B.n382 B.n234 256.663
R637 B.n376 B.n234 256.663
R638 B.n374 B.n234 256.663
R639 B.n367 B.n234 256.663
R640 B.n365 B.n234 256.663
R641 B.n359 B.n234 256.663
R642 B.n357 B.n234 256.663
R643 B.n351 B.n234 256.663
R644 B.n263 B.n234 256.663
R645 B.n345 B.n234 256.663
R646 B.n339 B.n234 256.663
R647 B.n337 B.n234 256.663
R648 B.n331 B.n234 256.663
R649 B.n329 B.n234 256.663
R650 B.n323 B.n234 256.663
R651 B.n321 B.n234 256.663
R652 B.n315 B.n234 256.663
R653 B.n313 B.n234 256.663
R654 B.n307 B.n234 256.663
R655 B.n305 B.n234 256.663
R656 B.n299 B.n234 256.663
R657 B.n297 B.n234 256.663
R658 B.n291 B.n234 256.663
R659 B.n289 B.n234 256.663
R660 B.n283 B.n234 256.663
R661 B.n281 B.n234 256.663
R662 B.n927 B.n926 256.663
R663 B.n120 B.t11 249.005
R664 B.n261 B.t17 249.005
R665 B.n114 B.t21 249.005
R666 B.n255 B.t14 249.005
R667 B.n820 B.n818 163.367
R668 B.n816 B.n96 163.367
R669 B.n812 B.n810 163.367
R670 B.n808 B.n98 163.367
R671 B.n804 B.n802 163.367
R672 B.n800 B.n100 163.367
R673 B.n796 B.n794 163.367
R674 B.n792 B.n102 163.367
R675 B.n788 B.n786 163.367
R676 B.n784 B.n104 163.367
R677 B.n780 B.n778 163.367
R678 B.n776 B.n106 163.367
R679 B.n772 B.n770 163.367
R680 B.n768 B.n108 163.367
R681 B.n764 B.n762 163.367
R682 B.n760 B.n110 163.367
R683 B.n756 B.n754 163.367
R684 B.n752 B.n112 163.367
R685 B.n747 B.n745 163.367
R686 B.n743 B.n116 163.367
R687 B.n739 B.n737 163.367
R688 B.n735 B.n118 163.367
R689 B.n730 B.n728 163.367
R690 B.n726 B.n122 163.367
R691 B.n722 B.n720 163.367
R692 B.n718 B.n124 163.367
R693 B.n714 B.n712 163.367
R694 B.n710 B.n126 163.367
R695 B.n706 B.n704 163.367
R696 B.n702 B.n128 163.367
R697 B.n698 B.n696 163.367
R698 B.n694 B.n130 163.367
R699 B.n690 B.n688 163.367
R700 B.n686 B.n132 163.367
R701 B.n682 B.n680 163.367
R702 B.n678 B.n134 163.367
R703 B.n674 B.n672 163.367
R704 B.n670 B.n136 163.367
R705 B.n666 B.n664 163.367
R706 B.n662 B.n138 163.367
R707 B.n444 B.n231 163.367
R708 B.n448 B.n231 163.367
R709 B.n448 B.n225 163.367
R710 B.n456 B.n225 163.367
R711 B.n456 B.n223 163.367
R712 B.n460 B.n223 163.367
R713 B.n460 B.n218 163.367
R714 B.n469 B.n218 163.367
R715 B.n469 B.n216 163.367
R716 B.n473 B.n216 163.367
R717 B.n473 B.n210 163.367
R718 B.n481 B.n210 163.367
R719 B.n481 B.n208 163.367
R720 B.n485 B.n208 163.367
R721 B.n485 B.n202 163.367
R722 B.n493 B.n202 163.367
R723 B.n493 B.n200 163.367
R724 B.n497 B.n200 163.367
R725 B.n497 B.n195 163.367
R726 B.n506 B.n195 163.367
R727 B.n506 B.n193 163.367
R728 B.n510 B.n193 163.367
R729 B.n510 B.n187 163.367
R730 B.n518 B.n187 163.367
R731 B.n518 B.n185 163.367
R732 B.n522 B.n185 163.367
R733 B.n522 B.n180 163.367
R734 B.n531 B.n180 163.367
R735 B.n531 B.n178 163.367
R736 B.n535 B.n178 163.367
R737 B.n535 B.n172 163.367
R738 B.n543 B.n172 163.367
R739 B.n543 B.n170 163.367
R740 B.n547 B.n170 163.367
R741 B.n547 B.n164 163.367
R742 B.n555 B.n164 163.367
R743 B.n555 B.n162 163.367
R744 B.n559 B.n162 163.367
R745 B.n559 B.n156 163.367
R746 B.n567 B.n156 163.367
R747 B.n567 B.n154 163.367
R748 B.n571 B.n154 163.367
R749 B.n571 B.n148 163.367
R750 B.n579 B.n148 163.367
R751 B.n579 B.n146 163.367
R752 B.n584 B.n146 163.367
R753 B.n584 B.n140 163.367
R754 B.n592 B.n140 163.367
R755 B.n593 B.n592 163.367
R756 B.n593 B.n5 163.367
R757 B.n6 B.n5 163.367
R758 B.n7 B.n6 163.367
R759 B.n599 B.n7 163.367
R760 B.n600 B.n599 163.367
R761 B.n600 B.n13 163.367
R762 B.n14 B.n13 163.367
R763 B.n15 B.n14 163.367
R764 B.n605 B.n15 163.367
R765 B.n605 B.n20 163.367
R766 B.n21 B.n20 163.367
R767 B.n22 B.n21 163.367
R768 B.n610 B.n22 163.367
R769 B.n610 B.n27 163.367
R770 B.n28 B.n27 163.367
R771 B.n29 B.n28 163.367
R772 B.n615 B.n29 163.367
R773 B.n615 B.n34 163.367
R774 B.n35 B.n34 163.367
R775 B.n36 B.n35 163.367
R776 B.n620 B.n36 163.367
R777 B.n620 B.n41 163.367
R778 B.n42 B.n41 163.367
R779 B.n43 B.n42 163.367
R780 B.n625 B.n43 163.367
R781 B.n625 B.n48 163.367
R782 B.n49 B.n48 163.367
R783 B.n50 B.n49 163.367
R784 B.n630 B.n50 163.367
R785 B.n630 B.n55 163.367
R786 B.n56 B.n55 163.367
R787 B.n57 B.n56 163.367
R788 B.n635 B.n57 163.367
R789 B.n635 B.n62 163.367
R790 B.n63 B.n62 163.367
R791 B.n64 B.n63 163.367
R792 B.n640 B.n64 163.367
R793 B.n640 B.n69 163.367
R794 B.n70 B.n69 163.367
R795 B.n71 B.n70 163.367
R796 B.n645 B.n71 163.367
R797 B.n645 B.n76 163.367
R798 B.n77 B.n76 163.367
R799 B.n78 B.n77 163.367
R800 B.n650 B.n78 163.367
R801 B.n650 B.n83 163.367
R802 B.n84 B.n83 163.367
R803 B.n85 B.n84 163.367
R804 B.n655 B.n85 163.367
R805 B.n655 B.n90 163.367
R806 B.n91 B.n90 163.367
R807 B.n92 B.n91 163.367
R808 B.n438 B.n436 163.367
R809 B.n436 B.n435 163.367
R810 B.n432 B.n431 163.367
R811 B.n429 B.n239 163.367
R812 B.n425 B.n423 163.367
R813 B.n421 B.n241 163.367
R814 B.n417 B.n415 163.367
R815 B.n413 B.n243 163.367
R816 B.n409 B.n407 163.367
R817 B.n405 B.n245 163.367
R818 B.n401 B.n399 163.367
R819 B.n397 B.n247 163.367
R820 B.n393 B.n391 163.367
R821 B.n389 B.n249 163.367
R822 B.n385 B.n383 163.367
R823 B.n381 B.n251 163.367
R824 B.n377 B.n375 163.367
R825 B.n373 B.n253 163.367
R826 B.n368 B.n366 163.367
R827 B.n364 B.n257 163.367
R828 B.n360 B.n358 163.367
R829 B.n356 B.n259 163.367
R830 B.n352 B.n350 163.367
R831 B.n347 B.n346 163.367
R832 B.n344 B.n265 163.367
R833 B.n340 B.n338 163.367
R834 B.n336 B.n267 163.367
R835 B.n332 B.n330 163.367
R836 B.n328 B.n269 163.367
R837 B.n324 B.n322 163.367
R838 B.n320 B.n271 163.367
R839 B.n316 B.n314 163.367
R840 B.n312 B.n273 163.367
R841 B.n308 B.n306 163.367
R842 B.n304 B.n275 163.367
R843 B.n300 B.n298 163.367
R844 B.n296 B.n277 163.367
R845 B.n292 B.n290 163.367
R846 B.n288 B.n279 163.367
R847 B.n284 B.n282 163.367
R848 B.n442 B.n229 163.367
R849 B.n450 B.n229 163.367
R850 B.n450 B.n227 163.367
R851 B.n454 B.n227 163.367
R852 B.n454 B.n221 163.367
R853 B.n463 B.n221 163.367
R854 B.n463 B.n219 163.367
R855 B.n467 B.n219 163.367
R856 B.n467 B.n214 163.367
R857 B.n475 B.n214 163.367
R858 B.n475 B.n212 163.367
R859 B.n479 B.n212 163.367
R860 B.n479 B.n206 163.367
R861 B.n487 B.n206 163.367
R862 B.n487 B.n204 163.367
R863 B.n491 B.n204 163.367
R864 B.n491 B.n198 163.367
R865 B.n500 B.n198 163.367
R866 B.n500 B.n196 163.367
R867 B.n504 B.n196 163.367
R868 B.n504 B.n191 163.367
R869 B.n512 B.n191 163.367
R870 B.n512 B.n189 163.367
R871 B.n516 B.n189 163.367
R872 B.n516 B.n183 163.367
R873 B.n525 B.n183 163.367
R874 B.n525 B.n181 163.367
R875 B.n529 B.n181 163.367
R876 B.n529 B.n176 163.367
R877 B.n537 B.n176 163.367
R878 B.n537 B.n174 163.367
R879 B.n541 B.n174 163.367
R880 B.n541 B.n168 163.367
R881 B.n549 B.n168 163.367
R882 B.n549 B.n166 163.367
R883 B.n553 B.n166 163.367
R884 B.n553 B.n160 163.367
R885 B.n561 B.n160 163.367
R886 B.n561 B.n158 163.367
R887 B.n565 B.n158 163.367
R888 B.n565 B.n152 163.367
R889 B.n573 B.n152 163.367
R890 B.n573 B.n150 163.367
R891 B.n577 B.n150 163.367
R892 B.n577 B.n144 163.367
R893 B.n586 B.n144 163.367
R894 B.n586 B.n142 163.367
R895 B.n590 B.n142 163.367
R896 B.n590 B.n3 163.367
R897 B.n925 B.n3 163.367
R898 B.n921 B.n2 163.367
R899 B.n921 B.n920 163.367
R900 B.n920 B.n9 163.367
R901 B.n916 B.n9 163.367
R902 B.n916 B.n11 163.367
R903 B.n912 B.n11 163.367
R904 B.n912 B.n17 163.367
R905 B.n908 B.n17 163.367
R906 B.n908 B.n19 163.367
R907 B.n904 B.n19 163.367
R908 B.n904 B.n24 163.367
R909 B.n900 B.n24 163.367
R910 B.n900 B.n26 163.367
R911 B.n896 B.n26 163.367
R912 B.n896 B.n31 163.367
R913 B.n892 B.n31 163.367
R914 B.n892 B.n33 163.367
R915 B.n888 B.n33 163.367
R916 B.n888 B.n38 163.367
R917 B.n884 B.n38 163.367
R918 B.n884 B.n40 163.367
R919 B.n880 B.n40 163.367
R920 B.n880 B.n44 163.367
R921 B.n876 B.n44 163.367
R922 B.n876 B.n46 163.367
R923 B.n872 B.n46 163.367
R924 B.n872 B.n52 163.367
R925 B.n868 B.n52 163.367
R926 B.n868 B.n54 163.367
R927 B.n864 B.n54 163.367
R928 B.n864 B.n58 163.367
R929 B.n860 B.n58 163.367
R930 B.n860 B.n60 163.367
R931 B.n856 B.n60 163.367
R932 B.n856 B.n66 163.367
R933 B.n852 B.n66 163.367
R934 B.n852 B.n68 163.367
R935 B.n848 B.n68 163.367
R936 B.n848 B.n73 163.367
R937 B.n844 B.n73 163.367
R938 B.n844 B.n75 163.367
R939 B.n840 B.n75 163.367
R940 B.n840 B.n79 163.367
R941 B.n836 B.n79 163.367
R942 B.n836 B.n81 163.367
R943 B.n832 B.n81 163.367
R944 B.n832 B.n87 163.367
R945 B.n828 B.n87 163.367
R946 B.n828 B.n89 163.367
R947 B.n824 B.n89 163.367
R948 B.n443 B.n234 101.076
R949 B.n825 B.n93 101.076
R950 B.n819 B.n94 71.676
R951 B.n818 B.n817 71.676
R952 B.n811 B.n96 71.676
R953 B.n810 B.n809 71.676
R954 B.n803 B.n98 71.676
R955 B.n802 B.n801 71.676
R956 B.n795 B.n100 71.676
R957 B.n794 B.n793 71.676
R958 B.n787 B.n102 71.676
R959 B.n786 B.n785 71.676
R960 B.n779 B.n104 71.676
R961 B.n778 B.n777 71.676
R962 B.n771 B.n106 71.676
R963 B.n770 B.n769 71.676
R964 B.n763 B.n108 71.676
R965 B.n762 B.n761 71.676
R966 B.n755 B.n110 71.676
R967 B.n754 B.n753 71.676
R968 B.n746 B.n112 71.676
R969 B.n745 B.n744 71.676
R970 B.n738 B.n116 71.676
R971 B.n737 B.n736 71.676
R972 B.n729 B.n118 71.676
R973 B.n728 B.n727 71.676
R974 B.n721 B.n122 71.676
R975 B.n720 B.n719 71.676
R976 B.n713 B.n124 71.676
R977 B.n712 B.n711 71.676
R978 B.n705 B.n126 71.676
R979 B.n704 B.n703 71.676
R980 B.n697 B.n128 71.676
R981 B.n696 B.n695 71.676
R982 B.n689 B.n130 71.676
R983 B.n688 B.n687 71.676
R984 B.n681 B.n132 71.676
R985 B.n680 B.n679 71.676
R986 B.n673 B.n134 71.676
R987 B.n672 B.n671 71.676
R988 B.n665 B.n136 71.676
R989 B.n664 B.n663 71.676
R990 B.n663 B.n662 71.676
R991 B.n666 B.n665 71.676
R992 B.n671 B.n670 71.676
R993 B.n674 B.n673 71.676
R994 B.n679 B.n678 71.676
R995 B.n682 B.n681 71.676
R996 B.n687 B.n686 71.676
R997 B.n690 B.n689 71.676
R998 B.n695 B.n694 71.676
R999 B.n698 B.n697 71.676
R1000 B.n703 B.n702 71.676
R1001 B.n706 B.n705 71.676
R1002 B.n711 B.n710 71.676
R1003 B.n714 B.n713 71.676
R1004 B.n719 B.n718 71.676
R1005 B.n722 B.n721 71.676
R1006 B.n727 B.n726 71.676
R1007 B.n730 B.n729 71.676
R1008 B.n736 B.n735 71.676
R1009 B.n739 B.n738 71.676
R1010 B.n744 B.n743 71.676
R1011 B.n747 B.n746 71.676
R1012 B.n753 B.n752 71.676
R1013 B.n756 B.n755 71.676
R1014 B.n761 B.n760 71.676
R1015 B.n764 B.n763 71.676
R1016 B.n769 B.n768 71.676
R1017 B.n772 B.n771 71.676
R1018 B.n777 B.n776 71.676
R1019 B.n780 B.n779 71.676
R1020 B.n785 B.n784 71.676
R1021 B.n788 B.n787 71.676
R1022 B.n793 B.n792 71.676
R1023 B.n796 B.n795 71.676
R1024 B.n801 B.n800 71.676
R1025 B.n804 B.n803 71.676
R1026 B.n809 B.n808 71.676
R1027 B.n812 B.n811 71.676
R1028 B.n817 B.n816 71.676
R1029 B.n820 B.n819 71.676
R1030 B.n437 B.n235 71.676
R1031 B.n435 B.n237 71.676
R1032 B.n431 B.n430 71.676
R1033 B.n424 B.n239 71.676
R1034 B.n423 B.n422 71.676
R1035 B.n416 B.n241 71.676
R1036 B.n415 B.n414 71.676
R1037 B.n408 B.n243 71.676
R1038 B.n407 B.n406 71.676
R1039 B.n400 B.n245 71.676
R1040 B.n399 B.n398 71.676
R1041 B.n392 B.n247 71.676
R1042 B.n391 B.n390 71.676
R1043 B.n384 B.n249 71.676
R1044 B.n383 B.n382 71.676
R1045 B.n376 B.n251 71.676
R1046 B.n375 B.n374 71.676
R1047 B.n367 B.n253 71.676
R1048 B.n366 B.n365 71.676
R1049 B.n359 B.n257 71.676
R1050 B.n358 B.n357 71.676
R1051 B.n351 B.n259 71.676
R1052 B.n350 B.n263 71.676
R1053 B.n346 B.n345 71.676
R1054 B.n339 B.n265 71.676
R1055 B.n338 B.n337 71.676
R1056 B.n331 B.n267 71.676
R1057 B.n330 B.n329 71.676
R1058 B.n323 B.n269 71.676
R1059 B.n322 B.n321 71.676
R1060 B.n315 B.n271 71.676
R1061 B.n314 B.n313 71.676
R1062 B.n307 B.n273 71.676
R1063 B.n306 B.n305 71.676
R1064 B.n299 B.n275 71.676
R1065 B.n298 B.n297 71.676
R1066 B.n291 B.n277 71.676
R1067 B.n290 B.n289 71.676
R1068 B.n283 B.n279 71.676
R1069 B.n282 B.n281 71.676
R1070 B.n438 B.n437 71.676
R1071 B.n432 B.n237 71.676
R1072 B.n430 B.n429 71.676
R1073 B.n425 B.n424 71.676
R1074 B.n422 B.n421 71.676
R1075 B.n417 B.n416 71.676
R1076 B.n414 B.n413 71.676
R1077 B.n409 B.n408 71.676
R1078 B.n406 B.n405 71.676
R1079 B.n401 B.n400 71.676
R1080 B.n398 B.n397 71.676
R1081 B.n393 B.n392 71.676
R1082 B.n390 B.n389 71.676
R1083 B.n385 B.n384 71.676
R1084 B.n382 B.n381 71.676
R1085 B.n377 B.n376 71.676
R1086 B.n374 B.n373 71.676
R1087 B.n368 B.n367 71.676
R1088 B.n365 B.n364 71.676
R1089 B.n360 B.n359 71.676
R1090 B.n357 B.n356 71.676
R1091 B.n352 B.n351 71.676
R1092 B.n347 B.n263 71.676
R1093 B.n345 B.n344 71.676
R1094 B.n340 B.n339 71.676
R1095 B.n337 B.n336 71.676
R1096 B.n332 B.n331 71.676
R1097 B.n329 B.n328 71.676
R1098 B.n324 B.n323 71.676
R1099 B.n321 B.n320 71.676
R1100 B.n316 B.n315 71.676
R1101 B.n313 B.n312 71.676
R1102 B.n308 B.n307 71.676
R1103 B.n305 B.n304 71.676
R1104 B.n300 B.n299 71.676
R1105 B.n297 B.n296 71.676
R1106 B.n292 B.n291 71.676
R1107 B.n289 B.n288 71.676
R1108 B.n284 B.n283 71.676
R1109 B.n281 B.n233 71.676
R1110 B.n926 B.n925 71.676
R1111 B.n926 B.n2 71.676
R1112 B.n750 B.n114 59.5399
R1113 B.n732 B.n120 59.5399
R1114 B.n262 B.n261 59.5399
R1115 B.n370 B.n255 59.5399
R1116 B.n114 B.n113 56.2429
R1117 B.n120 B.n119 56.2429
R1118 B.n261 B.n260 56.2429
R1119 B.n255 B.n254 56.2429
R1120 B.n443 B.n230 48.746
R1121 B.n449 B.n230 48.746
R1122 B.n449 B.n226 48.746
R1123 B.n455 B.n226 48.746
R1124 B.n455 B.n222 48.746
R1125 B.n462 B.n222 48.746
R1126 B.n462 B.n461 48.746
R1127 B.n468 B.n215 48.746
R1128 B.n474 B.n215 48.746
R1129 B.n474 B.n211 48.746
R1130 B.n480 B.n211 48.746
R1131 B.n480 B.n207 48.746
R1132 B.n486 B.n207 48.746
R1133 B.n486 B.n203 48.746
R1134 B.n492 B.n203 48.746
R1135 B.n492 B.n199 48.746
R1136 B.n499 B.n199 48.746
R1137 B.n499 B.n498 48.746
R1138 B.n505 B.n192 48.746
R1139 B.n511 B.n192 48.746
R1140 B.n511 B.n188 48.746
R1141 B.n517 B.n188 48.746
R1142 B.n517 B.n184 48.746
R1143 B.n524 B.n184 48.746
R1144 B.n524 B.n523 48.746
R1145 B.n530 B.n177 48.746
R1146 B.n536 B.n177 48.746
R1147 B.n536 B.n173 48.746
R1148 B.n542 B.n173 48.746
R1149 B.n542 B.n169 48.746
R1150 B.n548 B.n169 48.746
R1151 B.n548 B.n165 48.746
R1152 B.n554 B.n165 48.746
R1153 B.n560 B.n161 48.746
R1154 B.n560 B.n157 48.746
R1155 B.n566 B.n157 48.746
R1156 B.n566 B.n153 48.746
R1157 B.n572 B.n153 48.746
R1158 B.n572 B.n149 48.746
R1159 B.n578 B.n149 48.746
R1160 B.n585 B.n145 48.746
R1161 B.n585 B.n141 48.746
R1162 B.n591 B.n141 48.746
R1163 B.n591 B.n4 48.746
R1164 B.n924 B.n4 48.746
R1165 B.n924 B.n923 48.746
R1166 B.n923 B.n922 48.746
R1167 B.n922 B.n8 48.746
R1168 B.n12 B.n8 48.746
R1169 B.n915 B.n12 48.746
R1170 B.n915 B.n914 48.746
R1171 B.n913 B.n16 48.746
R1172 B.n907 B.n16 48.746
R1173 B.n907 B.n906 48.746
R1174 B.n906 B.n905 48.746
R1175 B.n905 B.n23 48.746
R1176 B.n899 B.n23 48.746
R1177 B.n899 B.n898 48.746
R1178 B.n897 B.n30 48.746
R1179 B.n891 B.n30 48.746
R1180 B.n891 B.n890 48.746
R1181 B.n890 B.n889 48.746
R1182 B.n889 B.n37 48.746
R1183 B.n883 B.n37 48.746
R1184 B.n883 B.n882 48.746
R1185 B.n882 B.n881 48.746
R1186 B.n875 B.n47 48.746
R1187 B.n875 B.n874 48.746
R1188 B.n874 B.n873 48.746
R1189 B.n873 B.n51 48.746
R1190 B.n867 B.n51 48.746
R1191 B.n867 B.n866 48.746
R1192 B.n866 B.n865 48.746
R1193 B.n859 B.n61 48.746
R1194 B.n859 B.n858 48.746
R1195 B.n858 B.n857 48.746
R1196 B.n857 B.n65 48.746
R1197 B.n851 B.n65 48.746
R1198 B.n851 B.n850 48.746
R1199 B.n850 B.n849 48.746
R1200 B.n849 B.n72 48.746
R1201 B.n843 B.n72 48.746
R1202 B.n843 B.n842 48.746
R1203 B.n842 B.n841 48.746
R1204 B.n835 B.n82 48.746
R1205 B.n835 B.n834 48.746
R1206 B.n834 B.n833 48.746
R1207 B.n833 B.n86 48.746
R1208 B.n827 B.n86 48.746
R1209 B.n827 B.n826 48.746
R1210 B.n826 B.n825 48.746
R1211 B.n505 B.t3 46.5955
R1212 B.n865 B.t4 46.5955
R1213 B.t5 B.n161 43.7281
R1214 B.n898 B.t2 43.7281
R1215 B.n441 B.n440 37.62
R1216 B.n445 B.n232 37.62
R1217 B.n660 B.n659 37.62
R1218 B.n823 B.n822 37.62
R1219 B.n468 B.t13 33.6923
R1220 B.n841 B.t9 33.6923
R1221 B.n578 B.t0 30.8249
R1222 B.t1 B.n913 30.8249
R1223 B.n523 B.t6 27.9575
R1224 B.n47 B.t7 27.9575
R1225 B.n530 B.t6 20.789
R1226 B.n881 B.t7 20.789
R1227 B B.n927 18.0485
R1228 B.t0 B.n145 17.9216
R1229 B.n914 B.t1 17.9216
R1230 B.n461 B.t13 15.0543
R1231 B.n82 B.t9 15.0543
R1232 B.n441 B.n228 10.6151
R1233 B.n451 B.n228 10.6151
R1234 B.n452 B.n451 10.6151
R1235 B.n453 B.n452 10.6151
R1236 B.n453 B.n220 10.6151
R1237 B.n464 B.n220 10.6151
R1238 B.n465 B.n464 10.6151
R1239 B.n466 B.n465 10.6151
R1240 B.n466 B.n213 10.6151
R1241 B.n476 B.n213 10.6151
R1242 B.n477 B.n476 10.6151
R1243 B.n478 B.n477 10.6151
R1244 B.n478 B.n205 10.6151
R1245 B.n488 B.n205 10.6151
R1246 B.n489 B.n488 10.6151
R1247 B.n490 B.n489 10.6151
R1248 B.n490 B.n197 10.6151
R1249 B.n501 B.n197 10.6151
R1250 B.n502 B.n501 10.6151
R1251 B.n503 B.n502 10.6151
R1252 B.n503 B.n190 10.6151
R1253 B.n513 B.n190 10.6151
R1254 B.n514 B.n513 10.6151
R1255 B.n515 B.n514 10.6151
R1256 B.n515 B.n182 10.6151
R1257 B.n526 B.n182 10.6151
R1258 B.n527 B.n526 10.6151
R1259 B.n528 B.n527 10.6151
R1260 B.n528 B.n175 10.6151
R1261 B.n538 B.n175 10.6151
R1262 B.n539 B.n538 10.6151
R1263 B.n540 B.n539 10.6151
R1264 B.n540 B.n167 10.6151
R1265 B.n550 B.n167 10.6151
R1266 B.n551 B.n550 10.6151
R1267 B.n552 B.n551 10.6151
R1268 B.n552 B.n159 10.6151
R1269 B.n562 B.n159 10.6151
R1270 B.n563 B.n562 10.6151
R1271 B.n564 B.n563 10.6151
R1272 B.n564 B.n151 10.6151
R1273 B.n574 B.n151 10.6151
R1274 B.n575 B.n574 10.6151
R1275 B.n576 B.n575 10.6151
R1276 B.n576 B.n143 10.6151
R1277 B.n587 B.n143 10.6151
R1278 B.n588 B.n587 10.6151
R1279 B.n589 B.n588 10.6151
R1280 B.n589 B.n0 10.6151
R1281 B.n440 B.n439 10.6151
R1282 B.n439 B.n236 10.6151
R1283 B.n434 B.n236 10.6151
R1284 B.n434 B.n433 10.6151
R1285 B.n433 B.n238 10.6151
R1286 B.n428 B.n238 10.6151
R1287 B.n428 B.n427 10.6151
R1288 B.n427 B.n426 10.6151
R1289 B.n426 B.n240 10.6151
R1290 B.n420 B.n240 10.6151
R1291 B.n420 B.n419 10.6151
R1292 B.n419 B.n418 10.6151
R1293 B.n418 B.n242 10.6151
R1294 B.n412 B.n242 10.6151
R1295 B.n412 B.n411 10.6151
R1296 B.n411 B.n410 10.6151
R1297 B.n410 B.n244 10.6151
R1298 B.n404 B.n244 10.6151
R1299 B.n404 B.n403 10.6151
R1300 B.n403 B.n402 10.6151
R1301 B.n402 B.n246 10.6151
R1302 B.n396 B.n246 10.6151
R1303 B.n396 B.n395 10.6151
R1304 B.n395 B.n394 10.6151
R1305 B.n394 B.n248 10.6151
R1306 B.n388 B.n248 10.6151
R1307 B.n388 B.n387 10.6151
R1308 B.n387 B.n386 10.6151
R1309 B.n386 B.n250 10.6151
R1310 B.n380 B.n250 10.6151
R1311 B.n380 B.n379 10.6151
R1312 B.n379 B.n378 10.6151
R1313 B.n378 B.n252 10.6151
R1314 B.n372 B.n252 10.6151
R1315 B.n372 B.n371 10.6151
R1316 B.n369 B.n256 10.6151
R1317 B.n363 B.n256 10.6151
R1318 B.n363 B.n362 10.6151
R1319 B.n362 B.n361 10.6151
R1320 B.n361 B.n258 10.6151
R1321 B.n355 B.n258 10.6151
R1322 B.n355 B.n354 10.6151
R1323 B.n354 B.n353 10.6151
R1324 B.n349 B.n348 10.6151
R1325 B.n348 B.n264 10.6151
R1326 B.n343 B.n264 10.6151
R1327 B.n343 B.n342 10.6151
R1328 B.n342 B.n341 10.6151
R1329 B.n341 B.n266 10.6151
R1330 B.n335 B.n266 10.6151
R1331 B.n335 B.n334 10.6151
R1332 B.n334 B.n333 10.6151
R1333 B.n333 B.n268 10.6151
R1334 B.n327 B.n268 10.6151
R1335 B.n327 B.n326 10.6151
R1336 B.n326 B.n325 10.6151
R1337 B.n325 B.n270 10.6151
R1338 B.n319 B.n270 10.6151
R1339 B.n319 B.n318 10.6151
R1340 B.n318 B.n317 10.6151
R1341 B.n317 B.n272 10.6151
R1342 B.n311 B.n272 10.6151
R1343 B.n311 B.n310 10.6151
R1344 B.n310 B.n309 10.6151
R1345 B.n309 B.n274 10.6151
R1346 B.n303 B.n274 10.6151
R1347 B.n303 B.n302 10.6151
R1348 B.n302 B.n301 10.6151
R1349 B.n301 B.n276 10.6151
R1350 B.n295 B.n276 10.6151
R1351 B.n295 B.n294 10.6151
R1352 B.n294 B.n293 10.6151
R1353 B.n293 B.n278 10.6151
R1354 B.n287 B.n278 10.6151
R1355 B.n287 B.n286 10.6151
R1356 B.n286 B.n285 10.6151
R1357 B.n285 B.n280 10.6151
R1358 B.n280 B.n232 10.6151
R1359 B.n446 B.n445 10.6151
R1360 B.n447 B.n446 10.6151
R1361 B.n447 B.n224 10.6151
R1362 B.n457 B.n224 10.6151
R1363 B.n458 B.n457 10.6151
R1364 B.n459 B.n458 10.6151
R1365 B.n459 B.n217 10.6151
R1366 B.n470 B.n217 10.6151
R1367 B.n471 B.n470 10.6151
R1368 B.n472 B.n471 10.6151
R1369 B.n472 B.n209 10.6151
R1370 B.n482 B.n209 10.6151
R1371 B.n483 B.n482 10.6151
R1372 B.n484 B.n483 10.6151
R1373 B.n484 B.n201 10.6151
R1374 B.n494 B.n201 10.6151
R1375 B.n495 B.n494 10.6151
R1376 B.n496 B.n495 10.6151
R1377 B.n496 B.n194 10.6151
R1378 B.n507 B.n194 10.6151
R1379 B.n508 B.n507 10.6151
R1380 B.n509 B.n508 10.6151
R1381 B.n509 B.n186 10.6151
R1382 B.n519 B.n186 10.6151
R1383 B.n520 B.n519 10.6151
R1384 B.n521 B.n520 10.6151
R1385 B.n521 B.n179 10.6151
R1386 B.n532 B.n179 10.6151
R1387 B.n533 B.n532 10.6151
R1388 B.n534 B.n533 10.6151
R1389 B.n534 B.n171 10.6151
R1390 B.n544 B.n171 10.6151
R1391 B.n545 B.n544 10.6151
R1392 B.n546 B.n545 10.6151
R1393 B.n546 B.n163 10.6151
R1394 B.n556 B.n163 10.6151
R1395 B.n557 B.n556 10.6151
R1396 B.n558 B.n557 10.6151
R1397 B.n558 B.n155 10.6151
R1398 B.n568 B.n155 10.6151
R1399 B.n569 B.n568 10.6151
R1400 B.n570 B.n569 10.6151
R1401 B.n570 B.n147 10.6151
R1402 B.n580 B.n147 10.6151
R1403 B.n581 B.n580 10.6151
R1404 B.n583 B.n581 10.6151
R1405 B.n583 B.n582 10.6151
R1406 B.n582 B.n139 10.6151
R1407 B.n594 B.n139 10.6151
R1408 B.n595 B.n594 10.6151
R1409 B.n596 B.n595 10.6151
R1410 B.n597 B.n596 10.6151
R1411 B.n598 B.n597 10.6151
R1412 B.n601 B.n598 10.6151
R1413 B.n602 B.n601 10.6151
R1414 B.n603 B.n602 10.6151
R1415 B.n604 B.n603 10.6151
R1416 B.n606 B.n604 10.6151
R1417 B.n607 B.n606 10.6151
R1418 B.n608 B.n607 10.6151
R1419 B.n609 B.n608 10.6151
R1420 B.n611 B.n609 10.6151
R1421 B.n612 B.n611 10.6151
R1422 B.n613 B.n612 10.6151
R1423 B.n614 B.n613 10.6151
R1424 B.n616 B.n614 10.6151
R1425 B.n617 B.n616 10.6151
R1426 B.n618 B.n617 10.6151
R1427 B.n619 B.n618 10.6151
R1428 B.n621 B.n619 10.6151
R1429 B.n622 B.n621 10.6151
R1430 B.n623 B.n622 10.6151
R1431 B.n624 B.n623 10.6151
R1432 B.n626 B.n624 10.6151
R1433 B.n627 B.n626 10.6151
R1434 B.n628 B.n627 10.6151
R1435 B.n629 B.n628 10.6151
R1436 B.n631 B.n629 10.6151
R1437 B.n632 B.n631 10.6151
R1438 B.n633 B.n632 10.6151
R1439 B.n634 B.n633 10.6151
R1440 B.n636 B.n634 10.6151
R1441 B.n637 B.n636 10.6151
R1442 B.n638 B.n637 10.6151
R1443 B.n639 B.n638 10.6151
R1444 B.n641 B.n639 10.6151
R1445 B.n642 B.n641 10.6151
R1446 B.n643 B.n642 10.6151
R1447 B.n644 B.n643 10.6151
R1448 B.n646 B.n644 10.6151
R1449 B.n647 B.n646 10.6151
R1450 B.n648 B.n647 10.6151
R1451 B.n649 B.n648 10.6151
R1452 B.n651 B.n649 10.6151
R1453 B.n652 B.n651 10.6151
R1454 B.n653 B.n652 10.6151
R1455 B.n654 B.n653 10.6151
R1456 B.n656 B.n654 10.6151
R1457 B.n657 B.n656 10.6151
R1458 B.n658 B.n657 10.6151
R1459 B.n659 B.n658 10.6151
R1460 B.n919 B.n1 10.6151
R1461 B.n919 B.n918 10.6151
R1462 B.n918 B.n917 10.6151
R1463 B.n917 B.n10 10.6151
R1464 B.n911 B.n10 10.6151
R1465 B.n911 B.n910 10.6151
R1466 B.n910 B.n909 10.6151
R1467 B.n909 B.n18 10.6151
R1468 B.n903 B.n18 10.6151
R1469 B.n903 B.n902 10.6151
R1470 B.n902 B.n901 10.6151
R1471 B.n901 B.n25 10.6151
R1472 B.n895 B.n25 10.6151
R1473 B.n895 B.n894 10.6151
R1474 B.n894 B.n893 10.6151
R1475 B.n893 B.n32 10.6151
R1476 B.n887 B.n32 10.6151
R1477 B.n887 B.n886 10.6151
R1478 B.n886 B.n885 10.6151
R1479 B.n885 B.n39 10.6151
R1480 B.n879 B.n39 10.6151
R1481 B.n879 B.n878 10.6151
R1482 B.n878 B.n877 10.6151
R1483 B.n877 B.n45 10.6151
R1484 B.n871 B.n45 10.6151
R1485 B.n871 B.n870 10.6151
R1486 B.n870 B.n869 10.6151
R1487 B.n869 B.n53 10.6151
R1488 B.n863 B.n53 10.6151
R1489 B.n863 B.n862 10.6151
R1490 B.n862 B.n861 10.6151
R1491 B.n861 B.n59 10.6151
R1492 B.n855 B.n59 10.6151
R1493 B.n855 B.n854 10.6151
R1494 B.n854 B.n853 10.6151
R1495 B.n853 B.n67 10.6151
R1496 B.n847 B.n67 10.6151
R1497 B.n847 B.n846 10.6151
R1498 B.n846 B.n845 10.6151
R1499 B.n845 B.n74 10.6151
R1500 B.n839 B.n74 10.6151
R1501 B.n839 B.n838 10.6151
R1502 B.n838 B.n837 10.6151
R1503 B.n837 B.n80 10.6151
R1504 B.n831 B.n80 10.6151
R1505 B.n831 B.n830 10.6151
R1506 B.n830 B.n829 10.6151
R1507 B.n829 B.n88 10.6151
R1508 B.n823 B.n88 10.6151
R1509 B.n822 B.n821 10.6151
R1510 B.n821 B.n95 10.6151
R1511 B.n815 B.n95 10.6151
R1512 B.n815 B.n814 10.6151
R1513 B.n814 B.n813 10.6151
R1514 B.n813 B.n97 10.6151
R1515 B.n807 B.n97 10.6151
R1516 B.n807 B.n806 10.6151
R1517 B.n806 B.n805 10.6151
R1518 B.n805 B.n99 10.6151
R1519 B.n799 B.n99 10.6151
R1520 B.n799 B.n798 10.6151
R1521 B.n798 B.n797 10.6151
R1522 B.n797 B.n101 10.6151
R1523 B.n791 B.n101 10.6151
R1524 B.n791 B.n790 10.6151
R1525 B.n790 B.n789 10.6151
R1526 B.n789 B.n103 10.6151
R1527 B.n783 B.n103 10.6151
R1528 B.n783 B.n782 10.6151
R1529 B.n782 B.n781 10.6151
R1530 B.n781 B.n105 10.6151
R1531 B.n775 B.n105 10.6151
R1532 B.n775 B.n774 10.6151
R1533 B.n774 B.n773 10.6151
R1534 B.n773 B.n107 10.6151
R1535 B.n767 B.n107 10.6151
R1536 B.n767 B.n766 10.6151
R1537 B.n766 B.n765 10.6151
R1538 B.n765 B.n109 10.6151
R1539 B.n759 B.n109 10.6151
R1540 B.n759 B.n758 10.6151
R1541 B.n758 B.n757 10.6151
R1542 B.n757 B.n111 10.6151
R1543 B.n751 B.n111 10.6151
R1544 B.n749 B.n748 10.6151
R1545 B.n748 B.n115 10.6151
R1546 B.n742 B.n115 10.6151
R1547 B.n742 B.n741 10.6151
R1548 B.n741 B.n740 10.6151
R1549 B.n740 B.n117 10.6151
R1550 B.n734 B.n117 10.6151
R1551 B.n734 B.n733 10.6151
R1552 B.n731 B.n121 10.6151
R1553 B.n725 B.n121 10.6151
R1554 B.n725 B.n724 10.6151
R1555 B.n724 B.n723 10.6151
R1556 B.n723 B.n123 10.6151
R1557 B.n717 B.n123 10.6151
R1558 B.n717 B.n716 10.6151
R1559 B.n716 B.n715 10.6151
R1560 B.n715 B.n125 10.6151
R1561 B.n709 B.n125 10.6151
R1562 B.n709 B.n708 10.6151
R1563 B.n708 B.n707 10.6151
R1564 B.n707 B.n127 10.6151
R1565 B.n701 B.n127 10.6151
R1566 B.n701 B.n700 10.6151
R1567 B.n700 B.n699 10.6151
R1568 B.n699 B.n129 10.6151
R1569 B.n693 B.n129 10.6151
R1570 B.n693 B.n692 10.6151
R1571 B.n692 B.n691 10.6151
R1572 B.n691 B.n131 10.6151
R1573 B.n685 B.n131 10.6151
R1574 B.n685 B.n684 10.6151
R1575 B.n684 B.n683 10.6151
R1576 B.n683 B.n133 10.6151
R1577 B.n677 B.n133 10.6151
R1578 B.n677 B.n676 10.6151
R1579 B.n676 B.n675 10.6151
R1580 B.n675 B.n135 10.6151
R1581 B.n669 B.n135 10.6151
R1582 B.n669 B.n668 10.6151
R1583 B.n668 B.n667 10.6151
R1584 B.n667 B.n137 10.6151
R1585 B.n661 B.n137 10.6151
R1586 B.n661 B.n660 10.6151
R1587 B.n927 B.n0 8.11757
R1588 B.n927 B.n1 8.11757
R1589 B.n370 B.n369 6.5566
R1590 B.n353 B.n262 6.5566
R1591 B.n750 B.n749 6.5566
R1592 B.n733 B.n732 6.5566
R1593 B.n554 B.t5 5.01842
R1594 B.t2 B.n897 5.01842
R1595 B.n371 B.n370 4.05904
R1596 B.n349 B.n262 4.05904
R1597 B.n751 B.n750 4.05904
R1598 B.n732 B.n731 4.05904
R1599 B.n498 B.t3 2.15104
R1600 B.n61 B.t4 2.15104
R1601 VP.n19 VP.n16 161.3
R1602 VP.n21 VP.n20 161.3
R1603 VP.n22 VP.n15 161.3
R1604 VP.n24 VP.n23 161.3
R1605 VP.n25 VP.n14 161.3
R1606 VP.n27 VP.n26 161.3
R1607 VP.n29 VP.n28 161.3
R1608 VP.n30 VP.n12 161.3
R1609 VP.n32 VP.n31 161.3
R1610 VP.n33 VP.n11 161.3
R1611 VP.n35 VP.n34 161.3
R1612 VP.n36 VP.n10 161.3
R1613 VP.n68 VP.n0 161.3
R1614 VP.n67 VP.n66 161.3
R1615 VP.n65 VP.n1 161.3
R1616 VP.n64 VP.n63 161.3
R1617 VP.n62 VP.n2 161.3
R1618 VP.n61 VP.n60 161.3
R1619 VP.n59 VP.n58 161.3
R1620 VP.n57 VP.n4 161.3
R1621 VP.n56 VP.n55 161.3
R1622 VP.n54 VP.n5 161.3
R1623 VP.n53 VP.n52 161.3
R1624 VP.n51 VP.n6 161.3
R1625 VP.n49 VP.n48 161.3
R1626 VP.n47 VP.n7 161.3
R1627 VP.n46 VP.n45 161.3
R1628 VP.n44 VP.n8 161.3
R1629 VP.n43 VP.n42 161.3
R1630 VP.n41 VP.n9 161.3
R1631 VP.n17 VP.t4 126.424
R1632 VP.n40 VP.n39 105.864
R1633 VP.n70 VP.n69 105.864
R1634 VP.n38 VP.n37 105.864
R1635 VP.n39 VP.t5 94.4312
R1636 VP.n50 VP.t7 94.4312
R1637 VP.n3 VP.t2 94.4312
R1638 VP.n69 VP.t3 94.4312
R1639 VP.n37 VP.t0 94.4312
R1640 VP.n13 VP.t6 94.4312
R1641 VP.n18 VP.t1 94.4312
R1642 VP.n18 VP.n17 62.5139
R1643 VP.n56 VP.n5 56.5193
R1644 VP.n24 VP.n15 56.5193
R1645 VP.n45 VP.n44 55.0624
R1646 VP.n63 VP.n1 55.0624
R1647 VP.n31 VP.n11 55.0624
R1648 VP.n40 VP.n38 49.2269
R1649 VP.n45 VP.n7 25.9244
R1650 VP.n63 VP.n62 25.9244
R1651 VP.n31 VP.n30 25.9244
R1652 VP.n43 VP.n9 24.4675
R1653 VP.n44 VP.n43 24.4675
R1654 VP.n49 VP.n7 24.4675
R1655 VP.n52 VP.n51 24.4675
R1656 VP.n52 VP.n5 24.4675
R1657 VP.n57 VP.n56 24.4675
R1658 VP.n58 VP.n57 24.4675
R1659 VP.n62 VP.n61 24.4675
R1660 VP.n67 VP.n1 24.4675
R1661 VP.n68 VP.n67 24.4675
R1662 VP.n35 VP.n11 24.4675
R1663 VP.n36 VP.n35 24.4675
R1664 VP.n25 VP.n24 24.4675
R1665 VP.n26 VP.n25 24.4675
R1666 VP.n30 VP.n29 24.4675
R1667 VP.n20 VP.n19 24.4675
R1668 VP.n20 VP.n15 24.4675
R1669 VP.n50 VP.n49 14.6807
R1670 VP.n61 VP.n3 14.6807
R1671 VP.n29 VP.n13 14.6807
R1672 VP.n51 VP.n50 9.7873
R1673 VP.n58 VP.n3 9.7873
R1674 VP.n26 VP.n13 9.7873
R1675 VP.n19 VP.n18 9.7873
R1676 VP.n17 VP.n16 7.17076
R1677 VP.n39 VP.n9 4.8939
R1678 VP.n69 VP.n68 4.8939
R1679 VP.n37 VP.n36 4.8939
R1680 VP.n38 VP.n10 0.278367
R1681 VP.n41 VP.n40 0.278367
R1682 VP.n70 VP.n0 0.278367
R1683 VP.n21 VP.n16 0.189894
R1684 VP.n22 VP.n21 0.189894
R1685 VP.n23 VP.n22 0.189894
R1686 VP.n23 VP.n14 0.189894
R1687 VP.n27 VP.n14 0.189894
R1688 VP.n28 VP.n27 0.189894
R1689 VP.n28 VP.n12 0.189894
R1690 VP.n32 VP.n12 0.189894
R1691 VP.n33 VP.n32 0.189894
R1692 VP.n34 VP.n33 0.189894
R1693 VP.n34 VP.n10 0.189894
R1694 VP.n42 VP.n41 0.189894
R1695 VP.n42 VP.n8 0.189894
R1696 VP.n46 VP.n8 0.189894
R1697 VP.n47 VP.n46 0.189894
R1698 VP.n48 VP.n47 0.189894
R1699 VP.n48 VP.n6 0.189894
R1700 VP.n53 VP.n6 0.189894
R1701 VP.n54 VP.n53 0.189894
R1702 VP.n55 VP.n54 0.189894
R1703 VP.n55 VP.n4 0.189894
R1704 VP.n59 VP.n4 0.189894
R1705 VP.n60 VP.n59 0.189894
R1706 VP.n60 VP.n2 0.189894
R1707 VP.n64 VP.n2 0.189894
R1708 VP.n65 VP.n64 0.189894
R1709 VP.n66 VP.n65 0.189894
R1710 VP.n66 VP.n0 0.189894
R1711 VP VP.n70 0.153454
R1712 VTAIL.n434 VTAIL.n386 289.615
R1713 VTAIL.n50 VTAIL.n2 289.615
R1714 VTAIL.n104 VTAIL.n56 289.615
R1715 VTAIL.n160 VTAIL.n112 289.615
R1716 VTAIL.n380 VTAIL.n332 289.615
R1717 VTAIL.n324 VTAIL.n276 289.615
R1718 VTAIL.n270 VTAIL.n222 289.615
R1719 VTAIL.n214 VTAIL.n166 289.615
R1720 VTAIL.n402 VTAIL.n401 185
R1721 VTAIL.n407 VTAIL.n406 185
R1722 VTAIL.n409 VTAIL.n408 185
R1723 VTAIL.n398 VTAIL.n397 185
R1724 VTAIL.n415 VTAIL.n414 185
R1725 VTAIL.n417 VTAIL.n416 185
R1726 VTAIL.n394 VTAIL.n393 185
R1727 VTAIL.n424 VTAIL.n423 185
R1728 VTAIL.n425 VTAIL.n392 185
R1729 VTAIL.n427 VTAIL.n426 185
R1730 VTAIL.n390 VTAIL.n389 185
R1731 VTAIL.n433 VTAIL.n432 185
R1732 VTAIL.n435 VTAIL.n434 185
R1733 VTAIL.n18 VTAIL.n17 185
R1734 VTAIL.n23 VTAIL.n22 185
R1735 VTAIL.n25 VTAIL.n24 185
R1736 VTAIL.n14 VTAIL.n13 185
R1737 VTAIL.n31 VTAIL.n30 185
R1738 VTAIL.n33 VTAIL.n32 185
R1739 VTAIL.n10 VTAIL.n9 185
R1740 VTAIL.n40 VTAIL.n39 185
R1741 VTAIL.n41 VTAIL.n8 185
R1742 VTAIL.n43 VTAIL.n42 185
R1743 VTAIL.n6 VTAIL.n5 185
R1744 VTAIL.n49 VTAIL.n48 185
R1745 VTAIL.n51 VTAIL.n50 185
R1746 VTAIL.n72 VTAIL.n71 185
R1747 VTAIL.n77 VTAIL.n76 185
R1748 VTAIL.n79 VTAIL.n78 185
R1749 VTAIL.n68 VTAIL.n67 185
R1750 VTAIL.n85 VTAIL.n84 185
R1751 VTAIL.n87 VTAIL.n86 185
R1752 VTAIL.n64 VTAIL.n63 185
R1753 VTAIL.n94 VTAIL.n93 185
R1754 VTAIL.n95 VTAIL.n62 185
R1755 VTAIL.n97 VTAIL.n96 185
R1756 VTAIL.n60 VTAIL.n59 185
R1757 VTAIL.n103 VTAIL.n102 185
R1758 VTAIL.n105 VTAIL.n104 185
R1759 VTAIL.n128 VTAIL.n127 185
R1760 VTAIL.n133 VTAIL.n132 185
R1761 VTAIL.n135 VTAIL.n134 185
R1762 VTAIL.n124 VTAIL.n123 185
R1763 VTAIL.n141 VTAIL.n140 185
R1764 VTAIL.n143 VTAIL.n142 185
R1765 VTAIL.n120 VTAIL.n119 185
R1766 VTAIL.n150 VTAIL.n149 185
R1767 VTAIL.n151 VTAIL.n118 185
R1768 VTAIL.n153 VTAIL.n152 185
R1769 VTAIL.n116 VTAIL.n115 185
R1770 VTAIL.n159 VTAIL.n158 185
R1771 VTAIL.n161 VTAIL.n160 185
R1772 VTAIL.n381 VTAIL.n380 185
R1773 VTAIL.n379 VTAIL.n378 185
R1774 VTAIL.n336 VTAIL.n335 185
R1775 VTAIL.n373 VTAIL.n372 185
R1776 VTAIL.n371 VTAIL.n338 185
R1777 VTAIL.n370 VTAIL.n369 185
R1778 VTAIL.n341 VTAIL.n339 185
R1779 VTAIL.n364 VTAIL.n363 185
R1780 VTAIL.n362 VTAIL.n361 185
R1781 VTAIL.n345 VTAIL.n344 185
R1782 VTAIL.n356 VTAIL.n355 185
R1783 VTAIL.n354 VTAIL.n353 185
R1784 VTAIL.n349 VTAIL.n348 185
R1785 VTAIL.n325 VTAIL.n324 185
R1786 VTAIL.n323 VTAIL.n322 185
R1787 VTAIL.n280 VTAIL.n279 185
R1788 VTAIL.n317 VTAIL.n316 185
R1789 VTAIL.n315 VTAIL.n282 185
R1790 VTAIL.n314 VTAIL.n313 185
R1791 VTAIL.n285 VTAIL.n283 185
R1792 VTAIL.n308 VTAIL.n307 185
R1793 VTAIL.n306 VTAIL.n305 185
R1794 VTAIL.n289 VTAIL.n288 185
R1795 VTAIL.n300 VTAIL.n299 185
R1796 VTAIL.n298 VTAIL.n297 185
R1797 VTAIL.n293 VTAIL.n292 185
R1798 VTAIL.n271 VTAIL.n270 185
R1799 VTAIL.n269 VTAIL.n268 185
R1800 VTAIL.n226 VTAIL.n225 185
R1801 VTAIL.n263 VTAIL.n262 185
R1802 VTAIL.n261 VTAIL.n228 185
R1803 VTAIL.n260 VTAIL.n259 185
R1804 VTAIL.n231 VTAIL.n229 185
R1805 VTAIL.n254 VTAIL.n253 185
R1806 VTAIL.n252 VTAIL.n251 185
R1807 VTAIL.n235 VTAIL.n234 185
R1808 VTAIL.n246 VTAIL.n245 185
R1809 VTAIL.n244 VTAIL.n243 185
R1810 VTAIL.n239 VTAIL.n238 185
R1811 VTAIL.n215 VTAIL.n214 185
R1812 VTAIL.n213 VTAIL.n212 185
R1813 VTAIL.n170 VTAIL.n169 185
R1814 VTAIL.n207 VTAIL.n206 185
R1815 VTAIL.n205 VTAIL.n172 185
R1816 VTAIL.n204 VTAIL.n203 185
R1817 VTAIL.n175 VTAIL.n173 185
R1818 VTAIL.n198 VTAIL.n197 185
R1819 VTAIL.n196 VTAIL.n195 185
R1820 VTAIL.n179 VTAIL.n178 185
R1821 VTAIL.n190 VTAIL.n189 185
R1822 VTAIL.n188 VTAIL.n187 185
R1823 VTAIL.n183 VTAIL.n182 185
R1824 VTAIL.n403 VTAIL.t3 149.524
R1825 VTAIL.n19 VTAIL.t0 149.524
R1826 VTAIL.n73 VTAIL.t8 149.524
R1827 VTAIL.n129 VTAIL.t9 149.524
R1828 VTAIL.n350 VTAIL.t12 149.524
R1829 VTAIL.n294 VTAIL.t11 149.524
R1830 VTAIL.n240 VTAIL.t4 149.524
R1831 VTAIL.n184 VTAIL.t2 149.524
R1832 VTAIL.n407 VTAIL.n401 104.615
R1833 VTAIL.n408 VTAIL.n407 104.615
R1834 VTAIL.n408 VTAIL.n397 104.615
R1835 VTAIL.n415 VTAIL.n397 104.615
R1836 VTAIL.n416 VTAIL.n415 104.615
R1837 VTAIL.n416 VTAIL.n393 104.615
R1838 VTAIL.n424 VTAIL.n393 104.615
R1839 VTAIL.n425 VTAIL.n424 104.615
R1840 VTAIL.n426 VTAIL.n425 104.615
R1841 VTAIL.n426 VTAIL.n389 104.615
R1842 VTAIL.n433 VTAIL.n389 104.615
R1843 VTAIL.n434 VTAIL.n433 104.615
R1844 VTAIL.n23 VTAIL.n17 104.615
R1845 VTAIL.n24 VTAIL.n23 104.615
R1846 VTAIL.n24 VTAIL.n13 104.615
R1847 VTAIL.n31 VTAIL.n13 104.615
R1848 VTAIL.n32 VTAIL.n31 104.615
R1849 VTAIL.n32 VTAIL.n9 104.615
R1850 VTAIL.n40 VTAIL.n9 104.615
R1851 VTAIL.n41 VTAIL.n40 104.615
R1852 VTAIL.n42 VTAIL.n41 104.615
R1853 VTAIL.n42 VTAIL.n5 104.615
R1854 VTAIL.n49 VTAIL.n5 104.615
R1855 VTAIL.n50 VTAIL.n49 104.615
R1856 VTAIL.n77 VTAIL.n71 104.615
R1857 VTAIL.n78 VTAIL.n77 104.615
R1858 VTAIL.n78 VTAIL.n67 104.615
R1859 VTAIL.n85 VTAIL.n67 104.615
R1860 VTAIL.n86 VTAIL.n85 104.615
R1861 VTAIL.n86 VTAIL.n63 104.615
R1862 VTAIL.n94 VTAIL.n63 104.615
R1863 VTAIL.n95 VTAIL.n94 104.615
R1864 VTAIL.n96 VTAIL.n95 104.615
R1865 VTAIL.n96 VTAIL.n59 104.615
R1866 VTAIL.n103 VTAIL.n59 104.615
R1867 VTAIL.n104 VTAIL.n103 104.615
R1868 VTAIL.n133 VTAIL.n127 104.615
R1869 VTAIL.n134 VTAIL.n133 104.615
R1870 VTAIL.n134 VTAIL.n123 104.615
R1871 VTAIL.n141 VTAIL.n123 104.615
R1872 VTAIL.n142 VTAIL.n141 104.615
R1873 VTAIL.n142 VTAIL.n119 104.615
R1874 VTAIL.n150 VTAIL.n119 104.615
R1875 VTAIL.n151 VTAIL.n150 104.615
R1876 VTAIL.n152 VTAIL.n151 104.615
R1877 VTAIL.n152 VTAIL.n115 104.615
R1878 VTAIL.n159 VTAIL.n115 104.615
R1879 VTAIL.n160 VTAIL.n159 104.615
R1880 VTAIL.n380 VTAIL.n379 104.615
R1881 VTAIL.n379 VTAIL.n335 104.615
R1882 VTAIL.n372 VTAIL.n335 104.615
R1883 VTAIL.n372 VTAIL.n371 104.615
R1884 VTAIL.n371 VTAIL.n370 104.615
R1885 VTAIL.n370 VTAIL.n339 104.615
R1886 VTAIL.n363 VTAIL.n339 104.615
R1887 VTAIL.n363 VTAIL.n362 104.615
R1888 VTAIL.n362 VTAIL.n344 104.615
R1889 VTAIL.n355 VTAIL.n344 104.615
R1890 VTAIL.n355 VTAIL.n354 104.615
R1891 VTAIL.n354 VTAIL.n348 104.615
R1892 VTAIL.n324 VTAIL.n323 104.615
R1893 VTAIL.n323 VTAIL.n279 104.615
R1894 VTAIL.n316 VTAIL.n279 104.615
R1895 VTAIL.n316 VTAIL.n315 104.615
R1896 VTAIL.n315 VTAIL.n314 104.615
R1897 VTAIL.n314 VTAIL.n283 104.615
R1898 VTAIL.n307 VTAIL.n283 104.615
R1899 VTAIL.n307 VTAIL.n306 104.615
R1900 VTAIL.n306 VTAIL.n288 104.615
R1901 VTAIL.n299 VTAIL.n288 104.615
R1902 VTAIL.n299 VTAIL.n298 104.615
R1903 VTAIL.n298 VTAIL.n292 104.615
R1904 VTAIL.n270 VTAIL.n269 104.615
R1905 VTAIL.n269 VTAIL.n225 104.615
R1906 VTAIL.n262 VTAIL.n225 104.615
R1907 VTAIL.n262 VTAIL.n261 104.615
R1908 VTAIL.n261 VTAIL.n260 104.615
R1909 VTAIL.n260 VTAIL.n229 104.615
R1910 VTAIL.n253 VTAIL.n229 104.615
R1911 VTAIL.n253 VTAIL.n252 104.615
R1912 VTAIL.n252 VTAIL.n234 104.615
R1913 VTAIL.n245 VTAIL.n234 104.615
R1914 VTAIL.n245 VTAIL.n244 104.615
R1915 VTAIL.n244 VTAIL.n238 104.615
R1916 VTAIL.n214 VTAIL.n213 104.615
R1917 VTAIL.n213 VTAIL.n169 104.615
R1918 VTAIL.n206 VTAIL.n169 104.615
R1919 VTAIL.n206 VTAIL.n205 104.615
R1920 VTAIL.n205 VTAIL.n204 104.615
R1921 VTAIL.n204 VTAIL.n173 104.615
R1922 VTAIL.n197 VTAIL.n173 104.615
R1923 VTAIL.n197 VTAIL.n196 104.615
R1924 VTAIL.n196 VTAIL.n178 104.615
R1925 VTAIL.n189 VTAIL.n178 104.615
R1926 VTAIL.n189 VTAIL.n188 104.615
R1927 VTAIL.n188 VTAIL.n182 104.615
R1928 VTAIL.t3 VTAIL.n401 52.3082
R1929 VTAIL.t0 VTAIL.n17 52.3082
R1930 VTAIL.t8 VTAIL.n71 52.3082
R1931 VTAIL.t9 VTAIL.n127 52.3082
R1932 VTAIL.t12 VTAIL.n348 52.3082
R1933 VTAIL.t11 VTAIL.n292 52.3082
R1934 VTAIL.t4 VTAIL.n238 52.3082
R1935 VTAIL.t2 VTAIL.n182 52.3082
R1936 VTAIL.n331 VTAIL.n330 48.0949
R1937 VTAIL.n221 VTAIL.n220 48.0949
R1938 VTAIL.n1 VTAIL.n0 48.0947
R1939 VTAIL.n111 VTAIL.n110 48.0947
R1940 VTAIL.n439 VTAIL.n438 34.3187
R1941 VTAIL.n55 VTAIL.n54 34.3187
R1942 VTAIL.n109 VTAIL.n108 34.3187
R1943 VTAIL.n165 VTAIL.n164 34.3187
R1944 VTAIL.n385 VTAIL.n384 34.3187
R1945 VTAIL.n329 VTAIL.n328 34.3187
R1946 VTAIL.n275 VTAIL.n274 34.3187
R1947 VTAIL.n219 VTAIL.n218 34.3187
R1948 VTAIL.n439 VTAIL.n385 23.5479
R1949 VTAIL.n219 VTAIL.n165 23.5479
R1950 VTAIL.n427 VTAIL.n392 13.1884
R1951 VTAIL.n43 VTAIL.n8 13.1884
R1952 VTAIL.n97 VTAIL.n62 13.1884
R1953 VTAIL.n153 VTAIL.n118 13.1884
R1954 VTAIL.n373 VTAIL.n338 13.1884
R1955 VTAIL.n317 VTAIL.n282 13.1884
R1956 VTAIL.n263 VTAIL.n228 13.1884
R1957 VTAIL.n207 VTAIL.n172 13.1884
R1958 VTAIL.n423 VTAIL.n422 12.8005
R1959 VTAIL.n428 VTAIL.n390 12.8005
R1960 VTAIL.n39 VTAIL.n38 12.8005
R1961 VTAIL.n44 VTAIL.n6 12.8005
R1962 VTAIL.n93 VTAIL.n92 12.8005
R1963 VTAIL.n98 VTAIL.n60 12.8005
R1964 VTAIL.n149 VTAIL.n148 12.8005
R1965 VTAIL.n154 VTAIL.n116 12.8005
R1966 VTAIL.n374 VTAIL.n336 12.8005
R1967 VTAIL.n369 VTAIL.n340 12.8005
R1968 VTAIL.n318 VTAIL.n280 12.8005
R1969 VTAIL.n313 VTAIL.n284 12.8005
R1970 VTAIL.n264 VTAIL.n226 12.8005
R1971 VTAIL.n259 VTAIL.n230 12.8005
R1972 VTAIL.n208 VTAIL.n170 12.8005
R1973 VTAIL.n203 VTAIL.n174 12.8005
R1974 VTAIL.n421 VTAIL.n394 12.0247
R1975 VTAIL.n432 VTAIL.n431 12.0247
R1976 VTAIL.n37 VTAIL.n10 12.0247
R1977 VTAIL.n48 VTAIL.n47 12.0247
R1978 VTAIL.n91 VTAIL.n64 12.0247
R1979 VTAIL.n102 VTAIL.n101 12.0247
R1980 VTAIL.n147 VTAIL.n120 12.0247
R1981 VTAIL.n158 VTAIL.n157 12.0247
R1982 VTAIL.n378 VTAIL.n377 12.0247
R1983 VTAIL.n368 VTAIL.n341 12.0247
R1984 VTAIL.n322 VTAIL.n321 12.0247
R1985 VTAIL.n312 VTAIL.n285 12.0247
R1986 VTAIL.n268 VTAIL.n267 12.0247
R1987 VTAIL.n258 VTAIL.n231 12.0247
R1988 VTAIL.n212 VTAIL.n211 12.0247
R1989 VTAIL.n202 VTAIL.n175 12.0247
R1990 VTAIL.n418 VTAIL.n417 11.249
R1991 VTAIL.n435 VTAIL.n388 11.249
R1992 VTAIL.n34 VTAIL.n33 11.249
R1993 VTAIL.n51 VTAIL.n4 11.249
R1994 VTAIL.n88 VTAIL.n87 11.249
R1995 VTAIL.n105 VTAIL.n58 11.249
R1996 VTAIL.n144 VTAIL.n143 11.249
R1997 VTAIL.n161 VTAIL.n114 11.249
R1998 VTAIL.n381 VTAIL.n334 11.249
R1999 VTAIL.n365 VTAIL.n364 11.249
R2000 VTAIL.n325 VTAIL.n278 11.249
R2001 VTAIL.n309 VTAIL.n308 11.249
R2002 VTAIL.n271 VTAIL.n224 11.249
R2003 VTAIL.n255 VTAIL.n254 11.249
R2004 VTAIL.n215 VTAIL.n168 11.249
R2005 VTAIL.n199 VTAIL.n198 11.249
R2006 VTAIL.n414 VTAIL.n396 10.4732
R2007 VTAIL.n436 VTAIL.n386 10.4732
R2008 VTAIL.n30 VTAIL.n12 10.4732
R2009 VTAIL.n52 VTAIL.n2 10.4732
R2010 VTAIL.n84 VTAIL.n66 10.4732
R2011 VTAIL.n106 VTAIL.n56 10.4732
R2012 VTAIL.n140 VTAIL.n122 10.4732
R2013 VTAIL.n162 VTAIL.n112 10.4732
R2014 VTAIL.n382 VTAIL.n332 10.4732
R2015 VTAIL.n361 VTAIL.n343 10.4732
R2016 VTAIL.n326 VTAIL.n276 10.4732
R2017 VTAIL.n305 VTAIL.n287 10.4732
R2018 VTAIL.n272 VTAIL.n222 10.4732
R2019 VTAIL.n251 VTAIL.n233 10.4732
R2020 VTAIL.n216 VTAIL.n166 10.4732
R2021 VTAIL.n195 VTAIL.n177 10.4732
R2022 VTAIL.n403 VTAIL.n402 10.2747
R2023 VTAIL.n19 VTAIL.n18 10.2747
R2024 VTAIL.n73 VTAIL.n72 10.2747
R2025 VTAIL.n129 VTAIL.n128 10.2747
R2026 VTAIL.n350 VTAIL.n349 10.2747
R2027 VTAIL.n294 VTAIL.n293 10.2747
R2028 VTAIL.n240 VTAIL.n239 10.2747
R2029 VTAIL.n184 VTAIL.n183 10.2747
R2030 VTAIL.n413 VTAIL.n398 9.69747
R2031 VTAIL.n29 VTAIL.n14 9.69747
R2032 VTAIL.n83 VTAIL.n68 9.69747
R2033 VTAIL.n139 VTAIL.n124 9.69747
R2034 VTAIL.n360 VTAIL.n345 9.69747
R2035 VTAIL.n304 VTAIL.n289 9.69747
R2036 VTAIL.n250 VTAIL.n235 9.69747
R2037 VTAIL.n194 VTAIL.n179 9.69747
R2038 VTAIL.n438 VTAIL.n437 9.45567
R2039 VTAIL.n54 VTAIL.n53 9.45567
R2040 VTAIL.n108 VTAIL.n107 9.45567
R2041 VTAIL.n164 VTAIL.n163 9.45567
R2042 VTAIL.n384 VTAIL.n383 9.45567
R2043 VTAIL.n328 VTAIL.n327 9.45567
R2044 VTAIL.n274 VTAIL.n273 9.45567
R2045 VTAIL.n218 VTAIL.n217 9.45567
R2046 VTAIL.n437 VTAIL.n436 9.3005
R2047 VTAIL.n388 VTAIL.n387 9.3005
R2048 VTAIL.n431 VTAIL.n430 9.3005
R2049 VTAIL.n429 VTAIL.n428 9.3005
R2050 VTAIL.n405 VTAIL.n404 9.3005
R2051 VTAIL.n400 VTAIL.n399 9.3005
R2052 VTAIL.n411 VTAIL.n410 9.3005
R2053 VTAIL.n413 VTAIL.n412 9.3005
R2054 VTAIL.n396 VTAIL.n395 9.3005
R2055 VTAIL.n419 VTAIL.n418 9.3005
R2056 VTAIL.n421 VTAIL.n420 9.3005
R2057 VTAIL.n422 VTAIL.n391 9.3005
R2058 VTAIL.n53 VTAIL.n52 9.3005
R2059 VTAIL.n4 VTAIL.n3 9.3005
R2060 VTAIL.n47 VTAIL.n46 9.3005
R2061 VTAIL.n45 VTAIL.n44 9.3005
R2062 VTAIL.n21 VTAIL.n20 9.3005
R2063 VTAIL.n16 VTAIL.n15 9.3005
R2064 VTAIL.n27 VTAIL.n26 9.3005
R2065 VTAIL.n29 VTAIL.n28 9.3005
R2066 VTAIL.n12 VTAIL.n11 9.3005
R2067 VTAIL.n35 VTAIL.n34 9.3005
R2068 VTAIL.n37 VTAIL.n36 9.3005
R2069 VTAIL.n38 VTAIL.n7 9.3005
R2070 VTAIL.n107 VTAIL.n106 9.3005
R2071 VTAIL.n58 VTAIL.n57 9.3005
R2072 VTAIL.n101 VTAIL.n100 9.3005
R2073 VTAIL.n99 VTAIL.n98 9.3005
R2074 VTAIL.n75 VTAIL.n74 9.3005
R2075 VTAIL.n70 VTAIL.n69 9.3005
R2076 VTAIL.n81 VTAIL.n80 9.3005
R2077 VTAIL.n83 VTAIL.n82 9.3005
R2078 VTAIL.n66 VTAIL.n65 9.3005
R2079 VTAIL.n89 VTAIL.n88 9.3005
R2080 VTAIL.n91 VTAIL.n90 9.3005
R2081 VTAIL.n92 VTAIL.n61 9.3005
R2082 VTAIL.n163 VTAIL.n162 9.3005
R2083 VTAIL.n114 VTAIL.n113 9.3005
R2084 VTAIL.n157 VTAIL.n156 9.3005
R2085 VTAIL.n155 VTAIL.n154 9.3005
R2086 VTAIL.n131 VTAIL.n130 9.3005
R2087 VTAIL.n126 VTAIL.n125 9.3005
R2088 VTAIL.n137 VTAIL.n136 9.3005
R2089 VTAIL.n139 VTAIL.n138 9.3005
R2090 VTAIL.n122 VTAIL.n121 9.3005
R2091 VTAIL.n145 VTAIL.n144 9.3005
R2092 VTAIL.n147 VTAIL.n146 9.3005
R2093 VTAIL.n148 VTAIL.n117 9.3005
R2094 VTAIL.n352 VTAIL.n351 9.3005
R2095 VTAIL.n347 VTAIL.n346 9.3005
R2096 VTAIL.n358 VTAIL.n357 9.3005
R2097 VTAIL.n360 VTAIL.n359 9.3005
R2098 VTAIL.n343 VTAIL.n342 9.3005
R2099 VTAIL.n366 VTAIL.n365 9.3005
R2100 VTAIL.n368 VTAIL.n367 9.3005
R2101 VTAIL.n340 VTAIL.n337 9.3005
R2102 VTAIL.n383 VTAIL.n382 9.3005
R2103 VTAIL.n334 VTAIL.n333 9.3005
R2104 VTAIL.n377 VTAIL.n376 9.3005
R2105 VTAIL.n375 VTAIL.n374 9.3005
R2106 VTAIL.n296 VTAIL.n295 9.3005
R2107 VTAIL.n291 VTAIL.n290 9.3005
R2108 VTAIL.n302 VTAIL.n301 9.3005
R2109 VTAIL.n304 VTAIL.n303 9.3005
R2110 VTAIL.n287 VTAIL.n286 9.3005
R2111 VTAIL.n310 VTAIL.n309 9.3005
R2112 VTAIL.n312 VTAIL.n311 9.3005
R2113 VTAIL.n284 VTAIL.n281 9.3005
R2114 VTAIL.n327 VTAIL.n326 9.3005
R2115 VTAIL.n278 VTAIL.n277 9.3005
R2116 VTAIL.n321 VTAIL.n320 9.3005
R2117 VTAIL.n319 VTAIL.n318 9.3005
R2118 VTAIL.n242 VTAIL.n241 9.3005
R2119 VTAIL.n237 VTAIL.n236 9.3005
R2120 VTAIL.n248 VTAIL.n247 9.3005
R2121 VTAIL.n250 VTAIL.n249 9.3005
R2122 VTAIL.n233 VTAIL.n232 9.3005
R2123 VTAIL.n256 VTAIL.n255 9.3005
R2124 VTAIL.n258 VTAIL.n257 9.3005
R2125 VTAIL.n230 VTAIL.n227 9.3005
R2126 VTAIL.n273 VTAIL.n272 9.3005
R2127 VTAIL.n224 VTAIL.n223 9.3005
R2128 VTAIL.n267 VTAIL.n266 9.3005
R2129 VTAIL.n265 VTAIL.n264 9.3005
R2130 VTAIL.n186 VTAIL.n185 9.3005
R2131 VTAIL.n181 VTAIL.n180 9.3005
R2132 VTAIL.n192 VTAIL.n191 9.3005
R2133 VTAIL.n194 VTAIL.n193 9.3005
R2134 VTAIL.n177 VTAIL.n176 9.3005
R2135 VTAIL.n200 VTAIL.n199 9.3005
R2136 VTAIL.n202 VTAIL.n201 9.3005
R2137 VTAIL.n174 VTAIL.n171 9.3005
R2138 VTAIL.n217 VTAIL.n216 9.3005
R2139 VTAIL.n168 VTAIL.n167 9.3005
R2140 VTAIL.n211 VTAIL.n210 9.3005
R2141 VTAIL.n209 VTAIL.n208 9.3005
R2142 VTAIL.n410 VTAIL.n409 8.92171
R2143 VTAIL.n26 VTAIL.n25 8.92171
R2144 VTAIL.n80 VTAIL.n79 8.92171
R2145 VTAIL.n136 VTAIL.n135 8.92171
R2146 VTAIL.n357 VTAIL.n356 8.92171
R2147 VTAIL.n301 VTAIL.n300 8.92171
R2148 VTAIL.n247 VTAIL.n246 8.92171
R2149 VTAIL.n191 VTAIL.n190 8.92171
R2150 VTAIL.n406 VTAIL.n400 8.14595
R2151 VTAIL.n22 VTAIL.n16 8.14595
R2152 VTAIL.n76 VTAIL.n70 8.14595
R2153 VTAIL.n132 VTAIL.n126 8.14595
R2154 VTAIL.n353 VTAIL.n347 8.14595
R2155 VTAIL.n297 VTAIL.n291 8.14595
R2156 VTAIL.n243 VTAIL.n237 8.14595
R2157 VTAIL.n187 VTAIL.n181 8.14595
R2158 VTAIL.n405 VTAIL.n402 7.3702
R2159 VTAIL.n21 VTAIL.n18 7.3702
R2160 VTAIL.n75 VTAIL.n72 7.3702
R2161 VTAIL.n131 VTAIL.n128 7.3702
R2162 VTAIL.n352 VTAIL.n349 7.3702
R2163 VTAIL.n296 VTAIL.n293 7.3702
R2164 VTAIL.n242 VTAIL.n239 7.3702
R2165 VTAIL.n186 VTAIL.n183 7.3702
R2166 VTAIL.n406 VTAIL.n405 5.81868
R2167 VTAIL.n22 VTAIL.n21 5.81868
R2168 VTAIL.n76 VTAIL.n75 5.81868
R2169 VTAIL.n132 VTAIL.n131 5.81868
R2170 VTAIL.n353 VTAIL.n352 5.81868
R2171 VTAIL.n297 VTAIL.n296 5.81868
R2172 VTAIL.n243 VTAIL.n242 5.81868
R2173 VTAIL.n187 VTAIL.n186 5.81868
R2174 VTAIL.n409 VTAIL.n400 5.04292
R2175 VTAIL.n25 VTAIL.n16 5.04292
R2176 VTAIL.n79 VTAIL.n70 5.04292
R2177 VTAIL.n135 VTAIL.n126 5.04292
R2178 VTAIL.n356 VTAIL.n347 5.04292
R2179 VTAIL.n300 VTAIL.n291 5.04292
R2180 VTAIL.n246 VTAIL.n237 5.04292
R2181 VTAIL.n190 VTAIL.n181 5.04292
R2182 VTAIL.n410 VTAIL.n398 4.26717
R2183 VTAIL.n26 VTAIL.n14 4.26717
R2184 VTAIL.n80 VTAIL.n68 4.26717
R2185 VTAIL.n136 VTAIL.n124 4.26717
R2186 VTAIL.n357 VTAIL.n345 4.26717
R2187 VTAIL.n301 VTAIL.n289 4.26717
R2188 VTAIL.n247 VTAIL.n235 4.26717
R2189 VTAIL.n191 VTAIL.n179 4.26717
R2190 VTAIL.n414 VTAIL.n413 3.49141
R2191 VTAIL.n438 VTAIL.n386 3.49141
R2192 VTAIL.n30 VTAIL.n29 3.49141
R2193 VTAIL.n54 VTAIL.n2 3.49141
R2194 VTAIL.n84 VTAIL.n83 3.49141
R2195 VTAIL.n108 VTAIL.n56 3.49141
R2196 VTAIL.n140 VTAIL.n139 3.49141
R2197 VTAIL.n164 VTAIL.n112 3.49141
R2198 VTAIL.n384 VTAIL.n332 3.49141
R2199 VTAIL.n361 VTAIL.n360 3.49141
R2200 VTAIL.n328 VTAIL.n276 3.49141
R2201 VTAIL.n305 VTAIL.n304 3.49141
R2202 VTAIL.n274 VTAIL.n222 3.49141
R2203 VTAIL.n251 VTAIL.n250 3.49141
R2204 VTAIL.n218 VTAIL.n166 3.49141
R2205 VTAIL.n195 VTAIL.n194 3.49141
R2206 VTAIL.n404 VTAIL.n403 2.84303
R2207 VTAIL.n20 VTAIL.n19 2.84303
R2208 VTAIL.n74 VTAIL.n73 2.84303
R2209 VTAIL.n130 VTAIL.n129 2.84303
R2210 VTAIL.n351 VTAIL.n350 2.84303
R2211 VTAIL.n295 VTAIL.n294 2.84303
R2212 VTAIL.n241 VTAIL.n240 2.84303
R2213 VTAIL.n185 VTAIL.n184 2.84303
R2214 VTAIL.n417 VTAIL.n396 2.71565
R2215 VTAIL.n436 VTAIL.n435 2.71565
R2216 VTAIL.n33 VTAIL.n12 2.71565
R2217 VTAIL.n52 VTAIL.n51 2.71565
R2218 VTAIL.n87 VTAIL.n66 2.71565
R2219 VTAIL.n106 VTAIL.n105 2.71565
R2220 VTAIL.n143 VTAIL.n122 2.71565
R2221 VTAIL.n162 VTAIL.n161 2.71565
R2222 VTAIL.n382 VTAIL.n381 2.71565
R2223 VTAIL.n364 VTAIL.n343 2.71565
R2224 VTAIL.n326 VTAIL.n325 2.71565
R2225 VTAIL.n308 VTAIL.n287 2.71565
R2226 VTAIL.n272 VTAIL.n271 2.71565
R2227 VTAIL.n254 VTAIL.n233 2.71565
R2228 VTAIL.n216 VTAIL.n215 2.71565
R2229 VTAIL.n198 VTAIL.n177 2.71565
R2230 VTAIL.n221 VTAIL.n219 2.5005
R2231 VTAIL.n275 VTAIL.n221 2.5005
R2232 VTAIL.n331 VTAIL.n329 2.5005
R2233 VTAIL.n385 VTAIL.n331 2.5005
R2234 VTAIL.n165 VTAIL.n111 2.5005
R2235 VTAIL.n111 VTAIL.n109 2.5005
R2236 VTAIL.n55 VTAIL.n1 2.5005
R2237 VTAIL VTAIL.n439 2.44231
R2238 VTAIL.n0 VTAIL.t1 1.96674
R2239 VTAIL.n0 VTAIL.t15 1.96674
R2240 VTAIL.n110 VTAIL.t14 1.96674
R2241 VTAIL.n110 VTAIL.t10 1.96674
R2242 VTAIL.n330 VTAIL.t7 1.96674
R2243 VTAIL.n330 VTAIL.t13 1.96674
R2244 VTAIL.n220 VTAIL.t6 1.96674
R2245 VTAIL.n220 VTAIL.t5 1.96674
R2246 VTAIL.n418 VTAIL.n394 1.93989
R2247 VTAIL.n432 VTAIL.n388 1.93989
R2248 VTAIL.n34 VTAIL.n10 1.93989
R2249 VTAIL.n48 VTAIL.n4 1.93989
R2250 VTAIL.n88 VTAIL.n64 1.93989
R2251 VTAIL.n102 VTAIL.n58 1.93989
R2252 VTAIL.n144 VTAIL.n120 1.93989
R2253 VTAIL.n158 VTAIL.n114 1.93989
R2254 VTAIL.n378 VTAIL.n334 1.93989
R2255 VTAIL.n365 VTAIL.n341 1.93989
R2256 VTAIL.n322 VTAIL.n278 1.93989
R2257 VTAIL.n309 VTAIL.n285 1.93989
R2258 VTAIL.n268 VTAIL.n224 1.93989
R2259 VTAIL.n255 VTAIL.n231 1.93989
R2260 VTAIL.n212 VTAIL.n168 1.93989
R2261 VTAIL.n199 VTAIL.n175 1.93989
R2262 VTAIL.n423 VTAIL.n421 1.16414
R2263 VTAIL.n431 VTAIL.n390 1.16414
R2264 VTAIL.n39 VTAIL.n37 1.16414
R2265 VTAIL.n47 VTAIL.n6 1.16414
R2266 VTAIL.n93 VTAIL.n91 1.16414
R2267 VTAIL.n101 VTAIL.n60 1.16414
R2268 VTAIL.n149 VTAIL.n147 1.16414
R2269 VTAIL.n157 VTAIL.n116 1.16414
R2270 VTAIL.n377 VTAIL.n336 1.16414
R2271 VTAIL.n369 VTAIL.n368 1.16414
R2272 VTAIL.n321 VTAIL.n280 1.16414
R2273 VTAIL.n313 VTAIL.n312 1.16414
R2274 VTAIL.n267 VTAIL.n226 1.16414
R2275 VTAIL.n259 VTAIL.n258 1.16414
R2276 VTAIL.n211 VTAIL.n170 1.16414
R2277 VTAIL.n203 VTAIL.n202 1.16414
R2278 VTAIL.n329 VTAIL.n275 0.470328
R2279 VTAIL.n109 VTAIL.n55 0.470328
R2280 VTAIL.n422 VTAIL.n392 0.388379
R2281 VTAIL.n428 VTAIL.n427 0.388379
R2282 VTAIL.n38 VTAIL.n8 0.388379
R2283 VTAIL.n44 VTAIL.n43 0.388379
R2284 VTAIL.n92 VTAIL.n62 0.388379
R2285 VTAIL.n98 VTAIL.n97 0.388379
R2286 VTAIL.n148 VTAIL.n118 0.388379
R2287 VTAIL.n154 VTAIL.n153 0.388379
R2288 VTAIL.n374 VTAIL.n373 0.388379
R2289 VTAIL.n340 VTAIL.n338 0.388379
R2290 VTAIL.n318 VTAIL.n317 0.388379
R2291 VTAIL.n284 VTAIL.n282 0.388379
R2292 VTAIL.n264 VTAIL.n263 0.388379
R2293 VTAIL.n230 VTAIL.n228 0.388379
R2294 VTAIL.n208 VTAIL.n207 0.388379
R2295 VTAIL.n174 VTAIL.n172 0.388379
R2296 VTAIL.n404 VTAIL.n399 0.155672
R2297 VTAIL.n411 VTAIL.n399 0.155672
R2298 VTAIL.n412 VTAIL.n411 0.155672
R2299 VTAIL.n412 VTAIL.n395 0.155672
R2300 VTAIL.n419 VTAIL.n395 0.155672
R2301 VTAIL.n420 VTAIL.n419 0.155672
R2302 VTAIL.n420 VTAIL.n391 0.155672
R2303 VTAIL.n429 VTAIL.n391 0.155672
R2304 VTAIL.n430 VTAIL.n429 0.155672
R2305 VTAIL.n430 VTAIL.n387 0.155672
R2306 VTAIL.n437 VTAIL.n387 0.155672
R2307 VTAIL.n20 VTAIL.n15 0.155672
R2308 VTAIL.n27 VTAIL.n15 0.155672
R2309 VTAIL.n28 VTAIL.n27 0.155672
R2310 VTAIL.n28 VTAIL.n11 0.155672
R2311 VTAIL.n35 VTAIL.n11 0.155672
R2312 VTAIL.n36 VTAIL.n35 0.155672
R2313 VTAIL.n36 VTAIL.n7 0.155672
R2314 VTAIL.n45 VTAIL.n7 0.155672
R2315 VTAIL.n46 VTAIL.n45 0.155672
R2316 VTAIL.n46 VTAIL.n3 0.155672
R2317 VTAIL.n53 VTAIL.n3 0.155672
R2318 VTAIL.n74 VTAIL.n69 0.155672
R2319 VTAIL.n81 VTAIL.n69 0.155672
R2320 VTAIL.n82 VTAIL.n81 0.155672
R2321 VTAIL.n82 VTAIL.n65 0.155672
R2322 VTAIL.n89 VTAIL.n65 0.155672
R2323 VTAIL.n90 VTAIL.n89 0.155672
R2324 VTAIL.n90 VTAIL.n61 0.155672
R2325 VTAIL.n99 VTAIL.n61 0.155672
R2326 VTAIL.n100 VTAIL.n99 0.155672
R2327 VTAIL.n100 VTAIL.n57 0.155672
R2328 VTAIL.n107 VTAIL.n57 0.155672
R2329 VTAIL.n130 VTAIL.n125 0.155672
R2330 VTAIL.n137 VTAIL.n125 0.155672
R2331 VTAIL.n138 VTAIL.n137 0.155672
R2332 VTAIL.n138 VTAIL.n121 0.155672
R2333 VTAIL.n145 VTAIL.n121 0.155672
R2334 VTAIL.n146 VTAIL.n145 0.155672
R2335 VTAIL.n146 VTAIL.n117 0.155672
R2336 VTAIL.n155 VTAIL.n117 0.155672
R2337 VTAIL.n156 VTAIL.n155 0.155672
R2338 VTAIL.n156 VTAIL.n113 0.155672
R2339 VTAIL.n163 VTAIL.n113 0.155672
R2340 VTAIL.n383 VTAIL.n333 0.155672
R2341 VTAIL.n376 VTAIL.n333 0.155672
R2342 VTAIL.n376 VTAIL.n375 0.155672
R2343 VTAIL.n375 VTAIL.n337 0.155672
R2344 VTAIL.n367 VTAIL.n337 0.155672
R2345 VTAIL.n367 VTAIL.n366 0.155672
R2346 VTAIL.n366 VTAIL.n342 0.155672
R2347 VTAIL.n359 VTAIL.n342 0.155672
R2348 VTAIL.n359 VTAIL.n358 0.155672
R2349 VTAIL.n358 VTAIL.n346 0.155672
R2350 VTAIL.n351 VTAIL.n346 0.155672
R2351 VTAIL.n327 VTAIL.n277 0.155672
R2352 VTAIL.n320 VTAIL.n277 0.155672
R2353 VTAIL.n320 VTAIL.n319 0.155672
R2354 VTAIL.n319 VTAIL.n281 0.155672
R2355 VTAIL.n311 VTAIL.n281 0.155672
R2356 VTAIL.n311 VTAIL.n310 0.155672
R2357 VTAIL.n310 VTAIL.n286 0.155672
R2358 VTAIL.n303 VTAIL.n286 0.155672
R2359 VTAIL.n303 VTAIL.n302 0.155672
R2360 VTAIL.n302 VTAIL.n290 0.155672
R2361 VTAIL.n295 VTAIL.n290 0.155672
R2362 VTAIL.n273 VTAIL.n223 0.155672
R2363 VTAIL.n266 VTAIL.n223 0.155672
R2364 VTAIL.n266 VTAIL.n265 0.155672
R2365 VTAIL.n265 VTAIL.n227 0.155672
R2366 VTAIL.n257 VTAIL.n227 0.155672
R2367 VTAIL.n257 VTAIL.n256 0.155672
R2368 VTAIL.n256 VTAIL.n232 0.155672
R2369 VTAIL.n249 VTAIL.n232 0.155672
R2370 VTAIL.n249 VTAIL.n248 0.155672
R2371 VTAIL.n248 VTAIL.n236 0.155672
R2372 VTAIL.n241 VTAIL.n236 0.155672
R2373 VTAIL.n217 VTAIL.n167 0.155672
R2374 VTAIL.n210 VTAIL.n167 0.155672
R2375 VTAIL.n210 VTAIL.n209 0.155672
R2376 VTAIL.n209 VTAIL.n171 0.155672
R2377 VTAIL.n201 VTAIL.n171 0.155672
R2378 VTAIL.n201 VTAIL.n200 0.155672
R2379 VTAIL.n200 VTAIL.n176 0.155672
R2380 VTAIL.n193 VTAIL.n176 0.155672
R2381 VTAIL.n193 VTAIL.n192 0.155672
R2382 VTAIL.n192 VTAIL.n180 0.155672
R2383 VTAIL.n185 VTAIL.n180 0.155672
R2384 VTAIL VTAIL.n1 0.0586897
R2385 VDD1 VDD1.n0 66.0818
R2386 VDD1.n3 VDD1.n2 65.9681
R2387 VDD1.n3 VDD1.n1 65.9681
R2388 VDD1.n5 VDD1.n4 64.7735
R2389 VDD1.n5 VDD1.n3 44.2293
R2390 VDD1.n4 VDD1.t1 1.96674
R2391 VDD1.n4 VDD1.t7 1.96674
R2392 VDD1.n0 VDD1.t3 1.96674
R2393 VDD1.n0 VDD1.t6 1.96674
R2394 VDD1.n2 VDD1.t5 1.96674
R2395 VDD1.n2 VDD1.t4 1.96674
R2396 VDD1.n1 VDD1.t2 1.96674
R2397 VDD1.n1 VDD1.t0 1.96674
R2398 VDD1 VDD1.n5 1.19231
R2399 VN.n55 VN.n29 161.3
R2400 VN.n54 VN.n53 161.3
R2401 VN.n52 VN.n30 161.3
R2402 VN.n51 VN.n50 161.3
R2403 VN.n49 VN.n31 161.3
R2404 VN.n48 VN.n47 161.3
R2405 VN.n46 VN.n45 161.3
R2406 VN.n44 VN.n33 161.3
R2407 VN.n43 VN.n42 161.3
R2408 VN.n41 VN.n34 161.3
R2409 VN.n40 VN.n39 161.3
R2410 VN.n38 VN.n35 161.3
R2411 VN.n26 VN.n0 161.3
R2412 VN.n25 VN.n24 161.3
R2413 VN.n23 VN.n1 161.3
R2414 VN.n22 VN.n21 161.3
R2415 VN.n20 VN.n2 161.3
R2416 VN.n19 VN.n18 161.3
R2417 VN.n17 VN.n16 161.3
R2418 VN.n15 VN.n4 161.3
R2419 VN.n14 VN.n13 161.3
R2420 VN.n12 VN.n5 161.3
R2421 VN.n11 VN.n10 161.3
R2422 VN.n9 VN.n6 161.3
R2423 VN.n7 VN.t5 126.424
R2424 VN.n36 VN.t6 126.424
R2425 VN.n28 VN.n27 105.864
R2426 VN.n57 VN.n56 105.864
R2427 VN.n8 VN.t3 94.4312
R2428 VN.n3 VN.t2 94.4312
R2429 VN.n27 VN.t7 94.4312
R2430 VN.n37 VN.t1 94.4312
R2431 VN.n32 VN.t0 94.4312
R2432 VN.n56 VN.t4 94.4312
R2433 VN.n8 VN.n7 62.5139
R2434 VN.n37 VN.n36 62.5139
R2435 VN.n14 VN.n5 56.5193
R2436 VN.n43 VN.n34 56.5193
R2437 VN.n21 VN.n1 55.0624
R2438 VN.n50 VN.n30 55.0624
R2439 VN VN.n57 49.5057
R2440 VN.n21 VN.n20 25.9244
R2441 VN.n50 VN.n49 25.9244
R2442 VN.n10 VN.n9 24.4675
R2443 VN.n10 VN.n5 24.4675
R2444 VN.n15 VN.n14 24.4675
R2445 VN.n16 VN.n15 24.4675
R2446 VN.n20 VN.n19 24.4675
R2447 VN.n25 VN.n1 24.4675
R2448 VN.n26 VN.n25 24.4675
R2449 VN.n39 VN.n34 24.4675
R2450 VN.n39 VN.n38 24.4675
R2451 VN.n49 VN.n48 24.4675
R2452 VN.n45 VN.n44 24.4675
R2453 VN.n44 VN.n43 24.4675
R2454 VN.n55 VN.n54 24.4675
R2455 VN.n54 VN.n30 24.4675
R2456 VN.n19 VN.n3 14.6807
R2457 VN.n48 VN.n32 14.6807
R2458 VN.n9 VN.n8 9.7873
R2459 VN.n16 VN.n3 9.7873
R2460 VN.n38 VN.n37 9.7873
R2461 VN.n45 VN.n32 9.7873
R2462 VN.n36 VN.n35 7.17076
R2463 VN.n7 VN.n6 7.17076
R2464 VN.n27 VN.n26 4.8939
R2465 VN.n56 VN.n55 4.8939
R2466 VN.n57 VN.n29 0.278367
R2467 VN.n28 VN.n0 0.278367
R2468 VN.n53 VN.n29 0.189894
R2469 VN.n53 VN.n52 0.189894
R2470 VN.n52 VN.n51 0.189894
R2471 VN.n51 VN.n31 0.189894
R2472 VN.n47 VN.n31 0.189894
R2473 VN.n47 VN.n46 0.189894
R2474 VN.n46 VN.n33 0.189894
R2475 VN.n42 VN.n33 0.189894
R2476 VN.n42 VN.n41 0.189894
R2477 VN.n41 VN.n40 0.189894
R2478 VN.n40 VN.n35 0.189894
R2479 VN.n11 VN.n6 0.189894
R2480 VN.n12 VN.n11 0.189894
R2481 VN.n13 VN.n12 0.189894
R2482 VN.n13 VN.n4 0.189894
R2483 VN.n17 VN.n4 0.189894
R2484 VN.n18 VN.n17 0.189894
R2485 VN.n18 VN.n2 0.189894
R2486 VN.n22 VN.n2 0.189894
R2487 VN.n23 VN.n22 0.189894
R2488 VN.n24 VN.n23 0.189894
R2489 VN.n24 VN.n0 0.189894
R2490 VN VN.n28 0.153454
R2491 VDD2.n2 VDD2.n1 65.9681
R2492 VDD2.n2 VDD2.n0 65.9681
R2493 VDD2 VDD2.n5 65.9653
R2494 VDD2.n4 VDD2.n3 64.7737
R2495 VDD2.n4 VDD2.n2 43.6463
R2496 VDD2.n5 VDD2.t6 1.96674
R2497 VDD2.n5 VDD2.t1 1.96674
R2498 VDD2.n3 VDD2.t3 1.96674
R2499 VDD2.n3 VDD2.t7 1.96674
R2500 VDD2.n1 VDD2.t5 1.96674
R2501 VDD2.n1 VDD2.t0 1.96674
R2502 VDD2.n0 VDD2.t2 1.96674
R2503 VDD2.n0 VDD2.t4 1.96674
R2504 VDD2 VDD2.n4 1.30869
C0 VDD2 VP 0.516513f
C1 VN VTAIL 7.81751f
C2 VDD1 VP 7.71013f
C3 VDD2 VN 7.34671f
C4 VDD2 VTAIL 7.47383f
C5 VDD1 VN 0.151708f
C6 VDD1 VTAIL 7.41962f
C7 VDD1 VDD2 1.76198f
C8 VN VP 7.27123f
C9 VTAIL VP 7.83162f
C10 VDD2 B 5.164683f
C11 VDD1 B 5.599508f
C12 VTAIL B 9.317338f
C13 VN B 15.230999f
C14 VP B 13.843868f
C15 VDD2.t2 B 0.192936f
C16 VDD2.t4 B 0.192936f
C17 VDD2.n0 B 1.71035f
C18 VDD2.t5 B 0.192936f
C19 VDD2.t0 B 0.192936f
C20 VDD2.n1 B 1.71035f
C21 VDD2.n2 B 3.03946f
C22 VDD2.t3 B 0.192936f
C23 VDD2.t7 B 0.192936f
C24 VDD2.n3 B 1.70139f
C25 VDD2.n4 B 2.70397f
C26 VDD2.t6 B 0.192936f
C27 VDD2.t1 B 0.192936f
C28 VDD2.n5 B 1.71031f
C29 VN.n0 B 0.030025f
C30 VN.t7 B 1.59707f
C31 VN.n1 B 0.039416f
C32 VN.n2 B 0.022774f
C33 VN.t2 B 1.59707f
C34 VN.n3 B 0.571536f
C35 VN.n4 B 0.022774f
C36 VN.n5 B 0.033246f
C37 VN.n6 B 0.219098f
C38 VN.t3 B 1.59707f
C39 VN.t5 B 1.77663f
C40 VN.n7 B 0.621525f
C41 VN.n8 B 0.634784f
C42 VN.n9 B 0.029872f
C43 VN.n10 B 0.042445f
C44 VN.n11 B 0.022774f
C45 VN.n12 B 0.022774f
C46 VN.n13 B 0.022774f
C47 VN.n14 B 0.033246f
C48 VN.n15 B 0.042445f
C49 VN.n16 B 0.029872f
C50 VN.n17 B 0.022774f
C51 VN.n18 B 0.022774f
C52 VN.n19 B 0.034063f
C53 VN.n20 B 0.043551f
C54 VN.n21 B 0.02597f
C55 VN.n22 B 0.022774f
C56 VN.n23 B 0.022774f
C57 VN.n24 B 0.022774f
C58 VN.n25 B 0.042445f
C59 VN.n26 B 0.025681f
C60 VN.n27 B 0.640766f
C61 VN.n28 B 0.039494f
C62 VN.n29 B 0.030025f
C63 VN.t4 B 1.59707f
C64 VN.n30 B 0.039416f
C65 VN.n31 B 0.022774f
C66 VN.t0 B 1.59707f
C67 VN.n32 B 0.571536f
C68 VN.n33 B 0.022774f
C69 VN.n34 B 0.033246f
C70 VN.n35 B 0.219098f
C71 VN.t1 B 1.59707f
C72 VN.t6 B 1.77663f
C73 VN.n36 B 0.621525f
C74 VN.n37 B 0.634784f
C75 VN.n38 B 0.029872f
C76 VN.n39 B 0.042445f
C77 VN.n40 B 0.022774f
C78 VN.n41 B 0.022774f
C79 VN.n42 B 0.022774f
C80 VN.n43 B 0.033246f
C81 VN.n44 B 0.042445f
C82 VN.n45 B 0.029872f
C83 VN.n46 B 0.022774f
C84 VN.n47 B 0.022774f
C85 VN.n48 B 0.034063f
C86 VN.n49 B 0.043551f
C87 VN.n50 B 0.02597f
C88 VN.n51 B 0.022774f
C89 VN.n52 B 0.022774f
C90 VN.n53 B 0.022774f
C91 VN.n54 B 0.042445f
C92 VN.n55 B 0.025681f
C93 VN.n56 B 0.640766f
C94 VN.n57 B 1.25239f
C95 VDD1.t3 B 0.195663f
C96 VDD1.t6 B 0.195663f
C97 VDD1.n0 B 1.73554f
C98 VDD1.t2 B 0.195663f
C99 VDD1.t0 B 0.195663f
C100 VDD1.n1 B 1.73452f
C101 VDD1.t5 B 0.195663f
C102 VDD1.t4 B 0.195663f
C103 VDD1.n2 B 1.73452f
C104 VDD1.n3 B 3.13371f
C105 VDD1.t1 B 0.195663f
C106 VDD1.t7 B 0.195663f
C107 VDD1.n4 B 1.72543f
C108 VDD1.n5 B 2.77249f
C109 VTAIL.t1 B 0.162508f
C110 VTAIL.t15 B 0.162508f
C111 VTAIL.n0 B 1.37711f
C112 VTAIL.n1 B 0.361716f
C113 VTAIL.n2 B 0.028567f
C114 VTAIL.n3 B 0.020422f
C115 VTAIL.n4 B 0.010974f
C116 VTAIL.n5 B 0.025938f
C117 VTAIL.n6 B 0.011619f
C118 VTAIL.n7 B 0.020422f
C119 VTAIL.n8 B 0.011297f
C120 VTAIL.n9 B 0.025938f
C121 VTAIL.n10 B 0.011619f
C122 VTAIL.n11 B 0.020422f
C123 VTAIL.n12 B 0.010974f
C124 VTAIL.n13 B 0.025938f
C125 VTAIL.n14 B 0.011619f
C126 VTAIL.n15 B 0.020422f
C127 VTAIL.n16 B 0.010974f
C128 VTAIL.n17 B 0.019453f
C129 VTAIL.n18 B 0.018336f
C130 VTAIL.t0 B 0.043597f
C131 VTAIL.n19 B 0.132109f
C132 VTAIL.n20 B 0.854926f
C133 VTAIL.n21 B 0.010974f
C134 VTAIL.n22 B 0.011619f
C135 VTAIL.n23 B 0.025938f
C136 VTAIL.n24 B 0.025938f
C137 VTAIL.n25 B 0.011619f
C138 VTAIL.n26 B 0.010974f
C139 VTAIL.n27 B 0.020422f
C140 VTAIL.n28 B 0.020422f
C141 VTAIL.n29 B 0.010974f
C142 VTAIL.n30 B 0.011619f
C143 VTAIL.n31 B 0.025938f
C144 VTAIL.n32 B 0.025938f
C145 VTAIL.n33 B 0.011619f
C146 VTAIL.n34 B 0.010974f
C147 VTAIL.n35 B 0.020422f
C148 VTAIL.n36 B 0.020422f
C149 VTAIL.n37 B 0.010974f
C150 VTAIL.n38 B 0.010974f
C151 VTAIL.n39 B 0.011619f
C152 VTAIL.n40 B 0.025938f
C153 VTAIL.n41 B 0.025938f
C154 VTAIL.n42 B 0.025938f
C155 VTAIL.n43 B 0.011297f
C156 VTAIL.n44 B 0.010974f
C157 VTAIL.n45 B 0.020422f
C158 VTAIL.n46 B 0.020422f
C159 VTAIL.n47 B 0.010974f
C160 VTAIL.n48 B 0.011619f
C161 VTAIL.n49 B 0.025938f
C162 VTAIL.n50 B 0.055908f
C163 VTAIL.n51 B 0.011619f
C164 VTAIL.n52 B 0.010974f
C165 VTAIL.n53 B 0.050273f
C166 VTAIL.n54 B 0.031349f
C167 VTAIL.n55 B 0.2146f
C168 VTAIL.n56 B 0.028567f
C169 VTAIL.n57 B 0.020422f
C170 VTAIL.n58 B 0.010974f
C171 VTAIL.n59 B 0.025938f
C172 VTAIL.n60 B 0.011619f
C173 VTAIL.n61 B 0.020422f
C174 VTAIL.n62 B 0.011297f
C175 VTAIL.n63 B 0.025938f
C176 VTAIL.n64 B 0.011619f
C177 VTAIL.n65 B 0.020422f
C178 VTAIL.n66 B 0.010974f
C179 VTAIL.n67 B 0.025938f
C180 VTAIL.n68 B 0.011619f
C181 VTAIL.n69 B 0.020422f
C182 VTAIL.n70 B 0.010974f
C183 VTAIL.n71 B 0.019453f
C184 VTAIL.n72 B 0.018336f
C185 VTAIL.t8 B 0.043597f
C186 VTAIL.n73 B 0.132109f
C187 VTAIL.n74 B 0.854926f
C188 VTAIL.n75 B 0.010974f
C189 VTAIL.n76 B 0.011619f
C190 VTAIL.n77 B 0.025938f
C191 VTAIL.n78 B 0.025938f
C192 VTAIL.n79 B 0.011619f
C193 VTAIL.n80 B 0.010974f
C194 VTAIL.n81 B 0.020422f
C195 VTAIL.n82 B 0.020422f
C196 VTAIL.n83 B 0.010974f
C197 VTAIL.n84 B 0.011619f
C198 VTAIL.n85 B 0.025938f
C199 VTAIL.n86 B 0.025938f
C200 VTAIL.n87 B 0.011619f
C201 VTAIL.n88 B 0.010974f
C202 VTAIL.n89 B 0.020422f
C203 VTAIL.n90 B 0.020422f
C204 VTAIL.n91 B 0.010974f
C205 VTAIL.n92 B 0.010974f
C206 VTAIL.n93 B 0.011619f
C207 VTAIL.n94 B 0.025938f
C208 VTAIL.n95 B 0.025938f
C209 VTAIL.n96 B 0.025938f
C210 VTAIL.n97 B 0.011297f
C211 VTAIL.n98 B 0.010974f
C212 VTAIL.n99 B 0.020422f
C213 VTAIL.n100 B 0.020422f
C214 VTAIL.n101 B 0.010974f
C215 VTAIL.n102 B 0.011619f
C216 VTAIL.n103 B 0.025938f
C217 VTAIL.n104 B 0.055908f
C218 VTAIL.n105 B 0.011619f
C219 VTAIL.n106 B 0.010974f
C220 VTAIL.n107 B 0.050273f
C221 VTAIL.n108 B 0.031349f
C222 VTAIL.n109 B 0.2146f
C223 VTAIL.t14 B 0.162508f
C224 VTAIL.t10 B 0.162508f
C225 VTAIL.n110 B 1.37711f
C226 VTAIL.n111 B 0.522395f
C227 VTAIL.n112 B 0.028567f
C228 VTAIL.n113 B 0.020422f
C229 VTAIL.n114 B 0.010974f
C230 VTAIL.n115 B 0.025938f
C231 VTAIL.n116 B 0.011619f
C232 VTAIL.n117 B 0.020422f
C233 VTAIL.n118 B 0.011297f
C234 VTAIL.n119 B 0.025938f
C235 VTAIL.n120 B 0.011619f
C236 VTAIL.n121 B 0.020422f
C237 VTAIL.n122 B 0.010974f
C238 VTAIL.n123 B 0.025938f
C239 VTAIL.n124 B 0.011619f
C240 VTAIL.n125 B 0.020422f
C241 VTAIL.n126 B 0.010974f
C242 VTAIL.n127 B 0.019453f
C243 VTAIL.n128 B 0.018336f
C244 VTAIL.t9 B 0.043597f
C245 VTAIL.n129 B 0.132109f
C246 VTAIL.n130 B 0.854926f
C247 VTAIL.n131 B 0.010974f
C248 VTAIL.n132 B 0.011619f
C249 VTAIL.n133 B 0.025938f
C250 VTAIL.n134 B 0.025938f
C251 VTAIL.n135 B 0.011619f
C252 VTAIL.n136 B 0.010974f
C253 VTAIL.n137 B 0.020422f
C254 VTAIL.n138 B 0.020422f
C255 VTAIL.n139 B 0.010974f
C256 VTAIL.n140 B 0.011619f
C257 VTAIL.n141 B 0.025938f
C258 VTAIL.n142 B 0.025938f
C259 VTAIL.n143 B 0.011619f
C260 VTAIL.n144 B 0.010974f
C261 VTAIL.n145 B 0.020422f
C262 VTAIL.n146 B 0.020422f
C263 VTAIL.n147 B 0.010974f
C264 VTAIL.n148 B 0.010974f
C265 VTAIL.n149 B 0.011619f
C266 VTAIL.n150 B 0.025938f
C267 VTAIL.n151 B 0.025938f
C268 VTAIL.n152 B 0.025938f
C269 VTAIL.n153 B 0.011297f
C270 VTAIL.n154 B 0.010974f
C271 VTAIL.n155 B 0.020422f
C272 VTAIL.n156 B 0.020422f
C273 VTAIL.n157 B 0.010974f
C274 VTAIL.n158 B 0.011619f
C275 VTAIL.n159 B 0.025938f
C276 VTAIL.n160 B 0.055908f
C277 VTAIL.n161 B 0.011619f
C278 VTAIL.n162 B 0.010974f
C279 VTAIL.n163 B 0.050273f
C280 VTAIL.n164 B 0.031349f
C281 VTAIL.n165 B 1.19684f
C282 VTAIL.n166 B 0.028567f
C283 VTAIL.n167 B 0.020422f
C284 VTAIL.n168 B 0.010974f
C285 VTAIL.n169 B 0.025938f
C286 VTAIL.n170 B 0.011619f
C287 VTAIL.n171 B 0.020422f
C288 VTAIL.n172 B 0.011297f
C289 VTAIL.n173 B 0.025938f
C290 VTAIL.n174 B 0.010974f
C291 VTAIL.n175 B 0.011619f
C292 VTAIL.n176 B 0.020422f
C293 VTAIL.n177 B 0.010974f
C294 VTAIL.n178 B 0.025938f
C295 VTAIL.n179 B 0.011619f
C296 VTAIL.n180 B 0.020422f
C297 VTAIL.n181 B 0.010974f
C298 VTAIL.n182 B 0.019453f
C299 VTAIL.n183 B 0.018336f
C300 VTAIL.t2 B 0.043597f
C301 VTAIL.n184 B 0.132109f
C302 VTAIL.n185 B 0.854925f
C303 VTAIL.n186 B 0.010974f
C304 VTAIL.n187 B 0.011619f
C305 VTAIL.n188 B 0.025938f
C306 VTAIL.n189 B 0.025938f
C307 VTAIL.n190 B 0.011619f
C308 VTAIL.n191 B 0.010974f
C309 VTAIL.n192 B 0.020422f
C310 VTAIL.n193 B 0.020422f
C311 VTAIL.n194 B 0.010974f
C312 VTAIL.n195 B 0.011619f
C313 VTAIL.n196 B 0.025938f
C314 VTAIL.n197 B 0.025938f
C315 VTAIL.n198 B 0.011619f
C316 VTAIL.n199 B 0.010974f
C317 VTAIL.n200 B 0.020422f
C318 VTAIL.n201 B 0.020422f
C319 VTAIL.n202 B 0.010974f
C320 VTAIL.n203 B 0.011619f
C321 VTAIL.n204 B 0.025938f
C322 VTAIL.n205 B 0.025938f
C323 VTAIL.n206 B 0.025938f
C324 VTAIL.n207 B 0.011297f
C325 VTAIL.n208 B 0.010974f
C326 VTAIL.n209 B 0.020422f
C327 VTAIL.n210 B 0.020422f
C328 VTAIL.n211 B 0.010974f
C329 VTAIL.n212 B 0.011619f
C330 VTAIL.n213 B 0.025938f
C331 VTAIL.n214 B 0.055908f
C332 VTAIL.n215 B 0.011619f
C333 VTAIL.n216 B 0.010974f
C334 VTAIL.n217 B 0.050273f
C335 VTAIL.n218 B 0.031349f
C336 VTAIL.n219 B 1.19684f
C337 VTAIL.t6 B 0.162508f
C338 VTAIL.t5 B 0.162508f
C339 VTAIL.n220 B 1.37712f
C340 VTAIL.n221 B 0.522387f
C341 VTAIL.n222 B 0.028567f
C342 VTAIL.n223 B 0.020422f
C343 VTAIL.n224 B 0.010974f
C344 VTAIL.n225 B 0.025938f
C345 VTAIL.n226 B 0.011619f
C346 VTAIL.n227 B 0.020422f
C347 VTAIL.n228 B 0.011297f
C348 VTAIL.n229 B 0.025938f
C349 VTAIL.n230 B 0.010974f
C350 VTAIL.n231 B 0.011619f
C351 VTAIL.n232 B 0.020422f
C352 VTAIL.n233 B 0.010974f
C353 VTAIL.n234 B 0.025938f
C354 VTAIL.n235 B 0.011619f
C355 VTAIL.n236 B 0.020422f
C356 VTAIL.n237 B 0.010974f
C357 VTAIL.n238 B 0.019453f
C358 VTAIL.n239 B 0.018336f
C359 VTAIL.t4 B 0.043597f
C360 VTAIL.n240 B 0.132109f
C361 VTAIL.n241 B 0.854925f
C362 VTAIL.n242 B 0.010974f
C363 VTAIL.n243 B 0.011619f
C364 VTAIL.n244 B 0.025938f
C365 VTAIL.n245 B 0.025938f
C366 VTAIL.n246 B 0.011619f
C367 VTAIL.n247 B 0.010974f
C368 VTAIL.n248 B 0.020422f
C369 VTAIL.n249 B 0.020422f
C370 VTAIL.n250 B 0.010974f
C371 VTAIL.n251 B 0.011619f
C372 VTAIL.n252 B 0.025938f
C373 VTAIL.n253 B 0.025938f
C374 VTAIL.n254 B 0.011619f
C375 VTAIL.n255 B 0.010974f
C376 VTAIL.n256 B 0.020422f
C377 VTAIL.n257 B 0.020422f
C378 VTAIL.n258 B 0.010974f
C379 VTAIL.n259 B 0.011619f
C380 VTAIL.n260 B 0.025938f
C381 VTAIL.n261 B 0.025938f
C382 VTAIL.n262 B 0.025938f
C383 VTAIL.n263 B 0.011297f
C384 VTAIL.n264 B 0.010974f
C385 VTAIL.n265 B 0.020422f
C386 VTAIL.n266 B 0.020422f
C387 VTAIL.n267 B 0.010974f
C388 VTAIL.n268 B 0.011619f
C389 VTAIL.n269 B 0.025938f
C390 VTAIL.n270 B 0.055908f
C391 VTAIL.n271 B 0.011619f
C392 VTAIL.n272 B 0.010974f
C393 VTAIL.n273 B 0.050273f
C394 VTAIL.n274 B 0.031349f
C395 VTAIL.n275 B 0.2146f
C396 VTAIL.n276 B 0.028567f
C397 VTAIL.n277 B 0.020422f
C398 VTAIL.n278 B 0.010974f
C399 VTAIL.n279 B 0.025938f
C400 VTAIL.n280 B 0.011619f
C401 VTAIL.n281 B 0.020422f
C402 VTAIL.n282 B 0.011297f
C403 VTAIL.n283 B 0.025938f
C404 VTAIL.n284 B 0.010974f
C405 VTAIL.n285 B 0.011619f
C406 VTAIL.n286 B 0.020422f
C407 VTAIL.n287 B 0.010974f
C408 VTAIL.n288 B 0.025938f
C409 VTAIL.n289 B 0.011619f
C410 VTAIL.n290 B 0.020422f
C411 VTAIL.n291 B 0.010974f
C412 VTAIL.n292 B 0.019453f
C413 VTAIL.n293 B 0.018336f
C414 VTAIL.t11 B 0.043597f
C415 VTAIL.n294 B 0.132109f
C416 VTAIL.n295 B 0.854925f
C417 VTAIL.n296 B 0.010974f
C418 VTAIL.n297 B 0.011619f
C419 VTAIL.n298 B 0.025938f
C420 VTAIL.n299 B 0.025938f
C421 VTAIL.n300 B 0.011619f
C422 VTAIL.n301 B 0.010974f
C423 VTAIL.n302 B 0.020422f
C424 VTAIL.n303 B 0.020422f
C425 VTAIL.n304 B 0.010974f
C426 VTAIL.n305 B 0.011619f
C427 VTAIL.n306 B 0.025938f
C428 VTAIL.n307 B 0.025938f
C429 VTAIL.n308 B 0.011619f
C430 VTAIL.n309 B 0.010974f
C431 VTAIL.n310 B 0.020422f
C432 VTAIL.n311 B 0.020422f
C433 VTAIL.n312 B 0.010974f
C434 VTAIL.n313 B 0.011619f
C435 VTAIL.n314 B 0.025938f
C436 VTAIL.n315 B 0.025938f
C437 VTAIL.n316 B 0.025938f
C438 VTAIL.n317 B 0.011297f
C439 VTAIL.n318 B 0.010974f
C440 VTAIL.n319 B 0.020422f
C441 VTAIL.n320 B 0.020422f
C442 VTAIL.n321 B 0.010974f
C443 VTAIL.n322 B 0.011619f
C444 VTAIL.n323 B 0.025938f
C445 VTAIL.n324 B 0.055908f
C446 VTAIL.n325 B 0.011619f
C447 VTAIL.n326 B 0.010974f
C448 VTAIL.n327 B 0.050273f
C449 VTAIL.n328 B 0.031349f
C450 VTAIL.n329 B 0.2146f
C451 VTAIL.t7 B 0.162508f
C452 VTAIL.t13 B 0.162508f
C453 VTAIL.n330 B 1.37712f
C454 VTAIL.n331 B 0.522387f
C455 VTAIL.n332 B 0.028567f
C456 VTAIL.n333 B 0.020422f
C457 VTAIL.n334 B 0.010974f
C458 VTAIL.n335 B 0.025938f
C459 VTAIL.n336 B 0.011619f
C460 VTAIL.n337 B 0.020422f
C461 VTAIL.n338 B 0.011297f
C462 VTAIL.n339 B 0.025938f
C463 VTAIL.n340 B 0.010974f
C464 VTAIL.n341 B 0.011619f
C465 VTAIL.n342 B 0.020422f
C466 VTAIL.n343 B 0.010974f
C467 VTAIL.n344 B 0.025938f
C468 VTAIL.n345 B 0.011619f
C469 VTAIL.n346 B 0.020422f
C470 VTAIL.n347 B 0.010974f
C471 VTAIL.n348 B 0.019453f
C472 VTAIL.n349 B 0.018336f
C473 VTAIL.t12 B 0.043597f
C474 VTAIL.n350 B 0.132109f
C475 VTAIL.n351 B 0.854925f
C476 VTAIL.n352 B 0.010974f
C477 VTAIL.n353 B 0.011619f
C478 VTAIL.n354 B 0.025938f
C479 VTAIL.n355 B 0.025938f
C480 VTAIL.n356 B 0.011619f
C481 VTAIL.n357 B 0.010974f
C482 VTAIL.n358 B 0.020422f
C483 VTAIL.n359 B 0.020422f
C484 VTAIL.n360 B 0.010974f
C485 VTAIL.n361 B 0.011619f
C486 VTAIL.n362 B 0.025938f
C487 VTAIL.n363 B 0.025938f
C488 VTAIL.n364 B 0.011619f
C489 VTAIL.n365 B 0.010974f
C490 VTAIL.n366 B 0.020422f
C491 VTAIL.n367 B 0.020422f
C492 VTAIL.n368 B 0.010974f
C493 VTAIL.n369 B 0.011619f
C494 VTAIL.n370 B 0.025938f
C495 VTAIL.n371 B 0.025938f
C496 VTAIL.n372 B 0.025938f
C497 VTAIL.n373 B 0.011297f
C498 VTAIL.n374 B 0.010974f
C499 VTAIL.n375 B 0.020422f
C500 VTAIL.n376 B 0.020422f
C501 VTAIL.n377 B 0.010974f
C502 VTAIL.n378 B 0.011619f
C503 VTAIL.n379 B 0.025938f
C504 VTAIL.n380 B 0.055908f
C505 VTAIL.n381 B 0.011619f
C506 VTAIL.n382 B 0.010974f
C507 VTAIL.n383 B 0.050273f
C508 VTAIL.n384 B 0.031349f
C509 VTAIL.n385 B 1.19684f
C510 VTAIL.n386 B 0.028567f
C511 VTAIL.n387 B 0.020422f
C512 VTAIL.n388 B 0.010974f
C513 VTAIL.n389 B 0.025938f
C514 VTAIL.n390 B 0.011619f
C515 VTAIL.n391 B 0.020422f
C516 VTAIL.n392 B 0.011297f
C517 VTAIL.n393 B 0.025938f
C518 VTAIL.n394 B 0.011619f
C519 VTAIL.n395 B 0.020422f
C520 VTAIL.n396 B 0.010974f
C521 VTAIL.n397 B 0.025938f
C522 VTAIL.n398 B 0.011619f
C523 VTAIL.n399 B 0.020422f
C524 VTAIL.n400 B 0.010974f
C525 VTAIL.n401 B 0.019453f
C526 VTAIL.n402 B 0.018336f
C527 VTAIL.t3 B 0.043597f
C528 VTAIL.n403 B 0.132109f
C529 VTAIL.n404 B 0.854926f
C530 VTAIL.n405 B 0.010974f
C531 VTAIL.n406 B 0.011619f
C532 VTAIL.n407 B 0.025938f
C533 VTAIL.n408 B 0.025938f
C534 VTAIL.n409 B 0.011619f
C535 VTAIL.n410 B 0.010974f
C536 VTAIL.n411 B 0.020422f
C537 VTAIL.n412 B 0.020422f
C538 VTAIL.n413 B 0.010974f
C539 VTAIL.n414 B 0.011619f
C540 VTAIL.n415 B 0.025938f
C541 VTAIL.n416 B 0.025938f
C542 VTAIL.n417 B 0.011619f
C543 VTAIL.n418 B 0.010974f
C544 VTAIL.n419 B 0.020422f
C545 VTAIL.n420 B 0.020422f
C546 VTAIL.n421 B 0.010974f
C547 VTAIL.n422 B 0.010974f
C548 VTAIL.n423 B 0.011619f
C549 VTAIL.n424 B 0.025938f
C550 VTAIL.n425 B 0.025938f
C551 VTAIL.n426 B 0.025938f
C552 VTAIL.n427 B 0.011297f
C553 VTAIL.n428 B 0.010974f
C554 VTAIL.n429 B 0.020422f
C555 VTAIL.n430 B 0.020422f
C556 VTAIL.n431 B 0.010974f
C557 VTAIL.n432 B 0.011619f
C558 VTAIL.n433 B 0.025938f
C559 VTAIL.n434 B 0.055908f
C560 VTAIL.n435 B 0.011619f
C561 VTAIL.n436 B 0.010974f
C562 VTAIL.n437 B 0.050273f
C563 VTAIL.n438 B 0.031349f
C564 VTAIL.n439 B 1.19301f
C565 VP.n0 B 0.030605f
C566 VP.t3 B 1.62791f
C567 VP.n1 B 0.040177f
C568 VP.n2 B 0.023214f
C569 VP.t2 B 1.62791f
C570 VP.n3 B 0.582575f
C571 VP.n4 B 0.023214f
C572 VP.n5 B 0.033888f
C573 VP.n6 B 0.023214f
C574 VP.t7 B 1.62791f
C575 VP.n7 B 0.044392f
C576 VP.n8 B 0.023214f
C577 VP.n9 B 0.026177f
C578 VP.n10 B 0.030605f
C579 VP.t0 B 1.62791f
C580 VP.n11 B 0.040177f
C581 VP.n12 B 0.023214f
C582 VP.t6 B 1.62791f
C583 VP.n13 B 0.582575f
C584 VP.n14 B 0.023214f
C585 VP.n15 B 0.033888f
C586 VP.n16 B 0.22333f
C587 VP.t1 B 1.62791f
C588 VP.t4 B 1.81094f
C589 VP.n17 B 0.633529f
C590 VP.n18 B 0.647044f
C591 VP.n19 B 0.030449f
C592 VP.n20 B 0.043265f
C593 VP.n21 B 0.023214f
C594 VP.n22 B 0.023214f
C595 VP.n23 B 0.023214f
C596 VP.n24 B 0.033888f
C597 VP.n25 B 0.043265f
C598 VP.n26 B 0.030449f
C599 VP.n27 B 0.023214f
C600 VP.n28 B 0.023214f
C601 VP.n29 B 0.034721f
C602 VP.n30 B 0.044392f
C603 VP.n31 B 0.026472f
C604 VP.n32 B 0.023214f
C605 VP.n33 B 0.023214f
C606 VP.n34 B 0.023214f
C607 VP.n35 B 0.043265f
C608 VP.n36 B 0.026177f
C609 VP.n37 B 0.653142f
C610 VP.n38 B 1.26407f
C611 VP.t5 B 1.62791f
C612 VP.n39 B 0.653142f
C613 VP.n40 B 1.28102f
C614 VP.n41 B 0.030605f
C615 VP.n42 B 0.023214f
C616 VP.n43 B 0.043265f
C617 VP.n44 B 0.040177f
C618 VP.n45 B 0.026472f
C619 VP.n46 B 0.023214f
C620 VP.n47 B 0.023214f
C621 VP.n48 B 0.023214f
C622 VP.n49 B 0.034721f
C623 VP.n50 B 0.582575f
C624 VP.n51 B 0.030449f
C625 VP.n52 B 0.043265f
C626 VP.n53 B 0.023214f
C627 VP.n54 B 0.023214f
C628 VP.n55 B 0.023214f
C629 VP.n56 B 0.033888f
C630 VP.n57 B 0.043265f
C631 VP.n58 B 0.030449f
C632 VP.n59 B 0.023214f
C633 VP.n60 B 0.023214f
C634 VP.n61 B 0.034721f
C635 VP.n62 B 0.044392f
C636 VP.n63 B 0.026472f
C637 VP.n64 B 0.023214f
C638 VP.n65 B 0.023214f
C639 VP.n66 B 0.023214f
C640 VP.n67 B 0.043265f
C641 VP.n68 B 0.026177f
C642 VP.n69 B 0.653142f
C643 VP.n70 B 0.040257f
.ends

