* NGSPICE file created from diff_pair_sample_1050.ext - technology: sky130A

.subckt diff_pair_sample_1050 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=0 ps=0 w=6.49 l=3.85
X1 VTAIL.t7 VP.t0 VDD1.t2 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=1.07085 ps=6.82 w=6.49 l=3.85
X2 VDD1.t3 VP.t1 VTAIL.t6 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=1.07085 pd=6.82 as=2.5311 ps=13.76 w=6.49 l=3.85
X3 VTAIL.t0 VN.t0 VDD2.t3 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=1.07085 ps=6.82 w=6.49 l=3.85
X4 VDD2.t2 VN.t1 VTAIL.t1 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=1.07085 pd=6.82 as=2.5311 ps=13.76 w=6.49 l=3.85
X5 VDD2.t1 VN.t2 VTAIL.t2 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=1.07085 pd=6.82 as=2.5311 ps=13.76 w=6.49 l=3.85
X6 VDD1.t0 VP.t2 VTAIL.t5 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=1.07085 pd=6.82 as=2.5311 ps=13.76 w=6.49 l=3.85
X7 B.t8 B.t6 B.t7 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=0 ps=0 w=6.49 l=3.85
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=1.07085 ps=6.82 w=6.49 l=3.85
X9 VTAIL.t4 VP.t3 VDD1.t1 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=1.07085 ps=6.82 w=6.49 l=3.85
X10 B.t5 B.t3 B.t4 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=0 ps=0 w=6.49 l=3.85
X11 B.t2 B.t0 B.t1 w_n3478_n2266# sky130_fd_pr__pfet_01v8 ad=2.5311 pd=13.76 as=0 ps=0 w=6.49 l=3.85
R0 B.n456 B.n455 585
R1 B.n457 B.n58 585
R2 B.n459 B.n458 585
R3 B.n460 B.n57 585
R4 B.n462 B.n461 585
R5 B.n463 B.n56 585
R6 B.n465 B.n464 585
R7 B.n466 B.n55 585
R8 B.n468 B.n467 585
R9 B.n469 B.n54 585
R10 B.n471 B.n470 585
R11 B.n472 B.n53 585
R12 B.n474 B.n473 585
R13 B.n475 B.n52 585
R14 B.n477 B.n476 585
R15 B.n478 B.n51 585
R16 B.n480 B.n479 585
R17 B.n481 B.n50 585
R18 B.n483 B.n482 585
R19 B.n484 B.n49 585
R20 B.n486 B.n485 585
R21 B.n487 B.n48 585
R22 B.n489 B.n488 585
R23 B.n490 B.n47 585
R24 B.n492 B.n491 585
R25 B.n494 B.n493 585
R26 B.n495 B.n43 585
R27 B.n497 B.n496 585
R28 B.n498 B.n42 585
R29 B.n500 B.n499 585
R30 B.n501 B.n41 585
R31 B.n503 B.n502 585
R32 B.n504 B.n40 585
R33 B.n506 B.n505 585
R34 B.n507 B.n37 585
R35 B.n510 B.n509 585
R36 B.n511 B.n36 585
R37 B.n513 B.n512 585
R38 B.n514 B.n35 585
R39 B.n516 B.n515 585
R40 B.n517 B.n34 585
R41 B.n519 B.n518 585
R42 B.n520 B.n33 585
R43 B.n522 B.n521 585
R44 B.n523 B.n32 585
R45 B.n525 B.n524 585
R46 B.n526 B.n31 585
R47 B.n528 B.n527 585
R48 B.n529 B.n30 585
R49 B.n531 B.n530 585
R50 B.n532 B.n29 585
R51 B.n534 B.n533 585
R52 B.n535 B.n28 585
R53 B.n537 B.n536 585
R54 B.n538 B.n27 585
R55 B.n540 B.n539 585
R56 B.n541 B.n26 585
R57 B.n543 B.n542 585
R58 B.n544 B.n25 585
R59 B.n546 B.n545 585
R60 B.n454 B.n59 585
R61 B.n453 B.n452 585
R62 B.n451 B.n60 585
R63 B.n450 B.n449 585
R64 B.n448 B.n61 585
R65 B.n447 B.n446 585
R66 B.n445 B.n62 585
R67 B.n444 B.n443 585
R68 B.n442 B.n63 585
R69 B.n441 B.n440 585
R70 B.n439 B.n64 585
R71 B.n438 B.n437 585
R72 B.n436 B.n65 585
R73 B.n435 B.n434 585
R74 B.n433 B.n66 585
R75 B.n432 B.n431 585
R76 B.n430 B.n67 585
R77 B.n429 B.n428 585
R78 B.n427 B.n68 585
R79 B.n426 B.n425 585
R80 B.n424 B.n69 585
R81 B.n423 B.n422 585
R82 B.n421 B.n70 585
R83 B.n420 B.n419 585
R84 B.n418 B.n71 585
R85 B.n417 B.n416 585
R86 B.n415 B.n72 585
R87 B.n414 B.n413 585
R88 B.n412 B.n73 585
R89 B.n411 B.n410 585
R90 B.n409 B.n74 585
R91 B.n408 B.n407 585
R92 B.n406 B.n75 585
R93 B.n405 B.n404 585
R94 B.n403 B.n76 585
R95 B.n402 B.n401 585
R96 B.n400 B.n77 585
R97 B.n399 B.n398 585
R98 B.n397 B.n78 585
R99 B.n396 B.n395 585
R100 B.n394 B.n79 585
R101 B.n393 B.n392 585
R102 B.n391 B.n80 585
R103 B.n390 B.n389 585
R104 B.n388 B.n81 585
R105 B.n387 B.n386 585
R106 B.n385 B.n82 585
R107 B.n384 B.n383 585
R108 B.n382 B.n83 585
R109 B.n381 B.n380 585
R110 B.n379 B.n84 585
R111 B.n378 B.n377 585
R112 B.n376 B.n85 585
R113 B.n375 B.n374 585
R114 B.n373 B.n86 585
R115 B.n372 B.n371 585
R116 B.n370 B.n87 585
R117 B.n369 B.n368 585
R118 B.n367 B.n88 585
R119 B.n366 B.n365 585
R120 B.n364 B.n89 585
R121 B.n363 B.n362 585
R122 B.n361 B.n90 585
R123 B.n360 B.n359 585
R124 B.n358 B.n91 585
R125 B.n357 B.n356 585
R126 B.n355 B.n92 585
R127 B.n354 B.n353 585
R128 B.n352 B.n93 585
R129 B.n351 B.n350 585
R130 B.n349 B.n94 585
R131 B.n348 B.n347 585
R132 B.n346 B.n95 585
R133 B.n345 B.n344 585
R134 B.n343 B.n96 585
R135 B.n342 B.n341 585
R136 B.n340 B.n97 585
R137 B.n339 B.n338 585
R138 B.n337 B.n98 585
R139 B.n336 B.n335 585
R140 B.n334 B.n99 585
R141 B.n333 B.n332 585
R142 B.n331 B.n100 585
R143 B.n330 B.n329 585
R144 B.n328 B.n101 585
R145 B.n327 B.n326 585
R146 B.n325 B.n102 585
R147 B.n324 B.n323 585
R148 B.n322 B.n103 585
R149 B.n321 B.n320 585
R150 B.n319 B.n104 585
R151 B.n228 B.n227 585
R152 B.n229 B.n138 585
R153 B.n231 B.n230 585
R154 B.n232 B.n137 585
R155 B.n234 B.n233 585
R156 B.n235 B.n136 585
R157 B.n237 B.n236 585
R158 B.n238 B.n135 585
R159 B.n240 B.n239 585
R160 B.n241 B.n134 585
R161 B.n243 B.n242 585
R162 B.n244 B.n133 585
R163 B.n246 B.n245 585
R164 B.n247 B.n132 585
R165 B.n249 B.n248 585
R166 B.n250 B.n131 585
R167 B.n252 B.n251 585
R168 B.n253 B.n130 585
R169 B.n255 B.n254 585
R170 B.n256 B.n129 585
R171 B.n258 B.n257 585
R172 B.n259 B.n128 585
R173 B.n261 B.n260 585
R174 B.n262 B.n127 585
R175 B.n264 B.n263 585
R176 B.n266 B.n265 585
R177 B.n267 B.n123 585
R178 B.n269 B.n268 585
R179 B.n270 B.n122 585
R180 B.n272 B.n271 585
R181 B.n273 B.n121 585
R182 B.n275 B.n274 585
R183 B.n276 B.n120 585
R184 B.n278 B.n277 585
R185 B.n279 B.n117 585
R186 B.n282 B.n281 585
R187 B.n283 B.n116 585
R188 B.n285 B.n284 585
R189 B.n286 B.n115 585
R190 B.n288 B.n287 585
R191 B.n289 B.n114 585
R192 B.n291 B.n290 585
R193 B.n292 B.n113 585
R194 B.n294 B.n293 585
R195 B.n295 B.n112 585
R196 B.n297 B.n296 585
R197 B.n298 B.n111 585
R198 B.n300 B.n299 585
R199 B.n301 B.n110 585
R200 B.n303 B.n302 585
R201 B.n304 B.n109 585
R202 B.n306 B.n305 585
R203 B.n307 B.n108 585
R204 B.n309 B.n308 585
R205 B.n310 B.n107 585
R206 B.n312 B.n311 585
R207 B.n313 B.n106 585
R208 B.n315 B.n314 585
R209 B.n316 B.n105 585
R210 B.n318 B.n317 585
R211 B.n226 B.n139 585
R212 B.n225 B.n224 585
R213 B.n223 B.n140 585
R214 B.n222 B.n221 585
R215 B.n220 B.n141 585
R216 B.n219 B.n218 585
R217 B.n217 B.n142 585
R218 B.n216 B.n215 585
R219 B.n214 B.n143 585
R220 B.n213 B.n212 585
R221 B.n211 B.n144 585
R222 B.n210 B.n209 585
R223 B.n208 B.n145 585
R224 B.n207 B.n206 585
R225 B.n205 B.n146 585
R226 B.n204 B.n203 585
R227 B.n202 B.n147 585
R228 B.n201 B.n200 585
R229 B.n199 B.n148 585
R230 B.n198 B.n197 585
R231 B.n196 B.n149 585
R232 B.n195 B.n194 585
R233 B.n193 B.n150 585
R234 B.n192 B.n191 585
R235 B.n190 B.n151 585
R236 B.n189 B.n188 585
R237 B.n187 B.n152 585
R238 B.n186 B.n185 585
R239 B.n184 B.n153 585
R240 B.n183 B.n182 585
R241 B.n181 B.n154 585
R242 B.n180 B.n179 585
R243 B.n178 B.n155 585
R244 B.n177 B.n176 585
R245 B.n175 B.n156 585
R246 B.n174 B.n173 585
R247 B.n172 B.n157 585
R248 B.n171 B.n170 585
R249 B.n169 B.n158 585
R250 B.n168 B.n167 585
R251 B.n166 B.n159 585
R252 B.n165 B.n164 585
R253 B.n163 B.n160 585
R254 B.n162 B.n161 585
R255 B.n2 B.n0 585
R256 B.n613 B.n1 585
R257 B.n612 B.n611 585
R258 B.n610 B.n3 585
R259 B.n609 B.n608 585
R260 B.n607 B.n4 585
R261 B.n606 B.n605 585
R262 B.n604 B.n5 585
R263 B.n603 B.n602 585
R264 B.n601 B.n6 585
R265 B.n600 B.n599 585
R266 B.n598 B.n7 585
R267 B.n597 B.n596 585
R268 B.n595 B.n8 585
R269 B.n594 B.n593 585
R270 B.n592 B.n9 585
R271 B.n591 B.n590 585
R272 B.n589 B.n10 585
R273 B.n588 B.n587 585
R274 B.n586 B.n11 585
R275 B.n585 B.n584 585
R276 B.n583 B.n12 585
R277 B.n582 B.n581 585
R278 B.n580 B.n13 585
R279 B.n579 B.n578 585
R280 B.n577 B.n14 585
R281 B.n576 B.n575 585
R282 B.n574 B.n15 585
R283 B.n573 B.n572 585
R284 B.n571 B.n16 585
R285 B.n570 B.n569 585
R286 B.n568 B.n17 585
R287 B.n567 B.n566 585
R288 B.n565 B.n18 585
R289 B.n564 B.n563 585
R290 B.n562 B.n19 585
R291 B.n561 B.n560 585
R292 B.n559 B.n20 585
R293 B.n558 B.n557 585
R294 B.n556 B.n21 585
R295 B.n555 B.n554 585
R296 B.n553 B.n22 585
R297 B.n552 B.n551 585
R298 B.n550 B.n23 585
R299 B.n549 B.n548 585
R300 B.n547 B.n24 585
R301 B.n615 B.n614 585
R302 B.n228 B.n139 530.939
R303 B.n547 B.n546 530.939
R304 B.n319 B.n318 530.939
R305 B.n456 B.n59 530.939
R306 B.n118 B.t8 357.568
R307 B.n44 B.t10 357.568
R308 B.n124 B.t5 357.568
R309 B.n38 B.t1 357.568
R310 B.n119 B.t7 276.502
R311 B.n45 B.t11 276.502
R312 B.n125 B.t4 276.502
R313 B.n39 B.t2 276.502
R314 B.n118 B.t6 250.007
R315 B.n124 B.t3 250.007
R316 B.n38 B.t0 250.007
R317 B.n44 B.t9 250.007
R318 B.n224 B.n139 163.367
R319 B.n224 B.n223 163.367
R320 B.n223 B.n222 163.367
R321 B.n222 B.n141 163.367
R322 B.n218 B.n141 163.367
R323 B.n218 B.n217 163.367
R324 B.n217 B.n216 163.367
R325 B.n216 B.n143 163.367
R326 B.n212 B.n143 163.367
R327 B.n212 B.n211 163.367
R328 B.n211 B.n210 163.367
R329 B.n210 B.n145 163.367
R330 B.n206 B.n145 163.367
R331 B.n206 B.n205 163.367
R332 B.n205 B.n204 163.367
R333 B.n204 B.n147 163.367
R334 B.n200 B.n147 163.367
R335 B.n200 B.n199 163.367
R336 B.n199 B.n198 163.367
R337 B.n198 B.n149 163.367
R338 B.n194 B.n149 163.367
R339 B.n194 B.n193 163.367
R340 B.n193 B.n192 163.367
R341 B.n192 B.n151 163.367
R342 B.n188 B.n151 163.367
R343 B.n188 B.n187 163.367
R344 B.n187 B.n186 163.367
R345 B.n186 B.n153 163.367
R346 B.n182 B.n153 163.367
R347 B.n182 B.n181 163.367
R348 B.n181 B.n180 163.367
R349 B.n180 B.n155 163.367
R350 B.n176 B.n155 163.367
R351 B.n176 B.n175 163.367
R352 B.n175 B.n174 163.367
R353 B.n174 B.n157 163.367
R354 B.n170 B.n157 163.367
R355 B.n170 B.n169 163.367
R356 B.n169 B.n168 163.367
R357 B.n168 B.n159 163.367
R358 B.n164 B.n159 163.367
R359 B.n164 B.n163 163.367
R360 B.n163 B.n162 163.367
R361 B.n162 B.n2 163.367
R362 B.n614 B.n2 163.367
R363 B.n614 B.n613 163.367
R364 B.n613 B.n612 163.367
R365 B.n612 B.n3 163.367
R366 B.n608 B.n3 163.367
R367 B.n608 B.n607 163.367
R368 B.n607 B.n606 163.367
R369 B.n606 B.n5 163.367
R370 B.n602 B.n5 163.367
R371 B.n602 B.n601 163.367
R372 B.n601 B.n600 163.367
R373 B.n600 B.n7 163.367
R374 B.n596 B.n7 163.367
R375 B.n596 B.n595 163.367
R376 B.n595 B.n594 163.367
R377 B.n594 B.n9 163.367
R378 B.n590 B.n9 163.367
R379 B.n590 B.n589 163.367
R380 B.n589 B.n588 163.367
R381 B.n588 B.n11 163.367
R382 B.n584 B.n11 163.367
R383 B.n584 B.n583 163.367
R384 B.n583 B.n582 163.367
R385 B.n582 B.n13 163.367
R386 B.n578 B.n13 163.367
R387 B.n578 B.n577 163.367
R388 B.n577 B.n576 163.367
R389 B.n576 B.n15 163.367
R390 B.n572 B.n15 163.367
R391 B.n572 B.n571 163.367
R392 B.n571 B.n570 163.367
R393 B.n570 B.n17 163.367
R394 B.n566 B.n17 163.367
R395 B.n566 B.n565 163.367
R396 B.n565 B.n564 163.367
R397 B.n564 B.n19 163.367
R398 B.n560 B.n19 163.367
R399 B.n560 B.n559 163.367
R400 B.n559 B.n558 163.367
R401 B.n558 B.n21 163.367
R402 B.n554 B.n21 163.367
R403 B.n554 B.n553 163.367
R404 B.n553 B.n552 163.367
R405 B.n552 B.n23 163.367
R406 B.n548 B.n23 163.367
R407 B.n548 B.n547 163.367
R408 B.n229 B.n228 163.367
R409 B.n230 B.n229 163.367
R410 B.n230 B.n137 163.367
R411 B.n234 B.n137 163.367
R412 B.n235 B.n234 163.367
R413 B.n236 B.n235 163.367
R414 B.n236 B.n135 163.367
R415 B.n240 B.n135 163.367
R416 B.n241 B.n240 163.367
R417 B.n242 B.n241 163.367
R418 B.n242 B.n133 163.367
R419 B.n246 B.n133 163.367
R420 B.n247 B.n246 163.367
R421 B.n248 B.n247 163.367
R422 B.n248 B.n131 163.367
R423 B.n252 B.n131 163.367
R424 B.n253 B.n252 163.367
R425 B.n254 B.n253 163.367
R426 B.n254 B.n129 163.367
R427 B.n258 B.n129 163.367
R428 B.n259 B.n258 163.367
R429 B.n260 B.n259 163.367
R430 B.n260 B.n127 163.367
R431 B.n264 B.n127 163.367
R432 B.n265 B.n264 163.367
R433 B.n265 B.n123 163.367
R434 B.n269 B.n123 163.367
R435 B.n270 B.n269 163.367
R436 B.n271 B.n270 163.367
R437 B.n271 B.n121 163.367
R438 B.n275 B.n121 163.367
R439 B.n276 B.n275 163.367
R440 B.n277 B.n276 163.367
R441 B.n277 B.n117 163.367
R442 B.n282 B.n117 163.367
R443 B.n283 B.n282 163.367
R444 B.n284 B.n283 163.367
R445 B.n284 B.n115 163.367
R446 B.n288 B.n115 163.367
R447 B.n289 B.n288 163.367
R448 B.n290 B.n289 163.367
R449 B.n290 B.n113 163.367
R450 B.n294 B.n113 163.367
R451 B.n295 B.n294 163.367
R452 B.n296 B.n295 163.367
R453 B.n296 B.n111 163.367
R454 B.n300 B.n111 163.367
R455 B.n301 B.n300 163.367
R456 B.n302 B.n301 163.367
R457 B.n302 B.n109 163.367
R458 B.n306 B.n109 163.367
R459 B.n307 B.n306 163.367
R460 B.n308 B.n307 163.367
R461 B.n308 B.n107 163.367
R462 B.n312 B.n107 163.367
R463 B.n313 B.n312 163.367
R464 B.n314 B.n313 163.367
R465 B.n314 B.n105 163.367
R466 B.n318 B.n105 163.367
R467 B.n320 B.n319 163.367
R468 B.n320 B.n103 163.367
R469 B.n324 B.n103 163.367
R470 B.n325 B.n324 163.367
R471 B.n326 B.n325 163.367
R472 B.n326 B.n101 163.367
R473 B.n330 B.n101 163.367
R474 B.n331 B.n330 163.367
R475 B.n332 B.n331 163.367
R476 B.n332 B.n99 163.367
R477 B.n336 B.n99 163.367
R478 B.n337 B.n336 163.367
R479 B.n338 B.n337 163.367
R480 B.n338 B.n97 163.367
R481 B.n342 B.n97 163.367
R482 B.n343 B.n342 163.367
R483 B.n344 B.n343 163.367
R484 B.n344 B.n95 163.367
R485 B.n348 B.n95 163.367
R486 B.n349 B.n348 163.367
R487 B.n350 B.n349 163.367
R488 B.n350 B.n93 163.367
R489 B.n354 B.n93 163.367
R490 B.n355 B.n354 163.367
R491 B.n356 B.n355 163.367
R492 B.n356 B.n91 163.367
R493 B.n360 B.n91 163.367
R494 B.n361 B.n360 163.367
R495 B.n362 B.n361 163.367
R496 B.n362 B.n89 163.367
R497 B.n366 B.n89 163.367
R498 B.n367 B.n366 163.367
R499 B.n368 B.n367 163.367
R500 B.n368 B.n87 163.367
R501 B.n372 B.n87 163.367
R502 B.n373 B.n372 163.367
R503 B.n374 B.n373 163.367
R504 B.n374 B.n85 163.367
R505 B.n378 B.n85 163.367
R506 B.n379 B.n378 163.367
R507 B.n380 B.n379 163.367
R508 B.n380 B.n83 163.367
R509 B.n384 B.n83 163.367
R510 B.n385 B.n384 163.367
R511 B.n386 B.n385 163.367
R512 B.n386 B.n81 163.367
R513 B.n390 B.n81 163.367
R514 B.n391 B.n390 163.367
R515 B.n392 B.n391 163.367
R516 B.n392 B.n79 163.367
R517 B.n396 B.n79 163.367
R518 B.n397 B.n396 163.367
R519 B.n398 B.n397 163.367
R520 B.n398 B.n77 163.367
R521 B.n402 B.n77 163.367
R522 B.n403 B.n402 163.367
R523 B.n404 B.n403 163.367
R524 B.n404 B.n75 163.367
R525 B.n408 B.n75 163.367
R526 B.n409 B.n408 163.367
R527 B.n410 B.n409 163.367
R528 B.n410 B.n73 163.367
R529 B.n414 B.n73 163.367
R530 B.n415 B.n414 163.367
R531 B.n416 B.n415 163.367
R532 B.n416 B.n71 163.367
R533 B.n420 B.n71 163.367
R534 B.n421 B.n420 163.367
R535 B.n422 B.n421 163.367
R536 B.n422 B.n69 163.367
R537 B.n426 B.n69 163.367
R538 B.n427 B.n426 163.367
R539 B.n428 B.n427 163.367
R540 B.n428 B.n67 163.367
R541 B.n432 B.n67 163.367
R542 B.n433 B.n432 163.367
R543 B.n434 B.n433 163.367
R544 B.n434 B.n65 163.367
R545 B.n438 B.n65 163.367
R546 B.n439 B.n438 163.367
R547 B.n440 B.n439 163.367
R548 B.n440 B.n63 163.367
R549 B.n444 B.n63 163.367
R550 B.n445 B.n444 163.367
R551 B.n446 B.n445 163.367
R552 B.n446 B.n61 163.367
R553 B.n450 B.n61 163.367
R554 B.n451 B.n450 163.367
R555 B.n452 B.n451 163.367
R556 B.n452 B.n59 163.367
R557 B.n546 B.n25 163.367
R558 B.n542 B.n25 163.367
R559 B.n542 B.n541 163.367
R560 B.n541 B.n540 163.367
R561 B.n540 B.n27 163.367
R562 B.n536 B.n27 163.367
R563 B.n536 B.n535 163.367
R564 B.n535 B.n534 163.367
R565 B.n534 B.n29 163.367
R566 B.n530 B.n29 163.367
R567 B.n530 B.n529 163.367
R568 B.n529 B.n528 163.367
R569 B.n528 B.n31 163.367
R570 B.n524 B.n31 163.367
R571 B.n524 B.n523 163.367
R572 B.n523 B.n522 163.367
R573 B.n522 B.n33 163.367
R574 B.n518 B.n33 163.367
R575 B.n518 B.n517 163.367
R576 B.n517 B.n516 163.367
R577 B.n516 B.n35 163.367
R578 B.n512 B.n35 163.367
R579 B.n512 B.n511 163.367
R580 B.n511 B.n510 163.367
R581 B.n510 B.n37 163.367
R582 B.n505 B.n37 163.367
R583 B.n505 B.n504 163.367
R584 B.n504 B.n503 163.367
R585 B.n503 B.n41 163.367
R586 B.n499 B.n41 163.367
R587 B.n499 B.n498 163.367
R588 B.n498 B.n497 163.367
R589 B.n497 B.n43 163.367
R590 B.n493 B.n43 163.367
R591 B.n493 B.n492 163.367
R592 B.n492 B.n47 163.367
R593 B.n488 B.n47 163.367
R594 B.n488 B.n487 163.367
R595 B.n487 B.n486 163.367
R596 B.n486 B.n49 163.367
R597 B.n482 B.n49 163.367
R598 B.n482 B.n481 163.367
R599 B.n481 B.n480 163.367
R600 B.n480 B.n51 163.367
R601 B.n476 B.n51 163.367
R602 B.n476 B.n475 163.367
R603 B.n475 B.n474 163.367
R604 B.n474 B.n53 163.367
R605 B.n470 B.n53 163.367
R606 B.n470 B.n469 163.367
R607 B.n469 B.n468 163.367
R608 B.n468 B.n55 163.367
R609 B.n464 B.n55 163.367
R610 B.n464 B.n463 163.367
R611 B.n463 B.n462 163.367
R612 B.n462 B.n57 163.367
R613 B.n458 B.n57 163.367
R614 B.n458 B.n457 163.367
R615 B.n457 B.n456 163.367
R616 B.n119 B.n118 81.0672
R617 B.n125 B.n124 81.0672
R618 B.n39 B.n38 81.0672
R619 B.n45 B.n44 81.0672
R620 B.n280 B.n119 59.5399
R621 B.n126 B.n125 59.5399
R622 B.n508 B.n39 59.5399
R623 B.n46 B.n45 59.5399
R624 B.n545 B.n24 34.4981
R625 B.n455 B.n454 34.4981
R626 B.n317 B.n104 34.4981
R627 B.n227 B.n226 34.4981
R628 B B.n615 18.0485
R629 B.n545 B.n544 10.6151
R630 B.n544 B.n543 10.6151
R631 B.n543 B.n26 10.6151
R632 B.n539 B.n26 10.6151
R633 B.n539 B.n538 10.6151
R634 B.n538 B.n537 10.6151
R635 B.n537 B.n28 10.6151
R636 B.n533 B.n28 10.6151
R637 B.n533 B.n532 10.6151
R638 B.n532 B.n531 10.6151
R639 B.n531 B.n30 10.6151
R640 B.n527 B.n30 10.6151
R641 B.n527 B.n526 10.6151
R642 B.n526 B.n525 10.6151
R643 B.n525 B.n32 10.6151
R644 B.n521 B.n32 10.6151
R645 B.n521 B.n520 10.6151
R646 B.n520 B.n519 10.6151
R647 B.n519 B.n34 10.6151
R648 B.n515 B.n34 10.6151
R649 B.n515 B.n514 10.6151
R650 B.n514 B.n513 10.6151
R651 B.n513 B.n36 10.6151
R652 B.n509 B.n36 10.6151
R653 B.n507 B.n506 10.6151
R654 B.n506 B.n40 10.6151
R655 B.n502 B.n40 10.6151
R656 B.n502 B.n501 10.6151
R657 B.n501 B.n500 10.6151
R658 B.n500 B.n42 10.6151
R659 B.n496 B.n42 10.6151
R660 B.n496 B.n495 10.6151
R661 B.n495 B.n494 10.6151
R662 B.n491 B.n490 10.6151
R663 B.n490 B.n489 10.6151
R664 B.n489 B.n48 10.6151
R665 B.n485 B.n48 10.6151
R666 B.n485 B.n484 10.6151
R667 B.n484 B.n483 10.6151
R668 B.n483 B.n50 10.6151
R669 B.n479 B.n50 10.6151
R670 B.n479 B.n478 10.6151
R671 B.n478 B.n477 10.6151
R672 B.n477 B.n52 10.6151
R673 B.n473 B.n52 10.6151
R674 B.n473 B.n472 10.6151
R675 B.n472 B.n471 10.6151
R676 B.n471 B.n54 10.6151
R677 B.n467 B.n54 10.6151
R678 B.n467 B.n466 10.6151
R679 B.n466 B.n465 10.6151
R680 B.n465 B.n56 10.6151
R681 B.n461 B.n56 10.6151
R682 B.n461 B.n460 10.6151
R683 B.n460 B.n459 10.6151
R684 B.n459 B.n58 10.6151
R685 B.n455 B.n58 10.6151
R686 B.n321 B.n104 10.6151
R687 B.n322 B.n321 10.6151
R688 B.n323 B.n322 10.6151
R689 B.n323 B.n102 10.6151
R690 B.n327 B.n102 10.6151
R691 B.n328 B.n327 10.6151
R692 B.n329 B.n328 10.6151
R693 B.n329 B.n100 10.6151
R694 B.n333 B.n100 10.6151
R695 B.n334 B.n333 10.6151
R696 B.n335 B.n334 10.6151
R697 B.n335 B.n98 10.6151
R698 B.n339 B.n98 10.6151
R699 B.n340 B.n339 10.6151
R700 B.n341 B.n340 10.6151
R701 B.n341 B.n96 10.6151
R702 B.n345 B.n96 10.6151
R703 B.n346 B.n345 10.6151
R704 B.n347 B.n346 10.6151
R705 B.n347 B.n94 10.6151
R706 B.n351 B.n94 10.6151
R707 B.n352 B.n351 10.6151
R708 B.n353 B.n352 10.6151
R709 B.n353 B.n92 10.6151
R710 B.n357 B.n92 10.6151
R711 B.n358 B.n357 10.6151
R712 B.n359 B.n358 10.6151
R713 B.n359 B.n90 10.6151
R714 B.n363 B.n90 10.6151
R715 B.n364 B.n363 10.6151
R716 B.n365 B.n364 10.6151
R717 B.n365 B.n88 10.6151
R718 B.n369 B.n88 10.6151
R719 B.n370 B.n369 10.6151
R720 B.n371 B.n370 10.6151
R721 B.n371 B.n86 10.6151
R722 B.n375 B.n86 10.6151
R723 B.n376 B.n375 10.6151
R724 B.n377 B.n376 10.6151
R725 B.n377 B.n84 10.6151
R726 B.n381 B.n84 10.6151
R727 B.n382 B.n381 10.6151
R728 B.n383 B.n382 10.6151
R729 B.n383 B.n82 10.6151
R730 B.n387 B.n82 10.6151
R731 B.n388 B.n387 10.6151
R732 B.n389 B.n388 10.6151
R733 B.n389 B.n80 10.6151
R734 B.n393 B.n80 10.6151
R735 B.n394 B.n393 10.6151
R736 B.n395 B.n394 10.6151
R737 B.n395 B.n78 10.6151
R738 B.n399 B.n78 10.6151
R739 B.n400 B.n399 10.6151
R740 B.n401 B.n400 10.6151
R741 B.n401 B.n76 10.6151
R742 B.n405 B.n76 10.6151
R743 B.n406 B.n405 10.6151
R744 B.n407 B.n406 10.6151
R745 B.n407 B.n74 10.6151
R746 B.n411 B.n74 10.6151
R747 B.n412 B.n411 10.6151
R748 B.n413 B.n412 10.6151
R749 B.n413 B.n72 10.6151
R750 B.n417 B.n72 10.6151
R751 B.n418 B.n417 10.6151
R752 B.n419 B.n418 10.6151
R753 B.n419 B.n70 10.6151
R754 B.n423 B.n70 10.6151
R755 B.n424 B.n423 10.6151
R756 B.n425 B.n424 10.6151
R757 B.n425 B.n68 10.6151
R758 B.n429 B.n68 10.6151
R759 B.n430 B.n429 10.6151
R760 B.n431 B.n430 10.6151
R761 B.n431 B.n66 10.6151
R762 B.n435 B.n66 10.6151
R763 B.n436 B.n435 10.6151
R764 B.n437 B.n436 10.6151
R765 B.n437 B.n64 10.6151
R766 B.n441 B.n64 10.6151
R767 B.n442 B.n441 10.6151
R768 B.n443 B.n442 10.6151
R769 B.n443 B.n62 10.6151
R770 B.n447 B.n62 10.6151
R771 B.n448 B.n447 10.6151
R772 B.n449 B.n448 10.6151
R773 B.n449 B.n60 10.6151
R774 B.n453 B.n60 10.6151
R775 B.n454 B.n453 10.6151
R776 B.n227 B.n138 10.6151
R777 B.n231 B.n138 10.6151
R778 B.n232 B.n231 10.6151
R779 B.n233 B.n232 10.6151
R780 B.n233 B.n136 10.6151
R781 B.n237 B.n136 10.6151
R782 B.n238 B.n237 10.6151
R783 B.n239 B.n238 10.6151
R784 B.n239 B.n134 10.6151
R785 B.n243 B.n134 10.6151
R786 B.n244 B.n243 10.6151
R787 B.n245 B.n244 10.6151
R788 B.n245 B.n132 10.6151
R789 B.n249 B.n132 10.6151
R790 B.n250 B.n249 10.6151
R791 B.n251 B.n250 10.6151
R792 B.n251 B.n130 10.6151
R793 B.n255 B.n130 10.6151
R794 B.n256 B.n255 10.6151
R795 B.n257 B.n256 10.6151
R796 B.n257 B.n128 10.6151
R797 B.n261 B.n128 10.6151
R798 B.n262 B.n261 10.6151
R799 B.n263 B.n262 10.6151
R800 B.n267 B.n266 10.6151
R801 B.n268 B.n267 10.6151
R802 B.n268 B.n122 10.6151
R803 B.n272 B.n122 10.6151
R804 B.n273 B.n272 10.6151
R805 B.n274 B.n273 10.6151
R806 B.n274 B.n120 10.6151
R807 B.n278 B.n120 10.6151
R808 B.n279 B.n278 10.6151
R809 B.n281 B.n116 10.6151
R810 B.n285 B.n116 10.6151
R811 B.n286 B.n285 10.6151
R812 B.n287 B.n286 10.6151
R813 B.n287 B.n114 10.6151
R814 B.n291 B.n114 10.6151
R815 B.n292 B.n291 10.6151
R816 B.n293 B.n292 10.6151
R817 B.n293 B.n112 10.6151
R818 B.n297 B.n112 10.6151
R819 B.n298 B.n297 10.6151
R820 B.n299 B.n298 10.6151
R821 B.n299 B.n110 10.6151
R822 B.n303 B.n110 10.6151
R823 B.n304 B.n303 10.6151
R824 B.n305 B.n304 10.6151
R825 B.n305 B.n108 10.6151
R826 B.n309 B.n108 10.6151
R827 B.n310 B.n309 10.6151
R828 B.n311 B.n310 10.6151
R829 B.n311 B.n106 10.6151
R830 B.n315 B.n106 10.6151
R831 B.n316 B.n315 10.6151
R832 B.n317 B.n316 10.6151
R833 B.n226 B.n225 10.6151
R834 B.n225 B.n140 10.6151
R835 B.n221 B.n140 10.6151
R836 B.n221 B.n220 10.6151
R837 B.n220 B.n219 10.6151
R838 B.n219 B.n142 10.6151
R839 B.n215 B.n142 10.6151
R840 B.n215 B.n214 10.6151
R841 B.n214 B.n213 10.6151
R842 B.n213 B.n144 10.6151
R843 B.n209 B.n144 10.6151
R844 B.n209 B.n208 10.6151
R845 B.n208 B.n207 10.6151
R846 B.n207 B.n146 10.6151
R847 B.n203 B.n146 10.6151
R848 B.n203 B.n202 10.6151
R849 B.n202 B.n201 10.6151
R850 B.n201 B.n148 10.6151
R851 B.n197 B.n148 10.6151
R852 B.n197 B.n196 10.6151
R853 B.n196 B.n195 10.6151
R854 B.n195 B.n150 10.6151
R855 B.n191 B.n150 10.6151
R856 B.n191 B.n190 10.6151
R857 B.n190 B.n189 10.6151
R858 B.n189 B.n152 10.6151
R859 B.n185 B.n152 10.6151
R860 B.n185 B.n184 10.6151
R861 B.n184 B.n183 10.6151
R862 B.n183 B.n154 10.6151
R863 B.n179 B.n154 10.6151
R864 B.n179 B.n178 10.6151
R865 B.n178 B.n177 10.6151
R866 B.n177 B.n156 10.6151
R867 B.n173 B.n156 10.6151
R868 B.n173 B.n172 10.6151
R869 B.n172 B.n171 10.6151
R870 B.n171 B.n158 10.6151
R871 B.n167 B.n158 10.6151
R872 B.n167 B.n166 10.6151
R873 B.n166 B.n165 10.6151
R874 B.n165 B.n160 10.6151
R875 B.n161 B.n160 10.6151
R876 B.n161 B.n0 10.6151
R877 B.n611 B.n1 10.6151
R878 B.n611 B.n610 10.6151
R879 B.n610 B.n609 10.6151
R880 B.n609 B.n4 10.6151
R881 B.n605 B.n4 10.6151
R882 B.n605 B.n604 10.6151
R883 B.n604 B.n603 10.6151
R884 B.n603 B.n6 10.6151
R885 B.n599 B.n6 10.6151
R886 B.n599 B.n598 10.6151
R887 B.n598 B.n597 10.6151
R888 B.n597 B.n8 10.6151
R889 B.n593 B.n8 10.6151
R890 B.n593 B.n592 10.6151
R891 B.n592 B.n591 10.6151
R892 B.n591 B.n10 10.6151
R893 B.n587 B.n10 10.6151
R894 B.n587 B.n586 10.6151
R895 B.n586 B.n585 10.6151
R896 B.n585 B.n12 10.6151
R897 B.n581 B.n12 10.6151
R898 B.n581 B.n580 10.6151
R899 B.n580 B.n579 10.6151
R900 B.n579 B.n14 10.6151
R901 B.n575 B.n14 10.6151
R902 B.n575 B.n574 10.6151
R903 B.n574 B.n573 10.6151
R904 B.n573 B.n16 10.6151
R905 B.n569 B.n16 10.6151
R906 B.n569 B.n568 10.6151
R907 B.n568 B.n567 10.6151
R908 B.n567 B.n18 10.6151
R909 B.n563 B.n18 10.6151
R910 B.n563 B.n562 10.6151
R911 B.n562 B.n561 10.6151
R912 B.n561 B.n20 10.6151
R913 B.n557 B.n20 10.6151
R914 B.n557 B.n556 10.6151
R915 B.n556 B.n555 10.6151
R916 B.n555 B.n22 10.6151
R917 B.n551 B.n22 10.6151
R918 B.n551 B.n550 10.6151
R919 B.n550 B.n549 10.6151
R920 B.n549 B.n24 10.6151
R921 B.n509 B.n508 9.36635
R922 B.n491 B.n46 9.36635
R923 B.n263 B.n126 9.36635
R924 B.n281 B.n280 9.36635
R925 B.n615 B.n0 2.81026
R926 B.n615 B.n1 2.81026
R927 B.n508 B.n507 1.24928
R928 B.n494 B.n46 1.24928
R929 B.n266 B.n126 1.24928
R930 B.n280 B.n279 1.24928
R931 VP.n21 VP.n20 161.3
R932 VP.n19 VP.n1 161.3
R933 VP.n18 VP.n17 161.3
R934 VP.n16 VP.n2 161.3
R935 VP.n15 VP.n14 161.3
R936 VP.n13 VP.n3 161.3
R937 VP.n12 VP.n11 161.3
R938 VP.n10 VP.n4 161.3
R939 VP.n9 VP.n8 161.3
R940 VP.n7 VP.n6 85.6633
R941 VP.n22 VP.n0 85.6633
R942 VP.n5 VP.t3 74.8689
R943 VP.n5 VP.t2 73.5067
R944 VP.n6 VP.n5 47.8773
R945 VP.n7 VP.t0 40.6262
R946 VP.n0 VP.t1 40.6262
R947 VP.n14 VP.n13 40.4934
R948 VP.n14 VP.n2 40.4934
R949 VP.n8 VP.n4 24.4675
R950 VP.n12 VP.n4 24.4675
R951 VP.n13 VP.n12 24.4675
R952 VP.n18 VP.n2 24.4675
R953 VP.n19 VP.n18 24.4675
R954 VP.n20 VP.n19 24.4675
R955 VP.n8 VP.n7 4.40456
R956 VP.n20 VP.n0 4.40456
R957 VP.n9 VP.n6 0.354971
R958 VP.n22 VP.n21 0.354971
R959 VP VP.n22 0.26696
R960 VP.n10 VP.n9 0.189894
R961 VP.n11 VP.n10 0.189894
R962 VP.n11 VP.n3 0.189894
R963 VP.n15 VP.n3 0.189894
R964 VP.n16 VP.n15 0.189894
R965 VP.n17 VP.n16 0.189894
R966 VP.n17 VP.n1 0.189894
R967 VP.n21 VP.n1 0.189894
R968 VDD1 VDD1.n1 131.022
R969 VDD1 VDD1.n0 90.4345
R970 VDD1.n0 VDD1.t1 5.00897
R971 VDD1.n0 VDD1.t0 5.00897
R972 VDD1.n1 VDD1.t2 5.00897
R973 VDD1.n1 VDD1.t3 5.00897
R974 VTAIL.n270 VTAIL.n269 756.745
R975 VTAIL.n32 VTAIL.n31 756.745
R976 VTAIL.n66 VTAIL.n65 756.745
R977 VTAIL.n100 VTAIL.n99 756.745
R978 VTAIL.n236 VTAIL.n235 756.745
R979 VTAIL.n202 VTAIL.n201 756.745
R980 VTAIL.n168 VTAIL.n167 756.745
R981 VTAIL.n134 VTAIL.n133 756.745
R982 VTAIL.n248 VTAIL.n247 585
R983 VTAIL.n253 VTAIL.n252 585
R984 VTAIL.n255 VTAIL.n254 585
R985 VTAIL.n244 VTAIL.n243 585
R986 VTAIL.n261 VTAIL.n260 585
R987 VTAIL.n263 VTAIL.n262 585
R988 VTAIL.n240 VTAIL.n239 585
R989 VTAIL.n269 VTAIL.n268 585
R990 VTAIL.n10 VTAIL.n9 585
R991 VTAIL.n15 VTAIL.n14 585
R992 VTAIL.n17 VTAIL.n16 585
R993 VTAIL.n6 VTAIL.n5 585
R994 VTAIL.n23 VTAIL.n22 585
R995 VTAIL.n25 VTAIL.n24 585
R996 VTAIL.n2 VTAIL.n1 585
R997 VTAIL.n31 VTAIL.n30 585
R998 VTAIL.n44 VTAIL.n43 585
R999 VTAIL.n49 VTAIL.n48 585
R1000 VTAIL.n51 VTAIL.n50 585
R1001 VTAIL.n40 VTAIL.n39 585
R1002 VTAIL.n57 VTAIL.n56 585
R1003 VTAIL.n59 VTAIL.n58 585
R1004 VTAIL.n36 VTAIL.n35 585
R1005 VTAIL.n65 VTAIL.n64 585
R1006 VTAIL.n78 VTAIL.n77 585
R1007 VTAIL.n83 VTAIL.n82 585
R1008 VTAIL.n85 VTAIL.n84 585
R1009 VTAIL.n74 VTAIL.n73 585
R1010 VTAIL.n91 VTAIL.n90 585
R1011 VTAIL.n93 VTAIL.n92 585
R1012 VTAIL.n70 VTAIL.n69 585
R1013 VTAIL.n99 VTAIL.n98 585
R1014 VTAIL.n235 VTAIL.n234 585
R1015 VTAIL.n206 VTAIL.n205 585
R1016 VTAIL.n229 VTAIL.n228 585
R1017 VTAIL.n227 VTAIL.n226 585
R1018 VTAIL.n210 VTAIL.n209 585
R1019 VTAIL.n221 VTAIL.n220 585
R1020 VTAIL.n219 VTAIL.n218 585
R1021 VTAIL.n214 VTAIL.n213 585
R1022 VTAIL.n201 VTAIL.n200 585
R1023 VTAIL.n172 VTAIL.n171 585
R1024 VTAIL.n195 VTAIL.n194 585
R1025 VTAIL.n193 VTAIL.n192 585
R1026 VTAIL.n176 VTAIL.n175 585
R1027 VTAIL.n187 VTAIL.n186 585
R1028 VTAIL.n185 VTAIL.n184 585
R1029 VTAIL.n180 VTAIL.n179 585
R1030 VTAIL.n167 VTAIL.n166 585
R1031 VTAIL.n138 VTAIL.n137 585
R1032 VTAIL.n161 VTAIL.n160 585
R1033 VTAIL.n159 VTAIL.n158 585
R1034 VTAIL.n142 VTAIL.n141 585
R1035 VTAIL.n153 VTAIL.n152 585
R1036 VTAIL.n151 VTAIL.n150 585
R1037 VTAIL.n146 VTAIL.n145 585
R1038 VTAIL.n133 VTAIL.n132 585
R1039 VTAIL.n104 VTAIL.n103 585
R1040 VTAIL.n127 VTAIL.n126 585
R1041 VTAIL.n125 VTAIL.n124 585
R1042 VTAIL.n108 VTAIL.n107 585
R1043 VTAIL.n119 VTAIL.n118 585
R1044 VTAIL.n117 VTAIL.n116 585
R1045 VTAIL.n112 VTAIL.n111 585
R1046 VTAIL.n249 VTAIL.t1 329.084
R1047 VTAIL.n11 VTAIL.t3 329.084
R1048 VTAIL.n45 VTAIL.t6 329.084
R1049 VTAIL.n79 VTAIL.t7 329.084
R1050 VTAIL.n215 VTAIL.t5 329.084
R1051 VTAIL.n181 VTAIL.t4 329.084
R1052 VTAIL.n147 VTAIL.t2 329.084
R1053 VTAIL.n113 VTAIL.t0 329.084
R1054 VTAIL.n253 VTAIL.n247 171.744
R1055 VTAIL.n254 VTAIL.n253 171.744
R1056 VTAIL.n254 VTAIL.n243 171.744
R1057 VTAIL.n261 VTAIL.n243 171.744
R1058 VTAIL.n262 VTAIL.n261 171.744
R1059 VTAIL.n262 VTAIL.n239 171.744
R1060 VTAIL.n269 VTAIL.n239 171.744
R1061 VTAIL.n15 VTAIL.n9 171.744
R1062 VTAIL.n16 VTAIL.n15 171.744
R1063 VTAIL.n16 VTAIL.n5 171.744
R1064 VTAIL.n23 VTAIL.n5 171.744
R1065 VTAIL.n24 VTAIL.n23 171.744
R1066 VTAIL.n24 VTAIL.n1 171.744
R1067 VTAIL.n31 VTAIL.n1 171.744
R1068 VTAIL.n49 VTAIL.n43 171.744
R1069 VTAIL.n50 VTAIL.n49 171.744
R1070 VTAIL.n50 VTAIL.n39 171.744
R1071 VTAIL.n57 VTAIL.n39 171.744
R1072 VTAIL.n58 VTAIL.n57 171.744
R1073 VTAIL.n58 VTAIL.n35 171.744
R1074 VTAIL.n65 VTAIL.n35 171.744
R1075 VTAIL.n83 VTAIL.n77 171.744
R1076 VTAIL.n84 VTAIL.n83 171.744
R1077 VTAIL.n84 VTAIL.n73 171.744
R1078 VTAIL.n91 VTAIL.n73 171.744
R1079 VTAIL.n92 VTAIL.n91 171.744
R1080 VTAIL.n92 VTAIL.n69 171.744
R1081 VTAIL.n99 VTAIL.n69 171.744
R1082 VTAIL.n235 VTAIL.n205 171.744
R1083 VTAIL.n228 VTAIL.n205 171.744
R1084 VTAIL.n228 VTAIL.n227 171.744
R1085 VTAIL.n227 VTAIL.n209 171.744
R1086 VTAIL.n220 VTAIL.n209 171.744
R1087 VTAIL.n220 VTAIL.n219 171.744
R1088 VTAIL.n219 VTAIL.n213 171.744
R1089 VTAIL.n201 VTAIL.n171 171.744
R1090 VTAIL.n194 VTAIL.n171 171.744
R1091 VTAIL.n194 VTAIL.n193 171.744
R1092 VTAIL.n193 VTAIL.n175 171.744
R1093 VTAIL.n186 VTAIL.n175 171.744
R1094 VTAIL.n186 VTAIL.n185 171.744
R1095 VTAIL.n185 VTAIL.n179 171.744
R1096 VTAIL.n167 VTAIL.n137 171.744
R1097 VTAIL.n160 VTAIL.n137 171.744
R1098 VTAIL.n160 VTAIL.n159 171.744
R1099 VTAIL.n159 VTAIL.n141 171.744
R1100 VTAIL.n152 VTAIL.n141 171.744
R1101 VTAIL.n152 VTAIL.n151 171.744
R1102 VTAIL.n151 VTAIL.n145 171.744
R1103 VTAIL.n133 VTAIL.n103 171.744
R1104 VTAIL.n126 VTAIL.n103 171.744
R1105 VTAIL.n126 VTAIL.n125 171.744
R1106 VTAIL.n125 VTAIL.n107 171.744
R1107 VTAIL.n118 VTAIL.n107 171.744
R1108 VTAIL.n118 VTAIL.n117 171.744
R1109 VTAIL.n117 VTAIL.n111 171.744
R1110 VTAIL.t1 VTAIL.n247 85.8723
R1111 VTAIL.t3 VTAIL.n9 85.8723
R1112 VTAIL.t6 VTAIL.n43 85.8723
R1113 VTAIL.t7 VTAIL.n77 85.8723
R1114 VTAIL.t5 VTAIL.n213 85.8723
R1115 VTAIL.t4 VTAIL.n179 85.8723
R1116 VTAIL.t2 VTAIL.n145 85.8723
R1117 VTAIL.t0 VTAIL.n111 85.8723
R1118 VTAIL.n271 VTAIL.n270 34.3187
R1119 VTAIL.n33 VTAIL.n32 34.3187
R1120 VTAIL.n67 VTAIL.n66 34.3187
R1121 VTAIL.n101 VTAIL.n100 34.3187
R1122 VTAIL.n237 VTAIL.n236 34.3187
R1123 VTAIL.n203 VTAIL.n202 34.3187
R1124 VTAIL.n169 VTAIL.n168 34.3187
R1125 VTAIL.n135 VTAIL.n134 34.3187
R1126 VTAIL.n271 VTAIL.n237 21.5652
R1127 VTAIL.n135 VTAIL.n101 21.5652
R1128 VTAIL.n268 VTAIL.n238 12.8005
R1129 VTAIL.n30 VTAIL.n0 12.8005
R1130 VTAIL.n64 VTAIL.n34 12.8005
R1131 VTAIL.n98 VTAIL.n68 12.8005
R1132 VTAIL.n234 VTAIL.n204 12.8005
R1133 VTAIL.n200 VTAIL.n170 12.8005
R1134 VTAIL.n166 VTAIL.n136 12.8005
R1135 VTAIL.n132 VTAIL.n102 12.8005
R1136 VTAIL.n267 VTAIL.n240 12.0247
R1137 VTAIL.n29 VTAIL.n2 12.0247
R1138 VTAIL.n63 VTAIL.n36 12.0247
R1139 VTAIL.n97 VTAIL.n70 12.0247
R1140 VTAIL.n233 VTAIL.n206 12.0247
R1141 VTAIL.n199 VTAIL.n172 12.0247
R1142 VTAIL.n165 VTAIL.n138 12.0247
R1143 VTAIL.n131 VTAIL.n104 12.0247
R1144 VTAIL.n264 VTAIL.n263 11.249
R1145 VTAIL.n26 VTAIL.n25 11.249
R1146 VTAIL.n60 VTAIL.n59 11.249
R1147 VTAIL.n94 VTAIL.n93 11.249
R1148 VTAIL.n230 VTAIL.n229 11.249
R1149 VTAIL.n196 VTAIL.n195 11.249
R1150 VTAIL.n162 VTAIL.n161 11.249
R1151 VTAIL.n128 VTAIL.n127 11.249
R1152 VTAIL.n249 VTAIL.n248 10.7233
R1153 VTAIL.n11 VTAIL.n10 10.7233
R1154 VTAIL.n45 VTAIL.n44 10.7233
R1155 VTAIL.n79 VTAIL.n78 10.7233
R1156 VTAIL.n215 VTAIL.n214 10.7233
R1157 VTAIL.n181 VTAIL.n180 10.7233
R1158 VTAIL.n147 VTAIL.n146 10.7233
R1159 VTAIL.n113 VTAIL.n112 10.7233
R1160 VTAIL.n260 VTAIL.n242 10.4732
R1161 VTAIL.n22 VTAIL.n4 10.4732
R1162 VTAIL.n56 VTAIL.n38 10.4732
R1163 VTAIL.n90 VTAIL.n72 10.4732
R1164 VTAIL.n226 VTAIL.n208 10.4732
R1165 VTAIL.n192 VTAIL.n174 10.4732
R1166 VTAIL.n158 VTAIL.n140 10.4732
R1167 VTAIL.n124 VTAIL.n106 10.4732
R1168 VTAIL.n259 VTAIL.n244 9.69747
R1169 VTAIL.n21 VTAIL.n6 9.69747
R1170 VTAIL.n55 VTAIL.n40 9.69747
R1171 VTAIL.n89 VTAIL.n74 9.69747
R1172 VTAIL.n225 VTAIL.n210 9.69747
R1173 VTAIL.n191 VTAIL.n176 9.69747
R1174 VTAIL.n157 VTAIL.n142 9.69747
R1175 VTAIL.n123 VTAIL.n108 9.69747
R1176 VTAIL.n266 VTAIL.n238 9.45567
R1177 VTAIL.n28 VTAIL.n0 9.45567
R1178 VTAIL.n62 VTAIL.n34 9.45567
R1179 VTAIL.n96 VTAIL.n68 9.45567
R1180 VTAIL.n232 VTAIL.n204 9.45567
R1181 VTAIL.n198 VTAIL.n170 9.45567
R1182 VTAIL.n164 VTAIL.n136 9.45567
R1183 VTAIL.n130 VTAIL.n102 9.45567
R1184 VTAIL.n251 VTAIL.n250 9.3005
R1185 VTAIL.n246 VTAIL.n245 9.3005
R1186 VTAIL.n257 VTAIL.n256 9.3005
R1187 VTAIL.n259 VTAIL.n258 9.3005
R1188 VTAIL.n242 VTAIL.n241 9.3005
R1189 VTAIL.n265 VTAIL.n264 9.3005
R1190 VTAIL.n267 VTAIL.n266 9.3005
R1191 VTAIL.n13 VTAIL.n12 9.3005
R1192 VTAIL.n8 VTAIL.n7 9.3005
R1193 VTAIL.n19 VTAIL.n18 9.3005
R1194 VTAIL.n21 VTAIL.n20 9.3005
R1195 VTAIL.n4 VTAIL.n3 9.3005
R1196 VTAIL.n27 VTAIL.n26 9.3005
R1197 VTAIL.n29 VTAIL.n28 9.3005
R1198 VTAIL.n47 VTAIL.n46 9.3005
R1199 VTAIL.n42 VTAIL.n41 9.3005
R1200 VTAIL.n53 VTAIL.n52 9.3005
R1201 VTAIL.n55 VTAIL.n54 9.3005
R1202 VTAIL.n38 VTAIL.n37 9.3005
R1203 VTAIL.n61 VTAIL.n60 9.3005
R1204 VTAIL.n63 VTAIL.n62 9.3005
R1205 VTAIL.n81 VTAIL.n80 9.3005
R1206 VTAIL.n76 VTAIL.n75 9.3005
R1207 VTAIL.n87 VTAIL.n86 9.3005
R1208 VTAIL.n89 VTAIL.n88 9.3005
R1209 VTAIL.n72 VTAIL.n71 9.3005
R1210 VTAIL.n95 VTAIL.n94 9.3005
R1211 VTAIL.n97 VTAIL.n96 9.3005
R1212 VTAIL.n233 VTAIL.n232 9.3005
R1213 VTAIL.n231 VTAIL.n230 9.3005
R1214 VTAIL.n208 VTAIL.n207 9.3005
R1215 VTAIL.n225 VTAIL.n224 9.3005
R1216 VTAIL.n223 VTAIL.n222 9.3005
R1217 VTAIL.n212 VTAIL.n211 9.3005
R1218 VTAIL.n217 VTAIL.n216 9.3005
R1219 VTAIL.n178 VTAIL.n177 9.3005
R1220 VTAIL.n189 VTAIL.n188 9.3005
R1221 VTAIL.n191 VTAIL.n190 9.3005
R1222 VTAIL.n174 VTAIL.n173 9.3005
R1223 VTAIL.n197 VTAIL.n196 9.3005
R1224 VTAIL.n199 VTAIL.n198 9.3005
R1225 VTAIL.n183 VTAIL.n182 9.3005
R1226 VTAIL.n144 VTAIL.n143 9.3005
R1227 VTAIL.n155 VTAIL.n154 9.3005
R1228 VTAIL.n157 VTAIL.n156 9.3005
R1229 VTAIL.n140 VTAIL.n139 9.3005
R1230 VTAIL.n163 VTAIL.n162 9.3005
R1231 VTAIL.n165 VTAIL.n164 9.3005
R1232 VTAIL.n149 VTAIL.n148 9.3005
R1233 VTAIL.n110 VTAIL.n109 9.3005
R1234 VTAIL.n121 VTAIL.n120 9.3005
R1235 VTAIL.n123 VTAIL.n122 9.3005
R1236 VTAIL.n106 VTAIL.n105 9.3005
R1237 VTAIL.n129 VTAIL.n128 9.3005
R1238 VTAIL.n131 VTAIL.n130 9.3005
R1239 VTAIL.n115 VTAIL.n114 9.3005
R1240 VTAIL.n256 VTAIL.n255 8.92171
R1241 VTAIL.n18 VTAIL.n17 8.92171
R1242 VTAIL.n52 VTAIL.n51 8.92171
R1243 VTAIL.n86 VTAIL.n85 8.92171
R1244 VTAIL.n222 VTAIL.n221 8.92171
R1245 VTAIL.n188 VTAIL.n187 8.92171
R1246 VTAIL.n154 VTAIL.n153 8.92171
R1247 VTAIL.n120 VTAIL.n119 8.92171
R1248 VTAIL.n252 VTAIL.n246 8.14595
R1249 VTAIL.n14 VTAIL.n8 8.14595
R1250 VTAIL.n48 VTAIL.n42 8.14595
R1251 VTAIL.n82 VTAIL.n76 8.14595
R1252 VTAIL.n218 VTAIL.n212 8.14595
R1253 VTAIL.n184 VTAIL.n178 8.14595
R1254 VTAIL.n150 VTAIL.n144 8.14595
R1255 VTAIL.n116 VTAIL.n110 8.14595
R1256 VTAIL.n251 VTAIL.n248 7.3702
R1257 VTAIL.n13 VTAIL.n10 7.3702
R1258 VTAIL.n47 VTAIL.n44 7.3702
R1259 VTAIL.n81 VTAIL.n78 7.3702
R1260 VTAIL.n217 VTAIL.n214 7.3702
R1261 VTAIL.n183 VTAIL.n180 7.3702
R1262 VTAIL.n149 VTAIL.n146 7.3702
R1263 VTAIL.n115 VTAIL.n112 7.3702
R1264 VTAIL.n252 VTAIL.n251 5.81868
R1265 VTAIL.n14 VTAIL.n13 5.81868
R1266 VTAIL.n48 VTAIL.n47 5.81868
R1267 VTAIL.n82 VTAIL.n81 5.81868
R1268 VTAIL.n218 VTAIL.n217 5.81868
R1269 VTAIL.n184 VTAIL.n183 5.81868
R1270 VTAIL.n150 VTAIL.n149 5.81868
R1271 VTAIL.n116 VTAIL.n115 5.81868
R1272 VTAIL.n255 VTAIL.n246 5.04292
R1273 VTAIL.n17 VTAIL.n8 5.04292
R1274 VTAIL.n51 VTAIL.n42 5.04292
R1275 VTAIL.n85 VTAIL.n76 5.04292
R1276 VTAIL.n221 VTAIL.n212 5.04292
R1277 VTAIL.n187 VTAIL.n178 5.04292
R1278 VTAIL.n153 VTAIL.n144 5.04292
R1279 VTAIL.n119 VTAIL.n110 5.04292
R1280 VTAIL.n256 VTAIL.n244 4.26717
R1281 VTAIL.n18 VTAIL.n6 4.26717
R1282 VTAIL.n52 VTAIL.n40 4.26717
R1283 VTAIL.n86 VTAIL.n74 4.26717
R1284 VTAIL.n222 VTAIL.n210 4.26717
R1285 VTAIL.n188 VTAIL.n176 4.26717
R1286 VTAIL.n154 VTAIL.n142 4.26717
R1287 VTAIL.n120 VTAIL.n108 4.26717
R1288 VTAIL.n169 VTAIL.n135 3.60395
R1289 VTAIL.n237 VTAIL.n203 3.60395
R1290 VTAIL.n101 VTAIL.n67 3.60395
R1291 VTAIL.n260 VTAIL.n259 3.49141
R1292 VTAIL.n22 VTAIL.n21 3.49141
R1293 VTAIL.n56 VTAIL.n55 3.49141
R1294 VTAIL.n90 VTAIL.n89 3.49141
R1295 VTAIL.n226 VTAIL.n225 3.49141
R1296 VTAIL.n192 VTAIL.n191 3.49141
R1297 VTAIL.n158 VTAIL.n157 3.49141
R1298 VTAIL.n124 VTAIL.n123 3.49141
R1299 VTAIL.n263 VTAIL.n242 2.71565
R1300 VTAIL.n25 VTAIL.n4 2.71565
R1301 VTAIL.n59 VTAIL.n38 2.71565
R1302 VTAIL.n93 VTAIL.n72 2.71565
R1303 VTAIL.n229 VTAIL.n208 2.71565
R1304 VTAIL.n195 VTAIL.n174 2.71565
R1305 VTAIL.n161 VTAIL.n140 2.71565
R1306 VTAIL.n127 VTAIL.n106 2.71565
R1307 VTAIL.n182 VTAIL.n181 2.41347
R1308 VTAIL.n148 VTAIL.n147 2.41347
R1309 VTAIL.n114 VTAIL.n113 2.41347
R1310 VTAIL.n250 VTAIL.n249 2.41347
R1311 VTAIL.n12 VTAIL.n11 2.41347
R1312 VTAIL.n46 VTAIL.n45 2.41347
R1313 VTAIL.n80 VTAIL.n79 2.41347
R1314 VTAIL.n216 VTAIL.n215 2.41347
R1315 VTAIL.n264 VTAIL.n240 1.93989
R1316 VTAIL.n26 VTAIL.n2 1.93989
R1317 VTAIL.n60 VTAIL.n36 1.93989
R1318 VTAIL.n94 VTAIL.n70 1.93989
R1319 VTAIL.n230 VTAIL.n206 1.93989
R1320 VTAIL.n196 VTAIL.n172 1.93989
R1321 VTAIL.n162 VTAIL.n138 1.93989
R1322 VTAIL.n128 VTAIL.n104 1.93989
R1323 VTAIL VTAIL.n33 1.86041
R1324 VTAIL VTAIL.n271 1.74403
R1325 VTAIL.n268 VTAIL.n267 1.16414
R1326 VTAIL.n30 VTAIL.n29 1.16414
R1327 VTAIL.n64 VTAIL.n63 1.16414
R1328 VTAIL.n98 VTAIL.n97 1.16414
R1329 VTAIL.n234 VTAIL.n233 1.16414
R1330 VTAIL.n200 VTAIL.n199 1.16414
R1331 VTAIL.n166 VTAIL.n165 1.16414
R1332 VTAIL.n132 VTAIL.n131 1.16414
R1333 VTAIL.n203 VTAIL.n169 0.470328
R1334 VTAIL.n67 VTAIL.n33 0.470328
R1335 VTAIL.n270 VTAIL.n238 0.388379
R1336 VTAIL.n32 VTAIL.n0 0.388379
R1337 VTAIL.n66 VTAIL.n34 0.388379
R1338 VTAIL.n100 VTAIL.n68 0.388379
R1339 VTAIL.n236 VTAIL.n204 0.388379
R1340 VTAIL.n202 VTAIL.n170 0.388379
R1341 VTAIL.n168 VTAIL.n136 0.388379
R1342 VTAIL.n134 VTAIL.n102 0.388379
R1343 VTAIL.n250 VTAIL.n245 0.155672
R1344 VTAIL.n257 VTAIL.n245 0.155672
R1345 VTAIL.n258 VTAIL.n257 0.155672
R1346 VTAIL.n258 VTAIL.n241 0.155672
R1347 VTAIL.n265 VTAIL.n241 0.155672
R1348 VTAIL.n266 VTAIL.n265 0.155672
R1349 VTAIL.n12 VTAIL.n7 0.155672
R1350 VTAIL.n19 VTAIL.n7 0.155672
R1351 VTAIL.n20 VTAIL.n19 0.155672
R1352 VTAIL.n20 VTAIL.n3 0.155672
R1353 VTAIL.n27 VTAIL.n3 0.155672
R1354 VTAIL.n28 VTAIL.n27 0.155672
R1355 VTAIL.n46 VTAIL.n41 0.155672
R1356 VTAIL.n53 VTAIL.n41 0.155672
R1357 VTAIL.n54 VTAIL.n53 0.155672
R1358 VTAIL.n54 VTAIL.n37 0.155672
R1359 VTAIL.n61 VTAIL.n37 0.155672
R1360 VTAIL.n62 VTAIL.n61 0.155672
R1361 VTAIL.n80 VTAIL.n75 0.155672
R1362 VTAIL.n87 VTAIL.n75 0.155672
R1363 VTAIL.n88 VTAIL.n87 0.155672
R1364 VTAIL.n88 VTAIL.n71 0.155672
R1365 VTAIL.n95 VTAIL.n71 0.155672
R1366 VTAIL.n96 VTAIL.n95 0.155672
R1367 VTAIL.n232 VTAIL.n231 0.155672
R1368 VTAIL.n231 VTAIL.n207 0.155672
R1369 VTAIL.n224 VTAIL.n207 0.155672
R1370 VTAIL.n224 VTAIL.n223 0.155672
R1371 VTAIL.n223 VTAIL.n211 0.155672
R1372 VTAIL.n216 VTAIL.n211 0.155672
R1373 VTAIL.n198 VTAIL.n197 0.155672
R1374 VTAIL.n197 VTAIL.n173 0.155672
R1375 VTAIL.n190 VTAIL.n173 0.155672
R1376 VTAIL.n190 VTAIL.n189 0.155672
R1377 VTAIL.n189 VTAIL.n177 0.155672
R1378 VTAIL.n182 VTAIL.n177 0.155672
R1379 VTAIL.n164 VTAIL.n163 0.155672
R1380 VTAIL.n163 VTAIL.n139 0.155672
R1381 VTAIL.n156 VTAIL.n139 0.155672
R1382 VTAIL.n156 VTAIL.n155 0.155672
R1383 VTAIL.n155 VTAIL.n143 0.155672
R1384 VTAIL.n148 VTAIL.n143 0.155672
R1385 VTAIL.n130 VTAIL.n129 0.155672
R1386 VTAIL.n129 VTAIL.n105 0.155672
R1387 VTAIL.n122 VTAIL.n105 0.155672
R1388 VTAIL.n122 VTAIL.n121 0.155672
R1389 VTAIL.n121 VTAIL.n109 0.155672
R1390 VTAIL.n114 VTAIL.n109 0.155672
R1391 VN.n1 VN.t2 74.869
R1392 VN.n0 VN.t3 74.869
R1393 VN.n0 VN.t1 73.5066
R1394 VN.n1 VN.t0 73.5066
R1395 VN VN.n1 48.0426
R1396 VN VN.n0 1.81916
R1397 VDD2.n2 VDD2.n0 130.496
R1398 VDD2.n2 VDD2.n1 90.3763
R1399 VDD2.n1 VDD2.t3 5.00897
R1400 VDD2.n1 VDD2.t1 5.00897
R1401 VDD2.n0 VDD2.t0 5.00897
R1402 VDD2.n0 VDD2.t2 5.00897
R1403 VDD2 VDD2.n2 0.0586897
C0 VN w_n3478_n2266# 6.01784f
C1 w_n3478_n2266# VDD1 1.5358f
C2 VN VDD1 0.149985f
C3 VDD2 B 1.40803f
C4 B VP 2.03058f
C5 B VTAIL 3.52377f
C6 VDD2 VP 0.4737f
C7 VDD2 VTAIL 4.68749f
C8 VTAIL VP 3.40728f
C9 B w_n3478_n2266# 9.247781f
C10 VDD2 w_n3478_n2266# 1.61947f
C11 w_n3478_n2266# VP 6.46811f
C12 B VN 1.27756f
C13 VTAIL w_n3478_n2266# 2.81862f
C14 B VDD1 1.3352f
C15 VDD2 VN 2.88538f
C16 VN VP 6.07032f
C17 VDD2 VDD1 1.3307f
C18 VDD1 VP 3.20804f
C19 VN VTAIL 3.39317f
C20 VTAIL VDD1 4.6249f
C21 VDD2 VSUBS 1.022532f
C22 VDD1 VSUBS 5.80267f
C23 VTAIL VSUBS 0.82318f
C24 VN VSUBS 6.0615f
C25 VP VSUBS 2.583526f
C26 B VSUBS 4.887981f
C27 w_n3478_n2266# VSUBS 98.204796f
C28 VDD2.t0 VSUBS 0.145999f
C29 VDD2.t2 VSUBS 0.145999f
C30 VDD2.n0 VSUBS 1.52786f
C31 VDD2.t3 VSUBS 0.145999f
C32 VDD2.t1 VSUBS 0.145999f
C33 VDD2.n1 VSUBS 1.0076f
C34 VDD2.n2 VSUBS 4.14388f
C35 VN.t1 VSUBS 2.73493f
C36 VN.t3 VSUBS 2.75422f
C37 VN.n0 VSUBS 1.6064f
C38 VN.t0 VSUBS 2.73493f
C39 VN.t2 VSUBS 2.75422f
C40 VN.n1 VSUBS 3.61851f
C41 VTAIL.n0 VSUBS 0.016071f
C42 VTAIL.n1 VSUBS 0.036307f
C43 VTAIL.n2 VSUBS 0.016264f
C44 VTAIL.n3 VSUBS 0.028586f
C45 VTAIL.n4 VSUBS 0.015361f
C46 VTAIL.n5 VSUBS 0.036307f
C47 VTAIL.n6 VSUBS 0.016264f
C48 VTAIL.n7 VSUBS 0.028586f
C49 VTAIL.n8 VSUBS 0.015361f
C50 VTAIL.n9 VSUBS 0.02723f
C51 VTAIL.n10 VSUBS 0.027308f
C52 VTAIL.t3 VSUBS 0.078023f
C53 VTAIL.n11 VSUBS 0.154166f
C54 VTAIL.n12 VSUBS 0.713799f
C55 VTAIL.n13 VSUBS 0.015361f
C56 VTAIL.n14 VSUBS 0.016264f
C57 VTAIL.n15 VSUBS 0.036307f
C58 VTAIL.n16 VSUBS 0.036307f
C59 VTAIL.n17 VSUBS 0.016264f
C60 VTAIL.n18 VSUBS 0.015361f
C61 VTAIL.n19 VSUBS 0.028586f
C62 VTAIL.n20 VSUBS 0.028586f
C63 VTAIL.n21 VSUBS 0.015361f
C64 VTAIL.n22 VSUBS 0.016264f
C65 VTAIL.n23 VSUBS 0.036307f
C66 VTAIL.n24 VSUBS 0.036307f
C67 VTAIL.n25 VSUBS 0.016264f
C68 VTAIL.n26 VSUBS 0.015361f
C69 VTAIL.n27 VSUBS 0.028586f
C70 VTAIL.n28 VSUBS 0.071151f
C71 VTAIL.n29 VSUBS 0.015361f
C72 VTAIL.n30 VSUBS 0.016264f
C73 VTAIL.n31 VSUBS 0.079646f
C74 VTAIL.n32 VSUBS 0.052293f
C75 VTAIL.n33 VSUBS 0.241434f
C76 VTAIL.n34 VSUBS 0.016071f
C77 VTAIL.n35 VSUBS 0.036307f
C78 VTAIL.n36 VSUBS 0.016264f
C79 VTAIL.n37 VSUBS 0.028586f
C80 VTAIL.n38 VSUBS 0.015361f
C81 VTAIL.n39 VSUBS 0.036307f
C82 VTAIL.n40 VSUBS 0.016264f
C83 VTAIL.n41 VSUBS 0.028586f
C84 VTAIL.n42 VSUBS 0.015361f
C85 VTAIL.n43 VSUBS 0.02723f
C86 VTAIL.n44 VSUBS 0.027308f
C87 VTAIL.t6 VSUBS 0.078023f
C88 VTAIL.n45 VSUBS 0.154166f
C89 VTAIL.n46 VSUBS 0.713799f
C90 VTAIL.n47 VSUBS 0.015361f
C91 VTAIL.n48 VSUBS 0.016264f
C92 VTAIL.n49 VSUBS 0.036307f
C93 VTAIL.n50 VSUBS 0.036307f
C94 VTAIL.n51 VSUBS 0.016264f
C95 VTAIL.n52 VSUBS 0.015361f
C96 VTAIL.n53 VSUBS 0.028586f
C97 VTAIL.n54 VSUBS 0.028586f
C98 VTAIL.n55 VSUBS 0.015361f
C99 VTAIL.n56 VSUBS 0.016264f
C100 VTAIL.n57 VSUBS 0.036307f
C101 VTAIL.n58 VSUBS 0.036307f
C102 VTAIL.n59 VSUBS 0.016264f
C103 VTAIL.n60 VSUBS 0.015361f
C104 VTAIL.n61 VSUBS 0.028586f
C105 VTAIL.n62 VSUBS 0.071151f
C106 VTAIL.n63 VSUBS 0.015361f
C107 VTAIL.n64 VSUBS 0.016264f
C108 VTAIL.n65 VSUBS 0.079646f
C109 VTAIL.n66 VSUBS 0.052293f
C110 VTAIL.n67 VSUBS 0.402029f
C111 VTAIL.n68 VSUBS 0.016071f
C112 VTAIL.n69 VSUBS 0.036307f
C113 VTAIL.n70 VSUBS 0.016264f
C114 VTAIL.n71 VSUBS 0.028586f
C115 VTAIL.n72 VSUBS 0.015361f
C116 VTAIL.n73 VSUBS 0.036307f
C117 VTAIL.n74 VSUBS 0.016264f
C118 VTAIL.n75 VSUBS 0.028586f
C119 VTAIL.n76 VSUBS 0.015361f
C120 VTAIL.n77 VSUBS 0.02723f
C121 VTAIL.n78 VSUBS 0.027308f
C122 VTAIL.t7 VSUBS 0.078023f
C123 VTAIL.n79 VSUBS 0.154166f
C124 VTAIL.n80 VSUBS 0.713799f
C125 VTAIL.n81 VSUBS 0.015361f
C126 VTAIL.n82 VSUBS 0.016264f
C127 VTAIL.n83 VSUBS 0.036307f
C128 VTAIL.n84 VSUBS 0.036307f
C129 VTAIL.n85 VSUBS 0.016264f
C130 VTAIL.n86 VSUBS 0.015361f
C131 VTAIL.n87 VSUBS 0.028586f
C132 VTAIL.n88 VSUBS 0.028586f
C133 VTAIL.n89 VSUBS 0.015361f
C134 VTAIL.n90 VSUBS 0.016264f
C135 VTAIL.n91 VSUBS 0.036307f
C136 VTAIL.n92 VSUBS 0.036307f
C137 VTAIL.n93 VSUBS 0.016264f
C138 VTAIL.n94 VSUBS 0.015361f
C139 VTAIL.n95 VSUBS 0.028586f
C140 VTAIL.n96 VSUBS 0.071151f
C141 VTAIL.n97 VSUBS 0.015361f
C142 VTAIL.n98 VSUBS 0.016264f
C143 VTAIL.n99 VSUBS 0.079646f
C144 VTAIL.n100 VSUBS 0.052293f
C145 VTAIL.n101 VSUBS 1.5943f
C146 VTAIL.n102 VSUBS 0.016071f
C147 VTAIL.n103 VSUBS 0.036307f
C148 VTAIL.n104 VSUBS 0.016264f
C149 VTAIL.n105 VSUBS 0.028586f
C150 VTAIL.n106 VSUBS 0.015361f
C151 VTAIL.n107 VSUBS 0.036307f
C152 VTAIL.n108 VSUBS 0.016264f
C153 VTAIL.n109 VSUBS 0.028586f
C154 VTAIL.n110 VSUBS 0.015361f
C155 VTAIL.n111 VSUBS 0.02723f
C156 VTAIL.n112 VSUBS 0.027308f
C157 VTAIL.t0 VSUBS 0.078023f
C158 VTAIL.n113 VSUBS 0.154166f
C159 VTAIL.n114 VSUBS 0.713799f
C160 VTAIL.n115 VSUBS 0.015361f
C161 VTAIL.n116 VSUBS 0.016264f
C162 VTAIL.n117 VSUBS 0.036307f
C163 VTAIL.n118 VSUBS 0.036307f
C164 VTAIL.n119 VSUBS 0.016264f
C165 VTAIL.n120 VSUBS 0.015361f
C166 VTAIL.n121 VSUBS 0.028586f
C167 VTAIL.n122 VSUBS 0.028586f
C168 VTAIL.n123 VSUBS 0.015361f
C169 VTAIL.n124 VSUBS 0.016264f
C170 VTAIL.n125 VSUBS 0.036307f
C171 VTAIL.n126 VSUBS 0.036307f
C172 VTAIL.n127 VSUBS 0.016264f
C173 VTAIL.n128 VSUBS 0.015361f
C174 VTAIL.n129 VSUBS 0.028586f
C175 VTAIL.n130 VSUBS 0.071151f
C176 VTAIL.n131 VSUBS 0.015361f
C177 VTAIL.n132 VSUBS 0.016264f
C178 VTAIL.n133 VSUBS 0.079646f
C179 VTAIL.n134 VSUBS 0.052293f
C180 VTAIL.n135 VSUBS 1.5943f
C181 VTAIL.n136 VSUBS 0.016071f
C182 VTAIL.n137 VSUBS 0.036307f
C183 VTAIL.n138 VSUBS 0.016264f
C184 VTAIL.n139 VSUBS 0.028586f
C185 VTAIL.n140 VSUBS 0.015361f
C186 VTAIL.n141 VSUBS 0.036307f
C187 VTAIL.n142 VSUBS 0.016264f
C188 VTAIL.n143 VSUBS 0.028586f
C189 VTAIL.n144 VSUBS 0.015361f
C190 VTAIL.n145 VSUBS 0.02723f
C191 VTAIL.n146 VSUBS 0.027308f
C192 VTAIL.t2 VSUBS 0.078023f
C193 VTAIL.n147 VSUBS 0.154166f
C194 VTAIL.n148 VSUBS 0.713799f
C195 VTAIL.n149 VSUBS 0.015361f
C196 VTAIL.n150 VSUBS 0.016264f
C197 VTAIL.n151 VSUBS 0.036307f
C198 VTAIL.n152 VSUBS 0.036307f
C199 VTAIL.n153 VSUBS 0.016264f
C200 VTAIL.n154 VSUBS 0.015361f
C201 VTAIL.n155 VSUBS 0.028586f
C202 VTAIL.n156 VSUBS 0.028586f
C203 VTAIL.n157 VSUBS 0.015361f
C204 VTAIL.n158 VSUBS 0.016264f
C205 VTAIL.n159 VSUBS 0.036307f
C206 VTAIL.n160 VSUBS 0.036307f
C207 VTAIL.n161 VSUBS 0.016264f
C208 VTAIL.n162 VSUBS 0.015361f
C209 VTAIL.n163 VSUBS 0.028586f
C210 VTAIL.n164 VSUBS 0.071151f
C211 VTAIL.n165 VSUBS 0.015361f
C212 VTAIL.n166 VSUBS 0.016264f
C213 VTAIL.n167 VSUBS 0.079646f
C214 VTAIL.n168 VSUBS 0.052293f
C215 VTAIL.n169 VSUBS 0.402029f
C216 VTAIL.n170 VSUBS 0.016071f
C217 VTAIL.n171 VSUBS 0.036307f
C218 VTAIL.n172 VSUBS 0.016264f
C219 VTAIL.n173 VSUBS 0.028586f
C220 VTAIL.n174 VSUBS 0.015361f
C221 VTAIL.n175 VSUBS 0.036307f
C222 VTAIL.n176 VSUBS 0.016264f
C223 VTAIL.n177 VSUBS 0.028586f
C224 VTAIL.n178 VSUBS 0.015361f
C225 VTAIL.n179 VSUBS 0.02723f
C226 VTAIL.n180 VSUBS 0.027308f
C227 VTAIL.t4 VSUBS 0.078023f
C228 VTAIL.n181 VSUBS 0.154166f
C229 VTAIL.n182 VSUBS 0.713799f
C230 VTAIL.n183 VSUBS 0.015361f
C231 VTAIL.n184 VSUBS 0.016264f
C232 VTAIL.n185 VSUBS 0.036307f
C233 VTAIL.n186 VSUBS 0.036307f
C234 VTAIL.n187 VSUBS 0.016264f
C235 VTAIL.n188 VSUBS 0.015361f
C236 VTAIL.n189 VSUBS 0.028586f
C237 VTAIL.n190 VSUBS 0.028586f
C238 VTAIL.n191 VSUBS 0.015361f
C239 VTAIL.n192 VSUBS 0.016264f
C240 VTAIL.n193 VSUBS 0.036307f
C241 VTAIL.n194 VSUBS 0.036307f
C242 VTAIL.n195 VSUBS 0.016264f
C243 VTAIL.n196 VSUBS 0.015361f
C244 VTAIL.n197 VSUBS 0.028586f
C245 VTAIL.n198 VSUBS 0.071151f
C246 VTAIL.n199 VSUBS 0.015361f
C247 VTAIL.n200 VSUBS 0.016264f
C248 VTAIL.n201 VSUBS 0.079646f
C249 VTAIL.n202 VSUBS 0.052293f
C250 VTAIL.n203 VSUBS 0.402029f
C251 VTAIL.n204 VSUBS 0.016071f
C252 VTAIL.n205 VSUBS 0.036307f
C253 VTAIL.n206 VSUBS 0.016264f
C254 VTAIL.n207 VSUBS 0.028586f
C255 VTAIL.n208 VSUBS 0.015361f
C256 VTAIL.n209 VSUBS 0.036307f
C257 VTAIL.n210 VSUBS 0.016264f
C258 VTAIL.n211 VSUBS 0.028586f
C259 VTAIL.n212 VSUBS 0.015361f
C260 VTAIL.n213 VSUBS 0.02723f
C261 VTAIL.n214 VSUBS 0.027308f
C262 VTAIL.t5 VSUBS 0.078023f
C263 VTAIL.n215 VSUBS 0.154166f
C264 VTAIL.n216 VSUBS 0.713799f
C265 VTAIL.n217 VSUBS 0.015361f
C266 VTAIL.n218 VSUBS 0.016264f
C267 VTAIL.n219 VSUBS 0.036307f
C268 VTAIL.n220 VSUBS 0.036307f
C269 VTAIL.n221 VSUBS 0.016264f
C270 VTAIL.n222 VSUBS 0.015361f
C271 VTAIL.n223 VSUBS 0.028586f
C272 VTAIL.n224 VSUBS 0.028586f
C273 VTAIL.n225 VSUBS 0.015361f
C274 VTAIL.n226 VSUBS 0.016264f
C275 VTAIL.n227 VSUBS 0.036307f
C276 VTAIL.n228 VSUBS 0.036307f
C277 VTAIL.n229 VSUBS 0.016264f
C278 VTAIL.n230 VSUBS 0.015361f
C279 VTAIL.n231 VSUBS 0.028586f
C280 VTAIL.n232 VSUBS 0.071151f
C281 VTAIL.n233 VSUBS 0.015361f
C282 VTAIL.n234 VSUBS 0.016264f
C283 VTAIL.n235 VSUBS 0.079646f
C284 VTAIL.n236 VSUBS 0.052293f
C285 VTAIL.n237 VSUBS 1.5943f
C286 VTAIL.n238 VSUBS 0.016071f
C287 VTAIL.n239 VSUBS 0.036307f
C288 VTAIL.n240 VSUBS 0.016264f
C289 VTAIL.n241 VSUBS 0.028586f
C290 VTAIL.n242 VSUBS 0.015361f
C291 VTAIL.n243 VSUBS 0.036307f
C292 VTAIL.n244 VSUBS 0.016264f
C293 VTAIL.n245 VSUBS 0.028586f
C294 VTAIL.n246 VSUBS 0.015361f
C295 VTAIL.n247 VSUBS 0.02723f
C296 VTAIL.n248 VSUBS 0.027308f
C297 VTAIL.t1 VSUBS 0.078023f
C298 VTAIL.n249 VSUBS 0.154166f
C299 VTAIL.n250 VSUBS 0.713799f
C300 VTAIL.n251 VSUBS 0.015361f
C301 VTAIL.n252 VSUBS 0.016264f
C302 VTAIL.n253 VSUBS 0.036307f
C303 VTAIL.n254 VSUBS 0.036307f
C304 VTAIL.n255 VSUBS 0.016264f
C305 VTAIL.n256 VSUBS 0.015361f
C306 VTAIL.n257 VSUBS 0.028586f
C307 VTAIL.n258 VSUBS 0.028586f
C308 VTAIL.n259 VSUBS 0.015361f
C309 VTAIL.n260 VSUBS 0.016264f
C310 VTAIL.n261 VSUBS 0.036307f
C311 VTAIL.n262 VSUBS 0.036307f
C312 VTAIL.n263 VSUBS 0.016264f
C313 VTAIL.n264 VSUBS 0.015361f
C314 VTAIL.n265 VSUBS 0.028586f
C315 VTAIL.n266 VSUBS 0.071151f
C316 VTAIL.n267 VSUBS 0.015361f
C317 VTAIL.n268 VSUBS 0.016264f
C318 VTAIL.n269 VSUBS 0.079646f
C319 VTAIL.n270 VSUBS 0.052293f
C320 VTAIL.n271 VSUBS 1.42299f
C321 VDD1.t1 VSUBS 0.147796f
C322 VDD1.t0 VSUBS 0.147796f
C323 VDD1.n0 VSUBS 1.02053f
C324 VDD1.t2 VSUBS 0.147796f
C325 VDD1.t3 VSUBS 0.147796f
C326 VDD1.n1 VSUBS 1.56919f
C327 VP.t1 VSUBS 2.5982f
C328 VP.n0 VSUBS 1.10083f
C329 VP.n1 VSUBS 0.039113f
C330 VP.n2 VSUBS 0.077738f
C331 VP.n3 VSUBS 0.039113f
C332 VP.n4 VSUBS 0.072898f
C333 VP.t3 VSUBS 3.18157f
C334 VP.t2 VSUBS 3.15929f
C335 VP.n5 VSUBS 4.1638f
C336 VP.n6 VSUBS 2.12719f
C337 VP.t0 VSUBS 2.5982f
C338 VP.n7 VSUBS 1.10083f
C339 VP.n8 VSUBS 0.043386f
C340 VP.n9 VSUBS 0.063128f
C341 VP.n10 VSUBS 0.039113f
C342 VP.n11 VSUBS 0.039113f
C343 VP.n12 VSUBS 0.072898f
C344 VP.n13 VSUBS 0.077738f
C345 VP.n14 VSUBS 0.031619f
C346 VP.n15 VSUBS 0.039113f
C347 VP.n16 VSUBS 0.039113f
C348 VP.n17 VSUBS 0.039113f
C349 VP.n18 VSUBS 0.072898f
C350 VP.n19 VSUBS 0.072898f
C351 VP.n20 VSUBS 0.043386f
C352 VP.n21 VSUBS 0.063128f
C353 VP.n22 VSUBS 0.119402f
C354 B.n0 VSUBS 0.005542f
C355 B.n1 VSUBS 0.005542f
C356 B.n2 VSUBS 0.008764f
C357 B.n3 VSUBS 0.008764f
C358 B.n4 VSUBS 0.008764f
C359 B.n5 VSUBS 0.008764f
C360 B.n6 VSUBS 0.008764f
C361 B.n7 VSUBS 0.008764f
C362 B.n8 VSUBS 0.008764f
C363 B.n9 VSUBS 0.008764f
C364 B.n10 VSUBS 0.008764f
C365 B.n11 VSUBS 0.008764f
C366 B.n12 VSUBS 0.008764f
C367 B.n13 VSUBS 0.008764f
C368 B.n14 VSUBS 0.008764f
C369 B.n15 VSUBS 0.008764f
C370 B.n16 VSUBS 0.008764f
C371 B.n17 VSUBS 0.008764f
C372 B.n18 VSUBS 0.008764f
C373 B.n19 VSUBS 0.008764f
C374 B.n20 VSUBS 0.008764f
C375 B.n21 VSUBS 0.008764f
C376 B.n22 VSUBS 0.008764f
C377 B.n23 VSUBS 0.008764f
C378 B.n24 VSUBS 0.020967f
C379 B.n25 VSUBS 0.008764f
C380 B.n26 VSUBS 0.008764f
C381 B.n27 VSUBS 0.008764f
C382 B.n28 VSUBS 0.008764f
C383 B.n29 VSUBS 0.008764f
C384 B.n30 VSUBS 0.008764f
C385 B.n31 VSUBS 0.008764f
C386 B.n32 VSUBS 0.008764f
C387 B.n33 VSUBS 0.008764f
C388 B.n34 VSUBS 0.008764f
C389 B.n35 VSUBS 0.008764f
C390 B.n36 VSUBS 0.008764f
C391 B.n37 VSUBS 0.008764f
C392 B.t2 VSUBS 0.122477f
C393 B.t1 VSUBS 0.168182f
C394 B.t0 VSUBS 1.50043f
C395 B.n38 VSUBS 0.27658f
C396 B.n39 VSUBS 0.214094f
C397 B.n40 VSUBS 0.008764f
C398 B.n41 VSUBS 0.008764f
C399 B.n42 VSUBS 0.008764f
C400 B.n43 VSUBS 0.008764f
C401 B.t11 VSUBS 0.12248f
C402 B.t10 VSUBS 0.168184f
C403 B.t9 VSUBS 1.50043f
C404 B.n44 VSUBS 0.276578f
C405 B.n45 VSUBS 0.214091f
C406 B.n46 VSUBS 0.020306f
C407 B.n47 VSUBS 0.008764f
C408 B.n48 VSUBS 0.008764f
C409 B.n49 VSUBS 0.008764f
C410 B.n50 VSUBS 0.008764f
C411 B.n51 VSUBS 0.008764f
C412 B.n52 VSUBS 0.008764f
C413 B.n53 VSUBS 0.008764f
C414 B.n54 VSUBS 0.008764f
C415 B.n55 VSUBS 0.008764f
C416 B.n56 VSUBS 0.008764f
C417 B.n57 VSUBS 0.008764f
C418 B.n58 VSUBS 0.008764f
C419 B.n59 VSUBS 0.020967f
C420 B.n60 VSUBS 0.008764f
C421 B.n61 VSUBS 0.008764f
C422 B.n62 VSUBS 0.008764f
C423 B.n63 VSUBS 0.008764f
C424 B.n64 VSUBS 0.008764f
C425 B.n65 VSUBS 0.008764f
C426 B.n66 VSUBS 0.008764f
C427 B.n67 VSUBS 0.008764f
C428 B.n68 VSUBS 0.008764f
C429 B.n69 VSUBS 0.008764f
C430 B.n70 VSUBS 0.008764f
C431 B.n71 VSUBS 0.008764f
C432 B.n72 VSUBS 0.008764f
C433 B.n73 VSUBS 0.008764f
C434 B.n74 VSUBS 0.008764f
C435 B.n75 VSUBS 0.008764f
C436 B.n76 VSUBS 0.008764f
C437 B.n77 VSUBS 0.008764f
C438 B.n78 VSUBS 0.008764f
C439 B.n79 VSUBS 0.008764f
C440 B.n80 VSUBS 0.008764f
C441 B.n81 VSUBS 0.008764f
C442 B.n82 VSUBS 0.008764f
C443 B.n83 VSUBS 0.008764f
C444 B.n84 VSUBS 0.008764f
C445 B.n85 VSUBS 0.008764f
C446 B.n86 VSUBS 0.008764f
C447 B.n87 VSUBS 0.008764f
C448 B.n88 VSUBS 0.008764f
C449 B.n89 VSUBS 0.008764f
C450 B.n90 VSUBS 0.008764f
C451 B.n91 VSUBS 0.008764f
C452 B.n92 VSUBS 0.008764f
C453 B.n93 VSUBS 0.008764f
C454 B.n94 VSUBS 0.008764f
C455 B.n95 VSUBS 0.008764f
C456 B.n96 VSUBS 0.008764f
C457 B.n97 VSUBS 0.008764f
C458 B.n98 VSUBS 0.008764f
C459 B.n99 VSUBS 0.008764f
C460 B.n100 VSUBS 0.008764f
C461 B.n101 VSUBS 0.008764f
C462 B.n102 VSUBS 0.008764f
C463 B.n103 VSUBS 0.008764f
C464 B.n104 VSUBS 0.020967f
C465 B.n105 VSUBS 0.008764f
C466 B.n106 VSUBS 0.008764f
C467 B.n107 VSUBS 0.008764f
C468 B.n108 VSUBS 0.008764f
C469 B.n109 VSUBS 0.008764f
C470 B.n110 VSUBS 0.008764f
C471 B.n111 VSUBS 0.008764f
C472 B.n112 VSUBS 0.008764f
C473 B.n113 VSUBS 0.008764f
C474 B.n114 VSUBS 0.008764f
C475 B.n115 VSUBS 0.008764f
C476 B.n116 VSUBS 0.008764f
C477 B.n117 VSUBS 0.008764f
C478 B.t7 VSUBS 0.12248f
C479 B.t8 VSUBS 0.168184f
C480 B.t6 VSUBS 1.50043f
C481 B.n118 VSUBS 0.276578f
C482 B.n119 VSUBS 0.214091f
C483 B.n120 VSUBS 0.008764f
C484 B.n121 VSUBS 0.008764f
C485 B.n122 VSUBS 0.008764f
C486 B.n123 VSUBS 0.008764f
C487 B.t4 VSUBS 0.122477f
C488 B.t5 VSUBS 0.168182f
C489 B.t3 VSUBS 1.50043f
C490 B.n124 VSUBS 0.27658f
C491 B.n125 VSUBS 0.214094f
C492 B.n126 VSUBS 0.020306f
C493 B.n127 VSUBS 0.008764f
C494 B.n128 VSUBS 0.008764f
C495 B.n129 VSUBS 0.008764f
C496 B.n130 VSUBS 0.008764f
C497 B.n131 VSUBS 0.008764f
C498 B.n132 VSUBS 0.008764f
C499 B.n133 VSUBS 0.008764f
C500 B.n134 VSUBS 0.008764f
C501 B.n135 VSUBS 0.008764f
C502 B.n136 VSUBS 0.008764f
C503 B.n137 VSUBS 0.008764f
C504 B.n138 VSUBS 0.008764f
C505 B.n139 VSUBS 0.020967f
C506 B.n140 VSUBS 0.008764f
C507 B.n141 VSUBS 0.008764f
C508 B.n142 VSUBS 0.008764f
C509 B.n143 VSUBS 0.008764f
C510 B.n144 VSUBS 0.008764f
C511 B.n145 VSUBS 0.008764f
C512 B.n146 VSUBS 0.008764f
C513 B.n147 VSUBS 0.008764f
C514 B.n148 VSUBS 0.008764f
C515 B.n149 VSUBS 0.008764f
C516 B.n150 VSUBS 0.008764f
C517 B.n151 VSUBS 0.008764f
C518 B.n152 VSUBS 0.008764f
C519 B.n153 VSUBS 0.008764f
C520 B.n154 VSUBS 0.008764f
C521 B.n155 VSUBS 0.008764f
C522 B.n156 VSUBS 0.008764f
C523 B.n157 VSUBS 0.008764f
C524 B.n158 VSUBS 0.008764f
C525 B.n159 VSUBS 0.008764f
C526 B.n160 VSUBS 0.008764f
C527 B.n161 VSUBS 0.008764f
C528 B.n162 VSUBS 0.008764f
C529 B.n163 VSUBS 0.008764f
C530 B.n164 VSUBS 0.008764f
C531 B.n165 VSUBS 0.008764f
C532 B.n166 VSUBS 0.008764f
C533 B.n167 VSUBS 0.008764f
C534 B.n168 VSUBS 0.008764f
C535 B.n169 VSUBS 0.008764f
C536 B.n170 VSUBS 0.008764f
C537 B.n171 VSUBS 0.008764f
C538 B.n172 VSUBS 0.008764f
C539 B.n173 VSUBS 0.008764f
C540 B.n174 VSUBS 0.008764f
C541 B.n175 VSUBS 0.008764f
C542 B.n176 VSUBS 0.008764f
C543 B.n177 VSUBS 0.008764f
C544 B.n178 VSUBS 0.008764f
C545 B.n179 VSUBS 0.008764f
C546 B.n180 VSUBS 0.008764f
C547 B.n181 VSUBS 0.008764f
C548 B.n182 VSUBS 0.008764f
C549 B.n183 VSUBS 0.008764f
C550 B.n184 VSUBS 0.008764f
C551 B.n185 VSUBS 0.008764f
C552 B.n186 VSUBS 0.008764f
C553 B.n187 VSUBS 0.008764f
C554 B.n188 VSUBS 0.008764f
C555 B.n189 VSUBS 0.008764f
C556 B.n190 VSUBS 0.008764f
C557 B.n191 VSUBS 0.008764f
C558 B.n192 VSUBS 0.008764f
C559 B.n193 VSUBS 0.008764f
C560 B.n194 VSUBS 0.008764f
C561 B.n195 VSUBS 0.008764f
C562 B.n196 VSUBS 0.008764f
C563 B.n197 VSUBS 0.008764f
C564 B.n198 VSUBS 0.008764f
C565 B.n199 VSUBS 0.008764f
C566 B.n200 VSUBS 0.008764f
C567 B.n201 VSUBS 0.008764f
C568 B.n202 VSUBS 0.008764f
C569 B.n203 VSUBS 0.008764f
C570 B.n204 VSUBS 0.008764f
C571 B.n205 VSUBS 0.008764f
C572 B.n206 VSUBS 0.008764f
C573 B.n207 VSUBS 0.008764f
C574 B.n208 VSUBS 0.008764f
C575 B.n209 VSUBS 0.008764f
C576 B.n210 VSUBS 0.008764f
C577 B.n211 VSUBS 0.008764f
C578 B.n212 VSUBS 0.008764f
C579 B.n213 VSUBS 0.008764f
C580 B.n214 VSUBS 0.008764f
C581 B.n215 VSUBS 0.008764f
C582 B.n216 VSUBS 0.008764f
C583 B.n217 VSUBS 0.008764f
C584 B.n218 VSUBS 0.008764f
C585 B.n219 VSUBS 0.008764f
C586 B.n220 VSUBS 0.008764f
C587 B.n221 VSUBS 0.008764f
C588 B.n222 VSUBS 0.008764f
C589 B.n223 VSUBS 0.008764f
C590 B.n224 VSUBS 0.008764f
C591 B.n225 VSUBS 0.008764f
C592 B.n226 VSUBS 0.020967f
C593 B.n227 VSUBS 0.021565f
C594 B.n228 VSUBS 0.021565f
C595 B.n229 VSUBS 0.008764f
C596 B.n230 VSUBS 0.008764f
C597 B.n231 VSUBS 0.008764f
C598 B.n232 VSUBS 0.008764f
C599 B.n233 VSUBS 0.008764f
C600 B.n234 VSUBS 0.008764f
C601 B.n235 VSUBS 0.008764f
C602 B.n236 VSUBS 0.008764f
C603 B.n237 VSUBS 0.008764f
C604 B.n238 VSUBS 0.008764f
C605 B.n239 VSUBS 0.008764f
C606 B.n240 VSUBS 0.008764f
C607 B.n241 VSUBS 0.008764f
C608 B.n242 VSUBS 0.008764f
C609 B.n243 VSUBS 0.008764f
C610 B.n244 VSUBS 0.008764f
C611 B.n245 VSUBS 0.008764f
C612 B.n246 VSUBS 0.008764f
C613 B.n247 VSUBS 0.008764f
C614 B.n248 VSUBS 0.008764f
C615 B.n249 VSUBS 0.008764f
C616 B.n250 VSUBS 0.008764f
C617 B.n251 VSUBS 0.008764f
C618 B.n252 VSUBS 0.008764f
C619 B.n253 VSUBS 0.008764f
C620 B.n254 VSUBS 0.008764f
C621 B.n255 VSUBS 0.008764f
C622 B.n256 VSUBS 0.008764f
C623 B.n257 VSUBS 0.008764f
C624 B.n258 VSUBS 0.008764f
C625 B.n259 VSUBS 0.008764f
C626 B.n260 VSUBS 0.008764f
C627 B.n261 VSUBS 0.008764f
C628 B.n262 VSUBS 0.008764f
C629 B.n263 VSUBS 0.008249f
C630 B.n264 VSUBS 0.008764f
C631 B.n265 VSUBS 0.008764f
C632 B.n266 VSUBS 0.004898f
C633 B.n267 VSUBS 0.008764f
C634 B.n268 VSUBS 0.008764f
C635 B.n269 VSUBS 0.008764f
C636 B.n270 VSUBS 0.008764f
C637 B.n271 VSUBS 0.008764f
C638 B.n272 VSUBS 0.008764f
C639 B.n273 VSUBS 0.008764f
C640 B.n274 VSUBS 0.008764f
C641 B.n275 VSUBS 0.008764f
C642 B.n276 VSUBS 0.008764f
C643 B.n277 VSUBS 0.008764f
C644 B.n278 VSUBS 0.008764f
C645 B.n279 VSUBS 0.004898f
C646 B.n280 VSUBS 0.020306f
C647 B.n281 VSUBS 0.008249f
C648 B.n282 VSUBS 0.008764f
C649 B.n283 VSUBS 0.008764f
C650 B.n284 VSUBS 0.008764f
C651 B.n285 VSUBS 0.008764f
C652 B.n286 VSUBS 0.008764f
C653 B.n287 VSUBS 0.008764f
C654 B.n288 VSUBS 0.008764f
C655 B.n289 VSUBS 0.008764f
C656 B.n290 VSUBS 0.008764f
C657 B.n291 VSUBS 0.008764f
C658 B.n292 VSUBS 0.008764f
C659 B.n293 VSUBS 0.008764f
C660 B.n294 VSUBS 0.008764f
C661 B.n295 VSUBS 0.008764f
C662 B.n296 VSUBS 0.008764f
C663 B.n297 VSUBS 0.008764f
C664 B.n298 VSUBS 0.008764f
C665 B.n299 VSUBS 0.008764f
C666 B.n300 VSUBS 0.008764f
C667 B.n301 VSUBS 0.008764f
C668 B.n302 VSUBS 0.008764f
C669 B.n303 VSUBS 0.008764f
C670 B.n304 VSUBS 0.008764f
C671 B.n305 VSUBS 0.008764f
C672 B.n306 VSUBS 0.008764f
C673 B.n307 VSUBS 0.008764f
C674 B.n308 VSUBS 0.008764f
C675 B.n309 VSUBS 0.008764f
C676 B.n310 VSUBS 0.008764f
C677 B.n311 VSUBS 0.008764f
C678 B.n312 VSUBS 0.008764f
C679 B.n313 VSUBS 0.008764f
C680 B.n314 VSUBS 0.008764f
C681 B.n315 VSUBS 0.008764f
C682 B.n316 VSUBS 0.008764f
C683 B.n317 VSUBS 0.021565f
C684 B.n318 VSUBS 0.021565f
C685 B.n319 VSUBS 0.020967f
C686 B.n320 VSUBS 0.008764f
C687 B.n321 VSUBS 0.008764f
C688 B.n322 VSUBS 0.008764f
C689 B.n323 VSUBS 0.008764f
C690 B.n324 VSUBS 0.008764f
C691 B.n325 VSUBS 0.008764f
C692 B.n326 VSUBS 0.008764f
C693 B.n327 VSUBS 0.008764f
C694 B.n328 VSUBS 0.008764f
C695 B.n329 VSUBS 0.008764f
C696 B.n330 VSUBS 0.008764f
C697 B.n331 VSUBS 0.008764f
C698 B.n332 VSUBS 0.008764f
C699 B.n333 VSUBS 0.008764f
C700 B.n334 VSUBS 0.008764f
C701 B.n335 VSUBS 0.008764f
C702 B.n336 VSUBS 0.008764f
C703 B.n337 VSUBS 0.008764f
C704 B.n338 VSUBS 0.008764f
C705 B.n339 VSUBS 0.008764f
C706 B.n340 VSUBS 0.008764f
C707 B.n341 VSUBS 0.008764f
C708 B.n342 VSUBS 0.008764f
C709 B.n343 VSUBS 0.008764f
C710 B.n344 VSUBS 0.008764f
C711 B.n345 VSUBS 0.008764f
C712 B.n346 VSUBS 0.008764f
C713 B.n347 VSUBS 0.008764f
C714 B.n348 VSUBS 0.008764f
C715 B.n349 VSUBS 0.008764f
C716 B.n350 VSUBS 0.008764f
C717 B.n351 VSUBS 0.008764f
C718 B.n352 VSUBS 0.008764f
C719 B.n353 VSUBS 0.008764f
C720 B.n354 VSUBS 0.008764f
C721 B.n355 VSUBS 0.008764f
C722 B.n356 VSUBS 0.008764f
C723 B.n357 VSUBS 0.008764f
C724 B.n358 VSUBS 0.008764f
C725 B.n359 VSUBS 0.008764f
C726 B.n360 VSUBS 0.008764f
C727 B.n361 VSUBS 0.008764f
C728 B.n362 VSUBS 0.008764f
C729 B.n363 VSUBS 0.008764f
C730 B.n364 VSUBS 0.008764f
C731 B.n365 VSUBS 0.008764f
C732 B.n366 VSUBS 0.008764f
C733 B.n367 VSUBS 0.008764f
C734 B.n368 VSUBS 0.008764f
C735 B.n369 VSUBS 0.008764f
C736 B.n370 VSUBS 0.008764f
C737 B.n371 VSUBS 0.008764f
C738 B.n372 VSUBS 0.008764f
C739 B.n373 VSUBS 0.008764f
C740 B.n374 VSUBS 0.008764f
C741 B.n375 VSUBS 0.008764f
C742 B.n376 VSUBS 0.008764f
C743 B.n377 VSUBS 0.008764f
C744 B.n378 VSUBS 0.008764f
C745 B.n379 VSUBS 0.008764f
C746 B.n380 VSUBS 0.008764f
C747 B.n381 VSUBS 0.008764f
C748 B.n382 VSUBS 0.008764f
C749 B.n383 VSUBS 0.008764f
C750 B.n384 VSUBS 0.008764f
C751 B.n385 VSUBS 0.008764f
C752 B.n386 VSUBS 0.008764f
C753 B.n387 VSUBS 0.008764f
C754 B.n388 VSUBS 0.008764f
C755 B.n389 VSUBS 0.008764f
C756 B.n390 VSUBS 0.008764f
C757 B.n391 VSUBS 0.008764f
C758 B.n392 VSUBS 0.008764f
C759 B.n393 VSUBS 0.008764f
C760 B.n394 VSUBS 0.008764f
C761 B.n395 VSUBS 0.008764f
C762 B.n396 VSUBS 0.008764f
C763 B.n397 VSUBS 0.008764f
C764 B.n398 VSUBS 0.008764f
C765 B.n399 VSUBS 0.008764f
C766 B.n400 VSUBS 0.008764f
C767 B.n401 VSUBS 0.008764f
C768 B.n402 VSUBS 0.008764f
C769 B.n403 VSUBS 0.008764f
C770 B.n404 VSUBS 0.008764f
C771 B.n405 VSUBS 0.008764f
C772 B.n406 VSUBS 0.008764f
C773 B.n407 VSUBS 0.008764f
C774 B.n408 VSUBS 0.008764f
C775 B.n409 VSUBS 0.008764f
C776 B.n410 VSUBS 0.008764f
C777 B.n411 VSUBS 0.008764f
C778 B.n412 VSUBS 0.008764f
C779 B.n413 VSUBS 0.008764f
C780 B.n414 VSUBS 0.008764f
C781 B.n415 VSUBS 0.008764f
C782 B.n416 VSUBS 0.008764f
C783 B.n417 VSUBS 0.008764f
C784 B.n418 VSUBS 0.008764f
C785 B.n419 VSUBS 0.008764f
C786 B.n420 VSUBS 0.008764f
C787 B.n421 VSUBS 0.008764f
C788 B.n422 VSUBS 0.008764f
C789 B.n423 VSUBS 0.008764f
C790 B.n424 VSUBS 0.008764f
C791 B.n425 VSUBS 0.008764f
C792 B.n426 VSUBS 0.008764f
C793 B.n427 VSUBS 0.008764f
C794 B.n428 VSUBS 0.008764f
C795 B.n429 VSUBS 0.008764f
C796 B.n430 VSUBS 0.008764f
C797 B.n431 VSUBS 0.008764f
C798 B.n432 VSUBS 0.008764f
C799 B.n433 VSUBS 0.008764f
C800 B.n434 VSUBS 0.008764f
C801 B.n435 VSUBS 0.008764f
C802 B.n436 VSUBS 0.008764f
C803 B.n437 VSUBS 0.008764f
C804 B.n438 VSUBS 0.008764f
C805 B.n439 VSUBS 0.008764f
C806 B.n440 VSUBS 0.008764f
C807 B.n441 VSUBS 0.008764f
C808 B.n442 VSUBS 0.008764f
C809 B.n443 VSUBS 0.008764f
C810 B.n444 VSUBS 0.008764f
C811 B.n445 VSUBS 0.008764f
C812 B.n446 VSUBS 0.008764f
C813 B.n447 VSUBS 0.008764f
C814 B.n448 VSUBS 0.008764f
C815 B.n449 VSUBS 0.008764f
C816 B.n450 VSUBS 0.008764f
C817 B.n451 VSUBS 0.008764f
C818 B.n452 VSUBS 0.008764f
C819 B.n453 VSUBS 0.008764f
C820 B.n454 VSUBS 0.021947f
C821 B.n455 VSUBS 0.020584f
C822 B.n456 VSUBS 0.021565f
C823 B.n457 VSUBS 0.008764f
C824 B.n458 VSUBS 0.008764f
C825 B.n459 VSUBS 0.008764f
C826 B.n460 VSUBS 0.008764f
C827 B.n461 VSUBS 0.008764f
C828 B.n462 VSUBS 0.008764f
C829 B.n463 VSUBS 0.008764f
C830 B.n464 VSUBS 0.008764f
C831 B.n465 VSUBS 0.008764f
C832 B.n466 VSUBS 0.008764f
C833 B.n467 VSUBS 0.008764f
C834 B.n468 VSUBS 0.008764f
C835 B.n469 VSUBS 0.008764f
C836 B.n470 VSUBS 0.008764f
C837 B.n471 VSUBS 0.008764f
C838 B.n472 VSUBS 0.008764f
C839 B.n473 VSUBS 0.008764f
C840 B.n474 VSUBS 0.008764f
C841 B.n475 VSUBS 0.008764f
C842 B.n476 VSUBS 0.008764f
C843 B.n477 VSUBS 0.008764f
C844 B.n478 VSUBS 0.008764f
C845 B.n479 VSUBS 0.008764f
C846 B.n480 VSUBS 0.008764f
C847 B.n481 VSUBS 0.008764f
C848 B.n482 VSUBS 0.008764f
C849 B.n483 VSUBS 0.008764f
C850 B.n484 VSUBS 0.008764f
C851 B.n485 VSUBS 0.008764f
C852 B.n486 VSUBS 0.008764f
C853 B.n487 VSUBS 0.008764f
C854 B.n488 VSUBS 0.008764f
C855 B.n489 VSUBS 0.008764f
C856 B.n490 VSUBS 0.008764f
C857 B.n491 VSUBS 0.008249f
C858 B.n492 VSUBS 0.008764f
C859 B.n493 VSUBS 0.008764f
C860 B.n494 VSUBS 0.004898f
C861 B.n495 VSUBS 0.008764f
C862 B.n496 VSUBS 0.008764f
C863 B.n497 VSUBS 0.008764f
C864 B.n498 VSUBS 0.008764f
C865 B.n499 VSUBS 0.008764f
C866 B.n500 VSUBS 0.008764f
C867 B.n501 VSUBS 0.008764f
C868 B.n502 VSUBS 0.008764f
C869 B.n503 VSUBS 0.008764f
C870 B.n504 VSUBS 0.008764f
C871 B.n505 VSUBS 0.008764f
C872 B.n506 VSUBS 0.008764f
C873 B.n507 VSUBS 0.004898f
C874 B.n508 VSUBS 0.020306f
C875 B.n509 VSUBS 0.008249f
C876 B.n510 VSUBS 0.008764f
C877 B.n511 VSUBS 0.008764f
C878 B.n512 VSUBS 0.008764f
C879 B.n513 VSUBS 0.008764f
C880 B.n514 VSUBS 0.008764f
C881 B.n515 VSUBS 0.008764f
C882 B.n516 VSUBS 0.008764f
C883 B.n517 VSUBS 0.008764f
C884 B.n518 VSUBS 0.008764f
C885 B.n519 VSUBS 0.008764f
C886 B.n520 VSUBS 0.008764f
C887 B.n521 VSUBS 0.008764f
C888 B.n522 VSUBS 0.008764f
C889 B.n523 VSUBS 0.008764f
C890 B.n524 VSUBS 0.008764f
C891 B.n525 VSUBS 0.008764f
C892 B.n526 VSUBS 0.008764f
C893 B.n527 VSUBS 0.008764f
C894 B.n528 VSUBS 0.008764f
C895 B.n529 VSUBS 0.008764f
C896 B.n530 VSUBS 0.008764f
C897 B.n531 VSUBS 0.008764f
C898 B.n532 VSUBS 0.008764f
C899 B.n533 VSUBS 0.008764f
C900 B.n534 VSUBS 0.008764f
C901 B.n535 VSUBS 0.008764f
C902 B.n536 VSUBS 0.008764f
C903 B.n537 VSUBS 0.008764f
C904 B.n538 VSUBS 0.008764f
C905 B.n539 VSUBS 0.008764f
C906 B.n540 VSUBS 0.008764f
C907 B.n541 VSUBS 0.008764f
C908 B.n542 VSUBS 0.008764f
C909 B.n543 VSUBS 0.008764f
C910 B.n544 VSUBS 0.008764f
C911 B.n545 VSUBS 0.021565f
C912 B.n546 VSUBS 0.021565f
C913 B.n547 VSUBS 0.020967f
C914 B.n548 VSUBS 0.008764f
C915 B.n549 VSUBS 0.008764f
C916 B.n550 VSUBS 0.008764f
C917 B.n551 VSUBS 0.008764f
C918 B.n552 VSUBS 0.008764f
C919 B.n553 VSUBS 0.008764f
C920 B.n554 VSUBS 0.008764f
C921 B.n555 VSUBS 0.008764f
C922 B.n556 VSUBS 0.008764f
C923 B.n557 VSUBS 0.008764f
C924 B.n558 VSUBS 0.008764f
C925 B.n559 VSUBS 0.008764f
C926 B.n560 VSUBS 0.008764f
C927 B.n561 VSUBS 0.008764f
C928 B.n562 VSUBS 0.008764f
C929 B.n563 VSUBS 0.008764f
C930 B.n564 VSUBS 0.008764f
C931 B.n565 VSUBS 0.008764f
C932 B.n566 VSUBS 0.008764f
C933 B.n567 VSUBS 0.008764f
C934 B.n568 VSUBS 0.008764f
C935 B.n569 VSUBS 0.008764f
C936 B.n570 VSUBS 0.008764f
C937 B.n571 VSUBS 0.008764f
C938 B.n572 VSUBS 0.008764f
C939 B.n573 VSUBS 0.008764f
C940 B.n574 VSUBS 0.008764f
C941 B.n575 VSUBS 0.008764f
C942 B.n576 VSUBS 0.008764f
C943 B.n577 VSUBS 0.008764f
C944 B.n578 VSUBS 0.008764f
C945 B.n579 VSUBS 0.008764f
C946 B.n580 VSUBS 0.008764f
C947 B.n581 VSUBS 0.008764f
C948 B.n582 VSUBS 0.008764f
C949 B.n583 VSUBS 0.008764f
C950 B.n584 VSUBS 0.008764f
C951 B.n585 VSUBS 0.008764f
C952 B.n586 VSUBS 0.008764f
C953 B.n587 VSUBS 0.008764f
C954 B.n588 VSUBS 0.008764f
C955 B.n589 VSUBS 0.008764f
C956 B.n590 VSUBS 0.008764f
C957 B.n591 VSUBS 0.008764f
C958 B.n592 VSUBS 0.008764f
C959 B.n593 VSUBS 0.008764f
C960 B.n594 VSUBS 0.008764f
C961 B.n595 VSUBS 0.008764f
C962 B.n596 VSUBS 0.008764f
C963 B.n597 VSUBS 0.008764f
C964 B.n598 VSUBS 0.008764f
C965 B.n599 VSUBS 0.008764f
C966 B.n600 VSUBS 0.008764f
C967 B.n601 VSUBS 0.008764f
C968 B.n602 VSUBS 0.008764f
C969 B.n603 VSUBS 0.008764f
C970 B.n604 VSUBS 0.008764f
C971 B.n605 VSUBS 0.008764f
C972 B.n606 VSUBS 0.008764f
C973 B.n607 VSUBS 0.008764f
C974 B.n608 VSUBS 0.008764f
C975 B.n609 VSUBS 0.008764f
C976 B.n610 VSUBS 0.008764f
C977 B.n611 VSUBS 0.008764f
C978 B.n612 VSUBS 0.008764f
C979 B.n613 VSUBS 0.008764f
C980 B.n614 VSUBS 0.008764f
C981 B.n615 VSUBS 0.019845f
.ends

