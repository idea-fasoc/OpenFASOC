* NGSPICE file created from diff_pair_sample_0909.ext - technology: sky130A

.subckt diff_pair_sample_0909 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=2.21
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=2.21
X2 VTAIL.t7 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=2.21
X3 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=2.21
X4 VDD1.t2 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=2.21
X5 VDD1.t0 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=2.21
X6 VDD2.t3 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=2.21
X7 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=2.21
X8 VTAIL.t3 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=2.21
X9 VTAIL.t4 VP.t3 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=2.21
X10 VDD2.t0 VN.t3 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=2.21
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=2.21
R0 B.n380 B.n83 585
R1 B.n83 B.n58 585
R2 B.n382 B.n381 585
R3 B.n384 B.n82 585
R4 B.n387 B.n386 585
R5 B.n388 B.n81 585
R6 B.n390 B.n389 585
R7 B.n392 B.n80 585
R8 B.n395 B.n394 585
R9 B.n396 B.n79 585
R10 B.n398 B.n397 585
R11 B.n400 B.n78 585
R12 B.n403 B.n402 585
R13 B.n404 B.n77 585
R14 B.n406 B.n405 585
R15 B.n408 B.n76 585
R16 B.n411 B.n410 585
R17 B.n413 B.n73 585
R18 B.n415 B.n414 585
R19 B.n417 B.n72 585
R20 B.n420 B.n419 585
R21 B.n421 B.n71 585
R22 B.n423 B.n422 585
R23 B.n425 B.n70 585
R24 B.n428 B.n427 585
R25 B.n429 B.n67 585
R26 B.n432 B.n431 585
R27 B.n434 B.n66 585
R28 B.n437 B.n436 585
R29 B.n438 B.n65 585
R30 B.n440 B.n439 585
R31 B.n442 B.n64 585
R32 B.n445 B.n444 585
R33 B.n446 B.n63 585
R34 B.n448 B.n447 585
R35 B.n450 B.n62 585
R36 B.n453 B.n452 585
R37 B.n454 B.n61 585
R38 B.n456 B.n455 585
R39 B.n458 B.n60 585
R40 B.n461 B.n460 585
R41 B.n462 B.n59 585
R42 B.n379 B.n57 585
R43 B.n465 B.n57 585
R44 B.n378 B.n56 585
R45 B.n466 B.n56 585
R46 B.n377 B.n55 585
R47 B.n467 B.n55 585
R48 B.n376 B.n375 585
R49 B.n375 B.n51 585
R50 B.n374 B.n50 585
R51 B.n473 B.n50 585
R52 B.n373 B.n49 585
R53 B.n474 B.n49 585
R54 B.n372 B.n48 585
R55 B.n475 B.n48 585
R56 B.n371 B.n370 585
R57 B.n370 B.n47 585
R58 B.n369 B.n43 585
R59 B.n481 B.n43 585
R60 B.n368 B.n42 585
R61 B.n482 B.n42 585
R62 B.n367 B.n41 585
R63 B.n483 B.n41 585
R64 B.n366 B.n365 585
R65 B.n365 B.n37 585
R66 B.n364 B.n36 585
R67 B.n489 B.n36 585
R68 B.n363 B.n35 585
R69 B.n490 B.n35 585
R70 B.n362 B.n34 585
R71 B.n491 B.n34 585
R72 B.n361 B.n360 585
R73 B.n360 B.n30 585
R74 B.n359 B.n29 585
R75 B.n497 B.n29 585
R76 B.n358 B.n28 585
R77 B.n498 B.n28 585
R78 B.n357 B.n27 585
R79 B.n499 B.n27 585
R80 B.n356 B.n355 585
R81 B.n355 B.n23 585
R82 B.n354 B.n22 585
R83 B.n505 B.n22 585
R84 B.n353 B.n21 585
R85 B.n506 B.n21 585
R86 B.n352 B.n20 585
R87 B.n507 B.n20 585
R88 B.n351 B.n350 585
R89 B.n350 B.n16 585
R90 B.n349 B.n15 585
R91 B.n513 B.n15 585
R92 B.n348 B.n14 585
R93 B.n514 B.n14 585
R94 B.n347 B.n13 585
R95 B.n515 B.n13 585
R96 B.n346 B.n345 585
R97 B.n345 B.n12 585
R98 B.n344 B.n343 585
R99 B.n344 B.n8 585
R100 B.n342 B.n7 585
R101 B.n522 B.n7 585
R102 B.n341 B.n6 585
R103 B.n523 B.n6 585
R104 B.n340 B.n5 585
R105 B.n524 B.n5 585
R106 B.n339 B.n338 585
R107 B.n338 B.n4 585
R108 B.n337 B.n84 585
R109 B.n337 B.n336 585
R110 B.n327 B.n85 585
R111 B.n86 B.n85 585
R112 B.n329 B.n328 585
R113 B.n330 B.n329 585
R114 B.n326 B.n90 585
R115 B.n94 B.n90 585
R116 B.n325 B.n324 585
R117 B.n324 B.n323 585
R118 B.n92 B.n91 585
R119 B.n93 B.n92 585
R120 B.n316 B.n315 585
R121 B.n317 B.n316 585
R122 B.n314 B.n99 585
R123 B.n99 B.n98 585
R124 B.n313 B.n312 585
R125 B.n312 B.n311 585
R126 B.n101 B.n100 585
R127 B.n102 B.n101 585
R128 B.n304 B.n303 585
R129 B.n305 B.n304 585
R130 B.n302 B.n106 585
R131 B.n110 B.n106 585
R132 B.n301 B.n300 585
R133 B.n300 B.n299 585
R134 B.n108 B.n107 585
R135 B.n109 B.n108 585
R136 B.n292 B.n291 585
R137 B.n293 B.n292 585
R138 B.n290 B.n115 585
R139 B.n115 B.n114 585
R140 B.n289 B.n288 585
R141 B.n288 B.n287 585
R142 B.n117 B.n116 585
R143 B.n118 B.n117 585
R144 B.n280 B.n279 585
R145 B.n281 B.n280 585
R146 B.n278 B.n123 585
R147 B.n123 B.n122 585
R148 B.n277 B.n276 585
R149 B.n276 B.n275 585
R150 B.n125 B.n124 585
R151 B.n268 B.n125 585
R152 B.n267 B.n266 585
R153 B.n269 B.n267 585
R154 B.n265 B.n130 585
R155 B.n130 B.n129 585
R156 B.n264 B.n263 585
R157 B.n263 B.n262 585
R158 B.n132 B.n131 585
R159 B.n133 B.n132 585
R160 B.n255 B.n254 585
R161 B.n256 B.n255 585
R162 B.n253 B.n138 585
R163 B.n138 B.n137 585
R164 B.n252 B.n251 585
R165 B.n251 B.n250 585
R166 B.n247 B.n142 585
R167 B.n246 B.n245 585
R168 B.n243 B.n143 585
R169 B.n243 B.n141 585
R170 B.n242 B.n241 585
R171 B.n240 B.n239 585
R172 B.n238 B.n145 585
R173 B.n236 B.n235 585
R174 B.n234 B.n146 585
R175 B.n233 B.n232 585
R176 B.n230 B.n147 585
R177 B.n228 B.n227 585
R178 B.n226 B.n148 585
R179 B.n225 B.n224 585
R180 B.n222 B.n149 585
R181 B.n220 B.n219 585
R182 B.n218 B.n150 585
R183 B.n216 B.n215 585
R184 B.n213 B.n153 585
R185 B.n211 B.n210 585
R186 B.n209 B.n154 585
R187 B.n208 B.n207 585
R188 B.n205 B.n155 585
R189 B.n203 B.n202 585
R190 B.n201 B.n156 585
R191 B.n200 B.n199 585
R192 B.n197 B.n196 585
R193 B.n195 B.n194 585
R194 B.n193 B.n161 585
R195 B.n191 B.n190 585
R196 B.n189 B.n162 585
R197 B.n188 B.n187 585
R198 B.n185 B.n163 585
R199 B.n183 B.n182 585
R200 B.n181 B.n164 585
R201 B.n180 B.n179 585
R202 B.n177 B.n165 585
R203 B.n175 B.n174 585
R204 B.n173 B.n166 585
R205 B.n172 B.n171 585
R206 B.n169 B.n167 585
R207 B.n140 B.n139 585
R208 B.n249 B.n248 585
R209 B.n250 B.n249 585
R210 B.n136 B.n135 585
R211 B.n137 B.n136 585
R212 B.n258 B.n257 585
R213 B.n257 B.n256 585
R214 B.n259 B.n134 585
R215 B.n134 B.n133 585
R216 B.n261 B.n260 585
R217 B.n262 B.n261 585
R218 B.n128 B.n127 585
R219 B.n129 B.n128 585
R220 B.n271 B.n270 585
R221 B.n270 B.n269 585
R222 B.n272 B.n126 585
R223 B.n268 B.n126 585
R224 B.n274 B.n273 585
R225 B.n275 B.n274 585
R226 B.n121 B.n120 585
R227 B.n122 B.n121 585
R228 B.n283 B.n282 585
R229 B.n282 B.n281 585
R230 B.n284 B.n119 585
R231 B.n119 B.n118 585
R232 B.n286 B.n285 585
R233 B.n287 B.n286 585
R234 B.n113 B.n112 585
R235 B.n114 B.n113 585
R236 B.n295 B.n294 585
R237 B.n294 B.n293 585
R238 B.n296 B.n111 585
R239 B.n111 B.n109 585
R240 B.n298 B.n297 585
R241 B.n299 B.n298 585
R242 B.n105 B.n104 585
R243 B.n110 B.n105 585
R244 B.n307 B.n306 585
R245 B.n306 B.n305 585
R246 B.n308 B.n103 585
R247 B.n103 B.n102 585
R248 B.n310 B.n309 585
R249 B.n311 B.n310 585
R250 B.n97 B.n96 585
R251 B.n98 B.n97 585
R252 B.n319 B.n318 585
R253 B.n318 B.n317 585
R254 B.n320 B.n95 585
R255 B.n95 B.n93 585
R256 B.n322 B.n321 585
R257 B.n323 B.n322 585
R258 B.n89 B.n88 585
R259 B.n94 B.n89 585
R260 B.n332 B.n331 585
R261 B.n331 B.n330 585
R262 B.n333 B.n87 585
R263 B.n87 B.n86 585
R264 B.n335 B.n334 585
R265 B.n336 B.n335 585
R266 B.n3 B.n0 585
R267 B.n4 B.n3 585
R268 B.n521 B.n1 585
R269 B.n522 B.n521 585
R270 B.n520 B.n519 585
R271 B.n520 B.n8 585
R272 B.n518 B.n9 585
R273 B.n12 B.n9 585
R274 B.n517 B.n516 585
R275 B.n516 B.n515 585
R276 B.n11 B.n10 585
R277 B.n514 B.n11 585
R278 B.n512 B.n511 585
R279 B.n513 B.n512 585
R280 B.n510 B.n17 585
R281 B.n17 B.n16 585
R282 B.n509 B.n508 585
R283 B.n508 B.n507 585
R284 B.n19 B.n18 585
R285 B.n506 B.n19 585
R286 B.n504 B.n503 585
R287 B.n505 B.n504 585
R288 B.n502 B.n24 585
R289 B.n24 B.n23 585
R290 B.n501 B.n500 585
R291 B.n500 B.n499 585
R292 B.n26 B.n25 585
R293 B.n498 B.n26 585
R294 B.n496 B.n495 585
R295 B.n497 B.n496 585
R296 B.n494 B.n31 585
R297 B.n31 B.n30 585
R298 B.n493 B.n492 585
R299 B.n492 B.n491 585
R300 B.n33 B.n32 585
R301 B.n490 B.n33 585
R302 B.n488 B.n487 585
R303 B.n489 B.n488 585
R304 B.n486 B.n38 585
R305 B.n38 B.n37 585
R306 B.n485 B.n484 585
R307 B.n484 B.n483 585
R308 B.n40 B.n39 585
R309 B.n482 B.n40 585
R310 B.n480 B.n479 585
R311 B.n481 B.n480 585
R312 B.n478 B.n44 585
R313 B.n47 B.n44 585
R314 B.n477 B.n476 585
R315 B.n476 B.n475 585
R316 B.n46 B.n45 585
R317 B.n474 B.n46 585
R318 B.n472 B.n471 585
R319 B.n473 B.n472 585
R320 B.n470 B.n52 585
R321 B.n52 B.n51 585
R322 B.n469 B.n468 585
R323 B.n468 B.n467 585
R324 B.n54 B.n53 585
R325 B.n466 B.n54 585
R326 B.n464 B.n463 585
R327 B.n465 B.n464 585
R328 B.n525 B.n524 585
R329 B.n523 B.n2 585
R330 B.n464 B.n59 540.549
R331 B.n83 B.n57 540.549
R332 B.n251 B.n140 540.549
R333 B.n249 B.n142 540.549
R334 B.n383 B.n58 256.663
R335 B.n385 B.n58 256.663
R336 B.n391 B.n58 256.663
R337 B.n393 B.n58 256.663
R338 B.n399 B.n58 256.663
R339 B.n401 B.n58 256.663
R340 B.n407 B.n58 256.663
R341 B.n409 B.n58 256.663
R342 B.n416 B.n58 256.663
R343 B.n418 B.n58 256.663
R344 B.n424 B.n58 256.663
R345 B.n426 B.n58 256.663
R346 B.n433 B.n58 256.663
R347 B.n435 B.n58 256.663
R348 B.n441 B.n58 256.663
R349 B.n443 B.n58 256.663
R350 B.n449 B.n58 256.663
R351 B.n451 B.n58 256.663
R352 B.n457 B.n58 256.663
R353 B.n459 B.n58 256.663
R354 B.n244 B.n141 256.663
R355 B.n144 B.n141 256.663
R356 B.n237 B.n141 256.663
R357 B.n231 B.n141 256.663
R358 B.n229 B.n141 256.663
R359 B.n223 B.n141 256.663
R360 B.n221 B.n141 256.663
R361 B.n214 B.n141 256.663
R362 B.n212 B.n141 256.663
R363 B.n206 B.n141 256.663
R364 B.n204 B.n141 256.663
R365 B.n198 B.n141 256.663
R366 B.n160 B.n141 256.663
R367 B.n192 B.n141 256.663
R368 B.n186 B.n141 256.663
R369 B.n184 B.n141 256.663
R370 B.n178 B.n141 256.663
R371 B.n176 B.n141 256.663
R372 B.n170 B.n141 256.663
R373 B.n168 B.n141 256.663
R374 B.n527 B.n526 256.663
R375 B.n68 B.t8 243.03
R376 B.n74 B.t4 243.03
R377 B.n157 B.t15 243.03
R378 B.n151 B.t11 243.03
R379 B.n74 B.t6 182.798
R380 B.n157 B.t17 182.798
R381 B.n68 B.t9 182.798
R382 B.n151 B.t14 182.798
R383 B.n460 B.n458 163.367
R384 B.n456 B.n61 163.367
R385 B.n452 B.n450 163.367
R386 B.n448 B.n63 163.367
R387 B.n444 B.n442 163.367
R388 B.n440 B.n65 163.367
R389 B.n436 B.n434 163.367
R390 B.n432 B.n67 163.367
R391 B.n427 B.n425 163.367
R392 B.n423 B.n71 163.367
R393 B.n419 B.n417 163.367
R394 B.n415 B.n73 163.367
R395 B.n410 B.n408 163.367
R396 B.n406 B.n77 163.367
R397 B.n402 B.n400 163.367
R398 B.n398 B.n79 163.367
R399 B.n394 B.n392 163.367
R400 B.n390 B.n81 163.367
R401 B.n386 B.n384 163.367
R402 B.n382 B.n83 163.367
R403 B.n251 B.n138 163.367
R404 B.n255 B.n138 163.367
R405 B.n255 B.n132 163.367
R406 B.n263 B.n132 163.367
R407 B.n263 B.n130 163.367
R408 B.n267 B.n130 163.367
R409 B.n267 B.n125 163.367
R410 B.n276 B.n125 163.367
R411 B.n276 B.n123 163.367
R412 B.n280 B.n123 163.367
R413 B.n280 B.n117 163.367
R414 B.n288 B.n117 163.367
R415 B.n288 B.n115 163.367
R416 B.n292 B.n115 163.367
R417 B.n292 B.n108 163.367
R418 B.n300 B.n108 163.367
R419 B.n300 B.n106 163.367
R420 B.n304 B.n106 163.367
R421 B.n304 B.n101 163.367
R422 B.n312 B.n101 163.367
R423 B.n312 B.n99 163.367
R424 B.n316 B.n99 163.367
R425 B.n316 B.n92 163.367
R426 B.n324 B.n92 163.367
R427 B.n324 B.n90 163.367
R428 B.n329 B.n90 163.367
R429 B.n329 B.n85 163.367
R430 B.n337 B.n85 163.367
R431 B.n338 B.n337 163.367
R432 B.n338 B.n5 163.367
R433 B.n6 B.n5 163.367
R434 B.n7 B.n6 163.367
R435 B.n344 B.n7 163.367
R436 B.n345 B.n344 163.367
R437 B.n345 B.n13 163.367
R438 B.n14 B.n13 163.367
R439 B.n15 B.n14 163.367
R440 B.n350 B.n15 163.367
R441 B.n350 B.n20 163.367
R442 B.n21 B.n20 163.367
R443 B.n22 B.n21 163.367
R444 B.n355 B.n22 163.367
R445 B.n355 B.n27 163.367
R446 B.n28 B.n27 163.367
R447 B.n29 B.n28 163.367
R448 B.n360 B.n29 163.367
R449 B.n360 B.n34 163.367
R450 B.n35 B.n34 163.367
R451 B.n36 B.n35 163.367
R452 B.n365 B.n36 163.367
R453 B.n365 B.n41 163.367
R454 B.n42 B.n41 163.367
R455 B.n43 B.n42 163.367
R456 B.n370 B.n43 163.367
R457 B.n370 B.n48 163.367
R458 B.n49 B.n48 163.367
R459 B.n50 B.n49 163.367
R460 B.n375 B.n50 163.367
R461 B.n375 B.n55 163.367
R462 B.n56 B.n55 163.367
R463 B.n57 B.n56 163.367
R464 B.n245 B.n243 163.367
R465 B.n243 B.n242 163.367
R466 B.n239 B.n238 163.367
R467 B.n236 B.n146 163.367
R468 B.n232 B.n230 163.367
R469 B.n228 B.n148 163.367
R470 B.n224 B.n222 163.367
R471 B.n220 B.n150 163.367
R472 B.n215 B.n213 163.367
R473 B.n211 B.n154 163.367
R474 B.n207 B.n205 163.367
R475 B.n203 B.n156 163.367
R476 B.n199 B.n197 163.367
R477 B.n194 B.n193 163.367
R478 B.n191 B.n162 163.367
R479 B.n187 B.n185 163.367
R480 B.n183 B.n164 163.367
R481 B.n179 B.n177 163.367
R482 B.n175 B.n166 163.367
R483 B.n171 B.n169 163.367
R484 B.n249 B.n136 163.367
R485 B.n257 B.n136 163.367
R486 B.n257 B.n134 163.367
R487 B.n261 B.n134 163.367
R488 B.n261 B.n128 163.367
R489 B.n270 B.n128 163.367
R490 B.n270 B.n126 163.367
R491 B.n274 B.n126 163.367
R492 B.n274 B.n121 163.367
R493 B.n282 B.n121 163.367
R494 B.n282 B.n119 163.367
R495 B.n286 B.n119 163.367
R496 B.n286 B.n113 163.367
R497 B.n294 B.n113 163.367
R498 B.n294 B.n111 163.367
R499 B.n298 B.n111 163.367
R500 B.n298 B.n105 163.367
R501 B.n306 B.n105 163.367
R502 B.n306 B.n103 163.367
R503 B.n310 B.n103 163.367
R504 B.n310 B.n97 163.367
R505 B.n318 B.n97 163.367
R506 B.n318 B.n95 163.367
R507 B.n322 B.n95 163.367
R508 B.n322 B.n89 163.367
R509 B.n331 B.n89 163.367
R510 B.n331 B.n87 163.367
R511 B.n335 B.n87 163.367
R512 B.n335 B.n3 163.367
R513 B.n525 B.n3 163.367
R514 B.n521 B.n2 163.367
R515 B.n521 B.n520 163.367
R516 B.n520 B.n9 163.367
R517 B.n516 B.n9 163.367
R518 B.n516 B.n11 163.367
R519 B.n512 B.n11 163.367
R520 B.n512 B.n17 163.367
R521 B.n508 B.n17 163.367
R522 B.n508 B.n19 163.367
R523 B.n504 B.n19 163.367
R524 B.n504 B.n24 163.367
R525 B.n500 B.n24 163.367
R526 B.n500 B.n26 163.367
R527 B.n496 B.n26 163.367
R528 B.n496 B.n31 163.367
R529 B.n492 B.n31 163.367
R530 B.n492 B.n33 163.367
R531 B.n488 B.n33 163.367
R532 B.n488 B.n38 163.367
R533 B.n484 B.n38 163.367
R534 B.n484 B.n40 163.367
R535 B.n480 B.n40 163.367
R536 B.n480 B.n44 163.367
R537 B.n476 B.n44 163.367
R538 B.n476 B.n46 163.367
R539 B.n472 B.n46 163.367
R540 B.n472 B.n52 163.367
R541 B.n468 B.n52 163.367
R542 B.n468 B.n54 163.367
R543 B.n464 B.n54 163.367
R544 B.n250 B.n141 160.913
R545 B.n465 B.n58 160.913
R546 B.n75 B.t7 133.536
R547 B.n158 B.t16 133.536
R548 B.n69 B.t10 133.536
R549 B.n152 B.t13 133.536
R550 B.n250 B.n137 87.5371
R551 B.n256 B.n137 87.5371
R552 B.n256 B.n133 87.5371
R553 B.n262 B.n133 87.5371
R554 B.n262 B.n129 87.5371
R555 B.n269 B.n129 87.5371
R556 B.n269 B.n268 87.5371
R557 B.n275 B.n122 87.5371
R558 B.n281 B.n122 87.5371
R559 B.n281 B.n118 87.5371
R560 B.n287 B.n118 87.5371
R561 B.n287 B.n114 87.5371
R562 B.n293 B.n114 87.5371
R563 B.n293 B.n109 87.5371
R564 B.n299 B.n109 87.5371
R565 B.n299 B.n110 87.5371
R566 B.n305 B.n102 87.5371
R567 B.n311 B.n102 87.5371
R568 B.n311 B.n98 87.5371
R569 B.n317 B.n98 87.5371
R570 B.n317 B.n93 87.5371
R571 B.n323 B.n93 87.5371
R572 B.n323 B.n94 87.5371
R573 B.n330 B.n86 87.5371
R574 B.n336 B.n86 87.5371
R575 B.n336 B.n4 87.5371
R576 B.n524 B.n4 87.5371
R577 B.n524 B.n523 87.5371
R578 B.n523 B.n522 87.5371
R579 B.n522 B.n8 87.5371
R580 B.n12 B.n8 87.5371
R581 B.n515 B.n12 87.5371
R582 B.n514 B.n513 87.5371
R583 B.n513 B.n16 87.5371
R584 B.n507 B.n16 87.5371
R585 B.n507 B.n506 87.5371
R586 B.n506 B.n505 87.5371
R587 B.n505 B.n23 87.5371
R588 B.n499 B.n23 87.5371
R589 B.n498 B.n497 87.5371
R590 B.n497 B.n30 87.5371
R591 B.n491 B.n30 87.5371
R592 B.n491 B.n490 87.5371
R593 B.n490 B.n489 87.5371
R594 B.n489 B.n37 87.5371
R595 B.n483 B.n37 87.5371
R596 B.n483 B.n482 87.5371
R597 B.n482 B.n481 87.5371
R598 B.n475 B.n47 87.5371
R599 B.n475 B.n474 87.5371
R600 B.n474 B.n473 87.5371
R601 B.n473 B.n51 87.5371
R602 B.n467 B.n51 87.5371
R603 B.n467 B.n466 87.5371
R604 B.n466 B.n465 87.5371
R605 B.n275 B.t12 86.2498
R606 B.n481 B.t5 86.2498
R607 B.n330 B.t3 73.3767
R608 B.n515 B.t0 73.3767
R609 B.n459 B.n59 71.676
R610 B.n458 B.n457 71.676
R611 B.n451 B.n61 71.676
R612 B.n450 B.n449 71.676
R613 B.n443 B.n63 71.676
R614 B.n442 B.n441 71.676
R615 B.n435 B.n65 71.676
R616 B.n434 B.n433 71.676
R617 B.n426 B.n67 71.676
R618 B.n425 B.n424 71.676
R619 B.n418 B.n71 71.676
R620 B.n417 B.n416 71.676
R621 B.n409 B.n73 71.676
R622 B.n408 B.n407 71.676
R623 B.n401 B.n77 71.676
R624 B.n400 B.n399 71.676
R625 B.n393 B.n79 71.676
R626 B.n392 B.n391 71.676
R627 B.n385 B.n81 71.676
R628 B.n384 B.n383 71.676
R629 B.n383 B.n382 71.676
R630 B.n386 B.n385 71.676
R631 B.n391 B.n390 71.676
R632 B.n394 B.n393 71.676
R633 B.n399 B.n398 71.676
R634 B.n402 B.n401 71.676
R635 B.n407 B.n406 71.676
R636 B.n410 B.n409 71.676
R637 B.n416 B.n415 71.676
R638 B.n419 B.n418 71.676
R639 B.n424 B.n423 71.676
R640 B.n427 B.n426 71.676
R641 B.n433 B.n432 71.676
R642 B.n436 B.n435 71.676
R643 B.n441 B.n440 71.676
R644 B.n444 B.n443 71.676
R645 B.n449 B.n448 71.676
R646 B.n452 B.n451 71.676
R647 B.n457 B.n456 71.676
R648 B.n460 B.n459 71.676
R649 B.n244 B.n142 71.676
R650 B.n242 B.n144 71.676
R651 B.n238 B.n237 71.676
R652 B.n231 B.n146 71.676
R653 B.n230 B.n229 71.676
R654 B.n223 B.n148 71.676
R655 B.n222 B.n221 71.676
R656 B.n214 B.n150 71.676
R657 B.n213 B.n212 71.676
R658 B.n206 B.n154 71.676
R659 B.n205 B.n204 71.676
R660 B.n198 B.n156 71.676
R661 B.n197 B.n160 71.676
R662 B.n193 B.n192 71.676
R663 B.n186 B.n162 71.676
R664 B.n185 B.n184 71.676
R665 B.n178 B.n164 71.676
R666 B.n177 B.n176 71.676
R667 B.n170 B.n166 71.676
R668 B.n169 B.n168 71.676
R669 B.n245 B.n244 71.676
R670 B.n239 B.n144 71.676
R671 B.n237 B.n236 71.676
R672 B.n232 B.n231 71.676
R673 B.n229 B.n228 71.676
R674 B.n224 B.n223 71.676
R675 B.n221 B.n220 71.676
R676 B.n215 B.n214 71.676
R677 B.n212 B.n211 71.676
R678 B.n207 B.n206 71.676
R679 B.n204 B.n203 71.676
R680 B.n199 B.n198 71.676
R681 B.n194 B.n160 71.676
R682 B.n192 B.n191 71.676
R683 B.n187 B.n186 71.676
R684 B.n184 B.n183 71.676
R685 B.n179 B.n178 71.676
R686 B.n176 B.n175 71.676
R687 B.n171 B.n170 71.676
R688 B.n168 B.n140 71.676
R689 B.n526 B.n525 71.676
R690 B.n526 B.n2 71.676
R691 B.n110 B.t2 60.5037
R692 B.t1 B.n498 60.5037
R693 B.n430 B.n69 59.5399
R694 B.n412 B.n75 59.5399
R695 B.n159 B.n158 59.5399
R696 B.n217 B.n152 59.5399
R697 B.n69 B.n68 49.2611
R698 B.n75 B.n74 49.2611
R699 B.n158 B.n157 49.2611
R700 B.n152 B.n151 49.2611
R701 B.n248 B.n247 35.1225
R702 B.n252 B.n139 35.1225
R703 B.n380 B.n379 35.1225
R704 B.n463 B.n462 35.1225
R705 B.n305 B.t2 27.0339
R706 B.n499 B.t1 27.0339
R707 B B.n527 18.0485
R708 B.n94 B.t3 14.1608
R709 B.t0 B.n514 14.1608
R710 B.n248 B.n135 10.6151
R711 B.n258 B.n135 10.6151
R712 B.n259 B.n258 10.6151
R713 B.n260 B.n259 10.6151
R714 B.n260 B.n127 10.6151
R715 B.n271 B.n127 10.6151
R716 B.n272 B.n271 10.6151
R717 B.n273 B.n272 10.6151
R718 B.n273 B.n120 10.6151
R719 B.n283 B.n120 10.6151
R720 B.n284 B.n283 10.6151
R721 B.n285 B.n284 10.6151
R722 B.n285 B.n112 10.6151
R723 B.n295 B.n112 10.6151
R724 B.n296 B.n295 10.6151
R725 B.n297 B.n296 10.6151
R726 B.n297 B.n104 10.6151
R727 B.n307 B.n104 10.6151
R728 B.n308 B.n307 10.6151
R729 B.n309 B.n308 10.6151
R730 B.n309 B.n96 10.6151
R731 B.n319 B.n96 10.6151
R732 B.n320 B.n319 10.6151
R733 B.n321 B.n320 10.6151
R734 B.n321 B.n88 10.6151
R735 B.n332 B.n88 10.6151
R736 B.n333 B.n332 10.6151
R737 B.n334 B.n333 10.6151
R738 B.n334 B.n0 10.6151
R739 B.n247 B.n246 10.6151
R740 B.n246 B.n143 10.6151
R741 B.n241 B.n143 10.6151
R742 B.n241 B.n240 10.6151
R743 B.n240 B.n145 10.6151
R744 B.n235 B.n145 10.6151
R745 B.n235 B.n234 10.6151
R746 B.n234 B.n233 10.6151
R747 B.n233 B.n147 10.6151
R748 B.n227 B.n147 10.6151
R749 B.n227 B.n226 10.6151
R750 B.n226 B.n225 10.6151
R751 B.n225 B.n149 10.6151
R752 B.n219 B.n149 10.6151
R753 B.n219 B.n218 10.6151
R754 B.n216 B.n153 10.6151
R755 B.n210 B.n153 10.6151
R756 B.n210 B.n209 10.6151
R757 B.n209 B.n208 10.6151
R758 B.n208 B.n155 10.6151
R759 B.n202 B.n155 10.6151
R760 B.n202 B.n201 10.6151
R761 B.n201 B.n200 10.6151
R762 B.n196 B.n195 10.6151
R763 B.n195 B.n161 10.6151
R764 B.n190 B.n161 10.6151
R765 B.n190 B.n189 10.6151
R766 B.n189 B.n188 10.6151
R767 B.n188 B.n163 10.6151
R768 B.n182 B.n163 10.6151
R769 B.n182 B.n181 10.6151
R770 B.n181 B.n180 10.6151
R771 B.n180 B.n165 10.6151
R772 B.n174 B.n165 10.6151
R773 B.n174 B.n173 10.6151
R774 B.n173 B.n172 10.6151
R775 B.n172 B.n167 10.6151
R776 B.n167 B.n139 10.6151
R777 B.n253 B.n252 10.6151
R778 B.n254 B.n253 10.6151
R779 B.n254 B.n131 10.6151
R780 B.n264 B.n131 10.6151
R781 B.n265 B.n264 10.6151
R782 B.n266 B.n265 10.6151
R783 B.n266 B.n124 10.6151
R784 B.n277 B.n124 10.6151
R785 B.n278 B.n277 10.6151
R786 B.n279 B.n278 10.6151
R787 B.n279 B.n116 10.6151
R788 B.n289 B.n116 10.6151
R789 B.n290 B.n289 10.6151
R790 B.n291 B.n290 10.6151
R791 B.n291 B.n107 10.6151
R792 B.n301 B.n107 10.6151
R793 B.n302 B.n301 10.6151
R794 B.n303 B.n302 10.6151
R795 B.n303 B.n100 10.6151
R796 B.n313 B.n100 10.6151
R797 B.n314 B.n313 10.6151
R798 B.n315 B.n314 10.6151
R799 B.n315 B.n91 10.6151
R800 B.n325 B.n91 10.6151
R801 B.n326 B.n325 10.6151
R802 B.n328 B.n326 10.6151
R803 B.n328 B.n327 10.6151
R804 B.n327 B.n84 10.6151
R805 B.n339 B.n84 10.6151
R806 B.n340 B.n339 10.6151
R807 B.n341 B.n340 10.6151
R808 B.n342 B.n341 10.6151
R809 B.n343 B.n342 10.6151
R810 B.n346 B.n343 10.6151
R811 B.n347 B.n346 10.6151
R812 B.n348 B.n347 10.6151
R813 B.n349 B.n348 10.6151
R814 B.n351 B.n349 10.6151
R815 B.n352 B.n351 10.6151
R816 B.n353 B.n352 10.6151
R817 B.n354 B.n353 10.6151
R818 B.n356 B.n354 10.6151
R819 B.n357 B.n356 10.6151
R820 B.n358 B.n357 10.6151
R821 B.n359 B.n358 10.6151
R822 B.n361 B.n359 10.6151
R823 B.n362 B.n361 10.6151
R824 B.n363 B.n362 10.6151
R825 B.n364 B.n363 10.6151
R826 B.n366 B.n364 10.6151
R827 B.n367 B.n366 10.6151
R828 B.n368 B.n367 10.6151
R829 B.n369 B.n368 10.6151
R830 B.n371 B.n369 10.6151
R831 B.n372 B.n371 10.6151
R832 B.n373 B.n372 10.6151
R833 B.n374 B.n373 10.6151
R834 B.n376 B.n374 10.6151
R835 B.n377 B.n376 10.6151
R836 B.n378 B.n377 10.6151
R837 B.n379 B.n378 10.6151
R838 B.n519 B.n1 10.6151
R839 B.n519 B.n518 10.6151
R840 B.n518 B.n517 10.6151
R841 B.n517 B.n10 10.6151
R842 B.n511 B.n10 10.6151
R843 B.n511 B.n510 10.6151
R844 B.n510 B.n509 10.6151
R845 B.n509 B.n18 10.6151
R846 B.n503 B.n18 10.6151
R847 B.n503 B.n502 10.6151
R848 B.n502 B.n501 10.6151
R849 B.n501 B.n25 10.6151
R850 B.n495 B.n25 10.6151
R851 B.n495 B.n494 10.6151
R852 B.n494 B.n493 10.6151
R853 B.n493 B.n32 10.6151
R854 B.n487 B.n32 10.6151
R855 B.n487 B.n486 10.6151
R856 B.n486 B.n485 10.6151
R857 B.n485 B.n39 10.6151
R858 B.n479 B.n39 10.6151
R859 B.n479 B.n478 10.6151
R860 B.n478 B.n477 10.6151
R861 B.n477 B.n45 10.6151
R862 B.n471 B.n45 10.6151
R863 B.n471 B.n470 10.6151
R864 B.n470 B.n469 10.6151
R865 B.n469 B.n53 10.6151
R866 B.n463 B.n53 10.6151
R867 B.n462 B.n461 10.6151
R868 B.n461 B.n60 10.6151
R869 B.n455 B.n60 10.6151
R870 B.n455 B.n454 10.6151
R871 B.n454 B.n453 10.6151
R872 B.n453 B.n62 10.6151
R873 B.n447 B.n62 10.6151
R874 B.n447 B.n446 10.6151
R875 B.n446 B.n445 10.6151
R876 B.n445 B.n64 10.6151
R877 B.n439 B.n64 10.6151
R878 B.n439 B.n438 10.6151
R879 B.n438 B.n437 10.6151
R880 B.n437 B.n66 10.6151
R881 B.n431 B.n66 10.6151
R882 B.n429 B.n428 10.6151
R883 B.n428 B.n70 10.6151
R884 B.n422 B.n70 10.6151
R885 B.n422 B.n421 10.6151
R886 B.n421 B.n420 10.6151
R887 B.n420 B.n72 10.6151
R888 B.n414 B.n72 10.6151
R889 B.n414 B.n413 10.6151
R890 B.n411 B.n76 10.6151
R891 B.n405 B.n76 10.6151
R892 B.n405 B.n404 10.6151
R893 B.n404 B.n403 10.6151
R894 B.n403 B.n78 10.6151
R895 B.n397 B.n78 10.6151
R896 B.n397 B.n396 10.6151
R897 B.n396 B.n395 10.6151
R898 B.n395 B.n80 10.6151
R899 B.n389 B.n80 10.6151
R900 B.n389 B.n388 10.6151
R901 B.n388 B.n387 10.6151
R902 B.n387 B.n82 10.6151
R903 B.n381 B.n82 10.6151
R904 B.n381 B.n380 10.6151
R905 B.n527 B.n0 8.11757
R906 B.n527 B.n1 8.11757
R907 B.n217 B.n216 6.5566
R908 B.n200 B.n159 6.5566
R909 B.n430 B.n429 6.5566
R910 B.n413 B.n412 6.5566
R911 B.n218 B.n217 4.05904
R912 B.n196 B.n159 4.05904
R913 B.n431 B.n430 4.05904
R914 B.n412 B.n411 4.05904
R915 B.n268 B.t12 1.2878
R916 B.n47 B.t5 1.2878
R917 VP.n12 VP.n0 161.3
R918 VP.n11 VP.n10 161.3
R919 VP.n9 VP.n1 161.3
R920 VP.n8 VP.n7 161.3
R921 VP.n6 VP.n2 161.3
R922 VP.n5 VP.n4 97.5443
R923 VP.n14 VP.n13 97.5443
R924 VP.n3 VP.t3 71.4101
R925 VP.n3 VP.t2 70.7721
R926 VP.n4 VP.n3 44.2426
R927 VP.n7 VP.n1 40.4934
R928 VP.n11 VP.n1 40.4934
R929 VP.n5 VP.t0 35.6598
R930 VP.n13 VP.t1 35.6598
R931 VP.n7 VP.n6 24.4675
R932 VP.n12 VP.n11 24.4675
R933 VP.n6 VP.n5 13.2127
R934 VP.n13 VP.n12 13.2127
R935 VP.n4 VP.n2 0.278367
R936 VP.n14 VP.n0 0.278367
R937 VP.n8 VP.n2 0.189894
R938 VP.n9 VP.n8 0.189894
R939 VP.n10 VP.n9 0.189894
R940 VP.n10 VP.n0 0.189894
R941 VP VP.n14 0.153454
R942 VDD1 VDD1.n1 114.285
R943 VDD1 VDD1.n0 80.7164
R944 VDD1.n0 VDD1.t1 6.05555
R945 VDD1.n0 VDD1.t0 6.05555
R946 VDD1.n1 VDD1.t3 6.05555
R947 VDD1.n1 VDD1.t2 6.05555
R948 VTAIL.n122 VTAIL.n112 289.615
R949 VTAIL.n10 VTAIL.n0 289.615
R950 VTAIL.n26 VTAIL.n16 289.615
R951 VTAIL.n42 VTAIL.n32 289.615
R952 VTAIL.n106 VTAIL.n96 289.615
R953 VTAIL.n90 VTAIL.n80 289.615
R954 VTAIL.n74 VTAIL.n64 289.615
R955 VTAIL.n58 VTAIL.n48 289.615
R956 VTAIL.n116 VTAIL.n115 185
R957 VTAIL.n121 VTAIL.n120 185
R958 VTAIL.n123 VTAIL.n122 185
R959 VTAIL.n4 VTAIL.n3 185
R960 VTAIL.n9 VTAIL.n8 185
R961 VTAIL.n11 VTAIL.n10 185
R962 VTAIL.n20 VTAIL.n19 185
R963 VTAIL.n25 VTAIL.n24 185
R964 VTAIL.n27 VTAIL.n26 185
R965 VTAIL.n36 VTAIL.n35 185
R966 VTAIL.n41 VTAIL.n40 185
R967 VTAIL.n43 VTAIL.n42 185
R968 VTAIL.n107 VTAIL.n106 185
R969 VTAIL.n105 VTAIL.n104 185
R970 VTAIL.n100 VTAIL.n99 185
R971 VTAIL.n91 VTAIL.n90 185
R972 VTAIL.n89 VTAIL.n88 185
R973 VTAIL.n84 VTAIL.n83 185
R974 VTAIL.n75 VTAIL.n74 185
R975 VTAIL.n73 VTAIL.n72 185
R976 VTAIL.n68 VTAIL.n67 185
R977 VTAIL.n59 VTAIL.n58 185
R978 VTAIL.n57 VTAIL.n56 185
R979 VTAIL.n52 VTAIL.n51 185
R980 VTAIL.n117 VTAIL.t1 148.606
R981 VTAIL.n5 VTAIL.t3 148.606
R982 VTAIL.n21 VTAIL.t6 148.606
R983 VTAIL.n37 VTAIL.t7 148.606
R984 VTAIL.n101 VTAIL.t5 148.606
R985 VTAIL.n85 VTAIL.t4 148.606
R986 VTAIL.n69 VTAIL.t0 148.606
R987 VTAIL.n53 VTAIL.t2 148.606
R988 VTAIL.n121 VTAIL.n115 104.615
R989 VTAIL.n122 VTAIL.n121 104.615
R990 VTAIL.n9 VTAIL.n3 104.615
R991 VTAIL.n10 VTAIL.n9 104.615
R992 VTAIL.n25 VTAIL.n19 104.615
R993 VTAIL.n26 VTAIL.n25 104.615
R994 VTAIL.n41 VTAIL.n35 104.615
R995 VTAIL.n42 VTAIL.n41 104.615
R996 VTAIL.n106 VTAIL.n105 104.615
R997 VTAIL.n105 VTAIL.n99 104.615
R998 VTAIL.n90 VTAIL.n89 104.615
R999 VTAIL.n89 VTAIL.n83 104.615
R1000 VTAIL.n74 VTAIL.n73 104.615
R1001 VTAIL.n73 VTAIL.n67 104.615
R1002 VTAIL.n58 VTAIL.n57 104.615
R1003 VTAIL.n57 VTAIL.n51 104.615
R1004 VTAIL.t1 VTAIL.n115 52.3082
R1005 VTAIL.t3 VTAIL.n3 52.3082
R1006 VTAIL.t6 VTAIL.n19 52.3082
R1007 VTAIL.t7 VTAIL.n35 52.3082
R1008 VTAIL.t5 VTAIL.n99 52.3082
R1009 VTAIL.t4 VTAIL.n83 52.3082
R1010 VTAIL.t0 VTAIL.n67 52.3082
R1011 VTAIL.t2 VTAIL.n51 52.3082
R1012 VTAIL.n127 VTAIL.n126 35.0944
R1013 VTAIL.n15 VTAIL.n14 35.0944
R1014 VTAIL.n31 VTAIL.n30 35.0944
R1015 VTAIL.n47 VTAIL.n46 35.0944
R1016 VTAIL.n111 VTAIL.n110 35.0944
R1017 VTAIL.n95 VTAIL.n94 35.0944
R1018 VTAIL.n79 VTAIL.n78 35.0944
R1019 VTAIL.n63 VTAIL.n62 35.0944
R1020 VTAIL.n127 VTAIL.n111 17.3755
R1021 VTAIL.n63 VTAIL.n47 17.3755
R1022 VTAIL.n117 VTAIL.n116 15.5966
R1023 VTAIL.n5 VTAIL.n4 15.5966
R1024 VTAIL.n21 VTAIL.n20 15.5966
R1025 VTAIL.n37 VTAIL.n36 15.5966
R1026 VTAIL.n101 VTAIL.n100 15.5966
R1027 VTAIL.n85 VTAIL.n84 15.5966
R1028 VTAIL.n69 VTAIL.n68 15.5966
R1029 VTAIL.n53 VTAIL.n52 15.5966
R1030 VTAIL.n120 VTAIL.n119 12.8005
R1031 VTAIL.n8 VTAIL.n7 12.8005
R1032 VTAIL.n24 VTAIL.n23 12.8005
R1033 VTAIL.n40 VTAIL.n39 12.8005
R1034 VTAIL.n104 VTAIL.n103 12.8005
R1035 VTAIL.n88 VTAIL.n87 12.8005
R1036 VTAIL.n72 VTAIL.n71 12.8005
R1037 VTAIL.n56 VTAIL.n55 12.8005
R1038 VTAIL.n123 VTAIL.n114 12.0247
R1039 VTAIL.n11 VTAIL.n2 12.0247
R1040 VTAIL.n27 VTAIL.n18 12.0247
R1041 VTAIL.n43 VTAIL.n34 12.0247
R1042 VTAIL.n107 VTAIL.n98 12.0247
R1043 VTAIL.n91 VTAIL.n82 12.0247
R1044 VTAIL.n75 VTAIL.n66 12.0247
R1045 VTAIL.n59 VTAIL.n50 12.0247
R1046 VTAIL.n124 VTAIL.n112 11.249
R1047 VTAIL.n12 VTAIL.n0 11.249
R1048 VTAIL.n28 VTAIL.n16 11.249
R1049 VTAIL.n44 VTAIL.n32 11.249
R1050 VTAIL.n108 VTAIL.n96 11.249
R1051 VTAIL.n92 VTAIL.n80 11.249
R1052 VTAIL.n76 VTAIL.n64 11.249
R1053 VTAIL.n60 VTAIL.n48 11.249
R1054 VTAIL.n126 VTAIL.n125 9.45567
R1055 VTAIL.n14 VTAIL.n13 9.45567
R1056 VTAIL.n30 VTAIL.n29 9.45567
R1057 VTAIL.n46 VTAIL.n45 9.45567
R1058 VTAIL.n110 VTAIL.n109 9.45567
R1059 VTAIL.n94 VTAIL.n93 9.45567
R1060 VTAIL.n78 VTAIL.n77 9.45567
R1061 VTAIL.n62 VTAIL.n61 9.45567
R1062 VTAIL.n125 VTAIL.n124 9.3005
R1063 VTAIL.n114 VTAIL.n113 9.3005
R1064 VTAIL.n119 VTAIL.n118 9.3005
R1065 VTAIL.n13 VTAIL.n12 9.3005
R1066 VTAIL.n2 VTAIL.n1 9.3005
R1067 VTAIL.n7 VTAIL.n6 9.3005
R1068 VTAIL.n29 VTAIL.n28 9.3005
R1069 VTAIL.n18 VTAIL.n17 9.3005
R1070 VTAIL.n23 VTAIL.n22 9.3005
R1071 VTAIL.n45 VTAIL.n44 9.3005
R1072 VTAIL.n34 VTAIL.n33 9.3005
R1073 VTAIL.n39 VTAIL.n38 9.3005
R1074 VTAIL.n109 VTAIL.n108 9.3005
R1075 VTAIL.n98 VTAIL.n97 9.3005
R1076 VTAIL.n103 VTAIL.n102 9.3005
R1077 VTAIL.n93 VTAIL.n92 9.3005
R1078 VTAIL.n82 VTAIL.n81 9.3005
R1079 VTAIL.n87 VTAIL.n86 9.3005
R1080 VTAIL.n77 VTAIL.n76 9.3005
R1081 VTAIL.n66 VTAIL.n65 9.3005
R1082 VTAIL.n71 VTAIL.n70 9.3005
R1083 VTAIL.n61 VTAIL.n60 9.3005
R1084 VTAIL.n50 VTAIL.n49 9.3005
R1085 VTAIL.n55 VTAIL.n54 9.3005
R1086 VTAIL.n118 VTAIL.n117 4.46457
R1087 VTAIL.n6 VTAIL.n5 4.46457
R1088 VTAIL.n22 VTAIL.n21 4.46457
R1089 VTAIL.n38 VTAIL.n37 4.46457
R1090 VTAIL.n102 VTAIL.n101 4.46457
R1091 VTAIL.n86 VTAIL.n85 4.46457
R1092 VTAIL.n70 VTAIL.n69 4.46457
R1093 VTAIL.n54 VTAIL.n53 4.46457
R1094 VTAIL.n126 VTAIL.n112 2.71565
R1095 VTAIL.n14 VTAIL.n0 2.71565
R1096 VTAIL.n30 VTAIL.n16 2.71565
R1097 VTAIL.n46 VTAIL.n32 2.71565
R1098 VTAIL.n110 VTAIL.n96 2.71565
R1099 VTAIL.n94 VTAIL.n80 2.71565
R1100 VTAIL.n78 VTAIL.n64 2.71565
R1101 VTAIL.n62 VTAIL.n48 2.71565
R1102 VTAIL.n79 VTAIL.n63 2.19016
R1103 VTAIL.n111 VTAIL.n95 2.19016
R1104 VTAIL.n47 VTAIL.n31 2.19016
R1105 VTAIL.n124 VTAIL.n123 1.93989
R1106 VTAIL.n12 VTAIL.n11 1.93989
R1107 VTAIL.n28 VTAIL.n27 1.93989
R1108 VTAIL.n44 VTAIL.n43 1.93989
R1109 VTAIL.n108 VTAIL.n107 1.93989
R1110 VTAIL.n92 VTAIL.n91 1.93989
R1111 VTAIL.n76 VTAIL.n75 1.93989
R1112 VTAIL.n60 VTAIL.n59 1.93989
R1113 VTAIL.n120 VTAIL.n114 1.16414
R1114 VTAIL.n8 VTAIL.n2 1.16414
R1115 VTAIL.n24 VTAIL.n18 1.16414
R1116 VTAIL.n40 VTAIL.n34 1.16414
R1117 VTAIL.n104 VTAIL.n98 1.16414
R1118 VTAIL.n88 VTAIL.n82 1.16414
R1119 VTAIL.n72 VTAIL.n66 1.16414
R1120 VTAIL.n56 VTAIL.n50 1.16414
R1121 VTAIL VTAIL.n15 1.15352
R1122 VTAIL VTAIL.n127 1.03714
R1123 VTAIL.n95 VTAIL.n79 0.470328
R1124 VTAIL.n31 VTAIL.n15 0.470328
R1125 VTAIL.n119 VTAIL.n116 0.388379
R1126 VTAIL.n7 VTAIL.n4 0.388379
R1127 VTAIL.n23 VTAIL.n20 0.388379
R1128 VTAIL.n39 VTAIL.n36 0.388379
R1129 VTAIL.n103 VTAIL.n100 0.388379
R1130 VTAIL.n87 VTAIL.n84 0.388379
R1131 VTAIL.n71 VTAIL.n68 0.388379
R1132 VTAIL.n55 VTAIL.n52 0.388379
R1133 VTAIL.n118 VTAIL.n113 0.155672
R1134 VTAIL.n125 VTAIL.n113 0.155672
R1135 VTAIL.n6 VTAIL.n1 0.155672
R1136 VTAIL.n13 VTAIL.n1 0.155672
R1137 VTAIL.n22 VTAIL.n17 0.155672
R1138 VTAIL.n29 VTAIL.n17 0.155672
R1139 VTAIL.n38 VTAIL.n33 0.155672
R1140 VTAIL.n45 VTAIL.n33 0.155672
R1141 VTAIL.n109 VTAIL.n97 0.155672
R1142 VTAIL.n102 VTAIL.n97 0.155672
R1143 VTAIL.n93 VTAIL.n81 0.155672
R1144 VTAIL.n86 VTAIL.n81 0.155672
R1145 VTAIL.n77 VTAIL.n65 0.155672
R1146 VTAIL.n70 VTAIL.n65 0.155672
R1147 VTAIL.n61 VTAIL.n49 0.155672
R1148 VTAIL.n54 VTAIL.n49 0.155672
R1149 VN.n0 VN.t2 71.4101
R1150 VN.n1 VN.t3 71.4101
R1151 VN.n0 VN.t0 70.7721
R1152 VN.n1 VN.t1 70.7721
R1153 VN VN.n1 44.5214
R1154 VN VN.n0 5.8131
R1155 VDD2.n2 VDD2.n0 113.76
R1156 VDD2.n2 VDD2.n1 80.6582
R1157 VDD2.n1 VDD2.t2 6.05555
R1158 VDD2.n1 VDD2.t0 6.05555
R1159 VDD2.n0 VDD2.t1 6.05555
R1160 VDD2.n0 VDD2.t3 6.05555
R1161 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 1.85717f
C1 VTAIL VDD1 3.15688f
C2 VDD1 VN 0.153189f
C3 VDD2 VTAIL 3.20847f
C4 VDD2 VN 1.48972f
C5 VDD2 VDD1 0.93437f
C6 VP VTAIL 1.87128f
C7 VP VN 4.30212f
C8 VP VDD1 1.70987f
C9 VP VDD2 0.374567f
C10 VDD2 B 2.793118f
C11 VDD1 B 4.95842f
C12 VTAIL B 4.321012f
C13 VN B 8.462637f
C14 VP B 7.339375f
C15 VDD2.t1 B 0.049307f
C16 VDD2.t3 B 0.049307f
C17 VDD2.n0 B 0.59215f
C18 VDD2.t2 B 0.049307f
C19 VDD2.t0 B 0.049307f
C20 VDD2.n1 B 0.372099f
C21 VDD2.n2 B 1.89978f
C22 VN.t2 B 0.479752f
C23 VN.t0 B 0.477468f
C24 VN.n0 B 0.316587f
C25 VN.t3 B 0.479752f
C26 VN.t1 B 0.477468f
C27 VN.n1 B 1.0706f
C28 VTAIL.n0 B 0.020166f
C29 VTAIL.n1 B 0.014416f
C30 VTAIL.n2 B 0.007746f
C31 VTAIL.n3 B 0.013732f
C32 VTAIL.n4 B 0.010677f
C33 VTAIL.t3 B 0.031073f
C34 VTAIL.n5 B 0.053954f
C35 VTAIL.n6 B 0.159288f
C36 VTAIL.n7 B 0.007746f
C37 VTAIL.n8 B 0.008202f
C38 VTAIL.n9 B 0.01831f
C39 VTAIL.n10 B 0.039466f
C40 VTAIL.n11 B 0.008202f
C41 VTAIL.n12 B 0.007746f
C42 VTAIL.n13 B 0.036276f
C43 VTAIL.n14 B 0.022152f
C44 VTAIL.n15 B 0.089366f
C45 VTAIL.n16 B 0.020166f
C46 VTAIL.n17 B 0.014416f
C47 VTAIL.n18 B 0.007746f
C48 VTAIL.n19 B 0.013732f
C49 VTAIL.n20 B 0.010677f
C50 VTAIL.t6 B 0.031073f
C51 VTAIL.n21 B 0.053954f
C52 VTAIL.n22 B 0.159288f
C53 VTAIL.n23 B 0.007746f
C54 VTAIL.n24 B 0.008202f
C55 VTAIL.n25 B 0.01831f
C56 VTAIL.n26 B 0.039466f
C57 VTAIL.n27 B 0.008202f
C58 VTAIL.n28 B 0.007746f
C59 VTAIL.n29 B 0.036276f
C60 VTAIL.n30 B 0.022152f
C61 VTAIL.n31 B 0.137519f
C62 VTAIL.n32 B 0.020166f
C63 VTAIL.n33 B 0.014416f
C64 VTAIL.n34 B 0.007746f
C65 VTAIL.n35 B 0.013732f
C66 VTAIL.n36 B 0.010677f
C67 VTAIL.t7 B 0.031073f
C68 VTAIL.n37 B 0.053954f
C69 VTAIL.n38 B 0.159288f
C70 VTAIL.n39 B 0.007746f
C71 VTAIL.n40 B 0.008202f
C72 VTAIL.n41 B 0.01831f
C73 VTAIL.n42 B 0.039466f
C74 VTAIL.n43 B 0.008202f
C75 VTAIL.n44 B 0.007746f
C76 VTAIL.n45 B 0.036276f
C77 VTAIL.n46 B 0.022152f
C78 VTAIL.n47 B 0.544175f
C79 VTAIL.n48 B 0.020166f
C80 VTAIL.n49 B 0.014416f
C81 VTAIL.n50 B 0.007746f
C82 VTAIL.n51 B 0.013732f
C83 VTAIL.n52 B 0.010677f
C84 VTAIL.t2 B 0.031073f
C85 VTAIL.n53 B 0.053954f
C86 VTAIL.n54 B 0.159288f
C87 VTAIL.n55 B 0.007746f
C88 VTAIL.n56 B 0.008202f
C89 VTAIL.n57 B 0.01831f
C90 VTAIL.n58 B 0.039466f
C91 VTAIL.n59 B 0.008202f
C92 VTAIL.n60 B 0.007746f
C93 VTAIL.n61 B 0.036276f
C94 VTAIL.n62 B 0.022152f
C95 VTAIL.n63 B 0.544175f
C96 VTAIL.n64 B 0.020166f
C97 VTAIL.n65 B 0.014416f
C98 VTAIL.n66 B 0.007746f
C99 VTAIL.n67 B 0.013732f
C100 VTAIL.n68 B 0.010677f
C101 VTAIL.t0 B 0.031073f
C102 VTAIL.n69 B 0.053954f
C103 VTAIL.n70 B 0.159288f
C104 VTAIL.n71 B 0.007746f
C105 VTAIL.n72 B 0.008202f
C106 VTAIL.n73 B 0.01831f
C107 VTAIL.n74 B 0.039466f
C108 VTAIL.n75 B 0.008202f
C109 VTAIL.n76 B 0.007746f
C110 VTAIL.n77 B 0.036276f
C111 VTAIL.n78 B 0.022152f
C112 VTAIL.n79 B 0.137519f
C113 VTAIL.n80 B 0.020166f
C114 VTAIL.n81 B 0.014416f
C115 VTAIL.n82 B 0.007746f
C116 VTAIL.n83 B 0.013732f
C117 VTAIL.n84 B 0.010677f
C118 VTAIL.t4 B 0.031073f
C119 VTAIL.n85 B 0.053954f
C120 VTAIL.n86 B 0.159288f
C121 VTAIL.n87 B 0.007746f
C122 VTAIL.n88 B 0.008202f
C123 VTAIL.n89 B 0.01831f
C124 VTAIL.n90 B 0.039466f
C125 VTAIL.n91 B 0.008202f
C126 VTAIL.n92 B 0.007746f
C127 VTAIL.n93 B 0.036276f
C128 VTAIL.n94 B 0.022152f
C129 VTAIL.n95 B 0.137519f
C130 VTAIL.n96 B 0.020166f
C131 VTAIL.n97 B 0.014416f
C132 VTAIL.n98 B 0.007746f
C133 VTAIL.n99 B 0.013732f
C134 VTAIL.n100 B 0.010677f
C135 VTAIL.t5 B 0.031073f
C136 VTAIL.n101 B 0.053954f
C137 VTAIL.n102 B 0.159288f
C138 VTAIL.n103 B 0.007746f
C139 VTAIL.n104 B 0.008202f
C140 VTAIL.n105 B 0.01831f
C141 VTAIL.n106 B 0.039466f
C142 VTAIL.n107 B 0.008202f
C143 VTAIL.n108 B 0.007746f
C144 VTAIL.n109 B 0.036276f
C145 VTAIL.n110 B 0.022152f
C146 VTAIL.n111 B 0.544175f
C147 VTAIL.n112 B 0.020166f
C148 VTAIL.n113 B 0.014416f
C149 VTAIL.n114 B 0.007746f
C150 VTAIL.n115 B 0.013732f
C151 VTAIL.n116 B 0.010677f
C152 VTAIL.t1 B 0.031073f
C153 VTAIL.n117 B 0.053954f
C154 VTAIL.n118 B 0.159288f
C155 VTAIL.n119 B 0.007746f
C156 VTAIL.n120 B 0.008202f
C157 VTAIL.n121 B 0.01831f
C158 VTAIL.n122 B 0.039466f
C159 VTAIL.n123 B 0.008202f
C160 VTAIL.n124 B 0.007746f
C161 VTAIL.n125 B 0.036276f
C162 VTAIL.n126 B 0.022152f
C163 VTAIL.n127 B 0.490616f
C164 VDD1.t1 B 0.048245f
C165 VDD1.t0 B 0.048245f
C166 VDD1.n0 B 0.364286f
C167 VDD1.t3 B 0.048245f
C168 VDD1.t2 B 0.048245f
C169 VDD1.n1 B 0.592956f
C170 VP.n0 B 0.025599f
C171 VP.t1 B 0.353152f
C172 VP.n1 B 0.015697f
C173 VP.n2 B 0.025599f
C174 VP.t0 B 0.353152f
C175 VP.t2 B 0.480498f
C176 VP.t3 B 0.482797f
C177 VP.n3 B 1.06716f
C178 VP.n4 B 0.841641f
C179 VP.n5 B 0.207081f
C180 VP.n6 B 0.027969f
C181 VP.n7 B 0.03859f
C182 VP.n8 B 0.019417f
C183 VP.n9 B 0.019417f
C184 VP.n10 B 0.019417f
C185 VP.n11 B 0.03859f
C186 VP.n12 B 0.027969f
C187 VP.n13 B 0.207081f
C188 VP.n14 B 0.027835f
.ends

