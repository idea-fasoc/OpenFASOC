* NGSPICE file created from diff_pair_sample_1380.ext - technology: sky130A

.subckt diff_pair_sample_1380 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=0 ps=0 w=12.17 l=1.59
X1 B.t8 B.t6 B.t7 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=0 ps=0 w=12.17 l=1.59
X2 VTAIL.t7 VP.t0 VDD1.t0 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=2.00805 ps=12.5 w=12.17 l=1.59
X3 B.t5 B.t3 B.t4 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=0 ps=0 w=12.17 l=1.59
X4 VDD1.t1 VP.t1 VTAIL.t6 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=2.00805 pd=12.5 as=4.7463 ps=25.12 w=12.17 l=1.59
X5 VDD2.t3 VN.t0 VTAIL.t2 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=2.00805 pd=12.5 as=4.7463 ps=25.12 w=12.17 l=1.59
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=2.00805 pd=12.5 as=4.7463 ps=25.12 w=12.17 l=1.59
X7 VTAIL.t0 VN.t2 VDD2.t1 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=2.00805 ps=12.5 w=12.17 l=1.59
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=2.00805 ps=12.5 w=12.17 l=1.59
X9 VDD1.t2 VP.t2 VTAIL.t5 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=2.00805 pd=12.5 as=4.7463 ps=25.12 w=12.17 l=1.59
X10 VTAIL.t4 VP.t3 VDD1.t3 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=2.00805 ps=12.5 w=12.17 l=1.59
X11 B.t2 B.t0 B.t1 w_n2122_n3402# sky130_fd_pr__pfet_01v8 ad=4.7463 pd=25.12 as=0 ps=0 w=12.17 l=1.59
R0 B.n411 B.n66 585
R1 B.n413 B.n412 585
R2 B.n414 B.n65 585
R3 B.n416 B.n415 585
R4 B.n417 B.n64 585
R5 B.n419 B.n418 585
R6 B.n420 B.n63 585
R7 B.n422 B.n421 585
R8 B.n423 B.n62 585
R9 B.n425 B.n424 585
R10 B.n426 B.n61 585
R11 B.n428 B.n427 585
R12 B.n429 B.n60 585
R13 B.n431 B.n430 585
R14 B.n432 B.n59 585
R15 B.n434 B.n433 585
R16 B.n435 B.n58 585
R17 B.n437 B.n436 585
R18 B.n438 B.n57 585
R19 B.n440 B.n439 585
R20 B.n441 B.n56 585
R21 B.n443 B.n442 585
R22 B.n444 B.n55 585
R23 B.n446 B.n445 585
R24 B.n447 B.n54 585
R25 B.n449 B.n448 585
R26 B.n450 B.n53 585
R27 B.n452 B.n451 585
R28 B.n453 B.n52 585
R29 B.n455 B.n454 585
R30 B.n456 B.n51 585
R31 B.n458 B.n457 585
R32 B.n459 B.n50 585
R33 B.n461 B.n460 585
R34 B.n462 B.n49 585
R35 B.n464 B.n463 585
R36 B.n465 B.n48 585
R37 B.n467 B.n466 585
R38 B.n468 B.n47 585
R39 B.n470 B.n469 585
R40 B.n471 B.n43 585
R41 B.n473 B.n472 585
R42 B.n474 B.n42 585
R43 B.n476 B.n475 585
R44 B.n477 B.n41 585
R45 B.n479 B.n478 585
R46 B.n480 B.n40 585
R47 B.n482 B.n481 585
R48 B.n483 B.n39 585
R49 B.n485 B.n484 585
R50 B.n486 B.n38 585
R51 B.n488 B.n487 585
R52 B.n490 B.n35 585
R53 B.n492 B.n491 585
R54 B.n493 B.n34 585
R55 B.n495 B.n494 585
R56 B.n496 B.n33 585
R57 B.n498 B.n497 585
R58 B.n499 B.n32 585
R59 B.n501 B.n500 585
R60 B.n502 B.n31 585
R61 B.n504 B.n503 585
R62 B.n505 B.n30 585
R63 B.n507 B.n506 585
R64 B.n508 B.n29 585
R65 B.n510 B.n509 585
R66 B.n511 B.n28 585
R67 B.n513 B.n512 585
R68 B.n514 B.n27 585
R69 B.n516 B.n515 585
R70 B.n517 B.n26 585
R71 B.n519 B.n518 585
R72 B.n520 B.n25 585
R73 B.n522 B.n521 585
R74 B.n523 B.n24 585
R75 B.n525 B.n524 585
R76 B.n526 B.n23 585
R77 B.n528 B.n527 585
R78 B.n529 B.n22 585
R79 B.n531 B.n530 585
R80 B.n532 B.n21 585
R81 B.n534 B.n533 585
R82 B.n535 B.n20 585
R83 B.n537 B.n536 585
R84 B.n538 B.n19 585
R85 B.n540 B.n539 585
R86 B.n541 B.n18 585
R87 B.n543 B.n542 585
R88 B.n544 B.n17 585
R89 B.n546 B.n545 585
R90 B.n547 B.n16 585
R91 B.n549 B.n548 585
R92 B.n550 B.n15 585
R93 B.n552 B.n551 585
R94 B.n410 B.n409 585
R95 B.n408 B.n67 585
R96 B.n407 B.n406 585
R97 B.n405 B.n68 585
R98 B.n404 B.n403 585
R99 B.n402 B.n69 585
R100 B.n401 B.n400 585
R101 B.n399 B.n70 585
R102 B.n398 B.n397 585
R103 B.n396 B.n71 585
R104 B.n395 B.n394 585
R105 B.n393 B.n72 585
R106 B.n392 B.n391 585
R107 B.n390 B.n73 585
R108 B.n389 B.n388 585
R109 B.n387 B.n74 585
R110 B.n386 B.n385 585
R111 B.n384 B.n75 585
R112 B.n383 B.n382 585
R113 B.n381 B.n76 585
R114 B.n380 B.n379 585
R115 B.n378 B.n77 585
R116 B.n377 B.n376 585
R117 B.n375 B.n78 585
R118 B.n374 B.n373 585
R119 B.n372 B.n79 585
R120 B.n371 B.n370 585
R121 B.n369 B.n80 585
R122 B.n368 B.n367 585
R123 B.n366 B.n81 585
R124 B.n365 B.n364 585
R125 B.n363 B.n82 585
R126 B.n362 B.n361 585
R127 B.n360 B.n83 585
R128 B.n359 B.n358 585
R129 B.n357 B.n84 585
R130 B.n356 B.n355 585
R131 B.n354 B.n85 585
R132 B.n353 B.n352 585
R133 B.n351 B.n86 585
R134 B.n350 B.n349 585
R135 B.n348 B.n87 585
R136 B.n347 B.n346 585
R137 B.n345 B.n88 585
R138 B.n344 B.n343 585
R139 B.n342 B.n89 585
R140 B.n341 B.n340 585
R141 B.n339 B.n90 585
R142 B.n338 B.n337 585
R143 B.n336 B.n91 585
R144 B.n335 B.n334 585
R145 B.n192 B.n143 585
R146 B.n194 B.n193 585
R147 B.n195 B.n142 585
R148 B.n197 B.n196 585
R149 B.n198 B.n141 585
R150 B.n200 B.n199 585
R151 B.n201 B.n140 585
R152 B.n203 B.n202 585
R153 B.n204 B.n139 585
R154 B.n206 B.n205 585
R155 B.n207 B.n138 585
R156 B.n209 B.n208 585
R157 B.n210 B.n137 585
R158 B.n212 B.n211 585
R159 B.n213 B.n136 585
R160 B.n215 B.n214 585
R161 B.n216 B.n135 585
R162 B.n218 B.n217 585
R163 B.n219 B.n134 585
R164 B.n221 B.n220 585
R165 B.n222 B.n133 585
R166 B.n224 B.n223 585
R167 B.n225 B.n132 585
R168 B.n227 B.n226 585
R169 B.n228 B.n131 585
R170 B.n230 B.n229 585
R171 B.n231 B.n130 585
R172 B.n233 B.n232 585
R173 B.n234 B.n129 585
R174 B.n236 B.n235 585
R175 B.n237 B.n128 585
R176 B.n239 B.n238 585
R177 B.n240 B.n127 585
R178 B.n242 B.n241 585
R179 B.n243 B.n126 585
R180 B.n245 B.n244 585
R181 B.n246 B.n125 585
R182 B.n248 B.n247 585
R183 B.n249 B.n124 585
R184 B.n251 B.n250 585
R185 B.n252 B.n123 585
R186 B.n254 B.n253 585
R187 B.n256 B.n120 585
R188 B.n258 B.n257 585
R189 B.n259 B.n119 585
R190 B.n261 B.n260 585
R191 B.n262 B.n118 585
R192 B.n264 B.n263 585
R193 B.n265 B.n117 585
R194 B.n267 B.n266 585
R195 B.n268 B.n116 585
R196 B.n270 B.n269 585
R197 B.n272 B.n271 585
R198 B.n273 B.n112 585
R199 B.n275 B.n274 585
R200 B.n276 B.n111 585
R201 B.n278 B.n277 585
R202 B.n279 B.n110 585
R203 B.n281 B.n280 585
R204 B.n282 B.n109 585
R205 B.n284 B.n283 585
R206 B.n285 B.n108 585
R207 B.n287 B.n286 585
R208 B.n288 B.n107 585
R209 B.n290 B.n289 585
R210 B.n291 B.n106 585
R211 B.n293 B.n292 585
R212 B.n294 B.n105 585
R213 B.n296 B.n295 585
R214 B.n297 B.n104 585
R215 B.n299 B.n298 585
R216 B.n300 B.n103 585
R217 B.n302 B.n301 585
R218 B.n303 B.n102 585
R219 B.n305 B.n304 585
R220 B.n306 B.n101 585
R221 B.n308 B.n307 585
R222 B.n309 B.n100 585
R223 B.n311 B.n310 585
R224 B.n312 B.n99 585
R225 B.n314 B.n313 585
R226 B.n315 B.n98 585
R227 B.n317 B.n316 585
R228 B.n318 B.n97 585
R229 B.n320 B.n319 585
R230 B.n321 B.n96 585
R231 B.n323 B.n322 585
R232 B.n324 B.n95 585
R233 B.n326 B.n325 585
R234 B.n327 B.n94 585
R235 B.n329 B.n328 585
R236 B.n330 B.n93 585
R237 B.n332 B.n331 585
R238 B.n333 B.n92 585
R239 B.n191 B.n190 585
R240 B.n189 B.n144 585
R241 B.n188 B.n187 585
R242 B.n186 B.n145 585
R243 B.n185 B.n184 585
R244 B.n183 B.n146 585
R245 B.n182 B.n181 585
R246 B.n180 B.n147 585
R247 B.n179 B.n178 585
R248 B.n177 B.n148 585
R249 B.n176 B.n175 585
R250 B.n174 B.n149 585
R251 B.n173 B.n172 585
R252 B.n171 B.n150 585
R253 B.n170 B.n169 585
R254 B.n168 B.n151 585
R255 B.n167 B.n166 585
R256 B.n165 B.n152 585
R257 B.n164 B.n163 585
R258 B.n162 B.n153 585
R259 B.n161 B.n160 585
R260 B.n159 B.n154 585
R261 B.n158 B.n157 585
R262 B.n156 B.n155 585
R263 B.n2 B.n0 585
R264 B.n589 B.n1 585
R265 B.n588 B.n587 585
R266 B.n586 B.n3 585
R267 B.n585 B.n584 585
R268 B.n583 B.n4 585
R269 B.n582 B.n581 585
R270 B.n580 B.n5 585
R271 B.n579 B.n578 585
R272 B.n577 B.n6 585
R273 B.n576 B.n575 585
R274 B.n574 B.n7 585
R275 B.n573 B.n572 585
R276 B.n571 B.n8 585
R277 B.n570 B.n569 585
R278 B.n568 B.n9 585
R279 B.n567 B.n566 585
R280 B.n565 B.n10 585
R281 B.n564 B.n563 585
R282 B.n562 B.n11 585
R283 B.n561 B.n560 585
R284 B.n559 B.n12 585
R285 B.n558 B.n557 585
R286 B.n556 B.n13 585
R287 B.n555 B.n554 585
R288 B.n553 B.n14 585
R289 B.n591 B.n590 585
R290 B.n192 B.n191 492.5
R291 B.n553 B.n552 492.5
R292 B.n335 B.n92 492.5
R293 B.n409 B.n66 492.5
R294 B.n113 B.t2 416.063
R295 B.n44 B.t10 416.063
R296 B.n121 B.t5 416.063
R297 B.n36 B.t7 416.063
R298 B.n113 B.t0 390.224
R299 B.n121 B.t3 390.224
R300 B.n36 B.t6 390.224
R301 B.n44 B.t9 390.224
R302 B.n114 B.t1 378.827
R303 B.n45 B.t11 378.827
R304 B.n122 B.t4 378.827
R305 B.n37 B.t8 378.827
R306 B.n191 B.n144 163.367
R307 B.n187 B.n144 163.367
R308 B.n187 B.n186 163.367
R309 B.n186 B.n185 163.367
R310 B.n185 B.n146 163.367
R311 B.n181 B.n146 163.367
R312 B.n181 B.n180 163.367
R313 B.n180 B.n179 163.367
R314 B.n179 B.n148 163.367
R315 B.n175 B.n148 163.367
R316 B.n175 B.n174 163.367
R317 B.n174 B.n173 163.367
R318 B.n173 B.n150 163.367
R319 B.n169 B.n150 163.367
R320 B.n169 B.n168 163.367
R321 B.n168 B.n167 163.367
R322 B.n167 B.n152 163.367
R323 B.n163 B.n152 163.367
R324 B.n163 B.n162 163.367
R325 B.n162 B.n161 163.367
R326 B.n161 B.n154 163.367
R327 B.n157 B.n154 163.367
R328 B.n157 B.n156 163.367
R329 B.n156 B.n2 163.367
R330 B.n590 B.n2 163.367
R331 B.n590 B.n589 163.367
R332 B.n589 B.n588 163.367
R333 B.n588 B.n3 163.367
R334 B.n584 B.n3 163.367
R335 B.n584 B.n583 163.367
R336 B.n583 B.n582 163.367
R337 B.n582 B.n5 163.367
R338 B.n578 B.n5 163.367
R339 B.n578 B.n577 163.367
R340 B.n577 B.n576 163.367
R341 B.n576 B.n7 163.367
R342 B.n572 B.n7 163.367
R343 B.n572 B.n571 163.367
R344 B.n571 B.n570 163.367
R345 B.n570 B.n9 163.367
R346 B.n566 B.n9 163.367
R347 B.n566 B.n565 163.367
R348 B.n565 B.n564 163.367
R349 B.n564 B.n11 163.367
R350 B.n560 B.n11 163.367
R351 B.n560 B.n559 163.367
R352 B.n559 B.n558 163.367
R353 B.n558 B.n13 163.367
R354 B.n554 B.n13 163.367
R355 B.n554 B.n553 163.367
R356 B.n193 B.n192 163.367
R357 B.n193 B.n142 163.367
R358 B.n197 B.n142 163.367
R359 B.n198 B.n197 163.367
R360 B.n199 B.n198 163.367
R361 B.n199 B.n140 163.367
R362 B.n203 B.n140 163.367
R363 B.n204 B.n203 163.367
R364 B.n205 B.n204 163.367
R365 B.n205 B.n138 163.367
R366 B.n209 B.n138 163.367
R367 B.n210 B.n209 163.367
R368 B.n211 B.n210 163.367
R369 B.n211 B.n136 163.367
R370 B.n215 B.n136 163.367
R371 B.n216 B.n215 163.367
R372 B.n217 B.n216 163.367
R373 B.n217 B.n134 163.367
R374 B.n221 B.n134 163.367
R375 B.n222 B.n221 163.367
R376 B.n223 B.n222 163.367
R377 B.n223 B.n132 163.367
R378 B.n227 B.n132 163.367
R379 B.n228 B.n227 163.367
R380 B.n229 B.n228 163.367
R381 B.n229 B.n130 163.367
R382 B.n233 B.n130 163.367
R383 B.n234 B.n233 163.367
R384 B.n235 B.n234 163.367
R385 B.n235 B.n128 163.367
R386 B.n239 B.n128 163.367
R387 B.n240 B.n239 163.367
R388 B.n241 B.n240 163.367
R389 B.n241 B.n126 163.367
R390 B.n245 B.n126 163.367
R391 B.n246 B.n245 163.367
R392 B.n247 B.n246 163.367
R393 B.n247 B.n124 163.367
R394 B.n251 B.n124 163.367
R395 B.n252 B.n251 163.367
R396 B.n253 B.n252 163.367
R397 B.n253 B.n120 163.367
R398 B.n258 B.n120 163.367
R399 B.n259 B.n258 163.367
R400 B.n260 B.n259 163.367
R401 B.n260 B.n118 163.367
R402 B.n264 B.n118 163.367
R403 B.n265 B.n264 163.367
R404 B.n266 B.n265 163.367
R405 B.n266 B.n116 163.367
R406 B.n270 B.n116 163.367
R407 B.n271 B.n270 163.367
R408 B.n271 B.n112 163.367
R409 B.n275 B.n112 163.367
R410 B.n276 B.n275 163.367
R411 B.n277 B.n276 163.367
R412 B.n277 B.n110 163.367
R413 B.n281 B.n110 163.367
R414 B.n282 B.n281 163.367
R415 B.n283 B.n282 163.367
R416 B.n283 B.n108 163.367
R417 B.n287 B.n108 163.367
R418 B.n288 B.n287 163.367
R419 B.n289 B.n288 163.367
R420 B.n289 B.n106 163.367
R421 B.n293 B.n106 163.367
R422 B.n294 B.n293 163.367
R423 B.n295 B.n294 163.367
R424 B.n295 B.n104 163.367
R425 B.n299 B.n104 163.367
R426 B.n300 B.n299 163.367
R427 B.n301 B.n300 163.367
R428 B.n301 B.n102 163.367
R429 B.n305 B.n102 163.367
R430 B.n306 B.n305 163.367
R431 B.n307 B.n306 163.367
R432 B.n307 B.n100 163.367
R433 B.n311 B.n100 163.367
R434 B.n312 B.n311 163.367
R435 B.n313 B.n312 163.367
R436 B.n313 B.n98 163.367
R437 B.n317 B.n98 163.367
R438 B.n318 B.n317 163.367
R439 B.n319 B.n318 163.367
R440 B.n319 B.n96 163.367
R441 B.n323 B.n96 163.367
R442 B.n324 B.n323 163.367
R443 B.n325 B.n324 163.367
R444 B.n325 B.n94 163.367
R445 B.n329 B.n94 163.367
R446 B.n330 B.n329 163.367
R447 B.n331 B.n330 163.367
R448 B.n331 B.n92 163.367
R449 B.n336 B.n335 163.367
R450 B.n337 B.n336 163.367
R451 B.n337 B.n90 163.367
R452 B.n341 B.n90 163.367
R453 B.n342 B.n341 163.367
R454 B.n343 B.n342 163.367
R455 B.n343 B.n88 163.367
R456 B.n347 B.n88 163.367
R457 B.n348 B.n347 163.367
R458 B.n349 B.n348 163.367
R459 B.n349 B.n86 163.367
R460 B.n353 B.n86 163.367
R461 B.n354 B.n353 163.367
R462 B.n355 B.n354 163.367
R463 B.n355 B.n84 163.367
R464 B.n359 B.n84 163.367
R465 B.n360 B.n359 163.367
R466 B.n361 B.n360 163.367
R467 B.n361 B.n82 163.367
R468 B.n365 B.n82 163.367
R469 B.n366 B.n365 163.367
R470 B.n367 B.n366 163.367
R471 B.n367 B.n80 163.367
R472 B.n371 B.n80 163.367
R473 B.n372 B.n371 163.367
R474 B.n373 B.n372 163.367
R475 B.n373 B.n78 163.367
R476 B.n377 B.n78 163.367
R477 B.n378 B.n377 163.367
R478 B.n379 B.n378 163.367
R479 B.n379 B.n76 163.367
R480 B.n383 B.n76 163.367
R481 B.n384 B.n383 163.367
R482 B.n385 B.n384 163.367
R483 B.n385 B.n74 163.367
R484 B.n389 B.n74 163.367
R485 B.n390 B.n389 163.367
R486 B.n391 B.n390 163.367
R487 B.n391 B.n72 163.367
R488 B.n395 B.n72 163.367
R489 B.n396 B.n395 163.367
R490 B.n397 B.n396 163.367
R491 B.n397 B.n70 163.367
R492 B.n401 B.n70 163.367
R493 B.n402 B.n401 163.367
R494 B.n403 B.n402 163.367
R495 B.n403 B.n68 163.367
R496 B.n407 B.n68 163.367
R497 B.n408 B.n407 163.367
R498 B.n409 B.n408 163.367
R499 B.n552 B.n15 163.367
R500 B.n548 B.n15 163.367
R501 B.n548 B.n547 163.367
R502 B.n547 B.n546 163.367
R503 B.n546 B.n17 163.367
R504 B.n542 B.n17 163.367
R505 B.n542 B.n541 163.367
R506 B.n541 B.n540 163.367
R507 B.n540 B.n19 163.367
R508 B.n536 B.n19 163.367
R509 B.n536 B.n535 163.367
R510 B.n535 B.n534 163.367
R511 B.n534 B.n21 163.367
R512 B.n530 B.n21 163.367
R513 B.n530 B.n529 163.367
R514 B.n529 B.n528 163.367
R515 B.n528 B.n23 163.367
R516 B.n524 B.n23 163.367
R517 B.n524 B.n523 163.367
R518 B.n523 B.n522 163.367
R519 B.n522 B.n25 163.367
R520 B.n518 B.n25 163.367
R521 B.n518 B.n517 163.367
R522 B.n517 B.n516 163.367
R523 B.n516 B.n27 163.367
R524 B.n512 B.n27 163.367
R525 B.n512 B.n511 163.367
R526 B.n511 B.n510 163.367
R527 B.n510 B.n29 163.367
R528 B.n506 B.n29 163.367
R529 B.n506 B.n505 163.367
R530 B.n505 B.n504 163.367
R531 B.n504 B.n31 163.367
R532 B.n500 B.n31 163.367
R533 B.n500 B.n499 163.367
R534 B.n499 B.n498 163.367
R535 B.n498 B.n33 163.367
R536 B.n494 B.n33 163.367
R537 B.n494 B.n493 163.367
R538 B.n493 B.n492 163.367
R539 B.n492 B.n35 163.367
R540 B.n487 B.n35 163.367
R541 B.n487 B.n486 163.367
R542 B.n486 B.n485 163.367
R543 B.n485 B.n39 163.367
R544 B.n481 B.n39 163.367
R545 B.n481 B.n480 163.367
R546 B.n480 B.n479 163.367
R547 B.n479 B.n41 163.367
R548 B.n475 B.n41 163.367
R549 B.n475 B.n474 163.367
R550 B.n474 B.n473 163.367
R551 B.n473 B.n43 163.367
R552 B.n469 B.n43 163.367
R553 B.n469 B.n468 163.367
R554 B.n468 B.n467 163.367
R555 B.n467 B.n48 163.367
R556 B.n463 B.n48 163.367
R557 B.n463 B.n462 163.367
R558 B.n462 B.n461 163.367
R559 B.n461 B.n50 163.367
R560 B.n457 B.n50 163.367
R561 B.n457 B.n456 163.367
R562 B.n456 B.n455 163.367
R563 B.n455 B.n52 163.367
R564 B.n451 B.n52 163.367
R565 B.n451 B.n450 163.367
R566 B.n450 B.n449 163.367
R567 B.n449 B.n54 163.367
R568 B.n445 B.n54 163.367
R569 B.n445 B.n444 163.367
R570 B.n444 B.n443 163.367
R571 B.n443 B.n56 163.367
R572 B.n439 B.n56 163.367
R573 B.n439 B.n438 163.367
R574 B.n438 B.n437 163.367
R575 B.n437 B.n58 163.367
R576 B.n433 B.n58 163.367
R577 B.n433 B.n432 163.367
R578 B.n432 B.n431 163.367
R579 B.n431 B.n60 163.367
R580 B.n427 B.n60 163.367
R581 B.n427 B.n426 163.367
R582 B.n426 B.n425 163.367
R583 B.n425 B.n62 163.367
R584 B.n421 B.n62 163.367
R585 B.n421 B.n420 163.367
R586 B.n420 B.n419 163.367
R587 B.n419 B.n64 163.367
R588 B.n415 B.n64 163.367
R589 B.n415 B.n414 163.367
R590 B.n414 B.n413 163.367
R591 B.n413 B.n66 163.367
R592 B.n115 B.n114 59.5399
R593 B.n255 B.n122 59.5399
R594 B.n489 B.n37 59.5399
R595 B.n46 B.n45 59.5399
R596 B.n114 B.n113 37.2369
R597 B.n122 B.n121 37.2369
R598 B.n37 B.n36 37.2369
R599 B.n45 B.n44 37.2369
R600 B.n551 B.n14 32.0005
R601 B.n411 B.n410 32.0005
R602 B.n334 B.n333 32.0005
R603 B.n190 B.n143 32.0005
R604 B B.n591 18.0485
R605 B.n551 B.n550 10.6151
R606 B.n550 B.n549 10.6151
R607 B.n549 B.n16 10.6151
R608 B.n545 B.n16 10.6151
R609 B.n545 B.n544 10.6151
R610 B.n544 B.n543 10.6151
R611 B.n543 B.n18 10.6151
R612 B.n539 B.n18 10.6151
R613 B.n539 B.n538 10.6151
R614 B.n538 B.n537 10.6151
R615 B.n537 B.n20 10.6151
R616 B.n533 B.n20 10.6151
R617 B.n533 B.n532 10.6151
R618 B.n532 B.n531 10.6151
R619 B.n531 B.n22 10.6151
R620 B.n527 B.n22 10.6151
R621 B.n527 B.n526 10.6151
R622 B.n526 B.n525 10.6151
R623 B.n525 B.n24 10.6151
R624 B.n521 B.n24 10.6151
R625 B.n521 B.n520 10.6151
R626 B.n520 B.n519 10.6151
R627 B.n519 B.n26 10.6151
R628 B.n515 B.n26 10.6151
R629 B.n515 B.n514 10.6151
R630 B.n514 B.n513 10.6151
R631 B.n513 B.n28 10.6151
R632 B.n509 B.n28 10.6151
R633 B.n509 B.n508 10.6151
R634 B.n508 B.n507 10.6151
R635 B.n507 B.n30 10.6151
R636 B.n503 B.n30 10.6151
R637 B.n503 B.n502 10.6151
R638 B.n502 B.n501 10.6151
R639 B.n501 B.n32 10.6151
R640 B.n497 B.n32 10.6151
R641 B.n497 B.n496 10.6151
R642 B.n496 B.n495 10.6151
R643 B.n495 B.n34 10.6151
R644 B.n491 B.n34 10.6151
R645 B.n491 B.n490 10.6151
R646 B.n488 B.n38 10.6151
R647 B.n484 B.n38 10.6151
R648 B.n484 B.n483 10.6151
R649 B.n483 B.n482 10.6151
R650 B.n482 B.n40 10.6151
R651 B.n478 B.n40 10.6151
R652 B.n478 B.n477 10.6151
R653 B.n477 B.n476 10.6151
R654 B.n476 B.n42 10.6151
R655 B.n472 B.n471 10.6151
R656 B.n471 B.n470 10.6151
R657 B.n470 B.n47 10.6151
R658 B.n466 B.n47 10.6151
R659 B.n466 B.n465 10.6151
R660 B.n465 B.n464 10.6151
R661 B.n464 B.n49 10.6151
R662 B.n460 B.n49 10.6151
R663 B.n460 B.n459 10.6151
R664 B.n459 B.n458 10.6151
R665 B.n458 B.n51 10.6151
R666 B.n454 B.n51 10.6151
R667 B.n454 B.n453 10.6151
R668 B.n453 B.n452 10.6151
R669 B.n452 B.n53 10.6151
R670 B.n448 B.n53 10.6151
R671 B.n448 B.n447 10.6151
R672 B.n447 B.n446 10.6151
R673 B.n446 B.n55 10.6151
R674 B.n442 B.n55 10.6151
R675 B.n442 B.n441 10.6151
R676 B.n441 B.n440 10.6151
R677 B.n440 B.n57 10.6151
R678 B.n436 B.n57 10.6151
R679 B.n436 B.n435 10.6151
R680 B.n435 B.n434 10.6151
R681 B.n434 B.n59 10.6151
R682 B.n430 B.n59 10.6151
R683 B.n430 B.n429 10.6151
R684 B.n429 B.n428 10.6151
R685 B.n428 B.n61 10.6151
R686 B.n424 B.n61 10.6151
R687 B.n424 B.n423 10.6151
R688 B.n423 B.n422 10.6151
R689 B.n422 B.n63 10.6151
R690 B.n418 B.n63 10.6151
R691 B.n418 B.n417 10.6151
R692 B.n417 B.n416 10.6151
R693 B.n416 B.n65 10.6151
R694 B.n412 B.n65 10.6151
R695 B.n412 B.n411 10.6151
R696 B.n334 B.n91 10.6151
R697 B.n338 B.n91 10.6151
R698 B.n339 B.n338 10.6151
R699 B.n340 B.n339 10.6151
R700 B.n340 B.n89 10.6151
R701 B.n344 B.n89 10.6151
R702 B.n345 B.n344 10.6151
R703 B.n346 B.n345 10.6151
R704 B.n346 B.n87 10.6151
R705 B.n350 B.n87 10.6151
R706 B.n351 B.n350 10.6151
R707 B.n352 B.n351 10.6151
R708 B.n352 B.n85 10.6151
R709 B.n356 B.n85 10.6151
R710 B.n357 B.n356 10.6151
R711 B.n358 B.n357 10.6151
R712 B.n358 B.n83 10.6151
R713 B.n362 B.n83 10.6151
R714 B.n363 B.n362 10.6151
R715 B.n364 B.n363 10.6151
R716 B.n364 B.n81 10.6151
R717 B.n368 B.n81 10.6151
R718 B.n369 B.n368 10.6151
R719 B.n370 B.n369 10.6151
R720 B.n370 B.n79 10.6151
R721 B.n374 B.n79 10.6151
R722 B.n375 B.n374 10.6151
R723 B.n376 B.n375 10.6151
R724 B.n376 B.n77 10.6151
R725 B.n380 B.n77 10.6151
R726 B.n381 B.n380 10.6151
R727 B.n382 B.n381 10.6151
R728 B.n382 B.n75 10.6151
R729 B.n386 B.n75 10.6151
R730 B.n387 B.n386 10.6151
R731 B.n388 B.n387 10.6151
R732 B.n388 B.n73 10.6151
R733 B.n392 B.n73 10.6151
R734 B.n393 B.n392 10.6151
R735 B.n394 B.n393 10.6151
R736 B.n394 B.n71 10.6151
R737 B.n398 B.n71 10.6151
R738 B.n399 B.n398 10.6151
R739 B.n400 B.n399 10.6151
R740 B.n400 B.n69 10.6151
R741 B.n404 B.n69 10.6151
R742 B.n405 B.n404 10.6151
R743 B.n406 B.n405 10.6151
R744 B.n406 B.n67 10.6151
R745 B.n410 B.n67 10.6151
R746 B.n194 B.n143 10.6151
R747 B.n195 B.n194 10.6151
R748 B.n196 B.n195 10.6151
R749 B.n196 B.n141 10.6151
R750 B.n200 B.n141 10.6151
R751 B.n201 B.n200 10.6151
R752 B.n202 B.n201 10.6151
R753 B.n202 B.n139 10.6151
R754 B.n206 B.n139 10.6151
R755 B.n207 B.n206 10.6151
R756 B.n208 B.n207 10.6151
R757 B.n208 B.n137 10.6151
R758 B.n212 B.n137 10.6151
R759 B.n213 B.n212 10.6151
R760 B.n214 B.n213 10.6151
R761 B.n214 B.n135 10.6151
R762 B.n218 B.n135 10.6151
R763 B.n219 B.n218 10.6151
R764 B.n220 B.n219 10.6151
R765 B.n220 B.n133 10.6151
R766 B.n224 B.n133 10.6151
R767 B.n225 B.n224 10.6151
R768 B.n226 B.n225 10.6151
R769 B.n226 B.n131 10.6151
R770 B.n230 B.n131 10.6151
R771 B.n231 B.n230 10.6151
R772 B.n232 B.n231 10.6151
R773 B.n232 B.n129 10.6151
R774 B.n236 B.n129 10.6151
R775 B.n237 B.n236 10.6151
R776 B.n238 B.n237 10.6151
R777 B.n238 B.n127 10.6151
R778 B.n242 B.n127 10.6151
R779 B.n243 B.n242 10.6151
R780 B.n244 B.n243 10.6151
R781 B.n244 B.n125 10.6151
R782 B.n248 B.n125 10.6151
R783 B.n249 B.n248 10.6151
R784 B.n250 B.n249 10.6151
R785 B.n250 B.n123 10.6151
R786 B.n254 B.n123 10.6151
R787 B.n257 B.n256 10.6151
R788 B.n257 B.n119 10.6151
R789 B.n261 B.n119 10.6151
R790 B.n262 B.n261 10.6151
R791 B.n263 B.n262 10.6151
R792 B.n263 B.n117 10.6151
R793 B.n267 B.n117 10.6151
R794 B.n268 B.n267 10.6151
R795 B.n269 B.n268 10.6151
R796 B.n273 B.n272 10.6151
R797 B.n274 B.n273 10.6151
R798 B.n274 B.n111 10.6151
R799 B.n278 B.n111 10.6151
R800 B.n279 B.n278 10.6151
R801 B.n280 B.n279 10.6151
R802 B.n280 B.n109 10.6151
R803 B.n284 B.n109 10.6151
R804 B.n285 B.n284 10.6151
R805 B.n286 B.n285 10.6151
R806 B.n286 B.n107 10.6151
R807 B.n290 B.n107 10.6151
R808 B.n291 B.n290 10.6151
R809 B.n292 B.n291 10.6151
R810 B.n292 B.n105 10.6151
R811 B.n296 B.n105 10.6151
R812 B.n297 B.n296 10.6151
R813 B.n298 B.n297 10.6151
R814 B.n298 B.n103 10.6151
R815 B.n302 B.n103 10.6151
R816 B.n303 B.n302 10.6151
R817 B.n304 B.n303 10.6151
R818 B.n304 B.n101 10.6151
R819 B.n308 B.n101 10.6151
R820 B.n309 B.n308 10.6151
R821 B.n310 B.n309 10.6151
R822 B.n310 B.n99 10.6151
R823 B.n314 B.n99 10.6151
R824 B.n315 B.n314 10.6151
R825 B.n316 B.n315 10.6151
R826 B.n316 B.n97 10.6151
R827 B.n320 B.n97 10.6151
R828 B.n321 B.n320 10.6151
R829 B.n322 B.n321 10.6151
R830 B.n322 B.n95 10.6151
R831 B.n326 B.n95 10.6151
R832 B.n327 B.n326 10.6151
R833 B.n328 B.n327 10.6151
R834 B.n328 B.n93 10.6151
R835 B.n332 B.n93 10.6151
R836 B.n333 B.n332 10.6151
R837 B.n190 B.n189 10.6151
R838 B.n189 B.n188 10.6151
R839 B.n188 B.n145 10.6151
R840 B.n184 B.n145 10.6151
R841 B.n184 B.n183 10.6151
R842 B.n183 B.n182 10.6151
R843 B.n182 B.n147 10.6151
R844 B.n178 B.n147 10.6151
R845 B.n178 B.n177 10.6151
R846 B.n177 B.n176 10.6151
R847 B.n176 B.n149 10.6151
R848 B.n172 B.n149 10.6151
R849 B.n172 B.n171 10.6151
R850 B.n171 B.n170 10.6151
R851 B.n170 B.n151 10.6151
R852 B.n166 B.n151 10.6151
R853 B.n166 B.n165 10.6151
R854 B.n165 B.n164 10.6151
R855 B.n164 B.n153 10.6151
R856 B.n160 B.n153 10.6151
R857 B.n160 B.n159 10.6151
R858 B.n159 B.n158 10.6151
R859 B.n158 B.n155 10.6151
R860 B.n155 B.n0 10.6151
R861 B.n587 B.n1 10.6151
R862 B.n587 B.n586 10.6151
R863 B.n586 B.n585 10.6151
R864 B.n585 B.n4 10.6151
R865 B.n581 B.n4 10.6151
R866 B.n581 B.n580 10.6151
R867 B.n580 B.n579 10.6151
R868 B.n579 B.n6 10.6151
R869 B.n575 B.n6 10.6151
R870 B.n575 B.n574 10.6151
R871 B.n574 B.n573 10.6151
R872 B.n573 B.n8 10.6151
R873 B.n569 B.n8 10.6151
R874 B.n569 B.n568 10.6151
R875 B.n568 B.n567 10.6151
R876 B.n567 B.n10 10.6151
R877 B.n563 B.n10 10.6151
R878 B.n563 B.n562 10.6151
R879 B.n562 B.n561 10.6151
R880 B.n561 B.n12 10.6151
R881 B.n557 B.n12 10.6151
R882 B.n557 B.n556 10.6151
R883 B.n556 B.n555 10.6151
R884 B.n555 B.n14 10.6151
R885 B.n490 B.n489 9.36635
R886 B.n472 B.n46 9.36635
R887 B.n255 B.n254 9.36635
R888 B.n272 B.n115 9.36635
R889 B.n591 B.n0 2.81026
R890 B.n591 B.n1 2.81026
R891 B.n489 B.n488 1.24928
R892 B.n46 B.n42 1.24928
R893 B.n256 B.n255 1.24928
R894 B.n269 B.n115 1.24928
R895 VP.n2 VP.t3 222.115
R896 VP.n2 VP.t2 221.791
R897 VP.n4 VP.t0 184.464
R898 VP.n11 VP.t1 184.464
R899 VP.n4 VP.n3 175.492
R900 VP.n12 VP.n11 175.492
R901 VP.n10 VP.n0 161.3
R902 VP.n9 VP.n8 161.3
R903 VP.n7 VP.n1 161.3
R904 VP.n6 VP.n5 161.3
R905 VP.n9 VP.n1 56.5193
R906 VP.n3 VP.n2 56.0376
R907 VP.n5 VP.n1 24.4675
R908 VP.n10 VP.n9 24.4675
R909 VP.n5 VP.n4 10.2766
R910 VP.n11 VP.n10 10.2766
R911 VP.n6 VP.n3 0.189894
R912 VP.n7 VP.n6 0.189894
R913 VP.n8 VP.n7 0.189894
R914 VP.n8 VP.n0 0.189894
R915 VP.n12 VP.n0 0.189894
R916 VP VP.n12 0.0516364
R917 VDD1 VDD1.n1 114.505
R918 VDD1 VDD1.n0 74.8669
R919 VDD1.n0 VDD1.t3 2.67141
R920 VDD1.n0 VDD1.t2 2.67141
R921 VDD1.n1 VDD1.t0 2.67141
R922 VDD1.n1 VDD1.t1 2.67141
R923 VTAIL.n522 VTAIL.n462 756.745
R924 VTAIL.n60 VTAIL.n0 756.745
R925 VTAIL.n126 VTAIL.n66 756.745
R926 VTAIL.n192 VTAIL.n132 756.745
R927 VTAIL.n456 VTAIL.n396 756.745
R928 VTAIL.n390 VTAIL.n330 756.745
R929 VTAIL.n324 VTAIL.n264 756.745
R930 VTAIL.n258 VTAIL.n198 756.745
R931 VTAIL.n482 VTAIL.n481 585
R932 VTAIL.n487 VTAIL.n486 585
R933 VTAIL.n489 VTAIL.n488 585
R934 VTAIL.n478 VTAIL.n477 585
R935 VTAIL.n495 VTAIL.n494 585
R936 VTAIL.n497 VTAIL.n496 585
R937 VTAIL.n474 VTAIL.n473 585
R938 VTAIL.n504 VTAIL.n503 585
R939 VTAIL.n505 VTAIL.n472 585
R940 VTAIL.n507 VTAIL.n506 585
R941 VTAIL.n470 VTAIL.n469 585
R942 VTAIL.n513 VTAIL.n512 585
R943 VTAIL.n515 VTAIL.n514 585
R944 VTAIL.n466 VTAIL.n465 585
R945 VTAIL.n521 VTAIL.n520 585
R946 VTAIL.n523 VTAIL.n522 585
R947 VTAIL.n20 VTAIL.n19 585
R948 VTAIL.n25 VTAIL.n24 585
R949 VTAIL.n27 VTAIL.n26 585
R950 VTAIL.n16 VTAIL.n15 585
R951 VTAIL.n33 VTAIL.n32 585
R952 VTAIL.n35 VTAIL.n34 585
R953 VTAIL.n12 VTAIL.n11 585
R954 VTAIL.n42 VTAIL.n41 585
R955 VTAIL.n43 VTAIL.n10 585
R956 VTAIL.n45 VTAIL.n44 585
R957 VTAIL.n8 VTAIL.n7 585
R958 VTAIL.n51 VTAIL.n50 585
R959 VTAIL.n53 VTAIL.n52 585
R960 VTAIL.n4 VTAIL.n3 585
R961 VTAIL.n59 VTAIL.n58 585
R962 VTAIL.n61 VTAIL.n60 585
R963 VTAIL.n86 VTAIL.n85 585
R964 VTAIL.n91 VTAIL.n90 585
R965 VTAIL.n93 VTAIL.n92 585
R966 VTAIL.n82 VTAIL.n81 585
R967 VTAIL.n99 VTAIL.n98 585
R968 VTAIL.n101 VTAIL.n100 585
R969 VTAIL.n78 VTAIL.n77 585
R970 VTAIL.n108 VTAIL.n107 585
R971 VTAIL.n109 VTAIL.n76 585
R972 VTAIL.n111 VTAIL.n110 585
R973 VTAIL.n74 VTAIL.n73 585
R974 VTAIL.n117 VTAIL.n116 585
R975 VTAIL.n119 VTAIL.n118 585
R976 VTAIL.n70 VTAIL.n69 585
R977 VTAIL.n125 VTAIL.n124 585
R978 VTAIL.n127 VTAIL.n126 585
R979 VTAIL.n152 VTAIL.n151 585
R980 VTAIL.n157 VTAIL.n156 585
R981 VTAIL.n159 VTAIL.n158 585
R982 VTAIL.n148 VTAIL.n147 585
R983 VTAIL.n165 VTAIL.n164 585
R984 VTAIL.n167 VTAIL.n166 585
R985 VTAIL.n144 VTAIL.n143 585
R986 VTAIL.n174 VTAIL.n173 585
R987 VTAIL.n175 VTAIL.n142 585
R988 VTAIL.n177 VTAIL.n176 585
R989 VTAIL.n140 VTAIL.n139 585
R990 VTAIL.n183 VTAIL.n182 585
R991 VTAIL.n185 VTAIL.n184 585
R992 VTAIL.n136 VTAIL.n135 585
R993 VTAIL.n191 VTAIL.n190 585
R994 VTAIL.n193 VTAIL.n192 585
R995 VTAIL.n457 VTAIL.n456 585
R996 VTAIL.n455 VTAIL.n454 585
R997 VTAIL.n400 VTAIL.n399 585
R998 VTAIL.n449 VTAIL.n448 585
R999 VTAIL.n447 VTAIL.n446 585
R1000 VTAIL.n404 VTAIL.n403 585
R1001 VTAIL.n441 VTAIL.n440 585
R1002 VTAIL.n439 VTAIL.n406 585
R1003 VTAIL.n438 VTAIL.n437 585
R1004 VTAIL.n409 VTAIL.n407 585
R1005 VTAIL.n432 VTAIL.n431 585
R1006 VTAIL.n430 VTAIL.n429 585
R1007 VTAIL.n413 VTAIL.n412 585
R1008 VTAIL.n424 VTAIL.n423 585
R1009 VTAIL.n422 VTAIL.n421 585
R1010 VTAIL.n417 VTAIL.n416 585
R1011 VTAIL.n391 VTAIL.n390 585
R1012 VTAIL.n389 VTAIL.n388 585
R1013 VTAIL.n334 VTAIL.n333 585
R1014 VTAIL.n383 VTAIL.n382 585
R1015 VTAIL.n381 VTAIL.n380 585
R1016 VTAIL.n338 VTAIL.n337 585
R1017 VTAIL.n375 VTAIL.n374 585
R1018 VTAIL.n373 VTAIL.n340 585
R1019 VTAIL.n372 VTAIL.n371 585
R1020 VTAIL.n343 VTAIL.n341 585
R1021 VTAIL.n366 VTAIL.n365 585
R1022 VTAIL.n364 VTAIL.n363 585
R1023 VTAIL.n347 VTAIL.n346 585
R1024 VTAIL.n358 VTAIL.n357 585
R1025 VTAIL.n356 VTAIL.n355 585
R1026 VTAIL.n351 VTAIL.n350 585
R1027 VTAIL.n325 VTAIL.n324 585
R1028 VTAIL.n323 VTAIL.n322 585
R1029 VTAIL.n268 VTAIL.n267 585
R1030 VTAIL.n317 VTAIL.n316 585
R1031 VTAIL.n315 VTAIL.n314 585
R1032 VTAIL.n272 VTAIL.n271 585
R1033 VTAIL.n309 VTAIL.n308 585
R1034 VTAIL.n307 VTAIL.n274 585
R1035 VTAIL.n306 VTAIL.n305 585
R1036 VTAIL.n277 VTAIL.n275 585
R1037 VTAIL.n300 VTAIL.n299 585
R1038 VTAIL.n298 VTAIL.n297 585
R1039 VTAIL.n281 VTAIL.n280 585
R1040 VTAIL.n292 VTAIL.n291 585
R1041 VTAIL.n290 VTAIL.n289 585
R1042 VTAIL.n285 VTAIL.n284 585
R1043 VTAIL.n259 VTAIL.n258 585
R1044 VTAIL.n257 VTAIL.n256 585
R1045 VTAIL.n202 VTAIL.n201 585
R1046 VTAIL.n251 VTAIL.n250 585
R1047 VTAIL.n249 VTAIL.n248 585
R1048 VTAIL.n206 VTAIL.n205 585
R1049 VTAIL.n243 VTAIL.n242 585
R1050 VTAIL.n241 VTAIL.n208 585
R1051 VTAIL.n240 VTAIL.n239 585
R1052 VTAIL.n211 VTAIL.n209 585
R1053 VTAIL.n234 VTAIL.n233 585
R1054 VTAIL.n232 VTAIL.n231 585
R1055 VTAIL.n215 VTAIL.n214 585
R1056 VTAIL.n226 VTAIL.n225 585
R1057 VTAIL.n224 VTAIL.n223 585
R1058 VTAIL.n219 VTAIL.n218 585
R1059 VTAIL.n483 VTAIL.t2 329.036
R1060 VTAIL.n21 VTAIL.t3 329.036
R1061 VTAIL.n87 VTAIL.t6 329.036
R1062 VTAIL.n153 VTAIL.t7 329.036
R1063 VTAIL.n418 VTAIL.t5 329.036
R1064 VTAIL.n352 VTAIL.t4 329.036
R1065 VTAIL.n286 VTAIL.t1 329.036
R1066 VTAIL.n220 VTAIL.t0 329.036
R1067 VTAIL.n487 VTAIL.n481 171.744
R1068 VTAIL.n488 VTAIL.n487 171.744
R1069 VTAIL.n488 VTAIL.n477 171.744
R1070 VTAIL.n495 VTAIL.n477 171.744
R1071 VTAIL.n496 VTAIL.n495 171.744
R1072 VTAIL.n496 VTAIL.n473 171.744
R1073 VTAIL.n504 VTAIL.n473 171.744
R1074 VTAIL.n505 VTAIL.n504 171.744
R1075 VTAIL.n506 VTAIL.n505 171.744
R1076 VTAIL.n506 VTAIL.n469 171.744
R1077 VTAIL.n513 VTAIL.n469 171.744
R1078 VTAIL.n514 VTAIL.n513 171.744
R1079 VTAIL.n514 VTAIL.n465 171.744
R1080 VTAIL.n521 VTAIL.n465 171.744
R1081 VTAIL.n522 VTAIL.n521 171.744
R1082 VTAIL.n25 VTAIL.n19 171.744
R1083 VTAIL.n26 VTAIL.n25 171.744
R1084 VTAIL.n26 VTAIL.n15 171.744
R1085 VTAIL.n33 VTAIL.n15 171.744
R1086 VTAIL.n34 VTAIL.n33 171.744
R1087 VTAIL.n34 VTAIL.n11 171.744
R1088 VTAIL.n42 VTAIL.n11 171.744
R1089 VTAIL.n43 VTAIL.n42 171.744
R1090 VTAIL.n44 VTAIL.n43 171.744
R1091 VTAIL.n44 VTAIL.n7 171.744
R1092 VTAIL.n51 VTAIL.n7 171.744
R1093 VTAIL.n52 VTAIL.n51 171.744
R1094 VTAIL.n52 VTAIL.n3 171.744
R1095 VTAIL.n59 VTAIL.n3 171.744
R1096 VTAIL.n60 VTAIL.n59 171.744
R1097 VTAIL.n91 VTAIL.n85 171.744
R1098 VTAIL.n92 VTAIL.n91 171.744
R1099 VTAIL.n92 VTAIL.n81 171.744
R1100 VTAIL.n99 VTAIL.n81 171.744
R1101 VTAIL.n100 VTAIL.n99 171.744
R1102 VTAIL.n100 VTAIL.n77 171.744
R1103 VTAIL.n108 VTAIL.n77 171.744
R1104 VTAIL.n109 VTAIL.n108 171.744
R1105 VTAIL.n110 VTAIL.n109 171.744
R1106 VTAIL.n110 VTAIL.n73 171.744
R1107 VTAIL.n117 VTAIL.n73 171.744
R1108 VTAIL.n118 VTAIL.n117 171.744
R1109 VTAIL.n118 VTAIL.n69 171.744
R1110 VTAIL.n125 VTAIL.n69 171.744
R1111 VTAIL.n126 VTAIL.n125 171.744
R1112 VTAIL.n157 VTAIL.n151 171.744
R1113 VTAIL.n158 VTAIL.n157 171.744
R1114 VTAIL.n158 VTAIL.n147 171.744
R1115 VTAIL.n165 VTAIL.n147 171.744
R1116 VTAIL.n166 VTAIL.n165 171.744
R1117 VTAIL.n166 VTAIL.n143 171.744
R1118 VTAIL.n174 VTAIL.n143 171.744
R1119 VTAIL.n175 VTAIL.n174 171.744
R1120 VTAIL.n176 VTAIL.n175 171.744
R1121 VTAIL.n176 VTAIL.n139 171.744
R1122 VTAIL.n183 VTAIL.n139 171.744
R1123 VTAIL.n184 VTAIL.n183 171.744
R1124 VTAIL.n184 VTAIL.n135 171.744
R1125 VTAIL.n191 VTAIL.n135 171.744
R1126 VTAIL.n192 VTAIL.n191 171.744
R1127 VTAIL.n456 VTAIL.n455 171.744
R1128 VTAIL.n455 VTAIL.n399 171.744
R1129 VTAIL.n448 VTAIL.n399 171.744
R1130 VTAIL.n448 VTAIL.n447 171.744
R1131 VTAIL.n447 VTAIL.n403 171.744
R1132 VTAIL.n440 VTAIL.n403 171.744
R1133 VTAIL.n440 VTAIL.n439 171.744
R1134 VTAIL.n439 VTAIL.n438 171.744
R1135 VTAIL.n438 VTAIL.n407 171.744
R1136 VTAIL.n431 VTAIL.n407 171.744
R1137 VTAIL.n431 VTAIL.n430 171.744
R1138 VTAIL.n430 VTAIL.n412 171.744
R1139 VTAIL.n423 VTAIL.n412 171.744
R1140 VTAIL.n423 VTAIL.n422 171.744
R1141 VTAIL.n422 VTAIL.n416 171.744
R1142 VTAIL.n390 VTAIL.n389 171.744
R1143 VTAIL.n389 VTAIL.n333 171.744
R1144 VTAIL.n382 VTAIL.n333 171.744
R1145 VTAIL.n382 VTAIL.n381 171.744
R1146 VTAIL.n381 VTAIL.n337 171.744
R1147 VTAIL.n374 VTAIL.n337 171.744
R1148 VTAIL.n374 VTAIL.n373 171.744
R1149 VTAIL.n373 VTAIL.n372 171.744
R1150 VTAIL.n372 VTAIL.n341 171.744
R1151 VTAIL.n365 VTAIL.n341 171.744
R1152 VTAIL.n365 VTAIL.n364 171.744
R1153 VTAIL.n364 VTAIL.n346 171.744
R1154 VTAIL.n357 VTAIL.n346 171.744
R1155 VTAIL.n357 VTAIL.n356 171.744
R1156 VTAIL.n356 VTAIL.n350 171.744
R1157 VTAIL.n324 VTAIL.n323 171.744
R1158 VTAIL.n323 VTAIL.n267 171.744
R1159 VTAIL.n316 VTAIL.n267 171.744
R1160 VTAIL.n316 VTAIL.n315 171.744
R1161 VTAIL.n315 VTAIL.n271 171.744
R1162 VTAIL.n308 VTAIL.n271 171.744
R1163 VTAIL.n308 VTAIL.n307 171.744
R1164 VTAIL.n307 VTAIL.n306 171.744
R1165 VTAIL.n306 VTAIL.n275 171.744
R1166 VTAIL.n299 VTAIL.n275 171.744
R1167 VTAIL.n299 VTAIL.n298 171.744
R1168 VTAIL.n298 VTAIL.n280 171.744
R1169 VTAIL.n291 VTAIL.n280 171.744
R1170 VTAIL.n291 VTAIL.n290 171.744
R1171 VTAIL.n290 VTAIL.n284 171.744
R1172 VTAIL.n258 VTAIL.n257 171.744
R1173 VTAIL.n257 VTAIL.n201 171.744
R1174 VTAIL.n250 VTAIL.n201 171.744
R1175 VTAIL.n250 VTAIL.n249 171.744
R1176 VTAIL.n249 VTAIL.n205 171.744
R1177 VTAIL.n242 VTAIL.n205 171.744
R1178 VTAIL.n242 VTAIL.n241 171.744
R1179 VTAIL.n241 VTAIL.n240 171.744
R1180 VTAIL.n240 VTAIL.n209 171.744
R1181 VTAIL.n233 VTAIL.n209 171.744
R1182 VTAIL.n233 VTAIL.n232 171.744
R1183 VTAIL.n232 VTAIL.n214 171.744
R1184 VTAIL.n225 VTAIL.n214 171.744
R1185 VTAIL.n225 VTAIL.n224 171.744
R1186 VTAIL.n224 VTAIL.n218 171.744
R1187 VTAIL.t2 VTAIL.n481 85.8723
R1188 VTAIL.t3 VTAIL.n19 85.8723
R1189 VTAIL.t6 VTAIL.n85 85.8723
R1190 VTAIL.t7 VTAIL.n151 85.8723
R1191 VTAIL.t5 VTAIL.n416 85.8723
R1192 VTAIL.t4 VTAIL.n350 85.8723
R1193 VTAIL.t1 VTAIL.n284 85.8723
R1194 VTAIL.t0 VTAIL.n218 85.8723
R1195 VTAIL.n527 VTAIL.n526 33.155
R1196 VTAIL.n65 VTAIL.n64 33.155
R1197 VTAIL.n131 VTAIL.n130 33.155
R1198 VTAIL.n197 VTAIL.n196 33.155
R1199 VTAIL.n461 VTAIL.n460 33.155
R1200 VTAIL.n395 VTAIL.n394 33.155
R1201 VTAIL.n329 VTAIL.n328 33.155
R1202 VTAIL.n263 VTAIL.n262 33.155
R1203 VTAIL.n527 VTAIL.n461 24.5134
R1204 VTAIL.n263 VTAIL.n197 24.5134
R1205 VTAIL.n507 VTAIL.n472 13.1884
R1206 VTAIL.n45 VTAIL.n10 13.1884
R1207 VTAIL.n111 VTAIL.n76 13.1884
R1208 VTAIL.n177 VTAIL.n142 13.1884
R1209 VTAIL.n441 VTAIL.n406 13.1884
R1210 VTAIL.n375 VTAIL.n340 13.1884
R1211 VTAIL.n309 VTAIL.n274 13.1884
R1212 VTAIL.n243 VTAIL.n208 13.1884
R1213 VTAIL.n503 VTAIL.n502 12.8005
R1214 VTAIL.n508 VTAIL.n470 12.8005
R1215 VTAIL.n41 VTAIL.n40 12.8005
R1216 VTAIL.n46 VTAIL.n8 12.8005
R1217 VTAIL.n107 VTAIL.n106 12.8005
R1218 VTAIL.n112 VTAIL.n74 12.8005
R1219 VTAIL.n173 VTAIL.n172 12.8005
R1220 VTAIL.n178 VTAIL.n140 12.8005
R1221 VTAIL.n442 VTAIL.n404 12.8005
R1222 VTAIL.n437 VTAIL.n408 12.8005
R1223 VTAIL.n376 VTAIL.n338 12.8005
R1224 VTAIL.n371 VTAIL.n342 12.8005
R1225 VTAIL.n310 VTAIL.n272 12.8005
R1226 VTAIL.n305 VTAIL.n276 12.8005
R1227 VTAIL.n244 VTAIL.n206 12.8005
R1228 VTAIL.n239 VTAIL.n210 12.8005
R1229 VTAIL.n501 VTAIL.n474 12.0247
R1230 VTAIL.n512 VTAIL.n511 12.0247
R1231 VTAIL.n39 VTAIL.n12 12.0247
R1232 VTAIL.n50 VTAIL.n49 12.0247
R1233 VTAIL.n105 VTAIL.n78 12.0247
R1234 VTAIL.n116 VTAIL.n115 12.0247
R1235 VTAIL.n171 VTAIL.n144 12.0247
R1236 VTAIL.n182 VTAIL.n181 12.0247
R1237 VTAIL.n446 VTAIL.n445 12.0247
R1238 VTAIL.n436 VTAIL.n409 12.0247
R1239 VTAIL.n380 VTAIL.n379 12.0247
R1240 VTAIL.n370 VTAIL.n343 12.0247
R1241 VTAIL.n314 VTAIL.n313 12.0247
R1242 VTAIL.n304 VTAIL.n277 12.0247
R1243 VTAIL.n248 VTAIL.n247 12.0247
R1244 VTAIL.n238 VTAIL.n211 12.0247
R1245 VTAIL.n498 VTAIL.n497 11.249
R1246 VTAIL.n515 VTAIL.n468 11.249
R1247 VTAIL.n36 VTAIL.n35 11.249
R1248 VTAIL.n53 VTAIL.n6 11.249
R1249 VTAIL.n102 VTAIL.n101 11.249
R1250 VTAIL.n119 VTAIL.n72 11.249
R1251 VTAIL.n168 VTAIL.n167 11.249
R1252 VTAIL.n185 VTAIL.n138 11.249
R1253 VTAIL.n449 VTAIL.n402 11.249
R1254 VTAIL.n433 VTAIL.n432 11.249
R1255 VTAIL.n383 VTAIL.n336 11.249
R1256 VTAIL.n367 VTAIL.n366 11.249
R1257 VTAIL.n317 VTAIL.n270 11.249
R1258 VTAIL.n301 VTAIL.n300 11.249
R1259 VTAIL.n251 VTAIL.n204 11.249
R1260 VTAIL.n235 VTAIL.n234 11.249
R1261 VTAIL.n483 VTAIL.n482 10.7239
R1262 VTAIL.n21 VTAIL.n20 10.7239
R1263 VTAIL.n87 VTAIL.n86 10.7239
R1264 VTAIL.n153 VTAIL.n152 10.7239
R1265 VTAIL.n418 VTAIL.n417 10.7239
R1266 VTAIL.n352 VTAIL.n351 10.7239
R1267 VTAIL.n286 VTAIL.n285 10.7239
R1268 VTAIL.n220 VTAIL.n219 10.7239
R1269 VTAIL.n494 VTAIL.n476 10.4732
R1270 VTAIL.n516 VTAIL.n466 10.4732
R1271 VTAIL.n32 VTAIL.n14 10.4732
R1272 VTAIL.n54 VTAIL.n4 10.4732
R1273 VTAIL.n98 VTAIL.n80 10.4732
R1274 VTAIL.n120 VTAIL.n70 10.4732
R1275 VTAIL.n164 VTAIL.n146 10.4732
R1276 VTAIL.n186 VTAIL.n136 10.4732
R1277 VTAIL.n450 VTAIL.n400 10.4732
R1278 VTAIL.n429 VTAIL.n411 10.4732
R1279 VTAIL.n384 VTAIL.n334 10.4732
R1280 VTAIL.n363 VTAIL.n345 10.4732
R1281 VTAIL.n318 VTAIL.n268 10.4732
R1282 VTAIL.n297 VTAIL.n279 10.4732
R1283 VTAIL.n252 VTAIL.n202 10.4732
R1284 VTAIL.n231 VTAIL.n213 10.4732
R1285 VTAIL.n493 VTAIL.n478 9.69747
R1286 VTAIL.n520 VTAIL.n519 9.69747
R1287 VTAIL.n31 VTAIL.n16 9.69747
R1288 VTAIL.n58 VTAIL.n57 9.69747
R1289 VTAIL.n97 VTAIL.n82 9.69747
R1290 VTAIL.n124 VTAIL.n123 9.69747
R1291 VTAIL.n163 VTAIL.n148 9.69747
R1292 VTAIL.n190 VTAIL.n189 9.69747
R1293 VTAIL.n454 VTAIL.n453 9.69747
R1294 VTAIL.n428 VTAIL.n413 9.69747
R1295 VTAIL.n388 VTAIL.n387 9.69747
R1296 VTAIL.n362 VTAIL.n347 9.69747
R1297 VTAIL.n322 VTAIL.n321 9.69747
R1298 VTAIL.n296 VTAIL.n281 9.69747
R1299 VTAIL.n256 VTAIL.n255 9.69747
R1300 VTAIL.n230 VTAIL.n215 9.69747
R1301 VTAIL.n526 VTAIL.n525 9.45567
R1302 VTAIL.n64 VTAIL.n63 9.45567
R1303 VTAIL.n130 VTAIL.n129 9.45567
R1304 VTAIL.n196 VTAIL.n195 9.45567
R1305 VTAIL.n460 VTAIL.n459 9.45567
R1306 VTAIL.n394 VTAIL.n393 9.45567
R1307 VTAIL.n328 VTAIL.n327 9.45567
R1308 VTAIL.n262 VTAIL.n261 9.45567
R1309 VTAIL.n525 VTAIL.n524 9.3005
R1310 VTAIL.n464 VTAIL.n463 9.3005
R1311 VTAIL.n519 VTAIL.n518 9.3005
R1312 VTAIL.n517 VTAIL.n516 9.3005
R1313 VTAIL.n468 VTAIL.n467 9.3005
R1314 VTAIL.n511 VTAIL.n510 9.3005
R1315 VTAIL.n509 VTAIL.n508 9.3005
R1316 VTAIL.n485 VTAIL.n484 9.3005
R1317 VTAIL.n480 VTAIL.n479 9.3005
R1318 VTAIL.n491 VTAIL.n490 9.3005
R1319 VTAIL.n493 VTAIL.n492 9.3005
R1320 VTAIL.n476 VTAIL.n475 9.3005
R1321 VTAIL.n499 VTAIL.n498 9.3005
R1322 VTAIL.n501 VTAIL.n500 9.3005
R1323 VTAIL.n502 VTAIL.n471 9.3005
R1324 VTAIL.n63 VTAIL.n62 9.3005
R1325 VTAIL.n2 VTAIL.n1 9.3005
R1326 VTAIL.n57 VTAIL.n56 9.3005
R1327 VTAIL.n55 VTAIL.n54 9.3005
R1328 VTAIL.n6 VTAIL.n5 9.3005
R1329 VTAIL.n49 VTAIL.n48 9.3005
R1330 VTAIL.n47 VTAIL.n46 9.3005
R1331 VTAIL.n23 VTAIL.n22 9.3005
R1332 VTAIL.n18 VTAIL.n17 9.3005
R1333 VTAIL.n29 VTAIL.n28 9.3005
R1334 VTAIL.n31 VTAIL.n30 9.3005
R1335 VTAIL.n14 VTAIL.n13 9.3005
R1336 VTAIL.n37 VTAIL.n36 9.3005
R1337 VTAIL.n39 VTAIL.n38 9.3005
R1338 VTAIL.n40 VTAIL.n9 9.3005
R1339 VTAIL.n129 VTAIL.n128 9.3005
R1340 VTAIL.n68 VTAIL.n67 9.3005
R1341 VTAIL.n123 VTAIL.n122 9.3005
R1342 VTAIL.n121 VTAIL.n120 9.3005
R1343 VTAIL.n72 VTAIL.n71 9.3005
R1344 VTAIL.n115 VTAIL.n114 9.3005
R1345 VTAIL.n113 VTAIL.n112 9.3005
R1346 VTAIL.n89 VTAIL.n88 9.3005
R1347 VTAIL.n84 VTAIL.n83 9.3005
R1348 VTAIL.n95 VTAIL.n94 9.3005
R1349 VTAIL.n97 VTAIL.n96 9.3005
R1350 VTAIL.n80 VTAIL.n79 9.3005
R1351 VTAIL.n103 VTAIL.n102 9.3005
R1352 VTAIL.n105 VTAIL.n104 9.3005
R1353 VTAIL.n106 VTAIL.n75 9.3005
R1354 VTAIL.n195 VTAIL.n194 9.3005
R1355 VTAIL.n134 VTAIL.n133 9.3005
R1356 VTAIL.n189 VTAIL.n188 9.3005
R1357 VTAIL.n187 VTAIL.n186 9.3005
R1358 VTAIL.n138 VTAIL.n137 9.3005
R1359 VTAIL.n181 VTAIL.n180 9.3005
R1360 VTAIL.n179 VTAIL.n178 9.3005
R1361 VTAIL.n155 VTAIL.n154 9.3005
R1362 VTAIL.n150 VTAIL.n149 9.3005
R1363 VTAIL.n161 VTAIL.n160 9.3005
R1364 VTAIL.n163 VTAIL.n162 9.3005
R1365 VTAIL.n146 VTAIL.n145 9.3005
R1366 VTAIL.n169 VTAIL.n168 9.3005
R1367 VTAIL.n171 VTAIL.n170 9.3005
R1368 VTAIL.n172 VTAIL.n141 9.3005
R1369 VTAIL.n420 VTAIL.n419 9.3005
R1370 VTAIL.n415 VTAIL.n414 9.3005
R1371 VTAIL.n426 VTAIL.n425 9.3005
R1372 VTAIL.n428 VTAIL.n427 9.3005
R1373 VTAIL.n411 VTAIL.n410 9.3005
R1374 VTAIL.n434 VTAIL.n433 9.3005
R1375 VTAIL.n436 VTAIL.n435 9.3005
R1376 VTAIL.n408 VTAIL.n405 9.3005
R1377 VTAIL.n459 VTAIL.n458 9.3005
R1378 VTAIL.n398 VTAIL.n397 9.3005
R1379 VTAIL.n453 VTAIL.n452 9.3005
R1380 VTAIL.n451 VTAIL.n450 9.3005
R1381 VTAIL.n402 VTAIL.n401 9.3005
R1382 VTAIL.n445 VTAIL.n444 9.3005
R1383 VTAIL.n443 VTAIL.n442 9.3005
R1384 VTAIL.n354 VTAIL.n353 9.3005
R1385 VTAIL.n349 VTAIL.n348 9.3005
R1386 VTAIL.n360 VTAIL.n359 9.3005
R1387 VTAIL.n362 VTAIL.n361 9.3005
R1388 VTAIL.n345 VTAIL.n344 9.3005
R1389 VTAIL.n368 VTAIL.n367 9.3005
R1390 VTAIL.n370 VTAIL.n369 9.3005
R1391 VTAIL.n342 VTAIL.n339 9.3005
R1392 VTAIL.n393 VTAIL.n392 9.3005
R1393 VTAIL.n332 VTAIL.n331 9.3005
R1394 VTAIL.n387 VTAIL.n386 9.3005
R1395 VTAIL.n385 VTAIL.n384 9.3005
R1396 VTAIL.n336 VTAIL.n335 9.3005
R1397 VTAIL.n379 VTAIL.n378 9.3005
R1398 VTAIL.n377 VTAIL.n376 9.3005
R1399 VTAIL.n288 VTAIL.n287 9.3005
R1400 VTAIL.n283 VTAIL.n282 9.3005
R1401 VTAIL.n294 VTAIL.n293 9.3005
R1402 VTAIL.n296 VTAIL.n295 9.3005
R1403 VTAIL.n279 VTAIL.n278 9.3005
R1404 VTAIL.n302 VTAIL.n301 9.3005
R1405 VTAIL.n304 VTAIL.n303 9.3005
R1406 VTAIL.n276 VTAIL.n273 9.3005
R1407 VTAIL.n327 VTAIL.n326 9.3005
R1408 VTAIL.n266 VTAIL.n265 9.3005
R1409 VTAIL.n321 VTAIL.n320 9.3005
R1410 VTAIL.n319 VTAIL.n318 9.3005
R1411 VTAIL.n270 VTAIL.n269 9.3005
R1412 VTAIL.n313 VTAIL.n312 9.3005
R1413 VTAIL.n311 VTAIL.n310 9.3005
R1414 VTAIL.n222 VTAIL.n221 9.3005
R1415 VTAIL.n217 VTAIL.n216 9.3005
R1416 VTAIL.n228 VTAIL.n227 9.3005
R1417 VTAIL.n230 VTAIL.n229 9.3005
R1418 VTAIL.n213 VTAIL.n212 9.3005
R1419 VTAIL.n236 VTAIL.n235 9.3005
R1420 VTAIL.n238 VTAIL.n237 9.3005
R1421 VTAIL.n210 VTAIL.n207 9.3005
R1422 VTAIL.n261 VTAIL.n260 9.3005
R1423 VTAIL.n200 VTAIL.n199 9.3005
R1424 VTAIL.n255 VTAIL.n254 9.3005
R1425 VTAIL.n253 VTAIL.n252 9.3005
R1426 VTAIL.n204 VTAIL.n203 9.3005
R1427 VTAIL.n247 VTAIL.n246 9.3005
R1428 VTAIL.n245 VTAIL.n244 9.3005
R1429 VTAIL.n490 VTAIL.n489 8.92171
R1430 VTAIL.n523 VTAIL.n464 8.92171
R1431 VTAIL.n28 VTAIL.n27 8.92171
R1432 VTAIL.n61 VTAIL.n2 8.92171
R1433 VTAIL.n94 VTAIL.n93 8.92171
R1434 VTAIL.n127 VTAIL.n68 8.92171
R1435 VTAIL.n160 VTAIL.n159 8.92171
R1436 VTAIL.n193 VTAIL.n134 8.92171
R1437 VTAIL.n457 VTAIL.n398 8.92171
R1438 VTAIL.n425 VTAIL.n424 8.92171
R1439 VTAIL.n391 VTAIL.n332 8.92171
R1440 VTAIL.n359 VTAIL.n358 8.92171
R1441 VTAIL.n325 VTAIL.n266 8.92171
R1442 VTAIL.n293 VTAIL.n292 8.92171
R1443 VTAIL.n259 VTAIL.n200 8.92171
R1444 VTAIL.n227 VTAIL.n226 8.92171
R1445 VTAIL.n486 VTAIL.n480 8.14595
R1446 VTAIL.n524 VTAIL.n462 8.14595
R1447 VTAIL.n24 VTAIL.n18 8.14595
R1448 VTAIL.n62 VTAIL.n0 8.14595
R1449 VTAIL.n90 VTAIL.n84 8.14595
R1450 VTAIL.n128 VTAIL.n66 8.14595
R1451 VTAIL.n156 VTAIL.n150 8.14595
R1452 VTAIL.n194 VTAIL.n132 8.14595
R1453 VTAIL.n458 VTAIL.n396 8.14595
R1454 VTAIL.n421 VTAIL.n415 8.14595
R1455 VTAIL.n392 VTAIL.n330 8.14595
R1456 VTAIL.n355 VTAIL.n349 8.14595
R1457 VTAIL.n326 VTAIL.n264 8.14595
R1458 VTAIL.n289 VTAIL.n283 8.14595
R1459 VTAIL.n260 VTAIL.n198 8.14595
R1460 VTAIL.n223 VTAIL.n217 8.14595
R1461 VTAIL.n485 VTAIL.n482 7.3702
R1462 VTAIL.n23 VTAIL.n20 7.3702
R1463 VTAIL.n89 VTAIL.n86 7.3702
R1464 VTAIL.n155 VTAIL.n152 7.3702
R1465 VTAIL.n420 VTAIL.n417 7.3702
R1466 VTAIL.n354 VTAIL.n351 7.3702
R1467 VTAIL.n288 VTAIL.n285 7.3702
R1468 VTAIL.n222 VTAIL.n219 7.3702
R1469 VTAIL.n486 VTAIL.n485 5.81868
R1470 VTAIL.n526 VTAIL.n462 5.81868
R1471 VTAIL.n24 VTAIL.n23 5.81868
R1472 VTAIL.n64 VTAIL.n0 5.81868
R1473 VTAIL.n90 VTAIL.n89 5.81868
R1474 VTAIL.n130 VTAIL.n66 5.81868
R1475 VTAIL.n156 VTAIL.n155 5.81868
R1476 VTAIL.n196 VTAIL.n132 5.81868
R1477 VTAIL.n460 VTAIL.n396 5.81868
R1478 VTAIL.n421 VTAIL.n420 5.81868
R1479 VTAIL.n394 VTAIL.n330 5.81868
R1480 VTAIL.n355 VTAIL.n354 5.81868
R1481 VTAIL.n328 VTAIL.n264 5.81868
R1482 VTAIL.n289 VTAIL.n288 5.81868
R1483 VTAIL.n262 VTAIL.n198 5.81868
R1484 VTAIL.n223 VTAIL.n222 5.81868
R1485 VTAIL.n489 VTAIL.n480 5.04292
R1486 VTAIL.n524 VTAIL.n523 5.04292
R1487 VTAIL.n27 VTAIL.n18 5.04292
R1488 VTAIL.n62 VTAIL.n61 5.04292
R1489 VTAIL.n93 VTAIL.n84 5.04292
R1490 VTAIL.n128 VTAIL.n127 5.04292
R1491 VTAIL.n159 VTAIL.n150 5.04292
R1492 VTAIL.n194 VTAIL.n193 5.04292
R1493 VTAIL.n458 VTAIL.n457 5.04292
R1494 VTAIL.n424 VTAIL.n415 5.04292
R1495 VTAIL.n392 VTAIL.n391 5.04292
R1496 VTAIL.n358 VTAIL.n349 5.04292
R1497 VTAIL.n326 VTAIL.n325 5.04292
R1498 VTAIL.n292 VTAIL.n283 5.04292
R1499 VTAIL.n260 VTAIL.n259 5.04292
R1500 VTAIL.n226 VTAIL.n217 5.04292
R1501 VTAIL.n490 VTAIL.n478 4.26717
R1502 VTAIL.n520 VTAIL.n464 4.26717
R1503 VTAIL.n28 VTAIL.n16 4.26717
R1504 VTAIL.n58 VTAIL.n2 4.26717
R1505 VTAIL.n94 VTAIL.n82 4.26717
R1506 VTAIL.n124 VTAIL.n68 4.26717
R1507 VTAIL.n160 VTAIL.n148 4.26717
R1508 VTAIL.n190 VTAIL.n134 4.26717
R1509 VTAIL.n454 VTAIL.n398 4.26717
R1510 VTAIL.n425 VTAIL.n413 4.26717
R1511 VTAIL.n388 VTAIL.n332 4.26717
R1512 VTAIL.n359 VTAIL.n347 4.26717
R1513 VTAIL.n322 VTAIL.n266 4.26717
R1514 VTAIL.n293 VTAIL.n281 4.26717
R1515 VTAIL.n256 VTAIL.n200 4.26717
R1516 VTAIL.n227 VTAIL.n215 4.26717
R1517 VTAIL.n494 VTAIL.n493 3.49141
R1518 VTAIL.n519 VTAIL.n466 3.49141
R1519 VTAIL.n32 VTAIL.n31 3.49141
R1520 VTAIL.n57 VTAIL.n4 3.49141
R1521 VTAIL.n98 VTAIL.n97 3.49141
R1522 VTAIL.n123 VTAIL.n70 3.49141
R1523 VTAIL.n164 VTAIL.n163 3.49141
R1524 VTAIL.n189 VTAIL.n136 3.49141
R1525 VTAIL.n453 VTAIL.n400 3.49141
R1526 VTAIL.n429 VTAIL.n428 3.49141
R1527 VTAIL.n387 VTAIL.n334 3.49141
R1528 VTAIL.n363 VTAIL.n362 3.49141
R1529 VTAIL.n321 VTAIL.n268 3.49141
R1530 VTAIL.n297 VTAIL.n296 3.49141
R1531 VTAIL.n255 VTAIL.n202 3.49141
R1532 VTAIL.n231 VTAIL.n230 3.49141
R1533 VTAIL.n497 VTAIL.n476 2.71565
R1534 VTAIL.n516 VTAIL.n515 2.71565
R1535 VTAIL.n35 VTAIL.n14 2.71565
R1536 VTAIL.n54 VTAIL.n53 2.71565
R1537 VTAIL.n101 VTAIL.n80 2.71565
R1538 VTAIL.n120 VTAIL.n119 2.71565
R1539 VTAIL.n167 VTAIL.n146 2.71565
R1540 VTAIL.n186 VTAIL.n185 2.71565
R1541 VTAIL.n450 VTAIL.n449 2.71565
R1542 VTAIL.n432 VTAIL.n411 2.71565
R1543 VTAIL.n384 VTAIL.n383 2.71565
R1544 VTAIL.n366 VTAIL.n345 2.71565
R1545 VTAIL.n318 VTAIL.n317 2.71565
R1546 VTAIL.n300 VTAIL.n279 2.71565
R1547 VTAIL.n252 VTAIL.n251 2.71565
R1548 VTAIL.n234 VTAIL.n213 2.71565
R1549 VTAIL.n419 VTAIL.n418 2.41282
R1550 VTAIL.n353 VTAIL.n352 2.41282
R1551 VTAIL.n287 VTAIL.n286 2.41282
R1552 VTAIL.n221 VTAIL.n220 2.41282
R1553 VTAIL.n484 VTAIL.n483 2.41282
R1554 VTAIL.n22 VTAIL.n21 2.41282
R1555 VTAIL.n88 VTAIL.n87 2.41282
R1556 VTAIL.n154 VTAIL.n153 2.41282
R1557 VTAIL.n498 VTAIL.n474 1.93989
R1558 VTAIL.n512 VTAIL.n468 1.93989
R1559 VTAIL.n36 VTAIL.n12 1.93989
R1560 VTAIL.n50 VTAIL.n6 1.93989
R1561 VTAIL.n102 VTAIL.n78 1.93989
R1562 VTAIL.n116 VTAIL.n72 1.93989
R1563 VTAIL.n168 VTAIL.n144 1.93989
R1564 VTAIL.n182 VTAIL.n138 1.93989
R1565 VTAIL.n446 VTAIL.n402 1.93989
R1566 VTAIL.n433 VTAIL.n409 1.93989
R1567 VTAIL.n380 VTAIL.n336 1.93989
R1568 VTAIL.n367 VTAIL.n343 1.93989
R1569 VTAIL.n314 VTAIL.n270 1.93989
R1570 VTAIL.n301 VTAIL.n277 1.93989
R1571 VTAIL.n248 VTAIL.n204 1.93989
R1572 VTAIL.n235 VTAIL.n211 1.93989
R1573 VTAIL.n329 VTAIL.n263 1.65567
R1574 VTAIL.n461 VTAIL.n395 1.65567
R1575 VTAIL.n197 VTAIL.n131 1.65567
R1576 VTAIL.n503 VTAIL.n501 1.16414
R1577 VTAIL.n511 VTAIL.n470 1.16414
R1578 VTAIL.n41 VTAIL.n39 1.16414
R1579 VTAIL.n49 VTAIL.n8 1.16414
R1580 VTAIL.n107 VTAIL.n105 1.16414
R1581 VTAIL.n115 VTAIL.n74 1.16414
R1582 VTAIL.n173 VTAIL.n171 1.16414
R1583 VTAIL.n181 VTAIL.n140 1.16414
R1584 VTAIL.n445 VTAIL.n404 1.16414
R1585 VTAIL.n437 VTAIL.n436 1.16414
R1586 VTAIL.n379 VTAIL.n338 1.16414
R1587 VTAIL.n371 VTAIL.n370 1.16414
R1588 VTAIL.n313 VTAIL.n272 1.16414
R1589 VTAIL.n305 VTAIL.n304 1.16414
R1590 VTAIL.n247 VTAIL.n206 1.16414
R1591 VTAIL.n239 VTAIL.n238 1.16414
R1592 VTAIL VTAIL.n65 0.886276
R1593 VTAIL VTAIL.n527 0.769897
R1594 VTAIL.n395 VTAIL.n329 0.470328
R1595 VTAIL.n131 VTAIL.n65 0.470328
R1596 VTAIL.n502 VTAIL.n472 0.388379
R1597 VTAIL.n508 VTAIL.n507 0.388379
R1598 VTAIL.n40 VTAIL.n10 0.388379
R1599 VTAIL.n46 VTAIL.n45 0.388379
R1600 VTAIL.n106 VTAIL.n76 0.388379
R1601 VTAIL.n112 VTAIL.n111 0.388379
R1602 VTAIL.n172 VTAIL.n142 0.388379
R1603 VTAIL.n178 VTAIL.n177 0.388379
R1604 VTAIL.n442 VTAIL.n441 0.388379
R1605 VTAIL.n408 VTAIL.n406 0.388379
R1606 VTAIL.n376 VTAIL.n375 0.388379
R1607 VTAIL.n342 VTAIL.n340 0.388379
R1608 VTAIL.n310 VTAIL.n309 0.388379
R1609 VTAIL.n276 VTAIL.n274 0.388379
R1610 VTAIL.n244 VTAIL.n243 0.388379
R1611 VTAIL.n210 VTAIL.n208 0.388379
R1612 VTAIL.n484 VTAIL.n479 0.155672
R1613 VTAIL.n491 VTAIL.n479 0.155672
R1614 VTAIL.n492 VTAIL.n491 0.155672
R1615 VTAIL.n492 VTAIL.n475 0.155672
R1616 VTAIL.n499 VTAIL.n475 0.155672
R1617 VTAIL.n500 VTAIL.n499 0.155672
R1618 VTAIL.n500 VTAIL.n471 0.155672
R1619 VTAIL.n509 VTAIL.n471 0.155672
R1620 VTAIL.n510 VTAIL.n509 0.155672
R1621 VTAIL.n510 VTAIL.n467 0.155672
R1622 VTAIL.n517 VTAIL.n467 0.155672
R1623 VTAIL.n518 VTAIL.n517 0.155672
R1624 VTAIL.n518 VTAIL.n463 0.155672
R1625 VTAIL.n525 VTAIL.n463 0.155672
R1626 VTAIL.n22 VTAIL.n17 0.155672
R1627 VTAIL.n29 VTAIL.n17 0.155672
R1628 VTAIL.n30 VTAIL.n29 0.155672
R1629 VTAIL.n30 VTAIL.n13 0.155672
R1630 VTAIL.n37 VTAIL.n13 0.155672
R1631 VTAIL.n38 VTAIL.n37 0.155672
R1632 VTAIL.n38 VTAIL.n9 0.155672
R1633 VTAIL.n47 VTAIL.n9 0.155672
R1634 VTAIL.n48 VTAIL.n47 0.155672
R1635 VTAIL.n48 VTAIL.n5 0.155672
R1636 VTAIL.n55 VTAIL.n5 0.155672
R1637 VTAIL.n56 VTAIL.n55 0.155672
R1638 VTAIL.n56 VTAIL.n1 0.155672
R1639 VTAIL.n63 VTAIL.n1 0.155672
R1640 VTAIL.n88 VTAIL.n83 0.155672
R1641 VTAIL.n95 VTAIL.n83 0.155672
R1642 VTAIL.n96 VTAIL.n95 0.155672
R1643 VTAIL.n96 VTAIL.n79 0.155672
R1644 VTAIL.n103 VTAIL.n79 0.155672
R1645 VTAIL.n104 VTAIL.n103 0.155672
R1646 VTAIL.n104 VTAIL.n75 0.155672
R1647 VTAIL.n113 VTAIL.n75 0.155672
R1648 VTAIL.n114 VTAIL.n113 0.155672
R1649 VTAIL.n114 VTAIL.n71 0.155672
R1650 VTAIL.n121 VTAIL.n71 0.155672
R1651 VTAIL.n122 VTAIL.n121 0.155672
R1652 VTAIL.n122 VTAIL.n67 0.155672
R1653 VTAIL.n129 VTAIL.n67 0.155672
R1654 VTAIL.n154 VTAIL.n149 0.155672
R1655 VTAIL.n161 VTAIL.n149 0.155672
R1656 VTAIL.n162 VTAIL.n161 0.155672
R1657 VTAIL.n162 VTAIL.n145 0.155672
R1658 VTAIL.n169 VTAIL.n145 0.155672
R1659 VTAIL.n170 VTAIL.n169 0.155672
R1660 VTAIL.n170 VTAIL.n141 0.155672
R1661 VTAIL.n179 VTAIL.n141 0.155672
R1662 VTAIL.n180 VTAIL.n179 0.155672
R1663 VTAIL.n180 VTAIL.n137 0.155672
R1664 VTAIL.n187 VTAIL.n137 0.155672
R1665 VTAIL.n188 VTAIL.n187 0.155672
R1666 VTAIL.n188 VTAIL.n133 0.155672
R1667 VTAIL.n195 VTAIL.n133 0.155672
R1668 VTAIL.n459 VTAIL.n397 0.155672
R1669 VTAIL.n452 VTAIL.n397 0.155672
R1670 VTAIL.n452 VTAIL.n451 0.155672
R1671 VTAIL.n451 VTAIL.n401 0.155672
R1672 VTAIL.n444 VTAIL.n401 0.155672
R1673 VTAIL.n444 VTAIL.n443 0.155672
R1674 VTAIL.n443 VTAIL.n405 0.155672
R1675 VTAIL.n435 VTAIL.n405 0.155672
R1676 VTAIL.n435 VTAIL.n434 0.155672
R1677 VTAIL.n434 VTAIL.n410 0.155672
R1678 VTAIL.n427 VTAIL.n410 0.155672
R1679 VTAIL.n427 VTAIL.n426 0.155672
R1680 VTAIL.n426 VTAIL.n414 0.155672
R1681 VTAIL.n419 VTAIL.n414 0.155672
R1682 VTAIL.n393 VTAIL.n331 0.155672
R1683 VTAIL.n386 VTAIL.n331 0.155672
R1684 VTAIL.n386 VTAIL.n385 0.155672
R1685 VTAIL.n385 VTAIL.n335 0.155672
R1686 VTAIL.n378 VTAIL.n335 0.155672
R1687 VTAIL.n378 VTAIL.n377 0.155672
R1688 VTAIL.n377 VTAIL.n339 0.155672
R1689 VTAIL.n369 VTAIL.n339 0.155672
R1690 VTAIL.n369 VTAIL.n368 0.155672
R1691 VTAIL.n368 VTAIL.n344 0.155672
R1692 VTAIL.n361 VTAIL.n344 0.155672
R1693 VTAIL.n361 VTAIL.n360 0.155672
R1694 VTAIL.n360 VTAIL.n348 0.155672
R1695 VTAIL.n353 VTAIL.n348 0.155672
R1696 VTAIL.n327 VTAIL.n265 0.155672
R1697 VTAIL.n320 VTAIL.n265 0.155672
R1698 VTAIL.n320 VTAIL.n319 0.155672
R1699 VTAIL.n319 VTAIL.n269 0.155672
R1700 VTAIL.n312 VTAIL.n269 0.155672
R1701 VTAIL.n312 VTAIL.n311 0.155672
R1702 VTAIL.n311 VTAIL.n273 0.155672
R1703 VTAIL.n303 VTAIL.n273 0.155672
R1704 VTAIL.n303 VTAIL.n302 0.155672
R1705 VTAIL.n302 VTAIL.n278 0.155672
R1706 VTAIL.n295 VTAIL.n278 0.155672
R1707 VTAIL.n295 VTAIL.n294 0.155672
R1708 VTAIL.n294 VTAIL.n282 0.155672
R1709 VTAIL.n287 VTAIL.n282 0.155672
R1710 VTAIL.n261 VTAIL.n199 0.155672
R1711 VTAIL.n254 VTAIL.n199 0.155672
R1712 VTAIL.n254 VTAIL.n253 0.155672
R1713 VTAIL.n253 VTAIL.n203 0.155672
R1714 VTAIL.n246 VTAIL.n203 0.155672
R1715 VTAIL.n246 VTAIL.n245 0.155672
R1716 VTAIL.n245 VTAIL.n207 0.155672
R1717 VTAIL.n237 VTAIL.n207 0.155672
R1718 VTAIL.n237 VTAIL.n236 0.155672
R1719 VTAIL.n236 VTAIL.n212 0.155672
R1720 VTAIL.n229 VTAIL.n212 0.155672
R1721 VTAIL.n229 VTAIL.n228 0.155672
R1722 VTAIL.n228 VTAIL.n216 0.155672
R1723 VTAIL.n221 VTAIL.n216 0.155672
R1724 VN.n0 VN.t3 222.115
R1725 VN.n1 VN.t1 222.115
R1726 VN.n0 VN.t0 221.791
R1727 VN.n1 VN.t2 221.791
R1728 VN VN.n1 56.4182
R1729 VN VN.n0 12.7478
R1730 VDD2.n2 VDD2.n0 113.981
R1731 VDD2.n2 VDD2.n1 74.8087
R1732 VDD2.n1 VDD2.t1 2.67141
R1733 VDD2.n1 VDD2.t2 2.67141
R1734 VDD2.n0 VDD2.t0 2.67141
R1735 VDD2.n0 VDD2.t3 2.67141
R1736 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 4.48848f
C1 VTAIL w_n2122_n3402# 4.041f
C2 VTAIL B 4.479741f
C3 VTAIL VDD2 5.58497f
C4 VTAIL VN 4.0658f
C5 VTAIL VP 4.07991f
C6 B w_n2122_n3402# 8.05067f
C7 VDD2 w_n2122_n3402# 1.29426f
C8 w_n2122_n3402# VN 3.40399f
C9 VTAIL VDD1 5.53754f
C10 VDD2 B 1.1243f
C11 B VN 0.918972f
C12 VDD2 VN 4.30701f
C13 VP w_n2122_n3402# 3.67423f
C14 VP B 1.36272f
C15 VDD2 VP 0.330157f
C16 VDD1 w_n2122_n3402# 1.26074f
C17 VP VN 5.49268f
C18 VDD1 B 1.08864f
C19 VDD1 VDD2 0.781878f
C20 VDD1 VN 0.148207f
C21 VDD2 VSUBS 0.795976f
C22 VDD1 VSUBS 5.208459f
C23 VTAIL VSUBS 1.068689f
C24 VN VSUBS 5.18652f
C25 VP VSUBS 1.752251f
C26 B VSUBS 3.416935f
C27 w_n2122_n3402# VSUBS 88.843895f
C28 VDD2.t0 VSUBS 0.256969f
C29 VDD2.t3 VSUBS 0.256969f
C30 VDD2.n0 VSUBS 2.66288f
C31 VDD2.t1 VSUBS 0.256969f
C32 VDD2.t2 VSUBS 0.256969f
C33 VDD2.n1 VSUBS 2.01314f
C34 VDD2.n2 VSUBS 4.04784f
C35 VN.t3 VSUBS 2.40602f
C36 VN.t0 VSUBS 2.40456f
C37 VN.n0 VSUBS 1.71037f
C38 VN.t1 VSUBS 2.40602f
C39 VN.t2 VSUBS 2.40456f
C40 VN.n1 VSUBS 3.34485f
C41 VTAIL.n0 VSUBS 0.025615f
C42 VTAIL.n1 VSUBS 0.022956f
C43 VTAIL.n2 VSUBS 0.012336f
C44 VTAIL.n3 VSUBS 0.029157f
C45 VTAIL.n4 VSUBS 0.013061f
C46 VTAIL.n5 VSUBS 0.022956f
C47 VTAIL.n6 VSUBS 0.012336f
C48 VTAIL.n7 VSUBS 0.029157f
C49 VTAIL.n8 VSUBS 0.013061f
C50 VTAIL.n9 VSUBS 0.022956f
C51 VTAIL.n10 VSUBS 0.012699f
C52 VTAIL.n11 VSUBS 0.029157f
C53 VTAIL.n12 VSUBS 0.013061f
C54 VTAIL.n13 VSUBS 0.022956f
C55 VTAIL.n14 VSUBS 0.012336f
C56 VTAIL.n15 VSUBS 0.029157f
C57 VTAIL.n16 VSUBS 0.013061f
C58 VTAIL.n17 VSUBS 0.022956f
C59 VTAIL.n18 VSUBS 0.012336f
C60 VTAIL.n19 VSUBS 0.021868f
C61 VTAIL.n20 VSUBS 0.021934f
C62 VTAIL.t3 VSUBS 0.062845f
C63 VTAIL.n21 VSUBS 0.182561f
C64 VTAIL.n22 VSUBS 1.14502f
C65 VTAIL.n23 VSUBS 0.012336f
C66 VTAIL.n24 VSUBS 0.013061f
C67 VTAIL.n25 VSUBS 0.029157f
C68 VTAIL.n26 VSUBS 0.029157f
C69 VTAIL.n27 VSUBS 0.013061f
C70 VTAIL.n28 VSUBS 0.012336f
C71 VTAIL.n29 VSUBS 0.022956f
C72 VTAIL.n30 VSUBS 0.022956f
C73 VTAIL.n31 VSUBS 0.012336f
C74 VTAIL.n32 VSUBS 0.013061f
C75 VTAIL.n33 VSUBS 0.029157f
C76 VTAIL.n34 VSUBS 0.029157f
C77 VTAIL.n35 VSUBS 0.013061f
C78 VTAIL.n36 VSUBS 0.012336f
C79 VTAIL.n37 VSUBS 0.022956f
C80 VTAIL.n38 VSUBS 0.022956f
C81 VTAIL.n39 VSUBS 0.012336f
C82 VTAIL.n40 VSUBS 0.012336f
C83 VTAIL.n41 VSUBS 0.013061f
C84 VTAIL.n42 VSUBS 0.029157f
C85 VTAIL.n43 VSUBS 0.029157f
C86 VTAIL.n44 VSUBS 0.029157f
C87 VTAIL.n45 VSUBS 0.012699f
C88 VTAIL.n46 VSUBS 0.012336f
C89 VTAIL.n47 VSUBS 0.022956f
C90 VTAIL.n48 VSUBS 0.022956f
C91 VTAIL.n49 VSUBS 0.012336f
C92 VTAIL.n50 VSUBS 0.013061f
C93 VTAIL.n51 VSUBS 0.029157f
C94 VTAIL.n52 VSUBS 0.029157f
C95 VTAIL.n53 VSUBS 0.013061f
C96 VTAIL.n54 VSUBS 0.012336f
C97 VTAIL.n55 VSUBS 0.022956f
C98 VTAIL.n56 VSUBS 0.022956f
C99 VTAIL.n57 VSUBS 0.012336f
C100 VTAIL.n58 VSUBS 0.013061f
C101 VTAIL.n59 VSUBS 0.029157f
C102 VTAIL.n60 VSUBS 0.071917f
C103 VTAIL.n61 VSUBS 0.013061f
C104 VTAIL.n62 VSUBS 0.012336f
C105 VTAIL.n63 VSUBS 0.054631f
C106 VTAIL.n64 VSUBS 0.036273f
C107 VTAIL.n65 VSUBS 0.120767f
C108 VTAIL.n66 VSUBS 0.025615f
C109 VTAIL.n67 VSUBS 0.022956f
C110 VTAIL.n68 VSUBS 0.012336f
C111 VTAIL.n69 VSUBS 0.029157f
C112 VTAIL.n70 VSUBS 0.013061f
C113 VTAIL.n71 VSUBS 0.022956f
C114 VTAIL.n72 VSUBS 0.012336f
C115 VTAIL.n73 VSUBS 0.029157f
C116 VTAIL.n74 VSUBS 0.013061f
C117 VTAIL.n75 VSUBS 0.022956f
C118 VTAIL.n76 VSUBS 0.012699f
C119 VTAIL.n77 VSUBS 0.029157f
C120 VTAIL.n78 VSUBS 0.013061f
C121 VTAIL.n79 VSUBS 0.022956f
C122 VTAIL.n80 VSUBS 0.012336f
C123 VTAIL.n81 VSUBS 0.029157f
C124 VTAIL.n82 VSUBS 0.013061f
C125 VTAIL.n83 VSUBS 0.022956f
C126 VTAIL.n84 VSUBS 0.012336f
C127 VTAIL.n85 VSUBS 0.021868f
C128 VTAIL.n86 VSUBS 0.021934f
C129 VTAIL.t6 VSUBS 0.062845f
C130 VTAIL.n87 VSUBS 0.182561f
C131 VTAIL.n88 VSUBS 1.14502f
C132 VTAIL.n89 VSUBS 0.012336f
C133 VTAIL.n90 VSUBS 0.013061f
C134 VTAIL.n91 VSUBS 0.029157f
C135 VTAIL.n92 VSUBS 0.029157f
C136 VTAIL.n93 VSUBS 0.013061f
C137 VTAIL.n94 VSUBS 0.012336f
C138 VTAIL.n95 VSUBS 0.022956f
C139 VTAIL.n96 VSUBS 0.022956f
C140 VTAIL.n97 VSUBS 0.012336f
C141 VTAIL.n98 VSUBS 0.013061f
C142 VTAIL.n99 VSUBS 0.029157f
C143 VTAIL.n100 VSUBS 0.029157f
C144 VTAIL.n101 VSUBS 0.013061f
C145 VTAIL.n102 VSUBS 0.012336f
C146 VTAIL.n103 VSUBS 0.022956f
C147 VTAIL.n104 VSUBS 0.022956f
C148 VTAIL.n105 VSUBS 0.012336f
C149 VTAIL.n106 VSUBS 0.012336f
C150 VTAIL.n107 VSUBS 0.013061f
C151 VTAIL.n108 VSUBS 0.029157f
C152 VTAIL.n109 VSUBS 0.029157f
C153 VTAIL.n110 VSUBS 0.029157f
C154 VTAIL.n111 VSUBS 0.012699f
C155 VTAIL.n112 VSUBS 0.012336f
C156 VTAIL.n113 VSUBS 0.022956f
C157 VTAIL.n114 VSUBS 0.022956f
C158 VTAIL.n115 VSUBS 0.012336f
C159 VTAIL.n116 VSUBS 0.013061f
C160 VTAIL.n117 VSUBS 0.029157f
C161 VTAIL.n118 VSUBS 0.029157f
C162 VTAIL.n119 VSUBS 0.013061f
C163 VTAIL.n120 VSUBS 0.012336f
C164 VTAIL.n121 VSUBS 0.022956f
C165 VTAIL.n122 VSUBS 0.022956f
C166 VTAIL.n123 VSUBS 0.012336f
C167 VTAIL.n124 VSUBS 0.013061f
C168 VTAIL.n125 VSUBS 0.029157f
C169 VTAIL.n126 VSUBS 0.071917f
C170 VTAIL.n127 VSUBS 0.013061f
C171 VTAIL.n128 VSUBS 0.012336f
C172 VTAIL.n129 VSUBS 0.054631f
C173 VTAIL.n130 VSUBS 0.036273f
C174 VTAIL.n131 VSUBS 0.17768f
C175 VTAIL.n132 VSUBS 0.025615f
C176 VTAIL.n133 VSUBS 0.022956f
C177 VTAIL.n134 VSUBS 0.012336f
C178 VTAIL.n135 VSUBS 0.029157f
C179 VTAIL.n136 VSUBS 0.013061f
C180 VTAIL.n137 VSUBS 0.022956f
C181 VTAIL.n138 VSUBS 0.012336f
C182 VTAIL.n139 VSUBS 0.029157f
C183 VTAIL.n140 VSUBS 0.013061f
C184 VTAIL.n141 VSUBS 0.022956f
C185 VTAIL.n142 VSUBS 0.012699f
C186 VTAIL.n143 VSUBS 0.029157f
C187 VTAIL.n144 VSUBS 0.013061f
C188 VTAIL.n145 VSUBS 0.022956f
C189 VTAIL.n146 VSUBS 0.012336f
C190 VTAIL.n147 VSUBS 0.029157f
C191 VTAIL.n148 VSUBS 0.013061f
C192 VTAIL.n149 VSUBS 0.022956f
C193 VTAIL.n150 VSUBS 0.012336f
C194 VTAIL.n151 VSUBS 0.021868f
C195 VTAIL.n152 VSUBS 0.021934f
C196 VTAIL.t7 VSUBS 0.062845f
C197 VTAIL.n153 VSUBS 0.182561f
C198 VTAIL.n154 VSUBS 1.14502f
C199 VTAIL.n155 VSUBS 0.012336f
C200 VTAIL.n156 VSUBS 0.013061f
C201 VTAIL.n157 VSUBS 0.029157f
C202 VTAIL.n158 VSUBS 0.029157f
C203 VTAIL.n159 VSUBS 0.013061f
C204 VTAIL.n160 VSUBS 0.012336f
C205 VTAIL.n161 VSUBS 0.022956f
C206 VTAIL.n162 VSUBS 0.022956f
C207 VTAIL.n163 VSUBS 0.012336f
C208 VTAIL.n164 VSUBS 0.013061f
C209 VTAIL.n165 VSUBS 0.029157f
C210 VTAIL.n166 VSUBS 0.029157f
C211 VTAIL.n167 VSUBS 0.013061f
C212 VTAIL.n168 VSUBS 0.012336f
C213 VTAIL.n169 VSUBS 0.022956f
C214 VTAIL.n170 VSUBS 0.022956f
C215 VTAIL.n171 VSUBS 0.012336f
C216 VTAIL.n172 VSUBS 0.012336f
C217 VTAIL.n173 VSUBS 0.013061f
C218 VTAIL.n174 VSUBS 0.029157f
C219 VTAIL.n175 VSUBS 0.029157f
C220 VTAIL.n176 VSUBS 0.029157f
C221 VTAIL.n177 VSUBS 0.012699f
C222 VTAIL.n178 VSUBS 0.012336f
C223 VTAIL.n179 VSUBS 0.022956f
C224 VTAIL.n180 VSUBS 0.022956f
C225 VTAIL.n181 VSUBS 0.012336f
C226 VTAIL.n182 VSUBS 0.013061f
C227 VTAIL.n183 VSUBS 0.029157f
C228 VTAIL.n184 VSUBS 0.029157f
C229 VTAIL.n185 VSUBS 0.013061f
C230 VTAIL.n186 VSUBS 0.012336f
C231 VTAIL.n187 VSUBS 0.022956f
C232 VTAIL.n188 VSUBS 0.022956f
C233 VTAIL.n189 VSUBS 0.012336f
C234 VTAIL.n190 VSUBS 0.013061f
C235 VTAIL.n191 VSUBS 0.029157f
C236 VTAIL.n192 VSUBS 0.071917f
C237 VTAIL.n193 VSUBS 0.013061f
C238 VTAIL.n194 VSUBS 0.012336f
C239 VTAIL.n195 VSUBS 0.054631f
C240 VTAIL.n196 VSUBS 0.036273f
C241 VTAIL.n197 VSUBS 1.35325f
C242 VTAIL.n198 VSUBS 0.025615f
C243 VTAIL.n199 VSUBS 0.022956f
C244 VTAIL.n200 VSUBS 0.012336f
C245 VTAIL.n201 VSUBS 0.029157f
C246 VTAIL.n202 VSUBS 0.013061f
C247 VTAIL.n203 VSUBS 0.022956f
C248 VTAIL.n204 VSUBS 0.012336f
C249 VTAIL.n205 VSUBS 0.029157f
C250 VTAIL.n206 VSUBS 0.013061f
C251 VTAIL.n207 VSUBS 0.022956f
C252 VTAIL.n208 VSUBS 0.012699f
C253 VTAIL.n209 VSUBS 0.029157f
C254 VTAIL.n210 VSUBS 0.012336f
C255 VTAIL.n211 VSUBS 0.013061f
C256 VTAIL.n212 VSUBS 0.022956f
C257 VTAIL.n213 VSUBS 0.012336f
C258 VTAIL.n214 VSUBS 0.029157f
C259 VTAIL.n215 VSUBS 0.013061f
C260 VTAIL.n216 VSUBS 0.022956f
C261 VTAIL.n217 VSUBS 0.012336f
C262 VTAIL.n218 VSUBS 0.021868f
C263 VTAIL.n219 VSUBS 0.021934f
C264 VTAIL.t0 VSUBS 0.062845f
C265 VTAIL.n220 VSUBS 0.182561f
C266 VTAIL.n221 VSUBS 1.14502f
C267 VTAIL.n222 VSUBS 0.012336f
C268 VTAIL.n223 VSUBS 0.013061f
C269 VTAIL.n224 VSUBS 0.029157f
C270 VTAIL.n225 VSUBS 0.029157f
C271 VTAIL.n226 VSUBS 0.013061f
C272 VTAIL.n227 VSUBS 0.012336f
C273 VTAIL.n228 VSUBS 0.022956f
C274 VTAIL.n229 VSUBS 0.022956f
C275 VTAIL.n230 VSUBS 0.012336f
C276 VTAIL.n231 VSUBS 0.013061f
C277 VTAIL.n232 VSUBS 0.029157f
C278 VTAIL.n233 VSUBS 0.029157f
C279 VTAIL.n234 VSUBS 0.013061f
C280 VTAIL.n235 VSUBS 0.012336f
C281 VTAIL.n236 VSUBS 0.022956f
C282 VTAIL.n237 VSUBS 0.022956f
C283 VTAIL.n238 VSUBS 0.012336f
C284 VTAIL.n239 VSUBS 0.013061f
C285 VTAIL.n240 VSUBS 0.029157f
C286 VTAIL.n241 VSUBS 0.029157f
C287 VTAIL.n242 VSUBS 0.029157f
C288 VTAIL.n243 VSUBS 0.012699f
C289 VTAIL.n244 VSUBS 0.012336f
C290 VTAIL.n245 VSUBS 0.022956f
C291 VTAIL.n246 VSUBS 0.022956f
C292 VTAIL.n247 VSUBS 0.012336f
C293 VTAIL.n248 VSUBS 0.013061f
C294 VTAIL.n249 VSUBS 0.029157f
C295 VTAIL.n250 VSUBS 0.029157f
C296 VTAIL.n251 VSUBS 0.013061f
C297 VTAIL.n252 VSUBS 0.012336f
C298 VTAIL.n253 VSUBS 0.022956f
C299 VTAIL.n254 VSUBS 0.022956f
C300 VTAIL.n255 VSUBS 0.012336f
C301 VTAIL.n256 VSUBS 0.013061f
C302 VTAIL.n257 VSUBS 0.029157f
C303 VTAIL.n258 VSUBS 0.071917f
C304 VTAIL.n259 VSUBS 0.013061f
C305 VTAIL.n260 VSUBS 0.012336f
C306 VTAIL.n261 VSUBS 0.054631f
C307 VTAIL.n262 VSUBS 0.036273f
C308 VTAIL.n263 VSUBS 1.35325f
C309 VTAIL.n264 VSUBS 0.025615f
C310 VTAIL.n265 VSUBS 0.022956f
C311 VTAIL.n266 VSUBS 0.012336f
C312 VTAIL.n267 VSUBS 0.029157f
C313 VTAIL.n268 VSUBS 0.013061f
C314 VTAIL.n269 VSUBS 0.022956f
C315 VTAIL.n270 VSUBS 0.012336f
C316 VTAIL.n271 VSUBS 0.029157f
C317 VTAIL.n272 VSUBS 0.013061f
C318 VTAIL.n273 VSUBS 0.022956f
C319 VTAIL.n274 VSUBS 0.012699f
C320 VTAIL.n275 VSUBS 0.029157f
C321 VTAIL.n276 VSUBS 0.012336f
C322 VTAIL.n277 VSUBS 0.013061f
C323 VTAIL.n278 VSUBS 0.022956f
C324 VTAIL.n279 VSUBS 0.012336f
C325 VTAIL.n280 VSUBS 0.029157f
C326 VTAIL.n281 VSUBS 0.013061f
C327 VTAIL.n282 VSUBS 0.022956f
C328 VTAIL.n283 VSUBS 0.012336f
C329 VTAIL.n284 VSUBS 0.021868f
C330 VTAIL.n285 VSUBS 0.021934f
C331 VTAIL.t1 VSUBS 0.062845f
C332 VTAIL.n286 VSUBS 0.182561f
C333 VTAIL.n287 VSUBS 1.14502f
C334 VTAIL.n288 VSUBS 0.012336f
C335 VTAIL.n289 VSUBS 0.013061f
C336 VTAIL.n290 VSUBS 0.029157f
C337 VTAIL.n291 VSUBS 0.029157f
C338 VTAIL.n292 VSUBS 0.013061f
C339 VTAIL.n293 VSUBS 0.012336f
C340 VTAIL.n294 VSUBS 0.022956f
C341 VTAIL.n295 VSUBS 0.022956f
C342 VTAIL.n296 VSUBS 0.012336f
C343 VTAIL.n297 VSUBS 0.013061f
C344 VTAIL.n298 VSUBS 0.029157f
C345 VTAIL.n299 VSUBS 0.029157f
C346 VTAIL.n300 VSUBS 0.013061f
C347 VTAIL.n301 VSUBS 0.012336f
C348 VTAIL.n302 VSUBS 0.022956f
C349 VTAIL.n303 VSUBS 0.022956f
C350 VTAIL.n304 VSUBS 0.012336f
C351 VTAIL.n305 VSUBS 0.013061f
C352 VTAIL.n306 VSUBS 0.029157f
C353 VTAIL.n307 VSUBS 0.029157f
C354 VTAIL.n308 VSUBS 0.029157f
C355 VTAIL.n309 VSUBS 0.012699f
C356 VTAIL.n310 VSUBS 0.012336f
C357 VTAIL.n311 VSUBS 0.022956f
C358 VTAIL.n312 VSUBS 0.022956f
C359 VTAIL.n313 VSUBS 0.012336f
C360 VTAIL.n314 VSUBS 0.013061f
C361 VTAIL.n315 VSUBS 0.029157f
C362 VTAIL.n316 VSUBS 0.029157f
C363 VTAIL.n317 VSUBS 0.013061f
C364 VTAIL.n318 VSUBS 0.012336f
C365 VTAIL.n319 VSUBS 0.022956f
C366 VTAIL.n320 VSUBS 0.022956f
C367 VTAIL.n321 VSUBS 0.012336f
C368 VTAIL.n322 VSUBS 0.013061f
C369 VTAIL.n323 VSUBS 0.029157f
C370 VTAIL.n324 VSUBS 0.071917f
C371 VTAIL.n325 VSUBS 0.013061f
C372 VTAIL.n326 VSUBS 0.012336f
C373 VTAIL.n327 VSUBS 0.054631f
C374 VTAIL.n328 VSUBS 0.036273f
C375 VTAIL.n329 VSUBS 0.17768f
C376 VTAIL.n330 VSUBS 0.025615f
C377 VTAIL.n331 VSUBS 0.022956f
C378 VTAIL.n332 VSUBS 0.012336f
C379 VTAIL.n333 VSUBS 0.029157f
C380 VTAIL.n334 VSUBS 0.013061f
C381 VTAIL.n335 VSUBS 0.022956f
C382 VTAIL.n336 VSUBS 0.012336f
C383 VTAIL.n337 VSUBS 0.029157f
C384 VTAIL.n338 VSUBS 0.013061f
C385 VTAIL.n339 VSUBS 0.022956f
C386 VTAIL.n340 VSUBS 0.012699f
C387 VTAIL.n341 VSUBS 0.029157f
C388 VTAIL.n342 VSUBS 0.012336f
C389 VTAIL.n343 VSUBS 0.013061f
C390 VTAIL.n344 VSUBS 0.022956f
C391 VTAIL.n345 VSUBS 0.012336f
C392 VTAIL.n346 VSUBS 0.029157f
C393 VTAIL.n347 VSUBS 0.013061f
C394 VTAIL.n348 VSUBS 0.022956f
C395 VTAIL.n349 VSUBS 0.012336f
C396 VTAIL.n350 VSUBS 0.021868f
C397 VTAIL.n351 VSUBS 0.021934f
C398 VTAIL.t4 VSUBS 0.062845f
C399 VTAIL.n352 VSUBS 0.182561f
C400 VTAIL.n353 VSUBS 1.14502f
C401 VTAIL.n354 VSUBS 0.012336f
C402 VTAIL.n355 VSUBS 0.013061f
C403 VTAIL.n356 VSUBS 0.029157f
C404 VTAIL.n357 VSUBS 0.029157f
C405 VTAIL.n358 VSUBS 0.013061f
C406 VTAIL.n359 VSUBS 0.012336f
C407 VTAIL.n360 VSUBS 0.022956f
C408 VTAIL.n361 VSUBS 0.022956f
C409 VTAIL.n362 VSUBS 0.012336f
C410 VTAIL.n363 VSUBS 0.013061f
C411 VTAIL.n364 VSUBS 0.029157f
C412 VTAIL.n365 VSUBS 0.029157f
C413 VTAIL.n366 VSUBS 0.013061f
C414 VTAIL.n367 VSUBS 0.012336f
C415 VTAIL.n368 VSUBS 0.022956f
C416 VTAIL.n369 VSUBS 0.022956f
C417 VTAIL.n370 VSUBS 0.012336f
C418 VTAIL.n371 VSUBS 0.013061f
C419 VTAIL.n372 VSUBS 0.029157f
C420 VTAIL.n373 VSUBS 0.029157f
C421 VTAIL.n374 VSUBS 0.029157f
C422 VTAIL.n375 VSUBS 0.012699f
C423 VTAIL.n376 VSUBS 0.012336f
C424 VTAIL.n377 VSUBS 0.022956f
C425 VTAIL.n378 VSUBS 0.022956f
C426 VTAIL.n379 VSUBS 0.012336f
C427 VTAIL.n380 VSUBS 0.013061f
C428 VTAIL.n381 VSUBS 0.029157f
C429 VTAIL.n382 VSUBS 0.029157f
C430 VTAIL.n383 VSUBS 0.013061f
C431 VTAIL.n384 VSUBS 0.012336f
C432 VTAIL.n385 VSUBS 0.022956f
C433 VTAIL.n386 VSUBS 0.022956f
C434 VTAIL.n387 VSUBS 0.012336f
C435 VTAIL.n388 VSUBS 0.013061f
C436 VTAIL.n389 VSUBS 0.029157f
C437 VTAIL.n390 VSUBS 0.071917f
C438 VTAIL.n391 VSUBS 0.013061f
C439 VTAIL.n392 VSUBS 0.012336f
C440 VTAIL.n393 VSUBS 0.054631f
C441 VTAIL.n394 VSUBS 0.036273f
C442 VTAIL.n395 VSUBS 0.17768f
C443 VTAIL.n396 VSUBS 0.025615f
C444 VTAIL.n397 VSUBS 0.022956f
C445 VTAIL.n398 VSUBS 0.012336f
C446 VTAIL.n399 VSUBS 0.029157f
C447 VTAIL.n400 VSUBS 0.013061f
C448 VTAIL.n401 VSUBS 0.022956f
C449 VTAIL.n402 VSUBS 0.012336f
C450 VTAIL.n403 VSUBS 0.029157f
C451 VTAIL.n404 VSUBS 0.013061f
C452 VTAIL.n405 VSUBS 0.022956f
C453 VTAIL.n406 VSUBS 0.012699f
C454 VTAIL.n407 VSUBS 0.029157f
C455 VTAIL.n408 VSUBS 0.012336f
C456 VTAIL.n409 VSUBS 0.013061f
C457 VTAIL.n410 VSUBS 0.022956f
C458 VTAIL.n411 VSUBS 0.012336f
C459 VTAIL.n412 VSUBS 0.029157f
C460 VTAIL.n413 VSUBS 0.013061f
C461 VTAIL.n414 VSUBS 0.022956f
C462 VTAIL.n415 VSUBS 0.012336f
C463 VTAIL.n416 VSUBS 0.021868f
C464 VTAIL.n417 VSUBS 0.021934f
C465 VTAIL.t5 VSUBS 0.062845f
C466 VTAIL.n418 VSUBS 0.182561f
C467 VTAIL.n419 VSUBS 1.14502f
C468 VTAIL.n420 VSUBS 0.012336f
C469 VTAIL.n421 VSUBS 0.013061f
C470 VTAIL.n422 VSUBS 0.029157f
C471 VTAIL.n423 VSUBS 0.029157f
C472 VTAIL.n424 VSUBS 0.013061f
C473 VTAIL.n425 VSUBS 0.012336f
C474 VTAIL.n426 VSUBS 0.022956f
C475 VTAIL.n427 VSUBS 0.022956f
C476 VTAIL.n428 VSUBS 0.012336f
C477 VTAIL.n429 VSUBS 0.013061f
C478 VTAIL.n430 VSUBS 0.029157f
C479 VTAIL.n431 VSUBS 0.029157f
C480 VTAIL.n432 VSUBS 0.013061f
C481 VTAIL.n433 VSUBS 0.012336f
C482 VTAIL.n434 VSUBS 0.022956f
C483 VTAIL.n435 VSUBS 0.022956f
C484 VTAIL.n436 VSUBS 0.012336f
C485 VTAIL.n437 VSUBS 0.013061f
C486 VTAIL.n438 VSUBS 0.029157f
C487 VTAIL.n439 VSUBS 0.029157f
C488 VTAIL.n440 VSUBS 0.029157f
C489 VTAIL.n441 VSUBS 0.012699f
C490 VTAIL.n442 VSUBS 0.012336f
C491 VTAIL.n443 VSUBS 0.022956f
C492 VTAIL.n444 VSUBS 0.022956f
C493 VTAIL.n445 VSUBS 0.012336f
C494 VTAIL.n446 VSUBS 0.013061f
C495 VTAIL.n447 VSUBS 0.029157f
C496 VTAIL.n448 VSUBS 0.029157f
C497 VTAIL.n449 VSUBS 0.013061f
C498 VTAIL.n450 VSUBS 0.012336f
C499 VTAIL.n451 VSUBS 0.022956f
C500 VTAIL.n452 VSUBS 0.022956f
C501 VTAIL.n453 VSUBS 0.012336f
C502 VTAIL.n454 VSUBS 0.013061f
C503 VTAIL.n455 VSUBS 0.029157f
C504 VTAIL.n456 VSUBS 0.071917f
C505 VTAIL.n457 VSUBS 0.013061f
C506 VTAIL.n458 VSUBS 0.012336f
C507 VTAIL.n459 VSUBS 0.054631f
C508 VTAIL.n460 VSUBS 0.036273f
C509 VTAIL.n461 VSUBS 1.35325f
C510 VTAIL.n462 VSUBS 0.025615f
C511 VTAIL.n463 VSUBS 0.022956f
C512 VTAIL.n464 VSUBS 0.012336f
C513 VTAIL.n465 VSUBS 0.029157f
C514 VTAIL.n466 VSUBS 0.013061f
C515 VTAIL.n467 VSUBS 0.022956f
C516 VTAIL.n468 VSUBS 0.012336f
C517 VTAIL.n469 VSUBS 0.029157f
C518 VTAIL.n470 VSUBS 0.013061f
C519 VTAIL.n471 VSUBS 0.022956f
C520 VTAIL.n472 VSUBS 0.012699f
C521 VTAIL.n473 VSUBS 0.029157f
C522 VTAIL.n474 VSUBS 0.013061f
C523 VTAIL.n475 VSUBS 0.022956f
C524 VTAIL.n476 VSUBS 0.012336f
C525 VTAIL.n477 VSUBS 0.029157f
C526 VTAIL.n478 VSUBS 0.013061f
C527 VTAIL.n479 VSUBS 0.022956f
C528 VTAIL.n480 VSUBS 0.012336f
C529 VTAIL.n481 VSUBS 0.021868f
C530 VTAIL.n482 VSUBS 0.021934f
C531 VTAIL.t2 VSUBS 0.062845f
C532 VTAIL.n483 VSUBS 0.182561f
C533 VTAIL.n484 VSUBS 1.14502f
C534 VTAIL.n485 VSUBS 0.012336f
C535 VTAIL.n486 VSUBS 0.013061f
C536 VTAIL.n487 VSUBS 0.029157f
C537 VTAIL.n488 VSUBS 0.029157f
C538 VTAIL.n489 VSUBS 0.013061f
C539 VTAIL.n490 VSUBS 0.012336f
C540 VTAIL.n491 VSUBS 0.022956f
C541 VTAIL.n492 VSUBS 0.022956f
C542 VTAIL.n493 VSUBS 0.012336f
C543 VTAIL.n494 VSUBS 0.013061f
C544 VTAIL.n495 VSUBS 0.029157f
C545 VTAIL.n496 VSUBS 0.029157f
C546 VTAIL.n497 VSUBS 0.013061f
C547 VTAIL.n498 VSUBS 0.012336f
C548 VTAIL.n499 VSUBS 0.022956f
C549 VTAIL.n500 VSUBS 0.022956f
C550 VTAIL.n501 VSUBS 0.012336f
C551 VTAIL.n502 VSUBS 0.012336f
C552 VTAIL.n503 VSUBS 0.013061f
C553 VTAIL.n504 VSUBS 0.029157f
C554 VTAIL.n505 VSUBS 0.029157f
C555 VTAIL.n506 VSUBS 0.029157f
C556 VTAIL.n507 VSUBS 0.012699f
C557 VTAIL.n508 VSUBS 0.012336f
C558 VTAIL.n509 VSUBS 0.022956f
C559 VTAIL.n510 VSUBS 0.022956f
C560 VTAIL.n511 VSUBS 0.012336f
C561 VTAIL.n512 VSUBS 0.013061f
C562 VTAIL.n513 VSUBS 0.029157f
C563 VTAIL.n514 VSUBS 0.029157f
C564 VTAIL.n515 VSUBS 0.013061f
C565 VTAIL.n516 VSUBS 0.012336f
C566 VTAIL.n517 VSUBS 0.022956f
C567 VTAIL.n518 VSUBS 0.022956f
C568 VTAIL.n519 VSUBS 0.012336f
C569 VTAIL.n520 VSUBS 0.013061f
C570 VTAIL.n521 VSUBS 0.029157f
C571 VTAIL.n522 VSUBS 0.071917f
C572 VTAIL.n523 VSUBS 0.013061f
C573 VTAIL.n524 VSUBS 0.012336f
C574 VTAIL.n525 VSUBS 0.054631f
C575 VTAIL.n526 VSUBS 0.036273f
C576 VTAIL.n527 VSUBS 1.28773f
C577 VDD1.t3 VSUBS 0.257003f
C578 VDD1.t2 VSUBS 0.257003f
C579 VDD1.n0 VSUBS 2.01391f
C580 VDD1.t0 VSUBS 0.257003f
C581 VDD1.t1 VSUBS 0.257003f
C582 VDD1.n1 VSUBS 2.68753f
C583 VP.n0 VSUBS 0.043822f
C584 VP.t1 VSUBS 2.31133f
C585 VP.n1 VSUBS 0.063973f
C586 VP.t3 VSUBS 2.48413f
C587 VP.t2 VSUBS 2.48262f
C588 VP.n2 VSUBS 3.42789f
C589 VP.n3 VSUBS 2.4372f
C590 VP.t0 VSUBS 2.31133f
C591 VP.n4 VSUBS 0.929768f
C592 VP.n5 VSUBS 0.058286f
C593 VP.n6 VSUBS 0.043822f
C594 VP.n7 VSUBS 0.043822f
C595 VP.n8 VSUBS 0.043822f
C596 VP.n9 VSUBS 0.063973f
C597 VP.n10 VSUBS 0.058286f
C598 VP.n11 VSUBS 0.929768f
C599 VP.n12 VSUBS 0.042521f
C600 B.n0 VSUBS 0.004679f
C601 B.n1 VSUBS 0.004679f
C602 B.n2 VSUBS 0.007399f
C603 B.n3 VSUBS 0.007399f
C604 B.n4 VSUBS 0.007399f
C605 B.n5 VSUBS 0.007399f
C606 B.n6 VSUBS 0.007399f
C607 B.n7 VSUBS 0.007399f
C608 B.n8 VSUBS 0.007399f
C609 B.n9 VSUBS 0.007399f
C610 B.n10 VSUBS 0.007399f
C611 B.n11 VSUBS 0.007399f
C612 B.n12 VSUBS 0.007399f
C613 B.n13 VSUBS 0.007399f
C614 B.n14 VSUBS 0.016549f
C615 B.n15 VSUBS 0.007399f
C616 B.n16 VSUBS 0.007399f
C617 B.n17 VSUBS 0.007399f
C618 B.n18 VSUBS 0.007399f
C619 B.n19 VSUBS 0.007399f
C620 B.n20 VSUBS 0.007399f
C621 B.n21 VSUBS 0.007399f
C622 B.n22 VSUBS 0.007399f
C623 B.n23 VSUBS 0.007399f
C624 B.n24 VSUBS 0.007399f
C625 B.n25 VSUBS 0.007399f
C626 B.n26 VSUBS 0.007399f
C627 B.n27 VSUBS 0.007399f
C628 B.n28 VSUBS 0.007399f
C629 B.n29 VSUBS 0.007399f
C630 B.n30 VSUBS 0.007399f
C631 B.n31 VSUBS 0.007399f
C632 B.n32 VSUBS 0.007399f
C633 B.n33 VSUBS 0.007399f
C634 B.n34 VSUBS 0.007399f
C635 B.n35 VSUBS 0.007399f
C636 B.t8 VSUBS 0.227214f
C637 B.t7 VSUBS 0.249904f
C638 B.t6 VSUBS 0.897761f
C639 B.n36 VSUBS 0.382714f
C640 B.n37 VSUBS 0.264088f
C641 B.n38 VSUBS 0.007399f
C642 B.n39 VSUBS 0.007399f
C643 B.n40 VSUBS 0.007399f
C644 B.n41 VSUBS 0.007399f
C645 B.n42 VSUBS 0.004135f
C646 B.n43 VSUBS 0.007399f
C647 B.t11 VSUBS 0.227217f
C648 B.t10 VSUBS 0.249907f
C649 B.t9 VSUBS 0.897761f
C650 B.n44 VSUBS 0.382711f
C651 B.n45 VSUBS 0.264085f
C652 B.n46 VSUBS 0.017142f
C653 B.n47 VSUBS 0.007399f
C654 B.n48 VSUBS 0.007399f
C655 B.n49 VSUBS 0.007399f
C656 B.n50 VSUBS 0.007399f
C657 B.n51 VSUBS 0.007399f
C658 B.n52 VSUBS 0.007399f
C659 B.n53 VSUBS 0.007399f
C660 B.n54 VSUBS 0.007399f
C661 B.n55 VSUBS 0.007399f
C662 B.n56 VSUBS 0.007399f
C663 B.n57 VSUBS 0.007399f
C664 B.n58 VSUBS 0.007399f
C665 B.n59 VSUBS 0.007399f
C666 B.n60 VSUBS 0.007399f
C667 B.n61 VSUBS 0.007399f
C668 B.n62 VSUBS 0.007399f
C669 B.n63 VSUBS 0.007399f
C670 B.n64 VSUBS 0.007399f
C671 B.n65 VSUBS 0.007399f
C672 B.n66 VSUBS 0.017616f
C673 B.n67 VSUBS 0.007399f
C674 B.n68 VSUBS 0.007399f
C675 B.n69 VSUBS 0.007399f
C676 B.n70 VSUBS 0.007399f
C677 B.n71 VSUBS 0.007399f
C678 B.n72 VSUBS 0.007399f
C679 B.n73 VSUBS 0.007399f
C680 B.n74 VSUBS 0.007399f
C681 B.n75 VSUBS 0.007399f
C682 B.n76 VSUBS 0.007399f
C683 B.n77 VSUBS 0.007399f
C684 B.n78 VSUBS 0.007399f
C685 B.n79 VSUBS 0.007399f
C686 B.n80 VSUBS 0.007399f
C687 B.n81 VSUBS 0.007399f
C688 B.n82 VSUBS 0.007399f
C689 B.n83 VSUBS 0.007399f
C690 B.n84 VSUBS 0.007399f
C691 B.n85 VSUBS 0.007399f
C692 B.n86 VSUBS 0.007399f
C693 B.n87 VSUBS 0.007399f
C694 B.n88 VSUBS 0.007399f
C695 B.n89 VSUBS 0.007399f
C696 B.n90 VSUBS 0.007399f
C697 B.n91 VSUBS 0.007399f
C698 B.n92 VSUBS 0.017616f
C699 B.n93 VSUBS 0.007399f
C700 B.n94 VSUBS 0.007399f
C701 B.n95 VSUBS 0.007399f
C702 B.n96 VSUBS 0.007399f
C703 B.n97 VSUBS 0.007399f
C704 B.n98 VSUBS 0.007399f
C705 B.n99 VSUBS 0.007399f
C706 B.n100 VSUBS 0.007399f
C707 B.n101 VSUBS 0.007399f
C708 B.n102 VSUBS 0.007399f
C709 B.n103 VSUBS 0.007399f
C710 B.n104 VSUBS 0.007399f
C711 B.n105 VSUBS 0.007399f
C712 B.n106 VSUBS 0.007399f
C713 B.n107 VSUBS 0.007399f
C714 B.n108 VSUBS 0.007399f
C715 B.n109 VSUBS 0.007399f
C716 B.n110 VSUBS 0.007399f
C717 B.n111 VSUBS 0.007399f
C718 B.n112 VSUBS 0.007399f
C719 B.t1 VSUBS 0.227217f
C720 B.t2 VSUBS 0.249907f
C721 B.t0 VSUBS 0.897761f
C722 B.n113 VSUBS 0.382711f
C723 B.n114 VSUBS 0.264085f
C724 B.n115 VSUBS 0.017142f
C725 B.n116 VSUBS 0.007399f
C726 B.n117 VSUBS 0.007399f
C727 B.n118 VSUBS 0.007399f
C728 B.n119 VSUBS 0.007399f
C729 B.n120 VSUBS 0.007399f
C730 B.t4 VSUBS 0.227214f
C731 B.t5 VSUBS 0.249904f
C732 B.t3 VSUBS 0.897761f
C733 B.n121 VSUBS 0.382714f
C734 B.n122 VSUBS 0.264088f
C735 B.n123 VSUBS 0.007399f
C736 B.n124 VSUBS 0.007399f
C737 B.n125 VSUBS 0.007399f
C738 B.n126 VSUBS 0.007399f
C739 B.n127 VSUBS 0.007399f
C740 B.n128 VSUBS 0.007399f
C741 B.n129 VSUBS 0.007399f
C742 B.n130 VSUBS 0.007399f
C743 B.n131 VSUBS 0.007399f
C744 B.n132 VSUBS 0.007399f
C745 B.n133 VSUBS 0.007399f
C746 B.n134 VSUBS 0.007399f
C747 B.n135 VSUBS 0.007399f
C748 B.n136 VSUBS 0.007399f
C749 B.n137 VSUBS 0.007399f
C750 B.n138 VSUBS 0.007399f
C751 B.n139 VSUBS 0.007399f
C752 B.n140 VSUBS 0.007399f
C753 B.n141 VSUBS 0.007399f
C754 B.n142 VSUBS 0.007399f
C755 B.n143 VSUBS 0.017616f
C756 B.n144 VSUBS 0.007399f
C757 B.n145 VSUBS 0.007399f
C758 B.n146 VSUBS 0.007399f
C759 B.n147 VSUBS 0.007399f
C760 B.n148 VSUBS 0.007399f
C761 B.n149 VSUBS 0.007399f
C762 B.n150 VSUBS 0.007399f
C763 B.n151 VSUBS 0.007399f
C764 B.n152 VSUBS 0.007399f
C765 B.n153 VSUBS 0.007399f
C766 B.n154 VSUBS 0.007399f
C767 B.n155 VSUBS 0.007399f
C768 B.n156 VSUBS 0.007399f
C769 B.n157 VSUBS 0.007399f
C770 B.n158 VSUBS 0.007399f
C771 B.n159 VSUBS 0.007399f
C772 B.n160 VSUBS 0.007399f
C773 B.n161 VSUBS 0.007399f
C774 B.n162 VSUBS 0.007399f
C775 B.n163 VSUBS 0.007399f
C776 B.n164 VSUBS 0.007399f
C777 B.n165 VSUBS 0.007399f
C778 B.n166 VSUBS 0.007399f
C779 B.n167 VSUBS 0.007399f
C780 B.n168 VSUBS 0.007399f
C781 B.n169 VSUBS 0.007399f
C782 B.n170 VSUBS 0.007399f
C783 B.n171 VSUBS 0.007399f
C784 B.n172 VSUBS 0.007399f
C785 B.n173 VSUBS 0.007399f
C786 B.n174 VSUBS 0.007399f
C787 B.n175 VSUBS 0.007399f
C788 B.n176 VSUBS 0.007399f
C789 B.n177 VSUBS 0.007399f
C790 B.n178 VSUBS 0.007399f
C791 B.n179 VSUBS 0.007399f
C792 B.n180 VSUBS 0.007399f
C793 B.n181 VSUBS 0.007399f
C794 B.n182 VSUBS 0.007399f
C795 B.n183 VSUBS 0.007399f
C796 B.n184 VSUBS 0.007399f
C797 B.n185 VSUBS 0.007399f
C798 B.n186 VSUBS 0.007399f
C799 B.n187 VSUBS 0.007399f
C800 B.n188 VSUBS 0.007399f
C801 B.n189 VSUBS 0.007399f
C802 B.n190 VSUBS 0.016549f
C803 B.n191 VSUBS 0.016549f
C804 B.n192 VSUBS 0.017616f
C805 B.n193 VSUBS 0.007399f
C806 B.n194 VSUBS 0.007399f
C807 B.n195 VSUBS 0.007399f
C808 B.n196 VSUBS 0.007399f
C809 B.n197 VSUBS 0.007399f
C810 B.n198 VSUBS 0.007399f
C811 B.n199 VSUBS 0.007399f
C812 B.n200 VSUBS 0.007399f
C813 B.n201 VSUBS 0.007399f
C814 B.n202 VSUBS 0.007399f
C815 B.n203 VSUBS 0.007399f
C816 B.n204 VSUBS 0.007399f
C817 B.n205 VSUBS 0.007399f
C818 B.n206 VSUBS 0.007399f
C819 B.n207 VSUBS 0.007399f
C820 B.n208 VSUBS 0.007399f
C821 B.n209 VSUBS 0.007399f
C822 B.n210 VSUBS 0.007399f
C823 B.n211 VSUBS 0.007399f
C824 B.n212 VSUBS 0.007399f
C825 B.n213 VSUBS 0.007399f
C826 B.n214 VSUBS 0.007399f
C827 B.n215 VSUBS 0.007399f
C828 B.n216 VSUBS 0.007399f
C829 B.n217 VSUBS 0.007399f
C830 B.n218 VSUBS 0.007399f
C831 B.n219 VSUBS 0.007399f
C832 B.n220 VSUBS 0.007399f
C833 B.n221 VSUBS 0.007399f
C834 B.n222 VSUBS 0.007399f
C835 B.n223 VSUBS 0.007399f
C836 B.n224 VSUBS 0.007399f
C837 B.n225 VSUBS 0.007399f
C838 B.n226 VSUBS 0.007399f
C839 B.n227 VSUBS 0.007399f
C840 B.n228 VSUBS 0.007399f
C841 B.n229 VSUBS 0.007399f
C842 B.n230 VSUBS 0.007399f
C843 B.n231 VSUBS 0.007399f
C844 B.n232 VSUBS 0.007399f
C845 B.n233 VSUBS 0.007399f
C846 B.n234 VSUBS 0.007399f
C847 B.n235 VSUBS 0.007399f
C848 B.n236 VSUBS 0.007399f
C849 B.n237 VSUBS 0.007399f
C850 B.n238 VSUBS 0.007399f
C851 B.n239 VSUBS 0.007399f
C852 B.n240 VSUBS 0.007399f
C853 B.n241 VSUBS 0.007399f
C854 B.n242 VSUBS 0.007399f
C855 B.n243 VSUBS 0.007399f
C856 B.n244 VSUBS 0.007399f
C857 B.n245 VSUBS 0.007399f
C858 B.n246 VSUBS 0.007399f
C859 B.n247 VSUBS 0.007399f
C860 B.n248 VSUBS 0.007399f
C861 B.n249 VSUBS 0.007399f
C862 B.n250 VSUBS 0.007399f
C863 B.n251 VSUBS 0.007399f
C864 B.n252 VSUBS 0.007399f
C865 B.n253 VSUBS 0.007399f
C866 B.n254 VSUBS 0.006964f
C867 B.n255 VSUBS 0.017142f
C868 B.n256 VSUBS 0.004135f
C869 B.n257 VSUBS 0.007399f
C870 B.n258 VSUBS 0.007399f
C871 B.n259 VSUBS 0.007399f
C872 B.n260 VSUBS 0.007399f
C873 B.n261 VSUBS 0.007399f
C874 B.n262 VSUBS 0.007399f
C875 B.n263 VSUBS 0.007399f
C876 B.n264 VSUBS 0.007399f
C877 B.n265 VSUBS 0.007399f
C878 B.n266 VSUBS 0.007399f
C879 B.n267 VSUBS 0.007399f
C880 B.n268 VSUBS 0.007399f
C881 B.n269 VSUBS 0.004135f
C882 B.n270 VSUBS 0.007399f
C883 B.n271 VSUBS 0.007399f
C884 B.n272 VSUBS 0.006964f
C885 B.n273 VSUBS 0.007399f
C886 B.n274 VSUBS 0.007399f
C887 B.n275 VSUBS 0.007399f
C888 B.n276 VSUBS 0.007399f
C889 B.n277 VSUBS 0.007399f
C890 B.n278 VSUBS 0.007399f
C891 B.n279 VSUBS 0.007399f
C892 B.n280 VSUBS 0.007399f
C893 B.n281 VSUBS 0.007399f
C894 B.n282 VSUBS 0.007399f
C895 B.n283 VSUBS 0.007399f
C896 B.n284 VSUBS 0.007399f
C897 B.n285 VSUBS 0.007399f
C898 B.n286 VSUBS 0.007399f
C899 B.n287 VSUBS 0.007399f
C900 B.n288 VSUBS 0.007399f
C901 B.n289 VSUBS 0.007399f
C902 B.n290 VSUBS 0.007399f
C903 B.n291 VSUBS 0.007399f
C904 B.n292 VSUBS 0.007399f
C905 B.n293 VSUBS 0.007399f
C906 B.n294 VSUBS 0.007399f
C907 B.n295 VSUBS 0.007399f
C908 B.n296 VSUBS 0.007399f
C909 B.n297 VSUBS 0.007399f
C910 B.n298 VSUBS 0.007399f
C911 B.n299 VSUBS 0.007399f
C912 B.n300 VSUBS 0.007399f
C913 B.n301 VSUBS 0.007399f
C914 B.n302 VSUBS 0.007399f
C915 B.n303 VSUBS 0.007399f
C916 B.n304 VSUBS 0.007399f
C917 B.n305 VSUBS 0.007399f
C918 B.n306 VSUBS 0.007399f
C919 B.n307 VSUBS 0.007399f
C920 B.n308 VSUBS 0.007399f
C921 B.n309 VSUBS 0.007399f
C922 B.n310 VSUBS 0.007399f
C923 B.n311 VSUBS 0.007399f
C924 B.n312 VSUBS 0.007399f
C925 B.n313 VSUBS 0.007399f
C926 B.n314 VSUBS 0.007399f
C927 B.n315 VSUBS 0.007399f
C928 B.n316 VSUBS 0.007399f
C929 B.n317 VSUBS 0.007399f
C930 B.n318 VSUBS 0.007399f
C931 B.n319 VSUBS 0.007399f
C932 B.n320 VSUBS 0.007399f
C933 B.n321 VSUBS 0.007399f
C934 B.n322 VSUBS 0.007399f
C935 B.n323 VSUBS 0.007399f
C936 B.n324 VSUBS 0.007399f
C937 B.n325 VSUBS 0.007399f
C938 B.n326 VSUBS 0.007399f
C939 B.n327 VSUBS 0.007399f
C940 B.n328 VSUBS 0.007399f
C941 B.n329 VSUBS 0.007399f
C942 B.n330 VSUBS 0.007399f
C943 B.n331 VSUBS 0.007399f
C944 B.n332 VSUBS 0.007399f
C945 B.n333 VSUBS 0.017616f
C946 B.n334 VSUBS 0.016549f
C947 B.n335 VSUBS 0.016549f
C948 B.n336 VSUBS 0.007399f
C949 B.n337 VSUBS 0.007399f
C950 B.n338 VSUBS 0.007399f
C951 B.n339 VSUBS 0.007399f
C952 B.n340 VSUBS 0.007399f
C953 B.n341 VSUBS 0.007399f
C954 B.n342 VSUBS 0.007399f
C955 B.n343 VSUBS 0.007399f
C956 B.n344 VSUBS 0.007399f
C957 B.n345 VSUBS 0.007399f
C958 B.n346 VSUBS 0.007399f
C959 B.n347 VSUBS 0.007399f
C960 B.n348 VSUBS 0.007399f
C961 B.n349 VSUBS 0.007399f
C962 B.n350 VSUBS 0.007399f
C963 B.n351 VSUBS 0.007399f
C964 B.n352 VSUBS 0.007399f
C965 B.n353 VSUBS 0.007399f
C966 B.n354 VSUBS 0.007399f
C967 B.n355 VSUBS 0.007399f
C968 B.n356 VSUBS 0.007399f
C969 B.n357 VSUBS 0.007399f
C970 B.n358 VSUBS 0.007399f
C971 B.n359 VSUBS 0.007399f
C972 B.n360 VSUBS 0.007399f
C973 B.n361 VSUBS 0.007399f
C974 B.n362 VSUBS 0.007399f
C975 B.n363 VSUBS 0.007399f
C976 B.n364 VSUBS 0.007399f
C977 B.n365 VSUBS 0.007399f
C978 B.n366 VSUBS 0.007399f
C979 B.n367 VSUBS 0.007399f
C980 B.n368 VSUBS 0.007399f
C981 B.n369 VSUBS 0.007399f
C982 B.n370 VSUBS 0.007399f
C983 B.n371 VSUBS 0.007399f
C984 B.n372 VSUBS 0.007399f
C985 B.n373 VSUBS 0.007399f
C986 B.n374 VSUBS 0.007399f
C987 B.n375 VSUBS 0.007399f
C988 B.n376 VSUBS 0.007399f
C989 B.n377 VSUBS 0.007399f
C990 B.n378 VSUBS 0.007399f
C991 B.n379 VSUBS 0.007399f
C992 B.n380 VSUBS 0.007399f
C993 B.n381 VSUBS 0.007399f
C994 B.n382 VSUBS 0.007399f
C995 B.n383 VSUBS 0.007399f
C996 B.n384 VSUBS 0.007399f
C997 B.n385 VSUBS 0.007399f
C998 B.n386 VSUBS 0.007399f
C999 B.n387 VSUBS 0.007399f
C1000 B.n388 VSUBS 0.007399f
C1001 B.n389 VSUBS 0.007399f
C1002 B.n390 VSUBS 0.007399f
C1003 B.n391 VSUBS 0.007399f
C1004 B.n392 VSUBS 0.007399f
C1005 B.n393 VSUBS 0.007399f
C1006 B.n394 VSUBS 0.007399f
C1007 B.n395 VSUBS 0.007399f
C1008 B.n396 VSUBS 0.007399f
C1009 B.n397 VSUBS 0.007399f
C1010 B.n398 VSUBS 0.007399f
C1011 B.n399 VSUBS 0.007399f
C1012 B.n400 VSUBS 0.007399f
C1013 B.n401 VSUBS 0.007399f
C1014 B.n402 VSUBS 0.007399f
C1015 B.n403 VSUBS 0.007399f
C1016 B.n404 VSUBS 0.007399f
C1017 B.n405 VSUBS 0.007399f
C1018 B.n406 VSUBS 0.007399f
C1019 B.n407 VSUBS 0.007399f
C1020 B.n408 VSUBS 0.007399f
C1021 B.n409 VSUBS 0.016549f
C1022 B.n410 VSUBS 0.017442f
C1023 B.n411 VSUBS 0.016723f
C1024 B.n412 VSUBS 0.007399f
C1025 B.n413 VSUBS 0.007399f
C1026 B.n414 VSUBS 0.007399f
C1027 B.n415 VSUBS 0.007399f
C1028 B.n416 VSUBS 0.007399f
C1029 B.n417 VSUBS 0.007399f
C1030 B.n418 VSUBS 0.007399f
C1031 B.n419 VSUBS 0.007399f
C1032 B.n420 VSUBS 0.007399f
C1033 B.n421 VSUBS 0.007399f
C1034 B.n422 VSUBS 0.007399f
C1035 B.n423 VSUBS 0.007399f
C1036 B.n424 VSUBS 0.007399f
C1037 B.n425 VSUBS 0.007399f
C1038 B.n426 VSUBS 0.007399f
C1039 B.n427 VSUBS 0.007399f
C1040 B.n428 VSUBS 0.007399f
C1041 B.n429 VSUBS 0.007399f
C1042 B.n430 VSUBS 0.007399f
C1043 B.n431 VSUBS 0.007399f
C1044 B.n432 VSUBS 0.007399f
C1045 B.n433 VSUBS 0.007399f
C1046 B.n434 VSUBS 0.007399f
C1047 B.n435 VSUBS 0.007399f
C1048 B.n436 VSUBS 0.007399f
C1049 B.n437 VSUBS 0.007399f
C1050 B.n438 VSUBS 0.007399f
C1051 B.n439 VSUBS 0.007399f
C1052 B.n440 VSUBS 0.007399f
C1053 B.n441 VSUBS 0.007399f
C1054 B.n442 VSUBS 0.007399f
C1055 B.n443 VSUBS 0.007399f
C1056 B.n444 VSUBS 0.007399f
C1057 B.n445 VSUBS 0.007399f
C1058 B.n446 VSUBS 0.007399f
C1059 B.n447 VSUBS 0.007399f
C1060 B.n448 VSUBS 0.007399f
C1061 B.n449 VSUBS 0.007399f
C1062 B.n450 VSUBS 0.007399f
C1063 B.n451 VSUBS 0.007399f
C1064 B.n452 VSUBS 0.007399f
C1065 B.n453 VSUBS 0.007399f
C1066 B.n454 VSUBS 0.007399f
C1067 B.n455 VSUBS 0.007399f
C1068 B.n456 VSUBS 0.007399f
C1069 B.n457 VSUBS 0.007399f
C1070 B.n458 VSUBS 0.007399f
C1071 B.n459 VSUBS 0.007399f
C1072 B.n460 VSUBS 0.007399f
C1073 B.n461 VSUBS 0.007399f
C1074 B.n462 VSUBS 0.007399f
C1075 B.n463 VSUBS 0.007399f
C1076 B.n464 VSUBS 0.007399f
C1077 B.n465 VSUBS 0.007399f
C1078 B.n466 VSUBS 0.007399f
C1079 B.n467 VSUBS 0.007399f
C1080 B.n468 VSUBS 0.007399f
C1081 B.n469 VSUBS 0.007399f
C1082 B.n470 VSUBS 0.007399f
C1083 B.n471 VSUBS 0.007399f
C1084 B.n472 VSUBS 0.006964f
C1085 B.n473 VSUBS 0.007399f
C1086 B.n474 VSUBS 0.007399f
C1087 B.n475 VSUBS 0.007399f
C1088 B.n476 VSUBS 0.007399f
C1089 B.n477 VSUBS 0.007399f
C1090 B.n478 VSUBS 0.007399f
C1091 B.n479 VSUBS 0.007399f
C1092 B.n480 VSUBS 0.007399f
C1093 B.n481 VSUBS 0.007399f
C1094 B.n482 VSUBS 0.007399f
C1095 B.n483 VSUBS 0.007399f
C1096 B.n484 VSUBS 0.007399f
C1097 B.n485 VSUBS 0.007399f
C1098 B.n486 VSUBS 0.007399f
C1099 B.n487 VSUBS 0.007399f
C1100 B.n488 VSUBS 0.004135f
C1101 B.n489 VSUBS 0.017142f
C1102 B.n490 VSUBS 0.006964f
C1103 B.n491 VSUBS 0.007399f
C1104 B.n492 VSUBS 0.007399f
C1105 B.n493 VSUBS 0.007399f
C1106 B.n494 VSUBS 0.007399f
C1107 B.n495 VSUBS 0.007399f
C1108 B.n496 VSUBS 0.007399f
C1109 B.n497 VSUBS 0.007399f
C1110 B.n498 VSUBS 0.007399f
C1111 B.n499 VSUBS 0.007399f
C1112 B.n500 VSUBS 0.007399f
C1113 B.n501 VSUBS 0.007399f
C1114 B.n502 VSUBS 0.007399f
C1115 B.n503 VSUBS 0.007399f
C1116 B.n504 VSUBS 0.007399f
C1117 B.n505 VSUBS 0.007399f
C1118 B.n506 VSUBS 0.007399f
C1119 B.n507 VSUBS 0.007399f
C1120 B.n508 VSUBS 0.007399f
C1121 B.n509 VSUBS 0.007399f
C1122 B.n510 VSUBS 0.007399f
C1123 B.n511 VSUBS 0.007399f
C1124 B.n512 VSUBS 0.007399f
C1125 B.n513 VSUBS 0.007399f
C1126 B.n514 VSUBS 0.007399f
C1127 B.n515 VSUBS 0.007399f
C1128 B.n516 VSUBS 0.007399f
C1129 B.n517 VSUBS 0.007399f
C1130 B.n518 VSUBS 0.007399f
C1131 B.n519 VSUBS 0.007399f
C1132 B.n520 VSUBS 0.007399f
C1133 B.n521 VSUBS 0.007399f
C1134 B.n522 VSUBS 0.007399f
C1135 B.n523 VSUBS 0.007399f
C1136 B.n524 VSUBS 0.007399f
C1137 B.n525 VSUBS 0.007399f
C1138 B.n526 VSUBS 0.007399f
C1139 B.n527 VSUBS 0.007399f
C1140 B.n528 VSUBS 0.007399f
C1141 B.n529 VSUBS 0.007399f
C1142 B.n530 VSUBS 0.007399f
C1143 B.n531 VSUBS 0.007399f
C1144 B.n532 VSUBS 0.007399f
C1145 B.n533 VSUBS 0.007399f
C1146 B.n534 VSUBS 0.007399f
C1147 B.n535 VSUBS 0.007399f
C1148 B.n536 VSUBS 0.007399f
C1149 B.n537 VSUBS 0.007399f
C1150 B.n538 VSUBS 0.007399f
C1151 B.n539 VSUBS 0.007399f
C1152 B.n540 VSUBS 0.007399f
C1153 B.n541 VSUBS 0.007399f
C1154 B.n542 VSUBS 0.007399f
C1155 B.n543 VSUBS 0.007399f
C1156 B.n544 VSUBS 0.007399f
C1157 B.n545 VSUBS 0.007399f
C1158 B.n546 VSUBS 0.007399f
C1159 B.n547 VSUBS 0.007399f
C1160 B.n548 VSUBS 0.007399f
C1161 B.n549 VSUBS 0.007399f
C1162 B.n550 VSUBS 0.007399f
C1163 B.n551 VSUBS 0.017616f
C1164 B.n552 VSUBS 0.017616f
C1165 B.n553 VSUBS 0.016549f
C1166 B.n554 VSUBS 0.007399f
C1167 B.n555 VSUBS 0.007399f
C1168 B.n556 VSUBS 0.007399f
C1169 B.n557 VSUBS 0.007399f
C1170 B.n558 VSUBS 0.007399f
C1171 B.n559 VSUBS 0.007399f
C1172 B.n560 VSUBS 0.007399f
C1173 B.n561 VSUBS 0.007399f
C1174 B.n562 VSUBS 0.007399f
C1175 B.n563 VSUBS 0.007399f
C1176 B.n564 VSUBS 0.007399f
C1177 B.n565 VSUBS 0.007399f
C1178 B.n566 VSUBS 0.007399f
C1179 B.n567 VSUBS 0.007399f
C1180 B.n568 VSUBS 0.007399f
C1181 B.n569 VSUBS 0.007399f
C1182 B.n570 VSUBS 0.007399f
C1183 B.n571 VSUBS 0.007399f
C1184 B.n572 VSUBS 0.007399f
C1185 B.n573 VSUBS 0.007399f
C1186 B.n574 VSUBS 0.007399f
C1187 B.n575 VSUBS 0.007399f
C1188 B.n576 VSUBS 0.007399f
C1189 B.n577 VSUBS 0.007399f
C1190 B.n578 VSUBS 0.007399f
C1191 B.n579 VSUBS 0.007399f
C1192 B.n580 VSUBS 0.007399f
C1193 B.n581 VSUBS 0.007399f
C1194 B.n582 VSUBS 0.007399f
C1195 B.n583 VSUBS 0.007399f
C1196 B.n584 VSUBS 0.007399f
C1197 B.n585 VSUBS 0.007399f
C1198 B.n586 VSUBS 0.007399f
C1199 B.n587 VSUBS 0.007399f
C1200 B.n588 VSUBS 0.007399f
C1201 B.n589 VSUBS 0.007399f
C1202 B.n590 VSUBS 0.007399f
C1203 B.n591 VSUBS 0.016753f
.ends

