* NGSPICE file created from diff_pair_sample_0459.ext - technology: sky130A

.subckt diff_pair_sample_0459 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=1.46
X1 VDD2.t5 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=1.46
X2 VTAIL.t9 VN.t2 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=1.46
X3 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=1.46
X4 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=1.46
X5 VDD2.t3 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=1.46
X6 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=1.46
X7 VTAIL.t0 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=1.46
X8 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=1.46
X9 VDD2.t2 VN.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=1.46
X10 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=1.46
X11 VDD2.t0 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=1.46
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=1.46
X13 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=1.46
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=1.46
X15 VDD1.t0 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=1.46
R0 VN.n9 VN.n8 171.524
R1 VN.n19 VN.n18 171.524
R2 VN.n17 VN.n10 161.3
R3 VN.n16 VN.n15 161.3
R4 VN.n14 VN.n11 161.3
R5 VN.n7 VN.n0 161.3
R6 VN.n6 VN.n5 161.3
R7 VN.n4 VN.n1 161.3
R8 VN.n3 VN.t1 66.583
R9 VN.n13 VN.t5 66.583
R10 VN.n6 VN.n1 50.6348
R11 VN.n16 VN.n11 50.6348
R12 VN.n3 VN.n2 41.7711
R13 VN.n13 VN.n12 41.7711
R14 VN VN.n19 36.8547
R15 VN.n7 VN.n6 30.1864
R16 VN.n17 VN.n16 30.1864
R17 VN.n2 VN.t0 30.043
R18 VN.n8 VN.t4 30.043
R19 VN.n12 VN.t2 30.043
R20 VN.n18 VN.t3 30.043
R21 VN.n2 VN.n1 24.3439
R22 VN.n12 VN.n11 24.3439
R23 VN.n14 VN.n13 17.3537
R24 VN.n4 VN.n3 17.3537
R25 VN.n8 VN.n7 14.1197
R26 VN.n18 VN.n17 14.1197
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n11 VDD2.n9 289.615
R35 VDD2.n2 VDD2.n0 289.615
R36 VDD2.n12 VDD2.n11 185
R37 VDD2.n3 VDD2.n2 185
R38 VDD2.t3 VDD2.n10 164.876
R39 VDD2.t5 VDD2.n1 164.876
R40 VDD2.n8 VDD2.n7 102.529
R41 VDD2 VDD2.n17 102.526
R42 VDD2.n8 VDD2.n6 52.6813
R43 VDD2.n11 VDD2.t3 52.3082
R44 VDD2.n2 VDD2.t5 52.3082
R45 VDD2.n16 VDD2.n15 51.5793
R46 VDD2.n16 VDD2.n8 30.2993
R47 VDD2.n12 VDD2.n10 14.7318
R48 VDD2.n3 VDD2.n1 14.7318
R49 VDD2.n13 VDD2.n9 12.8005
R50 VDD2.n4 VDD2.n0 12.8005
R51 VDD2.n17 VDD2.t4 10.8796
R52 VDD2.n17 VDD2.t0 10.8796
R53 VDD2.n7 VDD2.t1 10.8796
R54 VDD2.n7 VDD2.t2 10.8796
R55 VDD2.n15 VDD2.n14 9.45567
R56 VDD2.n6 VDD2.n5 9.45567
R57 VDD2.n14 VDD2.n13 9.3005
R58 VDD2.n5 VDD2.n4 9.3005
R59 VDD2.n14 VDD2.n10 5.62509
R60 VDD2.n5 VDD2.n1 5.62509
R61 VDD2 VDD2.n16 1.21602
R62 VDD2.n15 VDD2.n9 1.16414
R63 VDD2.n6 VDD2.n0 1.16414
R64 VDD2.n13 VDD2.n12 0.388379
R65 VDD2.n4 VDD2.n3 0.388379
R66 VTAIL.n34 VTAIL.n32 289.615
R67 VTAIL.n4 VTAIL.n2 289.615
R68 VTAIL.n26 VTAIL.n24 289.615
R69 VTAIL.n16 VTAIL.n14 289.615
R70 VTAIL.n35 VTAIL.n34 185
R71 VTAIL.n5 VTAIL.n4 185
R72 VTAIL.n27 VTAIL.n26 185
R73 VTAIL.n17 VTAIL.n16 185
R74 VTAIL.t7 VTAIL.n33 164.876
R75 VTAIL.t3 VTAIL.n3 164.876
R76 VTAIL.t4 VTAIL.n25 164.876
R77 VTAIL.t6 VTAIL.n15 164.876
R78 VTAIL.n23 VTAIL.n22 85.5201
R79 VTAIL.n13 VTAIL.n12 85.5201
R80 VTAIL.n1 VTAIL.n0 85.52
R81 VTAIL.n11 VTAIL.n10 85.52
R82 VTAIL.n34 VTAIL.t7 52.3082
R83 VTAIL.n4 VTAIL.t3 52.3082
R84 VTAIL.n26 VTAIL.t4 52.3082
R85 VTAIL.n16 VTAIL.t6 52.3082
R86 VTAIL.n39 VTAIL.n38 34.9005
R87 VTAIL.n9 VTAIL.n8 34.9005
R88 VTAIL.n31 VTAIL.n30 34.9005
R89 VTAIL.n21 VTAIL.n20 34.9005
R90 VTAIL.n13 VTAIL.n11 17.0221
R91 VTAIL.n39 VTAIL.n31 15.4789
R92 VTAIL.n35 VTAIL.n33 14.7318
R93 VTAIL.n5 VTAIL.n3 14.7318
R94 VTAIL.n27 VTAIL.n25 14.7318
R95 VTAIL.n17 VTAIL.n15 14.7318
R96 VTAIL.n36 VTAIL.n32 12.8005
R97 VTAIL.n6 VTAIL.n2 12.8005
R98 VTAIL.n28 VTAIL.n24 12.8005
R99 VTAIL.n18 VTAIL.n14 12.8005
R100 VTAIL.n0 VTAIL.t10 10.8796
R101 VTAIL.n0 VTAIL.t11 10.8796
R102 VTAIL.n10 VTAIL.t2 10.8796
R103 VTAIL.n10 VTAIL.t1 10.8796
R104 VTAIL.n22 VTAIL.t5 10.8796
R105 VTAIL.n22 VTAIL.t0 10.8796
R106 VTAIL.n12 VTAIL.t8 10.8796
R107 VTAIL.n12 VTAIL.t9 10.8796
R108 VTAIL.n38 VTAIL.n37 9.45567
R109 VTAIL.n8 VTAIL.n7 9.45567
R110 VTAIL.n30 VTAIL.n29 9.45567
R111 VTAIL.n20 VTAIL.n19 9.45567
R112 VTAIL.n37 VTAIL.n36 9.3005
R113 VTAIL.n7 VTAIL.n6 9.3005
R114 VTAIL.n29 VTAIL.n28 9.3005
R115 VTAIL.n19 VTAIL.n18 9.3005
R116 VTAIL.n37 VTAIL.n33 5.62509
R117 VTAIL.n7 VTAIL.n3 5.62509
R118 VTAIL.n29 VTAIL.n25 5.62509
R119 VTAIL.n19 VTAIL.n15 5.62509
R120 VTAIL.n21 VTAIL.n13 1.5436
R121 VTAIL.n31 VTAIL.n23 1.5436
R122 VTAIL.n11 VTAIL.n9 1.5436
R123 VTAIL.n23 VTAIL.n21 1.24188
R124 VTAIL.n9 VTAIL.n1 1.24188
R125 VTAIL.n38 VTAIL.n32 1.16414
R126 VTAIL.n8 VTAIL.n2 1.16414
R127 VTAIL.n30 VTAIL.n24 1.16414
R128 VTAIL.n20 VTAIL.n14 1.16414
R129 VTAIL VTAIL.n39 1.09964
R130 VTAIL VTAIL.n1 0.444466
R131 VTAIL.n36 VTAIL.n35 0.388379
R132 VTAIL.n6 VTAIL.n5 0.388379
R133 VTAIL.n28 VTAIL.n27 0.388379
R134 VTAIL.n18 VTAIL.n17 0.388379
R135 B.n411 B.n410 585
R136 B.n412 B.n411 585
R137 B.n141 B.n72 585
R138 B.n140 B.n139 585
R139 B.n138 B.n137 585
R140 B.n136 B.n135 585
R141 B.n134 B.n133 585
R142 B.n132 B.n131 585
R143 B.n130 B.n129 585
R144 B.n128 B.n127 585
R145 B.n126 B.n125 585
R146 B.n124 B.n123 585
R147 B.n122 B.n121 585
R148 B.n119 B.n118 585
R149 B.n117 B.n116 585
R150 B.n115 B.n114 585
R151 B.n113 B.n112 585
R152 B.n111 B.n110 585
R153 B.n109 B.n108 585
R154 B.n107 B.n106 585
R155 B.n105 B.n104 585
R156 B.n103 B.n102 585
R157 B.n101 B.n100 585
R158 B.n99 B.n98 585
R159 B.n97 B.n96 585
R160 B.n95 B.n94 585
R161 B.n93 B.n92 585
R162 B.n91 B.n90 585
R163 B.n89 B.n88 585
R164 B.n87 B.n86 585
R165 B.n85 B.n84 585
R166 B.n83 B.n82 585
R167 B.n81 B.n80 585
R168 B.n79 B.n78 585
R169 B.n409 B.n55 585
R170 B.n413 B.n55 585
R171 B.n408 B.n54 585
R172 B.n414 B.n54 585
R173 B.n407 B.n406 585
R174 B.n406 B.n50 585
R175 B.n405 B.n49 585
R176 B.n420 B.n49 585
R177 B.n404 B.n48 585
R178 B.n421 B.n48 585
R179 B.n403 B.n47 585
R180 B.n422 B.n47 585
R181 B.n402 B.n401 585
R182 B.n401 B.n43 585
R183 B.n400 B.n42 585
R184 B.n428 B.n42 585
R185 B.n399 B.n41 585
R186 B.n429 B.n41 585
R187 B.n398 B.n40 585
R188 B.n430 B.n40 585
R189 B.n397 B.n396 585
R190 B.n396 B.n36 585
R191 B.n395 B.n35 585
R192 B.n436 B.n35 585
R193 B.n394 B.n34 585
R194 B.n437 B.n34 585
R195 B.n393 B.n33 585
R196 B.n438 B.n33 585
R197 B.n392 B.n391 585
R198 B.n391 B.n32 585
R199 B.n390 B.n28 585
R200 B.n444 B.n28 585
R201 B.n389 B.n27 585
R202 B.n445 B.n27 585
R203 B.n388 B.n26 585
R204 B.n446 B.n26 585
R205 B.n387 B.n386 585
R206 B.n386 B.n22 585
R207 B.n385 B.n21 585
R208 B.n452 B.n21 585
R209 B.n384 B.n20 585
R210 B.n453 B.n20 585
R211 B.n383 B.n19 585
R212 B.n454 B.n19 585
R213 B.n382 B.n381 585
R214 B.n381 B.n15 585
R215 B.n380 B.n14 585
R216 B.n460 B.n14 585
R217 B.n379 B.n13 585
R218 B.n461 B.n13 585
R219 B.n378 B.n12 585
R220 B.n462 B.n12 585
R221 B.n377 B.n376 585
R222 B.n376 B.n8 585
R223 B.n375 B.n7 585
R224 B.n468 B.n7 585
R225 B.n374 B.n6 585
R226 B.n469 B.n6 585
R227 B.n373 B.n5 585
R228 B.n470 B.n5 585
R229 B.n372 B.n371 585
R230 B.n371 B.n4 585
R231 B.n370 B.n142 585
R232 B.n370 B.n369 585
R233 B.n360 B.n143 585
R234 B.n144 B.n143 585
R235 B.n362 B.n361 585
R236 B.n363 B.n362 585
R237 B.n359 B.n148 585
R238 B.n152 B.n148 585
R239 B.n358 B.n357 585
R240 B.n357 B.n356 585
R241 B.n150 B.n149 585
R242 B.n151 B.n150 585
R243 B.n349 B.n348 585
R244 B.n350 B.n349 585
R245 B.n347 B.n157 585
R246 B.n157 B.n156 585
R247 B.n346 B.n345 585
R248 B.n345 B.n344 585
R249 B.n159 B.n158 585
R250 B.n160 B.n159 585
R251 B.n337 B.n336 585
R252 B.n338 B.n337 585
R253 B.n335 B.n165 585
R254 B.n165 B.n164 585
R255 B.n334 B.n333 585
R256 B.n333 B.n332 585
R257 B.n167 B.n166 585
R258 B.n325 B.n167 585
R259 B.n324 B.n323 585
R260 B.n326 B.n324 585
R261 B.n322 B.n172 585
R262 B.n172 B.n171 585
R263 B.n321 B.n320 585
R264 B.n320 B.n319 585
R265 B.n174 B.n173 585
R266 B.n175 B.n174 585
R267 B.n312 B.n311 585
R268 B.n313 B.n312 585
R269 B.n310 B.n180 585
R270 B.n180 B.n179 585
R271 B.n309 B.n308 585
R272 B.n308 B.n307 585
R273 B.n182 B.n181 585
R274 B.n183 B.n182 585
R275 B.n300 B.n299 585
R276 B.n301 B.n300 585
R277 B.n298 B.n188 585
R278 B.n188 B.n187 585
R279 B.n297 B.n296 585
R280 B.n296 B.n295 585
R281 B.n190 B.n189 585
R282 B.n191 B.n190 585
R283 B.n288 B.n287 585
R284 B.n289 B.n288 585
R285 B.n286 B.n196 585
R286 B.n196 B.n195 585
R287 B.n280 B.n279 585
R288 B.n278 B.n214 585
R289 B.n277 B.n213 585
R290 B.n282 B.n213 585
R291 B.n276 B.n275 585
R292 B.n274 B.n273 585
R293 B.n272 B.n271 585
R294 B.n270 B.n269 585
R295 B.n268 B.n267 585
R296 B.n266 B.n265 585
R297 B.n264 B.n263 585
R298 B.n262 B.n261 585
R299 B.n260 B.n259 585
R300 B.n257 B.n256 585
R301 B.n255 B.n254 585
R302 B.n253 B.n252 585
R303 B.n251 B.n250 585
R304 B.n249 B.n248 585
R305 B.n247 B.n246 585
R306 B.n245 B.n244 585
R307 B.n243 B.n242 585
R308 B.n241 B.n240 585
R309 B.n239 B.n238 585
R310 B.n237 B.n236 585
R311 B.n235 B.n234 585
R312 B.n233 B.n232 585
R313 B.n231 B.n230 585
R314 B.n229 B.n228 585
R315 B.n227 B.n226 585
R316 B.n225 B.n224 585
R317 B.n223 B.n222 585
R318 B.n221 B.n220 585
R319 B.n198 B.n197 585
R320 B.n285 B.n284 585
R321 B.n194 B.n193 585
R322 B.n195 B.n194 585
R323 B.n291 B.n290 585
R324 B.n290 B.n289 585
R325 B.n292 B.n192 585
R326 B.n192 B.n191 585
R327 B.n294 B.n293 585
R328 B.n295 B.n294 585
R329 B.n186 B.n185 585
R330 B.n187 B.n186 585
R331 B.n303 B.n302 585
R332 B.n302 B.n301 585
R333 B.n304 B.n184 585
R334 B.n184 B.n183 585
R335 B.n306 B.n305 585
R336 B.n307 B.n306 585
R337 B.n178 B.n177 585
R338 B.n179 B.n178 585
R339 B.n315 B.n314 585
R340 B.n314 B.n313 585
R341 B.n316 B.n176 585
R342 B.n176 B.n175 585
R343 B.n318 B.n317 585
R344 B.n319 B.n318 585
R345 B.n170 B.n169 585
R346 B.n171 B.n170 585
R347 B.n328 B.n327 585
R348 B.n327 B.n326 585
R349 B.n329 B.n168 585
R350 B.n325 B.n168 585
R351 B.n331 B.n330 585
R352 B.n332 B.n331 585
R353 B.n163 B.n162 585
R354 B.n164 B.n163 585
R355 B.n340 B.n339 585
R356 B.n339 B.n338 585
R357 B.n341 B.n161 585
R358 B.n161 B.n160 585
R359 B.n343 B.n342 585
R360 B.n344 B.n343 585
R361 B.n155 B.n154 585
R362 B.n156 B.n155 585
R363 B.n352 B.n351 585
R364 B.n351 B.n350 585
R365 B.n353 B.n153 585
R366 B.n153 B.n151 585
R367 B.n355 B.n354 585
R368 B.n356 B.n355 585
R369 B.n147 B.n146 585
R370 B.n152 B.n147 585
R371 B.n365 B.n364 585
R372 B.n364 B.n363 585
R373 B.n366 B.n145 585
R374 B.n145 B.n144 585
R375 B.n368 B.n367 585
R376 B.n369 B.n368 585
R377 B.n2 B.n0 585
R378 B.n4 B.n2 585
R379 B.n3 B.n1 585
R380 B.n469 B.n3 585
R381 B.n467 B.n466 585
R382 B.n468 B.n467 585
R383 B.n465 B.n9 585
R384 B.n9 B.n8 585
R385 B.n464 B.n463 585
R386 B.n463 B.n462 585
R387 B.n11 B.n10 585
R388 B.n461 B.n11 585
R389 B.n459 B.n458 585
R390 B.n460 B.n459 585
R391 B.n457 B.n16 585
R392 B.n16 B.n15 585
R393 B.n456 B.n455 585
R394 B.n455 B.n454 585
R395 B.n18 B.n17 585
R396 B.n453 B.n18 585
R397 B.n451 B.n450 585
R398 B.n452 B.n451 585
R399 B.n449 B.n23 585
R400 B.n23 B.n22 585
R401 B.n448 B.n447 585
R402 B.n447 B.n446 585
R403 B.n25 B.n24 585
R404 B.n445 B.n25 585
R405 B.n443 B.n442 585
R406 B.n444 B.n443 585
R407 B.n441 B.n29 585
R408 B.n32 B.n29 585
R409 B.n440 B.n439 585
R410 B.n439 B.n438 585
R411 B.n31 B.n30 585
R412 B.n437 B.n31 585
R413 B.n435 B.n434 585
R414 B.n436 B.n435 585
R415 B.n433 B.n37 585
R416 B.n37 B.n36 585
R417 B.n432 B.n431 585
R418 B.n431 B.n430 585
R419 B.n39 B.n38 585
R420 B.n429 B.n39 585
R421 B.n427 B.n426 585
R422 B.n428 B.n427 585
R423 B.n425 B.n44 585
R424 B.n44 B.n43 585
R425 B.n424 B.n423 585
R426 B.n423 B.n422 585
R427 B.n46 B.n45 585
R428 B.n421 B.n46 585
R429 B.n419 B.n418 585
R430 B.n420 B.n419 585
R431 B.n417 B.n51 585
R432 B.n51 B.n50 585
R433 B.n416 B.n415 585
R434 B.n415 B.n414 585
R435 B.n53 B.n52 585
R436 B.n413 B.n53 585
R437 B.n472 B.n471 585
R438 B.n471 B.n470 585
R439 B.n280 B.n194 521.33
R440 B.n78 B.n53 521.33
R441 B.n284 B.n196 521.33
R442 B.n411 B.n55 521.33
R443 B.n412 B.n71 256.663
R444 B.n412 B.n70 256.663
R445 B.n412 B.n69 256.663
R446 B.n412 B.n68 256.663
R447 B.n412 B.n67 256.663
R448 B.n412 B.n66 256.663
R449 B.n412 B.n65 256.663
R450 B.n412 B.n64 256.663
R451 B.n412 B.n63 256.663
R452 B.n412 B.n62 256.663
R453 B.n412 B.n61 256.663
R454 B.n412 B.n60 256.663
R455 B.n412 B.n59 256.663
R456 B.n412 B.n58 256.663
R457 B.n412 B.n57 256.663
R458 B.n412 B.n56 256.663
R459 B.n282 B.n281 256.663
R460 B.n282 B.n199 256.663
R461 B.n282 B.n200 256.663
R462 B.n282 B.n201 256.663
R463 B.n282 B.n202 256.663
R464 B.n282 B.n203 256.663
R465 B.n282 B.n204 256.663
R466 B.n282 B.n205 256.663
R467 B.n282 B.n206 256.663
R468 B.n282 B.n207 256.663
R469 B.n282 B.n208 256.663
R470 B.n282 B.n209 256.663
R471 B.n282 B.n210 256.663
R472 B.n282 B.n211 256.663
R473 B.n282 B.n212 256.663
R474 B.n283 B.n282 256.663
R475 B.n217 B.t17 235.974
R476 B.n73 B.t10 235.974
R477 B.n215 B.t13 235.496
R478 B.n75 B.t6 235.496
R479 B.n282 B.n195 209.303
R480 B.n413 B.n412 209.303
R481 B.n290 B.n194 163.367
R482 B.n290 B.n192 163.367
R483 B.n294 B.n192 163.367
R484 B.n294 B.n186 163.367
R485 B.n302 B.n186 163.367
R486 B.n302 B.n184 163.367
R487 B.n306 B.n184 163.367
R488 B.n306 B.n178 163.367
R489 B.n314 B.n178 163.367
R490 B.n314 B.n176 163.367
R491 B.n318 B.n176 163.367
R492 B.n318 B.n170 163.367
R493 B.n327 B.n170 163.367
R494 B.n327 B.n168 163.367
R495 B.n331 B.n168 163.367
R496 B.n331 B.n163 163.367
R497 B.n339 B.n163 163.367
R498 B.n339 B.n161 163.367
R499 B.n343 B.n161 163.367
R500 B.n343 B.n155 163.367
R501 B.n351 B.n155 163.367
R502 B.n351 B.n153 163.367
R503 B.n355 B.n153 163.367
R504 B.n355 B.n147 163.367
R505 B.n364 B.n147 163.367
R506 B.n364 B.n145 163.367
R507 B.n368 B.n145 163.367
R508 B.n368 B.n2 163.367
R509 B.n471 B.n2 163.367
R510 B.n471 B.n3 163.367
R511 B.n467 B.n3 163.367
R512 B.n467 B.n9 163.367
R513 B.n463 B.n9 163.367
R514 B.n463 B.n11 163.367
R515 B.n459 B.n11 163.367
R516 B.n459 B.n16 163.367
R517 B.n455 B.n16 163.367
R518 B.n455 B.n18 163.367
R519 B.n451 B.n18 163.367
R520 B.n451 B.n23 163.367
R521 B.n447 B.n23 163.367
R522 B.n447 B.n25 163.367
R523 B.n443 B.n25 163.367
R524 B.n443 B.n29 163.367
R525 B.n439 B.n29 163.367
R526 B.n439 B.n31 163.367
R527 B.n435 B.n31 163.367
R528 B.n435 B.n37 163.367
R529 B.n431 B.n37 163.367
R530 B.n431 B.n39 163.367
R531 B.n427 B.n39 163.367
R532 B.n427 B.n44 163.367
R533 B.n423 B.n44 163.367
R534 B.n423 B.n46 163.367
R535 B.n419 B.n46 163.367
R536 B.n419 B.n51 163.367
R537 B.n415 B.n51 163.367
R538 B.n415 B.n53 163.367
R539 B.n214 B.n213 163.367
R540 B.n275 B.n213 163.367
R541 B.n273 B.n272 163.367
R542 B.n269 B.n268 163.367
R543 B.n265 B.n264 163.367
R544 B.n261 B.n260 163.367
R545 B.n256 B.n255 163.367
R546 B.n252 B.n251 163.367
R547 B.n248 B.n247 163.367
R548 B.n244 B.n243 163.367
R549 B.n240 B.n239 163.367
R550 B.n236 B.n235 163.367
R551 B.n232 B.n231 163.367
R552 B.n228 B.n227 163.367
R553 B.n224 B.n223 163.367
R554 B.n220 B.n198 163.367
R555 B.n288 B.n196 163.367
R556 B.n288 B.n190 163.367
R557 B.n296 B.n190 163.367
R558 B.n296 B.n188 163.367
R559 B.n300 B.n188 163.367
R560 B.n300 B.n182 163.367
R561 B.n308 B.n182 163.367
R562 B.n308 B.n180 163.367
R563 B.n312 B.n180 163.367
R564 B.n312 B.n174 163.367
R565 B.n320 B.n174 163.367
R566 B.n320 B.n172 163.367
R567 B.n324 B.n172 163.367
R568 B.n324 B.n167 163.367
R569 B.n333 B.n167 163.367
R570 B.n333 B.n165 163.367
R571 B.n337 B.n165 163.367
R572 B.n337 B.n159 163.367
R573 B.n345 B.n159 163.367
R574 B.n345 B.n157 163.367
R575 B.n349 B.n157 163.367
R576 B.n349 B.n150 163.367
R577 B.n357 B.n150 163.367
R578 B.n357 B.n148 163.367
R579 B.n362 B.n148 163.367
R580 B.n362 B.n143 163.367
R581 B.n370 B.n143 163.367
R582 B.n371 B.n370 163.367
R583 B.n371 B.n5 163.367
R584 B.n6 B.n5 163.367
R585 B.n7 B.n6 163.367
R586 B.n376 B.n7 163.367
R587 B.n376 B.n12 163.367
R588 B.n13 B.n12 163.367
R589 B.n14 B.n13 163.367
R590 B.n381 B.n14 163.367
R591 B.n381 B.n19 163.367
R592 B.n20 B.n19 163.367
R593 B.n21 B.n20 163.367
R594 B.n386 B.n21 163.367
R595 B.n386 B.n26 163.367
R596 B.n27 B.n26 163.367
R597 B.n28 B.n27 163.367
R598 B.n391 B.n28 163.367
R599 B.n391 B.n33 163.367
R600 B.n34 B.n33 163.367
R601 B.n35 B.n34 163.367
R602 B.n396 B.n35 163.367
R603 B.n396 B.n40 163.367
R604 B.n41 B.n40 163.367
R605 B.n42 B.n41 163.367
R606 B.n401 B.n42 163.367
R607 B.n401 B.n47 163.367
R608 B.n48 B.n47 163.367
R609 B.n49 B.n48 163.367
R610 B.n406 B.n49 163.367
R611 B.n406 B.n54 163.367
R612 B.n55 B.n54 163.367
R613 B.n82 B.n81 163.367
R614 B.n86 B.n85 163.367
R615 B.n90 B.n89 163.367
R616 B.n94 B.n93 163.367
R617 B.n98 B.n97 163.367
R618 B.n102 B.n101 163.367
R619 B.n106 B.n105 163.367
R620 B.n110 B.n109 163.367
R621 B.n114 B.n113 163.367
R622 B.n118 B.n117 163.367
R623 B.n123 B.n122 163.367
R624 B.n127 B.n126 163.367
R625 B.n131 B.n130 163.367
R626 B.n135 B.n134 163.367
R627 B.n139 B.n138 163.367
R628 B.n411 B.n72 163.367
R629 B.n217 B.t19 154.436
R630 B.n73 B.t11 154.436
R631 B.n215 B.t16 154.436
R632 B.n75 B.t8 154.436
R633 B.n218 B.t18 119.722
R634 B.n74 B.t12 119.722
R635 B.n216 B.t15 119.722
R636 B.n76 B.t9 119.722
R637 B.n289 B.n195 105.427
R638 B.n289 B.n191 105.427
R639 B.n295 B.n191 105.427
R640 B.n295 B.n187 105.427
R641 B.n301 B.n187 105.427
R642 B.n307 B.n183 105.427
R643 B.n307 B.n179 105.427
R644 B.n313 B.n179 105.427
R645 B.n313 B.n175 105.427
R646 B.n319 B.n175 105.427
R647 B.n319 B.n171 105.427
R648 B.n326 B.n171 105.427
R649 B.n326 B.n325 105.427
R650 B.n332 B.n164 105.427
R651 B.n338 B.n164 105.427
R652 B.n338 B.n160 105.427
R653 B.n344 B.n160 105.427
R654 B.n350 B.n156 105.427
R655 B.n350 B.n151 105.427
R656 B.n356 B.n151 105.427
R657 B.n356 B.n152 105.427
R658 B.n363 B.n144 105.427
R659 B.n369 B.n144 105.427
R660 B.n369 B.n4 105.427
R661 B.n470 B.n4 105.427
R662 B.n470 B.n469 105.427
R663 B.n469 B.n468 105.427
R664 B.n468 B.n8 105.427
R665 B.n462 B.n8 105.427
R666 B.n461 B.n460 105.427
R667 B.n460 B.n15 105.427
R668 B.n454 B.n15 105.427
R669 B.n454 B.n453 105.427
R670 B.n452 B.n22 105.427
R671 B.n446 B.n22 105.427
R672 B.n446 B.n445 105.427
R673 B.n445 B.n444 105.427
R674 B.n438 B.n32 105.427
R675 B.n438 B.n437 105.427
R676 B.n437 B.n436 105.427
R677 B.n436 B.n36 105.427
R678 B.n430 B.n36 105.427
R679 B.n430 B.n429 105.427
R680 B.n429 B.n428 105.427
R681 B.n428 B.n43 105.427
R682 B.n422 B.n421 105.427
R683 B.n421 B.n420 105.427
R684 B.n420 B.n50 105.427
R685 B.n414 B.n50 105.427
R686 B.n414 B.n413 105.427
R687 B.n301 B.t14 80.6207
R688 B.n332 B.t2 80.6207
R689 B.n152 B.t3 80.6207
R690 B.t5 B.n461 80.6207
R691 B.n444 B.t4 80.6207
R692 B.n422 B.t7 80.6207
R693 B.n281 B.n280 71.676
R694 B.n275 B.n199 71.676
R695 B.n272 B.n200 71.676
R696 B.n268 B.n201 71.676
R697 B.n264 B.n202 71.676
R698 B.n260 B.n203 71.676
R699 B.n255 B.n204 71.676
R700 B.n251 B.n205 71.676
R701 B.n247 B.n206 71.676
R702 B.n243 B.n207 71.676
R703 B.n239 B.n208 71.676
R704 B.n235 B.n209 71.676
R705 B.n231 B.n210 71.676
R706 B.n227 B.n211 71.676
R707 B.n223 B.n212 71.676
R708 B.n283 B.n198 71.676
R709 B.n78 B.n56 71.676
R710 B.n82 B.n57 71.676
R711 B.n86 B.n58 71.676
R712 B.n90 B.n59 71.676
R713 B.n94 B.n60 71.676
R714 B.n98 B.n61 71.676
R715 B.n102 B.n62 71.676
R716 B.n106 B.n63 71.676
R717 B.n110 B.n64 71.676
R718 B.n114 B.n65 71.676
R719 B.n118 B.n66 71.676
R720 B.n123 B.n67 71.676
R721 B.n127 B.n68 71.676
R722 B.n131 B.n69 71.676
R723 B.n135 B.n70 71.676
R724 B.n139 B.n71 71.676
R725 B.n72 B.n71 71.676
R726 B.n138 B.n70 71.676
R727 B.n134 B.n69 71.676
R728 B.n130 B.n68 71.676
R729 B.n126 B.n67 71.676
R730 B.n122 B.n66 71.676
R731 B.n117 B.n65 71.676
R732 B.n113 B.n64 71.676
R733 B.n109 B.n63 71.676
R734 B.n105 B.n62 71.676
R735 B.n101 B.n61 71.676
R736 B.n97 B.n60 71.676
R737 B.n93 B.n59 71.676
R738 B.n89 B.n58 71.676
R739 B.n85 B.n57 71.676
R740 B.n81 B.n56 71.676
R741 B.n281 B.n214 71.676
R742 B.n273 B.n199 71.676
R743 B.n269 B.n200 71.676
R744 B.n265 B.n201 71.676
R745 B.n261 B.n202 71.676
R746 B.n256 B.n203 71.676
R747 B.n252 B.n204 71.676
R748 B.n248 B.n205 71.676
R749 B.n244 B.n206 71.676
R750 B.n240 B.n207 71.676
R751 B.n236 B.n208 71.676
R752 B.n232 B.n209 71.676
R753 B.n228 B.n210 71.676
R754 B.n224 B.n211 71.676
R755 B.n220 B.n212 71.676
R756 B.n284 B.n283 71.676
R757 B.n219 B.n218 59.5399
R758 B.n258 B.n216 59.5399
R759 B.n77 B.n76 59.5399
R760 B.n120 B.n74 59.5399
R761 B.n344 B.t1 52.7137
R762 B.t1 B.n156 52.7137
R763 B.n453 B.t0 52.7137
R764 B.t0 B.n452 52.7137
R765 B.n218 B.n217 34.7157
R766 B.n216 B.n215 34.7157
R767 B.n76 B.n75 34.7157
R768 B.n74 B.n73 34.7157
R769 B.n79 B.n52 33.8737
R770 B.n410 B.n409 33.8737
R771 B.n286 B.n285 33.8737
R772 B.n279 B.n193 33.8737
R773 B.t14 B.n183 24.8067
R774 B.n325 B.t2 24.8067
R775 B.n363 B.t3 24.8067
R776 B.n462 B.t5 24.8067
R777 B.n32 B.t4 24.8067
R778 B.t7 B.n43 24.8067
R779 B B.n472 18.0485
R780 B.n80 B.n79 10.6151
R781 B.n83 B.n80 10.6151
R782 B.n84 B.n83 10.6151
R783 B.n87 B.n84 10.6151
R784 B.n88 B.n87 10.6151
R785 B.n91 B.n88 10.6151
R786 B.n92 B.n91 10.6151
R787 B.n95 B.n92 10.6151
R788 B.n96 B.n95 10.6151
R789 B.n99 B.n96 10.6151
R790 B.n100 B.n99 10.6151
R791 B.n104 B.n103 10.6151
R792 B.n107 B.n104 10.6151
R793 B.n108 B.n107 10.6151
R794 B.n111 B.n108 10.6151
R795 B.n112 B.n111 10.6151
R796 B.n115 B.n112 10.6151
R797 B.n116 B.n115 10.6151
R798 B.n119 B.n116 10.6151
R799 B.n124 B.n121 10.6151
R800 B.n125 B.n124 10.6151
R801 B.n128 B.n125 10.6151
R802 B.n129 B.n128 10.6151
R803 B.n132 B.n129 10.6151
R804 B.n133 B.n132 10.6151
R805 B.n136 B.n133 10.6151
R806 B.n137 B.n136 10.6151
R807 B.n140 B.n137 10.6151
R808 B.n141 B.n140 10.6151
R809 B.n410 B.n141 10.6151
R810 B.n287 B.n286 10.6151
R811 B.n287 B.n189 10.6151
R812 B.n297 B.n189 10.6151
R813 B.n298 B.n297 10.6151
R814 B.n299 B.n298 10.6151
R815 B.n299 B.n181 10.6151
R816 B.n309 B.n181 10.6151
R817 B.n310 B.n309 10.6151
R818 B.n311 B.n310 10.6151
R819 B.n311 B.n173 10.6151
R820 B.n321 B.n173 10.6151
R821 B.n322 B.n321 10.6151
R822 B.n323 B.n322 10.6151
R823 B.n323 B.n166 10.6151
R824 B.n334 B.n166 10.6151
R825 B.n335 B.n334 10.6151
R826 B.n336 B.n335 10.6151
R827 B.n336 B.n158 10.6151
R828 B.n346 B.n158 10.6151
R829 B.n347 B.n346 10.6151
R830 B.n348 B.n347 10.6151
R831 B.n348 B.n149 10.6151
R832 B.n358 B.n149 10.6151
R833 B.n359 B.n358 10.6151
R834 B.n361 B.n359 10.6151
R835 B.n361 B.n360 10.6151
R836 B.n360 B.n142 10.6151
R837 B.n372 B.n142 10.6151
R838 B.n373 B.n372 10.6151
R839 B.n374 B.n373 10.6151
R840 B.n375 B.n374 10.6151
R841 B.n377 B.n375 10.6151
R842 B.n378 B.n377 10.6151
R843 B.n379 B.n378 10.6151
R844 B.n380 B.n379 10.6151
R845 B.n382 B.n380 10.6151
R846 B.n383 B.n382 10.6151
R847 B.n384 B.n383 10.6151
R848 B.n385 B.n384 10.6151
R849 B.n387 B.n385 10.6151
R850 B.n388 B.n387 10.6151
R851 B.n389 B.n388 10.6151
R852 B.n390 B.n389 10.6151
R853 B.n392 B.n390 10.6151
R854 B.n393 B.n392 10.6151
R855 B.n394 B.n393 10.6151
R856 B.n395 B.n394 10.6151
R857 B.n397 B.n395 10.6151
R858 B.n398 B.n397 10.6151
R859 B.n399 B.n398 10.6151
R860 B.n400 B.n399 10.6151
R861 B.n402 B.n400 10.6151
R862 B.n403 B.n402 10.6151
R863 B.n404 B.n403 10.6151
R864 B.n405 B.n404 10.6151
R865 B.n407 B.n405 10.6151
R866 B.n408 B.n407 10.6151
R867 B.n409 B.n408 10.6151
R868 B.n279 B.n278 10.6151
R869 B.n278 B.n277 10.6151
R870 B.n277 B.n276 10.6151
R871 B.n276 B.n274 10.6151
R872 B.n274 B.n271 10.6151
R873 B.n271 B.n270 10.6151
R874 B.n270 B.n267 10.6151
R875 B.n267 B.n266 10.6151
R876 B.n266 B.n263 10.6151
R877 B.n263 B.n262 10.6151
R878 B.n262 B.n259 10.6151
R879 B.n257 B.n254 10.6151
R880 B.n254 B.n253 10.6151
R881 B.n253 B.n250 10.6151
R882 B.n250 B.n249 10.6151
R883 B.n249 B.n246 10.6151
R884 B.n246 B.n245 10.6151
R885 B.n245 B.n242 10.6151
R886 B.n242 B.n241 10.6151
R887 B.n238 B.n237 10.6151
R888 B.n237 B.n234 10.6151
R889 B.n234 B.n233 10.6151
R890 B.n233 B.n230 10.6151
R891 B.n230 B.n229 10.6151
R892 B.n229 B.n226 10.6151
R893 B.n226 B.n225 10.6151
R894 B.n225 B.n222 10.6151
R895 B.n222 B.n221 10.6151
R896 B.n221 B.n197 10.6151
R897 B.n285 B.n197 10.6151
R898 B.n291 B.n193 10.6151
R899 B.n292 B.n291 10.6151
R900 B.n293 B.n292 10.6151
R901 B.n293 B.n185 10.6151
R902 B.n303 B.n185 10.6151
R903 B.n304 B.n303 10.6151
R904 B.n305 B.n304 10.6151
R905 B.n305 B.n177 10.6151
R906 B.n315 B.n177 10.6151
R907 B.n316 B.n315 10.6151
R908 B.n317 B.n316 10.6151
R909 B.n317 B.n169 10.6151
R910 B.n328 B.n169 10.6151
R911 B.n329 B.n328 10.6151
R912 B.n330 B.n329 10.6151
R913 B.n330 B.n162 10.6151
R914 B.n340 B.n162 10.6151
R915 B.n341 B.n340 10.6151
R916 B.n342 B.n341 10.6151
R917 B.n342 B.n154 10.6151
R918 B.n352 B.n154 10.6151
R919 B.n353 B.n352 10.6151
R920 B.n354 B.n353 10.6151
R921 B.n354 B.n146 10.6151
R922 B.n365 B.n146 10.6151
R923 B.n366 B.n365 10.6151
R924 B.n367 B.n366 10.6151
R925 B.n367 B.n0 10.6151
R926 B.n466 B.n1 10.6151
R927 B.n466 B.n465 10.6151
R928 B.n465 B.n464 10.6151
R929 B.n464 B.n10 10.6151
R930 B.n458 B.n10 10.6151
R931 B.n458 B.n457 10.6151
R932 B.n457 B.n456 10.6151
R933 B.n456 B.n17 10.6151
R934 B.n450 B.n17 10.6151
R935 B.n450 B.n449 10.6151
R936 B.n449 B.n448 10.6151
R937 B.n448 B.n24 10.6151
R938 B.n442 B.n24 10.6151
R939 B.n442 B.n441 10.6151
R940 B.n441 B.n440 10.6151
R941 B.n440 B.n30 10.6151
R942 B.n434 B.n30 10.6151
R943 B.n434 B.n433 10.6151
R944 B.n433 B.n432 10.6151
R945 B.n432 B.n38 10.6151
R946 B.n426 B.n38 10.6151
R947 B.n426 B.n425 10.6151
R948 B.n425 B.n424 10.6151
R949 B.n424 B.n45 10.6151
R950 B.n418 B.n45 10.6151
R951 B.n418 B.n417 10.6151
R952 B.n417 B.n416 10.6151
R953 B.n416 B.n52 10.6151
R954 B.n103 B.n77 6.4005
R955 B.n120 B.n119 6.4005
R956 B.n258 B.n257 6.4005
R957 B.n241 B.n219 6.4005
R958 B.n100 B.n77 4.21513
R959 B.n121 B.n120 4.21513
R960 B.n259 B.n258 4.21513
R961 B.n238 B.n219 4.21513
R962 B.n472 B.n0 2.81026
R963 B.n472 B.n1 2.81026
R964 VP.n15 VP.n14 171.524
R965 VP.n27 VP.n26 171.524
R966 VP.n13 VP.n12 171.524
R967 VP.n8 VP.n5 161.3
R968 VP.n10 VP.n9 161.3
R969 VP.n11 VP.n4 161.3
R970 VP.n25 VP.n0 161.3
R971 VP.n24 VP.n23 161.3
R972 VP.n22 VP.n1 161.3
R973 VP.n21 VP.n20 161.3
R974 VP.n19 VP.n2 161.3
R975 VP.n18 VP.n17 161.3
R976 VP.n16 VP.n3 161.3
R977 VP.n7 VP.t0 66.583
R978 VP.n19 VP.n18 50.6348
R979 VP.n24 VP.n1 50.6348
R980 VP.n10 VP.n5 50.6348
R981 VP.n7 VP.n6 41.7711
R982 VP.n15 VP.n13 36.474
R983 VP.n18 VP.n3 30.1864
R984 VP.n25 VP.n24 30.1864
R985 VP.n11 VP.n10 30.1864
R986 VP.n20 VP.t3 30.043
R987 VP.n14 VP.t1 30.043
R988 VP.n26 VP.t4 30.043
R989 VP.n6 VP.t2 30.043
R990 VP.n12 VP.t5 30.043
R991 VP.n20 VP.n19 24.3439
R992 VP.n20 VP.n1 24.3439
R993 VP.n6 VP.n5 24.3439
R994 VP.n8 VP.n7 17.3537
R995 VP.n14 VP.n3 14.1197
R996 VP.n26 VP.n25 14.1197
R997 VP.n12 VP.n11 14.1197
R998 VP.n9 VP.n8 0.189894
R999 VP.n9 VP.n4 0.189894
R1000 VP.n13 VP.n4 0.189894
R1001 VP.n16 VP.n15 0.189894
R1002 VP.n17 VP.n16 0.189894
R1003 VP.n17 VP.n2 0.189894
R1004 VP.n21 VP.n2 0.189894
R1005 VP.n22 VP.n21 0.189894
R1006 VP.n23 VP.n22 0.189894
R1007 VP.n23 VP.n0 0.189894
R1008 VP.n27 VP.n0 0.189894
R1009 VP VP.n27 0.0516364
R1010 VDD1.n2 VDD1.n0 289.615
R1011 VDD1.n9 VDD1.n7 289.615
R1012 VDD1.n3 VDD1.n2 185
R1013 VDD1.n10 VDD1.n9 185
R1014 VDD1.t5 VDD1.n1 164.876
R1015 VDD1.t4 VDD1.n8 164.876
R1016 VDD1.n15 VDD1.n14 102.529
R1017 VDD1.n17 VDD1.n16 102.198
R1018 VDD1 VDD1.n6 52.7948
R1019 VDD1.n15 VDD1.n13 52.6813
R1020 VDD1.n2 VDD1.t5 52.3082
R1021 VDD1.n9 VDD1.t4 52.3082
R1022 VDD1.n17 VDD1.n15 31.6539
R1023 VDD1.n3 VDD1.n1 14.7318
R1024 VDD1.n10 VDD1.n8 14.7318
R1025 VDD1.n4 VDD1.n0 12.8005
R1026 VDD1.n11 VDD1.n7 12.8005
R1027 VDD1.n16 VDD1.t3 10.8796
R1028 VDD1.n16 VDD1.t0 10.8796
R1029 VDD1.n14 VDD1.t2 10.8796
R1030 VDD1.n14 VDD1.t1 10.8796
R1031 VDD1.n6 VDD1.n5 9.45567
R1032 VDD1.n13 VDD1.n12 9.45567
R1033 VDD1.n5 VDD1.n4 9.3005
R1034 VDD1.n12 VDD1.n11 9.3005
R1035 VDD1.n5 VDD1.n1 5.62509
R1036 VDD1.n12 VDD1.n8 5.62509
R1037 VDD1.n6 VDD1.n0 1.16414
R1038 VDD1.n13 VDD1.n7 1.16414
R1039 VDD1.n4 VDD1.n3 0.388379
R1040 VDD1.n11 VDD1.n10 0.388379
R1041 VDD1 VDD1.n17 0.328086
C0 VN VDD1 0.155446f
C1 VTAIL VDD2 3.353f
C2 VP VDD1 1.40448f
C3 VTAIL VDD1 3.30776f
C4 VDD1 VDD2 0.989825f
C5 VN VP 3.94276f
C6 VTAIL VN 1.67397f
C7 VN VDD2 1.19425f
C8 VTAIL VP 1.68813f
C9 VP VDD2 0.367805f
C10 VDD2 B 3.128894f
C11 VDD1 B 3.250491f
C12 VTAIL B 2.739053f
C13 VN B 8.077646f
C14 VP B 7.170011f
C15 VDD1.n0 B 0.021715f
C16 VDD1.n1 B 0.050896f
C17 VDD1.t5 B 0.036313f
C18 VDD1.n2 B 0.037531f
C19 VDD1.n3 B 0.010743f
C20 VDD1.n4 B 0.00872f
C21 VDD1.n5 B 0.099657f
C22 VDD1.n6 B 0.037183f
C23 VDD1.n7 B 0.021715f
C24 VDD1.n8 B 0.050896f
C25 VDD1.t4 B 0.036313f
C26 VDD1.n9 B 0.037531f
C27 VDD1.n10 B 0.010743f
C28 VDD1.n11 B 0.00872f
C29 VDD1.n12 B 0.099657f
C30 VDD1.n13 B 0.036863f
C31 VDD1.t2 B 0.023339f
C32 VDD1.t1 B 0.023339f
C33 VDD1.n14 B 0.150269f
C34 VDD1.n15 B 1.06861f
C35 VDD1.t3 B 0.023339f
C36 VDD1.t0 B 0.023339f
C37 VDD1.n16 B 0.149563f
C38 VDD1.n17 B 1.05795f
C39 VP.n0 B 0.023246f
C40 VP.t4 B 0.14077f
C41 VP.n1 B 0.042649f
C42 VP.n2 B 0.023246f
C43 VP.t3 B 0.14077f
C44 VP.n3 B 0.037675f
C45 VP.n4 B 0.023246f
C46 VP.t5 B 0.14077f
C47 VP.n5 B 0.042649f
C48 VP.t0 B 0.234071f
C49 VP.t2 B 0.14077f
C50 VP.n6 B 0.13355f
C51 VP.n7 B 0.10993f
C52 VP.n8 B 0.147853f
C53 VP.n9 B 0.023246f
C54 VP.n10 B 0.022354f
C55 VP.n11 B 0.037675f
C56 VP.n12 B 0.130257f
C57 VP.n13 B 0.752207f
C58 VP.t1 B 0.14077f
C59 VP.n14 B 0.130257f
C60 VP.n15 B 0.775051f
C61 VP.n16 B 0.023246f
C62 VP.n17 B 0.023246f
C63 VP.n18 B 0.022354f
C64 VP.n19 B 0.042649f
C65 VP.n20 B 0.101245f
C66 VP.n21 B 0.023246f
C67 VP.n22 B 0.023246f
C68 VP.n23 B 0.023246f
C69 VP.n24 B 0.022354f
C70 VP.n25 B 0.037675f
C71 VP.n26 B 0.130257f
C72 VP.n27 B 0.021251f
C73 VTAIL.t10 B 0.031457f
C74 VTAIL.t11 B 0.031457f
C75 VTAIL.n0 B 0.172476f
C76 VTAIL.n1 B 0.271545f
C77 VTAIL.n2 B 0.029267f
C78 VTAIL.n3 B 0.068598f
C79 VTAIL.t3 B 0.048943f
C80 VTAIL.n4 B 0.050585f
C81 VTAIL.n5 B 0.014479f
C82 VTAIL.n6 B 0.011753f
C83 VTAIL.n7 B 0.134318f
C84 VTAIL.n8 B 0.032046f
C85 VTAIL.n9 B 0.217288f
C86 VTAIL.t2 B 0.031457f
C87 VTAIL.t1 B 0.031457f
C88 VTAIL.n10 B 0.172476f
C89 VTAIL.n11 B 0.88671f
C90 VTAIL.t8 B 0.031457f
C91 VTAIL.t9 B 0.031457f
C92 VTAIL.n12 B 0.172477f
C93 VTAIL.n13 B 0.886709f
C94 VTAIL.n14 B 0.029267f
C95 VTAIL.n15 B 0.068598f
C96 VTAIL.t6 B 0.048943f
C97 VTAIL.n16 B 0.050585f
C98 VTAIL.n17 B 0.014479f
C99 VTAIL.n18 B 0.011753f
C100 VTAIL.n19 B 0.134318f
C101 VTAIL.n20 B 0.032046f
C102 VTAIL.n21 B 0.217288f
C103 VTAIL.t5 B 0.031457f
C104 VTAIL.t0 B 0.031457f
C105 VTAIL.n22 B 0.172477f
C106 VTAIL.n23 B 0.349008f
C107 VTAIL.n24 B 0.029267f
C108 VTAIL.n25 B 0.068598f
C109 VTAIL.t4 B 0.048943f
C110 VTAIL.n26 B 0.050585f
C111 VTAIL.n27 B 0.014479f
C112 VTAIL.n28 B 0.011753f
C113 VTAIL.n29 B 0.134318f
C114 VTAIL.n30 B 0.032046f
C115 VTAIL.n31 B 0.646235f
C116 VTAIL.n32 B 0.029267f
C117 VTAIL.n33 B 0.068598f
C118 VTAIL.t7 B 0.048943f
C119 VTAIL.n34 B 0.050585f
C120 VTAIL.n35 B 0.014479f
C121 VTAIL.n36 B 0.011753f
C122 VTAIL.n37 B 0.134318f
C123 VTAIL.n38 B 0.032046f
C124 VTAIL.n39 B 0.614946f
C125 VDD2.n0 B 0.022787f
C126 VDD2.n1 B 0.053408f
C127 VDD2.t5 B 0.038105f
C128 VDD2.n2 B 0.039384f
C129 VDD2.n3 B 0.011273f
C130 VDD2.n4 B 0.009151f
C131 VDD2.n5 B 0.104577f
C132 VDD2.n6 B 0.038682f
C133 VDD2.t1 B 0.024492f
C134 VDD2.t2 B 0.024492f
C135 VDD2.n7 B 0.157687f
C136 VDD2.n8 B 1.06196f
C137 VDD2.n9 B 0.022787f
C138 VDD2.n10 B 0.053408f
C139 VDD2.t3 B 0.038105f
C140 VDD2.n11 B 0.039384f
C141 VDD2.n12 B 0.011273f
C142 VDD2.n13 B 0.009151f
C143 VDD2.n14 B 0.104577f
C144 VDD2.n15 B 0.036685f
C145 VDD2.n16 B 0.979095f
C146 VDD2.t4 B 0.024492f
C147 VDD2.t0 B 0.024492f
C148 VDD2.n17 B 0.157677f
C149 VN.n0 B 0.023053f
C150 VN.t4 B 0.1396f
C151 VN.n1 B 0.042295f
C152 VN.t1 B 0.232126f
C153 VN.t0 B 0.1396f
C154 VN.n2 B 0.13244f
C155 VN.n3 B 0.109017f
C156 VN.n4 B 0.146624f
C157 VN.n5 B 0.023053f
C158 VN.n6 B 0.022169f
C159 VN.n7 B 0.037362f
C160 VN.n8 B 0.129174f
C161 VN.n9 B 0.021075f
C162 VN.n10 B 0.023053f
C163 VN.t3 B 0.1396f
C164 VN.n11 B 0.042295f
C165 VN.t5 B 0.232126f
C166 VN.t2 B 0.1396f
C167 VN.n12 B 0.13244f
C168 VN.n13 B 0.109017f
C169 VN.n14 B 0.146624f
C170 VN.n15 B 0.023053f
C171 VN.n16 B 0.022169f
C172 VN.n17 B 0.037362f
C173 VN.n18 B 0.129174f
C174 VN.n19 B 0.761232f
.ends

