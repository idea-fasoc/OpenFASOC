* NGSPICE file created from diff_pair_sample_1228.ext - technology: sky130A

.subckt diff_pair_sample_1228 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=4.8126 ps=25.46 w=12.34 l=1.08
X1 B.t11 B.t9 B.t10 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=0 ps=0 w=12.34 l=1.08
X2 B.t8 B.t6 B.t7 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=0 ps=0 w=12.34 l=1.08
X3 B.t5 B.t3 B.t4 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=0 ps=0 w=12.34 l=1.08
X4 B.t2 B.t0 B.t1 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=0 ps=0 w=12.34 l=1.08
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=4.8126 ps=25.46 w=12.34 l=1.08
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=4.8126 ps=25.46 w=12.34 l=1.08
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1534_n3440# sky130_fd_pr__pfet_01v8 ad=4.8126 pd=25.46 as=4.8126 ps=25.46 w=12.34 l=1.08
R0 VN VN.t1 514.317
R1 VN VN.t0 473.089
R2 VTAIL.n1 VTAIL.t3 63.2454
R3 VTAIL.n3 VTAIL.t2 63.2443
R4 VTAIL.n0 VTAIL.t0 63.2443
R5 VTAIL.n2 VTAIL.t1 63.2442
R6 VTAIL.n1 VTAIL.n0 25.4531
R7 VTAIL.n3 VTAIL.n2 24.2376
R8 VTAIL.n2 VTAIL.n1 1.07809
R9 VTAIL VTAIL.n0 0.832397
R10 VTAIL VTAIL.n3 0.24619
R11 VDD2.n0 VDD2.t1 116.668
R12 VDD2.n0 VDD2.t0 79.923
R13 VDD2 VDD2.n0 0.362569
R14 B.n304 B.n79 585
R15 B.n303 B.n302 585
R16 B.n301 B.n80 585
R17 B.n300 B.n299 585
R18 B.n298 B.n81 585
R19 B.n297 B.n296 585
R20 B.n295 B.n82 585
R21 B.n294 B.n293 585
R22 B.n292 B.n83 585
R23 B.n291 B.n290 585
R24 B.n289 B.n84 585
R25 B.n288 B.n287 585
R26 B.n286 B.n85 585
R27 B.n285 B.n284 585
R28 B.n283 B.n86 585
R29 B.n282 B.n281 585
R30 B.n280 B.n87 585
R31 B.n279 B.n278 585
R32 B.n277 B.n88 585
R33 B.n276 B.n275 585
R34 B.n274 B.n89 585
R35 B.n273 B.n272 585
R36 B.n271 B.n90 585
R37 B.n270 B.n269 585
R38 B.n268 B.n91 585
R39 B.n267 B.n266 585
R40 B.n265 B.n92 585
R41 B.n264 B.n263 585
R42 B.n262 B.n93 585
R43 B.n261 B.n260 585
R44 B.n259 B.n94 585
R45 B.n258 B.n257 585
R46 B.n256 B.n95 585
R47 B.n255 B.n254 585
R48 B.n253 B.n96 585
R49 B.n252 B.n251 585
R50 B.n250 B.n97 585
R51 B.n249 B.n248 585
R52 B.n247 B.n98 585
R53 B.n246 B.n245 585
R54 B.n244 B.n99 585
R55 B.n243 B.n242 585
R56 B.n241 B.n100 585
R57 B.n240 B.n239 585
R58 B.n235 B.n101 585
R59 B.n234 B.n233 585
R60 B.n232 B.n102 585
R61 B.n231 B.n230 585
R62 B.n229 B.n103 585
R63 B.n228 B.n227 585
R64 B.n226 B.n104 585
R65 B.n225 B.n224 585
R66 B.n222 B.n105 585
R67 B.n221 B.n220 585
R68 B.n219 B.n108 585
R69 B.n218 B.n217 585
R70 B.n216 B.n109 585
R71 B.n215 B.n214 585
R72 B.n213 B.n110 585
R73 B.n212 B.n211 585
R74 B.n210 B.n111 585
R75 B.n209 B.n208 585
R76 B.n207 B.n112 585
R77 B.n206 B.n205 585
R78 B.n204 B.n113 585
R79 B.n203 B.n202 585
R80 B.n201 B.n114 585
R81 B.n200 B.n199 585
R82 B.n198 B.n115 585
R83 B.n197 B.n196 585
R84 B.n195 B.n116 585
R85 B.n194 B.n193 585
R86 B.n192 B.n117 585
R87 B.n191 B.n190 585
R88 B.n189 B.n118 585
R89 B.n188 B.n187 585
R90 B.n186 B.n119 585
R91 B.n185 B.n184 585
R92 B.n183 B.n120 585
R93 B.n182 B.n181 585
R94 B.n180 B.n121 585
R95 B.n179 B.n178 585
R96 B.n177 B.n122 585
R97 B.n176 B.n175 585
R98 B.n174 B.n123 585
R99 B.n173 B.n172 585
R100 B.n171 B.n124 585
R101 B.n170 B.n169 585
R102 B.n168 B.n125 585
R103 B.n167 B.n166 585
R104 B.n165 B.n126 585
R105 B.n164 B.n163 585
R106 B.n162 B.n127 585
R107 B.n161 B.n160 585
R108 B.n159 B.n128 585
R109 B.n306 B.n305 585
R110 B.n307 B.n78 585
R111 B.n309 B.n308 585
R112 B.n310 B.n77 585
R113 B.n312 B.n311 585
R114 B.n313 B.n76 585
R115 B.n315 B.n314 585
R116 B.n316 B.n75 585
R117 B.n318 B.n317 585
R118 B.n319 B.n74 585
R119 B.n321 B.n320 585
R120 B.n322 B.n73 585
R121 B.n324 B.n323 585
R122 B.n325 B.n72 585
R123 B.n327 B.n326 585
R124 B.n328 B.n71 585
R125 B.n330 B.n329 585
R126 B.n331 B.n70 585
R127 B.n333 B.n332 585
R128 B.n334 B.n69 585
R129 B.n336 B.n335 585
R130 B.n337 B.n68 585
R131 B.n339 B.n338 585
R132 B.n340 B.n67 585
R133 B.n342 B.n341 585
R134 B.n343 B.n66 585
R135 B.n345 B.n344 585
R136 B.n346 B.n65 585
R137 B.n348 B.n347 585
R138 B.n349 B.n64 585
R139 B.n351 B.n350 585
R140 B.n352 B.n63 585
R141 B.n354 B.n353 585
R142 B.n355 B.n62 585
R143 B.n499 B.n10 585
R144 B.n498 B.n497 585
R145 B.n496 B.n11 585
R146 B.n495 B.n494 585
R147 B.n493 B.n12 585
R148 B.n492 B.n491 585
R149 B.n490 B.n13 585
R150 B.n489 B.n488 585
R151 B.n487 B.n14 585
R152 B.n486 B.n485 585
R153 B.n484 B.n15 585
R154 B.n483 B.n482 585
R155 B.n481 B.n16 585
R156 B.n480 B.n479 585
R157 B.n478 B.n17 585
R158 B.n477 B.n476 585
R159 B.n475 B.n18 585
R160 B.n474 B.n473 585
R161 B.n472 B.n19 585
R162 B.n471 B.n470 585
R163 B.n469 B.n20 585
R164 B.n468 B.n467 585
R165 B.n466 B.n21 585
R166 B.n465 B.n464 585
R167 B.n463 B.n22 585
R168 B.n462 B.n461 585
R169 B.n460 B.n23 585
R170 B.n459 B.n458 585
R171 B.n457 B.n24 585
R172 B.n456 B.n455 585
R173 B.n454 B.n25 585
R174 B.n453 B.n452 585
R175 B.n451 B.n26 585
R176 B.n450 B.n449 585
R177 B.n448 B.n27 585
R178 B.n447 B.n446 585
R179 B.n445 B.n28 585
R180 B.n444 B.n443 585
R181 B.n442 B.n29 585
R182 B.n441 B.n440 585
R183 B.n439 B.n30 585
R184 B.n438 B.n437 585
R185 B.n436 B.n31 585
R186 B.n434 B.n433 585
R187 B.n432 B.n34 585
R188 B.n431 B.n430 585
R189 B.n429 B.n35 585
R190 B.n428 B.n427 585
R191 B.n426 B.n36 585
R192 B.n425 B.n424 585
R193 B.n423 B.n37 585
R194 B.n422 B.n421 585
R195 B.n420 B.n419 585
R196 B.n418 B.n41 585
R197 B.n417 B.n416 585
R198 B.n415 B.n42 585
R199 B.n414 B.n413 585
R200 B.n412 B.n43 585
R201 B.n411 B.n410 585
R202 B.n409 B.n44 585
R203 B.n408 B.n407 585
R204 B.n406 B.n45 585
R205 B.n405 B.n404 585
R206 B.n403 B.n46 585
R207 B.n402 B.n401 585
R208 B.n400 B.n47 585
R209 B.n399 B.n398 585
R210 B.n397 B.n48 585
R211 B.n396 B.n395 585
R212 B.n394 B.n49 585
R213 B.n393 B.n392 585
R214 B.n391 B.n50 585
R215 B.n390 B.n389 585
R216 B.n388 B.n51 585
R217 B.n387 B.n386 585
R218 B.n385 B.n52 585
R219 B.n384 B.n383 585
R220 B.n382 B.n53 585
R221 B.n381 B.n380 585
R222 B.n379 B.n54 585
R223 B.n378 B.n377 585
R224 B.n376 B.n55 585
R225 B.n375 B.n374 585
R226 B.n373 B.n56 585
R227 B.n372 B.n371 585
R228 B.n370 B.n57 585
R229 B.n369 B.n368 585
R230 B.n367 B.n58 585
R231 B.n366 B.n365 585
R232 B.n364 B.n59 585
R233 B.n363 B.n362 585
R234 B.n361 B.n60 585
R235 B.n360 B.n359 585
R236 B.n358 B.n61 585
R237 B.n357 B.n356 585
R238 B.n501 B.n500 585
R239 B.n502 B.n9 585
R240 B.n504 B.n503 585
R241 B.n505 B.n8 585
R242 B.n507 B.n506 585
R243 B.n508 B.n7 585
R244 B.n510 B.n509 585
R245 B.n511 B.n6 585
R246 B.n513 B.n512 585
R247 B.n514 B.n5 585
R248 B.n516 B.n515 585
R249 B.n517 B.n4 585
R250 B.n519 B.n518 585
R251 B.n520 B.n3 585
R252 B.n522 B.n521 585
R253 B.n523 B.n0 585
R254 B.n2 B.n1 585
R255 B.n137 B.n136 585
R256 B.n138 B.n135 585
R257 B.n140 B.n139 585
R258 B.n141 B.n134 585
R259 B.n143 B.n142 585
R260 B.n144 B.n133 585
R261 B.n146 B.n145 585
R262 B.n147 B.n132 585
R263 B.n149 B.n148 585
R264 B.n150 B.n131 585
R265 B.n152 B.n151 585
R266 B.n153 B.n130 585
R267 B.n155 B.n154 585
R268 B.n156 B.n129 585
R269 B.n158 B.n157 585
R270 B.n106 B.t6 478.805
R271 B.n236 B.t0 478.805
R272 B.n38 B.t3 478.805
R273 B.n32 B.t9 478.805
R274 B.n159 B.n158 478.086
R275 B.n306 B.n79 478.086
R276 B.n356 B.n355 478.086
R277 B.n500 B.n499 478.086
R278 B.n525 B.n524 256.663
R279 B.n524 B.n523 235.042
R280 B.n524 B.n2 235.042
R281 B.n160 B.n159 163.367
R282 B.n160 B.n127 163.367
R283 B.n164 B.n127 163.367
R284 B.n165 B.n164 163.367
R285 B.n166 B.n165 163.367
R286 B.n166 B.n125 163.367
R287 B.n170 B.n125 163.367
R288 B.n171 B.n170 163.367
R289 B.n172 B.n171 163.367
R290 B.n172 B.n123 163.367
R291 B.n176 B.n123 163.367
R292 B.n177 B.n176 163.367
R293 B.n178 B.n177 163.367
R294 B.n178 B.n121 163.367
R295 B.n182 B.n121 163.367
R296 B.n183 B.n182 163.367
R297 B.n184 B.n183 163.367
R298 B.n184 B.n119 163.367
R299 B.n188 B.n119 163.367
R300 B.n189 B.n188 163.367
R301 B.n190 B.n189 163.367
R302 B.n190 B.n117 163.367
R303 B.n194 B.n117 163.367
R304 B.n195 B.n194 163.367
R305 B.n196 B.n195 163.367
R306 B.n196 B.n115 163.367
R307 B.n200 B.n115 163.367
R308 B.n201 B.n200 163.367
R309 B.n202 B.n201 163.367
R310 B.n202 B.n113 163.367
R311 B.n206 B.n113 163.367
R312 B.n207 B.n206 163.367
R313 B.n208 B.n207 163.367
R314 B.n208 B.n111 163.367
R315 B.n212 B.n111 163.367
R316 B.n213 B.n212 163.367
R317 B.n214 B.n213 163.367
R318 B.n214 B.n109 163.367
R319 B.n218 B.n109 163.367
R320 B.n219 B.n218 163.367
R321 B.n220 B.n219 163.367
R322 B.n220 B.n105 163.367
R323 B.n225 B.n105 163.367
R324 B.n226 B.n225 163.367
R325 B.n227 B.n226 163.367
R326 B.n227 B.n103 163.367
R327 B.n231 B.n103 163.367
R328 B.n232 B.n231 163.367
R329 B.n233 B.n232 163.367
R330 B.n233 B.n101 163.367
R331 B.n240 B.n101 163.367
R332 B.n241 B.n240 163.367
R333 B.n242 B.n241 163.367
R334 B.n242 B.n99 163.367
R335 B.n246 B.n99 163.367
R336 B.n247 B.n246 163.367
R337 B.n248 B.n247 163.367
R338 B.n248 B.n97 163.367
R339 B.n252 B.n97 163.367
R340 B.n253 B.n252 163.367
R341 B.n254 B.n253 163.367
R342 B.n254 B.n95 163.367
R343 B.n258 B.n95 163.367
R344 B.n259 B.n258 163.367
R345 B.n260 B.n259 163.367
R346 B.n260 B.n93 163.367
R347 B.n264 B.n93 163.367
R348 B.n265 B.n264 163.367
R349 B.n266 B.n265 163.367
R350 B.n266 B.n91 163.367
R351 B.n270 B.n91 163.367
R352 B.n271 B.n270 163.367
R353 B.n272 B.n271 163.367
R354 B.n272 B.n89 163.367
R355 B.n276 B.n89 163.367
R356 B.n277 B.n276 163.367
R357 B.n278 B.n277 163.367
R358 B.n278 B.n87 163.367
R359 B.n282 B.n87 163.367
R360 B.n283 B.n282 163.367
R361 B.n284 B.n283 163.367
R362 B.n284 B.n85 163.367
R363 B.n288 B.n85 163.367
R364 B.n289 B.n288 163.367
R365 B.n290 B.n289 163.367
R366 B.n290 B.n83 163.367
R367 B.n294 B.n83 163.367
R368 B.n295 B.n294 163.367
R369 B.n296 B.n295 163.367
R370 B.n296 B.n81 163.367
R371 B.n300 B.n81 163.367
R372 B.n301 B.n300 163.367
R373 B.n302 B.n301 163.367
R374 B.n302 B.n79 163.367
R375 B.n355 B.n354 163.367
R376 B.n354 B.n63 163.367
R377 B.n350 B.n63 163.367
R378 B.n350 B.n349 163.367
R379 B.n349 B.n348 163.367
R380 B.n348 B.n65 163.367
R381 B.n344 B.n65 163.367
R382 B.n344 B.n343 163.367
R383 B.n343 B.n342 163.367
R384 B.n342 B.n67 163.367
R385 B.n338 B.n67 163.367
R386 B.n338 B.n337 163.367
R387 B.n337 B.n336 163.367
R388 B.n336 B.n69 163.367
R389 B.n332 B.n69 163.367
R390 B.n332 B.n331 163.367
R391 B.n331 B.n330 163.367
R392 B.n330 B.n71 163.367
R393 B.n326 B.n71 163.367
R394 B.n326 B.n325 163.367
R395 B.n325 B.n324 163.367
R396 B.n324 B.n73 163.367
R397 B.n320 B.n73 163.367
R398 B.n320 B.n319 163.367
R399 B.n319 B.n318 163.367
R400 B.n318 B.n75 163.367
R401 B.n314 B.n75 163.367
R402 B.n314 B.n313 163.367
R403 B.n313 B.n312 163.367
R404 B.n312 B.n77 163.367
R405 B.n308 B.n77 163.367
R406 B.n308 B.n307 163.367
R407 B.n307 B.n306 163.367
R408 B.n499 B.n498 163.367
R409 B.n498 B.n11 163.367
R410 B.n494 B.n11 163.367
R411 B.n494 B.n493 163.367
R412 B.n493 B.n492 163.367
R413 B.n492 B.n13 163.367
R414 B.n488 B.n13 163.367
R415 B.n488 B.n487 163.367
R416 B.n487 B.n486 163.367
R417 B.n486 B.n15 163.367
R418 B.n482 B.n15 163.367
R419 B.n482 B.n481 163.367
R420 B.n481 B.n480 163.367
R421 B.n480 B.n17 163.367
R422 B.n476 B.n17 163.367
R423 B.n476 B.n475 163.367
R424 B.n475 B.n474 163.367
R425 B.n474 B.n19 163.367
R426 B.n470 B.n19 163.367
R427 B.n470 B.n469 163.367
R428 B.n469 B.n468 163.367
R429 B.n468 B.n21 163.367
R430 B.n464 B.n21 163.367
R431 B.n464 B.n463 163.367
R432 B.n463 B.n462 163.367
R433 B.n462 B.n23 163.367
R434 B.n458 B.n23 163.367
R435 B.n458 B.n457 163.367
R436 B.n457 B.n456 163.367
R437 B.n456 B.n25 163.367
R438 B.n452 B.n25 163.367
R439 B.n452 B.n451 163.367
R440 B.n451 B.n450 163.367
R441 B.n450 B.n27 163.367
R442 B.n446 B.n27 163.367
R443 B.n446 B.n445 163.367
R444 B.n445 B.n444 163.367
R445 B.n444 B.n29 163.367
R446 B.n440 B.n29 163.367
R447 B.n440 B.n439 163.367
R448 B.n439 B.n438 163.367
R449 B.n438 B.n31 163.367
R450 B.n433 B.n31 163.367
R451 B.n433 B.n432 163.367
R452 B.n432 B.n431 163.367
R453 B.n431 B.n35 163.367
R454 B.n427 B.n35 163.367
R455 B.n427 B.n426 163.367
R456 B.n426 B.n425 163.367
R457 B.n425 B.n37 163.367
R458 B.n421 B.n37 163.367
R459 B.n421 B.n420 163.367
R460 B.n420 B.n41 163.367
R461 B.n416 B.n41 163.367
R462 B.n416 B.n415 163.367
R463 B.n415 B.n414 163.367
R464 B.n414 B.n43 163.367
R465 B.n410 B.n43 163.367
R466 B.n410 B.n409 163.367
R467 B.n409 B.n408 163.367
R468 B.n408 B.n45 163.367
R469 B.n404 B.n45 163.367
R470 B.n404 B.n403 163.367
R471 B.n403 B.n402 163.367
R472 B.n402 B.n47 163.367
R473 B.n398 B.n47 163.367
R474 B.n398 B.n397 163.367
R475 B.n397 B.n396 163.367
R476 B.n396 B.n49 163.367
R477 B.n392 B.n49 163.367
R478 B.n392 B.n391 163.367
R479 B.n391 B.n390 163.367
R480 B.n390 B.n51 163.367
R481 B.n386 B.n51 163.367
R482 B.n386 B.n385 163.367
R483 B.n385 B.n384 163.367
R484 B.n384 B.n53 163.367
R485 B.n380 B.n53 163.367
R486 B.n380 B.n379 163.367
R487 B.n379 B.n378 163.367
R488 B.n378 B.n55 163.367
R489 B.n374 B.n55 163.367
R490 B.n374 B.n373 163.367
R491 B.n373 B.n372 163.367
R492 B.n372 B.n57 163.367
R493 B.n368 B.n57 163.367
R494 B.n368 B.n367 163.367
R495 B.n367 B.n366 163.367
R496 B.n366 B.n59 163.367
R497 B.n362 B.n59 163.367
R498 B.n362 B.n361 163.367
R499 B.n361 B.n360 163.367
R500 B.n360 B.n61 163.367
R501 B.n356 B.n61 163.367
R502 B.n500 B.n9 163.367
R503 B.n504 B.n9 163.367
R504 B.n505 B.n504 163.367
R505 B.n506 B.n505 163.367
R506 B.n506 B.n7 163.367
R507 B.n510 B.n7 163.367
R508 B.n511 B.n510 163.367
R509 B.n512 B.n511 163.367
R510 B.n512 B.n5 163.367
R511 B.n516 B.n5 163.367
R512 B.n517 B.n516 163.367
R513 B.n518 B.n517 163.367
R514 B.n518 B.n3 163.367
R515 B.n522 B.n3 163.367
R516 B.n523 B.n522 163.367
R517 B.n136 B.n2 163.367
R518 B.n136 B.n135 163.367
R519 B.n140 B.n135 163.367
R520 B.n141 B.n140 163.367
R521 B.n142 B.n141 163.367
R522 B.n142 B.n133 163.367
R523 B.n146 B.n133 163.367
R524 B.n147 B.n146 163.367
R525 B.n148 B.n147 163.367
R526 B.n148 B.n131 163.367
R527 B.n152 B.n131 163.367
R528 B.n153 B.n152 163.367
R529 B.n154 B.n153 163.367
R530 B.n154 B.n129 163.367
R531 B.n158 B.n129 163.367
R532 B.n236 B.t1 136.314
R533 B.n38 B.t5 136.314
R534 B.n106 B.t7 136.298
R535 B.n32 B.t11 136.298
R536 B.n237 B.t2 108.969
R537 B.n39 B.t4 108.969
R538 B.n107 B.t8 108.954
R539 B.n33 B.t10 108.954
R540 B.n223 B.n107 59.5399
R541 B.n238 B.n237 59.5399
R542 B.n40 B.n39 59.5399
R543 B.n435 B.n33 59.5399
R544 B.n501 B.n10 31.0639
R545 B.n357 B.n62 31.0639
R546 B.n305 B.n304 31.0639
R547 B.n157 B.n128 31.0639
R548 B.n107 B.n106 27.346
R549 B.n237 B.n236 27.346
R550 B.n39 B.n38 27.346
R551 B.n33 B.n32 27.346
R552 B B.n525 18.0485
R553 B.n502 B.n501 10.6151
R554 B.n503 B.n502 10.6151
R555 B.n503 B.n8 10.6151
R556 B.n507 B.n8 10.6151
R557 B.n508 B.n507 10.6151
R558 B.n509 B.n508 10.6151
R559 B.n509 B.n6 10.6151
R560 B.n513 B.n6 10.6151
R561 B.n514 B.n513 10.6151
R562 B.n515 B.n514 10.6151
R563 B.n515 B.n4 10.6151
R564 B.n519 B.n4 10.6151
R565 B.n520 B.n519 10.6151
R566 B.n521 B.n520 10.6151
R567 B.n521 B.n0 10.6151
R568 B.n497 B.n10 10.6151
R569 B.n497 B.n496 10.6151
R570 B.n496 B.n495 10.6151
R571 B.n495 B.n12 10.6151
R572 B.n491 B.n12 10.6151
R573 B.n491 B.n490 10.6151
R574 B.n490 B.n489 10.6151
R575 B.n489 B.n14 10.6151
R576 B.n485 B.n14 10.6151
R577 B.n485 B.n484 10.6151
R578 B.n484 B.n483 10.6151
R579 B.n483 B.n16 10.6151
R580 B.n479 B.n16 10.6151
R581 B.n479 B.n478 10.6151
R582 B.n478 B.n477 10.6151
R583 B.n477 B.n18 10.6151
R584 B.n473 B.n18 10.6151
R585 B.n473 B.n472 10.6151
R586 B.n472 B.n471 10.6151
R587 B.n471 B.n20 10.6151
R588 B.n467 B.n20 10.6151
R589 B.n467 B.n466 10.6151
R590 B.n466 B.n465 10.6151
R591 B.n465 B.n22 10.6151
R592 B.n461 B.n22 10.6151
R593 B.n461 B.n460 10.6151
R594 B.n460 B.n459 10.6151
R595 B.n459 B.n24 10.6151
R596 B.n455 B.n24 10.6151
R597 B.n455 B.n454 10.6151
R598 B.n454 B.n453 10.6151
R599 B.n453 B.n26 10.6151
R600 B.n449 B.n26 10.6151
R601 B.n449 B.n448 10.6151
R602 B.n448 B.n447 10.6151
R603 B.n447 B.n28 10.6151
R604 B.n443 B.n28 10.6151
R605 B.n443 B.n442 10.6151
R606 B.n442 B.n441 10.6151
R607 B.n441 B.n30 10.6151
R608 B.n437 B.n30 10.6151
R609 B.n437 B.n436 10.6151
R610 B.n434 B.n34 10.6151
R611 B.n430 B.n34 10.6151
R612 B.n430 B.n429 10.6151
R613 B.n429 B.n428 10.6151
R614 B.n428 B.n36 10.6151
R615 B.n424 B.n36 10.6151
R616 B.n424 B.n423 10.6151
R617 B.n423 B.n422 10.6151
R618 B.n419 B.n418 10.6151
R619 B.n418 B.n417 10.6151
R620 B.n417 B.n42 10.6151
R621 B.n413 B.n42 10.6151
R622 B.n413 B.n412 10.6151
R623 B.n412 B.n411 10.6151
R624 B.n411 B.n44 10.6151
R625 B.n407 B.n44 10.6151
R626 B.n407 B.n406 10.6151
R627 B.n406 B.n405 10.6151
R628 B.n405 B.n46 10.6151
R629 B.n401 B.n46 10.6151
R630 B.n401 B.n400 10.6151
R631 B.n400 B.n399 10.6151
R632 B.n399 B.n48 10.6151
R633 B.n395 B.n48 10.6151
R634 B.n395 B.n394 10.6151
R635 B.n394 B.n393 10.6151
R636 B.n393 B.n50 10.6151
R637 B.n389 B.n50 10.6151
R638 B.n389 B.n388 10.6151
R639 B.n388 B.n387 10.6151
R640 B.n387 B.n52 10.6151
R641 B.n383 B.n52 10.6151
R642 B.n383 B.n382 10.6151
R643 B.n382 B.n381 10.6151
R644 B.n381 B.n54 10.6151
R645 B.n377 B.n54 10.6151
R646 B.n377 B.n376 10.6151
R647 B.n376 B.n375 10.6151
R648 B.n375 B.n56 10.6151
R649 B.n371 B.n56 10.6151
R650 B.n371 B.n370 10.6151
R651 B.n370 B.n369 10.6151
R652 B.n369 B.n58 10.6151
R653 B.n365 B.n58 10.6151
R654 B.n365 B.n364 10.6151
R655 B.n364 B.n363 10.6151
R656 B.n363 B.n60 10.6151
R657 B.n359 B.n60 10.6151
R658 B.n359 B.n358 10.6151
R659 B.n358 B.n357 10.6151
R660 B.n353 B.n62 10.6151
R661 B.n353 B.n352 10.6151
R662 B.n352 B.n351 10.6151
R663 B.n351 B.n64 10.6151
R664 B.n347 B.n64 10.6151
R665 B.n347 B.n346 10.6151
R666 B.n346 B.n345 10.6151
R667 B.n345 B.n66 10.6151
R668 B.n341 B.n66 10.6151
R669 B.n341 B.n340 10.6151
R670 B.n340 B.n339 10.6151
R671 B.n339 B.n68 10.6151
R672 B.n335 B.n68 10.6151
R673 B.n335 B.n334 10.6151
R674 B.n334 B.n333 10.6151
R675 B.n333 B.n70 10.6151
R676 B.n329 B.n70 10.6151
R677 B.n329 B.n328 10.6151
R678 B.n328 B.n327 10.6151
R679 B.n327 B.n72 10.6151
R680 B.n323 B.n72 10.6151
R681 B.n323 B.n322 10.6151
R682 B.n322 B.n321 10.6151
R683 B.n321 B.n74 10.6151
R684 B.n317 B.n74 10.6151
R685 B.n317 B.n316 10.6151
R686 B.n316 B.n315 10.6151
R687 B.n315 B.n76 10.6151
R688 B.n311 B.n76 10.6151
R689 B.n311 B.n310 10.6151
R690 B.n310 B.n309 10.6151
R691 B.n309 B.n78 10.6151
R692 B.n305 B.n78 10.6151
R693 B.n137 B.n1 10.6151
R694 B.n138 B.n137 10.6151
R695 B.n139 B.n138 10.6151
R696 B.n139 B.n134 10.6151
R697 B.n143 B.n134 10.6151
R698 B.n144 B.n143 10.6151
R699 B.n145 B.n144 10.6151
R700 B.n145 B.n132 10.6151
R701 B.n149 B.n132 10.6151
R702 B.n150 B.n149 10.6151
R703 B.n151 B.n150 10.6151
R704 B.n151 B.n130 10.6151
R705 B.n155 B.n130 10.6151
R706 B.n156 B.n155 10.6151
R707 B.n157 B.n156 10.6151
R708 B.n161 B.n128 10.6151
R709 B.n162 B.n161 10.6151
R710 B.n163 B.n162 10.6151
R711 B.n163 B.n126 10.6151
R712 B.n167 B.n126 10.6151
R713 B.n168 B.n167 10.6151
R714 B.n169 B.n168 10.6151
R715 B.n169 B.n124 10.6151
R716 B.n173 B.n124 10.6151
R717 B.n174 B.n173 10.6151
R718 B.n175 B.n174 10.6151
R719 B.n175 B.n122 10.6151
R720 B.n179 B.n122 10.6151
R721 B.n180 B.n179 10.6151
R722 B.n181 B.n180 10.6151
R723 B.n181 B.n120 10.6151
R724 B.n185 B.n120 10.6151
R725 B.n186 B.n185 10.6151
R726 B.n187 B.n186 10.6151
R727 B.n187 B.n118 10.6151
R728 B.n191 B.n118 10.6151
R729 B.n192 B.n191 10.6151
R730 B.n193 B.n192 10.6151
R731 B.n193 B.n116 10.6151
R732 B.n197 B.n116 10.6151
R733 B.n198 B.n197 10.6151
R734 B.n199 B.n198 10.6151
R735 B.n199 B.n114 10.6151
R736 B.n203 B.n114 10.6151
R737 B.n204 B.n203 10.6151
R738 B.n205 B.n204 10.6151
R739 B.n205 B.n112 10.6151
R740 B.n209 B.n112 10.6151
R741 B.n210 B.n209 10.6151
R742 B.n211 B.n210 10.6151
R743 B.n211 B.n110 10.6151
R744 B.n215 B.n110 10.6151
R745 B.n216 B.n215 10.6151
R746 B.n217 B.n216 10.6151
R747 B.n217 B.n108 10.6151
R748 B.n221 B.n108 10.6151
R749 B.n222 B.n221 10.6151
R750 B.n224 B.n104 10.6151
R751 B.n228 B.n104 10.6151
R752 B.n229 B.n228 10.6151
R753 B.n230 B.n229 10.6151
R754 B.n230 B.n102 10.6151
R755 B.n234 B.n102 10.6151
R756 B.n235 B.n234 10.6151
R757 B.n239 B.n235 10.6151
R758 B.n243 B.n100 10.6151
R759 B.n244 B.n243 10.6151
R760 B.n245 B.n244 10.6151
R761 B.n245 B.n98 10.6151
R762 B.n249 B.n98 10.6151
R763 B.n250 B.n249 10.6151
R764 B.n251 B.n250 10.6151
R765 B.n251 B.n96 10.6151
R766 B.n255 B.n96 10.6151
R767 B.n256 B.n255 10.6151
R768 B.n257 B.n256 10.6151
R769 B.n257 B.n94 10.6151
R770 B.n261 B.n94 10.6151
R771 B.n262 B.n261 10.6151
R772 B.n263 B.n262 10.6151
R773 B.n263 B.n92 10.6151
R774 B.n267 B.n92 10.6151
R775 B.n268 B.n267 10.6151
R776 B.n269 B.n268 10.6151
R777 B.n269 B.n90 10.6151
R778 B.n273 B.n90 10.6151
R779 B.n274 B.n273 10.6151
R780 B.n275 B.n274 10.6151
R781 B.n275 B.n88 10.6151
R782 B.n279 B.n88 10.6151
R783 B.n280 B.n279 10.6151
R784 B.n281 B.n280 10.6151
R785 B.n281 B.n86 10.6151
R786 B.n285 B.n86 10.6151
R787 B.n286 B.n285 10.6151
R788 B.n287 B.n286 10.6151
R789 B.n287 B.n84 10.6151
R790 B.n291 B.n84 10.6151
R791 B.n292 B.n291 10.6151
R792 B.n293 B.n292 10.6151
R793 B.n293 B.n82 10.6151
R794 B.n297 B.n82 10.6151
R795 B.n298 B.n297 10.6151
R796 B.n299 B.n298 10.6151
R797 B.n299 B.n80 10.6151
R798 B.n303 B.n80 10.6151
R799 B.n304 B.n303 10.6151
R800 B.n525 B.n0 8.11757
R801 B.n525 B.n1 8.11757
R802 B.n435 B.n434 7.18099
R803 B.n422 B.n40 7.18099
R804 B.n224 B.n223 7.18099
R805 B.n239 B.n238 7.18099
R806 B.n436 B.n435 3.43465
R807 B.n419 B.n40 3.43465
R808 B.n223 B.n222 3.43465
R809 B.n238 B.n100 3.43465
R810 VP.n0 VP.t0 513.937
R811 VP.n0 VP.t1 473.038
R812 VP VP.n0 0.0516364
R813 VDD1 VDD1.t0 117.498
R814 VDD1 VDD1.t1 80.285
C0 VN VTAIL 1.88005f
C1 VP VN 4.79405f
C2 B VTAIL 2.99209f
C3 VDD2 VTAIL 5.39113f
C4 w_n1534_n3440# VN 1.98227f
C5 VP B 1.10897f
C6 VP VDD2 0.271181f
C7 w_n1534_n3440# B 7.2667f
C8 w_n1534_n3440# VDD2 1.64587f
C9 VDD1 VN 0.149095f
C10 VDD1 B 1.50702f
C11 VP VTAIL 1.89457f
C12 VDD1 VDD2 0.50054f
C13 w_n1534_n3440# VTAIL 2.91378f
C14 VP w_n1534_n3440# 2.17439f
C15 VN B 0.799203f
C16 VDD2 VN 2.34629f
C17 VDD1 VTAIL 5.35359f
C18 VDD2 B 1.52425f
C19 VDD1 VP 2.46449f
C20 VDD1 w_n1534_n3440# 1.6374f
C21 VDD2 VSUBS 0.784854f
C22 VDD1 VSUBS 4.114768f
C23 VTAIL VSUBS 0.8129f
C24 VN VSUBS 5.49454f
C25 VP VSUBS 1.232226f
C26 B VSUBS 2.803713f
C27 w_n1534_n3440# VSUBS 64.925f
C28 VDD1.t1 VSUBS 2.08302f
C29 VDD1.t0 VSUBS 2.592f
C30 VP.t0 VSUBS 2.39804f
C31 VP.t1 VSUBS 2.19667f
C32 VP.n0 VSUBS 4.87555f
C33 B.n0 VSUBS 0.006192f
C34 B.n1 VSUBS 0.006192f
C35 B.n2 VSUBS 0.009158f
C36 B.n3 VSUBS 0.007018f
C37 B.n4 VSUBS 0.007018f
C38 B.n5 VSUBS 0.007018f
C39 B.n6 VSUBS 0.007018f
C40 B.n7 VSUBS 0.007018f
C41 B.n8 VSUBS 0.007018f
C42 B.n9 VSUBS 0.007018f
C43 B.n10 VSUBS 0.016266f
C44 B.n11 VSUBS 0.007018f
C45 B.n12 VSUBS 0.007018f
C46 B.n13 VSUBS 0.007018f
C47 B.n14 VSUBS 0.007018f
C48 B.n15 VSUBS 0.007018f
C49 B.n16 VSUBS 0.007018f
C50 B.n17 VSUBS 0.007018f
C51 B.n18 VSUBS 0.007018f
C52 B.n19 VSUBS 0.007018f
C53 B.n20 VSUBS 0.007018f
C54 B.n21 VSUBS 0.007018f
C55 B.n22 VSUBS 0.007018f
C56 B.n23 VSUBS 0.007018f
C57 B.n24 VSUBS 0.007018f
C58 B.n25 VSUBS 0.007018f
C59 B.n26 VSUBS 0.007018f
C60 B.n27 VSUBS 0.007018f
C61 B.n28 VSUBS 0.007018f
C62 B.n29 VSUBS 0.007018f
C63 B.n30 VSUBS 0.007018f
C64 B.n31 VSUBS 0.007018f
C65 B.t10 VSUBS 0.404369f
C66 B.t11 VSUBS 0.415541f
C67 B.t9 VSUBS 0.568336f
C68 B.n32 VSUBS 0.164328f
C69 B.n33 VSUBS 0.065696f
C70 B.n34 VSUBS 0.007018f
C71 B.n35 VSUBS 0.007018f
C72 B.n36 VSUBS 0.007018f
C73 B.n37 VSUBS 0.007018f
C74 B.t4 VSUBS 0.40436f
C75 B.t5 VSUBS 0.415533f
C76 B.t3 VSUBS 0.568336f
C77 B.n38 VSUBS 0.164336f
C78 B.n39 VSUBS 0.065704f
C79 B.n40 VSUBS 0.01626f
C80 B.n41 VSUBS 0.007018f
C81 B.n42 VSUBS 0.007018f
C82 B.n43 VSUBS 0.007018f
C83 B.n44 VSUBS 0.007018f
C84 B.n45 VSUBS 0.007018f
C85 B.n46 VSUBS 0.007018f
C86 B.n47 VSUBS 0.007018f
C87 B.n48 VSUBS 0.007018f
C88 B.n49 VSUBS 0.007018f
C89 B.n50 VSUBS 0.007018f
C90 B.n51 VSUBS 0.007018f
C91 B.n52 VSUBS 0.007018f
C92 B.n53 VSUBS 0.007018f
C93 B.n54 VSUBS 0.007018f
C94 B.n55 VSUBS 0.007018f
C95 B.n56 VSUBS 0.007018f
C96 B.n57 VSUBS 0.007018f
C97 B.n58 VSUBS 0.007018f
C98 B.n59 VSUBS 0.007018f
C99 B.n60 VSUBS 0.007018f
C100 B.n61 VSUBS 0.007018f
C101 B.n62 VSUBS 0.015522f
C102 B.n63 VSUBS 0.007018f
C103 B.n64 VSUBS 0.007018f
C104 B.n65 VSUBS 0.007018f
C105 B.n66 VSUBS 0.007018f
C106 B.n67 VSUBS 0.007018f
C107 B.n68 VSUBS 0.007018f
C108 B.n69 VSUBS 0.007018f
C109 B.n70 VSUBS 0.007018f
C110 B.n71 VSUBS 0.007018f
C111 B.n72 VSUBS 0.007018f
C112 B.n73 VSUBS 0.007018f
C113 B.n74 VSUBS 0.007018f
C114 B.n75 VSUBS 0.007018f
C115 B.n76 VSUBS 0.007018f
C116 B.n77 VSUBS 0.007018f
C117 B.n78 VSUBS 0.007018f
C118 B.n79 VSUBS 0.016266f
C119 B.n80 VSUBS 0.007018f
C120 B.n81 VSUBS 0.007018f
C121 B.n82 VSUBS 0.007018f
C122 B.n83 VSUBS 0.007018f
C123 B.n84 VSUBS 0.007018f
C124 B.n85 VSUBS 0.007018f
C125 B.n86 VSUBS 0.007018f
C126 B.n87 VSUBS 0.007018f
C127 B.n88 VSUBS 0.007018f
C128 B.n89 VSUBS 0.007018f
C129 B.n90 VSUBS 0.007018f
C130 B.n91 VSUBS 0.007018f
C131 B.n92 VSUBS 0.007018f
C132 B.n93 VSUBS 0.007018f
C133 B.n94 VSUBS 0.007018f
C134 B.n95 VSUBS 0.007018f
C135 B.n96 VSUBS 0.007018f
C136 B.n97 VSUBS 0.007018f
C137 B.n98 VSUBS 0.007018f
C138 B.n99 VSUBS 0.007018f
C139 B.n100 VSUBS 0.004644f
C140 B.n101 VSUBS 0.007018f
C141 B.n102 VSUBS 0.007018f
C142 B.n103 VSUBS 0.007018f
C143 B.n104 VSUBS 0.007018f
C144 B.n105 VSUBS 0.007018f
C145 B.t8 VSUBS 0.404369f
C146 B.t7 VSUBS 0.415541f
C147 B.t6 VSUBS 0.568336f
C148 B.n106 VSUBS 0.164328f
C149 B.n107 VSUBS 0.065696f
C150 B.n108 VSUBS 0.007018f
C151 B.n109 VSUBS 0.007018f
C152 B.n110 VSUBS 0.007018f
C153 B.n111 VSUBS 0.007018f
C154 B.n112 VSUBS 0.007018f
C155 B.n113 VSUBS 0.007018f
C156 B.n114 VSUBS 0.007018f
C157 B.n115 VSUBS 0.007018f
C158 B.n116 VSUBS 0.007018f
C159 B.n117 VSUBS 0.007018f
C160 B.n118 VSUBS 0.007018f
C161 B.n119 VSUBS 0.007018f
C162 B.n120 VSUBS 0.007018f
C163 B.n121 VSUBS 0.007018f
C164 B.n122 VSUBS 0.007018f
C165 B.n123 VSUBS 0.007018f
C166 B.n124 VSUBS 0.007018f
C167 B.n125 VSUBS 0.007018f
C168 B.n126 VSUBS 0.007018f
C169 B.n127 VSUBS 0.007018f
C170 B.n128 VSUBS 0.016266f
C171 B.n129 VSUBS 0.007018f
C172 B.n130 VSUBS 0.007018f
C173 B.n131 VSUBS 0.007018f
C174 B.n132 VSUBS 0.007018f
C175 B.n133 VSUBS 0.007018f
C176 B.n134 VSUBS 0.007018f
C177 B.n135 VSUBS 0.007018f
C178 B.n136 VSUBS 0.007018f
C179 B.n137 VSUBS 0.007018f
C180 B.n138 VSUBS 0.007018f
C181 B.n139 VSUBS 0.007018f
C182 B.n140 VSUBS 0.007018f
C183 B.n141 VSUBS 0.007018f
C184 B.n142 VSUBS 0.007018f
C185 B.n143 VSUBS 0.007018f
C186 B.n144 VSUBS 0.007018f
C187 B.n145 VSUBS 0.007018f
C188 B.n146 VSUBS 0.007018f
C189 B.n147 VSUBS 0.007018f
C190 B.n148 VSUBS 0.007018f
C191 B.n149 VSUBS 0.007018f
C192 B.n150 VSUBS 0.007018f
C193 B.n151 VSUBS 0.007018f
C194 B.n152 VSUBS 0.007018f
C195 B.n153 VSUBS 0.007018f
C196 B.n154 VSUBS 0.007018f
C197 B.n155 VSUBS 0.007018f
C198 B.n156 VSUBS 0.007018f
C199 B.n157 VSUBS 0.015522f
C200 B.n158 VSUBS 0.015522f
C201 B.n159 VSUBS 0.016266f
C202 B.n160 VSUBS 0.007018f
C203 B.n161 VSUBS 0.007018f
C204 B.n162 VSUBS 0.007018f
C205 B.n163 VSUBS 0.007018f
C206 B.n164 VSUBS 0.007018f
C207 B.n165 VSUBS 0.007018f
C208 B.n166 VSUBS 0.007018f
C209 B.n167 VSUBS 0.007018f
C210 B.n168 VSUBS 0.007018f
C211 B.n169 VSUBS 0.007018f
C212 B.n170 VSUBS 0.007018f
C213 B.n171 VSUBS 0.007018f
C214 B.n172 VSUBS 0.007018f
C215 B.n173 VSUBS 0.007018f
C216 B.n174 VSUBS 0.007018f
C217 B.n175 VSUBS 0.007018f
C218 B.n176 VSUBS 0.007018f
C219 B.n177 VSUBS 0.007018f
C220 B.n178 VSUBS 0.007018f
C221 B.n179 VSUBS 0.007018f
C222 B.n180 VSUBS 0.007018f
C223 B.n181 VSUBS 0.007018f
C224 B.n182 VSUBS 0.007018f
C225 B.n183 VSUBS 0.007018f
C226 B.n184 VSUBS 0.007018f
C227 B.n185 VSUBS 0.007018f
C228 B.n186 VSUBS 0.007018f
C229 B.n187 VSUBS 0.007018f
C230 B.n188 VSUBS 0.007018f
C231 B.n189 VSUBS 0.007018f
C232 B.n190 VSUBS 0.007018f
C233 B.n191 VSUBS 0.007018f
C234 B.n192 VSUBS 0.007018f
C235 B.n193 VSUBS 0.007018f
C236 B.n194 VSUBS 0.007018f
C237 B.n195 VSUBS 0.007018f
C238 B.n196 VSUBS 0.007018f
C239 B.n197 VSUBS 0.007018f
C240 B.n198 VSUBS 0.007018f
C241 B.n199 VSUBS 0.007018f
C242 B.n200 VSUBS 0.007018f
C243 B.n201 VSUBS 0.007018f
C244 B.n202 VSUBS 0.007018f
C245 B.n203 VSUBS 0.007018f
C246 B.n204 VSUBS 0.007018f
C247 B.n205 VSUBS 0.007018f
C248 B.n206 VSUBS 0.007018f
C249 B.n207 VSUBS 0.007018f
C250 B.n208 VSUBS 0.007018f
C251 B.n209 VSUBS 0.007018f
C252 B.n210 VSUBS 0.007018f
C253 B.n211 VSUBS 0.007018f
C254 B.n212 VSUBS 0.007018f
C255 B.n213 VSUBS 0.007018f
C256 B.n214 VSUBS 0.007018f
C257 B.n215 VSUBS 0.007018f
C258 B.n216 VSUBS 0.007018f
C259 B.n217 VSUBS 0.007018f
C260 B.n218 VSUBS 0.007018f
C261 B.n219 VSUBS 0.007018f
C262 B.n220 VSUBS 0.007018f
C263 B.n221 VSUBS 0.007018f
C264 B.n222 VSUBS 0.004644f
C265 B.n223 VSUBS 0.01626f
C266 B.n224 VSUBS 0.005883f
C267 B.n225 VSUBS 0.007018f
C268 B.n226 VSUBS 0.007018f
C269 B.n227 VSUBS 0.007018f
C270 B.n228 VSUBS 0.007018f
C271 B.n229 VSUBS 0.007018f
C272 B.n230 VSUBS 0.007018f
C273 B.n231 VSUBS 0.007018f
C274 B.n232 VSUBS 0.007018f
C275 B.n233 VSUBS 0.007018f
C276 B.n234 VSUBS 0.007018f
C277 B.n235 VSUBS 0.007018f
C278 B.t2 VSUBS 0.40436f
C279 B.t1 VSUBS 0.415533f
C280 B.t0 VSUBS 0.568336f
C281 B.n236 VSUBS 0.164336f
C282 B.n237 VSUBS 0.065704f
C283 B.n238 VSUBS 0.01626f
C284 B.n239 VSUBS 0.005883f
C285 B.n240 VSUBS 0.007018f
C286 B.n241 VSUBS 0.007018f
C287 B.n242 VSUBS 0.007018f
C288 B.n243 VSUBS 0.007018f
C289 B.n244 VSUBS 0.007018f
C290 B.n245 VSUBS 0.007018f
C291 B.n246 VSUBS 0.007018f
C292 B.n247 VSUBS 0.007018f
C293 B.n248 VSUBS 0.007018f
C294 B.n249 VSUBS 0.007018f
C295 B.n250 VSUBS 0.007018f
C296 B.n251 VSUBS 0.007018f
C297 B.n252 VSUBS 0.007018f
C298 B.n253 VSUBS 0.007018f
C299 B.n254 VSUBS 0.007018f
C300 B.n255 VSUBS 0.007018f
C301 B.n256 VSUBS 0.007018f
C302 B.n257 VSUBS 0.007018f
C303 B.n258 VSUBS 0.007018f
C304 B.n259 VSUBS 0.007018f
C305 B.n260 VSUBS 0.007018f
C306 B.n261 VSUBS 0.007018f
C307 B.n262 VSUBS 0.007018f
C308 B.n263 VSUBS 0.007018f
C309 B.n264 VSUBS 0.007018f
C310 B.n265 VSUBS 0.007018f
C311 B.n266 VSUBS 0.007018f
C312 B.n267 VSUBS 0.007018f
C313 B.n268 VSUBS 0.007018f
C314 B.n269 VSUBS 0.007018f
C315 B.n270 VSUBS 0.007018f
C316 B.n271 VSUBS 0.007018f
C317 B.n272 VSUBS 0.007018f
C318 B.n273 VSUBS 0.007018f
C319 B.n274 VSUBS 0.007018f
C320 B.n275 VSUBS 0.007018f
C321 B.n276 VSUBS 0.007018f
C322 B.n277 VSUBS 0.007018f
C323 B.n278 VSUBS 0.007018f
C324 B.n279 VSUBS 0.007018f
C325 B.n280 VSUBS 0.007018f
C326 B.n281 VSUBS 0.007018f
C327 B.n282 VSUBS 0.007018f
C328 B.n283 VSUBS 0.007018f
C329 B.n284 VSUBS 0.007018f
C330 B.n285 VSUBS 0.007018f
C331 B.n286 VSUBS 0.007018f
C332 B.n287 VSUBS 0.007018f
C333 B.n288 VSUBS 0.007018f
C334 B.n289 VSUBS 0.007018f
C335 B.n290 VSUBS 0.007018f
C336 B.n291 VSUBS 0.007018f
C337 B.n292 VSUBS 0.007018f
C338 B.n293 VSUBS 0.007018f
C339 B.n294 VSUBS 0.007018f
C340 B.n295 VSUBS 0.007018f
C341 B.n296 VSUBS 0.007018f
C342 B.n297 VSUBS 0.007018f
C343 B.n298 VSUBS 0.007018f
C344 B.n299 VSUBS 0.007018f
C345 B.n300 VSUBS 0.007018f
C346 B.n301 VSUBS 0.007018f
C347 B.n302 VSUBS 0.007018f
C348 B.n303 VSUBS 0.007018f
C349 B.n304 VSUBS 0.015394f
C350 B.n305 VSUBS 0.016393f
C351 B.n306 VSUBS 0.015522f
C352 B.n307 VSUBS 0.007018f
C353 B.n308 VSUBS 0.007018f
C354 B.n309 VSUBS 0.007018f
C355 B.n310 VSUBS 0.007018f
C356 B.n311 VSUBS 0.007018f
C357 B.n312 VSUBS 0.007018f
C358 B.n313 VSUBS 0.007018f
C359 B.n314 VSUBS 0.007018f
C360 B.n315 VSUBS 0.007018f
C361 B.n316 VSUBS 0.007018f
C362 B.n317 VSUBS 0.007018f
C363 B.n318 VSUBS 0.007018f
C364 B.n319 VSUBS 0.007018f
C365 B.n320 VSUBS 0.007018f
C366 B.n321 VSUBS 0.007018f
C367 B.n322 VSUBS 0.007018f
C368 B.n323 VSUBS 0.007018f
C369 B.n324 VSUBS 0.007018f
C370 B.n325 VSUBS 0.007018f
C371 B.n326 VSUBS 0.007018f
C372 B.n327 VSUBS 0.007018f
C373 B.n328 VSUBS 0.007018f
C374 B.n329 VSUBS 0.007018f
C375 B.n330 VSUBS 0.007018f
C376 B.n331 VSUBS 0.007018f
C377 B.n332 VSUBS 0.007018f
C378 B.n333 VSUBS 0.007018f
C379 B.n334 VSUBS 0.007018f
C380 B.n335 VSUBS 0.007018f
C381 B.n336 VSUBS 0.007018f
C382 B.n337 VSUBS 0.007018f
C383 B.n338 VSUBS 0.007018f
C384 B.n339 VSUBS 0.007018f
C385 B.n340 VSUBS 0.007018f
C386 B.n341 VSUBS 0.007018f
C387 B.n342 VSUBS 0.007018f
C388 B.n343 VSUBS 0.007018f
C389 B.n344 VSUBS 0.007018f
C390 B.n345 VSUBS 0.007018f
C391 B.n346 VSUBS 0.007018f
C392 B.n347 VSUBS 0.007018f
C393 B.n348 VSUBS 0.007018f
C394 B.n349 VSUBS 0.007018f
C395 B.n350 VSUBS 0.007018f
C396 B.n351 VSUBS 0.007018f
C397 B.n352 VSUBS 0.007018f
C398 B.n353 VSUBS 0.007018f
C399 B.n354 VSUBS 0.007018f
C400 B.n355 VSUBS 0.015522f
C401 B.n356 VSUBS 0.016266f
C402 B.n357 VSUBS 0.016266f
C403 B.n358 VSUBS 0.007018f
C404 B.n359 VSUBS 0.007018f
C405 B.n360 VSUBS 0.007018f
C406 B.n361 VSUBS 0.007018f
C407 B.n362 VSUBS 0.007018f
C408 B.n363 VSUBS 0.007018f
C409 B.n364 VSUBS 0.007018f
C410 B.n365 VSUBS 0.007018f
C411 B.n366 VSUBS 0.007018f
C412 B.n367 VSUBS 0.007018f
C413 B.n368 VSUBS 0.007018f
C414 B.n369 VSUBS 0.007018f
C415 B.n370 VSUBS 0.007018f
C416 B.n371 VSUBS 0.007018f
C417 B.n372 VSUBS 0.007018f
C418 B.n373 VSUBS 0.007018f
C419 B.n374 VSUBS 0.007018f
C420 B.n375 VSUBS 0.007018f
C421 B.n376 VSUBS 0.007018f
C422 B.n377 VSUBS 0.007018f
C423 B.n378 VSUBS 0.007018f
C424 B.n379 VSUBS 0.007018f
C425 B.n380 VSUBS 0.007018f
C426 B.n381 VSUBS 0.007018f
C427 B.n382 VSUBS 0.007018f
C428 B.n383 VSUBS 0.007018f
C429 B.n384 VSUBS 0.007018f
C430 B.n385 VSUBS 0.007018f
C431 B.n386 VSUBS 0.007018f
C432 B.n387 VSUBS 0.007018f
C433 B.n388 VSUBS 0.007018f
C434 B.n389 VSUBS 0.007018f
C435 B.n390 VSUBS 0.007018f
C436 B.n391 VSUBS 0.007018f
C437 B.n392 VSUBS 0.007018f
C438 B.n393 VSUBS 0.007018f
C439 B.n394 VSUBS 0.007018f
C440 B.n395 VSUBS 0.007018f
C441 B.n396 VSUBS 0.007018f
C442 B.n397 VSUBS 0.007018f
C443 B.n398 VSUBS 0.007018f
C444 B.n399 VSUBS 0.007018f
C445 B.n400 VSUBS 0.007018f
C446 B.n401 VSUBS 0.007018f
C447 B.n402 VSUBS 0.007018f
C448 B.n403 VSUBS 0.007018f
C449 B.n404 VSUBS 0.007018f
C450 B.n405 VSUBS 0.007018f
C451 B.n406 VSUBS 0.007018f
C452 B.n407 VSUBS 0.007018f
C453 B.n408 VSUBS 0.007018f
C454 B.n409 VSUBS 0.007018f
C455 B.n410 VSUBS 0.007018f
C456 B.n411 VSUBS 0.007018f
C457 B.n412 VSUBS 0.007018f
C458 B.n413 VSUBS 0.007018f
C459 B.n414 VSUBS 0.007018f
C460 B.n415 VSUBS 0.007018f
C461 B.n416 VSUBS 0.007018f
C462 B.n417 VSUBS 0.007018f
C463 B.n418 VSUBS 0.007018f
C464 B.n419 VSUBS 0.004644f
C465 B.n420 VSUBS 0.007018f
C466 B.n421 VSUBS 0.007018f
C467 B.n422 VSUBS 0.005883f
C468 B.n423 VSUBS 0.007018f
C469 B.n424 VSUBS 0.007018f
C470 B.n425 VSUBS 0.007018f
C471 B.n426 VSUBS 0.007018f
C472 B.n427 VSUBS 0.007018f
C473 B.n428 VSUBS 0.007018f
C474 B.n429 VSUBS 0.007018f
C475 B.n430 VSUBS 0.007018f
C476 B.n431 VSUBS 0.007018f
C477 B.n432 VSUBS 0.007018f
C478 B.n433 VSUBS 0.007018f
C479 B.n434 VSUBS 0.005883f
C480 B.n435 VSUBS 0.01626f
C481 B.n436 VSUBS 0.004644f
C482 B.n437 VSUBS 0.007018f
C483 B.n438 VSUBS 0.007018f
C484 B.n439 VSUBS 0.007018f
C485 B.n440 VSUBS 0.007018f
C486 B.n441 VSUBS 0.007018f
C487 B.n442 VSUBS 0.007018f
C488 B.n443 VSUBS 0.007018f
C489 B.n444 VSUBS 0.007018f
C490 B.n445 VSUBS 0.007018f
C491 B.n446 VSUBS 0.007018f
C492 B.n447 VSUBS 0.007018f
C493 B.n448 VSUBS 0.007018f
C494 B.n449 VSUBS 0.007018f
C495 B.n450 VSUBS 0.007018f
C496 B.n451 VSUBS 0.007018f
C497 B.n452 VSUBS 0.007018f
C498 B.n453 VSUBS 0.007018f
C499 B.n454 VSUBS 0.007018f
C500 B.n455 VSUBS 0.007018f
C501 B.n456 VSUBS 0.007018f
C502 B.n457 VSUBS 0.007018f
C503 B.n458 VSUBS 0.007018f
C504 B.n459 VSUBS 0.007018f
C505 B.n460 VSUBS 0.007018f
C506 B.n461 VSUBS 0.007018f
C507 B.n462 VSUBS 0.007018f
C508 B.n463 VSUBS 0.007018f
C509 B.n464 VSUBS 0.007018f
C510 B.n465 VSUBS 0.007018f
C511 B.n466 VSUBS 0.007018f
C512 B.n467 VSUBS 0.007018f
C513 B.n468 VSUBS 0.007018f
C514 B.n469 VSUBS 0.007018f
C515 B.n470 VSUBS 0.007018f
C516 B.n471 VSUBS 0.007018f
C517 B.n472 VSUBS 0.007018f
C518 B.n473 VSUBS 0.007018f
C519 B.n474 VSUBS 0.007018f
C520 B.n475 VSUBS 0.007018f
C521 B.n476 VSUBS 0.007018f
C522 B.n477 VSUBS 0.007018f
C523 B.n478 VSUBS 0.007018f
C524 B.n479 VSUBS 0.007018f
C525 B.n480 VSUBS 0.007018f
C526 B.n481 VSUBS 0.007018f
C527 B.n482 VSUBS 0.007018f
C528 B.n483 VSUBS 0.007018f
C529 B.n484 VSUBS 0.007018f
C530 B.n485 VSUBS 0.007018f
C531 B.n486 VSUBS 0.007018f
C532 B.n487 VSUBS 0.007018f
C533 B.n488 VSUBS 0.007018f
C534 B.n489 VSUBS 0.007018f
C535 B.n490 VSUBS 0.007018f
C536 B.n491 VSUBS 0.007018f
C537 B.n492 VSUBS 0.007018f
C538 B.n493 VSUBS 0.007018f
C539 B.n494 VSUBS 0.007018f
C540 B.n495 VSUBS 0.007018f
C541 B.n496 VSUBS 0.007018f
C542 B.n497 VSUBS 0.007018f
C543 B.n498 VSUBS 0.007018f
C544 B.n499 VSUBS 0.016266f
C545 B.n500 VSUBS 0.015522f
C546 B.n501 VSUBS 0.015522f
C547 B.n502 VSUBS 0.007018f
C548 B.n503 VSUBS 0.007018f
C549 B.n504 VSUBS 0.007018f
C550 B.n505 VSUBS 0.007018f
C551 B.n506 VSUBS 0.007018f
C552 B.n507 VSUBS 0.007018f
C553 B.n508 VSUBS 0.007018f
C554 B.n509 VSUBS 0.007018f
C555 B.n510 VSUBS 0.007018f
C556 B.n511 VSUBS 0.007018f
C557 B.n512 VSUBS 0.007018f
C558 B.n513 VSUBS 0.007018f
C559 B.n514 VSUBS 0.007018f
C560 B.n515 VSUBS 0.007018f
C561 B.n516 VSUBS 0.007018f
C562 B.n517 VSUBS 0.007018f
C563 B.n518 VSUBS 0.007018f
C564 B.n519 VSUBS 0.007018f
C565 B.n520 VSUBS 0.007018f
C566 B.n521 VSUBS 0.007018f
C567 B.n522 VSUBS 0.007018f
C568 B.n523 VSUBS 0.009158f
C569 B.n524 VSUBS 0.009756f
C570 B.n525 VSUBS 0.0194f
C571 VDD2.t1 VSUBS 2.52634f
C572 VDD2.t0 VSUBS 2.04798f
C573 VDD2.n0 VSUBS 3.06169f
C574 VTAIL.t0 VSUBS 2.24025f
C575 VTAIL.n0 VSUBS 1.96214f
C576 VTAIL.t3 VSUBS 2.24025f
C577 VTAIL.n1 VSUBS 1.98072f
C578 VTAIL.t1 VSUBS 2.24024f
C579 VTAIL.n2 VSUBS 1.88878f
C580 VTAIL.t2 VSUBS 2.24025f
C581 VTAIL.n3 VSUBS 1.82584f
C582 VN.t0 VSUBS 1.62945f
C583 VN.t1 VSUBS 1.78206f
.ends

