* NGSPICE file created from diff_pair_sample_0026.ext - technology: sky130A

.subckt diff_pair_sample_0026 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2936 pd=8.17 as=3.0576 ps=16.46 w=7.84 l=1.47
X1 VTAIL.t4 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=1.2936 ps=8.17 w=7.84 l=1.47
X2 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=0 ps=0 w=7.84 l=1.47
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=0 ps=0 w=7.84 l=1.47
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=0 ps=0 w=7.84 l=1.47
X5 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=1.2936 ps=8.17 w=7.84 l=1.47
X6 VDD1.t1 VP.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2936 pd=8.17 as=3.0576 ps=16.46 w=7.84 l=1.47
X7 VTAIL.t5 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=1.2936 ps=8.17 w=7.84 l=1.47
X8 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=1.2936 ps=8.17 w=7.84 l=1.47
X9 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2936 pd=8.17 as=3.0576 ps=16.46 w=7.84 l=1.47
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.0576 pd=16.46 as=0 ps=0 w=7.84 l=1.47
X11 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2936 pd=8.17 as=3.0576 ps=16.46 w=7.84 l=1.47
R0 VP.n4 VP.n3 178.514
R1 VP.n12 VP.n11 178.514
R2 VP.n2 VP.t3 164.535
R3 VP.n2 VP.t0 164.22
R4 VP.n10 VP.n0 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n1 161.3
R7 VP.n6 VP.n5 161.3
R8 VP.n4 VP.t1 128.534
R9 VP.n11 VP.t2 128.534
R10 VP.n9 VP.n1 56.5617
R11 VP.n3 VP.n2 52.7045
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 7.37805
R15 VP.n11 VP.n10 7.37805
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VTAIL.n330 VTAIL.n294 289.615
R23 VTAIL.n36 VTAIL.n0 289.615
R24 VTAIL.n78 VTAIL.n42 289.615
R25 VTAIL.n120 VTAIL.n84 289.615
R26 VTAIL.n288 VTAIL.n252 289.615
R27 VTAIL.n246 VTAIL.n210 289.615
R28 VTAIL.n204 VTAIL.n168 289.615
R29 VTAIL.n162 VTAIL.n126 289.615
R30 VTAIL.n306 VTAIL.n305 185
R31 VTAIL.n311 VTAIL.n310 185
R32 VTAIL.n313 VTAIL.n312 185
R33 VTAIL.n302 VTAIL.n301 185
R34 VTAIL.n319 VTAIL.n318 185
R35 VTAIL.n321 VTAIL.n320 185
R36 VTAIL.n298 VTAIL.n297 185
R37 VTAIL.n328 VTAIL.n327 185
R38 VTAIL.n329 VTAIL.n296 185
R39 VTAIL.n331 VTAIL.n330 185
R40 VTAIL.n12 VTAIL.n11 185
R41 VTAIL.n17 VTAIL.n16 185
R42 VTAIL.n19 VTAIL.n18 185
R43 VTAIL.n8 VTAIL.n7 185
R44 VTAIL.n25 VTAIL.n24 185
R45 VTAIL.n27 VTAIL.n26 185
R46 VTAIL.n4 VTAIL.n3 185
R47 VTAIL.n34 VTAIL.n33 185
R48 VTAIL.n35 VTAIL.n2 185
R49 VTAIL.n37 VTAIL.n36 185
R50 VTAIL.n54 VTAIL.n53 185
R51 VTAIL.n59 VTAIL.n58 185
R52 VTAIL.n61 VTAIL.n60 185
R53 VTAIL.n50 VTAIL.n49 185
R54 VTAIL.n67 VTAIL.n66 185
R55 VTAIL.n69 VTAIL.n68 185
R56 VTAIL.n46 VTAIL.n45 185
R57 VTAIL.n76 VTAIL.n75 185
R58 VTAIL.n77 VTAIL.n44 185
R59 VTAIL.n79 VTAIL.n78 185
R60 VTAIL.n96 VTAIL.n95 185
R61 VTAIL.n101 VTAIL.n100 185
R62 VTAIL.n103 VTAIL.n102 185
R63 VTAIL.n92 VTAIL.n91 185
R64 VTAIL.n109 VTAIL.n108 185
R65 VTAIL.n111 VTAIL.n110 185
R66 VTAIL.n88 VTAIL.n87 185
R67 VTAIL.n118 VTAIL.n117 185
R68 VTAIL.n119 VTAIL.n86 185
R69 VTAIL.n121 VTAIL.n120 185
R70 VTAIL.n289 VTAIL.n288 185
R71 VTAIL.n287 VTAIL.n254 185
R72 VTAIL.n286 VTAIL.n285 185
R73 VTAIL.n257 VTAIL.n255 185
R74 VTAIL.n280 VTAIL.n279 185
R75 VTAIL.n278 VTAIL.n277 185
R76 VTAIL.n261 VTAIL.n260 185
R77 VTAIL.n272 VTAIL.n271 185
R78 VTAIL.n270 VTAIL.n269 185
R79 VTAIL.n265 VTAIL.n264 185
R80 VTAIL.n247 VTAIL.n246 185
R81 VTAIL.n245 VTAIL.n212 185
R82 VTAIL.n244 VTAIL.n243 185
R83 VTAIL.n215 VTAIL.n213 185
R84 VTAIL.n238 VTAIL.n237 185
R85 VTAIL.n236 VTAIL.n235 185
R86 VTAIL.n219 VTAIL.n218 185
R87 VTAIL.n230 VTAIL.n229 185
R88 VTAIL.n228 VTAIL.n227 185
R89 VTAIL.n223 VTAIL.n222 185
R90 VTAIL.n205 VTAIL.n204 185
R91 VTAIL.n203 VTAIL.n170 185
R92 VTAIL.n202 VTAIL.n201 185
R93 VTAIL.n173 VTAIL.n171 185
R94 VTAIL.n196 VTAIL.n195 185
R95 VTAIL.n194 VTAIL.n193 185
R96 VTAIL.n177 VTAIL.n176 185
R97 VTAIL.n188 VTAIL.n187 185
R98 VTAIL.n186 VTAIL.n185 185
R99 VTAIL.n181 VTAIL.n180 185
R100 VTAIL.n163 VTAIL.n162 185
R101 VTAIL.n161 VTAIL.n128 185
R102 VTAIL.n160 VTAIL.n159 185
R103 VTAIL.n131 VTAIL.n129 185
R104 VTAIL.n154 VTAIL.n153 185
R105 VTAIL.n152 VTAIL.n151 185
R106 VTAIL.n135 VTAIL.n134 185
R107 VTAIL.n146 VTAIL.n145 185
R108 VTAIL.n144 VTAIL.n143 185
R109 VTAIL.n139 VTAIL.n138 185
R110 VTAIL.n307 VTAIL.t1 149.524
R111 VTAIL.n13 VTAIL.t3 149.524
R112 VTAIL.n55 VTAIL.t6 149.524
R113 VTAIL.n97 VTAIL.t4 149.524
R114 VTAIL.n266 VTAIL.t7 149.524
R115 VTAIL.n224 VTAIL.t5 149.524
R116 VTAIL.n182 VTAIL.t0 149.524
R117 VTAIL.n140 VTAIL.t2 149.524
R118 VTAIL.n311 VTAIL.n305 104.615
R119 VTAIL.n312 VTAIL.n311 104.615
R120 VTAIL.n312 VTAIL.n301 104.615
R121 VTAIL.n319 VTAIL.n301 104.615
R122 VTAIL.n320 VTAIL.n319 104.615
R123 VTAIL.n320 VTAIL.n297 104.615
R124 VTAIL.n328 VTAIL.n297 104.615
R125 VTAIL.n329 VTAIL.n328 104.615
R126 VTAIL.n330 VTAIL.n329 104.615
R127 VTAIL.n17 VTAIL.n11 104.615
R128 VTAIL.n18 VTAIL.n17 104.615
R129 VTAIL.n18 VTAIL.n7 104.615
R130 VTAIL.n25 VTAIL.n7 104.615
R131 VTAIL.n26 VTAIL.n25 104.615
R132 VTAIL.n26 VTAIL.n3 104.615
R133 VTAIL.n34 VTAIL.n3 104.615
R134 VTAIL.n35 VTAIL.n34 104.615
R135 VTAIL.n36 VTAIL.n35 104.615
R136 VTAIL.n59 VTAIL.n53 104.615
R137 VTAIL.n60 VTAIL.n59 104.615
R138 VTAIL.n60 VTAIL.n49 104.615
R139 VTAIL.n67 VTAIL.n49 104.615
R140 VTAIL.n68 VTAIL.n67 104.615
R141 VTAIL.n68 VTAIL.n45 104.615
R142 VTAIL.n76 VTAIL.n45 104.615
R143 VTAIL.n77 VTAIL.n76 104.615
R144 VTAIL.n78 VTAIL.n77 104.615
R145 VTAIL.n101 VTAIL.n95 104.615
R146 VTAIL.n102 VTAIL.n101 104.615
R147 VTAIL.n102 VTAIL.n91 104.615
R148 VTAIL.n109 VTAIL.n91 104.615
R149 VTAIL.n110 VTAIL.n109 104.615
R150 VTAIL.n110 VTAIL.n87 104.615
R151 VTAIL.n118 VTAIL.n87 104.615
R152 VTAIL.n119 VTAIL.n118 104.615
R153 VTAIL.n120 VTAIL.n119 104.615
R154 VTAIL.n288 VTAIL.n287 104.615
R155 VTAIL.n287 VTAIL.n286 104.615
R156 VTAIL.n286 VTAIL.n255 104.615
R157 VTAIL.n279 VTAIL.n255 104.615
R158 VTAIL.n279 VTAIL.n278 104.615
R159 VTAIL.n278 VTAIL.n260 104.615
R160 VTAIL.n271 VTAIL.n260 104.615
R161 VTAIL.n271 VTAIL.n270 104.615
R162 VTAIL.n270 VTAIL.n264 104.615
R163 VTAIL.n246 VTAIL.n245 104.615
R164 VTAIL.n245 VTAIL.n244 104.615
R165 VTAIL.n244 VTAIL.n213 104.615
R166 VTAIL.n237 VTAIL.n213 104.615
R167 VTAIL.n237 VTAIL.n236 104.615
R168 VTAIL.n236 VTAIL.n218 104.615
R169 VTAIL.n229 VTAIL.n218 104.615
R170 VTAIL.n229 VTAIL.n228 104.615
R171 VTAIL.n228 VTAIL.n222 104.615
R172 VTAIL.n204 VTAIL.n203 104.615
R173 VTAIL.n203 VTAIL.n202 104.615
R174 VTAIL.n202 VTAIL.n171 104.615
R175 VTAIL.n195 VTAIL.n171 104.615
R176 VTAIL.n195 VTAIL.n194 104.615
R177 VTAIL.n194 VTAIL.n176 104.615
R178 VTAIL.n187 VTAIL.n176 104.615
R179 VTAIL.n187 VTAIL.n186 104.615
R180 VTAIL.n186 VTAIL.n180 104.615
R181 VTAIL.n162 VTAIL.n161 104.615
R182 VTAIL.n161 VTAIL.n160 104.615
R183 VTAIL.n160 VTAIL.n129 104.615
R184 VTAIL.n153 VTAIL.n129 104.615
R185 VTAIL.n153 VTAIL.n152 104.615
R186 VTAIL.n152 VTAIL.n134 104.615
R187 VTAIL.n145 VTAIL.n134 104.615
R188 VTAIL.n145 VTAIL.n144 104.615
R189 VTAIL.n144 VTAIL.n138 104.615
R190 VTAIL.t1 VTAIL.n305 52.3082
R191 VTAIL.t3 VTAIL.n11 52.3082
R192 VTAIL.t6 VTAIL.n53 52.3082
R193 VTAIL.t4 VTAIL.n95 52.3082
R194 VTAIL.t7 VTAIL.n264 52.3082
R195 VTAIL.t5 VTAIL.n222 52.3082
R196 VTAIL.t0 VTAIL.n180 52.3082
R197 VTAIL.t2 VTAIL.n138 52.3082
R198 VTAIL.n335 VTAIL.n334 32.9611
R199 VTAIL.n41 VTAIL.n40 32.9611
R200 VTAIL.n83 VTAIL.n82 32.9611
R201 VTAIL.n125 VTAIL.n124 32.9611
R202 VTAIL.n293 VTAIL.n292 32.9611
R203 VTAIL.n251 VTAIL.n250 32.9611
R204 VTAIL.n209 VTAIL.n208 32.9611
R205 VTAIL.n167 VTAIL.n166 32.9611
R206 VTAIL.n335 VTAIL.n293 20.6772
R207 VTAIL.n167 VTAIL.n125 20.6772
R208 VTAIL.n331 VTAIL.n296 13.1884
R209 VTAIL.n37 VTAIL.n2 13.1884
R210 VTAIL.n79 VTAIL.n44 13.1884
R211 VTAIL.n121 VTAIL.n86 13.1884
R212 VTAIL.n289 VTAIL.n254 13.1884
R213 VTAIL.n247 VTAIL.n212 13.1884
R214 VTAIL.n205 VTAIL.n170 13.1884
R215 VTAIL.n163 VTAIL.n128 13.1884
R216 VTAIL.n327 VTAIL.n326 12.8005
R217 VTAIL.n332 VTAIL.n294 12.8005
R218 VTAIL.n33 VTAIL.n32 12.8005
R219 VTAIL.n38 VTAIL.n0 12.8005
R220 VTAIL.n75 VTAIL.n74 12.8005
R221 VTAIL.n80 VTAIL.n42 12.8005
R222 VTAIL.n117 VTAIL.n116 12.8005
R223 VTAIL.n122 VTAIL.n84 12.8005
R224 VTAIL.n290 VTAIL.n252 12.8005
R225 VTAIL.n285 VTAIL.n256 12.8005
R226 VTAIL.n248 VTAIL.n210 12.8005
R227 VTAIL.n243 VTAIL.n214 12.8005
R228 VTAIL.n206 VTAIL.n168 12.8005
R229 VTAIL.n201 VTAIL.n172 12.8005
R230 VTAIL.n164 VTAIL.n126 12.8005
R231 VTAIL.n159 VTAIL.n130 12.8005
R232 VTAIL.n325 VTAIL.n298 12.0247
R233 VTAIL.n31 VTAIL.n4 12.0247
R234 VTAIL.n73 VTAIL.n46 12.0247
R235 VTAIL.n115 VTAIL.n88 12.0247
R236 VTAIL.n284 VTAIL.n257 12.0247
R237 VTAIL.n242 VTAIL.n215 12.0247
R238 VTAIL.n200 VTAIL.n173 12.0247
R239 VTAIL.n158 VTAIL.n131 12.0247
R240 VTAIL.n322 VTAIL.n321 11.249
R241 VTAIL.n28 VTAIL.n27 11.249
R242 VTAIL.n70 VTAIL.n69 11.249
R243 VTAIL.n112 VTAIL.n111 11.249
R244 VTAIL.n281 VTAIL.n280 11.249
R245 VTAIL.n239 VTAIL.n238 11.249
R246 VTAIL.n197 VTAIL.n196 11.249
R247 VTAIL.n155 VTAIL.n154 11.249
R248 VTAIL.n318 VTAIL.n300 10.4732
R249 VTAIL.n24 VTAIL.n6 10.4732
R250 VTAIL.n66 VTAIL.n48 10.4732
R251 VTAIL.n108 VTAIL.n90 10.4732
R252 VTAIL.n277 VTAIL.n259 10.4732
R253 VTAIL.n235 VTAIL.n217 10.4732
R254 VTAIL.n193 VTAIL.n175 10.4732
R255 VTAIL.n151 VTAIL.n133 10.4732
R256 VTAIL.n307 VTAIL.n306 10.2747
R257 VTAIL.n13 VTAIL.n12 10.2747
R258 VTAIL.n55 VTAIL.n54 10.2747
R259 VTAIL.n97 VTAIL.n96 10.2747
R260 VTAIL.n266 VTAIL.n265 10.2747
R261 VTAIL.n224 VTAIL.n223 10.2747
R262 VTAIL.n182 VTAIL.n181 10.2747
R263 VTAIL.n140 VTAIL.n139 10.2747
R264 VTAIL.n317 VTAIL.n302 9.69747
R265 VTAIL.n23 VTAIL.n8 9.69747
R266 VTAIL.n65 VTAIL.n50 9.69747
R267 VTAIL.n107 VTAIL.n92 9.69747
R268 VTAIL.n276 VTAIL.n261 9.69747
R269 VTAIL.n234 VTAIL.n219 9.69747
R270 VTAIL.n192 VTAIL.n177 9.69747
R271 VTAIL.n150 VTAIL.n135 9.69747
R272 VTAIL.n334 VTAIL.n333 9.45567
R273 VTAIL.n40 VTAIL.n39 9.45567
R274 VTAIL.n82 VTAIL.n81 9.45567
R275 VTAIL.n124 VTAIL.n123 9.45567
R276 VTAIL.n292 VTAIL.n291 9.45567
R277 VTAIL.n250 VTAIL.n249 9.45567
R278 VTAIL.n208 VTAIL.n207 9.45567
R279 VTAIL.n166 VTAIL.n165 9.45567
R280 VTAIL.n333 VTAIL.n332 9.3005
R281 VTAIL.n309 VTAIL.n308 9.3005
R282 VTAIL.n304 VTAIL.n303 9.3005
R283 VTAIL.n315 VTAIL.n314 9.3005
R284 VTAIL.n317 VTAIL.n316 9.3005
R285 VTAIL.n300 VTAIL.n299 9.3005
R286 VTAIL.n323 VTAIL.n322 9.3005
R287 VTAIL.n325 VTAIL.n324 9.3005
R288 VTAIL.n326 VTAIL.n295 9.3005
R289 VTAIL.n39 VTAIL.n38 9.3005
R290 VTAIL.n15 VTAIL.n14 9.3005
R291 VTAIL.n10 VTAIL.n9 9.3005
R292 VTAIL.n21 VTAIL.n20 9.3005
R293 VTAIL.n23 VTAIL.n22 9.3005
R294 VTAIL.n6 VTAIL.n5 9.3005
R295 VTAIL.n29 VTAIL.n28 9.3005
R296 VTAIL.n31 VTAIL.n30 9.3005
R297 VTAIL.n32 VTAIL.n1 9.3005
R298 VTAIL.n81 VTAIL.n80 9.3005
R299 VTAIL.n57 VTAIL.n56 9.3005
R300 VTAIL.n52 VTAIL.n51 9.3005
R301 VTAIL.n63 VTAIL.n62 9.3005
R302 VTAIL.n65 VTAIL.n64 9.3005
R303 VTAIL.n48 VTAIL.n47 9.3005
R304 VTAIL.n71 VTAIL.n70 9.3005
R305 VTAIL.n73 VTAIL.n72 9.3005
R306 VTAIL.n74 VTAIL.n43 9.3005
R307 VTAIL.n123 VTAIL.n122 9.3005
R308 VTAIL.n99 VTAIL.n98 9.3005
R309 VTAIL.n94 VTAIL.n93 9.3005
R310 VTAIL.n105 VTAIL.n104 9.3005
R311 VTAIL.n107 VTAIL.n106 9.3005
R312 VTAIL.n90 VTAIL.n89 9.3005
R313 VTAIL.n113 VTAIL.n112 9.3005
R314 VTAIL.n115 VTAIL.n114 9.3005
R315 VTAIL.n116 VTAIL.n85 9.3005
R316 VTAIL.n268 VTAIL.n267 9.3005
R317 VTAIL.n263 VTAIL.n262 9.3005
R318 VTAIL.n274 VTAIL.n273 9.3005
R319 VTAIL.n276 VTAIL.n275 9.3005
R320 VTAIL.n259 VTAIL.n258 9.3005
R321 VTAIL.n282 VTAIL.n281 9.3005
R322 VTAIL.n284 VTAIL.n283 9.3005
R323 VTAIL.n256 VTAIL.n253 9.3005
R324 VTAIL.n291 VTAIL.n290 9.3005
R325 VTAIL.n226 VTAIL.n225 9.3005
R326 VTAIL.n221 VTAIL.n220 9.3005
R327 VTAIL.n232 VTAIL.n231 9.3005
R328 VTAIL.n234 VTAIL.n233 9.3005
R329 VTAIL.n217 VTAIL.n216 9.3005
R330 VTAIL.n240 VTAIL.n239 9.3005
R331 VTAIL.n242 VTAIL.n241 9.3005
R332 VTAIL.n214 VTAIL.n211 9.3005
R333 VTAIL.n249 VTAIL.n248 9.3005
R334 VTAIL.n184 VTAIL.n183 9.3005
R335 VTAIL.n179 VTAIL.n178 9.3005
R336 VTAIL.n190 VTAIL.n189 9.3005
R337 VTAIL.n192 VTAIL.n191 9.3005
R338 VTAIL.n175 VTAIL.n174 9.3005
R339 VTAIL.n198 VTAIL.n197 9.3005
R340 VTAIL.n200 VTAIL.n199 9.3005
R341 VTAIL.n172 VTAIL.n169 9.3005
R342 VTAIL.n207 VTAIL.n206 9.3005
R343 VTAIL.n142 VTAIL.n141 9.3005
R344 VTAIL.n137 VTAIL.n136 9.3005
R345 VTAIL.n148 VTAIL.n147 9.3005
R346 VTAIL.n150 VTAIL.n149 9.3005
R347 VTAIL.n133 VTAIL.n132 9.3005
R348 VTAIL.n156 VTAIL.n155 9.3005
R349 VTAIL.n158 VTAIL.n157 9.3005
R350 VTAIL.n130 VTAIL.n127 9.3005
R351 VTAIL.n165 VTAIL.n164 9.3005
R352 VTAIL.n314 VTAIL.n313 8.92171
R353 VTAIL.n20 VTAIL.n19 8.92171
R354 VTAIL.n62 VTAIL.n61 8.92171
R355 VTAIL.n104 VTAIL.n103 8.92171
R356 VTAIL.n273 VTAIL.n272 8.92171
R357 VTAIL.n231 VTAIL.n230 8.92171
R358 VTAIL.n189 VTAIL.n188 8.92171
R359 VTAIL.n147 VTAIL.n146 8.92171
R360 VTAIL.n310 VTAIL.n304 8.14595
R361 VTAIL.n16 VTAIL.n10 8.14595
R362 VTAIL.n58 VTAIL.n52 8.14595
R363 VTAIL.n100 VTAIL.n94 8.14595
R364 VTAIL.n269 VTAIL.n263 8.14595
R365 VTAIL.n227 VTAIL.n221 8.14595
R366 VTAIL.n185 VTAIL.n179 8.14595
R367 VTAIL.n143 VTAIL.n137 8.14595
R368 VTAIL.n309 VTAIL.n306 7.3702
R369 VTAIL.n15 VTAIL.n12 7.3702
R370 VTAIL.n57 VTAIL.n54 7.3702
R371 VTAIL.n99 VTAIL.n96 7.3702
R372 VTAIL.n268 VTAIL.n265 7.3702
R373 VTAIL.n226 VTAIL.n223 7.3702
R374 VTAIL.n184 VTAIL.n181 7.3702
R375 VTAIL.n142 VTAIL.n139 7.3702
R376 VTAIL.n310 VTAIL.n309 5.81868
R377 VTAIL.n16 VTAIL.n15 5.81868
R378 VTAIL.n58 VTAIL.n57 5.81868
R379 VTAIL.n100 VTAIL.n99 5.81868
R380 VTAIL.n269 VTAIL.n268 5.81868
R381 VTAIL.n227 VTAIL.n226 5.81868
R382 VTAIL.n185 VTAIL.n184 5.81868
R383 VTAIL.n143 VTAIL.n142 5.81868
R384 VTAIL.n313 VTAIL.n304 5.04292
R385 VTAIL.n19 VTAIL.n10 5.04292
R386 VTAIL.n61 VTAIL.n52 5.04292
R387 VTAIL.n103 VTAIL.n94 5.04292
R388 VTAIL.n272 VTAIL.n263 5.04292
R389 VTAIL.n230 VTAIL.n221 5.04292
R390 VTAIL.n188 VTAIL.n179 5.04292
R391 VTAIL.n146 VTAIL.n137 5.04292
R392 VTAIL.n314 VTAIL.n302 4.26717
R393 VTAIL.n20 VTAIL.n8 4.26717
R394 VTAIL.n62 VTAIL.n50 4.26717
R395 VTAIL.n104 VTAIL.n92 4.26717
R396 VTAIL.n273 VTAIL.n261 4.26717
R397 VTAIL.n231 VTAIL.n219 4.26717
R398 VTAIL.n189 VTAIL.n177 4.26717
R399 VTAIL.n147 VTAIL.n135 4.26717
R400 VTAIL.n318 VTAIL.n317 3.49141
R401 VTAIL.n24 VTAIL.n23 3.49141
R402 VTAIL.n66 VTAIL.n65 3.49141
R403 VTAIL.n108 VTAIL.n107 3.49141
R404 VTAIL.n277 VTAIL.n276 3.49141
R405 VTAIL.n235 VTAIL.n234 3.49141
R406 VTAIL.n193 VTAIL.n192 3.49141
R407 VTAIL.n151 VTAIL.n150 3.49141
R408 VTAIL.n308 VTAIL.n307 2.84304
R409 VTAIL.n14 VTAIL.n13 2.84304
R410 VTAIL.n56 VTAIL.n55 2.84304
R411 VTAIL.n98 VTAIL.n97 2.84304
R412 VTAIL.n267 VTAIL.n266 2.84304
R413 VTAIL.n225 VTAIL.n224 2.84304
R414 VTAIL.n183 VTAIL.n182 2.84304
R415 VTAIL.n141 VTAIL.n140 2.84304
R416 VTAIL.n321 VTAIL.n300 2.71565
R417 VTAIL.n27 VTAIL.n6 2.71565
R418 VTAIL.n69 VTAIL.n48 2.71565
R419 VTAIL.n111 VTAIL.n90 2.71565
R420 VTAIL.n280 VTAIL.n259 2.71565
R421 VTAIL.n238 VTAIL.n217 2.71565
R422 VTAIL.n196 VTAIL.n175 2.71565
R423 VTAIL.n154 VTAIL.n133 2.71565
R424 VTAIL.n322 VTAIL.n298 1.93989
R425 VTAIL.n28 VTAIL.n4 1.93989
R426 VTAIL.n70 VTAIL.n46 1.93989
R427 VTAIL.n112 VTAIL.n88 1.93989
R428 VTAIL.n281 VTAIL.n257 1.93989
R429 VTAIL.n239 VTAIL.n215 1.93989
R430 VTAIL.n197 VTAIL.n173 1.93989
R431 VTAIL.n155 VTAIL.n131 1.93989
R432 VTAIL.n209 VTAIL.n167 1.55222
R433 VTAIL.n293 VTAIL.n251 1.55222
R434 VTAIL.n125 VTAIL.n83 1.55222
R435 VTAIL.n327 VTAIL.n325 1.16414
R436 VTAIL.n334 VTAIL.n294 1.16414
R437 VTAIL.n33 VTAIL.n31 1.16414
R438 VTAIL.n40 VTAIL.n0 1.16414
R439 VTAIL.n75 VTAIL.n73 1.16414
R440 VTAIL.n82 VTAIL.n42 1.16414
R441 VTAIL.n117 VTAIL.n115 1.16414
R442 VTAIL.n124 VTAIL.n84 1.16414
R443 VTAIL.n292 VTAIL.n252 1.16414
R444 VTAIL.n285 VTAIL.n284 1.16414
R445 VTAIL.n250 VTAIL.n210 1.16414
R446 VTAIL.n243 VTAIL.n242 1.16414
R447 VTAIL.n208 VTAIL.n168 1.16414
R448 VTAIL.n201 VTAIL.n200 1.16414
R449 VTAIL.n166 VTAIL.n126 1.16414
R450 VTAIL.n159 VTAIL.n158 1.16414
R451 VTAIL VTAIL.n41 0.834552
R452 VTAIL VTAIL.n335 0.718172
R453 VTAIL.n251 VTAIL.n209 0.470328
R454 VTAIL.n83 VTAIL.n41 0.470328
R455 VTAIL.n326 VTAIL.n296 0.388379
R456 VTAIL.n332 VTAIL.n331 0.388379
R457 VTAIL.n32 VTAIL.n2 0.388379
R458 VTAIL.n38 VTAIL.n37 0.388379
R459 VTAIL.n74 VTAIL.n44 0.388379
R460 VTAIL.n80 VTAIL.n79 0.388379
R461 VTAIL.n116 VTAIL.n86 0.388379
R462 VTAIL.n122 VTAIL.n121 0.388379
R463 VTAIL.n290 VTAIL.n289 0.388379
R464 VTAIL.n256 VTAIL.n254 0.388379
R465 VTAIL.n248 VTAIL.n247 0.388379
R466 VTAIL.n214 VTAIL.n212 0.388379
R467 VTAIL.n206 VTAIL.n205 0.388379
R468 VTAIL.n172 VTAIL.n170 0.388379
R469 VTAIL.n164 VTAIL.n163 0.388379
R470 VTAIL.n130 VTAIL.n128 0.388379
R471 VTAIL.n308 VTAIL.n303 0.155672
R472 VTAIL.n315 VTAIL.n303 0.155672
R473 VTAIL.n316 VTAIL.n315 0.155672
R474 VTAIL.n316 VTAIL.n299 0.155672
R475 VTAIL.n323 VTAIL.n299 0.155672
R476 VTAIL.n324 VTAIL.n323 0.155672
R477 VTAIL.n324 VTAIL.n295 0.155672
R478 VTAIL.n333 VTAIL.n295 0.155672
R479 VTAIL.n14 VTAIL.n9 0.155672
R480 VTAIL.n21 VTAIL.n9 0.155672
R481 VTAIL.n22 VTAIL.n21 0.155672
R482 VTAIL.n22 VTAIL.n5 0.155672
R483 VTAIL.n29 VTAIL.n5 0.155672
R484 VTAIL.n30 VTAIL.n29 0.155672
R485 VTAIL.n30 VTAIL.n1 0.155672
R486 VTAIL.n39 VTAIL.n1 0.155672
R487 VTAIL.n56 VTAIL.n51 0.155672
R488 VTAIL.n63 VTAIL.n51 0.155672
R489 VTAIL.n64 VTAIL.n63 0.155672
R490 VTAIL.n64 VTAIL.n47 0.155672
R491 VTAIL.n71 VTAIL.n47 0.155672
R492 VTAIL.n72 VTAIL.n71 0.155672
R493 VTAIL.n72 VTAIL.n43 0.155672
R494 VTAIL.n81 VTAIL.n43 0.155672
R495 VTAIL.n98 VTAIL.n93 0.155672
R496 VTAIL.n105 VTAIL.n93 0.155672
R497 VTAIL.n106 VTAIL.n105 0.155672
R498 VTAIL.n106 VTAIL.n89 0.155672
R499 VTAIL.n113 VTAIL.n89 0.155672
R500 VTAIL.n114 VTAIL.n113 0.155672
R501 VTAIL.n114 VTAIL.n85 0.155672
R502 VTAIL.n123 VTAIL.n85 0.155672
R503 VTAIL.n291 VTAIL.n253 0.155672
R504 VTAIL.n283 VTAIL.n253 0.155672
R505 VTAIL.n283 VTAIL.n282 0.155672
R506 VTAIL.n282 VTAIL.n258 0.155672
R507 VTAIL.n275 VTAIL.n258 0.155672
R508 VTAIL.n275 VTAIL.n274 0.155672
R509 VTAIL.n274 VTAIL.n262 0.155672
R510 VTAIL.n267 VTAIL.n262 0.155672
R511 VTAIL.n249 VTAIL.n211 0.155672
R512 VTAIL.n241 VTAIL.n211 0.155672
R513 VTAIL.n241 VTAIL.n240 0.155672
R514 VTAIL.n240 VTAIL.n216 0.155672
R515 VTAIL.n233 VTAIL.n216 0.155672
R516 VTAIL.n233 VTAIL.n232 0.155672
R517 VTAIL.n232 VTAIL.n220 0.155672
R518 VTAIL.n225 VTAIL.n220 0.155672
R519 VTAIL.n207 VTAIL.n169 0.155672
R520 VTAIL.n199 VTAIL.n169 0.155672
R521 VTAIL.n199 VTAIL.n198 0.155672
R522 VTAIL.n198 VTAIL.n174 0.155672
R523 VTAIL.n191 VTAIL.n174 0.155672
R524 VTAIL.n191 VTAIL.n190 0.155672
R525 VTAIL.n190 VTAIL.n178 0.155672
R526 VTAIL.n183 VTAIL.n178 0.155672
R527 VTAIL.n165 VTAIL.n127 0.155672
R528 VTAIL.n157 VTAIL.n127 0.155672
R529 VTAIL.n157 VTAIL.n156 0.155672
R530 VTAIL.n156 VTAIL.n132 0.155672
R531 VTAIL.n149 VTAIL.n132 0.155672
R532 VTAIL.n149 VTAIL.n148 0.155672
R533 VTAIL.n148 VTAIL.n136 0.155672
R534 VTAIL.n141 VTAIL.n136 0.155672
R535 VDD1 VDD1.n1 100.406
R536 VDD1 VDD1.n0 64.8117
R537 VDD1.n0 VDD1.t0 2.52601
R538 VDD1.n0 VDD1.t3 2.52601
R539 VDD1.n1 VDD1.t2 2.52601
R540 VDD1.n1 VDD1.t1 2.52601
R541 B.n544 B.n543 585
R542 B.n218 B.n81 585
R543 B.n217 B.n216 585
R544 B.n215 B.n214 585
R545 B.n213 B.n212 585
R546 B.n211 B.n210 585
R547 B.n209 B.n208 585
R548 B.n207 B.n206 585
R549 B.n205 B.n204 585
R550 B.n203 B.n202 585
R551 B.n201 B.n200 585
R552 B.n199 B.n198 585
R553 B.n197 B.n196 585
R554 B.n195 B.n194 585
R555 B.n193 B.n192 585
R556 B.n191 B.n190 585
R557 B.n189 B.n188 585
R558 B.n187 B.n186 585
R559 B.n185 B.n184 585
R560 B.n183 B.n182 585
R561 B.n181 B.n180 585
R562 B.n179 B.n178 585
R563 B.n177 B.n176 585
R564 B.n175 B.n174 585
R565 B.n173 B.n172 585
R566 B.n171 B.n170 585
R567 B.n169 B.n168 585
R568 B.n167 B.n166 585
R569 B.n165 B.n164 585
R570 B.n162 B.n161 585
R571 B.n160 B.n159 585
R572 B.n158 B.n157 585
R573 B.n156 B.n155 585
R574 B.n154 B.n153 585
R575 B.n152 B.n151 585
R576 B.n150 B.n149 585
R577 B.n148 B.n147 585
R578 B.n146 B.n145 585
R579 B.n144 B.n143 585
R580 B.n141 B.n140 585
R581 B.n139 B.n138 585
R582 B.n137 B.n136 585
R583 B.n135 B.n134 585
R584 B.n133 B.n132 585
R585 B.n131 B.n130 585
R586 B.n129 B.n128 585
R587 B.n127 B.n126 585
R588 B.n125 B.n124 585
R589 B.n123 B.n122 585
R590 B.n121 B.n120 585
R591 B.n119 B.n118 585
R592 B.n117 B.n116 585
R593 B.n115 B.n114 585
R594 B.n113 B.n112 585
R595 B.n111 B.n110 585
R596 B.n109 B.n108 585
R597 B.n107 B.n106 585
R598 B.n105 B.n104 585
R599 B.n103 B.n102 585
R600 B.n101 B.n100 585
R601 B.n99 B.n98 585
R602 B.n97 B.n96 585
R603 B.n95 B.n94 585
R604 B.n93 B.n92 585
R605 B.n91 B.n90 585
R606 B.n89 B.n88 585
R607 B.n87 B.n86 585
R608 B.n46 B.n45 585
R609 B.n542 B.n47 585
R610 B.n547 B.n47 585
R611 B.n541 B.n540 585
R612 B.n540 B.n43 585
R613 B.n539 B.n42 585
R614 B.n553 B.n42 585
R615 B.n538 B.n41 585
R616 B.n554 B.n41 585
R617 B.n537 B.n40 585
R618 B.n555 B.n40 585
R619 B.n536 B.n535 585
R620 B.n535 B.n39 585
R621 B.n534 B.n35 585
R622 B.n561 B.n35 585
R623 B.n533 B.n34 585
R624 B.n562 B.n34 585
R625 B.n532 B.n33 585
R626 B.n563 B.n33 585
R627 B.n531 B.n530 585
R628 B.n530 B.n29 585
R629 B.n529 B.n28 585
R630 B.n569 B.n28 585
R631 B.n528 B.n27 585
R632 B.n570 B.n27 585
R633 B.n527 B.n26 585
R634 B.n571 B.n26 585
R635 B.n526 B.n525 585
R636 B.n525 B.n22 585
R637 B.n524 B.n21 585
R638 B.n577 B.n21 585
R639 B.n523 B.n20 585
R640 B.n578 B.n20 585
R641 B.n522 B.n19 585
R642 B.n579 B.n19 585
R643 B.n521 B.n520 585
R644 B.n520 B.n15 585
R645 B.n519 B.n14 585
R646 B.n585 B.n14 585
R647 B.n518 B.n13 585
R648 B.n586 B.n13 585
R649 B.n517 B.n12 585
R650 B.n587 B.n12 585
R651 B.n516 B.n515 585
R652 B.n515 B.n8 585
R653 B.n514 B.n7 585
R654 B.n593 B.n7 585
R655 B.n513 B.n6 585
R656 B.n594 B.n6 585
R657 B.n512 B.n5 585
R658 B.n595 B.n5 585
R659 B.n511 B.n510 585
R660 B.n510 B.n4 585
R661 B.n509 B.n219 585
R662 B.n509 B.n508 585
R663 B.n499 B.n220 585
R664 B.n221 B.n220 585
R665 B.n501 B.n500 585
R666 B.n502 B.n501 585
R667 B.n498 B.n225 585
R668 B.n229 B.n225 585
R669 B.n497 B.n496 585
R670 B.n496 B.n495 585
R671 B.n227 B.n226 585
R672 B.n228 B.n227 585
R673 B.n488 B.n487 585
R674 B.n489 B.n488 585
R675 B.n486 B.n234 585
R676 B.n234 B.n233 585
R677 B.n485 B.n484 585
R678 B.n484 B.n483 585
R679 B.n236 B.n235 585
R680 B.n237 B.n236 585
R681 B.n476 B.n475 585
R682 B.n477 B.n476 585
R683 B.n474 B.n242 585
R684 B.n242 B.n241 585
R685 B.n473 B.n472 585
R686 B.n472 B.n471 585
R687 B.n244 B.n243 585
R688 B.n245 B.n244 585
R689 B.n464 B.n463 585
R690 B.n465 B.n464 585
R691 B.n462 B.n250 585
R692 B.n250 B.n249 585
R693 B.n461 B.n460 585
R694 B.n460 B.n459 585
R695 B.n252 B.n251 585
R696 B.n452 B.n252 585
R697 B.n451 B.n450 585
R698 B.n453 B.n451 585
R699 B.n449 B.n257 585
R700 B.n257 B.n256 585
R701 B.n448 B.n447 585
R702 B.n447 B.n446 585
R703 B.n259 B.n258 585
R704 B.n260 B.n259 585
R705 B.n439 B.n438 585
R706 B.n440 B.n439 585
R707 B.n263 B.n262 585
R708 B.n306 B.n305 585
R709 B.n307 B.n303 585
R710 B.n303 B.n264 585
R711 B.n309 B.n308 585
R712 B.n311 B.n302 585
R713 B.n314 B.n313 585
R714 B.n315 B.n301 585
R715 B.n317 B.n316 585
R716 B.n319 B.n300 585
R717 B.n322 B.n321 585
R718 B.n323 B.n299 585
R719 B.n325 B.n324 585
R720 B.n327 B.n298 585
R721 B.n330 B.n329 585
R722 B.n331 B.n297 585
R723 B.n333 B.n332 585
R724 B.n335 B.n296 585
R725 B.n338 B.n337 585
R726 B.n339 B.n295 585
R727 B.n341 B.n340 585
R728 B.n343 B.n294 585
R729 B.n346 B.n345 585
R730 B.n347 B.n293 585
R731 B.n349 B.n348 585
R732 B.n351 B.n292 585
R733 B.n354 B.n353 585
R734 B.n355 B.n291 585
R735 B.n357 B.n356 585
R736 B.n359 B.n290 585
R737 B.n362 B.n361 585
R738 B.n363 B.n286 585
R739 B.n365 B.n364 585
R740 B.n367 B.n285 585
R741 B.n370 B.n369 585
R742 B.n371 B.n284 585
R743 B.n373 B.n372 585
R744 B.n375 B.n283 585
R745 B.n378 B.n377 585
R746 B.n379 B.n280 585
R747 B.n382 B.n381 585
R748 B.n384 B.n279 585
R749 B.n387 B.n386 585
R750 B.n388 B.n278 585
R751 B.n390 B.n389 585
R752 B.n392 B.n277 585
R753 B.n395 B.n394 585
R754 B.n396 B.n276 585
R755 B.n398 B.n397 585
R756 B.n400 B.n275 585
R757 B.n403 B.n402 585
R758 B.n404 B.n274 585
R759 B.n406 B.n405 585
R760 B.n408 B.n273 585
R761 B.n411 B.n410 585
R762 B.n412 B.n272 585
R763 B.n414 B.n413 585
R764 B.n416 B.n271 585
R765 B.n419 B.n418 585
R766 B.n420 B.n270 585
R767 B.n422 B.n421 585
R768 B.n424 B.n269 585
R769 B.n427 B.n426 585
R770 B.n428 B.n268 585
R771 B.n430 B.n429 585
R772 B.n432 B.n267 585
R773 B.n433 B.n266 585
R774 B.n436 B.n435 585
R775 B.n437 B.n265 585
R776 B.n265 B.n264 585
R777 B.n442 B.n441 585
R778 B.n441 B.n440 585
R779 B.n443 B.n261 585
R780 B.n261 B.n260 585
R781 B.n445 B.n444 585
R782 B.n446 B.n445 585
R783 B.n255 B.n254 585
R784 B.n256 B.n255 585
R785 B.n455 B.n454 585
R786 B.n454 B.n453 585
R787 B.n456 B.n253 585
R788 B.n452 B.n253 585
R789 B.n458 B.n457 585
R790 B.n459 B.n458 585
R791 B.n248 B.n247 585
R792 B.n249 B.n248 585
R793 B.n467 B.n466 585
R794 B.n466 B.n465 585
R795 B.n468 B.n246 585
R796 B.n246 B.n245 585
R797 B.n470 B.n469 585
R798 B.n471 B.n470 585
R799 B.n240 B.n239 585
R800 B.n241 B.n240 585
R801 B.n479 B.n478 585
R802 B.n478 B.n477 585
R803 B.n480 B.n238 585
R804 B.n238 B.n237 585
R805 B.n482 B.n481 585
R806 B.n483 B.n482 585
R807 B.n232 B.n231 585
R808 B.n233 B.n232 585
R809 B.n491 B.n490 585
R810 B.n490 B.n489 585
R811 B.n492 B.n230 585
R812 B.n230 B.n228 585
R813 B.n494 B.n493 585
R814 B.n495 B.n494 585
R815 B.n224 B.n223 585
R816 B.n229 B.n224 585
R817 B.n504 B.n503 585
R818 B.n503 B.n502 585
R819 B.n505 B.n222 585
R820 B.n222 B.n221 585
R821 B.n507 B.n506 585
R822 B.n508 B.n507 585
R823 B.n2 B.n0 585
R824 B.n4 B.n2 585
R825 B.n3 B.n1 585
R826 B.n594 B.n3 585
R827 B.n592 B.n591 585
R828 B.n593 B.n592 585
R829 B.n590 B.n9 585
R830 B.n9 B.n8 585
R831 B.n589 B.n588 585
R832 B.n588 B.n587 585
R833 B.n11 B.n10 585
R834 B.n586 B.n11 585
R835 B.n584 B.n583 585
R836 B.n585 B.n584 585
R837 B.n582 B.n16 585
R838 B.n16 B.n15 585
R839 B.n581 B.n580 585
R840 B.n580 B.n579 585
R841 B.n18 B.n17 585
R842 B.n578 B.n18 585
R843 B.n576 B.n575 585
R844 B.n577 B.n576 585
R845 B.n574 B.n23 585
R846 B.n23 B.n22 585
R847 B.n573 B.n572 585
R848 B.n572 B.n571 585
R849 B.n25 B.n24 585
R850 B.n570 B.n25 585
R851 B.n568 B.n567 585
R852 B.n569 B.n568 585
R853 B.n566 B.n30 585
R854 B.n30 B.n29 585
R855 B.n565 B.n564 585
R856 B.n564 B.n563 585
R857 B.n32 B.n31 585
R858 B.n562 B.n32 585
R859 B.n560 B.n559 585
R860 B.n561 B.n560 585
R861 B.n558 B.n36 585
R862 B.n39 B.n36 585
R863 B.n557 B.n556 585
R864 B.n556 B.n555 585
R865 B.n38 B.n37 585
R866 B.n554 B.n38 585
R867 B.n552 B.n551 585
R868 B.n553 B.n552 585
R869 B.n550 B.n44 585
R870 B.n44 B.n43 585
R871 B.n549 B.n548 585
R872 B.n548 B.n547 585
R873 B.n597 B.n596 585
R874 B.n596 B.n595 585
R875 B.n441 B.n263 526.135
R876 B.n548 B.n46 526.135
R877 B.n439 B.n265 526.135
R878 B.n544 B.n47 526.135
R879 B.n281 B.t15 333.86
R880 B.n287 B.t4 333.86
R881 B.n84 B.t8 333.86
R882 B.n82 B.t12 333.86
R883 B.n546 B.n545 256.663
R884 B.n546 B.n80 256.663
R885 B.n546 B.n79 256.663
R886 B.n546 B.n78 256.663
R887 B.n546 B.n77 256.663
R888 B.n546 B.n76 256.663
R889 B.n546 B.n75 256.663
R890 B.n546 B.n74 256.663
R891 B.n546 B.n73 256.663
R892 B.n546 B.n72 256.663
R893 B.n546 B.n71 256.663
R894 B.n546 B.n70 256.663
R895 B.n546 B.n69 256.663
R896 B.n546 B.n68 256.663
R897 B.n546 B.n67 256.663
R898 B.n546 B.n66 256.663
R899 B.n546 B.n65 256.663
R900 B.n546 B.n64 256.663
R901 B.n546 B.n63 256.663
R902 B.n546 B.n62 256.663
R903 B.n546 B.n61 256.663
R904 B.n546 B.n60 256.663
R905 B.n546 B.n59 256.663
R906 B.n546 B.n58 256.663
R907 B.n546 B.n57 256.663
R908 B.n546 B.n56 256.663
R909 B.n546 B.n55 256.663
R910 B.n546 B.n54 256.663
R911 B.n546 B.n53 256.663
R912 B.n546 B.n52 256.663
R913 B.n546 B.n51 256.663
R914 B.n546 B.n50 256.663
R915 B.n546 B.n49 256.663
R916 B.n546 B.n48 256.663
R917 B.n304 B.n264 256.663
R918 B.n310 B.n264 256.663
R919 B.n312 B.n264 256.663
R920 B.n318 B.n264 256.663
R921 B.n320 B.n264 256.663
R922 B.n326 B.n264 256.663
R923 B.n328 B.n264 256.663
R924 B.n334 B.n264 256.663
R925 B.n336 B.n264 256.663
R926 B.n342 B.n264 256.663
R927 B.n344 B.n264 256.663
R928 B.n350 B.n264 256.663
R929 B.n352 B.n264 256.663
R930 B.n358 B.n264 256.663
R931 B.n360 B.n264 256.663
R932 B.n366 B.n264 256.663
R933 B.n368 B.n264 256.663
R934 B.n374 B.n264 256.663
R935 B.n376 B.n264 256.663
R936 B.n383 B.n264 256.663
R937 B.n385 B.n264 256.663
R938 B.n391 B.n264 256.663
R939 B.n393 B.n264 256.663
R940 B.n399 B.n264 256.663
R941 B.n401 B.n264 256.663
R942 B.n407 B.n264 256.663
R943 B.n409 B.n264 256.663
R944 B.n415 B.n264 256.663
R945 B.n417 B.n264 256.663
R946 B.n423 B.n264 256.663
R947 B.n425 B.n264 256.663
R948 B.n431 B.n264 256.663
R949 B.n434 B.n264 256.663
R950 B.n281 B.t17 245.097
R951 B.n82 B.t13 245.097
R952 B.n287 B.t7 245.097
R953 B.n84 B.t10 245.097
R954 B.n282 B.t16 210.189
R955 B.n83 B.t14 210.189
R956 B.n288 B.t6 210.189
R957 B.n85 B.t11 210.189
R958 B.n441 B.n261 163.367
R959 B.n445 B.n261 163.367
R960 B.n445 B.n255 163.367
R961 B.n454 B.n255 163.367
R962 B.n454 B.n253 163.367
R963 B.n458 B.n253 163.367
R964 B.n458 B.n248 163.367
R965 B.n466 B.n248 163.367
R966 B.n466 B.n246 163.367
R967 B.n470 B.n246 163.367
R968 B.n470 B.n240 163.367
R969 B.n478 B.n240 163.367
R970 B.n478 B.n238 163.367
R971 B.n482 B.n238 163.367
R972 B.n482 B.n232 163.367
R973 B.n490 B.n232 163.367
R974 B.n490 B.n230 163.367
R975 B.n494 B.n230 163.367
R976 B.n494 B.n224 163.367
R977 B.n503 B.n224 163.367
R978 B.n503 B.n222 163.367
R979 B.n507 B.n222 163.367
R980 B.n507 B.n2 163.367
R981 B.n596 B.n2 163.367
R982 B.n596 B.n3 163.367
R983 B.n592 B.n3 163.367
R984 B.n592 B.n9 163.367
R985 B.n588 B.n9 163.367
R986 B.n588 B.n11 163.367
R987 B.n584 B.n11 163.367
R988 B.n584 B.n16 163.367
R989 B.n580 B.n16 163.367
R990 B.n580 B.n18 163.367
R991 B.n576 B.n18 163.367
R992 B.n576 B.n23 163.367
R993 B.n572 B.n23 163.367
R994 B.n572 B.n25 163.367
R995 B.n568 B.n25 163.367
R996 B.n568 B.n30 163.367
R997 B.n564 B.n30 163.367
R998 B.n564 B.n32 163.367
R999 B.n560 B.n32 163.367
R1000 B.n560 B.n36 163.367
R1001 B.n556 B.n36 163.367
R1002 B.n556 B.n38 163.367
R1003 B.n552 B.n38 163.367
R1004 B.n552 B.n44 163.367
R1005 B.n548 B.n44 163.367
R1006 B.n305 B.n303 163.367
R1007 B.n309 B.n303 163.367
R1008 B.n313 B.n311 163.367
R1009 B.n317 B.n301 163.367
R1010 B.n321 B.n319 163.367
R1011 B.n325 B.n299 163.367
R1012 B.n329 B.n327 163.367
R1013 B.n333 B.n297 163.367
R1014 B.n337 B.n335 163.367
R1015 B.n341 B.n295 163.367
R1016 B.n345 B.n343 163.367
R1017 B.n349 B.n293 163.367
R1018 B.n353 B.n351 163.367
R1019 B.n357 B.n291 163.367
R1020 B.n361 B.n359 163.367
R1021 B.n365 B.n286 163.367
R1022 B.n369 B.n367 163.367
R1023 B.n373 B.n284 163.367
R1024 B.n377 B.n375 163.367
R1025 B.n382 B.n280 163.367
R1026 B.n386 B.n384 163.367
R1027 B.n390 B.n278 163.367
R1028 B.n394 B.n392 163.367
R1029 B.n398 B.n276 163.367
R1030 B.n402 B.n400 163.367
R1031 B.n406 B.n274 163.367
R1032 B.n410 B.n408 163.367
R1033 B.n414 B.n272 163.367
R1034 B.n418 B.n416 163.367
R1035 B.n422 B.n270 163.367
R1036 B.n426 B.n424 163.367
R1037 B.n430 B.n268 163.367
R1038 B.n433 B.n432 163.367
R1039 B.n435 B.n265 163.367
R1040 B.n439 B.n259 163.367
R1041 B.n447 B.n259 163.367
R1042 B.n447 B.n257 163.367
R1043 B.n451 B.n257 163.367
R1044 B.n451 B.n252 163.367
R1045 B.n460 B.n252 163.367
R1046 B.n460 B.n250 163.367
R1047 B.n464 B.n250 163.367
R1048 B.n464 B.n244 163.367
R1049 B.n472 B.n244 163.367
R1050 B.n472 B.n242 163.367
R1051 B.n476 B.n242 163.367
R1052 B.n476 B.n236 163.367
R1053 B.n484 B.n236 163.367
R1054 B.n484 B.n234 163.367
R1055 B.n488 B.n234 163.367
R1056 B.n488 B.n227 163.367
R1057 B.n496 B.n227 163.367
R1058 B.n496 B.n225 163.367
R1059 B.n501 B.n225 163.367
R1060 B.n501 B.n220 163.367
R1061 B.n509 B.n220 163.367
R1062 B.n510 B.n509 163.367
R1063 B.n510 B.n5 163.367
R1064 B.n6 B.n5 163.367
R1065 B.n7 B.n6 163.367
R1066 B.n515 B.n7 163.367
R1067 B.n515 B.n12 163.367
R1068 B.n13 B.n12 163.367
R1069 B.n14 B.n13 163.367
R1070 B.n520 B.n14 163.367
R1071 B.n520 B.n19 163.367
R1072 B.n20 B.n19 163.367
R1073 B.n21 B.n20 163.367
R1074 B.n525 B.n21 163.367
R1075 B.n525 B.n26 163.367
R1076 B.n27 B.n26 163.367
R1077 B.n28 B.n27 163.367
R1078 B.n530 B.n28 163.367
R1079 B.n530 B.n33 163.367
R1080 B.n34 B.n33 163.367
R1081 B.n35 B.n34 163.367
R1082 B.n535 B.n35 163.367
R1083 B.n535 B.n40 163.367
R1084 B.n41 B.n40 163.367
R1085 B.n42 B.n41 163.367
R1086 B.n540 B.n42 163.367
R1087 B.n540 B.n47 163.367
R1088 B.n88 B.n87 163.367
R1089 B.n92 B.n91 163.367
R1090 B.n96 B.n95 163.367
R1091 B.n100 B.n99 163.367
R1092 B.n104 B.n103 163.367
R1093 B.n108 B.n107 163.367
R1094 B.n112 B.n111 163.367
R1095 B.n116 B.n115 163.367
R1096 B.n120 B.n119 163.367
R1097 B.n124 B.n123 163.367
R1098 B.n128 B.n127 163.367
R1099 B.n132 B.n131 163.367
R1100 B.n136 B.n135 163.367
R1101 B.n140 B.n139 163.367
R1102 B.n145 B.n144 163.367
R1103 B.n149 B.n148 163.367
R1104 B.n153 B.n152 163.367
R1105 B.n157 B.n156 163.367
R1106 B.n161 B.n160 163.367
R1107 B.n166 B.n165 163.367
R1108 B.n170 B.n169 163.367
R1109 B.n174 B.n173 163.367
R1110 B.n178 B.n177 163.367
R1111 B.n182 B.n181 163.367
R1112 B.n186 B.n185 163.367
R1113 B.n190 B.n189 163.367
R1114 B.n194 B.n193 163.367
R1115 B.n198 B.n197 163.367
R1116 B.n202 B.n201 163.367
R1117 B.n206 B.n205 163.367
R1118 B.n210 B.n209 163.367
R1119 B.n214 B.n213 163.367
R1120 B.n216 B.n81 163.367
R1121 B.n440 B.n264 103.165
R1122 B.n547 B.n546 103.165
R1123 B.n304 B.n263 71.676
R1124 B.n310 B.n309 71.676
R1125 B.n313 B.n312 71.676
R1126 B.n318 B.n317 71.676
R1127 B.n321 B.n320 71.676
R1128 B.n326 B.n325 71.676
R1129 B.n329 B.n328 71.676
R1130 B.n334 B.n333 71.676
R1131 B.n337 B.n336 71.676
R1132 B.n342 B.n341 71.676
R1133 B.n345 B.n344 71.676
R1134 B.n350 B.n349 71.676
R1135 B.n353 B.n352 71.676
R1136 B.n358 B.n357 71.676
R1137 B.n361 B.n360 71.676
R1138 B.n366 B.n365 71.676
R1139 B.n369 B.n368 71.676
R1140 B.n374 B.n373 71.676
R1141 B.n377 B.n376 71.676
R1142 B.n383 B.n382 71.676
R1143 B.n386 B.n385 71.676
R1144 B.n391 B.n390 71.676
R1145 B.n394 B.n393 71.676
R1146 B.n399 B.n398 71.676
R1147 B.n402 B.n401 71.676
R1148 B.n407 B.n406 71.676
R1149 B.n410 B.n409 71.676
R1150 B.n415 B.n414 71.676
R1151 B.n418 B.n417 71.676
R1152 B.n423 B.n422 71.676
R1153 B.n426 B.n425 71.676
R1154 B.n431 B.n430 71.676
R1155 B.n434 B.n433 71.676
R1156 B.n48 B.n46 71.676
R1157 B.n88 B.n49 71.676
R1158 B.n92 B.n50 71.676
R1159 B.n96 B.n51 71.676
R1160 B.n100 B.n52 71.676
R1161 B.n104 B.n53 71.676
R1162 B.n108 B.n54 71.676
R1163 B.n112 B.n55 71.676
R1164 B.n116 B.n56 71.676
R1165 B.n120 B.n57 71.676
R1166 B.n124 B.n58 71.676
R1167 B.n128 B.n59 71.676
R1168 B.n132 B.n60 71.676
R1169 B.n136 B.n61 71.676
R1170 B.n140 B.n62 71.676
R1171 B.n145 B.n63 71.676
R1172 B.n149 B.n64 71.676
R1173 B.n153 B.n65 71.676
R1174 B.n157 B.n66 71.676
R1175 B.n161 B.n67 71.676
R1176 B.n166 B.n68 71.676
R1177 B.n170 B.n69 71.676
R1178 B.n174 B.n70 71.676
R1179 B.n178 B.n71 71.676
R1180 B.n182 B.n72 71.676
R1181 B.n186 B.n73 71.676
R1182 B.n190 B.n74 71.676
R1183 B.n194 B.n75 71.676
R1184 B.n198 B.n76 71.676
R1185 B.n202 B.n77 71.676
R1186 B.n206 B.n78 71.676
R1187 B.n210 B.n79 71.676
R1188 B.n214 B.n80 71.676
R1189 B.n545 B.n81 71.676
R1190 B.n545 B.n544 71.676
R1191 B.n216 B.n80 71.676
R1192 B.n213 B.n79 71.676
R1193 B.n209 B.n78 71.676
R1194 B.n205 B.n77 71.676
R1195 B.n201 B.n76 71.676
R1196 B.n197 B.n75 71.676
R1197 B.n193 B.n74 71.676
R1198 B.n189 B.n73 71.676
R1199 B.n185 B.n72 71.676
R1200 B.n181 B.n71 71.676
R1201 B.n177 B.n70 71.676
R1202 B.n173 B.n69 71.676
R1203 B.n169 B.n68 71.676
R1204 B.n165 B.n67 71.676
R1205 B.n160 B.n66 71.676
R1206 B.n156 B.n65 71.676
R1207 B.n152 B.n64 71.676
R1208 B.n148 B.n63 71.676
R1209 B.n144 B.n62 71.676
R1210 B.n139 B.n61 71.676
R1211 B.n135 B.n60 71.676
R1212 B.n131 B.n59 71.676
R1213 B.n127 B.n58 71.676
R1214 B.n123 B.n57 71.676
R1215 B.n119 B.n56 71.676
R1216 B.n115 B.n55 71.676
R1217 B.n111 B.n54 71.676
R1218 B.n107 B.n53 71.676
R1219 B.n103 B.n52 71.676
R1220 B.n99 B.n51 71.676
R1221 B.n95 B.n50 71.676
R1222 B.n91 B.n49 71.676
R1223 B.n87 B.n48 71.676
R1224 B.n305 B.n304 71.676
R1225 B.n311 B.n310 71.676
R1226 B.n312 B.n301 71.676
R1227 B.n319 B.n318 71.676
R1228 B.n320 B.n299 71.676
R1229 B.n327 B.n326 71.676
R1230 B.n328 B.n297 71.676
R1231 B.n335 B.n334 71.676
R1232 B.n336 B.n295 71.676
R1233 B.n343 B.n342 71.676
R1234 B.n344 B.n293 71.676
R1235 B.n351 B.n350 71.676
R1236 B.n352 B.n291 71.676
R1237 B.n359 B.n358 71.676
R1238 B.n360 B.n286 71.676
R1239 B.n367 B.n366 71.676
R1240 B.n368 B.n284 71.676
R1241 B.n375 B.n374 71.676
R1242 B.n376 B.n280 71.676
R1243 B.n384 B.n383 71.676
R1244 B.n385 B.n278 71.676
R1245 B.n392 B.n391 71.676
R1246 B.n393 B.n276 71.676
R1247 B.n400 B.n399 71.676
R1248 B.n401 B.n274 71.676
R1249 B.n408 B.n407 71.676
R1250 B.n409 B.n272 71.676
R1251 B.n416 B.n415 71.676
R1252 B.n417 B.n270 71.676
R1253 B.n424 B.n423 71.676
R1254 B.n425 B.n268 71.676
R1255 B.n432 B.n431 71.676
R1256 B.n435 B.n434 71.676
R1257 B.n380 B.n282 59.5399
R1258 B.n289 B.n288 59.5399
R1259 B.n142 B.n85 59.5399
R1260 B.n163 B.n83 59.5399
R1261 B.n440 B.n260 57.0344
R1262 B.n446 B.n260 57.0344
R1263 B.n446 B.n256 57.0344
R1264 B.n453 B.n256 57.0344
R1265 B.n453 B.n452 57.0344
R1266 B.n459 B.n249 57.0344
R1267 B.n465 B.n249 57.0344
R1268 B.n465 B.n245 57.0344
R1269 B.n471 B.n245 57.0344
R1270 B.n471 B.n241 57.0344
R1271 B.n477 B.n241 57.0344
R1272 B.n477 B.n237 57.0344
R1273 B.n483 B.n237 57.0344
R1274 B.n489 B.n233 57.0344
R1275 B.n489 B.n228 57.0344
R1276 B.n495 B.n228 57.0344
R1277 B.n495 B.n229 57.0344
R1278 B.n502 B.n221 57.0344
R1279 B.n508 B.n221 57.0344
R1280 B.n508 B.n4 57.0344
R1281 B.n595 B.n4 57.0344
R1282 B.n595 B.n594 57.0344
R1283 B.n594 B.n593 57.0344
R1284 B.n593 B.n8 57.0344
R1285 B.n587 B.n8 57.0344
R1286 B.n586 B.n585 57.0344
R1287 B.n585 B.n15 57.0344
R1288 B.n579 B.n15 57.0344
R1289 B.n579 B.n578 57.0344
R1290 B.n577 B.n22 57.0344
R1291 B.n571 B.n22 57.0344
R1292 B.n571 B.n570 57.0344
R1293 B.n570 B.n569 57.0344
R1294 B.n569 B.n29 57.0344
R1295 B.n563 B.n29 57.0344
R1296 B.n563 B.n562 57.0344
R1297 B.n562 B.n561 57.0344
R1298 B.n555 B.n39 57.0344
R1299 B.n555 B.n554 57.0344
R1300 B.n554 B.n553 57.0344
R1301 B.n553 B.n43 57.0344
R1302 B.n547 B.n43 57.0344
R1303 B.n452 B.t5 54.5182
R1304 B.n39 B.t9 54.5182
R1305 B.n229 B.t0 42.7759
R1306 B.t3 B.n586 42.7759
R1307 B.n282 B.n281 34.9096
R1308 B.n288 B.n287 34.9096
R1309 B.n85 B.n84 34.9096
R1310 B.n83 B.n82 34.9096
R1311 B.n549 B.n45 34.1859
R1312 B.n543 B.n542 34.1859
R1313 B.n438 B.n437 34.1859
R1314 B.n442 B.n262 34.1859
R1315 B.t2 B.n233 31.0337
R1316 B.n578 B.t1 31.0337
R1317 B.n483 B.t2 26.0013
R1318 B.t1 B.n577 26.0013
R1319 B B.n597 18.0485
R1320 B.n502 B.t0 14.259
R1321 B.n587 B.t3 14.259
R1322 B.n86 B.n45 10.6151
R1323 B.n89 B.n86 10.6151
R1324 B.n90 B.n89 10.6151
R1325 B.n93 B.n90 10.6151
R1326 B.n94 B.n93 10.6151
R1327 B.n97 B.n94 10.6151
R1328 B.n98 B.n97 10.6151
R1329 B.n101 B.n98 10.6151
R1330 B.n102 B.n101 10.6151
R1331 B.n105 B.n102 10.6151
R1332 B.n106 B.n105 10.6151
R1333 B.n109 B.n106 10.6151
R1334 B.n110 B.n109 10.6151
R1335 B.n113 B.n110 10.6151
R1336 B.n114 B.n113 10.6151
R1337 B.n117 B.n114 10.6151
R1338 B.n118 B.n117 10.6151
R1339 B.n121 B.n118 10.6151
R1340 B.n122 B.n121 10.6151
R1341 B.n125 B.n122 10.6151
R1342 B.n126 B.n125 10.6151
R1343 B.n129 B.n126 10.6151
R1344 B.n130 B.n129 10.6151
R1345 B.n133 B.n130 10.6151
R1346 B.n134 B.n133 10.6151
R1347 B.n137 B.n134 10.6151
R1348 B.n138 B.n137 10.6151
R1349 B.n141 B.n138 10.6151
R1350 B.n146 B.n143 10.6151
R1351 B.n147 B.n146 10.6151
R1352 B.n150 B.n147 10.6151
R1353 B.n151 B.n150 10.6151
R1354 B.n154 B.n151 10.6151
R1355 B.n155 B.n154 10.6151
R1356 B.n158 B.n155 10.6151
R1357 B.n159 B.n158 10.6151
R1358 B.n162 B.n159 10.6151
R1359 B.n167 B.n164 10.6151
R1360 B.n168 B.n167 10.6151
R1361 B.n171 B.n168 10.6151
R1362 B.n172 B.n171 10.6151
R1363 B.n175 B.n172 10.6151
R1364 B.n176 B.n175 10.6151
R1365 B.n179 B.n176 10.6151
R1366 B.n180 B.n179 10.6151
R1367 B.n183 B.n180 10.6151
R1368 B.n184 B.n183 10.6151
R1369 B.n187 B.n184 10.6151
R1370 B.n188 B.n187 10.6151
R1371 B.n191 B.n188 10.6151
R1372 B.n192 B.n191 10.6151
R1373 B.n195 B.n192 10.6151
R1374 B.n196 B.n195 10.6151
R1375 B.n199 B.n196 10.6151
R1376 B.n200 B.n199 10.6151
R1377 B.n203 B.n200 10.6151
R1378 B.n204 B.n203 10.6151
R1379 B.n207 B.n204 10.6151
R1380 B.n208 B.n207 10.6151
R1381 B.n211 B.n208 10.6151
R1382 B.n212 B.n211 10.6151
R1383 B.n215 B.n212 10.6151
R1384 B.n217 B.n215 10.6151
R1385 B.n218 B.n217 10.6151
R1386 B.n543 B.n218 10.6151
R1387 B.n438 B.n258 10.6151
R1388 B.n448 B.n258 10.6151
R1389 B.n449 B.n448 10.6151
R1390 B.n450 B.n449 10.6151
R1391 B.n450 B.n251 10.6151
R1392 B.n461 B.n251 10.6151
R1393 B.n462 B.n461 10.6151
R1394 B.n463 B.n462 10.6151
R1395 B.n463 B.n243 10.6151
R1396 B.n473 B.n243 10.6151
R1397 B.n474 B.n473 10.6151
R1398 B.n475 B.n474 10.6151
R1399 B.n475 B.n235 10.6151
R1400 B.n485 B.n235 10.6151
R1401 B.n486 B.n485 10.6151
R1402 B.n487 B.n486 10.6151
R1403 B.n487 B.n226 10.6151
R1404 B.n497 B.n226 10.6151
R1405 B.n498 B.n497 10.6151
R1406 B.n500 B.n498 10.6151
R1407 B.n500 B.n499 10.6151
R1408 B.n499 B.n219 10.6151
R1409 B.n511 B.n219 10.6151
R1410 B.n512 B.n511 10.6151
R1411 B.n513 B.n512 10.6151
R1412 B.n514 B.n513 10.6151
R1413 B.n516 B.n514 10.6151
R1414 B.n517 B.n516 10.6151
R1415 B.n518 B.n517 10.6151
R1416 B.n519 B.n518 10.6151
R1417 B.n521 B.n519 10.6151
R1418 B.n522 B.n521 10.6151
R1419 B.n523 B.n522 10.6151
R1420 B.n524 B.n523 10.6151
R1421 B.n526 B.n524 10.6151
R1422 B.n527 B.n526 10.6151
R1423 B.n528 B.n527 10.6151
R1424 B.n529 B.n528 10.6151
R1425 B.n531 B.n529 10.6151
R1426 B.n532 B.n531 10.6151
R1427 B.n533 B.n532 10.6151
R1428 B.n534 B.n533 10.6151
R1429 B.n536 B.n534 10.6151
R1430 B.n537 B.n536 10.6151
R1431 B.n538 B.n537 10.6151
R1432 B.n539 B.n538 10.6151
R1433 B.n541 B.n539 10.6151
R1434 B.n542 B.n541 10.6151
R1435 B.n306 B.n262 10.6151
R1436 B.n307 B.n306 10.6151
R1437 B.n308 B.n307 10.6151
R1438 B.n308 B.n302 10.6151
R1439 B.n314 B.n302 10.6151
R1440 B.n315 B.n314 10.6151
R1441 B.n316 B.n315 10.6151
R1442 B.n316 B.n300 10.6151
R1443 B.n322 B.n300 10.6151
R1444 B.n323 B.n322 10.6151
R1445 B.n324 B.n323 10.6151
R1446 B.n324 B.n298 10.6151
R1447 B.n330 B.n298 10.6151
R1448 B.n331 B.n330 10.6151
R1449 B.n332 B.n331 10.6151
R1450 B.n332 B.n296 10.6151
R1451 B.n338 B.n296 10.6151
R1452 B.n339 B.n338 10.6151
R1453 B.n340 B.n339 10.6151
R1454 B.n340 B.n294 10.6151
R1455 B.n346 B.n294 10.6151
R1456 B.n347 B.n346 10.6151
R1457 B.n348 B.n347 10.6151
R1458 B.n348 B.n292 10.6151
R1459 B.n354 B.n292 10.6151
R1460 B.n355 B.n354 10.6151
R1461 B.n356 B.n355 10.6151
R1462 B.n356 B.n290 10.6151
R1463 B.n363 B.n362 10.6151
R1464 B.n364 B.n363 10.6151
R1465 B.n364 B.n285 10.6151
R1466 B.n370 B.n285 10.6151
R1467 B.n371 B.n370 10.6151
R1468 B.n372 B.n371 10.6151
R1469 B.n372 B.n283 10.6151
R1470 B.n378 B.n283 10.6151
R1471 B.n379 B.n378 10.6151
R1472 B.n381 B.n279 10.6151
R1473 B.n387 B.n279 10.6151
R1474 B.n388 B.n387 10.6151
R1475 B.n389 B.n388 10.6151
R1476 B.n389 B.n277 10.6151
R1477 B.n395 B.n277 10.6151
R1478 B.n396 B.n395 10.6151
R1479 B.n397 B.n396 10.6151
R1480 B.n397 B.n275 10.6151
R1481 B.n403 B.n275 10.6151
R1482 B.n404 B.n403 10.6151
R1483 B.n405 B.n404 10.6151
R1484 B.n405 B.n273 10.6151
R1485 B.n411 B.n273 10.6151
R1486 B.n412 B.n411 10.6151
R1487 B.n413 B.n412 10.6151
R1488 B.n413 B.n271 10.6151
R1489 B.n419 B.n271 10.6151
R1490 B.n420 B.n419 10.6151
R1491 B.n421 B.n420 10.6151
R1492 B.n421 B.n269 10.6151
R1493 B.n427 B.n269 10.6151
R1494 B.n428 B.n427 10.6151
R1495 B.n429 B.n428 10.6151
R1496 B.n429 B.n267 10.6151
R1497 B.n267 B.n266 10.6151
R1498 B.n436 B.n266 10.6151
R1499 B.n437 B.n436 10.6151
R1500 B.n443 B.n442 10.6151
R1501 B.n444 B.n443 10.6151
R1502 B.n444 B.n254 10.6151
R1503 B.n455 B.n254 10.6151
R1504 B.n456 B.n455 10.6151
R1505 B.n457 B.n456 10.6151
R1506 B.n457 B.n247 10.6151
R1507 B.n467 B.n247 10.6151
R1508 B.n468 B.n467 10.6151
R1509 B.n469 B.n468 10.6151
R1510 B.n469 B.n239 10.6151
R1511 B.n479 B.n239 10.6151
R1512 B.n480 B.n479 10.6151
R1513 B.n481 B.n480 10.6151
R1514 B.n481 B.n231 10.6151
R1515 B.n491 B.n231 10.6151
R1516 B.n492 B.n491 10.6151
R1517 B.n493 B.n492 10.6151
R1518 B.n493 B.n223 10.6151
R1519 B.n504 B.n223 10.6151
R1520 B.n505 B.n504 10.6151
R1521 B.n506 B.n505 10.6151
R1522 B.n506 B.n0 10.6151
R1523 B.n591 B.n1 10.6151
R1524 B.n591 B.n590 10.6151
R1525 B.n590 B.n589 10.6151
R1526 B.n589 B.n10 10.6151
R1527 B.n583 B.n10 10.6151
R1528 B.n583 B.n582 10.6151
R1529 B.n582 B.n581 10.6151
R1530 B.n581 B.n17 10.6151
R1531 B.n575 B.n17 10.6151
R1532 B.n575 B.n574 10.6151
R1533 B.n574 B.n573 10.6151
R1534 B.n573 B.n24 10.6151
R1535 B.n567 B.n24 10.6151
R1536 B.n567 B.n566 10.6151
R1537 B.n566 B.n565 10.6151
R1538 B.n565 B.n31 10.6151
R1539 B.n559 B.n31 10.6151
R1540 B.n559 B.n558 10.6151
R1541 B.n558 B.n557 10.6151
R1542 B.n557 B.n37 10.6151
R1543 B.n551 B.n37 10.6151
R1544 B.n551 B.n550 10.6151
R1545 B.n550 B.n549 10.6151
R1546 B.n142 B.n141 9.36635
R1547 B.n164 B.n163 9.36635
R1548 B.n290 B.n289 9.36635
R1549 B.n381 B.n380 9.36635
R1550 B.n597 B.n0 2.81026
R1551 B.n597 B.n1 2.81026
R1552 B.n459 B.t5 2.5167
R1553 B.n561 B.t9 2.5167
R1554 B.n143 B.n142 1.24928
R1555 B.n163 B.n162 1.24928
R1556 B.n362 B.n289 1.24928
R1557 B.n380 B.n379 1.24928
R1558 VN.n0 VN.t1 164.535
R1559 VN.n1 VN.t2 164.535
R1560 VN.n0 VN.t3 164.22
R1561 VN.n1 VN.t0 164.22
R1562 VN VN.n1 53.0852
R1563 VN VN.n0 13.1495
R1564 VDD2.n2 VDD2.n0 99.8821
R1565 VDD2.n2 VDD2.n1 64.7536
R1566 VDD2.n1 VDD2.t3 2.52601
R1567 VDD2.n1 VDD2.t1 2.52601
R1568 VDD2.n0 VDD2.t2 2.52601
R1569 VDD2.n0 VDD2.t0 2.52601
R1570 VDD2 VDD2.n2 0.0586897
C0 VDD2 VDD1 0.752352f
C1 VDD1 VP 2.99261f
C2 VTAIL VDD1 4.28541f
C3 VDD2 VN 2.81864f
C4 VN VP 4.60518f
C5 VTAIL VN 2.73296f
C6 VDD2 VP 0.322852f
C7 VTAIL VDD2 4.33204f
C8 VN VDD1 0.148429f
C9 VTAIL VP 2.74706f
C10 VDD2 B 2.809163f
C11 VDD1 B 6.12279f
C12 VTAIL B 6.950037f
C13 VN B 8.360499f
C14 VP B 6.243456f
C15 VDD2.t2 B 0.165376f
C16 VDD2.t0 B 0.165376f
C17 VDD2.n0 B 1.89063f
C18 VDD2.t3 B 0.165376f
C19 VDD2.t1 B 0.165376f
C20 VDD2.n1 B 1.42923f
C21 VDD2.n2 B 2.97941f
C22 VN.t1 B 1.25312f
C23 VN.t3 B 1.25199f
C24 VN.n0 B 0.940937f
C25 VN.t2 B 1.25312f
C26 VN.t0 B 1.25199f
C27 VN.n1 B 2.1352f
C28 VDD1.t0 B 0.167706f
C29 VDD1.t3 B 0.167706f
C30 VDD1.n0 B 1.4497f
C31 VDD1.t2 B 0.167706f
C32 VDD1.t1 B 0.167706f
C33 VDD1.n1 B 1.94128f
C34 VTAIL.n0 B 0.021595f
C35 VTAIL.n1 B 0.016995f
C36 VTAIL.n2 B 0.009401f
C37 VTAIL.n3 B 0.021586f
C38 VTAIL.n4 B 0.00967f
C39 VTAIL.n5 B 0.016995f
C40 VTAIL.n6 B 0.009133f
C41 VTAIL.n7 B 0.021586f
C42 VTAIL.n8 B 0.00967f
C43 VTAIL.n9 B 0.016995f
C44 VTAIL.n10 B 0.009133f
C45 VTAIL.n11 B 0.01619f
C46 VTAIL.n12 B 0.01526f
C47 VTAIL.t3 B 0.036086f
C48 VTAIL.n13 B 0.095407f
C49 VTAIL.n14 B 0.542891f
C50 VTAIL.n15 B 0.009133f
C51 VTAIL.n16 B 0.00967f
C52 VTAIL.n17 B 0.021586f
C53 VTAIL.n18 B 0.021586f
C54 VTAIL.n19 B 0.00967f
C55 VTAIL.n20 B 0.009133f
C56 VTAIL.n21 B 0.016995f
C57 VTAIL.n22 B 0.016995f
C58 VTAIL.n23 B 0.009133f
C59 VTAIL.n24 B 0.00967f
C60 VTAIL.n25 B 0.021586f
C61 VTAIL.n26 B 0.021586f
C62 VTAIL.n27 B 0.00967f
C63 VTAIL.n28 B 0.009133f
C64 VTAIL.n29 B 0.016995f
C65 VTAIL.n30 B 0.016995f
C66 VTAIL.n31 B 0.009133f
C67 VTAIL.n32 B 0.009133f
C68 VTAIL.n33 B 0.00967f
C69 VTAIL.n34 B 0.021586f
C70 VTAIL.n35 B 0.021586f
C71 VTAIL.n36 B 0.042674f
C72 VTAIL.n37 B 0.009401f
C73 VTAIL.n38 B 0.009133f
C74 VTAIL.n39 B 0.040212f
C75 VTAIL.n40 B 0.02349f
C76 VTAIL.n41 B 0.086443f
C77 VTAIL.n42 B 0.021595f
C78 VTAIL.n43 B 0.016995f
C79 VTAIL.n44 B 0.009401f
C80 VTAIL.n45 B 0.021586f
C81 VTAIL.n46 B 0.00967f
C82 VTAIL.n47 B 0.016995f
C83 VTAIL.n48 B 0.009133f
C84 VTAIL.n49 B 0.021586f
C85 VTAIL.n50 B 0.00967f
C86 VTAIL.n51 B 0.016995f
C87 VTAIL.n52 B 0.009133f
C88 VTAIL.n53 B 0.01619f
C89 VTAIL.n54 B 0.01526f
C90 VTAIL.t6 B 0.036086f
C91 VTAIL.n55 B 0.095407f
C92 VTAIL.n56 B 0.542891f
C93 VTAIL.n57 B 0.009133f
C94 VTAIL.n58 B 0.00967f
C95 VTAIL.n59 B 0.021586f
C96 VTAIL.n60 B 0.021586f
C97 VTAIL.n61 B 0.00967f
C98 VTAIL.n62 B 0.009133f
C99 VTAIL.n63 B 0.016995f
C100 VTAIL.n64 B 0.016995f
C101 VTAIL.n65 B 0.009133f
C102 VTAIL.n66 B 0.00967f
C103 VTAIL.n67 B 0.021586f
C104 VTAIL.n68 B 0.021586f
C105 VTAIL.n69 B 0.00967f
C106 VTAIL.n70 B 0.009133f
C107 VTAIL.n71 B 0.016995f
C108 VTAIL.n72 B 0.016995f
C109 VTAIL.n73 B 0.009133f
C110 VTAIL.n74 B 0.009133f
C111 VTAIL.n75 B 0.00967f
C112 VTAIL.n76 B 0.021586f
C113 VTAIL.n77 B 0.021586f
C114 VTAIL.n78 B 0.042674f
C115 VTAIL.n79 B 0.009401f
C116 VTAIL.n80 B 0.009133f
C117 VTAIL.n81 B 0.040212f
C118 VTAIL.n82 B 0.02349f
C119 VTAIL.n83 B 0.125745f
C120 VTAIL.n84 B 0.021595f
C121 VTAIL.n85 B 0.016995f
C122 VTAIL.n86 B 0.009401f
C123 VTAIL.n87 B 0.021586f
C124 VTAIL.n88 B 0.00967f
C125 VTAIL.n89 B 0.016995f
C126 VTAIL.n90 B 0.009133f
C127 VTAIL.n91 B 0.021586f
C128 VTAIL.n92 B 0.00967f
C129 VTAIL.n93 B 0.016995f
C130 VTAIL.n94 B 0.009133f
C131 VTAIL.n95 B 0.01619f
C132 VTAIL.n96 B 0.01526f
C133 VTAIL.t4 B 0.036086f
C134 VTAIL.n97 B 0.095407f
C135 VTAIL.n98 B 0.542891f
C136 VTAIL.n99 B 0.009133f
C137 VTAIL.n100 B 0.00967f
C138 VTAIL.n101 B 0.021586f
C139 VTAIL.n102 B 0.021586f
C140 VTAIL.n103 B 0.00967f
C141 VTAIL.n104 B 0.009133f
C142 VTAIL.n105 B 0.016995f
C143 VTAIL.n106 B 0.016995f
C144 VTAIL.n107 B 0.009133f
C145 VTAIL.n108 B 0.00967f
C146 VTAIL.n109 B 0.021586f
C147 VTAIL.n110 B 0.021586f
C148 VTAIL.n111 B 0.00967f
C149 VTAIL.n112 B 0.009133f
C150 VTAIL.n113 B 0.016995f
C151 VTAIL.n114 B 0.016995f
C152 VTAIL.n115 B 0.009133f
C153 VTAIL.n116 B 0.009133f
C154 VTAIL.n117 B 0.00967f
C155 VTAIL.n118 B 0.021586f
C156 VTAIL.n119 B 0.021586f
C157 VTAIL.n120 B 0.042674f
C158 VTAIL.n121 B 0.009401f
C159 VTAIL.n122 B 0.009133f
C160 VTAIL.n123 B 0.040212f
C161 VTAIL.n124 B 0.02349f
C162 VTAIL.n125 B 0.785972f
C163 VTAIL.n126 B 0.021595f
C164 VTAIL.n127 B 0.016995f
C165 VTAIL.n128 B 0.009401f
C166 VTAIL.n129 B 0.021586f
C167 VTAIL.n130 B 0.009133f
C168 VTAIL.n131 B 0.00967f
C169 VTAIL.n132 B 0.016995f
C170 VTAIL.n133 B 0.009133f
C171 VTAIL.n134 B 0.021586f
C172 VTAIL.n135 B 0.00967f
C173 VTAIL.n136 B 0.016995f
C174 VTAIL.n137 B 0.009133f
C175 VTAIL.n138 B 0.01619f
C176 VTAIL.n139 B 0.01526f
C177 VTAIL.t2 B 0.036086f
C178 VTAIL.n140 B 0.095407f
C179 VTAIL.n141 B 0.542891f
C180 VTAIL.n142 B 0.009133f
C181 VTAIL.n143 B 0.00967f
C182 VTAIL.n144 B 0.021586f
C183 VTAIL.n145 B 0.021586f
C184 VTAIL.n146 B 0.00967f
C185 VTAIL.n147 B 0.009133f
C186 VTAIL.n148 B 0.016995f
C187 VTAIL.n149 B 0.016995f
C188 VTAIL.n150 B 0.009133f
C189 VTAIL.n151 B 0.00967f
C190 VTAIL.n152 B 0.021586f
C191 VTAIL.n153 B 0.021586f
C192 VTAIL.n154 B 0.00967f
C193 VTAIL.n155 B 0.009133f
C194 VTAIL.n156 B 0.016995f
C195 VTAIL.n157 B 0.016995f
C196 VTAIL.n158 B 0.009133f
C197 VTAIL.n159 B 0.00967f
C198 VTAIL.n160 B 0.021586f
C199 VTAIL.n161 B 0.021586f
C200 VTAIL.n162 B 0.042674f
C201 VTAIL.n163 B 0.009401f
C202 VTAIL.n164 B 0.009133f
C203 VTAIL.n165 B 0.040212f
C204 VTAIL.n166 B 0.02349f
C205 VTAIL.n167 B 0.785972f
C206 VTAIL.n168 B 0.021595f
C207 VTAIL.n169 B 0.016995f
C208 VTAIL.n170 B 0.009401f
C209 VTAIL.n171 B 0.021586f
C210 VTAIL.n172 B 0.009133f
C211 VTAIL.n173 B 0.00967f
C212 VTAIL.n174 B 0.016995f
C213 VTAIL.n175 B 0.009133f
C214 VTAIL.n176 B 0.021586f
C215 VTAIL.n177 B 0.00967f
C216 VTAIL.n178 B 0.016995f
C217 VTAIL.n179 B 0.009133f
C218 VTAIL.n180 B 0.01619f
C219 VTAIL.n181 B 0.01526f
C220 VTAIL.t0 B 0.036086f
C221 VTAIL.n182 B 0.095407f
C222 VTAIL.n183 B 0.542891f
C223 VTAIL.n184 B 0.009133f
C224 VTAIL.n185 B 0.00967f
C225 VTAIL.n186 B 0.021586f
C226 VTAIL.n187 B 0.021586f
C227 VTAIL.n188 B 0.00967f
C228 VTAIL.n189 B 0.009133f
C229 VTAIL.n190 B 0.016995f
C230 VTAIL.n191 B 0.016995f
C231 VTAIL.n192 B 0.009133f
C232 VTAIL.n193 B 0.00967f
C233 VTAIL.n194 B 0.021586f
C234 VTAIL.n195 B 0.021586f
C235 VTAIL.n196 B 0.00967f
C236 VTAIL.n197 B 0.009133f
C237 VTAIL.n198 B 0.016995f
C238 VTAIL.n199 B 0.016995f
C239 VTAIL.n200 B 0.009133f
C240 VTAIL.n201 B 0.00967f
C241 VTAIL.n202 B 0.021586f
C242 VTAIL.n203 B 0.021586f
C243 VTAIL.n204 B 0.042674f
C244 VTAIL.n205 B 0.009401f
C245 VTAIL.n206 B 0.009133f
C246 VTAIL.n207 B 0.040212f
C247 VTAIL.n208 B 0.02349f
C248 VTAIL.n209 B 0.125745f
C249 VTAIL.n210 B 0.021595f
C250 VTAIL.n211 B 0.016995f
C251 VTAIL.n212 B 0.009401f
C252 VTAIL.n213 B 0.021586f
C253 VTAIL.n214 B 0.009133f
C254 VTAIL.n215 B 0.00967f
C255 VTAIL.n216 B 0.016995f
C256 VTAIL.n217 B 0.009133f
C257 VTAIL.n218 B 0.021586f
C258 VTAIL.n219 B 0.00967f
C259 VTAIL.n220 B 0.016995f
C260 VTAIL.n221 B 0.009133f
C261 VTAIL.n222 B 0.01619f
C262 VTAIL.n223 B 0.01526f
C263 VTAIL.t5 B 0.036086f
C264 VTAIL.n224 B 0.095407f
C265 VTAIL.n225 B 0.542891f
C266 VTAIL.n226 B 0.009133f
C267 VTAIL.n227 B 0.00967f
C268 VTAIL.n228 B 0.021586f
C269 VTAIL.n229 B 0.021586f
C270 VTAIL.n230 B 0.00967f
C271 VTAIL.n231 B 0.009133f
C272 VTAIL.n232 B 0.016995f
C273 VTAIL.n233 B 0.016995f
C274 VTAIL.n234 B 0.009133f
C275 VTAIL.n235 B 0.00967f
C276 VTAIL.n236 B 0.021586f
C277 VTAIL.n237 B 0.021586f
C278 VTAIL.n238 B 0.00967f
C279 VTAIL.n239 B 0.009133f
C280 VTAIL.n240 B 0.016995f
C281 VTAIL.n241 B 0.016995f
C282 VTAIL.n242 B 0.009133f
C283 VTAIL.n243 B 0.00967f
C284 VTAIL.n244 B 0.021586f
C285 VTAIL.n245 B 0.021586f
C286 VTAIL.n246 B 0.042674f
C287 VTAIL.n247 B 0.009401f
C288 VTAIL.n248 B 0.009133f
C289 VTAIL.n249 B 0.040212f
C290 VTAIL.n250 B 0.02349f
C291 VTAIL.n251 B 0.125745f
C292 VTAIL.n252 B 0.021595f
C293 VTAIL.n253 B 0.016995f
C294 VTAIL.n254 B 0.009401f
C295 VTAIL.n255 B 0.021586f
C296 VTAIL.n256 B 0.009133f
C297 VTAIL.n257 B 0.00967f
C298 VTAIL.n258 B 0.016995f
C299 VTAIL.n259 B 0.009133f
C300 VTAIL.n260 B 0.021586f
C301 VTAIL.n261 B 0.00967f
C302 VTAIL.n262 B 0.016995f
C303 VTAIL.n263 B 0.009133f
C304 VTAIL.n264 B 0.01619f
C305 VTAIL.n265 B 0.01526f
C306 VTAIL.t7 B 0.036086f
C307 VTAIL.n266 B 0.095407f
C308 VTAIL.n267 B 0.542891f
C309 VTAIL.n268 B 0.009133f
C310 VTAIL.n269 B 0.00967f
C311 VTAIL.n270 B 0.021586f
C312 VTAIL.n271 B 0.021586f
C313 VTAIL.n272 B 0.00967f
C314 VTAIL.n273 B 0.009133f
C315 VTAIL.n274 B 0.016995f
C316 VTAIL.n275 B 0.016995f
C317 VTAIL.n276 B 0.009133f
C318 VTAIL.n277 B 0.00967f
C319 VTAIL.n278 B 0.021586f
C320 VTAIL.n279 B 0.021586f
C321 VTAIL.n280 B 0.00967f
C322 VTAIL.n281 B 0.009133f
C323 VTAIL.n282 B 0.016995f
C324 VTAIL.n283 B 0.016995f
C325 VTAIL.n284 B 0.009133f
C326 VTAIL.n285 B 0.00967f
C327 VTAIL.n286 B 0.021586f
C328 VTAIL.n287 B 0.021586f
C329 VTAIL.n288 B 0.042674f
C330 VTAIL.n289 B 0.009401f
C331 VTAIL.n290 B 0.009133f
C332 VTAIL.n291 B 0.040212f
C333 VTAIL.n292 B 0.02349f
C334 VTAIL.n293 B 0.785972f
C335 VTAIL.n294 B 0.021595f
C336 VTAIL.n295 B 0.016995f
C337 VTAIL.n296 B 0.009401f
C338 VTAIL.n297 B 0.021586f
C339 VTAIL.n298 B 0.00967f
C340 VTAIL.n299 B 0.016995f
C341 VTAIL.n300 B 0.009133f
C342 VTAIL.n301 B 0.021586f
C343 VTAIL.n302 B 0.00967f
C344 VTAIL.n303 B 0.016995f
C345 VTAIL.n304 B 0.009133f
C346 VTAIL.n305 B 0.01619f
C347 VTAIL.n306 B 0.01526f
C348 VTAIL.t1 B 0.036086f
C349 VTAIL.n307 B 0.095407f
C350 VTAIL.n308 B 0.542891f
C351 VTAIL.n309 B 0.009133f
C352 VTAIL.n310 B 0.00967f
C353 VTAIL.n311 B 0.021586f
C354 VTAIL.n312 B 0.021586f
C355 VTAIL.n313 B 0.00967f
C356 VTAIL.n314 B 0.009133f
C357 VTAIL.n315 B 0.016995f
C358 VTAIL.n316 B 0.016995f
C359 VTAIL.n317 B 0.009133f
C360 VTAIL.n318 B 0.00967f
C361 VTAIL.n319 B 0.021586f
C362 VTAIL.n320 B 0.021586f
C363 VTAIL.n321 B 0.00967f
C364 VTAIL.n322 B 0.009133f
C365 VTAIL.n323 B 0.016995f
C366 VTAIL.n324 B 0.016995f
C367 VTAIL.n325 B 0.009133f
C368 VTAIL.n326 B 0.009133f
C369 VTAIL.n327 B 0.00967f
C370 VTAIL.n328 B 0.021586f
C371 VTAIL.n329 B 0.021586f
C372 VTAIL.n330 B 0.042674f
C373 VTAIL.n331 B 0.009401f
C374 VTAIL.n332 B 0.009133f
C375 VTAIL.n333 B 0.040212f
C376 VTAIL.n334 B 0.02349f
C377 VTAIL.n335 B 0.740297f
C378 VP.n0 B 0.037408f
C379 VP.t2 B 1.15684f
C380 VP.n1 B 0.054379f
C381 VP.t3 B 1.28446f
C382 VP.t0 B 1.2833f
C383 VP.n2 B 2.16718f
C384 VP.n3 B 1.83692f
C385 VP.t1 B 1.15684f
C386 VP.n4 B 0.507088f
C387 VP.n5 B 0.045398f
C388 VP.n6 B 0.037408f
C389 VP.n7 B 0.037408f
C390 VP.n8 B 0.037408f
C391 VP.n9 B 0.054379f
C392 VP.n10 B 0.045398f
C393 VP.n11 B 0.507088f
C394 VP.n12 B 0.036472f
.ends

