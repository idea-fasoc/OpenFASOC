* NGSPICE file created from diff_pair_sample_1100.ext - technology: sky130A

.subckt diff_pair_sample_1100 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=0 ps=0 w=12.53 l=2.09
X1 B.t8 B.t6 B.t7 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=0 ps=0 w=12.53 l=2.09
X2 VDD1.t1 VP.t0 VTAIL.t3 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=4.8867 ps=25.84 w=12.53 l=2.09
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=4.8867 ps=25.84 w=12.53 l=2.09
X4 B.t5 B.t3 B.t4 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=0 ps=0 w=12.53 l=2.09
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=4.8867 ps=25.84 w=12.53 l=2.09
X6 B.t2 B.t0 B.t1 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=0 ps=0 w=12.53 l=2.09
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n1938_n3474# sky130_fd_pr__pfet_01v8 ad=4.8867 pd=25.84 as=4.8867 ps=25.84 w=12.53 l=2.09
R0 B.n328 B.n89 585
R1 B.n327 B.n326 585
R2 B.n325 B.n90 585
R3 B.n324 B.n323 585
R4 B.n322 B.n91 585
R5 B.n321 B.n320 585
R6 B.n319 B.n92 585
R7 B.n318 B.n317 585
R8 B.n316 B.n93 585
R9 B.n315 B.n314 585
R10 B.n313 B.n94 585
R11 B.n312 B.n311 585
R12 B.n310 B.n95 585
R13 B.n309 B.n308 585
R14 B.n307 B.n96 585
R15 B.n306 B.n305 585
R16 B.n304 B.n97 585
R17 B.n303 B.n302 585
R18 B.n301 B.n98 585
R19 B.n300 B.n299 585
R20 B.n298 B.n99 585
R21 B.n297 B.n296 585
R22 B.n295 B.n100 585
R23 B.n294 B.n293 585
R24 B.n292 B.n101 585
R25 B.n291 B.n290 585
R26 B.n289 B.n102 585
R27 B.n288 B.n287 585
R28 B.n286 B.n103 585
R29 B.n285 B.n284 585
R30 B.n283 B.n104 585
R31 B.n282 B.n281 585
R32 B.n280 B.n105 585
R33 B.n279 B.n278 585
R34 B.n277 B.n106 585
R35 B.n276 B.n275 585
R36 B.n274 B.n107 585
R37 B.n273 B.n272 585
R38 B.n271 B.n108 585
R39 B.n270 B.n269 585
R40 B.n268 B.n109 585
R41 B.n267 B.n266 585
R42 B.n265 B.n110 585
R43 B.n263 B.n262 585
R44 B.n261 B.n113 585
R45 B.n260 B.n259 585
R46 B.n258 B.n114 585
R47 B.n257 B.n256 585
R48 B.n255 B.n115 585
R49 B.n254 B.n253 585
R50 B.n252 B.n116 585
R51 B.n251 B.n250 585
R52 B.n249 B.n117 585
R53 B.n248 B.n247 585
R54 B.n243 B.n118 585
R55 B.n242 B.n241 585
R56 B.n240 B.n119 585
R57 B.n239 B.n238 585
R58 B.n237 B.n120 585
R59 B.n236 B.n235 585
R60 B.n234 B.n121 585
R61 B.n233 B.n232 585
R62 B.n231 B.n122 585
R63 B.n230 B.n229 585
R64 B.n228 B.n123 585
R65 B.n227 B.n226 585
R66 B.n225 B.n124 585
R67 B.n224 B.n223 585
R68 B.n222 B.n125 585
R69 B.n221 B.n220 585
R70 B.n219 B.n126 585
R71 B.n218 B.n217 585
R72 B.n216 B.n127 585
R73 B.n215 B.n214 585
R74 B.n213 B.n128 585
R75 B.n212 B.n211 585
R76 B.n210 B.n129 585
R77 B.n209 B.n208 585
R78 B.n207 B.n130 585
R79 B.n206 B.n205 585
R80 B.n204 B.n131 585
R81 B.n203 B.n202 585
R82 B.n201 B.n132 585
R83 B.n200 B.n199 585
R84 B.n198 B.n133 585
R85 B.n197 B.n196 585
R86 B.n195 B.n134 585
R87 B.n194 B.n193 585
R88 B.n192 B.n135 585
R89 B.n191 B.n190 585
R90 B.n189 B.n136 585
R91 B.n188 B.n187 585
R92 B.n186 B.n137 585
R93 B.n185 B.n184 585
R94 B.n183 B.n138 585
R95 B.n182 B.n181 585
R96 B.n330 B.n329 585
R97 B.n331 B.n88 585
R98 B.n333 B.n332 585
R99 B.n334 B.n87 585
R100 B.n336 B.n335 585
R101 B.n337 B.n86 585
R102 B.n339 B.n338 585
R103 B.n340 B.n85 585
R104 B.n342 B.n341 585
R105 B.n343 B.n84 585
R106 B.n345 B.n344 585
R107 B.n346 B.n83 585
R108 B.n348 B.n347 585
R109 B.n349 B.n82 585
R110 B.n351 B.n350 585
R111 B.n352 B.n81 585
R112 B.n354 B.n353 585
R113 B.n355 B.n80 585
R114 B.n357 B.n356 585
R115 B.n358 B.n79 585
R116 B.n360 B.n359 585
R117 B.n361 B.n78 585
R118 B.n363 B.n362 585
R119 B.n364 B.n77 585
R120 B.n366 B.n365 585
R121 B.n367 B.n76 585
R122 B.n369 B.n368 585
R123 B.n370 B.n75 585
R124 B.n372 B.n371 585
R125 B.n373 B.n74 585
R126 B.n375 B.n374 585
R127 B.n376 B.n73 585
R128 B.n378 B.n377 585
R129 B.n379 B.n72 585
R130 B.n381 B.n380 585
R131 B.n382 B.n71 585
R132 B.n384 B.n383 585
R133 B.n385 B.n70 585
R134 B.n387 B.n386 585
R135 B.n388 B.n69 585
R136 B.n390 B.n389 585
R137 B.n391 B.n68 585
R138 B.n393 B.n392 585
R139 B.n394 B.n67 585
R140 B.n396 B.n395 585
R141 B.n397 B.n66 585
R142 B.n542 B.n13 585
R143 B.n541 B.n540 585
R144 B.n539 B.n14 585
R145 B.n538 B.n537 585
R146 B.n536 B.n15 585
R147 B.n535 B.n534 585
R148 B.n533 B.n16 585
R149 B.n532 B.n531 585
R150 B.n530 B.n17 585
R151 B.n529 B.n528 585
R152 B.n527 B.n18 585
R153 B.n526 B.n525 585
R154 B.n524 B.n19 585
R155 B.n523 B.n522 585
R156 B.n521 B.n20 585
R157 B.n520 B.n519 585
R158 B.n518 B.n21 585
R159 B.n517 B.n516 585
R160 B.n515 B.n22 585
R161 B.n514 B.n513 585
R162 B.n512 B.n23 585
R163 B.n511 B.n510 585
R164 B.n509 B.n24 585
R165 B.n508 B.n507 585
R166 B.n506 B.n25 585
R167 B.n505 B.n504 585
R168 B.n503 B.n26 585
R169 B.n502 B.n501 585
R170 B.n500 B.n27 585
R171 B.n499 B.n498 585
R172 B.n497 B.n28 585
R173 B.n496 B.n495 585
R174 B.n494 B.n29 585
R175 B.n493 B.n492 585
R176 B.n491 B.n30 585
R177 B.n490 B.n489 585
R178 B.n488 B.n31 585
R179 B.n487 B.n486 585
R180 B.n485 B.n32 585
R181 B.n484 B.n483 585
R182 B.n482 B.n33 585
R183 B.n481 B.n480 585
R184 B.n479 B.n34 585
R185 B.n478 B.n477 585
R186 B.n476 B.n35 585
R187 B.n475 B.n474 585
R188 B.n473 B.n39 585
R189 B.n472 B.n471 585
R190 B.n470 B.n40 585
R191 B.n469 B.n468 585
R192 B.n467 B.n41 585
R193 B.n466 B.n465 585
R194 B.n464 B.n42 585
R195 B.n462 B.n461 585
R196 B.n460 B.n45 585
R197 B.n459 B.n458 585
R198 B.n457 B.n46 585
R199 B.n456 B.n455 585
R200 B.n454 B.n47 585
R201 B.n453 B.n452 585
R202 B.n451 B.n48 585
R203 B.n450 B.n449 585
R204 B.n448 B.n49 585
R205 B.n447 B.n446 585
R206 B.n445 B.n50 585
R207 B.n444 B.n443 585
R208 B.n442 B.n51 585
R209 B.n441 B.n440 585
R210 B.n439 B.n52 585
R211 B.n438 B.n437 585
R212 B.n436 B.n53 585
R213 B.n435 B.n434 585
R214 B.n433 B.n54 585
R215 B.n432 B.n431 585
R216 B.n430 B.n55 585
R217 B.n429 B.n428 585
R218 B.n427 B.n56 585
R219 B.n426 B.n425 585
R220 B.n424 B.n57 585
R221 B.n423 B.n422 585
R222 B.n421 B.n58 585
R223 B.n420 B.n419 585
R224 B.n418 B.n59 585
R225 B.n417 B.n416 585
R226 B.n415 B.n60 585
R227 B.n414 B.n413 585
R228 B.n412 B.n61 585
R229 B.n411 B.n410 585
R230 B.n409 B.n62 585
R231 B.n408 B.n407 585
R232 B.n406 B.n63 585
R233 B.n405 B.n404 585
R234 B.n403 B.n64 585
R235 B.n402 B.n401 585
R236 B.n400 B.n65 585
R237 B.n399 B.n398 585
R238 B.n544 B.n543 585
R239 B.n545 B.n12 585
R240 B.n547 B.n546 585
R241 B.n548 B.n11 585
R242 B.n550 B.n549 585
R243 B.n551 B.n10 585
R244 B.n553 B.n552 585
R245 B.n554 B.n9 585
R246 B.n556 B.n555 585
R247 B.n557 B.n8 585
R248 B.n559 B.n558 585
R249 B.n560 B.n7 585
R250 B.n562 B.n561 585
R251 B.n563 B.n6 585
R252 B.n565 B.n564 585
R253 B.n566 B.n5 585
R254 B.n568 B.n567 585
R255 B.n569 B.n4 585
R256 B.n571 B.n570 585
R257 B.n572 B.n3 585
R258 B.n574 B.n573 585
R259 B.n575 B.n0 585
R260 B.n2 B.n1 585
R261 B.n150 B.n149 585
R262 B.n152 B.n151 585
R263 B.n153 B.n148 585
R264 B.n155 B.n154 585
R265 B.n156 B.n147 585
R266 B.n158 B.n157 585
R267 B.n159 B.n146 585
R268 B.n161 B.n160 585
R269 B.n162 B.n145 585
R270 B.n164 B.n163 585
R271 B.n165 B.n144 585
R272 B.n167 B.n166 585
R273 B.n168 B.n143 585
R274 B.n170 B.n169 585
R275 B.n171 B.n142 585
R276 B.n173 B.n172 585
R277 B.n174 B.n141 585
R278 B.n176 B.n175 585
R279 B.n177 B.n140 585
R280 B.n179 B.n178 585
R281 B.n180 B.n139 585
R282 B.n181 B.n180 468.476
R283 B.n329 B.n328 468.476
R284 B.n399 B.n66 468.476
R285 B.n544 B.n13 468.476
R286 B.n244 B.t3 351.606
R287 B.n111 B.t9 351.606
R288 B.n43 B.t6 351.606
R289 B.n36 B.t0 351.606
R290 B.n577 B.n576 256.663
R291 B.n576 B.n575 235.042
R292 B.n576 B.n2 235.042
R293 B.n181 B.n138 163.367
R294 B.n185 B.n138 163.367
R295 B.n186 B.n185 163.367
R296 B.n187 B.n186 163.367
R297 B.n187 B.n136 163.367
R298 B.n191 B.n136 163.367
R299 B.n192 B.n191 163.367
R300 B.n193 B.n192 163.367
R301 B.n193 B.n134 163.367
R302 B.n197 B.n134 163.367
R303 B.n198 B.n197 163.367
R304 B.n199 B.n198 163.367
R305 B.n199 B.n132 163.367
R306 B.n203 B.n132 163.367
R307 B.n204 B.n203 163.367
R308 B.n205 B.n204 163.367
R309 B.n205 B.n130 163.367
R310 B.n209 B.n130 163.367
R311 B.n210 B.n209 163.367
R312 B.n211 B.n210 163.367
R313 B.n211 B.n128 163.367
R314 B.n215 B.n128 163.367
R315 B.n216 B.n215 163.367
R316 B.n217 B.n216 163.367
R317 B.n217 B.n126 163.367
R318 B.n221 B.n126 163.367
R319 B.n222 B.n221 163.367
R320 B.n223 B.n222 163.367
R321 B.n223 B.n124 163.367
R322 B.n227 B.n124 163.367
R323 B.n228 B.n227 163.367
R324 B.n229 B.n228 163.367
R325 B.n229 B.n122 163.367
R326 B.n233 B.n122 163.367
R327 B.n234 B.n233 163.367
R328 B.n235 B.n234 163.367
R329 B.n235 B.n120 163.367
R330 B.n239 B.n120 163.367
R331 B.n240 B.n239 163.367
R332 B.n241 B.n240 163.367
R333 B.n241 B.n118 163.367
R334 B.n248 B.n118 163.367
R335 B.n249 B.n248 163.367
R336 B.n250 B.n249 163.367
R337 B.n250 B.n116 163.367
R338 B.n254 B.n116 163.367
R339 B.n255 B.n254 163.367
R340 B.n256 B.n255 163.367
R341 B.n256 B.n114 163.367
R342 B.n260 B.n114 163.367
R343 B.n261 B.n260 163.367
R344 B.n262 B.n261 163.367
R345 B.n262 B.n110 163.367
R346 B.n267 B.n110 163.367
R347 B.n268 B.n267 163.367
R348 B.n269 B.n268 163.367
R349 B.n269 B.n108 163.367
R350 B.n273 B.n108 163.367
R351 B.n274 B.n273 163.367
R352 B.n275 B.n274 163.367
R353 B.n275 B.n106 163.367
R354 B.n279 B.n106 163.367
R355 B.n280 B.n279 163.367
R356 B.n281 B.n280 163.367
R357 B.n281 B.n104 163.367
R358 B.n285 B.n104 163.367
R359 B.n286 B.n285 163.367
R360 B.n287 B.n286 163.367
R361 B.n287 B.n102 163.367
R362 B.n291 B.n102 163.367
R363 B.n292 B.n291 163.367
R364 B.n293 B.n292 163.367
R365 B.n293 B.n100 163.367
R366 B.n297 B.n100 163.367
R367 B.n298 B.n297 163.367
R368 B.n299 B.n298 163.367
R369 B.n299 B.n98 163.367
R370 B.n303 B.n98 163.367
R371 B.n304 B.n303 163.367
R372 B.n305 B.n304 163.367
R373 B.n305 B.n96 163.367
R374 B.n309 B.n96 163.367
R375 B.n310 B.n309 163.367
R376 B.n311 B.n310 163.367
R377 B.n311 B.n94 163.367
R378 B.n315 B.n94 163.367
R379 B.n316 B.n315 163.367
R380 B.n317 B.n316 163.367
R381 B.n317 B.n92 163.367
R382 B.n321 B.n92 163.367
R383 B.n322 B.n321 163.367
R384 B.n323 B.n322 163.367
R385 B.n323 B.n90 163.367
R386 B.n327 B.n90 163.367
R387 B.n328 B.n327 163.367
R388 B.n395 B.n66 163.367
R389 B.n395 B.n394 163.367
R390 B.n394 B.n393 163.367
R391 B.n393 B.n68 163.367
R392 B.n389 B.n68 163.367
R393 B.n389 B.n388 163.367
R394 B.n388 B.n387 163.367
R395 B.n387 B.n70 163.367
R396 B.n383 B.n70 163.367
R397 B.n383 B.n382 163.367
R398 B.n382 B.n381 163.367
R399 B.n381 B.n72 163.367
R400 B.n377 B.n72 163.367
R401 B.n377 B.n376 163.367
R402 B.n376 B.n375 163.367
R403 B.n375 B.n74 163.367
R404 B.n371 B.n74 163.367
R405 B.n371 B.n370 163.367
R406 B.n370 B.n369 163.367
R407 B.n369 B.n76 163.367
R408 B.n365 B.n76 163.367
R409 B.n365 B.n364 163.367
R410 B.n364 B.n363 163.367
R411 B.n363 B.n78 163.367
R412 B.n359 B.n78 163.367
R413 B.n359 B.n358 163.367
R414 B.n358 B.n357 163.367
R415 B.n357 B.n80 163.367
R416 B.n353 B.n80 163.367
R417 B.n353 B.n352 163.367
R418 B.n352 B.n351 163.367
R419 B.n351 B.n82 163.367
R420 B.n347 B.n82 163.367
R421 B.n347 B.n346 163.367
R422 B.n346 B.n345 163.367
R423 B.n345 B.n84 163.367
R424 B.n341 B.n84 163.367
R425 B.n341 B.n340 163.367
R426 B.n340 B.n339 163.367
R427 B.n339 B.n86 163.367
R428 B.n335 B.n86 163.367
R429 B.n335 B.n334 163.367
R430 B.n334 B.n333 163.367
R431 B.n333 B.n88 163.367
R432 B.n329 B.n88 163.367
R433 B.n540 B.n13 163.367
R434 B.n540 B.n539 163.367
R435 B.n539 B.n538 163.367
R436 B.n538 B.n15 163.367
R437 B.n534 B.n15 163.367
R438 B.n534 B.n533 163.367
R439 B.n533 B.n532 163.367
R440 B.n532 B.n17 163.367
R441 B.n528 B.n17 163.367
R442 B.n528 B.n527 163.367
R443 B.n527 B.n526 163.367
R444 B.n526 B.n19 163.367
R445 B.n522 B.n19 163.367
R446 B.n522 B.n521 163.367
R447 B.n521 B.n520 163.367
R448 B.n520 B.n21 163.367
R449 B.n516 B.n21 163.367
R450 B.n516 B.n515 163.367
R451 B.n515 B.n514 163.367
R452 B.n514 B.n23 163.367
R453 B.n510 B.n23 163.367
R454 B.n510 B.n509 163.367
R455 B.n509 B.n508 163.367
R456 B.n508 B.n25 163.367
R457 B.n504 B.n25 163.367
R458 B.n504 B.n503 163.367
R459 B.n503 B.n502 163.367
R460 B.n502 B.n27 163.367
R461 B.n498 B.n27 163.367
R462 B.n498 B.n497 163.367
R463 B.n497 B.n496 163.367
R464 B.n496 B.n29 163.367
R465 B.n492 B.n29 163.367
R466 B.n492 B.n491 163.367
R467 B.n491 B.n490 163.367
R468 B.n490 B.n31 163.367
R469 B.n486 B.n31 163.367
R470 B.n486 B.n485 163.367
R471 B.n485 B.n484 163.367
R472 B.n484 B.n33 163.367
R473 B.n480 B.n33 163.367
R474 B.n480 B.n479 163.367
R475 B.n479 B.n478 163.367
R476 B.n478 B.n35 163.367
R477 B.n474 B.n35 163.367
R478 B.n474 B.n473 163.367
R479 B.n473 B.n472 163.367
R480 B.n472 B.n40 163.367
R481 B.n468 B.n40 163.367
R482 B.n468 B.n467 163.367
R483 B.n467 B.n466 163.367
R484 B.n466 B.n42 163.367
R485 B.n461 B.n42 163.367
R486 B.n461 B.n460 163.367
R487 B.n460 B.n459 163.367
R488 B.n459 B.n46 163.367
R489 B.n455 B.n46 163.367
R490 B.n455 B.n454 163.367
R491 B.n454 B.n453 163.367
R492 B.n453 B.n48 163.367
R493 B.n449 B.n48 163.367
R494 B.n449 B.n448 163.367
R495 B.n448 B.n447 163.367
R496 B.n447 B.n50 163.367
R497 B.n443 B.n50 163.367
R498 B.n443 B.n442 163.367
R499 B.n442 B.n441 163.367
R500 B.n441 B.n52 163.367
R501 B.n437 B.n52 163.367
R502 B.n437 B.n436 163.367
R503 B.n436 B.n435 163.367
R504 B.n435 B.n54 163.367
R505 B.n431 B.n54 163.367
R506 B.n431 B.n430 163.367
R507 B.n430 B.n429 163.367
R508 B.n429 B.n56 163.367
R509 B.n425 B.n56 163.367
R510 B.n425 B.n424 163.367
R511 B.n424 B.n423 163.367
R512 B.n423 B.n58 163.367
R513 B.n419 B.n58 163.367
R514 B.n419 B.n418 163.367
R515 B.n418 B.n417 163.367
R516 B.n417 B.n60 163.367
R517 B.n413 B.n60 163.367
R518 B.n413 B.n412 163.367
R519 B.n412 B.n411 163.367
R520 B.n411 B.n62 163.367
R521 B.n407 B.n62 163.367
R522 B.n407 B.n406 163.367
R523 B.n406 B.n405 163.367
R524 B.n405 B.n64 163.367
R525 B.n401 B.n64 163.367
R526 B.n401 B.n400 163.367
R527 B.n400 B.n399 163.367
R528 B.n545 B.n544 163.367
R529 B.n546 B.n545 163.367
R530 B.n546 B.n11 163.367
R531 B.n550 B.n11 163.367
R532 B.n551 B.n550 163.367
R533 B.n552 B.n551 163.367
R534 B.n552 B.n9 163.367
R535 B.n556 B.n9 163.367
R536 B.n557 B.n556 163.367
R537 B.n558 B.n557 163.367
R538 B.n558 B.n7 163.367
R539 B.n562 B.n7 163.367
R540 B.n563 B.n562 163.367
R541 B.n564 B.n563 163.367
R542 B.n564 B.n5 163.367
R543 B.n568 B.n5 163.367
R544 B.n569 B.n568 163.367
R545 B.n570 B.n569 163.367
R546 B.n570 B.n3 163.367
R547 B.n574 B.n3 163.367
R548 B.n575 B.n574 163.367
R549 B.n150 B.n2 163.367
R550 B.n151 B.n150 163.367
R551 B.n151 B.n148 163.367
R552 B.n155 B.n148 163.367
R553 B.n156 B.n155 163.367
R554 B.n157 B.n156 163.367
R555 B.n157 B.n146 163.367
R556 B.n161 B.n146 163.367
R557 B.n162 B.n161 163.367
R558 B.n163 B.n162 163.367
R559 B.n163 B.n144 163.367
R560 B.n167 B.n144 163.367
R561 B.n168 B.n167 163.367
R562 B.n169 B.n168 163.367
R563 B.n169 B.n142 163.367
R564 B.n173 B.n142 163.367
R565 B.n174 B.n173 163.367
R566 B.n175 B.n174 163.367
R567 B.n175 B.n140 163.367
R568 B.n179 B.n140 163.367
R569 B.n180 B.n179 163.367
R570 B.n111 B.t10 159.547
R571 B.n43 B.t8 159.547
R572 B.n244 B.t4 159.531
R573 B.n36 B.t2 159.531
R574 B.n112 B.t11 112.614
R575 B.n44 B.t7 112.614
R576 B.n245 B.t5 112.599
R577 B.n37 B.t1 112.599
R578 B.n246 B.n245 59.5399
R579 B.n264 B.n112 59.5399
R580 B.n463 B.n44 59.5399
R581 B.n38 B.n37 59.5399
R582 B.n245 B.n244 46.9338
R583 B.n112 B.n111 46.9338
R584 B.n44 B.n43 46.9338
R585 B.n37 B.n36 46.9338
R586 B.n543 B.n542 30.4395
R587 B.n398 B.n397 30.4395
R588 B.n330 B.n89 30.4395
R589 B.n182 B.n139 30.4395
R590 B B.n577 18.0485
R591 B.n543 B.n12 10.6151
R592 B.n547 B.n12 10.6151
R593 B.n548 B.n547 10.6151
R594 B.n549 B.n548 10.6151
R595 B.n549 B.n10 10.6151
R596 B.n553 B.n10 10.6151
R597 B.n554 B.n553 10.6151
R598 B.n555 B.n554 10.6151
R599 B.n555 B.n8 10.6151
R600 B.n559 B.n8 10.6151
R601 B.n560 B.n559 10.6151
R602 B.n561 B.n560 10.6151
R603 B.n561 B.n6 10.6151
R604 B.n565 B.n6 10.6151
R605 B.n566 B.n565 10.6151
R606 B.n567 B.n566 10.6151
R607 B.n567 B.n4 10.6151
R608 B.n571 B.n4 10.6151
R609 B.n572 B.n571 10.6151
R610 B.n573 B.n572 10.6151
R611 B.n573 B.n0 10.6151
R612 B.n542 B.n541 10.6151
R613 B.n541 B.n14 10.6151
R614 B.n537 B.n14 10.6151
R615 B.n537 B.n536 10.6151
R616 B.n536 B.n535 10.6151
R617 B.n535 B.n16 10.6151
R618 B.n531 B.n16 10.6151
R619 B.n531 B.n530 10.6151
R620 B.n530 B.n529 10.6151
R621 B.n529 B.n18 10.6151
R622 B.n525 B.n18 10.6151
R623 B.n525 B.n524 10.6151
R624 B.n524 B.n523 10.6151
R625 B.n523 B.n20 10.6151
R626 B.n519 B.n20 10.6151
R627 B.n519 B.n518 10.6151
R628 B.n518 B.n517 10.6151
R629 B.n517 B.n22 10.6151
R630 B.n513 B.n22 10.6151
R631 B.n513 B.n512 10.6151
R632 B.n512 B.n511 10.6151
R633 B.n511 B.n24 10.6151
R634 B.n507 B.n24 10.6151
R635 B.n507 B.n506 10.6151
R636 B.n506 B.n505 10.6151
R637 B.n505 B.n26 10.6151
R638 B.n501 B.n26 10.6151
R639 B.n501 B.n500 10.6151
R640 B.n500 B.n499 10.6151
R641 B.n499 B.n28 10.6151
R642 B.n495 B.n28 10.6151
R643 B.n495 B.n494 10.6151
R644 B.n494 B.n493 10.6151
R645 B.n493 B.n30 10.6151
R646 B.n489 B.n30 10.6151
R647 B.n489 B.n488 10.6151
R648 B.n488 B.n487 10.6151
R649 B.n487 B.n32 10.6151
R650 B.n483 B.n32 10.6151
R651 B.n483 B.n482 10.6151
R652 B.n482 B.n481 10.6151
R653 B.n481 B.n34 10.6151
R654 B.n477 B.n476 10.6151
R655 B.n476 B.n475 10.6151
R656 B.n475 B.n39 10.6151
R657 B.n471 B.n39 10.6151
R658 B.n471 B.n470 10.6151
R659 B.n470 B.n469 10.6151
R660 B.n469 B.n41 10.6151
R661 B.n465 B.n41 10.6151
R662 B.n465 B.n464 10.6151
R663 B.n462 B.n45 10.6151
R664 B.n458 B.n45 10.6151
R665 B.n458 B.n457 10.6151
R666 B.n457 B.n456 10.6151
R667 B.n456 B.n47 10.6151
R668 B.n452 B.n47 10.6151
R669 B.n452 B.n451 10.6151
R670 B.n451 B.n450 10.6151
R671 B.n450 B.n49 10.6151
R672 B.n446 B.n49 10.6151
R673 B.n446 B.n445 10.6151
R674 B.n445 B.n444 10.6151
R675 B.n444 B.n51 10.6151
R676 B.n440 B.n51 10.6151
R677 B.n440 B.n439 10.6151
R678 B.n439 B.n438 10.6151
R679 B.n438 B.n53 10.6151
R680 B.n434 B.n53 10.6151
R681 B.n434 B.n433 10.6151
R682 B.n433 B.n432 10.6151
R683 B.n432 B.n55 10.6151
R684 B.n428 B.n55 10.6151
R685 B.n428 B.n427 10.6151
R686 B.n427 B.n426 10.6151
R687 B.n426 B.n57 10.6151
R688 B.n422 B.n57 10.6151
R689 B.n422 B.n421 10.6151
R690 B.n421 B.n420 10.6151
R691 B.n420 B.n59 10.6151
R692 B.n416 B.n59 10.6151
R693 B.n416 B.n415 10.6151
R694 B.n415 B.n414 10.6151
R695 B.n414 B.n61 10.6151
R696 B.n410 B.n61 10.6151
R697 B.n410 B.n409 10.6151
R698 B.n409 B.n408 10.6151
R699 B.n408 B.n63 10.6151
R700 B.n404 B.n63 10.6151
R701 B.n404 B.n403 10.6151
R702 B.n403 B.n402 10.6151
R703 B.n402 B.n65 10.6151
R704 B.n398 B.n65 10.6151
R705 B.n397 B.n396 10.6151
R706 B.n396 B.n67 10.6151
R707 B.n392 B.n67 10.6151
R708 B.n392 B.n391 10.6151
R709 B.n391 B.n390 10.6151
R710 B.n390 B.n69 10.6151
R711 B.n386 B.n69 10.6151
R712 B.n386 B.n385 10.6151
R713 B.n385 B.n384 10.6151
R714 B.n384 B.n71 10.6151
R715 B.n380 B.n71 10.6151
R716 B.n380 B.n379 10.6151
R717 B.n379 B.n378 10.6151
R718 B.n378 B.n73 10.6151
R719 B.n374 B.n73 10.6151
R720 B.n374 B.n373 10.6151
R721 B.n373 B.n372 10.6151
R722 B.n372 B.n75 10.6151
R723 B.n368 B.n75 10.6151
R724 B.n368 B.n367 10.6151
R725 B.n367 B.n366 10.6151
R726 B.n366 B.n77 10.6151
R727 B.n362 B.n77 10.6151
R728 B.n362 B.n361 10.6151
R729 B.n361 B.n360 10.6151
R730 B.n360 B.n79 10.6151
R731 B.n356 B.n79 10.6151
R732 B.n356 B.n355 10.6151
R733 B.n355 B.n354 10.6151
R734 B.n354 B.n81 10.6151
R735 B.n350 B.n81 10.6151
R736 B.n350 B.n349 10.6151
R737 B.n349 B.n348 10.6151
R738 B.n348 B.n83 10.6151
R739 B.n344 B.n83 10.6151
R740 B.n344 B.n343 10.6151
R741 B.n343 B.n342 10.6151
R742 B.n342 B.n85 10.6151
R743 B.n338 B.n85 10.6151
R744 B.n338 B.n337 10.6151
R745 B.n337 B.n336 10.6151
R746 B.n336 B.n87 10.6151
R747 B.n332 B.n87 10.6151
R748 B.n332 B.n331 10.6151
R749 B.n331 B.n330 10.6151
R750 B.n149 B.n1 10.6151
R751 B.n152 B.n149 10.6151
R752 B.n153 B.n152 10.6151
R753 B.n154 B.n153 10.6151
R754 B.n154 B.n147 10.6151
R755 B.n158 B.n147 10.6151
R756 B.n159 B.n158 10.6151
R757 B.n160 B.n159 10.6151
R758 B.n160 B.n145 10.6151
R759 B.n164 B.n145 10.6151
R760 B.n165 B.n164 10.6151
R761 B.n166 B.n165 10.6151
R762 B.n166 B.n143 10.6151
R763 B.n170 B.n143 10.6151
R764 B.n171 B.n170 10.6151
R765 B.n172 B.n171 10.6151
R766 B.n172 B.n141 10.6151
R767 B.n176 B.n141 10.6151
R768 B.n177 B.n176 10.6151
R769 B.n178 B.n177 10.6151
R770 B.n178 B.n139 10.6151
R771 B.n183 B.n182 10.6151
R772 B.n184 B.n183 10.6151
R773 B.n184 B.n137 10.6151
R774 B.n188 B.n137 10.6151
R775 B.n189 B.n188 10.6151
R776 B.n190 B.n189 10.6151
R777 B.n190 B.n135 10.6151
R778 B.n194 B.n135 10.6151
R779 B.n195 B.n194 10.6151
R780 B.n196 B.n195 10.6151
R781 B.n196 B.n133 10.6151
R782 B.n200 B.n133 10.6151
R783 B.n201 B.n200 10.6151
R784 B.n202 B.n201 10.6151
R785 B.n202 B.n131 10.6151
R786 B.n206 B.n131 10.6151
R787 B.n207 B.n206 10.6151
R788 B.n208 B.n207 10.6151
R789 B.n208 B.n129 10.6151
R790 B.n212 B.n129 10.6151
R791 B.n213 B.n212 10.6151
R792 B.n214 B.n213 10.6151
R793 B.n214 B.n127 10.6151
R794 B.n218 B.n127 10.6151
R795 B.n219 B.n218 10.6151
R796 B.n220 B.n219 10.6151
R797 B.n220 B.n125 10.6151
R798 B.n224 B.n125 10.6151
R799 B.n225 B.n224 10.6151
R800 B.n226 B.n225 10.6151
R801 B.n226 B.n123 10.6151
R802 B.n230 B.n123 10.6151
R803 B.n231 B.n230 10.6151
R804 B.n232 B.n231 10.6151
R805 B.n232 B.n121 10.6151
R806 B.n236 B.n121 10.6151
R807 B.n237 B.n236 10.6151
R808 B.n238 B.n237 10.6151
R809 B.n238 B.n119 10.6151
R810 B.n242 B.n119 10.6151
R811 B.n243 B.n242 10.6151
R812 B.n247 B.n243 10.6151
R813 B.n251 B.n117 10.6151
R814 B.n252 B.n251 10.6151
R815 B.n253 B.n252 10.6151
R816 B.n253 B.n115 10.6151
R817 B.n257 B.n115 10.6151
R818 B.n258 B.n257 10.6151
R819 B.n259 B.n258 10.6151
R820 B.n259 B.n113 10.6151
R821 B.n263 B.n113 10.6151
R822 B.n266 B.n265 10.6151
R823 B.n266 B.n109 10.6151
R824 B.n270 B.n109 10.6151
R825 B.n271 B.n270 10.6151
R826 B.n272 B.n271 10.6151
R827 B.n272 B.n107 10.6151
R828 B.n276 B.n107 10.6151
R829 B.n277 B.n276 10.6151
R830 B.n278 B.n277 10.6151
R831 B.n278 B.n105 10.6151
R832 B.n282 B.n105 10.6151
R833 B.n283 B.n282 10.6151
R834 B.n284 B.n283 10.6151
R835 B.n284 B.n103 10.6151
R836 B.n288 B.n103 10.6151
R837 B.n289 B.n288 10.6151
R838 B.n290 B.n289 10.6151
R839 B.n290 B.n101 10.6151
R840 B.n294 B.n101 10.6151
R841 B.n295 B.n294 10.6151
R842 B.n296 B.n295 10.6151
R843 B.n296 B.n99 10.6151
R844 B.n300 B.n99 10.6151
R845 B.n301 B.n300 10.6151
R846 B.n302 B.n301 10.6151
R847 B.n302 B.n97 10.6151
R848 B.n306 B.n97 10.6151
R849 B.n307 B.n306 10.6151
R850 B.n308 B.n307 10.6151
R851 B.n308 B.n95 10.6151
R852 B.n312 B.n95 10.6151
R853 B.n313 B.n312 10.6151
R854 B.n314 B.n313 10.6151
R855 B.n314 B.n93 10.6151
R856 B.n318 B.n93 10.6151
R857 B.n319 B.n318 10.6151
R858 B.n320 B.n319 10.6151
R859 B.n320 B.n91 10.6151
R860 B.n324 B.n91 10.6151
R861 B.n325 B.n324 10.6151
R862 B.n326 B.n325 10.6151
R863 B.n326 B.n89 10.6151
R864 B.n38 B.n34 9.36635
R865 B.n463 B.n462 9.36635
R866 B.n247 B.n246 9.36635
R867 B.n265 B.n264 9.36635
R868 B.n577 B.n0 8.11757
R869 B.n577 B.n1 8.11757
R870 B.n477 B.n38 1.24928
R871 B.n464 B.n463 1.24928
R872 B.n246 B.n117 1.24928
R873 B.n264 B.n263 1.24928
R874 VP.n0 VP.t0 247.052
R875 VP.n0 VP.t1 203.345
R876 VP VP.n0 0.241678
R877 VTAIL.n1 VTAIL.t0 60.2968
R878 VTAIL.n3 VTAIL.t1 60.2967
R879 VTAIL.n0 VTAIL.t2 60.2967
R880 VTAIL.n2 VTAIL.t3 60.2967
R881 VTAIL.n1 VTAIL.n0 27.341
R882 VTAIL.n3 VTAIL.n2 25.2548
R883 VTAIL.n2 VTAIL.n1 1.51343
R884 VTAIL VTAIL.n0 1.05007
R885 VTAIL VTAIL.n3 0.463862
R886 VDD1 VDD1.t0 116.656
R887 VDD1 VDD1.t1 77.5552
R888 VN VN.t0 247.243
R889 VN VN.t1 203.588
R890 VDD2.n0 VDD2.t0 115.609
R891 VDD2.n0 VDD2.t1 76.9754
R892 VDD2 VDD2.n0 0.580241
C0 VP VTAIL 2.40118f
C1 VTAIL VN 2.38683f
C2 VDD2 VTAIL 5.21335f
C3 B VDD1 1.67701f
C4 w_n1938_n3474# VTAIL 2.851f
C5 B VP 1.37199f
C6 B VN 0.969988f
C7 VP VDD1 2.94791f
C8 VN VDD1 0.147888f
C9 VDD2 B 1.70258f
C10 VDD2 VDD1 0.613973f
C11 B w_n1938_n3474# 8.40723f
C12 w_n1938_n3474# VDD1 1.76142f
C13 VP VN 5.31084f
C14 VDD2 VP 0.311728f
C15 VDD2 VN 2.78702f
C16 B VTAIL 3.55536f
C17 VTAIL VDD1 5.16695f
C18 w_n1938_n3474# VP 2.88088f
C19 w_n1938_n3474# VN 2.63511f
C20 VDD2 w_n1938_n3474# 1.78118f
C21 VDD2 VSUBS 0.863691f
C22 VDD1 VSUBS 4.39374f
C23 VTAIL VSUBS 0.962329f
C24 VN VSUBS 7.79132f
C25 VP VSUBS 1.551677f
C26 B VSUBS 3.557402f
C27 w_n1938_n3474# VSUBS 82.8146f
C28 VDD2.t0 VSUBS 2.59606f
C29 VDD2.t1 VSUBS 2.05207f
C30 VDD2.n0 VSUBS 3.24584f
C31 VN.t1 VSUBS 3.50438f
C32 VN.t0 VSUBS 4.03898f
C33 VDD1.t1 VSUBS 2.06223f
C34 VDD1.t0 VSUBS 2.63558f
C35 VTAIL.t2 VSUBS 2.79522f
C36 VTAIL.n0 VSUBS 2.68434f
C37 VTAIL.t0 VSUBS 2.79524f
C38 VTAIL.n1 VSUBS 2.72793f
C39 VTAIL.t3 VSUBS 2.79522f
C40 VTAIL.n2 VSUBS 2.53162f
C41 VTAIL.t1 VSUBS 2.79522f
C42 VTAIL.n3 VSUBS 2.43285f
C43 VP.t0 VSUBS 4.1762f
C44 VP.t1 VSUBS 3.62698f
C45 VP.n0 VSUBS 5.61772f
C46 B.n0 VSUBS 0.005556f
C47 B.n1 VSUBS 0.005556f
C48 B.n2 VSUBS 0.008218f
C49 B.n3 VSUBS 0.006297f
C50 B.n4 VSUBS 0.006297f
C51 B.n5 VSUBS 0.006297f
C52 B.n6 VSUBS 0.006297f
C53 B.n7 VSUBS 0.006297f
C54 B.n8 VSUBS 0.006297f
C55 B.n9 VSUBS 0.006297f
C56 B.n10 VSUBS 0.006297f
C57 B.n11 VSUBS 0.006297f
C58 B.n12 VSUBS 0.006297f
C59 B.n13 VSUBS 0.014378f
C60 B.n14 VSUBS 0.006297f
C61 B.n15 VSUBS 0.006297f
C62 B.n16 VSUBS 0.006297f
C63 B.n17 VSUBS 0.006297f
C64 B.n18 VSUBS 0.006297f
C65 B.n19 VSUBS 0.006297f
C66 B.n20 VSUBS 0.006297f
C67 B.n21 VSUBS 0.006297f
C68 B.n22 VSUBS 0.006297f
C69 B.n23 VSUBS 0.006297f
C70 B.n24 VSUBS 0.006297f
C71 B.n25 VSUBS 0.006297f
C72 B.n26 VSUBS 0.006297f
C73 B.n27 VSUBS 0.006297f
C74 B.n28 VSUBS 0.006297f
C75 B.n29 VSUBS 0.006297f
C76 B.n30 VSUBS 0.006297f
C77 B.n31 VSUBS 0.006297f
C78 B.n32 VSUBS 0.006297f
C79 B.n33 VSUBS 0.006297f
C80 B.n34 VSUBS 0.005927f
C81 B.n35 VSUBS 0.006297f
C82 B.t1 VSUBS 0.36901f
C83 B.t2 VSUBS 0.384818f
C84 B.t0 VSUBS 1.05364f
C85 B.n36 VSUBS 0.190232f
C86 B.n37 VSUBS 0.062715f
C87 B.n38 VSUBS 0.01459f
C88 B.n39 VSUBS 0.006297f
C89 B.n40 VSUBS 0.006297f
C90 B.n41 VSUBS 0.006297f
C91 B.n42 VSUBS 0.006297f
C92 B.t7 VSUBS 0.369003f
C93 B.t8 VSUBS 0.384812f
C94 B.t6 VSUBS 1.05364f
C95 B.n43 VSUBS 0.190239f
C96 B.n44 VSUBS 0.062722f
C97 B.n45 VSUBS 0.006297f
C98 B.n46 VSUBS 0.006297f
C99 B.n47 VSUBS 0.006297f
C100 B.n48 VSUBS 0.006297f
C101 B.n49 VSUBS 0.006297f
C102 B.n50 VSUBS 0.006297f
C103 B.n51 VSUBS 0.006297f
C104 B.n52 VSUBS 0.006297f
C105 B.n53 VSUBS 0.006297f
C106 B.n54 VSUBS 0.006297f
C107 B.n55 VSUBS 0.006297f
C108 B.n56 VSUBS 0.006297f
C109 B.n57 VSUBS 0.006297f
C110 B.n58 VSUBS 0.006297f
C111 B.n59 VSUBS 0.006297f
C112 B.n60 VSUBS 0.006297f
C113 B.n61 VSUBS 0.006297f
C114 B.n62 VSUBS 0.006297f
C115 B.n63 VSUBS 0.006297f
C116 B.n64 VSUBS 0.006297f
C117 B.n65 VSUBS 0.006297f
C118 B.n66 VSUBS 0.013774f
C119 B.n67 VSUBS 0.006297f
C120 B.n68 VSUBS 0.006297f
C121 B.n69 VSUBS 0.006297f
C122 B.n70 VSUBS 0.006297f
C123 B.n71 VSUBS 0.006297f
C124 B.n72 VSUBS 0.006297f
C125 B.n73 VSUBS 0.006297f
C126 B.n74 VSUBS 0.006297f
C127 B.n75 VSUBS 0.006297f
C128 B.n76 VSUBS 0.006297f
C129 B.n77 VSUBS 0.006297f
C130 B.n78 VSUBS 0.006297f
C131 B.n79 VSUBS 0.006297f
C132 B.n80 VSUBS 0.006297f
C133 B.n81 VSUBS 0.006297f
C134 B.n82 VSUBS 0.006297f
C135 B.n83 VSUBS 0.006297f
C136 B.n84 VSUBS 0.006297f
C137 B.n85 VSUBS 0.006297f
C138 B.n86 VSUBS 0.006297f
C139 B.n87 VSUBS 0.006297f
C140 B.n88 VSUBS 0.006297f
C141 B.n89 VSUBS 0.01358f
C142 B.n90 VSUBS 0.006297f
C143 B.n91 VSUBS 0.006297f
C144 B.n92 VSUBS 0.006297f
C145 B.n93 VSUBS 0.006297f
C146 B.n94 VSUBS 0.006297f
C147 B.n95 VSUBS 0.006297f
C148 B.n96 VSUBS 0.006297f
C149 B.n97 VSUBS 0.006297f
C150 B.n98 VSUBS 0.006297f
C151 B.n99 VSUBS 0.006297f
C152 B.n100 VSUBS 0.006297f
C153 B.n101 VSUBS 0.006297f
C154 B.n102 VSUBS 0.006297f
C155 B.n103 VSUBS 0.006297f
C156 B.n104 VSUBS 0.006297f
C157 B.n105 VSUBS 0.006297f
C158 B.n106 VSUBS 0.006297f
C159 B.n107 VSUBS 0.006297f
C160 B.n108 VSUBS 0.006297f
C161 B.n109 VSUBS 0.006297f
C162 B.n110 VSUBS 0.006297f
C163 B.t11 VSUBS 0.369003f
C164 B.t10 VSUBS 0.384812f
C165 B.t9 VSUBS 1.05364f
C166 B.n111 VSUBS 0.190239f
C167 B.n112 VSUBS 0.062722f
C168 B.n113 VSUBS 0.006297f
C169 B.n114 VSUBS 0.006297f
C170 B.n115 VSUBS 0.006297f
C171 B.n116 VSUBS 0.006297f
C172 B.n117 VSUBS 0.003519f
C173 B.n118 VSUBS 0.006297f
C174 B.n119 VSUBS 0.006297f
C175 B.n120 VSUBS 0.006297f
C176 B.n121 VSUBS 0.006297f
C177 B.n122 VSUBS 0.006297f
C178 B.n123 VSUBS 0.006297f
C179 B.n124 VSUBS 0.006297f
C180 B.n125 VSUBS 0.006297f
C181 B.n126 VSUBS 0.006297f
C182 B.n127 VSUBS 0.006297f
C183 B.n128 VSUBS 0.006297f
C184 B.n129 VSUBS 0.006297f
C185 B.n130 VSUBS 0.006297f
C186 B.n131 VSUBS 0.006297f
C187 B.n132 VSUBS 0.006297f
C188 B.n133 VSUBS 0.006297f
C189 B.n134 VSUBS 0.006297f
C190 B.n135 VSUBS 0.006297f
C191 B.n136 VSUBS 0.006297f
C192 B.n137 VSUBS 0.006297f
C193 B.n138 VSUBS 0.006297f
C194 B.n139 VSUBS 0.013774f
C195 B.n140 VSUBS 0.006297f
C196 B.n141 VSUBS 0.006297f
C197 B.n142 VSUBS 0.006297f
C198 B.n143 VSUBS 0.006297f
C199 B.n144 VSUBS 0.006297f
C200 B.n145 VSUBS 0.006297f
C201 B.n146 VSUBS 0.006297f
C202 B.n147 VSUBS 0.006297f
C203 B.n148 VSUBS 0.006297f
C204 B.n149 VSUBS 0.006297f
C205 B.n150 VSUBS 0.006297f
C206 B.n151 VSUBS 0.006297f
C207 B.n152 VSUBS 0.006297f
C208 B.n153 VSUBS 0.006297f
C209 B.n154 VSUBS 0.006297f
C210 B.n155 VSUBS 0.006297f
C211 B.n156 VSUBS 0.006297f
C212 B.n157 VSUBS 0.006297f
C213 B.n158 VSUBS 0.006297f
C214 B.n159 VSUBS 0.006297f
C215 B.n160 VSUBS 0.006297f
C216 B.n161 VSUBS 0.006297f
C217 B.n162 VSUBS 0.006297f
C218 B.n163 VSUBS 0.006297f
C219 B.n164 VSUBS 0.006297f
C220 B.n165 VSUBS 0.006297f
C221 B.n166 VSUBS 0.006297f
C222 B.n167 VSUBS 0.006297f
C223 B.n168 VSUBS 0.006297f
C224 B.n169 VSUBS 0.006297f
C225 B.n170 VSUBS 0.006297f
C226 B.n171 VSUBS 0.006297f
C227 B.n172 VSUBS 0.006297f
C228 B.n173 VSUBS 0.006297f
C229 B.n174 VSUBS 0.006297f
C230 B.n175 VSUBS 0.006297f
C231 B.n176 VSUBS 0.006297f
C232 B.n177 VSUBS 0.006297f
C233 B.n178 VSUBS 0.006297f
C234 B.n179 VSUBS 0.006297f
C235 B.n180 VSUBS 0.013774f
C236 B.n181 VSUBS 0.014378f
C237 B.n182 VSUBS 0.014378f
C238 B.n183 VSUBS 0.006297f
C239 B.n184 VSUBS 0.006297f
C240 B.n185 VSUBS 0.006297f
C241 B.n186 VSUBS 0.006297f
C242 B.n187 VSUBS 0.006297f
C243 B.n188 VSUBS 0.006297f
C244 B.n189 VSUBS 0.006297f
C245 B.n190 VSUBS 0.006297f
C246 B.n191 VSUBS 0.006297f
C247 B.n192 VSUBS 0.006297f
C248 B.n193 VSUBS 0.006297f
C249 B.n194 VSUBS 0.006297f
C250 B.n195 VSUBS 0.006297f
C251 B.n196 VSUBS 0.006297f
C252 B.n197 VSUBS 0.006297f
C253 B.n198 VSUBS 0.006297f
C254 B.n199 VSUBS 0.006297f
C255 B.n200 VSUBS 0.006297f
C256 B.n201 VSUBS 0.006297f
C257 B.n202 VSUBS 0.006297f
C258 B.n203 VSUBS 0.006297f
C259 B.n204 VSUBS 0.006297f
C260 B.n205 VSUBS 0.006297f
C261 B.n206 VSUBS 0.006297f
C262 B.n207 VSUBS 0.006297f
C263 B.n208 VSUBS 0.006297f
C264 B.n209 VSUBS 0.006297f
C265 B.n210 VSUBS 0.006297f
C266 B.n211 VSUBS 0.006297f
C267 B.n212 VSUBS 0.006297f
C268 B.n213 VSUBS 0.006297f
C269 B.n214 VSUBS 0.006297f
C270 B.n215 VSUBS 0.006297f
C271 B.n216 VSUBS 0.006297f
C272 B.n217 VSUBS 0.006297f
C273 B.n218 VSUBS 0.006297f
C274 B.n219 VSUBS 0.006297f
C275 B.n220 VSUBS 0.006297f
C276 B.n221 VSUBS 0.006297f
C277 B.n222 VSUBS 0.006297f
C278 B.n223 VSUBS 0.006297f
C279 B.n224 VSUBS 0.006297f
C280 B.n225 VSUBS 0.006297f
C281 B.n226 VSUBS 0.006297f
C282 B.n227 VSUBS 0.006297f
C283 B.n228 VSUBS 0.006297f
C284 B.n229 VSUBS 0.006297f
C285 B.n230 VSUBS 0.006297f
C286 B.n231 VSUBS 0.006297f
C287 B.n232 VSUBS 0.006297f
C288 B.n233 VSUBS 0.006297f
C289 B.n234 VSUBS 0.006297f
C290 B.n235 VSUBS 0.006297f
C291 B.n236 VSUBS 0.006297f
C292 B.n237 VSUBS 0.006297f
C293 B.n238 VSUBS 0.006297f
C294 B.n239 VSUBS 0.006297f
C295 B.n240 VSUBS 0.006297f
C296 B.n241 VSUBS 0.006297f
C297 B.n242 VSUBS 0.006297f
C298 B.n243 VSUBS 0.006297f
C299 B.t5 VSUBS 0.36901f
C300 B.t4 VSUBS 0.384818f
C301 B.t3 VSUBS 1.05364f
C302 B.n244 VSUBS 0.190232f
C303 B.n245 VSUBS 0.062715f
C304 B.n246 VSUBS 0.01459f
C305 B.n247 VSUBS 0.005927f
C306 B.n248 VSUBS 0.006297f
C307 B.n249 VSUBS 0.006297f
C308 B.n250 VSUBS 0.006297f
C309 B.n251 VSUBS 0.006297f
C310 B.n252 VSUBS 0.006297f
C311 B.n253 VSUBS 0.006297f
C312 B.n254 VSUBS 0.006297f
C313 B.n255 VSUBS 0.006297f
C314 B.n256 VSUBS 0.006297f
C315 B.n257 VSUBS 0.006297f
C316 B.n258 VSUBS 0.006297f
C317 B.n259 VSUBS 0.006297f
C318 B.n260 VSUBS 0.006297f
C319 B.n261 VSUBS 0.006297f
C320 B.n262 VSUBS 0.006297f
C321 B.n263 VSUBS 0.003519f
C322 B.n264 VSUBS 0.01459f
C323 B.n265 VSUBS 0.005927f
C324 B.n266 VSUBS 0.006297f
C325 B.n267 VSUBS 0.006297f
C326 B.n268 VSUBS 0.006297f
C327 B.n269 VSUBS 0.006297f
C328 B.n270 VSUBS 0.006297f
C329 B.n271 VSUBS 0.006297f
C330 B.n272 VSUBS 0.006297f
C331 B.n273 VSUBS 0.006297f
C332 B.n274 VSUBS 0.006297f
C333 B.n275 VSUBS 0.006297f
C334 B.n276 VSUBS 0.006297f
C335 B.n277 VSUBS 0.006297f
C336 B.n278 VSUBS 0.006297f
C337 B.n279 VSUBS 0.006297f
C338 B.n280 VSUBS 0.006297f
C339 B.n281 VSUBS 0.006297f
C340 B.n282 VSUBS 0.006297f
C341 B.n283 VSUBS 0.006297f
C342 B.n284 VSUBS 0.006297f
C343 B.n285 VSUBS 0.006297f
C344 B.n286 VSUBS 0.006297f
C345 B.n287 VSUBS 0.006297f
C346 B.n288 VSUBS 0.006297f
C347 B.n289 VSUBS 0.006297f
C348 B.n290 VSUBS 0.006297f
C349 B.n291 VSUBS 0.006297f
C350 B.n292 VSUBS 0.006297f
C351 B.n293 VSUBS 0.006297f
C352 B.n294 VSUBS 0.006297f
C353 B.n295 VSUBS 0.006297f
C354 B.n296 VSUBS 0.006297f
C355 B.n297 VSUBS 0.006297f
C356 B.n298 VSUBS 0.006297f
C357 B.n299 VSUBS 0.006297f
C358 B.n300 VSUBS 0.006297f
C359 B.n301 VSUBS 0.006297f
C360 B.n302 VSUBS 0.006297f
C361 B.n303 VSUBS 0.006297f
C362 B.n304 VSUBS 0.006297f
C363 B.n305 VSUBS 0.006297f
C364 B.n306 VSUBS 0.006297f
C365 B.n307 VSUBS 0.006297f
C366 B.n308 VSUBS 0.006297f
C367 B.n309 VSUBS 0.006297f
C368 B.n310 VSUBS 0.006297f
C369 B.n311 VSUBS 0.006297f
C370 B.n312 VSUBS 0.006297f
C371 B.n313 VSUBS 0.006297f
C372 B.n314 VSUBS 0.006297f
C373 B.n315 VSUBS 0.006297f
C374 B.n316 VSUBS 0.006297f
C375 B.n317 VSUBS 0.006297f
C376 B.n318 VSUBS 0.006297f
C377 B.n319 VSUBS 0.006297f
C378 B.n320 VSUBS 0.006297f
C379 B.n321 VSUBS 0.006297f
C380 B.n322 VSUBS 0.006297f
C381 B.n323 VSUBS 0.006297f
C382 B.n324 VSUBS 0.006297f
C383 B.n325 VSUBS 0.006297f
C384 B.n326 VSUBS 0.006297f
C385 B.n327 VSUBS 0.006297f
C386 B.n328 VSUBS 0.014378f
C387 B.n329 VSUBS 0.013774f
C388 B.n330 VSUBS 0.014573f
C389 B.n331 VSUBS 0.006297f
C390 B.n332 VSUBS 0.006297f
C391 B.n333 VSUBS 0.006297f
C392 B.n334 VSUBS 0.006297f
C393 B.n335 VSUBS 0.006297f
C394 B.n336 VSUBS 0.006297f
C395 B.n337 VSUBS 0.006297f
C396 B.n338 VSUBS 0.006297f
C397 B.n339 VSUBS 0.006297f
C398 B.n340 VSUBS 0.006297f
C399 B.n341 VSUBS 0.006297f
C400 B.n342 VSUBS 0.006297f
C401 B.n343 VSUBS 0.006297f
C402 B.n344 VSUBS 0.006297f
C403 B.n345 VSUBS 0.006297f
C404 B.n346 VSUBS 0.006297f
C405 B.n347 VSUBS 0.006297f
C406 B.n348 VSUBS 0.006297f
C407 B.n349 VSUBS 0.006297f
C408 B.n350 VSUBS 0.006297f
C409 B.n351 VSUBS 0.006297f
C410 B.n352 VSUBS 0.006297f
C411 B.n353 VSUBS 0.006297f
C412 B.n354 VSUBS 0.006297f
C413 B.n355 VSUBS 0.006297f
C414 B.n356 VSUBS 0.006297f
C415 B.n357 VSUBS 0.006297f
C416 B.n358 VSUBS 0.006297f
C417 B.n359 VSUBS 0.006297f
C418 B.n360 VSUBS 0.006297f
C419 B.n361 VSUBS 0.006297f
C420 B.n362 VSUBS 0.006297f
C421 B.n363 VSUBS 0.006297f
C422 B.n364 VSUBS 0.006297f
C423 B.n365 VSUBS 0.006297f
C424 B.n366 VSUBS 0.006297f
C425 B.n367 VSUBS 0.006297f
C426 B.n368 VSUBS 0.006297f
C427 B.n369 VSUBS 0.006297f
C428 B.n370 VSUBS 0.006297f
C429 B.n371 VSUBS 0.006297f
C430 B.n372 VSUBS 0.006297f
C431 B.n373 VSUBS 0.006297f
C432 B.n374 VSUBS 0.006297f
C433 B.n375 VSUBS 0.006297f
C434 B.n376 VSUBS 0.006297f
C435 B.n377 VSUBS 0.006297f
C436 B.n378 VSUBS 0.006297f
C437 B.n379 VSUBS 0.006297f
C438 B.n380 VSUBS 0.006297f
C439 B.n381 VSUBS 0.006297f
C440 B.n382 VSUBS 0.006297f
C441 B.n383 VSUBS 0.006297f
C442 B.n384 VSUBS 0.006297f
C443 B.n385 VSUBS 0.006297f
C444 B.n386 VSUBS 0.006297f
C445 B.n387 VSUBS 0.006297f
C446 B.n388 VSUBS 0.006297f
C447 B.n389 VSUBS 0.006297f
C448 B.n390 VSUBS 0.006297f
C449 B.n391 VSUBS 0.006297f
C450 B.n392 VSUBS 0.006297f
C451 B.n393 VSUBS 0.006297f
C452 B.n394 VSUBS 0.006297f
C453 B.n395 VSUBS 0.006297f
C454 B.n396 VSUBS 0.006297f
C455 B.n397 VSUBS 0.013774f
C456 B.n398 VSUBS 0.014378f
C457 B.n399 VSUBS 0.014378f
C458 B.n400 VSUBS 0.006297f
C459 B.n401 VSUBS 0.006297f
C460 B.n402 VSUBS 0.006297f
C461 B.n403 VSUBS 0.006297f
C462 B.n404 VSUBS 0.006297f
C463 B.n405 VSUBS 0.006297f
C464 B.n406 VSUBS 0.006297f
C465 B.n407 VSUBS 0.006297f
C466 B.n408 VSUBS 0.006297f
C467 B.n409 VSUBS 0.006297f
C468 B.n410 VSUBS 0.006297f
C469 B.n411 VSUBS 0.006297f
C470 B.n412 VSUBS 0.006297f
C471 B.n413 VSUBS 0.006297f
C472 B.n414 VSUBS 0.006297f
C473 B.n415 VSUBS 0.006297f
C474 B.n416 VSUBS 0.006297f
C475 B.n417 VSUBS 0.006297f
C476 B.n418 VSUBS 0.006297f
C477 B.n419 VSUBS 0.006297f
C478 B.n420 VSUBS 0.006297f
C479 B.n421 VSUBS 0.006297f
C480 B.n422 VSUBS 0.006297f
C481 B.n423 VSUBS 0.006297f
C482 B.n424 VSUBS 0.006297f
C483 B.n425 VSUBS 0.006297f
C484 B.n426 VSUBS 0.006297f
C485 B.n427 VSUBS 0.006297f
C486 B.n428 VSUBS 0.006297f
C487 B.n429 VSUBS 0.006297f
C488 B.n430 VSUBS 0.006297f
C489 B.n431 VSUBS 0.006297f
C490 B.n432 VSUBS 0.006297f
C491 B.n433 VSUBS 0.006297f
C492 B.n434 VSUBS 0.006297f
C493 B.n435 VSUBS 0.006297f
C494 B.n436 VSUBS 0.006297f
C495 B.n437 VSUBS 0.006297f
C496 B.n438 VSUBS 0.006297f
C497 B.n439 VSUBS 0.006297f
C498 B.n440 VSUBS 0.006297f
C499 B.n441 VSUBS 0.006297f
C500 B.n442 VSUBS 0.006297f
C501 B.n443 VSUBS 0.006297f
C502 B.n444 VSUBS 0.006297f
C503 B.n445 VSUBS 0.006297f
C504 B.n446 VSUBS 0.006297f
C505 B.n447 VSUBS 0.006297f
C506 B.n448 VSUBS 0.006297f
C507 B.n449 VSUBS 0.006297f
C508 B.n450 VSUBS 0.006297f
C509 B.n451 VSUBS 0.006297f
C510 B.n452 VSUBS 0.006297f
C511 B.n453 VSUBS 0.006297f
C512 B.n454 VSUBS 0.006297f
C513 B.n455 VSUBS 0.006297f
C514 B.n456 VSUBS 0.006297f
C515 B.n457 VSUBS 0.006297f
C516 B.n458 VSUBS 0.006297f
C517 B.n459 VSUBS 0.006297f
C518 B.n460 VSUBS 0.006297f
C519 B.n461 VSUBS 0.006297f
C520 B.n462 VSUBS 0.005927f
C521 B.n463 VSUBS 0.01459f
C522 B.n464 VSUBS 0.003519f
C523 B.n465 VSUBS 0.006297f
C524 B.n466 VSUBS 0.006297f
C525 B.n467 VSUBS 0.006297f
C526 B.n468 VSUBS 0.006297f
C527 B.n469 VSUBS 0.006297f
C528 B.n470 VSUBS 0.006297f
C529 B.n471 VSUBS 0.006297f
C530 B.n472 VSUBS 0.006297f
C531 B.n473 VSUBS 0.006297f
C532 B.n474 VSUBS 0.006297f
C533 B.n475 VSUBS 0.006297f
C534 B.n476 VSUBS 0.006297f
C535 B.n477 VSUBS 0.003519f
C536 B.n478 VSUBS 0.006297f
C537 B.n479 VSUBS 0.006297f
C538 B.n480 VSUBS 0.006297f
C539 B.n481 VSUBS 0.006297f
C540 B.n482 VSUBS 0.006297f
C541 B.n483 VSUBS 0.006297f
C542 B.n484 VSUBS 0.006297f
C543 B.n485 VSUBS 0.006297f
C544 B.n486 VSUBS 0.006297f
C545 B.n487 VSUBS 0.006297f
C546 B.n488 VSUBS 0.006297f
C547 B.n489 VSUBS 0.006297f
C548 B.n490 VSUBS 0.006297f
C549 B.n491 VSUBS 0.006297f
C550 B.n492 VSUBS 0.006297f
C551 B.n493 VSUBS 0.006297f
C552 B.n494 VSUBS 0.006297f
C553 B.n495 VSUBS 0.006297f
C554 B.n496 VSUBS 0.006297f
C555 B.n497 VSUBS 0.006297f
C556 B.n498 VSUBS 0.006297f
C557 B.n499 VSUBS 0.006297f
C558 B.n500 VSUBS 0.006297f
C559 B.n501 VSUBS 0.006297f
C560 B.n502 VSUBS 0.006297f
C561 B.n503 VSUBS 0.006297f
C562 B.n504 VSUBS 0.006297f
C563 B.n505 VSUBS 0.006297f
C564 B.n506 VSUBS 0.006297f
C565 B.n507 VSUBS 0.006297f
C566 B.n508 VSUBS 0.006297f
C567 B.n509 VSUBS 0.006297f
C568 B.n510 VSUBS 0.006297f
C569 B.n511 VSUBS 0.006297f
C570 B.n512 VSUBS 0.006297f
C571 B.n513 VSUBS 0.006297f
C572 B.n514 VSUBS 0.006297f
C573 B.n515 VSUBS 0.006297f
C574 B.n516 VSUBS 0.006297f
C575 B.n517 VSUBS 0.006297f
C576 B.n518 VSUBS 0.006297f
C577 B.n519 VSUBS 0.006297f
C578 B.n520 VSUBS 0.006297f
C579 B.n521 VSUBS 0.006297f
C580 B.n522 VSUBS 0.006297f
C581 B.n523 VSUBS 0.006297f
C582 B.n524 VSUBS 0.006297f
C583 B.n525 VSUBS 0.006297f
C584 B.n526 VSUBS 0.006297f
C585 B.n527 VSUBS 0.006297f
C586 B.n528 VSUBS 0.006297f
C587 B.n529 VSUBS 0.006297f
C588 B.n530 VSUBS 0.006297f
C589 B.n531 VSUBS 0.006297f
C590 B.n532 VSUBS 0.006297f
C591 B.n533 VSUBS 0.006297f
C592 B.n534 VSUBS 0.006297f
C593 B.n535 VSUBS 0.006297f
C594 B.n536 VSUBS 0.006297f
C595 B.n537 VSUBS 0.006297f
C596 B.n538 VSUBS 0.006297f
C597 B.n539 VSUBS 0.006297f
C598 B.n540 VSUBS 0.006297f
C599 B.n541 VSUBS 0.006297f
C600 B.n542 VSUBS 0.014378f
C601 B.n543 VSUBS 0.013774f
C602 B.n544 VSUBS 0.013774f
C603 B.n545 VSUBS 0.006297f
C604 B.n546 VSUBS 0.006297f
C605 B.n547 VSUBS 0.006297f
C606 B.n548 VSUBS 0.006297f
C607 B.n549 VSUBS 0.006297f
C608 B.n550 VSUBS 0.006297f
C609 B.n551 VSUBS 0.006297f
C610 B.n552 VSUBS 0.006297f
C611 B.n553 VSUBS 0.006297f
C612 B.n554 VSUBS 0.006297f
C613 B.n555 VSUBS 0.006297f
C614 B.n556 VSUBS 0.006297f
C615 B.n557 VSUBS 0.006297f
C616 B.n558 VSUBS 0.006297f
C617 B.n559 VSUBS 0.006297f
C618 B.n560 VSUBS 0.006297f
C619 B.n561 VSUBS 0.006297f
C620 B.n562 VSUBS 0.006297f
C621 B.n563 VSUBS 0.006297f
C622 B.n564 VSUBS 0.006297f
C623 B.n565 VSUBS 0.006297f
C624 B.n566 VSUBS 0.006297f
C625 B.n567 VSUBS 0.006297f
C626 B.n568 VSUBS 0.006297f
C627 B.n569 VSUBS 0.006297f
C628 B.n570 VSUBS 0.006297f
C629 B.n571 VSUBS 0.006297f
C630 B.n572 VSUBS 0.006297f
C631 B.n573 VSUBS 0.006297f
C632 B.n574 VSUBS 0.006297f
C633 B.n575 VSUBS 0.008218f
C634 B.n576 VSUBS 0.008754f
C635 B.n577 VSUBS 0.017408f
.ends

