* NGSPICE file created from diff_pair_sample_0530.ext - technology: sky130A

.subckt diff_pair_sample_0530 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t2 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=3.2802 pd=20.21 as=7.7532 ps=40.54 w=19.88 l=2.12
X1 VDD1.t2 VP.t1 VTAIL.t5 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=3.2802 pd=20.21 as=7.7532 ps=40.54 w=19.88 l=2.12
X2 VDD2.t3 VN.t0 VTAIL.t6 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=3.2802 pd=20.21 as=7.7532 ps=40.54 w=19.88 l=2.12
X3 VTAIL.t0 VN.t1 VDD2.t2 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=3.2802 ps=20.21 w=19.88 l=2.12
X4 B.t11 B.t9 B.t10 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=0 ps=0 w=19.88 l=2.12
X5 VTAIL.t4 VP.t2 VDD1.t1 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=3.2802 ps=20.21 w=19.88 l=2.12
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=3.2802 ps=20.21 w=19.88 l=2.12
X7 VDD2.t0 VN.t3 VTAIL.t7 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=3.2802 pd=20.21 as=7.7532 ps=40.54 w=19.88 l=2.12
X8 B.t8 B.t6 B.t7 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=0 ps=0 w=19.88 l=2.12
X9 B.t5 B.t3 B.t4 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=0 ps=0 w=19.88 l=2.12
X10 B.t2 B.t0 B.t1 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=0 ps=0 w=19.88 l=2.12
X11 VTAIL.t3 VP.t3 VDD1.t0 w_n2440_n4944# sky130_fd_pr__pfet_01v8 ad=7.7532 pd=40.54 as=3.2802 ps=20.21 w=19.88 l=2.12
R0 VP.n2 VP.t2 262.272
R1 VP.n2 VP.t0 261.719
R2 VP.n4 VP.t3 225.994
R3 VP.n11 VP.t1 225.994
R4 VP.n10 VP.n0 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n1 161.3
R7 VP.n6 VP.n5 161.3
R8 VP.n4 VP.n3 87.546
R9 VP.n12 VP.n11 87.546
R10 VP.n3 VP.n2 57.6747
R11 VP.n9 VP.n1 56.5617
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 23.3627
R15 VP.n11 VP.n10 23.3627
R16 VP.n6 VP.n3 0.278335
R17 VP.n12 VP.n0 0.278335
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153485
R22 VTAIL.n5 VTAIL.t4 56.5573
R23 VTAIL.n4 VTAIL.t7 56.5573
R24 VTAIL.n3 VTAIL.t0 56.5573
R25 VTAIL.n7 VTAIL.t6 56.5571
R26 VTAIL.n0 VTAIL.t1 56.5571
R27 VTAIL.n1 VTAIL.t5 56.5571
R28 VTAIL.n2 VTAIL.t3 56.5571
R29 VTAIL.n6 VTAIL.t2 56.5571
R30 VTAIL.n7 VTAIL.n6 31.6169
R31 VTAIL.n3 VTAIL.n2 31.6169
R32 VTAIL.n4 VTAIL.n3 2.11257
R33 VTAIL.n6 VTAIL.n5 2.11257
R34 VTAIL.n2 VTAIL.n1 2.11257
R35 VTAIL VTAIL.n0 1.11472
R36 VTAIL VTAIL.n7 0.998345
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 119.314
R40 VDD1 VDD1.n0 71.659
R41 VDD1.n0 VDD1.t1 1.63556
R42 VDD1.n0 VDD1.t3 1.63556
R43 VDD1.n1 VDD1.t0 1.63556
R44 VDD1.n1 VDD1.t2 1.63556
R45 VN.n0 VN.t2 262.272
R46 VN.n1 VN.t3 262.272
R47 VN.n0 VN.t0 261.719
R48 VN.n1 VN.t1 261.719
R49 VN VN.n1 57.9536
R50 VN VN.n0 6.81341
R51 VDD2.n2 VDD2.n0 118.79
R52 VDD2.n2 VDD2.n1 71.6008
R53 VDD2.n1 VDD2.t2 1.63556
R54 VDD2.n1 VDD2.t0 1.63556
R55 VDD2.n0 VDD2.t1 1.63556
R56 VDD2.n0 VDD2.t3 1.63556
R57 VDD2 VDD2.n2 0.0586897
R58 B.n459 B.n120 585
R59 B.n458 B.n457 585
R60 B.n456 B.n121 585
R61 B.n455 B.n454 585
R62 B.n453 B.n122 585
R63 B.n452 B.n451 585
R64 B.n450 B.n123 585
R65 B.n449 B.n448 585
R66 B.n447 B.n124 585
R67 B.n446 B.n445 585
R68 B.n444 B.n125 585
R69 B.n443 B.n442 585
R70 B.n441 B.n126 585
R71 B.n440 B.n439 585
R72 B.n438 B.n127 585
R73 B.n437 B.n436 585
R74 B.n435 B.n128 585
R75 B.n434 B.n433 585
R76 B.n432 B.n129 585
R77 B.n431 B.n430 585
R78 B.n429 B.n130 585
R79 B.n428 B.n427 585
R80 B.n426 B.n131 585
R81 B.n425 B.n424 585
R82 B.n423 B.n132 585
R83 B.n422 B.n421 585
R84 B.n420 B.n133 585
R85 B.n419 B.n418 585
R86 B.n417 B.n134 585
R87 B.n416 B.n415 585
R88 B.n414 B.n135 585
R89 B.n413 B.n412 585
R90 B.n411 B.n136 585
R91 B.n410 B.n409 585
R92 B.n408 B.n137 585
R93 B.n407 B.n406 585
R94 B.n405 B.n138 585
R95 B.n404 B.n403 585
R96 B.n402 B.n139 585
R97 B.n401 B.n400 585
R98 B.n399 B.n140 585
R99 B.n398 B.n397 585
R100 B.n396 B.n141 585
R101 B.n395 B.n394 585
R102 B.n393 B.n142 585
R103 B.n392 B.n391 585
R104 B.n390 B.n143 585
R105 B.n389 B.n388 585
R106 B.n387 B.n144 585
R107 B.n386 B.n385 585
R108 B.n384 B.n145 585
R109 B.n383 B.n382 585
R110 B.n381 B.n146 585
R111 B.n380 B.n379 585
R112 B.n378 B.n147 585
R113 B.n377 B.n376 585
R114 B.n375 B.n148 585
R115 B.n374 B.n373 585
R116 B.n372 B.n149 585
R117 B.n371 B.n370 585
R118 B.n369 B.n150 585
R119 B.n368 B.n367 585
R120 B.n366 B.n151 585
R121 B.n365 B.n364 585
R122 B.n363 B.n152 585
R123 B.n362 B.n361 585
R124 B.n357 B.n153 585
R125 B.n356 B.n355 585
R126 B.n354 B.n154 585
R127 B.n353 B.n352 585
R128 B.n351 B.n155 585
R129 B.n350 B.n349 585
R130 B.n348 B.n156 585
R131 B.n347 B.n346 585
R132 B.n344 B.n157 585
R133 B.n343 B.n342 585
R134 B.n341 B.n160 585
R135 B.n340 B.n339 585
R136 B.n338 B.n161 585
R137 B.n337 B.n336 585
R138 B.n335 B.n162 585
R139 B.n334 B.n333 585
R140 B.n332 B.n163 585
R141 B.n331 B.n330 585
R142 B.n329 B.n164 585
R143 B.n328 B.n327 585
R144 B.n326 B.n165 585
R145 B.n325 B.n324 585
R146 B.n323 B.n166 585
R147 B.n322 B.n321 585
R148 B.n320 B.n167 585
R149 B.n319 B.n318 585
R150 B.n317 B.n168 585
R151 B.n316 B.n315 585
R152 B.n314 B.n169 585
R153 B.n313 B.n312 585
R154 B.n311 B.n170 585
R155 B.n310 B.n309 585
R156 B.n308 B.n171 585
R157 B.n307 B.n306 585
R158 B.n305 B.n172 585
R159 B.n304 B.n303 585
R160 B.n302 B.n173 585
R161 B.n301 B.n300 585
R162 B.n299 B.n174 585
R163 B.n298 B.n297 585
R164 B.n296 B.n175 585
R165 B.n295 B.n294 585
R166 B.n293 B.n176 585
R167 B.n292 B.n291 585
R168 B.n290 B.n177 585
R169 B.n289 B.n288 585
R170 B.n287 B.n178 585
R171 B.n286 B.n285 585
R172 B.n284 B.n179 585
R173 B.n283 B.n282 585
R174 B.n281 B.n180 585
R175 B.n280 B.n279 585
R176 B.n278 B.n181 585
R177 B.n277 B.n276 585
R178 B.n275 B.n182 585
R179 B.n274 B.n273 585
R180 B.n272 B.n183 585
R181 B.n271 B.n270 585
R182 B.n269 B.n184 585
R183 B.n268 B.n267 585
R184 B.n266 B.n185 585
R185 B.n265 B.n264 585
R186 B.n263 B.n186 585
R187 B.n262 B.n261 585
R188 B.n260 B.n187 585
R189 B.n259 B.n258 585
R190 B.n257 B.n188 585
R191 B.n256 B.n255 585
R192 B.n254 B.n189 585
R193 B.n253 B.n252 585
R194 B.n251 B.n190 585
R195 B.n250 B.n249 585
R196 B.n248 B.n191 585
R197 B.n461 B.n460 585
R198 B.n462 B.n119 585
R199 B.n464 B.n463 585
R200 B.n465 B.n118 585
R201 B.n467 B.n466 585
R202 B.n468 B.n117 585
R203 B.n470 B.n469 585
R204 B.n471 B.n116 585
R205 B.n473 B.n472 585
R206 B.n474 B.n115 585
R207 B.n476 B.n475 585
R208 B.n477 B.n114 585
R209 B.n479 B.n478 585
R210 B.n480 B.n113 585
R211 B.n482 B.n481 585
R212 B.n483 B.n112 585
R213 B.n485 B.n484 585
R214 B.n486 B.n111 585
R215 B.n488 B.n487 585
R216 B.n489 B.n110 585
R217 B.n491 B.n490 585
R218 B.n492 B.n109 585
R219 B.n494 B.n493 585
R220 B.n495 B.n108 585
R221 B.n497 B.n496 585
R222 B.n498 B.n107 585
R223 B.n500 B.n499 585
R224 B.n501 B.n106 585
R225 B.n503 B.n502 585
R226 B.n504 B.n105 585
R227 B.n506 B.n505 585
R228 B.n507 B.n104 585
R229 B.n509 B.n508 585
R230 B.n510 B.n103 585
R231 B.n512 B.n511 585
R232 B.n513 B.n102 585
R233 B.n515 B.n514 585
R234 B.n516 B.n101 585
R235 B.n518 B.n517 585
R236 B.n519 B.n100 585
R237 B.n521 B.n520 585
R238 B.n522 B.n99 585
R239 B.n524 B.n523 585
R240 B.n525 B.n98 585
R241 B.n527 B.n526 585
R242 B.n528 B.n97 585
R243 B.n530 B.n529 585
R244 B.n531 B.n96 585
R245 B.n533 B.n532 585
R246 B.n534 B.n95 585
R247 B.n536 B.n535 585
R248 B.n537 B.n94 585
R249 B.n539 B.n538 585
R250 B.n540 B.n93 585
R251 B.n542 B.n541 585
R252 B.n543 B.n92 585
R253 B.n545 B.n544 585
R254 B.n546 B.n91 585
R255 B.n548 B.n547 585
R256 B.n549 B.n90 585
R257 B.n760 B.n759 585
R258 B.n758 B.n17 585
R259 B.n757 B.n756 585
R260 B.n755 B.n18 585
R261 B.n754 B.n753 585
R262 B.n752 B.n19 585
R263 B.n751 B.n750 585
R264 B.n749 B.n20 585
R265 B.n748 B.n747 585
R266 B.n746 B.n21 585
R267 B.n745 B.n744 585
R268 B.n743 B.n22 585
R269 B.n742 B.n741 585
R270 B.n740 B.n23 585
R271 B.n739 B.n738 585
R272 B.n737 B.n24 585
R273 B.n736 B.n735 585
R274 B.n734 B.n25 585
R275 B.n733 B.n732 585
R276 B.n731 B.n26 585
R277 B.n730 B.n729 585
R278 B.n728 B.n27 585
R279 B.n727 B.n726 585
R280 B.n725 B.n28 585
R281 B.n724 B.n723 585
R282 B.n722 B.n29 585
R283 B.n721 B.n720 585
R284 B.n719 B.n30 585
R285 B.n718 B.n717 585
R286 B.n716 B.n31 585
R287 B.n715 B.n714 585
R288 B.n713 B.n32 585
R289 B.n712 B.n711 585
R290 B.n710 B.n33 585
R291 B.n709 B.n708 585
R292 B.n707 B.n34 585
R293 B.n706 B.n705 585
R294 B.n704 B.n35 585
R295 B.n703 B.n702 585
R296 B.n701 B.n36 585
R297 B.n700 B.n699 585
R298 B.n698 B.n37 585
R299 B.n697 B.n696 585
R300 B.n695 B.n38 585
R301 B.n694 B.n693 585
R302 B.n692 B.n39 585
R303 B.n691 B.n690 585
R304 B.n689 B.n40 585
R305 B.n688 B.n687 585
R306 B.n686 B.n41 585
R307 B.n685 B.n684 585
R308 B.n683 B.n42 585
R309 B.n682 B.n681 585
R310 B.n680 B.n43 585
R311 B.n679 B.n678 585
R312 B.n677 B.n44 585
R313 B.n676 B.n675 585
R314 B.n674 B.n45 585
R315 B.n673 B.n672 585
R316 B.n671 B.n46 585
R317 B.n670 B.n669 585
R318 B.n668 B.n47 585
R319 B.n667 B.n666 585
R320 B.n665 B.n48 585
R321 B.n664 B.n663 585
R322 B.n661 B.n49 585
R323 B.n660 B.n659 585
R324 B.n658 B.n52 585
R325 B.n657 B.n656 585
R326 B.n655 B.n53 585
R327 B.n654 B.n653 585
R328 B.n652 B.n54 585
R329 B.n651 B.n650 585
R330 B.n649 B.n55 585
R331 B.n647 B.n646 585
R332 B.n645 B.n58 585
R333 B.n644 B.n643 585
R334 B.n642 B.n59 585
R335 B.n641 B.n640 585
R336 B.n639 B.n60 585
R337 B.n638 B.n637 585
R338 B.n636 B.n61 585
R339 B.n635 B.n634 585
R340 B.n633 B.n62 585
R341 B.n632 B.n631 585
R342 B.n630 B.n63 585
R343 B.n629 B.n628 585
R344 B.n627 B.n64 585
R345 B.n626 B.n625 585
R346 B.n624 B.n65 585
R347 B.n623 B.n622 585
R348 B.n621 B.n66 585
R349 B.n620 B.n619 585
R350 B.n618 B.n67 585
R351 B.n617 B.n616 585
R352 B.n615 B.n68 585
R353 B.n614 B.n613 585
R354 B.n612 B.n69 585
R355 B.n611 B.n610 585
R356 B.n609 B.n70 585
R357 B.n608 B.n607 585
R358 B.n606 B.n71 585
R359 B.n605 B.n604 585
R360 B.n603 B.n72 585
R361 B.n602 B.n601 585
R362 B.n600 B.n73 585
R363 B.n599 B.n598 585
R364 B.n597 B.n74 585
R365 B.n596 B.n595 585
R366 B.n594 B.n75 585
R367 B.n593 B.n592 585
R368 B.n591 B.n76 585
R369 B.n590 B.n589 585
R370 B.n588 B.n77 585
R371 B.n587 B.n586 585
R372 B.n585 B.n78 585
R373 B.n584 B.n583 585
R374 B.n582 B.n79 585
R375 B.n581 B.n580 585
R376 B.n579 B.n80 585
R377 B.n578 B.n577 585
R378 B.n576 B.n81 585
R379 B.n575 B.n574 585
R380 B.n573 B.n82 585
R381 B.n572 B.n571 585
R382 B.n570 B.n83 585
R383 B.n569 B.n568 585
R384 B.n567 B.n84 585
R385 B.n566 B.n565 585
R386 B.n564 B.n85 585
R387 B.n563 B.n562 585
R388 B.n561 B.n86 585
R389 B.n560 B.n559 585
R390 B.n558 B.n87 585
R391 B.n557 B.n556 585
R392 B.n555 B.n88 585
R393 B.n554 B.n553 585
R394 B.n552 B.n89 585
R395 B.n551 B.n550 585
R396 B.n761 B.n16 585
R397 B.n763 B.n762 585
R398 B.n764 B.n15 585
R399 B.n766 B.n765 585
R400 B.n767 B.n14 585
R401 B.n769 B.n768 585
R402 B.n770 B.n13 585
R403 B.n772 B.n771 585
R404 B.n773 B.n12 585
R405 B.n775 B.n774 585
R406 B.n776 B.n11 585
R407 B.n778 B.n777 585
R408 B.n779 B.n10 585
R409 B.n781 B.n780 585
R410 B.n782 B.n9 585
R411 B.n784 B.n783 585
R412 B.n785 B.n8 585
R413 B.n787 B.n786 585
R414 B.n788 B.n7 585
R415 B.n790 B.n789 585
R416 B.n791 B.n6 585
R417 B.n793 B.n792 585
R418 B.n794 B.n5 585
R419 B.n796 B.n795 585
R420 B.n797 B.n4 585
R421 B.n799 B.n798 585
R422 B.n800 B.n3 585
R423 B.n802 B.n801 585
R424 B.n803 B.n0 585
R425 B.n2 B.n1 585
R426 B.n206 B.n205 585
R427 B.n208 B.n207 585
R428 B.n209 B.n204 585
R429 B.n211 B.n210 585
R430 B.n212 B.n203 585
R431 B.n214 B.n213 585
R432 B.n215 B.n202 585
R433 B.n217 B.n216 585
R434 B.n218 B.n201 585
R435 B.n220 B.n219 585
R436 B.n221 B.n200 585
R437 B.n223 B.n222 585
R438 B.n224 B.n199 585
R439 B.n226 B.n225 585
R440 B.n227 B.n198 585
R441 B.n229 B.n228 585
R442 B.n230 B.n197 585
R443 B.n232 B.n231 585
R444 B.n233 B.n196 585
R445 B.n235 B.n234 585
R446 B.n236 B.n195 585
R447 B.n238 B.n237 585
R448 B.n239 B.n194 585
R449 B.n241 B.n240 585
R450 B.n242 B.n193 585
R451 B.n244 B.n243 585
R452 B.n245 B.n192 585
R453 B.n247 B.n246 585
R454 B.n246 B.n191 550.159
R455 B.n460 B.n459 550.159
R456 B.n550 B.n549 550.159
R457 B.n761 B.n760 550.159
R458 B.n158 B.t9 433.18
R459 B.n358 B.t0 433.18
R460 B.n56 B.t6 433.18
R461 B.n50 B.t3 433.18
R462 B.n805 B.n804 256.663
R463 B.n804 B.n803 235.042
R464 B.n804 B.n2 235.042
R465 B.n250 B.n191 163.367
R466 B.n251 B.n250 163.367
R467 B.n252 B.n251 163.367
R468 B.n252 B.n189 163.367
R469 B.n256 B.n189 163.367
R470 B.n257 B.n256 163.367
R471 B.n258 B.n257 163.367
R472 B.n258 B.n187 163.367
R473 B.n262 B.n187 163.367
R474 B.n263 B.n262 163.367
R475 B.n264 B.n263 163.367
R476 B.n264 B.n185 163.367
R477 B.n268 B.n185 163.367
R478 B.n269 B.n268 163.367
R479 B.n270 B.n269 163.367
R480 B.n270 B.n183 163.367
R481 B.n274 B.n183 163.367
R482 B.n275 B.n274 163.367
R483 B.n276 B.n275 163.367
R484 B.n276 B.n181 163.367
R485 B.n280 B.n181 163.367
R486 B.n281 B.n280 163.367
R487 B.n282 B.n281 163.367
R488 B.n282 B.n179 163.367
R489 B.n286 B.n179 163.367
R490 B.n287 B.n286 163.367
R491 B.n288 B.n287 163.367
R492 B.n288 B.n177 163.367
R493 B.n292 B.n177 163.367
R494 B.n293 B.n292 163.367
R495 B.n294 B.n293 163.367
R496 B.n294 B.n175 163.367
R497 B.n298 B.n175 163.367
R498 B.n299 B.n298 163.367
R499 B.n300 B.n299 163.367
R500 B.n300 B.n173 163.367
R501 B.n304 B.n173 163.367
R502 B.n305 B.n304 163.367
R503 B.n306 B.n305 163.367
R504 B.n306 B.n171 163.367
R505 B.n310 B.n171 163.367
R506 B.n311 B.n310 163.367
R507 B.n312 B.n311 163.367
R508 B.n312 B.n169 163.367
R509 B.n316 B.n169 163.367
R510 B.n317 B.n316 163.367
R511 B.n318 B.n317 163.367
R512 B.n318 B.n167 163.367
R513 B.n322 B.n167 163.367
R514 B.n323 B.n322 163.367
R515 B.n324 B.n323 163.367
R516 B.n324 B.n165 163.367
R517 B.n328 B.n165 163.367
R518 B.n329 B.n328 163.367
R519 B.n330 B.n329 163.367
R520 B.n330 B.n163 163.367
R521 B.n334 B.n163 163.367
R522 B.n335 B.n334 163.367
R523 B.n336 B.n335 163.367
R524 B.n336 B.n161 163.367
R525 B.n340 B.n161 163.367
R526 B.n341 B.n340 163.367
R527 B.n342 B.n341 163.367
R528 B.n342 B.n157 163.367
R529 B.n347 B.n157 163.367
R530 B.n348 B.n347 163.367
R531 B.n349 B.n348 163.367
R532 B.n349 B.n155 163.367
R533 B.n353 B.n155 163.367
R534 B.n354 B.n353 163.367
R535 B.n355 B.n354 163.367
R536 B.n355 B.n153 163.367
R537 B.n362 B.n153 163.367
R538 B.n363 B.n362 163.367
R539 B.n364 B.n363 163.367
R540 B.n364 B.n151 163.367
R541 B.n368 B.n151 163.367
R542 B.n369 B.n368 163.367
R543 B.n370 B.n369 163.367
R544 B.n370 B.n149 163.367
R545 B.n374 B.n149 163.367
R546 B.n375 B.n374 163.367
R547 B.n376 B.n375 163.367
R548 B.n376 B.n147 163.367
R549 B.n380 B.n147 163.367
R550 B.n381 B.n380 163.367
R551 B.n382 B.n381 163.367
R552 B.n382 B.n145 163.367
R553 B.n386 B.n145 163.367
R554 B.n387 B.n386 163.367
R555 B.n388 B.n387 163.367
R556 B.n388 B.n143 163.367
R557 B.n392 B.n143 163.367
R558 B.n393 B.n392 163.367
R559 B.n394 B.n393 163.367
R560 B.n394 B.n141 163.367
R561 B.n398 B.n141 163.367
R562 B.n399 B.n398 163.367
R563 B.n400 B.n399 163.367
R564 B.n400 B.n139 163.367
R565 B.n404 B.n139 163.367
R566 B.n405 B.n404 163.367
R567 B.n406 B.n405 163.367
R568 B.n406 B.n137 163.367
R569 B.n410 B.n137 163.367
R570 B.n411 B.n410 163.367
R571 B.n412 B.n411 163.367
R572 B.n412 B.n135 163.367
R573 B.n416 B.n135 163.367
R574 B.n417 B.n416 163.367
R575 B.n418 B.n417 163.367
R576 B.n418 B.n133 163.367
R577 B.n422 B.n133 163.367
R578 B.n423 B.n422 163.367
R579 B.n424 B.n423 163.367
R580 B.n424 B.n131 163.367
R581 B.n428 B.n131 163.367
R582 B.n429 B.n428 163.367
R583 B.n430 B.n429 163.367
R584 B.n430 B.n129 163.367
R585 B.n434 B.n129 163.367
R586 B.n435 B.n434 163.367
R587 B.n436 B.n435 163.367
R588 B.n436 B.n127 163.367
R589 B.n440 B.n127 163.367
R590 B.n441 B.n440 163.367
R591 B.n442 B.n441 163.367
R592 B.n442 B.n125 163.367
R593 B.n446 B.n125 163.367
R594 B.n447 B.n446 163.367
R595 B.n448 B.n447 163.367
R596 B.n448 B.n123 163.367
R597 B.n452 B.n123 163.367
R598 B.n453 B.n452 163.367
R599 B.n454 B.n453 163.367
R600 B.n454 B.n121 163.367
R601 B.n458 B.n121 163.367
R602 B.n459 B.n458 163.367
R603 B.n549 B.n548 163.367
R604 B.n548 B.n91 163.367
R605 B.n544 B.n91 163.367
R606 B.n544 B.n543 163.367
R607 B.n543 B.n542 163.367
R608 B.n542 B.n93 163.367
R609 B.n538 B.n93 163.367
R610 B.n538 B.n537 163.367
R611 B.n537 B.n536 163.367
R612 B.n536 B.n95 163.367
R613 B.n532 B.n95 163.367
R614 B.n532 B.n531 163.367
R615 B.n531 B.n530 163.367
R616 B.n530 B.n97 163.367
R617 B.n526 B.n97 163.367
R618 B.n526 B.n525 163.367
R619 B.n525 B.n524 163.367
R620 B.n524 B.n99 163.367
R621 B.n520 B.n99 163.367
R622 B.n520 B.n519 163.367
R623 B.n519 B.n518 163.367
R624 B.n518 B.n101 163.367
R625 B.n514 B.n101 163.367
R626 B.n514 B.n513 163.367
R627 B.n513 B.n512 163.367
R628 B.n512 B.n103 163.367
R629 B.n508 B.n103 163.367
R630 B.n508 B.n507 163.367
R631 B.n507 B.n506 163.367
R632 B.n506 B.n105 163.367
R633 B.n502 B.n105 163.367
R634 B.n502 B.n501 163.367
R635 B.n501 B.n500 163.367
R636 B.n500 B.n107 163.367
R637 B.n496 B.n107 163.367
R638 B.n496 B.n495 163.367
R639 B.n495 B.n494 163.367
R640 B.n494 B.n109 163.367
R641 B.n490 B.n109 163.367
R642 B.n490 B.n489 163.367
R643 B.n489 B.n488 163.367
R644 B.n488 B.n111 163.367
R645 B.n484 B.n111 163.367
R646 B.n484 B.n483 163.367
R647 B.n483 B.n482 163.367
R648 B.n482 B.n113 163.367
R649 B.n478 B.n113 163.367
R650 B.n478 B.n477 163.367
R651 B.n477 B.n476 163.367
R652 B.n476 B.n115 163.367
R653 B.n472 B.n115 163.367
R654 B.n472 B.n471 163.367
R655 B.n471 B.n470 163.367
R656 B.n470 B.n117 163.367
R657 B.n466 B.n117 163.367
R658 B.n466 B.n465 163.367
R659 B.n465 B.n464 163.367
R660 B.n464 B.n119 163.367
R661 B.n460 B.n119 163.367
R662 B.n760 B.n17 163.367
R663 B.n756 B.n17 163.367
R664 B.n756 B.n755 163.367
R665 B.n755 B.n754 163.367
R666 B.n754 B.n19 163.367
R667 B.n750 B.n19 163.367
R668 B.n750 B.n749 163.367
R669 B.n749 B.n748 163.367
R670 B.n748 B.n21 163.367
R671 B.n744 B.n21 163.367
R672 B.n744 B.n743 163.367
R673 B.n743 B.n742 163.367
R674 B.n742 B.n23 163.367
R675 B.n738 B.n23 163.367
R676 B.n738 B.n737 163.367
R677 B.n737 B.n736 163.367
R678 B.n736 B.n25 163.367
R679 B.n732 B.n25 163.367
R680 B.n732 B.n731 163.367
R681 B.n731 B.n730 163.367
R682 B.n730 B.n27 163.367
R683 B.n726 B.n27 163.367
R684 B.n726 B.n725 163.367
R685 B.n725 B.n724 163.367
R686 B.n724 B.n29 163.367
R687 B.n720 B.n29 163.367
R688 B.n720 B.n719 163.367
R689 B.n719 B.n718 163.367
R690 B.n718 B.n31 163.367
R691 B.n714 B.n31 163.367
R692 B.n714 B.n713 163.367
R693 B.n713 B.n712 163.367
R694 B.n712 B.n33 163.367
R695 B.n708 B.n33 163.367
R696 B.n708 B.n707 163.367
R697 B.n707 B.n706 163.367
R698 B.n706 B.n35 163.367
R699 B.n702 B.n35 163.367
R700 B.n702 B.n701 163.367
R701 B.n701 B.n700 163.367
R702 B.n700 B.n37 163.367
R703 B.n696 B.n37 163.367
R704 B.n696 B.n695 163.367
R705 B.n695 B.n694 163.367
R706 B.n694 B.n39 163.367
R707 B.n690 B.n39 163.367
R708 B.n690 B.n689 163.367
R709 B.n689 B.n688 163.367
R710 B.n688 B.n41 163.367
R711 B.n684 B.n41 163.367
R712 B.n684 B.n683 163.367
R713 B.n683 B.n682 163.367
R714 B.n682 B.n43 163.367
R715 B.n678 B.n43 163.367
R716 B.n678 B.n677 163.367
R717 B.n677 B.n676 163.367
R718 B.n676 B.n45 163.367
R719 B.n672 B.n45 163.367
R720 B.n672 B.n671 163.367
R721 B.n671 B.n670 163.367
R722 B.n670 B.n47 163.367
R723 B.n666 B.n47 163.367
R724 B.n666 B.n665 163.367
R725 B.n665 B.n664 163.367
R726 B.n664 B.n49 163.367
R727 B.n659 B.n49 163.367
R728 B.n659 B.n658 163.367
R729 B.n658 B.n657 163.367
R730 B.n657 B.n53 163.367
R731 B.n653 B.n53 163.367
R732 B.n653 B.n652 163.367
R733 B.n652 B.n651 163.367
R734 B.n651 B.n55 163.367
R735 B.n646 B.n55 163.367
R736 B.n646 B.n645 163.367
R737 B.n645 B.n644 163.367
R738 B.n644 B.n59 163.367
R739 B.n640 B.n59 163.367
R740 B.n640 B.n639 163.367
R741 B.n639 B.n638 163.367
R742 B.n638 B.n61 163.367
R743 B.n634 B.n61 163.367
R744 B.n634 B.n633 163.367
R745 B.n633 B.n632 163.367
R746 B.n632 B.n63 163.367
R747 B.n628 B.n63 163.367
R748 B.n628 B.n627 163.367
R749 B.n627 B.n626 163.367
R750 B.n626 B.n65 163.367
R751 B.n622 B.n65 163.367
R752 B.n622 B.n621 163.367
R753 B.n621 B.n620 163.367
R754 B.n620 B.n67 163.367
R755 B.n616 B.n67 163.367
R756 B.n616 B.n615 163.367
R757 B.n615 B.n614 163.367
R758 B.n614 B.n69 163.367
R759 B.n610 B.n69 163.367
R760 B.n610 B.n609 163.367
R761 B.n609 B.n608 163.367
R762 B.n608 B.n71 163.367
R763 B.n604 B.n71 163.367
R764 B.n604 B.n603 163.367
R765 B.n603 B.n602 163.367
R766 B.n602 B.n73 163.367
R767 B.n598 B.n73 163.367
R768 B.n598 B.n597 163.367
R769 B.n597 B.n596 163.367
R770 B.n596 B.n75 163.367
R771 B.n592 B.n75 163.367
R772 B.n592 B.n591 163.367
R773 B.n591 B.n590 163.367
R774 B.n590 B.n77 163.367
R775 B.n586 B.n77 163.367
R776 B.n586 B.n585 163.367
R777 B.n585 B.n584 163.367
R778 B.n584 B.n79 163.367
R779 B.n580 B.n79 163.367
R780 B.n580 B.n579 163.367
R781 B.n579 B.n578 163.367
R782 B.n578 B.n81 163.367
R783 B.n574 B.n81 163.367
R784 B.n574 B.n573 163.367
R785 B.n573 B.n572 163.367
R786 B.n572 B.n83 163.367
R787 B.n568 B.n83 163.367
R788 B.n568 B.n567 163.367
R789 B.n567 B.n566 163.367
R790 B.n566 B.n85 163.367
R791 B.n562 B.n85 163.367
R792 B.n562 B.n561 163.367
R793 B.n561 B.n560 163.367
R794 B.n560 B.n87 163.367
R795 B.n556 B.n87 163.367
R796 B.n556 B.n555 163.367
R797 B.n555 B.n554 163.367
R798 B.n554 B.n89 163.367
R799 B.n550 B.n89 163.367
R800 B.n762 B.n761 163.367
R801 B.n762 B.n15 163.367
R802 B.n766 B.n15 163.367
R803 B.n767 B.n766 163.367
R804 B.n768 B.n767 163.367
R805 B.n768 B.n13 163.367
R806 B.n772 B.n13 163.367
R807 B.n773 B.n772 163.367
R808 B.n774 B.n773 163.367
R809 B.n774 B.n11 163.367
R810 B.n778 B.n11 163.367
R811 B.n779 B.n778 163.367
R812 B.n780 B.n779 163.367
R813 B.n780 B.n9 163.367
R814 B.n784 B.n9 163.367
R815 B.n785 B.n784 163.367
R816 B.n786 B.n785 163.367
R817 B.n786 B.n7 163.367
R818 B.n790 B.n7 163.367
R819 B.n791 B.n790 163.367
R820 B.n792 B.n791 163.367
R821 B.n792 B.n5 163.367
R822 B.n796 B.n5 163.367
R823 B.n797 B.n796 163.367
R824 B.n798 B.n797 163.367
R825 B.n798 B.n3 163.367
R826 B.n802 B.n3 163.367
R827 B.n803 B.n802 163.367
R828 B.n205 B.n2 163.367
R829 B.n208 B.n205 163.367
R830 B.n209 B.n208 163.367
R831 B.n210 B.n209 163.367
R832 B.n210 B.n203 163.367
R833 B.n214 B.n203 163.367
R834 B.n215 B.n214 163.367
R835 B.n216 B.n215 163.367
R836 B.n216 B.n201 163.367
R837 B.n220 B.n201 163.367
R838 B.n221 B.n220 163.367
R839 B.n222 B.n221 163.367
R840 B.n222 B.n199 163.367
R841 B.n226 B.n199 163.367
R842 B.n227 B.n226 163.367
R843 B.n228 B.n227 163.367
R844 B.n228 B.n197 163.367
R845 B.n232 B.n197 163.367
R846 B.n233 B.n232 163.367
R847 B.n234 B.n233 163.367
R848 B.n234 B.n195 163.367
R849 B.n238 B.n195 163.367
R850 B.n239 B.n238 163.367
R851 B.n240 B.n239 163.367
R852 B.n240 B.n193 163.367
R853 B.n244 B.n193 163.367
R854 B.n245 B.n244 163.367
R855 B.n246 B.n245 163.367
R856 B.n358 B.t1 156.655
R857 B.n56 B.t8 156.655
R858 B.n158 B.t10 156.629
R859 B.n50 B.t5 156.629
R860 B.n359 B.t2 109.138
R861 B.n57 B.t7 109.138
R862 B.n159 B.t11 109.114
R863 B.n51 B.t4 109.114
R864 B.n345 B.n159 59.5399
R865 B.n360 B.n359 59.5399
R866 B.n648 B.n57 59.5399
R867 B.n662 B.n51 59.5399
R868 B.n159 B.n158 47.5157
R869 B.n359 B.n358 47.5157
R870 B.n57 B.n56 47.5157
R871 B.n51 B.n50 47.5157
R872 B.n461 B.n120 35.7468
R873 B.n759 B.n16 35.7468
R874 B.n551 B.n90 35.7468
R875 B.n248 B.n247 35.7468
R876 B B.n805 18.0485
R877 B.n763 B.n16 10.6151
R878 B.n764 B.n763 10.6151
R879 B.n765 B.n764 10.6151
R880 B.n765 B.n14 10.6151
R881 B.n769 B.n14 10.6151
R882 B.n770 B.n769 10.6151
R883 B.n771 B.n770 10.6151
R884 B.n771 B.n12 10.6151
R885 B.n775 B.n12 10.6151
R886 B.n776 B.n775 10.6151
R887 B.n777 B.n776 10.6151
R888 B.n777 B.n10 10.6151
R889 B.n781 B.n10 10.6151
R890 B.n782 B.n781 10.6151
R891 B.n783 B.n782 10.6151
R892 B.n783 B.n8 10.6151
R893 B.n787 B.n8 10.6151
R894 B.n788 B.n787 10.6151
R895 B.n789 B.n788 10.6151
R896 B.n789 B.n6 10.6151
R897 B.n793 B.n6 10.6151
R898 B.n794 B.n793 10.6151
R899 B.n795 B.n794 10.6151
R900 B.n795 B.n4 10.6151
R901 B.n799 B.n4 10.6151
R902 B.n800 B.n799 10.6151
R903 B.n801 B.n800 10.6151
R904 B.n801 B.n0 10.6151
R905 B.n759 B.n758 10.6151
R906 B.n758 B.n757 10.6151
R907 B.n757 B.n18 10.6151
R908 B.n753 B.n18 10.6151
R909 B.n753 B.n752 10.6151
R910 B.n752 B.n751 10.6151
R911 B.n751 B.n20 10.6151
R912 B.n747 B.n20 10.6151
R913 B.n747 B.n746 10.6151
R914 B.n746 B.n745 10.6151
R915 B.n745 B.n22 10.6151
R916 B.n741 B.n22 10.6151
R917 B.n741 B.n740 10.6151
R918 B.n740 B.n739 10.6151
R919 B.n739 B.n24 10.6151
R920 B.n735 B.n24 10.6151
R921 B.n735 B.n734 10.6151
R922 B.n734 B.n733 10.6151
R923 B.n733 B.n26 10.6151
R924 B.n729 B.n26 10.6151
R925 B.n729 B.n728 10.6151
R926 B.n728 B.n727 10.6151
R927 B.n727 B.n28 10.6151
R928 B.n723 B.n28 10.6151
R929 B.n723 B.n722 10.6151
R930 B.n722 B.n721 10.6151
R931 B.n721 B.n30 10.6151
R932 B.n717 B.n30 10.6151
R933 B.n717 B.n716 10.6151
R934 B.n716 B.n715 10.6151
R935 B.n715 B.n32 10.6151
R936 B.n711 B.n32 10.6151
R937 B.n711 B.n710 10.6151
R938 B.n710 B.n709 10.6151
R939 B.n709 B.n34 10.6151
R940 B.n705 B.n34 10.6151
R941 B.n705 B.n704 10.6151
R942 B.n704 B.n703 10.6151
R943 B.n703 B.n36 10.6151
R944 B.n699 B.n36 10.6151
R945 B.n699 B.n698 10.6151
R946 B.n698 B.n697 10.6151
R947 B.n697 B.n38 10.6151
R948 B.n693 B.n38 10.6151
R949 B.n693 B.n692 10.6151
R950 B.n692 B.n691 10.6151
R951 B.n691 B.n40 10.6151
R952 B.n687 B.n40 10.6151
R953 B.n687 B.n686 10.6151
R954 B.n686 B.n685 10.6151
R955 B.n685 B.n42 10.6151
R956 B.n681 B.n42 10.6151
R957 B.n681 B.n680 10.6151
R958 B.n680 B.n679 10.6151
R959 B.n679 B.n44 10.6151
R960 B.n675 B.n44 10.6151
R961 B.n675 B.n674 10.6151
R962 B.n674 B.n673 10.6151
R963 B.n673 B.n46 10.6151
R964 B.n669 B.n46 10.6151
R965 B.n669 B.n668 10.6151
R966 B.n668 B.n667 10.6151
R967 B.n667 B.n48 10.6151
R968 B.n663 B.n48 10.6151
R969 B.n661 B.n660 10.6151
R970 B.n660 B.n52 10.6151
R971 B.n656 B.n52 10.6151
R972 B.n656 B.n655 10.6151
R973 B.n655 B.n654 10.6151
R974 B.n654 B.n54 10.6151
R975 B.n650 B.n54 10.6151
R976 B.n650 B.n649 10.6151
R977 B.n647 B.n58 10.6151
R978 B.n643 B.n58 10.6151
R979 B.n643 B.n642 10.6151
R980 B.n642 B.n641 10.6151
R981 B.n641 B.n60 10.6151
R982 B.n637 B.n60 10.6151
R983 B.n637 B.n636 10.6151
R984 B.n636 B.n635 10.6151
R985 B.n635 B.n62 10.6151
R986 B.n631 B.n62 10.6151
R987 B.n631 B.n630 10.6151
R988 B.n630 B.n629 10.6151
R989 B.n629 B.n64 10.6151
R990 B.n625 B.n64 10.6151
R991 B.n625 B.n624 10.6151
R992 B.n624 B.n623 10.6151
R993 B.n623 B.n66 10.6151
R994 B.n619 B.n66 10.6151
R995 B.n619 B.n618 10.6151
R996 B.n618 B.n617 10.6151
R997 B.n617 B.n68 10.6151
R998 B.n613 B.n68 10.6151
R999 B.n613 B.n612 10.6151
R1000 B.n612 B.n611 10.6151
R1001 B.n611 B.n70 10.6151
R1002 B.n607 B.n70 10.6151
R1003 B.n607 B.n606 10.6151
R1004 B.n606 B.n605 10.6151
R1005 B.n605 B.n72 10.6151
R1006 B.n601 B.n72 10.6151
R1007 B.n601 B.n600 10.6151
R1008 B.n600 B.n599 10.6151
R1009 B.n599 B.n74 10.6151
R1010 B.n595 B.n74 10.6151
R1011 B.n595 B.n594 10.6151
R1012 B.n594 B.n593 10.6151
R1013 B.n593 B.n76 10.6151
R1014 B.n589 B.n76 10.6151
R1015 B.n589 B.n588 10.6151
R1016 B.n588 B.n587 10.6151
R1017 B.n587 B.n78 10.6151
R1018 B.n583 B.n78 10.6151
R1019 B.n583 B.n582 10.6151
R1020 B.n582 B.n581 10.6151
R1021 B.n581 B.n80 10.6151
R1022 B.n577 B.n80 10.6151
R1023 B.n577 B.n576 10.6151
R1024 B.n576 B.n575 10.6151
R1025 B.n575 B.n82 10.6151
R1026 B.n571 B.n82 10.6151
R1027 B.n571 B.n570 10.6151
R1028 B.n570 B.n569 10.6151
R1029 B.n569 B.n84 10.6151
R1030 B.n565 B.n84 10.6151
R1031 B.n565 B.n564 10.6151
R1032 B.n564 B.n563 10.6151
R1033 B.n563 B.n86 10.6151
R1034 B.n559 B.n86 10.6151
R1035 B.n559 B.n558 10.6151
R1036 B.n558 B.n557 10.6151
R1037 B.n557 B.n88 10.6151
R1038 B.n553 B.n88 10.6151
R1039 B.n553 B.n552 10.6151
R1040 B.n552 B.n551 10.6151
R1041 B.n547 B.n90 10.6151
R1042 B.n547 B.n546 10.6151
R1043 B.n546 B.n545 10.6151
R1044 B.n545 B.n92 10.6151
R1045 B.n541 B.n92 10.6151
R1046 B.n541 B.n540 10.6151
R1047 B.n540 B.n539 10.6151
R1048 B.n539 B.n94 10.6151
R1049 B.n535 B.n94 10.6151
R1050 B.n535 B.n534 10.6151
R1051 B.n534 B.n533 10.6151
R1052 B.n533 B.n96 10.6151
R1053 B.n529 B.n96 10.6151
R1054 B.n529 B.n528 10.6151
R1055 B.n528 B.n527 10.6151
R1056 B.n527 B.n98 10.6151
R1057 B.n523 B.n98 10.6151
R1058 B.n523 B.n522 10.6151
R1059 B.n522 B.n521 10.6151
R1060 B.n521 B.n100 10.6151
R1061 B.n517 B.n100 10.6151
R1062 B.n517 B.n516 10.6151
R1063 B.n516 B.n515 10.6151
R1064 B.n515 B.n102 10.6151
R1065 B.n511 B.n102 10.6151
R1066 B.n511 B.n510 10.6151
R1067 B.n510 B.n509 10.6151
R1068 B.n509 B.n104 10.6151
R1069 B.n505 B.n104 10.6151
R1070 B.n505 B.n504 10.6151
R1071 B.n504 B.n503 10.6151
R1072 B.n503 B.n106 10.6151
R1073 B.n499 B.n106 10.6151
R1074 B.n499 B.n498 10.6151
R1075 B.n498 B.n497 10.6151
R1076 B.n497 B.n108 10.6151
R1077 B.n493 B.n108 10.6151
R1078 B.n493 B.n492 10.6151
R1079 B.n492 B.n491 10.6151
R1080 B.n491 B.n110 10.6151
R1081 B.n487 B.n110 10.6151
R1082 B.n487 B.n486 10.6151
R1083 B.n486 B.n485 10.6151
R1084 B.n485 B.n112 10.6151
R1085 B.n481 B.n112 10.6151
R1086 B.n481 B.n480 10.6151
R1087 B.n480 B.n479 10.6151
R1088 B.n479 B.n114 10.6151
R1089 B.n475 B.n114 10.6151
R1090 B.n475 B.n474 10.6151
R1091 B.n474 B.n473 10.6151
R1092 B.n473 B.n116 10.6151
R1093 B.n469 B.n116 10.6151
R1094 B.n469 B.n468 10.6151
R1095 B.n468 B.n467 10.6151
R1096 B.n467 B.n118 10.6151
R1097 B.n463 B.n118 10.6151
R1098 B.n463 B.n462 10.6151
R1099 B.n462 B.n461 10.6151
R1100 B.n206 B.n1 10.6151
R1101 B.n207 B.n206 10.6151
R1102 B.n207 B.n204 10.6151
R1103 B.n211 B.n204 10.6151
R1104 B.n212 B.n211 10.6151
R1105 B.n213 B.n212 10.6151
R1106 B.n213 B.n202 10.6151
R1107 B.n217 B.n202 10.6151
R1108 B.n218 B.n217 10.6151
R1109 B.n219 B.n218 10.6151
R1110 B.n219 B.n200 10.6151
R1111 B.n223 B.n200 10.6151
R1112 B.n224 B.n223 10.6151
R1113 B.n225 B.n224 10.6151
R1114 B.n225 B.n198 10.6151
R1115 B.n229 B.n198 10.6151
R1116 B.n230 B.n229 10.6151
R1117 B.n231 B.n230 10.6151
R1118 B.n231 B.n196 10.6151
R1119 B.n235 B.n196 10.6151
R1120 B.n236 B.n235 10.6151
R1121 B.n237 B.n236 10.6151
R1122 B.n237 B.n194 10.6151
R1123 B.n241 B.n194 10.6151
R1124 B.n242 B.n241 10.6151
R1125 B.n243 B.n242 10.6151
R1126 B.n243 B.n192 10.6151
R1127 B.n247 B.n192 10.6151
R1128 B.n249 B.n248 10.6151
R1129 B.n249 B.n190 10.6151
R1130 B.n253 B.n190 10.6151
R1131 B.n254 B.n253 10.6151
R1132 B.n255 B.n254 10.6151
R1133 B.n255 B.n188 10.6151
R1134 B.n259 B.n188 10.6151
R1135 B.n260 B.n259 10.6151
R1136 B.n261 B.n260 10.6151
R1137 B.n261 B.n186 10.6151
R1138 B.n265 B.n186 10.6151
R1139 B.n266 B.n265 10.6151
R1140 B.n267 B.n266 10.6151
R1141 B.n267 B.n184 10.6151
R1142 B.n271 B.n184 10.6151
R1143 B.n272 B.n271 10.6151
R1144 B.n273 B.n272 10.6151
R1145 B.n273 B.n182 10.6151
R1146 B.n277 B.n182 10.6151
R1147 B.n278 B.n277 10.6151
R1148 B.n279 B.n278 10.6151
R1149 B.n279 B.n180 10.6151
R1150 B.n283 B.n180 10.6151
R1151 B.n284 B.n283 10.6151
R1152 B.n285 B.n284 10.6151
R1153 B.n285 B.n178 10.6151
R1154 B.n289 B.n178 10.6151
R1155 B.n290 B.n289 10.6151
R1156 B.n291 B.n290 10.6151
R1157 B.n291 B.n176 10.6151
R1158 B.n295 B.n176 10.6151
R1159 B.n296 B.n295 10.6151
R1160 B.n297 B.n296 10.6151
R1161 B.n297 B.n174 10.6151
R1162 B.n301 B.n174 10.6151
R1163 B.n302 B.n301 10.6151
R1164 B.n303 B.n302 10.6151
R1165 B.n303 B.n172 10.6151
R1166 B.n307 B.n172 10.6151
R1167 B.n308 B.n307 10.6151
R1168 B.n309 B.n308 10.6151
R1169 B.n309 B.n170 10.6151
R1170 B.n313 B.n170 10.6151
R1171 B.n314 B.n313 10.6151
R1172 B.n315 B.n314 10.6151
R1173 B.n315 B.n168 10.6151
R1174 B.n319 B.n168 10.6151
R1175 B.n320 B.n319 10.6151
R1176 B.n321 B.n320 10.6151
R1177 B.n321 B.n166 10.6151
R1178 B.n325 B.n166 10.6151
R1179 B.n326 B.n325 10.6151
R1180 B.n327 B.n326 10.6151
R1181 B.n327 B.n164 10.6151
R1182 B.n331 B.n164 10.6151
R1183 B.n332 B.n331 10.6151
R1184 B.n333 B.n332 10.6151
R1185 B.n333 B.n162 10.6151
R1186 B.n337 B.n162 10.6151
R1187 B.n338 B.n337 10.6151
R1188 B.n339 B.n338 10.6151
R1189 B.n339 B.n160 10.6151
R1190 B.n343 B.n160 10.6151
R1191 B.n344 B.n343 10.6151
R1192 B.n346 B.n156 10.6151
R1193 B.n350 B.n156 10.6151
R1194 B.n351 B.n350 10.6151
R1195 B.n352 B.n351 10.6151
R1196 B.n352 B.n154 10.6151
R1197 B.n356 B.n154 10.6151
R1198 B.n357 B.n356 10.6151
R1199 B.n361 B.n357 10.6151
R1200 B.n365 B.n152 10.6151
R1201 B.n366 B.n365 10.6151
R1202 B.n367 B.n366 10.6151
R1203 B.n367 B.n150 10.6151
R1204 B.n371 B.n150 10.6151
R1205 B.n372 B.n371 10.6151
R1206 B.n373 B.n372 10.6151
R1207 B.n373 B.n148 10.6151
R1208 B.n377 B.n148 10.6151
R1209 B.n378 B.n377 10.6151
R1210 B.n379 B.n378 10.6151
R1211 B.n379 B.n146 10.6151
R1212 B.n383 B.n146 10.6151
R1213 B.n384 B.n383 10.6151
R1214 B.n385 B.n384 10.6151
R1215 B.n385 B.n144 10.6151
R1216 B.n389 B.n144 10.6151
R1217 B.n390 B.n389 10.6151
R1218 B.n391 B.n390 10.6151
R1219 B.n391 B.n142 10.6151
R1220 B.n395 B.n142 10.6151
R1221 B.n396 B.n395 10.6151
R1222 B.n397 B.n396 10.6151
R1223 B.n397 B.n140 10.6151
R1224 B.n401 B.n140 10.6151
R1225 B.n402 B.n401 10.6151
R1226 B.n403 B.n402 10.6151
R1227 B.n403 B.n138 10.6151
R1228 B.n407 B.n138 10.6151
R1229 B.n408 B.n407 10.6151
R1230 B.n409 B.n408 10.6151
R1231 B.n409 B.n136 10.6151
R1232 B.n413 B.n136 10.6151
R1233 B.n414 B.n413 10.6151
R1234 B.n415 B.n414 10.6151
R1235 B.n415 B.n134 10.6151
R1236 B.n419 B.n134 10.6151
R1237 B.n420 B.n419 10.6151
R1238 B.n421 B.n420 10.6151
R1239 B.n421 B.n132 10.6151
R1240 B.n425 B.n132 10.6151
R1241 B.n426 B.n425 10.6151
R1242 B.n427 B.n426 10.6151
R1243 B.n427 B.n130 10.6151
R1244 B.n431 B.n130 10.6151
R1245 B.n432 B.n431 10.6151
R1246 B.n433 B.n432 10.6151
R1247 B.n433 B.n128 10.6151
R1248 B.n437 B.n128 10.6151
R1249 B.n438 B.n437 10.6151
R1250 B.n439 B.n438 10.6151
R1251 B.n439 B.n126 10.6151
R1252 B.n443 B.n126 10.6151
R1253 B.n444 B.n443 10.6151
R1254 B.n445 B.n444 10.6151
R1255 B.n445 B.n124 10.6151
R1256 B.n449 B.n124 10.6151
R1257 B.n450 B.n449 10.6151
R1258 B.n451 B.n450 10.6151
R1259 B.n451 B.n122 10.6151
R1260 B.n455 B.n122 10.6151
R1261 B.n456 B.n455 10.6151
R1262 B.n457 B.n456 10.6151
R1263 B.n457 B.n120 10.6151
R1264 B.n805 B.n0 8.11757
R1265 B.n805 B.n1 8.11757
R1266 B.n662 B.n661 6.5566
R1267 B.n649 B.n648 6.5566
R1268 B.n346 B.n345 6.5566
R1269 B.n361 B.n360 6.5566
R1270 B.n663 B.n662 4.05904
R1271 B.n648 B.n647 4.05904
R1272 B.n345 B.n344 4.05904
R1273 B.n360 B.n152 4.05904
C0 VDD1 w_n2440_n4944# 1.57344f
C1 w_n2440_n4944# VN 4.1781f
C2 VDD2 w_n2440_n4944# 1.61882f
C3 VDD1 B 1.39054f
C4 B VN 1.11355f
C5 VDD2 B 1.43481f
C6 VDD1 VTAIL 7.40762f
C7 VDD1 VP 7.56882f
C8 VTAIL VN 6.86691f
C9 VP VN 7.29807f
C10 VDD2 VTAIL 7.45861f
C11 VDD2 VP 0.364223f
C12 B w_n2440_n4944# 10.8648f
C13 w_n2440_n4944# VTAIL 5.77442f
C14 VP w_n2440_n4944# 4.49056f
C15 B VTAIL 7.2228f
C16 VP B 1.62982f
C17 VDD1 VN 0.149027f
C18 VDD2 VDD1 0.913864f
C19 VP VTAIL 6.88102f
C20 VDD2 VN 7.35424f
C21 VDD2 VSUBS 1.055064f
C22 VDD1 VSUBS 6.474979f
C23 VTAIL VSUBS 1.543272f
C24 VN VSUBS 5.63517f
C25 VP VSUBS 2.333189f
C26 B VSUBS 4.523482f
C27 w_n2440_n4944# VSUBS 0.147308p
C28 B.n0 VSUBS 0.005508f
C29 B.n1 VSUBS 0.005508f
C30 B.n2 VSUBS 0.008146f
C31 B.n3 VSUBS 0.006242f
C32 B.n4 VSUBS 0.006242f
C33 B.n5 VSUBS 0.006242f
C34 B.n6 VSUBS 0.006242f
C35 B.n7 VSUBS 0.006242f
C36 B.n8 VSUBS 0.006242f
C37 B.n9 VSUBS 0.006242f
C38 B.n10 VSUBS 0.006242f
C39 B.n11 VSUBS 0.006242f
C40 B.n12 VSUBS 0.006242f
C41 B.n13 VSUBS 0.006242f
C42 B.n14 VSUBS 0.006242f
C43 B.n15 VSUBS 0.006242f
C44 B.n16 VSUBS 0.015112f
C45 B.n17 VSUBS 0.006242f
C46 B.n18 VSUBS 0.006242f
C47 B.n19 VSUBS 0.006242f
C48 B.n20 VSUBS 0.006242f
C49 B.n21 VSUBS 0.006242f
C50 B.n22 VSUBS 0.006242f
C51 B.n23 VSUBS 0.006242f
C52 B.n24 VSUBS 0.006242f
C53 B.n25 VSUBS 0.006242f
C54 B.n26 VSUBS 0.006242f
C55 B.n27 VSUBS 0.006242f
C56 B.n28 VSUBS 0.006242f
C57 B.n29 VSUBS 0.006242f
C58 B.n30 VSUBS 0.006242f
C59 B.n31 VSUBS 0.006242f
C60 B.n32 VSUBS 0.006242f
C61 B.n33 VSUBS 0.006242f
C62 B.n34 VSUBS 0.006242f
C63 B.n35 VSUBS 0.006242f
C64 B.n36 VSUBS 0.006242f
C65 B.n37 VSUBS 0.006242f
C66 B.n38 VSUBS 0.006242f
C67 B.n39 VSUBS 0.006242f
C68 B.n40 VSUBS 0.006242f
C69 B.n41 VSUBS 0.006242f
C70 B.n42 VSUBS 0.006242f
C71 B.n43 VSUBS 0.006242f
C72 B.n44 VSUBS 0.006242f
C73 B.n45 VSUBS 0.006242f
C74 B.n46 VSUBS 0.006242f
C75 B.n47 VSUBS 0.006242f
C76 B.n48 VSUBS 0.006242f
C77 B.n49 VSUBS 0.006242f
C78 B.t4 VSUBS 0.602474f
C79 B.t5 VSUBS 0.61876f
C80 B.t3 VSUBS 1.63029f
C81 B.n50 VSUBS 0.31741f
C82 B.n51 VSUBS 0.06259f
C83 B.n52 VSUBS 0.006242f
C84 B.n53 VSUBS 0.006242f
C85 B.n54 VSUBS 0.006242f
C86 B.n55 VSUBS 0.006242f
C87 B.t7 VSUBS 0.602448f
C88 B.t8 VSUBS 0.61874f
C89 B.t6 VSUBS 1.63029f
C90 B.n56 VSUBS 0.31743f
C91 B.n57 VSUBS 0.062615f
C92 B.n58 VSUBS 0.006242f
C93 B.n59 VSUBS 0.006242f
C94 B.n60 VSUBS 0.006242f
C95 B.n61 VSUBS 0.006242f
C96 B.n62 VSUBS 0.006242f
C97 B.n63 VSUBS 0.006242f
C98 B.n64 VSUBS 0.006242f
C99 B.n65 VSUBS 0.006242f
C100 B.n66 VSUBS 0.006242f
C101 B.n67 VSUBS 0.006242f
C102 B.n68 VSUBS 0.006242f
C103 B.n69 VSUBS 0.006242f
C104 B.n70 VSUBS 0.006242f
C105 B.n71 VSUBS 0.006242f
C106 B.n72 VSUBS 0.006242f
C107 B.n73 VSUBS 0.006242f
C108 B.n74 VSUBS 0.006242f
C109 B.n75 VSUBS 0.006242f
C110 B.n76 VSUBS 0.006242f
C111 B.n77 VSUBS 0.006242f
C112 B.n78 VSUBS 0.006242f
C113 B.n79 VSUBS 0.006242f
C114 B.n80 VSUBS 0.006242f
C115 B.n81 VSUBS 0.006242f
C116 B.n82 VSUBS 0.006242f
C117 B.n83 VSUBS 0.006242f
C118 B.n84 VSUBS 0.006242f
C119 B.n85 VSUBS 0.006242f
C120 B.n86 VSUBS 0.006242f
C121 B.n87 VSUBS 0.006242f
C122 B.n88 VSUBS 0.006242f
C123 B.n89 VSUBS 0.006242f
C124 B.n90 VSUBS 0.015112f
C125 B.n91 VSUBS 0.006242f
C126 B.n92 VSUBS 0.006242f
C127 B.n93 VSUBS 0.006242f
C128 B.n94 VSUBS 0.006242f
C129 B.n95 VSUBS 0.006242f
C130 B.n96 VSUBS 0.006242f
C131 B.n97 VSUBS 0.006242f
C132 B.n98 VSUBS 0.006242f
C133 B.n99 VSUBS 0.006242f
C134 B.n100 VSUBS 0.006242f
C135 B.n101 VSUBS 0.006242f
C136 B.n102 VSUBS 0.006242f
C137 B.n103 VSUBS 0.006242f
C138 B.n104 VSUBS 0.006242f
C139 B.n105 VSUBS 0.006242f
C140 B.n106 VSUBS 0.006242f
C141 B.n107 VSUBS 0.006242f
C142 B.n108 VSUBS 0.006242f
C143 B.n109 VSUBS 0.006242f
C144 B.n110 VSUBS 0.006242f
C145 B.n111 VSUBS 0.006242f
C146 B.n112 VSUBS 0.006242f
C147 B.n113 VSUBS 0.006242f
C148 B.n114 VSUBS 0.006242f
C149 B.n115 VSUBS 0.006242f
C150 B.n116 VSUBS 0.006242f
C151 B.n117 VSUBS 0.006242f
C152 B.n118 VSUBS 0.006242f
C153 B.n119 VSUBS 0.006242f
C154 B.n120 VSUBS 0.015243f
C155 B.n121 VSUBS 0.006242f
C156 B.n122 VSUBS 0.006242f
C157 B.n123 VSUBS 0.006242f
C158 B.n124 VSUBS 0.006242f
C159 B.n125 VSUBS 0.006242f
C160 B.n126 VSUBS 0.006242f
C161 B.n127 VSUBS 0.006242f
C162 B.n128 VSUBS 0.006242f
C163 B.n129 VSUBS 0.006242f
C164 B.n130 VSUBS 0.006242f
C165 B.n131 VSUBS 0.006242f
C166 B.n132 VSUBS 0.006242f
C167 B.n133 VSUBS 0.006242f
C168 B.n134 VSUBS 0.006242f
C169 B.n135 VSUBS 0.006242f
C170 B.n136 VSUBS 0.006242f
C171 B.n137 VSUBS 0.006242f
C172 B.n138 VSUBS 0.006242f
C173 B.n139 VSUBS 0.006242f
C174 B.n140 VSUBS 0.006242f
C175 B.n141 VSUBS 0.006242f
C176 B.n142 VSUBS 0.006242f
C177 B.n143 VSUBS 0.006242f
C178 B.n144 VSUBS 0.006242f
C179 B.n145 VSUBS 0.006242f
C180 B.n146 VSUBS 0.006242f
C181 B.n147 VSUBS 0.006242f
C182 B.n148 VSUBS 0.006242f
C183 B.n149 VSUBS 0.006242f
C184 B.n150 VSUBS 0.006242f
C185 B.n151 VSUBS 0.006242f
C186 B.n152 VSUBS 0.004315f
C187 B.n153 VSUBS 0.006242f
C188 B.n154 VSUBS 0.006242f
C189 B.n155 VSUBS 0.006242f
C190 B.n156 VSUBS 0.006242f
C191 B.n157 VSUBS 0.006242f
C192 B.t11 VSUBS 0.602474f
C193 B.t10 VSUBS 0.61876f
C194 B.t9 VSUBS 1.63029f
C195 B.n158 VSUBS 0.31741f
C196 B.n159 VSUBS 0.06259f
C197 B.n160 VSUBS 0.006242f
C198 B.n161 VSUBS 0.006242f
C199 B.n162 VSUBS 0.006242f
C200 B.n163 VSUBS 0.006242f
C201 B.n164 VSUBS 0.006242f
C202 B.n165 VSUBS 0.006242f
C203 B.n166 VSUBS 0.006242f
C204 B.n167 VSUBS 0.006242f
C205 B.n168 VSUBS 0.006242f
C206 B.n169 VSUBS 0.006242f
C207 B.n170 VSUBS 0.006242f
C208 B.n171 VSUBS 0.006242f
C209 B.n172 VSUBS 0.006242f
C210 B.n173 VSUBS 0.006242f
C211 B.n174 VSUBS 0.006242f
C212 B.n175 VSUBS 0.006242f
C213 B.n176 VSUBS 0.006242f
C214 B.n177 VSUBS 0.006242f
C215 B.n178 VSUBS 0.006242f
C216 B.n179 VSUBS 0.006242f
C217 B.n180 VSUBS 0.006242f
C218 B.n181 VSUBS 0.006242f
C219 B.n182 VSUBS 0.006242f
C220 B.n183 VSUBS 0.006242f
C221 B.n184 VSUBS 0.006242f
C222 B.n185 VSUBS 0.006242f
C223 B.n186 VSUBS 0.006242f
C224 B.n187 VSUBS 0.006242f
C225 B.n188 VSUBS 0.006242f
C226 B.n189 VSUBS 0.006242f
C227 B.n190 VSUBS 0.006242f
C228 B.n191 VSUBS 0.015917f
C229 B.n192 VSUBS 0.006242f
C230 B.n193 VSUBS 0.006242f
C231 B.n194 VSUBS 0.006242f
C232 B.n195 VSUBS 0.006242f
C233 B.n196 VSUBS 0.006242f
C234 B.n197 VSUBS 0.006242f
C235 B.n198 VSUBS 0.006242f
C236 B.n199 VSUBS 0.006242f
C237 B.n200 VSUBS 0.006242f
C238 B.n201 VSUBS 0.006242f
C239 B.n202 VSUBS 0.006242f
C240 B.n203 VSUBS 0.006242f
C241 B.n204 VSUBS 0.006242f
C242 B.n205 VSUBS 0.006242f
C243 B.n206 VSUBS 0.006242f
C244 B.n207 VSUBS 0.006242f
C245 B.n208 VSUBS 0.006242f
C246 B.n209 VSUBS 0.006242f
C247 B.n210 VSUBS 0.006242f
C248 B.n211 VSUBS 0.006242f
C249 B.n212 VSUBS 0.006242f
C250 B.n213 VSUBS 0.006242f
C251 B.n214 VSUBS 0.006242f
C252 B.n215 VSUBS 0.006242f
C253 B.n216 VSUBS 0.006242f
C254 B.n217 VSUBS 0.006242f
C255 B.n218 VSUBS 0.006242f
C256 B.n219 VSUBS 0.006242f
C257 B.n220 VSUBS 0.006242f
C258 B.n221 VSUBS 0.006242f
C259 B.n222 VSUBS 0.006242f
C260 B.n223 VSUBS 0.006242f
C261 B.n224 VSUBS 0.006242f
C262 B.n225 VSUBS 0.006242f
C263 B.n226 VSUBS 0.006242f
C264 B.n227 VSUBS 0.006242f
C265 B.n228 VSUBS 0.006242f
C266 B.n229 VSUBS 0.006242f
C267 B.n230 VSUBS 0.006242f
C268 B.n231 VSUBS 0.006242f
C269 B.n232 VSUBS 0.006242f
C270 B.n233 VSUBS 0.006242f
C271 B.n234 VSUBS 0.006242f
C272 B.n235 VSUBS 0.006242f
C273 B.n236 VSUBS 0.006242f
C274 B.n237 VSUBS 0.006242f
C275 B.n238 VSUBS 0.006242f
C276 B.n239 VSUBS 0.006242f
C277 B.n240 VSUBS 0.006242f
C278 B.n241 VSUBS 0.006242f
C279 B.n242 VSUBS 0.006242f
C280 B.n243 VSUBS 0.006242f
C281 B.n244 VSUBS 0.006242f
C282 B.n245 VSUBS 0.006242f
C283 B.n246 VSUBS 0.015112f
C284 B.n247 VSUBS 0.015112f
C285 B.n248 VSUBS 0.015917f
C286 B.n249 VSUBS 0.006242f
C287 B.n250 VSUBS 0.006242f
C288 B.n251 VSUBS 0.006242f
C289 B.n252 VSUBS 0.006242f
C290 B.n253 VSUBS 0.006242f
C291 B.n254 VSUBS 0.006242f
C292 B.n255 VSUBS 0.006242f
C293 B.n256 VSUBS 0.006242f
C294 B.n257 VSUBS 0.006242f
C295 B.n258 VSUBS 0.006242f
C296 B.n259 VSUBS 0.006242f
C297 B.n260 VSUBS 0.006242f
C298 B.n261 VSUBS 0.006242f
C299 B.n262 VSUBS 0.006242f
C300 B.n263 VSUBS 0.006242f
C301 B.n264 VSUBS 0.006242f
C302 B.n265 VSUBS 0.006242f
C303 B.n266 VSUBS 0.006242f
C304 B.n267 VSUBS 0.006242f
C305 B.n268 VSUBS 0.006242f
C306 B.n269 VSUBS 0.006242f
C307 B.n270 VSUBS 0.006242f
C308 B.n271 VSUBS 0.006242f
C309 B.n272 VSUBS 0.006242f
C310 B.n273 VSUBS 0.006242f
C311 B.n274 VSUBS 0.006242f
C312 B.n275 VSUBS 0.006242f
C313 B.n276 VSUBS 0.006242f
C314 B.n277 VSUBS 0.006242f
C315 B.n278 VSUBS 0.006242f
C316 B.n279 VSUBS 0.006242f
C317 B.n280 VSUBS 0.006242f
C318 B.n281 VSUBS 0.006242f
C319 B.n282 VSUBS 0.006242f
C320 B.n283 VSUBS 0.006242f
C321 B.n284 VSUBS 0.006242f
C322 B.n285 VSUBS 0.006242f
C323 B.n286 VSUBS 0.006242f
C324 B.n287 VSUBS 0.006242f
C325 B.n288 VSUBS 0.006242f
C326 B.n289 VSUBS 0.006242f
C327 B.n290 VSUBS 0.006242f
C328 B.n291 VSUBS 0.006242f
C329 B.n292 VSUBS 0.006242f
C330 B.n293 VSUBS 0.006242f
C331 B.n294 VSUBS 0.006242f
C332 B.n295 VSUBS 0.006242f
C333 B.n296 VSUBS 0.006242f
C334 B.n297 VSUBS 0.006242f
C335 B.n298 VSUBS 0.006242f
C336 B.n299 VSUBS 0.006242f
C337 B.n300 VSUBS 0.006242f
C338 B.n301 VSUBS 0.006242f
C339 B.n302 VSUBS 0.006242f
C340 B.n303 VSUBS 0.006242f
C341 B.n304 VSUBS 0.006242f
C342 B.n305 VSUBS 0.006242f
C343 B.n306 VSUBS 0.006242f
C344 B.n307 VSUBS 0.006242f
C345 B.n308 VSUBS 0.006242f
C346 B.n309 VSUBS 0.006242f
C347 B.n310 VSUBS 0.006242f
C348 B.n311 VSUBS 0.006242f
C349 B.n312 VSUBS 0.006242f
C350 B.n313 VSUBS 0.006242f
C351 B.n314 VSUBS 0.006242f
C352 B.n315 VSUBS 0.006242f
C353 B.n316 VSUBS 0.006242f
C354 B.n317 VSUBS 0.006242f
C355 B.n318 VSUBS 0.006242f
C356 B.n319 VSUBS 0.006242f
C357 B.n320 VSUBS 0.006242f
C358 B.n321 VSUBS 0.006242f
C359 B.n322 VSUBS 0.006242f
C360 B.n323 VSUBS 0.006242f
C361 B.n324 VSUBS 0.006242f
C362 B.n325 VSUBS 0.006242f
C363 B.n326 VSUBS 0.006242f
C364 B.n327 VSUBS 0.006242f
C365 B.n328 VSUBS 0.006242f
C366 B.n329 VSUBS 0.006242f
C367 B.n330 VSUBS 0.006242f
C368 B.n331 VSUBS 0.006242f
C369 B.n332 VSUBS 0.006242f
C370 B.n333 VSUBS 0.006242f
C371 B.n334 VSUBS 0.006242f
C372 B.n335 VSUBS 0.006242f
C373 B.n336 VSUBS 0.006242f
C374 B.n337 VSUBS 0.006242f
C375 B.n338 VSUBS 0.006242f
C376 B.n339 VSUBS 0.006242f
C377 B.n340 VSUBS 0.006242f
C378 B.n341 VSUBS 0.006242f
C379 B.n342 VSUBS 0.006242f
C380 B.n343 VSUBS 0.006242f
C381 B.n344 VSUBS 0.004315f
C382 B.n345 VSUBS 0.014463f
C383 B.n346 VSUBS 0.005049f
C384 B.n347 VSUBS 0.006242f
C385 B.n348 VSUBS 0.006242f
C386 B.n349 VSUBS 0.006242f
C387 B.n350 VSUBS 0.006242f
C388 B.n351 VSUBS 0.006242f
C389 B.n352 VSUBS 0.006242f
C390 B.n353 VSUBS 0.006242f
C391 B.n354 VSUBS 0.006242f
C392 B.n355 VSUBS 0.006242f
C393 B.n356 VSUBS 0.006242f
C394 B.n357 VSUBS 0.006242f
C395 B.t2 VSUBS 0.602448f
C396 B.t1 VSUBS 0.61874f
C397 B.t0 VSUBS 1.63029f
C398 B.n358 VSUBS 0.31743f
C399 B.n359 VSUBS 0.062615f
C400 B.n360 VSUBS 0.014463f
C401 B.n361 VSUBS 0.005049f
C402 B.n362 VSUBS 0.006242f
C403 B.n363 VSUBS 0.006242f
C404 B.n364 VSUBS 0.006242f
C405 B.n365 VSUBS 0.006242f
C406 B.n366 VSUBS 0.006242f
C407 B.n367 VSUBS 0.006242f
C408 B.n368 VSUBS 0.006242f
C409 B.n369 VSUBS 0.006242f
C410 B.n370 VSUBS 0.006242f
C411 B.n371 VSUBS 0.006242f
C412 B.n372 VSUBS 0.006242f
C413 B.n373 VSUBS 0.006242f
C414 B.n374 VSUBS 0.006242f
C415 B.n375 VSUBS 0.006242f
C416 B.n376 VSUBS 0.006242f
C417 B.n377 VSUBS 0.006242f
C418 B.n378 VSUBS 0.006242f
C419 B.n379 VSUBS 0.006242f
C420 B.n380 VSUBS 0.006242f
C421 B.n381 VSUBS 0.006242f
C422 B.n382 VSUBS 0.006242f
C423 B.n383 VSUBS 0.006242f
C424 B.n384 VSUBS 0.006242f
C425 B.n385 VSUBS 0.006242f
C426 B.n386 VSUBS 0.006242f
C427 B.n387 VSUBS 0.006242f
C428 B.n388 VSUBS 0.006242f
C429 B.n389 VSUBS 0.006242f
C430 B.n390 VSUBS 0.006242f
C431 B.n391 VSUBS 0.006242f
C432 B.n392 VSUBS 0.006242f
C433 B.n393 VSUBS 0.006242f
C434 B.n394 VSUBS 0.006242f
C435 B.n395 VSUBS 0.006242f
C436 B.n396 VSUBS 0.006242f
C437 B.n397 VSUBS 0.006242f
C438 B.n398 VSUBS 0.006242f
C439 B.n399 VSUBS 0.006242f
C440 B.n400 VSUBS 0.006242f
C441 B.n401 VSUBS 0.006242f
C442 B.n402 VSUBS 0.006242f
C443 B.n403 VSUBS 0.006242f
C444 B.n404 VSUBS 0.006242f
C445 B.n405 VSUBS 0.006242f
C446 B.n406 VSUBS 0.006242f
C447 B.n407 VSUBS 0.006242f
C448 B.n408 VSUBS 0.006242f
C449 B.n409 VSUBS 0.006242f
C450 B.n410 VSUBS 0.006242f
C451 B.n411 VSUBS 0.006242f
C452 B.n412 VSUBS 0.006242f
C453 B.n413 VSUBS 0.006242f
C454 B.n414 VSUBS 0.006242f
C455 B.n415 VSUBS 0.006242f
C456 B.n416 VSUBS 0.006242f
C457 B.n417 VSUBS 0.006242f
C458 B.n418 VSUBS 0.006242f
C459 B.n419 VSUBS 0.006242f
C460 B.n420 VSUBS 0.006242f
C461 B.n421 VSUBS 0.006242f
C462 B.n422 VSUBS 0.006242f
C463 B.n423 VSUBS 0.006242f
C464 B.n424 VSUBS 0.006242f
C465 B.n425 VSUBS 0.006242f
C466 B.n426 VSUBS 0.006242f
C467 B.n427 VSUBS 0.006242f
C468 B.n428 VSUBS 0.006242f
C469 B.n429 VSUBS 0.006242f
C470 B.n430 VSUBS 0.006242f
C471 B.n431 VSUBS 0.006242f
C472 B.n432 VSUBS 0.006242f
C473 B.n433 VSUBS 0.006242f
C474 B.n434 VSUBS 0.006242f
C475 B.n435 VSUBS 0.006242f
C476 B.n436 VSUBS 0.006242f
C477 B.n437 VSUBS 0.006242f
C478 B.n438 VSUBS 0.006242f
C479 B.n439 VSUBS 0.006242f
C480 B.n440 VSUBS 0.006242f
C481 B.n441 VSUBS 0.006242f
C482 B.n442 VSUBS 0.006242f
C483 B.n443 VSUBS 0.006242f
C484 B.n444 VSUBS 0.006242f
C485 B.n445 VSUBS 0.006242f
C486 B.n446 VSUBS 0.006242f
C487 B.n447 VSUBS 0.006242f
C488 B.n448 VSUBS 0.006242f
C489 B.n449 VSUBS 0.006242f
C490 B.n450 VSUBS 0.006242f
C491 B.n451 VSUBS 0.006242f
C492 B.n452 VSUBS 0.006242f
C493 B.n453 VSUBS 0.006242f
C494 B.n454 VSUBS 0.006242f
C495 B.n455 VSUBS 0.006242f
C496 B.n456 VSUBS 0.006242f
C497 B.n457 VSUBS 0.006242f
C498 B.n458 VSUBS 0.006242f
C499 B.n459 VSUBS 0.015917f
C500 B.n460 VSUBS 0.015112f
C501 B.n461 VSUBS 0.015786f
C502 B.n462 VSUBS 0.006242f
C503 B.n463 VSUBS 0.006242f
C504 B.n464 VSUBS 0.006242f
C505 B.n465 VSUBS 0.006242f
C506 B.n466 VSUBS 0.006242f
C507 B.n467 VSUBS 0.006242f
C508 B.n468 VSUBS 0.006242f
C509 B.n469 VSUBS 0.006242f
C510 B.n470 VSUBS 0.006242f
C511 B.n471 VSUBS 0.006242f
C512 B.n472 VSUBS 0.006242f
C513 B.n473 VSUBS 0.006242f
C514 B.n474 VSUBS 0.006242f
C515 B.n475 VSUBS 0.006242f
C516 B.n476 VSUBS 0.006242f
C517 B.n477 VSUBS 0.006242f
C518 B.n478 VSUBS 0.006242f
C519 B.n479 VSUBS 0.006242f
C520 B.n480 VSUBS 0.006242f
C521 B.n481 VSUBS 0.006242f
C522 B.n482 VSUBS 0.006242f
C523 B.n483 VSUBS 0.006242f
C524 B.n484 VSUBS 0.006242f
C525 B.n485 VSUBS 0.006242f
C526 B.n486 VSUBS 0.006242f
C527 B.n487 VSUBS 0.006242f
C528 B.n488 VSUBS 0.006242f
C529 B.n489 VSUBS 0.006242f
C530 B.n490 VSUBS 0.006242f
C531 B.n491 VSUBS 0.006242f
C532 B.n492 VSUBS 0.006242f
C533 B.n493 VSUBS 0.006242f
C534 B.n494 VSUBS 0.006242f
C535 B.n495 VSUBS 0.006242f
C536 B.n496 VSUBS 0.006242f
C537 B.n497 VSUBS 0.006242f
C538 B.n498 VSUBS 0.006242f
C539 B.n499 VSUBS 0.006242f
C540 B.n500 VSUBS 0.006242f
C541 B.n501 VSUBS 0.006242f
C542 B.n502 VSUBS 0.006242f
C543 B.n503 VSUBS 0.006242f
C544 B.n504 VSUBS 0.006242f
C545 B.n505 VSUBS 0.006242f
C546 B.n506 VSUBS 0.006242f
C547 B.n507 VSUBS 0.006242f
C548 B.n508 VSUBS 0.006242f
C549 B.n509 VSUBS 0.006242f
C550 B.n510 VSUBS 0.006242f
C551 B.n511 VSUBS 0.006242f
C552 B.n512 VSUBS 0.006242f
C553 B.n513 VSUBS 0.006242f
C554 B.n514 VSUBS 0.006242f
C555 B.n515 VSUBS 0.006242f
C556 B.n516 VSUBS 0.006242f
C557 B.n517 VSUBS 0.006242f
C558 B.n518 VSUBS 0.006242f
C559 B.n519 VSUBS 0.006242f
C560 B.n520 VSUBS 0.006242f
C561 B.n521 VSUBS 0.006242f
C562 B.n522 VSUBS 0.006242f
C563 B.n523 VSUBS 0.006242f
C564 B.n524 VSUBS 0.006242f
C565 B.n525 VSUBS 0.006242f
C566 B.n526 VSUBS 0.006242f
C567 B.n527 VSUBS 0.006242f
C568 B.n528 VSUBS 0.006242f
C569 B.n529 VSUBS 0.006242f
C570 B.n530 VSUBS 0.006242f
C571 B.n531 VSUBS 0.006242f
C572 B.n532 VSUBS 0.006242f
C573 B.n533 VSUBS 0.006242f
C574 B.n534 VSUBS 0.006242f
C575 B.n535 VSUBS 0.006242f
C576 B.n536 VSUBS 0.006242f
C577 B.n537 VSUBS 0.006242f
C578 B.n538 VSUBS 0.006242f
C579 B.n539 VSUBS 0.006242f
C580 B.n540 VSUBS 0.006242f
C581 B.n541 VSUBS 0.006242f
C582 B.n542 VSUBS 0.006242f
C583 B.n543 VSUBS 0.006242f
C584 B.n544 VSUBS 0.006242f
C585 B.n545 VSUBS 0.006242f
C586 B.n546 VSUBS 0.006242f
C587 B.n547 VSUBS 0.006242f
C588 B.n548 VSUBS 0.006242f
C589 B.n549 VSUBS 0.015112f
C590 B.n550 VSUBS 0.015917f
C591 B.n551 VSUBS 0.015917f
C592 B.n552 VSUBS 0.006242f
C593 B.n553 VSUBS 0.006242f
C594 B.n554 VSUBS 0.006242f
C595 B.n555 VSUBS 0.006242f
C596 B.n556 VSUBS 0.006242f
C597 B.n557 VSUBS 0.006242f
C598 B.n558 VSUBS 0.006242f
C599 B.n559 VSUBS 0.006242f
C600 B.n560 VSUBS 0.006242f
C601 B.n561 VSUBS 0.006242f
C602 B.n562 VSUBS 0.006242f
C603 B.n563 VSUBS 0.006242f
C604 B.n564 VSUBS 0.006242f
C605 B.n565 VSUBS 0.006242f
C606 B.n566 VSUBS 0.006242f
C607 B.n567 VSUBS 0.006242f
C608 B.n568 VSUBS 0.006242f
C609 B.n569 VSUBS 0.006242f
C610 B.n570 VSUBS 0.006242f
C611 B.n571 VSUBS 0.006242f
C612 B.n572 VSUBS 0.006242f
C613 B.n573 VSUBS 0.006242f
C614 B.n574 VSUBS 0.006242f
C615 B.n575 VSUBS 0.006242f
C616 B.n576 VSUBS 0.006242f
C617 B.n577 VSUBS 0.006242f
C618 B.n578 VSUBS 0.006242f
C619 B.n579 VSUBS 0.006242f
C620 B.n580 VSUBS 0.006242f
C621 B.n581 VSUBS 0.006242f
C622 B.n582 VSUBS 0.006242f
C623 B.n583 VSUBS 0.006242f
C624 B.n584 VSUBS 0.006242f
C625 B.n585 VSUBS 0.006242f
C626 B.n586 VSUBS 0.006242f
C627 B.n587 VSUBS 0.006242f
C628 B.n588 VSUBS 0.006242f
C629 B.n589 VSUBS 0.006242f
C630 B.n590 VSUBS 0.006242f
C631 B.n591 VSUBS 0.006242f
C632 B.n592 VSUBS 0.006242f
C633 B.n593 VSUBS 0.006242f
C634 B.n594 VSUBS 0.006242f
C635 B.n595 VSUBS 0.006242f
C636 B.n596 VSUBS 0.006242f
C637 B.n597 VSUBS 0.006242f
C638 B.n598 VSUBS 0.006242f
C639 B.n599 VSUBS 0.006242f
C640 B.n600 VSUBS 0.006242f
C641 B.n601 VSUBS 0.006242f
C642 B.n602 VSUBS 0.006242f
C643 B.n603 VSUBS 0.006242f
C644 B.n604 VSUBS 0.006242f
C645 B.n605 VSUBS 0.006242f
C646 B.n606 VSUBS 0.006242f
C647 B.n607 VSUBS 0.006242f
C648 B.n608 VSUBS 0.006242f
C649 B.n609 VSUBS 0.006242f
C650 B.n610 VSUBS 0.006242f
C651 B.n611 VSUBS 0.006242f
C652 B.n612 VSUBS 0.006242f
C653 B.n613 VSUBS 0.006242f
C654 B.n614 VSUBS 0.006242f
C655 B.n615 VSUBS 0.006242f
C656 B.n616 VSUBS 0.006242f
C657 B.n617 VSUBS 0.006242f
C658 B.n618 VSUBS 0.006242f
C659 B.n619 VSUBS 0.006242f
C660 B.n620 VSUBS 0.006242f
C661 B.n621 VSUBS 0.006242f
C662 B.n622 VSUBS 0.006242f
C663 B.n623 VSUBS 0.006242f
C664 B.n624 VSUBS 0.006242f
C665 B.n625 VSUBS 0.006242f
C666 B.n626 VSUBS 0.006242f
C667 B.n627 VSUBS 0.006242f
C668 B.n628 VSUBS 0.006242f
C669 B.n629 VSUBS 0.006242f
C670 B.n630 VSUBS 0.006242f
C671 B.n631 VSUBS 0.006242f
C672 B.n632 VSUBS 0.006242f
C673 B.n633 VSUBS 0.006242f
C674 B.n634 VSUBS 0.006242f
C675 B.n635 VSUBS 0.006242f
C676 B.n636 VSUBS 0.006242f
C677 B.n637 VSUBS 0.006242f
C678 B.n638 VSUBS 0.006242f
C679 B.n639 VSUBS 0.006242f
C680 B.n640 VSUBS 0.006242f
C681 B.n641 VSUBS 0.006242f
C682 B.n642 VSUBS 0.006242f
C683 B.n643 VSUBS 0.006242f
C684 B.n644 VSUBS 0.006242f
C685 B.n645 VSUBS 0.006242f
C686 B.n646 VSUBS 0.006242f
C687 B.n647 VSUBS 0.004315f
C688 B.n648 VSUBS 0.014463f
C689 B.n649 VSUBS 0.005049f
C690 B.n650 VSUBS 0.006242f
C691 B.n651 VSUBS 0.006242f
C692 B.n652 VSUBS 0.006242f
C693 B.n653 VSUBS 0.006242f
C694 B.n654 VSUBS 0.006242f
C695 B.n655 VSUBS 0.006242f
C696 B.n656 VSUBS 0.006242f
C697 B.n657 VSUBS 0.006242f
C698 B.n658 VSUBS 0.006242f
C699 B.n659 VSUBS 0.006242f
C700 B.n660 VSUBS 0.006242f
C701 B.n661 VSUBS 0.005049f
C702 B.n662 VSUBS 0.014463f
C703 B.n663 VSUBS 0.004315f
C704 B.n664 VSUBS 0.006242f
C705 B.n665 VSUBS 0.006242f
C706 B.n666 VSUBS 0.006242f
C707 B.n667 VSUBS 0.006242f
C708 B.n668 VSUBS 0.006242f
C709 B.n669 VSUBS 0.006242f
C710 B.n670 VSUBS 0.006242f
C711 B.n671 VSUBS 0.006242f
C712 B.n672 VSUBS 0.006242f
C713 B.n673 VSUBS 0.006242f
C714 B.n674 VSUBS 0.006242f
C715 B.n675 VSUBS 0.006242f
C716 B.n676 VSUBS 0.006242f
C717 B.n677 VSUBS 0.006242f
C718 B.n678 VSUBS 0.006242f
C719 B.n679 VSUBS 0.006242f
C720 B.n680 VSUBS 0.006242f
C721 B.n681 VSUBS 0.006242f
C722 B.n682 VSUBS 0.006242f
C723 B.n683 VSUBS 0.006242f
C724 B.n684 VSUBS 0.006242f
C725 B.n685 VSUBS 0.006242f
C726 B.n686 VSUBS 0.006242f
C727 B.n687 VSUBS 0.006242f
C728 B.n688 VSUBS 0.006242f
C729 B.n689 VSUBS 0.006242f
C730 B.n690 VSUBS 0.006242f
C731 B.n691 VSUBS 0.006242f
C732 B.n692 VSUBS 0.006242f
C733 B.n693 VSUBS 0.006242f
C734 B.n694 VSUBS 0.006242f
C735 B.n695 VSUBS 0.006242f
C736 B.n696 VSUBS 0.006242f
C737 B.n697 VSUBS 0.006242f
C738 B.n698 VSUBS 0.006242f
C739 B.n699 VSUBS 0.006242f
C740 B.n700 VSUBS 0.006242f
C741 B.n701 VSUBS 0.006242f
C742 B.n702 VSUBS 0.006242f
C743 B.n703 VSUBS 0.006242f
C744 B.n704 VSUBS 0.006242f
C745 B.n705 VSUBS 0.006242f
C746 B.n706 VSUBS 0.006242f
C747 B.n707 VSUBS 0.006242f
C748 B.n708 VSUBS 0.006242f
C749 B.n709 VSUBS 0.006242f
C750 B.n710 VSUBS 0.006242f
C751 B.n711 VSUBS 0.006242f
C752 B.n712 VSUBS 0.006242f
C753 B.n713 VSUBS 0.006242f
C754 B.n714 VSUBS 0.006242f
C755 B.n715 VSUBS 0.006242f
C756 B.n716 VSUBS 0.006242f
C757 B.n717 VSUBS 0.006242f
C758 B.n718 VSUBS 0.006242f
C759 B.n719 VSUBS 0.006242f
C760 B.n720 VSUBS 0.006242f
C761 B.n721 VSUBS 0.006242f
C762 B.n722 VSUBS 0.006242f
C763 B.n723 VSUBS 0.006242f
C764 B.n724 VSUBS 0.006242f
C765 B.n725 VSUBS 0.006242f
C766 B.n726 VSUBS 0.006242f
C767 B.n727 VSUBS 0.006242f
C768 B.n728 VSUBS 0.006242f
C769 B.n729 VSUBS 0.006242f
C770 B.n730 VSUBS 0.006242f
C771 B.n731 VSUBS 0.006242f
C772 B.n732 VSUBS 0.006242f
C773 B.n733 VSUBS 0.006242f
C774 B.n734 VSUBS 0.006242f
C775 B.n735 VSUBS 0.006242f
C776 B.n736 VSUBS 0.006242f
C777 B.n737 VSUBS 0.006242f
C778 B.n738 VSUBS 0.006242f
C779 B.n739 VSUBS 0.006242f
C780 B.n740 VSUBS 0.006242f
C781 B.n741 VSUBS 0.006242f
C782 B.n742 VSUBS 0.006242f
C783 B.n743 VSUBS 0.006242f
C784 B.n744 VSUBS 0.006242f
C785 B.n745 VSUBS 0.006242f
C786 B.n746 VSUBS 0.006242f
C787 B.n747 VSUBS 0.006242f
C788 B.n748 VSUBS 0.006242f
C789 B.n749 VSUBS 0.006242f
C790 B.n750 VSUBS 0.006242f
C791 B.n751 VSUBS 0.006242f
C792 B.n752 VSUBS 0.006242f
C793 B.n753 VSUBS 0.006242f
C794 B.n754 VSUBS 0.006242f
C795 B.n755 VSUBS 0.006242f
C796 B.n756 VSUBS 0.006242f
C797 B.n757 VSUBS 0.006242f
C798 B.n758 VSUBS 0.006242f
C799 B.n759 VSUBS 0.015917f
C800 B.n760 VSUBS 0.015917f
C801 B.n761 VSUBS 0.015112f
C802 B.n762 VSUBS 0.006242f
C803 B.n763 VSUBS 0.006242f
C804 B.n764 VSUBS 0.006242f
C805 B.n765 VSUBS 0.006242f
C806 B.n766 VSUBS 0.006242f
C807 B.n767 VSUBS 0.006242f
C808 B.n768 VSUBS 0.006242f
C809 B.n769 VSUBS 0.006242f
C810 B.n770 VSUBS 0.006242f
C811 B.n771 VSUBS 0.006242f
C812 B.n772 VSUBS 0.006242f
C813 B.n773 VSUBS 0.006242f
C814 B.n774 VSUBS 0.006242f
C815 B.n775 VSUBS 0.006242f
C816 B.n776 VSUBS 0.006242f
C817 B.n777 VSUBS 0.006242f
C818 B.n778 VSUBS 0.006242f
C819 B.n779 VSUBS 0.006242f
C820 B.n780 VSUBS 0.006242f
C821 B.n781 VSUBS 0.006242f
C822 B.n782 VSUBS 0.006242f
C823 B.n783 VSUBS 0.006242f
C824 B.n784 VSUBS 0.006242f
C825 B.n785 VSUBS 0.006242f
C826 B.n786 VSUBS 0.006242f
C827 B.n787 VSUBS 0.006242f
C828 B.n788 VSUBS 0.006242f
C829 B.n789 VSUBS 0.006242f
C830 B.n790 VSUBS 0.006242f
C831 B.n791 VSUBS 0.006242f
C832 B.n792 VSUBS 0.006242f
C833 B.n793 VSUBS 0.006242f
C834 B.n794 VSUBS 0.006242f
C835 B.n795 VSUBS 0.006242f
C836 B.n796 VSUBS 0.006242f
C837 B.n797 VSUBS 0.006242f
C838 B.n798 VSUBS 0.006242f
C839 B.n799 VSUBS 0.006242f
C840 B.n800 VSUBS 0.006242f
C841 B.n801 VSUBS 0.006242f
C842 B.n802 VSUBS 0.006242f
C843 B.n803 VSUBS 0.008146f
C844 B.n804 VSUBS 0.008678f
C845 B.n805 VSUBS 0.017256f
C846 VDD2.t1 VSUBS 0.417233f
C847 VDD2.t3 VSUBS 0.417233f
C848 VDD2.n0 VSUBS 4.50176f
C849 VDD2.t2 VSUBS 0.417233f
C850 VDD2.t0 VSUBS 0.417233f
C851 VDD2.n1 VSUBS 3.53261f
C852 VDD2.n2 VSUBS 5.01024f
C853 VN.t2 VSUBS 4.03874f
C854 VN.t0 VSUBS 4.03559f
C855 VN.n0 VSUBS 2.6978f
C856 VN.t3 VSUBS 4.03874f
C857 VN.t1 VSUBS 4.03559f
C858 VN.n1 VSUBS 4.56526f
C859 VDD1.t1 VSUBS 0.417286f
C860 VDD1.t3 VSUBS 0.417286f
C861 VDD1.n0 VSUBS 3.53363f
C862 VDD1.t0 VSUBS 0.417286f
C863 VDD1.t2 VSUBS 0.417286f
C864 VDD1.n1 VSUBS 4.52969f
C865 VTAIL.t1 VSUBS 3.61513f
C866 VTAIL.n0 VSUBS 0.71878f
C867 VTAIL.t5 VSUBS 3.61513f
C868 VTAIL.n1 VSUBS 0.788939f
C869 VTAIL.t3 VSUBS 3.61513f
C870 VTAIL.n2 VSUBS 2.4058f
C871 VTAIL.t0 VSUBS 3.61513f
C872 VTAIL.n3 VSUBS 2.4058f
C873 VTAIL.t7 VSUBS 3.61513f
C874 VTAIL.n4 VSUBS 0.788938f
C875 VTAIL.t4 VSUBS 3.61513f
C876 VTAIL.n5 VSUBS 0.788938f
C877 VTAIL.t2 VSUBS 3.61513f
C878 VTAIL.n6 VSUBS 2.4058f
C879 VTAIL.t6 VSUBS 3.61513f
C880 VTAIL.n7 VSUBS 2.32746f
C881 VP.n0 VSUBS 0.044392f
C882 VP.t1 VSUBS 3.91047f
C883 VP.n1 VSUBS 0.048949f
C884 VP.t0 VSUBS 4.1212f
C885 VP.t2 VSUBS 4.12442f
C886 VP.n2 VSUBS 4.64496f
C887 VP.n3 VSUBS 2.18418f
C888 VP.t3 VSUBS 3.91047f
C889 VP.n4 VSUBS 1.47272f
C890 VP.n5 VSUBS 0.060902f
C891 VP.n6 VSUBS 0.044392f
C892 VP.n7 VSUBS 0.033673f
C893 VP.n8 VSUBS 0.033673f
C894 VP.n9 VSUBS 0.048949f
C895 VP.n10 VSUBS 0.060902f
C896 VP.n11 VSUBS 1.47272f
C897 VP.n12 VSUBS 0.037647f
.ends

