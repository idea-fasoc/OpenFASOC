* NGSPICE file created from diff_pair_sample_0017.ext - technology: sky130A

.subckt diff_pair_sample_0017 VTAIL VN VP B VDD2 VDD1
X0 B.t22 B.t20 B.t21 B.t14 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=0.54
X1 VDD1.t9 VP.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X2 VDD2.t9 VN.t0 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X3 B.t19 B.t17 B.t18 B.t10 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=0.54
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=0.54
X5 VDD2.t8 VN.t1 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=0.54
X6 VDD1.t8 VP.t1 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=0.54
X7 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=0 ps=0 w=10.97 l=0.54
X8 VDD2.t7 VN.t2 VTAIL.t19 B.t1 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X9 VTAIL.t1 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X10 VTAIL.t0 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X11 VDD1.t7 VP.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=0.54
X12 VTAIL.t8 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X13 VTAIL.t4 VN.t5 VDD2.t4 B.t23 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X14 VDD1.t5 VP.t4 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X15 VDD1.t4 VP.t5 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=0.54
X16 VDD2.t3 VN.t6 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=0.54
X17 VDD2.t2 VN.t7 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=0.54
X18 VTAIL.t12 VP.t6 VDD1.t3 B.t23 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X19 VDD1.t2 VP.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=4.2783 ps=22.72 w=10.97 l=0.54
X20 VDD2.t1 VN.t8 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=4.2783 pd=22.72 as=1.81005 ps=11.3 w=10.97 l=0.54
X21 VTAIL.t14 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X22 VTAIL.t15 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
X23 VTAIL.t16 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.81005 pd=11.3 as=1.81005 ps=11.3 w=10.97 l=0.54
R0 B.n95 B.t13 695.102
R1 B.n92 B.t20 695.102
R2 B.n354 B.t17 695.102
R3 B.n351 B.t9 695.102
R4 B.n633 B.n632 585
R5 B.n634 B.n633 585
R6 B.n264 B.n90 585
R7 B.n263 B.n262 585
R8 B.n261 B.n260 585
R9 B.n259 B.n258 585
R10 B.n257 B.n256 585
R11 B.n255 B.n254 585
R12 B.n253 B.n252 585
R13 B.n251 B.n250 585
R14 B.n249 B.n248 585
R15 B.n247 B.n246 585
R16 B.n245 B.n244 585
R17 B.n243 B.n242 585
R18 B.n241 B.n240 585
R19 B.n239 B.n238 585
R20 B.n237 B.n236 585
R21 B.n235 B.n234 585
R22 B.n233 B.n232 585
R23 B.n231 B.n230 585
R24 B.n229 B.n228 585
R25 B.n227 B.n226 585
R26 B.n225 B.n224 585
R27 B.n223 B.n222 585
R28 B.n221 B.n220 585
R29 B.n219 B.n218 585
R30 B.n217 B.n216 585
R31 B.n215 B.n214 585
R32 B.n213 B.n212 585
R33 B.n211 B.n210 585
R34 B.n209 B.n208 585
R35 B.n207 B.n206 585
R36 B.n205 B.n204 585
R37 B.n203 B.n202 585
R38 B.n201 B.n200 585
R39 B.n199 B.n198 585
R40 B.n197 B.n196 585
R41 B.n195 B.n194 585
R42 B.n193 B.n192 585
R43 B.n191 B.n190 585
R44 B.n189 B.n188 585
R45 B.n187 B.n186 585
R46 B.n185 B.n184 585
R47 B.n183 B.n182 585
R48 B.n181 B.n180 585
R49 B.n179 B.n178 585
R50 B.n177 B.n176 585
R51 B.n175 B.n174 585
R52 B.n173 B.n172 585
R53 B.n170 B.n169 585
R54 B.n168 B.n167 585
R55 B.n166 B.n165 585
R56 B.n164 B.n163 585
R57 B.n162 B.n161 585
R58 B.n160 B.n159 585
R59 B.n158 B.n157 585
R60 B.n156 B.n155 585
R61 B.n154 B.n153 585
R62 B.n152 B.n151 585
R63 B.n150 B.n149 585
R64 B.n148 B.n147 585
R65 B.n146 B.n145 585
R66 B.n144 B.n143 585
R67 B.n142 B.n141 585
R68 B.n140 B.n139 585
R69 B.n138 B.n137 585
R70 B.n136 B.n135 585
R71 B.n134 B.n133 585
R72 B.n132 B.n131 585
R73 B.n130 B.n129 585
R74 B.n128 B.n127 585
R75 B.n126 B.n125 585
R76 B.n124 B.n123 585
R77 B.n122 B.n121 585
R78 B.n120 B.n119 585
R79 B.n118 B.n117 585
R80 B.n116 B.n115 585
R81 B.n114 B.n113 585
R82 B.n112 B.n111 585
R83 B.n110 B.n109 585
R84 B.n108 B.n107 585
R85 B.n106 B.n105 585
R86 B.n104 B.n103 585
R87 B.n102 B.n101 585
R88 B.n100 B.n99 585
R89 B.n98 B.n97 585
R90 B.n47 B.n46 585
R91 B.n637 B.n636 585
R92 B.n631 B.n91 585
R93 B.n91 B.n44 585
R94 B.n630 B.n43 585
R95 B.n641 B.n43 585
R96 B.n629 B.n42 585
R97 B.n642 B.n42 585
R98 B.n628 B.n41 585
R99 B.n643 B.n41 585
R100 B.n627 B.n626 585
R101 B.n626 B.n40 585
R102 B.n625 B.n36 585
R103 B.n649 B.n36 585
R104 B.n624 B.n35 585
R105 B.n650 B.n35 585
R106 B.n623 B.n34 585
R107 B.n651 B.n34 585
R108 B.n622 B.n621 585
R109 B.n621 B.n30 585
R110 B.n620 B.n29 585
R111 B.n657 B.n29 585
R112 B.n619 B.n28 585
R113 B.n658 B.n28 585
R114 B.n618 B.n27 585
R115 B.n659 B.n27 585
R116 B.n617 B.n616 585
R117 B.n616 B.n26 585
R118 B.n615 B.n22 585
R119 B.n665 B.n22 585
R120 B.n614 B.n21 585
R121 B.n666 B.n21 585
R122 B.n613 B.n20 585
R123 B.n667 B.n20 585
R124 B.n612 B.n611 585
R125 B.n611 B.n16 585
R126 B.n610 B.n15 585
R127 B.n673 B.n15 585
R128 B.n609 B.n14 585
R129 B.n674 B.n14 585
R130 B.n608 B.n13 585
R131 B.n675 B.n13 585
R132 B.n607 B.n606 585
R133 B.n606 B.n12 585
R134 B.n605 B.n604 585
R135 B.n605 B.n8 585
R136 B.n603 B.n7 585
R137 B.n682 B.n7 585
R138 B.n602 B.n6 585
R139 B.n683 B.n6 585
R140 B.n601 B.n5 585
R141 B.n684 B.n5 585
R142 B.n600 B.n599 585
R143 B.n599 B.n4 585
R144 B.n598 B.n265 585
R145 B.n598 B.n597 585
R146 B.n587 B.n266 585
R147 B.n590 B.n266 585
R148 B.n589 B.n588 585
R149 B.n591 B.n589 585
R150 B.n586 B.n270 585
R151 B.n274 B.n270 585
R152 B.n585 B.n584 585
R153 B.n584 B.n583 585
R154 B.n272 B.n271 585
R155 B.n273 B.n272 585
R156 B.n576 B.n575 585
R157 B.n577 B.n576 585
R158 B.n574 B.n279 585
R159 B.n279 B.n278 585
R160 B.n573 B.n572 585
R161 B.n572 B.n571 585
R162 B.n281 B.n280 585
R163 B.n564 B.n281 585
R164 B.n563 B.n562 585
R165 B.n565 B.n563 585
R166 B.n561 B.n285 585
R167 B.n289 B.n285 585
R168 B.n560 B.n559 585
R169 B.n559 B.n558 585
R170 B.n287 B.n286 585
R171 B.n288 B.n287 585
R172 B.n551 B.n550 585
R173 B.n552 B.n551 585
R174 B.n549 B.n294 585
R175 B.n294 B.n293 585
R176 B.n548 B.n547 585
R177 B.n547 B.n546 585
R178 B.n296 B.n295 585
R179 B.n539 B.n296 585
R180 B.n538 B.n537 585
R181 B.n540 B.n538 585
R182 B.n536 B.n301 585
R183 B.n301 B.n300 585
R184 B.n535 B.n534 585
R185 B.n534 B.n533 585
R186 B.n303 B.n302 585
R187 B.n304 B.n303 585
R188 B.n529 B.n528 585
R189 B.n307 B.n306 585
R190 B.n525 B.n524 585
R191 B.n526 B.n525 585
R192 B.n523 B.n350 585
R193 B.n522 B.n521 585
R194 B.n520 B.n519 585
R195 B.n518 B.n517 585
R196 B.n516 B.n515 585
R197 B.n514 B.n513 585
R198 B.n512 B.n511 585
R199 B.n510 B.n509 585
R200 B.n508 B.n507 585
R201 B.n506 B.n505 585
R202 B.n504 B.n503 585
R203 B.n502 B.n501 585
R204 B.n500 B.n499 585
R205 B.n498 B.n497 585
R206 B.n496 B.n495 585
R207 B.n494 B.n493 585
R208 B.n492 B.n491 585
R209 B.n490 B.n489 585
R210 B.n488 B.n487 585
R211 B.n486 B.n485 585
R212 B.n484 B.n483 585
R213 B.n482 B.n481 585
R214 B.n480 B.n479 585
R215 B.n478 B.n477 585
R216 B.n476 B.n475 585
R217 B.n474 B.n473 585
R218 B.n472 B.n471 585
R219 B.n470 B.n469 585
R220 B.n468 B.n467 585
R221 B.n466 B.n465 585
R222 B.n464 B.n463 585
R223 B.n462 B.n461 585
R224 B.n460 B.n459 585
R225 B.n458 B.n457 585
R226 B.n456 B.n455 585
R227 B.n454 B.n453 585
R228 B.n452 B.n451 585
R229 B.n450 B.n449 585
R230 B.n448 B.n447 585
R231 B.n446 B.n445 585
R232 B.n444 B.n443 585
R233 B.n442 B.n441 585
R234 B.n440 B.n439 585
R235 B.n438 B.n437 585
R236 B.n436 B.n435 585
R237 B.n433 B.n432 585
R238 B.n431 B.n430 585
R239 B.n429 B.n428 585
R240 B.n427 B.n426 585
R241 B.n425 B.n424 585
R242 B.n423 B.n422 585
R243 B.n421 B.n420 585
R244 B.n419 B.n418 585
R245 B.n417 B.n416 585
R246 B.n415 B.n414 585
R247 B.n413 B.n412 585
R248 B.n411 B.n410 585
R249 B.n409 B.n408 585
R250 B.n407 B.n406 585
R251 B.n405 B.n404 585
R252 B.n403 B.n402 585
R253 B.n401 B.n400 585
R254 B.n399 B.n398 585
R255 B.n397 B.n396 585
R256 B.n395 B.n394 585
R257 B.n393 B.n392 585
R258 B.n391 B.n390 585
R259 B.n389 B.n388 585
R260 B.n387 B.n386 585
R261 B.n385 B.n384 585
R262 B.n383 B.n382 585
R263 B.n381 B.n380 585
R264 B.n379 B.n378 585
R265 B.n377 B.n376 585
R266 B.n375 B.n374 585
R267 B.n373 B.n372 585
R268 B.n371 B.n370 585
R269 B.n369 B.n368 585
R270 B.n367 B.n366 585
R271 B.n365 B.n364 585
R272 B.n363 B.n362 585
R273 B.n361 B.n360 585
R274 B.n359 B.n358 585
R275 B.n357 B.n356 585
R276 B.n530 B.n305 585
R277 B.n305 B.n304 585
R278 B.n532 B.n531 585
R279 B.n533 B.n532 585
R280 B.n299 B.n298 585
R281 B.n300 B.n299 585
R282 B.n542 B.n541 585
R283 B.n541 B.n540 585
R284 B.n543 B.n297 585
R285 B.n539 B.n297 585
R286 B.n545 B.n544 585
R287 B.n546 B.n545 585
R288 B.n292 B.n291 585
R289 B.n293 B.n292 585
R290 B.n554 B.n553 585
R291 B.n553 B.n552 585
R292 B.n555 B.n290 585
R293 B.n290 B.n288 585
R294 B.n557 B.n556 585
R295 B.n558 B.n557 585
R296 B.n284 B.n283 585
R297 B.n289 B.n284 585
R298 B.n567 B.n566 585
R299 B.n566 B.n565 585
R300 B.n568 B.n282 585
R301 B.n564 B.n282 585
R302 B.n570 B.n569 585
R303 B.n571 B.n570 585
R304 B.n277 B.n276 585
R305 B.n278 B.n277 585
R306 B.n579 B.n578 585
R307 B.n578 B.n577 585
R308 B.n580 B.n275 585
R309 B.n275 B.n273 585
R310 B.n582 B.n581 585
R311 B.n583 B.n582 585
R312 B.n269 B.n268 585
R313 B.n274 B.n269 585
R314 B.n593 B.n592 585
R315 B.n592 B.n591 585
R316 B.n594 B.n267 585
R317 B.n590 B.n267 585
R318 B.n596 B.n595 585
R319 B.n597 B.n596 585
R320 B.n3 B.n0 585
R321 B.n4 B.n3 585
R322 B.n681 B.n1 585
R323 B.n682 B.n681 585
R324 B.n680 B.n679 585
R325 B.n680 B.n8 585
R326 B.n678 B.n9 585
R327 B.n12 B.n9 585
R328 B.n677 B.n676 585
R329 B.n676 B.n675 585
R330 B.n11 B.n10 585
R331 B.n674 B.n11 585
R332 B.n672 B.n671 585
R333 B.n673 B.n672 585
R334 B.n670 B.n17 585
R335 B.n17 B.n16 585
R336 B.n669 B.n668 585
R337 B.n668 B.n667 585
R338 B.n19 B.n18 585
R339 B.n666 B.n19 585
R340 B.n664 B.n663 585
R341 B.n665 B.n664 585
R342 B.n662 B.n23 585
R343 B.n26 B.n23 585
R344 B.n661 B.n660 585
R345 B.n660 B.n659 585
R346 B.n25 B.n24 585
R347 B.n658 B.n25 585
R348 B.n656 B.n655 585
R349 B.n657 B.n656 585
R350 B.n654 B.n31 585
R351 B.n31 B.n30 585
R352 B.n653 B.n652 585
R353 B.n652 B.n651 585
R354 B.n33 B.n32 585
R355 B.n650 B.n33 585
R356 B.n648 B.n647 585
R357 B.n649 B.n648 585
R358 B.n646 B.n37 585
R359 B.n40 B.n37 585
R360 B.n645 B.n644 585
R361 B.n644 B.n643 585
R362 B.n39 B.n38 585
R363 B.n642 B.n39 585
R364 B.n640 B.n639 585
R365 B.n641 B.n640 585
R366 B.n638 B.n45 585
R367 B.n45 B.n44 585
R368 B.n685 B.n684 585
R369 B.n683 B.n2 585
R370 B.n636 B.n45 473.281
R371 B.n633 B.n91 473.281
R372 B.n356 B.n303 473.281
R373 B.n528 B.n305 473.281
R374 B.n634 B.n89 256.663
R375 B.n634 B.n88 256.663
R376 B.n634 B.n87 256.663
R377 B.n634 B.n86 256.663
R378 B.n634 B.n85 256.663
R379 B.n634 B.n84 256.663
R380 B.n634 B.n83 256.663
R381 B.n634 B.n82 256.663
R382 B.n634 B.n81 256.663
R383 B.n634 B.n80 256.663
R384 B.n634 B.n79 256.663
R385 B.n634 B.n78 256.663
R386 B.n634 B.n77 256.663
R387 B.n634 B.n76 256.663
R388 B.n634 B.n75 256.663
R389 B.n634 B.n74 256.663
R390 B.n634 B.n73 256.663
R391 B.n634 B.n72 256.663
R392 B.n634 B.n71 256.663
R393 B.n634 B.n70 256.663
R394 B.n634 B.n69 256.663
R395 B.n634 B.n68 256.663
R396 B.n634 B.n67 256.663
R397 B.n634 B.n66 256.663
R398 B.n634 B.n65 256.663
R399 B.n634 B.n64 256.663
R400 B.n634 B.n63 256.663
R401 B.n634 B.n62 256.663
R402 B.n634 B.n61 256.663
R403 B.n634 B.n60 256.663
R404 B.n634 B.n59 256.663
R405 B.n634 B.n58 256.663
R406 B.n634 B.n57 256.663
R407 B.n634 B.n56 256.663
R408 B.n634 B.n55 256.663
R409 B.n634 B.n54 256.663
R410 B.n634 B.n53 256.663
R411 B.n634 B.n52 256.663
R412 B.n634 B.n51 256.663
R413 B.n634 B.n50 256.663
R414 B.n634 B.n49 256.663
R415 B.n634 B.n48 256.663
R416 B.n635 B.n634 256.663
R417 B.n527 B.n526 256.663
R418 B.n526 B.n308 256.663
R419 B.n526 B.n309 256.663
R420 B.n526 B.n310 256.663
R421 B.n526 B.n311 256.663
R422 B.n526 B.n312 256.663
R423 B.n526 B.n313 256.663
R424 B.n526 B.n314 256.663
R425 B.n526 B.n315 256.663
R426 B.n526 B.n316 256.663
R427 B.n526 B.n317 256.663
R428 B.n526 B.n318 256.663
R429 B.n526 B.n319 256.663
R430 B.n526 B.n320 256.663
R431 B.n526 B.n321 256.663
R432 B.n526 B.n322 256.663
R433 B.n526 B.n323 256.663
R434 B.n526 B.n324 256.663
R435 B.n526 B.n325 256.663
R436 B.n526 B.n326 256.663
R437 B.n526 B.n327 256.663
R438 B.n526 B.n328 256.663
R439 B.n526 B.n329 256.663
R440 B.n526 B.n330 256.663
R441 B.n526 B.n331 256.663
R442 B.n526 B.n332 256.663
R443 B.n526 B.n333 256.663
R444 B.n526 B.n334 256.663
R445 B.n526 B.n335 256.663
R446 B.n526 B.n336 256.663
R447 B.n526 B.n337 256.663
R448 B.n526 B.n338 256.663
R449 B.n526 B.n339 256.663
R450 B.n526 B.n340 256.663
R451 B.n526 B.n341 256.663
R452 B.n526 B.n342 256.663
R453 B.n526 B.n343 256.663
R454 B.n526 B.n344 256.663
R455 B.n526 B.n345 256.663
R456 B.n526 B.n346 256.663
R457 B.n526 B.n347 256.663
R458 B.n526 B.n348 256.663
R459 B.n526 B.n349 256.663
R460 B.n687 B.n686 256.663
R461 B.n97 B.n47 163.367
R462 B.n101 B.n100 163.367
R463 B.n105 B.n104 163.367
R464 B.n109 B.n108 163.367
R465 B.n113 B.n112 163.367
R466 B.n117 B.n116 163.367
R467 B.n121 B.n120 163.367
R468 B.n125 B.n124 163.367
R469 B.n129 B.n128 163.367
R470 B.n133 B.n132 163.367
R471 B.n137 B.n136 163.367
R472 B.n141 B.n140 163.367
R473 B.n145 B.n144 163.367
R474 B.n149 B.n148 163.367
R475 B.n153 B.n152 163.367
R476 B.n157 B.n156 163.367
R477 B.n161 B.n160 163.367
R478 B.n165 B.n164 163.367
R479 B.n169 B.n168 163.367
R480 B.n174 B.n173 163.367
R481 B.n178 B.n177 163.367
R482 B.n182 B.n181 163.367
R483 B.n186 B.n185 163.367
R484 B.n190 B.n189 163.367
R485 B.n194 B.n193 163.367
R486 B.n198 B.n197 163.367
R487 B.n202 B.n201 163.367
R488 B.n206 B.n205 163.367
R489 B.n210 B.n209 163.367
R490 B.n214 B.n213 163.367
R491 B.n218 B.n217 163.367
R492 B.n222 B.n221 163.367
R493 B.n226 B.n225 163.367
R494 B.n230 B.n229 163.367
R495 B.n234 B.n233 163.367
R496 B.n238 B.n237 163.367
R497 B.n242 B.n241 163.367
R498 B.n246 B.n245 163.367
R499 B.n250 B.n249 163.367
R500 B.n254 B.n253 163.367
R501 B.n258 B.n257 163.367
R502 B.n262 B.n261 163.367
R503 B.n633 B.n90 163.367
R504 B.n534 B.n303 163.367
R505 B.n534 B.n301 163.367
R506 B.n538 B.n301 163.367
R507 B.n538 B.n296 163.367
R508 B.n547 B.n296 163.367
R509 B.n547 B.n294 163.367
R510 B.n551 B.n294 163.367
R511 B.n551 B.n287 163.367
R512 B.n559 B.n287 163.367
R513 B.n559 B.n285 163.367
R514 B.n563 B.n285 163.367
R515 B.n563 B.n281 163.367
R516 B.n572 B.n281 163.367
R517 B.n572 B.n279 163.367
R518 B.n576 B.n279 163.367
R519 B.n576 B.n272 163.367
R520 B.n584 B.n272 163.367
R521 B.n584 B.n270 163.367
R522 B.n589 B.n270 163.367
R523 B.n589 B.n266 163.367
R524 B.n598 B.n266 163.367
R525 B.n599 B.n598 163.367
R526 B.n599 B.n5 163.367
R527 B.n6 B.n5 163.367
R528 B.n7 B.n6 163.367
R529 B.n605 B.n7 163.367
R530 B.n606 B.n605 163.367
R531 B.n606 B.n13 163.367
R532 B.n14 B.n13 163.367
R533 B.n15 B.n14 163.367
R534 B.n611 B.n15 163.367
R535 B.n611 B.n20 163.367
R536 B.n21 B.n20 163.367
R537 B.n22 B.n21 163.367
R538 B.n616 B.n22 163.367
R539 B.n616 B.n27 163.367
R540 B.n28 B.n27 163.367
R541 B.n29 B.n28 163.367
R542 B.n621 B.n29 163.367
R543 B.n621 B.n34 163.367
R544 B.n35 B.n34 163.367
R545 B.n36 B.n35 163.367
R546 B.n626 B.n36 163.367
R547 B.n626 B.n41 163.367
R548 B.n42 B.n41 163.367
R549 B.n43 B.n42 163.367
R550 B.n91 B.n43 163.367
R551 B.n525 B.n307 163.367
R552 B.n525 B.n350 163.367
R553 B.n521 B.n520 163.367
R554 B.n517 B.n516 163.367
R555 B.n513 B.n512 163.367
R556 B.n509 B.n508 163.367
R557 B.n505 B.n504 163.367
R558 B.n501 B.n500 163.367
R559 B.n497 B.n496 163.367
R560 B.n493 B.n492 163.367
R561 B.n489 B.n488 163.367
R562 B.n485 B.n484 163.367
R563 B.n481 B.n480 163.367
R564 B.n477 B.n476 163.367
R565 B.n473 B.n472 163.367
R566 B.n469 B.n468 163.367
R567 B.n465 B.n464 163.367
R568 B.n461 B.n460 163.367
R569 B.n457 B.n456 163.367
R570 B.n453 B.n452 163.367
R571 B.n449 B.n448 163.367
R572 B.n445 B.n444 163.367
R573 B.n441 B.n440 163.367
R574 B.n437 B.n436 163.367
R575 B.n432 B.n431 163.367
R576 B.n428 B.n427 163.367
R577 B.n424 B.n423 163.367
R578 B.n420 B.n419 163.367
R579 B.n416 B.n415 163.367
R580 B.n412 B.n411 163.367
R581 B.n408 B.n407 163.367
R582 B.n404 B.n403 163.367
R583 B.n400 B.n399 163.367
R584 B.n396 B.n395 163.367
R585 B.n392 B.n391 163.367
R586 B.n388 B.n387 163.367
R587 B.n384 B.n383 163.367
R588 B.n380 B.n379 163.367
R589 B.n376 B.n375 163.367
R590 B.n372 B.n371 163.367
R591 B.n368 B.n367 163.367
R592 B.n364 B.n363 163.367
R593 B.n360 B.n359 163.367
R594 B.n532 B.n305 163.367
R595 B.n532 B.n299 163.367
R596 B.n541 B.n299 163.367
R597 B.n541 B.n297 163.367
R598 B.n545 B.n297 163.367
R599 B.n545 B.n292 163.367
R600 B.n553 B.n292 163.367
R601 B.n553 B.n290 163.367
R602 B.n557 B.n290 163.367
R603 B.n557 B.n284 163.367
R604 B.n566 B.n284 163.367
R605 B.n566 B.n282 163.367
R606 B.n570 B.n282 163.367
R607 B.n570 B.n277 163.367
R608 B.n578 B.n277 163.367
R609 B.n578 B.n275 163.367
R610 B.n582 B.n275 163.367
R611 B.n582 B.n269 163.367
R612 B.n592 B.n269 163.367
R613 B.n592 B.n267 163.367
R614 B.n596 B.n267 163.367
R615 B.n596 B.n3 163.367
R616 B.n685 B.n3 163.367
R617 B.n681 B.n2 163.367
R618 B.n681 B.n680 163.367
R619 B.n680 B.n9 163.367
R620 B.n676 B.n9 163.367
R621 B.n676 B.n11 163.367
R622 B.n672 B.n11 163.367
R623 B.n672 B.n17 163.367
R624 B.n668 B.n17 163.367
R625 B.n668 B.n19 163.367
R626 B.n664 B.n19 163.367
R627 B.n664 B.n23 163.367
R628 B.n660 B.n23 163.367
R629 B.n660 B.n25 163.367
R630 B.n656 B.n25 163.367
R631 B.n656 B.n31 163.367
R632 B.n652 B.n31 163.367
R633 B.n652 B.n33 163.367
R634 B.n648 B.n33 163.367
R635 B.n648 B.n37 163.367
R636 B.n644 B.n37 163.367
R637 B.n644 B.n39 163.367
R638 B.n640 B.n39 163.367
R639 B.n640 B.n45 163.367
R640 B.n92 B.t21 86.5615
R641 B.n354 B.t19 86.5615
R642 B.n95 B.t15 86.5478
R643 B.n351 B.t12 86.5478
R644 B.n526 B.n304 81.9334
R645 B.n634 B.n44 81.9334
R646 B.n636 B.n635 71.676
R647 B.n97 B.n48 71.676
R648 B.n101 B.n49 71.676
R649 B.n105 B.n50 71.676
R650 B.n109 B.n51 71.676
R651 B.n113 B.n52 71.676
R652 B.n117 B.n53 71.676
R653 B.n121 B.n54 71.676
R654 B.n125 B.n55 71.676
R655 B.n129 B.n56 71.676
R656 B.n133 B.n57 71.676
R657 B.n137 B.n58 71.676
R658 B.n141 B.n59 71.676
R659 B.n145 B.n60 71.676
R660 B.n149 B.n61 71.676
R661 B.n153 B.n62 71.676
R662 B.n157 B.n63 71.676
R663 B.n161 B.n64 71.676
R664 B.n165 B.n65 71.676
R665 B.n169 B.n66 71.676
R666 B.n174 B.n67 71.676
R667 B.n178 B.n68 71.676
R668 B.n182 B.n69 71.676
R669 B.n186 B.n70 71.676
R670 B.n190 B.n71 71.676
R671 B.n194 B.n72 71.676
R672 B.n198 B.n73 71.676
R673 B.n202 B.n74 71.676
R674 B.n206 B.n75 71.676
R675 B.n210 B.n76 71.676
R676 B.n214 B.n77 71.676
R677 B.n218 B.n78 71.676
R678 B.n222 B.n79 71.676
R679 B.n226 B.n80 71.676
R680 B.n230 B.n81 71.676
R681 B.n234 B.n82 71.676
R682 B.n238 B.n83 71.676
R683 B.n242 B.n84 71.676
R684 B.n246 B.n85 71.676
R685 B.n250 B.n86 71.676
R686 B.n254 B.n87 71.676
R687 B.n258 B.n88 71.676
R688 B.n262 B.n89 71.676
R689 B.n90 B.n89 71.676
R690 B.n261 B.n88 71.676
R691 B.n257 B.n87 71.676
R692 B.n253 B.n86 71.676
R693 B.n249 B.n85 71.676
R694 B.n245 B.n84 71.676
R695 B.n241 B.n83 71.676
R696 B.n237 B.n82 71.676
R697 B.n233 B.n81 71.676
R698 B.n229 B.n80 71.676
R699 B.n225 B.n79 71.676
R700 B.n221 B.n78 71.676
R701 B.n217 B.n77 71.676
R702 B.n213 B.n76 71.676
R703 B.n209 B.n75 71.676
R704 B.n205 B.n74 71.676
R705 B.n201 B.n73 71.676
R706 B.n197 B.n72 71.676
R707 B.n193 B.n71 71.676
R708 B.n189 B.n70 71.676
R709 B.n185 B.n69 71.676
R710 B.n181 B.n68 71.676
R711 B.n177 B.n67 71.676
R712 B.n173 B.n66 71.676
R713 B.n168 B.n65 71.676
R714 B.n164 B.n64 71.676
R715 B.n160 B.n63 71.676
R716 B.n156 B.n62 71.676
R717 B.n152 B.n61 71.676
R718 B.n148 B.n60 71.676
R719 B.n144 B.n59 71.676
R720 B.n140 B.n58 71.676
R721 B.n136 B.n57 71.676
R722 B.n132 B.n56 71.676
R723 B.n128 B.n55 71.676
R724 B.n124 B.n54 71.676
R725 B.n120 B.n53 71.676
R726 B.n116 B.n52 71.676
R727 B.n112 B.n51 71.676
R728 B.n108 B.n50 71.676
R729 B.n104 B.n49 71.676
R730 B.n100 B.n48 71.676
R731 B.n635 B.n47 71.676
R732 B.n528 B.n527 71.676
R733 B.n350 B.n308 71.676
R734 B.n520 B.n309 71.676
R735 B.n516 B.n310 71.676
R736 B.n512 B.n311 71.676
R737 B.n508 B.n312 71.676
R738 B.n504 B.n313 71.676
R739 B.n500 B.n314 71.676
R740 B.n496 B.n315 71.676
R741 B.n492 B.n316 71.676
R742 B.n488 B.n317 71.676
R743 B.n484 B.n318 71.676
R744 B.n480 B.n319 71.676
R745 B.n476 B.n320 71.676
R746 B.n472 B.n321 71.676
R747 B.n468 B.n322 71.676
R748 B.n464 B.n323 71.676
R749 B.n460 B.n324 71.676
R750 B.n456 B.n325 71.676
R751 B.n452 B.n326 71.676
R752 B.n448 B.n327 71.676
R753 B.n444 B.n328 71.676
R754 B.n440 B.n329 71.676
R755 B.n436 B.n330 71.676
R756 B.n431 B.n331 71.676
R757 B.n427 B.n332 71.676
R758 B.n423 B.n333 71.676
R759 B.n419 B.n334 71.676
R760 B.n415 B.n335 71.676
R761 B.n411 B.n336 71.676
R762 B.n407 B.n337 71.676
R763 B.n403 B.n338 71.676
R764 B.n399 B.n339 71.676
R765 B.n395 B.n340 71.676
R766 B.n391 B.n341 71.676
R767 B.n387 B.n342 71.676
R768 B.n383 B.n343 71.676
R769 B.n379 B.n344 71.676
R770 B.n375 B.n345 71.676
R771 B.n371 B.n346 71.676
R772 B.n367 B.n347 71.676
R773 B.n363 B.n348 71.676
R774 B.n359 B.n349 71.676
R775 B.n527 B.n307 71.676
R776 B.n521 B.n308 71.676
R777 B.n517 B.n309 71.676
R778 B.n513 B.n310 71.676
R779 B.n509 B.n311 71.676
R780 B.n505 B.n312 71.676
R781 B.n501 B.n313 71.676
R782 B.n497 B.n314 71.676
R783 B.n493 B.n315 71.676
R784 B.n489 B.n316 71.676
R785 B.n485 B.n317 71.676
R786 B.n481 B.n318 71.676
R787 B.n477 B.n319 71.676
R788 B.n473 B.n320 71.676
R789 B.n469 B.n321 71.676
R790 B.n465 B.n322 71.676
R791 B.n461 B.n323 71.676
R792 B.n457 B.n324 71.676
R793 B.n453 B.n325 71.676
R794 B.n449 B.n326 71.676
R795 B.n445 B.n327 71.676
R796 B.n441 B.n328 71.676
R797 B.n437 B.n329 71.676
R798 B.n432 B.n330 71.676
R799 B.n428 B.n331 71.676
R800 B.n424 B.n332 71.676
R801 B.n420 B.n333 71.676
R802 B.n416 B.n334 71.676
R803 B.n412 B.n335 71.676
R804 B.n408 B.n336 71.676
R805 B.n404 B.n337 71.676
R806 B.n400 B.n338 71.676
R807 B.n396 B.n339 71.676
R808 B.n392 B.n340 71.676
R809 B.n388 B.n341 71.676
R810 B.n384 B.n342 71.676
R811 B.n380 B.n343 71.676
R812 B.n376 B.n344 71.676
R813 B.n372 B.n345 71.676
R814 B.n368 B.n346 71.676
R815 B.n364 B.n347 71.676
R816 B.n360 B.n348 71.676
R817 B.n356 B.n349 71.676
R818 B.n686 B.n685 71.676
R819 B.n686 B.n2 71.676
R820 B.n93 B.t22 69.6888
R821 B.n355 B.t18 69.6888
R822 B.n96 B.t16 69.675
R823 B.n352 B.t11 69.675
R824 B.n171 B.n96 59.5399
R825 B.n94 B.n93 59.5399
R826 B.n434 B.n355 59.5399
R827 B.n353 B.n352 59.5399
R828 B.n533 B.n304 46.0454
R829 B.n533 B.n300 46.0454
R830 B.n540 B.n300 46.0454
R831 B.n540 B.n539 46.0454
R832 B.n546 B.n293 46.0454
R833 B.n552 B.n293 46.0454
R834 B.n552 B.n288 46.0454
R835 B.n558 B.n288 46.0454
R836 B.n558 B.n289 46.0454
R837 B.n565 B.n564 46.0454
R838 B.n571 B.n278 46.0454
R839 B.n577 B.n278 46.0454
R840 B.n583 B.n273 46.0454
R841 B.n583 B.n274 46.0454
R842 B.n591 B.n590 46.0454
R843 B.n597 B.n4 46.0454
R844 B.n684 B.n4 46.0454
R845 B.n684 B.n683 46.0454
R846 B.n683 B.n682 46.0454
R847 B.n682 B.n8 46.0454
R848 B.n675 B.n12 46.0454
R849 B.n674 B.n673 46.0454
R850 B.n673 B.n16 46.0454
R851 B.n667 B.n666 46.0454
R852 B.n666 B.n665 46.0454
R853 B.n659 B.n26 46.0454
R854 B.n658 B.n657 46.0454
R855 B.n657 B.n30 46.0454
R856 B.n651 B.n30 46.0454
R857 B.n651 B.n650 46.0454
R858 B.n650 B.n649 46.0454
R859 B.n643 B.n40 46.0454
R860 B.n643 B.n642 46.0454
R861 B.n642 B.n641 46.0454
R862 B.n641 B.n44 46.0454
R863 B.n564 B.t2 43.3369
R864 B.n591 B.t23 43.3369
R865 B.n675 B.t4 43.3369
R866 B.n26 B.t5 43.3369
R867 B.n530 B.n529 30.7517
R868 B.n357 B.n302 30.7517
R869 B.n632 B.n631 30.7517
R870 B.n638 B.n637 30.7517
R871 B.n539 B.t10 28.44
R872 B.n565 B.t6 28.44
R873 B.n590 B.t0 28.44
R874 B.n12 B.t7 28.44
R875 B.n659 B.t3 28.44
R876 B.n40 B.t14 28.44
R877 B.n577 B.t8 23.023
R878 B.t8 B.n273 23.023
R879 B.t1 B.n16 23.023
R880 B.n667 B.t1 23.023
R881 B B.n687 18.0485
R882 B.n546 B.t10 17.6059
R883 B.n289 B.t6 17.6059
R884 B.n597 B.t0 17.6059
R885 B.t7 B.n8 17.6059
R886 B.t3 B.n658 17.6059
R887 B.n649 B.t14 17.6059
R888 B.n96 B.n95 16.8732
R889 B.n93 B.n92 16.8732
R890 B.n355 B.n354 16.8732
R891 B.n352 B.n351 16.8732
R892 B.n531 B.n530 10.6151
R893 B.n531 B.n298 10.6151
R894 B.n542 B.n298 10.6151
R895 B.n543 B.n542 10.6151
R896 B.n544 B.n543 10.6151
R897 B.n544 B.n291 10.6151
R898 B.n554 B.n291 10.6151
R899 B.n555 B.n554 10.6151
R900 B.n556 B.n555 10.6151
R901 B.n556 B.n283 10.6151
R902 B.n567 B.n283 10.6151
R903 B.n568 B.n567 10.6151
R904 B.n569 B.n568 10.6151
R905 B.n569 B.n276 10.6151
R906 B.n579 B.n276 10.6151
R907 B.n580 B.n579 10.6151
R908 B.n581 B.n580 10.6151
R909 B.n581 B.n268 10.6151
R910 B.n593 B.n268 10.6151
R911 B.n594 B.n593 10.6151
R912 B.n595 B.n594 10.6151
R913 B.n595 B.n0 10.6151
R914 B.n529 B.n306 10.6151
R915 B.n524 B.n306 10.6151
R916 B.n524 B.n523 10.6151
R917 B.n523 B.n522 10.6151
R918 B.n522 B.n519 10.6151
R919 B.n519 B.n518 10.6151
R920 B.n518 B.n515 10.6151
R921 B.n515 B.n514 10.6151
R922 B.n514 B.n511 10.6151
R923 B.n511 B.n510 10.6151
R924 B.n510 B.n507 10.6151
R925 B.n507 B.n506 10.6151
R926 B.n506 B.n503 10.6151
R927 B.n503 B.n502 10.6151
R928 B.n502 B.n499 10.6151
R929 B.n499 B.n498 10.6151
R930 B.n498 B.n495 10.6151
R931 B.n495 B.n494 10.6151
R932 B.n494 B.n491 10.6151
R933 B.n491 B.n490 10.6151
R934 B.n490 B.n487 10.6151
R935 B.n487 B.n486 10.6151
R936 B.n486 B.n483 10.6151
R937 B.n483 B.n482 10.6151
R938 B.n482 B.n479 10.6151
R939 B.n479 B.n478 10.6151
R940 B.n478 B.n475 10.6151
R941 B.n475 B.n474 10.6151
R942 B.n474 B.n471 10.6151
R943 B.n471 B.n470 10.6151
R944 B.n470 B.n467 10.6151
R945 B.n467 B.n466 10.6151
R946 B.n466 B.n463 10.6151
R947 B.n463 B.n462 10.6151
R948 B.n462 B.n459 10.6151
R949 B.n459 B.n458 10.6151
R950 B.n458 B.n455 10.6151
R951 B.n455 B.n454 10.6151
R952 B.n451 B.n450 10.6151
R953 B.n450 B.n447 10.6151
R954 B.n447 B.n446 10.6151
R955 B.n446 B.n443 10.6151
R956 B.n443 B.n442 10.6151
R957 B.n442 B.n439 10.6151
R958 B.n439 B.n438 10.6151
R959 B.n438 B.n435 10.6151
R960 B.n433 B.n430 10.6151
R961 B.n430 B.n429 10.6151
R962 B.n429 B.n426 10.6151
R963 B.n426 B.n425 10.6151
R964 B.n425 B.n422 10.6151
R965 B.n422 B.n421 10.6151
R966 B.n421 B.n418 10.6151
R967 B.n418 B.n417 10.6151
R968 B.n417 B.n414 10.6151
R969 B.n414 B.n413 10.6151
R970 B.n413 B.n410 10.6151
R971 B.n410 B.n409 10.6151
R972 B.n409 B.n406 10.6151
R973 B.n406 B.n405 10.6151
R974 B.n405 B.n402 10.6151
R975 B.n402 B.n401 10.6151
R976 B.n401 B.n398 10.6151
R977 B.n398 B.n397 10.6151
R978 B.n397 B.n394 10.6151
R979 B.n394 B.n393 10.6151
R980 B.n393 B.n390 10.6151
R981 B.n390 B.n389 10.6151
R982 B.n389 B.n386 10.6151
R983 B.n386 B.n385 10.6151
R984 B.n385 B.n382 10.6151
R985 B.n382 B.n381 10.6151
R986 B.n381 B.n378 10.6151
R987 B.n378 B.n377 10.6151
R988 B.n377 B.n374 10.6151
R989 B.n374 B.n373 10.6151
R990 B.n373 B.n370 10.6151
R991 B.n370 B.n369 10.6151
R992 B.n369 B.n366 10.6151
R993 B.n366 B.n365 10.6151
R994 B.n365 B.n362 10.6151
R995 B.n362 B.n361 10.6151
R996 B.n361 B.n358 10.6151
R997 B.n358 B.n357 10.6151
R998 B.n535 B.n302 10.6151
R999 B.n536 B.n535 10.6151
R1000 B.n537 B.n536 10.6151
R1001 B.n537 B.n295 10.6151
R1002 B.n548 B.n295 10.6151
R1003 B.n549 B.n548 10.6151
R1004 B.n550 B.n549 10.6151
R1005 B.n550 B.n286 10.6151
R1006 B.n560 B.n286 10.6151
R1007 B.n561 B.n560 10.6151
R1008 B.n562 B.n561 10.6151
R1009 B.n562 B.n280 10.6151
R1010 B.n573 B.n280 10.6151
R1011 B.n574 B.n573 10.6151
R1012 B.n575 B.n574 10.6151
R1013 B.n575 B.n271 10.6151
R1014 B.n585 B.n271 10.6151
R1015 B.n586 B.n585 10.6151
R1016 B.n588 B.n586 10.6151
R1017 B.n588 B.n587 10.6151
R1018 B.n587 B.n265 10.6151
R1019 B.n600 B.n265 10.6151
R1020 B.n601 B.n600 10.6151
R1021 B.n602 B.n601 10.6151
R1022 B.n603 B.n602 10.6151
R1023 B.n604 B.n603 10.6151
R1024 B.n607 B.n604 10.6151
R1025 B.n608 B.n607 10.6151
R1026 B.n609 B.n608 10.6151
R1027 B.n610 B.n609 10.6151
R1028 B.n612 B.n610 10.6151
R1029 B.n613 B.n612 10.6151
R1030 B.n614 B.n613 10.6151
R1031 B.n615 B.n614 10.6151
R1032 B.n617 B.n615 10.6151
R1033 B.n618 B.n617 10.6151
R1034 B.n619 B.n618 10.6151
R1035 B.n620 B.n619 10.6151
R1036 B.n622 B.n620 10.6151
R1037 B.n623 B.n622 10.6151
R1038 B.n624 B.n623 10.6151
R1039 B.n625 B.n624 10.6151
R1040 B.n627 B.n625 10.6151
R1041 B.n628 B.n627 10.6151
R1042 B.n629 B.n628 10.6151
R1043 B.n630 B.n629 10.6151
R1044 B.n631 B.n630 10.6151
R1045 B.n679 B.n1 10.6151
R1046 B.n679 B.n678 10.6151
R1047 B.n678 B.n677 10.6151
R1048 B.n677 B.n10 10.6151
R1049 B.n671 B.n10 10.6151
R1050 B.n671 B.n670 10.6151
R1051 B.n670 B.n669 10.6151
R1052 B.n669 B.n18 10.6151
R1053 B.n663 B.n18 10.6151
R1054 B.n663 B.n662 10.6151
R1055 B.n662 B.n661 10.6151
R1056 B.n661 B.n24 10.6151
R1057 B.n655 B.n24 10.6151
R1058 B.n655 B.n654 10.6151
R1059 B.n654 B.n653 10.6151
R1060 B.n653 B.n32 10.6151
R1061 B.n647 B.n32 10.6151
R1062 B.n647 B.n646 10.6151
R1063 B.n646 B.n645 10.6151
R1064 B.n645 B.n38 10.6151
R1065 B.n639 B.n38 10.6151
R1066 B.n639 B.n638 10.6151
R1067 B.n637 B.n46 10.6151
R1068 B.n98 B.n46 10.6151
R1069 B.n99 B.n98 10.6151
R1070 B.n102 B.n99 10.6151
R1071 B.n103 B.n102 10.6151
R1072 B.n106 B.n103 10.6151
R1073 B.n107 B.n106 10.6151
R1074 B.n110 B.n107 10.6151
R1075 B.n111 B.n110 10.6151
R1076 B.n114 B.n111 10.6151
R1077 B.n115 B.n114 10.6151
R1078 B.n118 B.n115 10.6151
R1079 B.n119 B.n118 10.6151
R1080 B.n122 B.n119 10.6151
R1081 B.n123 B.n122 10.6151
R1082 B.n126 B.n123 10.6151
R1083 B.n127 B.n126 10.6151
R1084 B.n130 B.n127 10.6151
R1085 B.n131 B.n130 10.6151
R1086 B.n134 B.n131 10.6151
R1087 B.n135 B.n134 10.6151
R1088 B.n138 B.n135 10.6151
R1089 B.n139 B.n138 10.6151
R1090 B.n142 B.n139 10.6151
R1091 B.n143 B.n142 10.6151
R1092 B.n146 B.n143 10.6151
R1093 B.n147 B.n146 10.6151
R1094 B.n150 B.n147 10.6151
R1095 B.n151 B.n150 10.6151
R1096 B.n154 B.n151 10.6151
R1097 B.n155 B.n154 10.6151
R1098 B.n158 B.n155 10.6151
R1099 B.n159 B.n158 10.6151
R1100 B.n162 B.n159 10.6151
R1101 B.n163 B.n162 10.6151
R1102 B.n166 B.n163 10.6151
R1103 B.n167 B.n166 10.6151
R1104 B.n170 B.n167 10.6151
R1105 B.n175 B.n172 10.6151
R1106 B.n176 B.n175 10.6151
R1107 B.n179 B.n176 10.6151
R1108 B.n180 B.n179 10.6151
R1109 B.n183 B.n180 10.6151
R1110 B.n184 B.n183 10.6151
R1111 B.n187 B.n184 10.6151
R1112 B.n188 B.n187 10.6151
R1113 B.n192 B.n191 10.6151
R1114 B.n195 B.n192 10.6151
R1115 B.n196 B.n195 10.6151
R1116 B.n199 B.n196 10.6151
R1117 B.n200 B.n199 10.6151
R1118 B.n203 B.n200 10.6151
R1119 B.n204 B.n203 10.6151
R1120 B.n207 B.n204 10.6151
R1121 B.n208 B.n207 10.6151
R1122 B.n211 B.n208 10.6151
R1123 B.n212 B.n211 10.6151
R1124 B.n215 B.n212 10.6151
R1125 B.n216 B.n215 10.6151
R1126 B.n219 B.n216 10.6151
R1127 B.n220 B.n219 10.6151
R1128 B.n223 B.n220 10.6151
R1129 B.n224 B.n223 10.6151
R1130 B.n227 B.n224 10.6151
R1131 B.n228 B.n227 10.6151
R1132 B.n231 B.n228 10.6151
R1133 B.n232 B.n231 10.6151
R1134 B.n235 B.n232 10.6151
R1135 B.n236 B.n235 10.6151
R1136 B.n239 B.n236 10.6151
R1137 B.n240 B.n239 10.6151
R1138 B.n243 B.n240 10.6151
R1139 B.n244 B.n243 10.6151
R1140 B.n247 B.n244 10.6151
R1141 B.n248 B.n247 10.6151
R1142 B.n251 B.n248 10.6151
R1143 B.n252 B.n251 10.6151
R1144 B.n255 B.n252 10.6151
R1145 B.n256 B.n255 10.6151
R1146 B.n259 B.n256 10.6151
R1147 B.n260 B.n259 10.6151
R1148 B.n263 B.n260 10.6151
R1149 B.n264 B.n263 10.6151
R1150 B.n632 B.n264 10.6151
R1151 B.n687 B.n0 8.11757
R1152 B.n687 B.n1 8.11757
R1153 B.n451 B.n353 6.5566
R1154 B.n435 B.n434 6.5566
R1155 B.n172 B.n171 6.5566
R1156 B.n188 B.n94 6.5566
R1157 B.n454 B.n353 4.05904
R1158 B.n434 B.n433 4.05904
R1159 B.n171 B.n170 4.05904
R1160 B.n191 B.n94 4.05904
R1161 B.n571 B.t2 2.70903
R1162 B.n274 B.t23 2.70903
R1163 B.t4 B.n674 2.70903
R1164 B.n665 B.t5 2.70903
R1165 VP.n5 VP.t5 583.761
R1166 VP.n16 VP.t1 562.78
R1167 VP.n17 VP.t8 562.78
R1168 VP.n1 VP.t4 562.78
R1169 VP.n23 VP.t6 562.78
R1170 VP.n24 VP.t2 562.78
R1171 VP.n13 VP.t7 562.78
R1172 VP.n12 VP.t9 562.78
R1173 VP.n4 VP.t0 562.78
R1174 VP.n6 VP.t3 562.78
R1175 VP.n25 VP.n24 161.3
R1176 VP.n8 VP.n7 161.3
R1177 VP.n9 VP.n4 161.3
R1178 VP.n11 VP.n10 161.3
R1179 VP.n12 VP.n3 161.3
R1180 VP.n14 VP.n13 161.3
R1181 VP.n23 VP.n0 161.3
R1182 VP.n22 VP.n21 161.3
R1183 VP.n20 VP.n1 161.3
R1184 VP.n19 VP.n18 161.3
R1185 VP.n17 VP.n2 161.3
R1186 VP.n16 VP.n15 161.3
R1187 VP.n8 VP.n5 70.4033
R1188 VP.n17 VP.n16 48.2005
R1189 VP.n24 VP.n23 48.2005
R1190 VP.n13 VP.n12 48.2005
R1191 VP.n15 VP.n14 41.2316
R1192 VP.n18 VP.n1 33.5944
R1193 VP.n22 VP.n1 33.5944
R1194 VP.n11 VP.n4 33.5944
R1195 VP.n7 VP.n4 33.5944
R1196 VP.n6 VP.n5 20.9576
R1197 VP.n18 VP.n17 14.6066
R1198 VP.n23 VP.n22 14.6066
R1199 VP.n12 VP.n11 14.6066
R1200 VP.n7 VP.n6 14.6066
R1201 VP.n9 VP.n8 0.189894
R1202 VP.n10 VP.n9 0.189894
R1203 VP.n10 VP.n3 0.189894
R1204 VP.n14 VP.n3 0.189894
R1205 VP.n15 VP.n2 0.189894
R1206 VP.n19 VP.n2 0.189894
R1207 VP.n20 VP.n19 0.189894
R1208 VP.n21 VP.n20 0.189894
R1209 VP.n21 VP.n0 0.189894
R1210 VP.n25 VP.n0 0.189894
R1211 VP VP.n25 0.0516364
R1212 VTAIL.n11 VTAIL.t2 45.9776
R1213 VTAIL.n17 VTAIL.t5 45.9775
R1214 VTAIL.n2 VTAIL.t7 45.9775
R1215 VTAIL.n16 VTAIL.t13 45.9775
R1216 VTAIL.n15 VTAIL.n14 44.1728
R1217 VTAIL.n13 VTAIL.n12 44.1728
R1218 VTAIL.n10 VTAIL.n9 44.1728
R1219 VTAIL.n8 VTAIL.n7 44.1728
R1220 VTAIL.n19 VTAIL.n18 44.1725
R1221 VTAIL.n1 VTAIL.n0 44.1725
R1222 VTAIL.n4 VTAIL.n3 44.1725
R1223 VTAIL.n6 VTAIL.n5 44.1725
R1224 VTAIL.n8 VTAIL.n6 23.3238
R1225 VTAIL.n17 VTAIL.n16 22.5738
R1226 VTAIL.n18 VTAIL.t19 1.80542
R1227 VTAIL.n18 VTAIL.t0 1.80542
R1228 VTAIL.n0 VTAIL.t18 1.80542
R1229 VTAIL.n0 VTAIL.t1 1.80542
R1230 VTAIL.n3 VTAIL.t10 1.80542
R1231 VTAIL.n3 VTAIL.t12 1.80542
R1232 VTAIL.n5 VTAIL.t9 1.80542
R1233 VTAIL.n5 VTAIL.t14 1.80542
R1234 VTAIL.n14 VTAIL.t6 1.80542
R1235 VTAIL.n14 VTAIL.t15 1.80542
R1236 VTAIL.n12 VTAIL.t11 1.80542
R1237 VTAIL.n12 VTAIL.t8 1.80542
R1238 VTAIL.n9 VTAIL.t17 1.80542
R1239 VTAIL.n9 VTAIL.t4 1.80542
R1240 VTAIL.n7 VTAIL.t3 1.80542
R1241 VTAIL.n7 VTAIL.t16 1.80542
R1242 VTAIL.n13 VTAIL.n11 0.845328
R1243 VTAIL.n2 VTAIL.n1 0.845328
R1244 VTAIL.n10 VTAIL.n8 0.7505
R1245 VTAIL.n11 VTAIL.n10 0.7505
R1246 VTAIL.n15 VTAIL.n13 0.7505
R1247 VTAIL.n16 VTAIL.n15 0.7505
R1248 VTAIL.n6 VTAIL.n4 0.7505
R1249 VTAIL.n4 VTAIL.n2 0.7505
R1250 VTAIL.n19 VTAIL.n17 0.7505
R1251 VTAIL VTAIL.n1 0.62119
R1252 VTAIL VTAIL.n19 0.12981
R1253 VDD1.n1 VDD1.t4 63.4064
R1254 VDD1.n3 VDD1.t8 63.4063
R1255 VDD1.n5 VDD1.n4 61.3585
R1256 VDD1.n1 VDD1.n0 60.8516
R1257 VDD1.n7 VDD1.n6 60.8514
R1258 VDD1.n3 VDD1.n2 60.8513
R1259 VDD1.n7 VDD1.n5 37.6927
R1260 VDD1.n6 VDD1.t0 1.80542
R1261 VDD1.n6 VDD1.t2 1.80542
R1262 VDD1.n0 VDD1.t6 1.80542
R1263 VDD1.n0 VDD1.t9 1.80542
R1264 VDD1.n4 VDD1.t3 1.80542
R1265 VDD1.n4 VDD1.t7 1.80542
R1266 VDD1.n2 VDD1.t1 1.80542
R1267 VDD1.n2 VDD1.t5 1.80542
R1268 VDD1 VDD1.n7 0.50481
R1269 VDD1 VDD1.n1 0.24619
R1270 VDD1.n5 VDD1.n3 0.132654
R1271 VN.n2 VN.t1 583.761
R1272 VN.n14 VN.t6 583.761
R1273 VN.n3 VN.t3 562.78
R1274 VN.n1 VN.t2 562.78
R1275 VN.n9 VN.t4 562.78
R1276 VN.n10 VN.t7 562.78
R1277 VN.n15 VN.t5 562.78
R1278 VN.n13 VN.t0 562.78
R1279 VN.n21 VN.t9 562.78
R1280 VN.n22 VN.t8 562.78
R1281 VN.n11 VN.n10 161.3
R1282 VN.n23 VN.n22 161.3
R1283 VN.n21 VN.n12 161.3
R1284 VN.n20 VN.n19 161.3
R1285 VN.n18 VN.n13 161.3
R1286 VN.n17 VN.n16 161.3
R1287 VN.n9 VN.n0 161.3
R1288 VN.n8 VN.n7 161.3
R1289 VN.n6 VN.n1 161.3
R1290 VN.n5 VN.n4 161.3
R1291 VN.n17 VN.n14 70.4033
R1292 VN.n5 VN.n2 70.4033
R1293 VN.n10 VN.n9 48.2005
R1294 VN.n22 VN.n21 48.2005
R1295 VN VN.n23 41.6122
R1296 VN.n4 VN.n1 33.5944
R1297 VN.n8 VN.n1 33.5944
R1298 VN.n16 VN.n13 33.5944
R1299 VN.n20 VN.n13 33.5944
R1300 VN.n15 VN.n14 20.9576
R1301 VN.n3 VN.n2 20.9576
R1302 VN.n4 VN.n3 14.6066
R1303 VN.n9 VN.n8 14.6066
R1304 VN.n16 VN.n15 14.6066
R1305 VN.n21 VN.n20 14.6066
R1306 VN.n23 VN.n12 0.189894
R1307 VN.n19 VN.n12 0.189894
R1308 VN.n19 VN.n18 0.189894
R1309 VN.n18 VN.n17 0.189894
R1310 VN.n6 VN.n5 0.189894
R1311 VN.n7 VN.n6 0.189894
R1312 VN.n7 VN.n0 0.189894
R1313 VN.n11 VN.n0 0.189894
R1314 VN VN.n11 0.0516364
R1315 VDD2.n1 VDD2.t8 63.4063
R1316 VDD2.n4 VDD2.t1 62.6564
R1317 VDD2.n3 VDD2.n2 61.3585
R1318 VDD2 VDD2.n7 61.3557
R1319 VDD2.n6 VDD2.n5 60.8516
R1320 VDD2.n1 VDD2.n0 60.8513
R1321 VDD2.n4 VDD2.n3 36.7347
R1322 VDD2.n7 VDD2.t4 1.80542
R1323 VDD2.n7 VDD2.t3 1.80542
R1324 VDD2.n5 VDD2.t0 1.80542
R1325 VDD2.n5 VDD2.t9 1.80542
R1326 VDD2.n2 VDD2.t5 1.80542
R1327 VDD2.n2 VDD2.t2 1.80542
R1328 VDD2.n0 VDD2.t6 1.80542
R1329 VDD2.n0 VDD2.t7 1.80542
R1330 VDD2.n6 VDD2.n4 0.7505
R1331 VDD2 VDD2.n6 0.24619
R1332 VDD2.n3 VDD2.n1 0.132654
C0 VTAIL VP 5.12228f
C1 VTAIL VDD1 14.799001f
C2 VP VDD1 5.4887f
C3 VTAIL VN 5.10766f
C4 VN VP 5.16802f
C5 VDD2 VTAIL 14.832099f
C6 VDD2 VP 0.321021f
C7 VN VDD1 0.148591f
C8 VDD2 VDD1 0.872221f
C9 VDD2 VN 5.32079f
C10 VDD2 B 4.611769f
C11 VDD1 B 4.51852f
C12 VTAIL B 5.987845f
C13 VN B 8.651791f
C14 VP B 6.655975f
C15 VDD2.t8 B 2.51103f
C16 VDD2.t6 B 0.222317f
C17 VDD2.t7 B 0.222317f
C18 VDD2.n0 B 1.96831f
C19 VDD2.n1 B 0.637941f
C20 VDD2.t5 B 0.222317f
C21 VDD2.t2 B 0.222317f
C22 VDD2.n2 B 1.97102f
C23 VDD2.n3 B 1.80141f
C24 VDD2.t1 B 2.50688f
C25 VDD2.n4 B 2.30538f
C26 VDD2.t0 B 0.222317f
C27 VDD2.t9 B 0.222317f
C28 VDD2.n5 B 1.96832f
C29 VDD2.n6 B 0.294595f
C30 VDD2.t4 B 0.222317f
C31 VDD2.t3 B 0.222317f
C32 VDD2.n7 B 1.97099f
C33 VN.n0 B 0.046606f
C34 VN.t2 B 0.788768f
C35 VN.n1 B 0.326292f
C36 VN.t1 B 0.800364f
C37 VN.n2 B 0.311323f
C38 VN.t3 B 0.788768f
C39 VN.n3 B 0.32543f
C40 VN.n4 B 0.010576f
C41 VN.n5 B 0.154398f
C42 VN.n6 B 0.046606f
C43 VN.n7 B 0.046606f
C44 VN.n8 B 0.010576f
C45 VN.t4 B 0.788768f
C46 VN.n9 B 0.32543f
C47 VN.t7 B 0.788768f
C48 VN.n10 B 0.322556f
C49 VN.n11 B 0.036118f
C50 VN.n12 B 0.046606f
C51 VN.t0 B 0.788768f
C52 VN.n13 B 0.326292f
C53 VN.t6 B 0.800364f
C54 VN.n14 B 0.311323f
C55 VN.t5 B 0.788768f
C56 VN.n15 B 0.32543f
C57 VN.n16 B 0.010576f
C58 VN.n17 B 0.154398f
C59 VN.n18 B 0.046606f
C60 VN.n19 B 0.046606f
C61 VN.n20 B 0.010576f
C62 VN.t9 B 0.788768f
C63 VN.n21 B 0.32543f
C64 VN.t8 B 0.788768f
C65 VN.n22 B 0.322556f
C66 VN.n23 B 1.89572f
C67 VDD1.t4 B 2.52413f
C68 VDD1.t6 B 0.223476f
C69 VDD1.t9 B 0.223476f
C70 VDD1.n0 B 1.97858f
C71 VDD1.n1 B 0.64616f
C72 VDD1.t8 B 2.52412f
C73 VDD1.t1 B 0.223476f
C74 VDD1.t5 B 0.223476f
C75 VDD1.n2 B 1.97857f
C76 VDD1.n3 B 0.641267f
C77 VDD1.t3 B 0.223476f
C78 VDD1.t7 B 0.223476f
C79 VDD1.n4 B 1.9813f
C80 VDD1.n5 B 1.88606f
C81 VDD1.t0 B 0.223476f
C82 VDD1.t2 B 0.223476f
C83 VDD1.n6 B 1.97857f
C84 VDD1.n7 B 2.31113f
C85 VTAIL.t18 B 0.2335f
C86 VTAIL.t1 B 0.2335f
C87 VTAIL.n0 B 1.98506f
C88 VTAIL.n1 B 0.395852f
C89 VTAIL.t7 B 2.52812f
C90 VTAIL.n2 B 0.500842f
C91 VTAIL.t10 B 0.2335f
C92 VTAIL.t12 B 0.2335f
C93 VTAIL.n3 B 1.98506f
C94 VTAIL.n4 B 0.398845f
C95 VTAIL.t9 B 0.2335f
C96 VTAIL.t14 B 0.2335f
C97 VTAIL.n5 B 1.98506f
C98 VTAIL.n6 B 1.65062f
C99 VTAIL.t3 B 0.2335f
C100 VTAIL.t16 B 0.2335f
C101 VTAIL.n7 B 1.98507f
C102 VTAIL.n8 B 1.65061f
C103 VTAIL.t17 B 0.2335f
C104 VTAIL.t4 B 0.2335f
C105 VTAIL.n9 B 1.98507f
C106 VTAIL.n10 B 0.398838f
C107 VTAIL.t2 B 2.52813f
C108 VTAIL.n11 B 0.500824f
C109 VTAIL.t11 B 0.2335f
C110 VTAIL.t8 B 0.2335f
C111 VTAIL.n12 B 1.98507f
C112 VTAIL.n13 B 0.407069f
C113 VTAIL.t6 B 0.2335f
C114 VTAIL.t15 B 0.2335f
C115 VTAIL.n14 B 1.98507f
C116 VTAIL.n15 B 0.398838f
C117 VTAIL.t13 B 2.52812f
C118 VTAIL.n16 B 1.67929f
C119 VTAIL.t5 B 2.52812f
C120 VTAIL.n17 B 1.67929f
C121 VTAIL.t19 B 0.2335f
C122 VTAIL.t0 B 0.2335f
C123 VTAIL.n18 B 1.98506f
C124 VTAIL.n19 B 0.344974f
C125 VP.n0 B 0.047403f
C126 VP.t4 B 0.802249f
C127 VP.n1 B 0.331869f
C128 VP.n2 B 0.047403f
C129 VP.n3 B 0.047403f
C130 VP.t7 B 0.802249f
C131 VP.t9 B 0.802249f
C132 VP.t0 B 0.802249f
C133 VP.n4 B 0.331869f
C134 VP.t5 B 0.814043f
C135 VP.n5 B 0.316644f
C136 VP.t3 B 0.802249f
C137 VP.n6 B 0.330992f
C138 VP.n7 B 0.010757f
C139 VP.n8 B 0.157037f
C140 VP.n9 B 0.047403f
C141 VP.n10 B 0.047403f
C142 VP.n11 B 0.010757f
C143 VP.n12 B 0.330992f
C144 VP.n13 B 0.328069f
C145 VP.n14 B 1.89697f
C146 VP.n15 B 1.9383f
C147 VP.t1 B 0.802249f
C148 VP.n16 B 0.328069f
C149 VP.t8 B 0.802249f
C150 VP.n17 B 0.330992f
C151 VP.n18 B 0.010757f
C152 VP.n19 B 0.047403f
C153 VP.n20 B 0.047403f
C154 VP.n21 B 0.047403f
C155 VP.n22 B 0.010757f
C156 VP.t6 B 0.802249f
C157 VP.n23 B 0.330992f
C158 VP.t2 B 0.802249f
C159 VP.n24 B 0.328069f
C160 VP.n25 B 0.036735f
.ends

