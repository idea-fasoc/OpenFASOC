* NGSPICE file created from diff_pair_sample_0136.ext - technology: sky130A

.subckt diff_pair_sample_0136 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=0 ps=0 w=18.47 l=3.29
X1 VDD2.t5 VN.t0 VTAIL.t10 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=7.2033 ps=37.72 w=18.47 l=3.29
X2 B.t8 B.t6 B.t7 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=0 ps=0 w=18.47 l=3.29
X3 VTAIL.t4 VP.t0 VDD1.t5 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=3.04755 ps=18.8 w=18.47 l=3.29
X4 VDD2.t4 VN.t1 VTAIL.t6 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=7.2033 ps=37.72 w=18.47 l=3.29
X5 B.t5 B.t3 B.t4 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=0 ps=0 w=18.47 l=3.29
X6 VTAIL.t8 VN.t2 VDD2.t3 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=3.04755 ps=18.8 w=18.47 l=3.29
X7 VTAIL.t7 VN.t3 VDD2.t2 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=3.04755 ps=18.8 w=18.47 l=3.29
X8 VDD1.t4 VP.t1 VTAIL.t2 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=3.04755 ps=18.8 w=18.47 l=3.29
X9 VDD1.t3 VP.t2 VTAIL.t3 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=3.04755 ps=18.8 w=18.47 l=3.29
X10 B.t2 B.t0 B.t1 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=0 ps=0 w=18.47 l=3.29
X11 VDD2.t1 VN.t4 VTAIL.t9 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=3.04755 ps=18.8 w=18.47 l=3.29
X12 VDD1.t2 VP.t3 VTAIL.t1 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=7.2033 ps=37.72 w=18.47 l=3.29
X13 VDD1.t1 VP.t4 VTAIL.t5 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=7.2033 ps=37.72 w=18.47 l=3.29
X14 VDD2.t0 VN.t5 VTAIL.t11 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=7.2033 pd=37.72 as=3.04755 ps=18.8 w=18.47 l=3.29
X15 VTAIL.t0 VP.t5 VDD1.t0 w_n3866_n4662# sky130_fd_pr__pfet_01v8 ad=3.04755 pd=18.8 as=3.04755 ps=18.8 w=18.47 l=3.29
R0 B.n513 B.n148 585
R1 B.n512 B.n511 585
R2 B.n510 B.n149 585
R3 B.n509 B.n508 585
R4 B.n507 B.n150 585
R5 B.n506 B.n505 585
R6 B.n504 B.n151 585
R7 B.n503 B.n502 585
R8 B.n501 B.n152 585
R9 B.n500 B.n499 585
R10 B.n498 B.n153 585
R11 B.n497 B.n496 585
R12 B.n495 B.n154 585
R13 B.n494 B.n493 585
R14 B.n492 B.n155 585
R15 B.n491 B.n490 585
R16 B.n489 B.n156 585
R17 B.n488 B.n487 585
R18 B.n486 B.n157 585
R19 B.n485 B.n484 585
R20 B.n483 B.n158 585
R21 B.n482 B.n481 585
R22 B.n480 B.n159 585
R23 B.n479 B.n478 585
R24 B.n477 B.n160 585
R25 B.n476 B.n475 585
R26 B.n474 B.n161 585
R27 B.n473 B.n472 585
R28 B.n471 B.n162 585
R29 B.n470 B.n469 585
R30 B.n468 B.n163 585
R31 B.n467 B.n466 585
R32 B.n465 B.n164 585
R33 B.n464 B.n463 585
R34 B.n462 B.n165 585
R35 B.n461 B.n460 585
R36 B.n459 B.n166 585
R37 B.n458 B.n457 585
R38 B.n456 B.n167 585
R39 B.n455 B.n454 585
R40 B.n453 B.n168 585
R41 B.n452 B.n451 585
R42 B.n450 B.n169 585
R43 B.n449 B.n448 585
R44 B.n447 B.n170 585
R45 B.n446 B.n445 585
R46 B.n444 B.n171 585
R47 B.n443 B.n442 585
R48 B.n441 B.n172 585
R49 B.n440 B.n439 585
R50 B.n438 B.n173 585
R51 B.n437 B.n436 585
R52 B.n435 B.n174 585
R53 B.n434 B.n433 585
R54 B.n432 B.n175 585
R55 B.n431 B.n430 585
R56 B.n429 B.n176 585
R57 B.n428 B.n427 585
R58 B.n426 B.n177 585
R59 B.n425 B.n424 585
R60 B.n423 B.n178 585
R61 B.n422 B.n421 585
R62 B.n417 B.n179 585
R63 B.n416 B.n415 585
R64 B.n414 B.n180 585
R65 B.n413 B.n412 585
R66 B.n411 B.n181 585
R67 B.n410 B.n409 585
R68 B.n408 B.n182 585
R69 B.n407 B.n406 585
R70 B.n404 B.n183 585
R71 B.n403 B.n402 585
R72 B.n401 B.n186 585
R73 B.n400 B.n399 585
R74 B.n398 B.n187 585
R75 B.n397 B.n396 585
R76 B.n395 B.n188 585
R77 B.n394 B.n393 585
R78 B.n392 B.n189 585
R79 B.n391 B.n390 585
R80 B.n389 B.n190 585
R81 B.n388 B.n387 585
R82 B.n386 B.n191 585
R83 B.n385 B.n384 585
R84 B.n383 B.n192 585
R85 B.n382 B.n381 585
R86 B.n380 B.n193 585
R87 B.n379 B.n378 585
R88 B.n377 B.n194 585
R89 B.n376 B.n375 585
R90 B.n374 B.n195 585
R91 B.n373 B.n372 585
R92 B.n371 B.n196 585
R93 B.n370 B.n369 585
R94 B.n368 B.n197 585
R95 B.n367 B.n366 585
R96 B.n365 B.n198 585
R97 B.n364 B.n363 585
R98 B.n362 B.n199 585
R99 B.n361 B.n360 585
R100 B.n359 B.n200 585
R101 B.n358 B.n357 585
R102 B.n356 B.n201 585
R103 B.n355 B.n354 585
R104 B.n353 B.n202 585
R105 B.n352 B.n351 585
R106 B.n350 B.n203 585
R107 B.n349 B.n348 585
R108 B.n347 B.n204 585
R109 B.n346 B.n345 585
R110 B.n344 B.n205 585
R111 B.n343 B.n342 585
R112 B.n341 B.n206 585
R113 B.n340 B.n339 585
R114 B.n338 B.n207 585
R115 B.n337 B.n336 585
R116 B.n335 B.n208 585
R117 B.n334 B.n333 585
R118 B.n332 B.n209 585
R119 B.n331 B.n330 585
R120 B.n329 B.n210 585
R121 B.n328 B.n327 585
R122 B.n326 B.n211 585
R123 B.n325 B.n324 585
R124 B.n323 B.n212 585
R125 B.n322 B.n321 585
R126 B.n320 B.n213 585
R127 B.n319 B.n318 585
R128 B.n317 B.n214 585
R129 B.n316 B.n315 585
R130 B.n314 B.n215 585
R131 B.n515 B.n514 585
R132 B.n516 B.n147 585
R133 B.n518 B.n517 585
R134 B.n519 B.n146 585
R135 B.n521 B.n520 585
R136 B.n522 B.n145 585
R137 B.n524 B.n523 585
R138 B.n525 B.n144 585
R139 B.n527 B.n526 585
R140 B.n528 B.n143 585
R141 B.n530 B.n529 585
R142 B.n531 B.n142 585
R143 B.n533 B.n532 585
R144 B.n534 B.n141 585
R145 B.n536 B.n535 585
R146 B.n537 B.n140 585
R147 B.n539 B.n538 585
R148 B.n540 B.n139 585
R149 B.n542 B.n541 585
R150 B.n543 B.n138 585
R151 B.n545 B.n544 585
R152 B.n546 B.n137 585
R153 B.n548 B.n547 585
R154 B.n549 B.n136 585
R155 B.n551 B.n550 585
R156 B.n552 B.n135 585
R157 B.n554 B.n553 585
R158 B.n555 B.n134 585
R159 B.n557 B.n556 585
R160 B.n558 B.n133 585
R161 B.n560 B.n559 585
R162 B.n561 B.n132 585
R163 B.n563 B.n562 585
R164 B.n564 B.n131 585
R165 B.n566 B.n565 585
R166 B.n567 B.n130 585
R167 B.n569 B.n568 585
R168 B.n570 B.n129 585
R169 B.n572 B.n571 585
R170 B.n573 B.n128 585
R171 B.n575 B.n574 585
R172 B.n576 B.n127 585
R173 B.n578 B.n577 585
R174 B.n579 B.n126 585
R175 B.n581 B.n580 585
R176 B.n582 B.n125 585
R177 B.n584 B.n583 585
R178 B.n585 B.n124 585
R179 B.n587 B.n586 585
R180 B.n588 B.n123 585
R181 B.n590 B.n589 585
R182 B.n591 B.n122 585
R183 B.n593 B.n592 585
R184 B.n594 B.n121 585
R185 B.n596 B.n595 585
R186 B.n597 B.n120 585
R187 B.n599 B.n598 585
R188 B.n600 B.n119 585
R189 B.n602 B.n601 585
R190 B.n603 B.n118 585
R191 B.n605 B.n604 585
R192 B.n606 B.n117 585
R193 B.n608 B.n607 585
R194 B.n609 B.n116 585
R195 B.n611 B.n610 585
R196 B.n612 B.n115 585
R197 B.n614 B.n613 585
R198 B.n615 B.n114 585
R199 B.n617 B.n616 585
R200 B.n618 B.n113 585
R201 B.n620 B.n619 585
R202 B.n621 B.n112 585
R203 B.n623 B.n622 585
R204 B.n624 B.n111 585
R205 B.n626 B.n625 585
R206 B.n627 B.n110 585
R207 B.n629 B.n628 585
R208 B.n630 B.n109 585
R209 B.n632 B.n631 585
R210 B.n633 B.n108 585
R211 B.n635 B.n634 585
R212 B.n636 B.n107 585
R213 B.n638 B.n637 585
R214 B.n639 B.n106 585
R215 B.n641 B.n640 585
R216 B.n642 B.n105 585
R217 B.n644 B.n643 585
R218 B.n645 B.n104 585
R219 B.n647 B.n646 585
R220 B.n648 B.n103 585
R221 B.n650 B.n649 585
R222 B.n651 B.n102 585
R223 B.n653 B.n652 585
R224 B.n654 B.n101 585
R225 B.n656 B.n655 585
R226 B.n657 B.n100 585
R227 B.n659 B.n658 585
R228 B.n660 B.n99 585
R229 B.n662 B.n661 585
R230 B.n663 B.n98 585
R231 B.n665 B.n664 585
R232 B.n666 B.n97 585
R233 B.n864 B.n27 585
R234 B.n863 B.n862 585
R235 B.n861 B.n28 585
R236 B.n860 B.n859 585
R237 B.n858 B.n29 585
R238 B.n857 B.n856 585
R239 B.n855 B.n30 585
R240 B.n854 B.n853 585
R241 B.n852 B.n31 585
R242 B.n851 B.n850 585
R243 B.n849 B.n32 585
R244 B.n848 B.n847 585
R245 B.n846 B.n33 585
R246 B.n845 B.n844 585
R247 B.n843 B.n34 585
R248 B.n842 B.n841 585
R249 B.n840 B.n35 585
R250 B.n839 B.n838 585
R251 B.n837 B.n36 585
R252 B.n836 B.n835 585
R253 B.n834 B.n37 585
R254 B.n833 B.n832 585
R255 B.n831 B.n38 585
R256 B.n830 B.n829 585
R257 B.n828 B.n39 585
R258 B.n827 B.n826 585
R259 B.n825 B.n40 585
R260 B.n824 B.n823 585
R261 B.n822 B.n41 585
R262 B.n821 B.n820 585
R263 B.n819 B.n42 585
R264 B.n818 B.n817 585
R265 B.n816 B.n43 585
R266 B.n815 B.n814 585
R267 B.n813 B.n44 585
R268 B.n812 B.n811 585
R269 B.n810 B.n45 585
R270 B.n809 B.n808 585
R271 B.n807 B.n46 585
R272 B.n806 B.n805 585
R273 B.n804 B.n47 585
R274 B.n803 B.n802 585
R275 B.n801 B.n48 585
R276 B.n800 B.n799 585
R277 B.n798 B.n49 585
R278 B.n797 B.n796 585
R279 B.n795 B.n50 585
R280 B.n794 B.n793 585
R281 B.n792 B.n51 585
R282 B.n791 B.n790 585
R283 B.n789 B.n52 585
R284 B.n788 B.n787 585
R285 B.n786 B.n53 585
R286 B.n785 B.n784 585
R287 B.n783 B.n54 585
R288 B.n782 B.n781 585
R289 B.n780 B.n55 585
R290 B.n779 B.n778 585
R291 B.n777 B.n56 585
R292 B.n776 B.n775 585
R293 B.n774 B.n57 585
R294 B.n772 B.n771 585
R295 B.n770 B.n60 585
R296 B.n769 B.n768 585
R297 B.n767 B.n61 585
R298 B.n766 B.n765 585
R299 B.n764 B.n62 585
R300 B.n763 B.n762 585
R301 B.n761 B.n63 585
R302 B.n760 B.n759 585
R303 B.n758 B.n757 585
R304 B.n756 B.n67 585
R305 B.n755 B.n754 585
R306 B.n753 B.n68 585
R307 B.n752 B.n751 585
R308 B.n750 B.n69 585
R309 B.n749 B.n748 585
R310 B.n747 B.n70 585
R311 B.n746 B.n745 585
R312 B.n744 B.n71 585
R313 B.n743 B.n742 585
R314 B.n741 B.n72 585
R315 B.n740 B.n739 585
R316 B.n738 B.n73 585
R317 B.n737 B.n736 585
R318 B.n735 B.n74 585
R319 B.n734 B.n733 585
R320 B.n732 B.n75 585
R321 B.n731 B.n730 585
R322 B.n729 B.n76 585
R323 B.n728 B.n727 585
R324 B.n726 B.n77 585
R325 B.n725 B.n724 585
R326 B.n723 B.n78 585
R327 B.n722 B.n721 585
R328 B.n720 B.n79 585
R329 B.n719 B.n718 585
R330 B.n717 B.n80 585
R331 B.n716 B.n715 585
R332 B.n714 B.n81 585
R333 B.n713 B.n712 585
R334 B.n711 B.n82 585
R335 B.n710 B.n709 585
R336 B.n708 B.n83 585
R337 B.n707 B.n706 585
R338 B.n705 B.n84 585
R339 B.n704 B.n703 585
R340 B.n702 B.n85 585
R341 B.n701 B.n700 585
R342 B.n699 B.n86 585
R343 B.n698 B.n697 585
R344 B.n696 B.n87 585
R345 B.n695 B.n694 585
R346 B.n693 B.n88 585
R347 B.n692 B.n691 585
R348 B.n690 B.n89 585
R349 B.n689 B.n688 585
R350 B.n687 B.n90 585
R351 B.n686 B.n685 585
R352 B.n684 B.n91 585
R353 B.n683 B.n682 585
R354 B.n681 B.n92 585
R355 B.n680 B.n679 585
R356 B.n678 B.n93 585
R357 B.n677 B.n676 585
R358 B.n675 B.n94 585
R359 B.n674 B.n673 585
R360 B.n672 B.n95 585
R361 B.n671 B.n670 585
R362 B.n669 B.n96 585
R363 B.n668 B.n667 585
R364 B.n866 B.n865 585
R365 B.n867 B.n26 585
R366 B.n869 B.n868 585
R367 B.n870 B.n25 585
R368 B.n872 B.n871 585
R369 B.n873 B.n24 585
R370 B.n875 B.n874 585
R371 B.n876 B.n23 585
R372 B.n878 B.n877 585
R373 B.n879 B.n22 585
R374 B.n881 B.n880 585
R375 B.n882 B.n21 585
R376 B.n884 B.n883 585
R377 B.n885 B.n20 585
R378 B.n887 B.n886 585
R379 B.n888 B.n19 585
R380 B.n890 B.n889 585
R381 B.n891 B.n18 585
R382 B.n893 B.n892 585
R383 B.n894 B.n17 585
R384 B.n896 B.n895 585
R385 B.n897 B.n16 585
R386 B.n899 B.n898 585
R387 B.n900 B.n15 585
R388 B.n902 B.n901 585
R389 B.n903 B.n14 585
R390 B.n905 B.n904 585
R391 B.n906 B.n13 585
R392 B.n908 B.n907 585
R393 B.n909 B.n12 585
R394 B.n911 B.n910 585
R395 B.n912 B.n11 585
R396 B.n914 B.n913 585
R397 B.n915 B.n10 585
R398 B.n917 B.n916 585
R399 B.n918 B.n9 585
R400 B.n920 B.n919 585
R401 B.n921 B.n8 585
R402 B.n923 B.n922 585
R403 B.n924 B.n7 585
R404 B.n926 B.n925 585
R405 B.n927 B.n6 585
R406 B.n929 B.n928 585
R407 B.n930 B.n5 585
R408 B.n932 B.n931 585
R409 B.n933 B.n4 585
R410 B.n935 B.n934 585
R411 B.n936 B.n3 585
R412 B.n938 B.n937 585
R413 B.n939 B.n0 585
R414 B.n2 B.n1 585
R415 B.n241 B.n240 585
R416 B.n242 B.n239 585
R417 B.n244 B.n243 585
R418 B.n245 B.n238 585
R419 B.n247 B.n246 585
R420 B.n248 B.n237 585
R421 B.n250 B.n249 585
R422 B.n251 B.n236 585
R423 B.n253 B.n252 585
R424 B.n254 B.n235 585
R425 B.n256 B.n255 585
R426 B.n257 B.n234 585
R427 B.n259 B.n258 585
R428 B.n260 B.n233 585
R429 B.n262 B.n261 585
R430 B.n263 B.n232 585
R431 B.n265 B.n264 585
R432 B.n266 B.n231 585
R433 B.n268 B.n267 585
R434 B.n269 B.n230 585
R435 B.n271 B.n270 585
R436 B.n272 B.n229 585
R437 B.n274 B.n273 585
R438 B.n275 B.n228 585
R439 B.n277 B.n276 585
R440 B.n278 B.n227 585
R441 B.n280 B.n279 585
R442 B.n281 B.n226 585
R443 B.n283 B.n282 585
R444 B.n284 B.n225 585
R445 B.n286 B.n285 585
R446 B.n287 B.n224 585
R447 B.n289 B.n288 585
R448 B.n290 B.n223 585
R449 B.n292 B.n291 585
R450 B.n293 B.n222 585
R451 B.n295 B.n294 585
R452 B.n296 B.n221 585
R453 B.n298 B.n297 585
R454 B.n299 B.n220 585
R455 B.n301 B.n300 585
R456 B.n302 B.n219 585
R457 B.n304 B.n303 585
R458 B.n305 B.n218 585
R459 B.n307 B.n306 585
R460 B.n308 B.n217 585
R461 B.n310 B.n309 585
R462 B.n311 B.n216 585
R463 B.n313 B.n312 585
R464 B.n312 B.n215 521.33
R465 B.n514 B.n513 521.33
R466 B.n668 B.n97 521.33
R467 B.n866 B.n27 521.33
R468 B.n184 B.t9 344.192
R469 B.n418 B.t0 344.192
R470 B.n64 B.t3 344.192
R471 B.n58 B.t6 344.192
R472 B.n941 B.n940 256.663
R473 B.n940 B.n939 235.042
R474 B.n940 B.n2 235.042
R475 B.n418 B.t1 178.499
R476 B.n64 B.t5 178.499
R477 B.n184 B.t10 178.475
R478 B.n58 B.t8 178.475
R479 B.n316 B.n215 163.367
R480 B.n317 B.n316 163.367
R481 B.n318 B.n317 163.367
R482 B.n318 B.n213 163.367
R483 B.n322 B.n213 163.367
R484 B.n323 B.n322 163.367
R485 B.n324 B.n323 163.367
R486 B.n324 B.n211 163.367
R487 B.n328 B.n211 163.367
R488 B.n329 B.n328 163.367
R489 B.n330 B.n329 163.367
R490 B.n330 B.n209 163.367
R491 B.n334 B.n209 163.367
R492 B.n335 B.n334 163.367
R493 B.n336 B.n335 163.367
R494 B.n336 B.n207 163.367
R495 B.n340 B.n207 163.367
R496 B.n341 B.n340 163.367
R497 B.n342 B.n341 163.367
R498 B.n342 B.n205 163.367
R499 B.n346 B.n205 163.367
R500 B.n347 B.n346 163.367
R501 B.n348 B.n347 163.367
R502 B.n348 B.n203 163.367
R503 B.n352 B.n203 163.367
R504 B.n353 B.n352 163.367
R505 B.n354 B.n353 163.367
R506 B.n354 B.n201 163.367
R507 B.n358 B.n201 163.367
R508 B.n359 B.n358 163.367
R509 B.n360 B.n359 163.367
R510 B.n360 B.n199 163.367
R511 B.n364 B.n199 163.367
R512 B.n365 B.n364 163.367
R513 B.n366 B.n365 163.367
R514 B.n366 B.n197 163.367
R515 B.n370 B.n197 163.367
R516 B.n371 B.n370 163.367
R517 B.n372 B.n371 163.367
R518 B.n372 B.n195 163.367
R519 B.n376 B.n195 163.367
R520 B.n377 B.n376 163.367
R521 B.n378 B.n377 163.367
R522 B.n378 B.n193 163.367
R523 B.n382 B.n193 163.367
R524 B.n383 B.n382 163.367
R525 B.n384 B.n383 163.367
R526 B.n384 B.n191 163.367
R527 B.n388 B.n191 163.367
R528 B.n389 B.n388 163.367
R529 B.n390 B.n389 163.367
R530 B.n390 B.n189 163.367
R531 B.n394 B.n189 163.367
R532 B.n395 B.n394 163.367
R533 B.n396 B.n395 163.367
R534 B.n396 B.n187 163.367
R535 B.n400 B.n187 163.367
R536 B.n401 B.n400 163.367
R537 B.n402 B.n401 163.367
R538 B.n402 B.n183 163.367
R539 B.n407 B.n183 163.367
R540 B.n408 B.n407 163.367
R541 B.n409 B.n408 163.367
R542 B.n409 B.n181 163.367
R543 B.n413 B.n181 163.367
R544 B.n414 B.n413 163.367
R545 B.n415 B.n414 163.367
R546 B.n415 B.n179 163.367
R547 B.n422 B.n179 163.367
R548 B.n423 B.n422 163.367
R549 B.n424 B.n423 163.367
R550 B.n424 B.n177 163.367
R551 B.n428 B.n177 163.367
R552 B.n429 B.n428 163.367
R553 B.n430 B.n429 163.367
R554 B.n430 B.n175 163.367
R555 B.n434 B.n175 163.367
R556 B.n435 B.n434 163.367
R557 B.n436 B.n435 163.367
R558 B.n436 B.n173 163.367
R559 B.n440 B.n173 163.367
R560 B.n441 B.n440 163.367
R561 B.n442 B.n441 163.367
R562 B.n442 B.n171 163.367
R563 B.n446 B.n171 163.367
R564 B.n447 B.n446 163.367
R565 B.n448 B.n447 163.367
R566 B.n448 B.n169 163.367
R567 B.n452 B.n169 163.367
R568 B.n453 B.n452 163.367
R569 B.n454 B.n453 163.367
R570 B.n454 B.n167 163.367
R571 B.n458 B.n167 163.367
R572 B.n459 B.n458 163.367
R573 B.n460 B.n459 163.367
R574 B.n460 B.n165 163.367
R575 B.n464 B.n165 163.367
R576 B.n465 B.n464 163.367
R577 B.n466 B.n465 163.367
R578 B.n466 B.n163 163.367
R579 B.n470 B.n163 163.367
R580 B.n471 B.n470 163.367
R581 B.n472 B.n471 163.367
R582 B.n472 B.n161 163.367
R583 B.n476 B.n161 163.367
R584 B.n477 B.n476 163.367
R585 B.n478 B.n477 163.367
R586 B.n478 B.n159 163.367
R587 B.n482 B.n159 163.367
R588 B.n483 B.n482 163.367
R589 B.n484 B.n483 163.367
R590 B.n484 B.n157 163.367
R591 B.n488 B.n157 163.367
R592 B.n489 B.n488 163.367
R593 B.n490 B.n489 163.367
R594 B.n490 B.n155 163.367
R595 B.n494 B.n155 163.367
R596 B.n495 B.n494 163.367
R597 B.n496 B.n495 163.367
R598 B.n496 B.n153 163.367
R599 B.n500 B.n153 163.367
R600 B.n501 B.n500 163.367
R601 B.n502 B.n501 163.367
R602 B.n502 B.n151 163.367
R603 B.n506 B.n151 163.367
R604 B.n507 B.n506 163.367
R605 B.n508 B.n507 163.367
R606 B.n508 B.n149 163.367
R607 B.n512 B.n149 163.367
R608 B.n513 B.n512 163.367
R609 B.n664 B.n97 163.367
R610 B.n664 B.n663 163.367
R611 B.n663 B.n662 163.367
R612 B.n662 B.n99 163.367
R613 B.n658 B.n99 163.367
R614 B.n658 B.n657 163.367
R615 B.n657 B.n656 163.367
R616 B.n656 B.n101 163.367
R617 B.n652 B.n101 163.367
R618 B.n652 B.n651 163.367
R619 B.n651 B.n650 163.367
R620 B.n650 B.n103 163.367
R621 B.n646 B.n103 163.367
R622 B.n646 B.n645 163.367
R623 B.n645 B.n644 163.367
R624 B.n644 B.n105 163.367
R625 B.n640 B.n105 163.367
R626 B.n640 B.n639 163.367
R627 B.n639 B.n638 163.367
R628 B.n638 B.n107 163.367
R629 B.n634 B.n107 163.367
R630 B.n634 B.n633 163.367
R631 B.n633 B.n632 163.367
R632 B.n632 B.n109 163.367
R633 B.n628 B.n109 163.367
R634 B.n628 B.n627 163.367
R635 B.n627 B.n626 163.367
R636 B.n626 B.n111 163.367
R637 B.n622 B.n111 163.367
R638 B.n622 B.n621 163.367
R639 B.n621 B.n620 163.367
R640 B.n620 B.n113 163.367
R641 B.n616 B.n113 163.367
R642 B.n616 B.n615 163.367
R643 B.n615 B.n614 163.367
R644 B.n614 B.n115 163.367
R645 B.n610 B.n115 163.367
R646 B.n610 B.n609 163.367
R647 B.n609 B.n608 163.367
R648 B.n608 B.n117 163.367
R649 B.n604 B.n117 163.367
R650 B.n604 B.n603 163.367
R651 B.n603 B.n602 163.367
R652 B.n602 B.n119 163.367
R653 B.n598 B.n119 163.367
R654 B.n598 B.n597 163.367
R655 B.n597 B.n596 163.367
R656 B.n596 B.n121 163.367
R657 B.n592 B.n121 163.367
R658 B.n592 B.n591 163.367
R659 B.n591 B.n590 163.367
R660 B.n590 B.n123 163.367
R661 B.n586 B.n123 163.367
R662 B.n586 B.n585 163.367
R663 B.n585 B.n584 163.367
R664 B.n584 B.n125 163.367
R665 B.n580 B.n125 163.367
R666 B.n580 B.n579 163.367
R667 B.n579 B.n578 163.367
R668 B.n578 B.n127 163.367
R669 B.n574 B.n127 163.367
R670 B.n574 B.n573 163.367
R671 B.n573 B.n572 163.367
R672 B.n572 B.n129 163.367
R673 B.n568 B.n129 163.367
R674 B.n568 B.n567 163.367
R675 B.n567 B.n566 163.367
R676 B.n566 B.n131 163.367
R677 B.n562 B.n131 163.367
R678 B.n562 B.n561 163.367
R679 B.n561 B.n560 163.367
R680 B.n560 B.n133 163.367
R681 B.n556 B.n133 163.367
R682 B.n556 B.n555 163.367
R683 B.n555 B.n554 163.367
R684 B.n554 B.n135 163.367
R685 B.n550 B.n135 163.367
R686 B.n550 B.n549 163.367
R687 B.n549 B.n548 163.367
R688 B.n548 B.n137 163.367
R689 B.n544 B.n137 163.367
R690 B.n544 B.n543 163.367
R691 B.n543 B.n542 163.367
R692 B.n542 B.n139 163.367
R693 B.n538 B.n139 163.367
R694 B.n538 B.n537 163.367
R695 B.n537 B.n536 163.367
R696 B.n536 B.n141 163.367
R697 B.n532 B.n141 163.367
R698 B.n532 B.n531 163.367
R699 B.n531 B.n530 163.367
R700 B.n530 B.n143 163.367
R701 B.n526 B.n143 163.367
R702 B.n526 B.n525 163.367
R703 B.n525 B.n524 163.367
R704 B.n524 B.n145 163.367
R705 B.n520 B.n145 163.367
R706 B.n520 B.n519 163.367
R707 B.n519 B.n518 163.367
R708 B.n518 B.n147 163.367
R709 B.n514 B.n147 163.367
R710 B.n862 B.n27 163.367
R711 B.n862 B.n861 163.367
R712 B.n861 B.n860 163.367
R713 B.n860 B.n29 163.367
R714 B.n856 B.n29 163.367
R715 B.n856 B.n855 163.367
R716 B.n855 B.n854 163.367
R717 B.n854 B.n31 163.367
R718 B.n850 B.n31 163.367
R719 B.n850 B.n849 163.367
R720 B.n849 B.n848 163.367
R721 B.n848 B.n33 163.367
R722 B.n844 B.n33 163.367
R723 B.n844 B.n843 163.367
R724 B.n843 B.n842 163.367
R725 B.n842 B.n35 163.367
R726 B.n838 B.n35 163.367
R727 B.n838 B.n837 163.367
R728 B.n837 B.n836 163.367
R729 B.n836 B.n37 163.367
R730 B.n832 B.n37 163.367
R731 B.n832 B.n831 163.367
R732 B.n831 B.n830 163.367
R733 B.n830 B.n39 163.367
R734 B.n826 B.n39 163.367
R735 B.n826 B.n825 163.367
R736 B.n825 B.n824 163.367
R737 B.n824 B.n41 163.367
R738 B.n820 B.n41 163.367
R739 B.n820 B.n819 163.367
R740 B.n819 B.n818 163.367
R741 B.n818 B.n43 163.367
R742 B.n814 B.n43 163.367
R743 B.n814 B.n813 163.367
R744 B.n813 B.n812 163.367
R745 B.n812 B.n45 163.367
R746 B.n808 B.n45 163.367
R747 B.n808 B.n807 163.367
R748 B.n807 B.n806 163.367
R749 B.n806 B.n47 163.367
R750 B.n802 B.n47 163.367
R751 B.n802 B.n801 163.367
R752 B.n801 B.n800 163.367
R753 B.n800 B.n49 163.367
R754 B.n796 B.n49 163.367
R755 B.n796 B.n795 163.367
R756 B.n795 B.n794 163.367
R757 B.n794 B.n51 163.367
R758 B.n790 B.n51 163.367
R759 B.n790 B.n789 163.367
R760 B.n789 B.n788 163.367
R761 B.n788 B.n53 163.367
R762 B.n784 B.n53 163.367
R763 B.n784 B.n783 163.367
R764 B.n783 B.n782 163.367
R765 B.n782 B.n55 163.367
R766 B.n778 B.n55 163.367
R767 B.n778 B.n777 163.367
R768 B.n777 B.n776 163.367
R769 B.n776 B.n57 163.367
R770 B.n771 B.n57 163.367
R771 B.n771 B.n770 163.367
R772 B.n770 B.n769 163.367
R773 B.n769 B.n61 163.367
R774 B.n765 B.n61 163.367
R775 B.n765 B.n764 163.367
R776 B.n764 B.n763 163.367
R777 B.n763 B.n63 163.367
R778 B.n759 B.n63 163.367
R779 B.n759 B.n758 163.367
R780 B.n758 B.n67 163.367
R781 B.n754 B.n67 163.367
R782 B.n754 B.n753 163.367
R783 B.n753 B.n752 163.367
R784 B.n752 B.n69 163.367
R785 B.n748 B.n69 163.367
R786 B.n748 B.n747 163.367
R787 B.n747 B.n746 163.367
R788 B.n746 B.n71 163.367
R789 B.n742 B.n71 163.367
R790 B.n742 B.n741 163.367
R791 B.n741 B.n740 163.367
R792 B.n740 B.n73 163.367
R793 B.n736 B.n73 163.367
R794 B.n736 B.n735 163.367
R795 B.n735 B.n734 163.367
R796 B.n734 B.n75 163.367
R797 B.n730 B.n75 163.367
R798 B.n730 B.n729 163.367
R799 B.n729 B.n728 163.367
R800 B.n728 B.n77 163.367
R801 B.n724 B.n77 163.367
R802 B.n724 B.n723 163.367
R803 B.n723 B.n722 163.367
R804 B.n722 B.n79 163.367
R805 B.n718 B.n79 163.367
R806 B.n718 B.n717 163.367
R807 B.n717 B.n716 163.367
R808 B.n716 B.n81 163.367
R809 B.n712 B.n81 163.367
R810 B.n712 B.n711 163.367
R811 B.n711 B.n710 163.367
R812 B.n710 B.n83 163.367
R813 B.n706 B.n83 163.367
R814 B.n706 B.n705 163.367
R815 B.n705 B.n704 163.367
R816 B.n704 B.n85 163.367
R817 B.n700 B.n85 163.367
R818 B.n700 B.n699 163.367
R819 B.n699 B.n698 163.367
R820 B.n698 B.n87 163.367
R821 B.n694 B.n87 163.367
R822 B.n694 B.n693 163.367
R823 B.n693 B.n692 163.367
R824 B.n692 B.n89 163.367
R825 B.n688 B.n89 163.367
R826 B.n688 B.n687 163.367
R827 B.n687 B.n686 163.367
R828 B.n686 B.n91 163.367
R829 B.n682 B.n91 163.367
R830 B.n682 B.n681 163.367
R831 B.n681 B.n680 163.367
R832 B.n680 B.n93 163.367
R833 B.n676 B.n93 163.367
R834 B.n676 B.n675 163.367
R835 B.n675 B.n674 163.367
R836 B.n674 B.n95 163.367
R837 B.n670 B.n95 163.367
R838 B.n670 B.n669 163.367
R839 B.n669 B.n668 163.367
R840 B.n867 B.n866 163.367
R841 B.n868 B.n867 163.367
R842 B.n868 B.n25 163.367
R843 B.n872 B.n25 163.367
R844 B.n873 B.n872 163.367
R845 B.n874 B.n873 163.367
R846 B.n874 B.n23 163.367
R847 B.n878 B.n23 163.367
R848 B.n879 B.n878 163.367
R849 B.n880 B.n879 163.367
R850 B.n880 B.n21 163.367
R851 B.n884 B.n21 163.367
R852 B.n885 B.n884 163.367
R853 B.n886 B.n885 163.367
R854 B.n886 B.n19 163.367
R855 B.n890 B.n19 163.367
R856 B.n891 B.n890 163.367
R857 B.n892 B.n891 163.367
R858 B.n892 B.n17 163.367
R859 B.n896 B.n17 163.367
R860 B.n897 B.n896 163.367
R861 B.n898 B.n897 163.367
R862 B.n898 B.n15 163.367
R863 B.n902 B.n15 163.367
R864 B.n903 B.n902 163.367
R865 B.n904 B.n903 163.367
R866 B.n904 B.n13 163.367
R867 B.n908 B.n13 163.367
R868 B.n909 B.n908 163.367
R869 B.n910 B.n909 163.367
R870 B.n910 B.n11 163.367
R871 B.n914 B.n11 163.367
R872 B.n915 B.n914 163.367
R873 B.n916 B.n915 163.367
R874 B.n916 B.n9 163.367
R875 B.n920 B.n9 163.367
R876 B.n921 B.n920 163.367
R877 B.n922 B.n921 163.367
R878 B.n922 B.n7 163.367
R879 B.n926 B.n7 163.367
R880 B.n927 B.n926 163.367
R881 B.n928 B.n927 163.367
R882 B.n928 B.n5 163.367
R883 B.n932 B.n5 163.367
R884 B.n933 B.n932 163.367
R885 B.n934 B.n933 163.367
R886 B.n934 B.n3 163.367
R887 B.n938 B.n3 163.367
R888 B.n939 B.n938 163.367
R889 B.n240 B.n2 163.367
R890 B.n240 B.n239 163.367
R891 B.n244 B.n239 163.367
R892 B.n245 B.n244 163.367
R893 B.n246 B.n245 163.367
R894 B.n246 B.n237 163.367
R895 B.n250 B.n237 163.367
R896 B.n251 B.n250 163.367
R897 B.n252 B.n251 163.367
R898 B.n252 B.n235 163.367
R899 B.n256 B.n235 163.367
R900 B.n257 B.n256 163.367
R901 B.n258 B.n257 163.367
R902 B.n258 B.n233 163.367
R903 B.n262 B.n233 163.367
R904 B.n263 B.n262 163.367
R905 B.n264 B.n263 163.367
R906 B.n264 B.n231 163.367
R907 B.n268 B.n231 163.367
R908 B.n269 B.n268 163.367
R909 B.n270 B.n269 163.367
R910 B.n270 B.n229 163.367
R911 B.n274 B.n229 163.367
R912 B.n275 B.n274 163.367
R913 B.n276 B.n275 163.367
R914 B.n276 B.n227 163.367
R915 B.n280 B.n227 163.367
R916 B.n281 B.n280 163.367
R917 B.n282 B.n281 163.367
R918 B.n282 B.n225 163.367
R919 B.n286 B.n225 163.367
R920 B.n287 B.n286 163.367
R921 B.n288 B.n287 163.367
R922 B.n288 B.n223 163.367
R923 B.n292 B.n223 163.367
R924 B.n293 B.n292 163.367
R925 B.n294 B.n293 163.367
R926 B.n294 B.n221 163.367
R927 B.n298 B.n221 163.367
R928 B.n299 B.n298 163.367
R929 B.n300 B.n299 163.367
R930 B.n300 B.n219 163.367
R931 B.n304 B.n219 163.367
R932 B.n305 B.n304 163.367
R933 B.n306 B.n305 163.367
R934 B.n306 B.n217 163.367
R935 B.n310 B.n217 163.367
R936 B.n311 B.n310 163.367
R937 B.n312 B.n311 163.367
R938 B.n419 B.t2 108.293
R939 B.n65 B.t4 108.293
R940 B.n185 B.t11 108.269
R941 B.n59 B.t7 108.269
R942 B.n185 B.n184 70.2066
R943 B.n419 B.n418 70.2066
R944 B.n65 B.n64 70.2066
R945 B.n59 B.n58 70.2066
R946 B.n405 B.n185 59.5399
R947 B.n420 B.n419 59.5399
R948 B.n66 B.n65 59.5399
R949 B.n773 B.n59 59.5399
R950 B.n865 B.n864 33.8737
R951 B.n667 B.n666 33.8737
R952 B.n515 B.n148 33.8737
R953 B.n314 B.n313 33.8737
R954 B B.n941 18.0485
R955 B.n865 B.n26 10.6151
R956 B.n869 B.n26 10.6151
R957 B.n870 B.n869 10.6151
R958 B.n871 B.n870 10.6151
R959 B.n871 B.n24 10.6151
R960 B.n875 B.n24 10.6151
R961 B.n876 B.n875 10.6151
R962 B.n877 B.n876 10.6151
R963 B.n877 B.n22 10.6151
R964 B.n881 B.n22 10.6151
R965 B.n882 B.n881 10.6151
R966 B.n883 B.n882 10.6151
R967 B.n883 B.n20 10.6151
R968 B.n887 B.n20 10.6151
R969 B.n888 B.n887 10.6151
R970 B.n889 B.n888 10.6151
R971 B.n889 B.n18 10.6151
R972 B.n893 B.n18 10.6151
R973 B.n894 B.n893 10.6151
R974 B.n895 B.n894 10.6151
R975 B.n895 B.n16 10.6151
R976 B.n899 B.n16 10.6151
R977 B.n900 B.n899 10.6151
R978 B.n901 B.n900 10.6151
R979 B.n901 B.n14 10.6151
R980 B.n905 B.n14 10.6151
R981 B.n906 B.n905 10.6151
R982 B.n907 B.n906 10.6151
R983 B.n907 B.n12 10.6151
R984 B.n911 B.n12 10.6151
R985 B.n912 B.n911 10.6151
R986 B.n913 B.n912 10.6151
R987 B.n913 B.n10 10.6151
R988 B.n917 B.n10 10.6151
R989 B.n918 B.n917 10.6151
R990 B.n919 B.n918 10.6151
R991 B.n919 B.n8 10.6151
R992 B.n923 B.n8 10.6151
R993 B.n924 B.n923 10.6151
R994 B.n925 B.n924 10.6151
R995 B.n925 B.n6 10.6151
R996 B.n929 B.n6 10.6151
R997 B.n930 B.n929 10.6151
R998 B.n931 B.n930 10.6151
R999 B.n931 B.n4 10.6151
R1000 B.n935 B.n4 10.6151
R1001 B.n936 B.n935 10.6151
R1002 B.n937 B.n936 10.6151
R1003 B.n937 B.n0 10.6151
R1004 B.n864 B.n863 10.6151
R1005 B.n863 B.n28 10.6151
R1006 B.n859 B.n28 10.6151
R1007 B.n859 B.n858 10.6151
R1008 B.n858 B.n857 10.6151
R1009 B.n857 B.n30 10.6151
R1010 B.n853 B.n30 10.6151
R1011 B.n853 B.n852 10.6151
R1012 B.n852 B.n851 10.6151
R1013 B.n851 B.n32 10.6151
R1014 B.n847 B.n32 10.6151
R1015 B.n847 B.n846 10.6151
R1016 B.n846 B.n845 10.6151
R1017 B.n845 B.n34 10.6151
R1018 B.n841 B.n34 10.6151
R1019 B.n841 B.n840 10.6151
R1020 B.n840 B.n839 10.6151
R1021 B.n839 B.n36 10.6151
R1022 B.n835 B.n36 10.6151
R1023 B.n835 B.n834 10.6151
R1024 B.n834 B.n833 10.6151
R1025 B.n833 B.n38 10.6151
R1026 B.n829 B.n38 10.6151
R1027 B.n829 B.n828 10.6151
R1028 B.n828 B.n827 10.6151
R1029 B.n827 B.n40 10.6151
R1030 B.n823 B.n40 10.6151
R1031 B.n823 B.n822 10.6151
R1032 B.n822 B.n821 10.6151
R1033 B.n821 B.n42 10.6151
R1034 B.n817 B.n42 10.6151
R1035 B.n817 B.n816 10.6151
R1036 B.n816 B.n815 10.6151
R1037 B.n815 B.n44 10.6151
R1038 B.n811 B.n44 10.6151
R1039 B.n811 B.n810 10.6151
R1040 B.n810 B.n809 10.6151
R1041 B.n809 B.n46 10.6151
R1042 B.n805 B.n46 10.6151
R1043 B.n805 B.n804 10.6151
R1044 B.n804 B.n803 10.6151
R1045 B.n803 B.n48 10.6151
R1046 B.n799 B.n48 10.6151
R1047 B.n799 B.n798 10.6151
R1048 B.n798 B.n797 10.6151
R1049 B.n797 B.n50 10.6151
R1050 B.n793 B.n50 10.6151
R1051 B.n793 B.n792 10.6151
R1052 B.n792 B.n791 10.6151
R1053 B.n791 B.n52 10.6151
R1054 B.n787 B.n52 10.6151
R1055 B.n787 B.n786 10.6151
R1056 B.n786 B.n785 10.6151
R1057 B.n785 B.n54 10.6151
R1058 B.n781 B.n54 10.6151
R1059 B.n781 B.n780 10.6151
R1060 B.n780 B.n779 10.6151
R1061 B.n779 B.n56 10.6151
R1062 B.n775 B.n56 10.6151
R1063 B.n775 B.n774 10.6151
R1064 B.n772 B.n60 10.6151
R1065 B.n768 B.n60 10.6151
R1066 B.n768 B.n767 10.6151
R1067 B.n767 B.n766 10.6151
R1068 B.n766 B.n62 10.6151
R1069 B.n762 B.n62 10.6151
R1070 B.n762 B.n761 10.6151
R1071 B.n761 B.n760 10.6151
R1072 B.n757 B.n756 10.6151
R1073 B.n756 B.n755 10.6151
R1074 B.n755 B.n68 10.6151
R1075 B.n751 B.n68 10.6151
R1076 B.n751 B.n750 10.6151
R1077 B.n750 B.n749 10.6151
R1078 B.n749 B.n70 10.6151
R1079 B.n745 B.n70 10.6151
R1080 B.n745 B.n744 10.6151
R1081 B.n744 B.n743 10.6151
R1082 B.n743 B.n72 10.6151
R1083 B.n739 B.n72 10.6151
R1084 B.n739 B.n738 10.6151
R1085 B.n738 B.n737 10.6151
R1086 B.n737 B.n74 10.6151
R1087 B.n733 B.n74 10.6151
R1088 B.n733 B.n732 10.6151
R1089 B.n732 B.n731 10.6151
R1090 B.n731 B.n76 10.6151
R1091 B.n727 B.n76 10.6151
R1092 B.n727 B.n726 10.6151
R1093 B.n726 B.n725 10.6151
R1094 B.n725 B.n78 10.6151
R1095 B.n721 B.n78 10.6151
R1096 B.n721 B.n720 10.6151
R1097 B.n720 B.n719 10.6151
R1098 B.n719 B.n80 10.6151
R1099 B.n715 B.n80 10.6151
R1100 B.n715 B.n714 10.6151
R1101 B.n714 B.n713 10.6151
R1102 B.n713 B.n82 10.6151
R1103 B.n709 B.n82 10.6151
R1104 B.n709 B.n708 10.6151
R1105 B.n708 B.n707 10.6151
R1106 B.n707 B.n84 10.6151
R1107 B.n703 B.n84 10.6151
R1108 B.n703 B.n702 10.6151
R1109 B.n702 B.n701 10.6151
R1110 B.n701 B.n86 10.6151
R1111 B.n697 B.n86 10.6151
R1112 B.n697 B.n696 10.6151
R1113 B.n696 B.n695 10.6151
R1114 B.n695 B.n88 10.6151
R1115 B.n691 B.n88 10.6151
R1116 B.n691 B.n690 10.6151
R1117 B.n690 B.n689 10.6151
R1118 B.n689 B.n90 10.6151
R1119 B.n685 B.n90 10.6151
R1120 B.n685 B.n684 10.6151
R1121 B.n684 B.n683 10.6151
R1122 B.n683 B.n92 10.6151
R1123 B.n679 B.n92 10.6151
R1124 B.n679 B.n678 10.6151
R1125 B.n678 B.n677 10.6151
R1126 B.n677 B.n94 10.6151
R1127 B.n673 B.n94 10.6151
R1128 B.n673 B.n672 10.6151
R1129 B.n672 B.n671 10.6151
R1130 B.n671 B.n96 10.6151
R1131 B.n667 B.n96 10.6151
R1132 B.n666 B.n665 10.6151
R1133 B.n665 B.n98 10.6151
R1134 B.n661 B.n98 10.6151
R1135 B.n661 B.n660 10.6151
R1136 B.n660 B.n659 10.6151
R1137 B.n659 B.n100 10.6151
R1138 B.n655 B.n100 10.6151
R1139 B.n655 B.n654 10.6151
R1140 B.n654 B.n653 10.6151
R1141 B.n653 B.n102 10.6151
R1142 B.n649 B.n102 10.6151
R1143 B.n649 B.n648 10.6151
R1144 B.n648 B.n647 10.6151
R1145 B.n647 B.n104 10.6151
R1146 B.n643 B.n104 10.6151
R1147 B.n643 B.n642 10.6151
R1148 B.n642 B.n641 10.6151
R1149 B.n641 B.n106 10.6151
R1150 B.n637 B.n106 10.6151
R1151 B.n637 B.n636 10.6151
R1152 B.n636 B.n635 10.6151
R1153 B.n635 B.n108 10.6151
R1154 B.n631 B.n108 10.6151
R1155 B.n631 B.n630 10.6151
R1156 B.n630 B.n629 10.6151
R1157 B.n629 B.n110 10.6151
R1158 B.n625 B.n110 10.6151
R1159 B.n625 B.n624 10.6151
R1160 B.n624 B.n623 10.6151
R1161 B.n623 B.n112 10.6151
R1162 B.n619 B.n112 10.6151
R1163 B.n619 B.n618 10.6151
R1164 B.n618 B.n617 10.6151
R1165 B.n617 B.n114 10.6151
R1166 B.n613 B.n114 10.6151
R1167 B.n613 B.n612 10.6151
R1168 B.n612 B.n611 10.6151
R1169 B.n611 B.n116 10.6151
R1170 B.n607 B.n116 10.6151
R1171 B.n607 B.n606 10.6151
R1172 B.n606 B.n605 10.6151
R1173 B.n605 B.n118 10.6151
R1174 B.n601 B.n118 10.6151
R1175 B.n601 B.n600 10.6151
R1176 B.n600 B.n599 10.6151
R1177 B.n599 B.n120 10.6151
R1178 B.n595 B.n120 10.6151
R1179 B.n595 B.n594 10.6151
R1180 B.n594 B.n593 10.6151
R1181 B.n593 B.n122 10.6151
R1182 B.n589 B.n122 10.6151
R1183 B.n589 B.n588 10.6151
R1184 B.n588 B.n587 10.6151
R1185 B.n587 B.n124 10.6151
R1186 B.n583 B.n124 10.6151
R1187 B.n583 B.n582 10.6151
R1188 B.n582 B.n581 10.6151
R1189 B.n581 B.n126 10.6151
R1190 B.n577 B.n126 10.6151
R1191 B.n577 B.n576 10.6151
R1192 B.n576 B.n575 10.6151
R1193 B.n575 B.n128 10.6151
R1194 B.n571 B.n128 10.6151
R1195 B.n571 B.n570 10.6151
R1196 B.n570 B.n569 10.6151
R1197 B.n569 B.n130 10.6151
R1198 B.n565 B.n130 10.6151
R1199 B.n565 B.n564 10.6151
R1200 B.n564 B.n563 10.6151
R1201 B.n563 B.n132 10.6151
R1202 B.n559 B.n132 10.6151
R1203 B.n559 B.n558 10.6151
R1204 B.n558 B.n557 10.6151
R1205 B.n557 B.n134 10.6151
R1206 B.n553 B.n134 10.6151
R1207 B.n553 B.n552 10.6151
R1208 B.n552 B.n551 10.6151
R1209 B.n551 B.n136 10.6151
R1210 B.n547 B.n136 10.6151
R1211 B.n547 B.n546 10.6151
R1212 B.n546 B.n545 10.6151
R1213 B.n545 B.n138 10.6151
R1214 B.n541 B.n138 10.6151
R1215 B.n541 B.n540 10.6151
R1216 B.n540 B.n539 10.6151
R1217 B.n539 B.n140 10.6151
R1218 B.n535 B.n140 10.6151
R1219 B.n535 B.n534 10.6151
R1220 B.n534 B.n533 10.6151
R1221 B.n533 B.n142 10.6151
R1222 B.n529 B.n142 10.6151
R1223 B.n529 B.n528 10.6151
R1224 B.n528 B.n527 10.6151
R1225 B.n527 B.n144 10.6151
R1226 B.n523 B.n144 10.6151
R1227 B.n523 B.n522 10.6151
R1228 B.n522 B.n521 10.6151
R1229 B.n521 B.n146 10.6151
R1230 B.n517 B.n146 10.6151
R1231 B.n517 B.n516 10.6151
R1232 B.n516 B.n515 10.6151
R1233 B.n241 B.n1 10.6151
R1234 B.n242 B.n241 10.6151
R1235 B.n243 B.n242 10.6151
R1236 B.n243 B.n238 10.6151
R1237 B.n247 B.n238 10.6151
R1238 B.n248 B.n247 10.6151
R1239 B.n249 B.n248 10.6151
R1240 B.n249 B.n236 10.6151
R1241 B.n253 B.n236 10.6151
R1242 B.n254 B.n253 10.6151
R1243 B.n255 B.n254 10.6151
R1244 B.n255 B.n234 10.6151
R1245 B.n259 B.n234 10.6151
R1246 B.n260 B.n259 10.6151
R1247 B.n261 B.n260 10.6151
R1248 B.n261 B.n232 10.6151
R1249 B.n265 B.n232 10.6151
R1250 B.n266 B.n265 10.6151
R1251 B.n267 B.n266 10.6151
R1252 B.n267 B.n230 10.6151
R1253 B.n271 B.n230 10.6151
R1254 B.n272 B.n271 10.6151
R1255 B.n273 B.n272 10.6151
R1256 B.n273 B.n228 10.6151
R1257 B.n277 B.n228 10.6151
R1258 B.n278 B.n277 10.6151
R1259 B.n279 B.n278 10.6151
R1260 B.n279 B.n226 10.6151
R1261 B.n283 B.n226 10.6151
R1262 B.n284 B.n283 10.6151
R1263 B.n285 B.n284 10.6151
R1264 B.n285 B.n224 10.6151
R1265 B.n289 B.n224 10.6151
R1266 B.n290 B.n289 10.6151
R1267 B.n291 B.n290 10.6151
R1268 B.n291 B.n222 10.6151
R1269 B.n295 B.n222 10.6151
R1270 B.n296 B.n295 10.6151
R1271 B.n297 B.n296 10.6151
R1272 B.n297 B.n220 10.6151
R1273 B.n301 B.n220 10.6151
R1274 B.n302 B.n301 10.6151
R1275 B.n303 B.n302 10.6151
R1276 B.n303 B.n218 10.6151
R1277 B.n307 B.n218 10.6151
R1278 B.n308 B.n307 10.6151
R1279 B.n309 B.n308 10.6151
R1280 B.n309 B.n216 10.6151
R1281 B.n313 B.n216 10.6151
R1282 B.n315 B.n314 10.6151
R1283 B.n315 B.n214 10.6151
R1284 B.n319 B.n214 10.6151
R1285 B.n320 B.n319 10.6151
R1286 B.n321 B.n320 10.6151
R1287 B.n321 B.n212 10.6151
R1288 B.n325 B.n212 10.6151
R1289 B.n326 B.n325 10.6151
R1290 B.n327 B.n326 10.6151
R1291 B.n327 B.n210 10.6151
R1292 B.n331 B.n210 10.6151
R1293 B.n332 B.n331 10.6151
R1294 B.n333 B.n332 10.6151
R1295 B.n333 B.n208 10.6151
R1296 B.n337 B.n208 10.6151
R1297 B.n338 B.n337 10.6151
R1298 B.n339 B.n338 10.6151
R1299 B.n339 B.n206 10.6151
R1300 B.n343 B.n206 10.6151
R1301 B.n344 B.n343 10.6151
R1302 B.n345 B.n344 10.6151
R1303 B.n345 B.n204 10.6151
R1304 B.n349 B.n204 10.6151
R1305 B.n350 B.n349 10.6151
R1306 B.n351 B.n350 10.6151
R1307 B.n351 B.n202 10.6151
R1308 B.n355 B.n202 10.6151
R1309 B.n356 B.n355 10.6151
R1310 B.n357 B.n356 10.6151
R1311 B.n357 B.n200 10.6151
R1312 B.n361 B.n200 10.6151
R1313 B.n362 B.n361 10.6151
R1314 B.n363 B.n362 10.6151
R1315 B.n363 B.n198 10.6151
R1316 B.n367 B.n198 10.6151
R1317 B.n368 B.n367 10.6151
R1318 B.n369 B.n368 10.6151
R1319 B.n369 B.n196 10.6151
R1320 B.n373 B.n196 10.6151
R1321 B.n374 B.n373 10.6151
R1322 B.n375 B.n374 10.6151
R1323 B.n375 B.n194 10.6151
R1324 B.n379 B.n194 10.6151
R1325 B.n380 B.n379 10.6151
R1326 B.n381 B.n380 10.6151
R1327 B.n381 B.n192 10.6151
R1328 B.n385 B.n192 10.6151
R1329 B.n386 B.n385 10.6151
R1330 B.n387 B.n386 10.6151
R1331 B.n387 B.n190 10.6151
R1332 B.n391 B.n190 10.6151
R1333 B.n392 B.n391 10.6151
R1334 B.n393 B.n392 10.6151
R1335 B.n393 B.n188 10.6151
R1336 B.n397 B.n188 10.6151
R1337 B.n398 B.n397 10.6151
R1338 B.n399 B.n398 10.6151
R1339 B.n399 B.n186 10.6151
R1340 B.n403 B.n186 10.6151
R1341 B.n404 B.n403 10.6151
R1342 B.n406 B.n182 10.6151
R1343 B.n410 B.n182 10.6151
R1344 B.n411 B.n410 10.6151
R1345 B.n412 B.n411 10.6151
R1346 B.n412 B.n180 10.6151
R1347 B.n416 B.n180 10.6151
R1348 B.n417 B.n416 10.6151
R1349 B.n421 B.n417 10.6151
R1350 B.n425 B.n178 10.6151
R1351 B.n426 B.n425 10.6151
R1352 B.n427 B.n426 10.6151
R1353 B.n427 B.n176 10.6151
R1354 B.n431 B.n176 10.6151
R1355 B.n432 B.n431 10.6151
R1356 B.n433 B.n432 10.6151
R1357 B.n433 B.n174 10.6151
R1358 B.n437 B.n174 10.6151
R1359 B.n438 B.n437 10.6151
R1360 B.n439 B.n438 10.6151
R1361 B.n439 B.n172 10.6151
R1362 B.n443 B.n172 10.6151
R1363 B.n444 B.n443 10.6151
R1364 B.n445 B.n444 10.6151
R1365 B.n445 B.n170 10.6151
R1366 B.n449 B.n170 10.6151
R1367 B.n450 B.n449 10.6151
R1368 B.n451 B.n450 10.6151
R1369 B.n451 B.n168 10.6151
R1370 B.n455 B.n168 10.6151
R1371 B.n456 B.n455 10.6151
R1372 B.n457 B.n456 10.6151
R1373 B.n457 B.n166 10.6151
R1374 B.n461 B.n166 10.6151
R1375 B.n462 B.n461 10.6151
R1376 B.n463 B.n462 10.6151
R1377 B.n463 B.n164 10.6151
R1378 B.n467 B.n164 10.6151
R1379 B.n468 B.n467 10.6151
R1380 B.n469 B.n468 10.6151
R1381 B.n469 B.n162 10.6151
R1382 B.n473 B.n162 10.6151
R1383 B.n474 B.n473 10.6151
R1384 B.n475 B.n474 10.6151
R1385 B.n475 B.n160 10.6151
R1386 B.n479 B.n160 10.6151
R1387 B.n480 B.n479 10.6151
R1388 B.n481 B.n480 10.6151
R1389 B.n481 B.n158 10.6151
R1390 B.n485 B.n158 10.6151
R1391 B.n486 B.n485 10.6151
R1392 B.n487 B.n486 10.6151
R1393 B.n487 B.n156 10.6151
R1394 B.n491 B.n156 10.6151
R1395 B.n492 B.n491 10.6151
R1396 B.n493 B.n492 10.6151
R1397 B.n493 B.n154 10.6151
R1398 B.n497 B.n154 10.6151
R1399 B.n498 B.n497 10.6151
R1400 B.n499 B.n498 10.6151
R1401 B.n499 B.n152 10.6151
R1402 B.n503 B.n152 10.6151
R1403 B.n504 B.n503 10.6151
R1404 B.n505 B.n504 10.6151
R1405 B.n505 B.n150 10.6151
R1406 B.n509 B.n150 10.6151
R1407 B.n510 B.n509 10.6151
R1408 B.n511 B.n510 10.6151
R1409 B.n511 B.n148 10.6151
R1410 B.n941 B.n0 8.11757
R1411 B.n941 B.n1 8.11757
R1412 B.n773 B.n772 6.5566
R1413 B.n760 B.n66 6.5566
R1414 B.n406 B.n405 6.5566
R1415 B.n421 B.n420 6.5566
R1416 B.n774 B.n773 4.05904
R1417 B.n757 B.n66 4.05904
R1418 B.n405 B.n404 4.05904
R1419 B.n420 B.n178 4.05904
R1420 VN.n23 VN.t1 168.543
R1421 VN.n5 VN.t5 168.543
R1422 VN.n34 VN.n33 161.3
R1423 VN.n32 VN.n19 161.3
R1424 VN.n31 VN.n30 161.3
R1425 VN.n29 VN.n20 161.3
R1426 VN.n28 VN.n27 161.3
R1427 VN.n26 VN.n21 161.3
R1428 VN.n25 VN.n24 161.3
R1429 VN.n16 VN.n15 161.3
R1430 VN.n14 VN.n1 161.3
R1431 VN.n13 VN.n12 161.3
R1432 VN.n11 VN.n2 161.3
R1433 VN.n10 VN.n9 161.3
R1434 VN.n8 VN.n3 161.3
R1435 VN.n7 VN.n6 161.3
R1436 VN.n4 VN.t3 135.298
R1437 VN.n0 VN.t0 135.298
R1438 VN.n22 VN.t2 135.298
R1439 VN.n18 VN.t4 135.298
R1440 VN.n17 VN.n0 71.9618
R1441 VN.n35 VN.n18 71.9618
R1442 VN.n5 VN.n4 62.0558
R1443 VN.n23 VN.n22 62.0558
R1444 VN VN.n35 56.6117
R1445 VN.n13 VN.n2 46.321
R1446 VN.n31 VN.n20 46.321
R1447 VN.n9 VN.n2 34.6658
R1448 VN.n27 VN.n20 34.6658
R1449 VN.n8 VN.n7 24.4675
R1450 VN.n9 VN.n8 24.4675
R1451 VN.n14 VN.n13 24.4675
R1452 VN.n15 VN.n14 24.4675
R1453 VN.n27 VN.n26 24.4675
R1454 VN.n26 VN.n25 24.4675
R1455 VN.n33 VN.n32 24.4675
R1456 VN.n32 VN.n31 24.4675
R1457 VN.n15 VN.n0 18.1061
R1458 VN.n33 VN.n18 18.1061
R1459 VN.n7 VN.n4 12.234
R1460 VN.n25 VN.n22 12.234
R1461 VN.n6 VN.n5 3.99399
R1462 VN.n24 VN.n23 3.99399
R1463 VN.n35 VN.n34 0.354971
R1464 VN.n17 VN.n16 0.354971
R1465 VN VN.n17 0.26696
R1466 VN.n34 VN.n19 0.189894
R1467 VN.n30 VN.n19 0.189894
R1468 VN.n30 VN.n29 0.189894
R1469 VN.n29 VN.n28 0.189894
R1470 VN.n28 VN.n21 0.189894
R1471 VN.n24 VN.n21 0.189894
R1472 VN.n6 VN.n3 0.189894
R1473 VN.n10 VN.n3 0.189894
R1474 VN.n11 VN.n10 0.189894
R1475 VN.n12 VN.n11 0.189894
R1476 VN.n12 VN.n1 0.189894
R1477 VN.n16 VN.n1 0.189894
R1478 VTAIL.n7 VTAIL.t6 57.7515
R1479 VTAIL.n11 VTAIL.t10 57.7504
R1480 VTAIL.n2 VTAIL.t1 57.7504
R1481 VTAIL.n10 VTAIL.t5 57.7503
R1482 VTAIL.n9 VTAIL.n8 55.9916
R1483 VTAIL.n6 VTAIL.n5 55.9916
R1484 VTAIL.n1 VTAIL.n0 55.9914
R1485 VTAIL.n4 VTAIL.n3 55.9914
R1486 VTAIL.n6 VTAIL.n4 34.5307
R1487 VTAIL.n11 VTAIL.n10 31.41
R1488 VTAIL.n7 VTAIL.n6 3.12119
R1489 VTAIL.n10 VTAIL.n9 3.12119
R1490 VTAIL.n4 VTAIL.n2 3.12119
R1491 VTAIL VTAIL.n11 2.28283
R1492 VTAIL.n9 VTAIL.n7 2.03067
R1493 VTAIL.n2 VTAIL.n1 2.03067
R1494 VTAIL.n0 VTAIL.t11 1.76038
R1495 VTAIL.n0 VTAIL.t7 1.76038
R1496 VTAIL.n3 VTAIL.t2 1.76038
R1497 VTAIL.n3 VTAIL.t4 1.76038
R1498 VTAIL.n8 VTAIL.t3 1.76038
R1499 VTAIL.n8 VTAIL.t0 1.76038
R1500 VTAIL.n5 VTAIL.t9 1.76038
R1501 VTAIL.n5 VTAIL.t8 1.76038
R1502 VTAIL VTAIL.n1 0.838862
R1503 VDD2.n1 VDD2.t0 76.7144
R1504 VDD2.n2 VDD2.t1 74.4302
R1505 VDD2.n1 VDD2.n0 73.395
R1506 VDD2 VDD2.n3 73.3912
R1507 VDD2.n2 VDD2.n1 49.7799
R1508 VDD2 VDD2.n2 2.39921
R1509 VDD2.n3 VDD2.t3 1.76038
R1510 VDD2.n3 VDD2.t4 1.76038
R1511 VDD2.n0 VDD2.t2 1.76038
R1512 VDD2.n0 VDD2.t5 1.76038
R1513 VP.n14 VP.t2 168.543
R1514 VP.n16 VP.n15 161.3
R1515 VP.n17 VP.n12 161.3
R1516 VP.n19 VP.n18 161.3
R1517 VP.n20 VP.n11 161.3
R1518 VP.n22 VP.n21 161.3
R1519 VP.n23 VP.n10 161.3
R1520 VP.n25 VP.n24 161.3
R1521 VP.n49 VP.n48 161.3
R1522 VP.n47 VP.n1 161.3
R1523 VP.n46 VP.n45 161.3
R1524 VP.n44 VP.n2 161.3
R1525 VP.n43 VP.n42 161.3
R1526 VP.n41 VP.n3 161.3
R1527 VP.n40 VP.n39 161.3
R1528 VP.n38 VP.n37 161.3
R1529 VP.n36 VP.n5 161.3
R1530 VP.n35 VP.n34 161.3
R1531 VP.n33 VP.n6 161.3
R1532 VP.n32 VP.n31 161.3
R1533 VP.n30 VP.n7 161.3
R1534 VP.n29 VP.n28 161.3
R1535 VP.n8 VP.t1 135.298
R1536 VP.n4 VP.t0 135.298
R1537 VP.n0 VP.t3 135.298
R1538 VP.n9 VP.t4 135.298
R1539 VP.n13 VP.t5 135.298
R1540 VP.n27 VP.n8 71.9618
R1541 VP.n50 VP.n0 71.9618
R1542 VP.n26 VP.n9 71.9618
R1543 VP.n14 VP.n13 62.0558
R1544 VP.n27 VP.n26 56.4463
R1545 VP.n31 VP.n6 46.321
R1546 VP.n46 VP.n2 46.321
R1547 VP.n22 VP.n11 46.321
R1548 VP.n35 VP.n6 34.6658
R1549 VP.n42 VP.n2 34.6658
R1550 VP.n18 VP.n11 34.6658
R1551 VP.n30 VP.n29 24.4675
R1552 VP.n31 VP.n30 24.4675
R1553 VP.n36 VP.n35 24.4675
R1554 VP.n37 VP.n36 24.4675
R1555 VP.n41 VP.n40 24.4675
R1556 VP.n42 VP.n41 24.4675
R1557 VP.n47 VP.n46 24.4675
R1558 VP.n48 VP.n47 24.4675
R1559 VP.n23 VP.n22 24.4675
R1560 VP.n24 VP.n23 24.4675
R1561 VP.n17 VP.n16 24.4675
R1562 VP.n18 VP.n17 24.4675
R1563 VP.n29 VP.n8 18.1061
R1564 VP.n48 VP.n0 18.1061
R1565 VP.n24 VP.n9 18.1061
R1566 VP.n37 VP.n4 12.234
R1567 VP.n40 VP.n4 12.234
R1568 VP.n16 VP.n13 12.234
R1569 VP.n15 VP.n14 3.99397
R1570 VP.n26 VP.n25 0.354971
R1571 VP.n28 VP.n27 0.354971
R1572 VP.n50 VP.n49 0.354971
R1573 VP VP.n50 0.26696
R1574 VP.n15 VP.n12 0.189894
R1575 VP.n19 VP.n12 0.189894
R1576 VP.n20 VP.n19 0.189894
R1577 VP.n21 VP.n20 0.189894
R1578 VP.n21 VP.n10 0.189894
R1579 VP.n25 VP.n10 0.189894
R1580 VP.n28 VP.n7 0.189894
R1581 VP.n32 VP.n7 0.189894
R1582 VP.n33 VP.n32 0.189894
R1583 VP.n34 VP.n33 0.189894
R1584 VP.n34 VP.n5 0.189894
R1585 VP.n38 VP.n5 0.189894
R1586 VP.n39 VP.n38 0.189894
R1587 VP.n39 VP.n3 0.189894
R1588 VP.n43 VP.n3 0.189894
R1589 VP.n44 VP.n43 0.189894
R1590 VP.n45 VP.n44 0.189894
R1591 VP.n45 VP.n1 0.189894
R1592 VP.n49 VP.n1 0.189894
R1593 VDD1 VDD1.t3 76.829
R1594 VDD1.n1 VDD1.t4 76.7144
R1595 VDD1.n1 VDD1.n0 73.395
R1596 VDD1.n3 VDD1.n2 72.6692
R1597 VDD1.n3 VDD1.n1 51.9233
R1598 VDD1.n2 VDD1.t0 1.76038
R1599 VDD1.n2 VDD1.t1 1.76038
R1600 VDD1.n0 VDD1.t5 1.76038
R1601 VDD1.n0 VDD1.t2 1.76038
R1602 VDD1 VDD1.n3 0.722483
C0 VDD2 VDD1 1.676f
C1 VTAIL VDD2 10.144401f
C2 VDD2 VP 0.51715f
C3 VDD2 w_n3866_n4662# 3.00847f
C4 VN B 1.38879f
C5 VN VDD1 0.151579f
C6 VN VTAIL 10.5898f
C7 VDD1 B 2.79178f
C8 VTAIL B 5.46906f
C9 VN VP 8.79427f
C10 B VP 2.22997f
C11 VN w_n3866_n4662# 7.60994f
C12 w_n3866_n4662# B 12.443001f
C13 VTAIL VDD1 10.089499f
C14 VDD1 VP 10.927f
C15 VN VDD2 10.5655f
C16 VTAIL VP 10.604099f
C17 w_n3866_n4662# VDD1 2.90135f
C18 VDD2 B 2.88242f
C19 VTAIL w_n3866_n4662# 3.91354f
C20 w_n3866_n4662# VP 8.11168f
C21 VDD2 VSUBS 2.23339f
C22 VDD1 VSUBS 2.78432f
C23 VTAIL VSUBS 1.558629f
C24 VN VSUBS 6.75575f
C25 VP VSUBS 3.713773f
C26 B VSUBS 5.865904f
C27 w_n3866_n4662# VSUBS 0.220316p
C28 VDD1.t3 VSUBS 4.33791f
C29 VDD1.t4 VSUBS 4.336451f
C30 VDD1.t5 VSUBS 0.39581f
C31 VDD1.t2 VSUBS 0.39581f
C32 VDD1.n0 VSUBS 3.33602f
C33 VDD1.n1 VSUBS 4.6587f
C34 VDD1.t0 VSUBS 0.39581f
C35 VDD1.t1 VSUBS 0.39581f
C36 VDD1.n2 VSUBS 3.32757f
C37 VDD1.n3 VSUBS 4.05013f
C38 VP.t3 VSUBS 4.27847f
C39 VP.n0 VSUBS 1.58216f
C40 VP.n1 VSUBS 0.025586f
C41 VP.n2 VSUBS 0.021892f
C42 VP.n3 VSUBS 0.025586f
C43 VP.t0 VSUBS 4.27847f
C44 VP.n4 VSUBS 1.47591f
C45 VP.n5 VSUBS 0.025586f
C46 VP.n6 VSUBS 0.021892f
C47 VP.n7 VSUBS 0.025586f
C48 VP.t1 VSUBS 4.27847f
C49 VP.n8 VSUBS 1.58216f
C50 VP.t4 VSUBS 4.27847f
C51 VP.n9 VSUBS 1.58216f
C52 VP.n10 VSUBS 0.025586f
C53 VP.n11 VSUBS 0.021892f
C54 VP.n12 VSUBS 0.025586f
C55 VP.t5 VSUBS 4.27847f
C56 VP.n13 VSUBS 1.56113f
C57 VP.t2 VSUBS 4.60638f
C58 VP.n14 VSUBS 1.49986f
C59 VP.n15 VSUBS 0.29854f
C60 VP.n16 VSUBS 0.035914f
C61 VP.n17 VSUBS 0.047685f
C62 VP.n18 VSUBS 0.0517f
C63 VP.n19 VSUBS 0.025586f
C64 VP.n20 VSUBS 0.025586f
C65 VP.n21 VSUBS 0.025586f
C66 VP.n22 VSUBS 0.048794f
C67 VP.n23 VSUBS 0.047685f
C68 VP.n24 VSUBS 0.041564f
C69 VP.n25 VSUBS 0.041294f
C70 VP.n26 VSUBS 1.72238f
C71 VP.n27 VSUBS 1.73867f
C72 VP.n28 VSUBS 0.041294f
C73 VP.n29 VSUBS 0.041564f
C74 VP.n30 VSUBS 0.047685f
C75 VP.n31 VSUBS 0.048794f
C76 VP.n32 VSUBS 0.025586f
C77 VP.n33 VSUBS 0.025586f
C78 VP.n34 VSUBS 0.025586f
C79 VP.n35 VSUBS 0.0517f
C80 VP.n36 VSUBS 0.047685f
C81 VP.n37 VSUBS 0.035914f
C82 VP.n38 VSUBS 0.025586f
C83 VP.n39 VSUBS 0.025586f
C84 VP.n40 VSUBS 0.035914f
C85 VP.n41 VSUBS 0.047685f
C86 VP.n42 VSUBS 0.0517f
C87 VP.n43 VSUBS 0.025586f
C88 VP.n44 VSUBS 0.025586f
C89 VP.n45 VSUBS 0.025586f
C90 VP.n46 VSUBS 0.048794f
C91 VP.n47 VSUBS 0.047685f
C92 VP.n48 VSUBS 0.041564f
C93 VP.n49 VSUBS 0.041294f
C94 VP.n50 VSUBS 0.058023f
C95 VDD2.t0 VSUBS 4.33647f
C96 VDD2.t2 VSUBS 0.395812f
C97 VDD2.t5 VSUBS 0.395812f
C98 VDD2.n0 VSUBS 3.33604f
C99 VDD2.n1 VSUBS 4.49901f
C100 VDD2.t1 VSUBS 4.31224f
C101 VDD2.n2 VSUBS 4.07836f
C102 VDD2.t3 VSUBS 0.395812f
C103 VDD2.t4 VSUBS 0.395812f
C104 VDD2.n3 VSUBS 3.33599f
C105 VTAIL.t11 VSUBS 0.406721f
C106 VTAIL.t7 VSUBS 0.406721f
C107 VTAIL.n0 VSUBS 3.2655f
C108 VTAIL.n1 VSUBS 0.895109f
C109 VTAIL.t1 VSUBS 4.25383f
C110 VTAIL.n2 VSUBS 1.22095f
C111 VTAIL.t2 VSUBS 0.406721f
C112 VTAIL.t4 VSUBS 0.406721f
C113 VTAIL.n3 VSUBS 3.2655f
C114 VTAIL.n4 VSUBS 3.28638f
C115 VTAIL.t9 VSUBS 0.406721f
C116 VTAIL.t8 VSUBS 0.406721f
C117 VTAIL.n5 VSUBS 3.26551f
C118 VTAIL.n6 VSUBS 3.28637f
C119 VTAIL.t6 VSUBS 4.25383f
C120 VTAIL.n7 VSUBS 1.22095f
C121 VTAIL.t3 VSUBS 0.406721f
C122 VTAIL.t0 VSUBS 0.406721f
C123 VTAIL.n8 VSUBS 3.26551f
C124 VTAIL.n9 VSUBS 1.10003f
C125 VTAIL.t5 VSUBS 4.25381f
C126 VTAIL.n10 VSUBS 3.1271f
C127 VTAIL.t10 VSUBS 4.25383f
C128 VTAIL.n11 VSUBS 3.05181f
C129 VN.t0 VSUBS 3.95882f
C130 VN.n0 VSUBS 1.46396f
C131 VN.n1 VSUBS 0.023674f
C132 VN.n2 VSUBS 0.020256f
C133 VN.n3 VSUBS 0.023674f
C134 VN.t3 VSUBS 3.95882f
C135 VN.n4 VSUBS 1.4445f
C136 VN.t5 VSUBS 4.26224f
C137 VN.n5 VSUBS 1.3878f
C138 VN.n6 VSUBS 0.276235f
C139 VN.n7 VSUBS 0.033231f
C140 VN.n8 VSUBS 0.044122f
C141 VN.n9 VSUBS 0.047838f
C142 VN.n10 VSUBS 0.023674f
C143 VN.n11 VSUBS 0.023674f
C144 VN.n12 VSUBS 0.023674f
C145 VN.n13 VSUBS 0.045148f
C146 VN.n14 VSUBS 0.044122f
C147 VN.n15 VSUBS 0.038459f
C148 VN.n16 VSUBS 0.038209f
C149 VN.n17 VSUBS 0.053688f
C150 VN.t4 VSUBS 3.95882f
C151 VN.n18 VSUBS 1.46396f
C152 VN.n19 VSUBS 0.023674f
C153 VN.n20 VSUBS 0.020256f
C154 VN.n21 VSUBS 0.023674f
C155 VN.t2 VSUBS 3.95882f
C156 VN.n22 VSUBS 1.4445f
C157 VN.t1 VSUBS 4.26224f
C158 VN.n23 VSUBS 1.3878f
C159 VN.n24 VSUBS 0.276235f
C160 VN.n25 VSUBS 0.033231f
C161 VN.n26 VSUBS 0.044122f
C162 VN.n27 VSUBS 0.047838f
C163 VN.n28 VSUBS 0.023674f
C164 VN.n29 VSUBS 0.023674f
C165 VN.n30 VSUBS 0.023674f
C166 VN.n31 VSUBS 0.045148f
C167 VN.n32 VSUBS 0.044122f
C168 VN.n33 VSUBS 0.038459f
C169 VN.n34 VSUBS 0.038209f
C170 VN.n35 VSUBS 1.60299f
C171 B.n0 VSUBS 0.006465f
C172 B.n1 VSUBS 0.006465f
C173 B.n2 VSUBS 0.009561f
C174 B.n3 VSUBS 0.007327f
C175 B.n4 VSUBS 0.007327f
C176 B.n5 VSUBS 0.007327f
C177 B.n6 VSUBS 0.007327f
C178 B.n7 VSUBS 0.007327f
C179 B.n8 VSUBS 0.007327f
C180 B.n9 VSUBS 0.007327f
C181 B.n10 VSUBS 0.007327f
C182 B.n11 VSUBS 0.007327f
C183 B.n12 VSUBS 0.007327f
C184 B.n13 VSUBS 0.007327f
C185 B.n14 VSUBS 0.007327f
C186 B.n15 VSUBS 0.007327f
C187 B.n16 VSUBS 0.007327f
C188 B.n17 VSUBS 0.007327f
C189 B.n18 VSUBS 0.007327f
C190 B.n19 VSUBS 0.007327f
C191 B.n20 VSUBS 0.007327f
C192 B.n21 VSUBS 0.007327f
C193 B.n22 VSUBS 0.007327f
C194 B.n23 VSUBS 0.007327f
C195 B.n24 VSUBS 0.007327f
C196 B.n25 VSUBS 0.007327f
C197 B.n26 VSUBS 0.007327f
C198 B.n27 VSUBS 0.018143f
C199 B.n28 VSUBS 0.007327f
C200 B.n29 VSUBS 0.007327f
C201 B.n30 VSUBS 0.007327f
C202 B.n31 VSUBS 0.007327f
C203 B.n32 VSUBS 0.007327f
C204 B.n33 VSUBS 0.007327f
C205 B.n34 VSUBS 0.007327f
C206 B.n35 VSUBS 0.007327f
C207 B.n36 VSUBS 0.007327f
C208 B.n37 VSUBS 0.007327f
C209 B.n38 VSUBS 0.007327f
C210 B.n39 VSUBS 0.007327f
C211 B.n40 VSUBS 0.007327f
C212 B.n41 VSUBS 0.007327f
C213 B.n42 VSUBS 0.007327f
C214 B.n43 VSUBS 0.007327f
C215 B.n44 VSUBS 0.007327f
C216 B.n45 VSUBS 0.007327f
C217 B.n46 VSUBS 0.007327f
C218 B.n47 VSUBS 0.007327f
C219 B.n48 VSUBS 0.007327f
C220 B.n49 VSUBS 0.007327f
C221 B.n50 VSUBS 0.007327f
C222 B.n51 VSUBS 0.007327f
C223 B.n52 VSUBS 0.007327f
C224 B.n53 VSUBS 0.007327f
C225 B.n54 VSUBS 0.007327f
C226 B.n55 VSUBS 0.007327f
C227 B.n56 VSUBS 0.007327f
C228 B.n57 VSUBS 0.007327f
C229 B.t7 VSUBS 0.653823f
C230 B.t8 VSUBS 0.680592f
C231 B.t6 VSUBS 2.8651f
C232 B.n58 VSUBS 0.407246f
C233 B.n59 VSUBS 0.078501f
C234 B.n60 VSUBS 0.007327f
C235 B.n61 VSUBS 0.007327f
C236 B.n62 VSUBS 0.007327f
C237 B.n63 VSUBS 0.007327f
C238 B.t4 VSUBS 0.653798f
C239 B.t5 VSUBS 0.680573f
C240 B.t3 VSUBS 2.8651f
C241 B.n64 VSUBS 0.407265f
C242 B.n65 VSUBS 0.078527f
C243 B.n66 VSUBS 0.016976f
C244 B.n67 VSUBS 0.007327f
C245 B.n68 VSUBS 0.007327f
C246 B.n69 VSUBS 0.007327f
C247 B.n70 VSUBS 0.007327f
C248 B.n71 VSUBS 0.007327f
C249 B.n72 VSUBS 0.007327f
C250 B.n73 VSUBS 0.007327f
C251 B.n74 VSUBS 0.007327f
C252 B.n75 VSUBS 0.007327f
C253 B.n76 VSUBS 0.007327f
C254 B.n77 VSUBS 0.007327f
C255 B.n78 VSUBS 0.007327f
C256 B.n79 VSUBS 0.007327f
C257 B.n80 VSUBS 0.007327f
C258 B.n81 VSUBS 0.007327f
C259 B.n82 VSUBS 0.007327f
C260 B.n83 VSUBS 0.007327f
C261 B.n84 VSUBS 0.007327f
C262 B.n85 VSUBS 0.007327f
C263 B.n86 VSUBS 0.007327f
C264 B.n87 VSUBS 0.007327f
C265 B.n88 VSUBS 0.007327f
C266 B.n89 VSUBS 0.007327f
C267 B.n90 VSUBS 0.007327f
C268 B.n91 VSUBS 0.007327f
C269 B.n92 VSUBS 0.007327f
C270 B.n93 VSUBS 0.007327f
C271 B.n94 VSUBS 0.007327f
C272 B.n95 VSUBS 0.007327f
C273 B.n96 VSUBS 0.007327f
C274 B.n97 VSUBS 0.016983f
C275 B.n98 VSUBS 0.007327f
C276 B.n99 VSUBS 0.007327f
C277 B.n100 VSUBS 0.007327f
C278 B.n101 VSUBS 0.007327f
C279 B.n102 VSUBS 0.007327f
C280 B.n103 VSUBS 0.007327f
C281 B.n104 VSUBS 0.007327f
C282 B.n105 VSUBS 0.007327f
C283 B.n106 VSUBS 0.007327f
C284 B.n107 VSUBS 0.007327f
C285 B.n108 VSUBS 0.007327f
C286 B.n109 VSUBS 0.007327f
C287 B.n110 VSUBS 0.007327f
C288 B.n111 VSUBS 0.007327f
C289 B.n112 VSUBS 0.007327f
C290 B.n113 VSUBS 0.007327f
C291 B.n114 VSUBS 0.007327f
C292 B.n115 VSUBS 0.007327f
C293 B.n116 VSUBS 0.007327f
C294 B.n117 VSUBS 0.007327f
C295 B.n118 VSUBS 0.007327f
C296 B.n119 VSUBS 0.007327f
C297 B.n120 VSUBS 0.007327f
C298 B.n121 VSUBS 0.007327f
C299 B.n122 VSUBS 0.007327f
C300 B.n123 VSUBS 0.007327f
C301 B.n124 VSUBS 0.007327f
C302 B.n125 VSUBS 0.007327f
C303 B.n126 VSUBS 0.007327f
C304 B.n127 VSUBS 0.007327f
C305 B.n128 VSUBS 0.007327f
C306 B.n129 VSUBS 0.007327f
C307 B.n130 VSUBS 0.007327f
C308 B.n131 VSUBS 0.007327f
C309 B.n132 VSUBS 0.007327f
C310 B.n133 VSUBS 0.007327f
C311 B.n134 VSUBS 0.007327f
C312 B.n135 VSUBS 0.007327f
C313 B.n136 VSUBS 0.007327f
C314 B.n137 VSUBS 0.007327f
C315 B.n138 VSUBS 0.007327f
C316 B.n139 VSUBS 0.007327f
C317 B.n140 VSUBS 0.007327f
C318 B.n141 VSUBS 0.007327f
C319 B.n142 VSUBS 0.007327f
C320 B.n143 VSUBS 0.007327f
C321 B.n144 VSUBS 0.007327f
C322 B.n145 VSUBS 0.007327f
C323 B.n146 VSUBS 0.007327f
C324 B.n147 VSUBS 0.007327f
C325 B.n148 VSUBS 0.017309f
C326 B.n149 VSUBS 0.007327f
C327 B.n150 VSUBS 0.007327f
C328 B.n151 VSUBS 0.007327f
C329 B.n152 VSUBS 0.007327f
C330 B.n153 VSUBS 0.007327f
C331 B.n154 VSUBS 0.007327f
C332 B.n155 VSUBS 0.007327f
C333 B.n156 VSUBS 0.007327f
C334 B.n157 VSUBS 0.007327f
C335 B.n158 VSUBS 0.007327f
C336 B.n159 VSUBS 0.007327f
C337 B.n160 VSUBS 0.007327f
C338 B.n161 VSUBS 0.007327f
C339 B.n162 VSUBS 0.007327f
C340 B.n163 VSUBS 0.007327f
C341 B.n164 VSUBS 0.007327f
C342 B.n165 VSUBS 0.007327f
C343 B.n166 VSUBS 0.007327f
C344 B.n167 VSUBS 0.007327f
C345 B.n168 VSUBS 0.007327f
C346 B.n169 VSUBS 0.007327f
C347 B.n170 VSUBS 0.007327f
C348 B.n171 VSUBS 0.007327f
C349 B.n172 VSUBS 0.007327f
C350 B.n173 VSUBS 0.007327f
C351 B.n174 VSUBS 0.007327f
C352 B.n175 VSUBS 0.007327f
C353 B.n176 VSUBS 0.007327f
C354 B.n177 VSUBS 0.007327f
C355 B.n178 VSUBS 0.005064f
C356 B.n179 VSUBS 0.007327f
C357 B.n180 VSUBS 0.007327f
C358 B.n181 VSUBS 0.007327f
C359 B.n182 VSUBS 0.007327f
C360 B.n183 VSUBS 0.007327f
C361 B.t11 VSUBS 0.653823f
C362 B.t10 VSUBS 0.680592f
C363 B.t9 VSUBS 2.8651f
C364 B.n184 VSUBS 0.407246f
C365 B.n185 VSUBS 0.078501f
C366 B.n186 VSUBS 0.007327f
C367 B.n187 VSUBS 0.007327f
C368 B.n188 VSUBS 0.007327f
C369 B.n189 VSUBS 0.007327f
C370 B.n190 VSUBS 0.007327f
C371 B.n191 VSUBS 0.007327f
C372 B.n192 VSUBS 0.007327f
C373 B.n193 VSUBS 0.007327f
C374 B.n194 VSUBS 0.007327f
C375 B.n195 VSUBS 0.007327f
C376 B.n196 VSUBS 0.007327f
C377 B.n197 VSUBS 0.007327f
C378 B.n198 VSUBS 0.007327f
C379 B.n199 VSUBS 0.007327f
C380 B.n200 VSUBS 0.007327f
C381 B.n201 VSUBS 0.007327f
C382 B.n202 VSUBS 0.007327f
C383 B.n203 VSUBS 0.007327f
C384 B.n204 VSUBS 0.007327f
C385 B.n205 VSUBS 0.007327f
C386 B.n206 VSUBS 0.007327f
C387 B.n207 VSUBS 0.007327f
C388 B.n208 VSUBS 0.007327f
C389 B.n209 VSUBS 0.007327f
C390 B.n210 VSUBS 0.007327f
C391 B.n211 VSUBS 0.007327f
C392 B.n212 VSUBS 0.007327f
C393 B.n213 VSUBS 0.007327f
C394 B.n214 VSUBS 0.007327f
C395 B.n215 VSUBS 0.018143f
C396 B.n216 VSUBS 0.007327f
C397 B.n217 VSUBS 0.007327f
C398 B.n218 VSUBS 0.007327f
C399 B.n219 VSUBS 0.007327f
C400 B.n220 VSUBS 0.007327f
C401 B.n221 VSUBS 0.007327f
C402 B.n222 VSUBS 0.007327f
C403 B.n223 VSUBS 0.007327f
C404 B.n224 VSUBS 0.007327f
C405 B.n225 VSUBS 0.007327f
C406 B.n226 VSUBS 0.007327f
C407 B.n227 VSUBS 0.007327f
C408 B.n228 VSUBS 0.007327f
C409 B.n229 VSUBS 0.007327f
C410 B.n230 VSUBS 0.007327f
C411 B.n231 VSUBS 0.007327f
C412 B.n232 VSUBS 0.007327f
C413 B.n233 VSUBS 0.007327f
C414 B.n234 VSUBS 0.007327f
C415 B.n235 VSUBS 0.007327f
C416 B.n236 VSUBS 0.007327f
C417 B.n237 VSUBS 0.007327f
C418 B.n238 VSUBS 0.007327f
C419 B.n239 VSUBS 0.007327f
C420 B.n240 VSUBS 0.007327f
C421 B.n241 VSUBS 0.007327f
C422 B.n242 VSUBS 0.007327f
C423 B.n243 VSUBS 0.007327f
C424 B.n244 VSUBS 0.007327f
C425 B.n245 VSUBS 0.007327f
C426 B.n246 VSUBS 0.007327f
C427 B.n247 VSUBS 0.007327f
C428 B.n248 VSUBS 0.007327f
C429 B.n249 VSUBS 0.007327f
C430 B.n250 VSUBS 0.007327f
C431 B.n251 VSUBS 0.007327f
C432 B.n252 VSUBS 0.007327f
C433 B.n253 VSUBS 0.007327f
C434 B.n254 VSUBS 0.007327f
C435 B.n255 VSUBS 0.007327f
C436 B.n256 VSUBS 0.007327f
C437 B.n257 VSUBS 0.007327f
C438 B.n258 VSUBS 0.007327f
C439 B.n259 VSUBS 0.007327f
C440 B.n260 VSUBS 0.007327f
C441 B.n261 VSUBS 0.007327f
C442 B.n262 VSUBS 0.007327f
C443 B.n263 VSUBS 0.007327f
C444 B.n264 VSUBS 0.007327f
C445 B.n265 VSUBS 0.007327f
C446 B.n266 VSUBS 0.007327f
C447 B.n267 VSUBS 0.007327f
C448 B.n268 VSUBS 0.007327f
C449 B.n269 VSUBS 0.007327f
C450 B.n270 VSUBS 0.007327f
C451 B.n271 VSUBS 0.007327f
C452 B.n272 VSUBS 0.007327f
C453 B.n273 VSUBS 0.007327f
C454 B.n274 VSUBS 0.007327f
C455 B.n275 VSUBS 0.007327f
C456 B.n276 VSUBS 0.007327f
C457 B.n277 VSUBS 0.007327f
C458 B.n278 VSUBS 0.007327f
C459 B.n279 VSUBS 0.007327f
C460 B.n280 VSUBS 0.007327f
C461 B.n281 VSUBS 0.007327f
C462 B.n282 VSUBS 0.007327f
C463 B.n283 VSUBS 0.007327f
C464 B.n284 VSUBS 0.007327f
C465 B.n285 VSUBS 0.007327f
C466 B.n286 VSUBS 0.007327f
C467 B.n287 VSUBS 0.007327f
C468 B.n288 VSUBS 0.007327f
C469 B.n289 VSUBS 0.007327f
C470 B.n290 VSUBS 0.007327f
C471 B.n291 VSUBS 0.007327f
C472 B.n292 VSUBS 0.007327f
C473 B.n293 VSUBS 0.007327f
C474 B.n294 VSUBS 0.007327f
C475 B.n295 VSUBS 0.007327f
C476 B.n296 VSUBS 0.007327f
C477 B.n297 VSUBS 0.007327f
C478 B.n298 VSUBS 0.007327f
C479 B.n299 VSUBS 0.007327f
C480 B.n300 VSUBS 0.007327f
C481 B.n301 VSUBS 0.007327f
C482 B.n302 VSUBS 0.007327f
C483 B.n303 VSUBS 0.007327f
C484 B.n304 VSUBS 0.007327f
C485 B.n305 VSUBS 0.007327f
C486 B.n306 VSUBS 0.007327f
C487 B.n307 VSUBS 0.007327f
C488 B.n308 VSUBS 0.007327f
C489 B.n309 VSUBS 0.007327f
C490 B.n310 VSUBS 0.007327f
C491 B.n311 VSUBS 0.007327f
C492 B.n312 VSUBS 0.016983f
C493 B.n313 VSUBS 0.016983f
C494 B.n314 VSUBS 0.018143f
C495 B.n315 VSUBS 0.007327f
C496 B.n316 VSUBS 0.007327f
C497 B.n317 VSUBS 0.007327f
C498 B.n318 VSUBS 0.007327f
C499 B.n319 VSUBS 0.007327f
C500 B.n320 VSUBS 0.007327f
C501 B.n321 VSUBS 0.007327f
C502 B.n322 VSUBS 0.007327f
C503 B.n323 VSUBS 0.007327f
C504 B.n324 VSUBS 0.007327f
C505 B.n325 VSUBS 0.007327f
C506 B.n326 VSUBS 0.007327f
C507 B.n327 VSUBS 0.007327f
C508 B.n328 VSUBS 0.007327f
C509 B.n329 VSUBS 0.007327f
C510 B.n330 VSUBS 0.007327f
C511 B.n331 VSUBS 0.007327f
C512 B.n332 VSUBS 0.007327f
C513 B.n333 VSUBS 0.007327f
C514 B.n334 VSUBS 0.007327f
C515 B.n335 VSUBS 0.007327f
C516 B.n336 VSUBS 0.007327f
C517 B.n337 VSUBS 0.007327f
C518 B.n338 VSUBS 0.007327f
C519 B.n339 VSUBS 0.007327f
C520 B.n340 VSUBS 0.007327f
C521 B.n341 VSUBS 0.007327f
C522 B.n342 VSUBS 0.007327f
C523 B.n343 VSUBS 0.007327f
C524 B.n344 VSUBS 0.007327f
C525 B.n345 VSUBS 0.007327f
C526 B.n346 VSUBS 0.007327f
C527 B.n347 VSUBS 0.007327f
C528 B.n348 VSUBS 0.007327f
C529 B.n349 VSUBS 0.007327f
C530 B.n350 VSUBS 0.007327f
C531 B.n351 VSUBS 0.007327f
C532 B.n352 VSUBS 0.007327f
C533 B.n353 VSUBS 0.007327f
C534 B.n354 VSUBS 0.007327f
C535 B.n355 VSUBS 0.007327f
C536 B.n356 VSUBS 0.007327f
C537 B.n357 VSUBS 0.007327f
C538 B.n358 VSUBS 0.007327f
C539 B.n359 VSUBS 0.007327f
C540 B.n360 VSUBS 0.007327f
C541 B.n361 VSUBS 0.007327f
C542 B.n362 VSUBS 0.007327f
C543 B.n363 VSUBS 0.007327f
C544 B.n364 VSUBS 0.007327f
C545 B.n365 VSUBS 0.007327f
C546 B.n366 VSUBS 0.007327f
C547 B.n367 VSUBS 0.007327f
C548 B.n368 VSUBS 0.007327f
C549 B.n369 VSUBS 0.007327f
C550 B.n370 VSUBS 0.007327f
C551 B.n371 VSUBS 0.007327f
C552 B.n372 VSUBS 0.007327f
C553 B.n373 VSUBS 0.007327f
C554 B.n374 VSUBS 0.007327f
C555 B.n375 VSUBS 0.007327f
C556 B.n376 VSUBS 0.007327f
C557 B.n377 VSUBS 0.007327f
C558 B.n378 VSUBS 0.007327f
C559 B.n379 VSUBS 0.007327f
C560 B.n380 VSUBS 0.007327f
C561 B.n381 VSUBS 0.007327f
C562 B.n382 VSUBS 0.007327f
C563 B.n383 VSUBS 0.007327f
C564 B.n384 VSUBS 0.007327f
C565 B.n385 VSUBS 0.007327f
C566 B.n386 VSUBS 0.007327f
C567 B.n387 VSUBS 0.007327f
C568 B.n388 VSUBS 0.007327f
C569 B.n389 VSUBS 0.007327f
C570 B.n390 VSUBS 0.007327f
C571 B.n391 VSUBS 0.007327f
C572 B.n392 VSUBS 0.007327f
C573 B.n393 VSUBS 0.007327f
C574 B.n394 VSUBS 0.007327f
C575 B.n395 VSUBS 0.007327f
C576 B.n396 VSUBS 0.007327f
C577 B.n397 VSUBS 0.007327f
C578 B.n398 VSUBS 0.007327f
C579 B.n399 VSUBS 0.007327f
C580 B.n400 VSUBS 0.007327f
C581 B.n401 VSUBS 0.007327f
C582 B.n402 VSUBS 0.007327f
C583 B.n403 VSUBS 0.007327f
C584 B.n404 VSUBS 0.005064f
C585 B.n405 VSUBS 0.016976f
C586 B.n406 VSUBS 0.005926f
C587 B.n407 VSUBS 0.007327f
C588 B.n408 VSUBS 0.007327f
C589 B.n409 VSUBS 0.007327f
C590 B.n410 VSUBS 0.007327f
C591 B.n411 VSUBS 0.007327f
C592 B.n412 VSUBS 0.007327f
C593 B.n413 VSUBS 0.007327f
C594 B.n414 VSUBS 0.007327f
C595 B.n415 VSUBS 0.007327f
C596 B.n416 VSUBS 0.007327f
C597 B.n417 VSUBS 0.007327f
C598 B.t2 VSUBS 0.653798f
C599 B.t1 VSUBS 0.680573f
C600 B.t0 VSUBS 2.8651f
C601 B.n418 VSUBS 0.407265f
C602 B.n419 VSUBS 0.078527f
C603 B.n420 VSUBS 0.016976f
C604 B.n421 VSUBS 0.005926f
C605 B.n422 VSUBS 0.007327f
C606 B.n423 VSUBS 0.007327f
C607 B.n424 VSUBS 0.007327f
C608 B.n425 VSUBS 0.007327f
C609 B.n426 VSUBS 0.007327f
C610 B.n427 VSUBS 0.007327f
C611 B.n428 VSUBS 0.007327f
C612 B.n429 VSUBS 0.007327f
C613 B.n430 VSUBS 0.007327f
C614 B.n431 VSUBS 0.007327f
C615 B.n432 VSUBS 0.007327f
C616 B.n433 VSUBS 0.007327f
C617 B.n434 VSUBS 0.007327f
C618 B.n435 VSUBS 0.007327f
C619 B.n436 VSUBS 0.007327f
C620 B.n437 VSUBS 0.007327f
C621 B.n438 VSUBS 0.007327f
C622 B.n439 VSUBS 0.007327f
C623 B.n440 VSUBS 0.007327f
C624 B.n441 VSUBS 0.007327f
C625 B.n442 VSUBS 0.007327f
C626 B.n443 VSUBS 0.007327f
C627 B.n444 VSUBS 0.007327f
C628 B.n445 VSUBS 0.007327f
C629 B.n446 VSUBS 0.007327f
C630 B.n447 VSUBS 0.007327f
C631 B.n448 VSUBS 0.007327f
C632 B.n449 VSUBS 0.007327f
C633 B.n450 VSUBS 0.007327f
C634 B.n451 VSUBS 0.007327f
C635 B.n452 VSUBS 0.007327f
C636 B.n453 VSUBS 0.007327f
C637 B.n454 VSUBS 0.007327f
C638 B.n455 VSUBS 0.007327f
C639 B.n456 VSUBS 0.007327f
C640 B.n457 VSUBS 0.007327f
C641 B.n458 VSUBS 0.007327f
C642 B.n459 VSUBS 0.007327f
C643 B.n460 VSUBS 0.007327f
C644 B.n461 VSUBS 0.007327f
C645 B.n462 VSUBS 0.007327f
C646 B.n463 VSUBS 0.007327f
C647 B.n464 VSUBS 0.007327f
C648 B.n465 VSUBS 0.007327f
C649 B.n466 VSUBS 0.007327f
C650 B.n467 VSUBS 0.007327f
C651 B.n468 VSUBS 0.007327f
C652 B.n469 VSUBS 0.007327f
C653 B.n470 VSUBS 0.007327f
C654 B.n471 VSUBS 0.007327f
C655 B.n472 VSUBS 0.007327f
C656 B.n473 VSUBS 0.007327f
C657 B.n474 VSUBS 0.007327f
C658 B.n475 VSUBS 0.007327f
C659 B.n476 VSUBS 0.007327f
C660 B.n477 VSUBS 0.007327f
C661 B.n478 VSUBS 0.007327f
C662 B.n479 VSUBS 0.007327f
C663 B.n480 VSUBS 0.007327f
C664 B.n481 VSUBS 0.007327f
C665 B.n482 VSUBS 0.007327f
C666 B.n483 VSUBS 0.007327f
C667 B.n484 VSUBS 0.007327f
C668 B.n485 VSUBS 0.007327f
C669 B.n486 VSUBS 0.007327f
C670 B.n487 VSUBS 0.007327f
C671 B.n488 VSUBS 0.007327f
C672 B.n489 VSUBS 0.007327f
C673 B.n490 VSUBS 0.007327f
C674 B.n491 VSUBS 0.007327f
C675 B.n492 VSUBS 0.007327f
C676 B.n493 VSUBS 0.007327f
C677 B.n494 VSUBS 0.007327f
C678 B.n495 VSUBS 0.007327f
C679 B.n496 VSUBS 0.007327f
C680 B.n497 VSUBS 0.007327f
C681 B.n498 VSUBS 0.007327f
C682 B.n499 VSUBS 0.007327f
C683 B.n500 VSUBS 0.007327f
C684 B.n501 VSUBS 0.007327f
C685 B.n502 VSUBS 0.007327f
C686 B.n503 VSUBS 0.007327f
C687 B.n504 VSUBS 0.007327f
C688 B.n505 VSUBS 0.007327f
C689 B.n506 VSUBS 0.007327f
C690 B.n507 VSUBS 0.007327f
C691 B.n508 VSUBS 0.007327f
C692 B.n509 VSUBS 0.007327f
C693 B.n510 VSUBS 0.007327f
C694 B.n511 VSUBS 0.007327f
C695 B.n512 VSUBS 0.007327f
C696 B.n513 VSUBS 0.018143f
C697 B.n514 VSUBS 0.016983f
C698 B.n515 VSUBS 0.017818f
C699 B.n516 VSUBS 0.007327f
C700 B.n517 VSUBS 0.007327f
C701 B.n518 VSUBS 0.007327f
C702 B.n519 VSUBS 0.007327f
C703 B.n520 VSUBS 0.007327f
C704 B.n521 VSUBS 0.007327f
C705 B.n522 VSUBS 0.007327f
C706 B.n523 VSUBS 0.007327f
C707 B.n524 VSUBS 0.007327f
C708 B.n525 VSUBS 0.007327f
C709 B.n526 VSUBS 0.007327f
C710 B.n527 VSUBS 0.007327f
C711 B.n528 VSUBS 0.007327f
C712 B.n529 VSUBS 0.007327f
C713 B.n530 VSUBS 0.007327f
C714 B.n531 VSUBS 0.007327f
C715 B.n532 VSUBS 0.007327f
C716 B.n533 VSUBS 0.007327f
C717 B.n534 VSUBS 0.007327f
C718 B.n535 VSUBS 0.007327f
C719 B.n536 VSUBS 0.007327f
C720 B.n537 VSUBS 0.007327f
C721 B.n538 VSUBS 0.007327f
C722 B.n539 VSUBS 0.007327f
C723 B.n540 VSUBS 0.007327f
C724 B.n541 VSUBS 0.007327f
C725 B.n542 VSUBS 0.007327f
C726 B.n543 VSUBS 0.007327f
C727 B.n544 VSUBS 0.007327f
C728 B.n545 VSUBS 0.007327f
C729 B.n546 VSUBS 0.007327f
C730 B.n547 VSUBS 0.007327f
C731 B.n548 VSUBS 0.007327f
C732 B.n549 VSUBS 0.007327f
C733 B.n550 VSUBS 0.007327f
C734 B.n551 VSUBS 0.007327f
C735 B.n552 VSUBS 0.007327f
C736 B.n553 VSUBS 0.007327f
C737 B.n554 VSUBS 0.007327f
C738 B.n555 VSUBS 0.007327f
C739 B.n556 VSUBS 0.007327f
C740 B.n557 VSUBS 0.007327f
C741 B.n558 VSUBS 0.007327f
C742 B.n559 VSUBS 0.007327f
C743 B.n560 VSUBS 0.007327f
C744 B.n561 VSUBS 0.007327f
C745 B.n562 VSUBS 0.007327f
C746 B.n563 VSUBS 0.007327f
C747 B.n564 VSUBS 0.007327f
C748 B.n565 VSUBS 0.007327f
C749 B.n566 VSUBS 0.007327f
C750 B.n567 VSUBS 0.007327f
C751 B.n568 VSUBS 0.007327f
C752 B.n569 VSUBS 0.007327f
C753 B.n570 VSUBS 0.007327f
C754 B.n571 VSUBS 0.007327f
C755 B.n572 VSUBS 0.007327f
C756 B.n573 VSUBS 0.007327f
C757 B.n574 VSUBS 0.007327f
C758 B.n575 VSUBS 0.007327f
C759 B.n576 VSUBS 0.007327f
C760 B.n577 VSUBS 0.007327f
C761 B.n578 VSUBS 0.007327f
C762 B.n579 VSUBS 0.007327f
C763 B.n580 VSUBS 0.007327f
C764 B.n581 VSUBS 0.007327f
C765 B.n582 VSUBS 0.007327f
C766 B.n583 VSUBS 0.007327f
C767 B.n584 VSUBS 0.007327f
C768 B.n585 VSUBS 0.007327f
C769 B.n586 VSUBS 0.007327f
C770 B.n587 VSUBS 0.007327f
C771 B.n588 VSUBS 0.007327f
C772 B.n589 VSUBS 0.007327f
C773 B.n590 VSUBS 0.007327f
C774 B.n591 VSUBS 0.007327f
C775 B.n592 VSUBS 0.007327f
C776 B.n593 VSUBS 0.007327f
C777 B.n594 VSUBS 0.007327f
C778 B.n595 VSUBS 0.007327f
C779 B.n596 VSUBS 0.007327f
C780 B.n597 VSUBS 0.007327f
C781 B.n598 VSUBS 0.007327f
C782 B.n599 VSUBS 0.007327f
C783 B.n600 VSUBS 0.007327f
C784 B.n601 VSUBS 0.007327f
C785 B.n602 VSUBS 0.007327f
C786 B.n603 VSUBS 0.007327f
C787 B.n604 VSUBS 0.007327f
C788 B.n605 VSUBS 0.007327f
C789 B.n606 VSUBS 0.007327f
C790 B.n607 VSUBS 0.007327f
C791 B.n608 VSUBS 0.007327f
C792 B.n609 VSUBS 0.007327f
C793 B.n610 VSUBS 0.007327f
C794 B.n611 VSUBS 0.007327f
C795 B.n612 VSUBS 0.007327f
C796 B.n613 VSUBS 0.007327f
C797 B.n614 VSUBS 0.007327f
C798 B.n615 VSUBS 0.007327f
C799 B.n616 VSUBS 0.007327f
C800 B.n617 VSUBS 0.007327f
C801 B.n618 VSUBS 0.007327f
C802 B.n619 VSUBS 0.007327f
C803 B.n620 VSUBS 0.007327f
C804 B.n621 VSUBS 0.007327f
C805 B.n622 VSUBS 0.007327f
C806 B.n623 VSUBS 0.007327f
C807 B.n624 VSUBS 0.007327f
C808 B.n625 VSUBS 0.007327f
C809 B.n626 VSUBS 0.007327f
C810 B.n627 VSUBS 0.007327f
C811 B.n628 VSUBS 0.007327f
C812 B.n629 VSUBS 0.007327f
C813 B.n630 VSUBS 0.007327f
C814 B.n631 VSUBS 0.007327f
C815 B.n632 VSUBS 0.007327f
C816 B.n633 VSUBS 0.007327f
C817 B.n634 VSUBS 0.007327f
C818 B.n635 VSUBS 0.007327f
C819 B.n636 VSUBS 0.007327f
C820 B.n637 VSUBS 0.007327f
C821 B.n638 VSUBS 0.007327f
C822 B.n639 VSUBS 0.007327f
C823 B.n640 VSUBS 0.007327f
C824 B.n641 VSUBS 0.007327f
C825 B.n642 VSUBS 0.007327f
C826 B.n643 VSUBS 0.007327f
C827 B.n644 VSUBS 0.007327f
C828 B.n645 VSUBS 0.007327f
C829 B.n646 VSUBS 0.007327f
C830 B.n647 VSUBS 0.007327f
C831 B.n648 VSUBS 0.007327f
C832 B.n649 VSUBS 0.007327f
C833 B.n650 VSUBS 0.007327f
C834 B.n651 VSUBS 0.007327f
C835 B.n652 VSUBS 0.007327f
C836 B.n653 VSUBS 0.007327f
C837 B.n654 VSUBS 0.007327f
C838 B.n655 VSUBS 0.007327f
C839 B.n656 VSUBS 0.007327f
C840 B.n657 VSUBS 0.007327f
C841 B.n658 VSUBS 0.007327f
C842 B.n659 VSUBS 0.007327f
C843 B.n660 VSUBS 0.007327f
C844 B.n661 VSUBS 0.007327f
C845 B.n662 VSUBS 0.007327f
C846 B.n663 VSUBS 0.007327f
C847 B.n664 VSUBS 0.007327f
C848 B.n665 VSUBS 0.007327f
C849 B.n666 VSUBS 0.016983f
C850 B.n667 VSUBS 0.018143f
C851 B.n668 VSUBS 0.018143f
C852 B.n669 VSUBS 0.007327f
C853 B.n670 VSUBS 0.007327f
C854 B.n671 VSUBS 0.007327f
C855 B.n672 VSUBS 0.007327f
C856 B.n673 VSUBS 0.007327f
C857 B.n674 VSUBS 0.007327f
C858 B.n675 VSUBS 0.007327f
C859 B.n676 VSUBS 0.007327f
C860 B.n677 VSUBS 0.007327f
C861 B.n678 VSUBS 0.007327f
C862 B.n679 VSUBS 0.007327f
C863 B.n680 VSUBS 0.007327f
C864 B.n681 VSUBS 0.007327f
C865 B.n682 VSUBS 0.007327f
C866 B.n683 VSUBS 0.007327f
C867 B.n684 VSUBS 0.007327f
C868 B.n685 VSUBS 0.007327f
C869 B.n686 VSUBS 0.007327f
C870 B.n687 VSUBS 0.007327f
C871 B.n688 VSUBS 0.007327f
C872 B.n689 VSUBS 0.007327f
C873 B.n690 VSUBS 0.007327f
C874 B.n691 VSUBS 0.007327f
C875 B.n692 VSUBS 0.007327f
C876 B.n693 VSUBS 0.007327f
C877 B.n694 VSUBS 0.007327f
C878 B.n695 VSUBS 0.007327f
C879 B.n696 VSUBS 0.007327f
C880 B.n697 VSUBS 0.007327f
C881 B.n698 VSUBS 0.007327f
C882 B.n699 VSUBS 0.007327f
C883 B.n700 VSUBS 0.007327f
C884 B.n701 VSUBS 0.007327f
C885 B.n702 VSUBS 0.007327f
C886 B.n703 VSUBS 0.007327f
C887 B.n704 VSUBS 0.007327f
C888 B.n705 VSUBS 0.007327f
C889 B.n706 VSUBS 0.007327f
C890 B.n707 VSUBS 0.007327f
C891 B.n708 VSUBS 0.007327f
C892 B.n709 VSUBS 0.007327f
C893 B.n710 VSUBS 0.007327f
C894 B.n711 VSUBS 0.007327f
C895 B.n712 VSUBS 0.007327f
C896 B.n713 VSUBS 0.007327f
C897 B.n714 VSUBS 0.007327f
C898 B.n715 VSUBS 0.007327f
C899 B.n716 VSUBS 0.007327f
C900 B.n717 VSUBS 0.007327f
C901 B.n718 VSUBS 0.007327f
C902 B.n719 VSUBS 0.007327f
C903 B.n720 VSUBS 0.007327f
C904 B.n721 VSUBS 0.007327f
C905 B.n722 VSUBS 0.007327f
C906 B.n723 VSUBS 0.007327f
C907 B.n724 VSUBS 0.007327f
C908 B.n725 VSUBS 0.007327f
C909 B.n726 VSUBS 0.007327f
C910 B.n727 VSUBS 0.007327f
C911 B.n728 VSUBS 0.007327f
C912 B.n729 VSUBS 0.007327f
C913 B.n730 VSUBS 0.007327f
C914 B.n731 VSUBS 0.007327f
C915 B.n732 VSUBS 0.007327f
C916 B.n733 VSUBS 0.007327f
C917 B.n734 VSUBS 0.007327f
C918 B.n735 VSUBS 0.007327f
C919 B.n736 VSUBS 0.007327f
C920 B.n737 VSUBS 0.007327f
C921 B.n738 VSUBS 0.007327f
C922 B.n739 VSUBS 0.007327f
C923 B.n740 VSUBS 0.007327f
C924 B.n741 VSUBS 0.007327f
C925 B.n742 VSUBS 0.007327f
C926 B.n743 VSUBS 0.007327f
C927 B.n744 VSUBS 0.007327f
C928 B.n745 VSUBS 0.007327f
C929 B.n746 VSUBS 0.007327f
C930 B.n747 VSUBS 0.007327f
C931 B.n748 VSUBS 0.007327f
C932 B.n749 VSUBS 0.007327f
C933 B.n750 VSUBS 0.007327f
C934 B.n751 VSUBS 0.007327f
C935 B.n752 VSUBS 0.007327f
C936 B.n753 VSUBS 0.007327f
C937 B.n754 VSUBS 0.007327f
C938 B.n755 VSUBS 0.007327f
C939 B.n756 VSUBS 0.007327f
C940 B.n757 VSUBS 0.005064f
C941 B.n758 VSUBS 0.007327f
C942 B.n759 VSUBS 0.007327f
C943 B.n760 VSUBS 0.005926f
C944 B.n761 VSUBS 0.007327f
C945 B.n762 VSUBS 0.007327f
C946 B.n763 VSUBS 0.007327f
C947 B.n764 VSUBS 0.007327f
C948 B.n765 VSUBS 0.007327f
C949 B.n766 VSUBS 0.007327f
C950 B.n767 VSUBS 0.007327f
C951 B.n768 VSUBS 0.007327f
C952 B.n769 VSUBS 0.007327f
C953 B.n770 VSUBS 0.007327f
C954 B.n771 VSUBS 0.007327f
C955 B.n772 VSUBS 0.005926f
C956 B.n773 VSUBS 0.016976f
C957 B.n774 VSUBS 0.005064f
C958 B.n775 VSUBS 0.007327f
C959 B.n776 VSUBS 0.007327f
C960 B.n777 VSUBS 0.007327f
C961 B.n778 VSUBS 0.007327f
C962 B.n779 VSUBS 0.007327f
C963 B.n780 VSUBS 0.007327f
C964 B.n781 VSUBS 0.007327f
C965 B.n782 VSUBS 0.007327f
C966 B.n783 VSUBS 0.007327f
C967 B.n784 VSUBS 0.007327f
C968 B.n785 VSUBS 0.007327f
C969 B.n786 VSUBS 0.007327f
C970 B.n787 VSUBS 0.007327f
C971 B.n788 VSUBS 0.007327f
C972 B.n789 VSUBS 0.007327f
C973 B.n790 VSUBS 0.007327f
C974 B.n791 VSUBS 0.007327f
C975 B.n792 VSUBS 0.007327f
C976 B.n793 VSUBS 0.007327f
C977 B.n794 VSUBS 0.007327f
C978 B.n795 VSUBS 0.007327f
C979 B.n796 VSUBS 0.007327f
C980 B.n797 VSUBS 0.007327f
C981 B.n798 VSUBS 0.007327f
C982 B.n799 VSUBS 0.007327f
C983 B.n800 VSUBS 0.007327f
C984 B.n801 VSUBS 0.007327f
C985 B.n802 VSUBS 0.007327f
C986 B.n803 VSUBS 0.007327f
C987 B.n804 VSUBS 0.007327f
C988 B.n805 VSUBS 0.007327f
C989 B.n806 VSUBS 0.007327f
C990 B.n807 VSUBS 0.007327f
C991 B.n808 VSUBS 0.007327f
C992 B.n809 VSUBS 0.007327f
C993 B.n810 VSUBS 0.007327f
C994 B.n811 VSUBS 0.007327f
C995 B.n812 VSUBS 0.007327f
C996 B.n813 VSUBS 0.007327f
C997 B.n814 VSUBS 0.007327f
C998 B.n815 VSUBS 0.007327f
C999 B.n816 VSUBS 0.007327f
C1000 B.n817 VSUBS 0.007327f
C1001 B.n818 VSUBS 0.007327f
C1002 B.n819 VSUBS 0.007327f
C1003 B.n820 VSUBS 0.007327f
C1004 B.n821 VSUBS 0.007327f
C1005 B.n822 VSUBS 0.007327f
C1006 B.n823 VSUBS 0.007327f
C1007 B.n824 VSUBS 0.007327f
C1008 B.n825 VSUBS 0.007327f
C1009 B.n826 VSUBS 0.007327f
C1010 B.n827 VSUBS 0.007327f
C1011 B.n828 VSUBS 0.007327f
C1012 B.n829 VSUBS 0.007327f
C1013 B.n830 VSUBS 0.007327f
C1014 B.n831 VSUBS 0.007327f
C1015 B.n832 VSUBS 0.007327f
C1016 B.n833 VSUBS 0.007327f
C1017 B.n834 VSUBS 0.007327f
C1018 B.n835 VSUBS 0.007327f
C1019 B.n836 VSUBS 0.007327f
C1020 B.n837 VSUBS 0.007327f
C1021 B.n838 VSUBS 0.007327f
C1022 B.n839 VSUBS 0.007327f
C1023 B.n840 VSUBS 0.007327f
C1024 B.n841 VSUBS 0.007327f
C1025 B.n842 VSUBS 0.007327f
C1026 B.n843 VSUBS 0.007327f
C1027 B.n844 VSUBS 0.007327f
C1028 B.n845 VSUBS 0.007327f
C1029 B.n846 VSUBS 0.007327f
C1030 B.n847 VSUBS 0.007327f
C1031 B.n848 VSUBS 0.007327f
C1032 B.n849 VSUBS 0.007327f
C1033 B.n850 VSUBS 0.007327f
C1034 B.n851 VSUBS 0.007327f
C1035 B.n852 VSUBS 0.007327f
C1036 B.n853 VSUBS 0.007327f
C1037 B.n854 VSUBS 0.007327f
C1038 B.n855 VSUBS 0.007327f
C1039 B.n856 VSUBS 0.007327f
C1040 B.n857 VSUBS 0.007327f
C1041 B.n858 VSUBS 0.007327f
C1042 B.n859 VSUBS 0.007327f
C1043 B.n860 VSUBS 0.007327f
C1044 B.n861 VSUBS 0.007327f
C1045 B.n862 VSUBS 0.007327f
C1046 B.n863 VSUBS 0.007327f
C1047 B.n864 VSUBS 0.018143f
C1048 B.n865 VSUBS 0.016983f
C1049 B.n866 VSUBS 0.016983f
C1050 B.n867 VSUBS 0.007327f
C1051 B.n868 VSUBS 0.007327f
C1052 B.n869 VSUBS 0.007327f
C1053 B.n870 VSUBS 0.007327f
C1054 B.n871 VSUBS 0.007327f
C1055 B.n872 VSUBS 0.007327f
C1056 B.n873 VSUBS 0.007327f
C1057 B.n874 VSUBS 0.007327f
C1058 B.n875 VSUBS 0.007327f
C1059 B.n876 VSUBS 0.007327f
C1060 B.n877 VSUBS 0.007327f
C1061 B.n878 VSUBS 0.007327f
C1062 B.n879 VSUBS 0.007327f
C1063 B.n880 VSUBS 0.007327f
C1064 B.n881 VSUBS 0.007327f
C1065 B.n882 VSUBS 0.007327f
C1066 B.n883 VSUBS 0.007327f
C1067 B.n884 VSUBS 0.007327f
C1068 B.n885 VSUBS 0.007327f
C1069 B.n886 VSUBS 0.007327f
C1070 B.n887 VSUBS 0.007327f
C1071 B.n888 VSUBS 0.007327f
C1072 B.n889 VSUBS 0.007327f
C1073 B.n890 VSUBS 0.007327f
C1074 B.n891 VSUBS 0.007327f
C1075 B.n892 VSUBS 0.007327f
C1076 B.n893 VSUBS 0.007327f
C1077 B.n894 VSUBS 0.007327f
C1078 B.n895 VSUBS 0.007327f
C1079 B.n896 VSUBS 0.007327f
C1080 B.n897 VSUBS 0.007327f
C1081 B.n898 VSUBS 0.007327f
C1082 B.n899 VSUBS 0.007327f
C1083 B.n900 VSUBS 0.007327f
C1084 B.n901 VSUBS 0.007327f
C1085 B.n902 VSUBS 0.007327f
C1086 B.n903 VSUBS 0.007327f
C1087 B.n904 VSUBS 0.007327f
C1088 B.n905 VSUBS 0.007327f
C1089 B.n906 VSUBS 0.007327f
C1090 B.n907 VSUBS 0.007327f
C1091 B.n908 VSUBS 0.007327f
C1092 B.n909 VSUBS 0.007327f
C1093 B.n910 VSUBS 0.007327f
C1094 B.n911 VSUBS 0.007327f
C1095 B.n912 VSUBS 0.007327f
C1096 B.n913 VSUBS 0.007327f
C1097 B.n914 VSUBS 0.007327f
C1098 B.n915 VSUBS 0.007327f
C1099 B.n916 VSUBS 0.007327f
C1100 B.n917 VSUBS 0.007327f
C1101 B.n918 VSUBS 0.007327f
C1102 B.n919 VSUBS 0.007327f
C1103 B.n920 VSUBS 0.007327f
C1104 B.n921 VSUBS 0.007327f
C1105 B.n922 VSUBS 0.007327f
C1106 B.n923 VSUBS 0.007327f
C1107 B.n924 VSUBS 0.007327f
C1108 B.n925 VSUBS 0.007327f
C1109 B.n926 VSUBS 0.007327f
C1110 B.n927 VSUBS 0.007327f
C1111 B.n928 VSUBS 0.007327f
C1112 B.n929 VSUBS 0.007327f
C1113 B.n930 VSUBS 0.007327f
C1114 B.n931 VSUBS 0.007327f
C1115 B.n932 VSUBS 0.007327f
C1116 B.n933 VSUBS 0.007327f
C1117 B.n934 VSUBS 0.007327f
C1118 B.n935 VSUBS 0.007327f
C1119 B.n936 VSUBS 0.007327f
C1120 B.n937 VSUBS 0.007327f
C1121 B.n938 VSUBS 0.007327f
C1122 B.n939 VSUBS 0.009561f
C1123 B.n940 VSUBS 0.010185f
C1124 B.n941 VSUBS 0.020254f
.ends

