VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ibex_wrapper
  CLASS BLOCK ;
  FOREIGN ibex_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 800.000 ;
  PIN EXT_IRQ
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 246.200 600.000 246.800 ;
    END
  END EXT_IRQ
  PIN HADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 796.000 148.490 800.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 796.000 581.810 800.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 796.000 271.770 800.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 796.000 24.290 800.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 223.080 600.000 223.680 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 108.840 600.000 109.440 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 360.440 600.000 361.040 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 796.000 426.330 800.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 796.000 596.530 800.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 199.960 600.000 200.560 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 703.160 600.000 703.760 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 17.720 600.000 18.320 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 337.320 600.000 337.920 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 796.000 101.570 800.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 520.920 600.000 521.520 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 796.000 457.610 800.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 451.560 600.000 452.160 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 635.160 600.000 635.760 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 542.680 600.000 543.280 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 796.000 132.850 800.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 176.840 600.000 177.440 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 269.320 600.000 269.920 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 796.000 504.530 800.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 406.680 600.000 407.280 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.080 600.000 291.680 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 62.600 600.000 63.200 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 796.000 71.210 800.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 565.800 600.000 566.400 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 796.000 85.930 800.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 796.000 225.770 800.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 796.000 8.650 800.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 749.400 600.000 750.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 796.000 256.130 800.000 ;
    END
  END HREADY
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 314.200 600.000 314.800 ;
    END
  END HRESETn
  PIN HSIZE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 796.000 364.690 800.000 ;
    END
  END HSIZE[0]
  PIN HSIZE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END HSIZE[1]
  PIN HSIZE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END HSIZE[2]
  PIN HTRANS[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 796.000 411.610 800.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 796.000 318.690 800.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 428.440 600.000 429.040 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 131.960 600.000 132.560 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 796.000 55.570 800.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 796.000 380.330 800.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 680.040 600.000 680.640 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 39.480 600.000 40.080 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 796.000 178.850 800.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 85.720 600.000 86.320 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 796.000 334.330 800.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 658.280 600.000 658.880 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 796.000 349.050 800.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 796.000 488.890 800.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 796.000 441.970 800.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 796.000 473.250 800.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END HWRITE
  PIN IRQ[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END IRQ[0]
  PIN IRQ[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END IRQ[10]
  PIN IRQ[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END IRQ[11]
  PIN IRQ[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 796.000 39.930 800.000 ;
    END
  END IRQ[12]
  PIN IRQ[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END IRQ[13]
  PIN IRQ[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 153.720 600.000 154.320 ;
    END
  END IRQ[14]
  PIN IRQ[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 796.000 194.490 800.000 ;
    END
  END IRQ[1]
  PIN IRQ[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 796.000 241.410 800.000 ;
    END
  END IRQ[2]
  PIN IRQ[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 796.000 395.970 800.000 ;
    END
  END IRQ[3]
  PIN IRQ[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END IRQ[4]
  PIN IRQ[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END IRQ[5]
  PIN IRQ[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END IRQ[6]
  PIN IRQ[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 796.000 534.890 800.000 ;
    END
  END IRQ[7]
  PIN IRQ[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 796.000 550.530 800.000 ;
    END
  END IRQ[8]
  PIN IRQ[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END IRQ[9]
  PIN NMI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END NMI
  PIN SYSTICKCLKDIV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 612.040 600.000 612.640 ;
    END
  END SYSTICKCLKDIV[0]
  PIN SYSTICKCLKDIV[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END SYSTICKCLKDIV[10]
  PIN SYSTICKCLKDIV[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 772.520 600.000 773.120 ;
    END
  END SYSTICKCLKDIV[11]
  PIN SYSTICKCLKDIV[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 588.920 600.000 589.520 ;
    END
  END SYSTICKCLKDIV[12]
  PIN SYSTICKCLKDIV[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END SYSTICKCLKDIV[13]
  PIN SYSTICKCLKDIV[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 796.000 117.210 800.000 ;
    END
  END SYSTICKCLKDIV[14]
  PIN SYSTICKCLKDIV[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 796.000 519.250 800.000 ;
    END
  END SYSTICKCLKDIV[15]
  PIN SYSTICKCLKDIV[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END SYSTICKCLKDIV[16]
  PIN SYSTICKCLKDIV[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 796.000 287.410 800.000 ;
    END
  END SYSTICKCLKDIV[17]
  PIN SYSTICKCLKDIV[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END SYSTICKCLKDIV[18]
  PIN SYSTICKCLKDIV[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END SYSTICKCLKDIV[19]
  PIN SYSTICKCLKDIV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 474.680 600.000 475.280 ;
    END
  END SYSTICKCLKDIV[1]
  PIN SYSTICKCLKDIV[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END SYSTICKCLKDIV[20]
  PIN SYSTICKCLKDIV[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END SYSTICKCLKDIV[21]
  PIN SYSTICKCLKDIV[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 796.000 210.130 800.000 ;
    END
  END SYSTICKCLKDIV[22]
  PIN SYSTICKCLKDIV[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 383.560 600.000 384.160 ;
    END
  END SYSTICKCLKDIV[23]
  PIN SYSTICKCLKDIV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 497.800 600.000 498.400 ;
    END
  END SYSTICKCLKDIV[2]
  PIN SYSTICKCLKDIV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END SYSTICKCLKDIV[3]
  PIN SYSTICKCLKDIV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END SYSTICKCLKDIV[4]
  PIN SYSTICKCLKDIV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 726.280 600.000 726.880 ;
    END
  END SYSTICKCLKDIV[5]
  PIN SYSTICKCLKDIV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 796.000 163.210 800.000 ;
    END
  END SYSTICKCLKDIV[6]
  PIN SYSTICKCLKDIV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END SYSTICKCLKDIV[7]
  PIN SYSTICKCLKDIV[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 796.000 566.170 800.000 ;
    END
  END SYSTICKCLKDIV[8]
  PIN SYSTICKCLKDIV[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 796.000 303.050 800.000 ;
    END
  END SYSTICKCLKDIV[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 788.885 ;
      LAYER met1 ;
        RECT 2.830 10.640 596.550 789.040 ;
      LAYER met2 ;
        RECT 2.860 795.720 8.090 796.010 ;
        RECT 8.930 795.720 23.730 796.010 ;
        RECT 24.570 795.720 39.370 796.010 ;
        RECT 40.210 795.720 55.010 796.010 ;
        RECT 55.850 795.720 70.650 796.010 ;
        RECT 71.490 795.720 85.370 796.010 ;
        RECT 86.210 795.720 101.010 796.010 ;
        RECT 101.850 795.720 116.650 796.010 ;
        RECT 117.490 795.720 132.290 796.010 ;
        RECT 133.130 795.720 147.930 796.010 ;
        RECT 148.770 795.720 162.650 796.010 ;
        RECT 163.490 795.720 178.290 796.010 ;
        RECT 179.130 795.720 193.930 796.010 ;
        RECT 194.770 795.720 209.570 796.010 ;
        RECT 210.410 795.720 225.210 796.010 ;
        RECT 226.050 795.720 240.850 796.010 ;
        RECT 241.690 795.720 255.570 796.010 ;
        RECT 256.410 795.720 271.210 796.010 ;
        RECT 272.050 795.720 286.850 796.010 ;
        RECT 287.690 795.720 302.490 796.010 ;
        RECT 303.330 795.720 318.130 796.010 ;
        RECT 318.970 795.720 333.770 796.010 ;
        RECT 334.610 795.720 348.490 796.010 ;
        RECT 349.330 795.720 364.130 796.010 ;
        RECT 364.970 795.720 379.770 796.010 ;
        RECT 380.610 795.720 395.410 796.010 ;
        RECT 396.250 795.720 411.050 796.010 ;
        RECT 411.890 795.720 425.770 796.010 ;
        RECT 426.610 795.720 441.410 796.010 ;
        RECT 442.250 795.720 457.050 796.010 ;
        RECT 457.890 795.720 472.690 796.010 ;
        RECT 473.530 795.720 488.330 796.010 ;
        RECT 489.170 795.720 503.970 796.010 ;
        RECT 504.810 795.720 518.690 796.010 ;
        RECT 519.530 795.720 534.330 796.010 ;
        RECT 535.170 795.720 549.970 796.010 ;
        RECT 550.810 795.720 565.610 796.010 ;
        RECT 566.450 795.720 581.250 796.010 ;
        RECT 582.090 795.720 595.970 796.010 ;
        RECT 2.860 4.280 596.520 795.720 ;
        RECT 3.410 4.000 17.290 4.280 ;
        RECT 18.130 4.000 32.930 4.280 ;
        RECT 33.770 4.000 48.570 4.280 ;
        RECT 49.410 4.000 64.210 4.280 ;
        RECT 65.050 4.000 79.850 4.280 ;
        RECT 80.690 4.000 94.570 4.280 ;
        RECT 95.410 4.000 110.210 4.280 ;
        RECT 111.050 4.000 125.850 4.280 ;
        RECT 126.690 4.000 141.490 4.280 ;
        RECT 142.330 4.000 157.130 4.280 ;
        RECT 157.970 4.000 172.770 4.280 ;
        RECT 173.610 4.000 187.490 4.280 ;
        RECT 188.330 4.000 203.130 4.280 ;
        RECT 203.970 4.000 218.770 4.280 ;
        RECT 219.610 4.000 234.410 4.280 ;
        RECT 235.250 4.000 250.050 4.280 ;
        RECT 250.890 4.000 264.770 4.280 ;
        RECT 265.610 4.000 280.410 4.280 ;
        RECT 281.250 4.000 296.050 4.280 ;
        RECT 296.890 4.000 311.690 4.280 ;
        RECT 312.530 4.000 327.330 4.280 ;
        RECT 328.170 4.000 342.970 4.280 ;
        RECT 343.810 4.000 357.690 4.280 ;
        RECT 358.530 4.000 373.330 4.280 ;
        RECT 374.170 4.000 388.970 4.280 ;
        RECT 389.810 4.000 404.610 4.280 ;
        RECT 405.450 4.000 420.250 4.280 ;
        RECT 421.090 4.000 435.890 4.280 ;
        RECT 436.730 4.000 450.610 4.280 ;
        RECT 451.450 4.000 466.250 4.280 ;
        RECT 467.090 4.000 481.890 4.280 ;
        RECT 482.730 4.000 497.530 4.280 ;
        RECT 498.370 4.000 513.170 4.280 ;
        RECT 514.010 4.000 527.890 4.280 ;
        RECT 528.730 4.000 543.530 4.280 ;
        RECT 544.370 4.000 559.170 4.280 ;
        RECT 560.010 4.000 574.810 4.280 ;
        RECT 575.650 4.000 590.450 4.280 ;
        RECT 591.290 4.000 596.520 4.280 ;
      LAYER met3 ;
        RECT 3.990 781.680 596.000 788.965 ;
        RECT 4.400 780.280 596.000 781.680 ;
        RECT 3.990 773.520 596.000 780.280 ;
        RECT 3.990 772.120 595.600 773.520 ;
        RECT 3.990 759.920 596.000 772.120 ;
        RECT 4.400 758.520 596.000 759.920 ;
        RECT 3.990 750.400 596.000 758.520 ;
        RECT 3.990 749.000 595.600 750.400 ;
        RECT 3.990 736.800 596.000 749.000 ;
        RECT 4.400 735.400 596.000 736.800 ;
        RECT 3.990 727.280 596.000 735.400 ;
        RECT 3.990 725.880 595.600 727.280 ;
        RECT 3.990 713.680 596.000 725.880 ;
        RECT 4.400 712.280 596.000 713.680 ;
        RECT 3.990 704.160 596.000 712.280 ;
        RECT 3.990 702.760 595.600 704.160 ;
        RECT 3.990 690.560 596.000 702.760 ;
        RECT 4.400 689.160 596.000 690.560 ;
        RECT 3.990 681.040 596.000 689.160 ;
        RECT 3.990 679.640 595.600 681.040 ;
        RECT 3.990 667.440 596.000 679.640 ;
        RECT 4.400 666.040 596.000 667.440 ;
        RECT 3.990 659.280 596.000 666.040 ;
        RECT 3.990 657.880 595.600 659.280 ;
        RECT 3.990 645.680 596.000 657.880 ;
        RECT 4.400 644.280 596.000 645.680 ;
        RECT 3.990 636.160 596.000 644.280 ;
        RECT 3.990 634.760 595.600 636.160 ;
        RECT 3.990 622.560 596.000 634.760 ;
        RECT 4.400 621.160 596.000 622.560 ;
        RECT 3.990 613.040 596.000 621.160 ;
        RECT 3.990 611.640 595.600 613.040 ;
        RECT 3.990 599.440 596.000 611.640 ;
        RECT 4.400 598.040 596.000 599.440 ;
        RECT 3.990 589.920 596.000 598.040 ;
        RECT 3.990 588.520 595.600 589.920 ;
        RECT 3.990 576.320 596.000 588.520 ;
        RECT 4.400 574.920 596.000 576.320 ;
        RECT 3.990 566.800 596.000 574.920 ;
        RECT 3.990 565.400 595.600 566.800 ;
        RECT 3.990 553.200 596.000 565.400 ;
        RECT 4.400 551.800 596.000 553.200 ;
        RECT 3.990 543.680 596.000 551.800 ;
        RECT 3.990 542.280 595.600 543.680 ;
        RECT 3.990 530.080 596.000 542.280 ;
        RECT 4.400 528.680 596.000 530.080 ;
        RECT 3.990 521.920 596.000 528.680 ;
        RECT 3.990 520.520 595.600 521.920 ;
        RECT 3.990 508.320 596.000 520.520 ;
        RECT 4.400 506.920 596.000 508.320 ;
        RECT 3.990 498.800 596.000 506.920 ;
        RECT 3.990 497.400 595.600 498.800 ;
        RECT 3.990 485.200 596.000 497.400 ;
        RECT 4.400 483.800 596.000 485.200 ;
        RECT 3.990 475.680 596.000 483.800 ;
        RECT 3.990 474.280 595.600 475.680 ;
        RECT 3.990 462.080 596.000 474.280 ;
        RECT 4.400 460.680 596.000 462.080 ;
        RECT 3.990 452.560 596.000 460.680 ;
        RECT 3.990 451.160 595.600 452.560 ;
        RECT 3.990 438.960 596.000 451.160 ;
        RECT 4.400 437.560 596.000 438.960 ;
        RECT 3.990 429.440 596.000 437.560 ;
        RECT 3.990 428.040 595.600 429.440 ;
        RECT 3.990 415.840 596.000 428.040 ;
        RECT 4.400 414.440 596.000 415.840 ;
        RECT 3.990 407.680 596.000 414.440 ;
        RECT 3.990 406.280 595.600 407.680 ;
        RECT 3.990 392.720 596.000 406.280 ;
        RECT 4.400 391.320 596.000 392.720 ;
        RECT 3.990 384.560 596.000 391.320 ;
        RECT 3.990 383.160 595.600 384.560 ;
        RECT 3.990 370.960 596.000 383.160 ;
        RECT 4.400 369.560 596.000 370.960 ;
        RECT 3.990 361.440 596.000 369.560 ;
        RECT 3.990 360.040 595.600 361.440 ;
        RECT 3.990 347.840 596.000 360.040 ;
        RECT 4.400 346.440 596.000 347.840 ;
        RECT 3.990 338.320 596.000 346.440 ;
        RECT 3.990 336.920 595.600 338.320 ;
        RECT 3.990 324.720 596.000 336.920 ;
        RECT 4.400 323.320 596.000 324.720 ;
        RECT 3.990 315.200 596.000 323.320 ;
        RECT 3.990 313.800 595.600 315.200 ;
        RECT 3.990 301.600 596.000 313.800 ;
        RECT 4.400 300.200 596.000 301.600 ;
        RECT 3.990 292.080 596.000 300.200 ;
        RECT 3.990 290.680 595.600 292.080 ;
        RECT 3.990 278.480 596.000 290.680 ;
        RECT 4.400 277.080 596.000 278.480 ;
        RECT 3.990 270.320 596.000 277.080 ;
        RECT 3.990 268.920 595.600 270.320 ;
        RECT 3.990 256.720 596.000 268.920 ;
        RECT 4.400 255.320 596.000 256.720 ;
        RECT 3.990 247.200 596.000 255.320 ;
        RECT 3.990 245.800 595.600 247.200 ;
        RECT 3.990 233.600 596.000 245.800 ;
        RECT 4.400 232.200 596.000 233.600 ;
        RECT 3.990 224.080 596.000 232.200 ;
        RECT 3.990 222.680 595.600 224.080 ;
        RECT 3.990 210.480 596.000 222.680 ;
        RECT 4.400 209.080 596.000 210.480 ;
        RECT 3.990 200.960 596.000 209.080 ;
        RECT 3.990 199.560 595.600 200.960 ;
        RECT 3.990 187.360 596.000 199.560 ;
        RECT 4.400 185.960 596.000 187.360 ;
        RECT 3.990 177.840 596.000 185.960 ;
        RECT 3.990 176.440 595.600 177.840 ;
        RECT 3.990 164.240 596.000 176.440 ;
        RECT 4.400 162.840 596.000 164.240 ;
        RECT 3.990 154.720 596.000 162.840 ;
        RECT 3.990 153.320 595.600 154.720 ;
        RECT 3.990 141.120 596.000 153.320 ;
        RECT 4.400 139.720 596.000 141.120 ;
        RECT 3.990 132.960 596.000 139.720 ;
        RECT 3.990 131.560 595.600 132.960 ;
        RECT 3.990 119.360 596.000 131.560 ;
        RECT 4.400 117.960 596.000 119.360 ;
        RECT 3.990 109.840 596.000 117.960 ;
        RECT 3.990 108.440 595.600 109.840 ;
        RECT 3.990 96.240 596.000 108.440 ;
        RECT 4.400 94.840 596.000 96.240 ;
        RECT 3.990 86.720 596.000 94.840 ;
        RECT 3.990 85.320 595.600 86.720 ;
        RECT 3.990 73.120 596.000 85.320 ;
        RECT 4.400 71.720 596.000 73.120 ;
        RECT 3.990 63.600 596.000 71.720 ;
        RECT 3.990 62.200 595.600 63.600 ;
        RECT 3.990 50.000 596.000 62.200 ;
        RECT 4.400 48.600 596.000 50.000 ;
        RECT 3.990 40.480 596.000 48.600 ;
        RECT 3.990 39.080 595.600 40.480 ;
        RECT 3.990 26.880 596.000 39.080 ;
        RECT 4.400 25.480 596.000 26.880 ;
        RECT 3.990 18.720 596.000 25.480 ;
        RECT 3.990 17.320 595.600 18.720 ;
        RECT 3.990 4.255 596.000 17.320 ;
      LAYER met4 ;
        RECT 13.175 12.415 20.640 787.265 ;
        RECT 23.040 12.415 97.440 787.265 ;
        RECT 99.840 12.415 174.240 787.265 ;
        RECT 176.640 12.415 251.040 787.265 ;
        RECT 253.440 12.415 327.840 787.265 ;
        RECT 330.240 12.415 404.640 787.265 ;
        RECT 407.040 12.415 481.440 787.265 ;
        RECT 483.840 12.415 558.240 787.265 ;
        RECT 560.640 12.415 586.665 787.265 ;
  END
END ibex_wrapper
END LIBRARY
