* NGSPICE file created from diff_pair_sample_0783.ext - technology: sky130A

.subckt diff_pair_sample_0783 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X1 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X2 VDD1.t6 VP.t1 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X3 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X4 VDD1.t5 VP.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=2.9562 ps=15.94 w=7.58 l=2.67
X5 VTAIL.t15 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X6 VTAIL.t7 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=1.2507 ps=7.91 w=7.58 l=2.67
X7 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=1.2507 ps=7.91 w=7.58 l=2.67
X8 VDD1.t3 VP.t4 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=2.9562 ps=15.94 w=7.58 l=2.67
X9 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=2.9562 ps=15.94 w=7.58 l=2.67
X10 VTAIL.t12 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=1.2507 ps=7.91 w=7.58 l=2.67
X11 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=2.9562 ps=15.94 w=7.58 l=2.67
X12 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=0 ps=0 w=7.58 l=2.67
X13 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X14 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=0 ps=0 w=7.58 l=2.67
X15 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X16 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=0 ps=0 w=7.58 l=2.67
X17 VTAIL.t14 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2507 pd=7.91 as=1.2507 ps=7.91 w=7.58 l=2.67
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=0 ps=0 w=7.58 l=2.67
X19 VTAIL.t9 VP.t7 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9562 pd=15.94 as=1.2507 ps=7.91 w=7.58 l=2.67
R0 VP.n18 VP.n17 161.3
R1 VP.n19 VP.n14 161.3
R2 VP.n21 VP.n20 161.3
R3 VP.n22 VP.n13 161.3
R4 VP.n24 VP.n23 161.3
R5 VP.n25 VP.n12 161.3
R6 VP.n27 VP.n26 161.3
R7 VP.n28 VP.n11 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n31 VP.n10 161.3
R10 VP.n33 VP.n32 161.3
R11 VP.n62 VP.n61 161.3
R12 VP.n60 VP.n1 161.3
R13 VP.n59 VP.n58 161.3
R14 VP.n57 VP.n2 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n54 VP.n3 161.3
R17 VP.n53 VP.n52 161.3
R18 VP.n51 VP.n4 161.3
R19 VP.n50 VP.n49 161.3
R20 VP.n48 VP.n5 161.3
R21 VP.n47 VP.n46 161.3
R22 VP.n45 VP.n6 161.3
R23 VP.n44 VP.n43 161.3
R24 VP.n42 VP.n7 161.3
R25 VP.n41 VP.n40 161.3
R26 VP.n39 VP.n8 161.3
R27 VP.n38 VP.n37 161.3
R28 VP.n16 VP.t7 100.642
R29 VP.n0 VP.t4 68.4192
R30 VP.n54 VP.t6 68.4192
R31 VP.n6 VP.t1 68.4192
R32 VP.n36 VP.t5 68.4192
R33 VP.n15 VP.t0 68.4192
R34 VP.n25 VP.t3 68.4192
R35 VP.n9 VP.t2 68.4192
R36 VP.n34 VP.n9 65.6537
R37 VP.n63 VP.n0 65.6537
R38 VP.n36 VP.n35 65.6537
R39 VP.n16 VP.n15 49.0352
R40 VP.n35 VP.n34 47.9844
R41 VP.n41 VP.n8 40.577
R42 VP.n42 VP.n41 40.577
R43 VP.n49 VP.n48 40.577
R44 VP.n49 VP.n4 40.577
R45 VP.n59 VP.n2 40.577
R46 VP.n60 VP.n59 40.577
R47 VP.n31 VP.n30 40.577
R48 VP.n30 VP.n11 40.577
R49 VP.n20 VP.n13 40.577
R50 VP.n20 VP.n19 40.577
R51 VP.n37 VP.n36 24.5923
R52 VP.n37 VP.n8 24.5923
R53 VP.n43 VP.n42 24.5923
R54 VP.n43 VP.n6 24.5923
R55 VP.n47 VP.n6 24.5923
R56 VP.n48 VP.n47 24.5923
R57 VP.n53 VP.n4 24.5923
R58 VP.n54 VP.n53 24.5923
R59 VP.n55 VP.n54 24.5923
R60 VP.n55 VP.n2 24.5923
R61 VP.n61 VP.n60 24.5923
R62 VP.n61 VP.n0 24.5923
R63 VP.n32 VP.n31 24.5923
R64 VP.n32 VP.n9 24.5923
R65 VP.n24 VP.n13 24.5923
R66 VP.n25 VP.n24 24.5923
R67 VP.n26 VP.n25 24.5923
R68 VP.n26 VP.n11 24.5923
R69 VP.n18 VP.n15 24.5923
R70 VP.n19 VP.n18 24.5923
R71 VP.n17 VP.n16 5.17217
R72 VP.n34 VP.n33 0.354861
R73 VP.n38 VP.n35 0.354861
R74 VP.n63 VP.n62 0.354861
R75 VP VP.n63 0.267071
R76 VP.n17 VP.n14 0.189894
R77 VP.n21 VP.n14 0.189894
R78 VP.n22 VP.n21 0.189894
R79 VP.n23 VP.n22 0.189894
R80 VP.n23 VP.n12 0.189894
R81 VP.n27 VP.n12 0.189894
R82 VP.n28 VP.n27 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n29 VP.n10 0.189894
R85 VP.n33 VP.n10 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n7 0.189894
R89 VP.n44 VP.n7 0.189894
R90 VP.n45 VP.n44 0.189894
R91 VP.n46 VP.n45 0.189894
R92 VP.n46 VP.n5 0.189894
R93 VP.n50 VP.n5 0.189894
R94 VP.n51 VP.n50 0.189894
R95 VP.n52 VP.n51 0.189894
R96 VP.n52 VP.n3 0.189894
R97 VP.n56 VP.n3 0.189894
R98 VP.n57 VP.n56 0.189894
R99 VP.n58 VP.n57 0.189894
R100 VP.n58 VP.n1 0.189894
R101 VP.n62 VP.n1 0.189894
R102 VTAIL.n11 VTAIL.t9 52.9398
R103 VTAIL.n10 VTAIL.t5 52.9398
R104 VTAIL.n7 VTAIL.t1 52.9398
R105 VTAIL.n15 VTAIL.t4 52.9396
R106 VTAIL.n2 VTAIL.t7 52.9396
R107 VTAIL.n3 VTAIL.t8 52.9396
R108 VTAIL.n6 VTAIL.t12 52.9396
R109 VTAIL.n14 VTAIL.t10 52.9396
R110 VTAIL.n13 VTAIL.n12 50.3276
R111 VTAIL.n9 VTAIL.n8 50.3276
R112 VTAIL.n1 VTAIL.n0 50.3274
R113 VTAIL.n5 VTAIL.n4 50.3274
R114 VTAIL.n15 VTAIL.n14 21.4876
R115 VTAIL.n7 VTAIL.n6 21.4876
R116 VTAIL.n0 VTAIL.t2 2.61264
R117 VTAIL.n0 VTAIL.t0 2.61264
R118 VTAIL.n4 VTAIL.t11 2.61264
R119 VTAIL.n4 VTAIL.t14 2.61264
R120 VTAIL.n12 VTAIL.t13 2.61264
R121 VTAIL.n12 VTAIL.t15 2.61264
R122 VTAIL.n8 VTAIL.t6 2.61264
R123 VTAIL.n8 VTAIL.t3 2.61264
R124 VTAIL.n9 VTAIL.n7 2.58671
R125 VTAIL.n10 VTAIL.n9 2.58671
R126 VTAIL.n13 VTAIL.n11 2.58671
R127 VTAIL.n14 VTAIL.n13 2.58671
R128 VTAIL.n6 VTAIL.n5 2.58671
R129 VTAIL.n5 VTAIL.n3 2.58671
R130 VTAIL.n2 VTAIL.n1 2.58671
R131 VTAIL VTAIL.n15 2.52852
R132 VTAIL.n11 VTAIL.n10 0.470328
R133 VTAIL.n3 VTAIL.n2 0.470328
R134 VTAIL VTAIL.n1 0.0586897
R135 VDD1 VDD1.n0 68.3577
R136 VDD1.n3 VDD1.n2 68.244
R137 VDD1.n3 VDD1.n1 68.244
R138 VDD1.n5 VDD1.n4 67.0062
R139 VDD1.n5 VDD1.n3 42.4707
R140 VDD1.n4 VDD1.t4 2.61264
R141 VDD1.n4 VDD1.t5 2.61264
R142 VDD1.n0 VDD1.t0 2.61264
R143 VDD1.n0 VDD1.t7 2.61264
R144 VDD1.n2 VDD1.t1 2.61264
R145 VDD1.n2 VDD1.t3 2.61264
R146 VDD1.n1 VDD1.t2 2.61264
R147 VDD1.n1 VDD1.t6 2.61264
R148 VDD1 VDD1.n5 1.23541
R149 B.n764 B.n763 585
R150 B.n765 B.n764 585
R151 B.n265 B.n130 585
R152 B.n264 B.n263 585
R153 B.n262 B.n261 585
R154 B.n260 B.n259 585
R155 B.n258 B.n257 585
R156 B.n256 B.n255 585
R157 B.n254 B.n253 585
R158 B.n252 B.n251 585
R159 B.n250 B.n249 585
R160 B.n248 B.n247 585
R161 B.n246 B.n245 585
R162 B.n244 B.n243 585
R163 B.n242 B.n241 585
R164 B.n240 B.n239 585
R165 B.n238 B.n237 585
R166 B.n236 B.n235 585
R167 B.n234 B.n233 585
R168 B.n232 B.n231 585
R169 B.n230 B.n229 585
R170 B.n228 B.n227 585
R171 B.n226 B.n225 585
R172 B.n224 B.n223 585
R173 B.n222 B.n221 585
R174 B.n220 B.n219 585
R175 B.n218 B.n217 585
R176 B.n216 B.n215 585
R177 B.n214 B.n213 585
R178 B.n212 B.n211 585
R179 B.n210 B.n209 585
R180 B.n208 B.n207 585
R181 B.n206 B.n205 585
R182 B.n204 B.n203 585
R183 B.n202 B.n201 585
R184 B.n200 B.n199 585
R185 B.n198 B.n197 585
R186 B.n196 B.n195 585
R187 B.n194 B.n193 585
R188 B.n191 B.n190 585
R189 B.n189 B.n188 585
R190 B.n187 B.n186 585
R191 B.n185 B.n184 585
R192 B.n183 B.n182 585
R193 B.n181 B.n180 585
R194 B.n179 B.n178 585
R195 B.n177 B.n176 585
R196 B.n175 B.n174 585
R197 B.n173 B.n172 585
R198 B.n171 B.n170 585
R199 B.n169 B.n168 585
R200 B.n167 B.n166 585
R201 B.n165 B.n164 585
R202 B.n163 B.n162 585
R203 B.n161 B.n160 585
R204 B.n159 B.n158 585
R205 B.n157 B.n156 585
R206 B.n155 B.n154 585
R207 B.n153 B.n152 585
R208 B.n151 B.n150 585
R209 B.n149 B.n148 585
R210 B.n147 B.n146 585
R211 B.n145 B.n144 585
R212 B.n143 B.n142 585
R213 B.n141 B.n140 585
R214 B.n139 B.n138 585
R215 B.n137 B.n136 585
R216 B.n95 B.n94 585
R217 B.n762 B.n96 585
R218 B.n766 B.n96 585
R219 B.n761 B.n760 585
R220 B.n760 B.n92 585
R221 B.n759 B.n91 585
R222 B.n772 B.n91 585
R223 B.n758 B.n90 585
R224 B.n773 B.n90 585
R225 B.n757 B.n89 585
R226 B.n774 B.n89 585
R227 B.n756 B.n755 585
R228 B.n755 B.n85 585
R229 B.n754 B.n84 585
R230 B.n780 B.n84 585
R231 B.n753 B.n83 585
R232 B.n781 B.n83 585
R233 B.n752 B.n82 585
R234 B.n782 B.n82 585
R235 B.n751 B.n750 585
R236 B.n750 B.n78 585
R237 B.n749 B.n77 585
R238 B.n788 B.n77 585
R239 B.n748 B.n76 585
R240 B.n789 B.n76 585
R241 B.n747 B.n75 585
R242 B.n790 B.n75 585
R243 B.n746 B.n745 585
R244 B.n745 B.n71 585
R245 B.n744 B.n70 585
R246 B.n796 B.n70 585
R247 B.n743 B.n69 585
R248 B.n797 B.n69 585
R249 B.n742 B.n68 585
R250 B.n798 B.n68 585
R251 B.n741 B.n740 585
R252 B.n740 B.n64 585
R253 B.n739 B.n63 585
R254 B.n804 B.n63 585
R255 B.n738 B.n62 585
R256 B.n805 B.n62 585
R257 B.n737 B.n61 585
R258 B.n806 B.n61 585
R259 B.n736 B.n735 585
R260 B.n735 B.n57 585
R261 B.n734 B.n56 585
R262 B.n812 B.n56 585
R263 B.n733 B.n55 585
R264 B.n813 B.n55 585
R265 B.n732 B.n54 585
R266 B.n814 B.n54 585
R267 B.n731 B.n730 585
R268 B.n730 B.n50 585
R269 B.n729 B.n49 585
R270 B.n820 B.n49 585
R271 B.n728 B.n48 585
R272 B.n821 B.n48 585
R273 B.n727 B.n47 585
R274 B.n822 B.n47 585
R275 B.n726 B.n725 585
R276 B.n725 B.n43 585
R277 B.n724 B.n42 585
R278 B.n828 B.n42 585
R279 B.n723 B.n41 585
R280 B.n829 B.n41 585
R281 B.n722 B.n40 585
R282 B.n830 B.n40 585
R283 B.n721 B.n720 585
R284 B.n720 B.n36 585
R285 B.n719 B.n35 585
R286 B.n836 B.n35 585
R287 B.n718 B.n34 585
R288 B.n837 B.n34 585
R289 B.n717 B.n33 585
R290 B.n838 B.n33 585
R291 B.n716 B.n715 585
R292 B.n715 B.n32 585
R293 B.n714 B.n28 585
R294 B.n844 B.n28 585
R295 B.n713 B.n27 585
R296 B.n845 B.n27 585
R297 B.n712 B.n26 585
R298 B.n846 B.n26 585
R299 B.n711 B.n710 585
R300 B.n710 B.n22 585
R301 B.n709 B.n21 585
R302 B.n852 B.n21 585
R303 B.n708 B.n20 585
R304 B.n853 B.n20 585
R305 B.n707 B.n19 585
R306 B.n854 B.n19 585
R307 B.n706 B.n705 585
R308 B.n705 B.n18 585
R309 B.n704 B.n14 585
R310 B.n860 B.n14 585
R311 B.n703 B.n13 585
R312 B.n861 B.n13 585
R313 B.n702 B.n12 585
R314 B.n862 B.n12 585
R315 B.n701 B.n700 585
R316 B.n700 B.n8 585
R317 B.n699 B.n7 585
R318 B.n868 B.n7 585
R319 B.n698 B.n6 585
R320 B.n869 B.n6 585
R321 B.n697 B.n5 585
R322 B.n870 B.n5 585
R323 B.n696 B.n695 585
R324 B.n695 B.n4 585
R325 B.n694 B.n266 585
R326 B.n694 B.n693 585
R327 B.n684 B.n267 585
R328 B.n268 B.n267 585
R329 B.n686 B.n685 585
R330 B.n687 B.n686 585
R331 B.n683 B.n273 585
R332 B.n273 B.n272 585
R333 B.n682 B.n681 585
R334 B.n681 B.n680 585
R335 B.n275 B.n274 585
R336 B.n673 B.n275 585
R337 B.n672 B.n671 585
R338 B.n674 B.n672 585
R339 B.n670 B.n280 585
R340 B.n280 B.n279 585
R341 B.n669 B.n668 585
R342 B.n668 B.n667 585
R343 B.n282 B.n281 585
R344 B.n283 B.n282 585
R345 B.n660 B.n659 585
R346 B.n661 B.n660 585
R347 B.n658 B.n288 585
R348 B.n288 B.n287 585
R349 B.n657 B.n656 585
R350 B.n656 B.n655 585
R351 B.n290 B.n289 585
R352 B.n648 B.n290 585
R353 B.n647 B.n646 585
R354 B.n649 B.n647 585
R355 B.n645 B.n295 585
R356 B.n295 B.n294 585
R357 B.n644 B.n643 585
R358 B.n643 B.n642 585
R359 B.n297 B.n296 585
R360 B.n298 B.n297 585
R361 B.n635 B.n634 585
R362 B.n636 B.n635 585
R363 B.n633 B.n303 585
R364 B.n303 B.n302 585
R365 B.n632 B.n631 585
R366 B.n631 B.n630 585
R367 B.n305 B.n304 585
R368 B.n306 B.n305 585
R369 B.n623 B.n622 585
R370 B.n624 B.n623 585
R371 B.n621 B.n311 585
R372 B.n311 B.n310 585
R373 B.n620 B.n619 585
R374 B.n619 B.n618 585
R375 B.n313 B.n312 585
R376 B.n314 B.n313 585
R377 B.n611 B.n610 585
R378 B.n612 B.n611 585
R379 B.n609 B.n319 585
R380 B.n319 B.n318 585
R381 B.n608 B.n607 585
R382 B.n607 B.n606 585
R383 B.n321 B.n320 585
R384 B.n322 B.n321 585
R385 B.n599 B.n598 585
R386 B.n600 B.n599 585
R387 B.n597 B.n326 585
R388 B.n330 B.n326 585
R389 B.n596 B.n595 585
R390 B.n595 B.n594 585
R391 B.n328 B.n327 585
R392 B.n329 B.n328 585
R393 B.n587 B.n586 585
R394 B.n588 B.n587 585
R395 B.n585 B.n335 585
R396 B.n335 B.n334 585
R397 B.n584 B.n583 585
R398 B.n583 B.n582 585
R399 B.n337 B.n336 585
R400 B.n338 B.n337 585
R401 B.n575 B.n574 585
R402 B.n576 B.n575 585
R403 B.n573 B.n343 585
R404 B.n343 B.n342 585
R405 B.n572 B.n571 585
R406 B.n571 B.n570 585
R407 B.n345 B.n344 585
R408 B.n346 B.n345 585
R409 B.n563 B.n562 585
R410 B.n564 B.n563 585
R411 B.n561 B.n350 585
R412 B.n354 B.n350 585
R413 B.n560 B.n559 585
R414 B.n559 B.n558 585
R415 B.n352 B.n351 585
R416 B.n353 B.n352 585
R417 B.n551 B.n550 585
R418 B.n552 B.n551 585
R419 B.n549 B.n359 585
R420 B.n359 B.n358 585
R421 B.n548 B.n547 585
R422 B.n547 B.n546 585
R423 B.n361 B.n360 585
R424 B.n362 B.n361 585
R425 B.n539 B.n538 585
R426 B.n540 B.n539 585
R427 B.n365 B.n364 585
R428 B.n407 B.n406 585
R429 B.n408 B.n404 585
R430 B.n404 B.n366 585
R431 B.n410 B.n409 585
R432 B.n412 B.n403 585
R433 B.n415 B.n414 585
R434 B.n416 B.n402 585
R435 B.n418 B.n417 585
R436 B.n420 B.n401 585
R437 B.n423 B.n422 585
R438 B.n424 B.n400 585
R439 B.n426 B.n425 585
R440 B.n428 B.n399 585
R441 B.n431 B.n430 585
R442 B.n432 B.n398 585
R443 B.n434 B.n433 585
R444 B.n436 B.n397 585
R445 B.n439 B.n438 585
R446 B.n440 B.n396 585
R447 B.n442 B.n441 585
R448 B.n444 B.n395 585
R449 B.n447 B.n446 585
R450 B.n448 B.n394 585
R451 B.n450 B.n449 585
R452 B.n452 B.n393 585
R453 B.n455 B.n454 585
R454 B.n456 B.n392 585
R455 B.n458 B.n457 585
R456 B.n460 B.n391 585
R457 B.n463 B.n462 585
R458 B.n464 B.n387 585
R459 B.n466 B.n465 585
R460 B.n468 B.n386 585
R461 B.n471 B.n470 585
R462 B.n472 B.n385 585
R463 B.n474 B.n473 585
R464 B.n476 B.n384 585
R465 B.n479 B.n478 585
R466 B.n481 B.n381 585
R467 B.n483 B.n482 585
R468 B.n485 B.n380 585
R469 B.n488 B.n487 585
R470 B.n489 B.n379 585
R471 B.n491 B.n490 585
R472 B.n493 B.n378 585
R473 B.n496 B.n495 585
R474 B.n497 B.n377 585
R475 B.n499 B.n498 585
R476 B.n501 B.n376 585
R477 B.n504 B.n503 585
R478 B.n505 B.n375 585
R479 B.n507 B.n506 585
R480 B.n509 B.n374 585
R481 B.n512 B.n511 585
R482 B.n513 B.n373 585
R483 B.n515 B.n514 585
R484 B.n517 B.n372 585
R485 B.n520 B.n519 585
R486 B.n521 B.n371 585
R487 B.n523 B.n522 585
R488 B.n525 B.n370 585
R489 B.n528 B.n527 585
R490 B.n529 B.n369 585
R491 B.n531 B.n530 585
R492 B.n533 B.n368 585
R493 B.n536 B.n535 585
R494 B.n537 B.n367 585
R495 B.n542 B.n541 585
R496 B.n541 B.n540 585
R497 B.n543 B.n363 585
R498 B.n363 B.n362 585
R499 B.n545 B.n544 585
R500 B.n546 B.n545 585
R501 B.n357 B.n356 585
R502 B.n358 B.n357 585
R503 B.n554 B.n553 585
R504 B.n553 B.n552 585
R505 B.n555 B.n355 585
R506 B.n355 B.n353 585
R507 B.n557 B.n556 585
R508 B.n558 B.n557 585
R509 B.n349 B.n348 585
R510 B.n354 B.n349 585
R511 B.n566 B.n565 585
R512 B.n565 B.n564 585
R513 B.n567 B.n347 585
R514 B.n347 B.n346 585
R515 B.n569 B.n568 585
R516 B.n570 B.n569 585
R517 B.n341 B.n340 585
R518 B.n342 B.n341 585
R519 B.n578 B.n577 585
R520 B.n577 B.n576 585
R521 B.n579 B.n339 585
R522 B.n339 B.n338 585
R523 B.n581 B.n580 585
R524 B.n582 B.n581 585
R525 B.n333 B.n332 585
R526 B.n334 B.n333 585
R527 B.n590 B.n589 585
R528 B.n589 B.n588 585
R529 B.n591 B.n331 585
R530 B.n331 B.n329 585
R531 B.n593 B.n592 585
R532 B.n594 B.n593 585
R533 B.n325 B.n324 585
R534 B.n330 B.n325 585
R535 B.n602 B.n601 585
R536 B.n601 B.n600 585
R537 B.n603 B.n323 585
R538 B.n323 B.n322 585
R539 B.n605 B.n604 585
R540 B.n606 B.n605 585
R541 B.n317 B.n316 585
R542 B.n318 B.n317 585
R543 B.n614 B.n613 585
R544 B.n613 B.n612 585
R545 B.n615 B.n315 585
R546 B.n315 B.n314 585
R547 B.n617 B.n616 585
R548 B.n618 B.n617 585
R549 B.n309 B.n308 585
R550 B.n310 B.n309 585
R551 B.n626 B.n625 585
R552 B.n625 B.n624 585
R553 B.n627 B.n307 585
R554 B.n307 B.n306 585
R555 B.n629 B.n628 585
R556 B.n630 B.n629 585
R557 B.n301 B.n300 585
R558 B.n302 B.n301 585
R559 B.n638 B.n637 585
R560 B.n637 B.n636 585
R561 B.n639 B.n299 585
R562 B.n299 B.n298 585
R563 B.n641 B.n640 585
R564 B.n642 B.n641 585
R565 B.n293 B.n292 585
R566 B.n294 B.n293 585
R567 B.n651 B.n650 585
R568 B.n650 B.n649 585
R569 B.n652 B.n291 585
R570 B.n648 B.n291 585
R571 B.n654 B.n653 585
R572 B.n655 B.n654 585
R573 B.n286 B.n285 585
R574 B.n287 B.n286 585
R575 B.n663 B.n662 585
R576 B.n662 B.n661 585
R577 B.n664 B.n284 585
R578 B.n284 B.n283 585
R579 B.n666 B.n665 585
R580 B.n667 B.n666 585
R581 B.n278 B.n277 585
R582 B.n279 B.n278 585
R583 B.n676 B.n675 585
R584 B.n675 B.n674 585
R585 B.n677 B.n276 585
R586 B.n673 B.n276 585
R587 B.n679 B.n678 585
R588 B.n680 B.n679 585
R589 B.n271 B.n270 585
R590 B.n272 B.n271 585
R591 B.n689 B.n688 585
R592 B.n688 B.n687 585
R593 B.n690 B.n269 585
R594 B.n269 B.n268 585
R595 B.n692 B.n691 585
R596 B.n693 B.n692 585
R597 B.n2 B.n0 585
R598 B.n4 B.n2 585
R599 B.n3 B.n1 585
R600 B.n869 B.n3 585
R601 B.n867 B.n866 585
R602 B.n868 B.n867 585
R603 B.n865 B.n9 585
R604 B.n9 B.n8 585
R605 B.n864 B.n863 585
R606 B.n863 B.n862 585
R607 B.n11 B.n10 585
R608 B.n861 B.n11 585
R609 B.n859 B.n858 585
R610 B.n860 B.n859 585
R611 B.n857 B.n15 585
R612 B.n18 B.n15 585
R613 B.n856 B.n855 585
R614 B.n855 B.n854 585
R615 B.n17 B.n16 585
R616 B.n853 B.n17 585
R617 B.n851 B.n850 585
R618 B.n852 B.n851 585
R619 B.n849 B.n23 585
R620 B.n23 B.n22 585
R621 B.n848 B.n847 585
R622 B.n847 B.n846 585
R623 B.n25 B.n24 585
R624 B.n845 B.n25 585
R625 B.n843 B.n842 585
R626 B.n844 B.n843 585
R627 B.n841 B.n29 585
R628 B.n32 B.n29 585
R629 B.n840 B.n839 585
R630 B.n839 B.n838 585
R631 B.n31 B.n30 585
R632 B.n837 B.n31 585
R633 B.n835 B.n834 585
R634 B.n836 B.n835 585
R635 B.n833 B.n37 585
R636 B.n37 B.n36 585
R637 B.n832 B.n831 585
R638 B.n831 B.n830 585
R639 B.n39 B.n38 585
R640 B.n829 B.n39 585
R641 B.n827 B.n826 585
R642 B.n828 B.n827 585
R643 B.n825 B.n44 585
R644 B.n44 B.n43 585
R645 B.n824 B.n823 585
R646 B.n823 B.n822 585
R647 B.n46 B.n45 585
R648 B.n821 B.n46 585
R649 B.n819 B.n818 585
R650 B.n820 B.n819 585
R651 B.n817 B.n51 585
R652 B.n51 B.n50 585
R653 B.n816 B.n815 585
R654 B.n815 B.n814 585
R655 B.n53 B.n52 585
R656 B.n813 B.n53 585
R657 B.n811 B.n810 585
R658 B.n812 B.n811 585
R659 B.n809 B.n58 585
R660 B.n58 B.n57 585
R661 B.n808 B.n807 585
R662 B.n807 B.n806 585
R663 B.n60 B.n59 585
R664 B.n805 B.n60 585
R665 B.n803 B.n802 585
R666 B.n804 B.n803 585
R667 B.n801 B.n65 585
R668 B.n65 B.n64 585
R669 B.n800 B.n799 585
R670 B.n799 B.n798 585
R671 B.n67 B.n66 585
R672 B.n797 B.n67 585
R673 B.n795 B.n794 585
R674 B.n796 B.n795 585
R675 B.n793 B.n72 585
R676 B.n72 B.n71 585
R677 B.n792 B.n791 585
R678 B.n791 B.n790 585
R679 B.n74 B.n73 585
R680 B.n789 B.n74 585
R681 B.n787 B.n786 585
R682 B.n788 B.n787 585
R683 B.n785 B.n79 585
R684 B.n79 B.n78 585
R685 B.n784 B.n783 585
R686 B.n783 B.n782 585
R687 B.n81 B.n80 585
R688 B.n781 B.n81 585
R689 B.n779 B.n778 585
R690 B.n780 B.n779 585
R691 B.n777 B.n86 585
R692 B.n86 B.n85 585
R693 B.n776 B.n775 585
R694 B.n775 B.n774 585
R695 B.n88 B.n87 585
R696 B.n773 B.n88 585
R697 B.n771 B.n770 585
R698 B.n772 B.n771 585
R699 B.n769 B.n93 585
R700 B.n93 B.n92 585
R701 B.n768 B.n767 585
R702 B.n767 B.n766 585
R703 B.n872 B.n871 585
R704 B.n871 B.n870 585
R705 B.n541 B.n365 521.33
R706 B.n767 B.n95 521.33
R707 B.n539 B.n367 521.33
R708 B.n764 B.n96 521.33
R709 B.n382 B.t8 276.57
R710 B.n388 B.t12 276.57
R711 B.n134 B.t19 276.57
R712 B.n131 B.t15 276.57
R713 B.n765 B.n129 256.663
R714 B.n765 B.n128 256.663
R715 B.n765 B.n127 256.663
R716 B.n765 B.n126 256.663
R717 B.n765 B.n125 256.663
R718 B.n765 B.n124 256.663
R719 B.n765 B.n123 256.663
R720 B.n765 B.n122 256.663
R721 B.n765 B.n121 256.663
R722 B.n765 B.n120 256.663
R723 B.n765 B.n119 256.663
R724 B.n765 B.n118 256.663
R725 B.n765 B.n117 256.663
R726 B.n765 B.n116 256.663
R727 B.n765 B.n115 256.663
R728 B.n765 B.n114 256.663
R729 B.n765 B.n113 256.663
R730 B.n765 B.n112 256.663
R731 B.n765 B.n111 256.663
R732 B.n765 B.n110 256.663
R733 B.n765 B.n109 256.663
R734 B.n765 B.n108 256.663
R735 B.n765 B.n107 256.663
R736 B.n765 B.n106 256.663
R737 B.n765 B.n105 256.663
R738 B.n765 B.n104 256.663
R739 B.n765 B.n103 256.663
R740 B.n765 B.n102 256.663
R741 B.n765 B.n101 256.663
R742 B.n765 B.n100 256.663
R743 B.n765 B.n99 256.663
R744 B.n765 B.n98 256.663
R745 B.n765 B.n97 256.663
R746 B.n405 B.n366 256.663
R747 B.n411 B.n366 256.663
R748 B.n413 B.n366 256.663
R749 B.n419 B.n366 256.663
R750 B.n421 B.n366 256.663
R751 B.n427 B.n366 256.663
R752 B.n429 B.n366 256.663
R753 B.n435 B.n366 256.663
R754 B.n437 B.n366 256.663
R755 B.n443 B.n366 256.663
R756 B.n445 B.n366 256.663
R757 B.n451 B.n366 256.663
R758 B.n453 B.n366 256.663
R759 B.n459 B.n366 256.663
R760 B.n461 B.n366 256.663
R761 B.n467 B.n366 256.663
R762 B.n469 B.n366 256.663
R763 B.n475 B.n366 256.663
R764 B.n477 B.n366 256.663
R765 B.n484 B.n366 256.663
R766 B.n486 B.n366 256.663
R767 B.n492 B.n366 256.663
R768 B.n494 B.n366 256.663
R769 B.n500 B.n366 256.663
R770 B.n502 B.n366 256.663
R771 B.n508 B.n366 256.663
R772 B.n510 B.n366 256.663
R773 B.n516 B.n366 256.663
R774 B.n518 B.n366 256.663
R775 B.n524 B.n366 256.663
R776 B.n526 B.n366 256.663
R777 B.n532 B.n366 256.663
R778 B.n534 B.n366 256.663
R779 B.n541 B.n363 163.367
R780 B.n545 B.n363 163.367
R781 B.n545 B.n357 163.367
R782 B.n553 B.n357 163.367
R783 B.n553 B.n355 163.367
R784 B.n557 B.n355 163.367
R785 B.n557 B.n349 163.367
R786 B.n565 B.n349 163.367
R787 B.n565 B.n347 163.367
R788 B.n569 B.n347 163.367
R789 B.n569 B.n341 163.367
R790 B.n577 B.n341 163.367
R791 B.n577 B.n339 163.367
R792 B.n581 B.n339 163.367
R793 B.n581 B.n333 163.367
R794 B.n589 B.n333 163.367
R795 B.n589 B.n331 163.367
R796 B.n593 B.n331 163.367
R797 B.n593 B.n325 163.367
R798 B.n601 B.n325 163.367
R799 B.n601 B.n323 163.367
R800 B.n605 B.n323 163.367
R801 B.n605 B.n317 163.367
R802 B.n613 B.n317 163.367
R803 B.n613 B.n315 163.367
R804 B.n617 B.n315 163.367
R805 B.n617 B.n309 163.367
R806 B.n625 B.n309 163.367
R807 B.n625 B.n307 163.367
R808 B.n629 B.n307 163.367
R809 B.n629 B.n301 163.367
R810 B.n637 B.n301 163.367
R811 B.n637 B.n299 163.367
R812 B.n641 B.n299 163.367
R813 B.n641 B.n293 163.367
R814 B.n650 B.n293 163.367
R815 B.n650 B.n291 163.367
R816 B.n654 B.n291 163.367
R817 B.n654 B.n286 163.367
R818 B.n662 B.n286 163.367
R819 B.n662 B.n284 163.367
R820 B.n666 B.n284 163.367
R821 B.n666 B.n278 163.367
R822 B.n675 B.n278 163.367
R823 B.n675 B.n276 163.367
R824 B.n679 B.n276 163.367
R825 B.n679 B.n271 163.367
R826 B.n688 B.n271 163.367
R827 B.n688 B.n269 163.367
R828 B.n692 B.n269 163.367
R829 B.n692 B.n2 163.367
R830 B.n871 B.n2 163.367
R831 B.n871 B.n3 163.367
R832 B.n867 B.n3 163.367
R833 B.n867 B.n9 163.367
R834 B.n863 B.n9 163.367
R835 B.n863 B.n11 163.367
R836 B.n859 B.n11 163.367
R837 B.n859 B.n15 163.367
R838 B.n855 B.n15 163.367
R839 B.n855 B.n17 163.367
R840 B.n851 B.n17 163.367
R841 B.n851 B.n23 163.367
R842 B.n847 B.n23 163.367
R843 B.n847 B.n25 163.367
R844 B.n843 B.n25 163.367
R845 B.n843 B.n29 163.367
R846 B.n839 B.n29 163.367
R847 B.n839 B.n31 163.367
R848 B.n835 B.n31 163.367
R849 B.n835 B.n37 163.367
R850 B.n831 B.n37 163.367
R851 B.n831 B.n39 163.367
R852 B.n827 B.n39 163.367
R853 B.n827 B.n44 163.367
R854 B.n823 B.n44 163.367
R855 B.n823 B.n46 163.367
R856 B.n819 B.n46 163.367
R857 B.n819 B.n51 163.367
R858 B.n815 B.n51 163.367
R859 B.n815 B.n53 163.367
R860 B.n811 B.n53 163.367
R861 B.n811 B.n58 163.367
R862 B.n807 B.n58 163.367
R863 B.n807 B.n60 163.367
R864 B.n803 B.n60 163.367
R865 B.n803 B.n65 163.367
R866 B.n799 B.n65 163.367
R867 B.n799 B.n67 163.367
R868 B.n795 B.n67 163.367
R869 B.n795 B.n72 163.367
R870 B.n791 B.n72 163.367
R871 B.n791 B.n74 163.367
R872 B.n787 B.n74 163.367
R873 B.n787 B.n79 163.367
R874 B.n783 B.n79 163.367
R875 B.n783 B.n81 163.367
R876 B.n779 B.n81 163.367
R877 B.n779 B.n86 163.367
R878 B.n775 B.n86 163.367
R879 B.n775 B.n88 163.367
R880 B.n771 B.n88 163.367
R881 B.n771 B.n93 163.367
R882 B.n767 B.n93 163.367
R883 B.n406 B.n404 163.367
R884 B.n410 B.n404 163.367
R885 B.n414 B.n412 163.367
R886 B.n418 B.n402 163.367
R887 B.n422 B.n420 163.367
R888 B.n426 B.n400 163.367
R889 B.n430 B.n428 163.367
R890 B.n434 B.n398 163.367
R891 B.n438 B.n436 163.367
R892 B.n442 B.n396 163.367
R893 B.n446 B.n444 163.367
R894 B.n450 B.n394 163.367
R895 B.n454 B.n452 163.367
R896 B.n458 B.n392 163.367
R897 B.n462 B.n460 163.367
R898 B.n466 B.n387 163.367
R899 B.n470 B.n468 163.367
R900 B.n474 B.n385 163.367
R901 B.n478 B.n476 163.367
R902 B.n483 B.n381 163.367
R903 B.n487 B.n485 163.367
R904 B.n491 B.n379 163.367
R905 B.n495 B.n493 163.367
R906 B.n499 B.n377 163.367
R907 B.n503 B.n501 163.367
R908 B.n507 B.n375 163.367
R909 B.n511 B.n509 163.367
R910 B.n515 B.n373 163.367
R911 B.n519 B.n517 163.367
R912 B.n523 B.n371 163.367
R913 B.n527 B.n525 163.367
R914 B.n531 B.n369 163.367
R915 B.n535 B.n533 163.367
R916 B.n539 B.n361 163.367
R917 B.n547 B.n361 163.367
R918 B.n547 B.n359 163.367
R919 B.n551 B.n359 163.367
R920 B.n551 B.n352 163.367
R921 B.n559 B.n352 163.367
R922 B.n559 B.n350 163.367
R923 B.n563 B.n350 163.367
R924 B.n563 B.n345 163.367
R925 B.n571 B.n345 163.367
R926 B.n571 B.n343 163.367
R927 B.n575 B.n343 163.367
R928 B.n575 B.n337 163.367
R929 B.n583 B.n337 163.367
R930 B.n583 B.n335 163.367
R931 B.n587 B.n335 163.367
R932 B.n587 B.n328 163.367
R933 B.n595 B.n328 163.367
R934 B.n595 B.n326 163.367
R935 B.n599 B.n326 163.367
R936 B.n599 B.n321 163.367
R937 B.n607 B.n321 163.367
R938 B.n607 B.n319 163.367
R939 B.n611 B.n319 163.367
R940 B.n611 B.n313 163.367
R941 B.n619 B.n313 163.367
R942 B.n619 B.n311 163.367
R943 B.n623 B.n311 163.367
R944 B.n623 B.n305 163.367
R945 B.n631 B.n305 163.367
R946 B.n631 B.n303 163.367
R947 B.n635 B.n303 163.367
R948 B.n635 B.n297 163.367
R949 B.n643 B.n297 163.367
R950 B.n643 B.n295 163.367
R951 B.n647 B.n295 163.367
R952 B.n647 B.n290 163.367
R953 B.n656 B.n290 163.367
R954 B.n656 B.n288 163.367
R955 B.n660 B.n288 163.367
R956 B.n660 B.n282 163.367
R957 B.n668 B.n282 163.367
R958 B.n668 B.n280 163.367
R959 B.n672 B.n280 163.367
R960 B.n672 B.n275 163.367
R961 B.n681 B.n275 163.367
R962 B.n681 B.n273 163.367
R963 B.n686 B.n273 163.367
R964 B.n686 B.n267 163.367
R965 B.n694 B.n267 163.367
R966 B.n695 B.n694 163.367
R967 B.n695 B.n5 163.367
R968 B.n6 B.n5 163.367
R969 B.n7 B.n6 163.367
R970 B.n700 B.n7 163.367
R971 B.n700 B.n12 163.367
R972 B.n13 B.n12 163.367
R973 B.n14 B.n13 163.367
R974 B.n705 B.n14 163.367
R975 B.n705 B.n19 163.367
R976 B.n20 B.n19 163.367
R977 B.n21 B.n20 163.367
R978 B.n710 B.n21 163.367
R979 B.n710 B.n26 163.367
R980 B.n27 B.n26 163.367
R981 B.n28 B.n27 163.367
R982 B.n715 B.n28 163.367
R983 B.n715 B.n33 163.367
R984 B.n34 B.n33 163.367
R985 B.n35 B.n34 163.367
R986 B.n720 B.n35 163.367
R987 B.n720 B.n40 163.367
R988 B.n41 B.n40 163.367
R989 B.n42 B.n41 163.367
R990 B.n725 B.n42 163.367
R991 B.n725 B.n47 163.367
R992 B.n48 B.n47 163.367
R993 B.n49 B.n48 163.367
R994 B.n730 B.n49 163.367
R995 B.n730 B.n54 163.367
R996 B.n55 B.n54 163.367
R997 B.n56 B.n55 163.367
R998 B.n735 B.n56 163.367
R999 B.n735 B.n61 163.367
R1000 B.n62 B.n61 163.367
R1001 B.n63 B.n62 163.367
R1002 B.n740 B.n63 163.367
R1003 B.n740 B.n68 163.367
R1004 B.n69 B.n68 163.367
R1005 B.n70 B.n69 163.367
R1006 B.n745 B.n70 163.367
R1007 B.n745 B.n75 163.367
R1008 B.n76 B.n75 163.367
R1009 B.n77 B.n76 163.367
R1010 B.n750 B.n77 163.367
R1011 B.n750 B.n82 163.367
R1012 B.n83 B.n82 163.367
R1013 B.n84 B.n83 163.367
R1014 B.n755 B.n84 163.367
R1015 B.n755 B.n89 163.367
R1016 B.n90 B.n89 163.367
R1017 B.n91 B.n90 163.367
R1018 B.n760 B.n91 163.367
R1019 B.n760 B.n96 163.367
R1020 B.n138 B.n137 163.367
R1021 B.n142 B.n141 163.367
R1022 B.n146 B.n145 163.367
R1023 B.n150 B.n149 163.367
R1024 B.n154 B.n153 163.367
R1025 B.n158 B.n157 163.367
R1026 B.n162 B.n161 163.367
R1027 B.n166 B.n165 163.367
R1028 B.n170 B.n169 163.367
R1029 B.n174 B.n173 163.367
R1030 B.n178 B.n177 163.367
R1031 B.n182 B.n181 163.367
R1032 B.n186 B.n185 163.367
R1033 B.n190 B.n189 163.367
R1034 B.n195 B.n194 163.367
R1035 B.n199 B.n198 163.367
R1036 B.n203 B.n202 163.367
R1037 B.n207 B.n206 163.367
R1038 B.n211 B.n210 163.367
R1039 B.n215 B.n214 163.367
R1040 B.n219 B.n218 163.367
R1041 B.n223 B.n222 163.367
R1042 B.n227 B.n226 163.367
R1043 B.n231 B.n230 163.367
R1044 B.n235 B.n234 163.367
R1045 B.n239 B.n238 163.367
R1046 B.n243 B.n242 163.367
R1047 B.n247 B.n246 163.367
R1048 B.n251 B.n250 163.367
R1049 B.n255 B.n254 163.367
R1050 B.n259 B.n258 163.367
R1051 B.n263 B.n262 163.367
R1052 B.n764 B.n130 163.367
R1053 B.n382 B.t11 128.869
R1054 B.n131 B.t17 128.869
R1055 B.n388 B.t14 128.859
R1056 B.n134 B.t20 128.859
R1057 B.n540 B.n366 118.942
R1058 B.n766 B.n765 118.942
R1059 B.n405 B.n365 71.676
R1060 B.n411 B.n410 71.676
R1061 B.n414 B.n413 71.676
R1062 B.n419 B.n418 71.676
R1063 B.n422 B.n421 71.676
R1064 B.n427 B.n426 71.676
R1065 B.n430 B.n429 71.676
R1066 B.n435 B.n434 71.676
R1067 B.n438 B.n437 71.676
R1068 B.n443 B.n442 71.676
R1069 B.n446 B.n445 71.676
R1070 B.n451 B.n450 71.676
R1071 B.n454 B.n453 71.676
R1072 B.n459 B.n458 71.676
R1073 B.n462 B.n461 71.676
R1074 B.n467 B.n466 71.676
R1075 B.n470 B.n469 71.676
R1076 B.n475 B.n474 71.676
R1077 B.n478 B.n477 71.676
R1078 B.n484 B.n483 71.676
R1079 B.n487 B.n486 71.676
R1080 B.n492 B.n491 71.676
R1081 B.n495 B.n494 71.676
R1082 B.n500 B.n499 71.676
R1083 B.n503 B.n502 71.676
R1084 B.n508 B.n507 71.676
R1085 B.n511 B.n510 71.676
R1086 B.n516 B.n515 71.676
R1087 B.n519 B.n518 71.676
R1088 B.n524 B.n523 71.676
R1089 B.n527 B.n526 71.676
R1090 B.n532 B.n531 71.676
R1091 B.n535 B.n534 71.676
R1092 B.n97 B.n95 71.676
R1093 B.n138 B.n98 71.676
R1094 B.n142 B.n99 71.676
R1095 B.n146 B.n100 71.676
R1096 B.n150 B.n101 71.676
R1097 B.n154 B.n102 71.676
R1098 B.n158 B.n103 71.676
R1099 B.n162 B.n104 71.676
R1100 B.n166 B.n105 71.676
R1101 B.n170 B.n106 71.676
R1102 B.n174 B.n107 71.676
R1103 B.n178 B.n108 71.676
R1104 B.n182 B.n109 71.676
R1105 B.n186 B.n110 71.676
R1106 B.n190 B.n111 71.676
R1107 B.n195 B.n112 71.676
R1108 B.n199 B.n113 71.676
R1109 B.n203 B.n114 71.676
R1110 B.n207 B.n115 71.676
R1111 B.n211 B.n116 71.676
R1112 B.n215 B.n117 71.676
R1113 B.n219 B.n118 71.676
R1114 B.n223 B.n119 71.676
R1115 B.n227 B.n120 71.676
R1116 B.n231 B.n121 71.676
R1117 B.n235 B.n122 71.676
R1118 B.n239 B.n123 71.676
R1119 B.n243 B.n124 71.676
R1120 B.n247 B.n125 71.676
R1121 B.n251 B.n126 71.676
R1122 B.n255 B.n127 71.676
R1123 B.n259 B.n128 71.676
R1124 B.n263 B.n129 71.676
R1125 B.n130 B.n129 71.676
R1126 B.n262 B.n128 71.676
R1127 B.n258 B.n127 71.676
R1128 B.n254 B.n126 71.676
R1129 B.n250 B.n125 71.676
R1130 B.n246 B.n124 71.676
R1131 B.n242 B.n123 71.676
R1132 B.n238 B.n122 71.676
R1133 B.n234 B.n121 71.676
R1134 B.n230 B.n120 71.676
R1135 B.n226 B.n119 71.676
R1136 B.n222 B.n118 71.676
R1137 B.n218 B.n117 71.676
R1138 B.n214 B.n116 71.676
R1139 B.n210 B.n115 71.676
R1140 B.n206 B.n114 71.676
R1141 B.n202 B.n113 71.676
R1142 B.n198 B.n112 71.676
R1143 B.n194 B.n111 71.676
R1144 B.n189 B.n110 71.676
R1145 B.n185 B.n109 71.676
R1146 B.n181 B.n108 71.676
R1147 B.n177 B.n107 71.676
R1148 B.n173 B.n106 71.676
R1149 B.n169 B.n105 71.676
R1150 B.n165 B.n104 71.676
R1151 B.n161 B.n103 71.676
R1152 B.n157 B.n102 71.676
R1153 B.n153 B.n101 71.676
R1154 B.n149 B.n100 71.676
R1155 B.n145 B.n99 71.676
R1156 B.n141 B.n98 71.676
R1157 B.n137 B.n97 71.676
R1158 B.n406 B.n405 71.676
R1159 B.n412 B.n411 71.676
R1160 B.n413 B.n402 71.676
R1161 B.n420 B.n419 71.676
R1162 B.n421 B.n400 71.676
R1163 B.n428 B.n427 71.676
R1164 B.n429 B.n398 71.676
R1165 B.n436 B.n435 71.676
R1166 B.n437 B.n396 71.676
R1167 B.n444 B.n443 71.676
R1168 B.n445 B.n394 71.676
R1169 B.n452 B.n451 71.676
R1170 B.n453 B.n392 71.676
R1171 B.n460 B.n459 71.676
R1172 B.n461 B.n387 71.676
R1173 B.n468 B.n467 71.676
R1174 B.n469 B.n385 71.676
R1175 B.n476 B.n475 71.676
R1176 B.n477 B.n381 71.676
R1177 B.n485 B.n484 71.676
R1178 B.n486 B.n379 71.676
R1179 B.n493 B.n492 71.676
R1180 B.n494 B.n377 71.676
R1181 B.n501 B.n500 71.676
R1182 B.n502 B.n375 71.676
R1183 B.n509 B.n508 71.676
R1184 B.n510 B.n373 71.676
R1185 B.n517 B.n516 71.676
R1186 B.n518 B.n371 71.676
R1187 B.n525 B.n524 71.676
R1188 B.n526 B.n369 71.676
R1189 B.n533 B.n532 71.676
R1190 B.n534 B.n367 71.676
R1191 B.n383 B.t10 70.6863
R1192 B.n132 B.t18 70.6863
R1193 B.n389 B.t13 70.6776
R1194 B.n135 B.t21 70.6776
R1195 B.n480 B.n383 59.5399
R1196 B.n390 B.n389 59.5399
R1197 B.n192 B.n135 59.5399
R1198 B.n133 B.n132 59.5399
R1199 B.n540 B.n362 58.188
R1200 B.n546 B.n362 58.188
R1201 B.n546 B.n358 58.188
R1202 B.n552 B.n358 58.188
R1203 B.n552 B.n353 58.188
R1204 B.n558 B.n353 58.188
R1205 B.n558 B.n354 58.188
R1206 B.n564 B.n346 58.188
R1207 B.n570 B.n346 58.188
R1208 B.n570 B.n342 58.188
R1209 B.n576 B.n342 58.188
R1210 B.n576 B.n338 58.188
R1211 B.n582 B.n338 58.188
R1212 B.n582 B.n334 58.188
R1213 B.n588 B.n334 58.188
R1214 B.n588 B.n329 58.188
R1215 B.n594 B.n329 58.188
R1216 B.n594 B.n330 58.188
R1217 B.n600 B.n322 58.188
R1218 B.n606 B.n322 58.188
R1219 B.n606 B.n318 58.188
R1220 B.n612 B.n318 58.188
R1221 B.n612 B.n314 58.188
R1222 B.n618 B.n314 58.188
R1223 B.n618 B.n310 58.188
R1224 B.n624 B.n310 58.188
R1225 B.n630 B.n306 58.188
R1226 B.n630 B.n302 58.188
R1227 B.n636 B.n302 58.188
R1228 B.n636 B.n298 58.188
R1229 B.n642 B.n298 58.188
R1230 B.n642 B.n294 58.188
R1231 B.n649 B.n294 58.188
R1232 B.n649 B.n648 58.188
R1233 B.n655 B.n287 58.188
R1234 B.n661 B.n287 58.188
R1235 B.n661 B.n283 58.188
R1236 B.n667 B.n283 58.188
R1237 B.n667 B.n279 58.188
R1238 B.n674 B.n279 58.188
R1239 B.n674 B.n673 58.188
R1240 B.n680 B.n272 58.188
R1241 B.n687 B.n272 58.188
R1242 B.n687 B.n268 58.188
R1243 B.n693 B.n268 58.188
R1244 B.n693 B.n4 58.188
R1245 B.n870 B.n4 58.188
R1246 B.n870 B.n869 58.188
R1247 B.n869 B.n868 58.188
R1248 B.n868 B.n8 58.188
R1249 B.n862 B.n8 58.188
R1250 B.n862 B.n861 58.188
R1251 B.n861 B.n860 58.188
R1252 B.n854 B.n18 58.188
R1253 B.n854 B.n853 58.188
R1254 B.n853 B.n852 58.188
R1255 B.n852 B.n22 58.188
R1256 B.n846 B.n22 58.188
R1257 B.n846 B.n845 58.188
R1258 B.n845 B.n844 58.188
R1259 B.n838 B.n32 58.188
R1260 B.n838 B.n837 58.188
R1261 B.n837 B.n836 58.188
R1262 B.n836 B.n36 58.188
R1263 B.n830 B.n36 58.188
R1264 B.n830 B.n829 58.188
R1265 B.n829 B.n828 58.188
R1266 B.n828 B.n43 58.188
R1267 B.n822 B.n821 58.188
R1268 B.n821 B.n820 58.188
R1269 B.n820 B.n50 58.188
R1270 B.n814 B.n50 58.188
R1271 B.n814 B.n813 58.188
R1272 B.n813 B.n812 58.188
R1273 B.n812 B.n57 58.188
R1274 B.n806 B.n57 58.188
R1275 B.n805 B.n804 58.188
R1276 B.n804 B.n64 58.188
R1277 B.n798 B.n64 58.188
R1278 B.n798 B.n797 58.188
R1279 B.n797 B.n796 58.188
R1280 B.n796 B.n71 58.188
R1281 B.n790 B.n71 58.188
R1282 B.n790 B.n789 58.188
R1283 B.n789 B.n788 58.188
R1284 B.n788 B.n78 58.188
R1285 B.n782 B.n78 58.188
R1286 B.n781 B.n780 58.188
R1287 B.n780 B.n85 58.188
R1288 B.n774 B.n85 58.188
R1289 B.n774 B.n773 58.188
R1290 B.n773 B.n772 58.188
R1291 B.n772 B.n92 58.188
R1292 B.n766 B.n92 58.188
R1293 B.n383 B.n382 58.1823
R1294 B.n389 B.n388 58.1823
R1295 B.n135 B.n134 58.1823
R1296 B.n132 B.n131 58.1823
R1297 B.n673 B.t5 57.3323
R1298 B.n18 B.t7 57.3323
R1299 B.n655 B.t3 48.7753
R1300 B.n844 B.t2 48.7753
R1301 B.t6 B.n306 38.5069
R1302 B.t0 B.n43 38.5069
R1303 B.n768 B.n94 33.8737
R1304 B.n763 B.n762 33.8737
R1305 B.n538 B.n537 33.8737
R1306 B.n542 B.n364 33.8737
R1307 B.n564 B.t9 29.9499
R1308 B.n330 B.t1 29.9499
R1309 B.t4 B.n805 29.9499
R1310 B.n782 B.t16 29.9499
R1311 B.n354 B.t9 28.2385
R1312 B.n600 B.t1 28.2385
R1313 B.n806 B.t4 28.2385
R1314 B.t16 B.n781 28.2385
R1315 B.n624 B.t6 19.6816
R1316 B.n822 B.t0 19.6816
R1317 B B.n872 18.0485
R1318 B.n136 B.n94 10.6151
R1319 B.n139 B.n136 10.6151
R1320 B.n140 B.n139 10.6151
R1321 B.n143 B.n140 10.6151
R1322 B.n144 B.n143 10.6151
R1323 B.n147 B.n144 10.6151
R1324 B.n148 B.n147 10.6151
R1325 B.n151 B.n148 10.6151
R1326 B.n152 B.n151 10.6151
R1327 B.n155 B.n152 10.6151
R1328 B.n156 B.n155 10.6151
R1329 B.n159 B.n156 10.6151
R1330 B.n160 B.n159 10.6151
R1331 B.n163 B.n160 10.6151
R1332 B.n164 B.n163 10.6151
R1333 B.n167 B.n164 10.6151
R1334 B.n168 B.n167 10.6151
R1335 B.n171 B.n168 10.6151
R1336 B.n172 B.n171 10.6151
R1337 B.n175 B.n172 10.6151
R1338 B.n176 B.n175 10.6151
R1339 B.n179 B.n176 10.6151
R1340 B.n180 B.n179 10.6151
R1341 B.n183 B.n180 10.6151
R1342 B.n184 B.n183 10.6151
R1343 B.n187 B.n184 10.6151
R1344 B.n188 B.n187 10.6151
R1345 B.n191 B.n188 10.6151
R1346 B.n196 B.n193 10.6151
R1347 B.n197 B.n196 10.6151
R1348 B.n200 B.n197 10.6151
R1349 B.n201 B.n200 10.6151
R1350 B.n204 B.n201 10.6151
R1351 B.n205 B.n204 10.6151
R1352 B.n208 B.n205 10.6151
R1353 B.n209 B.n208 10.6151
R1354 B.n213 B.n212 10.6151
R1355 B.n216 B.n213 10.6151
R1356 B.n217 B.n216 10.6151
R1357 B.n220 B.n217 10.6151
R1358 B.n221 B.n220 10.6151
R1359 B.n224 B.n221 10.6151
R1360 B.n225 B.n224 10.6151
R1361 B.n228 B.n225 10.6151
R1362 B.n229 B.n228 10.6151
R1363 B.n232 B.n229 10.6151
R1364 B.n233 B.n232 10.6151
R1365 B.n236 B.n233 10.6151
R1366 B.n237 B.n236 10.6151
R1367 B.n240 B.n237 10.6151
R1368 B.n241 B.n240 10.6151
R1369 B.n244 B.n241 10.6151
R1370 B.n245 B.n244 10.6151
R1371 B.n248 B.n245 10.6151
R1372 B.n249 B.n248 10.6151
R1373 B.n252 B.n249 10.6151
R1374 B.n253 B.n252 10.6151
R1375 B.n256 B.n253 10.6151
R1376 B.n257 B.n256 10.6151
R1377 B.n260 B.n257 10.6151
R1378 B.n261 B.n260 10.6151
R1379 B.n264 B.n261 10.6151
R1380 B.n265 B.n264 10.6151
R1381 B.n763 B.n265 10.6151
R1382 B.n538 B.n360 10.6151
R1383 B.n548 B.n360 10.6151
R1384 B.n549 B.n548 10.6151
R1385 B.n550 B.n549 10.6151
R1386 B.n550 B.n351 10.6151
R1387 B.n560 B.n351 10.6151
R1388 B.n561 B.n560 10.6151
R1389 B.n562 B.n561 10.6151
R1390 B.n562 B.n344 10.6151
R1391 B.n572 B.n344 10.6151
R1392 B.n573 B.n572 10.6151
R1393 B.n574 B.n573 10.6151
R1394 B.n574 B.n336 10.6151
R1395 B.n584 B.n336 10.6151
R1396 B.n585 B.n584 10.6151
R1397 B.n586 B.n585 10.6151
R1398 B.n586 B.n327 10.6151
R1399 B.n596 B.n327 10.6151
R1400 B.n597 B.n596 10.6151
R1401 B.n598 B.n597 10.6151
R1402 B.n598 B.n320 10.6151
R1403 B.n608 B.n320 10.6151
R1404 B.n609 B.n608 10.6151
R1405 B.n610 B.n609 10.6151
R1406 B.n610 B.n312 10.6151
R1407 B.n620 B.n312 10.6151
R1408 B.n621 B.n620 10.6151
R1409 B.n622 B.n621 10.6151
R1410 B.n622 B.n304 10.6151
R1411 B.n632 B.n304 10.6151
R1412 B.n633 B.n632 10.6151
R1413 B.n634 B.n633 10.6151
R1414 B.n634 B.n296 10.6151
R1415 B.n644 B.n296 10.6151
R1416 B.n645 B.n644 10.6151
R1417 B.n646 B.n645 10.6151
R1418 B.n646 B.n289 10.6151
R1419 B.n657 B.n289 10.6151
R1420 B.n658 B.n657 10.6151
R1421 B.n659 B.n658 10.6151
R1422 B.n659 B.n281 10.6151
R1423 B.n669 B.n281 10.6151
R1424 B.n670 B.n669 10.6151
R1425 B.n671 B.n670 10.6151
R1426 B.n671 B.n274 10.6151
R1427 B.n682 B.n274 10.6151
R1428 B.n683 B.n682 10.6151
R1429 B.n685 B.n683 10.6151
R1430 B.n685 B.n684 10.6151
R1431 B.n684 B.n266 10.6151
R1432 B.n696 B.n266 10.6151
R1433 B.n697 B.n696 10.6151
R1434 B.n698 B.n697 10.6151
R1435 B.n699 B.n698 10.6151
R1436 B.n701 B.n699 10.6151
R1437 B.n702 B.n701 10.6151
R1438 B.n703 B.n702 10.6151
R1439 B.n704 B.n703 10.6151
R1440 B.n706 B.n704 10.6151
R1441 B.n707 B.n706 10.6151
R1442 B.n708 B.n707 10.6151
R1443 B.n709 B.n708 10.6151
R1444 B.n711 B.n709 10.6151
R1445 B.n712 B.n711 10.6151
R1446 B.n713 B.n712 10.6151
R1447 B.n714 B.n713 10.6151
R1448 B.n716 B.n714 10.6151
R1449 B.n717 B.n716 10.6151
R1450 B.n718 B.n717 10.6151
R1451 B.n719 B.n718 10.6151
R1452 B.n721 B.n719 10.6151
R1453 B.n722 B.n721 10.6151
R1454 B.n723 B.n722 10.6151
R1455 B.n724 B.n723 10.6151
R1456 B.n726 B.n724 10.6151
R1457 B.n727 B.n726 10.6151
R1458 B.n728 B.n727 10.6151
R1459 B.n729 B.n728 10.6151
R1460 B.n731 B.n729 10.6151
R1461 B.n732 B.n731 10.6151
R1462 B.n733 B.n732 10.6151
R1463 B.n734 B.n733 10.6151
R1464 B.n736 B.n734 10.6151
R1465 B.n737 B.n736 10.6151
R1466 B.n738 B.n737 10.6151
R1467 B.n739 B.n738 10.6151
R1468 B.n741 B.n739 10.6151
R1469 B.n742 B.n741 10.6151
R1470 B.n743 B.n742 10.6151
R1471 B.n744 B.n743 10.6151
R1472 B.n746 B.n744 10.6151
R1473 B.n747 B.n746 10.6151
R1474 B.n748 B.n747 10.6151
R1475 B.n749 B.n748 10.6151
R1476 B.n751 B.n749 10.6151
R1477 B.n752 B.n751 10.6151
R1478 B.n753 B.n752 10.6151
R1479 B.n754 B.n753 10.6151
R1480 B.n756 B.n754 10.6151
R1481 B.n757 B.n756 10.6151
R1482 B.n758 B.n757 10.6151
R1483 B.n759 B.n758 10.6151
R1484 B.n761 B.n759 10.6151
R1485 B.n762 B.n761 10.6151
R1486 B.n407 B.n364 10.6151
R1487 B.n408 B.n407 10.6151
R1488 B.n409 B.n408 10.6151
R1489 B.n409 B.n403 10.6151
R1490 B.n415 B.n403 10.6151
R1491 B.n416 B.n415 10.6151
R1492 B.n417 B.n416 10.6151
R1493 B.n417 B.n401 10.6151
R1494 B.n423 B.n401 10.6151
R1495 B.n424 B.n423 10.6151
R1496 B.n425 B.n424 10.6151
R1497 B.n425 B.n399 10.6151
R1498 B.n431 B.n399 10.6151
R1499 B.n432 B.n431 10.6151
R1500 B.n433 B.n432 10.6151
R1501 B.n433 B.n397 10.6151
R1502 B.n439 B.n397 10.6151
R1503 B.n440 B.n439 10.6151
R1504 B.n441 B.n440 10.6151
R1505 B.n441 B.n395 10.6151
R1506 B.n447 B.n395 10.6151
R1507 B.n448 B.n447 10.6151
R1508 B.n449 B.n448 10.6151
R1509 B.n449 B.n393 10.6151
R1510 B.n455 B.n393 10.6151
R1511 B.n456 B.n455 10.6151
R1512 B.n457 B.n456 10.6151
R1513 B.n457 B.n391 10.6151
R1514 B.n464 B.n463 10.6151
R1515 B.n465 B.n464 10.6151
R1516 B.n465 B.n386 10.6151
R1517 B.n471 B.n386 10.6151
R1518 B.n472 B.n471 10.6151
R1519 B.n473 B.n472 10.6151
R1520 B.n473 B.n384 10.6151
R1521 B.n479 B.n384 10.6151
R1522 B.n482 B.n481 10.6151
R1523 B.n482 B.n380 10.6151
R1524 B.n488 B.n380 10.6151
R1525 B.n489 B.n488 10.6151
R1526 B.n490 B.n489 10.6151
R1527 B.n490 B.n378 10.6151
R1528 B.n496 B.n378 10.6151
R1529 B.n497 B.n496 10.6151
R1530 B.n498 B.n497 10.6151
R1531 B.n498 B.n376 10.6151
R1532 B.n504 B.n376 10.6151
R1533 B.n505 B.n504 10.6151
R1534 B.n506 B.n505 10.6151
R1535 B.n506 B.n374 10.6151
R1536 B.n512 B.n374 10.6151
R1537 B.n513 B.n512 10.6151
R1538 B.n514 B.n513 10.6151
R1539 B.n514 B.n372 10.6151
R1540 B.n520 B.n372 10.6151
R1541 B.n521 B.n520 10.6151
R1542 B.n522 B.n521 10.6151
R1543 B.n522 B.n370 10.6151
R1544 B.n528 B.n370 10.6151
R1545 B.n529 B.n528 10.6151
R1546 B.n530 B.n529 10.6151
R1547 B.n530 B.n368 10.6151
R1548 B.n536 B.n368 10.6151
R1549 B.n537 B.n536 10.6151
R1550 B.n543 B.n542 10.6151
R1551 B.n544 B.n543 10.6151
R1552 B.n544 B.n356 10.6151
R1553 B.n554 B.n356 10.6151
R1554 B.n555 B.n554 10.6151
R1555 B.n556 B.n555 10.6151
R1556 B.n556 B.n348 10.6151
R1557 B.n566 B.n348 10.6151
R1558 B.n567 B.n566 10.6151
R1559 B.n568 B.n567 10.6151
R1560 B.n568 B.n340 10.6151
R1561 B.n578 B.n340 10.6151
R1562 B.n579 B.n578 10.6151
R1563 B.n580 B.n579 10.6151
R1564 B.n580 B.n332 10.6151
R1565 B.n590 B.n332 10.6151
R1566 B.n591 B.n590 10.6151
R1567 B.n592 B.n591 10.6151
R1568 B.n592 B.n324 10.6151
R1569 B.n602 B.n324 10.6151
R1570 B.n603 B.n602 10.6151
R1571 B.n604 B.n603 10.6151
R1572 B.n604 B.n316 10.6151
R1573 B.n614 B.n316 10.6151
R1574 B.n615 B.n614 10.6151
R1575 B.n616 B.n615 10.6151
R1576 B.n616 B.n308 10.6151
R1577 B.n626 B.n308 10.6151
R1578 B.n627 B.n626 10.6151
R1579 B.n628 B.n627 10.6151
R1580 B.n628 B.n300 10.6151
R1581 B.n638 B.n300 10.6151
R1582 B.n639 B.n638 10.6151
R1583 B.n640 B.n639 10.6151
R1584 B.n640 B.n292 10.6151
R1585 B.n651 B.n292 10.6151
R1586 B.n652 B.n651 10.6151
R1587 B.n653 B.n652 10.6151
R1588 B.n653 B.n285 10.6151
R1589 B.n663 B.n285 10.6151
R1590 B.n664 B.n663 10.6151
R1591 B.n665 B.n664 10.6151
R1592 B.n665 B.n277 10.6151
R1593 B.n676 B.n277 10.6151
R1594 B.n677 B.n676 10.6151
R1595 B.n678 B.n677 10.6151
R1596 B.n678 B.n270 10.6151
R1597 B.n689 B.n270 10.6151
R1598 B.n690 B.n689 10.6151
R1599 B.n691 B.n690 10.6151
R1600 B.n691 B.n0 10.6151
R1601 B.n866 B.n1 10.6151
R1602 B.n866 B.n865 10.6151
R1603 B.n865 B.n864 10.6151
R1604 B.n864 B.n10 10.6151
R1605 B.n858 B.n10 10.6151
R1606 B.n858 B.n857 10.6151
R1607 B.n857 B.n856 10.6151
R1608 B.n856 B.n16 10.6151
R1609 B.n850 B.n16 10.6151
R1610 B.n850 B.n849 10.6151
R1611 B.n849 B.n848 10.6151
R1612 B.n848 B.n24 10.6151
R1613 B.n842 B.n24 10.6151
R1614 B.n842 B.n841 10.6151
R1615 B.n841 B.n840 10.6151
R1616 B.n840 B.n30 10.6151
R1617 B.n834 B.n30 10.6151
R1618 B.n834 B.n833 10.6151
R1619 B.n833 B.n832 10.6151
R1620 B.n832 B.n38 10.6151
R1621 B.n826 B.n38 10.6151
R1622 B.n826 B.n825 10.6151
R1623 B.n825 B.n824 10.6151
R1624 B.n824 B.n45 10.6151
R1625 B.n818 B.n45 10.6151
R1626 B.n818 B.n817 10.6151
R1627 B.n817 B.n816 10.6151
R1628 B.n816 B.n52 10.6151
R1629 B.n810 B.n52 10.6151
R1630 B.n810 B.n809 10.6151
R1631 B.n809 B.n808 10.6151
R1632 B.n808 B.n59 10.6151
R1633 B.n802 B.n59 10.6151
R1634 B.n802 B.n801 10.6151
R1635 B.n801 B.n800 10.6151
R1636 B.n800 B.n66 10.6151
R1637 B.n794 B.n66 10.6151
R1638 B.n794 B.n793 10.6151
R1639 B.n793 B.n792 10.6151
R1640 B.n792 B.n73 10.6151
R1641 B.n786 B.n73 10.6151
R1642 B.n786 B.n785 10.6151
R1643 B.n785 B.n784 10.6151
R1644 B.n784 B.n80 10.6151
R1645 B.n778 B.n80 10.6151
R1646 B.n778 B.n777 10.6151
R1647 B.n777 B.n776 10.6151
R1648 B.n776 B.n87 10.6151
R1649 B.n770 B.n87 10.6151
R1650 B.n770 B.n769 10.6151
R1651 B.n769 B.n768 10.6151
R1652 B.n648 B.t3 9.41318
R1653 B.n32 B.t2 9.41318
R1654 B.n193 B.n192 6.5566
R1655 B.n209 B.n133 6.5566
R1656 B.n463 B.n390 6.5566
R1657 B.n480 B.n479 6.5566
R1658 B.n192 B.n191 4.05904
R1659 B.n212 B.n133 4.05904
R1660 B.n391 B.n390 4.05904
R1661 B.n481 B.n480 4.05904
R1662 B.n872 B.n0 2.81026
R1663 B.n872 B.n1 2.81026
R1664 B.n680 B.t5 0.856198
R1665 B.n860 B.t7 0.856198
R1666 VN.n50 VN.n49 161.3
R1667 VN.n48 VN.n27 161.3
R1668 VN.n47 VN.n46 161.3
R1669 VN.n45 VN.n28 161.3
R1670 VN.n44 VN.n43 161.3
R1671 VN.n42 VN.n29 161.3
R1672 VN.n41 VN.n40 161.3
R1673 VN.n39 VN.n30 161.3
R1674 VN.n38 VN.n37 161.3
R1675 VN.n36 VN.n31 161.3
R1676 VN.n35 VN.n34 161.3
R1677 VN.n24 VN.n23 161.3
R1678 VN.n22 VN.n1 161.3
R1679 VN.n21 VN.n20 161.3
R1680 VN.n19 VN.n2 161.3
R1681 VN.n18 VN.n17 161.3
R1682 VN.n16 VN.n3 161.3
R1683 VN.n15 VN.n14 161.3
R1684 VN.n13 VN.n4 161.3
R1685 VN.n12 VN.n11 161.3
R1686 VN.n10 VN.n5 161.3
R1687 VN.n9 VN.n8 161.3
R1688 VN.n7 VN.t2 100.642
R1689 VN.n33 VN.t5 100.642
R1690 VN.n0 VN.t4 68.4192
R1691 VN.n16 VN.t1 68.4192
R1692 VN.n6 VN.t6 68.4192
R1693 VN.n26 VN.t3 68.4192
R1694 VN.n42 VN.t0 68.4192
R1695 VN.n32 VN.t7 68.4192
R1696 VN.n51 VN.n26 65.6537
R1697 VN.n25 VN.n0 65.6537
R1698 VN.n33 VN.n32 49.0351
R1699 VN.n7 VN.n6 49.0351
R1700 VN VN.n51 48.1496
R1701 VN.n11 VN.n10 40.577
R1702 VN.n11 VN.n4 40.577
R1703 VN.n21 VN.n2 40.577
R1704 VN.n22 VN.n21 40.577
R1705 VN.n37 VN.n36 40.577
R1706 VN.n37 VN.n30 40.577
R1707 VN.n47 VN.n28 40.577
R1708 VN.n48 VN.n47 40.577
R1709 VN.n9 VN.n6 24.5923
R1710 VN.n10 VN.n9 24.5923
R1711 VN.n15 VN.n4 24.5923
R1712 VN.n16 VN.n15 24.5923
R1713 VN.n17 VN.n16 24.5923
R1714 VN.n17 VN.n2 24.5923
R1715 VN.n23 VN.n22 24.5923
R1716 VN.n23 VN.n0 24.5923
R1717 VN.n36 VN.n35 24.5923
R1718 VN.n35 VN.n32 24.5923
R1719 VN.n43 VN.n28 24.5923
R1720 VN.n43 VN.n42 24.5923
R1721 VN.n42 VN.n41 24.5923
R1722 VN.n41 VN.n30 24.5923
R1723 VN.n49 VN.n26 24.5923
R1724 VN.n49 VN.n48 24.5923
R1725 VN.n34 VN.n33 5.17221
R1726 VN.n8 VN.n7 5.17221
R1727 VN.n51 VN.n50 0.354861
R1728 VN.n25 VN.n24 0.354861
R1729 VN VN.n25 0.267071
R1730 VN.n50 VN.n27 0.189894
R1731 VN.n46 VN.n27 0.189894
R1732 VN.n46 VN.n45 0.189894
R1733 VN.n45 VN.n44 0.189894
R1734 VN.n44 VN.n29 0.189894
R1735 VN.n40 VN.n29 0.189894
R1736 VN.n40 VN.n39 0.189894
R1737 VN.n39 VN.n38 0.189894
R1738 VN.n38 VN.n31 0.189894
R1739 VN.n34 VN.n31 0.189894
R1740 VN.n8 VN.n5 0.189894
R1741 VN.n12 VN.n5 0.189894
R1742 VN.n13 VN.n12 0.189894
R1743 VN.n14 VN.n13 0.189894
R1744 VN.n14 VN.n3 0.189894
R1745 VN.n18 VN.n3 0.189894
R1746 VN.n19 VN.n18 0.189894
R1747 VN.n20 VN.n19 0.189894
R1748 VN.n20 VN.n1 0.189894
R1749 VN.n24 VN.n1 0.189894
R1750 VDD2.n2 VDD2.n1 68.244
R1751 VDD2.n2 VDD2.n0 68.244
R1752 VDD2 VDD2.n5 68.2412
R1753 VDD2.n4 VDD2.n3 67.0064
R1754 VDD2.n4 VDD2.n2 41.8877
R1755 VDD2.n5 VDD2.t0 2.61264
R1756 VDD2.n5 VDD2.t2 2.61264
R1757 VDD2.n3 VDD2.t4 2.61264
R1758 VDD2.n3 VDD2.t7 2.61264
R1759 VDD2.n1 VDD2.t6 2.61264
R1760 VDD2.n1 VDD2.t3 2.61264
R1761 VDD2.n0 VDD2.t5 2.61264
R1762 VDD2.n0 VDD2.t1 2.61264
R1763 VDD2 VDD2.n4 1.35179
C0 VDD1 VN 0.151696f
C1 VDD2 VN 5.69472f
C2 VTAIL VP 6.31822f
C3 VDD2 VDD1 1.81036f
C4 VTAIL VN 6.30411f
C5 VTAIL VDD1 6.62722f
C6 VP VN 6.92807f
C7 VDD2 VTAIL 6.68211f
C8 VP VDD1 6.06856f
C9 VDD2 VP 0.526961f
C10 VDD2 B 5.056567f
C11 VDD1 B 5.503826f
C12 VTAIL B 7.889149f
C13 VN B 15.453069f
C14 VP B 14.090392f
C15 VDD2.t5 B 0.145523f
C16 VDD2.t1 B 0.145523f
C17 VDD2.n0 B 1.26403f
C18 VDD2.t6 B 0.145523f
C19 VDD2.t3 B 0.145523f
C20 VDD2.n1 B 1.26403f
C21 VDD2.n2 B 2.94351f
C22 VDD2.t4 B 0.145523f
C23 VDD2.t7 B 0.145523f
C24 VDD2.n3 B 1.25495f
C25 VDD2.n4 B 2.55144f
C26 VDD2.t0 B 0.145523f
C27 VDD2.t2 B 0.145523f
C28 VDD2.n5 B 1.264f
C29 VN.t4 B 1.25919f
C30 VN.n0 B 0.549576f
C31 VN.n1 B 0.023222f
C32 VN.n2 B 0.045911f
C33 VN.n3 B 0.023222f
C34 VN.t1 B 1.25919f
C35 VN.n4 B 0.045911f
C36 VN.n5 B 0.023222f
C37 VN.t6 B 1.25919f
C38 VN.n6 B 0.541439f
C39 VN.t2 B 1.45423f
C40 VN.n7 B 0.512245f
C41 VN.n8 B 0.240188f
C42 VN.n9 B 0.043063f
C43 VN.n10 B 0.045911f
C44 VN.n11 B 0.018756f
C45 VN.n12 B 0.023222f
C46 VN.n13 B 0.023222f
C47 VN.n14 B 0.023222f
C48 VN.n15 B 0.043063f
C49 VN.n16 B 0.4821f
C50 VN.n17 B 0.043063f
C51 VN.n18 B 0.023222f
C52 VN.n19 B 0.023222f
C53 VN.n20 B 0.023222f
C54 VN.n21 B 0.018756f
C55 VN.n22 B 0.045911f
C56 VN.n23 B 0.043063f
C57 VN.n24 B 0.037474f
C58 VN.n25 B 0.041209f
C59 VN.t3 B 1.25919f
C60 VN.n26 B 0.549576f
C61 VN.n27 B 0.023222f
C62 VN.n28 B 0.045911f
C63 VN.n29 B 0.023222f
C64 VN.t0 B 1.25919f
C65 VN.n30 B 0.045911f
C66 VN.n31 B 0.023222f
C67 VN.t7 B 1.25919f
C68 VN.n32 B 0.541439f
C69 VN.t5 B 1.45423f
C70 VN.n33 B 0.512245f
C71 VN.n34 B 0.240188f
C72 VN.n35 B 0.043063f
C73 VN.n36 B 0.045911f
C74 VN.n37 B 0.018756f
C75 VN.n38 B 0.023222f
C76 VN.n39 B 0.023222f
C77 VN.n40 B 0.023222f
C78 VN.n41 B 0.043063f
C79 VN.n42 B 0.4821f
C80 VN.n43 B 0.043063f
C81 VN.n44 B 0.023222f
C82 VN.n45 B 0.023222f
C83 VN.n46 B 0.023222f
C84 VN.n47 B 0.018756f
C85 VN.n48 B 0.045911f
C86 VN.n49 B 0.043063f
C87 VN.n50 B 0.037474f
C88 VN.n51 B 1.23738f
C89 VDD1.t0 B 0.147973f
C90 VDD1.t7 B 0.147973f
C91 VDD1.n0 B 1.28632f
C92 VDD1.t2 B 0.147973f
C93 VDD1.t6 B 0.147973f
C94 VDD1.n1 B 1.28531f
C95 VDD1.t1 B 0.147973f
C96 VDD1.t3 B 0.147973f
C97 VDD1.n2 B 1.28531f
C98 VDD1.n3 B 3.04462f
C99 VDD1.t4 B 0.147973f
C100 VDD1.t5 B 0.147973f
C101 VDD1.n4 B 1.27607f
C102 VDD1.n5 B 2.62481f
C103 VTAIL.t2 B 0.130583f
C104 VTAIL.t0 B 0.130583f
C105 VTAIL.n0 B 1.07052f
C106 VTAIL.n1 B 0.383595f
C107 VTAIL.t7 B 1.3627f
C108 VTAIL.n2 B 0.476462f
C109 VTAIL.t8 B 1.3627f
C110 VTAIL.n3 B 0.476462f
C111 VTAIL.t11 B 0.130583f
C112 VTAIL.t14 B 0.130583f
C113 VTAIL.n4 B 1.07052f
C114 VTAIL.n5 B 0.561177f
C115 VTAIL.t12 B 1.3627f
C116 VTAIL.n6 B 1.38028f
C117 VTAIL.t1 B 1.3627f
C118 VTAIL.n7 B 1.38027f
C119 VTAIL.t6 B 0.130583f
C120 VTAIL.t3 B 0.130583f
C121 VTAIL.n8 B 1.07052f
C122 VTAIL.n9 B 0.561174f
C123 VTAIL.t5 B 1.3627f
C124 VTAIL.n10 B 0.476459f
C125 VTAIL.t9 B 1.3627f
C126 VTAIL.n11 B 0.476459f
C127 VTAIL.t13 B 0.130583f
C128 VTAIL.t15 B 0.130583f
C129 VTAIL.n12 B 1.07052f
C130 VTAIL.n13 B 0.561174f
C131 VTAIL.t10 B 1.3627f
C132 VTAIL.n14 B 1.38028f
C133 VTAIL.t4 B 1.3627f
C134 VTAIL.n15 B 1.37619f
C135 VP.t4 B 1.28806f
C136 VP.n0 B 0.562179f
C137 VP.n1 B 0.023755f
C138 VP.n2 B 0.046963f
C139 VP.n3 B 0.023755f
C140 VP.t6 B 1.28806f
C141 VP.n4 B 0.046963f
C142 VP.n5 B 0.023755f
C143 VP.t1 B 1.28806f
C144 VP.n6 B 0.493155f
C145 VP.n7 B 0.023755f
C146 VP.n8 B 0.046963f
C147 VP.t2 B 1.28806f
C148 VP.n9 B 0.562179f
C149 VP.n10 B 0.023755f
C150 VP.n11 B 0.046963f
C151 VP.n12 B 0.023755f
C152 VP.t3 B 1.28806f
C153 VP.n13 B 0.046963f
C154 VP.n14 B 0.023755f
C155 VP.t0 B 1.28806f
C156 VP.n15 B 0.553854f
C157 VP.t7 B 1.48757f
C158 VP.n16 B 0.523992f
C159 VP.n17 B 0.245696f
C160 VP.n18 B 0.044051f
C161 VP.n19 B 0.046963f
C162 VP.n20 B 0.019186f
C163 VP.n21 B 0.023755f
C164 VP.n22 B 0.023755f
C165 VP.n23 B 0.023755f
C166 VP.n24 B 0.044051f
C167 VP.n25 B 0.493155f
C168 VP.n26 B 0.044051f
C169 VP.n27 B 0.023755f
C170 VP.n28 B 0.023755f
C171 VP.n29 B 0.023755f
C172 VP.n30 B 0.019186f
C173 VP.n31 B 0.046963f
C174 VP.n32 B 0.044051f
C175 VP.n33 B 0.038333f
C176 VP.n34 B 1.25588f
C177 VP.n35 B 1.27373f
C178 VP.t5 B 1.28806f
C179 VP.n36 B 0.562179f
C180 VP.n37 B 0.044051f
C181 VP.n38 B 0.038333f
C182 VP.n39 B 0.023755f
C183 VP.n40 B 0.023755f
C184 VP.n41 B 0.019186f
C185 VP.n42 B 0.046963f
C186 VP.n43 B 0.044051f
C187 VP.n44 B 0.023755f
C188 VP.n45 B 0.023755f
C189 VP.n46 B 0.023755f
C190 VP.n47 B 0.044051f
C191 VP.n48 B 0.046963f
C192 VP.n49 B 0.019186f
C193 VP.n50 B 0.023755f
C194 VP.n51 B 0.023755f
C195 VP.n52 B 0.023755f
C196 VP.n53 B 0.044051f
C197 VP.n54 B 0.493155f
C198 VP.n55 B 0.044051f
C199 VP.n56 B 0.023755f
C200 VP.n57 B 0.023755f
C201 VP.n58 B 0.023755f
C202 VP.n59 B 0.019186f
C203 VP.n60 B 0.046963f
C204 VP.n61 B 0.044051f
C205 VP.n62 B 0.038333f
C206 VP.n63 B 0.042154f
.ends

