* NGSPICE file created from diff_pair_sample_0865.ext - technology: sky130A

.subckt diff_pair_sample_0865 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=1.1517 ps=7.31 w=6.98 l=1.01
X1 B.t11 B.t9 B.t10 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=0 ps=0 w=6.98 l=1.01
X2 VDD2.t5 VN.t0 VTAIL.t1 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=1.1517 ps=7.31 w=6.98 l=1.01
X3 B.t8 B.t6 B.t7 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=0 ps=0 w=6.98 l=1.01
X4 VDD1.t4 VP.t1 VTAIL.t7 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=2.7222 ps=14.74 w=6.98 l=1.01
X5 VDD1.t3 VP.t2 VTAIL.t11 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=1.1517 ps=7.31 w=6.98 l=1.01
X6 VTAIL.t6 VP.t3 VDD1.t2 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=1.1517 ps=7.31 w=6.98 l=1.01
X7 VDD2.t4 VN.t1 VTAIL.t2 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=2.7222 ps=14.74 w=6.98 l=1.01
X8 VTAIL.t10 VP.t4 VDD1.t1 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=1.1517 ps=7.31 w=6.98 l=1.01
X9 B.t5 B.t3 B.t4 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=0 ps=0 w=6.98 l=1.01
X10 B.t2 B.t0 B.t1 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=0 ps=0 w=6.98 l=1.01
X11 VDD2.t3 VN.t2 VTAIL.t3 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=2.7222 pd=14.74 as=1.1517 ps=7.31 w=6.98 l=1.01
X12 VDD1.t0 VP.t5 VTAIL.t8 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=2.7222 ps=14.74 w=6.98 l=1.01
X13 VDD2.t2 VN.t3 VTAIL.t4 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=2.7222 ps=14.74 w=6.98 l=1.01
X14 VTAIL.t5 VN.t4 VDD2.t1 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=1.1517 ps=7.31 w=6.98 l=1.01
X15 VTAIL.t0 VN.t5 VDD2.t0 w_n2042_n2364# sky130_fd_pr__pfet_01v8 ad=1.1517 pd=7.31 as=1.1517 ps=7.31 w=6.98 l=1.01
R0 VP.n3 VP.t0 228.374
R1 VP.n8 VP.t2 205.924
R2 VP.n14 VP.t1 205.924
R3 VP.n6 VP.t5 205.924
R4 VP.n12 VP.t3 166.553
R5 VP.n4 VP.t4 166.553
R6 VP.n5 VP.n2 161.3
R7 VP.n13 VP.n0 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n10 VP.n1 161.3
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 48.4439
R14 VP.n14 VP.n13 48.4439
R15 VP.n6 VP.n5 48.4439
R16 VP.n9 VP.n7 38.7362
R17 VP.n4 VP.n3 32.0779
R18 VP.n3 VP.n2 28.4181
R19 VP.n12 VP.n1 24.3439
R20 VP.n13 VP.n12 24.3439
R21 VP.n5 VP.n4 24.3439
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n7 VTAIL.t2 72.8048
R29 VTAIL.n11 VTAIL.t4 72.8046
R30 VTAIL.n2 VTAIL.t7 72.8046
R31 VTAIL.n10 VTAIL.t8 72.8046
R32 VTAIL.n9 VTAIL.n8 68.1479
R33 VTAIL.n6 VTAIL.n5 68.1479
R34 VTAIL.n1 VTAIL.n0 68.1479
R35 VTAIL.n4 VTAIL.n3 68.1479
R36 VTAIL.n6 VTAIL.n4 20.6945
R37 VTAIL.n11 VTAIL.n10 19.5393
R38 VTAIL.n0 VTAIL.t3 4.65738
R39 VTAIL.n0 VTAIL.t5 4.65738
R40 VTAIL.n3 VTAIL.t11 4.65738
R41 VTAIL.n3 VTAIL.t6 4.65738
R42 VTAIL.n8 VTAIL.t9 4.65738
R43 VTAIL.n8 VTAIL.t10 4.65738
R44 VTAIL.n5 VTAIL.t1 4.65738
R45 VTAIL.n5 VTAIL.t0 4.65738
R46 VTAIL.n7 VTAIL.n6 1.15567
R47 VTAIL.n10 VTAIL.n9 1.15567
R48 VTAIL.n4 VTAIL.n2 1.15567
R49 VTAIL.n9 VTAIL.n7 1.04791
R50 VTAIL.n2 VTAIL.n1 1.04791
R51 VTAIL VTAIL.n11 0.80869
R52 VTAIL VTAIL.n1 0.347483
R53 VDD1 VDD1.t5 90.4082
R54 VDD1.n1 VDD1.t3 90.2944
R55 VDD1.n1 VDD1.n0 85.0601
R56 VDD1.n3 VDD1.n2 84.8266
R57 VDD1.n3 VDD1.n1 34.6474
R58 VDD1.n2 VDD1.t1 4.65738
R59 VDD1.n2 VDD1.t0 4.65738
R60 VDD1.n0 VDD1.t2 4.65738
R61 VDD1.n0 VDD1.t4 4.65738
R62 VDD1 VDD1.n3 0.231103
R63 B.n327 B.n326 585
R64 B.n328 B.n49 585
R65 B.n330 B.n329 585
R66 B.n331 B.n48 585
R67 B.n333 B.n332 585
R68 B.n334 B.n47 585
R69 B.n336 B.n335 585
R70 B.n337 B.n46 585
R71 B.n339 B.n338 585
R72 B.n340 B.n45 585
R73 B.n342 B.n341 585
R74 B.n343 B.n44 585
R75 B.n345 B.n344 585
R76 B.n346 B.n43 585
R77 B.n348 B.n347 585
R78 B.n349 B.n42 585
R79 B.n351 B.n350 585
R80 B.n352 B.n41 585
R81 B.n354 B.n353 585
R82 B.n355 B.n40 585
R83 B.n357 B.n356 585
R84 B.n358 B.n39 585
R85 B.n360 B.n359 585
R86 B.n361 B.n38 585
R87 B.n363 B.n362 585
R88 B.n364 B.n37 585
R89 B.n366 B.n365 585
R90 B.n368 B.n367 585
R91 B.n369 B.n33 585
R92 B.n371 B.n370 585
R93 B.n372 B.n32 585
R94 B.n374 B.n373 585
R95 B.n375 B.n31 585
R96 B.n377 B.n376 585
R97 B.n378 B.n30 585
R98 B.n380 B.n379 585
R99 B.n382 B.n27 585
R100 B.n384 B.n383 585
R101 B.n385 B.n26 585
R102 B.n387 B.n386 585
R103 B.n388 B.n25 585
R104 B.n390 B.n389 585
R105 B.n391 B.n24 585
R106 B.n393 B.n392 585
R107 B.n394 B.n23 585
R108 B.n396 B.n395 585
R109 B.n397 B.n22 585
R110 B.n399 B.n398 585
R111 B.n400 B.n21 585
R112 B.n402 B.n401 585
R113 B.n403 B.n20 585
R114 B.n405 B.n404 585
R115 B.n406 B.n19 585
R116 B.n408 B.n407 585
R117 B.n409 B.n18 585
R118 B.n411 B.n410 585
R119 B.n412 B.n17 585
R120 B.n414 B.n413 585
R121 B.n415 B.n16 585
R122 B.n417 B.n416 585
R123 B.n418 B.n15 585
R124 B.n420 B.n419 585
R125 B.n421 B.n14 585
R126 B.n325 B.n50 585
R127 B.n324 B.n323 585
R128 B.n322 B.n51 585
R129 B.n321 B.n320 585
R130 B.n319 B.n52 585
R131 B.n318 B.n317 585
R132 B.n316 B.n53 585
R133 B.n315 B.n314 585
R134 B.n313 B.n54 585
R135 B.n312 B.n311 585
R136 B.n310 B.n55 585
R137 B.n309 B.n308 585
R138 B.n307 B.n56 585
R139 B.n306 B.n305 585
R140 B.n304 B.n57 585
R141 B.n303 B.n302 585
R142 B.n301 B.n58 585
R143 B.n300 B.n299 585
R144 B.n298 B.n59 585
R145 B.n297 B.n296 585
R146 B.n295 B.n60 585
R147 B.n294 B.n293 585
R148 B.n292 B.n61 585
R149 B.n291 B.n290 585
R150 B.n289 B.n62 585
R151 B.n288 B.n287 585
R152 B.n286 B.n63 585
R153 B.n285 B.n284 585
R154 B.n283 B.n64 585
R155 B.n282 B.n281 585
R156 B.n280 B.n65 585
R157 B.n279 B.n278 585
R158 B.n277 B.n66 585
R159 B.n276 B.n275 585
R160 B.n274 B.n67 585
R161 B.n273 B.n272 585
R162 B.n271 B.n68 585
R163 B.n270 B.n269 585
R164 B.n268 B.n69 585
R165 B.n267 B.n266 585
R166 B.n265 B.n70 585
R167 B.n264 B.n263 585
R168 B.n262 B.n71 585
R169 B.n261 B.n260 585
R170 B.n259 B.n72 585
R171 B.n258 B.n257 585
R172 B.n256 B.n73 585
R173 B.n255 B.n254 585
R174 B.n253 B.n74 585
R175 B.n157 B.n110 585
R176 B.n159 B.n158 585
R177 B.n160 B.n109 585
R178 B.n162 B.n161 585
R179 B.n163 B.n108 585
R180 B.n165 B.n164 585
R181 B.n166 B.n107 585
R182 B.n168 B.n167 585
R183 B.n169 B.n106 585
R184 B.n171 B.n170 585
R185 B.n172 B.n105 585
R186 B.n174 B.n173 585
R187 B.n175 B.n104 585
R188 B.n177 B.n176 585
R189 B.n178 B.n103 585
R190 B.n180 B.n179 585
R191 B.n181 B.n102 585
R192 B.n183 B.n182 585
R193 B.n184 B.n101 585
R194 B.n186 B.n185 585
R195 B.n187 B.n100 585
R196 B.n189 B.n188 585
R197 B.n190 B.n99 585
R198 B.n192 B.n191 585
R199 B.n193 B.n98 585
R200 B.n195 B.n194 585
R201 B.n196 B.n95 585
R202 B.n199 B.n198 585
R203 B.n200 B.n94 585
R204 B.n202 B.n201 585
R205 B.n203 B.n93 585
R206 B.n205 B.n204 585
R207 B.n206 B.n92 585
R208 B.n208 B.n207 585
R209 B.n209 B.n91 585
R210 B.n211 B.n210 585
R211 B.n213 B.n212 585
R212 B.n214 B.n87 585
R213 B.n216 B.n215 585
R214 B.n217 B.n86 585
R215 B.n219 B.n218 585
R216 B.n220 B.n85 585
R217 B.n222 B.n221 585
R218 B.n223 B.n84 585
R219 B.n225 B.n224 585
R220 B.n226 B.n83 585
R221 B.n228 B.n227 585
R222 B.n229 B.n82 585
R223 B.n231 B.n230 585
R224 B.n232 B.n81 585
R225 B.n234 B.n233 585
R226 B.n235 B.n80 585
R227 B.n237 B.n236 585
R228 B.n238 B.n79 585
R229 B.n240 B.n239 585
R230 B.n241 B.n78 585
R231 B.n243 B.n242 585
R232 B.n244 B.n77 585
R233 B.n246 B.n245 585
R234 B.n247 B.n76 585
R235 B.n249 B.n248 585
R236 B.n250 B.n75 585
R237 B.n252 B.n251 585
R238 B.n156 B.n155 585
R239 B.n154 B.n111 585
R240 B.n153 B.n152 585
R241 B.n151 B.n112 585
R242 B.n150 B.n149 585
R243 B.n148 B.n113 585
R244 B.n147 B.n146 585
R245 B.n145 B.n114 585
R246 B.n144 B.n143 585
R247 B.n142 B.n115 585
R248 B.n141 B.n140 585
R249 B.n139 B.n116 585
R250 B.n138 B.n137 585
R251 B.n136 B.n117 585
R252 B.n135 B.n134 585
R253 B.n133 B.n118 585
R254 B.n132 B.n131 585
R255 B.n130 B.n119 585
R256 B.n129 B.n128 585
R257 B.n127 B.n120 585
R258 B.n126 B.n125 585
R259 B.n124 B.n121 585
R260 B.n123 B.n122 585
R261 B.n2 B.n0 585
R262 B.n457 B.n1 585
R263 B.n456 B.n455 585
R264 B.n454 B.n3 585
R265 B.n453 B.n452 585
R266 B.n451 B.n4 585
R267 B.n450 B.n449 585
R268 B.n448 B.n5 585
R269 B.n447 B.n446 585
R270 B.n445 B.n6 585
R271 B.n444 B.n443 585
R272 B.n442 B.n7 585
R273 B.n441 B.n440 585
R274 B.n439 B.n8 585
R275 B.n438 B.n437 585
R276 B.n436 B.n9 585
R277 B.n435 B.n434 585
R278 B.n433 B.n10 585
R279 B.n432 B.n431 585
R280 B.n430 B.n11 585
R281 B.n429 B.n428 585
R282 B.n427 B.n12 585
R283 B.n426 B.n425 585
R284 B.n424 B.n13 585
R285 B.n423 B.n422 585
R286 B.n459 B.n458 585
R287 B.n157 B.n156 502.111
R288 B.n422 B.n421 502.111
R289 B.n253 B.n252 502.111
R290 B.n326 B.n325 502.111
R291 B.n88 B.t9 369.546
R292 B.n96 B.t6 369.546
R293 B.n28 B.t0 369.546
R294 B.n34 B.t3 369.546
R295 B.n156 B.n111 163.367
R296 B.n152 B.n111 163.367
R297 B.n152 B.n151 163.367
R298 B.n151 B.n150 163.367
R299 B.n150 B.n113 163.367
R300 B.n146 B.n113 163.367
R301 B.n146 B.n145 163.367
R302 B.n145 B.n144 163.367
R303 B.n144 B.n115 163.367
R304 B.n140 B.n115 163.367
R305 B.n140 B.n139 163.367
R306 B.n139 B.n138 163.367
R307 B.n138 B.n117 163.367
R308 B.n134 B.n117 163.367
R309 B.n134 B.n133 163.367
R310 B.n133 B.n132 163.367
R311 B.n132 B.n119 163.367
R312 B.n128 B.n119 163.367
R313 B.n128 B.n127 163.367
R314 B.n127 B.n126 163.367
R315 B.n126 B.n121 163.367
R316 B.n122 B.n121 163.367
R317 B.n122 B.n2 163.367
R318 B.n458 B.n2 163.367
R319 B.n458 B.n457 163.367
R320 B.n457 B.n456 163.367
R321 B.n456 B.n3 163.367
R322 B.n452 B.n3 163.367
R323 B.n452 B.n451 163.367
R324 B.n451 B.n450 163.367
R325 B.n450 B.n5 163.367
R326 B.n446 B.n5 163.367
R327 B.n446 B.n445 163.367
R328 B.n445 B.n444 163.367
R329 B.n444 B.n7 163.367
R330 B.n440 B.n7 163.367
R331 B.n440 B.n439 163.367
R332 B.n439 B.n438 163.367
R333 B.n438 B.n9 163.367
R334 B.n434 B.n9 163.367
R335 B.n434 B.n433 163.367
R336 B.n433 B.n432 163.367
R337 B.n432 B.n11 163.367
R338 B.n428 B.n11 163.367
R339 B.n428 B.n427 163.367
R340 B.n427 B.n426 163.367
R341 B.n426 B.n13 163.367
R342 B.n422 B.n13 163.367
R343 B.n158 B.n157 163.367
R344 B.n158 B.n109 163.367
R345 B.n162 B.n109 163.367
R346 B.n163 B.n162 163.367
R347 B.n164 B.n163 163.367
R348 B.n164 B.n107 163.367
R349 B.n168 B.n107 163.367
R350 B.n169 B.n168 163.367
R351 B.n170 B.n169 163.367
R352 B.n170 B.n105 163.367
R353 B.n174 B.n105 163.367
R354 B.n175 B.n174 163.367
R355 B.n176 B.n175 163.367
R356 B.n176 B.n103 163.367
R357 B.n180 B.n103 163.367
R358 B.n181 B.n180 163.367
R359 B.n182 B.n181 163.367
R360 B.n182 B.n101 163.367
R361 B.n186 B.n101 163.367
R362 B.n187 B.n186 163.367
R363 B.n188 B.n187 163.367
R364 B.n188 B.n99 163.367
R365 B.n192 B.n99 163.367
R366 B.n193 B.n192 163.367
R367 B.n194 B.n193 163.367
R368 B.n194 B.n95 163.367
R369 B.n199 B.n95 163.367
R370 B.n200 B.n199 163.367
R371 B.n201 B.n200 163.367
R372 B.n201 B.n93 163.367
R373 B.n205 B.n93 163.367
R374 B.n206 B.n205 163.367
R375 B.n207 B.n206 163.367
R376 B.n207 B.n91 163.367
R377 B.n211 B.n91 163.367
R378 B.n212 B.n211 163.367
R379 B.n212 B.n87 163.367
R380 B.n216 B.n87 163.367
R381 B.n217 B.n216 163.367
R382 B.n218 B.n217 163.367
R383 B.n218 B.n85 163.367
R384 B.n222 B.n85 163.367
R385 B.n223 B.n222 163.367
R386 B.n224 B.n223 163.367
R387 B.n224 B.n83 163.367
R388 B.n228 B.n83 163.367
R389 B.n229 B.n228 163.367
R390 B.n230 B.n229 163.367
R391 B.n230 B.n81 163.367
R392 B.n234 B.n81 163.367
R393 B.n235 B.n234 163.367
R394 B.n236 B.n235 163.367
R395 B.n236 B.n79 163.367
R396 B.n240 B.n79 163.367
R397 B.n241 B.n240 163.367
R398 B.n242 B.n241 163.367
R399 B.n242 B.n77 163.367
R400 B.n246 B.n77 163.367
R401 B.n247 B.n246 163.367
R402 B.n248 B.n247 163.367
R403 B.n248 B.n75 163.367
R404 B.n252 B.n75 163.367
R405 B.n254 B.n253 163.367
R406 B.n254 B.n73 163.367
R407 B.n258 B.n73 163.367
R408 B.n259 B.n258 163.367
R409 B.n260 B.n259 163.367
R410 B.n260 B.n71 163.367
R411 B.n264 B.n71 163.367
R412 B.n265 B.n264 163.367
R413 B.n266 B.n265 163.367
R414 B.n266 B.n69 163.367
R415 B.n270 B.n69 163.367
R416 B.n271 B.n270 163.367
R417 B.n272 B.n271 163.367
R418 B.n272 B.n67 163.367
R419 B.n276 B.n67 163.367
R420 B.n277 B.n276 163.367
R421 B.n278 B.n277 163.367
R422 B.n278 B.n65 163.367
R423 B.n282 B.n65 163.367
R424 B.n283 B.n282 163.367
R425 B.n284 B.n283 163.367
R426 B.n284 B.n63 163.367
R427 B.n288 B.n63 163.367
R428 B.n289 B.n288 163.367
R429 B.n290 B.n289 163.367
R430 B.n290 B.n61 163.367
R431 B.n294 B.n61 163.367
R432 B.n295 B.n294 163.367
R433 B.n296 B.n295 163.367
R434 B.n296 B.n59 163.367
R435 B.n300 B.n59 163.367
R436 B.n301 B.n300 163.367
R437 B.n302 B.n301 163.367
R438 B.n302 B.n57 163.367
R439 B.n306 B.n57 163.367
R440 B.n307 B.n306 163.367
R441 B.n308 B.n307 163.367
R442 B.n308 B.n55 163.367
R443 B.n312 B.n55 163.367
R444 B.n313 B.n312 163.367
R445 B.n314 B.n313 163.367
R446 B.n314 B.n53 163.367
R447 B.n318 B.n53 163.367
R448 B.n319 B.n318 163.367
R449 B.n320 B.n319 163.367
R450 B.n320 B.n51 163.367
R451 B.n324 B.n51 163.367
R452 B.n325 B.n324 163.367
R453 B.n421 B.n420 163.367
R454 B.n420 B.n15 163.367
R455 B.n416 B.n15 163.367
R456 B.n416 B.n415 163.367
R457 B.n415 B.n414 163.367
R458 B.n414 B.n17 163.367
R459 B.n410 B.n17 163.367
R460 B.n410 B.n409 163.367
R461 B.n409 B.n408 163.367
R462 B.n408 B.n19 163.367
R463 B.n404 B.n19 163.367
R464 B.n404 B.n403 163.367
R465 B.n403 B.n402 163.367
R466 B.n402 B.n21 163.367
R467 B.n398 B.n21 163.367
R468 B.n398 B.n397 163.367
R469 B.n397 B.n396 163.367
R470 B.n396 B.n23 163.367
R471 B.n392 B.n23 163.367
R472 B.n392 B.n391 163.367
R473 B.n391 B.n390 163.367
R474 B.n390 B.n25 163.367
R475 B.n386 B.n25 163.367
R476 B.n386 B.n385 163.367
R477 B.n385 B.n384 163.367
R478 B.n384 B.n27 163.367
R479 B.n379 B.n27 163.367
R480 B.n379 B.n378 163.367
R481 B.n378 B.n377 163.367
R482 B.n377 B.n31 163.367
R483 B.n373 B.n31 163.367
R484 B.n373 B.n372 163.367
R485 B.n372 B.n371 163.367
R486 B.n371 B.n33 163.367
R487 B.n367 B.n33 163.367
R488 B.n367 B.n366 163.367
R489 B.n366 B.n37 163.367
R490 B.n362 B.n37 163.367
R491 B.n362 B.n361 163.367
R492 B.n361 B.n360 163.367
R493 B.n360 B.n39 163.367
R494 B.n356 B.n39 163.367
R495 B.n356 B.n355 163.367
R496 B.n355 B.n354 163.367
R497 B.n354 B.n41 163.367
R498 B.n350 B.n41 163.367
R499 B.n350 B.n349 163.367
R500 B.n349 B.n348 163.367
R501 B.n348 B.n43 163.367
R502 B.n344 B.n43 163.367
R503 B.n344 B.n343 163.367
R504 B.n343 B.n342 163.367
R505 B.n342 B.n45 163.367
R506 B.n338 B.n45 163.367
R507 B.n338 B.n337 163.367
R508 B.n337 B.n336 163.367
R509 B.n336 B.n47 163.367
R510 B.n332 B.n47 163.367
R511 B.n332 B.n331 163.367
R512 B.n331 B.n330 163.367
R513 B.n330 B.n49 163.367
R514 B.n326 B.n49 163.367
R515 B.n88 B.t11 139.109
R516 B.n34 B.t4 139.109
R517 B.n96 B.t8 139.101
R518 B.n28 B.t1 139.101
R519 B.n89 B.t10 113.121
R520 B.n35 B.t5 113.121
R521 B.n97 B.t7 113.115
R522 B.n29 B.t2 113.115
R523 B.n90 B.n89 59.5399
R524 B.n197 B.n97 59.5399
R525 B.n381 B.n29 59.5399
R526 B.n36 B.n35 59.5399
R527 B.n423 B.n14 32.6249
R528 B.n327 B.n50 32.6249
R529 B.n251 B.n74 32.6249
R530 B.n155 B.n110 32.6249
R531 B.n89 B.n88 25.9884
R532 B.n97 B.n96 25.9884
R533 B.n29 B.n28 25.9884
R534 B.n35 B.n34 25.9884
R535 B B.n459 18.0485
R536 B.n419 B.n14 10.6151
R537 B.n419 B.n418 10.6151
R538 B.n418 B.n417 10.6151
R539 B.n417 B.n16 10.6151
R540 B.n413 B.n16 10.6151
R541 B.n413 B.n412 10.6151
R542 B.n412 B.n411 10.6151
R543 B.n411 B.n18 10.6151
R544 B.n407 B.n18 10.6151
R545 B.n407 B.n406 10.6151
R546 B.n406 B.n405 10.6151
R547 B.n405 B.n20 10.6151
R548 B.n401 B.n20 10.6151
R549 B.n401 B.n400 10.6151
R550 B.n400 B.n399 10.6151
R551 B.n399 B.n22 10.6151
R552 B.n395 B.n22 10.6151
R553 B.n395 B.n394 10.6151
R554 B.n394 B.n393 10.6151
R555 B.n393 B.n24 10.6151
R556 B.n389 B.n24 10.6151
R557 B.n389 B.n388 10.6151
R558 B.n388 B.n387 10.6151
R559 B.n387 B.n26 10.6151
R560 B.n383 B.n26 10.6151
R561 B.n383 B.n382 10.6151
R562 B.n380 B.n30 10.6151
R563 B.n376 B.n30 10.6151
R564 B.n376 B.n375 10.6151
R565 B.n375 B.n374 10.6151
R566 B.n374 B.n32 10.6151
R567 B.n370 B.n32 10.6151
R568 B.n370 B.n369 10.6151
R569 B.n369 B.n368 10.6151
R570 B.n365 B.n364 10.6151
R571 B.n364 B.n363 10.6151
R572 B.n363 B.n38 10.6151
R573 B.n359 B.n38 10.6151
R574 B.n359 B.n358 10.6151
R575 B.n358 B.n357 10.6151
R576 B.n357 B.n40 10.6151
R577 B.n353 B.n40 10.6151
R578 B.n353 B.n352 10.6151
R579 B.n352 B.n351 10.6151
R580 B.n351 B.n42 10.6151
R581 B.n347 B.n42 10.6151
R582 B.n347 B.n346 10.6151
R583 B.n346 B.n345 10.6151
R584 B.n345 B.n44 10.6151
R585 B.n341 B.n44 10.6151
R586 B.n341 B.n340 10.6151
R587 B.n340 B.n339 10.6151
R588 B.n339 B.n46 10.6151
R589 B.n335 B.n46 10.6151
R590 B.n335 B.n334 10.6151
R591 B.n334 B.n333 10.6151
R592 B.n333 B.n48 10.6151
R593 B.n329 B.n48 10.6151
R594 B.n329 B.n328 10.6151
R595 B.n328 B.n327 10.6151
R596 B.n255 B.n74 10.6151
R597 B.n256 B.n255 10.6151
R598 B.n257 B.n256 10.6151
R599 B.n257 B.n72 10.6151
R600 B.n261 B.n72 10.6151
R601 B.n262 B.n261 10.6151
R602 B.n263 B.n262 10.6151
R603 B.n263 B.n70 10.6151
R604 B.n267 B.n70 10.6151
R605 B.n268 B.n267 10.6151
R606 B.n269 B.n268 10.6151
R607 B.n269 B.n68 10.6151
R608 B.n273 B.n68 10.6151
R609 B.n274 B.n273 10.6151
R610 B.n275 B.n274 10.6151
R611 B.n275 B.n66 10.6151
R612 B.n279 B.n66 10.6151
R613 B.n280 B.n279 10.6151
R614 B.n281 B.n280 10.6151
R615 B.n281 B.n64 10.6151
R616 B.n285 B.n64 10.6151
R617 B.n286 B.n285 10.6151
R618 B.n287 B.n286 10.6151
R619 B.n287 B.n62 10.6151
R620 B.n291 B.n62 10.6151
R621 B.n292 B.n291 10.6151
R622 B.n293 B.n292 10.6151
R623 B.n293 B.n60 10.6151
R624 B.n297 B.n60 10.6151
R625 B.n298 B.n297 10.6151
R626 B.n299 B.n298 10.6151
R627 B.n299 B.n58 10.6151
R628 B.n303 B.n58 10.6151
R629 B.n304 B.n303 10.6151
R630 B.n305 B.n304 10.6151
R631 B.n305 B.n56 10.6151
R632 B.n309 B.n56 10.6151
R633 B.n310 B.n309 10.6151
R634 B.n311 B.n310 10.6151
R635 B.n311 B.n54 10.6151
R636 B.n315 B.n54 10.6151
R637 B.n316 B.n315 10.6151
R638 B.n317 B.n316 10.6151
R639 B.n317 B.n52 10.6151
R640 B.n321 B.n52 10.6151
R641 B.n322 B.n321 10.6151
R642 B.n323 B.n322 10.6151
R643 B.n323 B.n50 10.6151
R644 B.n159 B.n110 10.6151
R645 B.n160 B.n159 10.6151
R646 B.n161 B.n160 10.6151
R647 B.n161 B.n108 10.6151
R648 B.n165 B.n108 10.6151
R649 B.n166 B.n165 10.6151
R650 B.n167 B.n166 10.6151
R651 B.n167 B.n106 10.6151
R652 B.n171 B.n106 10.6151
R653 B.n172 B.n171 10.6151
R654 B.n173 B.n172 10.6151
R655 B.n173 B.n104 10.6151
R656 B.n177 B.n104 10.6151
R657 B.n178 B.n177 10.6151
R658 B.n179 B.n178 10.6151
R659 B.n179 B.n102 10.6151
R660 B.n183 B.n102 10.6151
R661 B.n184 B.n183 10.6151
R662 B.n185 B.n184 10.6151
R663 B.n185 B.n100 10.6151
R664 B.n189 B.n100 10.6151
R665 B.n190 B.n189 10.6151
R666 B.n191 B.n190 10.6151
R667 B.n191 B.n98 10.6151
R668 B.n195 B.n98 10.6151
R669 B.n196 B.n195 10.6151
R670 B.n198 B.n94 10.6151
R671 B.n202 B.n94 10.6151
R672 B.n203 B.n202 10.6151
R673 B.n204 B.n203 10.6151
R674 B.n204 B.n92 10.6151
R675 B.n208 B.n92 10.6151
R676 B.n209 B.n208 10.6151
R677 B.n210 B.n209 10.6151
R678 B.n214 B.n213 10.6151
R679 B.n215 B.n214 10.6151
R680 B.n215 B.n86 10.6151
R681 B.n219 B.n86 10.6151
R682 B.n220 B.n219 10.6151
R683 B.n221 B.n220 10.6151
R684 B.n221 B.n84 10.6151
R685 B.n225 B.n84 10.6151
R686 B.n226 B.n225 10.6151
R687 B.n227 B.n226 10.6151
R688 B.n227 B.n82 10.6151
R689 B.n231 B.n82 10.6151
R690 B.n232 B.n231 10.6151
R691 B.n233 B.n232 10.6151
R692 B.n233 B.n80 10.6151
R693 B.n237 B.n80 10.6151
R694 B.n238 B.n237 10.6151
R695 B.n239 B.n238 10.6151
R696 B.n239 B.n78 10.6151
R697 B.n243 B.n78 10.6151
R698 B.n244 B.n243 10.6151
R699 B.n245 B.n244 10.6151
R700 B.n245 B.n76 10.6151
R701 B.n249 B.n76 10.6151
R702 B.n250 B.n249 10.6151
R703 B.n251 B.n250 10.6151
R704 B.n155 B.n154 10.6151
R705 B.n154 B.n153 10.6151
R706 B.n153 B.n112 10.6151
R707 B.n149 B.n112 10.6151
R708 B.n149 B.n148 10.6151
R709 B.n148 B.n147 10.6151
R710 B.n147 B.n114 10.6151
R711 B.n143 B.n114 10.6151
R712 B.n143 B.n142 10.6151
R713 B.n142 B.n141 10.6151
R714 B.n141 B.n116 10.6151
R715 B.n137 B.n116 10.6151
R716 B.n137 B.n136 10.6151
R717 B.n136 B.n135 10.6151
R718 B.n135 B.n118 10.6151
R719 B.n131 B.n118 10.6151
R720 B.n131 B.n130 10.6151
R721 B.n130 B.n129 10.6151
R722 B.n129 B.n120 10.6151
R723 B.n125 B.n120 10.6151
R724 B.n125 B.n124 10.6151
R725 B.n124 B.n123 10.6151
R726 B.n123 B.n0 10.6151
R727 B.n455 B.n1 10.6151
R728 B.n455 B.n454 10.6151
R729 B.n454 B.n453 10.6151
R730 B.n453 B.n4 10.6151
R731 B.n449 B.n4 10.6151
R732 B.n449 B.n448 10.6151
R733 B.n448 B.n447 10.6151
R734 B.n447 B.n6 10.6151
R735 B.n443 B.n6 10.6151
R736 B.n443 B.n442 10.6151
R737 B.n442 B.n441 10.6151
R738 B.n441 B.n8 10.6151
R739 B.n437 B.n8 10.6151
R740 B.n437 B.n436 10.6151
R741 B.n436 B.n435 10.6151
R742 B.n435 B.n10 10.6151
R743 B.n431 B.n10 10.6151
R744 B.n431 B.n430 10.6151
R745 B.n430 B.n429 10.6151
R746 B.n429 B.n12 10.6151
R747 B.n425 B.n12 10.6151
R748 B.n425 B.n424 10.6151
R749 B.n424 B.n423 10.6151
R750 B.n381 B.n380 6.5566
R751 B.n368 B.n36 6.5566
R752 B.n198 B.n197 6.5566
R753 B.n210 B.n90 6.5566
R754 B.n382 B.n381 4.05904
R755 B.n365 B.n36 4.05904
R756 B.n197 B.n196 4.05904
R757 B.n213 B.n90 4.05904
R758 B.n459 B.n0 2.81026
R759 B.n459 B.n1 2.81026
R760 VN.n1 VN.t2 228.374
R761 VN.n7 VN.t1 228.374
R762 VN.n4 VN.t3 205.924
R763 VN.n10 VN.t0 205.924
R764 VN.n2 VN.t4 166.553
R765 VN.n8 VN.t5 166.553
R766 VN.n9 VN.n6 161.3
R767 VN.n3 VN.n0 161.3
R768 VN.n11 VN.n10 80.6037
R769 VN.n5 VN.n4 80.6037
R770 VN.n4 VN.n3 48.4439
R771 VN.n10 VN.n9 48.4439
R772 VN VN.n11 39.0218
R773 VN.n2 VN.n1 32.0779
R774 VN.n8 VN.n7 32.0779
R775 VN.n7 VN.n6 28.4181
R776 VN.n1 VN.n0 28.4181
R777 VN.n3 VN.n2 24.3439
R778 VN.n9 VN.n8 24.3439
R779 VN.n11 VN.n6 0.285035
R780 VN.n5 VN.n0 0.285035
R781 VN VN.n5 0.146778
R782 VDD2.n1 VDD2.t3 90.2944
R783 VDD2.n2 VDD2.t5 89.4836
R784 VDD2.n1 VDD2.n0 85.0601
R785 VDD2 VDD2.n3 85.0572
R786 VDD2.n2 VDD2.n1 33.4868
R787 VDD2.n3 VDD2.t0 4.65738
R788 VDD2.n3 VDD2.t4 4.65738
R789 VDD2.n0 VDD2.t1 4.65738
R790 VDD2.n0 VDD2.t2 4.65738
R791 VDD2 VDD2.n2 0.925069
C0 VDD1 VN 0.148293f
C1 VDD1 B 1.28033f
C2 VP VTAIL 3.17013f
C3 VDD1 VDD2 0.82338f
C4 w_n2042_n2364# VTAIL 2.15869f
C5 VP w_n2042_n2364# 3.6584f
C6 VN B 0.768655f
C7 VDD2 VN 3.11318f
C8 VDD1 VTAIL 5.99067f
C9 VDD2 B 1.31659f
C10 VDD1 VP 3.2851f
C11 VDD1 w_n2042_n2364# 1.53023f
C12 VN VTAIL 3.15578f
C13 VP VN 4.45815f
C14 B VTAIL 1.95892f
C15 VDD2 VTAIL 6.03026f
C16 VP B 1.19403f
C17 w_n2042_n2364# VN 3.39883f
C18 VP VDD2 0.322831f
C19 w_n2042_n2364# B 6.07469f
C20 w_n2042_n2364# VDD2 1.56421f
C21 VDD2 VSUBS 1.154827f
C22 VDD1 VSUBS 1.474398f
C23 VTAIL VSUBS 0.52255f
C24 VN VSUBS 4.22588f
C25 VP VSUBS 1.463641f
C26 B VSUBS 2.640964f
C27 w_n2042_n2364# VSUBS 60.0593f
C28 VDD2.t3 VSUBS 1.13448f
C29 VDD2.t1 VSUBS 0.123494f
C30 VDD2.t2 VSUBS 0.123494f
C31 VDD2.n0 VSUBS 0.849732f
C32 VDD2.n1 VSUBS 2.11221f
C33 VDD2.t5 VSUBS 1.12993f
C34 VDD2.n2 VSUBS 1.95532f
C35 VDD2.t0 VSUBS 0.123494f
C36 VDD2.t4 VSUBS 0.123494f
C37 VDD2.n3 VSUBS 0.849707f
C38 VN.n0 VSUBS 0.292296f
C39 VN.t4 VSUBS 1.01743f
C40 VN.t2 VSUBS 1.15079f
C41 VN.n1 VSUBS 0.471011f
C42 VN.n2 VSUBS 0.490632f
C43 VN.n3 VSUBS 0.063229f
C44 VN.t3 VSUBS 1.10162f
C45 VN.n4 VSUBS 0.487617f
C46 VN.n5 VSUBS 0.050648f
C47 VN.n6 VSUBS 0.292296f
C48 VN.t5 VSUBS 1.01743f
C49 VN.t1 VSUBS 1.15079f
C50 VN.n7 VSUBS 0.471011f
C51 VN.n8 VSUBS 0.490632f
C52 VN.n9 VSUBS 0.063229f
C53 VN.t0 VSUBS 1.10162f
C54 VN.n10 VSUBS 0.487617f
C55 VN.n11 VSUBS 1.99313f
C56 B.n0 VSUBS 0.003863f
C57 B.n1 VSUBS 0.003863f
C58 B.n2 VSUBS 0.006109f
C59 B.n3 VSUBS 0.006109f
C60 B.n4 VSUBS 0.006109f
C61 B.n5 VSUBS 0.006109f
C62 B.n6 VSUBS 0.006109f
C63 B.n7 VSUBS 0.006109f
C64 B.n8 VSUBS 0.006109f
C65 B.n9 VSUBS 0.006109f
C66 B.n10 VSUBS 0.006109f
C67 B.n11 VSUBS 0.006109f
C68 B.n12 VSUBS 0.006109f
C69 B.n13 VSUBS 0.006109f
C70 B.n14 VSUBS 0.014469f
C71 B.n15 VSUBS 0.006109f
C72 B.n16 VSUBS 0.006109f
C73 B.n17 VSUBS 0.006109f
C74 B.n18 VSUBS 0.006109f
C75 B.n19 VSUBS 0.006109f
C76 B.n20 VSUBS 0.006109f
C77 B.n21 VSUBS 0.006109f
C78 B.n22 VSUBS 0.006109f
C79 B.n23 VSUBS 0.006109f
C80 B.n24 VSUBS 0.006109f
C81 B.n25 VSUBS 0.006109f
C82 B.n26 VSUBS 0.006109f
C83 B.n27 VSUBS 0.006109f
C84 B.t2 VSUBS 0.183405f
C85 B.t1 VSUBS 0.192312f
C86 B.t0 VSUBS 0.271032f
C87 B.n28 VSUBS 0.091137f
C88 B.n29 VSUBS 0.056388f
C89 B.n30 VSUBS 0.006109f
C90 B.n31 VSUBS 0.006109f
C91 B.n32 VSUBS 0.006109f
C92 B.n33 VSUBS 0.006109f
C93 B.t5 VSUBS 0.183404f
C94 B.t4 VSUBS 0.19231f
C95 B.t3 VSUBS 0.271032f
C96 B.n34 VSUBS 0.091138f
C97 B.n35 VSUBS 0.056389f
C98 B.n36 VSUBS 0.014154f
C99 B.n37 VSUBS 0.006109f
C100 B.n38 VSUBS 0.006109f
C101 B.n39 VSUBS 0.006109f
C102 B.n40 VSUBS 0.006109f
C103 B.n41 VSUBS 0.006109f
C104 B.n42 VSUBS 0.006109f
C105 B.n43 VSUBS 0.006109f
C106 B.n44 VSUBS 0.006109f
C107 B.n45 VSUBS 0.006109f
C108 B.n46 VSUBS 0.006109f
C109 B.n47 VSUBS 0.006109f
C110 B.n48 VSUBS 0.006109f
C111 B.n49 VSUBS 0.006109f
C112 B.n50 VSUBS 0.014821f
C113 B.n51 VSUBS 0.006109f
C114 B.n52 VSUBS 0.006109f
C115 B.n53 VSUBS 0.006109f
C116 B.n54 VSUBS 0.006109f
C117 B.n55 VSUBS 0.006109f
C118 B.n56 VSUBS 0.006109f
C119 B.n57 VSUBS 0.006109f
C120 B.n58 VSUBS 0.006109f
C121 B.n59 VSUBS 0.006109f
C122 B.n60 VSUBS 0.006109f
C123 B.n61 VSUBS 0.006109f
C124 B.n62 VSUBS 0.006109f
C125 B.n63 VSUBS 0.006109f
C126 B.n64 VSUBS 0.006109f
C127 B.n65 VSUBS 0.006109f
C128 B.n66 VSUBS 0.006109f
C129 B.n67 VSUBS 0.006109f
C130 B.n68 VSUBS 0.006109f
C131 B.n69 VSUBS 0.006109f
C132 B.n70 VSUBS 0.006109f
C133 B.n71 VSUBS 0.006109f
C134 B.n72 VSUBS 0.006109f
C135 B.n73 VSUBS 0.006109f
C136 B.n74 VSUBS 0.014099f
C137 B.n75 VSUBS 0.006109f
C138 B.n76 VSUBS 0.006109f
C139 B.n77 VSUBS 0.006109f
C140 B.n78 VSUBS 0.006109f
C141 B.n79 VSUBS 0.006109f
C142 B.n80 VSUBS 0.006109f
C143 B.n81 VSUBS 0.006109f
C144 B.n82 VSUBS 0.006109f
C145 B.n83 VSUBS 0.006109f
C146 B.n84 VSUBS 0.006109f
C147 B.n85 VSUBS 0.006109f
C148 B.n86 VSUBS 0.006109f
C149 B.n87 VSUBS 0.006109f
C150 B.t10 VSUBS 0.183404f
C151 B.t11 VSUBS 0.19231f
C152 B.t9 VSUBS 0.271032f
C153 B.n88 VSUBS 0.091138f
C154 B.n89 VSUBS 0.056389f
C155 B.n90 VSUBS 0.014154f
C156 B.n91 VSUBS 0.006109f
C157 B.n92 VSUBS 0.006109f
C158 B.n93 VSUBS 0.006109f
C159 B.n94 VSUBS 0.006109f
C160 B.n95 VSUBS 0.006109f
C161 B.t7 VSUBS 0.183405f
C162 B.t8 VSUBS 0.192312f
C163 B.t6 VSUBS 0.271032f
C164 B.n96 VSUBS 0.091137f
C165 B.n97 VSUBS 0.056388f
C166 B.n98 VSUBS 0.006109f
C167 B.n99 VSUBS 0.006109f
C168 B.n100 VSUBS 0.006109f
C169 B.n101 VSUBS 0.006109f
C170 B.n102 VSUBS 0.006109f
C171 B.n103 VSUBS 0.006109f
C172 B.n104 VSUBS 0.006109f
C173 B.n105 VSUBS 0.006109f
C174 B.n106 VSUBS 0.006109f
C175 B.n107 VSUBS 0.006109f
C176 B.n108 VSUBS 0.006109f
C177 B.n109 VSUBS 0.006109f
C178 B.n110 VSUBS 0.014469f
C179 B.n111 VSUBS 0.006109f
C180 B.n112 VSUBS 0.006109f
C181 B.n113 VSUBS 0.006109f
C182 B.n114 VSUBS 0.006109f
C183 B.n115 VSUBS 0.006109f
C184 B.n116 VSUBS 0.006109f
C185 B.n117 VSUBS 0.006109f
C186 B.n118 VSUBS 0.006109f
C187 B.n119 VSUBS 0.006109f
C188 B.n120 VSUBS 0.006109f
C189 B.n121 VSUBS 0.006109f
C190 B.n122 VSUBS 0.006109f
C191 B.n123 VSUBS 0.006109f
C192 B.n124 VSUBS 0.006109f
C193 B.n125 VSUBS 0.006109f
C194 B.n126 VSUBS 0.006109f
C195 B.n127 VSUBS 0.006109f
C196 B.n128 VSUBS 0.006109f
C197 B.n129 VSUBS 0.006109f
C198 B.n130 VSUBS 0.006109f
C199 B.n131 VSUBS 0.006109f
C200 B.n132 VSUBS 0.006109f
C201 B.n133 VSUBS 0.006109f
C202 B.n134 VSUBS 0.006109f
C203 B.n135 VSUBS 0.006109f
C204 B.n136 VSUBS 0.006109f
C205 B.n137 VSUBS 0.006109f
C206 B.n138 VSUBS 0.006109f
C207 B.n139 VSUBS 0.006109f
C208 B.n140 VSUBS 0.006109f
C209 B.n141 VSUBS 0.006109f
C210 B.n142 VSUBS 0.006109f
C211 B.n143 VSUBS 0.006109f
C212 B.n144 VSUBS 0.006109f
C213 B.n145 VSUBS 0.006109f
C214 B.n146 VSUBS 0.006109f
C215 B.n147 VSUBS 0.006109f
C216 B.n148 VSUBS 0.006109f
C217 B.n149 VSUBS 0.006109f
C218 B.n150 VSUBS 0.006109f
C219 B.n151 VSUBS 0.006109f
C220 B.n152 VSUBS 0.006109f
C221 B.n153 VSUBS 0.006109f
C222 B.n154 VSUBS 0.006109f
C223 B.n155 VSUBS 0.014099f
C224 B.n156 VSUBS 0.014099f
C225 B.n157 VSUBS 0.014469f
C226 B.n158 VSUBS 0.006109f
C227 B.n159 VSUBS 0.006109f
C228 B.n160 VSUBS 0.006109f
C229 B.n161 VSUBS 0.006109f
C230 B.n162 VSUBS 0.006109f
C231 B.n163 VSUBS 0.006109f
C232 B.n164 VSUBS 0.006109f
C233 B.n165 VSUBS 0.006109f
C234 B.n166 VSUBS 0.006109f
C235 B.n167 VSUBS 0.006109f
C236 B.n168 VSUBS 0.006109f
C237 B.n169 VSUBS 0.006109f
C238 B.n170 VSUBS 0.006109f
C239 B.n171 VSUBS 0.006109f
C240 B.n172 VSUBS 0.006109f
C241 B.n173 VSUBS 0.006109f
C242 B.n174 VSUBS 0.006109f
C243 B.n175 VSUBS 0.006109f
C244 B.n176 VSUBS 0.006109f
C245 B.n177 VSUBS 0.006109f
C246 B.n178 VSUBS 0.006109f
C247 B.n179 VSUBS 0.006109f
C248 B.n180 VSUBS 0.006109f
C249 B.n181 VSUBS 0.006109f
C250 B.n182 VSUBS 0.006109f
C251 B.n183 VSUBS 0.006109f
C252 B.n184 VSUBS 0.006109f
C253 B.n185 VSUBS 0.006109f
C254 B.n186 VSUBS 0.006109f
C255 B.n187 VSUBS 0.006109f
C256 B.n188 VSUBS 0.006109f
C257 B.n189 VSUBS 0.006109f
C258 B.n190 VSUBS 0.006109f
C259 B.n191 VSUBS 0.006109f
C260 B.n192 VSUBS 0.006109f
C261 B.n193 VSUBS 0.006109f
C262 B.n194 VSUBS 0.006109f
C263 B.n195 VSUBS 0.006109f
C264 B.n196 VSUBS 0.004222f
C265 B.n197 VSUBS 0.014154f
C266 B.n198 VSUBS 0.004941f
C267 B.n199 VSUBS 0.006109f
C268 B.n200 VSUBS 0.006109f
C269 B.n201 VSUBS 0.006109f
C270 B.n202 VSUBS 0.006109f
C271 B.n203 VSUBS 0.006109f
C272 B.n204 VSUBS 0.006109f
C273 B.n205 VSUBS 0.006109f
C274 B.n206 VSUBS 0.006109f
C275 B.n207 VSUBS 0.006109f
C276 B.n208 VSUBS 0.006109f
C277 B.n209 VSUBS 0.006109f
C278 B.n210 VSUBS 0.004941f
C279 B.n211 VSUBS 0.006109f
C280 B.n212 VSUBS 0.006109f
C281 B.n213 VSUBS 0.004222f
C282 B.n214 VSUBS 0.006109f
C283 B.n215 VSUBS 0.006109f
C284 B.n216 VSUBS 0.006109f
C285 B.n217 VSUBS 0.006109f
C286 B.n218 VSUBS 0.006109f
C287 B.n219 VSUBS 0.006109f
C288 B.n220 VSUBS 0.006109f
C289 B.n221 VSUBS 0.006109f
C290 B.n222 VSUBS 0.006109f
C291 B.n223 VSUBS 0.006109f
C292 B.n224 VSUBS 0.006109f
C293 B.n225 VSUBS 0.006109f
C294 B.n226 VSUBS 0.006109f
C295 B.n227 VSUBS 0.006109f
C296 B.n228 VSUBS 0.006109f
C297 B.n229 VSUBS 0.006109f
C298 B.n230 VSUBS 0.006109f
C299 B.n231 VSUBS 0.006109f
C300 B.n232 VSUBS 0.006109f
C301 B.n233 VSUBS 0.006109f
C302 B.n234 VSUBS 0.006109f
C303 B.n235 VSUBS 0.006109f
C304 B.n236 VSUBS 0.006109f
C305 B.n237 VSUBS 0.006109f
C306 B.n238 VSUBS 0.006109f
C307 B.n239 VSUBS 0.006109f
C308 B.n240 VSUBS 0.006109f
C309 B.n241 VSUBS 0.006109f
C310 B.n242 VSUBS 0.006109f
C311 B.n243 VSUBS 0.006109f
C312 B.n244 VSUBS 0.006109f
C313 B.n245 VSUBS 0.006109f
C314 B.n246 VSUBS 0.006109f
C315 B.n247 VSUBS 0.006109f
C316 B.n248 VSUBS 0.006109f
C317 B.n249 VSUBS 0.006109f
C318 B.n250 VSUBS 0.006109f
C319 B.n251 VSUBS 0.014469f
C320 B.n252 VSUBS 0.014469f
C321 B.n253 VSUBS 0.014099f
C322 B.n254 VSUBS 0.006109f
C323 B.n255 VSUBS 0.006109f
C324 B.n256 VSUBS 0.006109f
C325 B.n257 VSUBS 0.006109f
C326 B.n258 VSUBS 0.006109f
C327 B.n259 VSUBS 0.006109f
C328 B.n260 VSUBS 0.006109f
C329 B.n261 VSUBS 0.006109f
C330 B.n262 VSUBS 0.006109f
C331 B.n263 VSUBS 0.006109f
C332 B.n264 VSUBS 0.006109f
C333 B.n265 VSUBS 0.006109f
C334 B.n266 VSUBS 0.006109f
C335 B.n267 VSUBS 0.006109f
C336 B.n268 VSUBS 0.006109f
C337 B.n269 VSUBS 0.006109f
C338 B.n270 VSUBS 0.006109f
C339 B.n271 VSUBS 0.006109f
C340 B.n272 VSUBS 0.006109f
C341 B.n273 VSUBS 0.006109f
C342 B.n274 VSUBS 0.006109f
C343 B.n275 VSUBS 0.006109f
C344 B.n276 VSUBS 0.006109f
C345 B.n277 VSUBS 0.006109f
C346 B.n278 VSUBS 0.006109f
C347 B.n279 VSUBS 0.006109f
C348 B.n280 VSUBS 0.006109f
C349 B.n281 VSUBS 0.006109f
C350 B.n282 VSUBS 0.006109f
C351 B.n283 VSUBS 0.006109f
C352 B.n284 VSUBS 0.006109f
C353 B.n285 VSUBS 0.006109f
C354 B.n286 VSUBS 0.006109f
C355 B.n287 VSUBS 0.006109f
C356 B.n288 VSUBS 0.006109f
C357 B.n289 VSUBS 0.006109f
C358 B.n290 VSUBS 0.006109f
C359 B.n291 VSUBS 0.006109f
C360 B.n292 VSUBS 0.006109f
C361 B.n293 VSUBS 0.006109f
C362 B.n294 VSUBS 0.006109f
C363 B.n295 VSUBS 0.006109f
C364 B.n296 VSUBS 0.006109f
C365 B.n297 VSUBS 0.006109f
C366 B.n298 VSUBS 0.006109f
C367 B.n299 VSUBS 0.006109f
C368 B.n300 VSUBS 0.006109f
C369 B.n301 VSUBS 0.006109f
C370 B.n302 VSUBS 0.006109f
C371 B.n303 VSUBS 0.006109f
C372 B.n304 VSUBS 0.006109f
C373 B.n305 VSUBS 0.006109f
C374 B.n306 VSUBS 0.006109f
C375 B.n307 VSUBS 0.006109f
C376 B.n308 VSUBS 0.006109f
C377 B.n309 VSUBS 0.006109f
C378 B.n310 VSUBS 0.006109f
C379 B.n311 VSUBS 0.006109f
C380 B.n312 VSUBS 0.006109f
C381 B.n313 VSUBS 0.006109f
C382 B.n314 VSUBS 0.006109f
C383 B.n315 VSUBS 0.006109f
C384 B.n316 VSUBS 0.006109f
C385 B.n317 VSUBS 0.006109f
C386 B.n318 VSUBS 0.006109f
C387 B.n319 VSUBS 0.006109f
C388 B.n320 VSUBS 0.006109f
C389 B.n321 VSUBS 0.006109f
C390 B.n322 VSUBS 0.006109f
C391 B.n323 VSUBS 0.006109f
C392 B.n324 VSUBS 0.006109f
C393 B.n325 VSUBS 0.014099f
C394 B.n326 VSUBS 0.014469f
C395 B.n327 VSUBS 0.013746f
C396 B.n328 VSUBS 0.006109f
C397 B.n329 VSUBS 0.006109f
C398 B.n330 VSUBS 0.006109f
C399 B.n331 VSUBS 0.006109f
C400 B.n332 VSUBS 0.006109f
C401 B.n333 VSUBS 0.006109f
C402 B.n334 VSUBS 0.006109f
C403 B.n335 VSUBS 0.006109f
C404 B.n336 VSUBS 0.006109f
C405 B.n337 VSUBS 0.006109f
C406 B.n338 VSUBS 0.006109f
C407 B.n339 VSUBS 0.006109f
C408 B.n340 VSUBS 0.006109f
C409 B.n341 VSUBS 0.006109f
C410 B.n342 VSUBS 0.006109f
C411 B.n343 VSUBS 0.006109f
C412 B.n344 VSUBS 0.006109f
C413 B.n345 VSUBS 0.006109f
C414 B.n346 VSUBS 0.006109f
C415 B.n347 VSUBS 0.006109f
C416 B.n348 VSUBS 0.006109f
C417 B.n349 VSUBS 0.006109f
C418 B.n350 VSUBS 0.006109f
C419 B.n351 VSUBS 0.006109f
C420 B.n352 VSUBS 0.006109f
C421 B.n353 VSUBS 0.006109f
C422 B.n354 VSUBS 0.006109f
C423 B.n355 VSUBS 0.006109f
C424 B.n356 VSUBS 0.006109f
C425 B.n357 VSUBS 0.006109f
C426 B.n358 VSUBS 0.006109f
C427 B.n359 VSUBS 0.006109f
C428 B.n360 VSUBS 0.006109f
C429 B.n361 VSUBS 0.006109f
C430 B.n362 VSUBS 0.006109f
C431 B.n363 VSUBS 0.006109f
C432 B.n364 VSUBS 0.006109f
C433 B.n365 VSUBS 0.004222f
C434 B.n366 VSUBS 0.006109f
C435 B.n367 VSUBS 0.006109f
C436 B.n368 VSUBS 0.004941f
C437 B.n369 VSUBS 0.006109f
C438 B.n370 VSUBS 0.006109f
C439 B.n371 VSUBS 0.006109f
C440 B.n372 VSUBS 0.006109f
C441 B.n373 VSUBS 0.006109f
C442 B.n374 VSUBS 0.006109f
C443 B.n375 VSUBS 0.006109f
C444 B.n376 VSUBS 0.006109f
C445 B.n377 VSUBS 0.006109f
C446 B.n378 VSUBS 0.006109f
C447 B.n379 VSUBS 0.006109f
C448 B.n380 VSUBS 0.004941f
C449 B.n381 VSUBS 0.014154f
C450 B.n382 VSUBS 0.004222f
C451 B.n383 VSUBS 0.006109f
C452 B.n384 VSUBS 0.006109f
C453 B.n385 VSUBS 0.006109f
C454 B.n386 VSUBS 0.006109f
C455 B.n387 VSUBS 0.006109f
C456 B.n388 VSUBS 0.006109f
C457 B.n389 VSUBS 0.006109f
C458 B.n390 VSUBS 0.006109f
C459 B.n391 VSUBS 0.006109f
C460 B.n392 VSUBS 0.006109f
C461 B.n393 VSUBS 0.006109f
C462 B.n394 VSUBS 0.006109f
C463 B.n395 VSUBS 0.006109f
C464 B.n396 VSUBS 0.006109f
C465 B.n397 VSUBS 0.006109f
C466 B.n398 VSUBS 0.006109f
C467 B.n399 VSUBS 0.006109f
C468 B.n400 VSUBS 0.006109f
C469 B.n401 VSUBS 0.006109f
C470 B.n402 VSUBS 0.006109f
C471 B.n403 VSUBS 0.006109f
C472 B.n404 VSUBS 0.006109f
C473 B.n405 VSUBS 0.006109f
C474 B.n406 VSUBS 0.006109f
C475 B.n407 VSUBS 0.006109f
C476 B.n408 VSUBS 0.006109f
C477 B.n409 VSUBS 0.006109f
C478 B.n410 VSUBS 0.006109f
C479 B.n411 VSUBS 0.006109f
C480 B.n412 VSUBS 0.006109f
C481 B.n413 VSUBS 0.006109f
C482 B.n414 VSUBS 0.006109f
C483 B.n415 VSUBS 0.006109f
C484 B.n416 VSUBS 0.006109f
C485 B.n417 VSUBS 0.006109f
C486 B.n418 VSUBS 0.006109f
C487 B.n419 VSUBS 0.006109f
C488 B.n420 VSUBS 0.006109f
C489 B.n421 VSUBS 0.014469f
C490 B.n422 VSUBS 0.014099f
C491 B.n423 VSUBS 0.014099f
C492 B.n424 VSUBS 0.006109f
C493 B.n425 VSUBS 0.006109f
C494 B.n426 VSUBS 0.006109f
C495 B.n427 VSUBS 0.006109f
C496 B.n428 VSUBS 0.006109f
C497 B.n429 VSUBS 0.006109f
C498 B.n430 VSUBS 0.006109f
C499 B.n431 VSUBS 0.006109f
C500 B.n432 VSUBS 0.006109f
C501 B.n433 VSUBS 0.006109f
C502 B.n434 VSUBS 0.006109f
C503 B.n435 VSUBS 0.006109f
C504 B.n436 VSUBS 0.006109f
C505 B.n437 VSUBS 0.006109f
C506 B.n438 VSUBS 0.006109f
C507 B.n439 VSUBS 0.006109f
C508 B.n440 VSUBS 0.006109f
C509 B.n441 VSUBS 0.006109f
C510 B.n442 VSUBS 0.006109f
C511 B.n443 VSUBS 0.006109f
C512 B.n444 VSUBS 0.006109f
C513 B.n445 VSUBS 0.006109f
C514 B.n446 VSUBS 0.006109f
C515 B.n447 VSUBS 0.006109f
C516 B.n448 VSUBS 0.006109f
C517 B.n449 VSUBS 0.006109f
C518 B.n450 VSUBS 0.006109f
C519 B.n451 VSUBS 0.006109f
C520 B.n452 VSUBS 0.006109f
C521 B.n453 VSUBS 0.006109f
C522 B.n454 VSUBS 0.006109f
C523 B.n455 VSUBS 0.006109f
C524 B.n456 VSUBS 0.006109f
C525 B.n457 VSUBS 0.006109f
C526 B.n458 VSUBS 0.006109f
C527 B.n459 VSUBS 0.013833f
C528 VDD1.t5 VSUBS 1.14969f
C529 VDD1.t3 VSUBS 1.14897f
C530 VDD1.t2 VSUBS 0.125072f
C531 VDD1.t4 VSUBS 0.125072f
C532 VDD1.n0 VSUBS 0.860587f
C533 VDD1.n1 VSUBS 2.21343f
C534 VDD1.t1 VSUBS 0.125072f
C535 VDD1.t0 VSUBS 0.125072f
C536 VDD1.n2 VSUBS 0.859209f
C537 VDD1.n3 VSUBS 1.96755f
C538 VTAIL.t3 VSUBS 0.155406f
C539 VTAIL.t5 VSUBS 0.155406f
C540 VTAIL.n0 VSUBS 0.950749f
C541 VTAIL.n1 VSUBS 0.687949f
C542 VTAIL.t7 VSUBS 1.2966f
C543 VTAIL.n2 VSUBS 0.839306f
C544 VTAIL.t11 VSUBS 0.155406f
C545 VTAIL.t6 VSUBS 0.155406f
C546 VTAIL.n3 VSUBS 0.950749f
C547 VTAIL.n4 VSUBS 1.80497f
C548 VTAIL.t1 VSUBS 0.155406f
C549 VTAIL.t0 VSUBS 0.155406f
C550 VTAIL.n5 VSUBS 0.950754f
C551 VTAIL.n6 VSUBS 1.80497f
C552 VTAIL.t2 VSUBS 1.2966f
C553 VTAIL.n7 VSUBS 0.8393f
C554 VTAIL.t9 VSUBS 0.155406f
C555 VTAIL.t10 VSUBS 0.155406f
C556 VTAIL.n8 VSUBS 0.950754f
C557 VTAIL.n9 VSUBS 0.761316f
C558 VTAIL.t8 VSUBS 1.2966f
C559 VTAIL.n10 VSUBS 1.77808f
C560 VTAIL.t4 VSUBS 1.2966f
C561 VTAIL.n11 VSUBS 1.74658f
C562 VP.n0 VSUBS 0.075106f
C563 VP.t3 VSUBS 1.05892f
C564 VP.n1 VSUBS 0.065807f
C565 VP.n2 VSUBS 0.304217f
C566 VP.t5 VSUBS 1.14655f
C567 VP.t4 VSUBS 1.05892f
C568 VP.t0 VSUBS 1.19773f
C569 VP.n3 VSUBS 0.49022f
C570 VP.n4 VSUBS 0.510642f
C571 VP.n5 VSUBS 0.065807f
C572 VP.n6 VSUBS 0.507503f
C573 VP.n7 VSUBS 2.04237f
C574 VP.t2 VSUBS 1.14655f
C575 VP.n8 VSUBS 0.507503f
C576 VP.n9 VSUBS 2.09445f
C577 VP.n10 VSUBS 0.075106f
C578 VP.n11 VSUBS 0.056286f
C579 VP.n12 VSUBS 0.476105f
C580 VP.n13 VSUBS 0.065807f
C581 VP.t1 VSUBS 1.14655f
C582 VP.n14 VSUBS 0.507503f
C583 VP.n15 VSUBS 0.052714f
.ends

