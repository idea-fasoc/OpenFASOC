* NGSPICE file created from diff_pair_sample_1515.ext - technology: sky130A

.subckt diff_pair_sample_1515 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=6.0216 ps=31.66 w=15.44 l=1.53
X1 VTAIL.t15 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X2 VTAIL.t14 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=2.5476 ps=15.77 w=15.44 l=1.53
X3 VTAIL.t8 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X4 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X5 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=2.5476 ps=15.77 w=15.44 l=1.53
X6 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=0 ps=0 w=15.44 l=1.53
X7 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=6.0216 ps=31.66 w=15.44 l=1.53
X8 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X9 VDD1.t3 VP.t4 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=6.0216 ps=31.66 w=15.44 l=1.53
X10 VTAIL.t4 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X11 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X12 VDD1.t2 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X13 VDD1.t1 VP.t6 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=2.5476 ps=15.77 w=15.44 l=1.53
X14 VTAIL.t0 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=2.5476 ps=15.77 w=15.44 l=1.53
X15 VDD2.t0 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5476 pd=15.77 as=6.0216 ps=31.66 w=15.44 l=1.53
X16 VTAIL.t11 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=2.5476 ps=15.77 w=15.44 l=1.53
X17 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=0 ps=0 w=15.44 l=1.53
X18 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=0 ps=0 w=15.44 l=1.53
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.0216 pd=31.66 as=0 ps=0 w=15.44 l=1.53
R0 VP.n11 VP.t7 279.474
R1 VP.n25 VP.t2 243.206
R2 VP.n31 VP.t5 243.206
R3 VP.n38 VP.t1 243.206
R4 VP.n45 VP.t4 243.206
R5 VP.n23 VP.t0 243.206
R6 VP.n16 VP.t3 243.206
R7 VP.n10 VP.t6 243.206
R8 VP.n26 VP.n25 171.63
R9 VP.n46 VP.n45 171.63
R10 VP.n24 VP.n23 171.63
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n44 VP.n0 161.3
R19 VP.n43 VP.n42 161.3
R20 VP.n41 VP.n1 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n37 VP.n2 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n34 VP.n3 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n30 VP.n4 161.3
R27 VP.n29 VP.n28 161.3
R28 VP.n27 VP.n5 161.3
R29 VP.n30 VP.n29 54.1398
R30 VP.n43 VP.n1 54.1398
R31 VP.n21 VP.n7 54.1398
R32 VP.n26 VP.n24 48.4929
R33 VP.n11 VP.n10 45.6659
R34 VP.n36 VP.n3 40.577
R35 VP.n37 VP.n36 40.577
R36 VP.n15 VP.n14 40.577
R37 VP.n14 VP.n9 40.577
R38 VP.n29 VP.n5 27.0143
R39 VP.n44 VP.n43 27.0143
R40 VP.n22 VP.n21 27.0143
R41 VP.n32 VP.n30 24.5923
R42 VP.n39 VP.n1 24.5923
R43 VP.n17 VP.n7 24.5923
R44 VP.n31 VP.n3 21.1495
R45 VP.n38 VP.n37 21.1495
R46 VP.n16 VP.n15 21.1495
R47 VP.n10 VP.n9 21.1495
R48 VP.n12 VP.n11 17.3242
R49 VP.n25 VP.n5 14.2638
R50 VP.n45 VP.n44 14.2638
R51 VP.n23 VP.n22 14.2638
R52 VP.n32 VP.n31 3.44336
R53 VP.n39 VP.n38 3.44336
R54 VP.n17 VP.n16 3.44336
R55 VP.n13 VP.n12 0.189894
R56 VP.n13 VP.n8 0.189894
R57 VP.n18 VP.n8 0.189894
R58 VP.n19 VP.n18 0.189894
R59 VP.n20 VP.n19 0.189894
R60 VP.n20 VP.n6 0.189894
R61 VP.n24 VP.n6 0.189894
R62 VP.n27 VP.n26 0.189894
R63 VP.n28 VP.n27 0.189894
R64 VP.n28 VP.n4 0.189894
R65 VP.n33 VP.n4 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n35 VP.n34 0.189894
R68 VP.n35 VP.n2 0.189894
R69 VP.n40 VP.n2 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n42 VP.n41 0.189894
R72 VP.n42 VP.n0 0.189894
R73 VP.n46 VP.n0 0.189894
R74 VP VP.n46 0.0516364
R75 VTAIL.n690 VTAIL.n610 289.615
R76 VTAIL.n82 VTAIL.n2 289.615
R77 VTAIL.n168 VTAIL.n88 289.615
R78 VTAIL.n256 VTAIL.n176 289.615
R79 VTAIL.n604 VTAIL.n524 289.615
R80 VTAIL.n516 VTAIL.n436 289.615
R81 VTAIL.n430 VTAIL.n350 289.615
R82 VTAIL.n342 VTAIL.n262 289.615
R83 VTAIL.n639 VTAIL.n638 185
R84 VTAIL.n641 VTAIL.n640 185
R85 VTAIL.n634 VTAIL.n633 185
R86 VTAIL.n647 VTAIL.n646 185
R87 VTAIL.n649 VTAIL.n648 185
R88 VTAIL.n630 VTAIL.n629 185
R89 VTAIL.n655 VTAIL.n654 185
R90 VTAIL.n657 VTAIL.n656 185
R91 VTAIL.n626 VTAIL.n625 185
R92 VTAIL.n663 VTAIL.n662 185
R93 VTAIL.n665 VTAIL.n664 185
R94 VTAIL.n622 VTAIL.n621 185
R95 VTAIL.n671 VTAIL.n670 185
R96 VTAIL.n673 VTAIL.n672 185
R97 VTAIL.n618 VTAIL.n617 185
R98 VTAIL.n680 VTAIL.n679 185
R99 VTAIL.n681 VTAIL.n616 185
R100 VTAIL.n683 VTAIL.n682 185
R101 VTAIL.n614 VTAIL.n613 185
R102 VTAIL.n689 VTAIL.n688 185
R103 VTAIL.n691 VTAIL.n690 185
R104 VTAIL.n31 VTAIL.n30 185
R105 VTAIL.n33 VTAIL.n32 185
R106 VTAIL.n26 VTAIL.n25 185
R107 VTAIL.n39 VTAIL.n38 185
R108 VTAIL.n41 VTAIL.n40 185
R109 VTAIL.n22 VTAIL.n21 185
R110 VTAIL.n47 VTAIL.n46 185
R111 VTAIL.n49 VTAIL.n48 185
R112 VTAIL.n18 VTAIL.n17 185
R113 VTAIL.n55 VTAIL.n54 185
R114 VTAIL.n57 VTAIL.n56 185
R115 VTAIL.n14 VTAIL.n13 185
R116 VTAIL.n63 VTAIL.n62 185
R117 VTAIL.n65 VTAIL.n64 185
R118 VTAIL.n10 VTAIL.n9 185
R119 VTAIL.n72 VTAIL.n71 185
R120 VTAIL.n73 VTAIL.n8 185
R121 VTAIL.n75 VTAIL.n74 185
R122 VTAIL.n6 VTAIL.n5 185
R123 VTAIL.n81 VTAIL.n80 185
R124 VTAIL.n83 VTAIL.n82 185
R125 VTAIL.n117 VTAIL.n116 185
R126 VTAIL.n119 VTAIL.n118 185
R127 VTAIL.n112 VTAIL.n111 185
R128 VTAIL.n125 VTAIL.n124 185
R129 VTAIL.n127 VTAIL.n126 185
R130 VTAIL.n108 VTAIL.n107 185
R131 VTAIL.n133 VTAIL.n132 185
R132 VTAIL.n135 VTAIL.n134 185
R133 VTAIL.n104 VTAIL.n103 185
R134 VTAIL.n141 VTAIL.n140 185
R135 VTAIL.n143 VTAIL.n142 185
R136 VTAIL.n100 VTAIL.n99 185
R137 VTAIL.n149 VTAIL.n148 185
R138 VTAIL.n151 VTAIL.n150 185
R139 VTAIL.n96 VTAIL.n95 185
R140 VTAIL.n158 VTAIL.n157 185
R141 VTAIL.n159 VTAIL.n94 185
R142 VTAIL.n161 VTAIL.n160 185
R143 VTAIL.n92 VTAIL.n91 185
R144 VTAIL.n167 VTAIL.n166 185
R145 VTAIL.n169 VTAIL.n168 185
R146 VTAIL.n205 VTAIL.n204 185
R147 VTAIL.n207 VTAIL.n206 185
R148 VTAIL.n200 VTAIL.n199 185
R149 VTAIL.n213 VTAIL.n212 185
R150 VTAIL.n215 VTAIL.n214 185
R151 VTAIL.n196 VTAIL.n195 185
R152 VTAIL.n221 VTAIL.n220 185
R153 VTAIL.n223 VTAIL.n222 185
R154 VTAIL.n192 VTAIL.n191 185
R155 VTAIL.n229 VTAIL.n228 185
R156 VTAIL.n231 VTAIL.n230 185
R157 VTAIL.n188 VTAIL.n187 185
R158 VTAIL.n237 VTAIL.n236 185
R159 VTAIL.n239 VTAIL.n238 185
R160 VTAIL.n184 VTAIL.n183 185
R161 VTAIL.n246 VTAIL.n245 185
R162 VTAIL.n247 VTAIL.n182 185
R163 VTAIL.n249 VTAIL.n248 185
R164 VTAIL.n180 VTAIL.n179 185
R165 VTAIL.n255 VTAIL.n254 185
R166 VTAIL.n257 VTAIL.n256 185
R167 VTAIL.n605 VTAIL.n604 185
R168 VTAIL.n603 VTAIL.n602 185
R169 VTAIL.n528 VTAIL.n527 185
R170 VTAIL.n532 VTAIL.n530 185
R171 VTAIL.n597 VTAIL.n596 185
R172 VTAIL.n595 VTAIL.n594 185
R173 VTAIL.n534 VTAIL.n533 185
R174 VTAIL.n589 VTAIL.n588 185
R175 VTAIL.n587 VTAIL.n586 185
R176 VTAIL.n538 VTAIL.n537 185
R177 VTAIL.n581 VTAIL.n580 185
R178 VTAIL.n579 VTAIL.n578 185
R179 VTAIL.n542 VTAIL.n541 185
R180 VTAIL.n573 VTAIL.n572 185
R181 VTAIL.n571 VTAIL.n570 185
R182 VTAIL.n546 VTAIL.n545 185
R183 VTAIL.n565 VTAIL.n564 185
R184 VTAIL.n563 VTAIL.n562 185
R185 VTAIL.n550 VTAIL.n549 185
R186 VTAIL.n557 VTAIL.n556 185
R187 VTAIL.n555 VTAIL.n554 185
R188 VTAIL.n517 VTAIL.n516 185
R189 VTAIL.n515 VTAIL.n514 185
R190 VTAIL.n440 VTAIL.n439 185
R191 VTAIL.n444 VTAIL.n442 185
R192 VTAIL.n509 VTAIL.n508 185
R193 VTAIL.n507 VTAIL.n506 185
R194 VTAIL.n446 VTAIL.n445 185
R195 VTAIL.n501 VTAIL.n500 185
R196 VTAIL.n499 VTAIL.n498 185
R197 VTAIL.n450 VTAIL.n449 185
R198 VTAIL.n493 VTAIL.n492 185
R199 VTAIL.n491 VTAIL.n490 185
R200 VTAIL.n454 VTAIL.n453 185
R201 VTAIL.n485 VTAIL.n484 185
R202 VTAIL.n483 VTAIL.n482 185
R203 VTAIL.n458 VTAIL.n457 185
R204 VTAIL.n477 VTAIL.n476 185
R205 VTAIL.n475 VTAIL.n474 185
R206 VTAIL.n462 VTAIL.n461 185
R207 VTAIL.n469 VTAIL.n468 185
R208 VTAIL.n467 VTAIL.n466 185
R209 VTAIL.n431 VTAIL.n430 185
R210 VTAIL.n429 VTAIL.n428 185
R211 VTAIL.n354 VTAIL.n353 185
R212 VTAIL.n358 VTAIL.n356 185
R213 VTAIL.n423 VTAIL.n422 185
R214 VTAIL.n421 VTAIL.n420 185
R215 VTAIL.n360 VTAIL.n359 185
R216 VTAIL.n415 VTAIL.n414 185
R217 VTAIL.n413 VTAIL.n412 185
R218 VTAIL.n364 VTAIL.n363 185
R219 VTAIL.n407 VTAIL.n406 185
R220 VTAIL.n405 VTAIL.n404 185
R221 VTAIL.n368 VTAIL.n367 185
R222 VTAIL.n399 VTAIL.n398 185
R223 VTAIL.n397 VTAIL.n396 185
R224 VTAIL.n372 VTAIL.n371 185
R225 VTAIL.n391 VTAIL.n390 185
R226 VTAIL.n389 VTAIL.n388 185
R227 VTAIL.n376 VTAIL.n375 185
R228 VTAIL.n383 VTAIL.n382 185
R229 VTAIL.n381 VTAIL.n380 185
R230 VTAIL.n343 VTAIL.n342 185
R231 VTAIL.n341 VTAIL.n340 185
R232 VTAIL.n266 VTAIL.n265 185
R233 VTAIL.n270 VTAIL.n268 185
R234 VTAIL.n335 VTAIL.n334 185
R235 VTAIL.n333 VTAIL.n332 185
R236 VTAIL.n272 VTAIL.n271 185
R237 VTAIL.n327 VTAIL.n326 185
R238 VTAIL.n325 VTAIL.n324 185
R239 VTAIL.n276 VTAIL.n275 185
R240 VTAIL.n319 VTAIL.n318 185
R241 VTAIL.n317 VTAIL.n316 185
R242 VTAIL.n280 VTAIL.n279 185
R243 VTAIL.n311 VTAIL.n310 185
R244 VTAIL.n309 VTAIL.n308 185
R245 VTAIL.n284 VTAIL.n283 185
R246 VTAIL.n303 VTAIL.n302 185
R247 VTAIL.n301 VTAIL.n300 185
R248 VTAIL.n288 VTAIL.n287 185
R249 VTAIL.n295 VTAIL.n294 185
R250 VTAIL.n293 VTAIL.n292 185
R251 VTAIL.n637 VTAIL.t5 147.659
R252 VTAIL.n29 VTAIL.t0 147.659
R253 VTAIL.n115 VTAIL.t9 147.659
R254 VTAIL.n203 VTAIL.t14 147.659
R255 VTAIL.n553 VTAIL.t12 147.659
R256 VTAIL.n465 VTAIL.t11 147.659
R257 VTAIL.n379 VTAIL.t2 147.659
R258 VTAIL.n291 VTAIL.t7 147.659
R259 VTAIL.n640 VTAIL.n639 104.615
R260 VTAIL.n640 VTAIL.n633 104.615
R261 VTAIL.n647 VTAIL.n633 104.615
R262 VTAIL.n648 VTAIL.n647 104.615
R263 VTAIL.n648 VTAIL.n629 104.615
R264 VTAIL.n655 VTAIL.n629 104.615
R265 VTAIL.n656 VTAIL.n655 104.615
R266 VTAIL.n656 VTAIL.n625 104.615
R267 VTAIL.n663 VTAIL.n625 104.615
R268 VTAIL.n664 VTAIL.n663 104.615
R269 VTAIL.n664 VTAIL.n621 104.615
R270 VTAIL.n671 VTAIL.n621 104.615
R271 VTAIL.n672 VTAIL.n671 104.615
R272 VTAIL.n672 VTAIL.n617 104.615
R273 VTAIL.n680 VTAIL.n617 104.615
R274 VTAIL.n681 VTAIL.n680 104.615
R275 VTAIL.n682 VTAIL.n681 104.615
R276 VTAIL.n682 VTAIL.n613 104.615
R277 VTAIL.n689 VTAIL.n613 104.615
R278 VTAIL.n690 VTAIL.n689 104.615
R279 VTAIL.n32 VTAIL.n31 104.615
R280 VTAIL.n32 VTAIL.n25 104.615
R281 VTAIL.n39 VTAIL.n25 104.615
R282 VTAIL.n40 VTAIL.n39 104.615
R283 VTAIL.n40 VTAIL.n21 104.615
R284 VTAIL.n47 VTAIL.n21 104.615
R285 VTAIL.n48 VTAIL.n47 104.615
R286 VTAIL.n48 VTAIL.n17 104.615
R287 VTAIL.n55 VTAIL.n17 104.615
R288 VTAIL.n56 VTAIL.n55 104.615
R289 VTAIL.n56 VTAIL.n13 104.615
R290 VTAIL.n63 VTAIL.n13 104.615
R291 VTAIL.n64 VTAIL.n63 104.615
R292 VTAIL.n64 VTAIL.n9 104.615
R293 VTAIL.n72 VTAIL.n9 104.615
R294 VTAIL.n73 VTAIL.n72 104.615
R295 VTAIL.n74 VTAIL.n73 104.615
R296 VTAIL.n74 VTAIL.n5 104.615
R297 VTAIL.n81 VTAIL.n5 104.615
R298 VTAIL.n82 VTAIL.n81 104.615
R299 VTAIL.n118 VTAIL.n117 104.615
R300 VTAIL.n118 VTAIL.n111 104.615
R301 VTAIL.n125 VTAIL.n111 104.615
R302 VTAIL.n126 VTAIL.n125 104.615
R303 VTAIL.n126 VTAIL.n107 104.615
R304 VTAIL.n133 VTAIL.n107 104.615
R305 VTAIL.n134 VTAIL.n133 104.615
R306 VTAIL.n134 VTAIL.n103 104.615
R307 VTAIL.n141 VTAIL.n103 104.615
R308 VTAIL.n142 VTAIL.n141 104.615
R309 VTAIL.n142 VTAIL.n99 104.615
R310 VTAIL.n149 VTAIL.n99 104.615
R311 VTAIL.n150 VTAIL.n149 104.615
R312 VTAIL.n150 VTAIL.n95 104.615
R313 VTAIL.n158 VTAIL.n95 104.615
R314 VTAIL.n159 VTAIL.n158 104.615
R315 VTAIL.n160 VTAIL.n159 104.615
R316 VTAIL.n160 VTAIL.n91 104.615
R317 VTAIL.n167 VTAIL.n91 104.615
R318 VTAIL.n168 VTAIL.n167 104.615
R319 VTAIL.n206 VTAIL.n205 104.615
R320 VTAIL.n206 VTAIL.n199 104.615
R321 VTAIL.n213 VTAIL.n199 104.615
R322 VTAIL.n214 VTAIL.n213 104.615
R323 VTAIL.n214 VTAIL.n195 104.615
R324 VTAIL.n221 VTAIL.n195 104.615
R325 VTAIL.n222 VTAIL.n221 104.615
R326 VTAIL.n222 VTAIL.n191 104.615
R327 VTAIL.n229 VTAIL.n191 104.615
R328 VTAIL.n230 VTAIL.n229 104.615
R329 VTAIL.n230 VTAIL.n187 104.615
R330 VTAIL.n237 VTAIL.n187 104.615
R331 VTAIL.n238 VTAIL.n237 104.615
R332 VTAIL.n238 VTAIL.n183 104.615
R333 VTAIL.n246 VTAIL.n183 104.615
R334 VTAIL.n247 VTAIL.n246 104.615
R335 VTAIL.n248 VTAIL.n247 104.615
R336 VTAIL.n248 VTAIL.n179 104.615
R337 VTAIL.n255 VTAIL.n179 104.615
R338 VTAIL.n256 VTAIL.n255 104.615
R339 VTAIL.n604 VTAIL.n603 104.615
R340 VTAIL.n603 VTAIL.n527 104.615
R341 VTAIL.n532 VTAIL.n527 104.615
R342 VTAIL.n596 VTAIL.n532 104.615
R343 VTAIL.n596 VTAIL.n595 104.615
R344 VTAIL.n595 VTAIL.n533 104.615
R345 VTAIL.n588 VTAIL.n533 104.615
R346 VTAIL.n588 VTAIL.n587 104.615
R347 VTAIL.n587 VTAIL.n537 104.615
R348 VTAIL.n580 VTAIL.n537 104.615
R349 VTAIL.n580 VTAIL.n579 104.615
R350 VTAIL.n579 VTAIL.n541 104.615
R351 VTAIL.n572 VTAIL.n541 104.615
R352 VTAIL.n572 VTAIL.n571 104.615
R353 VTAIL.n571 VTAIL.n545 104.615
R354 VTAIL.n564 VTAIL.n545 104.615
R355 VTAIL.n564 VTAIL.n563 104.615
R356 VTAIL.n563 VTAIL.n549 104.615
R357 VTAIL.n556 VTAIL.n549 104.615
R358 VTAIL.n556 VTAIL.n555 104.615
R359 VTAIL.n516 VTAIL.n515 104.615
R360 VTAIL.n515 VTAIL.n439 104.615
R361 VTAIL.n444 VTAIL.n439 104.615
R362 VTAIL.n508 VTAIL.n444 104.615
R363 VTAIL.n508 VTAIL.n507 104.615
R364 VTAIL.n507 VTAIL.n445 104.615
R365 VTAIL.n500 VTAIL.n445 104.615
R366 VTAIL.n500 VTAIL.n499 104.615
R367 VTAIL.n499 VTAIL.n449 104.615
R368 VTAIL.n492 VTAIL.n449 104.615
R369 VTAIL.n492 VTAIL.n491 104.615
R370 VTAIL.n491 VTAIL.n453 104.615
R371 VTAIL.n484 VTAIL.n453 104.615
R372 VTAIL.n484 VTAIL.n483 104.615
R373 VTAIL.n483 VTAIL.n457 104.615
R374 VTAIL.n476 VTAIL.n457 104.615
R375 VTAIL.n476 VTAIL.n475 104.615
R376 VTAIL.n475 VTAIL.n461 104.615
R377 VTAIL.n468 VTAIL.n461 104.615
R378 VTAIL.n468 VTAIL.n467 104.615
R379 VTAIL.n430 VTAIL.n429 104.615
R380 VTAIL.n429 VTAIL.n353 104.615
R381 VTAIL.n358 VTAIL.n353 104.615
R382 VTAIL.n422 VTAIL.n358 104.615
R383 VTAIL.n422 VTAIL.n421 104.615
R384 VTAIL.n421 VTAIL.n359 104.615
R385 VTAIL.n414 VTAIL.n359 104.615
R386 VTAIL.n414 VTAIL.n413 104.615
R387 VTAIL.n413 VTAIL.n363 104.615
R388 VTAIL.n406 VTAIL.n363 104.615
R389 VTAIL.n406 VTAIL.n405 104.615
R390 VTAIL.n405 VTAIL.n367 104.615
R391 VTAIL.n398 VTAIL.n367 104.615
R392 VTAIL.n398 VTAIL.n397 104.615
R393 VTAIL.n397 VTAIL.n371 104.615
R394 VTAIL.n390 VTAIL.n371 104.615
R395 VTAIL.n390 VTAIL.n389 104.615
R396 VTAIL.n389 VTAIL.n375 104.615
R397 VTAIL.n382 VTAIL.n375 104.615
R398 VTAIL.n382 VTAIL.n381 104.615
R399 VTAIL.n342 VTAIL.n341 104.615
R400 VTAIL.n341 VTAIL.n265 104.615
R401 VTAIL.n270 VTAIL.n265 104.615
R402 VTAIL.n334 VTAIL.n270 104.615
R403 VTAIL.n334 VTAIL.n333 104.615
R404 VTAIL.n333 VTAIL.n271 104.615
R405 VTAIL.n326 VTAIL.n271 104.615
R406 VTAIL.n326 VTAIL.n325 104.615
R407 VTAIL.n325 VTAIL.n275 104.615
R408 VTAIL.n318 VTAIL.n275 104.615
R409 VTAIL.n318 VTAIL.n317 104.615
R410 VTAIL.n317 VTAIL.n279 104.615
R411 VTAIL.n310 VTAIL.n279 104.615
R412 VTAIL.n310 VTAIL.n309 104.615
R413 VTAIL.n309 VTAIL.n283 104.615
R414 VTAIL.n302 VTAIL.n283 104.615
R415 VTAIL.n302 VTAIL.n301 104.615
R416 VTAIL.n301 VTAIL.n287 104.615
R417 VTAIL.n294 VTAIL.n287 104.615
R418 VTAIL.n294 VTAIL.n293 104.615
R419 VTAIL.n639 VTAIL.t5 52.3082
R420 VTAIL.n31 VTAIL.t0 52.3082
R421 VTAIL.n117 VTAIL.t9 52.3082
R422 VTAIL.n205 VTAIL.t14 52.3082
R423 VTAIL.n555 VTAIL.t12 52.3082
R424 VTAIL.n467 VTAIL.t11 52.3082
R425 VTAIL.n381 VTAIL.t2 52.3082
R426 VTAIL.n293 VTAIL.t7 52.3082
R427 VTAIL.n523 VTAIL.n522 45.7153
R428 VTAIL.n349 VTAIL.n348 45.7153
R429 VTAIL.n1 VTAIL.n0 45.7151
R430 VTAIL.n175 VTAIL.n174 45.7151
R431 VTAIL.n695 VTAIL.n694 33.7369
R432 VTAIL.n87 VTAIL.n86 33.7369
R433 VTAIL.n173 VTAIL.n172 33.7369
R434 VTAIL.n261 VTAIL.n260 33.7369
R435 VTAIL.n609 VTAIL.n608 33.7369
R436 VTAIL.n521 VTAIL.n520 33.7369
R437 VTAIL.n435 VTAIL.n434 33.7369
R438 VTAIL.n347 VTAIL.n346 33.7369
R439 VTAIL.n695 VTAIL.n609 27.2807
R440 VTAIL.n347 VTAIL.n261 27.2807
R441 VTAIL.n638 VTAIL.n637 15.6677
R442 VTAIL.n30 VTAIL.n29 15.6677
R443 VTAIL.n116 VTAIL.n115 15.6677
R444 VTAIL.n204 VTAIL.n203 15.6677
R445 VTAIL.n554 VTAIL.n553 15.6677
R446 VTAIL.n466 VTAIL.n465 15.6677
R447 VTAIL.n380 VTAIL.n379 15.6677
R448 VTAIL.n292 VTAIL.n291 15.6677
R449 VTAIL.n683 VTAIL.n614 13.1884
R450 VTAIL.n75 VTAIL.n6 13.1884
R451 VTAIL.n161 VTAIL.n92 13.1884
R452 VTAIL.n249 VTAIL.n180 13.1884
R453 VTAIL.n530 VTAIL.n528 13.1884
R454 VTAIL.n442 VTAIL.n440 13.1884
R455 VTAIL.n356 VTAIL.n354 13.1884
R456 VTAIL.n268 VTAIL.n266 13.1884
R457 VTAIL.n641 VTAIL.n636 12.8005
R458 VTAIL.n684 VTAIL.n616 12.8005
R459 VTAIL.n688 VTAIL.n687 12.8005
R460 VTAIL.n33 VTAIL.n28 12.8005
R461 VTAIL.n76 VTAIL.n8 12.8005
R462 VTAIL.n80 VTAIL.n79 12.8005
R463 VTAIL.n119 VTAIL.n114 12.8005
R464 VTAIL.n162 VTAIL.n94 12.8005
R465 VTAIL.n166 VTAIL.n165 12.8005
R466 VTAIL.n207 VTAIL.n202 12.8005
R467 VTAIL.n250 VTAIL.n182 12.8005
R468 VTAIL.n254 VTAIL.n253 12.8005
R469 VTAIL.n602 VTAIL.n601 12.8005
R470 VTAIL.n598 VTAIL.n597 12.8005
R471 VTAIL.n557 VTAIL.n552 12.8005
R472 VTAIL.n514 VTAIL.n513 12.8005
R473 VTAIL.n510 VTAIL.n509 12.8005
R474 VTAIL.n469 VTAIL.n464 12.8005
R475 VTAIL.n428 VTAIL.n427 12.8005
R476 VTAIL.n424 VTAIL.n423 12.8005
R477 VTAIL.n383 VTAIL.n378 12.8005
R478 VTAIL.n340 VTAIL.n339 12.8005
R479 VTAIL.n336 VTAIL.n335 12.8005
R480 VTAIL.n295 VTAIL.n290 12.8005
R481 VTAIL.n642 VTAIL.n634 12.0247
R482 VTAIL.n679 VTAIL.n678 12.0247
R483 VTAIL.n691 VTAIL.n612 12.0247
R484 VTAIL.n34 VTAIL.n26 12.0247
R485 VTAIL.n71 VTAIL.n70 12.0247
R486 VTAIL.n83 VTAIL.n4 12.0247
R487 VTAIL.n120 VTAIL.n112 12.0247
R488 VTAIL.n157 VTAIL.n156 12.0247
R489 VTAIL.n169 VTAIL.n90 12.0247
R490 VTAIL.n208 VTAIL.n200 12.0247
R491 VTAIL.n245 VTAIL.n244 12.0247
R492 VTAIL.n257 VTAIL.n178 12.0247
R493 VTAIL.n605 VTAIL.n526 12.0247
R494 VTAIL.n594 VTAIL.n531 12.0247
R495 VTAIL.n558 VTAIL.n550 12.0247
R496 VTAIL.n517 VTAIL.n438 12.0247
R497 VTAIL.n506 VTAIL.n443 12.0247
R498 VTAIL.n470 VTAIL.n462 12.0247
R499 VTAIL.n431 VTAIL.n352 12.0247
R500 VTAIL.n420 VTAIL.n357 12.0247
R501 VTAIL.n384 VTAIL.n376 12.0247
R502 VTAIL.n343 VTAIL.n264 12.0247
R503 VTAIL.n332 VTAIL.n269 12.0247
R504 VTAIL.n296 VTAIL.n288 12.0247
R505 VTAIL.n646 VTAIL.n645 11.249
R506 VTAIL.n677 VTAIL.n618 11.249
R507 VTAIL.n692 VTAIL.n610 11.249
R508 VTAIL.n38 VTAIL.n37 11.249
R509 VTAIL.n69 VTAIL.n10 11.249
R510 VTAIL.n84 VTAIL.n2 11.249
R511 VTAIL.n124 VTAIL.n123 11.249
R512 VTAIL.n155 VTAIL.n96 11.249
R513 VTAIL.n170 VTAIL.n88 11.249
R514 VTAIL.n212 VTAIL.n211 11.249
R515 VTAIL.n243 VTAIL.n184 11.249
R516 VTAIL.n258 VTAIL.n176 11.249
R517 VTAIL.n606 VTAIL.n524 11.249
R518 VTAIL.n593 VTAIL.n534 11.249
R519 VTAIL.n562 VTAIL.n561 11.249
R520 VTAIL.n518 VTAIL.n436 11.249
R521 VTAIL.n505 VTAIL.n446 11.249
R522 VTAIL.n474 VTAIL.n473 11.249
R523 VTAIL.n432 VTAIL.n350 11.249
R524 VTAIL.n419 VTAIL.n360 11.249
R525 VTAIL.n388 VTAIL.n387 11.249
R526 VTAIL.n344 VTAIL.n262 11.249
R527 VTAIL.n331 VTAIL.n272 11.249
R528 VTAIL.n300 VTAIL.n299 11.249
R529 VTAIL.n649 VTAIL.n632 10.4732
R530 VTAIL.n674 VTAIL.n673 10.4732
R531 VTAIL.n41 VTAIL.n24 10.4732
R532 VTAIL.n66 VTAIL.n65 10.4732
R533 VTAIL.n127 VTAIL.n110 10.4732
R534 VTAIL.n152 VTAIL.n151 10.4732
R535 VTAIL.n215 VTAIL.n198 10.4732
R536 VTAIL.n240 VTAIL.n239 10.4732
R537 VTAIL.n590 VTAIL.n589 10.4732
R538 VTAIL.n565 VTAIL.n548 10.4732
R539 VTAIL.n502 VTAIL.n501 10.4732
R540 VTAIL.n477 VTAIL.n460 10.4732
R541 VTAIL.n416 VTAIL.n415 10.4732
R542 VTAIL.n391 VTAIL.n374 10.4732
R543 VTAIL.n328 VTAIL.n327 10.4732
R544 VTAIL.n303 VTAIL.n286 10.4732
R545 VTAIL.n650 VTAIL.n630 9.69747
R546 VTAIL.n670 VTAIL.n620 9.69747
R547 VTAIL.n42 VTAIL.n22 9.69747
R548 VTAIL.n62 VTAIL.n12 9.69747
R549 VTAIL.n128 VTAIL.n108 9.69747
R550 VTAIL.n148 VTAIL.n98 9.69747
R551 VTAIL.n216 VTAIL.n196 9.69747
R552 VTAIL.n236 VTAIL.n186 9.69747
R553 VTAIL.n586 VTAIL.n536 9.69747
R554 VTAIL.n566 VTAIL.n546 9.69747
R555 VTAIL.n498 VTAIL.n448 9.69747
R556 VTAIL.n478 VTAIL.n458 9.69747
R557 VTAIL.n412 VTAIL.n362 9.69747
R558 VTAIL.n392 VTAIL.n372 9.69747
R559 VTAIL.n324 VTAIL.n274 9.69747
R560 VTAIL.n304 VTAIL.n284 9.69747
R561 VTAIL.n694 VTAIL.n693 9.45567
R562 VTAIL.n86 VTAIL.n85 9.45567
R563 VTAIL.n172 VTAIL.n171 9.45567
R564 VTAIL.n260 VTAIL.n259 9.45567
R565 VTAIL.n608 VTAIL.n607 9.45567
R566 VTAIL.n520 VTAIL.n519 9.45567
R567 VTAIL.n434 VTAIL.n433 9.45567
R568 VTAIL.n346 VTAIL.n345 9.45567
R569 VTAIL.n693 VTAIL.n692 9.3005
R570 VTAIL.n612 VTAIL.n611 9.3005
R571 VTAIL.n687 VTAIL.n686 9.3005
R572 VTAIL.n659 VTAIL.n658 9.3005
R573 VTAIL.n628 VTAIL.n627 9.3005
R574 VTAIL.n653 VTAIL.n652 9.3005
R575 VTAIL.n651 VTAIL.n650 9.3005
R576 VTAIL.n632 VTAIL.n631 9.3005
R577 VTAIL.n645 VTAIL.n644 9.3005
R578 VTAIL.n643 VTAIL.n642 9.3005
R579 VTAIL.n636 VTAIL.n635 9.3005
R580 VTAIL.n661 VTAIL.n660 9.3005
R581 VTAIL.n624 VTAIL.n623 9.3005
R582 VTAIL.n667 VTAIL.n666 9.3005
R583 VTAIL.n669 VTAIL.n668 9.3005
R584 VTAIL.n620 VTAIL.n619 9.3005
R585 VTAIL.n675 VTAIL.n674 9.3005
R586 VTAIL.n677 VTAIL.n676 9.3005
R587 VTAIL.n678 VTAIL.n615 9.3005
R588 VTAIL.n685 VTAIL.n684 9.3005
R589 VTAIL.n85 VTAIL.n84 9.3005
R590 VTAIL.n4 VTAIL.n3 9.3005
R591 VTAIL.n79 VTAIL.n78 9.3005
R592 VTAIL.n51 VTAIL.n50 9.3005
R593 VTAIL.n20 VTAIL.n19 9.3005
R594 VTAIL.n45 VTAIL.n44 9.3005
R595 VTAIL.n43 VTAIL.n42 9.3005
R596 VTAIL.n24 VTAIL.n23 9.3005
R597 VTAIL.n37 VTAIL.n36 9.3005
R598 VTAIL.n35 VTAIL.n34 9.3005
R599 VTAIL.n28 VTAIL.n27 9.3005
R600 VTAIL.n53 VTAIL.n52 9.3005
R601 VTAIL.n16 VTAIL.n15 9.3005
R602 VTAIL.n59 VTAIL.n58 9.3005
R603 VTAIL.n61 VTAIL.n60 9.3005
R604 VTAIL.n12 VTAIL.n11 9.3005
R605 VTAIL.n67 VTAIL.n66 9.3005
R606 VTAIL.n69 VTAIL.n68 9.3005
R607 VTAIL.n70 VTAIL.n7 9.3005
R608 VTAIL.n77 VTAIL.n76 9.3005
R609 VTAIL.n171 VTAIL.n170 9.3005
R610 VTAIL.n90 VTAIL.n89 9.3005
R611 VTAIL.n165 VTAIL.n164 9.3005
R612 VTAIL.n137 VTAIL.n136 9.3005
R613 VTAIL.n106 VTAIL.n105 9.3005
R614 VTAIL.n131 VTAIL.n130 9.3005
R615 VTAIL.n129 VTAIL.n128 9.3005
R616 VTAIL.n110 VTAIL.n109 9.3005
R617 VTAIL.n123 VTAIL.n122 9.3005
R618 VTAIL.n121 VTAIL.n120 9.3005
R619 VTAIL.n114 VTAIL.n113 9.3005
R620 VTAIL.n139 VTAIL.n138 9.3005
R621 VTAIL.n102 VTAIL.n101 9.3005
R622 VTAIL.n145 VTAIL.n144 9.3005
R623 VTAIL.n147 VTAIL.n146 9.3005
R624 VTAIL.n98 VTAIL.n97 9.3005
R625 VTAIL.n153 VTAIL.n152 9.3005
R626 VTAIL.n155 VTAIL.n154 9.3005
R627 VTAIL.n156 VTAIL.n93 9.3005
R628 VTAIL.n163 VTAIL.n162 9.3005
R629 VTAIL.n259 VTAIL.n258 9.3005
R630 VTAIL.n178 VTAIL.n177 9.3005
R631 VTAIL.n253 VTAIL.n252 9.3005
R632 VTAIL.n225 VTAIL.n224 9.3005
R633 VTAIL.n194 VTAIL.n193 9.3005
R634 VTAIL.n219 VTAIL.n218 9.3005
R635 VTAIL.n217 VTAIL.n216 9.3005
R636 VTAIL.n198 VTAIL.n197 9.3005
R637 VTAIL.n211 VTAIL.n210 9.3005
R638 VTAIL.n209 VTAIL.n208 9.3005
R639 VTAIL.n202 VTAIL.n201 9.3005
R640 VTAIL.n227 VTAIL.n226 9.3005
R641 VTAIL.n190 VTAIL.n189 9.3005
R642 VTAIL.n233 VTAIL.n232 9.3005
R643 VTAIL.n235 VTAIL.n234 9.3005
R644 VTAIL.n186 VTAIL.n185 9.3005
R645 VTAIL.n241 VTAIL.n240 9.3005
R646 VTAIL.n243 VTAIL.n242 9.3005
R647 VTAIL.n244 VTAIL.n181 9.3005
R648 VTAIL.n251 VTAIL.n250 9.3005
R649 VTAIL.n540 VTAIL.n539 9.3005
R650 VTAIL.n583 VTAIL.n582 9.3005
R651 VTAIL.n585 VTAIL.n584 9.3005
R652 VTAIL.n536 VTAIL.n535 9.3005
R653 VTAIL.n591 VTAIL.n590 9.3005
R654 VTAIL.n593 VTAIL.n592 9.3005
R655 VTAIL.n531 VTAIL.n529 9.3005
R656 VTAIL.n599 VTAIL.n598 9.3005
R657 VTAIL.n607 VTAIL.n606 9.3005
R658 VTAIL.n526 VTAIL.n525 9.3005
R659 VTAIL.n601 VTAIL.n600 9.3005
R660 VTAIL.n577 VTAIL.n576 9.3005
R661 VTAIL.n575 VTAIL.n574 9.3005
R662 VTAIL.n544 VTAIL.n543 9.3005
R663 VTAIL.n569 VTAIL.n568 9.3005
R664 VTAIL.n567 VTAIL.n566 9.3005
R665 VTAIL.n548 VTAIL.n547 9.3005
R666 VTAIL.n561 VTAIL.n560 9.3005
R667 VTAIL.n559 VTAIL.n558 9.3005
R668 VTAIL.n552 VTAIL.n551 9.3005
R669 VTAIL.n452 VTAIL.n451 9.3005
R670 VTAIL.n495 VTAIL.n494 9.3005
R671 VTAIL.n497 VTAIL.n496 9.3005
R672 VTAIL.n448 VTAIL.n447 9.3005
R673 VTAIL.n503 VTAIL.n502 9.3005
R674 VTAIL.n505 VTAIL.n504 9.3005
R675 VTAIL.n443 VTAIL.n441 9.3005
R676 VTAIL.n511 VTAIL.n510 9.3005
R677 VTAIL.n519 VTAIL.n518 9.3005
R678 VTAIL.n438 VTAIL.n437 9.3005
R679 VTAIL.n513 VTAIL.n512 9.3005
R680 VTAIL.n489 VTAIL.n488 9.3005
R681 VTAIL.n487 VTAIL.n486 9.3005
R682 VTAIL.n456 VTAIL.n455 9.3005
R683 VTAIL.n481 VTAIL.n480 9.3005
R684 VTAIL.n479 VTAIL.n478 9.3005
R685 VTAIL.n460 VTAIL.n459 9.3005
R686 VTAIL.n473 VTAIL.n472 9.3005
R687 VTAIL.n471 VTAIL.n470 9.3005
R688 VTAIL.n464 VTAIL.n463 9.3005
R689 VTAIL.n366 VTAIL.n365 9.3005
R690 VTAIL.n409 VTAIL.n408 9.3005
R691 VTAIL.n411 VTAIL.n410 9.3005
R692 VTAIL.n362 VTAIL.n361 9.3005
R693 VTAIL.n417 VTAIL.n416 9.3005
R694 VTAIL.n419 VTAIL.n418 9.3005
R695 VTAIL.n357 VTAIL.n355 9.3005
R696 VTAIL.n425 VTAIL.n424 9.3005
R697 VTAIL.n433 VTAIL.n432 9.3005
R698 VTAIL.n352 VTAIL.n351 9.3005
R699 VTAIL.n427 VTAIL.n426 9.3005
R700 VTAIL.n403 VTAIL.n402 9.3005
R701 VTAIL.n401 VTAIL.n400 9.3005
R702 VTAIL.n370 VTAIL.n369 9.3005
R703 VTAIL.n395 VTAIL.n394 9.3005
R704 VTAIL.n393 VTAIL.n392 9.3005
R705 VTAIL.n374 VTAIL.n373 9.3005
R706 VTAIL.n387 VTAIL.n386 9.3005
R707 VTAIL.n385 VTAIL.n384 9.3005
R708 VTAIL.n378 VTAIL.n377 9.3005
R709 VTAIL.n278 VTAIL.n277 9.3005
R710 VTAIL.n321 VTAIL.n320 9.3005
R711 VTAIL.n323 VTAIL.n322 9.3005
R712 VTAIL.n274 VTAIL.n273 9.3005
R713 VTAIL.n329 VTAIL.n328 9.3005
R714 VTAIL.n331 VTAIL.n330 9.3005
R715 VTAIL.n269 VTAIL.n267 9.3005
R716 VTAIL.n337 VTAIL.n336 9.3005
R717 VTAIL.n345 VTAIL.n344 9.3005
R718 VTAIL.n264 VTAIL.n263 9.3005
R719 VTAIL.n339 VTAIL.n338 9.3005
R720 VTAIL.n315 VTAIL.n314 9.3005
R721 VTAIL.n313 VTAIL.n312 9.3005
R722 VTAIL.n282 VTAIL.n281 9.3005
R723 VTAIL.n307 VTAIL.n306 9.3005
R724 VTAIL.n305 VTAIL.n304 9.3005
R725 VTAIL.n286 VTAIL.n285 9.3005
R726 VTAIL.n299 VTAIL.n298 9.3005
R727 VTAIL.n297 VTAIL.n296 9.3005
R728 VTAIL.n290 VTAIL.n289 9.3005
R729 VTAIL.n654 VTAIL.n653 8.92171
R730 VTAIL.n669 VTAIL.n622 8.92171
R731 VTAIL.n46 VTAIL.n45 8.92171
R732 VTAIL.n61 VTAIL.n14 8.92171
R733 VTAIL.n132 VTAIL.n131 8.92171
R734 VTAIL.n147 VTAIL.n100 8.92171
R735 VTAIL.n220 VTAIL.n219 8.92171
R736 VTAIL.n235 VTAIL.n188 8.92171
R737 VTAIL.n585 VTAIL.n538 8.92171
R738 VTAIL.n570 VTAIL.n569 8.92171
R739 VTAIL.n497 VTAIL.n450 8.92171
R740 VTAIL.n482 VTAIL.n481 8.92171
R741 VTAIL.n411 VTAIL.n364 8.92171
R742 VTAIL.n396 VTAIL.n395 8.92171
R743 VTAIL.n323 VTAIL.n276 8.92171
R744 VTAIL.n308 VTAIL.n307 8.92171
R745 VTAIL.n657 VTAIL.n628 8.14595
R746 VTAIL.n666 VTAIL.n665 8.14595
R747 VTAIL.n49 VTAIL.n20 8.14595
R748 VTAIL.n58 VTAIL.n57 8.14595
R749 VTAIL.n135 VTAIL.n106 8.14595
R750 VTAIL.n144 VTAIL.n143 8.14595
R751 VTAIL.n223 VTAIL.n194 8.14595
R752 VTAIL.n232 VTAIL.n231 8.14595
R753 VTAIL.n582 VTAIL.n581 8.14595
R754 VTAIL.n573 VTAIL.n544 8.14595
R755 VTAIL.n494 VTAIL.n493 8.14595
R756 VTAIL.n485 VTAIL.n456 8.14595
R757 VTAIL.n408 VTAIL.n407 8.14595
R758 VTAIL.n399 VTAIL.n370 8.14595
R759 VTAIL.n320 VTAIL.n319 8.14595
R760 VTAIL.n311 VTAIL.n282 8.14595
R761 VTAIL.n658 VTAIL.n626 7.3702
R762 VTAIL.n662 VTAIL.n624 7.3702
R763 VTAIL.n50 VTAIL.n18 7.3702
R764 VTAIL.n54 VTAIL.n16 7.3702
R765 VTAIL.n136 VTAIL.n104 7.3702
R766 VTAIL.n140 VTAIL.n102 7.3702
R767 VTAIL.n224 VTAIL.n192 7.3702
R768 VTAIL.n228 VTAIL.n190 7.3702
R769 VTAIL.n578 VTAIL.n540 7.3702
R770 VTAIL.n574 VTAIL.n542 7.3702
R771 VTAIL.n490 VTAIL.n452 7.3702
R772 VTAIL.n486 VTAIL.n454 7.3702
R773 VTAIL.n404 VTAIL.n366 7.3702
R774 VTAIL.n400 VTAIL.n368 7.3702
R775 VTAIL.n316 VTAIL.n278 7.3702
R776 VTAIL.n312 VTAIL.n280 7.3702
R777 VTAIL.n661 VTAIL.n626 6.59444
R778 VTAIL.n662 VTAIL.n661 6.59444
R779 VTAIL.n53 VTAIL.n18 6.59444
R780 VTAIL.n54 VTAIL.n53 6.59444
R781 VTAIL.n139 VTAIL.n104 6.59444
R782 VTAIL.n140 VTAIL.n139 6.59444
R783 VTAIL.n227 VTAIL.n192 6.59444
R784 VTAIL.n228 VTAIL.n227 6.59444
R785 VTAIL.n578 VTAIL.n577 6.59444
R786 VTAIL.n577 VTAIL.n542 6.59444
R787 VTAIL.n490 VTAIL.n489 6.59444
R788 VTAIL.n489 VTAIL.n454 6.59444
R789 VTAIL.n404 VTAIL.n403 6.59444
R790 VTAIL.n403 VTAIL.n368 6.59444
R791 VTAIL.n316 VTAIL.n315 6.59444
R792 VTAIL.n315 VTAIL.n280 6.59444
R793 VTAIL.n658 VTAIL.n657 5.81868
R794 VTAIL.n665 VTAIL.n624 5.81868
R795 VTAIL.n50 VTAIL.n49 5.81868
R796 VTAIL.n57 VTAIL.n16 5.81868
R797 VTAIL.n136 VTAIL.n135 5.81868
R798 VTAIL.n143 VTAIL.n102 5.81868
R799 VTAIL.n224 VTAIL.n223 5.81868
R800 VTAIL.n231 VTAIL.n190 5.81868
R801 VTAIL.n581 VTAIL.n540 5.81868
R802 VTAIL.n574 VTAIL.n573 5.81868
R803 VTAIL.n493 VTAIL.n452 5.81868
R804 VTAIL.n486 VTAIL.n485 5.81868
R805 VTAIL.n407 VTAIL.n366 5.81868
R806 VTAIL.n400 VTAIL.n399 5.81868
R807 VTAIL.n319 VTAIL.n278 5.81868
R808 VTAIL.n312 VTAIL.n311 5.81868
R809 VTAIL.n654 VTAIL.n628 5.04292
R810 VTAIL.n666 VTAIL.n622 5.04292
R811 VTAIL.n46 VTAIL.n20 5.04292
R812 VTAIL.n58 VTAIL.n14 5.04292
R813 VTAIL.n132 VTAIL.n106 5.04292
R814 VTAIL.n144 VTAIL.n100 5.04292
R815 VTAIL.n220 VTAIL.n194 5.04292
R816 VTAIL.n232 VTAIL.n188 5.04292
R817 VTAIL.n582 VTAIL.n538 5.04292
R818 VTAIL.n570 VTAIL.n544 5.04292
R819 VTAIL.n494 VTAIL.n450 5.04292
R820 VTAIL.n482 VTAIL.n456 5.04292
R821 VTAIL.n408 VTAIL.n364 5.04292
R822 VTAIL.n396 VTAIL.n370 5.04292
R823 VTAIL.n320 VTAIL.n276 5.04292
R824 VTAIL.n308 VTAIL.n282 5.04292
R825 VTAIL.n637 VTAIL.n635 4.38563
R826 VTAIL.n29 VTAIL.n27 4.38563
R827 VTAIL.n115 VTAIL.n113 4.38563
R828 VTAIL.n203 VTAIL.n201 4.38563
R829 VTAIL.n553 VTAIL.n551 4.38563
R830 VTAIL.n465 VTAIL.n463 4.38563
R831 VTAIL.n379 VTAIL.n377 4.38563
R832 VTAIL.n291 VTAIL.n289 4.38563
R833 VTAIL.n653 VTAIL.n630 4.26717
R834 VTAIL.n670 VTAIL.n669 4.26717
R835 VTAIL.n45 VTAIL.n22 4.26717
R836 VTAIL.n62 VTAIL.n61 4.26717
R837 VTAIL.n131 VTAIL.n108 4.26717
R838 VTAIL.n148 VTAIL.n147 4.26717
R839 VTAIL.n219 VTAIL.n196 4.26717
R840 VTAIL.n236 VTAIL.n235 4.26717
R841 VTAIL.n586 VTAIL.n585 4.26717
R842 VTAIL.n569 VTAIL.n546 4.26717
R843 VTAIL.n498 VTAIL.n497 4.26717
R844 VTAIL.n481 VTAIL.n458 4.26717
R845 VTAIL.n412 VTAIL.n411 4.26717
R846 VTAIL.n395 VTAIL.n372 4.26717
R847 VTAIL.n324 VTAIL.n323 4.26717
R848 VTAIL.n307 VTAIL.n284 4.26717
R849 VTAIL.n650 VTAIL.n649 3.49141
R850 VTAIL.n673 VTAIL.n620 3.49141
R851 VTAIL.n42 VTAIL.n41 3.49141
R852 VTAIL.n65 VTAIL.n12 3.49141
R853 VTAIL.n128 VTAIL.n127 3.49141
R854 VTAIL.n151 VTAIL.n98 3.49141
R855 VTAIL.n216 VTAIL.n215 3.49141
R856 VTAIL.n239 VTAIL.n186 3.49141
R857 VTAIL.n589 VTAIL.n536 3.49141
R858 VTAIL.n566 VTAIL.n565 3.49141
R859 VTAIL.n501 VTAIL.n448 3.49141
R860 VTAIL.n478 VTAIL.n477 3.49141
R861 VTAIL.n415 VTAIL.n362 3.49141
R862 VTAIL.n392 VTAIL.n391 3.49141
R863 VTAIL.n327 VTAIL.n274 3.49141
R864 VTAIL.n304 VTAIL.n303 3.49141
R865 VTAIL.n646 VTAIL.n632 2.71565
R866 VTAIL.n674 VTAIL.n618 2.71565
R867 VTAIL.n694 VTAIL.n610 2.71565
R868 VTAIL.n38 VTAIL.n24 2.71565
R869 VTAIL.n66 VTAIL.n10 2.71565
R870 VTAIL.n86 VTAIL.n2 2.71565
R871 VTAIL.n124 VTAIL.n110 2.71565
R872 VTAIL.n152 VTAIL.n96 2.71565
R873 VTAIL.n172 VTAIL.n88 2.71565
R874 VTAIL.n212 VTAIL.n198 2.71565
R875 VTAIL.n240 VTAIL.n184 2.71565
R876 VTAIL.n260 VTAIL.n176 2.71565
R877 VTAIL.n608 VTAIL.n524 2.71565
R878 VTAIL.n590 VTAIL.n534 2.71565
R879 VTAIL.n562 VTAIL.n548 2.71565
R880 VTAIL.n520 VTAIL.n436 2.71565
R881 VTAIL.n502 VTAIL.n446 2.71565
R882 VTAIL.n474 VTAIL.n460 2.71565
R883 VTAIL.n434 VTAIL.n350 2.71565
R884 VTAIL.n416 VTAIL.n360 2.71565
R885 VTAIL.n388 VTAIL.n374 2.71565
R886 VTAIL.n346 VTAIL.n262 2.71565
R887 VTAIL.n328 VTAIL.n272 2.71565
R888 VTAIL.n300 VTAIL.n286 2.71565
R889 VTAIL.n645 VTAIL.n634 1.93989
R890 VTAIL.n679 VTAIL.n677 1.93989
R891 VTAIL.n692 VTAIL.n691 1.93989
R892 VTAIL.n37 VTAIL.n26 1.93989
R893 VTAIL.n71 VTAIL.n69 1.93989
R894 VTAIL.n84 VTAIL.n83 1.93989
R895 VTAIL.n123 VTAIL.n112 1.93989
R896 VTAIL.n157 VTAIL.n155 1.93989
R897 VTAIL.n170 VTAIL.n169 1.93989
R898 VTAIL.n211 VTAIL.n200 1.93989
R899 VTAIL.n245 VTAIL.n243 1.93989
R900 VTAIL.n258 VTAIL.n257 1.93989
R901 VTAIL.n606 VTAIL.n605 1.93989
R902 VTAIL.n594 VTAIL.n593 1.93989
R903 VTAIL.n561 VTAIL.n550 1.93989
R904 VTAIL.n518 VTAIL.n517 1.93989
R905 VTAIL.n506 VTAIL.n505 1.93989
R906 VTAIL.n473 VTAIL.n462 1.93989
R907 VTAIL.n432 VTAIL.n431 1.93989
R908 VTAIL.n420 VTAIL.n419 1.93989
R909 VTAIL.n387 VTAIL.n376 1.93989
R910 VTAIL.n344 VTAIL.n343 1.93989
R911 VTAIL.n332 VTAIL.n331 1.93989
R912 VTAIL.n299 VTAIL.n288 1.93989
R913 VTAIL.n349 VTAIL.n347 1.60395
R914 VTAIL.n435 VTAIL.n349 1.60395
R915 VTAIL.n523 VTAIL.n521 1.60395
R916 VTAIL.n609 VTAIL.n523 1.60395
R917 VTAIL.n261 VTAIL.n175 1.60395
R918 VTAIL.n175 VTAIL.n173 1.60395
R919 VTAIL.n87 VTAIL.n1 1.60395
R920 VTAIL VTAIL.n695 1.54576
R921 VTAIL.n0 VTAIL.t3 1.28288
R922 VTAIL.n0 VTAIL.t4 1.28288
R923 VTAIL.n174 VTAIL.t10 1.28288
R924 VTAIL.n174 VTAIL.t15 1.28288
R925 VTAIL.n522 VTAIL.t13 1.28288
R926 VTAIL.n522 VTAIL.t8 1.28288
R927 VTAIL.n348 VTAIL.t6 1.28288
R928 VTAIL.n348 VTAIL.t1 1.28288
R929 VTAIL.n642 VTAIL.n641 1.16414
R930 VTAIL.n678 VTAIL.n616 1.16414
R931 VTAIL.n688 VTAIL.n612 1.16414
R932 VTAIL.n34 VTAIL.n33 1.16414
R933 VTAIL.n70 VTAIL.n8 1.16414
R934 VTAIL.n80 VTAIL.n4 1.16414
R935 VTAIL.n120 VTAIL.n119 1.16414
R936 VTAIL.n156 VTAIL.n94 1.16414
R937 VTAIL.n166 VTAIL.n90 1.16414
R938 VTAIL.n208 VTAIL.n207 1.16414
R939 VTAIL.n244 VTAIL.n182 1.16414
R940 VTAIL.n254 VTAIL.n178 1.16414
R941 VTAIL.n602 VTAIL.n526 1.16414
R942 VTAIL.n597 VTAIL.n531 1.16414
R943 VTAIL.n558 VTAIL.n557 1.16414
R944 VTAIL.n514 VTAIL.n438 1.16414
R945 VTAIL.n509 VTAIL.n443 1.16414
R946 VTAIL.n470 VTAIL.n469 1.16414
R947 VTAIL.n428 VTAIL.n352 1.16414
R948 VTAIL.n423 VTAIL.n357 1.16414
R949 VTAIL.n384 VTAIL.n383 1.16414
R950 VTAIL.n340 VTAIL.n264 1.16414
R951 VTAIL.n335 VTAIL.n269 1.16414
R952 VTAIL.n296 VTAIL.n295 1.16414
R953 VTAIL.n521 VTAIL.n435 0.470328
R954 VTAIL.n173 VTAIL.n87 0.470328
R955 VTAIL.n638 VTAIL.n636 0.388379
R956 VTAIL.n684 VTAIL.n683 0.388379
R957 VTAIL.n687 VTAIL.n614 0.388379
R958 VTAIL.n30 VTAIL.n28 0.388379
R959 VTAIL.n76 VTAIL.n75 0.388379
R960 VTAIL.n79 VTAIL.n6 0.388379
R961 VTAIL.n116 VTAIL.n114 0.388379
R962 VTAIL.n162 VTAIL.n161 0.388379
R963 VTAIL.n165 VTAIL.n92 0.388379
R964 VTAIL.n204 VTAIL.n202 0.388379
R965 VTAIL.n250 VTAIL.n249 0.388379
R966 VTAIL.n253 VTAIL.n180 0.388379
R967 VTAIL.n601 VTAIL.n528 0.388379
R968 VTAIL.n598 VTAIL.n530 0.388379
R969 VTAIL.n554 VTAIL.n552 0.388379
R970 VTAIL.n513 VTAIL.n440 0.388379
R971 VTAIL.n510 VTAIL.n442 0.388379
R972 VTAIL.n466 VTAIL.n464 0.388379
R973 VTAIL.n427 VTAIL.n354 0.388379
R974 VTAIL.n424 VTAIL.n356 0.388379
R975 VTAIL.n380 VTAIL.n378 0.388379
R976 VTAIL.n339 VTAIL.n266 0.388379
R977 VTAIL.n336 VTAIL.n268 0.388379
R978 VTAIL.n292 VTAIL.n290 0.388379
R979 VTAIL.n643 VTAIL.n635 0.155672
R980 VTAIL.n644 VTAIL.n643 0.155672
R981 VTAIL.n644 VTAIL.n631 0.155672
R982 VTAIL.n651 VTAIL.n631 0.155672
R983 VTAIL.n652 VTAIL.n651 0.155672
R984 VTAIL.n652 VTAIL.n627 0.155672
R985 VTAIL.n659 VTAIL.n627 0.155672
R986 VTAIL.n660 VTAIL.n659 0.155672
R987 VTAIL.n660 VTAIL.n623 0.155672
R988 VTAIL.n667 VTAIL.n623 0.155672
R989 VTAIL.n668 VTAIL.n667 0.155672
R990 VTAIL.n668 VTAIL.n619 0.155672
R991 VTAIL.n675 VTAIL.n619 0.155672
R992 VTAIL.n676 VTAIL.n675 0.155672
R993 VTAIL.n676 VTAIL.n615 0.155672
R994 VTAIL.n685 VTAIL.n615 0.155672
R995 VTAIL.n686 VTAIL.n685 0.155672
R996 VTAIL.n686 VTAIL.n611 0.155672
R997 VTAIL.n693 VTAIL.n611 0.155672
R998 VTAIL.n35 VTAIL.n27 0.155672
R999 VTAIL.n36 VTAIL.n35 0.155672
R1000 VTAIL.n36 VTAIL.n23 0.155672
R1001 VTAIL.n43 VTAIL.n23 0.155672
R1002 VTAIL.n44 VTAIL.n43 0.155672
R1003 VTAIL.n44 VTAIL.n19 0.155672
R1004 VTAIL.n51 VTAIL.n19 0.155672
R1005 VTAIL.n52 VTAIL.n51 0.155672
R1006 VTAIL.n52 VTAIL.n15 0.155672
R1007 VTAIL.n59 VTAIL.n15 0.155672
R1008 VTAIL.n60 VTAIL.n59 0.155672
R1009 VTAIL.n60 VTAIL.n11 0.155672
R1010 VTAIL.n67 VTAIL.n11 0.155672
R1011 VTAIL.n68 VTAIL.n67 0.155672
R1012 VTAIL.n68 VTAIL.n7 0.155672
R1013 VTAIL.n77 VTAIL.n7 0.155672
R1014 VTAIL.n78 VTAIL.n77 0.155672
R1015 VTAIL.n78 VTAIL.n3 0.155672
R1016 VTAIL.n85 VTAIL.n3 0.155672
R1017 VTAIL.n121 VTAIL.n113 0.155672
R1018 VTAIL.n122 VTAIL.n121 0.155672
R1019 VTAIL.n122 VTAIL.n109 0.155672
R1020 VTAIL.n129 VTAIL.n109 0.155672
R1021 VTAIL.n130 VTAIL.n129 0.155672
R1022 VTAIL.n130 VTAIL.n105 0.155672
R1023 VTAIL.n137 VTAIL.n105 0.155672
R1024 VTAIL.n138 VTAIL.n137 0.155672
R1025 VTAIL.n138 VTAIL.n101 0.155672
R1026 VTAIL.n145 VTAIL.n101 0.155672
R1027 VTAIL.n146 VTAIL.n145 0.155672
R1028 VTAIL.n146 VTAIL.n97 0.155672
R1029 VTAIL.n153 VTAIL.n97 0.155672
R1030 VTAIL.n154 VTAIL.n153 0.155672
R1031 VTAIL.n154 VTAIL.n93 0.155672
R1032 VTAIL.n163 VTAIL.n93 0.155672
R1033 VTAIL.n164 VTAIL.n163 0.155672
R1034 VTAIL.n164 VTAIL.n89 0.155672
R1035 VTAIL.n171 VTAIL.n89 0.155672
R1036 VTAIL.n209 VTAIL.n201 0.155672
R1037 VTAIL.n210 VTAIL.n209 0.155672
R1038 VTAIL.n210 VTAIL.n197 0.155672
R1039 VTAIL.n217 VTAIL.n197 0.155672
R1040 VTAIL.n218 VTAIL.n217 0.155672
R1041 VTAIL.n218 VTAIL.n193 0.155672
R1042 VTAIL.n225 VTAIL.n193 0.155672
R1043 VTAIL.n226 VTAIL.n225 0.155672
R1044 VTAIL.n226 VTAIL.n189 0.155672
R1045 VTAIL.n233 VTAIL.n189 0.155672
R1046 VTAIL.n234 VTAIL.n233 0.155672
R1047 VTAIL.n234 VTAIL.n185 0.155672
R1048 VTAIL.n241 VTAIL.n185 0.155672
R1049 VTAIL.n242 VTAIL.n241 0.155672
R1050 VTAIL.n242 VTAIL.n181 0.155672
R1051 VTAIL.n251 VTAIL.n181 0.155672
R1052 VTAIL.n252 VTAIL.n251 0.155672
R1053 VTAIL.n252 VTAIL.n177 0.155672
R1054 VTAIL.n259 VTAIL.n177 0.155672
R1055 VTAIL.n607 VTAIL.n525 0.155672
R1056 VTAIL.n600 VTAIL.n525 0.155672
R1057 VTAIL.n600 VTAIL.n599 0.155672
R1058 VTAIL.n599 VTAIL.n529 0.155672
R1059 VTAIL.n592 VTAIL.n529 0.155672
R1060 VTAIL.n592 VTAIL.n591 0.155672
R1061 VTAIL.n591 VTAIL.n535 0.155672
R1062 VTAIL.n584 VTAIL.n535 0.155672
R1063 VTAIL.n584 VTAIL.n583 0.155672
R1064 VTAIL.n583 VTAIL.n539 0.155672
R1065 VTAIL.n576 VTAIL.n539 0.155672
R1066 VTAIL.n576 VTAIL.n575 0.155672
R1067 VTAIL.n575 VTAIL.n543 0.155672
R1068 VTAIL.n568 VTAIL.n543 0.155672
R1069 VTAIL.n568 VTAIL.n567 0.155672
R1070 VTAIL.n567 VTAIL.n547 0.155672
R1071 VTAIL.n560 VTAIL.n547 0.155672
R1072 VTAIL.n560 VTAIL.n559 0.155672
R1073 VTAIL.n559 VTAIL.n551 0.155672
R1074 VTAIL.n519 VTAIL.n437 0.155672
R1075 VTAIL.n512 VTAIL.n437 0.155672
R1076 VTAIL.n512 VTAIL.n511 0.155672
R1077 VTAIL.n511 VTAIL.n441 0.155672
R1078 VTAIL.n504 VTAIL.n441 0.155672
R1079 VTAIL.n504 VTAIL.n503 0.155672
R1080 VTAIL.n503 VTAIL.n447 0.155672
R1081 VTAIL.n496 VTAIL.n447 0.155672
R1082 VTAIL.n496 VTAIL.n495 0.155672
R1083 VTAIL.n495 VTAIL.n451 0.155672
R1084 VTAIL.n488 VTAIL.n451 0.155672
R1085 VTAIL.n488 VTAIL.n487 0.155672
R1086 VTAIL.n487 VTAIL.n455 0.155672
R1087 VTAIL.n480 VTAIL.n455 0.155672
R1088 VTAIL.n480 VTAIL.n479 0.155672
R1089 VTAIL.n479 VTAIL.n459 0.155672
R1090 VTAIL.n472 VTAIL.n459 0.155672
R1091 VTAIL.n472 VTAIL.n471 0.155672
R1092 VTAIL.n471 VTAIL.n463 0.155672
R1093 VTAIL.n433 VTAIL.n351 0.155672
R1094 VTAIL.n426 VTAIL.n351 0.155672
R1095 VTAIL.n426 VTAIL.n425 0.155672
R1096 VTAIL.n425 VTAIL.n355 0.155672
R1097 VTAIL.n418 VTAIL.n355 0.155672
R1098 VTAIL.n418 VTAIL.n417 0.155672
R1099 VTAIL.n417 VTAIL.n361 0.155672
R1100 VTAIL.n410 VTAIL.n361 0.155672
R1101 VTAIL.n410 VTAIL.n409 0.155672
R1102 VTAIL.n409 VTAIL.n365 0.155672
R1103 VTAIL.n402 VTAIL.n365 0.155672
R1104 VTAIL.n402 VTAIL.n401 0.155672
R1105 VTAIL.n401 VTAIL.n369 0.155672
R1106 VTAIL.n394 VTAIL.n369 0.155672
R1107 VTAIL.n394 VTAIL.n393 0.155672
R1108 VTAIL.n393 VTAIL.n373 0.155672
R1109 VTAIL.n386 VTAIL.n373 0.155672
R1110 VTAIL.n386 VTAIL.n385 0.155672
R1111 VTAIL.n385 VTAIL.n377 0.155672
R1112 VTAIL.n345 VTAIL.n263 0.155672
R1113 VTAIL.n338 VTAIL.n263 0.155672
R1114 VTAIL.n338 VTAIL.n337 0.155672
R1115 VTAIL.n337 VTAIL.n267 0.155672
R1116 VTAIL.n330 VTAIL.n267 0.155672
R1117 VTAIL.n330 VTAIL.n329 0.155672
R1118 VTAIL.n329 VTAIL.n273 0.155672
R1119 VTAIL.n322 VTAIL.n273 0.155672
R1120 VTAIL.n322 VTAIL.n321 0.155672
R1121 VTAIL.n321 VTAIL.n277 0.155672
R1122 VTAIL.n314 VTAIL.n277 0.155672
R1123 VTAIL.n314 VTAIL.n313 0.155672
R1124 VTAIL.n313 VTAIL.n281 0.155672
R1125 VTAIL.n306 VTAIL.n281 0.155672
R1126 VTAIL.n306 VTAIL.n305 0.155672
R1127 VTAIL.n305 VTAIL.n285 0.155672
R1128 VTAIL.n298 VTAIL.n285 0.155672
R1129 VTAIL.n298 VTAIL.n297 0.155672
R1130 VTAIL.n297 VTAIL.n289 0.155672
R1131 VTAIL VTAIL.n1 0.0586897
R1132 VDD1 VDD1.n0 63.254
R1133 VDD1.n3 VDD1.n2 63.1403
R1134 VDD1.n3 VDD1.n1 63.1403
R1135 VDD1.n5 VDD1.n4 62.3939
R1136 VDD1.n5 VDD1.n3 44.8242
R1137 VDD1.n4 VDD1.t4 1.28288
R1138 VDD1.n4 VDD1.t7 1.28288
R1139 VDD1.n0 VDD1.t0 1.28288
R1140 VDD1.n0 VDD1.t1 1.28288
R1141 VDD1.n2 VDD1.t6 1.28288
R1142 VDD1.n2 VDD1.t3 1.28288
R1143 VDD1.n1 VDD1.t5 1.28288
R1144 VDD1.n1 VDD1.t2 1.28288
R1145 VDD1 VDD1.n5 0.744035
R1146 B.n859 B.n858 585
R1147 B.n860 B.n859 585
R1148 B.n349 B.n123 585
R1149 B.n348 B.n347 585
R1150 B.n346 B.n345 585
R1151 B.n344 B.n343 585
R1152 B.n342 B.n341 585
R1153 B.n340 B.n339 585
R1154 B.n338 B.n337 585
R1155 B.n336 B.n335 585
R1156 B.n334 B.n333 585
R1157 B.n332 B.n331 585
R1158 B.n330 B.n329 585
R1159 B.n328 B.n327 585
R1160 B.n326 B.n325 585
R1161 B.n324 B.n323 585
R1162 B.n322 B.n321 585
R1163 B.n320 B.n319 585
R1164 B.n318 B.n317 585
R1165 B.n316 B.n315 585
R1166 B.n314 B.n313 585
R1167 B.n312 B.n311 585
R1168 B.n310 B.n309 585
R1169 B.n308 B.n307 585
R1170 B.n306 B.n305 585
R1171 B.n304 B.n303 585
R1172 B.n302 B.n301 585
R1173 B.n300 B.n299 585
R1174 B.n298 B.n297 585
R1175 B.n296 B.n295 585
R1176 B.n294 B.n293 585
R1177 B.n292 B.n291 585
R1178 B.n290 B.n289 585
R1179 B.n288 B.n287 585
R1180 B.n286 B.n285 585
R1181 B.n284 B.n283 585
R1182 B.n282 B.n281 585
R1183 B.n280 B.n279 585
R1184 B.n278 B.n277 585
R1185 B.n276 B.n275 585
R1186 B.n274 B.n273 585
R1187 B.n272 B.n271 585
R1188 B.n270 B.n269 585
R1189 B.n268 B.n267 585
R1190 B.n266 B.n265 585
R1191 B.n264 B.n263 585
R1192 B.n262 B.n261 585
R1193 B.n260 B.n259 585
R1194 B.n258 B.n257 585
R1195 B.n256 B.n255 585
R1196 B.n254 B.n253 585
R1197 B.n252 B.n251 585
R1198 B.n250 B.n249 585
R1199 B.n247 B.n246 585
R1200 B.n245 B.n244 585
R1201 B.n243 B.n242 585
R1202 B.n241 B.n240 585
R1203 B.n239 B.n238 585
R1204 B.n237 B.n236 585
R1205 B.n235 B.n234 585
R1206 B.n233 B.n232 585
R1207 B.n231 B.n230 585
R1208 B.n229 B.n228 585
R1209 B.n227 B.n226 585
R1210 B.n225 B.n224 585
R1211 B.n223 B.n222 585
R1212 B.n221 B.n220 585
R1213 B.n219 B.n218 585
R1214 B.n217 B.n216 585
R1215 B.n215 B.n214 585
R1216 B.n213 B.n212 585
R1217 B.n211 B.n210 585
R1218 B.n209 B.n208 585
R1219 B.n207 B.n206 585
R1220 B.n205 B.n204 585
R1221 B.n203 B.n202 585
R1222 B.n201 B.n200 585
R1223 B.n199 B.n198 585
R1224 B.n197 B.n196 585
R1225 B.n195 B.n194 585
R1226 B.n193 B.n192 585
R1227 B.n191 B.n190 585
R1228 B.n189 B.n188 585
R1229 B.n187 B.n186 585
R1230 B.n185 B.n184 585
R1231 B.n183 B.n182 585
R1232 B.n181 B.n180 585
R1233 B.n179 B.n178 585
R1234 B.n177 B.n176 585
R1235 B.n175 B.n174 585
R1236 B.n173 B.n172 585
R1237 B.n171 B.n170 585
R1238 B.n169 B.n168 585
R1239 B.n167 B.n166 585
R1240 B.n165 B.n164 585
R1241 B.n163 B.n162 585
R1242 B.n161 B.n160 585
R1243 B.n159 B.n158 585
R1244 B.n157 B.n156 585
R1245 B.n155 B.n154 585
R1246 B.n153 B.n152 585
R1247 B.n151 B.n150 585
R1248 B.n149 B.n148 585
R1249 B.n147 B.n146 585
R1250 B.n145 B.n144 585
R1251 B.n143 B.n142 585
R1252 B.n141 B.n140 585
R1253 B.n139 B.n138 585
R1254 B.n137 B.n136 585
R1255 B.n135 B.n134 585
R1256 B.n133 B.n132 585
R1257 B.n131 B.n130 585
R1258 B.n67 B.n66 585
R1259 B.n863 B.n862 585
R1260 B.n857 B.n124 585
R1261 B.n124 B.n64 585
R1262 B.n856 B.n63 585
R1263 B.n867 B.n63 585
R1264 B.n855 B.n62 585
R1265 B.n868 B.n62 585
R1266 B.n854 B.n61 585
R1267 B.n869 B.n61 585
R1268 B.n853 B.n852 585
R1269 B.n852 B.n57 585
R1270 B.n851 B.n56 585
R1271 B.n875 B.n56 585
R1272 B.n850 B.n55 585
R1273 B.n876 B.n55 585
R1274 B.n849 B.n54 585
R1275 B.n877 B.n54 585
R1276 B.n848 B.n847 585
R1277 B.n847 B.n50 585
R1278 B.n846 B.n49 585
R1279 B.n883 B.n49 585
R1280 B.n845 B.n48 585
R1281 B.n884 B.n48 585
R1282 B.n844 B.n47 585
R1283 B.n885 B.n47 585
R1284 B.n843 B.n842 585
R1285 B.n842 B.n43 585
R1286 B.n841 B.n42 585
R1287 B.n891 B.n42 585
R1288 B.n840 B.n41 585
R1289 B.n892 B.n41 585
R1290 B.n839 B.n40 585
R1291 B.n893 B.n40 585
R1292 B.n838 B.n837 585
R1293 B.n837 B.n36 585
R1294 B.n836 B.n35 585
R1295 B.n899 B.n35 585
R1296 B.n835 B.n34 585
R1297 B.n900 B.n34 585
R1298 B.n834 B.n33 585
R1299 B.n901 B.n33 585
R1300 B.n833 B.n832 585
R1301 B.n832 B.n32 585
R1302 B.n831 B.n28 585
R1303 B.n907 B.n28 585
R1304 B.n830 B.n27 585
R1305 B.n908 B.n27 585
R1306 B.n829 B.n26 585
R1307 B.n909 B.n26 585
R1308 B.n828 B.n827 585
R1309 B.n827 B.n22 585
R1310 B.n826 B.n21 585
R1311 B.n915 B.n21 585
R1312 B.n825 B.n20 585
R1313 B.n916 B.n20 585
R1314 B.n824 B.n19 585
R1315 B.n917 B.n19 585
R1316 B.n823 B.n822 585
R1317 B.n822 B.n15 585
R1318 B.n821 B.n14 585
R1319 B.n923 B.n14 585
R1320 B.n820 B.n13 585
R1321 B.n924 B.n13 585
R1322 B.n819 B.n12 585
R1323 B.n925 B.n12 585
R1324 B.n818 B.n817 585
R1325 B.n817 B.n816 585
R1326 B.n815 B.n814 585
R1327 B.n815 B.n8 585
R1328 B.n813 B.n7 585
R1329 B.n932 B.n7 585
R1330 B.n812 B.n6 585
R1331 B.n933 B.n6 585
R1332 B.n811 B.n5 585
R1333 B.n934 B.n5 585
R1334 B.n810 B.n809 585
R1335 B.n809 B.n4 585
R1336 B.n808 B.n350 585
R1337 B.n808 B.n807 585
R1338 B.n798 B.n351 585
R1339 B.n352 B.n351 585
R1340 B.n800 B.n799 585
R1341 B.n801 B.n800 585
R1342 B.n797 B.n357 585
R1343 B.n357 B.n356 585
R1344 B.n796 B.n795 585
R1345 B.n795 B.n794 585
R1346 B.n359 B.n358 585
R1347 B.n360 B.n359 585
R1348 B.n787 B.n786 585
R1349 B.n788 B.n787 585
R1350 B.n785 B.n365 585
R1351 B.n365 B.n364 585
R1352 B.n784 B.n783 585
R1353 B.n783 B.n782 585
R1354 B.n367 B.n366 585
R1355 B.n368 B.n367 585
R1356 B.n775 B.n774 585
R1357 B.n776 B.n775 585
R1358 B.n773 B.n373 585
R1359 B.n373 B.n372 585
R1360 B.n772 B.n771 585
R1361 B.n771 B.n770 585
R1362 B.n375 B.n374 585
R1363 B.n763 B.n375 585
R1364 B.n762 B.n761 585
R1365 B.n764 B.n762 585
R1366 B.n760 B.n380 585
R1367 B.n380 B.n379 585
R1368 B.n759 B.n758 585
R1369 B.n758 B.n757 585
R1370 B.n382 B.n381 585
R1371 B.n383 B.n382 585
R1372 B.n750 B.n749 585
R1373 B.n751 B.n750 585
R1374 B.n748 B.n387 585
R1375 B.n391 B.n387 585
R1376 B.n747 B.n746 585
R1377 B.n746 B.n745 585
R1378 B.n389 B.n388 585
R1379 B.n390 B.n389 585
R1380 B.n738 B.n737 585
R1381 B.n739 B.n738 585
R1382 B.n736 B.n396 585
R1383 B.n396 B.n395 585
R1384 B.n735 B.n734 585
R1385 B.n734 B.n733 585
R1386 B.n398 B.n397 585
R1387 B.n399 B.n398 585
R1388 B.n726 B.n725 585
R1389 B.n727 B.n726 585
R1390 B.n724 B.n403 585
R1391 B.n407 B.n403 585
R1392 B.n723 B.n722 585
R1393 B.n722 B.n721 585
R1394 B.n405 B.n404 585
R1395 B.n406 B.n405 585
R1396 B.n714 B.n713 585
R1397 B.n715 B.n714 585
R1398 B.n712 B.n412 585
R1399 B.n412 B.n411 585
R1400 B.n711 B.n710 585
R1401 B.n710 B.n709 585
R1402 B.n414 B.n413 585
R1403 B.n415 B.n414 585
R1404 B.n705 B.n704 585
R1405 B.n418 B.n417 585
R1406 B.n701 B.n700 585
R1407 B.n702 B.n701 585
R1408 B.n699 B.n474 585
R1409 B.n698 B.n697 585
R1410 B.n696 B.n695 585
R1411 B.n694 B.n693 585
R1412 B.n692 B.n691 585
R1413 B.n690 B.n689 585
R1414 B.n688 B.n687 585
R1415 B.n686 B.n685 585
R1416 B.n684 B.n683 585
R1417 B.n682 B.n681 585
R1418 B.n680 B.n679 585
R1419 B.n678 B.n677 585
R1420 B.n676 B.n675 585
R1421 B.n674 B.n673 585
R1422 B.n672 B.n671 585
R1423 B.n670 B.n669 585
R1424 B.n668 B.n667 585
R1425 B.n666 B.n665 585
R1426 B.n664 B.n663 585
R1427 B.n662 B.n661 585
R1428 B.n660 B.n659 585
R1429 B.n658 B.n657 585
R1430 B.n656 B.n655 585
R1431 B.n654 B.n653 585
R1432 B.n652 B.n651 585
R1433 B.n650 B.n649 585
R1434 B.n648 B.n647 585
R1435 B.n646 B.n645 585
R1436 B.n644 B.n643 585
R1437 B.n642 B.n641 585
R1438 B.n640 B.n639 585
R1439 B.n638 B.n637 585
R1440 B.n636 B.n635 585
R1441 B.n634 B.n633 585
R1442 B.n632 B.n631 585
R1443 B.n630 B.n629 585
R1444 B.n628 B.n627 585
R1445 B.n626 B.n625 585
R1446 B.n624 B.n623 585
R1447 B.n622 B.n621 585
R1448 B.n620 B.n619 585
R1449 B.n618 B.n617 585
R1450 B.n616 B.n615 585
R1451 B.n614 B.n613 585
R1452 B.n612 B.n611 585
R1453 B.n610 B.n609 585
R1454 B.n608 B.n607 585
R1455 B.n606 B.n605 585
R1456 B.n604 B.n603 585
R1457 B.n601 B.n600 585
R1458 B.n599 B.n598 585
R1459 B.n597 B.n596 585
R1460 B.n595 B.n594 585
R1461 B.n593 B.n592 585
R1462 B.n591 B.n590 585
R1463 B.n589 B.n588 585
R1464 B.n587 B.n586 585
R1465 B.n585 B.n584 585
R1466 B.n583 B.n582 585
R1467 B.n581 B.n580 585
R1468 B.n579 B.n578 585
R1469 B.n577 B.n576 585
R1470 B.n575 B.n574 585
R1471 B.n573 B.n572 585
R1472 B.n571 B.n570 585
R1473 B.n569 B.n568 585
R1474 B.n567 B.n566 585
R1475 B.n565 B.n564 585
R1476 B.n563 B.n562 585
R1477 B.n561 B.n560 585
R1478 B.n559 B.n558 585
R1479 B.n557 B.n556 585
R1480 B.n555 B.n554 585
R1481 B.n553 B.n552 585
R1482 B.n551 B.n550 585
R1483 B.n549 B.n548 585
R1484 B.n547 B.n546 585
R1485 B.n545 B.n544 585
R1486 B.n543 B.n542 585
R1487 B.n541 B.n540 585
R1488 B.n539 B.n538 585
R1489 B.n537 B.n536 585
R1490 B.n535 B.n534 585
R1491 B.n533 B.n532 585
R1492 B.n531 B.n530 585
R1493 B.n529 B.n528 585
R1494 B.n527 B.n526 585
R1495 B.n525 B.n524 585
R1496 B.n523 B.n522 585
R1497 B.n521 B.n520 585
R1498 B.n519 B.n518 585
R1499 B.n517 B.n516 585
R1500 B.n515 B.n514 585
R1501 B.n513 B.n512 585
R1502 B.n511 B.n510 585
R1503 B.n509 B.n508 585
R1504 B.n507 B.n506 585
R1505 B.n505 B.n504 585
R1506 B.n503 B.n502 585
R1507 B.n501 B.n500 585
R1508 B.n499 B.n498 585
R1509 B.n497 B.n496 585
R1510 B.n495 B.n494 585
R1511 B.n493 B.n492 585
R1512 B.n491 B.n490 585
R1513 B.n489 B.n488 585
R1514 B.n487 B.n486 585
R1515 B.n485 B.n484 585
R1516 B.n483 B.n482 585
R1517 B.n481 B.n480 585
R1518 B.n706 B.n416 585
R1519 B.n416 B.n415 585
R1520 B.n708 B.n707 585
R1521 B.n709 B.n708 585
R1522 B.n410 B.n409 585
R1523 B.n411 B.n410 585
R1524 B.n717 B.n716 585
R1525 B.n716 B.n715 585
R1526 B.n718 B.n408 585
R1527 B.n408 B.n406 585
R1528 B.n720 B.n719 585
R1529 B.n721 B.n720 585
R1530 B.n402 B.n401 585
R1531 B.n407 B.n402 585
R1532 B.n729 B.n728 585
R1533 B.n728 B.n727 585
R1534 B.n730 B.n400 585
R1535 B.n400 B.n399 585
R1536 B.n732 B.n731 585
R1537 B.n733 B.n732 585
R1538 B.n394 B.n393 585
R1539 B.n395 B.n394 585
R1540 B.n741 B.n740 585
R1541 B.n740 B.n739 585
R1542 B.n742 B.n392 585
R1543 B.n392 B.n390 585
R1544 B.n744 B.n743 585
R1545 B.n745 B.n744 585
R1546 B.n386 B.n385 585
R1547 B.n391 B.n386 585
R1548 B.n753 B.n752 585
R1549 B.n752 B.n751 585
R1550 B.n754 B.n384 585
R1551 B.n384 B.n383 585
R1552 B.n756 B.n755 585
R1553 B.n757 B.n756 585
R1554 B.n378 B.n377 585
R1555 B.n379 B.n378 585
R1556 B.n766 B.n765 585
R1557 B.n765 B.n764 585
R1558 B.n767 B.n376 585
R1559 B.n763 B.n376 585
R1560 B.n769 B.n768 585
R1561 B.n770 B.n769 585
R1562 B.n371 B.n370 585
R1563 B.n372 B.n371 585
R1564 B.n778 B.n777 585
R1565 B.n777 B.n776 585
R1566 B.n779 B.n369 585
R1567 B.n369 B.n368 585
R1568 B.n781 B.n780 585
R1569 B.n782 B.n781 585
R1570 B.n363 B.n362 585
R1571 B.n364 B.n363 585
R1572 B.n790 B.n789 585
R1573 B.n789 B.n788 585
R1574 B.n791 B.n361 585
R1575 B.n361 B.n360 585
R1576 B.n793 B.n792 585
R1577 B.n794 B.n793 585
R1578 B.n355 B.n354 585
R1579 B.n356 B.n355 585
R1580 B.n803 B.n802 585
R1581 B.n802 B.n801 585
R1582 B.n804 B.n353 585
R1583 B.n353 B.n352 585
R1584 B.n806 B.n805 585
R1585 B.n807 B.n806 585
R1586 B.n3 B.n0 585
R1587 B.n4 B.n3 585
R1588 B.n931 B.n1 585
R1589 B.n932 B.n931 585
R1590 B.n930 B.n929 585
R1591 B.n930 B.n8 585
R1592 B.n928 B.n9 585
R1593 B.n816 B.n9 585
R1594 B.n927 B.n926 585
R1595 B.n926 B.n925 585
R1596 B.n11 B.n10 585
R1597 B.n924 B.n11 585
R1598 B.n922 B.n921 585
R1599 B.n923 B.n922 585
R1600 B.n920 B.n16 585
R1601 B.n16 B.n15 585
R1602 B.n919 B.n918 585
R1603 B.n918 B.n917 585
R1604 B.n18 B.n17 585
R1605 B.n916 B.n18 585
R1606 B.n914 B.n913 585
R1607 B.n915 B.n914 585
R1608 B.n912 B.n23 585
R1609 B.n23 B.n22 585
R1610 B.n911 B.n910 585
R1611 B.n910 B.n909 585
R1612 B.n25 B.n24 585
R1613 B.n908 B.n25 585
R1614 B.n906 B.n905 585
R1615 B.n907 B.n906 585
R1616 B.n904 B.n29 585
R1617 B.n32 B.n29 585
R1618 B.n903 B.n902 585
R1619 B.n902 B.n901 585
R1620 B.n31 B.n30 585
R1621 B.n900 B.n31 585
R1622 B.n898 B.n897 585
R1623 B.n899 B.n898 585
R1624 B.n896 B.n37 585
R1625 B.n37 B.n36 585
R1626 B.n895 B.n894 585
R1627 B.n894 B.n893 585
R1628 B.n39 B.n38 585
R1629 B.n892 B.n39 585
R1630 B.n890 B.n889 585
R1631 B.n891 B.n890 585
R1632 B.n888 B.n44 585
R1633 B.n44 B.n43 585
R1634 B.n887 B.n886 585
R1635 B.n886 B.n885 585
R1636 B.n46 B.n45 585
R1637 B.n884 B.n46 585
R1638 B.n882 B.n881 585
R1639 B.n883 B.n882 585
R1640 B.n880 B.n51 585
R1641 B.n51 B.n50 585
R1642 B.n879 B.n878 585
R1643 B.n878 B.n877 585
R1644 B.n53 B.n52 585
R1645 B.n876 B.n53 585
R1646 B.n874 B.n873 585
R1647 B.n875 B.n874 585
R1648 B.n872 B.n58 585
R1649 B.n58 B.n57 585
R1650 B.n871 B.n870 585
R1651 B.n870 B.n869 585
R1652 B.n60 B.n59 585
R1653 B.n868 B.n60 585
R1654 B.n866 B.n865 585
R1655 B.n867 B.n866 585
R1656 B.n864 B.n65 585
R1657 B.n65 B.n64 585
R1658 B.n935 B.n934 585
R1659 B.n933 B.n2 585
R1660 B.n862 B.n65 497.305
R1661 B.n859 B.n124 497.305
R1662 B.n480 B.n414 497.305
R1663 B.n704 B.n416 497.305
R1664 B.n127 B.t19 448.755
R1665 B.n125 B.t8 448.755
R1666 B.n477 B.t12 448.755
R1667 B.n475 B.t16 448.755
R1668 B.n127 B.t20 377.418
R1669 B.n125 B.t10 377.418
R1670 B.n477 B.t15 377.418
R1671 B.n475 B.t18 377.418
R1672 B.n126 B.t11 341.346
R1673 B.n478 B.t14 341.346
R1674 B.n128 B.t21 341.346
R1675 B.n476 B.t17 341.346
R1676 B.n860 B.n122 256.663
R1677 B.n860 B.n121 256.663
R1678 B.n860 B.n120 256.663
R1679 B.n860 B.n119 256.663
R1680 B.n860 B.n118 256.663
R1681 B.n860 B.n117 256.663
R1682 B.n860 B.n116 256.663
R1683 B.n860 B.n115 256.663
R1684 B.n860 B.n114 256.663
R1685 B.n860 B.n113 256.663
R1686 B.n860 B.n112 256.663
R1687 B.n860 B.n111 256.663
R1688 B.n860 B.n110 256.663
R1689 B.n860 B.n109 256.663
R1690 B.n860 B.n108 256.663
R1691 B.n860 B.n107 256.663
R1692 B.n860 B.n106 256.663
R1693 B.n860 B.n105 256.663
R1694 B.n860 B.n104 256.663
R1695 B.n860 B.n103 256.663
R1696 B.n860 B.n102 256.663
R1697 B.n860 B.n101 256.663
R1698 B.n860 B.n100 256.663
R1699 B.n860 B.n99 256.663
R1700 B.n860 B.n98 256.663
R1701 B.n860 B.n97 256.663
R1702 B.n860 B.n96 256.663
R1703 B.n860 B.n95 256.663
R1704 B.n860 B.n94 256.663
R1705 B.n860 B.n93 256.663
R1706 B.n860 B.n92 256.663
R1707 B.n860 B.n91 256.663
R1708 B.n860 B.n90 256.663
R1709 B.n860 B.n89 256.663
R1710 B.n860 B.n88 256.663
R1711 B.n860 B.n87 256.663
R1712 B.n860 B.n86 256.663
R1713 B.n860 B.n85 256.663
R1714 B.n860 B.n84 256.663
R1715 B.n860 B.n83 256.663
R1716 B.n860 B.n82 256.663
R1717 B.n860 B.n81 256.663
R1718 B.n860 B.n80 256.663
R1719 B.n860 B.n79 256.663
R1720 B.n860 B.n78 256.663
R1721 B.n860 B.n77 256.663
R1722 B.n860 B.n76 256.663
R1723 B.n860 B.n75 256.663
R1724 B.n860 B.n74 256.663
R1725 B.n860 B.n73 256.663
R1726 B.n860 B.n72 256.663
R1727 B.n860 B.n71 256.663
R1728 B.n860 B.n70 256.663
R1729 B.n860 B.n69 256.663
R1730 B.n860 B.n68 256.663
R1731 B.n861 B.n860 256.663
R1732 B.n703 B.n702 256.663
R1733 B.n702 B.n419 256.663
R1734 B.n702 B.n420 256.663
R1735 B.n702 B.n421 256.663
R1736 B.n702 B.n422 256.663
R1737 B.n702 B.n423 256.663
R1738 B.n702 B.n424 256.663
R1739 B.n702 B.n425 256.663
R1740 B.n702 B.n426 256.663
R1741 B.n702 B.n427 256.663
R1742 B.n702 B.n428 256.663
R1743 B.n702 B.n429 256.663
R1744 B.n702 B.n430 256.663
R1745 B.n702 B.n431 256.663
R1746 B.n702 B.n432 256.663
R1747 B.n702 B.n433 256.663
R1748 B.n702 B.n434 256.663
R1749 B.n702 B.n435 256.663
R1750 B.n702 B.n436 256.663
R1751 B.n702 B.n437 256.663
R1752 B.n702 B.n438 256.663
R1753 B.n702 B.n439 256.663
R1754 B.n702 B.n440 256.663
R1755 B.n702 B.n441 256.663
R1756 B.n702 B.n442 256.663
R1757 B.n702 B.n443 256.663
R1758 B.n702 B.n444 256.663
R1759 B.n702 B.n445 256.663
R1760 B.n702 B.n446 256.663
R1761 B.n702 B.n447 256.663
R1762 B.n702 B.n448 256.663
R1763 B.n702 B.n449 256.663
R1764 B.n702 B.n450 256.663
R1765 B.n702 B.n451 256.663
R1766 B.n702 B.n452 256.663
R1767 B.n702 B.n453 256.663
R1768 B.n702 B.n454 256.663
R1769 B.n702 B.n455 256.663
R1770 B.n702 B.n456 256.663
R1771 B.n702 B.n457 256.663
R1772 B.n702 B.n458 256.663
R1773 B.n702 B.n459 256.663
R1774 B.n702 B.n460 256.663
R1775 B.n702 B.n461 256.663
R1776 B.n702 B.n462 256.663
R1777 B.n702 B.n463 256.663
R1778 B.n702 B.n464 256.663
R1779 B.n702 B.n465 256.663
R1780 B.n702 B.n466 256.663
R1781 B.n702 B.n467 256.663
R1782 B.n702 B.n468 256.663
R1783 B.n702 B.n469 256.663
R1784 B.n702 B.n470 256.663
R1785 B.n702 B.n471 256.663
R1786 B.n702 B.n472 256.663
R1787 B.n702 B.n473 256.663
R1788 B.n937 B.n936 256.663
R1789 B.n130 B.n67 163.367
R1790 B.n134 B.n133 163.367
R1791 B.n138 B.n137 163.367
R1792 B.n142 B.n141 163.367
R1793 B.n146 B.n145 163.367
R1794 B.n150 B.n149 163.367
R1795 B.n154 B.n153 163.367
R1796 B.n158 B.n157 163.367
R1797 B.n162 B.n161 163.367
R1798 B.n166 B.n165 163.367
R1799 B.n170 B.n169 163.367
R1800 B.n174 B.n173 163.367
R1801 B.n178 B.n177 163.367
R1802 B.n182 B.n181 163.367
R1803 B.n186 B.n185 163.367
R1804 B.n190 B.n189 163.367
R1805 B.n194 B.n193 163.367
R1806 B.n198 B.n197 163.367
R1807 B.n202 B.n201 163.367
R1808 B.n206 B.n205 163.367
R1809 B.n210 B.n209 163.367
R1810 B.n214 B.n213 163.367
R1811 B.n218 B.n217 163.367
R1812 B.n222 B.n221 163.367
R1813 B.n226 B.n225 163.367
R1814 B.n230 B.n229 163.367
R1815 B.n234 B.n233 163.367
R1816 B.n238 B.n237 163.367
R1817 B.n242 B.n241 163.367
R1818 B.n246 B.n245 163.367
R1819 B.n251 B.n250 163.367
R1820 B.n255 B.n254 163.367
R1821 B.n259 B.n258 163.367
R1822 B.n263 B.n262 163.367
R1823 B.n267 B.n266 163.367
R1824 B.n271 B.n270 163.367
R1825 B.n275 B.n274 163.367
R1826 B.n279 B.n278 163.367
R1827 B.n283 B.n282 163.367
R1828 B.n287 B.n286 163.367
R1829 B.n291 B.n290 163.367
R1830 B.n295 B.n294 163.367
R1831 B.n299 B.n298 163.367
R1832 B.n303 B.n302 163.367
R1833 B.n307 B.n306 163.367
R1834 B.n311 B.n310 163.367
R1835 B.n315 B.n314 163.367
R1836 B.n319 B.n318 163.367
R1837 B.n323 B.n322 163.367
R1838 B.n327 B.n326 163.367
R1839 B.n331 B.n330 163.367
R1840 B.n335 B.n334 163.367
R1841 B.n339 B.n338 163.367
R1842 B.n343 B.n342 163.367
R1843 B.n347 B.n346 163.367
R1844 B.n859 B.n123 163.367
R1845 B.n710 B.n414 163.367
R1846 B.n710 B.n412 163.367
R1847 B.n714 B.n412 163.367
R1848 B.n714 B.n405 163.367
R1849 B.n722 B.n405 163.367
R1850 B.n722 B.n403 163.367
R1851 B.n726 B.n403 163.367
R1852 B.n726 B.n398 163.367
R1853 B.n734 B.n398 163.367
R1854 B.n734 B.n396 163.367
R1855 B.n738 B.n396 163.367
R1856 B.n738 B.n389 163.367
R1857 B.n746 B.n389 163.367
R1858 B.n746 B.n387 163.367
R1859 B.n750 B.n387 163.367
R1860 B.n750 B.n382 163.367
R1861 B.n758 B.n382 163.367
R1862 B.n758 B.n380 163.367
R1863 B.n762 B.n380 163.367
R1864 B.n762 B.n375 163.367
R1865 B.n771 B.n375 163.367
R1866 B.n771 B.n373 163.367
R1867 B.n775 B.n373 163.367
R1868 B.n775 B.n367 163.367
R1869 B.n783 B.n367 163.367
R1870 B.n783 B.n365 163.367
R1871 B.n787 B.n365 163.367
R1872 B.n787 B.n359 163.367
R1873 B.n795 B.n359 163.367
R1874 B.n795 B.n357 163.367
R1875 B.n800 B.n357 163.367
R1876 B.n800 B.n351 163.367
R1877 B.n808 B.n351 163.367
R1878 B.n809 B.n808 163.367
R1879 B.n809 B.n5 163.367
R1880 B.n6 B.n5 163.367
R1881 B.n7 B.n6 163.367
R1882 B.n815 B.n7 163.367
R1883 B.n817 B.n815 163.367
R1884 B.n817 B.n12 163.367
R1885 B.n13 B.n12 163.367
R1886 B.n14 B.n13 163.367
R1887 B.n822 B.n14 163.367
R1888 B.n822 B.n19 163.367
R1889 B.n20 B.n19 163.367
R1890 B.n21 B.n20 163.367
R1891 B.n827 B.n21 163.367
R1892 B.n827 B.n26 163.367
R1893 B.n27 B.n26 163.367
R1894 B.n28 B.n27 163.367
R1895 B.n832 B.n28 163.367
R1896 B.n832 B.n33 163.367
R1897 B.n34 B.n33 163.367
R1898 B.n35 B.n34 163.367
R1899 B.n837 B.n35 163.367
R1900 B.n837 B.n40 163.367
R1901 B.n41 B.n40 163.367
R1902 B.n42 B.n41 163.367
R1903 B.n842 B.n42 163.367
R1904 B.n842 B.n47 163.367
R1905 B.n48 B.n47 163.367
R1906 B.n49 B.n48 163.367
R1907 B.n847 B.n49 163.367
R1908 B.n847 B.n54 163.367
R1909 B.n55 B.n54 163.367
R1910 B.n56 B.n55 163.367
R1911 B.n852 B.n56 163.367
R1912 B.n852 B.n61 163.367
R1913 B.n62 B.n61 163.367
R1914 B.n63 B.n62 163.367
R1915 B.n124 B.n63 163.367
R1916 B.n701 B.n418 163.367
R1917 B.n701 B.n474 163.367
R1918 B.n697 B.n696 163.367
R1919 B.n693 B.n692 163.367
R1920 B.n689 B.n688 163.367
R1921 B.n685 B.n684 163.367
R1922 B.n681 B.n680 163.367
R1923 B.n677 B.n676 163.367
R1924 B.n673 B.n672 163.367
R1925 B.n669 B.n668 163.367
R1926 B.n665 B.n664 163.367
R1927 B.n661 B.n660 163.367
R1928 B.n657 B.n656 163.367
R1929 B.n653 B.n652 163.367
R1930 B.n649 B.n648 163.367
R1931 B.n645 B.n644 163.367
R1932 B.n641 B.n640 163.367
R1933 B.n637 B.n636 163.367
R1934 B.n633 B.n632 163.367
R1935 B.n629 B.n628 163.367
R1936 B.n625 B.n624 163.367
R1937 B.n621 B.n620 163.367
R1938 B.n617 B.n616 163.367
R1939 B.n613 B.n612 163.367
R1940 B.n609 B.n608 163.367
R1941 B.n605 B.n604 163.367
R1942 B.n600 B.n599 163.367
R1943 B.n596 B.n595 163.367
R1944 B.n592 B.n591 163.367
R1945 B.n588 B.n587 163.367
R1946 B.n584 B.n583 163.367
R1947 B.n580 B.n579 163.367
R1948 B.n576 B.n575 163.367
R1949 B.n572 B.n571 163.367
R1950 B.n568 B.n567 163.367
R1951 B.n564 B.n563 163.367
R1952 B.n560 B.n559 163.367
R1953 B.n556 B.n555 163.367
R1954 B.n552 B.n551 163.367
R1955 B.n548 B.n547 163.367
R1956 B.n544 B.n543 163.367
R1957 B.n540 B.n539 163.367
R1958 B.n536 B.n535 163.367
R1959 B.n532 B.n531 163.367
R1960 B.n528 B.n527 163.367
R1961 B.n524 B.n523 163.367
R1962 B.n520 B.n519 163.367
R1963 B.n516 B.n515 163.367
R1964 B.n512 B.n511 163.367
R1965 B.n508 B.n507 163.367
R1966 B.n504 B.n503 163.367
R1967 B.n500 B.n499 163.367
R1968 B.n496 B.n495 163.367
R1969 B.n492 B.n491 163.367
R1970 B.n488 B.n487 163.367
R1971 B.n484 B.n483 163.367
R1972 B.n708 B.n416 163.367
R1973 B.n708 B.n410 163.367
R1974 B.n716 B.n410 163.367
R1975 B.n716 B.n408 163.367
R1976 B.n720 B.n408 163.367
R1977 B.n720 B.n402 163.367
R1978 B.n728 B.n402 163.367
R1979 B.n728 B.n400 163.367
R1980 B.n732 B.n400 163.367
R1981 B.n732 B.n394 163.367
R1982 B.n740 B.n394 163.367
R1983 B.n740 B.n392 163.367
R1984 B.n744 B.n392 163.367
R1985 B.n744 B.n386 163.367
R1986 B.n752 B.n386 163.367
R1987 B.n752 B.n384 163.367
R1988 B.n756 B.n384 163.367
R1989 B.n756 B.n378 163.367
R1990 B.n765 B.n378 163.367
R1991 B.n765 B.n376 163.367
R1992 B.n769 B.n376 163.367
R1993 B.n769 B.n371 163.367
R1994 B.n777 B.n371 163.367
R1995 B.n777 B.n369 163.367
R1996 B.n781 B.n369 163.367
R1997 B.n781 B.n363 163.367
R1998 B.n789 B.n363 163.367
R1999 B.n789 B.n361 163.367
R2000 B.n793 B.n361 163.367
R2001 B.n793 B.n355 163.367
R2002 B.n802 B.n355 163.367
R2003 B.n802 B.n353 163.367
R2004 B.n806 B.n353 163.367
R2005 B.n806 B.n3 163.367
R2006 B.n935 B.n3 163.367
R2007 B.n931 B.n2 163.367
R2008 B.n931 B.n930 163.367
R2009 B.n930 B.n9 163.367
R2010 B.n926 B.n9 163.367
R2011 B.n926 B.n11 163.367
R2012 B.n922 B.n11 163.367
R2013 B.n922 B.n16 163.367
R2014 B.n918 B.n16 163.367
R2015 B.n918 B.n18 163.367
R2016 B.n914 B.n18 163.367
R2017 B.n914 B.n23 163.367
R2018 B.n910 B.n23 163.367
R2019 B.n910 B.n25 163.367
R2020 B.n906 B.n25 163.367
R2021 B.n906 B.n29 163.367
R2022 B.n902 B.n29 163.367
R2023 B.n902 B.n31 163.367
R2024 B.n898 B.n31 163.367
R2025 B.n898 B.n37 163.367
R2026 B.n894 B.n37 163.367
R2027 B.n894 B.n39 163.367
R2028 B.n890 B.n39 163.367
R2029 B.n890 B.n44 163.367
R2030 B.n886 B.n44 163.367
R2031 B.n886 B.n46 163.367
R2032 B.n882 B.n46 163.367
R2033 B.n882 B.n51 163.367
R2034 B.n878 B.n51 163.367
R2035 B.n878 B.n53 163.367
R2036 B.n874 B.n53 163.367
R2037 B.n874 B.n58 163.367
R2038 B.n870 B.n58 163.367
R2039 B.n870 B.n60 163.367
R2040 B.n866 B.n60 163.367
R2041 B.n866 B.n65 163.367
R2042 B.n862 B.n861 71.676
R2043 B.n130 B.n68 71.676
R2044 B.n134 B.n69 71.676
R2045 B.n138 B.n70 71.676
R2046 B.n142 B.n71 71.676
R2047 B.n146 B.n72 71.676
R2048 B.n150 B.n73 71.676
R2049 B.n154 B.n74 71.676
R2050 B.n158 B.n75 71.676
R2051 B.n162 B.n76 71.676
R2052 B.n166 B.n77 71.676
R2053 B.n170 B.n78 71.676
R2054 B.n174 B.n79 71.676
R2055 B.n178 B.n80 71.676
R2056 B.n182 B.n81 71.676
R2057 B.n186 B.n82 71.676
R2058 B.n190 B.n83 71.676
R2059 B.n194 B.n84 71.676
R2060 B.n198 B.n85 71.676
R2061 B.n202 B.n86 71.676
R2062 B.n206 B.n87 71.676
R2063 B.n210 B.n88 71.676
R2064 B.n214 B.n89 71.676
R2065 B.n218 B.n90 71.676
R2066 B.n222 B.n91 71.676
R2067 B.n226 B.n92 71.676
R2068 B.n230 B.n93 71.676
R2069 B.n234 B.n94 71.676
R2070 B.n238 B.n95 71.676
R2071 B.n242 B.n96 71.676
R2072 B.n246 B.n97 71.676
R2073 B.n251 B.n98 71.676
R2074 B.n255 B.n99 71.676
R2075 B.n259 B.n100 71.676
R2076 B.n263 B.n101 71.676
R2077 B.n267 B.n102 71.676
R2078 B.n271 B.n103 71.676
R2079 B.n275 B.n104 71.676
R2080 B.n279 B.n105 71.676
R2081 B.n283 B.n106 71.676
R2082 B.n287 B.n107 71.676
R2083 B.n291 B.n108 71.676
R2084 B.n295 B.n109 71.676
R2085 B.n299 B.n110 71.676
R2086 B.n303 B.n111 71.676
R2087 B.n307 B.n112 71.676
R2088 B.n311 B.n113 71.676
R2089 B.n315 B.n114 71.676
R2090 B.n319 B.n115 71.676
R2091 B.n323 B.n116 71.676
R2092 B.n327 B.n117 71.676
R2093 B.n331 B.n118 71.676
R2094 B.n335 B.n119 71.676
R2095 B.n339 B.n120 71.676
R2096 B.n343 B.n121 71.676
R2097 B.n347 B.n122 71.676
R2098 B.n123 B.n122 71.676
R2099 B.n346 B.n121 71.676
R2100 B.n342 B.n120 71.676
R2101 B.n338 B.n119 71.676
R2102 B.n334 B.n118 71.676
R2103 B.n330 B.n117 71.676
R2104 B.n326 B.n116 71.676
R2105 B.n322 B.n115 71.676
R2106 B.n318 B.n114 71.676
R2107 B.n314 B.n113 71.676
R2108 B.n310 B.n112 71.676
R2109 B.n306 B.n111 71.676
R2110 B.n302 B.n110 71.676
R2111 B.n298 B.n109 71.676
R2112 B.n294 B.n108 71.676
R2113 B.n290 B.n107 71.676
R2114 B.n286 B.n106 71.676
R2115 B.n282 B.n105 71.676
R2116 B.n278 B.n104 71.676
R2117 B.n274 B.n103 71.676
R2118 B.n270 B.n102 71.676
R2119 B.n266 B.n101 71.676
R2120 B.n262 B.n100 71.676
R2121 B.n258 B.n99 71.676
R2122 B.n254 B.n98 71.676
R2123 B.n250 B.n97 71.676
R2124 B.n245 B.n96 71.676
R2125 B.n241 B.n95 71.676
R2126 B.n237 B.n94 71.676
R2127 B.n233 B.n93 71.676
R2128 B.n229 B.n92 71.676
R2129 B.n225 B.n91 71.676
R2130 B.n221 B.n90 71.676
R2131 B.n217 B.n89 71.676
R2132 B.n213 B.n88 71.676
R2133 B.n209 B.n87 71.676
R2134 B.n205 B.n86 71.676
R2135 B.n201 B.n85 71.676
R2136 B.n197 B.n84 71.676
R2137 B.n193 B.n83 71.676
R2138 B.n189 B.n82 71.676
R2139 B.n185 B.n81 71.676
R2140 B.n181 B.n80 71.676
R2141 B.n177 B.n79 71.676
R2142 B.n173 B.n78 71.676
R2143 B.n169 B.n77 71.676
R2144 B.n165 B.n76 71.676
R2145 B.n161 B.n75 71.676
R2146 B.n157 B.n74 71.676
R2147 B.n153 B.n73 71.676
R2148 B.n149 B.n72 71.676
R2149 B.n145 B.n71 71.676
R2150 B.n141 B.n70 71.676
R2151 B.n137 B.n69 71.676
R2152 B.n133 B.n68 71.676
R2153 B.n861 B.n67 71.676
R2154 B.n704 B.n703 71.676
R2155 B.n474 B.n419 71.676
R2156 B.n696 B.n420 71.676
R2157 B.n692 B.n421 71.676
R2158 B.n688 B.n422 71.676
R2159 B.n684 B.n423 71.676
R2160 B.n680 B.n424 71.676
R2161 B.n676 B.n425 71.676
R2162 B.n672 B.n426 71.676
R2163 B.n668 B.n427 71.676
R2164 B.n664 B.n428 71.676
R2165 B.n660 B.n429 71.676
R2166 B.n656 B.n430 71.676
R2167 B.n652 B.n431 71.676
R2168 B.n648 B.n432 71.676
R2169 B.n644 B.n433 71.676
R2170 B.n640 B.n434 71.676
R2171 B.n636 B.n435 71.676
R2172 B.n632 B.n436 71.676
R2173 B.n628 B.n437 71.676
R2174 B.n624 B.n438 71.676
R2175 B.n620 B.n439 71.676
R2176 B.n616 B.n440 71.676
R2177 B.n612 B.n441 71.676
R2178 B.n608 B.n442 71.676
R2179 B.n604 B.n443 71.676
R2180 B.n599 B.n444 71.676
R2181 B.n595 B.n445 71.676
R2182 B.n591 B.n446 71.676
R2183 B.n587 B.n447 71.676
R2184 B.n583 B.n448 71.676
R2185 B.n579 B.n449 71.676
R2186 B.n575 B.n450 71.676
R2187 B.n571 B.n451 71.676
R2188 B.n567 B.n452 71.676
R2189 B.n563 B.n453 71.676
R2190 B.n559 B.n454 71.676
R2191 B.n555 B.n455 71.676
R2192 B.n551 B.n456 71.676
R2193 B.n547 B.n457 71.676
R2194 B.n543 B.n458 71.676
R2195 B.n539 B.n459 71.676
R2196 B.n535 B.n460 71.676
R2197 B.n531 B.n461 71.676
R2198 B.n527 B.n462 71.676
R2199 B.n523 B.n463 71.676
R2200 B.n519 B.n464 71.676
R2201 B.n515 B.n465 71.676
R2202 B.n511 B.n466 71.676
R2203 B.n507 B.n467 71.676
R2204 B.n503 B.n468 71.676
R2205 B.n499 B.n469 71.676
R2206 B.n495 B.n470 71.676
R2207 B.n491 B.n471 71.676
R2208 B.n487 B.n472 71.676
R2209 B.n483 B.n473 71.676
R2210 B.n703 B.n418 71.676
R2211 B.n697 B.n419 71.676
R2212 B.n693 B.n420 71.676
R2213 B.n689 B.n421 71.676
R2214 B.n685 B.n422 71.676
R2215 B.n681 B.n423 71.676
R2216 B.n677 B.n424 71.676
R2217 B.n673 B.n425 71.676
R2218 B.n669 B.n426 71.676
R2219 B.n665 B.n427 71.676
R2220 B.n661 B.n428 71.676
R2221 B.n657 B.n429 71.676
R2222 B.n653 B.n430 71.676
R2223 B.n649 B.n431 71.676
R2224 B.n645 B.n432 71.676
R2225 B.n641 B.n433 71.676
R2226 B.n637 B.n434 71.676
R2227 B.n633 B.n435 71.676
R2228 B.n629 B.n436 71.676
R2229 B.n625 B.n437 71.676
R2230 B.n621 B.n438 71.676
R2231 B.n617 B.n439 71.676
R2232 B.n613 B.n440 71.676
R2233 B.n609 B.n441 71.676
R2234 B.n605 B.n442 71.676
R2235 B.n600 B.n443 71.676
R2236 B.n596 B.n444 71.676
R2237 B.n592 B.n445 71.676
R2238 B.n588 B.n446 71.676
R2239 B.n584 B.n447 71.676
R2240 B.n580 B.n448 71.676
R2241 B.n576 B.n449 71.676
R2242 B.n572 B.n450 71.676
R2243 B.n568 B.n451 71.676
R2244 B.n564 B.n452 71.676
R2245 B.n560 B.n453 71.676
R2246 B.n556 B.n454 71.676
R2247 B.n552 B.n455 71.676
R2248 B.n548 B.n456 71.676
R2249 B.n544 B.n457 71.676
R2250 B.n540 B.n458 71.676
R2251 B.n536 B.n459 71.676
R2252 B.n532 B.n460 71.676
R2253 B.n528 B.n461 71.676
R2254 B.n524 B.n462 71.676
R2255 B.n520 B.n463 71.676
R2256 B.n516 B.n464 71.676
R2257 B.n512 B.n465 71.676
R2258 B.n508 B.n466 71.676
R2259 B.n504 B.n467 71.676
R2260 B.n500 B.n468 71.676
R2261 B.n496 B.n469 71.676
R2262 B.n492 B.n470 71.676
R2263 B.n488 B.n471 71.676
R2264 B.n484 B.n472 71.676
R2265 B.n480 B.n473 71.676
R2266 B.n936 B.n935 71.676
R2267 B.n936 B.n2 71.676
R2268 B.n702 B.n415 64.2535
R2269 B.n860 B.n64 64.2535
R2270 B.n129 B.n128 59.5399
R2271 B.n248 B.n126 59.5399
R2272 B.n479 B.n478 59.5399
R2273 B.n602 B.n476 59.5399
R2274 B.n709 B.n415 36.1096
R2275 B.n709 B.n411 36.1096
R2276 B.n715 B.n411 36.1096
R2277 B.n715 B.n406 36.1096
R2278 B.n721 B.n406 36.1096
R2279 B.n721 B.n407 36.1096
R2280 B.n727 B.n399 36.1096
R2281 B.n733 B.n399 36.1096
R2282 B.n733 B.n395 36.1096
R2283 B.n739 B.n395 36.1096
R2284 B.n739 B.n390 36.1096
R2285 B.n745 B.n390 36.1096
R2286 B.n745 B.n391 36.1096
R2287 B.n751 B.n383 36.1096
R2288 B.n757 B.n383 36.1096
R2289 B.n757 B.n379 36.1096
R2290 B.n764 B.n379 36.1096
R2291 B.n764 B.n763 36.1096
R2292 B.n770 B.n372 36.1096
R2293 B.n776 B.n372 36.1096
R2294 B.n776 B.n368 36.1096
R2295 B.n782 B.n368 36.1096
R2296 B.n788 B.n364 36.1096
R2297 B.n788 B.n360 36.1096
R2298 B.n794 B.n360 36.1096
R2299 B.n794 B.n356 36.1096
R2300 B.n801 B.n356 36.1096
R2301 B.n807 B.n352 36.1096
R2302 B.n807 B.n4 36.1096
R2303 B.n934 B.n4 36.1096
R2304 B.n934 B.n933 36.1096
R2305 B.n933 B.n932 36.1096
R2306 B.n932 B.n8 36.1096
R2307 B.n816 B.n8 36.1096
R2308 B.n925 B.n924 36.1096
R2309 B.n924 B.n923 36.1096
R2310 B.n923 B.n15 36.1096
R2311 B.n917 B.n15 36.1096
R2312 B.n917 B.n916 36.1096
R2313 B.n915 B.n22 36.1096
R2314 B.n909 B.n22 36.1096
R2315 B.n909 B.n908 36.1096
R2316 B.n908 B.n907 36.1096
R2317 B.n901 B.n32 36.1096
R2318 B.n901 B.n900 36.1096
R2319 B.n900 B.n899 36.1096
R2320 B.n899 B.n36 36.1096
R2321 B.n893 B.n36 36.1096
R2322 B.n892 B.n891 36.1096
R2323 B.n891 B.n43 36.1096
R2324 B.n885 B.n43 36.1096
R2325 B.n885 B.n884 36.1096
R2326 B.n884 B.n883 36.1096
R2327 B.n883 B.n50 36.1096
R2328 B.n877 B.n50 36.1096
R2329 B.n876 B.n875 36.1096
R2330 B.n875 B.n57 36.1096
R2331 B.n869 B.n57 36.1096
R2332 B.n869 B.n868 36.1096
R2333 B.n868 B.n867 36.1096
R2334 B.n867 B.n64 36.1096
R2335 B.n128 B.n127 36.0732
R2336 B.n126 B.n125 36.0732
R2337 B.n478 B.n477 36.0732
R2338 B.n476 B.n475 36.0732
R2339 B.n727 B.t13 33.4545
R2340 B.n877 B.t9 33.4545
R2341 B.n706 B.n705 32.3127
R2342 B.n481 B.n413 32.3127
R2343 B.n858 B.n857 32.3127
R2344 B.n864 B.n863 32.3127
R2345 B.t2 B.n352 30.2684
R2346 B.n816 B.t0 30.2684
R2347 B.n770 B.t6 28.1444
R2348 B.n907 B.t4 28.1444
R2349 B.n391 B.t7 27.0823
R2350 B.t5 B.n892 27.0823
R2351 B.n782 B.t1 24.9583
R2352 B.t3 B.n915 24.9583
R2353 B B.n937 18.0485
R2354 B.t1 B.n364 11.1518
R2355 B.n916 B.t3 11.1518
R2356 B.n707 B.n706 10.6151
R2357 B.n707 B.n409 10.6151
R2358 B.n717 B.n409 10.6151
R2359 B.n718 B.n717 10.6151
R2360 B.n719 B.n718 10.6151
R2361 B.n719 B.n401 10.6151
R2362 B.n729 B.n401 10.6151
R2363 B.n730 B.n729 10.6151
R2364 B.n731 B.n730 10.6151
R2365 B.n731 B.n393 10.6151
R2366 B.n741 B.n393 10.6151
R2367 B.n742 B.n741 10.6151
R2368 B.n743 B.n742 10.6151
R2369 B.n743 B.n385 10.6151
R2370 B.n753 B.n385 10.6151
R2371 B.n754 B.n753 10.6151
R2372 B.n755 B.n754 10.6151
R2373 B.n755 B.n377 10.6151
R2374 B.n766 B.n377 10.6151
R2375 B.n767 B.n766 10.6151
R2376 B.n768 B.n767 10.6151
R2377 B.n768 B.n370 10.6151
R2378 B.n778 B.n370 10.6151
R2379 B.n779 B.n778 10.6151
R2380 B.n780 B.n779 10.6151
R2381 B.n780 B.n362 10.6151
R2382 B.n790 B.n362 10.6151
R2383 B.n791 B.n790 10.6151
R2384 B.n792 B.n791 10.6151
R2385 B.n792 B.n354 10.6151
R2386 B.n803 B.n354 10.6151
R2387 B.n804 B.n803 10.6151
R2388 B.n805 B.n804 10.6151
R2389 B.n805 B.n0 10.6151
R2390 B.n705 B.n417 10.6151
R2391 B.n700 B.n417 10.6151
R2392 B.n700 B.n699 10.6151
R2393 B.n699 B.n698 10.6151
R2394 B.n698 B.n695 10.6151
R2395 B.n695 B.n694 10.6151
R2396 B.n694 B.n691 10.6151
R2397 B.n691 B.n690 10.6151
R2398 B.n690 B.n687 10.6151
R2399 B.n687 B.n686 10.6151
R2400 B.n686 B.n683 10.6151
R2401 B.n683 B.n682 10.6151
R2402 B.n682 B.n679 10.6151
R2403 B.n679 B.n678 10.6151
R2404 B.n678 B.n675 10.6151
R2405 B.n675 B.n674 10.6151
R2406 B.n674 B.n671 10.6151
R2407 B.n671 B.n670 10.6151
R2408 B.n670 B.n667 10.6151
R2409 B.n667 B.n666 10.6151
R2410 B.n666 B.n663 10.6151
R2411 B.n663 B.n662 10.6151
R2412 B.n662 B.n659 10.6151
R2413 B.n659 B.n658 10.6151
R2414 B.n658 B.n655 10.6151
R2415 B.n655 B.n654 10.6151
R2416 B.n654 B.n651 10.6151
R2417 B.n651 B.n650 10.6151
R2418 B.n650 B.n647 10.6151
R2419 B.n647 B.n646 10.6151
R2420 B.n646 B.n643 10.6151
R2421 B.n643 B.n642 10.6151
R2422 B.n642 B.n639 10.6151
R2423 B.n639 B.n638 10.6151
R2424 B.n638 B.n635 10.6151
R2425 B.n635 B.n634 10.6151
R2426 B.n634 B.n631 10.6151
R2427 B.n631 B.n630 10.6151
R2428 B.n630 B.n627 10.6151
R2429 B.n627 B.n626 10.6151
R2430 B.n626 B.n623 10.6151
R2431 B.n623 B.n622 10.6151
R2432 B.n622 B.n619 10.6151
R2433 B.n619 B.n618 10.6151
R2434 B.n618 B.n615 10.6151
R2435 B.n615 B.n614 10.6151
R2436 B.n614 B.n611 10.6151
R2437 B.n611 B.n610 10.6151
R2438 B.n610 B.n607 10.6151
R2439 B.n607 B.n606 10.6151
R2440 B.n606 B.n603 10.6151
R2441 B.n601 B.n598 10.6151
R2442 B.n598 B.n597 10.6151
R2443 B.n597 B.n594 10.6151
R2444 B.n594 B.n593 10.6151
R2445 B.n593 B.n590 10.6151
R2446 B.n590 B.n589 10.6151
R2447 B.n589 B.n586 10.6151
R2448 B.n586 B.n585 10.6151
R2449 B.n582 B.n581 10.6151
R2450 B.n581 B.n578 10.6151
R2451 B.n578 B.n577 10.6151
R2452 B.n577 B.n574 10.6151
R2453 B.n574 B.n573 10.6151
R2454 B.n573 B.n570 10.6151
R2455 B.n570 B.n569 10.6151
R2456 B.n569 B.n566 10.6151
R2457 B.n566 B.n565 10.6151
R2458 B.n565 B.n562 10.6151
R2459 B.n562 B.n561 10.6151
R2460 B.n561 B.n558 10.6151
R2461 B.n558 B.n557 10.6151
R2462 B.n557 B.n554 10.6151
R2463 B.n554 B.n553 10.6151
R2464 B.n553 B.n550 10.6151
R2465 B.n550 B.n549 10.6151
R2466 B.n549 B.n546 10.6151
R2467 B.n546 B.n545 10.6151
R2468 B.n545 B.n542 10.6151
R2469 B.n542 B.n541 10.6151
R2470 B.n541 B.n538 10.6151
R2471 B.n538 B.n537 10.6151
R2472 B.n537 B.n534 10.6151
R2473 B.n534 B.n533 10.6151
R2474 B.n533 B.n530 10.6151
R2475 B.n530 B.n529 10.6151
R2476 B.n529 B.n526 10.6151
R2477 B.n526 B.n525 10.6151
R2478 B.n525 B.n522 10.6151
R2479 B.n522 B.n521 10.6151
R2480 B.n521 B.n518 10.6151
R2481 B.n518 B.n517 10.6151
R2482 B.n517 B.n514 10.6151
R2483 B.n514 B.n513 10.6151
R2484 B.n513 B.n510 10.6151
R2485 B.n510 B.n509 10.6151
R2486 B.n509 B.n506 10.6151
R2487 B.n506 B.n505 10.6151
R2488 B.n505 B.n502 10.6151
R2489 B.n502 B.n501 10.6151
R2490 B.n501 B.n498 10.6151
R2491 B.n498 B.n497 10.6151
R2492 B.n497 B.n494 10.6151
R2493 B.n494 B.n493 10.6151
R2494 B.n493 B.n490 10.6151
R2495 B.n490 B.n489 10.6151
R2496 B.n489 B.n486 10.6151
R2497 B.n486 B.n485 10.6151
R2498 B.n485 B.n482 10.6151
R2499 B.n482 B.n481 10.6151
R2500 B.n711 B.n413 10.6151
R2501 B.n712 B.n711 10.6151
R2502 B.n713 B.n712 10.6151
R2503 B.n713 B.n404 10.6151
R2504 B.n723 B.n404 10.6151
R2505 B.n724 B.n723 10.6151
R2506 B.n725 B.n724 10.6151
R2507 B.n725 B.n397 10.6151
R2508 B.n735 B.n397 10.6151
R2509 B.n736 B.n735 10.6151
R2510 B.n737 B.n736 10.6151
R2511 B.n737 B.n388 10.6151
R2512 B.n747 B.n388 10.6151
R2513 B.n748 B.n747 10.6151
R2514 B.n749 B.n748 10.6151
R2515 B.n749 B.n381 10.6151
R2516 B.n759 B.n381 10.6151
R2517 B.n760 B.n759 10.6151
R2518 B.n761 B.n760 10.6151
R2519 B.n761 B.n374 10.6151
R2520 B.n772 B.n374 10.6151
R2521 B.n773 B.n772 10.6151
R2522 B.n774 B.n773 10.6151
R2523 B.n774 B.n366 10.6151
R2524 B.n784 B.n366 10.6151
R2525 B.n785 B.n784 10.6151
R2526 B.n786 B.n785 10.6151
R2527 B.n786 B.n358 10.6151
R2528 B.n796 B.n358 10.6151
R2529 B.n797 B.n796 10.6151
R2530 B.n799 B.n797 10.6151
R2531 B.n799 B.n798 10.6151
R2532 B.n798 B.n350 10.6151
R2533 B.n810 B.n350 10.6151
R2534 B.n811 B.n810 10.6151
R2535 B.n812 B.n811 10.6151
R2536 B.n813 B.n812 10.6151
R2537 B.n814 B.n813 10.6151
R2538 B.n818 B.n814 10.6151
R2539 B.n819 B.n818 10.6151
R2540 B.n820 B.n819 10.6151
R2541 B.n821 B.n820 10.6151
R2542 B.n823 B.n821 10.6151
R2543 B.n824 B.n823 10.6151
R2544 B.n825 B.n824 10.6151
R2545 B.n826 B.n825 10.6151
R2546 B.n828 B.n826 10.6151
R2547 B.n829 B.n828 10.6151
R2548 B.n830 B.n829 10.6151
R2549 B.n831 B.n830 10.6151
R2550 B.n833 B.n831 10.6151
R2551 B.n834 B.n833 10.6151
R2552 B.n835 B.n834 10.6151
R2553 B.n836 B.n835 10.6151
R2554 B.n838 B.n836 10.6151
R2555 B.n839 B.n838 10.6151
R2556 B.n840 B.n839 10.6151
R2557 B.n841 B.n840 10.6151
R2558 B.n843 B.n841 10.6151
R2559 B.n844 B.n843 10.6151
R2560 B.n845 B.n844 10.6151
R2561 B.n846 B.n845 10.6151
R2562 B.n848 B.n846 10.6151
R2563 B.n849 B.n848 10.6151
R2564 B.n850 B.n849 10.6151
R2565 B.n851 B.n850 10.6151
R2566 B.n853 B.n851 10.6151
R2567 B.n854 B.n853 10.6151
R2568 B.n855 B.n854 10.6151
R2569 B.n856 B.n855 10.6151
R2570 B.n857 B.n856 10.6151
R2571 B.n929 B.n1 10.6151
R2572 B.n929 B.n928 10.6151
R2573 B.n928 B.n927 10.6151
R2574 B.n927 B.n10 10.6151
R2575 B.n921 B.n10 10.6151
R2576 B.n921 B.n920 10.6151
R2577 B.n920 B.n919 10.6151
R2578 B.n919 B.n17 10.6151
R2579 B.n913 B.n17 10.6151
R2580 B.n913 B.n912 10.6151
R2581 B.n912 B.n911 10.6151
R2582 B.n911 B.n24 10.6151
R2583 B.n905 B.n24 10.6151
R2584 B.n905 B.n904 10.6151
R2585 B.n904 B.n903 10.6151
R2586 B.n903 B.n30 10.6151
R2587 B.n897 B.n30 10.6151
R2588 B.n897 B.n896 10.6151
R2589 B.n896 B.n895 10.6151
R2590 B.n895 B.n38 10.6151
R2591 B.n889 B.n38 10.6151
R2592 B.n889 B.n888 10.6151
R2593 B.n888 B.n887 10.6151
R2594 B.n887 B.n45 10.6151
R2595 B.n881 B.n45 10.6151
R2596 B.n881 B.n880 10.6151
R2597 B.n880 B.n879 10.6151
R2598 B.n879 B.n52 10.6151
R2599 B.n873 B.n52 10.6151
R2600 B.n873 B.n872 10.6151
R2601 B.n872 B.n871 10.6151
R2602 B.n871 B.n59 10.6151
R2603 B.n865 B.n59 10.6151
R2604 B.n865 B.n864 10.6151
R2605 B.n863 B.n66 10.6151
R2606 B.n131 B.n66 10.6151
R2607 B.n132 B.n131 10.6151
R2608 B.n135 B.n132 10.6151
R2609 B.n136 B.n135 10.6151
R2610 B.n139 B.n136 10.6151
R2611 B.n140 B.n139 10.6151
R2612 B.n143 B.n140 10.6151
R2613 B.n144 B.n143 10.6151
R2614 B.n147 B.n144 10.6151
R2615 B.n148 B.n147 10.6151
R2616 B.n151 B.n148 10.6151
R2617 B.n152 B.n151 10.6151
R2618 B.n155 B.n152 10.6151
R2619 B.n156 B.n155 10.6151
R2620 B.n159 B.n156 10.6151
R2621 B.n160 B.n159 10.6151
R2622 B.n163 B.n160 10.6151
R2623 B.n164 B.n163 10.6151
R2624 B.n167 B.n164 10.6151
R2625 B.n168 B.n167 10.6151
R2626 B.n171 B.n168 10.6151
R2627 B.n172 B.n171 10.6151
R2628 B.n175 B.n172 10.6151
R2629 B.n176 B.n175 10.6151
R2630 B.n179 B.n176 10.6151
R2631 B.n180 B.n179 10.6151
R2632 B.n183 B.n180 10.6151
R2633 B.n184 B.n183 10.6151
R2634 B.n187 B.n184 10.6151
R2635 B.n188 B.n187 10.6151
R2636 B.n191 B.n188 10.6151
R2637 B.n192 B.n191 10.6151
R2638 B.n195 B.n192 10.6151
R2639 B.n196 B.n195 10.6151
R2640 B.n199 B.n196 10.6151
R2641 B.n200 B.n199 10.6151
R2642 B.n203 B.n200 10.6151
R2643 B.n204 B.n203 10.6151
R2644 B.n207 B.n204 10.6151
R2645 B.n208 B.n207 10.6151
R2646 B.n211 B.n208 10.6151
R2647 B.n212 B.n211 10.6151
R2648 B.n215 B.n212 10.6151
R2649 B.n216 B.n215 10.6151
R2650 B.n219 B.n216 10.6151
R2651 B.n220 B.n219 10.6151
R2652 B.n223 B.n220 10.6151
R2653 B.n224 B.n223 10.6151
R2654 B.n227 B.n224 10.6151
R2655 B.n228 B.n227 10.6151
R2656 B.n232 B.n231 10.6151
R2657 B.n235 B.n232 10.6151
R2658 B.n236 B.n235 10.6151
R2659 B.n239 B.n236 10.6151
R2660 B.n240 B.n239 10.6151
R2661 B.n243 B.n240 10.6151
R2662 B.n244 B.n243 10.6151
R2663 B.n247 B.n244 10.6151
R2664 B.n252 B.n249 10.6151
R2665 B.n253 B.n252 10.6151
R2666 B.n256 B.n253 10.6151
R2667 B.n257 B.n256 10.6151
R2668 B.n260 B.n257 10.6151
R2669 B.n261 B.n260 10.6151
R2670 B.n264 B.n261 10.6151
R2671 B.n265 B.n264 10.6151
R2672 B.n268 B.n265 10.6151
R2673 B.n269 B.n268 10.6151
R2674 B.n272 B.n269 10.6151
R2675 B.n273 B.n272 10.6151
R2676 B.n276 B.n273 10.6151
R2677 B.n277 B.n276 10.6151
R2678 B.n280 B.n277 10.6151
R2679 B.n281 B.n280 10.6151
R2680 B.n284 B.n281 10.6151
R2681 B.n285 B.n284 10.6151
R2682 B.n288 B.n285 10.6151
R2683 B.n289 B.n288 10.6151
R2684 B.n292 B.n289 10.6151
R2685 B.n293 B.n292 10.6151
R2686 B.n296 B.n293 10.6151
R2687 B.n297 B.n296 10.6151
R2688 B.n300 B.n297 10.6151
R2689 B.n301 B.n300 10.6151
R2690 B.n304 B.n301 10.6151
R2691 B.n305 B.n304 10.6151
R2692 B.n308 B.n305 10.6151
R2693 B.n309 B.n308 10.6151
R2694 B.n312 B.n309 10.6151
R2695 B.n313 B.n312 10.6151
R2696 B.n316 B.n313 10.6151
R2697 B.n317 B.n316 10.6151
R2698 B.n320 B.n317 10.6151
R2699 B.n321 B.n320 10.6151
R2700 B.n324 B.n321 10.6151
R2701 B.n325 B.n324 10.6151
R2702 B.n328 B.n325 10.6151
R2703 B.n329 B.n328 10.6151
R2704 B.n332 B.n329 10.6151
R2705 B.n333 B.n332 10.6151
R2706 B.n336 B.n333 10.6151
R2707 B.n337 B.n336 10.6151
R2708 B.n340 B.n337 10.6151
R2709 B.n341 B.n340 10.6151
R2710 B.n344 B.n341 10.6151
R2711 B.n345 B.n344 10.6151
R2712 B.n348 B.n345 10.6151
R2713 B.n349 B.n348 10.6151
R2714 B.n858 B.n349 10.6151
R2715 B.n751 B.t7 9.02778
R2716 B.n893 B.t5 9.02778
R2717 B.n937 B.n0 8.11757
R2718 B.n937 B.n1 8.11757
R2719 B.n763 B.t6 7.96574
R2720 B.n32 B.t4 7.96574
R2721 B.n602 B.n601 6.5566
R2722 B.n585 B.n479 6.5566
R2723 B.n231 B.n129 6.5566
R2724 B.n248 B.n247 6.5566
R2725 B.n801 B.t2 5.84168
R2726 B.n925 B.t0 5.84168
R2727 B.n603 B.n602 4.05904
R2728 B.n582 B.n479 4.05904
R2729 B.n228 B.n129 4.05904
R2730 B.n249 B.n248 4.05904
R2731 B.n407 B.t13 2.65558
R2732 B.t9 B.n876 2.65558
R2733 VN.n5 VN.t6 279.474
R2734 VN.n24 VN.t7 279.474
R2735 VN.n4 VN.t3 243.206
R2736 VN.n10 VN.t4 243.206
R2737 VN.n17 VN.t2 243.206
R2738 VN.n23 VN.t5 243.206
R2739 VN.n29 VN.t0 243.206
R2740 VN.n36 VN.t1 243.206
R2741 VN.n18 VN.n17 171.63
R2742 VN.n37 VN.n36 171.63
R2743 VN.n35 VN.n19 161.3
R2744 VN.n34 VN.n33 161.3
R2745 VN.n32 VN.n20 161.3
R2746 VN.n31 VN.n30 161.3
R2747 VN.n28 VN.n21 161.3
R2748 VN.n27 VN.n26 161.3
R2749 VN.n25 VN.n22 161.3
R2750 VN.n16 VN.n0 161.3
R2751 VN.n15 VN.n14 161.3
R2752 VN.n13 VN.n1 161.3
R2753 VN.n12 VN.n11 161.3
R2754 VN.n9 VN.n2 161.3
R2755 VN.n8 VN.n7 161.3
R2756 VN.n6 VN.n3 161.3
R2757 VN.n15 VN.n1 54.1398
R2758 VN.n34 VN.n20 54.1398
R2759 VN VN.n37 48.8736
R2760 VN.n5 VN.n4 45.6659
R2761 VN.n24 VN.n23 45.6659
R2762 VN.n8 VN.n3 40.577
R2763 VN.n9 VN.n8 40.577
R2764 VN.n27 VN.n22 40.577
R2765 VN.n28 VN.n27 40.577
R2766 VN.n16 VN.n15 27.0143
R2767 VN.n35 VN.n34 27.0143
R2768 VN.n11 VN.n1 24.5923
R2769 VN.n30 VN.n20 24.5923
R2770 VN.n4 VN.n3 21.1495
R2771 VN.n10 VN.n9 21.1495
R2772 VN.n23 VN.n22 21.1495
R2773 VN.n29 VN.n28 21.1495
R2774 VN.n25 VN.n24 17.3242
R2775 VN.n6 VN.n5 17.3242
R2776 VN.n17 VN.n16 14.2638
R2777 VN.n36 VN.n35 14.2638
R2778 VN.n11 VN.n10 3.44336
R2779 VN.n30 VN.n29 3.44336
R2780 VN.n37 VN.n19 0.189894
R2781 VN.n33 VN.n19 0.189894
R2782 VN.n33 VN.n32 0.189894
R2783 VN.n32 VN.n31 0.189894
R2784 VN.n31 VN.n21 0.189894
R2785 VN.n26 VN.n21 0.189894
R2786 VN.n26 VN.n25 0.189894
R2787 VN.n7 VN.n6 0.189894
R2788 VN.n7 VN.n2 0.189894
R2789 VN.n12 VN.n2 0.189894
R2790 VN.n13 VN.n12 0.189894
R2791 VN.n14 VN.n13 0.189894
R2792 VN.n14 VN.n0 0.189894
R2793 VN.n18 VN.n0 0.189894
R2794 VN VN.n18 0.0516364
R2795 VDD2.n2 VDD2.n1 63.1403
R2796 VDD2.n2 VDD2.n0 63.1403
R2797 VDD2 VDD2.n5 63.1375
R2798 VDD2.n4 VDD2.n3 62.3941
R2799 VDD2.n4 VDD2.n2 44.2412
R2800 VDD2.n5 VDD2.t2 1.28288
R2801 VDD2.n5 VDD2.t0 1.28288
R2802 VDD2.n3 VDD2.t6 1.28288
R2803 VDD2.n3 VDD2.t7 1.28288
R2804 VDD2.n1 VDD2.t3 1.28288
R2805 VDD2.n1 VDD2.t5 1.28288
R2806 VDD2.n0 VDD2.t1 1.28288
R2807 VDD2.n0 VDD2.t4 1.28288
R2808 VDD2 VDD2.n4 0.860414
C0 VN VDD2 9.672231f
C1 VN VP 6.983069f
C2 VTAIL VDD2 10.0549f
C3 VDD1 VDD2 1.23559f
C4 VTAIL VP 9.60435f
C5 VP VDD1 9.927401f
C6 VP VDD2 0.406108f
C7 VN VTAIL 9.59024f
C8 VN VDD1 0.15009f
C9 VTAIL VDD1 10.0077f
C10 VDD2 B 4.56867f
C11 VDD1 B 4.887232f
C12 VTAIL B 11.671393f
C13 VN B 11.8143f
C14 VP B 10.10477f
C15 VDD2.t1 B 0.305997f
C16 VDD2.t4 B 0.305997f
C17 VDD2.n0 B 2.77606f
C18 VDD2.t3 B 0.305997f
C19 VDD2.t5 B 0.305997f
C20 VDD2.n1 B 2.77606f
C21 VDD2.n2 B 2.87529f
C22 VDD2.t6 B 0.305997f
C23 VDD2.t7 B 0.305997f
C24 VDD2.n3 B 2.77129f
C25 VDD2.n4 B 2.84856f
C26 VDD2.t2 B 0.305997f
C27 VDD2.t0 B 0.305997f
C28 VDD2.n5 B 2.77603f
C29 VN.n0 B 0.030115f
C30 VN.t2 B 1.95069f
C31 VN.n1 B 0.052536f
C32 VN.n2 B 0.030115f
C33 VN.t4 B 1.95069f
C34 VN.n3 B 0.055679f
C35 VN.t6 B 2.05618f
C36 VN.t3 B 1.95069f
C37 VN.n4 B 0.7591f
C38 VN.n5 B 0.756122f
C39 VN.n6 B 0.193036f
C40 VN.n7 B 0.030115f
C41 VN.n8 B 0.024323f
C42 VN.n9 B 0.055679f
C43 VN.n10 B 0.692146f
C44 VN.n11 B 0.032136f
C45 VN.n12 B 0.030115f
C46 VN.n13 B 0.030115f
C47 VN.n14 B 0.030115f
C48 VN.n15 B 0.032794f
C49 VN.n16 B 0.046491f
C50 VN.n17 B 0.761214f
C51 VN.n18 B 0.027761f
C52 VN.n19 B 0.030115f
C53 VN.t1 B 1.95069f
C54 VN.n20 B 0.052536f
C55 VN.n21 B 0.030115f
C56 VN.t0 B 1.95069f
C57 VN.n22 B 0.055679f
C58 VN.t7 B 2.05618f
C59 VN.t5 B 1.95069f
C60 VN.n23 B 0.7591f
C61 VN.n24 B 0.756122f
C62 VN.n25 B 0.193036f
C63 VN.n26 B 0.030115f
C64 VN.n27 B 0.024323f
C65 VN.n28 B 0.055679f
C66 VN.n29 B 0.692146f
C67 VN.n30 B 0.032136f
C68 VN.n31 B 0.030115f
C69 VN.n32 B 0.030115f
C70 VN.n33 B 0.030115f
C71 VN.n34 B 0.032794f
C72 VN.n35 B 0.046491f
C73 VN.n36 B 0.761214f
C74 VN.n37 B 1.58706f
C75 VDD1.t0 B 0.30611f
C76 VDD1.t1 B 0.30611f
C77 VDD1.n0 B 2.77793f
C78 VDD1.t5 B 0.30611f
C79 VDD1.t2 B 0.30611f
C80 VDD1.n1 B 2.77709f
C81 VDD1.t6 B 0.30611f
C82 VDD1.t3 B 0.30611f
C83 VDD1.n2 B 2.77709f
C84 VDD1.n3 B 2.92911f
C85 VDD1.t4 B 0.30611f
C86 VDD1.t7 B 0.30611f
C87 VDD1.n4 B 2.7723f
C88 VDD1.n5 B 2.88013f
C89 VTAIL.t3 B 0.227635f
C90 VTAIL.t4 B 0.227635f
C91 VTAIL.n0 B 2.00747f
C92 VTAIL.n1 B 0.280512f
C93 VTAIL.n2 B 0.025217f
C94 VTAIL.n3 B 0.018657f
C95 VTAIL.n4 B 0.010025f
C96 VTAIL.n5 B 0.023696f
C97 VTAIL.n6 B 0.01032f
C98 VTAIL.n7 B 0.018657f
C99 VTAIL.n8 B 0.010615f
C100 VTAIL.n9 B 0.023696f
C101 VTAIL.n10 B 0.010615f
C102 VTAIL.n11 B 0.018657f
C103 VTAIL.n12 B 0.010025f
C104 VTAIL.n13 B 0.023696f
C105 VTAIL.n14 B 0.010615f
C106 VTAIL.n15 B 0.018657f
C107 VTAIL.n16 B 0.010025f
C108 VTAIL.n17 B 0.023696f
C109 VTAIL.n18 B 0.010615f
C110 VTAIL.n19 B 0.018657f
C111 VTAIL.n20 B 0.010025f
C112 VTAIL.n21 B 0.023696f
C113 VTAIL.n22 B 0.010615f
C114 VTAIL.n23 B 0.018657f
C115 VTAIL.n24 B 0.010025f
C116 VTAIL.n25 B 0.023696f
C117 VTAIL.n26 B 0.010615f
C118 VTAIL.n27 B 1.25146f
C119 VTAIL.n28 B 0.010025f
C120 VTAIL.t0 B 0.0391f
C121 VTAIL.n29 B 0.123742f
C122 VTAIL.n30 B 0.013998f
C123 VTAIL.n31 B 0.017772f
C124 VTAIL.n32 B 0.023696f
C125 VTAIL.n33 B 0.010615f
C126 VTAIL.n34 B 0.010025f
C127 VTAIL.n35 B 0.018657f
C128 VTAIL.n36 B 0.018657f
C129 VTAIL.n37 B 0.010025f
C130 VTAIL.n38 B 0.010615f
C131 VTAIL.n39 B 0.023696f
C132 VTAIL.n40 B 0.023696f
C133 VTAIL.n41 B 0.010615f
C134 VTAIL.n42 B 0.010025f
C135 VTAIL.n43 B 0.018657f
C136 VTAIL.n44 B 0.018657f
C137 VTAIL.n45 B 0.010025f
C138 VTAIL.n46 B 0.010615f
C139 VTAIL.n47 B 0.023696f
C140 VTAIL.n48 B 0.023696f
C141 VTAIL.n49 B 0.010615f
C142 VTAIL.n50 B 0.010025f
C143 VTAIL.n51 B 0.018657f
C144 VTAIL.n52 B 0.018657f
C145 VTAIL.n53 B 0.010025f
C146 VTAIL.n54 B 0.010615f
C147 VTAIL.n55 B 0.023696f
C148 VTAIL.n56 B 0.023696f
C149 VTAIL.n57 B 0.010615f
C150 VTAIL.n58 B 0.010025f
C151 VTAIL.n59 B 0.018657f
C152 VTAIL.n60 B 0.018657f
C153 VTAIL.n61 B 0.010025f
C154 VTAIL.n62 B 0.010615f
C155 VTAIL.n63 B 0.023696f
C156 VTAIL.n64 B 0.023696f
C157 VTAIL.n65 B 0.010615f
C158 VTAIL.n66 B 0.010025f
C159 VTAIL.n67 B 0.018657f
C160 VTAIL.n68 B 0.018657f
C161 VTAIL.n69 B 0.010025f
C162 VTAIL.n70 B 0.010025f
C163 VTAIL.n71 B 0.010615f
C164 VTAIL.n72 B 0.023696f
C165 VTAIL.n73 B 0.023696f
C166 VTAIL.n74 B 0.023696f
C167 VTAIL.n75 B 0.01032f
C168 VTAIL.n76 B 0.010025f
C169 VTAIL.n77 B 0.018657f
C170 VTAIL.n78 B 0.018657f
C171 VTAIL.n79 B 0.010025f
C172 VTAIL.n80 B 0.010615f
C173 VTAIL.n81 B 0.023696f
C174 VTAIL.n82 B 0.049518f
C175 VTAIL.n83 B 0.010615f
C176 VTAIL.n84 B 0.010025f
C177 VTAIL.n85 B 0.045163f
C178 VTAIL.n86 B 0.027585f
C179 VTAIL.n87 B 0.141724f
C180 VTAIL.n88 B 0.025217f
C181 VTAIL.n89 B 0.018657f
C182 VTAIL.n90 B 0.010025f
C183 VTAIL.n91 B 0.023696f
C184 VTAIL.n92 B 0.01032f
C185 VTAIL.n93 B 0.018657f
C186 VTAIL.n94 B 0.010615f
C187 VTAIL.n95 B 0.023696f
C188 VTAIL.n96 B 0.010615f
C189 VTAIL.n97 B 0.018657f
C190 VTAIL.n98 B 0.010025f
C191 VTAIL.n99 B 0.023696f
C192 VTAIL.n100 B 0.010615f
C193 VTAIL.n101 B 0.018657f
C194 VTAIL.n102 B 0.010025f
C195 VTAIL.n103 B 0.023696f
C196 VTAIL.n104 B 0.010615f
C197 VTAIL.n105 B 0.018657f
C198 VTAIL.n106 B 0.010025f
C199 VTAIL.n107 B 0.023696f
C200 VTAIL.n108 B 0.010615f
C201 VTAIL.n109 B 0.018657f
C202 VTAIL.n110 B 0.010025f
C203 VTAIL.n111 B 0.023696f
C204 VTAIL.n112 B 0.010615f
C205 VTAIL.n113 B 1.25146f
C206 VTAIL.n114 B 0.010025f
C207 VTAIL.t9 B 0.0391f
C208 VTAIL.n115 B 0.123742f
C209 VTAIL.n116 B 0.013998f
C210 VTAIL.n117 B 0.017772f
C211 VTAIL.n118 B 0.023696f
C212 VTAIL.n119 B 0.010615f
C213 VTAIL.n120 B 0.010025f
C214 VTAIL.n121 B 0.018657f
C215 VTAIL.n122 B 0.018657f
C216 VTAIL.n123 B 0.010025f
C217 VTAIL.n124 B 0.010615f
C218 VTAIL.n125 B 0.023696f
C219 VTAIL.n126 B 0.023696f
C220 VTAIL.n127 B 0.010615f
C221 VTAIL.n128 B 0.010025f
C222 VTAIL.n129 B 0.018657f
C223 VTAIL.n130 B 0.018657f
C224 VTAIL.n131 B 0.010025f
C225 VTAIL.n132 B 0.010615f
C226 VTAIL.n133 B 0.023696f
C227 VTAIL.n134 B 0.023696f
C228 VTAIL.n135 B 0.010615f
C229 VTAIL.n136 B 0.010025f
C230 VTAIL.n137 B 0.018657f
C231 VTAIL.n138 B 0.018657f
C232 VTAIL.n139 B 0.010025f
C233 VTAIL.n140 B 0.010615f
C234 VTAIL.n141 B 0.023696f
C235 VTAIL.n142 B 0.023696f
C236 VTAIL.n143 B 0.010615f
C237 VTAIL.n144 B 0.010025f
C238 VTAIL.n145 B 0.018657f
C239 VTAIL.n146 B 0.018657f
C240 VTAIL.n147 B 0.010025f
C241 VTAIL.n148 B 0.010615f
C242 VTAIL.n149 B 0.023696f
C243 VTAIL.n150 B 0.023696f
C244 VTAIL.n151 B 0.010615f
C245 VTAIL.n152 B 0.010025f
C246 VTAIL.n153 B 0.018657f
C247 VTAIL.n154 B 0.018657f
C248 VTAIL.n155 B 0.010025f
C249 VTAIL.n156 B 0.010025f
C250 VTAIL.n157 B 0.010615f
C251 VTAIL.n158 B 0.023696f
C252 VTAIL.n159 B 0.023696f
C253 VTAIL.n160 B 0.023696f
C254 VTAIL.n161 B 0.01032f
C255 VTAIL.n162 B 0.010025f
C256 VTAIL.n163 B 0.018657f
C257 VTAIL.n164 B 0.018657f
C258 VTAIL.n165 B 0.010025f
C259 VTAIL.n166 B 0.010615f
C260 VTAIL.n167 B 0.023696f
C261 VTAIL.n168 B 0.049518f
C262 VTAIL.n169 B 0.010615f
C263 VTAIL.n170 B 0.010025f
C264 VTAIL.n171 B 0.045163f
C265 VTAIL.n172 B 0.027585f
C266 VTAIL.n173 B 0.141724f
C267 VTAIL.t10 B 0.227635f
C268 VTAIL.t15 B 0.227635f
C269 VTAIL.n174 B 2.00747f
C270 VTAIL.n175 B 0.373407f
C271 VTAIL.n176 B 0.025217f
C272 VTAIL.n177 B 0.018657f
C273 VTAIL.n178 B 0.010025f
C274 VTAIL.n179 B 0.023696f
C275 VTAIL.n180 B 0.01032f
C276 VTAIL.n181 B 0.018657f
C277 VTAIL.n182 B 0.010615f
C278 VTAIL.n183 B 0.023696f
C279 VTAIL.n184 B 0.010615f
C280 VTAIL.n185 B 0.018657f
C281 VTAIL.n186 B 0.010025f
C282 VTAIL.n187 B 0.023696f
C283 VTAIL.n188 B 0.010615f
C284 VTAIL.n189 B 0.018657f
C285 VTAIL.n190 B 0.010025f
C286 VTAIL.n191 B 0.023696f
C287 VTAIL.n192 B 0.010615f
C288 VTAIL.n193 B 0.018657f
C289 VTAIL.n194 B 0.010025f
C290 VTAIL.n195 B 0.023696f
C291 VTAIL.n196 B 0.010615f
C292 VTAIL.n197 B 0.018657f
C293 VTAIL.n198 B 0.010025f
C294 VTAIL.n199 B 0.023696f
C295 VTAIL.n200 B 0.010615f
C296 VTAIL.n201 B 1.25146f
C297 VTAIL.n202 B 0.010025f
C298 VTAIL.t14 B 0.0391f
C299 VTAIL.n203 B 0.123742f
C300 VTAIL.n204 B 0.013998f
C301 VTAIL.n205 B 0.017772f
C302 VTAIL.n206 B 0.023696f
C303 VTAIL.n207 B 0.010615f
C304 VTAIL.n208 B 0.010025f
C305 VTAIL.n209 B 0.018657f
C306 VTAIL.n210 B 0.018657f
C307 VTAIL.n211 B 0.010025f
C308 VTAIL.n212 B 0.010615f
C309 VTAIL.n213 B 0.023696f
C310 VTAIL.n214 B 0.023696f
C311 VTAIL.n215 B 0.010615f
C312 VTAIL.n216 B 0.010025f
C313 VTAIL.n217 B 0.018657f
C314 VTAIL.n218 B 0.018657f
C315 VTAIL.n219 B 0.010025f
C316 VTAIL.n220 B 0.010615f
C317 VTAIL.n221 B 0.023696f
C318 VTAIL.n222 B 0.023696f
C319 VTAIL.n223 B 0.010615f
C320 VTAIL.n224 B 0.010025f
C321 VTAIL.n225 B 0.018657f
C322 VTAIL.n226 B 0.018657f
C323 VTAIL.n227 B 0.010025f
C324 VTAIL.n228 B 0.010615f
C325 VTAIL.n229 B 0.023696f
C326 VTAIL.n230 B 0.023696f
C327 VTAIL.n231 B 0.010615f
C328 VTAIL.n232 B 0.010025f
C329 VTAIL.n233 B 0.018657f
C330 VTAIL.n234 B 0.018657f
C331 VTAIL.n235 B 0.010025f
C332 VTAIL.n236 B 0.010615f
C333 VTAIL.n237 B 0.023696f
C334 VTAIL.n238 B 0.023696f
C335 VTAIL.n239 B 0.010615f
C336 VTAIL.n240 B 0.010025f
C337 VTAIL.n241 B 0.018657f
C338 VTAIL.n242 B 0.018657f
C339 VTAIL.n243 B 0.010025f
C340 VTAIL.n244 B 0.010025f
C341 VTAIL.n245 B 0.010615f
C342 VTAIL.n246 B 0.023696f
C343 VTAIL.n247 B 0.023696f
C344 VTAIL.n248 B 0.023696f
C345 VTAIL.n249 B 0.01032f
C346 VTAIL.n250 B 0.010025f
C347 VTAIL.n251 B 0.018657f
C348 VTAIL.n252 B 0.018657f
C349 VTAIL.n253 B 0.010025f
C350 VTAIL.n254 B 0.010615f
C351 VTAIL.n255 B 0.023696f
C352 VTAIL.n256 B 0.049518f
C353 VTAIL.n257 B 0.010615f
C354 VTAIL.n258 B 0.010025f
C355 VTAIL.n259 B 0.045163f
C356 VTAIL.n260 B 0.027585f
C357 VTAIL.n261 B 1.26347f
C358 VTAIL.n262 B 0.025217f
C359 VTAIL.n263 B 0.018657f
C360 VTAIL.n264 B 0.010025f
C361 VTAIL.n265 B 0.023696f
C362 VTAIL.n266 B 0.01032f
C363 VTAIL.n267 B 0.018657f
C364 VTAIL.n268 B 0.01032f
C365 VTAIL.n269 B 0.010025f
C366 VTAIL.n270 B 0.023696f
C367 VTAIL.n271 B 0.023696f
C368 VTAIL.n272 B 0.010615f
C369 VTAIL.n273 B 0.018657f
C370 VTAIL.n274 B 0.010025f
C371 VTAIL.n275 B 0.023696f
C372 VTAIL.n276 B 0.010615f
C373 VTAIL.n277 B 0.018657f
C374 VTAIL.n278 B 0.010025f
C375 VTAIL.n279 B 0.023696f
C376 VTAIL.n280 B 0.010615f
C377 VTAIL.n281 B 0.018657f
C378 VTAIL.n282 B 0.010025f
C379 VTAIL.n283 B 0.023696f
C380 VTAIL.n284 B 0.010615f
C381 VTAIL.n285 B 0.018657f
C382 VTAIL.n286 B 0.010025f
C383 VTAIL.n287 B 0.023696f
C384 VTAIL.n288 B 0.010615f
C385 VTAIL.n289 B 1.25146f
C386 VTAIL.n290 B 0.010025f
C387 VTAIL.t7 B 0.0391f
C388 VTAIL.n291 B 0.123742f
C389 VTAIL.n292 B 0.013998f
C390 VTAIL.n293 B 0.017772f
C391 VTAIL.n294 B 0.023696f
C392 VTAIL.n295 B 0.010615f
C393 VTAIL.n296 B 0.010025f
C394 VTAIL.n297 B 0.018657f
C395 VTAIL.n298 B 0.018657f
C396 VTAIL.n299 B 0.010025f
C397 VTAIL.n300 B 0.010615f
C398 VTAIL.n301 B 0.023696f
C399 VTAIL.n302 B 0.023696f
C400 VTAIL.n303 B 0.010615f
C401 VTAIL.n304 B 0.010025f
C402 VTAIL.n305 B 0.018657f
C403 VTAIL.n306 B 0.018657f
C404 VTAIL.n307 B 0.010025f
C405 VTAIL.n308 B 0.010615f
C406 VTAIL.n309 B 0.023696f
C407 VTAIL.n310 B 0.023696f
C408 VTAIL.n311 B 0.010615f
C409 VTAIL.n312 B 0.010025f
C410 VTAIL.n313 B 0.018657f
C411 VTAIL.n314 B 0.018657f
C412 VTAIL.n315 B 0.010025f
C413 VTAIL.n316 B 0.010615f
C414 VTAIL.n317 B 0.023696f
C415 VTAIL.n318 B 0.023696f
C416 VTAIL.n319 B 0.010615f
C417 VTAIL.n320 B 0.010025f
C418 VTAIL.n321 B 0.018657f
C419 VTAIL.n322 B 0.018657f
C420 VTAIL.n323 B 0.010025f
C421 VTAIL.n324 B 0.010615f
C422 VTAIL.n325 B 0.023696f
C423 VTAIL.n326 B 0.023696f
C424 VTAIL.n327 B 0.010615f
C425 VTAIL.n328 B 0.010025f
C426 VTAIL.n329 B 0.018657f
C427 VTAIL.n330 B 0.018657f
C428 VTAIL.n331 B 0.010025f
C429 VTAIL.n332 B 0.010615f
C430 VTAIL.n333 B 0.023696f
C431 VTAIL.n334 B 0.023696f
C432 VTAIL.n335 B 0.010615f
C433 VTAIL.n336 B 0.010025f
C434 VTAIL.n337 B 0.018657f
C435 VTAIL.n338 B 0.018657f
C436 VTAIL.n339 B 0.010025f
C437 VTAIL.n340 B 0.010615f
C438 VTAIL.n341 B 0.023696f
C439 VTAIL.n342 B 0.049518f
C440 VTAIL.n343 B 0.010615f
C441 VTAIL.n344 B 0.010025f
C442 VTAIL.n345 B 0.045163f
C443 VTAIL.n346 B 0.027585f
C444 VTAIL.n347 B 1.26347f
C445 VTAIL.t6 B 0.227635f
C446 VTAIL.t1 B 0.227635f
C447 VTAIL.n348 B 2.00748f
C448 VTAIL.n349 B 0.373397f
C449 VTAIL.n350 B 0.025217f
C450 VTAIL.n351 B 0.018657f
C451 VTAIL.n352 B 0.010025f
C452 VTAIL.n353 B 0.023696f
C453 VTAIL.n354 B 0.01032f
C454 VTAIL.n355 B 0.018657f
C455 VTAIL.n356 B 0.01032f
C456 VTAIL.n357 B 0.010025f
C457 VTAIL.n358 B 0.023696f
C458 VTAIL.n359 B 0.023696f
C459 VTAIL.n360 B 0.010615f
C460 VTAIL.n361 B 0.018657f
C461 VTAIL.n362 B 0.010025f
C462 VTAIL.n363 B 0.023696f
C463 VTAIL.n364 B 0.010615f
C464 VTAIL.n365 B 0.018657f
C465 VTAIL.n366 B 0.010025f
C466 VTAIL.n367 B 0.023696f
C467 VTAIL.n368 B 0.010615f
C468 VTAIL.n369 B 0.018657f
C469 VTAIL.n370 B 0.010025f
C470 VTAIL.n371 B 0.023696f
C471 VTAIL.n372 B 0.010615f
C472 VTAIL.n373 B 0.018657f
C473 VTAIL.n374 B 0.010025f
C474 VTAIL.n375 B 0.023696f
C475 VTAIL.n376 B 0.010615f
C476 VTAIL.n377 B 1.25146f
C477 VTAIL.n378 B 0.010025f
C478 VTAIL.t2 B 0.0391f
C479 VTAIL.n379 B 0.123742f
C480 VTAIL.n380 B 0.013998f
C481 VTAIL.n381 B 0.017772f
C482 VTAIL.n382 B 0.023696f
C483 VTAIL.n383 B 0.010615f
C484 VTAIL.n384 B 0.010025f
C485 VTAIL.n385 B 0.018657f
C486 VTAIL.n386 B 0.018657f
C487 VTAIL.n387 B 0.010025f
C488 VTAIL.n388 B 0.010615f
C489 VTAIL.n389 B 0.023696f
C490 VTAIL.n390 B 0.023696f
C491 VTAIL.n391 B 0.010615f
C492 VTAIL.n392 B 0.010025f
C493 VTAIL.n393 B 0.018657f
C494 VTAIL.n394 B 0.018657f
C495 VTAIL.n395 B 0.010025f
C496 VTAIL.n396 B 0.010615f
C497 VTAIL.n397 B 0.023696f
C498 VTAIL.n398 B 0.023696f
C499 VTAIL.n399 B 0.010615f
C500 VTAIL.n400 B 0.010025f
C501 VTAIL.n401 B 0.018657f
C502 VTAIL.n402 B 0.018657f
C503 VTAIL.n403 B 0.010025f
C504 VTAIL.n404 B 0.010615f
C505 VTAIL.n405 B 0.023696f
C506 VTAIL.n406 B 0.023696f
C507 VTAIL.n407 B 0.010615f
C508 VTAIL.n408 B 0.010025f
C509 VTAIL.n409 B 0.018657f
C510 VTAIL.n410 B 0.018657f
C511 VTAIL.n411 B 0.010025f
C512 VTAIL.n412 B 0.010615f
C513 VTAIL.n413 B 0.023696f
C514 VTAIL.n414 B 0.023696f
C515 VTAIL.n415 B 0.010615f
C516 VTAIL.n416 B 0.010025f
C517 VTAIL.n417 B 0.018657f
C518 VTAIL.n418 B 0.018657f
C519 VTAIL.n419 B 0.010025f
C520 VTAIL.n420 B 0.010615f
C521 VTAIL.n421 B 0.023696f
C522 VTAIL.n422 B 0.023696f
C523 VTAIL.n423 B 0.010615f
C524 VTAIL.n424 B 0.010025f
C525 VTAIL.n425 B 0.018657f
C526 VTAIL.n426 B 0.018657f
C527 VTAIL.n427 B 0.010025f
C528 VTAIL.n428 B 0.010615f
C529 VTAIL.n429 B 0.023696f
C530 VTAIL.n430 B 0.049518f
C531 VTAIL.n431 B 0.010615f
C532 VTAIL.n432 B 0.010025f
C533 VTAIL.n433 B 0.045163f
C534 VTAIL.n434 B 0.027585f
C535 VTAIL.n435 B 0.141724f
C536 VTAIL.n436 B 0.025217f
C537 VTAIL.n437 B 0.018657f
C538 VTAIL.n438 B 0.010025f
C539 VTAIL.n439 B 0.023696f
C540 VTAIL.n440 B 0.01032f
C541 VTAIL.n441 B 0.018657f
C542 VTAIL.n442 B 0.01032f
C543 VTAIL.n443 B 0.010025f
C544 VTAIL.n444 B 0.023696f
C545 VTAIL.n445 B 0.023696f
C546 VTAIL.n446 B 0.010615f
C547 VTAIL.n447 B 0.018657f
C548 VTAIL.n448 B 0.010025f
C549 VTAIL.n449 B 0.023696f
C550 VTAIL.n450 B 0.010615f
C551 VTAIL.n451 B 0.018657f
C552 VTAIL.n452 B 0.010025f
C553 VTAIL.n453 B 0.023696f
C554 VTAIL.n454 B 0.010615f
C555 VTAIL.n455 B 0.018657f
C556 VTAIL.n456 B 0.010025f
C557 VTAIL.n457 B 0.023696f
C558 VTAIL.n458 B 0.010615f
C559 VTAIL.n459 B 0.018657f
C560 VTAIL.n460 B 0.010025f
C561 VTAIL.n461 B 0.023696f
C562 VTAIL.n462 B 0.010615f
C563 VTAIL.n463 B 1.25146f
C564 VTAIL.n464 B 0.010025f
C565 VTAIL.t11 B 0.0391f
C566 VTAIL.n465 B 0.123742f
C567 VTAIL.n466 B 0.013998f
C568 VTAIL.n467 B 0.017772f
C569 VTAIL.n468 B 0.023696f
C570 VTAIL.n469 B 0.010615f
C571 VTAIL.n470 B 0.010025f
C572 VTAIL.n471 B 0.018657f
C573 VTAIL.n472 B 0.018657f
C574 VTAIL.n473 B 0.010025f
C575 VTAIL.n474 B 0.010615f
C576 VTAIL.n475 B 0.023696f
C577 VTAIL.n476 B 0.023696f
C578 VTAIL.n477 B 0.010615f
C579 VTAIL.n478 B 0.010025f
C580 VTAIL.n479 B 0.018657f
C581 VTAIL.n480 B 0.018657f
C582 VTAIL.n481 B 0.010025f
C583 VTAIL.n482 B 0.010615f
C584 VTAIL.n483 B 0.023696f
C585 VTAIL.n484 B 0.023696f
C586 VTAIL.n485 B 0.010615f
C587 VTAIL.n486 B 0.010025f
C588 VTAIL.n487 B 0.018657f
C589 VTAIL.n488 B 0.018657f
C590 VTAIL.n489 B 0.010025f
C591 VTAIL.n490 B 0.010615f
C592 VTAIL.n491 B 0.023696f
C593 VTAIL.n492 B 0.023696f
C594 VTAIL.n493 B 0.010615f
C595 VTAIL.n494 B 0.010025f
C596 VTAIL.n495 B 0.018657f
C597 VTAIL.n496 B 0.018657f
C598 VTAIL.n497 B 0.010025f
C599 VTAIL.n498 B 0.010615f
C600 VTAIL.n499 B 0.023696f
C601 VTAIL.n500 B 0.023696f
C602 VTAIL.n501 B 0.010615f
C603 VTAIL.n502 B 0.010025f
C604 VTAIL.n503 B 0.018657f
C605 VTAIL.n504 B 0.018657f
C606 VTAIL.n505 B 0.010025f
C607 VTAIL.n506 B 0.010615f
C608 VTAIL.n507 B 0.023696f
C609 VTAIL.n508 B 0.023696f
C610 VTAIL.n509 B 0.010615f
C611 VTAIL.n510 B 0.010025f
C612 VTAIL.n511 B 0.018657f
C613 VTAIL.n512 B 0.018657f
C614 VTAIL.n513 B 0.010025f
C615 VTAIL.n514 B 0.010615f
C616 VTAIL.n515 B 0.023696f
C617 VTAIL.n516 B 0.049518f
C618 VTAIL.n517 B 0.010615f
C619 VTAIL.n518 B 0.010025f
C620 VTAIL.n519 B 0.045163f
C621 VTAIL.n520 B 0.027585f
C622 VTAIL.n521 B 0.141724f
C623 VTAIL.t13 B 0.227635f
C624 VTAIL.t8 B 0.227635f
C625 VTAIL.n522 B 2.00748f
C626 VTAIL.n523 B 0.373397f
C627 VTAIL.n524 B 0.025217f
C628 VTAIL.n525 B 0.018657f
C629 VTAIL.n526 B 0.010025f
C630 VTAIL.n527 B 0.023696f
C631 VTAIL.n528 B 0.01032f
C632 VTAIL.n529 B 0.018657f
C633 VTAIL.n530 B 0.01032f
C634 VTAIL.n531 B 0.010025f
C635 VTAIL.n532 B 0.023696f
C636 VTAIL.n533 B 0.023696f
C637 VTAIL.n534 B 0.010615f
C638 VTAIL.n535 B 0.018657f
C639 VTAIL.n536 B 0.010025f
C640 VTAIL.n537 B 0.023696f
C641 VTAIL.n538 B 0.010615f
C642 VTAIL.n539 B 0.018657f
C643 VTAIL.n540 B 0.010025f
C644 VTAIL.n541 B 0.023696f
C645 VTAIL.n542 B 0.010615f
C646 VTAIL.n543 B 0.018657f
C647 VTAIL.n544 B 0.010025f
C648 VTAIL.n545 B 0.023696f
C649 VTAIL.n546 B 0.010615f
C650 VTAIL.n547 B 0.018657f
C651 VTAIL.n548 B 0.010025f
C652 VTAIL.n549 B 0.023696f
C653 VTAIL.n550 B 0.010615f
C654 VTAIL.n551 B 1.25146f
C655 VTAIL.n552 B 0.010025f
C656 VTAIL.t12 B 0.0391f
C657 VTAIL.n553 B 0.123742f
C658 VTAIL.n554 B 0.013998f
C659 VTAIL.n555 B 0.017772f
C660 VTAIL.n556 B 0.023696f
C661 VTAIL.n557 B 0.010615f
C662 VTAIL.n558 B 0.010025f
C663 VTAIL.n559 B 0.018657f
C664 VTAIL.n560 B 0.018657f
C665 VTAIL.n561 B 0.010025f
C666 VTAIL.n562 B 0.010615f
C667 VTAIL.n563 B 0.023696f
C668 VTAIL.n564 B 0.023696f
C669 VTAIL.n565 B 0.010615f
C670 VTAIL.n566 B 0.010025f
C671 VTAIL.n567 B 0.018657f
C672 VTAIL.n568 B 0.018657f
C673 VTAIL.n569 B 0.010025f
C674 VTAIL.n570 B 0.010615f
C675 VTAIL.n571 B 0.023696f
C676 VTAIL.n572 B 0.023696f
C677 VTAIL.n573 B 0.010615f
C678 VTAIL.n574 B 0.010025f
C679 VTAIL.n575 B 0.018657f
C680 VTAIL.n576 B 0.018657f
C681 VTAIL.n577 B 0.010025f
C682 VTAIL.n578 B 0.010615f
C683 VTAIL.n579 B 0.023696f
C684 VTAIL.n580 B 0.023696f
C685 VTAIL.n581 B 0.010615f
C686 VTAIL.n582 B 0.010025f
C687 VTAIL.n583 B 0.018657f
C688 VTAIL.n584 B 0.018657f
C689 VTAIL.n585 B 0.010025f
C690 VTAIL.n586 B 0.010615f
C691 VTAIL.n587 B 0.023696f
C692 VTAIL.n588 B 0.023696f
C693 VTAIL.n589 B 0.010615f
C694 VTAIL.n590 B 0.010025f
C695 VTAIL.n591 B 0.018657f
C696 VTAIL.n592 B 0.018657f
C697 VTAIL.n593 B 0.010025f
C698 VTAIL.n594 B 0.010615f
C699 VTAIL.n595 B 0.023696f
C700 VTAIL.n596 B 0.023696f
C701 VTAIL.n597 B 0.010615f
C702 VTAIL.n598 B 0.010025f
C703 VTAIL.n599 B 0.018657f
C704 VTAIL.n600 B 0.018657f
C705 VTAIL.n601 B 0.010025f
C706 VTAIL.n602 B 0.010615f
C707 VTAIL.n603 B 0.023696f
C708 VTAIL.n604 B 0.049518f
C709 VTAIL.n605 B 0.010615f
C710 VTAIL.n606 B 0.010025f
C711 VTAIL.n607 B 0.045163f
C712 VTAIL.n608 B 0.027585f
C713 VTAIL.n609 B 1.26347f
C714 VTAIL.n610 B 0.025217f
C715 VTAIL.n611 B 0.018657f
C716 VTAIL.n612 B 0.010025f
C717 VTAIL.n613 B 0.023696f
C718 VTAIL.n614 B 0.01032f
C719 VTAIL.n615 B 0.018657f
C720 VTAIL.n616 B 0.010615f
C721 VTAIL.n617 B 0.023696f
C722 VTAIL.n618 B 0.010615f
C723 VTAIL.n619 B 0.018657f
C724 VTAIL.n620 B 0.010025f
C725 VTAIL.n621 B 0.023696f
C726 VTAIL.n622 B 0.010615f
C727 VTAIL.n623 B 0.018657f
C728 VTAIL.n624 B 0.010025f
C729 VTAIL.n625 B 0.023696f
C730 VTAIL.n626 B 0.010615f
C731 VTAIL.n627 B 0.018657f
C732 VTAIL.n628 B 0.010025f
C733 VTAIL.n629 B 0.023696f
C734 VTAIL.n630 B 0.010615f
C735 VTAIL.n631 B 0.018657f
C736 VTAIL.n632 B 0.010025f
C737 VTAIL.n633 B 0.023696f
C738 VTAIL.n634 B 0.010615f
C739 VTAIL.n635 B 1.25146f
C740 VTAIL.n636 B 0.010025f
C741 VTAIL.t5 B 0.0391f
C742 VTAIL.n637 B 0.123742f
C743 VTAIL.n638 B 0.013998f
C744 VTAIL.n639 B 0.017772f
C745 VTAIL.n640 B 0.023696f
C746 VTAIL.n641 B 0.010615f
C747 VTAIL.n642 B 0.010025f
C748 VTAIL.n643 B 0.018657f
C749 VTAIL.n644 B 0.018657f
C750 VTAIL.n645 B 0.010025f
C751 VTAIL.n646 B 0.010615f
C752 VTAIL.n647 B 0.023696f
C753 VTAIL.n648 B 0.023696f
C754 VTAIL.n649 B 0.010615f
C755 VTAIL.n650 B 0.010025f
C756 VTAIL.n651 B 0.018657f
C757 VTAIL.n652 B 0.018657f
C758 VTAIL.n653 B 0.010025f
C759 VTAIL.n654 B 0.010615f
C760 VTAIL.n655 B 0.023696f
C761 VTAIL.n656 B 0.023696f
C762 VTAIL.n657 B 0.010615f
C763 VTAIL.n658 B 0.010025f
C764 VTAIL.n659 B 0.018657f
C765 VTAIL.n660 B 0.018657f
C766 VTAIL.n661 B 0.010025f
C767 VTAIL.n662 B 0.010615f
C768 VTAIL.n663 B 0.023696f
C769 VTAIL.n664 B 0.023696f
C770 VTAIL.n665 B 0.010615f
C771 VTAIL.n666 B 0.010025f
C772 VTAIL.n667 B 0.018657f
C773 VTAIL.n668 B 0.018657f
C774 VTAIL.n669 B 0.010025f
C775 VTAIL.n670 B 0.010615f
C776 VTAIL.n671 B 0.023696f
C777 VTAIL.n672 B 0.023696f
C778 VTAIL.n673 B 0.010615f
C779 VTAIL.n674 B 0.010025f
C780 VTAIL.n675 B 0.018657f
C781 VTAIL.n676 B 0.018657f
C782 VTAIL.n677 B 0.010025f
C783 VTAIL.n678 B 0.010025f
C784 VTAIL.n679 B 0.010615f
C785 VTAIL.n680 B 0.023696f
C786 VTAIL.n681 B 0.023696f
C787 VTAIL.n682 B 0.023696f
C788 VTAIL.n683 B 0.01032f
C789 VTAIL.n684 B 0.010025f
C790 VTAIL.n685 B 0.018657f
C791 VTAIL.n686 B 0.018657f
C792 VTAIL.n687 B 0.010025f
C793 VTAIL.n688 B 0.010615f
C794 VTAIL.n689 B 0.023696f
C795 VTAIL.n690 B 0.049518f
C796 VTAIL.n691 B 0.010615f
C797 VTAIL.n692 B 0.010025f
C798 VTAIL.n693 B 0.045163f
C799 VTAIL.n694 B 0.027585f
C800 VTAIL.n695 B 1.25998f
C801 VP.n0 B 0.030393f
C802 VP.t4 B 1.96869f
C803 VP.n1 B 0.05302f
C804 VP.n2 B 0.030393f
C805 VP.t1 B 1.96869f
C806 VP.n3 B 0.056193f
C807 VP.n4 B 0.030393f
C808 VP.n5 B 0.04692f
C809 VP.n6 B 0.030393f
C810 VP.t0 B 1.96869f
C811 VP.n7 B 0.05302f
C812 VP.n8 B 0.030393f
C813 VP.t3 B 1.96869f
C814 VP.n9 B 0.056193f
C815 VP.t7 B 2.07516f
C816 VP.t6 B 1.96869f
C817 VP.n10 B 0.766106f
C818 VP.n11 B 0.7631f
C819 VP.n12 B 0.194818f
C820 VP.n13 B 0.030393f
C821 VP.n14 B 0.024548f
C822 VP.n15 B 0.056193f
C823 VP.n16 B 0.698534f
C824 VP.n17 B 0.032433f
C825 VP.n18 B 0.030393f
C826 VP.n19 B 0.030393f
C827 VP.n20 B 0.030393f
C828 VP.n21 B 0.033097f
C829 VP.n22 B 0.04692f
C830 VP.n23 B 0.768239f
C831 VP.n24 B 1.58192f
C832 VP.t2 B 1.96869f
C833 VP.n25 B 0.768239f
C834 VP.n26 B 1.60451f
C835 VP.n27 B 0.030393f
C836 VP.n28 B 0.030393f
C837 VP.n29 B 0.033097f
C838 VP.n30 B 0.05302f
C839 VP.t5 B 1.96869f
C840 VP.n31 B 0.698534f
C841 VP.n32 B 0.032433f
C842 VP.n33 B 0.030393f
C843 VP.n34 B 0.030393f
C844 VP.n35 B 0.030393f
C845 VP.n36 B 0.024548f
C846 VP.n37 B 0.056193f
C847 VP.n38 B 0.698534f
C848 VP.n39 B 0.032433f
C849 VP.n40 B 0.030393f
C850 VP.n41 B 0.030393f
C851 VP.n42 B 0.030393f
C852 VP.n43 B 0.033097f
C853 VP.n44 B 0.04692f
C854 VP.n45 B 0.768239f
C855 VP.n46 B 0.028017f
.ends

