* NGSPICE file created from diff_pair_sample_1293.ext - technology: sky130A

.subckt diff_pair_sample_1293 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=1.05
X1 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=1.05
X2 VTAIL.t12 VP.t1 VDD1.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X3 VTAIL.t4 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X4 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=1.05
X5 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X6 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=1.05
X7 VDD2.t5 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X8 VDD1.t7 VP.t2 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=1.05
X9 VTAIL.t17 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X10 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=1.05
X11 VTAIL.t7 VN.t5 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=1.05
X13 VDD1.t5 VP.t4 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X14 VTAIL.t19 VN.t6 VDD2.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=1.05
X16 VTAIL.t10 VP.t5 VDD1.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X17 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=1.05
X18 VDD1.t3 VP.t6 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=1.05
X19 VTAIL.t8 VN.t8 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X20 VDD1.t2 VP.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=1.05
X21 VDD2.t0 VN.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=1.05
X22 VTAIL.t18 VP.t8 VDD1.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
X23 VDD1.t0 VP.t9 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.99165 pd=6.34 as=0.99165 ps=6.34 w=6.01 l=1.05
R0 VP.n9 VP.t6 190.731
R1 VP.n25 VP.t7 175.587
R2 VP.n41 VP.t2 175.587
R3 VP.n22 VP.t0 175.587
R4 VP.n10 VP.n7 161.3
R5 VP.n12 VP.n11 161.3
R6 VP.n13 VP.n6 161.3
R7 VP.n16 VP.n15 161.3
R8 VP.n17 VP.n5 161.3
R9 VP.n19 VP.n18 161.3
R10 VP.n21 VP.n4 161.3
R11 VP.n40 VP.n0 161.3
R12 VP.n38 VP.n37 161.3
R13 VP.n36 VP.n1 161.3
R14 VP.n35 VP.n34 161.3
R15 VP.n32 VP.n2 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n29 VP.n3 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.t3 137.945
R20 VP.n33 VP.t9 137.945
R21 VP.n39 VP.t8 137.945
R22 VP.n20 VP.t1 137.945
R23 VP.n14 VP.t4 137.945
R24 VP.n8 VP.t5 137.945
R25 VP.n23 VP.n22 80.6037
R26 VP.n42 VP.n41 80.6037
R27 VP.n25 VP.n24 80.6037
R28 VP.n27 VP.n25 55.7853
R29 VP.n41 VP.n40 55.7853
R30 VP.n22 VP.n21 55.7853
R31 VP.n9 VP.n8 48.3043
R32 VP.n32 VP.n31 46.321
R33 VP.n34 VP.n1 46.321
R34 VP.n15 VP.n5 46.321
R35 VP.n13 VP.n12 46.321
R36 VP.n10 VP.n9 43.9769
R37 VP.n24 VP.n23 40.3878
R38 VP.n31 VP.n3 34.6658
R39 VP.n38 VP.n1 34.6658
R40 VP.n19 VP.n5 34.6658
R41 VP.n12 VP.n7 34.6658
R42 VP.n27 VP.n26 18.1061
R43 VP.n40 VP.n39 18.1061
R44 VP.n21 VP.n20 18.1061
R45 VP.n33 VP.n32 12.234
R46 VP.n34 VP.n33 12.234
R47 VP.n14 VP.n13 12.234
R48 VP.n15 VP.n14 12.234
R49 VP.n26 VP.n3 6.36192
R50 VP.n39 VP.n38 6.36192
R51 VP.n20 VP.n19 6.36192
R52 VP.n8 VP.n7 6.36192
R53 VP.n23 VP.n4 0.285035
R54 VP.n28 VP.n24 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n11 VP.n10 0.189894
R57 VP.n11 VP.n6 0.189894
R58 VP.n16 VP.n6 0.189894
R59 VP.n17 VP.n16 0.189894
R60 VP.n18 VP.n17 0.189894
R61 VP.n18 VP.n4 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n30 VP.n29 0.189894
R64 VP.n30 VP.n2 0.189894
R65 VP.n35 VP.n2 0.189894
R66 VP.n36 VP.n35 0.189894
R67 VP.n37 VP.n36 0.189894
R68 VP.n37 VP.n0 0.189894
R69 VP VP.n42 0.146778
R70 VTAIL.n136 VTAIL.n110 289.615
R71 VTAIL.n28 VTAIL.n2 289.615
R72 VTAIL.n104 VTAIL.n78 289.615
R73 VTAIL.n68 VTAIL.n42 289.615
R74 VTAIL.n121 VTAIL.n120 185
R75 VTAIL.n118 VTAIL.n117 185
R76 VTAIL.n127 VTAIL.n126 185
R77 VTAIL.n129 VTAIL.n128 185
R78 VTAIL.n114 VTAIL.n113 185
R79 VTAIL.n135 VTAIL.n134 185
R80 VTAIL.n137 VTAIL.n136 185
R81 VTAIL.n13 VTAIL.n12 185
R82 VTAIL.n10 VTAIL.n9 185
R83 VTAIL.n19 VTAIL.n18 185
R84 VTAIL.n21 VTAIL.n20 185
R85 VTAIL.n6 VTAIL.n5 185
R86 VTAIL.n27 VTAIL.n26 185
R87 VTAIL.n29 VTAIL.n28 185
R88 VTAIL.n105 VTAIL.n104 185
R89 VTAIL.n103 VTAIL.n102 185
R90 VTAIL.n82 VTAIL.n81 185
R91 VTAIL.n97 VTAIL.n96 185
R92 VTAIL.n95 VTAIL.n94 185
R93 VTAIL.n86 VTAIL.n85 185
R94 VTAIL.n89 VTAIL.n88 185
R95 VTAIL.n69 VTAIL.n68 185
R96 VTAIL.n67 VTAIL.n66 185
R97 VTAIL.n46 VTAIL.n45 185
R98 VTAIL.n61 VTAIL.n60 185
R99 VTAIL.n59 VTAIL.n58 185
R100 VTAIL.n50 VTAIL.n49 185
R101 VTAIL.n53 VTAIL.n52 185
R102 VTAIL.t1 VTAIL.n119 147.661
R103 VTAIL.t16 VTAIL.n11 147.661
R104 VTAIL.t15 VTAIL.n87 147.661
R105 VTAIL.t2 VTAIL.n51 147.661
R106 VTAIL.n120 VTAIL.n117 104.615
R107 VTAIL.n127 VTAIL.n117 104.615
R108 VTAIL.n128 VTAIL.n127 104.615
R109 VTAIL.n128 VTAIL.n113 104.615
R110 VTAIL.n135 VTAIL.n113 104.615
R111 VTAIL.n136 VTAIL.n135 104.615
R112 VTAIL.n12 VTAIL.n9 104.615
R113 VTAIL.n19 VTAIL.n9 104.615
R114 VTAIL.n20 VTAIL.n19 104.615
R115 VTAIL.n20 VTAIL.n5 104.615
R116 VTAIL.n27 VTAIL.n5 104.615
R117 VTAIL.n28 VTAIL.n27 104.615
R118 VTAIL.n104 VTAIL.n103 104.615
R119 VTAIL.n103 VTAIL.n81 104.615
R120 VTAIL.n96 VTAIL.n81 104.615
R121 VTAIL.n96 VTAIL.n95 104.615
R122 VTAIL.n95 VTAIL.n85 104.615
R123 VTAIL.n88 VTAIL.n85 104.615
R124 VTAIL.n68 VTAIL.n67 104.615
R125 VTAIL.n67 VTAIL.n45 104.615
R126 VTAIL.n60 VTAIL.n45 104.615
R127 VTAIL.n60 VTAIL.n59 104.615
R128 VTAIL.n59 VTAIL.n49 104.615
R129 VTAIL.n52 VTAIL.n49 104.615
R130 VTAIL.n120 VTAIL.t1 52.3082
R131 VTAIL.n12 VTAIL.t16 52.3082
R132 VTAIL.n88 VTAIL.t15 52.3082
R133 VTAIL.n52 VTAIL.t2 52.3082
R134 VTAIL.n77 VTAIL.n76 50.706
R135 VTAIL.n75 VTAIL.n74 50.706
R136 VTAIL.n41 VTAIL.n40 50.706
R137 VTAIL.n39 VTAIL.n38 50.706
R138 VTAIL.n143 VTAIL.n142 50.7058
R139 VTAIL.n1 VTAIL.n0 50.7058
R140 VTAIL.n35 VTAIL.n34 50.7058
R141 VTAIL.n37 VTAIL.n36 50.7058
R142 VTAIL.n141 VTAIL.n140 32.3793
R143 VTAIL.n33 VTAIL.n32 32.3793
R144 VTAIL.n109 VTAIL.n108 32.3793
R145 VTAIL.n73 VTAIL.n72 32.3793
R146 VTAIL.n39 VTAIL.n37 19.9272
R147 VTAIL.n141 VTAIL.n109 18.7376
R148 VTAIL.n121 VTAIL.n119 15.6674
R149 VTAIL.n13 VTAIL.n11 15.6674
R150 VTAIL.n89 VTAIL.n87 15.6674
R151 VTAIL.n53 VTAIL.n51 15.6674
R152 VTAIL.n122 VTAIL.n118 12.8005
R153 VTAIL.n14 VTAIL.n10 12.8005
R154 VTAIL.n90 VTAIL.n86 12.8005
R155 VTAIL.n54 VTAIL.n50 12.8005
R156 VTAIL.n126 VTAIL.n125 12.0247
R157 VTAIL.n18 VTAIL.n17 12.0247
R158 VTAIL.n94 VTAIL.n93 12.0247
R159 VTAIL.n58 VTAIL.n57 12.0247
R160 VTAIL.n129 VTAIL.n116 11.249
R161 VTAIL.n21 VTAIL.n8 11.249
R162 VTAIL.n97 VTAIL.n84 11.249
R163 VTAIL.n61 VTAIL.n48 11.249
R164 VTAIL.n130 VTAIL.n114 10.4732
R165 VTAIL.n22 VTAIL.n6 10.4732
R166 VTAIL.n98 VTAIL.n82 10.4732
R167 VTAIL.n62 VTAIL.n46 10.4732
R168 VTAIL.n134 VTAIL.n133 9.69747
R169 VTAIL.n26 VTAIL.n25 9.69747
R170 VTAIL.n102 VTAIL.n101 9.69747
R171 VTAIL.n66 VTAIL.n65 9.69747
R172 VTAIL.n140 VTAIL.n139 9.45567
R173 VTAIL.n32 VTAIL.n31 9.45567
R174 VTAIL.n108 VTAIL.n107 9.45567
R175 VTAIL.n72 VTAIL.n71 9.45567
R176 VTAIL.n139 VTAIL.n138 9.3005
R177 VTAIL.n112 VTAIL.n111 9.3005
R178 VTAIL.n133 VTAIL.n132 9.3005
R179 VTAIL.n131 VTAIL.n130 9.3005
R180 VTAIL.n116 VTAIL.n115 9.3005
R181 VTAIL.n125 VTAIL.n124 9.3005
R182 VTAIL.n123 VTAIL.n122 9.3005
R183 VTAIL.n31 VTAIL.n30 9.3005
R184 VTAIL.n4 VTAIL.n3 9.3005
R185 VTAIL.n25 VTAIL.n24 9.3005
R186 VTAIL.n23 VTAIL.n22 9.3005
R187 VTAIL.n8 VTAIL.n7 9.3005
R188 VTAIL.n17 VTAIL.n16 9.3005
R189 VTAIL.n15 VTAIL.n14 9.3005
R190 VTAIL.n107 VTAIL.n106 9.3005
R191 VTAIL.n80 VTAIL.n79 9.3005
R192 VTAIL.n101 VTAIL.n100 9.3005
R193 VTAIL.n99 VTAIL.n98 9.3005
R194 VTAIL.n84 VTAIL.n83 9.3005
R195 VTAIL.n93 VTAIL.n92 9.3005
R196 VTAIL.n91 VTAIL.n90 9.3005
R197 VTAIL.n71 VTAIL.n70 9.3005
R198 VTAIL.n44 VTAIL.n43 9.3005
R199 VTAIL.n65 VTAIL.n64 9.3005
R200 VTAIL.n63 VTAIL.n62 9.3005
R201 VTAIL.n48 VTAIL.n47 9.3005
R202 VTAIL.n57 VTAIL.n56 9.3005
R203 VTAIL.n55 VTAIL.n54 9.3005
R204 VTAIL.n137 VTAIL.n112 8.92171
R205 VTAIL.n29 VTAIL.n4 8.92171
R206 VTAIL.n105 VTAIL.n80 8.92171
R207 VTAIL.n69 VTAIL.n44 8.92171
R208 VTAIL.n138 VTAIL.n110 8.14595
R209 VTAIL.n30 VTAIL.n2 8.14595
R210 VTAIL.n106 VTAIL.n78 8.14595
R211 VTAIL.n70 VTAIL.n42 8.14595
R212 VTAIL.n140 VTAIL.n110 5.81868
R213 VTAIL.n32 VTAIL.n2 5.81868
R214 VTAIL.n108 VTAIL.n78 5.81868
R215 VTAIL.n72 VTAIL.n42 5.81868
R216 VTAIL.n138 VTAIL.n137 5.04292
R217 VTAIL.n30 VTAIL.n29 5.04292
R218 VTAIL.n106 VTAIL.n105 5.04292
R219 VTAIL.n70 VTAIL.n69 5.04292
R220 VTAIL.n123 VTAIL.n119 4.38594
R221 VTAIL.n15 VTAIL.n11 4.38594
R222 VTAIL.n91 VTAIL.n87 4.38594
R223 VTAIL.n55 VTAIL.n51 4.38594
R224 VTAIL.n134 VTAIL.n112 4.26717
R225 VTAIL.n26 VTAIL.n4 4.26717
R226 VTAIL.n102 VTAIL.n80 4.26717
R227 VTAIL.n66 VTAIL.n44 4.26717
R228 VTAIL.n133 VTAIL.n114 3.49141
R229 VTAIL.n25 VTAIL.n6 3.49141
R230 VTAIL.n101 VTAIL.n82 3.49141
R231 VTAIL.n65 VTAIL.n46 3.49141
R232 VTAIL.n142 VTAIL.t6 3.29501
R233 VTAIL.n142 VTAIL.t7 3.29501
R234 VTAIL.n0 VTAIL.t0 3.29501
R235 VTAIL.n0 VTAIL.t8 3.29501
R236 VTAIL.n34 VTAIL.t9 3.29501
R237 VTAIL.n34 VTAIL.t18 3.29501
R238 VTAIL.n36 VTAIL.t13 3.29501
R239 VTAIL.n36 VTAIL.t17 3.29501
R240 VTAIL.n76 VTAIL.t14 3.29501
R241 VTAIL.n76 VTAIL.t12 3.29501
R242 VTAIL.n74 VTAIL.t11 3.29501
R243 VTAIL.n74 VTAIL.t10 3.29501
R244 VTAIL.n40 VTAIL.t5 3.29501
R245 VTAIL.n40 VTAIL.t19 3.29501
R246 VTAIL.n38 VTAIL.t3 3.29501
R247 VTAIL.n38 VTAIL.t4 3.29501
R248 VTAIL.n130 VTAIL.n129 2.71565
R249 VTAIL.n22 VTAIL.n21 2.71565
R250 VTAIL.n98 VTAIL.n97 2.71565
R251 VTAIL.n62 VTAIL.n61 2.71565
R252 VTAIL.n126 VTAIL.n116 1.93989
R253 VTAIL.n18 VTAIL.n8 1.93989
R254 VTAIL.n94 VTAIL.n84 1.93989
R255 VTAIL.n58 VTAIL.n48 1.93989
R256 VTAIL.n41 VTAIL.n39 1.19016
R257 VTAIL.n73 VTAIL.n41 1.19016
R258 VTAIL.n77 VTAIL.n75 1.19016
R259 VTAIL.n109 VTAIL.n77 1.19016
R260 VTAIL.n37 VTAIL.n35 1.19016
R261 VTAIL.n35 VTAIL.n33 1.19016
R262 VTAIL.n143 VTAIL.n141 1.19016
R263 VTAIL.n125 VTAIL.n118 1.16414
R264 VTAIL.n17 VTAIL.n10 1.16414
R265 VTAIL.n93 VTAIL.n86 1.16414
R266 VTAIL.n57 VTAIL.n50 1.16414
R267 VTAIL.n75 VTAIL.n73 1.06516
R268 VTAIL.n33 VTAIL.n1 1.06516
R269 VTAIL VTAIL.n1 0.950931
R270 VTAIL.n122 VTAIL.n121 0.388379
R271 VTAIL.n14 VTAIL.n13 0.388379
R272 VTAIL.n90 VTAIL.n89 0.388379
R273 VTAIL.n54 VTAIL.n53 0.388379
R274 VTAIL VTAIL.n143 0.239724
R275 VTAIL.n124 VTAIL.n123 0.155672
R276 VTAIL.n124 VTAIL.n115 0.155672
R277 VTAIL.n131 VTAIL.n115 0.155672
R278 VTAIL.n132 VTAIL.n131 0.155672
R279 VTAIL.n132 VTAIL.n111 0.155672
R280 VTAIL.n139 VTAIL.n111 0.155672
R281 VTAIL.n16 VTAIL.n15 0.155672
R282 VTAIL.n16 VTAIL.n7 0.155672
R283 VTAIL.n23 VTAIL.n7 0.155672
R284 VTAIL.n24 VTAIL.n23 0.155672
R285 VTAIL.n24 VTAIL.n3 0.155672
R286 VTAIL.n31 VTAIL.n3 0.155672
R287 VTAIL.n107 VTAIL.n79 0.155672
R288 VTAIL.n100 VTAIL.n79 0.155672
R289 VTAIL.n100 VTAIL.n99 0.155672
R290 VTAIL.n99 VTAIL.n83 0.155672
R291 VTAIL.n92 VTAIL.n83 0.155672
R292 VTAIL.n92 VTAIL.n91 0.155672
R293 VTAIL.n71 VTAIL.n43 0.155672
R294 VTAIL.n64 VTAIL.n43 0.155672
R295 VTAIL.n64 VTAIL.n63 0.155672
R296 VTAIL.n63 VTAIL.n47 0.155672
R297 VTAIL.n56 VTAIL.n47 0.155672
R298 VTAIL.n56 VTAIL.n55 0.155672
R299 VDD1.n26 VDD1.n0 289.615
R300 VDD1.n59 VDD1.n33 289.615
R301 VDD1.n27 VDD1.n26 185
R302 VDD1.n25 VDD1.n24 185
R303 VDD1.n4 VDD1.n3 185
R304 VDD1.n19 VDD1.n18 185
R305 VDD1.n17 VDD1.n16 185
R306 VDD1.n8 VDD1.n7 185
R307 VDD1.n11 VDD1.n10 185
R308 VDD1.n44 VDD1.n43 185
R309 VDD1.n41 VDD1.n40 185
R310 VDD1.n50 VDD1.n49 185
R311 VDD1.n52 VDD1.n51 185
R312 VDD1.n37 VDD1.n36 185
R313 VDD1.n58 VDD1.n57 185
R314 VDD1.n60 VDD1.n59 185
R315 VDD1.t3 VDD1.n9 147.661
R316 VDD1.t2 VDD1.n42 147.661
R317 VDD1.n26 VDD1.n25 104.615
R318 VDD1.n25 VDD1.n3 104.615
R319 VDD1.n18 VDD1.n3 104.615
R320 VDD1.n18 VDD1.n17 104.615
R321 VDD1.n17 VDD1.n7 104.615
R322 VDD1.n10 VDD1.n7 104.615
R323 VDD1.n43 VDD1.n40 104.615
R324 VDD1.n50 VDD1.n40 104.615
R325 VDD1.n51 VDD1.n50 104.615
R326 VDD1.n51 VDD1.n36 104.615
R327 VDD1.n58 VDD1.n36 104.615
R328 VDD1.n59 VDD1.n58 104.615
R329 VDD1.n67 VDD1.n66 68.2215
R330 VDD1.n32 VDD1.n31 67.3848
R331 VDD1.n69 VDD1.n68 67.3846
R332 VDD1.n65 VDD1.n64 67.3846
R333 VDD1.n10 VDD1.t3 52.3082
R334 VDD1.n43 VDD1.t2 52.3082
R335 VDD1.n32 VDD1.n30 50.2477
R336 VDD1.n65 VDD1.n63 50.2477
R337 VDD1.n69 VDD1.n67 35.725
R338 VDD1.n11 VDD1.n9 15.6674
R339 VDD1.n44 VDD1.n42 15.6674
R340 VDD1.n12 VDD1.n8 12.8005
R341 VDD1.n45 VDD1.n41 12.8005
R342 VDD1.n16 VDD1.n15 12.0247
R343 VDD1.n49 VDD1.n48 12.0247
R344 VDD1.n19 VDD1.n6 11.249
R345 VDD1.n52 VDD1.n39 11.249
R346 VDD1.n20 VDD1.n4 10.4732
R347 VDD1.n53 VDD1.n37 10.4732
R348 VDD1.n24 VDD1.n23 9.69747
R349 VDD1.n57 VDD1.n56 9.69747
R350 VDD1.n30 VDD1.n29 9.45567
R351 VDD1.n63 VDD1.n62 9.45567
R352 VDD1.n29 VDD1.n28 9.3005
R353 VDD1.n2 VDD1.n1 9.3005
R354 VDD1.n23 VDD1.n22 9.3005
R355 VDD1.n21 VDD1.n20 9.3005
R356 VDD1.n6 VDD1.n5 9.3005
R357 VDD1.n15 VDD1.n14 9.3005
R358 VDD1.n13 VDD1.n12 9.3005
R359 VDD1.n62 VDD1.n61 9.3005
R360 VDD1.n35 VDD1.n34 9.3005
R361 VDD1.n56 VDD1.n55 9.3005
R362 VDD1.n54 VDD1.n53 9.3005
R363 VDD1.n39 VDD1.n38 9.3005
R364 VDD1.n48 VDD1.n47 9.3005
R365 VDD1.n46 VDD1.n45 9.3005
R366 VDD1.n27 VDD1.n2 8.92171
R367 VDD1.n60 VDD1.n35 8.92171
R368 VDD1.n28 VDD1.n0 8.14595
R369 VDD1.n61 VDD1.n33 8.14595
R370 VDD1.n30 VDD1.n0 5.81868
R371 VDD1.n63 VDD1.n33 5.81868
R372 VDD1.n28 VDD1.n27 5.04292
R373 VDD1.n61 VDD1.n60 5.04292
R374 VDD1.n13 VDD1.n9 4.38594
R375 VDD1.n46 VDD1.n42 4.38594
R376 VDD1.n24 VDD1.n2 4.26717
R377 VDD1.n57 VDD1.n35 4.26717
R378 VDD1.n23 VDD1.n4 3.49141
R379 VDD1.n56 VDD1.n37 3.49141
R380 VDD1.n68 VDD1.t8 3.29501
R381 VDD1.n68 VDD1.t9 3.29501
R382 VDD1.n31 VDD1.t4 3.29501
R383 VDD1.n31 VDD1.t5 3.29501
R384 VDD1.n66 VDD1.t1 3.29501
R385 VDD1.n66 VDD1.t7 3.29501
R386 VDD1.n64 VDD1.t6 3.29501
R387 VDD1.n64 VDD1.t0 3.29501
R388 VDD1.n20 VDD1.n19 2.71565
R389 VDD1.n53 VDD1.n52 2.71565
R390 VDD1.n16 VDD1.n6 1.93989
R391 VDD1.n49 VDD1.n39 1.93989
R392 VDD1.n15 VDD1.n8 1.16414
R393 VDD1.n48 VDD1.n41 1.16414
R394 VDD1 VDD1.n69 0.834552
R395 VDD1.n12 VDD1.n11 0.388379
R396 VDD1.n45 VDD1.n44 0.388379
R397 VDD1 VDD1.n32 0.356103
R398 VDD1.n67 VDD1.n65 0.242568
R399 VDD1.n29 VDD1.n1 0.155672
R400 VDD1.n22 VDD1.n1 0.155672
R401 VDD1.n22 VDD1.n21 0.155672
R402 VDD1.n21 VDD1.n5 0.155672
R403 VDD1.n14 VDD1.n5 0.155672
R404 VDD1.n14 VDD1.n13 0.155672
R405 VDD1.n47 VDD1.n46 0.155672
R406 VDD1.n47 VDD1.n38 0.155672
R407 VDD1.n54 VDD1.n38 0.155672
R408 VDD1.n55 VDD1.n54 0.155672
R409 VDD1.n55 VDD1.n34 0.155672
R410 VDD1.n62 VDD1.n34 0.155672
R411 B.n561 B.n560 585
R412 B.n207 B.n90 585
R413 B.n206 B.n205 585
R414 B.n204 B.n203 585
R415 B.n202 B.n201 585
R416 B.n200 B.n199 585
R417 B.n198 B.n197 585
R418 B.n196 B.n195 585
R419 B.n194 B.n193 585
R420 B.n192 B.n191 585
R421 B.n190 B.n189 585
R422 B.n188 B.n187 585
R423 B.n186 B.n185 585
R424 B.n184 B.n183 585
R425 B.n182 B.n181 585
R426 B.n180 B.n179 585
R427 B.n178 B.n177 585
R428 B.n176 B.n175 585
R429 B.n174 B.n173 585
R430 B.n172 B.n171 585
R431 B.n170 B.n169 585
R432 B.n168 B.n167 585
R433 B.n166 B.n165 585
R434 B.n164 B.n163 585
R435 B.n162 B.n161 585
R436 B.n160 B.n159 585
R437 B.n158 B.n157 585
R438 B.n156 B.n155 585
R439 B.n154 B.n153 585
R440 B.n152 B.n151 585
R441 B.n150 B.n149 585
R442 B.n148 B.n147 585
R443 B.n146 B.n145 585
R444 B.n144 B.n143 585
R445 B.n142 B.n141 585
R446 B.n140 B.n139 585
R447 B.n138 B.n137 585
R448 B.n136 B.n135 585
R449 B.n134 B.n133 585
R450 B.n132 B.n131 585
R451 B.n130 B.n129 585
R452 B.n128 B.n127 585
R453 B.n126 B.n125 585
R454 B.n124 B.n123 585
R455 B.n122 B.n121 585
R456 B.n120 B.n119 585
R457 B.n118 B.n117 585
R458 B.n116 B.n115 585
R459 B.n114 B.n113 585
R460 B.n112 B.n111 585
R461 B.n110 B.n109 585
R462 B.n108 B.n107 585
R463 B.n106 B.n105 585
R464 B.n104 B.n103 585
R465 B.n102 B.n101 585
R466 B.n100 B.n99 585
R467 B.n98 B.n97 585
R468 B.n60 B.n59 585
R469 B.n559 B.n61 585
R470 B.n564 B.n61 585
R471 B.n558 B.n557 585
R472 B.n557 B.n57 585
R473 B.n556 B.n56 585
R474 B.n570 B.n56 585
R475 B.n555 B.n55 585
R476 B.n571 B.n55 585
R477 B.n554 B.n54 585
R478 B.n572 B.n54 585
R479 B.n553 B.n552 585
R480 B.n552 B.n53 585
R481 B.n551 B.n49 585
R482 B.n578 B.n49 585
R483 B.n550 B.n48 585
R484 B.n579 B.n48 585
R485 B.n549 B.n47 585
R486 B.n580 B.n47 585
R487 B.n548 B.n547 585
R488 B.n547 B.n43 585
R489 B.n546 B.n42 585
R490 B.n586 B.n42 585
R491 B.n545 B.n41 585
R492 B.n587 B.n41 585
R493 B.n544 B.n40 585
R494 B.n588 B.n40 585
R495 B.n543 B.n542 585
R496 B.n542 B.n36 585
R497 B.n541 B.n35 585
R498 B.n594 B.n35 585
R499 B.n540 B.n34 585
R500 B.n595 B.n34 585
R501 B.n539 B.n33 585
R502 B.n596 B.n33 585
R503 B.n538 B.n537 585
R504 B.n537 B.n29 585
R505 B.n536 B.n28 585
R506 B.n602 B.n28 585
R507 B.n535 B.n27 585
R508 B.n603 B.n27 585
R509 B.n534 B.n26 585
R510 B.n604 B.n26 585
R511 B.n533 B.n532 585
R512 B.n532 B.n22 585
R513 B.n531 B.n21 585
R514 B.n610 B.n21 585
R515 B.n530 B.n20 585
R516 B.n611 B.n20 585
R517 B.n529 B.n19 585
R518 B.n612 B.n19 585
R519 B.n528 B.n527 585
R520 B.n527 B.n15 585
R521 B.n526 B.n14 585
R522 B.n618 B.n14 585
R523 B.n525 B.n13 585
R524 B.n619 B.n13 585
R525 B.n524 B.n12 585
R526 B.n620 B.n12 585
R527 B.n523 B.n522 585
R528 B.n522 B.n521 585
R529 B.n520 B.n519 585
R530 B.n520 B.n8 585
R531 B.n518 B.n7 585
R532 B.n627 B.n7 585
R533 B.n517 B.n6 585
R534 B.n628 B.n6 585
R535 B.n516 B.n5 585
R536 B.n629 B.n5 585
R537 B.n515 B.n514 585
R538 B.n514 B.n4 585
R539 B.n513 B.n208 585
R540 B.n513 B.n512 585
R541 B.n503 B.n209 585
R542 B.n210 B.n209 585
R543 B.n505 B.n504 585
R544 B.n506 B.n505 585
R545 B.n502 B.n215 585
R546 B.n215 B.n214 585
R547 B.n501 B.n500 585
R548 B.n500 B.n499 585
R549 B.n217 B.n216 585
R550 B.n218 B.n217 585
R551 B.n492 B.n491 585
R552 B.n493 B.n492 585
R553 B.n490 B.n223 585
R554 B.n223 B.n222 585
R555 B.n489 B.n488 585
R556 B.n488 B.n487 585
R557 B.n225 B.n224 585
R558 B.n226 B.n225 585
R559 B.n480 B.n479 585
R560 B.n481 B.n480 585
R561 B.n478 B.n231 585
R562 B.n231 B.n230 585
R563 B.n477 B.n476 585
R564 B.n476 B.n475 585
R565 B.n233 B.n232 585
R566 B.n234 B.n233 585
R567 B.n468 B.n467 585
R568 B.n469 B.n468 585
R569 B.n466 B.n239 585
R570 B.n239 B.n238 585
R571 B.n465 B.n464 585
R572 B.n464 B.n463 585
R573 B.n241 B.n240 585
R574 B.n242 B.n241 585
R575 B.n456 B.n455 585
R576 B.n457 B.n456 585
R577 B.n454 B.n247 585
R578 B.n247 B.n246 585
R579 B.n453 B.n452 585
R580 B.n452 B.n451 585
R581 B.n249 B.n248 585
R582 B.n250 B.n249 585
R583 B.n444 B.n443 585
R584 B.n445 B.n444 585
R585 B.n442 B.n255 585
R586 B.n255 B.n254 585
R587 B.n441 B.n440 585
R588 B.n440 B.n439 585
R589 B.n257 B.n256 585
R590 B.n432 B.n257 585
R591 B.n431 B.n430 585
R592 B.n433 B.n431 585
R593 B.n429 B.n262 585
R594 B.n262 B.n261 585
R595 B.n428 B.n427 585
R596 B.n427 B.n426 585
R597 B.n264 B.n263 585
R598 B.n265 B.n264 585
R599 B.n419 B.n418 585
R600 B.n420 B.n419 585
R601 B.n268 B.n267 585
R602 B.n303 B.n301 585
R603 B.n304 B.n300 585
R604 B.n304 B.n269 585
R605 B.n307 B.n306 585
R606 B.n308 B.n299 585
R607 B.n310 B.n309 585
R608 B.n312 B.n298 585
R609 B.n315 B.n314 585
R610 B.n316 B.n297 585
R611 B.n318 B.n317 585
R612 B.n320 B.n296 585
R613 B.n323 B.n322 585
R614 B.n324 B.n295 585
R615 B.n326 B.n325 585
R616 B.n328 B.n294 585
R617 B.n331 B.n330 585
R618 B.n332 B.n293 585
R619 B.n334 B.n333 585
R620 B.n336 B.n292 585
R621 B.n339 B.n338 585
R622 B.n340 B.n291 585
R623 B.n342 B.n341 585
R624 B.n344 B.n290 585
R625 B.n347 B.n346 585
R626 B.n349 B.n287 585
R627 B.n351 B.n350 585
R628 B.n353 B.n286 585
R629 B.n356 B.n355 585
R630 B.n357 B.n285 585
R631 B.n359 B.n358 585
R632 B.n361 B.n284 585
R633 B.n364 B.n363 585
R634 B.n365 B.n283 585
R635 B.n370 B.n369 585
R636 B.n372 B.n282 585
R637 B.n375 B.n374 585
R638 B.n376 B.n281 585
R639 B.n378 B.n377 585
R640 B.n380 B.n280 585
R641 B.n383 B.n382 585
R642 B.n384 B.n279 585
R643 B.n386 B.n385 585
R644 B.n388 B.n278 585
R645 B.n391 B.n390 585
R646 B.n392 B.n277 585
R647 B.n394 B.n393 585
R648 B.n396 B.n276 585
R649 B.n399 B.n398 585
R650 B.n400 B.n275 585
R651 B.n402 B.n401 585
R652 B.n404 B.n274 585
R653 B.n407 B.n406 585
R654 B.n408 B.n273 585
R655 B.n410 B.n409 585
R656 B.n412 B.n272 585
R657 B.n413 B.n271 585
R658 B.n416 B.n415 585
R659 B.n417 B.n270 585
R660 B.n270 B.n269 585
R661 B.n422 B.n421 585
R662 B.n421 B.n420 585
R663 B.n423 B.n266 585
R664 B.n266 B.n265 585
R665 B.n425 B.n424 585
R666 B.n426 B.n425 585
R667 B.n260 B.n259 585
R668 B.n261 B.n260 585
R669 B.n435 B.n434 585
R670 B.n434 B.n433 585
R671 B.n436 B.n258 585
R672 B.n432 B.n258 585
R673 B.n438 B.n437 585
R674 B.n439 B.n438 585
R675 B.n253 B.n252 585
R676 B.n254 B.n253 585
R677 B.n447 B.n446 585
R678 B.n446 B.n445 585
R679 B.n448 B.n251 585
R680 B.n251 B.n250 585
R681 B.n450 B.n449 585
R682 B.n451 B.n450 585
R683 B.n245 B.n244 585
R684 B.n246 B.n245 585
R685 B.n459 B.n458 585
R686 B.n458 B.n457 585
R687 B.n460 B.n243 585
R688 B.n243 B.n242 585
R689 B.n462 B.n461 585
R690 B.n463 B.n462 585
R691 B.n237 B.n236 585
R692 B.n238 B.n237 585
R693 B.n471 B.n470 585
R694 B.n470 B.n469 585
R695 B.n472 B.n235 585
R696 B.n235 B.n234 585
R697 B.n474 B.n473 585
R698 B.n475 B.n474 585
R699 B.n229 B.n228 585
R700 B.n230 B.n229 585
R701 B.n483 B.n482 585
R702 B.n482 B.n481 585
R703 B.n484 B.n227 585
R704 B.n227 B.n226 585
R705 B.n486 B.n485 585
R706 B.n487 B.n486 585
R707 B.n221 B.n220 585
R708 B.n222 B.n221 585
R709 B.n495 B.n494 585
R710 B.n494 B.n493 585
R711 B.n496 B.n219 585
R712 B.n219 B.n218 585
R713 B.n498 B.n497 585
R714 B.n499 B.n498 585
R715 B.n213 B.n212 585
R716 B.n214 B.n213 585
R717 B.n508 B.n507 585
R718 B.n507 B.n506 585
R719 B.n509 B.n211 585
R720 B.n211 B.n210 585
R721 B.n511 B.n510 585
R722 B.n512 B.n511 585
R723 B.n3 B.n0 585
R724 B.n4 B.n3 585
R725 B.n626 B.n1 585
R726 B.n627 B.n626 585
R727 B.n625 B.n624 585
R728 B.n625 B.n8 585
R729 B.n623 B.n9 585
R730 B.n521 B.n9 585
R731 B.n622 B.n621 585
R732 B.n621 B.n620 585
R733 B.n11 B.n10 585
R734 B.n619 B.n11 585
R735 B.n617 B.n616 585
R736 B.n618 B.n617 585
R737 B.n615 B.n16 585
R738 B.n16 B.n15 585
R739 B.n614 B.n613 585
R740 B.n613 B.n612 585
R741 B.n18 B.n17 585
R742 B.n611 B.n18 585
R743 B.n609 B.n608 585
R744 B.n610 B.n609 585
R745 B.n607 B.n23 585
R746 B.n23 B.n22 585
R747 B.n606 B.n605 585
R748 B.n605 B.n604 585
R749 B.n25 B.n24 585
R750 B.n603 B.n25 585
R751 B.n601 B.n600 585
R752 B.n602 B.n601 585
R753 B.n599 B.n30 585
R754 B.n30 B.n29 585
R755 B.n598 B.n597 585
R756 B.n597 B.n596 585
R757 B.n32 B.n31 585
R758 B.n595 B.n32 585
R759 B.n593 B.n592 585
R760 B.n594 B.n593 585
R761 B.n591 B.n37 585
R762 B.n37 B.n36 585
R763 B.n590 B.n589 585
R764 B.n589 B.n588 585
R765 B.n39 B.n38 585
R766 B.n587 B.n39 585
R767 B.n585 B.n584 585
R768 B.n586 B.n585 585
R769 B.n583 B.n44 585
R770 B.n44 B.n43 585
R771 B.n582 B.n581 585
R772 B.n581 B.n580 585
R773 B.n46 B.n45 585
R774 B.n579 B.n46 585
R775 B.n577 B.n576 585
R776 B.n578 B.n577 585
R777 B.n575 B.n50 585
R778 B.n53 B.n50 585
R779 B.n574 B.n573 585
R780 B.n573 B.n572 585
R781 B.n52 B.n51 585
R782 B.n571 B.n52 585
R783 B.n569 B.n568 585
R784 B.n570 B.n569 585
R785 B.n567 B.n58 585
R786 B.n58 B.n57 585
R787 B.n566 B.n565 585
R788 B.n565 B.n564 585
R789 B.n630 B.n629 585
R790 B.n628 B.n2 585
R791 B.n565 B.n60 458.866
R792 B.n561 B.n61 458.866
R793 B.n419 B.n270 458.866
R794 B.n421 B.n268 458.866
R795 B.n94 B.t14 341.199
R796 B.n91 B.t18 341.199
R797 B.n366 B.t21 341.199
R798 B.n288 B.t10 341.199
R799 B.n563 B.n562 256.663
R800 B.n563 B.n89 256.663
R801 B.n563 B.n88 256.663
R802 B.n563 B.n87 256.663
R803 B.n563 B.n86 256.663
R804 B.n563 B.n85 256.663
R805 B.n563 B.n84 256.663
R806 B.n563 B.n83 256.663
R807 B.n563 B.n82 256.663
R808 B.n563 B.n81 256.663
R809 B.n563 B.n80 256.663
R810 B.n563 B.n79 256.663
R811 B.n563 B.n78 256.663
R812 B.n563 B.n77 256.663
R813 B.n563 B.n76 256.663
R814 B.n563 B.n75 256.663
R815 B.n563 B.n74 256.663
R816 B.n563 B.n73 256.663
R817 B.n563 B.n72 256.663
R818 B.n563 B.n71 256.663
R819 B.n563 B.n70 256.663
R820 B.n563 B.n69 256.663
R821 B.n563 B.n68 256.663
R822 B.n563 B.n67 256.663
R823 B.n563 B.n66 256.663
R824 B.n563 B.n65 256.663
R825 B.n563 B.n64 256.663
R826 B.n563 B.n63 256.663
R827 B.n563 B.n62 256.663
R828 B.n302 B.n269 256.663
R829 B.n305 B.n269 256.663
R830 B.n311 B.n269 256.663
R831 B.n313 B.n269 256.663
R832 B.n319 B.n269 256.663
R833 B.n321 B.n269 256.663
R834 B.n327 B.n269 256.663
R835 B.n329 B.n269 256.663
R836 B.n335 B.n269 256.663
R837 B.n337 B.n269 256.663
R838 B.n343 B.n269 256.663
R839 B.n345 B.n269 256.663
R840 B.n352 B.n269 256.663
R841 B.n354 B.n269 256.663
R842 B.n360 B.n269 256.663
R843 B.n362 B.n269 256.663
R844 B.n371 B.n269 256.663
R845 B.n373 B.n269 256.663
R846 B.n379 B.n269 256.663
R847 B.n381 B.n269 256.663
R848 B.n387 B.n269 256.663
R849 B.n389 B.n269 256.663
R850 B.n395 B.n269 256.663
R851 B.n397 B.n269 256.663
R852 B.n403 B.n269 256.663
R853 B.n405 B.n269 256.663
R854 B.n411 B.n269 256.663
R855 B.n414 B.n269 256.663
R856 B.n632 B.n631 256.663
R857 B.n91 B.t19 205.945
R858 B.n366 B.t23 205.945
R859 B.n94 B.t16 205.945
R860 B.n288 B.t13 205.945
R861 B.n92 B.t20 179.18
R862 B.n367 B.t22 179.18
R863 B.n95 B.t17 179.18
R864 B.n289 B.t12 179.18
R865 B.n99 B.n98 163.367
R866 B.n103 B.n102 163.367
R867 B.n107 B.n106 163.367
R868 B.n111 B.n110 163.367
R869 B.n115 B.n114 163.367
R870 B.n119 B.n118 163.367
R871 B.n123 B.n122 163.367
R872 B.n127 B.n126 163.367
R873 B.n131 B.n130 163.367
R874 B.n135 B.n134 163.367
R875 B.n139 B.n138 163.367
R876 B.n143 B.n142 163.367
R877 B.n147 B.n146 163.367
R878 B.n151 B.n150 163.367
R879 B.n155 B.n154 163.367
R880 B.n159 B.n158 163.367
R881 B.n163 B.n162 163.367
R882 B.n167 B.n166 163.367
R883 B.n171 B.n170 163.367
R884 B.n175 B.n174 163.367
R885 B.n179 B.n178 163.367
R886 B.n183 B.n182 163.367
R887 B.n187 B.n186 163.367
R888 B.n191 B.n190 163.367
R889 B.n195 B.n194 163.367
R890 B.n199 B.n198 163.367
R891 B.n203 B.n202 163.367
R892 B.n205 B.n90 163.367
R893 B.n419 B.n264 163.367
R894 B.n427 B.n264 163.367
R895 B.n427 B.n262 163.367
R896 B.n431 B.n262 163.367
R897 B.n431 B.n257 163.367
R898 B.n440 B.n257 163.367
R899 B.n440 B.n255 163.367
R900 B.n444 B.n255 163.367
R901 B.n444 B.n249 163.367
R902 B.n452 B.n249 163.367
R903 B.n452 B.n247 163.367
R904 B.n456 B.n247 163.367
R905 B.n456 B.n241 163.367
R906 B.n464 B.n241 163.367
R907 B.n464 B.n239 163.367
R908 B.n468 B.n239 163.367
R909 B.n468 B.n233 163.367
R910 B.n476 B.n233 163.367
R911 B.n476 B.n231 163.367
R912 B.n480 B.n231 163.367
R913 B.n480 B.n225 163.367
R914 B.n488 B.n225 163.367
R915 B.n488 B.n223 163.367
R916 B.n492 B.n223 163.367
R917 B.n492 B.n217 163.367
R918 B.n500 B.n217 163.367
R919 B.n500 B.n215 163.367
R920 B.n505 B.n215 163.367
R921 B.n505 B.n209 163.367
R922 B.n513 B.n209 163.367
R923 B.n514 B.n513 163.367
R924 B.n514 B.n5 163.367
R925 B.n6 B.n5 163.367
R926 B.n7 B.n6 163.367
R927 B.n520 B.n7 163.367
R928 B.n522 B.n520 163.367
R929 B.n522 B.n12 163.367
R930 B.n13 B.n12 163.367
R931 B.n14 B.n13 163.367
R932 B.n527 B.n14 163.367
R933 B.n527 B.n19 163.367
R934 B.n20 B.n19 163.367
R935 B.n21 B.n20 163.367
R936 B.n532 B.n21 163.367
R937 B.n532 B.n26 163.367
R938 B.n27 B.n26 163.367
R939 B.n28 B.n27 163.367
R940 B.n537 B.n28 163.367
R941 B.n537 B.n33 163.367
R942 B.n34 B.n33 163.367
R943 B.n35 B.n34 163.367
R944 B.n542 B.n35 163.367
R945 B.n542 B.n40 163.367
R946 B.n41 B.n40 163.367
R947 B.n42 B.n41 163.367
R948 B.n547 B.n42 163.367
R949 B.n547 B.n47 163.367
R950 B.n48 B.n47 163.367
R951 B.n49 B.n48 163.367
R952 B.n552 B.n49 163.367
R953 B.n552 B.n54 163.367
R954 B.n55 B.n54 163.367
R955 B.n56 B.n55 163.367
R956 B.n557 B.n56 163.367
R957 B.n557 B.n61 163.367
R958 B.n304 B.n303 163.367
R959 B.n306 B.n304 163.367
R960 B.n310 B.n299 163.367
R961 B.n314 B.n312 163.367
R962 B.n318 B.n297 163.367
R963 B.n322 B.n320 163.367
R964 B.n326 B.n295 163.367
R965 B.n330 B.n328 163.367
R966 B.n334 B.n293 163.367
R967 B.n338 B.n336 163.367
R968 B.n342 B.n291 163.367
R969 B.n346 B.n344 163.367
R970 B.n351 B.n287 163.367
R971 B.n355 B.n353 163.367
R972 B.n359 B.n285 163.367
R973 B.n363 B.n361 163.367
R974 B.n370 B.n283 163.367
R975 B.n374 B.n372 163.367
R976 B.n378 B.n281 163.367
R977 B.n382 B.n380 163.367
R978 B.n386 B.n279 163.367
R979 B.n390 B.n388 163.367
R980 B.n394 B.n277 163.367
R981 B.n398 B.n396 163.367
R982 B.n402 B.n275 163.367
R983 B.n406 B.n404 163.367
R984 B.n410 B.n273 163.367
R985 B.n413 B.n412 163.367
R986 B.n415 B.n270 163.367
R987 B.n421 B.n266 163.367
R988 B.n425 B.n266 163.367
R989 B.n425 B.n260 163.367
R990 B.n434 B.n260 163.367
R991 B.n434 B.n258 163.367
R992 B.n438 B.n258 163.367
R993 B.n438 B.n253 163.367
R994 B.n446 B.n253 163.367
R995 B.n446 B.n251 163.367
R996 B.n450 B.n251 163.367
R997 B.n450 B.n245 163.367
R998 B.n458 B.n245 163.367
R999 B.n458 B.n243 163.367
R1000 B.n462 B.n243 163.367
R1001 B.n462 B.n237 163.367
R1002 B.n470 B.n237 163.367
R1003 B.n470 B.n235 163.367
R1004 B.n474 B.n235 163.367
R1005 B.n474 B.n229 163.367
R1006 B.n482 B.n229 163.367
R1007 B.n482 B.n227 163.367
R1008 B.n486 B.n227 163.367
R1009 B.n486 B.n221 163.367
R1010 B.n494 B.n221 163.367
R1011 B.n494 B.n219 163.367
R1012 B.n498 B.n219 163.367
R1013 B.n498 B.n213 163.367
R1014 B.n507 B.n213 163.367
R1015 B.n507 B.n211 163.367
R1016 B.n511 B.n211 163.367
R1017 B.n511 B.n3 163.367
R1018 B.n630 B.n3 163.367
R1019 B.n626 B.n2 163.367
R1020 B.n626 B.n625 163.367
R1021 B.n625 B.n9 163.367
R1022 B.n621 B.n9 163.367
R1023 B.n621 B.n11 163.367
R1024 B.n617 B.n11 163.367
R1025 B.n617 B.n16 163.367
R1026 B.n613 B.n16 163.367
R1027 B.n613 B.n18 163.367
R1028 B.n609 B.n18 163.367
R1029 B.n609 B.n23 163.367
R1030 B.n605 B.n23 163.367
R1031 B.n605 B.n25 163.367
R1032 B.n601 B.n25 163.367
R1033 B.n601 B.n30 163.367
R1034 B.n597 B.n30 163.367
R1035 B.n597 B.n32 163.367
R1036 B.n593 B.n32 163.367
R1037 B.n593 B.n37 163.367
R1038 B.n589 B.n37 163.367
R1039 B.n589 B.n39 163.367
R1040 B.n585 B.n39 163.367
R1041 B.n585 B.n44 163.367
R1042 B.n581 B.n44 163.367
R1043 B.n581 B.n46 163.367
R1044 B.n577 B.n46 163.367
R1045 B.n577 B.n50 163.367
R1046 B.n573 B.n50 163.367
R1047 B.n573 B.n52 163.367
R1048 B.n569 B.n52 163.367
R1049 B.n569 B.n58 163.367
R1050 B.n565 B.n58 163.367
R1051 B.n420 B.n269 117.945
R1052 B.n564 B.n563 117.945
R1053 B.n62 B.n60 71.676
R1054 B.n99 B.n63 71.676
R1055 B.n103 B.n64 71.676
R1056 B.n107 B.n65 71.676
R1057 B.n111 B.n66 71.676
R1058 B.n115 B.n67 71.676
R1059 B.n119 B.n68 71.676
R1060 B.n123 B.n69 71.676
R1061 B.n127 B.n70 71.676
R1062 B.n131 B.n71 71.676
R1063 B.n135 B.n72 71.676
R1064 B.n139 B.n73 71.676
R1065 B.n143 B.n74 71.676
R1066 B.n147 B.n75 71.676
R1067 B.n151 B.n76 71.676
R1068 B.n155 B.n77 71.676
R1069 B.n159 B.n78 71.676
R1070 B.n163 B.n79 71.676
R1071 B.n167 B.n80 71.676
R1072 B.n171 B.n81 71.676
R1073 B.n175 B.n82 71.676
R1074 B.n179 B.n83 71.676
R1075 B.n183 B.n84 71.676
R1076 B.n187 B.n85 71.676
R1077 B.n191 B.n86 71.676
R1078 B.n195 B.n87 71.676
R1079 B.n199 B.n88 71.676
R1080 B.n203 B.n89 71.676
R1081 B.n562 B.n90 71.676
R1082 B.n562 B.n561 71.676
R1083 B.n205 B.n89 71.676
R1084 B.n202 B.n88 71.676
R1085 B.n198 B.n87 71.676
R1086 B.n194 B.n86 71.676
R1087 B.n190 B.n85 71.676
R1088 B.n186 B.n84 71.676
R1089 B.n182 B.n83 71.676
R1090 B.n178 B.n82 71.676
R1091 B.n174 B.n81 71.676
R1092 B.n170 B.n80 71.676
R1093 B.n166 B.n79 71.676
R1094 B.n162 B.n78 71.676
R1095 B.n158 B.n77 71.676
R1096 B.n154 B.n76 71.676
R1097 B.n150 B.n75 71.676
R1098 B.n146 B.n74 71.676
R1099 B.n142 B.n73 71.676
R1100 B.n138 B.n72 71.676
R1101 B.n134 B.n71 71.676
R1102 B.n130 B.n70 71.676
R1103 B.n126 B.n69 71.676
R1104 B.n122 B.n68 71.676
R1105 B.n118 B.n67 71.676
R1106 B.n114 B.n66 71.676
R1107 B.n110 B.n65 71.676
R1108 B.n106 B.n64 71.676
R1109 B.n102 B.n63 71.676
R1110 B.n98 B.n62 71.676
R1111 B.n302 B.n268 71.676
R1112 B.n306 B.n305 71.676
R1113 B.n311 B.n310 71.676
R1114 B.n314 B.n313 71.676
R1115 B.n319 B.n318 71.676
R1116 B.n322 B.n321 71.676
R1117 B.n327 B.n326 71.676
R1118 B.n330 B.n329 71.676
R1119 B.n335 B.n334 71.676
R1120 B.n338 B.n337 71.676
R1121 B.n343 B.n342 71.676
R1122 B.n346 B.n345 71.676
R1123 B.n352 B.n351 71.676
R1124 B.n355 B.n354 71.676
R1125 B.n360 B.n359 71.676
R1126 B.n363 B.n362 71.676
R1127 B.n371 B.n370 71.676
R1128 B.n374 B.n373 71.676
R1129 B.n379 B.n378 71.676
R1130 B.n382 B.n381 71.676
R1131 B.n387 B.n386 71.676
R1132 B.n390 B.n389 71.676
R1133 B.n395 B.n394 71.676
R1134 B.n398 B.n397 71.676
R1135 B.n403 B.n402 71.676
R1136 B.n406 B.n405 71.676
R1137 B.n411 B.n410 71.676
R1138 B.n414 B.n413 71.676
R1139 B.n303 B.n302 71.676
R1140 B.n305 B.n299 71.676
R1141 B.n312 B.n311 71.676
R1142 B.n313 B.n297 71.676
R1143 B.n320 B.n319 71.676
R1144 B.n321 B.n295 71.676
R1145 B.n328 B.n327 71.676
R1146 B.n329 B.n293 71.676
R1147 B.n336 B.n335 71.676
R1148 B.n337 B.n291 71.676
R1149 B.n344 B.n343 71.676
R1150 B.n345 B.n287 71.676
R1151 B.n353 B.n352 71.676
R1152 B.n354 B.n285 71.676
R1153 B.n361 B.n360 71.676
R1154 B.n362 B.n283 71.676
R1155 B.n372 B.n371 71.676
R1156 B.n373 B.n281 71.676
R1157 B.n380 B.n379 71.676
R1158 B.n381 B.n279 71.676
R1159 B.n388 B.n387 71.676
R1160 B.n389 B.n277 71.676
R1161 B.n396 B.n395 71.676
R1162 B.n397 B.n275 71.676
R1163 B.n404 B.n403 71.676
R1164 B.n405 B.n273 71.676
R1165 B.n412 B.n411 71.676
R1166 B.n415 B.n414 71.676
R1167 B.n631 B.n630 71.676
R1168 B.n631 B.n2 71.676
R1169 B.n420 B.n265 66.2832
R1170 B.n426 B.n265 66.2832
R1171 B.n426 B.n261 66.2832
R1172 B.n433 B.n261 66.2832
R1173 B.n433 B.n432 66.2832
R1174 B.n439 B.n254 66.2832
R1175 B.n445 B.n254 66.2832
R1176 B.n445 B.n250 66.2832
R1177 B.n451 B.n250 66.2832
R1178 B.n451 B.n246 66.2832
R1179 B.n457 B.n246 66.2832
R1180 B.n463 B.n242 66.2832
R1181 B.n463 B.n238 66.2832
R1182 B.n469 B.n238 66.2832
R1183 B.n475 B.n234 66.2832
R1184 B.n475 B.n230 66.2832
R1185 B.n481 B.n230 66.2832
R1186 B.n487 B.n226 66.2832
R1187 B.n487 B.n222 66.2832
R1188 B.n493 B.n222 66.2832
R1189 B.n499 B.n218 66.2832
R1190 B.n499 B.n214 66.2832
R1191 B.n506 B.n214 66.2832
R1192 B.n512 B.n210 66.2832
R1193 B.n512 B.n4 66.2832
R1194 B.n629 B.n4 66.2832
R1195 B.n629 B.n628 66.2832
R1196 B.n628 B.n627 66.2832
R1197 B.n627 B.n8 66.2832
R1198 B.n521 B.n8 66.2832
R1199 B.n620 B.n619 66.2832
R1200 B.n619 B.n618 66.2832
R1201 B.n618 B.n15 66.2832
R1202 B.n612 B.n611 66.2832
R1203 B.n611 B.n610 66.2832
R1204 B.n610 B.n22 66.2832
R1205 B.n604 B.n603 66.2832
R1206 B.n603 B.n602 66.2832
R1207 B.n602 B.n29 66.2832
R1208 B.n596 B.n595 66.2832
R1209 B.n595 B.n594 66.2832
R1210 B.n594 B.n36 66.2832
R1211 B.n588 B.n587 66.2832
R1212 B.n587 B.n586 66.2832
R1213 B.n586 B.n43 66.2832
R1214 B.n580 B.n43 66.2832
R1215 B.n580 B.n579 66.2832
R1216 B.n579 B.n578 66.2832
R1217 B.n572 B.n53 66.2832
R1218 B.n572 B.n571 66.2832
R1219 B.n571 B.n570 66.2832
R1220 B.n570 B.n57 66.2832
R1221 B.n564 B.n57 66.2832
R1222 B.n96 B.n95 59.5399
R1223 B.n93 B.n92 59.5399
R1224 B.n368 B.n367 59.5399
R1225 B.n348 B.n289 59.5399
R1226 B.n506 B.t2 57.5105
R1227 B.n620 B.t0 57.5105
R1228 B.n493 B.t9 53.6115
R1229 B.n612 B.t8 53.6115
R1230 B.n481 B.t5 49.7125
R1231 B.n604 B.t6 49.7125
R1232 B.n469 B.t4 45.8135
R1233 B.n596 B.t7 45.8135
R1234 B.n439 B.t11 41.9145
R1235 B.n457 B.t3 41.9145
R1236 B.n588 B.t1 41.9145
R1237 B.n578 B.t15 41.9145
R1238 B.n560 B.n559 29.8151
R1239 B.n422 B.n267 29.8151
R1240 B.n418 B.n417 29.8151
R1241 B.n566 B.n59 29.8151
R1242 B.n95 B.n94 26.7641
R1243 B.n92 B.n91 26.7641
R1244 B.n367 B.n366 26.7641
R1245 B.n289 B.n288 26.7641
R1246 B.n432 B.t11 24.3691
R1247 B.t3 B.n242 24.3691
R1248 B.t1 B.n36 24.3691
R1249 B.n53 B.t15 24.3691
R1250 B.t4 B.n234 20.4702
R1251 B.t7 B.n29 20.4702
R1252 B B.n632 18.0485
R1253 B.t5 B.n226 16.5712
R1254 B.t6 B.n22 16.5712
R1255 B.t9 B.n218 12.6722
R1256 B.t8 B.n15 12.6722
R1257 B.n423 B.n422 10.6151
R1258 B.n424 B.n423 10.6151
R1259 B.n424 B.n259 10.6151
R1260 B.n435 B.n259 10.6151
R1261 B.n436 B.n435 10.6151
R1262 B.n437 B.n436 10.6151
R1263 B.n437 B.n252 10.6151
R1264 B.n447 B.n252 10.6151
R1265 B.n448 B.n447 10.6151
R1266 B.n449 B.n448 10.6151
R1267 B.n449 B.n244 10.6151
R1268 B.n459 B.n244 10.6151
R1269 B.n460 B.n459 10.6151
R1270 B.n461 B.n460 10.6151
R1271 B.n461 B.n236 10.6151
R1272 B.n471 B.n236 10.6151
R1273 B.n472 B.n471 10.6151
R1274 B.n473 B.n472 10.6151
R1275 B.n473 B.n228 10.6151
R1276 B.n483 B.n228 10.6151
R1277 B.n484 B.n483 10.6151
R1278 B.n485 B.n484 10.6151
R1279 B.n485 B.n220 10.6151
R1280 B.n495 B.n220 10.6151
R1281 B.n496 B.n495 10.6151
R1282 B.n497 B.n496 10.6151
R1283 B.n497 B.n212 10.6151
R1284 B.n508 B.n212 10.6151
R1285 B.n509 B.n508 10.6151
R1286 B.n510 B.n509 10.6151
R1287 B.n510 B.n0 10.6151
R1288 B.n301 B.n267 10.6151
R1289 B.n301 B.n300 10.6151
R1290 B.n307 B.n300 10.6151
R1291 B.n308 B.n307 10.6151
R1292 B.n309 B.n308 10.6151
R1293 B.n309 B.n298 10.6151
R1294 B.n315 B.n298 10.6151
R1295 B.n316 B.n315 10.6151
R1296 B.n317 B.n316 10.6151
R1297 B.n317 B.n296 10.6151
R1298 B.n323 B.n296 10.6151
R1299 B.n324 B.n323 10.6151
R1300 B.n325 B.n324 10.6151
R1301 B.n325 B.n294 10.6151
R1302 B.n331 B.n294 10.6151
R1303 B.n332 B.n331 10.6151
R1304 B.n333 B.n332 10.6151
R1305 B.n333 B.n292 10.6151
R1306 B.n339 B.n292 10.6151
R1307 B.n340 B.n339 10.6151
R1308 B.n341 B.n340 10.6151
R1309 B.n341 B.n290 10.6151
R1310 B.n347 B.n290 10.6151
R1311 B.n350 B.n349 10.6151
R1312 B.n350 B.n286 10.6151
R1313 B.n356 B.n286 10.6151
R1314 B.n357 B.n356 10.6151
R1315 B.n358 B.n357 10.6151
R1316 B.n358 B.n284 10.6151
R1317 B.n364 B.n284 10.6151
R1318 B.n365 B.n364 10.6151
R1319 B.n369 B.n365 10.6151
R1320 B.n375 B.n282 10.6151
R1321 B.n376 B.n375 10.6151
R1322 B.n377 B.n376 10.6151
R1323 B.n377 B.n280 10.6151
R1324 B.n383 B.n280 10.6151
R1325 B.n384 B.n383 10.6151
R1326 B.n385 B.n384 10.6151
R1327 B.n385 B.n278 10.6151
R1328 B.n391 B.n278 10.6151
R1329 B.n392 B.n391 10.6151
R1330 B.n393 B.n392 10.6151
R1331 B.n393 B.n276 10.6151
R1332 B.n399 B.n276 10.6151
R1333 B.n400 B.n399 10.6151
R1334 B.n401 B.n400 10.6151
R1335 B.n401 B.n274 10.6151
R1336 B.n407 B.n274 10.6151
R1337 B.n408 B.n407 10.6151
R1338 B.n409 B.n408 10.6151
R1339 B.n409 B.n272 10.6151
R1340 B.n272 B.n271 10.6151
R1341 B.n416 B.n271 10.6151
R1342 B.n417 B.n416 10.6151
R1343 B.n418 B.n263 10.6151
R1344 B.n428 B.n263 10.6151
R1345 B.n429 B.n428 10.6151
R1346 B.n430 B.n429 10.6151
R1347 B.n430 B.n256 10.6151
R1348 B.n441 B.n256 10.6151
R1349 B.n442 B.n441 10.6151
R1350 B.n443 B.n442 10.6151
R1351 B.n443 B.n248 10.6151
R1352 B.n453 B.n248 10.6151
R1353 B.n454 B.n453 10.6151
R1354 B.n455 B.n454 10.6151
R1355 B.n455 B.n240 10.6151
R1356 B.n465 B.n240 10.6151
R1357 B.n466 B.n465 10.6151
R1358 B.n467 B.n466 10.6151
R1359 B.n467 B.n232 10.6151
R1360 B.n477 B.n232 10.6151
R1361 B.n478 B.n477 10.6151
R1362 B.n479 B.n478 10.6151
R1363 B.n479 B.n224 10.6151
R1364 B.n489 B.n224 10.6151
R1365 B.n490 B.n489 10.6151
R1366 B.n491 B.n490 10.6151
R1367 B.n491 B.n216 10.6151
R1368 B.n501 B.n216 10.6151
R1369 B.n502 B.n501 10.6151
R1370 B.n504 B.n502 10.6151
R1371 B.n504 B.n503 10.6151
R1372 B.n503 B.n208 10.6151
R1373 B.n515 B.n208 10.6151
R1374 B.n516 B.n515 10.6151
R1375 B.n517 B.n516 10.6151
R1376 B.n518 B.n517 10.6151
R1377 B.n519 B.n518 10.6151
R1378 B.n523 B.n519 10.6151
R1379 B.n524 B.n523 10.6151
R1380 B.n525 B.n524 10.6151
R1381 B.n526 B.n525 10.6151
R1382 B.n528 B.n526 10.6151
R1383 B.n529 B.n528 10.6151
R1384 B.n530 B.n529 10.6151
R1385 B.n531 B.n530 10.6151
R1386 B.n533 B.n531 10.6151
R1387 B.n534 B.n533 10.6151
R1388 B.n535 B.n534 10.6151
R1389 B.n536 B.n535 10.6151
R1390 B.n538 B.n536 10.6151
R1391 B.n539 B.n538 10.6151
R1392 B.n540 B.n539 10.6151
R1393 B.n541 B.n540 10.6151
R1394 B.n543 B.n541 10.6151
R1395 B.n544 B.n543 10.6151
R1396 B.n545 B.n544 10.6151
R1397 B.n546 B.n545 10.6151
R1398 B.n548 B.n546 10.6151
R1399 B.n549 B.n548 10.6151
R1400 B.n550 B.n549 10.6151
R1401 B.n551 B.n550 10.6151
R1402 B.n553 B.n551 10.6151
R1403 B.n554 B.n553 10.6151
R1404 B.n555 B.n554 10.6151
R1405 B.n556 B.n555 10.6151
R1406 B.n558 B.n556 10.6151
R1407 B.n559 B.n558 10.6151
R1408 B.n624 B.n1 10.6151
R1409 B.n624 B.n623 10.6151
R1410 B.n623 B.n622 10.6151
R1411 B.n622 B.n10 10.6151
R1412 B.n616 B.n10 10.6151
R1413 B.n616 B.n615 10.6151
R1414 B.n615 B.n614 10.6151
R1415 B.n614 B.n17 10.6151
R1416 B.n608 B.n17 10.6151
R1417 B.n608 B.n607 10.6151
R1418 B.n607 B.n606 10.6151
R1419 B.n606 B.n24 10.6151
R1420 B.n600 B.n24 10.6151
R1421 B.n600 B.n599 10.6151
R1422 B.n599 B.n598 10.6151
R1423 B.n598 B.n31 10.6151
R1424 B.n592 B.n31 10.6151
R1425 B.n592 B.n591 10.6151
R1426 B.n591 B.n590 10.6151
R1427 B.n590 B.n38 10.6151
R1428 B.n584 B.n38 10.6151
R1429 B.n584 B.n583 10.6151
R1430 B.n583 B.n582 10.6151
R1431 B.n582 B.n45 10.6151
R1432 B.n576 B.n45 10.6151
R1433 B.n576 B.n575 10.6151
R1434 B.n575 B.n574 10.6151
R1435 B.n574 B.n51 10.6151
R1436 B.n568 B.n51 10.6151
R1437 B.n568 B.n567 10.6151
R1438 B.n567 B.n566 10.6151
R1439 B.n97 B.n59 10.6151
R1440 B.n100 B.n97 10.6151
R1441 B.n101 B.n100 10.6151
R1442 B.n104 B.n101 10.6151
R1443 B.n105 B.n104 10.6151
R1444 B.n108 B.n105 10.6151
R1445 B.n109 B.n108 10.6151
R1446 B.n112 B.n109 10.6151
R1447 B.n113 B.n112 10.6151
R1448 B.n116 B.n113 10.6151
R1449 B.n117 B.n116 10.6151
R1450 B.n120 B.n117 10.6151
R1451 B.n121 B.n120 10.6151
R1452 B.n124 B.n121 10.6151
R1453 B.n125 B.n124 10.6151
R1454 B.n128 B.n125 10.6151
R1455 B.n129 B.n128 10.6151
R1456 B.n132 B.n129 10.6151
R1457 B.n133 B.n132 10.6151
R1458 B.n136 B.n133 10.6151
R1459 B.n137 B.n136 10.6151
R1460 B.n140 B.n137 10.6151
R1461 B.n141 B.n140 10.6151
R1462 B.n145 B.n144 10.6151
R1463 B.n148 B.n145 10.6151
R1464 B.n149 B.n148 10.6151
R1465 B.n152 B.n149 10.6151
R1466 B.n153 B.n152 10.6151
R1467 B.n156 B.n153 10.6151
R1468 B.n157 B.n156 10.6151
R1469 B.n160 B.n157 10.6151
R1470 B.n161 B.n160 10.6151
R1471 B.n165 B.n164 10.6151
R1472 B.n168 B.n165 10.6151
R1473 B.n169 B.n168 10.6151
R1474 B.n172 B.n169 10.6151
R1475 B.n173 B.n172 10.6151
R1476 B.n176 B.n173 10.6151
R1477 B.n177 B.n176 10.6151
R1478 B.n180 B.n177 10.6151
R1479 B.n181 B.n180 10.6151
R1480 B.n184 B.n181 10.6151
R1481 B.n185 B.n184 10.6151
R1482 B.n188 B.n185 10.6151
R1483 B.n189 B.n188 10.6151
R1484 B.n192 B.n189 10.6151
R1485 B.n193 B.n192 10.6151
R1486 B.n196 B.n193 10.6151
R1487 B.n197 B.n196 10.6151
R1488 B.n200 B.n197 10.6151
R1489 B.n201 B.n200 10.6151
R1490 B.n204 B.n201 10.6151
R1491 B.n206 B.n204 10.6151
R1492 B.n207 B.n206 10.6151
R1493 B.n560 B.n207 10.6151
R1494 B.n348 B.n347 9.36635
R1495 B.n368 B.n282 9.36635
R1496 B.n141 B.n96 9.36635
R1497 B.n164 B.n93 9.36635
R1498 B.t2 B.n210 8.77321
R1499 B.n521 B.t0 8.77321
R1500 B.n632 B.n0 8.11757
R1501 B.n632 B.n1 8.11757
R1502 B.n349 B.n348 1.24928
R1503 B.n369 B.n368 1.24928
R1504 B.n144 B.n96 1.24928
R1505 B.n161 B.n93 1.24928
R1506 VN.n5 VN.t0 190.731
R1507 VN.n25 VN.t7 190.731
R1508 VN.n18 VN.t9 175.587
R1509 VN.n38 VN.t2 175.587
R1510 VN.n37 VN.n20 161.3
R1511 VN.n35 VN.n34 161.3
R1512 VN.n33 VN.n21 161.3
R1513 VN.n32 VN.n31 161.3
R1514 VN.n29 VN.n22 161.3
R1515 VN.n28 VN.n27 161.3
R1516 VN.n26 VN.n23 161.3
R1517 VN.n17 VN.n0 161.3
R1518 VN.n15 VN.n14 161.3
R1519 VN.n13 VN.n1 161.3
R1520 VN.n12 VN.n11 161.3
R1521 VN.n9 VN.n2 161.3
R1522 VN.n8 VN.n7 161.3
R1523 VN.n6 VN.n3 161.3
R1524 VN.n4 VN.t8 137.945
R1525 VN.n10 VN.t3 137.945
R1526 VN.n16 VN.t5 137.945
R1527 VN.n24 VN.t6 137.945
R1528 VN.n30 VN.t4 137.945
R1529 VN.n36 VN.t1 137.945
R1530 VN.n39 VN.n38 80.6037
R1531 VN.n19 VN.n18 80.6037
R1532 VN.n18 VN.n17 55.7853
R1533 VN.n38 VN.n37 55.7853
R1534 VN.n5 VN.n4 48.3043
R1535 VN.n25 VN.n24 48.3043
R1536 VN.n9 VN.n8 46.321
R1537 VN.n11 VN.n1 46.321
R1538 VN.n29 VN.n28 46.321
R1539 VN.n31 VN.n21 46.321
R1540 VN.n26 VN.n25 43.9769
R1541 VN.n6 VN.n5 43.9769
R1542 VN VN.n39 40.6733
R1543 VN.n8 VN.n3 34.6658
R1544 VN.n15 VN.n1 34.6658
R1545 VN.n28 VN.n23 34.6658
R1546 VN.n35 VN.n21 34.6658
R1547 VN.n17 VN.n16 18.1061
R1548 VN.n37 VN.n36 18.1061
R1549 VN.n10 VN.n9 12.234
R1550 VN.n11 VN.n10 12.234
R1551 VN.n31 VN.n30 12.234
R1552 VN.n30 VN.n29 12.234
R1553 VN.n4 VN.n3 6.36192
R1554 VN.n16 VN.n15 6.36192
R1555 VN.n24 VN.n23 6.36192
R1556 VN.n36 VN.n35 6.36192
R1557 VN.n39 VN.n20 0.285035
R1558 VN.n19 VN.n0 0.285035
R1559 VN.n34 VN.n20 0.189894
R1560 VN.n34 VN.n33 0.189894
R1561 VN.n33 VN.n32 0.189894
R1562 VN.n32 VN.n22 0.189894
R1563 VN.n27 VN.n22 0.189894
R1564 VN.n27 VN.n26 0.189894
R1565 VN.n7 VN.n6 0.189894
R1566 VN.n7 VN.n2 0.189894
R1567 VN.n12 VN.n2 0.189894
R1568 VN.n13 VN.n12 0.189894
R1569 VN.n14 VN.n13 0.189894
R1570 VN.n14 VN.n0 0.189894
R1571 VN VN.n19 0.146778
R1572 VDD2.n61 VDD2.n35 289.615
R1573 VDD2.n26 VDD2.n0 289.615
R1574 VDD2.n62 VDD2.n61 185
R1575 VDD2.n60 VDD2.n59 185
R1576 VDD2.n39 VDD2.n38 185
R1577 VDD2.n54 VDD2.n53 185
R1578 VDD2.n52 VDD2.n51 185
R1579 VDD2.n43 VDD2.n42 185
R1580 VDD2.n46 VDD2.n45 185
R1581 VDD2.n11 VDD2.n10 185
R1582 VDD2.n8 VDD2.n7 185
R1583 VDD2.n17 VDD2.n16 185
R1584 VDD2.n19 VDD2.n18 185
R1585 VDD2.n4 VDD2.n3 185
R1586 VDD2.n25 VDD2.n24 185
R1587 VDD2.n27 VDD2.n26 185
R1588 VDD2.t7 VDD2.n44 147.661
R1589 VDD2.t9 VDD2.n9 147.661
R1590 VDD2.n61 VDD2.n60 104.615
R1591 VDD2.n60 VDD2.n38 104.615
R1592 VDD2.n53 VDD2.n38 104.615
R1593 VDD2.n53 VDD2.n52 104.615
R1594 VDD2.n52 VDD2.n42 104.615
R1595 VDD2.n45 VDD2.n42 104.615
R1596 VDD2.n10 VDD2.n7 104.615
R1597 VDD2.n17 VDD2.n7 104.615
R1598 VDD2.n18 VDD2.n17 104.615
R1599 VDD2.n18 VDD2.n3 104.615
R1600 VDD2.n25 VDD2.n3 104.615
R1601 VDD2.n26 VDD2.n25 104.615
R1602 VDD2.n34 VDD2.n33 68.2215
R1603 VDD2 VDD2.n69 68.2186
R1604 VDD2.n68 VDD2.n67 67.3848
R1605 VDD2.n32 VDD2.n31 67.3846
R1606 VDD2.n45 VDD2.t7 52.3082
R1607 VDD2.n10 VDD2.t9 52.3082
R1608 VDD2.n32 VDD2.n30 50.2477
R1609 VDD2.n66 VDD2.n65 49.0581
R1610 VDD2.n66 VDD2.n34 34.5472
R1611 VDD2.n46 VDD2.n44 15.6674
R1612 VDD2.n11 VDD2.n9 15.6674
R1613 VDD2.n47 VDD2.n43 12.8005
R1614 VDD2.n12 VDD2.n8 12.8005
R1615 VDD2.n51 VDD2.n50 12.0247
R1616 VDD2.n16 VDD2.n15 12.0247
R1617 VDD2.n54 VDD2.n41 11.249
R1618 VDD2.n19 VDD2.n6 11.249
R1619 VDD2.n55 VDD2.n39 10.4732
R1620 VDD2.n20 VDD2.n4 10.4732
R1621 VDD2.n59 VDD2.n58 9.69747
R1622 VDD2.n24 VDD2.n23 9.69747
R1623 VDD2.n65 VDD2.n64 9.45567
R1624 VDD2.n30 VDD2.n29 9.45567
R1625 VDD2.n64 VDD2.n63 9.3005
R1626 VDD2.n37 VDD2.n36 9.3005
R1627 VDD2.n58 VDD2.n57 9.3005
R1628 VDD2.n56 VDD2.n55 9.3005
R1629 VDD2.n41 VDD2.n40 9.3005
R1630 VDD2.n50 VDD2.n49 9.3005
R1631 VDD2.n48 VDD2.n47 9.3005
R1632 VDD2.n29 VDD2.n28 9.3005
R1633 VDD2.n2 VDD2.n1 9.3005
R1634 VDD2.n23 VDD2.n22 9.3005
R1635 VDD2.n21 VDD2.n20 9.3005
R1636 VDD2.n6 VDD2.n5 9.3005
R1637 VDD2.n15 VDD2.n14 9.3005
R1638 VDD2.n13 VDD2.n12 9.3005
R1639 VDD2.n62 VDD2.n37 8.92171
R1640 VDD2.n27 VDD2.n2 8.92171
R1641 VDD2.n63 VDD2.n35 8.14595
R1642 VDD2.n28 VDD2.n0 8.14595
R1643 VDD2.n65 VDD2.n35 5.81868
R1644 VDD2.n30 VDD2.n0 5.81868
R1645 VDD2.n63 VDD2.n62 5.04292
R1646 VDD2.n28 VDD2.n27 5.04292
R1647 VDD2.n48 VDD2.n44 4.38594
R1648 VDD2.n13 VDD2.n9 4.38594
R1649 VDD2.n59 VDD2.n37 4.26717
R1650 VDD2.n24 VDD2.n2 4.26717
R1651 VDD2.n58 VDD2.n39 3.49141
R1652 VDD2.n23 VDD2.n4 3.49141
R1653 VDD2.n69 VDD2.t3 3.29501
R1654 VDD2.n69 VDD2.t2 3.29501
R1655 VDD2.n67 VDD2.t8 3.29501
R1656 VDD2.n67 VDD2.t5 3.29501
R1657 VDD2.n33 VDD2.t4 3.29501
R1658 VDD2.n33 VDD2.t0 3.29501
R1659 VDD2.n31 VDD2.t1 3.29501
R1660 VDD2.n31 VDD2.t6 3.29501
R1661 VDD2.n55 VDD2.n54 2.71565
R1662 VDD2.n20 VDD2.n19 2.71565
R1663 VDD2.n51 VDD2.n41 1.93989
R1664 VDD2.n16 VDD2.n6 1.93989
R1665 VDD2.n68 VDD2.n66 1.19016
R1666 VDD2.n50 VDD2.n43 1.16414
R1667 VDD2.n15 VDD2.n8 1.16414
R1668 VDD2.n47 VDD2.n46 0.388379
R1669 VDD2.n12 VDD2.n11 0.388379
R1670 VDD2 VDD2.n68 0.356103
R1671 VDD2.n34 VDD2.n32 0.242568
R1672 VDD2.n64 VDD2.n36 0.155672
R1673 VDD2.n57 VDD2.n36 0.155672
R1674 VDD2.n57 VDD2.n56 0.155672
R1675 VDD2.n56 VDD2.n40 0.155672
R1676 VDD2.n49 VDD2.n40 0.155672
R1677 VDD2.n49 VDD2.n48 0.155672
R1678 VDD2.n14 VDD2.n13 0.155672
R1679 VDD2.n14 VDD2.n5 0.155672
R1680 VDD2.n21 VDD2.n5 0.155672
R1681 VDD2.n22 VDD2.n21 0.155672
R1682 VDD2.n22 VDD2.n1 0.155672
R1683 VDD2.n29 VDD2.n1 0.155672
C0 VTAIL VDD1 7.52815f
C1 VDD2 VP 0.385229f
C2 VDD2 VN 4.29198f
C3 VP VN 5.00086f
C4 VDD2 VTAIL 7.56863f
C5 VTAIL VP 4.63057f
C6 VTAIL VN 4.61626f
C7 VDD2 VDD1 1.19121f
C8 VP VDD1 4.52489f
C9 VDD1 VN 0.149756f
C10 VDD2 B 4.309072f
C11 VDD1 B 4.255907f
C12 VTAIL B 4.425582f
C13 VN B 10.27138f
C14 VP B 8.681831f
C15 VDD2.n0 B 0.033128f
C16 VDD2.n1 B 0.023456f
C17 VDD2.n2 B 0.012604f
C18 VDD2.n3 B 0.029792f
C19 VDD2.n4 B 0.013346f
C20 VDD2.n5 B 0.023456f
C21 VDD2.n6 B 0.012604f
C22 VDD2.n7 B 0.029792f
C23 VDD2.n8 B 0.013346f
C24 VDD2.n9 B 0.100442f
C25 VDD2.t9 B 0.048561f
C26 VDD2.n10 B 0.022344f
C27 VDD2.n11 B 0.017598f
C28 VDD2.n12 B 0.012604f
C29 VDD2.n13 B 0.559186f
C30 VDD2.n14 B 0.023456f
C31 VDD2.n15 B 0.012604f
C32 VDD2.n16 B 0.013346f
C33 VDD2.n17 B 0.029792f
C34 VDD2.n18 B 0.029792f
C35 VDD2.n19 B 0.013346f
C36 VDD2.n20 B 0.012604f
C37 VDD2.n21 B 0.023456f
C38 VDD2.n22 B 0.023456f
C39 VDD2.n23 B 0.012604f
C40 VDD2.n24 B 0.013346f
C41 VDD2.n25 B 0.029792f
C42 VDD2.n26 B 0.064775f
C43 VDD2.n27 B 0.013346f
C44 VDD2.n28 B 0.012604f
C45 VDD2.n29 B 0.054539f
C46 VDD2.n30 B 0.055679f
C47 VDD2.t1 B 0.111401f
C48 VDD2.t6 B 0.111401f
C49 VDD2.n31 B 0.929334f
C50 VDD2.n32 B 0.432868f
C51 VDD2.t4 B 0.111401f
C52 VDD2.t0 B 0.111401f
C53 VDD2.n33 B 0.933672f
C54 VDD2.n34 B 1.62233f
C55 VDD2.n35 B 0.033128f
C56 VDD2.n36 B 0.023456f
C57 VDD2.n37 B 0.012604f
C58 VDD2.n38 B 0.029792f
C59 VDD2.n39 B 0.013346f
C60 VDD2.n40 B 0.023456f
C61 VDD2.n41 B 0.012604f
C62 VDD2.n42 B 0.029792f
C63 VDD2.n43 B 0.013346f
C64 VDD2.n44 B 0.100442f
C65 VDD2.t7 B 0.048561f
C66 VDD2.n45 B 0.022344f
C67 VDD2.n46 B 0.017598f
C68 VDD2.n47 B 0.012604f
C69 VDD2.n48 B 0.559186f
C70 VDD2.n49 B 0.023456f
C71 VDD2.n50 B 0.012604f
C72 VDD2.n51 B 0.013346f
C73 VDD2.n52 B 0.029792f
C74 VDD2.n53 B 0.029792f
C75 VDD2.n54 B 0.013346f
C76 VDD2.n55 B 0.012604f
C77 VDD2.n56 B 0.023456f
C78 VDD2.n57 B 0.023456f
C79 VDD2.n58 B 0.012604f
C80 VDD2.n59 B 0.013346f
C81 VDD2.n60 B 0.029792f
C82 VDD2.n61 B 0.064775f
C83 VDD2.n62 B 0.013346f
C84 VDD2.n63 B 0.012604f
C85 VDD2.n64 B 0.054539f
C86 VDD2.n65 B 0.052476f
C87 VDD2.n66 B 1.70372f
C88 VDD2.t8 B 0.111401f
C89 VDD2.t5 B 0.111401f
C90 VDD2.n67 B 0.929338f
C91 VDD2.n68 B 0.307135f
C92 VDD2.t3 B 0.111401f
C93 VDD2.t2 B 0.111401f
C94 VDD2.n69 B 0.933647f
C95 VN.n0 B 0.050115f
C96 VN.t5 B 0.627355f
C97 VN.n1 B 0.032134f
C98 VN.n2 B 0.037557f
C99 VN.t3 B 0.627355f
C100 VN.n3 B 0.050318f
C101 VN.t0 B 0.713042f
C102 VN.t8 B 0.627355f
C103 VN.n4 B 0.289104f
C104 VN.n5 B 0.313434f
C105 VN.n6 B 0.162619f
C106 VN.n7 B 0.037557f
C107 VN.n8 B 0.032134f
C108 VN.n9 B 0.054345f
C109 VN.n10 B 0.255956f
C110 VN.n11 B 0.054345f
C111 VN.n12 B 0.037557f
C112 VN.n13 B 0.037557f
C113 VN.n14 B 0.037557f
C114 VN.n15 B 0.050318f
C115 VN.n16 B 0.255956f
C116 VN.n17 B 0.053022f
C117 VN.t9 B 0.68777f
C118 VN.n18 B 0.318025f
C119 VN.n19 B 0.035173f
C120 VN.n20 B 0.050115f
C121 VN.t1 B 0.627355f
C122 VN.n21 B 0.032134f
C123 VN.n22 B 0.037557f
C124 VN.t4 B 0.627355f
C125 VN.n23 B 0.050318f
C126 VN.t7 B 0.713042f
C127 VN.t6 B 0.627355f
C128 VN.n24 B 0.289104f
C129 VN.n25 B 0.313434f
C130 VN.n26 B 0.162619f
C131 VN.n27 B 0.037557f
C132 VN.n28 B 0.032134f
C133 VN.n29 B 0.054345f
C134 VN.n30 B 0.255956f
C135 VN.n31 B 0.054345f
C136 VN.n32 B 0.037557f
C137 VN.n33 B 0.037557f
C138 VN.n34 B 0.037557f
C139 VN.n35 B 0.050318f
C140 VN.n36 B 0.255956f
C141 VN.n37 B 0.053022f
C142 VN.t2 B 0.68777f
C143 VN.n38 B 0.318025f
C144 VN.n39 B 1.48562f
C145 VDD1.n0 B 0.033165f
C146 VDD1.n1 B 0.023482f
C147 VDD1.n2 B 0.012618f
C148 VDD1.n3 B 0.029825f
C149 VDD1.n4 B 0.013361f
C150 VDD1.n5 B 0.023482f
C151 VDD1.n6 B 0.012618f
C152 VDD1.n7 B 0.029825f
C153 VDD1.n8 B 0.013361f
C154 VDD1.n9 B 0.100554f
C155 VDD1.t3 B 0.048615f
C156 VDD1.n10 B 0.022369f
C157 VDD1.n11 B 0.017618f
C158 VDD1.n12 B 0.012618f
C159 VDD1.n13 B 0.55981f
C160 VDD1.n14 B 0.023482f
C161 VDD1.n15 B 0.012618f
C162 VDD1.n16 B 0.013361f
C163 VDD1.n17 B 0.029825f
C164 VDD1.n18 B 0.029825f
C165 VDD1.n19 B 0.013361f
C166 VDD1.n20 B 0.012618f
C167 VDD1.n21 B 0.023482f
C168 VDD1.n22 B 0.023482f
C169 VDD1.n23 B 0.012618f
C170 VDD1.n24 B 0.013361f
C171 VDD1.n25 B 0.029825f
C172 VDD1.n26 B 0.064847f
C173 VDD1.n27 B 0.013361f
C174 VDD1.n28 B 0.012618f
C175 VDD1.n29 B 0.054599f
C176 VDD1.n30 B 0.055741f
C177 VDD1.t4 B 0.111525f
C178 VDD1.t5 B 0.111525f
C179 VDD1.n31 B 0.930375f
C180 VDD1.n32 B 0.439688f
C181 VDD1.n33 B 0.033165f
C182 VDD1.n34 B 0.023482f
C183 VDD1.n35 B 0.012618f
C184 VDD1.n36 B 0.029825f
C185 VDD1.n37 B 0.013361f
C186 VDD1.n38 B 0.023482f
C187 VDD1.n39 B 0.012618f
C188 VDD1.n40 B 0.029825f
C189 VDD1.n41 B 0.013361f
C190 VDD1.n42 B 0.100554f
C191 VDD1.t2 B 0.048615f
C192 VDD1.n43 B 0.022369f
C193 VDD1.n44 B 0.017618f
C194 VDD1.n45 B 0.012618f
C195 VDD1.n46 B 0.55981f
C196 VDD1.n47 B 0.023482f
C197 VDD1.n48 B 0.012618f
C198 VDD1.n49 B 0.013361f
C199 VDD1.n50 B 0.029825f
C200 VDD1.n51 B 0.029825f
C201 VDD1.n52 B 0.013361f
C202 VDD1.n53 B 0.012618f
C203 VDD1.n54 B 0.023482f
C204 VDD1.n55 B 0.023482f
C205 VDD1.n56 B 0.012618f
C206 VDD1.n57 B 0.013361f
C207 VDD1.n58 B 0.029825f
C208 VDD1.n59 B 0.064847f
C209 VDD1.n60 B 0.013361f
C210 VDD1.n61 B 0.012618f
C211 VDD1.n62 B 0.054599f
C212 VDD1.n63 B 0.055741f
C213 VDD1.t6 B 0.111525f
C214 VDD1.t0 B 0.111525f
C215 VDD1.n64 B 0.93037f
C216 VDD1.n65 B 0.433351f
C217 VDD1.t1 B 0.111525f
C218 VDD1.t7 B 0.111525f
C219 VDD1.n66 B 0.934713f
C220 VDD1.n67 B 1.70142f
C221 VDD1.t8 B 0.111525f
C222 VDD1.t9 B 0.111525f
C223 VDD1.n68 B 0.93037f
C224 VDD1.n69 B 1.93279f
C225 VTAIL.t0 B 0.127738f
C226 VTAIL.t8 B 0.127738f
C227 VTAIL.n0 B 0.995512f
C228 VTAIL.n1 B 0.426451f
C229 VTAIL.n2 B 0.037986f
C230 VTAIL.n3 B 0.026896f
C231 VTAIL.n4 B 0.014453f
C232 VTAIL.n5 B 0.034161f
C233 VTAIL.n6 B 0.015303f
C234 VTAIL.n7 B 0.026896f
C235 VTAIL.n8 B 0.014453f
C236 VTAIL.n9 B 0.034161f
C237 VTAIL.n10 B 0.015303f
C238 VTAIL.n11 B 0.115171f
C239 VTAIL.t16 B 0.055683f
C240 VTAIL.n12 B 0.025621f
C241 VTAIL.n13 B 0.020179f
C242 VTAIL.n14 B 0.014453f
C243 VTAIL.n15 B 0.641191f
C244 VTAIL.n16 B 0.026896f
C245 VTAIL.n17 B 0.014453f
C246 VTAIL.n18 B 0.015303f
C247 VTAIL.n19 B 0.034161f
C248 VTAIL.n20 B 0.034161f
C249 VTAIL.n21 B 0.015303f
C250 VTAIL.n22 B 0.014453f
C251 VTAIL.n23 B 0.026896f
C252 VTAIL.n24 B 0.026896f
C253 VTAIL.n25 B 0.014453f
C254 VTAIL.n26 B 0.015303f
C255 VTAIL.n27 B 0.034161f
C256 VTAIL.n28 B 0.074274f
C257 VTAIL.n29 B 0.015303f
C258 VTAIL.n30 B 0.014453f
C259 VTAIL.n31 B 0.062537f
C260 VTAIL.n32 B 0.041604f
C261 VTAIL.n33 B 0.21855f
C262 VTAIL.t9 B 0.127738f
C263 VTAIL.t18 B 0.127738f
C264 VTAIL.n34 B 0.995512f
C265 VTAIL.n35 B 0.458017f
C266 VTAIL.t13 B 0.127738f
C267 VTAIL.t17 B 0.127738f
C268 VTAIL.n36 B 0.995512f
C269 VTAIL.n37 B 1.37549f
C270 VTAIL.t3 B 0.127738f
C271 VTAIL.t4 B 0.127738f
C272 VTAIL.n38 B 0.995519f
C273 VTAIL.n39 B 1.37548f
C274 VTAIL.t5 B 0.127738f
C275 VTAIL.t19 B 0.127738f
C276 VTAIL.n40 B 0.995519f
C277 VTAIL.n41 B 0.45801f
C278 VTAIL.n42 B 0.037986f
C279 VTAIL.n43 B 0.026896f
C280 VTAIL.n44 B 0.014453f
C281 VTAIL.n45 B 0.034161f
C282 VTAIL.n46 B 0.015303f
C283 VTAIL.n47 B 0.026896f
C284 VTAIL.n48 B 0.014453f
C285 VTAIL.n49 B 0.034161f
C286 VTAIL.n50 B 0.015303f
C287 VTAIL.n51 B 0.115171f
C288 VTAIL.t2 B 0.055683f
C289 VTAIL.n52 B 0.025621f
C290 VTAIL.n53 B 0.020179f
C291 VTAIL.n54 B 0.014453f
C292 VTAIL.n55 B 0.641191f
C293 VTAIL.n56 B 0.026896f
C294 VTAIL.n57 B 0.014453f
C295 VTAIL.n58 B 0.015303f
C296 VTAIL.n59 B 0.034161f
C297 VTAIL.n60 B 0.034161f
C298 VTAIL.n61 B 0.015303f
C299 VTAIL.n62 B 0.014453f
C300 VTAIL.n63 B 0.026896f
C301 VTAIL.n64 B 0.026896f
C302 VTAIL.n65 B 0.014453f
C303 VTAIL.n66 B 0.015303f
C304 VTAIL.n67 B 0.034161f
C305 VTAIL.n68 B 0.074274f
C306 VTAIL.n69 B 0.015303f
C307 VTAIL.n70 B 0.014453f
C308 VTAIL.n71 B 0.062537f
C309 VTAIL.n72 B 0.041604f
C310 VTAIL.n73 B 0.21855f
C311 VTAIL.t11 B 0.127738f
C312 VTAIL.t10 B 0.127738f
C313 VTAIL.n74 B 0.995519f
C314 VTAIL.n75 B 0.447177f
C315 VTAIL.t14 B 0.127738f
C316 VTAIL.t12 B 0.127738f
C317 VTAIL.n76 B 0.995519f
C318 VTAIL.n77 B 0.45801f
C319 VTAIL.n78 B 0.037986f
C320 VTAIL.n79 B 0.026896f
C321 VTAIL.n80 B 0.014453f
C322 VTAIL.n81 B 0.034161f
C323 VTAIL.n82 B 0.015303f
C324 VTAIL.n83 B 0.026896f
C325 VTAIL.n84 B 0.014453f
C326 VTAIL.n85 B 0.034161f
C327 VTAIL.n86 B 0.015303f
C328 VTAIL.n87 B 0.115171f
C329 VTAIL.t15 B 0.055683f
C330 VTAIL.n88 B 0.025621f
C331 VTAIL.n89 B 0.020179f
C332 VTAIL.n90 B 0.014453f
C333 VTAIL.n91 B 0.641191f
C334 VTAIL.n92 B 0.026896f
C335 VTAIL.n93 B 0.014453f
C336 VTAIL.n94 B 0.015303f
C337 VTAIL.n95 B 0.034161f
C338 VTAIL.n96 B 0.034161f
C339 VTAIL.n97 B 0.015303f
C340 VTAIL.n98 B 0.014453f
C341 VTAIL.n99 B 0.026896f
C342 VTAIL.n100 B 0.026896f
C343 VTAIL.n101 B 0.014453f
C344 VTAIL.n102 B 0.015303f
C345 VTAIL.n103 B 0.034161f
C346 VTAIL.n104 B 0.074274f
C347 VTAIL.n105 B 0.015303f
C348 VTAIL.n106 B 0.014453f
C349 VTAIL.n107 B 0.062537f
C350 VTAIL.n108 B 0.041604f
C351 VTAIL.n109 B 1.04375f
C352 VTAIL.n110 B 0.037986f
C353 VTAIL.n111 B 0.026896f
C354 VTAIL.n112 B 0.014453f
C355 VTAIL.n113 B 0.034161f
C356 VTAIL.n114 B 0.015303f
C357 VTAIL.n115 B 0.026896f
C358 VTAIL.n116 B 0.014453f
C359 VTAIL.n117 B 0.034161f
C360 VTAIL.n118 B 0.015303f
C361 VTAIL.n119 B 0.115171f
C362 VTAIL.t1 B 0.055683f
C363 VTAIL.n120 B 0.025621f
C364 VTAIL.n121 B 0.020179f
C365 VTAIL.n122 B 0.014453f
C366 VTAIL.n123 B 0.641191f
C367 VTAIL.n124 B 0.026896f
C368 VTAIL.n125 B 0.014453f
C369 VTAIL.n126 B 0.015303f
C370 VTAIL.n127 B 0.034161f
C371 VTAIL.n128 B 0.034161f
C372 VTAIL.n129 B 0.015303f
C373 VTAIL.n130 B 0.014453f
C374 VTAIL.n131 B 0.026896f
C375 VTAIL.n132 B 0.026896f
C376 VTAIL.n133 B 0.014453f
C377 VTAIL.n134 B 0.015303f
C378 VTAIL.n135 B 0.034161f
C379 VTAIL.n136 B 0.074274f
C380 VTAIL.n137 B 0.015303f
C381 VTAIL.n138 B 0.014453f
C382 VTAIL.n139 B 0.062537f
C383 VTAIL.n140 B 0.041604f
C384 VTAIL.n141 B 1.04375f
C385 VTAIL.t6 B 0.127738f
C386 VTAIL.t7 B 0.127738f
C387 VTAIL.n142 B 0.995512f
C388 VTAIL.n143 B 0.375648f
C389 VP.n0 B 0.05103f
C390 VP.t8 B 0.638808f
C391 VP.n1 B 0.032721f
C392 VP.n2 B 0.038243f
C393 VP.t9 B 0.638808f
C394 VP.n3 B 0.051237f
C395 VP.n4 B 0.05103f
C396 VP.t0 B 0.700326f
C397 VP.t1 B 0.638808f
C398 VP.n5 B 0.032721f
C399 VP.n6 B 0.038243f
C400 VP.t4 B 0.638808f
C401 VP.n7 B 0.051237f
C402 VP.t5 B 0.638808f
C403 VP.n8 B 0.294381f
C404 VP.t6 B 0.726059f
C405 VP.n9 B 0.319156f
C406 VP.n10 B 0.165588f
C407 VP.n11 B 0.038243f
C408 VP.n12 B 0.032721f
C409 VP.n13 B 0.055337f
C410 VP.n14 B 0.260628f
C411 VP.n15 B 0.055337f
C412 VP.n16 B 0.038243f
C413 VP.n17 B 0.038243f
C414 VP.n18 B 0.038243f
C415 VP.n19 B 0.051237f
C416 VP.n20 B 0.260628f
C417 VP.n21 B 0.05399f
C418 VP.n22 B 0.32383f
C419 VP.n23 B 1.49114f
C420 VP.n24 B 1.52517f
C421 VP.t7 B 0.700326f
C422 VP.n25 B 0.32383f
C423 VP.t3 B 0.638808f
C424 VP.n26 B 0.260628f
C425 VP.n27 B 0.05399f
C426 VP.n28 B 0.05103f
C427 VP.n29 B 0.038243f
C428 VP.n30 B 0.038243f
C429 VP.n31 B 0.032721f
C430 VP.n32 B 0.055337f
C431 VP.n33 B 0.260628f
C432 VP.n34 B 0.055337f
C433 VP.n35 B 0.038243f
C434 VP.n36 B 0.038243f
C435 VP.n37 B 0.038243f
C436 VP.n38 B 0.051237f
C437 VP.n39 B 0.260628f
C438 VP.n40 B 0.05399f
C439 VP.t2 B 0.700326f
C440 VP.n41 B 0.32383f
C441 VP.n42 B 0.035816f
.ends

