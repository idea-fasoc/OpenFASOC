* NGSPICE file created from diff_pair_sample_0699.ext - technology: sky130A

.subckt diff_pair_sample_0699 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=0 ps=0 w=15.77 l=2.08
X1 B.t8 B.t6 B.t7 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=0 ps=0 w=15.77 l=2.08
X2 B.t5 B.t3 B.t4 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=0 ps=0 w=15.77 l=2.08
X3 VDD1.t3 VP.t0 VTAIL.t6 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=2.60205 pd=16.1 as=6.1503 ps=32.32 w=15.77 l=2.08
X4 VTAIL.t1 VN.t0 VDD2.t3 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=2.60205 ps=16.1 w=15.77 l=2.08
X5 VDD2.t2 VN.t1 VTAIL.t2 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=2.60205 pd=16.1 as=6.1503 ps=32.32 w=15.77 l=2.08
X6 VDD1.t2 VP.t1 VTAIL.t4 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=2.60205 pd=16.1 as=6.1503 ps=32.32 w=15.77 l=2.08
X7 VDD2.t1 VN.t2 VTAIL.t0 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=2.60205 pd=16.1 as=6.1503 ps=32.32 w=15.77 l=2.08
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=2.60205 ps=16.1 w=15.77 l=2.08
X9 B.t2 B.t0 B.t1 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=0 ps=0 w=15.77 l=2.08
X10 VTAIL.t5 VP.t2 VDD1.t1 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=2.60205 ps=16.1 w=15.77 l=2.08
X11 VTAIL.t7 VP.t3 VDD1.t0 w_n2416_n4122# sky130_fd_pr__pfet_01v8 ad=6.1503 pd=32.32 as=2.60205 ps=16.1 w=15.77 l=2.08
R0 B.n399 B.n108 585
R1 B.n398 B.n397 585
R2 B.n396 B.n109 585
R3 B.n395 B.n394 585
R4 B.n393 B.n110 585
R5 B.n392 B.n391 585
R6 B.n390 B.n111 585
R7 B.n389 B.n388 585
R8 B.n387 B.n112 585
R9 B.n386 B.n385 585
R10 B.n384 B.n113 585
R11 B.n383 B.n382 585
R12 B.n381 B.n114 585
R13 B.n380 B.n379 585
R14 B.n378 B.n115 585
R15 B.n377 B.n376 585
R16 B.n375 B.n116 585
R17 B.n374 B.n373 585
R18 B.n372 B.n117 585
R19 B.n371 B.n370 585
R20 B.n369 B.n118 585
R21 B.n368 B.n367 585
R22 B.n366 B.n119 585
R23 B.n365 B.n364 585
R24 B.n363 B.n120 585
R25 B.n362 B.n361 585
R26 B.n360 B.n121 585
R27 B.n359 B.n358 585
R28 B.n357 B.n122 585
R29 B.n356 B.n355 585
R30 B.n354 B.n123 585
R31 B.n353 B.n352 585
R32 B.n351 B.n124 585
R33 B.n350 B.n349 585
R34 B.n348 B.n125 585
R35 B.n347 B.n346 585
R36 B.n345 B.n126 585
R37 B.n344 B.n343 585
R38 B.n342 B.n127 585
R39 B.n341 B.n340 585
R40 B.n339 B.n128 585
R41 B.n338 B.n337 585
R42 B.n336 B.n129 585
R43 B.n335 B.n334 585
R44 B.n333 B.n130 585
R45 B.n332 B.n331 585
R46 B.n330 B.n131 585
R47 B.n329 B.n328 585
R48 B.n327 B.n132 585
R49 B.n326 B.n325 585
R50 B.n324 B.n133 585
R51 B.n323 B.n322 585
R52 B.n321 B.n134 585
R53 B.n320 B.n319 585
R54 B.n315 B.n135 585
R55 B.n314 B.n313 585
R56 B.n312 B.n136 585
R57 B.n311 B.n310 585
R58 B.n309 B.n137 585
R59 B.n308 B.n307 585
R60 B.n306 B.n138 585
R61 B.n305 B.n304 585
R62 B.n302 B.n139 585
R63 B.n301 B.n300 585
R64 B.n299 B.n142 585
R65 B.n298 B.n297 585
R66 B.n296 B.n143 585
R67 B.n295 B.n294 585
R68 B.n293 B.n144 585
R69 B.n292 B.n291 585
R70 B.n290 B.n145 585
R71 B.n289 B.n288 585
R72 B.n287 B.n146 585
R73 B.n286 B.n285 585
R74 B.n284 B.n147 585
R75 B.n283 B.n282 585
R76 B.n281 B.n148 585
R77 B.n280 B.n279 585
R78 B.n278 B.n149 585
R79 B.n277 B.n276 585
R80 B.n275 B.n150 585
R81 B.n274 B.n273 585
R82 B.n272 B.n151 585
R83 B.n271 B.n270 585
R84 B.n269 B.n152 585
R85 B.n268 B.n267 585
R86 B.n266 B.n153 585
R87 B.n265 B.n264 585
R88 B.n263 B.n154 585
R89 B.n262 B.n261 585
R90 B.n260 B.n155 585
R91 B.n259 B.n258 585
R92 B.n257 B.n156 585
R93 B.n256 B.n255 585
R94 B.n254 B.n157 585
R95 B.n253 B.n252 585
R96 B.n251 B.n158 585
R97 B.n250 B.n249 585
R98 B.n248 B.n159 585
R99 B.n247 B.n246 585
R100 B.n245 B.n160 585
R101 B.n244 B.n243 585
R102 B.n242 B.n161 585
R103 B.n241 B.n240 585
R104 B.n239 B.n162 585
R105 B.n238 B.n237 585
R106 B.n236 B.n163 585
R107 B.n235 B.n234 585
R108 B.n233 B.n164 585
R109 B.n232 B.n231 585
R110 B.n230 B.n165 585
R111 B.n229 B.n228 585
R112 B.n227 B.n166 585
R113 B.n226 B.n225 585
R114 B.n224 B.n167 585
R115 B.n401 B.n400 585
R116 B.n402 B.n107 585
R117 B.n404 B.n403 585
R118 B.n405 B.n106 585
R119 B.n407 B.n406 585
R120 B.n408 B.n105 585
R121 B.n410 B.n409 585
R122 B.n411 B.n104 585
R123 B.n413 B.n412 585
R124 B.n414 B.n103 585
R125 B.n416 B.n415 585
R126 B.n417 B.n102 585
R127 B.n419 B.n418 585
R128 B.n420 B.n101 585
R129 B.n422 B.n421 585
R130 B.n423 B.n100 585
R131 B.n425 B.n424 585
R132 B.n426 B.n99 585
R133 B.n428 B.n427 585
R134 B.n429 B.n98 585
R135 B.n431 B.n430 585
R136 B.n432 B.n97 585
R137 B.n434 B.n433 585
R138 B.n435 B.n96 585
R139 B.n437 B.n436 585
R140 B.n438 B.n95 585
R141 B.n440 B.n439 585
R142 B.n441 B.n94 585
R143 B.n443 B.n442 585
R144 B.n444 B.n93 585
R145 B.n446 B.n445 585
R146 B.n447 B.n92 585
R147 B.n449 B.n448 585
R148 B.n450 B.n91 585
R149 B.n452 B.n451 585
R150 B.n453 B.n90 585
R151 B.n455 B.n454 585
R152 B.n456 B.n89 585
R153 B.n458 B.n457 585
R154 B.n459 B.n88 585
R155 B.n461 B.n460 585
R156 B.n462 B.n87 585
R157 B.n464 B.n463 585
R158 B.n465 B.n86 585
R159 B.n467 B.n466 585
R160 B.n468 B.n85 585
R161 B.n470 B.n469 585
R162 B.n471 B.n84 585
R163 B.n473 B.n472 585
R164 B.n474 B.n83 585
R165 B.n476 B.n475 585
R166 B.n477 B.n82 585
R167 B.n479 B.n478 585
R168 B.n480 B.n81 585
R169 B.n482 B.n481 585
R170 B.n483 B.n80 585
R171 B.n485 B.n484 585
R172 B.n486 B.n79 585
R173 B.n488 B.n487 585
R174 B.n489 B.n78 585
R175 B.n664 B.n663 585
R176 B.n662 B.n17 585
R177 B.n661 B.n660 585
R178 B.n659 B.n18 585
R179 B.n658 B.n657 585
R180 B.n656 B.n19 585
R181 B.n655 B.n654 585
R182 B.n653 B.n20 585
R183 B.n652 B.n651 585
R184 B.n650 B.n21 585
R185 B.n649 B.n648 585
R186 B.n647 B.n22 585
R187 B.n646 B.n645 585
R188 B.n644 B.n23 585
R189 B.n643 B.n642 585
R190 B.n641 B.n24 585
R191 B.n640 B.n639 585
R192 B.n638 B.n25 585
R193 B.n637 B.n636 585
R194 B.n635 B.n26 585
R195 B.n634 B.n633 585
R196 B.n632 B.n27 585
R197 B.n631 B.n630 585
R198 B.n629 B.n28 585
R199 B.n628 B.n627 585
R200 B.n626 B.n29 585
R201 B.n625 B.n624 585
R202 B.n623 B.n30 585
R203 B.n622 B.n621 585
R204 B.n620 B.n31 585
R205 B.n619 B.n618 585
R206 B.n617 B.n32 585
R207 B.n616 B.n615 585
R208 B.n614 B.n33 585
R209 B.n613 B.n612 585
R210 B.n611 B.n34 585
R211 B.n610 B.n609 585
R212 B.n608 B.n35 585
R213 B.n607 B.n606 585
R214 B.n605 B.n36 585
R215 B.n604 B.n603 585
R216 B.n602 B.n37 585
R217 B.n601 B.n600 585
R218 B.n599 B.n38 585
R219 B.n598 B.n597 585
R220 B.n596 B.n39 585
R221 B.n595 B.n594 585
R222 B.n593 B.n40 585
R223 B.n592 B.n591 585
R224 B.n590 B.n41 585
R225 B.n589 B.n588 585
R226 B.n587 B.n42 585
R227 B.n586 B.n585 585
R228 B.n583 B.n43 585
R229 B.n582 B.n581 585
R230 B.n580 B.n46 585
R231 B.n579 B.n578 585
R232 B.n577 B.n47 585
R233 B.n576 B.n575 585
R234 B.n574 B.n48 585
R235 B.n573 B.n572 585
R236 B.n571 B.n49 585
R237 B.n569 B.n568 585
R238 B.n567 B.n52 585
R239 B.n566 B.n565 585
R240 B.n564 B.n53 585
R241 B.n563 B.n562 585
R242 B.n561 B.n54 585
R243 B.n560 B.n559 585
R244 B.n558 B.n55 585
R245 B.n557 B.n556 585
R246 B.n555 B.n56 585
R247 B.n554 B.n553 585
R248 B.n552 B.n57 585
R249 B.n551 B.n550 585
R250 B.n549 B.n58 585
R251 B.n548 B.n547 585
R252 B.n546 B.n59 585
R253 B.n545 B.n544 585
R254 B.n543 B.n60 585
R255 B.n542 B.n541 585
R256 B.n540 B.n61 585
R257 B.n539 B.n538 585
R258 B.n537 B.n62 585
R259 B.n536 B.n535 585
R260 B.n534 B.n63 585
R261 B.n533 B.n532 585
R262 B.n531 B.n64 585
R263 B.n530 B.n529 585
R264 B.n528 B.n65 585
R265 B.n527 B.n526 585
R266 B.n525 B.n66 585
R267 B.n524 B.n523 585
R268 B.n522 B.n67 585
R269 B.n521 B.n520 585
R270 B.n519 B.n68 585
R271 B.n518 B.n517 585
R272 B.n516 B.n69 585
R273 B.n515 B.n514 585
R274 B.n513 B.n70 585
R275 B.n512 B.n511 585
R276 B.n510 B.n71 585
R277 B.n509 B.n508 585
R278 B.n507 B.n72 585
R279 B.n506 B.n505 585
R280 B.n504 B.n73 585
R281 B.n503 B.n502 585
R282 B.n501 B.n74 585
R283 B.n500 B.n499 585
R284 B.n498 B.n75 585
R285 B.n497 B.n496 585
R286 B.n495 B.n76 585
R287 B.n494 B.n493 585
R288 B.n492 B.n77 585
R289 B.n491 B.n490 585
R290 B.n665 B.n16 585
R291 B.n667 B.n666 585
R292 B.n668 B.n15 585
R293 B.n670 B.n669 585
R294 B.n671 B.n14 585
R295 B.n673 B.n672 585
R296 B.n674 B.n13 585
R297 B.n676 B.n675 585
R298 B.n677 B.n12 585
R299 B.n679 B.n678 585
R300 B.n680 B.n11 585
R301 B.n682 B.n681 585
R302 B.n683 B.n10 585
R303 B.n685 B.n684 585
R304 B.n686 B.n9 585
R305 B.n688 B.n687 585
R306 B.n689 B.n8 585
R307 B.n691 B.n690 585
R308 B.n692 B.n7 585
R309 B.n694 B.n693 585
R310 B.n695 B.n6 585
R311 B.n697 B.n696 585
R312 B.n698 B.n5 585
R313 B.n700 B.n699 585
R314 B.n701 B.n4 585
R315 B.n703 B.n702 585
R316 B.n704 B.n3 585
R317 B.n706 B.n705 585
R318 B.n707 B.n0 585
R319 B.n2 B.n1 585
R320 B.n182 B.n181 585
R321 B.n184 B.n183 585
R322 B.n185 B.n180 585
R323 B.n187 B.n186 585
R324 B.n188 B.n179 585
R325 B.n190 B.n189 585
R326 B.n191 B.n178 585
R327 B.n193 B.n192 585
R328 B.n194 B.n177 585
R329 B.n196 B.n195 585
R330 B.n197 B.n176 585
R331 B.n199 B.n198 585
R332 B.n200 B.n175 585
R333 B.n202 B.n201 585
R334 B.n203 B.n174 585
R335 B.n205 B.n204 585
R336 B.n206 B.n173 585
R337 B.n208 B.n207 585
R338 B.n209 B.n172 585
R339 B.n211 B.n210 585
R340 B.n212 B.n171 585
R341 B.n214 B.n213 585
R342 B.n215 B.n170 585
R343 B.n217 B.n216 585
R344 B.n218 B.n169 585
R345 B.n220 B.n219 585
R346 B.n221 B.n168 585
R347 B.n223 B.n222 585
R348 B.n222 B.n167 478.086
R349 B.n400 B.n399 478.086
R350 B.n490 B.n489 478.086
R351 B.n665 B.n664 478.086
R352 B.n140 B.t3 389.82
R353 B.n316 B.t6 389.82
R354 B.n50 B.t9 389.82
R355 B.n44 B.t0 389.82
R356 B.n709 B.n708 256.663
R357 B.n708 B.n707 235.042
R358 B.n708 B.n2 235.042
R359 B.n226 B.n167 163.367
R360 B.n227 B.n226 163.367
R361 B.n228 B.n227 163.367
R362 B.n228 B.n165 163.367
R363 B.n232 B.n165 163.367
R364 B.n233 B.n232 163.367
R365 B.n234 B.n233 163.367
R366 B.n234 B.n163 163.367
R367 B.n238 B.n163 163.367
R368 B.n239 B.n238 163.367
R369 B.n240 B.n239 163.367
R370 B.n240 B.n161 163.367
R371 B.n244 B.n161 163.367
R372 B.n245 B.n244 163.367
R373 B.n246 B.n245 163.367
R374 B.n246 B.n159 163.367
R375 B.n250 B.n159 163.367
R376 B.n251 B.n250 163.367
R377 B.n252 B.n251 163.367
R378 B.n252 B.n157 163.367
R379 B.n256 B.n157 163.367
R380 B.n257 B.n256 163.367
R381 B.n258 B.n257 163.367
R382 B.n258 B.n155 163.367
R383 B.n262 B.n155 163.367
R384 B.n263 B.n262 163.367
R385 B.n264 B.n263 163.367
R386 B.n264 B.n153 163.367
R387 B.n268 B.n153 163.367
R388 B.n269 B.n268 163.367
R389 B.n270 B.n269 163.367
R390 B.n270 B.n151 163.367
R391 B.n274 B.n151 163.367
R392 B.n275 B.n274 163.367
R393 B.n276 B.n275 163.367
R394 B.n276 B.n149 163.367
R395 B.n280 B.n149 163.367
R396 B.n281 B.n280 163.367
R397 B.n282 B.n281 163.367
R398 B.n282 B.n147 163.367
R399 B.n286 B.n147 163.367
R400 B.n287 B.n286 163.367
R401 B.n288 B.n287 163.367
R402 B.n288 B.n145 163.367
R403 B.n292 B.n145 163.367
R404 B.n293 B.n292 163.367
R405 B.n294 B.n293 163.367
R406 B.n294 B.n143 163.367
R407 B.n298 B.n143 163.367
R408 B.n299 B.n298 163.367
R409 B.n300 B.n299 163.367
R410 B.n300 B.n139 163.367
R411 B.n305 B.n139 163.367
R412 B.n306 B.n305 163.367
R413 B.n307 B.n306 163.367
R414 B.n307 B.n137 163.367
R415 B.n311 B.n137 163.367
R416 B.n312 B.n311 163.367
R417 B.n313 B.n312 163.367
R418 B.n313 B.n135 163.367
R419 B.n320 B.n135 163.367
R420 B.n321 B.n320 163.367
R421 B.n322 B.n321 163.367
R422 B.n322 B.n133 163.367
R423 B.n326 B.n133 163.367
R424 B.n327 B.n326 163.367
R425 B.n328 B.n327 163.367
R426 B.n328 B.n131 163.367
R427 B.n332 B.n131 163.367
R428 B.n333 B.n332 163.367
R429 B.n334 B.n333 163.367
R430 B.n334 B.n129 163.367
R431 B.n338 B.n129 163.367
R432 B.n339 B.n338 163.367
R433 B.n340 B.n339 163.367
R434 B.n340 B.n127 163.367
R435 B.n344 B.n127 163.367
R436 B.n345 B.n344 163.367
R437 B.n346 B.n345 163.367
R438 B.n346 B.n125 163.367
R439 B.n350 B.n125 163.367
R440 B.n351 B.n350 163.367
R441 B.n352 B.n351 163.367
R442 B.n352 B.n123 163.367
R443 B.n356 B.n123 163.367
R444 B.n357 B.n356 163.367
R445 B.n358 B.n357 163.367
R446 B.n358 B.n121 163.367
R447 B.n362 B.n121 163.367
R448 B.n363 B.n362 163.367
R449 B.n364 B.n363 163.367
R450 B.n364 B.n119 163.367
R451 B.n368 B.n119 163.367
R452 B.n369 B.n368 163.367
R453 B.n370 B.n369 163.367
R454 B.n370 B.n117 163.367
R455 B.n374 B.n117 163.367
R456 B.n375 B.n374 163.367
R457 B.n376 B.n375 163.367
R458 B.n376 B.n115 163.367
R459 B.n380 B.n115 163.367
R460 B.n381 B.n380 163.367
R461 B.n382 B.n381 163.367
R462 B.n382 B.n113 163.367
R463 B.n386 B.n113 163.367
R464 B.n387 B.n386 163.367
R465 B.n388 B.n387 163.367
R466 B.n388 B.n111 163.367
R467 B.n392 B.n111 163.367
R468 B.n393 B.n392 163.367
R469 B.n394 B.n393 163.367
R470 B.n394 B.n109 163.367
R471 B.n398 B.n109 163.367
R472 B.n399 B.n398 163.367
R473 B.n489 B.n488 163.367
R474 B.n488 B.n79 163.367
R475 B.n484 B.n79 163.367
R476 B.n484 B.n483 163.367
R477 B.n483 B.n482 163.367
R478 B.n482 B.n81 163.367
R479 B.n478 B.n81 163.367
R480 B.n478 B.n477 163.367
R481 B.n477 B.n476 163.367
R482 B.n476 B.n83 163.367
R483 B.n472 B.n83 163.367
R484 B.n472 B.n471 163.367
R485 B.n471 B.n470 163.367
R486 B.n470 B.n85 163.367
R487 B.n466 B.n85 163.367
R488 B.n466 B.n465 163.367
R489 B.n465 B.n464 163.367
R490 B.n464 B.n87 163.367
R491 B.n460 B.n87 163.367
R492 B.n460 B.n459 163.367
R493 B.n459 B.n458 163.367
R494 B.n458 B.n89 163.367
R495 B.n454 B.n89 163.367
R496 B.n454 B.n453 163.367
R497 B.n453 B.n452 163.367
R498 B.n452 B.n91 163.367
R499 B.n448 B.n91 163.367
R500 B.n448 B.n447 163.367
R501 B.n447 B.n446 163.367
R502 B.n446 B.n93 163.367
R503 B.n442 B.n93 163.367
R504 B.n442 B.n441 163.367
R505 B.n441 B.n440 163.367
R506 B.n440 B.n95 163.367
R507 B.n436 B.n95 163.367
R508 B.n436 B.n435 163.367
R509 B.n435 B.n434 163.367
R510 B.n434 B.n97 163.367
R511 B.n430 B.n97 163.367
R512 B.n430 B.n429 163.367
R513 B.n429 B.n428 163.367
R514 B.n428 B.n99 163.367
R515 B.n424 B.n99 163.367
R516 B.n424 B.n423 163.367
R517 B.n423 B.n422 163.367
R518 B.n422 B.n101 163.367
R519 B.n418 B.n101 163.367
R520 B.n418 B.n417 163.367
R521 B.n417 B.n416 163.367
R522 B.n416 B.n103 163.367
R523 B.n412 B.n103 163.367
R524 B.n412 B.n411 163.367
R525 B.n411 B.n410 163.367
R526 B.n410 B.n105 163.367
R527 B.n406 B.n105 163.367
R528 B.n406 B.n405 163.367
R529 B.n405 B.n404 163.367
R530 B.n404 B.n107 163.367
R531 B.n400 B.n107 163.367
R532 B.n664 B.n17 163.367
R533 B.n660 B.n17 163.367
R534 B.n660 B.n659 163.367
R535 B.n659 B.n658 163.367
R536 B.n658 B.n19 163.367
R537 B.n654 B.n19 163.367
R538 B.n654 B.n653 163.367
R539 B.n653 B.n652 163.367
R540 B.n652 B.n21 163.367
R541 B.n648 B.n21 163.367
R542 B.n648 B.n647 163.367
R543 B.n647 B.n646 163.367
R544 B.n646 B.n23 163.367
R545 B.n642 B.n23 163.367
R546 B.n642 B.n641 163.367
R547 B.n641 B.n640 163.367
R548 B.n640 B.n25 163.367
R549 B.n636 B.n25 163.367
R550 B.n636 B.n635 163.367
R551 B.n635 B.n634 163.367
R552 B.n634 B.n27 163.367
R553 B.n630 B.n27 163.367
R554 B.n630 B.n629 163.367
R555 B.n629 B.n628 163.367
R556 B.n628 B.n29 163.367
R557 B.n624 B.n29 163.367
R558 B.n624 B.n623 163.367
R559 B.n623 B.n622 163.367
R560 B.n622 B.n31 163.367
R561 B.n618 B.n31 163.367
R562 B.n618 B.n617 163.367
R563 B.n617 B.n616 163.367
R564 B.n616 B.n33 163.367
R565 B.n612 B.n33 163.367
R566 B.n612 B.n611 163.367
R567 B.n611 B.n610 163.367
R568 B.n610 B.n35 163.367
R569 B.n606 B.n35 163.367
R570 B.n606 B.n605 163.367
R571 B.n605 B.n604 163.367
R572 B.n604 B.n37 163.367
R573 B.n600 B.n37 163.367
R574 B.n600 B.n599 163.367
R575 B.n599 B.n598 163.367
R576 B.n598 B.n39 163.367
R577 B.n594 B.n39 163.367
R578 B.n594 B.n593 163.367
R579 B.n593 B.n592 163.367
R580 B.n592 B.n41 163.367
R581 B.n588 B.n41 163.367
R582 B.n588 B.n587 163.367
R583 B.n587 B.n586 163.367
R584 B.n586 B.n43 163.367
R585 B.n581 B.n43 163.367
R586 B.n581 B.n580 163.367
R587 B.n580 B.n579 163.367
R588 B.n579 B.n47 163.367
R589 B.n575 B.n47 163.367
R590 B.n575 B.n574 163.367
R591 B.n574 B.n573 163.367
R592 B.n573 B.n49 163.367
R593 B.n568 B.n49 163.367
R594 B.n568 B.n567 163.367
R595 B.n567 B.n566 163.367
R596 B.n566 B.n53 163.367
R597 B.n562 B.n53 163.367
R598 B.n562 B.n561 163.367
R599 B.n561 B.n560 163.367
R600 B.n560 B.n55 163.367
R601 B.n556 B.n55 163.367
R602 B.n556 B.n555 163.367
R603 B.n555 B.n554 163.367
R604 B.n554 B.n57 163.367
R605 B.n550 B.n57 163.367
R606 B.n550 B.n549 163.367
R607 B.n549 B.n548 163.367
R608 B.n548 B.n59 163.367
R609 B.n544 B.n59 163.367
R610 B.n544 B.n543 163.367
R611 B.n543 B.n542 163.367
R612 B.n542 B.n61 163.367
R613 B.n538 B.n61 163.367
R614 B.n538 B.n537 163.367
R615 B.n537 B.n536 163.367
R616 B.n536 B.n63 163.367
R617 B.n532 B.n63 163.367
R618 B.n532 B.n531 163.367
R619 B.n531 B.n530 163.367
R620 B.n530 B.n65 163.367
R621 B.n526 B.n65 163.367
R622 B.n526 B.n525 163.367
R623 B.n525 B.n524 163.367
R624 B.n524 B.n67 163.367
R625 B.n520 B.n67 163.367
R626 B.n520 B.n519 163.367
R627 B.n519 B.n518 163.367
R628 B.n518 B.n69 163.367
R629 B.n514 B.n69 163.367
R630 B.n514 B.n513 163.367
R631 B.n513 B.n512 163.367
R632 B.n512 B.n71 163.367
R633 B.n508 B.n71 163.367
R634 B.n508 B.n507 163.367
R635 B.n507 B.n506 163.367
R636 B.n506 B.n73 163.367
R637 B.n502 B.n73 163.367
R638 B.n502 B.n501 163.367
R639 B.n501 B.n500 163.367
R640 B.n500 B.n75 163.367
R641 B.n496 B.n75 163.367
R642 B.n496 B.n495 163.367
R643 B.n495 B.n494 163.367
R644 B.n494 B.n77 163.367
R645 B.n490 B.n77 163.367
R646 B.n666 B.n665 163.367
R647 B.n666 B.n15 163.367
R648 B.n670 B.n15 163.367
R649 B.n671 B.n670 163.367
R650 B.n672 B.n671 163.367
R651 B.n672 B.n13 163.367
R652 B.n676 B.n13 163.367
R653 B.n677 B.n676 163.367
R654 B.n678 B.n677 163.367
R655 B.n678 B.n11 163.367
R656 B.n682 B.n11 163.367
R657 B.n683 B.n682 163.367
R658 B.n684 B.n683 163.367
R659 B.n684 B.n9 163.367
R660 B.n688 B.n9 163.367
R661 B.n689 B.n688 163.367
R662 B.n690 B.n689 163.367
R663 B.n690 B.n7 163.367
R664 B.n694 B.n7 163.367
R665 B.n695 B.n694 163.367
R666 B.n696 B.n695 163.367
R667 B.n696 B.n5 163.367
R668 B.n700 B.n5 163.367
R669 B.n701 B.n700 163.367
R670 B.n702 B.n701 163.367
R671 B.n702 B.n3 163.367
R672 B.n706 B.n3 163.367
R673 B.n707 B.n706 163.367
R674 B.n181 B.n2 163.367
R675 B.n184 B.n181 163.367
R676 B.n185 B.n184 163.367
R677 B.n186 B.n185 163.367
R678 B.n186 B.n179 163.367
R679 B.n190 B.n179 163.367
R680 B.n191 B.n190 163.367
R681 B.n192 B.n191 163.367
R682 B.n192 B.n177 163.367
R683 B.n196 B.n177 163.367
R684 B.n197 B.n196 163.367
R685 B.n198 B.n197 163.367
R686 B.n198 B.n175 163.367
R687 B.n202 B.n175 163.367
R688 B.n203 B.n202 163.367
R689 B.n204 B.n203 163.367
R690 B.n204 B.n173 163.367
R691 B.n208 B.n173 163.367
R692 B.n209 B.n208 163.367
R693 B.n210 B.n209 163.367
R694 B.n210 B.n171 163.367
R695 B.n214 B.n171 163.367
R696 B.n215 B.n214 163.367
R697 B.n216 B.n215 163.367
R698 B.n216 B.n169 163.367
R699 B.n220 B.n169 163.367
R700 B.n221 B.n220 163.367
R701 B.n222 B.n221 163.367
R702 B.n316 B.t7 155.716
R703 B.n50 B.t11 155.716
R704 B.n140 B.t4 155.696
R705 B.n44 B.t2 155.696
R706 B.n317 B.t8 108.978
R707 B.n51 B.t10 108.978
R708 B.n141 B.t5 108.957
R709 B.n45 B.t1 108.957
R710 B.n303 B.n141 59.5399
R711 B.n318 B.n317 59.5399
R712 B.n570 B.n51 59.5399
R713 B.n584 B.n45 59.5399
R714 B.n141 B.n140 46.7399
R715 B.n317 B.n316 46.7399
R716 B.n51 B.n50 46.7399
R717 B.n45 B.n44 46.7399
R718 B.n663 B.n16 31.0639
R719 B.n491 B.n78 31.0639
R720 B.n401 B.n108 31.0639
R721 B.n224 B.n223 31.0639
R722 B B.n709 18.0485
R723 B.n667 B.n16 10.6151
R724 B.n668 B.n667 10.6151
R725 B.n669 B.n668 10.6151
R726 B.n669 B.n14 10.6151
R727 B.n673 B.n14 10.6151
R728 B.n674 B.n673 10.6151
R729 B.n675 B.n674 10.6151
R730 B.n675 B.n12 10.6151
R731 B.n679 B.n12 10.6151
R732 B.n680 B.n679 10.6151
R733 B.n681 B.n680 10.6151
R734 B.n681 B.n10 10.6151
R735 B.n685 B.n10 10.6151
R736 B.n686 B.n685 10.6151
R737 B.n687 B.n686 10.6151
R738 B.n687 B.n8 10.6151
R739 B.n691 B.n8 10.6151
R740 B.n692 B.n691 10.6151
R741 B.n693 B.n692 10.6151
R742 B.n693 B.n6 10.6151
R743 B.n697 B.n6 10.6151
R744 B.n698 B.n697 10.6151
R745 B.n699 B.n698 10.6151
R746 B.n699 B.n4 10.6151
R747 B.n703 B.n4 10.6151
R748 B.n704 B.n703 10.6151
R749 B.n705 B.n704 10.6151
R750 B.n705 B.n0 10.6151
R751 B.n663 B.n662 10.6151
R752 B.n662 B.n661 10.6151
R753 B.n661 B.n18 10.6151
R754 B.n657 B.n18 10.6151
R755 B.n657 B.n656 10.6151
R756 B.n656 B.n655 10.6151
R757 B.n655 B.n20 10.6151
R758 B.n651 B.n20 10.6151
R759 B.n651 B.n650 10.6151
R760 B.n650 B.n649 10.6151
R761 B.n649 B.n22 10.6151
R762 B.n645 B.n22 10.6151
R763 B.n645 B.n644 10.6151
R764 B.n644 B.n643 10.6151
R765 B.n643 B.n24 10.6151
R766 B.n639 B.n24 10.6151
R767 B.n639 B.n638 10.6151
R768 B.n638 B.n637 10.6151
R769 B.n637 B.n26 10.6151
R770 B.n633 B.n26 10.6151
R771 B.n633 B.n632 10.6151
R772 B.n632 B.n631 10.6151
R773 B.n631 B.n28 10.6151
R774 B.n627 B.n28 10.6151
R775 B.n627 B.n626 10.6151
R776 B.n626 B.n625 10.6151
R777 B.n625 B.n30 10.6151
R778 B.n621 B.n30 10.6151
R779 B.n621 B.n620 10.6151
R780 B.n620 B.n619 10.6151
R781 B.n619 B.n32 10.6151
R782 B.n615 B.n32 10.6151
R783 B.n615 B.n614 10.6151
R784 B.n614 B.n613 10.6151
R785 B.n613 B.n34 10.6151
R786 B.n609 B.n34 10.6151
R787 B.n609 B.n608 10.6151
R788 B.n608 B.n607 10.6151
R789 B.n607 B.n36 10.6151
R790 B.n603 B.n36 10.6151
R791 B.n603 B.n602 10.6151
R792 B.n602 B.n601 10.6151
R793 B.n601 B.n38 10.6151
R794 B.n597 B.n38 10.6151
R795 B.n597 B.n596 10.6151
R796 B.n596 B.n595 10.6151
R797 B.n595 B.n40 10.6151
R798 B.n591 B.n40 10.6151
R799 B.n591 B.n590 10.6151
R800 B.n590 B.n589 10.6151
R801 B.n589 B.n42 10.6151
R802 B.n585 B.n42 10.6151
R803 B.n583 B.n582 10.6151
R804 B.n582 B.n46 10.6151
R805 B.n578 B.n46 10.6151
R806 B.n578 B.n577 10.6151
R807 B.n577 B.n576 10.6151
R808 B.n576 B.n48 10.6151
R809 B.n572 B.n48 10.6151
R810 B.n572 B.n571 10.6151
R811 B.n569 B.n52 10.6151
R812 B.n565 B.n52 10.6151
R813 B.n565 B.n564 10.6151
R814 B.n564 B.n563 10.6151
R815 B.n563 B.n54 10.6151
R816 B.n559 B.n54 10.6151
R817 B.n559 B.n558 10.6151
R818 B.n558 B.n557 10.6151
R819 B.n557 B.n56 10.6151
R820 B.n553 B.n56 10.6151
R821 B.n553 B.n552 10.6151
R822 B.n552 B.n551 10.6151
R823 B.n551 B.n58 10.6151
R824 B.n547 B.n58 10.6151
R825 B.n547 B.n546 10.6151
R826 B.n546 B.n545 10.6151
R827 B.n545 B.n60 10.6151
R828 B.n541 B.n60 10.6151
R829 B.n541 B.n540 10.6151
R830 B.n540 B.n539 10.6151
R831 B.n539 B.n62 10.6151
R832 B.n535 B.n62 10.6151
R833 B.n535 B.n534 10.6151
R834 B.n534 B.n533 10.6151
R835 B.n533 B.n64 10.6151
R836 B.n529 B.n64 10.6151
R837 B.n529 B.n528 10.6151
R838 B.n528 B.n527 10.6151
R839 B.n527 B.n66 10.6151
R840 B.n523 B.n66 10.6151
R841 B.n523 B.n522 10.6151
R842 B.n522 B.n521 10.6151
R843 B.n521 B.n68 10.6151
R844 B.n517 B.n68 10.6151
R845 B.n517 B.n516 10.6151
R846 B.n516 B.n515 10.6151
R847 B.n515 B.n70 10.6151
R848 B.n511 B.n70 10.6151
R849 B.n511 B.n510 10.6151
R850 B.n510 B.n509 10.6151
R851 B.n509 B.n72 10.6151
R852 B.n505 B.n72 10.6151
R853 B.n505 B.n504 10.6151
R854 B.n504 B.n503 10.6151
R855 B.n503 B.n74 10.6151
R856 B.n499 B.n74 10.6151
R857 B.n499 B.n498 10.6151
R858 B.n498 B.n497 10.6151
R859 B.n497 B.n76 10.6151
R860 B.n493 B.n76 10.6151
R861 B.n493 B.n492 10.6151
R862 B.n492 B.n491 10.6151
R863 B.n487 B.n78 10.6151
R864 B.n487 B.n486 10.6151
R865 B.n486 B.n485 10.6151
R866 B.n485 B.n80 10.6151
R867 B.n481 B.n80 10.6151
R868 B.n481 B.n480 10.6151
R869 B.n480 B.n479 10.6151
R870 B.n479 B.n82 10.6151
R871 B.n475 B.n82 10.6151
R872 B.n475 B.n474 10.6151
R873 B.n474 B.n473 10.6151
R874 B.n473 B.n84 10.6151
R875 B.n469 B.n84 10.6151
R876 B.n469 B.n468 10.6151
R877 B.n468 B.n467 10.6151
R878 B.n467 B.n86 10.6151
R879 B.n463 B.n86 10.6151
R880 B.n463 B.n462 10.6151
R881 B.n462 B.n461 10.6151
R882 B.n461 B.n88 10.6151
R883 B.n457 B.n88 10.6151
R884 B.n457 B.n456 10.6151
R885 B.n456 B.n455 10.6151
R886 B.n455 B.n90 10.6151
R887 B.n451 B.n90 10.6151
R888 B.n451 B.n450 10.6151
R889 B.n450 B.n449 10.6151
R890 B.n449 B.n92 10.6151
R891 B.n445 B.n92 10.6151
R892 B.n445 B.n444 10.6151
R893 B.n444 B.n443 10.6151
R894 B.n443 B.n94 10.6151
R895 B.n439 B.n94 10.6151
R896 B.n439 B.n438 10.6151
R897 B.n438 B.n437 10.6151
R898 B.n437 B.n96 10.6151
R899 B.n433 B.n96 10.6151
R900 B.n433 B.n432 10.6151
R901 B.n432 B.n431 10.6151
R902 B.n431 B.n98 10.6151
R903 B.n427 B.n98 10.6151
R904 B.n427 B.n426 10.6151
R905 B.n426 B.n425 10.6151
R906 B.n425 B.n100 10.6151
R907 B.n421 B.n100 10.6151
R908 B.n421 B.n420 10.6151
R909 B.n420 B.n419 10.6151
R910 B.n419 B.n102 10.6151
R911 B.n415 B.n102 10.6151
R912 B.n415 B.n414 10.6151
R913 B.n414 B.n413 10.6151
R914 B.n413 B.n104 10.6151
R915 B.n409 B.n104 10.6151
R916 B.n409 B.n408 10.6151
R917 B.n408 B.n407 10.6151
R918 B.n407 B.n106 10.6151
R919 B.n403 B.n106 10.6151
R920 B.n403 B.n402 10.6151
R921 B.n402 B.n401 10.6151
R922 B.n182 B.n1 10.6151
R923 B.n183 B.n182 10.6151
R924 B.n183 B.n180 10.6151
R925 B.n187 B.n180 10.6151
R926 B.n188 B.n187 10.6151
R927 B.n189 B.n188 10.6151
R928 B.n189 B.n178 10.6151
R929 B.n193 B.n178 10.6151
R930 B.n194 B.n193 10.6151
R931 B.n195 B.n194 10.6151
R932 B.n195 B.n176 10.6151
R933 B.n199 B.n176 10.6151
R934 B.n200 B.n199 10.6151
R935 B.n201 B.n200 10.6151
R936 B.n201 B.n174 10.6151
R937 B.n205 B.n174 10.6151
R938 B.n206 B.n205 10.6151
R939 B.n207 B.n206 10.6151
R940 B.n207 B.n172 10.6151
R941 B.n211 B.n172 10.6151
R942 B.n212 B.n211 10.6151
R943 B.n213 B.n212 10.6151
R944 B.n213 B.n170 10.6151
R945 B.n217 B.n170 10.6151
R946 B.n218 B.n217 10.6151
R947 B.n219 B.n218 10.6151
R948 B.n219 B.n168 10.6151
R949 B.n223 B.n168 10.6151
R950 B.n225 B.n224 10.6151
R951 B.n225 B.n166 10.6151
R952 B.n229 B.n166 10.6151
R953 B.n230 B.n229 10.6151
R954 B.n231 B.n230 10.6151
R955 B.n231 B.n164 10.6151
R956 B.n235 B.n164 10.6151
R957 B.n236 B.n235 10.6151
R958 B.n237 B.n236 10.6151
R959 B.n237 B.n162 10.6151
R960 B.n241 B.n162 10.6151
R961 B.n242 B.n241 10.6151
R962 B.n243 B.n242 10.6151
R963 B.n243 B.n160 10.6151
R964 B.n247 B.n160 10.6151
R965 B.n248 B.n247 10.6151
R966 B.n249 B.n248 10.6151
R967 B.n249 B.n158 10.6151
R968 B.n253 B.n158 10.6151
R969 B.n254 B.n253 10.6151
R970 B.n255 B.n254 10.6151
R971 B.n255 B.n156 10.6151
R972 B.n259 B.n156 10.6151
R973 B.n260 B.n259 10.6151
R974 B.n261 B.n260 10.6151
R975 B.n261 B.n154 10.6151
R976 B.n265 B.n154 10.6151
R977 B.n266 B.n265 10.6151
R978 B.n267 B.n266 10.6151
R979 B.n267 B.n152 10.6151
R980 B.n271 B.n152 10.6151
R981 B.n272 B.n271 10.6151
R982 B.n273 B.n272 10.6151
R983 B.n273 B.n150 10.6151
R984 B.n277 B.n150 10.6151
R985 B.n278 B.n277 10.6151
R986 B.n279 B.n278 10.6151
R987 B.n279 B.n148 10.6151
R988 B.n283 B.n148 10.6151
R989 B.n284 B.n283 10.6151
R990 B.n285 B.n284 10.6151
R991 B.n285 B.n146 10.6151
R992 B.n289 B.n146 10.6151
R993 B.n290 B.n289 10.6151
R994 B.n291 B.n290 10.6151
R995 B.n291 B.n144 10.6151
R996 B.n295 B.n144 10.6151
R997 B.n296 B.n295 10.6151
R998 B.n297 B.n296 10.6151
R999 B.n297 B.n142 10.6151
R1000 B.n301 B.n142 10.6151
R1001 B.n302 B.n301 10.6151
R1002 B.n304 B.n138 10.6151
R1003 B.n308 B.n138 10.6151
R1004 B.n309 B.n308 10.6151
R1005 B.n310 B.n309 10.6151
R1006 B.n310 B.n136 10.6151
R1007 B.n314 B.n136 10.6151
R1008 B.n315 B.n314 10.6151
R1009 B.n319 B.n315 10.6151
R1010 B.n323 B.n134 10.6151
R1011 B.n324 B.n323 10.6151
R1012 B.n325 B.n324 10.6151
R1013 B.n325 B.n132 10.6151
R1014 B.n329 B.n132 10.6151
R1015 B.n330 B.n329 10.6151
R1016 B.n331 B.n330 10.6151
R1017 B.n331 B.n130 10.6151
R1018 B.n335 B.n130 10.6151
R1019 B.n336 B.n335 10.6151
R1020 B.n337 B.n336 10.6151
R1021 B.n337 B.n128 10.6151
R1022 B.n341 B.n128 10.6151
R1023 B.n342 B.n341 10.6151
R1024 B.n343 B.n342 10.6151
R1025 B.n343 B.n126 10.6151
R1026 B.n347 B.n126 10.6151
R1027 B.n348 B.n347 10.6151
R1028 B.n349 B.n348 10.6151
R1029 B.n349 B.n124 10.6151
R1030 B.n353 B.n124 10.6151
R1031 B.n354 B.n353 10.6151
R1032 B.n355 B.n354 10.6151
R1033 B.n355 B.n122 10.6151
R1034 B.n359 B.n122 10.6151
R1035 B.n360 B.n359 10.6151
R1036 B.n361 B.n360 10.6151
R1037 B.n361 B.n120 10.6151
R1038 B.n365 B.n120 10.6151
R1039 B.n366 B.n365 10.6151
R1040 B.n367 B.n366 10.6151
R1041 B.n367 B.n118 10.6151
R1042 B.n371 B.n118 10.6151
R1043 B.n372 B.n371 10.6151
R1044 B.n373 B.n372 10.6151
R1045 B.n373 B.n116 10.6151
R1046 B.n377 B.n116 10.6151
R1047 B.n378 B.n377 10.6151
R1048 B.n379 B.n378 10.6151
R1049 B.n379 B.n114 10.6151
R1050 B.n383 B.n114 10.6151
R1051 B.n384 B.n383 10.6151
R1052 B.n385 B.n384 10.6151
R1053 B.n385 B.n112 10.6151
R1054 B.n389 B.n112 10.6151
R1055 B.n390 B.n389 10.6151
R1056 B.n391 B.n390 10.6151
R1057 B.n391 B.n110 10.6151
R1058 B.n395 B.n110 10.6151
R1059 B.n396 B.n395 10.6151
R1060 B.n397 B.n396 10.6151
R1061 B.n397 B.n108 10.6151
R1062 B.n709 B.n0 8.11757
R1063 B.n709 B.n1 8.11757
R1064 B.n584 B.n583 6.5566
R1065 B.n571 B.n570 6.5566
R1066 B.n304 B.n303 6.5566
R1067 B.n319 B.n318 6.5566
R1068 B.n585 B.n584 4.05904
R1069 B.n570 B.n569 4.05904
R1070 B.n303 B.n302 4.05904
R1071 B.n318 B.n134 4.05904
R1072 VP.n2 VP.t3 218.73
R1073 VP.n2 VP.t0 218.185
R1074 VP.n4 VP.t2 182.72
R1075 VP.n11 VP.t1 182.72
R1076 VP.n10 VP.n0 161.3
R1077 VP.n9 VP.n8 161.3
R1078 VP.n7 VP.n1 161.3
R1079 VP.n6 VP.n5 161.3
R1080 VP.n4 VP.n3 88.4915
R1081 VP.n12 VP.n11 88.4915
R1082 VP.n9 VP.n1 56.5193
R1083 VP.n3 VP.n2 54.5752
R1084 VP.n5 VP.n1 24.4675
R1085 VP.n10 VP.n9 24.4675
R1086 VP.n5 VP.n4 22.2655
R1087 VP.n11 VP.n10 22.2655
R1088 VP.n6 VP.n3 0.278367
R1089 VP.n12 VP.n0 0.278367
R1090 VP.n7 VP.n6 0.189894
R1091 VP.n8 VP.n7 0.189894
R1092 VP.n8 VP.n0 0.189894
R1093 VP VP.n12 0.153454
R1094 VTAIL.n5 VTAIL.t7 56.3758
R1095 VTAIL.n4 VTAIL.t2 56.3758
R1096 VTAIL.n3 VTAIL.t3 56.3758
R1097 VTAIL.n6 VTAIL.t6 56.3757
R1098 VTAIL.n7 VTAIL.t0 56.3757
R1099 VTAIL.n0 VTAIL.t1 56.3757
R1100 VTAIL.n1 VTAIL.t4 56.3757
R1101 VTAIL.n2 VTAIL.t5 56.3757
R1102 VTAIL.n7 VTAIL.n6 28.0393
R1103 VTAIL.n3 VTAIL.n2 28.0393
R1104 VTAIL.n4 VTAIL.n3 2.07809
R1105 VTAIL.n6 VTAIL.n5 2.07809
R1106 VTAIL.n2 VTAIL.n1 2.07809
R1107 VTAIL VTAIL.n0 1.09748
R1108 VTAIL VTAIL.n7 0.981103
R1109 VTAIL.n5 VTAIL.n4 0.470328
R1110 VTAIL.n1 VTAIL.n0 0.470328
R1111 VDD1 VDD1.n1 115.061
R1112 VDD1 VDD1.n0 71.0515
R1113 VDD1.n0 VDD1.t0 2.06169
R1114 VDD1.n0 VDD1.t3 2.06169
R1115 VDD1.n1 VDD1.t1 2.06169
R1116 VDD1.n1 VDD1.t2 2.06169
R1117 VN.n0 VN.t0 218.73
R1118 VN.n1 VN.t1 218.73
R1119 VN.n0 VN.t2 218.185
R1120 VN.n1 VN.t3 218.185
R1121 VN VN.n1 54.8541
R1122 VN VN.n0 6.97905
R1123 VDD2.n2 VDD2.n0 114.535
R1124 VDD2.n2 VDD2.n1 70.9933
R1125 VDD2.n1 VDD2.t0 2.06169
R1126 VDD2.n1 VDD2.t2 2.06169
R1127 VDD2.n0 VDD2.t3 2.06169
R1128 VDD2.n0 VDD2.t1 2.06169
R1129 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 5.55487f
C1 B VTAIL 5.89219f
C2 VP w_n2416_n4122# 4.37034f
C3 VP VDD1 6.08415f
C4 B VN 1.05432f
C5 VDD2 VTAIL 6.40692f
C6 VDD2 VN 5.87207f
C7 w_n2416_n4122# VTAIL 4.83584f
C8 B VDD2 1.31632f
C9 VTAIL VDD1 6.3562f
C10 w_n2416_n4122# VN 4.06107f
C11 VN VDD1 0.148657f
C12 w_n2416_n4122# B 9.663219f
C13 B VDD1 1.2727f
C14 VP VTAIL 5.56898f
C15 w_n2416_n4122# VDD2 1.49988f
C16 VDD2 VDD1 0.903829f
C17 VP VN 6.51306f
C18 VP B 1.56512f
C19 w_n2416_n4122# VDD1 1.45539f
C20 VP VDD2 0.361344f
C21 VDD2 VSUBS 0.949729f
C22 VDD1 VSUBS 5.94616f
C23 VTAIL VSUBS 1.335473f
C24 VN VSUBS 5.41004f
C25 VP VSUBS 2.160237f
C26 B VSUBS 4.141731f
C27 w_n2416_n4122# VSUBS 0.122027p
C28 VDD2.t3 VSUBS 0.331183f
C29 VDD2.t1 VSUBS 0.331183f
C30 VDD2.n0 VSUBS 3.53206f
C31 VDD2.t0 VSUBS 0.331183f
C32 VDD2.t2 VSUBS 0.331183f
C33 VDD2.n1 VSUBS 2.70906f
C34 VDD2.n2 VSUBS 4.55052f
C35 VN.t0 VSUBS 3.36135f
C36 VN.t2 VSUBS 3.35814f
C37 VN.n0 VSUBS 2.25926f
C38 VN.t1 VSUBS 3.36135f
C39 VN.t3 VSUBS 3.35814f
C40 VN.n1 VSUBS 4.05555f
C41 VDD1.t0 VSUBS 0.333903f
C42 VDD1.t3 VSUBS 0.333903f
C43 VDD1.n0 VSUBS 2.7319f
C44 VDD1.t1 VSUBS 0.333903f
C45 VDD1.t2 VSUBS 0.333903f
C46 VDD1.n1 VSUBS 3.5876f
C47 VTAIL.t1 VSUBS 2.82351f
C48 VTAIL.n0 VSUBS 0.740849f
C49 VTAIL.t4 VSUBS 2.82351f
C50 VTAIL.n1 VSUBS 0.811772f
C51 VTAIL.t5 VSUBS 2.82351f
C52 VTAIL.n2 VSUBS 2.21621f
C53 VTAIL.t3 VSUBS 2.82353f
C54 VTAIL.n3 VSUBS 2.21619f
C55 VTAIL.t2 VSUBS 2.82353f
C56 VTAIL.n4 VSUBS 0.81175f
C57 VTAIL.t7 VSUBS 2.82353f
C58 VTAIL.n5 VSUBS 0.81175f
C59 VTAIL.t6 VSUBS 2.82351f
C60 VTAIL.n6 VSUBS 2.21621f
C61 VTAIL.t0 VSUBS 2.82351f
C62 VTAIL.n7 VSUBS 2.13687f
C63 VP.n0 VSUBS 0.047267f
C64 VP.t1 VSUBS 3.22602f
C65 VP.n1 VSUBS 0.052337f
C66 VP.t0 VSUBS 3.44177f
C67 VP.t3 VSUBS 3.44506f
C68 VP.n2 VSUBS 4.13823f
C69 VP.n3 VSUBS 2.13431f
C70 VP.t2 VSUBS 3.22602f
C71 VP.n4 VSUBS 1.25137f
C72 VP.n5 VSUBS 0.063848f
C73 VP.n6 VSUBS 0.047267f
C74 VP.n7 VSUBS 0.035852f
C75 VP.n8 VSUBS 0.035852f
C76 VP.n9 VSUBS 0.052337f
C77 VP.n10 VSUBS 0.063848f
C78 VP.n11 VSUBS 1.25137f
C79 VP.n12 VSUBS 0.041149f
C80 B.n0 VSUBS 0.005828f
C81 B.n1 VSUBS 0.005828f
C82 B.n2 VSUBS 0.00862f
C83 B.n3 VSUBS 0.006606f
C84 B.n4 VSUBS 0.006606f
C85 B.n5 VSUBS 0.006606f
C86 B.n6 VSUBS 0.006606f
C87 B.n7 VSUBS 0.006606f
C88 B.n8 VSUBS 0.006606f
C89 B.n9 VSUBS 0.006606f
C90 B.n10 VSUBS 0.006606f
C91 B.n11 VSUBS 0.006606f
C92 B.n12 VSUBS 0.006606f
C93 B.n13 VSUBS 0.006606f
C94 B.n14 VSUBS 0.006606f
C95 B.n15 VSUBS 0.006606f
C96 B.n16 VSUBS 0.014649f
C97 B.n17 VSUBS 0.006606f
C98 B.n18 VSUBS 0.006606f
C99 B.n19 VSUBS 0.006606f
C100 B.n20 VSUBS 0.006606f
C101 B.n21 VSUBS 0.006606f
C102 B.n22 VSUBS 0.006606f
C103 B.n23 VSUBS 0.006606f
C104 B.n24 VSUBS 0.006606f
C105 B.n25 VSUBS 0.006606f
C106 B.n26 VSUBS 0.006606f
C107 B.n27 VSUBS 0.006606f
C108 B.n28 VSUBS 0.006606f
C109 B.n29 VSUBS 0.006606f
C110 B.n30 VSUBS 0.006606f
C111 B.n31 VSUBS 0.006606f
C112 B.n32 VSUBS 0.006606f
C113 B.n33 VSUBS 0.006606f
C114 B.n34 VSUBS 0.006606f
C115 B.n35 VSUBS 0.006606f
C116 B.n36 VSUBS 0.006606f
C117 B.n37 VSUBS 0.006606f
C118 B.n38 VSUBS 0.006606f
C119 B.n39 VSUBS 0.006606f
C120 B.n40 VSUBS 0.006606f
C121 B.n41 VSUBS 0.006606f
C122 B.n42 VSUBS 0.006606f
C123 B.n43 VSUBS 0.006606f
C124 B.t1 VSUBS 0.497441f
C125 B.t2 VSUBS 0.514404f
C126 B.t0 VSUBS 1.36242f
C127 B.n44 VSUBS 0.255456f
C128 B.n45 VSUBS 0.065928f
C129 B.n46 VSUBS 0.006606f
C130 B.n47 VSUBS 0.006606f
C131 B.n48 VSUBS 0.006606f
C132 B.n49 VSUBS 0.006606f
C133 B.t10 VSUBS 0.497425f
C134 B.t11 VSUBS 0.514391f
C135 B.t9 VSUBS 1.36242f
C136 B.n50 VSUBS 0.255468f
C137 B.n51 VSUBS 0.065943f
C138 B.n52 VSUBS 0.006606f
C139 B.n53 VSUBS 0.006606f
C140 B.n54 VSUBS 0.006606f
C141 B.n55 VSUBS 0.006606f
C142 B.n56 VSUBS 0.006606f
C143 B.n57 VSUBS 0.006606f
C144 B.n58 VSUBS 0.006606f
C145 B.n59 VSUBS 0.006606f
C146 B.n60 VSUBS 0.006606f
C147 B.n61 VSUBS 0.006606f
C148 B.n62 VSUBS 0.006606f
C149 B.n63 VSUBS 0.006606f
C150 B.n64 VSUBS 0.006606f
C151 B.n65 VSUBS 0.006606f
C152 B.n66 VSUBS 0.006606f
C153 B.n67 VSUBS 0.006606f
C154 B.n68 VSUBS 0.006606f
C155 B.n69 VSUBS 0.006606f
C156 B.n70 VSUBS 0.006606f
C157 B.n71 VSUBS 0.006606f
C158 B.n72 VSUBS 0.006606f
C159 B.n73 VSUBS 0.006606f
C160 B.n74 VSUBS 0.006606f
C161 B.n75 VSUBS 0.006606f
C162 B.n76 VSUBS 0.006606f
C163 B.n77 VSUBS 0.006606f
C164 B.n78 VSUBS 0.014649f
C165 B.n79 VSUBS 0.006606f
C166 B.n80 VSUBS 0.006606f
C167 B.n81 VSUBS 0.006606f
C168 B.n82 VSUBS 0.006606f
C169 B.n83 VSUBS 0.006606f
C170 B.n84 VSUBS 0.006606f
C171 B.n85 VSUBS 0.006606f
C172 B.n86 VSUBS 0.006606f
C173 B.n87 VSUBS 0.006606f
C174 B.n88 VSUBS 0.006606f
C175 B.n89 VSUBS 0.006606f
C176 B.n90 VSUBS 0.006606f
C177 B.n91 VSUBS 0.006606f
C178 B.n92 VSUBS 0.006606f
C179 B.n93 VSUBS 0.006606f
C180 B.n94 VSUBS 0.006606f
C181 B.n95 VSUBS 0.006606f
C182 B.n96 VSUBS 0.006606f
C183 B.n97 VSUBS 0.006606f
C184 B.n98 VSUBS 0.006606f
C185 B.n99 VSUBS 0.006606f
C186 B.n100 VSUBS 0.006606f
C187 B.n101 VSUBS 0.006606f
C188 B.n102 VSUBS 0.006606f
C189 B.n103 VSUBS 0.006606f
C190 B.n104 VSUBS 0.006606f
C191 B.n105 VSUBS 0.006606f
C192 B.n106 VSUBS 0.006606f
C193 B.n107 VSUBS 0.006606f
C194 B.n108 VSUBS 0.014449f
C195 B.n109 VSUBS 0.006606f
C196 B.n110 VSUBS 0.006606f
C197 B.n111 VSUBS 0.006606f
C198 B.n112 VSUBS 0.006606f
C199 B.n113 VSUBS 0.006606f
C200 B.n114 VSUBS 0.006606f
C201 B.n115 VSUBS 0.006606f
C202 B.n116 VSUBS 0.006606f
C203 B.n117 VSUBS 0.006606f
C204 B.n118 VSUBS 0.006606f
C205 B.n119 VSUBS 0.006606f
C206 B.n120 VSUBS 0.006606f
C207 B.n121 VSUBS 0.006606f
C208 B.n122 VSUBS 0.006606f
C209 B.n123 VSUBS 0.006606f
C210 B.n124 VSUBS 0.006606f
C211 B.n125 VSUBS 0.006606f
C212 B.n126 VSUBS 0.006606f
C213 B.n127 VSUBS 0.006606f
C214 B.n128 VSUBS 0.006606f
C215 B.n129 VSUBS 0.006606f
C216 B.n130 VSUBS 0.006606f
C217 B.n131 VSUBS 0.006606f
C218 B.n132 VSUBS 0.006606f
C219 B.n133 VSUBS 0.006606f
C220 B.n134 VSUBS 0.004566f
C221 B.n135 VSUBS 0.006606f
C222 B.n136 VSUBS 0.006606f
C223 B.n137 VSUBS 0.006606f
C224 B.n138 VSUBS 0.006606f
C225 B.n139 VSUBS 0.006606f
C226 B.t5 VSUBS 0.497441f
C227 B.t4 VSUBS 0.514404f
C228 B.t3 VSUBS 1.36242f
C229 B.n140 VSUBS 0.255456f
C230 B.n141 VSUBS 0.065928f
C231 B.n142 VSUBS 0.006606f
C232 B.n143 VSUBS 0.006606f
C233 B.n144 VSUBS 0.006606f
C234 B.n145 VSUBS 0.006606f
C235 B.n146 VSUBS 0.006606f
C236 B.n147 VSUBS 0.006606f
C237 B.n148 VSUBS 0.006606f
C238 B.n149 VSUBS 0.006606f
C239 B.n150 VSUBS 0.006606f
C240 B.n151 VSUBS 0.006606f
C241 B.n152 VSUBS 0.006606f
C242 B.n153 VSUBS 0.006606f
C243 B.n154 VSUBS 0.006606f
C244 B.n155 VSUBS 0.006606f
C245 B.n156 VSUBS 0.006606f
C246 B.n157 VSUBS 0.006606f
C247 B.n158 VSUBS 0.006606f
C248 B.n159 VSUBS 0.006606f
C249 B.n160 VSUBS 0.006606f
C250 B.n161 VSUBS 0.006606f
C251 B.n162 VSUBS 0.006606f
C252 B.n163 VSUBS 0.006606f
C253 B.n164 VSUBS 0.006606f
C254 B.n165 VSUBS 0.006606f
C255 B.n166 VSUBS 0.006606f
C256 B.n167 VSUBS 0.01527f
C257 B.n168 VSUBS 0.006606f
C258 B.n169 VSUBS 0.006606f
C259 B.n170 VSUBS 0.006606f
C260 B.n171 VSUBS 0.006606f
C261 B.n172 VSUBS 0.006606f
C262 B.n173 VSUBS 0.006606f
C263 B.n174 VSUBS 0.006606f
C264 B.n175 VSUBS 0.006606f
C265 B.n176 VSUBS 0.006606f
C266 B.n177 VSUBS 0.006606f
C267 B.n178 VSUBS 0.006606f
C268 B.n179 VSUBS 0.006606f
C269 B.n180 VSUBS 0.006606f
C270 B.n181 VSUBS 0.006606f
C271 B.n182 VSUBS 0.006606f
C272 B.n183 VSUBS 0.006606f
C273 B.n184 VSUBS 0.006606f
C274 B.n185 VSUBS 0.006606f
C275 B.n186 VSUBS 0.006606f
C276 B.n187 VSUBS 0.006606f
C277 B.n188 VSUBS 0.006606f
C278 B.n189 VSUBS 0.006606f
C279 B.n190 VSUBS 0.006606f
C280 B.n191 VSUBS 0.006606f
C281 B.n192 VSUBS 0.006606f
C282 B.n193 VSUBS 0.006606f
C283 B.n194 VSUBS 0.006606f
C284 B.n195 VSUBS 0.006606f
C285 B.n196 VSUBS 0.006606f
C286 B.n197 VSUBS 0.006606f
C287 B.n198 VSUBS 0.006606f
C288 B.n199 VSUBS 0.006606f
C289 B.n200 VSUBS 0.006606f
C290 B.n201 VSUBS 0.006606f
C291 B.n202 VSUBS 0.006606f
C292 B.n203 VSUBS 0.006606f
C293 B.n204 VSUBS 0.006606f
C294 B.n205 VSUBS 0.006606f
C295 B.n206 VSUBS 0.006606f
C296 B.n207 VSUBS 0.006606f
C297 B.n208 VSUBS 0.006606f
C298 B.n209 VSUBS 0.006606f
C299 B.n210 VSUBS 0.006606f
C300 B.n211 VSUBS 0.006606f
C301 B.n212 VSUBS 0.006606f
C302 B.n213 VSUBS 0.006606f
C303 B.n214 VSUBS 0.006606f
C304 B.n215 VSUBS 0.006606f
C305 B.n216 VSUBS 0.006606f
C306 B.n217 VSUBS 0.006606f
C307 B.n218 VSUBS 0.006606f
C308 B.n219 VSUBS 0.006606f
C309 B.n220 VSUBS 0.006606f
C310 B.n221 VSUBS 0.006606f
C311 B.n222 VSUBS 0.014649f
C312 B.n223 VSUBS 0.014649f
C313 B.n224 VSUBS 0.01527f
C314 B.n225 VSUBS 0.006606f
C315 B.n226 VSUBS 0.006606f
C316 B.n227 VSUBS 0.006606f
C317 B.n228 VSUBS 0.006606f
C318 B.n229 VSUBS 0.006606f
C319 B.n230 VSUBS 0.006606f
C320 B.n231 VSUBS 0.006606f
C321 B.n232 VSUBS 0.006606f
C322 B.n233 VSUBS 0.006606f
C323 B.n234 VSUBS 0.006606f
C324 B.n235 VSUBS 0.006606f
C325 B.n236 VSUBS 0.006606f
C326 B.n237 VSUBS 0.006606f
C327 B.n238 VSUBS 0.006606f
C328 B.n239 VSUBS 0.006606f
C329 B.n240 VSUBS 0.006606f
C330 B.n241 VSUBS 0.006606f
C331 B.n242 VSUBS 0.006606f
C332 B.n243 VSUBS 0.006606f
C333 B.n244 VSUBS 0.006606f
C334 B.n245 VSUBS 0.006606f
C335 B.n246 VSUBS 0.006606f
C336 B.n247 VSUBS 0.006606f
C337 B.n248 VSUBS 0.006606f
C338 B.n249 VSUBS 0.006606f
C339 B.n250 VSUBS 0.006606f
C340 B.n251 VSUBS 0.006606f
C341 B.n252 VSUBS 0.006606f
C342 B.n253 VSUBS 0.006606f
C343 B.n254 VSUBS 0.006606f
C344 B.n255 VSUBS 0.006606f
C345 B.n256 VSUBS 0.006606f
C346 B.n257 VSUBS 0.006606f
C347 B.n258 VSUBS 0.006606f
C348 B.n259 VSUBS 0.006606f
C349 B.n260 VSUBS 0.006606f
C350 B.n261 VSUBS 0.006606f
C351 B.n262 VSUBS 0.006606f
C352 B.n263 VSUBS 0.006606f
C353 B.n264 VSUBS 0.006606f
C354 B.n265 VSUBS 0.006606f
C355 B.n266 VSUBS 0.006606f
C356 B.n267 VSUBS 0.006606f
C357 B.n268 VSUBS 0.006606f
C358 B.n269 VSUBS 0.006606f
C359 B.n270 VSUBS 0.006606f
C360 B.n271 VSUBS 0.006606f
C361 B.n272 VSUBS 0.006606f
C362 B.n273 VSUBS 0.006606f
C363 B.n274 VSUBS 0.006606f
C364 B.n275 VSUBS 0.006606f
C365 B.n276 VSUBS 0.006606f
C366 B.n277 VSUBS 0.006606f
C367 B.n278 VSUBS 0.006606f
C368 B.n279 VSUBS 0.006606f
C369 B.n280 VSUBS 0.006606f
C370 B.n281 VSUBS 0.006606f
C371 B.n282 VSUBS 0.006606f
C372 B.n283 VSUBS 0.006606f
C373 B.n284 VSUBS 0.006606f
C374 B.n285 VSUBS 0.006606f
C375 B.n286 VSUBS 0.006606f
C376 B.n287 VSUBS 0.006606f
C377 B.n288 VSUBS 0.006606f
C378 B.n289 VSUBS 0.006606f
C379 B.n290 VSUBS 0.006606f
C380 B.n291 VSUBS 0.006606f
C381 B.n292 VSUBS 0.006606f
C382 B.n293 VSUBS 0.006606f
C383 B.n294 VSUBS 0.006606f
C384 B.n295 VSUBS 0.006606f
C385 B.n296 VSUBS 0.006606f
C386 B.n297 VSUBS 0.006606f
C387 B.n298 VSUBS 0.006606f
C388 B.n299 VSUBS 0.006606f
C389 B.n300 VSUBS 0.006606f
C390 B.n301 VSUBS 0.006606f
C391 B.n302 VSUBS 0.004566f
C392 B.n303 VSUBS 0.015304f
C393 B.n304 VSUBS 0.005343f
C394 B.n305 VSUBS 0.006606f
C395 B.n306 VSUBS 0.006606f
C396 B.n307 VSUBS 0.006606f
C397 B.n308 VSUBS 0.006606f
C398 B.n309 VSUBS 0.006606f
C399 B.n310 VSUBS 0.006606f
C400 B.n311 VSUBS 0.006606f
C401 B.n312 VSUBS 0.006606f
C402 B.n313 VSUBS 0.006606f
C403 B.n314 VSUBS 0.006606f
C404 B.n315 VSUBS 0.006606f
C405 B.t8 VSUBS 0.497425f
C406 B.t7 VSUBS 0.514391f
C407 B.t6 VSUBS 1.36242f
C408 B.n316 VSUBS 0.255468f
C409 B.n317 VSUBS 0.065943f
C410 B.n318 VSUBS 0.015304f
C411 B.n319 VSUBS 0.005343f
C412 B.n320 VSUBS 0.006606f
C413 B.n321 VSUBS 0.006606f
C414 B.n322 VSUBS 0.006606f
C415 B.n323 VSUBS 0.006606f
C416 B.n324 VSUBS 0.006606f
C417 B.n325 VSUBS 0.006606f
C418 B.n326 VSUBS 0.006606f
C419 B.n327 VSUBS 0.006606f
C420 B.n328 VSUBS 0.006606f
C421 B.n329 VSUBS 0.006606f
C422 B.n330 VSUBS 0.006606f
C423 B.n331 VSUBS 0.006606f
C424 B.n332 VSUBS 0.006606f
C425 B.n333 VSUBS 0.006606f
C426 B.n334 VSUBS 0.006606f
C427 B.n335 VSUBS 0.006606f
C428 B.n336 VSUBS 0.006606f
C429 B.n337 VSUBS 0.006606f
C430 B.n338 VSUBS 0.006606f
C431 B.n339 VSUBS 0.006606f
C432 B.n340 VSUBS 0.006606f
C433 B.n341 VSUBS 0.006606f
C434 B.n342 VSUBS 0.006606f
C435 B.n343 VSUBS 0.006606f
C436 B.n344 VSUBS 0.006606f
C437 B.n345 VSUBS 0.006606f
C438 B.n346 VSUBS 0.006606f
C439 B.n347 VSUBS 0.006606f
C440 B.n348 VSUBS 0.006606f
C441 B.n349 VSUBS 0.006606f
C442 B.n350 VSUBS 0.006606f
C443 B.n351 VSUBS 0.006606f
C444 B.n352 VSUBS 0.006606f
C445 B.n353 VSUBS 0.006606f
C446 B.n354 VSUBS 0.006606f
C447 B.n355 VSUBS 0.006606f
C448 B.n356 VSUBS 0.006606f
C449 B.n357 VSUBS 0.006606f
C450 B.n358 VSUBS 0.006606f
C451 B.n359 VSUBS 0.006606f
C452 B.n360 VSUBS 0.006606f
C453 B.n361 VSUBS 0.006606f
C454 B.n362 VSUBS 0.006606f
C455 B.n363 VSUBS 0.006606f
C456 B.n364 VSUBS 0.006606f
C457 B.n365 VSUBS 0.006606f
C458 B.n366 VSUBS 0.006606f
C459 B.n367 VSUBS 0.006606f
C460 B.n368 VSUBS 0.006606f
C461 B.n369 VSUBS 0.006606f
C462 B.n370 VSUBS 0.006606f
C463 B.n371 VSUBS 0.006606f
C464 B.n372 VSUBS 0.006606f
C465 B.n373 VSUBS 0.006606f
C466 B.n374 VSUBS 0.006606f
C467 B.n375 VSUBS 0.006606f
C468 B.n376 VSUBS 0.006606f
C469 B.n377 VSUBS 0.006606f
C470 B.n378 VSUBS 0.006606f
C471 B.n379 VSUBS 0.006606f
C472 B.n380 VSUBS 0.006606f
C473 B.n381 VSUBS 0.006606f
C474 B.n382 VSUBS 0.006606f
C475 B.n383 VSUBS 0.006606f
C476 B.n384 VSUBS 0.006606f
C477 B.n385 VSUBS 0.006606f
C478 B.n386 VSUBS 0.006606f
C479 B.n387 VSUBS 0.006606f
C480 B.n388 VSUBS 0.006606f
C481 B.n389 VSUBS 0.006606f
C482 B.n390 VSUBS 0.006606f
C483 B.n391 VSUBS 0.006606f
C484 B.n392 VSUBS 0.006606f
C485 B.n393 VSUBS 0.006606f
C486 B.n394 VSUBS 0.006606f
C487 B.n395 VSUBS 0.006606f
C488 B.n396 VSUBS 0.006606f
C489 B.n397 VSUBS 0.006606f
C490 B.n398 VSUBS 0.006606f
C491 B.n399 VSUBS 0.01527f
C492 B.n400 VSUBS 0.014649f
C493 B.n401 VSUBS 0.01547f
C494 B.n402 VSUBS 0.006606f
C495 B.n403 VSUBS 0.006606f
C496 B.n404 VSUBS 0.006606f
C497 B.n405 VSUBS 0.006606f
C498 B.n406 VSUBS 0.006606f
C499 B.n407 VSUBS 0.006606f
C500 B.n408 VSUBS 0.006606f
C501 B.n409 VSUBS 0.006606f
C502 B.n410 VSUBS 0.006606f
C503 B.n411 VSUBS 0.006606f
C504 B.n412 VSUBS 0.006606f
C505 B.n413 VSUBS 0.006606f
C506 B.n414 VSUBS 0.006606f
C507 B.n415 VSUBS 0.006606f
C508 B.n416 VSUBS 0.006606f
C509 B.n417 VSUBS 0.006606f
C510 B.n418 VSUBS 0.006606f
C511 B.n419 VSUBS 0.006606f
C512 B.n420 VSUBS 0.006606f
C513 B.n421 VSUBS 0.006606f
C514 B.n422 VSUBS 0.006606f
C515 B.n423 VSUBS 0.006606f
C516 B.n424 VSUBS 0.006606f
C517 B.n425 VSUBS 0.006606f
C518 B.n426 VSUBS 0.006606f
C519 B.n427 VSUBS 0.006606f
C520 B.n428 VSUBS 0.006606f
C521 B.n429 VSUBS 0.006606f
C522 B.n430 VSUBS 0.006606f
C523 B.n431 VSUBS 0.006606f
C524 B.n432 VSUBS 0.006606f
C525 B.n433 VSUBS 0.006606f
C526 B.n434 VSUBS 0.006606f
C527 B.n435 VSUBS 0.006606f
C528 B.n436 VSUBS 0.006606f
C529 B.n437 VSUBS 0.006606f
C530 B.n438 VSUBS 0.006606f
C531 B.n439 VSUBS 0.006606f
C532 B.n440 VSUBS 0.006606f
C533 B.n441 VSUBS 0.006606f
C534 B.n442 VSUBS 0.006606f
C535 B.n443 VSUBS 0.006606f
C536 B.n444 VSUBS 0.006606f
C537 B.n445 VSUBS 0.006606f
C538 B.n446 VSUBS 0.006606f
C539 B.n447 VSUBS 0.006606f
C540 B.n448 VSUBS 0.006606f
C541 B.n449 VSUBS 0.006606f
C542 B.n450 VSUBS 0.006606f
C543 B.n451 VSUBS 0.006606f
C544 B.n452 VSUBS 0.006606f
C545 B.n453 VSUBS 0.006606f
C546 B.n454 VSUBS 0.006606f
C547 B.n455 VSUBS 0.006606f
C548 B.n456 VSUBS 0.006606f
C549 B.n457 VSUBS 0.006606f
C550 B.n458 VSUBS 0.006606f
C551 B.n459 VSUBS 0.006606f
C552 B.n460 VSUBS 0.006606f
C553 B.n461 VSUBS 0.006606f
C554 B.n462 VSUBS 0.006606f
C555 B.n463 VSUBS 0.006606f
C556 B.n464 VSUBS 0.006606f
C557 B.n465 VSUBS 0.006606f
C558 B.n466 VSUBS 0.006606f
C559 B.n467 VSUBS 0.006606f
C560 B.n468 VSUBS 0.006606f
C561 B.n469 VSUBS 0.006606f
C562 B.n470 VSUBS 0.006606f
C563 B.n471 VSUBS 0.006606f
C564 B.n472 VSUBS 0.006606f
C565 B.n473 VSUBS 0.006606f
C566 B.n474 VSUBS 0.006606f
C567 B.n475 VSUBS 0.006606f
C568 B.n476 VSUBS 0.006606f
C569 B.n477 VSUBS 0.006606f
C570 B.n478 VSUBS 0.006606f
C571 B.n479 VSUBS 0.006606f
C572 B.n480 VSUBS 0.006606f
C573 B.n481 VSUBS 0.006606f
C574 B.n482 VSUBS 0.006606f
C575 B.n483 VSUBS 0.006606f
C576 B.n484 VSUBS 0.006606f
C577 B.n485 VSUBS 0.006606f
C578 B.n486 VSUBS 0.006606f
C579 B.n487 VSUBS 0.006606f
C580 B.n488 VSUBS 0.006606f
C581 B.n489 VSUBS 0.014649f
C582 B.n490 VSUBS 0.01527f
C583 B.n491 VSUBS 0.01527f
C584 B.n492 VSUBS 0.006606f
C585 B.n493 VSUBS 0.006606f
C586 B.n494 VSUBS 0.006606f
C587 B.n495 VSUBS 0.006606f
C588 B.n496 VSUBS 0.006606f
C589 B.n497 VSUBS 0.006606f
C590 B.n498 VSUBS 0.006606f
C591 B.n499 VSUBS 0.006606f
C592 B.n500 VSUBS 0.006606f
C593 B.n501 VSUBS 0.006606f
C594 B.n502 VSUBS 0.006606f
C595 B.n503 VSUBS 0.006606f
C596 B.n504 VSUBS 0.006606f
C597 B.n505 VSUBS 0.006606f
C598 B.n506 VSUBS 0.006606f
C599 B.n507 VSUBS 0.006606f
C600 B.n508 VSUBS 0.006606f
C601 B.n509 VSUBS 0.006606f
C602 B.n510 VSUBS 0.006606f
C603 B.n511 VSUBS 0.006606f
C604 B.n512 VSUBS 0.006606f
C605 B.n513 VSUBS 0.006606f
C606 B.n514 VSUBS 0.006606f
C607 B.n515 VSUBS 0.006606f
C608 B.n516 VSUBS 0.006606f
C609 B.n517 VSUBS 0.006606f
C610 B.n518 VSUBS 0.006606f
C611 B.n519 VSUBS 0.006606f
C612 B.n520 VSUBS 0.006606f
C613 B.n521 VSUBS 0.006606f
C614 B.n522 VSUBS 0.006606f
C615 B.n523 VSUBS 0.006606f
C616 B.n524 VSUBS 0.006606f
C617 B.n525 VSUBS 0.006606f
C618 B.n526 VSUBS 0.006606f
C619 B.n527 VSUBS 0.006606f
C620 B.n528 VSUBS 0.006606f
C621 B.n529 VSUBS 0.006606f
C622 B.n530 VSUBS 0.006606f
C623 B.n531 VSUBS 0.006606f
C624 B.n532 VSUBS 0.006606f
C625 B.n533 VSUBS 0.006606f
C626 B.n534 VSUBS 0.006606f
C627 B.n535 VSUBS 0.006606f
C628 B.n536 VSUBS 0.006606f
C629 B.n537 VSUBS 0.006606f
C630 B.n538 VSUBS 0.006606f
C631 B.n539 VSUBS 0.006606f
C632 B.n540 VSUBS 0.006606f
C633 B.n541 VSUBS 0.006606f
C634 B.n542 VSUBS 0.006606f
C635 B.n543 VSUBS 0.006606f
C636 B.n544 VSUBS 0.006606f
C637 B.n545 VSUBS 0.006606f
C638 B.n546 VSUBS 0.006606f
C639 B.n547 VSUBS 0.006606f
C640 B.n548 VSUBS 0.006606f
C641 B.n549 VSUBS 0.006606f
C642 B.n550 VSUBS 0.006606f
C643 B.n551 VSUBS 0.006606f
C644 B.n552 VSUBS 0.006606f
C645 B.n553 VSUBS 0.006606f
C646 B.n554 VSUBS 0.006606f
C647 B.n555 VSUBS 0.006606f
C648 B.n556 VSUBS 0.006606f
C649 B.n557 VSUBS 0.006606f
C650 B.n558 VSUBS 0.006606f
C651 B.n559 VSUBS 0.006606f
C652 B.n560 VSUBS 0.006606f
C653 B.n561 VSUBS 0.006606f
C654 B.n562 VSUBS 0.006606f
C655 B.n563 VSUBS 0.006606f
C656 B.n564 VSUBS 0.006606f
C657 B.n565 VSUBS 0.006606f
C658 B.n566 VSUBS 0.006606f
C659 B.n567 VSUBS 0.006606f
C660 B.n568 VSUBS 0.006606f
C661 B.n569 VSUBS 0.004566f
C662 B.n570 VSUBS 0.015304f
C663 B.n571 VSUBS 0.005343f
C664 B.n572 VSUBS 0.006606f
C665 B.n573 VSUBS 0.006606f
C666 B.n574 VSUBS 0.006606f
C667 B.n575 VSUBS 0.006606f
C668 B.n576 VSUBS 0.006606f
C669 B.n577 VSUBS 0.006606f
C670 B.n578 VSUBS 0.006606f
C671 B.n579 VSUBS 0.006606f
C672 B.n580 VSUBS 0.006606f
C673 B.n581 VSUBS 0.006606f
C674 B.n582 VSUBS 0.006606f
C675 B.n583 VSUBS 0.005343f
C676 B.n584 VSUBS 0.015304f
C677 B.n585 VSUBS 0.004566f
C678 B.n586 VSUBS 0.006606f
C679 B.n587 VSUBS 0.006606f
C680 B.n588 VSUBS 0.006606f
C681 B.n589 VSUBS 0.006606f
C682 B.n590 VSUBS 0.006606f
C683 B.n591 VSUBS 0.006606f
C684 B.n592 VSUBS 0.006606f
C685 B.n593 VSUBS 0.006606f
C686 B.n594 VSUBS 0.006606f
C687 B.n595 VSUBS 0.006606f
C688 B.n596 VSUBS 0.006606f
C689 B.n597 VSUBS 0.006606f
C690 B.n598 VSUBS 0.006606f
C691 B.n599 VSUBS 0.006606f
C692 B.n600 VSUBS 0.006606f
C693 B.n601 VSUBS 0.006606f
C694 B.n602 VSUBS 0.006606f
C695 B.n603 VSUBS 0.006606f
C696 B.n604 VSUBS 0.006606f
C697 B.n605 VSUBS 0.006606f
C698 B.n606 VSUBS 0.006606f
C699 B.n607 VSUBS 0.006606f
C700 B.n608 VSUBS 0.006606f
C701 B.n609 VSUBS 0.006606f
C702 B.n610 VSUBS 0.006606f
C703 B.n611 VSUBS 0.006606f
C704 B.n612 VSUBS 0.006606f
C705 B.n613 VSUBS 0.006606f
C706 B.n614 VSUBS 0.006606f
C707 B.n615 VSUBS 0.006606f
C708 B.n616 VSUBS 0.006606f
C709 B.n617 VSUBS 0.006606f
C710 B.n618 VSUBS 0.006606f
C711 B.n619 VSUBS 0.006606f
C712 B.n620 VSUBS 0.006606f
C713 B.n621 VSUBS 0.006606f
C714 B.n622 VSUBS 0.006606f
C715 B.n623 VSUBS 0.006606f
C716 B.n624 VSUBS 0.006606f
C717 B.n625 VSUBS 0.006606f
C718 B.n626 VSUBS 0.006606f
C719 B.n627 VSUBS 0.006606f
C720 B.n628 VSUBS 0.006606f
C721 B.n629 VSUBS 0.006606f
C722 B.n630 VSUBS 0.006606f
C723 B.n631 VSUBS 0.006606f
C724 B.n632 VSUBS 0.006606f
C725 B.n633 VSUBS 0.006606f
C726 B.n634 VSUBS 0.006606f
C727 B.n635 VSUBS 0.006606f
C728 B.n636 VSUBS 0.006606f
C729 B.n637 VSUBS 0.006606f
C730 B.n638 VSUBS 0.006606f
C731 B.n639 VSUBS 0.006606f
C732 B.n640 VSUBS 0.006606f
C733 B.n641 VSUBS 0.006606f
C734 B.n642 VSUBS 0.006606f
C735 B.n643 VSUBS 0.006606f
C736 B.n644 VSUBS 0.006606f
C737 B.n645 VSUBS 0.006606f
C738 B.n646 VSUBS 0.006606f
C739 B.n647 VSUBS 0.006606f
C740 B.n648 VSUBS 0.006606f
C741 B.n649 VSUBS 0.006606f
C742 B.n650 VSUBS 0.006606f
C743 B.n651 VSUBS 0.006606f
C744 B.n652 VSUBS 0.006606f
C745 B.n653 VSUBS 0.006606f
C746 B.n654 VSUBS 0.006606f
C747 B.n655 VSUBS 0.006606f
C748 B.n656 VSUBS 0.006606f
C749 B.n657 VSUBS 0.006606f
C750 B.n658 VSUBS 0.006606f
C751 B.n659 VSUBS 0.006606f
C752 B.n660 VSUBS 0.006606f
C753 B.n661 VSUBS 0.006606f
C754 B.n662 VSUBS 0.006606f
C755 B.n663 VSUBS 0.01527f
C756 B.n664 VSUBS 0.01527f
C757 B.n665 VSUBS 0.014649f
C758 B.n666 VSUBS 0.006606f
C759 B.n667 VSUBS 0.006606f
C760 B.n668 VSUBS 0.006606f
C761 B.n669 VSUBS 0.006606f
C762 B.n670 VSUBS 0.006606f
C763 B.n671 VSUBS 0.006606f
C764 B.n672 VSUBS 0.006606f
C765 B.n673 VSUBS 0.006606f
C766 B.n674 VSUBS 0.006606f
C767 B.n675 VSUBS 0.006606f
C768 B.n676 VSUBS 0.006606f
C769 B.n677 VSUBS 0.006606f
C770 B.n678 VSUBS 0.006606f
C771 B.n679 VSUBS 0.006606f
C772 B.n680 VSUBS 0.006606f
C773 B.n681 VSUBS 0.006606f
C774 B.n682 VSUBS 0.006606f
C775 B.n683 VSUBS 0.006606f
C776 B.n684 VSUBS 0.006606f
C777 B.n685 VSUBS 0.006606f
C778 B.n686 VSUBS 0.006606f
C779 B.n687 VSUBS 0.006606f
C780 B.n688 VSUBS 0.006606f
C781 B.n689 VSUBS 0.006606f
C782 B.n690 VSUBS 0.006606f
C783 B.n691 VSUBS 0.006606f
C784 B.n692 VSUBS 0.006606f
C785 B.n693 VSUBS 0.006606f
C786 B.n694 VSUBS 0.006606f
C787 B.n695 VSUBS 0.006606f
C788 B.n696 VSUBS 0.006606f
C789 B.n697 VSUBS 0.006606f
C790 B.n698 VSUBS 0.006606f
C791 B.n699 VSUBS 0.006606f
C792 B.n700 VSUBS 0.006606f
C793 B.n701 VSUBS 0.006606f
C794 B.n702 VSUBS 0.006606f
C795 B.n703 VSUBS 0.006606f
C796 B.n704 VSUBS 0.006606f
C797 B.n705 VSUBS 0.006606f
C798 B.n706 VSUBS 0.006606f
C799 B.n707 VSUBS 0.00862f
C800 B.n708 VSUBS 0.009182f
C801 B.n709 VSUBS 0.01826f
.ends

