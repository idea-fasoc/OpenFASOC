* NGSPICE file created from diff_pair_sample_1311.ext - technology: sky130A

.subckt diff_pair_sample_1311 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.32
X1 VDD1.t3 VP.t0 VTAIL.t5 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.32
X2 VTAIL.t4 VP.t1 VDD1.t2 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.32
X3 B.t8 B.t6 B.t7 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.32
X4 B.t5 B.t3 B.t4 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.32
X5 B.t2 B.t0 B.t1 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.32
X6 VTAIL.t2 VN.t0 VDD2.t3 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.32
X7 VDD1.t1 VP.t2 VTAIL.t7 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.32
X8 VTAIL.t0 VN.t1 VDD2.t2 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.32
X9 VDD2.t1 VN.t2 VTAIL.t3 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.32
X10 VDD2.t0 VN.t3 VTAIL.t1 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.32
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n1360_n4668# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.32
R0 B.n124 B.t6 1605.53
R1 B.n132 B.t3 1605.53
R2 B.n40 B.t0 1605.53
R3 B.n46 B.t9 1605.53
R4 B.n432 B.n431 585
R5 B.n433 B.n78 585
R6 B.n435 B.n434 585
R7 B.n436 B.n77 585
R8 B.n438 B.n437 585
R9 B.n439 B.n76 585
R10 B.n441 B.n440 585
R11 B.n442 B.n75 585
R12 B.n444 B.n443 585
R13 B.n445 B.n74 585
R14 B.n447 B.n446 585
R15 B.n448 B.n73 585
R16 B.n450 B.n449 585
R17 B.n451 B.n72 585
R18 B.n453 B.n452 585
R19 B.n454 B.n71 585
R20 B.n456 B.n455 585
R21 B.n457 B.n70 585
R22 B.n459 B.n458 585
R23 B.n460 B.n69 585
R24 B.n462 B.n461 585
R25 B.n463 B.n68 585
R26 B.n465 B.n464 585
R27 B.n466 B.n67 585
R28 B.n468 B.n467 585
R29 B.n469 B.n66 585
R30 B.n471 B.n470 585
R31 B.n472 B.n65 585
R32 B.n474 B.n473 585
R33 B.n475 B.n64 585
R34 B.n477 B.n476 585
R35 B.n478 B.n63 585
R36 B.n480 B.n479 585
R37 B.n481 B.n62 585
R38 B.n483 B.n482 585
R39 B.n484 B.n61 585
R40 B.n486 B.n485 585
R41 B.n487 B.n60 585
R42 B.n489 B.n488 585
R43 B.n490 B.n59 585
R44 B.n492 B.n491 585
R45 B.n493 B.n58 585
R46 B.n495 B.n494 585
R47 B.n496 B.n57 585
R48 B.n498 B.n497 585
R49 B.n499 B.n56 585
R50 B.n501 B.n500 585
R51 B.n502 B.n55 585
R52 B.n504 B.n503 585
R53 B.n505 B.n54 585
R54 B.n507 B.n506 585
R55 B.n508 B.n53 585
R56 B.n510 B.n509 585
R57 B.n511 B.n52 585
R58 B.n513 B.n512 585
R59 B.n514 B.n51 585
R60 B.n516 B.n515 585
R61 B.n517 B.n50 585
R62 B.n519 B.n518 585
R63 B.n520 B.n49 585
R64 B.n522 B.n521 585
R65 B.n524 B.n523 585
R66 B.n525 B.n45 585
R67 B.n527 B.n526 585
R68 B.n528 B.n44 585
R69 B.n530 B.n529 585
R70 B.n531 B.n43 585
R71 B.n533 B.n532 585
R72 B.n534 B.n42 585
R73 B.n536 B.n535 585
R74 B.n538 B.n39 585
R75 B.n540 B.n539 585
R76 B.n541 B.n38 585
R77 B.n543 B.n542 585
R78 B.n544 B.n37 585
R79 B.n546 B.n545 585
R80 B.n547 B.n36 585
R81 B.n549 B.n548 585
R82 B.n550 B.n35 585
R83 B.n552 B.n551 585
R84 B.n553 B.n34 585
R85 B.n555 B.n554 585
R86 B.n556 B.n33 585
R87 B.n558 B.n557 585
R88 B.n559 B.n32 585
R89 B.n561 B.n560 585
R90 B.n562 B.n31 585
R91 B.n564 B.n563 585
R92 B.n565 B.n30 585
R93 B.n567 B.n566 585
R94 B.n568 B.n29 585
R95 B.n570 B.n569 585
R96 B.n571 B.n28 585
R97 B.n573 B.n572 585
R98 B.n574 B.n27 585
R99 B.n576 B.n575 585
R100 B.n577 B.n26 585
R101 B.n579 B.n578 585
R102 B.n580 B.n25 585
R103 B.n582 B.n581 585
R104 B.n583 B.n24 585
R105 B.n585 B.n584 585
R106 B.n586 B.n23 585
R107 B.n588 B.n587 585
R108 B.n589 B.n22 585
R109 B.n591 B.n590 585
R110 B.n592 B.n21 585
R111 B.n594 B.n593 585
R112 B.n595 B.n20 585
R113 B.n597 B.n596 585
R114 B.n598 B.n19 585
R115 B.n600 B.n599 585
R116 B.n601 B.n18 585
R117 B.n603 B.n602 585
R118 B.n604 B.n17 585
R119 B.n606 B.n605 585
R120 B.n607 B.n16 585
R121 B.n609 B.n608 585
R122 B.n610 B.n15 585
R123 B.n612 B.n611 585
R124 B.n613 B.n14 585
R125 B.n615 B.n614 585
R126 B.n616 B.n13 585
R127 B.n618 B.n617 585
R128 B.n619 B.n12 585
R129 B.n621 B.n620 585
R130 B.n622 B.n11 585
R131 B.n624 B.n623 585
R132 B.n625 B.n10 585
R133 B.n627 B.n626 585
R134 B.n628 B.n9 585
R135 B.n430 B.n79 585
R136 B.n429 B.n428 585
R137 B.n427 B.n80 585
R138 B.n426 B.n425 585
R139 B.n424 B.n81 585
R140 B.n423 B.n422 585
R141 B.n421 B.n82 585
R142 B.n420 B.n419 585
R143 B.n418 B.n83 585
R144 B.n417 B.n416 585
R145 B.n415 B.n84 585
R146 B.n414 B.n413 585
R147 B.n412 B.n85 585
R148 B.n411 B.n410 585
R149 B.n409 B.n86 585
R150 B.n408 B.n407 585
R151 B.n406 B.n87 585
R152 B.n405 B.n404 585
R153 B.n403 B.n88 585
R154 B.n402 B.n401 585
R155 B.n400 B.n89 585
R156 B.n399 B.n398 585
R157 B.n397 B.n90 585
R158 B.n396 B.n395 585
R159 B.n394 B.n91 585
R160 B.n393 B.n392 585
R161 B.n391 B.n92 585
R162 B.n390 B.n389 585
R163 B.n388 B.n93 585
R164 B.n190 B.n163 585
R165 B.n192 B.n191 585
R166 B.n193 B.n162 585
R167 B.n195 B.n194 585
R168 B.n196 B.n161 585
R169 B.n198 B.n197 585
R170 B.n199 B.n160 585
R171 B.n201 B.n200 585
R172 B.n202 B.n159 585
R173 B.n204 B.n203 585
R174 B.n205 B.n158 585
R175 B.n207 B.n206 585
R176 B.n208 B.n157 585
R177 B.n210 B.n209 585
R178 B.n211 B.n156 585
R179 B.n213 B.n212 585
R180 B.n214 B.n155 585
R181 B.n216 B.n215 585
R182 B.n217 B.n154 585
R183 B.n219 B.n218 585
R184 B.n220 B.n153 585
R185 B.n222 B.n221 585
R186 B.n223 B.n152 585
R187 B.n225 B.n224 585
R188 B.n226 B.n151 585
R189 B.n228 B.n227 585
R190 B.n229 B.n150 585
R191 B.n231 B.n230 585
R192 B.n232 B.n149 585
R193 B.n234 B.n233 585
R194 B.n235 B.n148 585
R195 B.n237 B.n236 585
R196 B.n238 B.n147 585
R197 B.n240 B.n239 585
R198 B.n241 B.n146 585
R199 B.n243 B.n242 585
R200 B.n244 B.n145 585
R201 B.n246 B.n245 585
R202 B.n247 B.n144 585
R203 B.n249 B.n248 585
R204 B.n250 B.n143 585
R205 B.n252 B.n251 585
R206 B.n253 B.n142 585
R207 B.n255 B.n254 585
R208 B.n256 B.n141 585
R209 B.n258 B.n257 585
R210 B.n259 B.n140 585
R211 B.n261 B.n260 585
R212 B.n262 B.n139 585
R213 B.n264 B.n263 585
R214 B.n265 B.n138 585
R215 B.n267 B.n266 585
R216 B.n268 B.n137 585
R217 B.n270 B.n269 585
R218 B.n271 B.n136 585
R219 B.n273 B.n272 585
R220 B.n274 B.n135 585
R221 B.n276 B.n275 585
R222 B.n277 B.n134 585
R223 B.n279 B.n278 585
R224 B.n280 B.n131 585
R225 B.n283 B.n282 585
R226 B.n284 B.n130 585
R227 B.n286 B.n285 585
R228 B.n287 B.n129 585
R229 B.n289 B.n288 585
R230 B.n290 B.n128 585
R231 B.n292 B.n291 585
R232 B.n293 B.n127 585
R233 B.n295 B.n294 585
R234 B.n297 B.n296 585
R235 B.n298 B.n123 585
R236 B.n300 B.n299 585
R237 B.n301 B.n122 585
R238 B.n303 B.n302 585
R239 B.n304 B.n121 585
R240 B.n306 B.n305 585
R241 B.n307 B.n120 585
R242 B.n309 B.n308 585
R243 B.n310 B.n119 585
R244 B.n312 B.n311 585
R245 B.n313 B.n118 585
R246 B.n315 B.n314 585
R247 B.n316 B.n117 585
R248 B.n318 B.n317 585
R249 B.n319 B.n116 585
R250 B.n321 B.n320 585
R251 B.n322 B.n115 585
R252 B.n324 B.n323 585
R253 B.n325 B.n114 585
R254 B.n327 B.n326 585
R255 B.n328 B.n113 585
R256 B.n330 B.n329 585
R257 B.n331 B.n112 585
R258 B.n333 B.n332 585
R259 B.n334 B.n111 585
R260 B.n336 B.n335 585
R261 B.n337 B.n110 585
R262 B.n339 B.n338 585
R263 B.n340 B.n109 585
R264 B.n342 B.n341 585
R265 B.n343 B.n108 585
R266 B.n345 B.n344 585
R267 B.n346 B.n107 585
R268 B.n348 B.n347 585
R269 B.n349 B.n106 585
R270 B.n351 B.n350 585
R271 B.n352 B.n105 585
R272 B.n354 B.n353 585
R273 B.n355 B.n104 585
R274 B.n357 B.n356 585
R275 B.n358 B.n103 585
R276 B.n360 B.n359 585
R277 B.n361 B.n102 585
R278 B.n363 B.n362 585
R279 B.n364 B.n101 585
R280 B.n366 B.n365 585
R281 B.n367 B.n100 585
R282 B.n369 B.n368 585
R283 B.n370 B.n99 585
R284 B.n372 B.n371 585
R285 B.n373 B.n98 585
R286 B.n375 B.n374 585
R287 B.n376 B.n97 585
R288 B.n378 B.n377 585
R289 B.n379 B.n96 585
R290 B.n381 B.n380 585
R291 B.n382 B.n95 585
R292 B.n384 B.n383 585
R293 B.n385 B.n94 585
R294 B.n387 B.n386 585
R295 B.n189 B.n188 585
R296 B.n187 B.n164 585
R297 B.n186 B.n185 585
R298 B.n184 B.n165 585
R299 B.n183 B.n182 585
R300 B.n181 B.n166 585
R301 B.n180 B.n179 585
R302 B.n178 B.n167 585
R303 B.n177 B.n176 585
R304 B.n175 B.n168 585
R305 B.n174 B.n173 585
R306 B.n172 B.n169 585
R307 B.n171 B.n170 585
R308 B.n2 B.n0 585
R309 B.n649 B.n1 585
R310 B.n648 B.n647 585
R311 B.n646 B.n3 585
R312 B.n645 B.n644 585
R313 B.n643 B.n4 585
R314 B.n642 B.n641 585
R315 B.n640 B.n5 585
R316 B.n639 B.n638 585
R317 B.n637 B.n6 585
R318 B.n636 B.n635 585
R319 B.n634 B.n7 585
R320 B.n633 B.n632 585
R321 B.n631 B.n8 585
R322 B.n630 B.n629 585
R323 B.n651 B.n650 585
R324 B.n188 B.n163 478.086
R325 B.n630 B.n9 478.086
R326 B.n386 B.n93 478.086
R327 B.n432 B.n79 478.086
R328 B.n188 B.n187 163.367
R329 B.n187 B.n186 163.367
R330 B.n186 B.n165 163.367
R331 B.n182 B.n165 163.367
R332 B.n182 B.n181 163.367
R333 B.n181 B.n180 163.367
R334 B.n180 B.n167 163.367
R335 B.n176 B.n167 163.367
R336 B.n176 B.n175 163.367
R337 B.n175 B.n174 163.367
R338 B.n174 B.n169 163.367
R339 B.n170 B.n169 163.367
R340 B.n170 B.n2 163.367
R341 B.n650 B.n2 163.367
R342 B.n650 B.n649 163.367
R343 B.n649 B.n648 163.367
R344 B.n648 B.n3 163.367
R345 B.n644 B.n3 163.367
R346 B.n644 B.n643 163.367
R347 B.n643 B.n642 163.367
R348 B.n642 B.n5 163.367
R349 B.n638 B.n5 163.367
R350 B.n638 B.n637 163.367
R351 B.n637 B.n636 163.367
R352 B.n636 B.n7 163.367
R353 B.n632 B.n7 163.367
R354 B.n632 B.n631 163.367
R355 B.n631 B.n630 163.367
R356 B.n192 B.n163 163.367
R357 B.n193 B.n192 163.367
R358 B.n194 B.n193 163.367
R359 B.n194 B.n161 163.367
R360 B.n198 B.n161 163.367
R361 B.n199 B.n198 163.367
R362 B.n200 B.n199 163.367
R363 B.n200 B.n159 163.367
R364 B.n204 B.n159 163.367
R365 B.n205 B.n204 163.367
R366 B.n206 B.n205 163.367
R367 B.n206 B.n157 163.367
R368 B.n210 B.n157 163.367
R369 B.n211 B.n210 163.367
R370 B.n212 B.n211 163.367
R371 B.n212 B.n155 163.367
R372 B.n216 B.n155 163.367
R373 B.n217 B.n216 163.367
R374 B.n218 B.n217 163.367
R375 B.n218 B.n153 163.367
R376 B.n222 B.n153 163.367
R377 B.n223 B.n222 163.367
R378 B.n224 B.n223 163.367
R379 B.n224 B.n151 163.367
R380 B.n228 B.n151 163.367
R381 B.n229 B.n228 163.367
R382 B.n230 B.n229 163.367
R383 B.n230 B.n149 163.367
R384 B.n234 B.n149 163.367
R385 B.n235 B.n234 163.367
R386 B.n236 B.n235 163.367
R387 B.n236 B.n147 163.367
R388 B.n240 B.n147 163.367
R389 B.n241 B.n240 163.367
R390 B.n242 B.n241 163.367
R391 B.n242 B.n145 163.367
R392 B.n246 B.n145 163.367
R393 B.n247 B.n246 163.367
R394 B.n248 B.n247 163.367
R395 B.n248 B.n143 163.367
R396 B.n252 B.n143 163.367
R397 B.n253 B.n252 163.367
R398 B.n254 B.n253 163.367
R399 B.n254 B.n141 163.367
R400 B.n258 B.n141 163.367
R401 B.n259 B.n258 163.367
R402 B.n260 B.n259 163.367
R403 B.n260 B.n139 163.367
R404 B.n264 B.n139 163.367
R405 B.n265 B.n264 163.367
R406 B.n266 B.n265 163.367
R407 B.n266 B.n137 163.367
R408 B.n270 B.n137 163.367
R409 B.n271 B.n270 163.367
R410 B.n272 B.n271 163.367
R411 B.n272 B.n135 163.367
R412 B.n276 B.n135 163.367
R413 B.n277 B.n276 163.367
R414 B.n278 B.n277 163.367
R415 B.n278 B.n131 163.367
R416 B.n283 B.n131 163.367
R417 B.n284 B.n283 163.367
R418 B.n285 B.n284 163.367
R419 B.n285 B.n129 163.367
R420 B.n289 B.n129 163.367
R421 B.n290 B.n289 163.367
R422 B.n291 B.n290 163.367
R423 B.n291 B.n127 163.367
R424 B.n295 B.n127 163.367
R425 B.n296 B.n295 163.367
R426 B.n296 B.n123 163.367
R427 B.n300 B.n123 163.367
R428 B.n301 B.n300 163.367
R429 B.n302 B.n301 163.367
R430 B.n302 B.n121 163.367
R431 B.n306 B.n121 163.367
R432 B.n307 B.n306 163.367
R433 B.n308 B.n307 163.367
R434 B.n308 B.n119 163.367
R435 B.n312 B.n119 163.367
R436 B.n313 B.n312 163.367
R437 B.n314 B.n313 163.367
R438 B.n314 B.n117 163.367
R439 B.n318 B.n117 163.367
R440 B.n319 B.n318 163.367
R441 B.n320 B.n319 163.367
R442 B.n320 B.n115 163.367
R443 B.n324 B.n115 163.367
R444 B.n325 B.n324 163.367
R445 B.n326 B.n325 163.367
R446 B.n326 B.n113 163.367
R447 B.n330 B.n113 163.367
R448 B.n331 B.n330 163.367
R449 B.n332 B.n331 163.367
R450 B.n332 B.n111 163.367
R451 B.n336 B.n111 163.367
R452 B.n337 B.n336 163.367
R453 B.n338 B.n337 163.367
R454 B.n338 B.n109 163.367
R455 B.n342 B.n109 163.367
R456 B.n343 B.n342 163.367
R457 B.n344 B.n343 163.367
R458 B.n344 B.n107 163.367
R459 B.n348 B.n107 163.367
R460 B.n349 B.n348 163.367
R461 B.n350 B.n349 163.367
R462 B.n350 B.n105 163.367
R463 B.n354 B.n105 163.367
R464 B.n355 B.n354 163.367
R465 B.n356 B.n355 163.367
R466 B.n356 B.n103 163.367
R467 B.n360 B.n103 163.367
R468 B.n361 B.n360 163.367
R469 B.n362 B.n361 163.367
R470 B.n362 B.n101 163.367
R471 B.n366 B.n101 163.367
R472 B.n367 B.n366 163.367
R473 B.n368 B.n367 163.367
R474 B.n368 B.n99 163.367
R475 B.n372 B.n99 163.367
R476 B.n373 B.n372 163.367
R477 B.n374 B.n373 163.367
R478 B.n374 B.n97 163.367
R479 B.n378 B.n97 163.367
R480 B.n379 B.n378 163.367
R481 B.n380 B.n379 163.367
R482 B.n380 B.n95 163.367
R483 B.n384 B.n95 163.367
R484 B.n385 B.n384 163.367
R485 B.n386 B.n385 163.367
R486 B.n390 B.n93 163.367
R487 B.n391 B.n390 163.367
R488 B.n392 B.n391 163.367
R489 B.n392 B.n91 163.367
R490 B.n396 B.n91 163.367
R491 B.n397 B.n396 163.367
R492 B.n398 B.n397 163.367
R493 B.n398 B.n89 163.367
R494 B.n402 B.n89 163.367
R495 B.n403 B.n402 163.367
R496 B.n404 B.n403 163.367
R497 B.n404 B.n87 163.367
R498 B.n408 B.n87 163.367
R499 B.n409 B.n408 163.367
R500 B.n410 B.n409 163.367
R501 B.n410 B.n85 163.367
R502 B.n414 B.n85 163.367
R503 B.n415 B.n414 163.367
R504 B.n416 B.n415 163.367
R505 B.n416 B.n83 163.367
R506 B.n420 B.n83 163.367
R507 B.n421 B.n420 163.367
R508 B.n422 B.n421 163.367
R509 B.n422 B.n81 163.367
R510 B.n426 B.n81 163.367
R511 B.n427 B.n426 163.367
R512 B.n428 B.n427 163.367
R513 B.n428 B.n79 163.367
R514 B.n626 B.n9 163.367
R515 B.n626 B.n625 163.367
R516 B.n625 B.n624 163.367
R517 B.n624 B.n11 163.367
R518 B.n620 B.n11 163.367
R519 B.n620 B.n619 163.367
R520 B.n619 B.n618 163.367
R521 B.n618 B.n13 163.367
R522 B.n614 B.n13 163.367
R523 B.n614 B.n613 163.367
R524 B.n613 B.n612 163.367
R525 B.n612 B.n15 163.367
R526 B.n608 B.n15 163.367
R527 B.n608 B.n607 163.367
R528 B.n607 B.n606 163.367
R529 B.n606 B.n17 163.367
R530 B.n602 B.n17 163.367
R531 B.n602 B.n601 163.367
R532 B.n601 B.n600 163.367
R533 B.n600 B.n19 163.367
R534 B.n596 B.n19 163.367
R535 B.n596 B.n595 163.367
R536 B.n595 B.n594 163.367
R537 B.n594 B.n21 163.367
R538 B.n590 B.n21 163.367
R539 B.n590 B.n589 163.367
R540 B.n589 B.n588 163.367
R541 B.n588 B.n23 163.367
R542 B.n584 B.n23 163.367
R543 B.n584 B.n583 163.367
R544 B.n583 B.n582 163.367
R545 B.n582 B.n25 163.367
R546 B.n578 B.n25 163.367
R547 B.n578 B.n577 163.367
R548 B.n577 B.n576 163.367
R549 B.n576 B.n27 163.367
R550 B.n572 B.n27 163.367
R551 B.n572 B.n571 163.367
R552 B.n571 B.n570 163.367
R553 B.n570 B.n29 163.367
R554 B.n566 B.n29 163.367
R555 B.n566 B.n565 163.367
R556 B.n565 B.n564 163.367
R557 B.n564 B.n31 163.367
R558 B.n560 B.n31 163.367
R559 B.n560 B.n559 163.367
R560 B.n559 B.n558 163.367
R561 B.n558 B.n33 163.367
R562 B.n554 B.n33 163.367
R563 B.n554 B.n553 163.367
R564 B.n553 B.n552 163.367
R565 B.n552 B.n35 163.367
R566 B.n548 B.n35 163.367
R567 B.n548 B.n547 163.367
R568 B.n547 B.n546 163.367
R569 B.n546 B.n37 163.367
R570 B.n542 B.n37 163.367
R571 B.n542 B.n541 163.367
R572 B.n541 B.n540 163.367
R573 B.n540 B.n39 163.367
R574 B.n535 B.n39 163.367
R575 B.n535 B.n534 163.367
R576 B.n534 B.n533 163.367
R577 B.n533 B.n43 163.367
R578 B.n529 B.n43 163.367
R579 B.n529 B.n528 163.367
R580 B.n528 B.n527 163.367
R581 B.n527 B.n45 163.367
R582 B.n523 B.n45 163.367
R583 B.n523 B.n522 163.367
R584 B.n522 B.n49 163.367
R585 B.n518 B.n49 163.367
R586 B.n518 B.n517 163.367
R587 B.n517 B.n516 163.367
R588 B.n516 B.n51 163.367
R589 B.n512 B.n51 163.367
R590 B.n512 B.n511 163.367
R591 B.n511 B.n510 163.367
R592 B.n510 B.n53 163.367
R593 B.n506 B.n53 163.367
R594 B.n506 B.n505 163.367
R595 B.n505 B.n504 163.367
R596 B.n504 B.n55 163.367
R597 B.n500 B.n55 163.367
R598 B.n500 B.n499 163.367
R599 B.n499 B.n498 163.367
R600 B.n498 B.n57 163.367
R601 B.n494 B.n57 163.367
R602 B.n494 B.n493 163.367
R603 B.n493 B.n492 163.367
R604 B.n492 B.n59 163.367
R605 B.n488 B.n59 163.367
R606 B.n488 B.n487 163.367
R607 B.n487 B.n486 163.367
R608 B.n486 B.n61 163.367
R609 B.n482 B.n61 163.367
R610 B.n482 B.n481 163.367
R611 B.n481 B.n480 163.367
R612 B.n480 B.n63 163.367
R613 B.n476 B.n63 163.367
R614 B.n476 B.n475 163.367
R615 B.n475 B.n474 163.367
R616 B.n474 B.n65 163.367
R617 B.n470 B.n65 163.367
R618 B.n470 B.n469 163.367
R619 B.n469 B.n468 163.367
R620 B.n468 B.n67 163.367
R621 B.n464 B.n67 163.367
R622 B.n464 B.n463 163.367
R623 B.n463 B.n462 163.367
R624 B.n462 B.n69 163.367
R625 B.n458 B.n69 163.367
R626 B.n458 B.n457 163.367
R627 B.n457 B.n456 163.367
R628 B.n456 B.n71 163.367
R629 B.n452 B.n71 163.367
R630 B.n452 B.n451 163.367
R631 B.n451 B.n450 163.367
R632 B.n450 B.n73 163.367
R633 B.n446 B.n73 163.367
R634 B.n446 B.n445 163.367
R635 B.n445 B.n444 163.367
R636 B.n444 B.n75 163.367
R637 B.n440 B.n75 163.367
R638 B.n440 B.n439 163.367
R639 B.n439 B.n438 163.367
R640 B.n438 B.n77 163.367
R641 B.n434 B.n77 163.367
R642 B.n434 B.n433 163.367
R643 B.n433 B.n432 163.367
R644 B.n124 B.t8 121.091
R645 B.n46 B.t10 121.091
R646 B.n132 B.t5 121.067
R647 B.n40 B.t1 121.067
R648 B.n125 B.t7 108.486
R649 B.n47 B.t11 108.486
R650 B.n133 B.t4 108.462
R651 B.n41 B.t2 108.462
R652 B.n126 B.n125 59.5399
R653 B.n281 B.n133 59.5399
R654 B.n537 B.n41 59.5399
R655 B.n48 B.n47 59.5399
R656 B.n629 B.n628 31.0639
R657 B.n431 B.n430 31.0639
R658 B.n388 B.n387 31.0639
R659 B.n190 B.n189 31.0639
R660 B B.n651 18.0485
R661 B.n125 B.n124 12.6066
R662 B.n133 B.n132 12.6066
R663 B.n41 B.n40 12.6066
R664 B.n47 B.n46 12.6066
R665 B.n628 B.n627 10.6151
R666 B.n627 B.n10 10.6151
R667 B.n623 B.n10 10.6151
R668 B.n623 B.n622 10.6151
R669 B.n622 B.n621 10.6151
R670 B.n621 B.n12 10.6151
R671 B.n617 B.n12 10.6151
R672 B.n617 B.n616 10.6151
R673 B.n616 B.n615 10.6151
R674 B.n615 B.n14 10.6151
R675 B.n611 B.n14 10.6151
R676 B.n611 B.n610 10.6151
R677 B.n610 B.n609 10.6151
R678 B.n609 B.n16 10.6151
R679 B.n605 B.n16 10.6151
R680 B.n605 B.n604 10.6151
R681 B.n604 B.n603 10.6151
R682 B.n603 B.n18 10.6151
R683 B.n599 B.n18 10.6151
R684 B.n599 B.n598 10.6151
R685 B.n598 B.n597 10.6151
R686 B.n597 B.n20 10.6151
R687 B.n593 B.n20 10.6151
R688 B.n593 B.n592 10.6151
R689 B.n592 B.n591 10.6151
R690 B.n591 B.n22 10.6151
R691 B.n587 B.n22 10.6151
R692 B.n587 B.n586 10.6151
R693 B.n586 B.n585 10.6151
R694 B.n585 B.n24 10.6151
R695 B.n581 B.n24 10.6151
R696 B.n581 B.n580 10.6151
R697 B.n580 B.n579 10.6151
R698 B.n579 B.n26 10.6151
R699 B.n575 B.n26 10.6151
R700 B.n575 B.n574 10.6151
R701 B.n574 B.n573 10.6151
R702 B.n573 B.n28 10.6151
R703 B.n569 B.n28 10.6151
R704 B.n569 B.n568 10.6151
R705 B.n568 B.n567 10.6151
R706 B.n567 B.n30 10.6151
R707 B.n563 B.n30 10.6151
R708 B.n563 B.n562 10.6151
R709 B.n562 B.n561 10.6151
R710 B.n561 B.n32 10.6151
R711 B.n557 B.n32 10.6151
R712 B.n557 B.n556 10.6151
R713 B.n556 B.n555 10.6151
R714 B.n555 B.n34 10.6151
R715 B.n551 B.n34 10.6151
R716 B.n551 B.n550 10.6151
R717 B.n550 B.n549 10.6151
R718 B.n549 B.n36 10.6151
R719 B.n545 B.n36 10.6151
R720 B.n545 B.n544 10.6151
R721 B.n544 B.n543 10.6151
R722 B.n543 B.n38 10.6151
R723 B.n539 B.n38 10.6151
R724 B.n539 B.n538 10.6151
R725 B.n536 B.n42 10.6151
R726 B.n532 B.n42 10.6151
R727 B.n532 B.n531 10.6151
R728 B.n531 B.n530 10.6151
R729 B.n530 B.n44 10.6151
R730 B.n526 B.n44 10.6151
R731 B.n526 B.n525 10.6151
R732 B.n525 B.n524 10.6151
R733 B.n521 B.n520 10.6151
R734 B.n520 B.n519 10.6151
R735 B.n519 B.n50 10.6151
R736 B.n515 B.n50 10.6151
R737 B.n515 B.n514 10.6151
R738 B.n514 B.n513 10.6151
R739 B.n513 B.n52 10.6151
R740 B.n509 B.n52 10.6151
R741 B.n509 B.n508 10.6151
R742 B.n508 B.n507 10.6151
R743 B.n507 B.n54 10.6151
R744 B.n503 B.n54 10.6151
R745 B.n503 B.n502 10.6151
R746 B.n502 B.n501 10.6151
R747 B.n501 B.n56 10.6151
R748 B.n497 B.n56 10.6151
R749 B.n497 B.n496 10.6151
R750 B.n496 B.n495 10.6151
R751 B.n495 B.n58 10.6151
R752 B.n491 B.n58 10.6151
R753 B.n491 B.n490 10.6151
R754 B.n490 B.n489 10.6151
R755 B.n489 B.n60 10.6151
R756 B.n485 B.n60 10.6151
R757 B.n485 B.n484 10.6151
R758 B.n484 B.n483 10.6151
R759 B.n483 B.n62 10.6151
R760 B.n479 B.n62 10.6151
R761 B.n479 B.n478 10.6151
R762 B.n478 B.n477 10.6151
R763 B.n477 B.n64 10.6151
R764 B.n473 B.n64 10.6151
R765 B.n473 B.n472 10.6151
R766 B.n472 B.n471 10.6151
R767 B.n471 B.n66 10.6151
R768 B.n467 B.n66 10.6151
R769 B.n467 B.n466 10.6151
R770 B.n466 B.n465 10.6151
R771 B.n465 B.n68 10.6151
R772 B.n461 B.n68 10.6151
R773 B.n461 B.n460 10.6151
R774 B.n460 B.n459 10.6151
R775 B.n459 B.n70 10.6151
R776 B.n455 B.n70 10.6151
R777 B.n455 B.n454 10.6151
R778 B.n454 B.n453 10.6151
R779 B.n453 B.n72 10.6151
R780 B.n449 B.n72 10.6151
R781 B.n449 B.n448 10.6151
R782 B.n448 B.n447 10.6151
R783 B.n447 B.n74 10.6151
R784 B.n443 B.n74 10.6151
R785 B.n443 B.n442 10.6151
R786 B.n442 B.n441 10.6151
R787 B.n441 B.n76 10.6151
R788 B.n437 B.n76 10.6151
R789 B.n437 B.n436 10.6151
R790 B.n436 B.n435 10.6151
R791 B.n435 B.n78 10.6151
R792 B.n431 B.n78 10.6151
R793 B.n389 B.n388 10.6151
R794 B.n389 B.n92 10.6151
R795 B.n393 B.n92 10.6151
R796 B.n394 B.n393 10.6151
R797 B.n395 B.n394 10.6151
R798 B.n395 B.n90 10.6151
R799 B.n399 B.n90 10.6151
R800 B.n400 B.n399 10.6151
R801 B.n401 B.n400 10.6151
R802 B.n401 B.n88 10.6151
R803 B.n405 B.n88 10.6151
R804 B.n406 B.n405 10.6151
R805 B.n407 B.n406 10.6151
R806 B.n407 B.n86 10.6151
R807 B.n411 B.n86 10.6151
R808 B.n412 B.n411 10.6151
R809 B.n413 B.n412 10.6151
R810 B.n413 B.n84 10.6151
R811 B.n417 B.n84 10.6151
R812 B.n418 B.n417 10.6151
R813 B.n419 B.n418 10.6151
R814 B.n419 B.n82 10.6151
R815 B.n423 B.n82 10.6151
R816 B.n424 B.n423 10.6151
R817 B.n425 B.n424 10.6151
R818 B.n425 B.n80 10.6151
R819 B.n429 B.n80 10.6151
R820 B.n430 B.n429 10.6151
R821 B.n191 B.n190 10.6151
R822 B.n191 B.n162 10.6151
R823 B.n195 B.n162 10.6151
R824 B.n196 B.n195 10.6151
R825 B.n197 B.n196 10.6151
R826 B.n197 B.n160 10.6151
R827 B.n201 B.n160 10.6151
R828 B.n202 B.n201 10.6151
R829 B.n203 B.n202 10.6151
R830 B.n203 B.n158 10.6151
R831 B.n207 B.n158 10.6151
R832 B.n208 B.n207 10.6151
R833 B.n209 B.n208 10.6151
R834 B.n209 B.n156 10.6151
R835 B.n213 B.n156 10.6151
R836 B.n214 B.n213 10.6151
R837 B.n215 B.n214 10.6151
R838 B.n215 B.n154 10.6151
R839 B.n219 B.n154 10.6151
R840 B.n220 B.n219 10.6151
R841 B.n221 B.n220 10.6151
R842 B.n221 B.n152 10.6151
R843 B.n225 B.n152 10.6151
R844 B.n226 B.n225 10.6151
R845 B.n227 B.n226 10.6151
R846 B.n227 B.n150 10.6151
R847 B.n231 B.n150 10.6151
R848 B.n232 B.n231 10.6151
R849 B.n233 B.n232 10.6151
R850 B.n233 B.n148 10.6151
R851 B.n237 B.n148 10.6151
R852 B.n238 B.n237 10.6151
R853 B.n239 B.n238 10.6151
R854 B.n239 B.n146 10.6151
R855 B.n243 B.n146 10.6151
R856 B.n244 B.n243 10.6151
R857 B.n245 B.n244 10.6151
R858 B.n245 B.n144 10.6151
R859 B.n249 B.n144 10.6151
R860 B.n250 B.n249 10.6151
R861 B.n251 B.n250 10.6151
R862 B.n251 B.n142 10.6151
R863 B.n255 B.n142 10.6151
R864 B.n256 B.n255 10.6151
R865 B.n257 B.n256 10.6151
R866 B.n257 B.n140 10.6151
R867 B.n261 B.n140 10.6151
R868 B.n262 B.n261 10.6151
R869 B.n263 B.n262 10.6151
R870 B.n263 B.n138 10.6151
R871 B.n267 B.n138 10.6151
R872 B.n268 B.n267 10.6151
R873 B.n269 B.n268 10.6151
R874 B.n269 B.n136 10.6151
R875 B.n273 B.n136 10.6151
R876 B.n274 B.n273 10.6151
R877 B.n275 B.n274 10.6151
R878 B.n275 B.n134 10.6151
R879 B.n279 B.n134 10.6151
R880 B.n280 B.n279 10.6151
R881 B.n282 B.n130 10.6151
R882 B.n286 B.n130 10.6151
R883 B.n287 B.n286 10.6151
R884 B.n288 B.n287 10.6151
R885 B.n288 B.n128 10.6151
R886 B.n292 B.n128 10.6151
R887 B.n293 B.n292 10.6151
R888 B.n294 B.n293 10.6151
R889 B.n298 B.n297 10.6151
R890 B.n299 B.n298 10.6151
R891 B.n299 B.n122 10.6151
R892 B.n303 B.n122 10.6151
R893 B.n304 B.n303 10.6151
R894 B.n305 B.n304 10.6151
R895 B.n305 B.n120 10.6151
R896 B.n309 B.n120 10.6151
R897 B.n310 B.n309 10.6151
R898 B.n311 B.n310 10.6151
R899 B.n311 B.n118 10.6151
R900 B.n315 B.n118 10.6151
R901 B.n316 B.n315 10.6151
R902 B.n317 B.n316 10.6151
R903 B.n317 B.n116 10.6151
R904 B.n321 B.n116 10.6151
R905 B.n322 B.n321 10.6151
R906 B.n323 B.n322 10.6151
R907 B.n323 B.n114 10.6151
R908 B.n327 B.n114 10.6151
R909 B.n328 B.n327 10.6151
R910 B.n329 B.n328 10.6151
R911 B.n329 B.n112 10.6151
R912 B.n333 B.n112 10.6151
R913 B.n334 B.n333 10.6151
R914 B.n335 B.n334 10.6151
R915 B.n335 B.n110 10.6151
R916 B.n339 B.n110 10.6151
R917 B.n340 B.n339 10.6151
R918 B.n341 B.n340 10.6151
R919 B.n341 B.n108 10.6151
R920 B.n345 B.n108 10.6151
R921 B.n346 B.n345 10.6151
R922 B.n347 B.n346 10.6151
R923 B.n347 B.n106 10.6151
R924 B.n351 B.n106 10.6151
R925 B.n352 B.n351 10.6151
R926 B.n353 B.n352 10.6151
R927 B.n353 B.n104 10.6151
R928 B.n357 B.n104 10.6151
R929 B.n358 B.n357 10.6151
R930 B.n359 B.n358 10.6151
R931 B.n359 B.n102 10.6151
R932 B.n363 B.n102 10.6151
R933 B.n364 B.n363 10.6151
R934 B.n365 B.n364 10.6151
R935 B.n365 B.n100 10.6151
R936 B.n369 B.n100 10.6151
R937 B.n370 B.n369 10.6151
R938 B.n371 B.n370 10.6151
R939 B.n371 B.n98 10.6151
R940 B.n375 B.n98 10.6151
R941 B.n376 B.n375 10.6151
R942 B.n377 B.n376 10.6151
R943 B.n377 B.n96 10.6151
R944 B.n381 B.n96 10.6151
R945 B.n382 B.n381 10.6151
R946 B.n383 B.n382 10.6151
R947 B.n383 B.n94 10.6151
R948 B.n387 B.n94 10.6151
R949 B.n189 B.n164 10.6151
R950 B.n185 B.n164 10.6151
R951 B.n185 B.n184 10.6151
R952 B.n184 B.n183 10.6151
R953 B.n183 B.n166 10.6151
R954 B.n179 B.n166 10.6151
R955 B.n179 B.n178 10.6151
R956 B.n178 B.n177 10.6151
R957 B.n177 B.n168 10.6151
R958 B.n173 B.n168 10.6151
R959 B.n173 B.n172 10.6151
R960 B.n172 B.n171 10.6151
R961 B.n171 B.n0 10.6151
R962 B.n647 B.n1 10.6151
R963 B.n647 B.n646 10.6151
R964 B.n646 B.n645 10.6151
R965 B.n645 B.n4 10.6151
R966 B.n641 B.n4 10.6151
R967 B.n641 B.n640 10.6151
R968 B.n640 B.n639 10.6151
R969 B.n639 B.n6 10.6151
R970 B.n635 B.n6 10.6151
R971 B.n635 B.n634 10.6151
R972 B.n634 B.n633 10.6151
R973 B.n633 B.n8 10.6151
R974 B.n629 B.n8 10.6151
R975 B.n537 B.n536 7.18099
R976 B.n524 B.n48 7.18099
R977 B.n282 B.n281 7.18099
R978 B.n294 B.n126 7.18099
R979 B.n538 B.n537 3.43465
R980 B.n521 B.n48 3.43465
R981 B.n281 B.n280 3.43465
R982 B.n297 B.n126 3.43465
R983 B.n651 B.n0 2.81026
R984 B.n651 B.n1 2.81026
R985 VP.n1 VP.t2 1537.15
R986 VP.n1 VP.t3 1537.15
R987 VP.n0 VP.t1 1537.15
R988 VP.n0 VP.t0 1537.15
R989 VP.n2 VP.n0 205.573
R990 VP.n2 VP.n1 161.3
R991 VP VP.n2 0.0516364
R992 VTAIL.n5 VTAIL.t4 51.2853
R993 VTAIL.n4 VTAIL.t3 51.2853
R994 VTAIL.n3 VTAIL.t0 51.2853
R995 VTAIL.n7 VTAIL.t1 51.2852
R996 VTAIL.n0 VTAIL.t2 51.2852
R997 VTAIL.n1 VTAIL.t7 51.2852
R998 VTAIL.n2 VTAIL.t6 51.2852
R999 VTAIL.n6 VTAIL.t5 51.2852
R1000 VTAIL.n7 VTAIL.n6 28.8755
R1001 VTAIL.n3 VTAIL.n2 28.8755
R1002 VTAIL.n4 VTAIL.n3 0.560845
R1003 VTAIL.n6 VTAIL.n5 0.560845
R1004 VTAIL.n2 VTAIL.n1 0.560845
R1005 VTAIL.n5 VTAIL.n4 0.470328
R1006 VTAIL.n1 VTAIL.n0 0.470328
R1007 VTAIL VTAIL.n0 0.338862
R1008 VTAIL VTAIL.n7 0.222483
R1009 VDD1 VDD1.n1 108.073
R1010 VDD1 VDD1.n0 66.2633
R1011 VDD1.n0 VDD1.t2 1.75943
R1012 VDD1.n0 VDD1.t3 1.75943
R1013 VDD1.n1 VDD1.t0 1.75943
R1014 VDD1.n1 VDD1.t1 1.75943
R1015 VN.n0 VN.t3 1537.15
R1016 VN.n0 VN.t0 1537.15
R1017 VN.n1 VN.t1 1537.15
R1018 VN.n1 VN.t2 1537.15
R1019 VN VN.n1 205.953
R1020 VN VN.n0 161.351
R1021 VDD2.n2 VDD2.n0 107.549
R1022 VDD2.n2 VDD2.n1 66.2051
R1023 VDD2.n1 VDD2.t2 1.75943
R1024 VDD2.n1 VDD2.t1 1.75943
R1025 VDD2.n0 VDD2.t3 1.75943
R1026 VDD2.n0 VDD2.t0 1.75943
R1027 VDD2 VDD2.n2 0.0586897
C0 B VDD2 1.04955f
C1 VN VDD2 3.16465f
C2 B VN 0.749758f
C3 VTAIL w_n1360_n4668# 5.98369f
C4 VP VTAIL 2.37289f
C5 VDD1 VTAIL 13.4762f
C6 VP w_n1360_n4668# 2.17042f
C7 VDD1 w_n1360_n4668# 1.14662f
C8 VTAIL VDD2 13.5152f
C9 B VTAIL 5.17782f
C10 VN VTAIL 2.35879f
C11 VP VDD1 3.26677f
C12 VDD2 w_n1360_n4668# 1.15382f
C13 B w_n1360_n4668# 8.26788f
C14 VN w_n1360_n4668# 2.00135f
C15 VP VDD2 0.250699f
C16 VDD1 VDD2 0.482688f
C17 VP B 1.01971f
C18 B VDD1 1.03327f
C19 VP VN 5.73968f
C20 VN VDD1 0.148413f
C21 VDD2 VSUBS 0.791467f
C22 VDD1 VSUBS 6.588283f
C23 VTAIL VSUBS 0.994173f
C24 VN VSUBS 7.78747f
C25 VP VSUBS 1.352215f
C26 B VSUBS 2.844211f
C27 w_n1360_n4668# VSUBS 77.6016f
C28 VDD2.t3 VSUBS 0.484968f
C29 VDD2.t0 VSUBS 0.484968f
C30 VDD2.n0 VSUBS 5.11007f
C31 VDD2.t2 VSUBS 0.484968f
C32 VDD2.t1 VSUBS 0.484968f
C33 VDD2.n1 VSUBS 4.02535f
C34 VDD2.n2 VSUBS 5.5576f
C35 VN.t0 VSUBS 1.2084f
C36 VN.t3 VSUBS 1.2084f
C37 VN.n0 VSUBS 0.907226f
C38 VN.t1 VSUBS 1.2084f
C39 VN.t2 VSUBS 1.2084f
C40 VN.n1 VSUBS 1.62117f
C41 VDD1.t2 VSUBS 0.484315f
C42 VDD1.t3 VSUBS 0.484315f
C43 VDD1.n0 VSUBS 4.02059f
C44 VDD1.t0 VSUBS 0.484315f
C45 VDD1.t1 VSUBS 0.484315f
C46 VDD1.n1 VSUBS 5.13739f
C47 VTAIL.t2 VSUBS 3.72114f
C48 VTAIL.n0 VSUBS 0.823719f
C49 VTAIL.t7 VSUBS 3.72114f
C50 VTAIL.n1 VSUBS 0.841524f
C51 VTAIL.t6 VSUBS 3.72114f
C52 VTAIL.n2 VSUBS 2.46619f
C53 VTAIL.t0 VSUBS 3.72117f
C54 VTAIL.n3 VSUBS 2.46616f
C55 VTAIL.t3 VSUBS 3.72117f
C56 VTAIL.n4 VSUBS 0.841495f
C57 VTAIL.t4 VSUBS 3.72117f
C58 VTAIL.n5 VSUBS 0.841495f
C59 VTAIL.t5 VSUBS 3.72114f
C60 VTAIL.n6 VSUBS 2.46619f
C61 VTAIL.t1 VSUBS 3.72114f
C62 VTAIL.n7 VSUBS 2.43905f
C63 VP.t1 VSUBS 1.24509f
C64 VP.t0 VSUBS 1.24509f
C65 VP.n0 VSUBS 1.65506f
C66 VP.t3 VSUBS 1.24509f
C67 VP.t2 VSUBS 1.24509f
C68 VP.n1 VSUBS 0.934747f
C69 VP.n2 VSUBS 5.99179f
C70 B.n0 VSUBS 0.005252f
C71 B.n1 VSUBS 0.005252f
C72 B.n2 VSUBS 0.008306f
C73 B.n3 VSUBS 0.008306f
C74 B.n4 VSUBS 0.008306f
C75 B.n5 VSUBS 0.008306f
C76 B.n6 VSUBS 0.008306f
C77 B.n7 VSUBS 0.008306f
C78 B.n8 VSUBS 0.008306f
C79 B.n9 VSUBS 0.019149f
C80 B.n10 VSUBS 0.008306f
C81 B.n11 VSUBS 0.008306f
C82 B.n12 VSUBS 0.008306f
C83 B.n13 VSUBS 0.008306f
C84 B.n14 VSUBS 0.008306f
C85 B.n15 VSUBS 0.008306f
C86 B.n16 VSUBS 0.008306f
C87 B.n17 VSUBS 0.008306f
C88 B.n18 VSUBS 0.008306f
C89 B.n19 VSUBS 0.008306f
C90 B.n20 VSUBS 0.008306f
C91 B.n21 VSUBS 0.008306f
C92 B.n22 VSUBS 0.008306f
C93 B.n23 VSUBS 0.008306f
C94 B.n24 VSUBS 0.008306f
C95 B.n25 VSUBS 0.008306f
C96 B.n26 VSUBS 0.008306f
C97 B.n27 VSUBS 0.008306f
C98 B.n28 VSUBS 0.008306f
C99 B.n29 VSUBS 0.008306f
C100 B.n30 VSUBS 0.008306f
C101 B.n31 VSUBS 0.008306f
C102 B.n32 VSUBS 0.008306f
C103 B.n33 VSUBS 0.008306f
C104 B.n34 VSUBS 0.008306f
C105 B.n35 VSUBS 0.008306f
C106 B.n36 VSUBS 0.008306f
C107 B.n37 VSUBS 0.008306f
C108 B.n38 VSUBS 0.008306f
C109 B.n39 VSUBS 0.008306f
C110 B.t2 VSUBS 0.741574f
C111 B.t1 VSUBS 0.748085f
C112 B.t0 VSUBS 0.27243f
C113 B.n40 VSUBS 0.14881f
C114 B.n41 VSUBS 0.074383f
C115 B.n42 VSUBS 0.008306f
C116 B.n43 VSUBS 0.008306f
C117 B.n44 VSUBS 0.008306f
C118 B.n45 VSUBS 0.008306f
C119 B.t11 VSUBS 0.741545f
C120 B.t10 VSUBS 0.748058f
C121 B.t9 VSUBS 0.27243f
C122 B.n46 VSUBS 0.148837f
C123 B.n47 VSUBS 0.074412f
C124 B.n48 VSUBS 0.019243f
C125 B.n49 VSUBS 0.008306f
C126 B.n50 VSUBS 0.008306f
C127 B.n51 VSUBS 0.008306f
C128 B.n52 VSUBS 0.008306f
C129 B.n53 VSUBS 0.008306f
C130 B.n54 VSUBS 0.008306f
C131 B.n55 VSUBS 0.008306f
C132 B.n56 VSUBS 0.008306f
C133 B.n57 VSUBS 0.008306f
C134 B.n58 VSUBS 0.008306f
C135 B.n59 VSUBS 0.008306f
C136 B.n60 VSUBS 0.008306f
C137 B.n61 VSUBS 0.008306f
C138 B.n62 VSUBS 0.008306f
C139 B.n63 VSUBS 0.008306f
C140 B.n64 VSUBS 0.008306f
C141 B.n65 VSUBS 0.008306f
C142 B.n66 VSUBS 0.008306f
C143 B.n67 VSUBS 0.008306f
C144 B.n68 VSUBS 0.008306f
C145 B.n69 VSUBS 0.008306f
C146 B.n70 VSUBS 0.008306f
C147 B.n71 VSUBS 0.008306f
C148 B.n72 VSUBS 0.008306f
C149 B.n73 VSUBS 0.008306f
C150 B.n74 VSUBS 0.008306f
C151 B.n75 VSUBS 0.008306f
C152 B.n76 VSUBS 0.008306f
C153 B.n77 VSUBS 0.008306f
C154 B.n78 VSUBS 0.008306f
C155 B.n79 VSUBS 0.01847f
C156 B.n80 VSUBS 0.008306f
C157 B.n81 VSUBS 0.008306f
C158 B.n82 VSUBS 0.008306f
C159 B.n83 VSUBS 0.008306f
C160 B.n84 VSUBS 0.008306f
C161 B.n85 VSUBS 0.008306f
C162 B.n86 VSUBS 0.008306f
C163 B.n87 VSUBS 0.008306f
C164 B.n88 VSUBS 0.008306f
C165 B.n89 VSUBS 0.008306f
C166 B.n90 VSUBS 0.008306f
C167 B.n91 VSUBS 0.008306f
C168 B.n92 VSUBS 0.008306f
C169 B.n93 VSUBS 0.01847f
C170 B.n94 VSUBS 0.008306f
C171 B.n95 VSUBS 0.008306f
C172 B.n96 VSUBS 0.008306f
C173 B.n97 VSUBS 0.008306f
C174 B.n98 VSUBS 0.008306f
C175 B.n99 VSUBS 0.008306f
C176 B.n100 VSUBS 0.008306f
C177 B.n101 VSUBS 0.008306f
C178 B.n102 VSUBS 0.008306f
C179 B.n103 VSUBS 0.008306f
C180 B.n104 VSUBS 0.008306f
C181 B.n105 VSUBS 0.008306f
C182 B.n106 VSUBS 0.008306f
C183 B.n107 VSUBS 0.008306f
C184 B.n108 VSUBS 0.008306f
C185 B.n109 VSUBS 0.008306f
C186 B.n110 VSUBS 0.008306f
C187 B.n111 VSUBS 0.008306f
C188 B.n112 VSUBS 0.008306f
C189 B.n113 VSUBS 0.008306f
C190 B.n114 VSUBS 0.008306f
C191 B.n115 VSUBS 0.008306f
C192 B.n116 VSUBS 0.008306f
C193 B.n117 VSUBS 0.008306f
C194 B.n118 VSUBS 0.008306f
C195 B.n119 VSUBS 0.008306f
C196 B.n120 VSUBS 0.008306f
C197 B.n121 VSUBS 0.008306f
C198 B.n122 VSUBS 0.008306f
C199 B.n123 VSUBS 0.008306f
C200 B.t7 VSUBS 0.741545f
C201 B.t8 VSUBS 0.748058f
C202 B.t6 VSUBS 0.27243f
C203 B.n124 VSUBS 0.148837f
C204 B.n125 VSUBS 0.074412f
C205 B.n126 VSUBS 0.019243f
C206 B.n127 VSUBS 0.008306f
C207 B.n128 VSUBS 0.008306f
C208 B.n129 VSUBS 0.008306f
C209 B.n130 VSUBS 0.008306f
C210 B.n131 VSUBS 0.008306f
C211 B.t4 VSUBS 0.741574f
C212 B.t5 VSUBS 0.748085f
C213 B.t3 VSUBS 0.27243f
C214 B.n132 VSUBS 0.14881f
C215 B.n133 VSUBS 0.074383f
C216 B.n134 VSUBS 0.008306f
C217 B.n135 VSUBS 0.008306f
C218 B.n136 VSUBS 0.008306f
C219 B.n137 VSUBS 0.008306f
C220 B.n138 VSUBS 0.008306f
C221 B.n139 VSUBS 0.008306f
C222 B.n140 VSUBS 0.008306f
C223 B.n141 VSUBS 0.008306f
C224 B.n142 VSUBS 0.008306f
C225 B.n143 VSUBS 0.008306f
C226 B.n144 VSUBS 0.008306f
C227 B.n145 VSUBS 0.008306f
C228 B.n146 VSUBS 0.008306f
C229 B.n147 VSUBS 0.008306f
C230 B.n148 VSUBS 0.008306f
C231 B.n149 VSUBS 0.008306f
C232 B.n150 VSUBS 0.008306f
C233 B.n151 VSUBS 0.008306f
C234 B.n152 VSUBS 0.008306f
C235 B.n153 VSUBS 0.008306f
C236 B.n154 VSUBS 0.008306f
C237 B.n155 VSUBS 0.008306f
C238 B.n156 VSUBS 0.008306f
C239 B.n157 VSUBS 0.008306f
C240 B.n158 VSUBS 0.008306f
C241 B.n159 VSUBS 0.008306f
C242 B.n160 VSUBS 0.008306f
C243 B.n161 VSUBS 0.008306f
C244 B.n162 VSUBS 0.008306f
C245 B.n163 VSUBS 0.019149f
C246 B.n164 VSUBS 0.008306f
C247 B.n165 VSUBS 0.008306f
C248 B.n166 VSUBS 0.008306f
C249 B.n167 VSUBS 0.008306f
C250 B.n168 VSUBS 0.008306f
C251 B.n169 VSUBS 0.008306f
C252 B.n170 VSUBS 0.008306f
C253 B.n171 VSUBS 0.008306f
C254 B.n172 VSUBS 0.008306f
C255 B.n173 VSUBS 0.008306f
C256 B.n174 VSUBS 0.008306f
C257 B.n175 VSUBS 0.008306f
C258 B.n176 VSUBS 0.008306f
C259 B.n177 VSUBS 0.008306f
C260 B.n178 VSUBS 0.008306f
C261 B.n179 VSUBS 0.008306f
C262 B.n180 VSUBS 0.008306f
C263 B.n181 VSUBS 0.008306f
C264 B.n182 VSUBS 0.008306f
C265 B.n183 VSUBS 0.008306f
C266 B.n184 VSUBS 0.008306f
C267 B.n185 VSUBS 0.008306f
C268 B.n186 VSUBS 0.008306f
C269 B.n187 VSUBS 0.008306f
C270 B.n188 VSUBS 0.01847f
C271 B.n189 VSUBS 0.01847f
C272 B.n190 VSUBS 0.019149f
C273 B.n191 VSUBS 0.008306f
C274 B.n192 VSUBS 0.008306f
C275 B.n193 VSUBS 0.008306f
C276 B.n194 VSUBS 0.008306f
C277 B.n195 VSUBS 0.008306f
C278 B.n196 VSUBS 0.008306f
C279 B.n197 VSUBS 0.008306f
C280 B.n198 VSUBS 0.008306f
C281 B.n199 VSUBS 0.008306f
C282 B.n200 VSUBS 0.008306f
C283 B.n201 VSUBS 0.008306f
C284 B.n202 VSUBS 0.008306f
C285 B.n203 VSUBS 0.008306f
C286 B.n204 VSUBS 0.008306f
C287 B.n205 VSUBS 0.008306f
C288 B.n206 VSUBS 0.008306f
C289 B.n207 VSUBS 0.008306f
C290 B.n208 VSUBS 0.008306f
C291 B.n209 VSUBS 0.008306f
C292 B.n210 VSUBS 0.008306f
C293 B.n211 VSUBS 0.008306f
C294 B.n212 VSUBS 0.008306f
C295 B.n213 VSUBS 0.008306f
C296 B.n214 VSUBS 0.008306f
C297 B.n215 VSUBS 0.008306f
C298 B.n216 VSUBS 0.008306f
C299 B.n217 VSUBS 0.008306f
C300 B.n218 VSUBS 0.008306f
C301 B.n219 VSUBS 0.008306f
C302 B.n220 VSUBS 0.008306f
C303 B.n221 VSUBS 0.008306f
C304 B.n222 VSUBS 0.008306f
C305 B.n223 VSUBS 0.008306f
C306 B.n224 VSUBS 0.008306f
C307 B.n225 VSUBS 0.008306f
C308 B.n226 VSUBS 0.008306f
C309 B.n227 VSUBS 0.008306f
C310 B.n228 VSUBS 0.008306f
C311 B.n229 VSUBS 0.008306f
C312 B.n230 VSUBS 0.008306f
C313 B.n231 VSUBS 0.008306f
C314 B.n232 VSUBS 0.008306f
C315 B.n233 VSUBS 0.008306f
C316 B.n234 VSUBS 0.008306f
C317 B.n235 VSUBS 0.008306f
C318 B.n236 VSUBS 0.008306f
C319 B.n237 VSUBS 0.008306f
C320 B.n238 VSUBS 0.008306f
C321 B.n239 VSUBS 0.008306f
C322 B.n240 VSUBS 0.008306f
C323 B.n241 VSUBS 0.008306f
C324 B.n242 VSUBS 0.008306f
C325 B.n243 VSUBS 0.008306f
C326 B.n244 VSUBS 0.008306f
C327 B.n245 VSUBS 0.008306f
C328 B.n246 VSUBS 0.008306f
C329 B.n247 VSUBS 0.008306f
C330 B.n248 VSUBS 0.008306f
C331 B.n249 VSUBS 0.008306f
C332 B.n250 VSUBS 0.008306f
C333 B.n251 VSUBS 0.008306f
C334 B.n252 VSUBS 0.008306f
C335 B.n253 VSUBS 0.008306f
C336 B.n254 VSUBS 0.008306f
C337 B.n255 VSUBS 0.008306f
C338 B.n256 VSUBS 0.008306f
C339 B.n257 VSUBS 0.008306f
C340 B.n258 VSUBS 0.008306f
C341 B.n259 VSUBS 0.008306f
C342 B.n260 VSUBS 0.008306f
C343 B.n261 VSUBS 0.008306f
C344 B.n262 VSUBS 0.008306f
C345 B.n263 VSUBS 0.008306f
C346 B.n264 VSUBS 0.008306f
C347 B.n265 VSUBS 0.008306f
C348 B.n266 VSUBS 0.008306f
C349 B.n267 VSUBS 0.008306f
C350 B.n268 VSUBS 0.008306f
C351 B.n269 VSUBS 0.008306f
C352 B.n270 VSUBS 0.008306f
C353 B.n271 VSUBS 0.008306f
C354 B.n272 VSUBS 0.008306f
C355 B.n273 VSUBS 0.008306f
C356 B.n274 VSUBS 0.008306f
C357 B.n275 VSUBS 0.008306f
C358 B.n276 VSUBS 0.008306f
C359 B.n277 VSUBS 0.008306f
C360 B.n278 VSUBS 0.008306f
C361 B.n279 VSUBS 0.008306f
C362 B.n280 VSUBS 0.005496f
C363 B.n281 VSUBS 0.019243f
C364 B.n282 VSUBS 0.006962f
C365 B.n283 VSUBS 0.008306f
C366 B.n284 VSUBS 0.008306f
C367 B.n285 VSUBS 0.008306f
C368 B.n286 VSUBS 0.008306f
C369 B.n287 VSUBS 0.008306f
C370 B.n288 VSUBS 0.008306f
C371 B.n289 VSUBS 0.008306f
C372 B.n290 VSUBS 0.008306f
C373 B.n291 VSUBS 0.008306f
C374 B.n292 VSUBS 0.008306f
C375 B.n293 VSUBS 0.008306f
C376 B.n294 VSUBS 0.006962f
C377 B.n295 VSUBS 0.008306f
C378 B.n296 VSUBS 0.008306f
C379 B.n297 VSUBS 0.005496f
C380 B.n298 VSUBS 0.008306f
C381 B.n299 VSUBS 0.008306f
C382 B.n300 VSUBS 0.008306f
C383 B.n301 VSUBS 0.008306f
C384 B.n302 VSUBS 0.008306f
C385 B.n303 VSUBS 0.008306f
C386 B.n304 VSUBS 0.008306f
C387 B.n305 VSUBS 0.008306f
C388 B.n306 VSUBS 0.008306f
C389 B.n307 VSUBS 0.008306f
C390 B.n308 VSUBS 0.008306f
C391 B.n309 VSUBS 0.008306f
C392 B.n310 VSUBS 0.008306f
C393 B.n311 VSUBS 0.008306f
C394 B.n312 VSUBS 0.008306f
C395 B.n313 VSUBS 0.008306f
C396 B.n314 VSUBS 0.008306f
C397 B.n315 VSUBS 0.008306f
C398 B.n316 VSUBS 0.008306f
C399 B.n317 VSUBS 0.008306f
C400 B.n318 VSUBS 0.008306f
C401 B.n319 VSUBS 0.008306f
C402 B.n320 VSUBS 0.008306f
C403 B.n321 VSUBS 0.008306f
C404 B.n322 VSUBS 0.008306f
C405 B.n323 VSUBS 0.008306f
C406 B.n324 VSUBS 0.008306f
C407 B.n325 VSUBS 0.008306f
C408 B.n326 VSUBS 0.008306f
C409 B.n327 VSUBS 0.008306f
C410 B.n328 VSUBS 0.008306f
C411 B.n329 VSUBS 0.008306f
C412 B.n330 VSUBS 0.008306f
C413 B.n331 VSUBS 0.008306f
C414 B.n332 VSUBS 0.008306f
C415 B.n333 VSUBS 0.008306f
C416 B.n334 VSUBS 0.008306f
C417 B.n335 VSUBS 0.008306f
C418 B.n336 VSUBS 0.008306f
C419 B.n337 VSUBS 0.008306f
C420 B.n338 VSUBS 0.008306f
C421 B.n339 VSUBS 0.008306f
C422 B.n340 VSUBS 0.008306f
C423 B.n341 VSUBS 0.008306f
C424 B.n342 VSUBS 0.008306f
C425 B.n343 VSUBS 0.008306f
C426 B.n344 VSUBS 0.008306f
C427 B.n345 VSUBS 0.008306f
C428 B.n346 VSUBS 0.008306f
C429 B.n347 VSUBS 0.008306f
C430 B.n348 VSUBS 0.008306f
C431 B.n349 VSUBS 0.008306f
C432 B.n350 VSUBS 0.008306f
C433 B.n351 VSUBS 0.008306f
C434 B.n352 VSUBS 0.008306f
C435 B.n353 VSUBS 0.008306f
C436 B.n354 VSUBS 0.008306f
C437 B.n355 VSUBS 0.008306f
C438 B.n356 VSUBS 0.008306f
C439 B.n357 VSUBS 0.008306f
C440 B.n358 VSUBS 0.008306f
C441 B.n359 VSUBS 0.008306f
C442 B.n360 VSUBS 0.008306f
C443 B.n361 VSUBS 0.008306f
C444 B.n362 VSUBS 0.008306f
C445 B.n363 VSUBS 0.008306f
C446 B.n364 VSUBS 0.008306f
C447 B.n365 VSUBS 0.008306f
C448 B.n366 VSUBS 0.008306f
C449 B.n367 VSUBS 0.008306f
C450 B.n368 VSUBS 0.008306f
C451 B.n369 VSUBS 0.008306f
C452 B.n370 VSUBS 0.008306f
C453 B.n371 VSUBS 0.008306f
C454 B.n372 VSUBS 0.008306f
C455 B.n373 VSUBS 0.008306f
C456 B.n374 VSUBS 0.008306f
C457 B.n375 VSUBS 0.008306f
C458 B.n376 VSUBS 0.008306f
C459 B.n377 VSUBS 0.008306f
C460 B.n378 VSUBS 0.008306f
C461 B.n379 VSUBS 0.008306f
C462 B.n380 VSUBS 0.008306f
C463 B.n381 VSUBS 0.008306f
C464 B.n382 VSUBS 0.008306f
C465 B.n383 VSUBS 0.008306f
C466 B.n384 VSUBS 0.008306f
C467 B.n385 VSUBS 0.008306f
C468 B.n386 VSUBS 0.019149f
C469 B.n387 VSUBS 0.019149f
C470 B.n388 VSUBS 0.01847f
C471 B.n389 VSUBS 0.008306f
C472 B.n390 VSUBS 0.008306f
C473 B.n391 VSUBS 0.008306f
C474 B.n392 VSUBS 0.008306f
C475 B.n393 VSUBS 0.008306f
C476 B.n394 VSUBS 0.008306f
C477 B.n395 VSUBS 0.008306f
C478 B.n396 VSUBS 0.008306f
C479 B.n397 VSUBS 0.008306f
C480 B.n398 VSUBS 0.008306f
C481 B.n399 VSUBS 0.008306f
C482 B.n400 VSUBS 0.008306f
C483 B.n401 VSUBS 0.008306f
C484 B.n402 VSUBS 0.008306f
C485 B.n403 VSUBS 0.008306f
C486 B.n404 VSUBS 0.008306f
C487 B.n405 VSUBS 0.008306f
C488 B.n406 VSUBS 0.008306f
C489 B.n407 VSUBS 0.008306f
C490 B.n408 VSUBS 0.008306f
C491 B.n409 VSUBS 0.008306f
C492 B.n410 VSUBS 0.008306f
C493 B.n411 VSUBS 0.008306f
C494 B.n412 VSUBS 0.008306f
C495 B.n413 VSUBS 0.008306f
C496 B.n414 VSUBS 0.008306f
C497 B.n415 VSUBS 0.008306f
C498 B.n416 VSUBS 0.008306f
C499 B.n417 VSUBS 0.008306f
C500 B.n418 VSUBS 0.008306f
C501 B.n419 VSUBS 0.008306f
C502 B.n420 VSUBS 0.008306f
C503 B.n421 VSUBS 0.008306f
C504 B.n422 VSUBS 0.008306f
C505 B.n423 VSUBS 0.008306f
C506 B.n424 VSUBS 0.008306f
C507 B.n425 VSUBS 0.008306f
C508 B.n426 VSUBS 0.008306f
C509 B.n427 VSUBS 0.008306f
C510 B.n428 VSUBS 0.008306f
C511 B.n429 VSUBS 0.008306f
C512 B.n430 VSUBS 0.019502f
C513 B.n431 VSUBS 0.018118f
C514 B.n432 VSUBS 0.019149f
C515 B.n433 VSUBS 0.008306f
C516 B.n434 VSUBS 0.008306f
C517 B.n435 VSUBS 0.008306f
C518 B.n436 VSUBS 0.008306f
C519 B.n437 VSUBS 0.008306f
C520 B.n438 VSUBS 0.008306f
C521 B.n439 VSUBS 0.008306f
C522 B.n440 VSUBS 0.008306f
C523 B.n441 VSUBS 0.008306f
C524 B.n442 VSUBS 0.008306f
C525 B.n443 VSUBS 0.008306f
C526 B.n444 VSUBS 0.008306f
C527 B.n445 VSUBS 0.008306f
C528 B.n446 VSUBS 0.008306f
C529 B.n447 VSUBS 0.008306f
C530 B.n448 VSUBS 0.008306f
C531 B.n449 VSUBS 0.008306f
C532 B.n450 VSUBS 0.008306f
C533 B.n451 VSUBS 0.008306f
C534 B.n452 VSUBS 0.008306f
C535 B.n453 VSUBS 0.008306f
C536 B.n454 VSUBS 0.008306f
C537 B.n455 VSUBS 0.008306f
C538 B.n456 VSUBS 0.008306f
C539 B.n457 VSUBS 0.008306f
C540 B.n458 VSUBS 0.008306f
C541 B.n459 VSUBS 0.008306f
C542 B.n460 VSUBS 0.008306f
C543 B.n461 VSUBS 0.008306f
C544 B.n462 VSUBS 0.008306f
C545 B.n463 VSUBS 0.008306f
C546 B.n464 VSUBS 0.008306f
C547 B.n465 VSUBS 0.008306f
C548 B.n466 VSUBS 0.008306f
C549 B.n467 VSUBS 0.008306f
C550 B.n468 VSUBS 0.008306f
C551 B.n469 VSUBS 0.008306f
C552 B.n470 VSUBS 0.008306f
C553 B.n471 VSUBS 0.008306f
C554 B.n472 VSUBS 0.008306f
C555 B.n473 VSUBS 0.008306f
C556 B.n474 VSUBS 0.008306f
C557 B.n475 VSUBS 0.008306f
C558 B.n476 VSUBS 0.008306f
C559 B.n477 VSUBS 0.008306f
C560 B.n478 VSUBS 0.008306f
C561 B.n479 VSUBS 0.008306f
C562 B.n480 VSUBS 0.008306f
C563 B.n481 VSUBS 0.008306f
C564 B.n482 VSUBS 0.008306f
C565 B.n483 VSUBS 0.008306f
C566 B.n484 VSUBS 0.008306f
C567 B.n485 VSUBS 0.008306f
C568 B.n486 VSUBS 0.008306f
C569 B.n487 VSUBS 0.008306f
C570 B.n488 VSUBS 0.008306f
C571 B.n489 VSUBS 0.008306f
C572 B.n490 VSUBS 0.008306f
C573 B.n491 VSUBS 0.008306f
C574 B.n492 VSUBS 0.008306f
C575 B.n493 VSUBS 0.008306f
C576 B.n494 VSUBS 0.008306f
C577 B.n495 VSUBS 0.008306f
C578 B.n496 VSUBS 0.008306f
C579 B.n497 VSUBS 0.008306f
C580 B.n498 VSUBS 0.008306f
C581 B.n499 VSUBS 0.008306f
C582 B.n500 VSUBS 0.008306f
C583 B.n501 VSUBS 0.008306f
C584 B.n502 VSUBS 0.008306f
C585 B.n503 VSUBS 0.008306f
C586 B.n504 VSUBS 0.008306f
C587 B.n505 VSUBS 0.008306f
C588 B.n506 VSUBS 0.008306f
C589 B.n507 VSUBS 0.008306f
C590 B.n508 VSUBS 0.008306f
C591 B.n509 VSUBS 0.008306f
C592 B.n510 VSUBS 0.008306f
C593 B.n511 VSUBS 0.008306f
C594 B.n512 VSUBS 0.008306f
C595 B.n513 VSUBS 0.008306f
C596 B.n514 VSUBS 0.008306f
C597 B.n515 VSUBS 0.008306f
C598 B.n516 VSUBS 0.008306f
C599 B.n517 VSUBS 0.008306f
C600 B.n518 VSUBS 0.008306f
C601 B.n519 VSUBS 0.008306f
C602 B.n520 VSUBS 0.008306f
C603 B.n521 VSUBS 0.005496f
C604 B.n522 VSUBS 0.008306f
C605 B.n523 VSUBS 0.008306f
C606 B.n524 VSUBS 0.006962f
C607 B.n525 VSUBS 0.008306f
C608 B.n526 VSUBS 0.008306f
C609 B.n527 VSUBS 0.008306f
C610 B.n528 VSUBS 0.008306f
C611 B.n529 VSUBS 0.008306f
C612 B.n530 VSUBS 0.008306f
C613 B.n531 VSUBS 0.008306f
C614 B.n532 VSUBS 0.008306f
C615 B.n533 VSUBS 0.008306f
C616 B.n534 VSUBS 0.008306f
C617 B.n535 VSUBS 0.008306f
C618 B.n536 VSUBS 0.006962f
C619 B.n537 VSUBS 0.019243f
C620 B.n538 VSUBS 0.005496f
C621 B.n539 VSUBS 0.008306f
C622 B.n540 VSUBS 0.008306f
C623 B.n541 VSUBS 0.008306f
C624 B.n542 VSUBS 0.008306f
C625 B.n543 VSUBS 0.008306f
C626 B.n544 VSUBS 0.008306f
C627 B.n545 VSUBS 0.008306f
C628 B.n546 VSUBS 0.008306f
C629 B.n547 VSUBS 0.008306f
C630 B.n548 VSUBS 0.008306f
C631 B.n549 VSUBS 0.008306f
C632 B.n550 VSUBS 0.008306f
C633 B.n551 VSUBS 0.008306f
C634 B.n552 VSUBS 0.008306f
C635 B.n553 VSUBS 0.008306f
C636 B.n554 VSUBS 0.008306f
C637 B.n555 VSUBS 0.008306f
C638 B.n556 VSUBS 0.008306f
C639 B.n557 VSUBS 0.008306f
C640 B.n558 VSUBS 0.008306f
C641 B.n559 VSUBS 0.008306f
C642 B.n560 VSUBS 0.008306f
C643 B.n561 VSUBS 0.008306f
C644 B.n562 VSUBS 0.008306f
C645 B.n563 VSUBS 0.008306f
C646 B.n564 VSUBS 0.008306f
C647 B.n565 VSUBS 0.008306f
C648 B.n566 VSUBS 0.008306f
C649 B.n567 VSUBS 0.008306f
C650 B.n568 VSUBS 0.008306f
C651 B.n569 VSUBS 0.008306f
C652 B.n570 VSUBS 0.008306f
C653 B.n571 VSUBS 0.008306f
C654 B.n572 VSUBS 0.008306f
C655 B.n573 VSUBS 0.008306f
C656 B.n574 VSUBS 0.008306f
C657 B.n575 VSUBS 0.008306f
C658 B.n576 VSUBS 0.008306f
C659 B.n577 VSUBS 0.008306f
C660 B.n578 VSUBS 0.008306f
C661 B.n579 VSUBS 0.008306f
C662 B.n580 VSUBS 0.008306f
C663 B.n581 VSUBS 0.008306f
C664 B.n582 VSUBS 0.008306f
C665 B.n583 VSUBS 0.008306f
C666 B.n584 VSUBS 0.008306f
C667 B.n585 VSUBS 0.008306f
C668 B.n586 VSUBS 0.008306f
C669 B.n587 VSUBS 0.008306f
C670 B.n588 VSUBS 0.008306f
C671 B.n589 VSUBS 0.008306f
C672 B.n590 VSUBS 0.008306f
C673 B.n591 VSUBS 0.008306f
C674 B.n592 VSUBS 0.008306f
C675 B.n593 VSUBS 0.008306f
C676 B.n594 VSUBS 0.008306f
C677 B.n595 VSUBS 0.008306f
C678 B.n596 VSUBS 0.008306f
C679 B.n597 VSUBS 0.008306f
C680 B.n598 VSUBS 0.008306f
C681 B.n599 VSUBS 0.008306f
C682 B.n600 VSUBS 0.008306f
C683 B.n601 VSUBS 0.008306f
C684 B.n602 VSUBS 0.008306f
C685 B.n603 VSUBS 0.008306f
C686 B.n604 VSUBS 0.008306f
C687 B.n605 VSUBS 0.008306f
C688 B.n606 VSUBS 0.008306f
C689 B.n607 VSUBS 0.008306f
C690 B.n608 VSUBS 0.008306f
C691 B.n609 VSUBS 0.008306f
C692 B.n610 VSUBS 0.008306f
C693 B.n611 VSUBS 0.008306f
C694 B.n612 VSUBS 0.008306f
C695 B.n613 VSUBS 0.008306f
C696 B.n614 VSUBS 0.008306f
C697 B.n615 VSUBS 0.008306f
C698 B.n616 VSUBS 0.008306f
C699 B.n617 VSUBS 0.008306f
C700 B.n618 VSUBS 0.008306f
C701 B.n619 VSUBS 0.008306f
C702 B.n620 VSUBS 0.008306f
C703 B.n621 VSUBS 0.008306f
C704 B.n622 VSUBS 0.008306f
C705 B.n623 VSUBS 0.008306f
C706 B.n624 VSUBS 0.008306f
C707 B.n625 VSUBS 0.008306f
C708 B.n626 VSUBS 0.008306f
C709 B.n627 VSUBS 0.008306f
C710 B.n628 VSUBS 0.019149f
C711 B.n629 VSUBS 0.01847f
C712 B.n630 VSUBS 0.01847f
C713 B.n631 VSUBS 0.008306f
C714 B.n632 VSUBS 0.008306f
C715 B.n633 VSUBS 0.008306f
C716 B.n634 VSUBS 0.008306f
C717 B.n635 VSUBS 0.008306f
C718 B.n636 VSUBS 0.008306f
C719 B.n637 VSUBS 0.008306f
C720 B.n638 VSUBS 0.008306f
C721 B.n639 VSUBS 0.008306f
C722 B.n640 VSUBS 0.008306f
C723 B.n641 VSUBS 0.008306f
C724 B.n642 VSUBS 0.008306f
C725 B.n643 VSUBS 0.008306f
C726 B.n644 VSUBS 0.008306f
C727 B.n645 VSUBS 0.008306f
C728 B.n646 VSUBS 0.008306f
C729 B.n647 VSUBS 0.008306f
C730 B.n648 VSUBS 0.008306f
C731 B.n649 VSUBS 0.008306f
C732 B.n650 VSUBS 0.008306f
C733 B.n651 VSUBS 0.018807f
.ends

