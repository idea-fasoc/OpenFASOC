* NGSPICE file created from diff_pair_sample_1067.ext - technology: sky130A

.subckt diff_pair_sample_1067 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=4.6605 ps=24.68 w=11.95 l=2.46
X1 VTAIL.t8 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=1.97175 ps=12.28 w=11.95 l=2.46
X2 VDD1.t3 VP.t2 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=4.6605 ps=24.68 w=11.95 l=2.46
X3 VTAIL.t10 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=1.97175 ps=12.28 w=11.95 l=2.46
X4 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=0 ps=0 w=11.95 l=2.46
X5 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=1.97175 ps=12.28 w=11.95 l=2.46
X6 VTAIL.t5 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=1.97175 ps=12.28 w=11.95 l=2.46
X7 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=0 ps=0 w=11.95 l=2.46
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=0 ps=0 w=11.95 l=2.46
X9 VTAIL.t2 VN.t2 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=1.97175 ps=12.28 w=11.95 l=2.46
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=4.6605 ps=24.68 w=11.95 l=2.46
X11 VDD1.t1 VP.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=1.97175 ps=12.28 w=11.95 l=2.46
X12 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.97175 pd=12.28 as=4.6605 ps=24.68 w=11.95 l=2.46
X13 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=1.97175 ps=12.28 w=11.95 l=2.46
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=0 ps=0 w=11.95 l=2.46
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6605 pd=24.68 as=1.97175 ps=12.28 w=11.95 l=2.46
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n37 VP.n0 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n34 VP.n1 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n31 VP.n2 161.3
R10 VP.n30 VP.n29 161.3
R11 VP.n28 VP.n3 161.3
R12 VP.n27 VP.n26 161.3
R13 VP.n25 VP.n4 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n5 161.3
R16 VP.n9 VP.t4 152.004
R17 VP.n30 VP.t3 117.072
R18 VP.n20 VP.t5 117.072
R19 VP.n38 VP.t2 117.072
R20 VP.n10 VP.t1 117.072
R21 VP.n18 VP.t0 117.072
R22 VP.n21 VP.n20 96.5656
R23 VP.n39 VP.n38 96.5656
R24 VP.n19 VP.n18 96.5656
R25 VP.n26 VP.n25 50.6917
R26 VP.n32 VP.n1 50.6917
R27 VP.n12 VP.n7 50.6917
R28 VP.n21 VP.n19 48.1397
R29 VP.n10 VP.n9 48.0623
R30 VP.n25 VP.n24 30.2951
R31 VP.n36 VP.n1 30.2951
R32 VP.n16 VP.n7 30.2951
R33 VP.n24 VP.n5 24.4675
R34 VP.n26 VP.n3 24.4675
R35 VP.n30 VP.n3 24.4675
R36 VP.n31 VP.n30 24.4675
R37 VP.n32 VP.n31 24.4675
R38 VP.n37 VP.n36 24.4675
R39 VP.n17 VP.n16 24.4675
R40 VP.n11 VP.n10 24.4675
R41 VP.n12 VP.n11 24.4675
R42 VP.n20 VP.n5 14.1914
R43 VP.n38 VP.n37 14.1914
R44 VP.n18 VP.n17 14.1914
R45 VP.n9 VP.n8 6.56002
R46 VP.n19 VP.n6 0.278367
R47 VP.n22 VP.n21 0.278367
R48 VP.n39 VP.n0 0.278367
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153454
R64 VTAIL.n270 VTAIL.n269 289.615
R65 VTAIL.n66 VTAIL.n65 289.615
R66 VTAIL.n204 VTAIL.n203 289.615
R67 VTAIL.n136 VTAIL.n135 289.615
R68 VTAIL.n229 VTAIL.n228 185
R69 VTAIL.n231 VTAIL.n230 185
R70 VTAIL.n224 VTAIL.n223 185
R71 VTAIL.n237 VTAIL.n236 185
R72 VTAIL.n239 VTAIL.n238 185
R73 VTAIL.n220 VTAIL.n219 185
R74 VTAIL.n245 VTAIL.n244 185
R75 VTAIL.n247 VTAIL.n246 185
R76 VTAIL.n216 VTAIL.n215 185
R77 VTAIL.n253 VTAIL.n252 185
R78 VTAIL.n255 VTAIL.n254 185
R79 VTAIL.n212 VTAIL.n211 185
R80 VTAIL.n261 VTAIL.n260 185
R81 VTAIL.n263 VTAIL.n262 185
R82 VTAIL.n208 VTAIL.n207 185
R83 VTAIL.n269 VTAIL.n268 185
R84 VTAIL.n25 VTAIL.n24 185
R85 VTAIL.n27 VTAIL.n26 185
R86 VTAIL.n20 VTAIL.n19 185
R87 VTAIL.n33 VTAIL.n32 185
R88 VTAIL.n35 VTAIL.n34 185
R89 VTAIL.n16 VTAIL.n15 185
R90 VTAIL.n41 VTAIL.n40 185
R91 VTAIL.n43 VTAIL.n42 185
R92 VTAIL.n12 VTAIL.n11 185
R93 VTAIL.n49 VTAIL.n48 185
R94 VTAIL.n51 VTAIL.n50 185
R95 VTAIL.n8 VTAIL.n7 185
R96 VTAIL.n57 VTAIL.n56 185
R97 VTAIL.n59 VTAIL.n58 185
R98 VTAIL.n4 VTAIL.n3 185
R99 VTAIL.n65 VTAIL.n64 185
R100 VTAIL.n203 VTAIL.n202 185
R101 VTAIL.n142 VTAIL.n141 185
R102 VTAIL.n197 VTAIL.n196 185
R103 VTAIL.n195 VTAIL.n194 185
R104 VTAIL.n146 VTAIL.n145 185
R105 VTAIL.n189 VTAIL.n188 185
R106 VTAIL.n187 VTAIL.n186 185
R107 VTAIL.n150 VTAIL.n149 185
R108 VTAIL.n181 VTAIL.n180 185
R109 VTAIL.n179 VTAIL.n178 185
R110 VTAIL.n154 VTAIL.n153 185
R111 VTAIL.n173 VTAIL.n172 185
R112 VTAIL.n171 VTAIL.n170 185
R113 VTAIL.n158 VTAIL.n157 185
R114 VTAIL.n165 VTAIL.n164 185
R115 VTAIL.n163 VTAIL.n162 185
R116 VTAIL.n135 VTAIL.n134 185
R117 VTAIL.n74 VTAIL.n73 185
R118 VTAIL.n129 VTAIL.n128 185
R119 VTAIL.n127 VTAIL.n126 185
R120 VTAIL.n78 VTAIL.n77 185
R121 VTAIL.n121 VTAIL.n120 185
R122 VTAIL.n119 VTAIL.n118 185
R123 VTAIL.n82 VTAIL.n81 185
R124 VTAIL.n113 VTAIL.n112 185
R125 VTAIL.n111 VTAIL.n110 185
R126 VTAIL.n86 VTAIL.n85 185
R127 VTAIL.n105 VTAIL.n104 185
R128 VTAIL.n103 VTAIL.n102 185
R129 VTAIL.n90 VTAIL.n89 185
R130 VTAIL.n97 VTAIL.n96 185
R131 VTAIL.n95 VTAIL.n94 185
R132 VTAIL.n93 VTAIL.t4 147.659
R133 VTAIL.n227 VTAIL.t0 147.659
R134 VTAIL.n23 VTAIL.t11 147.659
R135 VTAIL.n161 VTAIL.t9 147.659
R136 VTAIL.n230 VTAIL.n229 104.615
R137 VTAIL.n230 VTAIL.n223 104.615
R138 VTAIL.n237 VTAIL.n223 104.615
R139 VTAIL.n238 VTAIL.n237 104.615
R140 VTAIL.n238 VTAIL.n219 104.615
R141 VTAIL.n245 VTAIL.n219 104.615
R142 VTAIL.n246 VTAIL.n245 104.615
R143 VTAIL.n246 VTAIL.n215 104.615
R144 VTAIL.n253 VTAIL.n215 104.615
R145 VTAIL.n254 VTAIL.n253 104.615
R146 VTAIL.n254 VTAIL.n211 104.615
R147 VTAIL.n261 VTAIL.n211 104.615
R148 VTAIL.n262 VTAIL.n261 104.615
R149 VTAIL.n262 VTAIL.n207 104.615
R150 VTAIL.n269 VTAIL.n207 104.615
R151 VTAIL.n26 VTAIL.n25 104.615
R152 VTAIL.n26 VTAIL.n19 104.615
R153 VTAIL.n33 VTAIL.n19 104.615
R154 VTAIL.n34 VTAIL.n33 104.615
R155 VTAIL.n34 VTAIL.n15 104.615
R156 VTAIL.n41 VTAIL.n15 104.615
R157 VTAIL.n42 VTAIL.n41 104.615
R158 VTAIL.n42 VTAIL.n11 104.615
R159 VTAIL.n49 VTAIL.n11 104.615
R160 VTAIL.n50 VTAIL.n49 104.615
R161 VTAIL.n50 VTAIL.n7 104.615
R162 VTAIL.n57 VTAIL.n7 104.615
R163 VTAIL.n58 VTAIL.n57 104.615
R164 VTAIL.n58 VTAIL.n3 104.615
R165 VTAIL.n65 VTAIL.n3 104.615
R166 VTAIL.n203 VTAIL.n141 104.615
R167 VTAIL.n196 VTAIL.n141 104.615
R168 VTAIL.n196 VTAIL.n195 104.615
R169 VTAIL.n195 VTAIL.n145 104.615
R170 VTAIL.n188 VTAIL.n145 104.615
R171 VTAIL.n188 VTAIL.n187 104.615
R172 VTAIL.n187 VTAIL.n149 104.615
R173 VTAIL.n180 VTAIL.n149 104.615
R174 VTAIL.n180 VTAIL.n179 104.615
R175 VTAIL.n179 VTAIL.n153 104.615
R176 VTAIL.n172 VTAIL.n153 104.615
R177 VTAIL.n172 VTAIL.n171 104.615
R178 VTAIL.n171 VTAIL.n157 104.615
R179 VTAIL.n164 VTAIL.n157 104.615
R180 VTAIL.n164 VTAIL.n163 104.615
R181 VTAIL.n135 VTAIL.n73 104.615
R182 VTAIL.n128 VTAIL.n73 104.615
R183 VTAIL.n128 VTAIL.n127 104.615
R184 VTAIL.n127 VTAIL.n77 104.615
R185 VTAIL.n120 VTAIL.n77 104.615
R186 VTAIL.n120 VTAIL.n119 104.615
R187 VTAIL.n119 VTAIL.n81 104.615
R188 VTAIL.n112 VTAIL.n81 104.615
R189 VTAIL.n112 VTAIL.n111 104.615
R190 VTAIL.n111 VTAIL.n85 104.615
R191 VTAIL.n104 VTAIL.n85 104.615
R192 VTAIL.n104 VTAIL.n103 104.615
R193 VTAIL.n103 VTAIL.n89 104.615
R194 VTAIL.n96 VTAIL.n89 104.615
R195 VTAIL.n96 VTAIL.n95 104.615
R196 VTAIL.n229 VTAIL.t0 52.3082
R197 VTAIL.n25 VTAIL.t11 52.3082
R198 VTAIL.n163 VTAIL.t9 52.3082
R199 VTAIL.n95 VTAIL.t4 52.3082
R200 VTAIL.n139 VTAIL.n138 48.2906
R201 VTAIL.n71 VTAIL.n70 48.2906
R202 VTAIL.n1 VTAIL.n0 48.2905
R203 VTAIL.n69 VTAIL.n68 48.2905
R204 VTAIL.n271 VTAIL.n270 34.7066
R205 VTAIL.n67 VTAIL.n66 34.7066
R206 VTAIL.n205 VTAIL.n204 34.7066
R207 VTAIL.n137 VTAIL.n136 34.7066
R208 VTAIL.n71 VTAIL.n69 27.4789
R209 VTAIL.n271 VTAIL.n205 25.0738
R210 VTAIL.n228 VTAIL.n227 15.6677
R211 VTAIL.n24 VTAIL.n23 15.6677
R212 VTAIL.n162 VTAIL.n161 15.6677
R213 VTAIL.n94 VTAIL.n93 15.6677
R214 VTAIL.n231 VTAIL.n226 12.8005
R215 VTAIL.n27 VTAIL.n22 12.8005
R216 VTAIL.n165 VTAIL.n160 12.8005
R217 VTAIL.n97 VTAIL.n92 12.8005
R218 VTAIL.n232 VTAIL.n224 12.0247
R219 VTAIL.n268 VTAIL.n206 12.0247
R220 VTAIL.n28 VTAIL.n20 12.0247
R221 VTAIL.n64 VTAIL.n2 12.0247
R222 VTAIL.n202 VTAIL.n140 12.0247
R223 VTAIL.n166 VTAIL.n158 12.0247
R224 VTAIL.n134 VTAIL.n72 12.0247
R225 VTAIL.n98 VTAIL.n90 12.0247
R226 VTAIL.n236 VTAIL.n235 11.249
R227 VTAIL.n267 VTAIL.n208 11.249
R228 VTAIL.n32 VTAIL.n31 11.249
R229 VTAIL.n63 VTAIL.n4 11.249
R230 VTAIL.n201 VTAIL.n142 11.249
R231 VTAIL.n170 VTAIL.n169 11.249
R232 VTAIL.n133 VTAIL.n74 11.249
R233 VTAIL.n102 VTAIL.n101 11.249
R234 VTAIL.n239 VTAIL.n222 10.4732
R235 VTAIL.n264 VTAIL.n263 10.4732
R236 VTAIL.n35 VTAIL.n18 10.4732
R237 VTAIL.n60 VTAIL.n59 10.4732
R238 VTAIL.n198 VTAIL.n197 10.4732
R239 VTAIL.n173 VTAIL.n156 10.4732
R240 VTAIL.n130 VTAIL.n129 10.4732
R241 VTAIL.n105 VTAIL.n88 10.4732
R242 VTAIL.n240 VTAIL.n220 9.69747
R243 VTAIL.n260 VTAIL.n210 9.69747
R244 VTAIL.n36 VTAIL.n16 9.69747
R245 VTAIL.n56 VTAIL.n6 9.69747
R246 VTAIL.n194 VTAIL.n144 9.69747
R247 VTAIL.n174 VTAIL.n154 9.69747
R248 VTAIL.n126 VTAIL.n76 9.69747
R249 VTAIL.n106 VTAIL.n86 9.69747
R250 VTAIL.n266 VTAIL.n206 9.45567
R251 VTAIL.n62 VTAIL.n2 9.45567
R252 VTAIL.n200 VTAIL.n140 9.45567
R253 VTAIL.n132 VTAIL.n72 9.45567
R254 VTAIL.n251 VTAIL.n250 9.3005
R255 VTAIL.n214 VTAIL.n213 9.3005
R256 VTAIL.n257 VTAIL.n256 9.3005
R257 VTAIL.n259 VTAIL.n258 9.3005
R258 VTAIL.n210 VTAIL.n209 9.3005
R259 VTAIL.n265 VTAIL.n264 9.3005
R260 VTAIL.n267 VTAIL.n266 9.3005
R261 VTAIL.n218 VTAIL.n217 9.3005
R262 VTAIL.n243 VTAIL.n242 9.3005
R263 VTAIL.n241 VTAIL.n240 9.3005
R264 VTAIL.n222 VTAIL.n221 9.3005
R265 VTAIL.n235 VTAIL.n234 9.3005
R266 VTAIL.n233 VTAIL.n232 9.3005
R267 VTAIL.n226 VTAIL.n225 9.3005
R268 VTAIL.n249 VTAIL.n248 9.3005
R269 VTAIL.n47 VTAIL.n46 9.3005
R270 VTAIL.n10 VTAIL.n9 9.3005
R271 VTAIL.n53 VTAIL.n52 9.3005
R272 VTAIL.n55 VTAIL.n54 9.3005
R273 VTAIL.n6 VTAIL.n5 9.3005
R274 VTAIL.n61 VTAIL.n60 9.3005
R275 VTAIL.n63 VTAIL.n62 9.3005
R276 VTAIL.n14 VTAIL.n13 9.3005
R277 VTAIL.n39 VTAIL.n38 9.3005
R278 VTAIL.n37 VTAIL.n36 9.3005
R279 VTAIL.n18 VTAIL.n17 9.3005
R280 VTAIL.n31 VTAIL.n30 9.3005
R281 VTAIL.n29 VTAIL.n28 9.3005
R282 VTAIL.n22 VTAIL.n21 9.3005
R283 VTAIL.n45 VTAIL.n44 9.3005
R284 VTAIL.n201 VTAIL.n200 9.3005
R285 VTAIL.n199 VTAIL.n198 9.3005
R286 VTAIL.n144 VTAIL.n143 9.3005
R287 VTAIL.n193 VTAIL.n192 9.3005
R288 VTAIL.n191 VTAIL.n190 9.3005
R289 VTAIL.n148 VTAIL.n147 9.3005
R290 VTAIL.n185 VTAIL.n184 9.3005
R291 VTAIL.n183 VTAIL.n182 9.3005
R292 VTAIL.n152 VTAIL.n151 9.3005
R293 VTAIL.n177 VTAIL.n176 9.3005
R294 VTAIL.n175 VTAIL.n174 9.3005
R295 VTAIL.n156 VTAIL.n155 9.3005
R296 VTAIL.n169 VTAIL.n168 9.3005
R297 VTAIL.n167 VTAIL.n166 9.3005
R298 VTAIL.n160 VTAIL.n159 9.3005
R299 VTAIL.n80 VTAIL.n79 9.3005
R300 VTAIL.n123 VTAIL.n122 9.3005
R301 VTAIL.n125 VTAIL.n124 9.3005
R302 VTAIL.n76 VTAIL.n75 9.3005
R303 VTAIL.n131 VTAIL.n130 9.3005
R304 VTAIL.n133 VTAIL.n132 9.3005
R305 VTAIL.n117 VTAIL.n116 9.3005
R306 VTAIL.n115 VTAIL.n114 9.3005
R307 VTAIL.n84 VTAIL.n83 9.3005
R308 VTAIL.n109 VTAIL.n108 9.3005
R309 VTAIL.n107 VTAIL.n106 9.3005
R310 VTAIL.n88 VTAIL.n87 9.3005
R311 VTAIL.n101 VTAIL.n100 9.3005
R312 VTAIL.n99 VTAIL.n98 9.3005
R313 VTAIL.n92 VTAIL.n91 9.3005
R314 VTAIL.n244 VTAIL.n243 8.92171
R315 VTAIL.n259 VTAIL.n212 8.92171
R316 VTAIL.n40 VTAIL.n39 8.92171
R317 VTAIL.n55 VTAIL.n8 8.92171
R318 VTAIL.n193 VTAIL.n146 8.92171
R319 VTAIL.n178 VTAIL.n177 8.92171
R320 VTAIL.n125 VTAIL.n78 8.92171
R321 VTAIL.n110 VTAIL.n109 8.92171
R322 VTAIL.n247 VTAIL.n218 8.14595
R323 VTAIL.n256 VTAIL.n255 8.14595
R324 VTAIL.n43 VTAIL.n14 8.14595
R325 VTAIL.n52 VTAIL.n51 8.14595
R326 VTAIL.n190 VTAIL.n189 8.14595
R327 VTAIL.n181 VTAIL.n152 8.14595
R328 VTAIL.n122 VTAIL.n121 8.14595
R329 VTAIL.n113 VTAIL.n84 8.14595
R330 VTAIL.n248 VTAIL.n216 7.3702
R331 VTAIL.n252 VTAIL.n214 7.3702
R332 VTAIL.n44 VTAIL.n12 7.3702
R333 VTAIL.n48 VTAIL.n10 7.3702
R334 VTAIL.n186 VTAIL.n148 7.3702
R335 VTAIL.n182 VTAIL.n150 7.3702
R336 VTAIL.n118 VTAIL.n80 7.3702
R337 VTAIL.n114 VTAIL.n82 7.3702
R338 VTAIL.n251 VTAIL.n216 6.59444
R339 VTAIL.n252 VTAIL.n251 6.59444
R340 VTAIL.n47 VTAIL.n12 6.59444
R341 VTAIL.n48 VTAIL.n47 6.59444
R342 VTAIL.n186 VTAIL.n185 6.59444
R343 VTAIL.n185 VTAIL.n150 6.59444
R344 VTAIL.n118 VTAIL.n117 6.59444
R345 VTAIL.n117 VTAIL.n82 6.59444
R346 VTAIL.n248 VTAIL.n247 5.81868
R347 VTAIL.n255 VTAIL.n214 5.81868
R348 VTAIL.n44 VTAIL.n43 5.81868
R349 VTAIL.n51 VTAIL.n10 5.81868
R350 VTAIL.n189 VTAIL.n148 5.81868
R351 VTAIL.n182 VTAIL.n181 5.81868
R352 VTAIL.n121 VTAIL.n80 5.81868
R353 VTAIL.n114 VTAIL.n113 5.81868
R354 VTAIL.n244 VTAIL.n218 5.04292
R355 VTAIL.n256 VTAIL.n212 5.04292
R356 VTAIL.n40 VTAIL.n14 5.04292
R357 VTAIL.n52 VTAIL.n8 5.04292
R358 VTAIL.n190 VTAIL.n146 5.04292
R359 VTAIL.n178 VTAIL.n152 5.04292
R360 VTAIL.n122 VTAIL.n78 5.04292
R361 VTAIL.n110 VTAIL.n84 5.04292
R362 VTAIL.n93 VTAIL.n91 4.38563
R363 VTAIL.n227 VTAIL.n225 4.38563
R364 VTAIL.n23 VTAIL.n21 4.38563
R365 VTAIL.n161 VTAIL.n159 4.38563
R366 VTAIL.n243 VTAIL.n220 4.26717
R367 VTAIL.n260 VTAIL.n259 4.26717
R368 VTAIL.n39 VTAIL.n16 4.26717
R369 VTAIL.n56 VTAIL.n55 4.26717
R370 VTAIL.n194 VTAIL.n193 4.26717
R371 VTAIL.n177 VTAIL.n154 4.26717
R372 VTAIL.n126 VTAIL.n125 4.26717
R373 VTAIL.n109 VTAIL.n86 4.26717
R374 VTAIL.n240 VTAIL.n239 3.49141
R375 VTAIL.n263 VTAIL.n210 3.49141
R376 VTAIL.n36 VTAIL.n35 3.49141
R377 VTAIL.n59 VTAIL.n6 3.49141
R378 VTAIL.n197 VTAIL.n144 3.49141
R379 VTAIL.n174 VTAIL.n173 3.49141
R380 VTAIL.n129 VTAIL.n76 3.49141
R381 VTAIL.n106 VTAIL.n105 3.49141
R382 VTAIL.n236 VTAIL.n222 2.71565
R383 VTAIL.n264 VTAIL.n208 2.71565
R384 VTAIL.n32 VTAIL.n18 2.71565
R385 VTAIL.n60 VTAIL.n4 2.71565
R386 VTAIL.n198 VTAIL.n142 2.71565
R387 VTAIL.n170 VTAIL.n156 2.71565
R388 VTAIL.n130 VTAIL.n74 2.71565
R389 VTAIL.n102 VTAIL.n88 2.71565
R390 VTAIL.n137 VTAIL.n71 2.40567
R391 VTAIL.n205 VTAIL.n139 2.40567
R392 VTAIL.n69 VTAIL.n67 2.40567
R393 VTAIL.n235 VTAIL.n224 1.93989
R394 VTAIL.n268 VTAIL.n267 1.93989
R395 VTAIL.n31 VTAIL.n20 1.93989
R396 VTAIL.n64 VTAIL.n63 1.93989
R397 VTAIL.n202 VTAIL.n201 1.93989
R398 VTAIL.n169 VTAIL.n158 1.93989
R399 VTAIL.n134 VTAIL.n133 1.93989
R400 VTAIL.n101 VTAIL.n90 1.93989
R401 VTAIL VTAIL.n271 1.74619
R402 VTAIL.n139 VTAIL.n137 1.67291
R403 VTAIL.n67 VTAIL.n1 1.67291
R404 VTAIL.n0 VTAIL.t1 1.6574
R405 VTAIL.n0 VTAIL.t5 1.6574
R406 VTAIL.n68 VTAIL.t6 1.6574
R407 VTAIL.n68 VTAIL.t10 1.6574
R408 VTAIL.n138 VTAIL.t7 1.6574
R409 VTAIL.n138 VTAIL.t8 1.6574
R410 VTAIL.n70 VTAIL.t3 1.6574
R411 VTAIL.n70 VTAIL.t2 1.6574
R412 VTAIL.n232 VTAIL.n231 1.16414
R413 VTAIL.n270 VTAIL.n206 1.16414
R414 VTAIL.n28 VTAIL.n27 1.16414
R415 VTAIL.n66 VTAIL.n2 1.16414
R416 VTAIL.n204 VTAIL.n140 1.16414
R417 VTAIL.n166 VTAIL.n165 1.16414
R418 VTAIL.n136 VTAIL.n72 1.16414
R419 VTAIL.n98 VTAIL.n97 1.16414
R420 VTAIL VTAIL.n1 0.659983
R421 VTAIL.n228 VTAIL.n226 0.388379
R422 VTAIL.n24 VTAIL.n22 0.388379
R423 VTAIL.n162 VTAIL.n160 0.388379
R424 VTAIL.n94 VTAIL.n92 0.388379
R425 VTAIL.n233 VTAIL.n225 0.155672
R426 VTAIL.n234 VTAIL.n233 0.155672
R427 VTAIL.n234 VTAIL.n221 0.155672
R428 VTAIL.n241 VTAIL.n221 0.155672
R429 VTAIL.n242 VTAIL.n241 0.155672
R430 VTAIL.n242 VTAIL.n217 0.155672
R431 VTAIL.n249 VTAIL.n217 0.155672
R432 VTAIL.n250 VTAIL.n249 0.155672
R433 VTAIL.n250 VTAIL.n213 0.155672
R434 VTAIL.n257 VTAIL.n213 0.155672
R435 VTAIL.n258 VTAIL.n257 0.155672
R436 VTAIL.n258 VTAIL.n209 0.155672
R437 VTAIL.n265 VTAIL.n209 0.155672
R438 VTAIL.n266 VTAIL.n265 0.155672
R439 VTAIL.n29 VTAIL.n21 0.155672
R440 VTAIL.n30 VTAIL.n29 0.155672
R441 VTAIL.n30 VTAIL.n17 0.155672
R442 VTAIL.n37 VTAIL.n17 0.155672
R443 VTAIL.n38 VTAIL.n37 0.155672
R444 VTAIL.n38 VTAIL.n13 0.155672
R445 VTAIL.n45 VTAIL.n13 0.155672
R446 VTAIL.n46 VTAIL.n45 0.155672
R447 VTAIL.n46 VTAIL.n9 0.155672
R448 VTAIL.n53 VTAIL.n9 0.155672
R449 VTAIL.n54 VTAIL.n53 0.155672
R450 VTAIL.n54 VTAIL.n5 0.155672
R451 VTAIL.n61 VTAIL.n5 0.155672
R452 VTAIL.n62 VTAIL.n61 0.155672
R453 VTAIL.n200 VTAIL.n199 0.155672
R454 VTAIL.n199 VTAIL.n143 0.155672
R455 VTAIL.n192 VTAIL.n143 0.155672
R456 VTAIL.n192 VTAIL.n191 0.155672
R457 VTAIL.n191 VTAIL.n147 0.155672
R458 VTAIL.n184 VTAIL.n147 0.155672
R459 VTAIL.n184 VTAIL.n183 0.155672
R460 VTAIL.n183 VTAIL.n151 0.155672
R461 VTAIL.n176 VTAIL.n151 0.155672
R462 VTAIL.n176 VTAIL.n175 0.155672
R463 VTAIL.n175 VTAIL.n155 0.155672
R464 VTAIL.n168 VTAIL.n155 0.155672
R465 VTAIL.n168 VTAIL.n167 0.155672
R466 VTAIL.n167 VTAIL.n159 0.155672
R467 VTAIL.n132 VTAIL.n131 0.155672
R468 VTAIL.n131 VTAIL.n75 0.155672
R469 VTAIL.n124 VTAIL.n75 0.155672
R470 VTAIL.n124 VTAIL.n123 0.155672
R471 VTAIL.n123 VTAIL.n79 0.155672
R472 VTAIL.n116 VTAIL.n79 0.155672
R473 VTAIL.n116 VTAIL.n115 0.155672
R474 VTAIL.n115 VTAIL.n83 0.155672
R475 VTAIL.n108 VTAIL.n83 0.155672
R476 VTAIL.n108 VTAIL.n107 0.155672
R477 VTAIL.n107 VTAIL.n87 0.155672
R478 VTAIL.n100 VTAIL.n87 0.155672
R479 VTAIL.n100 VTAIL.n99 0.155672
R480 VTAIL.n99 VTAIL.n91 0.155672
R481 VDD1.n64 VDD1.n63 289.615
R482 VDD1.n129 VDD1.n128 289.615
R483 VDD1.n63 VDD1.n62 185
R484 VDD1.n2 VDD1.n1 185
R485 VDD1.n57 VDD1.n56 185
R486 VDD1.n55 VDD1.n54 185
R487 VDD1.n6 VDD1.n5 185
R488 VDD1.n49 VDD1.n48 185
R489 VDD1.n47 VDD1.n46 185
R490 VDD1.n10 VDD1.n9 185
R491 VDD1.n41 VDD1.n40 185
R492 VDD1.n39 VDD1.n38 185
R493 VDD1.n14 VDD1.n13 185
R494 VDD1.n33 VDD1.n32 185
R495 VDD1.n31 VDD1.n30 185
R496 VDD1.n18 VDD1.n17 185
R497 VDD1.n25 VDD1.n24 185
R498 VDD1.n23 VDD1.n22 185
R499 VDD1.n88 VDD1.n87 185
R500 VDD1.n90 VDD1.n89 185
R501 VDD1.n83 VDD1.n82 185
R502 VDD1.n96 VDD1.n95 185
R503 VDD1.n98 VDD1.n97 185
R504 VDD1.n79 VDD1.n78 185
R505 VDD1.n104 VDD1.n103 185
R506 VDD1.n106 VDD1.n105 185
R507 VDD1.n75 VDD1.n74 185
R508 VDD1.n112 VDD1.n111 185
R509 VDD1.n114 VDD1.n113 185
R510 VDD1.n71 VDD1.n70 185
R511 VDD1.n120 VDD1.n119 185
R512 VDD1.n122 VDD1.n121 185
R513 VDD1.n67 VDD1.n66 185
R514 VDD1.n128 VDD1.n127 185
R515 VDD1.n21 VDD1.t1 147.659
R516 VDD1.n86 VDD1.t0 147.659
R517 VDD1.n63 VDD1.n1 104.615
R518 VDD1.n56 VDD1.n1 104.615
R519 VDD1.n56 VDD1.n55 104.615
R520 VDD1.n55 VDD1.n5 104.615
R521 VDD1.n48 VDD1.n5 104.615
R522 VDD1.n48 VDD1.n47 104.615
R523 VDD1.n47 VDD1.n9 104.615
R524 VDD1.n40 VDD1.n9 104.615
R525 VDD1.n40 VDD1.n39 104.615
R526 VDD1.n39 VDD1.n13 104.615
R527 VDD1.n32 VDD1.n13 104.615
R528 VDD1.n32 VDD1.n31 104.615
R529 VDD1.n31 VDD1.n17 104.615
R530 VDD1.n24 VDD1.n17 104.615
R531 VDD1.n24 VDD1.n23 104.615
R532 VDD1.n89 VDD1.n88 104.615
R533 VDD1.n89 VDD1.n82 104.615
R534 VDD1.n96 VDD1.n82 104.615
R535 VDD1.n97 VDD1.n96 104.615
R536 VDD1.n97 VDD1.n78 104.615
R537 VDD1.n104 VDD1.n78 104.615
R538 VDD1.n105 VDD1.n104 104.615
R539 VDD1.n105 VDD1.n74 104.615
R540 VDD1.n112 VDD1.n74 104.615
R541 VDD1.n113 VDD1.n112 104.615
R542 VDD1.n113 VDD1.n70 104.615
R543 VDD1.n120 VDD1.n70 104.615
R544 VDD1.n121 VDD1.n120 104.615
R545 VDD1.n121 VDD1.n66 104.615
R546 VDD1.n128 VDD1.n66 104.615
R547 VDD1.n131 VDD1.n130 65.5152
R548 VDD1.n133 VDD1.n132 64.9684
R549 VDD1 VDD1.n64 53.2474
R550 VDD1.n131 VDD1.n129 53.1339
R551 VDD1.n23 VDD1.t1 52.3082
R552 VDD1.n88 VDD1.t0 52.3082
R553 VDD1.n133 VDD1.n131 43.6194
R554 VDD1.n22 VDD1.n21 15.6677
R555 VDD1.n87 VDD1.n86 15.6677
R556 VDD1.n25 VDD1.n20 12.8005
R557 VDD1.n90 VDD1.n85 12.8005
R558 VDD1.n62 VDD1.n0 12.0247
R559 VDD1.n26 VDD1.n18 12.0247
R560 VDD1.n91 VDD1.n83 12.0247
R561 VDD1.n127 VDD1.n65 12.0247
R562 VDD1.n61 VDD1.n2 11.249
R563 VDD1.n30 VDD1.n29 11.249
R564 VDD1.n95 VDD1.n94 11.249
R565 VDD1.n126 VDD1.n67 11.249
R566 VDD1.n58 VDD1.n57 10.4732
R567 VDD1.n33 VDD1.n16 10.4732
R568 VDD1.n98 VDD1.n81 10.4732
R569 VDD1.n123 VDD1.n122 10.4732
R570 VDD1.n54 VDD1.n4 9.69747
R571 VDD1.n34 VDD1.n14 9.69747
R572 VDD1.n99 VDD1.n79 9.69747
R573 VDD1.n119 VDD1.n69 9.69747
R574 VDD1.n60 VDD1.n0 9.45567
R575 VDD1.n125 VDD1.n65 9.45567
R576 VDD1.n8 VDD1.n7 9.3005
R577 VDD1.n51 VDD1.n50 9.3005
R578 VDD1.n53 VDD1.n52 9.3005
R579 VDD1.n4 VDD1.n3 9.3005
R580 VDD1.n59 VDD1.n58 9.3005
R581 VDD1.n61 VDD1.n60 9.3005
R582 VDD1.n45 VDD1.n44 9.3005
R583 VDD1.n43 VDD1.n42 9.3005
R584 VDD1.n12 VDD1.n11 9.3005
R585 VDD1.n37 VDD1.n36 9.3005
R586 VDD1.n35 VDD1.n34 9.3005
R587 VDD1.n16 VDD1.n15 9.3005
R588 VDD1.n29 VDD1.n28 9.3005
R589 VDD1.n27 VDD1.n26 9.3005
R590 VDD1.n20 VDD1.n19 9.3005
R591 VDD1.n110 VDD1.n109 9.3005
R592 VDD1.n73 VDD1.n72 9.3005
R593 VDD1.n116 VDD1.n115 9.3005
R594 VDD1.n118 VDD1.n117 9.3005
R595 VDD1.n69 VDD1.n68 9.3005
R596 VDD1.n124 VDD1.n123 9.3005
R597 VDD1.n126 VDD1.n125 9.3005
R598 VDD1.n77 VDD1.n76 9.3005
R599 VDD1.n102 VDD1.n101 9.3005
R600 VDD1.n100 VDD1.n99 9.3005
R601 VDD1.n81 VDD1.n80 9.3005
R602 VDD1.n94 VDD1.n93 9.3005
R603 VDD1.n92 VDD1.n91 9.3005
R604 VDD1.n85 VDD1.n84 9.3005
R605 VDD1.n108 VDD1.n107 9.3005
R606 VDD1.n53 VDD1.n6 8.92171
R607 VDD1.n38 VDD1.n37 8.92171
R608 VDD1.n103 VDD1.n102 8.92171
R609 VDD1.n118 VDD1.n71 8.92171
R610 VDD1.n50 VDD1.n49 8.14595
R611 VDD1.n41 VDD1.n12 8.14595
R612 VDD1.n106 VDD1.n77 8.14595
R613 VDD1.n115 VDD1.n114 8.14595
R614 VDD1.n46 VDD1.n8 7.3702
R615 VDD1.n42 VDD1.n10 7.3702
R616 VDD1.n107 VDD1.n75 7.3702
R617 VDD1.n111 VDD1.n73 7.3702
R618 VDD1.n46 VDD1.n45 6.59444
R619 VDD1.n45 VDD1.n10 6.59444
R620 VDD1.n110 VDD1.n75 6.59444
R621 VDD1.n111 VDD1.n110 6.59444
R622 VDD1.n49 VDD1.n8 5.81868
R623 VDD1.n42 VDD1.n41 5.81868
R624 VDD1.n107 VDD1.n106 5.81868
R625 VDD1.n114 VDD1.n73 5.81868
R626 VDD1.n50 VDD1.n6 5.04292
R627 VDD1.n38 VDD1.n12 5.04292
R628 VDD1.n103 VDD1.n77 5.04292
R629 VDD1.n115 VDD1.n71 5.04292
R630 VDD1.n21 VDD1.n19 4.38563
R631 VDD1.n86 VDD1.n84 4.38563
R632 VDD1.n54 VDD1.n53 4.26717
R633 VDD1.n37 VDD1.n14 4.26717
R634 VDD1.n102 VDD1.n79 4.26717
R635 VDD1.n119 VDD1.n118 4.26717
R636 VDD1.n57 VDD1.n4 3.49141
R637 VDD1.n34 VDD1.n33 3.49141
R638 VDD1.n99 VDD1.n98 3.49141
R639 VDD1.n122 VDD1.n69 3.49141
R640 VDD1.n58 VDD1.n2 2.71565
R641 VDD1.n30 VDD1.n16 2.71565
R642 VDD1.n95 VDD1.n81 2.71565
R643 VDD1.n123 VDD1.n67 2.71565
R644 VDD1.n62 VDD1.n61 1.93989
R645 VDD1.n29 VDD1.n18 1.93989
R646 VDD1.n94 VDD1.n83 1.93989
R647 VDD1.n127 VDD1.n126 1.93989
R648 VDD1.n132 VDD1.t4 1.6574
R649 VDD1.n132 VDD1.t5 1.6574
R650 VDD1.n130 VDD1.t2 1.6574
R651 VDD1.n130 VDD1.t3 1.6574
R652 VDD1.n64 VDD1.n0 1.16414
R653 VDD1.n26 VDD1.n25 1.16414
R654 VDD1.n91 VDD1.n90 1.16414
R655 VDD1.n129 VDD1.n65 1.16414
R656 VDD1 VDD1.n133 0.543603
R657 VDD1.n22 VDD1.n20 0.388379
R658 VDD1.n87 VDD1.n85 0.388379
R659 VDD1.n60 VDD1.n59 0.155672
R660 VDD1.n59 VDD1.n3 0.155672
R661 VDD1.n52 VDD1.n3 0.155672
R662 VDD1.n52 VDD1.n51 0.155672
R663 VDD1.n51 VDD1.n7 0.155672
R664 VDD1.n44 VDD1.n7 0.155672
R665 VDD1.n44 VDD1.n43 0.155672
R666 VDD1.n43 VDD1.n11 0.155672
R667 VDD1.n36 VDD1.n11 0.155672
R668 VDD1.n36 VDD1.n35 0.155672
R669 VDD1.n35 VDD1.n15 0.155672
R670 VDD1.n28 VDD1.n15 0.155672
R671 VDD1.n28 VDD1.n27 0.155672
R672 VDD1.n27 VDD1.n19 0.155672
R673 VDD1.n92 VDD1.n84 0.155672
R674 VDD1.n93 VDD1.n92 0.155672
R675 VDD1.n93 VDD1.n80 0.155672
R676 VDD1.n100 VDD1.n80 0.155672
R677 VDD1.n101 VDD1.n100 0.155672
R678 VDD1.n101 VDD1.n76 0.155672
R679 VDD1.n108 VDD1.n76 0.155672
R680 VDD1.n109 VDD1.n108 0.155672
R681 VDD1.n109 VDD1.n72 0.155672
R682 VDD1.n116 VDD1.n72 0.155672
R683 VDD1.n117 VDD1.n116 0.155672
R684 VDD1.n117 VDD1.n68 0.155672
R685 VDD1.n124 VDD1.n68 0.155672
R686 VDD1.n125 VDD1.n124 0.155672
R687 B.n807 B.n806 585
R688 B.n808 B.n807 585
R689 B.n312 B.n123 585
R690 B.n311 B.n310 585
R691 B.n309 B.n308 585
R692 B.n307 B.n306 585
R693 B.n305 B.n304 585
R694 B.n303 B.n302 585
R695 B.n301 B.n300 585
R696 B.n299 B.n298 585
R697 B.n297 B.n296 585
R698 B.n295 B.n294 585
R699 B.n293 B.n292 585
R700 B.n291 B.n290 585
R701 B.n289 B.n288 585
R702 B.n287 B.n286 585
R703 B.n285 B.n284 585
R704 B.n283 B.n282 585
R705 B.n281 B.n280 585
R706 B.n279 B.n278 585
R707 B.n277 B.n276 585
R708 B.n275 B.n274 585
R709 B.n273 B.n272 585
R710 B.n271 B.n270 585
R711 B.n269 B.n268 585
R712 B.n267 B.n266 585
R713 B.n265 B.n264 585
R714 B.n263 B.n262 585
R715 B.n261 B.n260 585
R716 B.n259 B.n258 585
R717 B.n257 B.n256 585
R718 B.n255 B.n254 585
R719 B.n253 B.n252 585
R720 B.n251 B.n250 585
R721 B.n249 B.n248 585
R722 B.n247 B.n246 585
R723 B.n245 B.n244 585
R724 B.n243 B.n242 585
R725 B.n241 B.n240 585
R726 B.n239 B.n238 585
R727 B.n237 B.n236 585
R728 B.n235 B.n234 585
R729 B.n233 B.n232 585
R730 B.n230 B.n229 585
R731 B.n228 B.n227 585
R732 B.n226 B.n225 585
R733 B.n224 B.n223 585
R734 B.n222 B.n221 585
R735 B.n220 B.n219 585
R736 B.n218 B.n217 585
R737 B.n216 B.n215 585
R738 B.n214 B.n213 585
R739 B.n212 B.n211 585
R740 B.n210 B.n209 585
R741 B.n208 B.n207 585
R742 B.n206 B.n205 585
R743 B.n204 B.n203 585
R744 B.n202 B.n201 585
R745 B.n200 B.n199 585
R746 B.n198 B.n197 585
R747 B.n196 B.n195 585
R748 B.n194 B.n193 585
R749 B.n192 B.n191 585
R750 B.n190 B.n189 585
R751 B.n188 B.n187 585
R752 B.n186 B.n185 585
R753 B.n184 B.n183 585
R754 B.n182 B.n181 585
R755 B.n180 B.n179 585
R756 B.n178 B.n177 585
R757 B.n176 B.n175 585
R758 B.n174 B.n173 585
R759 B.n172 B.n171 585
R760 B.n170 B.n169 585
R761 B.n168 B.n167 585
R762 B.n166 B.n165 585
R763 B.n164 B.n163 585
R764 B.n162 B.n161 585
R765 B.n160 B.n159 585
R766 B.n158 B.n157 585
R767 B.n156 B.n155 585
R768 B.n154 B.n153 585
R769 B.n152 B.n151 585
R770 B.n150 B.n149 585
R771 B.n148 B.n147 585
R772 B.n146 B.n145 585
R773 B.n144 B.n143 585
R774 B.n142 B.n141 585
R775 B.n140 B.n139 585
R776 B.n138 B.n137 585
R777 B.n136 B.n135 585
R778 B.n134 B.n133 585
R779 B.n132 B.n131 585
R780 B.n130 B.n129 585
R781 B.n805 B.n76 585
R782 B.n809 B.n76 585
R783 B.n804 B.n75 585
R784 B.n810 B.n75 585
R785 B.n803 B.n802 585
R786 B.n802 B.n71 585
R787 B.n801 B.n70 585
R788 B.n816 B.n70 585
R789 B.n800 B.n69 585
R790 B.n817 B.n69 585
R791 B.n799 B.n68 585
R792 B.n818 B.n68 585
R793 B.n798 B.n797 585
R794 B.n797 B.n64 585
R795 B.n796 B.n63 585
R796 B.n824 B.n63 585
R797 B.n795 B.n62 585
R798 B.n825 B.n62 585
R799 B.n794 B.n61 585
R800 B.n826 B.n61 585
R801 B.n793 B.n792 585
R802 B.n792 B.n57 585
R803 B.n791 B.n56 585
R804 B.n832 B.n56 585
R805 B.n790 B.n55 585
R806 B.n833 B.n55 585
R807 B.n789 B.n54 585
R808 B.n834 B.n54 585
R809 B.n788 B.n787 585
R810 B.n787 B.n50 585
R811 B.n786 B.n49 585
R812 B.n840 B.n49 585
R813 B.n785 B.n48 585
R814 B.n841 B.n48 585
R815 B.n784 B.n47 585
R816 B.n842 B.n47 585
R817 B.n783 B.n782 585
R818 B.n782 B.n46 585
R819 B.n781 B.n42 585
R820 B.n848 B.n42 585
R821 B.n780 B.n41 585
R822 B.n849 B.n41 585
R823 B.n779 B.n40 585
R824 B.n850 B.n40 585
R825 B.n778 B.n777 585
R826 B.n777 B.n36 585
R827 B.n776 B.n35 585
R828 B.n856 B.n35 585
R829 B.n775 B.n34 585
R830 B.n857 B.n34 585
R831 B.n774 B.n33 585
R832 B.n858 B.n33 585
R833 B.n773 B.n772 585
R834 B.n772 B.n29 585
R835 B.n771 B.n28 585
R836 B.n864 B.n28 585
R837 B.n770 B.n27 585
R838 B.n865 B.n27 585
R839 B.n769 B.n26 585
R840 B.n866 B.n26 585
R841 B.n768 B.n767 585
R842 B.n767 B.n22 585
R843 B.n766 B.n21 585
R844 B.n872 B.n21 585
R845 B.n765 B.n20 585
R846 B.n873 B.n20 585
R847 B.n764 B.n19 585
R848 B.n874 B.n19 585
R849 B.n763 B.n762 585
R850 B.n762 B.n15 585
R851 B.n761 B.n14 585
R852 B.n880 B.n14 585
R853 B.n760 B.n13 585
R854 B.n881 B.n13 585
R855 B.n759 B.n12 585
R856 B.n882 B.n12 585
R857 B.n758 B.n757 585
R858 B.n757 B.n8 585
R859 B.n756 B.n7 585
R860 B.n888 B.n7 585
R861 B.n755 B.n6 585
R862 B.n889 B.n6 585
R863 B.n754 B.n5 585
R864 B.n890 B.n5 585
R865 B.n753 B.n752 585
R866 B.n752 B.n4 585
R867 B.n751 B.n313 585
R868 B.n751 B.n750 585
R869 B.n741 B.n314 585
R870 B.n315 B.n314 585
R871 B.n743 B.n742 585
R872 B.n744 B.n743 585
R873 B.n740 B.n320 585
R874 B.n320 B.n319 585
R875 B.n739 B.n738 585
R876 B.n738 B.n737 585
R877 B.n322 B.n321 585
R878 B.n323 B.n322 585
R879 B.n730 B.n729 585
R880 B.n731 B.n730 585
R881 B.n728 B.n328 585
R882 B.n328 B.n327 585
R883 B.n727 B.n726 585
R884 B.n726 B.n725 585
R885 B.n330 B.n329 585
R886 B.n331 B.n330 585
R887 B.n718 B.n717 585
R888 B.n719 B.n718 585
R889 B.n716 B.n336 585
R890 B.n336 B.n335 585
R891 B.n715 B.n714 585
R892 B.n714 B.n713 585
R893 B.n338 B.n337 585
R894 B.n339 B.n338 585
R895 B.n706 B.n705 585
R896 B.n707 B.n706 585
R897 B.n704 B.n344 585
R898 B.n344 B.n343 585
R899 B.n703 B.n702 585
R900 B.n702 B.n701 585
R901 B.n346 B.n345 585
R902 B.n347 B.n346 585
R903 B.n694 B.n693 585
R904 B.n695 B.n694 585
R905 B.n692 B.n352 585
R906 B.n352 B.n351 585
R907 B.n691 B.n690 585
R908 B.n690 B.n689 585
R909 B.n354 B.n353 585
R910 B.n682 B.n354 585
R911 B.n681 B.n680 585
R912 B.n683 B.n681 585
R913 B.n679 B.n359 585
R914 B.n359 B.n358 585
R915 B.n678 B.n677 585
R916 B.n677 B.n676 585
R917 B.n361 B.n360 585
R918 B.n362 B.n361 585
R919 B.n669 B.n668 585
R920 B.n670 B.n669 585
R921 B.n667 B.n367 585
R922 B.n367 B.n366 585
R923 B.n666 B.n665 585
R924 B.n665 B.n664 585
R925 B.n369 B.n368 585
R926 B.n370 B.n369 585
R927 B.n657 B.n656 585
R928 B.n658 B.n657 585
R929 B.n655 B.n375 585
R930 B.n375 B.n374 585
R931 B.n654 B.n653 585
R932 B.n653 B.n652 585
R933 B.n377 B.n376 585
R934 B.n378 B.n377 585
R935 B.n645 B.n644 585
R936 B.n646 B.n645 585
R937 B.n643 B.n383 585
R938 B.n383 B.n382 585
R939 B.n642 B.n641 585
R940 B.n641 B.n640 585
R941 B.n385 B.n384 585
R942 B.n386 B.n385 585
R943 B.n633 B.n632 585
R944 B.n634 B.n633 585
R945 B.n631 B.n391 585
R946 B.n391 B.n390 585
R947 B.n625 B.n624 585
R948 B.n623 B.n439 585
R949 B.n622 B.n438 585
R950 B.n627 B.n438 585
R951 B.n621 B.n620 585
R952 B.n619 B.n618 585
R953 B.n617 B.n616 585
R954 B.n615 B.n614 585
R955 B.n613 B.n612 585
R956 B.n611 B.n610 585
R957 B.n609 B.n608 585
R958 B.n607 B.n606 585
R959 B.n605 B.n604 585
R960 B.n603 B.n602 585
R961 B.n601 B.n600 585
R962 B.n599 B.n598 585
R963 B.n597 B.n596 585
R964 B.n595 B.n594 585
R965 B.n593 B.n592 585
R966 B.n591 B.n590 585
R967 B.n589 B.n588 585
R968 B.n587 B.n586 585
R969 B.n585 B.n584 585
R970 B.n583 B.n582 585
R971 B.n581 B.n580 585
R972 B.n579 B.n578 585
R973 B.n577 B.n576 585
R974 B.n575 B.n574 585
R975 B.n573 B.n572 585
R976 B.n571 B.n570 585
R977 B.n569 B.n568 585
R978 B.n567 B.n566 585
R979 B.n565 B.n564 585
R980 B.n563 B.n562 585
R981 B.n561 B.n560 585
R982 B.n559 B.n558 585
R983 B.n557 B.n556 585
R984 B.n555 B.n554 585
R985 B.n553 B.n552 585
R986 B.n551 B.n550 585
R987 B.n549 B.n548 585
R988 B.n547 B.n546 585
R989 B.n545 B.n544 585
R990 B.n542 B.n541 585
R991 B.n540 B.n539 585
R992 B.n538 B.n537 585
R993 B.n536 B.n535 585
R994 B.n534 B.n533 585
R995 B.n532 B.n531 585
R996 B.n530 B.n529 585
R997 B.n528 B.n527 585
R998 B.n526 B.n525 585
R999 B.n524 B.n523 585
R1000 B.n522 B.n521 585
R1001 B.n520 B.n519 585
R1002 B.n518 B.n517 585
R1003 B.n516 B.n515 585
R1004 B.n514 B.n513 585
R1005 B.n512 B.n511 585
R1006 B.n510 B.n509 585
R1007 B.n508 B.n507 585
R1008 B.n506 B.n505 585
R1009 B.n504 B.n503 585
R1010 B.n502 B.n501 585
R1011 B.n500 B.n499 585
R1012 B.n498 B.n497 585
R1013 B.n496 B.n495 585
R1014 B.n494 B.n493 585
R1015 B.n492 B.n491 585
R1016 B.n490 B.n489 585
R1017 B.n488 B.n487 585
R1018 B.n486 B.n485 585
R1019 B.n484 B.n483 585
R1020 B.n482 B.n481 585
R1021 B.n480 B.n479 585
R1022 B.n478 B.n477 585
R1023 B.n476 B.n475 585
R1024 B.n474 B.n473 585
R1025 B.n472 B.n471 585
R1026 B.n470 B.n469 585
R1027 B.n468 B.n467 585
R1028 B.n466 B.n465 585
R1029 B.n464 B.n463 585
R1030 B.n462 B.n461 585
R1031 B.n460 B.n459 585
R1032 B.n458 B.n457 585
R1033 B.n456 B.n455 585
R1034 B.n454 B.n453 585
R1035 B.n452 B.n451 585
R1036 B.n450 B.n449 585
R1037 B.n448 B.n447 585
R1038 B.n446 B.n445 585
R1039 B.n393 B.n392 585
R1040 B.n630 B.n629 585
R1041 B.n389 B.n388 585
R1042 B.n390 B.n389 585
R1043 B.n636 B.n635 585
R1044 B.n635 B.n634 585
R1045 B.n637 B.n387 585
R1046 B.n387 B.n386 585
R1047 B.n639 B.n638 585
R1048 B.n640 B.n639 585
R1049 B.n381 B.n380 585
R1050 B.n382 B.n381 585
R1051 B.n648 B.n647 585
R1052 B.n647 B.n646 585
R1053 B.n649 B.n379 585
R1054 B.n379 B.n378 585
R1055 B.n651 B.n650 585
R1056 B.n652 B.n651 585
R1057 B.n373 B.n372 585
R1058 B.n374 B.n373 585
R1059 B.n660 B.n659 585
R1060 B.n659 B.n658 585
R1061 B.n661 B.n371 585
R1062 B.n371 B.n370 585
R1063 B.n663 B.n662 585
R1064 B.n664 B.n663 585
R1065 B.n365 B.n364 585
R1066 B.n366 B.n365 585
R1067 B.n672 B.n671 585
R1068 B.n671 B.n670 585
R1069 B.n673 B.n363 585
R1070 B.n363 B.n362 585
R1071 B.n675 B.n674 585
R1072 B.n676 B.n675 585
R1073 B.n357 B.n356 585
R1074 B.n358 B.n357 585
R1075 B.n685 B.n684 585
R1076 B.n684 B.n683 585
R1077 B.n686 B.n355 585
R1078 B.n682 B.n355 585
R1079 B.n688 B.n687 585
R1080 B.n689 B.n688 585
R1081 B.n350 B.n349 585
R1082 B.n351 B.n350 585
R1083 B.n697 B.n696 585
R1084 B.n696 B.n695 585
R1085 B.n698 B.n348 585
R1086 B.n348 B.n347 585
R1087 B.n700 B.n699 585
R1088 B.n701 B.n700 585
R1089 B.n342 B.n341 585
R1090 B.n343 B.n342 585
R1091 B.n709 B.n708 585
R1092 B.n708 B.n707 585
R1093 B.n710 B.n340 585
R1094 B.n340 B.n339 585
R1095 B.n712 B.n711 585
R1096 B.n713 B.n712 585
R1097 B.n334 B.n333 585
R1098 B.n335 B.n334 585
R1099 B.n721 B.n720 585
R1100 B.n720 B.n719 585
R1101 B.n722 B.n332 585
R1102 B.n332 B.n331 585
R1103 B.n724 B.n723 585
R1104 B.n725 B.n724 585
R1105 B.n326 B.n325 585
R1106 B.n327 B.n326 585
R1107 B.n733 B.n732 585
R1108 B.n732 B.n731 585
R1109 B.n734 B.n324 585
R1110 B.n324 B.n323 585
R1111 B.n736 B.n735 585
R1112 B.n737 B.n736 585
R1113 B.n318 B.n317 585
R1114 B.n319 B.n318 585
R1115 B.n746 B.n745 585
R1116 B.n745 B.n744 585
R1117 B.n747 B.n316 585
R1118 B.n316 B.n315 585
R1119 B.n749 B.n748 585
R1120 B.n750 B.n749 585
R1121 B.n2 B.n0 585
R1122 B.n4 B.n2 585
R1123 B.n3 B.n1 585
R1124 B.n889 B.n3 585
R1125 B.n887 B.n886 585
R1126 B.n888 B.n887 585
R1127 B.n885 B.n9 585
R1128 B.n9 B.n8 585
R1129 B.n884 B.n883 585
R1130 B.n883 B.n882 585
R1131 B.n11 B.n10 585
R1132 B.n881 B.n11 585
R1133 B.n879 B.n878 585
R1134 B.n880 B.n879 585
R1135 B.n877 B.n16 585
R1136 B.n16 B.n15 585
R1137 B.n876 B.n875 585
R1138 B.n875 B.n874 585
R1139 B.n18 B.n17 585
R1140 B.n873 B.n18 585
R1141 B.n871 B.n870 585
R1142 B.n872 B.n871 585
R1143 B.n869 B.n23 585
R1144 B.n23 B.n22 585
R1145 B.n868 B.n867 585
R1146 B.n867 B.n866 585
R1147 B.n25 B.n24 585
R1148 B.n865 B.n25 585
R1149 B.n863 B.n862 585
R1150 B.n864 B.n863 585
R1151 B.n861 B.n30 585
R1152 B.n30 B.n29 585
R1153 B.n860 B.n859 585
R1154 B.n859 B.n858 585
R1155 B.n32 B.n31 585
R1156 B.n857 B.n32 585
R1157 B.n855 B.n854 585
R1158 B.n856 B.n855 585
R1159 B.n853 B.n37 585
R1160 B.n37 B.n36 585
R1161 B.n852 B.n851 585
R1162 B.n851 B.n850 585
R1163 B.n39 B.n38 585
R1164 B.n849 B.n39 585
R1165 B.n847 B.n846 585
R1166 B.n848 B.n847 585
R1167 B.n845 B.n43 585
R1168 B.n46 B.n43 585
R1169 B.n844 B.n843 585
R1170 B.n843 B.n842 585
R1171 B.n45 B.n44 585
R1172 B.n841 B.n45 585
R1173 B.n839 B.n838 585
R1174 B.n840 B.n839 585
R1175 B.n837 B.n51 585
R1176 B.n51 B.n50 585
R1177 B.n836 B.n835 585
R1178 B.n835 B.n834 585
R1179 B.n53 B.n52 585
R1180 B.n833 B.n53 585
R1181 B.n831 B.n830 585
R1182 B.n832 B.n831 585
R1183 B.n829 B.n58 585
R1184 B.n58 B.n57 585
R1185 B.n828 B.n827 585
R1186 B.n827 B.n826 585
R1187 B.n60 B.n59 585
R1188 B.n825 B.n60 585
R1189 B.n823 B.n822 585
R1190 B.n824 B.n823 585
R1191 B.n821 B.n65 585
R1192 B.n65 B.n64 585
R1193 B.n820 B.n819 585
R1194 B.n819 B.n818 585
R1195 B.n67 B.n66 585
R1196 B.n817 B.n67 585
R1197 B.n815 B.n814 585
R1198 B.n816 B.n815 585
R1199 B.n813 B.n72 585
R1200 B.n72 B.n71 585
R1201 B.n812 B.n811 585
R1202 B.n811 B.n810 585
R1203 B.n74 B.n73 585
R1204 B.n809 B.n74 585
R1205 B.n892 B.n891 585
R1206 B.n891 B.n890 585
R1207 B.n625 B.n389 449.257
R1208 B.n129 B.n74 449.257
R1209 B.n629 B.n391 449.257
R1210 B.n807 B.n76 449.257
R1211 B.n442 B.t9 335.147
R1212 B.n124 B.t12 335.147
R1213 B.n440 B.t16 335.147
R1214 B.n126 B.t18 335.147
R1215 B.n442 B.t6 324.897
R1216 B.n440 B.t14 324.897
R1217 B.n126 B.t17 324.897
R1218 B.n124 B.t10 324.897
R1219 B.n443 B.t8 281.038
R1220 B.n125 B.t13 281.038
R1221 B.n441 B.t15 281.038
R1222 B.n127 B.t19 281.038
R1223 B.n808 B.n122 256.663
R1224 B.n808 B.n121 256.663
R1225 B.n808 B.n120 256.663
R1226 B.n808 B.n119 256.663
R1227 B.n808 B.n118 256.663
R1228 B.n808 B.n117 256.663
R1229 B.n808 B.n116 256.663
R1230 B.n808 B.n115 256.663
R1231 B.n808 B.n114 256.663
R1232 B.n808 B.n113 256.663
R1233 B.n808 B.n112 256.663
R1234 B.n808 B.n111 256.663
R1235 B.n808 B.n110 256.663
R1236 B.n808 B.n109 256.663
R1237 B.n808 B.n108 256.663
R1238 B.n808 B.n107 256.663
R1239 B.n808 B.n106 256.663
R1240 B.n808 B.n105 256.663
R1241 B.n808 B.n104 256.663
R1242 B.n808 B.n103 256.663
R1243 B.n808 B.n102 256.663
R1244 B.n808 B.n101 256.663
R1245 B.n808 B.n100 256.663
R1246 B.n808 B.n99 256.663
R1247 B.n808 B.n98 256.663
R1248 B.n808 B.n97 256.663
R1249 B.n808 B.n96 256.663
R1250 B.n808 B.n95 256.663
R1251 B.n808 B.n94 256.663
R1252 B.n808 B.n93 256.663
R1253 B.n808 B.n92 256.663
R1254 B.n808 B.n91 256.663
R1255 B.n808 B.n90 256.663
R1256 B.n808 B.n89 256.663
R1257 B.n808 B.n88 256.663
R1258 B.n808 B.n87 256.663
R1259 B.n808 B.n86 256.663
R1260 B.n808 B.n85 256.663
R1261 B.n808 B.n84 256.663
R1262 B.n808 B.n83 256.663
R1263 B.n808 B.n82 256.663
R1264 B.n808 B.n81 256.663
R1265 B.n808 B.n80 256.663
R1266 B.n808 B.n79 256.663
R1267 B.n808 B.n78 256.663
R1268 B.n808 B.n77 256.663
R1269 B.n627 B.n626 256.663
R1270 B.n627 B.n394 256.663
R1271 B.n627 B.n395 256.663
R1272 B.n627 B.n396 256.663
R1273 B.n627 B.n397 256.663
R1274 B.n627 B.n398 256.663
R1275 B.n627 B.n399 256.663
R1276 B.n627 B.n400 256.663
R1277 B.n627 B.n401 256.663
R1278 B.n627 B.n402 256.663
R1279 B.n627 B.n403 256.663
R1280 B.n627 B.n404 256.663
R1281 B.n627 B.n405 256.663
R1282 B.n627 B.n406 256.663
R1283 B.n627 B.n407 256.663
R1284 B.n627 B.n408 256.663
R1285 B.n627 B.n409 256.663
R1286 B.n627 B.n410 256.663
R1287 B.n627 B.n411 256.663
R1288 B.n627 B.n412 256.663
R1289 B.n627 B.n413 256.663
R1290 B.n627 B.n414 256.663
R1291 B.n627 B.n415 256.663
R1292 B.n627 B.n416 256.663
R1293 B.n627 B.n417 256.663
R1294 B.n627 B.n418 256.663
R1295 B.n627 B.n419 256.663
R1296 B.n627 B.n420 256.663
R1297 B.n627 B.n421 256.663
R1298 B.n627 B.n422 256.663
R1299 B.n627 B.n423 256.663
R1300 B.n627 B.n424 256.663
R1301 B.n627 B.n425 256.663
R1302 B.n627 B.n426 256.663
R1303 B.n627 B.n427 256.663
R1304 B.n627 B.n428 256.663
R1305 B.n627 B.n429 256.663
R1306 B.n627 B.n430 256.663
R1307 B.n627 B.n431 256.663
R1308 B.n627 B.n432 256.663
R1309 B.n627 B.n433 256.663
R1310 B.n627 B.n434 256.663
R1311 B.n627 B.n435 256.663
R1312 B.n627 B.n436 256.663
R1313 B.n627 B.n437 256.663
R1314 B.n628 B.n627 256.663
R1315 B.n635 B.n389 163.367
R1316 B.n635 B.n387 163.367
R1317 B.n639 B.n387 163.367
R1318 B.n639 B.n381 163.367
R1319 B.n647 B.n381 163.367
R1320 B.n647 B.n379 163.367
R1321 B.n651 B.n379 163.367
R1322 B.n651 B.n373 163.367
R1323 B.n659 B.n373 163.367
R1324 B.n659 B.n371 163.367
R1325 B.n663 B.n371 163.367
R1326 B.n663 B.n365 163.367
R1327 B.n671 B.n365 163.367
R1328 B.n671 B.n363 163.367
R1329 B.n675 B.n363 163.367
R1330 B.n675 B.n357 163.367
R1331 B.n684 B.n357 163.367
R1332 B.n684 B.n355 163.367
R1333 B.n688 B.n355 163.367
R1334 B.n688 B.n350 163.367
R1335 B.n696 B.n350 163.367
R1336 B.n696 B.n348 163.367
R1337 B.n700 B.n348 163.367
R1338 B.n700 B.n342 163.367
R1339 B.n708 B.n342 163.367
R1340 B.n708 B.n340 163.367
R1341 B.n712 B.n340 163.367
R1342 B.n712 B.n334 163.367
R1343 B.n720 B.n334 163.367
R1344 B.n720 B.n332 163.367
R1345 B.n724 B.n332 163.367
R1346 B.n724 B.n326 163.367
R1347 B.n732 B.n326 163.367
R1348 B.n732 B.n324 163.367
R1349 B.n736 B.n324 163.367
R1350 B.n736 B.n318 163.367
R1351 B.n745 B.n318 163.367
R1352 B.n745 B.n316 163.367
R1353 B.n749 B.n316 163.367
R1354 B.n749 B.n2 163.367
R1355 B.n891 B.n2 163.367
R1356 B.n891 B.n3 163.367
R1357 B.n887 B.n3 163.367
R1358 B.n887 B.n9 163.367
R1359 B.n883 B.n9 163.367
R1360 B.n883 B.n11 163.367
R1361 B.n879 B.n11 163.367
R1362 B.n879 B.n16 163.367
R1363 B.n875 B.n16 163.367
R1364 B.n875 B.n18 163.367
R1365 B.n871 B.n18 163.367
R1366 B.n871 B.n23 163.367
R1367 B.n867 B.n23 163.367
R1368 B.n867 B.n25 163.367
R1369 B.n863 B.n25 163.367
R1370 B.n863 B.n30 163.367
R1371 B.n859 B.n30 163.367
R1372 B.n859 B.n32 163.367
R1373 B.n855 B.n32 163.367
R1374 B.n855 B.n37 163.367
R1375 B.n851 B.n37 163.367
R1376 B.n851 B.n39 163.367
R1377 B.n847 B.n39 163.367
R1378 B.n847 B.n43 163.367
R1379 B.n843 B.n43 163.367
R1380 B.n843 B.n45 163.367
R1381 B.n839 B.n45 163.367
R1382 B.n839 B.n51 163.367
R1383 B.n835 B.n51 163.367
R1384 B.n835 B.n53 163.367
R1385 B.n831 B.n53 163.367
R1386 B.n831 B.n58 163.367
R1387 B.n827 B.n58 163.367
R1388 B.n827 B.n60 163.367
R1389 B.n823 B.n60 163.367
R1390 B.n823 B.n65 163.367
R1391 B.n819 B.n65 163.367
R1392 B.n819 B.n67 163.367
R1393 B.n815 B.n67 163.367
R1394 B.n815 B.n72 163.367
R1395 B.n811 B.n72 163.367
R1396 B.n811 B.n74 163.367
R1397 B.n439 B.n438 163.367
R1398 B.n620 B.n438 163.367
R1399 B.n618 B.n617 163.367
R1400 B.n614 B.n613 163.367
R1401 B.n610 B.n609 163.367
R1402 B.n606 B.n605 163.367
R1403 B.n602 B.n601 163.367
R1404 B.n598 B.n597 163.367
R1405 B.n594 B.n593 163.367
R1406 B.n590 B.n589 163.367
R1407 B.n586 B.n585 163.367
R1408 B.n582 B.n581 163.367
R1409 B.n578 B.n577 163.367
R1410 B.n574 B.n573 163.367
R1411 B.n570 B.n569 163.367
R1412 B.n566 B.n565 163.367
R1413 B.n562 B.n561 163.367
R1414 B.n558 B.n557 163.367
R1415 B.n554 B.n553 163.367
R1416 B.n550 B.n549 163.367
R1417 B.n546 B.n545 163.367
R1418 B.n541 B.n540 163.367
R1419 B.n537 B.n536 163.367
R1420 B.n533 B.n532 163.367
R1421 B.n529 B.n528 163.367
R1422 B.n525 B.n524 163.367
R1423 B.n521 B.n520 163.367
R1424 B.n517 B.n516 163.367
R1425 B.n513 B.n512 163.367
R1426 B.n509 B.n508 163.367
R1427 B.n505 B.n504 163.367
R1428 B.n501 B.n500 163.367
R1429 B.n497 B.n496 163.367
R1430 B.n493 B.n492 163.367
R1431 B.n489 B.n488 163.367
R1432 B.n485 B.n484 163.367
R1433 B.n481 B.n480 163.367
R1434 B.n477 B.n476 163.367
R1435 B.n473 B.n472 163.367
R1436 B.n469 B.n468 163.367
R1437 B.n465 B.n464 163.367
R1438 B.n461 B.n460 163.367
R1439 B.n457 B.n456 163.367
R1440 B.n453 B.n452 163.367
R1441 B.n449 B.n448 163.367
R1442 B.n445 B.n393 163.367
R1443 B.n633 B.n391 163.367
R1444 B.n633 B.n385 163.367
R1445 B.n641 B.n385 163.367
R1446 B.n641 B.n383 163.367
R1447 B.n645 B.n383 163.367
R1448 B.n645 B.n377 163.367
R1449 B.n653 B.n377 163.367
R1450 B.n653 B.n375 163.367
R1451 B.n657 B.n375 163.367
R1452 B.n657 B.n369 163.367
R1453 B.n665 B.n369 163.367
R1454 B.n665 B.n367 163.367
R1455 B.n669 B.n367 163.367
R1456 B.n669 B.n361 163.367
R1457 B.n677 B.n361 163.367
R1458 B.n677 B.n359 163.367
R1459 B.n681 B.n359 163.367
R1460 B.n681 B.n354 163.367
R1461 B.n690 B.n354 163.367
R1462 B.n690 B.n352 163.367
R1463 B.n694 B.n352 163.367
R1464 B.n694 B.n346 163.367
R1465 B.n702 B.n346 163.367
R1466 B.n702 B.n344 163.367
R1467 B.n706 B.n344 163.367
R1468 B.n706 B.n338 163.367
R1469 B.n714 B.n338 163.367
R1470 B.n714 B.n336 163.367
R1471 B.n718 B.n336 163.367
R1472 B.n718 B.n330 163.367
R1473 B.n726 B.n330 163.367
R1474 B.n726 B.n328 163.367
R1475 B.n730 B.n328 163.367
R1476 B.n730 B.n322 163.367
R1477 B.n738 B.n322 163.367
R1478 B.n738 B.n320 163.367
R1479 B.n743 B.n320 163.367
R1480 B.n743 B.n314 163.367
R1481 B.n751 B.n314 163.367
R1482 B.n752 B.n751 163.367
R1483 B.n752 B.n5 163.367
R1484 B.n6 B.n5 163.367
R1485 B.n7 B.n6 163.367
R1486 B.n757 B.n7 163.367
R1487 B.n757 B.n12 163.367
R1488 B.n13 B.n12 163.367
R1489 B.n14 B.n13 163.367
R1490 B.n762 B.n14 163.367
R1491 B.n762 B.n19 163.367
R1492 B.n20 B.n19 163.367
R1493 B.n21 B.n20 163.367
R1494 B.n767 B.n21 163.367
R1495 B.n767 B.n26 163.367
R1496 B.n27 B.n26 163.367
R1497 B.n28 B.n27 163.367
R1498 B.n772 B.n28 163.367
R1499 B.n772 B.n33 163.367
R1500 B.n34 B.n33 163.367
R1501 B.n35 B.n34 163.367
R1502 B.n777 B.n35 163.367
R1503 B.n777 B.n40 163.367
R1504 B.n41 B.n40 163.367
R1505 B.n42 B.n41 163.367
R1506 B.n782 B.n42 163.367
R1507 B.n782 B.n47 163.367
R1508 B.n48 B.n47 163.367
R1509 B.n49 B.n48 163.367
R1510 B.n787 B.n49 163.367
R1511 B.n787 B.n54 163.367
R1512 B.n55 B.n54 163.367
R1513 B.n56 B.n55 163.367
R1514 B.n792 B.n56 163.367
R1515 B.n792 B.n61 163.367
R1516 B.n62 B.n61 163.367
R1517 B.n63 B.n62 163.367
R1518 B.n797 B.n63 163.367
R1519 B.n797 B.n68 163.367
R1520 B.n69 B.n68 163.367
R1521 B.n70 B.n69 163.367
R1522 B.n802 B.n70 163.367
R1523 B.n802 B.n75 163.367
R1524 B.n76 B.n75 163.367
R1525 B.n133 B.n132 163.367
R1526 B.n137 B.n136 163.367
R1527 B.n141 B.n140 163.367
R1528 B.n145 B.n144 163.367
R1529 B.n149 B.n148 163.367
R1530 B.n153 B.n152 163.367
R1531 B.n157 B.n156 163.367
R1532 B.n161 B.n160 163.367
R1533 B.n165 B.n164 163.367
R1534 B.n169 B.n168 163.367
R1535 B.n173 B.n172 163.367
R1536 B.n177 B.n176 163.367
R1537 B.n181 B.n180 163.367
R1538 B.n185 B.n184 163.367
R1539 B.n189 B.n188 163.367
R1540 B.n193 B.n192 163.367
R1541 B.n197 B.n196 163.367
R1542 B.n201 B.n200 163.367
R1543 B.n205 B.n204 163.367
R1544 B.n209 B.n208 163.367
R1545 B.n213 B.n212 163.367
R1546 B.n217 B.n216 163.367
R1547 B.n221 B.n220 163.367
R1548 B.n225 B.n224 163.367
R1549 B.n229 B.n228 163.367
R1550 B.n234 B.n233 163.367
R1551 B.n238 B.n237 163.367
R1552 B.n242 B.n241 163.367
R1553 B.n246 B.n245 163.367
R1554 B.n250 B.n249 163.367
R1555 B.n254 B.n253 163.367
R1556 B.n258 B.n257 163.367
R1557 B.n262 B.n261 163.367
R1558 B.n266 B.n265 163.367
R1559 B.n270 B.n269 163.367
R1560 B.n274 B.n273 163.367
R1561 B.n278 B.n277 163.367
R1562 B.n282 B.n281 163.367
R1563 B.n286 B.n285 163.367
R1564 B.n290 B.n289 163.367
R1565 B.n294 B.n293 163.367
R1566 B.n298 B.n297 163.367
R1567 B.n302 B.n301 163.367
R1568 B.n306 B.n305 163.367
R1569 B.n310 B.n309 163.367
R1570 B.n807 B.n123 163.367
R1571 B.n627 B.n390 75.9947
R1572 B.n809 B.n808 75.9947
R1573 B.n626 B.n625 71.676
R1574 B.n620 B.n394 71.676
R1575 B.n617 B.n395 71.676
R1576 B.n613 B.n396 71.676
R1577 B.n609 B.n397 71.676
R1578 B.n605 B.n398 71.676
R1579 B.n601 B.n399 71.676
R1580 B.n597 B.n400 71.676
R1581 B.n593 B.n401 71.676
R1582 B.n589 B.n402 71.676
R1583 B.n585 B.n403 71.676
R1584 B.n581 B.n404 71.676
R1585 B.n577 B.n405 71.676
R1586 B.n573 B.n406 71.676
R1587 B.n569 B.n407 71.676
R1588 B.n565 B.n408 71.676
R1589 B.n561 B.n409 71.676
R1590 B.n557 B.n410 71.676
R1591 B.n553 B.n411 71.676
R1592 B.n549 B.n412 71.676
R1593 B.n545 B.n413 71.676
R1594 B.n540 B.n414 71.676
R1595 B.n536 B.n415 71.676
R1596 B.n532 B.n416 71.676
R1597 B.n528 B.n417 71.676
R1598 B.n524 B.n418 71.676
R1599 B.n520 B.n419 71.676
R1600 B.n516 B.n420 71.676
R1601 B.n512 B.n421 71.676
R1602 B.n508 B.n422 71.676
R1603 B.n504 B.n423 71.676
R1604 B.n500 B.n424 71.676
R1605 B.n496 B.n425 71.676
R1606 B.n492 B.n426 71.676
R1607 B.n488 B.n427 71.676
R1608 B.n484 B.n428 71.676
R1609 B.n480 B.n429 71.676
R1610 B.n476 B.n430 71.676
R1611 B.n472 B.n431 71.676
R1612 B.n468 B.n432 71.676
R1613 B.n464 B.n433 71.676
R1614 B.n460 B.n434 71.676
R1615 B.n456 B.n435 71.676
R1616 B.n452 B.n436 71.676
R1617 B.n448 B.n437 71.676
R1618 B.n628 B.n393 71.676
R1619 B.n129 B.n77 71.676
R1620 B.n133 B.n78 71.676
R1621 B.n137 B.n79 71.676
R1622 B.n141 B.n80 71.676
R1623 B.n145 B.n81 71.676
R1624 B.n149 B.n82 71.676
R1625 B.n153 B.n83 71.676
R1626 B.n157 B.n84 71.676
R1627 B.n161 B.n85 71.676
R1628 B.n165 B.n86 71.676
R1629 B.n169 B.n87 71.676
R1630 B.n173 B.n88 71.676
R1631 B.n177 B.n89 71.676
R1632 B.n181 B.n90 71.676
R1633 B.n185 B.n91 71.676
R1634 B.n189 B.n92 71.676
R1635 B.n193 B.n93 71.676
R1636 B.n197 B.n94 71.676
R1637 B.n201 B.n95 71.676
R1638 B.n205 B.n96 71.676
R1639 B.n209 B.n97 71.676
R1640 B.n213 B.n98 71.676
R1641 B.n217 B.n99 71.676
R1642 B.n221 B.n100 71.676
R1643 B.n225 B.n101 71.676
R1644 B.n229 B.n102 71.676
R1645 B.n234 B.n103 71.676
R1646 B.n238 B.n104 71.676
R1647 B.n242 B.n105 71.676
R1648 B.n246 B.n106 71.676
R1649 B.n250 B.n107 71.676
R1650 B.n254 B.n108 71.676
R1651 B.n258 B.n109 71.676
R1652 B.n262 B.n110 71.676
R1653 B.n266 B.n111 71.676
R1654 B.n270 B.n112 71.676
R1655 B.n274 B.n113 71.676
R1656 B.n278 B.n114 71.676
R1657 B.n282 B.n115 71.676
R1658 B.n286 B.n116 71.676
R1659 B.n290 B.n117 71.676
R1660 B.n294 B.n118 71.676
R1661 B.n298 B.n119 71.676
R1662 B.n302 B.n120 71.676
R1663 B.n306 B.n121 71.676
R1664 B.n310 B.n122 71.676
R1665 B.n123 B.n122 71.676
R1666 B.n309 B.n121 71.676
R1667 B.n305 B.n120 71.676
R1668 B.n301 B.n119 71.676
R1669 B.n297 B.n118 71.676
R1670 B.n293 B.n117 71.676
R1671 B.n289 B.n116 71.676
R1672 B.n285 B.n115 71.676
R1673 B.n281 B.n114 71.676
R1674 B.n277 B.n113 71.676
R1675 B.n273 B.n112 71.676
R1676 B.n269 B.n111 71.676
R1677 B.n265 B.n110 71.676
R1678 B.n261 B.n109 71.676
R1679 B.n257 B.n108 71.676
R1680 B.n253 B.n107 71.676
R1681 B.n249 B.n106 71.676
R1682 B.n245 B.n105 71.676
R1683 B.n241 B.n104 71.676
R1684 B.n237 B.n103 71.676
R1685 B.n233 B.n102 71.676
R1686 B.n228 B.n101 71.676
R1687 B.n224 B.n100 71.676
R1688 B.n220 B.n99 71.676
R1689 B.n216 B.n98 71.676
R1690 B.n212 B.n97 71.676
R1691 B.n208 B.n96 71.676
R1692 B.n204 B.n95 71.676
R1693 B.n200 B.n94 71.676
R1694 B.n196 B.n93 71.676
R1695 B.n192 B.n92 71.676
R1696 B.n188 B.n91 71.676
R1697 B.n184 B.n90 71.676
R1698 B.n180 B.n89 71.676
R1699 B.n176 B.n88 71.676
R1700 B.n172 B.n87 71.676
R1701 B.n168 B.n86 71.676
R1702 B.n164 B.n85 71.676
R1703 B.n160 B.n84 71.676
R1704 B.n156 B.n83 71.676
R1705 B.n152 B.n82 71.676
R1706 B.n148 B.n81 71.676
R1707 B.n144 B.n80 71.676
R1708 B.n140 B.n79 71.676
R1709 B.n136 B.n78 71.676
R1710 B.n132 B.n77 71.676
R1711 B.n626 B.n439 71.676
R1712 B.n618 B.n394 71.676
R1713 B.n614 B.n395 71.676
R1714 B.n610 B.n396 71.676
R1715 B.n606 B.n397 71.676
R1716 B.n602 B.n398 71.676
R1717 B.n598 B.n399 71.676
R1718 B.n594 B.n400 71.676
R1719 B.n590 B.n401 71.676
R1720 B.n586 B.n402 71.676
R1721 B.n582 B.n403 71.676
R1722 B.n578 B.n404 71.676
R1723 B.n574 B.n405 71.676
R1724 B.n570 B.n406 71.676
R1725 B.n566 B.n407 71.676
R1726 B.n562 B.n408 71.676
R1727 B.n558 B.n409 71.676
R1728 B.n554 B.n410 71.676
R1729 B.n550 B.n411 71.676
R1730 B.n546 B.n412 71.676
R1731 B.n541 B.n413 71.676
R1732 B.n537 B.n414 71.676
R1733 B.n533 B.n415 71.676
R1734 B.n529 B.n416 71.676
R1735 B.n525 B.n417 71.676
R1736 B.n521 B.n418 71.676
R1737 B.n517 B.n419 71.676
R1738 B.n513 B.n420 71.676
R1739 B.n509 B.n421 71.676
R1740 B.n505 B.n422 71.676
R1741 B.n501 B.n423 71.676
R1742 B.n497 B.n424 71.676
R1743 B.n493 B.n425 71.676
R1744 B.n489 B.n426 71.676
R1745 B.n485 B.n427 71.676
R1746 B.n481 B.n428 71.676
R1747 B.n477 B.n429 71.676
R1748 B.n473 B.n430 71.676
R1749 B.n469 B.n431 71.676
R1750 B.n465 B.n432 71.676
R1751 B.n461 B.n433 71.676
R1752 B.n457 B.n434 71.676
R1753 B.n453 B.n435 71.676
R1754 B.n449 B.n436 71.676
R1755 B.n445 B.n437 71.676
R1756 B.n629 B.n628 71.676
R1757 B.n444 B.n443 59.5399
R1758 B.n543 B.n441 59.5399
R1759 B.n128 B.n127 59.5399
R1760 B.n231 B.n125 59.5399
R1761 B.n443 B.n442 54.1096
R1762 B.n441 B.n440 54.1096
R1763 B.n127 B.n126 54.1096
R1764 B.n125 B.n124 54.1096
R1765 B.n634 B.n390 43.4258
R1766 B.n634 B.n386 43.4258
R1767 B.n640 B.n386 43.4258
R1768 B.n640 B.n382 43.4258
R1769 B.n646 B.n382 43.4258
R1770 B.n646 B.n378 43.4258
R1771 B.n652 B.n378 43.4258
R1772 B.n658 B.n374 43.4258
R1773 B.n658 B.n370 43.4258
R1774 B.n664 B.n370 43.4258
R1775 B.n664 B.n366 43.4258
R1776 B.n670 B.n366 43.4258
R1777 B.n670 B.n362 43.4258
R1778 B.n676 B.n362 43.4258
R1779 B.n676 B.n358 43.4258
R1780 B.n683 B.n358 43.4258
R1781 B.n683 B.n682 43.4258
R1782 B.n689 B.n351 43.4258
R1783 B.n695 B.n351 43.4258
R1784 B.n695 B.n347 43.4258
R1785 B.n701 B.n347 43.4258
R1786 B.n701 B.n343 43.4258
R1787 B.n707 B.n343 43.4258
R1788 B.n707 B.n339 43.4258
R1789 B.n713 B.n339 43.4258
R1790 B.n719 B.n335 43.4258
R1791 B.n719 B.n331 43.4258
R1792 B.n725 B.n331 43.4258
R1793 B.n725 B.n327 43.4258
R1794 B.n731 B.n327 43.4258
R1795 B.n731 B.n323 43.4258
R1796 B.n737 B.n323 43.4258
R1797 B.n744 B.n319 43.4258
R1798 B.n744 B.n315 43.4258
R1799 B.n750 B.n315 43.4258
R1800 B.n750 B.n4 43.4258
R1801 B.n890 B.n4 43.4258
R1802 B.n890 B.n889 43.4258
R1803 B.n889 B.n888 43.4258
R1804 B.n888 B.n8 43.4258
R1805 B.n882 B.n8 43.4258
R1806 B.n882 B.n881 43.4258
R1807 B.n880 B.n15 43.4258
R1808 B.n874 B.n15 43.4258
R1809 B.n874 B.n873 43.4258
R1810 B.n873 B.n872 43.4258
R1811 B.n872 B.n22 43.4258
R1812 B.n866 B.n22 43.4258
R1813 B.n866 B.n865 43.4258
R1814 B.n864 B.n29 43.4258
R1815 B.n858 B.n29 43.4258
R1816 B.n858 B.n857 43.4258
R1817 B.n857 B.n856 43.4258
R1818 B.n856 B.n36 43.4258
R1819 B.n850 B.n36 43.4258
R1820 B.n850 B.n849 43.4258
R1821 B.n849 B.n848 43.4258
R1822 B.n842 B.n46 43.4258
R1823 B.n842 B.n841 43.4258
R1824 B.n841 B.n840 43.4258
R1825 B.n840 B.n50 43.4258
R1826 B.n834 B.n50 43.4258
R1827 B.n834 B.n833 43.4258
R1828 B.n833 B.n832 43.4258
R1829 B.n832 B.n57 43.4258
R1830 B.n826 B.n57 43.4258
R1831 B.n826 B.n825 43.4258
R1832 B.n824 B.n64 43.4258
R1833 B.n818 B.n64 43.4258
R1834 B.n818 B.n817 43.4258
R1835 B.n817 B.n816 43.4258
R1836 B.n816 B.n71 43.4258
R1837 B.n810 B.n71 43.4258
R1838 B.n810 B.n809 43.4258
R1839 B.t2 B.n335 39.5941
R1840 B.n865 B.t5 39.5941
R1841 B.n682 B.t3 38.3169
R1842 B.n46 B.t0 38.3169
R1843 B.t4 B.n319 30.6536
R1844 B.n881 B.t1 30.6536
R1845 B.n806 B.n805 29.1907
R1846 B.n130 B.n73 29.1907
R1847 B.n631 B.n630 29.1907
R1848 B.n624 B.n388 29.1907
R1849 B.t7 B.n374 22.9903
R1850 B.n825 B.t11 22.9903
R1851 B.n652 B.t7 20.4359
R1852 B.t11 B.n824 20.4359
R1853 B B.n892 18.0485
R1854 B.n737 B.t4 12.7726
R1855 B.t1 B.n880 12.7726
R1856 B.n131 B.n130 10.6151
R1857 B.n134 B.n131 10.6151
R1858 B.n135 B.n134 10.6151
R1859 B.n138 B.n135 10.6151
R1860 B.n139 B.n138 10.6151
R1861 B.n142 B.n139 10.6151
R1862 B.n143 B.n142 10.6151
R1863 B.n146 B.n143 10.6151
R1864 B.n147 B.n146 10.6151
R1865 B.n150 B.n147 10.6151
R1866 B.n151 B.n150 10.6151
R1867 B.n154 B.n151 10.6151
R1868 B.n155 B.n154 10.6151
R1869 B.n158 B.n155 10.6151
R1870 B.n159 B.n158 10.6151
R1871 B.n162 B.n159 10.6151
R1872 B.n163 B.n162 10.6151
R1873 B.n166 B.n163 10.6151
R1874 B.n167 B.n166 10.6151
R1875 B.n170 B.n167 10.6151
R1876 B.n171 B.n170 10.6151
R1877 B.n174 B.n171 10.6151
R1878 B.n175 B.n174 10.6151
R1879 B.n178 B.n175 10.6151
R1880 B.n179 B.n178 10.6151
R1881 B.n182 B.n179 10.6151
R1882 B.n183 B.n182 10.6151
R1883 B.n186 B.n183 10.6151
R1884 B.n187 B.n186 10.6151
R1885 B.n190 B.n187 10.6151
R1886 B.n191 B.n190 10.6151
R1887 B.n194 B.n191 10.6151
R1888 B.n195 B.n194 10.6151
R1889 B.n198 B.n195 10.6151
R1890 B.n199 B.n198 10.6151
R1891 B.n202 B.n199 10.6151
R1892 B.n203 B.n202 10.6151
R1893 B.n206 B.n203 10.6151
R1894 B.n207 B.n206 10.6151
R1895 B.n210 B.n207 10.6151
R1896 B.n211 B.n210 10.6151
R1897 B.n215 B.n214 10.6151
R1898 B.n218 B.n215 10.6151
R1899 B.n219 B.n218 10.6151
R1900 B.n222 B.n219 10.6151
R1901 B.n223 B.n222 10.6151
R1902 B.n226 B.n223 10.6151
R1903 B.n227 B.n226 10.6151
R1904 B.n230 B.n227 10.6151
R1905 B.n235 B.n232 10.6151
R1906 B.n236 B.n235 10.6151
R1907 B.n239 B.n236 10.6151
R1908 B.n240 B.n239 10.6151
R1909 B.n243 B.n240 10.6151
R1910 B.n244 B.n243 10.6151
R1911 B.n247 B.n244 10.6151
R1912 B.n248 B.n247 10.6151
R1913 B.n251 B.n248 10.6151
R1914 B.n252 B.n251 10.6151
R1915 B.n255 B.n252 10.6151
R1916 B.n256 B.n255 10.6151
R1917 B.n259 B.n256 10.6151
R1918 B.n260 B.n259 10.6151
R1919 B.n263 B.n260 10.6151
R1920 B.n264 B.n263 10.6151
R1921 B.n267 B.n264 10.6151
R1922 B.n268 B.n267 10.6151
R1923 B.n271 B.n268 10.6151
R1924 B.n272 B.n271 10.6151
R1925 B.n275 B.n272 10.6151
R1926 B.n276 B.n275 10.6151
R1927 B.n279 B.n276 10.6151
R1928 B.n280 B.n279 10.6151
R1929 B.n283 B.n280 10.6151
R1930 B.n284 B.n283 10.6151
R1931 B.n287 B.n284 10.6151
R1932 B.n288 B.n287 10.6151
R1933 B.n291 B.n288 10.6151
R1934 B.n292 B.n291 10.6151
R1935 B.n295 B.n292 10.6151
R1936 B.n296 B.n295 10.6151
R1937 B.n299 B.n296 10.6151
R1938 B.n300 B.n299 10.6151
R1939 B.n303 B.n300 10.6151
R1940 B.n304 B.n303 10.6151
R1941 B.n307 B.n304 10.6151
R1942 B.n308 B.n307 10.6151
R1943 B.n311 B.n308 10.6151
R1944 B.n312 B.n311 10.6151
R1945 B.n806 B.n312 10.6151
R1946 B.n632 B.n631 10.6151
R1947 B.n632 B.n384 10.6151
R1948 B.n642 B.n384 10.6151
R1949 B.n643 B.n642 10.6151
R1950 B.n644 B.n643 10.6151
R1951 B.n644 B.n376 10.6151
R1952 B.n654 B.n376 10.6151
R1953 B.n655 B.n654 10.6151
R1954 B.n656 B.n655 10.6151
R1955 B.n656 B.n368 10.6151
R1956 B.n666 B.n368 10.6151
R1957 B.n667 B.n666 10.6151
R1958 B.n668 B.n667 10.6151
R1959 B.n668 B.n360 10.6151
R1960 B.n678 B.n360 10.6151
R1961 B.n679 B.n678 10.6151
R1962 B.n680 B.n679 10.6151
R1963 B.n680 B.n353 10.6151
R1964 B.n691 B.n353 10.6151
R1965 B.n692 B.n691 10.6151
R1966 B.n693 B.n692 10.6151
R1967 B.n693 B.n345 10.6151
R1968 B.n703 B.n345 10.6151
R1969 B.n704 B.n703 10.6151
R1970 B.n705 B.n704 10.6151
R1971 B.n705 B.n337 10.6151
R1972 B.n715 B.n337 10.6151
R1973 B.n716 B.n715 10.6151
R1974 B.n717 B.n716 10.6151
R1975 B.n717 B.n329 10.6151
R1976 B.n727 B.n329 10.6151
R1977 B.n728 B.n727 10.6151
R1978 B.n729 B.n728 10.6151
R1979 B.n729 B.n321 10.6151
R1980 B.n739 B.n321 10.6151
R1981 B.n740 B.n739 10.6151
R1982 B.n742 B.n740 10.6151
R1983 B.n742 B.n741 10.6151
R1984 B.n741 B.n313 10.6151
R1985 B.n753 B.n313 10.6151
R1986 B.n754 B.n753 10.6151
R1987 B.n755 B.n754 10.6151
R1988 B.n756 B.n755 10.6151
R1989 B.n758 B.n756 10.6151
R1990 B.n759 B.n758 10.6151
R1991 B.n760 B.n759 10.6151
R1992 B.n761 B.n760 10.6151
R1993 B.n763 B.n761 10.6151
R1994 B.n764 B.n763 10.6151
R1995 B.n765 B.n764 10.6151
R1996 B.n766 B.n765 10.6151
R1997 B.n768 B.n766 10.6151
R1998 B.n769 B.n768 10.6151
R1999 B.n770 B.n769 10.6151
R2000 B.n771 B.n770 10.6151
R2001 B.n773 B.n771 10.6151
R2002 B.n774 B.n773 10.6151
R2003 B.n775 B.n774 10.6151
R2004 B.n776 B.n775 10.6151
R2005 B.n778 B.n776 10.6151
R2006 B.n779 B.n778 10.6151
R2007 B.n780 B.n779 10.6151
R2008 B.n781 B.n780 10.6151
R2009 B.n783 B.n781 10.6151
R2010 B.n784 B.n783 10.6151
R2011 B.n785 B.n784 10.6151
R2012 B.n786 B.n785 10.6151
R2013 B.n788 B.n786 10.6151
R2014 B.n789 B.n788 10.6151
R2015 B.n790 B.n789 10.6151
R2016 B.n791 B.n790 10.6151
R2017 B.n793 B.n791 10.6151
R2018 B.n794 B.n793 10.6151
R2019 B.n795 B.n794 10.6151
R2020 B.n796 B.n795 10.6151
R2021 B.n798 B.n796 10.6151
R2022 B.n799 B.n798 10.6151
R2023 B.n800 B.n799 10.6151
R2024 B.n801 B.n800 10.6151
R2025 B.n803 B.n801 10.6151
R2026 B.n804 B.n803 10.6151
R2027 B.n805 B.n804 10.6151
R2028 B.n624 B.n623 10.6151
R2029 B.n623 B.n622 10.6151
R2030 B.n622 B.n621 10.6151
R2031 B.n621 B.n619 10.6151
R2032 B.n619 B.n616 10.6151
R2033 B.n616 B.n615 10.6151
R2034 B.n615 B.n612 10.6151
R2035 B.n612 B.n611 10.6151
R2036 B.n611 B.n608 10.6151
R2037 B.n608 B.n607 10.6151
R2038 B.n607 B.n604 10.6151
R2039 B.n604 B.n603 10.6151
R2040 B.n603 B.n600 10.6151
R2041 B.n600 B.n599 10.6151
R2042 B.n599 B.n596 10.6151
R2043 B.n596 B.n595 10.6151
R2044 B.n595 B.n592 10.6151
R2045 B.n592 B.n591 10.6151
R2046 B.n591 B.n588 10.6151
R2047 B.n588 B.n587 10.6151
R2048 B.n587 B.n584 10.6151
R2049 B.n584 B.n583 10.6151
R2050 B.n583 B.n580 10.6151
R2051 B.n580 B.n579 10.6151
R2052 B.n579 B.n576 10.6151
R2053 B.n576 B.n575 10.6151
R2054 B.n575 B.n572 10.6151
R2055 B.n572 B.n571 10.6151
R2056 B.n571 B.n568 10.6151
R2057 B.n568 B.n567 10.6151
R2058 B.n567 B.n564 10.6151
R2059 B.n564 B.n563 10.6151
R2060 B.n563 B.n560 10.6151
R2061 B.n560 B.n559 10.6151
R2062 B.n559 B.n556 10.6151
R2063 B.n556 B.n555 10.6151
R2064 B.n555 B.n552 10.6151
R2065 B.n552 B.n551 10.6151
R2066 B.n551 B.n548 10.6151
R2067 B.n548 B.n547 10.6151
R2068 B.n547 B.n544 10.6151
R2069 B.n542 B.n539 10.6151
R2070 B.n539 B.n538 10.6151
R2071 B.n538 B.n535 10.6151
R2072 B.n535 B.n534 10.6151
R2073 B.n534 B.n531 10.6151
R2074 B.n531 B.n530 10.6151
R2075 B.n530 B.n527 10.6151
R2076 B.n527 B.n526 10.6151
R2077 B.n523 B.n522 10.6151
R2078 B.n522 B.n519 10.6151
R2079 B.n519 B.n518 10.6151
R2080 B.n518 B.n515 10.6151
R2081 B.n515 B.n514 10.6151
R2082 B.n514 B.n511 10.6151
R2083 B.n511 B.n510 10.6151
R2084 B.n510 B.n507 10.6151
R2085 B.n507 B.n506 10.6151
R2086 B.n506 B.n503 10.6151
R2087 B.n503 B.n502 10.6151
R2088 B.n502 B.n499 10.6151
R2089 B.n499 B.n498 10.6151
R2090 B.n498 B.n495 10.6151
R2091 B.n495 B.n494 10.6151
R2092 B.n494 B.n491 10.6151
R2093 B.n491 B.n490 10.6151
R2094 B.n490 B.n487 10.6151
R2095 B.n487 B.n486 10.6151
R2096 B.n486 B.n483 10.6151
R2097 B.n483 B.n482 10.6151
R2098 B.n482 B.n479 10.6151
R2099 B.n479 B.n478 10.6151
R2100 B.n478 B.n475 10.6151
R2101 B.n475 B.n474 10.6151
R2102 B.n474 B.n471 10.6151
R2103 B.n471 B.n470 10.6151
R2104 B.n470 B.n467 10.6151
R2105 B.n467 B.n466 10.6151
R2106 B.n466 B.n463 10.6151
R2107 B.n463 B.n462 10.6151
R2108 B.n462 B.n459 10.6151
R2109 B.n459 B.n458 10.6151
R2110 B.n458 B.n455 10.6151
R2111 B.n455 B.n454 10.6151
R2112 B.n454 B.n451 10.6151
R2113 B.n451 B.n450 10.6151
R2114 B.n450 B.n447 10.6151
R2115 B.n447 B.n446 10.6151
R2116 B.n446 B.n392 10.6151
R2117 B.n630 B.n392 10.6151
R2118 B.n636 B.n388 10.6151
R2119 B.n637 B.n636 10.6151
R2120 B.n638 B.n637 10.6151
R2121 B.n638 B.n380 10.6151
R2122 B.n648 B.n380 10.6151
R2123 B.n649 B.n648 10.6151
R2124 B.n650 B.n649 10.6151
R2125 B.n650 B.n372 10.6151
R2126 B.n660 B.n372 10.6151
R2127 B.n661 B.n660 10.6151
R2128 B.n662 B.n661 10.6151
R2129 B.n662 B.n364 10.6151
R2130 B.n672 B.n364 10.6151
R2131 B.n673 B.n672 10.6151
R2132 B.n674 B.n673 10.6151
R2133 B.n674 B.n356 10.6151
R2134 B.n685 B.n356 10.6151
R2135 B.n686 B.n685 10.6151
R2136 B.n687 B.n686 10.6151
R2137 B.n687 B.n349 10.6151
R2138 B.n697 B.n349 10.6151
R2139 B.n698 B.n697 10.6151
R2140 B.n699 B.n698 10.6151
R2141 B.n699 B.n341 10.6151
R2142 B.n709 B.n341 10.6151
R2143 B.n710 B.n709 10.6151
R2144 B.n711 B.n710 10.6151
R2145 B.n711 B.n333 10.6151
R2146 B.n721 B.n333 10.6151
R2147 B.n722 B.n721 10.6151
R2148 B.n723 B.n722 10.6151
R2149 B.n723 B.n325 10.6151
R2150 B.n733 B.n325 10.6151
R2151 B.n734 B.n733 10.6151
R2152 B.n735 B.n734 10.6151
R2153 B.n735 B.n317 10.6151
R2154 B.n746 B.n317 10.6151
R2155 B.n747 B.n746 10.6151
R2156 B.n748 B.n747 10.6151
R2157 B.n748 B.n0 10.6151
R2158 B.n886 B.n1 10.6151
R2159 B.n886 B.n885 10.6151
R2160 B.n885 B.n884 10.6151
R2161 B.n884 B.n10 10.6151
R2162 B.n878 B.n10 10.6151
R2163 B.n878 B.n877 10.6151
R2164 B.n877 B.n876 10.6151
R2165 B.n876 B.n17 10.6151
R2166 B.n870 B.n17 10.6151
R2167 B.n870 B.n869 10.6151
R2168 B.n869 B.n868 10.6151
R2169 B.n868 B.n24 10.6151
R2170 B.n862 B.n24 10.6151
R2171 B.n862 B.n861 10.6151
R2172 B.n861 B.n860 10.6151
R2173 B.n860 B.n31 10.6151
R2174 B.n854 B.n31 10.6151
R2175 B.n854 B.n853 10.6151
R2176 B.n853 B.n852 10.6151
R2177 B.n852 B.n38 10.6151
R2178 B.n846 B.n38 10.6151
R2179 B.n846 B.n845 10.6151
R2180 B.n845 B.n844 10.6151
R2181 B.n844 B.n44 10.6151
R2182 B.n838 B.n44 10.6151
R2183 B.n838 B.n837 10.6151
R2184 B.n837 B.n836 10.6151
R2185 B.n836 B.n52 10.6151
R2186 B.n830 B.n52 10.6151
R2187 B.n830 B.n829 10.6151
R2188 B.n829 B.n828 10.6151
R2189 B.n828 B.n59 10.6151
R2190 B.n822 B.n59 10.6151
R2191 B.n822 B.n821 10.6151
R2192 B.n821 B.n820 10.6151
R2193 B.n820 B.n66 10.6151
R2194 B.n814 B.n66 10.6151
R2195 B.n814 B.n813 10.6151
R2196 B.n813 B.n812 10.6151
R2197 B.n812 B.n73 10.6151
R2198 B.n214 B.n128 6.5566
R2199 B.n231 B.n230 6.5566
R2200 B.n543 B.n542 6.5566
R2201 B.n526 B.n444 6.5566
R2202 B.n689 B.t3 5.10935
R2203 B.n848 B.t0 5.10935
R2204 B.n211 B.n128 4.05904
R2205 B.n232 B.n231 4.05904
R2206 B.n544 B.n543 4.05904
R2207 B.n523 B.n444 4.05904
R2208 B.n713 B.t2 3.83214
R2209 B.t5 B.n864 3.83214
R2210 B.n892 B.n0 2.81026
R2211 B.n892 B.n1 2.81026
R2212 VN.n25 VN.n14 161.3
R2213 VN.n24 VN.n23 161.3
R2214 VN.n22 VN.n15 161.3
R2215 VN.n21 VN.n20 161.3
R2216 VN.n19 VN.n16 161.3
R2217 VN.n11 VN.n0 161.3
R2218 VN.n10 VN.n9 161.3
R2219 VN.n8 VN.n1 161.3
R2220 VN.n7 VN.n6 161.3
R2221 VN.n5 VN.n2 161.3
R2222 VN.n3 VN.t5 152.004
R2223 VN.n17 VN.t4 152.004
R2224 VN.n4 VN.t1 117.072
R2225 VN.n12 VN.t3 117.072
R2226 VN.n18 VN.t2 117.072
R2227 VN.n26 VN.t0 117.072
R2228 VN.n13 VN.n12 96.5656
R2229 VN.n27 VN.n26 96.5656
R2230 VN.n6 VN.n1 50.6917
R2231 VN.n20 VN.n15 50.6917
R2232 VN VN.n27 48.4186
R2233 VN.n4 VN.n3 48.0623
R2234 VN.n18 VN.n17 48.0623
R2235 VN.n10 VN.n1 30.2951
R2236 VN.n24 VN.n15 30.2951
R2237 VN.n5 VN.n4 24.4675
R2238 VN.n6 VN.n5 24.4675
R2239 VN.n11 VN.n10 24.4675
R2240 VN.n20 VN.n19 24.4675
R2241 VN.n19 VN.n18 24.4675
R2242 VN.n25 VN.n24 24.4675
R2243 VN.n12 VN.n11 14.1914
R2244 VN.n26 VN.n25 14.1914
R2245 VN.n17 VN.n16 6.56002
R2246 VN.n3 VN.n2 6.56002
R2247 VN.n27 VN.n14 0.278367
R2248 VN.n13 VN.n0 0.278367
R2249 VN.n23 VN.n14 0.189894
R2250 VN.n23 VN.n22 0.189894
R2251 VN.n22 VN.n21 0.189894
R2252 VN.n21 VN.n16 0.189894
R2253 VN.n7 VN.n2 0.189894
R2254 VN.n8 VN.n7 0.189894
R2255 VN.n9 VN.n8 0.189894
R2256 VN.n9 VN.n0 0.189894
R2257 VN VN.n13 0.153454
R2258 VDD2.n131 VDD2.n130 289.615
R2259 VDD2.n64 VDD2.n63 289.615
R2260 VDD2.n130 VDD2.n129 185
R2261 VDD2.n69 VDD2.n68 185
R2262 VDD2.n124 VDD2.n123 185
R2263 VDD2.n122 VDD2.n121 185
R2264 VDD2.n73 VDD2.n72 185
R2265 VDD2.n116 VDD2.n115 185
R2266 VDD2.n114 VDD2.n113 185
R2267 VDD2.n77 VDD2.n76 185
R2268 VDD2.n108 VDD2.n107 185
R2269 VDD2.n106 VDD2.n105 185
R2270 VDD2.n81 VDD2.n80 185
R2271 VDD2.n100 VDD2.n99 185
R2272 VDD2.n98 VDD2.n97 185
R2273 VDD2.n85 VDD2.n84 185
R2274 VDD2.n92 VDD2.n91 185
R2275 VDD2.n90 VDD2.n89 185
R2276 VDD2.n23 VDD2.n22 185
R2277 VDD2.n25 VDD2.n24 185
R2278 VDD2.n18 VDD2.n17 185
R2279 VDD2.n31 VDD2.n30 185
R2280 VDD2.n33 VDD2.n32 185
R2281 VDD2.n14 VDD2.n13 185
R2282 VDD2.n39 VDD2.n38 185
R2283 VDD2.n41 VDD2.n40 185
R2284 VDD2.n10 VDD2.n9 185
R2285 VDD2.n47 VDD2.n46 185
R2286 VDD2.n49 VDD2.n48 185
R2287 VDD2.n6 VDD2.n5 185
R2288 VDD2.n55 VDD2.n54 185
R2289 VDD2.n57 VDD2.n56 185
R2290 VDD2.n2 VDD2.n1 185
R2291 VDD2.n63 VDD2.n62 185
R2292 VDD2.n88 VDD2.t5 147.659
R2293 VDD2.n21 VDD2.t0 147.659
R2294 VDD2.n130 VDD2.n68 104.615
R2295 VDD2.n123 VDD2.n68 104.615
R2296 VDD2.n123 VDD2.n122 104.615
R2297 VDD2.n122 VDD2.n72 104.615
R2298 VDD2.n115 VDD2.n72 104.615
R2299 VDD2.n115 VDD2.n114 104.615
R2300 VDD2.n114 VDD2.n76 104.615
R2301 VDD2.n107 VDD2.n76 104.615
R2302 VDD2.n107 VDD2.n106 104.615
R2303 VDD2.n106 VDD2.n80 104.615
R2304 VDD2.n99 VDD2.n80 104.615
R2305 VDD2.n99 VDD2.n98 104.615
R2306 VDD2.n98 VDD2.n84 104.615
R2307 VDD2.n91 VDD2.n84 104.615
R2308 VDD2.n91 VDD2.n90 104.615
R2309 VDD2.n24 VDD2.n23 104.615
R2310 VDD2.n24 VDD2.n17 104.615
R2311 VDD2.n31 VDD2.n17 104.615
R2312 VDD2.n32 VDD2.n31 104.615
R2313 VDD2.n32 VDD2.n13 104.615
R2314 VDD2.n39 VDD2.n13 104.615
R2315 VDD2.n40 VDD2.n39 104.615
R2316 VDD2.n40 VDD2.n9 104.615
R2317 VDD2.n47 VDD2.n9 104.615
R2318 VDD2.n48 VDD2.n47 104.615
R2319 VDD2.n48 VDD2.n5 104.615
R2320 VDD2.n55 VDD2.n5 104.615
R2321 VDD2.n56 VDD2.n55 104.615
R2322 VDD2.n56 VDD2.n1 104.615
R2323 VDD2.n63 VDD2.n1 104.615
R2324 VDD2.n66 VDD2.n65 65.5152
R2325 VDD2 VDD2.n133 65.5115
R2326 VDD2.n66 VDD2.n64 53.1339
R2327 VDD2.n90 VDD2.t5 52.3082
R2328 VDD2.n23 VDD2.t0 52.3082
R2329 VDD2.n132 VDD2.n131 51.3853
R2330 VDD2.n132 VDD2.n66 41.8338
R2331 VDD2.n89 VDD2.n88 15.6677
R2332 VDD2.n22 VDD2.n21 15.6677
R2333 VDD2.n92 VDD2.n87 12.8005
R2334 VDD2.n25 VDD2.n20 12.8005
R2335 VDD2.n129 VDD2.n67 12.0247
R2336 VDD2.n93 VDD2.n85 12.0247
R2337 VDD2.n26 VDD2.n18 12.0247
R2338 VDD2.n62 VDD2.n0 12.0247
R2339 VDD2.n128 VDD2.n69 11.249
R2340 VDD2.n97 VDD2.n96 11.249
R2341 VDD2.n30 VDD2.n29 11.249
R2342 VDD2.n61 VDD2.n2 11.249
R2343 VDD2.n125 VDD2.n124 10.4732
R2344 VDD2.n100 VDD2.n83 10.4732
R2345 VDD2.n33 VDD2.n16 10.4732
R2346 VDD2.n58 VDD2.n57 10.4732
R2347 VDD2.n121 VDD2.n71 9.69747
R2348 VDD2.n101 VDD2.n81 9.69747
R2349 VDD2.n34 VDD2.n14 9.69747
R2350 VDD2.n54 VDD2.n4 9.69747
R2351 VDD2.n127 VDD2.n67 9.45567
R2352 VDD2.n60 VDD2.n0 9.45567
R2353 VDD2.n75 VDD2.n74 9.3005
R2354 VDD2.n118 VDD2.n117 9.3005
R2355 VDD2.n120 VDD2.n119 9.3005
R2356 VDD2.n71 VDD2.n70 9.3005
R2357 VDD2.n126 VDD2.n125 9.3005
R2358 VDD2.n128 VDD2.n127 9.3005
R2359 VDD2.n112 VDD2.n111 9.3005
R2360 VDD2.n110 VDD2.n109 9.3005
R2361 VDD2.n79 VDD2.n78 9.3005
R2362 VDD2.n104 VDD2.n103 9.3005
R2363 VDD2.n102 VDD2.n101 9.3005
R2364 VDD2.n83 VDD2.n82 9.3005
R2365 VDD2.n96 VDD2.n95 9.3005
R2366 VDD2.n94 VDD2.n93 9.3005
R2367 VDD2.n87 VDD2.n86 9.3005
R2368 VDD2.n45 VDD2.n44 9.3005
R2369 VDD2.n8 VDD2.n7 9.3005
R2370 VDD2.n51 VDD2.n50 9.3005
R2371 VDD2.n53 VDD2.n52 9.3005
R2372 VDD2.n4 VDD2.n3 9.3005
R2373 VDD2.n59 VDD2.n58 9.3005
R2374 VDD2.n61 VDD2.n60 9.3005
R2375 VDD2.n12 VDD2.n11 9.3005
R2376 VDD2.n37 VDD2.n36 9.3005
R2377 VDD2.n35 VDD2.n34 9.3005
R2378 VDD2.n16 VDD2.n15 9.3005
R2379 VDD2.n29 VDD2.n28 9.3005
R2380 VDD2.n27 VDD2.n26 9.3005
R2381 VDD2.n20 VDD2.n19 9.3005
R2382 VDD2.n43 VDD2.n42 9.3005
R2383 VDD2.n120 VDD2.n73 8.92171
R2384 VDD2.n105 VDD2.n104 8.92171
R2385 VDD2.n38 VDD2.n37 8.92171
R2386 VDD2.n53 VDD2.n6 8.92171
R2387 VDD2.n117 VDD2.n116 8.14595
R2388 VDD2.n108 VDD2.n79 8.14595
R2389 VDD2.n41 VDD2.n12 8.14595
R2390 VDD2.n50 VDD2.n49 8.14595
R2391 VDD2.n113 VDD2.n75 7.3702
R2392 VDD2.n109 VDD2.n77 7.3702
R2393 VDD2.n42 VDD2.n10 7.3702
R2394 VDD2.n46 VDD2.n8 7.3702
R2395 VDD2.n113 VDD2.n112 6.59444
R2396 VDD2.n112 VDD2.n77 6.59444
R2397 VDD2.n45 VDD2.n10 6.59444
R2398 VDD2.n46 VDD2.n45 6.59444
R2399 VDD2.n116 VDD2.n75 5.81868
R2400 VDD2.n109 VDD2.n108 5.81868
R2401 VDD2.n42 VDD2.n41 5.81868
R2402 VDD2.n49 VDD2.n8 5.81868
R2403 VDD2.n117 VDD2.n73 5.04292
R2404 VDD2.n105 VDD2.n79 5.04292
R2405 VDD2.n38 VDD2.n12 5.04292
R2406 VDD2.n50 VDD2.n6 5.04292
R2407 VDD2.n88 VDD2.n86 4.38563
R2408 VDD2.n21 VDD2.n19 4.38563
R2409 VDD2.n121 VDD2.n120 4.26717
R2410 VDD2.n104 VDD2.n81 4.26717
R2411 VDD2.n37 VDD2.n14 4.26717
R2412 VDD2.n54 VDD2.n53 4.26717
R2413 VDD2.n124 VDD2.n71 3.49141
R2414 VDD2.n101 VDD2.n100 3.49141
R2415 VDD2.n34 VDD2.n33 3.49141
R2416 VDD2.n57 VDD2.n4 3.49141
R2417 VDD2.n125 VDD2.n69 2.71565
R2418 VDD2.n97 VDD2.n83 2.71565
R2419 VDD2.n30 VDD2.n16 2.71565
R2420 VDD2.n58 VDD2.n2 2.71565
R2421 VDD2.n129 VDD2.n128 1.93989
R2422 VDD2.n96 VDD2.n85 1.93989
R2423 VDD2.n29 VDD2.n18 1.93989
R2424 VDD2.n62 VDD2.n61 1.93989
R2425 VDD2 VDD2.n132 1.86257
R2426 VDD2.n133 VDD2.t3 1.6574
R2427 VDD2.n133 VDD2.t1 1.6574
R2428 VDD2.n65 VDD2.t4 1.6574
R2429 VDD2.n65 VDD2.t2 1.6574
R2430 VDD2.n131 VDD2.n67 1.16414
R2431 VDD2.n93 VDD2.n92 1.16414
R2432 VDD2.n26 VDD2.n25 1.16414
R2433 VDD2.n64 VDD2.n0 1.16414
R2434 VDD2.n89 VDD2.n87 0.388379
R2435 VDD2.n22 VDD2.n20 0.388379
R2436 VDD2.n127 VDD2.n126 0.155672
R2437 VDD2.n126 VDD2.n70 0.155672
R2438 VDD2.n119 VDD2.n70 0.155672
R2439 VDD2.n119 VDD2.n118 0.155672
R2440 VDD2.n118 VDD2.n74 0.155672
R2441 VDD2.n111 VDD2.n74 0.155672
R2442 VDD2.n111 VDD2.n110 0.155672
R2443 VDD2.n110 VDD2.n78 0.155672
R2444 VDD2.n103 VDD2.n78 0.155672
R2445 VDD2.n103 VDD2.n102 0.155672
R2446 VDD2.n102 VDD2.n82 0.155672
R2447 VDD2.n95 VDD2.n82 0.155672
R2448 VDD2.n95 VDD2.n94 0.155672
R2449 VDD2.n94 VDD2.n86 0.155672
R2450 VDD2.n27 VDD2.n19 0.155672
R2451 VDD2.n28 VDD2.n27 0.155672
R2452 VDD2.n28 VDD2.n15 0.155672
R2453 VDD2.n35 VDD2.n15 0.155672
R2454 VDD2.n36 VDD2.n35 0.155672
R2455 VDD2.n36 VDD2.n11 0.155672
R2456 VDD2.n43 VDD2.n11 0.155672
R2457 VDD2.n44 VDD2.n43 0.155672
R2458 VDD2.n44 VDD2.n7 0.155672
R2459 VDD2.n51 VDD2.n7 0.155672
R2460 VDD2.n52 VDD2.n51 0.155672
R2461 VDD2.n52 VDD2.n3 0.155672
R2462 VDD2.n59 VDD2.n3 0.155672
R2463 VDD2.n60 VDD2.n59 0.155672
C0 VDD2 VN 6.62588f
C1 VDD2 VTAIL 7.74169f
C2 VDD2 VDD1 1.35221f
C3 VP VN 6.77958f
C4 VP VTAIL 6.76631f
C5 VN VTAIL 6.75201f
C6 VP VDD1 6.91856f
C7 VN VDD1 0.150512f
C8 VTAIL VDD1 7.69194f
C9 VDD2 VP 0.446417f
C10 VDD2 B 5.862412f
C11 VDD1 B 5.993888f
C12 VTAIL B 7.699682f
C13 VN B 12.47679f
C14 VP B 11.081879f
C15 VDD2.n0 B 0.01201f
C16 VDD2.n1 B 0.027067f
C17 VDD2.n2 B 0.012125f
C18 VDD2.n3 B 0.021311f
C19 VDD2.n4 B 0.011451f
C20 VDD2.n5 B 0.027067f
C21 VDD2.n6 B 0.012125f
C22 VDD2.n7 B 0.021311f
C23 VDD2.n8 B 0.011451f
C24 VDD2.n9 B 0.027067f
C25 VDD2.n10 B 0.012125f
C26 VDD2.n11 B 0.021311f
C27 VDD2.n12 B 0.011451f
C28 VDD2.n13 B 0.027067f
C29 VDD2.n14 B 0.012125f
C30 VDD2.n15 B 0.021311f
C31 VDD2.n16 B 0.011451f
C32 VDD2.n17 B 0.027067f
C33 VDD2.n18 B 0.012125f
C34 VDD2.n19 B 1.08863f
C35 VDD2.n20 B 0.011451f
C36 VDD2.t0 B 0.044408f
C37 VDD2.n21 B 0.122698f
C38 VDD2.n22 B 0.01599f
C39 VDD2.n23 B 0.0203f
C40 VDD2.n24 B 0.027067f
C41 VDD2.n25 B 0.012125f
C42 VDD2.n26 B 0.011451f
C43 VDD2.n27 B 0.021311f
C44 VDD2.n28 B 0.021311f
C45 VDD2.n29 B 0.011451f
C46 VDD2.n30 B 0.012125f
C47 VDD2.n31 B 0.027067f
C48 VDD2.n32 B 0.027067f
C49 VDD2.n33 B 0.012125f
C50 VDD2.n34 B 0.011451f
C51 VDD2.n35 B 0.021311f
C52 VDD2.n36 B 0.021311f
C53 VDD2.n37 B 0.011451f
C54 VDD2.n38 B 0.012125f
C55 VDD2.n39 B 0.027067f
C56 VDD2.n40 B 0.027067f
C57 VDD2.n41 B 0.012125f
C58 VDD2.n42 B 0.011451f
C59 VDD2.n43 B 0.021311f
C60 VDD2.n44 B 0.021311f
C61 VDD2.n45 B 0.011451f
C62 VDD2.n46 B 0.012125f
C63 VDD2.n47 B 0.027067f
C64 VDD2.n48 B 0.027067f
C65 VDD2.n49 B 0.012125f
C66 VDD2.n50 B 0.011451f
C67 VDD2.n51 B 0.021311f
C68 VDD2.n52 B 0.021311f
C69 VDD2.n53 B 0.011451f
C70 VDD2.n54 B 0.012125f
C71 VDD2.n55 B 0.027067f
C72 VDD2.n56 B 0.027067f
C73 VDD2.n57 B 0.012125f
C74 VDD2.n58 B 0.011451f
C75 VDD2.n59 B 0.021311f
C76 VDD2.n60 B 0.054791f
C77 VDD2.n61 B 0.011451f
C78 VDD2.n62 B 0.012125f
C79 VDD2.n63 B 0.054274f
C80 VDD2.n64 B 0.065972f
C81 VDD2.t4 B 0.201244f
C82 VDD2.t2 B 0.201244f
C83 VDD2.n65 B 1.80458f
C84 VDD2.n66 B 2.22341f
C85 VDD2.n67 B 0.01201f
C86 VDD2.n68 B 0.027067f
C87 VDD2.n69 B 0.012125f
C88 VDD2.n70 B 0.021311f
C89 VDD2.n71 B 0.011451f
C90 VDD2.n72 B 0.027067f
C91 VDD2.n73 B 0.012125f
C92 VDD2.n74 B 0.021311f
C93 VDD2.n75 B 0.011451f
C94 VDD2.n76 B 0.027067f
C95 VDD2.n77 B 0.012125f
C96 VDD2.n78 B 0.021311f
C97 VDD2.n79 B 0.011451f
C98 VDD2.n80 B 0.027067f
C99 VDD2.n81 B 0.012125f
C100 VDD2.n82 B 0.021311f
C101 VDD2.n83 B 0.011451f
C102 VDD2.n84 B 0.027067f
C103 VDD2.n85 B 0.012125f
C104 VDD2.n86 B 1.08863f
C105 VDD2.n87 B 0.011451f
C106 VDD2.t5 B 0.044408f
C107 VDD2.n88 B 0.122698f
C108 VDD2.n89 B 0.01599f
C109 VDD2.n90 B 0.0203f
C110 VDD2.n91 B 0.027067f
C111 VDD2.n92 B 0.012125f
C112 VDD2.n93 B 0.011451f
C113 VDD2.n94 B 0.021311f
C114 VDD2.n95 B 0.021311f
C115 VDD2.n96 B 0.011451f
C116 VDD2.n97 B 0.012125f
C117 VDD2.n98 B 0.027067f
C118 VDD2.n99 B 0.027067f
C119 VDD2.n100 B 0.012125f
C120 VDD2.n101 B 0.011451f
C121 VDD2.n102 B 0.021311f
C122 VDD2.n103 B 0.021311f
C123 VDD2.n104 B 0.011451f
C124 VDD2.n105 B 0.012125f
C125 VDD2.n106 B 0.027067f
C126 VDD2.n107 B 0.027067f
C127 VDD2.n108 B 0.012125f
C128 VDD2.n109 B 0.011451f
C129 VDD2.n110 B 0.021311f
C130 VDD2.n111 B 0.021311f
C131 VDD2.n112 B 0.011451f
C132 VDD2.n113 B 0.012125f
C133 VDD2.n114 B 0.027067f
C134 VDD2.n115 B 0.027067f
C135 VDD2.n116 B 0.012125f
C136 VDD2.n117 B 0.011451f
C137 VDD2.n118 B 0.021311f
C138 VDD2.n119 B 0.021311f
C139 VDD2.n120 B 0.011451f
C140 VDD2.n121 B 0.012125f
C141 VDD2.n122 B 0.027067f
C142 VDD2.n123 B 0.027067f
C143 VDD2.n124 B 0.012125f
C144 VDD2.n125 B 0.011451f
C145 VDD2.n126 B 0.021311f
C146 VDD2.n127 B 0.054791f
C147 VDD2.n128 B 0.011451f
C148 VDD2.n129 B 0.012125f
C149 VDD2.n130 B 0.054274f
C150 VDD2.n131 B 0.060589f
C151 VDD2.n132 B 2.14972f
C152 VDD2.t3 B 0.201244f
C153 VDD2.t1 B 0.201244f
C154 VDD2.n133 B 1.80456f
C155 VN.n0 B 0.031904f
C156 VN.t3 B 1.938f
C157 VN.n1 B 0.023222f
C158 VN.n2 B 0.230359f
C159 VN.t1 B 1.938f
C160 VN.t5 B 2.12976f
C161 VN.n3 B 0.730643f
C162 VN.n4 B 0.767465f
C163 VN.n5 B 0.045101f
C164 VN.n6 B 0.044179f
C165 VN.n7 B 0.024199f
C166 VN.n8 B 0.024199f
C167 VN.n9 B 0.024199f
C168 VN.n10 B 0.048356f
C169 VN.n11 B 0.035749f
C170 VN.n12 B 0.769216f
C171 VN.n13 B 0.035623f
C172 VN.n14 B 0.031904f
C173 VN.t0 B 1.938f
C174 VN.n15 B 0.023222f
C175 VN.n16 B 0.230359f
C176 VN.t2 B 1.938f
C177 VN.t4 B 2.12976f
C178 VN.n17 B 0.730643f
C179 VN.n18 B 0.767465f
C180 VN.n19 B 0.045101f
C181 VN.n20 B 0.044179f
C182 VN.n21 B 0.024199f
C183 VN.n22 B 0.024199f
C184 VN.n23 B 0.024199f
C185 VN.n24 B 0.048356f
C186 VN.n25 B 0.035749f
C187 VN.n26 B 0.769216f
C188 VN.n27 B 1.28249f
C189 VDD1.n0 B 0.012195f
C190 VDD1.n1 B 0.027484f
C191 VDD1.n2 B 0.012312f
C192 VDD1.n3 B 0.021639f
C193 VDD1.n4 B 0.011628f
C194 VDD1.n5 B 0.027484f
C195 VDD1.n6 B 0.012312f
C196 VDD1.n7 B 0.021639f
C197 VDD1.n8 B 0.011628f
C198 VDD1.n9 B 0.027484f
C199 VDD1.n10 B 0.012312f
C200 VDD1.n11 B 0.021639f
C201 VDD1.n12 B 0.011628f
C202 VDD1.n13 B 0.027484f
C203 VDD1.n14 B 0.012312f
C204 VDD1.n15 B 0.021639f
C205 VDD1.n16 B 0.011628f
C206 VDD1.n17 B 0.027484f
C207 VDD1.n18 B 0.012312f
C208 VDD1.n19 B 1.10538f
C209 VDD1.n20 B 0.011628f
C210 VDD1.t1 B 0.045091f
C211 VDD1.n21 B 0.124586f
C212 VDD1.n22 B 0.016236f
C213 VDD1.n23 B 0.020613f
C214 VDD1.n24 B 0.027484f
C215 VDD1.n25 B 0.012312f
C216 VDD1.n26 B 0.011628f
C217 VDD1.n27 B 0.021639f
C218 VDD1.n28 B 0.021639f
C219 VDD1.n29 B 0.011628f
C220 VDD1.n30 B 0.012312f
C221 VDD1.n31 B 0.027484f
C222 VDD1.n32 B 0.027484f
C223 VDD1.n33 B 0.012312f
C224 VDD1.n34 B 0.011628f
C225 VDD1.n35 B 0.021639f
C226 VDD1.n36 B 0.021639f
C227 VDD1.n37 B 0.011628f
C228 VDD1.n38 B 0.012312f
C229 VDD1.n39 B 0.027484f
C230 VDD1.n40 B 0.027484f
C231 VDD1.n41 B 0.012312f
C232 VDD1.n42 B 0.011628f
C233 VDD1.n43 B 0.021639f
C234 VDD1.n44 B 0.021639f
C235 VDD1.n45 B 0.011628f
C236 VDD1.n46 B 0.012312f
C237 VDD1.n47 B 0.027484f
C238 VDD1.n48 B 0.027484f
C239 VDD1.n49 B 0.012312f
C240 VDD1.n50 B 0.011628f
C241 VDD1.n51 B 0.021639f
C242 VDD1.n52 B 0.021639f
C243 VDD1.n53 B 0.011628f
C244 VDD1.n54 B 0.012312f
C245 VDD1.n55 B 0.027484f
C246 VDD1.n56 B 0.027484f
C247 VDD1.n57 B 0.012312f
C248 VDD1.n58 B 0.011628f
C249 VDD1.n59 B 0.021639f
C250 VDD1.n60 B 0.055634f
C251 VDD1.n61 B 0.011628f
C252 VDD1.n62 B 0.012312f
C253 VDD1.n63 B 0.055109f
C254 VDD1.n64 B 0.067596f
C255 VDD1.n65 B 0.012195f
C256 VDD1.n66 B 0.027484f
C257 VDD1.n67 B 0.012312f
C258 VDD1.n68 B 0.021639f
C259 VDD1.n69 B 0.011628f
C260 VDD1.n70 B 0.027484f
C261 VDD1.n71 B 0.012312f
C262 VDD1.n72 B 0.021639f
C263 VDD1.n73 B 0.011628f
C264 VDD1.n74 B 0.027484f
C265 VDD1.n75 B 0.012312f
C266 VDD1.n76 B 0.021639f
C267 VDD1.n77 B 0.011628f
C268 VDD1.n78 B 0.027484f
C269 VDD1.n79 B 0.012312f
C270 VDD1.n80 B 0.021639f
C271 VDD1.n81 B 0.011628f
C272 VDD1.n82 B 0.027484f
C273 VDD1.n83 B 0.012312f
C274 VDD1.n84 B 1.10538f
C275 VDD1.n85 B 0.011628f
C276 VDD1.t0 B 0.045091f
C277 VDD1.n86 B 0.124586f
C278 VDD1.n87 B 0.016236f
C279 VDD1.n88 B 0.020613f
C280 VDD1.n89 B 0.027484f
C281 VDD1.n90 B 0.012312f
C282 VDD1.n91 B 0.011628f
C283 VDD1.n92 B 0.021639f
C284 VDD1.n93 B 0.021639f
C285 VDD1.n94 B 0.011628f
C286 VDD1.n95 B 0.012312f
C287 VDD1.n96 B 0.027484f
C288 VDD1.n97 B 0.027484f
C289 VDD1.n98 B 0.012312f
C290 VDD1.n99 B 0.011628f
C291 VDD1.n100 B 0.021639f
C292 VDD1.n101 B 0.021639f
C293 VDD1.n102 B 0.011628f
C294 VDD1.n103 B 0.012312f
C295 VDD1.n104 B 0.027484f
C296 VDD1.n105 B 0.027484f
C297 VDD1.n106 B 0.012312f
C298 VDD1.n107 B 0.011628f
C299 VDD1.n108 B 0.021639f
C300 VDD1.n109 B 0.021639f
C301 VDD1.n110 B 0.011628f
C302 VDD1.n111 B 0.012312f
C303 VDD1.n112 B 0.027484f
C304 VDD1.n113 B 0.027484f
C305 VDD1.n114 B 0.012312f
C306 VDD1.n115 B 0.011628f
C307 VDD1.n116 B 0.021639f
C308 VDD1.n117 B 0.021639f
C309 VDD1.n118 B 0.011628f
C310 VDD1.n119 B 0.012312f
C311 VDD1.n120 B 0.027484f
C312 VDD1.n121 B 0.027484f
C313 VDD1.n122 B 0.012312f
C314 VDD1.n123 B 0.011628f
C315 VDD1.n124 B 0.021639f
C316 VDD1.n125 B 0.055634f
C317 VDD1.n126 B 0.011628f
C318 VDD1.n127 B 0.012312f
C319 VDD1.n128 B 0.055109f
C320 VDD1.n129 B 0.066987f
C321 VDD1.t2 B 0.204341f
C322 VDD1.t3 B 0.204341f
C323 VDD1.n130 B 1.83235f
C324 VDD1.n131 B 2.36188f
C325 VDD1.t4 B 0.204341f
C326 VDD1.t5 B 0.204341f
C327 VDD1.n132 B 1.82914f
C328 VDD1.n133 B 2.36932f
C329 VTAIL.t1 B 0.223729f
C330 VTAIL.t5 B 0.223729f
C331 VTAIL.n0 B 1.93986f
C332 VTAIL.n1 B 0.395054f
C333 VTAIL.n2 B 0.013352f
C334 VTAIL.n3 B 0.030091f
C335 VTAIL.n4 B 0.01348f
C336 VTAIL.n5 B 0.023692f
C337 VTAIL.n6 B 0.012731f
C338 VTAIL.n7 B 0.030091f
C339 VTAIL.n8 B 0.01348f
C340 VTAIL.n9 B 0.023692f
C341 VTAIL.n10 B 0.012731f
C342 VTAIL.n11 B 0.030091f
C343 VTAIL.n12 B 0.01348f
C344 VTAIL.n13 B 0.023692f
C345 VTAIL.n14 B 0.012731f
C346 VTAIL.n15 B 0.030091f
C347 VTAIL.n16 B 0.01348f
C348 VTAIL.n17 B 0.023692f
C349 VTAIL.n18 B 0.012731f
C350 VTAIL.n19 B 0.030091f
C351 VTAIL.n20 B 0.01348f
C352 VTAIL.n21 B 1.21026f
C353 VTAIL.n22 B 0.012731f
C354 VTAIL.t11 B 0.049369f
C355 VTAIL.n23 B 0.136407f
C356 VTAIL.n24 B 0.017776f
C357 VTAIL.n25 B 0.022569f
C358 VTAIL.n26 B 0.030091f
C359 VTAIL.n27 B 0.01348f
C360 VTAIL.n28 B 0.012731f
C361 VTAIL.n29 B 0.023692f
C362 VTAIL.n30 B 0.023692f
C363 VTAIL.n31 B 0.012731f
C364 VTAIL.n32 B 0.01348f
C365 VTAIL.n33 B 0.030091f
C366 VTAIL.n34 B 0.030091f
C367 VTAIL.n35 B 0.01348f
C368 VTAIL.n36 B 0.012731f
C369 VTAIL.n37 B 0.023692f
C370 VTAIL.n38 B 0.023692f
C371 VTAIL.n39 B 0.012731f
C372 VTAIL.n40 B 0.01348f
C373 VTAIL.n41 B 0.030091f
C374 VTAIL.n42 B 0.030091f
C375 VTAIL.n43 B 0.01348f
C376 VTAIL.n44 B 0.012731f
C377 VTAIL.n45 B 0.023692f
C378 VTAIL.n46 B 0.023692f
C379 VTAIL.n47 B 0.012731f
C380 VTAIL.n48 B 0.01348f
C381 VTAIL.n49 B 0.030091f
C382 VTAIL.n50 B 0.030091f
C383 VTAIL.n51 B 0.01348f
C384 VTAIL.n52 B 0.012731f
C385 VTAIL.n53 B 0.023692f
C386 VTAIL.n54 B 0.023692f
C387 VTAIL.n55 B 0.012731f
C388 VTAIL.n56 B 0.01348f
C389 VTAIL.n57 B 0.030091f
C390 VTAIL.n58 B 0.030091f
C391 VTAIL.n59 B 0.01348f
C392 VTAIL.n60 B 0.012731f
C393 VTAIL.n61 B 0.023692f
C394 VTAIL.n62 B 0.060912f
C395 VTAIL.n63 B 0.012731f
C396 VTAIL.n64 B 0.01348f
C397 VTAIL.n65 B 0.060337f
C398 VTAIL.n66 B 0.051031f
C399 VTAIL.n67 B 0.333899f
C400 VTAIL.t6 B 0.223729f
C401 VTAIL.t10 B 0.223729f
C402 VTAIL.n68 B 1.93986f
C403 VTAIL.n69 B 1.87614f
C404 VTAIL.t3 B 0.223729f
C405 VTAIL.t2 B 0.223729f
C406 VTAIL.n70 B 1.93987f
C407 VTAIL.n71 B 1.87613f
C408 VTAIL.n72 B 0.013352f
C409 VTAIL.n73 B 0.030091f
C410 VTAIL.n74 B 0.01348f
C411 VTAIL.n75 B 0.023692f
C412 VTAIL.n76 B 0.012731f
C413 VTAIL.n77 B 0.030091f
C414 VTAIL.n78 B 0.01348f
C415 VTAIL.n79 B 0.023692f
C416 VTAIL.n80 B 0.012731f
C417 VTAIL.n81 B 0.030091f
C418 VTAIL.n82 B 0.01348f
C419 VTAIL.n83 B 0.023692f
C420 VTAIL.n84 B 0.012731f
C421 VTAIL.n85 B 0.030091f
C422 VTAIL.n86 B 0.01348f
C423 VTAIL.n87 B 0.023692f
C424 VTAIL.n88 B 0.012731f
C425 VTAIL.n89 B 0.030091f
C426 VTAIL.n90 B 0.01348f
C427 VTAIL.n91 B 1.21026f
C428 VTAIL.n92 B 0.012731f
C429 VTAIL.t4 B 0.049369f
C430 VTAIL.n93 B 0.136407f
C431 VTAIL.n94 B 0.017776f
C432 VTAIL.n95 B 0.022569f
C433 VTAIL.n96 B 0.030091f
C434 VTAIL.n97 B 0.01348f
C435 VTAIL.n98 B 0.012731f
C436 VTAIL.n99 B 0.023692f
C437 VTAIL.n100 B 0.023692f
C438 VTAIL.n101 B 0.012731f
C439 VTAIL.n102 B 0.01348f
C440 VTAIL.n103 B 0.030091f
C441 VTAIL.n104 B 0.030091f
C442 VTAIL.n105 B 0.01348f
C443 VTAIL.n106 B 0.012731f
C444 VTAIL.n107 B 0.023692f
C445 VTAIL.n108 B 0.023692f
C446 VTAIL.n109 B 0.012731f
C447 VTAIL.n110 B 0.01348f
C448 VTAIL.n111 B 0.030091f
C449 VTAIL.n112 B 0.030091f
C450 VTAIL.n113 B 0.01348f
C451 VTAIL.n114 B 0.012731f
C452 VTAIL.n115 B 0.023692f
C453 VTAIL.n116 B 0.023692f
C454 VTAIL.n117 B 0.012731f
C455 VTAIL.n118 B 0.01348f
C456 VTAIL.n119 B 0.030091f
C457 VTAIL.n120 B 0.030091f
C458 VTAIL.n121 B 0.01348f
C459 VTAIL.n122 B 0.012731f
C460 VTAIL.n123 B 0.023692f
C461 VTAIL.n124 B 0.023692f
C462 VTAIL.n125 B 0.012731f
C463 VTAIL.n126 B 0.01348f
C464 VTAIL.n127 B 0.030091f
C465 VTAIL.n128 B 0.030091f
C466 VTAIL.n129 B 0.01348f
C467 VTAIL.n130 B 0.012731f
C468 VTAIL.n131 B 0.023692f
C469 VTAIL.n132 B 0.060912f
C470 VTAIL.n133 B 0.012731f
C471 VTAIL.n134 B 0.01348f
C472 VTAIL.n135 B 0.060337f
C473 VTAIL.n136 B 0.051031f
C474 VTAIL.n137 B 0.333899f
C475 VTAIL.t7 B 0.223729f
C476 VTAIL.t8 B 0.223729f
C477 VTAIL.n138 B 1.93987f
C478 VTAIL.n139 B 0.528315f
C479 VTAIL.n140 B 0.013352f
C480 VTAIL.n141 B 0.030091f
C481 VTAIL.n142 B 0.01348f
C482 VTAIL.n143 B 0.023692f
C483 VTAIL.n144 B 0.012731f
C484 VTAIL.n145 B 0.030091f
C485 VTAIL.n146 B 0.01348f
C486 VTAIL.n147 B 0.023692f
C487 VTAIL.n148 B 0.012731f
C488 VTAIL.n149 B 0.030091f
C489 VTAIL.n150 B 0.01348f
C490 VTAIL.n151 B 0.023692f
C491 VTAIL.n152 B 0.012731f
C492 VTAIL.n153 B 0.030091f
C493 VTAIL.n154 B 0.01348f
C494 VTAIL.n155 B 0.023692f
C495 VTAIL.n156 B 0.012731f
C496 VTAIL.n157 B 0.030091f
C497 VTAIL.n158 B 0.01348f
C498 VTAIL.n159 B 1.21026f
C499 VTAIL.n160 B 0.012731f
C500 VTAIL.t9 B 0.049369f
C501 VTAIL.n161 B 0.136407f
C502 VTAIL.n162 B 0.017776f
C503 VTAIL.n163 B 0.022569f
C504 VTAIL.n164 B 0.030091f
C505 VTAIL.n165 B 0.01348f
C506 VTAIL.n166 B 0.012731f
C507 VTAIL.n167 B 0.023692f
C508 VTAIL.n168 B 0.023692f
C509 VTAIL.n169 B 0.012731f
C510 VTAIL.n170 B 0.01348f
C511 VTAIL.n171 B 0.030091f
C512 VTAIL.n172 B 0.030091f
C513 VTAIL.n173 B 0.01348f
C514 VTAIL.n174 B 0.012731f
C515 VTAIL.n175 B 0.023692f
C516 VTAIL.n176 B 0.023692f
C517 VTAIL.n177 B 0.012731f
C518 VTAIL.n178 B 0.01348f
C519 VTAIL.n179 B 0.030091f
C520 VTAIL.n180 B 0.030091f
C521 VTAIL.n181 B 0.01348f
C522 VTAIL.n182 B 0.012731f
C523 VTAIL.n183 B 0.023692f
C524 VTAIL.n184 B 0.023692f
C525 VTAIL.n185 B 0.012731f
C526 VTAIL.n186 B 0.01348f
C527 VTAIL.n187 B 0.030091f
C528 VTAIL.n188 B 0.030091f
C529 VTAIL.n189 B 0.01348f
C530 VTAIL.n190 B 0.012731f
C531 VTAIL.n191 B 0.023692f
C532 VTAIL.n192 B 0.023692f
C533 VTAIL.n193 B 0.012731f
C534 VTAIL.n194 B 0.01348f
C535 VTAIL.n195 B 0.030091f
C536 VTAIL.n196 B 0.030091f
C537 VTAIL.n197 B 0.01348f
C538 VTAIL.n198 B 0.012731f
C539 VTAIL.n199 B 0.023692f
C540 VTAIL.n200 B 0.060912f
C541 VTAIL.n201 B 0.012731f
C542 VTAIL.n202 B 0.01348f
C543 VTAIL.n203 B 0.060337f
C544 VTAIL.n204 B 0.051031f
C545 VTAIL.n205 B 1.4981f
C546 VTAIL.n206 B 0.013352f
C547 VTAIL.n207 B 0.030091f
C548 VTAIL.n208 B 0.01348f
C549 VTAIL.n209 B 0.023692f
C550 VTAIL.n210 B 0.012731f
C551 VTAIL.n211 B 0.030091f
C552 VTAIL.n212 B 0.01348f
C553 VTAIL.n213 B 0.023692f
C554 VTAIL.n214 B 0.012731f
C555 VTAIL.n215 B 0.030091f
C556 VTAIL.n216 B 0.01348f
C557 VTAIL.n217 B 0.023692f
C558 VTAIL.n218 B 0.012731f
C559 VTAIL.n219 B 0.030091f
C560 VTAIL.n220 B 0.01348f
C561 VTAIL.n221 B 0.023692f
C562 VTAIL.n222 B 0.012731f
C563 VTAIL.n223 B 0.030091f
C564 VTAIL.n224 B 0.01348f
C565 VTAIL.n225 B 1.21026f
C566 VTAIL.n226 B 0.012731f
C567 VTAIL.t0 B 0.049369f
C568 VTAIL.n227 B 0.136407f
C569 VTAIL.n228 B 0.017776f
C570 VTAIL.n229 B 0.022569f
C571 VTAIL.n230 B 0.030091f
C572 VTAIL.n231 B 0.01348f
C573 VTAIL.n232 B 0.012731f
C574 VTAIL.n233 B 0.023692f
C575 VTAIL.n234 B 0.023692f
C576 VTAIL.n235 B 0.012731f
C577 VTAIL.n236 B 0.01348f
C578 VTAIL.n237 B 0.030091f
C579 VTAIL.n238 B 0.030091f
C580 VTAIL.n239 B 0.01348f
C581 VTAIL.n240 B 0.012731f
C582 VTAIL.n241 B 0.023692f
C583 VTAIL.n242 B 0.023692f
C584 VTAIL.n243 B 0.012731f
C585 VTAIL.n244 B 0.01348f
C586 VTAIL.n245 B 0.030091f
C587 VTAIL.n246 B 0.030091f
C588 VTAIL.n247 B 0.01348f
C589 VTAIL.n248 B 0.012731f
C590 VTAIL.n249 B 0.023692f
C591 VTAIL.n250 B 0.023692f
C592 VTAIL.n251 B 0.012731f
C593 VTAIL.n252 B 0.01348f
C594 VTAIL.n253 B 0.030091f
C595 VTAIL.n254 B 0.030091f
C596 VTAIL.n255 B 0.01348f
C597 VTAIL.n256 B 0.012731f
C598 VTAIL.n257 B 0.023692f
C599 VTAIL.n258 B 0.023692f
C600 VTAIL.n259 B 0.012731f
C601 VTAIL.n260 B 0.01348f
C602 VTAIL.n261 B 0.030091f
C603 VTAIL.n262 B 0.030091f
C604 VTAIL.n263 B 0.01348f
C605 VTAIL.n264 B 0.012731f
C606 VTAIL.n265 B 0.023692f
C607 VTAIL.n266 B 0.060912f
C608 VTAIL.n267 B 0.012731f
C609 VTAIL.n268 B 0.01348f
C610 VTAIL.n269 B 0.060337f
C611 VTAIL.n270 B 0.051031f
C612 VTAIL.n271 B 1.44776f
C613 VP.n0 B 0.032432f
C614 VP.t2 B 1.9701f
C615 VP.n1 B 0.023607f
C616 VP.n2 B 0.0246f
C617 VP.t3 B 1.9701f
C618 VP.n3 B 0.045848f
C619 VP.n4 B 0.0246f
C620 VP.n5 B 0.036341f
C621 VP.n6 B 0.032432f
C622 VP.t0 B 1.9701f
C623 VP.n7 B 0.023607f
C624 VP.n8 B 0.234175f
C625 VP.t1 B 1.9701f
C626 VP.t4 B 2.16504f
C627 VP.n9 B 0.742745f
C628 VP.n10 B 0.780177f
C629 VP.n11 B 0.045848f
C630 VP.n12 B 0.044911f
C631 VP.n13 B 0.0246f
C632 VP.n14 B 0.0246f
C633 VP.n15 B 0.0246f
C634 VP.n16 B 0.049157f
C635 VP.n17 B 0.036341f
C636 VP.n18 B 0.781957f
C637 VP.n19 B 1.29043f
C638 VP.t5 B 1.9701f
C639 VP.n20 B 0.781957f
C640 VP.n21 B 1.3088f
C641 VP.n22 B 0.032432f
C642 VP.n23 B 0.0246f
C643 VP.n24 B 0.049157f
C644 VP.n25 B 0.023607f
C645 VP.n26 B 0.044911f
C646 VP.n27 B 0.0246f
C647 VP.n28 B 0.0246f
C648 VP.n29 B 0.0246f
C649 VP.n30 B 0.721391f
C650 VP.n31 B 0.045848f
C651 VP.n32 B 0.044911f
C652 VP.n33 B 0.0246f
C653 VP.n34 B 0.0246f
C654 VP.n35 B 0.0246f
C655 VP.n36 B 0.049157f
C656 VP.n37 B 0.036341f
C657 VP.n38 B 0.781957f
C658 VP.n39 B 0.036213f
.ends

