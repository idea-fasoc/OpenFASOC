* NGSPICE file created from diff_pair_sample_0864.ext - technology: sky130A

.subckt diff_pair_sample_0864 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.06095 pd=6.76 as=2.5077 ps=13.64 w=6.43 l=1.07
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=0 ps=0 w=6.43 l=1.07
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=0 ps=0 w=6.43 l=1.07
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.06095 pd=6.76 as=2.5077 ps=13.64 w=6.43 l=1.07
X4 VTAIL.t4 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=1.06095 ps=6.76 w=6.43 l=1.07
X5 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=1.06095 ps=6.76 w=6.43 l=1.07
X6 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=1.06095 ps=6.76 w=6.43 l=1.07
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=0 ps=0 w=6.43 l=1.07
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=0 ps=0 w=6.43 l=1.07
X9 VDD2.t1 VN.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.06095 pd=6.76 as=2.5077 ps=13.64 w=6.43 l=1.07
X10 VTAIL.t6 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5077 pd=13.64 as=1.06095 ps=6.76 w=6.43 l=1.07
X11 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.06095 pd=6.76 as=2.5077 ps=13.64 w=6.43 l=1.07
R0 VN.n0 VN.t3 200.37
R1 VN.n1 VN.t2 200.37
R2 VN.n1 VN.t1 200.284
R3 VN.n0 VN.t0 200.284
R4 VN VN.n1 68.9933
R5 VN VN.n0 31.2622
R6 VTAIL.n5 VTAIL.t1 54.3541
R7 VTAIL.n4 VTAIL.t7 54.3541
R8 VTAIL.n3 VTAIL.t4 54.3541
R9 VTAIL.n6 VTAIL.t3 54.354
R10 VTAIL.n7 VTAIL.t5 54.354
R11 VTAIL.n0 VTAIL.t6 54.354
R12 VTAIL.n1 VTAIL.t2 54.354
R13 VTAIL.n2 VTAIL.t0 54.354
R14 VTAIL.n7 VTAIL.n6 19.1169
R15 VTAIL.n3 VTAIL.n2 19.1169
R16 VTAIL.n4 VTAIL.n3 1.2074
R17 VTAIL.n6 VTAIL.n5 1.2074
R18 VTAIL.n2 VTAIL.n1 1.2074
R19 VTAIL VTAIL.n0 0.662138
R20 VTAIL VTAIL.n7 0.545759
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 100.832
R24 VDD2.n2 VDD2.n1 67.9535
R25 VDD2.n1 VDD2.t2 3.07982
R26 VDD2.n1 VDD2.t1 3.07982
R27 VDD2.n0 VDD2.t0 3.07982
R28 VDD2.n0 VDD2.t3 3.07982
R29 VDD2 VDD2.n2 0.0586897
R30 B.n475 B.n474 585
R31 B.n191 B.n70 585
R32 B.n190 B.n189 585
R33 B.n188 B.n187 585
R34 B.n186 B.n185 585
R35 B.n184 B.n183 585
R36 B.n182 B.n181 585
R37 B.n180 B.n179 585
R38 B.n178 B.n177 585
R39 B.n176 B.n175 585
R40 B.n174 B.n173 585
R41 B.n172 B.n171 585
R42 B.n170 B.n169 585
R43 B.n168 B.n167 585
R44 B.n166 B.n165 585
R45 B.n164 B.n163 585
R46 B.n162 B.n161 585
R47 B.n160 B.n159 585
R48 B.n158 B.n157 585
R49 B.n156 B.n155 585
R50 B.n154 B.n153 585
R51 B.n152 B.n151 585
R52 B.n150 B.n149 585
R53 B.n148 B.n147 585
R54 B.n146 B.n145 585
R55 B.n143 B.n142 585
R56 B.n141 B.n140 585
R57 B.n139 B.n138 585
R58 B.n137 B.n136 585
R59 B.n135 B.n134 585
R60 B.n133 B.n132 585
R61 B.n131 B.n130 585
R62 B.n129 B.n128 585
R63 B.n127 B.n126 585
R64 B.n125 B.n124 585
R65 B.n122 B.n121 585
R66 B.n120 B.n119 585
R67 B.n118 B.n117 585
R68 B.n116 B.n115 585
R69 B.n114 B.n113 585
R70 B.n112 B.n111 585
R71 B.n110 B.n109 585
R72 B.n108 B.n107 585
R73 B.n106 B.n105 585
R74 B.n104 B.n103 585
R75 B.n102 B.n101 585
R76 B.n100 B.n99 585
R77 B.n98 B.n97 585
R78 B.n96 B.n95 585
R79 B.n94 B.n93 585
R80 B.n92 B.n91 585
R81 B.n90 B.n89 585
R82 B.n88 B.n87 585
R83 B.n86 B.n85 585
R84 B.n84 B.n83 585
R85 B.n82 B.n81 585
R86 B.n80 B.n79 585
R87 B.n78 B.n77 585
R88 B.n76 B.n75 585
R89 B.n39 B.n38 585
R90 B.n473 B.n40 585
R91 B.n478 B.n40 585
R92 B.n472 B.n471 585
R93 B.n471 B.n36 585
R94 B.n470 B.n35 585
R95 B.n484 B.n35 585
R96 B.n469 B.n34 585
R97 B.n485 B.n34 585
R98 B.n468 B.n33 585
R99 B.n486 B.n33 585
R100 B.n467 B.n466 585
R101 B.n466 B.n32 585
R102 B.n465 B.n28 585
R103 B.n492 B.n28 585
R104 B.n464 B.n27 585
R105 B.n493 B.n27 585
R106 B.n463 B.n26 585
R107 B.n494 B.n26 585
R108 B.n462 B.n461 585
R109 B.n461 B.n22 585
R110 B.n460 B.n21 585
R111 B.n500 B.n21 585
R112 B.n459 B.n20 585
R113 B.n501 B.n20 585
R114 B.n458 B.n19 585
R115 B.n502 B.n19 585
R116 B.n457 B.n456 585
R117 B.n456 B.n15 585
R118 B.n455 B.n14 585
R119 B.n508 B.n14 585
R120 B.n454 B.n13 585
R121 B.n509 B.n13 585
R122 B.n453 B.n12 585
R123 B.n510 B.n12 585
R124 B.n452 B.n451 585
R125 B.n451 B.n450 585
R126 B.n449 B.n448 585
R127 B.n449 B.n8 585
R128 B.n447 B.n7 585
R129 B.n517 B.n7 585
R130 B.n446 B.n6 585
R131 B.n518 B.n6 585
R132 B.n445 B.n5 585
R133 B.n519 B.n5 585
R134 B.n444 B.n443 585
R135 B.n443 B.n4 585
R136 B.n442 B.n192 585
R137 B.n442 B.n441 585
R138 B.n432 B.n193 585
R139 B.n194 B.n193 585
R140 B.n434 B.n433 585
R141 B.n435 B.n434 585
R142 B.n431 B.n199 585
R143 B.n199 B.n198 585
R144 B.n430 B.n429 585
R145 B.n429 B.n428 585
R146 B.n201 B.n200 585
R147 B.n202 B.n201 585
R148 B.n421 B.n420 585
R149 B.n422 B.n421 585
R150 B.n419 B.n207 585
R151 B.n207 B.n206 585
R152 B.n418 B.n417 585
R153 B.n417 B.n416 585
R154 B.n209 B.n208 585
R155 B.n210 B.n209 585
R156 B.n409 B.n408 585
R157 B.n410 B.n409 585
R158 B.n407 B.n215 585
R159 B.n215 B.n214 585
R160 B.n406 B.n405 585
R161 B.n405 B.n404 585
R162 B.n217 B.n216 585
R163 B.n397 B.n217 585
R164 B.n396 B.n395 585
R165 B.n398 B.n396 585
R166 B.n394 B.n222 585
R167 B.n222 B.n221 585
R168 B.n393 B.n392 585
R169 B.n392 B.n391 585
R170 B.n224 B.n223 585
R171 B.n225 B.n224 585
R172 B.n384 B.n383 585
R173 B.n385 B.n384 585
R174 B.n228 B.n227 585
R175 B.n267 B.n266 585
R176 B.n268 B.n264 585
R177 B.n264 B.n229 585
R178 B.n270 B.n269 585
R179 B.n272 B.n263 585
R180 B.n275 B.n274 585
R181 B.n276 B.n262 585
R182 B.n278 B.n277 585
R183 B.n280 B.n261 585
R184 B.n283 B.n282 585
R185 B.n284 B.n260 585
R186 B.n286 B.n285 585
R187 B.n288 B.n259 585
R188 B.n291 B.n290 585
R189 B.n292 B.n258 585
R190 B.n294 B.n293 585
R191 B.n296 B.n257 585
R192 B.n299 B.n298 585
R193 B.n300 B.n256 585
R194 B.n302 B.n301 585
R195 B.n304 B.n255 585
R196 B.n307 B.n306 585
R197 B.n308 B.n254 585
R198 B.n310 B.n309 585
R199 B.n312 B.n253 585
R200 B.n315 B.n314 585
R201 B.n316 B.n249 585
R202 B.n318 B.n317 585
R203 B.n320 B.n248 585
R204 B.n323 B.n322 585
R205 B.n324 B.n247 585
R206 B.n326 B.n325 585
R207 B.n328 B.n246 585
R208 B.n331 B.n330 585
R209 B.n332 B.n243 585
R210 B.n335 B.n334 585
R211 B.n337 B.n242 585
R212 B.n340 B.n339 585
R213 B.n341 B.n241 585
R214 B.n343 B.n342 585
R215 B.n345 B.n240 585
R216 B.n348 B.n347 585
R217 B.n349 B.n239 585
R218 B.n351 B.n350 585
R219 B.n353 B.n238 585
R220 B.n356 B.n355 585
R221 B.n357 B.n237 585
R222 B.n359 B.n358 585
R223 B.n361 B.n236 585
R224 B.n364 B.n363 585
R225 B.n365 B.n235 585
R226 B.n367 B.n366 585
R227 B.n369 B.n234 585
R228 B.n372 B.n371 585
R229 B.n373 B.n233 585
R230 B.n375 B.n374 585
R231 B.n377 B.n232 585
R232 B.n378 B.n231 585
R233 B.n381 B.n380 585
R234 B.n382 B.n230 585
R235 B.n230 B.n229 585
R236 B.n387 B.n386 585
R237 B.n386 B.n385 585
R238 B.n388 B.n226 585
R239 B.n226 B.n225 585
R240 B.n390 B.n389 585
R241 B.n391 B.n390 585
R242 B.n220 B.n219 585
R243 B.n221 B.n220 585
R244 B.n400 B.n399 585
R245 B.n399 B.n398 585
R246 B.n401 B.n218 585
R247 B.n397 B.n218 585
R248 B.n403 B.n402 585
R249 B.n404 B.n403 585
R250 B.n213 B.n212 585
R251 B.n214 B.n213 585
R252 B.n412 B.n411 585
R253 B.n411 B.n410 585
R254 B.n413 B.n211 585
R255 B.n211 B.n210 585
R256 B.n415 B.n414 585
R257 B.n416 B.n415 585
R258 B.n205 B.n204 585
R259 B.n206 B.n205 585
R260 B.n424 B.n423 585
R261 B.n423 B.n422 585
R262 B.n425 B.n203 585
R263 B.n203 B.n202 585
R264 B.n427 B.n426 585
R265 B.n428 B.n427 585
R266 B.n197 B.n196 585
R267 B.n198 B.n197 585
R268 B.n437 B.n436 585
R269 B.n436 B.n435 585
R270 B.n438 B.n195 585
R271 B.n195 B.n194 585
R272 B.n440 B.n439 585
R273 B.n441 B.n440 585
R274 B.n3 B.n0 585
R275 B.n4 B.n3 585
R276 B.n516 B.n1 585
R277 B.n517 B.n516 585
R278 B.n515 B.n514 585
R279 B.n515 B.n8 585
R280 B.n513 B.n9 585
R281 B.n450 B.n9 585
R282 B.n512 B.n511 585
R283 B.n511 B.n510 585
R284 B.n11 B.n10 585
R285 B.n509 B.n11 585
R286 B.n507 B.n506 585
R287 B.n508 B.n507 585
R288 B.n505 B.n16 585
R289 B.n16 B.n15 585
R290 B.n504 B.n503 585
R291 B.n503 B.n502 585
R292 B.n18 B.n17 585
R293 B.n501 B.n18 585
R294 B.n499 B.n498 585
R295 B.n500 B.n499 585
R296 B.n497 B.n23 585
R297 B.n23 B.n22 585
R298 B.n496 B.n495 585
R299 B.n495 B.n494 585
R300 B.n25 B.n24 585
R301 B.n493 B.n25 585
R302 B.n491 B.n490 585
R303 B.n492 B.n491 585
R304 B.n489 B.n29 585
R305 B.n32 B.n29 585
R306 B.n488 B.n487 585
R307 B.n487 B.n486 585
R308 B.n31 B.n30 585
R309 B.n485 B.n31 585
R310 B.n483 B.n482 585
R311 B.n484 B.n483 585
R312 B.n481 B.n37 585
R313 B.n37 B.n36 585
R314 B.n480 B.n479 585
R315 B.n479 B.n478 585
R316 B.n520 B.n519 585
R317 B.n518 B.n2 585
R318 B.n479 B.n39 497.305
R319 B.n475 B.n40 497.305
R320 B.n384 B.n230 497.305
R321 B.n386 B.n228 497.305
R322 B.n73 B.t15 348.204
R323 B.n71 B.t11 348.204
R324 B.n244 B.t4 348.204
R325 B.n250 B.t8 348.204
R326 B.n477 B.n476 256.663
R327 B.n477 B.n69 256.663
R328 B.n477 B.n68 256.663
R329 B.n477 B.n67 256.663
R330 B.n477 B.n66 256.663
R331 B.n477 B.n65 256.663
R332 B.n477 B.n64 256.663
R333 B.n477 B.n63 256.663
R334 B.n477 B.n62 256.663
R335 B.n477 B.n61 256.663
R336 B.n477 B.n60 256.663
R337 B.n477 B.n59 256.663
R338 B.n477 B.n58 256.663
R339 B.n477 B.n57 256.663
R340 B.n477 B.n56 256.663
R341 B.n477 B.n55 256.663
R342 B.n477 B.n54 256.663
R343 B.n477 B.n53 256.663
R344 B.n477 B.n52 256.663
R345 B.n477 B.n51 256.663
R346 B.n477 B.n50 256.663
R347 B.n477 B.n49 256.663
R348 B.n477 B.n48 256.663
R349 B.n477 B.n47 256.663
R350 B.n477 B.n46 256.663
R351 B.n477 B.n45 256.663
R352 B.n477 B.n44 256.663
R353 B.n477 B.n43 256.663
R354 B.n477 B.n42 256.663
R355 B.n477 B.n41 256.663
R356 B.n265 B.n229 256.663
R357 B.n271 B.n229 256.663
R358 B.n273 B.n229 256.663
R359 B.n279 B.n229 256.663
R360 B.n281 B.n229 256.663
R361 B.n287 B.n229 256.663
R362 B.n289 B.n229 256.663
R363 B.n295 B.n229 256.663
R364 B.n297 B.n229 256.663
R365 B.n303 B.n229 256.663
R366 B.n305 B.n229 256.663
R367 B.n311 B.n229 256.663
R368 B.n313 B.n229 256.663
R369 B.n319 B.n229 256.663
R370 B.n321 B.n229 256.663
R371 B.n327 B.n229 256.663
R372 B.n329 B.n229 256.663
R373 B.n336 B.n229 256.663
R374 B.n338 B.n229 256.663
R375 B.n344 B.n229 256.663
R376 B.n346 B.n229 256.663
R377 B.n352 B.n229 256.663
R378 B.n354 B.n229 256.663
R379 B.n360 B.n229 256.663
R380 B.n362 B.n229 256.663
R381 B.n368 B.n229 256.663
R382 B.n370 B.n229 256.663
R383 B.n376 B.n229 256.663
R384 B.n379 B.n229 256.663
R385 B.n522 B.n521 256.663
R386 B.n77 B.n76 163.367
R387 B.n81 B.n80 163.367
R388 B.n85 B.n84 163.367
R389 B.n89 B.n88 163.367
R390 B.n93 B.n92 163.367
R391 B.n97 B.n96 163.367
R392 B.n101 B.n100 163.367
R393 B.n105 B.n104 163.367
R394 B.n109 B.n108 163.367
R395 B.n113 B.n112 163.367
R396 B.n117 B.n116 163.367
R397 B.n121 B.n120 163.367
R398 B.n126 B.n125 163.367
R399 B.n130 B.n129 163.367
R400 B.n134 B.n133 163.367
R401 B.n138 B.n137 163.367
R402 B.n142 B.n141 163.367
R403 B.n147 B.n146 163.367
R404 B.n151 B.n150 163.367
R405 B.n155 B.n154 163.367
R406 B.n159 B.n158 163.367
R407 B.n163 B.n162 163.367
R408 B.n167 B.n166 163.367
R409 B.n171 B.n170 163.367
R410 B.n175 B.n174 163.367
R411 B.n179 B.n178 163.367
R412 B.n183 B.n182 163.367
R413 B.n187 B.n186 163.367
R414 B.n189 B.n70 163.367
R415 B.n384 B.n224 163.367
R416 B.n392 B.n224 163.367
R417 B.n392 B.n222 163.367
R418 B.n396 B.n222 163.367
R419 B.n396 B.n217 163.367
R420 B.n405 B.n217 163.367
R421 B.n405 B.n215 163.367
R422 B.n409 B.n215 163.367
R423 B.n409 B.n209 163.367
R424 B.n417 B.n209 163.367
R425 B.n417 B.n207 163.367
R426 B.n421 B.n207 163.367
R427 B.n421 B.n201 163.367
R428 B.n429 B.n201 163.367
R429 B.n429 B.n199 163.367
R430 B.n434 B.n199 163.367
R431 B.n434 B.n193 163.367
R432 B.n442 B.n193 163.367
R433 B.n443 B.n442 163.367
R434 B.n443 B.n5 163.367
R435 B.n6 B.n5 163.367
R436 B.n7 B.n6 163.367
R437 B.n449 B.n7 163.367
R438 B.n451 B.n449 163.367
R439 B.n451 B.n12 163.367
R440 B.n13 B.n12 163.367
R441 B.n14 B.n13 163.367
R442 B.n456 B.n14 163.367
R443 B.n456 B.n19 163.367
R444 B.n20 B.n19 163.367
R445 B.n21 B.n20 163.367
R446 B.n461 B.n21 163.367
R447 B.n461 B.n26 163.367
R448 B.n27 B.n26 163.367
R449 B.n28 B.n27 163.367
R450 B.n466 B.n28 163.367
R451 B.n466 B.n33 163.367
R452 B.n34 B.n33 163.367
R453 B.n35 B.n34 163.367
R454 B.n471 B.n35 163.367
R455 B.n471 B.n40 163.367
R456 B.n266 B.n264 163.367
R457 B.n270 B.n264 163.367
R458 B.n274 B.n272 163.367
R459 B.n278 B.n262 163.367
R460 B.n282 B.n280 163.367
R461 B.n286 B.n260 163.367
R462 B.n290 B.n288 163.367
R463 B.n294 B.n258 163.367
R464 B.n298 B.n296 163.367
R465 B.n302 B.n256 163.367
R466 B.n306 B.n304 163.367
R467 B.n310 B.n254 163.367
R468 B.n314 B.n312 163.367
R469 B.n318 B.n249 163.367
R470 B.n322 B.n320 163.367
R471 B.n326 B.n247 163.367
R472 B.n330 B.n328 163.367
R473 B.n335 B.n243 163.367
R474 B.n339 B.n337 163.367
R475 B.n343 B.n241 163.367
R476 B.n347 B.n345 163.367
R477 B.n351 B.n239 163.367
R478 B.n355 B.n353 163.367
R479 B.n359 B.n237 163.367
R480 B.n363 B.n361 163.367
R481 B.n367 B.n235 163.367
R482 B.n371 B.n369 163.367
R483 B.n375 B.n233 163.367
R484 B.n378 B.n377 163.367
R485 B.n380 B.n230 163.367
R486 B.n386 B.n226 163.367
R487 B.n390 B.n226 163.367
R488 B.n390 B.n220 163.367
R489 B.n399 B.n220 163.367
R490 B.n399 B.n218 163.367
R491 B.n403 B.n218 163.367
R492 B.n403 B.n213 163.367
R493 B.n411 B.n213 163.367
R494 B.n411 B.n211 163.367
R495 B.n415 B.n211 163.367
R496 B.n415 B.n205 163.367
R497 B.n423 B.n205 163.367
R498 B.n423 B.n203 163.367
R499 B.n427 B.n203 163.367
R500 B.n427 B.n197 163.367
R501 B.n436 B.n197 163.367
R502 B.n436 B.n195 163.367
R503 B.n440 B.n195 163.367
R504 B.n440 B.n3 163.367
R505 B.n520 B.n3 163.367
R506 B.n516 B.n2 163.367
R507 B.n516 B.n515 163.367
R508 B.n515 B.n9 163.367
R509 B.n511 B.n9 163.367
R510 B.n511 B.n11 163.367
R511 B.n507 B.n11 163.367
R512 B.n507 B.n16 163.367
R513 B.n503 B.n16 163.367
R514 B.n503 B.n18 163.367
R515 B.n499 B.n18 163.367
R516 B.n499 B.n23 163.367
R517 B.n495 B.n23 163.367
R518 B.n495 B.n25 163.367
R519 B.n491 B.n25 163.367
R520 B.n491 B.n29 163.367
R521 B.n487 B.n29 163.367
R522 B.n487 B.n31 163.367
R523 B.n483 B.n31 163.367
R524 B.n483 B.n37 163.367
R525 B.n479 B.n37 163.367
R526 B.n385 B.n229 113.713
R527 B.n478 B.n477 113.713
R528 B.n71 B.t13 102.386
R529 B.n244 B.t7 102.386
R530 B.n73 B.t16 102.379
R531 B.n250 B.t10 102.379
R532 B.n72 B.t14 75.2346
R533 B.n245 B.t6 75.2346
R534 B.n74 B.t17 75.2278
R535 B.n251 B.t9 75.2278
R536 B.n41 B.n39 71.676
R537 B.n77 B.n42 71.676
R538 B.n81 B.n43 71.676
R539 B.n85 B.n44 71.676
R540 B.n89 B.n45 71.676
R541 B.n93 B.n46 71.676
R542 B.n97 B.n47 71.676
R543 B.n101 B.n48 71.676
R544 B.n105 B.n49 71.676
R545 B.n109 B.n50 71.676
R546 B.n113 B.n51 71.676
R547 B.n117 B.n52 71.676
R548 B.n121 B.n53 71.676
R549 B.n126 B.n54 71.676
R550 B.n130 B.n55 71.676
R551 B.n134 B.n56 71.676
R552 B.n138 B.n57 71.676
R553 B.n142 B.n58 71.676
R554 B.n147 B.n59 71.676
R555 B.n151 B.n60 71.676
R556 B.n155 B.n61 71.676
R557 B.n159 B.n62 71.676
R558 B.n163 B.n63 71.676
R559 B.n167 B.n64 71.676
R560 B.n171 B.n65 71.676
R561 B.n175 B.n66 71.676
R562 B.n179 B.n67 71.676
R563 B.n183 B.n68 71.676
R564 B.n187 B.n69 71.676
R565 B.n476 B.n70 71.676
R566 B.n476 B.n475 71.676
R567 B.n189 B.n69 71.676
R568 B.n186 B.n68 71.676
R569 B.n182 B.n67 71.676
R570 B.n178 B.n66 71.676
R571 B.n174 B.n65 71.676
R572 B.n170 B.n64 71.676
R573 B.n166 B.n63 71.676
R574 B.n162 B.n62 71.676
R575 B.n158 B.n61 71.676
R576 B.n154 B.n60 71.676
R577 B.n150 B.n59 71.676
R578 B.n146 B.n58 71.676
R579 B.n141 B.n57 71.676
R580 B.n137 B.n56 71.676
R581 B.n133 B.n55 71.676
R582 B.n129 B.n54 71.676
R583 B.n125 B.n53 71.676
R584 B.n120 B.n52 71.676
R585 B.n116 B.n51 71.676
R586 B.n112 B.n50 71.676
R587 B.n108 B.n49 71.676
R588 B.n104 B.n48 71.676
R589 B.n100 B.n47 71.676
R590 B.n96 B.n46 71.676
R591 B.n92 B.n45 71.676
R592 B.n88 B.n44 71.676
R593 B.n84 B.n43 71.676
R594 B.n80 B.n42 71.676
R595 B.n76 B.n41 71.676
R596 B.n265 B.n228 71.676
R597 B.n271 B.n270 71.676
R598 B.n274 B.n273 71.676
R599 B.n279 B.n278 71.676
R600 B.n282 B.n281 71.676
R601 B.n287 B.n286 71.676
R602 B.n290 B.n289 71.676
R603 B.n295 B.n294 71.676
R604 B.n298 B.n297 71.676
R605 B.n303 B.n302 71.676
R606 B.n306 B.n305 71.676
R607 B.n311 B.n310 71.676
R608 B.n314 B.n313 71.676
R609 B.n319 B.n318 71.676
R610 B.n322 B.n321 71.676
R611 B.n327 B.n326 71.676
R612 B.n330 B.n329 71.676
R613 B.n336 B.n335 71.676
R614 B.n339 B.n338 71.676
R615 B.n344 B.n343 71.676
R616 B.n347 B.n346 71.676
R617 B.n352 B.n351 71.676
R618 B.n355 B.n354 71.676
R619 B.n360 B.n359 71.676
R620 B.n363 B.n362 71.676
R621 B.n368 B.n367 71.676
R622 B.n371 B.n370 71.676
R623 B.n376 B.n375 71.676
R624 B.n379 B.n378 71.676
R625 B.n266 B.n265 71.676
R626 B.n272 B.n271 71.676
R627 B.n273 B.n262 71.676
R628 B.n280 B.n279 71.676
R629 B.n281 B.n260 71.676
R630 B.n288 B.n287 71.676
R631 B.n289 B.n258 71.676
R632 B.n296 B.n295 71.676
R633 B.n297 B.n256 71.676
R634 B.n304 B.n303 71.676
R635 B.n305 B.n254 71.676
R636 B.n312 B.n311 71.676
R637 B.n313 B.n249 71.676
R638 B.n320 B.n319 71.676
R639 B.n321 B.n247 71.676
R640 B.n328 B.n327 71.676
R641 B.n329 B.n243 71.676
R642 B.n337 B.n336 71.676
R643 B.n338 B.n241 71.676
R644 B.n345 B.n344 71.676
R645 B.n346 B.n239 71.676
R646 B.n353 B.n352 71.676
R647 B.n354 B.n237 71.676
R648 B.n361 B.n360 71.676
R649 B.n362 B.n235 71.676
R650 B.n369 B.n368 71.676
R651 B.n370 B.n233 71.676
R652 B.n377 B.n376 71.676
R653 B.n380 B.n379 71.676
R654 B.n521 B.n520 71.676
R655 B.n521 B.n2 71.676
R656 B.n385 B.n225 63.9048
R657 B.n391 B.n225 63.9048
R658 B.n391 B.n221 63.9048
R659 B.n398 B.n221 63.9048
R660 B.n398 B.n397 63.9048
R661 B.n404 B.n214 63.9048
R662 B.n410 B.n214 63.9048
R663 B.n410 B.n210 63.9048
R664 B.n416 B.n210 63.9048
R665 B.n416 B.n206 63.9048
R666 B.n422 B.n206 63.9048
R667 B.n428 B.n202 63.9048
R668 B.n428 B.n198 63.9048
R669 B.n435 B.n198 63.9048
R670 B.n441 B.n194 63.9048
R671 B.n441 B.n4 63.9048
R672 B.n519 B.n4 63.9048
R673 B.n519 B.n518 63.9048
R674 B.n518 B.n517 63.9048
R675 B.n517 B.n8 63.9048
R676 B.n450 B.n8 63.9048
R677 B.n510 B.n509 63.9048
R678 B.n509 B.n508 63.9048
R679 B.n508 B.n15 63.9048
R680 B.n502 B.n501 63.9048
R681 B.n501 B.n500 63.9048
R682 B.n500 B.n22 63.9048
R683 B.n494 B.n22 63.9048
R684 B.n494 B.n493 63.9048
R685 B.n493 B.n492 63.9048
R686 B.n486 B.n32 63.9048
R687 B.n486 B.n485 63.9048
R688 B.n485 B.n484 63.9048
R689 B.n484 B.n36 63.9048
R690 B.n478 B.n36 63.9048
R691 B.n123 B.n74 59.5399
R692 B.n144 B.n72 59.5399
R693 B.n333 B.n245 59.5399
R694 B.n252 B.n251 59.5399
R695 B.n435 B.t2 53.5674
R696 B.n510 B.t1 53.5674
R697 B.n422 B.t0 46.0492
R698 B.n502 B.t3 46.0492
R699 B.n404 B.t5 38.531
R700 B.n492 B.t12 38.531
R701 B.n387 B.n227 32.3127
R702 B.n383 B.n382 32.3127
R703 B.n474 B.n473 32.3127
R704 B.n480 B.n38 32.3127
R705 B.n74 B.n73 27.152
R706 B.n72 B.n71 27.152
R707 B.n245 B.n244 27.152
R708 B.n251 B.n250 27.152
R709 B.n397 B.t5 25.3743
R710 B.n32 B.t12 25.3743
R711 B B.n522 18.0485
R712 B.t0 B.n202 17.8561
R713 B.t3 B.n15 17.8561
R714 B.n388 B.n387 10.6151
R715 B.n389 B.n388 10.6151
R716 B.n389 B.n219 10.6151
R717 B.n400 B.n219 10.6151
R718 B.n401 B.n400 10.6151
R719 B.n402 B.n401 10.6151
R720 B.n402 B.n212 10.6151
R721 B.n412 B.n212 10.6151
R722 B.n413 B.n412 10.6151
R723 B.n414 B.n413 10.6151
R724 B.n414 B.n204 10.6151
R725 B.n424 B.n204 10.6151
R726 B.n425 B.n424 10.6151
R727 B.n426 B.n425 10.6151
R728 B.n426 B.n196 10.6151
R729 B.n437 B.n196 10.6151
R730 B.n438 B.n437 10.6151
R731 B.n439 B.n438 10.6151
R732 B.n439 B.n0 10.6151
R733 B.n267 B.n227 10.6151
R734 B.n268 B.n267 10.6151
R735 B.n269 B.n268 10.6151
R736 B.n269 B.n263 10.6151
R737 B.n275 B.n263 10.6151
R738 B.n276 B.n275 10.6151
R739 B.n277 B.n276 10.6151
R740 B.n277 B.n261 10.6151
R741 B.n283 B.n261 10.6151
R742 B.n284 B.n283 10.6151
R743 B.n285 B.n284 10.6151
R744 B.n285 B.n259 10.6151
R745 B.n291 B.n259 10.6151
R746 B.n292 B.n291 10.6151
R747 B.n293 B.n292 10.6151
R748 B.n293 B.n257 10.6151
R749 B.n299 B.n257 10.6151
R750 B.n300 B.n299 10.6151
R751 B.n301 B.n300 10.6151
R752 B.n301 B.n255 10.6151
R753 B.n307 B.n255 10.6151
R754 B.n308 B.n307 10.6151
R755 B.n309 B.n308 10.6151
R756 B.n309 B.n253 10.6151
R757 B.n316 B.n315 10.6151
R758 B.n317 B.n316 10.6151
R759 B.n317 B.n248 10.6151
R760 B.n323 B.n248 10.6151
R761 B.n324 B.n323 10.6151
R762 B.n325 B.n324 10.6151
R763 B.n325 B.n246 10.6151
R764 B.n331 B.n246 10.6151
R765 B.n332 B.n331 10.6151
R766 B.n334 B.n242 10.6151
R767 B.n340 B.n242 10.6151
R768 B.n341 B.n340 10.6151
R769 B.n342 B.n341 10.6151
R770 B.n342 B.n240 10.6151
R771 B.n348 B.n240 10.6151
R772 B.n349 B.n348 10.6151
R773 B.n350 B.n349 10.6151
R774 B.n350 B.n238 10.6151
R775 B.n356 B.n238 10.6151
R776 B.n357 B.n356 10.6151
R777 B.n358 B.n357 10.6151
R778 B.n358 B.n236 10.6151
R779 B.n364 B.n236 10.6151
R780 B.n365 B.n364 10.6151
R781 B.n366 B.n365 10.6151
R782 B.n366 B.n234 10.6151
R783 B.n372 B.n234 10.6151
R784 B.n373 B.n372 10.6151
R785 B.n374 B.n373 10.6151
R786 B.n374 B.n232 10.6151
R787 B.n232 B.n231 10.6151
R788 B.n381 B.n231 10.6151
R789 B.n382 B.n381 10.6151
R790 B.n383 B.n223 10.6151
R791 B.n393 B.n223 10.6151
R792 B.n394 B.n393 10.6151
R793 B.n395 B.n394 10.6151
R794 B.n395 B.n216 10.6151
R795 B.n406 B.n216 10.6151
R796 B.n407 B.n406 10.6151
R797 B.n408 B.n407 10.6151
R798 B.n408 B.n208 10.6151
R799 B.n418 B.n208 10.6151
R800 B.n419 B.n418 10.6151
R801 B.n420 B.n419 10.6151
R802 B.n420 B.n200 10.6151
R803 B.n430 B.n200 10.6151
R804 B.n431 B.n430 10.6151
R805 B.n433 B.n431 10.6151
R806 B.n433 B.n432 10.6151
R807 B.n432 B.n192 10.6151
R808 B.n444 B.n192 10.6151
R809 B.n445 B.n444 10.6151
R810 B.n446 B.n445 10.6151
R811 B.n447 B.n446 10.6151
R812 B.n448 B.n447 10.6151
R813 B.n452 B.n448 10.6151
R814 B.n453 B.n452 10.6151
R815 B.n454 B.n453 10.6151
R816 B.n455 B.n454 10.6151
R817 B.n457 B.n455 10.6151
R818 B.n458 B.n457 10.6151
R819 B.n459 B.n458 10.6151
R820 B.n460 B.n459 10.6151
R821 B.n462 B.n460 10.6151
R822 B.n463 B.n462 10.6151
R823 B.n464 B.n463 10.6151
R824 B.n465 B.n464 10.6151
R825 B.n467 B.n465 10.6151
R826 B.n468 B.n467 10.6151
R827 B.n469 B.n468 10.6151
R828 B.n470 B.n469 10.6151
R829 B.n472 B.n470 10.6151
R830 B.n473 B.n472 10.6151
R831 B.n514 B.n1 10.6151
R832 B.n514 B.n513 10.6151
R833 B.n513 B.n512 10.6151
R834 B.n512 B.n10 10.6151
R835 B.n506 B.n10 10.6151
R836 B.n506 B.n505 10.6151
R837 B.n505 B.n504 10.6151
R838 B.n504 B.n17 10.6151
R839 B.n498 B.n17 10.6151
R840 B.n498 B.n497 10.6151
R841 B.n497 B.n496 10.6151
R842 B.n496 B.n24 10.6151
R843 B.n490 B.n24 10.6151
R844 B.n490 B.n489 10.6151
R845 B.n489 B.n488 10.6151
R846 B.n488 B.n30 10.6151
R847 B.n482 B.n30 10.6151
R848 B.n482 B.n481 10.6151
R849 B.n481 B.n480 10.6151
R850 B.n75 B.n38 10.6151
R851 B.n78 B.n75 10.6151
R852 B.n79 B.n78 10.6151
R853 B.n82 B.n79 10.6151
R854 B.n83 B.n82 10.6151
R855 B.n86 B.n83 10.6151
R856 B.n87 B.n86 10.6151
R857 B.n90 B.n87 10.6151
R858 B.n91 B.n90 10.6151
R859 B.n94 B.n91 10.6151
R860 B.n95 B.n94 10.6151
R861 B.n98 B.n95 10.6151
R862 B.n99 B.n98 10.6151
R863 B.n102 B.n99 10.6151
R864 B.n103 B.n102 10.6151
R865 B.n106 B.n103 10.6151
R866 B.n107 B.n106 10.6151
R867 B.n110 B.n107 10.6151
R868 B.n111 B.n110 10.6151
R869 B.n114 B.n111 10.6151
R870 B.n115 B.n114 10.6151
R871 B.n118 B.n115 10.6151
R872 B.n119 B.n118 10.6151
R873 B.n122 B.n119 10.6151
R874 B.n127 B.n124 10.6151
R875 B.n128 B.n127 10.6151
R876 B.n131 B.n128 10.6151
R877 B.n132 B.n131 10.6151
R878 B.n135 B.n132 10.6151
R879 B.n136 B.n135 10.6151
R880 B.n139 B.n136 10.6151
R881 B.n140 B.n139 10.6151
R882 B.n143 B.n140 10.6151
R883 B.n148 B.n145 10.6151
R884 B.n149 B.n148 10.6151
R885 B.n152 B.n149 10.6151
R886 B.n153 B.n152 10.6151
R887 B.n156 B.n153 10.6151
R888 B.n157 B.n156 10.6151
R889 B.n160 B.n157 10.6151
R890 B.n161 B.n160 10.6151
R891 B.n164 B.n161 10.6151
R892 B.n165 B.n164 10.6151
R893 B.n168 B.n165 10.6151
R894 B.n169 B.n168 10.6151
R895 B.n172 B.n169 10.6151
R896 B.n173 B.n172 10.6151
R897 B.n176 B.n173 10.6151
R898 B.n177 B.n176 10.6151
R899 B.n180 B.n177 10.6151
R900 B.n181 B.n180 10.6151
R901 B.n184 B.n181 10.6151
R902 B.n185 B.n184 10.6151
R903 B.n188 B.n185 10.6151
R904 B.n190 B.n188 10.6151
R905 B.n191 B.n190 10.6151
R906 B.n474 B.n191 10.6151
R907 B.t2 B.n194 10.338
R908 B.n450 B.t1 10.338
R909 B.n253 B.n252 9.36635
R910 B.n334 B.n333 9.36635
R911 B.n123 B.n122 9.36635
R912 B.n145 B.n144 9.36635
R913 B.n522 B.n0 8.11757
R914 B.n522 B.n1 8.11757
R915 B.n315 B.n252 1.24928
R916 B.n333 B.n332 1.24928
R917 B.n124 B.n123 1.24928
R918 B.n144 B.n143 1.24928
R919 VP.n0 VP.t2 200.37
R920 VP.n0 VP.t3 200.284
R921 VP.n2 VP.t1 181.764
R922 VP.n3 VP.t0 181.764
R923 VP.n4 VP.n3 80.6037
R924 VP.n2 VP.n1 80.6037
R925 VP.n1 VP.n0 68.7077
R926 VP.n3 VP.n2 48.2005
R927 VP.n4 VP.n1 0.380177
R928 VP VP.n4 0.146778
R929 VDD1 VDD1.n1 101.356
R930 VDD1 VDD1.n0 68.0116
R931 VDD1.n0 VDD1.t1 3.07982
R932 VDD1.n0 VDD1.t0 3.07982
R933 VDD1.n1 VDD1.t2 3.07982
R934 VDD1.n1 VDD1.t3 3.07982
C0 VN VDD2 2.14606f
C1 VP VDD2 0.297061f
C2 VDD1 VDD2 0.65527f
C3 VN VP 4.05538f
C4 VDD1 VN 0.147729f
C5 VDD1 VP 2.29504f
C6 VTAIL VDD2 4.00339f
C7 VTAIL VN 2.10941f
C8 VTAIL VP 2.12352f
C9 VDD1 VTAIL 3.95944f
C10 VDD2 B 2.47203f
C11 VDD1 B 5.53995f
C12 VTAIL B 5.732608f
C13 VN B 7.72089f
C14 VP B 5.246064f
C15 VDD1.t1 B 0.138801f
C16 VDD1.t0 B 0.138801f
C17 VDD1.n0 B 1.16797f
C18 VDD1.t2 B 0.138801f
C19 VDD1.t3 B 0.138801f
C20 VDD1.n1 B 1.59198f
C21 VP.t3 B 0.925359f
C22 VP.t2 B 0.925562f
C23 VP.n0 B 1.6301f
C24 VP.n1 B 2.3396f
C25 VP.t1 B 0.888345f
C26 VP.n2 B 0.40029f
C27 VP.t0 B 0.888345f
C28 VP.n3 B 0.40029f
C29 VP.n4 B 0.056674f
C30 VDD2.t0 B 0.136582f
C31 VDD2.t3 B 0.136582f
C32 VDD2.n0 B 1.54419f
C33 VDD2.t2 B 0.136582f
C34 VDD2.t1 B 0.136582f
C35 VDD2.n1 B 1.14901f
C36 VDD2.n2 B 2.75015f
C37 VTAIL.t6 B 0.911807f
C38 VTAIL.n0 B 0.281038f
C39 VTAIL.t2 B 0.911807f
C40 VTAIL.n1 B 0.3123f
C41 VTAIL.t0 B 0.911807f
C42 VTAIL.n2 B 0.914085f
C43 VTAIL.t4 B 0.911813f
C44 VTAIL.n3 B 0.91408f
C45 VTAIL.t7 B 0.911813f
C46 VTAIL.n4 B 0.312295f
C47 VTAIL.t1 B 0.911813f
C48 VTAIL.n5 B 0.312295f
C49 VTAIL.t3 B 0.911807f
C50 VTAIL.n6 B 0.914085f
C51 VTAIL.t5 B 0.911807f
C52 VTAIL.n7 B 0.87615f
C53 VN.t3 B 0.897167f
C54 VN.t0 B 0.896971f
C55 VN.n0 B 0.705249f
C56 VN.t2 B 0.897167f
C57 VN.t1 B 0.896971f
C58 VN.n1 B 1.59668f
.ends

