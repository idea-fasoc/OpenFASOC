* NGSPICE file created from diff_pair_sample_0611.ext - technology: sky130A

.subckt diff_pair_sample_0611 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X1 VTAIL.t7 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=2.80005 ps=17.3 w=16.97 l=1.15
X2 VTAIL.t14 VN.t1 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=2.80005 ps=17.3 w=16.97 l=1.15
X3 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=0 ps=0 w=16.97 l=1.15
X4 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=0 ps=0 w=16.97 l=1.15
X5 VTAIL.t13 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X6 VDD1.t6 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=6.6183 ps=34.72 w=16.97 l=1.15
X7 VDD2.t2 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X8 VDD2.t5 VN.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=6.6183 ps=34.72 w=16.97 l=1.15
X9 VDD2.t4 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X10 VDD1.t5 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X11 VDD2.t7 VN.t6 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=6.6183 ps=34.72 w=16.97 l=1.15
X12 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=2.80005 ps=17.3 w=16.97 l=1.15
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=0 ps=0 w=16.97 l=1.15
X14 VDD1.t3 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=6.6183 ps=34.72 w=16.97 l=1.15
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=0 ps=0 w=16.97 l=1.15
X16 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X17 VTAIL.t8 VN.t7 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6183 pd=34.72 as=2.80005 ps=17.3 w=16.97 l=1.15
X18 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
X19 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.80005 pd=17.3 as=2.80005 ps=17.3 w=16.97 l=1.15
R0 VN.n3 VN.t1 413.253
R1 VN.n16 VN.t6 413.253
R2 VN.n11 VN.t4 390.002
R3 VN.n24 VN.t7 390.002
R4 VN.n4 VN.t3 355.632
R5 VN.n1 VN.t2 355.632
R6 VN.n17 VN.t0 355.632
R7 VN.n14 VN.t5 355.632
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN.n11 VN.n10 51.3812
R21 VN.n24 VN.n23 51.3812
R22 VN VN.n25 48.393
R23 VN.n4 VN.n3 33.3566
R24 VN.n17 VN.n16 33.3566
R25 VN.n16 VN.n15 28.0267
R26 VN.n3 VN.n2 28.0267
R27 VN.n10 VN.n9 24.4675
R28 VN.n23 VN.n22 24.4675
R29 VN.n5 VN.n4 23.9782
R30 VN.n6 VN.n1 23.9782
R31 VN.n18 VN.n17 23.9782
R32 VN.n19 VN.n14 23.9782
R33 VN.n9 VN.n1 0.48984
R34 VN.n22 VN.n14 0.48984
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 64.6042
R45 VDD2.n2 VDD2.n0 64.6042
R46 VDD2 VDD2.n5 64.6013
R47 VDD2.n4 VDD2.n3 64.0218
R48 VDD2.n4 VDD2.n2 44.086
R49 VDD2.n5 VDD2.t1 1.16726
R50 VDD2.n5 VDD2.t7 1.16726
R51 VDD2.n3 VDD2.t6 1.16726
R52 VDD2.n3 VDD2.t4 1.16726
R53 VDD2.n1 VDD2.t3 1.16726
R54 VDD2.n1 VDD2.t5 1.16726
R55 VDD2.n0 VDD2.t0 1.16726
R56 VDD2.n0 VDD2.t2 1.16726
R57 VDD2 VDD2.n4 0.696621
R58 VTAIL.n754 VTAIL.n666 289.615
R59 VTAIL.n90 VTAIL.n2 289.615
R60 VTAIL.n184 VTAIL.n96 289.615
R61 VTAIL.n280 VTAIL.n192 289.615
R62 VTAIL.n660 VTAIL.n572 289.615
R63 VTAIL.n564 VTAIL.n476 289.615
R64 VTAIL.n470 VTAIL.n382 289.615
R65 VTAIL.n374 VTAIL.n286 289.615
R66 VTAIL.n697 VTAIL.n696 185
R67 VTAIL.n694 VTAIL.n693 185
R68 VTAIL.n703 VTAIL.n702 185
R69 VTAIL.n705 VTAIL.n704 185
R70 VTAIL.n690 VTAIL.n689 185
R71 VTAIL.n711 VTAIL.n710 185
R72 VTAIL.n713 VTAIL.n712 185
R73 VTAIL.n686 VTAIL.n685 185
R74 VTAIL.n719 VTAIL.n718 185
R75 VTAIL.n721 VTAIL.n720 185
R76 VTAIL.n682 VTAIL.n681 185
R77 VTAIL.n727 VTAIL.n726 185
R78 VTAIL.n729 VTAIL.n728 185
R79 VTAIL.n678 VTAIL.n677 185
R80 VTAIL.n735 VTAIL.n734 185
R81 VTAIL.n738 VTAIL.n737 185
R82 VTAIL.n736 VTAIL.n674 185
R83 VTAIL.n743 VTAIL.n673 185
R84 VTAIL.n745 VTAIL.n744 185
R85 VTAIL.n747 VTAIL.n746 185
R86 VTAIL.n670 VTAIL.n669 185
R87 VTAIL.n753 VTAIL.n752 185
R88 VTAIL.n755 VTAIL.n754 185
R89 VTAIL.n33 VTAIL.n32 185
R90 VTAIL.n30 VTAIL.n29 185
R91 VTAIL.n39 VTAIL.n38 185
R92 VTAIL.n41 VTAIL.n40 185
R93 VTAIL.n26 VTAIL.n25 185
R94 VTAIL.n47 VTAIL.n46 185
R95 VTAIL.n49 VTAIL.n48 185
R96 VTAIL.n22 VTAIL.n21 185
R97 VTAIL.n55 VTAIL.n54 185
R98 VTAIL.n57 VTAIL.n56 185
R99 VTAIL.n18 VTAIL.n17 185
R100 VTAIL.n63 VTAIL.n62 185
R101 VTAIL.n65 VTAIL.n64 185
R102 VTAIL.n14 VTAIL.n13 185
R103 VTAIL.n71 VTAIL.n70 185
R104 VTAIL.n74 VTAIL.n73 185
R105 VTAIL.n72 VTAIL.n10 185
R106 VTAIL.n79 VTAIL.n9 185
R107 VTAIL.n81 VTAIL.n80 185
R108 VTAIL.n83 VTAIL.n82 185
R109 VTAIL.n6 VTAIL.n5 185
R110 VTAIL.n89 VTAIL.n88 185
R111 VTAIL.n91 VTAIL.n90 185
R112 VTAIL.n127 VTAIL.n126 185
R113 VTAIL.n124 VTAIL.n123 185
R114 VTAIL.n133 VTAIL.n132 185
R115 VTAIL.n135 VTAIL.n134 185
R116 VTAIL.n120 VTAIL.n119 185
R117 VTAIL.n141 VTAIL.n140 185
R118 VTAIL.n143 VTAIL.n142 185
R119 VTAIL.n116 VTAIL.n115 185
R120 VTAIL.n149 VTAIL.n148 185
R121 VTAIL.n151 VTAIL.n150 185
R122 VTAIL.n112 VTAIL.n111 185
R123 VTAIL.n157 VTAIL.n156 185
R124 VTAIL.n159 VTAIL.n158 185
R125 VTAIL.n108 VTAIL.n107 185
R126 VTAIL.n165 VTAIL.n164 185
R127 VTAIL.n168 VTAIL.n167 185
R128 VTAIL.n166 VTAIL.n104 185
R129 VTAIL.n173 VTAIL.n103 185
R130 VTAIL.n175 VTAIL.n174 185
R131 VTAIL.n177 VTAIL.n176 185
R132 VTAIL.n100 VTAIL.n99 185
R133 VTAIL.n183 VTAIL.n182 185
R134 VTAIL.n185 VTAIL.n184 185
R135 VTAIL.n223 VTAIL.n222 185
R136 VTAIL.n220 VTAIL.n219 185
R137 VTAIL.n229 VTAIL.n228 185
R138 VTAIL.n231 VTAIL.n230 185
R139 VTAIL.n216 VTAIL.n215 185
R140 VTAIL.n237 VTAIL.n236 185
R141 VTAIL.n239 VTAIL.n238 185
R142 VTAIL.n212 VTAIL.n211 185
R143 VTAIL.n245 VTAIL.n244 185
R144 VTAIL.n247 VTAIL.n246 185
R145 VTAIL.n208 VTAIL.n207 185
R146 VTAIL.n253 VTAIL.n252 185
R147 VTAIL.n255 VTAIL.n254 185
R148 VTAIL.n204 VTAIL.n203 185
R149 VTAIL.n261 VTAIL.n260 185
R150 VTAIL.n264 VTAIL.n263 185
R151 VTAIL.n262 VTAIL.n200 185
R152 VTAIL.n269 VTAIL.n199 185
R153 VTAIL.n271 VTAIL.n270 185
R154 VTAIL.n273 VTAIL.n272 185
R155 VTAIL.n196 VTAIL.n195 185
R156 VTAIL.n279 VTAIL.n278 185
R157 VTAIL.n281 VTAIL.n280 185
R158 VTAIL.n661 VTAIL.n660 185
R159 VTAIL.n659 VTAIL.n658 185
R160 VTAIL.n576 VTAIL.n575 185
R161 VTAIL.n653 VTAIL.n652 185
R162 VTAIL.n651 VTAIL.n650 185
R163 VTAIL.n649 VTAIL.n579 185
R164 VTAIL.n583 VTAIL.n580 185
R165 VTAIL.n644 VTAIL.n643 185
R166 VTAIL.n642 VTAIL.n641 185
R167 VTAIL.n585 VTAIL.n584 185
R168 VTAIL.n636 VTAIL.n635 185
R169 VTAIL.n634 VTAIL.n633 185
R170 VTAIL.n589 VTAIL.n588 185
R171 VTAIL.n628 VTAIL.n627 185
R172 VTAIL.n626 VTAIL.n625 185
R173 VTAIL.n593 VTAIL.n592 185
R174 VTAIL.n620 VTAIL.n619 185
R175 VTAIL.n618 VTAIL.n617 185
R176 VTAIL.n597 VTAIL.n596 185
R177 VTAIL.n612 VTAIL.n611 185
R178 VTAIL.n610 VTAIL.n609 185
R179 VTAIL.n601 VTAIL.n600 185
R180 VTAIL.n604 VTAIL.n603 185
R181 VTAIL.n565 VTAIL.n564 185
R182 VTAIL.n563 VTAIL.n562 185
R183 VTAIL.n480 VTAIL.n479 185
R184 VTAIL.n557 VTAIL.n556 185
R185 VTAIL.n555 VTAIL.n554 185
R186 VTAIL.n553 VTAIL.n483 185
R187 VTAIL.n487 VTAIL.n484 185
R188 VTAIL.n548 VTAIL.n547 185
R189 VTAIL.n546 VTAIL.n545 185
R190 VTAIL.n489 VTAIL.n488 185
R191 VTAIL.n540 VTAIL.n539 185
R192 VTAIL.n538 VTAIL.n537 185
R193 VTAIL.n493 VTAIL.n492 185
R194 VTAIL.n532 VTAIL.n531 185
R195 VTAIL.n530 VTAIL.n529 185
R196 VTAIL.n497 VTAIL.n496 185
R197 VTAIL.n524 VTAIL.n523 185
R198 VTAIL.n522 VTAIL.n521 185
R199 VTAIL.n501 VTAIL.n500 185
R200 VTAIL.n516 VTAIL.n515 185
R201 VTAIL.n514 VTAIL.n513 185
R202 VTAIL.n505 VTAIL.n504 185
R203 VTAIL.n508 VTAIL.n507 185
R204 VTAIL.n471 VTAIL.n470 185
R205 VTAIL.n469 VTAIL.n468 185
R206 VTAIL.n386 VTAIL.n385 185
R207 VTAIL.n463 VTAIL.n462 185
R208 VTAIL.n461 VTAIL.n460 185
R209 VTAIL.n459 VTAIL.n389 185
R210 VTAIL.n393 VTAIL.n390 185
R211 VTAIL.n454 VTAIL.n453 185
R212 VTAIL.n452 VTAIL.n451 185
R213 VTAIL.n395 VTAIL.n394 185
R214 VTAIL.n446 VTAIL.n445 185
R215 VTAIL.n444 VTAIL.n443 185
R216 VTAIL.n399 VTAIL.n398 185
R217 VTAIL.n438 VTAIL.n437 185
R218 VTAIL.n436 VTAIL.n435 185
R219 VTAIL.n403 VTAIL.n402 185
R220 VTAIL.n430 VTAIL.n429 185
R221 VTAIL.n428 VTAIL.n427 185
R222 VTAIL.n407 VTAIL.n406 185
R223 VTAIL.n422 VTAIL.n421 185
R224 VTAIL.n420 VTAIL.n419 185
R225 VTAIL.n411 VTAIL.n410 185
R226 VTAIL.n414 VTAIL.n413 185
R227 VTAIL.n375 VTAIL.n374 185
R228 VTAIL.n373 VTAIL.n372 185
R229 VTAIL.n290 VTAIL.n289 185
R230 VTAIL.n367 VTAIL.n366 185
R231 VTAIL.n365 VTAIL.n364 185
R232 VTAIL.n363 VTAIL.n293 185
R233 VTAIL.n297 VTAIL.n294 185
R234 VTAIL.n358 VTAIL.n357 185
R235 VTAIL.n356 VTAIL.n355 185
R236 VTAIL.n299 VTAIL.n298 185
R237 VTAIL.n350 VTAIL.n349 185
R238 VTAIL.n348 VTAIL.n347 185
R239 VTAIL.n303 VTAIL.n302 185
R240 VTAIL.n342 VTAIL.n341 185
R241 VTAIL.n340 VTAIL.n339 185
R242 VTAIL.n307 VTAIL.n306 185
R243 VTAIL.n334 VTAIL.n333 185
R244 VTAIL.n332 VTAIL.n331 185
R245 VTAIL.n311 VTAIL.n310 185
R246 VTAIL.n326 VTAIL.n325 185
R247 VTAIL.n324 VTAIL.n323 185
R248 VTAIL.n315 VTAIL.n314 185
R249 VTAIL.n318 VTAIL.n317 185
R250 VTAIL.t2 VTAIL.n602 147.659
R251 VTAIL.t7 VTAIL.n506 147.659
R252 VTAIL.t9 VTAIL.n412 147.659
R253 VTAIL.t8 VTAIL.n316 147.659
R254 VTAIL.t11 VTAIL.n695 147.659
R255 VTAIL.t14 VTAIL.n31 147.659
R256 VTAIL.t6 VTAIL.n125 147.659
R257 VTAIL.t4 VTAIL.n221 147.659
R258 VTAIL.n696 VTAIL.n693 104.615
R259 VTAIL.n703 VTAIL.n693 104.615
R260 VTAIL.n704 VTAIL.n703 104.615
R261 VTAIL.n704 VTAIL.n689 104.615
R262 VTAIL.n711 VTAIL.n689 104.615
R263 VTAIL.n712 VTAIL.n711 104.615
R264 VTAIL.n712 VTAIL.n685 104.615
R265 VTAIL.n719 VTAIL.n685 104.615
R266 VTAIL.n720 VTAIL.n719 104.615
R267 VTAIL.n720 VTAIL.n681 104.615
R268 VTAIL.n727 VTAIL.n681 104.615
R269 VTAIL.n728 VTAIL.n727 104.615
R270 VTAIL.n728 VTAIL.n677 104.615
R271 VTAIL.n735 VTAIL.n677 104.615
R272 VTAIL.n737 VTAIL.n735 104.615
R273 VTAIL.n737 VTAIL.n736 104.615
R274 VTAIL.n736 VTAIL.n673 104.615
R275 VTAIL.n745 VTAIL.n673 104.615
R276 VTAIL.n746 VTAIL.n745 104.615
R277 VTAIL.n746 VTAIL.n669 104.615
R278 VTAIL.n753 VTAIL.n669 104.615
R279 VTAIL.n754 VTAIL.n753 104.615
R280 VTAIL.n32 VTAIL.n29 104.615
R281 VTAIL.n39 VTAIL.n29 104.615
R282 VTAIL.n40 VTAIL.n39 104.615
R283 VTAIL.n40 VTAIL.n25 104.615
R284 VTAIL.n47 VTAIL.n25 104.615
R285 VTAIL.n48 VTAIL.n47 104.615
R286 VTAIL.n48 VTAIL.n21 104.615
R287 VTAIL.n55 VTAIL.n21 104.615
R288 VTAIL.n56 VTAIL.n55 104.615
R289 VTAIL.n56 VTAIL.n17 104.615
R290 VTAIL.n63 VTAIL.n17 104.615
R291 VTAIL.n64 VTAIL.n63 104.615
R292 VTAIL.n64 VTAIL.n13 104.615
R293 VTAIL.n71 VTAIL.n13 104.615
R294 VTAIL.n73 VTAIL.n71 104.615
R295 VTAIL.n73 VTAIL.n72 104.615
R296 VTAIL.n72 VTAIL.n9 104.615
R297 VTAIL.n81 VTAIL.n9 104.615
R298 VTAIL.n82 VTAIL.n81 104.615
R299 VTAIL.n82 VTAIL.n5 104.615
R300 VTAIL.n89 VTAIL.n5 104.615
R301 VTAIL.n90 VTAIL.n89 104.615
R302 VTAIL.n126 VTAIL.n123 104.615
R303 VTAIL.n133 VTAIL.n123 104.615
R304 VTAIL.n134 VTAIL.n133 104.615
R305 VTAIL.n134 VTAIL.n119 104.615
R306 VTAIL.n141 VTAIL.n119 104.615
R307 VTAIL.n142 VTAIL.n141 104.615
R308 VTAIL.n142 VTAIL.n115 104.615
R309 VTAIL.n149 VTAIL.n115 104.615
R310 VTAIL.n150 VTAIL.n149 104.615
R311 VTAIL.n150 VTAIL.n111 104.615
R312 VTAIL.n157 VTAIL.n111 104.615
R313 VTAIL.n158 VTAIL.n157 104.615
R314 VTAIL.n158 VTAIL.n107 104.615
R315 VTAIL.n165 VTAIL.n107 104.615
R316 VTAIL.n167 VTAIL.n165 104.615
R317 VTAIL.n167 VTAIL.n166 104.615
R318 VTAIL.n166 VTAIL.n103 104.615
R319 VTAIL.n175 VTAIL.n103 104.615
R320 VTAIL.n176 VTAIL.n175 104.615
R321 VTAIL.n176 VTAIL.n99 104.615
R322 VTAIL.n183 VTAIL.n99 104.615
R323 VTAIL.n184 VTAIL.n183 104.615
R324 VTAIL.n222 VTAIL.n219 104.615
R325 VTAIL.n229 VTAIL.n219 104.615
R326 VTAIL.n230 VTAIL.n229 104.615
R327 VTAIL.n230 VTAIL.n215 104.615
R328 VTAIL.n237 VTAIL.n215 104.615
R329 VTAIL.n238 VTAIL.n237 104.615
R330 VTAIL.n238 VTAIL.n211 104.615
R331 VTAIL.n245 VTAIL.n211 104.615
R332 VTAIL.n246 VTAIL.n245 104.615
R333 VTAIL.n246 VTAIL.n207 104.615
R334 VTAIL.n253 VTAIL.n207 104.615
R335 VTAIL.n254 VTAIL.n253 104.615
R336 VTAIL.n254 VTAIL.n203 104.615
R337 VTAIL.n261 VTAIL.n203 104.615
R338 VTAIL.n263 VTAIL.n261 104.615
R339 VTAIL.n263 VTAIL.n262 104.615
R340 VTAIL.n262 VTAIL.n199 104.615
R341 VTAIL.n271 VTAIL.n199 104.615
R342 VTAIL.n272 VTAIL.n271 104.615
R343 VTAIL.n272 VTAIL.n195 104.615
R344 VTAIL.n279 VTAIL.n195 104.615
R345 VTAIL.n280 VTAIL.n279 104.615
R346 VTAIL.n660 VTAIL.n659 104.615
R347 VTAIL.n659 VTAIL.n575 104.615
R348 VTAIL.n652 VTAIL.n575 104.615
R349 VTAIL.n652 VTAIL.n651 104.615
R350 VTAIL.n651 VTAIL.n579 104.615
R351 VTAIL.n583 VTAIL.n579 104.615
R352 VTAIL.n643 VTAIL.n583 104.615
R353 VTAIL.n643 VTAIL.n642 104.615
R354 VTAIL.n642 VTAIL.n584 104.615
R355 VTAIL.n635 VTAIL.n584 104.615
R356 VTAIL.n635 VTAIL.n634 104.615
R357 VTAIL.n634 VTAIL.n588 104.615
R358 VTAIL.n627 VTAIL.n588 104.615
R359 VTAIL.n627 VTAIL.n626 104.615
R360 VTAIL.n626 VTAIL.n592 104.615
R361 VTAIL.n619 VTAIL.n592 104.615
R362 VTAIL.n619 VTAIL.n618 104.615
R363 VTAIL.n618 VTAIL.n596 104.615
R364 VTAIL.n611 VTAIL.n596 104.615
R365 VTAIL.n611 VTAIL.n610 104.615
R366 VTAIL.n610 VTAIL.n600 104.615
R367 VTAIL.n603 VTAIL.n600 104.615
R368 VTAIL.n564 VTAIL.n563 104.615
R369 VTAIL.n563 VTAIL.n479 104.615
R370 VTAIL.n556 VTAIL.n479 104.615
R371 VTAIL.n556 VTAIL.n555 104.615
R372 VTAIL.n555 VTAIL.n483 104.615
R373 VTAIL.n487 VTAIL.n483 104.615
R374 VTAIL.n547 VTAIL.n487 104.615
R375 VTAIL.n547 VTAIL.n546 104.615
R376 VTAIL.n546 VTAIL.n488 104.615
R377 VTAIL.n539 VTAIL.n488 104.615
R378 VTAIL.n539 VTAIL.n538 104.615
R379 VTAIL.n538 VTAIL.n492 104.615
R380 VTAIL.n531 VTAIL.n492 104.615
R381 VTAIL.n531 VTAIL.n530 104.615
R382 VTAIL.n530 VTAIL.n496 104.615
R383 VTAIL.n523 VTAIL.n496 104.615
R384 VTAIL.n523 VTAIL.n522 104.615
R385 VTAIL.n522 VTAIL.n500 104.615
R386 VTAIL.n515 VTAIL.n500 104.615
R387 VTAIL.n515 VTAIL.n514 104.615
R388 VTAIL.n514 VTAIL.n504 104.615
R389 VTAIL.n507 VTAIL.n504 104.615
R390 VTAIL.n470 VTAIL.n469 104.615
R391 VTAIL.n469 VTAIL.n385 104.615
R392 VTAIL.n462 VTAIL.n385 104.615
R393 VTAIL.n462 VTAIL.n461 104.615
R394 VTAIL.n461 VTAIL.n389 104.615
R395 VTAIL.n393 VTAIL.n389 104.615
R396 VTAIL.n453 VTAIL.n393 104.615
R397 VTAIL.n453 VTAIL.n452 104.615
R398 VTAIL.n452 VTAIL.n394 104.615
R399 VTAIL.n445 VTAIL.n394 104.615
R400 VTAIL.n445 VTAIL.n444 104.615
R401 VTAIL.n444 VTAIL.n398 104.615
R402 VTAIL.n437 VTAIL.n398 104.615
R403 VTAIL.n437 VTAIL.n436 104.615
R404 VTAIL.n436 VTAIL.n402 104.615
R405 VTAIL.n429 VTAIL.n402 104.615
R406 VTAIL.n429 VTAIL.n428 104.615
R407 VTAIL.n428 VTAIL.n406 104.615
R408 VTAIL.n421 VTAIL.n406 104.615
R409 VTAIL.n421 VTAIL.n420 104.615
R410 VTAIL.n420 VTAIL.n410 104.615
R411 VTAIL.n413 VTAIL.n410 104.615
R412 VTAIL.n374 VTAIL.n373 104.615
R413 VTAIL.n373 VTAIL.n289 104.615
R414 VTAIL.n366 VTAIL.n289 104.615
R415 VTAIL.n366 VTAIL.n365 104.615
R416 VTAIL.n365 VTAIL.n293 104.615
R417 VTAIL.n297 VTAIL.n293 104.615
R418 VTAIL.n357 VTAIL.n297 104.615
R419 VTAIL.n357 VTAIL.n356 104.615
R420 VTAIL.n356 VTAIL.n298 104.615
R421 VTAIL.n349 VTAIL.n298 104.615
R422 VTAIL.n349 VTAIL.n348 104.615
R423 VTAIL.n348 VTAIL.n302 104.615
R424 VTAIL.n341 VTAIL.n302 104.615
R425 VTAIL.n341 VTAIL.n340 104.615
R426 VTAIL.n340 VTAIL.n306 104.615
R427 VTAIL.n333 VTAIL.n306 104.615
R428 VTAIL.n333 VTAIL.n332 104.615
R429 VTAIL.n332 VTAIL.n310 104.615
R430 VTAIL.n325 VTAIL.n310 104.615
R431 VTAIL.n325 VTAIL.n324 104.615
R432 VTAIL.n324 VTAIL.n314 104.615
R433 VTAIL.n317 VTAIL.n314 104.615
R434 VTAIL.n696 VTAIL.t11 52.3082
R435 VTAIL.n32 VTAIL.t14 52.3082
R436 VTAIL.n126 VTAIL.t6 52.3082
R437 VTAIL.n222 VTAIL.t4 52.3082
R438 VTAIL.n603 VTAIL.t2 52.3082
R439 VTAIL.n507 VTAIL.t7 52.3082
R440 VTAIL.n413 VTAIL.t9 52.3082
R441 VTAIL.n317 VTAIL.t8 52.3082
R442 VTAIL.n571 VTAIL.n570 47.343
R443 VTAIL.n381 VTAIL.n380 47.343
R444 VTAIL.n1 VTAIL.n0 47.3428
R445 VTAIL.n191 VTAIL.n190 47.3428
R446 VTAIL.n759 VTAIL.n758 35.4823
R447 VTAIL.n95 VTAIL.n94 35.4823
R448 VTAIL.n189 VTAIL.n188 35.4823
R449 VTAIL.n285 VTAIL.n284 35.4823
R450 VTAIL.n665 VTAIL.n664 35.4823
R451 VTAIL.n569 VTAIL.n568 35.4823
R452 VTAIL.n475 VTAIL.n474 35.4823
R453 VTAIL.n379 VTAIL.n378 35.4823
R454 VTAIL.n759 VTAIL.n665 28.2721
R455 VTAIL.n379 VTAIL.n285 28.2721
R456 VTAIL.n697 VTAIL.n695 15.6677
R457 VTAIL.n33 VTAIL.n31 15.6677
R458 VTAIL.n127 VTAIL.n125 15.6677
R459 VTAIL.n223 VTAIL.n221 15.6677
R460 VTAIL.n604 VTAIL.n602 15.6677
R461 VTAIL.n508 VTAIL.n506 15.6677
R462 VTAIL.n414 VTAIL.n412 15.6677
R463 VTAIL.n318 VTAIL.n316 15.6677
R464 VTAIL.n744 VTAIL.n743 13.1884
R465 VTAIL.n80 VTAIL.n79 13.1884
R466 VTAIL.n174 VTAIL.n173 13.1884
R467 VTAIL.n270 VTAIL.n269 13.1884
R468 VTAIL.n650 VTAIL.n649 13.1884
R469 VTAIL.n554 VTAIL.n553 13.1884
R470 VTAIL.n460 VTAIL.n459 13.1884
R471 VTAIL.n364 VTAIL.n363 13.1884
R472 VTAIL.n698 VTAIL.n694 12.8005
R473 VTAIL.n742 VTAIL.n674 12.8005
R474 VTAIL.n747 VTAIL.n672 12.8005
R475 VTAIL.n34 VTAIL.n30 12.8005
R476 VTAIL.n78 VTAIL.n10 12.8005
R477 VTAIL.n83 VTAIL.n8 12.8005
R478 VTAIL.n128 VTAIL.n124 12.8005
R479 VTAIL.n172 VTAIL.n104 12.8005
R480 VTAIL.n177 VTAIL.n102 12.8005
R481 VTAIL.n224 VTAIL.n220 12.8005
R482 VTAIL.n268 VTAIL.n200 12.8005
R483 VTAIL.n273 VTAIL.n198 12.8005
R484 VTAIL.n653 VTAIL.n578 12.8005
R485 VTAIL.n648 VTAIL.n580 12.8005
R486 VTAIL.n605 VTAIL.n601 12.8005
R487 VTAIL.n557 VTAIL.n482 12.8005
R488 VTAIL.n552 VTAIL.n484 12.8005
R489 VTAIL.n509 VTAIL.n505 12.8005
R490 VTAIL.n463 VTAIL.n388 12.8005
R491 VTAIL.n458 VTAIL.n390 12.8005
R492 VTAIL.n415 VTAIL.n411 12.8005
R493 VTAIL.n367 VTAIL.n292 12.8005
R494 VTAIL.n362 VTAIL.n294 12.8005
R495 VTAIL.n319 VTAIL.n315 12.8005
R496 VTAIL.n702 VTAIL.n701 12.0247
R497 VTAIL.n739 VTAIL.n738 12.0247
R498 VTAIL.n748 VTAIL.n670 12.0247
R499 VTAIL.n38 VTAIL.n37 12.0247
R500 VTAIL.n75 VTAIL.n74 12.0247
R501 VTAIL.n84 VTAIL.n6 12.0247
R502 VTAIL.n132 VTAIL.n131 12.0247
R503 VTAIL.n169 VTAIL.n168 12.0247
R504 VTAIL.n178 VTAIL.n100 12.0247
R505 VTAIL.n228 VTAIL.n227 12.0247
R506 VTAIL.n265 VTAIL.n264 12.0247
R507 VTAIL.n274 VTAIL.n196 12.0247
R508 VTAIL.n654 VTAIL.n576 12.0247
R509 VTAIL.n645 VTAIL.n644 12.0247
R510 VTAIL.n609 VTAIL.n608 12.0247
R511 VTAIL.n558 VTAIL.n480 12.0247
R512 VTAIL.n549 VTAIL.n548 12.0247
R513 VTAIL.n513 VTAIL.n512 12.0247
R514 VTAIL.n464 VTAIL.n386 12.0247
R515 VTAIL.n455 VTAIL.n454 12.0247
R516 VTAIL.n419 VTAIL.n418 12.0247
R517 VTAIL.n368 VTAIL.n290 12.0247
R518 VTAIL.n359 VTAIL.n358 12.0247
R519 VTAIL.n323 VTAIL.n322 12.0247
R520 VTAIL.n705 VTAIL.n692 11.249
R521 VTAIL.n734 VTAIL.n676 11.249
R522 VTAIL.n752 VTAIL.n751 11.249
R523 VTAIL.n41 VTAIL.n28 11.249
R524 VTAIL.n70 VTAIL.n12 11.249
R525 VTAIL.n88 VTAIL.n87 11.249
R526 VTAIL.n135 VTAIL.n122 11.249
R527 VTAIL.n164 VTAIL.n106 11.249
R528 VTAIL.n182 VTAIL.n181 11.249
R529 VTAIL.n231 VTAIL.n218 11.249
R530 VTAIL.n260 VTAIL.n202 11.249
R531 VTAIL.n278 VTAIL.n277 11.249
R532 VTAIL.n658 VTAIL.n657 11.249
R533 VTAIL.n641 VTAIL.n582 11.249
R534 VTAIL.n612 VTAIL.n599 11.249
R535 VTAIL.n562 VTAIL.n561 11.249
R536 VTAIL.n545 VTAIL.n486 11.249
R537 VTAIL.n516 VTAIL.n503 11.249
R538 VTAIL.n468 VTAIL.n467 11.249
R539 VTAIL.n451 VTAIL.n392 11.249
R540 VTAIL.n422 VTAIL.n409 11.249
R541 VTAIL.n372 VTAIL.n371 11.249
R542 VTAIL.n355 VTAIL.n296 11.249
R543 VTAIL.n326 VTAIL.n313 11.249
R544 VTAIL.n706 VTAIL.n690 10.4732
R545 VTAIL.n733 VTAIL.n678 10.4732
R546 VTAIL.n755 VTAIL.n668 10.4732
R547 VTAIL.n42 VTAIL.n26 10.4732
R548 VTAIL.n69 VTAIL.n14 10.4732
R549 VTAIL.n91 VTAIL.n4 10.4732
R550 VTAIL.n136 VTAIL.n120 10.4732
R551 VTAIL.n163 VTAIL.n108 10.4732
R552 VTAIL.n185 VTAIL.n98 10.4732
R553 VTAIL.n232 VTAIL.n216 10.4732
R554 VTAIL.n259 VTAIL.n204 10.4732
R555 VTAIL.n281 VTAIL.n194 10.4732
R556 VTAIL.n661 VTAIL.n574 10.4732
R557 VTAIL.n640 VTAIL.n585 10.4732
R558 VTAIL.n613 VTAIL.n597 10.4732
R559 VTAIL.n565 VTAIL.n478 10.4732
R560 VTAIL.n544 VTAIL.n489 10.4732
R561 VTAIL.n517 VTAIL.n501 10.4732
R562 VTAIL.n471 VTAIL.n384 10.4732
R563 VTAIL.n450 VTAIL.n395 10.4732
R564 VTAIL.n423 VTAIL.n407 10.4732
R565 VTAIL.n375 VTAIL.n288 10.4732
R566 VTAIL.n354 VTAIL.n299 10.4732
R567 VTAIL.n327 VTAIL.n311 10.4732
R568 VTAIL.n710 VTAIL.n709 9.69747
R569 VTAIL.n730 VTAIL.n729 9.69747
R570 VTAIL.n756 VTAIL.n666 9.69747
R571 VTAIL.n46 VTAIL.n45 9.69747
R572 VTAIL.n66 VTAIL.n65 9.69747
R573 VTAIL.n92 VTAIL.n2 9.69747
R574 VTAIL.n140 VTAIL.n139 9.69747
R575 VTAIL.n160 VTAIL.n159 9.69747
R576 VTAIL.n186 VTAIL.n96 9.69747
R577 VTAIL.n236 VTAIL.n235 9.69747
R578 VTAIL.n256 VTAIL.n255 9.69747
R579 VTAIL.n282 VTAIL.n192 9.69747
R580 VTAIL.n662 VTAIL.n572 9.69747
R581 VTAIL.n637 VTAIL.n636 9.69747
R582 VTAIL.n617 VTAIL.n616 9.69747
R583 VTAIL.n566 VTAIL.n476 9.69747
R584 VTAIL.n541 VTAIL.n540 9.69747
R585 VTAIL.n521 VTAIL.n520 9.69747
R586 VTAIL.n472 VTAIL.n382 9.69747
R587 VTAIL.n447 VTAIL.n446 9.69747
R588 VTAIL.n427 VTAIL.n426 9.69747
R589 VTAIL.n376 VTAIL.n286 9.69747
R590 VTAIL.n351 VTAIL.n350 9.69747
R591 VTAIL.n331 VTAIL.n330 9.69747
R592 VTAIL.n758 VTAIL.n757 9.45567
R593 VTAIL.n94 VTAIL.n93 9.45567
R594 VTAIL.n188 VTAIL.n187 9.45567
R595 VTAIL.n284 VTAIL.n283 9.45567
R596 VTAIL.n664 VTAIL.n663 9.45567
R597 VTAIL.n568 VTAIL.n567 9.45567
R598 VTAIL.n474 VTAIL.n473 9.45567
R599 VTAIL.n378 VTAIL.n377 9.45567
R600 VTAIL.n757 VTAIL.n756 9.3005
R601 VTAIL.n668 VTAIL.n667 9.3005
R602 VTAIL.n751 VTAIL.n750 9.3005
R603 VTAIL.n749 VTAIL.n748 9.3005
R604 VTAIL.n672 VTAIL.n671 9.3005
R605 VTAIL.n717 VTAIL.n716 9.3005
R606 VTAIL.n715 VTAIL.n714 9.3005
R607 VTAIL.n688 VTAIL.n687 9.3005
R608 VTAIL.n709 VTAIL.n708 9.3005
R609 VTAIL.n707 VTAIL.n706 9.3005
R610 VTAIL.n692 VTAIL.n691 9.3005
R611 VTAIL.n701 VTAIL.n700 9.3005
R612 VTAIL.n699 VTAIL.n698 9.3005
R613 VTAIL.n684 VTAIL.n683 9.3005
R614 VTAIL.n723 VTAIL.n722 9.3005
R615 VTAIL.n725 VTAIL.n724 9.3005
R616 VTAIL.n680 VTAIL.n679 9.3005
R617 VTAIL.n731 VTAIL.n730 9.3005
R618 VTAIL.n733 VTAIL.n732 9.3005
R619 VTAIL.n676 VTAIL.n675 9.3005
R620 VTAIL.n740 VTAIL.n739 9.3005
R621 VTAIL.n742 VTAIL.n741 9.3005
R622 VTAIL.n93 VTAIL.n92 9.3005
R623 VTAIL.n4 VTAIL.n3 9.3005
R624 VTAIL.n87 VTAIL.n86 9.3005
R625 VTAIL.n85 VTAIL.n84 9.3005
R626 VTAIL.n8 VTAIL.n7 9.3005
R627 VTAIL.n53 VTAIL.n52 9.3005
R628 VTAIL.n51 VTAIL.n50 9.3005
R629 VTAIL.n24 VTAIL.n23 9.3005
R630 VTAIL.n45 VTAIL.n44 9.3005
R631 VTAIL.n43 VTAIL.n42 9.3005
R632 VTAIL.n28 VTAIL.n27 9.3005
R633 VTAIL.n37 VTAIL.n36 9.3005
R634 VTAIL.n35 VTAIL.n34 9.3005
R635 VTAIL.n20 VTAIL.n19 9.3005
R636 VTAIL.n59 VTAIL.n58 9.3005
R637 VTAIL.n61 VTAIL.n60 9.3005
R638 VTAIL.n16 VTAIL.n15 9.3005
R639 VTAIL.n67 VTAIL.n66 9.3005
R640 VTAIL.n69 VTAIL.n68 9.3005
R641 VTAIL.n12 VTAIL.n11 9.3005
R642 VTAIL.n76 VTAIL.n75 9.3005
R643 VTAIL.n78 VTAIL.n77 9.3005
R644 VTAIL.n187 VTAIL.n186 9.3005
R645 VTAIL.n98 VTAIL.n97 9.3005
R646 VTAIL.n181 VTAIL.n180 9.3005
R647 VTAIL.n179 VTAIL.n178 9.3005
R648 VTAIL.n102 VTAIL.n101 9.3005
R649 VTAIL.n147 VTAIL.n146 9.3005
R650 VTAIL.n145 VTAIL.n144 9.3005
R651 VTAIL.n118 VTAIL.n117 9.3005
R652 VTAIL.n139 VTAIL.n138 9.3005
R653 VTAIL.n137 VTAIL.n136 9.3005
R654 VTAIL.n122 VTAIL.n121 9.3005
R655 VTAIL.n131 VTAIL.n130 9.3005
R656 VTAIL.n129 VTAIL.n128 9.3005
R657 VTAIL.n114 VTAIL.n113 9.3005
R658 VTAIL.n153 VTAIL.n152 9.3005
R659 VTAIL.n155 VTAIL.n154 9.3005
R660 VTAIL.n110 VTAIL.n109 9.3005
R661 VTAIL.n161 VTAIL.n160 9.3005
R662 VTAIL.n163 VTAIL.n162 9.3005
R663 VTAIL.n106 VTAIL.n105 9.3005
R664 VTAIL.n170 VTAIL.n169 9.3005
R665 VTAIL.n172 VTAIL.n171 9.3005
R666 VTAIL.n283 VTAIL.n282 9.3005
R667 VTAIL.n194 VTAIL.n193 9.3005
R668 VTAIL.n277 VTAIL.n276 9.3005
R669 VTAIL.n275 VTAIL.n274 9.3005
R670 VTAIL.n198 VTAIL.n197 9.3005
R671 VTAIL.n243 VTAIL.n242 9.3005
R672 VTAIL.n241 VTAIL.n240 9.3005
R673 VTAIL.n214 VTAIL.n213 9.3005
R674 VTAIL.n235 VTAIL.n234 9.3005
R675 VTAIL.n233 VTAIL.n232 9.3005
R676 VTAIL.n218 VTAIL.n217 9.3005
R677 VTAIL.n227 VTAIL.n226 9.3005
R678 VTAIL.n225 VTAIL.n224 9.3005
R679 VTAIL.n210 VTAIL.n209 9.3005
R680 VTAIL.n249 VTAIL.n248 9.3005
R681 VTAIL.n251 VTAIL.n250 9.3005
R682 VTAIL.n206 VTAIL.n205 9.3005
R683 VTAIL.n257 VTAIL.n256 9.3005
R684 VTAIL.n259 VTAIL.n258 9.3005
R685 VTAIL.n202 VTAIL.n201 9.3005
R686 VTAIL.n266 VTAIL.n265 9.3005
R687 VTAIL.n268 VTAIL.n267 9.3005
R688 VTAIL.n630 VTAIL.n629 9.3005
R689 VTAIL.n632 VTAIL.n631 9.3005
R690 VTAIL.n587 VTAIL.n586 9.3005
R691 VTAIL.n638 VTAIL.n637 9.3005
R692 VTAIL.n640 VTAIL.n639 9.3005
R693 VTAIL.n582 VTAIL.n581 9.3005
R694 VTAIL.n646 VTAIL.n645 9.3005
R695 VTAIL.n648 VTAIL.n647 9.3005
R696 VTAIL.n663 VTAIL.n662 9.3005
R697 VTAIL.n574 VTAIL.n573 9.3005
R698 VTAIL.n657 VTAIL.n656 9.3005
R699 VTAIL.n655 VTAIL.n654 9.3005
R700 VTAIL.n578 VTAIL.n577 9.3005
R701 VTAIL.n591 VTAIL.n590 9.3005
R702 VTAIL.n624 VTAIL.n623 9.3005
R703 VTAIL.n622 VTAIL.n621 9.3005
R704 VTAIL.n595 VTAIL.n594 9.3005
R705 VTAIL.n616 VTAIL.n615 9.3005
R706 VTAIL.n614 VTAIL.n613 9.3005
R707 VTAIL.n599 VTAIL.n598 9.3005
R708 VTAIL.n608 VTAIL.n607 9.3005
R709 VTAIL.n606 VTAIL.n605 9.3005
R710 VTAIL.n534 VTAIL.n533 9.3005
R711 VTAIL.n536 VTAIL.n535 9.3005
R712 VTAIL.n491 VTAIL.n490 9.3005
R713 VTAIL.n542 VTAIL.n541 9.3005
R714 VTAIL.n544 VTAIL.n543 9.3005
R715 VTAIL.n486 VTAIL.n485 9.3005
R716 VTAIL.n550 VTAIL.n549 9.3005
R717 VTAIL.n552 VTAIL.n551 9.3005
R718 VTAIL.n567 VTAIL.n566 9.3005
R719 VTAIL.n478 VTAIL.n477 9.3005
R720 VTAIL.n561 VTAIL.n560 9.3005
R721 VTAIL.n559 VTAIL.n558 9.3005
R722 VTAIL.n482 VTAIL.n481 9.3005
R723 VTAIL.n495 VTAIL.n494 9.3005
R724 VTAIL.n528 VTAIL.n527 9.3005
R725 VTAIL.n526 VTAIL.n525 9.3005
R726 VTAIL.n499 VTAIL.n498 9.3005
R727 VTAIL.n520 VTAIL.n519 9.3005
R728 VTAIL.n518 VTAIL.n517 9.3005
R729 VTAIL.n503 VTAIL.n502 9.3005
R730 VTAIL.n512 VTAIL.n511 9.3005
R731 VTAIL.n510 VTAIL.n509 9.3005
R732 VTAIL.n440 VTAIL.n439 9.3005
R733 VTAIL.n442 VTAIL.n441 9.3005
R734 VTAIL.n397 VTAIL.n396 9.3005
R735 VTAIL.n448 VTAIL.n447 9.3005
R736 VTAIL.n450 VTAIL.n449 9.3005
R737 VTAIL.n392 VTAIL.n391 9.3005
R738 VTAIL.n456 VTAIL.n455 9.3005
R739 VTAIL.n458 VTAIL.n457 9.3005
R740 VTAIL.n473 VTAIL.n472 9.3005
R741 VTAIL.n384 VTAIL.n383 9.3005
R742 VTAIL.n467 VTAIL.n466 9.3005
R743 VTAIL.n465 VTAIL.n464 9.3005
R744 VTAIL.n388 VTAIL.n387 9.3005
R745 VTAIL.n401 VTAIL.n400 9.3005
R746 VTAIL.n434 VTAIL.n433 9.3005
R747 VTAIL.n432 VTAIL.n431 9.3005
R748 VTAIL.n405 VTAIL.n404 9.3005
R749 VTAIL.n426 VTAIL.n425 9.3005
R750 VTAIL.n424 VTAIL.n423 9.3005
R751 VTAIL.n409 VTAIL.n408 9.3005
R752 VTAIL.n418 VTAIL.n417 9.3005
R753 VTAIL.n416 VTAIL.n415 9.3005
R754 VTAIL.n344 VTAIL.n343 9.3005
R755 VTAIL.n346 VTAIL.n345 9.3005
R756 VTAIL.n301 VTAIL.n300 9.3005
R757 VTAIL.n352 VTAIL.n351 9.3005
R758 VTAIL.n354 VTAIL.n353 9.3005
R759 VTAIL.n296 VTAIL.n295 9.3005
R760 VTAIL.n360 VTAIL.n359 9.3005
R761 VTAIL.n362 VTAIL.n361 9.3005
R762 VTAIL.n377 VTAIL.n376 9.3005
R763 VTAIL.n288 VTAIL.n287 9.3005
R764 VTAIL.n371 VTAIL.n370 9.3005
R765 VTAIL.n369 VTAIL.n368 9.3005
R766 VTAIL.n292 VTAIL.n291 9.3005
R767 VTAIL.n305 VTAIL.n304 9.3005
R768 VTAIL.n338 VTAIL.n337 9.3005
R769 VTAIL.n336 VTAIL.n335 9.3005
R770 VTAIL.n309 VTAIL.n308 9.3005
R771 VTAIL.n330 VTAIL.n329 9.3005
R772 VTAIL.n328 VTAIL.n327 9.3005
R773 VTAIL.n313 VTAIL.n312 9.3005
R774 VTAIL.n322 VTAIL.n321 9.3005
R775 VTAIL.n320 VTAIL.n319 9.3005
R776 VTAIL.n713 VTAIL.n688 8.92171
R777 VTAIL.n726 VTAIL.n680 8.92171
R778 VTAIL.n49 VTAIL.n24 8.92171
R779 VTAIL.n62 VTAIL.n16 8.92171
R780 VTAIL.n143 VTAIL.n118 8.92171
R781 VTAIL.n156 VTAIL.n110 8.92171
R782 VTAIL.n239 VTAIL.n214 8.92171
R783 VTAIL.n252 VTAIL.n206 8.92171
R784 VTAIL.n633 VTAIL.n587 8.92171
R785 VTAIL.n620 VTAIL.n595 8.92171
R786 VTAIL.n537 VTAIL.n491 8.92171
R787 VTAIL.n524 VTAIL.n499 8.92171
R788 VTAIL.n443 VTAIL.n397 8.92171
R789 VTAIL.n430 VTAIL.n405 8.92171
R790 VTAIL.n347 VTAIL.n301 8.92171
R791 VTAIL.n334 VTAIL.n309 8.92171
R792 VTAIL.n714 VTAIL.n686 8.14595
R793 VTAIL.n725 VTAIL.n682 8.14595
R794 VTAIL.n50 VTAIL.n22 8.14595
R795 VTAIL.n61 VTAIL.n18 8.14595
R796 VTAIL.n144 VTAIL.n116 8.14595
R797 VTAIL.n155 VTAIL.n112 8.14595
R798 VTAIL.n240 VTAIL.n212 8.14595
R799 VTAIL.n251 VTAIL.n208 8.14595
R800 VTAIL.n632 VTAIL.n589 8.14595
R801 VTAIL.n621 VTAIL.n593 8.14595
R802 VTAIL.n536 VTAIL.n493 8.14595
R803 VTAIL.n525 VTAIL.n497 8.14595
R804 VTAIL.n442 VTAIL.n399 8.14595
R805 VTAIL.n431 VTAIL.n403 8.14595
R806 VTAIL.n346 VTAIL.n303 8.14595
R807 VTAIL.n335 VTAIL.n307 8.14595
R808 VTAIL.n718 VTAIL.n717 7.3702
R809 VTAIL.n722 VTAIL.n721 7.3702
R810 VTAIL.n54 VTAIL.n53 7.3702
R811 VTAIL.n58 VTAIL.n57 7.3702
R812 VTAIL.n148 VTAIL.n147 7.3702
R813 VTAIL.n152 VTAIL.n151 7.3702
R814 VTAIL.n244 VTAIL.n243 7.3702
R815 VTAIL.n248 VTAIL.n247 7.3702
R816 VTAIL.n629 VTAIL.n628 7.3702
R817 VTAIL.n625 VTAIL.n624 7.3702
R818 VTAIL.n533 VTAIL.n532 7.3702
R819 VTAIL.n529 VTAIL.n528 7.3702
R820 VTAIL.n439 VTAIL.n438 7.3702
R821 VTAIL.n435 VTAIL.n434 7.3702
R822 VTAIL.n343 VTAIL.n342 7.3702
R823 VTAIL.n339 VTAIL.n338 7.3702
R824 VTAIL.n718 VTAIL.n684 6.59444
R825 VTAIL.n721 VTAIL.n684 6.59444
R826 VTAIL.n54 VTAIL.n20 6.59444
R827 VTAIL.n57 VTAIL.n20 6.59444
R828 VTAIL.n148 VTAIL.n114 6.59444
R829 VTAIL.n151 VTAIL.n114 6.59444
R830 VTAIL.n244 VTAIL.n210 6.59444
R831 VTAIL.n247 VTAIL.n210 6.59444
R832 VTAIL.n628 VTAIL.n591 6.59444
R833 VTAIL.n625 VTAIL.n591 6.59444
R834 VTAIL.n532 VTAIL.n495 6.59444
R835 VTAIL.n529 VTAIL.n495 6.59444
R836 VTAIL.n438 VTAIL.n401 6.59444
R837 VTAIL.n435 VTAIL.n401 6.59444
R838 VTAIL.n342 VTAIL.n305 6.59444
R839 VTAIL.n339 VTAIL.n305 6.59444
R840 VTAIL.n717 VTAIL.n686 5.81868
R841 VTAIL.n722 VTAIL.n682 5.81868
R842 VTAIL.n53 VTAIL.n22 5.81868
R843 VTAIL.n58 VTAIL.n18 5.81868
R844 VTAIL.n147 VTAIL.n116 5.81868
R845 VTAIL.n152 VTAIL.n112 5.81868
R846 VTAIL.n243 VTAIL.n212 5.81868
R847 VTAIL.n248 VTAIL.n208 5.81868
R848 VTAIL.n629 VTAIL.n589 5.81868
R849 VTAIL.n624 VTAIL.n593 5.81868
R850 VTAIL.n533 VTAIL.n493 5.81868
R851 VTAIL.n528 VTAIL.n497 5.81868
R852 VTAIL.n439 VTAIL.n399 5.81868
R853 VTAIL.n434 VTAIL.n403 5.81868
R854 VTAIL.n343 VTAIL.n303 5.81868
R855 VTAIL.n338 VTAIL.n307 5.81868
R856 VTAIL.n714 VTAIL.n713 5.04292
R857 VTAIL.n726 VTAIL.n725 5.04292
R858 VTAIL.n50 VTAIL.n49 5.04292
R859 VTAIL.n62 VTAIL.n61 5.04292
R860 VTAIL.n144 VTAIL.n143 5.04292
R861 VTAIL.n156 VTAIL.n155 5.04292
R862 VTAIL.n240 VTAIL.n239 5.04292
R863 VTAIL.n252 VTAIL.n251 5.04292
R864 VTAIL.n633 VTAIL.n632 5.04292
R865 VTAIL.n621 VTAIL.n620 5.04292
R866 VTAIL.n537 VTAIL.n536 5.04292
R867 VTAIL.n525 VTAIL.n524 5.04292
R868 VTAIL.n443 VTAIL.n442 5.04292
R869 VTAIL.n431 VTAIL.n430 5.04292
R870 VTAIL.n347 VTAIL.n346 5.04292
R871 VTAIL.n335 VTAIL.n334 5.04292
R872 VTAIL.n606 VTAIL.n602 4.38563
R873 VTAIL.n510 VTAIL.n506 4.38563
R874 VTAIL.n416 VTAIL.n412 4.38563
R875 VTAIL.n320 VTAIL.n316 4.38563
R876 VTAIL.n699 VTAIL.n695 4.38563
R877 VTAIL.n35 VTAIL.n31 4.38563
R878 VTAIL.n129 VTAIL.n125 4.38563
R879 VTAIL.n225 VTAIL.n221 4.38563
R880 VTAIL.n710 VTAIL.n688 4.26717
R881 VTAIL.n729 VTAIL.n680 4.26717
R882 VTAIL.n758 VTAIL.n666 4.26717
R883 VTAIL.n46 VTAIL.n24 4.26717
R884 VTAIL.n65 VTAIL.n16 4.26717
R885 VTAIL.n94 VTAIL.n2 4.26717
R886 VTAIL.n140 VTAIL.n118 4.26717
R887 VTAIL.n159 VTAIL.n110 4.26717
R888 VTAIL.n188 VTAIL.n96 4.26717
R889 VTAIL.n236 VTAIL.n214 4.26717
R890 VTAIL.n255 VTAIL.n206 4.26717
R891 VTAIL.n284 VTAIL.n192 4.26717
R892 VTAIL.n664 VTAIL.n572 4.26717
R893 VTAIL.n636 VTAIL.n587 4.26717
R894 VTAIL.n617 VTAIL.n595 4.26717
R895 VTAIL.n568 VTAIL.n476 4.26717
R896 VTAIL.n540 VTAIL.n491 4.26717
R897 VTAIL.n521 VTAIL.n499 4.26717
R898 VTAIL.n474 VTAIL.n382 4.26717
R899 VTAIL.n446 VTAIL.n397 4.26717
R900 VTAIL.n427 VTAIL.n405 4.26717
R901 VTAIL.n378 VTAIL.n286 4.26717
R902 VTAIL.n350 VTAIL.n301 4.26717
R903 VTAIL.n331 VTAIL.n309 4.26717
R904 VTAIL.n709 VTAIL.n690 3.49141
R905 VTAIL.n730 VTAIL.n678 3.49141
R906 VTAIL.n756 VTAIL.n755 3.49141
R907 VTAIL.n45 VTAIL.n26 3.49141
R908 VTAIL.n66 VTAIL.n14 3.49141
R909 VTAIL.n92 VTAIL.n91 3.49141
R910 VTAIL.n139 VTAIL.n120 3.49141
R911 VTAIL.n160 VTAIL.n108 3.49141
R912 VTAIL.n186 VTAIL.n185 3.49141
R913 VTAIL.n235 VTAIL.n216 3.49141
R914 VTAIL.n256 VTAIL.n204 3.49141
R915 VTAIL.n282 VTAIL.n281 3.49141
R916 VTAIL.n662 VTAIL.n661 3.49141
R917 VTAIL.n637 VTAIL.n585 3.49141
R918 VTAIL.n616 VTAIL.n597 3.49141
R919 VTAIL.n566 VTAIL.n565 3.49141
R920 VTAIL.n541 VTAIL.n489 3.49141
R921 VTAIL.n520 VTAIL.n501 3.49141
R922 VTAIL.n472 VTAIL.n471 3.49141
R923 VTAIL.n447 VTAIL.n395 3.49141
R924 VTAIL.n426 VTAIL.n407 3.49141
R925 VTAIL.n376 VTAIL.n375 3.49141
R926 VTAIL.n351 VTAIL.n299 3.49141
R927 VTAIL.n330 VTAIL.n311 3.49141
R928 VTAIL.n706 VTAIL.n705 2.71565
R929 VTAIL.n734 VTAIL.n733 2.71565
R930 VTAIL.n752 VTAIL.n668 2.71565
R931 VTAIL.n42 VTAIL.n41 2.71565
R932 VTAIL.n70 VTAIL.n69 2.71565
R933 VTAIL.n88 VTAIL.n4 2.71565
R934 VTAIL.n136 VTAIL.n135 2.71565
R935 VTAIL.n164 VTAIL.n163 2.71565
R936 VTAIL.n182 VTAIL.n98 2.71565
R937 VTAIL.n232 VTAIL.n231 2.71565
R938 VTAIL.n260 VTAIL.n259 2.71565
R939 VTAIL.n278 VTAIL.n194 2.71565
R940 VTAIL.n658 VTAIL.n574 2.71565
R941 VTAIL.n641 VTAIL.n640 2.71565
R942 VTAIL.n613 VTAIL.n612 2.71565
R943 VTAIL.n562 VTAIL.n478 2.71565
R944 VTAIL.n545 VTAIL.n544 2.71565
R945 VTAIL.n517 VTAIL.n516 2.71565
R946 VTAIL.n468 VTAIL.n384 2.71565
R947 VTAIL.n451 VTAIL.n450 2.71565
R948 VTAIL.n423 VTAIL.n422 2.71565
R949 VTAIL.n372 VTAIL.n288 2.71565
R950 VTAIL.n355 VTAIL.n354 2.71565
R951 VTAIL.n327 VTAIL.n326 2.71565
R952 VTAIL.n702 VTAIL.n692 1.93989
R953 VTAIL.n738 VTAIL.n676 1.93989
R954 VTAIL.n751 VTAIL.n670 1.93989
R955 VTAIL.n38 VTAIL.n28 1.93989
R956 VTAIL.n74 VTAIL.n12 1.93989
R957 VTAIL.n87 VTAIL.n6 1.93989
R958 VTAIL.n132 VTAIL.n122 1.93989
R959 VTAIL.n168 VTAIL.n106 1.93989
R960 VTAIL.n181 VTAIL.n100 1.93989
R961 VTAIL.n228 VTAIL.n218 1.93989
R962 VTAIL.n264 VTAIL.n202 1.93989
R963 VTAIL.n277 VTAIL.n196 1.93989
R964 VTAIL.n657 VTAIL.n576 1.93989
R965 VTAIL.n644 VTAIL.n582 1.93989
R966 VTAIL.n609 VTAIL.n599 1.93989
R967 VTAIL.n561 VTAIL.n480 1.93989
R968 VTAIL.n548 VTAIL.n486 1.93989
R969 VTAIL.n513 VTAIL.n503 1.93989
R970 VTAIL.n467 VTAIL.n386 1.93989
R971 VTAIL.n454 VTAIL.n392 1.93989
R972 VTAIL.n419 VTAIL.n409 1.93989
R973 VTAIL.n371 VTAIL.n290 1.93989
R974 VTAIL.n358 VTAIL.n296 1.93989
R975 VTAIL.n323 VTAIL.n313 1.93989
R976 VTAIL.n381 VTAIL.n379 1.27636
R977 VTAIL.n475 VTAIL.n381 1.27636
R978 VTAIL.n571 VTAIL.n569 1.27636
R979 VTAIL.n665 VTAIL.n571 1.27636
R980 VTAIL.n285 VTAIL.n191 1.27636
R981 VTAIL.n191 VTAIL.n189 1.27636
R982 VTAIL.n95 VTAIL.n1 1.27636
R983 VTAIL VTAIL.n759 1.21817
R984 VTAIL.n0 VTAIL.t12 1.16726
R985 VTAIL.n0 VTAIL.t13 1.16726
R986 VTAIL.n190 VTAIL.t0 1.16726
R987 VTAIL.n190 VTAIL.t3 1.16726
R988 VTAIL.n570 VTAIL.t5 1.16726
R989 VTAIL.n570 VTAIL.t1 1.16726
R990 VTAIL.n380 VTAIL.t10 1.16726
R991 VTAIL.n380 VTAIL.t15 1.16726
R992 VTAIL.n701 VTAIL.n694 1.16414
R993 VTAIL.n739 VTAIL.n674 1.16414
R994 VTAIL.n748 VTAIL.n747 1.16414
R995 VTAIL.n37 VTAIL.n30 1.16414
R996 VTAIL.n75 VTAIL.n10 1.16414
R997 VTAIL.n84 VTAIL.n83 1.16414
R998 VTAIL.n131 VTAIL.n124 1.16414
R999 VTAIL.n169 VTAIL.n104 1.16414
R1000 VTAIL.n178 VTAIL.n177 1.16414
R1001 VTAIL.n227 VTAIL.n220 1.16414
R1002 VTAIL.n265 VTAIL.n200 1.16414
R1003 VTAIL.n274 VTAIL.n273 1.16414
R1004 VTAIL.n654 VTAIL.n653 1.16414
R1005 VTAIL.n645 VTAIL.n580 1.16414
R1006 VTAIL.n608 VTAIL.n601 1.16414
R1007 VTAIL.n558 VTAIL.n557 1.16414
R1008 VTAIL.n549 VTAIL.n484 1.16414
R1009 VTAIL.n512 VTAIL.n505 1.16414
R1010 VTAIL.n464 VTAIL.n463 1.16414
R1011 VTAIL.n455 VTAIL.n390 1.16414
R1012 VTAIL.n418 VTAIL.n411 1.16414
R1013 VTAIL.n368 VTAIL.n367 1.16414
R1014 VTAIL.n359 VTAIL.n294 1.16414
R1015 VTAIL.n322 VTAIL.n315 1.16414
R1016 VTAIL.n569 VTAIL.n475 0.470328
R1017 VTAIL.n189 VTAIL.n95 0.470328
R1018 VTAIL.n698 VTAIL.n697 0.388379
R1019 VTAIL.n743 VTAIL.n742 0.388379
R1020 VTAIL.n744 VTAIL.n672 0.388379
R1021 VTAIL.n34 VTAIL.n33 0.388379
R1022 VTAIL.n79 VTAIL.n78 0.388379
R1023 VTAIL.n80 VTAIL.n8 0.388379
R1024 VTAIL.n128 VTAIL.n127 0.388379
R1025 VTAIL.n173 VTAIL.n172 0.388379
R1026 VTAIL.n174 VTAIL.n102 0.388379
R1027 VTAIL.n224 VTAIL.n223 0.388379
R1028 VTAIL.n269 VTAIL.n268 0.388379
R1029 VTAIL.n270 VTAIL.n198 0.388379
R1030 VTAIL.n650 VTAIL.n578 0.388379
R1031 VTAIL.n649 VTAIL.n648 0.388379
R1032 VTAIL.n605 VTAIL.n604 0.388379
R1033 VTAIL.n554 VTAIL.n482 0.388379
R1034 VTAIL.n553 VTAIL.n552 0.388379
R1035 VTAIL.n509 VTAIL.n508 0.388379
R1036 VTAIL.n460 VTAIL.n388 0.388379
R1037 VTAIL.n459 VTAIL.n458 0.388379
R1038 VTAIL.n415 VTAIL.n414 0.388379
R1039 VTAIL.n364 VTAIL.n292 0.388379
R1040 VTAIL.n363 VTAIL.n362 0.388379
R1041 VTAIL.n319 VTAIL.n318 0.388379
R1042 VTAIL.n700 VTAIL.n699 0.155672
R1043 VTAIL.n700 VTAIL.n691 0.155672
R1044 VTAIL.n707 VTAIL.n691 0.155672
R1045 VTAIL.n708 VTAIL.n707 0.155672
R1046 VTAIL.n708 VTAIL.n687 0.155672
R1047 VTAIL.n715 VTAIL.n687 0.155672
R1048 VTAIL.n716 VTAIL.n715 0.155672
R1049 VTAIL.n716 VTAIL.n683 0.155672
R1050 VTAIL.n723 VTAIL.n683 0.155672
R1051 VTAIL.n724 VTAIL.n723 0.155672
R1052 VTAIL.n724 VTAIL.n679 0.155672
R1053 VTAIL.n731 VTAIL.n679 0.155672
R1054 VTAIL.n732 VTAIL.n731 0.155672
R1055 VTAIL.n732 VTAIL.n675 0.155672
R1056 VTAIL.n740 VTAIL.n675 0.155672
R1057 VTAIL.n741 VTAIL.n740 0.155672
R1058 VTAIL.n741 VTAIL.n671 0.155672
R1059 VTAIL.n749 VTAIL.n671 0.155672
R1060 VTAIL.n750 VTAIL.n749 0.155672
R1061 VTAIL.n750 VTAIL.n667 0.155672
R1062 VTAIL.n757 VTAIL.n667 0.155672
R1063 VTAIL.n36 VTAIL.n35 0.155672
R1064 VTAIL.n36 VTAIL.n27 0.155672
R1065 VTAIL.n43 VTAIL.n27 0.155672
R1066 VTAIL.n44 VTAIL.n43 0.155672
R1067 VTAIL.n44 VTAIL.n23 0.155672
R1068 VTAIL.n51 VTAIL.n23 0.155672
R1069 VTAIL.n52 VTAIL.n51 0.155672
R1070 VTAIL.n52 VTAIL.n19 0.155672
R1071 VTAIL.n59 VTAIL.n19 0.155672
R1072 VTAIL.n60 VTAIL.n59 0.155672
R1073 VTAIL.n60 VTAIL.n15 0.155672
R1074 VTAIL.n67 VTAIL.n15 0.155672
R1075 VTAIL.n68 VTAIL.n67 0.155672
R1076 VTAIL.n68 VTAIL.n11 0.155672
R1077 VTAIL.n76 VTAIL.n11 0.155672
R1078 VTAIL.n77 VTAIL.n76 0.155672
R1079 VTAIL.n77 VTAIL.n7 0.155672
R1080 VTAIL.n85 VTAIL.n7 0.155672
R1081 VTAIL.n86 VTAIL.n85 0.155672
R1082 VTAIL.n86 VTAIL.n3 0.155672
R1083 VTAIL.n93 VTAIL.n3 0.155672
R1084 VTAIL.n130 VTAIL.n129 0.155672
R1085 VTAIL.n130 VTAIL.n121 0.155672
R1086 VTAIL.n137 VTAIL.n121 0.155672
R1087 VTAIL.n138 VTAIL.n137 0.155672
R1088 VTAIL.n138 VTAIL.n117 0.155672
R1089 VTAIL.n145 VTAIL.n117 0.155672
R1090 VTAIL.n146 VTAIL.n145 0.155672
R1091 VTAIL.n146 VTAIL.n113 0.155672
R1092 VTAIL.n153 VTAIL.n113 0.155672
R1093 VTAIL.n154 VTAIL.n153 0.155672
R1094 VTAIL.n154 VTAIL.n109 0.155672
R1095 VTAIL.n161 VTAIL.n109 0.155672
R1096 VTAIL.n162 VTAIL.n161 0.155672
R1097 VTAIL.n162 VTAIL.n105 0.155672
R1098 VTAIL.n170 VTAIL.n105 0.155672
R1099 VTAIL.n171 VTAIL.n170 0.155672
R1100 VTAIL.n171 VTAIL.n101 0.155672
R1101 VTAIL.n179 VTAIL.n101 0.155672
R1102 VTAIL.n180 VTAIL.n179 0.155672
R1103 VTAIL.n180 VTAIL.n97 0.155672
R1104 VTAIL.n187 VTAIL.n97 0.155672
R1105 VTAIL.n226 VTAIL.n225 0.155672
R1106 VTAIL.n226 VTAIL.n217 0.155672
R1107 VTAIL.n233 VTAIL.n217 0.155672
R1108 VTAIL.n234 VTAIL.n233 0.155672
R1109 VTAIL.n234 VTAIL.n213 0.155672
R1110 VTAIL.n241 VTAIL.n213 0.155672
R1111 VTAIL.n242 VTAIL.n241 0.155672
R1112 VTAIL.n242 VTAIL.n209 0.155672
R1113 VTAIL.n249 VTAIL.n209 0.155672
R1114 VTAIL.n250 VTAIL.n249 0.155672
R1115 VTAIL.n250 VTAIL.n205 0.155672
R1116 VTAIL.n257 VTAIL.n205 0.155672
R1117 VTAIL.n258 VTAIL.n257 0.155672
R1118 VTAIL.n258 VTAIL.n201 0.155672
R1119 VTAIL.n266 VTAIL.n201 0.155672
R1120 VTAIL.n267 VTAIL.n266 0.155672
R1121 VTAIL.n267 VTAIL.n197 0.155672
R1122 VTAIL.n275 VTAIL.n197 0.155672
R1123 VTAIL.n276 VTAIL.n275 0.155672
R1124 VTAIL.n276 VTAIL.n193 0.155672
R1125 VTAIL.n283 VTAIL.n193 0.155672
R1126 VTAIL.n663 VTAIL.n573 0.155672
R1127 VTAIL.n656 VTAIL.n573 0.155672
R1128 VTAIL.n656 VTAIL.n655 0.155672
R1129 VTAIL.n655 VTAIL.n577 0.155672
R1130 VTAIL.n647 VTAIL.n577 0.155672
R1131 VTAIL.n647 VTAIL.n646 0.155672
R1132 VTAIL.n646 VTAIL.n581 0.155672
R1133 VTAIL.n639 VTAIL.n581 0.155672
R1134 VTAIL.n639 VTAIL.n638 0.155672
R1135 VTAIL.n638 VTAIL.n586 0.155672
R1136 VTAIL.n631 VTAIL.n586 0.155672
R1137 VTAIL.n631 VTAIL.n630 0.155672
R1138 VTAIL.n630 VTAIL.n590 0.155672
R1139 VTAIL.n623 VTAIL.n590 0.155672
R1140 VTAIL.n623 VTAIL.n622 0.155672
R1141 VTAIL.n622 VTAIL.n594 0.155672
R1142 VTAIL.n615 VTAIL.n594 0.155672
R1143 VTAIL.n615 VTAIL.n614 0.155672
R1144 VTAIL.n614 VTAIL.n598 0.155672
R1145 VTAIL.n607 VTAIL.n598 0.155672
R1146 VTAIL.n607 VTAIL.n606 0.155672
R1147 VTAIL.n567 VTAIL.n477 0.155672
R1148 VTAIL.n560 VTAIL.n477 0.155672
R1149 VTAIL.n560 VTAIL.n559 0.155672
R1150 VTAIL.n559 VTAIL.n481 0.155672
R1151 VTAIL.n551 VTAIL.n481 0.155672
R1152 VTAIL.n551 VTAIL.n550 0.155672
R1153 VTAIL.n550 VTAIL.n485 0.155672
R1154 VTAIL.n543 VTAIL.n485 0.155672
R1155 VTAIL.n543 VTAIL.n542 0.155672
R1156 VTAIL.n542 VTAIL.n490 0.155672
R1157 VTAIL.n535 VTAIL.n490 0.155672
R1158 VTAIL.n535 VTAIL.n534 0.155672
R1159 VTAIL.n534 VTAIL.n494 0.155672
R1160 VTAIL.n527 VTAIL.n494 0.155672
R1161 VTAIL.n527 VTAIL.n526 0.155672
R1162 VTAIL.n526 VTAIL.n498 0.155672
R1163 VTAIL.n519 VTAIL.n498 0.155672
R1164 VTAIL.n519 VTAIL.n518 0.155672
R1165 VTAIL.n518 VTAIL.n502 0.155672
R1166 VTAIL.n511 VTAIL.n502 0.155672
R1167 VTAIL.n511 VTAIL.n510 0.155672
R1168 VTAIL.n473 VTAIL.n383 0.155672
R1169 VTAIL.n466 VTAIL.n383 0.155672
R1170 VTAIL.n466 VTAIL.n465 0.155672
R1171 VTAIL.n465 VTAIL.n387 0.155672
R1172 VTAIL.n457 VTAIL.n387 0.155672
R1173 VTAIL.n457 VTAIL.n456 0.155672
R1174 VTAIL.n456 VTAIL.n391 0.155672
R1175 VTAIL.n449 VTAIL.n391 0.155672
R1176 VTAIL.n449 VTAIL.n448 0.155672
R1177 VTAIL.n448 VTAIL.n396 0.155672
R1178 VTAIL.n441 VTAIL.n396 0.155672
R1179 VTAIL.n441 VTAIL.n440 0.155672
R1180 VTAIL.n440 VTAIL.n400 0.155672
R1181 VTAIL.n433 VTAIL.n400 0.155672
R1182 VTAIL.n433 VTAIL.n432 0.155672
R1183 VTAIL.n432 VTAIL.n404 0.155672
R1184 VTAIL.n425 VTAIL.n404 0.155672
R1185 VTAIL.n425 VTAIL.n424 0.155672
R1186 VTAIL.n424 VTAIL.n408 0.155672
R1187 VTAIL.n417 VTAIL.n408 0.155672
R1188 VTAIL.n417 VTAIL.n416 0.155672
R1189 VTAIL.n377 VTAIL.n287 0.155672
R1190 VTAIL.n370 VTAIL.n287 0.155672
R1191 VTAIL.n370 VTAIL.n369 0.155672
R1192 VTAIL.n369 VTAIL.n291 0.155672
R1193 VTAIL.n361 VTAIL.n291 0.155672
R1194 VTAIL.n361 VTAIL.n360 0.155672
R1195 VTAIL.n360 VTAIL.n295 0.155672
R1196 VTAIL.n353 VTAIL.n295 0.155672
R1197 VTAIL.n353 VTAIL.n352 0.155672
R1198 VTAIL.n352 VTAIL.n300 0.155672
R1199 VTAIL.n345 VTAIL.n300 0.155672
R1200 VTAIL.n345 VTAIL.n344 0.155672
R1201 VTAIL.n344 VTAIL.n304 0.155672
R1202 VTAIL.n337 VTAIL.n304 0.155672
R1203 VTAIL.n337 VTAIL.n336 0.155672
R1204 VTAIL.n336 VTAIL.n308 0.155672
R1205 VTAIL.n329 VTAIL.n308 0.155672
R1206 VTAIL.n329 VTAIL.n328 0.155672
R1207 VTAIL.n328 VTAIL.n312 0.155672
R1208 VTAIL.n321 VTAIL.n312 0.155672
R1209 VTAIL.n321 VTAIL.n320 0.155672
R1210 VTAIL VTAIL.n1 0.0586897
R1211 B.n621 B.n620 585
R1212 B.n623 B.n123 585
R1213 B.n626 B.n625 585
R1214 B.n627 B.n122 585
R1215 B.n629 B.n628 585
R1216 B.n631 B.n121 585
R1217 B.n634 B.n633 585
R1218 B.n635 B.n120 585
R1219 B.n637 B.n636 585
R1220 B.n639 B.n119 585
R1221 B.n642 B.n641 585
R1222 B.n643 B.n118 585
R1223 B.n645 B.n644 585
R1224 B.n647 B.n117 585
R1225 B.n650 B.n649 585
R1226 B.n651 B.n116 585
R1227 B.n653 B.n652 585
R1228 B.n655 B.n115 585
R1229 B.n658 B.n657 585
R1230 B.n659 B.n114 585
R1231 B.n661 B.n660 585
R1232 B.n663 B.n113 585
R1233 B.n666 B.n665 585
R1234 B.n667 B.n112 585
R1235 B.n669 B.n668 585
R1236 B.n671 B.n111 585
R1237 B.n674 B.n673 585
R1238 B.n675 B.n110 585
R1239 B.n677 B.n676 585
R1240 B.n679 B.n109 585
R1241 B.n682 B.n681 585
R1242 B.n683 B.n108 585
R1243 B.n685 B.n684 585
R1244 B.n687 B.n107 585
R1245 B.n690 B.n689 585
R1246 B.n691 B.n106 585
R1247 B.n693 B.n692 585
R1248 B.n695 B.n105 585
R1249 B.n698 B.n697 585
R1250 B.n699 B.n104 585
R1251 B.n701 B.n700 585
R1252 B.n703 B.n103 585
R1253 B.n706 B.n705 585
R1254 B.n707 B.n102 585
R1255 B.n709 B.n708 585
R1256 B.n711 B.n101 585
R1257 B.n714 B.n713 585
R1258 B.n715 B.n100 585
R1259 B.n717 B.n716 585
R1260 B.n719 B.n99 585
R1261 B.n722 B.n721 585
R1262 B.n723 B.n98 585
R1263 B.n725 B.n724 585
R1264 B.n727 B.n97 585
R1265 B.n729 B.n728 585
R1266 B.n731 B.n730 585
R1267 B.n734 B.n733 585
R1268 B.n735 B.n92 585
R1269 B.n737 B.n736 585
R1270 B.n739 B.n91 585
R1271 B.n742 B.n741 585
R1272 B.n743 B.n90 585
R1273 B.n745 B.n744 585
R1274 B.n747 B.n89 585
R1275 B.n750 B.n749 585
R1276 B.n751 B.n86 585
R1277 B.n754 B.n753 585
R1278 B.n756 B.n85 585
R1279 B.n759 B.n758 585
R1280 B.n760 B.n84 585
R1281 B.n762 B.n761 585
R1282 B.n764 B.n83 585
R1283 B.n767 B.n766 585
R1284 B.n768 B.n82 585
R1285 B.n770 B.n769 585
R1286 B.n772 B.n81 585
R1287 B.n775 B.n774 585
R1288 B.n776 B.n80 585
R1289 B.n778 B.n777 585
R1290 B.n780 B.n79 585
R1291 B.n783 B.n782 585
R1292 B.n784 B.n78 585
R1293 B.n786 B.n785 585
R1294 B.n788 B.n77 585
R1295 B.n791 B.n790 585
R1296 B.n792 B.n76 585
R1297 B.n794 B.n793 585
R1298 B.n796 B.n75 585
R1299 B.n799 B.n798 585
R1300 B.n800 B.n74 585
R1301 B.n802 B.n801 585
R1302 B.n804 B.n73 585
R1303 B.n807 B.n806 585
R1304 B.n808 B.n72 585
R1305 B.n810 B.n809 585
R1306 B.n812 B.n71 585
R1307 B.n815 B.n814 585
R1308 B.n816 B.n70 585
R1309 B.n818 B.n817 585
R1310 B.n820 B.n69 585
R1311 B.n823 B.n822 585
R1312 B.n824 B.n68 585
R1313 B.n826 B.n825 585
R1314 B.n828 B.n67 585
R1315 B.n831 B.n830 585
R1316 B.n832 B.n66 585
R1317 B.n834 B.n833 585
R1318 B.n836 B.n65 585
R1319 B.n839 B.n838 585
R1320 B.n840 B.n64 585
R1321 B.n842 B.n841 585
R1322 B.n844 B.n63 585
R1323 B.n847 B.n846 585
R1324 B.n848 B.n62 585
R1325 B.n850 B.n849 585
R1326 B.n852 B.n61 585
R1327 B.n855 B.n854 585
R1328 B.n856 B.n60 585
R1329 B.n858 B.n857 585
R1330 B.n860 B.n59 585
R1331 B.n863 B.n862 585
R1332 B.n864 B.n58 585
R1333 B.n619 B.n56 585
R1334 B.n867 B.n56 585
R1335 B.n618 B.n55 585
R1336 B.n868 B.n55 585
R1337 B.n617 B.n54 585
R1338 B.n869 B.n54 585
R1339 B.n616 B.n615 585
R1340 B.n615 B.n50 585
R1341 B.n614 B.n49 585
R1342 B.n875 B.n49 585
R1343 B.n613 B.n48 585
R1344 B.n876 B.n48 585
R1345 B.n612 B.n47 585
R1346 B.n877 B.n47 585
R1347 B.n611 B.n610 585
R1348 B.n610 B.n43 585
R1349 B.n609 B.n42 585
R1350 B.n883 B.n42 585
R1351 B.n608 B.n41 585
R1352 B.n884 B.n41 585
R1353 B.n607 B.n40 585
R1354 B.n885 B.n40 585
R1355 B.n606 B.n605 585
R1356 B.n605 B.n36 585
R1357 B.n604 B.n35 585
R1358 B.n891 B.n35 585
R1359 B.n603 B.n34 585
R1360 B.n892 B.n34 585
R1361 B.n602 B.n33 585
R1362 B.n893 B.n33 585
R1363 B.n601 B.n600 585
R1364 B.n600 B.n29 585
R1365 B.n599 B.n28 585
R1366 B.n899 B.n28 585
R1367 B.n598 B.n27 585
R1368 B.n900 B.n27 585
R1369 B.n597 B.n26 585
R1370 B.n901 B.n26 585
R1371 B.n596 B.n595 585
R1372 B.n595 B.n22 585
R1373 B.n594 B.n21 585
R1374 B.n907 B.n21 585
R1375 B.n593 B.n20 585
R1376 B.n908 B.n20 585
R1377 B.n592 B.n19 585
R1378 B.n909 B.n19 585
R1379 B.n591 B.n590 585
R1380 B.n590 B.n15 585
R1381 B.n589 B.n14 585
R1382 B.n915 B.n14 585
R1383 B.n588 B.n13 585
R1384 B.n916 B.n13 585
R1385 B.n587 B.n12 585
R1386 B.n917 B.n12 585
R1387 B.n586 B.n585 585
R1388 B.n585 B.n8 585
R1389 B.n584 B.n7 585
R1390 B.n923 B.n7 585
R1391 B.n583 B.n6 585
R1392 B.n924 B.n6 585
R1393 B.n582 B.n5 585
R1394 B.n925 B.n5 585
R1395 B.n581 B.n580 585
R1396 B.n580 B.n4 585
R1397 B.n579 B.n124 585
R1398 B.n579 B.n578 585
R1399 B.n569 B.n125 585
R1400 B.n126 B.n125 585
R1401 B.n571 B.n570 585
R1402 B.n572 B.n571 585
R1403 B.n568 B.n131 585
R1404 B.n131 B.n130 585
R1405 B.n567 B.n566 585
R1406 B.n566 B.n565 585
R1407 B.n133 B.n132 585
R1408 B.n134 B.n133 585
R1409 B.n558 B.n557 585
R1410 B.n559 B.n558 585
R1411 B.n556 B.n138 585
R1412 B.n142 B.n138 585
R1413 B.n555 B.n554 585
R1414 B.n554 B.n553 585
R1415 B.n140 B.n139 585
R1416 B.n141 B.n140 585
R1417 B.n546 B.n545 585
R1418 B.n547 B.n546 585
R1419 B.n544 B.n146 585
R1420 B.n150 B.n146 585
R1421 B.n543 B.n542 585
R1422 B.n542 B.n541 585
R1423 B.n148 B.n147 585
R1424 B.n149 B.n148 585
R1425 B.n534 B.n533 585
R1426 B.n535 B.n534 585
R1427 B.n532 B.n154 585
R1428 B.n158 B.n154 585
R1429 B.n531 B.n530 585
R1430 B.n530 B.n529 585
R1431 B.n156 B.n155 585
R1432 B.n157 B.n156 585
R1433 B.n522 B.n521 585
R1434 B.n523 B.n522 585
R1435 B.n520 B.n163 585
R1436 B.n163 B.n162 585
R1437 B.n519 B.n518 585
R1438 B.n518 B.n517 585
R1439 B.n165 B.n164 585
R1440 B.n166 B.n165 585
R1441 B.n510 B.n509 585
R1442 B.n511 B.n510 585
R1443 B.n508 B.n170 585
R1444 B.n174 B.n170 585
R1445 B.n507 B.n506 585
R1446 B.n506 B.n505 585
R1447 B.n172 B.n171 585
R1448 B.n173 B.n172 585
R1449 B.n498 B.n497 585
R1450 B.n499 B.n498 585
R1451 B.n496 B.n179 585
R1452 B.n179 B.n178 585
R1453 B.n495 B.n494 585
R1454 B.n494 B.n493 585
R1455 B.n490 B.n183 585
R1456 B.n489 B.n488 585
R1457 B.n486 B.n184 585
R1458 B.n486 B.n182 585
R1459 B.n485 B.n484 585
R1460 B.n483 B.n482 585
R1461 B.n481 B.n186 585
R1462 B.n479 B.n478 585
R1463 B.n477 B.n187 585
R1464 B.n476 B.n475 585
R1465 B.n473 B.n188 585
R1466 B.n471 B.n470 585
R1467 B.n469 B.n189 585
R1468 B.n468 B.n467 585
R1469 B.n465 B.n190 585
R1470 B.n463 B.n462 585
R1471 B.n461 B.n191 585
R1472 B.n460 B.n459 585
R1473 B.n457 B.n192 585
R1474 B.n455 B.n454 585
R1475 B.n453 B.n193 585
R1476 B.n452 B.n451 585
R1477 B.n449 B.n194 585
R1478 B.n447 B.n446 585
R1479 B.n445 B.n195 585
R1480 B.n444 B.n443 585
R1481 B.n441 B.n196 585
R1482 B.n439 B.n438 585
R1483 B.n437 B.n197 585
R1484 B.n436 B.n435 585
R1485 B.n433 B.n198 585
R1486 B.n431 B.n430 585
R1487 B.n429 B.n199 585
R1488 B.n428 B.n427 585
R1489 B.n425 B.n200 585
R1490 B.n423 B.n422 585
R1491 B.n421 B.n201 585
R1492 B.n420 B.n419 585
R1493 B.n417 B.n202 585
R1494 B.n415 B.n414 585
R1495 B.n413 B.n203 585
R1496 B.n412 B.n411 585
R1497 B.n409 B.n204 585
R1498 B.n407 B.n406 585
R1499 B.n405 B.n205 585
R1500 B.n404 B.n403 585
R1501 B.n401 B.n206 585
R1502 B.n399 B.n398 585
R1503 B.n397 B.n207 585
R1504 B.n396 B.n395 585
R1505 B.n393 B.n208 585
R1506 B.n391 B.n390 585
R1507 B.n389 B.n209 585
R1508 B.n388 B.n387 585
R1509 B.n385 B.n210 585
R1510 B.n383 B.n382 585
R1511 B.n381 B.n211 585
R1512 B.n379 B.n378 585
R1513 B.n376 B.n214 585
R1514 B.n374 B.n373 585
R1515 B.n372 B.n215 585
R1516 B.n371 B.n370 585
R1517 B.n368 B.n216 585
R1518 B.n366 B.n365 585
R1519 B.n364 B.n217 585
R1520 B.n363 B.n362 585
R1521 B.n360 B.n218 585
R1522 B.n358 B.n357 585
R1523 B.n356 B.n219 585
R1524 B.n355 B.n354 585
R1525 B.n352 B.n223 585
R1526 B.n350 B.n349 585
R1527 B.n348 B.n224 585
R1528 B.n347 B.n346 585
R1529 B.n344 B.n225 585
R1530 B.n342 B.n341 585
R1531 B.n340 B.n226 585
R1532 B.n339 B.n338 585
R1533 B.n336 B.n227 585
R1534 B.n334 B.n333 585
R1535 B.n332 B.n228 585
R1536 B.n331 B.n330 585
R1537 B.n328 B.n229 585
R1538 B.n326 B.n325 585
R1539 B.n324 B.n230 585
R1540 B.n323 B.n322 585
R1541 B.n320 B.n231 585
R1542 B.n318 B.n317 585
R1543 B.n316 B.n232 585
R1544 B.n315 B.n314 585
R1545 B.n312 B.n233 585
R1546 B.n310 B.n309 585
R1547 B.n308 B.n234 585
R1548 B.n307 B.n306 585
R1549 B.n304 B.n235 585
R1550 B.n302 B.n301 585
R1551 B.n300 B.n236 585
R1552 B.n299 B.n298 585
R1553 B.n296 B.n237 585
R1554 B.n294 B.n293 585
R1555 B.n292 B.n238 585
R1556 B.n291 B.n290 585
R1557 B.n288 B.n239 585
R1558 B.n286 B.n285 585
R1559 B.n284 B.n240 585
R1560 B.n283 B.n282 585
R1561 B.n280 B.n241 585
R1562 B.n278 B.n277 585
R1563 B.n276 B.n242 585
R1564 B.n275 B.n274 585
R1565 B.n272 B.n243 585
R1566 B.n270 B.n269 585
R1567 B.n268 B.n244 585
R1568 B.n267 B.n266 585
R1569 B.n264 B.n245 585
R1570 B.n262 B.n261 585
R1571 B.n260 B.n246 585
R1572 B.n259 B.n258 585
R1573 B.n256 B.n247 585
R1574 B.n254 B.n253 585
R1575 B.n252 B.n248 585
R1576 B.n251 B.n250 585
R1577 B.n181 B.n180 585
R1578 B.n182 B.n181 585
R1579 B.n492 B.n491 585
R1580 B.n493 B.n492 585
R1581 B.n177 B.n176 585
R1582 B.n178 B.n177 585
R1583 B.n501 B.n500 585
R1584 B.n500 B.n499 585
R1585 B.n502 B.n175 585
R1586 B.n175 B.n173 585
R1587 B.n504 B.n503 585
R1588 B.n505 B.n504 585
R1589 B.n169 B.n168 585
R1590 B.n174 B.n169 585
R1591 B.n513 B.n512 585
R1592 B.n512 B.n511 585
R1593 B.n514 B.n167 585
R1594 B.n167 B.n166 585
R1595 B.n516 B.n515 585
R1596 B.n517 B.n516 585
R1597 B.n161 B.n160 585
R1598 B.n162 B.n161 585
R1599 B.n525 B.n524 585
R1600 B.n524 B.n523 585
R1601 B.n526 B.n159 585
R1602 B.n159 B.n157 585
R1603 B.n528 B.n527 585
R1604 B.n529 B.n528 585
R1605 B.n153 B.n152 585
R1606 B.n158 B.n153 585
R1607 B.n537 B.n536 585
R1608 B.n536 B.n535 585
R1609 B.n538 B.n151 585
R1610 B.n151 B.n149 585
R1611 B.n540 B.n539 585
R1612 B.n541 B.n540 585
R1613 B.n145 B.n144 585
R1614 B.n150 B.n145 585
R1615 B.n549 B.n548 585
R1616 B.n548 B.n547 585
R1617 B.n550 B.n143 585
R1618 B.n143 B.n141 585
R1619 B.n552 B.n551 585
R1620 B.n553 B.n552 585
R1621 B.n137 B.n136 585
R1622 B.n142 B.n137 585
R1623 B.n561 B.n560 585
R1624 B.n560 B.n559 585
R1625 B.n562 B.n135 585
R1626 B.n135 B.n134 585
R1627 B.n564 B.n563 585
R1628 B.n565 B.n564 585
R1629 B.n129 B.n128 585
R1630 B.n130 B.n129 585
R1631 B.n574 B.n573 585
R1632 B.n573 B.n572 585
R1633 B.n575 B.n127 585
R1634 B.n127 B.n126 585
R1635 B.n577 B.n576 585
R1636 B.n578 B.n577 585
R1637 B.n2 B.n0 585
R1638 B.n4 B.n2 585
R1639 B.n3 B.n1 585
R1640 B.n924 B.n3 585
R1641 B.n922 B.n921 585
R1642 B.n923 B.n922 585
R1643 B.n920 B.n9 585
R1644 B.n9 B.n8 585
R1645 B.n919 B.n918 585
R1646 B.n918 B.n917 585
R1647 B.n11 B.n10 585
R1648 B.n916 B.n11 585
R1649 B.n914 B.n913 585
R1650 B.n915 B.n914 585
R1651 B.n912 B.n16 585
R1652 B.n16 B.n15 585
R1653 B.n911 B.n910 585
R1654 B.n910 B.n909 585
R1655 B.n18 B.n17 585
R1656 B.n908 B.n18 585
R1657 B.n906 B.n905 585
R1658 B.n907 B.n906 585
R1659 B.n904 B.n23 585
R1660 B.n23 B.n22 585
R1661 B.n903 B.n902 585
R1662 B.n902 B.n901 585
R1663 B.n25 B.n24 585
R1664 B.n900 B.n25 585
R1665 B.n898 B.n897 585
R1666 B.n899 B.n898 585
R1667 B.n896 B.n30 585
R1668 B.n30 B.n29 585
R1669 B.n895 B.n894 585
R1670 B.n894 B.n893 585
R1671 B.n32 B.n31 585
R1672 B.n892 B.n32 585
R1673 B.n890 B.n889 585
R1674 B.n891 B.n890 585
R1675 B.n888 B.n37 585
R1676 B.n37 B.n36 585
R1677 B.n887 B.n886 585
R1678 B.n886 B.n885 585
R1679 B.n39 B.n38 585
R1680 B.n884 B.n39 585
R1681 B.n882 B.n881 585
R1682 B.n883 B.n882 585
R1683 B.n880 B.n44 585
R1684 B.n44 B.n43 585
R1685 B.n879 B.n878 585
R1686 B.n878 B.n877 585
R1687 B.n46 B.n45 585
R1688 B.n876 B.n46 585
R1689 B.n874 B.n873 585
R1690 B.n875 B.n874 585
R1691 B.n872 B.n51 585
R1692 B.n51 B.n50 585
R1693 B.n871 B.n870 585
R1694 B.n870 B.n869 585
R1695 B.n53 B.n52 585
R1696 B.n868 B.n53 585
R1697 B.n866 B.n865 585
R1698 B.n867 B.n866 585
R1699 B.n927 B.n926 585
R1700 B.n926 B.n925 585
R1701 B.n220 B.t12 559.481
R1702 B.n212 B.t8 559.481
R1703 B.n87 B.t19 559.481
R1704 B.n93 B.t15 559.481
R1705 B.n492 B.n183 482.89
R1706 B.n866 B.n58 482.89
R1707 B.n494 B.n181 482.89
R1708 B.n621 B.n56 482.89
R1709 B.n220 B.t14 396.771
R1710 B.n93 B.t17 396.771
R1711 B.n212 B.t11 396.771
R1712 B.n87 B.t20 396.771
R1713 B.n221 B.t13 368.067
R1714 B.n94 B.t18 368.067
R1715 B.n213 B.t10 368.067
R1716 B.n88 B.t21 368.067
R1717 B.n622 B.n57 256.663
R1718 B.n624 B.n57 256.663
R1719 B.n630 B.n57 256.663
R1720 B.n632 B.n57 256.663
R1721 B.n638 B.n57 256.663
R1722 B.n640 B.n57 256.663
R1723 B.n646 B.n57 256.663
R1724 B.n648 B.n57 256.663
R1725 B.n654 B.n57 256.663
R1726 B.n656 B.n57 256.663
R1727 B.n662 B.n57 256.663
R1728 B.n664 B.n57 256.663
R1729 B.n670 B.n57 256.663
R1730 B.n672 B.n57 256.663
R1731 B.n678 B.n57 256.663
R1732 B.n680 B.n57 256.663
R1733 B.n686 B.n57 256.663
R1734 B.n688 B.n57 256.663
R1735 B.n694 B.n57 256.663
R1736 B.n696 B.n57 256.663
R1737 B.n702 B.n57 256.663
R1738 B.n704 B.n57 256.663
R1739 B.n710 B.n57 256.663
R1740 B.n712 B.n57 256.663
R1741 B.n718 B.n57 256.663
R1742 B.n720 B.n57 256.663
R1743 B.n726 B.n57 256.663
R1744 B.n96 B.n57 256.663
R1745 B.n732 B.n57 256.663
R1746 B.n738 B.n57 256.663
R1747 B.n740 B.n57 256.663
R1748 B.n746 B.n57 256.663
R1749 B.n748 B.n57 256.663
R1750 B.n755 B.n57 256.663
R1751 B.n757 B.n57 256.663
R1752 B.n763 B.n57 256.663
R1753 B.n765 B.n57 256.663
R1754 B.n771 B.n57 256.663
R1755 B.n773 B.n57 256.663
R1756 B.n779 B.n57 256.663
R1757 B.n781 B.n57 256.663
R1758 B.n787 B.n57 256.663
R1759 B.n789 B.n57 256.663
R1760 B.n795 B.n57 256.663
R1761 B.n797 B.n57 256.663
R1762 B.n803 B.n57 256.663
R1763 B.n805 B.n57 256.663
R1764 B.n811 B.n57 256.663
R1765 B.n813 B.n57 256.663
R1766 B.n819 B.n57 256.663
R1767 B.n821 B.n57 256.663
R1768 B.n827 B.n57 256.663
R1769 B.n829 B.n57 256.663
R1770 B.n835 B.n57 256.663
R1771 B.n837 B.n57 256.663
R1772 B.n843 B.n57 256.663
R1773 B.n845 B.n57 256.663
R1774 B.n851 B.n57 256.663
R1775 B.n853 B.n57 256.663
R1776 B.n859 B.n57 256.663
R1777 B.n861 B.n57 256.663
R1778 B.n487 B.n182 256.663
R1779 B.n185 B.n182 256.663
R1780 B.n480 B.n182 256.663
R1781 B.n474 B.n182 256.663
R1782 B.n472 B.n182 256.663
R1783 B.n466 B.n182 256.663
R1784 B.n464 B.n182 256.663
R1785 B.n458 B.n182 256.663
R1786 B.n456 B.n182 256.663
R1787 B.n450 B.n182 256.663
R1788 B.n448 B.n182 256.663
R1789 B.n442 B.n182 256.663
R1790 B.n440 B.n182 256.663
R1791 B.n434 B.n182 256.663
R1792 B.n432 B.n182 256.663
R1793 B.n426 B.n182 256.663
R1794 B.n424 B.n182 256.663
R1795 B.n418 B.n182 256.663
R1796 B.n416 B.n182 256.663
R1797 B.n410 B.n182 256.663
R1798 B.n408 B.n182 256.663
R1799 B.n402 B.n182 256.663
R1800 B.n400 B.n182 256.663
R1801 B.n394 B.n182 256.663
R1802 B.n392 B.n182 256.663
R1803 B.n386 B.n182 256.663
R1804 B.n384 B.n182 256.663
R1805 B.n377 B.n182 256.663
R1806 B.n375 B.n182 256.663
R1807 B.n369 B.n182 256.663
R1808 B.n367 B.n182 256.663
R1809 B.n361 B.n182 256.663
R1810 B.n359 B.n182 256.663
R1811 B.n353 B.n182 256.663
R1812 B.n351 B.n182 256.663
R1813 B.n345 B.n182 256.663
R1814 B.n343 B.n182 256.663
R1815 B.n337 B.n182 256.663
R1816 B.n335 B.n182 256.663
R1817 B.n329 B.n182 256.663
R1818 B.n327 B.n182 256.663
R1819 B.n321 B.n182 256.663
R1820 B.n319 B.n182 256.663
R1821 B.n313 B.n182 256.663
R1822 B.n311 B.n182 256.663
R1823 B.n305 B.n182 256.663
R1824 B.n303 B.n182 256.663
R1825 B.n297 B.n182 256.663
R1826 B.n295 B.n182 256.663
R1827 B.n289 B.n182 256.663
R1828 B.n287 B.n182 256.663
R1829 B.n281 B.n182 256.663
R1830 B.n279 B.n182 256.663
R1831 B.n273 B.n182 256.663
R1832 B.n271 B.n182 256.663
R1833 B.n265 B.n182 256.663
R1834 B.n263 B.n182 256.663
R1835 B.n257 B.n182 256.663
R1836 B.n255 B.n182 256.663
R1837 B.n249 B.n182 256.663
R1838 B.n492 B.n177 163.367
R1839 B.n500 B.n177 163.367
R1840 B.n500 B.n175 163.367
R1841 B.n504 B.n175 163.367
R1842 B.n504 B.n169 163.367
R1843 B.n512 B.n169 163.367
R1844 B.n512 B.n167 163.367
R1845 B.n516 B.n167 163.367
R1846 B.n516 B.n161 163.367
R1847 B.n524 B.n161 163.367
R1848 B.n524 B.n159 163.367
R1849 B.n528 B.n159 163.367
R1850 B.n528 B.n153 163.367
R1851 B.n536 B.n153 163.367
R1852 B.n536 B.n151 163.367
R1853 B.n540 B.n151 163.367
R1854 B.n540 B.n145 163.367
R1855 B.n548 B.n145 163.367
R1856 B.n548 B.n143 163.367
R1857 B.n552 B.n143 163.367
R1858 B.n552 B.n137 163.367
R1859 B.n560 B.n137 163.367
R1860 B.n560 B.n135 163.367
R1861 B.n564 B.n135 163.367
R1862 B.n564 B.n129 163.367
R1863 B.n573 B.n129 163.367
R1864 B.n573 B.n127 163.367
R1865 B.n577 B.n127 163.367
R1866 B.n577 B.n2 163.367
R1867 B.n926 B.n2 163.367
R1868 B.n926 B.n3 163.367
R1869 B.n922 B.n3 163.367
R1870 B.n922 B.n9 163.367
R1871 B.n918 B.n9 163.367
R1872 B.n918 B.n11 163.367
R1873 B.n914 B.n11 163.367
R1874 B.n914 B.n16 163.367
R1875 B.n910 B.n16 163.367
R1876 B.n910 B.n18 163.367
R1877 B.n906 B.n18 163.367
R1878 B.n906 B.n23 163.367
R1879 B.n902 B.n23 163.367
R1880 B.n902 B.n25 163.367
R1881 B.n898 B.n25 163.367
R1882 B.n898 B.n30 163.367
R1883 B.n894 B.n30 163.367
R1884 B.n894 B.n32 163.367
R1885 B.n890 B.n32 163.367
R1886 B.n890 B.n37 163.367
R1887 B.n886 B.n37 163.367
R1888 B.n886 B.n39 163.367
R1889 B.n882 B.n39 163.367
R1890 B.n882 B.n44 163.367
R1891 B.n878 B.n44 163.367
R1892 B.n878 B.n46 163.367
R1893 B.n874 B.n46 163.367
R1894 B.n874 B.n51 163.367
R1895 B.n870 B.n51 163.367
R1896 B.n870 B.n53 163.367
R1897 B.n866 B.n53 163.367
R1898 B.n488 B.n486 163.367
R1899 B.n486 B.n485 163.367
R1900 B.n482 B.n481 163.367
R1901 B.n479 B.n187 163.367
R1902 B.n475 B.n473 163.367
R1903 B.n471 B.n189 163.367
R1904 B.n467 B.n465 163.367
R1905 B.n463 B.n191 163.367
R1906 B.n459 B.n457 163.367
R1907 B.n455 B.n193 163.367
R1908 B.n451 B.n449 163.367
R1909 B.n447 B.n195 163.367
R1910 B.n443 B.n441 163.367
R1911 B.n439 B.n197 163.367
R1912 B.n435 B.n433 163.367
R1913 B.n431 B.n199 163.367
R1914 B.n427 B.n425 163.367
R1915 B.n423 B.n201 163.367
R1916 B.n419 B.n417 163.367
R1917 B.n415 B.n203 163.367
R1918 B.n411 B.n409 163.367
R1919 B.n407 B.n205 163.367
R1920 B.n403 B.n401 163.367
R1921 B.n399 B.n207 163.367
R1922 B.n395 B.n393 163.367
R1923 B.n391 B.n209 163.367
R1924 B.n387 B.n385 163.367
R1925 B.n383 B.n211 163.367
R1926 B.n378 B.n376 163.367
R1927 B.n374 B.n215 163.367
R1928 B.n370 B.n368 163.367
R1929 B.n366 B.n217 163.367
R1930 B.n362 B.n360 163.367
R1931 B.n358 B.n219 163.367
R1932 B.n354 B.n352 163.367
R1933 B.n350 B.n224 163.367
R1934 B.n346 B.n344 163.367
R1935 B.n342 B.n226 163.367
R1936 B.n338 B.n336 163.367
R1937 B.n334 B.n228 163.367
R1938 B.n330 B.n328 163.367
R1939 B.n326 B.n230 163.367
R1940 B.n322 B.n320 163.367
R1941 B.n318 B.n232 163.367
R1942 B.n314 B.n312 163.367
R1943 B.n310 B.n234 163.367
R1944 B.n306 B.n304 163.367
R1945 B.n302 B.n236 163.367
R1946 B.n298 B.n296 163.367
R1947 B.n294 B.n238 163.367
R1948 B.n290 B.n288 163.367
R1949 B.n286 B.n240 163.367
R1950 B.n282 B.n280 163.367
R1951 B.n278 B.n242 163.367
R1952 B.n274 B.n272 163.367
R1953 B.n270 B.n244 163.367
R1954 B.n266 B.n264 163.367
R1955 B.n262 B.n246 163.367
R1956 B.n258 B.n256 163.367
R1957 B.n254 B.n248 163.367
R1958 B.n250 B.n181 163.367
R1959 B.n494 B.n179 163.367
R1960 B.n498 B.n179 163.367
R1961 B.n498 B.n172 163.367
R1962 B.n506 B.n172 163.367
R1963 B.n506 B.n170 163.367
R1964 B.n510 B.n170 163.367
R1965 B.n510 B.n165 163.367
R1966 B.n518 B.n165 163.367
R1967 B.n518 B.n163 163.367
R1968 B.n522 B.n163 163.367
R1969 B.n522 B.n156 163.367
R1970 B.n530 B.n156 163.367
R1971 B.n530 B.n154 163.367
R1972 B.n534 B.n154 163.367
R1973 B.n534 B.n148 163.367
R1974 B.n542 B.n148 163.367
R1975 B.n542 B.n146 163.367
R1976 B.n546 B.n146 163.367
R1977 B.n546 B.n140 163.367
R1978 B.n554 B.n140 163.367
R1979 B.n554 B.n138 163.367
R1980 B.n558 B.n138 163.367
R1981 B.n558 B.n133 163.367
R1982 B.n566 B.n133 163.367
R1983 B.n566 B.n131 163.367
R1984 B.n571 B.n131 163.367
R1985 B.n571 B.n125 163.367
R1986 B.n579 B.n125 163.367
R1987 B.n580 B.n579 163.367
R1988 B.n580 B.n5 163.367
R1989 B.n6 B.n5 163.367
R1990 B.n7 B.n6 163.367
R1991 B.n585 B.n7 163.367
R1992 B.n585 B.n12 163.367
R1993 B.n13 B.n12 163.367
R1994 B.n14 B.n13 163.367
R1995 B.n590 B.n14 163.367
R1996 B.n590 B.n19 163.367
R1997 B.n20 B.n19 163.367
R1998 B.n21 B.n20 163.367
R1999 B.n595 B.n21 163.367
R2000 B.n595 B.n26 163.367
R2001 B.n27 B.n26 163.367
R2002 B.n28 B.n27 163.367
R2003 B.n600 B.n28 163.367
R2004 B.n600 B.n33 163.367
R2005 B.n34 B.n33 163.367
R2006 B.n35 B.n34 163.367
R2007 B.n605 B.n35 163.367
R2008 B.n605 B.n40 163.367
R2009 B.n41 B.n40 163.367
R2010 B.n42 B.n41 163.367
R2011 B.n610 B.n42 163.367
R2012 B.n610 B.n47 163.367
R2013 B.n48 B.n47 163.367
R2014 B.n49 B.n48 163.367
R2015 B.n615 B.n49 163.367
R2016 B.n615 B.n54 163.367
R2017 B.n55 B.n54 163.367
R2018 B.n56 B.n55 163.367
R2019 B.n862 B.n860 163.367
R2020 B.n858 B.n60 163.367
R2021 B.n854 B.n852 163.367
R2022 B.n850 B.n62 163.367
R2023 B.n846 B.n844 163.367
R2024 B.n842 B.n64 163.367
R2025 B.n838 B.n836 163.367
R2026 B.n834 B.n66 163.367
R2027 B.n830 B.n828 163.367
R2028 B.n826 B.n68 163.367
R2029 B.n822 B.n820 163.367
R2030 B.n818 B.n70 163.367
R2031 B.n814 B.n812 163.367
R2032 B.n810 B.n72 163.367
R2033 B.n806 B.n804 163.367
R2034 B.n802 B.n74 163.367
R2035 B.n798 B.n796 163.367
R2036 B.n794 B.n76 163.367
R2037 B.n790 B.n788 163.367
R2038 B.n786 B.n78 163.367
R2039 B.n782 B.n780 163.367
R2040 B.n778 B.n80 163.367
R2041 B.n774 B.n772 163.367
R2042 B.n770 B.n82 163.367
R2043 B.n766 B.n764 163.367
R2044 B.n762 B.n84 163.367
R2045 B.n758 B.n756 163.367
R2046 B.n754 B.n86 163.367
R2047 B.n749 B.n747 163.367
R2048 B.n745 B.n90 163.367
R2049 B.n741 B.n739 163.367
R2050 B.n737 B.n92 163.367
R2051 B.n733 B.n731 163.367
R2052 B.n728 B.n727 163.367
R2053 B.n725 B.n98 163.367
R2054 B.n721 B.n719 163.367
R2055 B.n717 B.n100 163.367
R2056 B.n713 B.n711 163.367
R2057 B.n709 B.n102 163.367
R2058 B.n705 B.n703 163.367
R2059 B.n701 B.n104 163.367
R2060 B.n697 B.n695 163.367
R2061 B.n693 B.n106 163.367
R2062 B.n689 B.n687 163.367
R2063 B.n685 B.n108 163.367
R2064 B.n681 B.n679 163.367
R2065 B.n677 B.n110 163.367
R2066 B.n673 B.n671 163.367
R2067 B.n669 B.n112 163.367
R2068 B.n665 B.n663 163.367
R2069 B.n661 B.n114 163.367
R2070 B.n657 B.n655 163.367
R2071 B.n653 B.n116 163.367
R2072 B.n649 B.n647 163.367
R2073 B.n645 B.n118 163.367
R2074 B.n641 B.n639 163.367
R2075 B.n637 B.n120 163.367
R2076 B.n633 B.n631 163.367
R2077 B.n629 B.n122 163.367
R2078 B.n625 B.n623 163.367
R2079 B.n487 B.n183 71.676
R2080 B.n485 B.n185 71.676
R2081 B.n481 B.n480 71.676
R2082 B.n474 B.n187 71.676
R2083 B.n473 B.n472 71.676
R2084 B.n466 B.n189 71.676
R2085 B.n465 B.n464 71.676
R2086 B.n458 B.n191 71.676
R2087 B.n457 B.n456 71.676
R2088 B.n450 B.n193 71.676
R2089 B.n449 B.n448 71.676
R2090 B.n442 B.n195 71.676
R2091 B.n441 B.n440 71.676
R2092 B.n434 B.n197 71.676
R2093 B.n433 B.n432 71.676
R2094 B.n426 B.n199 71.676
R2095 B.n425 B.n424 71.676
R2096 B.n418 B.n201 71.676
R2097 B.n417 B.n416 71.676
R2098 B.n410 B.n203 71.676
R2099 B.n409 B.n408 71.676
R2100 B.n402 B.n205 71.676
R2101 B.n401 B.n400 71.676
R2102 B.n394 B.n207 71.676
R2103 B.n393 B.n392 71.676
R2104 B.n386 B.n209 71.676
R2105 B.n385 B.n384 71.676
R2106 B.n377 B.n211 71.676
R2107 B.n376 B.n375 71.676
R2108 B.n369 B.n215 71.676
R2109 B.n368 B.n367 71.676
R2110 B.n361 B.n217 71.676
R2111 B.n360 B.n359 71.676
R2112 B.n353 B.n219 71.676
R2113 B.n352 B.n351 71.676
R2114 B.n345 B.n224 71.676
R2115 B.n344 B.n343 71.676
R2116 B.n337 B.n226 71.676
R2117 B.n336 B.n335 71.676
R2118 B.n329 B.n228 71.676
R2119 B.n328 B.n327 71.676
R2120 B.n321 B.n230 71.676
R2121 B.n320 B.n319 71.676
R2122 B.n313 B.n232 71.676
R2123 B.n312 B.n311 71.676
R2124 B.n305 B.n234 71.676
R2125 B.n304 B.n303 71.676
R2126 B.n297 B.n236 71.676
R2127 B.n296 B.n295 71.676
R2128 B.n289 B.n238 71.676
R2129 B.n288 B.n287 71.676
R2130 B.n281 B.n240 71.676
R2131 B.n280 B.n279 71.676
R2132 B.n273 B.n242 71.676
R2133 B.n272 B.n271 71.676
R2134 B.n265 B.n244 71.676
R2135 B.n264 B.n263 71.676
R2136 B.n257 B.n246 71.676
R2137 B.n256 B.n255 71.676
R2138 B.n249 B.n248 71.676
R2139 B.n861 B.n58 71.676
R2140 B.n860 B.n859 71.676
R2141 B.n853 B.n60 71.676
R2142 B.n852 B.n851 71.676
R2143 B.n845 B.n62 71.676
R2144 B.n844 B.n843 71.676
R2145 B.n837 B.n64 71.676
R2146 B.n836 B.n835 71.676
R2147 B.n829 B.n66 71.676
R2148 B.n828 B.n827 71.676
R2149 B.n821 B.n68 71.676
R2150 B.n820 B.n819 71.676
R2151 B.n813 B.n70 71.676
R2152 B.n812 B.n811 71.676
R2153 B.n805 B.n72 71.676
R2154 B.n804 B.n803 71.676
R2155 B.n797 B.n74 71.676
R2156 B.n796 B.n795 71.676
R2157 B.n789 B.n76 71.676
R2158 B.n788 B.n787 71.676
R2159 B.n781 B.n78 71.676
R2160 B.n780 B.n779 71.676
R2161 B.n773 B.n80 71.676
R2162 B.n772 B.n771 71.676
R2163 B.n765 B.n82 71.676
R2164 B.n764 B.n763 71.676
R2165 B.n757 B.n84 71.676
R2166 B.n756 B.n755 71.676
R2167 B.n748 B.n86 71.676
R2168 B.n747 B.n746 71.676
R2169 B.n740 B.n90 71.676
R2170 B.n739 B.n738 71.676
R2171 B.n732 B.n92 71.676
R2172 B.n731 B.n96 71.676
R2173 B.n727 B.n726 71.676
R2174 B.n720 B.n98 71.676
R2175 B.n719 B.n718 71.676
R2176 B.n712 B.n100 71.676
R2177 B.n711 B.n710 71.676
R2178 B.n704 B.n102 71.676
R2179 B.n703 B.n702 71.676
R2180 B.n696 B.n104 71.676
R2181 B.n695 B.n694 71.676
R2182 B.n688 B.n106 71.676
R2183 B.n687 B.n686 71.676
R2184 B.n680 B.n108 71.676
R2185 B.n679 B.n678 71.676
R2186 B.n672 B.n110 71.676
R2187 B.n671 B.n670 71.676
R2188 B.n664 B.n112 71.676
R2189 B.n663 B.n662 71.676
R2190 B.n656 B.n114 71.676
R2191 B.n655 B.n654 71.676
R2192 B.n648 B.n116 71.676
R2193 B.n647 B.n646 71.676
R2194 B.n640 B.n118 71.676
R2195 B.n639 B.n638 71.676
R2196 B.n632 B.n120 71.676
R2197 B.n631 B.n630 71.676
R2198 B.n624 B.n122 71.676
R2199 B.n623 B.n622 71.676
R2200 B.n622 B.n621 71.676
R2201 B.n625 B.n624 71.676
R2202 B.n630 B.n629 71.676
R2203 B.n633 B.n632 71.676
R2204 B.n638 B.n637 71.676
R2205 B.n641 B.n640 71.676
R2206 B.n646 B.n645 71.676
R2207 B.n649 B.n648 71.676
R2208 B.n654 B.n653 71.676
R2209 B.n657 B.n656 71.676
R2210 B.n662 B.n661 71.676
R2211 B.n665 B.n664 71.676
R2212 B.n670 B.n669 71.676
R2213 B.n673 B.n672 71.676
R2214 B.n678 B.n677 71.676
R2215 B.n681 B.n680 71.676
R2216 B.n686 B.n685 71.676
R2217 B.n689 B.n688 71.676
R2218 B.n694 B.n693 71.676
R2219 B.n697 B.n696 71.676
R2220 B.n702 B.n701 71.676
R2221 B.n705 B.n704 71.676
R2222 B.n710 B.n709 71.676
R2223 B.n713 B.n712 71.676
R2224 B.n718 B.n717 71.676
R2225 B.n721 B.n720 71.676
R2226 B.n726 B.n725 71.676
R2227 B.n728 B.n96 71.676
R2228 B.n733 B.n732 71.676
R2229 B.n738 B.n737 71.676
R2230 B.n741 B.n740 71.676
R2231 B.n746 B.n745 71.676
R2232 B.n749 B.n748 71.676
R2233 B.n755 B.n754 71.676
R2234 B.n758 B.n757 71.676
R2235 B.n763 B.n762 71.676
R2236 B.n766 B.n765 71.676
R2237 B.n771 B.n770 71.676
R2238 B.n774 B.n773 71.676
R2239 B.n779 B.n778 71.676
R2240 B.n782 B.n781 71.676
R2241 B.n787 B.n786 71.676
R2242 B.n790 B.n789 71.676
R2243 B.n795 B.n794 71.676
R2244 B.n798 B.n797 71.676
R2245 B.n803 B.n802 71.676
R2246 B.n806 B.n805 71.676
R2247 B.n811 B.n810 71.676
R2248 B.n814 B.n813 71.676
R2249 B.n819 B.n818 71.676
R2250 B.n822 B.n821 71.676
R2251 B.n827 B.n826 71.676
R2252 B.n830 B.n829 71.676
R2253 B.n835 B.n834 71.676
R2254 B.n838 B.n837 71.676
R2255 B.n843 B.n842 71.676
R2256 B.n846 B.n845 71.676
R2257 B.n851 B.n850 71.676
R2258 B.n854 B.n853 71.676
R2259 B.n859 B.n858 71.676
R2260 B.n862 B.n861 71.676
R2261 B.n488 B.n487 71.676
R2262 B.n482 B.n185 71.676
R2263 B.n480 B.n479 71.676
R2264 B.n475 B.n474 71.676
R2265 B.n472 B.n471 71.676
R2266 B.n467 B.n466 71.676
R2267 B.n464 B.n463 71.676
R2268 B.n459 B.n458 71.676
R2269 B.n456 B.n455 71.676
R2270 B.n451 B.n450 71.676
R2271 B.n448 B.n447 71.676
R2272 B.n443 B.n442 71.676
R2273 B.n440 B.n439 71.676
R2274 B.n435 B.n434 71.676
R2275 B.n432 B.n431 71.676
R2276 B.n427 B.n426 71.676
R2277 B.n424 B.n423 71.676
R2278 B.n419 B.n418 71.676
R2279 B.n416 B.n415 71.676
R2280 B.n411 B.n410 71.676
R2281 B.n408 B.n407 71.676
R2282 B.n403 B.n402 71.676
R2283 B.n400 B.n399 71.676
R2284 B.n395 B.n394 71.676
R2285 B.n392 B.n391 71.676
R2286 B.n387 B.n386 71.676
R2287 B.n384 B.n383 71.676
R2288 B.n378 B.n377 71.676
R2289 B.n375 B.n374 71.676
R2290 B.n370 B.n369 71.676
R2291 B.n367 B.n366 71.676
R2292 B.n362 B.n361 71.676
R2293 B.n359 B.n358 71.676
R2294 B.n354 B.n353 71.676
R2295 B.n351 B.n350 71.676
R2296 B.n346 B.n345 71.676
R2297 B.n343 B.n342 71.676
R2298 B.n338 B.n337 71.676
R2299 B.n335 B.n334 71.676
R2300 B.n330 B.n329 71.676
R2301 B.n327 B.n326 71.676
R2302 B.n322 B.n321 71.676
R2303 B.n319 B.n318 71.676
R2304 B.n314 B.n313 71.676
R2305 B.n311 B.n310 71.676
R2306 B.n306 B.n305 71.676
R2307 B.n303 B.n302 71.676
R2308 B.n298 B.n297 71.676
R2309 B.n295 B.n294 71.676
R2310 B.n290 B.n289 71.676
R2311 B.n287 B.n286 71.676
R2312 B.n282 B.n281 71.676
R2313 B.n279 B.n278 71.676
R2314 B.n274 B.n273 71.676
R2315 B.n271 B.n270 71.676
R2316 B.n266 B.n265 71.676
R2317 B.n263 B.n262 71.676
R2318 B.n258 B.n257 71.676
R2319 B.n255 B.n254 71.676
R2320 B.n250 B.n249 71.676
R2321 B.n222 B.n221 59.5399
R2322 B.n380 B.n213 59.5399
R2323 B.n752 B.n88 59.5399
R2324 B.n95 B.n94 59.5399
R2325 B.n493 B.n182 56.8672
R2326 B.n867 B.n57 56.8672
R2327 B.n493 B.n178 33.626
R2328 B.n499 B.n178 33.626
R2329 B.n499 B.n173 33.626
R2330 B.n505 B.n173 33.626
R2331 B.n505 B.n174 33.626
R2332 B.n511 B.n166 33.626
R2333 B.n517 B.n166 33.626
R2334 B.n517 B.n162 33.626
R2335 B.n523 B.n162 33.626
R2336 B.n523 B.n157 33.626
R2337 B.n529 B.n157 33.626
R2338 B.n529 B.n158 33.626
R2339 B.n535 B.n149 33.626
R2340 B.n541 B.n149 33.626
R2341 B.n541 B.n150 33.626
R2342 B.n547 B.n141 33.626
R2343 B.n553 B.n141 33.626
R2344 B.n553 B.n142 33.626
R2345 B.n559 B.n134 33.626
R2346 B.n565 B.n134 33.626
R2347 B.n565 B.n130 33.626
R2348 B.n572 B.n130 33.626
R2349 B.n578 B.n126 33.626
R2350 B.n578 B.n4 33.626
R2351 B.n925 B.n4 33.626
R2352 B.n925 B.n924 33.626
R2353 B.n924 B.n923 33.626
R2354 B.n923 B.n8 33.626
R2355 B.n917 B.n916 33.626
R2356 B.n916 B.n915 33.626
R2357 B.n915 B.n15 33.626
R2358 B.n909 B.n15 33.626
R2359 B.n908 B.n907 33.626
R2360 B.n907 B.n22 33.626
R2361 B.n901 B.n22 33.626
R2362 B.n900 B.n899 33.626
R2363 B.n899 B.n29 33.626
R2364 B.n893 B.n29 33.626
R2365 B.n892 B.n891 33.626
R2366 B.n891 B.n36 33.626
R2367 B.n885 B.n36 33.626
R2368 B.n885 B.n884 33.626
R2369 B.n884 B.n883 33.626
R2370 B.n883 B.n43 33.626
R2371 B.n877 B.n43 33.626
R2372 B.n876 B.n875 33.626
R2373 B.n875 B.n50 33.626
R2374 B.n869 B.n50 33.626
R2375 B.n869 B.n868 33.626
R2376 B.n868 B.n867 33.626
R2377 B.n865 B.n864 31.3761
R2378 B.n620 B.n619 31.3761
R2379 B.n495 B.n180 31.3761
R2380 B.n491 B.n490 31.3761
R2381 B.n142 B.t3 29.1756
R2382 B.t5 B.n908 29.1756
R2383 B.n221 B.n220 28.7035
R2384 B.n213 B.n212 28.7035
R2385 B.n88 B.n87 28.7035
R2386 B.n94 B.n93 28.7035
R2387 B.n535 B.t4 28.1866
R2388 B.n893 B.t2 28.1866
R2389 B.t6 B.n126 26.2086
R2390 B.t7 B.n8 26.2086
R2391 B.n174 B.t9 20.2747
R2392 B.t16 B.n876 20.2747
R2393 B B.n927 18.0485
R2394 B.n150 B.t0 17.3078
R2395 B.t1 B.n900 17.3078
R2396 B.n547 B.t0 16.3188
R2397 B.n901 B.t1 16.3188
R2398 B.n511 B.t9 13.3518
R2399 B.n877 B.t16 13.3518
R2400 B.n864 B.n863 10.6151
R2401 B.n863 B.n59 10.6151
R2402 B.n857 B.n59 10.6151
R2403 B.n857 B.n856 10.6151
R2404 B.n856 B.n855 10.6151
R2405 B.n855 B.n61 10.6151
R2406 B.n849 B.n61 10.6151
R2407 B.n849 B.n848 10.6151
R2408 B.n848 B.n847 10.6151
R2409 B.n847 B.n63 10.6151
R2410 B.n841 B.n63 10.6151
R2411 B.n841 B.n840 10.6151
R2412 B.n840 B.n839 10.6151
R2413 B.n839 B.n65 10.6151
R2414 B.n833 B.n65 10.6151
R2415 B.n833 B.n832 10.6151
R2416 B.n832 B.n831 10.6151
R2417 B.n831 B.n67 10.6151
R2418 B.n825 B.n67 10.6151
R2419 B.n825 B.n824 10.6151
R2420 B.n824 B.n823 10.6151
R2421 B.n823 B.n69 10.6151
R2422 B.n817 B.n69 10.6151
R2423 B.n817 B.n816 10.6151
R2424 B.n816 B.n815 10.6151
R2425 B.n815 B.n71 10.6151
R2426 B.n809 B.n71 10.6151
R2427 B.n809 B.n808 10.6151
R2428 B.n808 B.n807 10.6151
R2429 B.n807 B.n73 10.6151
R2430 B.n801 B.n73 10.6151
R2431 B.n801 B.n800 10.6151
R2432 B.n800 B.n799 10.6151
R2433 B.n799 B.n75 10.6151
R2434 B.n793 B.n75 10.6151
R2435 B.n793 B.n792 10.6151
R2436 B.n792 B.n791 10.6151
R2437 B.n791 B.n77 10.6151
R2438 B.n785 B.n77 10.6151
R2439 B.n785 B.n784 10.6151
R2440 B.n784 B.n783 10.6151
R2441 B.n783 B.n79 10.6151
R2442 B.n777 B.n79 10.6151
R2443 B.n777 B.n776 10.6151
R2444 B.n776 B.n775 10.6151
R2445 B.n775 B.n81 10.6151
R2446 B.n769 B.n81 10.6151
R2447 B.n769 B.n768 10.6151
R2448 B.n768 B.n767 10.6151
R2449 B.n767 B.n83 10.6151
R2450 B.n761 B.n83 10.6151
R2451 B.n761 B.n760 10.6151
R2452 B.n760 B.n759 10.6151
R2453 B.n759 B.n85 10.6151
R2454 B.n753 B.n85 10.6151
R2455 B.n751 B.n750 10.6151
R2456 B.n750 B.n89 10.6151
R2457 B.n744 B.n89 10.6151
R2458 B.n744 B.n743 10.6151
R2459 B.n743 B.n742 10.6151
R2460 B.n742 B.n91 10.6151
R2461 B.n736 B.n91 10.6151
R2462 B.n736 B.n735 10.6151
R2463 B.n735 B.n734 10.6151
R2464 B.n730 B.n729 10.6151
R2465 B.n729 B.n97 10.6151
R2466 B.n724 B.n97 10.6151
R2467 B.n724 B.n723 10.6151
R2468 B.n723 B.n722 10.6151
R2469 B.n722 B.n99 10.6151
R2470 B.n716 B.n99 10.6151
R2471 B.n716 B.n715 10.6151
R2472 B.n715 B.n714 10.6151
R2473 B.n714 B.n101 10.6151
R2474 B.n708 B.n101 10.6151
R2475 B.n708 B.n707 10.6151
R2476 B.n707 B.n706 10.6151
R2477 B.n706 B.n103 10.6151
R2478 B.n700 B.n103 10.6151
R2479 B.n700 B.n699 10.6151
R2480 B.n699 B.n698 10.6151
R2481 B.n698 B.n105 10.6151
R2482 B.n692 B.n105 10.6151
R2483 B.n692 B.n691 10.6151
R2484 B.n691 B.n690 10.6151
R2485 B.n690 B.n107 10.6151
R2486 B.n684 B.n107 10.6151
R2487 B.n684 B.n683 10.6151
R2488 B.n683 B.n682 10.6151
R2489 B.n682 B.n109 10.6151
R2490 B.n676 B.n109 10.6151
R2491 B.n676 B.n675 10.6151
R2492 B.n675 B.n674 10.6151
R2493 B.n674 B.n111 10.6151
R2494 B.n668 B.n111 10.6151
R2495 B.n668 B.n667 10.6151
R2496 B.n667 B.n666 10.6151
R2497 B.n666 B.n113 10.6151
R2498 B.n660 B.n113 10.6151
R2499 B.n660 B.n659 10.6151
R2500 B.n659 B.n658 10.6151
R2501 B.n658 B.n115 10.6151
R2502 B.n652 B.n115 10.6151
R2503 B.n652 B.n651 10.6151
R2504 B.n651 B.n650 10.6151
R2505 B.n650 B.n117 10.6151
R2506 B.n644 B.n117 10.6151
R2507 B.n644 B.n643 10.6151
R2508 B.n643 B.n642 10.6151
R2509 B.n642 B.n119 10.6151
R2510 B.n636 B.n119 10.6151
R2511 B.n636 B.n635 10.6151
R2512 B.n635 B.n634 10.6151
R2513 B.n634 B.n121 10.6151
R2514 B.n628 B.n121 10.6151
R2515 B.n628 B.n627 10.6151
R2516 B.n627 B.n626 10.6151
R2517 B.n626 B.n123 10.6151
R2518 B.n620 B.n123 10.6151
R2519 B.n496 B.n495 10.6151
R2520 B.n497 B.n496 10.6151
R2521 B.n497 B.n171 10.6151
R2522 B.n507 B.n171 10.6151
R2523 B.n508 B.n507 10.6151
R2524 B.n509 B.n508 10.6151
R2525 B.n509 B.n164 10.6151
R2526 B.n519 B.n164 10.6151
R2527 B.n520 B.n519 10.6151
R2528 B.n521 B.n520 10.6151
R2529 B.n521 B.n155 10.6151
R2530 B.n531 B.n155 10.6151
R2531 B.n532 B.n531 10.6151
R2532 B.n533 B.n532 10.6151
R2533 B.n533 B.n147 10.6151
R2534 B.n543 B.n147 10.6151
R2535 B.n544 B.n543 10.6151
R2536 B.n545 B.n544 10.6151
R2537 B.n545 B.n139 10.6151
R2538 B.n555 B.n139 10.6151
R2539 B.n556 B.n555 10.6151
R2540 B.n557 B.n556 10.6151
R2541 B.n557 B.n132 10.6151
R2542 B.n567 B.n132 10.6151
R2543 B.n568 B.n567 10.6151
R2544 B.n570 B.n568 10.6151
R2545 B.n570 B.n569 10.6151
R2546 B.n569 B.n124 10.6151
R2547 B.n581 B.n124 10.6151
R2548 B.n582 B.n581 10.6151
R2549 B.n583 B.n582 10.6151
R2550 B.n584 B.n583 10.6151
R2551 B.n586 B.n584 10.6151
R2552 B.n587 B.n586 10.6151
R2553 B.n588 B.n587 10.6151
R2554 B.n589 B.n588 10.6151
R2555 B.n591 B.n589 10.6151
R2556 B.n592 B.n591 10.6151
R2557 B.n593 B.n592 10.6151
R2558 B.n594 B.n593 10.6151
R2559 B.n596 B.n594 10.6151
R2560 B.n597 B.n596 10.6151
R2561 B.n598 B.n597 10.6151
R2562 B.n599 B.n598 10.6151
R2563 B.n601 B.n599 10.6151
R2564 B.n602 B.n601 10.6151
R2565 B.n603 B.n602 10.6151
R2566 B.n604 B.n603 10.6151
R2567 B.n606 B.n604 10.6151
R2568 B.n607 B.n606 10.6151
R2569 B.n608 B.n607 10.6151
R2570 B.n609 B.n608 10.6151
R2571 B.n611 B.n609 10.6151
R2572 B.n612 B.n611 10.6151
R2573 B.n613 B.n612 10.6151
R2574 B.n614 B.n613 10.6151
R2575 B.n616 B.n614 10.6151
R2576 B.n617 B.n616 10.6151
R2577 B.n618 B.n617 10.6151
R2578 B.n619 B.n618 10.6151
R2579 B.n490 B.n489 10.6151
R2580 B.n489 B.n184 10.6151
R2581 B.n484 B.n184 10.6151
R2582 B.n484 B.n483 10.6151
R2583 B.n483 B.n186 10.6151
R2584 B.n478 B.n186 10.6151
R2585 B.n478 B.n477 10.6151
R2586 B.n477 B.n476 10.6151
R2587 B.n476 B.n188 10.6151
R2588 B.n470 B.n188 10.6151
R2589 B.n470 B.n469 10.6151
R2590 B.n469 B.n468 10.6151
R2591 B.n468 B.n190 10.6151
R2592 B.n462 B.n190 10.6151
R2593 B.n462 B.n461 10.6151
R2594 B.n461 B.n460 10.6151
R2595 B.n460 B.n192 10.6151
R2596 B.n454 B.n192 10.6151
R2597 B.n454 B.n453 10.6151
R2598 B.n453 B.n452 10.6151
R2599 B.n452 B.n194 10.6151
R2600 B.n446 B.n194 10.6151
R2601 B.n446 B.n445 10.6151
R2602 B.n445 B.n444 10.6151
R2603 B.n444 B.n196 10.6151
R2604 B.n438 B.n196 10.6151
R2605 B.n438 B.n437 10.6151
R2606 B.n437 B.n436 10.6151
R2607 B.n436 B.n198 10.6151
R2608 B.n430 B.n198 10.6151
R2609 B.n430 B.n429 10.6151
R2610 B.n429 B.n428 10.6151
R2611 B.n428 B.n200 10.6151
R2612 B.n422 B.n200 10.6151
R2613 B.n422 B.n421 10.6151
R2614 B.n421 B.n420 10.6151
R2615 B.n420 B.n202 10.6151
R2616 B.n414 B.n202 10.6151
R2617 B.n414 B.n413 10.6151
R2618 B.n413 B.n412 10.6151
R2619 B.n412 B.n204 10.6151
R2620 B.n406 B.n204 10.6151
R2621 B.n406 B.n405 10.6151
R2622 B.n405 B.n404 10.6151
R2623 B.n404 B.n206 10.6151
R2624 B.n398 B.n206 10.6151
R2625 B.n398 B.n397 10.6151
R2626 B.n397 B.n396 10.6151
R2627 B.n396 B.n208 10.6151
R2628 B.n390 B.n208 10.6151
R2629 B.n390 B.n389 10.6151
R2630 B.n389 B.n388 10.6151
R2631 B.n388 B.n210 10.6151
R2632 B.n382 B.n210 10.6151
R2633 B.n382 B.n381 10.6151
R2634 B.n379 B.n214 10.6151
R2635 B.n373 B.n214 10.6151
R2636 B.n373 B.n372 10.6151
R2637 B.n372 B.n371 10.6151
R2638 B.n371 B.n216 10.6151
R2639 B.n365 B.n216 10.6151
R2640 B.n365 B.n364 10.6151
R2641 B.n364 B.n363 10.6151
R2642 B.n363 B.n218 10.6151
R2643 B.n357 B.n356 10.6151
R2644 B.n356 B.n355 10.6151
R2645 B.n355 B.n223 10.6151
R2646 B.n349 B.n223 10.6151
R2647 B.n349 B.n348 10.6151
R2648 B.n348 B.n347 10.6151
R2649 B.n347 B.n225 10.6151
R2650 B.n341 B.n225 10.6151
R2651 B.n341 B.n340 10.6151
R2652 B.n340 B.n339 10.6151
R2653 B.n339 B.n227 10.6151
R2654 B.n333 B.n227 10.6151
R2655 B.n333 B.n332 10.6151
R2656 B.n332 B.n331 10.6151
R2657 B.n331 B.n229 10.6151
R2658 B.n325 B.n229 10.6151
R2659 B.n325 B.n324 10.6151
R2660 B.n324 B.n323 10.6151
R2661 B.n323 B.n231 10.6151
R2662 B.n317 B.n231 10.6151
R2663 B.n317 B.n316 10.6151
R2664 B.n316 B.n315 10.6151
R2665 B.n315 B.n233 10.6151
R2666 B.n309 B.n233 10.6151
R2667 B.n309 B.n308 10.6151
R2668 B.n308 B.n307 10.6151
R2669 B.n307 B.n235 10.6151
R2670 B.n301 B.n235 10.6151
R2671 B.n301 B.n300 10.6151
R2672 B.n300 B.n299 10.6151
R2673 B.n299 B.n237 10.6151
R2674 B.n293 B.n237 10.6151
R2675 B.n293 B.n292 10.6151
R2676 B.n292 B.n291 10.6151
R2677 B.n291 B.n239 10.6151
R2678 B.n285 B.n239 10.6151
R2679 B.n285 B.n284 10.6151
R2680 B.n284 B.n283 10.6151
R2681 B.n283 B.n241 10.6151
R2682 B.n277 B.n241 10.6151
R2683 B.n277 B.n276 10.6151
R2684 B.n276 B.n275 10.6151
R2685 B.n275 B.n243 10.6151
R2686 B.n269 B.n243 10.6151
R2687 B.n269 B.n268 10.6151
R2688 B.n268 B.n267 10.6151
R2689 B.n267 B.n245 10.6151
R2690 B.n261 B.n245 10.6151
R2691 B.n261 B.n260 10.6151
R2692 B.n260 B.n259 10.6151
R2693 B.n259 B.n247 10.6151
R2694 B.n253 B.n247 10.6151
R2695 B.n253 B.n252 10.6151
R2696 B.n252 B.n251 10.6151
R2697 B.n251 B.n180 10.6151
R2698 B.n491 B.n176 10.6151
R2699 B.n501 B.n176 10.6151
R2700 B.n502 B.n501 10.6151
R2701 B.n503 B.n502 10.6151
R2702 B.n503 B.n168 10.6151
R2703 B.n513 B.n168 10.6151
R2704 B.n514 B.n513 10.6151
R2705 B.n515 B.n514 10.6151
R2706 B.n515 B.n160 10.6151
R2707 B.n525 B.n160 10.6151
R2708 B.n526 B.n525 10.6151
R2709 B.n527 B.n526 10.6151
R2710 B.n527 B.n152 10.6151
R2711 B.n537 B.n152 10.6151
R2712 B.n538 B.n537 10.6151
R2713 B.n539 B.n538 10.6151
R2714 B.n539 B.n144 10.6151
R2715 B.n549 B.n144 10.6151
R2716 B.n550 B.n549 10.6151
R2717 B.n551 B.n550 10.6151
R2718 B.n551 B.n136 10.6151
R2719 B.n561 B.n136 10.6151
R2720 B.n562 B.n561 10.6151
R2721 B.n563 B.n562 10.6151
R2722 B.n563 B.n128 10.6151
R2723 B.n574 B.n128 10.6151
R2724 B.n575 B.n574 10.6151
R2725 B.n576 B.n575 10.6151
R2726 B.n576 B.n0 10.6151
R2727 B.n921 B.n1 10.6151
R2728 B.n921 B.n920 10.6151
R2729 B.n920 B.n919 10.6151
R2730 B.n919 B.n10 10.6151
R2731 B.n913 B.n10 10.6151
R2732 B.n913 B.n912 10.6151
R2733 B.n912 B.n911 10.6151
R2734 B.n911 B.n17 10.6151
R2735 B.n905 B.n17 10.6151
R2736 B.n905 B.n904 10.6151
R2737 B.n904 B.n903 10.6151
R2738 B.n903 B.n24 10.6151
R2739 B.n897 B.n24 10.6151
R2740 B.n897 B.n896 10.6151
R2741 B.n896 B.n895 10.6151
R2742 B.n895 B.n31 10.6151
R2743 B.n889 B.n31 10.6151
R2744 B.n889 B.n888 10.6151
R2745 B.n888 B.n887 10.6151
R2746 B.n887 B.n38 10.6151
R2747 B.n881 B.n38 10.6151
R2748 B.n881 B.n880 10.6151
R2749 B.n880 B.n879 10.6151
R2750 B.n879 B.n45 10.6151
R2751 B.n873 B.n45 10.6151
R2752 B.n873 B.n872 10.6151
R2753 B.n872 B.n871 10.6151
R2754 B.n871 B.n52 10.6151
R2755 B.n865 B.n52 10.6151
R2756 B.n753 B.n752 9.36635
R2757 B.n730 B.n95 9.36635
R2758 B.n381 B.n380 9.36635
R2759 B.n357 B.n222 9.36635
R2760 B.n572 B.t6 7.4179
R2761 B.n917 B.t7 7.4179
R2762 B.n158 B.t4 5.43992
R2763 B.t2 B.n892 5.43992
R2764 B.n559 B.t3 4.45094
R2765 B.n909 B.t5 4.45094
R2766 B.n927 B.n0 2.81026
R2767 B.n927 B.n1 2.81026
R2768 B.n752 B.n751 1.24928
R2769 B.n734 B.n95 1.24928
R2770 B.n380 B.n379 1.24928
R2771 B.n222 B.n218 1.24928
R2772 VP.n7 VP.t0 413.253
R2773 VP.n17 VP.t3 390.002
R2774 VP.n29 VP.t4 390.002
R2775 VP.n15 VP.t1 390.002
R2776 VP.n22 VP.t5 355.632
R2777 VP.n1 VP.t7 355.632
R2778 VP.n5 VP.t6 355.632
R2779 VP.n8 VP.t2 355.632
R2780 VP.n9 VP.n6 161.3
R2781 VP.n11 VP.n10 161.3
R2782 VP.n13 VP.n12 161.3
R2783 VP.n14 VP.n4 161.3
R2784 VP.n28 VP.n0 161.3
R2785 VP.n27 VP.n26 161.3
R2786 VP.n25 VP.n24 161.3
R2787 VP.n23 VP.n2 161.3
R2788 VP.n21 VP.n20 161.3
R2789 VP.n19 VP.n3 161.3
R2790 VP.n16 VP.n15 80.6037
R2791 VP.n30 VP.n29 80.6037
R2792 VP.n18 VP.n17 80.6037
R2793 VP.n24 VP.n23 56.5193
R2794 VP.n10 VP.n9 56.5193
R2795 VP.n17 VP.n3 51.3812
R2796 VP.n29 VP.n28 51.3812
R2797 VP.n15 VP.n14 51.3812
R2798 VP.n18 VP.n16 48.1074
R2799 VP.n8 VP.n7 33.3566
R2800 VP.n7 VP.n6 28.0267
R2801 VP.n21 VP.n3 24.4675
R2802 VP.n28 VP.n27 24.4675
R2803 VP.n14 VP.n13 24.4675
R2804 VP.n23 VP.n22 23.9782
R2805 VP.n24 VP.n1 23.9782
R2806 VP.n10 VP.n5 23.9782
R2807 VP.n9 VP.n8 23.9782
R2808 VP.n22 VP.n21 0.48984
R2809 VP.n27 VP.n1 0.48984
R2810 VP.n13 VP.n5 0.48984
R2811 VP.n16 VP.n4 0.285035
R2812 VP.n19 VP.n18 0.285035
R2813 VP.n30 VP.n0 0.285035
R2814 VP.n11 VP.n6 0.189894
R2815 VP.n12 VP.n11 0.189894
R2816 VP.n12 VP.n4 0.189894
R2817 VP.n20 VP.n19 0.189894
R2818 VP.n20 VP.n2 0.189894
R2819 VP.n25 VP.n2 0.189894
R2820 VP.n26 VP.n25 0.189894
R2821 VP.n26 VP.n0 0.189894
R2822 VP VP.n30 0.146778
R2823 VDD1 VDD1.n0 64.7179
R2824 VDD1.n3 VDD1.n2 64.6042
R2825 VDD1.n3 VDD1.n1 64.6042
R2826 VDD1.n5 VDD1.n4 64.0216
R2827 VDD1.n5 VDD1.n3 44.669
R2828 VDD1.n4 VDD1.t1 1.16726
R2829 VDD1.n4 VDD1.t6 1.16726
R2830 VDD1.n0 VDD1.t7 1.16726
R2831 VDD1.n0 VDD1.t5 1.16726
R2832 VDD1.n2 VDD1.t0 1.16726
R2833 VDD1.n2 VDD1.t3 1.16726
R2834 VDD1.n1 VDD1.t4 1.16726
R2835 VDD1.n1 VDD1.t2 1.16726
R2836 VDD1 VDD1.n5 0.580241
C0 VDD2 VP 0.365433f
C1 VDD1 VDD2 1.05175f
C2 VN VTAIL 9.30977f
C3 VTAIL VP 9.32387f
C4 VDD1 VTAIL 11.8305f
C5 VN VP 6.80607f
C6 VDD2 VTAIL 11.8752f
C7 VDD1 VN 0.149164f
C8 VDD2 VN 9.57499f
C9 VDD1 VP 9.790589f
C10 VDD2 B 4.309605f
C11 VDD1 B 4.589297f
C12 VTAIL B 12.222091f
C13 VN B 10.66166f
C14 VP B 8.739177f
C15 VDD1.t7 B 0.344633f
C16 VDD1.t5 B 0.344633f
C17 VDD1.n0 B 3.1399f
C18 VDD1.t4 B 0.344633f
C19 VDD1.t2 B 0.344633f
C20 VDD1.n1 B 3.13915f
C21 VDD1.t0 B 0.344633f
C22 VDD1.t3 B 0.344633f
C23 VDD1.n2 B 3.13915f
C24 VDD1.n3 B 2.87032f
C25 VDD1.t1 B 0.344633f
C26 VDD1.t6 B 0.344633f
C27 VDD1.n4 B 3.13577f
C28 VDD1.n5 B 2.93462f
C29 VP.n0 B 0.047152f
C30 VP.t7 B 1.89465f
C31 VP.n1 B 0.676717f
C32 VP.n2 B 0.035336f
C33 VP.t5 B 1.89465f
C34 VP.n3 B 0.048277f
C35 VP.n4 B 0.047152f
C36 VP.t1 B 1.9569f
C37 VP.t6 B 1.89465f
C38 VP.n5 B 0.676717f
C39 VP.n6 B 0.187744f
C40 VP.t2 B 1.89465f
C41 VP.t0 B 1.99912f
C42 VP.n7 B 0.723936f
C43 VP.n8 B 0.735696f
C44 VP.n9 B 0.050935f
C45 VP.n10 B 0.050935f
C46 VP.n11 B 0.035336f
C47 VP.n12 B 0.035336f
C48 VP.n13 B 0.033994f
C49 VP.n14 B 0.048277f
C50 VP.n15 B 0.741068f
C51 VP.n16 B 1.82436f
C52 VP.t3 B 1.9569f
C53 VP.n17 B 0.741068f
C54 VP.n18 B 1.85076f
C55 VP.n19 B 0.047152f
C56 VP.n20 B 0.035336f
C57 VP.n21 B 0.033994f
C58 VP.n22 B 0.676717f
C59 VP.n23 B 0.050935f
C60 VP.n24 B 0.050935f
C61 VP.n25 B 0.035336f
C62 VP.n26 B 0.035336f
C63 VP.n27 B 0.033994f
C64 VP.n28 B 0.048277f
C65 VP.t4 B 1.9569f
C66 VP.n29 B 0.741068f
C67 VP.n30 B 0.033094f
C68 VTAIL.t12 B 0.249181f
C69 VTAIL.t13 B 0.249181f
C70 VTAIL.n0 B 2.21531f
C71 VTAIL.n1 B 0.257586f
C72 VTAIL.n2 B 0.027246f
C73 VTAIL.n3 B 0.018581f
C74 VTAIL.n4 B 0.009985f
C75 VTAIL.n5 B 0.023601f
C76 VTAIL.n6 B 0.010572f
C77 VTAIL.n7 B 0.018581f
C78 VTAIL.n8 B 0.009985f
C79 VTAIL.n9 B 0.023601f
C80 VTAIL.n10 B 0.010572f
C81 VTAIL.n11 B 0.018581f
C82 VTAIL.n12 B 0.009985f
C83 VTAIL.n13 B 0.023601f
C84 VTAIL.n14 B 0.010572f
C85 VTAIL.n15 B 0.018581f
C86 VTAIL.n16 B 0.009985f
C87 VTAIL.n17 B 0.023601f
C88 VTAIL.n18 B 0.010572f
C89 VTAIL.n19 B 0.018581f
C90 VTAIL.n20 B 0.009985f
C91 VTAIL.n21 B 0.023601f
C92 VTAIL.n22 B 0.010572f
C93 VTAIL.n23 B 0.018581f
C94 VTAIL.n24 B 0.009985f
C95 VTAIL.n25 B 0.023601f
C96 VTAIL.n26 B 0.010572f
C97 VTAIL.n27 B 0.018581f
C98 VTAIL.n28 B 0.009985f
C99 VTAIL.n29 B 0.023601f
C100 VTAIL.n30 B 0.010572f
C101 VTAIL.n31 B 0.13037f
C102 VTAIL.t14 B 0.03904f
C103 VTAIL.n32 B 0.017701f
C104 VTAIL.n33 B 0.013942f
C105 VTAIL.n34 B 0.009985f
C106 VTAIL.n35 B 1.3767f
C107 VTAIL.n36 B 0.018581f
C108 VTAIL.n37 B 0.009985f
C109 VTAIL.n38 B 0.010572f
C110 VTAIL.n39 B 0.023601f
C111 VTAIL.n40 B 0.023601f
C112 VTAIL.n41 B 0.010572f
C113 VTAIL.n42 B 0.009985f
C114 VTAIL.n43 B 0.018581f
C115 VTAIL.n44 B 0.018581f
C116 VTAIL.n45 B 0.009985f
C117 VTAIL.n46 B 0.010572f
C118 VTAIL.n47 B 0.023601f
C119 VTAIL.n48 B 0.023601f
C120 VTAIL.n49 B 0.010572f
C121 VTAIL.n50 B 0.009985f
C122 VTAIL.n51 B 0.018581f
C123 VTAIL.n52 B 0.018581f
C124 VTAIL.n53 B 0.009985f
C125 VTAIL.n54 B 0.010572f
C126 VTAIL.n55 B 0.023601f
C127 VTAIL.n56 B 0.023601f
C128 VTAIL.n57 B 0.010572f
C129 VTAIL.n58 B 0.009985f
C130 VTAIL.n59 B 0.018581f
C131 VTAIL.n60 B 0.018581f
C132 VTAIL.n61 B 0.009985f
C133 VTAIL.n62 B 0.010572f
C134 VTAIL.n63 B 0.023601f
C135 VTAIL.n64 B 0.023601f
C136 VTAIL.n65 B 0.010572f
C137 VTAIL.n66 B 0.009985f
C138 VTAIL.n67 B 0.018581f
C139 VTAIL.n68 B 0.018581f
C140 VTAIL.n69 B 0.009985f
C141 VTAIL.n70 B 0.010572f
C142 VTAIL.n71 B 0.023601f
C143 VTAIL.n72 B 0.023601f
C144 VTAIL.n73 B 0.023601f
C145 VTAIL.n74 B 0.010572f
C146 VTAIL.n75 B 0.009985f
C147 VTAIL.n76 B 0.018581f
C148 VTAIL.n77 B 0.018581f
C149 VTAIL.n78 B 0.009985f
C150 VTAIL.n79 B 0.010278f
C151 VTAIL.n80 B 0.010278f
C152 VTAIL.n81 B 0.023601f
C153 VTAIL.n82 B 0.023601f
C154 VTAIL.n83 B 0.010572f
C155 VTAIL.n84 B 0.009985f
C156 VTAIL.n85 B 0.018581f
C157 VTAIL.n86 B 0.018581f
C158 VTAIL.n87 B 0.009985f
C159 VTAIL.n88 B 0.010572f
C160 VTAIL.n89 B 0.023601f
C161 VTAIL.n90 B 0.053087f
C162 VTAIL.n91 B 0.010572f
C163 VTAIL.n92 B 0.009985f
C164 VTAIL.n93 B 0.047265f
C165 VTAIL.n94 B 0.030036f
C166 VTAIL.n95 B 0.122832f
C167 VTAIL.n96 B 0.027246f
C168 VTAIL.n97 B 0.018581f
C169 VTAIL.n98 B 0.009985f
C170 VTAIL.n99 B 0.023601f
C171 VTAIL.n100 B 0.010572f
C172 VTAIL.n101 B 0.018581f
C173 VTAIL.n102 B 0.009985f
C174 VTAIL.n103 B 0.023601f
C175 VTAIL.n104 B 0.010572f
C176 VTAIL.n105 B 0.018581f
C177 VTAIL.n106 B 0.009985f
C178 VTAIL.n107 B 0.023601f
C179 VTAIL.n108 B 0.010572f
C180 VTAIL.n109 B 0.018581f
C181 VTAIL.n110 B 0.009985f
C182 VTAIL.n111 B 0.023601f
C183 VTAIL.n112 B 0.010572f
C184 VTAIL.n113 B 0.018581f
C185 VTAIL.n114 B 0.009985f
C186 VTAIL.n115 B 0.023601f
C187 VTAIL.n116 B 0.010572f
C188 VTAIL.n117 B 0.018581f
C189 VTAIL.n118 B 0.009985f
C190 VTAIL.n119 B 0.023601f
C191 VTAIL.n120 B 0.010572f
C192 VTAIL.n121 B 0.018581f
C193 VTAIL.n122 B 0.009985f
C194 VTAIL.n123 B 0.023601f
C195 VTAIL.n124 B 0.010572f
C196 VTAIL.n125 B 0.13037f
C197 VTAIL.t6 B 0.03904f
C198 VTAIL.n126 B 0.017701f
C199 VTAIL.n127 B 0.013942f
C200 VTAIL.n128 B 0.009985f
C201 VTAIL.n129 B 1.3767f
C202 VTAIL.n130 B 0.018581f
C203 VTAIL.n131 B 0.009985f
C204 VTAIL.n132 B 0.010572f
C205 VTAIL.n133 B 0.023601f
C206 VTAIL.n134 B 0.023601f
C207 VTAIL.n135 B 0.010572f
C208 VTAIL.n136 B 0.009985f
C209 VTAIL.n137 B 0.018581f
C210 VTAIL.n138 B 0.018581f
C211 VTAIL.n139 B 0.009985f
C212 VTAIL.n140 B 0.010572f
C213 VTAIL.n141 B 0.023601f
C214 VTAIL.n142 B 0.023601f
C215 VTAIL.n143 B 0.010572f
C216 VTAIL.n144 B 0.009985f
C217 VTAIL.n145 B 0.018581f
C218 VTAIL.n146 B 0.018581f
C219 VTAIL.n147 B 0.009985f
C220 VTAIL.n148 B 0.010572f
C221 VTAIL.n149 B 0.023601f
C222 VTAIL.n150 B 0.023601f
C223 VTAIL.n151 B 0.010572f
C224 VTAIL.n152 B 0.009985f
C225 VTAIL.n153 B 0.018581f
C226 VTAIL.n154 B 0.018581f
C227 VTAIL.n155 B 0.009985f
C228 VTAIL.n156 B 0.010572f
C229 VTAIL.n157 B 0.023601f
C230 VTAIL.n158 B 0.023601f
C231 VTAIL.n159 B 0.010572f
C232 VTAIL.n160 B 0.009985f
C233 VTAIL.n161 B 0.018581f
C234 VTAIL.n162 B 0.018581f
C235 VTAIL.n163 B 0.009985f
C236 VTAIL.n164 B 0.010572f
C237 VTAIL.n165 B 0.023601f
C238 VTAIL.n166 B 0.023601f
C239 VTAIL.n167 B 0.023601f
C240 VTAIL.n168 B 0.010572f
C241 VTAIL.n169 B 0.009985f
C242 VTAIL.n170 B 0.018581f
C243 VTAIL.n171 B 0.018581f
C244 VTAIL.n172 B 0.009985f
C245 VTAIL.n173 B 0.010278f
C246 VTAIL.n174 B 0.010278f
C247 VTAIL.n175 B 0.023601f
C248 VTAIL.n176 B 0.023601f
C249 VTAIL.n177 B 0.010572f
C250 VTAIL.n178 B 0.009985f
C251 VTAIL.n179 B 0.018581f
C252 VTAIL.n180 B 0.018581f
C253 VTAIL.n181 B 0.009985f
C254 VTAIL.n182 B 0.010572f
C255 VTAIL.n183 B 0.023601f
C256 VTAIL.n184 B 0.053087f
C257 VTAIL.n185 B 0.010572f
C258 VTAIL.n186 B 0.009985f
C259 VTAIL.n187 B 0.047265f
C260 VTAIL.n188 B 0.030036f
C261 VTAIL.n189 B 0.122832f
C262 VTAIL.t0 B 0.249181f
C263 VTAIL.t3 B 0.249181f
C264 VTAIL.n190 B 2.21531f
C265 VTAIL.n191 B 0.330492f
C266 VTAIL.n192 B 0.027246f
C267 VTAIL.n193 B 0.018581f
C268 VTAIL.n194 B 0.009985f
C269 VTAIL.n195 B 0.023601f
C270 VTAIL.n196 B 0.010572f
C271 VTAIL.n197 B 0.018581f
C272 VTAIL.n198 B 0.009985f
C273 VTAIL.n199 B 0.023601f
C274 VTAIL.n200 B 0.010572f
C275 VTAIL.n201 B 0.018581f
C276 VTAIL.n202 B 0.009985f
C277 VTAIL.n203 B 0.023601f
C278 VTAIL.n204 B 0.010572f
C279 VTAIL.n205 B 0.018581f
C280 VTAIL.n206 B 0.009985f
C281 VTAIL.n207 B 0.023601f
C282 VTAIL.n208 B 0.010572f
C283 VTAIL.n209 B 0.018581f
C284 VTAIL.n210 B 0.009985f
C285 VTAIL.n211 B 0.023601f
C286 VTAIL.n212 B 0.010572f
C287 VTAIL.n213 B 0.018581f
C288 VTAIL.n214 B 0.009985f
C289 VTAIL.n215 B 0.023601f
C290 VTAIL.n216 B 0.010572f
C291 VTAIL.n217 B 0.018581f
C292 VTAIL.n218 B 0.009985f
C293 VTAIL.n219 B 0.023601f
C294 VTAIL.n220 B 0.010572f
C295 VTAIL.n221 B 0.13037f
C296 VTAIL.t4 B 0.03904f
C297 VTAIL.n222 B 0.017701f
C298 VTAIL.n223 B 0.013942f
C299 VTAIL.n224 B 0.009985f
C300 VTAIL.n225 B 1.3767f
C301 VTAIL.n226 B 0.018581f
C302 VTAIL.n227 B 0.009985f
C303 VTAIL.n228 B 0.010572f
C304 VTAIL.n229 B 0.023601f
C305 VTAIL.n230 B 0.023601f
C306 VTAIL.n231 B 0.010572f
C307 VTAIL.n232 B 0.009985f
C308 VTAIL.n233 B 0.018581f
C309 VTAIL.n234 B 0.018581f
C310 VTAIL.n235 B 0.009985f
C311 VTAIL.n236 B 0.010572f
C312 VTAIL.n237 B 0.023601f
C313 VTAIL.n238 B 0.023601f
C314 VTAIL.n239 B 0.010572f
C315 VTAIL.n240 B 0.009985f
C316 VTAIL.n241 B 0.018581f
C317 VTAIL.n242 B 0.018581f
C318 VTAIL.n243 B 0.009985f
C319 VTAIL.n244 B 0.010572f
C320 VTAIL.n245 B 0.023601f
C321 VTAIL.n246 B 0.023601f
C322 VTAIL.n247 B 0.010572f
C323 VTAIL.n248 B 0.009985f
C324 VTAIL.n249 B 0.018581f
C325 VTAIL.n250 B 0.018581f
C326 VTAIL.n251 B 0.009985f
C327 VTAIL.n252 B 0.010572f
C328 VTAIL.n253 B 0.023601f
C329 VTAIL.n254 B 0.023601f
C330 VTAIL.n255 B 0.010572f
C331 VTAIL.n256 B 0.009985f
C332 VTAIL.n257 B 0.018581f
C333 VTAIL.n258 B 0.018581f
C334 VTAIL.n259 B 0.009985f
C335 VTAIL.n260 B 0.010572f
C336 VTAIL.n261 B 0.023601f
C337 VTAIL.n262 B 0.023601f
C338 VTAIL.n263 B 0.023601f
C339 VTAIL.n264 B 0.010572f
C340 VTAIL.n265 B 0.009985f
C341 VTAIL.n266 B 0.018581f
C342 VTAIL.n267 B 0.018581f
C343 VTAIL.n268 B 0.009985f
C344 VTAIL.n269 B 0.010278f
C345 VTAIL.n270 B 0.010278f
C346 VTAIL.n271 B 0.023601f
C347 VTAIL.n272 B 0.023601f
C348 VTAIL.n273 B 0.010572f
C349 VTAIL.n274 B 0.009985f
C350 VTAIL.n275 B 0.018581f
C351 VTAIL.n276 B 0.018581f
C352 VTAIL.n277 B 0.009985f
C353 VTAIL.n278 B 0.010572f
C354 VTAIL.n279 B 0.023601f
C355 VTAIL.n280 B 0.053087f
C356 VTAIL.n281 B 0.010572f
C357 VTAIL.n282 B 0.009985f
C358 VTAIL.n283 B 0.047265f
C359 VTAIL.n284 B 0.030036f
C360 VTAIL.n285 B 1.29941f
C361 VTAIL.n286 B 0.027246f
C362 VTAIL.n287 B 0.018581f
C363 VTAIL.n288 B 0.009985f
C364 VTAIL.n289 B 0.023601f
C365 VTAIL.n290 B 0.010572f
C366 VTAIL.n291 B 0.018581f
C367 VTAIL.n292 B 0.009985f
C368 VTAIL.n293 B 0.023601f
C369 VTAIL.n294 B 0.010572f
C370 VTAIL.n295 B 0.018581f
C371 VTAIL.n296 B 0.009985f
C372 VTAIL.n297 B 0.023601f
C373 VTAIL.n298 B 0.023601f
C374 VTAIL.n299 B 0.010572f
C375 VTAIL.n300 B 0.018581f
C376 VTAIL.n301 B 0.009985f
C377 VTAIL.n302 B 0.023601f
C378 VTAIL.n303 B 0.010572f
C379 VTAIL.n304 B 0.018581f
C380 VTAIL.n305 B 0.009985f
C381 VTAIL.n306 B 0.023601f
C382 VTAIL.n307 B 0.010572f
C383 VTAIL.n308 B 0.018581f
C384 VTAIL.n309 B 0.009985f
C385 VTAIL.n310 B 0.023601f
C386 VTAIL.n311 B 0.010572f
C387 VTAIL.n312 B 0.018581f
C388 VTAIL.n313 B 0.009985f
C389 VTAIL.n314 B 0.023601f
C390 VTAIL.n315 B 0.010572f
C391 VTAIL.n316 B 0.13037f
C392 VTAIL.t8 B 0.03904f
C393 VTAIL.n317 B 0.017701f
C394 VTAIL.n318 B 0.013942f
C395 VTAIL.n319 B 0.009985f
C396 VTAIL.n320 B 1.3767f
C397 VTAIL.n321 B 0.018581f
C398 VTAIL.n322 B 0.009985f
C399 VTAIL.n323 B 0.010572f
C400 VTAIL.n324 B 0.023601f
C401 VTAIL.n325 B 0.023601f
C402 VTAIL.n326 B 0.010572f
C403 VTAIL.n327 B 0.009985f
C404 VTAIL.n328 B 0.018581f
C405 VTAIL.n329 B 0.018581f
C406 VTAIL.n330 B 0.009985f
C407 VTAIL.n331 B 0.010572f
C408 VTAIL.n332 B 0.023601f
C409 VTAIL.n333 B 0.023601f
C410 VTAIL.n334 B 0.010572f
C411 VTAIL.n335 B 0.009985f
C412 VTAIL.n336 B 0.018581f
C413 VTAIL.n337 B 0.018581f
C414 VTAIL.n338 B 0.009985f
C415 VTAIL.n339 B 0.010572f
C416 VTAIL.n340 B 0.023601f
C417 VTAIL.n341 B 0.023601f
C418 VTAIL.n342 B 0.010572f
C419 VTAIL.n343 B 0.009985f
C420 VTAIL.n344 B 0.018581f
C421 VTAIL.n345 B 0.018581f
C422 VTAIL.n346 B 0.009985f
C423 VTAIL.n347 B 0.010572f
C424 VTAIL.n348 B 0.023601f
C425 VTAIL.n349 B 0.023601f
C426 VTAIL.n350 B 0.010572f
C427 VTAIL.n351 B 0.009985f
C428 VTAIL.n352 B 0.018581f
C429 VTAIL.n353 B 0.018581f
C430 VTAIL.n354 B 0.009985f
C431 VTAIL.n355 B 0.010572f
C432 VTAIL.n356 B 0.023601f
C433 VTAIL.n357 B 0.023601f
C434 VTAIL.n358 B 0.010572f
C435 VTAIL.n359 B 0.009985f
C436 VTAIL.n360 B 0.018581f
C437 VTAIL.n361 B 0.018581f
C438 VTAIL.n362 B 0.009985f
C439 VTAIL.n363 B 0.010278f
C440 VTAIL.n364 B 0.010278f
C441 VTAIL.n365 B 0.023601f
C442 VTAIL.n366 B 0.023601f
C443 VTAIL.n367 B 0.010572f
C444 VTAIL.n368 B 0.009985f
C445 VTAIL.n369 B 0.018581f
C446 VTAIL.n370 B 0.018581f
C447 VTAIL.n371 B 0.009985f
C448 VTAIL.n372 B 0.010572f
C449 VTAIL.n373 B 0.023601f
C450 VTAIL.n374 B 0.053087f
C451 VTAIL.n375 B 0.010572f
C452 VTAIL.n376 B 0.009985f
C453 VTAIL.n377 B 0.047265f
C454 VTAIL.n378 B 0.030036f
C455 VTAIL.n379 B 1.29941f
C456 VTAIL.t10 B 0.249181f
C457 VTAIL.t15 B 0.249181f
C458 VTAIL.n380 B 2.21532f
C459 VTAIL.n381 B 0.330483f
C460 VTAIL.n382 B 0.027246f
C461 VTAIL.n383 B 0.018581f
C462 VTAIL.n384 B 0.009985f
C463 VTAIL.n385 B 0.023601f
C464 VTAIL.n386 B 0.010572f
C465 VTAIL.n387 B 0.018581f
C466 VTAIL.n388 B 0.009985f
C467 VTAIL.n389 B 0.023601f
C468 VTAIL.n390 B 0.010572f
C469 VTAIL.n391 B 0.018581f
C470 VTAIL.n392 B 0.009985f
C471 VTAIL.n393 B 0.023601f
C472 VTAIL.n394 B 0.023601f
C473 VTAIL.n395 B 0.010572f
C474 VTAIL.n396 B 0.018581f
C475 VTAIL.n397 B 0.009985f
C476 VTAIL.n398 B 0.023601f
C477 VTAIL.n399 B 0.010572f
C478 VTAIL.n400 B 0.018581f
C479 VTAIL.n401 B 0.009985f
C480 VTAIL.n402 B 0.023601f
C481 VTAIL.n403 B 0.010572f
C482 VTAIL.n404 B 0.018581f
C483 VTAIL.n405 B 0.009985f
C484 VTAIL.n406 B 0.023601f
C485 VTAIL.n407 B 0.010572f
C486 VTAIL.n408 B 0.018581f
C487 VTAIL.n409 B 0.009985f
C488 VTAIL.n410 B 0.023601f
C489 VTAIL.n411 B 0.010572f
C490 VTAIL.n412 B 0.13037f
C491 VTAIL.t9 B 0.03904f
C492 VTAIL.n413 B 0.017701f
C493 VTAIL.n414 B 0.013942f
C494 VTAIL.n415 B 0.009985f
C495 VTAIL.n416 B 1.3767f
C496 VTAIL.n417 B 0.018581f
C497 VTAIL.n418 B 0.009985f
C498 VTAIL.n419 B 0.010572f
C499 VTAIL.n420 B 0.023601f
C500 VTAIL.n421 B 0.023601f
C501 VTAIL.n422 B 0.010572f
C502 VTAIL.n423 B 0.009985f
C503 VTAIL.n424 B 0.018581f
C504 VTAIL.n425 B 0.018581f
C505 VTAIL.n426 B 0.009985f
C506 VTAIL.n427 B 0.010572f
C507 VTAIL.n428 B 0.023601f
C508 VTAIL.n429 B 0.023601f
C509 VTAIL.n430 B 0.010572f
C510 VTAIL.n431 B 0.009985f
C511 VTAIL.n432 B 0.018581f
C512 VTAIL.n433 B 0.018581f
C513 VTAIL.n434 B 0.009985f
C514 VTAIL.n435 B 0.010572f
C515 VTAIL.n436 B 0.023601f
C516 VTAIL.n437 B 0.023601f
C517 VTAIL.n438 B 0.010572f
C518 VTAIL.n439 B 0.009985f
C519 VTAIL.n440 B 0.018581f
C520 VTAIL.n441 B 0.018581f
C521 VTAIL.n442 B 0.009985f
C522 VTAIL.n443 B 0.010572f
C523 VTAIL.n444 B 0.023601f
C524 VTAIL.n445 B 0.023601f
C525 VTAIL.n446 B 0.010572f
C526 VTAIL.n447 B 0.009985f
C527 VTAIL.n448 B 0.018581f
C528 VTAIL.n449 B 0.018581f
C529 VTAIL.n450 B 0.009985f
C530 VTAIL.n451 B 0.010572f
C531 VTAIL.n452 B 0.023601f
C532 VTAIL.n453 B 0.023601f
C533 VTAIL.n454 B 0.010572f
C534 VTAIL.n455 B 0.009985f
C535 VTAIL.n456 B 0.018581f
C536 VTAIL.n457 B 0.018581f
C537 VTAIL.n458 B 0.009985f
C538 VTAIL.n459 B 0.010278f
C539 VTAIL.n460 B 0.010278f
C540 VTAIL.n461 B 0.023601f
C541 VTAIL.n462 B 0.023601f
C542 VTAIL.n463 B 0.010572f
C543 VTAIL.n464 B 0.009985f
C544 VTAIL.n465 B 0.018581f
C545 VTAIL.n466 B 0.018581f
C546 VTAIL.n467 B 0.009985f
C547 VTAIL.n468 B 0.010572f
C548 VTAIL.n469 B 0.023601f
C549 VTAIL.n470 B 0.053087f
C550 VTAIL.n471 B 0.010572f
C551 VTAIL.n472 B 0.009985f
C552 VTAIL.n473 B 0.047265f
C553 VTAIL.n474 B 0.030036f
C554 VTAIL.n475 B 0.122832f
C555 VTAIL.n476 B 0.027246f
C556 VTAIL.n477 B 0.018581f
C557 VTAIL.n478 B 0.009985f
C558 VTAIL.n479 B 0.023601f
C559 VTAIL.n480 B 0.010572f
C560 VTAIL.n481 B 0.018581f
C561 VTAIL.n482 B 0.009985f
C562 VTAIL.n483 B 0.023601f
C563 VTAIL.n484 B 0.010572f
C564 VTAIL.n485 B 0.018581f
C565 VTAIL.n486 B 0.009985f
C566 VTAIL.n487 B 0.023601f
C567 VTAIL.n488 B 0.023601f
C568 VTAIL.n489 B 0.010572f
C569 VTAIL.n490 B 0.018581f
C570 VTAIL.n491 B 0.009985f
C571 VTAIL.n492 B 0.023601f
C572 VTAIL.n493 B 0.010572f
C573 VTAIL.n494 B 0.018581f
C574 VTAIL.n495 B 0.009985f
C575 VTAIL.n496 B 0.023601f
C576 VTAIL.n497 B 0.010572f
C577 VTAIL.n498 B 0.018581f
C578 VTAIL.n499 B 0.009985f
C579 VTAIL.n500 B 0.023601f
C580 VTAIL.n501 B 0.010572f
C581 VTAIL.n502 B 0.018581f
C582 VTAIL.n503 B 0.009985f
C583 VTAIL.n504 B 0.023601f
C584 VTAIL.n505 B 0.010572f
C585 VTAIL.n506 B 0.13037f
C586 VTAIL.t7 B 0.03904f
C587 VTAIL.n507 B 0.017701f
C588 VTAIL.n508 B 0.013942f
C589 VTAIL.n509 B 0.009985f
C590 VTAIL.n510 B 1.3767f
C591 VTAIL.n511 B 0.018581f
C592 VTAIL.n512 B 0.009985f
C593 VTAIL.n513 B 0.010572f
C594 VTAIL.n514 B 0.023601f
C595 VTAIL.n515 B 0.023601f
C596 VTAIL.n516 B 0.010572f
C597 VTAIL.n517 B 0.009985f
C598 VTAIL.n518 B 0.018581f
C599 VTAIL.n519 B 0.018581f
C600 VTAIL.n520 B 0.009985f
C601 VTAIL.n521 B 0.010572f
C602 VTAIL.n522 B 0.023601f
C603 VTAIL.n523 B 0.023601f
C604 VTAIL.n524 B 0.010572f
C605 VTAIL.n525 B 0.009985f
C606 VTAIL.n526 B 0.018581f
C607 VTAIL.n527 B 0.018581f
C608 VTAIL.n528 B 0.009985f
C609 VTAIL.n529 B 0.010572f
C610 VTAIL.n530 B 0.023601f
C611 VTAIL.n531 B 0.023601f
C612 VTAIL.n532 B 0.010572f
C613 VTAIL.n533 B 0.009985f
C614 VTAIL.n534 B 0.018581f
C615 VTAIL.n535 B 0.018581f
C616 VTAIL.n536 B 0.009985f
C617 VTAIL.n537 B 0.010572f
C618 VTAIL.n538 B 0.023601f
C619 VTAIL.n539 B 0.023601f
C620 VTAIL.n540 B 0.010572f
C621 VTAIL.n541 B 0.009985f
C622 VTAIL.n542 B 0.018581f
C623 VTAIL.n543 B 0.018581f
C624 VTAIL.n544 B 0.009985f
C625 VTAIL.n545 B 0.010572f
C626 VTAIL.n546 B 0.023601f
C627 VTAIL.n547 B 0.023601f
C628 VTAIL.n548 B 0.010572f
C629 VTAIL.n549 B 0.009985f
C630 VTAIL.n550 B 0.018581f
C631 VTAIL.n551 B 0.018581f
C632 VTAIL.n552 B 0.009985f
C633 VTAIL.n553 B 0.010278f
C634 VTAIL.n554 B 0.010278f
C635 VTAIL.n555 B 0.023601f
C636 VTAIL.n556 B 0.023601f
C637 VTAIL.n557 B 0.010572f
C638 VTAIL.n558 B 0.009985f
C639 VTAIL.n559 B 0.018581f
C640 VTAIL.n560 B 0.018581f
C641 VTAIL.n561 B 0.009985f
C642 VTAIL.n562 B 0.010572f
C643 VTAIL.n563 B 0.023601f
C644 VTAIL.n564 B 0.053087f
C645 VTAIL.n565 B 0.010572f
C646 VTAIL.n566 B 0.009985f
C647 VTAIL.n567 B 0.047265f
C648 VTAIL.n568 B 0.030036f
C649 VTAIL.n569 B 0.122832f
C650 VTAIL.t5 B 0.249181f
C651 VTAIL.t1 B 0.249181f
C652 VTAIL.n570 B 2.21532f
C653 VTAIL.n571 B 0.330483f
C654 VTAIL.n572 B 0.027246f
C655 VTAIL.n573 B 0.018581f
C656 VTAIL.n574 B 0.009985f
C657 VTAIL.n575 B 0.023601f
C658 VTAIL.n576 B 0.010572f
C659 VTAIL.n577 B 0.018581f
C660 VTAIL.n578 B 0.009985f
C661 VTAIL.n579 B 0.023601f
C662 VTAIL.n580 B 0.010572f
C663 VTAIL.n581 B 0.018581f
C664 VTAIL.n582 B 0.009985f
C665 VTAIL.n583 B 0.023601f
C666 VTAIL.n584 B 0.023601f
C667 VTAIL.n585 B 0.010572f
C668 VTAIL.n586 B 0.018581f
C669 VTAIL.n587 B 0.009985f
C670 VTAIL.n588 B 0.023601f
C671 VTAIL.n589 B 0.010572f
C672 VTAIL.n590 B 0.018581f
C673 VTAIL.n591 B 0.009985f
C674 VTAIL.n592 B 0.023601f
C675 VTAIL.n593 B 0.010572f
C676 VTAIL.n594 B 0.018581f
C677 VTAIL.n595 B 0.009985f
C678 VTAIL.n596 B 0.023601f
C679 VTAIL.n597 B 0.010572f
C680 VTAIL.n598 B 0.018581f
C681 VTAIL.n599 B 0.009985f
C682 VTAIL.n600 B 0.023601f
C683 VTAIL.n601 B 0.010572f
C684 VTAIL.n602 B 0.13037f
C685 VTAIL.t2 B 0.03904f
C686 VTAIL.n603 B 0.017701f
C687 VTAIL.n604 B 0.013942f
C688 VTAIL.n605 B 0.009985f
C689 VTAIL.n606 B 1.3767f
C690 VTAIL.n607 B 0.018581f
C691 VTAIL.n608 B 0.009985f
C692 VTAIL.n609 B 0.010572f
C693 VTAIL.n610 B 0.023601f
C694 VTAIL.n611 B 0.023601f
C695 VTAIL.n612 B 0.010572f
C696 VTAIL.n613 B 0.009985f
C697 VTAIL.n614 B 0.018581f
C698 VTAIL.n615 B 0.018581f
C699 VTAIL.n616 B 0.009985f
C700 VTAIL.n617 B 0.010572f
C701 VTAIL.n618 B 0.023601f
C702 VTAIL.n619 B 0.023601f
C703 VTAIL.n620 B 0.010572f
C704 VTAIL.n621 B 0.009985f
C705 VTAIL.n622 B 0.018581f
C706 VTAIL.n623 B 0.018581f
C707 VTAIL.n624 B 0.009985f
C708 VTAIL.n625 B 0.010572f
C709 VTAIL.n626 B 0.023601f
C710 VTAIL.n627 B 0.023601f
C711 VTAIL.n628 B 0.010572f
C712 VTAIL.n629 B 0.009985f
C713 VTAIL.n630 B 0.018581f
C714 VTAIL.n631 B 0.018581f
C715 VTAIL.n632 B 0.009985f
C716 VTAIL.n633 B 0.010572f
C717 VTAIL.n634 B 0.023601f
C718 VTAIL.n635 B 0.023601f
C719 VTAIL.n636 B 0.010572f
C720 VTAIL.n637 B 0.009985f
C721 VTAIL.n638 B 0.018581f
C722 VTAIL.n639 B 0.018581f
C723 VTAIL.n640 B 0.009985f
C724 VTAIL.n641 B 0.010572f
C725 VTAIL.n642 B 0.023601f
C726 VTAIL.n643 B 0.023601f
C727 VTAIL.n644 B 0.010572f
C728 VTAIL.n645 B 0.009985f
C729 VTAIL.n646 B 0.018581f
C730 VTAIL.n647 B 0.018581f
C731 VTAIL.n648 B 0.009985f
C732 VTAIL.n649 B 0.010278f
C733 VTAIL.n650 B 0.010278f
C734 VTAIL.n651 B 0.023601f
C735 VTAIL.n652 B 0.023601f
C736 VTAIL.n653 B 0.010572f
C737 VTAIL.n654 B 0.009985f
C738 VTAIL.n655 B 0.018581f
C739 VTAIL.n656 B 0.018581f
C740 VTAIL.n657 B 0.009985f
C741 VTAIL.n658 B 0.010572f
C742 VTAIL.n659 B 0.023601f
C743 VTAIL.n660 B 0.053087f
C744 VTAIL.n661 B 0.010572f
C745 VTAIL.n662 B 0.009985f
C746 VTAIL.n663 B 0.047265f
C747 VTAIL.n664 B 0.030036f
C748 VTAIL.n665 B 1.29941f
C749 VTAIL.n666 B 0.027246f
C750 VTAIL.n667 B 0.018581f
C751 VTAIL.n668 B 0.009985f
C752 VTAIL.n669 B 0.023601f
C753 VTAIL.n670 B 0.010572f
C754 VTAIL.n671 B 0.018581f
C755 VTAIL.n672 B 0.009985f
C756 VTAIL.n673 B 0.023601f
C757 VTAIL.n674 B 0.010572f
C758 VTAIL.n675 B 0.018581f
C759 VTAIL.n676 B 0.009985f
C760 VTAIL.n677 B 0.023601f
C761 VTAIL.n678 B 0.010572f
C762 VTAIL.n679 B 0.018581f
C763 VTAIL.n680 B 0.009985f
C764 VTAIL.n681 B 0.023601f
C765 VTAIL.n682 B 0.010572f
C766 VTAIL.n683 B 0.018581f
C767 VTAIL.n684 B 0.009985f
C768 VTAIL.n685 B 0.023601f
C769 VTAIL.n686 B 0.010572f
C770 VTAIL.n687 B 0.018581f
C771 VTAIL.n688 B 0.009985f
C772 VTAIL.n689 B 0.023601f
C773 VTAIL.n690 B 0.010572f
C774 VTAIL.n691 B 0.018581f
C775 VTAIL.n692 B 0.009985f
C776 VTAIL.n693 B 0.023601f
C777 VTAIL.n694 B 0.010572f
C778 VTAIL.n695 B 0.13037f
C779 VTAIL.t11 B 0.03904f
C780 VTAIL.n696 B 0.017701f
C781 VTAIL.n697 B 0.013942f
C782 VTAIL.n698 B 0.009985f
C783 VTAIL.n699 B 1.3767f
C784 VTAIL.n700 B 0.018581f
C785 VTAIL.n701 B 0.009985f
C786 VTAIL.n702 B 0.010572f
C787 VTAIL.n703 B 0.023601f
C788 VTAIL.n704 B 0.023601f
C789 VTAIL.n705 B 0.010572f
C790 VTAIL.n706 B 0.009985f
C791 VTAIL.n707 B 0.018581f
C792 VTAIL.n708 B 0.018581f
C793 VTAIL.n709 B 0.009985f
C794 VTAIL.n710 B 0.010572f
C795 VTAIL.n711 B 0.023601f
C796 VTAIL.n712 B 0.023601f
C797 VTAIL.n713 B 0.010572f
C798 VTAIL.n714 B 0.009985f
C799 VTAIL.n715 B 0.018581f
C800 VTAIL.n716 B 0.018581f
C801 VTAIL.n717 B 0.009985f
C802 VTAIL.n718 B 0.010572f
C803 VTAIL.n719 B 0.023601f
C804 VTAIL.n720 B 0.023601f
C805 VTAIL.n721 B 0.010572f
C806 VTAIL.n722 B 0.009985f
C807 VTAIL.n723 B 0.018581f
C808 VTAIL.n724 B 0.018581f
C809 VTAIL.n725 B 0.009985f
C810 VTAIL.n726 B 0.010572f
C811 VTAIL.n727 B 0.023601f
C812 VTAIL.n728 B 0.023601f
C813 VTAIL.n729 B 0.010572f
C814 VTAIL.n730 B 0.009985f
C815 VTAIL.n731 B 0.018581f
C816 VTAIL.n732 B 0.018581f
C817 VTAIL.n733 B 0.009985f
C818 VTAIL.n734 B 0.010572f
C819 VTAIL.n735 B 0.023601f
C820 VTAIL.n736 B 0.023601f
C821 VTAIL.n737 B 0.023601f
C822 VTAIL.n738 B 0.010572f
C823 VTAIL.n739 B 0.009985f
C824 VTAIL.n740 B 0.018581f
C825 VTAIL.n741 B 0.018581f
C826 VTAIL.n742 B 0.009985f
C827 VTAIL.n743 B 0.010278f
C828 VTAIL.n744 B 0.010278f
C829 VTAIL.n745 B 0.023601f
C830 VTAIL.n746 B 0.023601f
C831 VTAIL.n747 B 0.010572f
C832 VTAIL.n748 B 0.009985f
C833 VTAIL.n749 B 0.018581f
C834 VTAIL.n750 B 0.018581f
C835 VTAIL.n751 B 0.009985f
C836 VTAIL.n752 B 0.010572f
C837 VTAIL.n753 B 0.023601f
C838 VTAIL.n754 B 0.053087f
C839 VTAIL.n755 B 0.010572f
C840 VTAIL.n756 B 0.009985f
C841 VTAIL.n757 B 0.047265f
C842 VTAIL.n758 B 0.030036f
C843 VTAIL.n759 B 1.29593f
C844 VDD2.t0 B 0.344552f
C845 VDD2.t2 B 0.344552f
C846 VDD2.n0 B 3.1384f
C847 VDD2.t3 B 0.344552f
C848 VDD2.t5 B 0.344552f
C849 VDD2.n1 B 3.1384f
C850 VDD2.n2 B 2.81544f
C851 VDD2.t6 B 0.344552f
C852 VDD2.t4 B 0.344552f
C853 VDD2.n3 B 3.13504f
C854 VDD2.n4 B 2.90285f
C855 VDD2.t1 B 0.344552f
C856 VDD2.t7 B 0.344552f
C857 VDD2.n5 B 3.13838f
C858 VN.n0 B 0.046698f
C859 VN.t2 B 1.87642f
C860 VN.n1 B 0.670206f
C861 VN.n2 B 0.185938f
C862 VN.t3 B 1.87642f
C863 VN.t1 B 1.97988f
C864 VN.n3 B 0.716971f
C865 VN.n4 B 0.728618f
C866 VN.n5 B 0.050445f
C867 VN.n6 B 0.050445f
C868 VN.n7 B 0.034996f
C869 VN.n8 B 0.034996f
C870 VN.n9 B 0.033667f
C871 VN.n10 B 0.047813f
C872 VN.t4 B 1.93807f
C873 VN.n11 B 0.733938f
C874 VN.n12 B 0.032776f
C875 VN.n13 B 0.046698f
C876 VN.t5 B 1.87642f
C877 VN.n14 B 0.670206f
C878 VN.n15 B 0.185938f
C879 VN.t0 B 1.87642f
C880 VN.t6 B 1.97988f
C881 VN.n16 B 0.716971f
C882 VN.n17 B 0.728618f
C883 VN.n18 B 0.050445f
C884 VN.n19 B 0.050445f
C885 VN.n20 B 0.034996f
C886 VN.n21 B 0.034996f
C887 VN.n22 B 0.033667f
C888 VN.n23 B 0.047813f
C889 VN.t7 B 1.93807f
C890 VN.n24 B 0.733938f
C891 VN.n25 B 1.826f
.ends

