* NGSPICE file created from diff_pair_sample_0727.ext - technology: sky130A

.subckt diff_pair_sample_0727 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=0 ps=0 w=8.89 l=0.31
X1 VDD2.t3 VN.t0 VTAIL.t4 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=1.46685 pd=9.22 as=3.4671 ps=18.56 w=8.89 l=0.31
X2 VDD1.t3 VP.t0 VTAIL.t2 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=1.46685 pd=9.22 as=3.4671 ps=18.56 w=8.89 l=0.31
X3 VTAIL.t5 VN.t1 VDD2.t2 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=1.46685 ps=9.22 w=8.89 l=0.31
X4 VTAIL.t6 VN.t2 VDD2.t1 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=1.46685 ps=9.22 w=8.89 l=0.31
X5 B.t8 B.t6 B.t7 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=0 ps=0 w=8.89 l=0.31
X6 VTAIL.t0 VP.t1 VDD1.t2 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=1.46685 ps=9.22 w=8.89 l=0.31
X7 VTAIL.t3 VP.t2 VDD1.t1 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=1.46685 ps=9.22 w=8.89 l=0.31
X8 B.t5 B.t3 B.t4 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=0 ps=0 w=8.89 l=0.31
X9 VDD1.t0 VP.t3 VTAIL.t1 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=1.46685 pd=9.22 as=3.4671 ps=18.56 w=8.89 l=0.31
X10 VDD2.t0 VN.t3 VTAIL.t7 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=1.46685 pd=9.22 as=3.4671 ps=18.56 w=8.89 l=0.31
X11 B.t2 B.t0 B.t1 w_n1354_n2750# sky130_fd_pr__pfet_01v8 ad=3.4671 pd=18.56 as=0 ps=0 w=8.89 l=0.31
R0 B.n86 B.t6 906.097
R1 B.n190 B.t9 906.097
R2 B.n32 B.t0 906.097
R3 B.n26 B.t3 906.097
R4 B.n243 B.n64 585
R5 B.n242 B.n241 585
R6 B.n240 B.n65 585
R7 B.n239 B.n238 585
R8 B.n237 B.n66 585
R9 B.n236 B.n235 585
R10 B.n234 B.n67 585
R11 B.n233 B.n232 585
R12 B.n231 B.n68 585
R13 B.n230 B.n229 585
R14 B.n228 B.n69 585
R15 B.n227 B.n226 585
R16 B.n225 B.n70 585
R17 B.n224 B.n223 585
R18 B.n222 B.n71 585
R19 B.n221 B.n220 585
R20 B.n219 B.n72 585
R21 B.n218 B.n217 585
R22 B.n216 B.n73 585
R23 B.n215 B.n214 585
R24 B.n213 B.n74 585
R25 B.n212 B.n211 585
R26 B.n210 B.n75 585
R27 B.n209 B.n208 585
R28 B.n207 B.n76 585
R29 B.n206 B.n205 585
R30 B.n204 B.n77 585
R31 B.n203 B.n202 585
R32 B.n201 B.n78 585
R33 B.n200 B.n199 585
R34 B.n198 B.n79 585
R35 B.n197 B.n196 585
R36 B.n195 B.n80 585
R37 B.n194 B.n193 585
R38 B.n189 B.n81 585
R39 B.n188 B.n187 585
R40 B.n186 B.n82 585
R41 B.n185 B.n184 585
R42 B.n183 B.n83 585
R43 B.n182 B.n181 585
R44 B.n180 B.n84 585
R45 B.n179 B.n178 585
R46 B.n176 B.n85 585
R47 B.n175 B.n174 585
R48 B.n173 B.n88 585
R49 B.n172 B.n171 585
R50 B.n170 B.n89 585
R51 B.n169 B.n168 585
R52 B.n167 B.n90 585
R53 B.n166 B.n165 585
R54 B.n164 B.n91 585
R55 B.n163 B.n162 585
R56 B.n161 B.n92 585
R57 B.n160 B.n159 585
R58 B.n158 B.n93 585
R59 B.n157 B.n156 585
R60 B.n155 B.n94 585
R61 B.n154 B.n153 585
R62 B.n152 B.n95 585
R63 B.n151 B.n150 585
R64 B.n149 B.n96 585
R65 B.n148 B.n147 585
R66 B.n146 B.n97 585
R67 B.n145 B.n144 585
R68 B.n143 B.n98 585
R69 B.n142 B.n141 585
R70 B.n140 B.n99 585
R71 B.n139 B.n138 585
R72 B.n137 B.n100 585
R73 B.n136 B.n135 585
R74 B.n134 B.n101 585
R75 B.n133 B.n132 585
R76 B.n131 B.n102 585
R77 B.n130 B.n129 585
R78 B.n128 B.n103 585
R79 B.n245 B.n244 585
R80 B.n246 B.n63 585
R81 B.n248 B.n247 585
R82 B.n249 B.n62 585
R83 B.n251 B.n250 585
R84 B.n252 B.n61 585
R85 B.n254 B.n253 585
R86 B.n255 B.n60 585
R87 B.n257 B.n256 585
R88 B.n258 B.n59 585
R89 B.n260 B.n259 585
R90 B.n261 B.n58 585
R91 B.n263 B.n262 585
R92 B.n264 B.n57 585
R93 B.n266 B.n265 585
R94 B.n267 B.n56 585
R95 B.n269 B.n268 585
R96 B.n270 B.n55 585
R97 B.n272 B.n271 585
R98 B.n273 B.n54 585
R99 B.n275 B.n274 585
R100 B.n276 B.n53 585
R101 B.n278 B.n277 585
R102 B.n279 B.n52 585
R103 B.n281 B.n280 585
R104 B.n282 B.n51 585
R105 B.n284 B.n283 585
R106 B.n285 B.n50 585
R107 B.n400 B.n399 585
R108 B.n398 B.n9 585
R109 B.n397 B.n396 585
R110 B.n395 B.n10 585
R111 B.n394 B.n393 585
R112 B.n392 B.n11 585
R113 B.n391 B.n390 585
R114 B.n389 B.n12 585
R115 B.n388 B.n387 585
R116 B.n386 B.n13 585
R117 B.n385 B.n384 585
R118 B.n383 B.n14 585
R119 B.n382 B.n381 585
R120 B.n380 B.n15 585
R121 B.n379 B.n378 585
R122 B.n377 B.n16 585
R123 B.n376 B.n375 585
R124 B.n374 B.n17 585
R125 B.n373 B.n372 585
R126 B.n371 B.n18 585
R127 B.n370 B.n369 585
R128 B.n368 B.n19 585
R129 B.n367 B.n366 585
R130 B.n365 B.n20 585
R131 B.n364 B.n363 585
R132 B.n362 B.n21 585
R133 B.n361 B.n360 585
R134 B.n359 B.n22 585
R135 B.n358 B.n357 585
R136 B.n356 B.n23 585
R137 B.n355 B.n354 585
R138 B.n353 B.n24 585
R139 B.n352 B.n351 585
R140 B.n349 B.n25 585
R141 B.n348 B.n347 585
R142 B.n346 B.n28 585
R143 B.n345 B.n344 585
R144 B.n343 B.n29 585
R145 B.n342 B.n341 585
R146 B.n340 B.n30 585
R147 B.n339 B.n338 585
R148 B.n337 B.n31 585
R149 B.n335 B.n334 585
R150 B.n333 B.n34 585
R151 B.n332 B.n331 585
R152 B.n330 B.n35 585
R153 B.n329 B.n328 585
R154 B.n327 B.n36 585
R155 B.n326 B.n325 585
R156 B.n324 B.n37 585
R157 B.n323 B.n322 585
R158 B.n321 B.n38 585
R159 B.n320 B.n319 585
R160 B.n318 B.n39 585
R161 B.n317 B.n316 585
R162 B.n315 B.n40 585
R163 B.n314 B.n313 585
R164 B.n312 B.n41 585
R165 B.n311 B.n310 585
R166 B.n309 B.n42 585
R167 B.n308 B.n307 585
R168 B.n306 B.n43 585
R169 B.n305 B.n304 585
R170 B.n303 B.n44 585
R171 B.n302 B.n301 585
R172 B.n300 B.n45 585
R173 B.n299 B.n298 585
R174 B.n297 B.n46 585
R175 B.n296 B.n295 585
R176 B.n294 B.n47 585
R177 B.n293 B.n292 585
R178 B.n291 B.n48 585
R179 B.n290 B.n289 585
R180 B.n288 B.n49 585
R181 B.n287 B.n286 585
R182 B.n401 B.n8 585
R183 B.n403 B.n402 585
R184 B.n404 B.n7 585
R185 B.n406 B.n405 585
R186 B.n407 B.n6 585
R187 B.n409 B.n408 585
R188 B.n410 B.n5 585
R189 B.n412 B.n411 585
R190 B.n413 B.n4 585
R191 B.n415 B.n414 585
R192 B.n416 B.n3 585
R193 B.n418 B.n417 585
R194 B.n419 B.n0 585
R195 B.n2 B.n1 585
R196 B.n110 B.n109 585
R197 B.n112 B.n111 585
R198 B.n113 B.n108 585
R199 B.n115 B.n114 585
R200 B.n116 B.n107 585
R201 B.n118 B.n117 585
R202 B.n119 B.n106 585
R203 B.n121 B.n120 585
R204 B.n122 B.n105 585
R205 B.n124 B.n123 585
R206 B.n125 B.n104 585
R207 B.n127 B.n126 585
R208 B.n126 B.n103 511.721
R209 B.n244 B.n243 511.721
R210 B.n286 B.n285 511.721
R211 B.n401 B.n400 511.721
R212 B.n421 B.n420 256.663
R213 B.n420 B.n419 235.042
R214 B.n420 B.n2 235.042
R215 B.n130 B.n103 163.367
R216 B.n131 B.n130 163.367
R217 B.n132 B.n131 163.367
R218 B.n132 B.n101 163.367
R219 B.n136 B.n101 163.367
R220 B.n137 B.n136 163.367
R221 B.n138 B.n137 163.367
R222 B.n138 B.n99 163.367
R223 B.n142 B.n99 163.367
R224 B.n143 B.n142 163.367
R225 B.n144 B.n143 163.367
R226 B.n144 B.n97 163.367
R227 B.n148 B.n97 163.367
R228 B.n149 B.n148 163.367
R229 B.n150 B.n149 163.367
R230 B.n150 B.n95 163.367
R231 B.n154 B.n95 163.367
R232 B.n155 B.n154 163.367
R233 B.n156 B.n155 163.367
R234 B.n156 B.n93 163.367
R235 B.n160 B.n93 163.367
R236 B.n161 B.n160 163.367
R237 B.n162 B.n161 163.367
R238 B.n162 B.n91 163.367
R239 B.n166 B.n91 163.367
R240 B.n167 B.n166 163.367
R241 B.n168 B.n167 163.367
R242 B.n168 B.n89 163.367
R243 B.n172 B.n89 163.367
R244 B.n173 B.n172 163.367
R245 B.n174 B.n173 163.367
R246 B.n174 B.n85 163.367
R247 B.n179 B.n85 163.367
R248 B.n180 B.n179 163.367
R249 B.n181 B.n180 163.367
R250 B.n181 B.n83 163.367
R251 B.n185 B.n83 163.367
R252 B.n186 B.n185 163.367
R253 B.n187 B.n186 163.367
R254 B.n187 B.n81 163.367
R255 B.n194 B.n81 163.367
R256 B.n195 B.n194 163.367
R257 B.n196 B.n195 163.367
R258 B.n196 B.n79 163.367
R259 B.n200 B.n79 163.367
R260 B.n201 B.n200 163.367
R261 B.n202 B.n201 163.367
R262 B.n202 B.n77 163.367
R263 B.n206 B.n77 163.367
R264 B.n207 B.n206 163.367
R265 B.n208 B.n207 163.367
R266 B.n208 B.n75 163.367
R267 B.n212 B.n75 163.367
R268 B.n213 B.n212 163.367
R269 B.n214 B.n213 163.367
R270 B.n214 B.n73 163.367
R271 B.n218 B.n73 163.367
R272 B.n219 B.n218 163.367
R273 B.n220 B.n219 163.367
R274 B.n220 B.n71 163.367
R275 B.n224 B.n71 163.367
R276 B.n225 B.n224 163.367
R277 B.n226 B.n225 163.367
R278 B.n226 B.n69 163.367
R279 B.n230 B.n69 163.367
R280 B.n231 B.n230 163.367
R281 B.n232 B.n231 163.367
R282 B.n232 B.n67 163.367
R283 B.n236 B.n67 163.367
R284 B.n237 B.n236 163.367
R285 B.n238 B.n237 163.367
R286 B.n238 B.n65 163.367
R287 B.n242 B.n65 163.367
R288 B.n243 B.n242 163.367
R289 B.n285 B.n284 163.367
R290 B.n284 B.n51 163.367
R291 B.n280 B.n51 163.367
R292 B.n280 B.n279 163.367
R293 B.n279 B.n278 163.367
R294 B.n278 B.n53 163.367
R295 B.n274 B.n53 163.367
R296 B.n274 B.n273 163.367
R297 B.n273 B.n272 163.367
R298 B.n272 B.n55 163.367
R299 B.n268 B.n55 163.367
R300 B.n268 B.n267 163.367
R301 B.n267 B.n266 163.367
R302 B.n266 B.n57 163.367
R303 B.n262 B.n57 163.367
R304 B.n262 B.n261 163.367
R305 B.n261 B.n260 163.367
R306 B.n260 B.n59 163.367
R307 B.n256 B.n59 163.367
R308 B.n256 B.n255 163.367
R309 B.n255 B.n254 163.367
R310 B.n254 B.n61 163.367
R311 B.n250 B.n61 163.367
R312 B.n250 B.n249 163.367
R313 B.n249 B.n248 163.367
R314 B.n248 B.n63 163.367
R315 B.n244 B.n63 163.367
R316 B.n400 B.n9 163.367
R317 B.n396 B.n9 163.367
R318 B.n396 B.n395 163.367
R319 B.n395 B.n394 163.367
R320 B.n394 B.n11 163.367
R321 B.n390 B.n11 163.367
R322 B.n390 B.n389 163.367
R323 B.n389 B.n388 163.367
R324 B.n388 B.n13 163.367
R325 B.n384 B.n13 163.367
R326 B.n384 B.n383 163.367
R327 B.n383 B.n382 163.367
R328 B.n382 B.n15 163.367
R329 B.n378 B.n15 163.367
R330 B.n378 B.n377 163.367
R331 B.n377 B.n376 163.367
R332 B.n376 B.n17 163.367
R333 B.n372 B.n17 163.367
R334 B.n372 B.n371 163.367
R335 B.n371 B.n370 163.367
R336 B.n370 B.n19 163.367
R337 B.n366 B.n19 163.367
R338 B.n366 B.n365 163.367
R339 B.n365 B.n364 163.367
R340 B.n364 B.n21 163.367
R341 B.n360 B.n21 163.367
R342 B.n360 B.n359 163.367
R343 B.n359 B.n358 163.367
R344 B.n358 B.n23 163.367
R345 B.n354 B.n23 163.367
R346 B.n354 B.n353 163.367
R347 B.n353 B.n352 163.367
R348 B.n352 B.n25 163.367
R349 B.n347 B.n25 163.367
R350 B.n347 B.n346 163.367
R351 B.n346 B.n345 163.367
R352 B.n345 B.n29 163.367
R353 B.n341 B.n29 163.367
R354 B.n341 B.n340 163.367
R355 B.n340 B.n339 163.367
R356 B.n339 B.n31 163.367
R357 B.n334 B.n31 163.367
R358 B.n334 B.n333 163.367
R359 B.n333 B.n332 163.367
R360 B.n332 B.n35 163.367
R361 B.n328 B.n35 163.367
R362 B.n328 B.n327 163.367
R363 B.n327 B.n326 163.367
R364 B.n326 B.n37 163.367
R365 B.n322 B.n37 163.367
R366 B.n322 B.n321 163.367
R367 B.n321 B.n320 163.367
R368 B.n320 B.n39 163.367
R369 B.n316 B.n39 163.367
R370 B.n316 B.n315 163.367
R371 B.n315 B.n314 163.367
R372 B.n314 B.n41 163.367
R373 B.n310 B.n41 163.367
R374 B.n310 B.n309 163.367
R375 B.n309 B.n308 163.367
R376 B.n308 B.n43 163.367
R377 B.n304 B.n43 163.367
R378 B.n304 B.n303 163.367
R379 B.n303 B.n302 163.367
R380 B.n302 B.n45 163.367
R381 B.n298 B.n45 163.367
R382 B.n298 B.n297 163.367
R383 B.n297 B.n296 163.367
R384 B.n296 B.n47 163.367
R385 B.n292 B.n47 163.367
R386 B.n292 B.n291 163.367
R387 B.n291 B.n290 163.367
R388 B.n290 B.n49 163.367
R389 B.n286 B.n49 163.367
R390 B.n402 B.n401 163.367
R391 B.n402 B.n7 163.367
R392 B.n406 B.n7 163.367
R393 B.n407 B.n406 163.367
R394 B.n408 B.n407 163.367
R395 B.n408 B.n5 163.367
R396 B.n412 B.n5 163.367
R397 B.n413 B.n412 163.367
R398 B.n414 B.n413 163.367
R399 B.n414 B.n3 163.367
R400 B.n418 B.n3 163.367
R401 B.n419 B.n418 163.367
R402 B.n109 B.n2 163.367
R403 B.n112 B.n109 163.367
R404 B.n113 B.n112 163.367
R405 B.n114 B.n113 163.367
R406 B.n114 B.n107 163.367
R407 B.n118 B.n107 163.367
R408 B.n119 B.n118 163.367
R409 B.n120 B.n119 163.367
R410 B.n120 B.n105 163.367
R411 B.n124 B.n105 163.367
R412 B.n125 B.n124 163.367
R413 B.n126 B.n125 163.367
R414 B.n190 B.t10 121.52
R415 B.n32 B.t2 121.52
R416 B.n86 B.t7 121.51
R417 B.n26 B.t5 121.51
R418 B.n191 B.t11 109.109
R419 B.n33 B.t1 109.109
R420 B.n87 B.t8 109.099
R421 B.n27 B.t4 109.099
R422 B.n177 B.n87 59.5399
R423 B.n192 B.n191 59.5399
R424 B.n336 B.n33 59.5399
R425 B.n350 B.n27 59.5399
R426 B.n399 B.n8 33.2493
R427 B.n287 B.n50 33.2493
R428 B.n245 B.n64 33.2493
R429 B.n128 B.n127 33.2493
R430 B B.n421 18.0485
R431 B.n87 B.n86 12.4126
R432 B.n191 B.n190 12.4126
R433 B.n33 B.n32 12.4126
R434 B.n27 B.n26 12.4126
R435 B.n403 B.n8 10.6151
R436 B.n404 B.n403 10.6151
R437 B.n405 B.n404 10.6151
R438 B.n405 B.n6 10.6151
R439 B.n409 B.n6 10.6151
R440 B.n410 B.n409 10.6151
R441 B.n411 B.n410 10.6151
R442 B.n411 B.n4 10.6151
R443 B.n415 B.n4 10.6151
R444 B.n416 B.n415 10.6151
R445 B.n417 B.n416 10.6151
R446 B.n417 B.n0 10.6151
R447 B.n399 B.n398 10.6151
R448 B.n398 B.n397 10.6151
R449 B.n397 B.n10 10.6151
R450 B.n393 B.n10 10.6151
R451 B.n393 B.n392 10.6151
R452 B.n392 B.n391 10.6151
R453 B.n391 B.n12 10.6151
R454 B.n387 B.n12 10.6151
R455 B.n387 B.n386 10.6151
R456 B.n386 B.n385 10.6151
R457 B.n385 B.n14 10.6151
R458 B.n381 B.n14 10.6151
R459 B.n381 B.n380 10.6151
R460 B.n380 B.n379 10.6151
R461 B.n379 B.n16 10.6151
R462 B.n375 B.n16 10.6151
R463 B.n375 B.n374 10.6151
R464 B.n374 B.n373 10.6151
R465 B.n373 B.n18 10.6151
R466 B.n369 B.n18 10.6151
R467 B.n369 B.n368 10.6151
R468 B.n368 B.n367 10.6151
R469 B.n367 B.n20 10.6151
R470 B.n363 B.n20 10.6151
R471 B.n363 B.n362 10.6151
R472 B.n362 B.n361 10.6151
R473 B.n361 B.n22 10.6151
R474 B.n357 B.n22 10.6151
R475 B.n357 B.n356 10.6151
R476 B.n356 B.n355 10.6151
R477 B.n355 B.n24 10.6151
R478 B.n351 B.n24 10.6151
R479 B.n349 B.n348 10.6151
R480 B.n348 B.n28 10.6151
R481 B.n344 B.n28 10.6151
R482 B.n344 B.n343 10.6151
R483 B.n343 B.n342 10.6151
R484 B.n342 B.n30 10.6151
R485 B.n338 B.n30 10.6151
R486 B.n338 B.n337 10.6151
R487 B.n335 B.n34 10.6151
R488 B.n331 B.n34 10.6151
R489 B.n331 B.n330 10.6151
R490 B.n330 B.n329 10.6151
R491 B.n329 B.n36 10.6151
R492 B.n325 B.n36 10.6151
R493 B.n325 B.n324 10.6151
R494 B.n324 B.n323 10.6151
R495 B.n323 B.n38 10.6151
R496 B.n319 B.n38 10.6151
R497 B.n319 B.n318 10.6151
R498 B.n318 B.n317 10.6151
R499 B.n317 B.n40 10.6151
R500 B.n313 B.n40 10.6151
R501 B.n313 B.n312 10.6151
R502 B.n312 B.n311 10.6151
R503 B.n311 B.n42 10.6151
R504 B.n307 B.n42 10.6151
R505 B.n307 B.n306 10.6151
R506 B.n306 B.n305 10.6151
R507 B.n305 B.n44 10.6151
R508 B.n301 B.n44 10.6151
R509 B.n301 B.n300 10.6151
R510 B.n300 B.n299 10.6151
R511 B.n299 B.n46 10.6151
R512 B.n295 B.n46 10.6151
R513 B.n295 B.n294 10.6151
R514 B.n294 B.n293 10.6151
R515 B.n293 B.n48 10.6151
R516 B.n289 B.n48 10.6151
R517 B.n289 B.n288 10.6151
R518 B.n288 B.n287 10.6151
R519 B.n283 B.n50 10.6151
R520 B.n283 B.n282 10.6151
R521 B.n282 B.n281 10.6151
R522 B.n281 B.n52 10.6151
R523 B.n277 B.n52 10.6151
R524 B.n277 B.n276 10.6151
R525 B.n276 B.n275 10.6151
R526 B.n275 B.n54 10.6151
R527 B.n271 B.n54 10.6151
R528 B.n271 B.n270 10.6151
R529 B.n270 B.n269 10.6151
R530 B.n269 B.n56 10.6151
R531 B.n265 B.n56 10.6151
R532 B.n265 B.n264 10.6151
R533 B.n264 B.n263 10.6151
R534 B.n263 B.n58 10.6151
R535 B.n259 B.n58 10.6151
R536 B.n259 B.n258 10.6151
R537 B.n258 B.n257 10.6151
R538 B.n257 B.n60 10.6151
R539 B.n253 B.n60 10.6151
R540 B.n253 B.n252 10.6151
R541 B.n252 B.n251 10.6151
R542 B.n251 B.n62 10.6151
R543 B.n247 B.n62 10.6151
R544 B.n247 B.n246 10.6151
R545 B.n246 B.n245 10.6151
R546 B.n110 B.n1 10.6151
R547 B.n111 B.n110 10.6151
R548 B.n111 B.n108 10.6151
R549 B.n115 B.n108 10.6151
R550 B.n116 B.n115 10.6151
R551 B.n117 B.n116 10.6151
R552 B.n117 B.n106 10.6151
R553 B.n121 B.n106 10.6151
R554 B.n122 B.n121 10.6151
R555 B.n123 B.n122 10.6151
R556 B.n123 B.n104 10.6151
R557 B.n127 B.n104 10.6151
R558 B.n129 B.n128 10.6151
R559 B.n129 B.n102 10.6151
R560 B.n133 B.n102 10.6151
R561 B.n134 B.n133 10.6151
R562 B.n135 B.n134 10.6151
R563 B.n135 B.n100 10.6151
R564 B.n139 B.n100 10.6151
R565 B.n140 B.n139 10.6151
R566 B.n141 B.n140 10.6151
R567 B.n141 B.n98 10.6151
R568 B.n145 B.n98 10.6151
R569 B.n146 B.n145 10.6151
R570 B.n147 B.n146 10.6151
R571 B.n147 B.n96 10.6151
R572 B.n151 B.n96 10.6151
R573 B.n152 B.n151 10.6151
R574 B.n153 B.n152 10.6151
R575 B.n153 B.n94 10.6151
R576 B.n157 B.n94 10.6151
R577 B.n158 B.n157 10.6151
R578 B.n159 B.n158 10.6151
R579 B.n159 B.n92 10.6151
R580 B.n163 B.n92 10.6151
R581 B.n164 B.n163 10.6151
R582 B.n165 B.n164 10.6151
R583 B.n165 B.n90 10.6151
R584 B.n169 B.n90 10.6151
R585 B.n170 B.n169 10.6151
R586 B.n171 B.n170 10.6151
R587 B.n171 B.n88 10.6151
R588 B.n175 B.n88 10.6151
R589 B.n176 B.n175 10.6151
R590 B.n178 B.n84 10.6151
R591 B.n182 B.n84 10.6151
R592 B.n183 B.n182 10.6151
R593 B.n184 B.n183 10.6151
R594 B.n184 B.n82 10.6151
R595 B.n188 B.n82 10.6151
R596 B.n189 B.n188 10.6151
R597 B.n193 B.n189 10.6151
R598 B.n197 B.n80 10.6151
R599 B.n198 B.n197 10.6151
R600 B.n199 B.n198 10.6151
R601 B.n199 B.n78 10.6151
R602 B.n203 B.n78 10.6151
R603 B.n204 B.n203 10.6151
R604 B.n205 B.n204 10.6151
R605 B.n205 B.n76 10.6151
R606 B.n209 B.n76 10.6151
R607 B.n210 B.n209 10.6151
R608 B.n211 B.n210 10.6151
R609 B.n211 B.n74 10.6151
R610 B.n215 B.n74 10.6151
R611 B.n216 B.n215 10.6151
R612 B.n217 B.n216 10.6151
R613 B.n217 B.n72 10.6151
R614 B.n221 B.n72 10.6151
R615 B.n222 B.n221 10.6151
R616 B.n223 B.n222 10.6151
R617 B.n223 B.n70 10.6151
R618 B.n227 B.n70 10.6151
R619 B.n228 B.n227 10.6151
R620 B.n229 B.n228 10.6151
R621 B.n229 B.n68 10.6151
R622 B.n233 B.n68 10.6151
R623 B.n234 B.n233 10.6151
R624 B.n235 B.n234 10.6151
R625 B.n235 B.n66 10.6151
R626 B.n239 B.n66 10.6151
R627 B.n240 B.n239 10.6151
R628 B.n241 B.n240 10.6151
R629 B.n241 B.n64 10.6151
R630 B.n421 B.n0 8.11757
R631 B.n421 B.n1 8.11757
R632 B.n350 B.n349 7.18099
R633 B.n337 B.n336 7.18099
R634 B.n178 B.n177 7.18099
R635 B.n193 B.n192 7.18099
R636 B.n351 B.n350 3.43465
R637 B.n336 B.n335 3.43465
R638 B.n177 B.n176 3.43465
R639 B.n192 B.n80 3.43465
R640 VN.n0 VN.t0 839.707
R641 VN.n0 VN.t1 839.707
R642 VN.n1 VN.t2 839.707
R643 VN.n1 VN.t3 839.707
R644 VN VN.n1 198.65
R645 VN VN.n0 161.351
R646 VTAIL.n5 VTAIL.t3 66.577
R647 VTAIL.n4 VTAIL.t7 66.577
R648 VTAIL.n3 VTAIL.t6 66.577
R649 VTAIL.n7 VTAIL.t4 66.5768
R650 VTAIL.n0 VTAIL.t5 66.5768
R651 VTAIL.n1 VTAIL.t1 66.5768
R652 VTAIL.n2 VTAIL.t0 66.5768
R653 VTAIL.n6 VTAIL.t2 66.5768
R654 VTAIL.n7 VTAIL.n6 20.5996
R655 VTAIL.n3 VTAIL.n2 20.5996
R656 VTAIL.n4 VTAIL.n3 0.552224
R657 VTAIL.n6 VTAIL.n5 0.552224
R658 VTAIL.n2 VTAIL.n1 0.552224
R659 VTAIL.n5 VTAIL.n4 0.470328
R660 VTAIL.n1 VTAIL.n0 0.470328
R661 VTAIL VTAIL.n0 0.334552
R662 VTAIL VTAIL.n7 0.218172
R663 VDD2.n2 VDD2.n0 112.65
R664 VDD2.n2 VDD2.n1 79.5993
R665 VDD2.n1 VDD2.t1 3.65686
R666 VDD2.n1 VDD2.t0 3.65686
R667 VDD2.n0 VDD2.t2 3.65686
R668 VDD2.n0 VDD2.t3 3.65686
R669 VDD2 VDD2.n2 0.0586897
R670 VP.n1 VP.t3 839.707
R671 VP.n1 VP.t1 839.707
R672 VP.n0 VP.t2 839.707
R673 VP.n0 VP.t0 839.707
R674 VP.n2 VP.n0 198.27
R675 VP.n2 VP.n1 161.3
R676 VP VP.n2 0.0516364
R677 VDD1 VDD1.n1 113.175
R678 VDD1 VDD1.n0 79.6575
R679 VDD1.n0 VDD1.t1 3.65686
R680 VDD1.n0 VDD1.t3 3.65686
R681 VDD1.n1 VDD1.t2 3.65686
R682 VDD1.n1 VDD1.t0 3.65686
C0 B VDD1 0.773109f
C1 VP VDD2 0.249729f
C2 w_n1354_n2750# VDD1 0.887135f
C3 VDD1 VDD2 0.480601f
C4 VTAIL VP 1.26526f
C5 VTAIL VDD1 7.230721f
C6 VP VDD1 1.73728f
C7 B VN 0.633339f
C8 VN w_n1354_n2750# 1.8126f
C9 VN VDD2 1.63578f
C10 VTAIL VN 1.25115f
C11 VN VP 3.959f
C12 VN VDD1 0.14807f
C13 B w_n1354_n2750# 5.57108f
C14 B VDD2 0.789254f
C15 w_n1354_n2750# VDD2 0.894138f
C16 B VTAIL 2.73666f
C17 VTAIL w_n1354_n2750# 3.42929f
C18 VTAIL VDD2 7.26958f
C19 B VP 0.901918f
C20 VP w_n1354_n2750# 1.98087f
C21 VDD2 VSUBS 0.543207f
C22 VDD1 VSUBS 3.977511f
C23 VTAIL VSUBS 0.628184f
C24 VN VSUBS 3.67202f
C25 VP VSUBS 0.968727f
C26 B VSUBS 2.025085f
C27 w_n1354_n2750# VSUBS 46.0956f
C28 VDD1.t1 VSUBS 0.181541f
C29 VDD1.t3 VSUBS 0.181541f
C30 VDD1.n0 VSUBS 1.33986f
C31 VDD1.t2 VSUBS 0.181541f
C32 VDD1.t0 VSUBS 0.181541f
C33 VDD1.n1 VSUBS 1.805f
C34 VP.t2 VSUBS 0.283034f
C35 VP.t0 VSUBS 0.283034f
C36 VP.n0 VSUBS 0.457868f
C37 VP.t1 VSUBS 0.283034f
C38 VP.t3 VSUBS 0.283034f
C39 VP.n1 VSUBS 0.238144f
C40 VP.n2 VSUBS 2.15407f
C41 VDD2.t2 VSUBS 0.186536f
C42 VDD2.t3 VSUBS 0.186536f
C43 VDD2.n0 VSUBS 1.83339f
C44 VDD2.t1 VSUBS 0.186536f
C45 VDD2.t0 VSUBS 0.186536f
C46 VDD2.n1 VSUBS 1.37633f
C47 VDD2.n2 VSUBS 3.29122f
C48 VTAIL.t5 VSUBS 1.48078f
C49 VTAIL.n0 VSUBS 0.625102f
C50 VTAIL.t1 VSUBS 1.48078f
C51 VTAIL.n1 VSUBS 0.641553f
C52 VTAIL.t0 VSUBS 1.48078f
C53 VTAIL.n2 VSUBS 1.5469f
C54 VTAIL.t6 VSUBS 1.48078f
C55 VTAIL.n3 VSUBS 1.54689f
C56 VTAIL.t7 VSUBS 1.48078f
C57 VTAIL.n4 VSUBS 0.641549f
C58 VTAIL.t3 VSUBS 1.48078f
C59 VTAIL.n5 VSUBS 0.641549f
C60 VTAIL.t2 VSUBS 1.48078f
C61 VTAIL.n6 VSUBS 1.5469f
C62 VTAIL.t4 VSUBS 1.48078f
C63 VTAIL.n7 VSUBS 1.52165f
C64 VN.t1 VSUBS 0.279558f
C65 VN.t0 VSUBS 0.279558f
C66 VN.n0 VSUBS 0.23523f
C67 VN.t2 VSUBS 0.279558f
C68 VN.t3 VSUBS 0.279558f
C69 VN.n1 VSUBS 0.458409f
C70 B.n0 VSUBS 0.008029f
C71 B.n1 VSUBS 0.008029f
C72 B.n2 VSUBS 0.011875f
C73 B.n3 VSUBS 0.0091f
C74 B.n4 VSUBS 0.0091f
C75 B.n5 VSUBS 0.0091f
C76 B.n6 VSUBS 0.0091f
C77 B.n7 VSUBS 0.0091f
C78 B.n8 VSUBS 0.020657f
C79 B.n9 VSUBS 0.0091f
C80 B.n10 VSUBS 0.0091f
C81 B.n11 VSUBS 0.0091f
C82 B.n12 VSUBS 0.0091f
C83 B.n13 VSUBS 0.0091f
C84 B.n14 VSUBS 0.0091f
C85 B.n15 VSUBS 0.0091f
C86 B.n16 VSUBS 0.0091f
C87 B.n17 VSUBS 0.0091f
C88 B.n18 VSUBS 0.0091f
C89 B.n19 VSUBS 0.0091f
C90 B.n20 VSUBS 0.0091f
C91 B.n21 VSUBS 0.0091f
C92 B.n22 VSUBS 0.0091f
C93 B.n23 VSUBS 0.0091f
C94 B.n24 VSUBS 0.0091f
C95 B.n25 VSUBS 0.0091f
C96 B.t4 VSUBS 0.36259f
C97 B.t5 VSUBS 0.369498f
C98 B.t3 VSUBS 0.142868f
C99 B.n26 VSUBS 0.111757f
C100 B.n27 VSUBS 0.08061f
C101 B.n28 VSUBS 0.0091f
C102 B.n29 VSUBS 0.0091f
C103 B.n30 VSUBS 0.0091f
C104 B.n31 VSUBS 0.0091f
C105 B.t1 VSUBS 0.362586f
C106 B.t2 VSUBS 0.369494f
C107 B.t0 VSUBS 0.142868f
C108 B.n32 VSUBS 0.111761f
C109 B.n33 VSUBS 0.080614f
C110 B.n34 VSUBS 0.0091f
C111 B.n35 VSUBS 0.0091f
C112 B.n36 VSUBS 0.0091f
C113 B.n37 VSUBS 0.0091f
C114 B.n38 VSUBS 0.0091f
C115 B.n39 VSUBS 0.0091f
C116 B.n40 VSUBS 0.0091f
C117 B.n41 VSUBS 0.0091f
C118 B.n42 VSUBS 0.0091f
C119 B.n43 VSUBS 0.0091f
C120 B.n44 VSUBS 0.0091f
C121 B.n45 VSUBS 0.0091f
C122 B.n46 VSUBS 0.0091f
C123 B.n47 VSUBS 0.0091f
C124 B.n48 VSUBS 0.0091f
C125 B.n49 VSUBS 0.0091f
C126 B.n50 VSUBS 0.020657f
C127 B.n51 VSUBS 0.0091f
C128 B.n52 VSUBS 0.0091f
C129 B.n53 VSUBS 0.0091f
C130 B.n54 VSUBS 0.0091f
C131 B.n55 VSUBS 0.0091f
C132 B.n56 VSUBS 0.0091f
C133 B.n57 VSUBS 0.0091f
C134 B.n58 VSUBS 0.0091f
C135 B.n59 VSUBS 0.0091f
C136 B.n60 VSUBS 0.0091f
C137 B.n61 VSUBS 0.0091f
C138 B.n62 VSUBS 0.0091f
C139 B.n63 VSUBS 0.0091f
C140 B.n64 VSUBS 0.021378f
C141 B.n65 VSUBS 0.0091f
C142 B.n66 VSUBS 0.0091f
C143 B.n67 VSUBS 0.0091f
C144 B.n68 VSUBS 0.0091f
C145 B.n69 VSUBS 0.0091f
C146 B.n70 VSUBS 0.0091f
C147 B.n71 VSUBS 0.0091f
C148 B.n72 VSUBS 0.0091f
C149 B.n73 VSUBS 0.0091f
C150 B.n74 VSUBS 0.0091f
C151 B.n75 VSUBS 0.0091f
C152 B.n76 VSUBS 0.0091f
C153 B.n77 VSUBS 0.0091f
C154 B.n78 VSUBS 0.0091f
C155 B.n79 VSUBS 0.0091f
C156 B.n80 VSUBS 0.006022f
C157 B.n81 VSUBS 0.0091f
C158 B.n82 VSUBS 0.0091f
C159 B.n83 VSUBS 0.0091f
C160 B.n84 VSUBS 0.0091f
C161 B.n85 VSUBS 0.0091f
C162 B.t8 VSUBS 0.36259f
C163 B.t7 VSUBS 0.369498f
C164 B.t6 VSUBS 0.142868f
C165 B.n86 VSUBS 0.111757f
C166 B.n87 VSUBS 0.08061f
C167 B.n88 VSUBS 0.0091f
C168 B.n89 VSUBS 0.0091f
C169 B.n90 VSUBS 0.0091f
C170 B.n91 VSUBS 0.0091f
C171 B.n92 VSUBS 0.0091f
C172 B.n93 VSUBS 0.0091f
C173 B.n94 VSUBS 0.0091f
C174 B.n95 VSUBS 0.0091f
C175 B.n96 VSUBS 0.0091f
C176 B.n97 VSUBS 0.0091f
C177 B.n98 VSUBS 0.0091f
C178 B.n99 VSUBS 0.0091f
C179 B.n100 VSUBS 0.0091f
C180 B.n101 VSUBS 0.0091f
C181 B.n102 VSUBS 0.0091f
C182 B.n103 VSUBS 0.022434f
C183 B.n104 VSUBS 0.0091f
C184 B.n105 VSUBS 0.0091f
C185 B.n106 VSUBS 0.0091f
C186 B.n107 VSUBS 0.0091f
C187 B.n108 VSUBS 0.0091f
C188 B.n109 VSUBS 0.0091f
C189 B.n110 VSUBS 0.0091f
C190 B.n111 VSUBS 0.0091f
C191 B.n112 VSUBS 0.0091f
C192 B.n113 VSUBS 0.0091f
C193 B.n114 VSUBS 0.0091f
C194 B.n115 VSUBS 0.0091f
C195 B.n116 VSUBS 0.0091f
C196 B.n117 VSUBS 0.0091f
C197 B.n118 VSUBS 0.0091f
C198 B.n119 VSUBS 0.0091f
C199 B.n120 VSUBS 0.0091f
C200 B.n121 VSUBS 0.0091f
C201 B.n122 VSUBS 0.0091f
C202 B.n123 VSUBS 0.0091f
C203 B.n124 VSUBS 0.0091f
C204 B.n125 VSUBS 0.0091f
C205 B.n126 VSUBS 0.020657f
C206 B.n127 VSUBS 0.020657f
C207 B.n128 VSUBS 0.022434f
C208 B.n129 VSUBS 0.0091f
C209 B.n130 VSUBS 0.0091f
C210 B.n131 VSUBS 0.0091f
C211 B.n132 VSUBS 0.0091f
C212 B.n133 VSUBS 0.0091f
C213 B.n134 VSUBS 0.0091f
C214 B.n135 VSUBS 0.0091f
C215 B.n136 VSUBS 0.0091f
C216 B.n137 VSUBS 0.0091f
C217 B.n138 VSUBS 0.0091f
C218 B.n139 VSUBS 0.0091f
C219 B.n140 VSUBS 0.0091f
C220 B.n141 VSUBS 0.0091f
C221 B.n142 VSUBS 0.0091f
C222 B.n143 VSUBS 0.0091f
C223 B.n144 VSUBS 0.0091f
C224 B.n145 VSUBS 0.0091f
C225 B.n146 VSUBS 0.0091f
C226 B.n147 VSUBS 0.0091f
C227 B.n148 VSUBS 0.0091f
C228 B.n149 VSUBS 0.0091f
C229 B.n150 VSUBS 0.0091f
C230 B.n151 VSUBS 0.0091f
C231 B.n152 VSUBS 0.0091f
C232 B.n153 VSUBS 0.0091f
C233 B.n154 VSUBS 0.0091f
C234 B.n155 VSUBS 0.0091f
C235 B.n156 VSUBS 0.0091f
C236 B.n157 VSUBS 0.0091f
C237 B.n158 VSUBS 0.0091f
C238 B.n159 VSUBS 0.0091f
C239 B.n160 VSUBS 0.0091f
C240 B.n161 VSUBS 0.0091f
C241 B.n162 VSUBS 0.0091f
C242 B.n163 VSUBS 0.0091f
C243 B.n164 VSUBS 0.0091f
C244 B.n165 VSUBS 0.0091f
C245 B.n166 VSUBS 0.0091f
C246 B.n167 VSUBS 0.0091f
C247 B.n168 VSUBS 0.0091f
C248 B.n169 VSUBS 0.0091f
C249 B.n170 VSUBS 0.0091f
C250 B.n171 VSUBS 0.0091f
C251 B.n172 VSUBS 0.0091f
C252 B.n173 VSUBS 0.0091f
C253 B.n174 VSUBS 0.0091f
C254 B.n175 VSUBS 0.0091f
C255 B.n176 VSUBS 0.006022f
C256 B.n177 VSUBS 0.021083f
C257 B.n178 VSUBS 0.007628f
C258 B.n179 VSUBS 0.0091f
C259 B.n180 VSUBS 0.0091f
C260 B.n181 VSUBS 0.0091f
C261 B.n182 VSUBS 0.0091f
C262 B.n183 VSUBS 0.0091f
C263 B.n184 VSUBS 0.0091f
C264 B.n185 VSUBS 0.0091f
C265 B.n186 VSUBS 0.0091f
C266 B.n187 VSUBS 0.0091f
C267 B.n188 VSUBS 0.0091f
C268 B.n189 VSUBS 0.0091f
C269 B.t11 VSUBS 0.362586f
C270 B.t10 VSUBS 0.369494f
C271 B.t9 VSUBS 0.142868f
C272 B.n190 VSUBS 0.111761f
C273 B.n191 VSUBS 0.080614f
C274 B.n192 VSUBS 0.021083f
C275 B.n193 VSUBS 0.007628f
C276 B.n194 VSUBS 0.0091f
C277 B.n195 VSUBS 0.0091f
C278 B.n196 VSUBS 0.0091f
C279 B.n197 VSUBS 0.0091f
C280 B.n198 VSUBS 0.0091f
C281 B.n199 VSUBS 0.0091f
C282 B.n200 VSUBS 0.0091f
C283 B.n201 VSUBS 0.0091f
C284 B.n202 VSUBS 0.0091f
C285 B.n203 VSUBS 0.0091f
C286 B.n204 VSUBS 0.0091f
C287 B.n205 VSUBS 0.0091f
C288 B.n206 VSUBS 0.0091f
C289 B.n207 VSUBS 0.0091f
C290 B.n208 VSUBS 0.0091f
C291 B.n209 VSUBS 0.0091f
C292 B.n210 VSUBS 0.0091f
C293 B.n211 VSUBS 0.0091f
C294 B.n212 VSUBS 0.0091f
C295 B.n213 VSUBS 0.0091f
C296 B.n214 VSUBS 0.0091f
C297 B.n215 VSUBS 0.0091f
C298 B.n216 VSUBS 0.0091f
C299 B.n217 VSUBS 0.0091f
C300 B.n218 VSUBS 0.0091f
C301 B.n219 VSUBS 0.0091f
C302 B.n220 VSUBS 0.0091f
C303 B.n221 VSUBS 0.0091f
C304 B.n222 VSUBS 0.0091f
C305 B.n223 VSUBS 0.0091f
C306 B.n224 VSUBS 0.0091f
C307 B.n225 VSUBS 0.0091f
C308 B.n226 VSUBS 0.0091f
C309 B.n227 VSUBS 0.0091f
C310 B.n228 VSUBS 0.0091f
C311 B.n229 VSUBS 0.0091f
C312 B.n230 VSUBS 0.0091f
C313 B.n231 VSUBS 0.0091f
C314 B.n232 VSUBS 0.0091f
C315 B.n233 VSUBS 0.0091f
C316 B.n234 VSUBS 0.0091f
C317 B.n235 VSUBS 0.0091f
C318 B.n236 VSUBS 0.0091f
C319 B.n237 VSUBS 0.0091f
C320 B.n238 VSUBS 0.0091f
C321 B.n239 VSUBS 0.0091f
C322 B.n240 VSUBS 0.0091f
C323 B.n241 VSUBS 0.0091f
C324 B.n242 VSUBS 0.0091f
C325 B.n243 VSUBS 0.022434f
C326 B.n244 VSUBS 0.020657f
C327 B.n245 VSUBS 0.021713f
C328 B.n246 VSUBS 0.0091f
C329 B.n247 VSUBS 0.0091f
C330 B.n248 VSUBS 0.0091f
C331 B.n249 VSUBS 0.0091f
C332 B.n250 VSUBS 0.0091f
C333 B.n251 VSUBS 0.0091f
C334 B.n252 VSUBS 0.0091f
C335 B.n253 VSUBS 0.0091f
C336 B.n254 VSUBS 0.0091f
C337 B.n255 VSUBS 0.0091f
C338 B.n256 VSUBS 0.0091f
C339 B.n257 VSUBS 0.0091f
C340 B.n258 VSUBS 0.0091f
C341 B.n259 VSUBS 0.0091f
C342 B.n260 VSUBS 0.0091f
C343 B.n261 VSUBS 0.0091f
C344 B.n262 VSUBS 0.0091f
C345 B.n263 VSUBS 0.0091f
C346 B.n264 VSUBS 0.0091f
C347 B.n265 VSUBS 0.0091f
C348 B.n266 VSUBS 0.0091f
C349 B.n267 VSUBS 0.0091f
C350 B.n268 VSUBS 0.0091f
C351 B.n269 VSUBS 0.0091f
C352 B.n270 VSUBS 0.0091f
C353 B.n271 VSUBS 0.0091f
C354 B.n272 VSUBS 0.0091f
C355 B.n273 VSUBS 0.0091f
C356 B.n274 VSUBS 0.0091f
C357 B.n275 VSUBS 0.0091f
C358 B.n276 VSUBS 0.0091f
C359 B.n277 VSUBS 0.0091f
C360 B.n278 VSUBS 0.0091f
C361 B.n279 VSUBS 0.0091f
C362 B.n280 VSUBS 0.0091f
C363 B.n281 VSUBS 0.0091f
C364 B.n282 VSUBS 0.0091f
C365 B.n283 VSUBS 0.0091f
C366 B.n284 VSUBS 0.0091f
C367 B.n285 VSUBS 0.020657f
C368 B.n286 VSUBS 0.022434f
C369 B.n287 VSUBS 0.022434f
C370 B.n288 VSUBS 0.0091f
C371 B.n289 VSUBS 0.0091f
C372 B.n290 VSUBS 0.0091f
C373 B.n291 VSUBS 0.0091f
C374 B.n292 VSUBS 0.0091f
C375 B.n293 VSUBS 0.0091f
C376 B.n294 VSUBS 0.0091f
C377 B.n295 VSUBS 0.0091f
C378 B.n296 VSUBS 0.0091f
C379 B.n297 VSUBS 0.0091f
C380 B.n298 VSUBS 0.0091f
C381 B.n299 VSUBS 0.0091f
C382 B.n300 VSUBS 0.0091f
C383 B.n301 VSUBS 0.0091f
C384 B.n302 VSUBS 0.0091f
C385 B.n303 VSUBS 0.0091f
C386 B.n304 VSUBS 0.0091f
C387 B.n305 VSUBS 0.0091f
C388 B.n306 VSUBS 0.0091f
C389 B.n307 VSUBS 0.0091f
C390 B.n308 VSUBS 0.0091f
C391 B.n309 VSUBS 0.0091f
C392 B.n310 VSUBS 0.0091f
C393 B.n311 VSUBS 0.0091f
C394 B.n312 VSUBS 0.0091f
C395 B.n313 VSUBS 0.0091f
C396 B.n314 VSUBS 0.0091f
C397 B.n315 VSUBS 0.0091f
C398 B.n316 VSUBS 0.0091f
C399 B.n317 VSUBS 0.0091f
C400 B.n318 VSUBS 0.0091f
C401 B.n319 VSUBS 0.0091f
C402 B.n320 VSUBS 0.0091f
C403 B.n321 VSUBS 0.0091f
C404 B.n322 VSUBS 0.0091f
C405 B.n323 VSUBS 0.0091f
C406 B.n324 VSUBS 0.0091f
C407 B.n325 VSUBS 0.0091f
C408 B.n326 VSUBS 0.0091f
C409 B.n327 VSUBS 0.0091f
C410 B.n328 VSUBS 0.0091f
C411 B.n329 VSUBS 0.0091f
C412 B.n330 VSUBS 0.0091f
C413 B.n331 VSUBS 0.0091f
C414 B.n332 VSUBS 0.0091f
C415 B.n333 VSUBS 0.0091f
C416 B.n334 VSUBS 0.0091f
C417 B.n335 VSUBS 0.006022f
C418 B.n336 VSUBS 0.021083f
C419 B.n337 VSUBS 0.007628f
C420 B.n338 VSUBS 0.0091f
C421 B.n339 VSUBS 0.0091f
C422 B.n340 VSUBS 0.0091f
C423 B.n341 VSUBS 0.0091f
C424 B.n342 VSUBS 0.0091f
C425 B.n343 VSUBS 0.0091f
C426 B.n344 VSUBS 0.0091f
C427 B.n345 VSUBS 0.0091f
C428 B.n346 VSUBS 0.0091f
C429 B.n347 VSUBS 0.0091f
C430 B.n348 VSUBS 0.0091f
C431 B.n349 VSUBS 0.007628f
C432 B.n350 VSUBS 0.021083f
C433 B.n351 VSUBS 0.006022f
C434 B.n352 VSUBS 0.0091f
C435 B.n353 VSUBS 0.0091f
C436 B.n354 VSUBS 0.0091f
C437 B.n355 VSUBS 0.0091f
C438 B.n356 VSUBS 0.0091f
C439 B.n357 VSUBS 0.0091f
C440 B.n358 VSUBS 0.0091f
C441 B.n359 VSUBS 0.0091f
C442 B.n360 VSUBS 0.0091f
C443 B.n361 VSUBS 0.0091f
C444 B.n362 VSUBS 0.0091f
C445 B.n363 VSUBS 0.0091f
C446 B.n364 VSUBS 0.0091f
C447 B.n365 VSUBS 0.0091f
C448 B.n366 VSUBS 0.0091f
C449 B.n367 VSUBS 0.0091f
C450 B.n368 VSUBS 0.0091f
C451 B.n369 VSUBS 0.0091f
C452 B.n370 VSUBS 0.0091f
C453 B.n371 VSUBS 0.0091f
C454 B.n372 VSUBS 0.0091f
C455 B.n373 VSUBS 0.0091f
C456 B.n374 VSUBS 0.0091f
C457 B.n375 VSUBS 0.0091f
C458 B.n376 VSUBS 0.0091f
C459 B.n377 VSUBS 0.0091f
C460 B.n378 VSUBS 0.0091f
C461 B.n379 VSUBS 0.0091f
C462 B.n380 VSUBS 0.0091f
C463 B.n381 VSUBS 0.0091f
C464 B.n382 VSUBS 0.0091f
C465 B.n383 VSUBS 0.0091f
C466 B.n384 VSUBS 0.0091f
C467 B.n385 VSUBS 0.0091f
C468 B.n386 VSUBS 0.0091f
C469 B.n387 VSUBS 0.0091f
C470 B.n388 VSUBS 0.0091f
C471 B.n389 VSUBS 0.0091f
C472 B.n390 VSUBS 0.0091f
C473 B.n391 VSUBS 0.0091f
C474 B.n392 VSUBS 0.0091f
C475 B.n393 VSUBS 0.0091f
C476 B.n394 VSUBS 0.0091f
C477 B.n395 VSUBS 0.0091f
C478 B.n396 VSUBS 0.0091f
C479 B.n397 VSUBS 0.0091f
C480 B.n398 VSUBS 0.0091f
C481 B.n399 VSUBS 0.022434f
C482 B.n400 VSUBS 0.022434f
C483 B.n401 VSUBS 0.020657f
C484 B.n402 VSUBS 0.0091f
C485 B.n403 VSUBS 0.0091f
C486 B.n404 VSUBS 0.0091f
C487 B.n405 VSUBS 0.0091f
C488 B.n406 VSUBS 0.0091f
C489 B.n407 VSUBS 0.0091f
C490 B.n408 VSUBS 0.0091f
C491 B.n409 VSUBS 0.0091f
C492 B.n410 VSUBS 0.0091f
C493 B.n411 VSUBS 0.0091f
C494 B.n412 VSUBS 0.0091f
C495 B.n413 VSUBS 0.0091f
C496 B.n414 VSUBS 0.0091f
C497 B.n415 VSUBS 0.0091f
C498 B.n416 VSUBS 0.0091f
C499 B.n417 VSUBS 0.0091f
C500 B.n418 VSUBS 0.0091f
C501 B.n419 VSUBS 0.011875f
C502 B.n420 VSUBS 0.01265f
C503 B.n421 VSUBS 0.025155f
.ends

