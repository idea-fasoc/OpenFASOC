* NGSPICE file created from diff_pair_sample_0175.ext - technology: sky130A

.subckt diff_pair_sample_0175 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t1 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X1 VDD2.t3 VN.t1 VTAIL.t18 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3
X2 B.t11 B.t9 B.t10 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3
X3 VDD2.t6 VN.t2 VTAIL.t17 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3
X4 B.t8 B.t6 B.t7 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3
X5 VDD2.t8 VN.t3 VTAIL.t16 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X6 VDD1.t9 VP.t0 VTAIL.t9 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3
X7 VDD1.t8 VP.t1 VTAIL.t7 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3
X8 VDD2.t2 VN.t4 VTAIL.t15 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3
X9 VTAIL.t14 VN.t5 VDD2.t5 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X10 VTAIL.t8 VP.t2 VDD1.t7 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X11 VDD2.t7 VN.t6 VTAIL.t13 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X12 VDD1.t6 VP.t3 VTAIL.t6 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3
X13 VDD1.t5 VP.t4 VTAIL.t0 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=3.5685 ps=19.08 w=9.15 l=3
X14 VTAIL.t12 VN.t7 VDD2.t9 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X15 B.t5 B.t3 B.t4 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3
X16 VDD1.t4 VP.t5 VTAIL.t3 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X17 VTAIL.t5 VP.t6 VDD1.t3 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X18 VTAIL.t2 VP.t7 VDD1.t2 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X19 VDD1.t1 VP.t8 VTAIL.t4 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X20 VTAIL.t1 VP.t9 VDD1.t0 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X21 VTAIL.t11 VN.t8 VDD2.t4 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=1.50975 pd=9.48 as=1.50975 ps=9.48 w=9.15 l=3
X22 VDD2.t0 VN.t9 VTAIL.t10 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=1.50975 ps=9.48 w=9.15 l=3
X23 B.t2 B.t0 B.t1 w_n4966_n2798# sky130_fd_pr__pfet_01v8 ad=3.5685 pd=19.08 as=0 ps=0 w=9.15 l=3
R0 VN.n90 VN.n89 161.3
R1 VN.n88 VN.n47 161.3
R2 VN.n87 VN.n86 161.3
R3 VN.n85 VN.n48 161.3
R4 VN.n84 VN.n83 161.3
R5 VN.n82 VN.n49 161.3
R6 VN.n80 VN.n79 161.3
R7 VN.n78 VN.n50 161.3
R8 VN.n77 VN.n76 161.3
R9 VN.n75 VN.n51 161.3
R10 VN.n74 VN.n73 161.3
R11 VN.n72 VN.n52 161.3
R12 VN.n71 VN.n70 161.3
R13 VN.n68 VN.n53 161.3
R14 VN.n67 VN.n66 161.3
R15 VN.n65 VN.n54 161.3
R16 VN.n64 VN.n63 161.3
R17 VN.n62 VN.n55 161.3
R18 VN.n61 VN.n60 161.3
R19 VN.n59 VN.n56 161.3
R20 VN.n44 VN.n43 161.3
R21 VN.n42 VN.n1 161.3
R22 VN.n41 VN.n40 161.3
R23 VN.n39 VN.n2 161.3
R24 VN.n38 VN.n37 161.3
R25 VN.n36 VN.n3 161.3
R26 VN.n34 VN.n33 161.3
R27 VN.n32 VN.n4 161.3
R28 VN.n31 VN.n30 161.3
R29 VN.n29 VN.n5 161.3
R30 VN.n28 VN.n27 161.3
R31 VN.n26 VN.n6 161.3
R32 VN.n25 VN.n24 161.3
R33 VN.n22 VN.n7 161.3
R34 VN.n21 VN.n20 161.3
R35 VN.n19 VN.n8 161.3
R36 VN.n18 VN.n17 161.3
R37 VN.n16 VN.n9 161.3
R38 VN.n15 VN.n14 161.3
R39 VN.n13 VN.n10 161.3
R40 VN.n58 VN.t4 105.207
R41 VN.n12 VN.t1 105.207
R42 VN.n11 VN.t7 73.5055
R43 VN.n23 VN.t6 73.5055
R44 VN.n35 VN.t0 73.5055
R45 VN.n0 VN.t2 73.5055
R46 VN.n57 VN.t5 73.5055
R47 VN.n69 VN.t3 73.5055
R48 VN.n81 VN.t8 73.5055
R49 VN.n46 VN.t9 73.5055
R50 VN.n45 VN.n0 70.0045
R51 VN.n91 VN.n46 70.0045
R52 VN.n12 VN.n11 69.746
R53 VN.n58 VN.n57 69.746
R54 VN.n41 VN.n2 56.5193
R55 VN.n87 VN.n48 56.5193
R56 VN VN.n91 53.4185
R57 VN.n17 VN.n8 48.7492
R58 VN.n29 VN.n28 48.7492
R59 VN.n63 VN.n54 48.7492
R60 VN.n75 VN.n74 48.7492
R61 VN.n17 VN.n16 32.2376
R62 VN.n30 VN.n29 32.2376
R63 VN.n63 VN.n62 32.2376
R64 VN.n76 VN.n75 32.2376
R65 VN.n15 VN.n10 24.4675
R66 VN.n16 VN.n15 24.4675
R67 VN.n21 VN.n8 24.4675
R68 VN.n22 VN.n21 24.4675
R69 VN.n24 VN.n6 24.4675
R70 VN.n28 VN.n6 24.4675
R71 VN.n30 VN.n4 24.4675
R72 VN.n34 VN.n4 24.4675
R73 VN.n37 VN.n36 24.4675
R74 VN.n37 VN.n2 24.4675
R75 VN.n42 VN.n41 24.4675
R76 VN.n43 VN.n42 24.4675
R77 VN.n62 VN.n61 24.4675
R78 VN.n61 VN.n56 24.4675
R79 VN.n74 VN.n52 24.4675
R80 VN.n70 VN.n52 24.4675
R81 VN.n68 VN.n67 24.4675
R82 VN.n67 VN.n54 24.4675
R83 VN.n83 VN.n48 24.4675
R84 VN.n83 VN.n82 24.4675
R85 VN.n80 VN.n50 24.4675
R86 VN.n76 VN.n50 24.4675
R87 VN.n89 VN.n88 24.4675
R88 VN.n88 VN.n87 24.4675
R89 VN.n36 VN.n35 20.5528
R90 VN.n82 VN.n81 20.5528
R91 VN.n43 VN.n0 20.0634
R92 VN.n89 VN.n46 20.0634
R93 VN.n23 VN.n22 12.234
R94 VN.n24 VN.n23 12.234
R95 VN.n70 VN.n69 12.234
R96 VN.n69 VN.n68 12.234
R97 VN.n59 VN.n58 5.54917
R98 VN.n13 VN.n12 5.54917
R99 VN.n11 VN.n10 3.91522
R100 VN.n35 VN.n34 3.91522
R101 VN.n57 VN.n56 3.91522
R102 VN.n81 VN.n80 3.91522
R103 VN.n91 VN.n90 0.354971
R104 VN.n45 VN.n44 0.354971
R105 VN VN.n45 0.26696
R106 VN.n90 VN.n47 0.189894
R107 VN.n86 VN.n47 0.189894
R108 VN.n86 VN.n85 0.189894
R109 VN.n85 VN.n84 0.189894
R110 VN.n84 VN.n49 0.189894
R111 VN.n79 VN.n49 0.189894
R112 VN.n79 VN.n78 0.189894
R113 VN.n78 VN.n77 0.189894
R114 VN.n77 VN.n51 0.189894
R115 VN.n73 VN.n51 0.189894
R116 VN.n73 VN.n72 0.189894
R117 VN.n72 VN.n71 0.189894
R118 VN.n71 VN.n53 0.189894
R119 VN.n66 VN.n53 0.189894
R120 VN.n66 VN.n65 0.189894
R121 VN.n65 VN.n64 0.189894
R122 VN.n64 VN.n55 0.189894
R123 VN.n60 VN.n55 0.189894
R124 VN.n60 VN.n59 0.189894
R125 VN.n14 VN.n13 0.189894
R126 VN.n14 VN.n9 0.189894
R127 VN.n18 VN.n9 0.189894
R128 VN.n19 VN.n18 0.189894
R129 VN.n20 VN.n19 0.189894
R130 VN.n20 VN.n7 0.189894
R131 VN.n25 VN.n7 0.189894
R132 VN.n26 VN.n25 0.189894
R133 VN.n27 VN.n26 0.189894
R134 VN.n27 VN.n5 0.189894
R135 VN.n31 VN.n5 0.189894
R136 VN.n32 VN.n31 0.189894
R137 VN.n33 VN.n32 0.189894
R138 VN.n33 VN.n3 0.189894
R139 VN.n38 VN.n3 0.189894
R140 VN.n39 VN.n38 0.189894
R141 VN.n40 VN.n39 0.189894
R142 VN.n40 VN.n1 0.189894
R143 VN.n44 VN.n1 0.189894
R144 VDD2.n1 VDD2.t3 84.4747
R145 VDD2.n4 VDD2.t0 81.6042
R146 VDD2.n3 VDD2.n2 80.1492
R147 VDD2 VDD2.n7 80.1466
R148 VDD2.n6 VDD2.n5 78.0517
R149 VDD2.n1 VDD2.n0 78.0515
R150 VDD2.n4 VDD2.n3 45.239
R151 VDD2.n7 VDD2.t5 3.55296
R152 VDD2.n7 VDD2.t2 3.55296
R153 VDD2.n5 VDD2.t4 3.55296
R154 VDD2.n5 VDD2.t8 3.55296
R155 VDD2.n2 VDD2.t1 3.55296
R156 VDD2.n2 VDD2.t6 3.55296
R157 VDD2.n0 VDD2.t9 3.55296
R158 VDD2.n0 VDD2.t7 3.55296
R159 VDD2.n6 VDD2.n4 2.87119
R160 VDD2 VDD2.n6 0.776362
R161 VDD2.n3 VDD2.n1 0.662826
R162 VTAIL.n16 VTAIL.t0 64.9254
R163 VTAIL.n11 VTAIL.t15 64.9254
R164 VTAIL.n17 VTAIL.t17 64.9252
R165 VTAIL.n2 VTAIL.t9 64.9252
R166 VTAIL.n15 VTAIL.n14 61.3729
R167 VTAIL.n13 VTAIL.n12 61.3729
R168 VTAIL.n10 VTAIL.n9 61.3729
R169 VTAIL.n8 VTAIL.n7 61.3729
R170 VTAIL.n19 VTAIL.n18 61.3727
R171 VTAIL.n1 VTAIL.n0 61.3727
R172 VTAIL.n4 VTAIL.n3 61.3727
R173 VTAIL.n6 VTAIL.n5 61.3727
R174 VTAIL.n8 VTAIL.n6 25.9962
R175 VTAIL.n17 VTAIL.n16 23.1255
R176 VTAIL.n18 VTAIL.t13 3.55296
R177 VTAIL.n18 VTAIL.t19 3.55296
R178 VTAIL.n0 VTAIL.t18 3.55296
R179 VTAIL.n0 VTAIL.t12 3.55296
R180 VTAIL.n3 VTAIL.t3 3.55296
R181 VTAIL.n3 VTAIL.t1 3.55296
R182 VTAIL.n5 VTAIL.t7 3.55296
R183 VTAIL.n5 VTAIL.t5 3.55296
R184 VTAIL.n14 VTAIL.t4 3.55296
R185 VTAIL.n14 VTAIL.t2 3.55296
R186 VTAIL.n12 VTAIL.t6 3.55296
R187 VTAIL.n12 VTAIL.t8 3.55296
R188 VTAIL.n9 VTAIL.t16 3.55296
R189 VTAIL.n9 VTAIL.t14 3.55296
R190 VTAIL.n7 VTAIL.t10 3.55296
R191 VTAIL.n7 VTAIL.t11 3.55296
R192 VTAIL.n10 VTAIL.n8 2.87119
R193 VTAIL.n11 VTAIL.n10 2.87119
R194 VTAIL.n15 VTAIL.n13 2.87119
R195 VTAIL.n16 VTAIL.n15 2.87119
R196 VTAIL.n6 VTAIL.n4 2.87119
R197 VTAIL.n4 VTAIL.n2 2.87119
R198 VTAIL.n19 VTAIL.n17 2.87119
R199 VTAIL VTAIL.n1 2.21171
R200 VTAIL.n13 VTAIL.n11 1.90567
R201 VTAIL.n2 VTAIL.n1 1.90567
R202 VTAIL VTAIL.n19 0.659983
R203 B.n639 B.n638 585
R204 B.n640 B.n77 585
R205 B.n642 B.n641 585
R206 B.n643 B.n76 585
R207 B.n645 B.n644 585
R208 B.n646 B.n75 585
R209 B.n648 B.n647 585
R210 B.n649 B.n74 585
R211 B.n651 B.n650 585
R212 B.n652 B.n73 585
R213 B.n654 B.n653 585
R214 B.n655 B.n72 585
R215 B.n657 B.n656 585
R216 B.n658 B.n71 585
R217 B.n660 B.n659 585
R218 B.n661 B.n70 585
R219 B.n663 B.n662 585
R220 B.n664 B.n69 585
R221 B.n666 B.n665 585
R222 B.n667 B.n68 585
R223 B.n669 B.n668 585
R224 B.n670 B.n67 585
R225 B.n672 B.n671 585
R226 B.n673 B.n66 585
R227 B.n675 B.n674 585
R228 B.n676 B.n65 585
R229 B.n678 B.n677 585
R230 B.n679 B.n64 585
R231 B.n681 B.n680 585
R232 B.n682 B.n63 585
R233 B.n684 B.n683 585
R234 B.n685 B.n62 585
R235 B.n687 B.n686 585
R236 B.n689 B.n59 585
R237 B.n691 B.n690 585
R238 B.n692 B.n58 585
R239 B.n694 B.n693 585
R240 B.n695 B.n57 585
R241 B.n697 B.n696 585
R242 B.n698 B.n56 585
R243 B.n700 B.n699 585
R244 B.n701 B.n55 585
R245 B.n703 B.n702 585
R246 B.n705 B.n704 585
R247 B.n706 B.n51 585
R248 B.n708 B.n707 585
R249 B.n709 B.n50 585
R250 B.n711 B.n710 585
R251 B.n712 B.n49 585
R252 B.n714 B.n713 585
R253 B.n715 B.n48 585
R254 B.n717 B.n716 585
R255 B.n718 B.n47 585
R256 B.n720 B.n719 585
R257 B.n721 B.n46 585
R258 B.n723 B.n722 585
R259 B.n724 B.n45 585
R260 B.n726 B.n725 585
R261 B.n727 B.n44 585
R262 B.n729 B.n728 585
R263 B.n730 B.n43 585
R264 B.n732 B.n731 585
R265 B.n733 B.n42 585
R266 B.n735 B.n734 585
R267 B.n736 B.n41 585
R268 B.n738 B.n737 585
R269 B.n739 B.n40 585
R270 B.n741 B.n740 585
R271 B.n742 B.n39 585
R272 B.n744 B.n743 585
R273 B.n745 B.n38 585
R274 B.n747 B.n746 585
R275 B.n748 B.n37 585
R276 B.n750 B.n749 585
R277 B.n751 B.n36 585
R278 B.n753 B.n752 585
R279 B.n637 B.n78 585
R280 B.n636 B.n635 585
R281 B.n634 B.n79 585
R282 B.n633 B.n632 585
R283 B.n631 B.n80 585
R284 B.n630 B.n629 585
R285 B.n628 B.n81 585
R286 B.n627 B.n626 585
R287 B.n625 B.n82 585
R288 B.n624 B.n623 585
R289 B.n622 B.n83 585
R290 B.n621 B.n620 585
R291 B.n619 B.n84 585
R292 B.n618 B.n617 585
R293 B.n616 B.n85 585
R294 B.n615 B.n614 585
R295 B.n613 B.n86 585
R296 B.n612 B.n611 585
R297 B.n610 B.n87 585
R298 B.n609 B.n608 585
R299 B.n607 B.n88 585
R300 B.n606 B.n605 585
R301 B.n604 B.n89 585
R302 B.n603 B.n602 585
R303 B.n601 B.n90 585
R304 B.n600 B.n599 585
R305 B.n598 B.n91 585
R306 B.n597 B.n596 585
R307 B.n595 B.n92 585
R308 B.n594 B.n593 585
R309 B.n592 B.n93 585
R310 B.n591 B.n590 585
R311 B.n589 B.n94 585
R312 B.n588 B.n587 585
R313 B.n586 B.n95 585
R314 B.n585 B.n584 585
R315 B.n583 B.n96 585
R316 B.n582 B.n581 585
R317 B.n580 B.n97 585
R318 B.n579 B.n578 585
R319 B.n577 B.n98 585
R320 B.n576 B.n575 585
R321 B.n574 B.n99 585
R322 B.n573 B.n572 585
R323 B.n571 B.n100 585
R324 B.n570 B.n569 585
R325 B.n568 B.n101 585
R326 B.n567 B.n566 585
R327 B.n565 B.n102 585
R328 B.n564 B.n563 585
R329 B.n562 B.n103 585
R330 B.n561 B.n560 585
R331 B.n559 B.n104 585
R332 B.n558 B.n557 585
R333 B.n556 B.n105 585
R334 B.n555 B.n554 585
R335 B.n553 B.n106 585
R336 B.n552 B.n551 585
R337 B.n550 B.n107 585
R338 B.n549 B.n548 585
R339 B.n547 B.n108 585
R340 B.n546 B.n545 585
R341 B.n544 B.n109 585
R342 B.n543 B.n542 585
R343 B.n541 B.n110 585
R344 B.n540 B.n539 585
R345 B.n538 B.n111 585
R346 B.n537 B.n536 585
R347 B.n535 B.n112 585
R348 B.n534 B.n533 585
R349 B.n532 B.n113 585
R350 B.n531 B.n530 585
R351 B.n529 B.n114 585
R352 B.n528 B.n527 585
R353 B.n526 B.n115 585
R354 B.n525 B.n524 585
R355 B.n523 B.n116 585
R356 B.n522 B.n521 585
R357 B.n520 B.n117 585
R358 B.n519 B.n518 585
R359 B.n517 B.n118 585
R360 B.n516 B.n515 585
R361 B.n514 B.n119 585
R362 B.n513 B.n512 585
R363 B.n511 B.n120 585
R364 B.n510 B.n509 585
R365 B.n508 B.n121 585
R366 B.n507 B.n506 585
R367 B.n505 B.n122 585
R368 B.n504 B.n503 585
R369 B.n502 B.n123 585
R370 B.n501 B.n500 585
R371 B.n499 B.n124 585
R372 B.n498 B.n497 585
R373 B.n496 B.n125 585
R374 B.n495 B.n494 585
R375 B.n493 B.n126 585
R376 B.n492 B.n491 585
R377 B.n490 B.n127 585
R378 B.n489 B.n488 585
R379 B.n487 B.n128 585
R380 B.n486 B.n485 585
R381 B.n484 B.n129 585
R382 B.n483 B.n482 585
R383 B.n481 B.n130 585
R384 B.n480 B.n479 585
R385 B.n478 B.n131 585
R386 B.n477 B.n476 585
R387 B.n475 B.n132 585
R388 B.n474 B.n473 585
R389 B.n472 B.n133 585
R390 B.n471 B.n470 585
R391 B.n469 B.n134 585
R392 B.n468 B.n467 585
R393 B.n466 B.n135 585
R394 B.n465 B.n464 585
R395 B.n463 B.n136 585
R396 B.n462 B.n461 585
R397 B.n460 B.n137 585
R398 B.n459 B.n458 585
R399 B.n457 B.n138 585
R400 B.n456 B.n455 585
R401 B.n454 B.n139 585
R402 B.n453 B.n452 585
R403 B.n451 B.n140 585
R404 B.n450 B.n449 585
R405 B.n448 B.n141 585
R406 B.n447 B.n446 585
R407 B.n445 B.n142 585
R408 B.n444 B.n443 585
R409 B.n442 B.n143 585
R410 B.n441 B.n440 585
R411 B.n439 B.n144 585
R412 B.n438 B.n437 585
R413 B.n436 B.n145 585
R414 B.n321 B.n320 585
R415 B.n322 B.n187 585
R416 B.n324 B.n323 585
R417 B.n325 B.n186 585
R418 B.n327 B.n326 585
R419 B.n328 B.n185 585
R420 B.n330 B.n329 585
R421 B.n331 B.n184 585
R422 B.n333 B.n332 585
R423 B.n334 B.n183 585
R424 B.n336 B.n335 585
R425 B.n337 B.n182 585
R426 B.n339 B.n338 585
R427 B.n340 B.n181 585
R428 B.n342 B.n341 585
R429 B.n343 B.n180 585
R430 B.n345 B.n344 585
R431 B.n346 B.n179 585
R432 B.n348 B.n347 585
R433 B.n349 B.n178 585
R434 B.n351 B.n350 585
R435 B.n352 B.n177 585
R436 B.n354 B.n353 585
R437 B.n355 B.n176 585
R438 B.n357 B.n356 585
R439 B.n358 B.n175 585
R440 B.n360 B.n359 585
R441 B.n361 B.n174 585
R442 B.n363 B.n362 585
R443 B.n364 B.n173 585
R444 B.n366 B.n365 585
R445 B.n367 B.n172 585
R446 B.n369 B.n368 585
R447 B.n371 B.n169 585
R448 B.n373 B.n372 585
R449 B.n374 B.n168 585
R450 B.n376 B.n375 585
R451 B.n377 B.n167 585
R452 B.n379 B.n378 585
R453 B.n380 B.n166 585
R454 B.n382 B.n381 585
R455 B.n383 B.n165 585
R456 B.n385 B.n384 585
R457 B.n387 B.n386 585
R458 B.n388 B.n161 585
R459 B.n390 B.n389 585
R460 B.n391 B.n160 585
R461 B.n393 B.n392 585
R462 B.n394 B.n159 585
R463 B.n396 B.n395 585
R464 B.n397 B.n158 585
R465 B.n399 B.n398 585
R466 B.n400 B.n157 585
R467 B.n402 B.n401 585
R468 B.n403 B.n156 585
R469 B.n405 B.n404 585
R470 B.n406 B.n155 585
R471 B.n408 B.n407 585
R472 B.n409 B.n154 585
R473 B.n411 B.n410 585
R474 B.n412 B.n153 585
R475 B.n414 B.n413 585
R476 B.n415 B.n152 585
R477 B.n417 B.n416 585
R478 B.n418 B.n151 585
R479 B.n420 B.n419 585
R480 B.n421 B.n150 585
R481 B.n423 B.n422 585
R482 B.n424 B.n149 585
R483 B.n426 B.n425 585
R484 B.n427 B.n148 585
R485 B.n429 B.n428 585
R486 B.n430 B.n147 585
R487 B.n432 B.n431 585
R488 B.n433 B.n146 585
R489 B.n435 B.n434 585
R490 B.n319 B.n188 585
R491 B.n318 B.n317 585
R492 B.n316 B.n189 585
R493 B.n315 B.n314 585
R494 B.n313 B.n190 585
R495 B.n312 B.n311 585
R496 B.n310 B.n191 585
R497 B.n309 B.n308 585
R498 B.n307 B.n192 585
R499 B.n306 B.n305 585
R500 B.n304 B.n193 585
R501 B.n303 B.n302 585
R502 B.n301 B.n194 585
R503 B.n300 B.n299 585
R504 B.n298 B.n195 585
R505 B.n297 B.n296 585
R506 B.n295 B.n196 585
R507 B.n294 B.n293 585
R508 B.n292 B.n197 585
R509 B.n291 B.n290 585
R510 B.n289 B.n198 585
R511 B.n288 B.n287 585
R512 B.n286 B.n199 585
R513 B.n285 B.n284 585
R514 B.n283 B.n200 585
R515 B.n282 B.n281 585
R516 B.n280 B.n201 585
R517 B.n279 B.n278 585
R518 B.n277 B.n202 585
R519 B.n276 B.n275 585
R520 B.n274 B.n203 585
R521 B.n273 B.n272 585
R522 B.n271 B.n204 585
R523 B.n270 B.n269 585
R524 B.n268 B.n205 585
R525 B.n267 B.n266 585
R526 B.n265 B.n206 585
R527 B.n264 B.n263 585
R528 B.n262 B.n207 585
R529 B.n261 B.n260 585
R530 B.n259 B.n208 585
R531 B.n258 B.n257 585
R532 B.n256 B.n209 585
R533 B.n255 B.n254 585
R534 B.n253 B.n210 585
R535 B.n252 B.n251 585
R536 B.n250 B.n211 585
R537 B.n249 B.n248 585
R538 B.n247 B.n212 585
R539 B.n246 B.n245 585
R540 B.n244 B.n213 585
R541 B.n243 B.n242 585
R542 B.n241 B.n214 585
R543 B.n240 B.n239 585
R544 B.n238 B.n215 585
R545 B.n237 B.n236 585
R546 B.n235 B.n216 585
R547 B.n234 B.n233 585
R548 B.n232 B.n217 585
R549 B.n231 B.n230 585
R550 B.n229 B.n218 585
R551 B.n228 B.n227 585
R552 B.n226 B.n219 585
R553 B.n225 B.n224 585
R554 B.n223 B.n220 585
R555 B.n222 B.n221 585
R556 B.n2 B.n0 585
R557 B.n853 B.n1 585
R558 B.n852 B.n851 585
R559 B.n850 B.n3 585
R560 B.n849 B.n848 585
R561 B.n847 B.n4 585
R562 B.n846 B.n845 585
R563 B.n844 B.n5 585
R564 B.n843 B.n842 585
R565 B.n841 B.n6 585
R566 B.n840 B.n839 585
R567 B.n838 B.n7 585
R568 B.n837 B.n836 585
R569 B.n835 B.n8 585
R570 B.n834 B.n833 585
R571 B.n832 B.n9 585
R572 B.n831 B.n830 585
R573 B.n829 B.n10 585
R574 B.n828 B.n827 585
R575 B.n826 B.n11 585
R576 B.n825 B.n824 585
R577 B.n823 B.n12 585
R578 B.n822 B.n821 585
R579 B.n820 B.n13 585
R580 B.n819 B.n818 585
R581 B.n817 B.n14 585
R582 B.n816 B.n815 585
R583 B.n814 B.n15 585
R584 B.n813 B.n812 585
R585 B.n811 B.n16 585
R586 B.n810 B.n809 585
R587 B.n808 B.n17 585
R588 B.n807 B.n806 585
R589 B.n805 B.n18 585
R590 B.n804 B.n803 585
R591 B.n802 B.n19 585
R592 B.n801 B.n800 585
R593 B.n799 B.n20 585
R594 B.n798 B.n797 585
R595 B.n796 B.n21 585
R596 B.n795 B.n794 585
R597 B.n793 B.n22 585
R598 B.n792 B.n791 585
R599 B.n790 B.n23 585
R600 B.n789 B.n788 585
R601 B.n787 B.n24 585
R602 B.n786 B.n785 585
R603 B.n784 B.n25 585
R604 B.n783 B.n782 585
R605 B.n781 B.n26 585
R606 B.n780 B.n779 585
R607 B.n778 B.n27 585
R608 B.n777 B.n776 585
R609 B.n775 B.n28 585
R610 B.n774 B.n773 585
R611 B.n772 B.n29 585
R612 B.n771 B.n770 585
R613 B.n769 B.n30 585
R614 B.n768 B.n767 585
R615 B.n766 B.n31 585
R616 B.n765 B.n764 585
R617 B.n763 B.n32 585
R618 B.n762 B.n761 585
R619 B.n760 B.n33 585
R620 B.n759 B.n758 585
R621 B.n757 B.n34 585
R622 B.n756 B.n755 585
R623 B.n754 B.n35 585
R624 B.n855 B.n854 585
R625 B.n320 B.n319 482.89
R626 B.n752 B.n35 482.89
R627 B.n434 B.n145 482.89
R628 B.n638 B.n637 482.89
R629 B.n162 B.t9 282.086
R630 B.n170 B.t0 282.086
R631 B.n52 B.t3 282.086
R632 B.n60 B.t6 282.086
R633 B.n162 B.t11 178.629
R634 B.n60 B.t7 178.629
R635 B.n170 B.t2 178.619
R636 B.n52 B.t4 178.619
R637 B.n319 B.n318 163.367
R638 B.n318 B.n189 163.367
R639 B.n314 B.n189 163.367
R640 B.n314 B.n313 163.367
R641 B.n313 B.n312 163.367
R642 B.n312 B.n191 163.367
R643 B.n308 B.n191 163.367
R644 B.n308 B.n307 163.367
R645 B.n307 B.n306 163.367
R646 B.n306 B.n193 163.367
R647 B.n302 B.n193 163.367
R648 B.n302 B.n301 163.367
R649 B.n301 B.n300 163.367
R650 B.n300 B.n195 163.367
R651 B.n296 B.n195 163.367
R652 B.n296 B.n295 163.367
R653 B.n295 B.n294 163.367
R654 B.n294 B.n197 163.367
R655 B.n290 B.n197 163.367
R656 B.n290 B.n289 163.367
R657 B.n289 B.n288 163.367
R658 B.n288 B.n199 163.367
R659 B.n284 B.n199 163.367
R660 B.n284 B.n283 163.367
R661 B.n283 B.n282 163.367
R662 B.n282 B.n201 163.367
R663 B.n278 B.n201 163.367
R664 B.n278 B.n277 163.367
R665 B.n277 B.n276 163.367
R666 B.n276 B.n203 163.367
R667 B.n272 B.n203 163.367
R668 B.n272 B.n271 163.367
R669 B.n271 B.n270 163.367
R670 B.n270 B.n205 163.367
R671 B.n266 B.n205 163.367
R672 B.n266 B.n265 163.367
R673 B.n265 B.n264 163.367
R674 B.n264 B.n207 163.367
R675 B.n260 B.n207 163.367
R676 B.n260 B.n259 163.367
R677 B.n259 B.n258 163.367
R678 B.n258 B.n209 163.367
R679 B.n254 B.n209 163.367
R680 B.n254 B.n253 163.367
R681 B.n253 B.n252 163.367
R682 B.n252 B.n211 163.367
R683 B.n248 B.n211 163.367
R684 B.n248 B.n247 163.367
R685 B.n247 B.n246 163.367
R686 B.n246 B.n213 163.367
R687 B.n242 B.n213 163.367
R688 B.n242 B.n241 163.367
R689 B.n241 B.n240 163.367
R690 B.n240 B.n215 163.367
R691 B.n236 B.n215 163.367
R692 B.n236 B.n235 163.367
R693 B.n235 B.n234 163.367
R694 B.n234 B.n217 163.367
R695 B.n230 B.n217 163.367
R696 B.n230 B.n229 163.367
R697 B.n229 B.n228 163.367
R698 B.n228 B.n219 163.367
R699 B.n224 B.n219 163.367
R700 B.n224 B.n223 163.367
R701 B.n223 B.n222 163.367
R702 B.n222 B.n2 163.367
R703 B.n854 B.n2 163.367
R704 B.n854 B.n853 163.367
R705 B.n853 B.n852 163.367
R706 B.n852 B.n3 163.367
R707 B.n848 B.n3 163.367
R708 B.n848 B.n847 163.367
R709 B.n847 B.n846 163.367
R710 B.n846 B.n5 163.367
R711 B.n842 B.n5 163.367
R712 B.n842 B.n841 163.367
R713 B.n841 B.n840 163.367
R714 B.n840 B.n7 163.367
R715 B.n836 B.n7 163.367
R716 B.n836 B.n835 163.367
R717 B.n835 B.n834 163.367
R718 B.n834 B.n9 163.367
R719 B.n830 B.n9 163.367
R720 B.n830 B.n829 163.367
R721 B.n829 B.n828 163.367
R722 B.n828 B.n11 163.367
R723 B.n824 B.n11 163.367
R724 B.n824 B.n823 163.367
R725 B.n823 B.n822 163.367
R726 B.n822 B.n13 163.367
R727 B.n818 B.n13 163.367
R728 B.n818 B.n817 163.367
R729 B.n817 B.n816 163.367
R730 B.n816 B.n15 163.367
R731 B.n812 B.n15 163.367
R732 B.n812 B.n811 163.367
R733 B.n811 B.n810 163.367
R734 B.n810 B.n17 163.367
R735 B.n806 B.n17 163.367
R736 B.n806 B.n805 163.367
R737 B.n805 B.n804 163.367
R738 B.n804 B.n19 163.367
R739 B.n800 B.n19 163.367
R740 B.n800 B.n799 163.367
R741 B.n799 B.n798 163.367
R742 B.n798 B.n21 163.367
R743 B.n794 B.n21 163.367
R744 B.n794 B.n793 163.367
R745 B.n793 B.n792 163.367
R746 B.n792 B.n23 163.367
R747 B.n788 B.n23 163.367
R748 B.n788 B.n787 163.367
R749 B.n787 B.n786 163.367
R750 B.n786 B.n25 163.367
R751 B.n782 B.n25 163.367
R752 B.n782 B.n781 163.367
R753 B.n781 B.n780 163.367
R754 B.n780 B.n27 163.367
R755 B.n776 B.n27 163.367
R756 B.n776 B.n775 163.367
R757 B.n775 B.n774 163.367
R758 B.n774 B.n29 163.367
R759 B.n770 B.n29 163.367
R760 B.n770 B.n769 163.367
R761 B.n769 B.n768 163.367
R762 B.n768 B.n31 163.367
R763 B.n764 B.n31 163.367
R764 B.n764 B.n763 163.367
R765 B.n763 B.n762 163.367
R766 B.n762 B.n33 163.367
R767 B.n758 B.n33 163.367
R768 B.n758 B.n757 163.367
R769 B.n757 B.n756 163.367
R770 B.n756 B.n35 163.367
R771 B.n320 B.n187 163.367
R772 B.n324 B.n187 163.367
R773 B.n325 B.n324 163.367
R774 B.n326 B.n325 163.367
R775 B.n326 B.n185 163.367
R776 B.n330 B.n185 163.367
R777 B.n331 B.n330 163.367
R778 B.n332 B.n331 163.367
R779 B.n332 B.n183 163.367
R780 B.n336 B.n183 163.367
R781 B.n337 B.n336 163.367
R782 B.n338 B.n337 163.367
R783 B.n338 B.n181 163.367
R784 B.n342 B.n181 163.367
R785 B.n343 B.n342 163.367
R786 B.n344 B.n343 163.367
R787 B.n344 B.n179 163.367
R788 B.n348 B.n179 163.367
R789 B.n349 B.n348 163.367
R790 B.n350 B.n349 163.367
R791 B.n350 B.n177 163.367
R792 B.n354 B.n177 163.367
R793 B.n355 B.n354 163.367
R794 B.n356 B.n355 163.367
R795 B.n356 B.n175 163.367
R796 B.n360 B.n175 163.367
R797 B.n361 B.n360 163.367
R798 B.n362 B.n361 163.367
R799 B.n362 B.n173 163.367
R800 B.n366 B.n173 163.367
R801 B.n367 B.n366 163.367
R802 B.n368 B.n367 163.367
R803 B.n368 B.n169 163.367
R804 B.n373 B.n169 163.367
R805 B.n374 B.n373 163.367
R806 B.n375 B.n374 163.367
R807 B.n375 B.n167 163.367
R808 B.n379 B.n167 163.367
R809 B.n380 B.n379 163.367
R810 B.n381 B.n380 163.367
R811 B.n381 B.n165 163.367
R812 B.n385 B.n165 163.367
R813 B.n386 B.n385 163.367
R814 B.n386 B.n161 163.367
R815 B.n390 B.n161 163.367
R816 B.n391 B.n390 163.367
R817 B.n392 B.n391 163.367
R818 B.n392 B.n159 163.367
R819 B.n396 B.n159 163.367
R820 B.n397 B.n396 163.367
R821 B.n398 B.n397 163.367
R822 B.n398 B.n157 163.367
R823 B.n402 B.n157 163.367
R824 B.n403 B.n402 163.367
R825 B.n404 B.n403 163.367
R826 B.n404 B.n155 163.367
R827 B.n408 B.n155 163.367
R828 B.n409 B.n408 163.367
R829 B.n410 B.n409 163.367
R830 B.n410 B.n153 163.367
R831 B.n414 B.n153 163.367
R832 B.n415 B.n414 163.367
R833 B.n416 B.n415 163.367
R834 B.n416 B.n151 163.367
R835 B.n420 B.n151 163.367
R836 B.n421 B.n420 163.367
R837 B.n422 B.n421 163.367
R838 B.n422 B.n149 163.367
R839 B.n426 B.n149 163.367
R840 B.n427 B.n426 163.367
R841 B.n428 B.n427 163.367
R842 B.n428 B.n147 163.367
R843 B.n432 B.n147 163.367
R844 B.n433 B.n432 163.367
R845 B.n434 B.n433 163.367
R846 B.n438 B.n145 163.367
R847 B.n439 B.n438 163.367
R848 B.n440 B.n439 163.367
R849 B.n440 B.n143 163.367
R850 B.n444 B.n143 163.367
R851 B.n445 B.n444 163.367
R852 B.n446 B.n445 163.367
R853 B.n446 B.n141 163.367
R854 B.n450 B.n141 163.367
R855 B.n451 B.n450 163.367
R856 B.n452 B.n451 163.367
R857 B.n452 B.n139 163.367
R858 B.n456 B.n139 163.367
R859 B.n457 B.n456 163.367
R860 B.n458 B.n457 163.367
R861 B.n458 B.n137 163.367
R862 B.n462 B.n137 163.367
R863 B.n463 B.n462 163.367
R864 B.n464 B.n463 163.367
R865 B.n464 B.n135 163.367
R866 B.n468 B.n135 163.367
R867 B.n469 B.n468 163.367
R868 B.n470 B.n469 163.367
R869 B.n470 B.n133 163.367
R870 B.n474 B.n133 163.367
R871 B.n475 B.n474 163.367
R872 B.n476 B.n475 163.367
R873 B.n476 B.n131 163.367
R874 B.n480 B.n131 163.367
R875 B.n481 B.n480 163.367
R876 B.n482 B.n481 163.367
R877 B.n482 B.n129 163.367
R878 B.n486 B.n129 163.367
R879 B.n487 B.n486 163.367
R880 B.n488 B.n487 163.367
R881 B.n488 B.n127 163.367
R882 B.n492 B.n127 163.367
R883 B.n493 B.n492 163.367
R884 B.n494 B.n493 163.367
R885 B.n494 B.n125 163.367
R886 B.n498 B.n125 163.367
R887 B.n499 B.n498 163.367
R888 B.n500 B.n499 163.367
R889 B.n500 B.n123 163.367
R890 B.n504 B.n123 163.367
R891 B.n505 B.n504 163.367
R892 B.n506 B.n505 163.367
R893 B.n506 B.n121 163.367
R894 B.n510 B.n121 163.367
R895 B.n511 B.n510 163.367
R896 B.n512 B.n511 163.367
R897 B.n512 B.n119 163.367
R898 B.n516 B.n119 163.367
R899 B.n517 B.n516 163.367
R900 B.n518 B.n517 163.367
R901 B.n518 B.n117 163.367
R902 B.n522 B.n117 163.367
R903 B.n523 B.n522 163.367
R904 B.n524 B.n523 163.367
R905 B.n524 B.n115 163.367
R906 B.n528 B.n115 163.367
R907 B.n529 B.n528 163.367
R908 B.n530 B.n529 163.367
R909 B.n530 B.n113 163.367
R910 B.n534 B.n113 163.367
R911 B.n535 B.n534 163.367
R912 B.n536 B.n535 163.367
R913 B.n536 B.n111 163.367
R914 B.n540 B.n111 163.367
R915 B.n541 B.n540 163.367
R916 B.n542 B.n541 163.367
R917 B.n542 B.n109 163.367
R918 B.n546 B.n109 163.367
R919 B.n547 B.n546 163.367
R920 B.n548 B.n547 163.367
R921 B.n548 B.n107 163.367
R922 B.n552 B.n107 163.367
R923 B.n553 B.n552 163.367
R924 B.n554 B.n553 163.367
R925 B.n554 B.n105 163.367
R926 B.n558 B.n105 163.367
R927 B.n559 B.n558 163.367
R928 B.n560 B.n559 163.367
R929 B.n560 B.n103 163.367
R930 B.n564 B.n103 163.367
R931 B.n565 B.n564 163.367
R932 B.n566 B.n565 163.367
R933 B.n566 B.n101 163.367
R934 B.n570 B.n101 163.367
R935 B.n571 B.n570 163.367
R936 B.n572 B.n571 163.367
R937 B.n572 B.n99 163.367
R938 B.n576 B.n99 163.367
R939 B.n577 B.n576 163.367
R940 B.n578 B.n577 163.367
R941 B.n578 B.n97 163.367
R942 B.n582 B.n97 163.367
R943 B.n583 B.n582 163.367
R944 B.n584 B.n583 163.367
R945 B.n584 B.n95 163.367
R946 B.n588 B.n95 163.367
R947 B.n589 B.n588 163.367
R948 B.n590 B.n589 163.367
R949 B.n590 B.n93 163.367
R950 B.n594 B.n93 163.367
R951 B.n595 B.n594 163.367
R952 B.n596 B.n595 163.367
R953 B.n596 B.n91 163.367
R954 B.n600 B.n91 163.367
R955 B.n601 B.n600 163.367
R956 B.n602 B.n601 163.367
R957 B.n602 B.n89 163.367
R958 B.n606 B.n89 163.367
R959 B.n607 B.n606 163.367
R960 B.n608 B.n607 163.367
R961 B.n608 B.n87 163.367
R962 B.n612 B.n87 163.367
R963 B.n613 B.n612 163.367
R964 B.n614 B.n613 163.367
R965 B.n614 B.n85 163.367
R966 B.n618 B.n85 163.367
R967 B.n619 B.n618 163.367
R968 B.n620 B.n619 163.367
R969 B.n620 B.n83 163.367
R970 B.n624 B.n83 163.367
R971 B.n625 B.n624 163.367
R972 B.n626 B.n625 163.367
R973 B.n626 B.n81 163.367
R974 B.n630 B.n81 163.367
R975 B.n631 B.n630 163.367
R976 B.n632 B.n631 163.367
R977 B.n632 B.n79 163.367
R978 B.n636 B.n79 163.367
R979 B.n637 B.n636 163.367
R980 B.n752 B.n751 163.367
R981 B.n751 B.n750 163.367
R982 B.n750 B.n37 163.367
R983 B.n746 B.n37 163.367
R984 B.n746 B.n745 163.367
R985 B.n745 B.n744 163.367
R986 B.n744 B.n39 163.367
R987 B.n740 B.n39 163.367
R988 B.n740 B.n739 163.367
R989 B.n739 B.n738 163.367
R990 B.n738 B.n41 163.367
R991 B.n734 B.n41 163.367
R992 B.n734 B.n733 163.367
R993 B.n733 B.n732 163.367
R994 B.n732 B.n43 163.367
R995 B.n728 B.n43 163.367
R996 B.n728 B.n727 163.367
R997 B.n727 B.n726 163.367
R998 B.n726 B.n45 163.367
R999 B.n722 B.n45 163.367
R1000 B.n722 B.n721 163.367
R1001 B.n721 B.n720 163.367
R1002 B.n720 B.n47 163.367
R1003 B.n716 B.n47 163.367
R1004 B.n716 B.n715 163.367
R1005 B.n715 B.n714 163.367
R1006 B.n714 B.n49 163.367
R1007 B.n710 B.n49 163.367
R1008 B.n710 B.n709 163.367
R1009 B.n709 B.n708 163.367
R1010 B.n708 B.n51 163.367
R1011 B.n704 B.n51 163.367
R1012 B.n704 B.n703 163.367
R1013 B.n703 B.n55 163.367
R1014 B.n699 B.n55 163.367
R1015 B.n699 B.n698 163.367
R1016 B.n698 B.n697 163.367
R1017 B.n697 B.n57 163.367
R1018 B.n693 B.n57 163.367
R1019 B.n693 B.n692 163.367
R1020 B.n692 B.n691 163.367
R1021 B.n691 B.n59 163.367
R1022 B.n686 B.n59 163.367
R1023 B.n686 B.n685 163.367
R1024 B.n685 B.n684 163.367
R1025 B.n684 B.n63 163.367
R1026 B.n680 B.n63 163.367
R1027 B.n680 B.n679 163.367
R1028 B.n679 B.n678 163.367
R1029 B.n678 B.n65 163.367
R1030 B.n674 B.n65 163.367
R1031 B.n674 B.n673 163.367
R1032 B.n673 B.n672 163.367
R1033 B.n672 B.n67 163.367
R1034 B.n668 B.n67 163.367
R1035 B.n668 B.n667 163.367
R1036 B.n667 B.n666 163.367
R1037 B.n666 B.n69 163.367
R1038 B.n662 B.n69 163.367
R1039 B.n662 B.n661 163.367
R1040 B.n661 B.n660 163.367
R1041 B.n660 B.n71 163.367
R1042 B.n656 B.n71 163.367
R1043 B.n656 B.n655 163.367
R1044 B.n655 B.n654 163.367
R1045 B.n654 B.n73 163.367
R1046 B.n650 B.n73 163.367
R1047 B.n650 B.n649 163.367
R1048 B.n649 B.n648 163.367
R1049 B.n648 B.n75 163.367
R1050 B.n644 B.n75 163.367
R1051 B.n644 B.n643 163.367
R1052 B.n643 B.n642 163.367
R1053 B.n642 B.n77 163.367
R1054 B.n638 B.n77 163.367
R1055 B.n163 B.t10 114.047
R1056 B.n61 B.t8 114.047
R1057 B.n171 B.t1 114.037
R1058 B.n53 B.t5 114.037
R1059 B.n163 B.n162 64.5823
R1060 B.n171 B.n170 64.5823
R1061 B.n53 B.n52 64.5823
R1062 B.n61 B.n60 64.5823
R1063 B.n164 B.n163 59.5399
R1064 B.n370 B.n171 59.5399
R1065 B.n54 B.n53 59.5399
R1066 B.n688 B.n61 59.5399
R1067 B.n754 B.n753 31.3761
R1068 B.n639 B.n78 31.3761
R1069 B.n436 B.n435 31.3761
R1070 B.n321 B.n188 31.3761
R1071 B B.n855 18.0485
R1072 B.n753 B.n36 10.6151
R1073 B.n749 B.n36 10.6151
R1074 B.n749 B.n748 10.6151
R1075 B.n748 B.n747 10.6151
R1076 B.n747 B.n38 10.6151
R1077 B.n743 B.n38 10.6151
R1078 B.n743 B.n742 10.6151
R1079 B.n742 B.n741 10.6151
R1080 B.n741 B.n40 10.6151
R1081 B.n737 B.n40 10.6151
R1082 B.n737 B.n736 10.6151
R1083 B.n736 B.n735 10.6151
R1084 B.n735 B.n42 10.6151
R1085 B.n731 B.n42 10.6151
R1086 B.n731 B.n730 10.6151
R1087 B.n730 B.n729 10.6151
R1088 B.n729 B.n44 10.6151
R1089 B.n725 B.n44 10.6151
R1090 B.n725 B.n724 10.6151
R1091 B.n724 B.n723 10.6151
R1092 B.n723 B.n46 10.6151
R1093 B.n719 B.n46 10.6151
R1094 B.n719 B.n718 10.6151
R1095 B.n718 B.n717 10.6151
R1096 B.n717 B.n48 10.6151
R1097 B.n713 B.n48 10.6151
R1098 B.n713 B.n712 10.6151
R1099 B.n712 B.n711 10.6151
R1100 B.n711 B.n50 10.6151
R1101 B.n707 B.n50 10.6151
R1102 B.n707 B.n706 10.6151
R1103 B.n706 B.n705 10.6151
R1104 B.n702 B.n701 10.6151
R1105 B.n701 B.n700 10.6151
R1106 B.n700 B.n56 10.6151
R1107 B.n696 B.n56 10.6151
R1108 B.n696 B.n695 10.6151
R1109 B.n695 B.n694 10.6151
R1110 B.n694 B.n58 10.6151
R1111 B.n690 B.n58 10.6151
R1112 B.n690 B.n689 10.6151
R1113 B.n687 B.n62 10.6151
R1114 B.n683 B.n62 10.6151
R1115 B.n683 B.n682 10.6151
R1116 B.n682 B.n681 10.6151
R1117 B.n681 B.n64 10.6151
R1118 B.n677 B.n64 10.6151
R1119 B.n677 B.n676 10.6151
R1120 B.n676 B.n675 10.6151
R1121 B.n675 B.n66 10.6151
R1122 B.n671 B.n66 10.6151
R1123 B.n671 B.n670 10.6151
R1124 B.n670 B.n669 10.6151
R1125 B.n669 B.n68 10.6151
R1126 B.n665 B.n68 10.6151
R1127 B.n665 B.n664 10.6151
R1128 B.n664 B.n663 10.6151
R1129 B.n663 B.n70 10.6151
R1130 B.n659 B.n70 10.6151
R1131 B.n659 B.n658 10.6151
R1132 B.n658 B.n657 10.6151
R1133 B.n657 B.n72 10.6151
R1134 B.n653 B.n72 10.6151
R1135 B.n653 B.n652 10.6151
R1136 B.n652 B.n651 10.6151
R1137 B.n651 B.n74 10.6151
R1138 B.n647 B.n74 10.6151
R1139 B.n647 B.n646 10.6151
R1140 B.n646 B.n645 10.6151
R1141 B.n645 B.n76 10.6151
R1142 B.n641 B.n76 10.6151
R1143 B.n641 B.n640 10.6151
R1144 B.n640 B.n639 10.6151
R1145 B.n437 B.n436 10.6151
R1146 B.n437 B.n144 10.6151
R1147 B.n441 B.n144 10.6151
R1148 B.n442 B.n441 10.6151
R1149 B.n443 B.n442 10.6151
R1150 B.n443 B.n142 10.6151
R1151 B.n447 B.n142 10.6151
R1152 B.n448 B.n447 10.6151
R1153 B.n449 B.n448 10.6151
R1154 B.n449 B.n140 10.6151
R1155 B.n453 B.n140 10.6151
R1156 B.n454 B.n453 10.6151
R1157 B.n455 B.n454 10.6151
R1158 B.n455 B.n138 10.6151
R1159 B.n459 B.n138 10.6151
R1160 B.n460 B.n459 10.6151
R1161 B.n461 B.n460 10.6151
R1162 B.n461 B.n136 10.6151
R1163 B.n465 B.n136 10.6151
R1164 B.n466 B.n465 10.6151
R1165 B.n467 B.n466 10.6151
R1166 B.n467 B.n134 10.6151
R1167 B.n471 B.n134 10.6151
R1168 B.n472 B.n471 10.6151
R1169 B.n473 B.n472 10.6151
R1170 B.n473 B.n132 10.6151
R1171 B.n477 B.n132 10.6151
R1172 B.n478 B.n477 10.6151
R1173 B.n479 B.n478 10.6151
R1174 B.n479 B.n130 10.6151
R1175 B.n483 B.n130 10.6151
R1176 B.n484 B.n483 10.6151
R1177 B.n485 B.n484 10.6151
R1178 B.n485 B.n128 10.6151
R1179 B.n489 B.n128 10.6151
R1180 B.n490 B.n489 10.6151
R1181 B.n491 B.n490 10.6151
R1182 B.n491 B.n126 10.6151
R1183 B.n495 B.n126 10.6151
R1184 B.n496 B.n495 10.6151
R1185 B.n497 B.n496 10.6151
R1186 B.n497 B.n124 10.6151
R1187 B.n501 B.n124 10.6151
R1188 B.n502 B.n501 10.6151
R1189 B.n503 B.n502 10.6151
R1190 B.n503 B.n122 10.6151
R1191 B.n507 B.n122 10.6151
R1192 B.n508 B.n507 10.6151
R1193 B.n509 B.n508 10.6151
R1194 B.n509 B.n120 10.6151
R1195 B.n513 B.n120 10.6151
R1196 B.n514 B.n513 10.6151
R1197 B.n515 B.n514 10.6151
R1198 B.n515 B.n118 10.6151
R1199 B.n519 B.n118 10.6151
R1200 B.n520 B.n519 10.6151
R1201 B.n521 B.n520 10.6151
R1202 B.n521 B.n116 10.6151
R1203 B.n525 B.n116 10.6151
R1204 B.n526 B.n525 10.6151
R1205 B.n527 B.n526 10.6151
R1206 B.n527 B.n114 10.6151
R1207 B.n531 B.n114 10.6151
R1208 B.n532 B.n531 10.6151
R1209 B.n533 B.n532 10.6151
R1210 B.n533 B.n112 10.6151
R1211 B.n537 B.n112 10.6151
R1212 B.n538 B.n537 10.6151
R1213 B.n539 B.n538 10.6151
R1214 B.n539 B.n110 10.6151
R1215 B.n543 B.n110 10.6151
R1216 B.n544 B.n543 10.6151
R1217 B.n545 B.n544 10.6151
R1218 B.n545 B.n108 10.6151
R1219 B.n549 B.n108 10.6151
R1220 B.n550 B.n549 10.6151
R1221 B.n551 B.n550 10.6151
R1222 B.n551 B.n106 10.6151
R1223 B.n555 B.n106 10.6151
R1224 B.n556 B.n555 10.6151
R1225 B.n557 B.n556 10.6151
R1226 B.n557 B.n104 10.6151
R1227 B.n561 B.n104 10.6151
R1228 B.n562 B.n561 10.6151
R1229 B.n563 B.n562 10.6151
R1230 B.n563 B.n102 10.6151
R1231 B.n567 B.n102 10.6151
R1232 B.n568 B.n567 10.6151
R1233 B.n569 B.n568 10.6151
R1234 B.n569 B.n100 10.6151
R1235 B.n573 B.n100 10.6151
R1236 B.n574 B.n573 10.6151
R1237 B.n575 B.n574 10.6151
R1238 B.n575 B.n98 10.6151
R1239 B.n579 B.n98 10.6151
R1240 B.n580 B.n579 10.6151
R1241 B.n581 B.n580 10.6151
R1242 B.n581 B.n96 10.6151
R1243 B.n585 B.n96 10.6151
R1244 B.n586 B.n585 10.6151
R1245 B.n587 B.n586 10.6151
R1246 B.n587 B.n94 10.6151
R1247 B.n591 B.n94 10.6151
R1248 B.n592 B.n591 10.6151
R1249 B.n593 B.n592 10.6151
R1250 B.n593 B.n92 10.6151
R1251 B.n597 B.n92 10.6151
R1252 B.n598 B.n597 10.6151
R1253 B.n599 B.n598 10.6151
R1254 B.n599 B.n90 10.6151
R1255 B.n603 B.n90 10.6151
R1256 B.n604 B.n603 10.6151
R1257 B.n605 B.n604 10.6151
R1258 B.n605 B.n88 10.6151
R1259 B.n609 B.n88 10.6151
R1260 B.n610 B.n609 10.6151
R1261 B.n611 B.n610 10.6151
R1262 B.n611 B.n86 10.6151
R1263 B.n615 B.n86 10.6151
R1264 B.n616 B.n615 10.6151
R1265 B.n617 B.n616 10.6151
R1266 B.n617 B.n84 10.6151
R1267 B.n621 B.n84 10.6151
R1268 B.n622 B.n621 10.6151
R1269 B.n623 B.n622 10.6151
R1270 B.n623 B.n82 10.6151
R1271 B.n627 B.n82 10.6151
R1272 B.n628 B.n627 10.6151
R1273 B.n629 B.n628 10.6151
R1274 B.n629 B.n80 10.6151
R1275 B.n633 B.n80 10.6151
R1276 B.n634 B.n633 10.6151
R1277 B.n635 B.n634 10.6151
R1278 B.n635 B.n78 10.6151
R1279 B.n322 B.n321 10.6151
R1280 B.n323 B.n322 10.6151
R1281 B.n323 B.n186 10.6151
R1282 B.n327 B.n186 10.6151
R1283 B.n328 B.n327 10.6151
R1284 B.n329 B.n328 10.6151
R1285 B.n329 B.n184 10.6151
R1286 B.n333 B.n184 10.6151
R1287 B.n334 B.n333 10.6151
R1288 B.n335 B.n334 10.6151
R1289 B.n335 B.n182 10.6151
R1290 B.n339 B.n182 10.6151
R1291 B.n340 B.n339 10.6151
R1292 B.n341 B.n340 10.6151
R1293 B.n341 B.n180 10.6151
R1294 B.n345 B.n180 10.6151
R1295 B.n346 B.n345 10.6151
R1296 B.n347 B.n346 10.6151
R1297 B.n347 B.n178 10.6151
R1298 B.n351 B.n178 10.6151
R1299 B.n352 B.n351 10.6151
R1300 B.n353 B.n352 10.6151
R1301 B.n353 B.n176 10.6151
R1302 B.n357 B.n176 10.6151
R1303 B.n358 B.n357 10.6151
R1304 B.n359 B.n358 10.6151
R1305 B.n359 B.n174 10.6151
R1306 B.n363 B.n174 10.6151
R1307 B.n364 B.n363 10.6151
R1308 B.n365 B.n364 10.6151
R1309 B.n365 B.n172 10.6151
R1310 B.n369 B.n172 10.6151
R1311 B.n372 B.n371 10.6151
R1312 B.n372 B.n168 10.6151
R1313 B.n376 B.n168 10.6151
R1314 B.n377 B.n376 10.6151
R1315 B.n378 B.n377 10.6151
R1316 B.n378 B.n166 10.6151
R1317 B.n382 B.n166 10.6151
R1318 B.n383 B.n382 10.6151
R1319 B.n384 B.n383 10.6151
R1320 B.n388 B.n387 10.6151
R1321 B.n389 B.n388 10.6151
R1322 B.n389 B.n160 10.6151
R1323 B.n393 B.n160 10.6151
R1324 B.n394 B.n393 10.6151
R1325 B.n395 B.n394 10.6151
R1326 B.n395 B.n158 10.6151
R1327 B.n399 B.n158 10.6151
R1328 B.n400 B.n399 10.6151
R1329 B.n401 B.n400 10.6151
R1330 B.n401 B.n156 10.6151
R1331 B.n405 B.n156 10.6151
R1332 B.n406 B.n405 10.6151
R1333 B.n407 B.n406 10.6151
R1334 B.n407 B.n154 10.6151
R1335 B.n411 B.n154 10.6151
R1336 B.n412 B.n411 10.6151
R1337 B.n413 B.n412 10.6151
R1338 B.n413 B.n152 10.6151
R1339 B.n417 B.n152 10.6151
R1340 B.n418 B.n417 10.6151
R1341 B.n419 B.n418 10.6151
R1342 B.n419 B.n150 10.6151
R1343 B.n423 B.n150 10.6151
R1344 B.n424 B.n423 10.6151
R1345 B.n425 B.n424 10.6151
R1346 B.n425 B.n148 10.6151
R1347 B.n429 B.n148 10.6151
R1348 B.n430 B.n429 10.6151
R1349 B.n431 B.n430 10.6151
R1350 B.n431 B.n146 10.6151
R1351 B.n435 B.n146 10.6151
R1352 B.n317 B.n188 10.6151
R1353 B.n317 B.n316 10.6151
R1354 B.n316 B.n315 10.6151
R1355 B.n315 B.n190 10.6151
R1356 B.n311 B.n190 10.6151
R1357 B.n311 B.n310 10.6151
R1358 B.n310 B.n309 10.6151
R1359 B.n309 B.n192 10.6151
R1360 B.n305 B.n192 10.6151
R1361 B.n305 B.n304 10.6151
R1362 B.n304 B.n303 10.6151
R1363 B.n303 B.n194 10.6151
R1364 B.n299 B.n194 10.6151
R1365 B.n299 B.n298 10.6151
R1366 B.n298 B.n297 10.6151
R1367 B.n297 B.n196 10.6151
R1368 B.n293 B.n196 10.6151
R1369 B.n293 B.n292 10.6151
R1370 B.n292 B.n291 10.6151
R1371 B.n291 B.n198 10.6151
R1372 B.n287 B.n198 10.6151
R1373 B.n287 B.n286 10.6151
R1374 B.n286 B.n285 10.6151
R1375 B.n285 B.n200 10.6151
R1376 B.n281 B.n200 10.6151
R1377 B.n281 B.n280 10.6151
R1378 B.n280 B.n279 10.6151
R1379 B.n279 B.n202 10.6151
R1380 B.n275 B.n202 10.6151
R1381 B.n275 B.n274 10.6151
R1382 B.n274 B.n273 10.6151
R1383 B.n273 B.n204 10.6151
R1384 B.n269 B.n204 10.6151
R1385 B.n269 B.n268 10.6151
R1386 B.n268 B.n267 10.6151
R1387 B.n267 B.n206 10.6151
R1388 B.n263 B.n206 10.6151
R1389 B.n263 B.n262 10.6151
R1390 B.n262 B.n261 10.6151
R1391 B.n261 B.n208 10.6151
R1392 B.n257 B.n208 10.6151
R1393 B.n257 B.n256 10.6151
R1394 B.n256 B.n255 10.6151
R1395 B.n255 B.n210 10.6151
R1396 B.n251 B.n210 10.6151
R1397 B.n251 B.n250 10.6151
R1398 B.n250 B.n249 10.6151
R1399 B.n249 B.n212 10.6151
R1400 B.n245 B.n212 10.6151
R1401 B.n245 B.n244 10.6151
R1402 B.n244 B.n243 10.6151
R1403 B.n243 B.n214 10.6151
R1404 B.n239 B.n214 10.6151
R1405 B.n239 B.n238 10.6151
R1406 B.n238 B.n237 10.6151
R1407 B.n237 B.n216 10.6151
R1408 B.n233 B.n216 10.6151
R1409 B.n233 B.n232 10.6151
R1410 B.n232 B.n231 10.6151
R1411 B.n231 B.n218 10.6151
R1412 B.n227 B.n218 10.6151
R1413 B.n227 B.n226 10.6151
R1414 B.n226 B.n225 10.6151
R1415 B.n225 B.n220 10.6151
R1416 B.n221 B.n220 10.6151
R1417 B.n221 B.n0 10.6151
R1418 B.n851 B.n1 10.6151
R1419 B.n851 B.n850 10.6151
R1420 B.n850 B.n849 10.6151
R1421 B.n849 B.n4 10.6151
R1422 B.n845 B.n4 10.6151
R1423 B.n845 B.n844 10.6151
R1424 B.n844 B.n843 10.6151
R1425 B.n843 B.n6 10.6151
R1426 B.n839 B.n6 10.6151
R1427 B.n839 B.n838 10.6151
R1428 B.n838 B.n837 10.6151
R1429 B.n837 B.n8 10.6151
R1430 B.n833 B.n8 10.6151
R1431 B.n833 B.n832 10.6151
R1432 B.n832 B.n831 10.6151
R1433 B.n831 B.n10 10.6151
R1434 B.n827 B.n10 10.6151
R1435 B.n827 B.n826 10.6151
R1436 B.n826 B.n825 10.6151
R1437 B.n825 B.n12 10.6151
R1438 B.n821 B.n12 10.6151
R1439 B.n821 B.n820 10.6151
R1440 B.n820 B.n819 10.6151
R1441 B.n819 B.n14 10.6151
R1442 B.n815 B.n14 10.6151
R1443 B.n815 B.n814 10.6151
R1444 B.n814 B.n813 10.6151
R1445 B.n813 B.n16 10.6151
R1446 B.n809 B.n16 10.6151
R1447 B.n809 B.n808 10.6151
R1448 B.n808 B.n807 10.6151
R1449 B.n807 B.n18 10.6151
R1450 B.n803 B.n18 10.6151
R1451 B.n803 B.n802 10.6151
R1452 B.n802 B.n801 10.6151
R1453 B.n801 B.n20 10.6151
R1454 B.n797 B.n20 10.6151
R1455 B.n797 B.n796 10.6151
R1456 B.n796 B.n795 10.6151
R1457 B.n795 B.n22 10.6151
R1458 B.n791 B.n22 10.6151
R1459 B.n791 B.n790 10.6151
R1460 B.n790 B.n789 10.6151
R1461 B.n789 B.n24 10.6151
R1462 B.n785 B.n24 10.6151
R1463 B.n785 B.n784 10.6151
R1464 B.n784 B.n783 10.6151
R1465 B.n783 B.n26 10.6151
R1466 B.n779 B.n26 10.6151
R1467 B.n779 B.n778 10.6151
R1468 B.n778 B.n777 10.6151
R1469 B.n777 B.n28 10.6151
R1470 B.n773 B.n28 10.6151
R1471 B.n773 B.n772 10.6151
R1472 B.n772 B.n771 10.6151
R1473 B.n771 B.n30 10.6151
R1474 B.n767 B.n30 10.6151
R1475 B.n767 B.n766 10.6151
R1476 B.n766 B.n765 10.6151
R1477 B.n765 B.n32 10.6151
R1478 B.n761 B.n32 10.6151
R1479 B.n761 B.n760 10.6151
R1480 B.n760 B.n759 10.6151
R1481 B.n759 B.n34 10.6151
R1482 B.n755 B.n34 10.6151
R1483 B.n755 B.n754 10.6151
R1484 B.n705 B.n54 9.36635
R1485 B.n688 B.n687 9.36635
R1486 B.n370 B.n369 9.36635
R1487 B.n387 B.n164 9.36635
R1488 B.n855 B.n0 2.81026
R1489 B.n855 B.n1 2.81026
R1490 B.n702 B.n54 1.24928
R1491 B.n689 B.n688 1.24928
R1492 B.n371 B.n370 1.24928
R1493 B.n384 B.n164 1.24928
R1494 VP.n27 VP.n24 161.3
R1495 VP.n29 VP.n28 161.3
R1496 VP.n30 VP.n23 161.3
R1497 VP.n32 VP.n31 161.3
R1498 VP.n33 VP.n22 161.3
R1499 VP.n35 VP.n34 161.3
R1500 VP.n36 VP.n21 161.3
R1501 VP.n39 VP.n38 161.3
R1502 VP.n40 VP.n20 161.3
R1503 VP.n42 VP.n41 161.3
R1504 VP.n43 VP.n19 161.3
R1505 VP.n45 VP.n44 161.3
R1506 VP.n46 VP.n18 161.3
R1507 VP.n48 VP.n47 161.3
R1508 VP.n50 VP.n17 161.3
R1509 VP.n52 VP.n51 161.3
R1510 VP.n53 VP.n16 161.3
R1511 VP.n55 VP.n54 161.3
R1512 VP.n56 VP.n15 161.3
R1513 VP.n58 VP.n57 161.3
R1514 VP.n103 VP.n102 161.3
R1515 VP.n101 VP.n1 161.3
R1516 VP.n100 VP.n99 161.3
R1517 VP.n98 VP.n2 161.3
R1518 VP.n97 VP.n96 161.3
R1519 VP.n95 VP.n3 161.3
R1520 VP.n93 VP.n92 161.3
R1521 VP.n91 VP.n4 161.3
R1522 VP.n90 VP.n89 161.3
R1523 VP.n88 VP.n5 161.3
R1524 VP.n87 VP.n86 161.3
R1525 VP.n85 VP.n6 161.3
R1526 VP.n84 VP.n83 161.3
R1527 VP.n81 VP.n7 161.3
R1528 VP.n80 VP.n79 161.3
R1529 VP.n78 VP.n8 161.3
R1530 VP.n77 VP.n76 161.3
R1531 VP.n75 VP.n9 161.3
R1532 VP.n74 VP.n73 161.3
R1533 VP.n72 VP.n10 161.3
R1534 VP.n71 VP.n70 161.3
R1535 VP.n68 VP.n11 161.3
R1536 VP.n67 VP.n66 161.3
R1537 VP.n65 VP.n12 161.3
R1538 VP.n64 VP.n63 161.3
R1539 VP.n62 VP.n13 161.3
R1540 VP.n26 VP.t3 105.207
R1541 VP.n61 VP.t1 73.5055
R1542 VP.n69 VP.t6 73.5055
R1543 VP.n82 VP.t5 73.5055
R1544 VP.n94 VP.t9 73.5055
R1545 VP.n0 VP.t0 73.5055
R1546 VP.n14 VP.t4 73.5055
R1547 VP.n49 VP.t7 73.5055
R1548 VP.n37 VP.t8 73.5055
R1549 VP.n25 VP.t2 73.5055
R1550 VP.n61 VP.n60 70.0045
R1551 VP.n104 VP.n0 70.0045
R1552 VP.n59 VP.n14 70.0045
R1553 VP.n26 VP.n25 69.7461
R1554 VP.n67 VP.n12 56.5193
R1555 VP.n100 VP.n2 56.5193
R1556 VP.n55 VP.n16 56.5193
R1557 VP.n60 VP.n59 53.2531
R1558 VP.n76 VP.n8 48.7492
R1559 VP.n88 VP.n87 48.7492
R1560 VP.n43 VP.n42 48.7492
R1561 VP.n31 VP.n22 48.7492
R1562 VP.n76 VP.n75 32.2376
R1563 VP.n89 VP.n88 32.2376
R1564 VP.n44 VP.n43 32.2376
R1565 VP.n31 VP.n30 32.2376
R1566 VP.n63 VP.n62 24.4675
R1567 VP.n63 VP.n12 24.4675
R1568 VP.n68 VP.n67 24.4675
R1569 VP.n70 VP.n68 24.4675
R1570 VP.n74 VP.n10 24.4675
R1571 VP.n75 VP.n74 24.4675
R1572 VP.n80 VP.n8 24.4675
R1573 VP.n81 VP.n80 24.4675
R1574 VP.n83 VP.n6 24.4675
R1575 VP.n87 VP.n6 24.4675
R1576 VP.n89 VP.n4 24.4675
R1577 VP.n93 VP.n4 24.4675
R1578 VP.n96 VP.n95 24.4675
R1579 VP.n96 VP.n2 24.4675
R1580 VP.n101 VP.n100 24.4675
R1581 VP.n102 VP.n101 24.4675
R1582 VP.n56 VP.n55 24.4675
R1583 VP.n57 VP.n56 24.4675
R1584 VP.n44 VP.n18 24.4675
R1585 VP.n48 VP.n18 24.4675
R1586 VP.n51 VP.n50 24.4675
R1587 VP.n51 VP.n16 24.4675
R1588 VP.n35 VP.n22 24.4675
R1589 VP.n36 VP.n35 24.4675
R1590 VP.n38 VP.n20 24.4675
R1591 VP.n42 VP.n20 24.4675
R1592 VP.n29 VP.n24 24.4675
R1593 VP.n30 VP.n29 24.4675
R1594 VP.n70 VP.n69 20.5528
R1595 VP.n95 VP.n94 20.5528
R1596 VP.n50 VP.n49 20.5528
R1597 VP.n62 VP.n61 20.0634
R1598 VP.n102 VP.n0 20.0634
R1599 VP.n57 VP.n14 20.0634
R1600 VP.n82 VP.n81 12.234
R1601 VP.n83 VP.n82 12.234
R1602 VP.n37 VP.n36 12.234
R1603 VP.n38 VP.n37 12.234
R1604 VP.n27 VP.n26 5.54913
R1605 VP.n69 VP.n10 3.91522
R1606 VP.n94 VP.n93 3.91522
R1607 VP.n49 VP.n48 3.91522
R1608 VP.n25 VP.n24 3.91522
R1609 VP.n59 VP.n58 0.354971
R1610 VP.n60 VP.n13 0.354971
R1611 VP.n104 VP.n103 0.354971
R1612 VP VP.n104 0.26696
R1613 VP.n28 VP.n27 0.189894
R1614 VP.n28 VP.n23 0.189894
R1615 VP.n32 VP.n23 0.189894
R1616 VP.n33 VP.n32 0.189894
R1617 VP.n34 VP.n33 0.189894
R1618 VP.n34 VP.n21 0.189894
R1619 VP.n39 VP.n21 0.189894
R1620 VP.n40 VP.n39 0.189894
R1621 VP.n41 VP.n40 0.189894
R1622 VP.n41 VP.n19 0.189894
R1623 VP.n45 VP.n19 0.189894
R1624 VP.n46 VP.n45 0.189894
R1625 VP.n47 VP.n46 0.189894
R1626 VP.n47 VP.n17 0.189894
R1627 VP.n52 VP.n17 0.189894
R1628 VP.n53 VP.n52 0.189894
R1629 VP.n54 VP.n53 0.189894
R1630 VP.n54 VP.n15 0.189894
R1631 VP.n58 VP.n15 0.189894
R1632 VP.n64 VP.n13 0.189894
R1633 VP.n65 VP.n64 0.189894
R1634 VP.n66 VP.n65 0.189894
R1635 VP.n66 VP.n11 0.189894
R1636 VP.n71 VP.n11 0.189894
R1637 VP.n72 VP.n71 0.189894
R1638 VP.n73 VP.n72 0.189894
R1639 VP.n73 VP.n9 0.189894
R1640 VP.n77 VP.n9 0.189894
R1641 VP.n78 VP.n77 0.189894
R1642 VP.n79 VP.n78 0.189894
R1643 VP.n79 VP.n7 0.189894
R1644 VP.n84 VP.n7 0.189894
R1645 VP.n85 VP.n84 0.189894
R1646 VP.n86 VP.n85 0.189894
R1647 VP.n86 VP.n5 0.189894
R1648 VP.n90 VP.n5 0.189894
R1649 VP.n91 VP.n90 0.189894
R1650 VP.n92 VP.n91 0.189894
R1651 VP.n92 VP.n3 0.189894
R1652 VP.n97 VP.n3 0.189894
R1653 VP.n98 VP.n97 0.189894
R1654 VP.n99 VP.n98 0.189894
R1655 VP.n99 VP.n1 0.189894
R1656 VP.n103 VP.n1 0.189894
R1657 VDD1.n1 VDD1.t6 84.4748
R1658 VDD1.n3 VDD1.t8 84.4747
R1659 VDD1.n5 VDD1.n4 80.1492
R1660 VDD1.n7 VDD1.n6 78.0517
R1661 VDD1.n1 VDD1.n0 78.0517
R1662 VDD1.n3 VDD1.n2 78.0515
R1663 VDD1.n7 VDD1.n5 47.2574
R1664 VDD1.n6 VDD1.t2 3.55296
R1665 VDD1.n6 VDD1.t5 3.55296
R1666 VDD1.n0 VDD1.t7 3.55296
R1667 VDD1.n0 VDD1.t1 3.55296
R1668 VDD1.n4 VDD1.t0 3.55296
R1669 VDD1.n4 VDD1.t9 3.55296
R1670 VDD1.n2 VDD1.t3 3.55296
R1671 VDD1.n2 VDD1.t4 3.55296
R1672 VDD1 VDD1.n7 2.09533
R1673 VDD1 VDD1.n1 0.776362
R1674 VDD1.n5 VDD1.n3 0.662826
C0 B w_n4966_n2798# 10.4206f
C1 w_n4966_n2798# VDD1 2.74475f
C2 w_n4966_n2798# VP 11.3412f
C3 VN w_n4966_n2798# 10.6934f
C4 B VDD1 2.40953f
C5 B VP 2.44308f
C6 VN B 1.35159f
C7 VP VDD1 8.9553f
C8 VN VDD1 0.15429f
C9 VN VP 8.46261f
C10 VDD2 VTAIL 9.35249f
C11 VTAIL w_n4966_n2798# 2.87531f
C12 VDD2 w_n4966_n2798# 2.90909f
C13 VTAIL B 3.23628f
C14 VDD2 B 2.54302f
C15 VTAIL VDD1 9.2979f
C16 VDD2 VDD1 2.43472f
C17 VTAIL VP 9.43821f
C18 VTAIL VN 9.42399f
C19 VDD2 VP 0.63442f
C20 VDD2 VN 8.4786f
C21 VDD2 VSUBS 2.294705f
C22 VDD1 VSUBS 2.055815f
C23 VTAIL VSUBS 1.310314f
C24 VN VSUBS 8.30615f
C25 VP VSUBS 4.658065f
C26 B VSUBS 5.623429f
C27 w_n4966_n2798# VSUBS 0.171923p
C28 VDD1.t6 VSUBS 2.25993f
C29 VDD1.t7 VSUBS 0.230554f
C30 VDD1.t1 VSUBS 0.230554f
C31 VDD1.n0 VSUBS 1.68851f
C32 VDD1.n1 VSUBS 1.91258f
C33 VDD1.t8 VSUBS 2.25992f
C34 VDD1.t3 VSUBS 0.230554f
C35 VDD1.t4 VSUBS 0.230554f
C36 VDD1.n2 VSUBS 1.68851f
C37 VDD1.n3 VSUBS 1.90205f
C38 VDD1.t0 VSUBS 0.230554f
C39 VDD1.t9 VSUBS 0.230554f
C40 VDD1.n4 VSUBS 1.71756f
C41 VDD1.n5 VSUBS 4.23841f
C42 VDD1.t2 VSUBS 0.230554f
C43 VDD1.t5 VSUBS 0.230554f
C44 VDD1.n6 VSUBS 1.68851f
C45 VDD1.n7 VSUBS 4.30464f
C46 VP.t0 VSUBS 2.32592f
C47 VP.n0 VSUBS 0.957591f
C48 VP.n1 VSUBS 0.031378f
C49 VP.n2 VSUBS 0.045372f
C50 VP.n3 VSUBS 0.031378f
C51 VP.t9 VSUBS 2.32592f
C52 VP.n4 VSUBS 0.058481f
C53 VP.n5 VSUBS 0.031378f
C54 VP.n6 VSUBS 0.058481f
C55 VP.n7 VSUBS 0.031378f
C56 VP.t5 VSUBS 2.32592f
C57 VP.n8 VSUBS 0.058481f
C58 VP.n9 VSUBS 0.031378f
C59 VP.n10 VSUBS 0.034228f
C60 VP.n11 VSUBS 0.031378f
C61 VP.n12 VSUBS 0.046247f
C62 VP.n13 VSUBS 0.050644f
C63 VP.t1 VSUBS 2.32592f
C64 VP.t4 VSUBS 2.32592f
C65 VP.n14 VSUBS 0.957591f
C66 VP.n15 VSUBS 0.031378f
C67 VP.n16 VSUBS 0.045372f
C68 VP.n17 VSUBS 0.031378f
C69 VP.t7 VSUBS 2.32592f
C70 VP.n18 VSUBS 0.058481f
C71 VP.n19 VSUBS 0.031378f
C72 VP.n20 VSUBS 0.058481f
C73 VP.n21 VSUBS 0.031378f
C74 VP.t8 VSUBS 2.32592f
C75 VP.n22 VSUBS 0.058481f
C76 VP.n23 VSUBS 0.031378f
C77 VP.n24 VSUBS 0.034228f
C78 VP.t3 VSUBS 2.64032f
C79 VP.t2 VSUBS 2.32592f
C80 VP.n25 VSUBS 0.92399f
C81 VP.n26 VSUBS 0.895199f
C82 VP.n27 VSUBS 0.33935f
C83 VP.n28 VSUBS 0.031378f
C84 VP.n29 VSUBS 0.058481f
C85 VP.n30 VSUBS 0.063213f
C86 VP.n31 VSUBS 0.028406f
C87 VP.n32 VSUBS 0.031378f
C88 VP.n33 VSUBS 0.031378f
C89 VP.n34 VSUBS 0.031378f
C90 VP.n35 VSUBS 0.058481f
C91 VP.n36 VSUBS 0.044045f
C92 VP.n37 VSUBS 0.833493f
C93 VP.n38 VSUBS 0.044045f
C94 VP.n39 VSUBS 0.031378f
C95 VP.n40 VSUBS 0.031378f
C96 VP.n41 VSUBS 0.031378f
C97 VP.n42 VSUBS 0.058481f
C98 VP.n43 VSUBS 0.028406f
C99 VP.n44 VSUBS 0.063213f
C100 VP.n45 VSUBS 0.031378f
C101 VP.n46 VSUBS 0.031378f
C102 VP.n47 VSUBS 0.031378f
C103 VP.n48 VSUBS 0.034228f
C104 VP.n49 VSUBS 0.833493f
C105 VP.n50 VSUBS 0.053862f
C106 VP.n51 VSUBS 0.058481f
C107 VP.n52 VSUBS 0.031378f
C108 VP.n53 VSUBS 0.031378f
C109 VP.n54 VSUBS 0.031378f
C110 VP.n55 VSUBS 0.046247f
C111 VP.n56 VSUBS 0.058481f
C112 VP.n57 VSUBS 0.053284f
C113 VP.n58 VSUBS 0.050644f
C114 VP.n59 VSUBS 1.94042f
C115 VP.n60 VSUBS 1.9616f
C116 VP.n61 VSUBS 0.957591f
C117 VP.n62 VSUBS 0.053284f
C118 VP.n63 VSUBS 0.058481f
C119 VP.n64 VSUBS 0.031378f
C120 VP.n65 VSUBS 0.031378f
C121 VP.n66 VSUBS 0.031378f
C122 VP.n67 VSUBS 0.045372f
C123 VP.n68 VSUBS 0.058481f
C124 VP.t6 VSUBS 2.32592f
C125 VP.n69 VSUBS 0.833493f
C126 VP.n70 VSUBS 0.053862f
C127 VP.n71 VSUBS 0.031378f
C128 VP.n72 VSUBS 0.031378f
C129 VP.n73 VSUBS 0.031378f
C130 VP.n74 VSUBS 0.058481f
C131 VP.n75 VSUBS 0.063213f
C132 VP.n76 VSUBS 0.028406f
C133 VP.n77 VSUBS 0.031378f
C134 VP.n78 VSUBS 0.031378f
C135 VP.n79 VSUBS 0.031378f
C136 VP.n80 VSUBS 0.058481f
C137 VP.n81 VSUBS 0.044045f
C138 VP.n82 VSUBS 0.833493f
C139 VP.n83 VSUBS 0.044045f
C140 VP.n84 VSUBS 0.031378f
C141 VP.n85 VSUBS 0.031378f
C142 VP.n86 VSUBS 0.031378f
C143 VP.n87 VSUBS 0.058481f
C144 VP.n88 VSUBS 0.028406f
C145 VP.n89 VSUBS 0.063213f
C146 VP.n90 VSUBS 0.031378f
C147 VP.n91 VSUBS 0.031378f
C148 VP.n92 VSUBS 0.031378f
C149 VP.n93 VSUBS 0.034228f
C150 VP.n94 VSUBS 0.833493f
C151 VP.n95 VSUBS 0.053862f
C152 VP.n96 VSUBS 0.058481f
C153 VP.n97 VSUBS 0.031378f
C154 VP.n98 VSUBS 0.031378f
C155 VP.n99 VSUBS 0.031378f
C156 VP.n100 VSUBS 0.046247f
C157 VP.n101 VSUBS 0.058481f
C158 VP.n102 VSUBS 0.053284f
C159 VP.n103 VSUBS 0.050644f
C160 VP.n104 VSUBS 0.065213f
C161 B.n0 VSUBS 0.006331f
C162 B.n1 VSUBS 0.006331f
C163 B.n2 VSUBS 0.010012f
C164 B.n3 VSUBS 0.010012f
C165 B.n4 VSUBS 0.010012f
C166 B.n5 VSUBS 0.010012f
C167 B.n6 VSUBS 0.010012f
C168 B.n7 VSUBS 0.010012f
C169 B.n8 VSUBS 0.010012f
C170 B.n9 VSUBS 0.010012f
C171 B.n10 VSUBS 0.010012f
C172 B.n11 VSUBS 0.010012f
C173 B.n12 VSUBS 0.010012f
C174 B.n13 VSUBS 0.010012f
C175 B.n14 VSUBS 0.010012f
C176 B.n15 VSUBS 0.010012f
C177 B.n16 VSUBS 0.010012f
C178 B.n17 VSUBS 0.010012f
C179 B.n18 VSUBS 0.010012f
C180 B.n19 VSUBS 0.010012f
C181 B.n20 VSUBS 0.010012f
C182 B.n21 VSUBS 0.010012f
C183 B.n22 VSUBS 0.010012f
C184 B.n23 VSUBS 0.010012f
C185 B.n24 VSUBS 0.010012f
C186 B.n25 VSUBS 0.010012f
C187 B.n26 VSUBS 0.010012f
C188 B.n27 VSUBS 0.010012f
C189 B.n28 VSUBS 0.010012f
C190 B.n29 VSUBS 0.010012f
C191 B.n30 VSUBS 0.010012f
C192 B.n31 VSUBS 0.010012f
C193 B.n32 VSUBS 0.010012f
C194 B.n33 VSUBS 0.010012f
C195 B.n34 VSUBS 0.010012f
C196 B.n35 VSUBS 0.022386f
C197 B.n36 VSUBS 0.010012f
C198 B.n37 VSUBS 0.010012f
C199 B.n38 VSUBS 0.010012f
C200 B.n39 VSUBS 0.010012f
C201 B.n40 VSUBS 0.010012f
C202 B.n41 VSUBS 0.010012f
C203 B.n42 VSUBS 0.010012f
C204 B.n43 VSUBS 0.010012f
C205 B.n44 VSUBS 0.010012f
C206 B.n45 VSUBS 0.010012f
C207 B.n46 VSUBS 0.010012f
C208 B.n47 VSUBS 0.010012f
C209 B.n48 VSUBS 0.010012f
C210 B.n49 VSUBS 0.010012f
C211 B.n50 VSUBS 0.010012f
C212 B.n51 VSUBS 0.010012f
C213 B.t5 VSUBS 0.412247f
C214 B.t4 VSUBS 0.444963f
C215 B.t3 VSUBS 1.83251f
C216 B.n52 VSUBS 0.244065f
C217 B.n53 VSUBS 0.104765f
C218 B.n54 VSUBS 0.023197f
C219 B.n55 VSUBS 0.010012f
C220 B.n56 VSUBS 0.010012f
C221 B.n57 VSUBS 0.010012f
C222 B.n58 VSUBS 0.010012f
C223 B.n59 VSUBS 0.010012f
C224 B.t8 VSUBS 0.412243f
C225 B.t7 VSUBS 0.444959f
C226 B.t6 VSUBS 1.83251f
C227 B.n60 VSUBS 0.24407f
C228 B.n61 VSUBS 0.104769f
C229 B.n62 VSUBS 0.010012f
C230 B.n63 VSUBS 0.010012f
C231 B.n64 VSUBS 0.010012f
C232 B.n65 VSUBS 0.010012f
C233 B.n66 VSUBS 0.010012f
C234 B.n67 VSUBS 0.010012f
C235 B.n68 VSUBS 0.010012f
C236 B.n69 VSUBS 0.010012f
C237 B.n70 VSUBS 0.010012f
C238 B.n71 VSUBS 0.010012f
C239 B.n72 VSUBS 0.010012f
C240 B.n73 VSUBS 0.010012f
C241 B.n74 VSUBS 0.010012f
C242 B.n75 VSUBS 0.010012f
C243 B.n76 VSUBS 0.010012f
C244 B.n77 VSUBS 0.010012f
C245 B.n78 VSUBS 0.023617f
C246 B.n79 VSUBS 0.010012f
C247 B.n80 VSUBS 0.010012f
C248 B.n81 VSUBS 0.010012f
C249 B.n82 VSUBS 0.010012f
C250 B.n83 VSUBS 0.010012f
C251 B.n84 VSUBS 0.010012f
C252 B.n85 VSUBS 0.010012f
C253 B.n86 VSUBS 0.010012f
C254 B.n87 VSUBS 0.010012f
C255 B.n88 VSUBS 0.010012f
C256 B.n89 VSUBS 0.010012f
C257 B.n90 VSUBS 0.010012f
C258 B.n91 VSUBS 0.010012f
C259 B.n92 VSUBS 0.010012f
C260 B.n93 VSUBS 0.010012f
C261 B.n94 VSUBS 0.010012f
C262 B.n95 VSUBS 0.010012f
C263 B.n96 VSUBS 0.010012f
C264 B.n97 VSUBS 0.010012f
C265 B.n98 VSUBS 0.010012f
C266 B.n99 VSUBS 0.010012f
C267 B.n100 VSUBS 0.010012f
C268 B.n101 VSUBS 0.010012f
C269 B.n102 VSUBS 0.010012f
C270 B.n103 VSUBS 0.010012f
C271 B.n104 VSUBS 0.010012f
C272 B.n105 VSUBS 0.010012f
C273 B.n106 VSUBS 0.010012f
C274 B.n107 VSUBS 0.010012f
C275 B.n108 VSUBS 0.010012f
C276 B.n109 VSUBS 0.010012f
C277 B.n110 VSUBS 0.010012f
C278 B.n111 VSUBS 0.010012f
C279 B.n112 VSUBS 0.010012f
C280 B.n113 VSUBS 0.010012f
C281 B.n114 VSUBS 0.010012f
C282 B.n115 VSUBS 0.010012f
C283 B.n116 VSUBS 0.010012f
C284 B.n117 VSUBS 0.010012f
C285 B.n118 VSUBS 0.010012f
C286 B.n119 VSUBS 0.010012f
C287 B.n120 VSUBS 0.010012f
C288 B.n121 VSUBS 0.010012f
C289 B.n122 VSUBS 0.010012f
C290 B.n123 VSUBS 0.010012f
C291 B.n124 VSUBS 0.010012f
C292 B.n125 VSUBS 0.010012f
C293 B.n126 VSUBS 0.010012f
C294 B.n127 VSUBS 0.010012f
C295 B.n128 VSUBS 0.010012f
C296 B.n129 VSUBS 0.010012f
C297 B.n130 VSUBS 0.010012f
C298 B.n131 VSUBS 0.010012f
C299 B.n132 VSUBS 0.010012f
C300 B.n133 VSUBS 0.010012f
C301 B.n134 VSUBS 0.010012f
C302 B.n135 VSUBS 0.010012f
C303 B.n136 VSUBS 0.010012f
C304 B.n137 VSUBS 0.010012f
C305 B.n138 VSUBS 0.010012f
C306 B.n139 VSUBS 0.010012f
C307 B.n140 VSUBS 0.010012f
C308 B.n141 VSUBS 0.010012f
C309 B.n142 VSUBS 0.010012f
C310 B.n143 VSUBS 0.010012f
C311 B.n144 VSUBS 0.010012f
C312 B.n145 VSUBS 0.022386f
C313 B.n146 VSUBS 0.010012f
C314 B.n147 VSUBS 0.010012f
C315 B.n148 VSUBS 0.010012f
C316 B.n149 VSUBS 0.010012f
C317 B.n150 VSUBS 0.010012f
C318 B.n151 VSUBS 0.010012f
C319 B.n152 VSUBS 0.010012f
C320 B.n153 VSUBS 0.010012f
C321 B.n154 VSUBS 0.010012f
C322 B.n155 VSUBS 0.010012f
C323 B.n156 VSUBS 0.010012f
C324 B.n157 VSUBS 0.010012f
C325 B.n158 VSUBS 0.010012f
C326 B.n159 VSUBS 0.010012f
C327 B.n160 VSUBS 0.010012f
C328 B.n161 VSUBS 0.010012f
C329 B.t10 VSUBS 0.412243f
C330 B.t11 VSUBS 0.444959f
C331 B.t9 VSUBS 1.83251f
C332 B.n162 VSUBS 0.24407f
C333 B.n163 VSUBS 0.104769f
C334 B.n164 VSUBS 0.023197f
C335 B.n165 VSUBS 0.010012f
C336 B.n166 VSUBS 0.010012f
C337 B.n167 VSUBS 0.010012f
C338 B.n168 VSUBS 0.010012f
C339 B.n169 VSUBS 0.010012f
C340 B.t1 VSUBS 0.412247f
C341 B.t2 VSUBS 0.444963f
C342 B.t0 VSUBS 1.83251f
C343 B.n170 VSUBS 0.244065f
C344 B.n171 VSUBS 0.104765f
C345 B.n172 VSUBS 0.010012f
C346 B.n173 VSUBS 0.010012f
C347 B.n174 VSUBS 0.010012f
C348 B.n175 VSUBS 0.010012f
C349 B.n176 VSUBS 0.010012f
C350 B.n177 VSUBS 0.010012f
C351 B.n178 VSUBS 0.010012f
C352 B.n179 VSUBS 0.010012f
C353 B.n180 VSUBS 0.010012f
C354 B.n181 VSUBS 0.010012f
C355 B.n182 VSUBS 0.010012f
C356 B.n183 VSUBS 0.010012f
C357 B.n184 VSUBS 0.010012f
C358 B.n185 VSUBS 0.010012f
C359 B.n186 VSUBS 0.010012f
C360 B.n187 VSUBS 0.010012f
C361 B.n188 VSUBS 0.022386f
C362 B.n189 VSUBS 0.010012f
C363 B.n190 VSUBS 0.010012f
C364 B.n191 VSUBS 0.010012f
C365 B.n192 VSUBS 0.010012f
C366 B.n193 VSUBS 0.010012f
C367 B.n194 VSUBS 0.010012f
C368 B.n195 VSUBS 0.010012f
C369 B.n196 VSUBS 0.010012f
C370 B.n197 VSUBS 0.010012f
C371 B.n198 VSUBS 0.010012f
C372 B.n199 VSUBS 0.010012f
C373 B.n200 VSUBS 0.010012f
C374 B.n201 VSUBS 0.010012f
C375 B.n202 VSUBS 0.010012f
C376 B.n203 VSUBS 0.010012f
C377 B.n204 VSUBS 0.010012f
C378 B.n205 VSUBS 0.010012f
C379 B.n206 VSUBS 0.010012f
C380 B.n207 VSUBS 0.010012f
C381 B.n208 VSUBS 0.010012f
C382 B.n209 VSUBS 0.010012f
C383 B.n210 VSUBS 0.010012f
C384 B.n211 VSUBS 0.010012f
C385 B.n212 VSUBS 0.010012f
C386 B.n213 VSUBS 0.010012f
C387 B.n214 VSUBS 0.010012f
C388 B.n215 VSUBS 0.010012f
C389 B.n216 VSUBS 0.010012f
C390 B.n217 VSUBS 0.010012f
C391 B.n218 VSUBS 0.010012f
C392 B.n219 VSUBS 0.010012f
C393 B.n220 VSUBS 0.010012f
C394 B.n221 VSUBS 0.010012f
C395 B.n222 VSUBS 0.010012f
C396 B.n223 VSUBS 0.010012f
C397 B.n224 VSUBS 0.010012f
C398 B.n225 VSUBS 0.010012f
C399 B.n226 VSUBS 0.010012f
C400 B.n227 VSUBS 0.010012f
C401 B.n228 VSUBS 0.010012f
C402 B.n229 VSUBS 0.010012f
C403 B.n230 VSUBS 0.010012f
C404 B.n231 VSUBS 0.010012f
C405 B.n232 VSUBS 0.010012f
C406 B.n233 VSUBS 0.010012f
C407 B.n234 VSUBS 0.010012f
C408 B.n235 VSUBS 0.010012f
C409 B.n236 VSUBS 0.010012f
C410 B.n237 VSUBS 0.010012f
C411 B.n238 VSUBS 0.010012f
C412 B.n239 VSUBS 0.010012f
C413 B.n240 VSUBS 0.010012f
C414 B.n241 VSUBS 0.010012f
C415 B.n242 VSUBS 0.010012f
C416 B.n243 VSUBS 0.010012f
C417 B.n244 VSUBS 0.010012f
C418 B.n245 VSUBS 0.010012f
C419 B.n246 VSUBS 0.010012f
C420 B.n247 VSUBS 0.010012f
C421 B.n248 VSUBS 0.010012f
C422 B.n249 VSUBS 0.010012f
C423 B.n250 VSUBS 0.010012f
C424 B.n251 VSUBS 0.010012f
C425 B.n252 VSUBS 0.010012f
C426 B.n253 VSUBS 0.010012f
C427 B.n254 VSUBS 0.010012f
C428 B.n255 VSUBS 0.010012f
C429 B.n256 VSUBS 0.010012f
C430 B.n257 VSUBS 0.010012f
C431 B.n258 VSUBS 0.010012f
C432 B.n259 VSUBS 0.010012f
C433 B.n260 VSUBS 0.010012f
C434 B.n261 VSUBS 0.010012f
C435 B.n262 VSUBS 0.010012f
C436 B.n263 VSUBS 0.010012f
C437 B.n264 VSUBS 0.010012f
C438 B.n265 VSUBS 0.010012f
C439 B.n266 VSUBS 0.010012f
C440 B.n267 VSUBS 0.010012f
C441 B.n268 VSUBS 0.010012f
C442 B.n269 VSUBS 0.010012f
C443 B.n270 VSUBS 0.010012f
C444 B.n271 VSUBS 0.010012f
C445 B.n272 VSUBS 0.010012f
C446 B.n273 VSUBS 0.010012f
C447 B.n274 VSUBS 0.010012f
C448 B.n275 VSUBS 0.010012f
C449 B.n276 VSUBS 0.010012f
C450 B.n277 VSUBS 0.010012f
C451 B.n278 VSUBS 0.010012f
C452 B.n279 VSUBS 0.010012f
C453 B.n280 VSUBS 0.010012f
C454 B.n281 VSUBS 0.010012f
C455 B.n282 VSUBS 0.010012f
C456 B.n283 VSUBS 0.010012f
C457 B.n284 VSUBS 0.010012f
C458 B.n285 VSUBS 0.010012f
C459 B.n286 VSUBS 0.010012f
C460 B.n287 VSUBS 0.010012f
C461 B.n288 VSUBS 0.010012f
C462 B.n289 VSUBS 0.010012f
C463 B.n290 VSUBS 0.010012f
C464 B.n291 VSUBS 0.010012f
C465 B.n292 VSUBS 0.010012f
C466 B.n293 VSUBS 0.010012f
C467 B.n294 VSUBS 0.010012f
C468 B.n295 VSUBS 0.010012f
C469 B.n296 VSUBS 0.010012f
C470 B.n297 VSUBS 0.010012f
C471 B.n298 VSUBS 0.010012f
C472 B.n299 VSUBS 0.010012f
C473 B.n300 VSUBS 0.010012f
C474 B.n301 VSUBS 0.010012f
C475 B.n302 VSUBS 0.010012f
C476 B.n303 VSUBS 0.010012f
C477 B.n304 VSUBS 0.010012f
C478 B.n305 VSUBS 0.010012f
C479 B.n306 VSUBS 0.010012f
C480 B.n307 VSUBS 0.010012f
C481 B.n308 VSUBS 0.010012f
C482 B.n309 VSUBS 0.010012f
C483 B.n310 VSUBS 0.010012f
C484 B.n311 VSUBS 0.010012f
C485 B.n312 VSUBS 0.010012f
C486 B.n313 VSUBS 0.010012f
C487 B.n314 VSUBS 0.010012f
C488 B.n315 VSUBS 0.010012f
C489 B.n316 VSUBS 0.010012f
C490 B.n317 VSUBS 0.010012f
C491 B.n318 VSUBS 0.010012f
C492 B.n319 VSUBS 0.022386f
C493 B.n320 VSUBS 0.023257f
C494 B.n321 VSUBS 0.023257f
C495 B.n322 VSUBS 0.010012f
C496 B.n323 VSUBS 0.010012f
C497 B.n324 VSUBS 0.010012f
C498 B.n325 VSUBS 0.010012f
C499 B.n326 VSUBS 0.010012f
C500 B.n327 VSUBS 0.010012f
C501 B.n328 VSUBS 0.010012f
C502 B.n329 VSUBS 0.010012f
C503 B.n330 VSUBS 0.010012f
C504 B.n331 VSUBS 0.010012f
C505 B.n332 VSUBS 0.010012f
C506 B.n333 VSUBS 0.010012f
C507 B.n334 VSUBS 0.010012f
C508 B.n335 VSUBS 0.010012f
C509 B.n336 VSUBS 0.010012f
C510 B.n337 VSUBS 0.010012f
C511 B.n338 VSUBS 0.010012f
C512 B.n339 VSUBS 0.010012f
C513 B.n340 VSUBS 0.010012f
C514 B.n341 VSUBS 0.010012f
C515 B.n342 VSUBS 0.010012f
C516 B.n343 VSUBS 0.010012f
C517 B.n344 VSUBS 0.010012f
C518 B.n345 VSUBS 0.010012f
C519 B.n346 VSUBS 0.010012f
C520 B.n347 VSUBS 0.010012f
C521 B.n348 VSUBS 0.010012f
C522 B.n349 VSUBS 0.010012f
C523 B.n350 VSUBS 0.010012f
C524 B.n351 VSUBS 0.010012f
C525 B.n352 VSUBS 0.010012f
C526 B.n353 VSUBS 0.010012f
C527 B.n354 VSUBS 0.010012f
C528 B.n355 VSUBS 0.010012f
C529 B.n356 VSUBS 0.010012f
C530 B.n357 VSUBS 0.010012f
C531 B.n358 VSUBS 0.010012f
C532 B.n359 VSUBS 0.010012f
C533 B.n360 VSUBS 0.010012f
C534 B.n361 VSUBS 0.010012f
C535 B.n362 VSUBS 0.010012f
C536 B.n363 VSUBS 0.010012f
C537 B.n364 VSUBS 0.010012f
C538 B.n365 VSUBS 0.010012f
C539 B.n366 VSUBS 0.010012f
C540 B.n367 VSUBS 0.010012f
C541 B.n368 VSUBS 0.010012f
C542 B.n369 VSUBS 0.009423f
C543 B.n370 VSUBS 0.023197f
C544 B.n371 VSUBS 0.005595f
C545 B.n372 VSUBS 0.010012f
C546 B.n373 VSUBS 0.010012f
C547 B.n374 VSUBS 0.010012f
C548 B.n375 VSUBS 0.010012f
C549 B.n376 VSUBS 0.010012f
C550 B.n377 VSUBS 0.010012f
C551 B.n378 VSUBS 0.010012f
C552 B.n379 VSUBS 0.010012f
C553 B.n380 VSUBS 0.010012f
C554 B.n381 VSUBS 0.010012f
C555 B.n382 VSUBS 0.010012f
C556 B.n383 VSUBS 0.010012f
C557 B.n384 VSUBS 0.005595f
C558 B.n385 VSUBS 0.010012f
C559 B.n386 VSUBS 0.010012f
C560 B.n387 VSUBS 0.009423f
C561 B.n388 VSUBS 0.010012f
C562 B.n389 VSUBS 0.010012f
C563 B.n390 VSUBS 0.010012f
C564 B.n391 VSUBS 0.010012f
C565 B.n392 VSUBS 0.010012f
C566 B.n393 VSUBS 0.010012f
C567 B.n394 VSUBS 0.010012f
C568 B.n395 VSUBS 0.010012f
C569 B.n396 VSUBS 0.010012f
C570 B.n397 VSUBS 0.010012f
C571 B.n398 VSUBS 0.010012f
C572 B.n399 VSUBS 0.010012f
C573 B.n400 VSUBS 0.010012f
C574 B.n401 VSUBS 0.010012f
C575 B.n402 VSUBS 0.010012f
C576 B.n403 VSUBS 0.010012f
C577 B.n404 VSUBS 0.010012f
C578 B.n405 VSUBS 0.010012f
C579 B.n406 VSUBS 0.010012f
C580 B.n407 VSUBS 0.010012f
C581 B.n408 VSUBS 0.010012f
C582 B.n409 VSUBS 0.010012f
C583 B.n410 VSUBS 0.010012f
C584 B.n411 VSUBS 0.010012f
C585 B.n412 VSUBS 0.010012f
C586 B.n413 VSUBS 0.010012f
C587 B.n414 VSUBS 0.010012f
C588 B.n415 VSUBS 0.010012f
C589 B.n416 VSUBS 0.010012f
C590 B.n417 VSUBS 0.010012f
C591 B.n418 VSUBS 0.010012f
C592 B.n419 VSUBS 0.010012f
C593 B.n420 VSUBS 0.010012f
C594 B.n421 VSUBS 0.010012f
C595 B.n422 VSUBS 0.010012f
C596 B.n423 VSUBS 0.010012f
C597 B.n424 VSUBS 0.010012f
C598 B.n425 VSUBS 0.010012f
C599 B.n426 VSUBS 0.010012f
C600 B.n427 VSUBS 0.010012f
C601 B.n428 VSUBS 0.010012f
C602 B.n429 VSUBS 0.010012f
C603 B.n430 VSUBS 0.010012f
C604 B.n431 VSUBS 0.010012f
C605 B.n432 VSUBS 0.010012f
C606 B.n433 VSUBS 0.010012f
C607 B.n434 VSUBS 0.023257f
C608 B.n435 VSUBS 0.023257f
C609 B.n436 VSUBS 0.022386f
C610 B.n437 VSUBS 0.010012f
C611 B.n438 VSUBS 0.010012f
C612 B.n439 VSUBS 0.010012f
C613 B.n440 VSUBS 0.010012f
C614 B.n441 VSUBS 0.010012f
C615 B.n442 VSUBS 0.010012f
C616 B.n443 VSUBS 0.010012f
C617 B.n444 VSUBS 0.010012f
C618 B.n445 VSUBS 0.010012f
C619 B.n446 VSUBS 0.010012f
C620 B.n447 VSUBS 0.010012f
C621 B.n448 VSUBS 0.010012f
C622 B.n449 VSUBS 0.010012f
C623 B.n450 VSUBS 0.010012f
C624 B.n451 VSUBS 0.010012f
C625 B.n452 VSUBS 0.010012f
C626 B.n453 VSUBS 0.010012f
C627 B.n454 VSUBS 0.010012f
C628 B.n455 VSUBS 0.010012f
C629 B.n456 VSUBS 0.010012f
C630 B.n457 VSUBS 0.010012f
C631 B.n458 VSUBS 0.010012f
C632 B.n459 VSUBS 0.010012f
C633 B.n460 VSUBS 0.010012f
C634 B.n461 VSUBS 0.010012f
C635 B.n462 VSUBS 0.010012f
C636 B.n463 VSUBS 0.010012f
C637 B.n464 VSUBS 0.010012f
C638 B.n465 VSUBS 0.010012f
C639 B.n466 VSUBS 0.010012f
C640 B.n467 VSUBS 0.010012f
C641 B.n468 VSUBS 0.010012f
C642 B.n469 VSUBS 0.010012f
C643 B.n470 VSUBS 0.010012f
C644 B.n471 VSUBS 0.010012f
C645 B.n472 VSUBS 0.010012f
C646 B.n473 VSUBS 0.010012f
C647 B.n474 VSUBS 0.010012f
C648 B.n475 VSUBS 0.010012f
C649 B.n476 VSUBS 0.010012f
C650 B.n477 VSUBS 0.010012f
C651 B.n478 VSUBS 0.010012f
C652 B.n479 VSUBS 0.010012f
C653 B.n480 VSUBS 0.010012f
C654 B.n481 VSUBS 0.010012f
C655 B.n482 VSUBS 0.010012f
C656 B.n483 VSUBS 0.010012f
C657 B.n484 VSUBS 0.010012f
C658 B.n485 VSUBS 0.010012f
C659 B.n486 VSUBS 0.010012f
C660 B.n487 VSUBS 0.010012f
C661 B.n488 VSUBS 0.010012f
C662 B.n489 VSUBS 0.010012f
C663 B.n490 VSUBS 0.010012f
C664 B.n491 VSUBS 0.010012f
C665 B.n492 VSUBS 0.010012f
C666 B.n493 VSUBS 0.010012f
C667 B.n494 VSUBS 0.010012f
C668 B.n495 VSUBS 0.010012f
C669 B.n496 VSUBS 0.010012f
C670 B.n497 VSUBS 0.010012f
C671 B.n498 VSUBS 0.010012f
C672 B.n499 VSUBS 0.010012f
C673 B.n500 VSUBS 0.010012f
C674 B.n501 VSUBS 0.010012f
C675 B.n502 VSUBS 0.010012f
C676 B.n503 VSUBS 0.010012f
C677 B.n504 VSUBS 0.010012f
C678 B.n505 VSUBS 0.010012f
C679 B.n506 VSUBS 0.010012f
C680 B.n507 VSUBS 0.010012f
C681 B.n508 VSUBS 0.010012f
C682 B.n509 VSUBS 0.010012f
C683 B.n510 VSUBS 0.010012f
C684 B.n511 VSUBS 0.010012f
C685 B.n512 VSUBS 0.010012f
C686 B.n513 VSUBS 0.010012f
C687 B.n514 VSUBS 0.010012f
C688 B.n515 VSUBS 0.010012f
C689 B.n516 VSUBS 0.010012f
C690 B.n517 VSUBS 0.010012f
C691 B.n518 VSUBS 0.010012f
C692 B.n519 VSUBS 0.010012f
C693 B.n520 VSUBS 0.010012f
C694 B.n521 VSUBS 0.010012f
C695 B.n522 VSUBS 0.010012f
C696 B.n523 VSUBS 0.010012f
C697 B.n524 VSUBS 0.010012f
C698 B.n525 VSUBS 0.010012f
C699 B.n526 VSUBS 0.010012f
C700 B.n527 VSUBS 0.010012f
C701 B.n528 VSUBS 0.010012f
C702 B.n529 VSUBS 0.010012f
C703 B.n530 VSUBS 0.010012f
C704 B.n531 VSUBS 0.010012f
C705 B.n532 VSUBS 0.010012f
C706 B.n533 VSUBS 0.010012f
C707 B.n534 VSUBS 0.010012f
C708 B.n535 VSUBS 0.010012f
C709 B.n536 VSUBS 0.010012f
C710 B.n537 VSUBS 0.010012f
C711 B.n538 VSUBS 0.010012f
C712 B.n539 VSUBS 0.010012f
C713 B.n540 VSUBS 0.010012f
C714 B.n541 VSUBS 0.010012f
C715 B.n542 VSUBS 0.010012f
C716 B.n543 VSUBS 0.010012f
C717 B.n544 VSUBS 0.010012f
C718 B.n545 VSUBS 0.010012f
C719 B.n546 VSUBS 0.010012f
C720 B.n547 VSUBS 0.010012f
C721 B.n548 VSUBS 0.010012f
C722 B.n549 VSUBS 0.010012f
C723 B.n550 VSUBS 0.010012f
C724 B.n551 VSUBS 0.010012f
C725 B.n552 VSUBS 0.010012f
C726 B.n553 VSUBS 0.010012f
C727 B.n554 VSUBS 0.010012f
C728 B.n555 VSUBS 0.010012f
C729 B.n556 VSUBS 0.010012f
C730 B.n557 VSUBS 0.010012f
C731 B.n558 VSUBS 0.010012f
C732 B.n559 VSUBS 0.010012f
C733 B.n560 VSUBS 0.010012f
C734 B.n561 VSUBS 0.010012f
C735 B.n562 VSUBS 0.010012f
C736 B.n563 VSUBS 0.010012f
C737 B.n564 VSUBS 0.010012f
C738 B.n565 VSUBS 0.010012f
C739 B.n566 VSUBS 0.010012f
C740 B.n567 VSUBS 0.010012f
C741 B.n568 VSUBS 0.010012f
C742 B.n569 VSUBS 0.010012f
C743 B.n570 VSUBS 0.010012f
C744 B.n571 VSUBS 0.010012f
C745 B.n572 VSUBS 0.010012f
C746 B.n573 VSUBS 0.010012f
C747 B.n574 VSUBS 0.010012f
C748 B.n575 VSUBS 0.010012f
C749 B.n576 VSUBS 0.010012f
C750 B.n577 VSUBS 0.010012f
C751 B.n578 VSUBS 0.010012f
C752 B.n579 VSUBS 0.010012f
C753 B.n580 VSUBS 0.010012f
C754 B.n581 VSUBS 0.010012f
C755 B.n582 VSUBS 0.010012f
C756 B.n583 VSUBS 0.010012f
C757 B.n584 VSUBS 0.010012f
C758 B.n585 VSUBS 0.010012f
C759 B.n586 VSUBS 0.010012f
C760 B.n587 VSUBS 0.010012f
C761 B.n588 VSUBS 0.010012f
C762 B.n589 VSUBS 0.010012f
C763 B.n590 VSUBS 0.010012f
C764 B.n591 VSUBS 0.010012f
C765 B.n592 VSUBS 0.010012f
C766 B.n593 VSUBS 0.010012f
C767 B.n594 VSUBS 0.010012f
C768 B.n595 VSUBS 0.010012f
C769 B.n596 VSUBS 0.010012f
C770 B.n597 VSUBS 0.010012f
C771 B.n598 VSUBS 0.010012f
C772 B.n599 VSUBS 0.010012f
C773 B.n600 VSUBS 0.010012f
C774 B.n601 VSUBS 0.010012f
C775 B.n602 VSUBS 0.010012f
C776 B.n603 VSUBS 0.010012f
C777 B.n604 VSUBS 0.010012f
C778 B.n605 VSUBS 0.010012f
C779 B.n606 VSUBS 0.010012f
C780 B.n607 VSUBS 0.010012f
C781 B.n608 VSUBS 0.010012f
C782 B.n609 VSUBS 0.010012f
C783 B.n610 VSUBS 0.010012f
C784 B.n611 VSUBS 0.010012f
C785 B.n612 VSUBS 0.010012f
C786 B.n613 VSUBS 0.010012f
C787 B.n614 VSUBS 0.010012f
C788 B.n615 VSUBS 0.010012f
C789 B.n616 VSUBS 0.010012f
C790 B.n617 VSUBS 0.010012f
C791 B.n618 VSUBS 0.010012f
C792 B.n619 VSUBS 0.010012f
C793 B.n620 VSUBS 0.010012f
C794 B.n621 VSUBS 0.010012f
C795 B.n622 VSUBS 0.010012f
C796 B.n623 VSUBS 0.010012f
C797 B.n624 VSUBS 0.010012f
C798 B.n625 VSUBS 0.010012f
C799 B.n626 VSUBS 0.010012f
C800 B.n627 VSUBS 0.010012f
C801 B.n628 VSUBS 0.010012f
C802 B.n629 VSUBS 0.010012f
C803 B.n630 VSUBS 0.010012f
C804 B.n631 VSUBS 0.010012f
C805 B.n632 VSUBS 0.010012f
C806 B.n633 VSUBS 0.010012f
C807 B.n634 VSUBS 0.010012f
C808 B.n635 VSUBS 0.010012f
C809 B.n636 VSUBS 0.010012f
C810 B.n637 VSUBS 0.022386f
C811 B.n638 VSUBS 0.023257f
C812 B.n639 VSUBS 0.022026f
C813 B.n640 VSUBS 0.010012f
C814 B.n641 VSUBS 0.010012f
C815 B.n642 VSUBS 0.010012f
C816 B.n643 VSUBS 0.010012f
C817 B.n644 VSUBS 0.010012f
C818 B.n645 VSUBS 0.010012f
C819 B.n646 VSUBS 0.010012f
C820 B.n647 VSUBS 0.010012f
C821 B.n648 VSUBS 0.010012f
C822 B.n649 VSUBS 0.010012f
C823 B.n650 VSUBS 0.010012f
C824 B.n651 VSUBS 0.010012f
C825 B.n652 VSUBS 0.010012f
C826 B.n653 VSUBS 0.010012f
C827 B.n654 VSUBS 0.010012f
C828 B.n655 VSUBS 0.010012f
C829 B.n656 VSUBS 0.010012f
C830 B.n657 VSUBS 0.010012f
C831 B.n658 VSUBS 0.010012f
C832 B.n659 VSUBS 0.010012f
C833 B.n660 VSUBS 0.010012f
C834 B.n661 VSUBS 0.010012f
C835 B.n662 VSUBS 0.010012f
C836 B.n663 VSUBS 0.010012f
C837 B.n664 VSUBS 0.010012f
C838 B.n665 VSUBS 0.010012f
C839 B.n666 VSUBS 0.010012f
C840 B.n667 VSUBS 0.010012f
C841 B.n668 VSUBS 0.010012f
C842 B.n669 VSUBS 0.010012f
C843 B.n670 VSUBS 0.010012f
C844 B.n671 VSUBS 0.010012f
C845 B.n672 VSUBS 0.010012f
C846 B.n673 VSUBS 0.010012f
C847 B.n674 VSUBS 0.010012f
C848 B.n675 VSUBS 0.010012f
C849 B.n676 VSUBS 0.010012f
C850 B.n677 VSUBS 0.010012f
C851 B.n678 VSUBS 0.010012f
C852 B.n679 VSUBS 0.010012f
C853 B.n680 VSUBS 0.010012f
C854 B.n681 VSUBS 0.010012f
C855 B.n682 VSUBS 0.010012f
C856 B.n683 VSUBS 0.010012f
C857 B.n684 VSUBS 0.010012f
C858 B.n685 VSUBS 0.010012f
C859 B.n686 VSUBS 0.010012f
C860 B.n687 VSUBS 0.009423f
C861 B.n688 VSUBS 0.023197f
C862 B.n689 VSUBS 0.005595f
C863 B.n690 VSUBS 0.010012f
C864 B.n691 VSUBS 0.010012f
C865 B.n692 VSUBS 0.010012f
C866 B.n693 VSUBS 0.010012f
C867 B.n694 VSUBS 0.010012f
C868 B.n695 VSUBS 0.010012f
C869 B.n696 VSUBS 0.010012f
C870 B.n697 VSUBS 0.010012f
C871 B.n698 VSUBS 0.010012f
C872 B.n699 VSUBS 0.010012f
C873 B.n700 VSUBS 0.010012f
C874 B.n701 VSUBS 0.010012f
C875 B.n702 VSUBS 0.005595f
C876 B.n703 VSUBS 0.010012f
C877 B.n704 VSUBS 0.010012f
C878 B.n705 VSUBS 0.009423f
C879 B.n706 VSUBS 0.010012f
C880 B.n707 VSUBS 0.010012f
C881 B.n708 VSUBS 0.010012f
C882 B.n709 VSUBS 0.010012f
C883 B.n710 VSUBS 0.010012f
C884 B.n711 VSUBS 0.010012f
C885 B.n712 VSUBS 0.010012f
C886 B.n713 VSUBS 0.010012f
C887 B.n714 VSUBS 0.010012f
C888 B.n715 VSUBS 0.010012f
C889 B.n716 VSUBS 0.010012f
C890 B.n717 VSUBS 0.010012f
C891 B.n718 VSUBS 0.010012f
C892 B.n719 VSUBS 0.010012f
C893 B.n720 VSUBS 0.010012f
C894 B.n721 VSUBS 0.010012f
C895 B.n722 VSUBS 0.010012f
C896 B.n723 VSUBS 0.010012f
C897 B.n724 VSUBS 0.010012f
C898 B.n725 VSUBS 0.010012f
C899 B.n726 VSUBS 0.010012f
C900 B.n727 VSUBS 0.010012f
C901 B.n728 VSUBS 0.010012f
C902 B.n729 VSUBS 0.010012f
C903 B.n730 VSUBS 0.010012f
C904 B.n731 VSUBS 0.010012f
C905 B.n732 VSUBS 0.010012f
C906 B.n733 VSUBS 0.010012f
C907 B.n734 VSUBS 0.010012f
C908 B.n735 VSUBS 0.010012f
C909 B.n736 VSUBS 0.010012f
C910 B.n737 VSUBS 0.010012f
C911 B.n738 VSUBS 0.010012f
C912 B.n739 VSUBS 0.010012f
C913 B.n740 VSUBS 0.010012f
C914 B.n741 VSUBS 0.010012f
C915 B.n742 VSUBS 0.010012f
C916 B.n743 VSUBS 0.010012f
C917 B.n744 VSUBS 0.010012f
C918 B.n745 VSUBS 0.010012f
C919 B.n746 VSUBS 0.010012f
C920 B.n747 VSUBS 0.010012f
C921 B.n748 VSUBS 0.010012f
C922 B.n749 VSUBS 0.010012f
C923 B.n750 VSUBS 0.010012f
C924 B.n751 VSUBS 0.010012f
C925 B.n752 VSUBS 0.023257f
C926 B.n753 VSUBS 0.023257f
C927 B.n754 VSUBS 0.022386f
C928 B.n755 VSUBS 0.010012f
C929 B.n756 VSUBS 0.010012f
C930 B.n757 VSUBS 0.010012f
C931 B.n758 VSUBS 0.010012f
C932 B.n759 VSUBS 0.010012f
C933 B.n760 VSUBS 0.010012f
C934 B.n761 VSUBS 0.010012f
C935 B.n762 VSUBS 0.010012f
C936 B.n763 VSUBS 0.010012f
C937 B.n764 VSUBS 0.010012f
C938 B.n765 VSUBS 0.010012f
C939 B.n766 VSUBS 0.010012f
C940 B.n767 VSUBS 0.010012f
C941 B.n768 VSUBS 0.010012f
C942 B.n769 VSUBS 0.010012f
C943 B.n770 VSUBS 0.010012f
C944 B.n771 VSUBS 0.010012f
C945 B.n772 VSUBS 0.010012f
C946 B.n773 VSUBS 0.010012f
C947 B.n774 VSUBS 0.010012f
C948 B.n775 VSUBS 0.010012f
C949 B.n776 VSUBS 0.010012f
C950 B.n777 VSUBS 0.010012f
C951 B.n778 VSUBS 0.010012f
C952 B.n779 VSUBS 0.010012f
C953 B.n780 VSUBS 0.010012f
C954 B.n781 VSUBS 0.010012f
C955 B.n782 VSUBS 0.010012f
C956 B.n783 VSUBS 0.010012f
C957 B.n784 VSUBS 0.010012f
C958 B.n785 VSUBS 0.010012f
C959 B.n786 VSUBS 0.010012f
C960 B.n787 VSUBS 0.010012f
C961 B.n788 VSUBS 0.010012f
C962 B.n789 VSUBS 0.010012f
C963 B.n790 VSUBS 0.010012f
C964 B.n791 VSUBS 0.010012f
C965 B.n792 VSUBS 0.010012f
C966 B.n793 VSUBS 0.010012f
C967 B.n794 VSUBS 0.010012f
C968 B.n795 VSUBS 0.010012f
C969 B.n796 VSUBS 0.010012f
C970 B.n797 VSUBS 0.010012f
C971 B.n798 VSUBS 0.010012f
C972 B.n799 VSUBS 0.010012f
C973 B.n800 VSUBS 0.010012f
C974 B.n801 VSUBS 0.010012f
C975 B.n802 VSUBS 0.010012f
C976 B.n803 VSUBS 0.010012f
C977 B.n804 VSUBS 0.010012f
C978 B.n805 VSUBS 0.010012f
C979 B.n806 VSUBS 0.010012f
C980 B.n807 VSUBS 0.010012f
C981 B.n808 VSUBS 0.010012f
C982 B.n809 VSUBS 0.010012f
C983 B.n810 VSUBS 0.010012f
C984 B.n811 VSUBS 0.010012f
C985 B.n812 VSUBS 0.010012f
C986 B.n813 VSUBS 0.010012f
C987 B.n814 VSUBS 0.010012f
C988 B.n815 VSUBS 0.010012f
C989 B.n816 VSUBS 0.010012f
C990 B.n817 VSUBS 0.010012f
C991 B.n818 VSUBS 0.010012f
C992 B.n819 VSUBS 0.010012f
C993 B.n820 VSUBS 0.010012f
C994 B.n821 VSUBS 0.010012f
C995 B.n822 VSUBS 0.010012f
C996 B.n823 VSUBS 0.010012f
C997 B.n824 VSUBS 0.010012f
C998 B.n825 VSUBS 0.010012f
C999 B.n826 VSUBS 0.010012f
C1000 B.n827 VSUBS 0.010012f
C1001 B.n828 VSUBS 0.010012f
C1002 B.n829 VSUBS 0.010012f
C1003 B.n830 VSUBS 0.010012f
C1004 B.n831 VSUBS 0.010012f
C1005 B.n832 VSUBS 0.010012f
C1006 B.n833 VSUBS 0.010012f
C1007 B.n834 VSUBS 0.010012f
C1008 B.n835 VSUBS 0.010012f
C1009 B.n836 VSUBS 0.010012f
C1010 B.n837 VSUBS 0.010012f
C1011 B.n838 VSUBS 0.010012f
C1012 B.n839 VSUBS 0.010012f
C1013 B.n840 VSUBS 0.010012f
C1014 B.n841 VSUBS 0.010012f
C1015 B.n842 VSUBS 0.010012f
C1016 B.n843 VSUBS 0.010012f
C1017 B.n844 VSUBS 0.010012f
C1018 B.n845 VSUBS 0.010012f
C1019 B.n846 VSUBS 0.010012f
C1020 B.n847 VSUBS 0.010012f
C1021 B.n848 VSUBS 0.010012f
C1022 B.n849 VSUBS 0.010012f
C1023 B.n850 VSUBS 0.010012f
C1024 B.n851 VSUBS 0.010012f
C1025 B.n852 VSUBS 0.010012f
C1026 B.n853 VSUBS 0.010012f
C1027 B.n854 VSUBS 0.010012f
C1028 B.n855 VSUBS 0.022671f
C1029 VTAIL.t18 VSUBS 0.222252f
C1030 VTAIL.t12 VSUBS 0.222252f
C1031 VTAIL.n0 VSUBS 1.47567f
C1032 VTAIL.n1 VSUBS 1.08323f
C1033 VTAIL.t9 VSUBS 1.98006f
C1034 VTAIL.n2 VSUBS 1.2503f
C1035 VTAIL.t3 VSUBS 0.222252f
C1036 VTAIL.t1 VSUBS 0.222252f
C1037 VTAIL.n3 VSUBS 1.47567f
C1038 VTAIL.n4 VSUBS 1.24417f
C1039 VTAIL.t7 VSUBS 0.222252f
C1040 VTAIL.t5 VSUBS 0.222252f
C1041 VTAIL.n5 VSUBS 1.47567f
C1042 VTAIL.n6 VSUBS 2.72728f
C1043 VTAIL.t10 VSUBS 0.222252f
C1044 VTAIL.t11 VSUBS 0.222252f
C1045 VTAIL.n7 VSUBS 1.47568f
C1046 VTAIL.n8 VSUBS 2.72727f
C1047 VTAIL.t16 VSUBS 0.222252f
C1048 VTAIL.t14 VSUBS 0.222252f
C1049 VTAIL.n9 VSUBS 1.47568f
C1050 VTAIL.n10 VSUBS 1.24416f
C1051 VTAIL.t15 VSUBS 1.98007f
C1052 VTAIL.n11 VSUBS 1.25028f
C1053 VTAIL.t6 VSUBS 0.222252f
C1054 VTAIL.t8 VSUBS 0.222252f
C1055 VTAIL.n12 VSUBS 1.47568f
C1056 VTAIL.n13 VSUBS 1.14854f
C1057 VTAIL.t4 VSUBS 0.222252f
C1058 VTAIL.t2 VSUBS 0.222252f
C1059 VTAIL.n14 VSUBS 1.47568f
C1060 VTAIL.n15 VSUBS 1.24416f
C1061 VTAIL.t0 VSUBS 1.98007f
C1062 VTAIL.n16 VSUBS 2.5447f
C1063 VTAIL.t17 VSUBS 1.98006f
C1064 VTAIL.n17 VSUBS 2.54471f
C1065 VTAIL.t13 VSUBS 0.222252f
C1066 VTAIL.t19 VSUBS 0.222252f
C1067 VTAIL.n18 VSUBS 1.47567f
C1068 VTAIL.n19 VSUBS 1.02517f
C1069 VDD2.t3 VSUBS 2.26148f
C1070 VDD2.t9 VSUBS 0.230714f
C1071 VDD2.t7 VSUBS 0.230714f
C1072 VDD2.n0 VSUBS 1.68967f
C1073 VDD2.n1 VSUBS 1.90336f
C1074 VDD2.t1 VSUBS 0.230714f
C1075 VDD2.t6 VSUBS 0.230714f
C1076 VDD2.n2 VSUBS 1.71875f
C1077 VDD2.n3 VSUBS 4.07074f
C1078 VDD2.t0 VSUBS 2.228f
C1079 VDD2.n4 VSUBS 4.2359f
C1080 VDD2.t4 VSUBS 0.230714f
C1081 VDD2.t8 VSUBS 0.230714f
C1082 VDD2.n5 VSUBS 1.68968f
C1083 VDD2.n6 VSUBS 0.961708f
C1084 VDD2.t5 VSUBS 0.230714f
C1085 VDD2.t2 VSUBS 0.230714f
C1086 VDD2.n7 VSUBS 1.7187f
C1087 VN.t2 VSUBS 2.12311f
C1088 VN.n0 VSUBS 0.874091f
C1089 VN.n1 VSUBS 0.028642f
C1090 VN.n2 VSUBS 0.041416f
C1091 VN.n3 VSUBS 0.028642f
C1092 VN.t0 VSUBS 2.12311f
C1093 VN.n4 VSUBS 0.053382f
C1094 VN.n5 VSUBS 0.028642f
C1095 VN.n6 VSUBS 0.053382f
C1096 VN.n7 VSUBS 0.028642f
C1097 VN.t6 VSUBS 2.12311f
C1098 VN.n8 VSUBS 0.053382f
C1099 VN.n9 VSUBS 0.028642f
C1100 VN.n10 VSUBS 0.031244f
C1101 VN.t7 VSUBS 2.12311f
C1102 VN.n11 VSUBS 0.843419f
C1103 VN.t1 VSUBS 2.41009f
C1104 VN.n12 VSUBS 0.817138f
C1105 VN.n13 VSUBS 0.309758f
C1106 VN.n14 VSUBS 0.028642f
C1107 VN.n15 VSUBS 0.053382f
C1108 VN.n16 VSUBS 0.057701f
C1109 VN.n17 VSUBS 0.025929f
C1110 VN.n18 VSUBS 0.028642f
C1111 VN.n19 VSUBS 0.028642f
C1112 VN.n20 VSUBS 0.028642f
C1113 VN.n21 VSUBS 0.053382f
C1114 VN.n22 VSUBS 0.040204f
C1115 VN.n23 VSUBS 0.760814f
C1116 VN.n24 VSUBS 0.040204f
C1117 VN.n25 VSUBS 0.028642f
C1118 VN.n26 VSUBS 0.028642f
C1119 VN.n27 VSUBS 0.028642f
C1120 VN.n28 VSUBS 0.053382f
C1121 VN.n29 VSUBS 0.025929f
C1122 VN.n30 VSUBS 0.057701f
C1123 VN.n31 VSUBS 0.028642f
C1124 VN.n32 VSUBS 0.028642f
C1125 VN.n33 VSUBS 0.028642f
C1126 VN.n34 VSUBS 0.031244f
C1127 VN.n35 VSUBS 0.760814f
C1128 VN.n36 VSUBS 0.049165f
C1129 VN.n37 VSUBS 0.053382f
C1130 VN.n38 VSUBS 0.028642f
C1131 VN.n39 VSUBS 0.028642f
C1132 VN.n40 VSUBS 0.028642f
C1133 VN.n41 VSUBS 0.042214f
C1134 VN.n42 VSUBS 0.053382f
C1135 VN.n43 VSUBS 0.048638f
C1136 VN.n44 VSUBS 0.046228f
C1137 VN.n45 VSUBS 0.059527f
C1138 VN.t9 VSUBS 2.12311f
C1139 VN.n46 VSUBS 0.874091f
C1140 VN.n47 VSUBS 0.028642f
C1141 VN.n48 VSUBS 0.041416f
C1142 VN.n49 VSUBS 0.028642f
C1143 VN.t8 VSUBS 2.12311f
C1144 VN.n50 VSUBS 0.053382f
C1145 VN.n51 VSUBS 0.028642f
C1146 VN.n52 VSUBS 0.053382f
C1147 VN.n53 VSUBS 0.028642f
C1148 VN.t3 VSUBS 2.12311f
C1149 VN.n54 VSUBS 0.053382f
C1150 VN.n55 VSUBS 0.028642f
C1151 VN.n56 VSUBS 0.031244f
C1152 VN.t4 VSUBS 2.41009f
C1153 VN.t5 VSUBS 2.12311f
C1154 VN.n57 VSUBS 0.843419f
C1155 VN.n58 VSUBS 0.817138f
C1156 VN.n59 VSUBS 0.309758f
C1157 VN.n60 VSUBS 0.028642f
C1158 VN.n61 VSUBS 0.053382f
C1159 VN.n62 VSUBS 0.057701f
C1160 VN.n63 VSUBS 0.025929f
C1161 VN.n64 VSUBS 0.028642f
C1162 VN.n65 VSUBS 0.028642f
C1163 VN.n66 VSUBS 0.028642f
C1164 VN.n67 VSUBS 0.053382f
C1165 VN.n68 VSUBS 0.040204f
C1166 VN.n69 VSUBS 0.760814f
C1167 VN.n70 VSUBS 0.040204f
C1168 VN.n71 VSUBS 0.028642f
C1169 VN.n72 VSUBS 0.028642f
C1170 VN.n73 VSUBS 0.028642f
C1171 VN.n74 VSUBS 0.053382f
C1172 VN.n75 VSUBS 0.025929f
C1173 VN.n76 VSUBS 0.057701f
C1174 VN.n77 VSUBS 0.028642f
C1175 VN.n78 VSUBS 0.028642f
C1176 VN.n79 VSUBS 0.028642f
C1177 VN.n80 VSUBS 0.031244f
C1178 VN.n81 VSUBS 0.760814f
C1179 VN.n82 VSUBS 0.049165f
C1180 VN.n83 VSUBS 0.053382f
C1181 VN.n84 VSUBS 0.028642f
C1182 VN.n85 VSUBS 0.028642f
C1183 VN.n86 VSUBS 0.028642f
C1184 VN.n87 VSUBS 0.042214f
C1185 VN.n88 VSUBS 0.053382f
C1186 VN.n89 VSUBS 0.048638f
C1187 VN.n90 VSUBS 0.046228f
C1188 VN.n91 VSUBS 1.78269f
.ends

