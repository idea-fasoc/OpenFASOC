* NGSPICE file created from diff_pair_sample_1375.ext - technology: sky130A

.subckt diff_pair_sample_1375 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=0 ps=0 w=6.39 l=0.68
X1 VDD2.t9 VN.t0 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X2 VTAIL.t5 VN.t1 VDD2.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X3 VDD2.t7 VN.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X4 VDD1.t9 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=2.4921 ps=13.56 w=6.39 l=0.68
X5 VTAIL.t4 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X6 VTAIL.t15 VP.t1 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X7 VTAIL.t1 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X8 VTAIL.t6 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X9 VDD2.t4 VN.t5 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=2.4921 ps=13.56 w=6.39 l=0.68
X10 VDD1.t6 VP.t3 VTAIL.t19 B.t5 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=2.4921 ps=13.56 w=6.39 l=0.68
X11 VDD1.t5 VP.t4 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=1.05435 ps=6.72 w=6.39 l=0.68
X12 VDD1.t4 VP.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X13 VDD2.t3 VN.t6 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=1.05435 ps=6.72 w=6.39 l=0.68
X14 VDD2.t2 VN.t7 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=2.4921 ps=13.56 w=6.39 l=0.68
X15 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=0 ps=0 w=6.39 l=0.68
X16 VTAIL.t16 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X17 VDD1.t2 VP.t7 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=1.05435 ps=6.72 w=6.39 l=0.68
X18 VTAIL.t17 VP.t8 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X19 VDD2.t1 VN.t8 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=1.05435 ps=6.72 w=6.39 l=0.68
X20 VTAIL.t8 VN.t9 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
X21 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=0 ps=0 w=6.39 l=0.68
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4921 pd=13.56 as=0 ps=0 w=6.39 l=0.68
X23 VDD1.t0 VP.t9 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.05435 pd=6.72 as=1.05435 ps=6.72 w=6.39 l=0.68
R0 B.n402 B.n401 585
R1 B.n404 B.n85 585
R2 B.n407 B.n406 585
R3 B.n408 B.n84 585
R4 B.n410 B.n409 585
R5 B.n412 B.n83 585
R6 B.n415 B.n414 585
R7 B.n416 B.n82 585
R8 B.n418 B.n417 585
R9 B.n420 B.n81 585
R10 B.n423 B.n422 585
R11 B.n424 B.n80 585
R12 B.n426 B.n425 585
R13 B.n428 B.n79 585
R14 B.n431 B.n430 585
R15 B.n432 B.n78 585
R16 B.n434 B.n433 585
R17 B.n436 B.n77 585
R18 B.n439 B.n438 585
R19 B.n440 B.n76 585
R20 B.n442 B.n441 585
R21 B.n444 B.n75 585
R22 B.n447 B.n446 585
R23 B.n448 B.n71 585
R24 B.n450 B.n449 585
R25 B.n452 B.n70 585
R26 B.n455 B.n454 585
R27 B.n456 B.n69 585
R28 B.n458 B.n457 585
R29 B.n460 B.n68 585
R30 B.n463 B.n462 585
R31 B.n464 B.n67 585
R32 B.n466 B.n465 585
R33 B.n468 B.n66 585
R34 B.n471 B.n470 585
R35 B.n473 B.n63 585
R36 B.n475 B.n474 585
R37 B.n477 B.n62 585
R38 B.n480 B.n479 585
R39 B.n481 B.n61 585
R40 B.n483 B.n482 585
R41 B.n485 B.n60 585
R42 B.n488 B.n487 585
R43 B.n489 B.n59 585
R44 B.n491 B.n490 585
R45 B.n493 B.n58 585
R46 B.n496 B.n495 585
R47 B.n497 B.n57 585
R48 B.n499 B.n498 585
R49 B.n501 B.n56 585
R50 B.n504 B.n503 585
R51 B.n505 B.n55 585
R52 B.n507 B.n506 585
R53 B.n509 B.n54 585
R54 B.n512 B.n511 585
R55 B.n513 B.n53 585
R56 B.n515 B.n514 585
R57 B.n517 B.n52 585
R58 B.n520 B.n519 585
R59 B.n521 B.n51 585
R60 B.n400 B.n49 585
R61 B.n524 B.n49 585
R62 B.n399 B.n48 585
R63 B.n525 B.n48 585
R64 B.n398 B.n47 585
R65 B.n526 B.n47 585
R66 B.n397 B.n396 585
R67 B.n396 B.n43 585
R68 B.n395 B.n42 585
R69 B.n532 B.n42 585
R70 B.n394 B.n41 585
R71 B.n533 B.n41 585
R72 B.n393 B.n40 585
R73 B.n534 B.n40 585
R74 B.n392 B.n391 585
R75 B.n391 B.n36 585
R76 B.n390 B.n35 585
R77 B.n540 B.n35 585
R78 B.n389 B.n34 585
R79 B.n541 B.n34 585
R80 B.n388 B.n33 585
R81 B.n542 B.n33 585
R82 B.n387 B.n386 585
R83 B.n386 B.n32 585
R84 B.n385 B.n28 585
R85 B.n548 B.n28 585
R86 B.n384 B.n27 585
R87 B.n549 B.n27 585
R88 B.n383 B.n26 585
R89 B.t0 B.n26 585
R90 B.n382 B.n381 585
R91 B.n381 B.n22 585
R92 B.n380 B.n21 585
R93 B.n555 B.n21 585
R94 B.n379 B.n20 585
R95 B.n556 B.n20 585
R96 B.n378 B.n19 585
R97 B.n557 B.n19 585
R98 B.n377 B.n376 585
R99 B.n376 B.n18 585
R100 B.n375 B.n14 585
R101 B.n563 B.n14 585
R102 B.n374 B.n13 585
R103 B.n564 B.n13 585
R104 B.n373 B.n12 585
R105 B.n565 B.n12 585
R106 B.n372 B.n371 585
R107 B.n371 B.n8 585
R108 B.n370 B.n7 585
R109 B.n571 B.n7 585
R110 B.n369 B.n6 585
R111 B.n572 B.n6 585
R112 B.n368 B.n5 585
R113 B.n573 B.n5 585
R114 B.n367 B.n366 585
R115 B.n366 B.n4 585
R116 B.n365 B.n86 585
R117 B.n365 B.n364 585
R118 B.n355 B.n87 585
R119 B.n88 B.n87 585
R120 B.n357 B.n356 585
R121 B.n358 B.n357 585
R122 B.n354 B.n93 585
R123 B.n93 B.n92 585
R124 B.n353 B.n352 585
R125 B.n352 B.n351 585
R126 B.n95 B.n94 585
R127 B.n344 B.n95 585
R128 B.n343 B.n342 585
R129 B.n345 B.n343 585
R130 B.n341 B.n100 585
R131 B.n100 B.n99 585
R132 B.n340 B.n339 585
R133 B.n339 B.n338 585
R134 B.n102 B.n101 585
R135 B.n103 B.n102 585
R136 B.n332 B.n331 585
R137 B.t4 B.n332 585
R138 B.n330 B.n108 585
R139 B.n108 B.n107 585
R140 B.n329 B.n328 585
R141 B.n328 B.n327 585
R142 B.n110 B.n109 585
R143 B.n320 B.n110 585
R144 B.n319 B.n318 585
R145 B.n321 B.n319 585
R146 B.n317 B.n115 585
R147 B.n115 B.n114 585
R148 B.n316 B.n315 585
R149 B.n315 B.n314 585
R150 B.n117 B.n116 585
R151 B.n118 B.n117 585
R152 B.n307 B.n306 585
R153 B.n308 B.n307 585
R154 B.n305 B.n123 585
R155 B.n123 B.n122 585
R156 B.n304 B.n303 585
R157 B.n303 B.n302 585
R158 B.n125 B.n124 585
R159 B.n126 B.n125 585
R160 B.n295 B.n294 585
R161 B.n296 B.n295 585
R162 B.n293 B.n131 585
R163 B.n131 B.n130 585
R164 B.n292 B.n291 585
R165 B.n291 B.n290 585
R166 B.n287 B.n135 585
R167 B.n286 B.n285 585
R168 B.n283 B.n136 585
R169 B.n283 B.n134 585
R170 B.n282 B.n281 585
R171 B.n280 B.n279 585
R172 B.n278 B.n138 585
R173 B.n276 B.n275 585
R174 B.n274 B.n139 585
R175 B.n273 B.n272 585
R176 B.n270 B.n140 585
R177 B.n268 B.n267 585
R178 B.n266 B.n141 585
R179 B.n265 B.n264 585
R180 B.n262 B.n142 585
R181 B.n260 B.n259 585
R182 B.n258 B.n143 585
R183 B.n257 B.n256 585
R184 B.n254 B.n144 585
R185 B.n252 B.n251 585
R186 B.n250 B.n145 585
R187 B.n249 B.n248 585
R188 B.n246 B.n146 585
R189 B.n244 B.n243 585
R190 B.n242 B.n147 585
R191 B.n241 B.n240 585
R192 B.n238 B.n237 585
R193 B.n236 B.n235 585
R194 B.n234 B.n152 585
R195 B.n232 B.n231 585
R196 B.n230 B.n153 585
R197 B.n229 B.n228 585
R198 B.n226 B.n154 585
R199 B.n224 B.n223 585
R200 B.n222 B.n155 585
R201 B.n221 B.n220 585
R202 B.n218 B.n217 585
R203 B.n216 B.n215 585
R204 B.n214 B.n160 585
R205 B.n212 B.n211 585
R206 B.n210 B.n161 585
R207 B.n209 B.n208 585
R208 B.n206 B.n162 585
R209 B.n204 B.n203 585
R210 B.n202 B.n163 585
R211 B.n201 B.n200 585
R212 B.n198 B.n164 585
R213 B.n196 B.n195 585
R214 B.n194 B.n165 585
R215 B.n193 B.n192 585
R216 B.n190 B.n166 585
R217 B.n188 B.n187 585
R218 B.n186 B.n167 585
R219 B.n185 B.n184 585
R220 B.n182 B.n168 585
R221 B.n180 B.n179 585
R222 B.n178 B.n169 585
R223 B.n177 B.n176 585
R224 B.n174 B.n170 585
R225 B.n172 B.n171 585
R226 B.n133 B.n132 585
R227 B.n134 B.n133 585
R228 B.n289 B.n288 585
R229 B.n290 B.n289 585
R230 B.n129 B.n128 585
R231 B.n130 B.n129 585
R232 B.n298 B.n297 585
R233 B.n297 B.n296 585
R234 B.n299 B.n127 585
R235 B.n127 B.n126 585
R236 B.n301 B.n300 585
R237 B.n302 B.n301 585
R238 B.n121 B.n120 585
R239 B.n122 B.n121 585
R240 B.n310 B.n309 585
R241 B.n309 B.n308 585
R242 B.n311 B.n119 585
R243 B.n119 B.n118 585
R244 B.n313 B.n312 585
R245 B.n314 B.n313 585
R246 B.n113 B.n112 585
R247 B.n114 B.n113 585
R248 B.n323 B.n322 585
R249 B.n322 B.n321 585
R250 B.n324 B.n111 585
R251 B.n320 B.n111 585
R252 B.n326 B.n325 585
R253 B.n327 B.n326 585
R254 B.n106 B.n105 585
R255 B.n107 B.n106 585
R256 B.n334 B.n333 585
R257 B.n333 B.t4 585
R258 B.n335 B.n104 585
R259 B.n104 B.n103 585
R260 B.n337 B.n336 585
R261 B.n338 B.n337 585
R262 B.n98 B.n97 585
R263 B.n99 B.n98 585
R264 B.n347 B.n346 585
R265 B.n346 B.n345 585
R266 B.n348 B.n96 585
R267 B.n344 B.n96 585
R268 B.n350 B.n349 585
R269 B.n351 B.n350 585
R270 B.n91 B.n90 585
R271 B.n92 B.n91 585
R272 B.n360 B.n359 585
R273 B.n359 B.n358 585
R274 B.n361 B.n89 585
R275 B.n89 B.n88 585
R276 B.n363 B.n362 585
R277 B.n364 B.n363 585
R278 B.n2 B.n0 585
R279 B.n4 B.n2 585
R280 B.n3 B.n1 585
R281 B.n572 B.n3 585
R282 B.n570 B.n569 585
R283 B.n571 B.n570 585
R284 B.n568 B.n9 585
R285 B.n9 B.n8 585
R286 B.n567 B.n566 585
R287 B.n566 B.n565 585
R288 B.n11 B.n10 585
R289 B.n564 B.n11 585
R290 B.n562 B.n561 585
R291 B.n563 B.n562 585
R292 B.n560 B.n15 585
R293 B.n18 B.n15 585
R294 B.n559 B.n558 585
R295 B.n558 B.n557 585
R296 B.n17 B.n16 585
R297 B.n556 B.n17 585
R298 B.n554 B.n553 585
R299 B.n555 B.n554 585
R300 B.n552 B.n23 585
R301 B.n23 B.n22 585
R302 B.n551 B.n550 585
R303 B.n550 B.t0 585
R304 B.n25 B.n24 585
R305 B.n549 B.n25 585
R306 B.n547 B.n546 585
R307 B.n548 B.n547 585
R308 B.n545 B.n29 585
R309 B.n32 B.n29 585
R310 B.n544 B.n543 585
R311 B.n543 B.n542 585
R312 B.n31 B.n30 585
R313 B.n541 B.n31 585
R314 B.n539 B.n538 585
R315 B.n540 B.n539 585
R316 B.n537 B.n37 585
R317 B.n37 B.n36 585
R318 B.n536 B.n535 585
R319 B.n535 B.n534 585
R320 B.n39 B.n38 585
R321 B.n533 B.n39 585
R322 B.n531 B.n530 585
R323 B.n532 B.n531 585
R324 B.n529 B.n44 585
R325 B.n44 B.n43 585
R326 B.n528 B.n527 585
R327 B.n527 B.n526 585
R328 B.n46 B.n45 585
R329 B.n525 B.n46 585
R330 B.n523 B.n522 585
R331 B.n524 B.n523 585
R332 B.n575 B.n574 585
R333 B.n574 B.n573 585
R334 B.n289 B.n135 473.281
R335 B.n523 B.n51 473.281
R336 B.n291 B.n133 473.281
R337 B.n402 B.n49 473.281
R338 B.n156 B.t17 429.688
R339 B.n148 B.t21 429.688
R340 B.n64 B.t10 429.688
R341 B.n72 B.t14 429.688
R342 B.n403 B.n50 256.663
R343 B.n405 B.n50 256.663
R344 B.n411 B.n50 256.663
R345 B.n413 B.n50 256.663
R346 B.n419 B.n50 256.663
R347 B.n421 B.n50 256.663
R348 B.n427 B.n50 256.663
R349 B.n429 B.n50 256.663
R350 B.n435 B.n50 256.663
R351 B.n437 B.n50 256.663
R352 B.n443 B.n50 256.663
R353 B.n445 B.n50 256.663
R354 B.n451 B.n50 256.663
R355 B.n453 B.n50 256.663
R356 B.n459 B.n50 256.663
R357 B.n461 B.n50 256.663
R358 B.n467 B.n50 256.663
R359 B.n469 B.n50 256.663
R360 B.n476 B.n50 256.663
R361 B.n478 B.n50 256.663
R362 B.n484 B.n50 256.663
R363 B.n486 B.n50 256.663
R364 B.n492 B.n50 256.663
R365 B.n494 B.n50 256.663
R366 B.n500 B.n50 256.663
R367 B.n502 B.n50 256.663
R368 B.n508 B.n50 256.663
R369 B.n510 B.n50 256.663
R370 B.n516 B.n50 256.663
R371 B.n518 B.n50 256.663
R372 B.n284 B.n134 256.663
R373 B.n137 B.n134 256.663
R374 B.n277 B.n134 256.663
R375 B.n271 B.n134 256.663
R376 B.n269 B.n134 256.663
R377 B.n263 B.n134 256.663
R378 B.n261 B.n134 256.663
R379 B.n255 B.n134 256.663
R380 B.n253 B.n134 256.663
R381 B.n247 B.n134 256.663
R382 B.n245 B.n134 256.663
R383 B.n239 B.n134 256.663
R384 B.n151 B.n134 256.663
R385 B.n233 B.n134 256.663
R386 B.n227 B.n134 256.663
R387 B.n225 B.n134 256.663
R388 B.n219 B.n134 256.663
R389 B.n159 B.n134 256.663
R390 B.n213 B.n134 256.663
R391 B.n207 B.n134 256.663
R392 B.n205 B.n134 256.663
R393 B.n199 B.n134 256.663
R394 B.n197 B.n134 256.663
R395 B.n191 B.n134 256.663
R396 B.n189 B.n134 256.663
R397 B.n183 B.n134 256.663
R398 B.n181 B.n134 256.663
R399 B.n175 B.n134 256.663
R400 B.n173 B.n134 256.663
R401 B.n289 B.n129 163.367
R402 B.n297 B.n129 163.367
R403 B.n297 B.n127 163.367
R404 B.n301 B.n127 163.367
R405 B.n301 B.n121 163.367
R406 B.n309 B.n121 163.367
R407 B.n309 B.n119 163.367
R408 B.n313 B.n119 163.367
R409 B.n313 B.n113 163.367
R410 B.n322 B.n113 163.367
R411 B.n322 B.n111 163.367
R412 B.n326 B.n111 163.367
R413 B.n326 B.n106 163.367
R414 B.n333 B.n106 163.367
R415 B.n333 B.n104 163.367
R416 B.n337 B.n104 163.367
R417 B.n337 B.n98 163.367
R418 B.n346 B.n98 163.367
R419 B.n346 B.n96 163.367
R420 B.n350 B.n96 163.367
R421 B.n350 B.n91 163.367
R422 B.n359 B.n91 163.367
R423 B.n359 B.n89 163.367
R424 B.n363 B.n89 163.367
R425 B.n363 B.n2 163.367
R426 B.n574 B.n2 163.367
R427 B.n574 B.n3 163.367
R428 B.n570 B.n3 163.367
R429 B.n570 B.n9 163.367
R430 B.n566 B.n9 163.367
R431 B.n566 B.n11 163.367
R432 B.n562 B.n11 163.367
R433 B.n562 B.n15 163.367
R434 B.n558 B.n15 163.367
R435 B.n558 B.n17 163.367
R436 B.n554 B.n17 163.367
R437 B.n554 B.n23 163.367
R438 B.n550 B.n23 163.367
R439 B.n550 B.n25 163.367
R440 B.n547 B.n25 163.367
R441 B.n547 B.n29 163.367
R442 B.n543 B.n29 163.367
R443 B.n543 B.n31 163.367
R444 B.n539 B.n31 163.367
R445 B.n539 B.n37 163.367
R446 B.n535 B.n37 163.367
R447 B.n535 B.n39 163.367
R448 B.n531 B.n39 163.367
R449 B.n531 B.n44 163.367
R450 B.n527 B.n44 163.367
R451 B.n527 B.n46 163.367
R452 B.n523 B.n46 163.367
R453 B.n285 B.n283 163.367
R454 B.n283 B.n282 163.367
R455 B.n279 B.n278 163.367
R456 B.n276 B.n139 163.367
R457 B.n272 B.n270 163.367
R458 B.n268 B.n141 163.367
R459 B.n264 B.n262 163.367
R460 B.n260 B.n143 163.367
R461 B.n256 B.n254 163.367
R462 B.n252 B.n145 163.367
R463 B.n248 B.n246 163.367
R464 B.n244 B.n147 163.367
R465 B.n240 B.n238 163.367
R466 B.n235 B.n234 163.367
R467 B.n232 B.n153 163.367
R468 B.n228 B.n226 163.367
R469 B.n224 B.n155 163.367
R470 B.n220 B.n218 163.367
R471 B.n215 B.n214 163.367
R472 B.n212 B.n161 163.367
R473 B.n208 B.n206 163.367
R474 B.n204 B.n163 163.367
R475 B.n200 B.n198 163.367
R476 B.n196 B.n165 163.367
R477 B.n192 B.n190 163.367
R478 B.n188 B.n167 163.367
R479 B.n184 B.n182 163.367
R480 B.n180 B.n169 163.367
R481 B.n176 B.n174 163.367
R482 B.n172 B.n133 163.367
R483 B.n291 B.n131 163.367
R484 B.n295 B.n131 163.367
R485 B.n295 B.n125 163.367
R486 B.n303 B.n125 163.367
R487 B.n303 B.n123 163.367
R488 B.n307 B.n123 163.367
R489 B.n307 B.n117 163.367
R490 B.n315 B.n117 163.367
R491 B.n315 B.n115 163.367
R492 B.n319 B.n115 163.367
R493 B.n319 B.n110 163.367
R494 B.n328 B.n110 163.367
R495 B.n328 B.n108 163.367
R496 B.n332 B.n108 163.367
R497 B.n332 B.n102 163.367
R498 B.n339 B.n102 163.367
R499 B.n339 B.n100 163.367
R500 B.n343 B.n100 163.367
R501 B.n343 B.n95 163.367
R502 B.n352 B.n95 163.367
R503 B.n352 B.n93 163.367
R504 B.n357 B.n93 163.367
R505 B.n357 B.n87 163.367
R506 B.n365 B.n87 163.367
R507 B.n366 B.n365 163.367
R508 B.n366 B.n5 163.367
R509 B.n6 B.n5 163.367
R510 B.n7 B.n6 163.367
R511 B.n371 B.n7 163.367
R512 B.n371 B.n12 163.367
R513 B.n13 B.n12 163.367
R514 B.n14 B.n13 163.367
R515 B.n376 B.n14 163.367
R516 B.n376 B.n19 163.367
R517 B.n20 B.n19 163.367
R518 B.n21 B.n20 163.367
R519 B.n381 B.n21 163.367
R520 B.n381 B.n26 163.367
R521 B.n27 B.n26 163.367
R522 B.n28 B.n27 163.367
R523 B.n386 B.n28 163.367
R524 B.n386 B.n33 163.367
R525 B.n34 B.n33 163.367
R526 B.n35 B.n34 163.367
R527 B.n391 B.n35 163.367
R528 B.n391 B.n40 163.367
R529 B.n41 B.n40 163.367
R530 B.n42 B.n41 163.367
R531 B.n396 B.n42 163.367
R532 B.n396 B.n47 163.367
R533 B.n48 B.n47 163.367
R534 B.n49 B.n48 163.367
R535 B.n519 B.n517 163.367
R536 B.n515 B.n53 163.367
R537 B.n511 B.n509 163.367
R538 B.n507 B.n55 163.367
R539 B.n503 B.n501 163.367
R540 B.n499 B.n57 163.367
R541 B.n495 B.n493 163.367
R542 B.n491 B.n59 163.367
R543 B.n487 B.n485 163.367
R544 B.n483 B.n61 163.367
R545 B.n479 B.n477 163.367
R546 B.n475 B.n63 163.367
R547 B.n470 B.n468 163.367
R548 B.n466 B.n67 163.367
R549 B.n462 B.n460 163.367
R550 B.n458 B.n69 163.367
R551 B.n454 B.n452 163.367
R552 B.n450 B.n71 163.367
R553 B.n446 B.n444 163.367
R554 B.n442 B.n76 163.367
R555 B.n438 B.n436 163.367
R556 B.n434 B.n78 163.367
R557 B.n430 B.n428 163.367
R558 B.n426 B.n80 163.367
R559 B.n422 B.n420 163.367
R560 B.n418 B.n82 163.367
R561 B.n414 B.n412 163.367
R562 B.n410 B.n84 163.367
R563 B.n406 B.n404 163.367
R564 B.n290 B.n134 112.216
R565 B.n524 B.n50 112.216
R566 B.n156 B.t20 94.066
R567 B.n72 B.t15 94.066
R568 B.n148 B.t23 94.0592
R569 B.n64 B.t12 94.0592
R570 B.n157 B.t19 74.4781
R571 B.n73 B.t16 74.4781
R572 B.n149 B.t22 74.4713
R573 B.n65 B.t13 74.4713
R574 B.n284 B.n135 71.676
R575 B.n282 B.n137 71.676
R576 B.n278 B.n277 71.676
R577 B.n271 B.n139 71.676
R578 B.n270 B.n269 71.676
R579 B.n263 B.n141 71.676
R580 B.n262 B.n261 71.676
R581 B.n255 B.n143 71.676
R582 B.n254 B.n253 71.676
R583 B.n247 B.n145 71.676
R584 B.n246 B.n245 71.676
R585 B.n239 B.n147 71.676
R586 B.n238 B.n151 71.676
R587 B.n234 B.n233 71.676
R588 B.n227 B.n153 71.676
R589 B.n226 B.n225 71.676
R590 B.n219 B.n155 71.676
R591 B.n218 B.n159 71.676
R592 B.n214 B.n213 71.676
R593 B.n207 B.n161 71.676
R594 B.n206 B.n205 71.676
R595 B.n199 B.n163 71.676
R596 B.n198 B.n197 71.676
R597 B.n191 B.n165 71.676
R598 B.n190 B.n189 71.676
R599 B.n183 B.n167 71.676
R600 B.n182 B.n181 71.676
R601 B.n175 B.n169 71.676
R602 B.n174 B.n173 71.676
R603 B.n518 B.n51 71.676
R604 B.n517 B.n516 71.676
R605 B.n510 B.n53 71.676
R606 B.n509 B.n508 71.676
R607 B.n502 B.n55 71.676
R608 B.n501 B.n500 71.676
R609 B.n494 B.n57 71.676
R610 B.n493 B.n492 71.676
R611 B.n486 B.n59 71.676
R612 B.n485 B.n484 71.676
R613 B.n478 B.n61 71.676
R614 B.n477 B.n476 71.676
R615 B.n469 B.n63 71.676
R616 B.n468 B.n467 71.676
R617 B.n461 B.n67 71.676
R618 B.n460 B.n459 71.676
R619 B.n453 B.n69 71.676
R620 B.n452 B.n451 71.676
R621 B.n445 B.n71 71.676
R622 B.n444 B.n443 71.676
R623 B.n437 B.n76 71.676
R624 B.n436 B.n435 71.676
R625 B.n429 B.n78 71.676
R626 B.n428 B.n427 71.676
R627 B.n421 B.n80 71.676
R628 B.n420 B.n419 71.676
R629 B.n413 B.n82 71.676
R630 B.n412 B.n411 71.676
R631 B.n405 B.n84 71.676
R632 B.n404 B.n403 71.676
R633 B.n403 B.n402 71.676
R634 B.n406 B.n405 71.676
R635 B.n411 B.n410 71.676
R636 B.n414 B.n413 71.676
R637 B.n419 B.n418 71.676
R638 B.n422 B.n421 71.676
R639 B.n427 B.n426 71.676
R640 B.n430 B.n429 71.676
R641 B.n435 B.n434 71.676
R642 B.n438 B.n437 71.676
R643 B.n443 B.n442 71.676
R644 B.n446 B.n445 71.676
R645 B.n451 B.n450 71.676
R646 B.n454 B.n453 71.676
R647 B.n459 B.n458 71.676
R648 B.n462 B.n461 71.676
R649 B.n467 B.n466 71.676
R650 B.n470 B.n469 71.676
R651 B.n476 B.n475 71.676
R652 B.n479 B.n478 71.676
R653 B.n484 B.n483 71.676
R654 B.n487 B.n486 71.676
R655 B.n492 B.n491 71.676
R656 B.n495 B.n494 71.676
R657 B.n500 B.n499 71.676
R658 B.n503 B.n502 71.676
R659 B.n508 B.n507 71.676
R660 B.n511 B.n510 71.676
R661 B.n516 B.n515 71.676
R662 B.n519 B.n518 71.676
R663 B.n285 B.n284 71.676
R664 B.n279 B.n137 71.676
R665 B.n277 B.n276 71.676
R666 B.n272 B.n271 71.676
R667 B.n269 B.n268 71.676
R668 B.n264 B.n263 71.676
R669 B.n261 B.n260 71.676
R670 B.n256 B.n255 71.676
R671 B.n253 B.n252 71.676
R672 B.n248 B.n247 71.676
R673 B.n245 B.n244 71.676
R674 B.n240 B.n239 71.676
R675 B.n235 B.n151 71.676
R676 B.n233 B.n232 71.676
R677 B.n228 B.n227 71.676
R678 B.n225 B.n224 71.676
R679 B.n220 B.n219 71.676
R680 B.n215 B.n159 71.676
R681 B.n213 B.n212 71.676
R682 B.n208 B.n207 71.676
R683 B.n205 B.n204 71.676
R684 B.n200 B.n199 71.676
R685 B.n197 B.n196 71.676
R686 B.n192 B.n191 71.676
R687 B.n189 B.n188 71.676
R688 B.n184 B.n183 71.676
R689 B.n181 B.n180 71.676
R690 B.n176 B.n175 71.676
R691 B.n173 B.n172 71.676
R692 B.n290 B.n130 64.1239
R693 B.n296 B.n130 64.1239
R694 B.n296 B.n126 64.1239
R695 B.n302 B.n126 64.1239
R696 B.n308 B.n122 64.1239
R697 B.n308 B.n118 64.1239
R698 B.n314 B.n118 64.1239
R699 B.n314 B.n114 64.1239
R700 B.n321 B.n114 64.1239
R701 B.n321 B.n320 64.1239
R702 B.n327 B.n107 64.1239
R703 B.t4 B.n107 64.1239
R704 B.t4 B.n103 64.1239
R705 B.n338 B.n103 64.1239
R706 B.n345 B.n99 64.1239
R707 B.n345 B.n344 64.1239
R708 B.n351 B.n92 64.1239
R709 B.n358 B.n92 64.1239
R710 B.n364 B.n88 64.1239
R711 B.n364 B.n4 64.1239
R712 B.n573 B.n4 64.1239
R713 B.n573 B.n572 64.1239
R714 B.n572 B.n571 64.1239
R715 B.n571 B.n8 64.1239
R716 B.n565 B.n564 64.1239
R717 B.n564 B.n563 64.1239
R718 B.n557 B.n18 64.1239
R719 B.n557 B.n556 64.1239
R720 B.n555 B.n22 64.1239
R721 B.t0 B.n22 64.1239
R722 B.t0 B.n549 64.1239
R723 B.n549 B.n548 64.1239
R724 B.n542 B.n32 64.1239
R725 B.n542 B.n541 64.1239
R726 B.n541 B.n540 64.1239
R727 B.n540 B.n36 64.1239
R728 B.n534 B.n36 64.1239
R729 B.n534 B.n533 64.1239
R730 B.n532 B.n43 64.1239
R731 B.n526 B.n43 64.1239
R732 B.n526 B.n525 64.1239
R733 B.n525 B.n524 64.1239
R734 B.n327 B.t7 62.238
R735 B.n338 B.t2 62.238
R736 B.t6 B.n555 62.238
R737 B.n548 B.t5 62.238
R738 B.n344 B.t3 60.352
R739 B.n18 B.t9 60.352
R740 B.n158 B.n157 59.5399
R741 B.n150 B.n149 59.5399
R742 B.n472 B.n65 59.5399
R743 B.n74 B.n73 59.5399
R744 B.n358 B.t1 58.466
R745 B.n565 B.t8 58.466
R746 B.n302 B.t18 54.694
R747 B.t11 B.n532 54.694
R748 B.n522 B.n521 30.7517
R749 B.n401 B.n400 30.7517
R750 B.n292 B.n132 30.7517
R751 B.n288 B.n287 30.7517
R752 B.n157 B.n156 19.5884
R753 B.n149 B.n148 19.5884
R754 B.n65 B.n64 19.5884
R755 B.n73 B.n72 19.5884
R756 B B.n575 18.0485
R757 B.n521 B.n520 10.6151
R758 B.n520 B.n52 10.6151
R759 B.n514 B.n52 10.6151
R760 B.n514 B.n513 10.6151
R761 B.n513 B.n512 10.6151
R762 B.n512 B.n54 10.6151
R763 B.n506 B.n54 10.6151
R764 B.n506 B.n505 10.6151
R765 B.n505 B.n504 10.6151
R766 B.n504 B.n56 10.6151
R767 B.n498 B.n56 10.6151
R768 B.n498 B.n497 10.6151
R769 B.n497 B.n496 10.6151
R770 B.n496 B.n58 10.6151
R771 B.n490 B.n58 10.6151
R772 B.n490 B.n489 10.6151
R773 B.n489 B.n488 10.6151
R774 B.n488 B.n60 10.6151
R775 B.n482 B.n60 10.6151
R776 B.n482 B.n481 10.6151
R777 B.n481 B.n480 10.6151
R778 B.n480 B.n62 10.6151
R779 B.n474 B.n62 10.6151
R780 B.n474 B.n473 10.6151
R781 B.n471 B.n66 10.6151
R782 B.n465 B.n66 10.6151
R783 B.n465 B.n464 10.6151
R784 B.n464 B.n463 10.6151
R785 B.n463 B.n68 10.6151
R786 B.n457 B.n68 10.6151
R787 B.n457 B.n456 10.6151
R788 B.n456 B.n455 10.6151
R789 B.n455 B.n70 10.6151
R790 B.n449 B.n448 10.6151
R791 B.n448 B.n447 10.6151
R792 B.n447 B.n75 10.6151
R793 B.n441 B.n75 10.6151
R794 B.n441 B.n440 10.6151
R795 B.n440 B.n439 10.6151
R796 B.n439 B.n77 10.6151
R797 B.n433 B.n77 10.6151
R798 B.n433 B.n432 10.6151
R799 B.n432 B.n431 10.6151
R800 B.n431 B.n79 10.6151
R801 B.n425 B.n79 10.6151
R802 B.n425 B.n424 10.6151
R803 B.n424 B.n423 10.6151
R804 B.n423 B.n81 10.6151
R805 B.n417 B.n81 10.6151
R806 B.n417 B.n416 10.6151
R807 B.n416 B.n415 10.6151
R808 B.n415 B.n83 10.6151
R809 B.n409 B.n83 10.6151
R810 B.n409 B.n408 10.6151
R811 B.n408 B.n407 10.6151
R812 B.n407 B.n85 10.6151
R813 B.n401 B.n85 10.6151
R814 B.n293 B.n292 10.6151
R815 B.n294 B.n293 10.6151
R816 B.n294 B.n124 10.6151
R817 B.n304 B.n124 10.6151
R818 B.n305 B.n304 10.6151
R819 B.n306 B.n305 10.6151
R820 B.n306 B.n116 10.6151
R821 B.n316 B.n116 10.6151
R822 B.n317 B.n316 10.6151
R823 B.n318 B.n317 10.6151
R824 B.n318 B.n109 10.6151
R825 B.n329 B.n109 10.6151
R826 B.n330 B.n329 10.6151
R827 B.n331 B.n330 10.6151
R828 B.n331 B.n101 10.6151
R829 B.n340 B.n101 10.6151
R830 B.n341 B.n340 10.6151
R831 B.n342 B.n341 10.6151
R832 B.n342 B.n94 10.6151
R833 B.n353 B.n94 10.6151
R834 B.n354 B.n353 10.6151
R835 B.n356 B.n354 10.6151
R836 B.n356 B.n355 10.6151
R837 B.n355 B.n86 10.6151
R838 B.n367 B.n86 10.6151
R839 B.n368 B.n367 10.6151
R840 B.n369 B.n368 10.6151
R841 B.n370 B.n369 10.6151
R842 B.n372 B.n370 10.6151
R843 B.n373 B.n372 10.6151
R844 B.n374 B.n373 10.6151
R845 B.n375 B.n374 10.6151
R846 B.n377 B.n375 10.6151
R847 B.n378 B.n377 10.6151
R848 B.n379 B.n378 10.6151
R849 B.n380 B.n379 10.6151
R850 B.n382 B.n380 10.6151
R851 B.n383 B.n382 10.6151
R852 B.n384 B.n383 10.6151
R853 B.n385 B.n384 10.6151
R854 B.n387 B.n385 10.6151
R855 B.n388 B.n387 10.6151
R856 B.n389 B.n388 10.6151
R857 B.n390 B.n389 10.6151
R858 B.n392 B.n390 10.6151
R859 B.n393 B.n392 10.6151
R860 B.n394 B.n393 10.6151
R861 B.n395 B.n394 10.6151
R862 B.n397 B.n395 10.6151
R863 B.n398 B.n397 10.6151
R864 B.n399 B.n398 10.6151
R865 B.n400 B.n399 10.6151
R866 B.n287 B.n286 10.6151
R867 B.n286 B.n136 10.6151
R868 B.n281 B.n136 10.6151
R869 B.n281 B.n280 10.6151
R870 B.n280 B.n138 10.6151
R871 B.n275 B.n138 10.6151
R872 B.n275 B.n274 10.6151
R873 B.n274 B.n273 10.6151
R874 B.n273 B.n140 10.6151
R875 B.n267 B.n140 10.6151
R876 B.n267 B.n266 10.6151
R877 B.n266 B.n265 10.6151
R878 B.n265 B.n142 10.6151
R879 B.n259 B.n142 10.6151
R880 B.n259 B.n258 10.6151
R881 B.n258 B.n257 10.6151
R882 B.n257 B.n144 10.6151
R883 B.n251 B.n144 10.6151
R884 B.n251 B.n250 10.6151
R885 B.n250 B.n249 10.6151
R886 B.n249 B.n146 10.6151
R887 B.n243 B.n146 10.6151
R888 B.n243 B.n242 10.6151
R889 B.n242 B.n241 10.6151
R890 B.n237 B.n236 10.6151
R891 B.n236 B.n152 10.6151
R892 B.n231 B.n152 10.6151
R893 B.n231 B.n230 10.6151
R894 B.n230 B.n229 10.6151
R895 B.n229 B.n154 10.6151
R896 B.n223 B.n154 10.6151
R897 B.n223 B.n222 10.6151
R898 B.n222 B.n221 10.6151
R899 B.n217 B.n216 10.6151
R900 B.n216 B.n160 10.6151
R901 B.n211 B.n160 10.6151
R902 B.n211 B.n210 10.6151
R903 B.n210 B.n209 10.6151
R904 B.n209 B.n162 10.6151
R905 B.n203 B.n162 10.6151
R906 B.n203 B.n202 10.6151
R907 B.n202 B.n201 10.6151
R908 B.n201 B.n164 10.6151
R909 B.n195 B.n164 10.6151
R910 B.n195 B.n194 10.6151
R911 B.n194 B.n193 10.6151
R912 B.n193 B.n166 10.6151
R913 B.n187 B.n166 10.6151
R914 B.n187 B.n186 10.6151
R915 B.n186 B.n185 10.6151
R916 B.n185 B.n168 10.6151
R917 B.n179 B.n168 10.6151
R918 B.n179 B.n178 10.6151
R919 B.n178 B.n177 10.6151
R920 B.n177 B.n170 10.6151
R921 B.n171 B.n170 10.6151
R922 B.n171 B.n132 10.6151
R923 B.n288 B.n128 10.6151
R924 B.n298 B.n128 10.6151
R925 B.n299 B.n298 10.6151
R926 B.n300 B.n299 10.6151
R927 B.n300 B.n120 10.6151
R928 B.n310 B.n120 10.6151
R929 B.n311 B.n310 10.6151
R930 B.n312 B.n311 10.6151
R931 B.n312 B.n112 10.6151
R932 B.n323 B.n112 10.6151
R933 B.n324 B.n323 10.6151
R934 B.n325 B.n324 10.6151
R935 B.n325 B.n105 10.6151
R936 B.n334 B.n105 10.6151
R937 B.n335 B.n334 10.6151
R938 B.n336 B.n335 10.6151
R939 B.n336 B.n97 10.6151
R940 B.n347 B.n97 10.6151
R941 B.n348 B.n347 10.6151
R942 B.n349 B.n348 10.6151
R943 B.n349 B.n90 10.6151
R944 B.n360 B.n90 10.6151
R945 B.n361 B.n360 10.6151
R946 B.n362 B.n361 10.6151
R947 B.n362 B.n0 10.6151
R948 B.n569 B.n1 10.6151
R949 B.n569 B.n568 10.6151
R950 B.n568 B.n567 10.6151
R951 B.n567 B.n10 10.6151
R952 B.n561 B.n10 10.6151
R953 B.n561 B.n560 10.6151
R954 B.n560 B.n559 10.6151
R955 B.n559 B.n16 10.6151
R956 B.n553 B.n16 10.6151
R957 B.n553 B.n552 10.6151
R958 B.n552 B.n551 10.6151
R959 B.n551 B.n24 10.6151
R960 B.n546 B.n24 10.6151
R961 B.n546 B.n545 10.6151
R962 B.n545 B.n544 10.6151
R963 B.n544 B.n30 10.6151
R964 B.n538 B.n30 10.6151
R965 B.n538 B.n537 10.6151
R966 B.n537 B.n536 10.6151
R967 B.n536 B.n38 10.6151
R968 B.n530 B.n38 10.6151
R969 B.n530 B.n529 10.6151
R970 B.n529 B.n528 10.6151
R971 B.n528 B.n45 10.6151
R972 B.n522 B.n45 10.6151
R973 B.t18 B.n122 9.43042
R974 B.n533 B.t11 9.43042
R975 B.n473 B.n472 9.36635
R976 B.n449 B.n74 9.36635
R977 B.n241 B.n150 9.36635
R978 B.n217 B.n158 9.36635
R979 B.t1 B.n88 5.65845
R980 B.t8 B.n8 5.65845
R981 B.n351 B.t3 3.77247
R982 B.n563 B.t9 3.77247
R983 B.n575 B.n0 2.81026
R984 B.n575 B.n1 2.81026
R985 B.n320 B.t7 1.88648
R986 B.t2 B.n99 1.88648
R987 B.n556 B.t6 1.88648
R988 B.n32 B.t5 1.88648
R989 B.n472 B.n471 1.24928
R990 B.n74 B.n70 1.24928
R991 B.n237 B.n150 1.24928
R992 B.n221 B.n158 1.24928
R993 VN.n3 VN.t8 306.188
R994 VN.n17 VN.t7 306.188
R995 VN.n4 VN.t1 284.594
R996 VN.n6 VN.t0 284.594
R997 VN.n10 VN.t3 284.594
R998 VN.n12 VN.t5 284.594
R999 VN.n18 VN.t4 284.594
R1000 VN.n20 VN.t2 284.594
R1001 VN.n24 VN.t9 284.594
R1002 VN.n26 VN.t6 284.594
R1003 VN.n13 VN.n12 161.3
R1004 VN.n27 VN.n26 161.3
R1005 VN.n25 VN.n14 161.3
R1006 VN.n24 VN.n23 161.3
R1007 VN.n22 VN.n15 161.3
R1008 VN.n21 VN.n20 161.3
R1009 VN.n19 VN.n16 161.3
R1010 VN.n11 VN.n0 161.3
R1011 VN.n10 VN.n9 161.3
R1012 VN.n8 VN.n1 161.3
R1013 VN.n7 VN.n6 161.3
R1014 VN.n5 VN.n2 161.3
R1015 VN.n17 VN.n16 44.8545
R1016 VN.n3 VN.n2 44.8545
R1017 VN VN.n27 38.7713
R1018 VN.n12 VN.n11 26.2914
R1019 VN.n26 VN.n25 26.2914
R1020 VN.n5 VN.n4 24.8308
R1021 VN.n10 VN.n1 24.8308
R1022 VN.n19 VN.n18 24.8308
R1023 VN.n24 VN.n15 24.8308
R1024 VN.n6 VN.n5 23.3702
R1025 VN.n6 VN.n1 23.3702
R1026 VN.n20 VN.n19 23.3702
R1027 VN.n20 VN.n15 23.3702
R1028 VN.n11 VN.n10 21.9096
R1029 VN.n25 VN.n24 21.9096
R1030 VN.n4 VN.n3 20.3348
R1031 VN.n18 VN.n17 20.3348
R1032 VN.n27 VN.n14 0.189894
R1033 VN.n23 VN.n14 0.189894
R1034 VN.n23 VN.n22 0.189894
R1035 VN.n22 VN.n21 0.189894
R1036 VN.n21 VN.n16 0.189894
R1037 VN.n7 VN.n2 0.189894
R1038 VN.n8 VN.n7 0.189894
R1039 VN.n9 VN.n8 0.189894
R1040 VN.n9 VN.n0 0.189894
R1041 VN.n13 VN.n0 0.189894
R1042 VN VN.n13 0.0516364
R1043 VTAIL.n11 VTAIL.t13 53.5976
R1044 VTAIL.n16 VTAIL.t19 53.5975
R1045 VTAIL.n17 VTAIL.t12 53.5975
R1046 VTAIL.n2 VTAIL.t2 53.5975
R1047 VTAIL.n15 VTAIL.n14 50.4991
R1048 VTAIL.n13 VTAIL.n12 50.4991
R1049 VTAIL.n10 VTAIL.n9 50.4991
R1050 VTAIL.n8 VTAIL.n7 50.4991
R1051 VTAIL.n19 VTAIL.n18 50.4989
R1052 VTAIL.n1 VTAIL.n0 50.4989
R1053 VTAIL.n4 VTAIL.n3 50.4989
R1054 VTAIL.n6 VTAIL.n5 50.4989
R1055 VTAIL.n8 VTAIL.n6 19.6169
R1056 VTAIL.n17 VTAIL.n16 18.7462
R1057 VTAIL.n18 VTAIL.t11 3.09909
R1058 VTAIL.n18 VTAIL.t4 3.09909
R1059 VTAIL.n0 VTAIL.t7 3.09909
R1060 VTAIL.n0 VTAIL.t5 3.09909
R1061 VTAIL.n3 VTAIL.t0 3.09909
R1062 VTAIL.n3 VTAIL.t1 3.09909
R1063 VTAIL.n5 VTAIL.t18 3.09909
R1064 VTAIL.n5 VTAIL.t17 3.09909
R1065 VTAIL.n14 VTAIL.t3 3.09909
R1066 VTAIL.n14 VTAIL.t16 3.09909
R1067 VTAIL.n12 VTAIL.t14 3.09909
R1068 VTAIL.n12 VTAIL.t15 3.09909
R1069 VTAIL.n9 VTAIL.t9 3.09909
R1070 VTAIL.n9 VTAIL.t6 3.09909
R1071 VTAIL.n7 VTAIL.t10 3.09909
R1072 VTAIL.n7 VTAIL.t8 3.09909
R1073 VTAIL.n13 VTAIL.n11 0.905672
R1074 VTAIL.n2 VTAIL.n1 0.905672
R1075 VTAIL.n10 VTAIL.n8 0.87119
R1076 VTAIL.n11 VTAIL.n10 0.87119
R1077 VTAIL.n15 VTAIL.n13 0.87119
R1078 VTAIL.n16 VTAIL.n15 0.87119
R1079 VTAIL.n6 VTAIL.n4 0.87119
R1080 VTAIL.n4 VTAIL.n2 0.87119
R1081 VTAIL.n19 VTAIL.n17 0.87119
R1082 VTAIL VTAIL.n1 0.711707
R1083 VTAIL VTAIL.n19 0.159983
R1084 VDD2.n1 VDD2.t1 71.147
R1085 VDD2.n4 VDD2.t3 70.2764
R1086 VDD2.n3 VDD2.n2 67.7753
R1087 VDD2 VDD2.n7 67.7725
R1088 VDD2.n6 VDD2.n5 67.1779
R1089 VDD2.n1 VDD2.n0 67.1777
R1090 VDD2.n4 VDD2.n3 33.3597
R1091 VDD2.n7 VDD2.t5 3.09909
R1092 VDD2.n7 VDD2.t2 3.09909
R1093 VDD2.n5 VDD2.t0 3.09909
R1094 VDD2.n5 VDD2.t7 3.09909
R1095 VDD2.n2 VDD2.t6 3.09909
R1096 VDD2.n2 VDD2.t4 3.09909
R1097 VDD2.n0 VDD2.t8 3.09909
R1098 VDD2.n0 VDD2.t9 3.09909
R1099 VDD2.n6 VDD2.n4 0.87119
R1100 VDD2 VDD2.n6 0.276362
R1101 VDD2.n3 VDD2.n1 0.162826
R1102 VP.n7 VP.t4 306.188
R1103 VP.n18 VP.t7 284.594
R1104 VP.n22 VP.t8 284.594
R1105 VP.n24 VP.t5 284.594
R1106 VP.n28 VP.t2 284.594
R1107 VP.n30 VP.t0 284.594
R1108 VP.n16 VP.t3 284.594
R1109 VP.n14 VP.t6 284.594
R1110 VP.n6 VP.t9 284.594
R1111 VP.n8 VP.t1 284.594
R1112 VP.n31 VP.n30 161.3
R1113 VP.n10 VP.n9 161.3
R1114 VP.n11 VP.n6 161.3
R1115 VP.n13 VP.n12 161.3
R1116 VP.n14 VP.n5 161.3
R1117 VP.n15 VP.n4 161.3
R1118 VP.n17 VP.n16 161.3
R1119 VP.n29 VP.n0 161.3
R1120 VP.n28 VP.n27 161.3
R1121 VP.n26 VP.n1 161.3
R1122 VP.n25 VP.n24 161.3
R1123 VP.n23 VP.n2 161.3
R1124 VP.n22 VP.n21 161.3
R1125 VP.n20 VP.n3 161.3
R1126 VP.n19 VP.n18 161.3
R1127 VP.n10 VP.n7 44.8545
R1128 VP.n19 VP.n17 38.3907
R1129 VP.n18 VP.n3 26.2914
R1130 VP.n30 VP.n29 26.2914
R1131 VP.n16 VP.n15 26.2914
R1132 VP.n23 VP.n22 24.8308
R1133 VP.n28 VP.n1 24.8308
R1134 VP.n14 VP.n13 24.8308
R1135 VP.n9 VP.n8 24.8308
R1136 VP.n24 VP.n23 23.3702
R1137 VP.n24 VP.n1 23.3702
R1138 VP.n13 VP.n6 23.3702
R1139 VP.n9 VP.n6 23.3702
R1140 VP.n22 VP.n3 21.9096
R1141 VP.n29 VP.n28 21.9096
R1142 VP.n15 VP.n14 21.9096
R1143 VP.n8 VP.n7 20.3348
R1144 VP.n11 VP.n10 0.189894
R1145 VP.n12 VP.n11 0.189894
R1146 VP.n12 VP.n5 0.189894
R1147 VP.n5 VP.n4 0.189894
R1148 VP.n17 VP.n4 0.189894
R1149 VP.n20 VP.n19 0.189894
R1150 VP.n21 VP.n20 0.189894
R1151 VP.n21 VP.n2 0.189894
R1152 VP.n25 VP.n2 0.189894
R1153 VP.n26 VP.n25 0.189894
R1154 VP.n27 VP.n26 0.189894
R1155 VP.n27 VP.n0 0.189894
R1156 VP.n31 VP.n0 0.189894
R1157 VP VP.n31 0.0516364
R1158 VDD1.n1 VDD1.t5 71.1471
R1159 VDD1.n3 VDD1.t2 71.147
R1160 VDD1.n5 VDD1.n4 67.7753
R1161 VDD1.n1 VDD1.n0 67.1779
R1162 VDD1.n7 VDD1.n6 67.1777
R1163 VDD1.n3 VDD1.n2 67.1777
R1164 VDD1.n7 VDD1.n5 34.378
R1165 VDD1.n6 VDD1.t3 3.09909
R1166 VDD1.n6 VDD1.t6 3.09909
R1167 VDD1.n0 VDD1.t8 3.09909
R1168 VDD1.n0 VDD1.t0 3.09909
R1169 VDD1.n4 VDD1.t7 3.09909
R1170 VDD1.n4 VDD1.t9 3.09909
R1171 VDD1.n2 VDD1.t1 3.09909
R1172 VDD1.n2 VDD1.t4 3.09909
R1173 VDD1 VDD1.n7 0.595328
R1174 VDD1 VDD1.n1 0.276362
R1175 VDD1.n5 VDD1.n3 0.162826
C0 VN VP 4.53132f
C1 VDD1 VN 0.148533f
C2 VTAIL VDD2 8.87f
C3 VTAIL VP 3.84592f
C4 VDD1 VTAIL 8.83287f
C5 VP VDD2 0.337737f
C6 VDD1 VDD2 0.955335f
C7 VDD1 VP 3.90621f
C8 VTAIL VN 3.83154f
C9 VN VDD2 3.71978f
C10 VDD2 B 3.94309f
C11 VDD1 B 3.866373f
C12 VTAIL B 4.284023f
C13 VN B 8.64116f
C14 VP B 6.94668f
C15 VDD1.t5 B 1.3365f
C16 VDD1.t8 B 0.1247f
C17 VDD1.t0 B 0.1247f
C18 VDD1.n0 B 1.048f
C19 VDD1.n1 B 0.624798f
C20 VDD1.t2 B 1.3365f
C21 VDD1.t1 B 0.1247f
C22 VDD1.t4 B 0.1247f
C23 VDD1.n2 B 1.048f
C24 VDD1.n3 B 0.6193f
C25 VDD1.t7 B 0.1247f
C26 VDD1.t9 B 0.1247f
C27 VDD1.n4 B 1.0509f
C28 VDD1.n5 B 1.61101f
C29 VDD1.t3 B 0.1247f
C30 VDD1.t6 B 0.1247f
C31 VDD1.n6 B 1.04799f
C32 VDD1.n7 B 1.91013f
C33 VP.n0 B 0.044746f
C34 VP.n1 B 0.010154f
C35 VP.n2 B 0.044746f
C36 VP.n3 B 0.010154f
C37 VP.n4 B 0.044746f
C38 VP.t3 B 0.563079f
C39 VP.t6 B 0.563079f
C40 VP.n5 B 0.044746f
C41 VP.t9 B 0.563079f
C42 VP.n6 B 0.256883f
C43 VP.t4 B 0.581137f
C44 VP.n7 B 0.242387f
C45 VP.t1 B 0.563079f
C46 VP.n8 B 0.260505f
C47 VP.n9 B 0.010154f
C48 VP.n10 B 0.184162f
C49 VP.n11 B 0.044746f
C50 VP.n12 B 0.044746f
C51 VP.n13 B 0.010154f
C52 VP.n14 B 0.256883f
C53 VP.n15 B 0.010154f
C54 VP.n16 B 0.25302f
C55 VP.n17 B 1.58231f
C56 VP.t7 B 0.563079f
C57 VP.n18 B 0.25302f
C58 VP.n19 B 1.62421f
C59 VP.n20 B 0.044746f
C60 VP.n21 B 0.044746f
C61 VP.t8 B 0.563079f
C62 VP.n22 B 0.256883f
C63 VP.n23 B 0.010154f
C64 VP.t5 B 0.563079f
C65 VP.n24 B 0.256883f
C66 VP.n25 B 0.044746f
C67 VP.n26 B 0.044746f
C68 VP.n27 B 0.044746f
C69 VP.t2 B 0.563079f
C70 VP.n28 B 0.256883f
C71 VP.n29 B 0.010154f
C72 VP.t0 B 0.563079f
C73 VP.n30 B 0.25302f
C74 VP.n31 B 0.034677f
C75 VDD2.t1 B 1.33556f
C76 VDD2.t8 B 0.124613f
C77 VDD2.t9 B 0.124613f
C78 VDD2.n0 B 1.04727f
C79 VDD2.n1 B 0.618869f
C80 VDD2.t6 B 0.124613f
C81 VDD2.t4 B 0.124613f
C82 VDD2.n2 B 1.05017f
C83 VDD2.n3 B 1.5365f
C84 VDD2.t3 B 1.33146f
C85 VDD2.n4 B 1.8994f
C86 VDD2.t0 B 0.124613f
C87 VDD2.t7 B 0.124613f
C88 VDD2.n5 B 1.04727f
C89 VDD2.n6 B 0.292403f
C90 VDD2.t5 B 0.124613f
C91 VDD2.t2 B 0.124613f
C92 VDD2.n7 B 1.05014f
C93 VTAIL.t7 B 0.138053f
C94 VTAIL.t5 B 0.138053f
C95 VTAIL.n0 B 1.08831f
C96 VTAIL.n1 B 0.40009f
C97 VTAIL.t2 B 1.38811f
C98 VTAIL.n2 B 0.490845f
C99 VTAIL.t0 B 0.138053f
C100 VTAIL.t1 B 0.138053f
C101 VTAIL.n3 B 1.08831f
C102 VTAIL.n4 B 0.411102f
C103 VTAIL.t18 B 0.138053f
C104 VTAIL.t17 B 0.138053f
C105 VTAIL.n5 B 1.08831f
C106 VTAIL.n6 B 1.34446f
C107 VTAIL.t10 B 0.138053f
C108 VTAIL.t8 B 0.138053f
C109 VTAIL.n7 B 1.08831f
C110 VTAIL.n8 B 1.34445f
C111 VTAIL.t9 B 0.138053f
C112 VTAIL.t6 B 0.138053f
C113 VTAIL.n9 B 1.08831f
C114 VTAIL.n10 B 0.411096f
C115 VTAIL.t13 B 1.38812f
C116 VTAIL.n11 B 0.490837f
C117 VTAIL.t14 B 0.138053f
C118 VTAIL.t15 B 0.138053f
C119 VTAIL.n12 B 1.08831f
C120 VTAIL.n13 B 0.414134f
C121 VTAIL.t3 B 0.138053f
C122 VTAIL.t16 B 0.138053f
C123 VTAIL.n14 B 1.08831f
C124 VTAIL.n15 B 0.411096f
C125 VTAIL.t19 B 1.38811f
C126 VTAIL.n16 B 1.34446f
C127 VTAIL.t12 B 1.38811f
C128 VTAIL.n17 B 1.34446f
C129 VTAIL.t11 B 0.138053f
C130 VTAIL.t4 B 0.138053f
C131 VTAIL.n18 B 1.08831f
C132 VTAIL.n19 B 0.348449f
C133 VN.n0 B 0.043787f
C134 VN.n1 B 0.009936f
C135 VN.n2 B 0.180214f
C136 VN.t8 B 0.568678f
C137 VN.n3 B 0.237191f
C138 VN.t1 B 0.551008f
C139 VN.n4 B 0.25492f
C140 VN.n5 B 0.009936f
C141 VN.t0 B 0.551008f
C142 VN.n6 B 0.251375f
C143 VN.n7 B 0.043787f
C144 VN.n8 B 0.043787f
C145 VN.n9 B 0.043787f
C146 VN.t3 B 0.551008f
C147 VN.n10 B 0.251375f
C148 VN.n11 B 0.009936f
C149 VN.t5 B 0.551008f
C150 VN.n12 B 0.247596f
C151 VN.n13 B 0.033933f
C152 VN.n14 B 0.043787f
C153 VN.n15 B 0.009936f
C154 VN.t9 B 0.551008f
C155 VN.n16 B 0.180214f
C156 VN.t7 B 0.568678f
C157 VN.n17 B 0.237191f
C158 VN.t4 B 0.551008f
C159 VN.n18 B 0.25492f
C160 VN.n19 B 0.009936f
C161 VN.t2 B 0.551008f
C162 VN.n20 B 0.251375f
C163 VN.n21 B 0.043787f
C164 VN.n22 B 0.043787f
C165 VN.n23 B 0.043787f
C166 VN.n24 B 0.251375f
C167 VN.n25 B 0.009936f
C168 VN.t6 B 0.551008f
C169 VN.n26 B 0.247596f
C170 VN.n27 B 1.5773f
.ends

