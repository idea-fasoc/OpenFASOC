* NGSPICE file created from diff_pair_sample_1555.ext - technology: sky130A

.subckt diff_pair_sample_1555 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=0 ps=0 w=10.66 l=3.57
X1 VTAIL.t11 VN.t0 VDD2.t1 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=1.7589 ps=10.99 w=10.66 l=3.57
X2 VDD1.t5 VP.t0 VTAIL.t0 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=4.1574 ps=22.1 w=10.66 l=3.57
X3 B.t8 B.t6 B.t7 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=0 ps=0 w=10.66 l=3.57
X4 B.t5 B.t3 B.t4 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=0 ps=0 w=10.66 l=3.57
X5 VDD2.t3 VN.t1 VTAIL.t10 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=1.7589 ps=10.99 w=10.66 l=3.57
X6 VDD2.t2 VN.t2 VTAIL.t9 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=4.1574 ps=22.1 w=10.66 l=3.57
X7 VDD1.t4 VP.t1 VTAIL.t5 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=1.7589 ps=10.99 w=10.66 l=3.57
X8 VTAIL.t8 VN.t3 VDD2.t5 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=1.7589 ps=10.99 w=10.66 l=3.57
X9 VDD1.t3 VP.t2 VTAIL.t4 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=4.1574 ps=22.1 w=10.66 l=3.57
X10 VDD1.t2 VP.t3 VTAIL.t1 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=1.7589 ps=10.99 w=10.66 l=3.57
X11 VDD2.t4 VN.t4 VTAIL.t7 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=4.1574 ps=22.1 w=10.66 l=3.57
X12 VTAIL.t2 VP.t4 VDD1.t1 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=1.7589 ps=10.99 w=10.66 l=3.57
X13 VDD2.t0 VN.t5 VTAIL.t6 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=1.7589 ps=10.99 w=10.66 l=3.57
X14 VTAIL.t3 VP.t5 VDD1.t0 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=10.99 as=1.7589 ps=10.99 w=10.66 l=3.57
X15 B.t2 B.t0 B.t1 w_n4090_n3100# sky130_fd_pr__pfet_01v8 ad=4.1574 pd=22.1 as=0 ps=0 w=10.66 l=3.57
R0 B.n577 B.n576 585
R1 B.n578 B.n75 585
R2 B.n580 B.n579 585
R3 B.n581 B.n74 585
R4 B.n583 B.n582 585
R5 B.n584 B.n73 585
R6 B.n586 B.n585 585
R7 B.n587 B.n72 585
R8 B.n589 B.n588 585
R9 B.n590 B.n71 585
R10 B.n592 B.n591 585
R11 B.n593 B.n70 585
R12 B.n595 B.n594 585
R13 B.n596 B.n69 585
R14 B.n598 B.n597 585
R15 B.n599 B.n68 585
R16 B.n601 B.n600 585
R17 B.n602 B.n67 585
R18 B.n604 B.n603 585
R19 B.n605 B.n66 585
R20 B.n607 B.n606 585
R21 B.n608 B.n65 585
R22 B.n610 B.n609 585
R23 B.n611 B.n64 585
R24 B.n613 B.n612 585
R25 B.n614 B.n63 585
R26 B.n616 B.n615 585
R27 B.n617 B.n62 585
R28 B.n619 B.n618 585
R29 B.n620 B.n61 585
R30 B.n622 B.n621 585
R31 B.n623 B.n60 585
R32 B.n625 B.n624 585
R33 B.n626 B.n59 585
R34 B.n628 B.n627 585
R35 B.n629 B.n58 585
R36 B.n631 B.n630 585
R37 B.n632 B.n55 585
R38 B.n635 B.n634 585
R39 B.n636 B.n54 585
R40 B.n638 B.n637 585
R41 B.n639 B.n53 585
R42 B.n641 B.n640 585
R43 B.n642 B.n52 585
R44 B.n644 B.n643 585
R45 B.n645 B.n51 585
R46 B.n647 B.n646 585
R47 B.n649 B.n648 585
R48 B.n650 B.n47 585
R49 B.n652 B.n651 585
R50 B.n653 B.n46 585
R51 B.n655 B.n654 585
R52 B.n656 B.n45 585
R53 B.n658 B.n657 585
R54 B.n659 B.n44 585
R55 B.n661 B.n660 585
R56 B.n662 B.n43 585
R57 B.n664 B.n663 585
R58 B.n665 B.n42 585
R59 B.n667 B.n666 585
R60 B.n668 B.n41 585
R61 B.n670 B.n669 585
R62 B.n671 B.n40 585
R63 B.n673 B.n672 585
R64 B.n674 B.n39 585
R65 B.n676 B.n675 585
R66 B.n677 B.n38 585
R67 B.n679 B.n678 585
R68 B.n680 B.n37 585
R69 B.n682 B.n681 585
R70 B.n683 B.n36 585
R71 B.n685 B.n684 585
R72 B.n686 B.n35 585
R73 B.n688 B.n687 585
R74 B.n689 B.n34 585
R75 B.n691 B.n690 585
R76 B.n692 B.n33 585
R77 B.n694 B.n693 585
R78 B.n695 B.n32 585
R79 B.n697 B.n696 585
R80 B.n698 B.n31 585
R81 B.n700 B.n699 585
R82 B.n701 B.n30 585
R83 B.n703 B.n702 585
R84 B.n704 B.n29 585
R85 B.n575 B.n76 585
R86 B.n574 B.n573 585
R87 B.n572 B.n77 585
R88 B.n571 B.n570 585
R89 B.n569 B.n78 585
R90 B.n568 B.n567 585
R91 B.n566 B.n79 585
R92 B.n565 B.n564 585
R93 B.n563 B.n80 585
R94 B.n562 B.n561 585
R95 B.n560 B.n81 585
R96 B.n559 B.n558 585
R97 B.n557 B.n82 585
R98 B.n556 B.n555 585
R99 B.n554 B.n83 585
R100 B.n553 B.n552 585
R101 B.n551 B.n84 585
R102 B.n550 B.n549 585
R103 B.n548 B.n85 585
R104 B.n547 B.n546 585
R105 B.n545 B.n86 585
R106 B.n544 B.n543 585
R107 B.n542 B.n87 585
R108 B.n541 B.n540 585
R109 B.n539 B.n88 585
R110 B.n538 B.n537 585
R111 B.n536 B.n89 585
R112 B.n535 B.n534 585
R113 B.n533 B.n90 585
R114 B.n532 B.n531 585
R115 B.n530 B.n91 585
R116 B.n529 B.n528 585
R117 B.n527 B.n92 585
R118 B.n526 B.n525 585
R119 B.n524 B.n93 585
R120 B.n523 B.n522 585
R121 B.n521 B.n94 585
R122 B.n520 B.n519 585
R123 B.n518 B.n95 585
R124 B.n517 B.n516 585
R125 B.n515 B.n96 585
R126 B.n514 B.n513 585
R127 B.n512 B.n97 585
R128 B.n511 B.n510 585
R129 B.n509 B.n98 585
R130 B.n508 B.n507 585
R131 B.n506 B.n99 585
R132 B.n505 B.n504 585
R133 B.n503 B.n100 585
R134 B.n502 B.n501 585
R135 B.n500 B.n101 585
R136 B.n499 B.n498 585
R137 B.n497 B.n102 585
R138 B.n496 B.n495 585
R139 B.n494 B.n103 585
R140 B.n493 B.n492 585
R141 B.n491 B.n104 585
R142 B.n490 B.n489 585
R143 B.n488 B.n105 585
R144 B.n487 B.n486 585
R145 B.n485 B.n106 585
R146 B.n484 B.n483 585
R147 B.n482 B.n107 585
R148 B.n481 B.n480 585
R149 B.n479 B.n108 585
R150 B.n478 B.n477 585
R151 B.n476 B.n109 585
R152 B.n475 B.n474 585
R153 B.n473 B.n110 585
R154 B.n472 B.n471 585
R155 B.n470 B.n111 585
R156 B.n469 B.n468 585
R157 B.n467 B.n112 585
R158 B.n466 B.n465 585
R159 B.n464 B.n113 585
R160 B.n463 B.n462 585
R161 B.n461 B.n114 585
R162 B.n460 B.n459 585
R163 B.n458 B.n115 585
R164 B.n457 B.n456 585
R165 B.n455 B.n116 585
R166 B.n454 B.n453 585
R167 B.n452 B.n117 585
R168 B.n451 B.n450 585
R169 B.n449 B.n118 585
R170 B.n448 B.n447 585
R171 B.n446 B.n119 585
R172 B.n445 B.n444 585
R173 B.n443 B.n120 585
R174 B.n442 B.n441 585
R175 B.n440 B.n121 585
R176 B.n439 B.n438 585
R177 B.n437 B.n122 585
R178 B.n436 B.n435 585
R179 B.n434 B.n123 585
R180 B.n433 B.n432 585
R181 B.n431 B.n124 585
R182 B.n430 B.n429 585
R183 B.n428 B.n125 585
R184 B.n427 B.n426 585
R185 B.n425 B.n126 585
R186 B.n424 B.n423 585
R187 B.n422 B.n127 585
R188 B.n421 B.n420 585
R189 B.n419 B.n128 585
R190 B.n418 B.n417 585
R191 B.n416 B.n129 585
R192 B.n415 B.n414 585
R193 B.n413 B.n130 585
R194 B.n284 B.n177 585
R195 B.n286 B.n285 585
R196 B.n287 B.n176 585
R197 B.n289 B.n288 585
R198 B.n290 B.n175 585
R199 B.n292 B.n291 585
R200 B.n293 B.n174 585
R201 B.n295 B.n294 585
R202 B.n296 B.n173 585
R203 B.n298 B.n297 585
R204 B.n299 B.n172 585
R205 B.n301 B.n300 585
R206 B.n302 B.n171 585
R207 B.n304 B.n303 585
R208 B.n305 B.n170 585
R209 B.n307 B.n306 585
R210 B.n308 B.n169 585
R211 B.n310 B.n309 585
R212 B.n311 B.n168 585
R213 B.n313 B.n312 585
R214 B.n314 B.n167 585
R215 B.n316 B.n315 585
R216 B.n317 B.n166 585
R217 B.n319 B.n318 585
R218 B.n320 B.n165 585
R219 B.n322 B.n321 585
R220 B.n323 B.n164 585
R221 B.n325 B.n324 585
R222 B.n326 B.n163 585
R223 B.n328 B.n327 585
R224 B.n329 B.n162 585
R225 B.n331 B.n330 585
R226 B.n332 B.n161 585
R227 B.n334 B.n333 585
R228 B.n335 B.n160 585
R229 B.n337 B.n336 585
R230 B.n338 B.n159 585
R231 B.n340 B.n339 585
R232 B.n342 B.n341 585
R233 B.n343 B.n155 585
R234 B.n345 B.n344 585
R235 B.n346 B.n154 585
R236 B.n348 B.n347 585
R237 B.n349 B.n153 585
R238 B.n351 B.n350 585
R239 B.n352 B.n152 585
R240 B.n354 B.n353 585
R241 B.n356 B.n149 585
R242 B.n358 B.n357 585
R243 B.n359 B.n148 585
R244 B.n361 B.n360 585
R245 B.n362 B.n147 585
R246 B.n364 B.n363 585
R247 B.n365 B.n146 585
R248 B.n367 B.n366 585
R249 B.n368 B.n145 585
R250 B.n370 B.n369 585
R251 B.n371 B.n144 585
R252 B.n373 B.n372 585
R253 B.n374 B.n143 585
R254 B.n376 B.n375 585
R255 B.n377 B.n142 585
R256 B.n379 B.n378 585
R257 B.n380 B.n141 585
R258 B.n382 B.n381 585
R259 B.n383 B.n140 585
R260 B.n385 B.n384 585
R261 B.n386 B.n139 585
R262 B.n388 B.n387 585
R263 B.n389 B.n138 585
R264 B.n391 B.n390 585
R265 B.n392 B.n137 585
R266 B.n394 B.n393 585
R267 B.n395 B.n136 585
R268 B.n397 B.n396 585
R269 B.n398 B.n135 585
R270 B.n400 B.n399 585
R271 B.n401 B.n134 585
R272 B.n403 B.n402 585
R273 B.n404 B.n133 585
R274 B.n406 B.n405 585
R275 B.n407 B.n132 585
R276 B.n409 B.n408 585
R277 B.n410 B.n131 585
R278 B.n412 B.n411 585
R279 B.n283 B.n282 585
R280 B.n281 B.n178 585
R281 B.n280 B.n279 585
R282 B.n278 B.n179 585
R283 B.n277 B.n276 585
R284 B.n275 B.n180 585
R285 B.n274 B.n273 585
R286 B.n272 B.n181 585
R287 B.n271 B.n270 585
R288 B.n269 B.n182 585
R289 B.n268 B.n267 585
R290 B.n266 B.n183 585
R291 B.n265 B.n264 585
R292 B.n263 B.n184 585
R293 B.n262 B.n261 585
R294 B.n260 B.n185 585
R295 B.n259 B.n258 585
R296 B.n257 B.n186 585
R297 B.n256 B.n255 585
R298 B.n254 B.n187 585
R299 B.n253 B.n252 585
R300 B.n251 B.n188 585
R301 B.n250 B.n249 585
R302 B.n248 B.n189 585
R303 B.n247 B.n246 585
R304 B.n245 B.n190 585
R305 B.n244 B.n243 585
R306 B.n242 B.n191 585
R307 B.n241 B.n240 585
R308 B.n239 B.n192 585
R309 B.n238 B.n237 585
R310 B.n236 B.n193 585
R311 B.n235 B.n234 585
R312 B.n233 B.n194 585
R313 B.n232 B.n231 585
R314 B.n230 B.n195 585
R315 B.n229 B.n228 585
R316 B.n227 B.n196 585
R317 B.n226 B.n225 585
R318 B.n224 B.n197 585
R319 B.n223 B.n222 585
R320 B.n221 B.n198 585
R321 B.n220 B.n219 585
R322 B.n218 B.n199 585
R323 B.n217 B.n216 585
R324 B.n215 B.n200 585
R325 B.n214 B.n213 585
R326 B.n212 B.n201 585
R327 B.n211 B.n210 585
R328 B.n209 B.n202 585
R329 B.n208 B.n207 585
R330 B.n206 B.n203 585
R331 B.n205 B.n204 585
R332 B.n2 B.n0 585
R333 B.n785 B.n1 585
R334 B.n784 B.n783 585
R335 B.n782 B.n3 585
R336 B.n781 B.n780 585
R337 B.n779 B.n4 585
R338 B.n778 B.n777 585
R339 B.n776 B.n5 585
R340 B.n775 B.n774 585
R341 B.n773 B.n6 585
R342 B.n772 B.n771 585
R343 B.n770 B.n7 585
R344 B.n769 B.n768 585
R345 B.n767 B.n8 585
R346 B.n766 B.n765 585
R347 B.n764 B.n9 585
R348 B.n763 B.n762 585
R349 B.n761 B.n10 585
R350 B.n760 B.n759 585
R351 B.n758 B.n11 585
R352 B.n757 B.n756 585
R353 B.n755 B.n12 585
R354 B.n754 B.n753 585
R355 B.n752 B.n13 585
R356 B.n751 B.n750 585
R357 B.n749 B.n14 585
R358 B.n748 B.n747 585
R359 B.n746 B.n15 585
R360 B.n745 B.n744 585
R361 B.n743 B.n16 585
R362 B.n742 B.n741 585
R363 B.n740 B.n17 585
R364 B.n739 B.n738 585
R365 B.n737 B.n18 585
R366 B.n736 B.n735 585
R367 B.n734 B.n19 585
R368 B.n733 B.n732 585
R369 B.n731 B.n20 585
R370 B.n730 B.n729 585
R371 B.n728 B.n21 585
R372 B.n727 B.n726 585
R373 B.n725 B.n22 585
R374 B.n724 B.n723 585
R375 B.n722 B.n23 585
R376 B.n721 B.n720 585
R377 B.n719 B.n24 585
R378 B.n718 B.n717 585
R379 B.n716 B.n25 585
R380 B.n715 B.n714 585
R381 B.n713 B.n26 585
R382 B.n712 B.n711 585
R383 B.n710 B.n27 585
R384 B.n709 B.n708 585
R385 B.n707 B.n28 585
R386 B.n706 B.n705 585
R387 B.n787 B.n786 585
R388 B.n282 B.n177 492.5
R389 B.n706 B.n29 492.5
R390 B.n413 B.n412 492.5
R391 B.n576 B.n575 492.5
R392 B.n150 B.t11 427.065
R393 B.n56 B.t4 427.065
R394 B.n156 B.t8 427.065
R395 B.n48 B.t1 427.065
R396 B.n151 B.t10 351.428
R397 B.n57 B.t5 351.428
R398 B.n157 B.t7 351.428
R399 B.n49 B.t2 351.428
R400 B.n150 B.t9 281.118
R401 B.n156 B.t6 281.118
R402 B.n48 B.t0 281.118
R403 B.n56 B.t3 281.118
R404 B.n282 B.n281 163.367
R405 B.n281 B.n280 163.367
R406 B.n280 B.n179 163.367
R407 B.n276 B.n179 163.367
R408 B.n276 B.n275 163.367
R409 B.n275 B.n274 163.367
R410 B.n274 B.n181 163.367
R411 B.n270 B.n181 163.367
R412 B.n270 B.n269 163.367
R413 B.n269 B.n268 163.367
R414 B.n268 B.n183 163.367
R415 B.n264 B.n183 163.367
R416 B.n264 B.n263 163.367
R417 B.n263 B.n262 163.367
R418 B.n262 B.n185 163.367
R419 B.n258 B.n185 163.367
R420 B.n258 B.n257 163.367
R421 B.n257 B.n256 163.367
R422 B.n256 B.n187 163.367
R423 B.n252 B.n187 163.367
R424 B.n252 B.n251 163.367
R425 B.n251 B.n250 163.367
R426 B.n250 B.n189 163.367
R427 B.n246 B.n189 163.367
R428 B.n246 B.n245 163.367
R429 B.n245 B.n244 163.367
R430 B.n244 B.n191 163.367
R431 B.n240 B.n191 163.367
R432 B.n240 B.n239 163.367
R433 B.n239 B.n238 163.367
R434 B.n238 B.n193 163.367
R435 B.n234 B.n193 163.367
R436 B.n234 B.n233 163.367
R437 B.n233 B.n232 163.367
R438 B.n232 B.n195 163.367
R439 B.n228 B.n195 163.367
R440 B.n228 B.n227 163.367
R441 B.n227 B.n226 163.367
R442 B.n226 B.n197 163.367
R443 B.n222 B.n197 163.367
R444 B.n222 B.n221 163.367
R445 B.n221 B.n220 163.367
R446 B.n220 B.n199 163.367
R447 B.n216 B.n199 163.367
R448 B.n216 B.n215 163.367
R449 B.n215 B.n214 163.367
R450 B.n214 B.n201 163.367
R451 B.n210 B.n201 163.367
R452 B.n210 B.n209 163.367
R453 B.n209 B.n208 163.367
R454 B.n208 B.n203 163.367
R455 B.n204 B.n203 163.367
R456 B.n204 B.n2 163.367
R457 B.n786 B.n2 163.367
R458 B.n786 B.n785 163.367
R459 B.n785 B.n784 163.367
R460 B.n784 B.n3 163.367
R461 B.n780 B.n3 163.367
R462 B.n780 B.n779 163.367
R463 B.n779 B.n778 163.367
R464 B.n778 B.n5 163.367
R465 B.n774 B.n5 163.367
R466 B.n774 B.n773 163.367
R467 B.n773 B.n772 163.367
R468 B.n772 B.n7 163.367
R469 B.n768 B.n7 163.367
R470 B.n768 B.n767 163.367
R471 B.n767 B.n766 163.367
R472 B.n766 B.n9 163.367
R473 B.n762 B.n9 163.367
R474 B.n762 B.n761 163.367
R475 B.n761 B.n760 163.367
R476 B.n760 B.n11 163.367
R477 B.n756 B.n11 163.367
R478 B.n756 B.n755 163.367
R479 B.n755 B.n754 163.367
R480 B.n754 B.n13 163.367
R481 B.n750 B.n13 163.367
R482 B.n750 B.n749 163.367
R483 B.n749 B.n748 163.367
R484 B.n748 B.n15 163.367
R485 B.n744 B.n15 163.367
R486 B.n744 B.n743 163.367
R487 B.n743 B.n742 163.367
R488 B.n742 B.n17 163.367
R489 B.n738 B.n17 163.367
R490 B.n738 B.n737 163.367
R491 B.n737 B.n736 163.367
R492 B.n736 B.n19 163.367
R493 B.n732 B.n19 163.367
R494 B.n732 B.n731 163.367
R495 B.n731 B.n730 163.367
R496 B.n730 B.n21 163.367
R497 B.n726 B.n21 163.367
R498 B.n726 B.n725 163.367
R499 B.n725 B.n724 163.367
R500 B.n724 B.n23 163.367
R501 B.n720 B.n23 163.367
R502 B.n720 B.n719 163.367
R503 B.n719 B.n718 163.367
R504 B.n718 B.n25 163.367
R505 B.n714 B.n25 163.367
R506 B.n714 B.n713 163.367
R507 B.n713 B.n712 163.367
R508 B.n712 B.n27 163.367
R509 B.n708 B.n27 163.367
R510 B.n708 B.n707 163.367
R511 B.n707 B.n706 163.367
R512 B.n286 B.n177 163.367
R513 B.n287 B.n286 163.367
R514 B.n288 B.n287 163.367
R515 B.n288 B.n175 163.367
R516 B.n292 B.n175 163.367
R517 B.n293 B.n292 163.367
R518 B.n294 B.n293 163.367
R519 B.n294 B.n173 163.367
R520 B.n298 B.n173 163.367
R521 B.n299 B.n298 163.367
R522 B.n300 B.n299 163.367
R523 B.n300 B.n171 163.367
R524 B.n304 B.n171 163.367
R525 B.n305 B.n304 163.367
R526 B.n306 B.n305 163.367
R527 B.n306 B.n169 163.367
R528 B.n310 B.n169 163.367
R529 B.n311 B.n310 163.367
R530 B.n312 B.n311 163.367
R531 B.n312 B.n167 163.367
R532 B.n316 B.n167 163.367
R533 B.n317 B.n316 163.367
R534 B.n318 B.n317 163.367
R535 B.n318 B.n165 163.367
R536 B.n322 B.n165 163.367
R537 B.n323 B.n322 163.367
R538 B.n324 B.n323 163.367
R539 B.n324 B.n163 163.367
R540 B.n328 B.n163 163.367
R541 B.n329 B.n328 163.367
R542 B.n330 B.n329 163.367
R543 B.n330 B.n161 163.367
R544 B.n334 B.n161 163.367
R545 B.n335 B.n334 163.367
R546 B.n336 B.n335 163.367
R547 B.n336 B.n159 163.367
R548 B.n340 B.n159 163.367
R549 B.n341 B.n340 163.367
R550 B.n341 B.n155 163.367
R551 B.n345 B.n155 163.367
R552 B.n346 B.n345 163.367
R553 B.n347 B.n346 163.367
R554 B.n347 B.n153 163.367
R555 B.n351 B.n153 163.367
R556 B.n352 B.n351 163.367
R557 B.n353 B.n352 163.367
R558 B.n353 B.n149 163.367
R559 B.n358 B.n149 163.367
R560 B.n359 B.n358 163.367
R561 B.n360 B.n359 163.367
R562 B.n360 B.n147 163.367
R563 B.n364 B.n147 163.367
R564 B.n365 B.n364 163.367
R565 B.n366 B.n365 163.367
R566 B.n366 B.n145 163.367
R567 B.n370 B.n145 163.367
R568 B.n371 B.n370 163.367
R569 B.n372 B.n371 163.367
R570 B.n372 B.n143 163.367
R571 B.n376 B.n143 163.367
R572 B.n377 B.n376 163.367
R573 B.n378 B.n377 163.367
R574 B.n378 B.n141 163.367
R575 B.n382 B.n141 163.367
R576 B.n383 B.n382 163.367
R577 B.n384 B.n383 163.367
R578 B.n384 B.n139 163.367
R579 B.n388 B.n139 163.367
R580 B.n389 B.n388 163.367
R581 B.n390 B.n389 163.367
R582 B.n390 B.n137 163.367
R583 B.n394 B.n137 163.367
R584 B.n395 B.n394 163.367
R585 B.n396 B.n395 163.367
R586 B.n396 B.n135 163.367
R587 B.n400 B.n135 163.367
R588 B.n401 B.n400 163.367
R589 B.n402 B.n401 163.367
R590 B.n402 B.n133 163.367
R591 B.n406 B.n133 163.367
R592 B.n407 B.n406 163.367
R593 B.n408 B.n407 163.367
R594 B.n408 B.n131 163.367
R595 B.n412 B.n131 163.367
R596 B.n414 B.n413 163.367
R597 B.n414 B.n129 163.367
R598 B.n418 B.n129 163.367
R599 B.n419 B.n418 163.367
R600 B.n420 B.n419 163.367
R601 B.n420 B.n127 163.367
R602 B.n424 B.n127 163.367
R603 B.n425 B.n424 163.367
R604 B.n426 B.n425 163.367
R605 B.n426 B.n125 163.367
R606 B.n430 B.n125 163.367
R607 B.n431 B.n430 163.367
R608 B.n432 B.n431 163.367
R609 B.n432 B.n123 163.367
R610 B.n436 B.n123 163.367
R611 B.n437 B.n436 163.367
R612 B.n438 B.n437 163.367
R613 B.n438 B.n121 163.367
R614 B.n442 B.n121 163.367
R615 B.n443 B.n442 163.367
R616 B.n444 B.n443 163.367
R617 B.n444 B.n119 163.367
R618 B.n448 B.n119 163.367
R619 B.n449 B.n448 163.367
R620 B.n450 B.n449 163.367
R621 B.n450 B.n117 163.367
R622 B.n454 B.n117 163.367
R623 B.n455 B.n454 163.367
R624 B.n456 B.n455 163.367
R625 B.n456 B.n115 163.367
R626 B.n460 B.n115 163.367
R627 B.n461 B.n460 163.367
R628 B.n462 B.n461 163.367
R629 B.n462 B.n113 163.367
R630 B.n466 B.n113 163.367
R631 B.n467 B.n466 163.367
R632 B.n468 B.n467 163.367
R633 B.n468 B.n111 163.367
R634 B.n472 B.n111 163.367
R635 B.n473 B.n472 163.367
R636 B.n474 B.n473 163.367
R637 B.n474 B.n109 163.367
R638 B.n478 B.n109 163.367
R639 B.n479 B.n478 163.367
R640 B.n480 B.n479 163.367
R641 B.n480 B.n107 163.367
R642 B.n484 B.n107 163.367
R643 B.n485 B.n484 163.367
R644 B.n486 B.n485 163.367
R645 B.n486 B.n105 163.367
R646 B.n490 B.n105 163.367
R647 B.n491 B.n490 163.367
R648 B.n492 B.n491 163.367
R649 B.n492 B.n103 163.367
R650 B.n496 B.n103 163.367
R651 B.n497 B.n496 163.367
R652 B.n498 B.n497 163.367
R653 B.n498 B.n101 163.367
R654 B.n502 B.n101 163.367
R655 B.n503 B.n502 163.367
R656 B.n504 B.n503 163.367
R657 B.n504 B.n99 163.367
R658 B.n508 B.n99 163.367
R659 B.n509 B.n508 163.367
R660 B.n510 B.n509 163.367
R661 B.n510 B.n97 163.367
R662 B.n514 B.n97 163.367
R663 B.n515 B.n514 163.367
R664 B.n516 B.n515 163.367
R665 B.n516 B.n95 163.367
R666 B.n520 B.n95 163.367
R667 B.n521 B.n520 163.367
R668 B.n522 B.n521 163.367
R669 B.n522 B.n93 163.367
R670 B.n526 B.n93 163.367
R671 B.n527 B.n526 163.367
R672 B.n528 B.n527 163.367
R673 B.n528 B.n91 163.367
R674 B.n532 B.n91 163.367
R675 B.n533 B.n532 163.367
R676 B.n534 B.n533 163.367
R677 B.n534 B.n89 163.367
R678 B.n538 B.n89 163.367
R679 B.n539 B.n538 163.367
R680 B.n540 B.n539 163.367
R681 B.n540 B.n87 163.367
R682 B.n544 B.n87 163.367
R683 B.n545 B.n544 163.367
R684 B.n546 B.n545 163.367
R685 B.n546 B.n85 163.367
R686 B.n550 B.n85 163.367
R687 B.n551 B.n550 163.367
R688 B.n552 B.n551 163.367
R689 B.n552 B.n83 163.367
R690 B.n556 B.n83 163.367
R691 B.n557 B.n556 163.367
R692 B.n558 B.n557 163.367
R693 B.n558 B.n81 163.367
R694 B.n562 B.n81 163.367
R695 B.n563 B.n562 163.367
R696 B.n564 B.n563 163.367
R697 B.n564 B.n79 163.367
R698 B.n568 B.n79 163.367
R699 B.n569 B.n568 163.367
R700 B.n570 B.n569 163.367
R701 B.n570 B.n77 163.367
R702 B.n574 B.n77 163.367
R703 B.n575 B.n574 163.367
R704 B.n702 B.n29 163.367
R705 B.n702 B.n701 163.367
R706 B.n701 B.n700 163.367
R707 B.n700 B.n31 163.367
R708 B.n696 B.n31 163.367
R709 B.n696 B.n695 163.367
R710 B.n695 B.n694 163.367
R711 B.n694 B.n33 163.367
R712 B.n690 B.n33 163.367
R713 B.n690 B.n689 163.367
R714 B.n689 B.n688 163.367
R715 B.n688 B.n35 163.367
R716 B.n684 B.n35 163.367
R717 B.n684 B.n683 163.367
R718 B.n683 B.n682 163.367
R719 B.n682 B.n37 163.367
R720 B.n678 B.n37 163.367
R721 B.n678 B.n677 163.367
R722 B.n677 B.n676 163.367
R723 B.n676 B.n39 163.367
R724 B.n672 B.n39 163.367
R725 B.n672 B.n671 163.367
R726 B.n671 B.n670 163.367
R727 B.n670 B.n41 163.367
R728 B.n666 B.n41 163.367
R729 B.n666 B.n665 163.367
R730 B.n665 B.n664 163.367
R731 B.n664 B.n43 163.367
R732 B.n660 B.n43 163.367
R733 B.n660 B.n659 163.367
R734 B.n659 B.n658 163.367
R735 B.n658 B.n45 163.367
R736 B.n654 B.n45 163.367
R737 B.n654 B.n653 163.367
R738 B.n653 B.n652 163.367
R739 B.n652 B.n47 163.367
R740 B.n648 B.n47 163.367
R741 B.n648 B.n647 163.367
R742 B.n647 B.n51 163.367
R743 B.n643 B.n51 163.367
R744 B.n643 B.n642 163.367
R745 B.n642 B.n641 163.367
R746 B.n641 B.n53 163.367
R747 B.n637 B.n53 163.367
R748 B.n637 B.n636 163.367
R749 B.n636 B.n635 163.367
R750 B.n635 B.n55 163.367
R751 B.n630 B.n55 163.367
R752 B.n630 B.n629 163.367
R753 B.n629 B.n628 163.367
R754 B.n628 B.n59 163.367
R755 B.n624 B.n59 163.367
R756 B.n624 B.n623 163.367
R757 B.n623 B.n622 163.367
R758 B.n622 B.n61 163.367
R759 B.n618 B.n61 163.367
R760 B.n618 B.n617 163.367
R761 B.n617 B.n616 163.367
R762 B.n616 B.n63 163.367
R763 B.n612 B.n63 163.367
R764 B.n612 B.n611 163.367
R765 B.n611 B.n610 163.367
R766 B.n610 B.n65 163.367
R767 B.n606 B.n65 163.367
R768 B.n606 B.n605 163.367
R769 B.n605 B.n604 163.367
R770 B.n604 B.n67 163.367
R771 B.n600 B.n67 163.367
R772 B.n600 B.n599 163.367
R773 B.n599 B.n598 163.367
R774 B.n598 B.n69 163.367
R775 B.n594 B.n69 163.367
R776 B.n594 B.n593 163.367
R777 B.n593 B.n592 163.367
R778 B.n592 B.n71 163.367
R779 B.n588 B.n71 163.367
R780 B.n588 B.n587 163.367
R781 B.n587 B.n586 163.367
R782 B.n586 B.n73 163.367
R783 B.n582 B.n73 163.367
R784 B.n582 B.n581 163.367
R785 B.n581 B.n580 163.367
R786 B.n580 B.n75 163.367
R787 B.n576 B.n75 163.367
R788 B.n151 B.n150 75.6369
R789 B.n157 B.n156 75.6369
R790 B.n49 B.n48 75.6369
R791 B.n57 B.n56 75.6369
R792 B.n355 B.n151 59.5399
R793 B.n158 B.n157 59.5399
R794 B.n50 B.n49 59.5399
R795 B.n633 B.n57 59.5399
R796 B.n705 B.n704 32.0005
R797 B.n577 B.n76 32.0005
R798 B.n411 B.n130 32.0005
R799 B.n284 B.n283 32.0005
R800 B B.n787 18.0485
R801 B.n704 B.n703 10.6151
R802 B.n703 B.n30 10.6151
R803 B.n699 B.n30 10.6151
R804 B.n699 B.n698 10.6151
R805 B.n698 B.n697 10.6151
R806 B.n697 B.n32 10.6151
R807 B.n693 B.n32 10.6151
R808 B.n693 B.n692 10.6151
R809 B.n692 B.n691 10.6151
R810 B.n691 B.n34 10.6151
R811 B.n687 B.n34 10.6151
R812 B.n687 B.n686 10.6151
R813 B.n686 B.n685 10.6151
R814 B.n685 B.n36 10.6151
R815 B.n681 B.n36 10.6151
R816 B.n681 B.n680 10.6151
R817 B.n680 B.n679 10.6151
R818 B.n679 B.n38 10.6151
R819 B.n675 B.n38 10.6151
R820 B.n675 B.n674 10.6151
R821 B.n674 B.n673 10.6151
R822 B.n673 B.n40 10.6151
R823 B.n669 B.n40 10.6151
R824 B.n669 B.n668 10.6151
R825 B.n668 B.n667 10.6151
R826 B.n667 B.n42 10.6151
R827 B.n663 B.n42 10.6151
R828 B.n663 B.n662 10.6151
R829 B.n662 B.n661 10.6151
R830 B.n661 B.n44 10.6151
R831 B.n657 B.n44 10.6151
R832 B.n657 B.n656 10.6151
R833 B.n656 B.n655 10.6151
R834 B.n655 B.n46 10.6151
R835 B.n651 B.n46 10.6151
R836 B.n651 B.n650 10.6151
R837 B.n650 B.n649 10.6151
R838 B.n646 B.n645 10.6151
R839 B.n645 B.n644 10.6151
R840 B.n644 B.n52 10.6151
R841 B.n640 B.n52 10.6151
R842 B.n640 B.n639 10.6151
R843 B.n639 B.n638 10.6151
R844 B.n638 B.n54 10.6151
R845 B.n634 B.n54 10.6151
R846 B.n632 B.n631 10.6151
R847 B.n631 B.n58 10.6151
R848 B.n627 B.n58 10.6151
R849 B.n627 B.n626 10.6151
R850 B.n626 B.n625 10.6151
R851 B.n625 B.n60 10.6151
R852 B.n621 B.n60 10.6151
R853 B.n621 B.n620 10.6151
R854 B.n620 B.n619 10.6151
R855 B.n619 B.n62 10.6151
R856 B.n615 B.n62 10.6151
R857 B.n615 B.n614 10.6151
R858 B.n614 B.n613 10.6151
R859 B.n613 B.n64 10.6151
R860 B.n609 B.n64 10.6151
R861 B.n609 B.n608 10.6151
R862 B.n608 B.n607 10.6151
R863 B.n607 B.n66 10.6151
R864 B.n603 B.n66 10.6151
R865 B.n603 B.n602 10.6151
R866 B.n602 B.n601 10.6151
R867 B.n601 B.n68 10.6151
R868 B.n597 B.n68 10.6151
R869 B.n597 B.n596 10.6151
R870 B.n596 B.n595 10.6151
R871 B.n595 B.n70 10.6151
R872 B.n591 B.n70 10.6151
R873 B.n591 B.n590 10.6151
R874 B.n590 B.n589 10.6151
R875 B.n589 B.n72 10.6151
R876 B.n585 B.n72 10.6151
R877 B.n585 B.n584 10.6151
R878 B.n584 B.n583 10.6151
R879 B.n583 B.n74 10.6151
R880 B.n579 B.n74 10.6151
R881 B.n579 B.n578 10.6151
R882 B.n578 B.n577 10.6151
R883 B.n415 B.n130 10.6151
R884 B.n416 B.n415 10.6151
R885 B.n417 B.n416 10.6151
R886 B.n417 B.n128 10.6151
R887 B.n421 B.n128 10.6151
R888 B.n422 B.n421 10.6151
R889 B.n423 B.n422 10.6151
R890 B.n423 B.n126 10.6151
R891 B.n427 B.n126 10.6151
R892 B.n428 B.n427 10.6151
R893 B.n429 B.n428 10.6151
R894 B.n429 B.n124 10.6151
R895 B.n433 B.n124 10.6151
R896 B.n434 B.n433 10.6151
R897 B.n435 B.n434 10.6151
R898 B.n435 B.n122 10.6151
R899 B.n439 B.n122 10.6151
R900 B.n440 B.n439 10.6151
R901 B.n441 B.n440 10.6151
R902 B.n441 B.n120 10.6151
R903 B.n445 B.n120 10.6151
R904 B.n446 B.n445 10.6151
R905 B.n447 B.n446 10.6151
R906 B.n447 B.n118 10.6151
R907 B.n451 B.n118 10.6151
R908 B.n452 B.n451 10.6151
R909 B.n453 B.n452 10.6151
R910 B.n453 B.n116 10.6151
R911 B.n457 B.n116 10.6151
R912 B.n458 B.n457 10.6151
R913 B.n459 B.n458 10.6151
R914 B.n459 B.n114 10.6151
R915 B.n463 B.n114 10.6151
R916 B.n464 B.n463 10.6151
R917 B.n465 B.n464 10.6151
R918 B.n465 B.n112 10.6151
R919 B.n469 B.n112 10.6151
R920 B.n470 B.n469 10.6151
R921 B.n471 B.n470 10.6151
R922 B.n471 B.n110 10.6151
R923 B.n475 B.n110 10.6151
R924 B.n476 B.n475 10.6151
R925 B.n477 B.n476 10.6151
R926 B.n477 B.n108 10.6151
R927 B.n481 B.n108 10.6151
R928 B.n482 B.n481 10.6151
R929 B.n483 B.n482 10.6151
R930 B.n483 B.n106 10.6151
R931 B.n487 B.n106 10.6151
R932 B.n488 B.n487 10.6151
R933 B.n489 B.n488 10.6151
R934 B.n489 B.n104 10.6151
R935 B.n493 B.n104 10.6151
R936 B.n494 B.n493 10.6151
R937 B.n495 B.n494 10.6151
R938 B.n495 B.n102 10.6151
R939 B.n499 B.n102 10.6151
R940 B.n500 B.n499 10.6151
R941 B.n501 B.n500 10.6151
R942 B.n501 B.n100 10.6151
R943 B.n505 B.n100 10.6151
R944 B.n506 B.n505 10.6151
R945 B.n507 B.n506 10.6151
R946 B.n507 B.n98 10.6151
R947 B.n511 B.n98 10.6151
R948 B.n512 B.n511 10.6151
R949 B.n513 B.n512 10.6151
R950 B.n513 B.n96 10.6151
R951 B.n517 B.n96 10.6151
R952 B.n518 B.n517 10.6151
R953 B.n519 B.n518 10.6151
R954 B.n519 B.n94 10.6151
R955 B.n523 B.n94 10.6151
R956 B.n524 B.n523 10.6151
R957 B.n525 B.n524 10.6151
R958 B.n525 B.n92 10.6151
R959 B.n529 B.n92 10.6151
R960 B.n530 B.n529 10.6151
R961 B.n531 B.n530 10.6151
R962 B.n531 B.n90 10.6151
R963 B.n535 B.n90 10.6151
R964 B.n536 B.n535 10.6151
R965 B.n537 B.n536 10.6151
R966 B.n537 B.n88 10.6151
R967 B.n541 B.n88 10.6151
R968 B.n542 B.n541 10.6151
R969 B.n543 B.n542 10.6151
R970 B.n543 B.n86 10.6151
R971 B.n547 B.n86 10.6151
R972 B.n548 B.n547 10.6151
R973 B.n549 B.n548 10.6151
R974 B.n549 B.n84 10.6151
R975 B.n553 B.n84 10.6151
R976 B.n554 B.n553 10.6151
R977 B.n555 B.n554 10.6151
R978 B.n555 B.n82 10.6151
R979 B.n559 B.n82 10.6151
R980 B.n560 B.n559 10.6151
R981 B.n561 B.n560 10.6151
R982 B.n561 B.n80 10.6151
R983 B.n565 B.n80 10.6151
R984 B.n566 B.n565 10.6151
R985 B.n567 B.n566 10.6151
R986 B.n567 B.n78 10.6151
R987 B.n571 B.n78 10.6151
R988 B.n572 B.n571 10.6151
R989 B.n573 B.n572 10.6151
R990 B.n573 B.n76 10.6151
R991 B.n285 B.n284 10.6151
R992 B.n285 B.n176 10.6151
R993 B.n289 B.n176 10.6151
R994 B.n290 B.n289 10.6151
R995 B.n291 B.n290 10.6151
R996 B.n291 B.n174 10.6151
R997 B.n295 B.n174 10.6151
R998 B.n296 B.n295 10.6151
R999 B.n297 B.n296 10.6151
R1000 B.n297 B.n172 10.6151
R1001 B.n301 B.n172 10.6151
R1002 B.n302 B.n301 10.6151
R1003 B.n303 B.n302 10.6151
R1004 B.n303 B.n170 10.6151
R1005 B.n307 B.n170 10.6151
R1006 B.n308 B.n307 10.6151
R1007 B.n309 B.n308 10.6151
R1008 B.n309 B.n168 10.6151
R1009 B.n313 B.n168 10.6151
R1010 B.n314 B.n313 10.6151
R1011 B.n315 B.n314 10.6151
R1012 B.n315 B.n166 10.6151
R1013 B.n319 B.n166 10.6151
R1014 B.n320 B.n319 10.6151
R1015 B.n321 B.n320 10.6151
R1016 B.n321 B.n164 10.6151
R1017 B.n325 B.n164 10.6151
R1018 B.n326 B.n325 10.6151
R1019 B.n327 B.n326 10.6151
R1020 B.n327 B.n162 10.6151
R1021 B.n331 B.n162 10.6151
R1022 B.n332 B.n331 10.6151
R1023 B.n333 B.n332 10.6151
R1024 B.n333 B.n160 10.6151
R1025 B.n337 B.n160 10.6151
R1026 B.n338 B.n337 10.6151
R1027 B.n339 B.n338 10.6151
R1028 B.n343 B.n342 10.6151
R1029 B.n344 B.n343 10.6151
R1030 B.n344 B.n154 10.6151
R1031 B.n348 B.n154 10.6151
R1032 B.n349 B.n348 10.6151
R1033 B.n350 B.n349 10.6151
R1034 B.n350 B.n152 10.6151
R1035 B.n354 B.n152 10.6151
R1036 B.n357 B.n356 10.6151
R1037 B.n357 B.n148 10.6151
R1038 B.n361 B.n148 10.6151
R1039 B.n362 B.n361 10.6151
R1040 B.n363 B.n362 10.6151
R1041 B.n363 B.n146 10.6151
R1042 B.n367 B.n146 10.6151
R1043 B.n368 B.n367 10.6151
R1044 B.n369 B.n368 10.6151
R1045 B.n369 B.n144 10.6151
R1046 B.n373 B.n144 10.6151
R1047 B.n374 B.n373 10.6151
R1048 B.n375 B.n374 10.6151
R1049 B.n375 B.n142 10.6151
R1050 B.n379 B.n142 10.6151
R1051 B.n380 B.n379 10.6151
R1052 B.n381 B.n380 10.6151
R1053 B.n381 B.n140 10.6151
R1054 B.n385 B.n140 10.6151
R1055 B.n386 B.n385 10.6151
R1056 B.n387 B.n386 10.6151
R1057 B.n387 B.n138 10.6151
R1058 B.n391 B.n138 10.6151
R1059 B.n392 B.n391 10.6151
R1060 B.n393 B.n392 10.6151
R1061 B.n393 B.n136 10.6151
R1062 B.n397 B.n136 10.6151
R1063 B.n398 B.n397 10.6151
R1064 B.n399 B.n398 10.6151
R1065 B.n399 B.n134 10.6151
R1066 B.n403 B.n134 10.6151
R1067 B.n404 B.n403 10.6151
R1068 B.n405 B.n404 10.6151
R1069 B.n405 B.n132 10.6151
R1070 B.n409 B.n132 10.6151
R1071 B.n410 B.n409 10.6151
R1072 B.n411 B.n410 10.6151
R1073 B.n283 B.n178 10.6151
R1074 B.n279 B.n178 10.6151
R1075 B.n279 B.n278 10.6151
R1076 B.n278 B.n277 10.6151
R1077 B.n277 B.n180 10.6151
R1078 B.n273 B.n180 10.6151
R1079 B.n273 B.n272 10.6151
R1080 B.n272 B.n271 10.6151
R1081 B.n271 B.n182 10.6151
R1082 B.n267 B.n182 10.6151
R1083 B.n267 B.n266 10.6151
R1084 B.n266 B.n265 10.6151
R1085 B.n265 B.n184 10.6151
R1086 B.n261 B.n184 10.6151
R1087 B.n261 B.n260 10.6151
R1088 B.n260 B.n259 10.6151
R1089 B.n259 B.n186 10.6151
R1090 B.n255 B.n186 10.6151
R1091 B.n255 B.n254 10.6151
R1092 B.n254 B.n253 10.6151
R1093 B.n253 B.n188 10.6151
R1094 B.n249 B.n188 10.6151
R1095 B.n249 B.n248 10.6151
R1096 B.n248 B.n247 10.6151
R1097 B.n247 B.n190 10.6151
R1098 B.n243 B.n190 10.6151
R1099 B.n243 B.n242 10.6151
R1100 B.n242 B.n241 10.6151
R1101 B.n241 B.n192 10.6151
R1102 B.n237 B.n192 10.6151
R1103 B.n237 B.n236 10.6151
R1104 B.n236 B.n235 10.6151
R1105 B.n235 B.n194 10.6151
R1106 B.n231 B.n194 10.6151
R1107 B.n231 B.n230 10.6151
R1108 B.n230 B.n229 10.6151
R1109 B.n229 B.n196 10.6151
R1110 B.n225 B.n196 10.6151
R1111 B.n225 B.n224 10.6151
R1112 B.n224 B.n223 10.6151
R1113 B.n223 B.n198 10.6151
R1114 B.n219 B.n198 10.6151
R1115 B.n219 B.n218 10.6151
R1116 B.n218 B.n217 10.6151
R1117 B.n217 B.n200 10.6151
R1118 B.n213 B.n200 10.6151
R1119 B.n213 B.n212 10.6151
R1120 B.n212 B.n211 10.6151
R1121 B.n211 B.n202 10.6151
R1122 B.n207 B.n202 10.6151
R1123 B.n207 B.n206 10.6151
R1124 B.n206 B.n205 10.6151
R1125 B.n205 B.n0 10.6151
R1126 B.n783 B.n1 10.6151
R1127 B.n783 B.n782 10.6151
R1128 B.n782 B.n781 10.6151
R1129 B.n781 B.n4 10.6151
R1130 B.n777 B.n4 10.6151
R1131 B.n777 B.n776 10.6151
R1132 B.n776 B.n775 10.6151
R1133 B.n775 B.n6 10.6151
R1134 B.n771 B.n6 10.6151
R1135 B.n771 B.n770 10.6151
R1136 B.n770 B.n769 10.6151
R1137 B.n769 B.n8 10.6151
R1138 B.n765 B.n8 10.6151
R1139 B.n765 B.n764 10.6151
R1140 B.n764 B.n763 10.6151
R1141 B.n763 B.n10 10.6151
R1142 B.n759 B.n10 10.6151
R1143 B.n759 B.n758 10.6151
R1144 B.n758 B.n757 10.6151
R1145 B.n757 B.n12 10.6151
R1146 B.n753 B.n12 10.6151
R1147 B.n753 B.n752 10.6151
R1148 B.n752 B.n751 10.6151
R1149 B.n751 B.n14 10.6151
R1150 B.n747 B.n14 10.6151
R1151 B.n747 B.n746 10.6151
R1152 B.n746 B.n745 10.6151
R1153 B.n745 B.n16 10.6151
R1154 B.n741 B.n16 10.6151
R1155 B.n741 B.n740 10.6151
R1156 B.n740 B.n739 10.6151
R1157 B.n739 B.n18 10.6151
R1158 B.n735 B.n18 10.6151
R1159 B.n735 B.n734 10.6151
R1160 B.n734 B.n733 10.6151
R1161 B.n733 B.n20 10.6151
R1162 B.n729 B.n20 10.6151
R1163 B.n729 B.n728 10.6151
R1164 B.n728 B.n727 10.6151
R1165 B.n727 B.n22 10.6151
R1166 B.n723 B.n22 10.6151
R1167 B.n723 B.n722 10.6151
R1168 B.n722 B.n721 10.6151
R1169 B.n721 B.n24 10.6151
R1170 B.n717 B.n24 10.6151
R1171 B.n717 B.n716 10.6151
R1172 B.n716 B.n715 10.6151
R1173 B.n715 B.n26 10.6151
R1174 B.n711 B.n26 10.6151
R1175 B.n711 B.n710 10.6151
R1176 B.n710 B.n709 10.6151
R1177 B.n709 B.n28 10.6151
R1178 B.n705 B.n28 10.6151
R1179 B.n646 B.n50 6.5566
R1180 B.n634 B.n633 6.5566
R1181 B.n342 B.n158 6.5566
R1182 B.n355 B.n354 6.5566
R1183 B.n649 B.n50 4.05904
R1184 B.n633 B.n632 4.05904
R1185 B.n339 B.n158 4.05904
R1186 B.n356 B.n355 4.05904
R1187 B.n787 B.n0 2.81026
R1188 B.n787 B.n1 2.81026
R1189 VN.n38 VN.n37 161.3
R1190 VN.n36 VN.n21 161.3
R1191 VN.n35 VN.n34 161.3
R1192 VN.n33 VN.n22 161.3
R1193 VN.n32 VN.n31 161.3
R1194 VN.n30 VN.n23 161.3
R1195 VN.n29 VN.n28 161.3
R1196 VN.n27 VN.n24 161.3
R1197 VN.n18 VN.n17 161.3
R1198 VN.n16 VN.n1 161.3
R1199 VN.n15 VN.n14 161.3
R1200 VN.n13 VN.n2 161.3
R1201 VN.n12 VN.n11 161.3
R1202 VN.n10 VN.n3 161.3
R1203 VN.n9 VN.n8 161.3
R1204 VN.n7 VN.n4 161.3
R1205 VN.n26 VN.t2 104.975
R1206 VN.n6 VN.t1 104.975
R1207 VN.n19 VN.n0 82.868
R1208 VN.n39 VN.n20 82.868
R1209 VN.n5 VN.t0 71.963
R1210 VN.n0 VN.t4 71.963
R1211 VN.n25 VN.t3 71.963
R1212 VN.n20 VN.t5 71.963
R1213 VN.n6 VN.n5 62.4546
R1214 VN.n26 VN.n25 62.4546
R1215 VN.n11 VN.n2 56.5617
R1216 VN.n31 VN.n22 56.5617
R1217 VN VN.n39 51.6951
R1218 VN.n9 VN.n4 24.5923
R1219 VN.n10 VN.n9 24.5923
R1220 VN.n11 VN.n10 24.5923
R1221 VN.n15 VN.n2 24.5923
R1222 VN.n16 VN.n15 24.5923
R1223 VN.n17 VN.n16 24.5923
R1224 VN.n31 VN.n30 24.5923
R1225 VN.n30 VN.n29 24.5923
R1226 VN.n29 VN.n24 24.5923
R1227 VN.n37 VN.n36 24.5923
R1228 VN.n36 VN.n35 24.5923
R1229 VN.n35 VN.n22 24.5923
R1230 VN.n5 VN.n4 12.2964
R1231 VN.n25 VN.n24 12.2964
R1232 VN.n17 VN.n0 7.37805
R1233 VN.n37 VN.n20 7.37805
R1234 VN.n27 VN.n26 3.23081
R1235 VN.n7 VN.n6 3.23081
R1236 VN.n39 VN.n38 0.354861
R1237 VN.n19 VN.n18 0.354861
R1238 VN VN.n19 0.267071
R1239 VN.n38 VN.n21 0.189894
R1240 VN.n34 VN.n21 0.189894
R1241 VN.n34 VN.n33 0.189894
R1242 VN.n33 VN.n32 0.189894
R1243 VN.n32 VN.n23 0.189894
R1244 VN.n28 VN.n23 0.189894
R1245 VN.n28 VN.n27 0.189894
R1246 VN.n8 VN.n7 0.189894
R1247 VN.n8 VN.n3 0.189894
R1248 VN.n12 VN.n3 0.189894
R1249 VN.n13 VN.n12 0.189894
R1250 VN.n14 VN.n13 0.189894
R1251 VN.n14 VN.n1 0.189894
R1252 VN.n18 VN.n1 0.189894
R1253 VDD2.n111 VDD2.n59 756.745
R1254 VDD2.n52 VDD2.n0 756.745
R1255 VDD2.n112 VDD2.n111 585
R1256 VDD2.n110 VDD2.n109 585
R1257 VDD2.n63 VDD2.n62 585
R1258 VDD2.n104 VDD2.n103 585
R1259 VDD2.n102 VDD2.n101 585
R1260 VDD2.n100 VDD2.n66 585
R1261 VDD2.n70 VDD2.n67 585
R1262 VDD2.n95 VDD2.n94 585
R1263 VDD2.n93 VDD2.n92 585
R1264 VDD2.n72 VDD2.n71 585
R1265 VDD2.n87 VDD2.n86 585
R1266 VDD2.n85 VDD2.n84 585
R1267 VDD2.n76 VDD2.n75 585
R1268 VDD2.n79 VDD2.n78 585
R1269 VDD2.n19 VDD2.n18 585
R1270 VDD2.n16 VDD2.n15 585
R1271 VDD2.n25 VDD2.n24 585
R1272 VDD2.n27 VDD2.n26 585
R1273 VDD2.n12 VDD2.n11 585
R1274 VDD2.n33 VDD2.n32 585
R1275 VDD2.n36 VDD2.n35 585
R1276 VDD2.n34 VDD2.n8 585
R1277 VDD2.n41 VDD2.n7 585
R1278 VDD2.n43 VDD2.n42 585
R1279 VDD2.n45 VDD2.n44 585
R1280 VDD2.n4 VDD2.n3 585
R1281 VDD2.n51 VDD2.n50 585
R1282 VDD2.n53 VDD2.n52 585
R1283 VDD2.t0 VDD2.n77 329.038
R1284 VDD2.t3 VDD2.n17 329.038
R1285 VDD2.n111 VDD2.n110 171.744
R1286 VDD2.n110 VDD2.n62 171.744
R1287 VDD2.n103 VDD2.n62 171.744
R1288 VDD2.n103 VDD2.n102 171.744
R1289 VDD2.n102 VDD2.n66 171.744
R1290 VDD2.n70 VDD2.n66 171.744
R1291 VDD2.n94 VDD2.n70 171.744
R1292 VDD2.n94 VDD2.n93 171.744
R1293 VDD2.n93 VDD2.n71 171.744
R1294 VDD2.n86 VDD2.n71 171.744
R1295 VDD2.n86 VDD2.n85 171.744
R1296 VDD2.n85 VDD2.n75 171.744
R1297 VDD2.n78 VDD2.n75 171.744
R1298 VDD2.n18 VDD2.n15 171.744
R1299 VDD2.n25 VDD2.n15 171.744
R1300 VDD2.n26 VDD2.n25 171.744
R1301 VDD2.n26 VDD2.n11 171.744
R1302 VDD2.n33 VDD2.n11 171.744
R1303 VDD2.n35 VDD2.n33 171.744
R1304 VDD2.n35 VDD2.n34 171.744
R1305 VDD2.n34 VDD2.n7 171.744
R1306 VDD2.n43 VDD2.n7 171.744
R1307 VDD2.n44 VDD2.n43 171.744
R1308 VDD2.n44 VDD2.n3 171.744
R1309 VDD2.n51 VDD2.n3 171.744
R1310 VDD2.n52 VDD2.n51 171.744
R1311 VDD2.n78 VDD2.t0 85.8723
R1312 VDD2.n18 VDD2.t3 85.8723
R1313 VDD2.n58 VDD2.n57 76.2633
R1314 VDD2 VDD2.n117 76.2604
R1315 VDD2.n58 VDD2.n56 50.9425
R1316 VDD2.n116 VDD2.n115 48.4763
R1317 VDD2.n116 VDD2.n58 43.8317
R1318 VDD2.n101 VDD2.n100 13.1884
R1319 VDD2.n42 VDD2.n41 13.1884
R1320 VDD2.n104 VDD2.n65 12.8005
R1321 VDD2.n99 VDD2.n67 12.8005
R1322 VDD2.n40 VDD2.n8 12.8005
R1323 VDD2.n45 VDD2.n6 12.8005
R1324 VDD2.n105 VDD2.n63 12.0247
R1325 VDD2.n96 VDD2.n95 12.0247
R1326 VDD2.n37 VDD2.n36 12.0247
R1327 VDD2.n46 VDD2.n4 12.0247
R1328 VDD2.n109 VDD2.n108 11.249
R1329 VDD2.n92 VDD2.n69 11.249
R1330 VDD2.n32 VDD2.n10 11.249
R1331 VDD2.n50 VDD2.n49 11.249
R1332 VDD2.n79 VDD2.n77 10.7239
R1333 VDD2.n19 VDD2.n17 10.7239
R1334 VDD2.n112 VDD2.n61 10.4732
R1335 VDD2.n91 VDD2.n72 10.4732
R1336 VDD2.n31 VDD2.n12 10.4732
R1337 VDD2.n53 VDD2.n2 10.4732
R1338 VDD2.n113 VDD2.n59 9.69747
R1339 VDD2.n88 VDD2.n87 9.69747
R1340 VDD2.n28 VDD2.n27 9.69747
R1341 VDD2.n54 VDD2.n0 9.69747
R1342 VDD2.n115 VDD2.n114 9.45567
R1343 VDD2.n56 VDD2.n55 9.45567
R1344 VDD2.n81 VDD2.n80 9.3005
R1345 VDD2.n83 VDD2.n82 9.3005
R1346 VDD2.n74 VDD2.n73 9.3005
R1347 VDD2.n89 VDD2.n88 9.3005
R1348 VDD2.n91 VDD2.n90 9.3005
R1349 VDD2.n69 VDD2.n68 9.3005
R1350 VDD2.n97 VDD2.n96 9.3005
R1351 VDD2.n99 VDD2.n98 9.3005
R1352 VDD2.n114 VDD2.n113 9.3005
R1353 VDD2.n61 VDD2.n60 9.3005
R1354 VDD2.n108 VDD2.n107 9.3005
R1355 VDD2.n106 VDD2.n105 9.3005
R1356 VDD2.n65 VDD2.n64 9.3005
R1357 VDD2.n55 VDD2.n54 9.3005
R1358 VDD2.n2 VDD2.n1 9.3005
R1359 VDD2.n49 VDD2.n48 9.3005
R1360 VDD2.n47 VDD2.n46 9.3005
R1361 VDD2.n6 VDD2.n5 9.3005
R1362 VDD2.n21 VDD2.n20 9.3005
R1363 VDD2.n23 VDD2.n22 9.3005
R1364 VDD2.n14 VDD2.n13 9.3005
R1365 VDD2.n29 VDD2.n28 9.3005
R1366 VDD2.n31 VDD2.n30 9.3005
R1367 VDD2.n10 VDD2.n9 9.3005
R1368 VDD2.n38 VDD2.n37 9.3005
R1369 VDD2.n40 VDD2.n39 9.3005
R1370 VDD2.n84 VDD2.n74 8.92171
R1371 VDD2.n24 VDD2.n14 8.92171
R1372 VDD2.n83 VDD2.n76 8.14595
R1373 VDD2.n23 VDD2.n16 8.14595
R1374 VDD2.n80 VDD2.n79 7.3702
R1375 VDD2.n20 VDD2.n19 7.3702
R1376 VDD2.n80 VDD2.n76 5.81868
R1377 VDD2.n20 VDD2.n16 5.81868
R1378 VDD2.n84 VDD2.n83 5.04292
R1379 VDD2.n24 VDD2.n23 5.04292
R1380 VDD2.n115 VDD2.n59 4.26717
R1381 VDD2.n87 VDD2.n74 4.26717
R1382 VDD2.n27 VDD2.n14 4.26717
R1383 VDD2.n56 VDD2.n0 4.26717
R1384 VDD2.n113 VDD2.n112 3.49141
R1385 VDD2.n88 VDD2.n72 3.49141
R1386 VDD2.n28 VDD2.n12 3.49141
R1387 VDD2.n54 VDD2.n53 3.49141
R1388 VDD2.n117 VDD2.t5 3.04975
R1389 VDD2.n117 VDD2.t2 3.04975
R1390 VDD2.n57 VDD2.t1 3.04975
R1391 VDD2.n57 VDD2.t4 3.04975
R1392 VDD2.n109 VDD2.n61 2.71565
R1393 VDD2.n92 VDD2.n91 2.71565
R1394 VDD2.n32 VDD2.n31 2.71565
R1395 VDD2.n50 VDD2.n2 2.71565
R1396 VDD2 VDD2.n116 2.58024
R1397 VDD2.n81 VDD2.n77 2.41282
R1398 VDD2.n21 VDD2.n17 2.41282
R1399 VDD2.n108 VDD2.n63 1.93989
R1400 VDD2.n95 VDD2.n69 1.93989
R1401 VDD2.n36 VDD2.n10 1.93989
R1402 VDD2.n49 VDD2.n4 1.93989
R1403 VDD2.n105 VDD2.n104 1.16414
R1404 VDD2.n96 VDD2.n67 1.16414
R1405 VDD2.n37 VDD2.n8 1.16414
R1406 VDD2.n46 VDD2.n45 1.16414
R1407 VDD2.n101 VDD2.n65 0.388379
R1408 VDD2.n100 VDD2.n99 0.388379
R1409 VDD2.n41 VDD2.n40 0.388379
R1410 VDD2.n42 VDD2.n6 0.388379
R1411 VDD2.n114 VDD2.n60 0.155672
R1412 VDD2.n107 VDD2.n60 0.155672
R1413 VDD2.n107 VDD2.n106 0.155672
R1414 VDD2.n106 VDD2.n64 0.155672
R1415 VDD2.n98 VDD2.n64 0.155672
R1416 VDD2.n98 VDD2.n97 0.155672
R1417 VDD2.n97 VDD2.n68 0.155672
R1418 VDD2.n90 VDD2.n68 0.155672
R1419 VDD2.n90 VDD2.n89 0.155672
R1420 VDD2.n89 VDD2.n73 0.155672
R1421 VDD2.n82 VDD2.n73 0.155672
R1422 VDD2.n82 VDD2.n81 0.155672
R1423 VDD2.n22 VDD2.n21 0.155672
R1424 VDD2.n22 VDD2.n13 0.155672
R1425 VDD2.n29 VDD2.n13 0.155672
R1426 VDD2.n30 VDD2.n29 0.155672
R1427 VDD2.n30 VDD2.n9 0.155672
R1428 VDD2.n38 VDD2.n9 0.155672
R1429 VDD2.n39 VDD2.n38 0.155672
R1430 VDD2.n39 VDD2.n5 0.155672
R1431 VDD2.n47 VDD2.n5 0.155672
R1432 VDD2.n48 VDD2.n47 0.155672
R1433 VDD2.n48 VDD2.n1 0.155672
R1434 VDD2.n55 VDD2.n1 0.155672
R1435 VTAIL.n234 VTAIL.n182 756.745
R1436 VTAIL.n54 VTAIL.n2 756.745
R1437 VTAIL.n176 VTAIL.n124 756.745
R1438 VTAIL.n116 VTAIL.n64 756.745
R1439 VTAIL.n201 VTAIL.n200 585
R1440 VTAIL.n198 VTAIL.n197 585
R1441 VTAIL.n207 VTAIL.n206 585
R1442 VTAIL.n209 VTAIL.n208 585
R1443 VTAIL.n194 VTAIL.n193 585
R1444 VTAIL.n215 VTAIL.n214 585
R1445 VTAIL.n218 VTAIL.n217 585
R1446 VTAIL.n216 VTAIL.n190 585
R1447 VTAIL.n223 VTAIL.n189 585
R1448 VTAIL.n225 VTAIL.n224 585
R1449 VTAIL.n227 VTAIL.n226 585
R1450 VTAIL.n186 VTAIL.n185 585
R1451 VTAIL.n233 VTAIL.n232 585
R1452 VTAIL.n235 VTAIL.n234 585
R1453 VTAIL.n21 VTAIL.n20 585
R1454 VTAIL.n18 VTAIL.n17 585
R1455 VTAIL.n27 VTAIL.n26 585
R1456 VTAIL.n29 VTAIL.n28 585
R1457 VTAIL.n14 VTAIL.n13 585
R1458 VTAIL.n35 VTAIL.n34 585
R1459 VTAIL.n38 VTAIL.n37 585
R1460 VTAIL.n36 VTAIL.n10 585
R1461 VTAIL.n43 VTAIL.n9 585
R1462 VTAIL.n45 VTAIL.n44 585
R1463 VTAIL.n47 VTAIL.n46 585
R1464 VTAIL.n6 VTAIL.n5 585
R1465 VTAIL.n53 VTAIL.n52 585
R1466 VTAIL.n55 VTAIL.n54 585
R1467 VTAIL.n177 VTAIL.n176 585
R1468 VTAIL.n175 VTAIL.n174 585
R1469 VTAIL.n128 VTAIL.n127 585
R1470 VTAIL.n169 VTAIL.n168 585
R1471 VTAIL.n167 VTAIL.n166 585
R1472 VTAIL.n165 VTAIL.n131 585
R1473 VTAIL.n135 VTAIL.n132 585
R1474 VTAIL.n160 VTAIL.n159 585
R1475 VTAIL.n158 VTAIL.n157 585
R1476 VTAIL.n137 VTAIL.n136 585
R1477 VTAIL.n152 VTAIL.n151 585
R1478 VTAIL.n150 VTAIL.n149 585
R1479 VTAIL.n141 VTAIL.n140 585
R1480 VTAIL.n144 VTAIL.n143 585
R1481 VTAIL.n117 VTAIL.n116 585
R1482 VTAIL.n115 VTAIL.n114 585
R1483 VTAIL.n68 VTAIL.n67 585
R1484 VTAIL.n109 VTAIL.n108 585
R1485 VTAIL.n107 VTAIL.n106 585
R1486 VTAIL.n105 VTAIL.n71 585
R1487 VTAIL.n75 VTAIL.n72 585
R1488 VTAIL.n100 VTAIL.n99 585
R1489 VTAIL.n98 VTAIL.n97 585
R1490 VTAIL.n77 VTAIL.n76 585
R1491 VTAIL.n92 VTAIL.n91 585
R1492 VTAIL.n90 VTAIL.n89 585
R1493 VTAIL.n81 VTAIL.n80 585
R1494 VTAIL.n84 VTAIL.n83 585
R1495 VTAIL.t4 VTAIL.n142 329.038
R1496 VTAIL.t9 VTAIL.n82 329.038
R1497 VTAIL.t7 VTAIL.n199 329.038
R1498 VTAIL.t0 VTAIL.n19 329.038
R1499 VTAIL.n200 VTAIL.n197 171.744
R1500 VTAIL.n207 VTAIL.n197 171.744
R1501 VTAIL.n208 VTAIL.n207 171.744
R1502 VTAIL.n208 VTAIL.n193 171.744
R1503 VTAIL.n215 VTAIL.n193 171.744
R1504 VTAIL.n217 VTAIL.n215 171.744
R1505 VTAIL.n217 VTAIL.n216 171.744
R1506 VTAIL.n216 VTAIL.n189 171.744
R1507 VTAIL.n225 VTAIL.n189 171.744
R1508 VTAIL.n226 VTAIL.n225 171.744
R1509 VTAIL.n226 VTAIL.n185 171.744
R1510 VTAIL.n233 VTAIL.n185 171.744
R1511 VTAIL.n234 VTAIL.n233 171.744
R1512 VTAIL.n20 VTAIL.n17 171.744
R1513 VTAIL.n27 VTAIL.n17 171.744
R1514 VTAIL.n28 VTAIL.n27 171.744
R1515 VTAIL.n28 VTAIL.n13 171.744
R1516 VTAIL.n35 VTAIL.n13 171.744
R1517 VTAIL.n37 VTAIL.n35 171.744
R1518 VTAIL.n37 VTAIL.n36 171.744
R1519 VTAIL.n36 VTAIL.n9 171.744
R1520 VTAIL.n45 VTAIL.n9 171.744
R1521 VTAIL.n46 VTAIL.n45 171.744
R1522 VTAIL.n46 VTAIL.n5 171.744
R1523 VTAIL.n53 VTAIL.n5 171.744
R1524 VTAIL.n54 VTAIL.n53 171.744
R1525 VTAIL.n176 VTAIL.n175 171.744
R1526 VTAIL.n175 VTAIL.n127 171.744
R1527 VTAIL.n168 VTAIL.n127 171.744
R1528 VTAIL.n168 VTAIL.n167 171.744
R1529 VTAIL.n167 VTAIL.n131 171.744
R1530 VTAIL.n135 VTAIL.n131 171.744
R1531 VTAIL.n159 VTAIL.n135 171.744
R1532 VTAIL.n159 VTAIL.n158 171.744
R1533 VTAIL.n158 VTAIL.n136 171.744
R1534 VTAIL.n151 VTAIL.n136 171.744
R1535 VTAIL.n151 VTAIL.n150 171.744
R1536 VTAIL.n150 VTAIL.n140 171.744
R1537 VTAIL.n143 VTAIL.n140 171.744
R1538 VTAIL.n116 VTAIL.n115 171.744
R1539 VTAIL.n115 VTAIL.n67 171.744
R1540 VTAIL.n108 VTAIL.n67 171.744
R1541 VTAIL.n108 VTAIL.n107 171.744
R1542 VTAIL.n107 VTAIL.n71 171.744
R1543 VTAIL.n75 VTAIL.n71 171.744
R1544 VTAIL.n99 VTAIL.n75 171.744
R1545 VTAIL.n99 VTAIL.n98 171.744
R1546 VTAIL.n98 VTAIL.n76 171.744
R1547 VTAIL.n91 VTAIL.n76 171.744
R1548 VTAIL.n91 VTAIL.n90 171.744
R1549 VTAIL.n90 VTAIL.n80 171.744
R1550 VTAIL.n83 VTAIL.n80 171.744
R1551 VTAIL.n200 VTAIL.t7 85.8723
R1552 VTAIL.n20 VTAIL.t0 85.8723
R1553 VTAIL.n143 VTAIL.t4 85.8723
R1554 VTAIL.n83 VTAIL.t9 85.8723
R1555 VTAIL.n123 VTAIL.n122 58.7995
R1556 VTAIL.n63 VTAIL.n62 58.7995
R1557 VTAIL.n1 VTAIL.n0 58.7993
R1558 VTAIL.n61 VTAIL.n60 58.7993
R1559 VTAIL.n239 VTAIL.n238 31.7975
R1560 VTAIL.n59 VTAIL.n58 31.7975
R1561 VTAIL.n181 VTAIL.n180 31.7975
R1562 VTAIL.n121 VTAIL.n120 31.7975
R1563 VTAIL.n63 VTAIL.n61 28.2807
R1564 VTAIL.n239 VTAIL.n181 24.9186
R1565 VTAIL.n224 VTAIL.n223 13.1884
R1566 VTAIL.n44 VTAIL.n43 13.1884
R1567 VTAIL.n166 VTAIL.n165 13.1884
R1568 VTAIL.n106 VTAIL.n105 13.1884
R1569 VTAIL.n222 VTAIL.n190 12.8005
R1570 VTAIL.n227 VTAIL.n188 12.8005
R1571 VTAIL.n42 VTAIL.n10 12.8005
R1572 VTAIL.n47 VTAIL.n8 12.8005
R1573 VTAIL.n169 VTAIL.n130 12.8005
R1574 VTAIL.n164 VTAIL.n132 12.8005
R1575 VTAIL.n109 VTAIL.n70 12.8005
R1576 VTAIL.n104 VTAIL.n72 12.8005
R1577 VTAIL.n219 VTAIL.n218 12.0247
R1578 VTAIL.n228 VTAIL.n186 12.0247
R1579 VTAIL.n39 VTAIL.n38 12.0247
R1580 VTAIL.n48 VTAIL.n6 12.0247
R1581 VTAIL.n170 VTAIL.n128 12.0247
R1582 VTAIL.n161 VTAIL.n160 12.0247
R1583 VTAIL.n110 VTAIL.n68 12.0247
R1584 VTAIL.n101 VTAIL.n100 12.0247
R1585 VTAIL.n214 VTAIL.n192 11.249
R1586 VTAIL.n232 VTAIL.n231 11.249
R1587 VTAIL.n34 VTAIL.n12 11.249
R1588 VTAIL.n52 VTAIL.n51 11.249
R1589 VTAIL.n174 VTAIL.n173 11.249
R1590 VTAIL.n157 VTAIL.n134 11.249
R1591 VTAIL.n114 VTAIL.n113 11.249
R1592 VTAIL.n97 VTAIL.n74 11.249
R1593 VTAIL.n201 VTAIL.n199 10.7239
R1594 VTAIL.n21 VTAIL.n19 10.7239
R1595 VTAIL.n144 VTAIL.n142 10.7239
R1596 VTAIL.n84 VTAIL.n82 10.7239
R1597 VTAIL.n213 VTAIL.n194 10.4732
R1598 VTAIL.n235 VTAIL.n184 10.4732
R1599 VTAIL.n33 VTAIL.n14 10.4732
R1600 VTAIL.n55 VTAIL.n4 10.4732
R1601 VTAIL.n177 VTAIL.n126 10.4732
R1602 VTAIL.n156 VTAIL.n137 10.4732
R1603 VTAIL.n117 VTAIL.n66 10.4732
R1604 VTAIL.n96 VTAIL.n77 10.4732
R1605 VTAIL.n210 VTAIL.n209 9.69747
R1606 VTAIL.n236 VTAIL.n182 9.69747
R1607 VTAIL.n30 VTAIL.n29 9.69747
R1608 VTAIL.n56 VTAIL.n2 9.69747
R1609 VTAIL.n178 VTAIL.n124 9.69747
R1610 VTAIL.n153 VTAIL.n152 9.69747
R1611 VTAIL.n118 VTAIL.n64 9.69747
R1612 VTAIL.n93 VTAIL.n92 9.69747
R1613 VTAIL.n238 VTAIL.n237 9.45567
R1614 VTAIL.n58 VTAIL.n57 9.45567
R1615 VTAIL.n180 VTAIL.n179 9.45567
R1616 VTAIL.n120 VTAIL.n119 9.45567
R1617 VTAIL.n237 VTAIL.n236 9.3005
R1618 VTAIL.n184 VTAIL.n183 9.3005
R1619 VTAIL.n231 VTAIL.n230 9.3005
R1620 VTAIL.n229 VTAIL.n228 9.3005
R1621 VTAIL.n188 VTAIL.n187 9.3005
R1622 VTAIL.n203 VTAIL.n202 9.3005
R1623 VTAIL.n205 VTAIL.n204 9.3005
R1624 VTAIL.n196 VTAIL.n195 9.3005
R1625 VTAIL.n211 VTAIL.n210 9.3005
R1626 VTAIL.n213 VTAIL.n212 9.3005
R1627 VTAIL.n192 VTAIL.n191 9.3005
R1628 VTAIL.n220 VTAIL.n219 9.3005
R1629 VTAIL.n222 VTAIL.n221 9.3005
R1630 VTAIL.n57 VTAIL.n56 9.3005
R1631 VTAIL.n4 VTAIL.n3 9.3005
R1632 VTAIL.n51 VTAIL.n50 9.3005
R1633 VTAIL.n49 VTAIL.n48 9.3005
R1634 VTAIL.n8 VTAIL.n7 9.3005
R1635 VTAIL.n23 VTAIL.n22 9.3005
R1636 VTAIL.n25 VTAIL.n24 9.3005
R1637 VTAIL.n16 VTAIL.n15 9.3005
R1638 VTAIL.n31 VTAIL.n30 9.3005
R1639 VTAIL.n33 VTAIL.n32 9.3005
R1640 VTAIL.n12 VTAIL.n11 9.3005
R1641 VTAIL.n40 VTAIL.n39 9.3005
R1642 VTAIL.n42 VTAIL.n41 9.3005
R1643 VTAIL.n146 VTAIL.n145 9.3005
R1644 VTAIL.n148 VTAIL.n147 9.3005
R1645 VTAIL.n139 VTAIL.n138 9.3005
R1646 VTAIL.n154 VTAIL.n153 9.3005
R1647 VTAIL.n156 VTAIL.n155 9.3005
R1648 VTAIL.n134 VTAIL.n133 9.3005
R1649 VTAIL.n162 VTAIL.n161 9.3005
R1650 VTAIL.n164 VTAIL.n163 9.3005
R1651 VTAIL.n179 VTAIL.n178 9.3005
R1652 VTAIL.n126 VTAIL.n125 9.3005
R1653 VTAIL.n173 VTAIL.n172 9.3005
R1654 VTAIL.n171 VTAIL.n170 9.3005
R1655 VTAIL.n130 VTAIL.n129 9.3005
R1656 VTAIL.n86 VTAIL.n85 9.3005
R1657 VTAIL.n88 VTAIL.n87 9.3005
R1658 VTAIL.n79 VTAIL.n78 9.3005
R1659 VTAIL.n94 VTAIL.n93 9.3005
R1660 VTAIL.n96 VTAIL.n95 9.3005
R1661 VTAIL.n74 VTAIL.n73 9.3005
R1662 VTAIL.n102 VTAIL.n101 9.3005
R1663 VTAIL.n104 VTAIL.n103 9.3005
R1664 VTAIL.n119 VTAIL.n118 9.3005
R1665 VTAIL.n66 VTAIL.n65 9.3005
R1666 VTAIL.n113 VTAIL.n112 9.3005
R1667 VTAIL.n111 VTAIL.n110 9.3005
R1668 VTAIL.n70 VTAIL.n69 9.3005
R1669 VTAIL.n206 VTAIL.n196 8.92171
R1670 VTAIL.n26 VTAIL.n16 8.92171
R1671 VTAIL.n149 VTAIL.n139 8.92171
R1672 VTAIL.n89 VTAIL.n79 8.92171
R1673 VTAIL.n205 VTAIL.n198 8.14595
R1674 VTAIL.n25 VTAIL.n18 8.14595
R1675 VTAIL.n148 VTAIL.n141 8.14595
R1676 VTAIL.n88 VTAIL.n81 8.14595
R1677 VTAIL.n202 VTAIL.n201 7.3702
R1678 VTAIL.n22 VTAIL.n21 7.3702
R1679 VTAIL.n145 VTAIL.n144 7.3702
R1680 VTAIL.n85 VTAIL.n84 7.3702
R1681 VTAIL.n202 VTAIL.n198 5.81868
R1682 VTAIL.n22 VTAIL.n18 5.81868
R1683 VTAIL.n145 VTAIL.n141 5.81868
R1684 VTAIL.n85 VTAIL.n81 5.81868
R1685 VTAIL.n206 VTAIL.n205 5.04292
R1686 VTAIL.n26 VTAIL.n25 5.04292
R1687 VTAIL.n149 VTAIL.n148 5.04292
R1688 VTAIL.n89 VTAIL.n88 5.04292
R1689 VTAIL.n209 VTAIL.n196 4.26717
R1690 VTAIL.n238 VTAIL.n182 4.26717
R1691 VTAIL.n29 VTAIL.n16 4.26717
R1692 VTAIL.n58 VTAIL.n2 4.26717
R1693 VTAIL.n180 VTAIL.n124 4.26717
R1694 VTAIL.n152 VTAIL.n139 4.26717
R1695 VTAIL.n120 VTAIL.n64 4.26717
R1696 VTAIL.n92 VTAIL.n79 4.26717
R1697 VTAIL.n210 VTAIL.n194 3.49141
R1698 VTAIL.n236 VTAIL.n235 3.49141
R1699 VTAIL.n30 VTAIL.n14 3.49141
R1700 VTAIL.n56 VTAIL.n55 3.49141
R1701 VTAIL.n178 VTAIL.n177 3.49141
R1702 VTAIL.n153 VTAIL.n137 3.49141
R1703 VTAIL.n118 VTAIL.n117 3.49141
R1704 VTAIL.n93 VTAIL.n77 3.49141
R1705 VTAIL.n121 VTAIL.n63 3.36257
R1706 VTAIL.n181 VTAIL.n123 3.36257
R1707 VTAIL.n61 VTAIL.n59 3.36257
R1708 VTAIL.n0 VTAIL.t10 3.04975
R1709 VTAIL.n0 VTAIL.t11 3.04975
R1710 VTAIL.n60 VTAIL.t5 3.04975
R1711 VTAIL.n60 VTAIL.t3 3.04975
R1712 VTAIL.n122 VTAIL.t1 3.04975
R1713 VTAIL.n122 VTAIL.t2 3.04975
R1714 VTAIL.n62 VTAIL.t6 3.04975
R1715 VTAIL.n62 VTAIL.t8 3.04975
R1716 VTAIL.n214 VTAIL.n213 2.71565
R1717 VTAIL.n232 VTAIL.n184 2.71565
R1718 VTAIL.n34 VTAIL.n33 2.71565
R1719 VTAIL.n52 VTAIL.n4 2.71565
R1720 VTAIL.n174 VTAIL.n126 2.71565
R1721 VTAIL.n157 VTAIL.n156 2.71565
R1722 VTAIL.n114 VTAIL.n66 2.71565
R1723 VTAIL.n97 VTAIL.n96 2.71565
R1724 VTAIL VTAIL.n239 2.46386
R1725 VTAIL.n203 VTAIL.n199 2.41282
R1726 VTAIL.n23 VTAIL.n19 2.41282
R1727 VTAIL.n146 VTAIL.n142 2.41282
R1728 VTAIL.n86 VTAIL.n82 2.41282
R1729 VTAIL.n123 VTAIL.n121 2.15136
R1730 VTAIL.n59 VTAIL.n1 2.15136
R1731 VTAIL.n218 VTAIL.n192 1.93989
R1732 VTAIL.n231 VTAIL.n186 1.93989
R1733 VTAIL.n38 VTAIL.n12 1.93989
R1734 VTAIL.n51 VTAIL.n6 1.93989
R1735 VTAIL.n173 VTAIL.n128 1.93989
R1736 VTAIL.n160 VTAIL.n134 1.93989
R1737 VTAIL.n113 VTAIL.n68 1.93989
R1738 VTAIL.n100 VTAIL.n74 1.93989
R1739 VTAIL.n219 VTAIL.n190 1.16414
R1740 VTAIL.n228 VTAIL.n227 1.16414
R1741 VTAIL.n39 VTAIL.n10 1.16414
R1742 VTAIL.n48 VTAIL.n47 1.16414
R1743 VTAIL.n170 VTAIL.n169 1.16414
R1744 VTAIL.n161 VTAIL.n132 1.16414
R1745 VTAIL.n110 VTAIL.n109 1.16414
R1746 VTAIL.n101 VTAIL.n72 1.16414
R1747 VTAIL VTAIL.n1 0.899207
R1748 VTAIL.n223 VTAIL.n222 0.388379
R1749 VTAIL.n224 VTAIL.n188 0.388379
R1750 VTAIL.n43 VTAIL.n42 0.388379
R1751 VTAIL.n44 VTAIL.n8 0.388379
R1752 VTAIL.n166 VTAIL.n130 0.388379
R1753 VTAIL.n165 VTAIL.n164 0.388379
R1754 VTAIL.n106 VTAIL.n70 0.388379
R1755 VTAIL.n105 VTAIL.n104 0.388379
R1756 VTAIL.n204 VTAIL.n203 0.155672
R1757 VTAIL.n204 VTAIL.n195 0.155672
R1758 VTAIL.n211 VTAIL.n195 0.155672
R1759 VTAIL.n212 VTAIL.n211 0.155672
R1760 VTAIL.n212 VTAIL.n191 0.155672
R1761 VTAIL.n220 VTAIL.n191 0.155672
R1762 VTAIL.n221 VTAIL.n220 0.155672
R1763 VTAIL.n221 VTAIL.n187 0.155672
R1764 VTAIL.n229 VTAIL.n187 0.155672
R1765 VTAIL.n230 VTAIL.n229 0.155672
R1766 VTAIL.n230 VTAIL.n183 0.155672
R1767 VTAIL.n237 VTAIL.n183 0.155672
R1768 VTAIL.n24 VTAIL.n23 0.155672
R1769 VTAIL.n24 VTAIL.n15 0.155672
R1770 VTAIL.n31 VTAIL.n15 0.155672
R1771 VTAIL.n32 VTAIL.n31 0.155672
R1772 VTAIL.n32 VTAIL.n11 0.155672
R1773 VTAIL.n40 VTAIL.n11 0.155672
R1774 VTAIL.n41 VTAIL.n40 0.155672
R1775 VTAIL.n41 VTAIL.n7 0.155672
R1776 VTAIL.n49 VTAIL.n7 0.155672
R1777 VTAIL.n50 VTAIL.n49 0.155672
R1778 VTAIL.n50 VTAIL.n3 0.155672
R1779 VTAIL.n57 VTAIL.n3 0.155672
R1780 VTAIL.n179 VTAIL.n125 0.155672
R1781 VTAIL.n172 VTAIL.n125 0.155672
R1782 VTAIL.n172 VTAIL.n171 0.155672
R1783 VTAIL.n171 VTAIL.n129 0.155672
R1784 VTAIL.n163 VTAIL.n129 0.155672
R1785 VTAIL.n163 VTAIL.n162 0.155672
R1786 VTAIL.n162 VTAIL.n133 0.155672
R1787 VTAIL.n155 VTAIL.n133 0.155672
R1788 VTAIL.n155 VTAIL.n154 0.155672
R1789 VTAIL.n154 VTAIL.n138 0.155672
R1790 VTAIL.n147 VTAIL.n138 0.155672
R1791 VTAIL.n147 VTAIL.n146 0.155672
R1792 VTAIL.n119 VTAIL.n65 0.155672
R1793 VTAIL.n112 VTAIL.n65 0.155672
R1794 VTAIL.n112 VTAIL.n111 0.155672
R1795 VTAIL.n111 VTAIL.n69 0.155672
R1796 VTAIL.n103 VTAIL.n69 0.155672
R1797 VTAIL.n103 VTAIL.n102 0.155672
R1798 VTAIL.n102 VTAIL.n73 0.155672
R1799 VTAIL.n95 VTAIL.n73 0.155672
R1800 VTAIL.n95 VTAIL.n94 0.155672
R1801 VTAIL.n94 VTAIL.n78 0.155672
R1802 VTAIL.n87 VTAIL.n78 0.155672
R1803 VTAIL.n87 VTAIL.n86 0.155672
R1804 VP.n16 VP.n13 161.3
R1805 VP.n18 VP.n17 161.3
R1806 VP.n19 VP.n12 161.3
R1807 VP.n21 VP.n20 161.3
R1808 VP.n22 VP.n11 161.3
R1809 VP.n24 VP.n23 161.3
R1810 VP.n25 VP.n10 161.3
R1811 VP.n27 VP.n26 161.3
R1812 VP.n55 VP.n54 161.3
R1813 VP.n53 VP.n1 161.3
R1814 VP.n52 VP.n51 161.3
R1815 VP.n50 VP.n2 161.3
R1816 VP.n49 VP.n48 161.3
R1817 VP.n47 VP.n3 161.3
R1818 VP.n46 VP.n45 161.3
R1819 VP.n44 VP.n4 161.3
R1820 VP.n43 VP.n42 161.3
R1821 VP.n40 VP.n5 161.3
R1822 VP.n39 VP.n38 161.3
R1823 VP.n37 VP.n6 161.3
R1824 VP.n36 VP.n35 161.3
R1825 VP.n34 VP.n7 161.3
R1826 VP.n33 VP.n32 161.3
R1827 VP.n31 VP.n8 161.3
R1828 VP.n15 VP.t3 104.975
R1829 VP.n30 VP.n29 82.868
R1830 VP.n56 VP.n0 82.868
R1831 VP.n28 VP.n9 82.868
R1832 VP.n29 VP.t1 71.963
R1833 VP.n41 VP.t5 71.963
R1834 VP.n0 VP.t0 71.963
R1835 VP.n9 VP.t2 71.963
R1836 VP.n14 VP.t4 71.963
R1837 VP.n15 VP.n14 62.4546
R1838 VP.n35 VP.n6 56.5617
R1839 VP.n48 VP.n2 56.5617
R1840 VP.n20 VP.n11 56.5617
R1841 VP.n30 VP.n28 51.5299
R1842 VP.n33 VP.n8 24.5923
R1843 VP.n34 VP.n33 24.5923
R1844 VP.n35 VP.n34 24.5923
R1845 VP.n39 VP.n6 24.5923
R1846 VP.n40 VP.n39 24.5923
R1847 VP.n42 VP.n40 24.5923
R1848 VP.n46 VP.n4 24.5923
R1849 VP.n47 VP.n46 24.5923
R1850 VP.n48 VP.n47 24.5923
R1851 VP.n52 VP.n2 24.5923
R1852 VP.n53 VP.n52 24.5923
R1853 VP.n54 VP.n53 24.5923
R1854 VP.n24 VP.n11 24.5923
R1855 VP.n25 VP.n24 24.5923
R1856 VP.n26 VP.n25 24.5923
R1857 VP.n18 VP.n13 24.5923
R1858 VP.n19 VP.n18 24.5923
R1859 VP.n20 VP.n19 24.5923
R1860 VP.n42 VP.n41 12.2964
R1861 VP.n41 VP.n4 12.2964
R1862 VP.n14 VP.n13 12.2964
R1863 VP.n29 VP.n8 7.37805
R1864 VP.n54 VP.n0 7.37805
R1865 VP.n26 VP.n9 7.37805
R1866 VP.n16 VP.n15 3.2308
R1867 VP.n28 VP.n27 0.354861
R1868 VP.n31 VP.n30 0.354861
R1869 VP.n56 VP.n55 0.354861
R1870 VP VP.n56 0.267071
R1871 VP.n17 VP.n16 0.189894
R1872 VP.n17 VP.n12 0.189894
R1873 VP.n21 VP.n12 0.189894
R1874 VP.n22 VP.n21 0.189894
R1875 VP.n23 VP.n22 0.189894
R1876 VP.n23 VP.n10 0.189894
R1877 VP.n27 VP.n10 0.189894
R1878 VP.n32 VP.n31 0.189894
R1879 VP.n32 VP.n7 0.189894
R1880 VP.n36 VP.n7 0.189894
R1881 VP.n37 VP.n36 0.189894
R1882 VP.n38 VP.n37 0.189894
R1883 VP.n38 VP.n5 0.189894
R1884 VP.n43 VP.n5 0.189894
R1885 VP.n44 VP.n43 0.189894
R1886 VP.n45 VP.n44 0.189894
R1887 VP.n45 VP.n3 0.189894
R1888 VP.n49 VP.n3 0.189894
R1889 VP.n50 VP.n49 0.189894
R1890 VP.n51 VP.n50 0.189894
R1891 VP.n51 VP.n1 0.189894
R1892 VP.n55 VP.n1 0.189894
R1893 VDD1.n52 VDD1.n0 756.745
R1894 VDD1.n109 VDD1.n57 756.745
R1895 VDD1.n53 VDD1.n52 585
R1896 VDD1.n51 VDD1.n50 585
R1897 VDD1.n4 VDD1.n3 585
R1898 VDD1.n45 VDD1.n44 585
R1899 VDD1.n43 VDD1.n42 585
R1900 VDD1.n41 VDD1.n7 585
R1901 VDD1.n11 VDD1.n8 585
R1902 VDD1.n36 VDD1.n35 585
R1903 VDD1.n34 VDD1.n33 585
R1904 VDD1.n13 VDD1.n12 585
R1905 VDD1.n28 VDD1.n27 585
R1906 VDD1.n26 VDD1.n25 585
R1907 VDD1.n17 VDD1.n16 585
R1908 VDD1.n20 VDD1.n19 585
R1909 VDD1.n76 VDD1.n75 585
R1910 VDD1.n73 VDD1.n72 585
R1911 VDD1.n82 VDD1.n81 585
R1912 VDD1.n84 VDD1.n83 585
R1913 VDD1.n69 VDD1.n68 585
R1914 VDD1.n90 VDD1.n89 585
R1915 VDD1.n93 VDD1.n92 585
R1916 VDD1.n91 VDD1.n65 585
R1917 VDD1.n98 VDD1.n64 585
R1918 VDD1.n100 VDD1.n99 585
R1919 VDD1.n102 VDD1.n101 585
R1920 VDD1.n61 VDD1.n60 585
R1921 VDD1.n108 VDD1.n107 585
R1922 VDD1.n110 VDD1.n109 585
R1923 VDD1.t2 VDD1.n18 329.038
R1924 VDD1.t4 VDD1.n74 329.038
R1925 VDD1.n52 VDD1.n51 171.744
R1926 VDD1.n51 VDD1.n3 171.744
R1927 VDD1.n44 VDD1.n3 171.744
R1928 VDD1.n44 VDD1.n43 171.744
R1929 VDD1.n43 VDD1.n7 171.744
R1930 VDD1.n11 VDD1.n7 171.744
R1931 VDD1.n35 VDD1.n11 171.744
R1932 VDD1.n35 VDD1.n34 171.744
R1933 VDD1.n34 VDD1.n12 171.744
R1934 VDD1.n27 VDD1.n12 171.744
R1935 VDD1.n27 VDD1.n26 171.744
R1936 VDD1.n26 VDD1.n16 171.744
R1937 VDD1.n19 VDD1.n16 171.744
R1938 VDD1.n75 VDD1.n72 171.744
R1939 VDD1.n82 VDD1.n72 171.744
R1940 VDD1.n83 VDD1.n82 171.744
R1941 VDD1.n83 VDD1.n68 171.744
R1942 VDD1.n90 VDD1.n68 171.744
R1943 VDD1.n92 VDD1.n90 171.744
R1944 VDD1.n92 VDD1.n91 171.744
R1945 VDD1.n91 VDD1.n64 171.744
R1946 VDD1.n100 VDD1.n64 171.744
R1947 VDD1.n101 VDD1.n100 171.744
R1948 VDD1.n101 VDD1.n60 171.744
R1949 VDD1.n108 VDD1.n60 171.744
R1950 VDD1.n109 VDD1.n108 171.744
R1951 VDD1.n19 VDD1.t2 85.8723
R1952 VDD1.n75 VDD1.t4 85.8723
R1953 VDD1.n115 VDD1.n114 76.2633
R1954 VDD1.n117 VDD1.n116 75.4781
R1955 VDD1 VDD1.n56 51.056
R1956 VDD1.n115 VDD1.n113 50.9425
R1957 VDD1.n117 VDD1.n115 46.0957
R1958 VDD1.n42 VDD1.n41 13.1884
R1959 VDD1.n99 VDD1.n98 13.1884
R1960 VDD1.n45 VDD1.n6 12.8005
R1961 VDD1.n40 VDD1.n8 12.8005
R1962 VDD1.n97 VDD1.n65 12.8005
R1963 VDD1.n102 VDD1.n63 12.8005
R1964 VDD1.n46 VDD1.n4 12.0247
R1965 VDD1.n37 VDD1.n36 12.0247
R1966 VDD1.n94 VDD1.n93 12.0247
R1967 VDD1.n103 VDD1.n61 12.0247
R1968 VDD1.n50 VDD1.n49 11.249
R1969 VDD1.n33 VDD1.n10 11.249
R1970 VDD1.n89 VDD1.n67 11.249
R1971 VDD1.n107 VDD1.n106 11.249
R1972 VDD1.n20 VDD1.n18 10.7239
R1973 VDD1.n76 VDD1.n74 10.7239
R1974 VDD1.n53 VDD1.n2 10.4732
R1975 VDD1.n32 VDD1.n13 10.4732
R1976 VDD1.n88 VDD1.n69 10.4732
R1977 VDD1.n110 VDD1.n59 10.4732
R1978 VDD1.n54 VDD1.n0 9.69747
R1979 VDD1.n29 VDD1.n28 9.69747
R1980 VDD1.n85 VDD1.n84 9.69747
R1981 VDD1.n111 VDD1.n57 9.69747
R1982 VDD1.n56 VDD1.n55 9.45567
R1983 VDD1.n113 VDD1.n112 9.45567
R1984 VDD1.n22 VDD1.n21 9.3005
R1985 VDD1.n24 VDD1.n23 9.3005
R1986 VDD1.n15 VDD1.n14 9.3005
R1987 VDD1.n30 VDD1.n29 9.3005
R1988 VDD1.n32 VDD1.n31 9.3005
R1989 VDD1.n10 VDD1.n9 9.3005
R1990 VDD1.n38 VDD1.n37 9.3005
R1991 VDD1.n40 VDD1.n39 9.3005
R1992 VDD1.n55 VDD1.n54 9.3005
R1993 VDD1.n2 VDD1.n1 9.3005
R1994 VDD1.n49 VDD1.n48 9.3005
R1995 VDD1.n47 VDD1.n46 9.3005
R1996 VDD1.n6 VDD1.n5 9.3005
R1997 VDD1.n112 VDD1.n111 9.3005
R1998 VDD1.n59 VDD1.n58 9.3005
R1999 VDD1.n106 VDD1.n105 9.3005
R2000 VDD1.n104 VDD1.n103 9.3005
R2001 VDD1.n63 VDD1.n62 9.3005
R2002 VDD1.n78 VDD1.n77 9.3005
R2003 VDD1.n80 VDD1.n79 9.3005
R2004 VDD1.n71 VDD1.n70 9.3005
R2005 VDD1.n86 VDD1.n85 9.3005
R2006 VDD1.n88 VDD1.n87 9.3005
R2007 VDD1.n67 VDD1.n66 9.3005
R2008 VDD1.n95 VDD1.n94 9.3005
R2009 VDD1.n97 VDD1.n96 9.3005
R2010 VDD1.n25 VDD1.n15 8.92171
R2011 VDD1.n81 VDD1.n71 8.92171
R2012 VDD1.n24 VDD1.n17 8.14595
R2013 VDD1.n80 VDD1.n73 8.14595
R2014 VDD1.n21 VDD1.n20 7.3702
R2015 VDD1.n77 VDD1.n76 7.3702
R2016 VDD1.n21 VDD1.n17 5.81868
R2017 VDD1.n77 VDD1.n73 5.81868
R2018 VDD1.n25 VDD1.n24 5.04292
R2019 VDD1.n81 VDD1.n80 5.04292
R2020 VDD1.n56 VDD1.n0 4.26717
R2021 VDD1.n28 VDD1.n15 4.26717
R2022 VDD1.n84 VDD1.n71 4.26717
R2023 VDD1.n113 VDD1.n57 4.26717
R2024 VDD1.n54 VDD1.n53 3.49141
R2025 VDD1.n29 VDD1.n13 3.49141
R2026 VDD1.n85 VDD1.n69 3.49141
R2027 VDD1.n111 VDD1.n110 3.49141
R2028 VDD1.n116 VDD1.t1 3.04975
R2029 VDD1.n116 VDD1.t3 3.04975
R2030 VDD1.n114 VDD1.t0 3.04975
R2031 VDD1.n114 VDD1.t5 3.04975
R2032 VDD1.n50 VDD1.n2 2.71565
R2033 VDD1.n33 VDD1.n32 2.71565
R2034 VDD1.n89 VDD1.n88 2.71565
R2035 VDD1.n107 VDD1.n59 2.71565
R2036 VDD1.n22 VDD1.n18 2.41282
R2037 VDD1.n78 VDD1.n74 2.41282
R2038 VDD1.n49 VDD1.n4 1.93989
R2039 VDD1.n36 VDD1.n10 1.93989
R2040 VDD1.n93 VDD1.n67 1.93989
R2041 VDD1.n106 VDD1.n61 1.93989
R2042 VDD1.n46 VDD1.n45 1.16414
R2043 VDD1.n37 VDD1.n8 1.16414
R2044 VDD1.n94 VDD1.n65 1.16414
R2045 VDD1.n103 VDD1.n102 1.16414
R2046 VDD1 VDD1.n117 0.782828
R2047 VDD1.n42 VDD1.n6 0.388379
R2048 VDD1.n41 VDD1.n40 0.388379
R2049 VDD1.n98 VDD1.n97 0.388379
R2050 VDD1.n99 VDD1.n63 0.388379
R2051 VDD1.n55 VDD1.n1 0.155672
R2052 VDD1.n48 VDD1.n1 0.155672
R2053 VDD1.n48 VDD1.n47 0.155672
R2054 VDD1.n47 VDD1.n5 0.155672
R2055 VDD1.n39 VDD1.n5 0.155672
R2056 VDD1.n39 VDD1.n38 0.155672
R2057 VDD1.n38 VDD1.n9 0.155672
R2058 VDD1.n31 VDD1.n9 0.155672
R2059 VDD1.n31 VDD1.n30 0.155672
R2060 VDD1.n30 VDD1.n14 0.155672
R2061 VDD1.n23 VDD1.n14 0.155672
R2062 VDD1.n23 VDD1.n22 0.155672
R2063 VDD1.n79 VDD1.n78 0.155672
R2064 VDD1.n79 VDD1.n70 0.155672
R2065 VDD1.n86 VDD1.n70 0.155672
R2066 VDD1.n87 VDD1.n86 0.155672
R2067 VDD1.n87 VDD1.n66 0.155672
R2068 VDD1.n95 VDD1.n66 0.155672
R2069 VDD1.n96 VDD1.n95 0.155672
R2070 VDD1.n96 VDD1.n62 0.155672
R2071 VDD1.n104 VDD1.n62 0.155672
R2072 VDD1.n105 VDD1.n104 0.155672
R2073 VDD1.n105 VDD1.n58 0.155672
R2074 VDD1.n112 VDD1.n58 0.155672
C0 w_n4090_n3100# VP 8.47953f
C1 VN VP 7.61679f
C2 VDD1 VP 6.72178f
C3 VTAIL VP 6.80689f
C4 VN w_n4090_n3100# 7.94805f
C5 VP VDD2 0.540908f
C6 w_n4090_n3100# VDD1 2.43636f
C7 w_n4090_n3100# VTAIL 2.88182f
C8 B VP 2.253f
C9 VN VDD1 0.152494f
C10 VN VTAIL 6.79266f
C11 VTAIL VDD1 7.61807f
C12 w_n4090_n3100# VDD2 2.55244f
C13 B w_n4090_n3100# 10.6401f
C14 VN VDD2 6.33623f
C15 VDD1 VDD2 1.78601f
C16 VTAIL VDD2 7.67645f
C17 VN B 1.36075f
C18 B VDD1 2.2376f
C19 B VTAIL 3.7411f
C20 B VDD2 2.33495f
C21 VDD2 VSUBS 2.13622f
C22 VDD1 VSUBS 2.131041f
C23 VTAIL VSUBS 1.330599f
C24 VN VSUBS 6.75572f
C25 VP VSUBS 3.643315f
C26 B VSUBS 5.482832f
C27 w_n4090_n3100# VSUBS 0.156418p
C28 VDD1.n0 VSUBS 0.030239f
C29 VDD1.n1 VSUBS 0.028739f
C30 VDD1.n2 VSUBS 0.015443f
C31 VDD1.n3 VSUBS 0.036501f
C32 VDD1.n4 VSUBS 0.016351f
C33 VDD1.n5 VSUBS 0.028739f
C34 VDD1.n6 VSUBS 0.015443f
C35 VDD1.n7 VSUBS 0.036501f
C36 VDD1.n8 VSUBS 0.016351f
C37 VDD1.n9 VSUBS 0.028739f
C38 VDD1.n10 VSUBS 0.015443f
C39 VDD1.n11 VSUBS 0.036501f
C40 VDD1.n12 VSUBS 0.036501f
C41 VDD1.n13 VSUBS 0.016351f
C42 VDD1.n14 VSUBS 0.028739f
C43 VDD1.n15 VSUBS 0.015443f
C44 VDD1.n16 VSUBS 0.036501f
C45 VDD1.n17 VSUBS 0.016351f
C46 VDD1.n18 VSUBS 0.208929f
C47 VDD1.t2 VSUBS 0.078535f
C48 VDD1.n19 VSUBS 0.027376f
C49 VDD1.n20 VSUBS 0.027458f
C50 VDD1.n21 VSUBS 0.015443f
C51 VDD1.n22 VSUBS 1.24327f
C52 VDD1.n23 VSUBS 0.028739f
C53 VDD1.n24 VSUBS 0.015443f
C54 VDD1.n25 VSUBS 0.016351f
C55 VDD1.n26 VSUBS 0.036501f
C56 VDD1.n27 VSUBS 0.036501f
C57 VDD1.n28 VSUBS 0.016351f
C58 VDD1.n29 VSUBS 0.015443f
C59 VDD1.n30 VSUBS 0.028739f
C60 VDD1.n31 VSUBS 0.028739f
C61 VDD1.n32 VSUBS 0.015443f
C62 VDD1.n33 VSUBS 0.016351f
C63 VDD1.n34 VSUBS 0.036501f
C64 VDD1.n35 VSUBS 0.036501f
C65 VDD1.n36 VSUBS 0.016351f
C66 VDD1.n37 VSUBS 0.015443f
C67 VDD1.n38 VSUBS 0.028739f
C68 VDD1.n39 VSUBS 0.028739f
C69 VDD1.n40 VSUBS 0.015443f
C70 VDD1.n41 VSUBS 0.015897f
C71 VDD1.n42 VSUBS 0.015897f
C72 VDD1.n43 VSUBS 0.036501f
C73 VDD1.n44 VSUBS 0.036501f
C74 VDD1.n45 VSUBS 0.016351f
C75 VDD1.n46 VSUBS 0.015443f
C76 VDD1.n47 VSUBS 0.028739f
C77 VDD1.n48 VSUBS 0.028739f
C78 VDD1.n49 VSUBS 0.015443f
C79 VDD1.n50 VSUBS 0.016351f
C80 VDD1.n51 VSUBS 0.036501f
C81 VDD1.n52 VSUBS 0.083807f
C82 VDD1.n53 VSUBS 0.016351f
C83 VDD1.n54 VSUBS 0.015443f
C84 VDD1.n55 VSUBS 0.065643f
C85 VDD1.n56 VSUBS 0.076613f
C86 VDD1.n57 VSUBS 0.030239f
C87 VDD1.n58 VSUBS 0.028739f
C88 VDD1.n59 VSUBS 0.015443f
C89 VDD1.n60 VSUBS 0.036501f
C90 VDD1.n61 VSUBS 0.016351f
C91 VDD1.n62 VSUBS 0.028739f
C92 VDD1.n63 VSUBS 0.015443f
C93 VDD1.n64 VSUBS 0.036501f
C94 VDD1.n65 VSUBS 0.016351f
C95 VDD1.n66 VSUBS 0.028739f
C96 VDD1.n67 VSUBS 0.015443f
C97 VDD1.n68 VSUBS 0.036501f
C98 VDD1.n69 VSUBS 0.016351f
C99 VDD1.n70 VSUBS 0.028739f
C100 VDD1.n71 VSUBS 0.015443f
C101 VDD1.n72 VSUBS 0.036501f
C102 VDD1.n73 VSUBS 0.016351f
C103 VDD1.n74 VSUBS 0.208929f
C104 VDD1.t4 VSUBS 0.078535f
C105 VDD1.n75 VSUBS 0.027376f
C106 VDD1.n76 VSUBS 0.027458f
C107 VDD1.n77 VSUBS 0.015443f
C108 VDD1.n78 VSUBS 1.24327f
C109 VDD1.n79 VSUBS 0.028739f
C110 VDD1.n80 VSUBS 0.015443f
C111 VDD1.n81 VSUBS 0.016351f
C112 VDD1.n82 VSUBS 0.036501f
C113 VDD1.n83 VSUBS 0.036501f
C114 VDD1.n84 VSUBS 0.016351f
C115 VDD1.n85 VSUBS 0.015443f
C116 VDD1.n86 VSUBS 0.028739f
C117 VDD1.n87 VSUBS 0.028739f
C118 VDD1.n88 VSUBS 0.015443f
C119 VDD1.n89 VSUBS 0.016351f
C120 VDD1.n90 VSUBS 0.036501f
C121 VDD1.n91 VSUBS 0.036501f
C122 VDD1.n92 VSUBS 0.036501f
C123 VDD1.n93 VSUBS 0.016351f
C124 VDD1.n94 VSUBS 0.015443f
C125 VDD1.n95 VSUBS 0.028739f
C126 VDD1.n96 VSUBS 0.028739f
C127 VDD1.n97 VSUBS 0.015443f
C128 VDD1.n98 VSUBS 0.015897f
C129 VDD1.n99 VSUBS 0.015897f
C130 VDD1.n100 VSUBS 0.036501f
C131 VDD1.n101 VSUBS 0.036501f
C132 VDD1.n102 VSUBS 0.016351f
C133 VDD1.n103 VSUBS 0.015443f
C134 VDD1.n104 VSUBS 0.028739f
C135 VDD1.n105 VSUBS 0.028739f
C136 VDD1.n106 VSUBS 0.015443f
C137 VDD1.n107 VSUBS 0.016351f
C138 VDD1.n108 VSUBS 0.036501f
C139 VDD1.n109 VSUBS 0.083807f
C140 VDD1.n110 VSUBS 0.016351f
C141 VDD1.n111 VSUBS 0.015443f
C142 VDD1.n112 VSUBS 0.065643f
C143 VDD1.n113 VSUBS 0.075495f
C144 VDD1.t0 VSUBS 0.24209f
C145 VDD1.t5 VSUBS 0.24209f
C146 VDD1.n114 VSUBS 1.85774f
C147 VDD1.n115 VSUBS 3.92436f
C148 VDD1.t1 VSUBS 0.24209f
C149 VDD1.t3 VSUBS 0.24209f
C150 VDD1.n116 VSUBS 1.84822f
C151 VDD1.n117 VSUBS 3.69531f
C152 VP.t0 VSUBS 3.0808f
C153 VP.n0 VSUBS 1.19919f
C154 VP.n1 VSUBS 0.029819f
C155 VP.n2 VSUBS 0.047472f
C156 VP.n3 VSUBS 0.029819f
C157 VP.n4 VSUBS 0.041647f
C158 VP.n5 VSUBS 0.029819f
C159 VP.n6 VSUBS 0.039222f
C160 VP.n7 VSUBS 0.029819f
C161 VP.n8 VSUBS 0.036188f
C162 VP.t2 VSUBS 3.0808f
C163 VP.n9 VSUBS 1.19919f
C164 VP.n10 VSUBS 0.029819f
C165 VP.n11 VSUBS 0.047472f
C166 VP.n12 VSUBS 0.029819f
C167 VP.n13 VSUBS 0.041647f
C168 VP.t3 VSUBS 3.49287f
C169 VP.t4 VSUBS 3.0808f
C170 VP.n14 VSUBS 1.18985f
C171 VP.n15 VSUBS 1.1291f
C172 VP.n16 VSUBS 0.371991f
C173 VP.n17 VSUBS 0.029819f
C174 VP.n18 VSUBS 0.055297f
C175 VP.n19 VSUBS 0.055297f
C176 VP.n20 VSUBS 0.039222f
C177 VP.n21 VSUBS 0.029819f
C178 VP.n22 VSUBS 0.029819f
C179 VP.n23 VSUBS 0.029819f
C180 VP.n24 VSUBS 0.055297f
C181 VP.n25 VSUBS 0.055297f
C182 VP.n26 VSUBS 0.036188f
C183 VP.n27 VSUBS 0.04812f
C184 VP.n28 VSUBS 1.78222f
C185 VP.t1 VSUBS 3.0808f
C186 VP.n29 VSUBS 1.19919f
C187 VP.n30 VSUBS 1.80309f
C188 VP.n31 VSUBS 0.04812f
C189 VP.n32 VSUBS 0.029819f
C190 VP.n33 VSUBS 0.055297f
C191 VP.n34 VSUBS 0.055297f
C192 VP.n35 VSUBS 0.047472f
C193 VP.n36 VSUBS 0.029819f
C194 VP.n37 VSUBS 0.029819f
C195 VP.n38 VSUBS 0.029819f
C196 VP.n39 VSUBS 0.055297f
C197 VP.n40 VSUBS 0.055297f
C198 VP.t5 VSUBS 3.0808f
C199 VP.n41 VSUBS 1.08738f
C200 VP.n42 VSUBS 0.041647f
C201 VP.n43 VSUBS 0.029819f
C202 VP.n44 VSUBS 0.029819f
C203 VP.n45 VSUBS 0.029819f
C204 VP.n46 VSUBS 0.055297f
C205 VP.n47 VSUBS 0.055297f
C206 VP.n48 VSUBS 0.039222f
C207 VP.n49 VSUBS 0.029819f
C208 VP.n50 VSUBS 0.029819f
C209 VP.n51 VSUBS 0.029819f
C210 VP.n52 VSUBS 0.055297f
C211 VP.n53 VSUBS 0.055297f
C212 VP.n54 VSUBS 0.036188f
C213 VP.n55 VSUBS 0.04812f
C214 VP.n56 VSUBS 0.083715f
C215 VTAIL.t10 VSUBS 0.257317f
C216 VTAIL.t11 VSUBS 0.257317f
C217 VTAIL.n0 VSUBS 1.8068f
C218 VTAIL.n1 VSUBS 0.977982f
C219 VTAIL.n2 VSUBS 0.032141f
C220 VTAIL.n3 VSUBS 0.030546f
C221 VTAIL.n4 VSUBS 0.016414f
C222 VTAIL.n5 VSUBS 0.038797f
C223 VTAIL.n6 VSUBS 0.01738f
C224 VTAIL.n7 VSUBS 0.030546f
C225 VTAIL.n8 VSUBS 0.016414f
C226 VTAIL.n9 VSUBS 0.038797f
C227 VTAIL.n10 VSUBS 0.01738f
C228 VTAIL.n11 VSUBS 0.030546f
C229 VTAIL.n12 VSUBS 0.016414f
C230 VTAIL.n13 VSUBS 0.038797f
C231 VTAIL.n14 VSUBS 0.01738f
C232 VTAIL.n15 VSUBS 0.030546f
C233 VTAIL.n16 VSUBS 0.016414f
C234 VTAIL.n17 VSUBS 0.038797f
C235 VTAIL.n18 VSUBS 0.01738f
C236 VTAIL.n19 VSUBS 0.22207f
C237 VTAIL.t0 VSUBS 0.083475f
C238 VTAIL.n20 VSUBS 0.029098f
C239 VTAIL.n21 VSUBS 0.029185f
C240 VTAIL.n22 VSUBS 0.016414f
C241 VTAIL.n23 VSUBS 1.32147f
C242 VTAIL.n24 VSUBS 0.030546f
C243 VTAIL.n25 VSUBS 0.016414f
C244 VTAIL.n26 VSUBS 0.01738f
C245 VTAIL.n27 VSUBS 0.038797f
C246 VTAIL.n28 VSUBS 0.038797f
C247 VTAIL.n29 VSUBS 0.01738f
C248 VTAIL.n30 VSUBS 0.016414f
C249 VTAIL.n31 VSUBS 0.030546f
C250 VTAIL.n32 VSUBS 0.030546f
C251 VTAIL.n33 VSUBS 0.016414f
C252 VTAIL.n34 VSUBS 0.01738f
C253 VTAIL.n35 VSUBS 0.038797f
C254 VTAIL.n36 VSUBS 0.038797f
C255 VTAIL.n37 VSUBS 0.038797f
C256 VTAIL.n38 VSUBS 0.01738f
C257 VTAIL.n39 VSUBS 0.016414f
C258 VTAIL.n40 VSUBS 0.030546f
C259 VTAIL.n41 VSUBS 0.030546f
C260 VTAIL.n42 VSUBS 0.016414f
C261 VTAIL.n43 VSUBS 0.016897f
C262 VTAIL.n44 VSUBS 0.016897f
C263 VTAIL.n45 VSUBS 0.038797f
C264 VTAIL.n46 VSUBS 0.038797f
C265 VTAIL.n47 VSUBS 0.01738f
C266 VTAIL.n48 VSUBS 0.016414f
C267 VTAIL.n49 VSUBS 0.030546f
C268 VTAIL.n50 VSUBS 0.030546f
C269 VTAIL.n51 VSUBS 0.016414f
C270 VTAIL.n52 VSUBS 0.01738f
C271 VTAIL.n53 VSUBS 0.038797f
C272 VTAIL.n54 VSUBS 0.089078f
C273 VTAIL.n55 VSUBS 0.01738f
C274 VTAIL.n56 VSUBS 0.016414f
C275 VTAIL.n57 VSUBS 0.069772f
C276 VTAIL.n58 VSUBS 0.044556f
C277 VTAIL.n59 VSUBS 0.568238f
C278 VTAIL.t5 VSUBS 0.257317f
C279 VTAIL.t3 VSUBS 0.257317f
C280 VTAIL.n60 VSUBS 1.8068f
C281 VTAIL.n61 VSUBS 2.99002f
C282 VTAIL.t6 VSUBS 0.257317f
C283 VTAIL.t8 VSUBS 0.257317f
C284 VTAIL.n62 VSUBS 1.80681f
C285 VTAIL.n63 VSUBS 2.99001f
C286 VTAIL.n64 VSUBS 0.032141f
C287 VTAIL.n65 VSUBS 0.030546f
C288 VTAIL.n66 VSUBS 0.016414f
C289 VTAIL.n67 VSUBS 0.038797f
C290 VTAIL.n68 VSUBS 0.01738f
C291 VTAIL.n69 VSUBS 0.030546f
C292 VTAIL.n70 VSUBS 0.016414f
C293 VTAIL.n71 VSUBS 0.038797f
C294 VTAIL.n72 VSUBS 0.01738f
C295 VTAIL.n73 VSUBS 0.030546f
C296 VTAIL.n74 VSUBS 0.016414f
C297 VTAIL.n75 VSUBS 0.038797f
C298 VTAIL.n76 VSUBS 0.038797f
C299 VTAIL.n77 VSUBS 0.01738f
C300 VTAIL.n78 VSUBS 0.030546f
C301 VTAIL.n79 VSUBS 0.016414f
C302 VTAIL.n80 VSUBS 0.038797f
C303 VTAIL.n81 VSUBS 0.01738f
C304 VTAIL.n82 VSUBS 0.22207f
C305 VTAIL.t9 VSUBS 0.083475f
C306 VTAIL.n83 VSUBS 0.029098f
C307 VTAIL.n84 VSUBS 0.029185f
C308 VTAIL.n85 VSUBS 0.016414f
C309 VTAIL.n86 VSUBS 1.32147f
C310 VTAIL.n87 VSUBS 0.030546f
C311 VTAIL.n88 VSUBS 0.016414f
C312 VTAIL.n89 VSUBS 0.01738f
C313 VTAIL.n90 VSUBS 0.038797f
C314 VTAIL.n91 VSUBS 0.038797f
C315 VTAIL.n92 VSUBS 0.01738f
C316 VTAIL.n93 VSUBS 0.016414f
C317 VTAIL.n94 VSUBS 0.030546f
C318 VTAIL.n95 VSUBS 0.030546f
C319 VTAIL.n96 VSUBS 0.016414f
C320 VTAIL.n97 VSUBS 0.01738f
C321 VTAIL.n98 VSUBS 0.038797f
C322 VTAIL.n99 VSUBS 0.038797f
C323 VTAIL.n100 VSUBS 0.01738f
C324 VTAIL.n101 VSUBS 0.016414f
C325 VTAIL.n102 VSUBS 0.030546f
C326 VTAIL.n103 VSUBS 0.030546f
C327 VTAIL.n104 VSUBS 0.016414f
C328 VTAIL.n105 VSUBS 0.016897f
C329 VTAIL.n106 VSUBS 0.016897f
C330 VTAIL.n107 VSUBS 0.038797f
C331 VTAIL.n108 VSUBS 0.038797f
C332 VTAIL.n109 VSUBS 0.01738f
C333 VTAIL.n110 VSUBS 0.016414f
C334 VTAIL.n111 VSUBS 0.030546f
C335 VTAIL.n112 VSUBS 0.030546f
C336 VTAIL.n113 VSUBS 0.016414f
C337 VTAIL.n114 VSUBS 0.01738f
C338 VTAIL.n115 VSUBS 0.038797f
C339 VTAIL.n116 VSUBS 0.089078f
C340 VTAIL.n117 VSUBS 0.01738f
C341 VTAIL.n118 VSUBS 0.016414f
C342 VTAIL.n119 VSUBS 0.069772f
C343 VTAIL.n120 VSUBS 0.044556f
C344 VTAIL.n121 VSUBS 0.568238f
C345 VTAIL.t1 VSUBS 0.257317f
C346 VTAIL.t2 VSUBS 0.257317f
C347 VTAIL.n122 VSUBS 1.80681f
C348 VTAIL.n123 VSUBS 1.22043f
C349 VTAIL.n124 VSUBS 0.032141f
C350 VTAIL.n125 VSUBS 0.030546f
C351 VTAIL.n126 VSUBS 0.016414f
C352 VTAIL.n127 VSUBS 0.038797f
C353 VTAIL.n128 VSUBS 0.01738f
C354 VTAIL.n129 VSUBS 0.030546f
C355 VTAIL.n130 VSUBS 0.016414f
C356 VTAIL.n131 VSUBS 0.038797f
C357 VTAIL.n132 VSUBS 0.01738f
C358 VTAIL.n133 VSUBS 0.030546f
C359 VTAIL.n134 VSUBS 0.016414f
C360 VTAIL.n135 VSUBS 0.038797f
C361 VTAIL.n136 VSUBS 0.038797f
C362 VTAIL.n137 VSUBS 0.01738f
C363 VTAIL.n138 VSUBS 0.030546f
C364 VTAIL.n139 VSUBS 0.016414f
C365 VTAIL.n140 VSUBS 0.038797f
C366 VTAIL.n141 VSUBS 0.01738f
C367 VTAIL.n142 VSUBS 0.22207f
C368 VTAIL.t4 VSUBS 0.083475f
C369 VTAIL.n143 VSUBS 0.029098f
C370 VTAIL.n144 VSUBS 0.029185f
C371 VTAIL.n145 VSUBS 0.016414f
C372 VTAIL.n146 VSUBS 1.32147f
C373 VTAIL.n147 VSUBS 0.030546f
C374 VTAIL.n148 VSUBS 0.016414f
C375 VTAIL.n149 VSUBS 0.01738f
C376 VTAIL.n150 VSUBS 0.038797f
C377 VTAIL.n151 VSUBS 0.038797f
C378 VTAIL.n152 VSUBS 0.01738f
C379 VTAIL.n153 VSUBS 0.016414f
C380 VTAIL.n154 VSUBS 0.030546f
C381 VTAIL.n155 VSUBS 0.030546f
C382 VTAIL.n156 VSUBS 0.016414f
C383 VTAIL.n157 VSUBS 0.01738f
C384 VTAIL.n158 VSUBS 0.038797f
C385 VTAIL.n159 VSUBS 0.038797f
C386 VTAIL.n160 VSUBS 0.01738f
C387 VTAIL.n161 VSUBS 0.016414f
C388 VTAIL.n162 VSUBS 0.030546f
C389 VTAIL.n163 VSUBS 0.030546f
C390 VTAIL.n164 VSUBS 0.016414f
C391 VTAIL.n165 VSUBS 0.016897f
C392 VTAIL.n166 VSUBS 0.016897f
C393 VTAIL.n167 VSUBS 0.038797f
C394 VTAIL.n168 VSUBS 0.038797f
C395 VTAIL.n169 VSUBS 0.01738f
C396 VTAIL.n170 VSUBS 0.016414f
C397 VTAIL.n171 VSUBS 0.030546f
C398 VTAIL.n172 VSUBS 0.030546f
C399 VTAIL.n173 VSUBS 0.016414f
C400 VTAIL.n174 VSUBS 0.01738f
C401 VTAIL.n175 VSUBS 0.038797f
C402 VTAIL.n176 VSUBS 0.089078f
C403 VTAIL.n177 VSUBS 0.01738f
C404 VTAIL.n178 VSUBS 0.016414f
C405 VTAIL.n179 VSUBS 0.069772f
C406 VTAIL.n180 VSUBS 0.044556f
C407 VTAIL.n181 VSUBS 2.0069f
C408 VTAIL.n182 VSUBS 0.032141f
C409 VTAIL.n183 VSUBS 0.030546f
C410 VTAIL.n184 VSUBS 0.016414f
C411 VTAIL.n185 VSUBS 0.038797f
C412 VTAIL.n186 VSUBS 0.01738f
C413 VTAIL.n187 VSUBS 0.030546f
C414 VTAIL.n188 VSUBS 0.016414f
C415 VTAIL.n189 VSUBS 0.038797f
C416 VTAIL.n190 VSUBS 0.01738f
C417 VTAIL.n191 VSUBS 0.030546f
C418 VTAIL.n192 VSUBS 0.016414f
C419 VTAIL.n193 VSUBS 0.038797f
C420 VTAIL.n194 VSUBS 0.01738f
C421 VTAIL.n195 VSUBS 0.030546f
C422 VTAIL.n196 VSUBS 0.016414f
C423 VTAIL.n197 VSUBS 0.038797f
C424 VTAIL.n198 VSUBS 0.01738f
C425 VTAIL.n199 VSUBS 0.22207f
C426 VTAIL.t7 VSUBS 0.083475f
C427 VTAIL.n200 VSUBS 0.029098f
C428 VTAIL.n201 VSUBS 0.029185f
C429 VTAIL.n202 VSUBS 0.016414f
C430 VTAIL.n203 VSUBS 1.32147f
C431 VTAIL.n204 VSUBS 0.030546f
C432 VTAIL.n205 VSUBS 0.016414f
C433 VTAIL.n206 VSUBS 0.01738f
C434 VTAIL.n207 VSUBS 0.038797f
C435 VTAIL.n208 VSUBS 0.038797f
C436 VTAIL.n209 VSUBS 0.01738f
C437 VTAIL.n210 VSUBS 0.016414f
C438 VTAIL.n211 VSUBS 0.030546f
C439 VTAIL.n212 VSUBS 0.030546f
C440 VTAIL.n213 VSUBS 0.016414f
C441 VTAIL.n214 VSUBS 0.01738f
C442 VTAIL.n215 VSUBS 0.038797f
C443 VTAIL.n216 VSUBS 0.038797f
C444 VTAIL.n217 VSUBS 0.038797f
C445 VTAIL.n218 VSUBS 0.01738f
C446 VTAIL.n219 VSUBS 0.016414f
C447 VTAIL.n220 VSUBS 0.030546f
C448 VTAIL.n221 VSUBS 0.030546f
C449 VTAIL.n222 VSUBS 0.016414f
C450 VTAIL.n223 VSUBS 0.016897f
C451 VTAIL.n224 VSUBS 0.016897f
C452 VTAIL.n225 VSUBS 0.038797f
C453 VTAIL.n226 VSUBS 0.038797f
C454 VTAIL.n227 VSUBS 0.01738f
C455 VTAIL.n228 VSUBS 0.016414f
C456 VTAIL.n229 VSUBS 0.030546f
C457 VTAIL.n230 VSUBS 0.030546f
C458 VTAIL.n231 VSUBS 0.016414f
C459 VTAIL.n232 VSUBS 0.01738f
C460 VTAIL.n233 VSUBS 0.038797f
C461 VTAIL.n234 VSUBS 0.089078f
C462 VTAIL.n235 VSUBS 0.01738f
C463 VTAIL.n236 VSUBS 0.016414f
C464 VTAIL.n237 VSUBS 0.069772f
C465 VTAIL.n238 VSUBS 0.044556f
C466 VTAIL.n239 VSUBS 1.91844f
C467 VDD2.n0 VSUBS 0.03041f
C468 VDD2.n1 VSUBS 0.028901f
C469 VDD2.n2 VSUBS 0.01553f
C470 VDD2.n3 VSUBS 0.036708f
C471 VDD2.n4 VSUBS 0.016444f
C472 VDD2.n5 VSUBS 0.028901f
C473 VDD2.n6 VSUBS 0.01553f
C474 VDD2.n7 VSUBS 0.036708f
C475 VDD2.n8 VSUBS 0.016444f
C476 VDD2.n9 VSUBS 0.028901f
C477 VDD2.n10 VSUBS 0.01553f
C478 VDD2.n11 VSUBS 0.036708f
C479 VDD2.n12 VSUBS 0.016444f
C480 VDD2.n13 VSUBS 0.028901f
C481 VDD2.n14 VSUBS 0.01553f
C482 VDD2.n15 VSUBS 0.036708f
C483 VDD2.n16 VSUBS 0.016444f
C484 VDD2.n17 VSUBS 0.210109f
C485 VDD2.t3 VSUBS 0.078979f
C486 VDD2.n18 VSUBS 0.027531f
C487 VDD2.n19 VSUBS 0.027613f
C488 VDD2.n20 VSUBS 0.01553f
C489 VDD2.n21 VSUBS 1.25029f
C490 VDD2.n22 VSUBS 0.028901f
C491 VDD2.n23 VSUBS 0.01553f
C492 VDD2.n24 VSUBS 0.016444f
C493 VDD2.n25 VSUBS 0.036708f
C494 VDD2.n26 VSUBS 0.036708f
C495 VDD2.n27 VSUBS 0.016444f
C496 VDD2.n28 VSUBS 0.01553f
C497 VDD2.n29 VSUBS 0.028901f
C498 VDD2.n30 VSUBS 0.028901f
C499 VDD2.n31 VSUBS 0.01553f
C500 VDD2.n32 VSUBS 0.016444f
C501 VDD2.n33 VSUBS 0.036708f
C502 VDD2.n34 VSUBS 0.036708f
C503 VDD2.n35 VSUBS 0.036708f
C504 VDD2.n36 VSUBS 0.016444f
C505 VDD2.n37 VSUBS 0.01553f
C506 VDD2.n38 VSUBS 0.028901f
C507 VDD2.n39 VSUBS 0.028901f
C508 VDD2.n40 VSUBS 0.01553f
C509 VDD2.n41 VSUBS 0.015987f
C510 VDD2.n42 VSUBS 0.015987f
C511 VDD2.n43 VSUBS 0.036708f
C512 VDD2.n44 VSUBS 0.036708f
C513 VDD2.n45 VSUBS 0.016444f
C514 VDD2.n46 VSUBS 0.01553f
C515 VDD2.n47 VSUBS 0.028901f
C516 VDD2.n48 VSUBS 0.028901f
C517 VDD2.n49 VSUBS 0.01553f
C518 VDD2.n50 VSUBS 0.016444f
C519 VDD2.n51 VSUBS 0.036708f
C520 VDD2.n52 VSUBS 0.08428f
C521 VDD2.n53 VSUBS 0.016444f
C522 VDD2.n54 VSUBS 0.01553f
C523 VDD2.n55 VSUBS 0.066014f
C524 VDD2.n56 VSUBS 0.075922f
C525 VDD2.t1 VSUBS 0.243458f
C526 VDD2.t4 VSUBS 0.243458f
C527 VDD2.n57 VSUBS 1.86824f
C528 VDD2.n58 VSUBS 3.77468f
C529 VDD2.n59 VSUBS 0.03041f
C530 VDD2.n60 VSUBS 0.028901f
C531 VDD2.n61 VSUBS 0.01553f
C532 VDD2.n62 VSUBS 0.036708f
C533 VDD2.n63 VSUBS 0.016444f
C534 VDD2.n64 VSUBS 0.028901f
C535 VDD2.n65 VSUBS 0.01553f
C536 VDD2.n66 VSUBS 0.036708f
C537 VDD2.n67 VSUBS 0.016444f
C538 VDD2.n68 VSUBS 0.028901f
C539 VDD2.n69 VSUBS 0.01553f
C540 VDD2.n70 VSUBS 0.036708f
C541 VDD2.n71 VSUBS 0.036708f
C542 VDD2.n72 VSUBS 0.016444f
C543 VDD2.n73 VSUBS 0.028901f
C544 VDD2.n74 VSUBS 0.01553f
C545 VDD2.n75 VSUBS 0.036708f
C546 VDD2.n76 VSUBS 0.016444f
C547 VDD2.n77 VSUBS 0.210109f
C548 VDD2.t0 VSUBS 0.078979f
C549 VDD2.n78 VSUBS 0.027531f
C550 VDD2.n79 VSUBS 0.027613f
C551 VDD2.n80 VSUBS 0.01553f
C552 VDD2.n81 VSUBS 1.25029f
C553 VDD2.n82 VSUBS 0.028901f
C554 VDD2.n83 VSUBS 0.01553f
C555 VDD2.n84 VSUBS 0.016444f
C556 VDD2.n85 VSUBS 0.036708f
C557 VDD2.n86 VSUBS 0.036708f
C558 VDD2.n87 VSUBS 0.016444f
C559 VDD2.n88 VSUBS 0.01553f
C560 VDD2.n89 VSUBS 0.028901f
C561 VDD2.n90 VSUBS 0.028901f
C562 VDD2.n91 VSUBS 0.01553f
C563 VDD2.n92 VSUBS 0.016444f
C564 VDD2.n93 VSUBS 0.036708f
C565 VDD2.n94 VSUBS 0.036708f
C566 VDD2.n95 VSUBS 0.016444f
C567 VDD2.n96 VSUBS 0.01553f
C568 VDD2.n97 VSUBS 0.028901f
C569 VDD2.n98 VSUBS 0.028901f
C570 VDD2.n99 VSUBS 0.01553f
C571 VDD2.n100 VSUBS 0.015987f
C572 VDD2.n101 VSUBS 0.015987f
C573 VDD2.n102 VSUBS 0.036708f
C574 VDD2.n103 VSUBS 0.036708f
C575 VDD2.n104 VSUBS 0.016444f
C576 VDD2.n105 VSUBS 0.01553f
C577 VDD2.n106 VSUBS 0.028901f
C578 VDD2.n107 VSUBS 0.028901f
C579 VDD2.n108 VSUBS 0.01553f
C580 VDD2.n109 VSUBS 0.016444f
C581 VDD2.n110 VSUBS 0.036708f
C582 VDD2.n111 VSUBS 0.08428f
C583 VDD2.n112 VSUBS 0.016444f
C584 VDD2.n113 VSUBS 0.01553f
C585 VDD2.n114 VSUBS 0.066014f
C586 VDD2.n115 VSUBS 0.062118f
C587 VDD2.n116 VSUBS 3.14771f
C588 VDD2.t5 VSUBS 0.243458f
C589 VDD2.t2 VSUBS 0.243458f
C590 VDD2.n117 VSUBS 1.86819f
C591 VN.t4 VSUBS 2.75847f
C592 VN.n0 VSUBS 1.07373f
C593 VN.n1 VSUBS 0.026699f
C594 VN.n2 VSUBS 0.042505f
C595 VN.n3 VSUBS 0.026699f
C596 VN.n4 VSUBS 0.03729f
C597 VN.t0 VSUBS 2.75847f
C598 VN.n5 VSUBS 1.06536f
C599 VN.t1 VSUBS 3.12744f
C600 VN.n6 VSUBS 1.01096f
C601 VN.n7 VSUBS 0.333071f
C602 VN.n8 VSUBS 0.026699f
C603 VN.n9 VSUBS 0.049511f
C604 VN.n10 VSUBS 0.049511f
C605 VN.n11 VSUBS 0.035118f
C606 VN.n12 VSUBS 0.026699f
C607 VN.n13 VSUBS 0.026699f
C608 VN.n14 VSUBS 0.026699f
C609 VN.n15 VSUBS 0.049511f
C610 VN.n16 VSUBS 0.049511f
C611 VN.n17 VSUBS 0.032402f
C612 VN.n18 VSUBS 0.043085f
C613 VN.n19 VSUBS 0.074956f
C614 VN.t5 VSUBS 2.75847f
C615 VN.n20 VSUBS 1.07373f
C616 VN.n21 VSUBS 0.026699f
C617 VN.n22 VSUBS 0.042505f
C618 VN.n23 VSUBS 0.026699f
C619 VN.n24 VSUBS 0.03729f
C620 VN.t2 VSUBS 3.12744f
C621 VN.t3 VSUBS 2.75847f
C622 VN.n25 VSUBS 1.06536f
C623 VN.n26 VSUBS 1.01096f
C624 VN.n27 VSUBS 0.333071f
C625 VN.n28 VSUBS 0.026699f
C626 VN.n29 VSUBS 0.049511f
C627 VN.n30 VSUBS 0.049511f
C628 VN.n31 VSUBS 0.035118f
C629 VN.n32 VSUBS 0.026699f
C630 VN.n33 VSUBS 0.026699f
C631 VN.n34 VSUBS 0.026699f
C632 VN.n35 VSUBS 0.049511f
C633 VN.n36 VSUBS 0.049511f
C634 VN.n37 VSUBS 0.032402f
C635 VN.n38 VSUBS 0.043085f
C636 VN.n39 VSUBS 1.60657f
C637 B.n0 VSUBS 0.005578f
C638 B.n1 VSUBS 0.005578f
C639 B.n2 VSUBS 0.008821f
C640 B.n3 VSUBS 0.008821f
C641 B.n4 VSUBS 0.008821f
C642 B.n5 VSUBS 0.008821f
C643 B.n6 VSUBS 0.008821f
C644 B.n7 VSUBS 0.008821f
C645 B.n8 VSUBS 0.008821f
C646 B.n9 VSUBS 0.008821f
C647 B.n10 VSUBS 0.008821f
C648 B.n11 VSUBS 0.008821f
C649 B.n12 VSUBS 0.008821f
C650 B.n13 VSUBS 0.008821f
C651 B.n14 VSUBS 0.008821f
C652 B.n15 VSUBS 0.008821f
C653 B.n16 VSUBS 0.008821f
C654 B.n17 VSUBS 0.008821f
C655 B.n18 VSUBS 0.008821f
C656 B.n19 VSUBS 0.008821f
C657 B.n20 VSUBS 0.008821f
C658 B.n21 VSUBS 0.008821f
C659 B.n22 VSUBS 0.008821f
C660 B.n23 VSUBS 0.008821f
C661 B.n24 VSUBS 0.008821f
C662 B.n25 VSUBS 0.008821f
C663 B.n26 VSUBS 0.008821f
C664 B.n27 VSUBS 0.008821f
C665 B.n28 VSUBS 0.008821f
C666 B.n29 VSUBS 0.020897f
C667 B.n30 VSUBS 0.008821f
C668 B.n31 VSUBS 0.008821f
C669 B.n32 VSUBS 0.008821f
C670 B.n33 VSUBS 0.008821f
C671 B.n34 VSUBS 0.008821f
C672 B.n35 VSUBS 0.008821f
C673 B.n36 VSUBS 0.008821f
C674 B.n37 VSUBS 0.008821f
C675 B.n38 VSUBS 0.008821f
C676 B.n39 VSUBS 0.008821f
C677 B.n40 VSUBS 0.008821f
C678 B.n41 VSUBS 0.008821f
C679 B.n42 VSUBS 0.008821f
C680 B.n43 VSUBS 0.008821f
C681 B.n44 VSUBS 0.008821f
C682 B.n45 VSUBS 0.008821f
C683 B.n46 VSUBS 0.008821f
C684 B.n47 VSUBS 0.008821f
C685 B.t2 VSUBS 0.228784f
C686 B.t1 VSUBS 0.279419f
C687 B.t0 VSUBS 2.2424f
C688 B.n48 VSUBS 0.448531f
C689 B.n49 VSUBS 0.298481f
C690 B.n50 VSUBS 0.020437f
C691 B.n51 VSUBS 0.008821f
C692 B.n52 VSUBS 0.008821f
C693 B.n53 VSUBS 0.008821f
C694 B.n54 VSUBS 0.008821f
C695 B.n55 VSUBS 0.008821f
C696 B.t5 VSUBS 0.228787f
C697 B.t4 VSUBS 0.279422f
C698 B.t3 VSUBS 2.2424f
C699 B.n56 VSUBS 0.448528f
C700 B.n57 VSUBS 0.298478f
C701 B.n58 VSUBS 0.008821f
C702 B.n59 VSUBS 0.008821f
C703 B.n60 VSUBS 0.008821f
C704 B.n61 VSUBS 0.008821f
C705 B.n62 VSUBS 0.008821f
C706 B.n63 VSUBS 0.008821f
C707 B.n64 VSUBS 0.008821f
C708 B.n65 VSUBS 0.008821f
C709 B.n66 VSUBS 0.008821f
C710 B.n67 VSUBS 0.008821f
C711 B.n68 VSUBS 0.008821f
C712 B.n69 VSUBS 0.008821f
C713 B.n70 VSUBS 0.008821f
C714 B.n71 VSUBS 0.008821f
C715 B.n72 VSUBS 0.008821f
C716 B.n73 VSUBS 0.008821f
C717 B.n74 VSUBS 0.008821f
C718 B.n75 VSUBS 0.008821f
C719 B.n76 VSUBS 0.020897f
C720 B.n77 VSUBS 0.008821f
C721 B.n78 VSUBS 0.008821f
C722 B.n79 VSUBS 0.008821f
C723 B.n80 VSUBS 0.008821f
C724 B.n81 VSUBS 0.008821f
C725 B.n82 VSUBS 0.008821f
C726 B.n83 VSUBS 0.008821f
C727 B.n84 VSUBS 0.008821f
C728 B.n85 VSUBS 0.008821f
C729 B.n86 VSUBS 0.008821f
C730 B.n87 VSUBS 0.008821f
C731 B.n88 VSUBS 0.008821f
C732 B.n89 VSUBS 0.008821f
C733 B.n90 VSUBS 0.008821f
C734 B.n91 VSUBS 0.008821f
C735 B.n92 VSUBS 0.008821f
C736 B.n93 VSUBS 0.008821f
C737 B.n94 VSUBS 0.008821f
C738 B.n95 VSUBS 0.008821f
C739 B.n96 VSUBS 0.008821f
C740 B.n97 VSUBS 0.008821f
C741 B.n98 VSUBS 0.008821f
C742 B.n99 VSUBS 0.008821f
C743 B.n100 VSUBS 0.008821f
C744 B.n101 VSUBS 0.008821f
C745 B.n102 VSUBS 0.008821f
C746 B.n103 VSUBS 0.008821f
C747 B.n104 VSUBS 0.008821f
C748 B.n105 VSUBS 0.008821f
C749 B.n106 VSUBS 0.008821f
C750 B.n107 VSUBS 0.008821f
C751 B.n108 VSUBS 0.008821f
C752 B.n109 VSUBS 0.008821f
C753 B.n110 VSUBS 0.008821f
C754 B.n111 VSUBS 0.008821f
C755 B.n112 VSUBS 0.008821f
C756 B.n113 VSUBS 0.008821f
C757 B.n114 VSUBS 0.008821f
C758 B.n115 VSUBS 0.008821f
C759 B.n116 VSUBS 0.008821f
C760 B.n117 VSUBS 0.008821f
C761 B.n118 VSUBS 0.008821f
C762 B.n119 VSUBS 0.008821f
C763 B.n120 VSUBS 0.008821f
C764 B.n121 VSUBS 0.008821f
C765 B.n122 VSUBS 0.008821f
C766 B.n123 VSUBS 0.008821f
C767 B.n124 VSUBS 0.008821f
C768 B.n125 VSUBS 0.008821f
C769 B.n126 VSUBS 0.008821f
C770 B.n127 VSUBS 0.008821f
C771 B.n128 VSUBS 0.008821f
C772 B.n129 VSUBS 0.008821f
C773 B.n130 VSUBS 0.019834f
C774 B.n131 VSUBS 0.008821f
C775 B.n132 VSUBS 0.008821f
C776 B.n133 VSUBS 0.008821f
C777 B.n134 VSUBS 0.008821f
C778 B.n135 VSUBS 0.008821f
C779 B.n136 VSUBS 0.008821f
C780 B.n137 VSUBS 0.008821f
C781 B.n138 VSUBS 0.008821f
C782 B.n139 VSUBS 0.008821f
C783 B.n140 VSUBS 0.008821f
C784 B.n141 VSUBS 0.008821f
C785 B.n142 VSUBS 0.008821f
C786 B.n143 VSUBS 0.008821f
C787 B.n144 VSUBS 0.008821f
C788 B.n145 VSUBS 0.008821f
C789 B.n146 VSUBS 0.008821f
C790 B.n147 VSUBS 0.008821f
C791 B.n148 VSUBS 0.008821f
C792 B.n149 VSUBS 0.008821f
C793 B.t10 VSUBS 0.228787f
C794 B.t11 VSUBS 0.279422f
C795 B.t9 VSUBS 2.2424f
C796 B.n150 VSUBS 0.448528f
C797 B.n151 VSUBS 0.298478f
C798 B.n152 VSUBS 0.008821f
C799 B.n153 VSUBS 0.008821f
C800 B.n154 VSUBS 0.008821f
C801 B.n155 VSUBS 0.008821f
C802 B.t7 VSUBS 0.228784f
C803 B.t8 VSUBS 0.279419f
C804 B.t6 VSUBS 2.2424f
C805 B.n156 VSUBS 0.448531f
C806 B.n157 VSUBS 0.298481f
C807 B.n158 VSUBS 0.020437f
C808 B.n159 VSUBS 0.008821f
C809 B.n160 VSUBS 0.008821f
C810 B.n161 VSUBS 0.008821f
C811 B.n162 VSUBS 0.008821f
C812 B.n163 VSUBS 0.008821f
C813 B.n164 VSUBS 0.008821f
C814 B.n165 VSUBS 0.008821f
C815 B.n166 VSUBS 0.008821f
C816 B.n167 VSUBS 0.008821f
C817 B.n168 VSUBS 0.008821f
C818 B.n169 VSUBS 0.008821f
C819 B.n170 VSUBS 0.008821f
C820 B.n171 VSUBS 0.008821f
C821 B.n172 VSUBS 0.008821f
C822 B.n173 VSUBS 0.008821f
C823 B.n174 VSUBS 0.008821f
C824 B.n175 VSUBS 0.008821f
C825 B.n176 VSUBS 0.008821f
C826 B.n177 VSUBS 0.020897f
C827 B.n178 VSUBS 0.008821f
C828 B.n179 VSUBS 0.008821f
C829 B.n180 VSUBS 0.008821f
C830 B.n181 VSUBS 0.008821f
C831 B.n182 VSUBS 0.008821f
C832 B.n183 VSUBS 0.008821f
C833 B.n184 VSUBS 0.008821f
C834 B.n185 VSUBS 0.008821f
C835 B.n186 VSUBS 0.008821f
C836 B.n187 VSUBS 0.008821f
C837 B.n188 VSUBS 0.008821f
C838 B.n189 VSUBS 0.008821f
C839 B.n190 VSUBS 0.008821f
C840 B.n191 VSUBS 0.008821f
C841 B.n192 VSUBS 0.008821f
C842 B.n193 VSUBS 0.008821f
C843 B.n194 VSUBS 0.008821f
C844 B.n195 VSUBS 0.008821f
C845 B.n196 VSUBS 0.008821f
C846 B.n197 VSUBS 0.008821f
C847 B.n198 VSUBS 0.008821f
C848 B.n199 VSUBS 0.008821f
C849 B.n200 VSUBS 0.008821f
C850 B.n201 VSUBS 0.008821f
C851 B.n202 VSUBS 0.008821f
C852 B.n203 VSUBS 0.008821f
C853 B.n204 VSUBS 0.008821f
C854 B.n205 VSUBS 0.008821f
C855 B.n206 VSUBS 0.008821f
C856 B.n207 VSUBS 0.008821f
C857 B.n208 VSUBS 0.008821f
C858 B.n209 VSUBS 0.008821f
C859 B.n210 VSUBS 0.008821f
C860 B.n211 VSUBS 0.008821f
C861 B.n212 VSUBS 0.008821f
C862 B.n213 VSUBS 0.008821f
C863 B.n214 VSUBS 0.008821f
C864 B.n215 VSUBS 0.008821f
C865 B.n216 VSUBS 0.008821f
C866 B.n217 VSUBS 0.008821f
C867 B.n218 VSUBS 0.008821f
C868 B.n219 VSUBS 0.008821f
C869 B.n220 VSUBS 0.008821f
C870 B.n221 VSUBS 0.008821f
C871 B.n222 VSUBS 0.008821f
C872 B.n223 VSUBS 0.008821f
C873 B.n224 VSUBS 0.008821f
C874 B.n225 VSUBS 0.008821f
C875 B.n226 VSUBS 0.008821f
C876 B.n227 VSUBS 0.008821f
C877 B.n228 VSUBS 0.008821f
C878 B.n229 VSUBS 0.008821f
C879 B.n230 VSUBS 0.008821f
C880 B.n231 VSUBS 0.008821f
C881 B.n232 VSUBS 0.008821f
C882 B.n233 VSUBS 0.008821f
C883 B.n234 VSUBS 0.008821f
C884 B.n235 VSUBS 0.008821f
C885 B.n236 VSUBS 0.008821f
C886 B.n237 VSUBS 0.008821f
C887 B.n238 VSUBS 0.008821f
C888 B.n239 VSUBS 0.008821f
C889 B.n240 VSUBS 0.008821f
C890 B.n241 VSUBS 0.008821f
C891 B.n242 VSUBS 0.008821f
C892 B.n243 VSUBS 0.008821f
C893 B.n244 VSUBS 0.008821f
C894 B.n245 VSUBS 0.008821f
C895 B.n246 VSUBS 0.008821f
C896 B.n247 VSUBS 0.008821f
C897 B.n248 VSUBS 0.008821f
C898 B.n249 VSUBS 0.008821f
C899 B.n250 VSUBS 0.008821f
C900 B.n251 VSUBS 0.008821f
C901 B.n252 VSUBS 0.008821f
C902 B.n253 VSUBS 0.008821f
C903 B.n254 VSUBS 0.008821f
C904 B.n255 VSUBS 0.008821f
C905 B.n256 VSUBS 0.008821f
C906 B.n257 VSUBS 0.008821f
C907 B.n258 VSUBS 0.008821f
C908 B.n259 VSUBS 0.008821f
C909 B.n260 VSUBS 0.008821f
C910 B.n261 VSUBS 0.008821f
C911 B.n262 VSUBS 0.008821f
C912 B.n263 VSUBS 0.008821f
C913 B.n264 VSUBS 0.008821f
C914 B.n265 VSUBS 0.008821f
C915 B.n266 VSUBS 0.008821f
C916 B.n267 VSUBS 0.008821f
C917 B.n268 VSUBS 0.008821f
C918 B.n269 VSUBS 0.008821f
C919 B.n270 VSUBS 0.008821f
C920 B.n271 VSUBS 0.008821f
C921 B.n272 VSUBS 0.008821f
C922 B.n273 VSUBS 0.008821f
C923 B.n274 VSUBS 0.008821f
C924 B.n275 VSUBS 0.008821f
C925 B.n276 VSUBS 0.008821f
C926 B.n277 VSUBS 0.008821f
C927 B.n278 VSUBS 0.008821f
C928 B.n279 VSUBS 0.008821f
C929 B.n280 VSUBS 0.008821f
C930 B.n281 VSUBS 0.008821f
C931 B.n282 VSUBS 0.019834f
C932 B.n283 VSUBS 0.019834f
C933 B.n284 VSUBS 0.020897f
C934 B.n285 VSUBS 0.008821f
C935 B.n286 VSUBS 0.008821f
C936 B.n287 VSUBS 0.008821f
C937 B.n288 VSUBS 0.008821f
C938 B.n289 VSUBS 0.008821f
C939 B.n290 VSUBS 0.008821f
C940 B.n291 VSUBS 0.008821f
C941 B.n292 VSUBS 0.008821f
C942 B.n293 VSUBS 0.008821f
C943 B.n294 VSUBS 0.008821f
C944 B.n295 VSUBS 0.008821f
C945 B.n296 VSUBS 0.008821f
C946 B.n297 VSUBS 0.008821f
C947 B.n298 VSUBS 0.008821f
C948 B.n299 VSUBS 0.008821f
C949 B.n300 VSUBS 0.008821f
C950 B.n301 VSUBS 0.008821f
C951 B.n302 VSUBS 0.008821f
C952 B.n303 VSUBS 0.008821f
C953 B.n304 VSUBS 0.008821f
C954 B.n305 VSUBS 0.008821f
C955 B.n306 VSUBS 0.008821f
C956 B.n307 VSUBS 0.008821f
C957 B.n308 VSUBS 0.008821f
C958 B.n309 VSUBS 0.008821f
C959 B.n310 VSUBS 0.008821f
C960 B.n311 VSUBS 0.008821f
C961 B.n312 VSUBS 0.008821f
C962 B.n313 VSUBS 0.008821f
C963 B.n314 VSUBS 0.008821f
C964 B.n315 VSUBS 0.008821f
C965 B.n316 VSUBS 0.008821f
C966 B.n317 VSUBS 0.008821f
C967 B.n318 VSUBS 0.008821f
C968 B.n319 VSUBS 0.008821f
C969 B.n320 VSUBS 0.008821f
C970 B.n321 VSUBS 0.008821f
C971 B.n322 VSUBS 0.008821f
C972 B.n323 VSUBS 0.008821f
C973 B.n324 VSUBS 0.008821f
C974 B.n325 VSUBS 0.008821f
C975 B.n326 VSUBS 0.008821f
C976 B.n327 VSUBS 0.008821f
C977 B.n328 VSUBS 0.008821f
C978 B.n329 VSUBS 0.008821f
C979 B.n330 VSUBS 0.008821f
C980 B.n331 VSUBS 0.008821f
C981 B.n332 VSUBS 0.008821f
C982 B.n333 VSUBS 0.008821f
C983 B.n334 VSUBS 0.008821f
C984 B.n335 VSUBS 0.008821f
C985 B.n336 VSUBS 0.008821f
C986 B.n337 VSUBS 0.008821f
C987 B.n338 VSUBS 0.008821f
C988 B.n339 VSUBS 0.006097f
C989 B.n340 VSUBS 0.008821f
C990 B.n341 VSUBS 0.008821f
C991 B.n342 VSUBS 0.007134f
C992 B.n343 VSUBS 0.008821f
C993 B.n344 VSUBS 0.008821f
C994 B.n345 VSUBS 0.008821f
C995 B.n346 VSUBS 0.008821f
C996 B.n347 VSUBS 0.008821f
C997 B.n348 VSUBS 0.008821f
C998 B.n349 VSUBS 0.008821f
C999 B.n350 VSUBS 0.008821f
C1000 B.n351 VSUBS 0.008821f
C1001 B.n352 VSUBS 0.008821f
C1002 B.n353 VSUBS 0.008821f
C1003 B.n354 VSUBS 0.007134f
C1004 B.n355 VSUBS 0.020437f
C1005 B.n356 VSUBS 0.006097f
C1006 B.n357 VSUBS 0.008821f
C1007 B.n358 VSUBS 0.008821f
C1008 B.n359 VSUBS 0.008821f
C1009 B.n360 VSUBS 0.008821f
C1010 B.n361 VSUBS 0.008821f
C1011 B.n362 VSUBS 0.008821f
C1012 B.n363 VSUBS 0.008821f
C1013 B.n364 VSUBS 0.008821f
C1014 B.n365 VSUBS 0.008821f
C1015 B.n366 VSUBS 0.008821f
C1016 B.n367 VSUBS 0.008821f
C1017 B.n368 VSUBS 0.008821f
C1018 B.n369 VSUBS 0.008821f
C1019 B.n370 VSUBS 0.008821f
C1020 B.n371 VSUBS 0.008821f
C1021 B.n372 VSUBS 0.008821f
C1022 B.n373 VSUBS 0.008821f
C1023 B.n374 VSUBS 0.008821f
C1024 B.n375 VSUBS 0.008821f
C1025 B.n376 VSUBS 0.008821f
C1026 B.n377 VSUBS 0.008821f
C1027 B.n378 VSUBS 0.008821f
C1028 B.n379 VSUBS 0.008821f
C1029 B.n380 VSUBS 0.008821f
C1030 B.n381 VSUBS 0.008821f
C1031 B.n382 VSUBS 0.008821f
C1032 B.n383 VSUBS 0.008821f
C1033 B.n384 VSUBS 0.008821f
C1034 B.n385 VSUBS 0.008821f
C1035 B.n386 VSUBS 0.008821f
C1036 B.n387 VSUBS 0.008821f
C1037 B.n388 VSUBS 0.008821f
C1038 B.n389 VSUBS 0.008821f
C1039 B.n390 VSUBS 0.008821f
C1040 B.n391 VSUBS 0.008821f
C1041 B.n392 VSUBS 0.008821f
C1042 B.n393 VSUBS 0.008821f
C1043 B.n394 VSUBS 0.008821f
C1044 B.n395 VSUBS 0.008821f
C1045 B.n396 VSUBS 0.008821f
C1046 B.n397 VSUBS 0.008821f
C1047 B.n398 VSUBS 0.008821f
C1048 B.n399 VSUBS 0.008821f
C1049 B.n400 VSUBS 0.008821f
C1050 B.n401 VSUBS 0.008821f
C1051 B.n402 VSUBS 0.008821f
C1052 B.n403 VSUBS 0.008821f
C1053 B.n404 VSUBS 0.008821f
C1054 B.n405 VSUBS 0.008821f
C1055 B.n406 VSUBS 0.008821f
C1056 B.n407 VSUBS 0.008821f
C1057 B.n408 VSUBS 0.008821f
C1058 B.n409 VSUBS 0.008821f
C1059 B.n410 VSUBS 0.008821f
C1060 B.n411 VSUBS 0.020897f
C1061 B.n412 VSUBS 0.020897f
C1062 B.n413 VSUBS 0.019834f
C1063 B.n414 VSUBS 0.008821f
C1064 B.n415 VSUBS 0.008821f
C1065 B.n416 VSUBS 0.008821f
C1066 B.n417 VSUBS 0.008821f
C1067 B.n418 VSUBS 0.008821f
C1068 B.n419 VSUBS 0.008821f
C1069 B.n420 VSUBS 0.008821f
C1070 B.n421 VSUBS 0.008821f
C1071 B.n422 VSUBS 0.008821f
C1072 B.n423 VSUBS 0.008821f
C1073 B.n424 VSUBS 0.008821f
C1074 B.n425 VSUBS 0.008821f
C1075 B.n426 VSUBS 0.008821f
C1076 B.n427 VSUBS 0.008821f
C1077 B.n428 VSUBS 0.008821f
C1078 B.n429 VSUBS 0.008821f
C1079 B.n430 VSUBS 0.008821f
C1080 B.n431 VSUBS 0.008821f
C1081 B.n432 VSUBS 0.008821f
C1082 B.n433 VSUBS 0.008821f
C1083 B.n434 VSUBS 0.008821f
C1084 B.n435 VSUBS 0.008821f
C1085 B.n436 VSUBS 0.008821f
C1086 B.n437 VSUBS 0.008821f
C1087 B.n438 VSUBS 0.008821f
C1088 B.n439 VSUBS 0.008821f
C1089 B.n440 VSUBS 0.008821f
C1090 B.n441 VSUBS 0.008821f
C1091 B.n442 VSUBS 0.008821f
C1092 B.n443 VSUBS 0.008821f
C1093 B.n444 VSUBS 0.008821f
C1094 B.n445 VSUBS 0.008821f
C1095 B.n446 VSUBS 0.008821f
C1096 B.n447 VSUBS 0.008821f
C1097 B.n448 VSUBS 0.008821f
C1098 B.n449 VSUBS 0.008821f
C1099 B.n450 VSUBS 0.008821f
C1100 B.n451 VSUBS 0.008821f
C1101 B.n452 VSUBS 0.008821f
C1102 B.n453 VSUBS 0.008821f
C1103 B.n454 VSUBS 0.008821f
C1104 B.n455 VSUBS 0.008821f
C1105 B.n456 VSUBS 0.008821f
C1106 B.n457 VSUBS 0.008821f
C1107 B.n458 VSUBS 0.008821f
C1108 B.n459 VSUBS 0.008821f
C1109 B.n460 VSUBS 0.008821f
C1110 B.n461 VSUBS 0.008821f
C1111 B.n462 VSUBS 0.008821f
C1112 B.n463 VSUBS 0.008821f
C1113 B.n464 VSUBS 0.008821f
C1114 B.n465 VSUBS 0.008821f
C1115 B.n466 VSUBS 0.008821f
C1116 B.n467 VSUBS 0.008821f
C1117 B.n468 VSUBS 0.008821f
C1118 B.n469 VSUBS 0.008821f
C1119 B.n470 VSUBS 0.008821f
C1120 B.n471 VSUBS 0.008821f
C1121 B.n472 VSUBS 0.008821f
C1122 B.n473 VSUBS 0.008821f
C1123 B.n474 VSUBS 0.008821f
C1124 B.n475 VSUBS 0.008821f
C1125 B.n476 VSUBS 0.008821f
C1126 B.n477 VSUBS 0.008821f
C1127 B.n478 VSUBS 0.008821f
C1128 B.n479 VSUBS 0.008821f
C1129 B.n480 VSUBS 0.008821f
C1130 B.n481 VSUBS 0.008821f
C1131 B.n482 VSUBS 0.008821f
C1132 B.n483 VSUBS 0.008821f
C1133 B.n484 VSUBS 0.008821f
C1134 B.n485 VSUBS 0.008821f
C1135 B.n486 VSUBS 0.008821f
C1136 B.n487 VSUBS 0.008821f
C1137 B.n488 VSUBS 0.008821f
C1138 B.n489 VSUBS 0.008821f
C1139 B.n490 VSUBS 0.008821f
C1140 B.n491 VSUBS 0.008821f
C1141 B.n492 VSUBS 0.008821f
C1142 B.n493 VSUBS 0.008821f
C1143 B.n494 VSUBS 0.008821f
C1144 B.n495 VSUBS 0.008821f
C1145 B.n496 VSUBS 0.008821f
C1146 B.n497 VSUBS 0.008821f
C1147 B.n498 VSUBS 0.008821f
C1148 B.n499 VSUBS 0.008821f
C1149 B.n500 VSUBS 0.008821f
C1150 B.n501 VSUBS 0.008821f
C1151 B.n502 VSUBS 0.008821f
C1152 B.n503 VSUBS 0.008821f
C1153 B.n504 VSUBS 0.008821f
C1154 B.n505 VSUBS 0.008821f
C1155 B.n506 VSUBS 0.008821f
C1156 B.n507 VSUBS 0.008821f
C1157 B.n508 VSUBS 0.008821f
C1158 B.n509 VSUBS 0.008821f
C1159 B.n510 VSUBS 0.008821f
C1160 B.n511 VSUBS 0.008821f
C1161 B.n512 VSUBS 0.008821f
C1162 B.n513 VSUBS 0.008821f
C1163 B.n514 VSUBS 0.008821f
C1164 B.n515 VSUBS 0.008821f
C1165 B.n516 VSUBS 0.008821f
C1166 B.n517 VSUBS 0.008821f
C1167 B.n518 VSUBS 0.008821f
C1168 B.n519 VSUBS 0.008821f
C1169 B.n520 VSUBS 0.008821f
C1170 B.n521 VSUBS 0.008821f
C1171 B.n522 VSUBS 0.008821f
C1172 B.n523 VSUBS 0.008821f
C1173 B.n524 VSUBS 0.008821f
C1174 B.n525 VSUBS 0.008821f
C1175 B.n526 VSUBS 0.008821f
C1176 B.n527 VSUBS 0.008821f
C1177 B.n528 VSUBS 0.008821f
C1178 B.n529 VSUBS 0.008821f
C1179 B.n530 VSUBS 0.008821f
C1180 B.n531 VSUBS 0.008821f
C1181 B.n532 VSUBS 0.008821f
C1182 B.n533 VSUBS 0.008821f
C1183 B.n534 VSUBS 0.008821f
C1184 B.n535 VSUBS 0.008821f
C1185 B.n536 VSUBS 0.008821f
C1186 B.n537 VSUBS 0.008821f
C1187 B.n538 VSUBS 0.008821f
C1188 B.n539 VSUBS 0.008821f
C1189 B.n540 VSUBS 0.008821f
C1190 B.n541 VSUBS 0.008821f
C1191 B.n542 VSUBS 0.008821f
C1192 B.n543 VSUBS 0.008821f
C1193 B.n544 VSUBS 0.008821f
C1194 B.n545 VSUBS 0.008821f
C1195 B.n546 VSUBS 0.008821f
C1196 B.n547 VSUBS 0.008821f
C1197 B.n548 VSUBS 0.008821f
C1198 B.n549 VSUBS 0.008821f
C1199 B.n550 VSUBS 0.008821f
C1200 B.n551 VSUBS 0.008821f
C1201 B.n552 VSUBS 0.008821f
C1202 B.n553 VSUBS 0.008821f
C1203 B.n554 VSUBS 0.008821f
C1204 B.n555 VSUBS 0.008821f
C1205 B.n556 VSUBS 0.008821f
C1206 B.n557 VSUBS 0.008821f
C1207 B.n558 VSUBS 0.008821f
C1208 B.n559 VSUBS 0.008821f
C1209 B.n560 VSUBS 0.008821f
C1210 B.n561 VSUBS 0.008821f
C1211 B.n562 VSUBS 0.008821f
C1212 B.n563 VSUBS 0.008821f
C1213 B.n564 VSUBS 0.008821f
C1214 B.n565 VSUBS 0.008821f
C1215 B.n566 VSUBS 0.008821f
C1216 B.n567 VSUBS 0.008821f
C1217 B.n568 VSUBS 0.008821f
C1218 B.n569 VSUBS 0.008821f
C1219 B.n570 VSUBS 0.008821f
C1220 B.n571 VSUBS 0.008821f
C1221 B.n572 VSUBS 0.008821f
C1222 B.n573 VSUBS 0.008821f
C1223 B.n574 VSUBS 0.008821f
C1224 B.n575 VSUBS 0.019834f
C1225 B.n576 VSUBS 0.020897f
C1226 B.n577 VSUBS 0.019834f
C1227 B.n578 VSUBS 0.008821f
C1228 B.n579 VSUBS 0.008821f
C1229 B.n580 VSUBS 0.008821f
C1230 B.n581 VSUBS 0.008821f
C1231 B.n582 VSUBS 0.008821f
C1232 B.n583 VSUBS 0.008821f
C1233 B.n584 VSUBS 0.008821f
C1234 B.n585 VSUBS 0.008821f
C1235 B.n586 VSUBS 0.008821f
C1236 B.n587 VSUBS 0.008821f
C1237 B.n588 VSUBS 0.008821f
C1238 B.n589 VSUBS 0.008821f
C1239 B.n590 VSUBS 0.008821f
C1240 B.n591 VSUBS 0.008821f
C1241 B.n592 VSUBS 0.008821f
C1242 B.n593 VSUBS 0.008821f
C1243 B.n594 VSUBS 0.008821f
C1244 B.n595 VSUBS 0.008821f
C1245 B.n596 VSUBS 0.008821f
C1246 B.n597 VSUBS 0.008821f
C1247 B.n598 VSUBS 0.008821f
C1248 B.n599 VSUBS 0.008821f
C1249 B.n600 VSUBS 0.008821f
C1250 B.n601 VSUBS 0.008821f
C1251 B.n602 VSUBS 0.008821f
C1252 B.n603 VSUBS 0.008821f
C1253 B.n604 VSUBS 0.008821f
C1254 B.n605 VSUBS 0.008821f
C1255 B.n606 VSUBS 0.008821f
C1256 B.n607 VSUBS 0.008821f
C1257 B.n608 VSUBS 0.008821f
C1258 B.n609 VSUBS 0.008821f
C1259 B.n610 VSUBS 0.008821f
C1260 B.n611 VSUBS 0.008821f
C1261 B.n612 VSUBS 0.008821f
C1262 B.n613 VSUBS 0.008821f
C1263 B.n614 VSUBS 0.008821f
C1264 B.n615 VSUBS 0.008821f
C1265 B.n616 VSUBS 0.008821f
C1266 B.n617 VSUBS 0.008821f
C1267 B.n618 VSUBS 0.008821f
C1268 B.n619 VSUBS 0.008821f
C1269 B.n620 VSUBS 0.008821f
C1270 B.n621 VSUBS 0.008821f
C1271 B.n622 VSUBS 0.008821f
C1272 B.n623 VSUBS 0.008821f
C1273 B.n624 VSUBS 0.008821f
C1274 B.n625 VSUBS 0.008821f
C1275 B.n626 VSUBS 0.008821f
C1276 B.n627 VSUBS 0.008821f
C1277 B.n628 VSUBS 0.008821f
C1278 B.n629 VSUBS 0.008821f
C1279 B.n630 VSUBS 0.008821f
C1280 B.n631 VSUBS 0.008821f
C1281 B.n632 VSUBS 0.006097f
C1282 B.n633 VSUBS 0.020437f
C1283 B.n634 VSUBS 0.007134f
C1284 B.n635 VSUBS 0.008821f
C1285 B.n636 VSUBS 0.008821f
C1286 B.n637 VSUBS 0.008821f
C1287 B.n638 VSUBS 0.008821f
C1288 B.n639 VSUBS 0.008821f
C1289 B.n640 VSUBS 0.008821f
C1290 B.n641 VSUBS 0.008821f
C1291 B.n642 VSUBS 0.008821f
C1292 B.n643 VSUBS 0.008821f
C1293 B.n644 VSUBS 0.008821f
C1294 B.n645 VSUBS 0.008821f
C1295 B.n646 VSUBS 0.007134f
C1296 B.n647 VSUBS 0.008821f
C1297 B.n648 VSUBS 0.008821f
C1298 B.n649 VSUBS 0.006097f
C1299 B.n650 VSUBS 0.008821f
C1300 B.n651 VSUBS 0.008821f
C1301 B.n652 VSUBS 0.008821f
C1302 B.n653 VSUBS 0.008821f
C1303 B.n654 VSUBS 0.008821f
C1304 B.n655 VSUBS 0.008821f
C1305 B.n656 VSUBS 0.008821f
C1306 B.n657 VSUBS 0.008821f
C1307 B.n658 VSUBS 0.008821f
C1308 B.n659 VSUBS 0.008821f
C1309 B.n660 VSUBS 0.008821f
C1310 B.n661 VSUBS 0.008821f
C1311 B.n662 VSUBS 0.008821f
C1312 B.n663 VSUBS 0.008821f
C1313 B.n664 VSUBS 0.008821f
C1314 B.n665 VSUBS 0.008821f
C1315 B.n666 VSUBS 0.008821f
C1316 B.n667 VSUBS 0.008821f
C1317 B.n668 VSUBS 0.008821f
C1318 B.n669 VSUBS 0.008821f
C1319 B.n670 VSUBS 0.008821f
C1320 B.n671 VSUBS 0.008821f
C1321 B.n672 VSUBS 0.008821f
C1322 B.n673 VSUBS 0.008821f
C1323 B.n674 VSUBS 0.008821f
C1324 B.n675 VSUBS 0.008821f
C1325 B.n676 VSUBS 0.008821f
C1326 B.n677 VSUBS 0.008821f
C1327 B.n678 VSUBS 0.008821f
C1328 B.n679 VSUBS 0.008821f
C1329 B.n680 VSUBS 0.008821f
C1330 B.n681 VSUBS 0.008821f
C1331 B.n682 VSUBS 0.008821f
C1332 B.n683 VSUBS 0.008821f
C1333 B.n684 VSUBS 0.008821f
C1334 B.n685 VSUBS 0.008821f
C1335 B.n686 VSUBS 0.008821f
C1336 B.n687 VSUBS 0.008821f
C1337 B.n688 VSUBS 0.008821f
C1338 B.n689 VSUBS 0.008821f
C1339 B.n690 VSUBS 0.008821f
C1340 B.n691 VSUBS 0.008821f
C1341 B.n692 VSUBS 0.008821f
C1342 B.n693 VSUBS 0.008821f
C1343 B.n694 VSUBS 0.008821f
C1344 B.n695 VSUBS 0.008821f
C1345 B.n696 VSUBS 0.008821f
C1346 B.n697 VSUBS 0.008821f
C1347 B.n698 VSUBS 0.008821f
C1348 B.n699 VSUBS 0.008821f
C1349 B.n700 VSUBS 0.008821f
C1350 B.n701 VSUBS 0.008821f
C1351 B.n702 VSUBS 0.008821f
C1352 B.n703 VSUBS 0.008821f
C1353 B.n704 VSUBS 0.020897f
C1354 B.n705 VSUBS 0.019834f
C1355 B.n706 VSUBS 0.019834f
C1356 B.n707 VSUBS 0.008821f
C1357 B.n708 VSUBS 0.008821f
C1358 B.n709 VSUBS 0.008821f
C1359 B.n710 VSUBS 0.008821f
C1360 B.n711 VSUBS 0.008821f
C1361 B.n712 VSUBS 0.008821f
C1362 B.n713 VSUBS 0.008821f
C1363 B.n714 VSUBS 0.008821f
C1364 B.n715 VSUBS 0.008821f
C1365 B.n716 VSUBS 0.008821f
C1366 B.n717 VSUBS 0.008821f
C1367 B.n718 VSUBS 0.008821f
C1368 B.n719 VSUBS 0.008821f
C1369 B.n720 VSUBS 0.008821f
C1370 B.n721 VSUBS 0.008821f
C1371 B.n722 VSUBS 0.008821f
C1372 B.n723 VSUBS 0.008821f
C1373 B.n724 VSUBS 0.008821f
C1374 B.n725 VSUBS 0.008821f
C1375 B.n726 VSUBS 0.008821f
C1376 B.n727 VSUBS 0.008821f
C1377 B.n728 VSUBS 0.008821f
C1378 B.n729 VSUBS 0.008821f
C1379 B.n730 VSUBS 0.008821f
C1380 B.n731 VSUBS 0.008821f
C1381 B.n732 VSUBS 0.008821f
C1382 B.n733 VSUBS 0.008821f
C1383 B.n734 VSUBS 0.008821f
C1384 B.n735 VSUBS 0.008821f
C1385 B.n736 VSUBS 0.008821f
C1386 B.n737 VSUBS 0.008821f
C1387 B.n738 VSUBS 0.008821f
C1388 B.n739 VSUBS 0.008821f
C1389 B.n740 VSUBS 0.008821f
C1390 B.n741 VSUBS 0.008821f
C1391 B.n742 VSUBS 0.008821f
C1392 B.n743 VSUBS 0.008821f
C1393 B.n744 VSUBS 0.008821f
C1394 B.n745 VSUBS 0.008821f
C1395 B.n746 VSUBS 0.008821f
C1396 B.n747 VSUBS 0.008821f
C1397 B.n748 VSUBS 0.008821f
C1398 B.n749 VSUBS 0.008821f
C1399 B.n750 VSUBS 0.008821f
C1400 B.n751 VSUBS 0.008821f
C1401 B.n752 VSUBS 0.008821f
C1402 B.n753 VSUBS 0.008821f
C1403 B.n754 VSUBS 0.008821f
C1404 B.n755 VSUBS 0.008821f
C1405 B.n756 VSUBS 0.008821f
C1406 B.n757 VSUBS 0.008821f
C1407 B.n758 VSUBS 0.008821f
C1408 B.n759 VSUBS 0.008821f
C1409 B.n760 VSUBS 0.008821f
C1410 B.n761 VSUBS 0.008821f
C1411 B.n762 VSUBS 0.008821f
C1412 B.n763 VSUBS 0.008821f
C1413 B.n764 VSUBS 0.008821f
C1414 B.n765 VSUBS 0.008821f
C1415 B.n766 VSUBS 0.008821f
C1416 B.n767 VSUBS 0.008821f
C1417 B.n768 VSUBS 0.008821f
C1418 B.n769 VSUBS 0.008821f
C1419 B.n770 VSUBS 0.008821f
C1420 B.n771 VSUBS 0.008821f
C1421 B.n772 VSUBS 0.008821f
C1422 B.n773 VSUBS 0.008821f
C1423 B.n774 VSUBS 0.008821f
C1424 B.n775 VSUBS 0.008821f
C1425 B.n776 VSUBS 0.008821f
C1426 B.n777 VSUBS 0.008821f
C1427 B.n778 VSUBS 0.008821f
C1428 B.n779 VSUBS 0.008821f
C1429 B.n780 VSUBS 0.008821f
C1430 B.n781 VSUBS 0.008821f
C1431 B.n782 VSUBS 0.008821f
C1432 B.n783 VSUBS 0.008821f
C1433 B.n784 VSUBS 0.008821f
C1434 B.n785 VSUBS 0.008821f
C1435 B.n786 VSUBS 0.008821f
C1436 B.n787 VSUBS 0.019973f
.ends

