* NGSPICE file created from diff_pair_sample_1266.ext - technology: sky130A

.subckt diff_pair_sample_1266 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0.19305 ps=1.5 w=1.17 l=3.01
X1 VTAIL.t0 VP.t0 VDD1.t5 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.19305 ps=1.5 w=1.17 l=3.01
X2 VDD1.t4 VP.t1 VTAIL.t1 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0.19305 ps=1.5 w=1.17 l=3.01
X3 VDD2.t4 VN.t1 VTAIL.t7 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.4563 ps=3.12 w=1.17 l=3.01
X4 B.t11 B.t9 B.t10 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0 ps=0 w=1.17 l=3.01
X5 VTAIL.t3 VP.t2 VDD1.t3 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.19305 ps=1.5 w=1.17 l=3.01
X6 B.t8 B.t6 B.t7 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0 ps=0 w=1.17 l=3.01
X7 VTAIL.t9 VN.t2 VDD2.t3 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.19305 ps=1.5 w=1.17 l=3.01
X8 VTAIL.t11 VN.t3 VDD2.t2 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.19305 ps=1.5 w=1.17 l=3.01
X9 B.t5 B.t3 B.t4 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0 ps=0 w=1.17 l=3.01
X10 VDD2.t1 VN.t4 VTAIL.t10 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.4563 ps=3.12 w=1.17 l=3.01
X11 VDD1.t2 VP.t3 VTAIL.t4 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.4563 ps=3.12 w=1.17 l=3.01
X12 VDD1.t1 VP.t4 VTAIL.t5 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0.19305 ps=1.5 w=1.17 l=3.01
X13 VDD2.t0 VN.t5 VTAIL.t6 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0.19305 ps=1.5 w=1.17 l=3.01
X14 VDD1.t0 VP.t5 VTAIL.t2 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.19305 pd=1.5 as=0.4563 ps=3.12 w=1.17 l=3.01
X15 B.t2 B.t0 B.t1 w_n3642_n1202# sky130_fd_pr__pfet_01v8 ad=0.4563 pd=3.12 as=0 ps=0 w=1.17 l=3.01
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n15 VN.n0 73.4298
R13 VN.n31 VN.n16 73.4298
R14 VN.n11 VN.n2 56.5193
R15 VN.n27 VN.n18 56.5193
R16 VN.n5 VN.n4 49.2372
R17 VN.n21 VN.n20 49.2372
R18 VN.n20 VN.t1 42.6169
R19 VN.n4 VN.t0 42.6169
R20 VN VN.n31 42.3162
R21 VN.n6 VN.n5 24.4675
R22 VN.n7 VN.n6 24.4675
R23 VN.n7 VN.n2 24.4675
R24 VN.n12 VN.n11 24.4675
R25 VN.n13 VN.n12 24.4675
R26 VN.n23 VN.n18 24.4675
R27 VN.n23 VN.n22 24.4675
R28 VN.n22 VN.n21 24.4675
R29 VN.n29 VN.n28 24.4675
R30 VN.n28 VN.n27 24.4675
R31 VN.n13 VN.n0 16.6381
R32 VN.n29 VN.n16 16.6381
R33 VN.n5 VN.t3 9.36827
R34 VN.n0 VN.t4 9.36827
R35 VN.n21 VN.t2 9.36827
R36 VN.n16 VN.t5 9.36827
R37 VN.n20 VN.n19 4.07659
R38 VN.n4 VN.n3 4.07659
R39 VN.n31 VN.n30 0.354971
R40 VN.n15 VN.n14 0.354971
R41 VN VN.n15 0.26696
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n11 VTAIL.t10 373.88
R53 VTAIL.n2 VTAIL.t4 373.88
R54 VTAIL.n10 VTAIL.t2 373.88
R55 VTAIL.n7 VTAIL.t7 373.88
R56 VTAIL.n1 VTAIL.n0 330.942
R57 VTAIL.n4 VTAIL.n3 330.942
R58 VTAIL.n9 VTAIL.n8 330.942
R59 VTAIL.n6 VTAIL.n5 330.942
R60 VTAIL.n0 VTAIL.t8 27.7826
R61 VTAIL.n0 VTAIL.t11 27.7826
R62 VTAIL.n3 VTAIL.t1 27.7826
R63 VTAIL.n3 VTAIL.t3 27.7826
R64 VTAIL.n8 VTAIL.t5 27.7826
R65 VTAIL.n8 VTAIL.t0 27.7826
R66 VTAIL.n5 VTAIL.t6 27.7826
R67 VTAIL.n5 VTAIL.t9 27.7826
R68 VTAIL.n6 VTAIL.n4 19.1341
R69 VTAIL.n11 VTAIL.n10 16.2548
R70 VTAIL.n7 VTAIL.n6 2.87981
R71 VTAIL.n10 VTAIL.n9 2.87981
R72 VTAIL.n4 VTAIL.n2 2.87981
R73 VTAIL VTAIL.n11 2.10179
R74 VTAIL.n9 VTAIL.n7 1.90998
R75 VTAIL.n2 VTAIL.n1 1.90998
R76 VTAIL VTAIL.n1 0.778517
R77 VDD2.n1 VDD2.t5 392.663
R78 VDD2.n2 VDD2.t0 390.558
R79 VDD2.n1 VDD2.n0 348.286
R80 VDD2 VDD2.n3 348.284
R81 VDD2.n2 VDD2.n1 34.0817
R82 VDD2.n3 VDD2.t3 27.7826
R83 VDD2.n3 VDD2.t4 27.7826
R84 VDD2.n0 VDD2.t2 27.7826
R85 VDD2.n0 VDD2.t1 27.7826
R86 VDD2 VDD2.n2 2.21817
R87 VP.n13 VP.n10 161.3
R88 VP.n15 VP.n14 161.3
R89 VP.n16 VP.n9 161.3
R90 VP.n18 VP.n17 161.3
R91 VP.n19 VP.n8 161.3
R92 VP.n21 VP.n20 161.3
R93 VP.n44 VP.n43 161.3
R94 VP.n42 VP.n1 161.3
R95 VP.n41 VP.n40 161.3
R96 VP.n39 VP.n2 161.3
R97 VP.n38 VP.n37 161.3
R98 VP.n36 VP.n3 161.3
R99 VP.n35 VP.n34 161.3
R100 VP.n33 VP.n4 161.3
R101 VP.n32 VP.n31 161.3
R102 VP.n30 VP.n5 161.3
R103 VP.n29 VP.n28 161.3
R104 VP.n27 VP.n6 161.3
R105 VP.n26 VP.n25 161.3
R106 VP.n24 VP.n23 73.4298
R107 VP.n45 VP.n0 73.4298
R108 VP.n22 VP.n7 73.4298
R109 VP.n30 VP.n29 56.5193
R110 VP.n41 VP.n2 56.5193
R111 VP.n18 VP.n9 56.5193
R112 VP.n12 VP.n11 49.2372
R113 VP.n11 VP.t4 42.6167
R114 VP.n23 VP.n22 42.1508
R115 VP.n25 VP.n6 24.4675
R116 VP.n29 VP.n6 24.4675
R117 VP.n31 VP.n30 24.4675
R118 VP.n31 VP.n4 24.4675
R119 VP.n35 VP.n4 24.4675
R120 VP.n36 VP.n35 24.4675
R121 VP.n37 VP.n36 24.4675
R122 VP.n37 VP.n2 24.4675
R123 VP.n42 VP.n41 24.4675
R124 VP.n43 VP.n42 24.4675
R125 VP.n19 VP.n18 24.4675
R126 VP.n20 VP.n19 24.4675
R127 VP.n13 VP.n12 24.4675
R128 VP.n14 VP.n13 24.4675
R129 VP.n14 VP.n9 24.4675
R130 VP.n25 VP.n24 16.6381
R131 VP.n43 VP.n0 16.6381
R132 VP.n20 VP.n7 16.6381
R133 VP.n35 VP.t2 9.36827
R134 VP.n24 VP.t1 9.36827
R135 VP.n0 VP.t3 9.36827
R136 VP.n12 VP.t0 9.36827
R137 VP.n7 VP.t5 9.36827
R138 VP.n11 VP.n10 4.07657
R139 VP.n22 VP.n21 0.354971
R140 VP.n26 VP.n23 0.354971
R141 VP.n45 VP.n44 0.354971
R142 VP VP.n45 0.26696
R143 VP.n15 VP.n10 0.189894
R144 VP.n16 VP.n15 0.189894
R145 VP.n17 VP.n16 0.189894
R146 VP.n17 VP.n8 0.189894
R147 VP.n21 VP.n8 0.189894
R148 VP.n27 VP.n26 0.189894
R149 VP.n28 VP.n27 0.189894
R150 VP.n28 VP.n5 0.189894
R151 VP.n32 VP.n5 0.189894
R152 VP.n33 VP.n32 0.189894
R153 VP.n34 VP.n33 0.189894
R154 VP.n34 VP.n3 0.189894
R155 VP.n38 VP.n3 0.189894
R156 VP.n39 VP.n38 0.189894
R157 VP.n40 VP.n39 0.189894
R158 VP.n40 VP.n1 0.189894
R159 VP.n44 VP.n1 0.189894
R160 VDD1 VDD1.t1 392.776
R161 VDD1.n1 VDD1.t4 392.663
R162 VDD1.n1 VDD1.n0 348.286
R163 VDD1.n3 VDD1.n2 347.622
R164 VDD1.n3 VDD1.n1 36.1043
R165 VDD1.n2 VDD1.t5 27.7826
R166 VDD1.n2 VDD1.t0 27.7826
R167 VDD1.n0 VDD1.t3 27.7826
R168 VDD1.n0 VDD1.t2 27.7826
R169 VDD1 VDD1.n3 0.662138
R170 B.n248 B.n93 585
R171 B.n247 B.n246 585
R172 B.n245 B.n94 585
R173 B.n244 B.n243 585
R174 B.n242 B.n95 585
R175 B.n241 B.n240 585
R176 B.n239 B.n96 585
R177 B.n238 B.n237 585
R178 B.n236 B.n97 585
R179 B.n235 B.n234 585
R180 B.n232 B.n98 585
R181 B.n231 B.n230 585
R182 B.n229 B.n101 585
R183 B.n228 B.n227 585
R184 B.n226 B.n102 585
R185 B.n225 B.n224 585
R186 B.n223 B.n103 585
R187 B.n222 B.n221 585
R188 B.n220 B.n104 585
R189 B.n218 B.n217 585
R190 B.n216 B.n107 585
R191 B.n215 B.n214 585
R192 B.n213 B.n108 585
R193 B.n212 B.n211 585
R194 B.n210 B.n109 585
R195 B.n209 B.n208 585
R196 B.n207 B.n110 585
R197 B.n206 B.n205 585
R198 B.n204 B.n111 585
R199 B.n250 B.n249 585
R200 B.n251 B.n92 585
R201 B.n253 B.n252 585
R202 B.n254 B.n91 585
R203 B.n256 B.n255 585
R204 B.n257 B.n90 585
R205 B.n259 B.n258 585
R206 B.n260 B.n89 585
R207 B.n262 B.n261 585
R208 B.n263 B.n88 585
R209 B.n265 B.n264 585
R210 B.n266 B.n87 585
R211 B.n268 B.n267 585
R212 B.n269 B.n86 585
R213 B.n271 B.n270 585
R214 B.n272 B.n85 585
R215 B.n274 B.n273 585
R216 B.n275 B.n84 585
R217 B.n277 B.n276 585
R218 B.n278 B.n83 585
R219 B.n280 B.n279 585
R220 B.n281 B.n82 585
R221 B.n283 B.n282 585
R222 B.n284 B.n81 585
R223 B.n286 B.n285 585
R224 B.n287 B.n80 585
R225 B.n289 B.n288 585
R226 B.n290 B.n79 585
R227 B.n292 B.n291 585
R228 B.n293 B.n78 585
R229 B.n295 B.n294 585
R230 B.n296 B.n77 585
R231 B.n298 B.n297 585
R232 B.n299 B.n76 585
R233 B.n301 B.n300 585
R234 B.n302 B.n75 585
R235 B.n304 B.n303 585
R236 B.n305 B.n74 585
R237 B.n307 B.n306 585
R238 B.n308 B.n73 585
R239 B.n310 B.n309 585
R240 B.n311 B.n72 585
R241 B.n313 B.n312 585
R242 B.n314 B.n71 585
R243 B.n316 B.n315 585
R244 B.n317 B.n70 585
R245 B.n319 B.n318 585
R246 B.n320 B.n69 585
R247 B.n322 B.n321 585
R248 B.n323 B.n68 585
R249 B.n325 B.n324 585
R250 B.n326 B.n67 585
R251 B.n328 B.n327 585
R252 B.n329 B.n66 585
R253 B.n331 B.n330 585
R254 B.n332 B.n65 585
R255 B.n334 B.n333 585
R256 B.n335 B.n64 585
R257 B.n337 B.n336 585
R258 B.n338 B.n63 585
R259 B.n340 B.n339 585
R260 B.n341 B.n62 585
R261 B.n343 B.n342 585
R262 B.n344 B.n61 585
R263 B.n346 B.n345 585
R264 B.n347 B.n60 585
R265 B.n349 B.n348 585
R266 B.n350 B.n59 585
R267 B.n352 B.n351 585
R268 B.n353 B.n58 585
R269 B.n355 B.n354 585
R270 B.n356 B.n57 585
R271 B.n358 B.n357 585
R272 B.n359 B.n56 585
R273 B.n361 B.n360 585
R274 B.n362 B.n55 585
R275 B.n364 B.n363 585
R276 B.n365 B.n54 585
R277 B.n367 B.n366 585
R278 B.n368 B.n53 585
R279 B.n370 B.n369 585
R280 B.n371 B.n52 585
R281 B.n373 B.n372 585
R282 B.n374 B.n51 585
R283 B.n376 B.n375 585
R284 B.n377 B.n50 585
R285 B.n379 B.n378 585
R286 B.n380 B.n49 585
R287 B.n382 B.n381 585
R288 B.n383 B.n48 585
R289 B.n385 B.n384 585
R290 B.n386 B.n47 585
R291 B.n388 B.n387 585
R292 B.n389 B.n46 585
R293 B.n391 B.n390 585
R294 B.n392 B.n45 585
R295 B.n437 B.n436 585
R296 B.n435 B.n26 585
R297 B.n434 B.n433 585
R298 B.n432 B.n27 585
R299 B.n431 B.n430 585
R300 B.n429 B.n28 585
R301 B.n428 B.n427 585
R302 B.n426 B.n29 585
R303 B.n425 B.n424 585
R304 B.n423 B.n30 585
R305 B.n422 B.n421 585
R306 B.n420 B.n31 585
R307 B.n419 B.n418 585
R308 B.n417 B.n35 585
R309 B.n416 B.n415 585
R310 B.n414 B.n36 585
R311 B.n413 B.n412 585
R312 B.n411 B.n37 585
R313 B.n410 B.n409 585
R314 B.n407 B.n38 585
R315 B.n406 B.n405 585
R316 B.n404 B.n41 585
R317 B.n403 B.n402 585
R318 B.n401 B.n42 585
R319 B.n400 B.n399 585
R320 B.n398 B.n43 585
R321 B.n397 B.n396 585
R322 B.n395 B.n44 585
R323 B.n394 B.n393 585
R324 B.n438 B.n25 585
R325 B.n440 B.n439 585
R326 B.n441 B.n24 585
R327 B.n443 B.n442 585
R328 B.n444 B.n23 585
R329 B.n446 B.n445 585
R330 B.n447 B.n22 585
R331 B.n449 B.n448 585
R332 B.n450 B.n21 585
R333 B.n452 B.n451 585
R334 B.n453 B.n20 585
R335 B.n455 B.n454 585
R336 B.n456 B.n19 585
R337 B.n458 B.n457 585
R338 B.n459 B.n18 585
R339 B.n461 B.n460 585
R340 B.n462 B.n17 585
R341 B.n464 B.n463 585
R342 B.n465 B.n16 585
R343 B.n467 B.n466 585
R344 B.n468 B.n15 585
R345 B.n470 B.n469 585
R346 B.n471 B.n14 585
R347 B.n473 B.n472 585
R348 B.n474 B.n13 585
R349 B.n476 B.n475 585
R350 B.n477 B.n12 585
R351 B.n479 B.n478 585
R352 B.n480 B.n11 585
R353 B.n482 B.n481 585
R354 B.n483 B.n10 585
R355 B.n485 B.n484 585
R356 B.n486 B.n9 585
R357 B.n488 B.n487 585
R358 B.n489 B.n8 585
R359 B.n491 B.n490 585
R360 B.n492 B.n7 585
R361 B.n494 B.n493 585
R362 B.n495 B.n6 585
R363 B.n497 B.n496 585
R364 B.n498 B.n5 585
R365 B.n500 B.n499 585
R366 B.n501 B.n4 585
R367 B.n503 B.n502 585
R368 B.n504 B.n3 585
R369 B.n506 B.n505 585
R370 B.n507 B.n0 585
R371 B.n2 B.n1 585
R372 B.n135 B.n134 585
R373 B.n137 B.n136 585
R374 B.n138 B.n133 585
R375 B.n140 B.n139 585
R376 B.n141 B.n132 585
R377 B.n143 B.n142 585
R378 B.n144 B.n131 585
R379 B.n146 B.n145 585
R380 B.n147 B.n130 585
R381 B.n149 B.n148 585
R382 B.n150 B.n129 585
R383 B.n152 B.n151 585
R384 B.n153 B.n128 585
R385 B.n155 B.n154 585
R386 B.n156 B.n127 585
R387 B.n158 B.n157 585
R388 B.n159 B.n126 585
R389 B.n161 B.n160 585
R390 B.n162 B.n125 585
R391 B.n164 B.n163 585
R392 B.n165 B.n124 585
R393 B.n167 B.n166 585
R394 B.n168 B.n123 585
R395 B.n170 B.n169 585
R396 B.n171 B.n122 585
R397 B.n173 B.n172 585
R398 B.n174 B.n121 585
R399 B.n176 B.n175 585
R400 B.n177 B.n120 585
R401 B.n179 B.n178 585
R402 B.n180 B.n119 585
R403 B.n182 B.n181 585
R404 B.n183 B.n118 585
R405 B.n185 B.n184 585
R406 B.n186 B.n117 585
R407 B.n188 B.n187 585
R408 B.n189 B.n116 585
R409 B.n191 B.n190 585
R410 B.n192 B.n115 585
R411 B.n194 B.n193 585
R412 B.n195 B.n114 585
R413 B.n197 B.n196 585
R414 B.n198 B.n113 585
R415 B.n200 B.n199 585
R416 B.n201 B.n112 585
R417 B.n203 B.n202 585
R418 B.n204 B.n203 492.5
R419 B.n249 B.n248 492.5
R420 B.n393 B.n392 492.5
R421 B.n436 B.n25 492.5
R422 B.n105 B.t4 429.272
R423 B.n99 B.t1 429.272
R424 B.n39 B.t8 429.272
R425 B.n32 B.t11 429.272
R426 B.n106 B.t5 364.497
R427 B.n100 B.t2 364.497
R428 B.n40 B.t7 364.497
R429 B.n33 B.t10 364.497
R430 B.n509 B.n508 256.663
R431 B.n508 B.n507 235.042
R432 B.n508 B.n2 235.042
R433 B.n105 B.t3 209.284
R434 B.n99 B.t0 209.284
R435 B.n39 B.t6 209.284
R436 B.n32 B.t9 209.284
R437 B.n205 B.n204 163.367
R438 B.n205 B.n110 163.367
R439 B.n209 B.n110 163.367
R440 B.n210 B.n209 163.367
R441 B.n211 B.n210 163.367
R442 B.n211 B.n108 163.367
R443 B.n215 B.n108 163.367
R444 B.n216 B.n215 163.367
R445 B.n217 B.n216 163.367
R446 B.n217 B.n104 163.367
R447 B.n222 B.n104 163.367
R448 B.n223 B.n222 163.367
R449 B.n224 B.n223 163.367
R450 B.n224 B.n102 163.367
R451 B.n228 B.n102 163.367
R452 B.n229 B.n228 163.367
R453 B.n230 B.n229 163.367
R454 B.n230 B.n98 163.367
R455 B.n235 B.n98 163.367
R456 B.n236 B.n235 163.367
R457 B.n237 B.n236 163.367
R458 B.n237 B.n96 163.367
R459 B.n241 B.n96 163.367
R460 B.n242 B.n241 163.367
R461 B.n243 B.n242 163.367
R462 B.n243 B.n94 163.367
R463 B.n247 B.n94 163.367
R464 B.n248 B.n247 163.367
R465 B.n392 B.n391 163.367
R466 B.n391 B.n46 163.367
R467 B.n387 B.n46 163.367
R468 B.n387 B.n386 163.367
R469 B.n386 B.n385 163.367
R470 B.n385 B.n48 163.367
R471 B.n381 B.n48 163.367
R472 B.n381 B.n380 163.367
R473 B.n380 B.n379 163.367
R474 B.n379 B.n50 163.367
R475 B.n375 B.n50 163.367
R476 B.n375 B.n374 163.367
R477 B.n374 B.n373 163.367
R478 B.n373 B.n52 163.367
R479 B.n369 B.n52 163.367
R480 B.n369 B.n368 163.367
R481 B.n368 B.n367 163.367
R482 B.n367 B.n54 163.367
R483 B.n363 B.n54 163.367
R484 B.n363 B.n362 163.367
R485 B.n362 B.n361 163.367
R486 B.n361 B.n56 163.367
R487 B.n357 B.n56 163.367
R488 B.n357 B.n356 163.367
R489 B.n356 B.n355 163.367
R490 B.n355 B.n58 163.367
R491 B.n351 B.n58 163.367
R492 B.n351 B.n350 163.367
R493 B.n350 B.n349 163.367
R494 B.n349 B.n60 163.367
R495 B.n345 B.n60 163.367
R496 B.n345 B.n344 163.367
R497 B.n344 B.n343 163.367
R498 B.n343 B.n62 163.367
R499 B.n339 B.n62 163.367
R500 B.n339 B.n338 163.367
R501 B.n338 B.n337 163.367
R502 B.n337 B.n64 163.367
R503 B.n333 B.n64 163.367
R504 B.n333 B.n332 163.367
R505 B.n332 B.n331 163.367
R506 B.n331 B.n66 163.367
R507 B.n327 B.n66 163.367
R508 B.n327 B.n326 163.367
R509 B.n326 B.n325 163.367
R510 B.n325 B.n68 163.367
R511 B.n321 B.n68 163.367
R512 B.n321 B.n320 163.367
R513 B.n320 B.n319 163.367
R514 B.n319 B.n70 163.367
R515 B.n315 B.n70 163.367
R516 B.n315 B.n314 163.367
R517 B.n314 B.n313 163.367
R518 B.n313 B.n72 163.367
R519 B.n309 B.n72 163.367
R520 B.n309 B.n308 163.367
R521 B.n308 B.n307 163.367
R522 B.n307 B.n74 163.367
R523 B.n303 B.n74 163.367
R524 B.n303 B.n302 163.367
R525 B.n302 B.n301 163.367
R526 B.n301 B.n76 163.367
R527 B.n297 B.n76 163.367
R528 B.n297 B.n296 163.367
R529 B.n296 B.n295 163.367
R530 B.n295 B.n78 163.367
R531 B.n291 B.n78 163.367
R532 B.n291 B.n290 163.367
R533 B.n290 B.n289 163.367
R534 B.n289 B.n80 163.367
R535 B.n285 B.n80 163.367
R536 B.n285 B.n284 163.367
R537 B.n284 B.n283 163.367
R538 B.n283 B.n82 163.367
R539 B.n279 B.n82 163.367
R540 B.n279 B.n278 163.367
R541 B.n278 B.n277 163.367
R542 B.n277 B.n84 163.367
R543 B.n273 B.n84 163.367
R544 B.n273 B.n272 163.367
R545 B.n272 B.n271 163.367
R546 B.n271 B.n86 163.367
R547 B.n267 B.n86 163.367
R548 B.n267 B.n266 163.367
R549 B.n266 B.n265 163.367
R550 B.n265 B.n88 163.367
R551 B.n261 B.n88 163.367
R552 B.n261 B.n260 163.367
R553 B.n260 B.n259 163.367
R554 B.n259 B.n90 163.367
R555 B.n255 B.n90 163.367
R556 B.n255 B.n254 163.367
R557 B.n254 B.n253 163.367
R558 B.n253 B.n92 163.367
R559 B.n249 B.n92 163.367
R560 B.n436 B.n435 163.367
R561 B.n435 B.n434 163.367
R562 B.n434 B.n27 163.367
R563 B.n430 B.n27 163.367
R564 B.n430 B.n429 163.367
R565 B.n429 B.n428 163.367
R566 B.n428 B.n29 163.367
R567 B.n424 B.n29 163.367
R568 B.n424 B.n423 163.367
R569 B.n423 B.n422 163.367
R570 B.n422 B.n31 163.367
R571 B.n418 B.n31 163.367
R572 B.n418 B.n417 163.367
R573 B.n417 B.n416 163.367
R574 B.n416 B.n36 163.367
R575 B.n412 B.n36 163.367
R576 B.n412 B.n411 163.367
R577 B.n411 B.n410 163.367
R578 B.n410 B.n38 163.367
R579 B.n405 B.n38 163.367
R580 B.n405 B.n404 163.367
R581 B.n404 B.n403 163.367
R582 B.n403 B.n42 163.367
R583 B.n399 B.n42 163.367
R584 B.n399 B.n398 163.367
R585 B.n398 B.n397 163.367
R586 B.n397 B.n44 163.367
R587 B.n393 B.n44 163.367
R588 B.n440 B.n25 163.367
R589 B.n441 B.n440 163.367
R590 B.n442 B.n441 163.367
R591 B.n442 B.n23 163.367
R592 B.n446 B.n23 163.367
R593 B.n447 B.n446 163.367
R594 B.n448 B.n447 163.367
R595 B.n448 B.n21 163.367
R596 B.n452 B.n21 163.367
R597 B.n453 B.n452 163.367
R598 B.n454 B.n453 163.367
R599 B.n454 B.n19 163.367
R600 B.n458 B.n19 163.367
R601 B.n459 B.n458 163.367
R602 B.n460 B.n459 163.367
R603 B.n460 B.n17 163.367
R604 B.n464 B.n17 163.367
R605 B.n465 B.n464 163.367
R606 B.n466 B.n465 163.367
R607 B.n466 B.n15 163.367
R608 B.n470 B.n15 163.367
R609 B.n471 B.n470 163.367
R610 B.n472 B.n471 163.367
R611 B.n472 B.n13 163.367
R612 B.n476 B.n13 163.367
R613 B.n477 B.n476 163.367
R614 B.n478 B.n477 163.367
R615 B.n478 B.n11 163.367
R616 B.n482 B.n11 163.367
R617 B.n483 B.n482 163.367
R618 B.n484 B.n483 163.367
R619 B.n484 B.n9 163.367
R620 B.n488 B.n9 163.367
R621 B.n489 B.n488 163.367
R622 B.n490 B.n489 163.367
R623 B.n490 B.n7 163.367
R624 B.n494 B.n7 163.367
R625 B.n495 B.n494 163.367
R626 B.n496 B.n495 163.367
R627 B.n496 B.n5 163.367
R628 B.n500 B.n5 163.367
R629 B.n501 B.n500 163.367
R630 B.n502 B.n501 163.367
R631 B.n502 B.n3 163.367
R632 B.n506 B.n3 163.367
R633 B.n507 B.n506 163.367
R634 B.n134 B.n2 163.367
R635 B.n137 B.n134 163.367
R636 B.n138 B.n137 163.367
R637 B.n139 B.n138 163.367
R638 B.n139 B.n132 163.367
R639 B.n143 B.n132 163.367
R640 B.n144 B.n143 163.367
R641 B.n145 B.n144 163.367
R642 B.n145 B.n130 163.367
R643 B.n149 B.n130 163.367
R644 B.n150 B.n149 163.367
R645 B.n151 B.n150 163.367
R646 B.n151 B.n128 163.367
R647 B.n155 B.n128 163.367
R648 B.n156 B.n155 163.367
R649 B.n157 B.n156 163.367
R650 B.n157 B.n126 163.367
R651 B.n161 B.n126 163.367
R652 B.n162 B.n161 163.367
R653 B.n163 B.n162 163.367
R654 B.n163 B.n124 163.367
R655 B.n167 B.n124 163.367
R656 B.n168 B.n167 163.367
R657 B.n169 B.n168 163.367
R658 B.n169 B.n122 163.367
R659 B.n173 B.n122 163.367
R660 B.n174 B.n173 163.367
R661 B.n175 B.n174 163.367
R662 B.n175 B.n120 163.367
R663 B.n179 B.n120 163.367
R664 B.n180 B.n179 163.367
R665 B.n181 B.n180 163.367
R666 B.n181 B.n118 163.367
R667 B.n185 B.n118 163.367
R668 B.n186 B.n185 163.367
R669 B.n187 B.n186 163.367
R670 B.n187 B.n116 163.367
R671 B.n191 B.n116 163.367
R672 B.n192 B.n191 163.367
R673 B.n193 B.n192 163.367
R674 B.n193 B.n114 163.367
R675 B.n197 B.n114 163.367
R676 B.n198 B.n197 163.367
R677 B.n199 B.n198 163.367
R678 B.n199 B.n112 163.367
R679 B.n203 B.n112 163.367
R680 B.n106 B.n105 64.7763
R681 B.n100 B.n99 64.7763
R682 B.n40 B.n39 64.7763
R683 B.n33 B.n32 64.7763
R684 B.n219 B.n106 59.5399
R685 B.n233 B.n100 59.5399
R686 B.n408 B.n40 59.5399
R687 B.n34 B.n33 59.5399
R688 B.n438 B.n437 32.0005
R689 B.n394 B.n45 32.0005
R690 B.n250 B.n93 32.0005
R691 B.n202 B.n111 32.0005
R692 B B.n509 18.0485
R693 B.n439 B.n438 10.6151
R694 B.n439 B.n24 10.6151
R695 B.n443 B.n24 10.6151
R696 B.n444 B.n443 10.6151
R697 B.n445 B.n444 10.6151
R698 B.n445 B.n22 10.6151
R699 B.n449 B.n22 10.6151
R700 B.n450 B.n449 10.6151
R701 B.n451 B.n450 10.6151
R702 B.n451 B.n20 10.6151
R703 B.n455 B.n20 10.6151
R704 B.n456 B.n455 10.6151
R705 B.n457 B.n456 10.6151
R706 B.n457 B.n18 10.6151
R707 B.n461 B.n18 10.6151
R708 B.n462 B.n461 10.6151
R709 B.n463 B.n462 10.6151
R710 B.n463 B.n16 10.6151
R711 B.n467 B.n16 10.6151
R712 B.n468 B.n467 10.6151
R713 B.n469 B.n468 10.6151
R714 B.n469 B.n14 10.6151
R715 B.n473 B.n14 10.6151
R716 B.n474 B.n473 10.6151
R717 B.n475 B.n474 10.6151
R718 B.n475 B.n12 10.6151
R719 B.n479 B.n12 10.6151
R720 B.n480 B.n479 10.6151
R721 B.n481 B.n480 10.6151
R722 B.n481 B.n10 10.6151
R723 B.n485 B.n10 10.6151
R724 B.n486 B.n485 10.6151
R725 B.n487 B.n486 10.6151
R726 B.n487 B.n8 10.6151
R727 B.n491 B.n8 10.6151
R728 B.n492 B.n491 10.6151
R729 B.n493 B.n492 10.6151
R730 B.n493 B.n6 10.6151
R731 B.n497 B.n6 10.6151
R732 B.n498 B.n497 10.6151
R733 B.n499 B.n498 10.6151
R734 B.n499 B.n4 10.6151
R735 B.n503 B.n4 10.6151
R736 B.n504 B.n503 10.6151
R737 B.n505 B.n504 10.6151
R738 B.n505 B.n0 10.6151
R739 B.n437 B.n26 10.6151
R740 B.n433 B.n26 10.6151
R741 B.n433 B.n432 10.6151
R742 B.n432 B.n431 10.6151
R743 B.n431 B.n28 10.6151
R744 B.n427 B.n28 10.6151
R745 B.n427 B.n426 10.6151
R746 B.n426 B.n425 10.6151
R747 B.n425 B.n30 10.6151
R748 B.n421 B.n420 10.6151
R749 B.n420 B.n419 10.6151
R750 B.n419 B.n35 10.6151
R751 B.n415 B.n35 10.6151
R752 B.n415 B.n414 10.6151
R753 B.n414 B.n413 10.6151
R754 B.n413 B.n37 10.6151
R755 B.n409 B.n37 10.6151
R756 B.n407 B.n406 10.6151
R757 B.n406 B.n41 10.6151
R758 B.n402 B.n41 10.6151
R759 B.n402 B.n401 10.6151
R760 B.n401 B.n400 10.6151
R761 B.n400 B.n43 10.6151
R762 B.n396 B.n43 10.6151
R763 B.n396 B.n395 10.6151
R764 B.n395 B.n394 10.6151
R765 B.n390 B.n45 10.6151
R766 B.n390 B.n389 10.6151
R767 B.n389 B.n388 10.6151
R768 B.n388 B.n47 10.6151
R769 B.n384 B.n47 10.6151
R770 B.n384 B.n383 10.6151
R771 B.n383 B.n382 10.6151
R772 B.n382 B.n49 10.6151
R773 B.n378 B.n49 10.6151
R774 B.n378 B.n377 10.6151
R775 B.n377 B.n376 10.6151
R776 B.n376 B.n51 10.6151
R777 B.n372 B.n51 10.6151
R778 B.n372 B.n371 10.6151
R779 B.n371 B.n370 10.6151
R780 B.n370 B.n53 10.6151
R781 B.n366 B.n53 10.6151
R782 B.n366 B.n365 10.6151
R783 B.n365 B.n364 10.6151
R784 B.n364 B.n55 10.6151
R785 B.n360 B.n55 10.6151
R786 B.n360 B.n359 10.6151
R787 B.n359 B.n358 10.6151
R788 B.n358 B.n57 10.6151
R789 B.n354 B.n57 10.6151
R790 B.n354 B.n353 10.6151
R791 B.n353 B.n352 10.6151
R792 B.n352 B.n59 10.6151
R793 B.n348 B.n59 10.6151
R794 B.n348 B.n347 10.6151
R795 B.n347 B.n346 10.6151
R796 B.n346 B.n61 10.6151
R797 B.n342 B.n61 10.6151
R798 B.n342 B.n341 10.6151
R799 B.n341 B.n340 10.6151
R800 B.n340 B.n63 10.6151
R801 B.n336 B.n63 10.6151
R802 B.n336 B.n335 10.6151
R803 B.n335 B.n334 10.6151
R804 B.n334 B.n65 10.6151
R805 B.n330 B.n65 10.6151
R806 B.n330 B.n329 10.6151
R807 B.n329 B.n328 10.6151
R808 B.n328 B.n67 10.6151
R809 B.n324 B.n67 10.6151
R810 B.n324 B.n323 10.6151
R811 B.n323 B.n322 10.6151
R812 B.n322 B.n69 10.6151
R813 B.n318 B.n69 10.6151
R814 B.n318 B.n317 10.6151
R815 B.n317 B.n316 10.6151
R816 B.n316 B.n71 10.6151
R817 B.n312 B.n71 10.6151
R818 B.n312 B.n311 10.6151
R819 B.n311 B.n310 10.6151
R820 B.n310 B.n73 10.6151
R821 B.n306 B.n73 10.6151
R822 B.n306 B.n305 10.6151
R823 B.n305 B.n304 10.6151
R824 B.n304 B.n75 10.6151
R825 B.n300 B.n75 10.6151
R826 B.n300 B.n299 10.6151
R827 B.n299 B.n298 10.6151
R828 B.n298 B.n77 10.6151
R829 B.n294 B.n77 10.6151
R830 B.n294 B.n293 10.6151
R831 B.n293 B.n292 10.6151
R832 B.n292 B.n79 10.6151
R833 B.n288 B.n79 10.6151
R834 B.n288 B.n287 10.6151
R835 B.n287 B.n286 10.6151
R836 B.n286 B.n81 10.6151
R837 B.n282 B.n81 10.6151
R838 B.n282 B.n281 10.6151
R839 B.n281 B.n280 10.6151
R840 B.n280 B.n83 10.6151
R841 B.n276 B.n83 10.6151
R842 B.n276 B.n275 10.6151
R843 B.n275 B.n274 10.6151
R844 B.n274 B.n85 10.6151
R845 B.n270 B.n85 10.6151
R846 B.n270 B.n269 10.6151
R847 B.n269 B.n268 10.6151
R848 B.n268 B.n87 10.6151
R849 B.n264 B.n87 10.6151
R850 B.n264 B.n263 10.6151
R851 B.n263 B.n262 10.6151
R852 B.n262 B.n89 10.6151
R853 B.n258 B.n89 10.6151
R854 B.n258 B.n257 10.6151
R855 B.n257 B.n256 10.6151
R856 B.n256 B.n91 10.6151
R857 B.n252 B.n91 10.6151
R858 B.n252 B.n251 10.6151
R859 B.n251 B.n250 10.6151
R860 B.n135 B.n1 10.6151
R861 B.n136 B.n135 10.6151
R862 B.n136 B.n133 10.6151
R863 B.n140 B.n133 10.6151
R864 B.n141 B.n140 10.6151
R865 B.n142 B.n141 10.6151
R866 B.n142 B.n131 10.6151
R867 B.n146 B.n131 10.6151
R868 B.n147 B.n146 10.6151
R869 B.n148 B.n147 10.6151
R870 B.n148 B.n129 10.6151
R871 B.n152 B.n129 10.6151
R872 B.n153 B.n152 10.6151
R873 B.n154 B.n153 10.6151
R874 B.n154 B.n127 10.6151
R875 B.n158 B.n127 10.6151
R876 B.n159 B.n158 10.6151
R877 B.n160 B.n159 10.6151
R878 B.n160 B.n125 10.6151
R879 B.n164 B.n125 10.6151
R880 B.n165 B.n164 10.6151
R881 B.n166 B.n165 10.6151
R882 B.n166 B.n123 10.6151
R883 B.n170 B.n123 10.6151
R884 B.n171 B.n170 10.6151
R885 B.n172 B.n171 10.6151
R886 B.n172 B.n121 10.6151
R887 B.n176 B.n121 10.6151
R888 B.n177 B.n176 10.6151
R889 B.n178 B.n177 10.6151
R890 B.n178 B.n119 10.6151
R891 B.n182 B.n119 10.6151
R892 B.n183 B.n182 10.6151
R893 B.n184 B.n183 10.6151
R894 B.n184 B.n117 10.6151
R895 B.n188 B.n117 10.6151
R896 B.n189 B.n188 10.6151
R897 B.n190 B.n189 10.6151
R898 B.n190 B.n115 10.6151
R899 B.n194 B.n115 10.6151
R900 B.n195 B.n194 10.6151
R901 B.n196 B.n195 10.6151
R902 B.n196 B.n113 10.6151
R903 B.n200 B.n113 10.6151
R904 B.n201 B.n200 10.6151
R905 B.n202 B.n201 10.6151
R906 B.n206 B.n111 10.6151
R907 B.n207 B.n206 10.6151
R908 B.n208 B.n207 10.6151
R909 B.n208 B.n109 10.6151
R910 B.n212 B.n109 10.6151
R911 B.n213 B.n212 10.6151
R912 B.n214 B.n213 10.6151
R913 B.n214 B.n107 10.6151
R914 B.n218 B.n107 10.6151
R915 B.n221 B.n220 10.6151
R916 B.n221 B.n103 10.6151
R917 B.n225 B.n103 10.6151
R918 B.n226 B.n225 10.6151
R919 B.n227 B.n226 10.6151
R920 B.n227 B.n101 10.6151
R921 B.n231 B.n101 10.6151
R922 B.n232 B.n231 10.6151
R923 B.n234 B.n97 10.6151
R924 B.n238 B.n97 10.6151
R925 B.n239 B.n238 10.6151
R926 B.n240 B.n239 10.6151
R927 B.n240 B.n95 10.6151
R928 B.n244 B.n95 10.6151
R929 B.n245 B.n244 10.6151
R930 B.n246 B.n245 10.6151
R931 B.n246 B.n93 10.6151
R932 B.n509 B.n0 8.11757
R933 B.n509 B.n1 8.11757
R934 B.n421 B.n34 6.5566
R935 B.n409 B.n408 6.5566
R936 B.n220 B.n219 6.5566
R937 B.n233 B.n232 6.5566
R938 B.n34 B.n30 4.05904
R939 B.n408 B.n407 4.05904
R940 B.n219 B.n218 4.05904
R941 B.n234 B.n233 4.05904
C0 B VN 1.0873f
C1 VDD2 VN 1.03129f
C2 VP VN 5.33266f
C3 B VDD2 1.42053f
C4 VP B 1.87628f
C5 VP VDD2 0.501648f
C6 w_n3642_n1202# VN 6.81738f
C7 w_n3642_n1202# B 7.28439f
C8 VDD1 VN 0.158984f
C9 w_n3642_n1202# VDD2 1.73326f
C10 B VDD1 1.33598f
C11 VP w_n3642_n1202# 7.28221f
C12 VDD1 VDD2 1.56642f
C13 VP VDD1 1.37052f
C14 w_n3642_n1202# VDD1 1.63611f
C15 VTAIL VN 2.14321f
C16 B VTAIL 1.19734f
C17 VDD2 VTAIL 4.16242f
C18 VP VTAIL 2.15733f
C19 w_n3642_n1202# VTAIL 1.44949f
C20 VDD1 VTAIL 4.10627f
C21 VDD2 VSUBS 1.118239f
C22 VDD1 VSUBS 1.591173f
C23 VTAIL VSUBS 0.580184f
C24 VN VSUBS 6.44243f
C25 VP VSUBS 2.657369f
C26 B VSUBS 3.873923f
C27 w_n3642_n1202# VSUBS 56.3345f
C28 B.n0 VSUBS 0.008851f
C29 B.n1 VSUBS 0.008851f
C30 B.n2 VSUBS 0.01309f
C31 B.n3 VSUBS 0.010031f
C32 B.n4 VSUBS 0.010031f
C33 B.n5 VSUBS 0.010031f
C34 B.n6 VSUBS 0.010031f
C35 B.n7 VSUBS 0.010031f
C36 B.n8 VSUBS 0.010031f
C37 B.n9 VSUBS 0.010031f
C38 B.n10 VSUBS 0.010031f
C39 B.n11 VSUBS 0.010031f
C40 B.n12 VSUBS 0.010031f
C41 B.n13 VSUBS 0.010031f
C42 B.n14 VSUBS 0.010031f
C43 B.n15 VSUBS 0.010031f
C44 B.n16 VSUBS 0.010031f
C45 B.n17 VSUBS 0.010031f
C46 B.n18 VSUBS 0.010031f
C47 B.n19 VSUBS 0.010031f
C48 B.n20 VSUBS 0.010031f
C49 B.n21 VSUBS 0.010031f
C50 B.n22 VSUBS 0.010031f
C51 B.n23 VSUBS 0.010031f
C52 B.n24 VSUBS 0.010031f
C53 B.n25 VSUBS 0.022733f
C54 B.n26 VSUBS 0.010031f
C55 B.n27 VSUBS 0.010031f
C56 B.n28 VSUBS 0.010031f
C57 B.n29 VSUBS 0.010031f
C58 B.n30 VSUBS 0.006933f
C59 B.n31 VSUBS 0.010031f
C60 B.t10 VSUBS 0.031606f
C61 B.t11 VSUBS 0.040464f
C62 B.t9 VSUBS 0.254747f
C63 B.n32 VSUBS 0.096013f
C64 B.n33 VSUBS 0.073005f
C65 B.n34 VSUBS 0.023242f
C66 B.n35 VSUBS 0.010031f
C67 B.n36 VSUBS 0.010031f
C68 B.n37 VSUBS 0.010031f
C69 B.n38 VSUBS 0.010031f
C70 B.t7 VSUBS 0.031606f
C71 B.t8 VSUBS 0.040464f
C72 B.t6 VSUBS 0.254747f
C73 B.n39 VSUBS 0.096013f
C74 B.n40 VSUBS 0.073005f
C75 B.n41 VSUBS 0.010031f
C76 B.n42 VSUBS 0.010031f
C77 B.n43 VSUBS 0.010031f
C78 B.n44 VSUBS 0.010031f
C79 B.n45 VSUBS 0.022733f
C80 B.n46 VSUBS 0.010031f
C81 B.n47 VSUBS 0.010031f
C82 B.n48 VSUBS 0.010031f
C83 B.n49 VSUBS 0.010031f
C84 B.n50 VSUBS 0.010031f
C85 B.n51 VSUBS 0.010031f
C86 B.n52 VSUBS 0.010031f
C87 B.n53 VSUBS 0.010031f
C88 B.n54 VSUBS 0.010031f
C89 B.n55 VSUBS 0.010031f
C90 B.n56 VSUBS 0.010031f
C91 B.n57 VSUBS 0.010031f
C92 B.n58 VSUBS 0.010031f
C93 B.n59 VSUBS 0.010031f
C94 B.n60 VSUBS 0.010031f
C95 B.n61 VSUBS 0.010031f
C96 B.n62 VSUBS 0.010031f
C97 B.n63 VSUBS 0.010031f
C98 B.n64 VSUBS 0.010031f
C99 B.n65 VSUBS 0.010031f
C100 B.n66 VSUBS 0.010031f
C101 B.n67 VSUBS 0.010031f
C102 B.n68 VSUBS 0.010031f
C103 B.n69 VSUBS 0.010031f
C104 B.n70 VSUBS 0.010031f
C105 B.n71 VSUBS 0.010031f
C106 B.n72 VSUBS 0.010031f
C107 B.n73 VSUBS 0.010031f
C108 B.n74 VSUBS 0.010031f
C109 B.n75 VSUBS 0.010031f
C110 B.n76 VSUBS 0.010031f
C111 B.n77 VSUBS 0.010031f
C112 B.n78 VSUBS 0.010031f
C113 B.n79 VSUBS 0.010031f
C114 B.n80 VSUBS 0.010031f
C115 B.n81 VSUBS 0.010031f
C116 B.n82 VSUBS 0.010031f
C117 B.n83 VSUBS 0.010031f
C118 B.n84 VSUBS 0.010031f
C119 B.n85 VSUBS 0.010031f
C120 B.n86 VSUBS 0.010031f
C121 B.n87 VSUBS 0.010031f
C122 B.n88 VSUBS 0.010031f
C123 B.n89 VSUBS 0.010031f
C124 B.n90 VSUBS 0.010031f
C125 B.n91 VSUBS 0.010031f
C126 B.n92 VSUBS 0.010031f
C127 B.n93 VSUBS 0.022379f
C128 B.n94 VSUBS 0.010031f
C129 B.n95 VSUBS 0.010031f
C130 B.n96 VSUBS 0.010031f
C131 B.n97 VSUBS 0.010031f
C132 B.n98 VSUBS 0.010031f
C133 B.t2 VSUBS 0.031606f
C134 B.t1 VSUBS 0.040464f
C135 B.t0 VSUBS 0.254747f
C136 B.n99 VSUBS 0.096013f
C137 B.n100 VSUBS 0.073005f
C138 B.n101 VSUBS 0.010031f
C139 B.n102 VSUBS 0.010031f
C140 B.n103 VSUBS 0.010031f
C141 B.n104 VSUBS 0.010031f
C142 B.t5 VSUBS 0.031606f
C143 B.t4 VSUBS 0.040464f
C144 B.t3 VSUBS 0.254747f
C145 B.n105 VSUBS 0.096013f
C146 B.n106 VSUBS 0.073005f
C147 B.n107 VSUBS 0.010031f
C148 B.n108 VSUBS 0.010031f
C149 B.n109 VSUBS 0.010031f
C150 B.n110 VSUBS 0.010031f
C151 B.n111 VSUBS 0.023588f
C152 B.n112 VSUBS 0.010031f
C153 B.n113 VSUBS 0.010031f
C154 B.n114 VSUBS 0.010031f
C155 B.n115 VSUBS 0.010031f
C156 B.n116 VSUBS 0.010031f
C157 B.n117 VSUBS 0.010031f
C158 B.n118 VSUBS 0.010031f
C159 B.n119 VSUBS 0.010031f
C160 B.n120 VSUBS 0.010031f
C161 B.n121 VSUBS 0.010031f
C162 B.n122 VSUBS 0.010031f
C163 B.n123 VSUBS 0.010031f
C164 B.n124 VSUBS 0.010031f
C165 B.n125 VSUBS 0.010031f
C166 B.n126 VSUBS 0.010031f
C167 B.n127 VSUBS 0.010031f
C168 B.n128 VSUBS 0.010031f
C169 B.n129 VSUBS 0.010031f
C170 B.n130 VSUBS 0.010031f
C171 B.n131 VSUBS 0.010031f
C172 B.n132 VSUBS 0.010031f
C173 B.n133 VSUBS 0.010031f
C174 B.n134 VSUBS 0.010031f
C175 B.n135 VSUBS 0.010031f
C176 B.n136 VSUBS 0.010031f
C177 B.n137 VSUBS 0.010031f
C178 B.n138 VSUBS 0.010031f
C179 B.n139 VSUBS 0.010031f
C180 B.n140 VSUBS 0.010031f
C181 B.n141 VSUBS 0.010031f
C182 B.n142 VSUBS 0.010031f
C183 B.n143 VSUBS 0.010031f
C184 B.n144 VSUBS 0.010031f
C185 B.n145 VSUBS 0.010031f
C186 B.n146 VSUBS 0.010031f
C187 B.n147 VSUBS 0.010031f
C188 B.n148 VSUBS 0.010031f
C189 B.n149 VSUBS 0.010031f
C190 B.n150 VSUBS 0.010031f
C191 B.n151 VSUBS 0.010031f
C192 B.n152 VSUBS 0.010031f
C193 B.n153 VSUBS 0.010031f
C194 B.n154 VSUBS 0.010031f
C195 B.n155 VSUBS 0.010031f
C196 B.n156 VSUBS 0.010031f
C197 B.n157 VSUBS 0.010031f
C198 B.n158 VSUBS 0.010031f
C199 B.n159 VSUBS 0.010031f
C200 B.n160 VSUBS 0.010031f
C201 B.n161 VSUBS 0.010031f
C202 B.n162 VSUBS 0.010031f
C203 B.n163 VSUBS 0.010031f
C204 B.n164 VSUBS 0.010031f
C205 B.n165 VSUBS 0.010031f
C206 B.n166 VSUBS 0.010031f
C207 B.n167 VSUBS 0.010031f
C208 B.n168 VSUBS 0.010031f
C209 B.n169 VSUBS 0.010031f
C210 B.n170 VSUBS 0.010031f
C211 B.n171 VSUBS 0.010031f
C212 B.n172 VSUBS 0.010031f
C213 B.n173 VSUBS 0.010031f
C214 B.n174 VSUBS 0.010031f
C215 B.n175 VSUBS 0.010031f
C216 B.n176 VSUBS 0.010031f
C217 B.n177 VSUBS 0.010031f
C218 B.n178 VSUBS 0.010031f
C219 B.n179 VSUBS 0.010031f
C220 B.n180 VSUBS 0.010031f
C221 B.n181 VSUBS 0.010031f
C222 B.n182 VSUBS 0.010031f
C223 B.n183 VSUBS 0.010031f
C224 B.n184 VSUBS 0.010031f
C225 B.n185 VSUBS 0.010031f
C226 B.n186 VSUBS 0.010031f
C227 B.n187 VSUBS 0.010031f
C228 B.n188 VSUBS 0.010031f
C229 B.n189 VSUBS 0.010031f
C230 B.n190 VSUBS 0.010031f
C231 B.n191 VSUBS 0.010031f
C232 B.n192 VSUBS 0.010031f
C233 B.n193 VSUBS 0.010031f
C234 B.n194 VSUBS 0.010031f
C235 B.n195 VSUBS 0.010031f
C236 B.n196 VSUBS 0.010031f
C237 B.n197 VSUBS 0.010031f
C238 B.n198 VSUBS 0.010031f
C239 B.n199 VSUBS 0.010031f
C240 B.n200 VSUBS 0.010031f
C241 B.n201 VSUBS 0.010031f
C242 B.n202 VSUBS 0.022733f
C243 B.n203 VSUBS 0.022733f
C244 B.n204 VSUBS 0.023588f
C245 B.n205 VSUBS 0.010031f
C246 B.n206 VSUBS 0.010031f
C247 B.n207 VSUBS 0.010031f
C248 B.n208 VSUBS 0.010031f
C249 B.n209 VSUBS 0.010031f
C250 B.n210 VSUBS 0.010031f
C251 B.n211 VSUBS 0.010031f
C252 B.n212 VSUBS 0.010031f
C253 B.n213 VSUBS 0.010031f
C254 B.n214 VSUBS 0.010031f
C255 B.n215 VSUBS 0.010031f
C256 B.n216 VSUBS 0.010031f
C257 B.n217 VSUBS 0.010031f
C258 B.n218 VSUBS 0.006933f
C259 B.n219 VSUBS 0.023242f
C260 B.n220 VSUBS 0.008114f
C261 B.n221 VSUBS 0.010031f
C262 B.n222 VSUBS 0.010031f
C263 B.n223 VSUBS 0.010031f
C264 B.n224 VSUBS 0.010031f
C265 B.n225 VSUBS 0.010031f
C266 B.n226 VSUBS 0.010031f
C267 B.n227 VSUBS 0.010031f
C268 B.n228 VSUBS 0.010031f
C269 B.n229 VSUBS 0.010031f
C270 B.n230 VSUBS 0.010031f
C271 B.n231 VSUBS 0.010031f
C272 B.n232 VSUBS 0.008114f
C273 B.n233 VSUBS 0.023242f
C274 B.n234 VSUBS 0.006933f
C275 B.n235 VSUBS 0.010031f
C276 B.n236 VSUBS 0.010031f
C277 B.n237 VSUBS 0.010031f
C278 B.n238 VSUBS 0.010031f
C279 B.n239 VSUBS 0.010031f
C280 B.n240 VSUBS 0.010031f
C281 B.n241 VSUBS 0.010031f
C282 B.n242 VSUBS 0.010031f
C283 B.n243 VSUBS 0.010031f
C284 B.n244 VSUBS 0.010031f
C285 B.n245 VSUBS 0.010031f
C286 B.n246 VSUBS 0.010031f
C287 B.n247 VSUBS 0.010031f
C288 B.n248 VSUBS 0.023588f
C289 B.n249 VSUBS 0.022733f
C290 B.n250 VSUBS 0.023943f
C291 B.n251 VSUBS 0.010031f
C292 B.n252 VSUBS 0.010031f
C293 B.n253 VSUBS 0.010031f
C294 B.n254 VSUBS 0.010031f
C295 B.n255 VSUBS 0.010031f
C296 B.n256 VSUBS 0.010031f
C297 B.n257 VSUBS 0.010031f
C298 B.n258 VSUBS 0.010031f
C299 B.n259 VSUBS 0.010031f
C300 B.n260 VSUBS 0.010031f
C301 B.n261 VSUBS 0.010031f
C302 B.n262 VSUBS 0.010031f
C303 B.n263 VSUBS 0.010031f
C304 B.n264 VSUBS 0.010031f
C305 B.n265 VSUBS 0.010031f
C306 B.n266 VSUBS 0.010031f
C307 B.n267 VSUBS 0.010031f
C308 B.n268 VSUBS 0.010031f
C309 B.n269 VSUBS 0.010031f
C310 B.n270 VSUBS 0.010031f
C311 B.n271 VSUBS 0.010031f
C312 B.n272 VSUBS 0.010031f
C313 B.n273 VSUBS 0.010031f
C314 B.n274 VSUBS 0.010031f
C315 B.n275 VSUBS 0.010031f
C316 B.n276 VSUBS 0.010031f
C317 B.n277 VSUBS 0.010031f
C318 B.n278 VSUBS 0.010031f
C319 B.n279 VSUBS 0.010031f
C320 B.n280 VSUBS 0.010031f
C321 B.n281 VSUBS 0.010031f
C322 B.n282 VSUBS 0.010031f
C323 B.n283 VSUBS 0.010031f
C324 B.n284 VSUBS 0.010031f
C325 B.n285 VSUBS 0.010031f
C326 B.n286 VSUBS 0.010031f
C327 B.n287 VSUBS 0.010031f
C328 B.n288 VSUBS 0.010031f
C329 B.n289 VSUBS 0.010031f
C330 B.n290 VSUBS 0.010031f
C331 B.n291 VSUBS 0.010031f
C332 B.n292 VSUBS 0.010031f
C333 B.n293 VSUBS 0.010031f
C334 B.n294 VSUBS 0.010031f
C335 B.n295 VSUBS 0.010031f
C336 B.n296 VSUBS 0.010031f
C337 B.n297 VSUBS 0.010031f
C338 B.n298 VSUBS 0.010031f
C339 B.n299 VSUBS 0.010031f
C340 B.n300 VSUBS 0.010031f
C341 B.n301 VSUBS 0.010031f
C342 B.n302 VSUBS 0.010031f
C343 B.n303 VSUBS 0.010031f
C344 B.n304 VSUBS 0.010031f
C345 B.n305 VSUBS 0.010031f
C346 B.n306 VSUBS 0.010031f
C347 B.n307 VSUBS 0.010031f
C348 B.n308 VSUBS 0.010031f
C349 B.n309 VSUBS 0.010031f
C350 B.n310 VSUBS 0.010031f
C351 B.n311 VSUBS 0.010031f
C352 B.n312 VSUBS 0.010031f
C353 B.n313 VSUBS 0.010031f
C354 B.n314 VSUBS 0.010031f
C355 B.n315 VSUBS 0.010031f
C356 B.n316 VSUBS 0.010031f
C357 B.n317 VSUBS 0.010031f
C358 B.n318 VSUBS 0.010031f
C359 B.n319 VSUBS 0.010031f
C360 B.n320 VSUBS 0.010031f
C361 B.n321 VSUBS 0.010031f
C362 B.n322 VSUBS 0.010031f
C363 B.n323 VSUBS 0.010031f
C364 B.n324 VSUBS 0.010031f
C365 B.n325 VSUBS 0.010031f
C366 B.n326 VSUBS 0.010031f
C367 B.n327 VSUBS 0.010031f
C368 B.n328 VSUBS 0.010031f
C369 B.n329 VSUBS 0.010031f
C370 B.n330 VSUBS 0.010031f
C371 B.n331 VSUBS 0.010031f
C372 B.n332 VSUBS 0.010031f
C373 B.n333 VSUBS 0.010031f
C374 B.n334 VSUBS 0.010031f
C375 B.n335 VSUBS 0.010031f
C376 B.n336 VSUBS 0.010031f
C377 B.n337 VSUBS 0.010031f
C378 B.n338 VSUBS 0.010031f
C379 B.n339 VSUBS 0.010031f
C380 B.n340 VSUBS 0.010031f
C381 B.n341 VSUBS 0.010031f
C382 B.n342 VSUBS 0.010031f
C383 B.n343 VSUBS 0.010031f
C384 B.n344 VSUBS 0.010031f
C385 B.n345 VSUBS 0.010031f
C386 B.n346 VSUBS 0.010031f
C387 B.n347 VSUBS 0.010031f
C388 B.n348 VSUBS 0.010031f
C389 B.n349 VSUBS 0.010031f
C390 B.n350 VSUBS 0.010031f
C391 B.n351 VSUBS 0.010031f
C392 B.n352 VSUBS 0.010031f
C393 B.n353 VSUBS 0.010031f
C394 B.n354 VSUBS 0.010031f
C395 B.n355 VSUBS 0.010031f
C396 B.n356 VSUBS 0.010031f
C397 B.n357 VSUBS 0.010031f
C398 B.n358 VSUBS 0.010031f
C399 B.n359 VSUBS 0.010031f
C400 B.n360 VSUBS 0.010031f
C401 B.n361 VSUBS 0.010031f
C402 B.n362 VSUBS 0.010031f
C403 B.n363 VSUBS 0.010031f
C404 B.n364 VSUBS 0.010031f
C405 B.n365 VSUBS 0.010031f
C406 B.n366 VSUBS 0.010031f
C407 B.n367 VSUBS 0.010031f
C408 B.n368 VSUBS 0.010031f
C409 B.n369 VSUBS 0.010031f
C410 B.n370 VSUBS 0.010031f
C411 B.n371 VSUBS 0.010031f
C412 B.n372 VSUBS 0.010031f
C413 B.n373 VSUBS 0.010031f
C414 B.n374 VSUBS 0.010031f
C415 B.n375 VSUBS 0.010031f
C416 B.n376 VSUBS 0.010031f
C417 B.n377 VSUBS 0.010031f
C418 B.n378 VSUBS 0.010031f
C419 B.n379 VSUBS 0.010031f
C420 B.n380 VSUBS 0.010031f
C421 B.n381 VSUBS 0.010031f
C422 B.n382 VSUBS 0.010031f
C423 B.n383 VSUBS 0.010031f
C424 B.n384 VSUBS 0.010031f
C425 B.n385 VSUBS 0.010031f
C426 B.n386 VSUBS 0.010031f
C427 B.n387 VSUBS 0.010031f
C428 B.n388 VSUBS 0.010031f
C429 B.n389 VSUBS 0.010031f
C430 B.n390 VSUBS 0.010031f
C431 B.n391 VSUBS 0.010031f
C432 B.n392 VSUBS 0.022733f
C433 B.n393 VSUBS 0.023588f
C434 B.n394 VSUBS 0.023588f
C435 B.n395 VSUBS 0.010031f
C436 B.n396 VSUBS 0.010031f
C437 B.n397 VSUBS 0.010031f
C438 B.n398 VSUBS 0.010031f
C439 B.n399 VSUBS 0.010031f
C440 B.n400 VSUBS 0.010031f
C441 B.n401 VSUBS 0.010031f
C442 B.n402 VSUBS 0.010031f
C443 B.n403 VSUBS 0.010031f
C444 B.n404 VSUBS 0.010031f
C445 B.n405 VSUBS 0.010031f
C446 B.n406 VSUBS 0.010031f
C447 B.n407 VSUBS 0.006933f
C448 B.n408 VSUBS 0.023242f
C449 B.n409 VSUBS 0.008114f
C450 B.n410 VSUBS 0.010031f
C451 B.n411 VSUBS 0.010031f
C452 B.n412 VSUBS 0.010031f
C453 B.n413 VSUBS 0.010031f
C454 B.n414 VSUBS 0.010031f
C455 B.n415 VSUBS 0.010031f
C456 B.n416 VSUBS 0.010031f
C457 B.n417 VSUBS 0.010031f
C458 B.n418 VSUBS 0.010031f
C459 B.n419 VSUBS 0.010031f
C460 B.n420 VSUBS 0.010031f
C461 B.n421 VSUBS 0.008114f
C462 B.n422 VSUBS 0.010031f
C463 B.n423 VSUBS 0.010031f
C464 B.n424 VSUBS 0.010031f
C465 B.n425 VSUBS 0.010031f
C466 B.n426 VSUBS 0.010031f
C467 B.n427 VSUBS 0.010031f
C468 B.n428 VSUBS 0.010031f
C469 B.n429 VSUBS 0.010031f
C470 B.n430 VSUBS 0.010031f
C471 B.n431 VSUBS 0.010031f
C472 B.n432 VSUBS 0.010031f
C473 B.n433 VSUBS 0.010031f
C474 B.n434 VSUBS 0.010031f
C475 B.n435 VSUBS 0.010031f
C476 B.n436 VSUBS 0.023588f
C477 B.n437 VSUBS 0.023588f
C478 B.n438 VSUBS 0.022733f
C479 B.n439 VSUBS 0.010031f
C480 B.n440 VSUBS 0.010031f
C481 B.n441 VSUBS 0.010031f
C482 B.n442 VSUBS 0.010031f
C483 B.n443 VSUBS 0.010031f
C484 B.n444 VSUBS 0.010031f
C485 B.n445 VSUBS 0.010031f
C486 B.n446 VSUBS 0.010031f
C487 B.n447 VSUBS 0.010031f
C488 B.n448 VSUBS 0.010031f
C489 B.n449 VSUBS 0.010031f
C490 B.n450 VSUBS 0.010031f
C491 B.n451 VSUBS 0.010031f
C492 B.n452 VSUBS 0.010031f
C493 B.n453 VSUBS 0.010031f
C494 B.n454 VSUBS 0.010031f
C495 B.n455 VSUBS 0.010031f
C496 B.n456 VSUBS 0.010031f
C497 B.n457 VSUBS 0.010031f
C498 B.n458 VSUBS 0.010031f
C499 B.n459 VSUBS 0.010031f
C500 B.n460 VSUBS 0.010031f
C501 B.n461 VSUBS 0.010031f
C502 B.n462 VSUBS 0.010031f
C503 B.n463 VSUBS 0.010031f
C504 B.n464 VSUBS 0.010031f
C505 B.n465 VSUBS 0.010031f
C506 B.n466 VSUBS 0.010031f
C507 B.n467 VSUBS 0.010031f
C508 B.n468 VSUBS 0.010031f
C509 B.n469 VSUBS 0.010031f
C510 B.n470 VSUBS 0.010031f
C511 B.n471 VSUBS 0.010031f
C512 B.n472 VSUBS 0.010031f
C513 B.n473 VSUBS 0.010031f
C514 B.n474 VSUBS 0.010031f
C515 B.n475 VSUBS 0.010031f
C516 B.n476 VSUBS 0.010031f
C517 B.n477 VSUBS 0.010031f
C518 B.n478 VSUBS 0.010031f
C519 B.n479 VSUBS 0.010031f
C520 B.n480 VSUBS 0.010031f
C521 B.n481 VSUBS 0.010031f
C522 B.n482 VSUBS 0.010031f
C523 B.n483 VSUBS 0.010031f
C524 B.n484 VSUBS 0.010031f
C525 B.n485 VSUBS 0.010031f
C526 B.n486 VSUBS 0.010031f
C527 B.n487 VSUBS 0.010031f
C528 B.n488 VSUBS 0.010031f
C529 B.n489 VSUBS 0.010031f
C530 B.n490 VSUBS 0.010031f
C531 B.n491 VSUBS 0.010031f
C532 B.n492 VSUBS 0.010031f
C533 B.n493 VSUBS 0.010031f
C534 B.n494 VSUBS 0.010031f
C535 B.n495 VSUBS 0.010031f
C536 B.n496 VSUBS 0.010031f
C537 B.n497 VSUBS 0.010031f
C538 B.n498 VSUBS 0.010031f
C539 B.n499 VSUBS 0.010031f
C540 B.n500 VSUBS 0.010031f
C541 B.n501 VSUBS 0.010031f
C542 B.n502 VSUBS 0.010031f
C543 B.n503 VSUBS 0.010031f
C544 B.n504 VSUBS 0.010031f
C545 B.n505 VSUBS 0.010031f
C546 B.n506 VSUBS 0.010031f
C547 B.n507 VSUBS 0.01309f
C548 B.n508 VSUBS 0.013945f
C549 B.n509 VSUBS 0.02773f
C550 VDD1.t1 VSUBS 0.092077f
C551 VDD1.t4 VSUBS 0.091959f
C552 VDD1.t3 VSUBS 0.016542f
C553 VDD1.t2 VSUBS 0.016542f
C554 VDD1.n0 VSUBS 0.055761f
C555 VDD1.n1 VSUBS 1.8067f
C556 VDD1.t5 VSUBS 0.016542f
C557 VDD1.t0 VSUBS 0.016542f
C558 VDD1.n2 VSUBS 0.055075f
C559 VDD1.n3 VSUBS 1.47523f
C560 VP.t3 VSUBS 0.418134f
C561 VP.n0 VSUBS 0.471055f
C562 VP.n1 VSUBS 0.059246f
C563 VP.n2 VSUBS 0.07328f
C564 VP.n3 VSUBS 0.059246f
C565 VP.t2 VSUBS 0.418134f
C566 VP.n4 VSUBS 0.110419f
C567 VP.n5 VSUBS 0.059246f
C568 VP.n6 VSUBS 0.110419f
C569 VP.t5 VSUBS 0.418134f
C570 VP.n7 VSUBS 0.471055f
C571 VP.n8 VSUBS 0.059246f
C572 VP.n9 VSUBS 0.07328f
C573 VP.n10 VSUBS 0.673453f
C574 VP.t0 VSUBS 0.418134f
C575 VP.t4 VSUBS 0.929366f
C576 VP.n11 VSUBS 0.471876f
C577 VP.n12 VSUBS 0.468938f
C578 VP.n13 VSUBS 0.110419f
C579 VP.n14 VSUBS 0.110419f
C580 VP.n15 VSUBS 0.059246f
C581 VP.n16 VSUBS 0.059246f
C582 VP.n17 VSUBS 0.059246f
C583 VP.n18 VSUBS 0.099695f
C584 VP.n19 VSUBS 0.110419f
C585 VP.n20 VSUBS 0.092974f
C586 VP.n21 VSUBS 0.095621f
C587 VP.n22 VSUBS 2.59397f
C588 VP.n23 VSUBS 2.64449f
C589 VP.t1 VSUBS 0.418134f
C590 VP.n24 VSUBS 0.471055f
C591 VP.n25 VSUBS 0.092974f
C592 VP.n26 VSUBS 0.095621f
C593 VP.n27 VSUBS 0.059246f
C594 VP.n28 VSUBS 0.059246f
C595 VP.n29 VSUBS 0.099695f
C596 VP.n30 VSUBS 0.07328f
C597 VP.n31 VSUBS 0.110419f
C598 VP.n32 VSUBS 0.059246f
C599 VP.n33 VSUBS 0.059246f
C600 VP.n34 VSUBS 0.059246f
C601 VP.n35 VSUBS 0.305326f
C602 VP.n36 VSUBS 0.110419f
C603 VP.n37 VSUBS 0.110419f
C604 VP.n38 VSUBS 0.059246f
C605 VP.n39 VSUBS 0.059246f
C606 VP.n40 VSUBS 0.059246f
C607 VP.n41 VSUBS 0.099695f
C608 VP.n42 VSUBS 0.110419f
C609 VP.n43 VSUBS 0.092974f
C610 VP.n44 VSUBS 0.095621f
C611 VP.n45 VSUBS 0.131932f
C612 VDD2.t5 VSUBS 0.095745f
C613 VDD2.t2 VSUBS 0.017223f
C614 VDD2.t1 VSUBS 0.017223f
C615 VDD2.n0 VSUBS 0.058057f
C616 VDD2.n1 VSUBS 1.79006f
C617 VDD2.t0 VSUBS 0.094148f
C618 VDD2.n2 VSUBS 1.48894f
C619 VDD2.t3 VSUBS 0.017223f
C620 VDD2.t4 VSUBS 0.017223f
C621 VDD2.n3 VSUBS 0.058053f
C622 VTAIL.t8 VSUBS 0.036498f
C623 VTAIL.t11 VSUBS 0.036498f
C624 VTAIL.n0 VSUBS 0.105453f
C625 VTAIL.n1 VSUBS 0.63048f
C626 VTAIL.t4 VSUBS 0.184332f
C627 VTAIL.n2 VSUBS 0.918428f
C628 VTAIL.t1 VSUBS 0.036498f
C629 VTAIL.t3 VSUBS 0.036498f
C630 VTAIL.n3 VSUBS 0.105453f
C631 VTAIL.n4 VSUBS 2.05191f
C632 VTAIL.t6 VSUBS 0.036498f
C633 VTAIL.t9 VSUBS 0.036498f
C634 VTAIL.n5 VSUBS 0.105453f
C635 VTAIL.n6 VSUBS 2.05192f
C636 VTAIL.t7 VSUBS 0.184332f
C637 VTAIL.n7 VSUBS 0.918428f
C638 VTAIL.t5 VSUBS 0.036498f
C639 VTAIL.t0 VSUBS 0.036498f
C640 VTAIL.n8 VSUBS 0.105453f
C641 VTAIL.n9 VSUBS 0.897767f
C642 VTAIL.t2 VSUBS 0.184332f
C643 VTAIL.n10 VSUBS 1.70633f
C644 VTAIL.t10 VSUBS 0.184332f
C645 VTAIL.n11 VSUBS 1.60736f
C646 VN.t4 VSUBS 0.398938f
C647 VN.n0 VSUBS 0.449429f
C648 VN.n1 VSUBS 0.056526f
C649 VN.n2 VSUBS 0.069916f
C650 VN.n3 VSUBS 0.642534f
C651 VN.t3 VSUBS 0.398938f
C652 VN.t0 VSUBS 0.886701f
C653 VN.n4 VSUBS 0.450212f
C654 VN.n5 VSUBS 0.447409f
C655 VN.n6 VSUBS 0.10535f
C656 VN.n7 VSUBS 0.10535f
C657 VN.n8 VSUBS 0.056526f
C658 VN.n9 VSUBS 0.056526f
C659 VN.n10 VSUBS 0.056526f
C660 VN.n11 VSUBS 0.095119f
C661 VN.n12 VSUBS 0.10535f
C662 VN.n13 VSUBS 0.088706f
C663 VN.n14 VSUBS 0.091231f
C664 VN.n15 VSUBS 0.125875f
C665 VN.t5 VSUBS 0.398938f
C666 VN.n16 VSUBS 0.449429f
C667 VN.n17 VSUBS 0.056526f
C668 VN.n18 VSUBS 0.069916f
C669 VN.n19 VSUBS 0.642534f
C670 VN.t2 VSUBS 0.398938f
C671 VN.t1 VSUBS 0.886701f
C672 VN.n20 VSUBS 0.450212f
C673 VN.n21 VSUBS 0.447409f
C674 VN.n22 VSUBS 0.10535f
C675 VN.n23 VSUBS 0.10535f
C676 VN.n24 VSUBS 0.056526f
C677 VN.n25 VSUBS 0.056526f
C678 VN.n26 VSUBS 0.056526f
C679 VN.n27 VSUBS 0.095119f
C680 VN.n28 VSUBS 0.10535f
C681 VN.n29 VSUBS 0.088706f
C682 VN.n30 VSUBS 0.091231f
C683 VN.n31 VSUBS 2.49951f
.ends

