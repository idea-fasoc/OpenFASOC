* NGSPICE file created from diff_pair_sample_1224.ext - technology: sky130A

.subckt diff_pair_sample_1224 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X1 B.t11 B.t9 B.t10 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=3.75
X2 VTAIL.t14 VP.t1 VDD1.t8 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X3 VDD2.t9 VN.t0 VTAIL.t0 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X4 VDD1.t7 VP.t2 VTAIL.t15 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=3.75
X5 VDD2.t8 VN.t1 VTAIL.t6 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=3.75
X6 VDD2.t7 VN.t2 VTAIL.t4 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=3.75
X7 VTAIL.t2 VN.t3 VDD2.t6 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X8 VTAIL.t18 VP.t3 VDD1.t6 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X9 B.t8 B.t6 B.t7 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=3.75
X10 VDD1.t5 VP.t4 VTAIL.t17 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X11 B.t5 B.t3 B.t4 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=3.75
X12 VDD2.t5 VN.t4 VTAIL.t1 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=3.75
X13 VTAIL.t11 VP.t5 VDD1.t4 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X14 VTAIL.t9 VN.t5 VDD2.t4 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X15 VDD2.t3 VN.t6 VTAIL.t8 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X16 VDD2.t2 VN.t7 VTAIL.t7 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=3.75
X17 B.t2 B.t0 B.t1 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=3.75
X18 VTAIL.t13 VP.t6 VDD1.t3 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X19 VDD1.t2 VP.t7 VTAIL.t10 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=3.75
X20 VTAIL.t3 VN.t8 VDD2.t1 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X21 VDD1.t1 VP.t8 VTAIL.t19 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=3.75
X22 VTAIL.t5 VN.t9 VDD2.t0 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=3.75
X23 VDD1.t0 VP.t9 VTAIL.t16 w_n5866_n3622# sky130_fd_pr__pfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=3.75
R0 VP.n33 VP.n32 161.3
R1 VP.n34 VP.n29 161.3
R2 VP.n36 VP.n35 161.3
R3 VP.n37 VP.n28 161.3
R4 VP.n39 VP.n38 161.3
R5 VP.n40 VP.n27 161.3
R6 VP.n42 VP.n41 161.3
R7 VP.n43 VP.n26 161.3
R8 VP.n45 VP.n44 161.3
R9 VP.n46 VP.n25 161.3
R10 VP.n48 VP.n47 161.3
R11 VP.n49 VP.n24 161.3
R12 VP.n51 VP.n50 161.3
R13 VP.n52 VP.n23 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n22 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n21 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n20 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n19 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n68 VP.n18 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n125 VP.n124 161.3
R26 VP.n123 VP.n1 161.3
R27 VP.n122 VP.n121 161.3
R28 VP.n120 VP.n2 161.3
R29 VP.n119 VP.n118 161.3
R30 VP.n117 VP.n3 161.3
R31 VP.n116 VP.n115 161.3
R32 VP.n114 VP.n4 161.3
R33 VP.n113 VP.n112 161.3
R34 VP.n110 VP.n5 161.3
R35 VP.n109 VP.n108 161.3
R36 VP.n107 VP.n6 161.3
R37 VP.n106 VP.n105 161.3
R38 VP.n104 VP.n7 161.3
R39 VP.n103 VP.n102 161.3
R40 VP.n101 VP.n8 161.3
R41 VP.n100 VP.n99 161.3
R42 VP.n98 VP.n9 161.3
R43 VP.n97 VP.n96 161.3
R44 VP.n95 VP.n10 161.3
R45 VP.n94 VP.n93 161.3
R46 VP.n92 VP.n11 161.3
R47 VP.n91 VP.n90 161.3
R48 VP.n89 VP.n12 161.3
R49 VP.n88 VP.n87 161.3
R50 VP.n85 VP.n13 161.3
R51 VP.n84 VP.n83 161.3
R52 VP.n82 VP.n14 161.3
R53 VP.n81 VP.n80 161.3
R54 VP.n79 VP.n15 161.3
R55 VP.n78 VP.n77 161.3
R56 VP.n76 VP.n16 161.3
R57 VP.n75 VP.n74 161.3
R58 VP.n30 VP.t7 118.285
R59 VP.n99 VP.t0 85.2824
R60 VP.n73 VP.t2 85.2824
R61 VP.n86 VP.t6 85.2824
R62 VP.n111 VP.t1 85.2824
R63 VP.n0 VP.t9 85.2824
R64 VP.n44 VP.t4 85.2824
R65 VP.n17 VP.t8 85.2824
R66 VP.n56 VP.t5 85.2824
R67 VP.n31 VP.t3 85.2824
R68 VP.n73 VP.n72 82.238
R69 VP.n126 VP.n0 82.238
R70 VP.n71 VP.n17 82.238
R71 VP.n31 VP.n30 70.8482
R72 VP.n72 VP.n71 60.4463
R73 VP.n80 VP.n79 52.1486
R74 VP.n118 VP.n2 52.1486
R75 VP.n63 VP.n19 52.1486
R76 VP.n93 VP.n92 44.3785
R77 VP.n105 VP.n6 44.3785
R78 VP.n50 VP.n23 44.3785
R79 VP.n38 VP.n37 44.3785
R80 VP.n93 VP.n10 36.6083
R81 VP.n105 VP.n104 36.6083
R82 VP.n50 VP.n49 36.6083
R83 VP.n38 VP.n27 36.6083
R84 VP.n80 VP.n14 28.8382
R85 VP.n118 VP.n117 28.8382
R86 VP.n63 VP.n62 28.8382
R87 VP.n74 VP.n16 24.4675
R88 VP.n78 VP.n16 24.4675
R89 VP.n79 VP.n78 24.4675
R90 VP.n84 VP.n14 24.4675
R91 VP.n85 VP.n84 24.4675
R92 VP.n87 VP.n12 24.4675
R93 VP.n91 VP.n12 24.4675
R94 VP.n92 VP.n91 24.4675
R95 VP.n97 VP.n10 24.4675
R96 VP.n98 VP.n97 24.4675
R97 VP.n99 VP.n98 24.4675
R98 VP.n99 VP.n8 24.4675
R99 VP.n103 VP.n8 24.4675
R100 VP.n104 VP.n103 24.4675
R101 VP.n109 VP.n6 24.4675
R102 VP.n110 VP.n109 24.4675
R103 VP.n112 VP.n110 24.4675
R104 VP.n116 VP.n4 24.4675
R105 VP.n117 VP.n116 24.4675
R106 VP.n122 VP.n2 24.4675
R107 VP.n123 VP.n122 24.4675
R108 VP.n124 VP.n123 24.4675
R109 VP.n67 VP.n19 24.4675
R110 VP.n68 VP.n67 24.4675
R111 VP.n69 VP.n68 24.4675
R112 VP.n54 VP.n23 24.4675
R113 VP.n55 VP.n54 24.4675
R114 VP.n57 VP.n55 24.4675
R115 VP.n61 VP.n21 24.4675
R116 VP.n62 VP.n61 24.4675
R117 VP.n42 VP.n27 24.4675
R118 VP.n43 VP.n42 24.4675
R119 VP.n44 VP.n43 24.4675
R120 VP.n44 VP.n25 24.4675
R121 VP.n48 VP.n25 24.4675
R122 VP.n49 VP.n48 24.4675
R123 VP.n32 VP.n29 24.4675
R124 VP.n36 VP.n29 24.4675
R125 VP.n37 VP.n36 24.4675
R126 VP.n86 VP.n85 20.5528
R127 VP.n111 VP.n4 20.5528
R128 VP.n56 VP.n21 20.5528
R129 VP.n74 VP.n73 7.82994
R130 VP.n124 VP.n0 7.82994
R131 VP.n69 VP.n17 7.82994
R132 VP.n87 VP.n86 3.91522
R133 VP.n112 VP.n111 3.91522
R134 VP.n57 VP.n56 3.91522
R135 VP.n32 VP.n31 3.91522
R136 VP.n33 VP.n30 3.22185
R137 VP.n71 VP.n70 0.354971
R138 VP.n75 VP.n72 0.354971
R139 VP.n126 VP.n125 0.354971
R140 VP VP.n126 0.26696
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n28 0.189894
R144 VP.n39 VP.n28 0.189894
R145 VP.n40 VP.n39 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n41 VP.n26 0.189894
R148 VP.n45 VP.n26 0.189894
R149 VP.n46 VP.n45 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n47 VP.n24 0.189894
R152 VP.n51 VP.n24 0.189894
R153 VP.n52 VP.n51 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n53 VP.n22 0.189894
R156 VP.n58 VP.n22 0.189894
R157 VP.n59 VP.n58 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n60 VP.n20 0.189894
R160 VP.n64 VP.n20 0.189894
R161 VP.n65 VP.n64 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n66 VP.n18 0.189894
R164 VP.n70 VP.n18 0.189894
R165 VP.n76 VP.n75 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n77 VP.n15 0.189894
R168 VP.n81 VP.n15 0.189894
R169 VP.n82 VP.n81 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n83 VP.n13 0.189894
R172 VP.n88 VP.n13 0.189894
R173 VP.n89 VP.n88 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n90 VP.n11 0.189894
R176 VP.n94 VP.n11 0.189894
R177 VP.n95 VP.n94 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n96 VP.n9 0.189894
R180 VP.n100 VP.n9 0.189894
R181 VP.n101 VP.n100 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n102 VP.n7 0.189894
R184 VP.n106 VP.n7 0.189894
R185 VP.n107 VP.n106 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n108 VP.n5 0.189894
R188 VP.n113 VP.n5 0.189894
R189 VP.n114 VP.n113 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n115 VP.n3 0.189894
R192 VP.n119 VP.n3 0.189894
R193 VP.n120 VP.n119 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n121 VP.n1 0.189894
R196 VP.n125 VP.n1 0.189894
R197 VTAIL.n255 VTAIL.n254 585
R198 VTAIL.n257 VTAIL.n256 585
R199 VTAIL.n250 VTAIL.n249 585
R200 VTAIL.n263 VTAIL.n262 585
R201 VTAIL.n265 VTAIL.n264 585
R202 VTAIL.n246 VTAIL.n245 585
R203 VTAIL.n271 VTAIL.n270 585
R204 VTAIL.n273 VTAIL.n272 585
R205 VTAIL.n242 VTAIL.n241 585
R206 VTAIL.n279 VTAIL.n278 585
R207 VTAIL.n281 VTAIL.n280 585
R208 VTAIL.n238 VTAIL.n237 585
R209 VTAIL.n287 VTAIL.n286 585
R210 VTAIL.n289 VTAIL.n288 585
R211 VTAIL.n234 VTAIL.n233 585
R212 VTAIL.n295 VTAIL.n294 585
R213 VTAIL.n297 VTAIL.n296 585
R214 VTAIL.n27 VTAIL.n26 585
R215 VTAIL.n29 VTAIL.n28 585
R216 VTAIL.n22 VTAIL.n21 585
R217 VTAIL.n35 VTAIL.n34 585
R218 VTAIL.n37 VTAIL.n36 585
R219 VTAIL.n18 VTAIL.n17 585
R220 VTAIL.n43 VTAIL.n42 585
R221 VTAIL.n45 VTAIL.n44 585
R222 VTAIL.n14 VTAIL.n13 585
R223 VTAIL.n51 VTAIL.n50 585
R224 VTAIL.n53 VTAIL.n52 585
R225 VTAIL.n10 VTAIL.n9 585
R226 VTAIL.n59 VTAIL.n58 585
R227 VTAIL.n61 VTAIL.n60 585
R228 VTAIL.n6 VTAIL.n5 585
R229 VTAIL.n67 VTAIL.n66 585
R230 VTAIL.n69 VTAIL.n68 585
R231 VTAIL.n225 VTAIL.n224 585
R232 VTAIL.n223 VTAIL.n222 585
R233 VTAIL.n162 VTAIL.n161 585
R234 VTAIL.n217 VTAIL.n216 585
R235 VTAIL.n215 VTAIL.n214 585
R236 VTAIL.n166 VTAIL.n165 585
R237 VTAIL.n209 VTAIL.n208 585
R238 VTAIL.n207 VTAIL.n206 585
R239 VTAIL.n170 VTAIL.n169 585
R240 VTAIL.n201 VTAIL.n200 585
R241 VTAIL.n199 VTAIL.n198 585
R242 VTAIL.n174 VTAIL.n173 585
R243 VTAIL.n193 VTAIL.n192 585
R244 VTAIL.n191 VTAIL.n190 585
R245 VTAIL.n178 VTAIL.n177 585
R246 VTAIL.n185 VTAIL.n184 585
R247 VTAIL.n183 VTAIL.n182 585
R248 VTAIL.n149 VTAIL.n148 585
R249 VTAIL.n147 VTAIL.n146 585
R250 VTAIL.n86 VTAIL.n85 585
R251 VTAIL.n141 VTAIL.n140 585
R252 VTAIL.n139 VTAIL.n138 585
R253 VTAIL.n90 VTAIL.n89 585
R254 VTAIL.n133 VTAIL.n132 585
R255 VTAIL.n131 VTAIL.n130 585
R256 VTAIL.n94 VTAIL.n93 585
R257 VTAIL.n125 VTAIL.n124 585
R258 VTAIL.n123 VTAIL.n122 585
R259 VTAIL.n98 VTAIL.n97 585
R260 VTAIL.n117 VTAIL.n116 585
R261 VTAIL.n115 VTAIL.n114 585
R262 VTAIL.n102 VTAIL.n101 585
R263 VTAIL.n109 VTAIL.n108 585
R264 VTAIL.n107 VTAIL.n106 585
R265 VTAIL.n296 VTAIL.n230 498.474
R266 VTAIL.n68 VTAIL.n2 498.474
R267 VTAIL.n224 VTAIL.n158 498.474
R268 VTAIL.n148 VTAIL.n82 498.474
R269 VTAIL.n253 VTAIL.t1 327.466
R270 VTAIL.n25 VTAIL.t16 327.466
R271 VTAIL.n181 VTAIL.t19 327.466
R272 VTAIL.n105 VTAIL.t6 327.466
R273 VTAIL.n256 VTAIL.n255 171.744
R274 VTAIL.n256 VTAIL.n249 171.744
R275 VTAIL.n263 VTAIL.n249 171.744
R276 VTAIL.n264 VTAIL.n263 171.744
R277 VTAIL.n264 VTAIL.n245 171.744
R278 VTAIL.n271 VTAIL.n245 171.744
R279 VTAIL.n272 VTAIL.n271 171.744
R280 VTAIL.n272 VTAIL.n241 171.744
R281 VTAIL.n279 VTAIL.n241 171.744
R282 VTAIL.n280 VTAIL.n279 171.744
R283 VTAIL.n280 VTAIL.n237 171.744
R284 VTAIL.n287 VTAIL.n237 171.744
R285 VTAIL.n288 VTAIL.n287 171.744
R286 VTAIL.n288 VTAIL.n233 171.744
R287 VTAIL.n295 VTAIL.n233 171.744
R288 VTAIL.n296 VTAIL.n295 171.744
R289 VTAIL.n28 VTAIL.n27 171.744
R290 VTAIL.n28 VTAIL.n21 171.744
R291 VTAIL.n35 VTAIL.n21 171.744
R292 VTAIL.n36 VTAIL.n35 171.744
R293 VTAIL.n36 VTAIL.n17 171.744
R294 VTAIL.n43 VTAIL.n17 171.744
R295 VTAIL.n44 VTAIL.n43 171.744
R296 VTAIL.n44 VTAIL.n13 171.744
R297 VTAIL.n51 VTAIL.n13 171.744
R298 VTAIL.n52 VTAIL.n51 171.744
R299 VTAIL.n52 VTAIL.n9 171.744
R300 VTAIL.n59 VTAIL.n9 171.744
R301 VTAIL.n60 VTAIL.n59 171.744
R302 VTAIL.n60 VTAIL.n5 171.744
R303 VTAIL.n67 VTAIL.n5 171.744
R304 VTAIL.n68 VTAIL.n67 171.744
R305 VTAIL.n224 VTAIL.n223 171.744
R306 VTAIL.n223 VTAIL.n161 171.744
R307 VTAIL.n216 VTAIL.n161 171.744
R308 VTAIL.n216 VTAIL.n215 171.744
R309 VTAIL.n215 VTAIL.n165 171.744
R310 VTAIL.n208 VTAIL.n165 171.744
R311 VTAIL.n208 VTAIL.n207 171.744
R312 VTAIL.n207 VTAIL.n169 171.744
R313 VTAIL.n200 VTAIL.n169 171.744
R314 VTAIL.n200 VTAIL.n199 171.744
R315 VTAIL.n199 VTAIL.n173 171.744
R316 VTAIL.n192 VTAIL.n173 171.744
R317 VTAIL.n192 VTAIL.n191 171.744
R318 VTAIL.n191 VTAIL.n177 171.744
R319 VTAIL.n184 VTAIL.n177 171.744
R320 VTAIL.n184 VTAIL.n183 171.744
R321 VTAIL.n148 VTAIL.n147 171.744
R322 VTAIL.n147 VTAIL.n85 171.744
R323 VTAIL.n140 VTAIL.n85 171.744
R324 VTAIL.n140 VTAIL.n139 171.744
R325 VTAIL.n139 VTAIL.n89 171.744
R326 VTAIL.n132 VTAIL.n89 171.744
R327 VTAIL.n132 VTAIL.n131 171.744
R328 VTAIL.n131 VTAIL.n93 171.744
R329 VTAIL.n124 VTAIL.n93 171.744
R330 VTAIL.n124 VTAIL.n123 171.744
R331 VTAIL.n123 VTAIL.n97 171.744
R332 VTAIL.n116 VTAIL.n97 171.744
R333 VTAIL.n116 VTAIL.n115 171.744
R334 VTAIL.n115 VTAIL.n101 171.744
R335 VTAIL.n108 VTAIL.n101 171.744
R336 VTAIL.n108 VTAIL.n107 171.744
R337 VTAIL.n255 VTAIL.t1 85.8723
R338 VTAIL.n27 VTAIL.t16 85.8723
R339 VTAIL.n183 VTAIL.t19 85.8723
R340 VTAIL.n107 VTAIL.t6 85.8723
R341 VTAIL.n157 VTAIL.n156 56.6453
R342 VTAIL.n155 VTAIL.n154 56.6453
R343 VTAIL.n81 VTAIL.n80 56.6453
R344 VTAIL.n79 VTAIL.n78 56.6453
R345 VTAIL.n303 VTAIL.n302 56.6452
R346 VTAIL.n1 VTAIL.n0 56.6452
R347 VTAIL.n75 VTAIL.n74 56.6452
R348 VTAIL.n77 VTAIL.n76 56.6452
R349 VTAIL.n301 VTAIL.n300 33.5429
R350 VTAIL.n73 VTAIL.n72 33.5429
R351 VTAIL.n229 VTAIL.n228 33.5429
R352 VTAIL.n153 VTAIL.n152 33.5429
R353 VTAIL.n79 VTAIL.n77 30.841
R354 VTAIL.n301 VTAIL.n229 27.3238
R355 VTAIL.n254 VTAIL.n253 16.3895
R356 VTAIL.n26 VTAIL.n25 16.3895
R357 VTAIL.n182 VTAIL.n181 16.3895
R358 VTAIL.n106 VTAIL.n105 16.3895
R359 VTAIL.n257 VTAIL.n252 12.8005
R360 VTAIL.n298 VTAIL.n297 12.8005
R361 VTAIL.n29 VTAIL.n24 12.8005
R362 VTAIL.n70 VTAIL.n69 12.8005
R363 VTAIL.n226 VTAIL.n225 12.8005
R364 VTAIL.n185 VTAIL.n180 12.8005
R365 VTAIL.n150 VTAIL.n149 12.8005
R366 VTAIL.n109 VTAIL.n104 12.8005
R367 VTAIL.n258 VTAIL.n250 12.0247
R368 VTAIL.n294 VTAIL.n232 12.0247
R369 VTAIL.n30 VTAIL.n22 12.0247
R370 VTAIL.n66 VTAIL.n4 12.0247
R371 VTAIL.n222 VTAIL.n160 12.0247
R372 VTAIL.n186 VTAIL.n178 12.0247
R373 VTAIL.n146 VTAIL.n84 12.0247
R374 VTAIL.n110 VTAIL.n102 12.0247
R375 VTAIL.n262 VTAIL.n261 11.249
R376 VTAIL.n293 VTAIL.n234 11.249
R377 VTAIL.n34 VTAIL.n33 11.249
R378 VTAIL.n65 VTAIL.n6 11.249
R379 VTAIL.n221 VTAIL.n162 11.249
R380 VTAIL.n190 VTAIL.n189 11.249
R381 VTAIL.n145 VTAIL.n86 11.249
R382 VTAIL.n114 VTAIL.n113 11.249
R383 VTAIL.n265 VTAIL.n248 10.4732
R384 VTAIL.n290 VTAIL.n289 10.4732
R385 VTAIL.n37 VTAIL.n20 10.4732
R386 VTAIL.n62 VTAIL.n61 10.4732
R387 VTAIL.n218 VTAIL.n217 10.4732
R388 VTAIL.n193 VTAIL.n176 10.4732
R389 VTAIL.n142 VTAIL.n141 10.4732
R390 VTAIL.n117 VTAIL.n100 10.4732
R391 VTAIL.n266 VTAIL.n246 9.69747
R392 VTAIL.n286 VTAIL.n236 9.69747
R393 VTAIL.n38 VTAIL.n18 9.69747
R394 VTAIL.n58 VTAIL.n8 9.69747
R395 VTAIL.n214 VTAIL.n164 9.69747
R396 VTAIL.n194 VTAIL.n174 9.69747
R397 VTAIL.n138 VTAIL.n88 9.69747
R398 VTAIL.n118 VTAIL.n98 9.69747
R399 VTAIL.n300 VTAIL.n299 9.45567
R400 VTAIL.n72 VTAIL.n71 9.45567
R401 VTAIL.n228 VTAIL.n227 9.45567
R402 VTAIL.n152 VTAIL.n151 9.45567
R403 VTAIL.n275 VTAIL.n274 9.3005
R404 VTAIL.n244 VTAIL.n243 9.3005
R405 VTAIL.n269 VTAIL.n268 9.3005
R406 VTAIL.n267 VTAIL.n266 9.3005
R407 VTAIL.n248 VTAIL.n247 9.3005
R408 VTAIL.n261 VTAIL.n260 9.3005
R409 VTAIL.n259 VTAIL.n258 9.3005
R410 VTAIL.n252 VTAIL.n251 9.3005
R411 VTAIL.n277 VTAIL.n276 9.3005
R412 VTAIL.n240 VTAIL.n239 9.3005
R413 VTAIL.n283 VTAIL.n282 9.3005
R414 VTAIL.n285 VTAIL.n284 9.3005
R415 VTAIL.n236 VTAIL.n235 9.3005
R416 VTAIL.n291 VTAIL.n290 9.3005
R417 VTAIL.n293 VTAIL.n292 9.3005
R418 VTAIL.n232 VTAIL.n231 9.3005
R419 VTAIL.n299 VTAIL.n298 9.3005
R420 VTAIL.n47 VTAIL.n46 9.3005
R421 VTAIL.n16 VTAIL.n15 9.3005
R422 VTAIL.n41 VTAIL.n40 9.3005
R423 VTAIL.n39 VTAIL.n38 9.3005
R424 VTAIL.n20 VTAIL.n19 9.3005
R425 VTAIL.n33 VTAIL.n32 9.3005
R426 VTAIL.n31 VTAIL.n30 9.3005
R427 VTAIL.n24 VTAIL.n23 9.3005
R428 VTAIL.n49 VTAIL.n48 9.3005
R429 VTAIL.n12 VTAIL.n11 9.3005
R430 VTAIL.n55 VTAIL.n54 9.3005
R431 VTAIL.n57 VTAIL.n56 9.3005
R432 VTAIL.n8 VTAIL.n7 9.3005
R433 VTAIL.n63 VTAIL.n62 9.3005
R434 VTAIL.n65 VTAIL.n64 9.3005
R435 VTAIL.n4 VTAIL.n3 9.3005
R436 VTAIL.n71 VTAIL.n70 9.3005
R437 VTAIL.n168 VTAIL.n167 9.3005
R438 VTAIL.n211 VTAIL.n210 9.3005
R439 VTAIL.n213 VTAIL.n212 9.3005
R440 VTAIL.n164 VTAIL.n163 9.3005
R441 VTAIL.n219 VTAIL.n218 9.3005
R442 VTAIL.n221 VTAIL.n220 9.3005
R443 VTAIL.n160 VTAIL.n159 9.3005
R444 VTAIL.n227 VTAIL.n226 9.3005
R445 VTAIL.n205 VTAIL.n204 9.3005
R446 VTAIL.n203 VTAIL.n202 9.3005
R447 VTAIL.n172 VTAIL.n171 9.3005
R448 VTAIL.n197 VTAIL.n196 9.3005
R449 VTAIL.n195 VTAIL.n194 9.3005
R450 VTAIL.n176 VTAIL.n175 9.3005
R451 VTAIL.n189 VTAIL.n188 9.3005
R452 VTAIL.n187 VTAIL.n186 9.3005
R453 VTAIL.n180 VTAIL.n179 9.3005
R454 VTAIL.n92 VTAIL.n91 9.3005
R455 VTAIL.n135 VTAIL.n134 9.3005
R456 VTAIL.n137 VTAIL.n136 9.3005
R457 VTAIL.n88 VTAIL.n87 9.3005
R458 VTAIL.n143 VTAIL.n142 9.3005
R459 VTAIL.n145 VTAIL.n144 9.3005
R460 VTAIL.n84 VTAIL.n83 9.3005
R461 VTAIL.n151 VTAIL.n150 9.3005
R462 VTAIL.n129 VTAIL.n128 9.3005
R463 VTAIL.n127 VTAIL.n126 9.3005
R464 VTAIL.n96 VTAIL.n95 9.3005
R465 VTAIL.n121 VTAIL.n120 9.3005
R466 VTAIL.n119 VTAIL.n118 9.3005
R467 VTAIL.n100 VTAIL.n99 9.3005
R468 VTAIL.n113 VTAIL.n112 9.3005
R469 VTAIL.n111 VTAIL.n110 9.3005
R470 VTAIL.n104 VTAIL.n103 9.3005
R471 VTAIL.n270 VTAIL.n269 8.92171
R472 VTAIL.n285 VTAIL.n238 8.92171
R473 VTAIL.n42 VTAIL.n41 8.92171
R474 VTAIL.n57 VTAIL.n10 8.92171
R475 VTAIL.n213 VTAIL.n166 8.92171
R476 VTAIL.n198 VTAIL.n197 8.92171
R477 VTAIL.n137 VTAIL.n90 8.92171
R478 VTAIL.n122 VTAIL.n121 8.92171
R479 VTAIL.n273 VTAIL.n244 8.14595
R480 VTAIL.n282 VTAIL.n281 8.14595
R481 VTAIL.n45 VTAIL.n16 8.14595
R482 VTAIL.n54 VTAIL.n53 8.14595
R483 VTAIL.n210 VTAIL.n209 8.14595
R484 VTAIL.n201 VTAIL.n172 8.14595
R485 VTAIL.n134 VTAIL.n133 8.14595
R486 VTAIL.n125 VTAIL.n96 8.14595
R487 VTAIL.n300 VTAIL.n230 7.75445
R488 VTAIL.n72 VTAIL.n2 7.75445
R489 VTAIL.n228 VTAIL.n158 7.75445
R490 VTAIL.n152 VTAIL.n82 7.75445
R491 VTAIL.n274 VTAIL.n242 7.3702
R492 VTAIL.n278 VTAIL.n240 7.3702
R493 VTAIL.n46 VTAIL.n14 7.3702
R494 VTAIL.n50 VTAIL.n12 7.3702
R495 VTAIL.n206 VTAIL.n168 7.3702
R496 VTAIL.n202 VTAIL.n170 7.3702
R497 VTAIL.n130 VTAIL.n92 7.3702
R498 VTAIL.n126 VTAIL.n94 7.3702
R499 VTAIL.n277 VTAIL.n242 6.59444
R500 VTAIL.n278 VTAIL.n277 6.59444
R501 VTAIL.n49 VTAIL.n14 6.59444
R502 VTAIL.n50 VTAIL.n49 6.59444
R503 VTAIL.n206 VTAIL.n205 6.59444
R504 VTAIL.n205 VTAIL.n170 6.59444
R505 VTAIL.n130 VTAIL.n129 6.59444
R506 VTAIL.n129 VTAIL.n94 6.59444
R507 VTAIL.n298 VTAIL.n230 6.08283
R508 VTAIL.n70 VTAIL.n2 6.08283
R509 VTAIL.n226 VTAIL.n158 6.08283
R510 VTAIL.n150 VTAIL.n82 6.08283
R511 VTAIL.n274 VTAIL.n273 5.81868
R512 VTAIL.n281 VTAIL.n240 5.81868
R513 VTAIL.n46 VTAIL.n45 5.81868
R514 VTAIL.n53 VTAIL.n12 5.81868
R515 VTAIL.n209 VTAIL.n168 5.81868
R516 VTAIL.n202 VTAIL.n201 5.81868
R517 VTAIL.n133 VTAIL.n92 5.81868
R518 VTAIL.n126 VTAIL.n125 5.81868
R519 VTAIL.n270 VTAIL.n244 5.04292
R520 VTAIL.n282 VTAIL.n238 5.04292
R521 VTAIL.n42 VTAIL.n16 5.04292
R522 VTAIL.n54 VTAIL.n10 5.04292
R523 VTAIL.n210 VTAIL.n166 5.04292
R524 VTAIL.n198 VTAIL.n172 5.04292
R525 VTAIL.n134 VTAIL.n90 5.04292
R526 VTAIL.n122 VTAIL.n96 5.04292
R527 VTAIL.n269 VTAIL.n246 4.26717
R528 VTAIL.n286 VTAIL.n285 4.26717
R529 VTAIL.n41 VTAIL.n18 4.26717
R530 VTAIL.n58 VTAIL.n57 4.26717
R531 VTAIL.n214 VTAIL.n213 4.26717
R532 VTAIL.n197 VTAIL.n174 4.26717
R533 VTAIL.n138 VTAIL.n137 4.26717
R534 VTAIL.n121 VTAIL.n98 4.26717
R535 VTAIL.n253 VTAIL.n251 3.70982
R536 VTAIL.n25 VTAIL.n23 3.70982
R537 VTAIL.n181 VTAIL.n179 3.70982
R538 VTAIL.n105 VTAIL.n103 3.70982
R539 VTAIL.n81 VTAIL.n79 3.51774
R540 VTAIL.n153 VTAIL.n81 3.51774
R541 VTAIL.n157 VTAIL.n155 3.51774
R542 VTAIL.n229 VTAIL.n157 3.51774
R543 VTAIL.n77 VTAIL.n75 3.51774
R544 VTAIL.n75 VTAIL.n73 3.51774
R545 VTAIL.n303 VTAIL.n301 3.51774
R546 VTAIL.n266 VTAIL.n265 3.49141
R547 VTAIL.n289 VTAIL.n236 3.49141
R548 VTAIL.n38 VTAIL.n37 3.49141
R549 VTAIL.n61 VTAIL.n8 3.49141
R550 VTAIL.n217 VTAIL.n164 3.49141
R551 VTAIL.n194 VTAIL.n193 3.49141
R552 VTAIL.n141 VTAIL.n88 3.49141
R553 VTAIL.n118 VTAIL.n117 3.49141
R554 VTAIL.n262 VTAIL.n248 2.71565
R555 VTAIL.n290 VTAIL.n234 2.71565
R556 VTAIL.n34 VTAIL.n20 2.71565
R557 VTAIL.n62 VTAIL.n6 2.71565
R558 VTAIL.n218 VTAIL.n162 2.71565
R559 VTAIL.n190 VTAIL.n176 2.71565
R560 VTAIL.n142 VTAIL.n86 2.71565
R561 VTAIL.n114 VTAIL.n100 2.71565
R562 VTAIL VTAIL.n1 2.69662
R563 VTAIL.n302 VTAIL.t8 2.45001
R564 VTAIL.n302 VTAIL.t3 2.45001
R565 VTAIL.n0 VTAIL.t4 2.45001
R566 VTAIL.n0 VTAIL.t5 2.45001
R567 VTAIL.n74 VTAIL.t12 2.45001
R568 VTAIL.n74 VTAIL.t14 2.45001
R569 VTAIL.n76 VTAIL.t15 2.45001
R570 VTAIL.n76 VTAIL.t13 2.45001
R571 VTAIL.n156 VTAIL.t17 2.45001
R572 VTAIL.n156 VTAIL.t11 2.45001
R573 VTAIL.n154 VTAIL.t10 2.45001
R574 VTAIL.n154 VTAIL.t18 2.45001
R575 VTAIL.n80 VTAIL.t0 2.45001
R576 VTAIL.n80 VTAIL.t9 2.45001
R577 VTAIL.n78 VTAIL.t7 2.45001
R578 VTAIL.n78 VTAIL.t2 2.45001
R579 VTAIL.n155 VTAIL.n153 2.22895
R580 VTAIL.n73 VTAIL.n1 2.22895
R581 VTAIL.n261 VTAIL.n250 1.93989
R582 VTAIL.n294 VTAIL.n293 1.93989
R583 VTAIL.n33 VTAIL.n22 1.93989
R584 VTAIL.n66 VTAIL.n65 1.93989
R585 VTAIL.n222 VTAIL.n221 1.93989
R586 VTAIL.n189 VTAIL.n178 1.93989
R587 VTAIL.n146 VTAIL.n145 1.93989
R588 VTAIL.n113 VTAIL.n102 1.93989
R589 VTAIL.n258 VTAIL.n257 1.16414
R590 VTAIL.n297 VTAIL.n232 1.16414
R591 VTAIL.n30 VTAIL.n29 1.16414
R592 VTAIL.n69 VTAIL.n4 1.16414
R593 VTAIL.n225 VTAIL.n160 1.16414
R594 VTAIL.n186 VTAIL.n185 1.16414
R595 VTAIL.n149 VTAIL.n84 1.16414
R596 VTAIL.n110 VTAIL.n109 1.16414
R597 VTAIL VTAIL.n303 0.821621
R598 VTAIL.n254 VTAIL.n252 0.388379
R599 VTAIL.n26 VTAIL.n24 0.388379
R600 VTAIL.n182 VTAIL.n180 0.388379
R601 VTAIL.n106 VTAIL.n104 0.388379
R602 VTAIL.n259 VTAIL.n251 0.155672
R603 VTAIL.n260 VTAIL.n259 0.155672
R604 VTAIL.n260 VTAIL.n247 0.155672
R605 VTAIL.n267 VTAIL.n247 0.155672
R606 VTAIL.n268 VTAIL.n267 0.155672
R607 VTAIL.n268 VTAIL.n243 0.155672
R608 VTAIL.n275 VTAIL.n243 0.155672
R609 VTAIL.n276 VTAIL.n275 0.155672
R610 VTAIL.n276 VTAIL.n239 0.155672
R611 VTAIL.n283 VTAIL.n239 0.155672
R612 VTAIL.n284 VTAIL.n283 0.155672
R613 VTAIL.n284 VTAIL.n235 0.155672
R614 VTAIL.n291 VTAIL.n235 0.155672
R615 VTAIL.n292 VTAIL.n291 0.155672
R616 VTAIL.n292 VTAIL.n231 0.155672
R617 VTAIL.n299 VTAIL.n231 0.155672
R618 VTAIL.n31 VTAIL.n23 0.155672
R619 VTAIL.n32 VTAIL.n31 0.155672
R620 VTAIL.n32 VTAIL.n19 0.155672
R621 VTAIL.n39 VTAIL.n19 0.155672
R622 VTAIL.n40 VTAIL.n39 0.155672
R623 VTAIL.n40 VTAIL.n15 0.155672
R624 VTAIL.n47 VTAIL.n15 0.155672
R625 VTAIL.n48 VTAIL.n47 0.155672
R626 VTAIL.n48 VTAIL.n11 0.155672
R627 VTAIL.n55 VTAIL.n11 0.155672
R628 VTAIL.n56 VTAIL.n55 0.155672
R629 VTAIL.n56 VTAIL.n7 0.155672
R630 VTAIL.n63 VTAIL.n7 0.155672
R631 VTAIL.n64 VTAIL.n63 0.155672
R632 VTAIL.n64 VTAIL.n3 0.155672
R633 VTAIL.n71 VTAIL.n3 0.155672
R634 VTAIL.n227 VTAIL.n159 0.155672
R635 VTAIL.n220 VTAIL.n159 0.155672
R636 VTAIL.n220 VTAIL.n219 0.155672
R637 VTAIL.n219 VTAIL.n163 0.155672
R638 VTAIL.n212 VTAIL.n163 0.155672
R639 VTAIL.n212 VTAIL.n211 0.155672
R640 VTAIL.n211 VTAIL.n167 0.155672
R641 VTAIL.n204 VTAIL.n167 0.155672
R642 VTAIL.n204 VTAIL.n203 0.155672
R643 VTAIL.n203 VTAIL.n171 0.155672
R644 VTAIL.n196 VTAIL.n171 0.155672
R645 VTAIL.n196 VTAIL.n195 0.155672
R646 VTAIL.n195 VTAIL.n175 0.155672
R647 VTAIL.n188 VTAIL.n175 0.155672
R648 VTAIL.n188 VTAIL.n187 0.155672
R649 VTAIL.n187 VTAIL.n179 0.155672
R650 VTAIL.n151 VTAIL.n83 0.155672
R651 VTAIL.n144 VTAIL.n83 0.155672
R652 VTAIL.n144 VTAIL.n143 0.155672
R653 VTAIL.n143 VTAIL.n87 0.155672
R654 VTAIL.n136 VTAIL.n87 0.155672
R655 VTAIL.n136 VTAIL.n135 0.155672
R656 VTAIL.n135 VTAIL.n91 0.155672
R657 VTAIL.n128 VTAIL.n91 0.155672
R658 VTAIL.n128 VTAIL.n127 0.155672
R659 VTAIL.n127 VTAIL.n95 0.155672
R660 VTAIL.n120 VTAIL.n95 0.155672
R661 VTAIL.n120 VTAIL.n119 0.155672
R662 VTAIL.n119 VTAIL.n99 0.155672
R663 VTAIL.n112 VTAIL.n99 0.155672
R664 VTAIL.n112 VTAIL.n111 0.155672
R665 VTAIL.n111 VTAIL.n103 0.155672
R666 VDD1.n67 VDD1.n66 585
R667 VDD1.n65 VDD1.n64 585
R668 VDD1.n4 VDD1.n3 585
R669 VDD1.n59 VDD1.n58 585
R670 VDD1.n57 VDD1.n56 585
R671 VDD1.n8 VDD1.n7 585
R672 VDD1.n51 VDD1.n50 585
R673 VDD1.n49 VDD1.n48 585
R674 VDD1.n12 VDD1.n11 585
R675 VDD1.n43 VDD1.n42 585
R676 VDD1.n41 VDD1.n40 585
R677 VDD1.n16 VDD1.n15 585
R678 VDD1.n35 VDD1.n34 585
R679 VDD1.n33 VDD1.n32 585
R680 VDD1.n20 VDD1.n19 585
R681 VDD1.n27 VDD1.n26 585
R682 VDD1.n25 VDD1.n24 585
R683 VDD1.n98 VDD1.n97 585
R684 VDD1.n100 VDD1.n99 585
R685 VDD1.n93 VDD1.n92 585
R686 VDD1.n106 VDD1.n105 585
R687 VDD1.n108 VDD1.n107 585
R688 VDD1.n89 VDD1.n88 585
R689 VDD1.n114 VDD1.n113 585
R690 VDD1.n116 VDD1.n115 585
R691 VDD1.n85 VDD1.n84 585
R692 VDD1.n122 VDD1.n121 585
R693 VDD1.n124 VDD1.n123 585
R694 VDD1.n81 VDD1.n80 585
R695 VDD1.n130 VDD1.n129 585
R696 VDD1.n132 VDD1.n131 585
R697 VDD1.n77 VDD1.n76 585
R698 VDD1.n138 VDD1.n137 585
R699 VDD1.n140 VDD1.n139 585
R700 VDD1.n66 VDD1.n0 498.474
R701 VDD1.n139 VDD1.n73 498.474
R702 VDD1.n23 VDD1.t2 327.466
R703 VDD1.n96 VDD1.t7 327.466
R704 VDD1.n66 VDD1.n65 171.744
R705 VDD1.n65 VDD1.n3 171.744
R706 VDD1.n58 VDD1.n3 171.744
R707 VDD1.n58 VDD1.n57 171.744
R708 VDD1.n57 VDD1.n7 171.744
R709 VDD1.n50 VDD1.n7 171.744
R710 VDD1.n50 VDD1.n49 171.744
R711 VDD1.n49 VDD1.n11 171.744
R712 VDD1.n42 VDD1.n11 171.744
R713 VDD1.n42 VDD1.n41 171.744
R714 VDD1.n41 VDD1.n15 171.744
R715 VDD1.n34 VDD1.n15 171.744
R716 VDD1.n34 VDD1.n33 171.744
R717 VDD1.n33 VDD1.n19 171.744
R718 VDD1.n26 VDD1.n19 171.744
R719 VDD1.n26 VDD1.n25 171.744
R720 VDD1.n99 VDD1.n98 171.744
R721 VDD1.n99 VDD1.n92 171.744
R722 VDD1.n106 VDD1.n92 171.744
R723 VDD1.n107 VDD1.n106 171.744
R724 VDD1.n107 VDD1.n88 171.744
R725 VDD1.n114 VDD1.n88 171.744
R726 VDD1.n115 VDD1.n114 171.744
R727 VDD1.n115 VDD1.n84 171.744
R728 VDD1.n122 VDD1.n84 171.744
R729 VDD1.n123 VDD1.n122 171.744
R730 VDD1.n123 VDD1.n80 171.744
R731 VDD1.n130 VDD1.n80 171.744
R732 VDD1.n131 VDD1.n130 171.744
R733 VDD1.n131 VDD1.n76 171.744
R734 VDD1.n138 VDD1.n76 171.744
R735 VDD1.n139 VDD1.n138 171.744
R736 VDD1.n25 VDD1.t2 85.8723
R737 VDD1.n98 VDD1.t7 85.8723
R738 VDD1.n147 VDD1.n146 75.9066
R739 VDD1.n72 VDD1.n71 73.3241
R740 VDD1.n149 VDD1.n148 73.324
R741 VDD1.n145 VDD1.n144 73.324
R742 VDD1.n149 VDD1.n147 54.2035
R743 VDD1.n72 VDD1.n70 53.739
R744 VDD1.n145 VDD1.n143 53.739
R745 VDD1.n24 VDD1.n23 16.3895
R746 VDD1.n97 VDD1.n96 16.3895
R747 VDD1.n68 VDD1.n67 12.8005
R748 VDD1.n27 VDD1.n22 12.8005
R749 VDD1.n100 VDD1.n95 12.8005
R750 VDD1.n141 VDD1.n140 12.8005
R751 VDD1.n64 VDD1.n2 12.0247
R752 VDD1.n28 VDD1.n20 12.0247
R753 VDD1.n101 VDD1.n93 12.0247
R754 VDD1.n137 VDD1.n75 12.0247
R755 VDD1.n63 VDD1.n4 11.249
R756 VDD1.n32 VDD1.n31 11.249
R757 VDD1.n105 VDD1.n104 11.249
R758 VDD1.n136 VDD1.n77 11.249
R759 VDD1.n60 VDD1.n59 10.4732
R760 VDD1.n35 VDD1.n18 10.4732
R761 VDD1.n108 VDD1.n91 10.4732
R762 VDD1.n133 VDD1.n132 10.4732
R763 VDD1.n56 VDD1.n6 9.69747
R764 VDD1.n36 VDD1.n16 9.69747
R765 VDD1.n109 VDD1.n89 9.69747
R766 VDD1.n129 VDD1.n79 9.69747
R767 VDD1.n70 VDD1.n69 9.45567
R768 VDD1.n143 VDD1.n142 9.45567
R769 VDD1.n10 VDD1.n9 9.3005
R770 VDD1.n53 VDD1.n52 9.3005
R771 VDD1.n55 VDD1.n54 9.3005
R772 VDD1.n6 VDD1.n5 9.3005
R773 VDD1.n61 VDD1.n60 9.3005
R774 VDD1.n63 VDD1.n62 9.3005
R775 VDD1.n2 VDD1.n1 9.3005
R776 VDD1.n69 VDD1.n68 9.3005
R777 VDD1.n47 VDD1.n46 9.3005
R778 VDD1.n45 VDD1.n44 9.3005
R779 VDD1.n14 VDD1.n13 9.3005
R780 VDD1.n39 VDD1.n38 9.3005
R781 VDD1.n37 VDD1.n36 9.3005
R782 VDD1.n18 VDD1.n17 9.3005
R783 VDD1.n31 VDD1.n30 9.3005
R784 VDD1.n29 VDD1.n28 9.3005
R785 VDD1.n22 VDD1.n21 9.3005
R786 VDD1.n118 VDD1.n117 9.3005
R787 VDD1.n87 VDD1.n86 9.3005
R788 VDD1.n112 VDD1.n111 9.3005
R789 VDD1.n110 VDD1.n109 9.3005
R790 VDD1.n91 VDD1.n90 9.3005
R791 VDD1.n104 VDD1.n103 9.3005
R792 VDD1.n102 VDD1.n101 9.3005
R793 VDD1.n95 VDD1.n94 9.3005
R794 VDD1.n120 VDD1.n119 9.3005
R795 VDD1.n83 VDD1.n82 9.3005
R796 VDD1.n126 VDD1.n125 9.3005
R797 VDD1.n128 VDD1.n127 9.3005
R798 VDD1.n79 VDD1.n78 9.3005
R799 VDD1.n134 VDD1.n133 9.3005
R800 VDD1.n136 VDD1.n135 9.3005
R801 VDD1.n75 VDD1.n74 9.3005
R802 VDD1.n142 VDD1.n141 9.3005
R803 VDD1.n55 VDD1.n8 8.92171
R804 VDD1.n40 VDD1.n39 8.92171
R805 VDD1.n113 VDD1.n112 8.92171
R806 VDD1.n128 VDD1.n81 8.92171
R807 VDD1.n52 VDD1.n51 8.14595
R808 VDD1.n43 VDD1.n14 8.14595
R809 VDD1.n116 VDD1.n87 8.14595
R810 VDD1.n125 VDD1.n124 8.14595
R811 VDD1.n70 VDD1.n0 7.75445
R812 VDD1.n143 VDD1.n73 7.75445
R813 VDD1.n48 VDD1.n10 7.3702
R814 VDD1.n44 VDD1.n12 7.3702
R815 VDD1.n117 VDD1.n85 7.3702
R816 VDD1.n121 VDD1.n83 7.3702
R817 VDD1.n48 VDD1.n47 6.59444
R818 VDD1.n47 VDD1.n12 6.59444
R819 VDD1.n120 VDD1.n85 6.59444
R820 VDD1.n121 VDD1.n120 6.59444
R821 VDD1.n68 VDD1.n0 6.08283
R822 VDD1.n141 VDD1.n73 6.08283
R823 VDD1.n51 VDD1.n10 5.81868
R824 VDD1.n44 VDD1.n43 5.81868
R825 VDD1.n117 VDD1.n116 5.81868
R826 VDD1.n124 VDD1.n83 5.81868
R827 VDD1.n52 VDD1.n8 5.04292
R828 VDD1.n40 VDD1.n14 5.04292
R829 VDD1.n113 VDD1.n87 5.04292
R830 VDD1.n125 VDD1.n81 5.04292
R831 VDD1.n56 VDD1.n55 4.26717
R832 VDD1.n39 VDD1.n16 4.26717
R833 VDD1.n112 VDD1.n89 4.26717
R834 VDD1.n129 VDD1.n128 4.26717
R835 VDD1.n23 VDD1.n21 3.70982
R836 VDD1.n96 VDD1.n94 3.70982
R837 VDD1.n59 VDD1.n6 3.49141
R838 VDD1.n36 VDD1.n35 3.49141
R839 VDD1.n109 VDD1.n108 3.49141
R840 VDD1.n132 VDD1.n79 3.49141
R841 VDD1.n60 VDD1.n4 2.71565
R842 VDD1.n32 VDD1.n18 2.71565
R843 VDD1.n105 VDD1.n91 2.71565
R844 VDD1.n133 VDD1.n77 2.71565
R845 VDD1 VDD1.n149 2.58024
R846 VDD1.n148 VDD1.t4 2.45001
R847 VDD1.n148 VDD1.t1 2.45001
R848 VDD1.n71 VDD1.t6 2.45001
R849 VDD1.n71 VDD1.t5 2.45001
R850 VDD1.n146 VDD1.t8 2.45001
R851 VDD1.n146 VDD1.t0 2.45001
R852 VDD1.n144 VDD1.t3 2.45001
R853 VDD1.n144 VDD1.t9 2.45001
R854 VDD1.n64 VDD1.n63 1.93989
R855 VDD1.n31 VDD1.n20 1.93989
R856 VDD1.n104 VDD1.n93 1.93989
R857 VDD1.n137 VDD1.n136 1.93989
R858 VDD1.n67 VDD1.n2 1.16414
R859 VDD1.n28 VDD1.n27 1.16414
R860 VDD1.n101 VDD1.n100 1.16414
R861 VDD1.n140 VDD1.n75 1.16414
R862 VDD1 VDD1.n72 0.938
R863 VDD1.n147 VDD1.n145 0.824464
R864 VDD1.n24 VDD1.n22 0.388379
R865 VDD1.n97 VDD1.n95 0.388379
R866 VDD1.n69 VDD1.n1 0.155672
R867 VDD1.n62 VDD1.n1 0.155672
R868 VDD1.n62 VDD1.n61 0.155672
R869 VDD1.n61 VDD1.n5 0.155672
R870 VDD1.n54 VDD1.n5 0.155672
R871 VDD1.n54 VDD1.n53 0.155672
R872 VDD1.n53 VDD1.n9 0.155672
R873 VDD1.n46 VDD1.n9 0.155672
R874 VDD1.n46 VDD1.n45 0.155672
R875 VDD1.n45 VDD1.n13 0.155672
R876 VDD1.n38 VDD1.n13 0.155672
R877 VDD1.n38 VDD1.n37 0.155672
R878 VDD1.n37 VDD1.n17 0.155672
R879 VDD1.n30 VDD1.n17 0.155672
R880 VDD1.n30 VDD1.n29 0.155672
R881 VDD1.n29 VDD1.n21 0.155672
R882 VDD1.n102 VDD1.n94 0.155672
R883 VDD1.n103 VDD1.n102 0.155672
R884 VDD1.n103 VDD1.n90 0.155672
R885 VDD1.n110 VDD1.n90 0.155672
R886 VDD1.n111 VDD1.n110 0.155672
R887 VDD1.n111 VDD1.n86 0.155672
R888 VDD1.n118 VDD1.n86 0.155672
R889 VDD1.n119 VDD1.n118 0.155672
R890 VDD1.n119 VDD1.n82 0.155672
R891 VDD1.n126 VDD1.n82 0.155672
R892 VDD1.n127 VDD1.n126 0.155672
R893 VDD1.n127 VDD1.n78 0.155672
R894 VDD1.n134 VDD1.n78 0.155672
R895 VDD1.n135 VDD1.n134 0.155672
R896 VDD1.n135 VDD1.n74 0.155672
R897 VDD1.n142 VDD1.n74 0.155672
R898 B.n784 B.n783 585
R899 B.n785 B.n96 585
R900 B.n787 B.n786 585
R901 B.n788 B.n95 585
R902 B.n790 B.n789 585
R903 B.n791 B.n94 585
R904 B.n793 B.n792 585
R905 B.n794 B.n93 585
R906 B.n796 B.n795 585
R907 B.n797 B.n92 585
R908 B.n799 B.n798 585
R909 B.n800 B.n91 585
R910 B.n802 B.n801 585
R911 B.n803 B.n90 585
R912 B.n805 B.n804 585
R913 B.n806 B.n89 585
R914 B.n808 B.n807 585
R915 B.n809 B.n88 585
R916 B.n811 B.n810 585
R917 B.n812 B.n87 585
R918 B.n814 B.n813 585
R919 B.n815 B.n86 585
R920 B.n817 B.n816 585
R921 B.n818 B.n85 585
R922 B.n820 B.n819 585
R923 B.n821 B.n84 585
R924 B.n823 B.n822 585
R925 B.n824 B.n83 585
R926 B.n826 B.n825 585
R927 B.n827 B.n82 585
R928 B.n829 B.n828 585
R929 B.n830 B.n81 585
R930 B.n832 B.n831 585
R931 B.n833 B.n80 585
R932 B.n835 B.n834 585
R933 B.n836 B.n79 585
R934 B.n838 B.n837 585
R935 B.n839 B.n78 585
R936 B.n841 B.n840 585
R937 B.n842 B.n77 585
R938 B.n844 B.n843 585
R939 B.n845 B.n76 585
R940 B.n847 B.n846 585
R941 B.n848 B.n75 585
R942 B.n850 B.n849 585
R943 B.n852 B.n72 585
R944 B.n854 B.n853 585
R945 B.n855 B.n71 585
R946 B.n857 B.n856 585
R947 B.n858 B.n70 585
R948 B.n860 B.n859 585
R949 B.n861 B.n69 585
R950 B.n863 B.n862 585
R951 B.n864 B.n65 585
R952 B.n866 B.n865 585
R953 B.n867 B.n64 585
R954 B.n869 B.n868 585
R955 B.n870 B.n63 585
R956 B.n872 B.n871 585
R957 B.n873 B.n62 585
R958 B.n875 B.n874 585
R959 B.n876 B.n61 585
R960 B.n878 B.n877 585
R961 B.n879 B.n60 585
R962 B.n881 B.n880 585
R963 B.n882 B.n59 585
R964 B.n884 B.n883 585
R965 B.n885 B.n58 585
R966 B.n887 B.n886 585
R967 B.n888 B.n57 585
R968 B.n890 B.n889 585
R969 B.n891 B.n56 585
R970 B.n893 B.n892 585
R971 B.n894 B.n55 585
R972 B.n896 B.n895 585
R973 B.n897 B.n54 585
R974 B.n899 B.n898 585
R975 B.n900 B.n53 585
R976 B.n902 B.n901 585
R977 B.n903 B.n52 585
R978 B.n905 B.n904 585
R979 B.n906 B.n51 585
R980 B.n908 B.n907 585
R981 B.n909 B.n50 585
R982 B.n911 B.n910 585
R983 B.n912 B.n49 585
R984 B.n914 B.n913 585
R985 B.n915 B.n48 585
R986 B.n917 B.n916 585
R987 B.n918 B.n47 585
R988 B.n920 B.n919 585
R989 B.n921 B.n46 585
R990 B.n923 B.n922 585
R991 B.n924 B.n45 585
R992 B.n926 B.n925 585
R993 B.n927 B.n44 585
R994 B.n929 B.n928 585
R995 B.n930 B.n43 585
R996 B.n932 B.n931 585
R997 B.n933 B.n42 585
R998 B.n782 B.n97 585
R999 B.n781 B.n780 585
R1000 B.n779 B.n98 585
R1001 B.n778 B.n777 585
R1002 B.n776 B.n99 585
R1003 B.n775 B.n774 585
R1004 B.n773 B.n100 585
R1005 B.n772 B.n771 585
R1006 B.n770 B.n101 585
R1007 B.n769 B.n768 585
R1008 B.n767 B.n102 585
R1009 B.n766 B.n765 585
R1010 B.n764 B.n103 585
R1011 B.n763 B.n762 585
R1012 B.n761 B.n104 585
R1013 B.n760 B.n759 585
R1014 B.n758 B.n105 585
R1015 B.n757 B.n756 585
R1016 B.n755 B.n106 585
R1017 B.n754 B.n753 585
R1018 B.n752 B.n107 585
R1019 B.n751 B.n750 585
R1020 B.n749 B.n108 585
R1021 B.n748 B.n747 585
R1022 B.n746 B.n109 585
R1023 B.n745 B.n744 585
R1024 B.n743 B.n110 585
R1025 B.n742 B.n741 585
R1026 B.n740 B.n111 585
R1027 B.n739 B.n738 585
R1028 B.n737 B.n112 585
R1029 B.n736 B.n735 585
R1030 B.n734 B.n113 585
R1031 B.n733 B.n732 585
R1032 B.n731 B.n114 585
R1033 B.n730 B.n729 585
R1034 B.n728 B.n115 585
R1035 B.n727 B.n726 585
R1036 B.n725 B.n116 585
R1037 B.n724 B.n723 585
R1038 B.n722 B.n117 585
R1039 B.n721 B.n720 585
R1040 B.n719 B.n118 585
R1041 B.n718 B.n717 585
R1042 B.n716 B.n119 585
R1043 B.n715 B.n714 585
R1044 B.n713 B.n120 585
R1045 B.n712 B.n711 585
R1046 B.n710 B.n121 585
R1047 B.n709 B.n708 585
R1048 B.n707 B.n122 585
R1049 B.n706 B.n705 585
R1050 B.n704 B.n123 585
R1051 B.n703 B.n702 585
R1052 B.n701 B.n124 585
R1053 B.n700 B.n699 585
R1054 B.n698 B.n125 585
R1055 B.n697 B.n696 585
R1056 B.n695 B.n126 585
R1057 B.n694 B.n693 585
R1058 B.n692 B.n127 585
R1059 B.n691 B.n690 585
R1060 B.n689 B.n128 585
R1061 B.n688 B.n687 585
R1062 B.n686 B.n129 585
R1063 B.n685 B.n684 585
R1064 B.n683 B.n130 585
R1065 B.n682 B.n681 585
R1066 B.n680 B.n131 585
R1067 B.n679 B.n678 585
R1068 B.n677 B.n132 585
R1069 B.n676 B.n675 585
R1070 B.n674 B.n133 585
R1071 B.n673 B.n672 585
R1072 B.n671 B.n134 585
R1073 B.n670 B.n669 585
R1074 B.n668 B.n135 585
R1075 B.n667 B.n666 585
R1076 B.n665 B.n136 585
R1077 B.n664 B.n663 585
R1078 B.n662 B.n137 585
R1079 B.n661 B.n660 585
R1080 B.n659 B.n138 585
R1081 B.n658 B.n657 585
R1082 B.n656 B.n139 585
R1083 B.n655 B.n654 585
R1084 B.n653 B.n140 585
R1085 B.n652 B.n651 585
R1086 B.n650 B.n141 585
R1087 B.n649 B.n648 585
R1088 B.n647 B.n142 585
R1089 B.n646 B.n645 585
R1090 B.n644 B.n143 585
R1091 B.n643 B.n642 585
R1092 B.n641 B.n144 585
R1093 B.n640 B.n639 585
R1094 B.n638 B.n145 585
R1095 B.n637 B.n636 585
R1096 B.n635 B.n146 585
R1097 B.n634 B.n633 585
R1098 B.n632 B.n147 585
R1099 B.n631 B.n630 585
R1100 B.n629 B.n148 585
R1101 B.n628 B.n627 585
R1102 B.n626 B.n149 585
R1103 B.n625 B.n624 585
R1104 B.n623 B.n150 585
R1105 B.n622 B.n621 585
R1106 B.n620 B.n151 585
R1107 B.n619 B.n618 585
R1108 B.n617 B.n152 585
R1109 B.n616 B.n615 585
R1110 B.n614 B.n153 585
R1111 B.n613 B.n612 585
R1112 B.n611 B.n154 585
R1113 B.n610 B.n609 585
R1114 B.n608 B.n155 585
R1115 B.n607 B.n606 585
R1116 B.n605 B.n156 585
R1117 B.n604 B.n603 585
R1118 B.n602 B.n157 585
R1119 B.n601 B.n600 585
R1120 B.n599 B.n158 585
R1121 B.n598 B.n597 585
R1122 B.n596 B.n159 585
R1123 B.n595 B.n594 585
R1124 B.n593 B.n160 585
R1125 B.n592 B.n591 585
R1126 B.n590 B.n161 585
R1127 B.n589 B.n588 585
R1128 B.n587 B.n162 585
R1129 B.n586 B.n585 585
R1130 B.n584 B.n163 585
R1131 B.n583 B.n582 585
R1132 B.n581 B.n164 585
R1133 B.n580 B.n579 585
R1134 B.n578 B.n165 585
R1135 B.n577 B.n576 585
R1136 B.n575 B.n166 585
R1137 B.n574 B.n573 585
R1138 B.n572 B.n167 585
R1139 B.n571 B.n570 585
R1140 B.n569 B.n168 585
R1141 B.n568 B.n567 585
R1142 B.n566 B.n169 585
R1143 B.n565 B.n564 585
R1144 B.n563 B.n170 585
R1145 B.n562 B.n561 585
R1146 B.n560 B.n171 585
R1147 B.n559 B.n558 585
R1148 B.n557 B.n172 585
R1149 B.n556 B.n555 585
R1150 B.n554 B.n173 585
R1151 B.n553 B.n552 585
R1152 B.n551 B.n174 585
R1153 B.n550 B.n549 585
R1154 B.n548 B.n175 585
R1155 B.n547 B.n546 585
R1156 B.n545 B.n176 585
R1157 B.n544 B.n543 585
R1158 B.n542 B.n177 585
R1159 B.n391 B.n390 585
R1160 B.n392 B.n231 585
R1161 B.n394 B.n393 585
R1162 B.n395 B.n230 585
R1163 B.n397 B.n396 585
R1164 B.n398 B.n229 585
R1165 B.n400 B.n399 585
R1166 B.n401 B.n228 585
R1167 B.n403 B.n402 585
R1168 B.n404 B.n227 585
R1169 B.n406 B.n405 585
R1170 B.n407 B.n226 585
R1171 B.n409 B.n408 585
R1172 B.n410 B.n225 585
R1173 B.n412 B.n411 585
R1174 B.n413 B.n224 585
R1175 B.n415 B.n414 585
R1176 B.n416 B.n223 585
R1177 B.n418 B.n417 585
R1178 B.n419 B.n222 585
R1179 B.n421 B.n420 585
R1180 B.n422 B.n221 585
R1181 B.n424 B.n423 585
R1182 B.n425 B.n220 585
R1183 B.n427 B.n426 585
R1184 B.n428 B.n219 585
R1185 B.n430 B.n429 585
R1186 B.n431 B.n218 585
R1187 B.n433 B.n432 585
R1188 B.n434 B.n217 585
R1189 B.n436 B.n435 585
R1190 B.n437 B.n216 585
R1191 B.n439 B.n438 585
R1192 B.n440 B.n215 585
R1193 B.n442 B.n441 585
R1194 B.n443 B.n214 585
R1195 B.n445 B.n444 585
R1196 B.n446 B.n213 585
R1197 B.n448 B.n447 585
R1198 B.n449 B.n212 585
R1199 B.n451 B.n450 585
R1200 B.n452 B.n211 585
R1201 B.n454 B.n453 585
R1202 B.n455 B.n210 585
R1203 B.n457 B.n456 585
R1204 B.n459 B.n458 585
R1205 B.n460 B.n206 585
R1206 B.n462 B.n461 585
R1207 B.n463 B.n205 585
R1208 B.n465 B.n464 585
R1209 B.n466 B.n204 585
R1210 B.n468 B.n467 585
R1211 B.n469 B.n203 585
R1212 B.n471 B.n470 585
R1213 B.n472 B.n200 585
R1214 B.n475 B.n474 585
R1215 B.n476 B.n199 585
R1216 B.n478 B.n477 585
R1217 B.n479 B.n198 585
R1218 B.n481 B.n480 585
R1219 B.n482 B.n197 585
R1220 B.n484 B.n483 585
R1221 B.n485 B.n196 585
R1222 B.n487 B.n486 585
R1223 B.n488 B.n195 585
R1224 B.n490 B.n489 585
R1225 B.n491 B.n194 585
R1226 B.n493 B.n492 585
R1227 B.n494 B.n193 585
R1228 B.n496 B.n495 585
R1229 B.n497 B.n192 585
R1230 B.n499 B.n498 585
R1231 B.n500 B.n191 585
R1232 B.n502 B.n501 585
R1233 B.n503 B.n190 585
R1234 B.n505 B.n504 585
R1235 B.n506 B.n189 585
R1236 B.n508 B.n507 585
R1237 B.n509 B.n188 585
R1238 B.n511 B.n510 585
R1239 B.n512 B.n187 585
R1240 B.n514 B.n513 585
R1241 B.n515 B.n186 585
R1242 B.n517 B.n516 585
R1243 B.n518 B.n185 585
R1244 B.n520 B.n519 585
R1245 B.n521 B.n184 585
R1246 B.n523 B.n522 585
R1247 B.n524 B.n183 585
R1248 B.n526 B.n525 585
R1249 B.n527 B.n182 585
R1250 B.n529 B.n528 585
R1251 B.n530 B.n181 585
R1252 B.n532 B.n531 585
R1253 B.n533 B.n180 585
R1254 B.n535 B.n534 585
R1255 B.n536 B.n179 585
R1256 B.n538 B.n537 585
R1257 B.n539 B.n178 585
R1258 B.n541 B.n540 585
R1259 B.n389 B.n232 585
R1260 B.n388 B.n387 585
R1261 B.n386 B.n233 585
R1262 B.n385 B.n384 585
R1263 B.n383 B.n234 585
R1264 B.n382 B.n381 585
R1265 B.n380 B.n235 585
R1266 B.n379 B.n378 585
R1267 B.n377 B.n236 585
R1268 B.n376 B.n375 585
R1269 B.n374 B.n237 585
R1270 B.n373 B.n372 585
R1271 B.n371 B.n238 585
R1272 B.n370 B.n369 585
R1273 B.n368 B.n239 585
R1274 B.n367 B.n366 585
R1275 B.n365 B.n240 585
R1276 B.n364 B.n363 585
R1277 B.n362 B.n241 585
R1278 B.n361 B.n360 585
R1279 B.n359 B.n242 585
R1280 B.n358 B.n357 585
R1281 B.n356 B.n243 585
R1282 B.n355 B.n354 585
R1283 B.n353 B.n244 585
R1284 B.n352 B.n351 585
R1285 B.n350 B.n245 585
R1286 B.n349 B.n348 585
R1287 B.n347 B.n246 585
R1288 B.n346 B.n345 585
R1289 B.n344 B.n247 585
R1290 B.n343 B.n342 585
R1291 B.n341 B.n248 585
R1292 B.n340 B.n339 585
R1293 B.n338 B.n249 585
R1294 B.n337 B.n336 585
R1295 B.n335 B.n250 585
R1296 B.n334 B.n333 585
R1297 B.n332 B.n251 585
R1298 B.n331 B.n330 585
R1299 B.n329 B.n252 585
R1300 B.n328 B.n327 585
R1301 B.n326 B.n253 585
R1302 B.n325 B.n324 585
R1303 B.n323 B.n254 585
R1304 B.n322 B.n321 585
R1305 B.n320 B.n255 585
R1306 B.n319 B.n318 585
R1307 B.n317 B.n256 585
R1308 B.n316 B.n315 585
R1309 B.n314 B.n257 585
R1310 B.n313 B.n312 585
R1311 B.n311 B.n258 585
R1312 B.n310 B.n309 585
R1313 B.n308 B.n259 585
R1314 B.n307 B.n306 585
R1315 B.n305 B.n260 585
R1316 B.n304 B.n303 585
R1317 B.n302 B.n261 585
R1318 B.n301 B.n300 585
R1319 B.n299 B.n262 585
R1320 B.n298 B.n297 585
R1321 B.n296 B.n263 585
R1322 B.n295 B.n294 585
R1323 B.n293 B.n264 585
R1324 B.n292 B.n291 585
R1325 B.n290 B.n265 585
R1326 B.n289 B.n288 585
R1327 B.n287 B.n266 585
R1328 B.n286 B.n285 585
R1329 B.n284 B.n267 585
R1330 B.n283 B.n282 585
R1331 B.n281 B.n268 585
R1332 B.n280 B.n279 585
R1333 B.n278 B.n269 585
R1334 B.n277 B.n276 585
R1335 B.n275 B.n270 585
R1336 B.n274 B.n273 585
R1337 B.n272 B.n271 585
R1338 B.n2 B.n0 585
R1339 B.n1053 B.n1 585
R1340 B.n1052 B.n1051 585
R1341 B.n1050 B.n3 585
R1342 B.n1049 B.n1048 585
R1343 B.n1047 B.n4 585
R1344 B.n1046 B.n1045 585
R1345 B.n1044 B.n5 585
R1346 B.n1043 B.n1042 585
R1347 B.n1041 B.n6 585
R1348 B.n1040 B.n1039 585
R1349 B.n1038 B.n7 585
R1350 B.n1037 B.n1036 585
R1351 B.n1035 B.n8 585
R1352 B.n1034 B.n1033 585
R1353 B.n1032 B.n9 585
R1354 B.n1031 B.n1030 585
R1355 B.n1029 B.n10 585
R1356 B.n1028 B.n1027 585
R1357 B.n1026 B.n11 585
R1358 B.n1025 B.n1024 585
R1359 B.n1023 B.n12 585
R1360 B.n1022 B.n1021 585
R1361 B.n1020 B.n13 585
R1362 B.n1019 B.n1018 585
R1363 B.n1017 B.n14 585
R1364 B.n1016 B.n1015 585
R1365 B.n1014 B.n15 585
R1366 B.n1013 B.n1012 585
R1367 B.n1011 B.n16 585
R1368 B.n1010 B.n1009 585
R1369 B.n1008 B.n17 585
R1370 B.n1007 B.n1006 585
R1371 B.n1005 B.n18 585
R1372 B.n1004 B.n1003 585
R1373 B.n1002 B.n19 585
R1374 B.n1001 B.n1000 585
R1375 B.n999 B.n20 585
R1376 B.n998 B.n997 585
R1377 B.n996 B.n21 585
R1378 B.n995 B.n994 585
R1379 B.n993 B.n22 585
R1380 B.n992 B.n991 585
R1381 B.n990 B.n23 585
R1382 B.n989 B.n988 585
R1383 B.n987 B.n24 585
R1384 B.n986 B.n985 585
R1385 B.n984 B.n25 585
R1386 B.n983 B.n982 585
R1387 B.n981 B.n26 585
R1388 B.n980 B.n979 585
R1389 B.n978 B.n27 585
R1390 B.n977 B.n976 585
R1391 B.n975 B.n28 585
R1392 B.n974 B.n973 585
R1393 B.n972 B.n29 585
R1394 B.n971 B.n970 585
R1395 B.n969 B.n30 585
R1396 B.n968 B.n967 585
R1397 B.n966 B.n31 585
R1398 B.n965 B.n964 585
R1399 B.n963 B.n32 585
R1400 B.n962 B.n961 585
R1401 B.n960 B.n33 585
R1402 B.n959 B.n958 585
R1403 B.n957 B.n34 585
R1404 B.n956 B.n955 585
R1405 B.n954 B.n35 585
R1406 B.n953 B.n952 585
R1407 B.n951 B.n36 585
R1408 B.n950 B.n949 585
R1409 B.n948 B.n37 585
R1410 B.n947 B.n946 585
R1411 B.n945 B.n38 585
R1412 B.n944 B.n943 585
R1413 B.n942 B.n39 585
R1414 B.n941 B.n940 585
R1415 B.n939 B.n40 585
R1416 B.n938 B.n937 585
R1417 B.n936 B.n41 585
R1418 B.n935 B.n934 585
R1419 B.n1055 B.n1054 585
R1420 B.n391 B.n232 540.549
R1421 B.n934 B.n933 540.549
R1422 B.n542 B.n541 540.549
R1423 B.n783 B.n782 540.549
R1424 B.n201 B.t11 477.406
R1425 B.n73 B.t1 477.406
R1426 B.n207 B.t8 477.406
R1427 B.n66 B.t4 477.406
R1428 B.n202 B.t10 398.279
R1429 B.n74 B.t2 398.279
R1430 B.n208 B.t7 398.279
R1431 B.n67 B.t5 398.279
R1432 B.n201 B.t9 294.587
R1433 B.n207 B.t6 294.587
R1434 B.n66 B.t3 294.587
R1435 B.n73 B.t0 294.587
R1436 B.n387 B.n232 163.367
R1437 B.n387 B.n386 163.367
R1438 B.n386 B.n385 163.367
R1439 B.n385 B.n234 163.367
R1440 B.n381 B.n234 163.367
R1441 B.n381 B.n380 163.367
R1442 B.n380 B.n379 163.367
R1443 B.n379 B.n236 163.367
R1444 B.n375 B.n236 163.367
R1445 B.n375 B.n374 163.367
R1446 B.n374 B.n373 163.367
R1447 B.n373 B.n238 163.367
R1448 B.n369 B.n238 163.367
R1449 B.n369 B.n368 163.367
R1450 B.n368 B.n367 163.367
R1451 B.n367 B.n240 163.367
R1452 B.n363 B.n240 163.367
R1453 B.n363 B.n362 163.367
R1454 B.n362 B.n361 163.367
R1455 B.n361 B.n242 163.367
R1456 B.n357 B.n242 163.367
R1457 B.n357 B.n356 163.367
R1458 B.n356 B.n355 163.367
R1459 B.n355 B.n244 163.367
R1460 B.n351 B.n244 163.367
R1461 B.n351 B.n350 163.367
R1462 B.n350 B.n349 163.367
R1463 B.n349 B.n246 163.367
R1464 B.n345 B.n246 163.367
R1465 B.n345 B.n344 163.367
R1466 B.n344 B.n343 163.367
R1467 B.n343 B.n248 163.367
R1468 B.n339 B.n248 163.367
R1469 B.n339 B.n338 163.367
R1470 B.n338 B.n337 163.367
R1471 B.n337 B.n250 163.367
R1472 B.n333 B.n250 163.367
R1473 B.n333 B.n332 163.367
R1474 B.n332 B.n331 163.367
R1475 B.n331 B.n252 163.367
R1476 B.n327 B.n252 163.367
R1477 B.n327 B.n326 163.367
R1478 B.n326 B.n325 163.367
R1479 B.n325 B.n254 163.367
R1480 B.n321 B.n254 163.367
R1481 B.n321 B.n320 163.367
R1482 B.n320 B.n319 163.367
R1483 B.n319 B.n256 163.367
R1484 B.n315 B.n256 163.367
R1485 B.n315 B.n314 163.367
R1486 B.n314 B.n313 163.367
R1487 B.n313 B.n258 163.367
R1488 B.n309 B.n258 163.367
R1489 B.n309 B.n308 163.367
R1490 B.n308 B.n307 163.367
R1491 B.n307 B.n260 163.367
R1492 B.n303 B.n260 163.367
R1493 B.n303 B.n302 163.367
R1494 B.n302 B.n301 163.367
R1495 B.n301 B.n262 163.367
R1496 B.n297 B.n262 163.367
R1497 B.n297 B.n296 163.367
R1498 B.n296 B.n295 163.367
R1499 B.n295 B.n264 163.367
R1500 B.n291 B.n264 163.367
R1501 B.n291 B.n290 163.367
R1502 B.n290 B.n289 163.367
R1503 B.n289 B.n266 163.367
R1504 B.n285 B.n266 163.367
R1505 B.n285 B.n284 163.367
R1506 B.n284 B.n283 163.367
R1507 B.n283 B.n268 163.367
R1508 B.n279 B.n268 163.367
R1509 B.n279 B.n278 163.367
R1510 B.n278 B.n277 163.367
R1511 B.n277 B.n270 163.367
R1512 B.n273 B.n270 163.367
R1513 B.n273 B.n272 163.367
R1514 B.n272 B.n2 163.367
R1515 B.n1054 B.n2 163.367
R1516 B.n1054 B.n1053 163.367
R1517 B.n1053 B.n1052 163.367
R1518 B.n1052 B.n3 163.367
R1519 B.n1048 B.n3 163.367
R1520 B.n1048 B.n1047 163.367
R1521 B.n1047 B.n1046 163.367
R1522 B.n1046 B.n5 163.367
R1523 B.n1042 B.n5 163.367
R1524 B.n1042 B.n1041 163.367
R1525 B.n1041 B.n1040 163.367
R1526 B.n1040 B.n7 163.367
R1527 B.n1036 B.n7 163.367
R1528 B.n1036 B.n1035 163.367
R1529 B.n1035 B.n1034 163.367
R1530 B.n1034 B.n9 163.367
R1531 B.n1030 B.n9 163.367
R1532 B.n1030 B.n1029 163.367
R1533 B.n1029 B.n1028 163.367
R1534 B.n1028 B.n11 163.367
R1535 B.n1024 B.n11 163.367
R1536 B.n1024 B.n1023 163.367
R1537 B.n1023 B.n1022 163.367
R1538 B.n1022 B.n13 163.367
R1539 B.n1018 B.n13 163.367
R1540 B.n1018 B.n1017 163.367
R1541 B.n1017 B.n1016 163.367
R1542 B.n1016 B.n15 163.367
R1543 B.n1012 B.n15 163.367
R1544 B.n1012 B.n1011 163.367
R1545 B.n1011 B.n1010 163.367
R1546 B.n1010 B.n17 163.367
R1547 B.n1006 B.n17 163.367
R1548 B.n1006 B.n1005 163.367
R1549 B.n1005 B.n1004 163.367
R1550 B.n1004 B.n19 163.367
R1551 B.n1000 B.n19 163.367
R1552 B.n1000 B.n999 163.367
R1553 B.n999 B.n998 163.367
R1554 B.n998 B.n21 163.367
R1555 B.n994 B.n21 163.367
R1556 B.n994 B.n993 163.367
R1557 B.n993 B.n992 163.367
R1558 B.n992 B.n23 163.367
R1559 B.n988 B.n23 163.367
R1560 B.n988 B.n987 163.367
R1561 B.n987 B.n986 163.367
R1562 B.n986 B.n25 163.367
R1563 B.n982 B.n25 163.367
R1564 B.n982 B.n981 163.367
R1565 B.n981 B.n980 163.367
R1566 B.n980 B.n27 163.367
R1567 B.n976 B.n27 163.367
R1568 B.n976 B.n975 163.367
R1569 B.n975 B.n974 163.367
R1570 B.n974 B.n29 163.367
R1571 B.n970 B.n29 163.367
R1572 B.n970 B.n969 163.367
R1573 B.n969 B.n968 163.367
R1574 B.n968 B.n31 163.367
R1575 B.n964 B.n31 163.367
R1576 B.n964 B.n963 163.367
R1577 B.n963 B.n962 163.367
R1578 B.n962 B.n33 163.367
R1579 B.n958 B.n33 163.367
R1580 B.n958 B.n957 163.367
R1581 B.n957 B.n956 163.367
R1582 B.n956 B.n35 163.367
R1583 B.n952 B.n35 163.367
R1584 B.n952 B.n951 163.367
R1585 B.n951 B.n950 163.367
R1586 B.n950 B.n37 163.367
R1587 B.n946 B.n37 163.367
R1588 B.n946 B.n945 163.367
R1589 B.n945 B.n944 163.367
R1590 B.n944 B.n39 163.367
R1591 B.n940 B.n39 163.367
R1592 B.n940 B.n939 163.367
R1593 B.n939 B.n938 163.367
R1594 B.n938 B.n41 163.367
R1595 B.n934 B.n41 163.367
R1596 B.n392 B.n391 163.367
R1597 B.n393 B.n392 163.367
R1598 B.n393 B.n230 163.367
R1599 B.n397 B.n230 163.367
R1600 B.n398 B.n397 163.367
R1601 B.n399 B.n398 163.367
R1602 B.n399 B.n228 163.367
R1603 B.n403 B.n228 163.367
R1604 B.n404 B.n403 163.367
R1605 B.n405 B.n404 163.367
R1606 B.n405 B.n226 163.367
R1607 B.n409 B.n226 163.367
R1608 B.n410 B.n409 163.367
R1609 B.n411 B.n410 163.367
R1610 B.n411 B.n224 163.367
R1611 B.n415 B.n224 163.367
R1612 B.n416 B.n415 163.367
R1613 B.n417 B.n416 163.367
R1614 B.n417 B.n222 163.367
R1615 B.n421 B.n222 163.367
R1616 B.n422 B.n421 163.367
R1617 B.n423 B.n422 163.367
R1618 B.n423 B.n220 163.367
R1619 B.n427 B.n220 163.367
R1620 B.n428 B.n427 163.367
R1621 B.n429 B.n428 163.367
R1622 B.n429 B.n218 163.367
R1623 B.n433 B.n218 163.367
R1624 B.n434 B.n433 163.367
R1625 B.n435 B.n434 163.367
R1626 B.n435 B.n216 163.367
R1627 B.n439 B.n216 163.367
R1628 B.n440 B.n439 163.367
R1629 B.n441 B.n440 163.367
R1630 B.n441 B.n214 163.367
R1631 B.n445 B.n214 163.367
R1632 B.n446 B.n445 163.367
R1633 B.n447 B.n446 163.367
R1634 B.n447 B.n212 163.367
R1635 B.n451 B.n212 163.367
R1636 B.n452 B.n451 163.367
R1637 B.n453 B.n452 163.367
R1638 B.n453 B.n210 163.367
R1639 B.n457 B.n210 163.367
R1640 B.n458 B.n457 163.367
R1641 B.n458 B.n206 163.367
R1642 B.n462 B.n206 163.367
R1643 B.n463 B.n462 163.367
R1644 B.n464 B.n463 163.367
R1645 B.n464 B.n204 163.367
R1646 B.n468 B.n204 163.367
R1647 B.n469 B.n468 163.367
R1648 B.n470 B.n469 163.367
R1649 B.n470 B.n200 163.367
R1650 B.n475 B.n200 163.367
R1651 B.n476 B.n475 163.367
R1652 B.n477 B.n476 163.367
R1653 B.n477 B.n198 163.367
R1654 B.n481 B.n198 163.367
R1655 B.n482 B.n481 163.367
R1656 B.n483 B.n482 163.367
R1657 B.n483 B.n196 163.367
R1658 B.n487 B.n196 163.367
R1659 B.n488 B.n487 163.367
R1660 B.n489 B.n488 163.367
R1661 B.n489 B.n194 163.367
R1662 B.n493 B.n194 163.367
R1663 B.n494 B.n493 163.367
R1664 B.n495 B.n494 163.367
R1665 B.n495 B.n192 163.367
R1666 B.n499 B.n192 163.367
R1667 B.n500 B.n499 163.367
R1668 B.n501 B.n500 163.367
R1669 B.n501 B.n190 163.367
R1670 B.n505 B.n190 163.367
R1671 B.n506 B.n505 163.367
R1672 B.n507 B.n506 163.367
R1673 B.n507 B.n188 163.367
R1674 B.n511 B.n188 163.367
R1675 B.n512 B.n511 163.367
R1676 B.n513 B.n512 163.367
R1677 B.n513 B.n186 163.367
R1678 B.n517 B.n186 163.367
R1679 B.n518 B.n517 163.367
R1680 B.n519 B.n518 163.367
R1681 B.n519 B.n184 163.367
R1682 B.n523 B.n184 163.367
R1683 B.n524 B.n523 163.367
R1684 B.n525 B.n524 163.367
R1685 B.n525 B.n182 163.367
R1686 B.n529 B.n182 163.367
R1687 B.n530 B.n529 163.367
R1688 B.n531 B.n530 163.367
R1689 B.n531 B.n180 163.367
R1690 B.n535 B.n180 163.367
R1691 B.n536 B.n535 163.367
R1692 B.n537 B.n536 163.367
R1693 B.n537 B.n178 163.367
R1694 B.n541 B.n178 163.367
R1695 B.n543 B.n542 163.367
R1696 B.n543 B.n176 163.367
R1697 B.n547 B.n176 163.367
R1698 B.n548 B.n547 163.367
R1699 B.n549 B.n548 163.367
R1700 B.n549 B.n174 163.367
R1701 B.n553 B.n174 163.367
R1702 B.n554 B.n553 163.367
R1703 B.n555 B.n554 163.367
R1704 B.n555 B.n172 163.367
R1705 B.n559 B.n172 163.367
R1706 B.n560 B.n559 163.367
R1707 B.n561 B.n560 163.367
R1708 B.n561 B.n170 163.367
R1709 B.n565 B.n170 163.367
R1710 B.n566 B.n565 163.367
R1711 B.n567 B.n566 163.367
R1712 B.n567 B.n168 163.367
R1713 B.n571 B.n168 163.367
R1714 B.n572 B.n571 163.367
R1715 B.n573 B.n572 163.367
R1716 B.n573 B.n166 163.367
R1717 B.n577 B.n166 163.367
R1718 B.n578 B.n577 163.367
R1719 B.n579 B.n578 163.367
R1720 B.n579 B.n164 163.367
R1721 B.n583 B.n164 163.367
R1722 B.n584 B.n583 163.367
R1723 B.n585 B.n584 163.367
R1724 B.n585 B.n162 163.367
R1725 B.n589 B.n162 163.367
R1726 B.n590 B.n589 163.367
R1727 B.n591 B.n590 163.367
R1728 B.n591 B.n160 163.367
R1729 B.n595 B.n160 163.367
R1730 B.n596 B.n595 163.367
R1731 B.n597 B.n596 163.367
R1732 B.n597 B.n158 163.367
R1733 B.n601 B.n158 163.367
R1734 B.n602 B.n601 163.367
R1735 B.n603 B.n602 163.367
R1736 B.n603 B.n156 163.367
R1737 B.n607 B.n156 163.367
R1738 B.n608 B.n607 163.367
R1739 B.n609 B.n608 163.367
R1740 B.n609 B.n154 163.367
R1741 B.n613 B.n154 163.367
R1742 B.n614 B.n613 163.367
R1743 B.n615 B.n614 163.367
R1744 B.n615 B.n152 163.367
R1745 B.n619 B.n152 163.367
R1746 B.n620 B.n619 163.367
R1747 B.n621 B.n620 163.367
R1748 B.n621 B.n150 163.367
R1749 B.n625 B.n150 163.367
R1750 B.n626 B.n625 163.367
R1751 B.n627 B.n626 163.367
R1752 B.n627 B.n148 163.367
R1753 B.n631 B.n148 163.367
R1754 B.n632 B.n631 163.367
R1755 B.n633 B.n632 163.367
R1756 B.n633 B.n146 163.367
R1757 B.n637 B.n146 163.367
R1758 B.n638 B.n637 163.367
R1759 B.n639 B.n638 163.367
R1760 B.n639 B.n144 163.367
R1761 B.n643 B.n144 163.367
R1762 B.n644 B.n643 163.367
R1763 B.n645 B.n644 163.367
R1764 B.n645 B.n142 163.367
R1765 B.n649 B.n142 163.367
R1766 B.n650 B.n649 163.367
R1767 B.n651 B.n650 163.367
R1768 B.n651 B.n140 163.367
R1769 B.n655 B.n140 163.367
R1770 B.n656 B.n655 163.367
R1771 B.n657 B.n656 163.367
R1772 B.n657 B.n138 163.367
R1773 B.n661 B.n138 163.367
R1774 B.n662 B.n661 163.367
R1775 B.n663 B.n662 163.367
R1776 B.n663 B.n136 163.367
R1777 B.n667 B.n136 163.367
R1778 B.n668 B.n667 163.367
R1779 B.n669 B.n668 163.367
R1780 B.n669 B.n134 163.367
R1781 B.n673 B.n134 163.367
R1782 B.n674 B.n673 163.367
R1783 B.n675 B.n674 163.367
R1784 B.n675 B.n132 163.367
R1785 B.n679 B.n132 163.367
R1786 B.n680 B.n679 163.367
R1787 B.n681 B.n680 163.367
R1788 B.n681 B.n130 163.367
R1789 B.n685 B.n130 163.367
R1790 B.n686 B.n685 163.367
R1791 B.n687 B.n686 163.367
R1792 B.n687 B.n128 163.367
R1793 B.n691 B.n128 163.367
R1794 B.n692 B.n691 163.367
R1795 B.n693 B.n692 163.367
R1796 B.n693 B.n126 163.367
R1797 B.n697 B.n126 163.367
R1798 B.n698 B.n697 163.367
R1799 B.n699 B.n698 163.367
R1800 B.n699 B.n124 163.367
R1801 B.n703 B.n124 163.367
R1802 B.n704 B.n703 163.367
R1803 B.n705 B.n704 163.367
R1804 B.n705 B.n122 163.367
R1805 B.n709 B.n122 163.367
R1806 B.n710 B.n709 163.367
R1807 B.n711 B.n710 163.367
R1808 B.n711 B.n120 163.367
R1809 B.n715 B.n120 163.367
R1810 B.n716 B.n715 163.367
R1811 B.n717 B.n716 163.367
R1812 B.n717 B.n118 163.367
R1813 B.n721 B.n118 163.367
R1814 B.n722 B.n721 163.367
R1815 B.n723 B.n722 163.367
R1816 B.n723 B.n116 163.367
R1817 B.n727 B.n116 163.367
R1818 B.n728 B.n727 163.367
R1819 B.n729 B.n728 163.367
R1820 B.n729 B.n114 163.367
R1821 B.n733 B.n114 163.367
R1822 B.n734 B.n733 163.367
R1823 B.n735 B.n734 163.367
R1824 B.n735 B.n112 163.367
R1825 B.n739 B.n112 163.367
R1826 B.n740 B.n739 163.367
R1827 B.n741 B.n740 163.367
R1828 B.n741 B.n110 163.367
R1829 B.n745 B.n110 163.367
R1830 B.n746 B.n745 163.367
R1831 B.n747 B.n746 163.367
R1832 B.n747 B.n108 163.367
R1833 B.n751 B.n108 163.367
R1834 B.n752 B.n751 163.367
R1835 B.n753 B.n752 163.367
R1836 B.n753 B.n106 163.367
R1837 B.n757 B.n106 163.367
R1838 B.n758 B.n757 163.367
R1839 B.n759 B.n758 163.367
R1840 B.n759 B.n104 163.367
R1841 B.n763 B.n104 163.367
R1842 B.n764 B.n763 163.367
R1843 B.n765 B.n764 163.367
R1844 B.n765 B.n102 163.367
R1845 B.n769 B.n102 163.367
R1846 B.n770 B.n769 163.367
R1847 B.n771 B.n770 163.367
R1848 B.n771 B.n100 163.367
R1849 B.n775 B.n100 163.367
R1850 B.n776 B.n775 163.367
R1851 B.n777 B.n776 163.367
R1852 B.n777 B.n98 163.367
R1853 B.n781 B.n98 163.367
R1854 B.n782 B.n781 163.367
R1855 B.n933 B.n932 163.367
R1856 B.n932 B.n43 163.367
R1857 B.n928 B.n43 163.367
R1858 B.n928 B.n927 163.367
R1859 B.n927 B.n926 163.367
R1860 B.n926 B.n45 163.367
R1861 B.n922 B.n45 163.367
R1862 B.n922 B.n921 163.367
R1863 B.n921 B.n920 163.367
R1864 B.n920 B.n47 163.367
R1865 B.n916 B.n47 163.367
R1866 B.n916 B.n915 163.367
R1867 B.n915 B.n914 163.367
R1868 B.n914 B.n49 163.367
R1869 B.n910 B.n49 163.367
R1870 B.n910 B.n909 163.367
R1871 B.n909 B.n908 163.367
R1872 B.n908 B.n51 163.367
R1873 B.n904 B.n51 163.367
R1874 B.n904 B.n903 163.367
R1875 B.n903 B.n902 163.367
R1876 B.n902 B.n53 163.367
R1877 B.n898 B.n53 163.367
R1878 B.n898 B.n897 163.367
R1879 B.n897 B.n896 163.367
R1880 B.n896 B.n55 163.367
R1881 B.n892 B.n55 163.367
R1882 B.n892 B.n891 163.367
R1883 B.n891 B.n890 163.367
R1884 B.n890 B.n57 163.367
R1885 B.n886 B.n57 163.367
R1886 B.n886 B.n885 163.367
R1887 B.n885 B.n884 163.367
R1888 B.n884 B.n59 163.367
R1889 B.n880 B.n59 163.367
R1890 B.n880 B.n879 163.367
R1891 B.n879 B.n878 163.367
R1892 B.n878 B.n61 163.367
R1893 B.n874 B.n61 163.367
R1894 B.n874 B.n873 163.367
R1895 B.n873 B.n872 163.367
R1896 B.n872 B.n63 163.367
R1897 B.n868 B.n63 163.367
R1898 B.n868 B.n867 163.367
R1899 B.n867 B.n866 163.367
R1900 B.n866 B.n65 163.367
R1901 B.n862 B.n65 163.367
R1902 B.n862 B.n861 163.367
R1903 B.n861 B.n860 163.367
R1904 B.n860 B.n70 163.367
R1905 B.n856 B.n70 163.367
R1906 B.n856 B.n855 163.367
R1907 B.n855 B.n854 163.367
R1908 B.n854 B.n72 163.367
R1909 B.n849 B.n72 163.367
R1910 B.n849 B.n848 163.367
R1911 B.n848 B.n847 163.367
R1912 B.n847 B.n76 163.367
R1913 B.n843 B.n76 163.367
R1914 B.n843 B.n842 163.367
R1915 B.n842 B.n841 163.367
R1916 B.n841 B.n78 163.367
R1917 B.n837 B.n78 163.367
R1918 B.n837 B.n836 163.367
R1919 B.n836 B.n835 163.367
R1920 B.n835 B.n80 163.367
R1921 B.n831 B.n80 163.367
R1922 B.n831 B.n830 163.367
R1923 B.n830 B.n829 163.367
R1924 B.n829 B.n82 163.367
R1925 B.n825 B.n82 163.367
R1926 B.n825 B.n824 163.367
R1927 B.n824 B.n823 163.367
R1928 B.n823 B.n84 163.367
R1929 B.n819 B.n84 163.367
R1930 B.n819 B.n818 163.367
R1931 B.n818 B.n817 163.367
R1932 B.n817 B.n86 163.367
R1933 B.n813 B.n86 163.367
R1934 B.n813 B.n812 163.367
R1935 B.n812 B.n811 163.367
R1936 B.n811 B.n88 163.367
R1937 B.n807 B.n88 163.367
R1938 B.n807 B.n806 163.367
R1939 B.n806 B.n805 163.367
R1940 B.n805 B.n90 163.367
R1941 B.n801 B.n90 163.367
R1942 B.n801 B.n800 163.367
R1943 B.n800 B.n799 163.367
R1944 B.n799 B.n92 163.367
R1945 B.n795 B.n92 163.367
R1946 B.n795 B.n794 163.367
R1947 B.n794 B.n793 163.367
R1948 B.n793 B.n94 163.367
R1949 B.n789 B.n94 163.367
R1950 B.n789 B.n788 163.367
R1951 B.n788 B.n787 163.367
R1952 B.n787 B.n96 163.367
R1953 B.n783 B.n96 163.367
R1954 B.n202 B.n201 79.1278
R1955 B.n208 B.n207 79.1278
R1956 B.n67 B.n66 79.1278
R1957 B.n74 B.n73 79.1278
R1958 B.n473 B.n202 59.5399
R1959 B.n209 B.n208 59.5399
R1960 B.n68 B.n67 59.5399
R1961 B.n851 B.n74 59.5399
R1962 B.n935 B.n42 35.1225
R1963 B.n540 B.n177 35.1225
R1964 B.n390 B.n389 35.1225
R1965 B.n784 B.n97 35.1224
R1966 B B.n1055 18.0485
R1967 B.n931 B.n42 10.6151
R1968 B.n931 B.n930 10.6151
R1969 B.n930 B.n929 10.6151
R1970 B.n929 B.n44 10.6151
R1971 B.n925 B.n44 10.6151
R1972 B.n925 B.n924 10.6151
R1973 B.n924 B.n923 10.6151
R1974 B.n923 B.n46 10.6151
R1975 B.n919 B.n46 10.6151
R1976 B.n919 B.n918 10.6151
R1977 B.n918 B.n917 10.6151
R1978 B.n917 B.n48 10.6151
R1979 B.n913 B.n48 10.6151
R1980 B.n913 B.n912 10.6151
R1981 B.n912 B.n911 10.6151
R1982 B.n911 B.n50 10.6151
R1983 B.n907 B.n50 10.6151
R1984 B.n907 B.n906 10.6151
R1985 B.n906 B.n905 10.6151
R1986 B.n905 B.n52 10.6151
R1987 B.n901 B.n52 10.6151
R1988 B.n901 B.n900 10.6151
R1989 B.n900 B.n899 10.6151
R1990 B.n899 B.n54 10.6151
R1991 B.n895 B.n54 10.6151
R1992 B.n895 B.n894 10.6151
R1993 B.n894 B.n893 10.6151
R1994 B.n893 B.n56 10.6151
R1995 B.n889 B.n56 10.6151
R1996 B.n889 B.n888 10.6151
R1997 B.n888 B.n887 10.6151
R1998 B.n887 B.n58 10.6151
R1999 B.n883 B.n58 10.6151
R2000 B.n883 B.n882 10.6151
R2001 B.n882 B.n881 10.6151
R2002 B.n881 B.n60 10.6151
R2003 B.n877 B.n60 10.6151
R2004 B.n877 B.n876 10.6151
R2005 B.n876 B.n875 10.6151
R2006 B.n875 B.n62 10.6151
R2007 B.n871 B.n62 10.6151
R2008 B.n871 B.n870 10.6151
R2009 B.n870 B.n869 10.6151
R2010 B.n869 B.n64 10.6151
R2011 B.n865 B.n864 10.6151
R2012 B.n864 B.n863 10.6151
R2013 B.n863 B.n69 10.6151
R2014 B.n859 B.n69 10.6151
R2015 B.n859 B.n858 10.6151
R2016 B.n858 B.n857 10.6151
R2017 B.n857 B.n71 10.6151
R2018 B.n853 B.n71 10.6151
R2019 B.n853 B.n852 10.6151
R2020 B.n850 B.n75 10.6151
R2021 B.n846 B.n75 10.6151
R2022 B.n846 B.n845 10.6151
R2023 B.n845 B.n844 10.6151
R2024 B.n844 B.n77 10.6151
R2025 B.n840 B.n77 10.6151
R2026 B.n840 B.n839 10.6151
R2027 B.n839 B.n838 10.6151
R2028 B.n838 B.n79 10.6151
R2029 B.n834 B.n79 10.6151
R2030 B.n834 B.n833 10.6151
R2031 B.n833 B.n832 10.6151
R2032 B.n832 B.n81 10.6151
R2033 B.n828 B.n81 10.6151
R2034 B.n828 B.n827 10.6151
R2035 B.n827 B.n826 10.6151
R2036 B.n826 B.n83 10.6151
R2037 B.n822 B.n83 10.6151
R2038 B.n822 B.n821 10.6151
R2039 B.n821 B.n820 10.6151
R2040 B.n820 B.n85 10.6151
R2041 B.n816 B.n85 10.6151
R2042 B.n816 B.n815 10.6151
R2043 B.n815 B.n814 10.6151
R2044 B.n814 B.n87 10.6151
R2045 B.n810 B.n87 10.6151
R2046 B.n810 B.n809 10.6151
R2047 B.n809 B.n808 10.6151
R2048 B.n808 B.n89 10.6151
R2049 B.n804 B.n89 10.6151
R2050 B.n804 B.n803 10.6151
R2051 B.n803 B.n802 10.6151
R2052 B.n802 B.n91 10.6151
R2053 B.n798 B.n91 10.6151
R2054 B.n798 B.n797 10.6151
R2055 B.n797 B.n796 10.6151
R2056 B.n796 B.n93 10.6151
R2057 B.n792 B.n93 10.6151
R2058 B.n792 B.n791 10.6151
R2059 B.n791 B.n790 10.6151
R2060 B.n790 B.n95 10.6151
R2061 B.n786 B.n95 10.6151
R2062 B.n786 B.n785 10.6151
R2063 B.n785 B.n784 10.6151
R2064 B.n544 B.n177 10.6151
R2065 B.n545 B.n544 10.6151
R2066 B.n546 B.n545 10.6151
R2067 B.n546 B.n175 10.6151
R2068 B.n550 B.n175 10.6151
R2069 B.n551 B.n550 10.6151
R2070 B.n552 B.n551 10.6151
R2071 B.n552 B.n173 10.6151
R2072 B.n556 B.n173 10.6151
R2073 B.n557 B.n556 10.6151
R2074 B.n558 B.n557 10.6151
R2075 B.n558 B.n171 10.6151
R2076 B.n562 B.n171 10.6151
R2077 B.n563 B.n562 10.6151
R2078 B.n564 B.n563 10.6151
R2079 B.n564 B.n169 10.6151
R2080 B.n568 B.n169 10.6151
R2081 B.n569 B.n568 10.6151
R2082 B.n570 B.n569 10.6151
R2083 B.n570 B.n167 10.6151
R2084 B.n574 B.n167 10.6151
R2085 B.n575 B.n574 10.6151
R2086 B.n576 B.n575 10.6151
R2087 B.n576 B.n165 10.6151
R2088 B.n580 B.n165 10.6151
R2089 B.n581 B.n580 10.6151
R2090 B.n582 B.n581 10.6151
R2091 B.n582 B.n163 10.6151
R2092 B.n586 B.n163 10.6151
R2093 B.n587 B.n586 10.6151
R2094 B.n588 B.n587 10.6151
R2095 B.n588 B.n161 10.6151
R2096 B.n592 B.n161 10.6151
R2097 B.n593 B.n592 10.6151
R2098 B.n594 B.n593 10.6151
R2099 B.n594 B.n159 10.6151
R2100 B.n598 B.n159 10.6151
R2101 B.n599 B.n598 10.6151
R2102 B.n600 B.n599 10.6151
R2103 B.n600 B.n157 10.6151
R2104 B.n604 B.n157 10.6151
R2105 B.n605 B.n604 10.6151
R2106 B.n606 B.n605 10.6151
R2107 B.n606 B.n155 10.6151
R2108 B.n610 B.n155 10.6151
R2109 B.n611 B.n610 10.6151
R2110 B.n612 B.n611 10.6151
R2111 B.n612 B.n153 10.6151
R2112 B.n616 B.n153 10.6151
R2113 B.n617 B.n616 10.6151
R2114 B.n618 B.n617 10.6151
R2115 B.n618 B.n151 10.6151
R2116 B.n622 B.n151 10.6151
R2117 B.n623 B.n622 10.6151
R2118 B.n624 B.n623 10.6151
R2119 B.n624 B.n149 10.6151
R2120 B.n628 B.n149 10.6151
R2121 B.n629 B.n628 10.6151
R2122 B.n630 B.n629 10.6151
R2123 B.n630 B.n147 10.6151
R2124 B.n634 B.n147 10.6151
R2125 B.n635 B.n634 10.6151
R2126 B.n636 B.n635 10.6151
R2127 B.n636 B.n145 10.6151
R2128 B.n640 B.n145 10.6151
R2129 B.n641 B.n640 10.6151
R2130 B.n642 B.n641 10.6151
R2131 B.n642 B.n143 10.6151
R2132 B.n646 B.n143 10.6151
R2133 B.n647 B.n646 10.6151
R2134 B.n648 B.n647 10.6151
R2135 B.n648 B.n141 10.6151
R2136 B.n652 B.n141 10.6151
R2137 B.n653 B.n652 10.6151
R2138 B.n654 B.n653 10.6151
R2139 B.n654 B.n139 10.6151
R2140 B.n658 B.n139 10.6151
R2141 B.n659 B.n658 10.6151
R2142 B.n660 B.n659 10.6151
R2143 B.n660 B.n137 10.6151
R2144 B.n664 B.n137 10.6151
R2145 B.n665 B.n664 10.6151
R2146 B.n666 B.n665 10.6151
R2147 B.n666 B.n135 10.6151
R2148 B.n670 B.n135 10.6151
R2149 B.n671 B.n670 10.6151
R2150 B.n672 B.n671 10.6151
R2151 B.n672 B.n133 10.6151
R2152 B.n676 B.n133 10.6151
R2153 B.n677 B.n676 10.6151
R2154 B.n678 B.n677 10.6151
R2155 B.n678 B.n131 10.6151
R2156 B.n682 B.n131 10.6151
R2157 B.n683 B.n682 10.6151
R2158 B.n684 B.n683 10.6151
R2159 B.n684 B.n129 10.6151
R2160 B.n688 B.n129 10.6151
R2161 B.n689 B.n688 10.6151
R2162 B.n690 B.n689 10.6151
R2163 B.n690 B.n127 10.6151
R2164 B.n694 B.n127 10.6151
R2165 B.n695 B.n694 10.6151
R2166 B.n696 B.n695 10.6151
R2167 B.n696 B.n125 10.6151
R2168 B.n700 B.n125 10.6151
R2169 B.n701 B.n700 10.6151
R2170 B.n702 B.n701 10.6151
R2171 B.n702 B.n123 10.6151
R2172 B.n706 B.n123 10.6151
R2173 B.n707 B.n706 10.6151
R2174 B.n708 B.n707 10.6151
R2175 B.n708 B.n121 10.6151
R2176 B.n712 B.n121 10.6151
R2177 B.n713 B.n712 10.6151
R2178 B.n714 B.n713 10.6151
R2179 B.n714 B.n119 10.6151
R2180 B.n718 B.n119 10.6151
R2181 B.n719 B.n718 10.6151
R2182 B.n720 B.n719 10.6151
R2183 B.n720 B.n117 10.6151
R2184 B.n724 B.n117 10.6151
R2185 B.n725 B.n724 10.6151
R2186 B.n726 B.n725 10.6151
R2187 B.n726 B.n115 10.6151
R2188 B.n730 B.n115 10.6151
R2189 B.n731 B.n730 10.6151
R2190 B.n732 B.n731 10.6151
R2191 B.n732 B.n113 10.6151
R2192 B.n736 B.n113 10.6151
R2193 B.n737 B.n736 10.6151
R2194 B.n738 B.n737 10.6151
R2195 B.n738 B.n111 10.6151
R2196 B.n742 B.n111 10.6151
R2197 B.n743 B.n742 10.6151
R2198 B.n744 B.n743 10.6151
R2199 B.n744 B.n109 10.6151
R2200 B.n748 B.n109 10.6151
R2201 B.n749 B.n748 10.6151
R2202 B.n750 B.n749 10.6151
R2203 B.n750 B.n107 10.6151
R2204 B.n754 B.n107 10.6151
R2205 B.n755 B.n754 10.6151
R2206 B.n756 B.n755 10.6151
R2207 B.n756 B.n105 10.6151
R2208 B.n760 B.n105 10.6151
R2209 B.n761 B.n760 10.6151
R2210 B.n762 B.n761 10.6151
R2211 B.n762 B.n103 10.6151
R2212 B.n766 B.n103 10.6151
R2213 B.n767 B.n766 10.6151
R2214 B.n768 B.n767 10.6151
R2215 B.n768 B.n101 10.6151
R2216 B.n772 B.n101 10.6151
R2217 B.n773 B.n772 10.6151
R2218 B.n774 B.n773 10.6151
R2219 B.n774 B.n99 10.6151
R2220 B.n778 B.n99 10.6151
R2221 B.n779 B.n778 10.6151
R2222 B.n780 B.n779 10.6151
R2223 B.n780 B.n97 10.6151
R2224 B.n390 B.n231 10.6151
R2225 B.n394 B.n231 10.6151
R2226 B.n395 B.n394 10.6151
R2227 B.n396 B.n395 10.6151
R2228 B.n396 B.n229 10.6151
R2229 B.n400 B.n229 10.6151
R2230 B.n401 B.n400 10.6151
R2231 B.n402 B.n401 10.6151
R2232 B.n402 B.n227 10.6151
R2233 B.n406 B.n227 10.6151
R2234 B.n407 B.n406 10.6151
R2235 B.n408 B.n407 10.6151
R2236 B.n408 B.n225 10.6151
R2237 B.n412 B.n225 10.6151
R2238 B.n413 B.n412 10.6151
R2239 B.n414 B.n413 10.6151
R2240 B.n414 B.n223 10.6151
R2241 B.n418 B.n223 10.6151
R2242 B.n419 B.n418 10.6151
R2243 B.n420 B.n419 10.6151
R2244 B.n420 B.n221 10.6151
R2245 B.n424 B.n221 10.6151
R2246 B.n425 B.n424 10.6151
R2247 B.n426 B.n425 10.6151
R2248 B.n426 B.n219 10.6151
R2249 B.n430 B.n219 10.6151
R2250 B.n431 B.n430 10.6151
R2251 B.n432 B.n431 10.6151
R2252 B.n432 B.n217 10.6151
R2253 B.n436 B.n217 10.6151
R2254 B.n437 B.n436 10.6151
R2255 B.n438 B.n437 10.6151
R2256 B.n438 B.n215 10.6151
R2257 B.n442 B.n215 10.6151
R2258 B.n443 B.n442 10.6151
R2259 B.n444 B.n443 10.6151
R2260 B.n444 B.n213 10.6151
R2261 B.n448 B.n213 10.6151
R2262 B.n449 B.n448 10.6151
R2263 B.n450 B.n449 10.6151
R2264 B.n450 B.n211 10.6151
R2265 B.n454 B.n211 10.6151
R2266 B.n455 B.n454 10.6151
R2267 B.n456 B.n455 10.6151
R2268 B.n460 B.n459 10.6151
R2269 B.n461 B.n460 10.6151
R2270 B.n461 B.n205 10.6151
R2271 B.n465 B.n205 10.6151
R2272 B.n466 B.n465 10.6151
R2273 B.n467 B.n466 10.6151
R2274 B.n467 B.n203 10.6151
R2275 B.n471 B.n203 10.6151
R2276 B.n472 B.n471 10.6151
R2277 B.n474 B.n199 10.6151
R2278 B.n478 B.n199 10.6151
R2279 B.n479 B.n478 10.6151
R2280 B.n480 B.n479 10.6151
R2281 B.n480 B.n197 10.6151
R2282 B.n484 B.n197 10.6151
R2283 B.n485 B.n484 10.6151
R2284 B.n486 B.n485 10.6151
R2285 B.n486 B.n195 10.6151
R2286 B.n490 B.n195 10.6151
R2287 B.n491 B.n490 10.6151
R2288 B.n492 B.n491 10.6151
R2289 B.n492 B.n193 10.6151
R2290 B.n496 B.n193 10.6151
R2291 B.n497 B.n496 10.6151
R2292 B.n498 B.n497 10.6151
R2293 B.n498 B.n191 10.6151
R2294 B.n502 B.n191 10.6151
R2295 B.n503 B.n502 10.6151
R2296 B.n504 B.n503 10.6151
R2297 B.n504 B.n189 10.6151
R2298 B.n508 B.n189 10.6151
R2299 B.n509 B.n508 10.6151
R2300 B.n510 B.n509 10.6151
R2301 B.n510 B.n187 10.6151
R2302 B.n514 B.n187 10.6151
R2303 B.n515 B.n514 10.6151
R2304 B.n516 B.n515 10.6151
R2305 B.n516 B.n185 10.6151
R2306 B.n520 B.n185 10.6151
R2307 B.n521 B.n520 10.6151
R2308 B.n522 B.n521 10.6151
R2309 B.n522 B.n183 10.6151
R2310 B.n526 B.n183 10.6151
R2311 B.n527 B.n526 10.6151
R2312 B.n528 B.n527 10.6151
R2313 B.n528 B.n181 10.6151
R2314 B.n532 B.n181 10.6151
R2315 B.n533 B.n532 10.6151
R2316 B.n534 B.n533 10.6151
R2317 B.n534 B.n179 10.6151
R2318 B.n538 B.n179 10.6151
R2319 B.n539 B.n538 10.6151
R2320 B.n540 B.n539 10.6151
R2321 B.n389 B.n388 10.6151
R2322 B.n388 B.n233 10.6151
R2323 B.n384 B.n233 10.6151
R2324 B.n384 B.n383 10.6151
R2325 B.n383 B.n382 10.6151
R2326 B.n382 B.n235 10.6151
R2327 B.n378 B.n235 10.6151
R2328 B.n378 B.n377 10.6151
R2329 B.n377 B.n376 10.6151
R2330 B.n376 B.n237 10.6151
R2331 B.n372 B.n237 10.6151
R2332 B.n372 B.n371 10.6151
R2333 B.n371 B.n370 10.6151
R2334 B.n370 B.n239 10.6151
R2335 B.n366 B.n239 10.6151
R2336 B.n366 B.n365 10.6151
R2337 B.n365 B.n364 10.6151
R2338 B.n364 B.n241 10.6151
R2339 B.n360 B.n241 10.6151
R2340 B.n360 B.n359 10.6151
R2341 B.n359 B.n358 10.6151
R2342 B.n358 B.n243 10.6151
R2343 B.n354 B.n243 10.6151
R2344 B.n354 B.n353 10.6151
R2345 B.n353 B.n352 10.6151
R2346 B.n352 B.n245 10.6151
R2347 B.n348 B.n245 10.6151
R2348 B.n348 B.n347 10.6151
R2349 B.n347 B.n346 10.6151
R2350 B.n346 B.n247 10.6151
R2351 B.n342 B.n247 10.6151
R2352 B.n342 B.n341 10.6151
R2353 B.n341 B.n340 10.6151
R2354 B.n340 B.n249 10.6151
R2355 B.n336 B.n249 10.6151
R2356 B.n336 B.n335 10.6151
R2357 B.n335 B.n334 10.6151
R2358 B.n334 B.n251 10.6151
R2359 B.n330 B.n251 10.6151
R2360 B.n330 B.n329 10.6151
R2361 B.n329 B.n328 10.6151
R2362 B.n328 B.n253 10.6151
R2363 B.n324 B.n253 10.6151
R2364 B.n324 B.n323 10.6151
R2365 B.n323 B.n322 10.6151
R2366 B.n322 B.n255 10.6151
R2367 B.n318 B.n255 10.6151
R2368 B.n318 B.n317 10.6151
R2369 B.n317 B.n316 10.6151
R2370 B.n316 B.n257 10.6151
R2371 B.n312 B.n257 10.6151
R2372 B.n312 B.n311 10.6151
R2373 B.n311 B.n310 10.6151
R2374 B.n310 B.n259 10.6151
R2375 B.n306 B.n259 10.6151
R2376 B.n306 B.n305 10.6151
R2377 B.n305 B.n304 10.6151
R2378 B.n304 B.n261 10.6151
R2379 B.n300 B.n261 10.6151
R2380 B.n300 B.n299 10.6151
R2381 B.n299 B.n298 10.6151
R2382 B.n298 B.n263 10.6151
R2383 B.n294 B.n263 10.6151
R2384 B.n294 B.n293 10.6151
R2385 B.n293 B.n292 10.6151
R2386 B.n292 B.n265 10.6151
R2387 B.n288 B.n265 10.6151
R2388 B.n288 B.n287 10.6151
R2389 B.n287 B.n286 10.6151
R2390 B.n286 B.n267 10.6151
R2391 B.n282 B.n267 10.6151
R2392 B.n282 B.n281 10.6151
R2393 B.n281 B.n280 10.6151
R2394 B.n280 B.n269 10.6151
R2395 B.n276 B.n269 10.6151
R2396 B.n276 B.n275 10.6151
R2397 B.n275 B.n274 10.6151
R2398 B.n274 B.n271 10.6151
R2399 B.n271 B.n0 10.6151
R2400 B.n1051 B.n1 10.6151
R2401 B.n1051 B.n1050 10.6151
R2402 B.n1050 B.n1049 10.6151
R2403 B.n1049 B.n4 10.6151
R2404 B.n1045 B.n4 10.6151
R2405 B.n1045 B.n1044 10.6151
R2406 B.n1044 B.n1043 10.6151
R2407 B.n1043 B.n6 10.6151
R2408 B.n1039 B.n6 10.6151
R2409 B.n1039 B.n1038 10.6151
R2410 B.n1038 B.n1037 10.6151
R2411 B.n1037 B.n8 10.6151
R2412 B.n1033 B.n8 10.6151
R2413 B.n1033 B.n1032 10.6151
R2414 B.n1032 B.n1031 10.6151
R2415 B.n1031 B.n10 10.6151
R2416 B.n1027 B.n10 10.6151
R2417 B.n1027 B.n1026 10.6151
R2418 B.n1026 B.n1025 10.6151
R2419 B.n1025 B.n12 10.6151
R2420 B.n1021 B.n12 10.6151
R2421 B.n1021 B.n1020 10.6151
R2422 B.n1020 B.n1019 10.6151
R2423 B.n1019 B.n14 10.6151
R2424 B.n1015 B.n14 10.6151
R2425 B.n1015 B.n1014 10.6151
R2426 B.n1014 B.n1013 10.6151
R2427 B.n1013 B.n16 10.6151
R2428 B.n1009 B.n16 10.6151
R2429 B.n1009 B.n1008 10.6151
R2430 B.n1008 B.n1007 10.6151
R2431 B.n1007 B.n18 10.6151
R2432 B.n1003 B.n18 10.6151
R2433 B.n1003 B.n1002 10.6151
R2434 B.n1002 B.n1001 10.6151
R2435 B.n1001 B.n20 10.6151
R2436 B.n997 B.n20 10.6151
R2437 B.n997 B.n996 10.6151
R2438 B.n996 B.n995 10.6151
R2439 B.n995 B.n22 10.6151
R2440 B.n991 B.n22 10.6151
R2441 B.n991 B.n990 10.6151
R2442 B.n990 B.n989 10.6151
R2443 B.n989 B.n24 10.6151
R2444 B.n985 B.n24 10.6151
R2445 B.n985 B.n984 10.6151
R2446 B.n984 B.n983 10.6151
R2447 B.n983 B.n26 10.6151
R2448 B.n979 B.n26 10.6151
R2449 B.n979 B.n978 10.6151
R2450 B.n978 B.n977 10.6151
R2451 B.n977 B.n28 10.6151
R2452 B.n973 B.n28 10.6151
R2453 B.n973 B.n972 10.6151
R2454 B.n972 B.n971 10.6151
R2455 B.n971 B.n30 10.6151
R2456 B.n967 B.n30 10.6151
R2457 B.n967 B.n966 10.6151
R2458 B.n966 B.n965 10.6151
R2459 B.n965 B.n32 10.6151
R2460 B.n961 B.n32 10.6151
R2461 B.n961 B.n960 10.6151
R2462 B.n960 B.n959 10.6151
R2463 B.n959 B.n34 10.6151
R2464 B.n955 B.n34 10.6151
R2465 B.n955 B.n954 10.6151
R2466 B.n954 B.n953 10.6151
R2467 B.n953 B.n36 10.6151
R2468 B.n949 B.n36 10.6151
R2469 B.n949 B.n948 10.6151
R2470 B.n948 B.n947 10.6151
R2471 B.n947 B.n38 10.6151
R2472 B.n943 B.n38 10.6151
R2473 B.n943 B.n942 10.6151
R2474 B.n942 B.n941 10.6151
R2475 B.n941 B.n40 10.6151
R2476 B.n937 B.n40 10.6151
R2477 B.n937 B.n936 10.6151
R2478 B.n936 B.n935 10.6151
R2479 B.n68 B.n64 9.36635
R2480 B.n851 B.n850 9.36635
R2481 B.n456 B.n209 9.36635
R2482 B.n474 B.n473 9.36635
R2483 B.n1055 B.n0 2.81026
R2484 B.n1055 B.n1 2.81026
R2485 B.n865 B.n68 1.24928
R2486 B.n852 B.n851 1.24928
R2487 B.n459 B.n209 1.24928
R2488 B.n473 B.n472 1.24928
R2489 VN.n108 VN.n107 161.3
R2490 VN.n106 VN.n56 161.3
R2491 VN.n105 VN.n104 161.3
R2492 VN.n103 VN.n57 161.3
R2493 VN.n102 VN.n101 161.3
R2494 VN.n100 VN.n58 161.3
R2495 VN.n99 VN.n98 161.3
R2496 VN.n97 VN.n59 161.3
R2497 VN.n96 VN.n95 161.3
R2498 VN.n94 VN.n60 161.3
R2499 VN.n93 VN.n92 161.3
R2500 VN.n91 VN.n62 161.3
R2501 VN.n90 VN.n89 161.3
R2502 VN.n88 VN.n63 161.3
R2503 VN.n87 VN.n86 161.3
R2504 VN.n85 VN.n64 161.3
R2505 VN.n84 VN.n83 161.3
R2506 VN.n82 VN.n65 161.3
R2507 VN.n81 VN.n80 161.3
R2508 VN.n79 VN.n66 161.3
R2509 VN.n78 VN.n77 161.3
R2510 VN.n76 VN.n67 161.3
R2511 VN.n75 VN.n74 161.3
R2512 VN.n73 VN.n68 161.3
R2513 VN.n72 VN.n71 161.3
R2514 VN.n53 VN.n52 161.3
R2515 VN.n51 VN.n1 161.3
R2516 VN.n50 VN.n49 161.3
R2517 VN.n48 VN.n2 161.3
R2518 VN.n47 VN.n46 161.3
R2519 VN.n45 VN.n3 161.3
R2520 VN.n44 VN.n43 161.3
R2521 VN.n42 VN.n4 161.3
R2522 VN.n41 VN.n40 161.3
R2523 VN.n38 VN.n5 161.3
R2524 VN.n37 VN.n36 161.3
R2525 VN.n35 VN.n6 161.3
R2526 VN.n34 VN.n33 161.3
R2527 VN.n32 VN.n7 161.3
R2528 VN.n31 VN.n30 161.3
R2529 VN.n29 VN.n8 161.3
R2530 VN.n28 VN.n27 161.3
R2531 VN.n26 VN.n9 161.3
R2532 VN.n25 VN.n24 161.3
R2533 VN.n23 VN.n10 161.3
R2534 VN.n22 VN.n21 161.3
R2535 VN.n20 VN.n11 161.3
R2536 VN.n19 VN.n18 161.3
R2537 VN.n17 VN.n12 161.3
R2538 VN.n16 VN.n15 161.3
R2539 VN.n69 VN.t1 118.285
R2540 VN.n13 VN.t2 118.285
R2541 VN.n27 VN.t6 85.2824
R2542 VN.n14 VN.t9 85.2824
R2543 VN.n39 VN.t8 85.2824
R2544 VN.n0 VN.t4 85.2824
R2545 VN.n83 VN.t0 85.2824
R2546 VN.n70 VN.t5 85.2824
R2547 VN.n61 VN.t3 85.2824
R2548 VN.n55 VN.t7 85.2824
R2549 VN.n54 VN.n0 82.238
R2550 VN.n109 VN.n55 82.238
R2551 VN.n14 VN.n13 70.8482
R2552 VN.n70 VN.n69 70.8482
R2553 VN VN.n109 60.6117
R2554 VN.n46 VN.n2 52.1486
R2555 VN.n101 VN.n57 52.1486
R2556 VN.n21 VN.n20 44.3785
R2557 VN.n33 VN.n6 44.3785
R2558 VN.n77 VN.n76 44.3785
R2559 VN.n89 VN.n62 44.3785
R2560 VN.n21 VN.n10 36.6083
R2561 VN.n33 VN.n32 36.6083
R2562 VN.n77 VN.n66 36.6083
R2563 VN.n89 VN.n88 36.6083
R2564 VN.n46 VN.n45 28.8382
R2565 VN.n101 VN.n100 28.8382
R2566 VN.n15 VN.n12 24.4675
R2567 VN.n19 VN.n12 24.4675
R2568 VN.n20 VN.n19 24.4675
R2569 VN.n25 VN.n10 24.4675
R2570 VN.n26 VN.n25 24.4675
R2571 VN.n27 VN.n26 24.4675
R2572 VN.n27 VN.n8 24.4675
R2573 VN.n31 VN.n8 24.4675
R2574 VN.n32 VN.n31 24.4675
R2575 VN.n37 VN.n6 24.4675
R2576 VN.n38 VN.n37 24.4675
R2577 VN.n40 VN.n38 24.4675
R2578 VN.n44 VN.n4 24.4675
R2579 VN.n45 VN.n44 24.4675
R2580 VN.n50 VN.n2 24.4675
R2581 VN.n51 VN.n50 24.4675
R2582 VN.n52 VN.n51 24.4675
R2583 VN.n76 VN.n75 24.4675
R2584 VN.n75 VN.n68 24.4675
R2585 VN.n71 VN.n68 24.4675
R2586 VN.n88 VN.n87 24.4675
R2587 VN.n87 VN.n64 24.4675
R2588 VN.n83 VN.n64 24.4675
R2589 VN.n83 VN.n82 24.4675
R2590 VN.n82 VN.n81 24.4675
R2591 VN.n81 VN.n66 24.4675
R2592 VN.n100 VN.n99 24.4675
R2593 VN.n99 VN.n59 24.4675
R2594 VN.n95 VN.n94 24.4675
R2595 VN.n94 VN.n93 24.4675
R2596 VN.n93 VN.n62 24.4675
R2597 VN.n107 VN.n106 24.4675
R2598 VN.n106 VN.n105 24.4675
R2599 VN.n105 VN.n57 24.4675
R2600 VN.n39 VN.n4 20.5528
R2601 VN.n61 VN.n59 20.5528
R2602 VN.n52 VN.n0 7.82994
R2603 VN.n107 VN.n55 7.82994
R2604 VN.n15 VN.n14 3.91522
R2605 VN.n40 VN.n39 3.91522
R2606 VN.n71 VN.n70 3.91522
R2607 VN.n95 VN.n61 3.91522
R2608 VN.n72 VN.n69 3.22187
R2609 VN.n16 VN.n13 3.22187
R2610 VN.n109 VN.n108 0.354971
R2611 VN.n54 VN.n53 0.354971
R2612 VN VN.n54 0.26696
R2613 VN.n108 VN.n56 0.189894
R2614 VN.n104 VN.n56 0.189894
R2615 VN.n104 VN.n103 0.189894
R2616 VN.n103 VN.n102 0.189894
R2617 VN.n102 VN.n58 0.189894
R2618 VN.n98 VN.n58 0.189894
R2619 VN.n98 VN.n97 0.189894
R2620 VN.n97 VN.n96 0.189894
R2621 VN.n96 VN.n60 0.189894
R2622 VN.n92 VN.n60 0.189894
R2623 VN.n92 VN.n91 0.189894
R2624 VN.n91 VN.n90 0.189894
R2625 VN.n90 VN.n63 0.189894
R2626 VN.n86 VN.n63 0.189894
R2627 VN.n86 VN.n85 0.189894
R2628 VN.n85 VN.n84 0.189894
R2629 VN.n84 VN.n65 0.189894
R2630 VN.n80 VN.n65 0.189894
R2631 VN.n80 VN.n79 0.189894
R2632 VN.n79 VN.n78 0.189894
R2633 VN.n78 VN.n67 0.189894
R2634 VN.n74 VN.n67 0.189894
R2635 VN.n74 VN.n73 0.189894
R2636 VN.n73 VN.n72 0.189894
R2637 VN.n17 VN.n16 0.189894
R2638 VN.n18 VN.n17 0.189894
R2639 VN.n18 VN.n11 0.189894
R2640 VN.n22 VN.n11 0.189894
R2641 VN.n23 VN.n22 0.189894
R2642 VN.n24 VN.n23 0.189894
R2643 VN.n24 VN.n9 0.189894
R2644 VN.n28 VN.n9 0.189894
R2645 VN.n29 VN.n28 0.189894
R2646 VN.n30 VN.n29 0.189894
R2647 VN.n30 VN.n7 0.189894
R2648 VN.n34 VN.n7 0.189894
R2649 VN.n35 VN.n34 0.189894
R2650 VN.n36 VN.n35 0.189894
R2651 VN.n36 VN.n5 0.189894
R2652 VN.n41 VN.n5 0.189894
R2653 VN.n42 VN.n41 0.189894
R2654 VN.n43 VN.n42 0.189894
R2655 VN.n43 VN.n3 0.189894
R2656 VN.n47 VN.n3 0.189894
R2657 VN.n48 VN.n47 0.189894
R2658 VN.n49 VN.n48 0.189894
R2659 VN.n49 VN.n1 0.189894
R2660 VN.n53 VN.n1 0.189894
R2661 VDD2.n142 VDD2.n141 585
R2662 VDD2.n140 VDD2.n139 585
R2663 VDD2.n79 VDD2.n78 585
R2664 VDD2.n134 VDD2.n133 585
R2665 VDD2.n132 VDD2.n131 585
R2666 VDD2.n83 VDD2.n82 585
R2667 VDD2.n126 VDD2.n125 585
R2668 VDD2.n124 VDD2.n123 585
R2669 VDD2.n87 VDD2.n86 585
R2670 VDD2.n118 VDD2.n117 585
R2671 VDD2.n116 VDD2.n115 585
R2672 VDD2.n91 VDD2.n90 585
R2673 VDD2.n110 VDD2.n109 585
R2674 VDD2.n108 VDD2.n107 585
R2675 VDD2.n95 VDD2.n94 585
R2676 VDD2.n102 VDD2.n101 585
R2677 VDD2.n100 VDD2.n99 585
R2678 VDD2.n25 VDD2.n24 585
R2679 VDD2.n27 VDD2.n26 585
R2680 VDD2.n20 VDD2.n19 585
R2681 VDD2.n33 VDD2.n32 585
R2682 VDD2.n35 VDD2.n34 585
R2683 VDD2.n16 VDD2.n15 585
R2684 VDD2.n41 VDD2.n40 585
R2685 VDD2.n43 VDD2.n42 585
R2686 VDD2.n12 VDD2.n11 585
R2687 VDD2.n49 VDD2.n48 585
R2688 VDD2.n51 VDD2.n50 585
R2689 VDD2.n8 VDD2.n7 585
R2690 VDD2.n57 VDD2.n56 585
R2691 VDD2.n59 VDD2.n58 585
R2692 VDD2.n4 VDD2.n3 585
R2693 VDD2.n65 VDD2.n64 585
R2694 VDD2.n67 VDD2.n66 585
R2695 VDD2.n141 VDD2.n75 498.474
R2696 VDD2.n66 VDD2.n0 498.474
R2697 VDD2.n98 VDD2.t2 327.466
R2698 VDD2.n23 VDD2.t7 327.466
R2699 VDD2.n141 VDD2.n140 171.744
R2700 VDD2.n140 VDD2.n78 171.744
R2701 VDD2.n133 VDD2.n78 171.744
R2702 VDD2.n133 VDD2.n132 171.744
R2703 VDD2.n132 VDD2.n82 171.744
R2704 VDD2.n125 VDD2.n82 171.744
R2705 VDD2.n125 VDD2.n124 171.744
R2706 VDD2.n124 VDD2.n86 171.744
R2707 VDD2.n117 VDD2.n86 171.744
R2708 VDD2.n117 VDD2.n116 171.744
R2709 VDD2.n116 VDD2.n90 171.744
R2710 VDD2.n109 VDD2.n90 171.744
R2711 VDD2.n109 VDD2.n108 171.744
R2712 VDD2.n108 VDD2.n94 171.744
R2713 VDD2.n101 VDD2.n94 171.744
R2714 VDD2.n101 VDD2.n100 171.744
R2715 VDD2.n26 VDD2.n25 171.744
R2716 VDD2.n26 VDD2.n19 171.744
R2717 VDD2.n33 VDD2.n19 171.744
R2718 VDD2.n34 VDD2.n33 171.744
R2719 VDD2.n34 VDD2.n15 171.744
R2720 VDD2.n41 VDD2.n15 171.744
R2721 VDD2.n42 VDD2.n41 171.744
R2722 VDD2.n42 VDD2.n11 171.744
R2723 VDD2.n49 VDD2.n11 171.744
R2724 VDD2.n50 VDD2.n49 171.744
R2725 VDD2.n50 VDD2.n7 171.744
R2726 VDD2.n57 VDD2.n7 171.744
R2727 VDD2.n58 VDD2.n57 171.744
R2728 VDD2.n58 VDD2.n3 171.744
R2729 VDD2.n65 VDD2.n3 171.744
R2730 VDD2.n66 VDD2.n65 171.744
R2731 VDD2.n100 VDD2.t2 85.8723
R2732 VDD2.n25 VDD2.t7 85.8723
R2733 VDD2.n74 VDD2.n73 75.9066
R2734 VDD2 VDD2.n149 75.9037
R2735 VDD2.n148 VDD2.n147 73.3241
R2736 VDD2.n72 VDD2.n71 73.324
R2737 VDD2.n72 VDD2.n70 53.739
R2738 VDD2.n146 VDD2.n74 51.8618
R2739 VDD2.n146 VDD2.n145 50.2217
R2740 VDD2.n99 VDD2.n98 16.3895
R2741 VDD2.n24 VDD2.n23 16.3895
R2742 VDD2.n143 VDD2.n142 12.8005
R2743 VDD2.n102 VDD2.n97 12.8005
R2744 VDD2.n27 VDD2.n22 12.8005
R2745 VDD2.n68 VDD2.n67 12.8005
R2746 VDD2.n139 VDD2.n77 12.0247
R2747 VDD2.n103 VDD2.n95 12.0247
R2748 VDD2.n28 VDD2.n20 12.0247
R2749 VDD2.n64 VDD2.n2 12.0247
R2750 VDD2.n138 VDD2.n79 11.249
R2751 VDD2.n107 VDD2.n106 11.249
R2752 VDD2.n32 VDD2.n31 11.249
R2753 VDD2.n63 VDD2.n4 11.249
R2754 VDD2.n135 VDD2.n134 10.4732
R2755 VDD2.n110 VDD2.n93 10.4732
R2756 VDD2.n35 VDD2.n18 10.4732
R2757 VDD2.n60 VDD2.n59 10.4732
R2758 VDD2.n131 VDD2.n81 9.69747
R2759 VDD2.n111 VDD2.n91 9.69747
R2760 VDD2.n36 VDD2.n16 9.69747
R2761 VDD2.n56 VDD2.n6 9.69747
R2762 VDD2.n145 VDD2.n144 9.45567
R2763 VDD2.n70 VDD2.n69 9.45567
R2764 VDD2.n85 VDD2.n84 9.3005
R2765 VDD2.n128 VDD2.n127 9.3005
R2766 VDD2.n130 VDD2.n129 9.3005
R2767 VDD2.n81 VDD2.n80 9.3005
R2768 VDD2.n136 VDD2.n135 9.3005
R2769 VDD2.n138 VDD2.n137 9.3005
R2770 VDD2.n77 VDD2.n76 9.3005
R2771 VDD2.n144 VDD2.n143 9.3005
R2772 VDD2.n122 VDD2.n121 9.3005
R2773 VDD2.n120 VDD2.n119 9.3005
R2774 VDD2.n89 VDD2.n88 9.3005
R2775 VDD2.n114 VDD2.n113 9.3005
R2776 VDD2.n112 VDD2.n111 9.3005
R2777 VDD2.n93 VDD2.n92 9.3005
R2778 VDD2.n106 VDD2.n105 9.3005
R2779 VDD2.n104 VDD2.n103 9.3005
R2780 VDD2.n97 VDD2.n96 9.3005
R2781 VDD2.n45 VDD2.n44 9.3005
R2782 VDD2.n14 VDD2.n13 9.3005
R2783 VDD2.n39 VDD2.n38 9.3005
R2784 VDD2.n37 VDD2.n36 9.3005
R2785 VDD2.n18 VDD2.n17 9.3005
R2786 VDD2.n31 VDD2.n30 9.3005
R2787 VDD2.n29 VDD2.n28 9.3005
R2788 VDD2.n22 VDD2.n21 9.3005
R2789 VDD2.n47 VDD2.n46 9.3005
R2790 VDD2.n10 VDD2.n9 9.3005
R2791 VDD2.n53 VDD2.n52 9.3005
R2792 VDD2.n55 VDD2.n54 9.3005
R2793 VDD2.n6 VDD2.n5 9.3005
R2794 VDD2.n61 VDD2.n60 9.3005
R2795 VDD2.n63 VDD2.n62 9.3005
R2796 VDD2.n2 VDD2.n1 9.3005
R2797 VDD2.n69 VDD2.n68 9.3005
R2798 VDD2.n130 VDD2.n83 8.92171
R2799 VDD2.n115 VDD2.n114 8.92171
R2800 VDD2.n40 VDD2.n39 8.92171
R2801 VDD2.n55 VDD2.n8 8.92171
R2802 VDD2.n127 VDD2.n126 8.14595
R2803 VDD2.n118 VDD2.n89 8.14595
R2804 VDD2.n43 VDD2.n14 8.14595
R2805 VDD2.n52 VDD2.n51 8.14595
R2806 VDD2.n145 VDD2.n75 7.75445
R2807 VDD2.n70 VDD2.n0 7.75445
R2808 VDD2.n123 VDD2.n85 7.3702
R2809 VDD2.n119 VDD2.n87 7.3702
R2810 VDD2.n44 VDD2.n12 7.3702
R2811 VDD2.n48 VDD2.n10 7.3702
R2812 VDD2.n123 VDD2.n122 6.59444
R2813 VDD2.n122 VDD2.n87 6.59444
R2814 VDD2.n47 VDD2.n12 6.59444
R2815 VDD2.n48 VDD2.n47 6.59444
R2816 VDD2.n143 VDD2.n75 6.08283
R2817 VDD2.n68 VDD2.n0 6.08283
R2818 VDD2.n126 VDD2.n85 5.81868
R2819 VDD2.n119 VDD2.n118 5.81868
R2820 VDD2.n44 VDD2.n43 5.81868
R2821 VDD2.n51 VDD2.n10 5.81868
R2822 VDD2.n127 VDD2.n83 5.04292
R2823 VDD2.n115 VDD2.n89 5.04292
R2824 VDD2.n40 VDD2.n14 5.04292
R2825 VDD2.n52 VDD2.n8 5.04292
R2826 VDD2.n131 VDD2.n130 4.26717
R2827 VDD2.n114 VDD2.n91 4.26717
R2828 VDD2.n39 VDD2.n16 4.26717
R2829 VDD2.n56 VDD2.n55 4.26717
R2830 VDD2.n98 VDD2.n96 3.70982
R2831 VDD2.n23 VDD2.n21 3.70982
R2832 VDD2.n148 VDD2.n146 3.51774
R2833 VDD2.n134 VDD2.n81 3.49141
R2834 VDD2.n111 VDD2.n110 3.49141
R2835 VDD2.n36 VDD2.n35 3.49141
R2836 VDD2.n59 VDD2.n6 3.49141
R2837 VDD2.n135 VDD2.n79 2.71565
R2838 VDD2.n107 VDD2.n93 2.71565
R2839 VDD2.n32 VDD2.n18 2.71565
R2840 VDD2.n60 VDD2.n4 2.71565
R2841 VDD2.n149 VDD2.t4 2.45001
R2842 VDD2.n149 VDD2.t8 2.45001
R2843 VDD2.n147 VDD2.t6 2.45001
R2844 VDD2.n147 VDD2.t9 2.45001
R2845 VDD2.n73 VDD2.t1 2.45001
R2846 VDD2.n73 VDD2.t5 2.45001
R2847 VDD2.n71 VDD2.t0 2.45001
R2848 VDD2.n71 VDD2.t3 2.45001
R2849 VDD2.n139 VDD2.n138 1.93989
R2850 VDD2.n106 VDD2.n95 1.93989
R2851 VDD2.n31 VDD2.n20 1.93989
R2852 VDD2.n64 VDD2.n63 1.93989
R2853 VDD2.n142 VDD2.n77 1.16414
R2854 VDD2.n103 VDD2.n102 1.16414
R2855 VDD2.n28 VDD2.n27 1.16414
R2856 VDD2.n67 VDD2.n2 1.16414
R2857 VDD2 VDD2.n148 0.938
R2858 VDD2.n74 VDD2.n72 0.824464
R2859 VDD2.n99 VDD2.n97 0.388379
R2860 VDD2.n24 VDD2.n22 0.388379
R2861 VDD2.n144 VDD2.n76 0.155672
R2862 VDD2.n137 VDD2.n76 0.155672
R2863 VDD2.n137 VDD2.n136 0.155672
R2864 VDD2.n136 VDD2.n80 0.155672
R2865 VDD2.n129 VDD2.n80 0.155672
R2866 VDD2.n129 VDD2.n128 0.155672
R2867 VDD2.n128 VDD2.n84 0.155672
R2868 VDD2.n121 VDD2.n84 0.155672
R2869 VDD2.n121 VDD2.n120 0.155672
R2870 VDD2.n120 VDD2.n88 0.155672
R2871 VDD2.n113 VDD2.n88 0.155672
R2872 VDD2.n113 VDD2.n112 0.155672
R2873 VDD2.n112 VDD2.n92 0.155672
R2874 VDD2.n105 VDD2.n92 0.155672
R2875 VDD2.n105 VDD2.n104 0.155672
R2876 VDD2.n104 VDD2.n96 0.155672
R2877 VDD2.n29 VDD2.n21 0.155672
R2878 VDD2.n30 VDD2.n29 0.155672
R2879 VDD2.n30 VDD2.n17 0.155672
R2880 VDD2.n37 VDD2.n17 0.155672
R2881 VDD2.n38 VDD2.n37 0.155672
R2882 VDD2.n38 VDD2.n13 0.155672
R2883 VDD2.n45 VDD2.n13 0.155672
R2884 VDD2.n46 VDD2.n45 0.155672
R2885 VDD2.n46 VDD2.n9 0.155672
R2886 VDD2.n53 VDD2.n9 0.155672
R2887 VDD2.n54 VDD2.n53 0.155672
R2888 VDD2.n54 VDD2.n5 0.155672
R2889 VDD2.n61 VDD2.n5 0.155672
R2890 VDD2.n62 VDD2.n61 0.155672
R2891 VDD2.n62 VDD2.n1 0.155672
R2892 VDD2.n69 VDD2.n1 0.155672
C0 VP VTAIL 13.587f
C1 VDD1 B 3.02934f
C2 VP B 2.88737f
C3 VP VDD1 13.0686f
C4 VN VTAIL 13.572299f
C5 VDD2 w_n5866_n3622# 3.51064f
C6 VN B 1.59082f
C7 VN VDD1 0.15585f
C8 VP VN 10.3276f
C9 VTAIL w_n5866_n3622# 3.54202f
C10 w_n5866_n3622# B 12.8361f
C11 VDD1 w_n5866_n3622# 3.30732f
C12 VP w_n5866_n3622# 13.6847f
C13 VDD2 VTAIL 11.528799f
C14 VDD2 B 3.19204f
C15 VN w_n5866_n3622# 12.9175f
C16 VDD2 VDD1 2.92277f
C17 VP VDD2 0.729821f
C18 VN VDD2 12.4983f
C19 VTAIL B 4.46731f
C20 VTAIL VDD1 11.469501f
C21 VDD2 VSUBS 2.60121f
C22 VDD1 VSUBS 2.468257f
C23 VTAIL VSUBS 1.619824f
C24 VN VSUBS 9.64729f
C25 VP VSUBS 5.748349f
C26 B VSUBS 6.89876f
C27 w_n5866_n3622# VSUBS 0.261084p
C28 VDD2.n0 VSUBS 0.031648f
C29 VDD2.n1 VSUBS 0.030584f
C30 VDD2.n2 VSUBS 0.016434f
C31 VDD2.n3 VSUBS 0.038844f
C32 VDD2.n4 VSUBS 0.017401f
C33 VDD2.n5 VSUBS 0.030584f
C34 VDD2.n6 VSUBS 0.016434f
C35 VDD2.n7 VSUBS 0.038844f
C36 VDD2.n8 VSUBS 0.017401f
C37 VDD2.n9 VSUBS 0.030584f
C38 VDD2.n10 VSUBS 0.016434f
C39 VDD2.n11 VSUBS 0.038844f
C40 VDD2.n12 VSUBS 0.017401f
C41 VDD2.n13 VSUBS 0.030584f
C42 VDD2.n14 VSUBS 0.016434f
C43 VDD2.n15 VSUBS 0.038844f
C44 VDD2.n16 VSUBS 0.017401f
C45 VDD2.n17 VSUBS 0.030584f
C46 VDD2.n18 VSUBS 0.016434f
C47 VDD2.n19 VSUBS 0.038844f
C48 VDD2.n20 VSUBS 0.017401f
C49 VDD2.n21 VSUBS 1.71262f
C50 VDD2.n22 VSUBS 0.016434f
C51 VDD2.t7 VSUBS 0.083028f
C52 VDD2.n23 VSUBS 0.199982f
C53 VDD2.n24 VSUBS 0.024711f
C54 VDD2.n25 VSUBS 0.029133f
C55 VDD2.n26 VSUBS 0.038844f
C56 VDD2.n27 VSUBS 0.017401f
C57 VDD2.n28 VSUBS 0.016434f
C58 VDD2.n29 VSUBS 0.030584f
C59 VDD2.n30 VSUBS 0.030584f
C60 VDD2.n31 VSUBS 0.016434f
C61 VDD2.n32 VSUBS 0.017401f
C62 VDD2.n33 VSUBS 0.038844f
C63 VDD2.n34 VSUBS 0.038844f
C64 VDD2.n35 VSUBS 0.017401f
C65 VDD2.n36 VSUBS 0.016434f
C66 VDD2.n37 VSUBS 0.030584f
C67 VDD2.n38 VSUBS 0.030584f
C68 VDD2.n39 VSUBS 0.016434f
C69 VDD2.n40 VSUBS 0.017401f
C70 VDD2.n41 VSUBS 0.038844f
C71 VDD2.n42 VSUBS 0.038844f
C72 VDD2.n43 VSUBS 0.017401f
C73 VDD2.n44 VSUBS 0.016434f
C74 VDD2.n45 VSUBS 0.030584f
C75 VDD2.n46 VSUBS 0.030584f
C76 VDD2.n47 VSUBS 0.016434f
C77 VDD2.n48 VSUBS 0.017401f
C78 VDD2.n49 VSUBS 0.038844f
C79 VDD2.n50 VSUBS 0.038844f
C80 VDD2.n51 VSUBS 0.017401f
C81 VDD2.n52 VSUBS 0.016434f
C82 VDD2.n53 VSUBS 0.030584f
C83 VDD2.n54 VSUBS 0.030584f
C84 VDD2.n55 VSUBS 0.016434f
C85 VDD2.n56 VSUBS 0.017401f
C86 VDD2.n57 VSUBS 0.038844f
C87 VDD2.n58 VSUBS 0.038844f
C88 VDD2.n59 VSUBS 0.017401f
C89 VDD2.n60 VSUBS 0.016434f
C90 VDD2.n61 VSUBS 0.030584f
C91 VDD2.n62 VSUBS 0.030584f
C92 VDD2.n63 VSUBS 0.016434f
C93 VDD2.n64 VSUBS 0.017401f
C94 VDD2.n65 VSUBS 0.038844f
C95 VDD2.n66 VSUBS 0.094119f
C96 VDD2.n67 VSUBS 0.017401f
C97 VDD2.n68 VSUBS 0.032273f
C98 VDD2.n69 VSUBS 0.073617f
C99 VDD2.n70 VSUBS 0.118567f
C100 VDD2.t0 VSUBS 0.320709f
C101 VDD2.t3 VSUBS 0.320709f
C102 VDD2.n71 VSUBS 2.5621f
C103 VDD2.n72 VSUBS 1.37651f
C104 VDD2.t1 VSUBS 0.320709f
C105 VDD2.t5 VSUBS 0.320709f
C106 VDD2.n73 VSUBS 2.60229f
C107 VDD2.n74 VSUBS 4.69262f
C108 VDD2.n75 VSUBS 0.031648f
C109 VDD2.n76 VSUBS 0.030584f
C110 VDD2.n77 VSUBS 0.016434f
C111 VDD2.n78 VSUBS 0.038844f
C112 VDD2.n79 VSUBS 0.017401f
C113 VDD2.n80 VSUBS 0.030584f
C114 VDD2.n81 VSUBS 0.016434f
C115 VDD2.n82 VSUBS 0.038844f
C116 VDD2.n83 VSUBS 0.017401f
C117 VDD2.n84 VSUBS 0.030584f
C118 VDD2.n85 VSUBS 0.016434f
C119 VDD2.n86 VSUBS 0.038844f
C120 VDD2.n87 VSUBS 0.017401f
C121 VDD2.n88 VSUBS 0.030584f
C122 VDD2.n89 VSUBS 0.016434f
C123 VDD2.n90 VSUBS 0.038844f
C124 VDD2.n91 VSUBS 0.017401f
C125 VDD2.n92 VSUBS 0.030584f
C126 VDD2.n93 VSUBS 0.016434f
C127 VDD2.n94 VSUBS 0.038844f
C128 VDD2.n95 VSUBS 0.017401f
C129 VDD2.n96 VSUBS 1.71262f
C130 VDD2.n97 VSUBS 0.016434f
C131 VDD2.t2 VSUBS 0.083028f
C132 VDD2.n98 VSUBS 0.199982f
C133 VDD2.n99 VSUBS 0.024711f
C134 VDD2.n100 VSUBS 0.029133f
C135 VDD2.n101 VSUBS 0.038844f
C136 VDD2.n102 VSUBS 0.017401f
C137 VDD2.n103 VSUBS 0.016434f
C138 VDD2.n104 VSUBS 0.030584f
C139 VDD2.n105 VSUBS 0.030584f
C140 VDD2.n106 VSUBS 0.016434f
C141 VDD2.n107 VSUBS 0.017401f
C142 VDD2.n108 VSUBS 0.038844f
C143 VDD2.n109 VSUBS 0.038844f
C144 VDD2.n110 VSUBS 0.017401f
C145 VDD2.n111 VSUBS 0.016434f
C146 VDD2.n112 VSUBS 0.030584f
C147 VDD2.n113 VSUBS 0.030584f
C148 VDD2.n114 VSUBS 0.016434f
C149 VDD2.n115 VSUBS 0.017401f
C150 VDD2.n116 VSUBS 0.038844f
C151 VDD2.n117 VSUBS 0.038844f
C152 VDD2.n118 VSUBS 0.017401f
C153 VDD2.n119 VSUBS 0.016434f
C154 VDD2.n120 VSUBS 0.030584f
C155 VDD2.n121 VSUBS 0.030584f
C156 VDD2.n122 VSUBS 0.016434f
C157 VDD2.n123 VSUBS 0.017401f
C158 VDD2.n124 VSUBS 0.038844f
C159 VDD2.n125 VSUBS 0.038844f
C160 VDD2.n126 VSUBS 0.017401f
C161 VDD2.n127 VSUBS 0.016434f
C162 VDD2.n128 VSUBS 0.030584f
C163 VDD2.n129 VSUBS 0.030584f
C164 VDD2.n130 VSUBS 0.016434f
C165 VDD2.n131 VSUBS 0.017401f
C166 VDD2.n132 VSUBS 0.038844f
C167 VDD2.n133 VSUBS 0.038844f
C168 VDD2.n134 VSUBS 0.017401f
C169 VDD2.n135 VSUBS 0.016434f
C170 VDD2.n136 VSUBS 0.030584f
C171 VDD2.n137 VSUBS 0.030584f
C172 VDD2.n138 VSUBS 0.016434f
C173 VDD2.n139 VSUBS 0.017401f
C174 VDD2.n140 VSUBS 0.038844f
C175 VDD2.n141 VSUBS 0.094119f
C176 VDD2.n142 VSUBS 0.017401f
C177 VDD2.n143 VSUBS 0.032273f
C178 VDD2.n144 VSUBS 0.073617f
C179 VDD2.n145 VSUBS 0.091917f
C180 VDD2.n146 VSUBS 4.2049f
C181 VDD2.t6 VSUBS 0.320709f
C182 VDD2.t9 VSUBS 0.320709f
C183 VDD2.n147 VSUBS 2.56212f
C184 VDD2.n148 VSUBS 1.0063f
C185 VDD2.t4 VSUBS 0.320709f
C186 VDD2.t8 VSUBS 0.320709f
C187 VDD2.n149 VSUBS 2.60223f
C188 VN.t4 VSUBS 3.06378f
C189 VN.n0 VSUBS 1.15804f
C190 VN.n1 VSUBS 0.022535f
C191 VN.n2 VSUBS 0.040457f
C192 VN.n3 VSUBS 0.022535f
C193 VN.n4 VSUBS 0.038682f
C194 VN.n5 VSUBS 0.022535f
C195 VN.n6 VSUBS 0.043673f
C196 VN.n7 VSUBS 0.022535f
C197 VN.n8 VSUBS 0.042f
C198 VN.n9 VSUBS 0.022535f
C199 VN.t6 VSUBS 3.06378f
C200 VN.n10 VSUBS 0.045437f
C201 VN.n11 VSUBS 0.022535f
C202 VN.n12 VSUBS 0.042f
C203 VN.t2 VSUBS 3.41062f
C204 VN.n13 VSUBS 1.08355f
C205 VN.t9 VSUBS 3.06378f
C206 VN.n14 VSUBS 1.14178f
C207 VN.n15 VSUBS 0.024582f
C208 VN.n16 VSUBS 0.286173f
C209 VN.n17 VSUBS 0.022535f
C210 VN.n18 VSUBS 0.022535f
C211 VN.n19 VSUBS 0.042f
C212 VN.n20 VSUBS 0.043673f
C213 VN.n21 VSUBS 0.018685f
C214 VN.n22 VSUBS 0.022535f
C215 VN.n23 VSUBS 0.022535f
C216 VN.n24 VSUBS 0.022535f
C217 VN.n25 VSUBS 0.042f
C218 VN.n26 VSUBS 0.042f
C219 VN.n27 VSUBS 1.08958f
C220 VN.n28 VSUBS 0.022535f
C221 VN.n29 VSUBS 0.022535f
C222 VN.n30 VSUBS 0.022535f
C223 VN.n31 VSUBS 0.042f
C224 VN.n32 VSUBS 0.045437f
C225 VN.n33 VSUBS 0.018685f
C226 VN.n34 VSUBS 0.022535f
C227 VN.n35 VSUBS 0.022535f
C228 VN.n36 VSUBS 0.022535f
C229 VN.n37 VSUBS 0.042f
C230 VN.n38 VSUBS 0.042f
C231 VN.t8 VSUBS 3.06378f
C232 VN.n39 VSUBS 1.06831f
C233 VN.n40 VSUBS 0.024582f
C234 VN.n41 VSUBS 0.022535f
C235 VN.n42 VSUBS 0.022535f
C236 VN.n43 VSUBS 0.022535f
C237 VN.n44 VSUBS 0.042f
C238 VN.n45 VSUBS 0.044576f
C239 VN.n46 VSUBS 0.022762f
C240 VN.n47 VSUBS 0.022535f
C241 VN.n48 VSUBS 0.022535f
C242 VN.n49 VSUBS 0.022535f
C243 VN.n50 VSUBS 0.042f
C244 VN.n51 VSUBS 0.042f
C245 VN.n52 VSUBS 0.0279f
C246 VN.n53 VSUBS 0.036371f
C247 VN.n54 VSUBS 0.065013f
C248 VN.t7 VSUBS 3.06378f
C249 VN.n55 VSUBS 1.15804f
C250 VN.n56 VSUBS 0.022535f
C251 VN.n57 VSUBS 0.040457f
C252 VN.n58 VSUBS 0.022535f
C253 VN.n59 VSUBS 0.038682f
C254 VN.n60 VSUBS 0.022535f
C255 VN.t3 VSUBS 3.06378f
C256 VN.n61 VSUBS 1.06831f
C257 VN.n62 VSUBS 0.043673f
C258 VN.n63 VSUBS 0.022535f
C259 VN.n64 VSUBS 0.042f
C260 VN.n65 VSUBS 0.022535f
C261 VN.t0 VSUBS 3.06378f
C262 VN.n66 VSUBS 0.045437f
C263 VN.n67 VSUBS 0.022535f
C264 VN.n68 VSUBS 0.042f
C265 VN.t1 VSUBS 3.41062f
C266 VN.n69 VSUBS 1.08355f
C267 VN.t5 VSUBS 3.06378f
C268 VN.n70 VSUBS 1.14178f
C269 VN.n71 VSUBS 0.024582f
C270 VN.n72 VSUBS 0.286173f
C271 VN.n73 VSUBS 0.022535f
C272 VN.n74 VSUBS 0.022535f
C273 VN.n75 VSUBS 0.042f
C274 VN.n76 VSUBS 0.043673f
C275 VN.n77 VSUBS 0.018685f
C276 VN.n78 VSUBS 0.022535f
C277 VN.n79 VSUBS 0.022535f
C278 VN.n80 VSUBS 0.022535f
C279 VN.n81 VSUBS 0.042f
C280 VN.n82 VSUBS 0.042f
C281 VN.n83 VSUBS 1.08958f
C282 VN.n84 VSUBS 0.022535f
C283 VN.n85 VSUBS 0.022535f
C284 VN.n86 VSUBS 0.022535f
C285 VN.n87 VSUBS 0.042f
C286 VN.n88 VSUBS 0.045437f
C287 VN.n89 VSUBS 0.018685f
C288 VN.n90 VSUBS 0.022535f
C289 VN.n91 VSUBS 0.022535f
C290 VN.n92 VSUBS 0.022535f
C291 VN.n93 VSUBS 0.042f
C292 VN.n94 VSUBS 0.042f
C293 VN.n95 VSUBS 0.024582f
C294 VN.n96 VSUBS 0.022535f
C295 VN.n97 VSUBS 0.022535f
C296 VN.n98 VSUBS 0.022535f
C297 VN.n99 VSUBS 0.042f
C298 VN.n100 VSUBS 0.044576f
C299 VN.n101 VSUBS 0.022762f
C300 VN.n102 VSUBS 0.022535f
C301 VN.n103 VSUBS 0.022535f
C302 VN.n104 VSUBS 0.022535f
C303 VN.n105 VSUBS 0.042f
C304 VN.n106 VSUBS 0.042f
C305 VN.n107 VSUBS 0.0279f
C306 VN.n108 VSUBS 0.036371f
C307 VN.n109 VSUBS 1.68712f
C308 B.n0 VSUBS 0.005372f
C309 B.n1 VSUBS 0.005372f
C310 B.n2 VSUBS 0.008494f
C311 B.n3 VSUBS 0.008494f
C312 B.n4 VSUBS 0.008494f
C313 B.n5 VSUBS 0.008494f
C314 B.n6 VSUBS 0.008494f
C315 B.n7 VSUBS 0.008494f
C316 B.n8 VSUBS 0.008494f
C317 B.n9 VSUBS 0.008494f
C318 B.n10 VSUBS 0.008494f
C319 B.n11 VSUBS 0.008494f
C320 B.n12 VSUBS 0.008494f
C321 B.n13 VSUBS 0.008494f
C322 B.n14 VSUBS 0.008494f
C323 B.n15 VSUBS 0.008494f
C324 B.n16 VSUBS 0.008494f
C325 B.n17 VSUBS 0.008494f
C326 B.n18 VSUBS 0.008494f
C327 B.n19 VSUBS 0.008494f
C328 B.n20 VSUBS 0.008494f
C329 B.n21 VSUBS 0.008494f
C330 B.n22 VSUBS 0.008494f
C331 B.n23 VSUBS 0.008494f
C332 B.n24 VSUBS 0.008494f
C333 B.n25 VSUBS 0.008494f
C334 B.n26 VSUBS 0.008494f
C335 B.n27 VSUBS 0.008494f
C336 B.n28 VSUBS 0.008494f
C337 B.n29 VSUBS 0.008494f
C338 B.n30 VSUBS 0.008494f
C339 B.n31 VSUBS 0.008494f
C340 B.n32 VSUBS 0.008494f
C341 B.n33 VSUBS 0.008494f
C342 B.n34 VSUBS 0.008494f
C343 B.n35 VSUBS 0.008494f
C344 B.n36 VSUBS 0.008494f
C345 B.n37 VSUBS 0.008494f
C346 B.n38 VSUBS 0.008494f
C347 B.n39 VSUBS 0.008494f
C348 B.n40 VSUBS 0.008494f
C349 B.n41 VSUBS 0.008494f
C350 B.n42 VSUBS 0.021283f
C351 B.n43 VSUBS 0.008494f
C352 B.n44 VSUBS 0.008494f
C353 B.n45 VSUBS 0.008494f
C354 B.n46 VSUBS 0.008494f
C355 B.n47 VSUBS 0.008494f
C356 B.n48 VSUBS 0.008494f
C357 B.n49 VSUBS 0.008494f
C358 B.n50 VSUBS 0.008494f
C359 B.n51 VSUBS 0.008494f
C360 B.n52 VSUBS 0.008494f
C361 B.n53 VSUBS 0.008494f
C362 B.n54 VSUBS 0.008494f
C363 B.n55 VSUBS 0.008494f
C364 B.n56 VSUBS 0.008494f
C365 B.n57 VSUBS 0.008494f
C366 B.n58 VSUBS 0.008494f
C367 B.n59 VSUBS 0.008494f
C368 B.n60 VSUBS 0.008494f
C369 B.n61 VSUBS 0.008494f
C370 B.n62 VSUBS 0.008494f
C371 B.n63 VSUBS 0.008494f
C372 B.n64 VSUBS 0.007995f
C373 B.n65 VSUBS 0.008494f
C374 B.t5 VSUBS 0.2905f
C375 B.t4 VSUBS 0.343631f
C376 B.t3 VSUBS 2.79896f
C377 B.n66 VSUBS 0.548462f
C378 B.n67 VSUBS 0.33268f
C379 B.n68 VSUBS 0.019681f
C380 B.n69 VSUBS 0.008494f
C381 B.n70 VSUBS 0.008494f
C382 B.n71 VSUBS 0.008494f
C383 B.n72 VSUBS 0.008494f
C384 B.t2 VSUBS 0.290504f
C385 B.t1 VSUBS 0.343635f
C386 B.t0 VSUBS 2.79896f
C387 B.n73 VSUBS 0.548459f
C388 B.n74 VSUBS 0.332676f
C389 B.n75 VSUBS 0.008494f
C390 B.n76 VSUBS 0.008494f
C391 B.n77 VSUBS 0.008494f
C392 B.n78 VSUBS 0.008494f
C393 B.n79 VSUBS 0.008494f
C394 B.n80 VSUBS 0.008494f
C395 B.n81 VSUBS 0.008494f
C396 B.n82 VSUBS 0.008494f
C397 B.n83 VSUBS 0.008494f
C398 B.n84 VSUBS 0.008494f
C399 B.n85 VSUBS 0.008494f
C400 B.n86 VSUBS 0.008494f
C401 B.n87 VSUBS 0.008494f
C402 B.n88 VSUBS 0.008494f
C403 B.n89 VSUBS 0.008494f
C404 B.n90 VSUBS 0.008494f
C405 B.n91 VSUBS 0.008494f
C406 B.n92 VSUBS 0.008494f
C407 B.n93 VSUBS 0.008494f
C408 B.n94 VSUBS 0.008494f
C409 B.n95 VSUBS 0.008494f
C410 B.n96 VSUBS 0.008494f
C411 B.n97 VSUBS 0.021374f
C412 B.n98 VSUBS 0.008494f
C413 B.n99 VSUBS 0.008494f
C414 B.n100 VSUBS 0.008494f
C415 B.n101 VSUBS 0.008494f
C416 B.n102 VSUBS 0.008494f
C417 B.n103 VSUBS 0.008494f
C418 B.n104 VSUBS 0.008494f
C419 B.n105 VSUBS 0.008494f
C420 B.n106 VSUBS 0.008494f
C421 B.n107 VSUBS 0.008494f
C422 B.n108 VSUBS 0.008494f
C423 B.n109 VSUBS 0.008494f
C424 B.n110 VSUBS 0.008494f
C425 B.n111 VSUBS 0.008494f
C426 B.n112 VSUBS 0.008494f
C427 B.n113 VSUBS 0.008494f
C428 B.n114 VSUBS 0.008494f
C429 B.n115 VSUBS 0.008494f
C430 B.n116 VSUBS 0.008494f
C431 B.n117 VSUBS 0.008494f
C432 B.n118 VSUBS 0.008494f
C433 B.n119 VSUBS 0.008494f
C434 B.n120 VSUBS 0.008494f
C435 B.n121 VSUBS 0.008494f
C436 B.n122 VSUBS 0.008494f
C437 B.n123 VSUBS 0.008494f
C438 B.n124 VSUBS 0.008494f
C439 B.n125 VSUBS 0.008494f
C440 B.n126 VSUBS 0.008494f
C441 B.n127 VSUBS 0.008494f
C442 B.n128 VSUBS 0.008494f
C443 B.n129 VSUBS 0.008494f
C444 B.n130 VSUBS 0.008494f
C445 B.n131 VSUBS 0.008494f
C446 B.n132 VSUBS 0.008494f
C447 B.n133 VSUBS 0.008494f
C448 B.n134 VSUBS 0.008494f
C449 B.n135 VSUBS 0.008494f
C450 B.n136 VSUBS 0.008494f
C451 B.n137 VSUBS 0.008494f
C452 B.n138 VSUBS 0.008494f
C453 B.n139 VSUBS 0.008494f
C454 B.n140 VSUBS 0.008494f
C455 B.n141 VSUBS 0.008494f
C456 B.n142 VSUBS 0.008494f
C457 B.n143 VSUBS 0.008494f
C458 B.n144 VSUBS 0.008494f
C459 B.n145 VSUBS 0.008494f
C460 B.n146 VSUBS 0.008494f
C461 B.n147 VSUBS 0.008494f
C462 B.n148 VSUBS 0.008494f
C463 B.n149 VSUBS 0.008494f
C464 B.n150 VSUBS 0.008494f
C465 B.n151 VSUBS 0.008494f
C466 B.n152 VSUBS 0.008494f
C467 B.n153 VSUBS 0.008494f
C468 B.n154 VSUBS 0.008494f
C469 B.n155 VSUBS 0.008494f
C470 B.n156 VSUBS 0.008494f
C471 B.n157 VSUBS 0.008494f
C472 B.n158 VSUBS 0.008494f
C473 B.n159 VSUBS 0.008494f
C474 B.n160 VSUBS 0.008494f
C475 B.n161 VSUBS 0.008494f
C476 B.n162 VSUBS 0.008494f
C477 B.n163 VSUBS 0.008494f
C478 B.n164 VSUBS 0.008494f
C479 B.n165 VSUBS 0.008494f
C480 B.n166 VSUBS 0.008494f
C481 B.n167 VSUBS 0.008494f
C482 B.n168 VSUBS 0.008494f
C483 B.n169 VSUBS 0.008494f
C484 B.n170 VSUBS 0.008494f
C485 B.n171 VSUBS 0.008494f
C486 B.n172 VSUBS 0.008494f
C487 B.n173 VSUBS 0.008494f
C488 B.n174 VSUBS 0.008494f
C489 B.n175 VSUBS 0.008494f
C490 B.n176 VSUBS 0.008494f
C491 B.n177 VSUBS 0.02044f
C492 B.n178 VSUBS 0.008494f
C493 B.n179 VSUBS 0.008494f
C494 B.n180 VSUBS 0.008494f
C495 B.n181 VSUBS 0.008494f
C496 B.n182 VSUBS 0.008494f
C497 B.n183 VSUBS 0.008494f
C498 B.n184 VSUBS 0.008494f
C499 B.n185 VSUBS 0.008494f
C500 B.n186 VSUBS 0.008494f
C501 B.n187 VSUBS 0.008494f
C502 B.n188 VSUBS 0.008494f
C503 B.n189 VSUBS 0.008494f
C504 B.n190 VSUBS 0.008494f
C505 B.n191 VSUBS 0.008494f
C506 B.n192 VSUBS 0.008494f
C507 B.n193 VSUBS 0.008494f
C508 B.n194 VSUBS 0.008494f
C509 B.n195 VSUBS 0.008494f
C510 B.n196 VSUBS 0.008494f
C511 B.n197 VSUBS 0.008494f
C512 B.n198 VSUBS 0.008494f
C513 B.n199 VSUBS 0.008494f
C514 B.n200 VSUBS 0.008494f
C515 B.t10 VSUBS 0.290504f
C516 B.t11 VSUBS 0.343635f
C517 B.t9 VSUBS 2.79896f
C518 B.n201 VSUBS 0.548459f
C519 B.n202 VSUBS 0.332676f
C520 B.n203 VSUBS 0.008494f
C521 B.n204 VSUBS 0.008494f
C522 B.n205 VSUBS 0.008494f
C523 B.n206 VSUBS 0.008494f
C524 B.t7 VSUBS 0.2905f
C525 B.t8 VSUBS 0.343631f
C526 B.t6 VSUBS 2.79896f
C527 B.n207 VSUBS 0.548462f
C528 B.n208 VSUBS 0.33268f
C529 B.n209 VSUBS 0.019681f
C530 B.n210 VSUBS 0.008494f
C531 B.n211 VSUBS 0.008494f
C532 B.n212 VSUBS 0.008494f
C533 B.n213 VSUBS 0.008494f
C534 B.n214 VSUBS 0.008494f
C535 B.n215 VSUBS 0.008494f
C536 B.n216 VSUBS 0.008494f
C537 B.n217 VSUBS 0.008494f
C538 B.n218 VSUBS 0.008494f
C539 B.n219 VSUBS 0.008494f
C540 B.n220 VSUBS 0.008494f
C541 B.n221 VSUBS 0.008494f
C542 B.n222 VSUBS 0.008494f
C543 B.n223 VSUBS 0.008494f
C544 B.n224 VSUBS 0.008494f
C545 B.n225 VSUBS 0.008494f
C546 B.n226 VSUBS 0.008494f
C547 B.n227 VSUBS 0.008494f
C548 B.n228 VSUBS 0.008494f
C549 B.n229 VSUBS 0.008494f
C550 B.n230 VSUBS 0.008494f
C551 B.n231 VSUBS 0.008494f
C552 B.n232 VSUBS 0.02044f
C553 B.n233 VSUBS 0.008494f
C554 B.n234 VSUBS 0.008494f
C555 B.n235 VSUBS 0.008494f
C556 B.n236 VSUBS 0.008494f
C557 B.n237 VSUBS 0.008494f
C558 B.n238 VSUBS 0.008494f
C559 B.n239 VSUBS 0.008494f
C560 B.n240 VSUBS 0.008494f
C561 B.n241 VSUBS 0.008494f
C562 B.n242 VSUBS 0.008494f
C563 B.n243 VSUBS 0.008494f
C564 B.n244 VSUBS 0.008494f
C565 B.n245 VSUBS 0.008494f
C566 B.n246 VSUBS 0.008494f
C567 B.n247 VSUBS 0.008494f
C568 B.n248 VSUBS 0.008494f
C569 B.n249 VSUBS 0.008494f
C570 B.n250 VSUBS 0.008494f
C571 B.n251 VSUBS 0.008494f
C572 B.n252 VSUBS 0.008494f
C573 B.n253 VSUBS 0.008494f
C574 B.n254 VSUBS 0.008494f
C575 B.n255 VSUBS 0.008494f
C576 B.n256 VSUBS 0.008494f
C577 B.n257 VSUBS 0.008494f
C578 B.n258 VSUBS 0.008494f
C579 B.n259 VSUBS 0.008494f
C580 B.n260 VSUBS 0.008494f
C581 B.n261 VSUBS 0.008494f
C582 B.n262 VSUBS 0.008494f
C583 B.n263 VSUBS 0.008494f
C584 B.n264 VSUBS 0.008494f
C585 B.n265 VSUBS 0.008494f
C586 B.n266 VSUBS 0.008494f
C587 B.n267 VSUBS 0.008494f
C588 B.n268 VSUBS 0.008494f
C589 B.n269 VSUBS 0.008494f
C590 B.n270 VSUBS 0.008494f
C591 B.n271 VSUBS 0.008494f
C592 B.n272 VSUBS 0.008494f
C593 B.n273 VSUBS 0.008494f
C594 B.n274 VSUBS 0.008494f
C595 B.n275 VSUBS 0.008494f
C596 B.n276 VSUBS 0.008494f
C597 B.n277 VSUBS 0.008494f
C598 B.n278 VSUBS 0.008494f
C599 B.n279 VSUBS 0.008494f
C600 B.n280 VSUBS 0.008494f
C601 B.n281 VSUBS 0.008494f
C602 B.n282 VSUBS 0.008494f
C603 B.n283 VSUBS 0.008494f
C604 B.n284 VSUBS 0.008494f
C605 B.n285 VSUBS 0.008494f
C606 B.n286 VSUBS 0.008494f
C607 B.n287 VSUBS 0.008494f
C608 B.n288 VSUBS 0.008494f
C609 B.n289 VSUBS 0.008494f
C610 B.n290 VSUBS 0.008494f
C611 B.n291 VSUBS 0.008494f
C612 B.n292 VSUBS 0.008494f
C613 B.n293 VSUBS 0.008494f
C614 B.n294 VSUBS 0.008494f
C615 B.n295 VSUBS 0.008494f
C616 B.n296 VSUBS 0.008494f
C617 B.n297 VSUBS 0.008494f
C618 B.n298 VSUBS 0.008494f
C619 B.n299 VSUBS 0.008494f
C620 B.n300 VSUBS 0.008494f
C621 B.n301 VSUBS 0.008494f
C622 B.n302 VSUBS 0.008494f
C623 B.n303 VSUBS 0.008494f
C624 B.n304 VSUBS 0.008494f
C625 B.n305 VSUBS 0.008494f
C626 B.n306 VSUBS 0.008494f
C627 B.n307 VSUBS 0.008494f
C628 B.n308 VSUBS 0.008494f
C629 B.n309 VSUBS 0.008494f
C630 B.n310 VSUBS 0.008494f
C631 B.n311 VSUBS 0.008494f
C632 B.n312 VSUBS 0.008494f
C633 B.n313 VSUBS 0.008494f
C634 B.n314 VSUBS 0.008494f
C635 B.n315 VSUBS 0.008494f
C636 B.n316 VSUBS 0.008494f
C637 B.n317 VSUBS 0.008494f
C638 B.n318 VSUBS 0.008494f
C639 B.n319 VSUBS 0.008494f
C640 B.n320 VSUBS 0.008494f
C641 B.n321 VSUBS 0.008494f
C642 B.n322 VSUBS 0.008494f
C643 B.n323 VSUBS 0.008494f
C644 B.n324 VSUBS 0.008494f
C645 B.n325 VSUBS 0.008494f
C646 B.n326 VSUBS 0.008494f
C647 B.n327 VSUBS 0.008494f
C648 B.n328 VSUBS 0.008494f
C649 B.n329 VSUBS 0.008494f
C650 B.n330 VSUBS 0.008494f
C651 B.n331 VSUBS 0.008494f
C652 B.n332 VSUBS 0.008494f
C653 B.n333 VSUBS 0.008494f
C654 B.n334 VSUBS 0.008494f
C655 B.n335 VSUBS 0.008494f
C656 B.n336 VSUBS 0.008494f
C657 B.n337 VSUBS 0.008494f
C658 B.n338 VSUBS 0.008494f
C659 B.n339 VSUBS 0.008494f
C660 B.n340 VSUBS 0.008494f
C661 B.n341 VSUBS 0.008494f
C662 B.n342 VSUBS 0.008494f
C663 B.n343 VSUBS 0.008494f
C664 B.n344 VSUBS 0.008494f
C665 B.n345 VSUBS 0.008494f
C666 B.n346 VSUBS 0.008494f
C667 B.n347 VSUBS 0.008494f
C668 B.n348 VSUBS 0.008494f
C669 B.n349 VSUBS 0.008494f
C670 B.n350 VSUBS 0.008494f
C671 B.n351 VSUBS 0.008494f
C672 B.n352 VSUBS 0.008494f
C673 B.n353 VSUBS 0.008494f
C674 B.n354 VSUBS 0.008494f
C675 B.n355 VSUBS 0.008494f
C676 B.n356 VSUBS 0.008494f
C677 B.n357 VSUBS 0.008494f
C678 B.n358 VSUBS 0.008494f
C679 B.n359 VSUBS 0.008494f
C680 B.n360 VSUBS 0.008494f
C681 B.n361 VSUBS 0.008494f
C682 B.n362 VSUBS 0.008494f
C683 B.n363 VSUBS 0.008494f
C684 B.n364 VSUBS 0.008494f
C685 B.n365 VSUBS 0.008494f
C686 B.n366 VSUBS 0.008494f
C687 B.n367 VSUBS 0.008494f
C688 B.n368 VSUBS 0.008494f
C689 B.n369 VSUBS 0.008494f
C690 B.n370 VSUBS 0.008494f
C691 B.n371 VSUBS 0.008494f
C692 B.n372 VSUBS 0.008494f
C693 B.n373 VSUBS 0.008494f
C694 B.n374 VSUBS 0.008494f
C695 B.n375 VSUBS 0.008494f
C696 B.n376 VSUBS 0.008494f
C697 B.n377 VSUBS 0.008494f
C698 B.n378 VSUBS 0.008494f
C699 B.n379 VSUBS 0.008494f
C700 B.n380 VSUBS 0.008494f
C701 B.n381 VSUBS 0.008494f
C702 B.n382 VSUBS 0.008494f
C703 B.n383 VSUBS 0.008494f
C704 B.n384 VSUBS 0.008494f
C705 B.n385 VSUBS 0.008494f
C706 B.n386 VSUBS 0.008494f
C707 B.n387 VSUBS 0.008494f
C708 B.n388 VSUBS 0.008494f
C709 B.n389 VSUBS 0.02044f
C710 B.n390 VSUBS 0.021283f
C711 B.n391 VSUBS 0.021283f
C712 B.n392 VSUBS 0.008494f
C713 B.n393 VSUBS 0.008494f
C714 B.n394 VSUBS 0.008494f
C715 B.n395 VSUBS 0.008494f
C716 B.n396 VSUBS 0.008494f
C717 B.n397 VSUBS 0.008494f
C718 B.n398 VSUBS 0.008494f
C719 B.n399 VSUBS 0.008494f
C720 B.n400 VSUBS 0.008494f
C721 B.n401 VSUBS 0.008494f
C722 B.n402 VSUBS 0.008494f
C723 B.n403 VSUBS 0.008494f
C724 B.n404 VSUBS 0.008494f
C725 B.n405 VSUBS 0.008494f
C726 B.n406 VSUBS 0.008494f
C727 B.n407 VSUBS 0.008494f
C728 B.n408 VSUBS 0.008494f
C729 B.n409 VSUBS 0.008494f
C730 B.n410 VSUBS 0.008494f
C731 B.n411 VSUBS 0.008494f
C732 B.n412 VSUBS 0.008494f
C733 B.n413 VSUBS 0.008494f
C734 B.n414 VSUBS 0.008494f
C735 B.n415 VSUBS 0.008494f
C736 B.n416 VSUBS 0.008494f
C737 B.n417 VSUBS 0.008494f
C738 B.n418 VSUBS 0.008494f
C739 B.n419 VSUBS 0.008494f
C740 B.n420 VSUBS 0.008494f
C741 B.n421 VSUBS 0.008494f
C742 B.n422 VSUBS 0.008494f
C743 B.n423 VSUBS 0.008494f
C744 B.n424 VSUBS 0.008494f
C745 B.n425 VSUBS 0.008494f
C746 B.n426 VSUBS 0.008494f
C747 B.n427 VSUBS 0.008494f
C748 B.n428 VSUBS 0.008494f
C749 B.n429 VSUBS 0.008494f
C750 B.n430 VSUBS 0.008494f
C751 B.n431 VSUBS 0.008494f
C752 B.n432 VSUBS 0.008494f
C753 B.n433 VSUBS 0.008494f
C754 B.n434 VSUBS 0.008494f
C755 B.n435 VSUBS 0.008494f
C756 B.n436 VSUBS 0.008494f
C757 B.n437 VSUBS 0.008494f
C758 B.n438 VSUBS 0.008494f
C759 B.n439 VSUBS 0.008494f
C760 B.n440 VSUBS 0.008494f
C761 B.n441 VSUBS 0.008494f
C762 B.n442 VSUBS 0.008494f
C763 B.n443 VSUBS 0.008494f
C764 B.n444 VSUBS 0.008494f
C765 B.n445 VSUBS 0.008494f
C766 B.n446 VSUBS 0.008494f
C767 B.n447 VSUBS 0.008494f
C768 B.n448 VSUBS 0.008494f
C769 B.n449 VSUBS 0.008494f
C770 B.n450 VSUBS 0.008494f
C771 B.n451 VSUBS 0.008494f
C772 B.n452 VSUBS 0.008494f
C773 B.n453 VSUBS 0.008494f
C774 B.n454 VSUBS 0.008494f
C775 B.n455 VSUBS 0.008494f
C776 B.n456 VSUBS 0.007995f
C777 B.n457 VSUBS 0.008494f
C778 B.n458 VSUBS 0.008494f
C779 B.n459 VSUBS 0.004747f
C780 B.n460 VSUBS 0.008494f
C781 B.n461 VSUBS 0.008494f
C782 B.n462 VSUBS 0.008494f
C783 B.n463 VSUBS 0.008494f
C784 B.n464 VSUBS 0.008494f
C785 B.n465 VSUBS 0.008494f
C786 B.n466 VSUBS 0.008494f
C787 B.n467 VSUBS 0.008494f
C788 B.n468 VSUBS 0.008494f
C789 B.n469 VSUBS 0.008494f
C790 B.n470 VSUBS 0.008494f
C791 B.n471 VSUBS 0.008494f
C792 B.n472 VSUBS 0.004747f
C793 B.n473 VSUBS 0.019681f
C794 B.n474 VSUBS 0.007995f
C795 B.n475 VSUBS 0.008494f
C796 B.n476 VSUBS 0.008494f
C797 B.n477 VSUBS 0.008494f
C798 B.n478 VSUBS 0.008494f
C799 B.n479 VSUBS 0.008494f
C800 B.n480 VSUBS 0.008494f
C801 B.n481 VSUBS 0.008494f
C802 B.n482 VSUBS 0.008494f
C803 B.n483 VSUBS 0.008494f
C804 B.n484 VSUBS 0.008494f
C805 B.n485 VSUBS 0.008494f
C806 B.n486 VSUBS 0.008494f
C807 B.n487 VSUBS 0.008494f
C808 B.n488 VSUBS 0.008494f
C809 B.n489 VSUBS 0.008494f
C810 B.n490 VSUBS 0.008494f
C811 B.n491 VSUBS 0.008494f
C812 B.n492 VSUBS 0.008494f
C813 B.n493 VSUBS 0.008494f
C814 B.n494 VSUBS 0.008494f
C815 B.n495 VSUBS 0.008494f
C816 B.n496 VSUBS 0.008494f
C817 B.n497 VSUBS 0.008494f
C818 B.n498 VSUBS 0.008494f
C819 B.n499 VSUBS 0.008494f
C820 B.n500 VSUBS 0.008494f
C821 B.n501 VSUBS 0.008494f
C822 B.n502 VSUBS 0.008494f
C823 B.n503 VSUBS 0.008494f
C824 B.n504 VSUBS 0.008494f
C825 B.n505 VSUBS 0.008494f
C826 B.n506 VSUBS 0.008494f
C827 B.n507 VSUBS 0.008494f
C828 B.n508 VSUBS 0.008494f
C829 B.n509 VSUBS 0.008494f
C830 B.n510 VSUBS 0.008494f
C831 B.n511 VSUBS 0.008494f
C832 B.n512 VSUBS 0.008494f
C833 B.n513 VSUBS 0.008494f
C834 B.n514 VSUBS 0.008494f
C835 B.n515 VSUBS 0.008494f
C836 B.n516 VSUBS 0.008494f
C837 B.n517 VSUBS 0.008494f
C838 B.n518 VSUBS 0.008494f
C839 B.n519 VSUBS 0.008494f
C840 B.n520 VSUBS 0.008494f
C841 B.n521 VSUBS 0.008494f
C842 B.n522 VSUBS 0.008494f
C843 B.n523 VSUBS 0.008494f
C844 B.n524 VSUBS 0.008494f
C845 B.n525 VSUBS 0.008494f
C846 B.n526 VSUBS 0.008494f
C847 B.n527 VSUBS 0.008494f
C848 B.n528 VSUBS 0.008494f
C849 B.n529 VSUBS 0.008494f
C850 B.n530 VSUBS 0.008494f
C851 B.n531 VSUBS 0.008494f
C852 B.n532 VSUBS 0.008494f
C853 B.n533 VSUBS 0.008494f
C854 B.n534 VSUBS 0.008494f
C855 B.n535 VSUBS 0.008494f
C856 B.n536 VSUBS 0.008494f
C857 B.n537 VSUBS 0.008494f
C858 B.n538 VSUBS 0.008494f
C859 B.n539 VSUBS 0.008494f
C860 B.n540 VSUBS 0.021283f
C861 B.n541 VSUBS 0.021283f
C862 B.n542 VSUBS 0.02044f
C863 B.n543 VSUBS 0.008494f
C864 B.n544 VSUBS 0.008494f
C865 B.n545 VSUBS 0.008494f
C866 B.n546 VSUBS 0.008494f
C867 B.n547 VSUBS 0.008494f
C868 B.n548 VSUBS 0.008494f
C869 B.n549 VSUBS 0.008494f
C870 B.n550 VSUBS 0.008494f
C871 B.n551 VSUBS 0.008494f
C872 B.n552 VSUBS 0.008494f
C873 B.n553 VSUBS 0.008494f
C874 B.n554 VSUBS 0.008494f
C875 B.n555 VSUBS 0.008494f
C876 B.n556 VSUBS 0.008494f
C877 B.n557 VSUBS 0.008494f
C878 B.n558 VSUBS 0.008494f
C879 B.n559 VSUBS 0.008494f
C880 B.n560 VSUBS 0.008494f
C881 B.n561 VSUBS 0.008494f
C882 B.n562 VSUBS 0.008494f
C883 B.n563 VSUBS 0.008494f
C884 B.n564 VSUBS 0.008494f
C885 B.n565 VSUBS 0.008494f
C886 B.n566 VSUBS 0.008494f
C887 B.n567 VSUBS 0.008494f
C888 B.n568 VSUBS 0.008494f
C889 B.n569 VSUBS 0.008494f
C890 B.n570 VSUBS 0.008494f
C891 B.n571 VSUBS 0.008494f
C892 B.n572 VSUBS 0.008494f
C893 B.n573 VSUBS 0.008494f
C894 B.n574 VSUBS 0.008494f
C895 B.n575 VSUBS 0.008494f
C896 B.n576 VSUBS 0.008494f
C897 B.n577 VSUBS 0.008494f
C898 B.n578 VSUBS 0.008494f
C899 B.n579 VSUBS 0.008494f
C900 B.n580 VSUBS 0.008494f
C901 B.n581 VSUBS 0.008494f
C902 B.n582 VSUBS 0.008494f
C903 B.n583 VSUBS 0.008494f
C904 B.n584 VSUBS 0.008494f
C905 B.n585 VSUBS 0.008494f
C906 B.n586 VSUBS 0.008494f
C907 B.n587 VSUBS 0.008494f
C908 B.n588 VSUBS 0.008494f
C909 B.n589 VSUBS 0.008494f
C910 B.n590 VSUBS 0.008494f
C911 B.n591 VSUBS 0.008494f
C912 B.n592 VSUBS 0.008494f
C913 B.n593 VSUBS 0.008494f
C914 B.n594 VSUBS 0.008494f
C915 B.n595 VSUBS 0.008494f
C916 B.n596 VSUBS 0.008494f
C917 B.n597 VSUBS 0.008494f
C918 B.n598 VSUBS 0.008494f
C919 B.n599 VSUBS 0.008494f
C920 B.n600 VSUBS 0.008494f
C921 B.n601 VSUBS 0.008494f
C922 B.n602 VSUBS 0.008494f
C923 B.n603 VSUBS 0.008494f
C924 B.n604 VSUBS 0.008494f
C925 B.n605 VSUBS 0.008494f
C926 B.n606 VSUBS 0.008494f
C927 B.n607 VSUBS 0.008494f
C928 B.n608 VSUBS 0.008494f
C929 B.n609 VSUBS 0.008494f
C930 B.n610 VSUBS 0.008494f
C931 B.n611 VSUBS 0.008494f
C932 B.n612 VSUBS 0.008494f
C933 B.n613 VSUBS 0.008494f
C934 B.n614 VSUBS 0.008494f
C935 B.n615 VSUBS 0.008494f
C936 B.n616 VSUBS 0.008494f
C937 B.n617 VSUBS 0.008494f
C938 B.n618 VSUBS 0.008494f
C939 B.n619 VSUBS 0.008494f
C940 B.n620 VSUBS 0.008494f
C941 B.n621 VSUBS 0.008494f
C942 B.n622 VSUBS 0.008494f
C943 B.n623 VSUBS 0.008494f
C944 B.n624 VSUBS 0.008494f
C945 B.n625 VSUBS 0.008494f
C946 B.n626 VSUBS 0.008494f
C947 B.n627 VSUBS 0.008494f
C948 B.n628 VSUBS 0.008494f
C949 B.n629 VSUBS 0.008494f
C950 B.n630 VSUBS 0.008494f
C951 B.n631 VSUBS 0.008494f
C952 B.n632 VSUBS 0.008494f
C953 B.n633 VSUBS 0.008494f
C954 B.n634 VSUBS 0.008494f
C955 B.n635 VSUBS 0.008494f
C956 B.n636 VSUBS 0.008494f
C957 B.n637 VSUBS 0.008494f
C958 B.n638 VSUBS 0.008494f
C959 B.n639 VSUBS 0.008494f
C960 B.n640 VSUBS 0.008494f
C961 B.n641 VSUBS 0.008494f
C962 B.n642 VSUBS 0.008494f
C963 B.n643 VSUBS 0.008494f
C964 B.n644 VSUBS 0.008494f
C965 B.n645 VSUBS 0.008494f
C966 B.n646 VSUBS 0.008494f
C967 B.n647 VSUBS 0.008494f
C968 B.n648 VSUBS 0.008494f
C969 B.n649 VSUBS 0.008494f
C970 B.n650 VSUBS 0.008494f
C971 B.n651 VSUBS 0.008494f
C972 B.n652 VSUBS 0.008494f
C973 B.n653 VSUBS 0.008494f
C974 B.n654 VSUBS 0.008494f
C975 B.n655 VSUBS 0.008494f
C976 B.n656 VSUBS 0.008494f
C977 B.n657 VSUBS 0.008494f
C978 B.n658 VSUBS 0.008494f
C979 B.n659 VSUBS 0.008494f
C980 B.n660 VSUBS 0.008494f
C981 B.n661 VSUBS 0.008494f
C982 B.n662 VSUBS 0.008494f
C983 B.n663 VSUBS 0.008494f
C984 B.n664 VSUBS 0.008494f
C985 B.n665 VSUBS 0.008494f
C986 B.n666 VSUBS 0.008494f
C987 B.n667 VSUBS 0.008494f
C988 B.n668 VSUBS 0.008494f
C989 B.n669 VSUBS 0.008494f
C990 B.n670 VSUBS 0.008494f
C991 B.n671 VSUBS 0.008494f
C992 B.n672 VSUBS 0.008494f
C993 B.n673 VSUBS 0.008494f
C994 B.n674 VSUBS 0.008494f
C995 B.n675 VSUBS 0.008494f
C996 B.n676 VSUBS 0.008494f
C997 B.n677 VSUBS 0.008494f
C998 B.n678 VSUBS 0.008494f
C999 B.n679 VSUBS 0.008494f
C1000 B.n680 VSUBS 0.008494f
C1001 B.n681 VSUBS 0.008494f
C1002 B.n682 VSUBS 0.008494f
C1003 B.n683 VSUBS 0.008494f
C1004 B.n684 VSUBS 0.008494f
C1005 B.n685 VSUBS 0.008494f
C1006 B.n686 VSUBS 0.008494f
C1007 B.n687 VSUBS 0.008494f
C1008 B.n688 VSUBS 0.008494f
C1009 B.n689 VSUBS 0.008494f
C1010 B.n690 VSUBS 0.008494f
C1011 B.n691 VSUBS 0.008494f
C1012 B.n692 VSUBS 0.008494f
C1013 B.n693 VSUBS 0.008494f
C1014 B.n694 VSUBS 0.008494f
C1015 B.n695 VSUBS 0.008494f
C1016 B.n696 VSUBS 0.008494f
C1017 B.n697 VSUBS 0.008494f
C1018 B.n698 VSUBS 0.008494f
C1019 B.n699 VSUBS 0.008494f
C1020 B.n700 VSUBS 0.008494f
C1021 B.n701 VSUBS 0.008494f
C1022 B.n702 VSUBS 0.008494f
C1023 B.n703 VSUBS 0.008494f
C1024 B.n704 VSUBS 0.008494f
C1025 B.n705 VSUBS 0.008494f
C1026 B.n706 VSUBS 0.008494f
C1027 B.n707 VSUBS 0.008494f
C1028 B.n708 VSUBS 0.008494f
C1029 B.n709 VSUBS 0.008494f
C1030 B.n710 VSUBS 0.008494f
C1031 B.n711 VSUBS 0.008494f
C1032 B.n712 VSUBS 0.008494f
C1033 B.n713 VSUBS 0.008494f
C1034 B.n714 VSUBS 0.008494f
C1035 B.n715 VSUBS 0.008494f
C1036 B.n716 VSUBS 0.008494f
C1037 B.n717 VSUBS 0.008494f
C1038 B.n718 VSUBS 0.008494f
C1039 B.n719 VSUBS 0.008494f
C1040 B.n720 VSUBS 0.008494f
C1041 B.n721 VSUBS 0.008494f
C1042 B.n722 VSUBS 0.008494f
C1043 B.n723 VSUBS 0.008494f
C1044 B.n724 VSUBS 0.008494f
C1045 B.n725 VSUBS 0.008494f
C1046 B.n726 VSUBS 0.008494f
C1047 B.n727 VSUBS 0.008494f
C1048 B.n728 VSUBS 0.008494f
C1049 B.n729 VSUBS 0.008494f
C1050 B.n730 VSUBS 0.008494f
C1051 B.n731 VSUBS 0.008494f
C1052 B.n732 VSUBS 0.008494f
C1053 B.n733 VSUBS 0.008494f
C1054 B.n734 VSUBS 0.008494f
C1055 B.n735 VSUBS 0.008494f
C1056 B.n736 VSUBS 0.008494f
C1057 B.n737 VSUBS 0.008494f
C1058 B.n738 VSUBS 0.008494f
C1059 B.n739 VSUBS 0.008494f
C1060 B.n740 VSUBS 0.008494f
C1061 B.n741 VSUBS 0.008494f
C1062 B.n742 VSUBS 0.008494f
C1063 B.n743 VSUBS 0.008494f
C1064 B.n744 VSUBS 0.008494f
C1065 B.n745 VSUBS 0.008494f
C1066 B.n746 VSUBS 0.008494f
C1067 B.n747 VSUBS 0.008494f
C1068 B.n748 VSUBS 0.008494f
C1069 B.n749 VSUBS 0.008494f
C1070 B.n750 VSUBS 0.008494f
C1071 B.n751 VSUBS 0.008494f
C1072 B.n752 VSUBS 0.008494f
C1073 B.n753 VSUBS 0.008494f
C1074 B.n754 VSUBS 0.008494f
C1075 B.n755 VSUBS 0.008494f
C1076 B.n756 VSUBS 0.008494f
C1077 B.n757 VSUBS 0.008494f
C1078 B.n758 VSUBS 0.008494f
C1079 B.n759 VSUBS 0.008494f
C1080 B.n760 VSUBS 0.008494f
C1081 B.n761 VSUBS 0.008494f
C1082 B.n762 VSUBS 0.008494f
C1083 B.n763 VSUBS 0.008494f
C1084 B.n764 VSUBS 0.008494f
C1085 B.n765 VSUBS 0.008494f
C1086 B.n766 VSUBS 0.008494f
C1087 B.n767 VSUBS 0.008494f
C1088 B.n768 VSUBS 0.008494f
C1089 B.n769 VSUBS 0.008494f
C1090 B.n770 VSUBS 0.008494f
C1091 B.n771 VSUBS 0.008494f
C1092 B.n772 VSUBS 0.008494f
C1093 B.n773 VSUBS 0.008494f
C1094 B.n774 VSUBS 0.008494f
C1095 B.n775 VSUBS 0.008494f
C1096 B.n776 VSUBS 0.008494f
C1097 B.n777 VSUBS 0.008494f
C1098 B.n778 VSUBS 0.008494f
C1099 B.n779 VSUBS 0.008494f
C1100 B.n780 VSUBS 0.008494f
C1101 B.n781 VSUBS 0.008494f
C1102 B.n782 VSUBS 0.02044f
C1103 B.n783 VSUBS 0.021283f
C1104 B.n784 VSUBS 0.020349f
C1105 B.n785 VSUBS 0.008494f
C1106 B.n786 VSUBS 0.008494f
C1107 B.n787 VSUBS 0.008494f
C1108 B.n788 VSUBS 0.008494f
C1109 B.n789 VSUBS 0.008494f
C1110 B.n790 VSUBS 0.008494f
C1111 B.n791 VSUBS 0.008494f
C1112 B.n792 VSUBS 0.008494f
C1113 B.n793 VSUBS 0.008494f
C1114 B.n794 VSUBS 0.008494f
C1115 B.n795 VSUBS 0.008494f
C1116 B.n796 VSUBS 0.008494f
C1117 B.n797 VSUBS 0.008494f
C1118 B.n798 VSUBS 0.008494f
C1119 B.n799 VSUBS 0.008494f
C1120 B.n800 VSUBS 0.008494f
C1121 B.n801 VSUBS 0.008494f
C1122 B.n802 VSUBS 0.008494f
C1123 B.n803 VSUBS 0.008494f
C1124 B.n804 VSUBS 0.008494f
C1125 B.n805 VSUBS 0.008494f
C1126 B.n806 VSUBS 0.008494f
C1127 B.n807 VSUBS 0.008494f
C1128 B.n808 VSUBS 0.008494f
C1129 B.n809 VSUBS 0.008494f
C1130 B.n810 VSUBS 0.008494f
C1131 B.n811 VSUBS 0.008494f
C1132 B.n812 VSUBS 0.008494f
C1133 B.n813 VSUBS 0.008494f
C1134 B.n814 VSUBS 0.008494f
C1135 B.n815 VSUBS 0.008494f
C1136 B.n816 VSUBS 0.008494f
C1137 B.n817 VSUBS 0.008494f
C1138 B.n818 VSUBS 0.008494f
C1139 B.n819 VSUBS 0.008494f
C1140 B.n820 VSUBS 0.008494f
C1141 B.n821 VSUBS 0.008494f
C1142 B.n822 VSUBS 0.008494f
C1143 B.n823 VSUBS 0.008494f
C1144 B.n824 VSUBS 0.008494f
C1145 B.n825 VSUBS 0.008494f
C1146 B.n826 VSUBS 0.008494f
C1147 B.n827 VSUBS 0.008494f
C1148 B.n828 VSUBS 0.008494f
C1149 B.n829 VSUBS 0.008494f
C1150 B.n830 VSUBS 0.008494f
C1151 B.n831 VSUBS 0.008494f
C1152 B.n832 VSUBS 0.008494f
C1153 B.n833 VSUBS 0.008494f
C1154 B.n834 VSUBS 0.008494f
C1155 B.n835 VSUBS 0.008494f
C1156 B.n836 VSUBS 0.008494f
C1157 B.n837 VSUBS 0.008494f
C1158 B.n838 VSUBS 0.008494f
C1159 B.n839 VSUBS 0.008494f
C1160 B.n840 VSUBS 0.008494f
C1161 B.n841 VSUBS 0.008494f
C1162 B.n842 VSUBS 0.008494f
C1163 B.n843 VSUBS 0.008494f
C1164 B.n844 VSUBS 0.008494f
C1165 B.n845 VSUBS 0.008494f
C1166 B.n846 VSUBS 0.008494f
C1167 B.n847 VSUBS 0.008494f
C1168 B.n848 VSUBS 0.008494f
C1169 B.n849 VSUBS 0.008494f
C1170 B.n850 VSUBS 0.007995f
C1171 B.n851 VSUBS 0.019681f
C1172 B.n852 VSUBS 0.004747f
C1173 B.n853 VSUBS 0.008494f
C1174 B.n854 VSUBS 0.008494f
C1175 B.n855 VSUBS 0.008494f
C1176 B.n856 VSUBS 0.008494f
C1177 B.n857 VSUBS 0.008494f
C1178 B.n858 VSUBS 0.008494f
C1179 B.n859 VSUBS 0.008494f
C1180 B.n860 VSUBS 0.008494f
C1181 B.n861 VSUBS 0.008494f
C1182 B.n862 VSUBS 0.008494f
C1183 B.n863 VSUBS 0.008494f
C1184 B.n864 VSUBS 0.008494f
C1185 B.n865 VSUBS 0.004747f
C1186 B.n866 VSUBS 0.008494f
C1187 B.n867 VSUBS 0.008494f
C1188 B.n868 VSUBS 0.008494f
C1189 B.n869 VSUBS 0.008494f
C1190 B.n870 VSUBS 0.008494f
C1191 B.n871 VSUBS 0.008494f
C1192 B.n872 VSUBS 0.008494f
C1193 B.n873 VSUBS 0.008494f
C1194 B.n874 VSUBS 0.008494f
C1195 B.n875 VSUBS 0.008494f
C1196 B.n876 VSUBS 0.008494f
C1197 B.n877 VSUBS 0.008494f
C1198 B.n878 VSUBS 0.008494f
C1199 B.n879 VSUBS 0.008494f
C1200 B.n880 VSUBS 0.008494f
C1201 B.n881 VSUBS 0.008494f
C1202 B.n882 VSUBS 0.008494f
C1203 B.n883 VSUBS 0.008494f
C1204 B.n884 VSUBS 0.008494f
C1205 B.n885 VSUBS 0.008494f
C1206 B.n886 VSUBS 0.008494f
C1207 B.n887 VSUBS 0.008494f
C1208 B.n888 VSUBS 0.008494f
C1209 B.n889 VSUBS 0.008494f
C1210 B.n890 VSUBS 0.008494f
C1211 B.n891 VSUBS 0.008494f
C1212 B.n892 VSUBS 0.008494f
C1213 B.n893 VSUBS 0.008494f
C1214 B.n894 VSUBS 0.008494f
C1215 B.n895 VSUBS 0.008494f
C1216 B.n896 VSUBS 0.008494f
C1217 B.n897 VSUBS 0.008494f
C1218 B.n898 VSUBS 0.008494f
C1219 B.n899 VSUBS 0.008494f
C1220 B.n900 VSUBS 0.008494f
C1221 B.n901 VSUBS 0.008494f
C1222 B.n902 VSUBS 0.008494f
C1223 B.n903 VSUBS 0.008494f
C1224 B.n904 VSUBS 0.008494f
C1225 B.n905 VSUBS 0.008494f
C1226 B.n906 VSUBS 0.008494f
C1227 B.n907 VSUBS 0.008494f
C1228 B.n908 VSUBS 0.008494f
C1229 B.n909 VSUBS 0.008494f
C1230 B.n910 VSUBS 0.008494f
C1231 B.n911 VSUBS 0.008494f
C1232 B.n912 VSUBS 0.008494f
C1233 B.n913 VSUBS 0.008494f
C1234 B.n914 VSUBS 0.008494f
C1235 B.n915 VSUBS 0.008494f
C1236 B.n916 VSUBS 0.008494f
C1237 B.n917 VSUBS 0.008494f
C1238 B.n918 VSUBS 0.008494f
C1239 B.n919 VSUBS 0.008494f
C1240 B.n920 VSUBS 0.008494f
C1241 B.n921 VSUBS 0.008494f
C1242 B.n922 VSUBS 0.008494f
C1243 B.n923 VSUBS 0.008494f
C1244 B.n924 VSUBS 0.008494f
C1245 B.n925 VSUBS 0.008494f
C1246 B.n926 VSUBS 0.008494f
C1247 B.n927 VSUBS 0.008494f
C1248 B.n928 VSUBS 0.008494f
C1249 B.n929 VSUBS 0.008494f
C1250 B.n930 VSUBS 0.008494f
C1251 B.n931 VSUBS 0.008494f
C1252 B.n932 VSUBS 0.008494f
C1253 B.n933 VSUBS 0.021283f
C1254 B.n934 VSUBS 0.02044f
C1255 B.n935 VSUBS 0.02044f
C1256 B.n936 VSUBS 0.008494f
C1257 B.n937 VSUBS 0.008494f
C1258 B.n938 VSUBS 0.008494f
C1259 B.n939 VSUBS 0.008494f
C1260 B.n940 VSUBS 0.008494f
C1261 B.n941 VSUBS 0.008494f
C1262 B.n942 VSUBS 0.008494f
C1263 B.n943 VSUBS 0.008494f
C1264 B.n944 VSUBS 0.008494f
C1265 B.n945 VSUBS 0.008494f
C1266 B.n946 VSUBS 0.008494f
C1267 B.n947 VSUBS 0.008494f
C1268 B.n948 VSUBS 0.008494f
C1269 B.n949 VSUBS 0.008494f
C1270 B.n950 VSUBS 0.008494f
C1271 B.n951 VSUBS 0.008494f
C1272 B.n952 VSUBS 0.008494f
C1273 B.n953 VSUBS 0.008494f
C1274 B.n954 VSUBS 0.008494f
C1275 B.n955 VSUBS 0.008494f
C1276 B.n956 VSUBS 0.008494f
C1277 B.n957 VSUBS 0.008494f
C1278 B.n958 VSUBS 0.008494f
C1279 B.n959 VSUBS 0.008494f
C1280 B.n960 VSUBS 0.008494f
C1281 B.n961 VSUBS 0.008494f
C1282 B.n962 VSUBS 0.008494f
C1283 B.n963 VSUBS 0.008494f
C1284 B.n964 VSUBS 0.008494f
C1285 B.n965 VSUBS 0.008494f
C1286 B.n966 VSUBS 0.008494f
C1287 B.n967 VSUBS 0.008494f
C1288 B.n968 VSUBS 0.008494f
C1289 B.n969 VSUBS 0.008494f
C1290 B.n970 VSUBS 0.008494f
C1291 B.n971 VSUBS 0.008494f
C1292 B.n972 VSUBS 0.008494f
C1293 B.n973 VSUBS 0.008494f
C1294 B.n974 VSUBS 0.008494f
C1295 B.n975 VSUBS 0.008494f
C1296 B.n976 VSUBS 0.008494f
C1297 B.n977 VSUBS 0.008494f
C1298 B.n978 VSUBS 0.008494f
C1299 B.n979 VSUBS 0.008494f
C1300 B.n980 VSUBS 0.008494f
C1301 B.n981 VSUBS 0.008494f
C1302 B.n982 VSUBS 0.008494f
C1303 B.n983 VSUBS 0.008494f
C1304 B.n984 VSUBS 0.008494f
C1305 B.n985 VSUBS 0.008494f
C1306 B.n986 VSUBS 0.008494f
C1307 B.n987 VSUBS 0.008494f
C1308 B.n988 VSUBS 0.008494f
C1309 B.n989 VSUBS 0.008494f
C1310 B.n990 VSUBS 0.008494f
C1311 B.n991 VSUBS 0.008494f
C1312 B.n992 VSUBS 0.008494f
C1313 B.n993 VSUBS 0.008494f
C1314 B.n994 VSUBS 0.008494f
C1315 B.n995 VSUBS 0.008494f
C1316 B.n996 VSUBS 0.008494f
C1317 B.n997 VSUBS 0.008494f
C1318 B.n998 VSUBS 0.008494f
C1319 B.n999 VSUBS 0.008494f
C1320 B.n1000 VSUBS 0.008494f
C1321 B.n1001 VSUBS 0.008494f
C1322 B.n1002 VSUBS 0.008494f
C1323 B.n1003 VSUBS 0.008494f
C1324 B.n1004 VSUBS 0.008494f
C1325 B.n1005 VSUBS 0.008494f
C1326 B.n1006 VSUBS 0.008494f
C1327 B.n1007 VSUBS 0.008494f
C1328 B.n1008 VSUBS 0.008494f
C1329 B.n1009 VSUBS 0.008494f
C1330 B.n1010 VSUBS 0.008494f
C1331 B.n1011 VSUBS 0.008494f
C1332 B.n1012 VSUBS 0.008494f
C1333 B.n1013 VSUBS 0.008494f
C1334 B.n1014 VSUBS 0.008494f
C1335 B.n1015 VSUBS 0.008494f
C1336 B.n1016 VSUBS 0.008494f
C1337 B.n1017 VSUBS 0.008494f
C1338 B.n1018 VSUBS 0.008494f
C1339 B.n1019 VSUBS 0.008494f
C1340 B.n1020 VSUBS 0.008494f
C1341 B.n1021 VSUBS 0.008494f
C1342 B.n1022 VSUBS 0.008494f
C1343 B.n1023 VSUBS 0.008494f
C1344 B.n1024 VSUBS 0.008494f
C1345 B.n1025 VSUBS 0.008494f
C1346 B.n1026 VSUBS 0.008494f
C1347 B.n1027 VSUBS 0.008494f
C1348 B.n1028 VSUBS 0.008494f
C1349 B.n1029 VSUBS 0.008494f
C1350 B.n1030 VSUBS 0.008494f
C1351 B.n1031 VSUBS 0.008494f
C1352 B.n1032 VSUBS 0.008494f
C1353 B.n1033 VSUBS 0.008494f
C1354 B.n1034 VSUBS 0.008494f
C1355 B.n1035 VSUBS 0.008494f
C1356 B.n1036 VSUBS 0.008494f
C1357 B.n1037 VSUBS 0.008494f
C1358 B.n1038 VSUBS 0.008494f
C1359 B.n1039 VSUBS 0.008494f
C1360 B.n1040 VSUBS 0.008494f
C1361 B.n1041 VSUBS 0.008494f
C1362 B.n1042 VSUBS 0.008494f
C1363 B.n1043 VSUBS 0.008494f
C1364 B.n1044 VSUBS 0.008494f
C1365 B.n1045 VSUBS 0.008494f
C1366 B.n1046 VSUBS 0.008494f
C1367 B.n1047 VSUBS 0.008494f
C1368 B.n1048 VSUBS 0.008494f
C1369 B.n1049 VSUBS 0.008494f
C1370 B.n1050 VSUBS 0.008494f
C1371 B.n1051 VSUBS 0.008494f
C1372 B.n1052 VSUBS 0.008494f
C1373 B.n1053 VSUBS 0.008494f
C1374 B.n1054 VSUBS 0.008494f
C1375 B.n1055 VSUBS 0.019235f
C1376 VDD1.n0 VSUBS 0.03173f
C1377 VDD1.n1 VSUBS 0.030662f
C1378 VDD1.n2 VSUBS 0.016477f
C1379 VDD1.n3 VSUBS 0.038945f
C1380 VDD1.n4 VSUBS 0.017446f
C1381 VDD1.n5 VSUBS 0.030662f
C1382 VDD1.n6 VSUBS 0.016477f
C1383 VDD1.n7 VSUBS 0.038945f
C1384 VDD1.n8 VSUBS 0.017446f
C1385 VDD1.n9 VSUBS 0.030662f
C1386 VDD1.n10 VSUBS 0.016477f
C1387 VDD1.n11 VSUBS 0.038945f
C1388 VDD1.n12 VSUBS 0.017446f
C1389 VDD1.n13 VSUBS 0.030662f
C1390 VDD1.n14 VSUBS 0.016477f
C1391 VDD1.n15 VSUBS 0.038945f
C1392 VDD1.n16 VSUBS 0.017446f
C1393 VDD1.n17 VSUBS 0.030662f
C1394 VDD1.n18 VSUBS 0.016477f
C1395 VDD1.n19 VSUBS 0.038945f
C1396 VDD1.n20 VSUBS 0.017446f
C1397 VDD1.n21 VSUBS 1.71704f
C1398 VDD1.n22 VSUBS 0.016477f
C1399 VDD1.t2 VSUBS 0.083242f
C1400 VDD1.n23 VSUBS 0.200498f
C1401 VDD1.n24 VSUBS 0.024775f
C1402 VDD1.n25 VSUBS 0.029209f
C1403 VDD1.n26 VSUBS 0.038945f
C1404 VDD1.n27 VSUBS 0.017446f
C1405 VDD1.n28 VSUBS 0.016477f
C1406 VDD1.n29 VSUBS 0.030662f
C1407 VDD1.n30 VSUBS 0.030662f
C1408 VDD1.n31 VSUBS 0.016477f
C1409 VDD1.n32 VSUBS 0.017446f
C1410 VDD1.n33 VSUBS 0.038945f
C1411 VDD1.n34 VSUBS 0.038945f
C1412 VDD1.n35 VSUBS 0.017446f
C1413 VDD1.n36 VSUBS 0.016477f
C1414 VDD1.n37 VSUBS 0.030662f
C1415 VDD1.n38 VSUBS 0.030662f
C1416 VDD1.n39 VSUBS 0.016477f
C1417 VDD1.n40 VSUBS 0.017446f
C1418 VDD1.n41 VSUBS 0.038945f
C1419 VDD1.n42 VSUBS 0.038945f
C1420 VDD1.n43 VSUBS 0.017446f
C1421 VDD1.n44 VSUBS 0.016477f
C1422 VDD1.n45 VSUBS 0.030662f
C1423 VDD1.n46 VSUBS 0.030662f
C1424 VDD1.n47 VSUBS 0.016477f
C1425 VDD1.n48 VSUBS 0.017446f
C1426 VDD1.n49 VSUBS 0.038945f
C1427 VDD1.n50 VSUBS 0.038945f
C1428 VDD1.n51 VSUBS 0.017446f
C1429 VDD1.n52 VSUBS 0.016477f
C1430 VDD1.n53 VSUBS 0.030662f
C1431 VDD1.n54 VSUBS 0.030662f
C1432 VDD1.n55 VSUBS 0.016477f
C1433 VDD1.n56 VSUBS 0.017446f
C1434 VDD1.n57 VSUBS 0.038945f
C1435 VDD1.n58 VSUBS 0.038945f
C1436 VDD1.n59 VSUBS 0.017446f
C1437 VDD1.n60 VSUBS 0.016477f
C1438 VDD1.n61 VSUBS 0.030662f
C1439 VDD1.n62 VSUBS 0.030662f
C1440 VDD1.n63 VSUBS 0.016477f
C1441 VDD1.n64 VSUBS 0.017446f
C1442 VDD1.n65 VSUBS 0.038945f
C1443 VDD1.n66 VSUBS 0.094362f
C1444 VDD1.n67 VSUBS 0.017446f
C1445 VDD1.n68 VSUBS 0.032356f
C1446 VDD1.n69 VSUBS 0.073807f
C1447 VDD1.n70 VSUBS 0.118874f
C1448 VDD1.t6 VSUBS 0.321537f
C1449 VDD1.t5 VSUBS 0.321537f
C1450 VDD1.n71 VSUBS 2.56873f
C1451 VDD1.n72 VSUBS 1.3904f
C1452 VDD1.n73 VSUBS 0.03173f
C1453 VDD1.n74 VSUBS 0.030662f
C1454 VDD1.n75 VSUBS 0.016477f
C1455 VDD1.n76 VSUBS 0.038945f
C1456 VDD1.n77 VSUBS 0.017446f
C1457 VDD1.n78 VSUBS 0.030662f
C1458 VDD1.n79 VSUBS 0.016477f
C1459 VDD1.n80 VSUBS 0.038945f
C1460 VDD1.n81 VSUBS 0.017446f
C1461 VDD1.n82 VSUBS 0.030662f
C1462 VDD1.n83 VSUBS 0.016477f
C1463 VDD1.n84 VSUBS 0.038945f
C1464 VDD1.n85 VSUBS 0.017446f
C1465 VDD1.n86 VSUBS 0.030662f
C1466 VDD1.n87 VSUBS 0.016477f
C1467 VDD1.n88 VSUBS 0.038945f
C1468 VDD1.n89 VSUBS 0.017446f
C1469 VDD1.n90 VSUBS 0.030662f
C1470 VDD1.n91 VSUBS 0.016477f
C1471 VDD1.n92 VSUBS 0.038945f
C1472 VDD1.n93 VSUBS 0.017446f
C1473 VDD1.n94 VSUBS 1.71704f
C1474 VDD1.n95 VSUBS 0.016477f
C1475 VDD1.t7 VSUBS 0.083242f
C1476 VDD1.n96 VSUBS 0.200498f
C1477 VDD1.n97 VSUBS 0.024775f
C1478 VDD1.n98 VSUBS 0.029209f
C1479 VDD1.n99 VSUBS 0.038945f
C1480 VDD1.n100 VSUBS 0.017446f
C1481 VDD1.n101 VSUBS 0.016477f
C1482 VDD1.n102 VSUBS 0.030662f
C1483 VDD1.n103 VSUBS 0.030662f
C1484 VDD1.n104 VSUBS 0.016477f
C1485 VDD1.n105 VSUBS 0.017446f
C1486 VDD1.n106 VSUBS 0.038945f
C1487 VDD1.n107 VSUBS 0.038945f
C1488 VDD1.n108 VSUBS 0.017446f
C1489 VDD1.n109 VSUBS 0.016477f
C1490 VDD1.n110 VSUBS 0.030662f
C1491 VDD1.n111 VSUBS 0.030662f
C1492 VDD1.n112 VSUBS 0.016477f
C1493 VDD1.n113 VSUBS 0.017446f
C1494 VDD1.n114 VSUBS 0.038945f
C1495 VDD1.n115 VSUBS 0.038945f
C1496 VDD1.n116 VSUBS 0.017446f
C1497 VDD1.n117 VSUBS 0.016477f
C1498 VDD1.n118 VSUBS 0.030662f
C1499 VDD1.n119 VSUBS 0.030662f
C1500 VDD1.n120 VSUBS 0.016477f
C1501 VDD1.n121 VSUBS 0.017446f
C1502 VDD1.n122 VSUBS 0.038945f
C1503 VDD1.n123 VSUBS 0.038945f
C1504 VDD1.n124 VSUBS 0.017446f
C1505 VDD1.n125 VSUBS 0.016477f
C1506 VDD1.n126 VSUBS 0.030662f
C1507 VDD1.n127 VSUBS 0.030662f
C1508 VDD1.n128 VSUBS 0.016477f
C1509 VDD1.n129 VSUBS 0.017446f
C1510 VDD1.n130 VSUBS 0.038945f
C1511 VDD1.n131 VSUBS 0.038945f
C1512 VDD1.n132 VSUBS 0.017446f
C1513 VDD1.n133 VSUBS 0.016477f
C1514 VDD1.n134 VSUBS 0.030662f
C1515 VDD1.n135 VSUBS 0.030662f
C1516 VDD1.n136 VSUBS 0.016477f
C1517 VDD1.n137 VSUBS 0.017446f
C1518 VDD1.n138 VSUBS 0.038945f
C1519 VDD1.n139 VSUBS 0.094362f
C1520 VDD1.n140 VSUBS 0.017446f
C1521 VDD1.n141 VSUBS 0.032356f
C1522 VDD1.n142 VSUBS 0.073807f
C1523 VDD1.n143 VSUBS 0.118874f
C1524 VDD1.t3 VSUBS 0.321537f
C1525 VDD1.t9 VSUBS 0.321537f
C1526 VDD1.n144 VSUBS 2.56872f
C1527 VDD1.n145 VSUBS 1.38006f
C1528 VDD1.t8 VSUBS 0.321537f
C1529 VDD1.t0 VSUBS 0.321537f
C1530 VDD1.n146 VSUBS 2.60901f
C1531 VDD1.n147 VSUBS 4.89825f
C1532 VDD1.t4 VSUBS 0.321537f
C1533 VDD1.t1 VSUBS 0.321537f
C1534 VDD1.n148 VSUBS 2.56872f
C1535 VDD1.n149 VSUBS 4.91078f
C1536 VTAIL.t4 VSUBS 0.309237f
C1537 VTAIL.t5 VSUBS 0.309237f
C1538 VTAIL.n0 VSUBS 2.31104f
C1539 VTAIL.n1 VSUBS 1.13429f
C1540 VTAIL.n2 VSUBS 0.030516f
C1541 VTAIL.n3 VSUBS 0.029489f
C1542 VTAIL.n4 VSUBS 0.015846f
C1543 VTAIL.n5 VSUBS 0.037455f
C1544 VTAIL.n6 VSUBS 0.016779f
C1545 VTAIL.n7 VSUBS 0.029489f
C1546 VTAIL.n8 VSUBS 0.015846f
C1547 VTAIL.n9 VSUBS 0.037455f
C1548 VTAIL.n10 VSUBS 0.016779f
C1549 VTAIL.n11 VSUBS 0.029489f
C1550 VTAIL.n12 VSUBS 0.015846f
C1551 VTAIL.n13 VSUBS 0.037455f
C1552 VTAIL.n14 VSUBS 0.016779f
C1553 VTAIL.n15 VSUBS 0.029489f
C1554 VTAIL.n16 VSUBS 0.015846f
C1555 VTAIL.n17 VSUBS 0.037455f
C1556 VTAIL.n18 VSUBS 0.016779f
C1557 VTAIL.n19 VSUBS 0.029489f
C1558 VTAIL.n20 VSUBS 0.015846f
C1559 VTAIL.n21 VSUBS 0.037455f
C1560 VTAIL.n22 VSUBS 0.016779f
C1561 VTAIL.n23 VSUBS 1.65136f
C1562 VTAIL.n24 VSUBS 0.015846f
C1563 VTAIL.t16 VSUBS 0.080058f
C1564 VTAIL.n25 VSUBS 0.192828f
C1565 VTAIL.n26 VSUBS 0.023827f
C1566 VTAIL.n27 VSUBS 0.028091f
C1567 VTAIL.n28 VSUBS 0.037455f
C1568 VTAIL.n29 VSUBS 0.016779f
C1569 VTAIL.n30 VSUBS 0.015846f
C1570 VTAIL.n31 VSUBS 0.029489f
C1571 VTAIL.n32 VSUBS 0.029489f
C1572 VTAIL.n33 VSUBS 0.015846f
C1573 VTAIL.n34 VSUBS 0.016779f
C1574 VTAIL.n35 VSUBS 0.037455f
C1575 VTAIL.n36 VSUBS 0.037455f
C1576 VTAIL.n37 VSUBS 0.016779f
C1577 VTAIL.n38 VSUBS 0.015846f
C1578 VTAIL.n39 VSUBS 0.029489f
C1579 VTAIL.n40 VSUBS 0.029489f
C1580 VTAIL.n41 VSUBS 0.015846f
C1581 VTAIL.n42 VSUBS 0.016779f
C1582 VTAIL.n43 VSUBS 0.037455f
C1583 VTAIL.n44 VSUBS 0.037455f
C1584 VTAIL.n45 VSUBS 0.016779f
C1585 VTAIL.n46 VSUBS 0.015846f
C1586 VTAIL.n47 VSUBS 0.029489f
C1587 VTAIL.n48 VSUBS 0.029489f
C1588 VTAIL.n49 VSUBS 0.015846f
C1589 VTAIL.n50 VSUBS 0.016779f
C1590 VTAIL.n51 VSUBS 0.037455f
C1591 VTAIL.n52 VSUBS 0.037455f
C1592 VTAIL.n53 VSUBS 0.016779f
C1593 VTAIL.n54 VSUBS 0.015846f
C1594 VTAIL.n55 VSUBS 0.029489f
C1595 VTAIL.n56 VSUBS 0.029489f
C1596 VTAIL.n57 VSUBS 0.015846f
C1597 VTAIL.n58 VSUBS 0.016779f
C1598 VTAIL.n59 VSUBS 0.037455f
C1599 VTAIL.n60 VSUBS 0.037455f
C1600 VTAIL.n61 VSUBS 0.016779f
C1601 VTAIL.n62 VSUBS 0.015846f
C1602 VTAIL.n63 VSUBS 0.029489f
C1603 VTAIL.n64 VSUBS 0.029489f
C1604 VTAIL.n65 VSUBS 0.015846f
C1605 VTAIL.n66 VSUBS 0.016779f
C1606 VTAIL.n67 VSUBS 0.037455f
C1607 VTAIL.n68 VSUBS 0.090752f
C1608 VTAIL.n69 VSUBS 0.016779f
C1609 VTAIL.n70 VSUBS 0.031118f
C1610 VTAIL.n71 VSUBS 0.070983f
C1611 VTAIL.n72 VSUBS 0.068289f
C1612 VTAIL.n73 VSUBS 0.572743f
C1613 VTAIL.t12 VSUBS 0.309237f
C1614 VTAIL.t14 VSUBS 0.309237f
C1615 VTAIL.n74 VSUBS 2.31104f
C1616 VTAIL.n75 VSUBS 1.33477f
C1617 VTAIL.t15 VSUBS 0.309237f
C1618 VTAIL.t13 VSUBS 0.309237f
C1619 VTAIL.n76 VSUBS 2.31104f
C1620 VTAIL.n77 VSUBS 3.15658f
C1621 VTAIL.t7 VSUBS 0.309237f
C1622 VTAIL.t2 VSUBS 0.309237f
C1623 VTAIL.n78 VSUBS 2.31106f
C1624 VTAIL.n79 VSUBS 3.15656f
C1625 VTAIL.t0 VSUBS 0.309237f
C1626 VTAIL.t9 VSUBS 0.309237f
C1627 VTAIL.n80 VSUBS 2.31106f
C1628 VTAIL.n81 VSUBS 1.33476f
C1629 VTAIL.n82 VSUBS 0.030516f
C1630 VTAIL.n83 VSUBS 0.029489f
C1631 VTAIL.n84 VSUBS 0.015846f
C1632 VTAIL.n85 VSUBS 0.037455f
C1633 VTAIL.n86 VSUBS 0.016779f
C1634 VTAIL.n87 VSUBS 0.029489f
C1635 VTAIL.n88 VSUBS 0.015846f
C1636 VTAIL.n89 VSUBS 0.037455f
C1637 VTAIL.n90 VSUBS 0.016779f
C1638 VTAIL.n91 VSUBS 0.029489f
C1639 VTAIL.n92 VSUBS 0.015846f
C1640 VTAIL.n93 VSUBS 0.037455f
C1641 VTAIL.n94 VSUBS 0.016779f
C1642 VTAIL.n95 VSUBS 0.029489f
C1643 VTAIL.n96 VSUBS 0.015846f
C1644 VTAIL.n97 VSUBS 0.037455f
C1645 VTAIL.n98 VSUBS 0.016779f
C1646 VTAIL.n99 VSUBS 0.029489f
C1647 VTAIL.n100 VSUBS 0.015846f
C1648 VTAIL.n101 VSUBS 0.037455f
C1649 VTAIL.n102 VSUBS 0.016779f
C1650 VTAIL.n103 VSUBS 1.65136f
C1651 VTAIL.n104 VSUBS 0.015846f
C1652 VTAIL.t6 VSUBS 0.080058f
C1653 VTAIL.n105 VSUBS 0.192828f
C1654 VTAIL.n106 VSUBS 0.023827f
C1655 VTAIL.n107 VSUBS 0.028091f
C1656 VTAIL.n108 VSUBS 0.037455f
C1657 VTAIL.n109 VSUBS 0.016779f
C1658 VTAIL.n110 VSUBS 0.015846f
C1659 VTAIL.n111 VSUBS 0.029489f
C1660 VTAIL.n112 VSUBS 0.029489f
C1661 VTAIL.n113 VSUBS 0.015846f
C1662 VTAIL.n114 VSUBS 0.016779f
C1663 VTAIL.n115 VSUBS 0.037455f
C1664 VTAIL.n116 VSUBS 0.037455f
C1665 VTAIL.n117 VSUBS 0.016779f
C1666 VTAIL.n118 VSUBS 0.015846f
C1667 VTAIL.n119 VSUBS 0.029489f
C1668 VTAIL.n120 VSUBS 0.029489f
C1669 VTAIL.n121 VSUBS 0.015846f
C1670 VTAIL.n122 VSUBS 0.016779f
C1671 VTAIL.n123 VSUBS 0.037455f
C1672 VTAIL.n124 VSUBS 0.037455f
C1673 VTAIL.n125 VSUBS 0.016779f
C1674 VTAIL.n126 VSUBS 0.015846f
C1675 VTAIL.n127 VSUBS 0.029489f
C1676 VTAIL.n128 VSUBS 0.029489f
C1677 VTAIL.n129 VSUBS 0.015846f
C1678 VTAIL.n130 VSUBS 0.016779f
C1679 VTAIL.n131 VSUBS 0.037455f
C1680 VTAIL.n132 VSUBS 0.037455f
C1681 VTAIL.n133 VSUBS 0.016779f
C1682 VTAIL.n134 VSUBS 0.015846f
C1683 VTAIL.n135 VSUBS 0.029489f
C1684 VTAIL.n136 VSUBS 0.029489f
C1685 VTAIL.n137 VSUBS 0.015846f
C1686 VTAIL.n138 VSUBS 0.016779f
C1687 VTAIL.n139 VSUBS 0.037455f
C1688 VTAIL.n140 VSUBS 0.037455f
C1689 VTAIL.n141 VSUBS 0.016779f
C1690 VTAIL.n142 VSUBS 0.015846f
C1691 VTAIL.n143 VSUBS 0.029489f
C1692 VTAIL.n144 VSUBS 0.029489f
C1693 VTAIL.n145 VSUBS 0.015846f
C1694 VTAIL.n146 VSUBS 0.016779f
C1695 VTAIL.n147 VSUBS 0.037455f
C1696 VTAIL.n148 VSUBS 0.090752f
C1697 VTAIL.n149 VSUBS 0.016779f
C1698 VTAIL.n150 VSUBS 0.031118f
C1699 VTAIL.n151 VSUBS 0.070983f
C1700 VTAIL.n152 VSUBS 0.068289f
C1701 VTAIL.n153 VSUBS 0.572743f
C1702 VTAIL.t10 VSUBS 0.309237f
C1703 VTAIL.t18 VSUBS 0.309237f
C1704 VTAIL.n154 VSUBS 2.31106f
C1705 VTAIL.n155 VSUBS 1.21229f
C1706 VTAIL.t17 VSUBS 0.309237f
C1707 VTAIL.t11 VSUBS 0.309237f
C1708 VTAIL.n156 VSUBS 2.31106f
C1709 VTAIL.n157 VSUBS 1.33476f
C1710 VTAIL.n158 VSUBS 0.030516f
C1711 VTAIL.n159 VSUBS 0.029489f
C1712 VTAIL.n160 VSUBS 0.015846f
C1713 VTAIL.n161 VSUBS 0.037455f
C1714 VTAIL.n162 VSUBS 0.016779f
C1715 VTAIL.n163 VSUBS 0.029489f
C1716 VTAIL.n164 VSUBS 0.015846f
C1717 VTAIL.n165 VSUBS 0.037455f
C1718 VTAIL.n166 VSUBS 0.016779f
C1719 VTAIL.n167 VSUBS 0.029489f
C1720 VTAIL.n168 VSUBS 0.015846f
C1721 VTAIL.n169 VSUBS 0.037455f
C1722 VTAIL.n170 VSUBS 0.016779f
C1723 VTAIL.n171 VSUBS 0.029489f
C1724 VTAIL.n172 VSUBS 0.015846f
C1725 VTAIL.n173 VSUBS 0.037455f
C1726 VTAIL.n174 VSUBS 0.016779f
C1727 VTAIL.n175 VSUBS 0.029489f
C1728 VTAIL.n176 VSUBS 0.015846f
C1729 VTAIL.n177 VSUBS 0.037455f
C1730 VTAIL.n178 VSUBS 0.016779f
C1731 VTAIL.n179 VSUBS 1.65136f
C1732 VTAIL.n180 VSUBS 0.015846f
C1733 VTAIL.t19 VSUBS 0.080058f
C1734 VTAIL.n181 VSUBS 0.192828f
C1735 VTAIL.n182 VSUBS 0.023827f
C1736 VTAIL.n183 VSUBS 0.028091f
C1737 VTAIL.n184 VSUBS 0.037455f
C1738 VTAIL.n185 VSUBS 0.016779f
C1739 VTAIL.n186 VSUBS 0.015846f
C1740 VTAIL.n187 VSUBS 0.029489f
C1741 VTAIL.n188 VSUBS 0.029489f
C1742 VTAIL.n189 VSUBS 0.015846f
C1743 VTAIL.n190 VSUBS 0.016779f
C1744 VTAIL.n191 VSUBS 0.037455f
C1745 VTAIL.n192 VSUBS 0.037455f
C1746 VTAIL.n193 VSUBS 0.016779f
C1747 VTAIL.n194 VSUBS 0.015846f
C1748 VTAIL.n195 VSUBS 0.029489f
C1749 VTAIL.n196 VSUBS 0.029489f
C1750 VTAIL.n197 VSUBS 0.015846f
C1751 VTAIL.n198 VSUBS 0.016779f
C1752 VTAIL.n199 VSUBS 0.037455f
C1753 VTAIL.n200 VSUBS 0.037455f
C1754 VTAIL.n201 VSUBS 0.016779f
C1755 VTAIL.n202 VSUBS 0.015846f
C1756 VTAIL.n203 VSUBS 0.029489f
C1757 VTAIL.n204 VSUBS 0.029489f
C1758 VTAIL.n205 VSUBS 0.015846f
C1759 VTAIL.n206 VSUBS 0.016779f
C1760 VTAIL.n207 VSUBS 0.037455f
C1761 VTAIL.n208 VSUBS 0.037455f
C1762 VTAIL.n209 VSUBS 0.016779f
C1763 VTAIL.n210 VSUBS 0.015846f
C1764 VTAIL.n211 VSUBS 0.029489f
C1765 VTAIL.n212 VSUBS 0.029489f
C1766 VTAIL.n213 VSUBS 0.015846f
C1767 VTAIL.n214 VSUBS 0.016779f
C1768 VTAIL.n215 VSUBS 0.037455f
C1769 VTAIL.n216 VSUBS 0.037455f
C1770 VTAIL.n217 VSUBS 0.016779f
C1771 VTAIL.n218 VSUBS 0.015846f
C1772 VTAIL.n219 VSUBS 0.029489f
C1773 VTAIL.n220 VSUBS 0.029489f
C1774 VTAIL.n221 VSUBS 0.015846f
C1775 VTAIL.n222 VSUBS 0.016779f
C1776 VTAIL.n223 VSUBS 0.037455f
C1777 VTAIL.n224 VSUBS 0.090752f
C1778 VTAIL.n225 VSUBS 0.016779f
C1779 VTAIL.n226 VSUBS 0.031118f
C1780 VTAIL.n227 VSUBS 0.070983f
C1781 VTAIL.n228 VSUBS 0.068289f
C1782 VTAIL.n229 VSUBS 2.1828f
C1783 VTAIL.n230 VSUBS 0.030516f
C1784 VTAIL.n231 VSUBS 0.029489f
C1785 VTAIL.n232 VSUBS 0.015846f
C1786 VTAIL.n233 VSUBS 0.037455f
C1787 VTAIL.n234 VSUBS 0.016779f
C1788 VTAIL.n235 VSUBS 0.029489f
C1789 VTAIL.n236 VSUBS 0.015846f
C1790 VTAIL.n237 VSUBS 0.037455f
C1791 VTAIL.n238 VSUBS 0.016779f
C1792 VTAIL.n239 VSUBS 0.029489f
C1793 VTAIL.n240 VSUBS 0.015846f
C1794 VTAIL.n241 VSUBS 0.037455f
C1795 VTAIL.n242 VSUBS 0.016779f
C1796 VTAIL.n243 VSUBS 0.029489f
C1797 VTAIL.n244 VSUBS 0.015846f
C1798 VTAIL.n245 VSUBS 0.037455f
C1799 VTAIL.n246 VSUBS 0.016779f
C1800 VTAIL.n247 VSUBS 0.029489f
C1801 VTAIL.n248 VSUBS 0.015846f
C1802 VTAIL.n249 VSUBS 0.037455f
C1803 VTAIL.n250 VSUBS 0.016779f
C1804 VTAIL.n251 VSUBS 1.65136f
C1805 VTAIL.n252 VSUBS 0.015846f
C1806 VTAIL.t1 VSUBS 0.080058f
C1807 VTAIL.n253 VSUBS 0.192828f
C1808 VTAIL.n254 VSUBS 0.023827f
C1809 VTAIL.n255 VSUBS 0.028091f
C1810 VTAIL.n256 VSUBS 0.037455f
C1811 VTAIL.n257 VSUBS 0.016779f
C1812 VTAIL.n258 VSUBS 0.015846f
C1813 VTAIL.n259 VSUBS 0.029489f
C1814 VTAIL.n260 VSUBS 0.029489f
C1815 VTAIL.n261 VSUBS 0.015846f
C1816 VTAIL.n262 VSUBS 0.016779f
C1817 VTAIL.n263 VSUBS 0.037455f
C1818 VTAIL.n264 VSUBS 0.037455f
C1819 VTAIL.n265 VSUBS 0.016779f
C1820 VTAIL.n266 VSUBS 0.015846f
C1821 VTAIL.n267 VSUBS 0.029489f
C1822 VTAIL.n268 VSUBS 0.029489f
C1823 VTAIL.n269 VSUBS 0.015846f
C1824 VTAIL.n270 VSUBS 0.016779f
C1825 VTAIL.n271 VSUBS 0.037455f
C1826 VTAIL.n272 VSUBS 0.037455f
C1827 VTAIL.n273 VSUBS 0.016779f
C1828 VTAIL.n274 VSUBS 0.015846f
C1829 VTAIL.n275 VSUBS 0.029489f
C1830 VTAIL.n276 VSUBS 0.029489f
C1831 VTAIL.n277 VSUBS 0.015846f
C1832 VTAIL.n278 VSUBS 0.016779f
C1833 VTAIL.n279 VSUBS 0.037455f
C1834 VTAIL.n280 VSUBS 0.037455f
C1835 VTAIL.n281 VSUBS 0.016779f
C1836 VTAIL.n282 VSUBS 0.015846f
C1837 VTAIL.n283 VSUBS 0.029489f
C1838 VTAIL.n284 VSUBS 0.029489f
C1839 VTAIL.n285 VSUBS 0.015846f
C1840 VTAIL.n286 VSUBS 0.016779f
C1841 VTAIL.n287 VSUBS 0.037455f
C1842 VTAIL.n288 VSUBS 0.037455f
C1843 VTAIL.n289 VSUBS 0.016779f
C1844 VTAIL.n290 VSUBS 0.015846f
C1845 VTAIL.n291 VSUBS 0.029489f
C1846 VTAIL.n292 VSUBS 0.029489f
C1847 VTAIL.n293 VSUBS 0.015846f
C1848 VTAIL.n294 VSUBS 0.016779f
C1849 VTAIL.n295 VSUBS 0.037455f
C1850 VTAIL.n296 VSUBS 0.090752f
C1851 VTAIL.n297 VSUBS 0.016779f
C1852 VTAIL.n298 VSUBS 0.031118f
C1853 VTAIL.n299 VSUBS 0.070983f
C1854 VTAIL.n300 VSUBS 0.068289f
C1855 VTAIL.n301 VSUBS 2.1828f
C1856 VTAIL.t8 VSUBS 0.309237f
C1857 VTAIL.t3 VSUBS 0.309237f
C1858 VTAIL.n302 VSUBS 2.31104f
C1859 VTAIL.n303 VSUBS 1.07858f
C1860 VP.t9 VSUBS 3.33315f
C1861 VP.n0 VSUBS 1.25986f
C1862 VP.n1 VSUBS 0.024517f
C1863 VP.n2 VSUBS 0.044014f
C1864 VP.n3 VSUBS 0.024517f
C1865 VP.n4 VSUBS 0.042083f
C1866 VP.n5 VSUBS 0.024517f
C1867 VP.n6 VSUBS 0.047513f
C1868 VP.n7 VSUBS 0.024517f
C1869 VP.n8 VSUBS 0.045693f
C1870 VP.n9 VSUBS 0.024517f
C1871 VP.t0 VSUBS 3.33315f
C1872 VP.n10 VSUBS 0.049432f
C1873 VP.n11 VSUBS 0.024517f
C1874 VP.n12 VSUBS 0.045693f
C1875 VP.n13 VSUBS 0.024517f
C1876 VP.t6 VSUBS 3.33315f
C1877 VP.n14 VSUBS 0.048495f
C1878 VP.n15 VSUBS 0.024517f
C1879 VP.n16 VSUBS 0.045693f
C1880 VP.t8 VSUBS 3.33315f
C1881 VP.n17 VSUBS 1.25986f
C1882 VP.n18 VSUBS 0.024517f
C1883 VP.n19 VSUBS 0.044014f
C1884 VP.n20 VSUBS 0.024517f
C1885 VP.n21 VSUBS 0.042083f
C1886 VP.n22 VSUBS 0.024517f
C1887 VP.n23 VSUBS 0.047513f
C1888 VP.n24 VSUBS 0.024517f
C1889 VP.n25 VSUBS 0.045693f
C1890 VP.n26 VSUBS 0.024517f
C1891 VP.t4 VSUBS 3.33315f
C1892 VP.n27 VSUBS 0.049432f
C1893 VP.n28 VSUBS 0.024517f
C1894 VP.n29 VSUBS 0.045693f
C1895 VP.t7 VSUBS 3.71048f
C1896 VP.n30 VSUBS 1.17882f
C1897 VP.t3 VSUBS 3.33315f
C1898 VP.n31 VSUBS 1.24217f
C1899 VP.n32 VSUBS 0.026743f
C1900 VP.n33 VSUBS 0.311334f
C1901 VP.n34 VSUBS 0.024517f
C1902 VP.n35 VSUBS 0.024517f
C1903 VP.n36 VSUBS 0.045693f
C1904 VP.n37 VSUBS 0.047513f
C1905 VP.n38 VSUBS 0.020328f
C1906 VP.n39 VSUBS 0.024517f
C1907 VP.n40 VSUBS 0.024517f
C1908 VP.n41 VSUBS 0.024517f
C1909 VP.n42 VSUBS 0.045693f
C1910 VP.n43 VSUBS 0.045693f
C1911 VP.n44 VSUBS 1.18537f
C1912 VP.n45 VSUBS 0.024517f
C1913 VP.n46 VSUBS 0.024517f
C1914 VP.n47 VSUBS 0.024517f
C1915 VP.n48 VSUBS 0.045693f
C1916 VP.n49 VSUBS 0.049432f
C1917 VP.n50 VSUBS 0.020328f
C1918 VP.n51 VSUBS 0.024517f
C1919 VP.n52 VSUBS 0.024517f
C1920 VP.n53 VSUBS 0.024517f
C1921 VP.n54 VSUBS 0.045693f
C1922 VP.n55 VSUBS 0.045693f
C1923 VP.t5 VSUBS 3.33315f
C1924 VP.n56 VSUBS 1.16224f
C1925 VP.n57 VSUBS 0.026743f
C1926 VP.n58 VSUBS 0.024517f
C1927 VP.n59 VSUBS 0.024517f
C1928 VP.n60 VSUBS 0.024517f
C1929 VP.n61 VSUBS 0.045693f
C1930 VP.n62 VSUBS 0.048495f
C1931 VP.n63 VSUBS 0.024763f
C1932 VP.n64 VSUBS 0.024517f
C1933 VP.n65 VSUBS 0.024517f
C1934 VP.n66 VSUBS 0.024517f
C1935 VP.n67 VSUBS 0.045693f
C1936 VP.n68 VSUBS 0.045693f
C1937 VP.n69 VSUBS 0.030353f
C1938 VP.n70 VSUBS 0.039569f
C1939 VP.n71 VSUBS 1.82602f
C1940 VP.n72 VSUBS 1.8406f
C1941 VP.t2 VSUBS 3.33315f
C1942 VP.n73 VSUBS 1.25986f
C1943 VP.n74 VSUBS 0.030353f
C1944 VP.n75 VSUBS 0.039569f
C1945 VP.n76 VSUBS 0.024517f
C1946 VP.n77 VSUBS 0.024517f
C1947 VP.n78 VSUBS 0.045693f
C1948 VP.n79 VSUBS 0.044014f
C1949 VP.n80 VSUBS 0.024763f
C1950 VP.n81 VSUBS 0.024517f
C1951 VP.n82 VSUBS 0.024517f
C1952 VP.n83 VSUBS 0.024517f
C1953 VP.n84 VSUBS 0.045693f
C1954 VP.n85 VSUBS 0.042083f
C1955 VP.n86 VSUBS 1.16224f
C1956 VP.n87 VSUBS 0.026743f
C1957 VP.n88 VSUBS 0.024517f
C1958 VP.n89 VSUBS 0.024517f
C1959 VP.n90 VSUBS 0.024517f
C1960 VP.n91 VSUBS 0.045693f
C1961 VP.n92 VSUBS 0.047513f
C1962 VP.n93 VSUBS 0.020328f
C1963 VP.n94 VSUBS 0.024517f
C1964 VP.n95 VSUBS 0.024517f
C1965 VP.n96 VSUBS 0.024517f
C1966 VP.n97 VSUBS 0.045693f
C1967 VP.n98 VSUBS 0.045693f
C1968 VP.n99 VSUBS 1.18537f
C1969 VP.n100 VSUBS 0.024517f
C1970 VP.n101 VSUBS 0.024517f
C1971 VP.n102 VSUBS 0.024517f
C1972 VP.n103 VSUBS 0.045693f
C1973 VP.n104 VSUBS 0.049432f
C1974 VP.n105 VSUBS 0.020328f
C1975 VP.n106 VSUBS 0.024517f
C1976 VP.n107 VSUBS 0.024517f
C1977 VP.n108 VSUBS 0.024517f
C1978 VP.n109 VSUBS 0.045693f
C1979 VP.n110 VSUBS 0.045693f
C1980 VP.t1 VSUBS 3.33315f
C1981 VP.n111 VSUBS 1.16224f
C1982 VP.n112 VSUBS 0.026743f
C1983 VP.n113 VSUBS 0.024517f
C1984 VP.n114 VSUBS 0.024517f
C1985 VP.n115 VSUBS 0.024517f
C1986 VP.n116 VSUBS 0.045693f
C1987 VP.n117 VSUBS 0.048495f
C1988 VP.n118 VSUBS 0.024763f
C1989 VP.n119 VSUBS 0.024517f
C1990 VP.n120 VSUBS 0.024517f
C1991 VP.n121 VSUBS 0.024517f
C1992 VP.n122 VSUBS 0.045693f
C1993 VP.n123 VSUBS 0.045693f
C1994 VP.n124 VSUBS 0.030353f
C1995 VP.n125 VSUBS 0.039569f
C1996 VP.n126 VSUBS 0.070729f
.ends

