* NGSPICE file created from diff_pair_sample_1491.ext - technology: sky130A

.subckt diff_pair_sample_1491 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0 ps=0 w=3.46 l=3.71
X1 VDD1.t5 VP.t0 VTAIL.t6 B.t19 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=1.3494 ps=7.7 w=3.46 l=3.71
X2 VDD2.t5 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0.5709 ps=3.79 w=3.46 l=3.71
X3 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0 ps=0 w=3.46 l=3.71
X4 VDD1.t4 VP.t1 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0.5709 ps=3.79 w=3.46 l=3.71
X5 VDD1.t3 VP.t2 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=1.3494 ps=7.7 w=3.46 l=3.71
X6 VDD2.t4 VN.t1 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=1.3494 ps=7.7 w=3.46 l=3.71
X7 VTAIL.t0 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=0.5709 ps=3.79 w=3.46 l=3.71
X8 VDD2.t2 VN.t3 VTAIL.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=1.3494 ps=7.7 w=3.46 l=3.71
X9 VTAIL.t10 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=0.5709 ps=3.79 w=3.46 l=3.71
X10 VTAIL.t9 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=0.5709 ps=3.79 w=3.46 l=3.71
X11 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0.5709 ps=3.79 w=3.46 l=3.71
X12 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5709 pd=3.79 as=0.5709 ps=3.79 w=3.46 l=3.71
X13 VDD1.t0 VP.t5 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0.5709 ps=3.79 w=3.46 l=3.71
X14 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0 ps=0 w=3.46 l=3.71
X15 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3494 pd=7.7 as=0 ps=0 w=3.46 l=3.71
R0 B.n669 B.n668 585
R1 B.n670 B.n669 585
R2 B.n210 B.n124 585
R3 B.n209 B.n208 585
R4 B.n207 B.n206 585
R5 B.n205 B.n204 585
R6 B.n203 B.n202 585
R7 B.n201 B.n200 585
R8 B.n199 B.n198 585
R9 B.n197 B.n196 585
R10 B.n195 B.n194 585
R11 B.n193 B.n192 585
R12 B.n191 B.n190 585
R13 B.n189 B.n188 585
R14 B.n187 B.n186 585
R15 B.n185 B.n184 585
R16 B.n183 B.n182 585
R17 B.n181 B.n180 585
R18 B.n179 B.n178 585
R19 B.n177 B.n176 585
R20 B.n175 B.n174 585
R21 B.n173 B.n172 585
R22 B.n171 B.n170 585
R23 B.n169 B.n168 585
R24 B.n167 B.n166 585
R25 B.n165 B.n164 585
R26 B.n163 B.n162 585
R27 B.n160 B.n159 585
R28 B.n158 B.n157 585
R29 B.n156 B.n155 585
R30 B.n154 B.n153 585
R31 B.n152 B.n151 585
R32 B.n150 B.n149 585
R33 B.n148 B.n147 585
R34 B.n146 B.n145 585
R35 B.n144 B.n143 585
R36 B.n142 B.n141 585
R37 B.n140 B.n139 585
R38 B.n138 B.n137 585
R39 B.n136 B.n135 585
R40 B.n134 B.n133 585
R41 B.n132 B.n131 585
R42 B.n103 B.n102 585
R43 B.n673 B.n672 585
R44 B.n667 B.n125 585
R45 B.n125 B.n100 585
R46 B.n666 B.n99 585
R47 B.n677 B.n99 585
R48 B.n665 B.n98 585
R49 B.n678 B.n98 585
R50 B.n664 B.n97 585
R51 B.n679 B.n97 585
R52 B.n663 B.n662 585
R53 B.n662 B.n93 585
R54 B.n661 B.n92 585
R55 B.n685 B.n92 585
R56 B.n660 B.n91 585
R57 B.n686 B.n91 585
R58 B.n659 B.n90 585
R59 B.n687 B.n90 585
R60 B.n658 B.n657 585
R61 B.n657 B.n86 585
R62 B.n656 B.n85 585
R63 B.n693 B.n85 585
R64 B.n655 B.n84 585
R65 B.n694 B.n84 585
R66 B.n654 B.n83 585
R67 B.n695 B.n83 585
R68 B.n653 B.n652 585
R69 B.n652 B.n79 585
R70 B.n651 B.n78 585
R71 B.n701 B.n78 585
R72 B.n650 B.n77 585
R73 B.n702 B.n77 585
R74 B.n649 B.n76 585
R75 B.n703 B.n76 585
R76 B.n648 B.n647 585
R77 B.n647 B.n72 585
R78 B.n646 B.n71 585
R79 B.n709 B.n71 585
R80 B.n645 B.n70 585
R81 B.n710 B.n70 585
R82 B.n644 B.n69 585
R83 B.n711 B.n69 585
R84 B.n643 B.n642 585
R85 B.n642 B.n65 585
R86 B.n641 B.n64 585
R87 B.n717 B.n64 585
R88 B.n640 B.n63 585
R89 B.n718 B.n63 585
R90 B.n639 B.n62 585
R91 B.n719 B.n62 585
R92 B.n638 B.n637 585
R93 B.n637 B.n61 585
R94 B.n636 B.n57 585
R95 B.n725 B.n57 585
R96 B.n635 B.n56 585
R97 B.n726 B.n56 585
R98 B.n634 B.n55 585
R99 B.n727 B.n55 585
R100 B.n633 B.n632 585
R101 B.n632 B.n51 585
R102 B.n631 B.n50 585
R103 B.n733 B.n50 585
R104 B.n630 B.n49 585
R105 B.n734 B.n49 585
R106 B.n629 B.n48 585
R107 B.n735 B.n48 585
R108 B.n628 B.n627 585
R109 B.n627 B.n44 585
R110 B.n626 B.n43 585
R111 B.n741 B.n43 585
R112 B.n625 B.n42 585
R113 B.n742 B.n42 585
R114 B.n624 B.n41 585
R115 B.n743 B.n41 585
R116 B.n623 B.n622 585
R117 B.n622 B.n40 585
R118 B.n621 B.n36 585
R119 B.n749 B.n36 585
R120 B.n620 B.n35 585
R121 B.n750 B.n35 585
R122 B.n619 B.n34 585
R123 B.n751 B.n34 585
R124 B.n618 B.n617 585
R125 B.n617 B.n30 585
R126 B.n616 B.n29 585
R127 B.n757 B.n29 585
R128 B.n615 B.n28 585
R129 B.n758 B.n28 585
R130 B.n614 B.n27 585
R131 B.n759 B.n27 585
R132 B.n613 B.n612 585
R133 B.n612 B.n23 585
R134 B.n611 B.n22 585
R135 B.n765 B.n22 585
R136 B.n610 B.n21 585
R137 B.n766 B.n21 585
R138 B.n609 B.n20 585
R139 B.n767 B.n20 585
R140 B.n608 B.n607 585
R141 B.n607 B.n16 585
R142 B.n606 B.n15 585
R143 B.n773 B.n15 585
R144 B.n605 B.n14 585
R145 B.n774 B.n14 585
R146 B.n604 B.n13 585
R147 B.n775 B.n13 585
R148 B.n603 B.n602 585
R149 B.n602 B.n12 585
R150 B.n601 B.n600 585
R151 B.n601 B.n8 585
R152 B.n599 B.n7 585
R153 B.n782 B.n7 585
R154 B.n598 B.n6 585
R155 B.n783 B.n6 585
R156 B.n597 B.n5 585
R157 B.n784 B.n5 585
R158 B.n596 B.n595 585
R159 B.n595 B.n4 585
R160 B.n594 B.n211 585
R161 B.n594 B.n593 585
R162 B.n584 B.n212 585
R163 B.n213 B.n212 585
R164 B.n586 B.n585 585
R165 B.n587 B.n586 585
R166 B.n583 B.n218 585
R167 B.n218 B.n217 585
R168 B.n582 B.n581 585
R169 B.n581 B.n580 585
R170 B.n220 B.n219 585
R171 B.n221 B.n220 585
R172 B.n573 B.n572 585
R173 B.n574 B.n573 585
R174 B.n571 B.n226 585
R175 B.n226 B.n225 585
R176 B.n570 B.n569 585
R177 B.n569 B.n568 585
R178 B.n228 B.n227 585
R179 B.n229 B.n228 585
R180 B.n561 B.n560 585
R181 B.n562 B.n561 585
R182 B.n559 B.n234 585
R183 B.n234 B.n233 585
R184 B.n558 B.n557 585
R185 B.n557 B.n556 585
R186 B.n236 B.n235 585
R187 B.n237 B.n236 585
R188 B.n549 B.n548 585
R189 B.n550 B.n549 585
R190 B.n547 B.n242 585
R191 B.n242 B.n241 585
R192 B.n546 B.n545 585
R193 B.n545 B.n544 585
R194 B.n244 B.n243 585
R195 B.n537 B.n244 585
R196 B.n536 B.n535 585
R197 B.n538 B.n536 585
R198 B.n534 B.n249 585
R199 B.n249 B.n248 585
R200 B.n533 B.n532 585
R201 B.n532 B.n531 585
R202 B.n251 B.n250 585
R203 B.n252 B.n251 585
R204 B.n524 B.n523 585
R205 B.n525 B.n524 585
R206 B.n522 B.n257 585
R207 B.n257 B.n256 585
R208 B.n521 B.n520 585
R209 B.n520 B.n519 585
R210 B.n259 B.n258 585
R211 B.n260 B.n259 585
R212 B.n512 B.n511 585
R213 B.n513 B.n512 585
R214 B.n510 B.n265 585
R215 B.n265 B.n264 585
R216 B.n509 B.n508 585
R217 B.n508 B.n507 585
R218 B.n267 B.n266 585
R219 B.n500 B.n267 585
R220 B.n499 B.n498 585
R221 B.n501 B.n499 585
R222 B.n497 B.n272 585
R223 B.n272 B.n271 585
R224 B.n496 B.n495 585
R225 B.n495 B.n494 585
R226 B.n274 B.n273 585
R227 B.n275 B.n274 585
R228 B.n487 B.n486 585
R229 B.n488 B.n487 585
R230 B.n485 B.n280 585
R231 B.n280 B.n279 585
R232 B.n484 B.n483 585
R233 B.n483 B.n482 585
R234 B.n282 B.n281 585
R235 B.n283 B.n282 585
R236 B.n475 B.n474 585
R237 B.n476 B.n475 585
R238 B.n473 B.n288 585
R239 B.n288 B.n287 585
R240 B.n472 B.n471 585
R241 B.n471 B.n470 585
R242 B.n290 B.n289 585
R243 B.n291 B.n290 585
R244 B.n463 B.n462 585
R245 B.n464 B.n463 585
R246 B.n461 B.n296 585
R247 B.n296 B.n295 585
R248 B.n460 B.n459 585
R249 B.n459 B.n458 585
R250 B.n298 B.n297 585
R251 B.n299 B.n298 585
R252 B.n451 B.n450 585
R253 B.n452 B.n451 585
R254 B.n449 B.n304 585
R255 B.n304 B.n303 585
R256 B.n448 B.n447 585
R257 B.n447 B.n446 585
R258 B.n306 B.n305 585
R259 B.n307 B.n306 585
R260 B.n439 B.n438 585
R261 B.n440 B.n439 585
R262 B.n437 B.n312 585
R263 B.n312 B.n311 585
R264 B.n436 B.n435 585
R265 B.n435 B.n434 585
R266 B.n314 B.n313 585
R267 B.n315 B.n314 585
R268 B.n430 B.n429 585
R269 B.n318 B.n317 585
R270 B.n426 B.n425 585
R271 B.n427 B.n426 585
R272 B.n424 B.n339 585
R273 B.n423 B.n422 585
R274 B.n421 B.n420 585
R275 B.n419 B.n418 585
R276 B.n417 B.n416 585
R277 B.n415 B.n414 585
R278 B.n413 B.n412 585
R279 B.n411 B.n410 585
R280 B.n409 B.n408 585
R281 B.n407 B.n406 585
R282 B.n405 B.n404 585
R283 B.n403 B.n402 585
R284 B.n401 B.n400 585
R285 B.n399 B.n398 585
R286 B.n397 B.n396 585
R287 B.n395 B.n394 585
R288 B.n393 B.n392 585
R289 B.n391 B.n390 585
R290 B.n389 B.n388 585
R291 B.n387 B.n386 585
R292 B.n385 B.n384 585
R293 B.n383 B.n382 585
R294 B.n381 B.n380 585
R295 B.n378 B.n377 585
R296 B.n376 B.n375 585
R297 B.n374 B.n373 585
R298 B.n372 B.n371 585
R299 B.n370 B.n369 585
R300 B.n368 B.n367 585
R301 B.n366 B.n365 585
R302 B.n364 B.n363 585
R303 B.n362 B.n361 585
R304 B.n360 B.n359 585
R305 B.n358 B.n357 585
R306 B.n356 B.n355 585
R307 B.n354 B.n353 585
R308 B.n352 B.n351 585
R309 B.n350 B.n349 585
R310 B.n348 B.n347 585
R311 B.n346 B.n345 585
R312 B.n431 B.n316 585
R313 B.n316 B.n315 585
R314 B.n433 B.n432 585
R315 B.n434 B.n433 585
R316 B.n310 B.n309 585
R317 B.n311 B.n310 585
R318 B.n442 B.n441 585
R319 B.n441 B.n440 585
R320 B.n443 B.n308 585
R321 B.n308 B.n307 585
R322 B.n445 B.n444 585
R323 B.n446 B.n445 585
R324 B.n302 B.n301 585
R325 B.n303 B.n302 585
R326 B.n454 B.n453 585
R327 B.n453 B.n452 585
R328 B.n455 B.n300 585
R329 B.n300 B.n299 585
R330 B.n457 B.n456 585
R331 B.n458 B.n457 585
R332 B.n294 B.n293 585
R333 B.n295 B.n294 585
R334 B.n466 B.n465 585
R335 B.n465 B.n464 585
R336 B.n467 B.n292 585
R337 B.n292 B.n291 585
R338 B.n469 B.n468 585
R339 B.n470 B.n469 585
R340 B.n286 B.n285 585
R341 B.n287 B.n286 585
R342 B.n478 B.n477 585
R343 B.n477 B.n476 585
R344 B.n479 B.n284 585
R345 B.n284 B.n283 585
R346 B.n481 B.n480 585
R347 B.n482 B.n481 585
R348 B.n278 B.n277 585
R349 B.n279 B.n278 585
R350 B.n490 B.n489 585
R351 B.n489 B.n488 585
R352 B.n491 B.n276 585
R353 B.n276 B.n275 585
R354 B.n493 B.n492 585
R355 B.n494 B.n493 585
R356 B.n270 B.n269 585
R357 B.n271 B.n270 585
R358 B.n503 B.n502 585
R359 B.n502 B.n501 585
R360 B.n504 B.n268 585
R361 B.n500 B.n268 585
R362 B.n506 B.n505 585
R363 B.n507 B.n506 585
R364 B.n263 B.n262 585
R365 B.n264 B.n263 585
R366 B.n515 B.n514 585
R367 B.n514 B.n513 585
R368 B.n516 B.n261 585
R369 B.n261 B.n260 585
R370 B.n518 B.n517 585
R371 B.n519 B.n518 585
R372 B.n255 B.n254 585
R373 B.n256 B.n255 585
R374 B.n527 B.n526 585
R375 B.n526 B.n525 585
R376 B.n528 B.n253 585
R377 B.n253 B.n252 585
R378 B.n530 B.n529 585
R379 B.n531 B.n530 585
R380 B.n247 B.n246 585
R381 B.n248 B.n247 585
R382 B.n540 B.n539 585
R383 B.n539 B.n538 585
R384 B.n541 B.n245 585
R385 B.n537 B.n245 585
R386 B.n543 B.n542 585
R387 B.n544 B.n543 585
R388 B.n240 B.n239 585
R389 B.n241 B.n240 585
R390 B.n552 B.n551 585
R391 B.n551 B.n550 585
R392 B.n553 B.n238 585
R393 B.n238 B.n237 585
R394 B.n555 B.n554 585
R395 B.n556 B.n555 585
R396 B.n232 B.n231 585
R397 B.n233 B.n232 585
R398 B.n564 B.n563 585
R399 B.n563 B.n562 585
R400 B.n565 B.n230 585
R401 B.n230 B.n229 585
R402 B.n567 B.n566 585
R403 B.n568 B.n567 585
R404 B.n224 B.n223 585
R405 B.n225 B.n224 585
R406 B.n576 B.n575 585
R407 B.n575 B.n574 585
R408 B.n577 B.n222 585
R409 B.n222 B.n221 585
R410 B.n579 B.n578 585
R411 B.n580 B.n579 585
R412 B.n216 B.n215 585
R413 B.n217 B.n216 585
R414 B.n589 B.n588 585
R415 B.n588 B.n587 585
R416 B.n590 B.n214 585
R417 B.n214 B.n213 585
R418 B.n592 B.n591 585
R419 B.n593 B.n592 585
R420 B.n3 B.n0 585
R421 B.n4 B.n3 585
R422 B.n781 B.n1 585
R423 B.n782 B.n781 585
R424 B.n780 B.n779 585
R425 B.n780 B.n8 585
R426 B.n778 B.n9 585
R427 B.n12 B.n9 585
R428 B.n777 B.n776 585
R429 B.n776 B.n775 585
R430 B.n11 B.n10 585
R431 B.n774 B.n11 585
R432 B.n772 B.n771 585
R433 B.n773 B.n772 585
R434 B.n770 B.n17 585
R435 B.n17 B.n16 585
R436 B.n769 B.n768 585
R437 B.n768 B.n767 585
R438 B.n19 B.n18 585
R439 B.n766 B.n19 585
R440 B.n764 B.n763 585
R441 B.n765 B.n764 585
R442 B.n762 B.n24 585
R443 B.n24 B.n23 585
R444 B.n761 B.n760 585
R445 B.n760 B.n759 585
R446 B.n26 B.n25 585
R447 B.n758 B.n26 585
R448 B.n756 B.n755 585
R449 B.n757 B.n756 585
R450 B.n754 B.n31 585
R451 B.n31 B.n30 585
R452 B.n753 B.n752 585
R453 B.n752 B.n751 585
R454 B.n33 B.n32 585
R455 B.n750 B.n33 585
R456 B.n748 B.n747 585
R457 B.n749 B.n748 585
R458 B.n746 B.n37 585
R459 B.n40 B.n37 585
R460 B.n745 B.n744 585
R461 B.n744 B.n743 585
R462 B.n39 B.n38 585
R463 B.n742 B.n39 585
R464 B.n740 B.n739 585
R465 B.n741 B.n740 585
R466 B.n738 B.n45 585
R467 B.n45 B.n44 585
R468 B.n737 B.n736 585
R469 B.n736 B.n735 585
R470 B.n47 B.n46 585
R471 B.n734 B.n47 585
R472 B.n732 B.n731 585
R473 B.n733 B.n732 585
R474 B.n730 B.n52 585
R475 B.n52 B.n51 585
R476 B.n729 B.n728 585
R477 B.n728 B.n727 585
R478 B.n54 B.n53 585
R479 B.n726 B.n54 585
R480 B.n724 B.n723 585
R481 B.n725 B.n724 585
R482 B.n722 B.n58 585
R483 B.n61 B.n58 585
R484 B.n721 B.n720 585
R485 B.n720 B.n719 585
R486 B.n60 B.n59 585
R487 B.n718 B.n60 585
R488 B.n716 B.n715 585
R489 B.n717 B.n716 585
R490 B.n714 B.n66 585
R491 B.n66 B.n65 585
R492 B.n713 B.n712 585
R493 B.n712 B.n711 585
R494 B.n68 B.n67 585
R495 B.n710 B.n68 585
R496 B.n708 B.n707 585
R497 B.n709 B.n708 585
R498 B.n706 B.n73 585
R499 B.n73 B.n72 585
R500 B.n705 B.n704 585
R501 B.n704 B.n703 585
R502 B.n75 B.n74 585
R503 B.n702 B.n75 585
R504 B.n700 B.n699 585
R505 B.n701 B.n700 585
R506 B.n698 B.n80 585
R507 B.n80 B.n79 585
R508 B.n697 B.n696 585
R509 B.n696 B.n695 585
R510 B.n82 B.n81 585
R511 B.n694 B.n82 585
R512 B.n692 B.n691 585
R513 B.n693 B.n692 585
R514 B.n690 B.n87 585
R515 B.n87 B.n86 585
R516 B.n689 B.n688 585
R517 B.n688 B.n687 585
R518 B.n89 B.n88 585
R519 B.n686 B.n89 585
R520 B.n684 B.n683 585
R521 B.n685 B.n684 585
R522 B.n682 B.n94 585
R523 B.n94 B.n93 585
R524 B.n681 B.n680 585
R525 B.n680 B.n679 585
R526 B.n96 B.n95 585
R527 B.n678 B.n96 585
R528 B.n676 B.n675 585
R529 B.n677 B.n676 585
R530 B.n674 B.n101 585
R531 B.n101 B.n100 585
R532 B.n785 B.n784 585
R533 B.n783 B.n2 585
R534 B.n672 B.n101 487.695
R535 B.n669 B.n125 487.695
R536 B.n345 B.n314 487.695
R537 B.n429 B.n316 487.695
R538 B.n670 B.n123 256.663
R539 B.n670 B.n122 256.663
R540 B.n670 B.n121 256.663
R541 B.n670 B.n120 256.663
R542 B.n670 B.n119 256.663
R543 B.n670 B.n118 256.663
R544 B.n670 B.n117 256.663
R545 B.n670 B.n116 256.663
R546 B.n670 B.n115 256.663
R547 B.n670 B.n114 256.663
R548 B.n670 B.n113 256.663
R549 B.n670 B.n112 256.663
R550 B.n670 B.n111 256.663
R551 B.n670 B.n110 256.663
R552 B.n670 B.n109 256.663
R553 B.n670 B.n108 256.663
R554 B.n670 B.n107 256.663
R555 B.n670 B.n106 256.663
R556 B.n670 B.n105 256.663
R557 B.n670 B.n104 256.663
R558 B.n671 B.n670 256.663
R559 B.n428 B.n427 256.663
R560 B.n427 B.n319 256.663
R561 B.n427 B.n320 256.663
R562 B.n427 B.n321 256.663
R563 B.n427 B.n322 256.663
R564 B.n427 B.n323 256.663
R565 B.n427 B.n324 256.663
R566 B.n427 B.n325 256.663
R567 B.n427 B.n326 256.663
R568 B.n427 B.n327 256.663
R569 B.n427 B.n328 256.663
R570 B.n427 B.n329 256.663
R571 B.n427 B.n330 256.663
R572 B.n427 B.n331 256.663
R573 B.n427 B.n332 256.663
R574 B.n427 B.n333 256.663
R575 B.n427 B.n334 256.663
R576 B.n427 B.n335 256.663
R577 B.n427 B.n336 256.663
R578 B.n427 B.n337 256.663
R579 B.n427 B.n338 256.663
R580 B.n787 B.n786 256.663
R581 B.n129 B.t5 231.749
R582 B.n126 B.t13 231.749
R583 B.n343 B.t9 231.749
R584 B.n340 B.t16 231.749
R585 B.n427 B.n315 167.488
R586 B.n670 B.n100 167.488
R587 B.n131 B.n103 163.367
R588 B.n135 B.n134 163.367
R589 B.n139 B.n138 163.367
R590 B.n143 B.n142 163.367
R591 B.n147 B.n146 163.367
R592 B.n151 B.n150 163.367
R593 B.n155 B.n154 163.367
R594 B.n159 B.n158 163.367
R595 B.n164 B.n163 163.367
R596 B.n168 B.n167 163.367
R597 B.n172 B.n171 163.367
R598 B.n176 B.n175 163.367
R599 B.n180 B.n179 163.367
R600 B.n184 B.n183 163.367
R601 B.n188 B.n187 163.367
R602 B.n192 B.n191 163.367
R603 B.n196 B.n195 163.367
R604 B.n200 B.n199 163.367
R605 B.n204 B.n203 163.367
R606 B.n208 B.n207 163.367
R607 B.n669 B.n124 163.367
R608 B.n435 B.n314 163.367
R609 B.n435 B.n312 163.367
R610 B.n439 B.n312 163.367
R611 B.n439 B.n306 163.367
R612 B.n447 B.n306 163.367
R613 B.n447 B.n304 163.367
R614 B.n451 B.n304 163.367
R615 B.n451 B.n298 163.367
R616 B.n459 B.n298 163.367
R617 B.n459 B.n296 163.367
R618 B.n463 B.n296 163.367
R619 B.n463 B.n290 163.367
R620 B.n471 B.n290 163.367
R621 B.n471 B.n288 163.367
R622 B.n475 B.n288 163.367
R623 B.n475 B.n282 163.367
R624 B.n483 B.n282 163.367
R625 B.n483 B.n280 163.367
R626 B.n487 B.n280 163.367
R627 B.n487 B.n274 163.367
R628 B.n495 B.n274 163.367
R629 B.n495 B.n272 163.367
R630 B.n499 B.n272 163.367
R631 B.n499 B.n267 163.367
R632 B.n508 B.n267 163.367
R633 B.n508 B.n265 163.367
R634 B.n512 B.n265 163.367
R635 B.n512 B.n259 163.367
R636 B.n520 B.n259 163.367
R637 B.n520 B.n257 163.367
R638 B.n524 B.n257 163.367
R639 B.n524 B.n251 163.367
R640 B.n532 B.n251 163.367
R641 B.n532 B.n249 163.367
R642 B.n536 B.n249 163.367
R643 B.n536 B.n244 163.367
R644 B.n545 B.n244 163.367
R645 B.n545 B.n242 163.367
R646 B.n549 B.n242 163.367
R647 B.n549 B.n236 163.367
R648 B.n557 B.n236 163.367
R649 B.n557 B.n234 163.367
R650 B.n561 B.n234 163.367
R651 B.n561 B.n228 163.367
R652 B.n569 B.n228 163.367
R653 B.n569 B.n226 163.367
R654 B.n573 B.n226 163.367
R655 B.n573 B.n220 163.367
R656 B.n581 B.n220 163.367
R657 B.n581 B.n218 163.367
R658 B.n586 B.n218 163.367
R659 B.n586 B.n212 163.367
R660 B.n594 B.n212 163.367
R661 B.n595 B.n594 163.367
R662 B.n595 B.n5 163.367
R663 B.n6 B.n5 163.367
R664 B.n7 B.n6 163.367
R665 B.n601 B.n7 163.367
R666 B.n602 B.n601 163.367
R667 B.n602 B.n13 163.367
R668 B.n14 B.n13 163.367
R669 B.n15 B.n14 163.367
R670 B.n607 B.n15 163.367
R671 B.n607 B.n20 163.367
R672 B.n21 B.n20 163.367
R673 B.n22 B.n21 163.367
R674 B.n612 B.n22 163.367
R675 B.n612 B.n27 163.367
R676 B.n28 B.n27 163.367
R677 B.n29 B.n28 163.367
R678 B.n617 B.n29 163.367
R679 B.n617 B.n34 163.367
R680 B.n35 B.n34 163.367
R681 B.n36 B.n35 163.367
R682 B.n622 B.n36 163.367
R683 B.n622 B.n41 163.367
R684 B.n42 B.n41 163.367
R685 B.n43 B.n42 163.367
R686 B.n627 B.n43 163.367
R687 B.n627 B.n48 163.367
R688 B.n49 B.n48 163.367
R689 B.n50 B.n49 163.367
R690 B.n632 B.n50 163.367
R691 B.n632 B.n55 163.367
R692 B.n56 B.n55 163.367
R693 B.n57 B.n56 163.367
R694 B.n637 B.n57 163.367
R695 B.n637 B.n62 163.367
R696 B.n63 B.n62 163.367
R697 B.n64 B.n63 163.367
R698 B.n642 B.n64 163.367
R699 B.n642 B.n69 163.367
R700 B.n70 B.n69 163.367
R701 B.n71 B.n70 163.367
R702 B.n647 B.n71 163.367
R703 B.n647 B.n76 163.367
R704 B.n77 B.n76 163.367
R705 B.n78 B.n77 163.367
R706 B.n652 B.n78 163.367
R707 B.n652 B.n83 163.367
R708 B.n84 B.n83 163.367
R709 B.n85 B.n84 163.367
R710 B.n657 B.n85 163.367
R711 B.n657 B.n90 163.367
R712 B.n91 B.n90 163.367
R713 B.n92 B.n91 163.367
R714 B.n662 B.n92 163.367
R715 B.n662 B.n97 163.367
R716 B.n98 B.n97 163.367
R717 B.n99 B.n98 163.367
R718 B.n125 B.n99 163.367
R719 B.n426 B.n318 163.367
R720 B.n426 B.n339 163.367
R721 B.n422 B.n421 163.367
R722 B.n418 B.n417 163.367
R723 B.n414 B.n413 163.367
R724 B.n410 B.n409 163.367
R725 B.n406 B.n405 163.367
R726 B.n402 B.n401 163.367
R727 B.n398 B.n397 163.367
R728 B.n394 B.n393 163.367
R729 B.n390 B.n389 163.367
R730 B.n386 B.n385 163.367
R731 B.n382 B.n381 163.367
R732 B.n377 B.n376 163.367
R733 B.n373 B.n372 163.367
R734 B.n369 B.n368 163.367
R735 B.n365 B.n364 163.367
R736 B.n361 B.n360 163.367
R737 B.n357 B.n356 163.367
R738 B.n353 B.n352 163.367
R739 B.n349 B.n348 163.367
R740 B.n433 B.n316 163.367
R741 B.n433 B.n310 163.367
R742 B.n441 B.n310 163.367
R743 B.n441 B.n308 163.367
R744 B.n445 B.n308 163.367
R745 B.n445 B.n302 163.367
R746 B.n453 B.n302 163.367
R747 B.n453 B.n300 163.367
R748 B.n457 B.n300 163.367
R749 B.n457 B.n294 163.367
R750 B.n465 B.n294 163.367
R751 B.n465 B.n292 163.367
R752 B.n469 B.n292 163.367
R753 B.n469 B.n286 163.367
R754 B.n477 B.n286 163.367
R755 B.n477 B.n284 163.367
R756 B.n481 B.n284 163.367
R757 B.n481 B.n278 163.367
R758 B.n489 B.n278 163.367
R759 B.n489 B.n276 163.367
R760 B.n493 B.n276 163.367
R761 B.n493 B.n270 163.367
R762 B.n502 B.n270 163.367
R763 B.n502 B.n268 163.367
R764 B.n506 B.n268 163.367
R765 B.n506 B.n263 163.367
R766 B.n514 B.n263 163.367
R767 B.n514 B.n261 163.367
R768 B.n518 B.n261 163.367
R769 B.n518 B.n255 163.367
R770 B.n526 B.n255 163.367
R771 B.n526 B.n253 163.367
R772 B.n530 B.n253 163.367
R773 B.n530 B.n247 163.367
R774 B.n539 B.n247 163.367
R775 B.n539 B.n245 163.367
R776 B.n543 B.n245 163.367
R777 B.n543 B.n240 163.367
R778 B.n551 B.n240 163.367
R779 B.n551 B.n238 163.367
R780 B.n555 B.n238 163.367
R781 B.n555 B.n232 163.367
R782 B.n563 B.n232 163.367
R783 B.n563 B.n230 163.367
R784 B.n567 B.n230 163.367
R785 B.n567 B.n224 163.367
R786 B.n575 B.n224 163.367
R787 B.n575 B.n222 163.367
R788 B.n579 B.n222 163.367
R789 B.n579 B.n216 163.367
R790 B.n588 B.n216 163.367
R791 B.n588 B.n214 163.367
R792 B.n592 B.n214 163.367
R793 B.n592 B.n3 163.367
R794 B.n785 B.n3 163.367
R795 B.n781 B.n2 163.367
R796 B.n781 B.n780 163.367
R797 B.n780 B.n9 163.367
R798 B.n776 B.n9 163.367
R799 B.n776 B.n11 163.367
R800 B.n772 B.n11 163.367
R801 B.n772 B.n17 163.367
R802 B.n768 B.n17 163.367
R803 B.n768 B.n19 163.367
R804 B.n764 B.n19 163.367
R805 B.n764 B.n24 163.367
R806 B.n760 B.n24 163.367
R807 B.n760 B.n26 163.367
R808 B.n756 B.n26 163.367
R809 B.n756 B.n31 163.367
R810 B.n752 B.n31 163.367
R811 B.n752 B.n33 163.367
R812 B.n748 B.n33 163.367
R813 B.n748 B.n37 163.367
R814 B.n744 B.n37 163.367
R815 B.n744 B.n39 163.367
R816 B.n740 B.n39 163.367
R817 B.n740 B.n45 163.367
R818 B.n736 B.n45 163.367
R819 B.n736 B.n47 163.367
R820 B.n732 B.n47 163.367
R821 B.n732 B.n52 163.367
R822 B.n728 B.n52 163.367
R823 B.n728 B.n54 163.367
R824 B.n724 B.n54 163.367
R825 B.n724 B.n58 163.367
R826 B.n720 B.n58 163.367
R827 B.n720 B.n60 163.367
R828 B.n716 B.n60 163.367
R829 B.n716 B.n66 163.367
R830 B.n712 B.n66 163.367
R831 B.n712 B.n68 163.367
R832 B.n708 B.n68 163.367
R833 B.n708 B.n73 163.367
R834 B.n704 B.n73 163.367
R835 B.n704 B.n75 163.367
R836 B.n700 B.n75 163.367
R837 B.n700 B.n80 163.367
R838 B.n696 B.n80 163.367
R839 B.n696 B.n82 163.367
R840 B.n692 B.n82 163.367
R841 B.n692 B.n87 163.367
R842 B.n688 B.n87 163.367
R843 B.n688 B.n89 163.367
R844 B.n684 B.n89 163.367
R845 B.n684 B.n94 163.367
R846 B.n680 B.n94 163.367
R847 B.n680 B.n96 163.367
R848 B.n676 B.n96 163.367
R849 B.n676 B.n101 163.367
R850 B.n126 B.t14 152.2
R851 B.n343 B.t12 152.2
R852 B.n129 B.t7 152.196
R853 B.n340 B.t18 152.196
R854 B.n434 B.n315 85.633
R855 B.n434 B.n311 85.633
R856 B.n440 B.n311 85.633
R857 B.n440 B.n307 85.633
R858 B.n446 B.n307 85.633
R859 B.n446 B.n303 85.633
R860 B.n452 B.n303 85.633
R861 B.n452 B.n299 85.633
R862 B.n458 B.n299 85.633
R863 B.n464 B.n295 85.633
R864 B.n464 B.n291 85.633
R865 B.n470 B.n291 85.633
R866 B.n470 B.n287 85.633
R867 B.n476 B.n287 85.633
R868 B.n476 B.n283 85.633
R869 B.n482 B.n283 85.633
R870 B.n482 B.n279 85.633
R871 B.n488 B.n279 85.633
R872 B.n488 B.n275 85.633
R873 B.n494 B.n275 85.633
R874 B.n494 B.n271 85.633
R875 B.n501 B.n271 85.633
R876 B.n501 B.n500 85.633
R877 B.n507 B.n264 85.633
R878 B.n513 B.n264 85.633
R879 B.n513 B.n260 85.633
R880 B.n519 B.n260 85.633
R881 B.n519 B.n256 85.633
R882 B.n525 B.n256 85.633
R883 B.n525 B.n252 85.633
R884 B.n531 B.n252 85.633
R885 B.n531 B.n248 85.633
R886 B.n538 B.n248 85.633
R887 B.n538 B.n537 85.633
R888 B.n544 B.n241 85.633
R889 B.n550 B.n241 85.633
R890 B.n550 B.n237 85.633
R891 B.n556 B.n237 85.633
R892 B.n556 B.n233 85.633
R893 B.n562 B.n233 85.633
R894 B.n562 B.n229 85.633
R895 B.n568 B.n229 85.633
R896 B.n568 B.n225 85.633
R897 B.n574 B.n225 85.633
R898 B.n580 B.n221 85.633
R899 B.n580 B.n217 85.633
R900 B.n587 B.n217 85.633
R901 B.n587 B.n213 85.633
R902 B.n593 B.n213 85.633
R903 B.n593 B.n4 85.633
R904 B.n784 B.n4 85.633
R905 B.n784 B.n783 85.633
R906 B.n783 B.n782 85.633
R907 B.n782 B.n8 85.633
R908 B.n12 B.n8 85.633
R909 B.n775 B.n12 85.633
R910 B.n775 B.n774 85.633
R911 B.n774 B.n773 85.633
R912 B.n773 B.n16 85.633
R913 B.n767 B.n766 85.633
R914 B.n766 B.n765 85.633
R915 B.n765 B.n23 85.633
R916 B.n759 B.n23 85.633
R917 B.n759 B.n758 85.633
R918 B.n758 B.n757 85.633
R919 B.n757 B.n30 85.633
R920 B.n751 B.n30 85.633
R921 B.n751 B.n750 85.633
R922 B.n750 B.n749 85.633
R923 B.n743 B.n40 85.633
R924 B.n743 B.n742 85.633
R925 B.n742 B.n741 85.633
R926 B.n741 B.n44 85.633
R927 B.n735 B.n44 85.633
R928 B.n735 B.n734 85.633
R929 B.n734 B.n733 85.633
R930 B.n733 B.n51 85.633
R931 B.n727 B.n51 85.633
R932 B.n727 B.n726 85.633
R933 B.n726 B.n725 85.633
R934 B.n719 B.n61 85.633
R935 B.n719 B.n718 85.633
R936 B.n718 B.n717 85.633
R937 B.n717 B.n65 85.633
R938 B.n711 B.n65 85.633
R939 B.n711 B.n710 85.633
R940 B.n710 B.n709 85.633
R941 B.n709 B.n72 85.633
R942 B.n703 B.n72 85.633
R943 B.n703 B.n702 85.633
R944 B.n702 B.n701 85.633
R945 B.n701 B.n79 85.633
R946 B.n695 B.n79 85.633
R947 B.n695 B.n694 85.633
R948 B.n693 B.n86 85.633
R949 B.n687 B.n86 85.633
R950 B.n687 B.n686 85.633
R951 B.n686 B.n685 85.633
R952 B.n685 B.n93 85.633
R953 B.n679 B.n93 85.633
R954 B.n679 B.n678 85.633
R955 B.n678 B.n677 85.633
R956 B.n677 B.n100 85.633
R957 B.n574 B.t19 81.8551
R958 B.n767 B.t0 81.8551
R959 B.n544 B.t1 79.3365
R960 B.n749 B.t3 79.3365
R961 B.n130 B.n129 78.352
R962 B.n127 B.n126 78.352
R963 B.n344 B.n343 78.352
R964 B.n341 B.n340 78.352
R965 B.t10 B.n295 76.8179
R966 B.n694 B.t6 76.8179
R967 B.n127 B.t15 73.8477
R968 B.n344 B.t11 73.8477
R969 B.n130 B.t8 73.8448
R970 B.n341 B.t17 73.8448
R971 B.n672 B.n671 71.676
R972 B.n131 B.n104 71.676
R973 B.n135 B.n105 71.676
R974 B.n139 B.n106 71.676
R975 B.n143 B.n107 71.676
R976 B.n147 B.n108 71.676
R977 B.n151 B.n109 71.676
R978 B.n155 B.n110 71.676
R979 B.n159 B.n111 71.676
R980 B.n164 B.n112 71.676
R981 B.n168 B.n113 71.676
R982 B.n172 B.n114 71.676
R983 B.n176 B.n115 71.676
R984 B.n180 B.n116 71.676
R985 B.n184 B.n117 71.676
R986 B.n188 B.n118 71.676
R987 B.n192 B.n119 71.676
R988 B.n196 B.n120 71.676
R989 B.n200 B.n121 71.676
R990 B.n204 B.n122 71.676
R991 B.n208 B.n123 71.676
R992 B.n124 B.n123 71.676
R993 B.n207 B.n122 71.676
R994 B.n203 B.n121 71.676
R995 B.n199 B.n120 71.676
R996 B.n195 B.n119 71.676
R997 B.n191 B.n118 71.676
R998 B.n187 B.n117 71.676
R999 B.n183 B.n116 71.676
R1000 B.n179 B.n115 71.676
R1001 B.n175 B.n114 71.676
R1002 B.n171 B.n113 71.676
R1003 B.n167 B.n112 71.676
R1004 B.n163 B.n111 71.676
R1005 B.n158 B.n110 71.676
R1006 B.n154 B.n109 71.676
R1007 B.n150 B.n108 71.676
R1008 B.n146 B.n107 71.676
R1009 B.n142 B.n106 71.676
R1010 B.n138 B.n105 71.676
R1011 B.n134 B.n104 71.676
R1012 B.n671 B.n103 71.676
R1013 B.n429 B.n428 71.676
R1014 B.n339 B.n319 71.676
R1015 B.n421 B.n320 71.676
R1016 B.n417 B.n321 71.676
R1017 B.n413 B.n322 71.676
R1018 B.n409 B.n323 71.676
R1019 B.n405 B.n324 71.676
R1020 B.n401 B.n325 71.676
R1021 B.n397 B.n326 71.676
R1022 B.n393 B.n327 71.676
R1023 B.n389 B.n328 71.676
R1024 B.n385 B.n329 71.676
R1025 B.n381 B.n330 71.676
R1026 B.n376 B.n331 71.676
R1027 B.n372 B.n332 71.676
R1028 B.n368 B.n333 71.676
R1029 B.n364 B.n334 71.676
R1030 B.n360 B.n335 71.676
R1031 B.n356 B.n336 71.676
R1032 B.n352 B.n337 71.676
R1033 B.n348 B.n338 71.676
R1034 B.n428 B.n318 71.676
R1035 B.n422 B.n319 71.676
R1036 B.n418 B.n320 71.676
R1037 B.n414 B.n321 71.676
R1038 B.n410 B.n322 71.676
R1039 B.n406 B.n323 71.676
R1040 B.n402 B.n324 71.676
R1041 B.n398 B.n325 71.676
R1042 B.n394 B.n326 71.676
R1043 B.n390 B.n327 71.676
R1044 B.n386 B.n328 71.676
R1045 B.n382 B.n329 71.676
R1046 B.n377 B.n330 71.676
R1047 B.n373 B.n331 71.676
R1048 B.n369 B.n332 71.676
R1049 B.n365 B.n333 71.676
R1050 B.n361 B.n334 71.676
R1051 B.n357 B.n335 71.676
R1052 B.n353 B.n336 71.676
R1053 B.n349 B.n337 71.676
R1054 B.n345 B.n338 71.676
R1055 B.n786 B.n785 71.676
R1056 B.n786 B.n2 71.676
R1057 B.n507 B.t4 69.2621
R1058 B.n725 B.t2 69.2621
R1059 B.n161 B.n130 59.5399
R1060 B.n128 B.n127 59.5399
R1061 B.n379 B.n344 59.5399
R1062 B.n342 B.n341 59.5399
R1063 B.n431 B.n430 31.6883
R1064 B.n346 B.n313 31.6883
R1065 B.n668 B.n667 31.6883
R1066 B.n674 B.n673 31.6883
R1067 B B.n787 18.0485
R1068 B.n500 B.t4 16.3714
R1069 B.n61 B.t2 16.3714
R1070 B.n432 B.n431 10.6151
R1071 B.n432 B.n309 10.6151
R1072 B.n442 B.n309 10.6151
R1073 B.n443 B.n442 10.6151
R1074 B.n444 B.n443 10.6151
R1075 B.n444 B.n301 10.6151
R1076 B.n454 B.n301 10.6151
R1077 B.n455 B.n454 10.6151
R1078 B.n456 B.n455 10.6151
R1079 B.n456 B.n293 10.6151
R1080 B.n466 B.n293 10.6151
R1081 B.n467 B.n466 10.6151
R1082 B.n468 B.n467 10.6151
R1083 B.n468 B.n285 10.6151
R1084 B.n478 B.n285 10.6151
R1085 B.n479 B.n478 10.6151
R1086 B.n480 B.n479 10.6151
R1087 B.n480 B.n277 10.6151
R1088 B.n490 B.n277 10.6151
R1089 B.n491 B.n490 10.6151
R1090 B.n492 B.n491 10.6151
R1091 B.n492 B.n269 10.6151
R1092 B.n503 B.n269 10.6151
R1093 B.n504 B.n503 10.6151
R1094 B.n505 B.n504 10.6151
R1095 B.n505 B.n262 10.6151
R1096 B.n515 B.n262 10.6151
R1097 B.n516 B.n515 10.6151
R1098 B.n517 B.n516 10.6151
R1099 B.n517 B.n254 10.6151
R1100 B.n527 B.n254 10.6151
R1101 B.n528 B.n527 10.6151
R1102 B.n529 B.n528 10.6151
R1103 B.n529 B.n246 10.6151
R1104 B.n540 B.n246 10.6151
R1105 B.n541 B.n540 10.6151
R1106 B.n542 B.n541 10.6151
R1107 B.n542 B.n239 10.6151
R1108 B.n552 B.n239 10.6151
R1109 B.n553 B.n552 10.6151
R1110 B.n554 B.n553 10.6151
R1111 B.n554 B.n231 10.6151
R1112 B.n564 B.n231 10.6151
R1113 B.n565 B.n564 10.6151
R1114 B.n566 B.n565 10.6151
R1115 B.n566 B.n223 10.6151
R1116 B.n576 B.n223 10.6151
R1117 B.n577 B.n576 10.6151
R1118 B.n578 B.n577 10.6151
R1119 B.n578 B.n215 10.6151
R1120 B.n589 B.n215 10.6151
R1121 B.n590 B.n589 10.6151
R1122 B.n591 B.n590 10.6151
R1123 B.n591 B.n0 10.6151
R1124 B.n430 B.n317 10.6151
R1125 B.n425 B.n317 10.6151
R1126 B.n425 B.n424 10.6151
R1127 B.n424 B.n423 10.6151
R1128 B.n423 B.n420 10.6151
R1129 B.n420 B.n419 10.6151
R1130 B.n419 B.n416 10.6151
R1131 B.n416 B.n415 10.6151
R1132 B.n415 B.n412 10.6151
R1133 B.n412 B.n411 10.6151
R1134 B.n411 B.n408 10.6151
R1135 B.n408 B.n407 10.6151
R1136 B.n407 B.n404 10.6151
R1137 B.n404 B.n403 10.6151
R1138 B.n403 B.n400 10.6151
R1139 B.n400 B.n399 10.6151
R1140 B.n396 B.n395 10.6151
R1141 B.n395 B.n392 10.6151
R1142 B.n392 B.n391 10.6151
R1143 B.n391 B.n388 10.6151
R1144 B.n388 B.n387 10.6151
R1145 B.n387 B.n384 10.6151
R1146 B.n384 B.n383 10.6151
R1147 B.n383 B.n380 10.6151
R1148 B.n378 B.n375 10.6151
R1149 B.n375 B.n374 10.6151
R1150 B.n374 B.n371 10.6151
R1151 B.n371 B.n370 10.6151
R1152 B.n370 B.n367 10.6151
R1153 B.n367 B.n366 10.6151
R1154 B.n366 B.n363 10.6151
R1155 B.n363 B.n362 10.6151
R1156 B.n362 B.n359 10.6151
R1157 B.n359 B.n358 10.6151
R1158 B.n358 B.n355 10.6151
R1159 B.n355 B.n354 10.6151
R1160 B.n354 B.n351 10.6151
R1161 B.n351 B.n350 10.6151
R1162 B.n350 B.n347 10.6151
R1163 B.n347 B.n346 10.6151
R1164 B.n436 B.n313 10.6151
R1165 B.n437 B.n436 10.6151
R1166 B.n438 B.n437 10.6151
R1167 B.n438 B.n305 10.6151
R1168 B.n448 B.n305 10.6151
R1169 B.n449 B.n448 10.6151
R1170 B.n450 B.n449 10.6151
R1171 B.n450 B.n297 10.6151
R1172 B.n460 B.n297 10.6151
R1173 B.n461 B.n460 10.6151
R1174 B.n462 B.n461 10.6151
R1175 B.n462 B.n289 10.6151
R1176 B.n472 B.n289 10.6151
R1177 B.n473 B.n472 10.6151
R1178 B.n474 B.n473 10.6151
R1179 B.n474 B.n281 10.6151
R1180 B.n484 B.n281 10.6151
R1181 B.n485 B.n484 10.6151
R1182 B.n486 B.n485 10.6151
R1183 B.n486 B.n273 10.6151
R1184 B.n496 B.n273 10.6151
R1185 B.n497 B.n496 10.6151
R1186 B.n498 B.n497 10.6151
R1187 B.n498 B.n266 10.6151
R1188 B.n509 B.n266 10.6151
R1189 B.n510 B.n509 10.6151
R1190 B.n511 B.n510 10.6151
R1191 B.n511 B.n258 10.6151
R1192 B.n521 B.n258 10.6151
R1193 B.n522 B.n521 10.6151
R1194 B.n523 B.n522 10.6151
R1195 B.n523 B.n250 10.6151
R1196 B.n533 B.n250 10.6151
R1197 B.n534 B.n533 10.6151
R1198 B.n535 B.n534 10.6151
R1199 B.n535 B.n243 10.6151
R1200 B.n546 B.n243 10.6151
R1201 B.n547 B.n546 10.6151
R1202 B.n548 B.n547 10.6151
R1203 B.n548 B.n235 10.6151
R1204 B.n558 B.n235 10.6151
R1205 B.n559 B.n558 10.6151
R1206 B.n560 B.n559 10.6151
R1207 B.n560 B.n227 10.6151
R1208 B.n570 B.n227 10.6151
R1209 B.n571 B.n570 10.6151
R1210 B.n572 B.n571 10.6151
R1211 B.n572 B.n219 10.6151
R1212 B.n582 B.n219 10.6151
R1213 B.n583 B.n582 10.6151
R1214 B.n585 B.n583 10.6151
R1215 B.n585 B.n584 10.6151
R1216 B.n584 B.n211 10.6151
R1217 B.n596 B.n211 10.6151
R1218 B.n597 B.n596 10.6151
R1219 B.n598 B.n597 10.6151
R1220 B.n599 B.n598 10.6151
R1221 B.n600 B.n599 10.6151
R1222 B.n603 B.n600 10.6151
R1223 B.n604 B.n603 10.6151
R1224 B.n605 B.n604 10.6151
R1225 B.n606 B.n605 10.6151
R1226 B.n608 B.n606 10.6151
R1227 B.n609 B.n608 10.6151
R1228 B.n610 B.n609 10.6151
R1229 B.n611 B.n610 10.6151
R1230 B.n613 B.n611 10.6151
R1231 B.n614 B.n613 10.6151
R1232 B.n615 B.n614 10.6151
R1233 B.n616 B.n615 10.6151
R1234 B.n618 B.n616 10.6151
R1235 B.n619 B.n618 10.6151
R1236 B.n620 B.n619 10.6151
R1237 B.n621 B.n620 10.6151
R1238 B.n623 B.n621 10.6151
R1239 B.n624 B.n623 10.6151
R1240 B.n625 B.n624 10.6151
R1241 B.n626 B.n625 10.6151
R1242 B.n628 B.n626 10.6151
R1243 B.n629 B.n628 10.6151
R1244 B.n630 B.n629 10.6151
R1245 B.n631 B.n630 10.6151
R1246 B.n633 B.n631 10.6151
R1247 B.n634 B.n633 10.6151
R1248 B.n635 B.n634 10.6151
R1249 B.n636 B.n635 10.6151
R1250 B.n638 B.n636 10.6151
R1251 B.n639 B.n638 10.6151
R1252 B.n640 B.n639 10.6151
R1253 B.n641 B.n640 10.6151
R1254 B.n643 B.n641 10.6151
R1255 B.n644 B.n643 10.6151
R1256 B.n645 B.n644 10.6151
R1257 B.n646 B.n645 10.6151
R1258 B.n648 B.n646 10.6151
R1259 B.n649 B.n648 10.6151
R1260 B.n650 B.n649 10.6151
R1261 B.n651 B.n650 10.6151
R1262 B.n653 B.n651 10.6151
R1263 B.n654 B.n653 10.6151
R1264 B.n655 B.n654 10.6151
R1265 B.n656 B.n655 10.6151
R1266 B.n658 B.n656 10.6151
R1267 B.n659 B.n658 10.6151
R1268 B.n660 B.n659 10.6151
R1269 B.n661 B.n660 10.6151
R1270 B.n663 B.n661 10.6151
R1271 B.n664 B.n663 10.6151
R1272 B.n665 B.n664 10.6151
R1273 B.n666 B.n665 10.6151
R1274 B.n667 B.n666 10.6151
R1275 B.n779 B.n1 10.6151
R1276 B.n779 B.n778 10.6151
R1277 B.n778 B.n777 10.6151
R1278 B.n777 B.n10 10.6151
R1279 B.n771 B.n10 10.6151
R1280 B.n771 B.n770 10.6151
R1281 B.n770 B.n769 10.6151
R1282 B.n769 B.n18 10.6151
R1283 B.n763 B.n18 10.6151
R1284 B.n763 B.n762 10.6151
R1285 B.n762 B.n761 10.6151
R1286 B.n761 B.n25 10.6151
R1287 B.n755 B.n25 10.6151
R1288 B.n755 B.n754 10.6151
R1289 B.n754 B.n753 10.6151
R1290 B.n753 B.n32 10.6151
R1291 B.n747 B.n32 10.6151
R1292 B.n747 B.n746 10.6151
R1293 B.n746 B.n745 10.6151
R1294 B.n745 B.n38 10.6151
R1295 B.n739 B.n38 10.6151
R1296 B.n739 B.n738 10.6151
R1297 B.n738 B.n737 10.6151
R1298 B.n737 B.n46 10.6151
R1299 B.n731 B.n46 10.6151
R1300 B.n731 B.n730 10.6151
R1301 B.n730 B.n729 10.6151
R1302 B.n729 B.n53 10.6151
R1303 B.n723 B.n53 10.6151
R1304 B.n723 B.n722 10.6151
R1305 B.n722 B.n721 10.6151
R1306 B.n721 B.n59 10.6151
R1307 B.n715 B.n59 10.6151
R1308 B.n715 B.n714 10.6151
R1309 B.n714 B.n713 10.6151
R1310 B.n713 B.n67 10.6151
R1311 B.n707 B.n67 10.6151
R1312 B.n707 B.n706 10.6151
R1313 B.n706 B.n705 10.6151
R1314 B.n705 B.n74 10.6151
R1315 B.n699 B.n74 10.6151
R1316 B.n699 B.n698 10.6151
R1317 B.n698 B.n697 10.6151
R1318 B.n697 B.n81 10.6151
R1319 B.n691 B.n81 10.6151
R1320 B.n691 B.n690 10.6151
R1321 B.n690 B.n689 10.6151
R1322 B.n689 B.n88 10.6151
R1323 B.n683 B.n88 10.6151
R1324 B.n683 B.n682 10.6151
R1325 B.n682 B.n681 10.6151
R1326 B.n681 B.n95 10.6151
R1327 B.n675 B.n95 10.6151
R1328 B.n675 B.n674 10.6151
R1329 B.n673 B.n102 10.6151
R1330 B.n132 B.n102 10.6151
R1331 B.n133 B.n132 10.6151
R1332 B.n136 B.n133 10.6151
R1333 B.n137 B.n136 10.6151
R1334 B.n140 B.n137 10.6151
R1335 B.n141 B.n140 10.6151
R1336 B.n144 B.n141 10.6151
R1337 B.n145 B.n144 10.6151
R1338 B.n148 B.n145 10.6151
R1339 B.n149 B.n148 10.6151
R1340 B.n152 B.n149 10.6151
R1341 B.n153 B.n152 10.6151
R1342 B.n156 B.n153 10.6151
R1343 B.n157 B.n156 10.6151
R1344 B.n160 B.n157 10.6151
R1345 B.n165 B.n162 10.6151
R1346 B.n166 B.n165 10.6151
R1347 B.n169 B.n166 10.6151
R1348 B.n170 B.n169 10.6151
R1349 B.n173 B.n170 10.6151
R1350 B.n174 B.n173 10.6151
R1351 B.n177 B.n174 10.6151
R1352 B.n178 B.n177 10.6151
R1353 B.n182 B.n181 10.6151
R1354 B.n185 B.n182 10.6151
R1355 B.n186 B.n185 10.6151
R1356 B.n189 B.n186 10.6151
R1357 B.n190 B.n189 10.6151
R1358 B.n193 B.n190 10.6151
R1359 B.n194 B.n193 10.6151
R1360 B.n197 B.n194 10.6151
R1361 B.n198 B.n197 10.6151
R1362 B.n201 B.n198 10.6151
R1363 B.n202 B.n201 10.6151
R1364 B.n205 B.n202 10.6151
R1365 B.n206 B.n205 10.6151
R1366 B.n209 B.n206 10.6151
R1367 B.n210 B.n209 10.6151
R1368 B.n668 B.n210 10.6151
R1369 B.n458 B.t10 8.81561
R1370 B.t6 B.n693 8.81561
R1371 B.n787 B.n0 8.11757
R1372 B.n787 B.n1 8.11757
R1373 B.n396 B.n342 6.5566
R1374 B.n380 B.n379 6.5566
R1375 B.n162 B.n161 6.5566
R1376 B.n178 B.n128 6.5566
R1377 B.n537 B.t1 6.29701
R1378 B.n40 B.t3 6.29701
R1379 B.n399 B.n342 4.05904
R1380 B.n379 B.n378 4.05904
R1381 B.n161 B.n160 4.05904
R1382 B.n181 B.n128 4.05904
R1383 B.t19 B.n221 3.7784
R1384 B.t0 B.n16 3.7784
R1385 VP.n16 VP.n13 161.3
R1386 VP.n18 VP.n17 161.3
R1387 VP.n19 VP.n12 161.3
R1388 VP.n21 VP.n20 161.3
R1389 VP.n22 VP.n11 161.3
R1390 VP.n24 VP.n23 161.3
R1391 VP.n25 VP.n10 161.3
R1392 VP.n27 VP.n26 161.3
R1393 VP.n56 VP.n55 161.3
R1394 VP.n54 VP.n1 161.3
R1395 VP.n53 VP.n52 161.3
R1396 VP.n51 VP.n2 161.3
R1397 VP.n50 VP.n49 161.3
R1398 VP.n48 VP.n3 161.3
R1399 VP.n47 VP.n46 161.3
R1400 VP.n45 VP.n4 161.3
R1401 VP.n44 VP.n43 161.3
R1402 VP.n42 VP.n5 161.3
R1403 VP.n41 VP.n40 161.3
R1404 VP.n39 VP.n6 161.3
R1405 VP.n38 VP.n37 161.3
R1406 VP.n36 VP.n7 161.3
R1407 VP.n35 VP.n34 161.3
R1408 VP.n33 VP.n8 161.3
R1409 VP.n32 VP.n31 161.3
R1410 VP.n30 VP.n29 88.2782
R1411 VP.n57 VP.n0 88.2782
R1412 VP.n28 VP.n9 88.2782
R1413 VP.n15 VP.t5 55.2165
R1414 VP.n15 VP.n14 50.5906
R1415 VP.n29 VP.n28 46.5753
R1416 VP.n37 VP.n36 42.5146
R1417 VP.n49 VP.n2 42.5146
R1418 VP.n20 VP.n11 42.5146
R1419 VP.n37 VP.n6 38.6395
R1420 VP.n49 VP.n48 38.6395
R1421 VP.n20 VP.n19 38.6395
R1422 VP.n31 VP.n8 24.5923
R1423 VP.n35 VP.n8 24.5923
R1424 VP.n36 VP.n35 24.5923
R1425 VP.n41 VP.n6 24.5923
R1426 VP.n42 VP.n41 24.5923
R1427 VP.n43 VP.n42 24.5923
R1428 VP.n43 VP.n4 24.5923
R1429 VP.n47 VP.n4 24.5923
R1430 VP.n48 VP.n47 24.5923
R1431 VP.n53 VP.n2 24.5923
R1432 VP.n54 VP.n53 24.5923
R1433 VP.n55 VP.n54 24.5923
R1434 VP.n24 VP.n11 24.5923
R1435 VP.n25 VP.n24 24.5923
R1436 VP.n26 VP.n25 24.5923
R1437 VP.n14 VP.n13 24.5923
R1438 VP.n18 VP.n13 24.5923
R1439 VP.n19 VP.n18 24.5923
R1440 VP.n43 VP.t4 22.4765
R1441 VP.n30 VP.t1 22.4765
R1442 VP.n0 VP.t0 22.4765
R1443 VP.n14 VP.t3 22.4765
R1444 VP.n9 VP.t2 22.4765
R1445 VP.n16 VP.n15 2.47297
R1446 VP.n31 VP.n30 1.96785
R1447 VP.n55 VP.n0 1.96785
R1448 VP.n26 VP.n9 1.96785
R1449 VP.n28 VP.n27 0.354861
R1450 VP.n32 VP.n29 0.354861
R1451 VP.n57 VP.n56 0.354861
R1452 VP VP.n57 0.267071
R1453 VP.n17 VP.n16 0.189894
R1454 VP.n17 VP.n12 0.189894
R1455 VP.n21 VP.n12 0.189894
R1456 VP.n22 VP.n21 0.189894
R1457 VP.n23 VP.n22 0.189894
R1458 VP.n23 VP.n10 0.189894
R1459 VP.n27 VP.n10 0.189894
R1460 VP.n33 VP.n32 0.189894
R1461 VP.n34 VP.n33 0.189894
R1462 VP.n34 VP.n7 0.189894
R1463 VP.n38 VP.n7 0.189894
R1464 VP.n39 VP.n38 0.189894
R1465 VP.n40 VP.n39 0.189894
R1466 VP.n40 VP.n5 0.189894
R1467 VP.n44 VP.n5 0.189894
R1468 VP.n45 VP.n44 0.189894
R1469 VP.n46 VP.n45 0.189894
R1470 VP.n46 VP.n3 0.189894
R1471 VP.n50 VP.n3 0.189894
R1472 VP.n51 VP.n50 0.189894
R1473 VP.n52 VP.n51 0.189894
R1474 VP.n52 VP.n1 0.189894
R1475 VP.n56 VP.n1 0.189894
R1476 VTAIL.n7 VTAIL.t5 64.0164
R1477 VTAIL.n11 VTAIL.t1 64.0164
R1478 VTAIL.n2 VTAIL.t6 64.0164
R1479 VTAIL.n10 VTAIL.t8 64.0164
R1480 VTAIL.n9 VTAIL.n8 58.294
R1481 VTAIL.n6 VTAIL.n5 58.294
R1482 VTAIL.n1 VTAIL.n0 58.2937
R1483 VTAIL.n4 VTAIL.n3 58.2937
R1484 VTAIL.n6 VTAIL.n4 22.3152
R1485 VTAIL.n11 VTAIL.n10 18.8324
R1486 VTAIL.n0 VTAIL.t2 5.72304
R1487 VTAIL.n0 VTAIL.t3 5.72304
R1488 VTAIL.n3 VTAIL.t11 5.72304
R1489 VTAIL.n3 VTAIL.t9 5.72304
R1490 VTAIL.n8 VTAIL.t7 5.72304
R1491 VTAIL.n8 VTAIL.t10 5.72304
R1492 VTAIL.n5 VTAIL.t4 5.72304
R1493 VTAIL.n5 VTAIL.t0 5.72304
R1494 VTAIL.n7 VTAIL.n6 3.48326
R1495 VTAIL.n10 VTAIL.n9 3.48326
R1496 VTAIL.n4 VTAIL.n2 3.48326
R1497 VTAIL VTAIL.n11 2.55438
R1498 VTAIL.n9 VTAIL.n7 2.21171
R1499 VTAIL.n2 VTAIL.n1 2.21171
R1500 VTAIL VTAIL.n1 0.929379
R1501 VDD1 VDD1.t0 83.3655
R1502 VDD1.n1 VDD1.t4 83.2519
R1503 VDD1.n1 VDD1.n0 75.7879
R1504 VDD1.n3 VDD1.n2 74.9726
R1505 VDD1.n3 VDD1.n1 40.3414
R1506 VDD1.n2 VDD1.t2 5.72304
R1507 VDD1.n2 VDD1.t3 5.72304
R1508 VDD1.n0 VDD1.t1 5.72304
R1509 VDD1.n0 VDD1.t5 5.72304
R1510 VDD1 VDD1.n3 0.813
R1511 VN.n38 VN.n37 161.3
R1512 VN.n36 VN.n21 161.3
R1513 VN.n35 VN.n34 161.3
R1514 VN.n33 VN.n22 161.3
R1515 VN.n32 VN.n31 161.3
R1516 VN.n30 VN.n23 161.3
R1517 VN.n29 VN.n28 161.3
R1518 VN.n27 VN.n24 161.3
R1519 VN.n18 VN.n17 161.3
R1520 VN.n16 VN.n1 161.3
R1521 VN.n15 VN.n14 161.3
R1522 VN.n13 VN.n2 161.3
R1523 VN.n12 VN.n11 161.3
R1524 VN.n10 VN.n3 161.3
R1525 VN.n9 VN.n8 161.3
R1526 VN.n7 VN.n4 161.3
R1527 VN.n19 VN.n0 88.2782
R1528 VN.n39 VN.n20 88.2782
R1529 VN.n26 VN.t3 55.2166
R1530 VN.n6 VN.t0 55.2166
R1531 VN.n6 VN.n5 50.5906
R1532 VN.n26 VN.n25 50.5906
R1533 VN VN.n39 46.7406
R1534 VN.n11 VN.n2 42.5146
R1535 VN.n31 VN.n22 42.5146
R1536 VN.n11 VN.n10 38.6395
R1537 VN.n31 VN.n30 38.6395
R1538 VN.n5 VN.n4 24.5923
R1539 VN.n9 VN.n4 24.5923
R1540 VN.n10 VN.n9 24.5923
R1541 VN.n15 VN.n2 24.5923
R1542 VN.n16 VN.n15 24.5923
R1543 VN.n17 VN.n16 24.5923
R1544 VN.n30 VN.n29 24.5923
R1545 VN.n29 VN.n24 24.5923
R1546 VN.n25 VN.n24 24.5923
R1547 VN.n37 VN.n36 24.5923
R1548 VN.n36 VN.n35 24.5923
R1549 VN.n35 VN.n22 24.5923
R1550 VN.n5 VN.t5 22.4765
R1551 VN.n0 VN.t1 22.4765
R1552 VN.n25 VN.t2 22.4765
R1553 VN.n20 VN.t4 22.4765
R1554 VN.n27 VN.n26 2.47298
R1555 VN.n7 VN.n6 2.47298
R1556 VN.n17 VN.n0 1.96785
R1557 VN.n37 VN.n20 1.96785
R1558 VN.n39 VN.n38 0.354861
R1559 VN.n19 VN.n18 0.354861
R1560 VN VN.n19 0.267071
R1561 VN.n38 VN.n21 0.189894
R1562 VN.n34 VN.n21 0.189894
R1563 VN.n34 VN.n33 0.189894
R1564 VN.n33 VN.n32 0.189894
R1565 VN.n32 VN.n23 0.189894
R1566 VN.n28 VN.n23 0.189894
R1567 VN.n28 VN.n27 0.189894
R1568 VN.n8 VN.n7 0.189894
R1569 VN.n8 VN.n3 0.189894
R1570 VN.n12 VN.n3 0.189894
R1571 VN.n13 VN.n12 0.189894
R1572 VN.n14 VN.n13 0.189894
R1573 VN.n14 VN.n1 0.189894
R1574 VN.n18 VN.n1 0.189894
R1575 VDD2.n1 VDD2.t5 83.2519
R1576 VDD2.n2 VDD2.t1 80.6952
R1577 VDD2.n1 VDD2.n0 75.7879
R1578 VDD2 VDD2.n3 75.7851
R1579 VDD2.n2 VDD2.n1 38.017
R1580 VDD2.n3 VDD2.t3 5.72304
R1581 VDD2.n3 VDD2.t2 5.72304
R1582 VDD2.n0 VDD2.t0 5.72304
R1583 VDD2.n0 VDD2.t4 5.72304
R1584 VDD2 VDD2.n2 2.67076
C0 VP VDD1 2.74648f
C1 VTAIL VDD1 5.38005f
C2 VN VP 6.4268f
C3 VN VTAIL 3.4352f
C4 VDD1 VDD2 1.83827f
C5 VN VDD2 2.3489f
C6 VP VTAIL 3.44943f
C7 VP VDD2 0.557447f
C8 VTAIL VDD2 5.4406f
C9 VN VDD1 0.157122f
C10 VDD2 B 5.30405f
C11 VDD1 B 5.681793f
C12 VTAIL B 4.573576f
C13 VN B 15.42387f
C14 VP B 14.033503f
C15 VDD2.t5 B 0.599855f
C16 VDD2.t0 B 0.060416f
C17 VDD2.t4 B 0.060416f
C18 VDD2.n0 B 0.46826f
C19 VDD2.n1 B 2.49264f
C20 VDD2.t1 B 0.587591f
C21 VDD2.n2 B 2.11621f
C22 VDD2.t3 B 0.060416f
C23 VDD2.t2 B 0.060416f
C24 VDD2.n3 B 0.468232f
C25 VN.t1 B 0.796446f
C26 VN.n0 B 0.404316f
C27 VN.n1 B 0.0245f
C28 VN.n2 B 0.047891f
C29 VN.n3 B 0.0245f
C30 VN.n4 B 0.045432f
C31 VN.t5 B 0.796446f
C32 VN.n5 B 0.415867f
C33 VN.t0 B 1.09755f
C34 VN.n6 B 0.419716f
C35 VN.n7 B 0.312323f
C36 VN.n8 B 0.0245f
C37 VN.n9 B 0.045432f
C38 VN.n10 B 0.048857f
C39 VN.n11 B 0.019913f
C40 VN.n12 B 0.0245f
C41 VN.n13 B 0.0245f
C42 VN.n14 B 0.0245f
C43 VN.n15 B 0.045432f
C44 VN.n16 B 0.045432f
C45 VN.n17 B 0.024798f
C46 VN.n18 B 0.039536f
C47 VN.n19 B 0.074567f
C48 VN.t4 B 0.796446f
C49 VN.n20 B 0.404316f
C50 VN.n21 B 0.0245f
C51 VN.n22 B 0.047891f
C52 VN.n23 B 0.0245f
C53 VN.n24 B 0.045432f
C54 VN.t3 B 1.09755f
C55 VN.t2 B 0.796446f
C56 VN.n25 B 0.415867f
C57 VN.n26 B 0.419716f
C58 VN.n27 B 0.312323f
C59 VN.n28 B 0.0245f
C60 VN.n29 B 0.045432f
C61 VN.n30 B 0.048857f
C62 VN.n31 B 0.019913f
C63 VN.n32 B 0.0245f
C64 VN.n33 B 0.0245f
C65 VN.n34 B 0.0245f
C66 VN.n35 B 0.045432f
C67 VN.n36 B 0.045432f
C68 VN.n37 B 0.024798f
C69 VN.n38 B 0.039536f
C70 VN.n39 B 1.28119f
C71 VDD1.t0 B 0.625213f
C72 VDD1.t4 B 0.624398f
C73 VDD1.t1 B 0.062888f
C74 VDD1.t5 B 0.062888f
C75 VDD1.n0 B 0.487419f
C76 VDD1.n1 B 2.72673f
C77 VDD1.t2 B 0.062888f
C78 VDD1.t3 B 0.062888f
C79 VDD1.n2 B 0.482003f
C80 VDD1.n3 B 2.2342f
C81 VTAIL.t2 B 0.087861f
C82 VTAIL.t3 B 0.087861f
C83 VTAIL.n0 B 0.605242f
C84 VTAIL.n1 B 0.593992f
C85 VTAIL.t6 B 0.777191f
C86 VTAIL.n2 B 0.9261f
C87 VTAIL.t11 B 0.087861f
C88 VTAIL.t9 B 0.087861f
C89 VTAIL.n3 B 0.605242f
C90 VTAIL.n4 B 2.09605f
C91 VTAIL.t4 B 0.087861f
C92 VTAIL.t0 B 0.087861f
C93 VTAIL.n5 B 0.605245f
C94 VTAIL.n6 B 2.09605f
C95 VTAIL.t5 B 0.777197f
C96 VTAIL.n7 B 0.926095f
C97 VTAIL.t7 B 0.087861f
C98 VTAIL.t10 B 0.087861f
C99 VTAIL.n8 B 0.605245f
C100 VTAIL.n9 B 0.858425f
C101 VTAIL.t8 B 0.777191f
C102 VTAIL.n10 B 1.80311f
C103 VTAIL.t1 B 0.777191f
C104 VTAIL.n11 B 1.70693f
C105 VP.t0 B 0.825124f
C106 VP.n0 B 0.418874f
C107 VP.n1 B 0.025382f
C108 VP.n2 B 0.049615f
C109 VP.n3 B 0.025382f
C110 VP.n4 B 0.047068f
C111 VP.n5 B 0.025382f
C112 VP.t4 B 0.825124f
C113 VP.n6 B 0.050616f
C114 VP.n7 B 0.025382f
C115 VP.n8 B 0.047068f
C116 VP.t2 B 0.825124f
C117 VP.n9 B 0.418874f
C118 VP.n10 B 0.025382f
C119 VP.n11 B 0.049615f
C120 VP.n12 B 0.025382f
C121 VP.n13 B 0.047068f
C122 VP.t5 B 1.13706f
C123 VP.t3 B 0.825124f
C124 VP.n14 B 0.430841f
C125 VP.n15 B 0.434829f
C126 VP.n16 B 0.323569f
C127 VP.n17 B 0.025382f
C128 VP.n18 B 0.047068f
C129 VP.n19 B 0.050616f
C130 VP.n20 B 0.02063f
C131 VP.n21 B 0.025382f
C132 VP.n22 B 0.025382f
C133 VP.n23 B 0.025382f
C134 VP.n24 B 0.047068f
C135 VP.n25 B 0.047068f
C136 VP.n26 B 0.025691f
C137 VP.n27 B 0.040959f
C138 VP.n28 B 1.31668f
C139 VP.n29 B 1.33632f
C140 VP.t1 B 0.825124f
C141 VP.n30 B 0.418874f
C142 VP.n31 B 0.025691f
C143 VP.n32 B 0.040959f
C144 VP.n33 B 0.025382f
C145 VP.n34 B 0.025382f
C146 VP.n35 B 0.047068f
C147 VP.n36 B 0.049615f
C148 VP.n37 B 0.02063f
C149 VP.n38 B 0.025382f
C150 VP.n39 B 0.025382f
C151 VP.n40 B 0.025382f
C152 VP.n41 B 0.047068f
C153 VP.n42 B 0.047068f
C154 VP.n43 B 0.351432f
C155 VP.n44 B 0.025382f
C156 VP.n45 B 0.025382f
C157 VP.n46 B 0.025382f
C158 VP.n47 B 0.047068f
C159 VP.n48 B 0.050616f
C160 VP.n49 B 0.02063f
C161 VP.n50 B 0.025382f
C162 VP.n51 B 0.025382f
C163 VP.n52 B 0.025382f
C164 VP.n53 B 0.047068f
C165 VP.n54 B 0.047068f
C166 VP.n55 B 0.025691f
C167 VP.n56 B 0.040959f
C168 VP.n57 B 0.077252f
.ends

