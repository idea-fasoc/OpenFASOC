* NGSPICE file created from diff_pair_sample_0196.ext - technology: sky130A

.subckt diff_pair_sample_0196 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=2.24895 ps=13.96 w=13.63 l=0.81
X1 VTAIL.t6 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=2.24895 ps=13.96 w=13.63 l=0.81
X2 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=2.24895 ps=13.96 w=13.63 l=0.81
X3 VDD1.t3 VP.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=2.24895 ps=13.96 w=13.63 l=0.81
X4 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=0 ps=0 w=13.63 l=0.81
X5 VDD1.t2 VP.t3 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=5.3157 ps=28.04 w=13.63 l=0.81
X6 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=0 ps=0 w=13.63 l=0.81
X7 VTAIL.t11 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=2.24895 ps=13.96 w=13.63 l=0.81
X8 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=5.3157 ps=28.04 w=13.63 l=0.81
X9 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=5.3157 ps=28.04 w=13.63 l=0.81
X10 VTAIL.t4 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=2.24895 ps=13.96 w=13.63 l=0.81
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=0 ps=0 w=13.63 l=0.81
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=0 ps=0 w=13.63 l=0.81
X13 VDD1.t0 VP.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=5.3157 ps=28.04 w=13.63 l=0.81
X14 VTAIL.t2 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.24895 pd=13.96 as=2.24895 ps=13.96 w=13.63 l=0.81
X15 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3157 pd=28.04 as=2.24895 ps=13.96 w=13.63 l=0.81
R0 VP.n3 VP.t2 477.998
R1 VP.n8 VP.t0 454.33
R2 VP.n12 VP.t1 454.33
R3 VP.n14 VP.t3 454.33
R4 VP.n6 VP.t5 454.33
R5 VP.n4 VP.t4 454.33
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.9044
R14 VP.n9 VP.n7 42.9778
R15 VP.n8 VP.n1 34.3247
R16 VP.n14 VP.n13 34.3247
R17 VP.n6 VP.n5 34.3247
R18 VP.n4 VP.n3 17.9645
R19 VP.n12 VP.n1 13.8763
R20 VP.n13 VP.n12 13.8763
R21 VP.n5 VP.n4 13.8763
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VTAIL.n7 VTAIL.t5 47.1986
R29 VTAIL.n11 VTAIL.t3 47.1984
R30 VTAIL.n2 VTAIL.t9 47.1984
R31 VTAIL.n10 VTAIL.t10 47.1984
R32 VTAIL.n9 VTAIL.n8 45.7459
R33 VTAIL.n6 VTAIL.n5 45.7459
R34 VTAIL.n1 VTAIL.n0 45.7457
R35 VTAIL.n4 VTAIL.n3 45.7457
R36 VTAIL.n6 VTAIL.n4 26.0824
R37 VTAIL.n11 VTAIL.n10 25.0996
R38 VTAIL.n0 VTAIL.t0 1.45318
R39 VTAIL.n0 VTAIL.t4 1.45318
R40 VTAIL.n3 VTAIL.t8 1.45318
R41 VTAIL.n3 VTAIL.t6 1.45318
R42 VTAIL.n8 VTAIL.t7 1.45318
R43 VTAIL.n8 VTAIL.t11 1.45318
R44 VTAIL.n5 VTAIL.t1 1.45318
R45 VTAIL.n5 VTAIL.t2 1.45318
R46 VTAIL.n7 VTAIL.n6 0.983259
R47 VTAIL.n10 VTAIL.n9 0.983259
R48 VTAIL.n4 VTAIL.n2 0.983259
R49 VTAIL.n9 VTAIL.n7 0.961707
R50 VTAIL.n2 VTAIL.n1 0.961707
R51 VTAIL VTAIL.n11 0.679379
R52 VTAIL VTAIL.n1 0.304379
R53 VDD1 VDD1.t3 64.6726
R54 VDD1.n1 VDD1.t5 64.5589
R55 VDD1.n1 VDD1.n0 62.6148
R56 VDD1.n3 VDD1.n2 62.4245
R57 VDD1.n3 VDD1.n1 39.7336
R58 VDD1.n2 VDD1.t1 1.45318
R59 VDD1.n2 VDD1.t0 1.45318
R60 VDD1.n0 VDD1.t4 1.45318
R61 VDD1.n0 VDD1.t2 1.45318
R62 VDD1 VDD1.n3 0.188
R63 B.n97 B.t6 607.331
R64 B.n94 B.t14 607.331
R65 B.n394 B.t10 607.331
R66 B.n392 B.t17 607.331
R67 B.n694 B.n693 585
R68 B.n300 B.n93 585
R69 B.n299 B.n298 585
R70 B.n297 B.n296 585
R71 B.n295 B.n294 585
R72 B.n293 B.n292 585
R73 B.n291 B.n290 585
R74 B.n289 B.n288 585
R75 B.n287 B.n286 585
R76 B.n285 B.n284 585
R77 B.n283 B.n282 585
R78 B.n281 B.n280 585
R79 B.n279 B.n278 585
R80 B.n277 B.n276 585
R81 B.n275 B.n274 585
R82 B.n273 B.n272 585
R83 B.n271 B.n270 585
R84 B.n269 B.n268 585
R85 B.n267 B.n266 585
R86 B.n265 B.n264 585
R87 B.n263 B.n262 585
R88 B.n261 B.n260 585
R89 B.n259 B.n258 585
R90 B.n257 B.n256 585
R91 B.n255 B.n254 585
R92 B.n253 B.n252 585
R93 B.n251 B.n250 585
R94 B.n249 B.n248 585
R95 B.n247 B.n246 585
R96 B.n245 B.n244 585
R97 B.n243 B.n242 585
R98 B.n241 B.n240 585
R99 B.n239 B.n238 585
R100 B.n237 B.n236 585
R101 B.n235 B.n234 585
R102 B.n233 B.n232 585
R103 B.n231 B.n230 585
R104 B.n229 B.n228 585
R105 B.n227 B.n226 585
R106 B.n225 B.n224 585
R107 B.n223 B.n222 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n179 B.n178 585
R130 B.n177 B.n176 585
R131 B.n175 B.n174 585
R132 B.n173 B.n172 585
R133 B.n171 B.n170 585
R134 B.n169 B.n168 585
R135 B.n167 B.n166 585
R136 B.n165 B.n164 585
R137 B.n163 B.n162 585
R138 B.n161 B.n160 585
R139 B.n159 B.n158 585
R140 B.n157 B.n156 585
R141 B.n155 B.n154 585
R142 B.n153 B.n152 585
R143 B.n151 B.n150 585
R144 B.n149 B.n148 585
R145 B.n147 B.n146 585
R146 B.n145 B.n144 585
R147 B.n143 B.n142 585
R148 B.n141 B.n140 585
R149 B.n139 B.n138 585
R150 B.n137 B.n136 585
R151 B.n135 B.n134 585
R152 B.n133 B.n132 585
R153 B.n131 B.n130 585
R154 B.n129 B.n128 585
R155 B.n127 B.n126 585
R156 B.n125 B.n124 585
R157 B.n123 B.n122 585
R158 B.n121 B.n120 585
R159 B.n119 B.n118 585
R160 B.n117 B.n116 585
R161 B.n115 B.n114 585
R162 B.n113 B.n112 585
R163 B.n111 B.n110 585
R164 B.n109 B.n108 585
R165 B.n107 B.n106 585
R166 B.n105 B.n104 585
R167 B.n103 B.n102 585
R168 B.n101 B.n100 585
R169 B.n692 B.n42 585
R170 B.n697 B.n42 585
R171 B.n691 B.n41 585
R172 B.n698 B.n41 585
R173 B.n690 B.n689 585
R174 B.n689 B.n37 585
R175 B.n688 B.n36 585
R176 B.n704 B.n36 585
R177 B.n687 B.n35 585
R178 B.n705 B.n35 585
R179 B.n686 B.n34 585
R180 B.n706 B.n34 585
R181 B.n685 B.n684 585
R182 B.n684 B.n30 585
R183 B.n683 B.n29 585
R184 B.n712 B.n29 585
R185 B.n682 B.n28 585
R186 B.n713 B.n28 585
R187 B.n681 B.n27 585
R188 B.n714 B.n27 585
R189 B.n680 B.n679 585
R190 B.n679 B.n23 585
R191 B.n678 B.n22 585
R192 B.n720 B.n22 585
R193 B.n677 B.n21 585
R194 B.n721 B.n21 585
R195 B.n676 B.n20 585
R196 B.n722 B.n20 585
R197 B.n675 B.n674 585
R198 B.n674 B.n19 585
R199 B.n673 B.n15 585
R200 B.n728 B.n15 585
R201 B.n672 B.n14 585
R202 B.n729 B.n14 585
R203 B.n671 B.n13 585
R204 B.n730 B.n13 585
R205 B.n670 B.n669 585
R206 B.n669 B.n12 585
R207 B.n668 B.n667 585
R208 B.n668 B.n8 585
R209 B.n666 B.n7 585
R210 B.n737 B.n7 585
R211 B.n665 B.n6 585
R212 B.n738 B.n6 585
R213 B.n664 B.n5 585
R214 B.n739 B.n5 585
R215 B.n663 B.n662 585
R216 B.n662 B.n4 585
R217 B.n661 B.n301 585
R218 B.n661 B.n660 585
R219 B.n650 B.n302 585
R220 B.n653 B.n302 585
R221 B.n652 B.n651 585
R222 B.n654 B.n652 585
R223 B.n649 B.n307 585
R224 B.n307 B.n306 585
R225 B.n648 B.n647 585
R226 B.n647 B.n646 585
R227 B.n309 B.n308 585
R228 B.n639 B.n309 585
R229 B.n638 B.n637 585
R230 B.n640 B.n638 585
R231 B.n636 B.n314 585
R232 B.n314 B.n313 585
R233 B.n635 B.n634 585
R234 B.n634 B.n633 585
R235 B.n316 B.n315 585
R236 B.n317 B.n316 585
R237 B.n626 B.n625 585
R238 B.n627 B.n626 585
R239 B.n624 B.n322 585
R240 B.n322 B.n321 585
R241 B.n623 B.n622 585
R242 B.n622 B.n621 585
R243 B.n324 B.n323 585
R244 B.n325 B.n324 585
R245 B.n614 B.n613 585
R246 B.n615 B.n614 585
R247 B.n612 B.n329 585
R248 B.n333 B.n329 585
R249 B.n611 B.n610 585
R250 B.n610 B.n609 585
R251 B.n331 B.n330 585
R252 B.n332 B.n331 585
R253 B.n602 B.n601 585
R254 B.n603 B.n602 585
R255 B.n600 B.n338 585
R256 B.n338 B.n337 585
R257 B.n595 B.n594 585
R258 B.n593 B.n391 585
R259 B.n592 B.n390 585
R260 B.n597 B.n390 585
R261 B.n591 B.n590 585
R262 B.n589 B.n588 585
R263 B.n587 B.n586 585
R264 B.n585 B.n584 585
R265 B.n583 B.n582 585
R266 B.n581 B.n580 585
R267 B.n579 B.n578 585
R268 B.n577 B.n576 585
R269 B.n575 B.n574 585
R270 B.n573 B.n572 585
R271 B.n571 B.n570 585
R272 B.n569 B.n568 585
R273 B.n567 B.n566 585
R274 B.n565 B.n564 585
R275 B.n563 B.n562 585
R276 B.n561 B.n560 585
R277 B.n559 B.n558 585
R278 B.n557 B.n556 585
R279 B.n555 B.n554 585
R280 B.n553 B.n552 585
R281 B.n551 B.n550 585
R282 B.n549 B.n548 585
R283 B.n547 B.n546 585
R284 B.n545 B.n544 585
R285 B.n543 B.n542 585
R286 B.n541 B.n540 585
R287 B.n539 B.n538 585
R288 B.n537 B.n536 585
R289 B.n535 B.n534 585
R290 B.n533 B.n532 585
R291 B.n531 B.n530 585
R292 B.n529 B.n528 585
R293 B.n527 B.n526 585
R294 B.n525 B.n524 585
R295 B.n523 B.n522 585
R296 B.n521 B.n520 585
R297 B.n519 B.n518 585
R298 B.n517 B.n516 585
R299 B.n515 B.n514 585
R300 B.n513 B.n512 585
R301 B.n511 B.n510 585
R302 B.n509 B.n508 585
R303 B.n507 B.n506 585
R304 B.n504 B.n503 585
R305 B.n502 B.n501 585
R306 B.n500 B.n499 585
R307 B.n498 B.n497 585
R308 B.n496 B.n495 585
R309 B.n494 B.n493 585
R310 B.n492 B.n491 585
R311 B.n490 B.n489 585
R312 B.n488 B.n487 585
R313 B.n486 B.n485 585
R314 B.n483 B.n482 585
R315 B.n481 B.n480 585
R316 B.n479 B.n478 585
R317 B.n477 B.n476 585
R318 B.n475 B.n474 585
R319 B.n473 B.n472 585
R320 B.n471 B.n470 585
R321 B.n469 B.n468 585
R322 B.n467 B.n466 585
R323 B.n465 B.n464 585
R324 B.n463 B.n462 585
R325 B.n461 B.n460 585
R326 B.n459 B.n458 585
R327 B.n457 B.n456 585
R328 B.n455 B.n454 585
R329 B.n453 B.n452 585
R330 B.n451 B.n450 585
R331 B.n449 B.n448 585
R332 B.n447 B.n446 585
R333 B.n445 B.n444 585
R334 B.n443 B.n442 585
R335 B.n441 B.n440 585
R336 B.n439 B.n438 585
R337 B.n437 B.n436 585
R338 B.n435 B.n434 585
R339 B.n433 B.n432 585
R340 B.n431 B.n430 585
R341 B.n429 B.n428 585
R342 B.n427 B.n426 585
R343 B.n425 B.n424 585
R344 B.n423 B.n422 585
R345 B.n421 B.n420 585
R346 B.n419 B.n418 585
R347 B.n417 B.n416 585
R348 B.n415 B.n414 585
R349 B.n413 B.n412 585
R350 B.n411 B.n410 585
R351 B.n409 B.n408 585
R352 B.n407 B.n406 585
R353 B.n405 B.n404 585
R354 B.n403 B.n402 585
R355 B.n401 B.n400 585
R356 B.n399 B.n398 585
R357 B.n397 B.n396 585
R358 B.n340 B.n339 585
R359 B.n599 B.n598 585
R360 B.n598 B.n597 585
R361 B.n336 B.n335 585
R362 B.n337 B.n336 585
R363 B.n605 B.n604 585
R364 B.n604 B.n603 585
R365 B.n606 B.n334 585
R366 B.n334 B.n332 585
R367 B.n608 B.n607 585
R368 B.n609 B.n608 585
R369 B.n328 B.n327 585
R370 B.n333 B.n328 585
R371 B.n617 B.n616 585
R372 B.n616 B.n615 585
R373 B.n618 B.n326 585
R374 B.n326 B.n325 585
R375 B.n620 B.n619 585
R376 B.n621 B.n620 585
R377 B.n320 B.n319 585
R378 B.n321 B.n320 585
R379 B.n629 B.n628 585
R380 B.n628 B.n627 585
R381 B.n630 B.n318 585
R382 B.n318 B.n317 585
R383 B.n632 B.n631 585
R384 B.n633 B.n632 585
R385 B.n312 B.n311 585
R386 B.n313 B.n312 585
R387 B.n642 B.n641 585
R388 B.n641 B.n640 585
R389 B.n643 B.n310 585
R390 B.n639 B.n310 585
R391 B.n645 B.n644 585
R392 B.n646 B.n645 585
R393 B.n305 B.n304 585
R394 B.n306 B.n305 585
R395 B.n656 B.n655 585
R396 B.n655 B.n654 585
R397 B.n657 B.n303 585
R398 B.n653 B.n303 585
R399 B.n659 B.n658 585
R400 B.n660 B.n659 585
R401 B.n3 B.n0 585
R402 B.n4 B.n3 585
R403 B.n736 B.n1 585
R404 B.n737 B.n736 585
R405 B.n735 B.n734 585
R406 B.n735 B.n8 585
R407 B.n733 B.n9 585
R408 B.n12 B.n9 585
R409 B.n732 B.n731 585
R410 B.n731 B.n730 585
R411 B.n11 B.n10 585
R412 B.n729 B.n11 585
R413 B.n727 B.n726 585
R414 B.n728 B.n727 585
R415 B.n725 B.n16 585
R416 B.n19 B.n16 585
R417 B.n724 B.n723 585
R418 B.n723 B.n722 585
R419 B.n18 B.n17 585
R420 B.n721 B.n18 585
R421 B.n719 B.n718 585
R422 B.n720 B.n719 585
R423 B.n717 B.n24 585
R424 B.n24 B.n23 585
R425 B.n716 B.n715 585
R426 B.n715 B.n714 585
R427 B.n26 B.n25 585
R428 B.n713 B.n26 585
R429 B.n711 B.n710 585
R430 B.n712 B.n711 585
R431 B.n709 B.n31 585
R432 B.n31 B.n30 585
R433 B.n708 B.n707 585
R434 B.n707 B.n706 585
R435 B.n33 B.n32 585
R436 B.n705 B.n33 585
R437 B.n703 B.n702 585
R438 B.n704 B.n703 585
R439 B.n701 B.n38 585
R440 B.n38 B.n37 585
R441 B.n700 B.n699 585
R442 B.n699 B.n698 585
R443 B.n40 B.n39 585
R444 B.n697 B.n40 585
R445 B.n740 B.n739 585
R446 B.n738 B.n2 585
R447 B.n100 B.n40 535.745
R448 B.n694 B.n42 535.745
R449 B.n598 B.n338 535.745
R450 B.n595 B.n336 535.745
R451 B.n696 B.n695 256.663
R452 B.n696 B.n92 256.663
R453 B.n696 B.n91 256.663
R454 B.n696 B.n90 256.663
R455 B.n696 B.n89 256.663
R456 B.n696 B.n88 256.663
R457 B.n696 B.n87 256.663
R458 B.n696 B.n86 256.663
R459 B.n696 B.n85 256.663
R460 B.n696 B.n84 256.663
R461 B.n696 B.n83 256.663
R462 B.n696 B.n82 256.663
R463 B.n696 B.n81 256.663
R464 B.n696 B.n80 256.663
R465 B.n696 B.n79 256.663
R466 B.n696 B.n78 256.663
R467 B.n696 B.n77 256.663
R468 B.n696 B.n76 256.663
R469 B.n696 B.n75 256.663
R470 B.n696 B.n74 256.663
R471 B.n696 B.n73 256.663
R472 B.n696 B.n72 256.663
R473 B.n696 B.n71 256.663
R474 B.n696 B.n70 256.663
R475 B.n696 B.n69 256.663
R476 B.n696 B.n68 256.663
R477 B.n696 B.n67 256.663
R478 B.n696 B.n66 256.663
R479 B.n696 B.n65 256.663
R480 B.n696 B.n64 256.663
R481 B.n696 B.n63 256.663
R482 B.n696 B.n62 256.663
R483 B.n696 B.n61 256.663
R484 B.n696 B.n60 256.663
R485 B.n696 B.n59 256.663
R486 B.n696 B.n58 256.663
R487 B.n696 B.n57 256.663
R488 B.n696 B.n56 256.663
R489 B.n696 B.n55 256.663
R490 B.n696 B.n54 256.663
R491 B.n696 B.n53 256.663
R492 B.n696 B.n52 256.663
R493 B.n696 B.n51 256.663
R494 B.n696 B.n50 256.663
R495 B.n696 B.n49 256.663
R496 B.n696 B.n48 256.663
R497 B.n696 B.n47 256.663
R498 B.n696 B.n46 256.663
R499 B.n696 B.n45 256.663
R500 B.n696 B.n44 256.663
R501 B.n696 B.n43 256.663
R502 B.n597 B.n596 256.663
R503 B.n597 B.n341 256.663
R504 B.n597 B.n342 256.663
R505 B.n597 B.n343 256.663
R506 B.n597 B.n344 256.663
R507 B.n597 B.n345 256.663
R508 B.n597 B.n346 256.663
R509 B.n597 B.n347 256.663
R510 B.n597 B.n348 256.663
R511 B.n597 B.n349 256.663
R512 B.n597 B.n350 256.663
R513 B.n597 B.n351 256.663
R514 B.n597 B.n352 256.663
R515 B.n597 B.n353 256.663
R516 B.n597 B.n354 256.663
R517 B.n597 B.n355 256.663
R518 B.n597 B.n356 256.663
R519 B.n597 B.n357 256.663
R520 B.n597 B.n358 256.663
R521 B.n597 B.n359 256.663
R522 B.n597 B.n360 256.663
R523 B.n597 B.n361 256.663
R524 B.n597 B.n362 256.663
R525 B.n597 B.n363 256.663
R526 B.n597 B.n364 256.663
R527 B.n597 B.n365 256.663
R528 B.n597 B.n366 256.663
R529 B.n597 B.n367 256.663
R530 B.n597 B.n368 256.663
R531 B.n597 B.n369 256.663
R532 B.n597 B.n370 256.663
R533 B.n597 B.n371 256.663
R534 B.n597 B.n372 256.663
R535 B.n597 B.n373 256.663
R536 B.n597 B.n374 256.663
R537 B.n597 B.n375 256.663
R538 B.n597 B.n376 256.663
R539 B.n597 B.n377 256.663
R540 B.n597 B.n378 256.663
R541 B.n597 B.n379 256.663
R542 B.n597 B.n380 256.663
R543 B.n597 B.n381 256.663
R544 B.n597 B.n382 256.663
R545 B.n597 B.n383 256.663
R546 B.n597 B.n384 256.663
R547 B.n597 B.n385 256.663
R548 B.n597 B.n386 256.663
R549 B.n597 B.n387 256.663
R550 B.n597 B.n388 256.663
R551 B.n597 B.n389 256.663
R552 B.n742 B.n741 256.663
R553 B.n104 B.n103 163.367
R554 B.n108 B.n107 163.367
R555 B.n112 B.n111 163.367
R556 B.n116 B.n115 163.367
R557 B.n120 B.n119 163.367
R558 B.n124 B.n123 163.367
R559 B.n128 B.n127 163.367
R560 B.n132 B.n131 163.367
R561 B.n136 B.n135 163.367
R562 B.n140 B.n139 163.367
R563 B.n144 B.n143 163.367
R564 B.n148 B.n147 163.367
R565 B.n152 B.n151 163.367
R566 B.n156 B.n155 163.367
R567 B.n160 B.n159 163.367
R568 B.n164 B.n163 163.367
R569 B.n168 B.n167 163.367
R570 B.n172 B.n171 163.367
R571 B.n176 B.n175 163.367
R572 B.n180 B.n179 163.367
R573 B.n184 B.n183 163.367
R574 B.n188 B.n187 163.367
R575 B.n192 B.n191 163.367
R576 B.n196 B.n195 163.367
R577 B.n200 B.n199 163.367
R578 B.n204 B.n203 163.367
R579 B.n208 B.n207 163.367
R580 B.n212 B.n211 163.367
R581 B.n216 B.n215 163.367
R582 B.n220 B.n219 163.367
R583 B.n224 B.n223 163.367
R584 B.n228 B.n227 163.367
R585 B.n232 B.n231 163.367
R586 B.n236 B.n235 163.367
R587 B.n240 B.n239 163.367
R588 B.n244 B.n243 163.367
R589 B.n248 B.n247 163.367
R590 B.n252 B.n251 163.367
R591 B.n256 B.n255 163.367
R592 B.n260 B.n259 163.367
R593 B.n264 B.n263 163.367
R594 B.n268 B.n267 163.367
R595 B.n272 B.n271 163.367
R596 B.n276 B.n275 163.367
R597 B.n280 B.n279 163.367
R598 B.n284 B.n283 163.367
R599 B.n288 B.n287 163.367
R600 B.n292 B.n291 163.367
R601 B.n296 B.n295 163.367
R602 B.n298 B.n93 163.367
R603 B.n602 B.n338 163.367
R604 B.n602 B.n331 163.367
R605 B.n610 B.n331 163.367
R606 B.n610 B.n329 163.367
R607 B.n614 B.n329 163.367
R608 B.n614 B.n324 163.367
R609 B.n622 B.n324 163.367
R610 B.n622 B.n322 163.367
R611 B.n626 B.n322 163.367
R612 B.n626 B.n316 163.367
R613 B.n634 B.n316 163.367
R614 B.n634 B.n314 163.367
R615 B.n638 B.n314 163.367
R616 B.n638 B.n309 163.367
R617 B.n647 B.n309 163.367
R618 B.n647 B.n307 163.367
R619 B.n652 B.n307 163.367
R620 B.n652 B.n302 163.367
R621 B.n661 B.n302 163.367
R622 B.n662 B.n661 163.367
R623 B.n662 B.n5 163.367
R624 B.n6 B.n5 163.367
R625 B.n7 B.n6 163.367
R626 B.n668 B.n7 163.367
R627 B.n669 B.n668 163.367
R628 B.n669 B.n13 163.367
R629 B.n14 B.n13 163.367
R630 B.n15 B.n14 163.367
R631 B.n674 B.n15 163.367
R632 B.n674 B.n20 163.367
R633 B.n21 B.n20 163.367
R634 B.n22 B.n21 163.367
R635 B.n679 B.n22 163.367
R636 B.n679 B.n27 163.367
R637 B.n28 B.n27 163.367
R638 B.n29 B.n28 163.367
R639 B.n684 B.n29 163.367
R640 B.n684 B.n34 163.367
R641 B.n35 B.n34 163.367
R642 B.n36 B.n35 163.367
R643 B.n689 B.n36 163.367
R644 B.n689 B.n41 163.367
R645 B.n42 B.n41 163.367
R646 B.n391 B.n390 163.367
R647 B.n590 B.n390 163.367
R648 B.n588 B.n587 163.367
R649 B.n584 B.n583 163.367
R650 B.n580 B.n579 163.367
R651 B.n576 B.n575 163.367
R652 B.n572 B.n571 163.367
R653 B.n568 B.n567 163.367
R654 B.n564 B.n563 163.367
R655 B.n560 B.n559 163.367
R656 B.n556 B.n555 163.367
R657 B.n552 B.n551 163.367
R658 B.n548 B.n547 163.367
R659 B.n544 B.n543 163.367
R660 B.n540 B.n539 163.367
R661 B.n536 B.n535 163.367
R662 B.n532 B.n531 163.367
R663 B.n528 B.n527 163.367
R664 B.n524 B.n523 163.367
R665 B.n520 B.n519 163.367
R666 B.n516 B.n515 163.367
R667 B.n512 B.n511 163.367
R668 B.n508 B.n507 163.367
R669 B.n503 B.n502 163.367
R670 B.n499 B.n498 163.367
R671 B.n495 B.n494 163.367
R672 B.n491 B.n490 163.367
R673 B.n487 B.n486 163.367
R674 B.n482 B.n481 163.367
R675 B.n478 B.n477 163.367
R676 B.n474 B.n473 163.367
R677 B.n470 B.n469 163.367
R678 B.n466 B.n465 163.367
R679 B.n462 B.n461 163.367
R680 B.n458 B.n457 163.367
R681 B.n454 B.n453 163.367
R682 B.n450 B.n449 163.367
R683 B.n446 B.n445 163.367
R684 B.n442 B.n441 163.367
R685 B.n438 B.n437 163.367
R686 B.n434 B.n433 163.367
R687 B.n430 B.n429 163.367
R688 B.n426 B.n425 163.367
R689 B.n422 B.n421 163.367
R690 B.n418 B.n417 163.367
R691 B.n414 B.n413 163.367
R692 B.n410 B.n409 163.367
R693 B.n406 B.n405 163.367
R694 B.n402 B.n401 163.367
R695 B.n398 B.n397 163.367
R696 B.n598 B.n340 163.367
R697 B.n604 B.n336 163.367
R698 B.n604 B.n334 163.367
R699 B.n608 B.n334 163.367
R700 B.n608 B.n328 163.367
R701 B.n616 B.n328 163.367
R702 B.n616 B.n326 163.367
R703 B.n620 B.n326 163.367
R704 B.n620 B.n320 163.367
R705 B.n628 B.n320 163.367
R706 B.n628 B.n318 163.367
R707 B.n632 B.n318 163.367
R708 B.n632 B.n312 163.367
R709 B.n641 B.n312 163.367
R710 B.n641 B.n310 163.367
R711 B.n645 B.n310 163.367
R712 B.n645 B.n305 163.367
R713 B.n655 B.n305 163.367
R714 B.n655 B.n303 163.367
R715 B.n659 B.n303 163.367
R716 B.n659 B.n3 163.367
R717 B.n740 B.n3 163.367
R718 B.n736 B.n2 163.367
R719 B.n736 B.n735 163.367
R720 B.n735 B.n9 163.367
R721 B.n731 B.n9 163.367
R722 B.n731 B.n11 163.367
R723 B.n727 B.n11 163.367
R724 B.n727 B.n16 163.367
R725 B.n723 B.n16 163.367
R726 B.n723 B.n18 163.367
R727 B.n719 B.n18 163.367
R728 B.n719 B.n24 163.367
R729 B.n715 B.n24 163.367
R730 B.n715 B.n26 163.367
R731 B.n711 B.n26 163.367
R732 B.n711 B.n31 163.367
R733 B.n707 B.n31 163.367
R734 B.n707 B.n33 163.367
R735 B.n703 B.n33 163.367
R736 B.n703 B.n38 163.367
R737 B.n699 B.n38 163.367
R738 B.n699 B.n40 163.367
R739 B.n94 B.t15 90.286
R740 B.n394 B.t13 90.286
R741 B.n97 B.t8 90.2683
R742 B.n392 B.t19 90.2683
R743 B.n597 B.n337 72.7326
R744 B.n697 B.n696 72.7326
R745 B.n100 B.n43 71.676
R746 B.n104 B.n44 71.676
R747 B.n108 B.n45 71.676
R748 B.n112 B.n46 71.676
R749 B.n116 B.n47 71.676
R750 B.n120 B.n48 71.676
R751 B.n124 B.n49 71.676
R752 B.n128 B.n50 71.676
R753 B.n132 B.n51 71.676
R754 B.n136 B.n52 71.676
R755 B.n140 B.n53 71.676
R756 B.n144 B.n54 71.676
R757 B.n148 B.n55 71.676
R758 B.n152 B.n56 71.676
R759 B.n156 B.n57 71.676
R760 B.n160 B.n58 71.676
R761 B.n164 B.n59 71.676
R762 B.n168 B.n60 71.676
R763 B.n172 B.n61 71.676
R764 B.n176 B.n62 71.676
R765 B.n180 B.n63 71.676
R766 B.n184 B.n64 71.676
R767 B.n188 B.n65 71.676
R768 B.n192 B.n66 71.676
R769 B.n196 B.n67 71.676
R770 B.n200 B.n68 71.676
R771 B.n204 B.n69 71.676
R772 B.n208 B.n70 71.676
R773 B.n212 B.n71 71.676
R774 B.n216 B.n72 71.676
R775 B.n220 B.n73 71.676
R776 B.n224 B.n74 71.676
R777 B.n228 B.n75 71.676
R778 B.n232 B.n76 71.676
R779 B.n236 B.n77 71.676
R780 B.n240 B.n78 71.676
R781 B.n244 B.n79 71.676
R782 B.n248 B.n80 71.676
R783 B.n252 B.n81 71.676
R784 B.n256 B.n82 71.676
R785 B.n260 B.n83 71.676
R786 B.n264 B.n84 71.676
R787 B.n268 B.n85 71.676
R788 B.n272 B.n86 71.676
R789 B.n276 B.n87 71.676
R790 B.n280 B.n88 71.676
R791 B.n284 B.n89 71.676
R792 B.n288 B.n90 71.676
R793 B.n292 B.n91 71.676
R794 B.n296 B.n92 71.676
R795 B.n695 B.n93 71.676
R796 B.n695 B.n694 71.676
R797 B.n298 B.n92 71.676
R798 B.n295 B.n91 71.676
R799 B.n291 B.n90 71.676
R800 B.n287 B.n89 71.676
R801 B.n283 B.n88 71.676
R802 B.n279 B.n87 71.676
R803 B.n275 B.n86 71.676
R804 B.n271 B.n85 71.676
R805 B.n267 B.n84 71.676
R806 B.n263 B.n83 71.676
R807 B.n259 B.n82 71.676
R808 B.n255 B.n81 71.676
R809 B.n251 B.n80 71.676
R810 B.n247 B.n79 71.676
R811 B.n243 B.n78 71.676
R812 B.n239 B.n77 71.676
R813 B.n235 B.n76 71.676
R814 B.n231 B.n75 71.676
R815 B.n227 B.n74 71.676
R816 B.n223 B.n73 71.676
R817 B.n219 B.n72 71.676
R818 B.n215 B.n71 71.676
R819 B.n211 B.n70 71.676
R820 B.n207 B.n69 71.676
R821 B.n203 B.n68 71.676
R822 B.n199 B.n67 71.676
R823 B.n195 B.n66 71.676
R824 B.n191 B.n65 71.676
R825 B.n187 B.n64 71.676
R826 B.n183 B.n63 71.676
R827 B.n179 B.n62 71.676
R828 B.n175 B.n61 71.676
R829 B.n171 B.n60 71.676
R830 B.n167 B.n59 71.676
R831 B.n163 B.n58 71.676
R832 B.n159 B.n57 71.676
R833 B.n155 B.n56 71.676
R834 B.n151 B.n55 71.676
R835 B.n147 B.n54 71.676
R836 B.n143 B.n53 71.676
R837 B.n139 B.n52 71.676
R838 B.n135 B.n51 71.676
R839 B.n131 B.n50 71.676
R840 B.n127 B.n49 71.676
R841 B.n123 B.n48 71.676
R842 B.n119 B.n47 71.676
R843 B.n115 B.n46 71.676
R844 B.n111 B.n45 71.676
R845 B.n107 B.n44 71.676
R846 B.n103 B.n43 71.676
R847 B.n596 B.n595 71.676
R848 B.n590 B.n341 71.676
R849 B.n587 B.n342 71.676
R850 B.n583 B.n343 71.676
R851 B.n579 B.n344 71.676
R852 B.n575 B.n345 71.676
R853 B.n571 B.n346 71.676
R854 B.n567 B.n347 71.676
R855 B.n563 B.n348 71.676
R856 B.n559 B.n349 71.676
R857 B.n555 B.n350 71.676
R858 B.n551 B.n351 71.676
R859 B.n547 B.n352 71.676
R860 B.n543 B.n353 71.676
R861 B.n539 B.n354 71.676
R862 B.n535 B.n355 71.676
R863 B.n531 B.n356 71.676
R864 B.n527 B.n357 71.676
R865 B.n523 B.n358 71.676
R866 B.n519 B.n359 71.676
R867 B.n515 B.n360 71.676
R868 B.n511 B.n361 71.676
R869 B.n507 B.n362 71.676
R870 B.n502 B.n363 71.676
R871 B.n498 B.n364 71.676
R872 B.n494 B.n365 71.676
R873 B.n490 B.n366 71.676
R874 B.n486 B.n367 71.676
R875 B.n481 B.n368 71.676
R876 B.n477 B.n369 71.676
R877 B.n473 B.n370 71.676
R878 B.n469 B.n371 71.676
R879 B.n465 B.n372 71.676
R880 B.n461 B.n373 71.676
R881 B.n457 B.n374 71.676
R882 B.n453 B.n375 71.676
R883 B.n449 B.n376 71.676
R884 B.n445 B.n377 71.676
R885 B.n441 B.n378 71.676
R886 B.n437 B.n379 71.676
R887 B.n433 B.n380 71.676
R888 B.n429 B.n381 71.676
R889 B.n425 B.n382 71.676
R890 B.n421 B.n383 71.676
R891 B.n417 B.n384 71.676
R892 B.n413 B.n385 71.676
R893 B.n409 B.n386 71.676
R894 B.n405 B.n387 71.676
R895 B.n401 B.n388 71.676
R896 B.n397 B.n389 71.676
R897 B.n596 B.n391 71.676
R898 B.n588 B.n341 71.676
R899 B.n584 B.n342 71.676
R900 B.n580 B.n343 71.676
R901 B.n576 B.n344 71.676
R902 B.n572 B.n345 71.676
R903 B.n568 B.n346 71.676
R904 B.n564 B.n347 71.676
R905 B.n560 B.n348 71.676
R906 B.n556 B.n349 71.676
R907 B.n552 B.n350 71.676
R908 B.n548 B.n351 71.676
R909 B.n544 B.n352 71.676
R910 B.n540 B.n353 71.676
R911 B.n536 B.n354 71.676
R912 B.n532 B.n355 71.676
R913 B.n528 B.n356 71.676
R914 B.n524 B.n357 71.676
R915 B.n520 B.n358 71.676
R916 B.n516 B.n359 71.676
R917 B.n512 B.n360 71.676
R918 B.n508 B.n361 71.676
R919 B.n503 B.n362 71.676
R920 B.n499 B.n363 71.676
R921 B.n495 B.n364 71.676
R922 B.n491 B.n365 71.676
R923 B.n487 B.n366 71.676
R924 B.n482 B.n367 71.676
R925 B.n478 B.n368 71.676
R926 B.n474 B.n369 71.676
R927 B.n470 B.n370 71.676
R928 B.n466 B.n371 71.676
R929 B.n462 B.n372 71.676
R930 B.n458 B.n373 71.676
R931 B.n454 B.n374 71.676
R932 B.n450 B.n375 71.676
R933 B.n446 B.n376 71.676
R934 B.n442 B.n377 71.676
R935 B.n438 B.n378 71.676
R936 B.n434 B.n379 71.676
R937 B.n430 B.n380 71.676
R938 B.n426 B.n381 71.676
R939 B.n422 B.n382 71.676
R940 B.n418 B.n383 71.676
R941 B.n414 B.n384 71.676
R942 B.n410 B.n385 71.676
R943 B.n406 B.n386 71.676
R944 B.n402 B.n387 71.676
R945 B.n398 B.n388 71.676
R946 B.n389 B.n340 71.676
R947 B.n741 B.n740 71.676
R948 B.n741 B.n2 71.676
R949 B.n95 B.t16 68.1769
R950 B.n395 B.t12 68.1769
R951 B.n98 B.t9 68.1592
R952 B.n393 B.t18 68.1592
R953 B.n99 B.n98 59.5399
R954 B.n96 B.n95 59.5399
R955 B.n484 B.n395 59.5399
R956 B.n505 B.n393 59.5399
R957 B.n603 B.n337 39.5668
R958 B.n603 B.n332 39.5668
R959 B.n609 B.n332 39.5668
R960 B.n609 B.n333 39.5668
R961 B.n615 B.n325 39.5668
R962 B.n621 B.n325 39.5668
R963 B.n621 B.n321 39.5668
R964 B.n627 B.n321 39.5668
R965 B.n627 B.n317 39.5668
R966 B.n633 B.n317 39.5668
R967 B.n640 B.n313 39.5668
R968 B.n640 B.n639 39.5668
R969 B.n646 B.n306 39.5668
R970 B.n654 B.n306 39.5668
R971 B.n654 B.n653 39.5668
R972 B.n660 B.n4 39.5668
R973 B.n739 B.n4 39.5668
R974 B.n739 B.n738 39.5668
R975 B.n738 B.n737 39.5668
R976 B.n737 B.n8 39.5668
R977 B.n730 B.n12 39.5668
R978 B.n730 B.n729 39.5668
R979 B.n729 B.n728 39.5668
R980 B.n722 B.n19 39.5668
R981 B.n722 B.n721 39.5668
R982 B.n720 B.n23 39.5668
R983 B.n714 B.n23 39.5668
R984 B.n714 B.n713 39.5668
R985 B.n713 B.n712 39.5668
R986 B.n712 B.n30 39.5668
R987 B.n706 B.n30 39.5668
R988 B.n705 B.n704 39.5668
R989 B.n704 B.n37 39.5668
R990 B.n698 B.n37 39.5668
R991 B.n698 B.n697 39.5668
R992 B.n333 B.t11 37.8212
R993 B.t7 B.n705 37.8212
R994 B.n594 B.n335 34.8103
R995 B.n600 B.n599 34.8103
R996 B.n693 B.n692 34.8103
R997 B.n101 B.n39 34.8103
R998 B.n639 B.t2 34.33
R999 B.n19 B.t4 34.33
R1000 B.n660 B.t5 30.8389
R1001 B.t0 B.n8 30.8389
R1002 B.n98 B.n97 22.1096
R1003 B.n95 B.n94 22.1096
R1004 B.n395 B.n394 22.1096
R1005 B.n393 B.n392 22.1096
R1006 B.n633 B.t1 20.3655
R1007 B.t3 B.n720 20.3655
R1008 B.t1 B.n313 19.2018
R1009 B.n721 B.t3 19.2018
R1010 B B.n742 18.0485
R1011 B.n605 B.n335 10.6151
R1012 B.n606 B.n605 10.6151
R1013 B.n607 B.n606 10.6151
R1014 B.n607 B.n327 10.6151
R1015 B.n617 B.n327 10.6151
R1016 B.n618 B.n617 10.6151
R1017 B.n619 B.n618 10.6151
R1018 B.n619 B.n319 10.6151
R1019 B.n629 B.n319 10.6151
R1020 B.n630 B.n629 10.6151
R1021 B.n631 B.n630 10.6151
R1022 B.n631 B.n311 10.6151
R1023 B.n642 B.n311 10.6151
R1024 B.n643 B.n642 10.6151
R1025 B.n644 B.n643 10.6151
R1026 B.n644 B.n304 10.6151
R1027 B.n656 B.n304 10.6151
R1028 B.n657 B.n656 10.6151
R1029 B.n658 B.n657 10.6151
R1030 B.n658 B.n0 10.6151
R1031 B.n594 B.n593 10.6151
R1032 B.n593 B.n592 10.6151
R1033 B.n592 B.n591 10.6151
R1034 B.n591 B.n589 10.6151
R1035 B.n589 B.n586 10.6151
R1036 B.n586 B.n585 10.6151
R1037 B.n585 B.n582 10.6151
R1038 B.n582 B.n581 10.6151
R1039 B.n581 B.n578 10.6151
R1040 B.n578 B.n577 10.6151
R1041 B.n577 B.n574 10.6151
R1042 B.n574 B.n573 10.6151
R1043 B.n573 B.n570 10.6151
R1044 B.n570 B.n569 10.6151
R1045 B.n569 B.n566 10.6151
R1046 B.n566 B.n565 10.6151
R1047 B.n565 B.n562 10.6151
R1048 B.n562 B.n561 10.6151
R1049 B.n561 B.n558 10.6151
R1050 B.n558 B.n557 10.6151
R1051 B.n557 B.n554 10.6151
R1052 B.n554 B.n553 10.6151
R1053 B.n553 B.n550 10.6151
R1054 B.n550 B.n549 10.6151
R1055 B.n549 B.n546 10.6151
R1056 B.n546 B.n545 10.6151
R1057 B.n545 B.n542 10.6151
R1058 B.n542 B.n541 10.6151
R1059 B.n541 B.n538 10.6151
R1060 B.n538 B.n537 10.6151
R1061 B.n537 B.n534 10.6151
R1062 B.n534 B.n533 10.6151
R1063 B.n533 B.n530 10.6151
R1064 B.n530 B.n529 10.6151
R1065 B.n529 B.n526 10.6151
R1066 B.n526 B.n525 10.6151
R1067 B.n525 B.n522 10.6151
R1068 B.n522 B.n521 10.6151
R1069 B.n521 B.n518 10.6151
R1070 B.n518 B.n517 10.6151
R1071 B.n517 B.n514 10.6151
R1072 B.n514 B.n513 10.6151
R1073 B.n513 B.n510 10.6151
R1074 B.n510 B.n509 10.6151
R1075 B.n509 B.n506 10.6151
R1076 B.n504 B.n501 10.6151
R1077 B.n501 B.n500 10.6151
R1078 B.n500 B.n497 10.6151
R1079 B.n497 B.n496 10.6151
R1080 B.n496 B.n493 10.6151
R1081 B.n493 B.n492 10.6151
R1082 B.n492 B.n489 10.6151
R1083 B.n489 B.n488 10.6151
R1084 B.n488 B.n485 10.6151
R1085 B.n483 B.n480 10.6151
R1086 B.n480 B.n479 10.6151
R1087 B.n479 B.n476 10.6151
R1088 B.n476 B.n475 10.6151
R1089 B.n475 B.n472 10.6151
R1090 B.n472 B.n471 10.6151
R1091 B.n471 B.n468 10.6151
R1092 B.n468 B.n467 10.6151
R1093 B.n467 B.n464 10.6151
R1094 B.n464 B.n463 10.6151
R1095 B.n463 B.n460 10.6151
R1096 B.n460 B.n459 10.6151
R1097 B.n459 B.n456 10.6151
R1098 B.n456 B.n455 10.6151
R1099 B.n455 B.n452 10.6151
R1100 B.n452 B.n451 10.6151
R1101 B.n451 B.n448 10.6151
R1102 B.n448 B.n447 10.6151
R1103 B.n447 B.n444 10.6151
R1104 B.n444 B.n443 10.6151
R1105 B.n443 B.n440 10.6151
R1106 B.n440 B.n439 10.6151
R1107 B.n439 B.n436 10.6151
R1108 B.n436 B.n435 10.6151
R1109 B.n435 B.n432 10.6151
R1110 B.n432 B.n431 10.6151
R1111 B.n431 B.n428 10.6151
R1112 B.n428 B.n427 10.6151
R1113 B.n427 B.n424 10.6151
R1114 B.n424 B.n423 10.6151
R1115 B.n423 B.n420 10.6151
R1116 B.n420 B.n419 10.6151
R1117 B.n419 B.n416 10.6151
R1118 B.n416 B.n415 10.6151
R1119 B.n415 B.n412 10.6151
R1120 B.n412 B.n411 10.6151
R1121 B.n411 B.n408 10.6151
R1122 B.n408 B.n407 10.6151
R1123 B.n407 B.n404 10.6151
R1124 B.n404 B.n403 10.6151
R1125 B.n403 B.n400 10.6151
R1126 B.n400 B.n399 10.6151
R1127 B.n399 B.n396 10.6151
R1128 B.n396 B.n339 10.6151
R1129 B.n599 B.n339 10.6151
R1130 B.n601 B.n600 10.6151
R1131 B.n601 B.n330 10.6151
R1132 B.n611 B.n330 10.6151
R1133 B.n612 B.n611 10.6151
R1134 B.n613 B.n612 10.6151
R1135 B.n613 B.n323 10.6151
R1136 B.n623 B.n323 10.6151
R1137 B.n624 B.n623 10.6151
R1138 B.n625 B.n624 10.6151
R1139 B.n625 B.n315 10.6151
R1140 B.n635 B.n315 10.6151
R1141 B.n636 B.n635 10.6151
R1142 B.n637 B.n636 10.6151
R1143 B.n637 B.n308 10.6151
R1144 B.n648 B.n308 10.6151
R1145 B.n649 B.n648 10.6151
R1146 B.n651 B.n649 10.6151
R1147 B.n651 B.n650 10.6151
R1148 B.n650 B.n301 10.6151
R1149 B.n663 B.n301 10.6151
R1150 B.n664 B.n663 10.6151
R1151 B.n665 B.n664 10.6151
R1152 B.n666 B.n665 10.6151
R1153 B.n667 B.n666 10.6151
R1154 B.n670 B.n667 10.6151
R1155 B.n671 B.n670 10.6151
R1156 B.n672 B.n671 10.6151
R1157 B.n673 B.n672 10.6151
R1158 B.n675 B.n673 10.6151
R1159 B.n676 B.n675 10.6151
R1160 B.n677 B.n676 10.6151
R1161 B.n678 B.n677 10.6151
R1162 B.n680 B.n678 10.6151
R1163 B.n681 B.n680 10.6151
R1164 B.n682 B.n681 10.6151
R1165 B.n683 B.n682 10.6151
R1166 B.n685 B.n683 10.6151
R1167 B.n686 B.n685 10.6151
R1168 B.n687 B.n686 10.6151
R1169 B.n688 B.n687 10.6151
R1170 B.n690 B.n688 10.6151
R1171 B.n691 B.n690 10.6151
R1172 B.n692 B.n691 10.6151
R1173 B.n734 B.n1 10.6151
R1174 B.n734 B.n733 10.6151
R1175 B.n733 B.n732 10.6151
R1176 B.n732 B.n10 10.6151
R1177 B.n726 B.n10 10.6151
R1178 B.n726 B.n725 10.6151
R1179 B.n725 B.n724 10.6151
R1180 B.n724 B.n17 10.6151
R1181 B.n718 B.n17 10.6151
R1182 B.n718 B.n717 10.6151
R1183 B.n717 B.n716 10.6151
R1184 B.n716 B.n25 10.6151
R1185 B.n710 B.n25 10.6151
R1186 B.n710 B.n709 10.6151
R1187 B.n709 B.n708 10.6151
R1188 B.n708 B.n32 10.6151
R1189 B.n702 B.n32 10.6151
R1190 B.n702 B.n701 10.6151
R1191 B.n701 B.n700 10.6151
R1192 B.n700 B.n39 10.6151
R1193 B.n102 B.n101 10.6151
R1194 B.n105 B.n102 10.6151
R1195 B.n106 B.n105 10.6151
R1196 B.n109 B.n106 10.6151
R1197 B.n110 B.n109 10.6151
R1198 B.n113 B.n110 10.6151
R1199 B.n114 B.n113 10.6151
R1200 B.n117 B.n114 10.6151
R1201 B.n118 B.n117 10.6151
R1202 B.n121 B.n118 10.6151
R1203 B.n122 B.n121 10.6151
R1204 B.n125 B.n122 10.6151
R1205 B.n126 B.n125 10.6151
R1206 B.n129 B.n126 10.6151
R1207 B.n130 B.n129 10.6151
R1208 B.n133 B.n130 10.6151
R1209 B.n134 B.n133 10.6151
R1210 B.n137 B.n134 10.6151
R1211 B.n138 B.n137 10.6151
R1212 B.n141 B.n138 10.6151
R1213 B.n142 B.n141 10.6151
R1214 B.n145 B.n142 10.6151
R1215 B.n146 B.n145 10.6151
R1216 B.n149 B.n146 10.6151
R1217 B.n150 B.n149 10.6151
R1218 B.n153 B.n150 10.6151
R1219 B.n154 B.n153 10.6151
R1220 B.n157 B.n154 10.6151
R1221 B.n158 B.n157 10.6151
R1222 B.n161 B.n158 10.6151
R1223 B.n162 B.n161 10.6151
R1224 B.n165 B.n162 10.6151
R1225 B.n166 B.n165 10.6151
R1226 B.n169 B.n166 10.6151
R1227 B.n170 B.n169 10.6151
R1228 B.n173 B.n170 10.6151
R1229 B.n174 B.n173 10.6151
R1230 B.n177 B.n174 10.6151
R1231 B.n178 B.n177 10.6151
R1232 B.n181 B.n178 10.6151
R1233 B.n182 B.n181 10.6151
R1234 B.n185 B.n182 10.6151
R1235 B.n186 B.n185 10.6151
R1236 B.n189 B.n186 10.6151
R1237 B.n190 B.n189 10.6151
R1238 B.n194 B.n193 10.6151
R1239 B.n197 B.n194 10.6151
R1240 B.n198 B.n197 10.6151
R1241 B.n201 B.n198 10.6151
R1242 B.n202 B.n201 10.6151
R1243 B.n205 B.n202 10.6151
R1244 B.n206 B.n205 10.6151
R1245 B.n209 B.n206 10.6151
R1246 B.n210 B.n209 10.6151
R1247 B.n214 B.n213 10.6151
R1248 B.n217 B.n214 10.6151
R1249 B.n218 B.n217 10.6151
R1250 B.n221 B.n218 10.6151
R1251 B.n222 B.n221 10.6151
R1252 B.n225 B.n222 10.6151
R1253 B.n226 B.n225 10.6151
R1254 B.n229 B.n226 10.6151
R1255 B.n230 B.n229 10.6151
R1256 B.n233 B.n230 10.6151
R1257 B.n234 B.n233 10.6151
R1258 B.n237 B.n234 10.6151
R1259 B.n238 B.n237 10.6151
R1260 B.n241 B.n238 10.6151
R1261 B.n242 B.n241 10.6151
R1262 B.n245 B.n242 10.6151
R1263 B.n246 B.n245 10.6151
R1264 B.n249 B.n246 10.6151
R1265 B.n250 B.n249 10.6151
R1266 B.n253 B.n250 10.6151
R1267 B.n254 B.n253 10.6151
R1268 B.n257 B.n254 10.6151
R1269 B.n258 B.n257 10.6151
R1270 B.n261 B.n258 10.6151
R1271 B.n262 B.n261 10.6151
R1272 B.n265 B.n262 10.6151
R1273 B.n266 B.n265 10.6151
R1274 B.n269 B.n266 10.6151
R1275 B.n270 B.n269 10.6151
R1276 B.n273 B.n270 10.6151
R1277 B.n274 B.n273 10.6151
R1278 B.n277 B.n274 10.6151
R1279 B.n278 B.n277 10.6151
R1280 B.n281 B.n278 10.6151
R1281 B.n282 B.n281 10.6151
R1282 B.n285 B.n282 10.6151
R1283 B.n286 B.n285 10.6151
R1284 B.n289 B.n286 10.6151
R1285 B.n290 B.n289 10.6151
R1286 B.n293 B.n290 10.6151
R1287 B.n294 B.n293 10.6151
R1288 B.n297 B.n294 10.6151
R1289 B.n299 B.n297 10.6151
R1290 B.n300 B.n299 10.6151
R1291 B.n693 B.n300 10.6151
R1292 B.n506 B.n505 9.36635
R1293 B.n484 B.n483 9.36635
R1294 B.n190 B.n99 9.36635
R1295 B.n213 B.n96 9.36635
R1296 B.n653 B.t5 8.72835
R1297 B.n12 B.t0 8.72835
R1298 B.n742 B.n0 8.11757
R1299 B.n742 B.n1 8.11757
R1300 B.n646 B.t2 5.23721
R1301 B.n728 B.t4 5.23721
R1302 B.n615 B.t11 1.74607
R1303 B.n706 B.t7 1.74607
R1304 B.n505 B.n504 1.24928
R1305 B.n485 B.n484 1.24928
R1306 B.n193 B.n99 1.24928
R1307 B.n210 B.n96 1.24928
R1308 VN.n1 VN.t5 477.998
R1309 VN.n7 VN.t2 477.998
R1310 VN.n2 VN.t3 454.33
R1311 VN.n4 VN.t1 454.33
R1312 VN.n8 VN.t4 454.33
R1313 VN.n10 VN.t0 454.33
R1314 VN.n5 VN.n4 161.3
R1315 VN.n11 VN.n10 161.3
R1316 VN.n9 VN.n6 161.3
R1317 VN.n3 VN.n0 161.3
R1318 VN.n7 VN.n6 44.9044
R1319 VN.n1 VN.n0 44.9044
R1320 VN VN.n11 43.3585
R1321 VN.n4 VN.n3 34.3247
R1322 VN.n10 VN.n9 34.3247
R1323 VN.n2 VN.n1 17.9645
R1324 VN.n8 VN.n7 17.9645
R1325 VN.n3 VN.n2 13.8763
R1326 VN.n9 VN.n8 13.8763
R1327 VN.n11 VN.n6 0.189894
R1328 VN.n5 VN.n0 0.189894
R1329 VN VN.n5 0.0516364
R1330 VDD2.n1 VDD2.t0 64.5589
R1331 VDD2.n2 VDD2.t5 63.8774
R1332 VDD2.n1 VDD2.n0 62.6148
R1333 VDD2 VDD2.n3 62.612
R1334 VDD2.n2 VDD2.n1 38.6593
R1335 VDD2.n3 VDD2.t1 1.45318
R1336 VDD2.n3 VDD2.t3 1.45318
R1337 VDD2.n0 VDD2.t2 1.45318
R1338 VDD2.n0 VDD2.t4 1.45318
R1339 VDD2 VDD2.n2 0.795759
C0 VDD1 VN 0.148173f
C1 VTAIL VP 4.90225f
C2 VDD1 VTAIL 10.4415f
C3 VTAIL VN 4.887609f
C4 VDD2 VP 0.307021f
C5 VDD1 VDD2 0.750287f
C6 VDD2 VN 5.23501f
C7 VDD2 VTAIL 10.475901f
C8 VDD1 VP 5.38894f
C9 VN VP 5.48535f
C10 VDD2 B 4.864525f
C11 VDD1 B 5.102574f
C12 VTAIL B 7.09354f
C13 VN B 8.18454f
C14 VP B 6.201552f
C15 VDD2.t0 B 2.834f
C16 VDD2.t2 B 0.246454f
C17 VDD2.t4 B 0.246454f
C18 VDD2.n0 B 2.21963f
C19 VDD2.n1 B 2.03459f
C20 VDD2.t5 B 2.83078f
C21 VDD2.n2 B 2.22395f
C22 VDD2.t1 B 0.246454f
C23 VDD2.t3 B 0.246454f
C24 VDD2.n3 B 2.21961f
C25 VN.n0 B 0.188433f
C26 VN.t5 B 1.39013f
C27 VN.n1 B 0.509673f
C28 VN.t3 B 1.36378f
C29 VN.n2 B 0.534416f
C30 VN.n3 B 0.009848f
C31 VN.t1 B 1.36378f
C32 VN.n4 B 0.530423f
C33 VN.n5 B 0.033632f
C34 VN.n6 B 0.188433f
C35 VN.t2 B 1.39013f
C36 VN.n7 B 0.509673f
C37 VN.t4 B 1.36378f
C38 VN.n8 B 0.534416f
C39 VN.n9 B 0.009848f
C40 VN.t0 B 1.36378f
C41 VN.n10 B 0.530423f
C42 VN.n11 B 1.88931f
C43 VDD1.t3 B 2.83741f
C44 VDD1.t5 B 2.83678f
C45 VDD1.t4 B 0.246696f
C46 VDD1.t2 B 0.246696f
C47 VDD1.n0 B 2.22181f
C48 VDD1.n1 B 2.1101f
C49 VDD1.t1 B 0.246696f
C50 VDD1.t0 B 0.246696f
C51 VDD1.n2 B 2.22095f
C52 VDD1.n3 B 2.2047f
C53 VTAIL.t0 B 0.255233f
C54 VTAIL.t4 B 0.255233f
C55 VTAIL.n0 B 2.22979f
C56 VTAIL.n1 B 0.323474f
C57 VTAIL.t9 B 2.84368f
C58 VTAIL.n2 B 0.457509f
C59 VTAIL.t8 B 0.255233f
C60 VTAIL.t6 B 0.255233f
C61 VTAIL.n3 B 2.22979f
C62 VTAIL.n4 B 1.67107f
C63 VTAIL.t1 B 0.255233f
C64 VTAIL.t2 B 0.255233f
C65 VTAIL.n5 B 2.22979f
C66 VTAIL.n6 B 1.67107f
C67 VTAIL.t5 B 2.84369f
C68 VTAIL.n7 B 0.457506f
C69 VTAIL.t7 B 0.255233f
C70 VTAIL.t11 B 0.255233f
C71 VTAIL.n8 B 2.22979f
C72 VTAIL.n9 B 0.375308f
C73 VTAIL.t10 B 2.84368f
C74 VTAIL.n10 B 1.67823f
C75 VTAIL.t3 B 2.84368f
C76 VTAIL.n11 B 1.65503f
C77 VP.n0 B 0.044128f
C78 VP.n1 B 0.010014f
C79 VP.n2 B 0.191598f
C80 VP.t5 B 1.38669f
C81 VP.t4 B 1.38669f
C82 VP.t2 B 1.41348f
C83 VP.n3 B 0.518234f
C84 VP.n4 B 0.543392f
C85 VP.n5 B 0.010014f
C86 VP.n6 B 0.539332f
C87 VP.n7 B 1.89212f
C88 VP.t0 B 1.38669f
C89 VP.n8 B 0.539332f
C90 VP.n9 B 1.92903f
C91 VP.n10 B 0.044128f
C92 VP.n11 B 0.044128f
C93 VP.t1 B 1.38669f
C94 VP.n12 B 0.538108f
C95 VP.n13 B 0.010014f
C96 VP.t3 B 1.38669f
C97 VP.n14 B 0.539332f
C98 VP.n15 B 0.034197f
.ends

