* NGSPICE file created from diff_pair_sample_0036.ext - technology: sky130A

.subckt diff_pair_sample_0036 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0 ps=0 w=4.35 l=1.4
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0 ps=0 w=4.35 l=1.4
X2 VTAIL.t7 VP.t0 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0.71775 ps=4.68 w=4.35 l=1.4
X3 VDD1.t2 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.71775 pd=4.68 as=1.6965 ps=9.48 w=4.35 l=1.4
X4 VTAIL.t5 VP.t2 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0.71775 ps=4.68 w=4.35 l=1.4
X5 VDD1.t1 VP.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.71775 pd=4.68 as=1.6965 ps=9.48 w=4.35 l=1.4
X6 VDD2.t3 VN.t0 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.71775 pd=4.68 as=1.6965 ps=9.48 w=4.35 l=1.4
X7 VTAIL.t0 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0.71775 ps=4.68 w=4.35 l=1.4
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0 ps=0 w=4.35 l=1.4
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0 ps=0 w=4.35 l=1.4
X10 VDD2.t1 VN.t2 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.71775 pd=4.68 as=1.6965 ps=9.48 w=4.35 l=1.4
X11 VTAIL.t3 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6965 pd=9.48 as=0.71775 ps=4.68 w=4.35 l=1.4
R0 B.n437 B.n436 585
R1 B.n165 B.n69 585
R2 B.n164 B.n163 585
R3 B.n162 B.n161 585
R4 B.n160 B.n159 585
R5 B.n158 B.n157 585
R6 B.n156 B.n155 585
R7 B.n154 B.n153 585
R8 B.n152 B.n151 585
R9 B.n150 B.n149 585
R10 B.n148 B.n147 585
R11 B.n146 B.n145 585
R12 B.n144 B.n143 585
R13 B.n142 B.n141 585
R14 B.n140 B.n139 585
R15 B.n138 B.n137 585
R16 B.n136 B.n135 585
R17 B.n134 B.n133 585
R18 B.n132 B.n131 585
R19 B.n129 B.n128 585
R20 B.n127 B.n126 585
R21 B.n125 B.n124 585
R22 B.n123 B.n122 585
R23 B.n121 B.n120 585
R24 B.n119 B.n118 585
R25 B.n117 B.n116 585
R26 B.n115 B.n114 585
R27 B.n113 B.n112 585
R28 B.n111 B.n110 585
R29 B.n108 B.n107 585
R30 B.n106 B.n105 585
R31 B.n104 B.n103 585
R32 B.n102 B.n101 585
R33 B.n100 B.n99 585
R34 B.n98 B.n97 585
R35 B.n96 B.n95 585
R36 B.n94 B.n93 585
R37 B.n92 B.n91 585
R38 B.n90 B.n89 585
R39 B.n88 B.n87 585
R40 B.n86 B.n85 585
R41 B.n84 B.n83 585
R42 B.n82 B.n81 585
R43 B.n80 B.n79 585
R44 B.n78 B.n77 585
R45 B.n76 B.n75 585
R46 B.n46 B.n45 585
R47 B.n442 B.n441 585
R48 B.n435 B.n70 585
R49 B.n70 B.n43 585
R50 B.n434 B.n42 585
R51 B.n446 B.n42 585
R52 B.n433 B.n41 585
R53 B.n447 B.n41 585
R54 B.n432 B.n40 585
R55 B.n448 B.n40 585
R56 B.n431 B.n430 585
R57 B.n430 B.n36 585
R58 B.n429 B.n35 585
R59 B.n454 B.n35 585
R60 B.n428 B.n34 585
R61 B.n455 B.n34 585
R62 B.n427 B.n33 585
R63 B.n456 B.n33 585
R64 B.n426 B.n425 585
R65 B.n425 B.n29 585
R66 B.n424 B.n28 585
R67 B.n462 B.n28 585
R68 B.n423 B.n27 585
R69 B.n463 B.n27 585
R70 B.n422 B.n26 585
R71 B.n464 B.n26 585
R72 B.n421 B.n420 585
R73 B.n420 B.n22 585
R74 B.n419 B.n21 585
R75 B.n470 B.n21 585
R76 B.n418 B.n20 585
R77 B.n471 B.n20 585
R78 B.n417 B.n19 585
R79 B.n472 B.n19 585
R80 B.n416 B.n415 585
R81 B.n415 B.n15 585
R82 B.n414 B.n14 585
R83 B.n478 B.n14 585
R84 B.n413 B.n13 585
R85 B.n479 B.n13 585
R86 B.n412 B.n12 585
R87 B.n480 B.n12 585
R88 B.n411 B.n410 585
R89 B.n410 B.n409 585
R90 B.n408 B.n407 585
R91 B.n408 B.n8 585
R92 B.n406 B.n7 585
R93 B.n487 B.n7 585
R94 B.n405 B.n6 585
R95 B.n488 B.n6 585
R96 B.n404 B.n5 585
R97 B.n489 B.n5 585
R98 B.n403 B.n402 585
R99 B.n402 B.n4 585
R100 B.n401 B.n166 585
R101 B.n401 B.n400 585
R102 B.n391 B.n167 585
R103 B.n168 B.n167 585
R104 B.n393 B.n392 585
R105 B.n394 B.n393 585
R106 B.n390 B.n173 585
R107 B.n173 B.n172 585
R108 B.n389 B.n388 585
R109 B.n388 B.n387 585
R110 B.n175 B.n174 585
R111 B.n176 B.n175 585
R112 B.n380 B.n379 585
R113 B.n381 B.n380 585
R114 B.n378 B.n180 585
R115 B.n184 B.n180 585
R116 B.n377 B.n376 585
R117 B.n376 B.n375 585
R118 B.n182 B.n181 585
R119 B.n183 B.n182 585
R120 B.n368 B.n367 585
R121 B.n369 B.n368 585
R122 B.n366 B.n189 585
R123 B.n189 B.n188 585
R124 B.n365 B.n364 585
R125 B.n364 B.n363 585
R126 B.n191 B.n190 585
R127 B.n192 B.n191 585
R128 B.n356 B.n355 585
R129 B.n357 B.n356 585
R130 B.n354 B.n197 585
R131 B.n197 B.n196 585
R132 B.n353 B.n352 585
R133 B.n352 B.n351 585
R134 B.n199 B.n198 585
R135 B.n200 B.n199 585
R136 B.n344 B.n343 585
R137 B.n345 B.n344 585
R138 B.n342 B.n205 585
R139 B.n205 B.n204 585
R140 B.n341 B.n340 585
R141 B.n340 B.n339 585
R142 B.n207 B.n206 585
R143 B.n208 B.n207 585
R144 B.n335 B.n334 585
R145 B.n211 B.n210 585
R146 B.n331 B.n330 585
R147 B.n332 B.n331 585
R148 B.n329 B.n235 585
R149 B.n328 B.n327 585
R150 B.n326 B.n325 585
R151 B.n324 B.n323 585
R152 B.n322 B.n321 585
R153 B.n320 B.n319 585
R154 B.n318 B.n317 585
R155 B.n316 B.n315 585
R156 B.n314 B.n313 585
R157 B.n312 B.n311 585
R158 B.n310 B.n309 585
R159 B.n308 B.n307 585
R160 B.n306 B.n305 585
R161 B.n304 B.n303 585
R162 B.n302 B.n301 585
R163 B.n300 B.n299 585
R164 B.n298 B.n297 585
R165 B.n296 B.n295 585
R166 B.n294 B.n293 585
R167 B.n292 B.n291 585
R168 B.n290 B.n289 585
R169 B.n288 B.n287 585
R170 B.n286 B.n285 585
R171 B.n284 B.n283 585
R172 B.n282 B.n281 585
R173 B.n280 B.n279 585
R174 B.n278 B.n277 585
R175 B.n276 B.n275 585
R176 B.n274 B.n273 585
R177 B.n272 B.n271 585
R178 B.n270 B.n269 585
R179 B.n268 B.n267 585
R180 B.n266 B.n265 585
R181 B.n264 B.n263 585
R182 B.n262 B.n261 585
R183 B.n260 B.n259 585
R184 B.n258 B.n257 585
R185 B.n256 B.n255 585
R186 B.n254 B.n253 585
R187 B.n252 B.n251 585
R188 B.n250 B.n249 585
R189 B.n248 B.n247 585
R190 B.n246 B.n245 585
R191 B.n244 B.n243 585
R192 B.n242 B.n234 585
R193 B.n332 B.n234 585
R194 B.n336 B.n209 585
R195 B.n209 B.n208 585
R196 B.n338 B.n337 585
R197 B.n339 B.n338 585
R198 B.n203 B.n202 585
R199 B.n204 B.n203 585
R200 B.n347 B.n346 585
R201 B.n346 B.n345 585
R202 B.n348 B.n201 585
R203 B.n201 B.n200 585
R204 B.n350 B.n349 585
R205 B.n351 B.n350 585
R206 B.n195 B.n194 585
R207 B.n196 B.n195 585
R208 B.n359 B.n358 585
R209 B.n358 B.n357 585
R210 B.n360 B.n193 585
R211 B.n193 B.n192 585
R212 B.n362 B.n361 585
R213 B.n363 B.n362 585
R214 B.n187 B.n186 585
R215 B.n188 B.n187 585
R216 B.n371 B.n370 585
R217 B.n370 B.n369 585
R218 B.n372 B.n185 585
R219 B.n185 B.n183 585
R220 B.n374 B.n373 585
R221 B.n375 B.n374 585
R222 B.n179 B.n178 585
R223 B.n184 B.n179 585
R224 B.n383 B.n382 585
R225 B.n382 B.n381 585
R226 B.n384 B.n177 585
R227 B.n177 B.n176 585
R228 B.n386 B.n385 585
R229 B.n387 B.n386 585
R230 B.n171 B.n170 585
R231 B.n172 B.n171 585
R232 B.n396 B.n395 585
R233 B.n395 B.n394 585
R234 B.n397 B.n169 585
R235 B.n169 B.n168 585
R236 B.n399 B.n398 585
R237 B.n400 B.n399 585
R238 B.n3 B.n0 585
R239 B.n4 B.n3 585
R240 B.n486 B.n1 585
R241 B.n487 B.n486 585
R242 B.n485 B.n484 585
R243 B.n485 B.n8 585
R244 B.n483 B.n9 585
R245 B.n409 B.n9 585
R246 B.n482 B.n481 585
R247 B.n481 B.n480 585
R248 B.n11 B.n10 585
R249 B.n479 B.n11 585
R250 B.n477 B.n476 585
R251 B.n478 B.n477 585
R252 B.n475 B.n16 585
R253 B.n16 B.n15 585
R254 B.n474 B.n473 585
R255 B.n473 B.n472 585
R256 B.n18 B.n17 585
R257 B.n471 B.n18 585
R258 B.n469 B.n468 585
R259 B.n470 B.n469 585
R260 B.n467 B.n23 585
R261 B.n23 B.n22 585
R262 B.n466 B.n465 585
R263 B.n465 B.n464 585
R264 B.n25 B.n24 585
R265 B.n463 B.n25 585
R266 B.n461 B.n460 585
R267 B.n462 B.n461 585
R268 B.n459 B.n30 585
R269 B.n30 B.n29 585
R270 B.n458 B.n457 585
R271 B.n457 B.n456 585
R272 B.n32 B.n31 585
R273 B.n455 B.n32 585
R274 B.n453 B.n452 585
R275 B.n454 B.n453 585
R276 B.n451 B.n37 585
R277 B.n37 B.n36 585
R278 B.n450 B.n449 585
R279 B.n449 B.n448 585
R280 B.n39 B.n38 585
R281 B.n447 B.n39 585
R282 B.n445 B.n444 585
R283 B.n446 B.n445 585
R284 B.n443 B.n44 585
R285 B.n44 B.n43 585
R286 B.n490 B.n489 585
R287 B.n488 B.n2 585
R288 B.n441 B.n44 463.671
R289 B.n437 B.n70 463.671
R290 B.n234 B.n207 463.671
R291 B.n334 B.n209 463.671
R292 B.n73 B.t15 279.93
R293 B.n71 B.t4 279.93
R294 B.n239 B.t12 279.93
R295 B.n236 B.t8 279.93
R296 B.n439 B.n438 256.663
R297 B.n439 B.n68 256.663
R298 B.n439 B.n67 256.663
R299 B.n439 B.n66 256.663
R300 B.n439 B.n65 256.663
R301 B.n439 B.n64 256.663
R302 B.n439 B.n63 256.663
R303 B.n439 B.n62 256.663
R304 B.n439 B.n61 256.663
R305 B.n439 B.n60 256.663
R306 B.n439 B.n59 256.663
R307 B.n439 B.n58 256.663
R308 B.n439 B.n57 256.663
R309 B.n439 B.n56 256.663
R310 B.n439 B.n55 256.663
R311 B.n439 B.n54 256.663
R312 B.n439 B.n53 256.663
R313 B.n439 B.n52 256.663
R314 B.n439 B.n51 256.663
R315 B.n439 B.n50 256.663
R316 B.n439 B.n49 256.663
R317 B.n439 B.n48 256.663
R318 B.n439 B.n47 256.663
R319 B.n440 B.n439 256.663
R320 B.n333 B.n332 256.663
R321 B.n332 B.n212 256.663
R322 B.n332 B.n213 256.663
R323 B.n332 B.n214 256.663
R324 B.n332 B.n215 256.663
R325 B.n332 B.n216 256.663
R326 B.n332 B.n217 256.663
R327 B.n332 B.n218 256.663
R328 B.n332 B.n219 256.663
R329 B.n332 B.n220 256.663
R330 B.n332 B.n221 256.663
R331 B.n332 B.n222 256.663
R332 B.n332 B.n223 256.663
R333 B.n332 B.n224 256.663
R334 B.n332 B.n225 256.663
R335 B.n332 B.n226 256.663
R336 B.n332 B.n227 256.663
R337 B.n332 B.n228 256.663
R338 B.n332 B.n229 256.663
R339 B.n332 B.n230 256.663
R340 B.n332 B.n231 256.663
R341 B.n332 B.n232 256.663
R342 B.n332 B.n233 256.663
R343 B.n492 B.n491 256.663
R344 B.n75 B.n46 163.367
R345 B.n79 B.n78 163.367
R346 B.n83 B.n82 163.367
R347 B.n87 B.n86 163.367
R348 B.n91 B.n90 163.367
R349 B.n95 B.n94 163.367
R350 B.n99 B.n98 163.367
R351 B.n103 B.n102 163.367
R352 B.n107 B.n106 163.367
R353 B.n112 B.n111 163.367
R354 B.n116 B.n115 163.367
R355 B.n120 B.n119 163.367
R356 B.n124 B.n123 163.367
R357 B.n128 B.n127 163.367
R358 B.n133 B.n132 163.367
R359 B.n137 B.n136 163.367
R360 B.n141 B.n140 163.367
R361 B.n145 B.n144 163.367
R362 B.n149 B.n148 163.367
R363 B.n153 B.n152 163.367
R364 B.n157 B.n156 163.367
R365 B.n161 B.n160 163.367
R366 B.n163 B.n69 163.367
R367 B.n340 B.n207 163.367
R368 B.n340 B.n205 163.367
R369 B.n344 B.n205 163.367
R370 B.n344 B.n199 163.367
R371 B.n352 B.n199 163.367
R372 B.n352 B.n197 163.367
R373 B.n356 B.n197 163.367
R374 B.n356 B.n191 163.367
R375 B.n364 B.n191 163.367
R376 B.n364 B.n189 163.367
R377 B.n368 B.n189 163.367
R378 B.n368 B.n182 163.367
R379 B.n376 B.n182 163.367
R380 B.n376 B.n180 163.367
R381 B.n380 B.n180 163.367
R382 B.n380 B.n175 163.367
R383 B.n388 B.n175 163.367
R384 B.n388 B.n173 163.367
R385 B.n393 B.n173 163.367
R386 B.n393 B.n167 163.367
R387 B.n401 B.n167 163.367
R388 B.n402 B.n401 163.367
R389 B.n402 B.n5 163.367
R390 B.n6 B.n5 163.367
R391 B.n7 B.n6 163.367
R392 B.n408 B.n7 163.367
R393 B.n410 B.n408 163.367
R394 B.n410 B.n12 163.367
R395 B.n13 B.n12 163.367
R396 B.n14 B.n13 163.367
R397 B.n415 B.n14 163.367
R398 B.n415 B.n19 163.367
R399 B.n20 B.n19 163.367
R400 B.n21 B.n20 163.367
R401 B.n420 B.n21 163.367
R402 B.n420 B.n26 163.367
R403 B.n27 B.n26 163.367
R404 B.n28 B.n27 163.367
R405 B.n425 B.n28 163.367
R406 B.n425 B.n33 163.367
R407 B.n34 B.n33 163.367
R408 B.n35 B.n34 163.367
R409 B.n430 B.n35 163.367
R410 B.n430 B.n40 163.367
R411 B.n41 B.n40 163.367
R412 B.n42 B.n41 163.367
R413 B.n70 B.n42 163.367
R414 B.n331 B.n211 163.367
R415 B.n331 B.n235 163.367
R416 B.n327 B.n326 163.367
R417 B.n323 B.n322 163.367
R418 B.n319 B.n318 163.367
R419 B.n315 B.n314 163.367
R420 B.n311 B.n310 163.367
R421 B.n307 B.n306 163.367
R422 B.n303 B.n302 163.367
R423 B.n299 B.n298 163.367
R424 B.n295 B.n294 163.367
R425 B.n291 B.n290 163.367
R426 B.n287 B.n286 163.367
R427 B.n283 B.n282 163.367
R428 B.n279 B.n278 163.367
R429 B.n275 B.n274 163.367
R430 B.n271 B.n270 163.367
R431 B.n267 B.n266 163.367
R432 B.n263 B.n262 163.367
R433 B.n259 B.n258 163.367
R434 B.n255 B.n254 163.367
R435 B.n251 B.n250 163.367
R436 B.n247 B.n246 163.367
R437 B.n243 B.n234 163.367
R438 B.n338 B.n209 163.367
R439 B.n338 B.n203 163.367
R440 B.n346 B.n203 163.367
R441 B.n346 B.n201 163.367
R442 B.n350 B.n201 163.367
R443 B.n350 B.n195 163.367
R444 B.n358 B.n195 163.367
R445 B.n358 B.n193 163.367
R446 B.n362 B.n193 163.367
R447 B.n362 B.n187 163.367
R448 B.n370 B.n187 163.367
R449 B.n370 B.n185 163.367
R450 B.n374 B.n185 163.367
R451 B.n374 B.n179 163.367
R452 B.n382 B.n179 163.367
R453 B.n382 B.n177 163.367
R454 B.n386 B.n177 163.367
R455 B.n386 B.n171 163.367
R456 B.n395 B.n171 163.367
R457 B.n395 B.n169 163.367
R458 B.n399 B.n169 163.367
R459 B.n399 B.n3 163.367
R460 B.n490 B.n3 163.367
R461 B.n486 B.n2 163.367
R462 B.n486 B.n485 163.367
R463 B.n485 B.n9 163.367
R464 B.n481 B.n9 163.367
R465 B.n481 B.n11 163.367
R466 B.n477 B.n11 163.367
R467 B.n477 B.n16 163.367
R468 B.n473 B.n16 163.367
R469 B.n473 B.n18 163.367
R470 B.n469 B.n18 163.367
R471 B.n469 B.n23 163.367
R472 B.n465 B.n23 163.367
R473 B.n465 B.n25 163.367
R474 B.n461 B.n25 163.367
R475 B.n461 B.n30 163.367
R476 B.n457 B.n30 163.367
R477 B.n457 B.n32 163.367
R478 B.n453 B.n32 163.367
R479 B.n453 B.n37 163.367
R480 B.n449 B.n37 163.367
R481 B.n449 B.n39 163.367
R482 B.n445 B.n39 163.367
R483 B.n445 B.n44 163.367
R484 B.n332 B.n208 131.429
R485 B.n439 B.n43 131.429
R486 B.n71 B.t6 109.754
R487 B.n239 B.t14 109.754
R488 B.n73 B.t16 109.751
R489 B.n236 B.t11 109.751
R490 B.n339 B.n208 77.7148
R491 B.n339 B.n204 77.7148
R492 B.n345 B.n204 77.7148
R493 B.n345 B.n200 77.7148
R494 B.n351 B.n200 77.7148
R495 B.n357 B.n196 77.7148
R496 B.n357 B.n192 77.7148
R497 B.n363 B.n192 77.7148
R498 B.n363 B.n188 77.7148
R499 B.n369 B.n188 77.7148
R500 B.n369 B.n183 77.7148
R501 B.n375 B.n183 77.7148
R502 B.n375 B.n184 77.7148
R503 B.n381 B.n176 77.7148
R504 B.n387 B.n176 77.7148
R505 B.n387 B.n172 77.7148
R506 B.n394 B.n172 77.7148
R507 B.n400 B.n168 77.7148
R508 B.n400 B.n4 77.7148
R509 B.n489 B.n4 77.7148
R510 B.n489 B.n488 77.7148
R511 B.n488 B.n487 77.7148
R512 B.n487 B.n8 77.7148
R513 B.n409 B.n8 77.7148
R514 B.n480 B.n479 77.7148
R515 B.n479 B.n478 77.7148
R516 B.n478 B.n15 77.7148
R517 B.n472 B.n15 77.7148
R518 B.n471 B.n470 77.7148
R519 B.n470 B.n22 77.7148
R520 B.n464 B.n22 77.7148
R521 B.n464 B.n463 77.7148
R522 B.n463 B.n462 77.7148
R523 B.n462 B.n29 77.7148
R524 B.n456 B.n29 77.7148
R525 B.n456 B.n455 77.7148
R526 B.n454 B.n36 77.7148
R527 B.n448 B.n36 77.7148
R528 B.n448 B.n447 77.7148
R529 B.n447 B.n446 77.7148
R530 B.n446 B.n43 77.7148
R531 B.n72 B.t7 76.2026
R532 B.n240 B.t13 76.2026
R533 B.n74 B.t17 76.1987
R534 B.n237 B.t10 76.1987
R535 B.n351 B.t9 75.4291
R536 B.t5 B.n454 75.4291
R537 B.n441 B.n440 71.676
R538 B.n75 B.n47 71.676
R539 B.n79 B.n48 71.676
R540 B.n83 B.n49 71.676
R541 B.n87 B.n50 71.676
R542 B.n91 B.n51 71.676
R543 B.n95 B.n52 71.676
R544 B.n99 B.n53 71.676
R545 B.n103 B.n54 71.676
R546 B.n107 B.n55 71.676
R547 B.n112 B.n56 71.676
R548 B.n116 B.n57 71.676
R549 B.n120 B.n58 71.676
R550 B.n124 B.n59 71.676
R551 B.n128 B.n60 71.676
R552 B.n133 B.n61 71.676
R553 B.n137 B.n62 71.676
R554 B.n141 B.n63 71.676
R555 B.n145 B.n64 71.676
R556 B.n149 B.n65 71.676
R557 B.n153 B.n66 71.676
R558 B.n157 B.n67 71.676
R559 B.n161 B.n68 71.676
R560 B.n438 B.n69 71.676
R561 B.n438 B.n437 71.676
R562 B.n163 B.n68 71.676
R563 B.n160 B.n67 71.676
R564 B.n156 B.n66 71.676
R565 B.n152 B.n65 71.676
R566 B.n148 B.n64 71.676
R567 B.n144 B.n63 71.676
R568 B.n140 B.n62 71.676
R569 B.n136 B.n61 71.676
R570 B.n132 B.n60 71.676
R571 B.n127 B.n59 71.676
R572 B.n123 B.n58 71.676
R573 B.n119 B.n57 71.676
R574 B.n115 B.n56 71.676
R575 B.n111 B.n55 71.676
R576 B.n106 B.n54 71.676
R577 B.n102 B.n53 71.676
R578 B.n98 B.n52 71.676
R579 B.n94 B.n51 71.676
R580 B.n90 B.n50 71.676
R581 B.n86 B.n49 71.676
R582 B.n82 B.n48 71.676
R583 B.n78 B.n47 71.676
R584 B.n440 B.n46 71.676
R585 B.n334 B.n333 71.676
R586 B.n235 B.n212 71.676
R587 B.n326 B.n213 71.676
R588 B.n322 B.n214 71.676
R589 B.n318 B.n215 71.676
R590 B.n314 B.n216 71.676
R591 B.n310 B.n217 71.676
R592 B.n306 B.n218 71.676
R593 B.n302 B.n219 71.676
R594 B.n298 B.n220 71.676
R595 B.n294 B.n221 71.676
R596 B.n290 B.n222 71.676
R597 B.n286 B.n223 71.676
R598 B.n282 B.n224 71.676
R599 B.n278 B.n225 71.676
R600 B.n274 B.n226 71.676
R601 B.n270 B.n227 71.676
R602 B.n266 B.n228 71.676
R603 B.n262 B.n229 71.676
R604 B.n258 B.n230 71.676
R605 B.n254 B.n231 71.676
R606 B.n250 B.n232 71.676
R607 B.n246 B.n233 71.676
R608 B.n333 B.n211 71.676
R609 B.n327 B.n212 71.676
R610 B.n323 B.n213 71.676
R611 B.n319 B.n214 71.676
R612 B.n315 B.n215 71.676
R613 B.n311 B.n216 71.676
R614 B.n307 B.n217 71.676
R615 B.n303 B.n218 71.676
R616 B.n299 B.n219 71.676
R617 B.n295 B.n220 71.676
R618 B.n291 B.n221 71.676
R619 B.n287 B.n222 71.676
R620 B.n283 B.n223 71.676
R621 B.n279 B.n224 71.676
R622 B.n275 B.n225 71.676
R623 B.n271 B.n226 71.676
R624 B.n267 B.n227 71.676
R625 B.n263 B.n228 71.676
R626 B.n259 B.n229 71.676
R627 B.n255 B.n230 71.676
R628 B.n251 B.n231 71.676
R629 B.n247 B.n232 71.676
R630 B.n243 B.n233 71.676
R631 B.n491 B.n490 71.676
R632 B.n491 B.n2 71.676
R633 B.n109 B.n74 59.5399
R634 B.n130 B.n72 59.5399
R635 B.n241 B.n240 59.5399
R636 B.n238 B.n237 59.5399
R637 B.n381 B.t2 57.1434
R638 B.n472 B.t1 57.1434
R639 B.t3 B.n168 50.2862
R640 B.n409 B.t0 50.2862
R641 B.n74 B.n73 33.552
R642 B.n72 B.n71 33.552
R643 B.n240 B.n239 33.552
R644 B.n237 B.n236 33.552
R645 B.n336 B.n335 30.1273
R646 B.n242 B.n206 30.1273
R647 B.n436 B.n435 30.1273
R648 B.n443 B.n442 30.1273
R649 B.n394 B.t3 27.4291
R650 B.n480 B.t0 27.4291
R651 B.n184 B.t2 20.5719
R652 B.t1 B.n471 20.5719
R653 B B.n492 18.0485
R654 B.n337 B.n336 10.6151
R655 B.n337 B.n202 10.6151
R656 B.n347 B.n202 10.6151
R657 B.n348 B.n347 10.6151
R658 B.n349 B.n348 10.6151
R659 B.n349 B.n194 10.6151
R660 B.n359 B.n194 10.6151
R661 B.n360 B.n359 10.6151
R662 B.n361 B.n360 10.6151
R663 B.n361 B.n186 10.6151
R664 B.n371 B.n186 10.6151
R665 B.n372 B.n371 10.6151
R666 B.n373 B.n372 10.6151
R667 B.n373 B.n178 10.6151
R668 B.n383 B.n178 10.6151
R669 B.n384 B.n383 10.6151
R670 B.n385 B.n384 10.6151
R671 B.n385 B.n170 10.6151
R672 B.n396 B.n170 10.6151
R673 B.n397 B.n396 10.6151
R674 B.n398 B.n397 10.6151
R675 B.n398 B.n0 10.6151
R676 B.n335 B.n210 10.6151
R677 B.n330 B.n210 10.6151
R678 B.n330 B.n329 10.6151
R679 B.n329 B.n328 10.6151
R680 B.n328 B.n325 10.6151
R681 B.n325 B.n324 10.6151
R682 B.n324 B.n321 10.6151
R683 B.n321 B.n320 10.6151
R684 B.n320 B.n317 10.6151
R685 B.n317 B.n316 10.6151
R686 B.n316 B.n313 10.6151
R687 B.n313 B.n312 10.6151
R688 B.n312 B.n309 10.6151
R689 B.n309 B.n308 10.6151
R690 B.n308 B.n305 10.6151
R691 B.n305 B.n304 10.6151
R692 B.n304 B.n301 10.6151
R693 B.n301 B.n300 10.6151
R694 B.n297 B.n296 10.6151
R695 B.n296 B.n293 10.6151
R696 B.n293 B.n292 10.6151
R697 B.n292 B.n289 10.6151
R698 B.n289 B.n288 10.6151
R699 B.n288 B.n285 10.6151
R700 B.n285 B.n284 10.6151
R701 B.n284 B.n281 10.6151
R702 B.n281 B.n280 10.6151
R703 B.n277 B.n276 10.6151
R704 B.n276 B.n273 10.6151
R705 B.n273 B.n272 10.6151
R706 B.n272 B.n269 10.6151
R707 B.n269 B.n268 10.6151
R708 B.n268 B.n265 10.6151
R709 B.n265 B.n264 10.6151
R710 B.n264 B.n261 10.6151
R711 B.n261 B.n260 10.6151
R712 B.n260 B.n257 10.6151
R713 B.n257 B.n256 10.6151
R714 B.n256 B.n253 10.6151
R715 B.n253 B.n252 10.6151
R716 B.n252 B.n249 10.6151
R717 B.n249 B.n248 10.6151
R718 B.n248 B.n245 10.6151
R719 B.n245 B.n244 10.6151
R720 B.n244 B.n242 10.6151
R721 B.n341 B.n206 10.6151
R722 B.n342 B.n341 10.6151
R723 B.n343 B.n342 10.6151
R724 B.n343 B.n198 10.6151
R725 B.n353 B.n198 10.6151
R726 B.n354 B.n353 10.6151
R727 B.n355 B.n354 10.6151
R728 B.n355 B.n190 10.6151
R729 B.n365 B.n190 10.6151
R730 B.n366 B.n365 10.6151
R731 B.n367 B.n366 10.6151
R732 B.n367 B.n181 10.6151
R733 B.n377 B.n181 10.6151
R734 B.n378 B.n377 10.6151
R735 B.n379 B.n378 10.6151
R736 B.n379 B.n174 10.6151
R737 B.n389 B.n174 10.6151
R738 B.n390 B.n389 10.6151
R739 B.n392 B.n390 10.6151
R740 B.n392 B.n391 10.6151
R741 B.n391 B.n166 10.6151
R742 B.n403 B.n166 10.6151
R743 B.n404 B.n403 10.6151
R744 B.n405 B.n404 10.6151
R745 B.n406 B.n405 10.6151
R746 B.n407 B.n406 10.6151
R747 B.n411 B.n407 10.6151
R748 B.n412 B.n411 10.6151
R749 B.n413 B.n412 10.6151
R750 B.n414 B.n413 10.6151
R751 B.n416 B.n414 10.6151
R752 B.n417 B.n416 10.6151
R753 B.n418 B.n417 10.6151
R754 B.n419 B.n418 10.6151
R755 B.n421 B.n419 10.6151
R756 B.n422 B.n421 10.6151
R757 B.n423 B.n422 10.6151
R758 B.n424 B.n423 10.6151
R759 B.n426 B.n424 10.6151
R760 B.n427 B.n426 10.6151
R761 B.n428 B.n427 10.6151
R762 B.n429 B.n428 10.6151
R763 B.n431 B.n429 10.6151
R764 B.n432 B.n431 10.6151
R765 B.n433 B.n432 10.6151
R766 B.n434 B.n433 10.6151
R767 B.n435 B.n434 10.6151
R768 B.n484 B.n1 10.6151
R769 B.n484 B.n483 10.6151
R770 B.n483 B.n482 10.6151
R771 B.n482 B.n10 10.6151
R772 B.n476 B.n10 10.6151
R773 B.n476 B.n475 10.6151
R774 B.n475 B.n474 10.6151
R775 B.n474 B.n17 10.6151
R776 B.n468 B.n17 10.6151
R777 B.n468 B.n467 10.6151
R778 B.n467 B.n466 10.6151
R779 B.n466 B.n24 10.6151
R780 B.n460 B.n24 10.6151
R781 B.n460 B.n459 10.6151
R782 B.n459 B.n458 10.6151
R783 B.n458 B.n31 10.6151
R784 B.n452 B.n31 10.6151
R785 B.n452 B.n451 10.6151
R786 B.n451 B.n450 10.6151
R787 B.n450 B.n38 10.6151
R788 B.n444 B.n38 10.6151
R789 B.n444 B.n443 10.6151
R790 B.n442 B.n45 10.6151
R791 B.n76 B.n45 10.6151
R792 B.n77 B.n76 10.6151
R793 B.n80 B.n77 10.6151
R794 B.n81 B.n80 10.6151
R795 B.n84 B.n81 10.6151
R796 B.n85 B.n84 10.6151
R797 B.n88 B.n85 10.6151
R798 B.n89 B.n88 10.6151
R799 B.n92 B.n89 10.6151
R800 B.n93 B.n92 10.6151
R801 B.n96 B.n93 10.6151
R802 B.n97 B.n96 10.6151
R803 B.n100 B.n97 10.6151
R804 B.n101 B.n100 10.6151
R805 B.n104 B.n101 10.6151
R806 B.n105 B.n104 10.6151
R807 B.n108 B.n105 10.6151
R808 B.n113 B.n110 10.6151
R809 B.n114 B.n113 10.6151
R810 B.n117 B.n114 10.6151
R811 B.n118 B.n117 10.6151
R812 B.n121 B.n118 10.6151
R813 B.n122 B.n121 10.6151
R814 B.n125 B.n122 10.6151
R815 B.n126 B.n125 10.6151
R816 B.n129 B.n126 10.6151
R817 B.n134 B.n131 10.6151
R818 B.n135 B.n134 10.6151
R819 B.n138 B.n135 10.6151
R820 B.n139 B.n138 10.6151
R821 B.n142 B.n139 10.6151
R822 B.n143 B.n142 10.6151
R823 B.n146 B.n143 10.6151
R824 B.n147 B.n146 10.6151
R825 B.n150 B.n147 10.6151
R826 B.n151 B.n150 10.6151
R827 B.n154 B.n151 10.6151
R828 B.n155 B.n154 10.6151
R829 B.n158 B.n155 10.6151
R830 B.n159 B.n158 10.6151
R831 B.n162 B.n159 10.6151
R832 B.n164 B.n162 10.6151
R833 B.n165 B.n164 10.6151
R834 B.n436 B.n165 10.6151
R835 B.n300 B.n238 9.36635
R836 B.n277 B.n241 9.36635
R837 B.n109 B.n108 9.36635
R838 B.n131 B.n130 9.36635
R839 B.n492 B.n0 8.11757
R840 B.n492 B.n1 8.11757
R841 B.t9 B.n196 2.28621
R842 B.n455 B.t5 2.28621
R843 B.n297 B.n238 1.24928
R844 B.n280 B.n241 1.24928
R845 B.n110 B.n109 1.24928
R846 B.n130 B.n129 1.24928
R847 VP.n4 VP.n3 180.141
R848 VP.n12 VP.n11 180.141
R849 VP.n10 VP.n0 161.3
R850 VP.n9 VP.n8 161.3
R851 VP.n7 VP.n1 161.3
R852 VP.n6 VP.n5 161.3
R853 VP.n2 VP.t0 109.757
R854 VP.n2 VP.t1 109.45
R855 VP.n4 VP.t2 74.8826
R856 VP.n11 VP.t3 74.8826
R857 VP.n9 VP.n1 56.5193
R858 VP.n3 VP.n2 50.0666
R859 VP.n5 VP.n1 24.4675
R860 VP.n10 VP.n9 24.4675
R861 VP.n5 VP.n4 5.62791
R862 VP.n11 VP.n10 5.62791
R863 VP.n6 VP.n3 0.189894
R864 VP.n7 VP.n6 0.189894
R865 VP.n8 VP.n7 0.189894
R866 VP.n8 VP.n0 0.189894
R867 VP.n12 VP.n0 0.189894
R868 VP VP.n12 0.0516364
R869 VDD1 VDD1.n1 107.291
R870 VDD1 VDD1.n0 74.8856
R871 VDD1.n0 VDD1.t0 4.55222
R872 VDD1.n0 VDD1.t2 4.55222
R873 VDD1.n1 VDD1.t3 4.55222
R874 VDD1.n1 VDD1.t1 4.55222
R875 VTAIL.n5 VTAIL.t7 62.7005
R876 VTAIL.n4 VTAIL.t1 62.7005
R877 VTAIL.n3 VTAIL.t0 62.7005
R878 VTAIL.n7 VTAIL.t2 62.7002
R879 VTAIL.n0 VTAIL.t3 62.7002
R880 VTAIL.n1 VTAIL.t4 62.7002
R881 VTAIL.n2 VTAIL.t5 62.7002
R882 VTAIL.n6 VTAIL.t6 62.7002
R883 VTAIL.n7 VTAIL.n6 17.6083
R884 VTAIL.n3 VTAIL.n2 17.6083
R885 VTAIL.n4 VTAIL.n3 1.49188
R886 VTAIL.n6 VTAIL.n5 1.49188
R887 VTAIL.n2 VTAIL.n1 1.49188
R888 VTAIL VTAIL.n0 0.804379
R889 VTAIL VTAIL.n7 0.688
R890 VTAIL.n5 VTAIL.n4 0.470328
R891 VTAIL.n1 VTAIL.n0 0.470328
R892 VN.n0 VN.t3 109.757
R893 VN.n1 VN.t0 109.757
R894 VN.n0 VN.t2 109.45
R895 VN.n1 VN.t1 109.45
R896 VN VN.n1 50.4473
R897 VN VN.n0 13.4208
R898 VDD2.n2 VDD2.n0 106.766
R899 VDD2.n2 VDD2.n1 74.8274
R900 VDD2.n1 VDD2.t2 4.55222
R901 VDD2.n1 VDD2.t3 4.55222
R902 VDD2.n0 VDD2.t0 4.55222
R903 VDD2.n0 VDD2.t1 4.55222
R904 VDD2 VDD2.n2 0.0586897
C0 VDD1 VTAIL 3.21492f
C1 VDD2 VTAIL 3.26108f
C2 VN VTAIL 1.81051f
C3 VDD1 VP 1.84746f
C4 VDD2 VP 0.322491f
C5 VN VP 3.91911f
C6 VDD1 VDD2 0.735181f
C7 VDD1 VN 0.152101f
C8 VN VDD2 1.67789f
C9 VTAIL VP 1.82462f
C10 VDD2 B 2.446563f
C11 VDD1 B 4.36386f
C12 VTAIL B 4.640734f
C13 VN B 6.90646f
C14 VP B 5.731505f
C15 VDD2.t0 B 0.062292f
C16 VDD2.t1 B 0.062292f
C17 VDD2.n0 B 0.716675f
C18 VDD2.t2 B 0.062292f
C19 VDD2.t3 B 0.062292f
C20 VDD2.n1 B 0.49631f
C21 VDD2.n2 B 1.74686f
C22 VN.t3 B 0.401105f
C23 VN.t2 B 0.400462f
C24 VN.n0 B 0.324524f
C25 VN.t0 B 0.401105f
C26 VN.t1 B 0.400462f
C27 VN.n1 B 0.921747f
C28 VTAIL.t3 B 0.409661f
C29 VTAIL.n0 B 0.191118f
C30 VTAIL.t4 B 0.409661f
C31 VTAIL.n1 B 0.219212f
C32 VTAIL.t5 B 0.409661f
C33 VTAIL.n2 B 0.586466f
C34 VTAIL.t0 B 0.409663f
C35 VTAIL.n3 B 0.586464f
C36 VTAIL.t1 B 0.409663f
C37 VTAIL.n4 B 0.219211f
C38 VTAIL.t7 B 0.409663f
C39 VTAIL.n5 B 0.219211f
C40 VTAIL.t6 B 0.409661f
C41 VTAIL.n6 B 0.586466f
C42 VTAIL.t2 B 0.409661f
C43 VTAIL.n7 B 0.553616f
C44 VDD1.t0 B 0.059203f
C45 VDD1.t2 B 0.059203f
C46 VDD1.n0 B 0.471881f
C47 VDD1.t3 B 0.059203f
C48 VDD1.t1 B 0.059203f
C49 VDD1.n1 B 0.694199f
C50 VP.n0 B 0.021218f
C51 VP.t3 B 0.334378f
C52 VP.n1 B 0.030974f
C53 VP.t0 B 0.404173f
C54 VP.t1 B 0.403525f
C55 VP.n2 B 0.916844f
C56 VP.n3 B 0.931419f
C57 VP.t2 B 0.334378f
C58 VP.n4 B 0.176163f
C59 VP.n5 B 0.024511f
C60 VP.n6 B 0.021218f
C61 VP.n7 B 0.021218f
C62 VP.n8 B 0.021218f
C63 VP.n9 B 0.030974f
C64 VP.n10 B 0.024511f
C65 VP.n11 B 0.176163f
C66 VP.n12 B 0.02064f
.ends

