* NGSPICE file created from diff_pair_sample_1364.ext - technology: sky130A

.subckt diff_pair_sample_1364 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0 ps=0 w=2.08 l=0.3
X1 VDD2.t7 VN.t0 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X2 VDD1.t7 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X3 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0.3432 ps=2.41 w=2.08 l=0.3
X4 VTAIL.t14 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X5 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0 ps=0 w=2.08 l=0.3
X7 VDD2.t5 VN.t2 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X8 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X9 VTAIL.t11 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0.3432 ps=2.41 w=2.08 l=0.3
X10 VDD2.t3 VN.t4 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.8112 ps=4.94 w=2.08 l=0.3
X11 VDD1.t3 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.8112 ps=4.94 w=2.08 l=0.3
X12 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X13 VTAIL.t8 VN.t5 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0.3432 ps=2.41 w=2.08 l=0.3
X14 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0.3432 ps=2.41 w=2.08 l=0.3
X15 VTAIL.t15 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.3432 ps=2.41 w=2.08 l=0.3
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0 ps=0 w=2.08 l=0.3
X17 VDD2.t0 VN.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.8112 ps=4.94 w=2.08 l=0.3
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8112 pd=4.94 as=0 ps=0 w=2.08 l=0.3
X19 VDD1.t0 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3432 pd=2.41 as=0.8112 ps=4.94 w=2.08 l=0.3
R0 B.n322 B.n321 585
R1 B.n122 B.n51 585
R2 B.n121 B.n120 585
R3 B.n119 B.n118 585
R4 B.n117 B.n116 585
R5 B.n115 B.n114 585
R6 B.n113 B.n112 585
R7 B.n111 B.n110 585
R8 B.n109 B.n108 585
R9 B.n107 B.n106 585
R10 B.n105 B.n104 585
R11 B.n103 B.n102 585
R12 B.n101 B.n100 585
R13 B.n99 B.n98 585
R14 B.n97 B.n96 585
R15 B.n95 B.n94 585
R16 B.n93 B.n92 585
R17 B.n91 B.n90 585
R18 B.n89 B.n88 585
R19 B.n87 B.n86 585
R20 B.n85 B.n84 585
R21 B.n83 B.n82 585
R22 B.n81 B.n80 585
R23 B.n79 B.n78 585
R24 B.n77 B.n76 585
R25 B.n75 B.n74 585
R26 B.n73 B.n72 585
R27 B.n71 B.n70 585
R28 B.n69 B.n68 585
R29 B.n67 B.n66 585
R30 B.n65 B.n64 585
R31 B.n63 B.n62 585
R32 B.n61 B.n60 585
R33 B.n59 B.n58 585
R34 B.n320 B.n34 585
R35 B.n325 B.n34 585
R36 B.n319 B.n33 585
R37 B.n326 B.n33 585
R38 B.n318 B.n317 585
R39 B.n317 B.n29 585
R40 B.n316 B.n28 585
R41 B.n332 B.n28 585
R42 B.n315 B.n27 585
R43 B.n333 B.n27 585
R44 B.n314 B.n26 585
R45 B.n334 B.n26 585
R46 B.n313 B.n312 585
R47 B.n312 B.n22 585
R48 B.n311 B.n21 585
R49 B.n340 B.n21 585
R50 B.n310 B.n20 585
R51 B.n341 B.n20 585
R52 B.n309 B.n19 585
R53 B.n342 B.n19 585
R54 B.n308 B.n307 585
R55 B.n307 B.n15 585
R56 B.n306 B.n14 585
R57 B.n348 B.n14 585
R58 B.n305 B.n13 585
R59 B.n349 B.n13 585
R60 B.n304 B.n12 585
R61 B.n350 B.n12 585
R62 B.n303 B.n302 585
R63 B.n302 B.n301 585
R64 B.n300 B.n299 585
R65 B.n300 B.n8 585
R66 B.n298 B.n7 585
R67 B.n357 B.n7 585
R68 B.n297 B.n6 585
R69 B.n358 B.n6 585
R70 B.n296 B.n5 585
R71 B.n359 B.n5 585
R72 B.n295 B.n294 585
R73 B.n294 B.n4 585
R74 B.n293 B.n123 585
R75 B.n293 B.n292 585
R76 B.n282 B.n124 585
R77 B.n285 B.n124 585
R78 B.n284 B.n283 585
R79 B.n286 B.n284 585
R80 B.n281 B.n129 585
R81 B.n129 B.n128 585
R82 B.n280 B.n279 585
R83 B.n279 B.n278 585
R84 B.n131 B.n130 585
R85 B.n132 B.n131 585
R86 B.n271 B.n270 585
R87 B.n272 B.n271 585
R88 B.n269 B.n137 585
R89 B.n137 B.n136 585
R90 B.n268 B.n267 585
R91 B.n267 B.n266 585
R92 B.n139 B.n138 585
R93 B.n140 B.n139 585
R94 B.n259 B.n258 585
R95 B.n260 B.n259 585
R96 B.n257 B.n144 585
R97 B.n148 B.n144 585
R98 B.n256 B.n255 585
R99 B.n255 B.n254 585
R100 B.n146 B.n145 585
R101 B.n147 B.n146 585
R102 B.n247 B.n246 585
R103 B.n248 B.n247 585
R104 B.n245 B.n153 585
R105 B.n153 B.n152 585
R106 B.n240 B.n239 585
R107 B.n238 B.n172 585
R108 B.n237 B.n171 585
R109 B.n242 B.n171 585
R110 B.n236 B.n235 585
R111 B.n234 B.n233 585
R112 B.n232 B.n231 585
R113 B.n230 B.n229 585
R114 B.n228 B.n227 585
R115 B.n226 B.n225 585
R116 B.n224 B.n223 585
R117 B.n222 B.n221 585
R118 B.n220 B.n219 585
R119 B.n217 B.n216 585
R120 B.n215 B.n214 585
R121 B.n213 B.n212 585
R122 B.n211 B.n210 585
R123 B.n209 B.n208 585
R124 B.n207 B.n206 585
R125 B.n205 B.n204 585
R126 B.n203 B.n202 585
R127 B.n201 B.n200 585
R128 B.n199 B.n198 585
R129 B.n196 B.n195 585
R130 B.n194 B.n193 585
R131 B.n192 B.n191 585
R132 B.n190 B.n189 585
R133 B.n188 B.n187 585
R134 B.n186 B.n185 585
R135 B.n184 B.n183 585
R136 B.n182 B.n181 585
R137 B.n180 B.n179 585
R138 B.n178 B.n177 585
R139 B.n155 B.n154 585
R140 B.n244 B.n243 585
R141 B.n243 B.n242 585
R142 B.n151 B.n150 585
R143 B.n152 B.n151 585
R144 B.n250 B.n249 585
R145 B.n249 B.n248 585
R146 B.n251 B.n149 585
R147 B.n149 B.n147 585
R148 B.n253 B.n252 585
R149 B.n254 B.n253 585
R150 B.n143 B.n142 585
R151 B.n148 B.n143 585
R152 B.n262 B.n261 585
R153 B.n261 B.n260 585
R154 B.n263 B.n141 585
R155 B.n141 B.n140 585
R156 B.n265 B.n264 585
R157 B.n266 B.n265 585
R158 B.n135 B.n134 585
R159 B.n136 B.n135 585
R160 B.n274 B.n273 585
R161 B.n273 B.n272 585
R162 B.n275 B.n133 585
R163 B.n133 B.n132 585
R164 B.n277 B.n276 585
R165 B.n278 B.n277 585
R166 B.n127 B.n126 585
R167 B.n128 B.n127 585
R168 B.n288 B.n287 585
R169 B.n287 B.n286 585
R170 B.n289 B.n125 585
R171 B.n285 B.n125 585
R172 B.n291 B.n290 585
R173 B.n292 B.n291 585
R174 B.n3 B.n0 585
R175 B.n4 B.n3 585
R176 B.n356 B.n1 585
R177 B.n357 B.n356 585
R178 B.n355 B.n354 585
R179 B.n355 B.n8 585
R180 B.n353 B.n9 585
R181 B.n301 B.n9 585
R182 B.n352 B.n351 585
R183 B.n351 B.n350 585
R184 B.n11 B.n10 585
R185 B.n349 B.n11 585
R186 B.n347 B.n346 585
R187 B.n348 B.n347 585
R188 B.n345 B.n16 585
R189 B.n16 B.n15 585
R190 B.n344 B.n343 585
R191 B.n343 B.n342 585
R192 B.n18 B.n17 585
R193 B.n341 B.n18 585
R194 B.n339 B.n338 585
R195 B.n340 B.n339 585
R196 B.n337 B.n23 585
R197 B.n23 B.n22 585
R198 B.n336 B.n335 585
R199 B.n335 B.n334 585
R200 B.n25 B.n24 585
R201 B.n333 B.n25 585
R202 B.n331 B.n330 585
R203 B.n332 B.n331 585
R204 B.n329 B.n30 585
R205 B.n30 B.n29 585
R206 B.n328 B.n327 585
R207 B.n327 B.n326 585
R208 B.n32 B.n31 585
R209 B.n325 B.n32 585
R210 B.n360 B.n359 585
R211 B.n358 B.n2 585
R212 B.n58 B.n32 516.524
R213 B.n322 B.n34 516.524
R214 B.n243 B.n153 516.524
R215 B.n240 B.n151 516.524
R216 B.n55 B.t8 383.361
R217 B.n52 B.t19 383.361
R218 B.n175 B.t12 383.361
R219 B.n173 B.t16 383.361
R220 B.n324 B.n323 256.663
R221 B.n324 B.n50 256.663
R222 B.n324 B.n49 256.663
R223 B.n324 B.n48 256.663
R224 B.n324 B.n47 256.663
R225 B.n324 B.n46 256.663
R226 B.n324 B.n45 256.663
R227 B.n324 B.n44 256.663
R228 B.n324 B.n43 256.663
R229 B.n324 B.n42 256.663
R230 B.n324 B.n41 256.663
R231 B.n324 B.n40 256.663
R232 B.n324 B.n39 256.663
R233 B.n324 B.n38 256.663
R234 B.n324 B.n37 256.663
R235 B.n324 B.n36 256.663
R236 B.n324 B.n35 256.663
R237 B.n242 B.n241 256.663
R238 B.n242 B.n156 256.663
R239 B.n242 B.n157 256.663
R240 B.n242 B.n158 256.663
R241 B.n242 B.n159 256.663
R242 B.n242 B.n160 256.663
R243 B.n242 B.n161 256.663
R244 B.n242 B.n162 256.663
R245 B.n242 B.n163 256.663
R246 B.n242 B.n164 256.663
R247 B.n242 B.n165 256.663
R248 B.n242 B.n166 256.663
R249 B.n242 B.n167 256.663
R250 B.n242 B.n168 256.663
R251 B.n242 B.n169 256.663
R252 B.n242 B.n170 256.663
R253 B.n362 B.n361 256.663
R254 B.n242 B.n152 171.993
R255 B.n325 B.n324 171.993
R256 B.n62 B.n61 163.367
R257 B.n66 B.n65 163.367
R258 B.n70 B.n69 163.367
R259 B.n74 B.n73 163.367
R260 B.n78 B.n77 163.367
R261 B.n82 B.n81 163.367
R262 B.n86 B.n85 163.367
R263 B.n90 B.n89 163.367
R264 B.n94 B.n93 163.367
R265 B.n98 B.n97 163.367
R266 B.n102 B.n101 163.367
R267 B.n106 B.n105 163.367
R268 B.n110 B.n109 163.367
R269 B.n114 B.n113 163.367
R270 B.n118 B.n117 163.367
R271 B.n120 B.n51 163.367
R272 B.n247 B.n153 163.367
R273 B.n247 B.n146 163.367
R274 B.n255 B.n146 163.367
R275 B.n255 B.n144 163.367
R276 B.n259 B.n144 163.367
R277 B.n259 B.n139 163.367
R278 B.n267 B.n139 163.367
R279 B.n267 B.n137 163.367
R280 B.n271 B.n137 163.367
R281 B.n271 B.n131 163.367
R282 B.n279 B.n131 163.367
R283 B.n279 B.n129 163.367
R284 B.n284 B.n129 163.367
R285 B.n284 B.n124 163.367
R286 B.n293 B.n124 163.367
R287 B.n294 B.n293 163.367
R288 B.n294 B.n5 163.367
R289 B.n6 B.n5 163.367
R290 B.n7 B.n6 163.367
R291 B.n300 B.n7 163.367
R292 B.n302 B.n300 163.367
R293 B.n302 B.n12 163.367
R294 B.n13 B.n12 163.367
R295 B.n14 B.n13 163.367
R296 B.n307 B.n14 163.367
R297 B.n307 B.n19 163.367
R298 B.n20 B.n19 163.367
R299 B.n21 B.n20 163.367
R300 B.n312 B.n21 163.367
R301 B.n312 B.n26 163.367
R302 B.n27 B.n26 163.367
R303 B.n28 B.n27 163.367
R304 B.n317 B.n28 163.367
R305 B.n317 B.n33 163.367
R306 B.n34 B.n33 163.367
R307 B.n172 B.n171 163.367
R308 B.n235 B.n171 163.367
R309 B.n233 B.n232 163.367
R310 B.n229 B.n228 163.367
R311 B.n225 B.n224 163.367
R312 B.n221 B.n220 163.367
R313 B.n216 B.n215 163.367
R314 B.n212 B.n211 163.367
R315 B.n208 B.n207 163.367
R316 B.n204 B.n203 163.367
R317 B.n200 B.n199 163.367
R318 B.n195 B.n194 163.367
R319 B.n191 B.n190 163.367
R320 B.n187 B.n186 163.367
R321 B.n183 B.n182 163.367
R322 B.n179 B.n178 163.367
R323 B.n243 B.n155 163.367
R324 B.n249 B.n151 163.367
R325 B.n249 B.n149 163.367
R326 B.n253 B.n149 163.367
R327 B.n253 B.n143 163.367
R328 B.n261 B.n143 163.367
R329 B.n261 B.n141 163.367
R330 B.n265 B.n141 163.367
R331 B.n265 B.n135 163.367
R332 B.n273 B.n135 163.367
R333 B.n273 B.n133 163.367
R334 B.n277 B.n133 163.367
R335 B.n277 B.n127 163.367
R336 B.n287 B.n127 163.367
R337 B.n287 B.n125 163.367
R338 B.n291 B.n125 163.367
R339 B.n291 B.n3 163.367
R340 B.n360 B.n3 163.367
R341 B.n356 B.n2 163.367
R342 B.n356 B.n355 163.367
R343 B.n355 B.n9 163.367
R344 B.n351 B.n9 163.367
R345 B.n351 B.n11 163.367
R346 B.n347 B.n11 163.367
R347 B.n347 B.n16 163.367
R348 B.n343 B.n16 163.367
R349 B.n343 B.n18 163.367
R350 B.n339 B.n18 163.367
R351 B.n339 B.n23 163.367
R352 B.n335 B.n23 163.367
R353 B.n335 B.n25 163.367
R354 B.n331 B.n25 163.367
R355 B.n331 B.n30 163.367
R356 B.n327 B.n30 163.367
R357 B.n327 B.n32 163.367
R358 B.n248 B.n152 101.701
R359 B.n248 B.n147 101.701
R360 B.n254 B.n147 101.701
R361 B.n254 B.n148 101.701
R362 B.n260 B.n140 101.701
R363 B.n266 B.n140 101.701
R364 B.n266 B.n136 101.701
R365 B.n272 B.n136 101.701
R366 B.n278 B.n132 101.701
R367 B.n286 B.n128 101.701
R368 B.n292 B.n4 101.701
R369 B.n359 B.n4 101.701
R370 B.n359 B.n358 101.701
R371 B.n358 B.n357 101.701
R372 B.n357 B.n8 101.701
R373 B.n350 B.n349 101.701
R374 B.n348 B.n15 101.701
R375 B.n342 B.n341 101.701
R376 B.n341 B.n340 101.701
R377 B.n340 B.n22 101.701
R378 B.n334 B.n22 101.701
R379 B.n333 B.n332 101.701
R380 B.n332 B.n29 101.701
R381 B.n326 B.n29 101.701
R382 B.n326 B.n325 101.701
R383 B.n285 B.t5 98.7089
R384 B.n301 B.t2 98.7089
R385 B.n52 B.t20 96.1179
R386 B.n175 B.t15 96.1179
R387 B.n55 B.t10 96.1176
R388 B.n173 B.t18 96.1176
R389 B.t1 B.n285 89.7354
R390 B.n301 B.t6 89.7354
R391 B.n53 B.t21 83.8997
R392 B.n176 B.t14 83.8997
R393 B.n56 B.t11 83.8994
R394 B.n174 B.t17 83.8994
R395 B.t7 B.n128 74.7796
R396 B.n349 B.t0 74.7796
R397 B.n58 B.n35 71.676
R398 B.n62 B.n36 71.676
R399 B.n66 B.n37 71.676
R400 B.n70 B.n38 71.676
R401 B.n74 B.n39 71.676
R402 B.n78 B.n40 71.676
R403 B.n82 B.n41 71.676
R404 B.n86 B.n42 71.676
R405 B.n90 B.n43 71.676
R406 B.n94 B.n44 71.676
R407 B.n98 B.n45 71.676
R408 B.n102 B.n46 71.676
R409 B.n106 B.n47 71.676
R410 B.n110 B.n48 71.676
R411 B.n114 B.n49 71.676
R412 B.n118 B.n50 71.676
R413 B.n323 B.n51 71.676
R414 B.n323 B.n322 71.676
R415 B.n120 B.n50 71.676
R416 B.n117 B.n49 71.676
R417 B.n113 B.n48 71.676
R418 B.n109 B.n47 71.676
R419 B.n105 B.n46 71.676
R420 B.n101 B.n45 71.676
R421 B.n97 B.n44 71.676
R422 B.n93 B.n43 71.676
R423 B.n89 B.n42 71.676
R424 B.n85 B.n41 71.676
R425 B.n81 B.n40 71.676
R426 B.n77 B.n39 71.676
R427 B.n73 B.n38 71.676
R428 B.n69 B.n37 71.676
R429 B.n65 B.n36 71.676
R430 B.n61 B.n35 71.676
R431 B.n241 B.n240 71.676
R432 B.n235 B.n156 71.676
R433 B.n232 B.n157 71.676
R434 B.n228 B.n158 71.676
R435 B.n224 B.n159 71.676
R436 B.n220 B.n160 71.676
R437 B.n215 B.n161 71.676
R438 B.n211 B.n162 71.676
R439 B.n207 B.n163 71.676
R440 B.n203 B.n164 71.676
R441 B.n199 B.n165 71.676
R442 B.n194 B.n166 71.676
R443 B.n190 B.n167 71.676
R444 B.n186 B.n168 71.676
R445 B.n182 B.n169 71.676
R446 B.n178 B.n170 71.676
R447 B.n241 B.n172 71.676
R448 B.n233 B.n156 71.676
R449 B.n229 B.n157 71.676
R450 B.n225 B.n158 71.676
R451 B.n221 B.n159 71.676
R452 B.n216 B.n160 71.676
R453 B.n212 B.n161 71.676
R454 B.n208 B.n162 71.676
R455 B.n204 B.n163 71.676
R456 B.n200 B.n164 71.676
R457 B.n195 B.n165 71.676
R458 B.n191 B.n166 71.676
R459 B.n187 B.n167 71.676
R460 B.n183 B.n168 71.676
R461 B.n179 B.n169 71.676
R462 B.n170 B.n155 71.676
R463 B.n361 B.n360 71.676
R464 B.n361 B.n2 71.676
R465 B.n260 B.t13 65.8061
R466 B.n334 B.t9 65.8061
R467 B.t4 B.n132 59.8237
R468 B.t3 B.n15 59.8237
R469 B.n57 B.n56 59.5399
R470 B.n54 B.n53 59.5399
R471 B.n197 B.n176 59.5399
R472 B.n218 B.n174 59.5399
R473 B.n272 B.t4 41.8768
R474 B.n342 B.t3 41.8768
R475 B.n148 B.t13 35.8944
R476 B.t9 B.n333 35.8944
R477 B.n239 B.n150 33.5615
R478 B.n245 B.n244 33.5615
R479 B.n321 B.n320 33.5615
R480 B.n59 B.n31 33.5615
R481 B.n278 B.t7 26.921
R482 B.t0 B.n348 26.921
R483 B B.n362 18.0485
R484 B.n56 B.n55 12.2187
R485 B.n53 B.n52 12.2187
R486 B.n176 B.n175 12.2187
R487 B.n174 B.n173 12.2187
R488 B.n286 B.t1 11.9651
R489 B.n350 B.t6 11.9651
R490 B.n250 B.n150 10.6151
R491 B.n251 B.n250 10.6151
R492 B.n252 B.n251 10.6151
R493 B.n252 B.n142 10.6151
R494 B.n262 B.n142 10.6151
R495 B.n263 B.n262 10.6151
R496 B.n264 B.n263 10.6151
R497 B.n264 B.n134 10.6151
R498 B.n274 B.n134 10.6151
R499 B.n275 B.n274 10.6151
R500 B.n276 B.n275 10.6151
R501 B.n276 B.n126 10.6151
R502 B.n288 B.n126 10.6151
R503 B.n289 B.n288 10.6151
R504 B.n290 B.n289 10.6151
R505 B.n290 B.n0 10.6151
R506 B.n239 B.n238 10.6151
R507 B.n238 B.n237 10.6151
R508 B.n237 B.n236 10.6151
R509 B.n236 B.n234 10.6151
R510 B.n234 B.n231 10.6151
R511 B.n231 B.n230 10.6151
R512 B.n230 B.n227 10.6151
R513 B.n227 B.n226 10.6151
R514 B.n226 B.n223 10.6151
R515 B.n223 B.n222 10.6151
R516 B.n222 B.n219 10.6151
R517 B.n217 B.n214 10.6151
R518 B.n214 B.n213 10.6151
R519 B.n213 B.n210 10.6151
R520 B.n210 B.n209 10.6151
R521 B.n209 B.n206 10.6151
R522 B.n206 B.n205 10.6151
R523 B.n205 B.n202 10.6151
R524 B.n202 B.n201 10.6151
R525 B.n201 B.n198 10.6151
R526 B.n196 B.n193 10.6151
R527 B.n193 B.n192 10.6151
R528 B.n192 B.n189 10.6151
R529 B.n189 B.n188 10.6151
R530 B.n188 B.n185 10.6151
R531 B.n185 B.n184 10.6151
R532 B.n184 B.n181 10.6151
R533 B.n181 B.n180 10.6151
R534 B.n180 B.n177 10.6151
R535 B.n177 B.n154 10.6151
R536 B.n244 B.n154 10.6151
R537 B.n246 B.n245 10.6151
R538 B.n246 B.n145 10.6151
R539 B.n256 B.n145 10.6151
R540 B.n257 B.n256 10.6151
R541 B.n258 B.n257 10.6151
R542 B.n258 B.n138 10.6151
R543 B.n268 B.n138 10.6151
R544 B.n269 B.n268 10.6151
R545 B.n270 B.n269 10.6151
R546 B.n270 B.n130 10.6151
R547 B.n280 B.n130 10.6151
R548 B.n281 B.n280 10.6151
R549 B.n283 B.n281 10.6151
R550 B.n283 B.n282 10.6151
R551 B.n282 B.n123 10.6151
R552 B.n295 B.n123 10.6151
R553 B.n296 B.n295 10.6151
R554 B.n297 B.n296 10.6151
R555 B.n298 B.n297 10.6151
R556 B.n299 B.n298 10.6151
R557 B.n303 B.n299 10.6151
R558 B.n304 B.n303 10.6151
R559 B.n305 B.n304 10.6151
R560 B.n306 B.n305 10.6151
R561 B.n308 B.n306 10.6151
R562 B.n309 B.n308 10.6151
R563 B.n310 B.n309 10.6151
R564 B.n311 B.n310 10.6151
R565 B.n313 B.n311 10.6151
R566 B.n314 B.n313 10.6151
R567 B.n315 B.n314 10.6151
R568 B.n316 B.n315 10.6151
R569 B.n318 B.n316 10.6151
R570 B.n319 B.n318 10.6151
R571 B.n320 B.n319 10.6151
R572 B.n354 B.n1 10.6151
R573 B.n354 B.n353 10.6151
R574 B.n353 B.n352 10.6151
R575 B.n352 B.n10 10.6151
R576 B.n346 B.n10 10.6151
R577 B.n346 B.n345 10.6151
R578 B.n345 B.n344 10.6151
R579 B.n344 B.n17 10.6151
R580 B.n338 B.n17 10.6151
R581 B.n338 B.n337 10.6151
R582 B.n337 B.n336 10.6151
R583 B.n336 B.n24 10.6151
R584 B.n330 B.n24 10.6151
R585 B.n330 B.n329 10.6151
R586 B.n329 B.n328 10.6151
R587 B.n328 B.n31 10.6151
R588 B.n60 B.n59 10.6151
R589 B.n63 B.n60 10.6151
R590 B.n64 B.n63 10.6151
R591 B.n67 B.n64 10.6151
R592 B.n68 B.n67 10.6151
R593 B.n71 B.n68 10.6151
R594 B.n72 B.n71 10.6151
R595 B.n75 B.n72 10.6151
R596 B.n76 B.n75 10.6151
R597 B.n79 B.n76 10.6151
R598 B.n80 B.n79 10.6151
R599 B.n84 B.n83 10.6151
R600 B.n87 B.n84 10.6151
R601 B.n88 B.n87 10.6151
R602 B.n91 B.n88 10.6151
R603 B.n92 B.n91 10.6151
R604 B.n95 B.n92 10.6151
R605 B.n96 B.n95 10.6151
R606 B.n99 B.n96 10.6151
R607 B.n100 B.n99 10.6151
R608 B.n104 B.n103 10.6151
R609 B.n107 B.n104 10.6151
R610 B.n108 B.n107 10.6151
R611 B.n111 B.n108 10.6151
R612 B.n112 B.n111 10.6151
R613 B.n115 B.n112 10.6151
R614 B.n116 B.n115 10.6151
R615 B.n119 B.n116 10.6151
R616 B.n121 B.n119 10.6151
R617 B.n122 B.n121 10.6151
R618 B.n321 B.n122 10.6151
R619 B.n219 B.n218 9.36635
R620 B.n197 B.n196 9.36635
R621 B.n80 B.n57 9.36635
R622 B.n103 B.n54 9.36635
R623 B.n362 B.n0 8.11757
R624 B.n362 B.n1 8.11757
R625 B.n292 B.t5 2.99166
R626 B.t2 B.n8 2.99166
R627 B.n218 B.n217 1.24928
R628 B.n198 B.n197 1.24928
R629 B.n83 B.n57 1.24928
R630 B.n100 B.n54 1.24928
R631 VN.n7 VN.t7 300.01
R632 VN.n2 VN.t5 300.01
R633 VN.n16 VN.t3 300.01
R634 VN.n11 VN.t4 300.01
R635 VN.n6 VN.t1 271.527
R636 VN.n1 VN.t2 271.527
R637 VN.n15 VN.t0 271.527
R638 VN.n10 VN.t6 271.527
R639 VN.n12 VN.n11 161.489
R640 VN.n3 VN.n2 161.489
R641 VN.n8 VN.n7 161.3
R642 VN.n17 VN.n16 161.3
R643 VN.n14 VN.n9 161.3
R644 VN.n13 VN.n12 161.3
R645 VN.n5 VN.n0 161.3
R646 VN.n4 VN.n3 161.3
R647 VN.n5 VN.n4 73.0308
R648 VN.n14 VN.n13 73.0308
R649 VN.n2 VN.n1 63.5369
R650 VN.n7 VN.n6 63.5369
R651 VN.n16 VN.n15 63.5369
R652 VN.n11 VN.n10 63.5369
R653 VN VN.n17 33.0024
R654 VN.n4 VN.n1 9.49444
R655 VN.n6 VN.n5 9.49444
R656 VN.n15 VN.n14 9.49444
R657 VN.n13 VN.n10 9.49444
R658 VN.n17 VN.n9 0.189894
R659 VN.n12 VN.n9 0.189894
R660 VN.n3 VN.n0 0.189894
R661 VN.n8 VN.n0 0.189894
R662 VN VN.n8 0.0516364
R663 VTAIL.n15 VTAIL.t13 84.3687
R664 VTAIL.n2 VTAIL.t8 84.3687
R665 VTAIL.n3 VTAIL.t5 84.3687
R666 VTAIL.n6 VTAIL.t4 84.3687
R667 VTAIL.n14 VTAIL.t3 84.3687
R668 VTAIL.n11 VTAIL.t2 84.3685
R669 VTAIL.n10 VTAIL.t9 84.3685
R670 VTAIL.n7 VTAIL.t11 84.3685
R671 VTAIL.n13 VTAIL.n12 74.8495
R672 VTAIL.n9 VTAIL.n8 74.8495
R673 VTAIL.n1 VTAIL.n0 74.8492
R674 VTAIL.n5 VTAIL.n4 74.8492
R675 VTAIL.n15 VTAIL.n14 14.7031
R676 VTAIL.n7 VTAIL.n6 14.7031
R677 VTAIL.n0 VTAIL.t12 9.51973
R678 VTAIL.n0 VTAIL.t14 9.51973
R679 VTAIL.n4 VTAIL.t7 9.51973
R680 VTAIL.n4 VTAIL.t1 9.51973
R681 VTAIL.n12 VTAIL.t6 9.51973
R682 VTAIL.n12 VTAIL.t0 9.51973
R683 VTAIL.n8 VTAIL.t10 9.51973
R684 VTAIL.n8 VTAIL.t15 9.51973
R685 VTAIL.n9 VTAIL.n7 0.543603
R686 VTAIL.n10 VTAIL.n9 0.543603
R687 VTAIL.n13 VTAIL.n11 0.543603
R688 VTAIL.n14 VTAIL.n13 0.543603
R689 VTAIL.n6 VTAIL.n5 0.543603
R690 VTAIL.n5 VTAIL.n3 0.543603
R691 VTAIL.n2 VTAIL.n1 0.543603
R692 VTAIL VTAIL.n15 0.485414
R693 VTAIL.n11 VTAIL.n10 0.470328
R694 VTAIL.n3 VTAIL.n2 0.470328
R695 VTAIL VTAIL.n1 0.0586897
R696 VDD2.n2 VDD2.n1 91.7442
R697 VDD2.n2 VDD2.n0 91.7442
R698 VDD2 VDD2.n5 91.7416
R699 VDD2.n4 VDD2.n3 91.5283
R700 VDD2.n4 VDD2.n2 27.9524
R701 VDD2.n5 VDD2.t1 9.51973
R702 VDD2.n5 VDD2.t3 9.51973
R703 VDD2.n3 VDD2.t4 9.51973
R704 VDD2.n3 VDD2.t7 9.51973
R705 VDD2.n1 VDD2.t6 9.51973
R706 VDD2.n1 VDD2.t0 9.51973
R707 VDD2.n0 VDD2.t2 9.51973
R708 VDD2.n0 VDD2.t5 9.51973
R709 VDD2 VDD2.n4 0.330241
R710 VP.n17 VP.t4 300.01
R711 VP.n11 VP.t6 300.01
R712 VP.n4 VP.t1 300.01
R713 VP.n9 VP.t7 300.01
R714 VP.n16 VP.t2 271.527
R715 VP.n1 VP.t0 271.527
R716 VP.n3 VP.t3 271.527
R717 VP.n8 VP.t5 271.527
R718 VP.n5 VP.n4 161.489
R719 VP.n18 VP.n17 161.3
R720 VP.n6 VP.n5 161.3
R721 VP.n7 VP.n2 161.3
R722 VP.n10 VP.n9 161.3
R723 VP.n15 VP.n0 161.3
R724 VP.n14 VP.n13 161.3
R725 VP.n12 VP.n11 161.3
R726 VP.n15 VP.n14 73.0308
R727 VP.n7 VP.n6 73.0308
R728 VP.n11 VP.n1 63.5369
R729 VP.n17 VP.n16 63.5369
R730 VP.n4 VP.n3 63.5369
R731 VP.n9 VP.n8 63.5369
R732 VP.n12 VP.n10 32.6217
R733 VP.n14 VP.n1 9.49444
R734 VP.n16 VP.n15 9.49444
R735 VP.n6 VP.n3 9.49444
R736 VP.n8 VP.n7 9.49444
R737 VP.n5 VP.n2 0.189894
R738 VP.n10 VP.n2 0.189894
R739 VP.n13 VP.n12 0.189894
R740 VP.n13 VP.n0 0.189894
R741 VP.n18 VP.n0 0.189894
R742 VP VP.n18 0.0516364
R743 VDD1 VDD1.n0 91.858
R744 VDD1.n3 VDD1.n2 91.7442
R745 VDD1.n3 VDD1.n1 91.7442
R746 VDD1.n5 VDD1.n4 91.5282
R747 VDD1.n5 VDD1.n3 28.5354
R748 VDD1.n4 VDD1.t2 9.51973
R749 VDD1.n4 VDD1.t0 9.51973
R750 VDD1.n0 VDD1.t6 9.51973
R751 VDD1.n0 VDD1.t4 9.51973
R752 VDD1.n2 VDD1.t5 9.51973
R753 VDD1.n2 VDD1.t3 9.51973
R754 VDD1.n1 VDD1.t1 9.51973
R755 VDD1.n1 VDD1.t7 9.51973
R756 VDD1 VDD1.n5 0.213862
C0 VDD2 VP 0.281524f
C1 VDD2 VTAIL 4.34813f
C2 VDD2 VN 0.86999f
C3 VDD1 VDD2 0.631433f
C4 VP VTAIL 0.950835f
C5 VP VN 3.02013f
C6 VDD1 VP 0.99709f
C7 VTAIL VN 0.936728f
C8 VDD1 VTAIL 4.30913f
C9 VDD1 VN 0.153505f
C10 VDD2 B 2.222754f
C11 VDD1 B 2.393531f
C12 VTAIL B 2.91821f
C13 VN B 5.288109f
C14 VP B 4.255057f
C15 VDD1.t6 B 0.039703f
C16 VDD1.t4 B 0.039703f
C17 VDD1.n0 B 0.269884f
C18 VDD1.t1 B 0.039703f
C19 VDD1.t7 B 0.039703f
C20 VDD1.n1 B 0.269563f
C21 VDD1.t5 B 0.039703f
C22 VDD1.t3 B 0.039703f
C23 VDD1.n2 B 0.269563f
C24 VDD1.n3 B 1.31036f
C25 VDD1.t2 B 0.039703f
C26 VDD1.t0 B 0.039703f
C27 VDD1.n4 B 0.268993f
C28 VDD1.n5 B 1.30471f
C29 VP.n0 B 0.034505f
C30 VP.t2 B 0.063242f
C31 VP.t0 B 0.063242f
C32 VP.n1 B 0.043322f
C33 VP.n2 B 0.034505f
C34 VP.t5 B 0.063242f
C35 VP.t3 B 0.063242f
C36 VP.n3 B 0.043322f
C37 VP.t1 B 0.067344f
C38 VP.n4 B 0.05337f
C39 VP.n5 B 0.073007f
C40 VP.n6 B 0.012829f
C41 VP.n7 B 0.012829f
C42 VP.n8 B 0.043322f
C43 VP.t7 B 0.067344f
C44 VP.n9 B 0.053325f
C45 VP.n10 B 0.893254f
C46 VP.t6 B 0.067344f
C47 VP.n11 B 0.053325f
C48 VP.n12 B 0.931386f
C49 VP.n13 B 0.034505f
C50 VP.n14 B 0.012829f
C51 VP.n15 B 0.012829f
C52 VP.n16 B 0.043322f
C53 VP.t4 B 0.067344f
C54 VP.n17 B 0.053325f
C55 VP.n18 B 0.02674f
C56 VDD2.t2 B 0.040545f
C57 VDD2.t5 B 0.040545f
C58 VDD2.n0 B 0.275274f
C59 VDD2.t6 B 0.040545f
C60 VDD2.t0 B 0.040545f
C61 VDD2.n1 B 0.275274f
C62 VDD2.n2 B 1.28495f
C63 VDD2.t4 B 0.040545f
C64 VDD2.t7 B 0.040545f
C65 VDD2.n3 B 0.274693f
C66 VDD2.n4 B 1.30367f
C67 VDD2.t1 B 0.040545f
C68 VDD2.t3 B 0.040545f
C69 VDD2.n5 B 0.275259f
C70 VTAIL.t12 B 0.038265f
C71 VTAIL.t14 B 0.038265f
C72 VTAIL.n0 B 0.223671f
C73 VTAIL.n1 B 0.213125f
C74 VTAIL.t8 B 0.295335f
C75 VTAIL.n2 B 0.276698f
C76 VTAIL.t5 B 0.295335f
C77 VTAIL.n3 B 0.276698f
C78 VTAIL.t7 B 0.038265f
C79 VTAIL.t1 B 0.038265f
C80 VTAIL.n4 B 0.223671f
C81 VTAIL.n5 B 0.2495f
C82 VTAIL.t4 B 0.295335f
C83 VTAIL.n6 B 0.732932f
C84 VTAIL.t11 B 0.295337f
C85 VTAIL.n7 B 0.73293f
C86 VTAIL.t10 B 0.038265f
C87 VTAIL.t15 B 0.038265f
C88 VTAIL.n8 B 0.223672f
C89 VTAIL.n9 B 0.249499f
C90 VTAIL.t9 B 0.295337f
C91 VTAIL.n10 B 0.276696f
C92 VTAIL.t2 B 0.295337f
C93 VTAIL.n11 B 0.276696f
C94 VTAIL.t6 B 0.038265f
C95 VTAIL.t0 B 0.038265f
C96 VTAIL.n12 B 0.223672f
C97 VTAIL.n13 B 0.249499f
C98 VTAIL.t3 B 0.295335f
C99 VTAIL.n14 B 0.732932f
C100 VTAIL.t13 B 0.295335f
C101 VTAIL.n15 B 0.728567f
C102 VN.n0 B 0.033956f
C103 VN.t1 B 0.062235f
C104 VN.t2 B 0.062235f
C105 VN.n1 B 0.042632f
C106 VN.t5 B 0.066273f
C107 VN.n2 B 0.052521f
C108 VN.n3 B 0.071846f
C109 VN.n4 B 0.012625f
C110 VN.n5 B 0.012625f
C111 VN.n6 B 0.042632f
C112 VN.t7 B 0.066273f
C113 VN.n7 B 0.052476f
C114 VN.n8 B 0.026315f
C115 VN.n9 B 0.033956f
C116 VN.t3 B 0.066273f
C117 VN.t0 B 0.062235f
C118 VN.t6 B 0.062235f
C119 VN.n10 B 0.042632f
C120 VN.t4 B 0.066273f
C121 VN.n11 B 0.052521f
C122 VN.n12 B 0.071846f
C123 VN.n13 B 0.012625f
C124 VN.n14 B 0.012625f
C125 VN.n15 B 0.042632f
C126 VN.n16 B 0.052476f
C127 VN.n17 B 0.901737f
.ends

