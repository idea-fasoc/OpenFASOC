* NGSPICE file created from diff_pair_sample_0948.ext - technology: sky130A

.subckt diff_pair_sample_0948 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X1 VTAIL.t14 VN.t1 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=2.15655 ps=13.4 w=13.07 l=0.74
X2 VDD2.t4 VN.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=5.0973 ps=26.92 w=13.07 l=0.74
X3 VTAIL.t12 VN.t3 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=2.15655 ps=13.4 w=13.07 l=0.74
X4 VDD2.t2 VN.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X5 VTAIL.t6 VP.t0 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=2.15655 ps=13.4 w=13.07 l=0.74
X6 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=5.0973 ps=26.92 w=13.07 l=0.74
X7 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=5.0973 ps=26.92 w=13.07 l=0.74
X8 VTAIL.t10 VN.t5 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X9 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=0 ps=0 w=13.07 l=0.74
X10 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X11 VTAIL.t2 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=2.15655 ps=13.4 w=13.07 l=0.74
X12 VDD2.t7 VN.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=5.0973 ps=26.92 w=13.07 l=0.74
X13 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=0 ps=0 w=13.07 l=0.74
X14 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X15 VDD2.t6 VN.t7 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X16 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=0 ps=0 w=13.07 l=0.74
X17 VTAIL.t7 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0973 pd=26.92 as=0 ps=0 w=13.07 l=0.74
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.15655 pd=13.4 as=2.15655 ps=13.4 w=13.07 l=0.74
R0 VN.n3 VN.t3 502.736
R1 VN.n13 VN.t6 502.736
R2 VN.n2 VN.t7 479.07
R3 VN.n6 VN.t0 479.07
R4 VN.n8 VN.t2 479.07
R5 VN.n12 VN.t5 479.07
R6 VN.n16 VN.t4 479.07
R7 VN.n18 VN.t1 479.07
R8 VN.n9 VN.n8 161.3
R9 VN.n19 VN.n18 161.3
R10 VN.n17 VN.n10 161.3
R11 VN.n16 VN.n15 161.3
R12 VN.n14 VN.n11 161.3
R13 VN.n7 VN.n0 161.3
R14 VN.n6 VN.n5 161.3
R15 VN.n4 VN.n1 161.3
R16 VN.n14 VN.n13 44.9044
R17 VN.n4 VN.n3 44.9044
R18 VN VN.n19 43.4266
R19 VN.n8 VN.n7 34.3247
R20 VN.n18 VN.n17 34.3247
R21 VN.n2 VN.n1 24.1005
R22 VN.n6 VN.n1 24.1005
R23 VN.n16 VN.n11 24.1005
R24 VN.n12 VN.n11 24.1005
R25 VN.n3 VN.n2 17.9645
R26 VN.n13 VN.n12 17.9645
R27 VN.n7 VN.n6 13.8763
R28 VN.n17 VN.n16 13.8763
R29 VN.n19 VN.n10 0.189894
R30 VN.n15 VN.n10 0.189894
R31 VN.n15 VN.n14 0.189894
R32 VN.n5 VN.n4 0.189894
R33 VN.n5 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VDD2.n2 VDD2.n1 66.0422
R37 VDD2.n2 VDD2.n0 66.0422
R38 VDD2 VDD2.n5 66.0394
R39 VDD2.n4 VDD2.n3 65.6376
R40 VDD2.n4 VDD2.n2 39.1334
R41 VDD2.n5 VDD2.t5 1.51542
R42 VDD2.n5 VDD2.t7 1.51542
R43 VDD2.n3 VDD2.t1 1.51542
R44 VDD2.n3 VDD2.t2 1.51542
R45 VDD2.n1 VDD2.t0 1.51542
R46 VDD2.n1 VDD2.t4 1.51542
R47 VDD2.n0 VDD2.t3 1.51542
R48 VDD2.n0 VDD2.t6 1.51542
R49 VDD2 VDD2.n4 0.519897
R50 VTAIL.n11 VTAIL.t2 50.4737
R51 VTAIL.n10 VTAIL.t9 50.4737
R52 VTAIL.n7 VTAIL.t14 50.4737
R53 VTAIL.n15 VTAIL.t13 50.4725
R54 VTAIL.n2 VTAIL.t12 50.4725
R55 VTAIL.n3 VTAIL.t1 50.4725
R56 VTAIL.n6 VTAIL.t6 50.4725
R57 VTAIL.n14 VTAIL.t5 50.4725
R58 VTAIL.n13 VTAIL.n12 48.9588
R59 VTAIL.n9 VTAIL.n8 48.9588
R60 VTAIL.n1 VTAIL.n0 48.9576
R61 VTAIL.n5 VTAIL.n4 48.9576
R62 VTAIL.n15 VTAIL.n14 24.5565
R63 VTAIL.n7 VTAIL.n6 24.5565
R64 VTAIL.n0 VTAIL.t8 1.51542
R65 VTAIL.n0 VTAIL.t15 1.51542
R66 VTAIL.n4 VTAIL.t0 1.51542
R67 VTAIL.n4 VTAIL.t7 1.51542
R68 VTAIL.n12 VTAIL.t3 1.51542
R69 VTAIL.n12 VTAIL.t4 1.51542
R70 VTAIL.n8 VTAIL.t11 1.51542
R71 VTAIL.n8 VTAIL.t10 1.51542
R72 VTAIL.n9 VTAIL.n7 0.922914
R73 VTAIL.n10 VTAIL.n9 0.922914
R74 VTAIL.n13 VTAIL.n11 0.922914
R75 VTAIL.n14 VTAIL.n13 0.922914
R76 VTAIL.n6 VTAIL.n5 0.922914
R77 VTAIL.n5 VTAIL.n3 0.922914
R78 VTAIL.n2 VTAIL.n1 0.922914
R79 VTAIL VTAIL.n15 0.864724
R80 VTAIL.n11 VTAIL.n10 0.470328
R81 VTAIL.n3 VTAIL.n2 0.470328
R82 VTAIL VTAIL.n1 0.0586897
R83 B.n365 B.t12 628.159
R84 B.n371 B.t8 628.159
R85 B.n101 B.t15 628.159
R86 B.n98 B.t19 628.159
R87 B.n700 B.n699 585
R88 B.n701 B.n700 585
R89 B.n296 B.n97 585
R90 B.n295 B.n294 585
R91 B.n293 B.n292 585
R92 B.n291 B.n290 585
R93 B.n289 B.n288 585
R94 B.n287 B.n286 585
R95 B.n285 B.n284 585
R96 B.n283 B.n282 585
R97 B.n281 B.n280 585
R98 B.n279 B.n278 585
R99 B.n277 B.n276 585
R100 B.n275 B.n274 585
R101 B.n273 B.n272 585
R102 B.n271 B.n270 585
R103 B.n269 B.n268 585
R104 B.n267 B.n266 585
R105 B.n265 B.n264 585
R106 B.n263 B.n262 585
R107 B.n261 B.n260 585
R108 B.n259 B.n258 585
R109 B.n257 B.n256 585
R110 B.n255 B.n254 585
R111 B.n253 B.n252 585
R112 B.n251 B.n250 585
R113 B.n249 B.n248 585
R114 B.n247 B.n246 585
R115 B.n245 B.n244 585
R116 B.n243 B.n242 585
R117 B.n241 B.n240 585
R118 B.n239 B.n238 585
R119 B.n237 B.n236 585
R120 B.n235 B.n234 585
R121 B.n233 B.n232 585
R122 B.n231 B.n230 585
R123 B.n229 B.n228 585
R124 B.n227 B.n226 585
R125 B.n225 B.n224 585
R126 B.n223 B.n222 585
R127 B.n221 B.n220 585
R128 B.n219 B.n218 585
R129 B.n217 B.n216 585
R130 B.n215 B.n214 585
R131 B.n213 B.n212 585
R132 B.n211 B.n210 585
R133 B.n209 B.n208 585
R134 B.n207 B.n206 585
R135 B.n205 B.n204 585
R136 B.n203 B.n202 585
R137 B.n201 B.n200 585
R138 B.n199 B.n198 585
R139 B.n197 B.n196 585
R140 B.n195 B.n194 585
R141 B.n193 B.n192 585
R142 B.n190 B.n189 585
R143 B.n188 B.n187 585
R144 B.n186 B.n185 585
R145 B.n184 B.n183 585
R146 B.n182 B.n181 585
R147 B.n180 B.n179 585
R148 B.n178 B.n177 585
R149 B.n176 B.n175 585
R150 B.n174 B.n173 585
R151 B.n172 B.n171 585
R152 B.n170 B.n169 585
R153 B.n168 B.n167 585
R154 B.n166 B.n165 585
R155 B.n164 B.n163 585
R156 B.n162 B.n161 585
R157 B.n160 B.n159 585
R158 B.n158 B.n157 585
R159 B.n156 B.n155 585
R160 B.n154 B.n153 585
R161 B.n152 B.n151 585
R162 B.n150 B.n149 585
R163 B.n148 B.n147 585
R164 B.n146 B.n145 585
R165 B.n144 B.n143 585
R166 B.n142 B.n141 585
R167 B.n140 B.n139 585
R168 B.n138 B.n137 585
R169 B.n136 B.n135 585
R170 B.n134 B.n133 585
R171 B.n132 B.n131 585
R172 B.n130 B.n129 585
R173 B.n128 B.n127 585
R174 B.n126 B.n125 585
R175 B.n124 B.n123 585
R176 B.n122 B.n121 585
R177 B.n120 B.n119 585
R178 B.n118 B.n117 585
R179 B.n116 B.n115 585
R180 B.n114 B.n113 585
R181 B.n112 B.n111 585
R182 B.n110 B.n109 585
R183 B.n108 B.n107 585
R184 B.n106 B.n105 585
R185 B.n104 B.n103 585
R186 B.n46 B.n45 585
R187 B.n698 B.n47 585
R188 B.n702 B.n47 585
R189 B.n697 B.n696 585
R190 B.n696 B.n43 585
R191 B.n695 B.n42 585
R192 B.n708 B.n42 585
R193 B.n694 B.n41 585
R194 B.n709 B.n41 585
R195 B.n693 B.n40 585
R196 B.n710 B.n40 585
R197 B.n692 B.n691 585
R198 B.n691 B.n39 585
R199 B.n690 B.n35 585
R200 B.n716 B.n35 585
R201 B.n689 B.n34 585
R202 B.n717 B.n34 585
R203 B.n688 B.n33 585
R204 B.n718 B.n33 585
R205 B.n687 B.n686 585
R206 B.n686 B.n29 585
R207 B.n685 B.n28 585
R208 B.n724 B.n28 585
R209 B.n684 B.n27 585
R210 B.n725 B.n27 585
R211 B.n683 B.n26 585
R212 B.n726 B.n26 585
R213 B.n682 B.n681 585
R214 B.n681 B.n22 585
R215 B.n680 B.n21 585
R216 B.n732 B.n21 585
R217 B.n679 B.n20 585
R218 B.n733 B.n20 585
R219 B.n678 B.n19 585
R220 B.n734 B.n19 585
R221 B.n677 B.n676 585
R222 B.n676 B.n18 585
R223 B.n675 B.n14 585
R224 B.n740 B.n14 585
R225 B.n674 B.n13 585
R226 B.n741 B.n13 585
R227 B.n673 B.n12 585
R228 B.n742 B.n12 585
R229 B.n672 B.n671 585
R230 B.n671 B.n8 585
R231 B.n670 B.n7 585
R232 B.n748 B.n7 585
R233 B.n669 B.n6 585
R234 B.n749 B.n6 585
R235 B.n668 B.n5 585
R236 B.n750 B.n5 585
R237 B.n667 B.n666 585
R238 B.n666 B.n4 585
R239 B.n665 B.n297 585
R240 B.n665 B.n664 585
R241 B.n655 B.n298 585
R242 B.n299 B.n298 585
R243 B.n657 B.n656 585
R244 B.n658 B.n657 585
R245 B.n654 B.n304 585
R246 B.n304 B.n303 585
R247 B.n653 B.n652 585
R248 B.n652 B.n651 585
R249 B.n306 B.n305 585
R250 B.n644 B.n306 585
R251 B.n643 B.n642 585
R252 B.n645 B.n643 585
R253 B.n641 B.n311 585
R254 B.n311 B.n310 585
R255 B.n640 B.n639 585
R256 B.n639 B.n638 585
R257 B.n313 B.n312 585
R258 B.n314 B.n313 585
R259 B.n631 B.n630 585
R260 B.n632 B.n631 585
R261 B.n629 B.n318 585
R262 B.n322 B.n318 585
R263 B.n628 B.n627 585
R264 B.n627 B.n626 585
R265 B.n320 B.n319 585
R266 B.n321 B.n320 585
R267 B.n619 B.n618 585
R268 B.n620 B.n619 585
R269 B.n617 B.n327 585
R270 B.n327 B.n326 585
R271 B.n616 B.n615 585
R272 B.n615 B.n614 585
R273 B.n329 B.n328 585
R274 B.n607 B.n329 585
R275 B.n606 B.n605 585
R276 B.n608 B.n606 585
R277 B.n604 B.n334 585
R278 B.n334 B.n333 585
R279 B.n603 B.n602 585
R280 B.n602 B.n601 585
R281 B.n336 B.n335 585
R282 B.n337 B.n336 585
R283 B.n594 B.n593 585
R284 B.n595 B.n594 585
R285 B.n340 B.n339 585
R286 B.n398 B.n397 585
R287 B.n399 B.n395 585
R288 B.n395 B.n341 585
R289 B.n401 B.n400 585
R290 B.n403 B.n394 585
R291 B.n406 B.n405 585
R292 B.n407 B.n393 585
R293 B.n409 B.n408 585
R294 B.n411 B.n392 585
R295 B.n414 B.n413 585
R296 B.n415 B.n391 585
R297 B.n417 B.n416 585
R298 B.n419 B.n390 585
R299 B.n422 B.n421 585
R300 B.n423 B.n389 585
R301 B.n425 B.n424 585
R302 B.n427 B.n388 585
R303 B.n430 B.n429 585
R304 B.n431 B.n387 585
R305 B.n433 B.n432 585
R306 B.n435 B.n386 585
R307 B.n438 B.n437 585
R308 B.n439 B.n385 585
R309 B.n441 B.n440 585
R310 B.n443 B.n384 585
R311 B.n446 B.n445 585
R312 B.n447 B.n383 585
R313 B.n449 B.n448 585
R314 B.n451 B.n382 585
R315 B.n454 B.n453 585
R316 B.n455 B.n381 585
R317 B.n457 B.n456 585
R318 B.n459 B.n380 585
R319 B.n462 B.n461 585
R320 B.n463 B.n379 585
R321 B.n465 B.n464 585
R322 B.n467 B.n378 585
R323 B.n470 B.n469 585
R324 B.n471 B.n377 585
R325 B.n473 B.n472 585
R326 B.n475 B.n376 585
R327 B.n478 B.n477 585
R328 B.n479 B.n375 585
R329 B.n481 B.n480 585
R330 B.n483 B.n374 585
R331 B.n486 B.n485 585
R332 B.n487 B.n370 585
R333 B.n489 B.n488 585
R334 B.n491 B.n369 585
R335 B.n494 B.n493 585
R336 B.n495 B.n368 585
R337 B.n497 B.n496 585
R338 B.n499 B.n367 585
R339 B.n502 B.n501 585
R340 B.n504 B.n364 585
R341 B.n506 B.n505 585
R342 B.n508 B.n363 585
R343 B.n511 B.n510 585
R344 B.n512 B.n362 585
R345 B.n514 B.n513 585
R346 B.n516 B.n361 585
R347 B.n519 B.n518 585
R348 B.n520 B.n360 585
R349 B.n522 B.n521 585
R350 B.n524 B.n359 585
R351 B.n527 B.n526 585
R352 B.n528 B.n358 585
R353 B.n530 B.n529 585
R354 B.n532 B.n357 585
R355 B.n535 B.n534 585
R356 B.n536 B.n356 585
R357 B.n538 B.n537 585
R358 B.n540 B.n355 585
R359 B.n543 B.n542 585
R360 B.n544 B.n354 585
R361 B.n546 B.n545 585
R362 B.n548 B.n353 585
R363 B.n551 B.n550 585
R364 B.n552 B.n352 585
R365 B.n554 B.n553 585
R366 B.n556 B.n351 585
R367 B.n559 B.n558 585
R368 B.n560 B.n350 585
R369 B.n562 B.n561 585
R370 B.n564 B.n349 585
R371 B.n567 B.n566 585
R372 B.n568 B.n348 585
R373 B.n570 B.n569 585
R374 B.n572 B.n347 585
R375 B.n575 B.n574 585
R376 B.n576 B.n346 585
R377 B.n578 B.n577 585
R378 B.n580 B.n345 585
R379 B.n583 B.n582 585
R380 B.n584 B.n344 585
R381 B.n586 B.n585 585
R382 B.n588 B.n343 585
R383 B.n591 B.n590 585
R384 B.n592 B.n342 585
R385 B.n597 B.n596 585
R386 B.n596 B.n595 585
R387 B.n598 B.n338 585
R388 B.n338 B.n337 585
R389 B.n600 B.n599 585
R390 B.n601 B.n600 585
R391 B.n332 B.n331 585
R392 B.n333 B.n332 585
R393 B.n610 B.n609 585
R394 B.n609 B.n608 585
R395 B.n611 B.n330 585
R396 B.n607 B.n330 585
R397 B.n613 B.n612 585
R398 B.n614 B.n613 585
R399 B.n325 B.n324 585
R400 B.n326 B.n325 585
R401 B.n622 B.n621 585
R402 B.n621 B.n620 585
R403 B.n623 B.n323 585
R404 B.n323 B.n321 585
R405 B.n625 B.n624 585
R406 B.n626 B.n625 585
R407 B.n317 B.n316 585
R408 B.n322 B.n317 585
R409 B.n634 B.n633 585
R410 B.n633 B.n632 585
R411 B.n635 B.n315 585
R412 B.n315 B.n314 585
R413 B.n637 B.n636 585
R414 B.n638 B.n637 585
R415 B.n309 B.n308 585
R416 B.n310 B.n309 585
R417 B.n647 B.n646 585
R418 B.n646 B.n645 585
R419 B.n648 B.n307 585
R420 B.n644 B.n307 585
R421 B.n650 B.n649 585
R422 B.n651 B.n650 585
R423 B.n302 B.n301 585
R424 B.n303 B.n302 585
R425 B.n660 B.n659 585
R426 B.n659 B.n658 585
R427 B.n661 B.n300 585
R428 B.n300 B.n299 585
R429 B.n663 B.n662 585
R430 B.n664 B.n663 585
R431 B.n2 B.n0 585
R432 B.n4 B.n2 585
R433 B.n3 B.n1 585
R434 B.n749 B.n3 585
R435 B.n747 B.n746 585
R436 B.n748 B.n747 585
R437 B.n745 B.n9 585
R438 B.n9 B.n8 585
R439 B.n744 B.n743 585
R440 B.n743 B.n742 585
R441 B.n11 B.n10 585
R442 B.n741 B.n11 585
R443 B.n739 B.n738 585
R444 B.n740 B.n739 585
R445 B.n737 B.n15 585
R446 B.n18 B.n15 585
R447 B.n736 B.n735 585
R448 B.n735 B.n734 585
R449 B.n17 B.n16 585
R450 B.n733 B.n17 585
R451 B.n731 B.n730 585
R452 B.n732 B.n731 585
R453 B.n729 B.n23 585
R454 B.n23 B.n22 585
R455 B.n728 B.n727 585
R456 B.n727 B.n726 585
R457 B.n25 B.n24 585
R458 B.n725 B.n25 585
R459 B.n723 B.n722 585
R460 B.n724 B.n723 585
R461 B.n721 B.n30 585
R462 B.n30 B.n29 585
R463 B.n720 B.n719 585
R464 B.n719 B.n718 585
R465 B.n32 B.n31 585
R466 B.n717 B.n32 585
R467 B.n715 B.n714 585
R468 B.n716 B.n715 585
R469 B.n713 B.n36 585
R470 B.n39 B.n36 585
R471 B.n712 B.n711 585
R472 B.n711 B.n710 585
R473 B.n38 B.n37 585
R474 B.n709 B.n38 585
R475 B.n707 B.n706 585
R476 B.n708 B.n707 585
R477 B.n705 B.n44 585
R478 B.n44 B.n43 585
R479 B.n704 B.n703 585
R480 B.n703 B.n702 585
R481 B.n752 B.n751 585
R482 B.n751 B.n750 585
R483 B.n596 B.n340 482.89
R484 B.n703 B.n46 482.89
R485 B.n594 B.n342 482.89
R486 B.n700 B.n47 482.89
R487 B.n701 B.n96 256.663
R488 B.n701 B.n95 256.663
R489 B.n701 B.n94 256.663
R490 B.n701 B.n93 256.663
R491 B.n701 B.n92 256.663
R492 B.n701 B.n91 256.663
R493 B.n701 B.n90 256.663
R494 B.n701 B.n89 256.663
R495 B.n701 B.n88 256.663
R496 B.n701 B.n87 256.663
R497 B.n701 B.n86 256.663
R498 B.n701 B.n85 256.663
R499 B.n701 B.n84 256.663
R500 B.n701 B.n83 256.663
R501 B.n701 B.n82 256.663
R502 B.n701 B.n81 256.663
R503 B.n701 B.n80 256.663
R504 B.n701 B.n79 256.663
R505 B.n701 B.n78 256.663
R506 B.n701 B.n77 256.663
R507 B.n701 B.n76 256.663
R508 B.n701 B.n75 256.663
R509 B.n701 B.n74 256.663
R510 B.n701 B.n73 256.663
R511 B.n701 B.n72 256.663
R512 B.n701 B.n71 256.663
R513 B.n701 B.n70 256.663
R514 B.n701 B.n69 256.663
R515 B.n701 B.n68 256.663
R516 B.n701 B.n67 256.663
R517 B.n701 B.n66 256.663
R518 B.n701 B.n65 256.663
R519 B.n701 B.n64 256.663
R520 B.n701 B.n63 256.663
R521 B.n701 B.n62 256.663
R522 B.n701 B.n61 256.663
R523 B.n701 B.n60 256.663
R524 B.n701 B.n59 256.663
R525 B.n701 B.n58 256.663
R526 B.n701 B.n57 256.663
R527 B.n701 B.n56 256.663
R528 B.n701 B.n55 256.663
R529 B.n701 B.n54 256.663
R530 B.n701 B.n53 256.663
R531 B.n701 B.n52 256.663
R532 B.n701 B.n51 256.663
R533 B.n701 B.n50 256.663
R534 B.n701 B.n49 256.663
R535 B.n701 B.n48 256.663
R536 B.n396 B.n341 256.663
R537 B.n402 B.n341 256.663
R538 B.n404 B.n341 256.663
R539 B.n410 B.n341 256.663
R540 B.n412 B.n341 256.663
R541 B.n418 B.n341 256.663
R542 B.n420 B.n341 256.663
R543 B.n426 B.n341 256.663
R544 B.n428 B.n341 256.663
R545 B.n434 B.n341 256.663
R546 B.n436 B.n341 256.663
R547 B.n442 B.n341 256.663
R548 B.n444 B.n341 256.663
R549 B.n450 B.n341 256.663
R550 B.n452 B.n341 256.663
R551 B.n458 B.n341 256.663
R552 B.n460 B.n341 256.663
R553 B.n466 B.n341 256.663
R554 B.n468 B.n341 256.663
R555 B.n474 B.n341 256.663
R556 B.n476 B.n341 256.663
R557 B.n482 B.n341 256.663
R558 B.n484 B.n341 256.663
R559 B.n490 B.n341 256.663
R560 B.n492 B.n341 256.663
R561 B.n498 B.n341 256.663
R562 B.n500 B.n341 256.663
R563 B.n507 B.n341 256.663
R564 B.n509 B.n341 256.663
R565 B.n515 B.n341 256.663
R566 B.n517 B.n341 256.663
R567 B.n523 B.n341 256.663
R568 B.n525 B.n341 256.663
R569 B.n531 B.n341 256.663
R570 B.n533 B.n341 256.663
R571 B.n539 B.n341 256.663
R572 B.n541 B.n341 256.663
R573 B.n547 B.n341 256.663
R574 B.n549 B.n341 256.663
R575 B.n555 B.n341 256.663
R576 B.n557 B.n341 256.663
R577 B.n563 B.n341 256.663
R578 B.n565 B.n341 256.663
R579 B.n571 B.n341 256.663
R580 B.n573 B.n341 256.663
R581 B.n579 B.n341 256.663
R582 B.n581 B.n341 256.663
R583 B.n587 B.n341 256.663
R584 B.n589 B.n341 256.663
R585 B.n596 B.n338 163.367
R586 B.n600 B.n338 163.367
R587 B.n600 B.n332 163.367
R588 B.n609 B.n332 163.367
R589 B.n609 B.n330 163.367
R590 B.n613 B.n330 163.367
R591 B.n613 B.n325 163.367
R592 B.n621 B.n325 163.367
R593 B.n621 B.n323 163.367
R594 B.n625 B.n323 163.367
R595 B.n625 B.n317 163.367
R596 B.n633 B.n317 163.367
R597 B.n633 B.n315 163.367
R598 B.n637 B.n315 163.367
R599 B.n637 B.n309 163.367
R600 B.n646 B.n309 163.367
R601 B.n646 B.n307 163.367
R602 B.n650 B.n307 163.367
R603 B.n650 B.n302 163.367
R604 B.n659 B.n302 163.367
R605 B.n659 B.n300 163.367
R606 B.n663 B.n300 163.367
R607 B.n663 B.n2 163.367
R608 B.n751 B.n2 163.367
R609 B.n751 B.n3 163.367
R610 B.n747 B.n3 163.367
R611 B.n747 B.n9 163.367
R612 B.n743 B.n9 163.367
R613 B.n743 B.n11 163.367
R614 B.n739 B.n11 163.367
R615 B.n739 B.n15 163.367
R616 B.n735 B.n15 163.367
R617 B.n735 B.n17 163.367
R618 B.n731 B.n17 163.367
R619 B.n731 B.n23 163.367
R620 B.n727 B.n23 163.367
R621 B.n727 B.n25 163.367
R622 B.n723 B.n25 163.367
R623 B.n723 B.n30 163.367
R624 B.n719 B.n30 163.367
R625 B.n719 B.n32 163.367
R626 B.n715 B.n32 163.367
R627 B.n715 B.n36 163.367
R628 B.n711 B.n36 163.367
R629 B.n711 B.n38 163.367
R630 B.n707 B.n38 163.367
R631 B.n707 B.n44 163.367
R632 B.n703 B.n44 163.367
R633 B.n397 B.n395 163.367
R634 B.n401 B.n395 163.367
R635 B.n405 B.n403 163.367
R636 B.n409 B.n393 163.367
R637 B.n413 B.n411 163.367
R638 B.n417 B.n391 163.367
R639 B.n421 B.n419 163.367
R640 B.n425 B.n389 163.367
R641 B.n429 B.n427 163.367
R642 B.n433 B.n387 163.367
R643 B.n437 B.n435 163.367
R644 B.n441 B.n385 163.367
R645 B.n445 B.n443 163.367
R646 B.n449 B.n383 163.367
R647 B.n453 B.n451 163.367
R648 B.n457 B.n381 163.367
R649 B.n461 B.n459 163.367
R650 B.n465 B.n379 163.367
R651 B.n469 B.n467 163.367
R652 B.n473 B.n377 163.367
R653 B.n477 B.n475 163.367
R654 B.n481 B.n375 163.367
R655 B.n485 B.n483 163.367
R656 B.n489 B.n370 163.367
R657 B.n493 B.n491 163.367
R658 B.n497 B.n368 163.367
R659 B.n501 B.n499 163.367
R660 B.n506 B.n364 163.367
R661 B.n510 B.n508 163.367
R662 B.n514 B.n362 163.367
R663 B.n518 B.n516 163.367
R664 B.n522 B.n360 163.367
R665 B.n526 B.n524 163.367
R666 B.n530 B.n358 163.367
R667 B.n534 B.n532 163.367
R668 B.n538 B.n356 163.367
R669 B.n542 B.n540 163.367
R670 B.n546 B.n354 163.367
R671 B.n550 B.n548 163.367
R672 B.n554 B.n352 163.367
R673 B.n558 B.n556 163.367
R674 B.n562 B.n350 163.367
R675 B.n566 B.n564 163.367
R676 B.n570 B.n348 163.367
R677 B.n574 B.n572 163.367
R678 B.n578 B.n346 163.367
R679 B.n582 B.n580 163.367
R680 B.n586 B.n344 163.367
R681 B.n590 B.n588 163.367
R682 B.n594 B.n336 163.367
R683 B.n602 B.n336 163.367
R684 B.n602 B.n334 163.367
R685 B.n606 B.n334 163.367
R686 B.n606 B.n329 163.367
R687 B.n615 B.n329 163.367
R688 B.n615 B.n327 163.367
R689 B.n619 B.n327 163.367
R690 B.n619 B.n320 163.367
R691 B.n627 B.n320 163.367
R692 B.n627 B.n318 163.367
R693 B.n631 B.n318 163.367
R694 B.n631 B.n313 163.367
R695 B.n639 B.n313 163.367
R696 B.n639 B.n311 163.367
R697 B.n643 B.n311 163.367
R698 B.n643 B.n306 163.367
R699 B.n652 B.n306 163.367
R700 B.n652 B.n304 163.367
R701 B.n657 B.n304 163.367
R702 B.n657 B.n298 163.367
R703 B.n665 B.n298 163.367
R704 B.n666 B.n665 163.367
R705 B.n666 B.n5 163.367
R706 B.n6 B.n5 163.367
R707 B.n7 B.n6 163.367
R708 B.n671 B.n7 163.367
R709 B.n671 B.n12 163.367
R710 B.n13 B.n12 163.367
R711 B.n14 B.n13 163.367
R712 B.n676 B.n14 163.367
R713 B.n676 B.n19 163.367
R714 B.n20 B.n19 163.367
R715 B.n21 B.n20 163.367
R716 B.n681 B.n21 163.367
R717 B.n681 B.n26 163.367
R718 B.n27 B.n26 163.367
R719 B.n28 B.n27 163.367
R720 B.n686 B.n28 163.367
R721 B.n686 B.n33 163.367
R722 B.n34 B.n33 163.367
R723 B.n35 B.n34 163.367
R724 B.n691 B.n35 163.367
R725 B.n691 B.n40 163.367
R726 B.n41 B.n40 163.367
R727 B.n42 B.n41 163.367
R728 B.n696 B.n42 163.367
R729 B.n696 B.n47 163.367
R730 B.n105 B.n104 163.367
R731 B.n109 B.n108 163.367
R732 B.n113 B.n112 163.367
R733 B.n117 B.n116 163.367
R734 B.n121 B.n120 163.367
R735 B.n125 B.n124 163.367
R736 B.n129 B.n128 163.367
R737 B.n133 B.n132 163.367
R738 B.n137 B.n136 163.367
R739 B.n141 B.n140 163.367
R740 B.n145 B.n144 163.367
R741 B.n149 B.n148 163.367
R742 B.n153 B.n152 163.367
R743 B.n157 B.n156 163.367
R744 B.n161 B.n160 163.367
R745 B.n165 B.n164 163.367
R746 B.n169 B.n168 163.367
R747 B.n173 B.n172 163.367
R748 B.n177 B.n176 163.367
R749 B.n181 B.n180 163.367
R750 B.n185 B.n184 163.367
R751 B.n189 B.n188 163.367
R752 B.n194 B.n193 163.367
R753 B.n198 B.n197 163.367
R754 B.n202 B.n201 163.367
R755 B.n206 B.n205 163.367
R756 B.n210 B.n209 163.367
R757 B.n214 B.n213 163.367
R758 B.n218 B.n217 163.367
R759 B.n222 B.n221 163.367
R760 B.n226 B.n225 163.367
R761 B.n230 B.n229 163.367
R762 B.n234 B.n233 163.367
R763 B.n238 B.n237 163.367
R764 B.n242 B.n241 163.367
R765 B.n246 B.n245 163.367
R766 B.n250 B.n249 163.367
R767 B.n254 B.n253 163.367
R768 B.n258 B.n257 163.367
R769 B.n262 B.n261 163.367
R770 B.n266 B.n265 163.367
R771 B.n270 B.n269 163.367
R772 B.n274 B.n273 163.367
R773 B.n278 B.n277 163.367
R774 B.n282 B.n281 163.367
R775 B.n286 B.n285 163.367
R776 B.n290 B.n289 163.367
R777 B.n294 B.n293 163.367
R778 B.n700 B.n97 163.367
R779 B.n365 B.t14 91.3169
R780 B.n98 B.t20 91.3169
R781 B.n371 B.t11 91.3002
R782 B.n101 B.t17 91.3002
R783 B.n396 B.n340 71.676
R784 B.n402 B.n401 71.676
R785 B.n405 B.n404 71.676
R786 B.n410 B.n409 71.676
R787 B.n413 B.n412 71.676
R788 B.n418 B.n417 71.676
R789 B.n421 B.n420 71.676
R790 B.n426 B.n425 71.676
R791 B.n429 B.n428 71.676
R792 B.n434 B.n433 71.676
R793 B.n437 B.n436 71.676
R794 B.n442 B.n441 71.676
R795 B.n445 B.n444 71.676
R796 B.n450 B.n449 71.676
R797 B.n453 B.n452 71.676
R798 B.n458 B.n457 71.676
R799 B.n461 B.n460 71.676
R800 B.n466 B.n465 71.676
R801 B.n469 B.n468 71.676
R802 B.n474 B.n473 71.676
R803 B.n477 B.n476 71.676
R804 B.n482 B.n481 71.676
R805 B.n485 B.n484 71.676
R806 B.n490 B.n489 71.676
R807 B.n493 B.n492 71.676
R808 B.n498 B.n497 71.676
R809 B.n501 B.n500 71.676
R810 B.n507 B.n506 71.676
R811 B.n510 B.n509 71.676
R812 B.n515 B.n514 71.676
R813 B.n518 B.n517 71.676
R814 B.n523 B.n522 71.676
R815 B.n526 B.n525 71.676
R816 B.n531 B.n530 71.676
R817 B.n534 B.n533 71.676
R818 B.n539 B.n538 71.676
R819 B.n542 B.n541 71.676
R820 B.n547 B.n546 71.676
R821 B.n550 B.n549 71.676
R822 B.n555 B.n554 71.676
R823 B.n558 B.n557 71.676
R824 B.n563 B.n562 71.676
R825 B.n566 B.n565 71.676
R826 B.n571 B.n570 71.676
R827 B.n574 B.n573 71.676
R828 B.n579 B.n578 71.676
R829 B.n582 B.n581 71.676
R830 B.n587 B.n586 71.676
R831 B.n590 B.n589 71.676
R832 B.n48 B.n46 71.676
R833 B.n105 B.n49 71.676
R834 B.n109 B.n50 71.676
R835 B.n113 B.n51 71.676
R836 B.n117 B.n52 71.676
R837 B.n121 B.n53 71.676
R838 B.n125 B.n54 71.676
R839 B.n129 B.n55 71.676
R840 B.n133 B.n56 71.676
R841 B.n137 B.n57 71.676
R842 B.n141 B.n58 71.676
R843 B.n145 B.n59 71.676
R844 B.n149 B.n60 71.676
R845 B.n153 B.n61 71.676
R846 B.n157 B.n62 71.676
R847 B.n161 B.n63 71.676
R848 B.n165 B.n64 71.676
R849 B.n169 B.n65 71.676
R850 B.n173 B.n66 71.676
R851 B.n177 B.n67 71.676
R852 B.n181 B.n68 71.676
R853 B.n185 B.n69 71.676
R854 B.n189 B.n70 71.676
R855 B.n194 B.n71 71.676
R856 B.n198 B.n72 71.676
R857 B.n202 B.n73 71.676
R858 B.n206 B.n74 71.676
R859 B.n210 B.n75 71.676
R860 B.n214 B.n76 71.676
R861 B.n218 B.n77 71.676
R862 B.n222 B.n78 71.676
R863 B.n226 B.n79 71.676
R864 B.n230 B.n80 71.676
R865 B.n234 B.n81 71.676
R866 B.n238 B.n82 71.676
R867 B.n242 B.n83 71.676
R868 B.n246 B.n84 71.676
R869 B.n250 B.n85 71.676
R870 B.n254 B.n86 71.676
R871 B.n258 B.n87 71.676
R872 B.n262 B.n88 71.676
R873 B.n266 B.n89 71.676
R874 B.n270 B.n90 71.676
R875 B.n274 B.n91 71.676
R876 B.n278 B.n92 71.676
R877 B.n282 B.n93 71.676
R878 B.n286 B.n94 71.676
R879 B.n290 B.n95 71.676
R880 B.n294 B.n96 71.676
R881 B.n97 B.n96 71.676
R882 B.n293 B.n95 71.676
R883 B.n289 B.n94 71.676
R884 B.n285 B.n93 71.676
R885 B.n281 B.n92 71.676
R886 B.n277 B.n91 71.676
R887 B.n273 B.n90 71.676
R888 B.n269 B.n89 71.676
R889 B.n265 B.n88 71.676
R890 B.n261 B.n87 71.676
R891 B.n257 B.n86 71.676
R892 B.n253 B.n85 71.676
R893 B.n249 B.n84 71.676
R894 B.n245 B.n83 71.676
R895 B.n241 B.n82 71.676
R896 B.n237 B.n81 71.676
R897 B.n233 B.n80 71.676
R898 B.n229 B.n79 71.676
R899 B.n225 B.n78 71.676
R900 B.n221 B.n77 71.676
R901 B.n217 B.n76 71.676
R902 B.n213 B.n75 71.676
R903 B.n209 B.n74 71.676
R904 B.n205 B.n73 71.676
R905 B.n201 B.n72 71.676
R906 B.n197 B.n71 71.676
R907 B.n193 B.n70 71.676
R908 B.n188 B.n69 71.676
R909 B.n184 B.n68 71.676
R910 B.n180 B.n67 71.676
R911 B.n176 B.n66 71.676
R912 B.n172 B.n65 71.676
R913 B.n168 B.n64 71.676
R914 B.n164 B.n63 71.676
R915 B.n160 B.n62 71.676
R916 B.n156 B.n61 71.676
R917 B.n152 B.n60 71.676
R918 B.n148 B.n59 71.676
R919 B.n144 B.n58 71.676
R920 B.n140 B.n57 71.676
R921 B.n136 B.n56 71.676
R922 B.n132 B.n55 71.676
R923 B.n128 B.n54 71.676
R924 B.n124 B.n53 71.676
R925 B.n120 B.n52 71.676
R926 B.n116 B.n51 71.676
R927 B.n112 B.n50 71.676
R928 B.n108 B.n49 71.676
R929 B.n104 B.n48 71.676
R930 B.n397 B.n396 71.676
R931 B.n403 B.n402 71.676
R932 B.n404 B.n393 71.676
R933 B.n411 B.n410 71.676
R934 B.n412 B.n391 71.676
R935 B.n419 B.n418 71.676
R936 B.n420 B.n389 71.676
R937 B.n427 B.n426 71.676
R938 B.n428 B.n387 71.676
R939 B.n435 B.n434 71.676
R940 B.n436 B.n385 71.676
R941 B.n443 B.n442 71.676
R942 B.n444 B.n383 71.676
R943 B.n451 B.n450 71.676
R944 B.n452 B.n381 71.676
R945 B.n459 B.n458 71.676
R946 B.n460 B.n379 71.676
R947 B.n467 B.n466 71.676
R948 B.n468 B.n377 71.676
R949 B.n475 B.n474 71.676
R950 B.n476 B.n375 71.676
R951 B.n483 B.n482 71.676
R952 B.n484 B.n370 71.676
R953 B.n491 B.n490 71.676
R954 B.n492 B.n368 71.676
R955 B.n499 B.n498 71.676
R956 B.n500 B.n364 71.676
R957 B.n508 B.n507 71.676
R958 B.n509 B.n362 71.676
R959 B.n516 B.n515 71.676
R960 B.n517 B.n360 71.676
R961 B.n524 B.n523 71.676
R962 B.n525 B.n358 71.676
R963 B.n532 B.n531 71.676
R964 B.n533 B.n356 71.676
R965 B.n540 B.n539 71.676
R966 B.n541 B.n354 71.676
R967 B.n548 B.n547 71.676
R968 B.n549 B.n352 71.676
R969 B.n556 B.n555 71.676
R970 B.n557 B.n350 71.676
R971 B.n564 B.n563 71.676
R972 B.n565 B.n348 71.676
R973 B.n572 B.n571 71.676
R974 B.n573 B.n346 71.676
R975 B.n580 B.n579 71.676
R976 B.n581 B.n344 71.676
R977 B.n588 B.n587 71.676
R978 B.n589 B.n342 71.676
R979 B.n366 B.t13 70.5654
R980 B.n99 B.t21 70.5654
R981 B.n372 B.t10 70.5487
R982 B.n102 B.t18 70.5487
R983 B.n595 B.n341 67.7574
R984 B.n702 B.n701 67.7574
R985 B.n503 B.n366 59.5399
R986 B.n373 B.n372 59.5399
R987 B.n191 B.n102 59.5399
R988 B.n100 B.n99 59.5399
R989 B.n595 B.n337 40.7746
R990 B.n601 B.n337 40.7746
R991 B.n601 B.n333 40.7746
R992 B.n608 B.n333 40.7746
R993 B.n608 B.n607 40.7746
R994 B.n614 B.n326 40.7746
R995 B.n620 B.n326 40.7746
R996 B.n620 B.n321 40.7746
R997 B.n626 B.n321 40.7746
R998 B.n626 B.n322 40.7746
R999 B.n632 B.n314 40.7746
R1000 B.n638 B.n314 40.7746
R1001 B.n645 B.n310 40.7746
R1002 B.n645 B.n644 40.7746
R1003 B.n651 B.n303 40.7746
R1004 B.n658 B.n303 40.7746
R1005 B.n664 B.n299 40.7746
R1006 B.n664 B.n4 40.7746
R1007 B.n750 B.n4 40.7746
R1008 B.n750 B.n749 40.7746
R1009 B.n749 B.n748 40.7746
R1010 B.n748 B.n8 40.7746
R1011 B.n742 B.n741 40.7746
R1012 B.n741 B.n740 40.7746
R1013 B.n734 B.n18 40.7746
R1014 B.n734 B.n733 40.7746
R1015 B.n732 B.n22 40.7746
R1016 B.n726 B.n22 40.7746
R1017 B.n725 B.n724 40.7746
R1018 B.n724 B.n29 40.7746
R1019 B.n718 B.n29 40.7746
R1020 B.n718 B.n717 40.7746
R1021 B.n717 B.n716 40.7746
R1022 B.n710 B.n39 40.7746
R1023 B.n710 B.n709 40.7746
R1024 B.n709 B.n708 40.7746
R1025 B.n708 B.n43 40.7746
R1026 B.n702 B.n43 40.7746
R1027 B.n614 B.t9 39.5753
R1028 B.n716 B.t16 39.5753
R1029 B.n658 B.t1 33.5791
R1030 B.n742 B.t2 33.5791
R1031 B.n704 B.n45 31.3761
R1032 B.n699 B.n698 31.3761
R1033 B.n593 B.n592 31.3761
R1034 B.n597 B.n339 31.3761
R1035 B.n644 B.t7 27.5829
R1036 B.n18 B.t3 27.5829
R1037 B.n632 B.t6 25.1845
R1038 B.n726 B.t5 25.1845
R1039 B.n638 B.t0 21.5868
R1040 B.t4 B.n732 21.5868
R1041 B.n366 B.n365 20.752
R1042 B.n372 B.n371 20.752
R1043 B.n102 B.n101 20.752
R1044 B.n99 B.n98 20.752
R1045 B.t0 B.n310 19.1883
R1046 B.n733 B.t4 19.1883
R1047 B B.n752 18.0485
R1048 B.n322 B.t6 15.5906
R1049 B.t5 B.n725 15.5906
R1050 B.n651 B.t7 13.1921
R1051 B.n740 B.t3 13.1921
R1052 B.n103 B.n45 10.6151
R1053 B.n106 B.n103 10.6151
R1054 B.n107 B.n106 10.6151
R1055 B.n110 B.n107 10.6151
R1056 B.n111 B.n110 10.6151
R1057 B.n114 B.n111 10.6151
R1058 B.n115 B.n114 10.6151
R1059 B.n118 B.n115 10.6151
R1060 B.n119 B.n118 10.6151
R1061 B.n122 B.n119 10.6151
R1062 B.n123 B.n122 10.6151
R1063 B.n126 B.n123 10.6151
R1064 B.n127 B.n126 10.6151
R1065 B.n130 B.n127 10.6151
R1066 B.n131 B.n130 10.6151
R1067 B.n134 B.n131 10.6151
R1068 B.n135 B.n134 10.6151
R1069 B.n138 B.n135 10.6151
R1070 B.n139 B.n138 10.6151
R1071 B.n142 B.n139 10.6151
R1072 B.n143 B.n142 10.6151
R1073 B.n146 B.n143 10.6151
R1074 B.n147 B.n146 10.6151
R1075 B.n150 B.n147 10.6151
R1076 B.n151 B.n150 10.6151
R1077 B.n154 B.n151 10.6151
R1078 B.n155 B.n154 10.6151
R1079 B.n158 B.n155 10.6151
R1080 B.n159 B.n158 10.6151
R1081 B.n162 B.n159 10.6151
R1082 B.n163 B.n162 10.6151
R1083 B.n166 B.n163 10.6151
R1084 B.n167 B.n166 10.6151
R1085 B.n170 B.n167 10.6151
R1086 B.n171 B.n170 10.6151
R1087 B.n174 B.n171 10.6151
R1088 B.n175 B.n174 10.6151
R1089 B.n178 B.n175 10.6151
R1090 B.n179 B.n178 10.6151
R1091 B.n182 B.n179 10.6151
R1092 B.n183 B.n182 10.6151
R1093 B.n186 B.n183 10.6151
R1094 B.n187 B.n186 10.6151
R1095 B.n190 B.n187 10.6151
R1096 B.n195 B.n192 10.6151
R1097 B.n196 B.n195 10.6151
R1098 B.n199 B.n196 10.6151
R1099 B.n200 B.n199 10.6151
R1100 B.n203 B.n200 10.6151
R1101 B.n204 B.n203 10.6151
R1102 B.n207 B.n204 10.6151
R1103 B.n208 B.n207 10.6151
R1104 B.n212 B.n211 10.6151
R1105 B.n215 B.n212 10.6151
R1106 B.n216 B.n215 10.6151
R1107 B.n219 B.n216 10.6151
R1108 B.n220 B.n219 10.6151
R1109 B.n223 B.n220 10.6151
R1110 B.n224 B.n223 10.6151
R1111 B.n227 B.n224 10.6151
R1112 B.n228 B.n227 10.6151
R1113 B.n231 B.n228 10.6151
R1114 B.n232 B.n231 10.6151
R1115 B.n235 B.n232 10.6151
R1116 B.n236 B.n235 10.6151
R1117 B.n239 B.n236 10.6151
R1118 B.n240 B.n239 10.6151
R1119 B.n243 B.n240 10.6151
R1120 B.n244 B.n243 10.6151
R1121 B.n247 B.n244 10.6151
R1122 B.n248 B.n247 10.6151
R1123 B.n251 B.n248 10.6151
R1124 B.n252 B.n251 10.6151
R1125 B.n255 B.n252 10.6151
R1126 B.n256 B.n255 10.6151
R1127 B.n259 B.n256 10.6151
R1128 B.n260 B.n259 10.6151
R1129 B.n263 B.n260 10.6151
R1130 B.n264 B.n263 10.6151
R1131 B.n267 B.n264 10.6151
R1132 B.n268 B.n267 10.6151
R1133 B.n271 B.n268 10.6151
R1134 B.n272 B.n271 10.6151
R1135 B.n275 B.n272 10.6151
R1136 B.n276 B.n275 10.6151
R1137 B.n279 B.n276 10.6151
R1138 B.n280 B.n279 10.6151
R1139 B.n283 B.n280 10.6151
R1140 B.n284 B.n283 10.6151
R1141 B.n287 B.n284 10.6151
R1142 B.n288 B.n287 10.6151
R1143 B.n291 B.n288 10.6151
R1144 B.n292 B.n291 10.6151
R1145 B.n295 B.n292 10.6151
R1146 B.n296 B.n295 10.6151
R1147 B.n699 B.n296 10.6151
R1148 B.n593 B.n335 10.6151
R1149 B.n603 B.n335 10.6151
R1150 B.n604 B.n603 10.6151
R1151 B.n605 B.n604 10.6151
R1152 B.n605 B.n328 10.6151
R1153 B.n616 B.n328 10.6151
R1154 B.n617 B.n616 10.6151
R1155 B.n618 B.n617 10.6151
R1156 B.n618 B.n319 10.6151
R1157 B.n628 B.n319 10.6151
R1158 B.n629 B.n628 10.6151
R1159 B.n630 B.n629 10.6151
R1160 B.n630 B.n312 10.6151
R1161 B.n640 B.n312 10.6151
R1162 B.n641 B.n640 10.6151
R1163 B.n642 B.n641 10.6151
R1164 B.n642 B.n305 10.6151
R1165 B.n653 B.n305 10.6151
R1166 B.n654 B.n653 10.6151
R1167 B.n656 B.n654 10.6151
R1168 B.n656 B.n655 10.6151
R1169 B.n655 B.n297 10.6151
R1170 B.n667 B.n297 10.6151
R1171 B.n668 B.n667 10.6151
R1172 B.n669 B.n668 10.6151
R1173 B.n670 B.n669 10.6151
R1174 B.n672 B.n670 10.6151
R1175 B.n673 B.n672 10.6151
R1176 B.n674 B.n673 10.6151
R1177 B.n675 B.n674 10.6151
R1178 B.n677 B.n675 10.6151
R1179 B.n678 B.n677 10.6151
R1180 B.n679 B.n678 10.6151
R1181 B.n680 B.n679 10.6151
R1182 B.n682 B.n680 10.6151
R1183 B.n683 B.n682 10.6151
R1184 B.n684 B.n683 10.6151
R1185 B.n685 B.n684 10.6151
R1186 B.n687 B.n685 10.6151
R1187 B.n688 B.n687 10.6151
R1188 B.n689 B.n688 10.6151
R1189 B.n690 B.n689 10.6151
R1190 B.n692 B.n690 10.6151
R1191 B.n693 B.n692 10.6151
R1192 B.n694 B.n693 10.6151
R1193 B.n695 B.n694 10.6151
R1194 B.n697 B.n695 10.6151
R1195 B.n698 B.n697 10.6151
R1196 B.n398 B.n339 10.6151
R1197 B.n399 B.n398 10.6151
R1198 B.n400 B.n399 10.6151
R1199 B.n400 B.n394 10.6151
R1200 B.n406 B.n394 10.6151
R1201 B.n407 B.n406 10.6151
R1202 B.n408 B.n407 10.6151
R1203 B.n408 B.n392 10.6151
R1204 B.n414 B.n392 10.6151
R1205 B.n415 B.n414 10.6151
R1206 B.n416 B.n415 10.6151
R1207 B.n416 B.n390 10.6151
R1208 B.n422 B.n390 10.6151
R1209 B.n423 B.n422 10.6151
R1210 B.n424 B.n423 10.6151
R1211 B.n424 B.n388 10.6151
R1212 B.n430 B.n388 10.6151
R1213 B.n431 B.n430 10.6151
R1214 B.n432 B.n431 10.6151
R1215 B.n432 B.n386 10.6151
R1216 B.n438 B.n386 10.6151
R1217 B.n439 B.n438 10.6151
R1218 B.n440 B.n439 10.6151
R1219 B.n440 B.n384 10.6151
R1220 B.n446 B.n384 10.6151
R1221 B.n447 B.n446 10.6151
R1222 B.n448 B.n447 10.6151
R1223 B.n448 B.n382 10.6151
R1224 B.n454 B.n382 10.6151
R1225 B.n455 B.n454 10.6151
R1226 B.n456 B.n455 10.6151
R1227 B.n456 B.n380 10.6151
R1228 B.n462 B.n380 10.6151
R1229 B.n463 B.n462 10.6151
R1230 B.n464 B.n463 10.6151
R1231 B.n464 B.n378 10.6151
R1232 B.n470 B.n378 10.6151
R1233 B.n471 B.n470 10.6151
R1234 B.n472 B.n471 10.6151
R1235 B.n472 B.n376 10.6151
R1236 B.n478 B.n376 10.6151
R1237 B.n479 B.n478 10.6151
R1238 B.n480 B.n479 10.6151
R1239 B.n480 B.n374 10.6151
R1240 B.n487 B.n486 10.6151
R1241 B.n488 B.n487 10.6151
R1242 B.n488 B.n369 10.6151
R1243 B.n494 B.n369 10.6151
R1244 B.n495 B.n494 10.6151
R1245 B.n496 B.n495 10.6151
R1246 B.n496 B.n367 10.6151
R1247 B.n502 B.n367 10.6151
R1248 B.n505 B.n504 10.6151
R1249 B.n505 B.n363 10.6151
R1250 B.n511 B.n363 10.6151
R1251 B.n512 B.n511 10.6151
R1252 B.n513 B.n512 10.6151
R1253 B.n513 B.n361 10.6151
R1254 B.n519 B.n361 10.6151
R1255 B.n520 B.n519 10.6151
R1256 B.n521 B.n520 10.6151
R1257 B.n521 B.n359 10.6151
R1258 B.n527 B.n359 10.6151
R1259 B.n528 B.n527 10.6151
R1260 B.n529 B.n528 10.6151
R1261 B.n529 B.n357 10.6151
R1262 B.n535 B.n357 10.6151
R1263 B.n536 B.n535 10.6151
R1264 B.n537 B.n536 10.6151
R1265 B.n537 B.n355 10.6151
R1266 B.n543 B.n355 10.6151
R1267 B.n544 B.n543 10.6151
R1268 B.n545 B.n544 10.6151
R1269 B.n545 B.n353 10.6151
R1270 B.n551 B.n353 10.6151
R1271 B.n552 B.n551 10.6151
R1272 B.n553 B.n552 10.6151
R1273 B.n553 B.n351 10.6151
R1274 B.n559 B.n351 10.6151
R1275 B.n560 B.n559 10.6151
R1276 B.n561 B.n560 10.6151
R1277 B.n561 B.n349 10.6151
R1278 B.n567 B.n349 10.6151
R1279 B.n568 B.n567 10.6151
R1280 B.n569 B.n568 10.6151
R1281 B.n569 B.n347 10.6151
R1282 B.n575 B.n347 10.6151
R1283 B.n576 B.n575 10.6151
R1284 B.n577 B.n576 10.6151
R1285 B.n577 B.n345 10.6151
R1286 B.n583 B.n345 10.6151
R1287 B.n584 B.n583 10.6151
R1288 B.n585 B.n584 10.6151
R1289 B.n585 B.n343 10.6151
R1290 B.n591 B.n343 10.6151
R1291 B.n592 B.n591 10.6151
R1292 B.n598 B.n597 10.6151
R1293 B.n599 B.n598 10.6151
R1294 B.n599 B.n331 10.6151
R1295 B.n610 B.n331 10.6151
R1296 B.n611 B.n610 10.6151
R1297 B.n612 B.n611 10.6151
R1298 B.n612 B.n324 10.6151
R1299 B.n622 B.n324 10.6151
R1300 B.n623 B.n622 10.6151
R1301 B.n624 B.n623 10.6151
R1302 B.n624 B.n316 10.6151
R1303 B.n634 B.n316 10.6151
R1304 B.n635 B.n634 10.6151
R1305 B.n636 B.n635 10.6151
R1306 B.n636 B.n308 10.6151
R1307 B.n647 B.n308 10.6151
R1308 B.n648 B.n647 10.6151
R1309 B.n649 B.n648 10.6151
R1310 B.n649 B.n301 10.6151
R1311 B.n660 B.n301 10.6151
R1312 B.n661 B.n660 10.6151
R1313 B.n662 B.n661 10.6151
R1314 B.n662 B.n0 10.6151
R1315 B.n746 B.n1 10.6151
R1316 B.n746 B.n745 10.6151
R1317 B.n745 B.n744 10.6151
R1318 B.n744 B.n10 10.6151
R1319 B.n738 B.n10 10.6151
R1320 B.n738 B.n737 10.6151
R1321 B.n737 B.n736 10.6151
R1322 B.n736 B.n16 10.6151
R1323 B.n730 B.n16 10.6151
R1324 B.n730 B.n729 10.6151
R1325 B.n729 B.n728 10.6151
R1326 B.n728 B.n24 10.6151
R1327 B.n722 B.n24 10.6151
R1328 B.n722 B.n721 10.6151
R1329 B.n721 B.n720 10.6151
R1330 B.n720 B.n31 10.6151
R1331 B.n714 B.n31 10.6151
R1332 B.n714 B.n713 10.6151
R1333 B.n713 B.n712 10.6151
R1334 B.n712 B.n37 10.6151
R1335 B.n706 B.n37 10.6151
R1336 B.n706 B.n705 10.6151
R1337 B.n705 B.n704 10.6151
R1338 B.t1 B.n299 7.19592
R1339 B.t2 B.n8 7.19592
R1340 B.n192 B.n191 6.5566
R1341 B.n208 B.n100 6.5566
R1342 B.n486 B.n373 6.5566
R1343 B.n503 B.n502 6.5566
R1344 B.n191 B.n190 4.05904
R1345 B.n211 B.n100 4.05904
R1346 B.n374 B.n373 4.05904
R1347 B.n504 B.n503 4.05904
R1348 B.n752 B.n0 2.81026
R1349 B.n752 B.n1 2.81026
R1350 B.n607 B.t9 1.19974
R1351 B.n39 B.t16 1.19974
R1352 VP.n6 VP.t4 502.736
R1353 VP.n14 VP.t0 479.07
R1354 VP.n16 VP.t7 479.07
R1355 VP.n20 VP.t6 479.07
R1356 VP.n22 VP.t2 479.07
R1357 VP.n11 VP.t1 479.07
R1358 VP.n9 VP.t3 479.07
R1359 VP.n5 VP.t5 479.07
R1360 VP.n23 VP.n22 161.3
R1361 VP.n8 VP.n7 161.3
R1362 VP.n9 VP.n4 161.3
R1363 VP.n10 VP.n3 161.3
R1364 VP.n12 VP.n11 161.3
R1365 VP.n21 VP.n0 161.3
R1366 VP.n20 VP.n19 161.3
R1367 VP.n18 VP.n1 161.3
R1368 VP.n17 VP.n16 161.3
R1369 VP.n15 VP.n2 161.3
R1370 VP.n14 VP.n13 161.3
R1371 VP.n7 VP.n6 44.9044
R1372 VP.n13 VP.n12 43.046
R1373 VP.n15 VP.n14 34.3247
R1374 VP.n22 VP.n21 34.3247
R1375 VP.n11 VP.n10 34.3247
R1376 VP.n16 VP.n1 24.1005
R1377 VP.n20 VP.n1 24.1005
R1378 VP.n8 VP.n5 24.1005
R1379 VP.n9 VP.n8 24.1005
R1380 VP.n6 VP.n5 17.9645
R1381 VP.n16 VP.n15 13.8763
R1382 VP.n21 VP.n20 13.8763
R1383 VP.n10 VP.n9 13.8763
R1384 VP.n7 VP.n4 0.189894
R1385 VP.n4 VP.n3 0.189894
R1386 VP.n12 VP.n3 0.189894
R1387 VP.n13 VP.n2 0.189894
R1388 VP.n17 VP.n2 0.189894
R1389 VP.n18 VP.n17 0.189894
R1390 VP.n19 VP.n18 0.189894
R1391 VP.n19 VP.n0 0.189894
R1392 VP.n23 VP.n0 0.189894
R1393 VP VP.n23 0.0516364
R1394 VDD1 VDD1.n0 66.157
R1395 VDD1.n3 VDD1.n2 66.0422
R1396 VDD1.n3 VDD1.n1 66.0422
R1397 VDD1.n5 VDD1.n4 65.6364
R1398 VDD1.n5 VDD1.n3 39.7164
R1399 VDD1.n4 VDD1.t4 1.51542
R1400 VDD1.n4 VDD1.t6 1.51542
R1401 VDD1.n0 VDD1.t3 1.51542
R1402 VDD1.n0 VDD1.t2 1.51542
R1403 VDD1.n2 VDD1.t1 1.51542
R1404 VDD1.n2 VDD1.t5 1.51542
R1405 VDD1.n1 VDD1.t7 1.51542
R1406 VDD1.n1 VDD1.t0 1.51542
R1407 VDD1 VDD1.n5 0.403517
C0 VP VDD2 0.321437f
C1 VP VTAIL 5.88698f
C2 VP VDD1 6.31475f
C3 VN VDD2 6.14183f
C4 VTAIL VN 5.87288f
C5 VN VDD1 0.148056f
C6 VTAIL VDD2 11.6248f
C7 VP VN 5.58449f
C8 VDD1 VDD2 0.843884f
C9 VTAIL VDD1 11.5828f
C10 VDD2 B 3.600393f
C11 VDD1 B 3.840803f
C12 VTAIL B 9.586477f
C13 VN B 8.842549f
C14 VP B 6.861428f
C15 VDD1.t3 B 0.280692f
C16 VDD1.t2 B 0.280692f
C17 VDD1.n0 B 2.52754f
C18 VDD1.t7 B 0.280692f
C19 VDD1.t0 B 0.280692f
C20 VDD1.n1 B 2.52688f
C21 VDD1.t1 B 0.280692f
C22 VDD1.t5 B 0.280692f
C23 VDD1.n2 B 2.52688f
C24 VDD1.n3 B 2.49923f
C25 VDD1.t4 B 0.280692f
C26 VDD1.t6 B 0.280692f
C27 VDD1.n4 B 2.52477f
C28 VDD1.n5 B 2.61875f
C29 VP.n0 B 0.043679f
C30 VP.n1 B 0.009912f
C31 VP.n2 B 0.043679f
C32 VP.n3 B 0.043679f
C33 VP.t1 B 1.20324f
C34 VP.t3 B 1.20324f
C35 VP.n4 B 0.043679f
C36 VP.t5 B 1.20324f
C37 VP.n5 B 0.477344f
C38 VP.t4 B 1.22552f
C39 VP.n6 B 0.45477f
C40 VP.n7 B 0.18591f
C41 VP.n8 B 0.009912f
C42 VP.n9 B 0.472113f
C43 VP.n10 B 0.009912f
C44 VP.n11 B 0.47144f
C45 VP.n12 B 1.87776f
C46 VP.n13 B 1.91423f
C47 VP.t0 B 1.20324f
C48 VP.n14 B 0.47144f
C49 VP.n15 B 0.009912f
C50 VP.t7 B 1.20324f
C51 VP.n16 B 0.472113f
C52 VP.n17 B 0.043679f
C53 VP.n18 B 0.043679f
C54 VP.n19 B 0.043679f
C55 VP.t6 B 1.20324f
C56 VP.n20 B 0.472113f
C57 VP.n21 B 0.009912f
C58 VP.t2 B 1.20324f
C59 VP.n22 B 0.47144f
C60 VP.n23 B 0.03385f
C61 VTAIL.t8 B 0.20463f
C62 VTAIL.t15 B 0.20463f
C63 VTAIL.n0 B 1.78844f
C64 VTAIL.n1 B 0.244735f
C65 VTAIL.t12 B 2.28223f
C66 VTAIL.n2 B 0.335305f
C67 VTAIL.t1 B 2.28223f
C68 VTAIL.n3 B 0.335305f
C69 VTAIL.t0 B 0.20463f
C70 VTAIL.t7 B 0.20463f
C71 VTAIL.n4 B 1.78844f
C72 VTAIL.n5 B 0.299908f
C73 VTAIL.t6 B 2.28223f
C74 VTAIL.n6 B 1.35263f
C75 VTAIL.t14 B 2.28224f
C76 VTAIL.n7 B 1.35262f
C77 VTAIL.t11 B 0.20463f
C78 VTAIL.t10 B 0.20463f
C79 VTAIL.n8 B 1.78845f
C80 VTAIL.n9 B 0.299899f
C81 VTAIL.t9 B 2.28224f
C82 VTAIL.n10 B 0.335292f
C83 VTAIL.t2 B 2.28224f
C84 VTAIL.n11 B 0.335292f
C85 VTAIL.t3 B 0.20463f
C86 VTAIL.t4 B 0.20463f
C87 VTAIL.n12 B 1.78845f
C88 VTAIL.n13 B 0.299899f
C89 VTAIL.t5 B 2.28223f
C90 VTAIL.n14 B 1.35263f
C91 VTAIL.t13 B 2.28223f
C92 VTAIL.n15 B 1.34892f
C93 VDD2.t3 B 0.279121f
C94 VDD2.t6 B 0.279121f
C95 VDD2.n0 B 2.51274f
C96 VDD2.t0 B 0.279121f
C97 VDD2.t4 B 0.279121f
C98 VDD2.n1 B 2.51274f
C99 VDD2.n2 B 2.42767f
C100 VDD2.t1 B 0.279121f
C101 VDD2.t2 B 0.279121f
C102 VDD2.n3 B 2.51064f
C103 VDD2.n4 B 2.57197f
C104 VDD2.t5 B 0.279121f
C105 VDD2.t7 B 0.279121f
C106 VDD2.n5 B 2.51271f
C107 VN.n0 B 0.04304f
C108 VN.n1 B 0.009767f
C109 VN.t3 B 1.20758f
C110 VN.t7 B 1.18563f
C111 VN.n2 B 0.470358f
C112 VN.n3 B 0.448114f
C113 VN.n4 B 0.183189f
C114 VN.n5 B 0.04304f
C115 VN.t0 B 1.18563f
C116 VN.n6 B 0.465204f
C117 VN.n7 B 0.009767f
C118 VN.t2 B 1.18563f
C119 VN.n8 B 0.46454f
C120 VN.n9 B 0.033354f
C121 VN.n10 B 0.04304f
C122 VN.n11 B 0.009767f
C123 VN.t4 B 1.18563f
C124 VN.t6 B 1.20758f
C125 VN.t5 B 1.18563f
C126 VN.n12 B 0.470358f
C127 VN.n13 B 0.448114f
C128 VN.n14 B 0.183189f
C129 VN.n15 B 0.04304f
C130 VN.n16 B 0.465204f
C131 VN.n17 B 0.009767f
C132 VN.t1 B 1.18563f
C133 VN.n18 B 0.46454f
C134 VN.n19 B 1.87849f
.ends

