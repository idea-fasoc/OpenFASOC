* NGSPICE file created from diff_pair_sample_1508.ext - technology: sky130A

.subckt diff_pair_sample_1508 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=0.91
X1 VDD1.t3 VP.t0 VTAIL.t1 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=0.91
X2 VDD2.t0 VN.t1 VTAIL.t6 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=0.91
X3 B.t11 B.t9 B.t10 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=0.91
X4 B.t8 B.t6 B.t7 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=0.91
X5 VTAIL.t3 VP.t1 VDD1.t2 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=0.91
X6 VTAIL.t5 VN.t2 VDD2.t3 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=0.91
X7 VDD1.t1 VP.t2 VTAIL.t2 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=0.91
X8 B.t5 B.t3 B.t4 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=0.91
X9 VDD2.t1 VN.t3 VTAIL.t4 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=0.91
X10 VTAIL.t0 VP.t3 VDD1.t0 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=0.91
X11 B.t2 B.t0 B.t1 w_n1714_n4616# sky130_fd_pr__pfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=0.91
R0 VN.n0 VN.t2 544.835
R1 VN.n1 VN.t1 544.835
R2 VN.n1 VN.t0 544.747
R3 VN.n0 VN.t3 544.747
R4 VN VN.n1 77.3342
R5 VN VN.n0 31.2622
R6 VDD2.n2 VDD2.n0 111.334
R7 VDD2.n2 VDD2.n1 68.6877
R8 VDD2.n1 VDD2.t2 1.78257
R9 VDD2.n1 VDD2.t0 1.78257
R10 VDD2.n0 VDD2.t3 1.78257
R11 VDD2.n0 VDD2.t1 1.78257
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n810 VTAIL.n714 756.745
R14 VTAIL.n96 VTAIL.n0 756.745
R15 VTAIL.n198 VTAIL.n102 756.745
R16 VTAIL.n300 VTAIL.n204 756.745
R17 VTAIL.n708 VTAIL.n612 756.745
R18 VTAIL.n606 VTAIL.n510 756.745
R19 VTAIL.n504 VTAIL.n408 756.745
R20 VTAIL.n402 VTAIL.n306 756.745
R21 VTAIL.n746 VTAIL.n745 585
R22 VTAIL.n751 VTAIL.n750 585
R23 VTAIL.n753 VTAIL.n752 585
R24 VTAIL.n742 VTAIL.n741 585
R25 VTAIL.n759 VTAIL.n758 585
R26 VTAIL.n761 VTAIL.n760 585
R27 VTAIL.n738 VTAIL.n737 585
R28 VTAIL.n767 VTAIL.n766 585
R29 VTAIL.n769 VTAIL.n768 585
R30 VTAIL.n734 VTAIL.n733 585
R31 VTAIL.n775 VTAIL.n774 585
R32 VTAIL.n777 VTAIL.n776 585
R33 VTAIL.n730 VTAIL.n729 585
R34 VTAIL.n783 VTAIL.n782 585
R35 VTAIL.n785 VTAIL.n784 585
R36 VTAIL.n726 VTAIL.n725 585
R37 VTAIL.n792 VTAIL.n791 585
R38 VTAIL.n793 VTAIL.n724 585
R39 VTAIL.n795 VTAIL.n794 585
R40 VTAIL.n722 VTAIL.n721 585
R41 VTAIL.n801 VTAIL.n800 585
R42 VTAIL.n803 VTAIL.n802 585
R43 VTAIL.n718 VTAIL.n717 585
R44 VTAIL.n809 VTAIL.n808 585
R45 VTAIL.n811 VTAIL.n810 585
R46 VTAIL.n32 VTAIL.n31 585
R47 VTAIL.n37 VTAIL.n36 585
R48 VTAIL.n39 VTAIL.n38 585
R49 VTAIL.n28 VTAIL.n27 585
R50 VTAIL.n45 VTAIL.n44 585
R51 VTAIL.n47 VTAIL.n46 585
R52 VTAIL.n24 VTAIL.n23 585
R53 VTAIL.n53 VTAIL.n52 585
R54 VTAIL.n55 VTAIL.n54 585
R55 VTAIL.n20 VTAIL.n19 585
R56 VTAIL.n61 VTAIL.n60 585
R57 VTAIL.n63 VTAIL.n62 585
R58 VTAIL.n16 VTAIL.n15 585
R59 VTAIL.n69 VTAIL.n68 585
R60 VTAIL.n71 VTAIL.n70 585
R61 VTAIL.n12 VTAIL.n11 585
R62 VTAIL.n78 VTAIL.n77 585
R63 VTAIL.n79 VTAIL.n10 585
R64 VTAIL.n81 VTAIL.n80 585
R65 VTAIL.n8 VTAIL.n7 585
R66 VTAIL.n87 VTAIL.n86 585
R67 VTAIL.n89 VTAIL.n88 585
R68 VTAIL.n4 VTAIL.n3 585
R69 VTAIL.n95 VTAIL.n94 585
R70 VTAIL.n97 VTAIL.n96 585
R71 VTAIL.n134 VTAIL.n133 585
R72 VTAIL.n139 VTAIL.n138 585
R73 VTAIL.n141 VTAIL.n140 585
R74 VTAIL.n130 VTAIL.n129 585
R75 VTAIL.n147 VTAIL.n146 585
R76 VTAIL.n149 VTAIL.n148 585
R77 VTAIL.n126 VTAIL.n125 585
R78 VTAIL.n155 VTAIL.n154 585
R79 VTAIL.n157 VTAIL.n156 585
R80 VTAIL.n122 VTAIL.n121 585
R81 VTAIL.n163 VTAIL.n162 585
R82 VTAIL.n165 VTAIL.n164 585
R83 VTAIL.n118 VTAIL.n117 585
R84 VTAIL.n171 VTAIL.n170 585
R85 VTAIL.n173 VTAIL.n172 585
R86 VTAIL.n114 VTAIL.n113 585
R87 VTAIL.n180 VTAIL.n179 585
R88 VTAIL.n181 VTAIL.n112 585
R89 VTAIL.n183 VTAIL.n182 585
R90 VTAIL.n110 VTAIL.n109 585
R91 VTAIL.n189 VTAIL.n188 585
R92 VTAIL.n191 VTAIL.n190 585
R93 VTAIL.n106 VTAIL.n105 585
R94 VTAIL.n197 VTAIL.n196 585
R95 VTAIL.n199 VTAIL.n198 585
R96 VTAIL.n236 VTAIL.n235 585
R97 VTAIL.n241 VTAIL.n240 585
R98 VTAIL.n243 VTAIL.n242 585
R99 VTAIL.n232 VTAIL.n231 585
R100 VTAIL.n249 VTAIL.n248 585
R101 VTAIL.n251 VTAIL.n250 585
R102 VTAIL.n228 VTAIL.n227 585
R103 VTAIL.n257 VTAIL.n256 585
R104 VTAIL.n259 VTAIL.n258 585
R105 VTAIL.n224 VTAIL.n223 585
R106 VTAIL.n265 VTAIL.n264 585
R107 VTAIL.n267 VTAIL.n266 585
R108 VTAIL.n220 VTAIL.n219 585
R109 VTAIL.n273 VTAIL.n272 585
R110 VTAIL.n275 VTAIL.n274 585
R111 VTAIL.n216 VTAIL.n215 585
R112 VTAIL.n282 VTAIL.n281 585
R113 VTAIL.n283 VTAIL.n214 585
R114 VTAIL.n285 VTAIL.n284 585
R115 VTAIL.n212 VTAIL.n211 585
R116 VTAIL.n291 VTAIL.n290 585
R117 VTAIL.n293 VTAIL.n292 585
R118 VTAIL.n208 VTAIL.n207 585
R119 VTAIL.n299 VTAIL.n298 585
R120 VTAIL.n301 VTAIL.n300 585
R121 VTAIL.n709 VTAIL.n708 585
R122 VTAIL.n707 VTAIL.n706 585
R123 VTAIL.n616 VTAIL.n615 585
R124 VTAIL.n701 VTAIL.n700 585
R125 VTAIL.n699 VTAIL.n698 585
R126 VTAIL.n620 VTAIL.n619 585
R127 VTAIL.n693 VTAIL.n692 585
R128 VTAIL.n691 VTAIL.n622 585
R129 VTAIL.n690 VTAIL.n689 585
R130 VTAIL.n625 VTAIL.n623 585
R131 VTAIL.n684 VTAIL.n683 585
R132 VTAIL.n682 VTAIL.n681 585
R133 VTAIL.n629 VTAIL.n628 585
R134 VTAIL.n676 VTAIL.n675 585
R135 VTAIL.n674 VTAIL.n673 585
R136 VTAIL.n633 VTAIL.n632 585
R137 VTAIL.n668 VTAIL.n667 585
R138 VTAIL.n666 VTAIL.n665 585
R139 VTAIL.n637 VTAIL.n636 585
R140 VTAIL.n660 VTAIL.n659 585
R141 VTAIL.n658 VTAIL.n657 585
R142 VTAIL.n641 VTAIL.n640 585
R143 VTAIL.n652 VTAIL.n651 585
R144 VTAIL.n650 VTAIL.n649 585
R145 VTAIL.n645 VTAIL.n644 585
R146 VTAIL.n607 VTAIL.n606 585
R147 VTAIL.n605 VTAIL.n604 585
R148 VTAIL.n514 VTAIL.n513 585
R149 VTAIL.n599 VTAIL.n598 585
R150 VTAIL.n597 VTAIL.n596 585
R151 VTAIL.n518 VTAIL.n517 585
R152 VTAIL.n591 VTAIL.n590 585
R153 VTAIL.n589 VTAIL.n520 585
R154 VTAIL.n588 VTAIL.n587 585
R155 VTAIL.n523 VTAIL.n521 585
R156 VTAIL.n582 VTAIL.n581 585
R157 VTAIL.n580 VTAIL.n579 585
R158 VTAIL.n527 VTAIL.n526 585
R159 VTAIL.n574 VTAIL.n573 585
R160 VTAIL.n572 VTAIL.n571 585
R161 VTAIL.n531 VTAIL.n530 585
R162 VTAIL.n566 VTAIL.n565 585
R163 VTAIL.n564 VTAIL.n563 585
R164 VTAIL.n535 VTAIL.n534 585
R165 VTAIL.n558 VTAIL.n557 585
R166 VTAIL.n556 VTAIL.n555 585
R167 VTAIL.n539 VTAIL.n538 585
R168 VTAIL.n550 VTAIL.n549 585
R169 VTAIL.n548 VTAIL.n547 585
R170 VTAIL.n543 VTAIL.n542 585
R171 VTAIL.n505 VTAIL.n504 585
R172 VTAIL.n503 VTAIL.n502 585
R173 VTAIL.n412 VTAIL.n411 585
R174 VTAIL.n497 VTAIL.n496 585
R175 VTAIL.n495 VTAIL.n494 585
R176 VTAIL.n416 VTAIL.n415 585
R177 VTAIL.n489 VTAIL.n488 585
R178 VTAIL.n487 VTAIL.n418 585
R179 VTAIL.n486 VTAIL.n485 585
R180 VTAIL.n421 VTAIL.n419 585
R181 VTAIL.n480 VTAIL.n479 585
R182 VTAIL.n478 VTAIL.n477 585
R183 VTAIL.n425 VTAIL.n424 585
R184 VTAIL.n472 VTAIL.n471 585
R185 VTAIL.n470 VTAIL.n469 585
R186 VTAIL.n429 VTAIL.n428 585
R187 VTAIL.n464 VTAIL.n463 585
R188 VTAIL.n462 VTAIL.n461 585
R189 VTAIL.n433 VTAIL.n432 585
R190 VTAIL.n456 VTAIL.n455 585
R191 VTAIL.n454 VTAIL.n453 585
R192 VTAIL.n437 VTAIL.n436 585
R193 VTAIL.n448 VTAIL.n447 585
R194 VTAIL.n446 VTAIL.n445 585
R195 VTAIL.n441 VTAIL.n440 585
R196 VTAIL.n403 VTAIL.n402 585
R197 VTAIL.n401 VTAIL.n400 585
R198 VTAIL.n310 VTAIL.n309 585
R199 VTAIL.n395 VTAIL.n394 585
R200 VTAIL.n393 VTAIL.n392 585
R201 VTAIL.n314 VTAIL.n313 585
R202 VTAIL.n387 VTAIL.n386 585
R203 VTAIL.n385 VTAIL.n316 585
R204 VTAIL.n384 VTAIL.n383 585
R205 VTAIL.n319 VTAIL.n317 585
R206 VTAIL.n378 VTAIL.n377 585
R207 VTAIL.n376 VTAIL.n375 585
R208 VTAIL.n323 VTAIL.n322 585
R209 VTAIL.n370 VTAIL.n369 585
R210 VTAIL.n368 VTAIL.n367 585
R211 VTAIL.n327 VTAIL.n326 585
R212 VTAIL.n362 VTAIL.n361 585
R213 VTAIL.n360 VTAIL.n359 585
R214 VTAIL.n331 VTAIL.n330 585
R215 VTAIL.n354 VTAIL.n353 585
R216 VTAIL.n352 VTAIL.n351 585
R217 VTAIL.n335 VTAIL.n334 585
R218 VTAIL.n346 VTAIL.n345 585
R219 VTAIL.n344 VTAIL.n343 585
R220 VTAIL.n339 VTAIL.n338 585
R221 VTAIL.n747 VTAIL.t4 327.466
R222 VTAIL.n33 VTAIL.t5 327.466
R223 VTAIL.n135 VTAIL.t2 327.466
R224 VTAIL.n237 VTAIL.t0 327.466
R225 VTAIL.n646 VTAIL.t1 327.466
R226 VTAIL.n544 VTAIL.t3 327.466
R227 VTAIL.n442 VTAIL.t6 327.466
R228 VTAIL.n340 VTAIL.t7 327.466
R229 VTAIL.n751 VTAIL.n745 171.744
R230 VTAIL.n752 VTAIL.n751 171.744
R231 VTAIL.n752 VTAIL.n741 171.744
R232 VTAIL.n759 VTAIL.n741 171.744
R233 VTAIL.n760 VTAIL.n759 171.744
R234 VTAIL.n760 VTAIL.n737 171.744
R235 VTAIL.n767 VTAIL.n737 171.744
R236 VTAIL.n768 VTAIL.n767 171.744
R237 VTAIL.n768 VTAIL.n733 171.744
R238 VTAIL.n775 VTAIL.n733 171.744
R239 VTAIL.n776 VTAIL.n775 171.744
R240 VTAIL.n776 VTAIL.n729 171.744
R241 VTAIL.n783 VTAIL.n729 171.744
R242 VTAIL.n784 VTAIL.n783 171.744
R243 VTAIL.n784 VTAIL.n725 171.744
R244 VTAIL.n792 VTAIL.n725 171.744
R245 VTAIL.n793 VTAIL.n792 171.744
R246 VTAIL.n794 VTAIL.n793 171.744
R247 VTAIL.n794 VTAIL.n721 171.744
R248 VTAIL.n801 VTAIL.n721 171.744
R249 VTAIL.n802 VTAIL.n801 171.744
R250 VTAIL.n802 VTAIL.n717 171.744
R251 VTAIL.n809 VTAIL.n717 171.744
R252 VTAIL.n810 VTAIL.n809 171.744
R253 VTAIL.n37 VTAIL.n31 171.744
R254 VTAIL.n38 VTAIL.n37 171.744
R255 VTAIL.n38 VTAIL.n27 171.744
R256 VTAIL.n45 VTAIL.n27 171.744
R257 VTAIL.n46 VTAIL.n45 171.744
R258 VTAIL.n46 VTAIL.n23 171.744
R259 VTAIL.n53 VTAIL.n23 171.744
R260 VTAIL.n54 VTAIL.n53 171.744
R261 VTAIL.n54 VTAIL.n19 171.744
R262 VTAIL.n61 VTAIL.n19 171.744
R263 VTAIL.n62 VTAIL.n61 171.744
R264 VTAIL.n62 VTAIL.n15 171.744
R265 VTAIL.n69 VTAIL.n15 171.744
R266 VTAIL.n70 VTAIL.n69 171.744
R267 VTAIL.n70 VTAIL.n11 171.744
R268 VTAIL.n78 VTAIL.n11 171.744
R269 VTAIL.n79 VTAIL.n78 171.744
R270 VTAIL.n80 VTAIL.n79 171.744
R271 VTAIL.n80 VTAIL.n7 171.744
R272 VTAIL.n87 VTAIL.n7 171.744
R273 VTAIL.n88 VTAIL.n87 171.744
R274 VTAIL.n88 VTAIL.n3 171.744
R275 VTAIL.n95 VTAIL.n3 171.744
R276 VTAIL.n96 VTAIL.n95 171.744
R277 VTAIL.n139 VTAIL.n133 171.744
R278 VTAIL.n140 VTAIL.n139 171.744
R279 VTAIL.n140 VTAIL.n129 171.744
R280 VTAIL.n147 VTAIL.n129 171.744
R281 VTAIL.n148 VTAIL.n147 171.744
R282 VTAIL.n148 VTAIL.n125 171.744
R283 VTAIL.n155 VTAIL.n125 171.744
R284 VTAIL.n156 VTAIL.n155 171.744
R285 VTAIL.n156 VTAIL.n121 171.744
R286 VTAIL.n163 VTAIL.n121 171.744
R287 VTAIL.n164 VTAIL.n163 171.744
R288 VTAIL.n164 VTAIL.n117 171.744
R289 VTAIL.n171 VTAIL.n117 171.744
R290 VTAIL.n172 VTAIL.n171 171.744
R291 VTAIL.n172 VTAIL.n113 171.744
R292 VTAIL.n180 VTAIL.n113 171.744
R293 VTAIL.n181 VTAIL.n180 171.744
R294 VTAIL.n182 VTAIL.n181 171.744
R295 VTAIL.n182 VTAIL.n109 171.744
R296 VTAIL.n189 VTAIL.n109 171.744
R297 VTAIL.n190 VTAIL.n189 171.744
R298 VTAIL.n190 VTAIL.n105 171.744
R299 VTAIL.n197 VTAIL.n105 171.744
R300 VTAIL.n198 VTAIL.n197 171.744
R301 VTAIL.n241 VTAIL.n235 171.744
R302 VTAIL.n242 VTAIL.n241 171.744
R303 VTAIL.n242 VTAIL.n231 171.744
R304 VTAIL.n249 VTAIL.n231 171.744
R305 VTAIL.n250 VTAIL.n249 171.744
R306 VTAIL.n250 VTAIL.n227 171.744
R307 VTAIL.n257 VTAIL.n227 171.744
R308 VTAIL.n258 VTAIL.n257 171.744
R309 VTAIL.n258 VTAIL.n223 171.744
R310 VTAIL.n265 VTAIL.n223 171.744
R311 VTAIL.n266 VTAIL.n265 171.744
R312 VTAIL.n266 VTAIL.n219 171.744
R313 VTAIL.n273 VTAIL.n219 171.744
R314 VTAIL.n274 VTAIL.n273 171.744
R315 VTAIL.n274 VTAIL.n215 171.744
R316 VTAIL.n282 VTAIL.n215 171.744
R317 VTAIL.n283 VTAIL.n282 171.744
R318 VTAIL.n284 VTAIL.n283 171.744
R319 VTAIL.n284 VTAIL.n211 171.744
R320 VTAIL.n291 VTAIL.n211 171.744
R321 VTAIL.n292 VTAIL.n291 171.744
R322 VTAIL.n292 VTAIL.n207 171.744
R323 VTAIL.n299 VTAIL.n207 171.744
R324 VTAIL.n300 VTAIL.n299 171.744
R325 VTAIL.n708 VTAIL.n707 171.744
R326 VTAIL.n707 VTAIL.n615 171.744
R327 VTAIL.n700 VTAIL.n615 171.744
R328 VTAIL.n700 VTAIL.n699 171.744
R329 VTAIL.n699 VTAIL.n619 171.744
R330 VTAIL.n692 VTAIL.n619 171.744
R331 VTAIL.n692 VTAIL.n691 171.744
R332 VTAIL.n691 VTAIL.n690 171.744
R333 VTAIL.n690 VTAIL.n623 171.744
R334 VTAIL.n683 VTAIL.n623 171.744
R335 VTAIL.n683 VTAIL.n682 171.744
R336 VTAIL.n682 VTAIL.n628 171.744
R337 VTAIL.n675 VTAIL.n628 171.744
R338 VTAIL.n675 VTAIL.n674 171.744
R339 VTAIL.n674 VTAIL.n632 171.744
R340 VTAIL.n667 VTAIL.n632 171.744
R341 VTAIL.n667 VTAIL.n666 171.744
R342 VTAIL.n666 VTAIL.n636 171.744
R343 VTAIL.n659 VTAIL.n636 171.744
R344 VTAIL.n659 VTAIL.n658 171.744
R345 VTAIL.n658 VTAIL.n640 171.744
R346 VTAIL.n651 VTAIL.n640 171.744
R347 VTAIL.n651 VTAIL.n650 171.744
R348 VTAIL.n650 VTAIL.n644 171.744
R349 VTAIL.n606 VTAIL.n605 171.744
R350 VTAIL.n605 VTAIL.n513 171.744
R351 VTAIL.n598 VTAIL.n513 171.744
R352 VTAIL.n598 VTAIL.n597 171.744
R353 VTAIL.n597 VTAIL.n517 171.744
R354 VTAIL.n590 VTAIL.n517 171.744
R355 VTAIL.n590 VTAIL.n589 171.744
R356 VTAIL.n589 VTAIL.n588 171.744
R357 VTAIL.n588 VTAIL.n521 171.744
R358 VTAIL.n581 VTAIL.n521 171.744
R359 VTAIL.n581 VTAIL.n580 171.744
R360 VTAIL.n580 VTAIL.n526 171.744
R361 VTAIL.n573 VTAIL.n526 171.744
R362 VTAIL.n573 VTAIL.n572 171.744
R363 VTAIL.n572 VTAIL.n530 171.744
R364 VTAIL.n565 VTAIL.n530 171.744
R365 VTAIL.n565 VTAIL.n564 171.744
R366 VTAIL.n564 VTAIL.n534 171.744
R367 VTAIL.n557 VTAIL.n534 171.744
R368 VTAIL.n557 VTAIL.n556 171.744
R369 VTAIL.n556 VTAIL.n538 171.744
R370 VTAIL.n549 VTAIL.n538 171.744
R371 VTAIL.n549 VTAIL.n548 171.744
R372 VTAIL.n548 VTAIL.n542 171.744
R373 VTAIL.n504 VTAIL.n503 171.744
R374 VTAIL.n503 VTAIL.n411 171.744
R375 VTAIL.n496 VTAIL.n411 171.744
R376 VTAIL.n496 VTAIL.n495 171.744
R377 VTAIL.n495 VTAIL.n415 171.744
R378 VTAIL.n488 VTAIL.n415 171.744
R379 VTAIL.n488 VTAIL.n487 171.744
R380 VTAIL.n487 VTAIL.n486 171.744
R381 VTAIL.n486 VTAIL.n419 171.744
R382 VTAIL.n479 VTAIL.n419 171.744
R383 VTAIL.n479 VTAIL.n478 171.744
R384 VTAIL.n478 VTAIL.n424 171.744
R385 VTAIL.n471 VTAIL.n424 171.744
R386 VTAIL.n471 VTAIL.n470 171.744
R387 VTAIL.n470 VTAIL.n428 171.744
R388 VTAIL.n463 VTAIL.n428 171.744
R389 VTAIL.n463 VTAIL.n462 171.744
R390 VTAIL.n462 VTAIL.n432 171.744
R391 VTAIL.n455 VTAIL.n432 171.744
R392 VTAIL.n455 VTAIL.n454 171.744
R393 VTAIL.n454 VTAIL.n436 171.744
R394 VTAIL.n447 VTAIL.n436 171.744
R395 VTAIL.n447 VTAIL.n446 171.744
R396 VTAIL.n446 VTAIL.n440 171.744
R397 VTAIL.n402 VTAIL.n401 171.744
R398 VTAIL.n401 VTAIL.n309 171.744
R399 VTAIL.n394 VTAIL.n309 171.744
R400 VTAIL.n394 VTAIL.n393 171.744
R401 VTAIL.n393 VTAIL.n313 171.744
R402 VTAIL.n386 VTAIL.n313 171.744
R403 VTAIL.n386 VTAIL.n385 171.744
R404 VTAIL.n385 VTAIL.n384 171.744
R405 VTAIL.n384 VTAIL.n317 171.744
R406 VTAIL.n377 VTAIL.n317 171.744
R407 VTAIL.n377 VTAIL.n376 171.744
R408 VTAIL.n376 VTAIL.n322 171.744
R409 VTAIL.n369 VTAIL.n322 171.744
R410 VTAIL.n369 VTAIL.n368 171.744
R411 VTAIL.n368 VTAIL.n326 171.744
R412 VTAIL.n361 VTAIL.n326 171.744
R413 VTAIL.n361 VTAIL.n360 171.744
R414 VTAIL.n360 VTAIL.n330 171.744
R415 VTAIL.n353 VTAIL.n330 171.744
R416 VTAIL.n353 VTAIL.n352 171.744
R417 VTAIL.n352 VTAIL.n334 171.744
R418 VTAIL.n345 VTAIL.n334 171.744
R419 VTAIL.n345 VTAIL.n344 171.744
R420 VTAIL.n344 VTAIL.n338 171.744
R421 VTAIL.t4 VTAIL.n745 85.8723
R422 VTAIL.t5 VTAIL.n31 85.8723
R423 VTAIL.t2 VTAIL.n133 85.8723
R424 VTAIL.t0 VTAIL.n235 85.8723
R425 VTAIL.t1 VTAIL.n644 85.8723
R426 VTAIL.t3 VTAIL.n542 85.8723
R427 VTAIL.t6 VTAIL.n440 85.8723
R428 VTAIL.t7 VTAIL.n338 85.8723
R429 VTAIL.n815 VTAIL.n814 32.1853
R430 VTAIL.n101 VTAIL.n100 32.1853
R431 VTAIL.n203 VTAIL.n202 32.1853
R432 VTAIL.n305 VTAIL.n304 32.1853
R433 VTAIL.n713 VTAIL.n712 32.1853
R434 VTAIL.n611 VTAIL.n610 32.1853
R435 VTAIL.n509 VTAIL.n508 32.1853
R436 VTAIL.n407 VTAIL.n406 32.1853
R437 VTAIL.n815 VTAIL.n713 29.16
R438 VTAIL.n407 VTAIL.n305 29.16
R439 VTAIL.n747 VTAIL.n746 16.3895
R440 VTAIL.n33 VTAIL.n32 16.3895
R441 VTAIL.n135 VTAIL.n134 16.3895
R442 VTAIL.n237 VTAIL.n236 16.3895
R443 VTAIL.n646 VTAIL.n645 16.3895
R444 VTAIL.n544 VTAIL.n543 16.3895
R445 VTAIL.n442 VTAIL.n441 16.3895
R446 VTAIL.n340 VTAIL.n339 16.3895
R447 VTAIL.n795 VTAIL.n724 13.1884
R448 VTAIL.n81 VTAIL.n10 13.1884
R449 VTAIL.n183 VTAIL.n112 13.1884
R450 VTAIL.n285 VTAIL.n214 13.1884
R451 VTAIL.n693 VTAIL.n622 13.1884
R452 VTAIL.n591 VTAIL.n520 13.1884
R453 VTAIL.n489 VTAIL.n418 13.1884
R454 VTAIL.n387 VTAIL.n316 13.1884
R455 VTAIL.n750 VTAIL.n749 12.8005
R456 VTAIL.n791 VTAIL.n790 12.8005
R457 VTAIL.n796 VTAIL.n722 12.8005
R458 VTAIL.n36 VTAIL.n35 12.8005
R459 VTAIL.n77 VTAIL.n76 12.8005
R460 VTAIL.n82 VTAIL.n8 12.8005
R461 VTAIL.n138 VTAIL.n137 12.8005
R462 VTAIL.n179 VTAIL.n178 12.8005
R463 VTAIL.n184 VTAIL.n110 12.8005
R464 VTAIL.n240 VTAIL.n239 12.8005
R465 VTAIL.n281 VTAIL.n280 12.8005
R466 VTAIL.n286 VTAIL.n212 12.8005
R467 VTAIL.n694 VTAIL.n620 12.8005
R468 VTAIL.n689 VTAIL.n624 12.8005
R469 VTAIL.n649 VTAIL.n648 12.8005
R470 VTAIL.n592 VTAIL.n518 12.8005
R471 VTAIL.n587 VTAIL.n522 12.8005
R472 VTAIL.n547 VTAIL.n546 12.8005
R473 VTAIL.n490 VTAIL.n416 12.8005
R474 VTAIL.n485 VTAIL.n420 12.8005
R475 VTAIL.n445 VTAIL.n444 12.8005
R476 VTAIL.n388 VTAIL.n314 12.8005
R477 VTAIL.n383 VTAIL.n318 12.8005
R478 VTAIL.n343 VTAIL.n342 12.8005
R479 VTAIL.n753 VTAIL.n744 12.0247
R480 VTAIL.n789 VTAIL.n726 12.0247
R481 VTAIL.n800 VTAIL.n799 12.0247
R482 VTAIL.n39 VTAIL.n30 12.0247
R483 VTAIL.n75 VTAIL.n12 12.0247
R484 VTAIL.n86 VTAIL.n85 12.0247
R485 VTAIL.n141 VTAIL.n132 12.0247
R486 VTAIL.n177 VTAIL.n114 12.0247
R487 VTAIL.n188 VTAIL.n187 12.0247
R488 VTAIL.n243 VTAIL.n234 12.0247
R489 VTAIL.n279 VTAIL.n216 12.0247
R490 VTAIL.n290 VTAIL.n289 12.0247
R491 VTAIL.n698 VTAIL.n697 12.0247
R492 VTAIL.n688 VTAIL.n625 12.0247
R493 VTAIL.n652 VTAIL.n643 12.0247
R494 VTAIL.n596 VTAIL.n595 12.0247
R495 VTAIL.n586 VTAIL.n523 12.0247
R496 VTAIL.n550 VTAIL.n541 12.0247
R497 VTAIL.n494 VTAIL.n493 12.0247
R498 VTAIL.n484 VTAIL.n421 12.0247
R499 VTAIL.n448 VTAIL.n439 12.0247
R500 VTAIL.n392 VTAIL.n391 12.0247
R501 VTAIL.n382 VTAIL.n319 12.0247
R502 VTAIL.n346 VTAIL.n337 12.0247
R503 VTAIL.n754 VTAIL.n742 11.249
R504 VTAIL.n786 VTAIL.n785 11.249
R505 VTAIL.n803 VTAIL.n720 11.249
R506 VTAIL.n40 VTAIL.n28 11.249
R507 VTAIL.n72 VTAIL.n71 11.249
R508 VTAIL.n89 VTAIL.n6 11.249
R509 VTAIL.n142 VTAIL.n130 11.249
R510 VTAIL.n174 VTAIL.n173 11.249
R511 VTAIL.n191 VTAIL.n108 11.249
R512 VTAIL.n244 VTAIL.n232 11.249
R513 VTAIL.n276 VTAIL.n275 11.249
R514 VTAIL.n293 VTAIL.n210 11.249
R515 VTAIL.n701 VTAIL.n618 11.249
R516 VTAIL.n685 VTAIL.n684 11.249
R517 VTAIL.n653 VTAIL.n641 11.249
R518 VTAIL.n599 VTAIL.n516 11.249
R519 VTAIL.n583 VTAIL.n582 11.249
R520 VTAIL.n551 VTAIL.n539 11.249
R521 VTAIL.n497 VTAIL.n414 11.249
R522 VTAIL.n481 VTAIL.n480 11.249
R523 VTAIL.n449 VTAIL.n437 11.249
R524 VTAIL.n395 VTAIL.n312 11.249
R525 VTAIL.n379 VTAIL.n378 11.249
R526 VTAIL.n347 VTAIL.n335 11.249
R527 VTAIL.n758 VTAIL.n757 10.4732
R528 VTAIL.n782 VTAIL.n728 10.4732
R529 VTAIL.n804 VTAIL.n718 10.4732
R530 VTAIL.n44 VTAIL.n43 10.4732
R531 VTAIL.n68 VTAIL.n14 10.4732
R532 VTAIL.n90 VTAIL.n4 10.4732
R533 VTAIL.n146 VTAIL.n145 10.4732
R534 VTAIL.n170 VTAIL.n116 10.4732
R535 VTAIL.n192 VTAIL.n106 10.4732
R536 VTAIL.n248 VTAIL.n247 10.4732
R537 VTAIL.n272 VTAIL.n218 10.4732
R538 VTAIL.n294 VTAIL.n208 10.4732
R539 VTAIL.n702 VTAIL.n616 10.4732
R540 VTAIL.n681 VTAIL.n627 10.4732
R541 VTAIL.n657 VTAIL.n656 10.4732
R542 VTAIL.n600 VTAIL.n514 10.4732
R543 VTAIL.n579 VTAIL.n525 10.4732
R544 VTAIL.n555 VTAIL.n554 10.4732
R545 VTAIL.n498 VTAIL.n412 10.4732
R546 VTAIL.n477 VTAIL.n423 10.4732
R547 VTAIL.n453 VTAIL.n452 10.4732
R548 VTAIL.n396 VTAIL.n310 10.4732
R549 VTAIL.n375 VTAIL.n321 10.4732
R550 VTAIL.n351 VTAIL.n350 10.4732
R551 VTAIL.n761 VTAIL.n740 9.69747
R552 VTAIL.n781 VTAIL.n730 9.69747
R553 VTAIL.n808 VTAIL.n807 9.69747
R554 VTAIL.n47 VTAIL.n26 9.69747
R555 VTAIL.n67 VTAIL.n16 9.69747
R556 VTAIL.n94 VTAIL.n93 9.69747
R557 VTAIL.n149 VTAIL.n128 9.69747
R558 VTAIL.n169 VTAIL.n118 9.69747
R559 VTAIL.n196 VTAIL.n195 9.69747
R560 VTAIL.n251 VTAIL.n230 9.69747
R561 VTAIL.n271 VTAIL.n220 9.69747
R562 VTAIL.n298 VTAIL.n297 9.69747
R563 VTAIL.n706 VTAIL.n705 9.69747
R564 VTAIL.n680 VTAIL.n629 9.69747
R565 VTAIL.n660 VTAIL.n639 9.69747
R566 VTAIL.n604 VTAIL.n603 9.69747
R567 VTAIL.n578 VTAIL.n527 9.69747
R568 VTAIL.n558 VTAIL.n537 9.69747
R569 VTAIL.n502 VTAIL.n501 9.69747
R570 VTAIL.n476 VTAIL.n425 9.69747
R571 VTAIL.n456 VTAIL.n435 9.69747
R572 VTAIL.n400 VTAIL.n399 9.69747
R573 VTAIL.n374 VTAIL.n323 9.69747
R574 VTAIL.n354 VTAIL.n333 9.69747
R575 VTAIL.n814 VTAIL.n813 9.45567
R576 VTAIL.n100 VTAIL.n99 9.45567
R577 VTAIL.n202 VTAIL.n201 9.45567
R578 VTAIL.n304 VTAIL.n303 9.45567
R579 VTAIL.n712 VTAIL.n711 9.45567
R580 VTAIL.n610 VTAIL.n609 9.45567
R581 VTAIL.n508 VTAIL.n507 9.45567
R582 VTAIL.n406 VTAIL.n405 9.45567
R583 VTAIL.n813 VTAIL.n812 9.3005
R584 VTAIL.n716 VTAIL.n715 9.3005
R585 VTAIL.n807 VTAIL.n806 9.3005
R586 VTAIL.n805 VTAIL.n804 9.3005
R587 VTAIL.n720 VTAIL.n719 9.3005
R588 VTAIL.n799 VTAIL.n798 9.3005
R589 VTAIL.n797 VTAIL.n796 9.3005
R590 VTAIL.n736 VTAIL.n735 9.3005
R591 VTAIL.n765 VTAIL.n764 9.3005
R592 VTAIL.n763 VTAIL.n762 9.3005
R593 VTAIL.n740 VTAIL.n739 9.3005
R594 VTAIL.n757 VTAIL.n756 9.3005
R595 VTAIL.n755 VTAIL.n754 9.3005
R596 VTAIL.n744 VTAIL.n743 9.3005
R597 VTAIL.n749 VTAIL.n748 9.3005
R598 VTAIL.n771 VTAIL.n770 9.3005
R599 VTAIL.n773 VTAIL.n772 9.3005
R600 VTAIL.n732 VTAIL.n731 9.3005
R601 VTAIL.n779 VTAIL.n778 9.3005
R602 VTAIL.n781 VTAIL.n780 9.3005
R603 VTAIL.n728 VTAIL.n727 9.3005
R604 VTAIL.n787 VTAIL.n786 9.3005
R605 VTAIL.n789 VTAIL.n788 9.3005
R606 VTAIL.n790 VTAIL.n723 9.3005
R607 VTAIL.n99 VTAIL.n98 9.3005
R608 VTAIL.n2 VTAIL.n1 9.3005
R609 VTAIL.n93 VTAIL.n92 9.3005
R610 VTAIL.n91 VTAIL.n90 9.3005
R611 VTAIL.n6 VTAIL.n5 9.3005
R612 VTAIL.n85 VTAIL.n84 9.3005
R613 VTAIL.n83 VTAIL.n82 9.3005
R614 VTAIL.n22 VTAIL.n21 9.3005
R615 VTAIL.n51 VTAIL.n50 9.3005
R616 VTAIL.n49 VTAIL.n48 9.3005
R617 VTAIL.n26 VTAIL.n25 9.3005
R618 VTAIL.n43 VTAIL.n42 9.3005
R619 VTAIL.n41 VTAIL.n40 9.3005
R620 VTAIL.n30 VTAIL.n29 9.3005
R621 VTAIL.n35 VTAIL.n34 9.3005
R622 VTAIL.n57 VTAIL.n56 9.3005
R623 VTAIL.n59 VTAIL.n58 9.3005
R624 VTAIL.n18 VTAIL.n17 9.3005
R625 VTAIL.n65 VTAIL.n64 9.3005
R626 VTAIL.n67 VTAIL.n66 9.3005
R627 VTAIL.n14 VTAIL.n13 9.3005
R628 VTAIL.n73 VTAIL.n72 9.3005
R629 VTAIL.n75 VTAIL.n74 9.3005
R630 VTAIL.n76 VTAIL.n9 9.3005
R631 VTAIL.n201 VTAIL.n200 9.3005
R632 VTAIL.n104 VTAIL.n103 9.3005
R633 VTAIL.n195 VTAIL.n194 9.3005
R634 VTAIL.n193 VTAIL.n192 9.3005
R635 VTAIL.n108 VTAIL.n107 9.3005
R636 VTAIL.n187 VTAIL.n186 9.3005
R637 VTAIL.n185 VTAIL.n184 9.3005
R638 VTAIL.n124 VTAIL.n123 9.3005
R639 VTAIL.n153 VTAIL.n152 9.3005
R640 VTAIL.n151 VTAIL.n150 9.3005
R641 VTAIL.n128 VTAIL.n127 9.3005
R642 VTAIL.n145 VTAIL.n144 9.3005
R643 VTAIL.n143 VTAIL.n142 9.3005
R644 VTAIL.n132 VTAIL.n131 9.3005
R645 VTAIL.n137 VTAIL.n136 9.3005
R646 VTAIL.n159 VTAIL.n158 9.3005
R647 VTAIL.n161 VTAIL.n160 9.3005
R648 VTAIL.n120 VTAIL.n119 9.3005
R649 VTAIL.n167 VTAIL.n166 9.3005
R650 VTAIL.n169 VTAIL.n168 9.3005
R651 VTAIL.n116 VTAIL.n115 9.3005
R652 VTAIL.n175 VTAIL.n174 9.3005
R653 VTAIL.n177 VTAIL.n176 9.3005
R654 VTAIL.n178 VTAIL.n111 9.3005
R655 VTAIL.n303 VTAIL.n302 9.3005
R656 VTAIL.n206 VTAIL.n205 9.3005
R657 VTAIL.n297 VTAIL.n296 9.3005
R658 VTAIL.n295 VTAIL.n294 9.3005
R659 VTAIL.n210 VTAIL.n209 9.3005
R660 VTAIL.n289 VTAIL.n288 9.3005
R661 VTAIL.n287 VTAIL.n286 9.3005
R662 VTAIL.n226 VTAIL.n225 9.3005
R663 VTAIL.n255 VTAIL.n254 9.3005
R664 VTAIL.n253 VTAIL.n252 9.3005
R665 VTAIL.n230 VTAIL.n229 9.3005
R666 VTAIL.n247 VTAIL.n246 9.3005
R667 VTAIL.n245 VTAIL.n244 9.3005
R668 VTAIL.n234 VTAIL.n233 9.3005
R669 VTAIL.n239 VTAIL.n238 9.3005
R670 VTAIL.n261 VTAIL.n260 9.3005
R671 VTAIL.n263 VTAIL.n262 9.3005
R672 VTAIL.n222 VTAIL.n221 9.3005
R673 VTAIL.n269 VTAIL.n268 9.3005
R674 VTAIL.n271 VTAIL.n270 9.3005
R675 VTAIL.n218 VTAIL.n217 9.3005
R676 VTAIL.n277 VTAIL.n276 9.3005
R677 VTAIL.n279 VTAIL.n278 9.3005
R678 VTAIL.n280 VTAIL.n213 9.3005
R679 VTAIL.n672 VTAIL.n671 9.3005
R680 VTAIL.n631 VTAIL.n630 9.3005
R681 VTAIL.n678 VTAIL.n677 9.3005
R682 VTAIL.n680 VTAIL.n679 9.3005
R683 VTAIL.n627 VTAIL.n626 9.3005
R684 VTAIL.n686 VTAIL.n685 9.3005
R685 VTAIL.n688 VTAIL.n687 9.3005
R686 VTAIL.n624 VTAIL.n621 9.3005
R687 VTAIL.n711 VTAIL.n710 9.3005
R688 VTAIL.n614 VTAIL.n613 9.3005
R689 VTAIL.n705 VTAIL.n704 9.3005
R690 VTAIL.n703 VTAIL.n702 9.3005
R691 VTAIL.n618 VTAIL.n617 9.3005
R692 VTAIL.n697 VTAIL.n696 9.3005
R693 VTAIL.n695 VTAIL.n694 9.3005
R694 VTAIL.n670 VTAIL.n669 9.3005
R695 VTAIL.n635 VTAIL.n634 9.3005
R696 VTAIL.n664 VTAIL.n663 9.3005
R697 VTAIL.n662 VTAIL.n661 9.3005
R698 VTAIL.n639 VTAIL.n638 9.3005
R699 VTAIL.n656 VTAIL.n655 9.3005
R700 VTAIL.n654 VTAIL.n653 9.3005
R701 VTAIL.n643 VTAIL.n642 9.3005
R702 VTAIL.n648 VTAIL.n647 9.3005
R703 VTAIL.n570 VTAIL.n569 9.3005
R704 VTAIL.n529 VTAIL.n528 9.3005
R705 VTAIL.n576 VTAIL.n575 9.3005
R706 VTAIL.n578 VTAIL.n577 9.3005
R707 VTAIL.n525 VTAIL.n524 9.3005
R708 VTAIL.n584 VTAIL.n583 9.3005
R709 VTAIL.n586 VTAIL.n585 9.3005
R710 VTAIL.n522 VTAIL.n519 9.3005
R711 VTAIL.n609 VTAIL.n608 9.3005
R712 VTAIL.n512 VTAIL.n511 9.3005
R713 VTAIL.n603 VTAIL.n602 9.3005
R714 VTAIL.n601 VTAIL.n600 9.3005
R715 VTAIL.n516 VTAIL.n515 9.3005
R716 VTAIL.n595 VTAIL.n594 9.3005
R717 VTAIL.n593 VTAIL.n592 9.3005
R718 VTAIL.n568 VTAIL.n567 9.3005
R719 VTAIL.n533 VTAIL.n532 9.3005
R720 VTAIL.n562 VTAIL.n561 9.3005
R721 VTAIL.n560 VTAIL.n559 9.3005
R722 VTAIL.n537 VTAIL.n536 9.3005
R723 VTAIL.n554 VTAIL.n553 9.3005
R724 VTAIL.n552 VTAIL.n551 9.3005
R725 VTAIL.n541 VTAIL.n540 9.3005
R726 VTAIL.n546 VTAIL.n545 9.3005
R727 VTAIL.n468 VTAIL.n467 9.3005
R728 VTAIL.n427 VTAIL.n426 9.3005
R729 VTAIL.n474 VTAIL.n473 9.3005
R730 VTAIL.n476 VTAIL.n475 9.3005
R731 VTAIL.n423 VTAIL.n422 9.3005
R732 VTAIL.n482 VTAIL.n481 9.3005
R733 VTAIL.n484 VTAIL.n483 9.3005
R734 VTAIL.n420 VTAIL.n417 9.3005
R735 VTAIL.n507 VTAIL.n506 9.3005
R736 VTAIL.n410 VTAIL.n409 9.3005
R737 VTAIL.n501 VTAIL.n500 9.3005
R738 VTAIL.n499 VTAIL.n498 9.3005
R739 VTAIL.n414 VTAIL.n413 9.3005
R740 VTAIL.n493 VTAIL.n492 9.3005
R741 VTAIL.n491 VTAIL.n490 9.3005
R742 VTAIL.n466 VTAIL.n465 9.3005
R743 VTAIL.n431 VTAIL.n430 9.3005
R744 VTAIL.n460 VTAIL.n459 9.3005
R745 VTAIL.n458 VTAIL.n457 9.3005
R746 VTAIL.n435 VTAIL.n434 9.3005
R747 VTAIL.n452 VTAIL.n451 9.3005
R748 VTAIL.n450 VTAIL.n449 9.3005
R749 VTAIL.n439 VTAIL.n438 9.3005
R750 VTAIL.n444 VTAIL.n443 9.3005
R751 VTAIL.n366 VTAIL.n365 9.3005
R752 VTAIL.n325 VTAIL.n324 9.3005
R753 VTAIL.n372 VTAIL.n371 9.3005
R754 VTAIL.n374 VTAIL.n373 9.3005
R755 VTAIL.n321 VTAIL.n320 9.3005
R756 VTAIL.n380 VTAIL.n379 9.3005
R757 VTAIL.n382 VTAIL.n381 9.3005
R758 VTAIL.n318 VTAIL.n315 9.3005
R759 VTAIL.n405 VTAIL.n404 9.3005
R760 VTAIL.n308 VTAIL.n307 9.3005
R761 VTAIL.n399 VTAIL.n398 9.3005
R762 VTAIL.n397 VTAIL.n396 9.3005
R763 VTAIL.n312 VTAIL.n311 9.3005
R764 VTAIL.n391 VTAIL.n390 9.3005
R765 VTAIL.n389 VTAIL.n388 9.3005
R766 VTAIL.n364 VTAIL.n363 9.3005
R767 VTAIL.n329 VTAIL.n328 9.3005
R768 VTAIL.n358 VTAIL.n357 9.3005
R769 VTAIL.n356 VTAIL.n355 9.3005
R770 VTAIL.n333 VTAIL.n332 9.3005
R771 VTAIL.n350 VTAIL.n349 9.3005
R772 VTAIL.n348 VTAIL.n347 9.3005
R773 VTAIL.n337 VTAIL.n336 9.3005
R774 VTAIL.n342 VTAIL.n341 9.3005
R775 VTAIL.n762 VTAIL.n738 8.92171
R776 VTAIL.n778 VTAIL.n777 8.92171
R777 VTAIL.n811 VTAIL.n716 8.92171
R778 VTAIL.n48 VTAIL.n24 8.92171
R779 VTAIL.n64 VTAIL.n63 8.92171
R780 VTAIL.n97 VTAIL.n2 8.92171
R781 VTAIL.n150 VTAIL.n126 8.92171
R782 VTAIL.n166 VTAIL.n165 8.92171
R783 VTAIL.n199 VTAIL.n104 8.92171
R784 VTAIL.n252 VTAIL.n228 8.92171
R785 VTAIL.n268 VTAIL.n267 8.92171
R786 VTAIL.n301 VTAIL.n206 8.92171
R787 VTAIL.n709 VTAIL.n614 8.92171
R788 VTAIL.n677 VTAIL.n676 8.92171
R789 VTAIL.n661 VTAIL.n637 8.92171
R790 VTAIL.n607 VTAIL.n512 8.92171
R791 VTAIL.n575 VTAIL.n574 8.92171
R792 VTAIL.n559 VTAIL.n535 8.92171
R793 VTAIL.n505 VTAIL.n410 8.92171
R794 VTAIL.n473 VTAIL.n472 8.92171
R795 VTAIL.n457 VTAIL.n433 8.92171
R796 VTAIL.n403 VTAIL.n308 8.92171
R797 VTAIL.n371 VTAIL.n370 8.92171
R798 VTAIL.n355 VTAIL.n331 8.92171
R799 VTAIL.n766 VTAIL.n765 8.14595
R800 VTAIL.n774 VTAIL.n732 8.14595
R801 VTAIL.n812 VTAIL.n714 8.14595
R802 VTAIL.n52 VTAIL.n51 8.14595
R803 VTAIL.n60 VTAIL.n18 8.14595
R804 VTAIL.n98 VTAIL.n0 8.14595
R805 VTAIL.n154 VTAIL.n153 8.14595
R806 VTAIL.n162 VTAIL.n120 8.14595
R807 VTAIL.n200 VTAIL.n102 8.14595
R808 VTAIL.n256 VTAIL.n255 8.14595
R809 VTAIL.n264 VTAIL.n222 8.14595
R810 VTAIL.n302 VTAIL.n204 8.14595
R811 VTAIL.n710 VTAIL.n612 8.14595
R812 VTAIL.n673 VTAIL.n631 8.14595
R813 VTAIL.n665 VTAIL.n664 8.14595
R814 VTAIL.n608 VTAIL.n510 8.14595
R815 VTAIL.n571 VTAIL.n529 8.14595
R816 VTAIL.n563 VTAIL.n562 8.14595
R817 VTAIL.n506 VTAIL.n408 8.14595
R818 VTAIL.n469 VTAIL.n427 8.14595
R819 VTAIL.n461 VTAIL.n460 8.14595
R820 VTAIL.n404 VTAIL.n306 8.14595
R821 VTAIL.n367 VTAIL.n325 8.14595
R822 VTAIL.n359 VTAIL.n358 8.14595
R823 VTAIL.n769 VTAIL.n736 7.3702
R824 VTAIL.n773 VTAIL.n734 7.3702
R825 VTAIL.n55 VTAIL.n22 7.3702
R826 VTAIL.n59 VTAIL.n20 7.3702
R827 VTAIL.n157 VTAIL.n124 7.3702
R828 VTAIL.n161 VTAIL.n122 7.3702
R829 VTAIL.n259 VTAIL.n226 7.3702
R830 VTAIL.n263 VTAIL.n224 7.3702
R831 VTAIL.n672 VTAIL.n633 7.3702
R832 VTAIL.n668 VTAIL.n635 7.3702
R833 VTAIL.n570 VTAIL.n531 7.3702
R834 VTAIL.n566 VTAIL.n533 7.3702
R835 VTAIL.n468 VTAIL.n429 7.3702
R836 VTAIL.n464 VTAIL.n431 7.3702
R837 VTAIL.n366 VTAIL.n327 7.3702
R838 VTAIL.n362 VTAIL.n329 7.3702
R839 VTAIL.n770 VTAIL.n769 6.59444
R840 VTAIL.n770 VTAIL.n734 6.59444
R841 VTAIL.n56 VTAIL.n55 6.59444
R842 VTAIL.n56 VTAIL.n20 6.59444
R843 VTAIL.n158 VTAIL.n157 6.59444
R844 VTAIL.n158 VTAIL.n122 6.59444
R845 VTAIL.n260 VTAIL.n259 6.59444
R846 VTAIL.n260 VTAIL.n224 6.59444
R847 VTAIL.n669 VTAIL.n633 6.59444
R848 VTAIL.n669 VTAIL.n668 6.59444
R849 VTAIL.n567 VTAIL.n531 6.59444
R850 VTAIL.n567 VTAIL.n566 6.59444
R851 VTAIL.n465 VTAIL.n429 6.59444
R852 VTAIL.n465 VTAIL.n464 6.59444
R853 VTAIL.n363 VTAIL.n327 6.59444
R854 VTAIL.n363 VTAIL.n362 6.59444
R855 VTAIL.n766 VTAIL.n736 5.81868
R856 VTAIL.n774 VTAIL.n773 5.81868
R857 VTAIL.n814 VTAIL.n714 5.81868
R858 VTAIL.n52 VTAIL.n22 5.81868
R859 VTAIL.n60 VTAIL.n59 5.81868
R860 VTAIL.n100 VTAIL.n0 5.81868
R861 VTAIL.n154 VTAIL.n124 5.81868
R862 VTAIL.n162 VTAIL.n161 5.81868
R863 VTAIL.n202 VTAIL.n102 5.81868
R864 VTAIL.n256 VTAIL.n226 5.81868
R865 VTAIL.n264 VTAIL.n263 5.81868
R866 VTAIL.n304 VTAIL.n204 5.81868
R867 VTAIL.n712 VTAIL.n612 5.81868
R868 VTAIL.n673 VTAIL.n672 5.81868
R869 VTAIL.n665 VTAIL.n635 5.81868
R870 VTAIL.n610 VTAIL.n510 5.81868
R871 VTAIL.n571 VTAIL.n570 5.81868
R872 VTAIL.n563 VTAIL.n533 5.81868
R873 VTAIL.n508 VTAIL.n408 5.81868
R874 VTAIL.n469 VTAIL.n468 5.81868
R875 VTAIL.n461 VTAIL.n431 5.81868
R876 VTAIL.n406 VTAIL.n306 5.81868
R877 VTAIL.n367 VTAIL.n366 5.81868
R878 VTAIL.n359 VTAIL.n329 5.81868
R879 VTAIL.n765 VTAIL.n738 5.04292
R880 VTAIL.n777 VTAIL.n732 5.04292
R881 VTAIL.n812 VTAIL.n811 5.04292
R882 VTAIL.n51 VTAIL.n24 5.04292
R883 VTAIL.n63 VTAIL.n18 5.04292
R884 VTAIL.n98 VTAIL.n97 5.04292
R885 VTAIL.n153 VTAIL.n126 5.04292
R886 VTAIL.n165 VTAIL.n120 5.04292
R887 VTAIL.n200 VTAIL.n199 5.04292
R888 VTAIL.n255 VTAIL.n228 5.04292
R889 VTAIL.n267 VTAIL.n222 5.04292
R890 VTAIL.n302 VTAIL.n301 5.04292
R891 VTAIL.n710 VTAIL.n709 5.04292
R892 VTAIL.n676 VTAIL.n631 5.04292
R893 VTAIL.n664 VTAIL.n637 5.04292
R894 VTAIL.n608 VTAIL.n607 5.04292
R895 VTAIL.n574 VTAIL.n529 5.04292
R896 VTAIL.n562 VTAIL.n535 5.04292
R897 VTAIL.n506 VTAIL.n505 5.04292
R898 VTAIL.n472 VTAIL.n427 5.04292
R899 VTAIL.n460 VTAIL.n433 5.04292
R900 VTAIL.n404 VTAIL.n403 5.04292
R901 VTAIL.n370 VTAIL.n325 5.04292
R902 VTAIL.n358 VTAIL.n331 5.04292
R903 VTAIL.n762 VTAIL.n761 4.26717
R904 VTAIL.n778 VTAIL.n730 4.26717
R905 VTAIL.n808 VTAIL.n716 4.26717
R906 VTAIL.n48 VTAIL.n47 4.26717
R907 VTAIL.n64 VTAIL.n16 4.26717
R908 VTAIL.n94 VTAIL.n2 4.26717
R909 VTAIL.n150 VTAIL.n149 4.26717
R910 VTAIL.n166 VTAIL.n118 4.26717
R911 VTAIL.n196 VTAIL.n104 4.26717
R912 VTAIL.n252 VTAIL.n251 4.26717
R913 VTAIL.n268 VTAIL.n220 4.26717
R914 VTAIL.n298 VTAIL.n206 4.26717
R915 VTAIL.n706 VTAIL.n614 4.26717
R916 VTAIL.n677 VTAIL.n629 4.26717
R917 VTAIL.n661 VTAIL.n660 4.26717
R918 VTAIL.n604 VTAIL.n512 4.26717
R919 VTAIL.n575 VTAIL.n527 4.26717
R920 VTAIL.n559 VTAIL.n558 4.26717
R921 VTAIL.n502 VTAIL.n410 4.26717
R922 VTAIL.n473 VTAIL.n425 4.26717
R923 VTAIL.n457 VTAIL.n456 4.26717
R924 VTAIL.n400 VTAIL.n308 4.26717
R925 VTAIL.n371 VTAIL.n323 4.26717
R926 VTAIL.n355 VTAIL.n354 4.26717
R927 VTAIL.n748 VTAIL.n747 3.70982
R928 VTAIL.n34 VTAIL.n33 3.70982
R929 VTAIL.n136 VTAIL.n135 3.70982
R930 VTAIL.n238 VTAIL.n237 3.70982
R931 VTAIL.n647 VTAIL.n646 3.70982
R932 VTAIL.n545 VTAIL.n544 3.70982
R933 VTAIL.n443 VTAIL.n442 3.70982
R934 VTAIL.n341 VTAIL.n340 3.70982
R935 VTAIL.n758 VTAIL.n740 3.49141
R936 VTAIL.n782 VTAIL.n781 3.49141
R937 VTAIL.n807 VTAIL.n718 3.49141
R938 VTAIL.n44 VTAIL.n26 3.49141
R939 VTAIL.n68 VTAIL.n67 3.49141
R940 VTAIL.n93 VTAIL.n4 3.49141
R941 VTAIL.n146 VTAIL.n128 3.49141
R942 VTAIL.n170 VTAIL.n169 3.49141
R943 VTAIL.n195 VTAIL.n106 3.49141
R944 VTAIL.n248 VTAIL.n230 3.49141
R945 VTAIL.n272 VTAIL.n271 3.49141
R946 VTAIL.n297 VTAIL.n208 3.49141
R947 VTAIL.n705 VTAIL.n616 3.49141
R948 VTAIL.n681 VTAIL.n680 3.49141
R949 VTAIL.n657 VTAIL.n639 3.49141
R950 VTAIL.n603 VTAIL.n514 3.49141
R951 VTAIL.n579 VTAIL.n578 3.49141
R952 VTAIL.n555 VTAIL.n537 3.49141
R953 VTAIL.n501 VTAIL.n412 3.49141
R954 VTAIL.n477 VTAIL.n476 3.49141
R955 VTAIL.n453 VTAIL.n435 3.49141
R956 VTAIL.n399 VTAIL.n310 3.49141
R957 VTAIL.n375 VTAIL.n374 3.49141
R958 VTAIL.n351 VTAIL.n333 3.49141
R959 VTAIL.n757 VTAIL.n742 2.71565
R960 VTAIL.n785 VTAIL.n728 2.71565
R961 VTAIL.n804 VTAIL.n803 2.71565
R962 VTAIL.n43 VTAIL.n28 2.71565
R963 VTAIL.n71 VTAIL.n14 2.71565
R964 VTAIL.n90 VTAIL.n89 2.71565
R965 VTAIL.n145 VTAIL.n130 2.71565
R966 VTAIL.n173 VTAIL.n116 2.71565
R967 VTAIL.n192 VTAIL.n191 2.71565
R968 VTAIL.n247 VTAIL.n232 2.71565
R969 VTAIL.n275 VTAIL.n218 2.71565
R970 VTAIL.n294 VTAIL.n293 2.71565
R971 VTAIL.n702 VTAIL.n701 2.71565
R972 VTAIL.n684 VTAIL.n627 2.71565
R973 VTAIL.n656 VTAIL.n641 2.71565
R974 VTAIL.n600 VTAIL.n599 2.71565
R975 VTAIL.n582 VTAIL.n525 2.71565
R976 VTAIL.n554 VTAIL.n539 2.71565
R977 VTAIL.n498 VTAIL.n497 2.71565
R978 VTAIL.n480 VTAIL.n423 2.71565
R979 VTAIL.n452 VTAIL.n437 2.71565
R980 VTAIL.n396 VTAIL.n395 2.71565
R981 VTAIL.n378 VTAIL.n321 2.71565
R982 VTAIL.n350 VTAIL.n335 2.71565
R983 VTAIL.n754 VTAIL.n753 1.93989
R984 VTAIL.n786 VTAIL.n726 1.93989
R985 VTAIL.n800 VTAIL.n720 1.93989
R986 VTAIL.n40 VTAIL.n39 1.93989
R987 VTAIL.n72 VTAIL.n12 1.93989
R988 VTAIL.n86 VTAIL.n6 1.93989
R989 VTAIL.n142 VTAIL.n141 1.93989
R990 VTAIL.n174 VTAIL.n114 1.93989
R991 VTAIL.n188 VTAIL.n108 1.93989
R992 VTAIL.n244 VTAIL.n243 1.93989
R993 VTAIL.n276 VTAIL.n216 1.93989
R994 VTAIL.n290 VTAIL.n210 1.93989
R995 VTAIL.n698 VTAIL.n618 1.93989
R996 VTAIL.n685 VTAIL.n625 1.93989
R997 VTAIL.n653 VTAIL.n652 1.93989
R998 VTAIL.n596 VTAIL.n516 1.93989
R999 VTAIL.n583 VTAIL.n523 1.93989
R1000 VTAIL.n551 VTAIL.n550 1.93989
R1001 VTAIL.n494 VTAIL.n414 1.93989
R1002 VTAIL.n481 VTAIL.n421 1.93989
R1003 VTAIL.n449 VTAIL.n448 1.93989
R1004 VTAIL.n392 VTAIL.n312 1.93989
R1005 VTAIL.n379 VTAIL.n319 1.93989
R1006 VTAIL.n347 VTAIL.n346 1.93989
R1007 VTAIL.n750 VTAIL.n744 1.16414
R1008 VTAIL.n791 VTAIL.n789 1.16414
R1009 VTAIL.n799 VTAIL.n722 1.16414
R1010 VTAIL.n36 VTAIL.n30 1.16414
R1011 VTAIL.n77 VTAIL.n75 1.16414
R1012 VTAIL.n85 VTAIL.n8 1.16414
R1013 VTAIL.n138 VTAIL.n132 1.16414
R1014 VTAIL.n179 VTAIL.n177 1.16414
R1015 VTAIL.n187 VTAIL.n110 1.16414
R1016 VTAIL.n240 VTAIL.n234 1.16414
R1017 VTAIL.n281 VTAIL.n279 1.16414
R1018 VTAIL.n289 VTAIL.n212 1.16414
R1019 VTAIL.n697 VTAIL.n620 1.16414
R1020 VTAIL.n689 VTAIL.n688 1.16414
R1021 VTAIL.n649 VTAIL.n643 1.16414
R1022 VTAIL.n595 VTAIL.n518 1.16414
R1023 VTAIL.n587 VTAIL.n586 1.16414
R1024 VTAIL.n547 VTAIL.n541 1.16414
R1025 VTAIL.n493 VTAIL.n416 1.16414
R1026 VTAIL.n485 VTAIL.n484 1.16414
R1027 VTAIL.n445 VTAIL.n439 1.16414
R1028 VTAIL.n391 VTAIL.n314 1.16414
R1029 VTAIL.n383 VTAIL.n382 1.16414
R1030 VTAIL.n343 VTAIL.n337 1.16414
R1031 VTAIL.n509 VTAIL.n407 1.06947
R1032 VTAIL.n713 VTAIL.n611 1.06947
R1033 VTAIL.n305 VTAIL.n203 1.06947
R1034 VTAIL VTAIL.n101 0.593172
R1035 VTAIL VTAIL.n815 0.476793
R1036 VTAIL.n611 VTAIL.n509 0.470328
R1037 VTAIL.n203 VTAIL.n101 0.470328
R1038 VTAIL.n749 VTAIL.n746 0.388379
R1039 VTAIL.n790 VTAIL.n724 0.388379
R1040 VTAIL.n796 VTAIL.n795 0.388379
R1041 VTAIL.n35 VTAIL.n32 0.388379
R1042 VTAIL.n76 VTAIL.n10 0.388379
R1043 VTAIL.n82 VTAIL.n81 0.388379
R1044 VTAIL.n137 VTAIL.n134 0.388379
R1045 VTAIL.n178 VTAIL.n112 0.388379
R1046 VTAIL.n184 VTAIL.n183 0.388379
R1047 VTAIL.n239 VTAIL.n236 0.388379
R1048 VTAIL.n280 VTAIL.n214 0.388379
R1049 VTAIL.n286 VTAIL.n285 0.388379
R1050 VTAIL.n694 VTAIL.n693 0.388379
R1051 VTAIL.n624 VTAIL.n622 0.388379
R1052 VTAIL.n648 VTAIL.n645 0.388379
R1053 VTAIL.n592 VTAIL.n591 0.388379
R1054 VTAIL.n522 VTAIL.n520 0.388379
R1055 VTAIL.n546 VTAIL.n543 0.388379
R1056 VTAIL.n490 VTAIL.n489 0.388379
R1057 VTAIL.n420 VTAIL.n418 0.388379
R1058 VTAIL.n444 VTAIL.n441 0.388379
R1059 VTAIL.n388 VTAIL.n387 0.388379
R1060 VTAIL.n318 VTAIL.n316 0.388379
R1061 VTAIL.n342 VTAIL.n339 0.388379
R1062 VTAIL.n748 VTAIL.n743 0.155672
R1063 VTAIL.n755 VTAIL.n743 0.155672
R1064 VTAIL.n756 VTAIL.n755 0.155672
R1065 VTAIL.n756 VTAIL.n739 0.155672
R1066 VTAIL.n763 VTAIL.n739 0.155672
R1067 VTAIL.n764 VTAIL.n763 0.155672
R1068 VTAIL.n764 VTAIL.n735 0.155672
R1069 VTAIL.n771 VTAIL.n735 0.155672
R1070 VTAIL.n772 VTAIL.n771 0.155672
R1071 VTAIL.n772 VTAIL.n731 0.155672
R1072 VTAIL.n779 VTAIL.n731 0.155672
R1073 VTAIL.n780 VTAIL.n779 0.155672
R1074 VTAIL.n780 VTAIL.n727 0.155672
R1075 VTAIL.n787 VTAIL.n727 0.155672
R1076 VTAIL.n788 VTAIL.n787 0.155672
R1077 VTAIL.n788 VTAIL.n723 0.155672
R1078 VTAIL.n797 VTAIL.n723 0.155672
R1079 VTAIL.n798 VTAIL.n797 0.155672
R1080 VTAIL.n798 VTAIL.n719 0.155672
R1081 VTAIL.n805 VTAIL.n719 0.155672
R1082 VTAIL.n806 VTAIL.n805 0.155672
R1083 VTAIL.n806 VTAIL.n715 0.155672
R1084 VTAIL.n813 VTAIL.n715 0.155672
R1085 VTAIL.n34 VTAIL.n29 0.155672
R1086 VTAIL.n41 VTAIL.n29 0.155672
R1087 VTAIL.n42 VTAIL.n41 0.155672
R1088 VTAIL.n42 VTAIL.n25 0.155672
R1089 VTAIL.n49 VTAIL.n25 0.155672
R1090 VTAIL.n50 VTAIL.n49 0.155672
R1091 VTAIL.n50 VTAIL.n21 0.155672
R1092 VTAIL.n57 VTAIL.n21 0.155672
R1093 VTAIL.n58 VTAIL.n57 0.155672
R1094 VTAIL.n58 VTAIL.n17 0.155672
R1095 VTAIL.n65 VTAIL.n17 0.155672
R1096 VTAIL.n66 VTAIL.n65 0.155672
R1097 VTAIL.n66 VTAIL.n13 0.155672
R1098 VTAIL.n73 VTAIL.n13 0.155672
R1099 VTAIL.n74 VTAIL.n73 0.155672
R1100 VTAIL.n74 VTAIL.n9 0.155672
R1101 VTAIL.n83 VTAIL.n9 0.155672
R1102 VTAIL.n84 VTAIL.n83 0.155672
R1103 VTAIL.n84 VTAIL.n5 0.155672
R1104 VTAIL.n91 VTAIL.n5 0.155672
R1105 VTAIL.n92 VTAIL.n91 0.155672
R1106 VTAIL.n92 VTAIL.n1 0.155672
R1107 VTAIL.n99 VTAIL.n1 0.155672
R1108 VTAIL.n136 VTAIL.n131 0.155672
R1109 VTAIL.n143 VTAIL.n131 0.155672
R1110 VTAIL.n144 VTAIL.n143 0.155672
R1111 VTAIL.n144 VTAIL.n127 0.155672
R1112 VTAIL.n151 VTAIL.n127 0.155672
R1113 VTAIL.n152 VTAIL.n151 0.155672
R1114 VTAIL.n152 VTAIL.n123 0.155672
R1115 VTAIL.n159 VTAIL.n123 0.155672
R1116 VTAIL.n160 VTAIL.n159 0.155672
R1117 VTAIL.n160 VTAIL.n119 0.155672
R1118 VTAIL.n167 VTAIL.n119 0.155672
R1119 VTAIL.n168 VTAIL.n167 0.155672
R1120 VTAIL.n168 VTAIL.n115 0.155672
R1121 VTAIL.n175 VTAIL.n115 0.155672
R1122 VTAIL.n176 VTAIL.n175 0.155672
R1123 VTAIL.n176 VTAIL.n111 0.155672
R1124 VTAIL.n185 VTAIL.n111 0.155672
R1125 VTAIL.n186 VTAIL.n185 0.155672
R1126 VTAIL.n186 VTAIL.n107 0.155672
R1127 VTAIL.n193 VTAIL.n107 0.155672
R1128 VTAIL.n194 VTAIL.n193 0.155672
R1129 VTAIL.n194 VTAIL.n103 0.155672
R1130 VTAIL.n201 VTAIL.n103 0.155672
R1131 VTAIL.n238 VTAIL.n233 0.155672
R1132 VTAIL.n245 VTAIL.n233 0.155672
R1133 VTAIL.n246 VTAIL.n245 0.155672
R1134 VTAIL.n246 VTAIL.n229 0.155672
R1135 VTAIL.n253 VTAIL.n229 0.155672
R1136 VTAIL.n254 VTAIL.n253 0.155672
R1137 VTAIL.n254 VTAIL.n225 0.155672
R1138 VTAIL.n261 VTAIL.n225 0.155672
R1139 VTAIL.n262 VTAIL.n261 0.155672
R1140 VTAIL.n262 VTAIL.n221 0.155672
R1141 VTAIL.n269 VTAIL.n221 0.155672
R1142 VTAIL.n270 VTAIL.n269 0.155672
R1143 VTAIL.n270 VTAIL.n217 0.155672
R1144 VTAIL.n277 VTAIL.n217 0.155672
R1145 VTAIL.n278 VTAIL.n277 0.155672
R1146 VTAIL.n278 VTAIL.n213 0.155672
R1147 VTAIL.n287 VTAIL.n213 0.155672
R1148 VTAIL.n288 VTAIL.n287 0.155672
R1149 VTAIL.n288 VTAIL.n209 0.155672
R1150 VTAIL.n295 VTAIL.n209 0.155672
R1151 VTAIL.n296 VTAIL.n295 0.155672
R1152 VTAIL.n296 VTAIL.n205 0.155672
R1153 VTAIL.n303 VTAIL.n205 0.155672
R1154 VTAIL.n711 VTAIL.n613 0.155672
R1155 VTAIL.n704 VTAIL.n613 0.155672
R1156 VTAIL.n704 VTAIL.n703 0.155672
R1157 VTAIL.n703 VTAIL.n617 0.155672
R1158 VTAIL.n696 VTAIL.n617 0.155672
R1159 VTAIL.n696 VTAIL.n695 0.155672
R1160 VTAIL.n695 VTAIL.n621 0.155672
R1161 VTAIL.n687 VTAIL.n621 0.155672
R1162 VTAIL.n687 VTAIL.n686 0.155672
R1163 VTAIL.n686 VTAIL.n626 0.155672
R1164 VTAIL.n679 VTAIL.n626 0.155672
R1165 VTAIL.n679 VTAIL.n678 0.155672
R1166 VTAIL.n678 VTAIL.n630 0.155672
R1167 VTAIL.n671 VTAIL.n630 0.155672
R1168 VTAIL.n671 VTAIL.n670 0.155672
R1169 VTAIL.n670 VTAIL.n634 0.155672
R1170 VTAIL.n663 VTAIL.n634 0.155672
R1171 VTAIL.n663 VTAIL.n662 0.155672
R1172 VTAIL.n662 VTAIL.n638 0.155672
R1173 VTAIL.n655 VTAIL.n638 0.155672
R1174 VTAIL.n655 VTAIL.n654 0.155672
R1175 VTAIL.n654 VTAIL.n642 0.155672
R1176 VTAIL.n647 VTAIL.n642 0.155672
R1177 VTAIL.n609 VTAIL.n511 0.155672
R1178 VTAIL.n602 VTAIL.n511 0.155672
R1179 VTAIL.n602 VTAIL.n601 0.155672
R1180 VTAIL.n601 VTAIL.n515 0.155672
R1181 VTAIL.n594 VTAIL.n515 0.155672
R1182 VTAIL.n594 VTAIL.n593 0.155672
R1183 VTAIL.n593 VTAIL.n519 0.155672
R1184 VTAIL.n585 VTAIL.n519 0.155672
R1185 VTAIL.n585 VTAIL.n584 0.155672
R1186 VTAIL.n584 VTAIL.n524 0.155672
R1187 VTAIL.n577 VTAIL.n524 0.155672
R1188 VTAIL.n577 VTAIL.n576 0.155672
R1189 VTAIL.n576 VTAIL.n528 0.155672
R1190 VTAIL.n569 VTAIL.n528 0.155672
R1191 VTAIL.n569 VTAIL.n568 0.155672
R1192 VTAIL.n568 VTAIL.n532 0.155672
R1193 VTAIL.n561 VTAIL.n532 0.155672
R1194 VTAIL.n561 VTAIL.n560 0.155672
R1195 VTAIL.n560 VTAIL.n536 0.155672
R1196 VTAIL.n553 VTAIL.n536 0.155672
R1197 VTAIL.n553 VTAIL.n552 0.155672
R1198 VTAIL.n552 VTAIL.n540 0.155672
R1199 VTAIL.n545 VTAIL.n540 0.155672
R1200 VTAIL.n507 VTAIL.n409 0.155672
R1201 VTAIL.n500 VTAIL.n409 0.155672
R1202 VTAIL.n500 VTAIL.n499 0.155672
R1203 VTAIL.n499 VTAIL.n413 0.155672
R1204 VTAIL.n492 VTAIL.n413 0.155672
R1205 VTAIL.n492 VTAIL.n491 0.155672
R1206 VTAIL.n491 VTAIL.n417 0.155672
R1207 VTAIL.n483 VTAIL.n417 0.155672
R1208 VTAIL.n483 VTAIL.n482 0.155672
R1209 VTAIL.n482 VTAIL.n422 0.155672
R1210 VTAIL.n475 VTAIL.n422 0.155672
R1211 VTAIL.n475 VTAIL.n474 0.155672
R1212 VTAIL.n474 VTAIL.n426 0.155672
R1213 VTAIL.n467 VTAIL.n426 0.155672
R1214 VTAIL.n467 VTAIL.n466 0.155672
R1215 VTAIL.n466 VTAIL.n430 0.155672
R1216 VTAIL.n459 VTAIL.n430 0.155672
R1217 VTAIL.n459 VTAIL.n458 0.155672
R1218 VTAIL.n458 VTAIL.n434 0.155672
R1219 VTAIL.n451 VTAIL.n434 0.155672
R1220 VTAIL.n451 VTAIL.n450 0.155672
R1221 VTAIL.n450 VTAIL.n438 0.155672
R1222 VTAIL.n443 VTAIL.n438 0.155672
R1223 VTAIL.n405 VTAIL.n307 0.155672
R1224 VTAIL.n398 VTAIL.n307 0.155672
R1225 VTAIL.n398 VTAIL.n397 0.155672
R1226 VTAIL.n397 VTAIL.n311 0.155672
R1227 VTAIL.n390 VTAIL.n311 0.155672
R1228 VTAIL.n390 VTAIL.n389 0.155672
R1229 VTAIL.n389 VTAIL.n315 0.155672
R1230 VTAIL.n381 VTAIL.n315 0.155672
R1231 VTAIL.n381 VTAIL.n380 0.155672
R1232 VTAIL.n380 VTAIL.n320 0.155672
R1233 VTAIL.n373 VTAIL.n320 0.155672
R1234 VTAIL.n373 VTAIL.n372 0.155672
R1235 VTAIL.n372 VTAIL.n324 0.155672
R1236 VTAIL.n365 VTAIL.n324 0.155672
R1237 VTAIL.n365 VTAIL.n364 0.155672
R1238 VTAIL.n364 VTAIL.n328 0.155672
R1239 VTAIL.n357 VTAIL.n328 0.155672
R1240 VTAIL.n357 VTAIL.n356 0.155672
R1241 VTAIL.n356 VTAIL.n332 0.155672
R1242 VTAIL.n349 VTAIL.n332 0.155672
R1243 VTAIL.n349 VTAIL.n348 0.155672
R1244 VTAIL.n348 VTAIL.n336 0.155672
R1245 VTAIL.n341 VTAIL.n336 0.155672
R1246 VP.n0 VP.t1 544.835
R1247 VP.n0 VP.t0 544.747
R1248 VP.n2 VP.t3 526.227
R1249 VP.n3 VP.t2 526.227
R1250 VP.n4 VP.n3 80.6037
R1251 VP.n2 VP.n1 80.6037
R1252 VP.n1 VP.n0 77.0486
R1253 VP.n3 VP.n2 48.2005
R1254 VP.n4 VP.n1 0.380177
R1255 VP VP.n4 0.146778
R1256 VDD1 VDD1.n1 111.859
R1257 VDD1 VDD1.n0 68.7459
R1258 VDD1.n0 VDD1.t2 1.78257
R1259 VDD1.n0 VDD1.t3 1.78257
R1260 VDD1.n1 VDD1.t0 1.78257
R1261 VDD1.n1 VDD1.t1 1.78257
R1262 B.n131 B.t6 685.335
R1263 B.n139 B.t3 685.335
R1264 B.n42 B.t0 685.335
R1265 B.n50 B.t9 685.335
R1266 B.n462 B.n81 585
R1267 B.n464 B.n463 585
R1268 B.n465 B.n80 585
R1269 B.n467 B.n466 585
R1270 B.n468 B.n79 585
R1271 B.n470 B.n469 585
R1272 B.n471 B.n78 585
R1273 B.n473 B.n472 585
R1274 B.n474 B.n77 585
R1275 B.n476 B.n475 585
R1276 B.n477 B.n76 585
R1277 B.n479 B.n478 585
R1278 B.n480 B.n75 585
R1279 B.n482 B.n481 585
R1280 B.n483 B.n74 585
R1281 B.n485 B.n484 585
R1282 B.n486 B.n73 585
R1283 B.n488 B.n487 585
R1284 B.n489 B.n72 585
R1285 B.n491 B.n490 585
R1286 B.n492 B.n71 585
R1287 B.n494 B.n493 585
R1288 B.n495 B.n70 585
R1289 B.n497 B.n496 585
R1290 B.n498 B.n69 585
R1291 B.n500 B.n499 585
R1292 B.n501 B.n68 585
R1293 B.n503 B.n502 585
R1294 B.n504 B.n67 585
R1295 B.n506 B.n505 585
R1296 B.n507 B.n66 585
R1297 B.n509 B.n508 585
R1298 B.n510 B.n65 585
R1299 B.n512 B.n511 585
R1300 B.n513 B.n64 585
R1301 B.n515 B.n514 585
R1302 B.n516 B.n63 585
R1303 B.n518 B.n517 585
R1304 B.n519 B.n62 585
R1305 B.n521 B.n520 585
R1306 B.n522 B.n61 585
R1307 B.n524 B.n523 585
R1308 B.n525 B.n60 585
R1309 B.n527 B.n526 585
R1310 B.n528 B.n59 585
R1311 B.n530 B.n529 585
R1312 B.n531 B.n58 585
R1313 B.n533 B.n532 585
R1314 B.n534 B.n57 585
R1315 B.n536 B.n535 585
R1316 B.n537 B.n56 585
R1317 B.n539 B.n538 585
R1318 B.n540 B.n55 585
R1319 B.n542 B.n541 585
R1320 B.n543 B.n54 585
R1321 B.n545 B.n544 585
R1322 B.n546 B.n53 585
R1323 B.n548 B.n547 585
R1324 B.n549 B.n49 585
R1325 B.n551 B.n550 585
R1326 B.n552 B.n48 585
R1327 B.n554 B.n553 585
R1328 B.n555 B.n47 585
R1329 B.n557 B.n556 585
R1330 B.n558 B.n46 585
R1331 B.n560 B.n559 585
R1332 B.n561 B.n45 585
R1333 B.n563 B.n562 585
R1334 B.n564 B.n44 585
R1335 B.n566 B.n565 585
R1336 B.n568 B.n41 585
R1337 B.n570 B.n569 585
R1338 B.n571 B.n40 585
R1339 B.n573 B.n572 585
R1340 B.n574 B.n39 585
R1341 B.n576 B.n575 585
R1342 B.n577 B.n38 585
R1343 B.n579 B.n578 585
R1344 B.n580 B.n37 585
R1345 B.n582 B.n581 585
R1346 B.n583 B.n36 585
R1347 B.n585 B.n584 585
R1348 B.n586 B.n35 585
R1349 B.n588 B.n587 585
R1350 B.n589 B.n34 585
R1351 B.n591 B.n590 585
R1352 B.n592 B.n33 585
R1353 B.n594 B.n593 585
R1354 B.n595 B.n32 585
R1355 B.n597 B.n596 585
R1356 B.n598 B.n31 585
R1357 B.n600 B.n599 585
R1358 B.n601 B.n30 585
R1359 B.n603 B.n602 585
R1360 B.n604 B.n29 585
R1361 B.n606 B.n605 585
R1362 B.n607 B.n28 585
R1363 B.n609 B.n608 585
R1364 B.n610 B.n27 585
R1365 B.n612 B.n611 585
R1366 B.n613 B.n26 585
R1367 B.n615 B.n614 585
R1368 B.n616 B.n25 585
R1369 B.n618 B.n617 585
R1370 B.n619 B.n24 585
R1371 B.n621 B.n620 585
R1372 B.n622 B.n23 585
R1373 B.n624 B.n623 585
R1374 B.n625 B.n22 585
R1375 B.n627 B.n626 585
R1376 B.n628 B.n21 585
R1377 B.n630 B.n629 585
R1378 B.n631 B.n20 585
R1379 B.n633 B.n632 585
R1380 B.n634 B.n19 585
R1381 B.n636 B.n635 585
R1382 B.n637 B.n18 585
R1383 B.n639 B.n638 585
R1384 B.n640 B.n17 585
R1385 B.n642 B.n641 585
R1386 B.n643 B.n16 585
R1387 B.n645 B.n644 585
R1388 B.n646 B.n15 585
R1389 B.n648 B.n647 585
R1390 B.n649 B.n14 585
R1391 B.n651 B.n650 585
R1392 B.n652 B.n13 585
R1393 B.n654 B.n653 585
R1394 B.n655 B.n12 585
R1395 B.n657 B.n656 585
R1396 B.n461 B.n460 585
R1397 B.n459 B.n82 585
R1398 B.n458 B.n457 585
R1399 B.n456 B.n83 585
R1400 B.n455 B.n454 585
R1401 B.n453 B.n84 585
R1402 B.n452 B.n451 585
R1403 B.n450 B.n85 585
R1404 B.n449 B.n448 585
R1405 B.n447 B.n86 585
R1406 B.n446 B.n445 585
R1407 B.n444 B.n87 585
R1408 B.n443 B.n442 585
R1409 B.n441 B.n88 585
R1410 B.n440 B.n439 585
R1411 B.n438 B.n89 585
R1412 B.n437 B.n436 585
R1413 B.n435 B.n90 585
R1414 B.n434 B.n433 585
R1415 B.n432 B.n91 585
R1416 B.n431 B.n430 585
R1417 B.n429 B.n92 585
R1418 B.n428 B.n427 585
R1419 B.n426 B.n93 585
R1420 B.n425 B.n424 585
R1421 B.n423 B.n94 585
R1422 B.n422 B.n421 585
R1423 B.n420 B.n95 585
R1424 B.n419 B.n418 585
R1425 B.n417 B.n96 585
R1426 B.n416 B.n415 585
R1427 B.n414 B.n97 585
R1428 B.n413 B.n412 585
R1429 B.n411 B.n98 585
R1430 B.n410 B.n409 585
R1431 B.n408 B.n99 585
R1432 B.n407 B.n406 585
R1433 B.n405 B.n100 585
R1434 B.n404 B.n403 585
R1435 B.n207 B.n170 585
R1436 B.n209 B.n208 585
R1437 B.n210 B.n169 585
R1438 B.n212 B.n211 585
R1439 B.n213 B.n168 585
R1440 B.n215 B.n214 585
R1441 B.n216 B.n167 585
R1442 B.n218 B.n217 585
R1443 B.n219 B.n166 585
R1444 B.n221 B.n220 585
R1445 B.n222 B.n165 585
R1446 B.n224 B.n223 585
R1447 B.n225 B.n164 585
R1448 B.n227 B.n226 585
R1449 B.n228 B.n163 585
R1450 B.n230 B.n229 585
R1451 B.n231 B.n162 585
R1452 B.n233 B.n232 585
R1453 B.n234 B.n161 585
R1454 B.n236 B.n235 585
R1455 B.n237 B.n160 585
R1456 B.n239 B.n238 585
R1457 B.n240 B.n159 585
R1458 B.n242 B.n241 585
R1459 B.n243 B.n158 585
R1460 B.n245 B.n244 585
R1461 B.n246 B.n157 585
R1462 B.n248 B.n247 585
R1463 B.n249 B.n156 585
R1464 B.n251 B.n250 585
R1465 B.n252 B.n155 585
R1466 B.n254 B.n253 585
R1467 B.n255 B.n154 585
R1468 B.n257 B.n256 585
R1469 B.n258 B.n153 585
R1470 B.n260 B.n259 585
R1471 B.n261 B.n152 585
R1472 B.n263 B.n262 585
R1473 B.n264 B.n151 585
R1474 B.n266 B.n265 585
R1475 B.n267 B.n150 585
R1476 B.n269 B.n268 585
R1477 B.n270 B.n149 585
R1478 B.n272 B.n271 585
R1479 B.n273 B.n148 585
R1480 B.n275 B.n274 585
R1481 B.n276 B.n147 585
R1482 B.n278 B.n277 585
R1483 B.n279 B.n146 585
R1484 B.n281 B.n280 585
R1485 B.n282 B.n145 585
R1486 B.n284 B.n283 585
R1487 B.n285 B.n144 585
R1488 B.n287 B.n286 585
R1489 B.n288 B.n143 585
R1490 B.n290 B.n289 585
R1491 B.n291 B.n142 585
R1492 B.n293 B.n292 585
R1493 B.n294 B.n141 585
R1494 B.n296 B.n295 585
R1495 B.n298 B.n138 585
R1496 B.n300 B.n299 585
R1497 B.n301 B.n137 585
R1498 B.n303 B.n302 585
R1499 B.n304 B.n136 585
R1500 B.n306 B.n305 585
R1501 B.n307 B.n135 585
R1502 B.n309 B.n308 585
R1503 B.n310 B.n134 585
R1504 B.n312 B.n311 585
R1505 B.n314 B.n313 585
R1506 B.n315 B.n130 585
R1507 B.n317 B.n316 585
R1508 B.n318 B.n129 585
R1509 B.n320 B.n319 585
R1510 B.n321 B.n128 585
R1511 B.n323 B.n322 585
R1512 B.n324 B.n127 585
R1513 B.n326 B.n325 585
R1514 B.n327 B.n126 585
R1515 B.n329 B.n328 585
R1516 B.n330 B.n125 585
R1517 B.n332 B.n331 585
R1518 B.n333 B.n124 585
R1519 B.n335 B.n334 585
R1520 B.n336 B.n123 585
R1521 B.n338 B.n337 585
R1522 B.n339 B.n122 585
R1523 B.n341 B.n340 585
R1524 B.n342 B.n121 585
R1525 B.n344 B.n343 585
R1526 B.n345 B.n120 585
R1527 B.n347 B.n346 585
R1528 B.n348 B.n119 585
R1529 B.n350 B.n349 585
R1530 B.n351 B.n118 585
R1531 B.n353 B.n352 585
R1532 B.n354 B.n117 585
R1533 B.n356 B.n355 585
R1534 B.n357 B.n116 585
R1535 B.n359 B.n358 585
R1536 B.n360 B.n115 585
R1537 B.n362 B.n361 585
R1538 B.n363 B.n114 585
R1539 B.n365 B.n364 585
R1540 B.n366 B.n113 585
R1541 B.n368 B.n367 585
R1542 B.n369 B.n112 585
R1543 B.n371 B.n370 585
R1544 B.n372 B.n111 585
R1545 B.n374 B.n373 585
R1546 B.n375 B.n110 585
R1547 B.n377 B.n376 585
R1548 B.n378 B.n109 585
R1549 B.n380 B.n379 585
R1550 B.n381 B.n108 585
R1551 B.n383 B.n382 585
R1552 B.n384 B.n107 585
R1553 B.n386 B.n385 585
R1554 B.n387 B.n106 585
R1555 B.n389 B.n388 585
R1556 B.n390 B.n105 585
R1557 B.n392 B.n391 585
R1558 B.n393 B.n104 585
R1559 B.n395 B.n394 585
R1560 B.n396 B.n103 585
R1561 B.n398 B.n397 585
R1562 B.n399 B.n102 585
R1563 B.n401 B.n400 585
R1564 B.n402 B.n101 585
R1565 B.n206 B.n205 585
R1566 B.n204 B.n171 585
R1567 B.n203 B.n202 585
R1568 B.n201 B.n172 585
R1569 B.n200 B.n199 585
R1570 B.n198 B.n173 585
R1571 B.n197 B.n196 585
R1572 B.n195 B.n174 585
R1573 B.n194 B.n193 585
R1574 B.n192 B.n175 585
R1575 B.n191 B.n190 585
R1576 B.n189 B.n176 585
R1577 B.n188 B.n187 585
R1578 B.n186 B.n177 585
R1579 B.n185 B.n184 585
R1580 B.n183 B.n178 585
R1581 B.n182 B.n181 585
R1582 B.n180 B.n179 585
R1583 B.n2 B.n0 585
R1584 B.n685 B.n1 585
R1585 B.n684 B.n683 585
R1586 B.n682 B.n3 585
R1587 B.n681 B.n680 585
R1588 B.n679 B.n4 585
R1589 B.n678 B.n677 585
R1590 B.n676 B.n5 585
R1591 B.n675 B.n674 585
R1592 B.n673 B.n6 585
R1593 B.n672 B.n671 585
R1594 B.n670 B.n7 585
R1595 B.n669 B.n668 585
R1596 B.n667 B.n8 585
R1597 B.n666 B.n665 585
R1598 B.n664 B.n9 585
R1599 B.n663 B.n662 585
R1600 B.n661 B.n10 585
R1601 B.n660 B.n659 585
R1602 B.n658 B.n11 585
R1603 B.n687 B.n686 585
R1604 B.n131 B.t8 512.138
R1605 B.n50 B.t10 512.138
R1606 B.n139 B.t5 512.138
R1607 B.n42 B.t1 512.138
R1608 B.n132 B.t7 488.089
R1609 B.n51 B.t11 488.089
R1610 B.n140 B.t4 488.089
R1611 B.n43 B.t2 488.089
R1612 B.n205 B.n170 468.476
R1613 B.n656 B.n11 468.476
R1614 B.n403 B.n402 468.476
R1615 B.n462 B.n461 468.476
R1616 B.n205 B.n204 163.367
R1617 B.n204 B.n203 163.367
R1618 B.n203 B.n172 163.367
R1619 B.n199 B.n172 163.367
R1620 B.n199 B.n198 163.367
R1621 B.n198 B.n197 163.367
R1622 B.n197 B.n174 163.367
R1623 B.n193 B.n174 163.367
R1624 B.n193 B.n192 163.367
R1625 B.n192 B.n191 163.367
R1626 B.n191 B.n176 163.367
R1627 B.n187 B.n176 163.367
R1628 B.n187 B.n186 163.367
R1629 B.n186 B.n185 163.367
R1630 B.n185 B.n178 163.367
R1631 B.n181 B.n178 163.367
R1632 B.n181 B.n180 163.367
R1633 B.n180 B.n2 163.367
R1634 B.n686 B.n2 163.367
R1635 B.n686 B.n685 163.367
R1636 B.n685 B.n684 163.367
R1637 B.n684 B.n3 163.367
R1638 B.n680 B.n3 163.367
R1639 B.n680 B.n679 163.367
R1640 B.n679 B.n678 163.367
R1641 B.n678 B.n5 163.367
R1642 B.n674 B.n5 163.367
R1643 B.n674 B.n673 163.367
R1644 B.n673 B.n672 163.367
R1645 B.n672 B.n7 163.367
R1646 B.n668 B.n7 163.367
R1647 B.n668 B.n667 163.367
R1648 B.n667 B.n666 163.367
R1649 B.n666 B.n9 163.367
R1650 B.n662 B.n9 163.367
R1651 B.n662 B.n661 163.367
R1652 B.n661 B.n660 163.367
R1653 B.n660 B.n11 163.367
R1654 B.n209 B.n170 163.367
R1655 B.n210 B.n209 163.367
R1656 B.n211 B.n210 163.367
R1657 B.n211 B.n168 163.367
R1658 B.n215 B.n168 163.367
R1659 B.n216 B.n215 163.367
R1660 B.n217 B.n216 163.367
R1661 B.n217 B.n166 163.367
R1662 B.n221 B.n166 163.367
R1663 B.n222 B.n221 163.367
R1664 B.n223 B.n222 163.367
R1665 B.n223 B.n164 163.367
R1666 B.n227 B.n164 163.367
R1667 B.n228 B.n227 163.367
R1668 B.n229 B.n228 163.367
R1669 B.n229 B.n162 163.367
R1670 B.n233 B.n162 163.367
R1671 B.n234 B.n233 163.367
R1672 B.n235 B.n234 163.367
R1673 B.n235 B.n160 163.367
R1674 B.n239 B.n160 163.367
R1675 B.n240 B.n239 163.367
R1676 B.n241 B.n240 163.367
R1677 B.n241 B.n158 163.367
R1678 B.n245 B.n158 163.367
R1679 B.n246 B.n245 163.367
R1680 B.n247 B.n246 163.367
R1681 B.n247 B.n156 163.367
R1682 B.n251 B.n156 163.367
R1683 B.n252 B.n251 163.367
R1684 B.n253 B.n252 163.367
R1685 B.n253 B.n154 163.367
R1686 B.n257 B.n154 163.367
R1687 B.n258 B.n257 163.367
R1688 B.n259 B.n258 163.367
R1689 B.n259 B.n152 163.367
R1690 B.n263 B.n152 163.367
R1691 B.n264 B.n263 163.367
R1692 B.n265 B.n264 163.367
R1693 B.n265 B.n150 163.367
R1694 B.n269 B.n150 163.367
R1695 B.n270 B.n269 163.367
R1696 B.n271 B.n270 163.367
R1697 B.n271 B.n148 163.367
R1698 B.n275 B.n148 163.367
R1699 B.n276 B.n275 163.367
R1700 B.n277 B.n276 163.367
R1701 B.n277 B.n146 163.367
R1702 B.n281 B.n146 163.367
R1703 B.n282 B.n281 163.367
R1704 B.n283 B.n282 163.367
R1705 B.n283 B.n144 163.367
R1706 B.n287 B.n144 163.367
R1707 B.n288 B.n287 163.367
R1708 B.n289 B.n288 163.367
R1709 B.n289 B.n142 163.367
R1710 B.n293 B.n142 163.367
R1711 B.n294 B.n293 163.367
R1712 B.n295 B.n294 163.367
R1713 B.n295 B.n138 163.367
R1714 B.n300 B.n138 163.367
R1715 B.n301 B.n300 163.367
R1716 B.n302 B.n301 163.367
R1717 B.n302 B.n136 163.367
R1718 B.n306 B.n136 163.367
R1719 B.n307 B.n306 163.367
R1720 B.n308 B.n307 163.367
R1721 B.n308 B.n134 163.367
R1722 B.n312 B.n134 163.367
R1723 B.n313 B.n312 163.367
R1724 B.n313 B.n130 163.367
R1725 B.n317 B.n130 163.367
R1726 B.n318 B.n317 163.367
R1727 B.n319 B.n318 163.367
R1728 B.n319 B.n128 163.367
R1729 B.n323 B.n128 163.367
R1730 B.n324 B.n323 163.367
R1731 B.n325 B.n324 163.367
R1732 B.n325 B.n126 163.367
R1733 B.n329 B.n126 163.367
R1734 B.n330 B.n329 163.367
R1735 B.n331 B.n330 163.367
R1736 B.n331 B.n124 163.367
R1737 B.n335 B.n124 163.367
R1738 B.n336 B.n335 163.367
R1739 B.n337 B.n336 163.367
R1740 B.n337 B.n122 163.367
R1741 B.n341 B.n122 163.367
R1742 B.n342 B.n341 163.367
R1743 B.n343 B.n342 163.367
R1744 B.n343 B.n120 163.367
R1745 B.n347 B.n120 163.367
R1746 B.n348 B.n347 163.367
R1747 B.n349 B.n348 163.367
R1748 B.n349 B.n118 163.367
R1749 B.n353 B.n118 163.367
R1750 B.n354 B.n353 163.367
R1751 B.n355 B.n354 163.367
R1752 B.n355 B.n116 163.367
R1753 B.n359 B.n116 163.367
R1754 B.n360 B.n359 163.367
R1755 B.n361 B.n360 163.367
R1756 B.n361 B.n114 163.367
R1757 B.n365 B.n114 163.367
R1758 B.n366 B.n365 163.367
R1759 B.n367 B.n366 163.367
R1760 B.n367 B.n112 163.367
R1761 B.n371 B.n112 163.367
R1762 B.n372 B.n371 163.367
R1763 B.n373 B.n372 163.367
R1764 B.n373 B.n110 163.367
R1765 B.n377 B.n110 163.367
R1766 B.n378 B.n377 163.367
R1767 B.n379 B.n378 163.367
R1768 B.n379 B.n108 163.367
R1769 B.n383 B.n108 163.367
R1770 B.n384 B.n383 163.367
R1771 B.n385 B.n384 163.367
R1772 B.n385 B.n106 163.367
R1773 B.n389 B.n106 163.367
R1774 B.n390 B.n389 163.367
R1775 B.n391 B.n390 163.367
R1776 B.n391 B.n104 163.367
R1777 B.n395 B.n104 163.367
R1778 B.n396 B.n395 163.367
R1779 B.n397 B.n396 163.367
R1780 B.n397 B.n102 163.367
R1781 B.n401 B.n102 163.367
R1782 B.n402 B.n401 163.367
R1783 B.n403 B.n100 163.367
R1784 B.n407 B.n100 163.367
R1785 B.n408 B.n407 163.367
R1786 B.n409 B.n408 163.367
R1787 B.n409 B.n98 163.367
R1788 B.n413 B.n98 163.367
R1789 B.n414 B.n413 163.367
R1790 B.n415 B.n414 163.367
R1791 B.n415 B.n96 163.367
R1792 B.n419 B.n96 163.367
R1793 B.n420 B.n419 163.367
R1794 B.n421 B.n420 163.367
R1795 B.n421 B.n94 163.367
R1796 B.n425 B.n94 163.367
R1797 B.n426 B.n425 163.367
R1798 B.n427 B.n426 163.367
R1799 B.n427 B.n92 163.367
R1800 B.n431 B.n92 163.367
R1801 B.n432 B.n431 163.367
R1802 B.n433 B.n432 163.367
R1803 B.n433 B.n90 163.367
R1804 B.n437 B.n90 163.367
R1805 B.n438 B.n437 163.367
R1806 B.n439 B.n438 163.367
R1807 B.n439 B.n88 163.367
R1808 B.n443 B.n88 163.367
R1809 B.n444 B.n443 163.367
R1810 B.n445 B.n444 163.367
R1811 B.n445 B.n86 163.367
R1812 B.n449 B.n86 163.367
R1813 B.n450 B.n449 163.367
R1814 B.n451 B.n450 163.367
R1815 B.n451 B.n84 163.367
R1816 B.n455 B.n84 163.367
R1817 B.n456 B.n455 163.367
R1818 B.n457 B.n456 163.367
R1819 B.n457 B.n82 163.367
R1820 B.n461 B.n82 163.367
R1821 B.n656 B.n655 163.367
R1822 B.n655 B.n654 163.367
R1823 B.n654 B.n13 163.367
R1824 B.n650 B.n13 163.367
R1825 B.n650 B.n649 163.367
R1826 B.n649 B.n648 163.367
R1827 B.n648 B.n15 163.367
R1828 B.n644 B.n15 163.367
R1829 B.n644 B.n643 163.367
R1830 B.n643 B.n642 163.367
R1831 B.n642 B.n17 163.367
R1832 B.n638 B.n17 163.367
R1833 B.n638 B.n637 163.367
R1834 B.n637 B.n636 163.367
R1835 B.n636 B.n19 163.367
R1836 B.n632 B.n19 163.367
R1837 B.n632 B.n631 163.367
R1838 B.n631 B.n630 163.367
R1839 B.n630 B.n21 163.367
R1840 B.n626 B.n21 163.367
R1841 B.n626 B.n625 163.367
R1842 B.n625 B.n624 163.367
R1843 B.n624 B.n23 163.367
R1844 B.n620 B.n23 163.367
R1845 B.n620 B.n619 163.367
R1846 B.n619 B.n618 163.367
R1847 B.n618 B.n25 163.367
R1848 B.n614 B.n25 163.367
R1849 B.n614 B.n613 163.367
R1850 B.n613 B.n612 163.367
R1851 B.n612 B.n27 163.367
R1852 B.n608 B.n27 163.367
R1853 B.n608 B.n607 163.367
R1854 B.n607 B.n606 163.367
R1855 B.n606 B.n29 163.367
R1856 B.n602 B.n29 163.367
R1857 B.n602 B.n601 163.367
R1858 B.n601 B.n600 163.367
R1859 B.n600 B.n31 163.367
R1860 B.n596 B.n31 163.367
R1861 B.n596 B.n595 163.367
R1862 B.n595 B.n594 163.367
R1863 B.n594 B.n33 163.367
R1864 B.n590 B.n33 163.367
R1865 B.n590 B.n589 163.367
R1866 B.n589 B.n588 163.367
R1867 B.n588 B.n35 163.367
R1868 B.n584 B.n35 163.367
R1869 B.n584 B.n583 163.367
R1870 B.n583 B.n582 163.367
R1871 B.n582 B.n37 163.367
R1872 B.n578 B.n37 163.367
R1873 B.n578 B.n577 163.367
R1874 B.n577 B.n576 163.367
R1875 B.n576 B.n39 163.367
R1876 B.n572 B.n39 163.367
R1877 B.n572 B.n571 163.367
R1878 B.n571 B.n570 163.367
R1879 B.n570 B.n41 163.367
R1880 B.n565 B.n41 163.367
R1881 B.n565 B.n564 163.367
R1882 B.n564 B.n563 163.367
R1883 B.n563 B.n45 163.367
R1884 B.n559 B.n45 163.367
R1885 B.n559 B.n558 163.367
R1886 B.n558 B.n557 163.367
R1887 B.n557 B.n47 163.367
R1888 B.n553 B.n47 163.367
R1889 B.n553 B.n552 163.367
R1890 B.n552 B.n551 163.367
R1891 B.n551 B.n49 163.367
R1892 B.n547 B.n49 163.367
R1893 B.n547 B.n546 163.367
R1894 B.n546 B.n545 163.367
R1895 B.n545 B.n54 163.367
R1896 B.n541 B.n54 163.367
R1897 B.n541 B.n540 163.367
R1898 B.n540 B.n539 163.367
R1899 B.n539 B.n56 163.367
R1900 B.n535 B.n56 163.367
R1901 B.n535 B.n534 163.367
R1902 B.n534 B.n533 163.367
R1903 B.n533 B.n58 163.367
R1904 B.n529 B.n58 163.367
R1905 B.n529 B.n528 163.367
R1906 B.n528 B.n527 163.367
R1907 B.n527 B.n60 163.367
R1908 B.n523 B.n60 163.367
R1909 B.n523 B.n522 163.367
R1910 B.n522 B.n521 163.367
R1911 B.n521 B.n62 163.367
R1912 B.n517 B.n62 163.367
R1913 B.n517 B.n516 163.367
R1914 B.n516 B.n515 163.367
R1915 B.n515 B.n64 163.367
R1916 B.n511 B.n64 163.367
R1917 B.n511 B.n510 163.367
R1918 B.n510 B.n509 163.367
R1919 B.n509 B.n66 163.367
R1920 B.n505 B.n66 163.367
R1921 B.n505 B.n504 163.367
R1922 B.n504 B.n503 163.367
R1923 B.n503 B.n68 163.367
R1924 B.n499 B.n68 163.367
R1925 B.n499 B.n498 163.367
R1926 B.n498 B.n497 163.367
R1927 B.n497 B.n70 163.367
R1928 B.n493 B.n70 163.367
R1929 B.n493 B.n492 163.367
R1930 B.n492 B.n491 163.367
R1931 B.n491 B.n72 163.367
R1932 B.n487 B.n72 163.367
R1933 B.n487 B.n486 163.367
R1934 B.n486 B.n485 163.367
R1935 B.n485 B.n74 163.367
R1936 B.n481 B.n74 163.367
R1937 B.n481 B.n480 163.367
R1938 B.n480 B.n479 163.367
R1939 B.n479 B.n76 163.367
R1940 B.n475 B.n76 163.367
R1941 B.n475 B.n474 163.367
R1942 B.n474 B.n473 163.367
R1943 B.n473 B.n78 163.367
R1944 B.n469 B.n78 163.367
R1945 B.n469 B.n468 163.367
R1946 B.n468 B.n467 163.367
R1947 B.n467 B.n80 163.367
R1948 B.n463 B.n80 163.367
R1949 B.n463 B.n462 163.367
R1950 B.n133 B.n132 59.5399
R1951 B.n297 B.n140 59.5399
R1952 B.n567 B.n43 59.5399
R1953 B.n52 B.n51 59.5399
R1954 B.n460 B.n81 30.4395
R1955 B.n658 B.n657 30.4395
R1956 B.n404 B.n101 30.4395
R1957 B.n207 B.n206 30.4395
R1958 B.n132 B.n131 24.049
R1959 B.n140 B.n139 24.049
R1960 B.n43 B.n42 24.049
R1961 B.n51 B.n50 24.049
R1962 B B.n687 18.0485
R1963 B.n657 B.n12 10.6151
R1964 B.n653 B.n12 10.6151
R1965 B.n653 B.n652 10.6151
R1966 B.n652 B.n651 10.6151
R1967 B.n651 B.n14 10.6151
R1968 B.n647 B.n14 10.6151
R1969 B.n647 B.n646 10.6151
R1970 B.n646 B.n645 10.6151
R1971 B.n645 B.n16 10.6151
R1972 B.n641 B.n16 10.6151
R1973 B.n641 B.n640 10.6151
R1974 B.n640 B.n639 10.6151
R1975 B.n639 B.n18 10.6151
R1976 B.n635 B.n18 10.6151
R1977 B.n635 B.n634 10.6151
R1978 B.n634 B.n633 10.6151
R1979 B.n633 B.n20 10.6151
R1980 B.n629 B.n20 10.6151
R1981 B.n629 B.n628 10.6151
R1982 B.n628 B.n627 10.6151
R1983 B.n627 B.n22 10.6151
R1984 B.n623 B.n22 10.6151
R1985 B.n623 B.n622 10.6151
R1986 B.n622 B.n621 10.6151
R1987 B.n621 B.n24 10.6151
R1988 B.n617 B.n24 10.6151
R1989 B.n617 B.n616 10.6151
R1990 B.n616 B.n615 10.6151
R1991 B.n615 B.n26 10.6151
R1992 B.n611 B.n26 10.6151
R1993 B.n611 B.n610 10.6151
R1994 B.n610 B.n609 10.6151
R1995 B.n609 B.n28 10.6151
R1996 B.n605 B.n28 10.6151
R1997 B.n605 B.n604 10.6151
R1998 B.n604 B.n603 10.6151
R1999 B.n603 B.n30 10.6151
R2000 B.n599 B.n30 10.6151
R2001 B.n599 B.n598 10.6151
R2002 B.n598 B.n597 10.6151
R2003 B.n597 B.n32 10.6151
R2004 B.n593 B.n32 10.6151
R2005 B.n593 B.n592 10.6151
R2006 B.n592 B.n591 10.6151
R2007 B.n591 B.n34 10.6151
R2008 B.n587 B.n34 10.6151
R2009 B.n587 B.n586 10.6151
R2010 B.n586 B.n585 10.6151
R2011 B.n585 B.n36 10.6151
R2012 B.n581 B.n36 10.6151
R2013 B.n581 B.n580 10.6151
R2014 B.n580 B.n579 10.6151
R2015 B.n579 B.n38 10.6151
R2016 B.n575 B.n38 10.6151
R2017 B.n575 B.n574 10.6151
R2018 B.n574 B.n573 10.6151
R2019 B.n573 B.n40 10.6151
R2020 B.n569 B.n40 10.6151
R2021 B.n569 B.n568 10.6151
R2022 B.n566 B.n44 10.6151
R2023 B.n562 B.n44 10.6151
R2024 B.n562 B.n561 10.6151
R2025 B.n561 B.n560 10.6151
R2026 B.n560 B.n46 10.6151
R2027 B.n556 B.n46 10.6151
R2028 B.n556 B.n555 10.6151
R2029 B.n555 B.n554 10.6151
R2030 B.n554 B.n48 10.6151
R2031 B.n550 B.n549 10.6151
R2032 B.n549 B.n548 10.6151
R2033 B.n548 B.n53 10.6151
R2034 B.n544 B.n53 10.6151
R2035 B.n544 B.n543 10.6151
R2036 B.n543 B.n542 10.6151
R2037 B.n542 B.n55 10.6151
R2038 B.n538 B.n55 10.6151
R2039 B.n538 B.n537 10.6151
R2040 B.n537 B.n536 10.6151
R2041 B.n536 B.n57 10.6151
R2042 B.n532 B.n57 10.6151
R2043 B.n532 B.n531 10.6151
R2044 B.n531 B.n530 10.6151
R2045 B.n530 B.n59 10.6151
R2046 B.n526 B.n59 10.6151
R2047 B.n526 B.n525 10.6151
R2048 B.n525 B.n524 10.6151
R2049 B.n524 B.n61 10.6151
R2050 B.n520 B.n61 10.6151
R2051 B.n520 B.n519 10.6151
R2052 B.n519 B.n518 10.6151
R2053 B.n518 B.n63 10.6151
R2054 B.n514 B.n63 10.6151
R2055 B.n514 B.n513 10.6151
R2056 B.n513 B.n512 10.6151
R2057 B.n512 B.n65 10.6151
R2058 B.n508 B.n65 10.6151
R2059 B.n508 B.n507 10.6151
R2060 B.n507 B.n506 10.6151
R2061 B.n506 B.n67 10.6151
R2062 B.n502 B.n67 10.6151
R2063 B.n502 B.n501 10.6151
R2064 B.n501 B.n500 10.6151
R2065 B.n500 B.n69 10.6151
R2066 B.n496 B.n69 10.6151
R2067 B.n496 B.n495 10.6151
R2068 B.n495 B.n494 10.6151
R2069 B.n494 B.n71 10.6151
R2070 B.n490 B.n71 10.6151
R2071 B.n490 B.n489 10.6151
R2072 B.n489 B.n488 10.6151
R2073 B.n488 B.n73 10.6151
R2074 B.n484 B.n73 10.6151
R2075 B.n484 B.n483 10.6151
R2076 B.n483 B.n482 10.6151
R2077 B.n482 B.n75 10.6151
R2078 B.n478 B.n75 10.6151
R2079 B.n478 B.n477 10.6151
R2080 B.n477 B.n476 10.6151
R2081 B.n476 B.n77 10.6151
R2082 B.n472 B.n77 10.6151
R2083 B.n472 B.n471 10.6151
R2084 B.n471 B.n470 10.6151
R2085 B.n470 B.n79 10.6151
R2086 B.n466 B.n79 10.6151
R2087 B.n466 B.n465 10.6151
R2088 B.n465 B.n464 10.6151
R2089 B.n464 B.n81 10.6151
R2090 B.n405 B.n404 10.6151
R2091 B.n406 B.n405 10.6151
R2092 B.n406 B.n99 10.6151
R2093 B.n410 B.n99 10.6151
R2094 B.n411 B.n410 10.6151
R2095 B.n412 B.n411 10.6151
R2096 B.n412 B.n97 10.6151
R2097 B.n416 B.n97 10.6151
R2098 B.n417 B.n416 10.6151
R2099 B.n418 B.n417 10.6151
R2100 B.n418 B.n95 10.6151
R2101 B.n422 B.n95 10.6151
R2102 B.n423 B.n422 10.6151
R2103 B.n424 B.n423 10.6151
R2104 B.n424 B.n93 10.6151
R2105 B.n428 B.n93 10.6151
R2106 B.n429 B.n428 10.6151
R2107 B.n430 B.n429 10.6151
R2108 B.n430 B.n91 10.6151
R2109 B.n434 B.n91 10.6151
R2110 B.n435 B.n434 10.6151
R2111 B.n436 B.n435 10.6151
R2112 B.n436 B.n89 10.6151
R2113 B.n440 B.n89 10.6151
R2114 B.n441 B.n440 10.6151
R2115 B.n442 B.n441 10.6151
R2116 B.n442 B.n87 10.6151
R2117 B.n446 B.n87 10.6151
R2118 B.n447 B.n446 10.6151
R2119 B.n448 B.n447 10.6151
R2120 B.n448 B.n85 10.6151
R2121 B.n452 B.n85 10.6151
R2122 B.n453 B.n452 10.6151
R2123 B.n454 B.n453 10.6151
R2124 B.n454 B.n83 10.6151
R2125 B.n458 B.n83 10.6151
R2126 B.n459 B.n458 10.6151
R2127 B.n460 B.n459 10.6151
R2128 B.n208 B.n207 10.6151
R2129 B.n208 B.n169 10.6151
R2130 B.n212 B.n169 10.6151
R2131 B.n213 B.n212 10.6151
R2132 B.n214 B.n213 10.6151
R2133 B.n214 B.n167 10.6151
R2134 B.n218 B.n167 10.6151
R2135 B.n219 B.n218 10.6151
R2136 B.n220 B.n219 10.6151
R2137 B.n220 B.n165 10.6151
R2138 B.n224 B.n165 10.6151
R2139 B.n225 B.n224 10.6151
R2140 B.n226 B.n225 10.6151
R2141 B.n226 B.n163 10.6151
R2142 B.n230 B.n163 10.6151
R2143 B.n231 B.n230 10.6151
R2144 B.n232 B.n231 10.6151
R2145 B.n232 B.n161 10.6151
R2146 B.n236 B.n161 10.6151
R2147 B.n237 B.n236 10.6151
R2148 B.n238 B.n237 10.6151
R2149 B.n238 B.n159 10.6151
R2150 B.n242 B.n159 10.6151
R2151 B.n243 B.n242 10.6151
R2152 B.n244 B.n243 10.6151
R2153 B.n244 B.n157 10.6151
R2154 B.n248 B.n157 10.6151
R2155 B.n249 B.n248 10.6151
R2156 B.n250 B.n249 10.6151
R2157 B.n250 B.n155 10.6151
R2158 B.n254 B.n155 10.6151
R2159 B.n255 B.n254 10.6151
R2160 B.n256 B.n255 10.6151
R2161 B.n256 B.n153 10.6151
R2162 B.n260 B.n153 10.6151
R2163 B.n261 B.n260 10.6151
R2164 B.n262 B.n261 10.6151
R2165 B.n262 B.n151 10.6151
R2166 B.n266 B.n151 10.6151
R2167 B.n267 B.n266 10.6151
R2168 B.n268 B.n267 10.6151
R2169 B.n268 B.n149 10.6151
R2170 B.n272 B.n149 10.6151
R2171 B.n273 B.n272 10.6151
R2172 B.n274 B.n273 10.6151
R2173 B.n274 B.n147 10.6151
R2174 B.n278 B.n147 10.6151
R2175 B.n279 B.n278 10.6151
R2176 B.n280 B.n279 10.6151
R2177 B.n280 B.n145 10.6151
R2178 B.n284 B.n145 10.6151
R2179 B.n285 B.n284 10.6151
R2180 B.n286 B.n285 10.6151
R2181 B.n286 B.n143 10.6151
R2182 B.n290 B.n143 10.6151
R2183 B.n291 B.n290 10.6151
R2184 B.n292 B.n291 10.6151
R2185 B.n292 B.n141 10.6151
R2186 B.n296 B.n141 10.6151
R2187 B.n299 B.n298 10.6151
R2188 B.n299 B.n137 10.6151
R2189 B.n303 B.n137 10.6151
R2190 B.n304 B.n303 10.6151
R2191 B.n305 B.n304 10.6151
R2192 B.n305 B.n135 10.6151
R2193 B.n309 B.n135 10.6151
R2194 B.n310 B.n309 10.6151
R2195 B.n311 B.n310 10.6151
R2196 B.n315 B.n314 10.6151
R2197 B.n316 B.n315 10.6151
R2198 B.n316 B.n129 10.6151
R2199 B.n320 B.n129 10.6151
R2200 B.n321 B.n320 10.6151
R2201 B.n322 B.n321 10.6151
R2202 B.n322 B.n127 10.6151
R2203 B.n326 B.n127 10.6151
R2204 B.n327 B.n326 10.6151
R2205 B.n328 B.n327 10.6151
R2206 B.n328 B.n125 10.6151
R2207 B.n332 B.n125 10.6151
R2208 B.n333 B.n332 10.6151
R2209 B.n334 B.n333 10.6151
R2210 B.n334 B.n123 10.6151
R2211 B.n338 B.n123 10.6151
R2212 B.n339 B.n338 10.6151
R2213 B.n340 B.n339 10.6151
R2214 B.n340 B.n121 10.6151
R2215 B.n344 B.n121 10.6151
R2216 B.n345 B.n344 10.6151
R2217 B.n346 B.n345 10.6151
R2218 B.n346 B.n119 10.6151
R2219 B.n350 B.n119 10.6151
R2220 B.n351 B.n350 10.6151
R2221 B.n352 B.n351 10.6151
R2222 B.n352 B.n117 10.6151
R2223 B.n356 B.n117 10.6151
R2224 B.n357 B.n356 10.6151
R2225 B.n358 B.n357 10.6151
R2226 B.n358 B.n115 10.6151
R2227 B.n362 B.n115 10.6151
R2228 B.n363 B.n362 10.6151
R2229 B.n364 B.n363 10.6151
R2230 B.n364 B.n113 10.6151
R2231 B.n368 B.n113 10.6151
R2232 B.n369 B.n368 10.6151
R2233 B.n370 B.n369 10.6151
R2234 B.n370 B.n111 10.6151
R2235 B.n374 B.n111 10.6151
R2236 B.n375 B.n374 10.6151
R2237 B.n376 B.n375 10.6151
R2238 B.n376 B.n109 10.6151
R2239 B.n380 B.n109 10.6151
R2240 B.n381 B.n380 10.6151
R2241 B.n382 B.n381 10.6151
R2242 B.n382 B.n107 10.6151
R2243 B.n386 B.n107 10.6151
R2244 B.n387 B.n386 10.6151
R2245 B.n388 B.n387 10.6151
R2246 B.n388 B.n105 10.6151
R2247 B.n392 B.n105 10.6151
R2248 B.n393 B.n392 10.6151
R2249 B.n394 B.n393 10.6151
R2250 B.n394 B.n103 10.6151
R2251 B.n398 B.n103 10.6151
R2252 B.n399 B.n398 10.6151
R2253 B.n400 B.n399 10.6151
R2254 B.n400 B.n101 10.6151
R2255 B.n206 B.n171 10.6151
R2256 B.n202 B.n171 10.6151
R2257 B.n202 B.n201 10.6151
R2258 B.n201 B.n200 10.6151
R2259 B.n200 B.n173 10.6151
R2260 B.n196 B.n173 10.6151
R2261 B.n196 B.n195 10.6151
R2262 B.n195 B.n194 10.6151
R2263 B.n194 B.n175 10.6151
R2264 B.n190 B.n175 10.6151
R2265 B.n190 B.n189 10.6151
R2266 B.n189 B.n188 10.6151
R2267 B.n188 B.n177 10.6151
R2268 B.n184 B.n177 10.6151
R2269 B.n184 B.n183 10.6151
R2270 B.n183 B.n182 10.6151
R2271 B.n182 B.n179 10.6151
R2272 B.n179 B.n0 10.6151
R2273 B.n683 B.n1 10.6151
R2274 B.n683 B.n682 10.6151
R2275 B.n682 B.n681 10.6151
R2276 B.n681 B.n4 10.6151
R2277 B.n677 B.n4 10.6151
R2278 B.n677 B.n676 10.6151
R2279 B.n676 B.n675 10.6151
R2280 B.n675 B.n6 10.6151
R2281 B.n671 B.n6 10.6151
R2282 B.n671 B.n670 10.6151
R2283 B.n670 B.n669 10.6151
R2284 B.n669 B.n8 10.6151
R2285 B.n665 B.n8 10.6151
R2286 B.n665 B.n664 10.6151
R2287 B.n664 B.n663 10.6151
R2288 B.n663 B.n10 10.6151
R2289 B.n659 B.n10 10.6151
R2290 B.n659 B.n658 10.6151
R2291 B.n568 B.n567 9.36635
R2292 B.n550 B.n52 9.36635
R2293 B.n297 B.n296 9.36635
R2294 B.n314 B.n133 9.36635
R2295 B.n687 B.n0 2.81026
R2296 B.n687 B.n1 2.81026
R2297 B.n567 B.n566 1.24928
R2298 B.n52 B.n48 1.24928
R2299 B.n298 B.n297 1.24928
R2300 B.n311 B.n133 1.24928
C0 VTAIL B 5.72052f
C1 VP B 1.21337f
C2 VN VDD2 5.21238f
C3 w_n1714_n4616# B 8.91569f
C4 VDD1 B 1.13153f
C5 VTAIL VN 4.60987f
C6 VP VN 6.12965f
C7 VTAIL VDD2 8.677299f
C8 VP VDD2 0.28721f
C9 VN w_n1714_n4616# 2.71218f
C10 VDD2 w_n1714_n4616# 1.29907f
C11 VDD1 VN 0.147915f
C12 VTAIL VP 4.62397f
C13 VDD1 VDD2 0.617301f
C14 VTAIL w_n1714_n4616# 5.63772f
C15 VP w_n1714_n4616# 2.92825f
C16 VTAIL VDD1 8.634429f
C17 VDD1 VP 5.35137f
C18 VN B 0.862677f
C19 VDD2 B 1.15619f
C20 VDD1 w_n1714_n4616# 1.28027f
C21 VDD2 VSUBS 0.854721f
C22 VDD1 VSUBS 5.872586f
C23 VTAIL VSUBS 1.201484f
C24 VN VSUBS 6.01392f
C25 VP VSUBS 1.652454f
C26 B VSUBS 3.327603f
C27 w_n1714_n4616# VSUBS 96.7313f
C28 B.n0 VSUBS 0.004703f
C29 B.n1 VSUBS 0.004703f
C30 B.n2 VSUBS 0.007437f
C31 B.n3 VSUBS 0.007437f
C32 B.n4 VSUBS 0.007437f
C33 B.n5 VSUBS 0.007437f
C34 B.n6 VSUBS 0.007437f
C35 B.n7 VSUBS 0.007437f
C36 B.n8 VSUBS 0.007437f
C37 B.n9 VSUBS 0.007437f
C38 B.n10 VSUBS 0.007437f
C39 B.n11 VSUBS 0.015945f
C40 B.n12 VSUBS 0.007437f
C41 B.n13 VSUBS 0.007437f
C42 B.n14 VSUBS 0.007437f
C43 B.n15 VSUBS 0.007437f
C44 B.n16 VSUBS 0.007437f
C45 B.n17 VSUBS 0.007437f
C46 B.n18 VSUBS 0.007437f
C47 B.n19 VSUBS 0.007437f
C48 B.n20 VSUBS 0.007437f
C49 B.n21 VSUBS 0.007437f
C50 B.n22 VSUBS 0.007437f
C51 B.n23 VSUBS 0.007437f
C52 B.n24 VSUBS 0.007437f
C53 B.n25 VSUBS 0.007437f
C54 B.n26 VSUBS 0.007437f
C55 B.n27 VSUBS 0.007437f
C56 B.n28 VSUBS 0.007437f
C57 B.n29 VSUBS 0.007437f
C58 B.n30 VSUBS 0.007437f
C59 B.n31 VSUBS 0.007437f
C60 B.n32 VSUBS 0.007437f
C61 B.n33 VSUBS 0.007437f
C62 B.n34 VSUBS 0.007437f
C63 B.n35 VSUBS 0.007437f
C64 B.n36 VSUBS 0.007437f
C65 B.n37 VSUBS 0.007437f
C66 B.n38 VSUBS 0.007437f
C67 B.n39 VSUBS 0.007437f
C68 B.n40 VSUBS 0.007437f
C69 B.n41 VSUBS 0.007437f
C70 B.t2 VSUBS 0.379227f
C71 B.t1 VSUBS 0.394918f
C72 B.t0 VSUBS 0.722159f
C73 B.n42 VSUBS 0.498528f
C74 B.n43 VSUBS 0.344759f
C75 B.n44 VSUBS 0.007437f
C76 B.n45 VSUBS 0.007437f
C77 B.n46 VSUBS 0.007437f
C78 B.n47 VSUBS 0.007437f
C79 B.n48 VSUBS 0.004156f
C80 B.n49 VSUBS 0.007437f
C81 B.t11 VSUBS 0.379231f
C82 B.t10 VSUBS 0.394921f
C83 B.t9 VSUBS 0.722159f
C84 B.n50 VSUBS 0.498524f
C85 B.n51 VSUBS 0.344755f
C86 B.n52 VSUBS 0.01723f
C87 B.n53 VSUBS 0.007437f
C88 B.n54 VSUBS 0.007437f
C89 B.n55 VSUBS 0.007437f
C90 B.n56 VSUBS 0.007437f
C91 B.n57 VSUBS 0.007437f
C92 B.n58 VSUBS 0.007437f
C93 B.n59 VSUBS 0.007437f
C94 B.n60 VSUBS 0.007437f
C95 B.n61 VSUBS 0.007437f
C96 B.n62 VSUBS 0.007437f
C97 B.n63 VSUBS 0.007437f
C98 B.n64 VSUBS 0.007437f
C99 B.n65 VSUBS 0.007437f
C100 B.n66 VSUBS 0.007437f
C101 B.n67 VSUBS 0.007437f
C102 B.n68 VSUBS 0.007437f
C103 B.n69 VSUBS 0.007437f
C104 B.n70 VSUBS 0.007437f
C105 B.n71 VSUBS 0.007437f
C106 B.n72 VSUBS 0.007437f
C107 B.n73 VSUBS 0.007437f
C108 B.n74 VSUBS 0.007437f
C109 B.n75 VSUBS 0.007437f
C110 B.n76 VSUBS 0.007437f
C111 B.n77 VSUBS 0.007437f
C112 B.n78 VSUBS 0.007437f
C113 B.n79 VSUBS 0.007437f
C114 B.n80 VSUBS 0.007437f
C115 B.n81 VSUBS 0.016359f
C116 B.n82 VSUBS 0.007437f
C117 B.n83 VSUBS 0.007437f
C118 B.n84 VSUBS 0.007437f
C119 B.n85 VSUBS 0.007437f
C120 B.n86 VSUBS 0.007437f
C121 B.n87 VSUBS 0.007437f
C122 B.n88 VSUBS 0.007437f
C123 B.n89 VSUBS 0.007437f
C124 B.n90 VSUBS 0.007437f
C125 B.n91 VSUBS 0.007437f
C126 B.n92 VSUBS 0.007437f
C127 B.n93 VSUBS 0.007437f
C128 B.n94 VSUBS 0.007437f
C129 B.n95 VSUBS 0.007437f
C130 B.n96 VSUBS 0.007437f
C131 B.n97 VSUBS 0.007437f
C132 B.n98 VSUBS 0.007437f
C133 B.n99 VSUBS 0.007437f
C134 B.n100 VSUBS 0.007437f
C135 B.n101 VSUBS 0.017302f
C136 B.n102 VSUBS 0.007437f
C137 B.n103 VSUBS 0.007437f
C138 B.n104 VSUBS 0.007437f
C139 B.n105 VSUBS 0.007437f
C140 B.n106 VSUBS 0.007437f
C141 B.n107 VSUBS 0.007437f
C142 B.n108 VSUBS 0.007437f
C143 B.n109 VSUBS 0.007437f
C144 B.n110 VSUBS 0.007437f
C145 B.n111 VSUBS 0.007437f
C146 B.n112 VSUBS 0.007437f
C147 B.n113 VSUBS 0.007437f
C148 B.n114 VSUBS 0.007437f
C149 B.n115 VSUBS 0.007437f
C150 B.n116 VSUBS 0.007437f
C151 B.n117 VSUBS 0.007437f
C152 B.n118 VSUBS 0.007437f
C153 B.n119 VSUBS 0.007437f
C154 B.n120 VSUBS 0.007437f
C155 B.n121 VSUBS 0.007437f
C156 B.n122 VSUBS 0.007437f
C157 B.n123 VSUBS 0.007437f
C158 B.n124 VSUBS 0.007437f
C159 B.n125 VSUBS 0.007437f
C160 B.n126 VSUBS 0.007437f
C161 B.n127 VSUBS 0.007437f
C162 B.n128 VSUBS 0.007437f
C163 B.n129 VSUBS 0.007437f
C164 B.n130 VSUBS 0.007437f
C165 B.t7 VSUBS 0.379231f
C166 B.t8 VSUBS 0.394921f
C167 B.t6 VSUBS 0.722159f
C168 B.n131 VSUBS 0.498524f
C169 B.n132 VSUBS 0.344755f
C170 B.n133 VSUBS 0.01723f
C171 B.n134 VSUBS 0.007437f
C172 B.n135 VSUBS 0.007437f
C173 B.n136 VSUBS 0.007437f
C174 B.n137 VSUBS 0.007437f
C175 B.n138 VSUBS 0.007437f
C176 B.t4 VSUBS 0.379227f
C177 B.t5 VSUBS 0.394918f
C178 B.t3 VSUBS 0.722159f
C179 B.n139 VSUBS 0.498528f
C180 B.n140 VSUBS 0.344759f
C181 B.n141 VSUBS 0.007437f
C182 B.n142 VSUBS 0.007437f
C183 B.n143 VSUBS 0.007437f
C184 B.n144 VSUBS 0.007437f
C185 B.n145 VSUBS 0.007437f
C186 B.n146 VSUBS 0.007437f
C187 B.n147 VSUBS 0.007437f
C188 B.n148 VSUBS 0.007437f
C189 B.n149 VSUBS 0.007437f
C190 B.n150 VSUBS 0.007437f
C191 B.n151 VSUBS 0.007437f
C192 B.n152 VSUBS 0.007437f
C193 B.n153 VSUBS 0.007437f
C194 B.n154 VSUBS 0.007437f
C195 B.n155 VSUBS 0.007437f
C196 B.n156 VSUBS 0.007437f
C197 B.n157 VSUBS 0.007437f
C198 B.n158 VSUBS 0.007437f
C199 B.n159 VSUBS 0.007437f
C200 B.n160 VSUBS 0.007437f
C201 B.n161 VSUBS 0.007437f
C202 B.n162 VSUBS 0.007437f
C203 B.n163 VSUBS 0.007437f
C204 B.n164 VSUBS 0.007437f
C205 B.n165 VSUBS 0.007437f
C206 B.n166 VSUBS 0.007437f
C207 B.n167 VSUBS 0.007437f
C208 B.n168 VSUBS 0.007437f
C209 B.n169 VSUBS 0.007437f
C210 B.n170 VSUBS 0.017302f
C211 B.n171 VSUBS 0.007437f
C212 B.n172 VSUBS 0.007437f
C213 B.n173 VSUBS 0.007437f
C214 B.n174 VSUBS 0.007437f
C215 B.n175 VSUBS 0.007437f
C216 B.n176 VSUBS 0.007437f
C217 B.n177 VSUBS 0.007437f
C218 B.n178 VSUBS 0.007437f
C219 B.n179 VSUBS 0.007437f
C220 B.n180 VSUBS 0.007437f
C221 B.n181 VSUBS 0.007437f
C222 B.n182 VSUBS 0.007437f
C223 B.n183 VSUBS 0.007437f
C224 B.n184 VSUBS 0.007437f
C225 B.n185 VSUBS 0.007437f
C226 B.n186 VSUBS 0.007437f
C227 B.n187 VSUBS 0.007437f
C228 B.n188 VSUBS 0.007437f
C229 B.n189 VSUBS 0.007437f
C230 B.n190 VSUBS 0.007437f
C231 B.n191 VSUBS 0.007437f
C232 B.n192 VSUBS 0.007437f
C233 B.n193 VSUBS 0.007437f
C234 B.n194 VSUBS 0.007437f
C235 B.n195 VSUBS 0.007437f
C236 B.n196 VSUBS 0.007437f
C237 B.n197 VSUBS 0.007437f
C238 B.n198 VSUBS 0.007437f
C239 B.n199 VSUBS 0.007437f
C240 B.n200 VSUBS 0.007437f
C241 B.n201 VSUBS 0.007437f
C242 B.n202 VSUBS 0.007437f
C243 B.n203 VSUBS 0.007437f
C244 B.n204 VSUBS 0.007437f
C245 B.n205 VSUBS 0.015945f
C246 B.n206 VSUBS 0.015945f
C247 B.n207 VSUBS 0.017302f
C248 B.n208 VSUBS 0.007437f
C249 B.n209 VSUBS 0.007437f
C250 B.n210 VSUBS 0.007437f
C251 B.n211 VSUBS 0.007437f
C252 B.n212 VSUBS 0.007437f
C253 B.n213 VSUBS 0.007437f
C254 B.n214 VSUBS 0.007437f
C255 B.n215 VSUBS 0.007437f
C256 B.n216 VSUBS 0.007437f
C257 B.n217 VSUBS 0.007437f
C258 B.n218 VSUBS 0.007437f
C259 B.n219 VSUBS 0.007437f
C260 B.n220 VSUBS 0.007437f
C261 B.n221 VSUBS 0.007437f
C262 B.n222 VSUBS 0.007437f
C263 B.n223 VSUBS 0.007437f
C264 B.n224 VSUBS 0.007437f
C265 B.n225 VSUBS 0.007437f
C266 B.n226 VSUBS 0.007437f
C267 B.n227 VSUBS 0.007437f
C268 B.n228 VSUBS 0.007437f
C269 B.n229 VSUBS 0.007437f
C270 B.n230 VSUBS 0.007437f
C271 B.n231 VSUBS 0.007437f
C272 B.n232 VSUBS 0.007437f
C273 B.n233 VSUBS 0.007437f
C274 B.n234 VSUBS 0.007437f
C275 B.n235 VSUBS 0.007437f
C276 B.n236 VSUBS 0.007437f
C277 B.n237 VSUBS 0.007437f
C278 B.n238 VSUBS 0.007437f
C279 B.n239 VSUBS 0.007437f
C280 B.n240 VSUBS 0.007437f
C281 B.n241 VSUBS 0.007437f
C282 B.n242 VSUBS 0.007437f
C283 B.n243 VSUBS 0.007437f
C284 B.n244 VSUBS 0.007437f
C285 B.n245 VSUBS 0.007437f
C286 B.n246 VSUBS 0.007437f
C287 B.n247 VSUBS 0.007437f
C288 B.n248 VSUBS 0.007437f
C289 B.n249 VSUBS 0.007437f
C290 B.n250 VSUBS 0.007437f
C291 B.n251 VSUBS 0.007437f
C292 B.n252 VSUBS 0.007437f
C293 B.n253 VSUBS 0.007437f
C294 B.n254 VSUBS 0.007437f
C295 B.n255 VSUBS 0.007437f
C296 B.n256 VSUBS 0.007437f
C297 B.n257 VSUBS 0.007437f
C298 B.n258 VSUBS 0.007437f
C299 B.n259 VSUBS 0.007437f
C300 B.n260 VSUBS 0.007437f
C301 B.n261 VSUBS 0.007437f
C302 B.n262 VSUBS 0.007437f
C303 B.n263 VSUBS 0.007437f
C304 B.n264 VSUBS 0.007437f
C305 B.n265 VSUBS 0.007437f
C306 B.n266 VSUBS 0.007437f
C307 B.n267 VSUBS 0.007437f
C308 B.n268 VSUBS 0.007437f
C309 B.n269 VSUBS 0.007437f
C310 B.n270 VSUBS 0.007437f
C311 B.n271 VSUBS 0.007437f
C312 B.n272 VSUBS 0.007437f
C313 B.n273 VSUBS 0.007437f
C314 B.n274 VSUBS 0.007437f
C315 B.n275 VSUBS 0.007437f
C316 B.n276 VSUBS 0.007437f
C317 B.n277 VSUBS 0.007437f
C318 B.n278 VSUBS 0.007437f
C319 B.n279 VSUBS 0.007437f
C320 B.n280 VSUBS 0.007437f
C321 B.n281 VSUBS 0.007437f
C322 B.n282 VSUBS 0.007437f
C323 B.n283 VSUBS 0.007437f
C324 B.n284 VSUBS 0.007437f
C325 B.n285 VSUBS 0.007437f
C326 B.n286 VSUBS 0.007437f
C327 B.n287 VSUBS 0.007437f
C328 B.n288 VSUBS 0.007437f
C329 B.n289 VSUBS 0.007437f
C330 B.n290 VSUBS 0.007437f
C331 B.n291 VSUBS 0.007437f
C332 B.n292 VSUBS 0.007437f
C333 B.n293 VSUBS 0.007437f
C334 B.n294 VSUBS 0.007437f
C335 B.n295 VSUBS 0.007437f
C336 B.n296 VSUBS 0.006999f
C337 B.n297 VSUBS 0.01723f
C338 B.n298 VSUBS 0.004156f
C339 B.n299 VSUBS 0.007437f
C340 B.n300 VSUBS 0.007437f
C341 B.n301 VSUBS 0.007437f
C342 B.n302 VSUBS 0.007437f
C343 B.n303 VSUBS 0.007437f
C344 B.n304 VSUBS 0.007437f
C345 B.n305 VSUBS 0.007437f
C346 B.n306 VSUBS 0.007437f
C347 B.n307 VSUBS 0.007437f
C348 B.n308 VSUBS 0.007437f
C349 B.n309 VSUBS 0.007437f
C350 B.n310 VSUBS 0.007437f
C351 B.n311 VSUBS 0.004156f
C352 B.n312 VSUBS 0.007437f
C353 B.n313 VSUBS 0.007437f
C354 B.n314 VSUBS 0.006999f
C355 B.n315 VSUBS 0.007437f
C356 B.n316 VSUBS 0.007437f
C357 B.n317 VSUBS 0.007437f
C358 B.n318 VSUBS 0.007437f
C359 B.n319 VSUBS 0.007437f
C360 B.n320 VSUBS 0.007437f
C361 B.n321 VSUBS 0.007437f
C362 B.n322 VSUBS 0.007437f
C363 B.n323 VSUBS 0.007437f
C364 B.n324 VSUBS 0.007437f
C365 B.n325 VSUBS 0.007437f
C366 B.n326 VSUBS 0.007437f
C367 B.n327 VSUBS 0.007437f
C368 B.n328 VSUBS 0.007437f
C369 B.n329 VSUBS 0.007437f
C370 B.n330 VSUBS 0.007437f
C371 B.n331 VSUBS 0.007437f
C372 B.n332 VSUBS 0.007437f
C373 B.n333 VSUBS 0.007437f
C374 B.n334 VSUBS 0.007437f
C375 B.n335 VSUBS 0.007437f
C376 B.n336 VSUBS 0.007437f
C377 B.n337 VSUBS 0.007437f
C378 B.n338 VSUBS 0.007437f
C379 B.n339 VSUBS 0.007437f
C380 B.n340 VSUBS 0.007437f
C381 B.n341 VSUBS 0.007437f
C382 B.n342 VSUBS 0.007437f
C383 B.n343 VSUBS 0.007437f
C384 B.n344 VSUBS 0.007437f
C385 B.n345 VSUBS 0.007437f
C386 B.n346 VSUBS 0.007437f
C387 B.n347 VSUBS 0.007437f
C388 B.n348 VSUBS 0.007437f
C389 B.n349 VSUBS 0.007437f
C390 B.n350 VSUBS 0.007437f
C391 B.n351 VSUBS 0.007437f
C392 B.n352 VSUBS 0.007437f
C393 B.n353 VSUBS 0.007437f
C394 B.n354 VSUBS 0.007437f
C395 B.n355 VSUBS 0.007437f
C396 B.n356 VSUBS 0.007437f
C397 B.n357 VSUBS 0.007437f
C398 B.n358 VSUBS 0.007437f
C399 B.n359 VSUBS 0.007437f
C400 B.n360 VSUBS 0.007437f
C401 B.n361 VSUBS 0.007437f
C402 B.n362 VSUBS 0.007437f
C403 B.n363 VSUBS 0.007437f
C404 B.n364 VSUBS 0.007437f
C405 B.n365 VSUBS 0.007437f
C406 B.n366 VSUBS 0.007437f
C407 B.n367 VSUBS 0.007437f
C408 B.n368 VSUBS 0.007437f
C409 B.n369 VSUBS 0.007437f
C410 B.n370 VSUBS 0.007437f
C411 B.n371 VSUBS 0.007437f
C412 B.n372 VSUBS 0.007437f
C413 B.n373 VSUBS 0.007437f
C414 B.n374 VSUBS 0.007437f
C415 B.n375 VSUBS 0.007437f
C416 B.n376 VSUBS 0.007437f
C417 B.n377 VSUBS 0.007437f
C418 B.n378 VSUBS 0.007437f
C419 B.n379 VSUBS 0.007437f
C420 B.n380 VSUBS 0.007437f
C421 B.n381 VSUBS 0.007437f
C422 B.n382 VSUBS 0.007437f
C423 B.n383 VSUBS 0.007437f
C424 B.n384 VSUBS 0.007437f
C425 B.n385 VSUBS 0.007437f
C426 B.n386 VSUBS 0.007437f
C427 B.n387 VSUBS 0.007437f
C428 B.n388 VSUBS 0.007437f
C429 B.n389 VSUBS 0.007437f
C430 B.n390 VSUBS 0.007437f
C431 B.n391 VSUBS 0.007437f
C432 B.n392 VSUBS 0.007437f
C433 B.n393 VSUBS 0.007437f
C434 B.n394 VSUBS 0.007437f
C435 B.n395 VSUBS 0.007437f
C436 B.n396 VSUBS 0.007437f
C437 B.n397 VSUBS 0.007437f
C438 B.n398 VSUBS 0.007437f
C439 B.n399 VSUBS 0.007437f
C440 B.n400 VSUBS 0.007437f
C441 B.n401 VSUBS 0.007437f
C442 B.n402 VSUBS 0.017302f
C443 B.n403 VSUBS 0.015945f
C444 B.n404 VSUBS 0.015945f
C445 B.n405 VSUBS 0.007437f
C446 B.n406 VSUBS 0.007437f
C447 B.n407 VSUBS 0.007437f
C448 B.n408 VSUBS 0.007437f
C449 B.n409 VSUBS 0.007437f
C450 B.n410 VSUBS 0.007437f
C451 B.n411 VSUBS 0.007437f
C452 B.n412 VSUBS 0.007437f
C453 B.n413 VSUBS 0.007437f
C454 B.n414 VSUBS 0.007437f
C455 B.n415 VSUBS 0.007437f
C456 B.n416 VSUBS 0.007437f
C457 B.n417 VSUBS 0.007437f
C458 B.n418 VSUBS 0.007437f
C459 B.n419 VSUBS 0.007437f
C460 B.n420 VSUBS 0.007437f
C461 B.n421 VSUBS 0.007437f
C462 B.n422 VSUBS 0.007437f
C463 B.n423 VSUBS 0.007437f
C464 B.n424 VSUBS 0.007437f
C465 B.n425 VSUBS 0.007437f
C466 B.n426 VSUBS 0.007437f
C467 B.n427 VSUBS 0.007437f
C468 B.n428 VSUBS 0.007437f
C469 B.n429 VSUBS 0.007437f
C470 B.n430 VSUBS 0.007437f
C471 B.n431 VSUBS 0.007437f
C472 B.n432 VSUBS 0.007437f
C473 B.n433 VSUBS 0.007437f
C474 B.n434 VSUBS 0.007437f
C475 B.n435 VSUBS 0.007437f
C476 B.n436 VSUBS 0.007437f
C477 B.n437 VSUBS 0.007437f
C478 B.n438 VSUBS 0.007437f
C479 B.n439 VSUBS 0.007437f
C480 B.n440 VSUBS 0.007437f
C481 B.n441 VSUBS 0.007437f
C482 B.n442 VSUBS 0.007437f
C483 B.n443 VSUBS 0.007437f
C484 B.n444 VSUBS 0.007437f
C485 B.n445 VSUBS 0.007437f
C486 B.n446 VSUBS 0.007437f
C487 B.n447 VSUBS 0.007437f
C488 B.n448 VSUBS 0.007437f
C489 B.n449 VSUBS 0.007437f
C490 B.n450 VSUBS 0.007437f
C491 B.n451 VSUBS 0.007437f
C492 B.n452 VSUBS 0.007437f
C493 B.n453 VSUBS 0.007437f
C494 B.n454 VSUBS 0.007437f
C495 B.n455 VSUBS 0.007437f
C496 B.n456 VSUBS 0.007437f
C497 B.n457 VSUBS 0.007437f
C498 B.n458 VSUBS 0.007437f
C499 B.n459 VSUBS 0.007437f
C500 B.n460 VSUBS 0.016888f
C501 B.n461 VSUBS 0.015945f
C502 B.n462 VSUBS 0.017302f
C503 B.n463 VSUBS 0.007437f
C504 B.n464 VSUBS 0.007437f
C505 B.n465 VSUBS 0.007437f
C506 B.n466 VSUBS 0.007437f
C507 B.n467 VSUBS 0.007437f
C508 B.n468 VSUBS 0.007437f
C509 B.n469 VSUBS 0.007437f
C510 B.n470 VSUBS 0.007437f
C511 B.n471 VSUBS 0.007437f
C512 B.n472 VSUBS 0.007437f
C513 B.n473 VSUBS 0.007437f
C514 B.n474 VSUBS 0.007437f
C515 B.n475 VSUBS 0.007437f
C516 B.n476 VSUBS 0.007437f
C517 B.n477 VSUBS 0.007437f
C518 B.n478 VSUBS 0.007437f
C519 B.n479 VSUBS 0.007437f
C520 B.n480 VSUBS 0.007437f
C521 B.n481 VSUBS 0.007437f
C522 B.n482 VSUBS 0.007437f
C523 B.n483 VSUBS 0.007437f
C524 B.n484 VSUBS 0.007437f
C525 B.n485 VSUBS 0.007437f
C526 B.n486 VSUBS 0.007437f
C527 B.n487 VSUBS 0.007437f
C528 B.n488 VSUBS 0.007437f
C529 B.n489 VSUBS 0.007437f
C530 B.n490 VSUBS 0.007437f
C531 B.n491 VSUBS 0.007437f
C532 B.n492 VSUBS 0.007437f
C533 B.n493 VSUBS 0.007437f
C534 B.n494 VSUBS 0.007437f
C535 B.n495 VSUBS 0.007437f
C536 B.n496 VSUBS 0.007437f
C537 B.n497 VSUBS 0.007437f
C538 B.n498 VSUBS 0.007437f
C539 B.n499 VSUBS 0.007437f
C540 B.n500 VSUBS 0.007437f
C541 B.n501 VSUBS 0.007437f
C542 B.n502 VSUBS 0.007437f
C543 B.n503 VSUBS 0.007437f
C544 B.n504 VSUBS 0.007437f
C545 B.n505 VSUBS 0.007437f
C546 B.n506 VSUBS 0.007437f
C547 B.n507 VSUBS 0.007437f
C548 B.n508 VSUBS 0.007437f
C549 B.n509 VSUBS 0.007437f
C550 B.n510 VSUBS 0.007437f
C551 B.n511 VSUBS 0.007437f
C552 B.n512 VSUBS 0.007437f
C553 B.n513 VSUBS 0.007437f
C554 B.n514 VSUBS 0.007437f
C555 B.n515 VSUBS 0.007437f
C556 B.n516 VSUBS 0.007437f
C557 B.n517 VSUBS 0.007437f
C558 B.n518 VSUBS 0.007437f
C559 B.n519 VSUBS 0.007437f
C560 B.n520 VSUBS 0.007437f
C561 B.n521 VSUBS 0.007437f
C562 B.n522 VSUBS 0.007437f
C563 B.n523 VSUBS 0.007437f
C564 B.n524 VSUBS 0.007437f
C565 B.n525 VSUBS 0.007437f
C566 B.n526 VSUBS 0.007437f
C567 B.n527 VSUBS 0.007437f
C568 B.n528 VSUBS 0.007437f
C569 B.n529 VSUBS 0.007437f
C570 B.n530 VSUBS 0.007437f
C571 B.n531 VSUBS 0.007437f
C572 B.n532 VSUBS 0.007437f
C573 B.n533 VSUBS 0.007437f
C574 B.n534 VSUBS 0.007437f
C575 B.n535 VSUBS 0.007437f
C576 B.n536 VSUBS 0.007437f
C577 B.n537 VSUBS 0.007437f
C578 B.n538 VSUBS 0.007437f
C579 B.n539 VSUBS 0.007437f
C580 B.n540 VSUBS 0.007437f
C581 B.n541 VSUBS 0.007437f
C582 B.n542 VSUBS 0.007437f
C583 B.n543 VSUBS 0.007437f
C584 B.n544 VSUBS 0.007437f
C585 B.n545 VSUBS 0.007437f
C586 B.n546 VSUBS 0.007437f
C587 B.n547 VSUBS 0.007437f
C588 B.n548 VSUBS 0.007437f
C589 B.n549 VSUBS 0.007437f
C590 B.n550 VSUBS 0.006999f
C591 B.n551 VSUBS 0.007437f
C592 B.n552 VSUBS 0.007437f
C593 B.n553 VSUBS 0.007437f
C594 B.n554 VSUBS 0.007437f
C595 B.n555 VSUBS 0.007437f
C596 B.n556 VSUBS 0.007437f
C597 B.n557 VSUBS 0.007437f
C598 B.n558 VSUBS 0.007437f
C599 B.n559 VSUBS 0.007437f
C600 B.n560 VSUBS 0.007437f
C601 B.n561 VSUBS 0.007437f
C602 B.n562 VSUBS 0.007437f
C603 B.n563 VSUBS 0.007437f
C604 B.n564 VSUBS 0.007437f
C605 B.n565 VSUBS 0.007437f
C606 B.n566 VSUBS 0.004156f
C607 B.n567 VSUBS 0.01723f
C608 B.n568 VSUBS 0.006999f
C609 B.n569 VSUBS 0.007437f
C610 B.n570 VSUBS 0.007437f
C611 B.n571 VSUBS 0.007437f
C612 B.n572 VSUBS 0.007437f
C613 B.n573 VSUBS 0.007437f
C614 B.n574 VSUBS 0.007437f
C615 B.n575 VSUBS 0.007437f
C616 B.n576 VSUBS 0.007437f
C617 B.n577 VSUBS 0.007437f
C618 B.n578 VSUBS 0.007437f
C619 B.n579 VSUBS 0.007437f
C620 B.n580 VSUBS 0.007437f
C621 B.n581 VSUBS 0.007437f
C622 B.n582 VSUBS 0.007437f
C623 B.n583 VSUBS 0.007437f
C624 B.n584 VSUBS 0.007437f
C625 B.n585 VSUBS 0.007437f
C626 B.n586 VSUBS 0.007437f
C627 B.n587 VSUBS 0.007437f
C628 B.n588 VSUBS 0.007437f
C629 B.n589 VSUBS 0.007437f
C630 B.n590 VSUBS 0.007437f
C631 B.n591 VSUBS 0.007437f
C632 B.n592 VSUBS 0.007437f
C633 B.n593 VSUBS 0.007437f
C634 B.n594 VSUBS 0.007437f
C635 B.n595 VSUBS 0.007437f
C636 B.n596 VSUBS 0.007437f
C637 B.n597 VSUBS 0.007437f
C638 B.n598 VSUBS 0.007437f
C639 B.n599 VSUBS 0.007437f
C640 B.n600 VSUBS 0.007437f
C641 B.n601 VSUBS 0.007437f
C642 B.n602 VSUBS 0.007437f
C643 B.n603 VSUBS 0.007437f
C644 B.n604 VSUBS 0.007437f
C645 B.n605 VSUBS 0.007437f
C646 B.n606 VSUBS 0.007437f
C647 B.n607 VSUBS 0.007437f
C648 B.n608 VSUBS 0.007437f
C649 B.n609 VSUBS 0.007437f
C650 B.n610 VSUBS 0.007437f
C651 B.n611 VSUBS 0.007437f
C652 B.n612 VSUBS 0.007437f
C653 B.n613 VSUBS 0.007437f
C654 B.n614 VSUBS 0.007437f
C655 B.n615 VSUBS 0.007437f
C656 B.n616 VSUBS 0.007437f
C657 B.n617 VSUBS 0.007437f
C658 B.n618 VSUBS 0.007437f
C659 B.n619 VSUBS 0.007437f
C660 B.n620 VSUBS 0.007437f
C661 B.n621 VSUBS 0.007437f
C662 B.n622 VSUBS 0.007437f
C663 B.n623 VSUBS 0.007437f
C664 B.n624 VSUBS 0.007437f
C665 B.n625 VSUBS 0.007437f
C666 B.n626 VSUBS 0.007437f
C667 B.n627 VSUBS 0.007437f
C668 B.n628 VSUBS 0.007437f
C669 B.n629 VSUBS 0.007437f
C670 B.n630 VSUBS 0.007437f
C671 B.n631 VSUBS 0.007437f
C672 B.n632 VSUBS 0.007437f
C673 B.n633 VSUBS 0.007437f
C674 B.n634 VSUBS 0.007437f
C675 B.n635 VSUBS 0.007437f
C676 B.n636 VSUBS 0.007437f
C677 B.n637 VSUBS 0.007437f
C678 B.n638 VSUBS 0.007437f
C679 B.n639 VSUBS 0.007437f
C680 B.n640 VSUBS 0.007437f
C681 B.n641 VSUBS 0.007437f
C682 B.n642 VSUBS 0.007437f
C683 B.n643 VSUBS 0.007437f
C684 B.n644 VSUBS 0.007437f
C685 B.n645 VSUBS 0.007437f
C686 B.n646 VSUBS 0.007437f
C687 B.n647 VSUBS 0.007437f
C688 B.n648 VSUBS 0.007437f
C689 B.n649 VSUBS 0.007437f
C690 B.n650 VSUBS 0.007437f
C691 B.n651 VSUBS 0.007437f
C692 B.n652 VSUBS 0.007437f
C693 B.n653 VSUBS 0.007437f
C694 B.n654 VSUBS 0.007437f
C695 B.n655 VSUBS 0.007437f
C696 B.n656 VSUBS 0.017302f
C697 B.n657 VSUBS 0.017302f
C698 B.n658 VSUBS 0.015945f
C699 B.n659 VSUBS 0.007437f
C700 B.n660 VSUBS 0.007437f
C701 B.n661 VSUBS 0.007437f
C702 B.n662 VSUBS 0.007437f
C703 B.n663 VSUBS 0.007437f
C704 B.n664 VSUBS 0.007437f
C705 B.n665 VSUBS 0.007437f
C706 B.n666 VSUBS 0.007437f
C707 B.n667 VSUBS 0.007437f
C708 B.n668 VSUBS 0.007437f
C709 B.n669 VSUBS 0.007437f
C710 B.n670 VSUBS 0.007437f
C711 B.n671 VSUBS 0.007437f
C712 B.n672 VSUBS 0.007437f
C713 B.n673 VSUBS 0.007437f
C714 B.n674 VSUBS 0.007437f
C715 B.n675 VSUBS 0.007437f
C716 B.n676 VSUBS 0.007437f
C717 B.n677 VSUBS 0.007437f
C718 B.n678 VSUBS 0.007437f
C719 B.n679 VSUBS 0.007437f
C720 B.n680 VSUBS 0.007437f
C721 B.n681 VSUBS 0.007437f
C722 B.n682 VSUBS 0.007437f
C723 B.n683 VSUBS 0.007437f
C724 B.n684 VSUBS 0.007437f
C725 B.n685 VSUBS 0.007437f
C726 B.n686 VSUBS 0.007437f
C727 B.n687 VSUBS 0.01684f
C728 VDD1.t2 VSUBS 0.39649f
C729 VDD1.t3 VSUBS 0.39649f
C730 VDD1.n0 VSUBS 3.29869f
C731 VDD1.t0 VSUBS 0.39649f
C732 VDD1.t1 VSUBS 0.39649f
C733 VDD1.n1 VSUBS 4.22518f
C734 VP.t0 VSUBS 2.50951f
C735 VP.t1 VSUBS 2.50967f
C736 VP.n0 VSUBS 3.38645f
C737 VP.n1 VSUBS 3.66408f
C738 VP.t3 VSUBS 2.47781f
C739 VP.n2 VSUBS 0.932237f
C740 VP.t2 VSUBS 2.47781f
C741 VP.n3 VSUBS 0.932237f
C742 VP.n4 VSUBS 0.066928f
C743 VTAIL.n0 VSUBS 0.023978f
C744 VTAIL.n1 VSUBS 0.021906f
C745 VTAIL.n2 VSUBS 0.011771f
C746 VTAIL.n3 VSUBS 0.027823f
C747 VTAIL.n4 VSUBS 0.012464f
C748 VTAIL.n5 VSUBS 0.021906f
C749 VTAIL.n6 VSUBS 0.011771f
C750 VTAIL.n7 VSUBS 0.027823f
C751 VTAIL.n8 VSUBS 0.012464f
C752 VTAIL.n9 VSUBS 0.021906f
C753 VTAIL.n10 VSUBS 0.012118f
C754 VTAIL.n11 VSUBS 0.027823f
C755 VTAIL.n12 VSUBS 0.012464f
C756 VTAIL.n13 VSUBS 0.021906f
C757 VTAIL.n14 VSUBS 0.011771f
C758 VTAIL.n15 VSUBS 0.027823f
C759 VTAIL.n16 VSUBS 0.012464f
C760 VTAIL.n17 VSUBS 0.021906f
C761 VTAIL.n18 VSUBS 0.011771f
C762 VTAIL.n19 VSUBS 0.027823f
C763 VTAIL.n20 VSUBS 0.012464f
C764 VTAIL.n21 VSUBS 0.021906f
C765 VTAIL.n22 VSUBS 0.011771f
C766 VTAIL.n23 VSUBS 0.027823f
C767 VTAIL.n24 VSUBS 0.012464f
C768 VTAIL.n25 VSUBS 0.021906f
C769 VTAIL.n26 VSUBS 0.011771f
C770 VTAIL.n27 VSUBS 0.027823f
C771 VTAIL.n28 VSUBS 0.012464f
C772 VTAIL.n29 VSUBS 0.021906f
C773 VTAIL.n30 VSUBS 0.011771f
C774 VTAIL.n31 VSUBS 0.020867f
C775 VTAIL.n32 VSUBS 0.0177f
C776 VTAIL.t5 VSUBS 0.05974f
C777 VTAIL.n33 VSUBS 0.175353f
C778 VTAIL.n34 VSUBS 1.72095f
C779 VTAIL.n35 VSUBS 0.011771f
C780 VTAIL.n36 VSUBS 0.012464f
C781 VTAIL.n37 VSUBS 0.027823f
C782 VTAIL.n38 VSUBS 0.027823f
C783 VTAIL.n39 VSUBS 0.012464f
C784 VTAIL.n40 VSUBS 0.011771f
C785 VTAIL.n41 VSUBS 0.021906f
C786 VTAIL.n42 VSUBS 0.021906f
C787 VTAIL.n43 VSUBS 0.011771f
C788 VTAIL.n44 VSUBS 0.012464f
C789 VTAIL.n45 VSUBS 0.027823f
C790 VTAIL.n46 VSUBS 0.027823f
C791 VTAIL.n47 VSUBS 0.012464f
C792 VTAIL.n48 VSUBS 0.011771f
C793 VTAIL.n49 VSUBS 0.021906f
C794 VTAIL.n50 VSUBS 0.021906f
C795 VTAIL.n51 VSUBS 0.011771f
C796 VTAIL.n52 VSUBS 0.012464f
C797 VTAIL.n53 VSUBS 0.027823f
C798 VTAIL.n54 VSUBS 0.027823f
C799 VTAIL.n55 VSUBS 0.012464f
C800 VTAIL.n56 VSUBS 0.011771f
C801 VTAIL.n57 VSUBS 0.021906f
C802 VTAIL.n58 VSUBS 0.021906f
C803 VTAIL.n59 VSUBS 0.011771f
C804 VTAIL.n60 VSUBS 0.012464f
C805 VTAIL.n61 VSUBS 0.027823f
C806 VTAIL.n62 VSUBS 0.027823f
C807 VTAIL.n63 VSUBS 0.012464f
C808 VTAIL.n64 VSUBS 0.011771f
C809 VTAIL.n65 VSUBS 0.021906f
C810 VTAIL.n66 VSUBS 0.021906f
C811 VTAIL.n67 VSUBS 0.011771f
C812 VTAIL.n68 VSUBS 0.012464f
C813 VTAIL.n69 VSUBS 0.027823f
C814 VTAIL.n70 VSUBS 0.027823f
C815 VTAIL.n71 VSUBS 0.012464f
C816 VTAIL.n72 VSUBS 0.011771f
C817 VTAIL.n73 VSUBS 0.021906f
C818 VTAIL.n74 VSUBS 0.021906f
C819 VTAIL.n75 VSUBS 0.011771f
C820 VTAIL.n76 VSUBS 0.011771f
C821 VTAIL.n77 VSUBS 0.012464f
C822 VTAIL.n78 VSUBS 0.027823f
C823 VTAIL.n79 VSUBS 0.027823f
C824 VTAIL.n80 VSUBS 0.027823f
C825 VTAIL.n81 VSUBS 0.012118f
C826 VTAIL.n82 VSUBS 0.011771f
C827 VTAIL.n83 VSUBS 0.021906f
C828 VTAIL.n84 VSUBS 0.021906f
C829 VTAIL.n85 VSUBS 0.011771f
C830 VTAIL.n86 VSUBS 0.012464f
C831 VTAIL.n87 VSUBS 0.027823f
C832 VTAIL.n88 VSUBS 0.027823f
C833 VTAIL.n89 VSUBS 0.012464f
C834 VTAIL.n90 VSUBS 0.011771f
C835 VTAIL.n91 VSUBS 0.021906f
C836 VTAIL.n92 VSUBS 0.021906f
C837 VTAIL.n93 VSUBS 0.011771f
C838 VTAIL.n94 VSUBS 0.012464f
C839 VTAIL.n95 VSUBS 0.027823f
C840 VTAIL.n96 VSUBS 0.067045f
C841 VTAIL.n97 VSUBS 0.012464f
C842 VTAIL.n98 VSUBS 0.011771f
C843 VTAIL.n99 VSUBS 0.050635f
C844 VTAIL.n100 VSUBS 0.033702f
C845 VTAIL.n101 VSUBS 0.093707f
C846 VTAIL.n102 VSUBS 0.023978f
C847 VTAIL.n103 VSUBS 0.021906f
C848 VTAIL.n104 VSUBS 0.011771f
C849 VTAIL.n105 VSUBS 0.027823f
C850 VTAIL.n106 VSUBS 0.012464f
C851 VTAIL.n107 VSUBS 0.021906f
C852 VTAIL.n108 VSUBS 0.011771f
C853 VTAIL.n109 VSUBS 0.027823f
C854 VTAIL.n110 VSUBS 0.012464f
C855 VTAIL.n111 VSUBS 0.021906f
C856 VTAIL.n112 VSUBS 0.012118f
C857 VTAIL.n113 VSUBS 0.027823f
C858 VTAIL.n114 VSUBS 0.012464f
C859 VTAIL.n115 VSUBS 0.021906f
C860 VTAIL.n116 VSUBS 0.011771f
C861 VTAIL.n117 VSUBS 0.027823f
C862 VTAIL.n118 VSUBS 0.012464f
C863 VTAIL.n119 VSUBS 0.021906f
C864 VTAIL.n120 VSUBS 0.011771f
C865 VTAIL.n121 VSUBS 0.027823f
C866 VTAIL.n122 VSUBS 0.012464f
C867 VTAIL.n123 VSUBS 0.021906f
C868 VTAIL.n124 VSUBS 0.011771f
C869 VTAIL.n125 VSUBS 0.027823f
C870 VTAIL.n126 VSUBS 0.012464f
C871 VTAIL.n127 VSUBS 0.021906f
C872 VTAIL.n128 VSUBS 0.011771f
C873 VTAIL.n129 VSUBS 0.027823f
C874 VTAIL.n130 VSUBS 0.012464f
C875 VTAIL.n131 VSUBS 0.021906f
C876 VTAIL.n132 VSUBS 0.011771f
C877 VTAIL.n133 VSUBS 0.020867f
C878 VTAIL.n134 VSUBS 0.0177f
C879 VTAIL.t2 VSUBS 0.05974f
C880 VTAIL.n135 VSUBS 0.175353f
C881 VTAIL.n136 VSUBS 1.72095f
C882 VTAIL.n137 VSUBS 0.011771f
C883 VTAIL.n138 VSUBS 0.012464f
C884 VTAIL.n139 VSUBS 0.027823f
C885 VTAIL.n140 VSUBS 0.027823f
C886 VTAIL.n141 VSUBS 0.012464f
C887 VTAIL.n142 VSUBS 0.011771f
C888 VTAIL.n143 VSUBS 0.021906f
C889 VTAIL.n144 VSUBS 0.021906f
C890 VTAIL.n145 VSUBS 0.011771f
C891 VTAIL.n146 VSUBS 0.012464f
C892 VTAIL.n147 VSUBS 0.027823f
C893 VTAIL.n148 VSUBS 0.027823f
C894 VTAIL.n149 VSUBS 0.012464f
C895 VTAIL.n150 VSUBS 0.011771f
C896 VTAIL.n151 VSUBS 0.021906f
C897 VTAIL.n152 VSUBS 0.021906f
C898 VTAIL.n153 VSUBS 0.011771f
C899 VTAIL.n154 VSUBS 0.012464f
C900 VTAIL.n155 VSUBS 0.027823f
C901 VTAIL.n156 VSUBS 0.027823f
C902 VTAIL.n157 VSUBS 0.012464f
C903 VTAIL.n158 VSUBS 0.011771f
C904 VTAIL.n159 VSUBS 0.021906f
C905 VTAIL.n160 VSUBS 0.021906f
C906 VTAIL.n161 VSUBS 0.011771f
C907 VTAIL.n162 VSUBS 0.012464f
C908 VTAIL.n163 VSUBS 0.027823f
C909 VTAIL.n164 VSUBS 0.027823f
C910 VTAIL.n165 VSUBS 0.012464f
C911 VTAIL.n166 VSUBS 0.011771f
C912 VTAIL.n167 VSUBS 0.021906f
C913 VTAIL.n168 VSUBS 0.021906f
C914 VTAIL.n169 VSUBS 0.011771f
C915 VTAIL.n170 VSUBS 0.012464f
C916 VTAIL.n171 VSUBS 0.027823f
C917 VTAIL.n172 VSUBS 0.027823f
C918 VTAIL.n173 VSUBS 0.012464f
C919 VTAIL.n174 VSUBS 0.011771f
C920 VTAIL.n175 VSUBS 0.021906f
C921 VTAIL.n176 VSUBS 0.021906f
C922 VTAIL.n177 VSUBS 0.011771f
C923 VTAIL.n178 VSUBS 0.011771f
C924 VTAIL.n179 VSUBS 0.012464f
C925 VTAIL.n180 VSUBS 0.027823f
C926 VTAIL.n181 VSUBS 0.027823f
C927 VTAIL.n182 VSUBS 0.027823f
C928 VTAIL.n183 VSUBS 0.012118f
C929 VTAIL.n184 VSUBS 0.011771f
C930 VTAIL.n185 VSUBS 0.021906f
C931 VTAIL.n186 VSUBS 0.021906f
C932 VTAIL.n187 VSUBS 0.011771f
C933 VTAIL.n188 VSUBS 0.012464f
C934 VTAIL.n189 VSUBS 0.027823f
C935 VTAIL.n190 VSUBS 0.027823f
C936 VTAIL.n191 VSUBS 0.012464f
C937 VTAIL.n192 VSUBS 0.011771f
C938 VTAIL.n193 VSUBS 0.021906f
C939 VTAIL.n194 VSUBS 0.021906f
C940 VTAIL.n195 VSUBS 0.011771f
C941 VTAIL.n196 VSUBS 0.012464f
C942 VTAIL.n197 VSUBS 0.027823f
C943 VTAIL.n198 VSUBS 0.067045f
C944 VTAIL.n199 VSUBS 0.012464f
C945 VTAIL.n200 VSUBS 0.011771f
C946 VTAIL.n201 VSUBS 0.050635f
C947 VTAIL.n202 VSUBS 0.033702f
C948 VTAIL.n203 VSUBS 0.127327f
C949 VTAIL.n204 VSUBS 0.023978f
C950 VTAIL.n205 VSUBS 0.021906f
C951 VTAIL.n206 VSUBS 0.011771f
C952 VTAIL.n207 VSUBS 0.027823f
C953 VTAIL.n208 VSUBS 0.012464f
C954 VTAIL.n209 VSUBS 0.021906f
C955 VTAIL.n210 VSUBS 0.011771f
C956 VTAIL.n211 VSUBS 0.027823f
C957 VTAIL.n212 VSUBS 0.012464f
C958 VTAIL.n213 VSUBS 0.021906f
C959 VTAIL.n214 VSUBS 0.012118f
C960 VTAIL.n215 VSUBS 0.027823f
C961 VTAIL.n216 VSUBS 0.012464f
C962 VTAIL.n217 VSUBS 0.021906f
C963 VTAIL.n218 VSUBS 0.011771f
C964 VTAIL.n219 VSUBS 0.027823f
C965 VTAIL.n220 VSUBS 0.012464f
C966 VTAIL.n221 VSUBS 0.021906f
C967 VTAIL.n222 VSUBS 0.011771f
C968 VTAIL.n223 VSUBS 0.027823f
C969 VTAIL.n224 VSUBS 0.012464f
C970 VTAIL.n225 VSUBS 0.021906f
C971 VTAIL.n226 VSUBS 0.011771f
C972 VTAIL.n227 VSUBS 0.027823f
C973 VTAIL.n228 VSUBS 0.012464f
C974 VTAIL.n229 VSUBS 0.021906f
C975 VTAIL.n230 VSUBS 0.011771f
C976 VTAIL.n231 VSUBS 0.027823f
C977 VTAIL.n232 VSUBS 0.012464f
C978 VTAIL.n233 VSUBS 0.021906f
C979 VTAIL.n234 VSUBS 0.011771f
C980 VTAIL.n235 VSUBS 0.020867f
C981 VTAIL.n236 VSUBS 0.0177f
C982 VTAIL.t0 VSUBS 0.05974f
C983 VTAIL.n237 VSUBS 0.175353f
C984 VTAIL.n238 VSUBS 1.72095f
C985 VTAIL.n239 VSUBS 0.011771f
C986 VTAIL.n240 VSUBS 0.012464f
C987 VTAIL.n241 VSUBS 0.027823f
C988 VTAIL.n242 VSUBS 0.027823f
C989 VTAIL.n243 VSUBS 0.012464f
C990 VTAIL.n244 VSUBS 0.011771f
C991 VTAIL.n245 VSUBS 0.021906f
C992 VTAIL.n246 VSUBS 0.021906f
C993 VTAIL.n247 VSUBS 0.011771f
C994 VTAIL.n248 VSUBS 0.012464f
C995 VTAIL.n249 VSUBS 0.027823f
C996 VTAIL.n250 VSUBS 0.027823f
C997 VTAIL.n251 VSUBS 0.012464f
C998 VTAIL.n252 VSUBS 0.011771f
C999 VTAIL.n253 VSUBS 0.021906f
C1000 VTAIL.n254 VSUBS 0.021906f
C1001 VTAIL.n255 VSUBS 0.011771f
C1002 VTAIL.n256 VSUBS 0.012464f
C1003 VTAIL.n257 VSUBS 0.027823f
C1004 VTAIL.n258 VSUBS 0.027823f
C1005 VTAIL.n259 VSUBS 0.012464f
C1006 VTAIL.n260 VSUBS 0.011771f
C1007 VTAIL.n261 VSUBS 0.021906f
C1008 VTAIL.n262 VSUBS 0.021906f
C1009 VTAIL.n263 VSUBS 0.011771f
C1010 VTAIL.n264 VSUBS 0.012464f
C1011 VTAIL.n265 VSUBS 0.027823f
C1012 VTAIL.n266 VSUBS 0.027823f
C1013 VTAIL.n267 VSUBS 0.012464f
C1014 VTAIL.n268 VSUBS 0.011771f
C1015 VTAIL.n269 VSUBS 0.021906f
C1016 VTAIL.n270 VSUBS 0.021906f
C1017 VTAIL.n271 VSUBS 0.011771f
C1018 VTAIL.n272 VSUBS 0.012464f
C1019 VTAIL.n273 VSUBS 0.027823f
C1020 VTAIL.n274 VSUBS 0.027823f
C1021 VTAIL.n275 VSUBS 0.012464f
C1022 VTAIL.n276 VSUBS 0.011771f
C1023 VTAIL.n277 VSUBS 0.021906f
C1024 VTAIL.n278 VSUBS 0.021906f
C1025 VTAIL.n279 VSUBS 0.011771f
C1026 VTAIL.n280 VSUBS 0.011771f
C1027 VTAIL.n281 VSUBS 0.012464f
C1028 VTAIL.n282 VSUBS 0.027823f
C1029 VTAIL.n283 VSUBS 0.027823f
C1030 VTAIL.n284 VSUBS 0.027823f
C1031 VTAIL.n285 VSUBS 0.012118f
C1032 VTAIL.n286 VSUBS 0.011771f
C1033 VTAIL.n287 VSUBS 0.021906f
C1034 VTAIL.n288 VSUBS 0.021906f
C1035 VTAIL.n289 VSUBS 0.011771f
C1036 VTAIL.n290 VSUBS 0.012464f
C1037 VTAIL.n291 VSUBS 0.027823f
C1038 VTAIL.n292 VSUBS 0.027823f
C1039 VTAIL.n293 VSUBS 0.012464f
C1040 VTAIL.n294 VSUBS 0.011771f
C1041 VTAIL.n295 VSUBS 0.021906f
C1042 VTAIL.n296 VSUBS 0.021906f
C1043 VTAIL.n297 VSUBS 0.011771f
C1044 VTAIL.n298 VSUBS 0.012464f
C1045 VTAIL.n299 VSUBS 0.027823f
C1046 VTAIL.n300 VSUBS 0.067045f
C1047 VTAIL.n301 VSUBS 0.012464f
C1048 VTAIL.n302 VSUBS 0.011771f
C1049 VTAIL.n303 VSUBS 0.050635f
C1050 VTAIL.n304 VSUBS 0.033702f
C1051 VTAIL.n305 VSUBS 1.57709f
C1052 VTAIL.n306 VSUBS 0.023978f
C1053 VTAIL.n307 VSUBS 0.021906f
C1054 VTAIL.n308 VSUBS 0.011771f
C1055 VTAIL.n309 VSUBS 0.027823f
C1056 VTAIL.n310 VSUBS 0.012464f
C1057 VTAIL.n311 VSUBS 0.021906f
C1058 VTAIL.n312 VSUBS 0.011771f
C1059 VTAIL.n313 VSUBS 0.027823f
C1060 VTAIL.n314 VSUBS 0.012464f
C1061 VTAIL.n315 VSUBS 0.021906f
C1062 VTAIL.n316 VSUBS 0.012118f
C1063 VTAIL.n317 VSUBS 0.027823f
C1064 VTAIL.n318 VSUBS 0.011771f
C1065 VTAIL.n319 VSUBS 0.012464f
C1066 VTAIL.n320 VSUBS 0.021906f
C1067 VTAIL.n321 VSUBS 0.011771f
C1068 VTAIL.n322 VSUBS 0.027823f
C1069 VTAIL.n323 VSUBS 0.012464f
C1070 VTAIL.n324 VSUBS 0.021906f
C1071 VTAIL.n325 VSUBS 0.011771f
C1072 VTAIL.n326 VSUBS 0.027823f
C1073 VTAIL.n327 VSUBS 0.012464f
C1074 VTAIL.n328 VSUBS 0.021906f
C1075 VTAIL.n329 VSUBS 0.011771f
C1076 VTAIL.n330 VSUBS 0.027823f
C1077 VTAIL.n331 VSUBS 0.012464f
C1078 VTAIL.n332 VSUBS 0.021906f
C1079 VTAIL.n333 VSUBS 0.011771f
C1080 VTAIL.n334 VSUBS 0.027823f
C1081 VTAIL.n335 VSUBS 0.012464f
C1082 VTAIL.n336 VSUBS 0.021906f
C1083 VTAIL.n337 VSUBS 0.011771f
C1084 VTAIL.n338 VSUBS 0.020867f
C1085 VTAIL.n339 VSUBS 0.0177f
C1086 VTAIL.t7 VSUBS 0.05974f
C1087 VTAIL.n340 VSUBS 0.175353f
C1088 VTAIL.n341 VSUBS 1.72095f
C1089 VTAIL.n342 VSUBS 0.011771f
C1090 VTAIL.n343 VSUBS 0.012464f
C1091 VTAIL.n344 VSUBS 0.027823f
C1092 VTAIL.n345 VSUBS 0.027823f
C1093 VTAIL.n346 VSUBS 0.012464f
C1094 VTAIL.n347 VSUBS 0.011771f
C1095 VTAIL.n348 VSUBS 0.021906f
C1096 VTAIL.n349 VSUBS 0.021906f
C1097 VTAIL.n350 VSUBS 0.011771f
C1098 VTAIL.n351 VSUBS 0.012464f
C1099 VTAIL.n352 VSUBS 0.027823f
C1100 VTAIL.n353 VSUBS 0.027823f
C1101 VTAIL.n354 VSUBS 0.012464f
C1102 VTAIL.n355 VSUBS 0.011771f
C1103 VTAIL.n356 VSUBS 0.021906f
C1104 VTAIL.n357 VSUBS 0.021906f
C1105 VTAIL.n358 VSUBS 0.011771f
C1106 VTAIL.n359 VSUBS 0.012464f
C1107 VTAIL.n360 VSUBS 0.027823f
C1108 VTAIL.n361 VSUBS 0.027823f
C1109 VTAIL.n362 VSUBS 0.012464f
C1110 VTAIL.n363 VSUBS 0.011771f
C1111 VTAIL.n364 VSUBS 0.021906f
C1112 VTAIL.n365 VSUBS 0.021906f
C1113 VTAIL.n366 VSUBS 0.011771f
C1114 VTAIL.n367 VSUBS 0.012464f
C1115 VTAIL.n368 VSUBS 0.027823f
C1116 VTAIL.n369 VSUBS 0.027823f
C1117 VTAIL.n370 VSUBS 0.012464f
C1118 VTAIL.n371 VSUBS 0.011771f
C1119 VTAIL.n372 VSUBS 0.021906f
C1120 VTAIL.n373 VSUBS 0.021906f
C1121 VTAIL.n374 VSUBS 0.011771f
C1122 VTAIL.n375 VSUBS 0.012464f
C1123 VTAIL.n376 VSUBS 0.027823f
C1124 VTAIL.n377 VSUBS 0.027823f
C1125 VTAIL.n378 VSUBS 0.012464f
C1126 VTAIL.n379 VSUBS 0.011771f
C1127 VTAIL.n380 VSUBS 0.021906f
C1128 VTAIL.n381 VSUBS 0.021906f
C1129 VTAIL.n382 VSUBS 0.011771f
C1130 VTAIL.n383 VSUBS 0.012464f
C1131 VTAIL.n384 VSUBS 0.027823f
C1132 VTAIL.n385 VSUBS 0.027823f
C1133 VTAIL.n386 VSUBS 0.027823f
C1134 VTAIL.n387 VSUBS 0.012118f
C1135 VTAIL.n388 VSUBS 0.011771f
C1136 VTAIL.n389 VSUBS 0.021906f
C1137 VTAIL.n390 VSUBS 0.021906f
C1138 VTAIL.n391 VSUBS 0.011771f
C1139 VTAIL.n392 VSUBS 0.012464f
C1140 VTAIL.n393 VSUBS 0.027823f
C1141 VTAIL.n394 VSUBS 0.027823f
C1142 VTAIL.n395 VSUBS 0.012464f
C1143 VTAIL.n396 VSUBS 0.011771f
C1144 VTAIL.n397 VSUBS 0.021906f
C1145 VTAIL.n398 VSUBS 0.021906f
C1146 VTAIL.n399 VSUBS 0.011771f
C1147 VTAIL.n400 VSUBS 0.012464f
C1148 VTAIL.n401 VSUBS 0.027823f
C1149 VTAIL.n402 VSUBS 0.067045f
C1150 VTAIL.n403 VSUBS 0.012464f
C1151 VTAIL.n404 VSUBS 0.011771f
C1152 VTAIL.n405 VSUBS 0.050635f
C1153 VTAIL.n406 VSUBS 0.033702f
C1154 VTAIL.n407 VSUBS 1.57709f
C1155 VTAIL.n408 VSUBS 0.023978f
C1156 VTAIL.n409 VSUBS 0.021906f
C1157 VTAIL.n410 VSUBS 0.011771f
C1158 VTAIL.n411 VSUBS 0.027823f
C1159 VTAIL.n412 VSUBS 0.012464f
C1160 VTAIL.n413 VSUBS 0.021906f
C1161 VTAIL.n414 VSUBS 0.011771f
C1162 VTAIL.n415 VSUBS 0.027823f
C1163 VTAIL.n416 VSUBS 0.012464f
C1164 VTAIL.n417 VSUBS 0.021906f
C1165 VTAIL.n418 VSUBS 0.012118f
C1166 VTAIL.n419 VSUBS 0.027823f
C1167 VTAIL.n420 VSUBS 0.011771f
C1168 VTAIL.n421 VSUBS 0.012464f
C1169 VTAIL.n422 VSUBS 0.021906f
C1170 VTAIL.n423 VSUBS 0.011771f
C1171 VTAIL.n424 VSUBS 0.027823f
C1172 VTAIL.n425 VSUBS 0.012464f
C1173 VTAIL.n426 VSUBS 0.021906f
C1174 VTAIL.n427 VSUBS 0.011771f
C1175 VTAIL.n428 VSUBS 0.027823f
C1176 VTAIL.n429 VSUBS 0.012464f
C1177 VTAIL.n430 VSUBS 0.021906f
C1178 VTAIL.n431 VSUBS 0.011771f
C1179 VTAIL.n432 VSUBS 0.027823f
C1180 VTAIL.n433 VSUBS 0.012464f
C1181 VTAIL.n434 VSUBS 0.021906f
C1182 VTAIL.n435 VSUBS 0.011771f
C1183 VTAIL.n436 VSUBS 0.027823f
C1184 VTAIL.n437 VSUBS 0.012464f
C1185 VTAIL.n438 VSUBS 0.021906f
C1186 VTAIL.n439 VSUBS 0.011771f
C1187 VTAIL.n440 VSUBS 0.020867f
C1188 VTAIL.n441 VSUBS 0.0177f
C1189 VTAIL.t6 VSUBS 0.05974f
C1190 VTAIL.n442 VSUBS 0.175353f
C1191 VTAIL.n443 VSUBS 1.72095f
C1192 VTAIL.n444 VSUBS 0.011771f
C1193 VTAIL.n445 VSUBS 0.012464f
C1194 VTAIL.n446 VSUBS 0.027823f
C1195 VTAIL.n447 VSUBS 0.027823f
C1196 VTAIL.n448 VSUBS 0.012464f
C1197 VTAIL.n449 VSUBS 0.011771f
C1198 VTAIL.n450 VSUBS 0.021906f
C1199 VTAIL.n451 VSUBS 0.021906f
C1200 VTAIL.n452 VSUBS 0.011771f
C1201 VTAIL.n453 VSUBS 0.012464f
C1202 VTAIL.n454 VSUBS 0.027823f
C1203 VTAIL.n455 VSUBS 0.027823f
C1204 VTAIL.n456 VSUBS 0.012464f
C1205 VTAIL.n457 VSUBS 0.011771f
C1206 VTAIL.n458 VSUBS 0.021906f
C1207 VTAIL.n459 VSUBS 0.021906f
C1208 VTAIL.n460 VSUBS 0.011771f
C1209 VTAIL.n461 VSUBS 0.012464f
C1210 VTAIL.n462 VSUBS 0.027823f
C1211 VTAIL.n463 VSUBS 0.027823f
C1212 VTAIL.n464 VSUBS 0.012464f
C1213 VTAIL.n465 VSUBS 0.011771f
C1214 VTAIL.n466 VSUBS 0.021906f
C1215 VTAIL.n467 VSUBS 0.021906f
C1216 VTAIL.n468 VSUBS 0.011771f
C1217 VTAIL.n469 VSUBS 0.012464f
C1218 VTAIL.n470 VSUBS 0.027823f
C1219 VTAIL.n471 VSUBS 0.027823f
C1220 VTAIL.n472 VSUBS 0.012464f
C1221 VTAIL.n473 VSUBS 0.011771f
C1222 VTAIL.n474 VSUBS 0.021906f
C1223 VTAIL.n475 VSUBS 0.021906f
C1224 VTAIL.n476 VSUBS 0.011771f
C1225 VTAIL.n477 VSUBS 0.012464f
C1226 VTAIL.n478 VSUBS 0.027823f
C1227 VTAIL.n479 VSUBS 0.027823f
C1228 VTAIL.n480 VSUBS 0.012464f
C1229 VTAIL.n481 VSUBS 0.011771f
C1230 VTAIL.n482 VSUBS 0.021906f
C1231 VTAIL.n483 VSUBS 0.021906f
C1232 VTAIL.n484 VSUBS 0.011771f
C1233 VTAIL.n485 VSUBS 0.012464f
C1234 VTAIL.n486 VSUBS 0.027823f
C1235 VTAIL.n487 VSUBS 0.027823f
C1236 VTAIL.n488 VSUBS 0.027823f
C1237 VTAIL.n489 VSUBS 0.012118f
C1238 VTAIL.n490 VSUBS 0.011771f
C1239 VTAIL.n491 VSUBS 0.021906f
C1240 VTAIL.n492 VSUBS 0.021906f
C1241 VTAIL.n493 VSUBS 0.011771f
C1242 VTAIL.n494 VSUBS 0.012464f
C1243 VTAIL.n495 VSUBS 0.027823f
C1244 VTAIL.n496 VSUBS 0.027823f
C1245 VTAIL.n497 VSUBS 0.012464f
C1246 VTAIL.n498 VSUBS 0.011771f
C1247 VTAIL.n499 VSUBS 0.021906f
C1248 VTAIL.n500 VSUBS 0.021906f
C1249 VTAIL.n501 VSUBS 0.011771f
C1250 VTAIL.n502 VSUBS 0.012464f
C1251 VTAIL.n503 VSUBS 0.027823f
C1252 VTAIL.n504 VSUBS 0.067045f
C1253 VTAIL.n505 VSUBS 0.012464f
C1254 VTAIL.n506 VSUBS 0.011771f
C1255 VTAIL.n507 VSUBS 0.050635f
C1256 VTAIL.n508 VSUBS 0.033702f
C1257 VTAIL.n509 VSUBS 0.127327f
C1258 VTAIL.n510 VSUBS 0.023978f
C1259 VTAIL.n511 VSUBS 0.021906f
C1260 VTAIL.n512 VSUBS 0.011771f
C1261 VTAIL.n513 VSUBS 0.027823f
C1262 VTAIL.n514 VSUBS 0.012464f
C1263 VTAIL.n515 VSUBS 0.021906f
C1264 VTAIL.n516 VSUBS 0.011771f
C1265 VTAIL.n517 VSUBS 0.027823f
C1266 VTAIL.n518 VSUBS 0.012464f
C1267 VTAIL.n519 VSUBS 0.021906f
C1268 VTAIL.n520 VSUBS 0.012118f
C1269 VTAIL.n521 VSUBS 0.027823f
C1270 VTAIL.n522 VSUBS 0.011771f
C1271 VTAIL.n523 VSUBS 0.012464f
C1272 VTAIL.n524 VSUBS 0.021906f
C1273 VTAIL.n525 VSUBS 0.011771f
C1274 VTAIL.n526 VSUBS 0.027823f
C1275 VTAIL.n527 VSUBS 0.012464f
C1276 VTAIL.n528 VSUBS 0.021906f
C1277 VTAIL.n529 VSUBS 0.011771f
C1278 VTAIL.n530 VSUBS 0.027823f
C1279 VTAIL.n531 VSUBS 0.012464f
C1280 VTAIL.n532 VSUBS 0.021906f
C1281 VTAIL.n533 VSUBS 0.011771f
C1282 VTAIL.n534 VSUBS 0.027823f
C1283 VTAIL.n535 VSUBS 0.012464f
C1284 VTAIL.n536 VSUBS 0.021906f
C1285 VTAIL.n537 VSUBS 0.011771f
C1286 VTAIL.n538 VSUBS 0.027823f
C1287 VTAIL.n539 VSUBS 0.012464f
C1288 VTAIL.n540 VSUBS 0.021906f
C1289 VTAIL.n541 VSUBS 0.011771f
C1290 VTAIL.n542 VSUBS 0.020867f
C1291 VTAIL.n543 VSUBS 0.0177f
C1292 VTAIL.t3 VSUBS 0.05974f
C1293 VTAIL.n544 VSUBS 0.175353f
C1294 VTAIL.n545 VSUBS 1.72095f
C1295 VTAIL.n546 VSUBS 0.011771f
C1296 VTAIL.n547 VSUBS 0.012464f
C1297 VTAIL.n548 VSUBS 0.027823f
C1298 VTAIL.n549 VSUBS 0.027823f
C1299 VTAIL.n550 VSUBS 0.012464f
C1300 VTAIL.n551 VSUBS 0.011771f
C1301 VTAIL.n552 VSUBS 0.021906f
C1302 VTAIL.n553 VSUBS 0.021906f
C1303 VTAIL.n554 VSUBS 0.011771f
C1304 VTAIL.n555 VSUBS 0.012464f
C1305 VTAIL.n556 VSUBS 0.027823f
C1306 VTAIL.n557 VSUBS 0.027823f
C1307 VTAIL.n558 VSUBS 0.012464f
C1308 VTAIL.n559 VSUBS 0.011771f
C1309 VTAIL.n560 VSUBS 0.021906f
C1310 VTAIL.n561 VSUBS 0.021906f
C1311 VTAIL.n562 VSUBS 0.011771f
C1312 VTAIL.n563 VSUBS 0.012464f
C1313 VTAIL.n564 VSUBS 0.027823f
C1314 VTAIL.n565 VSUBS 0.027823f
C1315 VTAIL.n566 VSUBS 0.012464f
C1316 VTAIL.n567 VSUBS 0.011771f
C1317 VTAIL.n568 VSUBS 0.021906f
C1318 VTAIL.n569 VSUBS 0.021906f
C1319 VTAIL.n570 VSUBS 0.011771f
C1320 VTAIL.n571 VSUBS 0.012464f
C1321 VTAIL.n572 VSUBS 0.027823f
C1322 VTAIL.n573 VSUBS 0.027823f
C1323 VTAIL.n574 VSUBS 0.012464f
C1324 VTAIL.n575 VSUBS 0.011771f
C1325 VTAIL.n576 VSUBS 0.021906f
C1326 VTAIL.n577 VSUBS 0.021906f
C1327 VTAIL.n578 VSUBS 0.011771f
C1328 VTAIL.n579 VSUBS 0.012464f
C1329 VTAIL.n580 VSUBS 0.027823f
C1330 VTAIL.n581 VSUBS 0.027823f
C1331 VTAIL.n582 VSUBS 0.012464f
C1332 VTAIL.n583 VSUBS 0.011771f
C1333 VTAIL.n584 VSUBS 0.021906f
C1334 VTAIL.n585 VSUBS 0.021906f
C1335 VTAIL.n586 VSUBS 0.011771f
C1336 VTAIL.n587 VSUBS 0.012464f
C1337 VTAIL.n588 VSUBS 0.027823f
C1338 VTAIL.n589 VSUBS 0.027823f
C1339 VTAIL.n590 VSUBS 0.027823f
C1340 VTAIL.n591 VSUBS 0.012118f
C1341 VTAIL.n592 VSUBS 0.011771f
C1342 VTAIL.n593 VSUBS 0.021906f
C1343 VTAIL.n594 VSUBS 0.021906f
C1344 VTAIL.n595 VSUBS 0.011771f
C1345 VTAIL.n596 VSUBS 0.012464f
C1346 VTAIL.n597 VSUBS 0.027823f
C1347 VTAIL.n598 VSUBS 0.027823f
C1348 VTAIL.n599 VSUBS 0.012464f
C1349 VTAIL.n600 VSUBS 0.011771f
C1350 VTAIL.n601 VSUBS 0.021906f
C1351 VTAIL.n602 VSUBS 0.021906f
C1352 VTAIL.n603 VSUBS 0.011771f
C1353 VTAIL.n604 VSUBS 0.012464f
C1354 VTAIL.n605 VSUBS 0.027823f
C1355 VTAIL.n606 VSUBS 0.067045f
C1356 VTAIL.n607 VSUBS 0.012464f
C1357 VTAIL.n608 VSUBS 0.011771f
C1358 VTAIL.n609 VSUBS 0.050635f
C1359 VTAIL.n610 VSUBS 0.033702f
C1360 VTAIL.n611 VSUBS 0.127327f
C1361 VTAIL.n612 VSUBS 0.023978f
C1362 VTAIL.n613 VSUBS 0.021906f
C1363 VTAIL.n614 VSUBS 0.011771f
C1364 VTAIL.n615 VSUBS 0.027823f
C1365 VTAIL.n616 VSUBS 0.012464f
C1366 VTAIL.n617 VSUBS 0.021906f
C1367 VTAIL.n618 VSUBS 0.011771f
C1368 VTAIL.n619 VSUBS 0.027823f
C1369 VTAIL.n620 VSUBS 0.012464f
C1370 VTAIL.n621 VSUBS 0.021906f
C1371 VTAIL.n622 VSUBS 0.012118f
C1372 VTAIL.n623 VSUBS 0.027823f
C1373 VTAIL.n624 VSUBS 0.011771f
C1374 VTAIL.n625 VSUBS 0.012464f
C1375 VTAIL.n626 VSUBS 0.021906f
C1376 VTAIL.n627 VSUBS 0.011771f
C1377 VTAIL.n628 VSUBS 0.027823f
C1378 VTAIL.n629 VSUBS 0.012464f
C1379 VTAIL.n630 VSUBS 0.021906f
C1380 VTAIL.n631 VSUBS 0.011771f
C1381 VTAIL.n632 VSUBS 0.027823f
C1382 VTAIL.n633 VSUBS 0.012464f
C1383 VTAIL.n634 VSUBS 0.021906f
C1384 VTAIL.n635 VSUBS 0.011771f
C1385 VTAIL.n636 VSUBS 0.027823f
C1386 VTAIL.n637 VSUBS 0.012464f
C1387 VTAIL.n638 VSUBS 0.021906f
C1388 VTAIL.n639 VSUBS 0.011771f
C1389 VTAIL.n640 VSUBS 0.027823f
C1390 VTAIL.n641 VSUBS 0.012464f
C1391 VTAIL.n642 VSUBS 0.021906f
C1392 VTAIL.n643 VSUBS 0.011771f
C1393 VTAIL.n644 VSUBS 0.020867f
C1394 VTAIL.n645 VSUBS 0.0177f
C1395 VTAIL.t1 VSUBS 0.05974f
C1396 VTAIL.n646 VSUBS 0.175353f
C1397 VTAIL.n647 VSUBS 1.72095f
C1398 VTAIL.n648 VSUBS 0.011771f
C1399 VTAIL.n649 VSUBS 0.012464f
C1400 VTAIL.n650 VSUBS 0.027823f
C1401 VTAIL.n651 VSUBS 0.027823f
C1402 VTAIL.n652 VSUBS 0.012464f
C1403 VTAIL.n653 VSUBS 0.011771f
C1404 VTAIL.n654 VSUBS 0.021906f
C1405 VTAIL.n655 VSUBS 0.021906f
C1406 VTAIL.n656 VSUBS 0.011771f
C1407 VTAIL.n657 VSUBS 0.012464f
C1408 VTAIL.n658 VSUBS 0.027823f
C1409 VTAIL.n659 VSUBS 0.027823f
C1410 VTAIL.n660 VSUBS 0.012464f
C1411 VTAIL.n661 VSUBS 0.011771f
C1412 VTAIL.n662 VSUBS 0.021906f
C1413 VTAIL.n663 VSUBS 0.021906f
C1414 VTAIL.n664 VSUBS 0.011771f
C1415 VTAIL.n665 VSUBS 0.012464f
C1416 VTAIL.n666 VSUBS 0.027823f
C1417 VTAIL.n667 VSUBS 0.027823f
C1418 VTAIL.n668 VSUBS 0.012464f
C1419 VTAIL.n669 VSUBS 0.011771f
C1420 VTAIL.n670 VSUBS 0.021906f
C1421 VTAIL.n671 VSUBS 0.021906f
C1422 VTAIL.n672 VSUBS 0.011771f
C1423 VTAIL.n673 VSUBS 0.012464f
C1424 VTAIL.n674 VSUBS 0.027823f
C1425 VTAIL.n675 VSUBS 0.027823f
C1426 VTAIL.n676 VSUBS 0.012464f
C1427 VTAIL.n677 VSUBS 0.011771f
C1428 VTAIL.n678 VSUBS 0.021906f
C1429 VTAIL.n679 VSUBS 0.021906f
C1430 VTAIL.n680 VSUBS 0.011771f
C1431 VTAIL.n681 VSUBS 0.012464f
C1432 VTAIL.n682 VSUBS 0.027823f
C1433 VTAIL.n683 VSUBS 0.027823f
C1434 VTAIL.n684 VSUBS 0.012464f
C1435 VTAIL.n685 VSUBS 0.011771f
C1436 VTAIL.n686 VSUBS 0.021906f
C1437 VTAIL.n687 VSUBS 0.021906f
C1438 VTAIL.n688 VSUBS 0.011771f
C1439 VTAIL.n689 VSUBS 0.012464f
C1440 VTAIL.n690 VSUBS 0.027823f
C1441 VTAIL.n691 VSUBS 0.027823f
C1442 VTAIL.n692 VSUBS 0.027823f
C1443 VTAIL.n693 VSUBS 0.012118f
C1444 VTAIL.n694 VSUBS 0.011771f
C1445 VTAIL.n695 VSUBS 0.021906f
C1446 VTAIL.n696 VSUBS 0.021906f
C1447 VTAIL.n697 VSUBS 0.011771f
C1448 VTAIL.n698 VSUBS 0.012464f
C1449 VTAIL.n699 VSUBS 0.027823f
C1450 VTAIL.n700 VSUBS 0.027823f
C1451 VTAIL.n701 VSUBS 0.012464f
C1452 VTAIL.n702 VSUBS 0.011771f
C1453 VTAIL.n703 VSUBS 0.021906f
C1454 VTAIL.n704 VSUBS 0.021906f
C1455 VTAIL.n705 VSUBS 0.011771f
C1456 VTAIL.n706 VSUBS 0.012464f
C1457 VTAIL.n707 VSUBS 0.027823f
C1458 VTAIL.n708 VSUBS 0.067045f
C1459 VTAIL.n709 VSUBS 0.012464f
C1460 VTAIL.n710 VSUBS 0.011771f
C1461 VTAIL.n711 VSUBS 0.050635f
C1462 VTAIL.n712 VSUBS 0.033702f
C1463 VTAIL.n713 VSUBS 1.57709f
C1464 VTAIL.n714 VSUBS 0.023978f
C1465 VTAIL.n715 VSUBS 0.021906f
C1466 VTAIL.n716 VSUBS 0.011771f
C1467 VTAIL.n717 VSUBS 0.027823f
C1468 VTAIL.n718 VSUBS 0.012464f
C1469 VTAIL.n719 VSUBS 0.021906f
C1470 VTAIL.n720 VSUBS 0.011771f
C1471 VTAIL.n721 VSUBS 0.027823f
C1472 VTAIL.n722 VSUBS 0.012464f
C1473 VTAIL.n723 VSUBS 0.021906f
C1474 VTAIL.n724 VSUBS 0.012118f
C1475 VTAIL.n725 VSUBS 0.027823f
C1476 VTAIL.n726 VSUBS 0.012464f
C1477 VTAIL.n727 VSUBS 0.021906f
C1478 VTAIL.n728 VSUBS 0.011771f
C1479 VTAIL.n729 VSUBS 0.027823f
C1480 VTAIL.n730 VSUBS 0.012464f
C1481 VTAIL.n731 VSUBS 0.021906f
C1482 VTAIL.n732 VSUBS 0.011771f
C1483 VTAIL.n733 VSUBS 0.027823f
C1484 VTAIL.n734 VSUBS 0.012464f
C1485 VTAIL.n735 VSUBS 0.021906f
C1486 VTAIL.n736 VSUBS 0.011771f
C1487 VTAIL.n737 VSUBS 0.027823f
C1488 VTAIL.n738 VSUBS 0.012464f
C1489 VTAIL.n739 VSUBS 0.021906f
C1490 VTAIL.n740 VSUBS 0.011771f
C1491 VTAIL.n741 VSUBS 0.027823f
C1492 VTAIL.n742 VSUBS 0.012464f
C1493 VTAIL.n743 VSUBS 0.021906f
C1494 VTAIL.n744 VSUBS 0.011771f
C1495 VTAIL.n745 VSUBS 0.020867f
C1496 VTAIL.n746 VSUBS 0.0177f
C1497 VTAIL.t4 VSUBS 0.05974f
C1498 VTAIL.n747 VSUBS 0.175353f
C1499 VTAIL.n748 VSUBS 1.72095f
C1500 VTAIL.n749 VSUBS 0.011771f
C1501 VTAIL.n750 VSUBS 0.012464f
C1502 VTAIL.n751 VSUBS 0.027823f
C1503 VTAIL.n752 VSUBS 0.027823f
C1504 VTAIL.n753 VSUBS 0.012464f
C1505 VTAIL.n754 VSUBS 0.011771f
C1506 VTAIL.n755 VSUBS 0.021906f
C1507 VTAIL.n756 VSUBS 0.021906f
C1508 VTAIL.n757 VSUBS 0.011771f
C1509 VTAIL.n758 VSUBS 0.012464f
C1510 VTAIL.n759 VSUBS 0.027823f
C1511 VTAIL.n760 VSUBS 0.027823f
C1512 VTAIL.n761 VSUBS 0.012464f
C1513 VTAIL.n762 VSUBS 0.011771f
C1514 VTAIL.n763 VSUBS 0.021906f
C1515 VTAIL.n764 VSUBS 0.021906f
C1516 VTAIL.n765 VSUBS 0.011771f
C1517 VTAIL.n766 VSUBS 0.012464f
C1518 VTAIL.n767 VSUBS 0.027823f
C1519 VTAIL.n768 VSUBS 0.027823f
C1520 VTAIL.n769 VSUBS 0.012464f
C1521 VTAIL.n770 VSUBS 0.011771f
C1522 VTAIL.n771 VSUBS 0.021906f
C1523 VTAIL.n772 VSUBS 0.021906f
C1524 VTAIL.n773 VSUBS 0.011771f
C1525 VTAIL.n774 VSUBS 0.012464f
C1526 VTAIL.n775 VSUBS 0.027823f
C1527 VTAIL.n776 VSUBS 0.027823f
C1528 VTAIL.n777 VSUBS 0.012464f
C1529 VTAIL.n778 VSUBS 0.011771f
C1530 VTAIL.n779 VSUBS 0.021906f
C1531 VTAIL.n780 VSUBS 0.021906f
C1532 VTAIL.n781 VSUBS 0.011771f
C1533 VTAIL.n782 VSUBS 0.012464f
C1534 VTAIL.n783 VSUBS 0.027823f
C1535 VTAIL.n784 VSUBS 0.027823f
C1536 VTAIL.n785 VSUBS 0.012464f
C1537 VTAIL.n786 VSUBS 0.011771f
C1538 VTAIL.n787 VSUBS 0.021906f
C1539 VTAIL.n788 VSUBS 0.021906f
C1540 VTAIL.n789 VSUBS 0.011771f
C1541 VTAIL.n790 VSUBS 0.011771f
C1542 VTAIL.n791 VSUBS 0.012464f
C1543 VTAIL.n792 VSUBS 0.027823f
C1544 VTAIL.n793 VSUBS 0.027823f
C1545 VTAIL.n794 VSUBS 0.027823f
C1546 VTAIL.n795 VSUBS 0.012118f
C1547 VTAIL.n796 VSUBS 0.011771f
C1548 VTAIL.n797 VSUBS 0.021906f
C1549 VTAIL.n798 VSUBS 0.021906f
C1550 VTAIL.n799 VSUBS 0.011771f
C1551 VTAIL.n800 VSUBS 0.012464f
C1552 VTAIL.n801 VSUBS 0.027823f
C1553 VTAIL.n802 VSUBS 0.027823f
C1554 VTAIL.n803 VSUBS 0.012464f
C1555 VTAIL.n804 VSUBS 0.011771f
C1556 VTAIL.n805 VSUBS 0.021906f
C1557 VTAIL.n806 VSUBS 0.021906f
C1558 VTAIL.n807 VSUBS 0.011771f
C1559 VTAIL.n808 VSUBS 0.012464f
C1560 VTAIL.n809 VSUBS 0.027823f
C1561 VTAIL.n810 VSUBS 0.067045f
C1562 VTAIL.n811 VSUBS 0.012464f
C1563 VTAIL.n812 VSUBS 0.011771f
C1564 VTAIL.n813 VSUBS 0.050635f
C1565 VTAIL.n814 VSUBS 0.033702f
C1566 VTAIL.n815 VSUBS 1.53526f
C1567 VDD2.t3 VSUBS 0.396535f
C1568 VDD2.t1 VSUBS 0.396535f
C1569 VDD2.n0 VSUBS 4.19769f
C1570 VDD2.t2 VSUBS 0.396535f
C1571 VDD2.t0 VSUBS 0.396535f
C1572 VDD2.n1 VSUBS 3.29851f
C1573 VDD2.n2 VSUBS 4.71698f
C1574 VN.t2 VSUBS 2.4473f
C1575 VN.t3 VSUBS 2.44714f
C1576 VN.n0 VSUBS 1.75748f
C1577 VN.t1 VSUBS 2.4473f
C1578 VN.t0 VSUBS 2.44714f
C1579 VN.n1 VSUBS 3.32312f
.ends

