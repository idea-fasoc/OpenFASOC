* NGSPICE file created from diff_pair_sample_1277.ext - technology: sky130A

.subckt diff_pair_sample_1277 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X1 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=3.54
X2 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X3 VTAIL.t3 VP.t1 VDD1.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X4 VDD2.t8 VN.t1 VTAIL.t19 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=3.54
X5 VDD2.t7 VN.t2 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=3.54
X6 VDD1.t7 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=3.54
X7 VDD1.t6 VP.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X8 VTAIL.t14 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X9 VTAIL.t1 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X10 VDD2.t5 VN.t4 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=3.54
X11 VTAIL.t13 VN.t5 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X12 VTAIL.t12 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X13 VDD2.t2 VN.t7 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X14 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=3.54
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=3.54
X16 VDD2.t1 VN.t8 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=3.54
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=3.54
X18 VTAIL.t10 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X19 VDD1.t4 VP.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=3.54
X20 VTAIL.t2 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X21 VTAIL.t4 VP.t7 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=3.54
X22 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=3.54
X23 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=3.54
R0 VN.n100 VN.n99 161.3
R1 VN.n98 VN.n52 161.3
R2 VN.n97 VN.n96 161.3
R3 VN.n95 VN.n53 161.3
R4 VN.n94 VN.n93 161.3
R5 VN.n92 VN.n54 161.3
R6 VN.n91 VN.n90 161.3
R7 VN.n89 VN.n55 161.3
R8 VN.n88 VN.n87 161.3
R9 VN.n86 VN.n56 161.3
R10 VN.n85 VN.n84 161.3
R11 VN.n83 VN.n58 161.3
R12 VN.n82 VN.n81 161.3
R13 VN.n80 VN.n59 161.3
R14 VN.n79 VN.n78 161.3
R15 VN.n77 VN.n60 161.3
R16 VN.n76 VN.n75 161.3
R17 VN.n74 VN.n61 161.3
R18 VN.n73 VN.n72 161.3
R19 VN.n71 VN.n62 161.3
R20 VN.n70 VN.n69 161.3
R21 VN.n68 VN.n63 161.3
R22 VN.n67 VN.n66 161.3
R23 VN.n49 VN.n48 161.3
R24 VN.n47 VN.n1 161.3
R25 VN.n46 VN.n45 161.3
R26 VN.n44 VN.n2 161.3
R27 VN.n43 VN.n42 161.3
R28 VN.n41 VN.n3 161.3
R29 VN.n40 VN.n39 161.3
R30 VN.n38 VN.n4 161.3
R31 VN.n37 VN.n36 161.3
R32 VN.n34 VN.n5 161.3
R33 VN.n33 VN.n32 161.3
R34 VN.n31 VN.n6 161.3
R35 VN.n30 VN.n29 161.3
R36 VN.n28 VN.n7 161.3
R37 VN.n27 VN.n26 161.3
R38 VN.n25 VN.n8 161.3
R39 VN.n24 VN.n23 161.3
R40 VN.n22 VN.n9 161.3
R41 VN.n21 VN.n20 161.3
R42 VN.n19 VN.n10 161.3
R43 VN.n18 VN.n17 161.3
R44 VN.n16 VN.n11 161.3
R45 VN.n15 VN.n14 161.3
R46 VN.n50 VN.n0 78.3232
R47 VN.n101 VN.n51 78.3232
R48 VN.n13 VN.n12 56.5559
R49 VN.n65 VN.n64 56.5559
R50 VN.n42 VN.n2 56.5193
R51 VN.n93 VN.n53 56.5193
R52 VN.n65 VN.t8 52.0972
R53 VN.n13 VN.t1 52.0972
R54 VN VN.n101 51.4791
R55 VN.n21 VN.n10 46.8066
R56 VN.n29 VN.n6 46.8066
R57 VN.n73 VN.n62 46.8066
R58 VN.n81 VN.n58 46.8066
R59 VN.n17 VN.n10 34.1802
R60 VN.n33 VN.n6 34.1802
R61 VN.n69 VN.n62 34.1802
R62 VN.n85 VN.n58 34.1802
R63 VN.n16 VN.n15 24.4675
R64 VN.n17 VN.n16 24.4675
R65 VN.n22 VN.n21 24.4675
R66 VN.n23 VN.n22 24.4675
R67 VN.n23 VN.n8 24.4675
R68 VN.n27 VN.n8 24.4675
R69 VN.n28 VN.n27 24.4675
R70 VN.n29 VN.n28 24.4675
R71 VN.n34 VN.n33 24.4675
R72 VN.n36 VN.n34 24.4675
R73 VN.n40 VN.n4 24.4675
R74 VN.n41 VN.n40 24.4675
R75 VN.n42 VN.n41 24.4675
R76 VN.n46 VN.n2 24.4675
R77 VN.n47 VN.n46 24.4675
R78 VN.n48 VN.n47 24.4675
R79 VN.n69 VN.n68 24.4675
R80 VN.n68 VN.n67 24.4675
R81 VN.n81 VN.n80 24.4675
R82 VN.n80 VN.n79 24.4675
R83 VN.n79 VN.n60 24.4675
R84 VN.n75 VN.n60 24.4675
R85 VN.n75 VN.n74 24.4675
R86 VN.n74 VN.n73 24.4675
R87 VN.n93 VN.n92 24.4675
R88 VN.n92 VN.n91 24.4675
R89 VN.n91 VN.n55 24.4675
R90 VN.n87 VN.n86 24.4675
R91 VN.n86 VN.n85 24.4675
R92 VN.n99 VN.n98 24.4675
R93 VN.n98 VN.n97 24.4675
R94 VN.n97 VN.n53 24.4675
R95 VN.n8 VN.t0 18.4499
R96 VN.n12 VN.t5 18.4499
R97 VN.n35 VN.t6 18.4499
R98 VN.n0 VN.t4 18.4499
R99 VN.n60 VN.t7 18.4499
R100 VN.n64 VN.t9 18.4499
R101 VN.n57 VN.t3 18.4499
R102 VN.n51 VN.t2 18.4499
R103 VN.n15 VN.n12 18.1061
R104 VN.n36 VN.n35 18.1061
R105 VN.n67 VN.n64 18.1061
R106 VN.n87 VN.n57 18.1061
R107 VN.n48 VN.n0 11.7447
R108 VN.n99 VN.n51 11.7447
R109 VN.n35 VN.n4 6.36192
R110 VN.n57 VN.n55 6.36192
R111 VN.n66 VN.n65 3.10014
R112 VN.n14 VN.n13 3.10014
R113 VN.n101 VN.n100 0.354971
R114 VN.n50 VN.n49 0.354971
R115 VN VN.n50 0.26696
R116 VN.n100 VN.n52 0.189894
R117 VN.n96 VN.n52 0.189894
R118 VN.n96 VN.n95 0.189894
R119 VN.n95 VN.n94 0.189894
R120 VN.n94 VN.n54 0.189894
R121 VN.n90 VN.n54 0.189894
R122 VN.n90 VN.n89 0.189894
R123 VN.n89 VN.n88 0.189894
R124 VN.n88 VN.n56 0.189894
R125 VN.n84 VN.n56 0.189894
R126 VN.n84 VN.n83 0.189894
R127 VN.n83 VN.n82 0.189894
R128 VN.n82 VN.n59 0.189894
R129 VN.n78 VN.n59 0.189894
R130 VN.n78 VN.n77 0.189894
R131 VN.n77 VN.n76 0.189894
R132 VN.n76 VN.n61 0.189894
R133 VN.n72 VN.n61 0.189894
R134 VN.n72 VN.n71 0.189894
R135 VN.n71 VN.n70 0.189894
R136 VN.n70 VN.n63 0.189894
R137 VN.n66 VN.n63 0.189894
R138 VN.n14 VN.n11 0.189894
R139 VN.n18 VN.n11 0.189894
R140 VN.n19 VN.n18 0.189894
R141 VN.n20 VN.n19 0.189894
R142 VN.n20 VN.n9 0.189894
R143 VN.n24 VN.n9 0.189894
R144 VN.n25 VN.n24 0.189894
R145 VN.n26 VN.n25 0.189894
R146 VN.n26 VN.n7 0.189894
R147 VN.n30 VN.n7 0.189894
R148 VN.n31 VN.n30 0.189894
R149 VN.n32 VN.n31 0.189894
R150 VN.n32 VN.n5 0.189894
R151 VN.n37 VN.n5 0.189894
R152 VN.n38 VN.n37 0.189894
R153 VN.n39 VN.n38 0.189894
R154 VN.n39 VN.n3 0.189894
R155 VN.n43 VN.n3 0.189894
R156 VN.n44 VN.n43 0.189894
R157 VN.n45 VN.n44 0.189894
R158 VN.n45 VN.n1 0.189894
R159 VN.n49 VN.n1 0.189894
R160 VTAIL.n56 VTAIL.n50 289.615
R161 VTAIL.n8 VTAIL.n2 289.615
R162 VTAIL.n44 VTAIL.n38 289.615
R163 VTAIL.n28 VTAIL.n22 289.615
R164 VTAIL.n55 VTAIL.n54 185
R165 VTAIL.n57 VTAIL.n56 185
R166 VTAIL.n7 VTAIL.n6 185
R167 VTAIL.n9 VTAIL.n8 185
R168 VTAIL.n45 VTAIL.n44 185
R169 VTAIL.n43 VTAIL.n42 185
R170 VTAIL.n29 VTAIL.n28 185
R171 VTAIL.n27 VTAIL.n26 185
R172 VTAIL.n53 VTAIL.t17 153.582
R173 VTAIL.n5 VTAIL.t5 153.582
R174 VTAIL.n41 VTAIL.t6 153.582
R175 VTAIL.n25 VTAIL.t18 153.582
R176 VTAIL.n56 VTAIL.n55 104.615
R177 VTAIL.n8 VTAIL.n7 104.615
R178 VTAIL.n44 VTAIL.n43 104.615
R179 VTAIL.n28 VTAIL.n27 104.615
R180 VTAIL.n63 VTAIL.n62 68.7696
R181 VTAIL.n1 VTAIL.n0 68.7696
R182 VTAIL.n15 VTAIL.n14 68.7696
R183 VTAIL.n17 VTAIL.n16 68.7696
R184 VTAIL.n37 VTAIL.n36 68.7696
R185 VTAIL.n35 VTAIL.n34 68.7696
R186 VTAIL.n21 VTAIL.n20 68.7696
R187 VTAIL.n19 VTAIL.n18 68.7696
R188 VTAIL.n55 VTAIL.t17 52.3082
R189 VTAIL.n7 VTAIL.t5 52.3082
R190 VTAIL.n43 VTAIL.t6 52.3082
R191 VTAIL.n27 VTAIL.t18 52.3082
R192 VTAIL.n61 VTAIL.n60 31.2157
R193 VTAIL.n13 VTAIL.n12 31.2157
R194 VTAIL.n49 VTAIL.n48 31.2157
R195 VTAIL.n33 VTAIL.n32 31.2157
R196 VTAIL.n19 VTAIL.n17 21.3755
R197 VTAIL.n61 VTAIL.n49 18.0393
R198 VTAIL.n54 VTAIL.n53 10.1164
R199 VTAIL.n6 VTAIL.n5 10.1164
R200 VTAIL.n42 VTAIL.n41 10.1164
R201 VTAIL.n26 VTAIL.n25 10.1164
R202 VTAIL.n60 VTAIL.n59 9.45567
R203 VTAIL.n12 VTAIL.n11 9.45567
R204 VTAIL.n48 VTAIL.n47 9.45567
R205 VTAIL.n32 VTAIL.n31 9.45567
R206 VTAIL.n52 VTAIL.n51 9.3005
R207 VTAIL.n59 VTAIL.n58 9.3005
R208 VTAIL.n4 VTAIL.n3 9.3005
R209 VTAIL.n11 VTAIL.n10 9.3005
R210 VTAIL.n40 VTAIL.n39 9.3005
R211 VTAIL.n47 VTAIL.n46 9.3005
R212 VTAIL.n31 VTAIL.n30 9.3005
R213 VTAIL.n24 VTAIL.n23 9.3005
R214 VTAIL.n60 VTAIL.n50 8.92171
R215 VTAIL.n12 VTAIL.n2 8.92171
R216 VTAIL.n48 VTAIL.n38 8.92171
R217 VTAIL.n32 VTAIL.n22 8.92171
R218 VTAIL.n58 VTAIL.n57 8.14595
R219 VTAIL.n10 VTAIL.n9 8.14595
R220 VTAIL.n46 VTAIL.n45 8.14595
R221 VTAIL.n30 VTAIL.n29 8.14595
R222 VTAIL.n54 VTAIL.n52 7.3702
R223 VTAIL.n6 VTAIL.n4 7.3702
R224 VTAIL.n42 VTAIL.n40 7.3702
R225 VTAIL.n26 VTAIL.n24 7.3702
R226 VTAIL.n62 VTAIL.t16 7.30677
R227 VTAIL.n62 VTAIL.t12 7.30677
R228 VTAIL.n0 VTAIL.t19 7.30677
R229 VTAIL.n0 VTAIL.t13 7.30677
R230 VTAIL.n14 VTAIL.t7 7.30677
R231 VTAIL.n14 VTAIL.t2 7.30677
R232 VTAIL.n16 VTAIL.t8 7.30677
R233 VTAIL.n16 VTAIL.t1 7.30677
R234 VTAIL.n36 VTAIL.t9 7.30677
R235 VTAIL.n36 VTAIL.t3 7.30677
R236 VTAIL.n34 VTAIL.t0 7.30677
R237 VTAIL.n34 VTAIL.t4 7.30677
R238 VTAIL.n20 VTAIL.t11 7.30677
R239 VTAIL.n20 VTAIL.t10 7.30677
R240 VTAIL.n18 VTAIL.t15 7.30677
R241 VTAIL.n18 VTAIL.t14 7.30677
R242 VTAIL.n57 VTAIL.n52 5.81868
R243 VTAIL.n9 VTAIL.n4 5.81868
R244 VTAIL.n45 VTAIL.n40 5.81868
R245 VTAIL.n29 VTAIL.n24 5.81868
R246 VTAIL.n58 VTAIL.n50 5.04292
R247 VTAIL.n10 VTAIL.n2 5.04292
R248 VTAIL.n46 VTAIL.n38 5.04292
R249 VTAIL.n30 VTAIL.n22 5.04292
R250 VTAIL.n21 VTAIL.n19 3.33671
R251 VTAIL.n33 VTAIL.n21 3.33671
R252 VTAIL.n37 VTAIL.n35 3.33671
R253 VTAIL.n49 VTAIL.n37 3.33671
R254 VTAIL.n17 VTAIL.n15 3.33671
R255 VTAIL.n15 VTAIL.n13 3.33671
R256 VTAIL.n63 VTAIL.n61 3.33671
R257 VTAIL.n25 VTAIL.n23 3.00987
R258 VTAIL.n53 VTAIL.n51 3.00987
R259 VTAIL.n5 VTAIL.n3 3.00987
R260 VTAIL.n41 VTAIL.n39 3.00987
R261 VTAIL VTAIL.n1 2.56084
R262 VTAIL.n35 VTAIL.n33 2.13843
R263 VTAIL.n13 VTAIL.n1 2.13843
R264 VTAIL VTAIL.n63 0.776362
R265 VTAIL.n59 VTAIL.n51 0.155672
R266 VTAIL.n11 VTAIL.n3 0.155672
R267 VTAIL.n47 VTAIL.n39 0.155672
R268 VTAIL.n31 VTAIL.n23 0.155672
R269 VDD2.n21 VDD2.n15 289.615
R270 VDD2.n6 VDD2.n0 289.615
R271 VDD2.n22 VDD2.n21 185
R272 VDD2.n20 VDD2.n19 185
R273 VDD2.n5 VDD2.n4 185
R274 VDD2.n7 VDD2.n6 185
R275 VDD2.n3 VDD2.t8 153.582
R276 VDD2.n18 VDD2.t7 153.582
R277 VDD2.n21 VDD2.n20 104.615
R278 VDD2.n6 VDD2.n5 104.615
R279 VDD2.n14 VDD2.n13 87.8952
R280 VDD2 VDD2.n29 87.8924
R281 VDD2.n28 VDD2.n27 85.4484
R282 VDD2.n12 VDD2.n11 85.4484
R283 VDD2.n20 VDD2.t7 52.3082
R284 VDD2.n5 VDD2.t8 52.3082
R285 VDD2.n12 VDD2.n10 51.2306
R286 VDD2.n26 VDD2.n25 47.8944
R287 VDD2.n26 VDD2.n14 41.8985
R288 VDD2.n19 VDD2.n18 10.1164
R289 VDD2.n4 VDD2.n3 10.1164
R290 VDD2.n25 VDD2.n24 9.45567
R291 VDD2.n10 VDD2.n9 9.45567
R292 VDD2.n24 VDD2.n23 9.3005
R293 VDD2.n17 VDD2.n16 9.3005
R294 VDD2.n2 VDD2.n1 9.3005
R295 VDD2.n9 VDD2.n8 9.3005
R296 VDD2.n25 VDD2.n15 8.92171
R297 VDD2.n10 VDD2.n0 8.92171
R298 VDD2.n23 VDD2.n22 8.14595
R299 VDD2.n8 VDD2.n7 8.14595
R300 VDD2.n19 VDD2.n17 7.3702
R301 VDD2.n4 VDD2.n2 7.3702
R302 VDD2.n29 VDD2.t0 7.30677
R303 VDD2.n29 VDD2.t1 7.30677
R304 VDD2.n27 VDD2.t6 7.30677
R305 VDD2.n27 VDD2.t2 7.30677
R306 VDD2.n13 VDD2.t3 7.30677
R307 VDD2.n13 VDD2.t5 7.30677
R308 VDD2.n11 VDD2.t4 7.30677
R309 VDD2.n11 VDD2.t9 7.30677
R310 VDD2.n22 VDD2.n17 5.81868
R311 VDD2.n7 VDD2.n2 5.81868
R312 VDD2.n23 VDD2.n15 5.04292
R313 VDD2.n8 VDD2.n0 5.04292
R314 VDD2.n28 VDD2.n26 3.33671
R315 VDD2.n18 VDD2.n16 3.00987
R316 VDD2.n3 VDD2.n1 3.00987
R317 VDD2 VDD2.n28 0.892741
R318 VDD2.n14 VDD2.n12 0.779206
R319 VDD2.n24 VDD2.n16 0.155672
R320 VDD2.n9 VDD2.n1 0.155672
R321 B.n813 B.n812 585
R322 B.n235 B.n158 585
R323 B.n234 B.n233 585
R324 B.n232 B.n231 585
R325 B.n230 B.n229 585
R326 B.n228 B.n227 585
R327 B.n226 B.n225 585
R328 B.n224 B.n223 585
R329 B.n222 B.n221 585
R330 B.n220 B.n219 585
R331 B.n218 B.n217 585
R332 B.n216 B.n215 585
R333 B.n214 B.n213 585
R334 B.n212 B.n211 585
R335 B.n210 B.n209 585
R336 B.n208 B.n207 585
R337 B.n206 B.n205 585
R338 B.n204 B.n203 585
R339 B.n202 B.n201 585
R340 B.n200 B.n199 585
R341 B.n198 B.n197 585
R342 B.n196 B.n195 585
R343 B.n194 B.n193 585
R344 B.n192 B.n191 585
R345 B.n190 B.n189 585
R346 B.n188 B.n187 585
R347 B.n186 B.n185 585
R348 B.n184 B.n183 585
R349 B.n182 B.n181 585
R350 B.n180 B.n179 585
R351 B.n178 B.n177 585
R352 B.n176 B.n175 585
R353 B.n174 B.n173 585
R354 B.n172 B.n171 585
R355 B.n170 B.n169 585
R356 B.n168 B.n167 585
R357 B.n166 B.n165 585
R358 B.n138 B.n137 585
R359 B.n811 B.n139 585
R360 B.n816 B.n139 585
R361 B.n810 B.n809 585
R362 B.n809 B.n135 585
R363 B.n808 B.n134 585
R364 B.n822 B.n134 585
R365 B.n807 B.n133 585
R366 B.n823 B.n133 585
R367 B.n806 B.n132 585
R368 B.n824 B.n132 585
R369 B.n805 B.n804 585
R370 B.n804 B.n128 585
R371 B.n803 B.n127 585
R372 B.n830 B.n127 585
R373 B.n802 B.n126 585
R374 B.n831 B.n126 585
R375 B.n801 B.n125 585
R376 B.n832 B.n125 585
R377 B.n800 B.n799 585
R378 B.n799 B.n124 585
R379 B.n798 B.n120 585
R380 B.n838 B.n120 585
R381 B.n797 B.n119 585
R382 B.n839 B.n119 585
R383 B.n796 B.n118 585
R384 B.n840 B.n118 585
R385 B.n795 B.n794 585
R386 B.n794 B.n114 585
R387 B.n793 B.n113 585
R388 B.n846 B.n113 585
R389 B.n792 B.n112 585
R390 B.n847 B.n112 585
R391 B.n791 B.n111 585
R392 B.n848 B.n111 585
R393 B.n790 B.n789 585
R394 B.n789 B.n107 585
R395 B.n788 B.n106 585
R396 B.n854 B.n106 585
R397 B.n787 B.n105 585
R398 B.n855 B.n105 585
R399 B.n786 B.n104 585
R400 B.n856 B.n104 585
R401 B.n785 B.n784 585
R402 B.n784 B.n100 585
R403 B.n783 B.n99 585
R404 B.n862 B.n99 585
R405 B.n782 B.n98 585
R406 B.n863 B.n98 585
R407 B.n781 B.n97 585
R408 B.n864 B.n97 585
R409 B.n780 B.n779 585
R410 B.n779 B.n93 585
R411 B.n778 B.n92 585
R412 B.n870 B.n92 585
R413 B.n777 B.n91 585
R414 B.n871 B.n91 585
R415 B.n776 B.n90 585
R416 B.n872 B.n90 585
R417 B.n775 B.n774 585
R418 B.n774 B.n86 585
R419 B.n773 B.n85 585
R420 B.n878 B.n85 585
R421 B.n772 B.n84 585
R422 B.n879 B.n84 585
R423 B.n771 B.n83 585
R424 B.n880 B.n83 585
R425 B.n770 B.n769 585
R426 B.n769 B.n79 585
R427 B.n768 B.n78 585
R428 B.n886 B.n78 585
R429 B.n767 B.n77 585
R430 B.n887 B.n77 585
R431 B.n766 B.n76 585
R432 B.n888 B.n76 585
R433 B.n765 B.n764 585
R434 B.n764 B.n72 585
R435 B.n763 B.n71 585
R436 B.n894 B.n71 585
R437 B.n762 B.n70 585
R438 B.n895 B.n70 585
R439 B.n761 B.n69 585
R440 B.n896 B.n69 585
R441 B.n760 B.n759 585
R442 B.n759 B.n65 585
R443 B.n758 B.n64 585
R444 B.n902 B.n64 585
R445 B.n757 B.n63 585
R446 B.n903 B.n63 585
R447 B.n756 B.n62 585
R448 B.n904 B.n62 585
R449 B.n755 B.n754 585
R450 B.n754 B.n58 585
R451 B.n753 B.n57 585
R452 B.n910 B.n57 585
R453 B.n752 B.n56 585
R454 B.n911 B.n56 585
R455 B.n751 B.n55 585
R456 B.n912 B.n55 585
R457 B.n750 B.n749 585
R458 B.n749 B.n51 585
R459 B.n748 B.n50 585
R460 B.n918 B.n50 585
R461 B.n747 B.n49 585
R462 B.n919 B.n49 585
R463 B.n746 B.n48 585
R464 B.n920 B.n48 585
R465 B.n745 B.n744 585
R466 B.n744 B.n44 585
R467 B.n743 B.n43 585
R468 B.n926 B.n43 585
R469 B.n742 B.n42 585
R470 B.n927 B.n42 585
R471 B.n741 B.n41 585
R472 B.n928 B.n41 585
R473 B.n740 B.n739 585
R474 B.n739 B.n40 585
R475 B.n738 B.n36 585
R476 B.n934 B.n36 585
R477 B.n737 B.n35 585
R478 B.n935 B.n35 585
R479 B.n736 B.n34 585
R480 B.n936 B.n34 585
R481 B.n735 B.n734 585
R482 B.n734 B.n30 585
R483 B.n733 B.n29 585
R484 B.n942 B.n29 585
R485 B.n732 B.n28 585
R486 B.n943 B.n28 585
R487 B.n731 B.n27 585
R488 B.n944 B.n27 585
R489 B.n730 B.n729 585
R490 B.n729 B.n23 585
R491 B.n728 B.n22 585
R492 B.n950 B.n22 585
R493 B.n727 B.n21 585
R494 B.n951 B.n21 585
R495 B.n726 B.n20 585
R496 B.n952 B.n20 585
R497 B.n725 B.n724 585
R498 B.n724 B.n19 585
R499 B.n723 B.n15 585
R500 B.n958 B.n15 585
R501 B.n722 B.n14 585
R502 B.n959 B.n14 585
R503 B.n721 B.n13 585
R504 B.n960 B.n13 585
R505 B.n720 B.n719 585
R506 B.n719 B.n12 585
R507 B.n718 B.n717 585
R508 B.n718 B.n8 585
R509 B.n716 B.n7 585
R510 B.n967 B.n7 585
R511 B.n715 B.n6 585
R512 B.n968 B.n6 585
R513 B.n714 B.n5 585
R514 B.n969 B.n5 585
R515 B.n713 B.n712 585
R516 B.n712 B.n4 585
R517 B.n711 B.n236 585
R518 B.n711 B.n710 585
R519 B.n701 B.n237 585
R520 B.n238 B.n237 585
R521 B.n703 B.n702 585
R522 B.n704 B.n703 585
R523 B.n700 B.n243 585
R524 B.n243 B.n242 585
R525 B.n699 B.n698 585
R526 B.n698 B.n697 585
R527 B.n245 B.n244 585
R528 B.n690 B.n245 585
R529 B.n689 B.n688 585
R530 B.n691 B.n689 585
R531 B.n687 B.n250 585
R532 B.n250 B.n249 585
R533 B.n686 B.n685 585
R534 B.n685 B.n684 585
R535 B.n252 B.n251 585
R536 B.n253 B.n252 585
R537 B.n677 B.n676 585
R538 B.n678 B.n677 585
R539 B.n675 B.n258 585
R540 B.n258 B.n257 585
R541 B.n674 B.n673 585
R542 B.n673 B.n672 585
R543 B.n260 B.n259 585
R544 B.n261 B.n260 585
R545 B.n665 B.n664 585
R546 B.n666 B.n665 585
R547 B.n663 B.n266 585
R548 B.n266 B.n265 585
R549 B.n662 B.n661 585
R550 B.n661 B.n660 585
R551 B.n268 B.n267 585
R552 B.n653 B.n268 585
R553 B.n652 B.n651 585
R554 B.n654 B.n652 585
R555 B.n650 B.n273 585
R556 B.n273 B.n272 585
R557 B.n649 B.n648 585
R558 B.n648 B.n647 585
R559 B.n275 B.n274 585
R560 B.n276 B.n275 585
R561 B.n640 B.n639 585
R562 B.n641 B.n640 585
R563 B.n638 B.n281 585
R564 B.n281 B.n280 585
R565 B.n637 B.n636 585
R566 B.n636 B.n635 585
R567 B.n283 B.n282 585
R568 B.n284 B.n283 585
R569 B.n628 B.n627 585
R570 B.n629 B.n628 585
R571 B.n626 B.n289 585
R572 B.n289 B.n288 585
R573 B.n625 B.n624 585
R574 B.n624 B.n623 585
R575 B.n291 B.n290 585
R576 B.n292 B.n291 585
R577 B.n616 B.n615 585
R578 B.n617 B.n616 585
R579 B.n614 B.n297 585
R580 B.n297 B.n296 585
R581 B.n613 B.n612 585
R582 B.n612 B.n611 585
R583 B.n299 B.n298 585
R584 B.n300 B.n299 585
R585 B.n604 B.n603 585
R586 B.n605 B.n604 585
R587 B.n602 B.n305 585
R588 B.n305 B.n304 585
R589 B.n601 B.n600 585
R590 B.n600 B.n599 585
R591 B.n307 B.n306 585
R592 B.n308 B.n307 585
R593 B.n592 B.n591 585
R594 B.n593 B.n592 585
R595 B.n590 B.n312 585
R596 B.n316 B.n312 585
R597 B.n589 B.n588 585
R598 B.n588 B.n587 585
R599 B.n314 B.n313 585
R600 B.n315 B.n314 585
R601 B.n580 B.n579 585
R602 B.n581 B.n580 585
R603 B.n578 B.n321 585
R604 B.n321 B.n320 585
R605 B.n577 B.n576 585
R606 B.n576 B.n575 585
R607 B.n323 B.n322 585
R608 B.n324 B.n323 585
R609 B.n568 B.n567 585
R610 B.n569 B.n568 585
R611 B.n566 B.n329 585
R612 B.n329 B.n328 585
R613 B.n565 B.n564 585
R614 B.n564 B.n563 585
R615 B.n331 B.n330 585
R616 B.n332 B.n331 585
R617 B.n556 B.n555 585
R618 B.n557 B.n556 585
R619 B.n554 B.n336 585
R620 B.n340 B.n336 585
R621 B.n553 B.n552 585
R622 B.n552 B.n551 585
R623 B.n338 B.n337 585
R624 B.n339 B.n338 585
R625 B.n544 B.n543 585
R626 B.n545 B.n544 585
R627 B.n542 B.n345 585
R628 B.n345 B.n344 585
R629 B.n541 B.n540 585
R630 B.n540 B.n539 585
R631 B.n347 B.n346 585
R632 B.n348 B.n347 585
R633 B.n532 B.n531 585
R634 B.n533 B.n532 585
R635 B.n530 B.n353 585
R636 B.n353 B.n352 585
R637 B.n529 B.n528 585
R638 B.n528 B.n527 585
R639 B.n355 B.n354 585
R640 B.n356 B.n355 585
R641 B.n520 B.n519 585
R642 B.n521 B.n520 585
R643 B.n518 B.n361 585
R644 B.n361 B.n360 585
R645 B.n517 B.n516 585
R646 B.n516 B.n515 585
R647 B.n363 B.n362 585
R648 B.n508 B.n363 585
R649 B.n507 B.n506 585
R650 B.n509 B.n507 585
R651 B.n505 B.n368 585
R652 B.n368 B.n367 585
R653 B.n504 B.n503 585
R654 B.n503 B.n502 585
R655 B.n370 B.n369 585
R656 B.n371 B.n370 585
R657 B.n495 B.n494 585
R658 B.n496 B.n495 585
R659 B.n493 B.n376 585
R660 B.n376 B.n375 585
R661 B.n492 B.n491 585
R662 B.n491 B.n490 585
R663 B.n378 B.n377 585
R664 B.n379 B.n378 585
R665 B.n483 B.n482 585
R666 B.n484 B.n483 585
R667 B.n382 B.n381 585
R668 B.n407 B.n405 585
R669 B.n408 B.n404 585
R670 B.n408 B.n383 585
R671 B.n411 B.n410 585
R672 B.n412 B.n403 585
R673 B.n414 B.n413 585
R674 B.n416 B.n402 585
R675 B.n419 B.n418 585
R676 B.n420 B.n401 585
R677 B.n422 B.n421 585
R678 B.n424 B.n400 585
R679 B.n427 B.n426 585
R680 B.n428 B.n399 585
R681 B.n433 B.n432 585
R682 B.n435 B.n398 585
R683 B.n438 B.n437 585
R684 B.n439 B.n397 585
R685 B.n441 B.n440 585
R686 B.n443 B.n396 585
R687 B.n446 B.n445 585
R688 B.n447 B.n395 585
R689 B.n449 B.n448 585
R690 B.n451 B.n394 585
R691 B.n454 B.n453 585
R692 B.n456 B.n391 585
R693 B.n458 B.n457 585
R694 B.n460 B.n390 585
R695 B.n463 B.n462 585
R696 B.n464 B.n389 585
R697 B.n466 B.n465 585
R698 B.n468 B.n388 585
R699 B.n471 B.n470 585
R700 B.n472 B.n387 585
R701 B.n474 B.n473 585
R702 B.n476 B.n386 585
R703 B.n477 B.n385 585
R704 B.n480 B.n479 585
R705 B.n481 B.n384 585
R706 B.n384 B.n383 585
R707 B.n486 B.n485 585
R708 B.n485 B.n484 585
R709 B.n487 B.n380 585
R710 B.n380 B.n379 585
R711 B.n489 B.n488 585
R712 B.n490 B.n489 585
R713 B.n374 B.n373 585
R714 B.n375 B.n374 585
R715 B.n498 B.n497 585
R716 B.n497 B.n496 585
R717 B.n499 B.n372 585
R718 B.n372 B.n371 585
R719 B.n501 B.n500 585
R720 B.n502 B.n501 585
R721 B.n366 B.n365 585
R722 B.n367 B.n366 585
R723 B.n511 B.n510 585
R724 B.n510 B.n509 585
R725 B.n512 B.n364 585
R726 B.n508 B.n364 585
R727 B.n514 B.n513 585
R728 B.n515 B.n514 585
R729 B.n359 B.n358 585
R730 B.n360 B.n359 585
R731 B.n523 B.n522 585
R732 B.n522 B.n521 585
R733 B.n524 B.n357 585
R734 B.n357 B.n356 585
R735 B.n526 B.n525 585
R736 B.n527 B.n526 585
R737 B.n351 B.n350 585
R738 B.n352 B.n351 585
R739 B.n535 B.n534 585
R740 B.n534 B.n533 585
R741 B.n536 B.n349 585
R742 B.n349 B.n348 585
R743 B.n538 B.n537 585
R744 B.n539 B.n538 585
R745 B.n343 B.n342 585
R746 B.n344 B.n343 585
R747 B.n547 B.n546 585
R748 B.n546 B.n545 585
R749 B.n548 B.n341 585
R750 B.n341 B.n339 585
R751 B.n550 B.n549 585
R752 B.n551 B.n550 585
R753 B.n335 B.n334 585
R754 B.n340 B.n335 585
R755 B.n559 B.n558 585
R756 B.n558 B.n557 585
R757 B.n560 B.n333 585
R758 B.n333 B.n332 585
R759 B.n562 B.n561 585
R760 B.n563 B.n562 585
R761 B.n327 B.n326 585
R762 B.n328 B.n327 585
R763 B.n571 B.n570 585
R764 B.n570 B.n569 585
R765 B.n572 B.n325 585
R766 B.n325 B.n324 585
R767 B.n574 B.n573 585
R768 B.n575 B.n574 585
R769 B.n319 B.n318 585
R770 B.n320 B.n319 585
R771 B.n583 B.n582 585
R772 B.n582 B.n581 585
R773 B.n584 B.n317 585
R774 B.n317 B.n315 585
R775 B.n586 B.n585 585
R776 B.n587 B.n586 585
R777 B.n311 B.n310 585
R778 B.n316 B.n311 585
R779 B.n595 B.n594 585
R780 B.n594 B.n593 585
R781 B.n596 B.n309 585
R782 B.n309 B.n308 585
R783 B.n598 B.n597 585
R784 B.n599 B.n598 585
R785 B.n303 B.n302 585
R786 B.n304 B.n303 585
R787 B.n607 B.n606 585
R788 B.n606 B.n605 585
R789 B.n608 B.n301 585
R790 B.n301 B.n300 585
R791 B.n610 B.n609 585
R792 B.n611 B.n610 585
R793 B.n295 B.n294 585
R794 B.n296 B.n295 585
R795 B.n619 B.n618 585
R796 B.n618 B.n617 585
R797 B.n620 B.n293 585
R798 B.n293 B.n292 585
R799 B.n622 B.n621 585
R800 B.n623 B.n622 585
R801 B.n287 B.n286 585
R802 B.n288 B.n287 585
R803 B.n631 B.n630 585
R804 B.n630 B.n629 585
R805 B.n632 B.n285 585
R806 B.n285 B.n284 585
R807 B.n634 B.n633 585
R808 B.n635 B.n634 585
R809 B.n279 B.n278 585
R810 B.n280 B.n279 585
R811 B.n643 B.n642 585
R812 B.n642 B.n641 585
R813 B.n644 B.n277 585
R814 B.n277 B.n276 585
R815 B.n646 B.n645 585
R816 B.n647 B.n646 585
R817 B.n271 B.n270 585
R818 B.n272 B.n271 585
R819 B.n656 B.n655 585
R820 B.n655 B.n654 585
R821 B.n657 B.n269 585
R822 B.n653 B.n269 585
R823 B.n659 B.n658 585
R824 B.n660 B.n659 585
R825 B.n264 B.n263 585
R826 B.n265 B.n264 585
R827 B.n668 B.n667 585
R828 B.n667 B.n666 585
R829 B.n669 B.n262 585
R830 B.n262 B.n261 585
R831 B.n671 B.n670 585
R832 B.n672 B.n671 585
R833 B.n256 B.n255 585
R834 B.n257 B.n256 585
R835 B.n680 B.n679 585
R836 B.n679 B.n678 585
R837 B.n681 B.n254 585
R838 B.n254 B.n253 585
R839 B.n683 B.n682 585
R840 B.n684 B.n683 585
R841 B.n248 B.n247 585
R842 B.n249 B.n248 585
R843 B.n693 B.n692 585
R844 B.n692 B.n691 585
R845 B.n694 B.n246 585
R846 B.n690 B.n246 585
R847 B.n696 B.n695 585
R848 B.n697 B.n696 585
R849 B.n241 B.n240 585
R850 B.n242 B.n241 585
R851 B.n706 B.n705 585
R852 B.n705 B.n704 585
R853 B.n707 B.n239 585
R854 B.n239 B.n238 585
R855 B.n709 B.n708 585
R856 B.n710 B.n709 585
R857 B.n3 B.n0 585
R858 B.n4 B.n3 585
R859 B.n966 B.n1 585
R860 B.n967 B.n966 585
R861 B.n965 B.n964 585
R862 B.n965 B.n8 585
R863 B.n963 B.n9 585
R864 B.n12 B.n9 585
R865 B.n962 B.n961 585
R866 B.n961 B.n960 585
R867 B.n11 B.n10 585
R868 B.n959 B.n11 585
R869 B.n957 B.n956 585
R870 B.n958 B.n957 585
R871 B.n955 B.n16 585
R872 B.n19 B.n16 585
R873 B.n954 B.n953 585
R874 B.n953 B.n952 585
R875 B.n18 B.n17 585
R876 B.n951 B.n18 585
R877 B.n949 B.n948 585
R878 B.n950 B.n949 585
R879 B.n947 B.n24 585
R880 B.n24 B.n23 585
R881 B.n946 B.n945 585
R882 B.n945 B.n944 585
R883 B.n26 B.n25 585
R884 B.n943 B.n26 585
R885 B.n941 B.n940 585
R886 B.n942 B.n941 585
R887 B.n939 B.n31 585
R888 B.n31 B.n30 585
R889 B.n938 B.n937 585
R890 B.n937 B.n936 585
R891 B.n33 B.n32 585
R892 B.n935 B.n33 585
R893 B.n933 B.n932 585
R894 B.n934 B.n933 585
R895 B.n931 B.n37 585
R896 B.n40 B.n37 585
R897 B.n930 B.n929 585
R898 B.n929 B.n928 585
R899 B.n39 B.n38 585
R900 B.n927 B.n39 585
R901 B.n925 B.n924 585
R902 B.n926 B.n925 585
R903 B.n923 B.n45 585
R904 B.n45 B.n44 585
R905 B.n922 B.n921 585
R906 B.n921 B.n920 585
R907 B.n47 B.n46 585
R908 B.n919 B.n47 585
R909 B.n917 B.n916 585
R910 B.n918 B.n917 585
R911 B.n915 B.n52 585
R912 B.n52 B.n51 585
R913 B.n914 B.n913 585
R914 B.n913 B.n912 585
R915 B.n54 B.n53 585
R916 B.n911 B.n54 585
R917 B.n909 B.n908 585
R918 B.n910 B.n909 585
R919 B.n907 B.n59 585
R920 B.n59 B.n58 585
R921 B.n906 B.n905 585
R922 B.n905 B.n904 585
R923 B.n61 B.n60 585
R924 B.n903 B.n61 585
R925 B.n901 B.n900 585
R926 B.n902 B.n901 585
R927 B.n899 B.n66 585
R928 B.n66 B.n65 585
R929 B.n898 B.n897 585
R930 B.n897 B.n896 585
R931 B.n68 B.n67 585
R932 B.n895 B.n68 585
R933 B.n893 B.n892 585
R934 B.n894 B.n893 585
R935 B.n891 B.n73 585
R936 B.n73 B.n72 585
R937 B.n890 B.n889 585
R938 B.n889 B.n888 585
R939 B.n75 B.n74 585
R940 B.n887 B.n75 585
R941 B.n885 B.n884 585
R942 B.n886 B.n885 585
R943 B.n883 B.n80 585
R944 B.n80 B.n79 585
R945 B.n882 B.n881 585
R946 B.n881 B.n880 585
R947 B.n82 B.n81 585
R948 B.n879 B.n82 585
R949 B.n877 B.n876 585
R950 B.n878 B.n877 585
R951 B.n875 B.n87 585
R952 B.n87 B.n86 585
R953 B.n874 B.n873 585
R954 B.n873 B.n872 585
R955 B.n89 B.n88 585
R956 B.n871 B.n89 585
R957 B.n869 B.n868 585
R958 B.n870 B.n869 585
R959 B.n867 B.n94 585
R960 B.n94 B.n93 585
R961 B.n866 B.n865 585
R962 B.n865 B.n864 585
R963 B.n96 B.n95 585
R964 B.n863 B.n96 585
R965 B.n861 B.n860 585
R966 B.n862 B.n861 585
R967 B.n859 B.n101 585
R968 B.n101 B.n100 585
R969 B.n858 B.n857 585
R970 B.n857 B.n856 585
R971 B.n103 B.n102 585
R972 B.n855 B.n103 585
R973 B.n853 B.n852 585
R974 B.n854 B.n853 585
R975 B.n851 B.n108 585
R976 B.n108 B.n107 585
R977 B.n850 B.n849 585
R978 B.n849 B.n848 585
R979 B.n110 B.n109 585
R980 B.n847 B.n110 585
R981 B.n845 B.n844 585
R982 B.n846 B.n845 585
R983 B.n843 B.n115 585
R984 B.n115 B.n114 585
R985 B.n842 B.n841 585
R986 B.n841 B.n840 585
R987 B.n117 B.n116 585
R988 B.n839 B.n117 585
R989 B.n837 B.n836 585
R990 B.n838 B.n837 585
R991 B.n835 B.n121 585
R992 B.n124 B.n121 585
R993 B.n834 B.n833 585
R994 B.n833 B.n832 585
R995 B.n123 B.n122 585
R996 B.n831 B.n123 585
R997 B.n829 B.n828 585
R998 B.n830 B.n829 585
R999 B.n827 B.n129 585
R1000 B.n129 B.n128 585
R1001 B.n826 B.n825 585
R1002 B.n825 B.n824 585
R1003 B.n131 B.n130 585
R1004 B.n823 B.n131 585
R1005 B.n821 B.n820 585
R1006 B.n822 B.n821 585
R1007 B.n819 B.n136 585
R1008 B.n136 B.n135 585
R1009 B.n818 B.n817 585
R1010 B.n817 B.n816 585
R1011 B.n970 B.n969 585
R1012 B.n968 B.n2 585
R1013 B.n817 B.n138 497.305
R1014 B.n813 B.n139 497.305
R1015 B.n483 B.n384 497.305
R1016 B.n485 B.n382 497.305
R1017 B.n815 B.n814 256.663
R1018 B.n815 B.n157 256.663
R1019 B.n815 B.n156 256.663
R1020 B.n815 B.n155 256.663
R1021 B.n815 B.n154 256.663
R1022 B.n815 B.n153 256.663
R1023 B.n815 B.n152 256.663
R1024 B.n815 B.n151 256.663
R1025 B.n815 B.n150 256.663
R1026 B.n815 B.n149 256.663
R1027 B.n815 B.n148 256.663
R1028 B.n815 B.n147 256.663
R1029 B.n815 B.n146 256.663
R1030 B.n815 B.n145 256.663
R1031 B.n815 B.n144 256.663
R1032 B.n815 B.n143 256.663
R1033 B.n815 B.n142 256.663
R1034 B.n815 B.n141 256.663
R1035 B.n815 B.n140 256.663
R1036 B.n406 B.n383 256.663
R1037 B.n409 B.n383 256.663
R1038 B.n415 B.n383 256.663
R1039 B.n417 B.n383 256.663
R1040 B.n423 B.n383 256.663
R1041 B.n425 B.n383 256.663
R1042 B.n434 B.n383 256.663
R1043 B.n436 B.n383 256.663
R1044 B.n442 B.n383 256.663
R1045 B.n444 B.n383 256.663
R1046 B.n450 B.n383 256.663
R1047 B.n452 B.n383 256.663
R1048 B.n459 B.n383 256.663
R1049 B.n461 B.n383 256.663
R1050 B.n467 B.n383 256.663
R1051 B.n469 B.n383 256.663
R1052 B.n475 B.n383 256.663
R1053 B.n478 B.n383 256.663
R1054 B.n972 B.n971 256.663
R1055 B.n162 B.t14 227.578
R1056 B.n159 B.t21 227.578
R1057 B.n392 B.t10 227.578
R1058 B.n429 B.t18 227.578
R1059 B.n159 B.t22 201.827
R1060 B.n392 B.t13 201.827
R1061 B.n162 B.t16 201.827
R1062 B.n429 B.t20 201.827
R1063 B.n167 B.n166 163.367
R1064 B.n171 B.n170 163.367
R1065 B.n175 B.n174 163.367
R1066 B.n179 B.n178 163.367
R1067 B.n183 B.n182 163.367
R1068 B.n187 B.n186 163.367
R1069 B.n191 B.n190 163.367
R1070 B.n195 B.n194 163.367
R1071 B.n199 B.n198 163.367
R1072 B.n203 B.n202 163.367
R1073 B.n207 B.n206 163.367
R1074 B.n211 B.n210 163.367
R1075 B.n215 B.n214 163.367
R1076 B.n219 B.n218 163.367
R1077 B.n223 B.n222 163.367
R1078 B.n227 B.n226 163.367
R1079 B.n231 B.n230 163.367
R1080 B.n233 B.n158 163.367
R1081 B.n483 B.n378 163.367
R1082 B.n491 B.n378 163.367
R1083 B.n491 B.n376 163.367
R1084 B.n495 B.n376 163.367
R1085 B.n495 B.n370 163.367
R1086 B.n503 B.n370 163.367
R1087 B.n503 B.n368 163.367
R1088 B.n507 B.n368 163.367
R1089 B.n507 B.n363 163.367
R1090 B.n516 B.n363 163.367
R1091 B.n516 B.n361 163.367
R1092 B.n520 B.n361 163.367
R1093 B.n520 B.n355 163.367
R1094 B.n528 B.n355 163.367
R1095 B.n528 B.n353 163.367
R1096 B.n532 B.n353 163.367
R1097 B.n532 B.n347 163.367
R1098 B.n540 B.n347 163.367
R1099 B.n540 B.n345 163.367
R1100 B.n544 B.n345 163.367
R1101 B.n544 B.n338 163.367
R1102 B.n552 B.n338 163.367
R1103 B.n552 B.n336 163.367
R1104 B.n556 B.n336 163.367
R1105 B.n556 B.n331 163.367
R1106 B.n564 B.n331 163.367
R1107 B.n564 B.n329 163.367
R1108 B.n568 B.n329 163.367
R1109 B.n568 B.n323 163.367
R1110 B.n576 B.n323 163.367
R1111 B.n576 B.n321 163.367
R1112 B.n580 B.n321 163.367
R1113 B.n580 B.n314 163.367
R1114 B.n588 B.n314 163.367
R1115 B.n588 B.n312 163.367
R1116 B.n592 B.n312 163.367
R1117 B.n592 B.n307 163.367
R1118 B.n600 B.n307 163.367
R1119 B.n600 B.n305 163.367
R1120 B.n604 B.n305 163.367
R1121 B.n604 B.n299 163.367
R1122 B.n612 B.n299 163.367
R1123 B.n612 B.n297 163.367
R1124 B.n616 B.n297 163.367
R1125 B.n616 B.n291 163.367
R1126 B.n624 B.n291 163.367
R1127 B.n624 B.n289 163.367
R1128 B.n628 B.n289 163.367
R1129 B.n628 B.n283 163.367
R1130 B.n636 B.n283 163.367
R1131 B.n636 B.n281 163.367
R1132 B.n640 B.n281 163.367
R1133 B.n640 B.n275 163.367
R1134 B.n648 B.n275 163.367
R1135 B.n648 B.n273 163.367
R1136 B.n652 B.n273 163.367
R1137 B.n652 B.n268 163.367
R1138 B.n661 B.n268 163.367
R1139 B.n661 B.n266 163.367
R1140 B.n665 B.n266 163.367
R1141 B.n665 B.n260 163.367
R1142 B.n673 B.n260 163.367
R1143 B.n673 B.n258 163.367
R1144 B.n677 B.n258 163.367
R1145 B.n677 B.n252 163.367
R1146 B.n685 B.n252 163.367
R1147 B.n685 B.n250 163.367
R1148 B.n689 B.n250 163.367
R1149 B.n689 B.n245 163.367
R1150 B.n698 B.n245 163.367
R1151 B.n698 B.n243 163.367
R1152 B.n703 B.n243 163.367
R1153 B.n703 B.n237 163.367
R1154 B.n711 B.n237 163.367
R1155 B.n712 B.n711 163.367
R1156 B.n712 B.n5 163.367
R1157 B.n6 B.n5 163.367
R1158 B.n7 B.n6 163.367
R1159 B.n718 B.n7 163.367
R1160 B.n719 B.n718 163.367
R1161 B.n719 B.n13 163.367
R1162 B.n14 B.n13 163.367
R1163 B.n15 B.n14 163.367
R1164 B.n724 B.n15 163.367
R1165 B.n724 B.n20 163.367
R1166 B.n21 B.n20 163.367
R1167 B.n22 B.n21 163.367
R1168 B.n729 B.n22 163.367
R1169 B.n729 B.n27 163.367
R1170 B.n28 B.n27 163.367
R1171 B.n29 B.n28 163.367
R1172 B.n734 B.n29 163.367
R1173 B.n734 B.n34 163.367
R1174 B.n35 B.n34 163.367
R1175 B.n36 B.n35 163.367
R1176 B.n739 B.n36 163.367
R1177 B.n739 B.n41 163.367
R1178 B.n42 B.n41 163.367
R1179 B.n43 B.n42 163.367
R1180 B.n744 B.n43 163.367
R1181 B.n744 B.n48 163.367
R1182 B.n49 B.n48 163.367
R1183 B.n50 B.n49 163.367
R1184 B.n749 B.n50 163.367
R1185 B.n749 B.n55 163.367
R1186 B.n56 B.n55 163.367
R1187 B.n57 B.n56 163.367
R1188 B.n754 B.n57 163.367
R1189 B.n754 B.n62 163.367
R1190 B.n63 B.n62 163.367
R1191 B.n64 B.n63 163.367
R1192 B.n759 B.n64 163.367
R1193 B.n759 B.n69 163.367
R1194 B.n70 B.n69 163.367
R1195 B.n71 B.n70 163.367
R1196 B.n764 B.n71 163.367
R1197 B.n764 B.n76 163.367
R1198 B.n77 B.n76 163.367
R1199 B.n78 B.n77 163.367
R1200 B.n769 B.n78 163.367
R1201 B.n769 B.n83 163.367
R1202 B.n84 B.n83 163.367
R1203 B.n85 B.n84 163.367
R1204 B.n774 B.n85 163.367
R1205 B.n774 B.n90 163.367
R1206 B.n91 B.n90 163.367
R1207 B.n92 B.n91 163.367
R1208 B.n779 B.n92 163.367
R1209 B.n779 B.n97 163.367
R1210 B.n98 B.n97 163.367
R1211 B.n99 B.n98 163.367
R1212 B.n784 B.n99 163.367
R1213 B.n784 B.n104 163.367
R1214 B.n105 B.n104 163.367
R1215 B.n106 B.n105 163.367
R1216 B.n789 B.n106 163.367
R1217 B.n789 B.n111 163.367
R1218 B.n112 B.n111 163.367
R1219 B.n113 B.n112 163.367
R1220 B.n794 B.n113 163.367
R1221 B.n794 B.n118 163.367
R1222 B.n119 B.n118 163.367
R1223 B.n120 B.n119 163.367
R1224 B.n799 B.n120 163.367
R1225 B.n799 B.n125 163.367
R1226 B.n126 B.n125 163.367
R1227 B.n127 B.n126 163.367
R1228 B.n804 B.n127 163.367
R1229 B.n804 B.n132 163.367
R1230 B.n133 B.n132 163.367
R1231 B.n134 B.n133 163.367
R1232 B.n809 B.n134 163.367
R1233 B.n809 B.n139 163.367
R1234 B.n408 B.n407 163.367
R1235 B.n410 B.n408 163.367
R1236 B.n414 B.n403 163.367
R1237 B.n418 B.n416 163.367
R1238 B.n422 B.n401 163.367
R1239 B.n426 B.n424 163.367
R1240 B.n433 B.n399 163.367
R1241 B.n437 B.n435 163.367
R1242 B.n441 B.n397 163.367
R1243 B.n445 B.n443 163.367
R1244 B.n449 B.n395 163.367
R1245 B.n453 B.n451 163.367
R1246 B.n458 B.n391 163.367
R1247 B.n462 B.n460 163.367
R1248 B.n466 B.n389 163.367
R1249 B.n470 B.n468 163.367
R1250 B.n474 B.n387 163.367
R1251 B.n477 B.n476 163.367
R1252 B.n479 B.n384 163.367
R1253 B.n485 B.n380 163.367
R1254 B.n489 B.n380 163.367
R1255 B.n489 B.n374 163.367
R1256 B.n497 B.n374 163.367
R1257 B.n497 B.n372 163.367
R1258 B.n501 B.n372 163.367
R1259 B.n501 B.n366 163.367
R1260 B.n510 B.n366 163.367
R1261 B.n510 B.n364 163.367
R1262 B.n514 B.n364 163.367
R1263 B.n514 B.n359 163.367
R1264 B.n522 B.n359 163.367
R1265 B.n522 B.n357 163.367
R1266 B.n526 B.n357 163.367
R1267 B.n526 B.n351 163.367
R1268 B.n534 B.n351 163.367
R1269 B.n534 B.n349 163.367
R1270 B.n538 B.n349 163.367
R1271 B.n538 B.n343 163.367
R1272 B.n546 B.n343 163.367
R1273 B.n546 B.n341 163.367
R1274 B.n550 B.n341 163.367
R1275 B.n550 B.n335 163.367
R1276 B.n558 B.n335 163.367
R1277 B.n558 B.n333 163.367
R1278 B.n562 B.n333 163.367
R1279 B.n562 B.n327 163.367
R1280 B.n570 B.n327 163.367
R1281 B.n570 B.n325 163.367
R1282 B.n574 B.n325 163.367
R1283 B.n574 B.n319 163.367
R1284 B.n582 B.n319 163.367
R1285 B.n582 B.n317 163.367
R1286 B.n586 B.n317 163.367
R1287 B.n586 B.n311 163.367
R1288 B.n594 B.n311 163.367
R1289 B.n594 B.n309 163.367
R1290 B.n598 B.n309 163.367
R1291 B.n598 B.n303 163.367
R1292 B.n606 B.n303 163.367
R1293 B.n606 B.n301 163.367
R1294 B.n610 B.n301 163.367
R1295 B.n610 B.n295 163.367
R1296 B.n618 B.n295 163.367
R1297 B.n618 B.n293 163.367
R1298 B.n622 B.n293 163.367
R1299 B.n622 B.n287 163.367
R1300 B.n630 B.n287 163.367
R1301 B.n630 B.n285 163.367
R1302 B.n634 B.n285 163.367
R1303 B.n634 B.n279 163.367
R1304 B.n642 B.n279 163.367
R1305 B.n642 B.n277 163.367
R1306 B.n646 B.n277 163.367
R1307 B.n646 B.n271 163.367
R1308 B.n655 B.n271 163.367
R1309 B.n655 B.n269 163.367
R1310 B.n659 B.n269 163.367
R1311 B.n659 B.n264 163.367
R1312 B.n667 B.n264 163.367
R1313 B.n667 B.n262 163.367
R1314 B.n671 B.n262 163.367
R1315 B.n671 B.n256 163.367
R1316 B.n679 B.n256 163.367
R1317 B.n679 B.n254 163.367
R1318 B.n683 B.n254 163.367
R1319 B.n683 B.n248 163.367
R1320 B.n692 B.n248 163.367
R1321 B.n692 B.n246 163.367
R1322 B.n696 B.n246 163.367
R1323 B.n696 B.n241 163.367
R1324 B.n705 B.n241 163.367
R1325 B.n705 B.n239 163.367
R1326 B.n709 B.n239 163.367
R1327 B.n709 B.n3 163.367
R1328 B.n970 B.n3 163.367
R1329 B.n966 B.n2 163.367
R1330 B.n966 B.n965 163.367
R1331 B.n965 B.n9 163.367
R1332 B.n961 B.n9 163.367
R1333 B.n961 B.n11 163.367
R1334 B.n957 B.n11 163.367
R1335 B.n957 B.n16 163.367
R1336 B.n953 B.n16 163.367
R1337 B.n953 B.n18 163.367
R1338 B.n949 B.n18 163.367
R1339 B.n949 B.n24 163.367
R1340 B.n945 B.n24 163.367
R1341 B.n945 B.n26 163.367
R1342 B.n941 B.n26 163.367
R1343 B.n941 B.n31 163.367
R1344 B.n937 B.n31 163.367
R1345 B.n937 B.n33 163.367
R1346 B.n933 B.n33 163.367
R1347 B.n933 B.n37 163.367
R1348 B.n929 B.n37 163.367
R1349 B.n929 B.n39 163.367
R1350 B.n925 B.n39 163.367
R1351 B.n925 B.n45 163.367
R1352 B.n921 B.n45 163.367
R1353 B.n921 B.n47 163.367
R1354 B.n917 B.n47 163.367
R1355 B.n917 B.n52 163.367
R1356 B.n913 B.n52 163.367
R1357 B.n913 B.n54 163.367
R1358 B.n909 B.n54 163.367
R1359 B.n909 B.n59 163.367
R1360 B.n905 B.n59 163.367
R1361 B.n905 B.n61 163.367
R1362 B.n901 B.n61 163.367
R1363 B.n901 B.n66 163.367
R1364 B.n897 B.n66 163.367
R1365 B.n897 B.n68 163.367
R1366 B.n893 B.n68 163.367
R1367 B.n893 B.n73 163.367
R1368 B.n889 B.n73 163.367
R1369 B.n889 B.n75 163.367
R1370 B.n885 B.n75 163.367
R1371 B.n885 B.n80 163.367
R1372 B.n881 B.n80 163.367
R1373 B.n881 B.n82 163.367
R1374 B.n877 B.n82 163.367
R1375 B.n877 B.n87 163.367
R1376 B.n873 B.n87 163.367
R1377 B.n873 B.n89 163.367
R1378 B.n869 B.n89 163.367
R1379 B.n869 B.n94 163.367
R1380 B.n865 B.n94 163.367
R1381 B.n865 B.n96 163.367
R1382 B.n861 B.n96 163.367
R1383 B.n861 B.n101 163.367
R1384 B.n857 B.n101 163.367
R1385 B.n857 B.n103 163.367
R1386 B.n853 B.n103 163.367
R1387 B.n853 B.n108 163.367
R1388 B.n849 B.n108 163.367
R1389 B.n849 B.n110 163.367
R1390 B.n845 B.n110 163.367
R1391 B.n845 B.n115 163.367
R1392 B.n841 B.n115 163.367
R1393 B.n841 B.n117 163.367
R1394 B.n837 B.n117 163.367
R1395 B.n837 B.n121 163.367
R1396 B.n833 B.n121 163.367
R1397 B.n833 B.n123 163.367
R1398 B.n829 B.n123 163.367
R1399 B.n829 B.n129 163.367
R1400 B.n825 B.n129 163.367
R1401 B.n825 B.n131 163.367
R1402 B.n821 B.n131 163.367
R1403 B.n821 B.n136 163.367
R1404 B.n817 B.n136 163.367
R1405 B.n484 B.n383 161.178
R1406 B.n816 B.n815 161.178
R1407 B.n160 B.t23 126.772
R1408 B.n393 B.t12 126.772
R1409 B.n163 B.t17 126.772
R1410 B.n430 B.t19 126.772
R1411 B.n484 B.n379 93.6761
R1412 B.n490 B.n379 93.6761
R1413 B.n490 B.n375 93.6761
R1414 B.n496 B.n375 93.6761
R1415 B.n496 B.n371 93.6761
R1416 B.n502 B.n371 93.6761
R1417 B.n502 B.n367 93.6761
R1418 B.n509 B.n367 93.6761
R1419 B.n509 B.n508 93.6761
R1420 B.n515 B.n360 93.6761
R1421 B.n521 B.n360 93.6761
R1422 B.n521 B.n356 93.6761
R1423 B.n527 B.n356 93.6761
R1424 B.n527 B.n352 93.6761
R1425 B.n533 B.n352 93.6761
R1426 B.n533 B.n348 93.6761
R1427 B.n539 B.n348 93.6761
R1428 B.n539 B.n344 93.6761
R1429 B.n545 B.n344 93.6761
R1430 B.n545 B.n339 93.6761
R1431 B.n551 B.n339 93.6761
R1432 B.n551 B.n340 93.6761
R1433 B.n557 B.n332 93.6761
R1434 B.n563 B.n332 93.6761
R1435 B.n563 B.n328 93.6761
R1436 B.n569 B.n328 93.6761
R1437 B.n569 B.n324 93.6761
R1438 B.n575 B.n324 93.6761
R1439 B.n575 B.n320 93.6761
R1440 B.n581 B.n320 93.6761
R1441 B.n581 B.n315 93.6761
R1442 B.n587 B.n315 93.6761
R1443 B.n587 B.n316 93.6761
R1444 B.n593 B.n308 93.6761
R1445 B.n599 B.n308 93.6761
R1446 B.n599 B.n304 93.6761
R1447 B.n605 B.n304 93.6761
R1448 B.n605 B.n300 93.6761
R1449 B.n611 B.n300 93.6761
R1450 B.n611 B.n296 93.6761
R1451 B.n617 B.n296 93.6761
R1452 B.n617 B.n292 93.6761
R1453 B.n623 B.n292 93.6761
R1454 B.n629 B.n288 93.6761
R1455 B.n629 B.n284 93.6761
R1456 B.n635 B.n284 93.6761
R1457 B.n635 B.n280 93.6761
R1458 B.n641 B.n280 93.6761
R1459 B.n641 B.n276 93.6761
R1460 B.n647 B.n276 93.6761
R1461 B.n647 B.n272 93.6761
R1462 B.n654 B.n272 93.6761
R1463 B.n654 B.n653 93.6761
R1464 B.n660 B.n265 93.6761
R1465 B.n666 B.n265 93.6761
R1466 B.n666 B.n261 93.6761
R1467 B.n672 B.n261 93.6761
R1468 B.n672 B.n257 93.6761
R1469 B.n678 B.n257 93.6761
R1470 B.n678 B.n253 93.6761
R1471 B.n684 B.n253 93.6761
R1472 B.n684 B.n249 93.6761
R1473 B.n691 B.n249 93.6761
R1474 B.n691 B.n690 93.6761
R1475 B.n697 B.n242 93.6761
R1476 B.n704 B.n242 93.6761
R1477 B.n704 B.n238 93.6761
R1478 B.n710 B.n238 93.6761
R1479 B.n710 B.n4 93.6761
R1480 B.n969 B.n4 93.6761
R1481 B.n969 B.n968 93.6761
R1482 B.n968 B.n967 93.6761
R1483 B.n967 B.n8 93.6761
R1484 B.n12 B.n8 93.6761
R1485 B.n960 B.n12 93.6761
R1486 B.n960 B.n959 93.6761
R1487 B.n959 B.n958 93.6761
R1488 B.n952 B.n19 93.6761
R1489 B.n952 B.n951 93.6761
R1490 B.n951 B.n950 93.6761
R1491 B.n950 B.n23 93.6761
R1492 B.n944 B.n23 93.6761
R1493 B.n944 B.n943 93.6761
R1494 B.n943 B.n942 93.6761
R1495 B.n942 B.n30 93.6761
R1496 B.n936 B.n30 93.6761
R1497 B.n936 B.n935 93.6761
R1498 B.n935 B.n934 93.6761
R1499 B.n928 B.n40 93.6761
R1500 B.n928 B.n927 93.6761
R1501 B.n927 B.n926 93.6761
R1502 B.n926 B.n44 93.6761
R1503 B.n920 B.n44 93.6761
R1504 B.n920 B.n919 93.6761
R1505 B.n919 B.n918 93.6761
R1506 B.n918 B.n51 93.6761
R1507 B.n912 B.n51 93.6761
R1508 B.n912 B.n911 93.6761
R1509 B.n910 B.n58 93.6761
R1510 B.n904 B.n58 93.6761
R1511 B.n904 B.n903 93.6761
R1512 B.n903 B.n902 93.6761
R1513 B.n902 B.n65 93.6761
R1514 B.n896 B.n65 93.6761
R1515 B.n896 B.n895 93.6761
R1516 B.n895 B.n894 93.6761
R1517 B.n894 B.n72 93.6761
R1518 B.n888 B.n72 93.6761
R1519 B.n887 B.n886 93.6761
R1520 B.n886 B.n79 93.6761
R1521 B.n880 B.n79 93.6761
R1522 B.n880 B.n879 93.6761
R1523 B.n879 B.n878 93.6761
R1524 B.n878 B.n86 93.6761
R1525 B.n872 B.n86 93.6761
R1526 B.n872 B.n871 93.6761
R1527 B.n871 B.n870 93.6761
R1528 B.n870 B.n93 93.6761
R1529 B.n864 B.n93 93.6761
R1530 B.n863 B.n862 93.6761
R1531 B.n862 B.n100 93.6761
R1532 B.n856 B.n100 93.6761
R1533 B.n856 B.n855 93.6761
R1534 B.n855 B.n854 93.6761
R1535 B.n854 B.n107 93.6761
R1536 B.n848 B.n107 93.6761
R1537 B.n848 B.n847 93.6761
R1538 B.n847 B.n846 93.6761
R1539 B.n846 B.n114 93.6761
R1540 B.n840 B.n114 93.6761
R1541 B.n840 B.n839 93.6761
R1542 B.n839 B.n838 93.6761
R1543 B.n832 B.n124 93.6761
R1544 B.n832 B.n831 93.6761
R1545 B.n831 B.n830 93.6761
R1546 B.n830 B.n128 93.6761
R1547 B.n824 B.n128 93.6761
R1548 B.n824 B.n823 93.6761
R1549 B.n823 B.n822 93.6761
R1550 B.n822 B.n135 93.6761
R1551 B.n816 B.n135 93.6761
R1552 B.n593 B.t1 88.1658
R1553 B.n888 B.t3 88.1658
R1554 B.n515 B.t11 85.4106
R1555 B.n838 B.t15 85.4106
R1556 B.n653 B.t2 77.1451
R1557 B.n40 B.t4 77.1451
R1558 B.n163 B.n162 75.0551
R1559 B.n160 B.n159 75.0551
R1560 B.n393 B.n392 75.0551
R1561 B.n430 B.n429 75.0551
R1562 B.n697 B.t5 74.39
R1563 B.n958 B.t0 74.39
R1564 B.n140 B.n138 71.676
R1565 B.n167 B.n141 71.676
R1566 B.n171 B.n142 71.676
R1567 B.n175 B.n143 71.676
R1568 B.n179 B.n144 71.676
R1569 B.n183 B.n145 71.676
R1570 B.n187 B.n146 71.676
R1571 B.n191 B.n147 71.676
R1572 B.n195 B.n148 71.676
R1573 B.n199 B.n149 71.676
R1574 B.n203 B.n150 71.676
R1575 B.n207 B.n151 71.676
R1576 B.n211 B.n152 71.676
R1577 B.n215 B.n153 71.676
R1578 B.n219 B.n154 71.676
R1579 B.n223 B.n155 71.676
R1580 B.n227 B.n156 71.676
R1581 B.n231 B.n157 71.676
R1582 B.n814 B.n158 71.676
R1583 B.n814 B.n813 71.676
R1584 B.n233 B.n157 71.676
R1585 B.n230 B.n156 71.676
R1586 B.n226 B.n155 71.676
R1587 B.n222 B.n154 71.676
R1588 B.n218 B.n153 71.676
R1589 B.n214 B.n152 71.676
R1590 B.n210 B.n151 71.676
R1591 B.n206 B.n150 71.676
R1592 B.n202 B.n149 71.676
R1593 B.n198 B.n148 71.676
R1594 B.n194 B.n147 71.676
R1595 B.n190 B.n146 71.676
R1596 B.n186 B.n145 71.676
R1597 B.n182 B.n144 71.676
R1598 B.n178 B.n143 71.676
R1599 B.n174 B.n142 71.676
R1600 B.n170 B.n141 71.676
R1601 B.n166 B.n140 71.676
R1602 B.n406 B.n382 71.676
R1603 B.n410 B.n409 71.676
R1604 B.n415 B.n414 71.676
R1605 B.n418 B.n417 71.676
R1606 B.n423 B.n422 71.676
R1607 B.n426 B.n425 71.676
R1608 B.n434 B.n433 71.676
R1609 B.n437 B.n436 71.676
R1610 B.n442 B.n441 71.676
R1611 B.n445 B.n444 71.676
R1612 B.n450 B.n449 71.676
R1613 B.n453 B.n452 71.676
R1614 B.n459 B.n458 71.676
R1615 B.n462 B.n461 71.676
R1616 B.n467 B.n466 71.676
R1617 B.n470 B.n469 71.676
R1618 B.n475 B.n474 71.676
R1619 B.n478 B.n477 71.676
R1620 B.n407 B.n406 71.676
R1621 B.n409 B.n403 71.676
R1622 B.n416 B.n415 71.676
R1623 B.n417 B.n401 71.676
R1624 B.n424 B.n423 71.676
R1625 B.n425 B.n399 71.676
R1626 B.n435 B.n434 71.676
R1627 B.n436 B.n397 71.676
R1628 B.n443 B.n442 71.676
R1629 B.n444 B.n395 71.676
R1630 B.n451 B.n450 71.676
R1631 B.n452 B.n391 71.676
R1632 B.n460 B.n459 71.676
R1633 B.n461 B.n389 71.676
R1634 B.n468 B.n467 71.676
R1635 B.n469 B.n387 71.676
R1636 B.n476 B.n475 71.676
R1637 B.n479 B.n478 71.676
R1638 B.n971 B.n970 71.676
R1639 B.n971 B.n2 71.676
R1640 B.n340 B.t8 63.3693
R1641 B.t6 B.n863 63.3693
R1642 B.n164 B.n163 59.5399
R1643 B.n161 B.n160 59.5399
R1644 B.n455 B.n393 59.5399
R1645 B.n431 B.n430 59.5399
R1646 B.t7 B.n288 52.3487
R1647 B.n911 B.t9 52.3487
R1648 B.n623 B.t7 41.328
R1649 B.t9 B.n910 41.328
R1650 B.n486 B.n381 32.3127
R1651 B.n482 B.n481 32.3127
R1652 B.n812 B.n811 32.3127
R1653 B.n818 B.n137 32.3127
R1654 B.n557 B.t8 30.3073
R1655 B.n864 B.t6 30.3073
R1656 B.n690 B.t5 19.2867
R1657 B.n19 B.t0 19.2867
R1658 B B.n972 18.0485
R1659 B.n660 B.t2 16.5315
R1660 B.n934 B.t4 16.5315
R1661 B.n487 B.n486 10.6151
R1662 B.n488 B.n487 10.6151
R1663 B.n488 B.n373 10.6151
R1664 B.n498 B.n373 10.6151
R1665 B.n499 B.n498 10.6151
R1666 B.n500 B.n499 10.6151
R1667 B.n500 B.n365 10.6151
R1668 B.n511 B.n365 10.6151
R1669 B.n512 B.n511 10.6151
R1670 B.n513 B.n512 10.6151
R1671 B.n513 B.n358 10.6151
R1672 B.n523 B.n358 10.6151
R1673 B.n524 B.n523 10.6151
R1674 B.n525 B.n524 10.6151
R1675 B.n525 B.n350 10.6151
R1676 B.n535 B.n350 10.6151
R1677 B.n536 B.n535 10.6151
R1678 B.n537 B.n536 10.6151
R1679 B.n537 B.n342 10.6151
R1680 B.n547 B.n342 10.6151
R1681 B.n548 B.n547 10.6151
R1682 B.n549 B.n548 10.6151
R1683 B.n549 B.n334 10.6151
R1684 B.n559 B.n334 10.6151
R1685 B.n560 B.n559 10.6151
R1686 B.n561 B.n560 10.6151
R1687 B.n561 B.n326 10.6151
R1688 B.n571 B.n326 10.6151
R1689 B.n572 B.n571 10.6151
R1690 B.n573 B.n572 10.6151
R1691 B.n573 B.n318 10.6151
R1692 B.n583 B.n318 10.6151
R1693 B.n584 B.n583 10.6151
R1694 B.n585 B.n584 10.6151
R1695 B.n585 B.n310 10.6151
R1696 B.n595 B.n310 10.6151
R1697 B.n596 B.n595 10.6151
R1698 B.n597 B.n596 10.6151
R1699 B.n597 B.n302 10.6151
R1700 B.n607 B.n302 10.6151
R1701 B.n608 B.n607 10.6151
R1702 B.n609 B.n608 10.6151
R1703 B.n609 B.n294 10.6151
R1704 B.n619 B.n294 10.6151
R1705 B.n620 B.n619 10.6151
R1706 B.n621 B.n620 10.6151
R1707 B.n621 B.n286 10.6151
R1708 B.n631 B.n286 10.6151
R1709 B.n632 B.n631 10.6151
R1710 B.n633 B.n632 10.6151
R1711 B.n633 B.n278 10.6151
R1712 B.n643 B.n278 10.6151
R1713 B.n644 B.n643 10.6151
R1714 B.n645 B.n644 10.6151
R1715 B.n645 B.n270 10.6151
R1716 B.n656 B.n270 10.6151
R1717 B.n657 B.n656 10.6151
R1718 B.n658 B.n657 10.6151
R1719 B.n658 B.n263 10.6151
R1720 B.n668 B.n263 10.6151
R1721 B.n669 B.n668 10.6151
R1722 B.n670 B.n669 10.6151
R1723 B.n670 B.n255 10.6151
R1724 B.n680 B.n255 10.6151
R1725 B.n681 B.n680 10.6151
R1726 B.n682 B.n681 10.6151
R1727 B.n682 B.n247 10.6151
R1728 B.n693 B.n247 10.6151
R1729 B.n694 B.n693 10.6151
R1730 B.n695 B.n694 10.6151
R1731 B.n695 B.n240 10.6151
R1732 B.n706 B.n240 10.6151
R1733 B.n707 B.n706 10.6151
R1734 B.n708 B.n707 10.6151
R1735 B.n708 B.n0 10.6151
R1736 B.n405 B.n381 10.6151
R1737 B.n405 B.n404 10.6151
R1738 B.n411 B.n404 10.6151
R1739 B.n412 B.n411 10.6151
R1740 B.n413 B.n412 10.6151
R1741 B.n413 B.n402 10.6151
R1742 B.n419 B.n402 10.6151
R1743 B.n420 B.n419 10.6151
R1744 B.n421 B.n420 10.6151
R1745 B.n421 B.n400 10.6151
R1746 B.n427 B.n400 10.6151
R1747 B.n428 B.n427 10.6151
R1748 B.n432 B.n428 10.6151
R1749 B.n438 B.n398 10.6151
R1750 B.n439 B.n438 10.6151
R1751 B.n440 B.n439 10.6151
R1752 B.n440 B.n396 10.6151
R1753 B.n446 B.n396 10.6151
R1754 B.n447 B.n446 10.6151
R1755 B.n448 B.n447 10.6151
R1756 B.n448 B.n394 10.6151
R1757 B.n454 B.n394 10.6151
R1758 B.n457 B.n456 10.6151
R1759 B.n457 B.n390 10.6151
R1760 B.n463 B.n390 10.6151
R1761 B.n464 B.n463 10.6151
R1762 B.n465 B.n464 10.6151
R1763 B.n465 B.n388 10.6151
R1764 B.n471 B.n388 10.6151
R1765 B.n472 B.n471 10.6151
R1766 B.n473 B.n472 10.6151
R1767 B.n473 B.n386 10.6151
R1768 B.n386 B.n385 10.6151
R1769 B.n480 B.n385 10.6151
R1770 B.n481 B.n480 10.6151
R1771 B.n482 B.n377 10.6151
R1772 B.n492 B.n377 10.6151
R1773 B.n493 B.n492 10.6151
R1774 B.n494 B.n493 10.6151
R1775 B.n494 B.n369 10.6151
R1776 B.n504 B.n369 10.6151
R1777 B.n505 B.n504 10.6151
R1778 B.n506 B.n505 10.6151
R1779 B.n506 B.n362 10.6151
R1780 B.n517 B.n362 10.6151
R1781 B.n518 B.n517 10.6151
R1782 B.n519 B.n518 10.6151
R1783 B.n519 B.n354 10.6151
R1784 B.n529 B.n354 10.6151
R1785 B.n530 B.n529 10.6151
R1786 B.n531 B.n530 10.6151
R1787 B.n531 B.n346 10.6151
R1788 B.n541 B.n346 10.6151
R1789 B.n542 B.n541 10.6151
R1790 B.n543 B.n542 10.6151
R1791 B.n543 B.n337 10.6151
R1792 B.n553 B.n337 10.6151
R1793 B.n554 B.n553 10.6151
R1794 B.n555 B.n554 10.6151
R1795 B.n555 B.n330 10.6151
R1796 B.n565 B.n330 10.6151
R1797 B.n566 B.n565 10.6151
R1798 B.n567 B.n566 10.6151
R1799 B.n567 B.n322 10.6151
R1800 B.n577 B.n322 10.6151
R1801 B.n578 B.n577 10.6151
R1802 B.n579 B.n578 10.6151
R1803 B.n579 B.n313 10.6151
R1804 B.n589 B.n313 10.6151
R1805 B.n590 B.n589 10.6151
R1806 B.n591 B.n590 10.6151
R1807 B.n591 B.n306 10.6151
R1808 B.n601 B.n306 10.6151
R1809 B.n602 B.n601 10.6151
R1810 B.n603 B.n602 10.6151
R1811 B.n603 B.n298 10.6151
R1812 B.n613 B.n298 10.6151
R1813 B.n614 B.n613 10.6151
R1814 B.n615 B.n614 10.6151
R1815 B.n615 B.n290 10.6151
R1816 B.n625 B.n290 10.6151
R1817 B.n626 B.n625 10.6151
R1818 B.n627 B.n626 10.6151
R1819 B.n627 B.n282 10.6151
R1820 B.n637 B.n282 10.6151
R1821 B.n638 B.n637 10.6151
R1822 B.n639 B.n638 10.6151
R1823 B.n639 B.n274 10.6151
R1824 B.n649 B.n274 10.6151
R1825 B.n650 B.n649 10.6151
R1826 B.n651 B.n650 10.6151
R1827 B.n651 B.n267 10.6151
R1828 B.n662 B.n267 10.6151
R1829 B.n663 B.n662 10.6151
R1830 B.n664 B.n663 10.6151
R1831 B.n664 B.n259 10.6151
R1832 B.n674 B.n259 10.6151
R1833 B.n675 B.n674 10.6151
R1834 B.n676 B.n675 10.6151
R1835 B.n676 B.n251 10.6151
R1836 B.n686 B.n251 10.6151
R1837 B.n687 B.n686 10.6151
R1838 B.n688 B.n687 10.6151
R1839 B.n688 B.n244 10.6151
R1840 B.n699 B.n244 10.6151
R1841 B.n700 B.n699 10.6151
R1842 B.n702 B.n700 10.6151
R1843 B.n702 B.n701 10.6151
R1844 B.n701 B.n236 10.6151
R1845 B.n713 B.n236 10.6151
R1846 B.n714 B.n713 10.6151
R1847 B.n715 B.n714 10.6151
R1848 B.n716 B.n715 10.6151
R1849 B.n717 B.n716 10.6151
R1850 B.n720 B.n717 10.6151
R1851 B.n721 B.n720 10.6151
R1852 B.n722 B.n721 10.6151
R1853 B.n723 B.n722 10.6151
R1854 B.n725 B.n723 10.6151
R1855 B.n726 B.n725 10.6151
R1856 B.n727 B.n726 10.6151
R1857 B.n728 B.n727 10.6151
R1858 B.n730 B.n728 10.6151
R1859 B.n731 B.n730 10.6151
R1860 B.n732 B.n731 10.6151
R1861 B.n733 B.n732 10.6151
R1862 B.n735 B.n733 10.6151
R1863 B.n736 B.n735 10.6151
R1864 B.n737 B.n736 10.6151
R1865 B.n738 B.n737 10.6151
R1866 B.n740 B.n738 10.6151
R1867 B.n741 B.n740 10.6151
R1868 B.n742 B.n741 10.6151
R1869 B.n743 B.n742 10.6151
R1870 B.n745 B.n743 10.6151
R1871 B.n746 B.n745 10.6151
R1872 B.n747 B.n746 10.6151
R1873 B.n748 B.n747 10.6151
R1874 B.n750 B.n748 10.6151
R1875 B.n751 B.n750 10.6151
R1876 B.n752 B.n751 10.6151
R1877 B.n753 B.n752 10.6151
R1878 B.n755 B.n753 10.6151
R1879 B.n756 B.n755 10.6151
R1880 B.n757 B.n756 10.6151
R1881 B.n758 B.n757 10.6151
R1882 B.n760 B.n758 10.6151
R1883 B.n761 B.n760 10.6151
R1884 B.n762 B.n761 10.6151
R1885 B.n763 B.n762 10.6151
R1886 B.n765 B.n763 10.6151
R1887 B.n766 B.n765 10.6151
R1888 B.n767 B.n766 10.6151
R1889 B.n768 B.n767 10.6151
R1890 B.n770 B.n768 10.6151
R1891 B.n771 B.n770 10.6151
R1892 B.n772 B.n771 10.6151
R1893 B.n773 B.n772 10.6151
R1894 B.n775 B.n773 10.6151
R1895 B.n776 B.n775 10.6151
R1896 B.n777 B.n776 10.6151
R1897 B.n778 B.n777 10.6151
R1898 B.n780 B.n778 10.6151
R1899 B.n781 B.n780 10.6151
R1900 B.n782 B.n781 10.6151
R1901 B.n783 B.n782 10.6151
R1902 B.n785 B.n783 10.6151
R1903 B.n786 B.n785 10.6151
R1904 B.n787 B.n786 10.6151
R1905 B.n788 B.n787 10.6151
R1906 B.n790 B.n788 10.6151
R1907 B.n791 B.n790 10.6151
R1908 B.n792 B.n791 10.6151
R1909 B.n793 B.n792 10.6151
R1910 B.n795 B.n793 10.6151
R1911 B.n796 B.n795 10.6151
R1912 B.n797 B.n796 10.6151
R1913 B.n798 B.n797 10.6151
R1914 B.n800 B.n798 10.6151
R1915 B.n801 B.n800 10.6151
R1916 B.n802 B.n801 10.6151
R1917 B.n803 B.n802 10.6151
R1918 B.n805 B.n803 10.6151
R1919 B.n806 B.n805 10.6151
R1920 B.n807 B.n806 10.6151
R1921 B.n808 B.n807 10.6151
R1922 B.n810 B.n808 10.6151
R1923 B.n811 B.n810 10.6151
R1924 B.n964 B.n1 10.6151
R1925 B.n964 B.n963 10.6151
R1926 B.n963 B.n962 10.6151
R1927 B.n962 B.n10 10.6151
R1928 B.n956 B.n10 10.6151
R1929 B.n956 B.n955 10.6151
R1930 B.n955 B.n954 10.6151
R1931 B.n954 B.n17 10.6151
R1932 B.n948 B.n17 10.6151
R1933 B.n948 B.n947 10.6151
R1934 B.n947 B.n946 10.6151
R1935 B.n946 B.n25 10.6151
R1936 B.n940 B.n25 10.6151
R1937 B.n940 B.n939 10.6151
R1938 B.n939 B.n938 10.6151
R1939 B.n938 B.n32 10.6151
R1940 B.n932 B.n32 10.6151
R1941 B.n932 B.n931 10.6151
R1942 B.n931 B.n930 10.6151
R1943 B.n930 B.n38 10.6151
R1944 B.n924 B.n38 10.6151
R1945 B.n924 B.n923 10.6151
R1946 B.n923 B.n922 10.6151
R1947 B.n922 B.n46 10.6151
R1948 B.n916 B.n46 10.6151
R1949 B.n916 B.n915 10.6151
R1950 B.n915 B.n914 10.6151
R1951 B.n914 B.n53 10.6151
R1952 B.n908 B.n53 10.6151
R1953 B.n908 B.n907 10.6151
R1954 B.n907 B.n906 10.6151
R1955 B.n906 B.n60 10.6151
R1956 B.n900 B.n60 10.6151
R1957 B.n900 B.n899 10.6151
R1958 B.n899 B.n898 10.6151
R1959 B.n898 B.n67 10.6151
R1960 B.n892 B.n67 10.6151
R1961 B.n892 B.n891 10.6151
R1962 B.n891 B.n890 10.6151
R1963 B.n890 B.n74 10.6151
R1964 B.n884 B.n74 10.6151
R1965 B.n884 B.n883 10.6151
R1966 B.n883 B.n882 10.6151
R1967 B.n882 B.n81 10.6151
R1968 B.n876 B.n81 10.6151
R1969 B.n876 B.n875 10.6151
R1970 B.n875 B.n874 10.6151
R1971 B.n874 B.n88 10.6151
R1972 B.n868 B.n88 10.6151
R1973 B.n868 B.n867 10.6151
R1974 B.n867 B.n866 10.6151
R1975 B.n866 B.n95 10.6151
R1976 B.n860 B.n95 10.6151
R1977 B.n860 B.n859 10.6151
R1978 B.n859 B.n858 10.6151
R1979 B.n858 B.n102 10.6151
R1980 B.n852 B.n102 10.6151
R1981 B.n852 B.n851 10.6151
R1982 B.n851 B.n850 10.6151
R1983 B.n850 B.n109 10.6151
R1984 B.n844 B.n109 10.6151
R1985 B.n844 B.n843 10.6151
R1986 B.n843 B.n842 10.6151
R1987 B.n842 B.n116 10.6151
R1988 B.n836 B.n116 10.6151
R1989 B.n836 B.n835 10.6151
R1990 B.n835 B.n834 10.6151
R1991 B.n834 B.n122 10.6151
R1992 B.n828 B.n122 10.6151
R1993 B.n828 B.n827 10.6151
R1994 B.n827 B.n826 10.6151
R1995 B.n826 B.n130 10.6151
R1996 B.n820 B.n130 10.6151
R1997 B.n820 B.n819 10.6151
R1998 B.n819 B.n818 10.6151
R1999 B.n165 B.n137 10.6151
R2000 B.n168 B.n165 10.6151
R2001 B.n169 B.n168 10.6151
R2002 B.n172 B.n169 10.6151
R2003 B.n173 B.n172 10.6151
R2004 B.n176 B.n173 10.6151
R2005 B.n177 B.n176 10.6151
R2006 B.n180 B.n177 10.6151
R2007 B.n181 B.n180 10.6151
R2008 B.n184 B.n181 10.6151
R2009 B.n185 B.n184 10.6151
R2010 B.n188 B.n185 10.6151
R2011 B.n189 B.n188 10.6151
R2012 B.n193 B.n192 10.6151
R2013 B.n196 B.n193 10.6151
R2014 B.n197 B.n196 10.6151
R2015 B.n200 B.n197 10.6151
R2016 B.n201 B.n200 10.6151
R2017 B.n204 B.n201 10.6151
R2018 B.n205 B.n204 10.6151
R2019 B.n208 B.n205 10.6151
R2020 B.n209 B.n208 10.6151
R2021 B.n213 B.n212 10.6151
R2022 B.n216 B.n213 10.6151
R2023 B.n217 B.n216 10.6151
R2024 B.n220 B.n217 10.6151
R2025 B.n221 B.n220 10.6151
R2026 B.n224 B.n221 10.6151
R2027 B.n225 B.n224 10.6151
R2028 B.n228 B.n225 10.6151
R2029 B.n229 B.n228 10.6151
R2030 B.n232 B.n229 10.6151
R2031 B.n234 B.n232 10.6151
R2032 B.n235 B.n234 10.6151
R2033 B.n812 B.n235 10.6151
R2034 B.n432 B.n431 9.36635
R2035 B.n456 B.n455 9.36635
R2036 B.n189 B.n164 9.36635
R2037 B.n212 B.n161 9.36635
R2038 B.n508 B.t11 8.266
R2039 B.n124 B.t15 8.266
R2040 B.n972 B.n0 8.11757
R2041 B.n972 B.n1 8.11757
R2042 B.n316 B.t1 5.51083
R2043 B.t3 B.n887 5.51083
R2044 B.n431 B.n398 1.24928
R2045 B.n455 B.n454 1.24928
R2046 B.n192 B.n164 1.24928
R2047 B.n209 B.n161 1.24928
R2048 VP.n32 VP.n31 161.3
R2049 VP.n33 VP.n28 161.3
R2050 VP.n35 VP.n34 161.3
R2051 VP.n36 VP.n27 161.3
R2052 VP.n38 VP.n37 161.3
R2053 VP.n39 VP.n26 161.3
R2054 VP.n41 VP.n40 161.3
R2055 VP.n42 VP.n25 161.3
R2056 VP.n44 VP.n43 161.3
R2057 VP.n45 VP.n24 161.3
R2058 VP.n47 VP.n46 161.3
R2059 VP.n48 VP.n23 161.3
R2060 VP.n50 VP.n49 161.3
R2061 VP.n51 VP.n22 161.3
R2062 VP.n54 VP.n53 161.3
R2063 VP.n55 VP.n21 161.3
R2064 VP.n57 VP.n56 161.3
R2065 VP.n58 VP.n20 161.3
R2066 VP.n60 VP.n59 161.3
R2067 VP.n61 VP.n19 161.3
R2068 VP.n63 VP.n62 161.3
R2069 VP.n64 VP.n18 161.3
R2070 VP.n66 VP.n65 161.3
R2071 VP.n117 VP.n116 161.3
R2072 VP.n115 VP.n1 161.3
R2073 VP.n114 VP.n113 161.3
R2074 VP.n112 VP.n2 161.3
R2075 VP.n111 VP.n110 161.3
R2076 VP.n109 VP.n3 161.3
R2077 VP.n108 VP.n107 161.3
R2078 VP.n106 VP.n4 161.3
R2079 VP.n105 VP.n104 161.3
R2080 VP.n102 VP.n5 161.3
R2081 VP.n101 VP.n100 161.3
R2082 VP.n99 VP.n6 161.3
R2083 VP.n98 VP.n97 161.3
R2084 VP.n96 VP.n7 161.3
R2085 VP.n95 VP.n94 161.3
R2086 VP.n93 VP.n8 161.3
R2087 VP.n92 VP.n91 161.3
R2088 VP.n90 VP.n9 161.3
R2089 VP.n89 VP.n88 161.3
R2090 VP.n87 VP.n10 161.3
R2091 VP.n86 VP.n85 161.3
R2092 VP.n84 VP.n11 161.3
R2093 VP.n83 VP.n82 161.3
R2094 VP.n81 VP.n80 161.3
R2095 VP.n79 VP.n13 161.3
R2096 VP.n78 VP.n77 161.3
R2097 VP.n76 VP.n14 161.3
R2098 VP.n75 VP.n74 161.3
R2099 VP.n73 VP.n15 161.3
R2100 VP.n72 VP.n71 161.3
R2101 VP.n70 VP.n16 161.3
R2102 VP.n69 VP.n68 78.3232
R2103 VP.n118 VP.n0 78.3232
R2104 VP.n67 VP.n17 78.3232
R2105 VP.n30 VP.n29 56.5559
R2106 VP.n74 VP.n14 56.5193
R2107 VP.n110 VP.n2 56.5193
R2108 VP.n59 VP.n19 56.5193
R2109 VP.n30 VP.t9 52.097
R2110 VP.n69 VP.n67 51.3137
R2111 VP.n89 VP.n10 46.8066
R2112 VP.n97 VP.n6 46.8066
R2113 VP.n46 VP.n23 46.8066
R2114 VP.n38 VP.n27 46.8066
R2115 VP.n85 VP.n10 34.1802
R2116 VP.n101 VP.n6 34.1802
R2117 VP.n50 VP.n23 34.1802
R2118 VP.n34 VP.n27 34.1802
R2119 VP.n72 VP.n16 24.4675
R2120 VP.n73 VP.n72 24.4675
R2121 VP.n74 VP.n73 24.4675
R2122 VP.n78 VP.n14 24.4675
R2123 VP.n79 VP.n78 24.4675
R2124 VP.n80 VP.n79 24.4675
R2125 VP.n84 VP.n83 24.4675
R2126 VP.n85 VP.n84 24.4675
R2127 VP.n90 VP.n89 24.4675
R2128 VP.n91 VP.n90 24.4675
R2129 VP.n91 VP.n8 24.4675
R2130 VP.n95 VP.n8 24.4675
R2131 VP.n96 VP.n95 24.4675
R2132 VP.n97 VP.n96 24.4675
R2133 VP.n102 VP.n101 24.4675
R2134 VP.n104 VP.n102 24.4675
R2135 VP.n108 VP.n4 24.4675
R2136 VP.n109 VP.n108 24.4675
R2137 VP.n110 VP.n109 24.4675
R2138 VP.n114 VP.n2 24.4675
R2139 VP.n115 VP.n114 24.4675
R2140 VP.n116 VP.n115 24.4675
R2141 VP.n63 VP.n19 24.4675
R2142 VP.n64 VP.n63 24.4675
R2143 VP.n65 VP.n64 24.4675
R2144 VP.n51 VP.n50 24.4675
R2145 VP.n53 VP.n51 24.4675
R2146 VP.n57 VP.n21 24.4675
R2147 VP.n58 VP.n57 24.4675
R2148 VP.n59 VP.n58 24.4675
R2149 VP.n39 VP.n38 24.4675
R2150 VP.n40 VP.n39 24.4675
R2151 VP.n40 VP.n25 24.4675
R2152 VP.n44 VP.n25 24.4675
R2153 VP.n45 VP.n44 24.4675
R2154 VP.n46 VP.n45 24.4675
R2155 VP.n33 VP.n32 24.4675
R2156 VP.n34 VP.n33 24.4675
R2157 VP.n8 VP.t0 18.4499
R2158 VP.n68 VP.t5 18.4499
R2159 VP.n12 VP.t4 18.4499
R2160 VP.n103 VP.t6 18.4499
R2161 VP.n0 VP.t8 18.4499
R2162 VP.n25 VP.t3 18.4499
R2163 VP.n17 VP.t2 18.4499
R2164 VP.n52 VP.t1 18.4499
R2165 VP.n29 VP.t7 18.4499
R2166 VP.n83 VP.n12 18.1061
R2167 VP.n104 VP.n103 18.1061
R2168 VP.n53 VP.n52 18.1061
R2169 VP.n32 VP.n29 18.1061
R2170 VP.n68 VP.n16 11.7447
R2171 VP.n116 VP.n0 11.7447
R2172 VP.n65 VP.n17 11.7447
R2173 VP.n80 VP.n12 6.36192
R2174 VP.n103 VP.n4 6.36192
R2175 VP.n52 VP.n21 6.36192
R2176 VP.n31 VP.n30 3.10013
R2177 VP.n67 VP.n66 0.354971
R2178 VP.n70 VP.n69 0.354971
R2179 VP.n118 VP.n117 0.354971
R2180 VP VP.n118 0.26696
R2181 VP.n31 VP.n28 0.189894
R2182 VP.n35 VP.n28 0.189894
R2183 VP.n36 VP.n35 0.189894
R2184 VP.n37 VP.n36 0.189894
R2185 VP.n37 VP.n26 0.189894
R2186 VP.n41 VP.n26 0.189894
R2187 VP.n42 VP.n41 0.189894
R2188 VP.n43 VP.n42 0.189894
R2189 VP.n43 VP.n24 0.189894
R2190 VP.n47 VP.n24 0.189894
R2191 VP.n48 VP.n47 0.189894
R2192 VP.n49 VP.n48 0.189894
R2193 VP.n49 VP.n22 0.189894
R2194 VP.n54 VP.n22 0.189894
R2195 VP.n55 VP.n54 0.189894
R2196 VP.n56 VP.n55 0.189894
R2197 VP.n56 VP.n20 0.189894
R2198 VP.n60 VP.n20 0.189894
R2199 VP.n61 VP.n60 0.189894
R2200 VP.n62 VP.n61 0.189894
R2201 VP.n62 VP.n18 0.189894
R2202 VP.n66 VP.n18 0.189894
R2203 VP.n71 VP.n70 0.189894
R2204 VP.n71 VP.n15 0.189894
R2205 VP.n75 VP.n15 0.189894
R2206 VP.n76 VP.n75 0.189894
R2207 VP.n77 VP.n76 0.189894
R2208 VP.n77 VP.n13 0.189894
R2209 VP.n81 VP.n13 0.189894
R2210 VP.n82 VP.n81 0.189894
R2211 VP.n82 VP.n11 0.189894
R2212 VP.n86 VP.n11 0.189894
R2213 VP.n87 VP.n86 0.189894
R2214 VP.n88 VP.n87 0.189894
R2215 VP.n88 VP.n9 0.189894
R2216 VP.n92 VP.n9 0.189894
R2217 VP.n93 VP.n92 0.189894
R2218 VP.n94 VP.n93 0.189894
R2219 VP.n94 VP.n7 0.189894
R2220 VP.n98 VP.n7 0.189894
R2221 VP.n99 VP.n98 0.189894
R2222 VP.n100 VP.n99 0.189894
R2223 VP.n100 VP.n5 0.189894
R2224 VP.n105 VP.n5 0.189894
R2225 VP.n106 VP.n105 0.189894
R2226 VP.n107 VP.n106 0.189894
R2227 VP.n107 VP.n3 0.189894
R2228 VP.n111 VP.n3 0.189894
R2229 VP.n112 VP.n111 0.189894
R2230 VP.n113 VP.n112 0.189894
R2231 VP.n113 VP.n1 0.189894
R2232 VP.n117 VP.n1 0.189894
R2233 VDD1.n6 VDD1.n0 289.615
R2234 VDD1.n19 VDD1.n13 289.615
R2235 VDD1.n7 VDD1.n6 185
R2236 VDD1.n5 VDD1.n4 185
R2237 VDD1.n18 VDD1.n17 185
R2238 VDD1.n20 VDD1.n19 185
R2239 VDD1.n16 VDD1.t4 153.582
R2240 VDD1.n3 VDD1.t0 153.582
R2241 VDD1.n6 VDD1.n5 104.615
R2242 VDD1.n19 VDD1.n18 104.615
R2243 VDD1.n27 VDD1.n26 87.8952
R2244 VDD1.n29 VDD1.n28 85.4484
R2245 VDD1.n12 VDD1.n11 85.4484
R2246 VDD1.n25 VDD1.n24 85.4484
R2247 VDD1.n5 VDD1.t0 52.3082
R2248 VDD1.n18 VDD1.t4 52.3082
R2249 VDD1.n12 VDD1.n10 51.2306
R2250 VDD1.n25 VDD1.n23 51.2306
R2251 VDD1.n29 VDD1.n27 44.1496
R2252 VDD1.n4 VDD1.n3 10.1164
R2253 VDD1.n17 VDD1.n16 10.1164
R2254 VDD1.n10 VDD1.n9 9.45567
R2255 VDD1.n23 VDD1.n22 9.45567
R2256 VDD1.n9 VDD1.n8 9.3005
R2257 VDD1.n2 VDD1.n1 9.3005
R2258 VDD1.n15 VDD1.n14 9.3005
R2259 VDD1.n22 VDD1.n21 9.3005
R2260 VDD1.n10 VDD1.n0 8.92171
R2261 VDD1.n23 VDD1.n13 8.92171
R2262 VDD1.n8 VDD1.n7 8.14595
R2263 VDD1.n21 VDD1.n20 8.14595
R2264 VDD1.n4 VDD1.n2 7.3702
R2265 VDD1.n17 VDD1.n15 7.3702
R2266 VDD1.n28 VDD1.t8 7.30677
R2267 VDD1.n28 VDD1.t7 7.30677
R2268 VDD1.n11 VDD1.t2 7.30677
R2269 VDD1.n11 VDD1.t6 7.30677
R2270 VDD1.n26 VDD1.t3 7.30677
R2271 VDD1.n26 VDD1.t1 7.30677
R2272 VDD1.n24 VDD1.t5 7.30677
R2273 VDD1.n24 VDD1.t9 7.30677
R2274 VDD1.n7 VDD1.n2 5.81868
R2275 VDD1.n20 VDD1.n15 5.81868
R2276 VDD1.n8 VDD1.n0 5.04292
R2277 VDD1.n21 VDD1.n13 5.04292
R2278 VDD1.n3 VDD1.n1 3.00987
R2279 VDD1.n16 VDD1.n14 3.00987
R2280 VDD1 VDD1.n29 2.44447
R2281 VDD1 VDD1.n12 0.892741
R2282 VDD1.n27 VDD1.n25 0.779206
R2283 VDD1.n9 VDD1.n1 0.155672
R2284 VDD1.n22 VDD1.n14 0.155672
C0 VN VDD1 0.161014f
C1 VN VDD2 2.9679f
C2 VDD1 VTAIL 7.11812f
C3 VDD2 VTAIL 7.17773f
C4 VDD1 VDD2 2.78591f
C5 VP VN 8.06994f
C6 VP VTAIL 4.83532f
C7 VP VDD1 3.51227f
C8 VP VDD2 0.709656f
C9 VN VTAIL 4.82118f
C10 VDD2 B 6.825221f
C11 VDD1 B 6.670863f
C12 VTAIL B 4.535096f
C13 VN B 21.872019f
C14 VP B 20.246176f
C15 VDD1.n0 B 0.044701f
C16 VDD1.n1 B 0.265422f
C17 VDD1.n2 B 0.016232f
C18 VDD1.t0 B 0.070255f
C19 VDD1.n3 B 0.114244f
C20 VDD1.n4 B 0.02627f
C21 VDD1.n5 B 0.028776f
C22 VDD1.n6 B 0.087023f
C23 VDD1.n7 B 0.017187f
C24 VDD1.n8 B 0.016232f
C25 VDD1.n9 B 0.06776f
C26 VDD1.n10 B 0.094769f
C27 VDD1.t2 B 0.064691f
C28 VDD1.t6 B 0.064691f
C29 VDD1.n11 B 0.452006f
C30 VDD1.n12 B 1.00884f
C31 VDD1.n13 B 0.044701f
C32 VDD1.n14 B 0.265422f
C33 VDD1.n15 B 0.016232f
C34 VDD1.t4 B 0.070255f
C35 VDD1.n16 B 0.114244f
C36 VDD1.n17 B 0.02627f
C37 VDD1.n18 B 0.028776f
C38 VDD1.n19 B 0.087023f
C39 VDD1.n20 B 0.017187f
C40 VDD1.n21 B 0.016232f
C41 VDD1.n22 B 0.06776f
C42 VDD1.n23 B 0.094769f
C43 VDD1.t5 B 0.064691f
C44 VDD1.t9 B 0.064691f
C45 VDD1.n24 B 0.452005f
C46 VDD1.n25 B 0.99869f
C47 VDD1.t3 B 0.064691f
C48 VDD1.t1 B 0.064691f
C49 VDD1.n26 B 0.474713f
C50 VDD1.n27 B 3.58882f
C51 VDD1.t8 B 0.064691f
C52 VDD1.t7 B 0.064691f
C53 VDD1.n28 B 0.452006f
C54 VDD1.n29 B 3.43292f
C55 VP.t8 B 0.598904f
C56 VP.n0 B 0.352747f
C57 VP.n1 B 0.025401f
C58 VP.n2 B 0.03319f
C59 VP.n3 B 0.025401f
C60 VP.n4 B 0.030045f
C61 VP.n5 B 0.025401f
C62 VP.n6 B 0.021948f
C63 VP.n7 B 0.025401f
C64 VP.t0 B 0.598904f
C65 VP.n8 B 0.274975f
C66 VP.n9 B 0.025401f
C67 VP.n10 B 0.021948f
C68 VP.n11 B 0.025401f
C69 VP.t4 B 0.598904f
C70 VP.n12 B 0.251006f
C71 VP.n13 B 0.025401f
C72 VP.n14 B 0.040976f
C73 VP.n15 B 0.025401f
C74 VP.n16 B 0.035187f
C75 VP.t2 B 0.598904f
C76 VP.n17 B 0.352747f
C77 VP.n18 B 0.025401f
C78 VP.n19 B 0.03319f
C79 VP.n20 B 0.025401f
C80 VP.n21 B 0.030045f
C81 VP.n22 B 0.025401f
C82 VP.n23 B 0.021948f
C83 VP.n24 B 0.025401f
C84 VP.t3 B 0.598904f
C85 VP.n25 B 0.274975f
C86 VP.n26 B 0.025401f
C87 VP.n27 B 0.021948f
C88 VP.n28 B 0.025401f
C89 VP.t7 B 0.598904f
C90 VP.n29 B 0.344925f
C91 VP.t9 B 0.885577f
C92 VP.n30 B 0.35301f
C93 VP.n31 B 0.314226f
C94 VP.n32 B 0.041264f
C95 VP.n33 B 0.047341f
C96 VP.n34 B 0.051325f
C97 VP.n35 B 0.025401f
C98 VP.n36 B 0.025401f
C99 VP.n37 B 0.025401f
C100 VP.n38 B 0.048233f
C101 VP.n39 B 0.047341f
C102 VP.n40 B 0.047341f
C103 VP.n41 B 0.025401f
C104 VP.n42 B 0.025401f
C105 VP.n43 B 0.025401f
C106 VP.n44 B 0.047341f
C107 VP.n45 B 0.047341f
C108 VP.n46 B 0.048233f
C109 VP.n47 B 0.025401f
C110 VP.n48 B 0.025401f
C111 VP.n49 B 0.025401f
C112 VP.n50 B 0.051325f
C113 VP.n51 B 0.047341f
C114 VP.t1 B 0.598904f
C115 VP.n52 B 0.251006f
C116 VP.n53 B 0.041264f
C117 VP.n54 B 0.025401f
C118 VP.n55 B 0.025401f
C119 VP.n56 B 0.025401f
C120 VP.n57 B 0.047341f
C121 VP.n58 B 0.047341f
C122 VP.n59 B 0.040976f
C123 VP.n60 B 0.025401f
C124 VP.n61 B 0.025401f
C125 VP.n62 B 0.025401f
C126 VP.n63 B 0.047341f
C127 VP.n64 B 0.047341f
C128 VP.n65 B 0.035187f
C129 VP.n66 B 0.040996f
C130 VP.n67 B 1.50627f
C131 VP.t5 B 0.598904f
C132 VP.n68 B 0.352747f
C133 VP.n69 B 1.52407f
C134 VP.n70 B 0.040996f
C135 VP.n71 B 0.025401f
C136 VP.n72 B 0.047341f
C137 VP.n73 B 0.047341f
C138 VP.n74 B 0.03319f
C139 VP.n75 B 0.025401f
C140 VP.n76 B 0.025401f
C141 VP.n77 B 0.025401f
C142 VP.n78 B 0.047341f
C143 VP.n79 B 0.047341f
C144 VP.n80 B 0.030045f
C145 VP.n81 B 0.025401f
C146 VP.n82 B 0.025401f
C147 VP.n83 B 0.041264f
C148 VP.n84 B 0.047341f
C149 VP.n85 B 0.051325f
C150 VP.n86 B 0.025401f
C151 VP.n87 B 0.025401f
C152 VP.n88 B 0.025401f
C153 VP.n89 B 0.048233f
C154 VP.n90 B 0.047341f
C155 VP.n91 B 0.047341f
C156 VP.n92 B 0.025401f
C157 VP.n93 B 0.025401f
C158 VP.n94 B 0.025401f
C159 VP.n95 B 0.047341f
C160 VP.n96 B 0.047341f
C161 VP.n97 B 0.048233f
C162 VP.n98 B 0.025401f
C163 VP.n99 B 0.025401f
C164 VP.n100 B 0.025401f
C165 VP.n101 B 0.051325f
C166 VP.n102 B 0.047341f
C167 VP.t6 B 0.598904f
C168 VP.n103 B 0.251006f
C169 VP.n104 B 0.041264f
C170 VP.n105 B 0.025401f
C171 VP.n106 B 0.025401f
C172 VP.n107 B 0.025401f
C173 VP.n108 B 0.047341f
C174 VP.n109 B 0.047341f
C175 VP.n110 B 0.040976f
C176 VP.n111 B 0.025401f
C177 VP.n112 B 0.025401f
C178 VP.n113 B 0.025401f
C179 VP.n114 B 0.047341f
C180 VP.n115 B 0.047341f
C181 VP.n116 B 0.035187f
C182 VP.n117 B 0.040996f
C183 VP.n118 B 0.067044f
C184 VDD2.n0 B 0.043731f
C185 VDD2.n1 B 0.259661f
C186 VDD2.n2 B 0.01588f
C187 VDD2.t8 B 0.06873f
C188 VDD2.n3 B 0.111764f
C189 VDD2.n4 B 0.0257f
C190 VDD2.n5 B 0.028151f
C191 VDD2.n6 B 0.085134f
C192 VDD2.n7 B 0.016814f
C193 VDD2.n8 B 0.01588f
C194 VDD2.n9 B 0.06629f
C195 VDD2.n10 B 0.092712f
C196 VDD2.t4 B 0.063286f
C197 VDD2.t9 B 0.063286f
C198 VDD2.n11 B 0.442194f
C199 VDD2.n12 B 0.977013f
C200 VDD2.t3 B 0.063286f
C201 VDD2.t5 B 0.063286f
C202 VDD2.n13 B 0.46441f
C203 VDD2.n14 B 3.34352f
C204 VDD2.n15 B 0.043731f
C205 VDD2.n16 B 0.259661f
C206 VDD2.n17 B 0.01588f
C207 VDD2.t7 B 0.06873f
C208 VDD2.n18 B 0.111764f
C209 VDD2.n19 B 0.0257f
C210 VDD2.n20 B 0.028151f
C211 VDD2.n21 B 0.085134f
C212 VDD2.n22 B 0.016814f
C213 VDD2.n23 B 0.01588f
C214 VDD2.n24 B 0.06629f
C215 VDD2.n25 B 0.068393f
C216 VDD2.n26 B 2.9926f
C217 VDD2.t6 B 0.063286f
C218 VDD2.t2 B 0.063286f
C219 VDD2.n27 B 0.442195f
C220 VDD2.n28 B 0.637827f
C221 VDD2.t0 B 0.063286f
C222 VDD2.t1 B 0.063286f
C223 VDD2.n29 B 0.464371f
C224 VTAIL.t19 B 0.07698f
C225 VTAIL.t13 B 0.07698f
C226 VTAIL.n0 B 0.470155f
C227 VTAIL.n1 B 0.849126f
C228 VTAIL.n2 B 0.053194f
C229 VTAIL.n3 B 0.315847f
C230 VTAIL.n4 B 0.019316f
C231 VTAIL.t5 B 0.083602f
C232 VTAIL.n5 B 0.135948f
C233 VTAIL.n6 B 0.031261f
C234 VTAIL.n7 B 0.034242f
C235 VTAIL.n8 B 0.103556f
C236 VTAIL.n9 B 0.020452f
C237 VTAIL.n10 B 0.019316f
C238 VTAIL.n11 B 0.080633f
C239 VTAIL.n12 B 0.058352f
C240 VTAIL.n13 B 0.663374f
C241 VTAIL.t7 B 0.07698f
C242 VTAIL.t2 B 0.07698f
C243 VTAIL.n14 B 0.470155f
C244 VTAIL.n15 B 1.07779f
C245 VTAIL.t8 B 0.07698f
C246 VTAIL.t1 B 0.07698f
C247 VTAIL.n16 B 0.470155f
C248 VTAIL.n17 B 2.2231f
C249 VTAIL.t15 B 0.07698f
C250 VTAIL.t14 B 0.07698f
C251 VTAIL.n18 B 0.470157f
C252 VTAIL.n19 B 2.2231f
C253 VTAIL.t11 B 0.07698f
C254 VTAIL.t10 B 0.07698f
C255 VTAIL.n20 B 0.470157f
C256 VTAIL.n21 B 1.07778f
C257 VTAIL.n22 B 0.053194f
C258 VTAIL.n23 B 0.315847f
C259 VTAIL.n24 B 0.019316f
C260 VTAIL.t18 B 0.083602f
C261 VTAIL.n25 B 0.135948f
C262 VTAIL.n26 B 0.031261f
C263 VTAIL.n27 B 0.034242f
C264 VTAIL.n28 B 0.103556f
C265 VTAIL.n29 B 0.020452f
C266 VTAIL.n30 B 0.019316f
C267 VTAIL.n31 B 0.080633f
C268 VTAIL.n32 B 0.058352f
C269 VTAIL.n33 B 0.663374f
C270 VTAIL.t0 B 0.07698f
C271 VTAIL.t4 B 0.07698f
C272 VTAIL.n34 B 0.470157f
C273 VTAIL.n35 B 0.93899f
C274 VTAIL.t9 B 0.07698f
C275 VTAIL.t3 B 0.07698f
C276 VTAIL.n36 B 0.470157f
C277 VTAIL.n37 B 1.07778f
C278 VTAIL.n38 B 0.053194f
C279 VTAIL.n39 B 0.315847f
C280 VTAIL.n40 B 0.019316f
C281 VTAIL.t6 B 0.083602f
C282 VTAIL.n41 B 0.135948f
C283 VTAIL.n42 B 0.031261f
C284 VTAIL.n43 B 0.034242f
C285 VTAIL.n44 B 0.103556f
C286 VTAIL.n45 B 0.020452f
C287 VTAIL.n46 B 0.019316f
C288 VTAIL.n47 B 0.080633f
C289 VTAIL.n48 B 0.058352f
C290 VTAIL.n49 B 1.56106f
C291 VTAIL.n50 B 0.053194f
C292 VTAIL.n51 B 0.315847f
C293 VTAIL.n52 B 0.019316f
C294 VTAIL.t17 B 0.083602f
C295 VTAIL.n53 B 0.135948f
C296 VTAIL.n54 B 0.031261f
C297 VTAIL.n55 B 0.034242f
C298 VTAIL.n56 B 0.103556f
C299 VTAIL.n57 B 0.020452f
C300 VTAIL.n58 B 0.019316f
C301 VTAIL.n59 B 0.080633f
C302 VTAIL.n60 B 0.058352f
C303 VTAIL.n61 B 1.56106f
C304 VTAIL.t16 B 0.07698f
C305 VTAIL.t12 B 0.07698f
C306 VTAIL.n62 B 0.470155f
C307 VTAIL.n63 B 0.781227f
C308 VN.t4 B 0.579384f
C309 VN.n0 B 0.341249f
C310 VN.n1 B 0.024573f
C311 VN.n2 B 0.032108f
C312 VN.n3 B 0.024573f
C313 VN.n4 B 0.029066f
C314 VN.n5 B 0.024573f
C315 VN.n6 B 0.021232f
C316 VN.n7 B 0.024573f
C317 VN.t0 B 0.579384f
C318 VN.n8 B 0.266012f
C319 VN.n9 B 0.024573f
C320 VN.n10 B 0.021232f
C321 VN.n11 B 0.024573f
C322 VN.t5 B 0.579384f
C323 VN.n12 B 0.333683f
C324 VN.t1 B 0.856714f
C325 VN.n13 B 0.341503f
C326 VN.n14 B 0.303984f
C327 VN.n15 B 0.039919f
C328 VN.n16 B 0.045798f
C329 VN.n17 B 0.049652f
C330 VN.n18 B 0.024573f
C331 VN.n19 B 0.024573f
C332 VN.n20 B 0.024573f
C333 VN.n21 B 0.046661f
C334 VN.n22 B 0.045798f
C335 VN.n23 B 0.045798f
C336 VN.n24 B 0.024573f
C337 VN.n25 B 0.024573f
C338 VN.n26 B 0.024573f
C339 VN.n27 B 0.045798f
C340 VN.n28 B 0.045798f
C341 VN.n29 B 0.046661f
C342 VN.n30 B 0.024573f
C343 VN.n31 B 0.024573f
C344 VN.n32 B 0.024573f
C345 VN.n33 B 0.049652f
C346 VN.n34 B 0.045798f
C347 VN.t6 B 0.579384f
C348 VN.n35 B 0.242825f
C349 VN.n36 B 0.039919f
C350 VN.n37 B 0.024573f
C351 VN.n38 B 0.024573f
C352 VN.n39 B 0.024573f
C353 VN.n40 B 0.045798f
C354 VN.n41 B 0.045798f
C355 VN.n42 B 0.03964f
C356 VN.n43 B 0.024573f
C357 VN.n44 B 0.024573f
C358 VN.n45 B 0.024573f
C359 VN.n46 B 0.045798f
C360 VN.n47 B 0.045798f
C361 VN.n48 B 0.03404f
C362 VN.n49 B 0.03966f
C363 VN.n50 B 0.064858f
C364 VN.t2 B 0.579384f
C365 VN.n51 B 0.341249f
C366 VN.n52 B 0.024573f
C367 VN.n53 B 0.032108f
C368 VN.n54 B 0.024573f
C369 VN.n55 B 0.029066f
C370 VN.n56 B 0.024573f
C371 VN.t3 B 0.579384f
C372 VN.n57 B 0.242825f
C373 VN.n58 B 0.021232f
C374 VN.n59 B 0.024573f
C375 VN.t7 B 0.579384f
C376 VN.n60 B 0.266012f
C377 VN.n61 B 0.024573f
C378 VN.n62 B 0.021232f
C379 VN.n63 B 0.024573f
C380 VN.t9 B 0.579384f
C381 VN.n64 B 0.333683f
C382 VN.t8 B 0.856714f
C383 VN.n65 B 0.341503f
C384 VN.n66 B 0.303984f
C385 VN.n67 B 0.039919f
C386 VN.n68 B 0.045798f
C387 VN.n69 B 0.049652f
C388 VN.n70 B 0.024573f
C389 VN.n71 B 0.024573f
C390 VN.n72 B 0.024573f
C391 VN.n73 B 0.046661f
C392 VN.n74 B 0.045798f
C393 VN.n75 B 0.045798f
C394 VN.n76 B 0.024573f
C395 VN.n77 B 0.024573f
C396 VN.n78 B 0.024573f
C397 VN.n79 B 0.045798f
C398 VN.n80 B 0.045798f
C399 VN.n81 B 0.046661f
C400 VN.n82 B 0.024573f
C401 VN.n83 B 0.024573f
C402 VN.n84 B 0.024573f
C403 VN.n85 B 0.049652f
C404 VN.n86 B 0.045798f
C405 VN.n87 B 0.039919f
C406 VN.n88 B 0.024573f
C407 VN.n89 B 0.024573f
C408 VN.n90 B 0.024573f
C409 VN.n91 B 0.045798f
C410 VN.n92 B 0.045798f
C411 VN.n93 B 0.03964f
C412 VN.n94 B 0.024573f
C413 VN.n95 B 0.024573f
C414 VN.n96 B 0.024573f
C415 VN.n97 B 0.045798f
C416 VN.n98 B 0.045798f
C417 VN.n99 B 0.03404f
C418 VN.n100 B 0.03966f
C419 VN.n101 B 1.46713f
.ends

