* NGSPICE file created from diff_pair_sample_0916.ext - technology: sky130A

.subckt diff_pair_sample_0916 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=0 ps=0 w=18.96 l=1.89
X1 VDD1.t5 VP.t0 VTAIL.t8 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=3.1284 ps=19.29 w=18.96 l=1.89
X2 VDD1.t4 VP.t1 VTAIL.t5 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=3.1284 ps=19.29 w=18.96 l=1.89
X3 VDD2.t5 VN.t0 VTAIL.t11 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=7.3944 ps=38.7 w=18.96 l=1.89
X4 VDD1.t3 VP.t2 VTAIL.t4 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=7.3944 ps=38.7 w=18.96 l=1.89
X5 VDD1.t2 VP.t3 VTAIL.t9 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=7.3944 ps=38.7 w=18.96 l=1.89
X6 B.t8 B.t6 B.t7 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=0 ps=0 w=18.96 l=1.89
X7 VDD2.t4 VN.t1 VTAIL.t0 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=7.3944 ps=38.7 w=18.96 l=1.89
X8 VDD2.t3 VN.t2 VTAIL.t1 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=3.1284 ps=19.29 w=18.96 l=1.89
X9 VDD2.t2 VN.t3 VTAIL.t2 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=3.1284 ps=19.29 w=18.96 l=1.89
X10 VTAIL.t7 VP.t4 VDD1.t1 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=3.1284 ps=19.29 w=18.96 l=1.89
X11 B.t5 B.t3 B.t4 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=0 ps=0 w=18.96 l=1.89
X12 VTAIL.t6 VP.t5 VDD1.t0 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=3.1284 ps=19.29 w=18.96 l=1.89
X13 VTAIL.t3 VN.t4 VDD2.t1 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=3.1284 ps=19.29 w=18.96 l=1.89
X14 VTAIL.t10 VN.t5 VDD2.t0 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=3.1284 pd=19.29 as=3.1284 ps=19.29 w=18.96 l=1.89
X15 B.t2 B.t0 B.t1 w_n2746_n4760# sky130_fd_pr__pfet_01v8 ad=7.3944 pd=38.7 as=0 ps=0 w=18.96 l=1.89
R0 B.n569 B.n90 585
R1 B.n571 B.n570 585
R2 B.n572 B.n89 585
R3 B.n574 B.n573 585
R4 B.n575 B.n88 585
R5 B.n577 B.n576 585
R6 B.n578 B.n87 585
R7 B.n580 B.n579 585
R8 B.n581 B.n86 585
R9 B.n583 B.n582 585
R10 B.n584 B.n85 585
R11 B.n586 B.n585 585
R12 B.n587 B.n84 585
R13 B.n589 B.n588 585
R14 B.n590 B.n83 585
R15 B.n592 B.n591 585
R16 B.n593 B.n82 585
R17 B.n595 B.n594 585
R18 B.n596 B.n81 585
R19 B.n598 B.n597 585
R20 B.n599 B.n80 585
R21 B.n601 B.n600 585
R22 B.n602 B.n79 585
R23 B.n604 B.n603 585
R24 B.n605 B.n78 585
R25 B.n607 B.n606 585
R26 B.n608 B.n77 585
R27 B.n610 B.n609 585
R28 B.n611 B.n76 585
R29 B.n613 B.n612 585
R30 B.n614 B.n75 585
R31 B.n616 B.n615 585
R32 B.n617 B.n74 585
R33 B.n619 B.n618 585
R34 B.n620 B.n73 585
R35 B.n622 B.n621 585
R36 B.n623 B.n72 585
R37 B.n625 B.n624 585
R38 B.n626 B.n71 585
R39 B.n628 B.n627 585
R40 B.n629 B.n70 585
R41 B.n631 B.n630 585
R42 B.n632 B.n69 585
R43 B.n634 B.n633 585
R44 B.n635 B.n68 585
R45 B.n637 B.n636 585
R46 B.n638 B.n67 585
R47 B.n640 B.n639 585
R48 B.n641 B.n66 585
R49 B.n643 B.n642 585
R50 B.n644 B.n65 585
R51 B.n646 B.n645 585
R52 B.n647 B.n64 585
R53 B.n649 B.n648 585
R54 B.n650 B.n63 585
R55 B.n652 B.n651 585
R56 B.n653 B.n62 585
R57 B.n655 B.n654 585
R58 B.n656 B.n61 585
R59 B.n658 B.n657 585
R60 B.n659 B.n60 585
R61 B.n661 B.n660 585
R62 B.n663 B.n57 585
R63 B.n665 B.n664 585
R64 B.n666 B.n56 585
R65 B.n668 B.n667 585
R66 B.n669 B.n55 585
R67 B.n671 B.n670 585
R68 B.n672 B.n54 585
R69 B.n674 B.n673 585
R70 B.n675 B.n53 585
R71 B.n677 B.n676 585
R72 B.n679 B.n678 585
R73 B.n680 B.n49 585
R74 B.n682 B.n681 585
R75 B.n683 B.n48 585
R76 B.n685 B.n684 585
R77 B.n686 B.n47 585
R78 B.n688 B.n687 585
R79 B.n689 B.n46 585
R80 B.n691 B.n690 585
R81 B.n692 B.n45 585
R82 B.n694 B.n693 585
R83 B.n695 B.n44 585
R84 B.n697 B.n696 585
R85 B.n698 B.n43 585
R86 B.n700 B.n699 585
R87 B.n701 B.n42 585
R88 B.n703 B.n702 585
R89 B.n704 B.n41 585
R90 B.n706 B.n705 585
R91 B.n707 B.n40 585
R92 B.n709 B.n708 585
R93 B.n710 B.n39 585
R94 B.n712 B.n711 585
R95 B.n713 B.n38 585
R96 B.n715 B.n714 585
R97 B.n716 B.n37 585
R98 B.n718 B.n717 585
R99 B.n719 B.n36 585
R100 B.n721 B.n720 585
R101 B.n722 B.n35 585
R102 B.n724 B.n723 585
R103 B.n725 B.n34 585
R104 B.n727 B.n726 585
R105 B.n728 B.n33 585
R106 B.n730 B.n729 585
R107 B.n731 B.n32 585
R108 B.n733 B.n732 585
R109 B.n734 B.n31 585
R110 B.n736 B.n735 585
R111 B.n737 B.n30 585
R112 B.n739 B.n738 585
R113 B.n740 B.n29 585
R114 B.n742 B.n741 585
R115 B.n743 B.n28 585
R116 B.n745 B.n744 585
R117 B.n746 B.n27 585
R118 B.n748 B.n747 585
R119 B.n749 B.n26 585
R120 B.n751 B.n750 585
R121 B.n752 B.n25 585
R122 B.n754 B.n753 585
R123 B.n755 B.n24 585
R124 B.n757 B.n756 585
R125 B.n758 B.n23 585
R126 B.n760 B.n759 585
R127 B.n761 B.n22 585
R128 B.n763 B.n762 585
R129 B.n764 B.n21 585
R130 B.n766 B.n765 585
R131 B.n767 B.n20 585
R132 B.n769 B.n768 585
R133 B.n770 B.n19 585
R134 B.n568 B.n567 585
R135 B.n566 B.n91 585
R136 B.n565 B.n564 585
R137 B.n563 B.n92 585
R138 B.n562 B.n561 585
R139 B.n560 B.n93 585
R140 B.n559 B.n558 585
R141 B.n557 B.n94 585
R142 B.n556 B.n555 585
R143 B.n554 B.n95 585
R144 B.n553 B.n552 585
R145 B.n551 B.n96 585
R146 B.n550 B.n549 585
R147 B.n548 B.n97 585
R148 B.n547 B.n546 585
R149 B.n545 B.n98 585
R150 B.n544 B.n543 585
R151 B.n542 B.n99 585
R152 B.n541 B.n540 585
R153 B.n539 B.n100 585
R154 B.n538 B.n537 585
R155 B.n536 B.n101 585
R156 B.n535 B.n534 585
R157 B.n533 B.n102 585
R158 B.n532 B.n531 585
R159 B.n530 B.n103 585
R160 B.n529 B.n528 585
R161 B.n527 B.n104 585
R162 B.n526 B.n525 585
R163 B.n524 B.n105 585
R164 B.n523 B.n522 585
R165 B.n521 B.n106 585
R166 B.n520 B.n519 585
R167 B.n518 B.n107 585
R168 B.n517 B.n516 585
R169 B.n515 B.n108 585
R170 B.n514 B.n513 585
R171 B.n512 B.n109 585
R172 B.n511 B.n510 585
R173 B.n509 B.n110 585
R174 B.n508 B.n507 585
R175 B.n506 B.n111 585
R176 B.n505 B.n504 585
R177 B.n503 B.n112 585
R178 B.n502 B.n501 585
R179 B.n500 B.n113 585
R180 B.n499 B.n498 585
R181 B.n497 B.n114 585
R182 B.n496 B.n495 585
R183 B.n494 B.n115 585
R184 B.n493 B.n492 585
R185 B.n491 B.n116 585
R186 B.n490 B.n489 585
R187 B.n488 B.n117 585
R188 B.n487 B.n486 585
R189 B.n485 B.n118 585
R190 B.n484 B.n483 585
R191 B.n482 B.n119 585
R192 B.n481 B.n480 585
R193 B.n479 B.n120 585
R194 B.n478 B.n477 585
R195 B.n476 B.n121 585
R196 B.n475 B.n474 585
R197 B.n473 B.n122 585
R198 B.n472 B.n471 585
R199 B.n470 B.n123 585
R200 B.n469 B.n468 585
R201 B.n467 B.n124 585
R202 B.n466 B.n465 585
R203 B.n263 B.n196 585
R204 B.n265 B.n264 585
R205 B.n266 B.n195 585
R206 B.n268 B.n267 585
R207 B.n269 B.n194 585
R208 B.n271 B.n270 585
R209 B.n272 B.n193 585
R210 B.n274 B.n273 585
R211 B.n275 B.n192 585
R212 B.n277 B.n276 585
R213 B.n278 B.n191 585
R214 B.n280 B.n279 585
R215 B.n281 B.n190 585
R216 B.n283 B.n282 585
R217 B.n284 B.n189 585
R218 B.n286 B.n285 585
R219 B.n287 B.n188 585
R220 B.n289 B.n288 585
R221 B.n290 B.n187 585
R222 B.n292 B.n291 585
R223 B.n293 B.n186 585
R224 B.n295 B.n294 585
R225 B.n296 B.n185 585
R226 B.n298 B.n297 585
R227 B.n299 B.n184 585
R228 B.n301 B.n300 585
R229 B.n302 B.n183 585
R230 B.n304 B.n303 585
R231 B.n305 B.n182 585
R232 B.n307 B.n306 585
R233 B.n308 B.n181 585
R234 B.n310 B.n309 585
R235 B.n311 B.n180 585
R236 B.n313 B.n312 585
R237 B.n314 B.n179 585
R238 B.n316 B.n315 585
R239 B.n317 B.n178 585
R240 B.n319 B.n318 585
R241 B.n320 B.n177 585
R242 B.n322 B.n321 585
R243 B.n323 B.n176 585
R244 B.n325 B.n324 585
R245 B.n326 B.n175 585
R246 B.n328 B.n327 585
R247 B.n329 B.n174 585
R248 B.n331 B.n330 585
R249 B.n332 B.n173 585
R250 B.n334 B.n333 585
R251 B.n335 B.n172 585
R252 B.n337 B.n336 585
R253 B.n338 B.n171 585
R254 B.n340 B.n339 585
R255 B.n341 B.n170 585
R256 B.n343 B.n342 585
R257 B.n344 B.n169 585
R258 B.n346 B.n345 585
R259 B.n347 B.n168 585
R260 B.n349 B.n348 585
R261 B.n350 B.n167 585
R262 B.n352 B.n351 585
R263 B.n353 B.n166 585
R264 B.n355 B.n354 585
R265 B.n357 B.n163 585
R266 B.n359 B.n358 585
R267 B.n360 B.n162 585
R268 B.n362 B.n361 585
R269 B.n363 B.n161 585
R270 B.n365 B.n364 585
R271 B.n366 B.n160 585
R272 B.n368 B.n367 585
R273 B.n369 B.n159 585
R274 B.n371 B.n370 585
R275 B.n373 B.n372 585
R276 B.n374 B.n155 585
R277 B.n376 B.n375 585
R278 B.n377 B.n154 585
R279 B.n379 B.n378 585
R280 B.n380 B.n153 585
R281 B.n382 B.n381 585
R282 B.n383 B.n152 585
R283 B.n385 B.n384 585
R284 B.n386 B.n151 585
R285 B.n388 B.n387 585
R286 B.n389 B.n150 585
R287 B.n391 B.n390 585
R288 B.n392 B.n149 585
R289 B.n394 B.n393 585
R290 B.n395 B.n148 585
R291 B.n397 B.n396 585
R292 B.n398 B.n147 585
R293 B.n400 B.n399 585
R294 B.n401 B.n146 585
R295 B.n403 B.n402 585
R296 B.n404 B.n145 585
R297 B.n406 B.n405 585
R298 B.n407 B.n144 585
R299 B.n409 B.n408 585
R300 B.n410 B.n143 585
R301 B.n412 B.n411 585
R302 B.n413 B.n142 585
R303 B.n415 B.n414 585
R304 B.n416 B.n141 585
R305 B.n418 B.n417 585
R306 B.n419 B.n140 585
R307 B.n421 B.n420 585
R308 B.n422 B.n139 585
R309 B.n424 B.n423 585
R310 B.n425 B.n138 585
R311 B.n427 B.n426 585
R312 B.n428 B.n137 585
R313 B.n430 B.n429 585
R314 B.n431 B.n136 585
R315 B.n433 B.n432 585
R316 B.n434 B.n135 585
R317 B.n436 B.n435 585
R318 B.n437 B.n134 585
R319 B.n439 B.n438 585
R320 B.n440 B.n133 585
R321 B.n442 B.n441 585
R322 B.n443 B.n132 585
R323 B.n445 B.n444 585
R324 B.n446 B.n131 585
R325 B.n448 B.n447 585
R326 B.n449 B.n130 585
R327 B.n451 B.n450 585
R328 B.n452 B.n129 585
R329 B.n454 B.n453 585
R330 B.n455 B.n128 585
R331 B.n457 B.n456 585
R332 B.n458 B.n127 585
R333 B.n460 B.n459 585
R334 B.n461 B.n126 585
R335 B.n463 B.n462 585
R336 B.n464 B.n125 585
R337 B.n262 B.n261 585
R338 B.n260 B.n197 585
R339 B.n259 B.n258 585
R340 B.n257 B.n198 585
R341 B.n256 B.n255 585
R342 B.n254 B.n199 585
R343 B.n253 B.n252 585
R344 B.n251 B.n200 585
R345 B.n250 B.n249 585
R346 B.n248 B.n201 585
R347 B.n247 B.n246 585
R348 B.n245 B.n202 585
R349 B.n244 B.n243 585
R350 B.n242 B.n203 585
R351 B.n241 B.n240 585
R352 B.n239 B.n204 585
R353 B.n238 B.n237 585
R354 B.n236 B.n205 585
R355 B.n235 B.n234 585
R356 B.n233 B.n206 585
R357 B.n232 B.n231 585
R358 B.n230 B.n207 585
R359 B.n229 B.n228 585
R360 B.n227 B.n208 585
R361 B.n226 B.n225 585
R362 B.n224 B.n209 585
R363 B.n223 B.n222 585
R364 B.n221 B.n210 585
R365 B.n220 B.n219 585
R366 B.n218 B.n211 585
R367 B.n217 B.n216 585
R368 B.n215 B.n212 585
R369 B.n214 B.n213 585
R370 B.n2 B.n0 585
R371 B.n821 B.n1 585
R372 B.n820 B.n819 585
R373 B.n818 B.n3 585
R374 B.n817 B.n816 585
R375 B.n815 B.n4 585
R376 B.n814 B.n813 585
R377 B.n812 B.n5 585
R378 B.n811 B.n810 585
R379 B.n809 B.n6 585
R380 B.n808 B.n807 585
R381 B.n806 B.n7 585
R382 B.n805 B.n804 585
R383 B.n803 B.n8 585
R384 B.n802 B.n801 585
R385 B.n800 B.n9 585
R386 B.n799 B.n798 585
R387 B.n797 B.n10 585
R388 B.n796 B.n795 585
R389 B.n794 B.n11 585
R390 B.n793 B.n792 585
R391 B.n791 B.n12 585
R392 B.n790 B.n789 585
R393 B.n788 B.n13 585
R394 B.n787 B.n786 585
R395 B.n785 B.n14 585
R396 B.n784 B.n783 585
R397 B.n782 B.n15 585
R398 B.n781 B.n780 585
R399 B.n779 B.n16 585
R400 B.n778 B.n777 585
R401 B.n776 B.n17 585
R402 B.n775 B.n774 585
R403 B.n773 B.n18 585
R404 B.n772 B.n771 585
R405 B.n823 B.n822 585
R406 B.n156 B.t8 544.168
R407 B.n58 B.t1 544.168
R408 B.n164 B.t5 544.168
R409 B.n50 B.t10 544.168
R410 B.n263 B.n262 516.524
R411 B.n772 B.n19 516.524
R412 B.n466 B.n125 516.524
R413 B.n569 B.n568 516.524
R414 B.n157 B.t7 501.113
R415 B.n59 B.t2 501.113
R416 B.n165 B.t4 501.113
R417 B.n51 B.t11 501.113
R418 B.n156 B.t6 448.413
R419 B.n164 B.t3 448.413
R420 B.n50 B.t9 448.413
R421 B.n58 B.t0 448.413
R422 B.n262 B.n197 163.367
R423 B.n258 B.n197 163.367
R424 B.n258 B.n257 163.367
R425 B.n257 B.n256 163.367
R426 B.n256 B.n199 163.367
R427 B.n252 B.n199 163.367
R428 B.n252 B.n251 163.367
R429 B.n251 B.n250 163.367
R430 B.n250 B.n201 163.367
R431 B.n246 B.n201 163.367
R432 B.n246 B.n245 163.367
R433 B.n245 B.n244 163.367
R434 B.n244 B.n203 163.367
R435 B.n240 B.n203 163.367
R436 B.n240 B.n239 163.367
R437 B.n239 B.n238 163.367
R438 B.n238 B.n205 163.367
R439 B.n234 B.n205 163.367
R440 B.n234 B.n233 163.367
R441 B.n233 B.n232 163.367
R442 B.n232 B.n207 163.367
R443 B.n228 B.n207 163.367
R444 B.n228 B.n227 163.367
R445 B.n227 B.n226 163.367
R446 B.n226 B.n209 163.367
R447 B.n222 B.n209 163.367
R448 B.n222 B.n221 163.367
R449 B.n221 B.n220 163.367
R450 B.n220 B.n211 163.367
R451 B.n216 B.n211 163.367
R452 B.n216 B.n215 163.367
R453 B.n215 B.n214 163.367
R454 B.n214 B.n2 163.367
R455 B.n822 B.n2 163.367
R456 B.n822 B.n821 163.367
R457 B.n821 B.n820 163.367
R458 B.n820 B.n3 163.367
R459 B.n816 B.n3 163.367
R460 B.n816 B.n815 163.367
R461 B.n815 B.n814 163.367
R462 B.n814 B.n5 163.367
R463 B.n810 B.n5 163.367
R464 B.n810 B.n809 163.367
R465 B.n809 B.n808 163.367
R466 B.n808 B.n7 163.367
R467 B.n804 B.n7 163.367
R468 B.n804 B.n803 163.367
R469 B.n803 B.n802 163.367
R470 B.n802 B.n9 163.367
R471 B.n798 B.n9 163.367
R472 B.n798 B.n797 163.367
R473 B.n797 B.n796 163.367
R474 B.n796 B.n11 163.367
R475 B.n792 B.n11 163.367
R476 B.n792 B.n791 163.367
R477 B.n791 B.n790 163.367
R478 B.n790 B.n13 163.367
R479 B.n786 B.n13 163.367
R480 B.n786 B.n785 163.367
R481 B.n785 B.n784 163.367
R482 B.n784 B.n15 163.367
R483 B.n780 B.n15 163.367
R484 B.n780 B.n779 163.367
R485 B.n779 B.n778 163.367
R486 B.n778 B.n17 163.367
R487 B.n774 B.n17 163.367
R488 B.n774 B.n773 163.367
R489 B.n773 B.n772 163.367
R490 B.n264 B.n263 163.367
R491 B.n264 B.n195 163.367
R492 B.n268 B.n195 163.367
R493 B.n269 B.n268 163.367
R494 B.n270 B.n269 163.367
R495 B.n270 B.n193 163.367
R496 B.n274 B.n193 163.367
R497 B.n275 B.n274 163.367
R498 B.n276 B.n275 163.367
R499 B.n276 B.n191 163.367
R500 B.n280 B.n191 163.367
R501 B.n281 B.n280 163.367
R502 B.n282 B.n281 163.367
R503 B.n282 B.n189 163.367
R504 B.n286 B.n189 163.367
R505 B.n287 B.n286 163.367
R506 B.n288 B.n287 163.367
R507 B.n288 B.n187 163.367
R508 B.n292 B.n187 163.367
R509 B.n293 B.n292 163.367
R510 B.n294 B.n293 163.367
R511 B.n294 B.n185 163.367
R512 B.n298 B.n185 163.367
R513 B.n299 B.n298 163.367
R514 B.n300 B.n299 163.367
R515 B.n300 B.n183 163.367
R516 B.n304 B.n183 163.367
R517 B.n305 B.n304 163.367
R518 B.n306 B.n305 163.367
R519 B.n306 B.n181 163.367
R520 B.n310 B.n181 163.367
R521 B.n311 B.n310 163.367
R522 B.n312 B.n311 163.367
R523 B.n312 B.n179 163.367
R524 B.n316 B.n179 163.367
R525 B.n317 B.n316 163.367
R526 B.n318 B.n317 163.367
R527 B.n318 B.n177 163.367
R528 B.n322 B.n177 163.367
R529 B.n323 B.n322 163.367
R530 B.n324 B.n323 163.367
R531 B.n324 B.n175 163.367
R532 B.n328 B.n175 163.367
R533 B.n329 B.n328 163.367
R534 B.n330 B.n329 163.367
R535 B.n330 B.n173 163.367
R536 B.n334 B.n173 163.367
R537 B.n335 B.n334 163.367
R538 B.n336 B.n335 163.367
R539 B.n336 B.n171 163.367
R540 B.n340 B.n171 163.367
R541 B.n341 B.n340 163.367
R542 B.n342 B.n341 163.367
R543 B.n342 B.n169 163.367
R544 B.n346 B.n169 163.367
R545 B.n347 B.n346 163.367
R546 B.n348 B.n347 163.367
R547 B.n348 B.n167 163.367
R548 B.n352 B.n167 163.367
R549 B.n353 B.n352 163.367
R550 B.n354 B.n353 163.367
R551 B.n354 B.n163 163.367
R552 B.n359 B.n163 163.367
R553 B.n360 B.n359 163.367
R554 B.n361 B.n360 163.367
R555 B.n361 B.n161 163.367
R556 B.n365 B.n161 163.367
R557 B.n366 B.n365 163.367
R558 B.n367 B.n366 163.367
R559 B.n367 B.n159 163.367
R560 B.n371 B.n159 163.367
R561 B.n372 B.n371 163.367
R562 B.n372 B.n155 163.367
R563 B.n376 B.n155 163.367
R564 B.n377 B.n376 163.367
R565 B.n378 B.n377 163.367
R566 B.n378 B.n153 163.367
R567 B.n382 B.n153 163.367
R568 B.n383 B.n382 163.367
R569 B.n384 B.n383 163.367
R570 B.n384 B.n151 163.367
R571 B.n388 B.n151 163.367
R572 B.n389 B.n388 163.367
R573 B.n390 B.n389 163.367
R574 B.n390 B.n149 163.367
R575 B.n394 B.n149 163.367
R576 B.n395 B.n394 163.367
R577 B.n396 B.n395 163.367
R578 B.n396 B.n147 163.367
R579 B.n400 B.n147 163.367
R580 B.n401 B.n400 163.367
R581 B.n402 B.n401 163.367
R582 B.n402 B.n145 163.367
R583 B.n406 B.n145 163.367
R584 B.n407 B.n406 163.367
R585 B.n408 B.n407 163.367
R586 B.n408 B.n143 163.367
R587 B.n412 B.n143 163.367
R588 B.n413 B.n412 163.367
R589 B.n414 B.n413 163.367
R590 B.n414 B.n141 163.367
R591 B.n418 B.n141 163.367
R592 B.n419 B.n418 163.367
R593 B.n420 B.n419 163.367
R594 B.n420 B.n139 163.367
R595 B.n424 B.n139 163.367
R596 B.n425 B.n424 163.367
R597 B.n426 B.n425 163.367
R598 B.n426 B.n137 163.367
R599 B.n430 B.n137 163.367
R600 B.n431 B.n430 163.367
R601 B.n432 B.n431 163.367
R602 B.n432 B.n135 163.367
R603 B.n436 B.n135 163.367
R604 B.n437 B.n436 163.367
R605 B.n438 B.n437 163.367
R606 B.n438 B.n133 163.367
R607 B.n442 B.n133 163.367
R608 B.n443 B.n442 163.367
R609 B.n444 B.n443 163.367
R610 B.n444 B.n131 163.367
R611 B.n448 B.n131 163.367
R612 B.n449 B.n448 163.367
R613 B.n450 B.n449 163.367
R614 B.n450 B.n129 163.367
R615 B.n454 B.n129 163.367
R616 B.n455 B.n454 163.367
R617 B.n456 B.n455 163.367
R618 B.n456 B.n127 163.367
R619 B.n460 B.n127 163.367
R620 B.n461 B.n460 163.367
R621 B.n462 B.n461 163.367
R622 B.n462 B.n125 163.367
R623 B.n467 B.n466 163.367
R624 B.n468 B.n467 163.367
R625 B.n468 B.n123 163.367
R626 B.n472 B.n123 163.367
R627 B.n473 B.n472 163.367
R628 B.n474 B.n473 163.367
R629 B.n474 B.n121 163.367
R630 B.n478 B.n121 163.367
R631 B.n479 B.n478 163.367
R632 B.n480 B.n479 163.367
R633 B.n480 B.n119 163.367
R634 B.n484 B.n119 163.367
R635 B.n485 B.n484 163.367
R636 B.n486 B.n485 163.367
R637 B.n486 B.n117 163.367
R638 B.n490 B.n117 163.367
R639 B.n491 B.n490 163.367
R640 B.n492 B.n491 163.367
R641 B.n492 B.n115 163.367
R642 B.n496 B.n115 163.367
R643 B.n497 B.n496 163.367
R644 B.n498 B.n497 163.367
R645 B.n498 B.n113 163.367
R646 B.n502 B.n113 163.367
R647 B.n503 B.n502 163.367
R648 B.n504 B.n503 163.367
R649 B.n504 B.n111 163.367
R650 B.n508 B.n111 163.367
R651 B.n509 B.n508 163.367
R652 B.n510 B.n509 163.367
R653 B.n510 B.n109 163.367
R654 B.n514 B.n109 163.367
R655 B.n515 B.n514 163.367
R656 B.n516 B.n515 163.367
R657 B.n516 B.n107 163.367
R658 B.n520 B.n107 163.367
R659 B.n521 B.n520 163.367
R660 B.n522 B.n521 163.367
R661 B.n522 B.n105 163.367
R662 B.n526 B.n105 163.367
R663 B.n527 B.n526 163.367
R664 B.n528 B.n527 163.367
R665 B.n528 B.n103 163.367
R666 B.n532 B.n103 163.367
R667 B.n533 B.n532 163.367
R668 B.n534 B.n533 163.367
R669 B.n534 B.n101 163.367
R670 B.n538 B.n101 163.367
R671 B.n539 B.n538 163.367
R672 B.n540 B.n539 163.367
R673 B.n540 B.n99 163.367
R674 B.n544 B.n99 163.367
R675 B.n545 B.n544 163.367
R676 B.n546 B.n545 163.367
R677 B.n546 B.n97 163.367
R678 B.n550 B.n97 163.367
R679 B.n551 B.n550 163.367
R680 B.n552 B.n551 163.367
R681 B.n552 B.n95 163.367
R682 B.n556 B.n95 163.367
R683 B.n557 B.n556 163.367
R684 B.n558 B.n557 163.367
R685 B.n558 B.n93 163.367
R686 B.n562 B.n93 163.367
R687 B.n563 B.n562 163.367
R688 B.n564 B.n563 163.367
R689 B.n564 B.n91 163.367
R690 B.n568 B.n91 163.367
R691 B.n768 B.n19 163.367
R692 B.n768 B.n767 163.367
R693 B.n767 B.n766 163.367
R694 B.n766 B.n21 163.367
R695 B.n762 B.n21 163.367
R696 B.n762 B.n761 163.367
R697 B.n761 B.n760 163.367
R698 B.n760 B.n23 163.367
R699 B.n756 B.n23 163.367
R700 B.n756 B.n755 163.367
R701 B.n755 B.n754 163.367
R702 B.n754 B.n25 163.367
R703 B.n750 B.n25 163.367
R704 B.n750 B.n749 163.367
R705 B.n749 B.n748 163.367
R706 B.n748 B.n27 163.367
R707 B.n744 B.n27 163.367
R708 B.n744 B.n743 163.367
R709 B.n743 B.n742 163.367
R710 B.n742 B.n29 163.367
R711 B.n738 B.n29 163.367
R712 B.n738 B.n737 163.367
R713 B.n737 B.n736 163.367
R714 B.n736 B.n31 163.367
R715 B.n732 B.n31 163.367
R716 B.n732 B.n731 163.367
R717 B.n731 B.n730 163.367
R718 B.n730 B.n33 163.367
R719 B.n726 B.n33 163.367
R720 B.n726 B.n725 163.367
R721 B.n725 B.n724 163.367
R722 B.n724 B.n35 163.367
R723 B.n720 B.n35 163.367
R724 B.n720 B.n719 163.367
R725 B.n719 B.n718 163.367
R726 B.n718 B.n37 163.367
R727 B.n714 B.n37 163.367
R728 B.n714 B.n713 163.367
R729 B.n713 B.n712 163.367
R730 B.n712 B.n39 163.367
R731 B.n708 B.n39 163.367
R732 B.n708 B.n707 163.367
R733 B.n707 B.n706 163.367
R734 B.n706 B.n41 163.367
R735 B.n702 B.n41 163.367
R736 B.n702 B.n701 163.367
R737 B.n701 B.n700 163.367
R738 B.n700 B.n43 163.367
R739 B.n696 B.n43 163.367
R740 B.n696 B.n695 163.367
R741 B.n695 B.n694 163.367
R742 B.n694 B.n45 163.367
R743 B.n690 B.n45 163.367
R744 B.n690 B.n689 163.367
R745 B.n689 B.n688 163.367
R746 B.n688 B.n47 163.367
R747 B.n684 B.n47 163.367
R748 B.n684 B.n683 163.367
R749 B.n683 B.n682 163.367
R750 B.n682 B.n49 163.367
R751 B.n678 B.n49 163.367
R752 B.n678 B.n677 163.367
R753 B.n677 B.n53 163.367
R754 B.n673 B.n53 163.367
R755 B.n673 B.n672 163.367
R756 B.n672 B.n671 163.367
R757 B.n671 B.n55 163.367
R758 B.n667 B.n55 163.367
R759 B.n667 B.n666 163.367
R760 B.n666 B.n665 163.367
R761 B.n665 B.n57 163.367
R762 B.n660 B.n57 163.367
R763 B.n660 B.n659 163.367
R764 B.n659 B.n658 163.367
R765 B.n658 B.n61 163.367
R766 B.n654 B.n61 163.367
R767 B.n654 B.n653 163.367
R768 B.n653 B.n652 163.367
R769 B.n652 B.n63 163.367
R770 B.n648 B.n63 163.367
R771 B.n648 B.n647 163.367
R772 B.n647 B.n646 163.367
R773 B.n646 B.n65 163.367
R774 B.n642 B.n65 163.367
R775 B.n642 B.n641 163.367
R776 B.n641 B.n640 163.367
R777 B.n640 B.n67 163.367
R778 B.n636 B.n67 163.367
R779 B.n636 B.n635 163.367
R780 B.n635 B.n634 163.367
R781 B.n634 B.n69 163.367
R782 B.n630 B.n69 163.367
R783 B.n630 B.n629 163.367
R784 B.n629 B.n628 163.367
R785 B.n628 B.n71 163.367
R786 B.n624 B.n71 163.367
R787 B.n624 B.n623 163.367
R788 B.n623 B.n622 163.367
R789 B.n622 B.n73 163.367
R790 B.n618 B.n73 163.367
R791 B.n618 B.n617 163.367
R792 B.n617 B.n616 163.367
R793 B.n616 B.n75 163.367
R794 B.n612 B.n75 163.367
R795 B.n612 B.n611 163.367
R796 B.n611 B.n610 163.367
R797 B.n610 B.n77 163.367
R798 B.n606 B.n77 163.367
R799 B.n606 B.n605 163.367
R800 B.n605 B.n604 163.367
R801 B.n604 B.n79 163.367
R802 B.n600 B.n79 163.367
R803 B.n600 B.n599 163.367
R804 B.n599 B.n598 163.367
R805 B.n598 B.n81 163.367
R806 B.n594 B.n81 163.367
R807 B.n594 B.n593 163.367
R808 B.n593 B.n592 163.367
R809 B.n592 B.n83 163.367
R810 B.n588 B.n83 163.367
R811 B.n588 B.n587 163.367
R812 B.n587 B.n586 163.367
R813 B.n586 B.n85 163.367
R814 B.n582 B.n85 163.367
R815 B.n582 B.n581 163.367
R816 B.n581 B.n580 163.367
R817 B.n580 B.n87 163.367
R818 B.n576 B.n87 163.367
R819 B.n576 B.n575 163.367
R820 B.n575 B.n574 163.367
R821 B.n574 B.n89 163.367
R822 B.n570 B.n89 163.367
R823 B.n570 B.n569 163.367
R824 B.n158 B.n157 59.5399
R825 B.n356 B.n165 59.5399
R826 B.n52 B.n51 59.5399
R827 B.n662 B.n59 59.5399
R828 B.n157 B.n156 43.055
R829 B.n165 B.n164 43.055
R830 B.n51 B.n50 43.055
R831 B.n59 B.n58 43.055
R832 B.n771 B.n770 33.5615
R833 B.n567 B.n90 33.5615
R834 B.n465 B.n464 33.5615
R835 B.n261 B.n196 33.5615
R836 B B.n823 18.0485
R837 B.n770 B.n769 10.6151
R838 B.n769 B.n20 10.6151
R839 B.n765 B.n20 10.6151
R840 B.n765 B.n764 10.6151
R841 B.n764 B.n763 10.6151
R842 B.n763 B.n22 10.6151
R843 B.n759 B.n22 10.6151
R844 B.n759 B.n758 10.6151
R845 B.n758 B.n757 10.6151
R846 B.n757 B.n24 10.6151
R847 B.n753 B.n24 10.6151
R848 B.n753 B.n752 10.6151
R849 B.n752 B.n751 10.6151
R850 B.n751 B.n26 10.6151
R851 B.n747 B.n26 10.6151
R852 B.n747 B.n746 10.6151
R853 B.n746 B.n745 10.6151
R854 B.n745 B.n28 10.6151
R855 B.n741 B.n28 10.6151
R856 B.n741 B.n740 10.6151
R857 B.n740 B.n739 10.6151
R858 B.n739 B.n30 10.6151
R859 B.n735 B.n30 10.6151
R860 B.n735 B.n734 10.6151
R861 B.n734 B.n733 10.6151
R862 B.n733 B.n32 10.6151
R863 B.n729 B.n32 10.6151
R864 B.n729 B.n728 10.6151
R865 B.n728 B.n727 10.6151
R866 B.n727 B.n34 10.6151
R867 B.n723 B.n34 10.6151
R868 B.n723 B.n722 10.6151
R869 B.n722 B.n721 10.6151
R870 B.n721 B.n36 10.6151
R871 B.n717 B.n36 10.6151
R872 B.n717 B.n716 10.6151
R873 B.n716 B.n715 10.6151
R874 B.n715 B.n38 10.6151
R875 B.n711 B.n38 10.6151
R876 B.n711 B.n710 10.6151
R877 B.n710 B.n709 10.6151
R878 B.n709 B.n40 10.6151
R879 B.n705 B.n40 10.6151
R880 B.n705 B.n704 10.6151
R881 B.n704 B.n703 10.6151
R882 B.n703 B.n42 10.6151
R883 B.n699 B.n42 10.6151
R884 B.n699 B.n698 10.6151
R885 B.n698 B.n697 10.6151
R886 B.n697 B.n44 10.6151
R887 B.n693 B.n44 10.6151
R888 B.n693 B.n692 10.6151
R889 B.n692 B.n691 10.6151
R890 B.n691 B.n46 10.6151
R891 B.n687 B.n46 10.6151
R892 B.n687 B.n686 10.6151
R893 B.n686 B.n685 10.6151
R894 B.n685 B.n48 10.6151
R895 B.n681 B.n48 10.6151
R896 B.n681 B.n680 10.6151
R897 B.n680 B.n679 10.6151
R898 B.n676 B.n675 10.6151
R899 B.n675 B.n674 10.6151
R900 B.n674 B.n54 10.6151
R901 B.n670 B.n54 10.6151
R902 B.n670 B.n669 10.6151
R903 B.n669 B.n668 10.6151
R904 B.n668 B.n56 10.6151
R905 B.n664 B.n56 10.6151
R906 B.n664 B.n663 10.6151
R907 B.n661 B.n60 10.6151
R908 B.n657 B.n60 10.6151
R909 B.n657 B.n656 10.6151
R910 B.n656 B.n655 10.6151
R911 B.n655 B.n62 10.6151
R912 B.n651 B.n62 10.6151
R913 B.n651 B.n650 10.6151
R914 B.n650 B.n649 10.6151
R915 B.n649 B.n64 10.6151
R916 B.n645 B.n64 10.6151
R917 B.n645 B.n644 10.6151
R918 B.n644 B.n643 10.6151
R919 B.n643 B.n66 10.6151
R920 B.n639 B.n66 10.6151
R921 B.n639 B.n638 10.6151
R922 B.n638 B.n637 10.6151
R923 B.n637 B.n68 10.6151
R924 B.n633 B.n68 10.6151
R925 B.n633 B.n632 10.6151
R926 B.n632 B.n631 10.6151
R927 B.n631 B.n70 10.6151
R928 B.n627 B.n70 10.6151
R929 B.n627 B.n626 10.6151
R930 B.n626 B.n625 10.6151
R931 B.n625 B.n72 10.6151
R932 B.n621 B.n72 10.6151
R933 B.n621 B.n620 10.6151
R934 B.n620 B.n619 10.6151
R935 B.n619 B.n74 10.6151
R936 B.n615 B.n74 10.6151
R937 B.n615 B.n614 10.6151
R938 B.n614 B.n613 10.6151
R939 B.n613 B.n76 10.6151
R940 B.n609 B.n76 10.6151
R941 B.n609 B.n608 10.6151
R942 B.n608 B.n607 10.6151
R943 B.n607 B.n78 10.6151
R944 B.n603 B.n78 10.6151
R945 B.n603 B.n602 10.6151
R946 B.n602 B.n601 10.6151
R947 B.n601 B.n80 10.6151
R948 B.n597 B.n80 10.6151
R949 B.n597 B.n596 10.6151
R950 B.n596 B.n595 10.6151
R951 B.n595 B.n82 10.6151
R952 B.n591 B.n82 10.6151
R953 B.n591 B.n590 10.6151
R954 B.n590 B.n589 10.6151
R955 B.n589 B.n84 10.6151
R956 B.n585 B.n84 10.6151
R957 B.n585 B.n584 10.6151
R958 B.n584 B.n583 10.6151
R959 B.n583 B.n86 10.6151
R960 B.n579 B.n86 10.6151
R961 B.n579 B.n578 10.6151
R962 B.n578 B.n577 10.6151
R963 B.n577 B.n88 10.6151
R964 B.n573 B.n88 10.6151
R965 B.n573 B.n572 10.6151
R966 B.n572 B.n571 10.6151
R967 B.n571 B.n90 10.6151
R968 B.n465 B.n124 10.6151
R969 B.n469 B.n124 10.6151
R970 B.n470 B.n469 10.6151
R971 B.n471 B.n470 10.6151
R972 B.n471 B.n122 10.6151
R973 B.n475 B.n122 10.6151
R974 B.n476 B.n475 10.6151
R975 B.n477 B.n476 10.6151
R976 B.n477 B.n120 10.6151
R977 B.n481 B.n120 10.6151
R978 B.n482 B.n481 10.6151
R979 B.n483 B.n482 10.6151
R980 B.n483 B.n118 10.6151
R981 B.n487 B.n118 10.6151
R982 B.n488 B.n487 10.6151
R983 B.n489 B.n488 10.6151
R984 B.n489 B.n116 10.6151
R985 B.n493 B.n116 10.6151
R986 B.n494 B.n493 10.6151
R987 B.n495 B.n494 10.6151
R988 B.n495 B.n114 10.6151
R989 B.n499 B.n114 10.6151
R990 B.n500 B.n499 10.6151
R991 B.n501 B.n500 10.6151
R992 B.n501 B.n112 10.6151
R993 B.n505 B.n112 10.6151
R994 B.n506 B.n505 10.6151
R995 B.n507 B.n506 10.6151
R996 B.n507 B.n110 10.6151
R997 B.n511 B.n110 10.6151
R998 B.n512 B.n511 10.6151
R999 B.n513 B.n512 10.6151
R1000 B.n513 B.n108 10.6151
R1001 B.n517 B.n108 10.6151
R1002 B.n518 B.n517 10.6151
R1003 B.n519 B.n518 10.6151
R1004 B.n519 B.n106 10.6151
R1005 B.n523 B.n106 10.6151
R1006 B.n524 B.n523 10.6151
R1007 B.n525 B.n524 10.6151
R1008 B.n525 B.n104 10.6151
R1009 B.n529 B.n104 10.6151
R1010 B.n530 B.n529 10.6151
R1011 B.n531 B.n530 10.6151
R1012 B.n531 B.n102 10.6151
R1013 B.n535 B.n102 10.6151
R1014 B.n536 B.n535 10.6151
R1015 B.n537 B.n536 10.6151
R1016 B.n537 B.n100 10.6151
R1017 B.n541 B.n100 10.6151
R1018 B.n542 B.n541 10.6151
R1019 B.n543 B.n542 10.6151
R1020 B.n543 B.n98 10.6151
R1021 B.n547 B.n98 10.6151
R1022 B.n548 B.n547 10.6151
R1023 B.n549 B.n548 10.6151
R1024 B.n549 B.n96 10.6151
R1025 B.n553 B.n96 10.6151
R1026 B.n554 B.n553 10.6151
R1027 B.n555 B.n554 10.6151
R1028 B.n555 B.n94 10.6151
R1029 B.n559 B.n94 10.6151
R1030 B.n560 B.n559 10.6151
R1031 B.n561 B.n560 10.6151
R1032 B.n561 B.n92 10.6151
R1033 B.n565 B.n92 10.6151
R1034 B.n566 B.n565 10.6151
R1035 B.n567 B.n566 10.6151
R1036 B.n265 B.n196 10.6151
R1037 B.n266 B.n265 10.6151
R1038 B.n267 B.n266 10.6151
R1039 B.n267 B.n194 10.6151
R1040 B.n271 B.n194 10.6151
R1041 B.n272 B.n271 10.6151
R1042 B.n273 B.n272 10.6151
R1043 B.n273 B.n192 10.6151
R1044 B.n277 B.n192 10.6151
R1045 B.n278 B.n277 10.6151
R1046 B.n279 B.n278 10.6151
R1047 B.n279 B.n190 10.6151
R1048 B.n283 B.n190 10.6151
R1049 B.n284 B.n283 10.6151
R1050 B.n285 B.n284 10.6151
R1051 B.n285 B.n188 10.6151
R1052 B.n289 B.n188 10.6151
R1053 B.n290 B.n289 10.6151
R1054 B.n291 B.n290 10.6151
R1055 B.n291 B.n186 10.6151
R1056 B.n295 B.n186 10.6151
R1057 B.n296 B.n295 10.6151
R1058 B.n297 B.n296 10.6151
R1059 B.n297 B.n184 10.6151
R1060 B.n301 B.n184 10.6151
R1061 B.n302 B.n301 10.6151
R1062 B.n303 B.n302 10.6151
R1063 B.n303 B.n182 10.6151
R1064 B.n307 B.n182 10.6151
R1065 B.n308 B.n307 10.6151
R1066 B.n309 B.n308 10.6151
R1067 B.n309 B.n180 10.6151
R1068 B.n313 B.n180 10.6151
R1069 B.n314 B.n313 10.6151
R1070 B.n315 B.n314 10.6151
R1071 B.n315 B.n178 10.6151
R1072 B.n319 B.n178 10.6151
R1073 B.n320 B.n319 10.6151
R1074 B.n321 B.n320 10.6151
R1075 B.n321 B.n176 10.6151
R1076 B.n325 B.n176 10.6151
R1077 B.n326 B.n325 10.6151
R1078 B.n327 B.n326 10.6151
R1079 B.n327 B.n174 10.6151
R1080 B.n331 B.n174 10.6151
R1081 B.n332 B.n331 10.6151
R1082 B.n333 B.n332 10.6151
R1083 B.n333 B.n172 10.6151
R1084 B.n337 B.n172 10.6151
R1085 B.n338 B.n337 10.6151
R1086 B.n339 B.n338 10.6151
R1087 B.n339 B.n170 10.6151
R1088 B.n343 B.n170 10.6151
R1089 B.n344 B.n343 10.6151
R1090 B.n345 B.n344 10.6151
R1091 B.n345 B.n168 10.6151
R1092 B.n349 B.n168 10.6151
R1093 B.n350 B.n349 10.6151
R1094 B.n351 B.n350 10.6151
R1095 B.n351 B.n166 10.6151
R1096 B.n355 B.n166 10.6151
R1097 B.n358 B.n357 10.6151
R1098 B.n358 B.n162 10.6151
R1099 B.n362 B.n162 10.6151
R1100 B.n363 B.n362 10.6151
R1101 B.n364 B.n363 10.6151
R1102 B.n364 B.n160 10.6151
R1103 B.n368 B.n160 10.6151
R1104 B.n369 B.n368 10.6151
R1105 B.n370 B.n369 10.6151
R1106 B.n374 B.n373 10.6151
R1107 B.n375 B.n374 10.6151
R1108 B.n375 B.n154 10.6151
R1109 B.n379 B.n154 10.6151
R1110 B.n380 B.n379 10.6151
R1111 B.n381 B.n380 10.6151
R1112 B.n381 B.n152 10.6151
R1113 B.n385 B.n152 10.6151
R1114 B.n386 B.n385 10.6151
R1115 B.n387 B.n386 10.6151
R1116 B.n387 B.n150 10.6151
R1117 B.n391 B.n150 10.6151
R1118 B.n392 B.n391 10.6151
R1119 B.n393 B.n392 10.6151
R1120 B.n393 B.n148 10.6151
R1121 B.n397 B.n148 10.6151
R1122 B.n398 B.n397 10.6151
R1123 B.n399 B.n398 10.6151
R1124 B.n399 B.n146 10.6151
R1125 B.n403 B.n146 10.6151
R1126 B.n404 B.n403 10.6151
R1127 B.n405 B.n404 10.6151
R1128 B.n405 B.n144 10.6151
R1129 B.n409 B.n144 10.6151
R1130 B.n410 B.n409 10.6151
R1131 B.n411 B.n410 10.6151
R1132 B.n411 B.n142 10.6151
R1133 B.n415 B.n142 10.6151
R1134 B.n416 B.n415 10.6151
R1135 B.n417 B.n416 10.6151
R1136 B.n417 B.n140 10.6151
R1137 B.n421 B.n140 10.6151
R1138 B.n422 B.n421 10.6151
R1139 B.n423 B.n422 10.6151
R1140 B.n423 B.n138 10.6151
R1141 B.n427 B.n138 10.6151
R1142 B.n428 B.n427 10.6151
R1143 B.n429 B.n428 10.6151
R1144 B.n429 B.n136 10.6151
R1145 B.n433 B.n136 10.6151
R1146 B.n434 B.n433 10.6151
R1147 B.n435 B.n434 10.6151
R1148 B.n435 B.n134 10.6151
R1149 B.n439 B.n134 10.6151
R1150 B.n440 B.n439 10.6151
R1151 B.n441 B.n440 10.6151
R1152 B.n441 B.n132 10.6151
R1153 B.n445 B.n132 10.6151
R1154 B.n446 B.n445 10.6151
R1155 B.n447 B.n446 10.6151
R1156 B.n447 B.n130 10.6151
R1157 B.n451 B.n130 10.6151
R1158 B.n452 B.n451 10.6151
R1159 B.n453 B.n452 10.6151
R1160 B.n453 B.n128 10.6151
R1161 B.n457 B.n128 10.6151
R1162 B.n458 B.n457 10.6151
R1163 B.n459 B.n458 10.6151
R1164 B.n459 B.n126 10.6151
R1165 B.n463 B.n126 10.6151
R1166 B.n464 B.n463 10.6151
R1167 B.n261 B.n260 10.6151
R1168 B.n260 B.n259 10.6151
R1169 B.n259 B.n198 10.6151
R1170 B.n255 B.n198 10.6151
R1171 B.n255 B.n254 10.6151
R1172 B.n254 B.n253 10.6151
R1173 B.n253 B.n200 10.6151
R1174 B.n249 B.n200 10.6151
R1175 B.n249 B.n248 10.6151
R1176 B.n248 B.n247 10.6151
R1177 B.n247 B.n202 10.6151
R1178 B.n243 B.n202 10.6151
R1179 B.n243 B.n242 10.6151
R1180 B.n242 B.n241 10.6151
R1181 B.n241 B.n204 10.6151
R1182 B.n237 B.n204 10.6151
R1183 B.n237 B.n236 10.6151
R1184 B.n236 B.n235 10.6151
R1185 B.n235 B.n206 10.6151
R1186 B.n231 B.n206 10.6151
R1187 B.n231 B.n230 10.6151
R1188 B.n230 B.n229 10.6151
R1189 B.n229 B.n208 10.6151
R1190 B.n225 B.n208 10.6151
R1191 B.n225 B.n224 10.6151
R1192 B.n224 B.n223 10.6151
R1193 B.n223 B.n210 10.6151
R1194 B.n219 B.n210 10.6151
R1195 B.n219 B.n218 10.6151
R1196 B.n218 B.n217 10.6151
R1197 B.n217 B.n212 10.6151
R1198 B.n213 B.n212 10.6151
R1199 B.n213 B.n0 10.6151
R1200 B.n819 B.n1 10.6151
R1201 B.n819 B.n818 10.6151
R1202 B.n818 B.n817 10.6151
R1203 B.n817 B.n4 10.6151
R1204 B.n813 B.n4 10.6151
R1205 B.n813 B.n812 10.6151
R1206 B.n812 B.n811 10.6151
R1207 B.n811 B.n6 10.6151
R1208 B.n807 B.n6 10.6151
R1209 B.n807 B.n806 10.6151
R1210 B.n806 B.n805 10.6151
R1211 B.n805 B.n8 10.6151
R1212 B.n801 B.n8 10.6151
R1213 B.n801 B.n800 10.6151
R1214 B.n800 B.n799 10.6151
R1215 B.n799 B.n10 10.6151
R1216 B.n795 B.n10 10.6151
R1217 B.n795 B.n794 10.6151
R1218 B.n794 B.n793 10.6151
R1219 B.n793 B.n12 10.6151
R1220 B.n789 B.n12 10.6151
R1221 B.n789 B.n788 10.6151
R1222 B.n788 B.n787 10.6151
R1223 B.n787 B.n14 10.6151
R1224 B.n783 B.n14 10.6151
R1225 B.n783 B.n782 10.6151
R1226 B.n782 B.n781 10.6151
R1227 B.n781 B.n16 10.6151
R1228 B.n777 B.n16 10.6151
R1229 B.n777 B.n776 10.6151
R1230 B.n776 B.n775 10.6151
R1231 B.n775 B.n18 10.6151
R1232 B.n771 B.n18 10.6151
R1233 B.n679 B.n52 9.36635
R1234 B.n662 B.n661 9.36635
R1235 B.n356 B.n355 9.36635
R1236 B.n373 B.n158 9.36635
R1237 B.n823 B.n0 2.81026
R1238 B.n823 B.n1 2.81026
R1239 B.n676 B.n52 1.24928
R1240 B.n663 B.n662 1.24928
R1241 B.n357 B.n356 1.24928
R1242 B.n370 B.n158 1.24928
R1243 VP.n6 VP.t1 272.935
R1244 VP.n17 VP.t0 241.766
R1245 VP.n24 VP.t5 241.766
R1246 VP.n31 VP.t3 241.766
R1247 VP.n14 VP.t2 241.766
R1248 VP.n7 VP.t4 241.766
R1249 VP.n9 VP.n8 161.3
R1250 VP.n10 VP.n5 161.3
R1251 VP.n12 VP.n11 161.3
R1252 VP.n13 VP.n4 161.3
R1253 VP.n30 VP.n0 161.3
R1254 VP.n29 VP.n28 161.3
R1255 VP.n27 VP.n1 161.3
R1256 VP.n26 VP.n25 161.3
R1257 VP.n23 VP.n2 161.3
R1258 VP.n22 VP.n21 161.3
R1259 VP.n20 VP.n3 161.3
R1260 VP.n19 VP.n18 161.3
R1261 VP.n17 VP.n16 87.7919
R1262 VP.n32 VP.n31 87.7919
R1263 VP.n15 VP.n14 87.7919
R1264 VP.n7 VP.n6 57.9788
R1265 VP.n22 VP.n3 54.1398
R1266 VP.n29 VP.n1 54.1398
R1267 VP.n12 VP.n5 54.1398
R1268 VP.n16 VP.n15 51.2118
R1269 VP.n18 VP.n3 27.0143
R1270 VP.n30 VP.n29 27.0143
R1271 VP.n13 VP.n12 27.0143
R1272 VP.n23 VP.n22 24.5923
R1273 VP.n25 VP.n1 24.5923
R1274 VP.n8 VP.n5 24.5923
R1275 VP.n18 VP.n17 23.1168
R1276 VP.n31 VP.n30 23.1168
R1277 VP.n14 VP.n13 23.1168
R1278 VP.n9 VP.n6 12.8269
R1279 VP.n24 VP.n23 12.2964
R1280 VP.n25 VP.n24 12.2964
R1281 VP.n8 VP.n7 12.2964
R1282 VP.n15 VP.n4 0.278335
R1283 VP.n19 VP.n16 0.278335
R1284 VP.n32 VP.n0 0.278335
R1285 VP.n10 VP.n9 0.189894
R1286 VP.n11 VP.n10 0.189894
R1287 VP.n11 VP.n4 0.189894
R1288 VP.n20 VP.n19 0.189894
R1289 VP.n21 VP.n20 0.189894
R1290 VP.n21 VP.n2 0.189894
R1291 VP.n26 VP.n2 0.189894
R1292 VP.n27 VP.n26 0.189894
R1293 VP.n28 VP.n27 0.189894
R1294 VP.n28 VP.n0 0.189894
R1295 VP VP.n32 0.153485
R1296 VTAIL.n426 VTAIL.n326 756.745
R1297 VTAIL.n102 VTAIL.n2 756.745
R1298 VTAIL.n320 VTAIL.n220 756.745
R1299 VTAIL.n212 VTAIL.n112 756.745
R1300 VTAIL.n361 VTAIL.n360 585
R1301 VTAIL.n358 VTAIL.n357 585
R1302 VTAIL.n367 VTAIL.n366 585
R1303 VTAIL.n369 VTAIL.n368 585
R1304 VTAIL.n354 VTAIL.n353 585
R1305 VTAIL.n375 VTAIL.n374 585
R1306 VTAIL.n377 VTAIL.n376 585
R1307 VTAIL.n350 VTAIL.n349 585
R1308 VTAIL.n383 VTAIL.n382 585
R1309 VTAIL.n385 VTAIL.n384 585
R1310 VTAIL.n346 VTAIL.n345 585
R1311 VTAIL.n391 VTAIL.n390 585
R1312 VTAIL.n393 VTAIL.n392 585
R1313 VTAIL.n342 VTAIL.n341 585
R1314 VTAIL.n399 VTAIL.n398 585
R1315 VTAIL.n402 VTAIL.n401 585
R1316 VTAIL.n400 VTAIL.n338 585
R1317 VTAIL.n407 VTAIL.n337 585
R1318 VTAIL.n409 VTAIL.n408 585
R1319 VTAIL.n411 VTAIL.n410 585
R1320 VTAIL.n334 VTAIL.n333 585
R1321 VTAIL.n417 VTAIL.n416 585
R1322 VTAIL.n419 VTAIL.n418 585
R1323 VTAIL.n330 VTAIL.n329 585
R1324 VTAIL.n425 VTAIL.n424 585
R1325 VTAIL.n427 VTAIL.n426 585
R1326 VTAIL.n37 VTAIL.n36 585
R1327 VTAIL.n34 VTAIL.n33 585
R1328 VTAIL.n43 VTAIL.n42 585
R1329 VTAIL.n45 VTAIL.n44 585
R1330 VTAIL.n30 VTAIL.n29 585
R1331 VTAIL.n51 VTAIL.n50 585
R1332 VTAIL.n53 VTAIL.n52 585
R1333 VTAIL.n26 VTAIL.n25 585
R1334 VTAIL.n59 VTAIL.n58 585
R1335 VTAIL.n61 VTAIL.n60 585
R1336 VTAIL.n22 VTAIL.n21 585
R1337 VTAIL.n67 VTAIL.n66 585
R1338 VTAIL.n69 VTAIL.n68 585
R1339 VTAIL.n18 VTAIL.n17 585
R1340 VTAIL.n75 VTAIL.n74 585
R1341 VTAIL.n78 VTAIL.n77 585
R1342 VTAIL.n76 VTAIL.n14 585
R1343 VTAIL.n83 VTAIL.n13 585
R1344 VTAIL.n85 VTAIL.n84 585
R1345 VTAIL.n87 VTAIL.n86 585
R1346 VTAIL.n10 VTAIL.n9 585
R1347 VTAIL.n93 VTAIL.n92 585
R1348 VTAIL.n95 VTAIL.n94 585
R1349 VTAIL.n6 VTAIL.n5 585
R1350 VTAIL.n101 VTAIL.n100 585
R1351 VTAIL.n103 VTAIL.n102 585
R1352 VTAIL.n321 VTAIL.n320 585
R1353 VTAIL.n319 VTAIL.n318 585
R1354 VTAIL.n224 VTAIL.n223 585
R1355 VTAIL.n313 VTAIL.n312 585
R1356 VTAIL.n311 VTAIL.n310 585
R1357 VTAIL.n228 VTAIL.n227 585
R1358 VTAIL.n305 VTAIL.n304 585
R1359 VTAIL.n303 VTAIL.n302 585
R1360 VTAIL.n301 VTAIL.n231 585
R1361 VTAIL.n235 VTAIL.n232 585
R1362 VTAIL.n296 VTAIL.n295 585
R1363 VTAIL.n294 VTAIL.n293 585
R1364 VTAIL.n237 VTAIL.n236 585
R1365 VTAIL.n288 VTAIL.n287 585
R1366 VTAIL.n286 VTAIL.n285 585
R1367 VTAIL.n241 VTAIL.n240 585
R1368 VTAIL.n280 VTAIL.n279 585
R1369 VTAIL.n278 VTAIL.n277 585
R1370 VTAIL.n245 VTAIL.n244 585
R1371 VTAIL.n272 VTAIL.n271 585
R1372 VTAIL.n270 VTAIL.n269 585
R1373 VTAIL.n249 VTAIL.n248 585
R1374 VTAIL.n264 VTAIL.n263 585
R1375 VTAIL.n262 VTAIL.n261 585
R1376 VTAIL.n253 VTAIL.n252 585
R1377 VTAIL.n256 VTAIL.n255 585
R1378 VTAIL.n213 VTAIL.n212 585
R1379 VTAIL.n211 VTAIL.n210 585
R1380 VTAIL.n116 VTAIL.n115 585
R1381 VTAIL.n205 VTAIL.n204 585
R1382 VTAIL.n203 VTAIL.n202 585
R1383 VTAIL.n120 VTAIL.n119 585
R1384 VTAIL.n197 VTAIL.n196 585
R1385 VTAIL.n195 VTAIL.n194 585
R1386 VTAIL.n193 VTAIL.n123 585
R1387 VTAIL.n127 VTAIL.n124 585
R1388 VTAIL.n188 VTAIL.n187 585
R1389 VTAIL.n186 VTAIL.n185 585
R1390 VTAIL.n129 VTAIL.n128 585
R1391 VTAIL.n180 VTAIL.n179 585
R1392 VTAIL.n178 VTAIL.n177 585
R1393 VTAIL.n133 VTAIL.n132 585
R1394 VTAIL.n172 VTAIL.n171 585
R1395 VTAIL.n170 VTAIL.n169 585
R1396 VTAIL.n137 VTAIL.n136 585
R1397 VTAIL.n164 VTAIL.n163 585
R1398 VTAIL.n162 VTAIL.n161 585
R1399 VTAIL.n141 VTAIL.n140 585
R1400 VTAIL.n156 VTAIL.n155 585
R1401 VTAIL.n154 VTAIL.n153 585
R1402 VTAIL.n145 VTAIL.n144 585
R1403 VTAIL.n148 VTAIL.n147 585
R1404 VTAIL.t4 VTAIL.n254 327.466
R1405 VTAIL.t11 VTAIL.n146 327.466
R1406 VTAIL.t0 VTAIL.n359 327.466
R1407 VTAIL.t9 VTAIL.n35 327.466
R1408 VTAIL.n360 VTAIL.n357 171.744
R1409 VTAIL.n367 VTAIL.n357 171.744
R1410 VTAIL.n368 VTAIL.n367 171.744
R1411 VTAIL.n368 VTAIL.n353 171.744
R1412 VTAIL.n375 VTAIL.n353 171.744
R1413 VTAIL.n376 VTAIL.n375 171.744
R1414 VTAIL.n376 VTAIL.n349 171.744
R1415 VTAIL.n383 VTAIL.n349 171.744
R1416 VTAIL.n384 VTAIL.n383 171.744
R1417 VTAIL.n384 VTAIL.n345 171.744
R1418 VTAIL.n391 VTAIL.n345 171.744
R1419 VTAIL.n392 VTAIL.n391 171.744
R1420 VTAIL.n392 VTAIL.n341 171.744
R1421 VTAIL.n399 VTAIL.n341 171.744
R1422 VTAIL.n401 VTAIL.n399 171.744
R1423 VTAIL.n401 VTAIL.n400 171.744
R1424 VTAIL.n400 VTAIL.n337 171.744
R1425 VTAIL.n409 VTAIL.n337 171.744
R1426 VTAIL.n410 VTAIL.n409 171.744
R1427 VTAIL.n410 VTAIL.n333 171.744
R1428 VTAIL.n417 VTAIL.n333 171.744
R1429 VTAIL.n418 VTAIL.n417 171.744
R1430 VTAIL.n418 VTAIL.n329 171.744
R1431 VTAIL.n425 VTAIL.n329 171.744
R1432 VTAIL.n426 VTAIL.n425 171.744
R1433 VTAIL.n36 VTAIL.n33 171.744
R1434 VTAIL.n43 VTAIL.n33 171.744
R1435 VTAIL.n44 VTAIL.n43 171.744
R1436 VTAIL.n44 VTAIL.n29 171.744
R1437 VTAIL.n51 VTAIL.n29 171.744
R1438 VTAIL.n52 VTAIL.n51 171.744
R1439 VTAIL.n52 VTAIL.n25 171.744
R1440 VTAIL.n59 VTAIL.n25 171.744
R1441 VTAIL.n60 VTAIL.n59 171.744
R1442 VTAIL.n60 VTAIL.n21 171.744
R1443 VTAIL.n67 VTAIL.n21 171.744
R1444 VTAIL.n68 VTAIL.n67 171.744
R1445 VTAIL.n68 VTAIL.n17 171.744
R1446 VTAIL.n75 VTAIL.n17 171.744
R1447 VTAIL.n77 VTAIL.n75 171.744
R1448 VTAIL.n77 VTAIL.n76 171.744
R1449 VTAIL.n76 VTAIL.n13 171.744
R1450 VTAIL.n85 VTAIL.n13 171.744
R1451 VTAIL.n86 VTAIL.n85 171.744
R1452 VTAIL.n86 VTAIL.n9 171.744
R1453 VTAIL.n93 VTAIL.n9 171.744
R1454 VTAIL.n94 VTAIL.n93 171.744
R1455 VTAIL.n94 VTAIL.n5 171.744
R1456 VTAIL.n101 VTAIL.n5 171.744
R1457 VTAIL.n102 VTAIL.n101 171.744
R1458 VTAIL.n320 VTAIL.n319 171.744
R1459 VTAIL.n319 VTAIL.n223 171.744
R1460 VTAIL.n312 VTAIL.n223 171.744
R1461 VTAIL.n312 VTAIL.n311 171.744
R1462 VTAIL.n311 VTAIL.n227 171.744
R1463 VTAIL.n304 VTAIL.n227 171.744
R1464 VTAIL.n304 VTAIL.n303 171.744
R1465 VTAIL.n303 VTAIL.n231 171.744
R1466 VTAIL.n235 VTAIL.n231 171.744
R1467 VTAIL.n295 VTAIL.n235 171.744
R1468 VTAIL.n295 VTAIL.n294 171.744
R1469 VTAIL.n294 VTAIL.n236 171.744
R1470 VTAIL.n287 VTAIL.n236 171.744
R1471 VTAIL.n287 VTAIL.n286 171.744
R1472 VTAIL.n286 VTAIL.n240 171.744
R1473 VTAIL.n279 VTAIL.n240 171.744
R1474 VTAIL.n279 VTAIL.n278 171.744
R1475 VTAIL.n278 VTAIL.n244 171.744
R1476 VTAIL.n271 VTAIL.n244 171.744
R1477 VTAIL.n271 VTAIL.n270 171.744
R1478 VTAIL.n270 VTAIL.n248 171.744
R1479 VTAIL.n263 VTAIL.n248 171.744
R1480 VTAIL.n263 VTAIL.n262 171.744
R1481 VTAIL.n262 VTAIL.n252 171.744
R1482 VTAIL.n255 VTAIL.n252 171.744
R1483 VTAIL.n212 VTAIL.n211 171.744
R1484 VTAIL.n211 VTAIL.n115 171.744
R1485 VTAIL.n204 VTAIL.n115 171.744
R1486 VTAIL.n204 VTAIL.n203 171.744
R1487 VTAIL.n203 VTAIL.n119 171.744
R1488 VTAIL.n196 VTAIL.n119 171.744
R1489 VTAIL.n196 VTAIL.n195 171.744
R1490 VTAIL.n195 VTAIL.n123 171.744
R1491 VTAIL.n127 VTAIL.n123 171.744
R1492 VTAIL.n187 VTAIL.n127 171.744
R1493 VTAIL.n187 VTAIL.n186 171.744
R1494 VTAIL.n186 VTAIL.n128 171.744
R1495 VTAIL.n179 VTAIL.n128 171.744
R1496 VTAIL.n179 VTAIL.n178 171.744
R1497 VTAIL.n178 VTAIL.n132 171.744
R1498 VTAIL.n171 VTAIL.n132 171.744
R1499 VTAIL.n171 VTAIL.n170 171.744
R1500 VTAIL.n170 VTAIL.n136 171.744
R1501 VTAIL.n163 VTAIL.n136 171.744
R1502 VTAIL.n163 VTAIL.n162 171.744
R1503 VTAIL.n162 VTAIL.n140 171.744
R1504 VTAIL.n155 VTAIL.n140 171.744
R1505 VTAIL.n155 VTAIL.n154 171.744
R1506 VTAIL.n154 VTAIL.n144 171.744
R1507 VTAIL.n147 VTAIL.n144 171.744
R1508 VTAIL.n360 VTAIL.t0 85.8723
R1509 VTAIL.n36 VTAIL.t9 85.8723
R1510 VTAIL.n255 VTAIL.t4 85.8723
R1511 VTAIL.n147 VTAIL.t11 85.8723
R1512 VTAIL.n1 VTAIL.n0 51.7061
R1513 VTAIL.n109 VTAIL.n108 51.7061
R1514 VTAIL.n219 VTAIL.n218 51.7061
R1515 VTAIL.n111 VTAIL.n110 51.7061
R1516 VTAIL.n111 VTAIL.n109 32.5393
R1517 VTAIL.n431 VTAIL.n430 32.1853
R1518 VTAIL.n107 VTAIL.n106 32.1853
R1519 VTAIL.n325 VTAIL.n324 32.1853
R1520 VTAIL.n217 VTAIL.n216 32.1853
R1521 VTAIL.n431 VTAIL.n325 30.6255
R1522 VTAIL.n361 VTAIL.n359 16.3895
R1523 VTAIL.n37 VTAIL.n35 16.3895
R1524 VTAIL.n256 VTAIL.n254 16.3895
R1525 VTAIL.n148 VTAIL.n146 16.3895
R1526 VTAIL.n408 VTAIL.n407 13.1884
R1527 VTAIL.n84 VTAIL.n83 13.1884
R1528 VTAIL.n302 VTAIL.n301 13.1884
R1529 VTAIL.n194 VTAIL.n193 13.1884
R1530 VTAIL.n362 VTAIL.n358 12.8005
R1531 VTAIL.n406 VTAIL.n338 12.8005
R1532 VTAIL.n411 VTAIL.n336 12.8005
R1533 VTAIL.n38 VTAIL.n34 12.8005
R1534 VTAIL.n82 VTAIL.n14 12.8005
R1535 VTAIL.n87 VTAIL.n12 12.8005
R1536 VTAIL.n305 VTAIL.n230 12.8005
R1537 VTAIL.n300 VTAIL.n232 12.8005
R1538 VTAIL.n257 VTAIL.n253 12.8005
R1539 VTAIL.n197 VTAIL.n122 12.8005
R1540 VTAIL.n192 VTAIL.n124 12.8005
R1541 VTAIL.n149 VTAIL.n145 12.8005
R1542 VTAIL.n366 VTAIL.n365 12.0247
R1543 VTAIL.n403 VTAIL.n402 12.0247
R1544 VTAIL.n412 VTAIL.n334 12.0247
R1545 VTAIL.n42 VTAIL.n41 12.0247
R1546 VTAIL.n79 VTAIL.n78 12.0247
R1547 VTAIL.n88 VTAIL.n10 12.0247
R1548 VTAIL.n306 VTAIL.n228 12.0247
R1549 VTAIL.n297 VTAIL.n296 12.0247
R1550 VTAIL.n261 VTAIL.n260 12.0247
R1551 VTAIL.n198 VTAIL.n120 12.0247
R1552 VTAIL.n189 VTAIL.n188 12.0247
R1553 VTAIL.n153 VTAIL.n152 12.0247
R1554 VTAIL.n369 VTAIL.n356 11.249
R1555 VTAIL.n398 VTAIL.n340 11.249
R1556 VTAIL.n416 VTAIL.n415 11.249
R1557 VTAIL.n45 VTAIL.n32 11.249
R1558 VTAIL.n74 VTAIL.n16 11.249
R1559 VTAIL.n92 VTAIL.n91 11.249
R1560 VTAIL.n310 VTAIL.n309 11.249
R1561 VTAIL.n293 VTAIL.n234 11.249
R1562 VTAIL.n264 VTAIL.n251 11.249
R1563 VTAIL.n202 VTAIL.n201 11.249
R1564 VTAIL.n185 VTAIL.n126 11.249
R1565 VTAIL.n156 VTAIL.n143 11.249
R1566 VTAIL.n370 VTAIL.n354 10.4732
R1567 VTAIL.n397 VTAIL.n342 10.4732
R1568 VTAIL.n419 VTAIL.n332 10.4732
R1569 VTAIL.n46 VTAIL.n30 10.4732
R1570 VTAIL.n73 VTAIL.n18 10.4732
R1571 VTAIL.n95 VTAIL.n8 10.4732
R1572 VTAIL.n313 VTAIL.n226 10.4732
R1573 VTAIL.n292 VTAIL.n237 10.4732
R1574 VTAIL.n265 VTAIL.n249 10.4732
R1575 VTAIL.n205 VTAIL.n118 10.4732
R1576 VTAIL.n184 VTAIL.n129 10.4732
R1577 VTAIL.n157 VTAIL.n141 10.4732
R1578 VTAIL.n374 VTAIL.n373 9.69747
R1579 VTAIL.n394 VTAIL.n393 9.69747
R1580 VTAIL.n420 VTAIL.n330 9.69747
R1581 VTAIL.n50 VTAIL.n49 9.69747
R1582 VTAIL.n70 VTAIL.n69 9.69747
R1583 VTAIL.n96 VTAIL.n6 9.69747
R1584 VTAIL.n314 VTAIL.n224 9.69747
R1585 VTAIL.n289 VTAIL.n288 9.69747
R1586 VTAIL.n269 VTAIL.n268 9.69747
R1587 VTAIL.n206 VTAIL.n116 9.69747
R1588 VTAIL.n181 VTAIL.n180 9.69747
R1589 VTAIL.n161 VTAIL.n160 9.69747
R1590 VTAIL.n430 VTAIL.n429 9.45567
R1591 VTAIL.n106 VTAIL.n105 9.45567
R1592 VTAIL.n324 VTAIL.n323 9.45567
R1593 VTAIL.n216 VTAIL.n215 9.45567
R1594 VTAIL.n328 VTAIL.n327 9.3005
R1595 VTAIL.n423 VTAIL.n422 9.3005
R1596 VTAIL.n421 VTAIL.n420 9.3005
R1597 VTAIL.n332 VTAIL.n331 9.3005
R1598 VTAIL.n415 VTAIL.n414 9.3005
R1599 VTAIL.n413 VTAIL.n412 9.3005
R1600 VTAIL.n336 VTAIL.n335 9.3005
R1601 VTAIL.n381 VTAIL.n380 9.3005
R1602 VTAIL.n379 VTAIL.n378 9.3005
R1603 VTAIL.n352 VTAIL.n351 9.3005
R1604 VTAIL.n373 VTAIL.n372 9.3005
R1605 VTAIL.n371 VTAIL.n370 9.3005
R1606 VTAIL.n356 VTAIL.n355 9.3005
R1607 VTAIL.n365 VTAIL.n364 9.3005
R1608 VTAIL.n363 VTAIL.n362 9.3005
R1609 VTAIL.n348 VTAIL.n347 9.3005
R1610 VTAIL.n387 VTAIL.n386 9.3005
R1611 VTAIL.n389 VTAIL.n388 9.3005
R1612 VTAIL.n344 VTAIL.n343 9.3005
R1613 VTAIL.n395 VTAIL.n394 9.3005
R1614 VTAIL.n397 VTAIL.n396 9.3005
R1615 VTAIL.n340 VTAIL.n339 9.3005
R1616 VTAIL.n404 VTAIL.n403 9.3005
R1617 VTAIL.n406 VTAIL.n405 9.3005
R1618 VTAIL.n429 VTAIL.n428 9.3005
R1619 VTAIL.n4 VTAIL.n3 9.3005
R1620 VTAIL.n99 VTAIL.n98 9.3005
R1621 VTAIL.n97 VTAIL.n96 9.3005
R1622 VTAIL.n8 VTAIL.n7 9.3005
R1623 VTAIL.n91 VTAIL.n90 9.3005
R1624 VTAIL.n89 VTAIL.n88 9.3005
R1625 VTAIL.n12 VTAIL.n11 9.3005
R1626 VTAIL.n57 VTAIL.n56 9.3005
R1627 VTAIL.n55 VTAIL.n54 9.3005
R1628 VTAIL.n28 VTAIL.n27 9.3005
R1629 VTAIL.n49 VTAIL.n48 9.3005
R1630 VTAIL.n47 VTAIL.n46 9.3005
R1631 VTAIL.n32 VTAIL.n31 9.3005
R1632 VTAIL.n41 VTAIL.n40 9.3005
R1633 VTAIL.n39 VTAIL.n38 9.3005
R1634 VTAIL.n24 VTAIL.n23 9.3005
R1635 VTAIL.n63 VTAIL.n62 9.3005
R1636 VTAIL.n65 VTAIL.n64 9.3005
R1637 VTAIL.n20 VTAIL.n19 9.3005
R1638 VTAIL.n71 VTAIL.n70 9.3005
R1639 VTAIL.n73 VTAIL.n72 9.3005
R1640 VTAIL.n16 VTAIL.n15 9.3005
R1641 VTAIL.n80 VTAIL.n79 9.3005
R1642 VTAIL.n82 VTAIL.n81 9.3005
R1643 VTAIL.n105 VTAIL.n104 9.3005
R1644 VTAIL.n282 VTAIL.n281 9.3005
R1645 VTAIL.n284 VTAIL.n283 9.3005
R1646 VTAIL.n239 VTAIL.n238 9.3005
R1647 VTAIL.n290 VTAIL.n289 9.3005
R1648 VTAIL.n292 VTAIL.n291 9.3005
R1649 VTAIL.n234 VTAIL.n233 9.3005
R1650 VTAIL.n298 VTAIL.n297 9.3005
R1651 VTAIL.n300 VTAIL.n299 9.3005
R1652 VTAIL.n323 VTAIL.n322 9.3005
R1653 VTAIL.n222 VTAIL.n221 9.3005
R1654 VTAIL.n317 VTAIL.n316 9.3005
R1655 VTAIL.n315 VTAIL.n314 9.3005
R1656 VTAIL.n226 VTAIL.n225 9.3005
R1657 VTAIL.n309 VTAIL.n308 9.3005
R1658 VTAIL.n307 VTAIL.n306 9.3005
R1659 VTAIL.n230 VTAIL.n229 9.3005
R1660 VTAIL.n243 VTAIL.n242 9.3005
R1661 VTAIL.n276 VTAIL.n275 9.3005
R1662 VTAIL.n274 VTAIL.n273 9.3005
R1663 VTAIL.n247 VTAIL.n246 9.3005
R1664 VTAIL.n268 VTAIL.n267 9.3005
R1665 VTAIL.n266 VTAIL.n265 9.3005
R1666 VTAIL.n251 VTAIL.n250 9.3005
R1667 VTAIL.n260 VTAIL.n259 9.3005
R1668 VTAIL.n258 VTAIL.n257 9.3005
R1669 VTAIL.n174 VTAIL.n173 9.3005
R1670 VTAIL.n176 VTAIL.n175 9.3005
R1671 VTAIL.n131 VTAIL.n130 9.3005
R1672 VTAIL.n182 VTAIL.n181 9.3005
R1673 VTAIL.n184 VTAIL.n183 9.3005
R1674 VTAIL.n126 VTAIL.n125 9.3005
R1675 VTAIL.n190 VTAIL.n189 9.3005
R1676 VTAIL.n192 VTAIL.n191 9.3005
R1677 VTAIL.n215 VTAIL.n214 9.3005
R1678 VTAIL.n114 VTAIL.n113 9.3005
R1679 VTAIL.n209 VTAIL.n208 9.3005
R1680 VTAIL.n207 VTAIL.n206 9.3005
R1681 VTAIL.n118 VTAIL.n117 9.3005
R1682 VTAIL.n201 VTAIL.n200 9.3005
R1683 VTAIL.n199 VTAIL.n198 9.3005
R1684 VTAIL.n122 VTAIL.n121 9.3005
R1685 VTAIL.n135 VTAIL.n134 9.3005
R1686 VTAIL.n168 VTAIL.n167 9.3005
R1687 VTAIL.n166 VTAIL.n165 9.3005
R1688 VTAIL.n139 VTAIL.n138 9.3005
R1689 VTAIL.n160 VTAIL.n159 9.3005
R1690 VTAIL.n158 VTAIL.n157 9.3005
R1691 VTAIL.n143 VTAIL.n142 9.3005
R1692 VTAIL.n152 VTAIL.n151 9.3005
R1693 VTAIL.n150 VTAIL.n149 9.3005
R1694 VTAIL.n377 VTAIL.n352 8.92171
R1695 VTAIL.n390 VTAIL.n344 8.92171
R1696 VTAIL.n424 VTAIL.n423 8.92171
R1697 VTAIL.n53 VTAIL.n28 8.92171
R1698 VTAIL.n66 VTAIL.n20 8.92171
R1699 VTAIL.n100 VTAIL.n99 8.92171
R1700 VTAIL.n318 VTAIL.n317 8.92171
R1701 VTAIL.n285 VTAIL.n239 8.92171
R1702 VTAIL.n272 VTAIL.n247 8.92171
R1703 VTAIL.n210 VTAIL.n209 8.92171
R1704 VTAIL.n177 VTAIL.n131 8.92171
R1705 VTAIL.n164 VTAIL.n139 8.92171
R1706 VTAIL.n378 VTAIL.n350 8.14595
R1707 VTAIL.n389 VTAIL.n346 8.14595
R1708 VTAIL.n427 VTAIL.n328 8.14595
R1709 VTAIL.n54 VTAIL.n26 8.14595
R1710 VTAIL.n65 VTAIL.n22 8.14595
R1711 VTAIL.n103 VTAIL.n4 8.14595
R1712 VTAIL.n321 VTAIL.n222 8.14595
R1713 VTAIL.n284 VTAIL.n241 8.14595
R1714 VTAIL.n273 VTAIL.n245 8.14595
R1715 VTAIL.n213 VTAIL.n114 8.14595
R1716 VTAIL.n176 VTAIL.n133 8.14595
R1717 VTAIL.n165 VTAIL.n137 8.14595
R1718 VTAIL.n382 VTAIL.n381 7.3702
R1719 VTAIL.n386 VTAIL.n385 7.3702
R1720 VTAIL.n428 VTAIL.n326 7.3702
R1721 VTAIL.n58 VTAIL.n57 7.3702
R1722 VTAIL.n62 VTAIL.n61 7.3702
R1723 VTAIL.n104 VTAIL.n2 7.3702
R1724 VTAIL.n322 VTAIL.n220 7.3702
R1725 VTAIL.n281 VTAIL.n280 7.3702
R1726 VTAIL.n277 VTAIL.n276 7.3702
R1727 VTAIL.n214 VTAIL.n112 7.3702
R1728 VTAIL.n173 VTAIL.n172 7.3702
R1729 VTAIL.n169 VTAIL.n168 7.3702
R1730 VTAIL.n382 VTAIL.n348 6.59444
R1731 VTAIL.n385 VTAIL.n348 6.59444
R1732 VTAIL.n430 VTAIL.n326 6.59444
R1733 VTAIL.n58 VTAIL.n24 6.59444
R1734 VTAIL.n61 VTAIL.n24 6.59444
R1735 VTAIL.n106 VTAIL.n2 6.59444
R1736 VTAIL.n324 VTAIL.n220 6.59444
R1737 VTAIL.n280 VTAIL.n243 6.59444
R1738 VTAIL.n277 VTAIL.n243 6.59444
R1739 VTAIL.n216 VTAIL.n112 6.59444
R1740 VTAIL.n172 VTAIL.n135 6.59444
R1741 VTAIL.n169 VTAIL.n135 6.59444
R1742 VTAIL.n381 VTAIL.n350 5.81868
R1743 VTAIL.n386 VTAIL.n346 5.81868
R1744 VTAIL.n428 VTAIL.n427 5.81868
R1745 VTAIL.n57 VTAIL.n26 5.81868
R1746 VTAIL.n62 VTAIL.n22 5.81868
R1747 VTAIL.n104 VTAIL.n103 5.81868
R1748 VTAIL.n322 VTAIL.n321 5.81868
R1749 VTAIL.n281 VTAIL.n241 5.81868
R1750 VTAIL.n276 VTAIL.n245 5.81868
R1751 VTAIL.n214 VTAIL.n213 5.81868
R1752 VTAIL.n173 VTAIL.n133 5.81868
R1753 VTAIL.n168 VTAIL.n137 5.81868
R1754 VTAIL.n378 VTAIL.n377 5.04292
R1755 VTAIL.n390 VTAIL.n389 5.04292
R1756 VTAIL.n424 VTAIL.n328 5.04292
R1757 VTAIL.n54 VTAIL.n53 5.04292
R1758 VTAIL.n66 VTAIL.n65 5.04292
R1759 VTAIL.n100 VTAIL.n4 5.04292
R1760 VTAIL.n318 VTAIL.n222 5.04292
R1761 VTAIL.n285 VTAIL.n284 5.04292
R1762 VTAIL.n273 VTAIL.n272 5.04292
R1763 VTAIL.n210 VTAIL.n114 5.04292
R1764 VTAIL.n177 VTAIL.n176 5.04292
R1765 VTAIL.n165 VTAIL.n164 5.04292
R1766 VTAIL.n374 VTAIL.n352 4.26717
R1767 VTAIL.n393 VTAIL.n344 4.26717
R1768 VTAIL.n423 VTAIL.n330 4.26717
R1769 VTAIL.n50 VTAIL.n28 4.26717
R1770 VTAIL.n69 VTAIL.n20 4.26717
R1771 VTAIL.n99 VTAIL.n6 4.26717
R1772 VTAIL.n317 VTAIL.n224 4.26717
R1773 VTAIL.n288 VTAIL.n239 4.26717
R1774 VTAIL.n269 VTAIL.n247 4.26717
R1775 VTAIL.n209 VTAIL.n116 4.26717
R1776 VTAIL.n180 VTAIL.n131 4.26717
R1777 VTAIL.n161 VTAIL.n139 4.26717
R1778 VTAIL.n363 VTAIL.n359 3.70982
R1779 VTAIL.n39 VTAIL.n35 3.70982
R1780 VTAIL.n258 VTAIL.n254 3.70982
R1781 VTAIL.n150 VTAIL.n146 3.70982
R1782 VTAIL.n373 VTAIL.n354 3.49141
R1783 VTAIL.n394 VTAIL.n342 3.49141
R1784 VTAIL.n420 VTAIL.n419 3.49141
R1785 VTAIL.n49 VTAIL.n30 3.49141
R1786 VTAIL.n70 VTAIL.n18 3.49141
R1787 VTAIL.n96 VTAIL.n95 3.49141
R1788 VTAIL.n314 VTAIL.n313 3.49141
R1789 VTAIL.n289 VTAIL.n237 3.49141
R1790 VTAIL.n268 VTAIL.n249 3.49141
R1791 VTAIL.n206 VTAIL.n205 3.49141
R1792 VTAIL.n181 VTAIL.n129 3.49141
R1793 VTAIL.n160 VTAIL.n141 3.49141
R1794 VTAIL.n370 VTAIL.n369 2.71565
R1795 VTAIL.n398 VTAIL.n397 2.71565
R1796 VTAIL.n416 VTAIL.n332 2.71565
R1797 VTAIL.n46 VTAIL.n45 2.71565
R1798 VTAIL.n74 VTAIL.n73 2.71565
R1799 VTAIL.n92 VTAIL.n8 2.71565
R1800 VTAIL.n310 VTAIL.n226 2.71565
R1801 VTAIL.n293 VTAIL.n292 2.71565
R1802 VTAIL.n265 VTAIL.n264 2.71565
R1803 VTAIL.n202 VTAIL.n118 2.71565
R1804 VTAIL.n185 VTAIL.n184 2.71565
R1805 VTAIL.n157 VTAIL.n156 2.71565
R1806 VTAIL.n366 VTAIL.n356 1.93989
R1807 VTAIL.n402 VTAIL.n340 1.93989
R1808 VTAIL.n415 VTAIL.n334 1.93989
R1809 VTAIL.n42 VTAIL.n32 1.93989
R1810 VTAIL.n78 VTAIL.n16 1.93989
R1811 VTAIL.n91 VTAIL.n10 1.93989
R1812 VTAIL.n309 VTAIL.n228 1.93989
R1813 VTAIL.n296 VTAIL.n234 1.93989
R1814 VTAIL.n261 VTAIL.n251 1.93989
R1815 VTAIL.n201 VTAIL.n120 1.93989
R1816 VTAIL.n188 VTAIL.n126 1.93989
R1817 VTAIL.n153 VTAIL.n143 1.93989
R1818 VTAIL.n217 VTAIL.n111 1.91429
R1819 VTAIL.n325 VTAIL.n219 1.91429
R1820 VTAIL.n109 VTAIL.n107 1.91429
R1821 VTAIL.n0 VTAIL.t1 1.7149
R1822 VTAIL.n0 VTAIL.t10 1.7149
R1823 VTAIL.n108 VTAIL.t8 1.7149
R1824 VTAIL.n108 VTAIL.t6 1.7149
R1825 VTAIL.n218 VTAIL.t5 1.7149
R1826 VTAIL.n218 VTAIL.t7 1.7149
R1827 VTAIL.n110 VTAIL.t2 1.7149
R1828 VTAIL.n110 VTAIL.t3 1.7149
R1829 VTAIL.n219 VTAIL.n217 1.42722
R1830 VTAIL.n107 VTAIL.n1 1.42722
R1831 VTAIL VTAIL.n431 1.37766
R1832 VTAIL.n365 VTAIL.n358 1.16414
R1833 VTAIL.n403 VTAIL.n338 1.16414
R1834 VTAIL.n412 VTAIL.n411 1.16414
R1835 VTAIL.n41 VTAIL.n34 1.16414
R1836 VTAIL.n79 VTAIL.n14 1.16414
R1837 VTAIL.n88 VTAIL.n87 1.16414
R1838 VTAIL.n306 VTAIL.n305 1.16414
R1839 VTAIL.n297 VTAIL.n232 1.16414
R1840 VTAIL.n260 VTAIL.n253 1.16414
R1841 VTAIL.n198 VTAIL.n197 1.16414
R1842 VTAIL.n189 VTAIL.n124 1.16414
R1843 VTAIL.n152 VTAIL.n145 1.16414
R1844 VTAIL VTAIL.n1 0.537138
R1845 VTAIL.n362 VTAIL.n361 0.388379
R1846 VTAIL.n407 VTAIL.n406 0.388379
R1847 VTAIL.n408 VTAIL.n336 0.388379
R1848 VTAIL.n38 VTAIL.n37 0.388379
R1849 VTAIL.n83 VTAIL.n82 0.388379
R1850 VTAIL.n84 VTAIL.n12 0.388379
R1851 VTAIL.n302 VTAIL.n230 0.388379
R1852 VTAIL.n301 VTAIL.n300 0.388379
R1853 VTAIL.n257 VTAIL.n256 0.388379
R1854 VTAIL.n194 VTAIL.n122 0.388379
R1855 VTAIL.n193 VTAIL.n192 0.388379
R1856 VTAIL.n149 VTAIL.n148 0.388379
R1857 VTAIL.n364 VTAIL.n363 0.155672
R1858 VTAIL.n364 VTAIL.n355 0.155672
R1859 VTAIL.n371 VTAIL.n355 0.155672
R1860 VTAIL.n372 VTAIL.n371 0.155672
R1861 VTAIL.n372 VTAIL.n351 0.155672
R1862 VTAIL.n379 VTAIL.n351 0.155672
R1863 VTAIL.n380 VTAIL.n379 0.155672
R1864 VTAIL.n380 VTAIL.n347 0.155672
R1865 VTAIL.n387 VTAIL.n347 0.155672
R1866 VTAIL.n388 VTAIL.n387 0.155672
R1867 VTAIL.n388 VTAIL.n343 0.155672
R1868 VTAIL.n395 VTAIL.n343 0.155672
R1869 VTAIL.n396 VTAIL.n395 0.155672
R1870 VTAIL.n396 VTAIL.n339 0.155672
R1871 VTAIL.n404 VTAIL.n339 0.155672
R1872 VTAIL.n405 VTAIL.n404 0.155672
R1873 VTAIL.n405 VTAIL.n335 0.155672
R1874 VTAIL.n413 VTAIL.n335 0.155672
R1875 VTAIL.n414 VTAIL.n413 0.155672
R1876 VTAIL.n414 VTAIL.n331 0.155672
R1877 VTAIL.n421 VTAIL.n331 0.155672
R1878 VTAIL.n422 VTAIL.n421 0.155672
R1879 VTAIL.n422 VTAIL.n327 0.155672
R1880 VTAIL.n429 VTAIL.n327 0.155672
R1881 VTAIL.n40 VTAIL.n39 0.155672
R1882 VTAIL.n40 VTAIL.n31 0.155672
R1883 VTAIL.n47 VTAIL.n31 0.155672
R1884 VTAIL.n48 VTAIL.n47 0.155672
R1885 VTAIL.n48 VTAIL.n27 0.155672
R1886 VTAIL.n55 VTAIL.n27 0.155672
R1887 VTAIL.n56 VTAIL.n55 0.155672
R1888 VTAIL.n56 VTAIL.n23 0.155672
R1889 VTAIL.n63 VTAIL.n23 0.155672
R1890 VTAIL.n64 VTAIL.n63 0.155672
R1891 VTAIL.n64 VTAIL.n19 0.155672
R1892 VTAIL.n71 VTAIL.n19 0.155672
R1893 VTAIL.n72 VTAIL.n71 0.155672
R1894 VTAIL.n72 VTAIL.n15 0.155672
R1895 VTAIL.n80 VTAIL.n15 0.155672
R1896 VTAIL.n81 VTAIL.n80 0.155672
R1897 VTAIL.n81 VTAIL.n11 0.155672
R1898 VTAIL.n89 VTAIL.n11 0.155672
R1899 VTAIL.n90 VTAIL.n89 0.155672
R1900 VTAIL.n90 VTAIL.n7 0.155672
R1901 VTAIL.n97 VTAIL.n7 0.155672
R1902 VTAIL.n98 VTAIL.n97 0.155672
R1903 VTAIL.n98 VTAIL.n3 0.155672
R1904 VTAIL.n105 VTAIL.n3 0.155672
R1905 VTAIL.n323 VTAIL.n221 0.155672
R1906 VTAIL.n316 VTAIL.n221 0.155672
R1907 VTAIL.n316 VTAIL.n315 0.155672
R1908 VTAIL.n315 VTAIL.n225 0.155672
R1909 VTAIL.n308 VTAIL.n225 0.155672
R1910 VTAIL.n308 VTAIL.n307 0.155672
R1911 VTAIL.n307 VTAIL.n229 0.155672
R1912 VTAIL.n299 VTAIL.n229 0.155672
R1913 VTAIL.n299 VTAIL.n298 0.155672
R1914 VTAIL.n298 VTAIL.n233 0.155672
R1915 VTAIL.n291 VTAIL.n233 0.155672
R1916 VTAIL.n291 VTAIL.n290 0.155672
R1917 VTAIL.n290 VTAIL.n238 0.155672
R1918 VTAIL.n283 VTAIL.n238 0.155672
R1919 VTAIL.n283 VTAIL.n282 0.155672
R1920 VTAIL.n282 VTAIL.n242 0.155672
R1921 VTAIL.n275 VTAIL.n242 0.155672
R1922 VTAIL.n275 VTAIL.n274 0.155672
R1923 VTAIL.n274 VTAIL.n246 0.155672
R1924 VTAIL.n267 VTAIL.n246 0.155672
R1925 VTAIL.n267 VTAIL.n266 0.155672
R1926 VTAIL.n266 VTAIL.n250 0.155672
R1927 VTAIL.n259 VTAIL.n250 0.155672
R1928 VTAIL.n259 VTAIL.n258 0.155672
R1929 VTAIL.n215 VTAIL.n113 0.155672
R1930 VTAIL.n208 VTAIL.n113 0.155672
R1931 VTAIL.n208 VTAIL.n207 0.155672
R1932 VTAIL.n207 VTAIL.n117 0.155672
R1933 VTAIL.n200 VTAIL.n117 0.155672
R1934 VTAIL.n200 VTAIL.n199 0.155672
R1935 VTAIL.n199 VTAIL.n121 0.155672
R1936 VTAIL.n191 VTAIL.n121 0.155672
R1937 VTAIL.n191 VTAIL.n190 0.155672
R1938 VTAIL.n190 VTAIL.n125 0.155672
R1939 VTAIL.n183 VTAIL.n125 0.155672
R1940 VTAIL.n183 VTAIL.n182 0.155672
R1941 VTAIL.n182 VTAIL.n130 0.155672
R1942 VTAIL.n175 VTAIL.n130 0.155672
R1943 VTAIL.n175 VTAIL.n174 0.155672
R1944 VTAIL.n174 VTAIL.n134 0.155672
R1945 VTAIL.n167 VTAIL.n134 0.155672
R1946 VTAIL.n167 VTAIL.n166 0.155672
R1947 VTAIL.n166 VTAIL.n138 0.155672
R1948 VTAIL.n159 VTAIL.n138 0.155672
R1949 VTAIL.n159 VTAIL.n158 0.155672
R1950 VTAIL.n158 VTAIL.n142 0.155672
R1951 VTAIL.n151 VTAIL.n142 0.155672
R1952 VTAIL.n151 VTAIL.n150 0.155672
R1953 VDD1.n100 VDD1.n0 756.745
R1954 VDD1.n205 VDD1.n105 756.745
R1955 VDD1.n101 VDD1.n100 585
R1956 VDD1.n99 VDD1.n98 585
R1957 VDD1.n4 VDD1.n3 585
R1958 VDD1.n93 VDD1.n92 585
R1959 VDD1.n91 VDD1.n90 585
R1960 VDD1.n8 VDD1.n7 585
R1961 VDD1.n85 VDD1.n84 585
R1962 VDD1.n83 VDD1.n82 585
R1963 VDD1.n81 VDD1.n11 585
R1964 VDD1.n15 VDD1.n12 585
R1965 VDD1.n76 VDD1.n75 585
R1966 VDD1.n74 VDD1.n73 585
R1967 VDD1.n17 VDD1.n16 585
R1968 VDD1.n68 VDD1.n67 585
R1969 VDD1.n66 VDD1.n65 585
R1970 VDD1.n21 VDD1.n20 585
R1971 VDD1.n60 VDD1.n59 585
R1972 VDD1.n58 VDD1.n57 585
R1973 VDD1.n25 VDD1.n24 585
R1974 VDD1.n52 VDD1.n51 585
R1975 VDD1.n50 VDD1.n49 585
R1976 VDD1.n29 VDD1.n28 585
R1977 VDD1.n44 VDD1.n43 585
R1978 VDD1.n42 VDD1.n41 585
R1979 VDD1.n33 VDD1.n32 585
R1980 VDD1.n36 VDD1.n35 585
R1981 VDD1.n140 VDD1.n139 585
R1982 VDD1.n137 VDD1.n136 585
R1983 VDD1.n146 VDD1.n145 585
R1984 VDD1.n148 VDD1.n147 585
R1985 VDD1.n133 VDD1.n132 585
R1986 VDD1.n154 VDD1.n153 585
R1987 VDD1.n156 VDD1.n155 585
R1988 VDD1.n129 VDD1.n128 585
R1989 VDD1.n162 VDD1.n161 585
R1990 VDD1.n164 VDD1.n163 585
R1991 VDD1.n125 VDD1.n124 585
R1992 VDD1.n170 VDD1.n169 585
R1993 VDD1.n172 VDD1.n171 585
R1994 VDD1.n121 VDD1.n120 585
R1995 VDD1.n178 VDD1.n177 585
R1996 VDD1.n181 VDD1.n180 585
R1997 VDD1.n179 VDD1.n117 585
R1998 VDD1.n186 VDD1.n116 585
R1999 VDD1.n188 VDD1.n187 585
R2000 VDD1.n190 VDD1.n189 585
R2001 VDD1.n113 VDD1.n112 585
R2002 VDD1.n196 VDD1.n195 585
R2003 VDD1.n198 VDD1.n197 585
R2004 VDD1.n109 VDD1.n108 585
R2005 VDD1.n204 VDD1.n203 585
R2006 VDD1.n206 VDD1.n205 585
R2007 VDD1.t4 VDD1.n34 327.466
R2008 VDD1.t5 VDD1.n138 327.466
R2009 VDD1.n100 VDD1.n99 171.744
R2010 VDD1.n99 VDD1.n3 171.744
R2011 VDD1.n92 VDD1.n3 171.744
R2012 VDD1.n92 VDD1.n91 171.744
R2013 VDD1.n91 VDD1.n7 171.744
R2014 VDD1.n84 VDD1.n7 171.744
R2015 VDD1.n84 VDD1.n83 171.744
R2016 VDD1.n83 VDD1.n11 171.744
R2017 VDD1.n15 VDD1.n11 171.744
R2018 VDD1.n75 VDD1.n15 171.744
R2019 VDD1.n75 VDD1.n74 171.744
R2020 VDD1.n74 VDD1.n16 171.744
R2021 VDD1.n67 VDD1.n16 171.744
R2022 VDD1.n67 VDD1.n66 171.744
R2023 VDD1.n66 VDD1.n20 171.744
R2024 VDD1.n59 VDD1.n20 171.744
R2025 VDD1.n59 VDD1.n58 171.744
R2026 VDD1.n58 VDD1.n24 171.744
R2027 VDD1.n51 VDD1.n24 171.744
R2028 VDD1.n51 VDD1.n50 171.744
R2029 VDD1.n50 VDD1.n28 171.744
R2030 VDD1.n43 VDD1.n28 171.744
R2031 VDD1.n43 VDD1.n42 171.744
R2032 VDD1.n42 VDD1.n32 171.744
R2033 VDD1.n35 VDD1.n32 171.744
R2034 VDD1.n139 VDD1.n136 171.744
R2035 VDD1.n146 VDD1.n136 171.744
R2036 VDD1.n147 VDD1.n146 171.744
R2037 VDD1.n147 VDD1.n132 171.744
R2038 VDD1.n154 VDD1.n132 171.744
R2039 VDD1.n155 VDD1.n154 171.744
R2040 VDD1.n155 VDD1.n128 171.744
R2041 VDD1.n162 VDD1.n128 171.744
R2042 VDD1.n163 VDD1.n162 171.744
R2043 VDD1.n163 VDD1.n124 171.744
R2044 VDD1.n170 VDD1.n124 171.744
R2045 VDD1.n171 VDD1.n170 171.744
R2046 VDD1.n171 VDD1.n120 171.744
R2047 VDD1.n178 VDD1.n120 171.744
R2048 VDD1.n180 VDD1.n178 171.744
R2049 VDD1.n180 VDD1.n179 171.744
R2050 VDD1.n179 VDD1.n116 171.744
R2051 VDD1.n188 VDD1.n116 171.744
R2052 VDD1.n189 VDD1.n188 171.744
R2053 VDD1.n189 VDD1.n112 171.744
R2054 VDD1.n196 VDD1.n112 171.744
R2055 VDD1.n197 VDD1.n196 171.744
R2056 VDD1.n197 VDD1.n108 171.744
R2057 VDD1.n204 VDD1.n108 171.744
R2058 VDD1.n205 VDD1.n204 171.744
R2059 VDD1.n35 VDD1.t4 85.8723
R2060 VDD1.n139 VDD1.t5 85.8723
R2061 VDD1.n211 VDD1.n210 68.808
R2062 VDD1.n213 VDD1.n212 68.3847
R2063 VDD1 VDD1.n104 50.3577
R2064 VDD1.n211 VDD1.n209 50.2441
R2065 VDD1.n213 VDD1.n211 47.8199
R2066 VDD1.n36 VDD1.n34 16.3895
R2067 VDD1.n140 VDD1.n138 16.3895
R2068 VDD1.n82 VDD1.n81 13.1884
R2069 VDD1.n187 VDD1.n186 13.1884
R2070 VDD1.n85 VDD1.n10 12.8005
R2071 VDD1.n80 VDD1.n12 12.8005
R2072 VDD1.n37 VDD1.n33 12.8005
R2073 VDD1.n141 VDD1.n137 12.8005
R2074 VDD1.n185 VDD1.n117 12.8005
R2075 VDD1.n190 VDD1.n115 12.8005
R2076 VDD1.n86 VDD1.n8 12.0247
R2077 VDD1.n77 VDD1.n76 12.0247
R2078 VDD1.n41 VDD1.n40 12.0247
R2079 VDD1.n145 VDD1.n144 12.0247
R2080 VDD1.n182 VDD1.n181 12.0247
R2081 VDD1.n191 VDD1.n113 12.0247
R2082 VDD1.n90 VDD1.n89 11.249
R2083 VDD1.n73 VDD1.n14 11.249
R2084 VDD1.n44 VDD1.n31 11.249
R2085 VDD1.n148 VDD1.n135 11.249
R2086 VDD1.n177 VDD1.n119 11.249
R2087 VDD1.n195 VDD1.n194 11.249
R2088 VDD1.n93 VDD1.n6 10.4732
R2089 VDD1.n72 VDD1.n17 10.4732
R2090 VDD1.n45 VDD1.n29 10.4732
R2091 VDD1.n149 VDD1.n133 10.4732
R2092 VDD1.n176 VDD1.n121 10.4732
R2093 VDD1.n198 VDD1.n111 10.4732
R2094 VDD1.n94 VDD1.n4 9.69747
R2095 VDD1.n69 VDD1.n68 9.69747
R2096 VDD1.n49 VDD1.n48 9.69747
R2097 VDD1.n153 VDD1.n152 9.69747
R2098 VDD1.n173 VDD1.n172 9.69747
R2099 VDD1.n199 VDD1.n109 9.69747
R2100 VDD1.n104 VDD1.n103 9.45567
R2101 VDD1.n209 VDD1.n208 9.45567
R2102 VDD1.n62 VDD1.n61 9.3005
R2103 VDD1.n64 VDD1.n63 9.3005
R2104 VDD1.n19 VDD1.n18 9.3005
R2105 VDD1.n70 VDD1.n69 9.3005
R2106 VDD1.n72 VDD1.n71 9.3005
R2107 VDD1.n14 VDD1.n13 9.3005
R2108 VDD1.n78 VDD1.n77 9.3005
R2109 VDD1.n80 VDD1.n79 9.3005
R2110 VDD1.n103 VDD1.n102 9.3005
R2111 VDD1.n2 VDD1.n1 9.3005
R2112 VDD1.n97 VDD1.n96 9.3005
R2113 VDD1.n95 VDD1.n94 9.3005
R2114 VDD1.n6 VDD1.n5 9.3005
R2115 VDD1.n89 VDD1.n88 9.3005
R2116 VDD1.n87 VDD1.n86 9.3005
R2117 VDD1.n10 VDD1.n9 9.3005
R2118 VDD1.n23 VDD1.n22 9.3005
R2119 VDD1.n56 VDD1.n55 9.3005
R2120 VDD1.n54 VDD1.n53 9.3005
R2121 VDD1.n27 VDD1.n26 9.3005
R2122 VDD1.n48 VDD1.n47 9.3005
R2123 VDD1.n46 VDD1.n45 9.3005
R2124 VDD1.n31 VDD1.n30 9.3005
R2125 VDD1.n40 VDD1.n39 9.3005
R2126 VDD1.n38 VDD1.n37 9.3005
R2127 VDD1.n107 VDD1.n106 9.3005
R2128 VDD1.n202 VDD1.n201 9.3005
R2129 VDD1.n200 VDD1.n199 9.3005
R2130 VDD1.n111 VDD1.n110 9.3005
R2131 VDD1.n194 VDD1.n193 9.3005
R2132 VDD1.n192 VDD1.n191 9.3005
R2133 VDD1.n115 VDD1.n114 9.3005
R2134 VDD1.n160 VDD1.n159 9.3005
R2135 VDD1.n158 VDD1.n157 9.3005
R2136 VDD1.n131 VDD1.n130 9.3005
R2137 VDD1.n152 VDD1.n151 9.3005
R2138 VDD1.n150 VDD1.n149 9.3005
R2139 VDD1.n135 VDD1.n134 9.3005
R2140 VDD1.n144 VDD1.n143 9.3005
R2141 VDD1.n142 VDD1.n141 9.3005
R2142 VDD1.n127 VDD1.n126 9.3005
R2143 VDD1.n166 VDD1.n165 9.3005
R2144 VDD1.n168 VDD1.n167 9.3005
R2145 VDD1.n123 VDD1.n122 9.3005
R2146 VDD1.n174 VDD1.n173 9.3005
R2147 VDD1.n176 VDD1.n175 9.3005
R2148 VDD1.n119 VDD1.n118 9.3005
R2149 VDD1.n183 VDD1.n182 9.3005
R2150 VDD1.n185 VDD1.n184 9.3005
R2151 VDD1.n208 VDD1.n207 9.3005
R2152 VDD1.n98 VDD1.n97 8.92171
R2153 VDD1.n65 VDD1.n19 8.92171
R2154 VDD1.n52 VDD1.n27 8.92171
R2155 VDD1.n156 VDD1.n131 8.92171
R2156 VDD1.n169 VDD1.n123 8.92171
R2157 VDD1.n203 VDD1.n202 8.92171
R2158 VDD1.n101 VDD1.n2 8.14595
R2159 VDD1.n64 VDD1.n21 8.14595
R2160 VDD1.n53 VDD1.n25 8.14595
R2161 VDD1.n157 VDD1.n129 8.14595
R2162 VDD1.n168 VDD1.n125 8.14595
R2163 VDD1.n206 VDD1.n107 8.14595
R2164 VDD1.n102 VDD1.n0 7.3702
R2165 VDD1.n61 VDD1.n60 7.3702
R2166 VDD1.n57 VDD1.n56 7.3702
R2167 VDD1.n161 VDD1.n160 7.3702
R2168 VDD1.n165 VDD1.n164 7.3702
R2169 VDD1.n207 VDD1.n105 7.3702
R2170 VDD1.n104 VDD1.n0 6.59444
R2171 VDD1.n60 VDD1.n23 6.59444
R2172 VDD1.n57 VDD1.n23 6.59444
R2173 VDD1.n161 VDD1.n127 6.59444
R2174 VDD1.n164 VDD1.n127 6.59444
R2175 VDD1.n209 VDD1.n105 6.59444
R2176 VDD1.n102 VDD1.n101 5.81868
R2177 VDD1.n61 VDD1.n21 5.81868
R2178 VDD1.n56 VDD1.n25 5.81868
R2179 VDD1.n160 VDD1.n129 5.81868
R2180 VDD1.n165 VDD1.n125 5.81868
R2181 VDD1.n207 VDD1.n206 5.81868
R2182 VDD1.n98 VDD1.n2 5.04292
R2183 VDD1.n65 VDD1.n64 5.04292
R2184 VDD1.n53 VDD1.n52 5.04292
R2185 VDD1.n157 VDD1.n156 5.04292
R2186 VDD1.n169 VDD1.n168 5.04292
R2187 VDD1.n203 VDD1.n107 5.04292
R2188 VDD1.n97 VDD1.n4 4.26717
R2189 VDD1.n68 VDD1.n19 4.26717
R2190 VDD1.n49 VDD1.n27 4.26717
R2191 VDD1.n153 VDD1.n131 4.26717
R2192 VDD1.n172 VDD1.n123 4.26717
R2193 VDD1.n202 VDD1.n109 4.26717
R2194 VDD1.n38 VDD1.n34 3.70982
R2195 VDD1.n142 VDD1.n138 3.70982
R2196 VDD1.n94 VDD1.n93 3.49141
R2197 VDD1.n69 VDD1.n17 3.49141
R2198 VDD1.n48 VDD1.n29 3.49141
R2199 VDD1.n152 VDD1.n133 3.49141
R2200 VDD1.n173 VDD1.n121 3.49141
R2201 VDD1.n199 VDD1.n198 3.49141
R2202 VDD1.n90 VDD1.n6 2.71565
R2203 VDD1.n73 VDD1.n72 2.71565
R2204 VDD1.n45 VDD1.n44 2.71565
R2205 VDD1.n149 VDD1.n148 2.71565
R2206 VDD1.n177 VDD1.n176 2.71565
R2207 VDD1.n195 VDD1.n111 2.71565
R2208 VDD1.n89 VDD1.n8 1.93989
R2209 VDD1.n76 VDD1.n14 1.93989
R2210 VDD1.n41 VDD1.n31 1.93989
R2211 VDD1.n145 VDD1.n135 1.93989
R2212 VDD1.n181 VDD1.n119 1.93989
R2213 VDD1.n194 VDD1.n113 1.93989
R2214 VDD1.n212 VDD1.t1 1.7149
R2215 VDD1.n212 VDD1.t3 1.7149
R2216 VDD1.n210 VDD1.t0 1.7149
R2217 VDD1.n210 VDD1.t2 1.7149
R2218 VDD1.n86 VDD1.n85 1.16414
R2219 VDD1.n77 VDD1.n12 1.16414
R2220 VDD1.n40 VDD1.n33 1.16414
R2221 VDD1.n144 VDD1.n137 1.16414
R2222 VDD1.n182 VDD1.n117 1.16414
R2223 VDD1.n191 VDD1.n190 1.16414
R2224 VDD1 VDD1.n213 0.420759
R2225 VDD1.n82 VDD1.n10 0.388379
R2226 VDD1.n81 VDD1.n80 0.388379
R2227 VDD1.n37 VDD1.n36 0.388379
R2228 VDD1.n141 VDD1.n140 0.388379
R2229 VDD1.n186 VDD1.n185 0.388379
R2230 VDD1.n187 VDD1.n115 0.388379
R2231 VDD1.n103 VDD1.n1 0.155672
R2232 VDD1.n96 VDD1.n1 0.155672
R2233 VDD1.n96 VDD1.n95 0.155672
R2234 VDD1.n95 VDD1.n5 0.155672
R2235 VDD1.n88 VDD1.n5 0.155672
R2236 VDD1.n88 VDD1.n87 0.155672
R2237 VDD1.n87 VDD1.n9 0.155672
R2238 VDD1.n79 VDD1.n9 0.155672
R2239 VDD1.n79 VDD1.n78 0.155672
R2240 VDD1.n78 VDD1.n13 0.155672
R2241 VDD1.n71 VDD1.n13 0.155672
R2242 VDD1.n71 VDD1.n70 0.155672
R2243 VDD1.n70 VDD1.n18 0.155672
R2244 VDD1.n63 VDD1.n18 0.155672
R2245 VDD1.n63 VDD1.n62 0.155672
R2246 VDD1.n62 VDD1.n22 0.155672
R2247 VDD1.n55 VDD1.n22 0.155672
R2248 VDD1.n55 VDD1.n54 0.155672
R2249 VDD1.n54 VDD1.n26 0.155672
R2250 VDD1.n47 VDD1.n26 0.155672
R2251 VDD1.n47 VDD1.n46 0.155672
R2252 VDD1.n46 VDD1.n30 0.155672
R2253 VDD1.n39 VDD1.n30 0.155672
R2254 VDD1.n39 VDD1.n38 0.155672
R2255 VDD1.n143 VDD1.n142 0.155672
R2256 VDD1.n143 VDD1.n134 0.155672
R2257 VDD1.n150 VDD1.n134 0.155672
R2258 VDD1.n151 VDD1.n150 0.155672
R2259 VDD1.n151 VDD1.n130 0.155672
R2260 VDD1.n158 VDD1.n130 0.155672
R2261 VDD1.n159 VDD1.n158 0.155672
R2262 VDD1.n159 VDD1.n126 0.155672
R2263 VDD1.n166 VDD1.n126 0.155672
R2264 VDD1.n167 VDD1.n166 0.155672
R2265 VDD1.n167 VDD1.n122 0.155672
R2266 VDD1.n174 VDD1.n122 0.155672
R2267 VDD1.n175 VDD1.n174 0.155672
R2268 VDD1.n175 VDD1.n118 0.155672
R2269 VDD1.n183 VDD1.n118 0.155672
R2270 VDD1.n184 VDD1.n183 0.155672
R2271 VDD1.n184 VDD1.n114 0.155672
R2272 VDD1.n192 VDD1.n114 0.155672
R2273 VDD1.n193 VDD1.n192 0.155672
R2274 VDD1.n193 VDD1.n110 0.155672
R2275 VDD1.n200 VDD1.n110 0.155672
R2276 VDD1.n201 VDD1.n200 0.155672
R2277 VDD1.n201 VDD1.n106 0.155672
R2278 VDD1.n208 VDD1.n106 0.155672
R2279 VN.n2 VN.t2 272.935
R2280 VN.n14 VN.t0 272.935
R2281 VN.n3 VN.t5 241.766
R2282 VN.n10 VN.t1 241.766
R2283 VN.n15 VN.t4 241.766
R2284 VN.n22 VN.t3 241.766
R2285 VN.n21 VN.n12 161.3
R2286 VN.n20 VN.n19 161.3
R2287 VN.n18 VN.n13 161.3
R2288 VN.n17 VN.n16 161.3
R2289 VN.n9 VN.n0 161.3
R2290 VN.n8 VN.n7 161.3
R2291 VN.n6 VN.n1 161.3
R2292 VN.n5 VN.n4 161.3
R2293 VN.n11 VN.n10 87.7919
R2294 VN.n23 VN.n22 87.7919
R2295 VN.n3 VN.n2 57.9788
R2296 VN.n15 VN.n14 57.9788
R2297 VN.n8 VN.n1 54.1398
R2298 VN.n20 VN.n13 54.1398
R2299 VN VN.n23 51.4906
R2300 VN.n9 VN.n8 27.0143
R2301 VN.n21 VN.n20 27.0143
R2302 VN.n4 VN.n1 24.5923
R2303 VN.n16 VN.n13 24.5923
R2304 VN.n10 VN.n9 23.1168
R2305 VN.n22 VN.n21 23.1168
R2306 VN.n17 VN.n14 12.8269
R2307 VN.n5 VN.n2 12.8269
R2308 VN.n4 VN.n3 12.2964
R2309 VN.n16 VN.n15 12.2964
R2310 VN.n23 VN.n12 0.278335
R2311 VN.n11 VN.n0 0.278335
R2312 VN.n19 VN.n12 0.189894
R2313 VN.n19 VN.n18 0.189894
R2314 VN.n18 VN.n17 0.189894
R2315 VN.n6 VN.n5 0.189894
R2316 VN.n7 VN.n6 0.189894
R2317 VN.n7 VN.n0 0.189894
R2318 VN VN.n11 0.153485
R2319 VDD2.n207 VDD2.n107 756.745
R2320 VDD2.n100 VDD2.n0 756.745
R2321 VDD2.n208 VDD2.n207 585
R2322 VDD2.n206 VDD2.n205 585
R2323 VDD2.n111 VDD2.n110 585
R2324 VDD2.n200 VDD2.n199 585
R2325 VDD2.n198 VDD2.n197 585
R2326 VDD2.n115 VDD2.n114 585
R2327 VDD2.n192 VDD2.n191 585
R2328 VDD2.n190 VDD2.n189 585
R2329 VDD2.n188 VDD2.n118 585
R2330 VDD2.n122 VDD2.n119 585
R2331 VDD2.n183 VDD2.n182 585
R2332 VDD2.n181 VDD2.n180 585
R2333 VDD2.n124 VDD2.n123 585
R2334 VDD2.n175 VDD2.n174 585
R2335 VDD2.n173 VDD2.n172 585
R2336 VDD2.n128 VDD2.n127 585
R2337 VDD2.n167 VDD2.n166 585
R2338 VDD2.n165 VDD2.n164 585
R2339 VDD2.n132 VDD2.n131 585
R2340 VDD2.n159 VDD2.n158 585
R2341 VDD2.n157 VDD2.n156 585
R2342 VDD2.n136 VDD2.n135 585
R2343 VDD2.n151 VDD2.n150 585
R2344 VDD2.n149 VDD2.n148 585
R2345 VDD2.n140 VDD2.n139 585
R2346 VDD2.n143 VDD2.n142 585
R2347 VDD2.n35 VDD2.n34 585
R2348 VDD2.n32 VDD2.n31 585
R2349 VDD2.n41 VDD2.n40 585
R2350 VDD2.n43 VDD2.n42 585
R2351 VDD2.n28 VDD2.n27 585
R2352 VDD2.n49 VDD2.n48 585
R2353 VDD2.n51 VDD2.n50 585
R2354 VDD2.n24 VDD2.n23 585
R2355 VDD2.n57 VDD2.n56 585
R2356 VDD2.n59 VDD2.n58 585
R2357 VDD2.n20 VDD2.n19 585
R2358 VDD2.n65 VDD2.n64 585
R2359 VDD2.n67 VDD2.n66 585
R2360 VDD2.n16 VDD2.n15 585
R2361 VDD2.n73 VDD2.n72 585
R2362 VDD2.n76 VDD2.n75 585
R2363 VDD2.n74 VDD2.n12 585
R2364 VDD2.n81 VDD2.n11 585
R2365 VDD2.n83 VDD2.n82 585
R2366 VDD2.n85 VDD2.n84 585
R2367 VDD2.n8 VDD2.n7 585
R2368 VDD2.n91 VDD2.n90 585
R2369 VDD2.n93 VDD2.n92 585
R2370 VDD2.n4 VDD2.n3 585
R2371 VDD2.n99 VDD2.n98 585
R2372 VDD2.n101 VDD2.n100 585
R2373 VDD2.t2 VDD2.n141 327.466
R2374 VDD2.t3 VDD2.n33 327.466
R2375 VDD2.n207 VDD2.n206 171.744
R2376 VDD2.n206 VDD2.n110 171.744
R2377 VDD2.n199 VDD2.n110 171.744
R2378 VDD2.n199 VDD2.n198 171.744
R2379 VDD2.n198 VDD2.n114 171.744
R2380 VDD2.n191 VDD2.n114 171.744
R2381 VDD2.n191 VDD2.n190 171.744
R2382 VDD2.n190 VDD2.n118 171.744
R2383 VDD2.n122 VDD2.n118 171.744
R2384 VDD2.n182 VDD2.n122 171.744
R2385 VDD2.n182 VDD2.n181 171.744
R2386 VDD2.n181 VDD2.n123 171.744
R2387 VDD2.n174 VDD2.n123 171.744
R2388 VDD2.n174 VDD2.n173 171.744
R2389 VDD2.n173 VDD2.n127 171.744
R2390 VDD2.n166 VDD2.n127 171.744
R2391 VDD2.n166 VDD2.n165 171.744
R2392 VDD2.n165 VDD2.n131 171.744
R2393 VDD2.n158 VDD2.n131 171.744
R2394 VDD2.n158 VDD2.n157 171.744
R2395 VDD2.n157 VDD2.n135 171.744
R2396 VDD2.n150 VDD2.n135 171.744
R2397 VDD2.n150 VDD2.n149 171.744
R2398 VDD2.n149 VDD2.n139 171.744
R2399 VDD2.n142 VDD2.n139 171.744
R2400 VDD2.n34 VDD2.n31 171.744
R2401 VDD2.n41 VDD2.n31 171.744
R2402 VDD2.n42 VDD2.n41 171.744
R2403 VDD2.n42 VDD2.n27 171.744
R2404 VDD2.n49 VDD2.n27 171.744
R2405 VDD2.n50 VDD2.n49 171.744
R2406 VDD2.n50 VDD2.n23 171.744
R2407 VDD2.n57 VDD2.n23 171.744
R2408 VDD2.n58 VDD2.n57 171.744
R2409 VDD2.n58 VDD2.n19 171.744
R2410 VDD2.n65 VDD2.n19 171.744
R2411 VDD2.n66 VDD2.n65 171.744
R2412 VDD2.n66 VDD2.n15 171.744
R2413 VDD2.n73 VDD2.n15 171.744
R2414 VDD2.n75 VDD2.n73 171.744
R2415 VDD2.n75 VDD2.n74 171.744
R2416 VDD2.n74 VDD2.n11 171.744
R2417 VDD2.n83 VDD2.n11 171.744
R2418 VDD2.n84 VDD2.n83 171.744
R2419 VDD2.n84 VDD2.n7 171.744
R2420 VDD2.n91 VDD2.n7 171.744
R2421 VDD2.n92 VDD2.n91 171.744
R2422 VDD2.n92 VDD2.n3 171.744
R2423 VDD2.n99 VDD2.n3 171.744
R2424 VDD2.n100 VDD2.n99 171.744
R2425 VDD2.n142 VDD2.t2 85.8723
R2426 VDD2.n34 VDD2.t3 85.8723
R2427 VDD2.n106 VDD2.n105 68.808
R2428 VDD2 VDD2.n213 68.805
R2429 VDD2.n106 VDD2.n104 50.2441
R2430 VDD2.n212 VDD2.n211 48.8641
R2431 VDD2.n212 VDD2.n106 46.2799
R2432 VDD2.n143 VDD2.n141 16.3895
R2433 VDD2.n35 VDD2.n33 16.3895
R2434 VDD2.n189 VDD2.n188 13.1884
R2435 VDD2.n82 VDD2.n81 13.1884
R2436 VDD2.n192 VDD2.n117 12.8005
R2437 VDD2.n187 VDD2.n119 12.8005
R2438 VDD2.n144 VDD2.n140 12.8005
R2439 VDD2.n36 VDD2.n32 12.8005
R2440 VDD2.n80 VDD2.n12 12.8005
R2441 VDD2.n85 VDD2.n10 12.8005
R2442 VDD2.n193 VDD2.n115 12.0247
R2443 VDD2.n184 VDD2.n183 12.0247
R2444 VDD2.n148 VDD2.n147 12.0247
R2445 VDD2.n40 VDD2.n39 12.0247
R2446 VDD2.n77 VDD2.n76 12.0247
R2447 VDD2.n86 VDD2.n8 12.0247
R2448 VDD2.n197 VDD2.n196 11.249
R2449 VDD2.n180 VDD2.n121 11.249
R2450 VDD2.n151 VDD2.n138 11.249
R2451 VDD2.n43 VDD2.n30 11.249
R2452 VDD2.n72 VDD2.n14 11.249
R2453 VDD2.n90 VDD2.n89 11.249
R2454 VDD2.n200 VDD2.n113 10.4732
R2455 VDD2.n179 VDD2.n124 10.4732
R2456 VDD2.n152 VDD2.n136 10.4732
R2457 VDD2.n44 VDD2.n28 10.4732
R2458 VDD2.n71 VDD2.n16 10.4732
R2459 VDD2.n93 VDD2.n6 10.4732
R2460 VDD2.n201 VDD2.n111 9.69747
R2461 VDD2.n176 VDD2.n175 9.69747
R2462 VDD2.n156 VDD2.n155 9.69747
R2463 VDD2.n48 VDD2.n47 9.69747
R2464 VDD2.n68 VDD2.n67 9.69747
R2465 VDD2.n94 VDD2.n4 9.69747
R2466 VDD2.n211 VDD2.n210 9.45567
R2467 VDD2.n104 VDD2.n103 9.45567
R2468 VDD2.n169 VDD2.n168 9.3005
R2469 VDD2.n171 VDD2.n170 9.3005
R2470 VDD2.n126 VDD2.n125 9.3005
R2471 VDD2.n177 VDD2.n176 9.3005
R2472 VDD2.n179 VDD2.n178 9.3005
R2473 VDD2.n121 VDD2.n120 9.3005
R2474 VDD2.n185 VDD2.n184 9.3005
R2475 VDD2.n187 VDD2.n186 9.3005
R2476 VDD2.n210 VDD2.n209 9.3005
R2477 VDD2.n109 VDD2.n108 9.3005
R2478 VDD2.n204 VDD2.n203 9.3005
R2479 VDD2.n202 VDD2.n201 9.3005
R2480 VDD2.n113 VDD2.n112 9.3005
R2481 VDD2.n196 VDD2.n195 9.3005
R2482 VDD2.n194 VDD2.n193 9.3005
R2483 VDD2.n117 VDD2.n116 9.3005
R2484 VDD2.n130 VDD2.n129 9.3005
R2485 VDD2.n163 VDD2.n162 9.3005
R2486 VDD2.n161 VDD2.n160 9.3005
R2487 VDD2.n134 VDD2.n133 9.3005
R2488 VDD2.n155 VDD2.n154 9.3005
R2489 VDD2.n153 VDD2.n152 9.3005
R2490 VDD2.n138 VDD2.n137 9.3005
R2491 VDD2.n147 VDD2.n146 9.3005
R2492 VDD2.n145 VDD2.n144 9.3005
R2493 VDD2.n2 VDD2.n1 9.3005
R2494 VDD2.n97 VDD2.n96 9.3005
R2495 VDD2.n95 VDD2.n94 9.3005
R2496 VDD2.n6 VDD2.n5 9.3005
R2497 VDD2.n89 VDD2.n88 9.3005
R2498 VDD2.n87 VDD2.n86 9.3005
R2499 VDD2.n10 VDD2.n9 9.3005
R2500 VDD2.n55 VDD2.n54 9.3005
R2501 VDD2.n53 VDD2.n52 9.3005
R2502 VDD2.n26 VDD2.n25 9.3005
R2503 VDD2.n47 VDD2.n46 9.3005
R2504 VDD2.n45 VDD2.n44 9.3005
R2505 VDD2.n30 VDD2.n29 9.3005
R2506 VDD2.n39 VDD2.n38 9.3005
R2507 VDD2.n37 VDD2.n36 9.3005
R2508 VDD2.n22 VDD2.n21 9.3005
R2509 VDD2.n61 VDD2.n60 9.3005
R2510 VDD2.n63 VDD2.n62 9.3005
R2511 VDD2.n18 VDD2.n17 9.3005
R2512 VDD2.n69 VDD2.n68 9.3005
R2513 VDD2.n71 VDD2.n70 9.3005
R2514 VDD2.n14 VDD2.n13 9.3005
R2515 VDD2.n78 VDD2.n77 9.3005
R2516 VDD2.n80 VDD2.n79 9.3005
R2517 VDD2.n103 VDD2.n102 9.3005
R2518 VDD2.n205 VDD2.n204 8.92171
R2519 VDD2.n172 VDD2.n126 8.92171
R2520 VDD2.n159 VDD2.n134 8.92171
R2521 VDD2.n51 VDD2.n26 8.92171
R2522 VDD2.n64 VDD2.n18 8.92171
R2523 VDD2.n98 VDD2.n97 8.92171
R2524 VDD2.n208 VDD2.n109 8.14595
R2525 VDD2.n171 VDD2.n128 8.14595
R2526 VDD2.n160 VDD2.n132 8.14595
R2527 VDD2.n52 VDD2.n24 8.14595
R2528 VDD2.n63 VDD2.n20 8.14595
R2529 VDD2.n101 VDD2.n2 8.14595
R2530 VDD2.n209 VDD2.n107 7.3702
R2531 VDD2.n168 VDD2.n167 7.3702
R2532 VDD2.n164 VDD2.n163 7.3702
R2533 VDD2.n56 VDD2.n55 7.3702
R2534 VDD2.n60 VDD2.n59 7.3702
R2535 VDD2.n102 VDD2.n0 7.3702
R2536 VDD2.n211 VDD2.n107 6.59444
R2537 VDD2.n167 VDD2.n130 6.59444
R2538 VDD2.n164 VDD2.n130 6.59444
R2539 VDD2.n56 VDD2.n22 6.59444
R2540 VDD2.n59 VDD2.n22 6.59444
R2541 VDD2.n104 VDD2.n0 6.59444
R2542 VDD2.n209 VDD2.n208 5.81868
R2543 VDD2.n168 VDD2.n128 5.81868
R2544 VDD2.n163 VDD2.n132 5.81868
R2545 VDD2.n55 VDD2.n24 5.81868
R2546 VDD2.n60 VDD2.n20 5.81868
R2547 VDD2.n102 VDD2.n101 5.81868
R2548 VDD2.n205 VDD2.n109 5.04292
R2549 VDD2.n172 VDD2.n171 5.04292
R2550 VDD2.n160 VDD2.n159 5.04292
R2551 VDD2.n52 VDD2.n51 5.04292
R2552 VDD2.n64 VDD2.n63 5.04292
R2553 VDD2.n98 VDD2.n2 5.04292
R2554 VDD2.n204 VDD2.n111 4.26717
R2555 VDD2.n175 VDD2.n126 4.26717
R2556 VDD2.n156 VDD2.n134 4.26717
R2557 VDD2.n48 VDD2.n26 4.26717
R2558 VDD2.n67 VDD2.n18 4.26717
R2559 VDD2.n97 VDD2.n4 4.26717
R2560 VDD2.n145 VDD2.n141 3.70982
R2561 VDD2.n37 VDD2.n33 3.70982
R2562 VDD2.n201 VDD2.n200 3.49141
R2563 VDD2.n176 VDD2.n124 3.49141
R2564 VDD2.n155 VDD2.n136 3.49141
R2565 VDD2.n47 VDD2.n28 3.49141
R2566 VDD2.n68 VDD2.n16 3.49141
R2567 VDD2.n94 VDD2.n93 3.49141
R2568 VDD2.n197 VDD2.n113 2.71565
R2569 VDD2.n180 VDD2.n179 2.71565
R2570 VDD2.n152 VDD2.n151 2.71565
R2571 VDD2.n44 VDD2.n43 2.71565
R2572 VDD2.n72 VDD2.n71 2.71565
R2573 VDD2.n90 VDD2.n6 2.71565
R2574 VDD2.n196 VDD2.n115 1.93989
R2575 VDD2.n183 VDD2.n121 1.93989
R2576 VDD2.n148 VDD2.n138 1.93989
R2577 VDD2.n40 VDD2.n30 1.93989
R2578 VDD2.n76 VDD2.n14 1.93989
R2579 VDD2.n89 VDD2.n8 1.93989
R2580 VDD2.n213 VDD2.t1 1.7149
R2581 VDD2.n213 VDD2.t5 1.7149
R2582 VDD2.n105 VDD2.t0 1.7149
R2583 VDD2.n105 VDD2.t4 1.7149
R2584 VDD2 VDD2.n212 1.49403
R2585 VDD2.n193 VDD2.n192 1.16414
R2586 VDD2.n184 VDD2.n119 1.16414
R2587 VDD2.n147 VDD2.n140 1.16414
R2588 VDD2.n39 VDD2.n32 1.16414
R2589 VDD2.n77 VDD2.n12 1.16414
R2590 VDD2.n86 VDD2.n85 1.16414
R2591 VDD2.n189 VDD2.n117 0.388379
R2592 VDD2.n188 VDD2.n187 0.388379
R2593 VDD2.n144 VDD2.n143 0.388379
R2594 VDD2.n36 VDD2.n35 0.388379
R2595 VDD2.n81 VDD2.n80 0.388379
R2596 VDD2.n82 VDD2.n10 0.388379
R2597 VDD2.n210 VDD2.n108 0.155672
R2598 VDD2.n203 VDD2.n108 0.155672
R2599 VDD2.n203 VDD2.n202 0.155672
R2600 VDD2.n202 VDD2.n112 0.155672
R2601 VDD2.n195 VDD2.n112 0.155672
R2602 VDD2.n195 VDD2.n194 0.155672
R2603 VDD2.n194 VDD2.n116 0.155672
R2604 VDD2.n186 VDD2.n116 0.155672
R2605 VDD2.n186 VDD2.n185 0.155672
R2606 VDD2.n185 VDD2.n120 0.155672
R2607 VDD2.n178 VDD2.n120 0.155672
R2608 VDD2.n178 VDD2.n177 0.155672
R2609 VDD2.n177 VDD2.n125 0.155672
R2610 VDD2.n170 VDD2.n125 0.155672
R2611 VDD2.n170 VDD2.n169 0.155672
R2612 VDD2.n169 VDD2.n129 0.155672
R2613 VDD2.n162 VDD2.n129 0.155672
R2614 VDD2.n162 VDD2.n161 0.155672
R2615 VDD2.n161 VDD2.n133 0.155672
R2616 VDD2.n154 VDD2.n133 0.155672
R2617 VDD2.n154 VDD2.n153 0.155672
R2618 VDD2.n153 VDD2.n137 0.155672
R2619 VDD2.n146 VDD2.n137 0.155672
R2620 VDD2.n146 VDD2.n145 0.155672
R2621 VDD2.n38 VDD2.n37 0.155672
R2622 VDD2.n38 VDD2.n29 0.155672
R2623 VDD2.n45 VDD2.n29 0.155672
R2624 VDD2.n46 VDD2.n45 0.155672
R2625 VDD2.n46 VDD2.n25 0.155672
R2626 VDD2.n53 VDD2.n25 0.155672
R2627 VDD2.n54 VDD2.n53 0.155672
R2628 VDD2.n54 VDD2.n21 0.155672
R2629 VDD2.n61 VDD2.n21 0.155672
R2630 VDD2.n62 VDD2.n61 0.155672
R2631 VDD2.n62 VDD2.n17 0.155672
R2632 VDD2.n69 VDD2.n17 0.155672
R2633 VDD2.n70 VDD2.n69 0.155672
R2634 VDD2.n70 VDD2.n13 0.155672
R2635 VDD2.n78 VDD2.n13 0.155672
R2636 VDD2.n79 VDD2.n78 0.155672
R2637 VDD2.n79 VDD2.n9 0.155672
R2638 VDD2.n87 VDD2.n9 0.155672
R2639 VDD2.n88 VDD2.n87 0.155672
R2640 VDD2.n88 VDD2.n5 0.155672
R2641 VDD2.n95 VDD2.n5 0.155672
R2642 VDD2.n96 VDD2.n95 0.155672
R2643 VDD2.n96 VDD2.n1 0.155672
R2644 VDD2.n103 VDD2.n1 0.155672
C0 w_n2746_n4760# VP 5.50952f
C1 w_n2746_n4760# VDD1 2.61007f
C2 VN VTAIL 9.395491f
C3 w_n2746_n4760# VDD2 2.67251f
C4 B VP 1.68792f
C5 VDD1 B 2.44193f
C6 w_n2746_n4760# VTAIL 3.92611f
C7 VDD2 B 2.499f
C8 VDD1 VP 9.93398f
C9 w_n2746_n4760# VN 5.15648f
C10 VDD2 VP 0.399223f
C11 VDD1 VDD2 1.15612f
C12 B VTAIL 4.85126f
C13 VP VTAIL 9.41f
C14 VDD1 VTAIL 10.633901f
C15 B VN 1.10205f
C16 VDD2 VTAIL 10.6769f
C17 VP VN 7.52278f
C18 VDD1 VN 0.15012f
C19 VDD2 VN 9.68987f
C20 w_n2746_n4760# B 10.6466f
C21 VDD2 VSUBS 1.91943f
C22 VDD1 VSUBS 1.761355f
C23 VTAIL VSUBS 1.316827f
C24 VN VSUBS 5.5714f
C25 VP VSUBS 2.650193f
C26 B VSUBS 4.523979f
C27 w_n2746_n4760# VSUBS 0.159718p
C28 VDD2.n0 VSUBS 0.029847f
C29 VDD2.n1 VSUBS 0.026852f
C30 VDD2.n2 VSUBS 0.014429f
C31 VDD2.n3 VSUBS 0.034105f
C32 VDD2.n4 VSUBS 0.015278f
C33 VDD2.n5 VSUBS 0.026852f
C34 VDD2.n6 VSUBS 0.014429f
C35 VDD2.n7 VSUBS 0.034105f
C36 VDD2.n8 VSUBS 0.015278f
C37 VDD2.n9 VSUBS 0.026852f
C38 VDD2.n10 VSUBS 0.014429f
C39 VDD2.n11 VSUBS 0.034105f
C40 VDD2.n12 VSUBS 0.015278f
C41 VDD2.n13 VSUBS 0.026852f
C42 VDD2.n14 VSUBS 0.014429f
C43 VDD2.n15 VSUBS 0.034105f
C44 VDD2.n16 VSUBS 0.015278f
C45 VDD2.n17 VSUBS 0.026852f
C46 VDD2.n18 VSUBS 0.014429f
C47 VDD2.n19 VSUBS 0.034105f
C48 VDD2.n20 VSUBS 0.015278f
C49 VDD2.n21 VSUBS 0.026852f
C50 VDD2.n22 VSUBS 0.014429f
C51 VDD2.n23 VSUBS 0.034105f
C52 VDD2.n24 VSUBS 0.015278f
C53 VDD2.n25 VSUBS 0.026852f
C54 VDD2.n26 VSUBS 0.014429f
C55 VDD2.n27 VSUBS 0.034105f
C56 VDD2.n28 VSUBS 0.015278f
C57 VDD2.n29 VSUBS 0.026852f
C58 VDD2.n30 VSUBS 0.014429f
C59 VDD2.n31 VSUBS 0.034105f
C60 VDD2.n32 VSUBS 0.015278f
C61 VDD2.n33 VSUBS 0.220645f
C62 VDD2.t3 VSUBS 0.073276f
C63 VDD2.n34 VSUBS 0.025579f
C64 VDD2.n35 VSUBS 0.021696f
C65 VDD2.n36 VSUBS 0.014429f
C66 VDD2.n37 VSUBS 2.19726f
C67 VDD2.n38 VSUBS 0.026852f
C68 VDD2.n39 VSUBS 0.014429f
C69 VDD2.n40 VSUBS 0.015278f
C70 VDD2.n41 VSUBS 0.034105f
C71 VDD2.n42 VSUBS 0.034105f
C72 VDD2.n43 VSUBS 0.015278f
C73 VDD2.n44 VSUBS 0.014429f
C74 VDD2.n45 VSUBS 0.026852f
C75 VDD2.n46 VSUBS 0.026852f
C76 VDD2.n47 VSUBS 0.014429f
C77 VDD2.n48 VSUBS 0.015278f
C78 VDD2.n49 VSUBS 0.034105f
C79 VDD2.n50 VSUBS 0.034105f
C80 VDD2.n51 VSUBS 0.015278f
C81 VDD2.n52 VSUBS 0.014429f
C82 VDD2.n53 VSUBS 0.026852f
C83 VDD2.n54 VSUBS 0.026852f
C84 VDD2.n55 VSUBS 0.014429f
C85 VDD2.n56 VSUBS 0.015278f
C86 VDD2.n57 VSUBS 0.034105f
C87 VDD2.n58 VSUBS 0.034105f
C88 VDD2.n59 VSUBS 0.015278f
C89 VDD2.n60 VSUBS 0.014429f
C90 VDD2.n61 VSUBS 0.026852f
C91 VDD2.n62 VSUBS 0.026852f
C92 VDD2.n63 VSUBS 0.014429f
C93 VDD2.n64 VSUBS 0.015278f
C94 VDD2.n65 VSUBS 0.034105f
C95 VDD2.n66 VSUBS 0.034105f
C96 VDD2.n67 VSUBS 0.015278f
C97 VDD2.n68 VSUBS 0.014429f
C98 VDD2.n69 VSUBS 0.026852f
C99 VDD2.n70 VSUBS 0.026852f
C100 VDD2.n71 VSUBS 0.014429f
C101 VDD2.n72 VSUBS 0.015278f
C102 VDD2.n73 VSUBS 0.034105f
C103 VDD2.n74 VSUBS 0.034105f
C104 VDD2.n75 VSUBS 0.034105f
C105 VDD2.n76 VSUBS 0.015278f
C106 VDD2.n77 VSUBS 0.014429f
C107 VDD2.n78 VSUBS 0.026852f
C108 VDD2.n79 VSUBS 0.026852f
C109 VDD2.n80 VSUBS 0.014429f
C110 VDD2.n81 VSUBS 0.014853f
C111 VDD2.n82 VSUBS 0.014853f
C112 VDD2.n83 VSUBS 0.034105f
C113 VDD2.n84 VSUBS 0.034105f
C114 VDD2.n85 VSUBS 0.015278f
C115 VDD2.n86 VSUBS 0.014429f
C116 VDD2.n87 VSUBS 0.026852f
C117 VDD2.n88 VSUBS 0.026852f
C118 VDD2.n89 VSUBS 0.014429f
C119 VDD2.n90 VSUBS 0.015278f
C120 VDD2.n91 VSUBS 0.034105f
C121 VDD2.n92 VSUBS 0.034105f
C122 VDD2.n93 VSUBS 0.015278f
C123 VDD2.n94 VSUBS 0.014429f
C124 VDD2.n95 VSUBS 0.026852f
C125 VDD2.n96 VSUBS 0.026852f
C126 VDD2.n97 VSUBS 0.014429f
C127 VDD2.n98 VSUBS 0.015278f
C128 VDD2.n99 VSUBS 0.034105f
C129 VDD2.n100 VSUBS 0.083732f
C130 VDD2.n101 VSUBS 0.015278f
C131 VDD2.n102 VSUBS 0.014429f
C132 VDD2.n103 VSUBS 0.062067f
C133 VDD2.n104 VSUBS 0.065413f
C134 VDD2.t0 VSUBS 0.402314f
C135 VDD2.t4 VSUBS 0.402314f
C136 VDD2.n105 VSUBS 3.36648f
C137 VDD2.n106 VSUBS 3.32435f
C138 VDD2.n107 VSUBS 0.029847f
C139 VDD2.n108 VSUBS 0.026852f
C140 VDD2.n109 VSUBS 0.014429f
C141 VDD2.n110 VSUBS 0.034105f
C142 VDD2.n111 VSUBS 0.015278f
C143 VDD2.n112 VSUBS 0.026852f
C144 VDD2.n113 VSUBS 0.014429f
C145 VDD2.n114 VSUBS 0.034105f
C146 VDD2.n115 VSUBS 0.015278f
C147 VDD2.n116 VSUBS 0.026852f
C148 VDD2.n117 VSUBS 0.014429f
C149 VDD2.n118 VSUBS 0.034105f
C150 VDD2.n119 VSUBS 0.015278f
C151 VDD2.n120 VSUBS 0.026852f
C152 VDD2.n121 VSUBS 0.014429f
C153 VDD2.n122 VSUBS 0.034105f
C154 VDD2.n123 VSUBS 0.034105f
C155 VDD2.n124 VSUBS 0.015278f
C156 VDD2.n125 VSUBS 0.026852f
C157 VDD2.n126 VSUBS 0.014429f
C158 VDD2.n127 VSUBS 0.034105f
C159 VDD2.n128 VSUBS 0.015278f
C160 VDD2.n129 VSUBS 0.026852f
C161 VDD2.n130 VSUBS 0.014429f
C162 VDD2.n131 VSUBS 0.034105f
C163 VDD2.n132 VSUBS 0.015278f
C164 VDD2.n133 VSUBS 0.026852f
C165 VDD2.n134 VSUBS 0.014429f
C166 VDD2.n135 VSUBS 0.034105f
C167 VDD2.n136 VSUBS 0.015278f
C168 VDD2.n137 VSUBS 0.026852f
C169 VDD2.n138 VSUBS 0.014429f
C170 VDD2.n139 VSUBS 0.034105f
C171 VDD2.n140 VSUBS 0.015278f
C172 VDD2.n141 VSUBS 0.220645f
C173 VDD2.t2 VSUBS 0.073276f
C174 VDD2.n142 VSUBS 0.025579f
C175 VDD2.n143 VSUBS 0.021696f
C176 VDD2.n144 VSUBS 0.014429f
C177 VDD2.n145 VSUBS 2.19726f
C178 VDD2.n146 VSUBS 0.026852f
C179 VDD2.n147 VSUBS 0.014429f
C180 VDD2.n148 VSUBS 0.015278f
C181 VDD2.n149 VSUBS 0.034105f
C182 VDD2.n150 VSUBS 0.034105f
C183 VDD2.n151 VSUBS 0.015278f
C184 VDD2.n152 VSUBS 0.014429f
C185 VDD2.n153 VSUBS 0.026852f
C186 VDD2.n154 VSUBS 0.026852f
C187 VDD2.n155 VSUBS 0.014429f
C188 VDD2.n156 VSUBS 0.015278f
C189 VDD2.n157 VSUBS 0.034105f
C190 VDD2.n158 VSUBS 0.034105f
C191 VDD2.n159 VSUBS 0.015278f
C192 VDD2.n160 VSUBS 0.014429f
C193 VDD2.n161 VSUBS 0.026852f
C194 VDD2.n162 VSUBS 0.026852f
C195 VDD2.n163 VSUBS 0.014429f
C196 VDD2.n164 VSUBS 0.015278f
C197 VDD2.n165 VSUBS 0.034105f
C198 VDD2.n166 VSUBS 0.034105f
C199 VDD2.n167 VSUBS 0.015278f
C200 VDD2.n168 VSUBS 0.014429f
C201 VDD2.n169 VSUBS 0.026852f
C202 VDD2.n170 VSUBS 0.026852f
C203 VDD2.n171 VSUBS 0.014429f
C204 VDD2.n172 VSUBS 0.015278f
C205 VDD2.n173 VSUBS 0.034105f
C206 VDD2.n174 VSUBS 0.034105f
C207 VDD2.n175 VSUBS 0.015278f
C208 VDD2.n176 VSUBS 0.014429f
C209 VDD2.n177 VSUBS 0.026852f
C210 VDD2.n178 VSUBS 0.026852f
C211 VDD2.n179 VSUBS 0.014429f
C212 VDD2.n180 VSUBS 0.015278f
C213 VDD2.n181 VSUBS 0.034105f
C214 VDD2.n182 VSUBS 0.034105f
C215 VDD2.n183 VSUBS 0.015278f
C216 VDD2.n184 VSUBS 0.014429f
C217 VDD2.n185 VSUBS 0.026852f
C218 VDD2.n186 VSUBS 0.026852f
C219 VDD2.n187 VSUBS 0.014429f
C220 VDD2.n188 VSUBS 0.014853f
C221 VDD2.n189 VSUBS 0.014853f
C222 VDD2.n190 VSUBS 0.034105f
C223 VDD2.n191 VSUBS 0.034105f
C224 VDD2.n192 VSUBS 0.015278f
C225 VDD2.n193 VSUBS 0.014429f
C226 VDD2.n194 VSUBS 0.026852f
C227 VDD2.n195 VSUBS 0.026852f
C228 VDD2.n196 VSUBS 0.014429f
C229 VDD2.n197 VSUBS 0.015278f
C230 VDD2.n198 VSUBS 0.034105f
C231 VDD2.n199 VSUBS 0.034105f
C232 VDD2.n200 VSUBS 0.015278f
C233 VDD2.n201 VSUBS 0.014429f
C234 VDD2.n202 VSUBS 0.026852f
C235 VDD2.n203 VSUBS 0.026852f
C236 VDD2.n204 VSUBS 0.014429f
C237 VDD2.n205 VSUBS 0.015278f
C238 VDD2.n206 VSUBS 0.034105f
C239 VDD2.n207 VSUBS 0.083732f
C240 VDD2.n208 VSUBS 0.015278f
C241 VDD2.n209 VSUBS 0.014429f
C242 VDD2.n210 VSUBS 0.062067f
C243 VDD2.n211 VSUBS 0.060701f
C244 VDD2.n212 VSUBS 3.115f
C245 VDD2.t1 VSUBS 0.402314f
C246 VDD2.t5 VSUBS 0.402314f
C247 VDD2.n213 VSUBS 3.36643f
C248 VN.n0 VSUBS 0.043083f
C249 VN.t1 VSUBS 3.2242f
C250 VN.n1 VSUBS 0.05701f
C251 VN.t2 VSUBS 3.37036f
C252 VN.n2 VSUBS 1.2092f
C253 VN.t5 VSUBS 3.2242f
C254 VN.n3 VSUBS 1.19871f
C255 VN.n4 VSUBS 0.045643f
C256 VN.n5 VSUBS 0.241396f
C257 VN.n6 VSUBS 0.03268f
C258 VN.n7 VSUBS 0.03268f
C259 VN.n8 VSUBS 0.035587f
C260 VN.n9 VSUBS 0.061221f
C261 VN.n10 VSUBS 1.22436f
C262 VN.n11 VSUBS 0.036013f
C263 VN.n12 VSUBS 0.043083f
C264 VN.t3 VSUBS 3.2242f
C265 VN.n13 VSUBS 0.05701f
C266 VN.t0 VSUBS 3.37036f
C267 VN.n14 VSUBS 1.2092f
C268 VN.t4 VSUBS 3.2242f
C269 VN.n15 VSUBS 1.19871f
C270 VN.n16 VSUBS 0.045643f
C271 VN.n17 VSUBS 0.241396f
C272 VN.n18 VSUBS 0.03268f
C273 VN.n19 VSUBS 0.03268f
C274 VN.n20 VSUBS 0.035587f
C275 VN.n21 VSUBS 0.061221f
C276 VN.n22 VSUBS 1.22436f
C277 VN.n23 VSUBS 1.8827f
C278 VDD1.n0 VSUBS 0.029616f
C279 VDD1.n1 VSUBS 0.026644f
C280 VDD1.n2 VSUBS 0.014317f
C281 VDD1.n3 VSUBS 0.03384f
C282 VDD1.n4 VSUBS 0.015159f
C283 VDD1.n5 VSUBS 0.026644f
C284 VDD1.n6 VSUBS 0.014317f
C285 VDD1.n7 VSUBS 0.03384f
C286 VDD1.n8 VSUBS 0.015159f
C287 VDD1.n9 VSUBS 0.026644f
C288 VDD1.n10 VSUBS 0.014317f
C289 VDD1.n11 VSUBS 0.03384f
C290 VDD1.n12 VSUBS 0.015159f
C291 VDD1.n13 VSUBS 0.026644f
C292 VDD1.n14 VSUBS 0.014317f
C293 VDD1.n15 VSUBS 0.03384f
C294 VDD1.n16 VSUBS 0.03384f
C295 VDD1.n17 VSUBS 0.015159f
C296 VDD1.n18 VSUBS 0.026644f
C297 VDD1.n19 VSUBS 0.014317f
C298 VDD1.n20 VSUBS 0.03384f
C299 VDD1.n21 VSUBS 0.015159f
C300 VDD1.n22 VSUBS 0.026644f
C301 VDD1.n23 VSUBS 0.014317f
C302 VDD1.n24 VSUBS 0.03384f
C303 VDD1.n25 VSUBS 0.015159f
C304 VDD1.n26 VSUBS 0.026644f
C305 VDD1.n27 VSUBS 0.014317f
C306 VDD1.n28 VSUBS 0.03384f
C307 VDD1.n29 VSUBS 0.015159f
C308 VDD1.n30 VSUBS 0.026644f
C309 VDD1.n31 VSUBS 0.014317f
C310 VDD1.n32 VSUBS 0.03384f
C311 VDD1.n33 VSUBS 0.015159f
C312 VDD1.n34 VSUBS 0.218935f
C313 VDD1.t4 VSUBS 0.072708f
C314 VDD1.n35 VSUBS 0.02538f
C315 VDD1.n36 VSUBS 0.021528f
C316 VDD1.n37 VSUBS 0.014317f
C317 VDD1.n38 VSUBS 2.18023f
C318 VDD1.n39 VSUBS 0.026644f
C319 VDD1.n40 VSUBS 0.014317f
C320 VDD1.n41 VSUBS 0.015159f
C321 VDD1.n42 VSUBS 0.03384f
C322 VDD1.n43 VSUBS 0.03384f
C323 VDD1.n44 VSUBS 0.015159f
C324 VDD1.n45 VSUBS 0.014317f
C325 VDD1.n46 VSUBS 0.026644f
C326 VDD1.n47 VSUBS 0.026644f
C327 VDD1.n48 VSUBS 0.014317f
C328 VDD1.n49 VSUBS 0.015159f
C329 VDD1.n50 VSUBS 0.03384f
C330 VDD1.n51 VSUBS 0.03384f
C331 VDD1.n52 VSUBS 0.015159f
C332 VDD1.n53 VSUBS 0.014317f
C333 VDD1.n54 VSUBS 0.026644f
C334 VDD1.n55 VSUBS 0.026644f
C335 VDD1.n56 VSUBS 0.014317f
C336 VDD1.n57 VSUBS 0.015159f
C337 VDD1.n58 VSUBS 0.03384f
C338 VDD1.n59 VSUBS 0.03384f
C339 VDD1.n60 VSUBS 0.015159f
C340 VDD1.n61 VSUBS 0.014317f
C341 VDD1.n62 VSUBS 0.026644f
C342 VDD1.n63 VSUBS 0.026644f
C343 VDD1.n64 VSUBS 0.014317f
C344 VDD1.n65 VSUBS 0.015159f
C345 VDD1.n66 VSUBS 0.03384f
C346 VDD1.n67 VSUBS 0.03384f
C347 VDD1.n68 VSUBS 0.015159f
C348 VDD1.n69 VSUBS 0.014317f
C349 VDD1.n70 VSUBS 0.026644f
C350 VDD1.n71 VSUBS 0.026644f
C351 VDD1.n72 VSUBS 0.014317f
C352 VDD1.n73 VSUBS 0.015159f
C353 VDD1.n74 VSUBS 0.03384f
C354 VDD1.n75 VSUBS 0.03384f
C355 VDD1.n76 VSUBS 0.015159f
C356 VDD1.n77 VSUBS 0.014317f
C357 VDD1.n78 VSUBS 0.026644f
C358 VDD1.n79 VSUBS 0.026644f
C359 VDD1.n80 VSUBS 0.014317f
C360 VDD1.n81 VSUBS 0.014738f
C361 VDD1.n82 VSUBS 0.014738f
C362 VDD1.n83 VSUBS 0.03384f
C363 VDD1.n84 VSUBS 0.03384f
C364 VDD1.n85 VSUBS 0.015159f
C365 VDD1.n86 VSUBS 0.014317f
C366 VDD1.n87 VSUBS 0.026644f
C367 VDD1.n88 VSUBS 0.026644f
C368 VDD1.n89 VSUBS 0.014317f
C369 VDD1.n90 VSUBS 0.015159f
C370 VDD1.n91 VSUBS 0.03384f
C371 VDD1.n92 VSUBS 0.03384f
C372 VDD1.n93 VSUBS 0.015159f
C373 VDD1.n94 VSUBS 0.014317f
C374 VDD1.n95 VSUBS 0.026644f
C375 VDD1.n96 VSUBS 0.026644f
C376 VDD1.n97 VSUBS 0.014317f
C377 VDD1.n98 VSUBS 0.015159f
C378 VDD1.n99 VSUBS 0.03384f
C379 VDD1.n100 VSUBS 0.083084f
C380 VDD1.n101 VSUBS 0.015159f
C381 VDD1.n102 VSUBS 0.014317f
C382 VDD1.n103 VSUBS 0.061585f
C383 VDD1.n104 VSUBS 0.065555f
C384 VDD1.n105 VSUBS 0.029616f
C385 VDD1.n106 VSUBS 0.026644f
C386 VDD1.n107 VSUBS 0.014317f
C387 VDD1.n108 VSUBS 0.03384f
C388 VDD1.n109 VSUBS 0.015159f
C389 VDD1.n110 VSUBS 0.026644f
C390 VDD1.n111 VSUBS 0.014317f
C391 VDD1.n112 VSUBS 0.03384f
C392 VDD1.n113 VSUBS 0.015159f
C393 VDD1.n114 VSUBS 0.026644f
C394 VDD1.n115 VSUBS 0.014317f
C395 VDD1.n116 VSUBS 0.03384f
C396 VDD1.n117 VSUBS 0.015159f
C397 VDD1.n118 VSUBS 0.026644f
C398 VDD1.n119 VSUBS 0.014317f
C399 VDD1.n120 VSUBS 0.03384f
C400 VDD1.n121 VSUBS 0.015159f
C401 VDD1.n122 VSUBS 0.026644f
C402 VDD1.n123 VSUBS 0.014317f
C403 VDD1.n124 VSUBS 0.03384f
C404 VDD1.n125 VSUBS 0.015159f
C405 VDD1.n126 VSUBS 0.026644f
C406 VDD1.n127 VSUBS 0.014317f
C407 VDD1.n128 VSUBS 0.03384f
C408 VDD1.n129 VSUBS 0.015159f
C409 VDD1.n130 VSUBS 0.026644f
C410 VDD1.n131 VSUBS 0.014317f
C411 VDD1.n132 VSUBS 0.03384f
C412 VDD1.n133 VSUBS 0.015159f
C413 VDD1.n134 VSUBS 0.026644f
C414 VDD1.n135 VSUBS 0.014317f
C415 VDD1.n136 VSUBS 0.03384f
C416 VDD1.n137 VSUBS 0.015159f
C417 VDD1.n138 VSUBS 0.218935f
C418 VDD1.t5 VSUBS 0.072708f
C419 VDD1.n139 VSUBS 0.02538f
C420 VDD1.n140 VSUBS 0.021528f
C421 VDD1.n141 VSUBS 0.014317f
C422 VDD1.n142 VSUBS 2.18023f
C423 VDD1.n143 VSUBS 0.026644f
C424 VDD1.n144 VSUBS 0.014317f
C425 VDD1.n145 VSUBS 0.015159f
C426 VDD1.n146 VSUBS 0.03384f
C427 VDD1.n147 VSUBS 0.03384f
C428 VDD1.n148 VSUBS 0.015159f
C429 VDD1.n149 VSUBS 0.014317f
C430 VDD1.n150 VSUBS 0.026644f
C431 VDD1.n151 VSUBS 0.026644f
C432 VDD1.n152 VSUBS 0.014317f
C433 VDD1.n153 VSUBS 0.015159f
C434 VDD1.n154 VSUBS 0.03384f
C435 VDD1.n155 VSUBS 0.03384f
C436 VDD1.n156 VSUBS 0.015159f
C437 VDD1.n157 VSUBS 0.014317f
C438 VDD1.n158 VSUBS 0.026644f
C439 VDD1.n159 VSUBS 0.026644f
C440 VDD1.n160 VSUBS 0.014317f
C441 VDD1.n161 VSUBS 0.015159f
C442 VDD1.n162 VSUBS 0.03384f
C443 VDD1.n163 VSUBS 0.03384f
C444 VDD1.n164 VSUBS 0.015159f
C445 VDD1.n165 VSUBS 0.014317f
C446 VDD1.n166 VSUBS 0.026644f
C447 VDD1.n167 VSUBS 0.026644f
C448 VDD1.n168 VSUBS 0.014317f
C449 VDD1.n169 VSUBS 0.015159f
C450 VDD1.n170 VSUBS 0.03384f
C451 VDD1.n171 VSUBS 0.03384f
C452 VDD1.n172 VSUBS 0.015159f
C453 VDD1.n173 VSUBS 0.014317f
C454 VDD1.n174 VSUBS 0.026644f
C455 VDD1.n175 VSUBS 0.026644f
C456 VDD1.n176 VSUBS 0.014317f
C457 VDD1.n177 VSUBS 0.015159f
C458 VDD1.n178 VSUBS 0.03384f
C459 VDD1.n179 VSUBS 0.03384f
C460 VDD1.n180 VSUBS 0.03384f
C461 VDD1.n181 VSUBS 0.015159f
C462 VDD1.n182 VSUBS 0.014317f
C463 VDD1.n183 VSUBS 0.026644f
C464 VDD1.n184 VSUBS 0.026644f
C465 VDD1.n185 VSUBS 0.014317f
C466 VDD1.n186 VSUBS 0.014738f
C467 VDD1.n187 VSUBS 0.014738f
C468 VDD1.n188 VSUBS 0.03384f
C469 VDD1.n189 VSUBS 0.03384f
C470 VDD1.n190 VSUBS 0.015159f
C471 VDD1.n191 VSUBS 0.014317f
C472 VDD1.n192 VSUBS 0.026644f
C473 VDD1.n193 VSUBS 0.026644f
C474 VDD1.n194 VSUBS 0.014317f
C475 VDD1.n195 VSUBS 0.015159f
C476 VDD1.n196 VSUBS 0.03384f
C477 VDD1.n197 VSUBS 0.03384f
C478 VDD1.n198 VSUBS 0.015159f
C479 VDD1.n199 VSUBS 0.014317f
C480 VDD1.n200 VSUBS 0.026644f
C481 VDD1.n201 VSUBS 0.026644f
C482 VDD1.n202 VSUBS 0.014317f
C483 VDD1.n203 VSUBS 0.015159f
C484 VDD1.n204 VSUBS 0.03384f
C485 VDD1.n205 VSUBS 0.083084f
C486 VDD1.n206 VSUBS 0.015159f
C487 VDD1.n207 VSUBS 0.014317f
C488 VDD1.n208 VSUBS 0.061585f
C489 VDD1.n209 VSUBS 0.064906f
C490 VDD1.t0 VSUBS 0.399196f
C491 VDD1.t2 VSUBS 0.399196f
C492 VDD1.n210 VSUBS 3.34039f
C493 VDD1.n211 VSUBS 3.41538f
C494 VDD1.t1 VSUBS 0.399196f
C495 VDD1.t3 VSUBS 0.399196f
C496 VDD1.n212 VSUBS 3.33581f
C497 VDD1.n213 VSUBS 3.63445f
C498 VTAIL.t1 VSUBS 0.406349f
C499 VTAIL.t10 VSUBS 0.406349f
C500 VTAIL.n0 VSUBS 3.2231f
C501 VTAIL.n1 VSUBS 0.847096f
C502 VTAIL.n2 VSUBS 0.030147f
C503 VTAIL.n3 VSUBS 0.027121f
C504 VTAIL.n4 VSUBS 0.014574f
C505 VTAIL.n5 VSUBS 0.034447f
C506 VTAIL.n6 VSUBS 0.015431f
C507 VTAIL.n7 VSUBS 0.027121f
C508 VTAIL.n8 VSUBS 0.014574f
C509 VTAIL.n9 VSUBS 0.034447f
C510 VTAIL.n10 VSUBS 0.015431f
C511 VTAIL.n11 VSUBS 0.027121f
C512 VTAIL.n12 VSUBS 0.014574f
C513 VTAIL.n13 VSUBS 0.034447f
C514 VTAIL.n14 VSUBS 0.015431f
C515 VTAIL.n15 VSUBS 0.027121f
C516 VTAIL.n16 VSUBS 0.014574f
C517 VTAIL.n17 VSUBS 0.034447f
C518 VTAIL.n18 VSUBS 0.015431f
C519 VTAIL.n19 VSUBS 0.027121f
C520 VTAIL.n20 VSUBS 0.014574f
C521 VTAIL.n21 VSUBS 0.034447f
C522 VTAIL.n22 VSUBS 0.015431f
C523 VTAIL.n23 VSUBS 0.027121f
C524 VTAIL.n24 VSUBS 0.014574f
C525 VTAIL.n25 VSUBS 0.034447f
C526 VTAIL.n26 VSUBS 0.015431f
C527 VTAIL.n27 VSUBS 0.027121f
C528 VTAIL.n28 VSUBS 0.014574f
C529 VTAIL.n29 VSUBS 0.034447f
C530 VTAIL.n30 VSUBS 0.015431f
C531 VTAIL.n31 VSUBS 0.027121f
C532 VTAIL.n32 VSUBS 0.014574f
C533 VTAIL.n33 VSUBS 0.034447f
C534 VTAIL.n34 VSUBS 0.015431f
C535 VTAIL.n35 VSUBS 0.222859f
C536 VTAIL.t9 VSUBS 0.074011f
C537 VTAIL.n36 VSUBS 0.025835f
C538 VTAIL.n37 VSUBS 0.021914f
C539 VTAIL.n38 VSUBS 0.014574f
C540 VTAIL.n39 VSUBS 2.2193f
C541 VTAIL.n40 VSUBS 0.027121f
C542 VTAIL.n41 VSUBS 0.014574f
C543 VTAIL.n42 VSUBS 0.015431f
C544 VTAIL.n43 VSUBS 0.034447f
C545 VTAIL.n44 VSUBS 0.034447f
C546 VTAIL.n45 VSUBS 0.015431f
C547 VTAIL.n46 VSUBS 0.014574f
C548 VTAIL.n47 VSUBS 0.027121f
C549 VTAIL.n48 VSUBS 0.027121f
C550 VTAIL.n49 VSUBS 0.014574f
C551 VTAIL.n50 VSUBS 0.015431f
C552 VTAIL.n51 VSUBS 0.034447f
C553 VTAIL.n52 VSUBS 0.034447f
C554 VTAIL.n53 VSUBS 0.015431f
C555 VTAIL.n54 VSUBS 0.014574f
C556 VTAIL.n55 VSUBS 0.027121f
C557 VTAIL.n56 VSUBS 0.027121f
C558 VTAIL.n57 VSUBS 0.014574f
C559 VTAIL.n58 VSUBS 0.015431f
C560 VTAIL.n59 VSUBS 0.034447f
C561 VTAIL.n60 VSUBS 0.034447f
C562 VTAIL.n61 VSUBS 0.015431f
C563 VTAIL.n62 VSUBS 0.014574f
C564 VTAIL.n63 VSUBS 0.027121f
C565 VTAIL.n64 VSUBS 0.027121f
C566 VTAIL.n65 VSUBS 0.014574f
C567 VTAIL.n66 VSUBS 0.015431f
C568 VTAIL.n67 VSUBS 0.034447f
C569 VTAIL.n68 VSUBS 0.034447f
C570 VTAIL.n69 VSUBS 0.015431f
C571 VTAIL.n70 VSUBS 0.014574f
C572 VTAIL.n71 VSUBS 0.027121f
C573 VTAIL.n72 VSUBS 0.027121f
C574 VTAIL.n73 VSUBS 0.014574f
C575 VTAIL.n74 VSUBS 0.015431f
C576 VTAIL.n75 VSUBS 0.034447f
C577 VTAIL.n76 VSUBS 0.034447f
C578 VTAIL.n77 VSUBS 0.034447f
C579 VTAIL.n78 VSUBS 0.015431f
C580 VTAIL.n79 VSUBS 0.014574f
C581 VTAIL.n80 VSUBS 0.027121f
C582 VTAIL.n81 VSUBS 0.027121f
C583 VTAIL.n82 VSUBS 0.014574f
C584 VTAIL.n83 VSUBS 0.015002f
C585 VTAIL.n84 VSUBS 0.015002f
C586 VTAIL.n85 VSUBS 0.034447f
C587 VTAIL.n86 VSUBS 0.034447f
C588 VTAIL.n87 VSUBS 0.015431f
C589 VTAIL.n88 VSUBS 0.014574f
C590 VTAIL.n89 VSUBS 0.027121f
C591 VTAIL.n90 VSUBS 0.027121f
C592 VTAIL.n91 VSUBS 0.014574f
C593 VTAIL.n92 VSUBS 0.015431f
C594 VTAIL.n93 VSUBS 0.034447f
C595 VTAIL.n94 VSUBS 0.034447f
C596 VTAIL.n95 VSUBS 0.015431f
C597 VTAIL.n96 VSUBS 0.014574f
C598 VTAIL.n97 VSUBS 0.027121f
C599 VTAIL.n98 VSUBS 0.027121f
C600 VTAIL.n99 VSUBS 0.014574f
C601 VTAIL.n100 VSUBS 0.015431f
C602 VTAIL.n101 VSUBS 0.034447f
C603 VTAIL.n102 VSUBS 0.084572f
C604 VTAIL.n103 VSUBS 0.015431f
C605 VTAIL.n104 VSUBS 0.014574f
C606 VTAIL.n105 VSUBS 0.062689f
C607 VTAIL.n106 VSUBS 0.042583f
C608 VTAIL.n107 VSUBS 0.315092f
C609 VTAIL.t8 VSUBS 0.406349f
C610 VTAIL.t6 VSUBS 0.406349f
C611 VTAIL.n108 VSUBS 3.2231f
C612 VTAIL.n109 VSUBS 2.97404f
C613 VTAIL.t2 VSUBS 0.406349f
C614 VTAIL.t3 VSUBS 0.406349f
C615 VTAIL.n110 VSUBS 3.22312f
C616 VTAIL.n111 VSUBS 2.97403f
C617 VTAIL.n112 VSUBS 0.030147f
C618 VTAIL.n113 VSUBS 0.027121f
C619 VTAIL.n114 VSUBS 0.014574f
C620 VTAIL.n115 VSUBS 0.034447f
C621 VTAIL.n116 VSUBS 0.015431f
C622 VTAIL.n117 VSUBS 0.027121f
C623 VTAIL.n118 VSUBS 0.014574f
C624 VTAIL.n119 VSUBS 0.034447f
C625 VTAIL.n120 VSUBS 0.015431f
C626 VTAIL.n121 VSUBS 0.027121f
C627 VTAIL.n122 VSUBS 0.014574f
C628 VTAIL.n123 VSUBS 0.034447f
C629 VTAIL.n124 VSUBS 0.015431f
C630 VTAIL.n125 VSUBS 0.027121f
C631 VTAIL.n126 VSUBS 0.014574f
C632 VTAIL.n127 VSUBS 0.034447f
C633 VTAIL.n128 VSUBS 0.034447f
C634 VTAIL.n129 VSUBS 0.015431f
C635 VTAIL.n130 VSUBS 0.027121f
C636 VTAIL.n131 VSUBS 0.014574f
C637 VTAIL.n132 VSUBS 0.034447f
C638 VTAIL.n133 VSUBS 0.015431f
C639 VTAIL.n134 VSUBS 0.027121f
C640 VTAIL.n135 VSUBS 0.014574f
C641 VTAIL.n136 VSUBS 0.034447f
C642 VTAIL.n137 VSUBS 0.015431f
C643 VTAIL.n138 VSUBS 0.027121f
C644 VTAIL.n139 VSUBS 0.014574f
C645 VTAIL.n140 VSUBS 0.034447f
C646 VTAIL.n141 VSUBS 0.015431f
C647 VTAIL.n142 VSUBS 0.027121f
C648 VTAIL.n143 VSUBS 0.014574f
C649 VTAIL.n144 VSUBS 0.034447f
C650 VTAIL.n145 VSUBS 0.015431f
C651 VTAIL.n146 VSUBS 0.222859f
C652 VTAIL.t11 VSUBS 0.074011f
C653 VTAIL.n147 VSUBS 0.025835f
C654 VTAIL.n148 VSUBS 0.021914f
C655 VTAIL.n149 VSUBS 0.014574f
C656 VTAIL.n150 VSUBS 2.2193f
C657 VTAIL.n151 VSUBS 0.027121f
C658 VTAIL.n152 VSUBS 0.014574f
C659 VTAIL.n153 VSUBS 0.015431f
C660 VTAIL.n154 VSUBS 0.034447f
C661 VTAIL.n155 VSUBS 0.034447f
C662 VTAIL.n156 VSUBS 0.015431f
C663 VTAIL.n157 VSUBS 0.014574f
C664 VTAIL.n158 VSUBS 0.027121f
C665 VTAIL.n159 VSUBS 0.027121f
C666 VTAIL.n160 VSUBS 0.014574f
C667 VTAIL.n161 VSUBS 0.015431f
C668 VTAIL.n162 VSUBS 0.034447f
C669 VTAIL.n163 VSUBS 0.034447f
C670 VTAIL.n164 VSUBS 0.015431f
C671 VTAIL.n165 VSUBS 0.014574f
C672 VTAIL.n166 VSUBS 0.027121f
C673 VTAIL.n167 VSUBS 0.027121f
C674 VTAIL.n168 VSUBS 0.014574f
C675 VTAIL.n169 VSUBS 0.015431f
C676 VTAIL.n170 VSUBS 0.034447f
C677 VTAIL.n171 VSUBS 0.034447f
C678 VTAIL.n172 VSUBS 0.015431f
C679 VTAIL.n173 VSUBS 0.014574f
C680 VTAIL.n174 VSUBS 0.027121f
C681 VTAIL.n175 VSUBS 0.027121f
C682 VTAIL.n176 VSUBS 0.014574f
C683 VTAIL.n177 VSUBS 0.015431f
C684 VTAIL.n178 VSUBS 0.034447f
C685 VTAIL.n179 VSUBS 0.034447f
C686 VTAIL.n180 VSUBS 0.015431f
C687 VTAIL.n181 VSUBS 0.014574f
C688 VTAIL.n182 VSUBS 0.027121f
C689 VTAIL.n183 VSUBS 0.027121f
C690 VTAIL.n184 VSUBS 0.014574f
C691 VTAIL.n185 VSUBS 0.015431f
C692 VTAIL.n186 VSUBS 0.034447f
C693 VTAIL.n187 VSUBS 0.034447f
C694 VTAIL.n188 VSUBS 0.015431f
C695 VTAIL.n189 VSUBS 0.014574f
C696 VTAIL.n190 VSUBS 0.027121f
C697 VTAIL.n191 VSUBS 0.027121f
C698 VTAIL.n192 VSUBS 0.014574f
C699 VTAIL.n193 VSUBS 0.015002f
C700 VTAIL.n194 VSUBS 0.015002f
C701 VTAIL.n195 VSUBS 0.034447f
C702 VTAIL.n196 VSUBS 0.034447f
C703 VTAIL.n197 VSUBS 0.015431f
C704 VTAIL.n198 VSUBS 0.014574f
C705 VTAIL.n199 VSUBS 0.027121f
C706 VTAIL.n200 VSUBS 0.027121f
C707 VTAIL.n201 VSUBS 0.014574f
C708 VTAIL.n202 VSUBS 0.015431f
C709 VTAIL.n203 VSUBS 0.034447f
C710 VTAIL.n204 VSUBS 0.034447f
C711 VTAIL.n205 VSUBS 0.015431f
C712 VTAIL.n206 VSUBS 0.014574f
C713 VTAIL.n207 VSUBS 0.027121f
C714 VTAIL.n208 VSUBS 0.027121f
C715 VTAIL.n209 VSUBS 0.014574f
C716 VTAIL.n210 VSUBS 0.015431f
C717 VTAIL.n211 VSUBS 0.034447f
C718 VTAIL.n212 VSUBS 0.084572f
C719 VTAIL.n213 VSUBS 0.015431f
C720 VTAIL.n214 VSUBS 0.014574f
C721 VTAIL.n215 VSUBS 0.062689f
C722 VTAIL.n216 VSUBS 0.042583f
C723 VTAIL.n217 VSUBS 0.315092f
C724 VTAIL.t5 VSUBS 0.406349f
C725 VTAIL.t7 VSUBS 0.406349f
C726 VTAIL.n218 VSUBS 3.22312f
C727 VTAIL.n219 VSUBS 0.967435f
C728 VTAIL.n220 VSUBS 0.030147f
C729 VTAIL.n221 VSUBS 0.027121f
C730 VTAIL.n222 VSUBS 0.014574f
C731 VTAIL.n223 VSUBS 0.034447f
C732 VTAIL.n224 VSUBS 0.015431f
C733 VTAIL.n225 VSUBS 0.027121f
C734 VTAIL.n226 VSUBS 0.014574f
C735 VTAIL.n227 VSUBS 0.034447f
C736 VTAIL.n228 VSUBS 0.015431f
C737 VTAIL.n229 VSUBS 0.027121f
C738 VTAIL.n230 VSUBS 0.014574f
C739 VTAIL.n231 VSUBS 0.034447f
C740 VTAIL.n232 VSUBS 0.015431f
C741 VTAIL.n233 VSUBS 0.027121f
C742 VTAIL.n234 VSUBS 0.014574f
C743 VTAIL.n235 VSUBS 0.034447f
C744 VTAIL.n236 VSUBS 0.034447f
C745 VTAIL.n237 VSUBS 0.015431f
C746 VTAIL.n238 VSUBS 0.027121f
C747 VTAIL.n239 VSUBS 0.014574f
C748 VTAIL.n240 VSUBS 0.034447f
C749 VTAIL.n241 VSUBS 0.015431f
C750 VTAIL.n242 VSUBS 0.027121f
C751 VTAIL.n243 VSUBS 0.014574f
C752 VTAIL.n244 VSUBS 0.034447f
C753 VTAIL.n245 VSUBS 0.015431f
C754 VTAIL.n246 VSUBS 0.027121f
C755 VTAIL.n247 VSUBS 0.014574f
C756 VTAIL.n248 VSUBS 0.034447f
C757 VTAIL.n249 VSUBS 0.015431f
C758 VTAIL.n250 VSUBS 0.027121f
C759 VTAIL.n251 VSUBS 0.014574f
C760 VTAIL.n252 VSUBS 0.034447f
C761 VTAIL.n253 VSUBS 0.015431f
C762 VTAIL.n254 VSUBS 0.222859f
C763 VTAIL.t4 VSUBS 0.074011f
C764 VTAIL.n255 VSUBS 0.025835f
C765 VTAIL.n256 VSUBS 0.021914f
C766 VTAIL.n257 VSUBS 0.014574f
C767 VTAIL.n258 VSUBS 2.2193f
C768 VTAIL.n259 VSUBS 0.027121f
C769 VTAIL.n260 VSUBS 0.014574f
C770 VTAIL.n261 VSUBS 0.015431f
C771 VTAIL.n262 VSUBS 0.034447f
C772 VTAIL.n263 VSUBS 0.034447f
C773 VTAIL.n264 VSUBS 0.015431f
C774 VTAIL.n265 VSUBS 0.014574f
C775 VTAIL.n266 VSUBS 0.027121f
C776 VTAIL.n267 VSUBS 0.027121f
C777 VTAIL.n268 VSUBS 0.014574f
C778 VTAIL.n269 VSUBS 0.015431f
C779 VTAIL.n270 VSUBS 0.034447f
C780 VTAIL.n271 VSUBS 0.034447f
C781 VTAIL.n272 VSUBS 0.015431f
C782 VTAIL.n273 VSUBS 0.014574f
C783 VTAIL.n274 VSUBS 0.027121f
C784 VTAIL.n275 VSUBS 0.027121f
C785 VTAIL.n276 VSUBS 0.014574f
C786 VTAIL.n277 VSUBS 0.015431f
C787 VTAIL.n278 VSUBS 0.034447f
C788 VTAIL.n279 VSUBS 0.034447f
C789 VTAIL.n280 VSUBS 0.015431f
C790 VTAIL.n281 VSUBS 0.014574f
C791 VTAIL.n282 VSUBS 0.027121f
C792 VTAIL.n283 VSUBS 0.027121f
C793 VTAIL.n284 VSUBS 0.014574f
C794 VTAIL.n285 VSUBS 0.015431f
C795 VTAIL.n286 VSUBS 0.034447f
C796 VTAIL.n287 VSUBS 0.034447f
C797 VTAIL.n288 VSUBS 0.015431f
C798 VTAIL.n289 VSUBS 0.014574f
C799 VTAIL.n290 VSUBS 0.027121f
C800 VTAIL.n291 VSUBS 0.027121f
C801 VTAIL.n292 VSUBS 0.014574f
C802 VTAIL.n293 VSUBS 0.015431f
C803 VTAIL.n294 VSUBS 0.034447f
C804 VTAIL.n295 VSUBS 0.034447f
C805 VTAIL.n296 VSUBS 0.015431f
C806 VTAIL.n297 VSUBS 0.014574f
C807 VTAIL.n298 VSUBS 0.027121f
C808 VTAIL.n299 VSUBS 0.027121f
C809 VTAIL.n300 VSUBS 0.014574f
C810 VTAIL.n301 VSUBS 0.015002f
C811 VTAIL.n302 VSUBS 0.015002f
C812 VTAIL.n303 VSUBS 0.034447f
C813 VTAIL.n304 VSUBS 0.034447f
C814 VTAIL.n305 VSUBS 0.015431f
C815 VTAIL.n306 VSUBS 0.014574f
C816 VTAIL.n307 VSUBS 0.027121f
C817 VTAIL.n308 VSUBS 0.027121f
C818 VTAIL.n309 VSUBS 0.014574f
C819 VTAIL.n310 VSUBS 0.015431f
C820 VTAIL.n311 VSUBS 0.034447f
C821 VTAIL.n312 VSUBS 0.034447f
C822 VTAIL.n313 VSUBS 0.015431f
C823 VTAIL.n314 VSUBS 0.014574f
C824 VTAIL.n315 VSUBS 0.027121f
C825 VTAIL.n316 VSUBS 0.027121f
C826 VTAIL.n317 VSUBS 0.014574f
C827 VTAIL.n318 VSUBS 0.015431f
C828 VTAIL.n319 VSUBS 0.034447f
C829 VTAIL.n320 VSUBS 0.084572f
C830 VTAIL.n321 VSUBS 0.015431f
C831 VTAIL.n322 VSUBS 0.014574f
C832 VTAIL.n323 VSUBS 0.062689f
C833 VTAIL.n324 VSUBS 0.042583f
C834 VTAIL.n325 VSUBS 2.15444f
C835 VTAIL.n326 VSUBS 0.030147f
C836 VTAIL.n327 VSUBS 0.027121f
C837 VTAIL.n328 VSUBS 0.014574f
C838 VTAIL.n329 VSUBS 0.034447f
C839 VTAIL.n330 VSUBS 0.015431f
C840 VTAIL.n331 VSUBS 0.027121f
C841 VTAIL.n332 VSUBS 0.014574f
C842 VTAIL.n333 VSUBS 0.034447f
C843 VTAIL.n334 VSUBS 0.015431f
C844 VTAIL.n335 VSUBS 0.027121f
C845 VTAIL.n336 VSUBS 0.014574f
C846 VTAIL.n337 VSUBS 0.034447f
C847 VTAIL.n338 VSUBS 0.015431f
C848 VTAIL.n339 VSUBS 0.027121f
C849 VTAIL.n340 VSUBS 0.014574f
C850 VTAIL.n341 VSUBS 0.034447f
C851 VTAIL.n342 VSUBS 0.015431f
C852 VTAIL.n343 VSUBS 0.027121f
C853 VTAIL.n344 VSUBS 0.014574f
C854 VTAIL.n345 VSUBS 0.034447f
C855 VTAIL.n346 VSUBS 0.015431f
C856 VTAIL.n347 VSUBS 0.027121f
C857 VTAIL.n348 VSUBS 0.014574f
C858 VTAIL.n349 VSUBS 0.034447f
C859 VTAIL.n350 VSUBS 0.015431f
C860 VTAIL.n351 VSUBS 0.027121f
C861 VTAIL.n352 VSUBS 0.014574f
C862 VTAIL.n353 VSUBS 0.034447f
C863 VTAIL.n354 VSUBS 0.015431f
C864 VTAIL.n355 VSUBS 0.027121f
C865 VTAIL.n356 VSUBS 0.014574f
C866 VTAIL.n357 VSUBS 0.034447f
C867 VTAIL.n358 VSUBS 0.015431f
C868 VTAIL.n359 VSUBS 0.222859f
C869 VTAIL.t0 VSUBS 0.074011f
C870 VTAIL.n360 VSUBS 0.025835f
C871 VTAIL.n361 VSUBS 0.021914f
C872 VTAIL.n362 VSUBS 0.014574f
C873 VTAIL.n363 VSUBS 2.2193f
C874 VTAIL.n364 VSUBS 0.027121f
C875 VTAIL.n365 VSUBS 0.014574f
C876 VTAIL.n366 VSUBS 0.015431f
C877 VTAIL.n367 VSUBS 0.034447f
C878 VTAIL.n368 VSUBS 0.034447f
C879 VTAIL.n369 VSUBS 0.015431f
C880 VTAIL.n370 VSUBS 0.014574f
C881 VTAIL.n371 VSUBS 0.027121f
C882 VTAIL.n372 VSUBS 0.027121f
C883 VTAIL.n373 VSUBS 0.014574f
C884 VTAIL.n374 VSUBS 0.015431f
C885 VTAIL.n375 VSUBS 0.034447f
C886 VTAIL.n376 VSUBS 0.034447f
C887 VTAIL.n377 VSUBS 0.015431f
C888 VTAIL.n378 VSUBS 0.014574f
C889 VTAIL.n379 VSUBS 0.027121f
C890 VTAIL.n380 VSUBS 0.027121f
C891 VTAIL.n381 VSUBS 0.014574f
C892 VTAIL.n382 VSUBS 0.015431f
C893 VTAIL.n383 VSUBS 0.034447f
C894 VTAIL.n384 VSUBS 0.034447f
C895 VTAIL.n385 VSUBS 0.015431f
C896 VTAIL.n386 VSUBS 0.014574f
C897 VTAIL.n387 VSUBS 0.027121f
C898 VTAIL.n388 VSUBS 0.027121f
C899 VTAIL.n389 VSUBS 0.014574f
C900 VTAIL.n390 VSUBS 0.015431f
C901 VTAIL.n391 VSUBS 0.034447f
C902 VTAIL.n392 VSUBS 0.034447f
C903 VTAIL.n393 VSUBS 0.015431f
C904 VTAIL.n394 VSUBS 0.014574f
C905 VTAIL.n395 VSUBS 0.027121f
C906 VTAIL.n396 VSUBS 0.027121f
C907 VTAIL.n397 VSUBS 0.014574f
C908 VTAIL.n398 VSUBS 0.015431f
C909 VTAIL.n399 VSUBS 0.034447f
C910 VTAIL.n400 VSUBS 0.034447f
C911 VTAIL.n401 VSUBS 0.034447f
C912 VTAIL.n402 VSUBS 0.015431f
C913 VTAIL.n403 VSUBS 0.014574f
C914 VTAIL.n404 VSUBS 0.027121f
C915 VTAIL.n405 VSUBS 0.027121f
C916 VTAIL.n406 VSUBS 0.014574f
C917 VTAIL.n407 VSUBS 0.015002f
C918 VTAIL.n408 VSUBS 0.015002f
C919 VTAIL.n409 VSUBS 0.034447f
C920 VTAIL.n410 VSUBS 0.034447f
C921 VTAIL.n411 VSUBS 0.015431f
C922 VTAIL.n412 VSUBS 0.014574f
C923 VTAIL.n413 VSUBS 0.027121f
C924 VTAIL.n414 VSUBS 0.027121f
C925 VTAIL.n415 VSUBS 0.014574f
C926 VTAIL.n416 VSUBS 0.015431f
C927 VTAIL.n417 VSUBS 0.034447f
C928 VTAIL.n418 VSUBS 0.034447f
C929 VTAIL.n419 VSUBS 0.015431f
C930 VTAIL.n420 VSUBS 0.014574f
C931 VTAIL.n421 VSUBS 0.027121f
C932 VTAIL.n422 VSUBS 0.027121f
C933 VTAIL.n423 VSUBS 0.014574f
C934 VTAIL.n424 VSUBS 0.015431f
C935 VTAIL.n425 VSUBS 0.034447f
C936 VTAIL.n426 VSUBS 0.084572f
C937 VTAIL.n427 VSUBS 0.015431f
C938 VTAIL.n428 VSUBS 0.014574f
C939 VTAIL.n429 VSUBS 0.062689f
C940 VTAIL.n430 VSUBS 0.042583f
C941 VTAIL.n431 VSUBS 2.10755f
C942 VP.n0 VSUBS 0.043824f
C943 VP.t3 VSUBS 3.27963f
C944 VP.n1 VSUBS 0.05799f
C945 VP.n2 VSUBS 0.033242f
C946 VP.t5 VSUBS 3.27963f
C947 VP.n3 VSUBS 0.036199f
C948 VP.n4 VSUBS 0.043824f
C949 VP.t2 VSUBS 3.27963f
C950 VP.n5 VSUBS 0.05799f
C951 VP.t1 VSUBS 3.4283f
C952 VP.n6 VSUBS 1.22999f
C953 VP.t4 VSUBS 3.27963f
C954 VP.n7 VSUBS 1.21931f
C955 VP.n8 VSUBS 0.046428f
C956 VP.n9 VSUBS 0.245546f
C957 VP.n10 VSUBS 0.033242f
C958 VP.n11 VSUBS 0.033242f
C959 VP.n12 VSUBS 0.036199f
C960 VP.n13 VSUBS 0.062274f
C961 VP.n14 VSUBS 1.24541f
C962 VP.n15 VSUBS 1.89727f
C963 VP.n16 VSUBS 1.92067f
C964 VP.t0 VSUBS 3.27963f
C965 VP.n17 VSUBS 1.24541f
C966 VP.n18 VSUBS 0.062274f
C967 VP.n19 VSUBS 0.043824f
C968 VP.n20 VSUBS 0.033242f
C969 VP.n21 VSUBS 0.033242f
C970 VP.n22 VSUBS 0.05799f
C971 VP.n23 VSUBS 0.046428f
C972 VP.n24 VSUBS 1.14321f
C973 VP.n25 VSUBS 0.046428f
C974 VP.n26 VSUBS 0.033242f
C975 VP.n27 VSUBS 0.033242f
C976 VP.n28 VSUBS 0.033242f
C977 VP.n29 VSUBS 0.036199f
C978 VP.n30 VSUBS 0.062274f
C979 VP.n31 VSUBS 1.24541f
C980 VP.n32 VSUBS 0.036632f
C981 B.n0 VSUBS 0.004791f
C982 B.n1 VSUBS 0.004791f
C983 B.n2 VSUBS 0.007576f
C984 B.n3 VSUBS 0.007576f
C985 B.n4 VSUBS 0.007576f
C986 B.n5 VSUBS 0.007576f
C987 B.n6 VSUBS 0.007576f
C988 B.n7 VSUBS 0.007576f
C989 B.n8 VSUBS 0.007576f
C990 B.n9 VSUBS 0.007576f
C991 B.n10 VSUBS 0.007576f
C992 B.n11 VSUBS 0.007576f
C993 B.n12 VSUBS 0.007576f
C994 B.n13 VSUBS 0.007576f
C995 B.n14 VSUBS 0.007576f
C996 B.n15 VSUBS 0.007576f
C997 B.n16 VSUBS 0.007576f
C998 B.n17 VSUBS 0.007576f
C999 B.n18 VSUBS 0.007576f
C1000 B.n19 VSUBS 0.018719f
C1001 B.n20 VSUBS 0.007576f
C1002 B.n21 VSUBS 0.007576f
C1003 B.n22 VSUBS 0.007576f
C1004 B.n23 VSUBS 0.007576f
C1005 B.n24 VSUBS 0.007576f
C1006 B.n25 VSUBS 0.007576f
C1007 B.n26 VSUBS 0.007576f
C1008 B.n27 VSUBS 0.007576f
C1009 B.n28 VSUBS 0.007576f
C1010 B.n29 VSUBS 0.007576f
C1011 B.n30 VSUBS 0.007576f
C1012 B.n31 VSUBS 0.007576f
C1013 B.n32 VSUBS 0.007576f
C1014 B.n33 VSUBS 0.007576f
C1015 B.n34 VSUBS 0.007576f
C1016 B.n35 VSUBS 0.007576f
C1017 B.n36 VSUBS 0.007576f
C1018 B.n37 VSUBS 0.007576f
C1019 B.n38 VSUBS 0.007576f
C1020 B.n39 VSUBS 0.007576f
C1021 B.n40 VSUBS 0.007576f
C1022 B.n41 VSUBS 0.007576f
C1023 B.n42 VSUBS 0.007576f
C1024 B.n43 VSUBS 0.007576f
C1025 B.n44 VSUBS 0.007576f
C1026 B.n45 VSUBS 0.007576f
C1027 B.n46 VSUBS 0.007576f
C1028 B.n47 VSUBS 0.007576f
C1029 B.n48 VSUBS 0.007576f
C1030 B.n49 VSUBS 0.007576f
C1031 B.t11 VSUBS 0.405356f
C1032 B.t10 VSUBS 0.433364f
C1033 B.t9 VSUBS 1.67305f
C1034 B.n50 VSUBS 0.626368f
C1035 B.n51 VSUBS 0.364794f
C1036 B.n52 VSUBS 0.017554f
C1037 B.n53 VSUBS 0.007576f
C1038 B.n54 VSUBS 0.007576f
C1039 B.n55 VSUBS 0.007576f
C1040 B.n56 VSUBS 0.007576f
C1041 B.n57 VSUBS 0.007576f
C1042 B.t2 VSUBS 0.40536f
C1043 B.t1 VSUBS 0.433367f
C1044 B.t0 VSUBS 1.67305f
C1045 B.n58 VSUBS 0.626364f
C1046 B.n59 VSUBS 0.36479f
C1047 B.n60 VSUBS 0.007576f
C1048 B.n61 VSUBS 0.007576f
C1049 B.n62 VSUBS 0.007576f
C1050 B.n63 VSUBS 0.007576f
C1051 B.n64 VSUBS 0.007576f
C1052 B.n65 VSUBS 0.007576f
C1053 B.n66 VSUBS 0.007576f
C1054 B.n67 VSUBS 0.007576f
C1055 B.n68 VSUBS 0.007576f
C1056 B.n69 VSUBS 0.007576f
C1057 B.n70 VSUBS 0.007576f
C1058 B.n71 VSUBS 0.007576f
C1059 B.n72 VSUBS 0.007576f
C1060 B.n73 VSUBS 0.007576f
C1061 B.n74 VSUBS 0.007576f
C1062 B.n75 VSUBS 0.007576f
C1063 B.n76 VSUBS 0.007576f
C1064 B.n77 VSUBS 0.007576f
C1065 B.n78 VSUBS 0.007576f
C1066 B.n79 VSUBS 0.007576f
C1067 B.n80 VSUBS 0.007576f
C1068 B.n81 VSUBS 0.007576f
C1069 B.n82 VSUBS 0.007576f
C1070 B.n83 VSUBS 0.007576f
C1071 B.n84 VSUBS 0.007576f
C1072 B.n85 VSUBS 0.007576f
C1073 B.n86 VSUBS 0.007576f
C1074 B.n87 VSUBS 0.007576f
C1075 B.n88 VSUBS 0.007576f
C1076 B.n89 VSUBS 0.007576f
C1077 B.n90 VSUBS 0.017848f
C1078 B.n91 VSUBS 0.007576f
C1079 B.n92 VSUBS 0.007576f
C1080 B.n93 VSUBS 0.007576f
C1081 B.n94 VSUBS 0.007576f
C1082 B.n95 VSUBS 0.007576f
C1083 B.n96 VSUBS 0.007576f
C1084 B.n97 VSUBS 0.007576f
C1085 B.n98 VSUBS 0.007576f
C1086 B.n99 VSUBS 0.007576f
C1087 B.n100 VSUBS 0.007576f
C1088 B.n101 VSUBS 0.007576f
C1089 B.n102 VSUBS 0.007576f
C1090 B.n103 VSUBS 0.007576f
C1091 B.n104 VSUBS 0.007576f
C1092 B.n105 VSUBS 0.007576f
C1093 B.n106 VSUBS 0.007576f
C1094 B.n107 VSUBS 0.007576f
C1095 B.n108 VSUBS 0.007576f
C1096 B.n109 VSUBS 0.007576f
C1097 B.n110 VSUBS 0.007576f
C1098 B.n111 VSUBS 0.007576f
C1099 B.n112 VSUBS 0.007576f
C1100 B.n113 VSUBS 0.007576f
C1101 B.n114 VSUBS 0.007576f
C1102 B.n115 VSUBS 0.007576f
C1103 B.n116 VSUBS 0.007576f
C1104 B.n117 VSUBS 0.007576f
C1105 B.n118 VSUBS 0.007576f
C1106 B.n119 VSUBS 0.007576f
C1107 B.n120 VSUBS 0.007576f
C1108 B.n121 VSUBS 0.007576f
C1109 B.n122 VSUBS 0.007576f
C1110 B.n123 VSUBS 0.007576f
C1111 B.n124 VSUBS 0.007576f
C1112 B.n125 VSUBS 0.018719f
C1113 B.n126 VSUBS 0.007576f
C1114 B.n127 VSUBS 0.007576f
C1115 B.n128 VSUBS 0.007576f
C1116 B.n129 VSUBS 0.007576f
C1117 B.n130 VSUBS 0.007576f
C1118 B.n131 VSUBS 0.007576f
C1119 B.n132 VSUBS 0.007576f
C1120 B.n133 VSUBS 0.007576f
C1121 B.n134 VSUBS 0.007576f
C1122 B.n135 VSUBS 0.007576f
C1123 B.n136 VSUBS 0.007576f
C1124 B.n137 VSUBS 0.007576f
C1125 B.n138 VSUBS 0.007576f
C1126 B.n139 VSUBS 0.007576f
C1127 B.n140 VSUBS 0.007576f
C1128 B.n141 VSUBS 0.007576f
C1129 B.n142 VSUBS 0.007576f
C1130 B.n143 VSUBS 0.007576f
C1131 B.n144 VSUBS 0.007576f
C1132 B.n145 VSUBS 0.007576f
C1133 B.n146 VSUBS 0.007576f
C1134 B.n147 VSUBS 0.007576f
C1135 B.n148 VSUBS 0.007576f
C1136 B.n149 VSUBS 0.007576f
C1137 B.n150 VSUBS 0.007576f
C1138 B.n151 VSUBS 0.007576f
C1139 B.n152 VSUBS 0.007576f
C1140 B.n153 VSUBS 0.007576f
C1141 B.n154 VSUBS 0.007576f
C1142 B.n155 VSUBS 0.007576f
C1143 B.t7 VSUBS 0.40536f
C1144 B.t8 VSUBS 0.433367f
C1145 B.t6 VSUBS 1.67305f
C1146 B.n156 VSUBS 0.626364f
C1147 B.n157 VSUBS 0.36479f
C1148 B.n158 VSUBS 0.017554f
C1149 B.n159 VSUBS 0.007576f
C1150 B.n160 VSUBS 0.007576f
C1151 B.n161 VSUBS 0.007576f
C1152 B.n162 VSUBS 0.007576f
C1153 B.n163 VSUBS 0.007576f
C1154 B.t4 VSUBS 0.405356f
C1155 B.t5 VSUBS 0.433364f
C1156 B.t3 VSUBS 1.67305f
C1157 B.n164 VSUBS 0.626368f
C1158 B.n165 VSUBS 0.364794f
C1159 B.n166 VSUBS 0.007576f
C1160 B.n167 VSUBS 0.007576f
C1161 B.n168 VSUBS 0.007576f
C1162 B.n169 VSUBS 0.007576f
C1163 B.n170 VSUBS 0.007576f
C1164 B.n171 VSUBS 0.007576f
C1165 B.n172 VSUBS 0.007576f
C1166 B.n173 VSUBS 0.007576f
C1167 B.n174 VSUBS 0.007576f
C1168 B.n175 VSUBS 0.007576f
C1169 B.n176 VSUBS 0.007576f
C1170 B.n177 VSUBS 0.007576f
C1171 B.n178 VSUBS 0.007576f
C1172 B.n179 VSUBS 0.007576f
C1173 B.n180 VSUBS 0.007576f
C1174 B.n181 VSUBS 0.007576f
C1175 B.n182 VSUBS 0.007576f
C1176 B.n183 VSUBS 0.007576f
C1177 B.n184 VSUBS 0.007576f
C1178 B.n185 VSUBS 0.007576f
C1179 B.n186 VSUBS 0.007576f
C1180 B.n187 VSUBS 0.007576f
C1181 B.n188 VSUBS 0.007576f
C1182 B.n189 VSUBS 0.007576f
C1183 B.n190 VSUBS 0.007576f
C1184 B.n191 VSUBS 0.007576f
C1185 B.n192 VSUBS 0.007576f
C1186 B.n193 VSUBS 0.007576f
C1187 B.n194 VSUBS 0.007576f
C1188 B.n195 VSUBS 0.007576f
C1189 B.n196 VSUBS 0.018719f
C1190 B.n197 VSUBS 0.007576f
C1191 B.n198 VSUBS 0.007576f
C1192 B.n199 VSUBS 0.007576f
C1193 B.n200 VSUBS 0.007576f
C1194 B.n201 VSUBS 0.007576f
C1195 B.n202 VSUBS 0.007576f
C1196 B.n203 VSUBS 0.007576f
C1197 B.n204 VSUBS 0.007576f
C1198 B.n205 VSUBS 0.007576f
C1199 B.n206 VSUBS 0.007576f
C1200 B.n207 VSUBS 0.007576f
C1201 B.n208 VSUBS 0.007576f
C1202 B.n209 VSUBS 0.007576f
C1203 B.n210 VSUBS 0.007576f
C1204 B.n211 VSUBS 0.007576f
C1205 B.n212 VSUBS 0.007576f
C1206 B.n213 VSUBS 0.007576f
C1207 B.n214 VSUBS 0.007576f
C1208 B.n215 VSUBS 0.007576f
C1209 B.n216 VSUBS 0.007576f
C1210 B.n217 VSUBS 0.007576f
C1211 B.n218 VSUBS 0.007576f
C1212 B.n219 VSUBS 0.007576f
C1213 B.n220 VSUBS 0.007576f
C1214 B.n221 VSUBS 0.007576f
C1215 B.n222 VSUBS 0.007576f
C1216 B.n223 VSUBS 0.007576f
C1217 B.n224 VSUBS 0.007576f
C1218 B.n225 VSUBS 0.007576f
C1219 B.n226 VSUBS 0.007576f
C1220 B.n227 VSUBS 0.007576f
C1221 B.n228 VSUBS 0.007576f
C1222 B.n229 VSUBS 0.007576f
C1223 B.n230 VSUBS 0.007576f
C1224 B.n231 VSUBS 0.007576f
C1225 B.n232 VSUBS 0.007576f
C1226 B.n233 VSUBS 0.007576f
C1227 B.n234 VSUBS 0.007576f
C1228 B.n235 VSUBS 0.007576f
C1229 B.n236 VSUBS 0.007576f
C1230 B.n237 VSUBS 0.007576f
C1231 B.n238 VSUBS 0.007576f
C1232 B.n239 VSUBS 0.007576f
C1233 B.n240 VSUBS 0.007576f
C1234 B.n241 VSUBS 0.007576f
C1235 B.n242 VSUBS 0.007576f
C1236 B.n243 VSUBS 0.007576f
C1237 B.n244 VSUBS 0.007576f
C1238 B.n245 VSUBS 0.007576f
C1239 B.n246 VSUBS 0.007576f
C1240 B.n247 VSUBS 0.007576f
C1241 B.n248 VSUBS 0.007576f
C1242 B.n249 VSUBS 0.007576f
C1243 B.n250 VSUBS 0.007576f
C1244 B.n251 VSUBS 0.007576f
C1245 B.n252 VSUBS 0.007576f
C1246 B.n253 VSUBS 0.007576f
C1247 B.n254 VSUBS 0.007576f
C1248 B.n255 VSUBS 0.007576f
C1249 B.n256 VSUBS 0.007576f
C1250 B.n257 VSUBS 0.007576f
C1251 B.n258 VSUBS 0.007576f
C1252 B.n259 VSUBS 0.007576f
C1253 B.n260 VSUBS 0.007576f
C1254 B.n261 VSUBS 0.01738f
C1255 B.n262 VSUBS 0.01738f
C1256 B.n263 VSUBS 0.018719f
C1257 B.n264 VSUBS 0.007576f
C1258 B.n265 VSUBS 0.007576f
C1259 B.n266 VSUBS 0.007576f
C1260 B.n267 VSUBS 0.007576f
C1261 B.n268 VSUBS 0.007576f
C1262 B.n269 VSUBS 0.007576f
C1263 B.n270 VSUBS 0.007576f
C1264 B.n271 VSUBS 0.007576f
C1265 B.n272 VSUBS 0.007576f
C1266 B.n273 VSUBS 0.007576f
C1267 B.n274 VSUBS 0.007576f
C1268 B.n275 VSUBS 0.007576f
C1269 B.n276 VSUBS 0.007576f
C1270 B.n277 VSUBS 0.007576f
C1271 B.n278 VSUBS 0.007576f
C1272 B.n279 VSUBS 0.007576f
C1273 B.n280 VSUBS 0.007576f
C1274 B.n281 VSUBS 0.007576f
C1275 B.n282 VSUBS 0.007576f
C1276 B.n283 VSUBS 0.007576f
C1277 B.n284 VSUBS 0.007576f
C1278 B.n285 VSUBS 0.007576f
C1279 B.n286 VSUBS 0.007576f
C1280 B.n287 VSUBS 0.007576f
C1281 B.n288 VSUBS 0.007576f
C1282 B.n289 VSUBS 0.007576f
C1283 B.n290 VSUBS 0.007576f
C1284 B.n291 VSUBS 0.007576f
C1285 B.n292 VSUBS 0.007576f
C1286 B.n293 VSUBS 0.007576f
C1287 B.n294 VSUBS 0.007576f
C1288 B.n295 VSUBS 0.007576f
C1289 B.n296 VSUBS 0.007576f
C1290 B.n297 VSUBS 0.007576f
C1291 B.n298 VSUBS 0.007576f
C1292 B.n299 VSUBS 0.007576f
C1293 B.n300 VSUBS 0.007576f
C1294 B.n301 VSUBS 0.007576f
C1295 B.n302 VSUBS 0.007576f
C1296 B.n303 VSUBS 0.007576f
C1297 B.n304 VSUBS 0.007576f
C1298 B.n305 VSUBS 0.007576f
C1299 B.n306 VSUBS 0.007576f
C1300 B.n307 VSUBS 0.007576f
C1301 B.n308 VSUBS 0.007576f
C1302 B.n309 VSUBS 0.007576f
C1303 B.n310 VSUBS 0.007576f
C1304 B.n311 VSUBS 0.007576f
C1305 B.n312 VSUBS 0.007576f
C1306 B.n313 VSUBS 0.007576f
C1307 B.n314 VSUBS 0.007576f
C1308 B.n315 VSUBS 0.007576f
C1309 B.n316 VSUBS 0.007576f
C1310 B.n317 VSUBS 0.007576f
C1311 B.n318 VSUBS 0.007576f
C1312 B.n319 VSUBS 0.007576f
C1313 B.n320 VSUBS 0.007576f
C1314 B.n321 VSUBS 0.007576f
C1315 B.n322 VSUBS 0.007576f
C1316 B.n323 VSUBS 0.007576f
C1317 B.n324 VSUBS 0.007576f
C1318 B.n325 VSUBS 0.007576f
C1319 B.n326 VSUBS 0.007576f
C1320 B.n327 VSUBS 0.007576f
C1321 B.n328 VSUBS 0.007576f
C1322 B.n329 VSUBS 0.007576f
C1323 B.n330 VSUBS 0.007576f
C1324 B.n331 VSUBS 0.007576f
C1325 B.n332 VSUBS 0.007576f
C1326 B.n333 VSUBS 0.007576f
C1327 B.n334 VSUBS 0.007576f
C1328 B.n335 VSUBS 0.007576f
C1329 B.n336 VSUBS 0.007576f
C1330 B.n337 VSUBS 0.007576f
C1331 B.n338 VSUBS 0.007576f
C1332 B.n339 VSUBS 0.007576f
C1333 B.n340 VSUBS 0.007576f
C1334 B.n341 VSUBS 0.007576f
C1335 B.n342 VSUBS 0.007576f
C1336 B.n343 VSUBS 0.007576f
C1337 B.n344 VSUBS 0.007576f
C1338 B.n345 VSUBS 0.007576f
C1339 B.n346 VSUBS 0.007576f
C1340 B.n347 VSUBS 0.007576f
C1341 B.n348 VSUBS 0.007576f
C1342 B.n349 VSUBS 0.007576f
C1343 B.n350 VSUBS 0.007576f
C1344 B.n351 VSUBS 0.007576f
C1345 B.n352 VSUBS 0.007576f
C1346 B.n353 VSUBS 0.007576f
C1347 B.n354 VSUBS 0.007576f
C1348 B.n355 VSUBS 0.007131f
C1349 B.n356 VSUBS 0.017554f
C1350 B.n357 VSUBS 0.004234f
C1351 B.n358 VSUBS 0.007576f
C1352 B.n359 VSUBS 0.007576f
C1353 B.n360 VSUBS 0.007576f
C1354 B.n361 VSUBS 0.007576f
C1355 B.n362 VSUBS 0.007576f
C1356 B.n363 VSUBS 0.007576f
C1357 B.n364 VSUBS 0.007576f
C1358 B.n365 VSUBS 0.007576f
C1359 B.n366 VSUBS 0.007576f
C1360 B.n367 VSUBS 0.007576f
C1361 B.n368 VSUBS 0.007576f
C1362 B.n369 VSUBS 0.007576f
C1363 B.n370 VSUBS 0.004234f
C1364 B.n371 VSUBS 0.007576f
C1365 B.n372 VSUBS 0.007576f
C1366 B.n373 VSUBS 0.007131f
C1367 B.n374 VSUBS 0.007576f
C1368 B.n375 VSUBS 0.007576f
C1369 B.n376 VSUBS 0.007576f
C1370 B.n377 VSUBS 0.007576f
C1371 B.n378 VSUBS 0.007576f
C1372 B.n379 VSUBS 0.007576f
C1373 B.n380 VSUBS 0.007576f
C1374 B.n381 VSUBS 0.007576f
C1375 B.n382 VSUBS 0.007576f
C1376 B.n383 VSUBS 0.007576f
C1377 B.n384 VSUBS 0.007576f
C1378 B.n385 VSUBS 0.007576f
C1379 B.n386 VSUBS 0.007576f
C1380 B.n387 VSUBS 0.007576f
C1381 B.n388 VSUBS 0.007576f
C1382 B.n389 VSUBS 0.007576f
C1383 B.n390 VSUBS 0.007576f
C1384 B.n391 VSUBS 0.007576f
C1385 B.n392 VSUBS 0.007576f
C1386 B.n393 VSUBS 0.007576f
C1387 B.n394 VSUBS 0.007576f
C1388 B.n395 VSUBS 0.007576f
C1389 B.n396 VSUBS 0.007576f
C1390 B.n397 VSUBS 0.007576f
C1391 B.n398 VSUBS 0.007576f
C1392 B.n399 VSUBS 0.007576f
C1393 B.n400 VSUBS 0.007576f
C1394 B.n401 VSUBS 0.007576f
C1395 B.n402 VSUBS 0.007576f
C1396 B.n403 VSUBS 0.007576f
C1397 B.n404 VSUBS 0.007576f
C1398 B.n405 VSUBS 0.007576f
C1399 B.n406 VSUBS 0.007576f
C1400 B.n407 VSUBS 0.007576f
C1401 B.n408 VSUBS 0.007576f
C1402 B.n409 VSUBS 0.007576f
C1403 B.n410 VSUBS 0.007576f
C1404 B.n411 VSUBS 0.007576f
C1405 B.n412 VSUBS 0.007576f
C1406 B.n413 VSUBS 0.007576f
C1407 B.n414 VSUBS 0.007576f
C1408 B.n415 VSUBS 0.007576f
C1409 B.n416 VSUBS 0.007576f
C1410 B.n417 VSUBS 0.007576f
C1411 B.n418 VSUBS 0.007576f
C1412 B.n419 VSUBS 0.007576f
C1413 B.n420 VSUBS 0.007576f
C1414 B.n421 VSUBS 0.007576f
C1415 B.n422 VSUBS 0.007576f
C1416 B.n423 VSUBS 0.007576f
C1417 B.n424 VSUBS 0.007576f
C1418 B.n425 VSUBS 0.007576f
C1419 B.n426 VSUBS 0.007576f
C1420 B.n427 VSUBS 0.007576f
C1421 B.n428 VSUBS 0.007576f
C1422 B.n429 VSUBS 0.007576f
C1423 B.n430 VSUBS 0.007576f
C1424 B.n431 VSUBS 0.007576f
C1425 B.n432 VSUBS 0.007576f
C1426 B.n433 VSUBS 0.007576f
C1427 B.n434 VSUBS 0.007576f
C1428 B.n435 VSUBS 0.007576f
C1429 B.n436 VSUBS 0.007576f
C1430 B.n437 VSUBS 0.007576f
C1431 B.n438 VSUBS 0.007576f
C1432 B.n439 VSUBS 0.007576f
C1433 B.n440 VSUBS 0.007576f
C1434 B.n441 VSUBS 0.007576f
C1435 B.n442 VSUBS 0.007576f
C1436 B.n443 VSUBS 0.007576f
C1437 B.n444 VSUBS 0.007576f
C1438 B.n445 VSUBS 0.007576f
C1439 B.n446 VSUBS 0.007576f
C1440 B.n447 VSUBS 0.007576f
C1441 B.n448 VSUBS 0.007576f
C1442 B.n449 VSUBS 0.007576f
C1443 B.n450 VSUBS 0.007576f
C1444 B.n451 VSUBS 0.007576f
C1445 B.n452 VSUBS 0.007576f
C1446 B.n453 VSUBS 0.007576f
C1447 B.n454 VSUBS 0.007576f
C1448 B.n455 VSUBS 0.007576f
C1449 B.n456 VSUBS 0.007576f
C1450 B.n457 VSUBS 0.007576f
C1451 B.n458 VSUBS 0.007576f
C1452 B.n459 VSUBS 0.007576f
C1453 B.n460 VSUBS 0.007576f
C1454 B.n461 VSUBS 0.007576f
C1455 B.n462 VSUBS 0.007576f
C1456 B.n463 VSUBS 0.007576f
C1457 B.n464 VSUBS 0.018719f
C1458 B.n465 VSUBS 0.01738f
C1459 B.n466 VSUBS 0.01738f
C1460 B.n467 VSUBS 0.007576f
C1461 B.n468 VSUBS 0.007576f
C1462 B.n469 VSUBS 0.007576f
C1463 B.n470 VSUBS 0.007576f
C1464 B.n471 VSUBS 0.007576f
C1465 B.n472 VSUBS 0.007576f
C1466 B.n473 VSUBS 0.007576f
C1467 B.n474 VSUBS 0.007576f
C1468 B.n475 VSUBS 0.007576f
C1469 B.n476 VSUBS 0.007576f
C1470 B.n477 VSUBS 0.007576f
C1471 B.n478 VSUBS 0.007576f
C1472 B.n479 VSUBS 0.007576f
C1473 B.n480 VSUBS 0.007576f
C1474 B.n481 VSUBS 0.007576f
C1475 B.n482 VSUBS 0.007576f
C1476 B.n483 VSUBS 0.007576f
C1477 B.n484 VSUBS 0.007576f
C1478 B.n485 VSUBS 0.007576f
C1479 B.n486 VSUBS 0.007576f
C1480 B.n487 VSUBS 0.007576f
C1481 B.n488 VSUBS 0.007576f
C1482 B.n489 VSUBS 0.007576f
C1483 B.n490 VSUBS 0.007576f
C1484 B.n491 VSUBS 0.007576f
C1485 B.n492 VSUBS 0.007576f
C1486 B.n493 VSUBS 0.007576f
C1487 B.n494 VSUBS 0.007576f
C1488 B.n495 VSUBS 0.007576f
C1489 B.n496 VSUBS 0.007576f
C1490 B.n497 VSUBS 0.007576f
C1491 B.n498 VSUBS 0.007576f
C1492 B.n499 VSUBS 0.007576f
C1493 B.n500 VSUBS 0.007576f
C1494 B.n501 VSUBS 0.007576f
C1495 B.n502 VSUBS 0.007576f
C1496 B.n503 VSUBS 0.007576f
C1497 B.n504 VSUBS 0.007576f
C1498 B.n505 VSUBS 0.007576f
C1499 B.n506 VSUBS 0.007576f
C1500 B.n507 VSUBS 0.007576f
C1501 B.n508 VSUBS 0.007576f
C1502 B.n509 VSUBS 0.007576f
C1503 B.n510 VSUBS 0.007576f
C1504 B.n511 VSUBS 0.007576f
C1505 B.n512 VSUBS 0.007576f
C1506 B.n513 VSUBS 0.007576f
C1507 B.n514 VSUBS 0.007576f
C1508 B.n515 VSUBS 0.007576f
C1509 B.n516 VSUBS 0.007576f
C1510 B.n517 VSUBS 0.007576f
C1511 B.n518 VSUBS 0.007576f
C1512 B.n519 VSUBS 0.007576f
C1513 B.n520 VSUBS 0.007576f
C1514 B.n521 VSUBS 0.007576f
C1515 B.n522 VSUBS 0.007576f
C1516 B.n523 VSUBS 0.007576f
C1517 B.n524 VSUBS 0.007576f
C1518 B.n525 VSUBS 0.007576f
C1519 B.n526 VSUBS 0.007576f
C1520 B.n527 VSUBS 0.007576f
C1521 B.n528 VSUBS 0.007576f
C1522 B.n529 VSUBS 0.007576f
C1523 B.n530 VSUBS 0.007576f
C1524 B.n531 VSUBS 0.007576f
C1525 B.n532 VSUBS 0.007576f
C1526 B.n533 VSUBS 0.007576f
C1527 B.n534 VSUBS 0.007576f
C1528 B.n535 VSUBS 0.007576f
C1529 B.n536 VSUBS 0.007576f
C1530 B.n537 VSUBS 0.007576f
C1531 B.n538 VSUBS 0.007576f
C1532 B.n539 VSUBS 0.007576f
C1533 B.n540 VSUBS 0.007576f
C1534 B.n541 VSUBS 0.007576f
C1535 B.n542 VSUBS 0.007576f
C1536 B.n543 VSUBS 0.007576f
C1537 B.n544 VSUBS 0.007576f
C1538 B.n545 VSUBS 0.007576f
C1539 B.n546 VSUBS 0.007576f
C1540 B.n547 VSUBS 0.007576f
C1541 B.n548 VSUBS 0.007576f
C1542 B.n549 VSUBS 0.007576f
C1543 B.n550 VSUBS 0.007576f
C1544 B.n551 VSUBS 0.007576f
C1545 B.n552 VSUBS 0.007576f
C1546 B.n553 VSUBS 0.007576f
C1547 B.n554 VSUBS 0.007576f
C1548 B.n555 VSUBS 0.007576f
C1549 B.n556 VSUBS 0.007576f
C1550 B.n557 VSUBS 0.007576f
C1551 B.n558 VSUBS 0.007576f
C1552 B.n559 VSUBS 0.007576f
C1553 B.n560 VSUBS 0.007576f
C1554 B.n561 VSUBS 0.007576f
C1555 B.n562 VSUBS 0.007576f
C1556 B.n563 VSUBS 0.007576f
C1557 B.n564 VSUBS 0.007576f
C1558 B.n565 VSUBS 0.007576f
C1559 B.n566 VSUBS 0.007576f
C1560 B.n567 VSUBS 0.018252f
C1561 B.n568 VSUBS 0.01738f
C1562 B.n569 VSUBS 0.018719f
C1563 B.n570 VSUBS 0.007576f
C1564 B.n571 VSUBS 0.007576f
C1565 B.n572 VSUBS 0.007576f
C1566 B.n573 VSUBS 0.007576f
C1567 B.n574 VSUBS 0.007576f
C1568 B.n575 VSUBS 0.007576f
C1569 B.n576 VSUBS 0.007576f
C1570 B.n577 VSUBS 0.007576f
C1571 B.n578 VSUBS 0.007576f
C1572 B.n579 VSUBS 0.007576f
C1573 B.n580 VSUBS 0.007576f
C1574 B.n581 VSUBS 0.007576f
C1575 B.n582 VSUBS 0.007576f
C1576 B.n583 VSUBS 0.007576f
C1577 B.n584 VSUBS 0.007576f
C1578 B.n585 VSUBS 0.007576f
C1579 B.n586 VSUBS 0.007576f
C1580 B.n587 VSUBS 0.007576f
C1581 B.n588 VSUBS 0.007576f
C1582 B.n589 VSUBS 0.007576f
C1583 B.n590 VSUBS 0.007576f
C1584 B.n591 VSUBS 0.007576f
C1585 B.n592 VSUBS 0.007576f
C1586 B.n593 VSUBS 0.007576f
C1587 B.n594 VSUBS 0.007576f
C1588 B.n595 VSUBS 0.007576f
C1589 B.n596 VSUBS 0.007576f
C1590 B.n597 VSUBS 0.007576f
C1591 B.n598 VSUBS 0.007576f
C1592 B.n599 VSUBS 0.007576f
C1593 B.n600 VSUBS 0.007576f
C1594 B.n601 VSUBS 0.007576f
C1595 B.n602 VSUBS 0.007576f
C1596 B.n603 VSUBS 0.007576f
C1597 B.n604 VSUBS 0.007576f
C1598 B.n605 VSUBS 0.007576f
C1599 B.n606 VSUBS 0.007576f
C1600 B.n607 VSUBS 0.007576f
C1601 B.n608 VSUBS 0.007576f
C1602 B.n609 VSUBS 0.007576f
C1603 B.n610 VSUBS 0.007576f
C1604 B.n611 VSUBS 0.007576f
C1605 B.n612 VSUBS 0.007576f
C1606 B.n613 VSUBS 0.007576f
C1607 B.n614 VSUBS 0.007576f
C1608 B.n615 VSUBS 0.007576f
C1609 B.n616 VSUBS 0.007576f
C1610 B.n617 VSUBS 0.007576f
C1611 B.n618 VSUBS 0.007576f
C1612 B.n619 VSUBS 0.007576f
C1613 B.n620 VSUBS 0.007576f
C1614 B.n621 VSUBS 0.007576f
C1615 B.n622 VSUBS 0.007576f
C1616 B.n623 VSUBS 0.007576f
C1617 B.n624 VSUBS 0.007576f
C1618 B.n625 VSUBS 0.007576f
C1619 B.n626 VSUBS 0.007576f
C1620 B.n627 VSUBS 0.007576f
C1621 B.n628 VSUBS 0.007576f
C1622 B.n629 VSUBS 0.007576f
C1623 B.n630 VSUBS 0.007576f
C1624 B.n631 VSUBS 0.007576f
C1625 B.n632 VSUBS 0.007576f
C1626 B.n633 VSUBS 0.007576f
C1627 B.n634 VSUBS 0.007576f
C1628 B.n635 VSUBS 0.007576f
C1629 B.n636 VSUBS 0.007576f
C1630 B.n637 VSUBS 0.007576f
C1631 B.n638 VSUBS 0.007576f
C1632 B.n639 VSUBS 0.007576f
C1633 B.n640 VSUBS 0.007576f
C1634 B.n641 VSUBS 0.007576f
C1635 B.n642 VSUBS 0.007576f
C1636 B.n643 VSUBS 0.007576f
C1637 B.n644 VSUBS 0.007576f
C1638 B.n645 VSUBS 0.007576f
C1639 B.n646 VSUBS 0.007576f
C1640 B.n647 VSUBS 0.007576f
C1641 B.n648 VSUBS 0.007576f
C1642 B.n649 VSUBS 0.007576f
C1643 B.n650 VSUBS 0.007576f
C1644 B.n651 VSUBS 0.007576f
C1645 B.n652 VSUBS 0.007576f
C1646 B.n653 VSUBS 0.007576f
C1647 B.n654 VSUBS 0.007576f
C1648 B.n655 VSUBS 0.007576f
C1649 B.n656 VSUBS 0.007576f
C1650 B.n657 VSUBS 0.007576f
C1651 B.n658 VSUBS 0.007576f
C1652 B.n659 VSUBS 0.007576f
C1653 B.n660 VSUBS 0.007576f
C1654 B.n661 VSUBS 0.007131f
C1655 B.n662 VSUBS 0.017554f
C1656 B.n663 VSUBS 0.004234f
C1657 B.n664 VSUBS 0.007576f
C1658 B.n665 VSUBS 0.007576f
C1659 B.n666 VSUBS 0.007576f
C1660 B.n667 VSUBS 0.007576f
C1661 B.n668 VSUBS 0.007576f
C1662 B.n669 VSUBS 0.007576f
C1663 B.n670 VSUBS 0.007576f
C1664 B.n671 VSUBS 0.007576f
C1665 B.n672 VSUBS 0.007576f
C1666 B.n673 VSUBS 0.007576f
C1667 B.n674 VSUBS 0.007576f
C1668 B.n675 VSUBS 0.007576f
C1669 B.n676 VSUBS 0.004234f
C1670 B.n677 VSUBS 0.007576f
C1671 B.n678 VSUBS 0.007576f
C1672 B.n679 VSUBS 0.007131f
C1673 B.n680 VSUBS 0.007576f
C1674 B.n681 VSUBS 0.007576f
C1675 B.n682 VSUBS 0.007576f
C1676 B.n683 VSUBS 0.007576f
C1677 B.n684 VSUBS 0.007576f
C1678 B.n685 VSUBS 0.007576f
C1679 B.n686 VSUBS 0.007576f
C1680 B.n687 VSUBS 0.007576f
C1681 B.n688 VSUBS 0.007576f
C1682 B.n689 VSUBS 0.007576f
C1683 B.n690 VSUBS 0.007576f
C1684 B.n691 VSUBS 0.007576f
C1685 B.n692 VSUBS 0.007576f
C1686 B.n693 VSUBS 0.007576f
C1687 B.n694 VSUBS 0.007576f
C1688 B.n695 VSUBS 0.007576f
C1689 B.n696 VSUBS 0.007576f
C1690 B.n697 VSUBS 0.007576f
C1691 B.n698 VSUBS 0.007576f
C1692 B.n699 VSUBS 0.007576f
C1693 B.n700 VSUBS 0.007576f
C1694 B.n701 VSUBS 0.007576f
C1695 B.n702 VSUBS 0.007576f
C1696 B.n703 VSUBS 0.007576f
C1697 B.n704 VSUBS 0.007576f
C1698 B.n705 VSUBS 0.007576f
C1699 B.n706 VSUBS 0.007576f
C1700 B.n707 VSUBS 0.007576f
C1701 B.n708 VSUBS 0.007576f
C1702 B.n709 VSUBS 0.007576f
C1703 B.n710 VSUBS 0.007576f
C1704 B.n711 VSUBS 0.007576f
C1705 B.n712 VSUBS 0.007576f
C1706 B.n713 VSUBS 0.007576f
C1707 B.n714 VSUBS 0.007576f
C1708 B.n715 VSUBS 0.007576f
C1709 B.n716 VSUBS 0.007576f
C1710 B.n717 VSUBS 0.007576f
C1711 B.n718 VSUBS 0.007576f
C1712 B.n719 VSUBS 0.007576f
C1713 B.n720 VSUBS 0.007576f
C1714 B.n721 VSUBS 0.007576f
C1715 B.n722 VSUBS 0.007576f
C1716 B.n723 VSUBS 0.007576f
C1717 B.n724 VSUBS 0.007576f
C1718 B.n725 VSUBS 0.007576f
C1719 B.n726 VSUBS 0.007576f
C1720 B.n727 VSUBS 0.007576f
C1721 B.n728 VSUBS 0.007576f
C1722 B.n729 VSUBS 0.007576f
C1723 B.n730 VSUBS 0.007576f
C1724 B.n731 VSUBS 0.007576f
C1725 B.n732 VSUBS 0.007576f
C1726 B.n733 VSUBS 0.007576f
C1727 B.n734 VSUBS 0.007576f
C1728 B.n735 VSUBS 0.007576f
C1729 B.n736 VSUBS 0.007576f
C1730 B.n737 VSUBS 0.007576f
C1731 B.n738 VSUBS 0.007576f
C1732 B.n739 VSUBS 0.007576f
C1733 B.n740 VSUBS 0.007576f
C1734 B.n741 VSUBS 0.007576f
C1735 B.n742 VSUBS 0.007576f
C1736 B.n743 VSUBS 0.007576f
C1737 B.n744 VSUBS 0.007576f
C1738 B.n745 VSUBS 0.007576f
C1739 B.n746 VSUBS 0.007576f
C1740 B.n747 VSUBS 0.007576f
C1741 B.n748 VSUBS 0.007576f
C1742 B.n749 VSUBS 0.007576f
C1743 B.n750 VSUBS 0.007576f
C1744 B.n751 VSUBS 0.007576f
C1745 B.n752 VSUBS 0.007576f
C1746 B.n753 VSUBS 0.007576f
C1747 B.n754 VSUBS 0.007576f
C1748 B.n755 VSUBS 0.007576f
C1749 B.n756 VSUBS 0.007576f
C1750 B.n757 VSUBS 0.007576f
C1751 B.n758 VSUBS 0.007576f
C1752 B.n759 VSUBS 0.007576f
C1753 B.n760 VSUBS 0.007576f
C1754 B.n761 VSUBS 0.007576f
C1755 B.n762 VSUBS 0.007576f
C1756 B.n763 VSUBS 0.007576f
C1757 B.n764 VSUBS 0.007576f
C1758 B.n765 VSUBS 0.007576f
C1759 B.n766 VSUBS 0.007576f
C1760 B.n767 VSUBS 0.007576f
C1761 B.n768 VSUBS 0.007576f
C1762 B.n769 VSUBS 0.007576f
C1763 B.n770 VSUBS 0.018719f
C1764 B.n771 VSUBS 0.01738f
C1765 B.n772 VSUBS 0.01738f
C1766 B.n773 VSUBS 0.007576f
C1767 B.n774 VSUBS 0.007576f
C1768 B.n775 VSUBS 0.007576f
C1769 B.n776 VSUBS 0.007576f
C1770 B.n777 VSUBS 0.007576f
C1771 B.n778 VSUBS 0.007576f
C1772 B.n779 VSUBS 0.007576f
C1773 B.n780 VSUBS 0.007576f
C1774 B.n781 VSUBS 0.007576f
C1775 B.n782 VSUBS 0.007576f
C1776 B.n783 VSUBS 0.007576f
C1777 B.n784 VSUBS 0.007576f
C1778 B.n785 VSUBS 0.007576f
C1779 B.n786 VSUBS 0.007576f
C1780 B.n787 VSUBS 0.007576f
C1781 B.n788 VSUBS 0.007576f
C1782 B.n789 VSUBS 0.007576f
C1783 B.n790 VSUBS 0.007576f
C1784 B.n791 VSUBS 0.007576f
C1785 B.n792 VSUBS 0.007576f
C1786 B.n793 VSUBS 0.007576f
C1787 B.n794 VSUBS 0.007576f
C1788 B.n795 VSUBS 0.007576f
C1789 B.n796 VSUBS 0.007576f
C1790 B.n797 VSUBS 0.007576f
C1791 B.n798 VSUBS 0.007576f
C1792 B.n799 VSUBS 0.007576f
C1793 B.n800 VSUBS 0.007576f
C1794 B.n801 VSUBS 0.007576f
C1795 B.n802 VSUBS 0.007576f
C1796 B.n803 VSUBS 0.007576f
C1797 B.n804 VSUBS 0.007576f
C1798 B.n805 VSUBS 0.007576f
C1799 B.n806 VSUBS 0.007576f
C1800 B.n807 VSUBS 0.007576f
C1801 B.n808 VSUBS 0.007576f
C1802 B.n809 VSUBS 0.007576f
C1803 B.n810 VSUBS 0.007576f
C1804 B.n811 VSUBS 0.007576f
C1805 B.n812 VSUBS 0.007576f
C1806 B.n813 VSUBS 0.007576f
C1807 B.n814 VSUBS 0.007576f
C1808 B.n815 VSUBS 0.007576f
C1809 B.n816 VSUBS 0.007576f
C1810 B.n817 VSUBS 0.007576f
C1811 B.n818 VSUBS 0.007576f
C1812 B.n819 VSUBS 0.007576f
C1813 B.n820 VSUBS 0.007576f
C1814 B.n821 VSUBS 0.007576f
C1815 B.n822 VSUBS 0.007576f
C1816 B.n823 VSUBS 0.017156f
.ends

