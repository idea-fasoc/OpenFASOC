* NGSPICE file created from diff_pair_sample_0653.ext - technology: sky130A

.subckt diff_pair_sample_0653 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.69
X1 VDD1.t4 VP.t1 VTAIL.t7 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.69
X2 VDD2.t5 VN.t0 VTAIL.t5 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.69
X3 B.t11 B.t9 B.t10 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.69
X4 B.t8 B.t6 B.t7 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.69
X5 VTAIL.t0 VN.t1 VDD2.t4 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.69
X6 VDD2.t3 VN.t2 VTAIL.t3 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.69
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.69
X8 VDD2.t1 VN.t4 VTAIL.t2 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.69
X9 VTAIL.t8 VP.t2 VDD1.t3 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.69
X10 B.t5 B.t3 B.t4 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.69
X11 B.t2 B.t0 B.t1 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0 ps=0 w=2.68 l=1.69
X12 VDD1.t2 VP.t3 VTAIL.t9 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=1.0452 ps=6.14 w=2.68 l=1.69
X13 VTAIL.t10 VP.t4 VDD1.t1 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.69
X14 VDD1.t0 VP.t5 VTAIL.t11 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=1.0452 pd=6.14 as=0.4422 ps=3.01 w=2.68 l=1.69
X15 VTAIL.t1 VN.t5 VDD2.t0 w_n2586_n1504# sky130_fd_pr__pfet_01v8 ad=0.4422 pd=3.01 as=0.4422 ps=3.01 w=2.68 l=1.69
R0 VP.n18 VP.n17 184.671
R1 VP.n33 VP.n32 184.671
R2 VP.n16 VP.n15 184.671
R3 VP.n10 VP.n9 161.3
R4 VP.n11 VP.n6 161.3
R5 VP.n13 VP.n12 161.3
R6 VP.n14 VP.n5 161.3
R7 VP.n31 VP.n0 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n28 VP.n1 161.3
R10 VP.n27 VP.n26 161.3
R11 VP.n25 VP.n2 161.3
R12 VP.n24 VP.n23 161.3
R13 VP.n22 VP.n3 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n19 VP.n4 161.3
R16 VP.n7 VP.t1 71.0458
R17 VP.n8 VP.n7 44.5457
R18 VP.n20 VP.n3 41.3843
R19 VP.n30 VP.n1 41.3843
R20 VP.n13 VP.n6 41.3843
R21 VP.n24 VP.n3 39.4369
R22 VP.n26 VP.n1 39.4369
R23 VP.n9 VP.n6 39.4369
R24 VP.n25 VP.t4 38.2183
R25 VP.n18 VP.t5 38.2183
R26 VP.n32 VP.t3 38.2183
R27 VP.n8 VP.t2 38.2183
R28 VP.n15 VP.t0 38.2183
R29 VP.n17 VP.n16 37.8793
R30 VP.n20 VP.n19 24.3439
R31 VP.n25 VP.n24 24.3439
R32 VP.n26 VP.n25 24.3439
R33 VP.n31 VP.n30 24.3439
R34 VP.n14 VP.n13 24.3439
R35 VP.n9 VP.n8 24.3439
R36 VP.n10 VP.n7 12.4931
R37 VP.n19 VP.n18 0.974237
R38 VP.n32 VP.n31 0.974237
R39 VP.n15 VP.n14 0.974237
R40 VP.n11 VP.n10 0.189894
R41 VP.n12 VP.n11 0.189894
R42 VP.n12 VP.n5 0.189894
R43 VP.n16 VP.n5 0.189894
R44 VP.n17 VP.n4 0.189894
R45 VP.n21 VP.n4 0.189894
R46 VP.n22 VP.n21 0.189894
R47 VP.n23 VP.n22 0.189894
R48 VP.n23 VP.n2 0.189894
R49 VP.n27 VP.n2 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n29 VP.n28 0.189894
R52 VP.n29 VP.n0 0.189894
R53 VP.n33 VP.n0 0.189894
R54 VP VP.n33 0.0516364
R55 VTAIL.n50 VTAIL.n44 756.745
R56 VTAIL.n8 VTAIL.n2 756.745
R57 VTAIL.n38 VTAIL.n32 756.745
R58 VTAIL.n24 VTAIL.n18 756.745
R59 VTAIL.n49 VTAIL.n48 585
R60 VTAIL.n51 VTAIL.n50 585
R61 VTAIL.n7 VTAIL.n6 585
R62 VTAIL.n9 VTAIL.n8 585
R63 VTAIL.n39 VTAIL.n38 585
R64 VTAIL.n37 VTAIL.n36 585
R65 VTAIL.n25 VTAIL.n24 585
R66 VTAIL.n23 VTAIL.n22 585
R67 VTAIL.n47 VTAIL.t2 357.269
R68 VTAIL.n5 VTAIL.t9 357.269
R69 VTAIL.n35 VTAIL.t6 357.269
R70 VTAIL.n21 VTAIL.t3 357.269
R71 VTAIL.n50 VTAIL.n49 171.744
R72 VTAIL.n8 VTAIL.n7 171.744
R73 VTAIL.n38 VTAIL.n37 171.744
R74 VTAIL.n24 VTAIL.n23 171.744
R75 VTAIL.n1 VTAIL.n0 134.899
R76 VTAIL.n15 VTAIL.n14 134.899
R77 VTAIL.n31 VTAIL.n30 134.899
R78 VTAIL.n17 VTAIL.n16 134.899
R79 VTAIL.n49 VTAIL.t2 85.8723
R80 VTAIL.n7 VTAIL.t9 85.8723
R81 VTAIL.n37 VTAIL.t6 85.8723
R82 VTAIL.n23 VTAIL.t3 85.8723
R83 VTAIL.n55 VTAIL.n54 30.6338
R84 VTAIL.n13 VTAIL.n12 30.6338
R85 VTAIL.n43 VTAIL.n42 30.6338
R86 VTAIL.n29 VTAIL.n28 30.6338
R87 VTAIL.n17 VTAIL.n15 18.16
R88 VTAIL.n55 VTAIL.n43 16.4186
R89 VTAIL.n0 VTAIL.t5 12.1292
R90 VTAIL.n0 VTAIL.t0 12.1292
R91 VTAIL.n14 VTAIL.t11 12.1292
R92 VTAIL.n14 VTAIL.t10 12.1292
R93 VTAIL.n30 VTAIL.t7 12.1292
R94 VTAIL.n30 VTAIL.t8 12.1292
R95 VTAIL.n16 VTAIL.t4 12.1292
R96 VTAIL.n16 VTAIL.t1 12.1292
R97 VTAIL.n48 VTAIL.n47 10.3978
R98 VTAIL.n6 VTAIL.n5 10.3978
R99 VTAIL.n36 VTAIL.n35 10.3978
R100 VTAIL.n22 VTAIL.n21 10.3978
R101 VTAIL.n54 VTAIL.n53 9.45567
R102 VTAIL.n12 VTAIL.n11 9.45567
R103 VTAIL.n42 VTAIL.n41 9.45567
R104 VTAIL.n28 VTAIL.n27 9.45567
R105 VTAIL.n46 VTAIL.n45 9.3005
R106 VTAIL.n53 VTAIL.n52 9.3005
R107 VTAIL.n4 VTAIL.n3 9.3005
R108 VTAIL.n11 VTAIL.n10 9.3005
R109 VTAIL.n34 VTAIL.n33 9.3005
R110 VTAIL.n41 VTAIL.n40 9.3005
R111 VTAIL.n27 VTAIL.n26 9.3005
R112 VTAIL.n20 VTAIL.n19 9.3005
R113 VTAIL.n54 VTAIL.n44 8.92171
R114 VTAIL.n12 VTAIL.n2 8.92171
R115 VTAIL.n42 VTAIL.n32 8.92171
R116 VTAIL.n28 VTAIL.n18 8.92171
R117 VTAIL.n52 VTAIL.n51 8.14595
R118 VTAIL.n10 VTAIL.n9 8.14595
R119 VTAIL.n40 VTAIL.n39 8.14595
R120 VTAIL.n26 VTAIL.n25 8.14595
R121 VTAIL.n48 VTAIL.n46 7.3702
R122 VTAIL.n6 VTAIL.n4 7.3702
R123 VTAIL.n36 VTAIL.n34 7.3702
R124 VTAIL.n22 VTAIL.n20 7.3702
R125 VTAIL.n51 VTAIL.n46 5.81868
R126 VTAIL.n9 VTAIL.n4 5.81868
R127 VTAIL.n39 VTAIL.n34 5.81868
R128 VTAIL.n25 VTAIL.n20 5.81868
R129 VTAIL.n52 VTAIL.n44 5.04292
R130 VTAIL.n10 VTAIL.n2 5.04292
R131 VTAIL.n40 VTAIL.n32 5.04292
R132 VTAIL.n26 VTAIL.n18 5.04292
R133 VTAIL.n47 VTAIL.n45 2.74506
R134 VTAIL.n5 VTAIL.n3 2.74506
R135 VTAIL.n35 VTAIL.n33 2.74506
R136 VTAIL.n21 VTAIL.n19 2.74506
R137 VTAIL.n29 VTAIL.n17 1.74188
R138 VTAIL.n43 VTAIL.n31 1.74188
R139 VTAIL.n15 VTAIL.n13 1.74188
R140 VTAIL.n31 VTAIL.n29 1.34102
R141 VTAIL.n13 VTAIL.n1 1.34102
R142 VTAIL VTAIL.n55 1.24834
R143 VTAIL VTAIL.n1 0.494034
R144 VTAIL.n53 VTAIL.n45 0.155672
R145 VTAIL.n11 VTAIL.n3 0.155672
R146 VTAIL.n41 VTAIL.n33 0.155672
R147 VTAIL.n27 VTAIL.n19 0.155672
R148 VDD1.n6 VDD1.n0 756.745
R149 VDD1.n17 VDD1.n11 756.745
R150 VDD1.n7 VDD1.n6 585
R151 VDD1.n5 VDD1.n4 585
R152 VDD1.n16 VDD1.n15 585
R153 VDD1.n18 VDD1.n17 585
R154 VDD1.n14 VDD1.t0 357.269
R155 VDD1.n3 VDD1.t4 357.269
R156 VDD1.n6 VDD1.n5 171.744
R157 VDD1.n17 VDD1.n16 171.744
R158 VDD1.n23 VDD1.n22 151.958
R159 VDD1.n25 VDD1.n24 151.577
R160 VDD1.n5 VDD1.t4 85.8723
R161 VDD1.n16 VDD1.t0 85.8723
R162 VDD1 VDD1.n10 48.6768
R163 VDD1.n23 VDD1.n21 48.5633
R164 VDD1.n25 VDD1.n23 33.1388
R165 VDD1.n24 VDD1.t3 12.1292
R166 VDD1.n24 VDD1.t5 12.1292
R167 VDD1.n22 VDD1.t1 12.1292
R168 VDD1.n22 VDD1.t2 12.1292
R169 VDD1.n4 VDD1.n3 10.3978
R170 VDD1.n15 VDD1.n14 10.3978
R171 VDD1.n10 VDD1.n9 9.45567
R172 VDD1.n21 VDD1.n20 9.45567
R173 VDD1.n9 VDD1.n8 9.3005
R174 VDD1.n2 VDD1.n1 9.3005
R175 VDD1.n13 VDD1.n12 9.3005
R176 VDD1.n20 VDD1.n19 9.3005
R177 VDD1.n10 VDD1.n0 8.92171
R178 VDD1.n21 VDD1.n11 8.92171
R179 VDD1.n8 VDD1.n7 8.14595
R180 VDD1.n19 VDD1.n18 8.14595
R181 VDD1.n4 VDD1.n2 7.3702
R182 VDD1.n15 VDD1.n13 7.3702
R183 VDD1.n7 VDD1.n2 5.81868
R184 VDD1.n18 VDD1.n13 5.81868
R185 VDD1.n8 VDD1.n0 5.04292
R186 VDD1.n19 VDD1.n11 5.04292
R187 VDD1.n3 VDD1.n1 2.74506
R188 VDD1.n14 VDD1.n12 2.74506
R189 VDD1 VDD1.n25 0.377655
R190 VDD1.n9 VDD1.n1 0.155672
R191 VDD1.n20 VDD1.n12 0.155672
R192 VN.n11 VN.n10 184.671
R193 VN.n23 VN.n22 184.671
R194 VN.n21 VN.n12 161.3
R195 VN.n20 VN.n19 161.3
R196 VN.n18 VN.n13 161.3
R197 VN.n17 VN.n16 161.3
R198 VN.n9 VN.n0 161.3
R199 VN.n8 VN.n7 161.3
R200 VN.n6 VN.n1 161.3
R201 VN.n5 VN.n4 161.3
R202 VN.n2 VN.t0 71.0458
R203 VN.n14 VN.t2 71.0458
R204 VN.n15 VN.n14 44.5457
R205 VN.n3 VN.n2 44.5457
R206 VN.n8 VN.n1 41.3843
R207 VN.n20 VN.n13 41.3843
R208 VN.n4 VN.n1 39.4369
R209 VN.n16 VN.n13 39.4369
R210 VN VN.n23 38.26
R211 VN.n3 VN.t1 38.2183
R212 VN.n10 VN.t4 38.2183
R213 VN.n15 VN.t5 38.2183
R214 VN.n22 VN.t3 38.2183
R215 VN.n4 VN.n3 24.3439
R216 VN.n9 VN.n8 24.3439
R217 VN.n16 VN.n15 24.3439
R218 VN.n21 VN.n20 24.3439
R219 VN.n17 VN.n14 12.4931
R220 VN.n5 VN.n2 12.4931
R221 VN.n10 VN.n9 0.974237
R222 VN.n22 VN.n21 0.974237
R223 VN.n23 VN.n12 0.189894
R224 VN.n19 VN.n12 0.189894
R225 VN.n19 VN.n18 0.189894
R226 VN.n18 VN.n17 0.189894
R227 VN.n6 VN.n5 0.189894
R228 VN.n7 VN.n6 0.189894
R229 VN.n7 VN.n0 0.189894
R230 VN.n11 VN.n0 0.189894
R231 VN VN.n11 0.0516364
R232 VDD2.n19 VDD2.n13 756.745
R233 VDD2.n6 VDD2.n0 756.745
R234 VDD2.n20 VDD2.n19 585
R235 VDD2.n18 VDD2.n17 585
R236 VDD2.n5 VDD2.n4 585
R237 VDD2.n7 VDD2.n6 585
R238 VDD2.n3 VDD2.t5 357.269
R239 VDD2.n16 VDD2.t2 357.269
R240 VDD2.n19 VDD2.n18 171.744
R241 VDD2.n6 VDD2.n5 171.744
R242 VDD2.n12 VDD2.n11 151.958
R243 VDD2 VDD2.n25 151.954
R244 VDD2.n18 VDD2.t2 85.8723
R245 VDD2.n5 VDD2.t5 85.8723
R246 VDD2.n12 VDD2.n10 48.5633
R247 VDD2.n24 VDD2.n23 47.3126
R248 VDD2.n24 VDD2.n12 31.6851
R249 VDD2.n25 VDD2.t0 12.1292
R250 VDD2.n25 VDD2.t3 12.1292
R251 VDD2.n11 VDD2.t4 12.1292
R252 VDD2.n11 VDD2.t1 12.1292
R253 VDD2.n17 VDD2.n16 10.3978
R254 VDD2.n4 VDD2.n3 10.3978
R255 VDD2.n23 VDD2.n22 9.45567
R256 VDD2.n10 VDD2.n9 9.45567
R257 VDD2.n22 VDD2.n21 9.3005
R258 VDD2.n15 VDD2.n14 9.3005
R259 VDD2.n2 VDD2.n1 9.3005
R260 VDD2.n9 VDD2.n8 9.3005
R261 VDD2.n23 VDD2.n13 8.92171
R262 VDD2.n10 VDD2.n0 8.92171
R263 VDD2.n21 VDD2.n20 8.14595
R264 VDD2.n8 VDD2.n7 8.14595
R265 VDD2.n17 VDD2.n15 7.3702
R266 VDD2.n4 VDD2.n2 7.3702
R267 VDD2.n20 VDD2.n15 5.81868
R268 VDD2.n7 VDD2.n2 5.81868
R269 VDD2.n21 VDD2.n13 5.04292
R270 VDD2.n8 VDD2.n0 5.04292
R271 VDD2.n16 VDD2.n14 2.74506
R272 VDD2.n3 VDD2.n1 2.74506
R273 VDD2 VDD2.n24 1.36472
R274 VDD2.n22 VDD2.n14 0.155672
R275 VDD2.n9 VDD2.n1 0.155672
R276 B.n316 B.n41 585
R277 B.n318 B.n317 585
R278 B.n319 B.n40 585
R279 B.n321 B.n320 585
R280 B.n322 B.n39 585
R281 B.n324 B.n323 585
R282 B.n325 B.n38 585
R283 B.n327 B.n326 585
R284 B.n328 B.n37 585
R285 B.n330 B.n329 585
R286 B.n331 B.n36 585
R287 B.n333 B.n332 585
R288 B.n334 B.n35 585
R289 B.n336 B.n335 585
R290 B.n338 B.n337 585
R291 B.n339 B.n31 585
R292 B.n341 B.n340 585
R293 B.n342 B.n30 585
R294 B.n344 B.n343 585
R295 B.n345 B.n29 585
R296 B.n347 B.n346 585
R297 B.n348 B.n28 585
R298 B.n350 B.n349 585
R299 B.n351 B.n25 585
R300 B.n354 B.n353 585
R301 B.n355 B.n24 585
R302 B.n357 B.n356 585
R303 B.n358 B.n23 585
R304 B.n360 B.n359 585
R305 B.n361 B.n22 585
R306 B.n363 B.n362 585
R307 B.n364 B.n21 585
R308 B.n366 B.n365 585
R309 B.n367 B.n20 585
R310 B.n369 B.n368 585
R311 B.n370 B.n19 585
R312 B.n372 B.n371 585
R313 B.n373 B.n18 585
R314 B.n315 B.n314 585
R315 B.n313 B.n42 585
R316 B.n312 B.n311 585
R317 B.n310 B.n43 585
R318 B.n309 B.n308 585
R319 B.n307 B.n44 585
R320 B.n306 B.n305 585
R321 B.n304 B.n45 585
R322 B.n303 B.n302 585
R323 B.n301 B.n46 585
R324 B.n300 B.n299 585
R325 B.n298 B.n47 585
R326 B.n297 B.n296 585
R327 B.n295 B.n48 585
R328 B.n294 B.n293 585
R329 B.n292 B.n49 585
R330 B.n291 B.n290 585
R331 B.n289 B.n50 585
R332 B.n288 B.n287 585
R333 B.n286 B.n51 585
R334 B.n285 B.n284 585
R335 B.n283 B.n52 585
R336 B.n282 B.n281 585
R337 B.n280 B.n53 585
R338 B.n279 B.n278 585
R339 B.n277 B.n54 585
R340 B.n276 B.n275 585
R341 B.n274 B.n55 585
R342 B.n273 B.n272 585
R343 B.n271 B.n56 585
R344 B.n270 B.n269 585
R345 B.n268 B.n57 585
R346 B.n267 B.n266 585
R347 B.n265 B.n58 585
R348 B.n264 B.n263 585
R349 B.n262 B.n59 585
R350 B.n261 B.n260 585
R351 B.n259 B.n60 585
R352 B.n258 B.n257 585
R353 B.n256 B.n61 585
R354 B.n255 B.n254 585
R355 B.n253 B.n62 585
R356 B.n252 B.n251 585
R357 B.n250 B.n63 585
R358 B.n249 B.n248 585
R359 B.n247 B.n64 585
R360 B.n246 B.n245 585
R361 B.n244 B.n65 585
R362 B.n243 B.n242 585
R363 B.n241 B.n66 585
R364 B.n240 B.n239 585
R365 B.n238 B.n67 585
R366 B.n237 B.n236 585
R367 B.n235 B.n68 585
R368 B.n234 B.n233 585
R369 B.n232 B.n69 585
R370 B.n231 B.n230 585
R371 B.n229 B.n70 585
R372 B.n228 B.n227 585
R373 B.n226 B.n71 585
R374 B.n225 B.n224 585
R375 B.n223 B.n72 585
R376 B.n222 B.n221 585
R377 B.n220 B.n73 585
R378 B.n219 B.n218 585
R379 B.n160 B.n97 585
R380 B.n162 B.n161 585
R381 B.n163 B.n96 585
R382 B.n165 B.n164 585
R383 B.n166 B.n95 585
R384 B.n168 B.n167 585
R385 B.n169 B.n94 585
R386 B.n171 B.n170 585
R387 B.n172 B.n93 585
R388 B.n174 B.n173 585
R389 B.n175 B.n92 585
R390 B.n177 B.n176 585
R391 B.n178 B.n91 585
R392 B.n180 B.n179 585
R393 B.n182 B.n181 585
R394 B.n183 B.n87 585
R395 B.n185 B.n184 585
R396 B.n186 B.n86 585
R397 B.n188 B.n187 585
R398 B.n189 B.n85 585
R399 B.n191 B.n190 585
R400 B.n192 B.n84 585
R401 B.n194 B.n193 585
R402 B.n195 B.n81 585
R403 B.n198 B.n197 585
R404 B.n199 B.n80 585
R405 B.n201 B.n200 585
R406 B.n202 B.n79 585
R407 B.n204 B.n203 585
R408 B.n205 B.n78 585
R409 B.n207 B.n206 585
R410 B.n208 B.n77 585
R411 B.n210 B.n209 585
R412 B.n211 B.n76 585
R413 B.n213 B.n212 585
R414 B.n214 B.n75 585
R415 B.n216 B.n215 585
R416 B.n217 B.n74 585
R417 B.n159 B.n158 585
R418 B.n157 B.n98 585
R419 B.n156 B.n155 585
R420 B.n154 B.n99 585
R421 B.n153 B.n152 585
R422 B.n151 B.n100 585
R423 B.n150 B.n149 585
R424 B.n148 B.n101 585
R425 B.n147 B.n146 585
R426 B.n145 B.n102 585
R427 B.n144 B.n143 585
R428 B.n142 B.n103 585
R429 B.n141 B.n140 585
R430 B.n139 B.n104 585
R431 B.n138 B.n137 585
R432 B.n136 B.n105 585
R433 B.n135 B.n134 585
R434 B.n133 B.n106 585
R435 B.n132 B.n131 585
R436 B.n130 B.n107 585
R437 B.n129 B.n128 585
R438 B.n127 B.n108 585
R439 B.n126 B.n125 585
R440 B.n124 B.n109 585
R441 B.n123 B.n122 585
R442 B.n121 B.n110 585
R443 B.n120 B.n119 585
R444 B.n118 B.n111 585
R445 B.n117 B.n116 585
R446 B.n115 B.n112 585
R447 B.n114 B.n113 585
R448 B.n2 B.n0 585
R449 B.n421 B.n1 585
R450 B.n420 B.n419 585
R451 B.n418 B.n3 585
R452 B.n417 B.n416 585
R453 B.n415 B.n4 585
R454 B.n414 B.n413 585
R455 B.n412 B.n5 585
R456 B.n411 B.n410 585
R457 B.n409 B.n6 585
R458 B.n408 B.n407 585
R459 B.n406 B.n7 585
R460 B.n405 B.n404 585
R461 B.n403 B.n8 585
R462 B.n402 B.n401 585
R463 B.n400 B.n9 585
R464 B.n399 B.n398 585
R465 B.n397 B.n10 585
R466 B.n396 B.n395 585
R467 B.n394 B.n11 585
R468 B.n393 B.n392 585
R469 B.n391 B.n12 585
R470 B.n390 B.n389 585
R471 B.n388 B.n13 585
R472 B.n387 B.n386 585
R473 B.n385 B.n14 585
R474 B.n384 B.n383 585
R475 B.n382 B.n15 585
R476 B.n381 B.n380 585
R477 B.n379 B.n16 585
R478 B.n378 B.n377 585
R479 B.n376 B.n17 585
R480 B.n375 B.n374 585
R481 B.n423 B.n422 585
R482 B.n158 B.n97 478.086
R483 B.n374 B.n373 478.086
R484 B.n218 B.n217 478.086
R485 B.n314 B.n41 478.086
R486 B.n82 B.t11 266.918
R487 B.n32 B.t1 266.918
R488 B.n88 B.t5 266.918
R489 B.n26 B.t7 266.918
R490 B.n82 B.t9 244.302
R491 B.n88 B.t3 244.302
R492 B.n26 B.t6 244.302
R493 B.n32 B.t0 244.302
R494 B.n83 B.t10 227.743
R495 B.n33 B.t2 227.743
R496 B.n89 B.t4 227.743
R497 B.n27 B.t8 227.743
R498 B.n158 B.n157 163.367
R499 B.n157 B.n156 163.367
R500 B.n156 B.n99 163.367
R501 B.n152 B.n99 163.367
R502 B.n152 B.n151 163.367
R503 B.n151 B.n150 163.367
R504 B.n150 B.n101 163.367
R505 B.n146 B.n101 163.367
R506 B.n146 B.n145 163.367
R507 B.n145 B.n144 163.367
R508 B.n144 B.n103 163.367
R509 B.n140 B.n103 163.367
R510 B.n140 B.n139 163.367
R511 B.n139 B.n138 163.367
R512 B.n138 B.n105 163.367
R513 B.n134 B.n105 163.367
R514 B.n134 B.n133 163.367
R515 B.n133 B.n132 163.367
R516 B.n132 B.n107 163.367
R517 B.n128 B.n107 163.367
R518 B.n128 B.n127 163.367
R519 B.n127 B.n126 163.367
R520 B.n126 B.n109 163.367
R521 B.n122 B.n109 163.367
R522 B.n122 B.n121 163.367
R523 B.n121 B.n120 163.367
R524 B.n120 B.n111 163.367
R525 B.n116 B.n111 163.367
R526 B.n116 B.n115 163.367
R527 B.n115 B.n114 163.367
R528 B.n114 B.n2 163.367
R529 B.n422 B.n2 163.367
R530 B.n422 B.n421 163.367
R531 B.n421 B.n420 163.367
R532 B.n420 B.n3 163.367
R533 B.n416 B.n3 163.367
R534 B.n416 B.n415 163.367
R535 B.n415 B.n414 163.367
R536 B.n414 B.n5 163.367
R537 B.n410 B.n5 163.367
R538 B.n410 B.n409 163.367
R539 B.n409 B.n408 163.367
R540 B.n408 B.n7 163.367
R541 B.n404 B.n7 163.367
R542 B.n404 B.n403 163.367
R543 B.n403 B.n402 163.367
R544 B.n402 B.n9 163.367
R545 B.n398 B.n9 163.367
R546 B.n398 B.n397 163.367
R547 B.n397 B.n396 163.367
R548 B.n396 B.n11 163.367
R549 B.n392 B.n11 163.367
R550 B.n392 B.n391 163.367
R551 B.n391 B.n390 163.367
R552 B.n390 B.n13 163.367
R553 B.n386 B.n13 163.367
R554 B.n386 B.n385 163.367
R555 B.n385 B.n384 163.367
R556 B.n384 B.n15 163.367
R557 B.n380 B.n15 163.367
R558 B.n380 B.n379 163.367
R559 B.n379 B.n378 163.367
R560 B.n378 B.n17 163.367
R561 B.n374 B.n17 163.367
R562 B.n162 B.n97 163.367
R563 B.n163 B.n162 163.367
R564 B.n164 B.n163 163.367
R565 B.n164 B.n95 163.367
R566 B.n168 B.n95 163.367
R567 B.n169 B.n168 163.367
R568 B.n170 B.n169 163.367
R569 B.n170 B.n93 163.367
R570 B.n174 B.n93 163.367
R571 B.n175 B.n174 163.367
R572 B.n176 B.n175 163.367
R573 B.n176 B.n91 163.367
R574 B.n180 B.n91 163.367
R575 B.n181 B.n180 163.367
R576 B.n181 B.n87 163.367
R577 B.n185 B.n87 163.367
R578 B.n186 B.n185 163.367
R579 B.n187 B.n186 163.367
R580 B.n187 B.n85 163.367
R581 B.n191 B.n85 163.367
R582 B.n192 B.n191 163.367
R583 B.n193 B.n192 163.367
R584 B.n193 B.n81 163.367
R585 B.n198 B.n81 163.367
R586 B.n199 B.n198 163.367
R587 B.n200 B.n199 163.367
R588 B.n200 B.n79 163.367
R589 B.n204 B.n79 163.367
R590 B.n205 B.n204 163.367
R591 B.n206 B.n205 163.367
R592 B.n206 B.n77 163.367
R593 B.n210 B.n77 163.367
R594 B.n211 B.n210 163.367
R595 B.n212 B.n211 163.367
R596 B.n212 B.n75 163.367
R597 B.n216 B.n75 163.367
R598 B.n217 B.n216 163.367
R599 B.n218 B.n73 163.367
R600 B.n222 B.n73 163.367
R601 B.n223 B.n222 163.367
R602 B.n224 B.n223 163.367
R603 B.n224 B.n71 163.367
R604 B.n228 B.n71 163.367
R605 B.n229 B.n228 163.367
R606 B.n230 B.n229 163.367
R607 B.n230 B.n69 163.367
R608 B.n234 B.n69 163.367
R609 B.n235 B.n234 163.367
R610 B.n236 B.n235 163.367
R611 B.n236 B.n67 163.367
R612 B.n240 B.n67 163.367
R613 B.n241 B.n240 163.367
R614 B.n242 B.n241 163.367
R615 B.n242 B.n65 163.367
R616 B.n246 B.n65 163.367
R617 B.n247 B.n246 163.367
R618 B.n248 B.n247 163.367
R619 B.n248 B.n63 163.367
R620 B.n252 B.n63 163.367
R621 B.n253 B.n252 163.367
R622 B.n254 B.n253 163.367
R623 B.n254 B.n61 163.367
R624 B.n258 B.n61 163.367
R625 B.n259 B.n258 163.367
R626 B.n260 B.n259 163.367
R627 B.n260 B.n59 163.367
R628 B.n264 B.n59 163.367
R629 B.n265 B.n264 163.367
R630 B.n266 B.n265 163.367
R631 B.n266 B.n57 163.367
R632 B.n270 B.n57 163.367
R633 B.n271 B.n270 163.367
R634 B.n272 B.n271 163.367
R635 B.n272 B.n55 163.367
R636 B.n276 B.n55 163.367
R637 B.n277 B.n276 163.367
R638 B.n278 B.n277 163.367
R639 B.n278 B.n53 163.367
R640 B.n282 B.n53 163.367
R641 B.n283 B.n282 163.367
R642 B.n284 B.n283 163.367
R643 B.n284 B.n51 163.367
R644 B.n288 B.n51 163.367
R645 B.n289 B.n288 163.367
R646 B.n290 B.n289 163.367
R647 B.n290 B.n49 163.367
R648 B.n294 B.n49 163.367
R649 B.n295 B.n294 163.367
R650 B.n296 B.n295 163.367
R651 B.n296 B.n47 163.367
R652 B.n300 B.n47 163.367
R653 B.n301 B.n300 163.367
R654 B.n302 B.n301 163.367
R655 B.n302 B.n45 163.367
R656 B.n306 B.n45 163.367
R657 B.n307 B.n306 163.367
R658 B.n308 B.n307 163.367
R659 B.n308 B.n43 163.367
R660 B.n312 B.n43 163.367
R661 B.n313 B.n312 163.367
R662 B.n314 B.n313 163.367
R663 B.n373 B.n372 163.367
R664 B.n372 B.n19 163.367
R665 B.n368 B.n19 163.367
R666 B.n368 B.n367 163.367
R667 B.n367 B.n366 163.367
R668 B.n366 B.n21 163.367
R669 B.n362 B.n21 163.367
R670 B.n362 B.n361 163.367
R671 B.n361 B.n360 163.367
R672 B.n360 B.n23 163.367
R673 B.n356 B.n23 163.367
R674 B.n356 B.n355 163.367
R675 B.n355 B.n354 163.367
R676 B.n354 B.n25 163.367
R677 B.n349 B.n25 163.367
R678 B.n349 B.n348 163.367
R679 B.n348 B.n347 163.367
R680 B.n347 B.n29 163.367
R681 B.n343 B.n29 163.367
R682 B.n343 B.n342 163.367
R683 B.n342 B.n341 163.367
R684 B.n341 B.n31 163.367
R685 B.n337 B.n31 163.367
R686 B.n337 B.n336 163.367
R687 B.n336 B.n35 163.367
R688 B.n332 B.n35 163.367
R689 B.n332 B.n331 163.367
R690 B.n331 B.n330 163.367
R691 B.n330 B.n37 163.367
R692 B.n326 B.n37 163.367
R693 B.n326 B.n325 163.367
R694 B.n325 B.n324 163.367
R695 B.n324 B.n39 163.367
R696 B.n320 B.n39 163.367
R697 B.n320 B.n319 163.367
R698 B.n319 B.n318 163.367
R699 B.n318 B.n41 163.367
R700 B.n196 B.n83 59.5399
R701 B.n90 B.n89 59.5399
R702 B.n352 B.n27 59.5399
R703 B.n34 B.n33 59.5399
R704 B.n83 B.n82 39.1763
R705 B.n89 B.n88 39.1763
R706 B.n27 B.n26 39.1763
R707 B.n33 B.n32 39.1763
R708 B.n375 B.n18 31.0639
R709 B.n316 B.n315 31.0639
R710 B.n219 B.n74 31.0639
R711 B.n160 B.n159 31.0639
R712 B B.n423 18.0485
R713 B.n371 B.n18 10.6151
R714 B.n371 B.n370 10.6151
R715 B.n370 B.n369 10.6151
R716 B.n369 B.n20 10.6151
R717 B.n365 B.n20 10.6151
R718 B.n365 B.n364 10.6151
R719 B.n364 B.n363 10.6151
R720 B.n363 B.n22 10.6151
R721 B.n359 B.n22 10.6151
R722 B.n359 B.n358 10.6151
R723 B.n358 B.n357 10.6151
R724 B.n357 B.n24 10.6151
R725 B.n353 B.n24 10.6151
R726 B.n351 B.n350 10.6151
R727 B.n350 B.n28 10.6151
R728 B.n346 B.n28 10.6151
R729 B.n346 B.n345 10.6151
R730 B.n345 B.n344 10.6151
R731 B.n344 B.n30 10.6151
R732 B.n340 B.n30 10.6151
R733 B.n340 B.n339 10.6151
R734 B.n339 B.n338 10.6151
R735 B.n335 B.n334 10.6151
R736 B.n334 B.n333 10.6151
R737 B.n333 B.n36 10.6151
R738 B.n329 B.n36 10.6151
R739 B.n329 B.n328 10.6151
R740 B.n328 B.n327 10.6151
R741 B.n327 B.n38 10.6151
R742 B.n323 B.n38 10.6151
R743 B.n323 B.n322 10.6151
R744 B.n322 B.n321 10.6151
R745 B.n321 B.n40 10.6151
R746 B.n317 B.n40 10.6151
R747 B.n317 B.n316 10.6151
R748 B.n220 B.n219 10.6151
R749 B.n221 B.n220 10.6151
R750 B.n221 B.n72 10.6151
R751 B.n225 B.n72 10.6151
R752 B.n226 B.n225 10.6151
R753 B.n227 B.n226 10.6151
R754 B.n227 B.n70 10.6151
R755 B.n231 B.n70 10.6151
R756 B.n232 B.n231 10.6151
R757 B.n233 B.n232 10.6151
R758 B.n233 B.n68 10.6151
R759 B.n237 B.n68 10.6151
R760 B.n238 B.n237 10.6151
R761 B.n239 B.n238 10.6151
R762 B.n239 B.n66 10.6151
R763 B.n243 B.n66 10.6151
R764 B.n244 B.n243 10.6151
R765 B.n245 B.n244 10.6151
R766 B.n245 B.n64 10.6151
R767 B.n249 B.n64 10.6151
R768 B.n250 B.n249 10.6151
R769 B.n251 B.n250 10.6151
R770 B.n251 B.n62 10.6151
R771 B.n255 B.n62 10.6151
R772 B.n256 B.n255 10.6151
R773 B.n257 B.n256 10.6151
R774 B.n257 B.n60 10.6151
R775 B.n261 B.n60 10.6151
R776 B.n262 B.n261 10.6151
R777 B.n263 B.n262 10.6151
R778 B.n263 B.n58 10.6151
R779 B.n267 B.n58 10.6151
R780 B.n268 B.n267 10.6151
R781 B.n269 B.n268 10.6151
R782 B.n269 B.n56 10.6151
R783 B.n273 B.n56 10.6151
R784 B.n274 B.n273 10.6151
R785 B.n275 B.n274 10.6151
R786 B.n275 B.n54 10.6151
R787 B.n279 B.n54 10.6151
R788 B.n280 B.n279 10.6151
R789 B.n281 B.n280 10.6151
R790 B.n281 B.n52 10.6151
R791 B.n285 B.n52 10.6151
R792 B.n286 B.n285 10.6151
R793 B.n287 B.n286 10.6151
R794 B.n287 B.n50 10.6151
R795 B.n291 B.n50 10.6151
R796 B.n292 B.n291 10.6151
R797 B.n293 B.n292 10.6151
R798 B.n293 B.n48 10.6151
R799 B.n297 B.n48 10.6151
R800 B.n298 B.n297 10.6151
R801 B.n299 B.n298 10.6151
R802 B.n299 B.n46 10.6151
R803 B.n303 B.n46 10.6151
R804 B.n304 B.n303 10.6151
R805 B.n305 B.n304 10.6151
R806 B.n305 B.n44 10.6151
R807 B.n309 B.n44 10.6151
R808 B.n310 B.n309 10.6151
R809 B.n311 B.n310 10.6151
R810 B.n311 B.n42 10.6151
R811 B.n315 B.n42 10.6151
R812 B.n161 B.n160 10.6151
R813 B.n161 B.n96 10.6151
R814 B.n165 B.n96 10.6151
R815 B.n166 B.n165 10.6151
R816 B.n167 B.n166 10.6151
R817 B.n167 B.n94 10.6151
R818 B.n171 B.n94 10.6151
R819 B.n172 B.n171 10.6151
R820 B.n173 B.n172 10.6151
R821 B.n173 B.n92 10.6151
R822 B.n177 B.n92 10.6151
R823 B.n178 B.n177 10.6151
R824 B.n179 B.n178 10.6151
R825 B.n183 B.n182 10.6151
R826 B.n184 B.n183 10.6151
R827 B.n184 B.n86 10.6151
R828 B.n188 B.n86 10.6151
R829 B.n189 B.n188 10.6151
R830 B.n190 B.n189 10.6151
R831 B.n190 B.n84 10.6151
R832 B.n194 B.n84 10.6151
R833 B.n195 B.n194 10.6151
R834 B.n197 B.n80 10.6151
R835 B.n201 B.n80 10.6151
R836 B.n202 B.n201 10.6151
R837 B.n203 B.n202 10.6151
R838 B.n203 B.n78 10.6151
R839 B.n207 B.n78 10.6151
R840 B.n208 B.n207 10.6151
R841 B.n209 B.n208 10.6151
R842 B.n209 B.n76 10.6151
R843 B.n213 B.n76 10.6151
R844 B.n214 B.n213 10.6151
R845 B.n215 B.n214 10.6151
R846 B.n215 B.n74 10.6151
R847 B.n159 B.n98 10.6151
R848 B.n155 B.n98 10.6151
R849 B.n155 B.n154 10.6151
R850 B.n154 B.n153 10.6151
R851 B.n153 B.n100 10.6151
R852 B.n149 B.n100 10.6151
R853 B.n149 B.n148 10.6151
R854 B.n148 B.n147 10.6151
R855 B.n147 B.n102 10.6151
R856 B.n143 B.n102 10.6151
R857 B.n143 B.n142 10.6151
R858 B.n142 B.n141 10.6151
R859 B.n141 B.n104 10.6151
R860 B.n137 B.n104 10.6151
R861 B.n137 B.n136 10.6151
R862 B.n136 B.n135 10.6151
R863 B.n135 B.n106 10.6151
R864 B.n131 B.n106 10.6151
R865 B.n131 B.n130 10.6151
R866 B.n130 B.n129 10.6151
R867 B.n129 B.n108 10.6151
R868 B.n125 B.n108 10.6151
R869 B.n125 B.n124 10.6151
R870 B.n124 B.n123 10.6151
R871 B.n123 B.n110 10.6151
R872 B.n119 B.n110 10.6151
R873 B.n119 B.n118 10.6151
R874 B.n118 B.n117 10.6151
R875 B.n117 B.n112 10.6151
R876 B.n113 B.n112 10.6151
R877 B.n113 B.n0 10.6151
R878 B.n419 B.n1 10.6151
R879 B.n419 B.n418 10.6151
R880 B.n418 B.n417 10.6151
R881 B.n417 B.n4 10.6151
R882 B.n413 B.n4 10.6151
R883 B.n413 B.n412 10.6151
R884 B.n412 B.n411 10.6151
R885 B.n411 B.n6 10.6151
R886 B.n407 B.n6 10.6151
R887 B.n407 B.n406 10.6151
R888 B.n406 B.n405 10.6151
R889 B.n405 B.n8 10.6151
R890 B.n401 B.n8 10.6151
R891 B.n401 B.n400 10.6151
R892 B.n400 B.n399 10.6151
R893 B.n399 B.n10 10.6151
R894 B.n395 B.n10 10.6151
R895 B.n395 B.n394 10.6151
R896 B.n394 B.n393 10.6151
R897 B.n393 B.n12 10.6151
R898 B.n389 B.n12 10.6151
R899 B.n389 B.n388 10.6151
R900 B.n388 B.n387 10.6151
R901 B.n387 B.n14 10.6151
R902 B.n383 B.n14 10.6151
R903 B.n383 B.n382 10.6151
R904 B.n382 B.n381 10.6151
R905 B.n381 B.n16 10.6151
R906 B.n377 B.n16 10.6151
R907 B.n377 B.n376 10.6151
R908 B.n376 B.n375 10.6151
R909 B.n353 B.n352 9.36635
R910 B.n335 B.n34 9.36635
R911 B.n179 B.n90 9.36635
R912 B.n197 B.n196 9.36635
R913 B.n423 B.n0 2.81026
R914 B.n423 B.n1 2.81026
R915 B.n352 B.n351 1.24928
R916 B.n338 B.n34 1.24928
R917 B.n182 B.n90 1.24928
R918 B.n196 B.n195 1.24928
C0 VDD2 VTAIL 3.85625f
C1 B VDD1 1.13076f
C2 VP B 1.40685f
C3 VP VDD1 1.8792f
C4 B VTAIL 1.30472f
C5 VDD1 VTAIL 3.80968f
C6 VN w_n2586_n1504# 4.51113f
C7 VP VTAIL 2.15012f
C8 VDD2 w_n2586_n1504# 1.45426f
C9 VN VDD2 1.6499f
C10 B w_n2586_n1504# 5.81956f
C11 VN B 0.857976f
C12 w_n2586_n1504# VDD1 1.39896f
C13 B VDD2 1.18327f
C14 VN VDD1 0.154439f
C15 VDD2 VDD1 1.07588f
C16 VP w_n2586_n1504# 4.84006f
C17 VN VP 4.32997f
C18 VP VDD2 0.385887f
C19 w_n2586_n1504# VTAIL 1.52103f
C20 VN VTAIL 2.13595f
C21 VDD2 VSUBS 0.888155f
C22 VDD1 VSUBS 1.048041f
C23 VTAIL VSUBS 0.451448f
C24 VN VSUBS 4.44485f
C25 VP VSUBS 1.706112f
C26 B VSUBS 2.791616f
C27 w_n2586_n1504# VSUBS 49.3719f
C28 B.n0 VSUBS 0.005109f
C29 B.n1 VSUBS 0.005109f
C30 B.n2 VSUBS 0.00808f
C31 B.n3 VSUBS 0.00808f
C32 B.n4 VSUBS 0.00808f
C33 B.n5 VSUBS 0.00808f
C34 B.n6 VSUBS 0.00808f
C35 B.n7 VSUBS 0.00808f
C36 B.n8 VSUBS 0.00808f
C37 B.n9 VSUBS 0.00808f
C38 B.n10 VSUBS 0.00808f
C39 B.n11 VSUBS 0.00808f
C40 B.n12 VSUBS 0.00808f
C41 B.n13 VSUBS 0.00808f
C42 B.n14 VSUBS 0.00808f
C43 B.n15 VSUBS 0.00808f
C44 B.n16 VSUBS 0.00808f
C45 B.n17 VSUBS 0.00808f
C46 B.n18 VSUBS 0.018678f
C47 B.n19 VSUBS 0.00808f
C48 B.n20 VSUBS 0.00808f
C49 B.n21 VSUBS 0.00808f
C50 B.n22 VSUBS 0.00808f
C51 B.n23 VSUBS 0.00808f
C52 B.n24 VSUBS 0.00808f
C53 B.n25 VSUBS 0.00808f
C54 B.t8 VSUBS 0.048261f
C55 B.t7 VSUBS 0.060176f
C56 B.t6 VSUBS 0.252014f
C57 B.n26 VSUBS 0.105412f
C58 B.n27 VSUBS 0.092707f
C59 B.n28 VSUBS 0.00808f
C60 B.n29 VSUBS 0.00808f
C61 B.n30 VSUBS 0.00808f
C62 B.n31 VSUBS 0.00808f
C63 B.t2 VSUBS 0.048262f
C64 B.t1 VSUBS 0.060177f
C65 B.t0 VSUBS 0.252014f
C66 B.n32 VSUBS 0.105412f
C67 B.n33 VSUBS 0.092707f
C68 B.n34 VSUBS 0.018721f
C69 B.n35 VSUBS 0.00808f
C70 B.n36 VSUBS 0.00808f
C71 B.n37 VSUBS 0.00808f
C72 B.n38 VSUBS 0.00808f
C73 B.n39 VSUBS 0.00808f
C74 B.n40 VSUBS 0.00808f
C75 B.n41 VSUBS 0.018678f
C76 B.n42 VSUBS 0.00808f
C77 B.n43 VSUBS 0.00808f
C78 B.n44 VSUBS 0.00808f
C79 B.n45 VSUBS 0.00808f
C80 B.n46 VSUBS 0.00808f
C81 B.n47 VSUBS 0.00808f
C82 B.n48 VSUBS 0.00808f
C83 B.n49 VSUBS 0.00808f
C84 B.n50 VSUBS 0.00808f
C85 B.n51 VSUBS 0.00808f
C86 B.n52 VSUBS 0.00808f
C87 B.n53 VSUBS 0.00808f
C88 B.n54 VSUBS 0.00808f
C89 B.n55 VSUBS 0.00808f
C90 B.n56 VSUBS 0.00808f
C91 B.n57 VSUBS 0.00808f
C92 B.n58 VSUBS 0.00808f
C93 B.n59 VSUBS 0.00808f
C94 B.n60 VSUBS 0.00808f
C95 B.n61 VSUBS 0.00808f
C96 B.n62 VSUBS 0.00808f
C97 B.n63 VSUBS 0.00808f
C98 B.n64 VSUBS 0.00808f
C99 B.n65 VSUBS 0.00808f
C100 B.n66 VSUBS 0.00808f
C101 B.n67 VSUBS 0.00808f
C102 B.n68 VSUBS 0.00808f
C103 B.n69 VSUBS 0.00808f
C104 B.n70 VSUBS 0.00808f
C105 B.n71 VSUBS 0.00808f
C106 B.n72 VSUBS 0.00808f
C107 B.n73 VSUBS 0.00808f
C108 B.n74 VSUBS 0.018678f
C109 B.n75 VSUBS 0.00808f
C110 B.n76 VSUBS 0.00808f
C111 B.n77 VSUBS 0.00808f
C112 B.n78 VSUBS 0.00808f
C113 B.n79 VSUBS 0.00808f
C114 B.n80 VSUBS 0.00808f
C115 B.n81 VSUBS 0.00808f
C116 B.t10 VSUBS 0.048262f
C117 B.t11 VSUBS 0.060177f
C118 B.t9 VSUBS 0.252014f
C119 B.n82 VSUBS 0.105412f
C120 B.n83 VSUBS 0.092707f
C121 B.n84 VSUBS 0.00808f
C122 B.n85 VSUBS 0.00808f
C123 B.n86 VSUBS 0.00808f
C124 B.n87 VSUBS 0.00808f
C125 B.t4 VSUBS 0.048261f
C126 B.t5 VSUBS 0.060176f
C127 B.t3 VSUBS 0.252014f
C128 B.n88 VSUBS 0.105412f
C129 B.n89 VSUBS 0.092707f
C130 B.n90 VSUBS 0.018721f
C131 B.n91 VSUBS 0.00808f
C132 B.n92 VSUBS 0.00808f
C133 B.n93 VSUBS 0.00808f
C134 B.n94 VSUBS 0.00808f
C135 B.n95 VSUBS 0.00808f
C136 B.n96 VSUBS 0.00808f
C137 B.n97 VSUBS 0.018678f
C138 B.n98 VSUBS 0.00808f
C139 B.n99 VSUBS 0.00808f
C140 B.n100 VSUBS 0.00808f
C141 B.n101 VSUBS 0.00808f
C142 B.n102 VSUBS 0.00808f
C143 B.n103 VSUBS 0.00808f
C144 B.n104 VSUBS 0.00808f
C145 B.n105 VSUBS 0.00808f
C146 B.n106 VSUBS 0.00808f
C147 B.n107 VSUBS 0.00808f
C148 B.n108 VSUBS 0.00808f
C149 B.n109 VSUBS 0.00808f
C150 B.n110 VSUBS 0.00808f
C151 B.n111 VSUBS 0.00808f
C152 B.n112 VSUBS 0.00808f
C153 B.n113 VSUBS 0.00808f
C154 B.n114 VSUBS 0.00808f
C155 B.n115 VSUBS 0.00808f
C156 B.n116 VSUBS 0.00808f
C157 B.n117 VSUBS 0.00808f
C158 B.n118 VSUBS 0.00808f
C159 B.n119 VSUBS 0.00808f
C160 B.n120 VSUBS 0.00808f
C161 B.n121 VSUBS 0.00808f
C162 B.n122 VSUBS 0.00808f
C163 B.n123 VSUBS 0.00808f
C164 B.n124 VSUBS 0.00808f
C165 B.n125 VSUBS 0.00808f
C166 B.n126 VSUBS 0.00808f
C167 B.n127 VSUBS 0.00808f
C168 B.n128 VSUBS 0.00808f
C169 B.n129 VSUBS 0.00808f
C170 B.n130 VSUBS 0.00808f
C171 B.n131 VSUBS 0.00808f
C172 B.n132 VSUBS 0.00808f
C173 B.n133 VSUBS 0.00808f
C174 B.n134 VSUBS 0.00808f
C175 B.n135 VSUBS 0.00808f
C176 B.n136 VSUBS 0.00808f
C177 B.n137 VSUBS 0.00808f
C178 B.n138 VSUBS 0.00808f
C179 B.n139 VSUBS 0.00808f
C180 B.n140 VSUBS 0.00808f
C181 B.n141 VSUBS 0.00808f
C182 B.n142 VSUBS 0.00808f
C183 B.n143 VSUBS 0.00808f
C184 B.n144 VSUBS 0.00808f
C185 B.n145 VSUBS 0.00808f
C186 B.n146 VSUBS 0.00808f
C187 B.n147 VSUBS 0.00808f
C188 B.n148 VSUBS 0.00808f
C189 B.n149 VSUBS 0.00808f
C190 B.n150 VSUBS 0.00808f
C191 B.n151 VSUBS 0.00808f
C192 B.n152 VSUBS 0.00808f
C193 B.n153 VSUBS 0.00808f
C194 B.n154 VSUBS 0.00808f
C195 B.n155 VSUBS 0.00808f
C196 B.n156 VSUBS 0.00808f
C197 B.n157 VSUBS 0.00808f
C198 B.n158 VSUBS 0.01792f
C199 B.n159 VSUBS 0.01792f
C200 B.n160 VSUBS 0.018678f
C201 B.n161 VSUBS 0.00808f
C202 B.n162 VSUBS 0.00808f
C203 B.n163 VSUBS 0.00808f
C204 B.n164 VSUBS 0.00808f
C205 B.n165 VSUBS 0.00808f
C206 B.n166 VSUBS 0.00808f
C207 B.n167 VSUBS 0.00808f
C208 B.n168 VSUBS 0.00808f
C209 B.n169 VSUBS 0.00808f
C210 B.n170 VSUBS 0.00808f
C211 B.n171 VSUBS 0.00808f
C212 B.n172 VSUBS 0.00808f
C213 B.n173 VSUBS 0.00808f
C214 B.n174 VSUBS 0.00808f
C215 B.n175 VSUBS 0.00808f
C216 B.n176 VSUBS 0.00808f
C217 B.n177 VSUBS 0.00808f
C218 B.n178 VSUBS 0.00808f
C219 B.n179 VSUBS 0.007605f
C220 B.n180 VSUBS 0.00808f
C221 B.n181 VSUBS 0.00808f
C222 B.n182 VSUBS 0.004515f
C223 B.n183 VSUBS 0.00808f
C224 B.n184 VSUBS 0.00808f
C225 B.n185 VSUBS 0.00808f
C226 B.n186 VSUBS 0.00808f
C227 B.n187 VSUBS 0.00808f
C228 B.n188 VSUBS 0.00808f
C229 B.n189 VSUBS 0.00808f
C230 B.n190 VSUBS 0.00808f
C231 B.n191 VSUBS 0.00808f
C232 B.n192 VSUBS 0.00808f
C233 B.n193 VSUBS 0.00808f
C234 B.n194 VSUBS 0.00808f
C235 B.n195 VSUBS 0.004515f
C236 B.n196 VSUBS 0.018721f
C237 B.n197 VSUBS 0.007605f
C238 B.n198 VSUBS 0.00808f
C239 B.n199 VSUBS 0.00808f
C240 B.n200 VSUBS 0.00808f
C241 B.n201 VSUBS 0.00808f
C242 B.n202 VSUBS 0.00808f
C243 B.n203 VSUBS 0.00808f
C244 B.n204 VSUBS 0.00808f
C245 B.n205 VSUBS 0.00808f
C246 B.n206 VSUBS 0.00808f
C247 B.n207 VSUBS 0.00808f
C248 B.n208 VSUBS 0.00808f
C249 B.n209 VSUBS 0.00808f
C250 B.n210 VSUBS 0.00808f
C251 B.n211 VSUBS 0.00808f
C252 B.n212 VSUBS 0.00808f
C253 B.n213 VSUBS 0.00808f
C254 B.n214 VSUBS 0.00808f
C255 B.n215 VSUBS 0.00808f
C256 B.n216 VSUBS 0.00808f
C257 B.n217 VSUBS 0.018678f
C258 B.n218 VSUBS 0.01792f
C259 B.n219 VSUBS 0.01792f
C260 B.n220 VSUBS 0.00808f
C261 B.n221 VSUBS 0.00808f
C262 B.n222 VSUBS 0.00808f
C263 B.n223 VSUBS 0.00808f
C264 B.n224 VSUBS 0.00808f
C265 B.n225 VSUBS 0.00808f
C266 B.n226 VSUBS 0.00808f
C267 B.n227 VSUBS 0.00808f
C268 B.n228 VSUBS 0.00808f
C269 B.n229 VSUBS 0.00808f
C270 B.n230 VSUBS 0.00808f
C271 B.n231 VSUBS 0.00808f
C272 B.n232 VSUBS 0.00808f
C273 B.n233 VSUBS 0.00808f
C274 B.n234 VSUBS 0.00808f
C275 B.n235 VSUBS 0.00808f
C276 B.n236 VSUBS 0.00808f
C277 B.n237 VSUBS 0.00808f
C278 B.n238 VSUBS 0.00808f
C279 B.n239 VSUBS 0.00808f
C280 B.n240 VSUBS 0.00808f
C281 B.n241 VSUBS 0.00808f
C282 B.n242 VSUBS 0.00808f
C283 B.n243 VSUBS 0.00808f
C284 B.n244 VSUBS 0.00808f
C285 B.n245 VSUBS 0.00808f
C286 B.n246 VSUBS 0.00808f
C287 B.n247 VSUBS 0.00808f
C288 B.n248 VSUBS 0.00808f
C289 B.n249 VSUBS 0.00808f
C290 B.n250 VSUBS 0.00808f
C291 B.n251 VSUBS 0.00808f
C292 B.n252 VSUBS 0.00808f
C293 B.n253 VSUBS 0.00808f
C294 B.n254 VSUBS 0.00808f
C295 B.n255 VSUBS 0.00808f
C296 B.n256 VSUBS 0.00808f
C297 B.n257 VSUBS 0.00808f
C298 B.n258 VSUBS 0.00808f
C299 B.n259 VSUBS 0.00808f
C300 B.n260 VSUBS 0.00808f
C301 B.n261 VSUBS 0.00808f
C302 B.n262 VSUBS 0.00808f
C303 B.n263 VSUBS 0.00808f
C304 B.n264 VSUBS 0.00808f
C305 B.n265 VSUBS 0.00808f
C306 B.n266 VSUBS 0.00808f
C307 B.n267 VSUBS 0.00808f
C308 B.n268 VSUBS 0.00808f
C309 B.n269 VSUBS 0.00808f
C310 B.n270 VSUBS 0.00808f
C311 B.n271 VSUBS 0.00808f
C312 B.n272 VSUBS 0.00808f
C313 B.n273 VSUBS 0.00808f
C314 B.n274 VSUBS 0.00808f
C315 B.n275 VSUBS 0.00808f
C316 B.n276 VSUBS 0.00808f
C317 B.n277 VSUBS 0.00808f
C318 B.n278 VSUBS 0.00808f
C319 B.n279 VSUBS 0.00808f
C320 B.n280 VSUBS 0.00808f
C321 B.n281 VSUBS 0.00808f
C322 B.n282 VSUBS 0.00808f
C323 B.n283 VSUBS 0.00808f
C324 B.n284 VSUBS 0.00808f
C325 B.n285 VSUBS 0.00808f
C326 B.n286 VSUBS 0.00808f
C327 B.n287 VSUBS 0.00808f
C328 B.n288 VSUBS 0.00808f
C329 B.n289 VSUBS 0.00808f
C330 B.n290 VSUBS 0.00808f
C331 B.n291 VSUBS 0.00808f
C332 B.n292 VSUBS 0.00808f
C333 B.n293 VSUBS 0.00808f
C334 B.n294 VSUBS 0.00808f
C335 B.n295 VSUBS 0.00808f
C336 B.n296 VSUBS 0.00808f
C337 B.n297 VSUBS 0.00808f
C338 B.n298 VSUBS 0.00808f
C339 B.n299 VSUBS 0.00808f
C340 B.n300 VSUBS 0.00808f
C341 B.n301 VSUBS 0.00808f
C342 B.n302 VSUBS 0.00808f
C343 B.n303 VSUBS 0.00808f
C344 B.n304 VSUBS 0.00808f
C345 B.n305 VSUBS 0.00808f
C346 B.n306 VSUBS 0.00808f
C347 B.n307 VSUBS 0.00808f
C348 B.n308 VSUBS 0.00808f
C349 B.n309 VSUBS 0.00808f
C350 B.n310 VSUBS 0.00808f
C351 B.n311 VSUBS 0.00808f
C352 B.n312 VSUBS 0.00808f
C353 B.n313 VSUBS 0.00808f
C354 B.n314 VSUBS 0.01792f
C355 B.n315 VSUBS 0.018923f
C356 B.n316 VSUBS 0.017675f
C357 B.n317 VSUBS 0.00808f
C358 B.n318 VSUBS 0.00808f
C359 B.n319 VSUBS 0.00808f
C360 B.n320 VSUBS 0.00808f
C361 B.n321 VSUBS 0.00808f
C362 B.n322 VSUBS 0.00808f
C363 B.n323 VSUBS 0.00808f
C364 B.n324 VSUBS 0.00808f
C365 B.n325 VSUBS 0.00808f
C366 B.n326 VSUBS 0.00808f
C367 B.n327 VSUBS 0.00808f
C368 B.n328 VSUBS 0.00808f
C369 B.n329 VSUBS 0.00808f
C370 B.n330 VSUBS 0.00808f
C371 B.n331 VSUBS 0.00808f
C372 B.n332 VSUBS 0.00808f
C373 B.n333 VSUBS 0.00808f
C374 B.n334 VSUBS 0.00808f
C375 B.n335 VSUBS 0.007605f
C376 B.n336 VSUBS 0.00808f
C377 B.n337 VSUBS 0.00808f
C378 B.n338 VSUBS 0.004515f
C379 B.n339 VSUBS 0.00808f
C380 B.n340 VSUBS 0.00808f
C381 B.n341 VSUBS 0.00808f
C382 B.n342 VSUBS 0.00808f
C383 B.n343 VSUBS 0.00808f
C384 B.n344 VSUBS 0.00808f
C385 B.n345 VSUBS 0.00808f
C386 B.n346 VSUBS 0.00808f
C387 B.n347 VSUBS 0.00808f
C388 B.n348 VSUBS 0.00808f
C389 B.n349 VSUBS 0.00808f
C390 B.n350 VSUBS 0.00808f
C391 B.n351 VSUBS 0.004515f
C392 B.n352 VSUBS 0.018721f
C393 B.n353 VSUBS 0.007605f
C394 B.n354 VSUBS 0.00808f
C395 B.n355 VSUBS 0.00808f
C396 B.n356 VSUBS 0.00808f
C397 B.n357 VSUBS 0.00808f
C398 B.n358 VSUBS 0.00808f
C399 B.n359 VSUBS 0.00808f
C400 B.n360 VSUBS 0.00808f
C401 B.n361 VSUBS 0.00808f
C402 B.n362 VSUBS 0.00808f
C403 B.n363 VSUBS 0.00808f
C404 B.n364 VSUBS 0.00808f
C405 B.n365 VSUBS 0.00808f
C406 B.n366 VSUBS 0.00808f
C407 B.n367 VSUBS 0.00808f
C408 B.n368 VSUBS 0.00808f
C409 B.n369 VSUBS 0.00808f
C410 B.n370 VSUBS 0.00808f
C411 B.n371 VSUBS 0.00808f
C412 B.n372 VSUBS 0.00808f
C413 B.n373 VSUBS 0.018678f
C414 B.n374 VSUBS 0.01792f
C415 B.n375 VSUBS 0.01792f
C416 B.n376 VSUBS 0.00808f
C417 B.n377 VSUBS 0.00808f
C418 B.n378 VSUBS 0.00808f
C419 B.n379 VSUBS 0.00808f
C420 B.n380 VSUBS 0.00808f
C421 B.n381 VSUBS 0.00808f
C422 B.n382 VSUBS 0.00808f
C423 B.n383 VSUBS 0.00808f
C424 B.n384 VSUBS 0.00808f
C425 B.n385 VSUBS 0.00808f
C426 B.n386 VSUBS 0.00808f
C427 B.n387 VSUBS 0.00808f
C428 B.n388 VSUBS 0.00808f
C429 B.n389 VSUBS 0.00808f
C430 B.n390 VSUBS 0.00808f
C431 B.n391 VSUBS 0.00808f
C432 B.n392 VSUBS 0.00808f
C433 B.n393 VSUBS 0.00808f
C434 B.n394 VSUBS 0.00808f
C435 B.n395 VSUBS 0.00808f
C436 B.n396 VSUBS 0.00808f
C437 B.n397 VSUBS 0.00808f
C438 B.n398 VSUBS 0.00808f
C439 B.n399 VSUBS 0.00808f
C440 B.n400 VSUBS 0.00808f
C441 B.n401 VSUBS 0.00808f
C442 B.n402 VSUBS 0.00808f
C443 B.n403 VSUBS 0.00808f
C444 B.n404 VSUBS 0.00808f
C445 B.n405 VSUBS 0.00808f
C446 B.n406 VSUBS 0.00808f
C447 B.n407 VSUBS 0.00808f
C448 B.n408 VSUBS 0.00808f
C449 B.n409 VSUBS 0.00808f
C450 B.n410 VSUBS 0.00808f
C451 B.n411 VSUBS 0.00808f
C452 B.n412 VSUBS 0.00808f
C453 B.n413 VSUBS 0.00808f
C454 B.n414 VSUBS 0.00808f
C455 B.n415 VSUBS 0.00808f
C456 B.n416 VSUBS 0.00808f
C457 B.n417 VSUBS 0.00808f
C458 B.n418 VSUBS 0.00808f
C459 B.n419 VSUBS 0.00808f
C460 B.n420 VSUBS 0.00808f
C461 B.n421 VSUBS 0.00808f
C462 B.n422 VSUBS 0.00808f
C463 B.n423 VSUBS 0.018296f
C464 VDD2.n0 VSUBS 0.017985f
C465 VDD2.n1 VSUBS 0.130001f
C466 VDD2.n2 VSUBS 0.008564f
C467 VDD2.t5 VSUBS 0.047451f
C468 VDD2.n3 VSUBS 0.057109f
C469 VDD2.n4 VSUBS 0.014354f
C470 VDD2.n5 VSUBS 0.015181f
C471 VDD2.n6 VSUBS 0.050617f
C472 VDD2.n7 VSUBS 0.009068f
C473 VDD2.n8 VSUBS 0.008564f
C474 VDD2.n9 VSUBS 0.035096f
C475 VDD2.n10 VSUBS 0.038917f
C476 VDD2.t4 VSUBS 0.033752f
C477 VDD2.t1 VSUBS 0.033752f
C478 VDD2.n11 VSUBS 0.162413f
C479 VDD2.n12 VSUBS 1.17284f
C480 VDD2.n13 VSUBS 0.017985f
C481 VDD2.n14 VSUBS 0.130001f
C482 VDD2.n15 VSUBS 0.008564f
C483 VDD2.t2 VSUBS 0.047451f
C484 VDD2.n16 VSUBS 0.057109f
C485 VDD2.n17 VSUBS 0.014354f
C486 VDD2.n18 VSUBS 0.015181f
C487 VDD2.n19 VSUBS 0.050617f
C488 VDD2.n20 VSUBS 0.009068f
C489 VDD2.n21 VSUBS 0.008564f
C490 VDD2.n22 VSUBS 0.035096f
C491 VDD2.n23 VSUBS 0.036491f
C492 VDD2.n24 VSUBS 1.00001f
C493 VDD2.t0 VSUBS 0.033752f
C494 VDD2.t3 VSUBS 0.033752f
C495 VDD2.n25 VSUBS 0.162405f
C496 VN.n0 VSUBS 0.048789f
C497 VN.t4 VSUBS 0.542253f
C498 VN.n1 VSUBS 0.039544f
C499 VN.t0 VSUBS 0.760313f
C500 VN.n2 VSUBS 0.339264f
C501 VN.t1 VSUBS 0.542253f
C502 VN.n3 VSUBS 0.380497f
C503 VN.n4 VSUBS 0.097949f
C504 VN.n5 VSUBS 0.352842f
C505 VN.n6 VSUBS 0.048789f
C506 VN.n7 VSUBS 0.048789f
C507 VN.n8 VSUBS 0.09696f
C508 VN.n9 VSUBS 0.04807f
C509 VN.n10 VSUBS 0.347921f
C510 VN.n11 VSUBS 0.051773f
C511 VN.n12 VSUBS 0.048789f
C512 VN.t3 VSUBS 0.542253f
C513 VN.n13 VSUBS 0.039544f
C514 VN.t2 VSUBS 0.760313f
C515 VN.n14 VSUBS 0.339264f
C516 VN.t5 VSUBS 0.542253f
C517 VN.n15 VSUBS 0.380497f
C518 VN.n16 VSUBS 0.097949f
C519 VN.n17 VSUBS 0.352842f
C520 VN.n18 VSUBS 0.048789f
C521 VN.n19 VSUBS 0.048789f
C522 VN.n20 VSUBS 0.09696f
C523 VN.n21 VSUBS 0.04807f
C524 VN.n22 VSUBS 0.347921f
C525 VN.n23 VSUBS 1.73063f
C526 VDD1.n0 VSUBS 0.017264f
C527 VDD1.n1 VSUBS 0.124785f
C528 VDD1.n2 VSUBS 0.00822f
C529 VDD1.t4 VSUBS 0.045547f
C530 VDD1.n3 VSUBS 0.054818f
C531 VDD1.n4 VSUBS 0.013778f
C532 VDD1.n5 VSUBS 0.014572f
C533 VDD1.n6 VSUBS 0.048586f
C534 VDD1.n7 VSUBS 0.008704f
C535 VDD1.n8 VSUBS 0.00822f
C536 VDD1.n9 VSUBS 0.033687f
C537 VDD1.n10 VSUBS 0.03771f
C538 VDD1.n11 VSUBS 0.017264f
C539 VDD1.n12 VSUBS 0.124785f
C540 VDD1.n13 VSUBS 0.00822f
C541 VDD1.t0 VSUBS 0.045547f
C542 VDD1.n14 VSUBS 0.054818f
C543 VDD1.n15 VSUBS 0.013778f
C544 VDD1.n16 VSUBS 0.014572f
C545 VDD1.n17 VSUBS 0.048586f
C546 VDD1.n18 VSUBS 0.008704f
C547 VDD1.n19 VSUBS 0.00822f
C548 VDD1.n20 VSUBS 0.033687f
C549 VDD1.n21 VSUBS 0.037355f
C550 VDD1.t1 VSUBS 0.032397f
C551 VDD1.t2 VSUBS 0.032397f
C552 VDD1.n22 VSUBS 0.155896f
C553 VDD1.n23 VSUBS 1.18282f
C554 VDD1.t3 VSUBS 0.032397f
C555 VDD1.t5 VSUBS 0.032397f
C556 VDD1.n24 VSUBS 0.155137f
C557 VDD1.n25 VSUBS 1.16624f
C558 VTAIL.t5 VSUBS 0.065049f
C559 VTAIL.t0 VSUBS 0.065049f
C560 VTAIL.n0 VSUBS 0.264538f
C561 VTAIL.n1 VSUBS 0.572341f
C562 VTAIL.n2 VSUBS 0.034663f
C563 VTAIL.n3 VSUBS 0.250551f
C564 VTAIL.n4 VSUBS 0.016505f
C565 VTAIL.t9 VSUBS 0.091452f
C566 VTAIL.n5 VSUBS 0.110066f
C567 VTAIL.n6 VSUBS 0.027665f
C568 VTAIL.n7 VSUBS 0.029259f
C569 VTAIL.n8 VSUBS 0.097554f
C570 VTAIL.n9 VSUBS 0.017476f
C571 VTAIL.n10 VSUBS 0.016505f
C572 VTAIL.n11 VSUBS 0.06764f
C573 VTAIL.n12 VSUBS 0.049092f
C574 VTAIL.n13 VSUBS 0.32936f
C575 VTAIL.t11 VSUBS 0.065049f
C576 VTAIL.t10 VSUBS 0.065049f
C577 VTAIL.n14 VSUBS 0.264538f
C578 VTAIL.n15 VSUBS 1.55375f
C579 VTAIL.t4 VSUBS 0.065049f
C580 VTAIL.t1 VSUBS 0.065049f
C581 VTAIL.n16 VSUBS 0.264539f
C582 VTAIL.n17 VSUBS 1.55375f
C583 VTAIL.n18 VSUBS 0.034663f
C584 VTAIL.n19 VSUBS 0.250551f
C585 VTAIL.n20 VSUBS 0.016505f
C586 VTAIL.t3 VSUBS 0.091452f
C587 VTAIL.n21 VSUBS 0.110066f
C588 VTAIL.n22 VSUBS 0.027665f
C589 VTAIL.n23 VSUBS 0.029259f
C590 VTAIL.n24 VSUBS 0.097554f
C591 VTAIL.n25 VSUBS 0.017476f
C592 VTAIL.n26 VSUBS 0.016505f
C593 VTAIL.n27 VSUBS 0.06764f
C594 VTAIL.n28 VSUBS 0.049092f
C595 VTAIL.n29 VSUBS 0.32936f
C596 VTAIL.t7 VSUBS 0.065049f
C597 VTAIL.t8 VSUBS 0.065049f
C598 VTAIL.n30 VSUBS 0.264539f
C599 VTAIL.n31 VSUBS 0.695841f
C600 VTAIL.n32 VSUBS 0.034663f
C601 VTAIL.n33 VSUBS 0.250551f
C602 VTAIL.n34 VSUBS 0.016505f
C603 VTAIL.t6 VSUBS 0.091452f
C604 VTAIL.n35 VSUBS 0.110066f
C605 VTAIL.n36 VSUBS 0.027665f
C606 VTAIL.n37 VSUBS 0.029259f
C607 VTAIL.n38 VSUBS 0.097554f
C608 VTAIL.n39 VSUBS 0.017476f
C609 VTAIL.n40 VSUBS 0.016505f
C610 VTAIL.n41 VSUBS 0.06764f
C611 VTAIL.n42 VSUBS 0.049092f
C612 VTAIL.n43 VSUBS 1.01492f
C613 VTAIL.n44 VSUBS 0.034663f
C614 VTAIL.n45 VSUBS 0.250551f
C615 VTAIL.n46 VSUBS 0.016505f
C616 VTAIL.t2 VSUBS 0.091452f
C617 VTAIL.n47 VSUBS 0.110066f
C618 VTAIL.n48 VSUBS 0.027665f
C619 VTAIL.n49 VSUBS 0.029259f
C620 VTAIL.n50 VSUBS 0.097554f
C621 VTAIL.n51 VSUBS 0.017476f
C622 VTAIL.n52 VSUBS 0.016505f
C623 VTAIL.n53 VSUBS 0.06764f
C624 VTAIL.n54 VSUBS 0.049092f
C625 VTAIL.n55 VSUBS 0.966075f
C626 VP.n0 VSUBS 0.0509f
C627 VP.t3 VSUBS 0.565712f
C628 VP.n1 VSUBS 0.041255f
C629 VP.n2 VSUBS 0.0509f
C630 VP.t4 VSUBS 0.565712f
C631 VP.n3 VSUBS 0.041255f
C632 VP.n4 VSUBS 0.0509f
C633 VP.t5 VSUBS 0.565712f
C634 VP.n5 VSUBS 0.0509f
C635 VP.t0 VSUBS 0.565712f
C636 VP.n6 VSUBS 0.041255f
C637 VP.t1 VSUBS 0.793206f
C638 VP.n7 VSUBS 0.353941f
C639 VP.t2 VSUBS 0.565712f
C640 VP.n8 VSUBS 0.396958f
C641 VP.n9 VSUBS 0.102186f
C642 VP.n10 VSUBS 0.368107f
C643 VP.n11 VSUBS 0.0509f
C644 VP.n12 VSUBS 0.0509f
C645 VP.n13 VSUBS 0.101155f
C646 VP.n14 VSUBS 0.05015f
C647 VP.n15 VSUBS 0.362973f
C648 VP.n16 VSUBS 1.77186f
C649 VP.n17 VSUBS 1.82003f
C650 VP.n18 VSUBS 0.362973f
C651 VP.n19 VSUBS 0.05015f
C652 VP.n20 VSUBS 0.101155f
C653 VP.n21 VSUBS 0.0509f
C654 VP.n22 VSUBS 0.0509f
C655 VP.n23 VSUBS 0.0509f
C656 VP.n24 VSUBS 0.102186f
C657 VP.n25 VSUBS 0.310696f
C658 VP.n26 VSUBS 0.102186f
C659 VP.n27 VSUBS 0.0509f
C660 VP.n28 VSUBS 0.0509f
C661 VP.n29 VSUBS 0.0509f
C662 VP.n30 VSUBS 0.101155f
C663 VP.n31 VSUBS 0.05015f
C664 VP.n32 VSUBS 0.362973f
C665 VP.n33 VSUBS 0.054013f
.ends

