* NGSPICE file created from diff_pair_sample_0012.ext - technology: sky130A

.subckt diff_pair_sample_0012 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=2.99
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=2.99
X2 VTAIL.t1 VN.t0 VDD2.t5 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=2.99
X3 VDD2.t4 VN.t1 VTAIL.t4 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=2.99
X4 VDD1.t4 VP.t1 VTAIL.t8 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=2.99
X5 VDD2.t3 VN.t2 VTAIL.t0 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=2.99
X6 B.t8 B.t6 B.t7 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=2.99
X7 VDD2.t2 VN.t3 VTAIL.t3 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=2.99
X8 VDD1.t3 VP.t2 VTAIL.t9 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=2.99
X9 VDD2.t1 VN.t4 VTAIL.t11 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=2.99
X10 VTAIL.t6 VP.t3 VDD1.t2 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=2.99
X11 VTAIL.t7 VP.t4 VDD1.t1 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=2.99
X12 B.t5 B.t3 B.t4 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=2.99
X13 VDD1.t0 VP.t5 VTAIL.t10 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=2.99
X14 VTAIL.t2 VN.t5 VDD2.t0 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=2.99
X15 B.t2 B.t0 B.t1 w_n3626_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=2.99
R0 B.n646 B.n95 585
R1 B.n648 B.n647 585
R2 B.n649 B.n94 585
R3 B.n651 B.n650 585
R4 B.n652 B.n93 585
R5 B.n654 B.n653 585
R6 B.n655 B.n92 585
R7 B.n657 B.n656 585
R8 B.n658 B.n91 585
R9 B.n660 B.n659 585
R10 B.n661 B.n90 585
R11 B.n663 B.n662 585
R12 B.n664 B.n89 585
R13 B.n666 B.n665 585
R14 B.n667 B.n88 585
R15 B.n669 B.n668 585
R16 B.n670 B.n87 585
R17 B.n672 B.n671 585
R18 B.n673 B.n86 585
R19 B.n675 B.n674 585
R20 B.n676 B.n85 585
R21 B.n678 B.n677 585
R22 B.n679 B.n84 585
R23 B.n681 B.n680 585
R24 B.n682 B.n83 585
R25 B.n684 B.n683 585
R26 B.n685 B.n82 585
R27 B.n687 B.n686 585
R28 B.n688 B.n81 585
R29 B.n690 B.n689 585
R30 B.n691 B.n80 585
R31 B.n693 B.n692 585
R32 B.n694 B.n79 585
R33 B.n696 B.n695 585
R34 B.n697 B.n78 585
R35 B.n699 B.n698 585
R36 B.n700 B.n77 585
R37 B.n702 B.n701 585
R38 B.n703 B.n76 585
R39 B.n705 B.n704 585
R40 B.n706 B.n75 585
R41 B.n708 B.n707 585
R42 B.n709 B.n74 585
R43 B.n711 B.n710 585
R44 B.n712 B.n73 585
R45 B.n714 B.n713 585
R46 B.n715 B.n72 585
R47 B.n717 B.n716 585
R48 B.n718 B.n71 585
R49 B.n720 B.n719 585
R50 B.n721 B.n70 585
R51 B.n723 B.n722 585
R52 B.n724 B.n69 585
R53 B.n726 B.n725 585
R54 B.n727 B.n68 585
R55 B.n729 B.n728 585
R56 B.n730 B.n67 585
R57 B.n732 B.n731 585
R58 B.n733 B.n66 585
R59 B.n735 B.n734 585
R60 B.n736 B.n63 585
R61 B.n739 B.n738 585
R62 B.n740 B.n62 585
R63 B.n742 B.n741 585
R64 B.n743 B.n61 585
R65 B.n745 B.n744 585
R66 B.n746 B.n60 585
R67 B.n748 B.n747 585
R68 B.n749 B.n59 585
R69 B.n751 B.n750 585
R70 B.n753 B.n752 585
R71 B.n754 B.n55 585
R72 B.n756 B.n755 585
R73 B.n757 B.n54 585
R74 B.n759 B.n758 585
R75 B.n760 B.n53 585
R76 B.n762 B.n761 585
R77 B.n763 B.n52 585
R78 B.n765 B.n764 585
R79 B.n766 B.n51 585
R80 B.n768 B.n767 585
R81 B.n769 B.n50 585
R82 B.n771 B.n770 585
R83 B.n772 B.n49 585
R84 B.n774 B.n773 585
R85 B.n775 B.n48 585
R86 B.n777 B.n776 585
R87 B.n778 B.n47 585
R88 B.n780 B.n779 585
R89 B.n781 B.n46 585
R90 B.n783 B.n782 585
R91 B.n784 B.n45 585
R92 B.n786 B.n785 585
R93 B.n787 B.n44 585
R94 B.n789 B.n788 585
R95 B.n790 B.n43 585
R96 B.n792 B.n791 585
R97 B.n793 B.n42 585
R98 B.n795 B.n794 585
R99 B.n796 B.n41 585
R100 B.n798 B.n797 585
R101 B.n799 B.n40 585
R102 B.n801 B.n800 585
R103 B.n802 B.n39 585
R104 B.n804 B.n803 585
R105 B.n805 B.n38 585
R106 B.n807 B.n806 585
R107 B.n808 B.n37 585
R108 B.n810 B.n809 585
R109 B.n811 B.n36 585
R110 B.n813 B.n812 585
R111 B.n814 B.n35 585
R112 B.n816 B.n815 585
R113 B.n817 B.n34 585
R114 B.n819 B.n818 585
R115 B.n820 B.n33 585
R116 B.n822 B.n821 585
R117 B.n823 B.n32 585
R118 B.n825 B.n824 585
R119 B.n826 B.n31 585
R120 B.n828 B.n827 585
R121 B.n829 B.n30 585
R122 B.n831 B.n830 585
R123 B.n832 B.n29 585
R124 B.n834 B.n833 585
R125 B.n835 B.n28 585
R126 B.n837 B.n836 585
R127 B.n838 B.n27 585
R128 B.n840 B.n839 585
R129 B.n841 B.n26 585
R130 B.n843 B.n842 585
R131 B.n645 B.n644 585
R132 B.n643 B.n96 585
R133 B.n642 B.n641 585
R134 B.n640 B.n97 585
R135 B.n639 B.n638 585
R136 B.n637 B.n98 585
R137 B.n636 B.n635 585
R138 B.n634 B.n99 585
R139 B.n633 B.n632 585
R140 B.n631 B.n100 585
R141 B.n630 B.n629 585
R142 B.n628 B.n101 585
R143 B.n627 B.n626 585
R144 B.n625 B.n102 585
R145 B.n624 B.n623 585
R146 B.n622 B.n103 585
R147 B.n621 B.n620 585
R148 B.n619 B.n104 585
R149 B.n618 B.n617 585
R150 B.n616 B.n105 585
R151 B.n615 B.n614 585
R152 B.n613 B.n106 585
R153 B.n612 B.n611 585
R154 B.n610 B.n107 585
R155 B.n609 B.n608 585
R156 B.n607 B.n108 585
R157 B.n606 B.n605 585
R158 B.n604 B.n109 585
R159 B.n603 B.n602 585
R160 B.n601 B.n110 585
R161 B.n600 B.n599 585
R162 B.n598 B.n111 585
R163 B.n597 B.n596 585
R164 B.n595 B.n112 585
R165 B.n594 B.n593 585
R166 B.n592 B.n113 585
R167 B.n591 B.n590 585
R168 B.n589 B.n114 585
R169 B.n588 B.n587 585
R170 B.n586 B.n115 585
R171 B.n585 B.n584 585
R172 B.n583 B.n116 585
R173 B.n582 B.n581 585
R174 B.n580 B.n117 585
R175 B.n579 B.n578 585
R176 B.n577 B.n118 585
R177 B.n576 B.n575 585
R178 B.n574 B.n119 585
R179 B.n573 B.n572 585
R180 B.n571 B.n120 585
R181 B.n570 B.n569 585
R182 B.n568 B.n121 585
R183 B.n567 B.n566 585
R184 B.n565 B.n122 585
R185 B.n564 B.n563 585
R186 B.n562 B.n123 585
R187 B.n561 B.n560 585
R188 B.n559 B.n124 585
R189 B.n558 B.n557 585
R190 B.n556 B.n125 585
R191 B.n555 B.n554 585
R192 B.n553 B.n126 585
R193 B.n552 B.n551 585
R194 B.n550 B.n127 585
R195 B.n549 B.n548 585
R196 B.n547 B.n128 585
R197 B.n546 B.n545 585
R198 B.n544 B.n129 585
R199 B.n543 B.n542 585
R200 B.n541 B.n130 585
R201 B.n540 B.n539 585
R202 B.n538 B.n131 585
R203 B.n537 B.n536 585
R204 B.n535 B.n132 585
R205 B.n534 B.n533 585
R206 B.n532 B.n133 585
R207 B.n531 B.n530 585
R208 B.n529 B.n134 585
R209 B.n528 B.n527 585
R210 B.n526 B.n135 585
R211 B.n525 B.n524 585
R212 B.n523 B.n136 585
R213 B.n522 B.n521 585
R214 B.n520 B.n137 585
R215 B.n519 B.n518 585
R216 B.n517 B.n138 585
R217 B.n516 B.n515 585
R218 B.n514 B.n139 585
R219 B.n513 B.n512 585
R220 B.n511 B.n140 585
R221 B.n510 B.n509 585
R222 B.n508 B.n141 585
R223 B.n507 B.n506 585
R224 B.n505 B.n142 585
R225 B.n504 B.n503 585
R226 B.n306 B.n305 585
R227 B.n307 B.n212 585
R228 B.n309 B.n308 585
R229 B.n310 B.n211 585
R230 B.n312 B.n311 585
R231 B.n313 B.n210 585
R232 B.n315 B.n314 585
R233 B.n316 B.n209 585
R234 B.n318 B.n317 585
R235 B.n319 B.n208 585
R236 B.n321 B.n320 585
R237 B.n322 B.n207 585
R238 B.n324 B.n323 585
R239 B.n325 B.n206 585
R240 B.n327 B.n326 585
R241 B.n328 B.n205 585
R242 B.n330 B.n329 585
R243 B.n331 B.n204 585
R244 B.n333 B.n332 585
R245 B.n334 B.n203 585
R246 B.n336 B.n335 585
R247 B.n337 B.n202 585
R248 B.n339 B.n338 585
R249 B.n340 B.n201 585
R250 B.n342 B.n341 585
R251 B.n343 B.n200 585
R252 B.n345 B.n344 585
R253 B.n346 B.n199 585
R254 B.n348 B.n347 585
R255 B.n349 B.n198 585
R256 B.n351 B.n350 585
R257 B.n352 B.n197 585
R258 B.n354 B.n353 585
R259 B.n355 B.n196 585
R260 B.n357 B.n356 585
R261 B.n358 B.n195 585
R262 B.n360 B.n359 585
R263 B.n361 B.n194 585
R264 B.n363 B.n362 585
R265 B.n364 B.n193 585
R266 B.n366 B.n365 585
R267 B.n367 B.n192 585
R268 B.n369 B.n368 585
R269 B.n370 B.n191 585
R270 B.n372 B.n371 585
R271 B.n373 B.n190 585
R272 B.n375 B.n374 585
R273 B.n376 B.n189 585
R274 B.n378 B.n377 585
R275 B.n379 B.n188 585
R276 B.n381 B.n380 585
R277 B.n382 B.n187 585
R278 B.n384 B.n383 585
R279 B.n385 B.n186 585
R280 B.n387 B.n386 585
R281 B.n388 B.n185 585
R282 B.n390 B.n389 585
R283 B.n391 B.n184 585
R284 B.n393 B.n392 585
R285 B.n394 B.n183 585
R286 B.n396 B.n395 585
R287 B.n398 B.n397 585
R288 B.n399 B.n179 585
R289 B.n401 B.n400 585
R290 B.n402 B.n178 585
R291 B.n404 B.n403 585
R292 B.n405 B.n177 585
R293 B.n407 B.n406 585
R294 B.n408 B.n176 585
R295 B.n410 B.n409 585
R296 B.n412 B.n173 585
R297 B.n414 B.n413 585
R298 B.n415 B.n172 585
R299 B.n417 B.n416 585
R300 B.n418 B.n171 585
R301 B.n420 B.n419 585
R302 B.n421 B.n170 585
R303 B.n423 B.n422 585
R304 B.n424 B.n169 585
R305 B.n426 B.n425 585
R306 B.n427 B.n168 585
R307 B.n429 B.n428 585
R308 B.n430 B.n167 585
R309 B.n432 B.n431 585
R310 B.n433 B.n166 585
R311 B.n435 B.n434 585
R312 B.n436 B.n165 585
R313 B.n438 B.n437 585
R314 B.n439 B.n164 585
R315 B.n441 B.n440 585
R316 B.n442 B.n163 585
R317 B.n444 B.n443 585
R318 B.n445 B.n162 585
R319 B.n447 B.n446 585
R320 B.n448 B.n161 585
R321 B.n450 B.n449 585
R322 B.n451 B.n160 585
R323 B.n453 B.n452 585
R324 B.n454 B.n159 585
R325 B.n456 B.n455 585
R326 B.n457 B.n158 585
R327 B.n459 B.n458 585
R328 B.n460 B.n157 585
R329 B.n462 B.n461 585
R330 B.n463 B.n156 585
R331 B.n465 B.n464 585
R332 B.n466 B.n155 585
R333 B.n468 B.n467 585
R334 B.n469 B.n154 585
R335 B.n471 B.n470 585
R336 B.n472 B.n153 585
R337 B.n474 B.n473 585
R338 B.n475 B.n152 585
R339 B.n477 B.n476 585
R340 B.n478 B.n151 585
R341 B.n480 B.n479 585
R342 B.n481 B.n150 585
R343 B.n483 B.n482 585
R344 B.n484 B.n149 585
R345 B.n486 B.n485 585
R346 B.n487 B.n148 585
R347 B.n489 B.n488 585
R348 B.n490 B.n147 585
R349 B.n492 B.n491 585
R350 B.n493 B.n146 585
R351 B.n495 B.n494 585
R352 B.n496 B.n145 585
R353 B.n498 B.n497 585
R354 B.n499 B.n144 585
R355 B.n501 B.n500 585
R356 B.n502 B.n143 585
R357 B.n304 B.n213 585
R358 B.n303 B.n302 585
R359 B.n301 B.n214 585
R360 B.n300 B.n299 585
R361 B.n298 B.n215 585
R362 B.n297 B.n296 585
R363 B.n295 B.n216 585
R364 B.n294 B.n293 585
R365 B.n292 B.n217 585
R366 B.n291 B.n290 585
R367 B.n289 B.n218 585
R368 B.n288 B.n287 585
R369 B.n286 B.n219 585
R370 B.n285 B.n284 585
R371 B.n283 B.n220 585
R372 B.n282 B.n281 585
R373 B.n280 B.n221 585
R374 B.n279 B.n278 585
R375 B.n277 B.n222 585
R376 B.n276 B.n275 585
R377 B.n274 B.n223 585
R378 B.n273 B.n272 585
R379 B.n271 B.n224 585
R380 B.n270 B.n269 585
R381 B.n268 B.n225 585
R382 B.n267 B.n266 585
R383 B.n265 B.n226 585
R384 B.n264 B.n263 585
R385 B.n262 B.n227 585
R386 B.n261 B.n260 585
R387 B.n259 B.n228 585
R388 B.n258 B.n257 585
R389 B.n256 B.n229 585
R390 B.n255 B.n254 585
R391 B.n253 B.n230 585
R392 B.n252 B.n251 585
R393 B.n250 B.n231 585
R394 B.n249 B.n248 585
R395 B.n247 B.n232 585
R396 B.n246 B.n245 585
R397 B.n244 B.n233 585
R398 B.n243 B.n242 585
R399 B.n241 B.n234 585
R400 B.n240 B.n239 585
R401 B.n238 B.n235 585
R402 B.n237 B.n236 585
R403 B.n2 B.n0 585
R404 B.n913 B.n1 585
R405 B.n912 B.n911 585
R406 B.n910 B.n3 585
R407 B.n909 B.n908 585
R408 B.n907 B.n4 585
R409 B.n906 B.n905 585
R410 B.n904 B.n5 585
R411 B.n903 B.n902 585
R412 B.n901 B.n6 585
R413 B.n900 B.n899 585
R414 B.n898 B.n7 585
R415 B.n897 B.n896 585
R416 B.n895 B.n8 585
R417 B.n894 B.n893 585
R418 B.n892 B.n9 585
R419 B.n891 B.n890 585
R420 B.n889 B.n10 585
R421 B.n888 B.n887 585
R422 B.n886 B.n11 585
R423 B.n885 B.n884 585
R424 B.n883 B.n12 585
R425 B.n882 B.n881 585
R426 B.n880 B.n13 585
R427 B.n879 B.n878 585
R428 B.n877 B.n14 585
R429 B.n876 B.n875 585
R430 B.n874 B.n15 585
R431 B.n873 B.n872 585
R432 B.n871 B.n16 585
R433 B.n870 B.n869 585
R434 B.n868 B.n17 585
R435 B.n867 B.n866 585
R436 B.n865 B.n18 585
R437 B.n864 B.n863 585
R438 B.n862 B.n19 585
R439 B.n861 B.n860 585
R440 B.n859 B.n20 585
R441 B.n858 B.n857 585
R442 B.n856 B.n21 585
R443 B.n855 B.n854 585
R444 B.n853 B.n22 585
R445 B.n852 B.n851 585
R446 B.n850 B.n23 585
R447 B.n849 B.n848 585
R448 B.n847 B.n24 585
R449 B.n846 B.n845 585
R450 B.n844 B.n25 585
R451 B.n915 B.n914 585
R452 B.n306 B.n213 550.159
R453 B.n842 B.n25 550.159
R454 B.n504 B.n143 550.159
R455 B.n644 B.n95 550.159
R456 B.n174 B.t0 358.005
R457 B.n180 B.t6 358.005
R458 B.n56 B.t9 358.005
R459 B.n64 B.t3 358.005
R460 B.n174 B.t2 174.03
R461 B.n64 B.t4 174.03
R462 B.n180 B.t8 174.006
R463 B.n56 B.t10 174.006
R464 B.n302 B.n213 163.367
R465 B.n302 B.n301 163.367
R466 B.n301 B.n300 163.367
R467 B.n300 B.n215 163.367
R468 B.n296 B.n215 163.367
R469 B.n296 B.n295 163.367
R470 B.n295 B.n294 163.367
R471 B.n294 B.n217 163.367
R472 B.n290 B.n217 163.367
R473 B.n290 B.n289 163.367
R474 B.n289 B.n288 163.367
R475 B.n288 B.n219 163.367
R476 B.n284 B.n219 163.367
R477 B.n284 B.n283 163.367
R478 B.n283 B.n282 163.367
R479 B.n282 B.n221 163.367
R480 B.n278 B.n221 163.367
R481 B.n278 B.n277 163.367
R482 B.n277 B.n276 163.367
R483 B.n276 B.n223 163.367
R484 B.n272 B.n223 163.367
R485 B.n272 B.n271 163.367
R486 B.n271 B.n270 163.367
R487 B.n270 B.n225 163.367
R488 B.n266 B.n225 163.367
R489 B.n266 B.n265 163.367
R490 B.n265 B.n264 163.367
R491 B.n264 B.n227 163.367
R492 B.n260 B.n227 163.367
R493 B.n260 B.n259 163.367
R494 B.n259 B.n258 163.367
R495 B.n258 B.n229 163.367
R496 B.n254 B.n229 163.367
R497 B.n254 B.n253 163.367
R498 B.n253 B.n252 163.367
R499 B.n252 B.n231 163.367
R500 B.n248 B.n231 163.367
R501 B.n248 B.n247 163.367
R502 B.n247 B.n246 163.367
R503 B.n246 B.n233 163.367
R504 B.n242 B.n233 163.367
R505 B.n242 B.n241 163.367
R506 B.n241 B.n240 163.367
R507 B.n240 B.n235 163.367
R508 B.n236 B.n235 163.367
R509 B.n236 B.n2 163.367
R510 B.n914 B.n2 163.367
R511 B.n914 B.n913 163.367
R512 B.n913 B.n912 163.367
R513 B.n912 B.n3 163.367
R514 B.n908 B.n3 163.367
R515 B.n908 B.n907 163.367
R516 B.n907 B.n906 163.367
R517 B.n906 B.n5 163.367
R518 B.n902 B.n5 163.367
R519 B.n902 B.n901 163.367
R520 B.n901 B.n900 163.367
R521 B.n900 B.n7 163.367
R522 B.n896 B.n7 163.367
R523 B.n896 B.n895 163.367
R524 B.n895 B.n894 163.367
R525 B.n894 B.n9 163.367
R526 B.n890 B.n9 163.367
R527 B.n890 B.n889 163.367
R528 B.n889 B.n888 163.367
R529 B.n888 B.n11 163.367
R530 B.n884 B.n11 163.367
R531 B.n884 B.n883 163.367
R532 B.n883 B.n882 163.367
R533 B.n882 B.n13 163.367
R534 B.n878 B.n13 163.367
R535 B.n878 B.n877 163.367
R536 B.n877 B.n876 163.367
R537 B.n876 B.n15 163.367
R538 B.n872 B.n15 163.367
R539 B.n872 B.n871 163.367
R540 B.n871 B.n870 163.367
R541 B.n870 B.n17 163.367
R542 B.n866 B.n17 163.367
R543 B.n866 B.n865 163.367
R544 B.n865 B.n864 163.367
R545 B.n864 B.n19 163.367
R546 B.n860 B.n19 163.367
R547 B.n860 B.n859 163.367
R548 B.n859 B.n858 163.367
R549 B.n858 B.n21 163.367
R550 B.n854 B.n21 163.367
R551 B.n854 B.n853 163.367
R552 B.n853 B.n852 163.367
R553 B.n852 B.n23 163.367
R554 B.n848 B.n23 163.367
R555 B.n848 B.n847 163.367
R556 B.n847 B.n846 163.367
R557 B.n846 B.n25 163.367
R558 B.n307 B.n306 163.367
R559 B.n308 B.n307 163.367
R560 B.n308 B.n211 163.367
R561 B.n312 B.n211 163.367
R562 B.n313 B.n312 163.367
R563 B.n314 B.n313 163.367
R564 B.n314 B.n209 163.367
R565 B.n318 B.n209 163.367
R566 B.n319 B.n318 163.367
R567 B.n320 B.n319 163.367
R568 B.n320 B.n207 163.367
R569 B.n324 B.n207 163.367
R570 B.n325 B.n324 163.367
R571 B.n326 B.n325 163.367
R572 B.n326 B.n205 163.367
R573 B.n330 B.n205 163.367
R574 B.n331 B.n330 163.367
R575 B.n332 B.n331 163.367
R576 B.n332 B.n203 163.367
R577 B.n336 B.n203 163.367
R578 B.n337 B.n336 163.367
R579 B.n338 B.n337 163.367
R580 B.n338 B.n201 163.367
R581 B.n342 B.n201 163.367
R582 B.n343 B.n342 163.367
R583 B.n344 B.n343 163.367
R584 B.n344 B.n199 163.367
R585 B.n348 B.n199 163.367
R586 B.n349 B.n348 163.367
R587 B.n350 B.n349 163.367
R588 B.n350 B.n197 163.367
R589 B.n354 B.n197 163.367
R590 B.n355 B.n354 163.367
R591 B.n356 B.n355 163.367
R592 B.n356 B.n195 163.367
R593 B.n360 B.n195 163.367
R594 B.n361 B.n360 163.367
R595 B.n362 B.n361 163.367
R596 B.n362 B.n193 163.367
R597 B.n366 B.n193 163.367
R598 B.n367 B.n366 163.367
R599 B.n368 B.n367 163.367
R600 B.n368 B.n191 163.367
R601 B.n372 B.n191 163.367
R602 B.n373 B.n372 163.367
R603 B.n374 B.n373 163.367
R604 B.n374 B.n189 163.367
R605 B.n378 B.n189 163.367
R606 B.n379 B.n378 163.367
R607 B.n380 B.n379 163.367
R608 B.n380 B.n187 163.367
R609 B.n384 B.n187 163.367
R610 B.n385 B.n384 163.367
R611 B.n386 B.n385 163.367
R612 B.n386 B.n185 163.367
R613 B.n390 B.n185 163.367
R614 B.n391 B.n390 163.367
R615 B.n392 B.n391 163.367
R616 B.n392 B.n183 163.367
R617 B.n396 B.n183 163.367
R618 B.n397 B.n396 163.367
R619 B.n397 B.n179 163.367
R620 B.n401 B.n179 163.367
R621 B.n402 B.n401 163.367
R622 B.n403 B.n402 163.367
R623 B.n403 B.n177 163.367
R624 B.n407 B.n177 163.367
R625 B.n408 B.n407 163.367
R626 B.n409 B.n408 163.367
R627 B.n409 B.n173 163.367
R628 B.n414 B.n173 163.367
R629 B.n415 B.n414 163.367
R630 B.n416 B.n415 163.367
R631 B.n416 B.n171 163.367
R632 B.n420 B.n171 163.367
R633 B.n421 B.n420 163.367
R634 B.n422 B.n421 163.367
R635 B.n422 B.n169 163.367
R636 B.n426 B.n169 163.367
R637 B.n427 B.n426 163.367
R638 B.n428 B.n427 163.367
R639 B.n428 B.n167 163.367
R640 B.n432 B.n167 163.367
R641 B.n433 B.n432 163.367
R642 B.n434 B.n433 163.367
R643 B.n434 B.n165 163.367
R644 B.n438 B.n165 163.367
R645 B.n439 B.n438 163.367
R646 B.n440 B.n439 163.367
R647 B.n440 B.n163 163.367
R648 B.n444 B.n163 163.367
R649 B.n445 B.n444 163.367
R650 B.n446 B.n445 163.367
R651 B.n446 B.n161 163.367
R652 B.n450 B.n161 163.367
R653 B.n451 B.n450 163.367
R654 B.n452 B.n451 163.367
R655 B.n452 B.n159 163.367
R656 B.n456 B.n159 163.367
R657 B.n457 B.n456 163.367
R658 B.n458 B.n457 163.367
R659 B.n458 B.n157 163.367
R660 B.n462 B.n157 163.367
R661 B.n463 B.n462 163.367
R662 B.n464 B.n463 163.367
R663 B.n464 B.n155 163.367
R664 B.n468 B.n155 163.367
R665 B.n469 B.n468 163.367
R666 B.n470 B.n469 163.367
R667 B.n470 B.n153 163.367
R668 B.n474 B.n153 163.367
R669 B.n475 B.n474 163.367
R670 B.n476 B.n475 163.367
R671 B.n476 B.n151 163.367
R672 B.n480 B.n151 163.367
R673 B.n481 B.n480 163.367
R674 B.n482 B.n481 163.367
R675 B.n482 B.n149 163.367
R676 B.n486 B.n149 163.367
R677 B.n487 B.n486 163.367
R678 B.n488 B.n487 163.367
R679 B.n488 B.n147 163.367
R680 B.n492 B.n147 163.367
R681 B.n493 B.n492 163.367
R682 B.n494 B.n493 163.367
R683 B.n494 B.n145 163.367
R684 B.n498 B.n145 163.367
R685 B.n499 B.n498 163.367
R686 B.n500 B.n499 163.367
R687 B.n500 B.n143 163.367
R688 B.n505 B.n504 163.367
R689 B.n506 B.n505 163.367
R690 B.n506 B.n141 163.367
R691 B.n510 B.n141 163.367
R692 B.n511 B.n510 163.367
R693 B.n512 B.n511 163.367
R694 B.n512 B.n139 163.367
R695 B.n516 B.n139 163.367
R696 B.n517 B.n516 163.367
R697 B.n518 B.n517 163.367
R698 B.n518 B.n137 163.367
R699 B.n522 B.n137 163.367
R700 B.n523 B.n522 163.367
R701 B.n524 B.n523 163.367
R702 B.n524 B.n135 163.367
R703 B.n528 B.n135 163.367
R704 B.n529 B.n528 163.367
R705 B.n530 B.n529 163.367
R706 B.n530 B.n133 163.367
R707 B.n534 B.n133 163.367
R708 B.n535 B.n534 163.367
R709 B.n536 B.n535 163.367
R710 B.n536 B.n131 163.367
R711 B.n540 B.n131 163.367
R712 B.n541 B.n540 163.367
R713 B.n542 B.n541 163.367
R714 B.n542 B.n129 163.367
R715 B.n546 B.n129 163.367
R716 B.n547 B.n546 163.367
R717 B.n548 B.n547 163.367
R718 B.n548 B.n127 163.367
R719 B.n552 B.n127 163.367
R720 B.n553 B.n552 163.367
R721 B.n554 B.n553 163.367
R722 B.n554 B.n125 163.367
R723 B.n558 B.n125 163.367
R724 B.n559 B.n558 163.367
R725 B.n560 B.n559 163.367
R726 B.n560 B.n123 163.367
R727 B.n564 B.n123 163.367
R728 B.n565 B.n564 163.367
R729 B.n566 B.n565 163.367
R730 B.n566 B.n121 163.367
R731 B.n570 B.n121 163.367
R732 B.n571 B.n570 163.367
R733 B.n572 B.n571 163.367
R734 B.n572 B.n119 163.367
R735 B.n576 B.n119 163.367
R736 B.n577 B.n576 163.367
R737 B.n578 B.n577 163.367
R738 B.n578 B.n117 163.367
R739 B.n582 B.n117 163.367
R740 B.n583 B.n582 163.367
R741 B.n584 B.n583 163.367
R742 B.n584 B.n115 163.367
R743 B.n588 B.n115 163.367
R744 B.n589 B.n588 163.367
R745 B.n590 B.n589 163.367
R746 B.n590 B.n113 163.367
R747 B.n594 B.n113 163.367
R748 B.n595 B.n594 163.367
R749 B.n596 B.n595 163.367
R750 B.n596 B.n111 163.367
R751 B.n600 B.n111 163.367
R752 B.n601 B.n600 163.367
R753 B.n602 B.n601 163.367
R754 B.n602 B.n109 163.367
R755 B.n606 B.n109 163.367
R756 B.n607 B.n606 163.367
R757 B.n608 B.n607 163.367
R758 B.n608 B.n107 163.367
R759 B.n612 B.n107 163.367
R760 B.n613 B.n612 163.367
R761 B.n614 B.n613 163.367
R762 B.n614 B.n105 163.367
R763 B.n618 B.n105 163.367
R764 B.n619 B.n618 163.367
R765 B.n620 B.n619 163.367
R766 B.n620 B.n103 163.367
R767 B.n624 B.n103 163.367
R768 B.n625 B.n624 163.367
R769 B.n626 B.n625 163.367
R770 B.n626 B.n101 163.367
R771 B.n630 B.n101 163.367
R772 B.n631 B.n630 163.367
R773 B.n632 B.n631 163.367
R774 B.n632 B.n99 163.367
R775 B.n636 B.n99 163.367
R776 B.n637 B.n636 163.367
R777 B.n638 B.n637 163.367
R778 B.n638 B.n97 163.367
R779 B.n642 B.n97 163.367
R780 B.n643 B.n642 163.367
R781 B.n644 B.n643 163.367
R782 B.n842 B.n841 163.367
R783 B.n841 B.n840 163.367
R784 B.n840 B.n27 163.367
R785 B.n836 B.n27 163.367
R786 B.n836 B.n835 163.367
R787 B.n835 B.n834 163.367
R788 B.n834 B.n29 163.367
R789 B.n830 B.n29 163.367
R790 B.n830 B.n829 163.367
R791 B.n829 B.n828 163.367
R792 B.n828 B.n31 163.367
R793 B.n824 B.n31 163.367
R794 B.n824 B.n823 163.367
R795 B.n823 B.n822 163.367
R796 B.n822 B.n33 163.367
R797 B.n818 B.n33 163.367
R798 B.n818 B.n817 163.367
R799 B.n817 B.n816 163.367
R800 B.n816 B.n35 163.367
R801 B.n812 B.n35 163.367
R802 B.n812 B.n811 163.367
R803 B.n811 B.n810 163.367
R804 B.n810 B.n37 163.367
R805 B.n806 B.n37 163.367
R806 B.n806 B.n805 163.367
R807 B.n805 B.n804 163.367
R808 B.n804 B.n39 163.367
R809 B.n800 B.n39 163.367
R810 B.n800 B.n799 163.367
R811 B.n799 B.n798 163.367
R812 B.n798 B.n41 163.367
R813 B.n794 B.n41 163.367
R814 B.n794 B.n793 163.367
R815 B.n793 B.n792 163.367
R816 B.n792 B.n43 163.367
R817 B.n788 B.n43 163.367
R818 B.n788 B.n787 163.367
R819 B.n787 B.n786 163.367
R820 B.n786 B.n45 163.367
R821 B.n782 B.n45 163.367
R822 B.n782 B.n781 163.367
R823 B.n781 B.n780 163.367
R824 B.n780 B.n47 163.367
R825 B.n776 B.n47 163.367
R826 B.n776 B.n775 163.367
R827 B.n775 B.n774 163.367
R828 B.n774 B.n49 163.367
R829 B.n770 B.n49 163.367
R830 B.n770 B.n769 163.367
R831 B.n769 B.n768 163.367
R832 B.n768 B.n51 163.367
R833 B.n764 B.n51 163.367
R834 B.n764 B.n763 163.367
R835 B.n763 B.n762 163.367
R836 B.n762 B.n53 163.367
R837 B.n758 B.n53 163.367
R838 B.n758 B.n757 163.367
R839 B.n757 B.n756 163.367
R840 B.n756 B.n55 163.367
R841 B.n752 B.n55 163.367
R842 B.n752 B.n751 163.367
R843 B.n751 B.n59 163.367
R844 B.n747 B.n59 163.367
R845 B.n747 B.n746 163.367
R846 B.n746 B.n745 163.367
R847 B.n745 B.n61 163.367
R848 B.n741 B.n61 163.367
R849 B.n741 B.n740 163.367
R850 B.n740 B.n739 163.367
R851 B.n739 B.n63 163.367
R852 B.n734 B.n63 163.367
R853 B.n734 B.n733 163.367
R854 B.n733 B.n732 163.367
R855 B.n732 B.n67 163.367
R856 B.n728 B.n67 163.367
R857 B.n728 B.n727 163.367
R858 B.n727 B.n726 163.367
R859 B.n726 B.n69 163.367
R860 B.n722 B.n69 163.367
R861 B.n722 B.n721 163.367
R862 B.n721 B.n720 163.367
R863 B.n720 B.n71 163.367
R864 B.n716 B.n71 163.367
R865 B.n716 B.n715 163.367
R866 B.n715 B.n714 163.367
R867 B.n714 B.n73 163.367
R868 B.n710 B.n73 163.367
R869 B.n710 B.n709 163.367
R870 B.n709 B.n708 163.367
R871 B.n708 B.n75 163.367
R872 B.n704 B.n75 163.367
R873 B.n704 B.n703 163.367
R874 B.n703 B.n702 163.367
R875 B.n702 B.n77 163.367
R876 B.n698 B.n77 163.367
R877 B.n698 B.n697 163.367
R878 B.n697 B.n696 163.367
R879 B.n696 B.n79 163.367
R880 B.n692 B.n79 163.367
R881 B.n692 B.n691 163.367
R882 B.n691 B.n690 163.367
R883 B.n690 B.n81 163.367
R884 B.n686 B.n81 163.367
R885 B.n686 B.n685 163.367
R886 B.n685 B.n684 163.367
R887 B.n684 B.n83 163.367
R888 B.n680 B.n83 163.367
R889 B.n680 B.n679 163.367
R890 B.n679 B.n678 163.367
R891 B.n678 B.n85 163.367
R892 B.n674 B.n85 163.367
R893 B.n674 B.n673 163.367
R894 B.n673 B.n672 163.367
R895 B.n672 B.n87 163.367
R896 B.n668 B.n87 163.367
R897 B.n668 B.n667 163.367
R898 B.n667 B.n666 163.367
R899 B.n666 B.n89 163.367
R900 B.n662 B.n89 163.367
R901 B.n662 B.n661 163.367
R902 B.n661 B.n660 163.367
R903 B.n660 B.n91 163.367
R904 B.n656 B.n91 163.367
R905 B.n656 B.n655 163.367
R906 B.n655 B.n654 163.367
R907 B.n654 B.n93 163.367
R908 B.n650 B.n93 163.367
R909 B.n650 B.n649 163.367
R910 B.n649 B.n648 163.367
R911 B.n648 B.n95 163.367
R912 B.n175 B.t1 109.644
R913 B.n65 B.t5 109.644
R914 B.n181 B.t7 109.62
R915 B.n57 B.t11 109.62
R916 B.n175 B.n174 64.3884
R917 B.n181 B.n180 64.3884
R918 B.n57 B.n56 64.3884
R919 B.n65 B.n64 64.3884
R920 B.n411 B.n175 59.5399
R921 B.n182 B.n181 59.5399
R922 B.n58 B.n57 59.5399
R923 B.n737 B.n65 59.5399
R924 B.n844 B.n843 35.7468
R925 B.n646 B.n645 35.7468
R926 B.n503 B.n502 35.7468
R927 B.n305 B.n304 35.7468
R928 B B.n915 18.0485
R929 B.n843 B.n26 10.6151
R930 B.n839 B.n26 10.6151
R931 B.n839 B.n838 10.6151
R932 B.n838 B.n837 10.6151
R933 B.n837 B.n28 10.6151
R934 B.n833 B.n28 10.6151
R935 B.n833 B.n832 10.6151
R936 B.n832 B.n831 10.6151
R937 B.n831 B.n30 10.6151
R938 B.n827 B.n30 10.6151
R939 B.n827 B.n826 10.6151
R940 B.n826 B.n825 10.6151
R941 B.n825 B.n32 10.6151
R942 B.n821 B.n32 10.6151
R943 B.n821 B.n820 10.6151
R944 B.n820 B.n819 10.6151
R945 B.n819 B.n34 10.6151
R946 B.n815 B.n34 10.6151
R947 B.n815 B.n814 10.6151
R948 B.n814 B.n813 10.6151
R949 B.n813 B.n36 10.6151
R950 B.n809 B.n36 10.6151
R951 B.n809 B.n808 10.6151
R952 B.n808 B.n807 10.6151
R953 B.n807 B.n38 10.6151
R954 B.n803 B.n38 10.6151
R955 B.n803 B.n802 10.6151
R956 B.n802 B.n801 10.6151
R957 B.n801 B.n40 10.6151
R958 B.n797 B.n40 10.6151
R959 B.n797 B.n796 10.6151
R960 B.n796 B.n795 10.6151
R961 B.n795 B.n42 10.6151
R962 B.n791 B.n42 10.6151
R963 B.n791 B.n790 10.6151
R964 B.n790 B.n789 10.6151
R965 B.n789 B.n44 10.6151
R966 B.n785 B.n44 10.6151
R967 B.n785 B.n784 10.6151
R968 B.n784 B.n783 10.6151
R969 B.n783 B.n46 10.6151
R970 B.n779 B.n46 10.6151
R971 B.n779 B.n778 10.6151
R972 B.n778 B.n777 10.6151
R973 B.n777 B.n48 10.6151
R974 B.n773 B.n48 10.6151
R975 B.n773 B.n772 10.6151
R976 B.n772 B.n771 10.6151
R977 B.n771 B.n50 10.6151
R978 B.n767 B.n50 10.6151
R979 B.n767 B.n766 10.6151
R980 B.n766 B.n765 10.6151
R981 B.n765 B.n52 10.6151
R982 B.n761 B.n52 10.6151
R983 B.n761 B.n760 10.6151
R984 B.n760 B.n759 10.6151
R985 B.n759 B.n54 10.6151
R986 B.n755 B.n54 10.6151
R987 B.n755 B.n754 10.6151
R988 B.n754 B.n753 10.6151
R989 B.n750 B.n749 10.6151
R990 B.n749 B.n748 10.6151
R991 B.n748 B.n60 10.6151
R992 B.n744 B.n60 10.6151
R993 B.n744 B.n743 10.6151
R994 B.n743 B.n742 10.6151
R995 B.n742 B.n62 10.6151
R996 B.n738 B.n62 10.6151
R997 B.n736 B.n735 10.6151
R998 B.n735 B.n66 10.6151
R999 B.n731 B.n66 10.6151
R1000 B.n731 B.n730 10.6151
R1001 B.n730 B.n729 10.6151
R1002 B.n729 B.n68 10.6151
R1003 B.n725 B.n68 10.6151
R1004 B.n725 B.n724 10.6151
R1005 B.n724 B.n723 10.6151
R1006 B.n723 B.n70 10.6151
R1007 B.n719 B.n70 10.6151
R1008 B.n719 B.n718 10.6151
R1009 B.n718 B.n717 10.6151
R1010 B.n717 B.n72 10.6151
R1011 B.n713 B.n72 10.6151
R1012 B.n713 B.n712 10.6151
R1013 B.n712 B.n711 10.6151
R1014 B.n711 B.n74 10.6151
R1015 B.n707 B.n74 10.6151
R1016 B.n707 B.n706 10.6151
R1017 B.n706 B.n705 10.6151
R1018 B.n705 B.n76 10.6151
R1019 B.n701 B.n76 10.6151
R1020 B.n701 B.n700 10.6151
R1021 B.n700 B.n699 10.6151
R1022 B.n699 B.n78 10.6151
R1023 B.n695 B.n78 10.6151
R1024 B.n695 B.n694 10.6151
R1025 B.n694 B.n693 10.6151
R1026 B.n693 B.n80 10.6151
R1027 B.n689 B.n80 10.6151
R1028 B.n689 B.n688 10.6151
R1029 B.n688 B.n687 10.6151
R1030 B.n687 B.n82 10.6151
R1031 B.n683 B.n82 10.6151
R1032 B.n683 B.n682 10.6151
R1033 B.n682 B.n681 10.6151
R1034 B.n681 B.n84 10.6151
R1035 B.n677 B.n84 10.6151
R1036 B.n677 B.n676 10.6151
R1037 B.n676 B.n675 10.6151
R1038 B.n675 B.n86 10.6151
R1039 B.n671 B.n86 10.6151
R1040 B.n671 B.n670 10.6151
R1041 B.n670 B.n669 10.6151
R1042 B.n669 B.n88 10.6151
R1043 B.n665 B.n88 10.6151
R1044 B.n665 B.n664 10.6151
R1045 B.n664 B.n663 10.6151
R1046 B.n663 B.n90 10.6151
R1047 B.n659 B.n90 10.6151
R1048 B.n659 B.n658 10.6151
R1049 B.n658 B.n657 10.6151
R1050 B.n657 B.n92 10.6151
R1051 B.n653 B.n92 10.6151
R1052 B.n653 B.n652 10.6151
R1053 B.n652 B.n651 10.6151
R1054 B.n651 B.n94 10.6151
R1055 B.n647 B.n94 10.6151
R1056 B.n647 B.n646 10.6151
R1057 B.n503 B.n142 10.6151
R1058 B.n507 B.n142 10.6151
R1059 B.n508 B.n507 10.6151
R1060 B.n509 B.n508 10.6151
R1061 B.n509 B.n140 10.6151
R1062 B.n513 B.n140 10.6151
R1063 B.n514 B.n513 10.6151
R1064 B.n515 B.n514 10.6151
R1065 B.n515 B.n138 10.6151
R1066 B.n519 B.n138 10.6151
R1067 B.n520 B.n519 10.6151
R1068 B.n521 B.n520 10.6151
R1069 B.n521 B.n136 10.6151
R1070 B.n525 B.n136 10.6151
R1071 B.n526 B.n525 10.6151
R1072 B.n527 B.n526 10.6151
R1073 B.n527 B.n134 10.6151
R1074 B.n531 B.n134 10.6151
R1075 B.n532 B.n531 10.6151
R1076 B.n533 B.n532 10.6151
R1077 B.n533 B.n132 10.6151
R1078 B.n537 B.n132 10.6151
R1079 B.n538 B.n537 10.6151
R1080 B.n539 B.n538 10.6151
R1081 B.n539 B.n130 10.6151
R1082 B.n543 B.n130 10.6151
R1083 B.n544 B.n543 10.6151
R1084 B.n545 B.n544 10.6151
R1085 B.n545 B.n128 10.6151
R1086 B.n549 B.n128 10.6151
R1087 B.n550 B.n549 10.6151
R1088 B.n551 B.n550 10.6151
R1089 B.n551 B.n126 10.6151
R1090 B.n555 B.n126 10.6151
R1091 B.n556 B.n555 10.6151
R1092 B.n557 B.n556 10.6151
R1093 B.n557 B.n124 10.6151
R1094 B.n561 B.n124 10.6151
R1095 B.n562 B.n561 10.6151
R1096 B.n563 B.n562 10.6151
R1097 B.n563 B.n122 10.6151
R1098 B.n567 B.n122 10.6151
R1099 B.n568 B.n567 10.6151
R1100 B.n569 B.n568 10.6151
R1101 B.n569 B.n120 10.6151
R1102 B.n573 B.n120 10.6151
R1103 B.n574 B.n573 10.6151
R1104 B.n575 B.n574 10.6151
R1105 B.n575 B.n118 10.6151
R1106 B.n579 B.n118 10.6151
R1107 B.n580 B.n579 10.6151
R1108 B.n581 B.n580 10.6151
R1109 B.n581 B.n116 10.6151
R1110 B.n585 B.n116 10.6151
R1111 B.n586 B.n585 10.6151
R1112 B.n587 B.n586 10.6151
R1113 B.n587 B.n114 10.6151
R1114 B.n591 B.n114 10.6151
R1115 B.n592 B.n591 10.6151
R1116 B.n593 B.n592 10.6151
R1117 B.n593 B.n112 10.6151
R1118 B.n597 B.n112 10.6151
R1119 B.n598 B.n597 10.6151
R1120 B.n599 B.n598 10.6151
R1121 B.n599 B.n110 10.6151
R1122 B.n603 B.n110 10.6151
R1123 B.n604 B.n603 10.6151
R1124 B.n605 B.n604 10.6151
R1125 B.n605 B.n108 10.6151
R1126 B.n609 B.n108 10.6151
R1127 B.n610 B.n609 10.6151
R1128 B.n611 B.n610 10.6151
R1129 B.n611 B.n106 10.6151
R1130 B.n615 B.n106 10.6151
R1131 B.n616 B.n615 10.6151
R1132 B.n617 B.n616 10.6151
R1133 B.n617 B.n104 10.6151
R1134 B.n621 B.n104 10.6151
R1135 B.n622 B.n621 10.6151
R1136 B.n623 B.n622 10.6151
R1137 B.n623 B.n102 10.6151
R1138 B.n627 B.n102 10.6151
R1139 B.n628 B.n627 10.6151
R1140 B.n629 B.n628 10.6151
R1141 B.n629 B.n100 10.6151
R1142 B.n633 B.n100 10.6151
R1143 B.n634 B.n633 10.6151
R1144 B.n635 B.n634 10.6151
R1145 B.n635 B.n98 10.6151
R1146 B.n639 B.n98 10.6151
R1147 B.n640 B.n639 10.6151
R1148 B.n641 B.n640 10.6151
R1149 B.n641 B.n96 10.6151
R1150 B.n645 B.n96 10.6151
R1151 B.n305 B.n212 10.6151
R1152 B.n309 B.n212 10.6151
R1153 B.n310 B.n309 10.6151
R1154 B.n311 B.n310 10.6151
R1155 B.n311 B.n210 10.6151
R1156 B.n315 B.n210 10.6151
R1157 B.n316 B.n315 10.6151
R1158 B.n317 B.n316 10.6151
R1159 B.n317 B.n208 10.6151
R1160 B.n321 B.n208 10.6151
R1161 B.n322 B.n321 10.6151
R1162 B.n323 B.n322 10.6151
R1163 B.n323 B.n206 10.6151
R1164 B.n327 B.n206 10.6151
R1165 B.n328 B.n327 10.6151
R1166 B.n329 B.n328 10.6151
R1167 B.n329 B.n204 10.6151
R1168 B.n333 B.n204 10.6151
R1169 B.n334 B.n333 10.6151
R1170 B.n335 B.n334 10.6151
R1171 B.n335 B.n202 10.6151
R1172 B.n339 B.n202 10.6151
R1173 B.n340 B.n339 10.6151
R1174 B.n341 B.n340 10.6151
R1175 B.n341 B.n200 10.6151
R1176 B.n345 B.n200 10.6151
R1177 B.n346 B.n345 10.6151
R1178 B.n347 B.n346 10.6151
R1179 B.n347 B.n198 10.6151
R1180 B.n351 B.n198 10.6151
R1181 B.n352 B.n351 10.6151
R1182 B.n353 B.n352 10.6151
R1183 B.n353 B.n196 10.6151
R1184 B.n357 B.n196 10.6151
R1185 B.n358 B.n357 10.6151
R1186 B.n359 B.n358 10.6151
R1187 B.n359 B.n194 10.6151
R1188 B.n363 B.n194 10.6151
R1189 B.n364 B.n363 10.6151
R1190 B.n365 B.n364 10.6151
R1191 B.n365 B.n192 10.6151
R1192 B.n369 B.n192 10.6151
R1193 B.n370 B.n369 10.6151
R1194 B.n371 B.n370 10.6151
R1195 B.n371 B.n190 10.6151
R1196 B.n375 B.n190 10.6151
R1197 B.n376 B.n375 10.6151
R1198 B.n377 B.n376 10.6151
R1199 B.n377 B.n188 10.6151
R1200 B.n381 B.n188 10.6151
R1201 B.n382 B.n381 10.6151
R1202 B.n383 B.n382 10.6151
R1203 B.n383 B.n186 10.6151
R1204 B.n387 B.n186 10.6151
R1205 B.n388 B.n387 10.6151
R1206 B.n389 B.n388 10.6151
R1207 B.n389 B.n184 10.6151
R1208 B.n393 B.n184 10.6151
R1209 B.n394 B.n393 10.6151
R1210 B.n395 B.n394 10.6151
R1211 B.n399 B.n398 10.6151
R1212 B.n400 B.n399 10.6151
R1213 B.n400 B.n178 10.6151
R1214 B.n404 B.n178 10.6151
R1215 B.n405 B.n404 10.6151
R1216 B.n406 B.n405 10.6151
R1217 B.n406 B.n176 10.6151
R1218 B.n410 B.n176 10.6151
R1219 B.n413 B.n412 10.6151
R1220 B.n413 B.n172 10.6151
R1221 B.n417 B.n172 10.6151
R1222 B.n418 B.n417 10.6151
R1223 B.n419 B.n418 10.6151
R1224 B.n419 B.n170 10.6151
R1225 B.n423 B.n170 10.6151
R1226 B.n424 B.n423 10.6151
R1227 B.n425 B.n424 10.6151
R1228 B.n425 B.n168 10.6151
R1229 B.n429 B.n168 10.6151
R1230 B.n430 B.n429 10.6151
R1231 B.n431 B.n430 10.6151
R1232 B.n431 B.n166 10.6151
R1233 B.n435 B.n166 10.6151
R1234 B.n436 B.n435 10.6151
R1235 B.n437 B.n436 10.6151
R1236 B.n437 B.n164 10.6151
R1237 B.n441 B.n164 10.6151
R1238 B.n442 B.n441 10.6151
R1239 B.n443 B.n442 10.6151
R1240 B.n443 B.n162 10.6151
R1241 B.n447 B.n162 10.6151
R1242 B.n448 B.n447 10.6151
R1243 B.n449 B.n448 10.6151
R1244 B.n449 B.n160 10.6151
R1245 B.n453 B.n160 10.6151
R1246 B.n454 B.n453 10.6151
R1247 B.n455 B.n454 10.6151
R1248 B.n455 B.n158 10.6151
R1249 B.n459 B.n158 10.6151
R1250 B.n460 B.n459 10.6151
R1251 B.n461 B.n460 10.6151
R1252 B.n461 B.n156 10.6151
R1253 B.n465 B.n156 10.6151
R1254 B.n466 B.n465 10.6151
R1255 B.n467 B.n466 10.6151
R1256 B.n467 B.n154 10.6151
R1257 B.n471 B.n154 10.6151
R1258 B.n472 B.n471 10.6151
R1259 B.n473 B.n472 10.6151
R1260 B.n473 B.n152 10.6151
R1261 B.n477 B.n152 10.6151
R1262 B.n478 B.n477 10.6151
R1263 B.n479 B.n478 10.6151
R1264 B.n479 B.n150 10.6151
R1265 B.n483 B.n150 10.6151
R1266 B.n484 B.n483 10.6151
R1267 B.n485 B.n484 10.6151
R1268 B.n485 B.n148 10.6151
R1269 B.n489 B.n148 10.6151
R1270 B.n490 B.n489 10.6151
R1271 B.n491 B.n490 10.6151
R1272 B.n491 B.n146 10.6151
R1273 B.n495 B.n146 10.6151
R1274 B.n496 B.n495 10.6151
R1275 B.n497 B.n496 10.6151
R1276 B.n497 B.n144 10.6151
R1277 B.n501 B.n144 10.6151
R1278 B.n502 B.n501 10.6151
R1279 B.n304 B.n303 10.6151
R1280 B.n303 B.n214 10.6151
R1281 B.n299 B.n214 10.6151
R1282 B.n299 B.n298 10.6151
R1283 B.n298 B.n297 10.6151
R1284 B.n297 B.n216 10.6151
R1285 B.n293 B.n216 10.6151
R1286 B.n293 B.n292 10.6151
R1287 B.n292 B.n291 10.6151
R1288 B.n291 B.n218 10.6151
R1289 B.n287 B.n218 10.6151
R1290 B.n287 B.n286 10.6151
R1291 B.n286 B.n285 10.6151
R1292 B.n285 B.n220 10.6151
R1293 B.n281 B.n220 10.6151
R1294 B.n281 B.n280 10.6151
R1295 B.n280 B.n279 10.6151
R1296 B.n279 B.n222 10.6151
R1297 B.n275 B.n222 10.6151
R1298 B.n275 B.n274 10.6151
R1299 B.n274 B.n273 10.6151
R1300 B.n273 B.n224 10.6151
R1301 B.n269 B.n224 10.6151
R1302 B.n269 B.n268 10.6151
R1303 B.n268 B.n267 10.6151
R1304 B.n267 B.n226 10.6151
R1305 B.n263 B.n226 10.6151
R1306 B.n263 B.n262 10.6151
R1307 B.n262 B.n261 10.6151
R1308 B.n261 B.n228 10.6151
R1309 B.n257 B.n228 10.6151
R1310 B.n257 B.n256 10.6151
R1311 B.n256 B.n255 10.6151
R1312 B.n255 B.n230 10.6151
R1313 B.n251 B.n230 10.6151
R1314 B.n251 B.n250 10.6151
R1315 B.n250 B.n249 10.6151
R1316 B.n249 B.n232 10.6151
R1317 B.n245 B.n232 10.6151
R1318 B.n245 B.n244 10.6151
R1319 B.n244 B.n243 10.6151
R1320 B.n243 B.n234 10.6151
R1321 B.n239 B.n234 10.6151
R1322 B.n239 B.n238 10.6151
R1323 B.n238 B.n237 10.6151
R1324 B.n237 B.n0 10.6151
R1325 B.n911 B.n1 10.6151
R1326 B.n911 B.n910 10.6151
R1327 B.n910 B.n909 10.6151
R1328 B.n909 B.n4 10.6151
R1329 B.n905 B.n4 10.6151
R1330 B.n905 B.n904 10.6151
R1331 B.n904 B.n903 10.6151
R1332 B.n903 B.n6 10.6151
R1333 B.n899 B.n6 10.6151
R1334 B.n899 B.n898 10.6151
R1335 B.n898 B.n897 10.6151
R1336 B.n897 B.n8 10.6151
R1337 B.n893 B.n8 10.6151
R1338 B.n893 B.n892 10.6151
R1339 B.n892 B.n891 10.6151
R1340 B.n891 B.n10 10.6151
R1341 B.n887 B.n10 10.6151
R1342 B.n887 B.n886 10.6151
R1343 B.n886 B.n885 10.6151
R1344 B.n885 B.n12 10.6151
R1345 B.n881 B.n12 10.6151
R1346 B.n881 B.n880 10.6151
R1347 B.n880 B.n879 10.6151
R1348 B.n879 B.n14 10.6151
R1349 B.n875 B.n14 10.6151
R1350 B.n875 B.n874 10.6151
R1351 B.n874 B.n873 10.6151
R1352 B.n873 B.n16 10.6151
R1353 B.n869 B.n16 10.6151
R1354 B.n869 B.n868 10.6151
R1355 B.n868 B.n867 10.6151
R1356 B.n867 B.n18 10.6151
R1357 B.n863 B.n18 10.6151
R1358 B.n863 B.n862 10.6151
R1359 B.n862 B.n861 10.6151
R1360 B.n861 B.n20 10.6151
R1361 B.n857 B.n20 10.6151
R1362 B.n857 B.n856 10.6151
R1363 B.n856 B.n855 10.6151
R1364 B.n855 B.n22 10.6151
R1365 B.n851 B.n22 10.6151
R1366 B.n851 B.n850 10.6151
R1367 B.n850 B.n849 10.6151
R1368 B.n849 B.n24 10.6151
R1369 B.n845 B.n24 10.6151
R1370 B.n845 B.n844 10.6151
R1371 B.n750 B.n58 6.5566
R1372 B.n738 B.n737 6.5566
R1373 B.n398 B.n182 6.5566
R1374 B.n411 B.n410 6.5566
R1375 B.n753 B.n58 4.05904
R1376 B.n737 B.n736 4.05904
R1377 B.n395 B.n182 4.05904
R1378 B.n412 B.n411 4.05904
R1379 B.n915 B.n0 2.81026
R1380 B.n915 B.n1 2.81026
R1381 VP.n11 VP.t1 182.69
R1382 VP.n13 VP.n10 161.3
R1383 VP.n15 VP.n14 161.3
R1384 VP.n16 VP.n9 161.3
R1385 VP.n18 VP.n17 161.3
R1386 VP.n19 VP.n8 161.3
R1387 VP.n21 VP.n20 161.3
R1388 VP.n44 VP.n43 161.3
R1389 VP.n42 VP.n1 161.3
R1390 VP.n41 VP.n40 161.3
R1391 VP.n39 VP.n2 161.3
R1392 VP.n38 VP.n37 161.3
R1393 VP.n36 VP.n3 161.3
R1394 VP.n35 VP.n34 161.3
R1395 VP.n33 VP.n4 161.3
R1396 VP.n32 VP.n31 161.3
R1397 VP.n30 VP.n5 161.3
R1398 VP.n29 VP.n28 161.3
R1399 VP.n27 VP.n6 161.3
R1400 VP.n26 VP.n25 161.3
R1401 VP.n35 VP.t3 149.436
R1402 VP.n24 VP.t0 149.436
R1403 VP.n0 VP.t2 149.436
R1404 VP.n12 VP.t4 149.436
R1405 VP.n7 VP.t5 149.436
R1406 VP.n24 VP.n23 74.5068
R1407 VP.n45 VP.n0 74.5068
R1408 VP.n22 VP.n7 74.5068
R1409 VP.n30 VP.n29 56.0773
R1410 VP.n41 VP.n2 56.0773
R1411 VP.n18 VP.n9 56.0773
R1412 VP.n23 VP.n22 55.2117
R1413 VP.n12 VP.n11 49.3258
R1414 VP.n31 VP.n30 25.0767
R1415 VP.n37 VP.n2 25.0767
R1416 VP.n14 VP.n9 25.0767
R1417 VP.n25 VP.n6 24.5923
R1418 VP.n29 VP.n6 24.5923
R1419 VP.n31 VP.n4 24.5923
R1420 VP.n35 VP.n4 24.5923
R1421 VP.n36 VP.n35 24.5923
R1422 VP.n37 VP.n36 24.5923
R1423 VP.n42 VP.n41 24.5923
R1424 VP.n43 VP.n42 24.5923
R1425 VP.n19 VP.n18 24.5923
R1426 VP.n20 VP.n19 24.5923
R1427 VP.n13 VP.n12 24.5923
R1428 VP.n14 VP.n13 24.5923
R1429 VP.n25 VP.n24 15.7393
R1430 VP.n43 VP.n0 15.7393
R1431 VP.n20 VP.n7 15.7393
R1432 VP.n11 VP.n10 4.10785
R1433 VP.n22 VP.n21 0.354861
R1434 VP.n26 VP.n23 0.354861
R1435 VP.n45 VP.n44 0.354861
R1436 VP VP.n45 0.267071
R1437 VP.n15 VP.n10 0.189894
R1438 VP.n16 VP.n15 0.189894
R1439 VP.n17 VP.n16 0.189894
R1440 VP.n17 VP.n8 0.189894
R1441 VP.n21 VP.n8 0.189894
R1442 VP.n27 VP.n26 0.189894
R1443 VP.n28 VP.n27 0.189894
R1444 VP.n28 VP.n5 0.189894
R1445 VP.n32 VP.n5 0.189894
R1446 VP.n33 VP.n32 0.189894
R1447 VP.n34 VP.n33 0.189894
R1448 VP.n34 VP.n3 0.189894
R1449 VP.n38 VP.n3 0.189894
R1450 VP.n39 VP.n38 0.189894
R1451 VP.n40 VP.n39 0.189894
R1452 VP.n40 VP.n1 0.189894
R1453 VP.n44 VP.n1 0.189894
R1454 VTAIL.n7 VTAIL.t0 52.4433
R1455 VTAIL.n11 VTAIL.t11 52.4431
R1456 VTAIL.n2 VTAIL.t9 52.4431
R1457 VTAIL.n10 VTAIL.t10 52.4431
R1458 VTAIL.n9 VTAIL.n8 50.6901
R1459 VTAIL.n6 VTAIL.n5 50.6901
R1460 VTAIL.n1 VTAIL.n0 50.6899
R1461 VTAIL.n4 VTAIL.n3 50.6899
R1462 VTAIL.n6 VTAIL.n4 34.0738
R1463 VTAIL.n11 VTAIL.n10 31.2117
R1464 VTAIL.n7 VTAIL.n6 2.86257
R1465 VTAIL.n10 VTAIL.n9 2.86257
R1466 VTAIL.n4 VTAIL.n2 2.86257
R1467 VTAIL VTAIL.n11 2.08886
R1468 VTAIL.n9 VTAIL.n7 1.90136
R1469 VTAIL.n2 VTAIL.n1 1.90136
R1470 VTAIL.n0 VTAIL.t4 1.75374
R1471 VTAIL.n0 VTAIL.t2 1.75374
R1472 VTAIL.n3 VTAIL.t5 1.75374
R1473 VTAIL.n3 VTAIL.t6 1.75374
R1474 VTAIL.n8 VTAIL.t8 1.75374
R1475 VTAIL.n8 VTAIL.t7 1.75374
R1476 VTAIL.n5 VTAIL.t3 1.75374
R1477 VTAIL.n5 VTAIL.t1 1.75374
R1478 VTAIL VTAIL.n1 0.774207
R1479 VDD1 VDD1.t4 71.3268
R1480 VDD1.n1 VDD1.t5 71.2131
R1481 VDD1.n1 VDD1.n0 68.0288
R1482 VDD1.n3 VDD1.n2 67.3687
R1483 VDD1.n3 VDD1.n1 51.0138
R1484 VDD1.n2 VDD1.t1 1.75374
R1485 VDD1.n2 VDD1.t0 1.75374
R1486 VDD1.n0 VDD1.t2 1.75374
R1487 VDD1.n0 VDD1.t3 1.75374
R1488 VDD1 VDD1.n3 0.657828
R1489 VN.n20 VN.t2 182.69
R1490 VN.n4 VN.t1 182.69
R1491 VN.n30 VN.n29 161.3
R1492 VN.n28 VN.n17 161.3
R1493 VN.n27 VN.n26 161.3
R1494 VN.n25 VN.n18 161.3
R1495 VN.n24 VN.n23 161.3
R1496 VN.n22 VN.n19 161.3
R1497 VN.n14 VN.n13 161.3
R1498 VN.n12 VN.n1 161.3
R1499 VN.n11 VN.n10 161.3
R1500 VN.n9 VN.n2 161.3
R1501 VN.n8 VN.n7 161.3
R1502 VN.n6 VN.n3 161.3
R1503 VN.n5 VN.t5 149.436
R1504 VN.n0 VN.t4 149.436
R1505 VN.n21 VN.t0 149.436
R1506 VN.n16 VN.t3 149.436
R1507 VN.n15 VN.n0 74.5068
R1508 VN.n31 VN.n16 74.5068
R1509 VN.n11 VN.n2 56.0773
R1510 VN.n27 VN.n18 56.0773
R1511 VN VN.n31 55.3769
R1512 VN.n5 VN.n4 49.3258
R1513 VN.n21 VN.n20 49.3258
R1514 VN.n7 VN.n2 25.0767
R1515 VN.n23 VN.n18 25.0767
R1516 VN.n6 VN.n5 24.5923
R1517 VN.n7 VN.n6 24.5923
R1518 VN.n12 VN.n11 24.5923
R1519 VN.n13 VN.n12 24.5923
R1520 VN.n23 VN.n22 24.5923
R1521 VN.n22 VN.n21 24.5923
R1522 VN.n29 VN.n28 24.5923
R1523 VN.n28 VN.n27 24.5923
R1524 VN.n13 VN.n0 15.7393
R1525 VN.n29 VN.n16 15.7393
R1526 VN.n4 VN.n3 4.10787
R1527 VN.n20 VN.n19 4.10787
R1528 VN.n31 VN.n30 0.354861
R1529 VN.n15 VN.n14 0.354861
R1530 VN VN.n15 0.267071
R1531 VN.n30 VN.n17 0.189894
R1532 VN.n26 VN.n17 0.189894
R1533 VN.n26 VN.n25 0.189894
R1534 VN.n25 VN.n24 0.189894
R1535 VN.n24 VN.n19 0.189894
R1536 VN.n8 VN.n3 0.189894
R1537 VN.n9 VN.n8 0.189894
R1538 VN.n10 VN.n9 0.189894
R1539 VN.n10 VN.n1 0.189894
R1540 VN.n14 VN.n1 0.189894
R1541 VDD2.n1 VDD2.t4 71.2131
R1542 VDD2.n2 VDD2.t2 69.1221
R1543 VDD2.n1 VDD2.n0 68.0288
R1544 VDD2 VDD2.n3 68.026
R1545 VDD2.n2 VDD2.n1 48.9998
R1546 VDD2 VDD2.n2 2.20524
R1547 VDD2.n3 VDD2.t5 1.75374
R1548 VDD2.n3 VDD2.t3 1.75374
R1549 VDD2.n0 VDD2.t0 1.75374
R1550 VDD2.n0 VDD2.t1 1.75374
C0 VP VDD2 0.492254f
C1 VN VDD1 0.151675f
C2 w_n3626_n4676# VN 7.08789f
C3 w_n3626_n4676# VDD1 2.83815f
C4 VP VN 8.51665f
C5 VP VDD1 10.7745f
C6 B VTAIL 5.34964f
C7 VP w_n3626_n4676# 7.55776f
C8 B VDD2 2.7999f
C9 VDD2 VTAIL 10.1307f
C10 B VN 1.33031f
C11 VN VTAIL 10.3949f
C12 B VDD1 2.71646f
C13 VDD1 VTAIL 10.0782f
C14 B w_n3626_n4676# 12.0486f
C15 w_n3626_n4676# VTAIL 3.90919f
C16 VP B 2.11678f
C17 VP VTAIL 10.409201f
C18 VDD2 VN 10.438f
C19 VDD2 VDD1 1.56021f
C20 w_n3626_n4676# VDD2 2.93567f
C21 VDD2 VSUBS 2.19364f
C22 VDD1 VSUBS 2.72573f
C23 VTAIL VSUBS 1.511553f
C24 VN VSUBS 6.47349f
C25 VP VSUBS 3.484611f
C26 B VSUBS 5.576251f
C27 w_n3626_n4676# VSUBS 0.207248p
C28 VDD2.t4 VSUBS 4.27979f
C29 VDD2.t0 VSUBS 0.394312f
C30 VDD2.t1 VSUBS 0.394312f
C31 VDD2.n0 VSUBS 3.28874f
C32 VDD2.n1 VSUBS 4.40602f
C33 VDD2.t2 VSUBS 4.25535f
C34 VDD2.n2 VSUBS 4.00818f
C35 VDD2.t5 VSUBS 0.394312f
C36 VDD2.t3 VSUBS 0.394312f
C37 VDD2.n3 VSUBS 3.28868f
C38 VN.t4 VSUBS 3.81175f
C39 VN.n0 VSUBS 1.40753f
C40 VN.n1 VSUBS 0.024985f
C41 VN.n2 VSUBS 0.029727f
C42 VN.n3 VSUBS 0.283644f
C43 VN.t5 VSUBS 3.81175f
C44 VN.t1 VSUBS 4.0821f
C45 VN.n4 VSUBS 1.35133f
C46 VN.n5 VSUBS 1.40845f
C47 VN.n6 VSUBS 0.046333f
C48 VN.n7 VSUBS 0.046766f
C49 VN.n8 VSUBS 0.024985f
C50 VN.n9 VSUBS 0.024985f
C51 VN.n10 VSUBS 0.024985f
C52 VN.n11 VSUBS 0.04248f
C53 VN.n12 VSUBS 0.046333f
C54 VN.n13 VSUBS 0.038098f
C55 VN.n14 VSUBS 0.040319f
C56 VN.n15 VSUBS 0.056334f
C57 VN.t3 VSUBS 3.81175f
C58 VN.n16 VSUBS 1.40753f
C59 VN.n17 VSUBS 0.024985f
C60 VN.n18 VSUBS 0.029727f
C61 VN.n19 VSUBS 0.283644f
C62 VN.t0 VSUBS 3.81175f
C63 VN.t2 VSUBS 4.0821f
C64 VN.n20 VSUBS 1.35133f
C65 VN.n21 VSUBS 1.40845f
C66 VN.n22 VSUBS 0.046333f
C67 VN.n23 VSUBS 0.046766f
C68 VN.n24 VSUBS 0.024985f
C69 VN.n25 VSUBS 0.024985f
C70 VN.n26 VSUBS 0.024985f
C71 VN.n27 VSUBS 0.04248f
C72 VN.n28 VSUBS 0.046333f
C73 VN.n29 VSUBS 0.038098f
C74 VN.n30 VSUBS 0.040319f
C75 VN.n31 VSUBS 1.63764f
C76 VDD1.t4 VSUBS 4.29777f
C77 VDD1.t5 VSUBS 4.29616f
C78 VDD1.t2 VSUBS 0.395821f
C79 VDD1.t3 VSUBS 0.395821f
C80 VDD1.n0 VSUBS 3.30131f
C81 VDD1.n1 VSUBS 4.57311f
C82 VDD1.t1 VSUBS 0.395821f
C83 VDD1.t0 VSUBS 0.395821f
C84 VDD1.n2 VSUBS 3.29296f
C85 VDD1.n3 VSUBS 3.98666f
C86 VTAIL.t4 VSUBS 0.405062f
C87 VTAIL.t2 VSUBS 0.405062f
C88 VTAIL.n0 VSUBS 3.18905f
C89 VTAIL.n1 VSUBS 0.936218f
C90 VTAIL.t9 VSUBS 4.16375f
C91 VTAIL.n2 VSUBS 1.25228f
C92 VTAIL.t5 VSUBS 0.405062f
C93 VTAIL.t6 VSUBS 0.405062f
C94 VTAIL.n3 VSUBS 3.18905f
C95 VTAIL.n4 VSUBS 3.26228f
C96 VTAIL.t3 VSUBS 0.405062f
C97 VTAIL.t1 VSUBS 0.405062f
C98 VTAIL.n5 VSUBS 3.18906f
C99 VTAIL.n6 VSUBS 3.26228f
C100 VTAIL.t0 VSUBS 4.16378f
C101 VTAIL.n7 VSUBS 1.25225f
C102 VTAIL.t8 VSUBS 0.405062f
C103 VTAIL.t7 VSUBS 0.405062f
C104 VTAIL.n8 VSUBS 3.18906f
C105 VTAIL.n9 VSUBS 1.12226f
C106 VTAIL.t10 VSUBS 4.16375f
C107 VTAIL.n10 VSUBS 3.13733f
C108 VTAIL.t11 VSUBS 4.16375f
C109 VTAIL.n11 VSUBS 3.0684f
C110 VP.t2 VSUBS 4.12989f
C111 VP.n0 VSUBS 1.52501f
C112 VP.n1 VSUBS 0.02707f
C113 VP.n2 VSUBS 0.032208f
C114 VP.n3 VSUBS 0.02707f
C115 VP.t3 VSUBS 4.12989f
C116 VP.n4 VSUBS 0.0502f
C117 VP.n5 VSUBS 0.02707f
C118 VP.n6 VSUBS 0.0502f
C119 VP.t5 VSUBS 4.12989f
C120 VP.n7 VSUBS 1.52501f
C121 VP.n8 VSUBS 0.02707f
C122 VP.n9 VSUBS 0.032208f
C123 VP.n10 VSUBS 0.307318f
C124 VP.t4 VSUBS 4.12989f
C125 VP.t1 VSUBS 4.4228f
C126 VP.n11 VSUBS 1.46412f
C127 VP.n12 VSUBS 1.52601f
C128 VP.n13 VSUBS 0.0502f
C129 VP.n14 VSUBS 0.050669f
C130 VP.n15 VSUBS 0.02707f
C131 VP.n16 VSUBS 0.02707f
C132 VP.n17 VSUBS 0.02707f
C133 VP.n18 VSUBS 0.046025f
C134 VP.n19 VSUBS 0.0502f
C135 VP.n20 VSUBS 0.041278f
C136 VP.n21 VSUBS 0.043684f
C137 VP.n22 VSUBS 1.7636f
C138 VP.n23 VSUBS 1.78127f
C139 VP.t0 VSUBS 4.12989f
C140 VP.n24 VSUBS 1.52501f
C141 VP.n25 VSUBS 0.041278f
C142 VP.n26 VSUBS 0.043684f
C143 VP.n27 VSUBS 0.02707f
C144 VP.n28 VSUBS 0.02707f
C145 VP.n29 VSUBS 0.046025f
C146 VP.n30 VSUBS 0.032208f
C147 VP.n31 VSUBS 0.050669f
C148 VP.n32 VSUBS 0.02707f
C149 VP.n33 VSUBS 0.02707f
C150 VP.n34 VSUBS 0.02707f
C151 VP.n35 VSUBS 1.45203f
C152 VP.n36 VSUBS 0.0502f
C153 VP.n37 VSUBS 0.050669f
C154 VP.n38 VSUBS 0.02707f
C155 VP.n39 VSUBS 0.02707f
C156 VP.n40 VSUBS 0.02707f
C157 VP.n41 VSUBS 0.046025f
C158 VP.n42 VSUBS 0.0502f
C159 VP.n43 VSUBS 0.041278f
C160 VP.n44 VSUBS 0.043684f
C161 VP.n45 VSUBS 0.061036f
C162 B.n0 VSUBS 0.004712f
C163 B.n1 VSUBS 0.004712f
C164 B.n2 VSUBS 0.007451f
C165 B.n3 VSUBS 0.007451f
C166 B.n4 VSUBS 0.007451f
C167 B.n5 VSUBS 0.007451f
C168 B.n6 VSUBS 0.007451f
C169 B.n7 VSUBS 0.007451f
C170 B.n8 VSUBS 0.007451f
C171 B.n9 VSUBS 0.007451f
C172 B.n10 VSUBS 0.007451f
C173 B.n11 VSUBS 0.007451f
C174 B.n12 VSUBS 0.007451f
C175 B.n13 VSUBS 0.007451f
C176 B.n14 VSUBS 0.007451f
C177 B.n15 VSUBS 0.007451f
C178 B.n16 VSUBS 0.007451f
C179 B.n17 VSUBS 0.007451f
C180 B.n18 VSUBS 0.007451f
C181 B.n19 VSUBS 0.007451f
C182 B.n20 VSUBS 0.007451f
C183 B.n21 VSUBS 0.007451f
C184 B.n22 VSUBS 0.007451f
C185 B.n23 VSUBS 0.007451f
C186 B.n24 VSUBS 0.007451f
C187 B.n25 VSUBS 0.018117f
C188 B.n26 VSUBS 0.007451f
C189 B.n27 VSUBS 0.007451f
C190 B.n28 VSUBS 0.007451f
C191 B.n29 VSUBS 0.007451f
C192 B.n30 VSUBS 0.007451f
C193 B.n31 VSUBS 0.007451f
C194 B.n32 VSUBS 0.007451f
C195 B.n33 VSUBS 0.007451f
C196 B.n34 VSUBS 0.007451f
C197 B.n35 VSUBS 0.007451f
C198 B.n36 VSUBS 0.007451f
C199 B.n37 VSUBS 0.007451f
C200 B.n38 VSUBS 0.007451f
C201 B.n39 VSUBS 0.007451f
C202 B.n40 VSUBS 0.007451f
C203 B.n41 VSUBS 0.007451f
C204 B.n42 VSUBS 0.007451f
C205 B.n43 VSUBS 0.007451f
C206 B.n44 VSUBS 0.007451f
C207 B.n45 VSUBS 0.007451f
C208 B.n46 VSUBS 0.007451f
C209 B.n47 VSUBS 0.007451f
C210 B.n48 VSUBS 0.007451f
C211 B.n49 VSUBS 0.007451f
C212 B.n50 VSUBS 0.007451f
C213 B.n51 VSUBS 0.007451f
C214 B.n52 VSUBS 0.007451f
C215 B.n53 VSUBS 0.007451f
C216 B.n54 VSUBS 0.007451f
C217 B.n55 VSUBS 0.007451f
C218 B.t11 VSUBS 0.667626f
C219 B.t10 VSUBS 0.692739f
C220 B.t9 VSUBS 2.63927f
C221 B.n56 VSUBS 0.401719f
C222 B.n57 VSUBS 0.078494f
C223 B.n58 VSUBS 0.017264f
C224 B.n59 VSUBS 0.007451f
C225 B.n60 VSUBS 0.007451f
C226 B.n61 VSUBS 0.007451f
C227 B.n62 VSUBS 0.007451f
C228 B.n63 VSUBS 0.007451f
C229 B.t5 VSUBS 0.667601f
C230 B.t4 VSUBS 0.692719f
C231 B.t3 VSUBS 2.63927f
C232 B.n64 VSUBS 0.401739f
C233 B.n65 VSUBS 0.078519f
C234 B.n66 VSUBS 0.007451f
C235 B.n67 VSUBS 0.007451f
C236 B.n68 VSUBS 0.007451f
C237 B.n69 VSUBS 0.007451f
C238 B.n70 VSUBS 0.007451f
C239 B.n71 VSUBS 0.007451f
C240 B.n72 VSUBS 0.007451f
C241 B.n73 VSUBS 0.007451f
C242 B.n74 VSUBS 0.007451f
C243 B.n75 VSUBS 0.007451f
C244 B.n76 VSUBS 0.007451f
C245 B.n77 VSUBS 0.007451f
C246 B.n78 VSUBS 0.007451f
C247 B.n79 VSUBS 0.007451f
C248 B.n80 VSUBS 0.007451f
C249 B.n81 VSUBS 0.007451f
C250 B.n82 VSUBS 0.007451f
C251 B.n83 VSUBS 0.007451f
C252 B.n84 VSUBS 0.007451f
C253 B.n85 VSUBS 0.007451f
C254 B.n86 VSUBS 0.007451f
C255 B.n87 VSUBS 0.007451f
C256 B.n88 VSUBS 0.007451f
C257 B.n89 VSUBS 0.007451f
C258 B.n90 VSUBS 0.007451f
C259 B.n91 VSUBS 0.007451f
C260 B.n92 VSUBS 0.007451f
C261 B.n93 VSUBS 0.007451f
C262 B.n94 VSUBS 0.007451f
C263 B.n95 VSUBS 0.018921f
C264 B.n96 VSUBS 0.007451f
C265 B.n97 VSUBS 0.007451f
C266 B.n98 VSUBS 0.007451f
C267 B.n99 VSUBS 0.007451f
C268 B.n100 VSUBS 0.007451f
C269 B.n101 VSUBS 0.007451f
C270 B.n102 VSUBS 0.007451f
C271 B.n103 VSUBS 0.007451f
C272 B.n104 VSUBS 0.007451f
C273 B.n105 VSUBS 0.007451f
C274 B.n106 VSUBS 0.007451f
C275 B.n107 VSUBS 0.007451f
C276 B.n108 VSUBS 0.007451f
C277 B.n109 VSUBS 0.007451f
C278 B.n110 VSUBS 0.007451f
C279 B.n111 VSUBS 0.007451f
C280 B.n112 VSUBS 0.007451f
C281 B.n113 VSUBS 0.007451f
C282 B.n114 VSUBS 0.007451f
C283 B.n115 VSUBS 0.007451f
C284 B.n116 VSUBS 0.007451f
C285 B.n117 VSUBS 0.007451f
C286 B.n118 VSUBS 0.007451f
C287 B.n119 VSUBS 0.007451f
C288 B.n120 VSUBS 0.007451f
C289 B.n121 VSUBS 0.007451f
C290 B.n122 VSUBS 0.007451f
C291 B.n123 VSUBS 0.007451f
C292 B.n124 VSUBS 0.007451f
C293 B.n125 VSUBS 0.007451f
C294 B.n126 VSUBS 0.007451f
C295 B.n127 VSUBS 0.007451f
C296 B.n128 VSUBS 0.007451f
C297 B.n129 VSUBS 0.007451f
C298 B.n130 VSUBS 0.007451f
C299 B.n131 VSUBS 0.007451f
C300 B.n132 VSUBS 0.007451f
C301 B.n133 VSUBS 0.007451f
C302 B.n134 VSUBS 0.007451f
C303 B.n135 VSUBS 0.007451f
C304 B.n136 VSUBS 0.007451f
C305 B.n137 VSUBS 0.007451f
C306 B.n138 VSUBS 0.007451f
C307 B.n139 VSUBS 0.007451f
C308 B.n140 VSUBS 0.007451f
C309 B.n141 VSUBS 0.007451f
C310 B.n142 VSUBS 0.007451f
C311 B.n143 VSUBS 0.018921f
C312 B.n144 VSUBS 0.007451f
C313 B.n145 VSUBS 0.007451f
C314 B.n146 VSUBS 0.007451f
C315 B.n147 VSUBS 0.007451f
C316 B.n148 VSUBS 0.007451f
C317 B.n149 VSUBS 0.007451f
C318 B.n150 VSUBS 0.007451f
C319 B.n151 VSUBS 0.007451f
C320 B.n152 VSUBS 0.007451f
C321 B.n153 VSUBS 0.007451f
C322 B.n154 VSUBS 0.007451f
C323 B.n155 VSUBS 0.007451f
C324 B.n156 VSUBS 0.007451f
C325 B.n157 VSUBS 0.007451f
C326 B.n158 VSUBS 0.007451f
C327 B.n159 VSUBS 0.007451f
C328 B.n160 VSUBS 0.007451f
C329 B.n161 VSUBS 0.007451f
C330 B.n162 VSUBS 0.007451f
C331 B.n163 VSUBS 0.007451f
C332 B.n164 VSUBS 0.007451f
C333 B.n165 VSUBS 0.007451f
C334 B.n166 VSUBS 0.007451f
C335 B.n167 VSUBS 0.007451f
C336 B.n168 VSUBS 0.007451f
C337 B.n169 VSUBS 0.007451f
C338 B.n170 VSUBS 0.007451f
C339 B.n171 VSUBS 0.007451f
C340 B.n172 VSUBS 0.007451f
C341 B.n173 VSUBS 0.007451f
C342 B.t1 VSUBS 0.667601f
C343 B.t2 VSUBS 0.692719f
C344 B.t0 VSUBS 2.63927f
C345 B.n174 VSUBS 0.401739f
C346 B.n175 VSUBS 0.078519f
C347 B.n176 VSUBS 0.007451f
C348 B.n177 VSUBS 0.007451f
C349 B.n178 VSUBS 0.007451f
C350 B.n179 VSUBS 0.007451f
C351 B.t7 VSUBS 0.667626f
C352 B.t8 VSUBS 0.692739f
C353 B.t6 VSUBS 2.63927f
C354 B.n180 VSUBS 0.401719f
C355 B.n181 VSUBS 0.078494f
C356 B.n182 VSUBS 0.017264f
C357 B.n183 VSUBS 0.007451f
C358 B.n184 VSUBS 0.007451f
C359 B.n185 VSUBS 0.007451f
C360 B.n186 VSUBS 0.007451f
C361 B.n187 VSUBS 0.007451f
C362 B.n188 VSUBS 0.007451f
C363 B.n189 VSUBS 0.007451f
C364 B.n190 VSUBS 0.007451f
C365 B.n191 VSUBS 0.007451f
C366 B.n192 VSUBS 0.007451f
C367 B.n193 VSUBS 0.007451f
C368 B.n194 VSUBS 0.007451f
C369 B.n195 VSUBS 0.007451f
C370 B.n196 VSUBS 0.007451f
C371 B.n197 VSUBS 0.007451f
C372 B.n198 VSUBS 0.007451f
C373 B.n199 VSUBS 0.007451f
C374 B.n200 VSUBS 0.007451f
C375 B.n201 VSUBS 0.007451f
C376 B.n202 VSUBS 0.007451f
C377 B.n203 VSUBS 0.007451f
C378 B.n204 VSUBS 0.007451f
C379 B.n205 VSUBS 0.007451f
C380 B.n206 VSUBS 0.007451f
C381 B.n207 VSUBS 0.007451f
C382 B.n208 VSUBS 0.007451f
C383 B.n209 VSUBS 0.007451f
C384 B.n210 VSUBS 0.007451f
C385 B.n211 VSUBS 0.007451f
C386 B.n212 VSUBS 0.007451f
C387 B.n213 VSUBS 0.018117f
C388 B.n214 VSUBS 0.007451f
C389 B.n215 VSUBS 0.007451f
C390 B.n216 VSUBS 0.007451f
C391 B.n217 VSUBS 0.007451f
C392 B.n218 VSUBS 0.007451f
C393 B.n219 VSUBS 0.007451f
C394 B.n220 VSUBS 0.007451f
C395 B.n221 VSUBS 0.007451f
C396 B.n222 VSUBS 0.007451f
C397 B.n223 VSUBS 0.007451f
C398 B.n224 VSUBS 0.007451f
C399 B.n225 VSUBS 0.007451f
C400 B.n226 VSUBS 0.007451f
C401 B.n227 VSUBS 0.007451f
C402 B.n228 VSUBS 0.007451f
C403 B.n229 VSUBS 0.007451f
C404 B.n230 VSUBS 0.007451f
C405 B.n231 VSUBS 0.007451f
C406 B.n232 VSUBS 0.007451f
C407 B.n233 VSUBS 0.007451f
C408 B.n234 VSUBS 0.007451f
C409 B.n235 VSUBS 0.007451f
C410 B.n236 VSUBS 0.007451f
C411 B.n237 VSUBS 0.007451f
C412 B.n238 VSUBS 0.007451f
C413 B.n239 VSUBS 0.007451f
C414 B.n240 VSUBS 0.007451f
C415 B.n241 VSUBS 0.007451f
C416 B.n242 VSUBS 0.007451f
C417 B.n243 VSUBS 0.007451f
C418 B.n244 VSUBS 0.007451f
C419 B.n245 VSUBS 0.007451f
C420 B.n246 VSUBS 0.007451f
C421 B.n247 VSUBS 0.007451f
C422 B.n248 VSUBS 0.007451f
C423 B.n249 VSUBS 0.007451f
C424 B.n250 VSUBS 0.007451f
C425 B.n251 VSUBS 0.007451f
C426 B.n252 VSUBS 0.007451f
C427 B.n253 VSUBS 0.007451f
C428 B.n254 VSUBS 0.007451f
C429 B.n255 VSUBS 0.007451f
C430 B.n256 VSUBS 0.007451f
C431 B.n257 VSUBS 0.007451f
C432 B.n258 VSUBS 0.007451f
C433 B.n259 VSUBS 0.007451f
C434 B.n260 VSUBS 0.007451f
C435 B.n261 VSUBS 0.007451f
C436 B.n262 VSUBS 0.007451f
C437 B.n263 VSUBS 0.007451f
C438 B.n264 VSUBS 0.007451f
C439 B.n265 VSUBS 0.007451f
C440 B.n266 VSUBS 0.007451f
C441 B.n267 VSUBS 0.007451f
C442 B.n268 VSUBS 0.007451f
C443 B.n269 VSUBS 0.007451f
C444 B.n270 VSUBS 0.007451f
C445 B.n271 VSUBS 0.007451f
C446 B.n272 VSUBS 0.007451f
C447 B.n273 VSUBS 0.007451f
C448 B.n274 VSUBS 0.007451f
C449 B.n275 VSUBS 0.007451f
C450 B.n276 VSUBS 0.007451f
C451 B.n277 VSUBS 0.007451f
C452 B.n278 VSUBS 0.007451f
C453 B.n279 VSUBS 0.007451f
C454 B.n280 VSUBS 0.007451f
C455 B.n281 VSUBS 0.007451f
C456 B.n282 VSUBS 0.007451f
C457 B.n283 VSUBS 0.007451f
C458 B.n284 VSUBS 0.007451f
C459 B.n285 VSUBS 0.007451f
C460 B.n286 VSUBS 0.007451f
C461 B.n287 VSUBS 0.007451f
C462 B.n288 VSUBS 0.007451f
C463 B.n289 VSUBS 0.007451f
C464 B.n290 VSUBS 0.007451f
C465 B.n291 VSUBS 0.007451f
C466 B.n292 VSUBS 0.007451f
C467 B.n293 VSUBS 0.007451f
C468 B.n294 VSUBS 0.007451f
C469 B.n295 VSUBS 0.007451f
C470 B.n296 VSUBS 0.007451f
C471 B.n297 VSUBS 0.007451f
C472 B.n298 VSUBS 0.007451f
C473 B.n299 VSUBS 0.007451f
C474 B.n300 VSUBS 0.007451f
C475 B.n301 VSUBS 0.007451f
C476 B.n302 VSUBS 0.007451f
C477 B.n303 VSUBS 0.007451f
C478 B.n304 VSUBS 0.018117f
C479 B.n305 VSUBS 0.018921f
C480 B.n306 VSUBS 0.018921f
C481 B.n307 VSUBS 0.007451f
C482 B.n308 VSUBS 0.007451f
C483 B.n309 VSUBS 0.007451f
C484 B.n310 VSUBS 0.007451f
C485 B.n311 VSUBS 0.007451f
C486 B.n312 VSUBS 0.007451f
C487 B.n313 VSUBS 0.007451f
C488 B.n314 VSUBS 0.007451f
C489 B.n315 VSUBS 0.007451f
C490 B.n316 VSUBS 0.007451f
C491 B.n317 VSUBS 0.007451f
C492 B.n318 VSUBS 0.007451f
C493 B.n319 VSUBS 0.007451f
C494 B.n320 VSUBS 0.007451f
C495 B.n321 VSUBS 0.007451f
C496 B.n322 VSUBS 0.007451f
C497 B.n323 VSUBS 0.007451f
C498 B.n324 VSUBS 0.007451f
C499 B.n325 VSUBS 0.007451f
C500 B.n326 VSUBS 0.007451f
C501 B.n327 VSUBS 0.007451f
C502 B.n328 VSUBS 0.007451f
C503 B.n329 VSUBS 0.007451f
C504 B.n330 VSUBS 0.007451f
C505 B.n331 VSUBS 0.007451f
C506 B.n332 VSUBS 0.007451f
C507 B.n333 VSUBS 0.007451f
C508 B.n334 VSUBS 0.007451f
C509 B.n335 VSUBS 0.007451f
C510 B.n336 VSUBS 0.007451f
C511 B.n337 VSUBS 0.007451f
C512 B.n338 VSUBS 0.007451f
C513 B.n339 VSUBS 0.007451f
C514 B.n340 VSUBS 0.007451f
C515 B.n341 VSUBS 0.007451f
C516 B.n342 VSUBS 0.007451f
C517 B.n343 VSUBS 0.007451f
C518 B.n344 VSUBS 0.007451f
C519 B.n345 VSUBS 0.007451f
C520 B.n346 VSUBS 0.007451f
C521 B.n347 VSUBS 0.007451f
C522 B.n348 VSUBS 0.007451f
C523 B.n349 VSUBS 0.007451f
C524 B.n350 VSUBS 0.007451f
C525 B.n351 VSUBS 0.007451f
C526 B.n352 VSUBS 0.007451f
C527 B.n353 VSUBS 0.007451f
C528 B.n354 VSUBS 0.007451f
C529 B.n355 VSUBS 0.007451f
C530 B.n356 VSUBS 0.007451f
C531 B.n357 VSUBS 0.007451f
C532 B.n358 VSUBS 0.007451f
C533 B.n359 VSUBS 0.007451f
C534 B.n360 VSUBS 0.007451f
C535 B.n361 VSUBS 0.007451f
C536 B.n362 VSUBS 0.007451f
C537 B.n363 VSUBS 0.007451f
C538 B.n364 VSUBS 0.007451f
C539 B.n365 VSUBS 0.007451f
C540 B.n366 VSUBS 0.007451f
C541 B.n367 VSUBS 0.007451f
C542 B.n368 VSUBS 0.007451f
C543 B.n369 VSUBS 0.007451f
C544 B.n370 VSUBS 0.007451f
C545 B.n371 VSUBS 0.007451f
C546 B.n372 VSUBS 0.007451f
C547 B.n373 VSUBS 0.007451f
C548 B.n374 VSUBS 0.007451f
C549 B.n375 VSUBS 0.007451f
C550 B.n376 VSUBS 0.007451f
C551 B.n377 VSUBS 0.007451f
C552 B.n378 VSUBS 0.007451f
C553 B.n379 VSUBS 0.007451f
C554 B.n380 VSUBS 0.007451f
C555 B.n381 VSUBS 0.007451f
C556 B.n382 VSUBS 0.007451f
C557 B.n383 VSUBS 0.007451f
C558 B.n384 VSUBS 0.007451f
C559 B.n385 VSUBS 0.007451f
C560 B.n386 VSUBS 0.007451f
C561 B.n387 VSUBS 0.007451f
C562 B.n388 VSUBS 0.007451f
C563 B.n389 VSUBS 0.007451f
C564 B.n390 VSUBS 0.007451f
C565 B.n391 VSUBS 0.007451f
C566 B.n392 VSUBS 0.007451f
C567 B.n393 VSUBS 0.007451f
C568 B.n394 VSUBS 0.007451f
C569 B.n395 VSUBS 0.00515f
C570 B.n396 VSUBS 0.007451f
C571 B.n397 VSUBS 0.007451f
C572 B.n398 VSUBS 0.006027f
C573 B.n399 VSUBS 0.007451f
C574 B.n400 VSUBS 0.007451f
C575 B.n401 VSUBS 0.007451f
C576 B.n402 VSUBS 0.007451f
C577 B.n403 VSUBS 0.007451f
C578 B.n404 VSUBS 0.007451f
C579 B.n405 VSUBS 0.007451f
C580 B.n406 VSUBS 0.007451f
C581 B.n407 VSUBS 0.007451f
C582 B.n408 VSUBS 0.007451f
C583 B.n409 VSUBS 0.007451f
C584 B.n410 VSUBS 0.006027f
C585 B.n411 VSUBS 0.017264f
C586 B.n412 VSUBS 0.00515f
C587 B.n413 VSUBS 0.007451f
C588 B.n414 VSUBS 0.007451f
C589 B.n415 VSUBS 0.007451f
C590 B.n416 VSUBS 0.007451f
C591 B.n417 VSUBS 0.007451f
C592 B.n418 VSUBS 0.007451f
C593 B.n419 VSUBS 0.007451f
C594 B.n420 VSUBS 0.007451f
C595 B.n421 VSUBS 0.007451f
C596 B.n422 VSUBS 0.007451f
C597 B.n423 VSUBS 0.007451f
C598 B.n424 VSUBS 0.007451f
C599 B.n425 VSUBS 0.007451f
C600 B.n426 VSUBS 0.007451f
C601 B.n427 VSUBS 0.007451f
C602 B.n428 VSUBS 0.007451f
C603 B.n429 VSUBS 0.007451f
C604 B.n430 VSUBS 0.007451f
C605 B.n431 VSUBS 0.007451f
C606 B.n432 VSUBS 0.007451f
C607 B.n433 VSUBS 0.007451f
C608 B.n434 VSUBS 0.007451f
C609 B.n435 VSUBS 0.007451f
C610 B.n436 VSUBS 0.007451f
C611 B.n437 VSUBS 0.007451f
C612 B.n438 VSUBS 0.007451f
C613 B.n439 VSUBS 0.007451f
C614 B.n440 VSUBS 0.007451f
C615 B.n441 VSUBS 0.007451f
C616 B.n442 VSUBS 0.007451f
C617 B.n443 VSUBS 0.007451f
C618 B.n444 VSUBS 0.007451f
C619 B.n445 VSUBS 0.007451f
C620 B.n446 VSUBS 0.007451f
C621 B.n447 VSUBS 0.007451f
C622 B.n448 VSUBS 0.007451f
C623 B.n449 VSUBS 0.007451f
C624 B.n450 VSUBS 0.007451f
C625 B.n451 VSUBS 0.007451f
C626 B.n452 VSUBS 0.007451f
C627 B.n453 VSUBS 0.007451f
C628 B.n454 VSUBS 0.007451f
C629 B.n455 VSUBS 0.007451f
C630 B.n456 VSUBS 0.007451f
C631 B.n457 VSUBS 0.007451f
C632 B.n458 VSUBS 0.007451f
C633 B.n459 VSUBS 0.007451f
C634 B.n460 VSUBS 0.007451f
C635 B.n461 VSUBS 0.007451f
C636 B.n462 VSUBS 0.007451f
C637 B.n463 VSUBS 0.007451f
C638 B.n464 VSUBS 0.007451f
C639 B.n465 VSUBS 0.007451f
C640 B.n466 VSUBS 0.007451f
C641 B.n467 VSUBS 0.007451f
C642 B.n468 VSUBS 0.007451f
C643 B.n469 VSUBS 0.007451f
C644 B.n470 VSUBS 0.007451f
C645 B.n471 VSUBS 0.007451f
C646 B.n472 VSUBS 0.007451f
C647 B.n473 VSUBS 0.007451f
C648 B.n474 VSUBS 0.007451f
C649 B.n475 VSUBS 0.007451f
C650 B.n476 VSUBS 0.007451f
C651 B.n477 VSUBS 0.007451f
C652 B.n478 VSUBS 0.007451f
C653 B.n479 VSUBS 0.007451f
C654 B.n480 VSUBS 0.007451f
C655 B.n481 VSUBS 0.007451f
C656 B.n482 VSUBS 0.007451f
C657 B.n483 VSUBS 0.007451f
C658 B.n484 VSUBS 0.007451f
C659 B.n485 VSUBS 0.007451f
C660 B.n486 VSUBS 0.007451f
C661 B.n487 VSUBS 0.007451f
C662 B.n488 VSUBS 0.007451f
C663 B.n489 VSUBS 0.007451f
C664 B.n490 VSUBS 0.007451f
C665 B.n491 VSUBS 0.007451f
C666 B.n492 VSUBS 0.007451f
C667 B.n493 VSUBS 0.007451f
C668 B.n494 VSUBS 0.007451f
C669 B.n495 VSUBS 0.007451f
C670 B.n496 VSUBS 0.007451f
C671 B.n497 VSUBS 0.007451f
C672 B.n498 VSUBS 0.007451f
C673 B.n499 VSUBS 0.007451f
C674 B.n500 VSUBS 0.007451f
C675 B.n501 VSUBS 0.007451f
C676 B.n502 VSUBS 0.018921f
C677 B.n503 VSUBS 0.018117f
C678 B.n504 VSUBS 0.018117f
C679 B.n505 VSUBS 0.007451f
C680 B.n506 VSUBS 0.007451f
C681 B.n507 VSUBS 0.007451f
C682 B.n508 VSUBS 0.007451f
C683 B.n509 VSUBS 0.007451f
C684 B.n510 VSUBS 0.007451f
C685 B.n511 VSUBS 0.007451f
C686 B.n512 VSUBS 0.007451f
C687 B.n513 VSUBS 0.007451f
C688 B.n514 VSUBS 0.007451f
C689 B.n515 VSUBS 0.007451f
C690 B.n516 VSUBS 0.007451f
C691 B.n517 VSUBS 0.007451f
C692 B.n518 VSUBS 0.007451f
C693 B.n519 VSUBS 0.007451f
C694 B.n520 VSUBS 0.007451f
C695 B.n521 VSUBS 0.007451f
C696 B.n522 VSUBS 0.007451f
C697 B.n523 VSUBS 0.007451f
C698 B.n524 VSUBS 0.007451f
C699 B.n525 VSUBS 0.007451f
C700 B.n526 VSUBS 0.007451f
C701 B.n527 VSUBS 0.007451f
C702 B.n528 VSUBS 0.007451f
C703 B.n529 VSUBS 0.007451f
C704 B.n530 VSUBS 0.007451f
C705 B.n531 VSUBS 0.007451f
C706 B.n532 VSUBS 0.007451f
C707 B.n533 VSUBS 0.007451f
C708 B.n534 VSUBS 0.007451f
C709 B.n535 VSUBS 0.007451f
C710 B.n536 VSUBS 0.007451f
C711 B.n537 VSUBS 0.007451f
C712 B.n538 VSUBS 0.007451f
C713 B.n539 VSUBS 0.007451f
C714 B.n540 VSUBS 0.007451f
C715 B.n541 VSUBS 0.007451f
C716 B.n542 VSUBS 0.007451f
C717 B.n543 VSUBS 0.007451f
C718 B.n544 VSUBS 0.007451f
C719 B.n545 VSUBS 0.007451f
C720 B.n546 VSUBS 0.007451f
C721 B.n547 VSUBS 0.007451f
C722 B.n548 VSUBS 0.007451f
C723 B.n549 VSUBS 0.007451f
C724 B.n550 VSUBS 0.007451f
C725 B.n551 VSUBS 0.007451f
C726 B.n552 VSUBS 0.007451f
C727 B.n553 VSUBS 0.007451f
C728 B.n554 VSUBS 0.007451f
C729 B.n555 VSUBS 0.007451f
C730 B.n556 VSUBS 0.007451f
C731 B.n557 VSUBS 0.007451f
C732 B.n558 VSUBS 0.007451f
C733 B.n559 VSUBS 0.007451f
C734 B.n560 VSUBS 0.007451f
C735 B.n561 VSUBS 0.007451f
C736 B.n562 VSUBS 0.007451f
C737 B.n563 VSUBS 0.007451f
C738 B.n564 VSUBS 0.007451f
C739 B.n565 VSUBS 0.007451f
C740 B.n566 VSUBS 0.007451f
C741 B.n567 VSUBS 0.007451f
C742 B.n568 VSUBS 0.007451f
C743 B.n569 VSUBS 0.007451f
C744 B.n570 VSUBS 0.007451f
C745 B.n571 VSUBS 0.007451f
C746 B.n572 VSUBS 0.007451f
C747 B.n573 VSUBS 0.007451f
C748 B.n574 VSUBS 0.007451f
C749 B.n575 VSUBS 0.007451f
C750 B.n576 VSUBS 0.007451f
C751 B.n577 VSUBS 0.007451f
C752 B.n578 VSUBS 0.007451f
C753 B.n579 VSUBS 0.007451f
C754 B.n580 VSUBS 0.007451f
C755 B.n581 VSUBS 0.007451f
C756 B.n582 VSUBS 0.007451f
C757 B.n583 VSUBS 0.007451f
C758 B.n584 VSUBS 0.007451f
C759 B.n585 VSUBS 0.007451f
C760 B.n586 VSUBS 0.007451f
C761 B.n587 VSUBS 0.007451f
C762 B.n588 VSUBS 0.007451f
C763 B.n589 VSUBS 0.007451f
C764 B.n590 VSUBS 0.007451f
C765 B.n591 VSUBS 0.007451f
C766 B.n592 VSUBS 0.007451f
C767 B.n593 VSUBS 0.007451f
C768 B.n594 VSUBS 0.007451f
C769 B.n595 VSUBS 0.007451f
C770 B.n596 VSUBS 0.007451f
C771 B.n597 VSUBS 0.007451f
C772 B.n598 VSUBS 0.007451f
C773 B.n599 VSUBS 0.007451f
C774 B.n600 VSUBS 0.007451f
C775 B.n601 VSUBS 0.007451f
C776 B.n602 VSUBS 0.007451f
C777 B.n603 VSUBS 0.007451f
C778 B.n604 VSUBS 0.007451f
C779 B.n605 VSUBS 0.007451f
C780 B.n606 VSUBS 0.007451f
C781 B.n607 VSUBS 0.007451f
C782 B.n608 VSUBS 0.007451f
C783 B.n609 VSUBS 0.007451f
C784 B.n610 VSUBS 0.007451f
C785 B.n611 VSUBS 0.007451f
C786 B.n612 VSUBS 0.007451f
C787 B.n613 VSUBS 0.007451f
C788 B.n614 VSUBS 0.007451f
C789 B.n615 VSUBS 0.007451f
C790 B.n616 VSUBS 0.007451f
C791 B.n617 VSUBS 0.007451f
C792 B.n618 VSUBS 0.007451f
C793 B.n619 VSUBS 0.007451f
C794 B.n620 VSUBS 0.007451f
C795 B.n621 VSUBS 0.007451f
C796 B.n622 VSUBS 0.007451f
C797 B.n623 VSUBS 0.007451f
C798 B.n624 VSUBS 0.007451f
C799 B.n625 VSUBS 0.007451f
C800 B.n626 VSUBS 0.007451f
C801 B.n627 VSUBS 0.007451f
C802 B.n628 VSUBS 0.007451f
C803 B.n629 VSUBS 0.007451f
C804 B.n630 VSUBS 0.007451f
C805 B.n631 VSUBS 0.007451f
C806 B.n632 VSUBS 0.007451f
C807 B.n633 VSUBS 0.007451f
C808 B.n634 VSUBS 0.007451f
C809 B.n635 VSUBS 0.007451f
C810 B.n636 VSUBS 0.007451f
C811 B.n637 VSUBS 0.007451f
C812 B.n638 VSUBS 0.007451f
C813 B.n639 VSUBS 0.007451f
C814 B.n640 VSUBS 0.007451f
C815 B.n641 VSUBS 0.007451f
C816 B.n642 VSUBS 0.007451f
C817 B.n643 VSUBS 0.007451f
C818 B.n644 VSUBS 0.018117f
C819 B.n645 VSUBS 0.018921f
C820 B.n646 VSUBS 0.018117f
C821 B.n647 VSUBS 0.007451f
C822 B.n648 VSUBS 0.007451f
C823 B.n649 VSUBS 0.007451f
C824 B.n650 VSUBS 0.007451f
C825 B.n651 VSUBS 0.007451f
C826 B.n652 VSUBS 0.007451f
C827 B.n653 VSUBS 0.007451f
C828 B.n654 VSUBS 0.007451f
C829 B.n655 VSUBS 0.007451f
C830 B.n656 VSUBS 0.007451f
C831 B.n657 VSUBS 0.007451f
C832 B.n658 VSUBS 0.007451f
C833 B.n659 VSUBS 0.007451f
C834 B.n660 VSUBS 0.007451f
C835 B.n661 VSUBS 0.007451f
C836 B.n662 VSUBS 0.007451f
C837 B.n663 VSUBS 0.007451f
C838 B.n664 VSUBS 0.007451f
C839 B.n665 VSUBS 0.007451f
C840 B.n666 VSUBS 0.007451f
C841 B.n667 VSUBS 0.007451f
C842 B.n668 VSUBS 0.007451f
C843 B.n669 VSUBS 0.007451f
C844 B.n670 VSUBS 0.007451f
C845 B.n671 VSUBS 0.007451f
C846 B.n672 VSUBS 0.007451f
C847 B.n673 VSUBS 0.007451f
C848 B.n674 VSUBS 0.007451f
C849 B.n675 VSUBS 0.007451f
C850 B.n676 VSUBS 0.007451f
C851 B.n677 VSUBS 0.007451f
C852 B.n678 VSUBS 0.007451f
C853 B.n679 VSUBS 0.007451f
C854 B.n680 VSUBS 0.007451f
C855 B.n681 VSUBS 0.007451f
C856 B.n682 VSUBS 0.007451f
C857 B.n683 VSUBS 0.007451f
C858 B.n684 VSUBS 0.007451f
C859 B.n685 VSUBS 0.007451f
C860 B.n686 VSUBS 0.007451f
C861 B.n687 VSUBS 0.007451f
C862 B.n688 VSUBS 0.007451f
C863 B.n689 VSUBS 0.007451f
C864 B.n690 VSUBS 0.007451f
C865 B.n691 VSUBS 0.007451f
C866 B.n692 VSUBS 0.007451f
C867 B.n693 VSUBS 0.007451f
C868 B.n694 VSUBS 0.007451f
C869 B.n695 VSUBS 0.007451f
C870 B.n696 VSUBS 0.007451f
C871 B.n697 VSUBS 0.007451f
C872 B.n698 VSUBS 0.007451f
C873 B.n699 VSUBS 0.007451f
C874 B.n700 VSUBS 0.007451f
C875 B.n701 VSUBS 0.007451f
C876 B.n702 VSUBS 0.007451f
C877 B.n703 VSUBS 0.007451f
C878 B.n704 VSUBS 0.007451f
C879 B.n705 VSUBS 0.007451f
C880 B.n706 VSUBS 0.007451f
C881 B.n707 VSUBS 0.007451f
C882 B.n708 VSUBS 0.007451f
C883 B.n709 VSUBS 0.007451f
C884 B.n710 VSUBS 0.007451f
C885 B.n711 VSUBS 0.007451f
C886 B.n712 VSUBS 0.007451f
C887 B.n713 VSUBS 0.007451f
C888 B.n714 VSUBS 0.007451f
C889 B.n715 VSUBS 0.007451f
C890 B.n716 VSUBS 0.007451f
C891 B.n717 VSUBS 0.007451f
C892 B.n718 VSUBS 0.007451f
C893 B.n719 VSUBS 0.007451f
C894 B.n720 VSUBS 0.007451f
C895 B.n721 VSUBS 0.007451f
C896 B.n722 VSUBS 0.007451f
C897 B.n723 VSUBS 0.007451f
C898 B.n724 VSUBS 0.007451f
C899 B.n725 VSUBS 0.007451f
C900 B.n726 VSUBS 0.007451f
C901 B.n727 VSUBS 0.007451f
C902 B.n728 VSUBS 0.007451f
C903 B.n729 VSUBS 0.007451f
C904 B.n730 VSUBS 0.007451f
C905 B.n731 VSUBS 0.007451f
C906 B.n732 VSUBS 0.007451f
C907 B.n733 VSUBS 0.007451f
C908 B.n734 VSUBS 0.007451f
C909 B.n735 VSUBS 0.007451f
C910 B.n736 VSUBS 0.00515f
C911 B.n737 VSUBS 0.017264f
C912 B.n738 VSUBS 0.006027f
C913 B.n739 VSUBS 0.007451f
C914 B.n740 VSUBS 0.007451f
C915 B.n741 VSUBS 0.007451f
C916 B.n742 VSUBS 0.007451f
C917 B.n743 VSUBS 0.007451f
C918 B.n744 VSUBS 0.007451f
C919 B.n745 VSUBS 0.007451f
C920 B.n746 VSUBS 0.007451f
C921 B.n747 VSUBS 0.007451f
C922 B.n748 VSUBS 0.007451f
C923 B.n749 VSUBS 0.007451f
C924 B.n750 VSUBS 0.006027f
C925 B.n751 VSUBS 0.007451f
C926 B.n752 VSUBS 0.007451f
C927 B.n753 VSUBS 0.00515f
C928 B.n754 VSUBS 0.007451f
C929 B.n755 VSUBS 0.007451f
C930 B.n756 VSUBS 0.007451f
C931 B.n757 VSUBS 0.007451f
C932 B.n758 VSUBS 0.007451f
C933 B.n759 VSUBS 0.007451f
C934 B.n760 VSUBS 0.007451f
C935 B.n761 VSUBS 0.007451f
C936 B.n762 VSUBS 0.007451f
C937 B.n763 VSUBS 0.007451f
C938 B.n764 VSUBS 0.007451f
C939 B.n765 VSUBS 0.007451f
C940 B.n766 VSUBS 0.007451f
C941 B.n767 VSUBS 0.007451f
C942 B.n768 VSUBS 0.007451f
C943 B.n769 VSUBS 0.007451f
C944 B.n770 VSUBS 0.007451f
C945 B.n771 VSUBS 0.007451f
C946 B.n772 VSUBS 0.007451f
C947 B.n773 VSUBS 0.007451f
C948 B.n774 VSUBS 0.007451f
C949 B.n775 VSUBS 0.007451f
C950 B.n776 VSUBS 0.007451f
C951 B.n777 VSUBS 0.007451f
C952 B.n778 VSUBS 0.007451f
C953 B.n779 VSUBS 0.007451f
C954 B.n780 VSUBS 0.007451f
C955 B.n781 VSUBS 0.007451f
C956 B.n782 VSUBS 0.007451f
C957 B.n783 VSUBS 0.007451f
C958 B.n784 VSUBS 0.007451f
C959 B.n785 VSUBS 0.007451f
C960 B.n786 VSUBS 0.007451f
C961 B.n787 VSUBS 0.007451f
C962 B.n788 VSUBS 0.007451f
C963 B.n789 VSUBS 0.007451f
C964 B.n790 VSUBS 0.007451f
C965 B.n791 VSUBS 0.007451f
C966 B.n792 VSUBS 0.007451f
C967 B.n793 VSUBS 0.007451f
C968 B.n794 VSUBS 0.007451f
C969 B.n795 VSUBS 0.007451f
C970 B.n796 VSUBS 0.007451f
C971 B.n797 VSUBS 0.007451f
C972 B.n798 VSUBS 0.007451f
C973 B.n799 VSUBS 0.007451f
C974 B.n800 VSUBS 0.007451f
C975 B.n801 VSUBS 0.007451f
C976 B.n802 VSUBS 0.007451f
C977 B.n803 VSUBS 0.007451f
C978 B.n804 VSUBS 0.007451f
C979 B.n805 VSUBS 0.007451f
C980 B.n806 VSUBS 0.007451f
C981 B.n807 VSUBS 0.007451f
C982 B.n808 VSUBS 0.007451f
C983 B.n809 VSUBS 0.007451f
C984 B.n810 VSUBS 0.007451f
C985 B.n811 VSUBS 0.007451f
C986 B.n812 VSUBS 0.007451f
C987 B.n813 VSUBS 0.007451f
C988 B.n814 VSUBS 0.007451f
C989 B.n815 VSUBS 0.007451f
C990 B.n816 VSUBS 0.007451f
C991 B.n817 VSUBS 0.007451f
C992 B.n818 VSUBS 0.007451f
C993 B.n819 VSUBS 0.007451f
C994 B.n820 VSUBS 0.007451f
C995 B.n821 VSUBS 0.007451f
C996 B.n822 VSUBS 0.007451f
C997 B.n823 VSUBS 0.007451f
C998 B.n824 VSUBS 0.007451f
C999 B.n825 VSUBS 0.007451f
C1000 B.n826 VSUBS 0.007451f
C1001 B.n827 VSUBS 0.007451f
C1002 B.n828 VSUBS 0.007451f
C1003 B.n829 VSUBS 0.007451f
C1004 B.n830 VSUBS 0.007451f
C1005 B.n831 VSUBS 0.007451f
C1006 B.n832 VSUBS 0.007451f
C1007 B.n833 VSUBS 0.007451f
C1008 B.n834 VSUBS 0.007451f
C1009 B.n835 VSUBS 0.007451f
C1010 B.n836 VSUBS 0.007451f
C1011 B.n837 VSUBS 0.007451f
C1012 B.n838 VSUBS 0.007451f
C1013 B.n839 VSUBS 0.007451f
C1014 B.n840 VSUBS 0.007451f
C1015 B.n841 VSUBS 0.007451f
C1016 B.n842 VSUBS 0.018921f
C1017 B.n843 VSUBS 0.018921f
C1018 B.n844 VSUBS 0.018117f
C1019 B.n845 VSUBS 0.007451f
C1020 B.n846 VSUBS 0.007451f
C1021 B.n847 VSUBS 0.007451f
C1022 B.n848 VSUBS 0.007451f
C1023 B.n849 VSUBS 0.007451f
C1024 B.n850 VSUBS 0.007451f
C1025 B.n851 VSUBS 0.007451f
C1026 B.n852 VSUBS 0.007451f
C1027 B.n853 VSUBS 0.007451f
C1028 B.n854 VSUBS 0.007451f
C1029 B.n855 VSUBS 0.007451f
C1030 B.n856 VSUBS 0.007451f
C1031 B.n857 VSUBS 0.007451f
C1032 B.n858 VSUBS 0.007451f
C1033 B.n859 VSUBS 0.007451f
C1034 B.n860 VSUBS 0.007451f
C1035 B.n861 VSUBS 0.007451f
C1036 B.n862 VSUBS 0.007451f
C1037 B.n863 VSUBS 0.007451f
C1038 B.n864 VSUBS 0.007451f
C1039 B.n865 VSUBS 0.007451f
C1040 B.n866 VSUBS 0.007451f
C1041 B.n867 VSUBS 0.007451f
C1042 B.n868 VSUBS 0.007451f
C1043 B.n869 VSUBS 0.007451f
C1044 B.n870 VSUBS 0.007451f
C1045 B.n871 VSUBS 0.007451f
C1046 B.n872 VSUBS 0.007451f
C1047 B.n873 VSUBS 0.007451f
C1048 B.n874 VSUBS 0.007451f
C1049 B.n875 VSUBS 0.007451f
C1050 B.n876 VSUBS 0.007451f
C1051 B.n877 VSUBS 0.007451f
C1052 B.n878 VSUBS 0.007451f
C1053 B.n879 VSUBS 0.007451f
C1054 B.n880 VSUBS 0.007451f
C1055 B.n881 VSUBS 0.007451f
C1056 B.n882 VSUBS 0.007451f
C1057 B.n883 VSUBS 0.007451f
C1058 B.n884 VSUBS 0.007451f
C1059 B.n885 VSUBS 0.007451f
C1060 B.n886 VSUBS 0.007451f
C1061 B.n887 VSUBS 0.007451f
C1062 B.n888 VSUBS 0.007451f
C1063 B.n889 VSUBS 0.007451f
C1064 B.n890 VSUBS 0.007451f
C1065 B.n891 VSUBS 0.007451f
C1066 B.n892 VSUBS 0.007451f
C1067 B.n893 VSUBS 0.007451f
C1068 B.n894 VSUBS 0.007451f
C1069 B.n895 VSUBS 0.007451f
C1070 B.n896 VSUBS 0.007451f
C1071 B.n897 VSUBS 0.007451f
C1072 B.n898 VSUBS 0.007451f
C1073 B.n899 VSUBS 0.007451f
C1074 B.n900 VSUBS 0.007451f
C1075 B.n901 VSUBS 0.007451f
C1076 B.n902 VSUBS 0.007451f
C1077 B.n903 VSUBS 0.007451f
C1078 B.n904 VSUBS 0.007451f
C1079 B.n905 VSUBS 0.007451f
C1080 B.n906 VSUBS 0.007451f
C1081 B.n907 VSUBS 0.007451f
C1082 B.n908 VSUBS 0.007451f
C1083 B.n909 VSUBS 0.007451f
C1084 B.n910 VSUBS 0.007451f
C1085 B.n911 VSUBS 0.007451f
C1086 B.n912 VSUBS 0.007451f
C1087 B.n913 VSUBS 0.007451f
C1088 B.n914 VSUBS 0.007451f
C1089 B.n915 VSUBS 0.016872f
.ends

