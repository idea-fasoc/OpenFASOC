* NGSPICE file created from diff_pair_sample_1495.ext - technology: sky130A

.subckt diff_pair_sample_1495 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=2.4222 ps=15.01 w=14.68 l=0.8
X1 VTAIL.t1 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=2.4222 ps=15.01 w=14.68 l=0.8
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=0 ps=0 w=14.68 l=0.8
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=0 ps=0 w=14.68 l=0.8
X4 VDD1.t4 VP.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=2.4222 ps=15.01 w=14.68 l=0.8
X5 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=5.7252 ps=30.14 w=14.68 l=0.8
X6 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=2.4222 ps=15.01 w=14.68 l=0.8
X7 VDD1.t1 VP.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=5.7252 ps=30.14 w=14.68 l=0.8
X8 VTAIL.t4 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=2.4222 ps=15.01 w=14.68 l=0.8
X9 VDD2.t1 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=5.7252 ps=30.14 w=14.68 l=0.8
X10 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=2.4222 ps=15.01 w=14.68 l=0.8
X11 VDD1.t3 VP.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=5.7252 ps=30.14 w=14.68 l=0.8
X12 VTAIL.t7 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4222 pd=15.01 as=2.4222 ps=15.01 w=14.68 l=0.8
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=0 ps=0 w=14.68 l=0.8
X14 VDD1.t0 VP.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=2.4222 ps=15.01 w=14.68 l=0.8
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7252 pd=30.14 as=0 ps=0 w=14.68 l=0.8
R0 VP.n3 VP.t5 514.826
R1 VP.n8 VP.t1 491.339
R2 VP.n12 VP.t0 491.339
R3 VP.n14 VP.t2 491.339
R4 VP.n6 VP.t3 491.339
R5 VP.n4 VP.t4 491.339
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.8973
R14 VP.n9 VP.n7 43.724
R15 VP.n8 VP.n1 33.5944
R16 VP.n14 VP.n13 33.5944
R17 VP.n6 VP.n5 33.5944
R18 VP.n4 VP.n3 18.1882
R19 VP.n12 VP.n1 14.6066
R20 VP.n13 VP.n12 14.6066
R21 VP.n5 VP.n4 14.6066
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VDD1.n76 VDD1.n0 289.615
R29 VDD1.n157 VDD1.n81 289.615
R30 VDD1.n77 VDD1.n76 185
R31 VDD1.n75 VDD1.n74 185
R32 VDD1.n73 VDD1.n3 185
R33 VDD1.n7 VDD1.n4 185
R34 VDD1.n68 VDD1.n67 185
R35 VDD1.n66 VDD1.n65 185
R36 VDD1.n9 VDD1.n8 185
R37 VDD1.n60 VDD1.n59 185
R38 VDD1.n58 VDD1.n57 185
R39 VDD1.n13 VDD1.n12 185
R40 VDD1.n52 VDD1.n51 185
R41 VDD1.n50 VDD1.n49 185
R42 VDD1.n17 VDD1.n16 185
R43 VDD1.n44 VDD1.n43 185
R44 VDD1.n42 VDD1.n41 185
R45 VDD1.n21 VDD1.n20 185
R46 VDD1.n36 VDD1.n35 185
R47 VDD1.n34 VDD1.n33 185
R48 VDD1.n25 VDD1.n24 185
R49 VDD1.n28 VDD1.n27 185
R50 VDD1.n108 VDD1.n107 185
R51 VDD1.n105 VDD1.n104 185
R52 VDD1.n114 VDD1.n113 185
R53 VDD1.n116 VDD1.n115 185
R54 VDD1.n101 VDD1.n100 185
R55 VDD1.n122 VDD1.n121 185
R56 VDD1.n124 VDD1.n123 185
R57 VDD1.n97 VDD1.n96 185
R58 VDD1.n130 VDD1.n129 185
R59 VDD1.n132 VDD1.n131 185
R60 VDD1.n93 VDD1.n92 185
R61 VDD1.n138 VDD1.n137 185
R62 VDD1.n140 VDD1.n139 185
R63 VDD1.n89 VDD1.n88 185
R64 VDD1.n146 VDD1.n145 185
R65 VDD1.n149 VDD1.n148 185
R66 VDD1.n147 VDD1.n85 185
R67 VDD1.n154 VDD1.n84 185
R68 VDD1.n156 VDD1.n155 185
R69 VDD1.n158 VDD1.n157 185
R70 VDD1.t0 VDD1.n26 147.659
R71 VDD1.t4 VDD1.n106 147.659
R72 VDD1.n76 VDD1.n75 104.615
R73 VDD1.n75 VDD1.n3 104.615
R74 VDD1.n7 VDD1.n3 104.615
R75 VDD1.n67 VDD1.n7 104.615
R76 VDD1.n67 VDD1.n66 104.615
R77 VDD1.n66 VDD1.n8 104.615
R78 VDD1.n59 VDD1.n8 104.615
R79 VDD1.n59 VDD1.n58 104.615
R80 VDD1.n58 VDD1.n12 104.615
R81 VDD1.n51 VDD1.n12 104.615
R82 VDD1.n51 VDD1.n50 104.615
R83 VDD1.n50 VDD1.n16 104.615
R84 VDD1.n43 VDD1.n16 104.615
R85 VDD1.n43 VDD1.n42 104.615
R86 VDD1.n42 VDD1.n20 104.615
R87 VDD1.n35 VDD1.n20 104.615
R88 VDD1.n35 VDD1.n34 104.615
R89 VDD1.n34 VDD1.n24 104.615
R90 VDD1.n27 VDD1.n24 104.615
R91 VDD1.n107 VDD1.n104 104.615
R92 VDD1.n114 VDD1.n104 104.615
R93 VDD1.n115 VDD1.n114 104.615
R94 VDD1.n115 VDD1.n100 104.615
R95 VDD1.n122 VDD1.n100 104.615
R96 VDD1.n123 VDD1.n122 104.615
R97 VDD1.n123 VDD1.n96 104.615
R98 VDD1.n130 VDD1.n96 104.615
R99 VDD1.n131 VDD1.n130 104.615
R100 VDD1.n131 VDD1.n92 104.615
R101 VDD1.n138 VDD1.n92 104.615
R102 VDD1.n139 VDD1.n138 104.615
R103 VDD1.n139 VDD1.n88 104.615
R104 VDD1.n146 VDD1.n88 104.615
R105 VDD1.n148 VDD1.n146 104.615
R106 VDD1.n148 VDD1.n147 104.615
R107 VDD1.n147 VDD1.n84 104.615
R108 VDD1.n156 VDD1.n84 104.615
R109 VDD1.n157 VDD1.n156 104.615
R110 VDD1.n163 VDD1.n162 61.8849
R111 VDD1.n165 VDD1.n164 61.6967
R112 VDD1.n27 VDD1.t0 52.3082
R113 VDD1.n107 VDD1.t4 52.3082
R114 VDD1 VDD1.n80 50.4287
R115 VDD1.n163 VDD1.n161 50.3152
R116 VDD1.n165 VDD1.n163 40.6065
R117 VDD1.n28 VDD1.n26 15.6677
R118 VDD1.n108 VDD1.n106 15.6677
R119 VDD1.n74 VDD1.n73 13.1884
R120 VDD1.n155 VDD1.n154 13.1884
R121 VDD1.n77 VDD1.n2 12.8005
R122 VDD1.n72 VDD1.n4 12.8005
R123 VDD1.n29 VDD1.n25 12.8005
R124 VDD1.n109 VDD1.n105 12.8005
R125 VDD1.n153 VDD1.n85 12.8005
R126 VDD1.n158 VDD1.n83 12.8005
R127 VDD1.n78 VDD1.n0 12.0247
R128 VDD1.n69 VDD1.n68 12.0247
R129 VDD1.n33 VDD1.n32 12.0247
R130 VDD1.n113 VDD1.n112 12.0247
R131 VDD1.n150 VDD1.n149 12.0247
R132 VDD1.n159 VDD1.n81 12.0247
R133 VDD1.n65 VDD1.n6 11.249
R134 VDD1.n36 VDD1.n23 11.249
R135 VDD1.n116 VDD1.n103 11.249
R136 VDD1.n145 VDD1.n87 11.249
R137 VDD1.n64 VDD1.n9 10.4732
R138 VDD1.n37 VDD1.n21 10.4732
R139 VDD1.n117 VDD1.n101 10.4732
R140 VDD1.n144 VDD1.n89 10.4732
R141 VDD1.n61 VDD1.n60 9.69747
R142 VDD1.n41 VDD1.n40 9.69747
R143 VDD1.n121 VDD1.n120 9.69747
R144 VDD1.n141 VDD1.n140 9.69747
R145 VDD1.n80 VDD1.n79 9.45567
R146 VDD1.n161 VDD1.n160 9.45567
R147 VDD1.n54 VDD1.n53 9.3005
R148 VDD1.n56 VDD1.n55 9.3005
R149 VDD1.n11 VDD1.n10 9.3005
R150 VDD1.n62 VDD1.n61 9.3005
R151 VDD1.n64 VDD1.n63 9.3005
R152 VDD1.n6 VDD1.n5 9.3005
R153 VDD1.n70 VDD1.n69 9.3005
R154 VDD1.n72 VDD1.n71 9.3005
R155 VDD1.n79 VDD1.n78 9.3005
R156 VDD1.n2 VDD1.n1 9.3005
R157 VDD1.n15 VDD1.n14 9.3005
R158 VDD1.n48 VDD1.n47 9.3005
R159 VDD1.n46 VDD1.n45 9.3005
R160 VDD1.n19 VDD1.n18 9.3005
R161 VDD1.n40 VDD1.n39 9.3005
R162 VDD1.n38 VDD1.n37 9.3005
R163 VDD1.n23 VDD1.n22 9.3005
R164 VDD1.n32 VDD1.n31 9.3005
R165 VDD1.n30 VDD1.n29 9.3005
R166 VDD1.n160 VDD1.n159 9.3005
R167 VDD1.n83 VDD1.n82 9.3005
R168 VDD1.n128 VDD1.n127 9.3005
R169 VDD1.n126 VDD1.n125 9.3005
R170 VDD1.n99 VDD1.n98 9.3005
R171 VDD1.n120 VDD1.n119 9.3005
R172 VDD1.n118 VDD1.n117 9.3005
R173 VDD1.n103 VDD1.n102 9.3005
R174 VDD1.n112 VDD1.n111 9.3005
R175 VDD1.n110 VDD1.n109 9.3005
R176 VDD1.n95 VDD1.n94 9.3005
R177 VDD1.n134 VDD1.n133 9.3005
R178 VDD1.n136 VDD1.n135 9.3005
R179 VDD1.n91 VDD1.n90 9.3005
R180 VDD1.n142 VDD1.n141 9.3005
R181 VDD1.n144 VDD1.n143 9.3005
R182 VDD1.n87 VDD1.n86 9.3005
R183 VDD1.n151 VDD1.n150 9.3005
R184 VDD1.n153 VDD1.n152 9.3005
R185 VDD1.n57 VDD1.n11 8.92171
R186 VDD1.n44 VDD1.n19 8.92171
R187 VDD1.n124 VDD1.n99 8.92171
R188 VDD1.n137 VDD1.n91 8.92171
R189 VDD1.n56 VDD1.n13 8.14595
R190 VDD1.n45 VDD1.n17 8.14595
R191 VDD1.n125 VDD1.n97 8.14595
R192 VDD1.n136 VDD1.n93 8.14595
R193 VDD1.n53 VDD1.n52 7.3702
R194 VDD1.n49 VDD1.n48 7.3702
R195 VDD1.n129 VDD1.n128 7.3702
R196 VDD1.n133 VDD1.n132 7.3702
R197 VDD1.n52 VDD1.n15 6.59444
R198 VDD1.n49 VDD1.n15 6.59444
R199 VDD1.n129 VDD1.n95 6.59444
R200 VDD1.n132 VDD1.n95 6.59444
R201 VDD1.n53 VDD1.n13 5.81868
R202 VDD1.n48 VDD1.n17 5.81868
R203 VDD1.n128 VDD1.n97 5.81868
R204 VDD1.n133 VDD1.n93 5.81868
R205 VDD1.n57 VDD1.n56 5.04292
R206 VDD1.n45 VDD1.n44 5.04292
R207 VDD1.n125 VDD1.n124 5.04292
R208 VDD1.n137 VDD1.n136 5.04292
R209 VDD1.n30 VDD1.n26 4.38563
R210 VDD1.n110 VDD1.n106 4.38563
R211 VDD1.n60 VDD1.n11 4.26717
R212 VDD1.n41 VDD1.n19 4.26717
R213 VDD1.n121 VDD1.n99 4.26717
R214 VDD1.n140 VDD1.n91 4.26717
R215 VDD1.n61 VDD1.n9 3.49141
R216 VDD1.n40 VDD1.n21 3.49141
R217 VDD1.n120 VDD1.n101 3.49141
R218 VDD1.n141 VDD1.n89 3.49141
R219 VDD1.n65 VDD1.n64 2.71565
R220 VDD1.n37 VDD1.n36 2.71565
R221 VDD1.n117 VDD1.n116 2.71565
R222 VDD1.n145 VDD1.n144 2.71565
R223 VDD1.n80 VDD1.n0 1.93989
R224 VDD1.n68 VDD1.n6 1.93989
R225 VDD1.n33 VDD1.n23 1.93989
R226 VDD1.n113 VDD1.n103 1.93989
R227 VDD1.n149 VDD1.n87 1.93989
R228 VDD1.n161 VDD1.n81 1.93989
R229 VDD1.n164 VDD1.t5 1.34927
R230 VDD1.n164 VDD1.t3 1.34927
R231 VDD1.n162 VDD1.t2 1.34927
R232 VDD1.n162 VDD1.t1 1.34927
R233 VDD1.n78 VDD1.n77 1.16414
R234 VDD1.n69 VDD1.n4 1.16414
R235 VDD1.n32 VDD1.n25 1.16414
R236 VDD1.n112 VDD1.n105 1.16414
R237 VDD1.n150 VDD1.n85 1.16414
R238 VDD1.n159 VDD1.n158 1.16414
R239 VDD1.n74 VDD1.n2 0.388379
R240 VDD1.n73 VDD1.n72 0.388379
R241 VDD1.n29 VDD1.n28 0.388379
R242 VDD1.n109 VDD1.n108 0.388379
R243 VDD1.n154 VDD1.n153 0.388379
R244 VDD1.n155 VDD1.n83 0.388379
R245 VDD1 VDD1.n165 0.185845
R246 VDD1.n79 VDD1.n1 0.155672
R247 VDD1.n71 VDD1.n1 0.155672
R248 VDD1.n71 VDD1.n70 0.155672
R249 VDD1.n70 VDD1.n5 0.155672
R250 VDD1.n63 VDD1.n5 0.155672
R251 VDD1.n63 VDD1.n62 0.155672
R252 VDD1.n62 VDD1.n10 0.155672
R253 VDD1.n55 VDD1.n10 0.155672
R254 VDD1.n55 VDD1.n54 0.155672
R255 VDD1.n54 VDD1.n14 0.155672
R256 VDD1.n47 VDD1.n14 0.155672
R257 VDD1.n47 VDD1.n46 0.155672
R258 VDD1.n46 VDD1.n18 0.155672
R259 VDD1.n39 VDD1.n18 0.155672
R260 VDD1.n39 VDD1.n38 0.155672
R261 VDD1.n38 VDD1.n22 0.155672
R262 VDD1.n31 VDD1.n22 0.155672
R263 VDD1.n31 VDD1.n30 0.155672
R264 VDD1.n111 VDD1.n110 0.155672
R265 VDD1.n111 VDD1.n102 0.155672
R266 VDD1.n118 VDD1.n102 0.155672
R267 VDD1.n119 VDD1.n118 0.155672
R268 VDD1.n119 VDD1.n98 0.155672
R269 VDD1.n126 VDD1.n98 0.155672
R270 VDD1.n127 VDD1.n126 0.155672
R271 VDD1.n127 VDD1.n94 0.155672
R272 VDD1.n134 VDD1.n94 0.155672
R273 VDD1.n135 VDD1.n134 0.155672
R274 VDD1.n135 VDD1.n90 0.155672
R275 VDD1.n142 VDD1.n90 0.155672
R276 VDD1.n143 VDD1.n142 0.155672
R277 VDD1.n143 VDD1.n86 0.155672
R278 VDD1.n151 VDD1.n86 0.155672
R279 VDD1.n152 VDD1.n151 0.155672
R280 VDD1.n152 VDD1.n82 0.155672
R281 VDD1.n160 VDD1.n82 0.155672
R282 VTAIL.n330 VTAIL.n254 289.615
R283 VTAIL.n78 VTAIL.n2 289.615
R284 VTAIL.n248 VTAIL.n172 289.615
R285 VTAIL.n164 VTAIL.n88 289.615
R286 VTAIL.n281 VTAIL.n280 185
R287 VTAIL.n278 VTAIL.n277 185
R288 VTAIL.n287 VTAIL.n286 185
R289 VTAIL.n289 VTAIL.n288 185
R290 VTAIL.n274 VTAIL.n273 185
R291 VTAIL.n295 VTAIL.n294 185
R292 VTAIL.n297 VTAIL.n296 185
R293 VTAIL.n270 VTAIL.n269 185
R294 VTAIL.n303 VTAIL.n302 185
R295 VTAIL.n305 VTAIL.n304 185
R296 VTAIL.n266 VTAIL.n265 185
R297 VTAIL.n311 VTAIL.n310 185
R298 VTAIL.n313 VTAIL.n312 185
R299 VTAIL.n262 VTAIL.n261 185
R300 VTAIL.n319 VTAIL.n318 185
R301 VTAIL.n322 VTAIL.n321 185
R302 VTAIL.n320 VTAIL.n258 185
R303 VTAIL.n327 VTAIL.n257 185
R304 VTAIL.n329 VTAIL.n328 185
R305 VTAIL.n331 VTAIL.n330 185
R306 VTAIL.n29 VTAIL.n28 185
R307 VTAIL.n26 VTAIL.n25 185
R308 VTAIL.n35 VTAIL.n34 185
R309 VTAIL.n37 VTAIL.n36 185
R310 VTAIL.n22 VTAIL.n21 185
R311 VTAIL.n43 VTAIL.n42 185
R312 VTAIL.n45 VTAIL.n44 185
R313 VTAIL.n18 VTAIL.n17 185
R314 VTAIL.n51 VTAIL.n50 185
R315 VTAIL.n53 VTAIL.n52 185
R316 VTAIL.n14 VTAIL.n13 185
R317 VTAIL.n59 VTAIL.n58 185
R318 VTAIL.n61 VTAIL.n60 185
R319 VTAIL.n10 VTAIL.n9 185
R320 VTAIL.n67 VTAIL.n66 185
R321 VTAIL.n70 VTAIL.n69 185
R322 VTAIL.n68 VTAIL.n6 185
R323 VTAIL.n75 VTAIL.n5 185
R324 VTAIL.n77 VTAIL.n76 185
R325 VTAIL.n79 VTAIL.n78 185
R326 VTAIL.n249 VTAIL.n248 185
R327 VTAIL.n247 VTAIL.n246 185
R328 VTAIL.n245 VTAIL.n175 185
R329 VTAIL.n179 VTAIL.n176 185
R330 VTAIL.n240 VTAIL.n239 185
R331 VTAIL.n238 VTAIL.n237 185
R332 VTAIL.n181 VTAIL.n180 185
R333 VTAIL.n232 VTAIL.n231 185
R334 VTAIL.n230 VTAIL.n229 185
R335 VTAIL.n185 VTAIL.n184 185
R336 VTAIL.n224 VTAIL.n223 185
R337 VTAIL.n222 VTAIL.n221 185
R338 VTAIL.n189 VTAIL.n188 185
R339 VTAIL.n216 VTAIL.n215 185
R340 VTAIL.n214 VTAIL.n213 185
R341 VTAIL.n193 VTAIL.n192 185
R342 VTAIL.n208 VTAIL.n207 185
R343 VTAIL.n206 VTAIL.n205 185
R344 VTAIL.n197 VTAIL.n196 185
R345 VTAIL.n200 VTAIL.n199 185
R346 VTAIL.n165 VTAIL.n164 185
R347 VTAIL.n163 VTAIL.n162 185
R348 VTAIL.n161 VTAIL.n91 185
R349 VTAIL.n95 VTAIL.n92 185
R350 VTAIL.n156 VTAIL.n155 185
R351 VTAIL.n154 VTAIL.n153 185
R352 VTAIL.n97 VTAIL.n96 185
R353 VTAIL.n148 VTAIL.n147 185
R354 VTAIL.n146 VTAIL.n145 185
R355 VTAIL.n101 VTAIL.n100 185
R356 VTAIL.n140 VTAIL.n139 185
R357 VTAIL.n138 VTAIL.n137 185
R358 VTAIL.n105 VTAIL.n104 185
R359 VTAIL.n132 VTAIL.n131 185
R360 VTAIL.n130 VTAIL.n129 185
R361 VTAIL.n109 VTAIL.n108 185
R362 VTAIL.n124 VTAIL.n123 185
R363 VTAIL.n122 VTAIL.n121 185
R364 VTAIL.n113 VTAIL.n112 185
R365 VTAIL.n116 VTAIL.n115 185
R366 VTAIL.t8 VTAIL.n198 147.659
R367 VTAIL.t2 VTAIL.n114 147.659
R368 VTAIL.t3 VTAIL.n279 147.659
R369 VTAIL.t9 VTAIL.n27 147.659
R370 VTAIL.n280 VTAIL.n277 104.615
R371 VTAIL.n287 VTAIL.n277 104.615
R372 VTAIL.n288 VTAIL.n287 104.615
R373 VTAIL.n288 VTAIL.n273 104.615
R374 VTAIL.n295 VTAIL.n273 104.615
R375 VTAIL.n296 VTAIL.n295 104.615
R376 VTAIL.n296 VTAIL.n269 104.615
R377 VTAIL.n303 VTAIL.n269 104.615
R378 VTAIL.n304 VTAIL.n303 104.615
R379 VTAIL.n304 VTAIL.n265 104.615
R380 VTAIL.n311 VTAIL.n265 104.615
R381 VTAIL.n312 VTAIL.n311 104.615
R382 VTAIL.n312 VTAIL.n261 104.615
R383 VTAIL.n319 VTAIL.n261 104.615
R384 VTAIL.n321 VTAIL.n319 104.615
R385 VTAIL.n321 VTAIL.n320 104.615
R386 VTAIL.n320 VTAIL.n257 104.615
R387 VTAIL.n329 VTAIL.n257 104.615
R388 VTAIL.n330 VTAIL.n329 104.615
R389 VTAIL.n28 VTAIL.n25 104.615
R390 VTAIL.n35 VTAIL.n25 104.615
R391 VTAIL.n36 VTAIL.n35 104.615
R392 VTAIL.n36 VTAIL.n21 104.615
R393 VTAIL.n43 VTAIL.n21 104.615
R394 VTAIL.n44 VTAIL.n43 104.615
R395 VTAIL.n44 VTAIL.n17 104.615
R396 VTAIL.n51 VTAIL.n17 104.615
R397 VTAIL.n52 VTAIL.n51 104.615
R398 VTAIL.n52 VTAIL.n13 104.615
R399 VTAIL.n59 VTAIL.n13 104.615
R400 VTAIL.n60 VTAIL.n59 104.615
R401 VTAIL.n60 VTAIL.n9 104.615
R402 VTAIL.n67 VTAIL.n9 104.615
R403 VTAIL.n69 VTAIL.n67 104.615
R404 VTAIL.n69 VTAIL.n68 104.615
R405 VTAIL.n68 VTAIL.n5 104.615
R406 VTAIL.n77 VTAIL.n5 104.615
R407 VTAIL.n78 VTAIL.n77 104.615
R408 VTAIL.n248 VTAIL.n247 104.615
R409 VTAIL.n247 VTAIL.n175 104.615
R410 VTAIL.n179 VTAIL.n175 104.615
R411 VTAIL.n239 VTAIL.n179 104.615
R412 VTAIL.n239 VTAIL.n238 104.615
R413 VTAIL.n238 VTAIL.n180 104.615
R414 VTAIL.n231 VTAIL.n180 104.615
R415 VTAIL.n231 VTAIL.n230 104.615
R416 VTAIL.n230 VTAIL.n184 104.615
R417 VTAIL.n223 VTAIL.n184 104.615
R418 VTAIL.n223 VTAIL.n222 104.615
R419 VTAIL.n222 VTAIL.n188 104.615
R420 VTAIL.n215 VTAIL.n188 104.615
R421 VTAIL.n215 VTAIL.n214 104.615
R422 VTAIL.n214 VTAIL.n192 104.615
R423 VTAIL.n207 VTAIL.n192 104.615
R424 VTAIL.n207 VTAIL.n206 104.615
R425 VTAIL.n206 VTAIL.n196 104.615
R426 VTAIL.n199 VTAIL.n196 104.615
R427 VTAIL.n164 VTAIL.n163 104.615
R428 VTAIL.n163 VTAIL.n91 104.615
R429 VTAIL.n95 VTAIL.n91 104.615
R430 VTAIL.n155 VTAIL.n95 104.615
R431 VTAIL.n155 VTAIL.n154 104.615
R432 VTAIL.n154 VTAIL.n96 104.615
R433 VTAIL.n147 VTAIL.n96 104.615
R434 VTAIL.n147 VTAIL.n146 104.615
R435 VTAIL.n146 VTAIL.n100 104.615
R436 VTAIL.n139 VTAIL.n100 104.615
R437 VTAIL.n139 VTAIL.n138 104.615
R438 VTAIL.n138 VTAIL.n104 104.615
R439 VTAIL.n131 VTAIL.n104 104.615
R440 VTAIL.n131 VTAIL.n130 104.615
R441 VTAIL.n130 VTAIL.n108 104.615
R442 VTAIL.n123 VTAIL.n108 104.615
R443 VTAIL.n123 VTAIL.n122 104.615
R444 VTAIL.n122 VTAIL.n112 104.615
R445 VTAIL.n115 VTAIL.n112 104.615
R446 VTAIL.n280 VTAIL.t3 52.3082
R447 VTAIL.n28 VTAIL.t9 52.3082
R448 VTAIL.n199 VTAIL.t8 52.3082
R449 VTAIL.n115 VTAIL.t2 52.3082
R450 VTAIL.n171 VTAIL.n170 45.0181
R451 VTAIL.n87 VTAIL.n86 45.0181
R452 VTAIL.n1 VTAIL.n0 45.0179
R453 VTAIL.n85 VTAIL.n84 45.0179
R454 VTAIL.n335 VTAIL.n334 32.9611
R455 VTAIL.n83 VTAIL.n82 32.9611
R456 VTAIL.n253 VTAIL.n252 32.9611
R457 VTAIL.n169 VTAIL.n168 32.9611
R458 VTAIL.n87 VTAIL.n85 26.9703
R459 VTAIL.n335 VTAIL.n253 25.9962
R460 VTAIL.n281 VTAIL.n279 15.6677
R461 VTAIL.n29 VTAIL.n27 15.6677
R462 VTAIL.n200 VTAIL.n198 15.6677
R463 VTAIL.n116 VTAIL.n114 15.6677
R464 VTAIL.n328 VTAIL.n327 13.1884
R465 VTAIL.n76 VTAIL.n75 13.1884
R466 VTAIL.n246 VTAIL.n245 13.1884
R467 VTAIL.n162 VTAIL.n161 13.1884
R468 VTAIL.n282 VTAIL.n278 12.8005
R469 VTAIL.n326 VTAIL.n258 12.8005
R470 VTAIL.n331 VTAIL.n256 12.8005
R471 VTAIL.n30 VTAIL.n26 12.8005
R472 VTAIL.n74 VTAIL.n6 12.8005
R473 VTAIL.n79 VTAIL.n4 12.8005
R474 VTAIL.n249 VTAIL.n174 12.8005
R475 VTAIL.n244 VTAIL.n176 12.8005
R476 VTAIL.n201 VTAIL.n197 12.8005
R477 VTAIL.n165 VTAIL.n90 12.8005
R478 VTAIL.n160 VTAIL.n92 12.8005
R479 VTAIL.n117 VTAIL.n113 12.8005
R480 VTAIL.n286 VTAIL.n285 12.0247
R481 VTAIL.n323 VTAIL.n322 12.0247
R482 VTAIL.n332 VTAIL.n254 12.0247
R483 VTAIL.n34 VTAIL.n33 12.0247
R484 VTAIL.n71 VTAIL.n70 12.0247
R485 VTAIL.n80 VTAIL.n2 12.0247
R486 VTAIL.n250 VTAIL.n172 12.0247
R487 VTAIL.n241 VTAIL.n240 12.0247
R488 VTAIL.n205 VTAIL.n204 12.0247
R489 VTAIL.n166 VTAIL.n88 12.0247
R490 VTAIL.n157 VTAIL.n156 12.0247
R491 VTAIL.n121 VTAIL.n120 12.0247
R492 VTAIL.n289 VTAIL.n276 11.249
R493 VTAIL.n318 VTAIL.n260 11.249
R494 VTAIL.n37 VTAIL.n24 11.249
R495 VTAIL.n66 VTAIL.n8 11.249
R496 VTAIL.n237 VTAIL.n178 11.249
R497 VTAIL.n208 VTAIL.n195 11.249
R498 VTAIL.n153 VTAIL.n94 11.249
R499 VTAIL.n124 VTAIL.n111 11.249
R500 VTAIL.n290 VTAIL.n274 10.4732
R501 VTAIL.n317 VTAIL.n262 10.4732
R502 VTAIL.n38 VTAIL.n22 10.4732
R503 VTAIL.n65 VTAIL.n10 10.4732
R504 VTAIL.n236 VTAIL.n181 10.4732
R505 VTAIL.n209 VTAIL.n193 10.4732
R506 VTAIL.n152 VTAIL.n97 10.4732
R507 VTAIL.n125 VTAIL.n109 10.4732
R508 VTAIL.n294 VTAIL.n293 9.69747
R509 VTAIL.n314 VTAIL.n313 9.69747
R510 VTAIL.n42 VTAIL.n41 9.69747
R511 VTAIL.n62 VTAIL.n61 9.69747
R512 VTAIL.n233 VTAIL.n232 9.69747
R513 VTAIL.n213 VTAIL.n212 9.69747
R514 VTAIL.n149 VTAIL.n148 9.69747
R515 VTAIL.n129 VTAIL.n128 9.69747
R516 VTAIL.n334 VTAIL.n333 9.45567
R517 VTAIL.n82 VTAIL.n81 9.45567
R518 VTAIL.n252 VTAIL.n251 9.45567
R519 VTAIL.n168 VTAIL.n167 9.45567
R520 VTAIL.n333 VTAIL.n332 9.3005
R521 VTAIL.n256 VTAIL.n255 9.3005
R522 VTAIL.n301 VTAIL.n300 9.3005
R523 VTAIL.n299 VTAIL.n298 9.3005
R524 VTAIL.n272 VTAIL.n271 9.3005
R525 VTAIL.n293 VTAIL.n292 9.3005
R526 VTAIL.n291 VTAIL.n290 9.3005
R527 VTAIL.n276 VTAIL.n275 9.3005
R528 VTAIL.n285 VTAIL.n284 9.3005
R529 VTAIL.n283 VTAIL.n282 9.3005
R530 VTAIL.n268 VTAIL.n267 9.3005
R531 VTAIL.n307 VTAIL.n306 9.3005
R532 VTAIL.n309 VTAIL.n308 9.3005
R533 VTAIL.n264 VTAIL.n263 9.3005
R534 VTAIL.n315 VTAIL.n314 9.3005
R535 VTAIL.n317 VTAIL.n316 9.3005
R536 VTAIL.n260 VTAIL.n259 9.3005
R537 VTAIL.n324 VTAIL.n323 9.3005
R538 VTAIL.n326 VTAIL.n325 9.3005
R539 VTAIL.n81 VTAIL.n80 9.3005
R540 VTAIL.n4 VTAIL.n3 9.3005
R541 VTAIL.n49 VTAIL.n48 9.3005
R542 VTAIL.n47 VTAIL.n46 9.3005
R543 VTAIL.n20 VTAIL.n19 9.3005
R544 VTAIL.n41 VTAIL.n40 9.3005
R545 VTAIL.n39 VTAIL.n38 9.3005
R546 VTAIL.n24 VTAIL.n23 9.3005
R547 VTAIL.n33 VTAIL.n32 9.3005
R548 VTAIL.n31 VTAIL.n30 9.3005
R549 VTAIL.n16 VTAIL.n15 9.3005
R550 VTAIL.n55 VTAIL.n54 9.3005
R551 VTAIL.n57 VTAIL.n56 9.3005
R552 VTAIL.n12 VTAIL.n11 9.3005
R553 VTAIL.n63 VTAIL.n62 9.3005
R554 VTAIL.n65 VTAIL.n64 9.3005
R555 VTAIL.n8 VTAIL.n7 9.3005
R556 VTAIL.n72 VTAIL.n71 9.3005
R557 VTAIL.n74 VTAIL.n73 9.3005
R558 VTAIL.n226 VTAIL.n225 9.3005
R559 VTAIL.n228 VTAIL.n227 9.3005
R560 VTAIL.n183 VTAIL.n182 9.3005
R561 VTAIL.n234 VTAIL.n233 9.3005
R562 VTAIL.n236 VTAIL.n235 9.3005
R563 VTAIL.n178 VTAIL.n177 9.3005
R564 VTAIL.n242 VTAIL.n241 9.3005
R565 VTAIL.n244 VTAIL.n243 9.3005
R566 VTAIL.n251 VTAIL.n250 9.3005
R567 VTAIL.n174 VTAIL.n173 9.3005
R568 VTAIL.n187 VTAIL.n186 9.3005
R569 VTAIL.n220 VTAIL.n219 9.3005
R570 VTAIL.n218 VTAIL.n217 9.3005
R571 VTAIL.n191 VTAIL.n190 9.3005
R572 VTAIL.n212 VTAIL.n211 9.3005
R573 VTAIL.n210 VTAIL.n209 9.3005
R574 VTAIL.n195 VTAIL.n194 9.3005
R575 VTAIL.n204 VTAIL.n203 9.3005
R576 VTAIL.n202 VTAIL.n201 9.3005
R577 VTAIL.n142 VTAIL.n141 9.3005
R578 VTAIL.n144 VTAIL.n143 9.3005
R579 VTAIL.n99 VTAIL.n98 9.3005
R580 VTAIL.n150 VTAIL.n149 9.3005
R581 VTAIL.n152 VTAIL.n151 9.3005
R582 VTAIL.n94 VTAIL.n93 9.3005
R583 VTAIL.n158 VTAIL.n157 9.3005
R584 VTAIL.n160 VTAIL.n159 9.3005
R585 VTAIL.n167 VTAIL.n166 9.3005
R586 VTAIL.n90 VTAIL.n89 9.3005
R587 VTAIL.n103 VTAIL.n102 9.3005
R588 VTAIL.n136 VTAIL.n135 9.3005
R589 VTAIL.n134 VTAIL.n133 9.3005
R590 VTAIL.n107 VTAIL.n106 9.3005
R591 VTAIL.n128 VTAIL.n127 9.3005
R592 VTAIL.n126 VTAIL.n125 9.3005
R593 VTAIL.n111 VTAIL.n110 9.3005
R594 VTAIL.n120 VTAIL.n119 9.3005
R595 VTAIL.n118 VTAIL.n117 9.3005
R596 VTAIL.n297 VTAIL.n272 8.92171
R597 VTAIL.n310 VTAIL.n264 8.92171
R598 VTAIL.n45 VTAIL.n20 8.92171
R599 VTAIL.n58 VTAIL.n12 8.92171
R600 VTAIL.n229 VTAIL.n183 8.92171
R601 VTAIL.n216 VTAIL.n191 8.92171
R602 VTAIL.n145 VTAIL.n99 8.92171
R603 VTAIL.n132 VTAIL.n107 8.92171
R604 VTAIL.n298 VTAIL.n270 8.14595
R605 VTAIL.n309 VTAIL.n266 8.14595
R606 VTAIL.n46 VTAIL.n18 8.14595
R607 VTAIL.n57 VTAIL.n14 8.14595
R608 VTAIL.n228 VTAIL.n185 8.14595
R609 VTAIL.n217 VTAIL.n189 8.14595
R610 VTAIL.n144 VTAIL.n101 8.14595
R611 VTAIL.n133 VTAIL.n105 8.14595
R612 VTAIL.n302 VTAIL.n301 7.3702
R613 VTAIL.n306 VTAIL.n305 7.3702
R614 VTAIL.n50 VTAIL.n49 7.3702
R615 VTAIL.n54 VTAIL.n53 7.3702
R616 VTAIL.n225 VTAIL.n224 7.3702
R617 VTAIL.n221 VTAIL.n220 7.3702
R618 VTAIL.n141 VTAIL.n140 7.3702
R619 VTAIL.n137 VTAIL.n136 7.3702
R620 VTAIL.n302 VTAIL.n268 6.59444
R621 VTAIL.n305 VTAIL.n268 6.59444
R622 VTAIL.n50 VTAIL.n16 6.59444
R623 VTAIL.n53 VTAIL.n16 6.59444
R624 VTAIL.n224 VTAIL.n187 6.59444
R625 VTAIL.n221 VTAIL.n187 6.59444
R626 VTAIL.n140 VTAIL.n103 6.59444
R627 VTAIL.n137 VTAIL.n103 6.59444
R628 VTAIL.n301 VTAIL.n270 5.81868
R629 VTAIL.n306 VTAIL.n266 5.81868
R630 VTAIL.n49 VTAIL.n18 5.81868
R631 VTAIL.n54 VTAIL.n14 5.81868
R632 VTAIL.n225 VTAIL.n185 5.81868
R633 VTAIL.n220 VTAIL.n189 5.81868
R634 VTAIL.n141 VTAIL.n101 5.81868
R635 VTAIL.n136 VTAIL.n105 5.81868
R636 VTAIL.n298 VTAIL.n297 5.04292
R637 VTAIL.n310 VTAIL.n309 5.04292
R638 VTAIL.n46 VTAIL.n45 5.04292
R639 VTAIL.n58 VTAIL.n57 5.04292
R640 VTAIL.n229 VTAIL.n228 5.04292
R641 VTAIL.n217 VTAIL.n216 5.04292
R642 VTAIL.n145 VTAIL.n144 5.04292
R643 VTAIL.n133 VTAIL.n132 5.04292
R644 VTAIL.n202 VTAIL.n198 4.38563
R645 VTAIL.n118 VTAIL.n114 4.38563
R646 VTAIL.n283 VTAIL.n279 4.38563
R647 VTAIL.n31 VTAIL.n27 4.38563
R648 VTAIL.n294 VTAIL.n272 4.26717
R649 VTAIL.n313 VTAIL.n264 4.26717
R650 VTAIL.n42 VTAIL.n20 4.26717
R651 VTAIL.n61 VTAIL.n12 4.26717
R652 VTAIL.n232 VTAIL.n183 4.26717
R653 VTAIL.n213 VTAIL.n191 4.26717
R654 VTAIL.n148 VTAIL.n99 4.26717
R655 VTAIL.n129 VTAIL.n107 4.26717
R656 VTAIL.n293 VTAIL.n274 3.49141
R657 VTAIL.n314 VTAIL.n262 3.49141
R658 VTAIL.n41 VTAIL.n22 3.49141
R659 VTAIL.n62 VTAIL.n10 3.49141
R660 VTAIL.n233 VTAIL.n181 3.49141
R661 VTAIL.n212 VTAIL.n193 3.49141
R662 VTAIL.n149 VTAIL.n97 3.49141
R663 VTAIL.n128 VTAIL.n109 3.49141
R664 VTAIL.n290 VTAIL.n289 2.71565
R665 VTAIL.n318 VTAIL.n317 2.71565
R666 VTAIL.n38 VTAIL.n37 2.71565
R667 VTAIL.n66 VTAIL.n65 2.71565
R668 VTAIL.n237 VTAIL.n236 2.71565
R669 VTAIL.n209 VTAIL.n208 2.71565
R670 VTAIL.n153 VTAIL.n152 2.71565
R671 VTAIL.n125 VTAIL.n124 2.71565
R672 VTAIL.n286 VTAIL.n276 1.93989
R673 VTAIL.n322 VTAIL.n260 1.93989
R674 VTAIL.n334 VTAIL.n254 1.93989
R675 VTAIL.n34 VTAIL.n24 1.93989
R676 VTAIL.n70 VTAIL.n8 1.93989
R677 VTAIL.n82 VTAIL.n2 1.93989
R678 VTAIL.n252 VTAIL.n172 1.93989
R679 VTAIL.n240 VTAIL.n178 1.93989
R680 VTAIL.n205 VTAIL.n195 1.93989
R681 VTAIL.n168 VTAIL.n88 1.93989
R682 VTAIL.n156 VTAIL.n94 1.93989
R683 VTAIL.n121 VTAIL.n111 1.93989
R684 VTAIL.n0 VTAIL.t0 1.34927
R685 VTAIL.n0 VTAIL.t1 1.34927
R686 VTAIL.n84 VTAIL.t10 1.34927
R687 VTAIL.n84 VTAIL.t11 1.34927
R688 VTAIL.n170 VTAIL.t6 1.34927
R689 VTAIL.n170 VTAIL.t7 1.34927
R690 VTAIL.n86 VTAIL.t5 1.34927
R691 VTAIL.n86 VTAIL.t4 1.34927
R692 VTAIL.n285 VTAIL.n278 1.16414
R693 VTAIL.n323 VTAIL.n258 1.16414
R694 VTAIL.n332 VTAIL.n331 1.16414
R695 VTAIL.n33 VTAIL.n26 1.16414
R696 VTAIL.n71 VTAIL.n6 1.16414
R697 VTAIL.n80 VTAIL.n79 1.16414
R698 VTAIL.n250 VTAIL.n249 1.16414
R699 VTAIL.n241 VTAIL.n176 1.16414
R700 VTAIL.n204 VTAIL.n197 1.16414
R701 VTAIL.n166 VTAIL.n165 1.16414
R702 VTAIL.n157 VTAIL.n92 1.16414
R703 VTAIL.n120 VTAIL.n113 1.16414
R704 VTAIL.n169 VTAIL.n87 0.974638
R705 VTAIL.n253 VTAIL.n171 0.974638
R706 VTAIL.n85 VTAIL.n83 0.974638
R707 VTAIL.n171 VTAIL.n169 0.957397
R708 VTAIL.n83 VTAIL.n1 0.957397
R709 VTAIL VTAIL.n335 0.672914
R710 VTAIL.n282 VTAIL.n281 0.388379
R711 VTAIL.n327 VTAIL.n326 0.388379
R712 VTAIL.n328 VTAIL.n256 0.388379
R713 VTAIL.n30 VTAIL.n29 0.388379
R714 VTAIL.n75 VTAIL.n74 0.388379
R715 VTAIL.n76 VTAIL.n4 0.388379
R716 VTAIL.n246 VTAIL.n174 0.388379
R717 VTAIL.n245 VTAIL.n244 0.388379
R718 VTAIL.n201 VTAIL.n200 0.388379
R719 VTAIL.n162 VTAIL.n90 0.388379
R720 VTAIL.n161 VTAIL.n160 0.388379
R721 VTAIL.n117 VTAIL.n116 0.388379
R722 VTAIL VTAIL.n1 0.302224
R723 VTAIL.n284 VTAIL.n283 0.155672
R724 VTAIL.n284 VTAIL.n275 0.155672
R725 VTAIL.n291 VTAIL.n275 0.155672
R726 VTAIL.n292 VTAIL.n291 0.155672
R727 VTAIL.n292 VTAIL.n271 0.155672
R728 VTAIL.n299 VTAIL.n271 0.155672
R729 VTAIL.n300 VTAIL.n299 0.155672
R730 VTAIL.n300 VTAIL.n267 0.155672
R731 VTAIL.n307 VTAIL.n267 0.155672
R732 VTAIL.n308 VTAIL.n307 0.155672
R733 VTAIL.n308 VTAIL.n263 0.155672
R734 VTAIL.n315 VTAIL.n263 0.155672
R735 VTAIL.n316 VTAIL.n315 0.155672
R736 VTAIL.n316 VTAIL.n259 0.155672
R737 VTAIL.n324 VTAIL.n259 0.155672
R738 VTAIL.n325 VTAIL.n324 0.155672
R739 VTAIL.n325 VTAIL.n255 0.155672
R740 VTAIL.n333 VTAIL.n255 0.155672
R741 VTAIL.n32 VTAIL.n31 0.155672
R742 VTAIL.n32 VTAIL.n23 0.155672
R743 VTAIL.n39 VTAIL.n23 0.155672
R744 VTAIL.n40 VTAIL.n39 0.155672
R745 VTAIL.n40 VTAIL.n19 0.155672
R746 VTAIL.n47 VTAIL.n19 0.155672
R747 VTAIL.n48 VTAIL.n47 0.155672
R748 VTAIL.n48 VTAIL.n15 0.155672
R749 VTAIL.n55 VTAIL.n15 0.155672
R750 VTAIL.n56 VTAIL.n55 0.155672
R751 VTAIL.n56 VTAIL.n11 0.155672
R752 VTAIL.n63 VTAIL.n11 0.155672
R753 VTAIL.n64 VTAIL.n63 0.155672
R754 VTAIL.n64 VTAIL.n7 0.155672
R755 VTAIL.n72 VTAIL.n7 0.155672
R756 VTAIL.n73 VTAIL.n72 0.155672
R757 VTAIL.n73 VTAIL.n3 0.155672
R758 VTAIL.n81 VTAIL.n3 0.155672
R759 VTAIL.n251 VTAIL.n173 0.155672
R760 VTAIL.n243 VTAIL.n173 0.155672
R761 VTAIL.n243 VTAIL.n242 0.155672
R762 VTAIL.n242 VTAIL.n177 0.155672
R763 VTAIL.n235 VTAIL.n177 0.155672
R764 VTAIL.n235 VTAIL.n234 0.155672
R765 VTAIL.n234 VTAIL.n182 0.155672
R766 VTAIL.n227 VTAIL.n182 0.155672
R767 VTAIL.n227 VTAIL.n226 0.155672
R768 VTAIL.n226 VTAIL.n186 0.155672
R769 VTAIL.n219 VTAIL.n186 0.155672
R770 VTAIL.n219 VTAIL.n218 0.155672
R771 VTAIL.n218 VTAIL.n190 0.155672
R772 VTAIL.n211 VTAIL.n190 0.155672
R773 VTAIL.n211 VTAIL.n210 0.155672
R774 VTAIL.n210 VTAIL.n194 0.155672
R775 VTAIL.n203 VTAIL.n194 0.155672
R776 VTAIL.n203 VTAIL.n202 0.155672
R777 VTAIL.n167 VTAIL.n89 0.155672
R778 VTAIL.n159 VTAIL.n89 0.155672
R779 VTAIL.n159 VTAIL.n158 0.155672
R780 VTAIL.n158 VTAIL.n93 0.155672
R781 VTAIL.n151 VTAIL.n93 0.155672
R782 VTAIL.n151 VTAIL.n150 0.155672
R783 VTAIL.n150 VTAIL.n98 0.155672
R784 VTAIL.n143 VTAIL.n98 0.155672
R785 VTAIL.n143 VTAIL.n142 0.155672
R786 VTAIL.n142 VTAIL.n102 0.155672
R787 VTAIL.n135 VTAIL.n102 0.155672
R788 VTAIL.n135 VTAIL.n134 0.155672
R789 VTAIL.n134 VTAIL.n106 0.155672
R790 VTAIL.n127 VTAIL.n106 0.155672
R791 VTAIL.n127 VTAIL.n126 0.155672
R792 VTAIL.n126 VTAIL.n110 0.155672
R793 VTAIL.n119 VTAIL.n110 0.155672
R794 VTAIL.n119 VTAIL.n118 0.155672
R795 B.n100 B.t17 644.125
R796 B.n98 B.t10 644.125
R797 B.n415 B.t6 644.125
R798 B.n413 B.t14 644.125
R799 B.n730 B.n729 585
R800 B.n731 B.n730 585
R801 B.n318 B.n97 585
R802 B.n317 B.n316 585
R803 B.n315 B.n314 585
R804 B.n313 B.n312 585
R805 B.n311 B.n310 585
R806 B.n309 B.n308 585
R807 B.n307 B.n306 585
R808 B.n305 B.n304 585
R809 B.n303 B.n302 585
R810 B.n301 B.n300 585
R811 B.n299 B.n298 585
R812 B.n297 B.n296 585
R813 B.n295 B.n294 585
R814 B.n293 B.n292 585
R815 B.n291 B.n290 585
R816 B.n289 B.n288 585
R817 B.n287 B.n286 585
R818 B.n285 B.n284 585
R819 B.n283 B.n282 585
R820 B.n281 B.n280 585
R821 B.n279 B.n278 585
R822 B.n277 B.n276 585
R823 B.n275 B.n274 585
R824 B.n273 B.n272 585
R825 B.n271 B.n270 585
R826 B.n269 B.n268 585
R827 B.n267 B.n266 585
R828 B.n265 B.n264 585
R829 B.n263 B.n262 585
R830 B.n261 B.n260 585
R831 B.n259 B.n258 585
R832 B.n257 B.n256 585
R833 B.n255 B.n254 585
R834 B.n253 B.n252 585
R835 B.n251 B.n250 585
R836 B.n249 B.n248 585
R837 B.n247 B.n246 585
R838 B.n245 B.n244 585
R839 B.n243 B.n242 585
R840 B.n241 B.n240 585
R841 B.n239 B.n238 585
R842 B.n237 B.n236 585
R843 B.n235 B.n234 585
R844 B.n233 B.n232 585
R845 B.n231 B.n230 585
R846 B.n229 B.n228 585
R847 B.n227 B.n226 585
R848 B.n225 B.n224 585
R849 B.n223 B.n222 585
R850 B.n220 B.n219 585
R851 B.n218 B.n217 585
R852 B.n216 B.n215 585
R853 B.n214 B.n213 585
R854 B.n212 B.n211 585
R855 B.n210 B.n209 585
R856 B.n208 B.n207 585
R857 B.n206 B.n205 585
R858 B.n204 B.n203 585
R859 B.n202 B.n201 585
R860 B.n200 B.n199 585
R861 B.n198 B.n197 585
R862 B.n196 B.n195 585
R863 B.n194 B.n193 585
R864 B.n192 B.n191 585
R865 B.n190 B.n189 585
R866 B.n188 B.n187 585
R867 B.n186 B.n185 585
R868 B.n184 B.n183 585
R869 B.n182 B.n181 585
R870 B.n180 B.n179 585
R871 B.n178 B.n177 585
R872 B.n176 B.n175 585
R873 B.n174 B.n173 585
R874 B.n172 B.n171 585
R875 B.n170 B.n169 585
R876 B.n168 B.n167 585
R877 B.n166 B.n165 585
R878 B.n164 B.n163 585
R879 B.n162 B.n161 585
R880 B.n160 B.n159 585
R881 B.n158 B.n157 585
R882 B.n156 B.n155 585
R883 B.n154 B.n153 585
R884 B.n152 B.n151 585
R885 B.n150 B.n149 585
R886 B.n148 B.n147 585
R887 B.n146 B.n145 585
R888 B.n144 B.n143 585
R889 B.n142 B.n141 585
R890 B.n140 B.n139 585
R891 B.n138 B.n137 585
R892 B.n136 B.n135 585
R893 B.n134 B.n133 585
R894 B.n132 B.n131 585
R895 B.n130 B.n129 585
R896 B.n128 B.n127 585
R897 B.n126 B.n125 585
R898 B.n124 B.n123 585
R899 B.n122 B.n121 585
R900 B.n120 B.n119 585
R901 B.n118 B.n117 585
R902 B.n116 B.n115 585
R903 B.n114 B.n113 585
R904 B.n112 B.n111 585
R905 B.n110 B.n109 585
R906 B.n108 B.n107 585
R907 B.n106 B.n105 585
R908 B.n104 B.n103 585
R909 B.n728 B.n42 585
R910 B.n732 B.n42 585
R911 B.n727 B.n41 585
R912 B.n733 B.n41 585
R913 B.n726 B.n725 585
R914 B.n725 B.n37 585
R915 B.n724 B.n36 585
R916 B.n739 B.n36 585
R917 B.n723 B.n35 585
R918 B.n740 B.n35 585
R919 B.n722 B.n34 585
R920 B.n741 B.n34 585
R921 B.n721 B.n720 585
R922 B.n720 B.n30 585
R923 B.n719 B.n29 585
R924 B.n747 B.n29 585
R925 B.n718 B.n28 585
R926 B.n748 B.n28 585
R927 B.n717 B.n27 585
R928 B.n749 B.n27 585
R929 B.n716 B.n715 585
R930 B.n715 B.n23 585
R931 B.n714 B.n22 585
R932 B.n755 B.n22 585
R933 B.n713 B.n21 585
R934 B.n756 B.n21 585
R935 B.n712 B.n20 585
R936 B.n757 B.n20 585
R937 B.n711 B.n710 585
R938 B.n710 B.n19 585
R939 B.n709 B.n15 585
R940 B.n763 B.n15 585
R941 B.n708 B.n14 585
R942 B.n764 B.n14 585
R943 B.n707 B.n13 585
R944 B.n765 B.n13 585
R945 B.n706 B.n705 585
R946 B.n705 B.n12 585
R947 B.n704 B.n703 585
R948 B.n704 B.n8 585
R949 B.n702 B.n7 585
R950 B.n772 B.n7 585
R951 B.n701 B.n6 585
R952 B.n773 B.n6 585
R953 B.n700 B.n5 585
R954 B.n774 B.n5 585
R955 B.n699 B.n698 585
R956 B.n698 B.n4 585
R957 B.n697 B.n319 585
R958 B.n697 B.n696 585
R959 B.n686 B.n320 585
R960 B.n689 B.n320 585
R961 B.n688 B.n687 585
R962 B.n690 B.n688 585
R963 B.n685 B.n325 585
R964 B.n325 B.n324 585
R965 B.n684 B.n683 585
R966 B.n683 B.n682 585
R967 B.n327 B.n326 585
R968 B.n675 B.n327 585
R969 B.n674 B.n673 585
R970 B.n676 B.n674 585
R971 B.n672 B.n332 585
R972 B.n332 B.n331 585
R973 B.n671 B.n670 585
R974 B.n670 B.n669 585
R975 B.n334 B.n333 585
R976 B.n335 B.n334 585
R977 B.n662 B.n661 585
R978 B.n663 B.n662 585
R979 B.n660 B.n340 585
R980 B.n340 B.n339 585
R981 B.n659 B.n658 585
R982 B.n658 B.n657 585
R983 B.n342 B.n341 585
R984 B.n343 B.n342 585
R985 B.n650 B.n649 585
R986 B.n651 B.n650 585
R987 B.n648 B.n348 585
R988 B.n348 B.n347 585
R989 B.n647 B.n646 585
R990 B.n646 B.n645 585
R991 B.n350 B.n349 585
R992 B.n351 B.n350 585
R993 B.n638 B.n637 585
R994 B.n639 B.n638 585
R995 B.n636 B.n356 585
R996 B.n356 B.n355 585
R997 B.n630 B.n629 585
R998 B.n628 B.n412 585
R999 B.n627 B.n411 585
R1000 B.n632 B.n411 585
R1001 B.n626 B.n625 585
R1002 B.n624 B.n623 585
R1003 B.n622 B.n621 585
R1004 B.n620 B.n619 585
R1005 B.n618 B.n617 585
R1006 B.n616 B.n615 585
R1007 B.n614 B.n613 585
R1008 B.n612 B.n611 585
R1009 B.n610 B.n609 585
R1010 B.n608 B.n607 585
R1011 B.n606 B.n605 585
R1012 B.n604 B.n603 585
R1013 B.n602 B.n601 585
R1014 B.n600 B.n599 585
R1015 B.n598 B.n597 585
R1016 B.n596 B.n595 585
R1017 B.n594 B.n593 585
R1018 B.n592 B.n591 585
R1019 B.n590 B.n589 585
R1020 B.n588 B.n587 585
R1021 B.n586 B.n585 585
R1022 B.n584 B.n583 585
R1023 B.n582 B.n581 585
R1024 B.n580 B.n579 585
R1025 B.n578 B.n577 585
R1026 B.n576 B.n575 585
R1027 B.n574 B.n573 585
R1028 B.n572 B.n571 585
R1029 B.n570 B.n569 585
R1030 B.n568 B.n567 585
R1031 B.n566 B.n565 585
R1032 B.n564 B.n563 585
R1033 B.n562 B.n561 585
R1034 B.n560 B.n559 585
R1035 B.n558 B.n557 585
R1036 B.n556 B.n555 585
R1037 B.n554 B.n553 585
R1038 B.n552 B.n551 585
R1039 B.n550 B.n549 585
R1040 B.n548 B.n547 585
R1041 B.n546 B.n545 585
R1042 B.n544 B.n543 585
R1043 B.n542 B.n541 585
R1044 B.n540 B.n539 585
R1045 B.n538 B.n537 585
R1046 B.n536 B.n535 585
R1047 B.n534 B.n533 585
R1048 B.n531 B.n530 585
R1049 B.n529 B.n528 585
R1050 B.n527 B.n526 585
R1051 B.n525 B.n524 585
R1052 B.n523 B.n522 585
R1053 B.n521 B.n520 585
R1054 B.n519 B.n518 585
R1055 B.n517 B.n516 585
R1056 B.n515 B.n514 585
R1057 B.n513 B.n512 585
R1058 B.n511 B.n510 585
R1059 B.n509 B.n508 585
R1060 B.n507 B.n506 585
R1061 B.n505 B.n504 585
R1062 B.n503 B.n502 585
R1063 B.n501 B.n500 585
R1064 B.n499 B.n498 585
R1065 B.n497 B.n496 585
R1066 B.n495 B.n494 585
R1067 B.n493 B.n492 585
R1068 B.n491 B.n490 585
R1069 B.n489 B.n488 585
R1070 B.n487 B.n486 585
R1071 B.n485 B.n484 585
R1072 B.n483 B.n482 585
R1073 B.n481 B.n480 585
R1074 B.n479 B.n478 585
R1075 B.n477 B.n476 585
R1076 B.n475 B.n474 585
R1077 B.n473 B.n472 585
R1078 B.n471 B.n470 585
R1079 B.n469 B.n468 585
R1080 B.n467 B.n466 585
R1081 B.n465 B.n464 585
R1082 B.n463 B.n462 585
R1083 B.n461 B.n460 585
R1084 B.n459 B.n458 585
R1085 B.n457 B.n456 585
R1086 B.n455 B.n454 585
R1087 B.n453 B.n452 585
R1088 B.n451 B.n450 585
R1089 B.n449 B.n448 585
R1090 B.n447 B.n446 585
R1091 B.n445 B.n444 585
R1092 B.n443 B.n442 585
R1093 B.n441 B.n440 585
R1094 B.n439 B.n438 585
R1095 B.n437 B.n436 585
R1096 B.n435 B.n434 585
R1097 B.n433 B.n432 585
R1098 B.n431 B.n430 585
R1099 B.n429 B.n428 585
R1100 B.n427 B.n426 585
R1101 B.n425 B.n424 585
R1102 B.n423 B.n422 585
R1103 B.n421 B.n420 585
R1104 B.n419 B.n418 585
R1105 B.n358 B.n357 585
R1106 B.n635 B.n634 585
R1107 B.n354 B.n353 585
R1108 B.n355 B.n354 585
R1109 B.n641 B.n640 585
R1110 B.n640 B.n639 585
R1111 B.n642 B.n352 585
R1112 B.n352 B.n351 585
R1113 B.n644 B.n643 585
R1114 B.n645 B.n644 585
R1115 B.n346 B.n345 585
R1116 B.n347 B.n346 585
R1117 B.n653 B.n652 585
R1118 B.n652 B.n651 585
R1119 B.n654 B.n344 585
R1120 B.n344 B.n343 585
R1121 B.n656 B.n655 585
R1122 B.n657 B.n656 585
R1123 B.n338 B.n337 585
R1124 B.n339 B.n338 585
R1125 B.n665 B.n664 585
R1126 B.n664 B.n663 585
R1127 B.n666 B.n336 585
R1128 B.n336 B.n335 585
R1129 B.n668 B.n667 585
R1130 B.n669 B.n668 585
R1131 B.n330 B.n329 585
R1132 B.n331 B.n330 585
R1133 B.n678 B.n677 585
R1134 B.n677 B.n676 585
R1135 B.n679 B.n328 585
R1136 B.n675 B.n328 585
R1137 B.n681 B.n680 585
R1138 B.n682 B.n681 585
R1139 B.n323 B.n322 585
R1140 B.n324 B.n323 585
R1141 B.n692 B.n691 585
R1142 B.n691 B.n690 585
R1143 B.n693 B.n321 585
R1144 B.n689 B.n321 585
R1145 B.n695 B.n694 585
R1146 B.n696 B.n695 585
R1147 B.n3 B.n0 585
R1148 B.n4 B.n3 585
R1149 B.n771 B.n1 585
R1150 B.n772 B.n771 585
R1151 B.n770 B.n769 585
R1152 B.n770 B.n8 585
R1153 B.n768 B.n9 585
R1154 B.n12 B.n9 585
R1155 B.n767 B.n766 585
R1156 B.n766 B.n765 585
R1157 B.n11 B.n10 585
R1158 B.n764 B.n11 585
R1159 B.n762 B.n761 585
R1160 B.n763 B.n762 585
R1161 B.n760 B.n16 585
R1162 B.n19 B.n16 585
R1163 B.n759 B.n758 585
R1164 B.n758 B.n757 585
R1165 B.n18 B.n17 585
R1166 B.n756 B.n18 585
R1167 B.n754 B.n753 585
R1168 B.n755 B.n754 585
R1169 B.n752 B.n24 585
R1170 B.n24 B.n23 585
R1171 B.n751 B.n750 585
R1172 B.n750 B.n749 585
R1173 B.n26 B.n25 585
R1174 B.n748 B.n26 585
R1175 B.n746 B.n745 585
R1176 B.n747 B.n746 585
R1177 B.n744 B.n31 585
R1178 B.n31 B.n30 585
R1179 B.n743 B.n742 585
R1180 B.n742 B.n741 585
R1181 B.n33 B.n32 585
R1182 B.n740 B.n33 585
R1183 B.n738 B.n737 585
R1184 B.n739 B.n738 585
R1185 B.n736 B.n38 585
R1186 B.n38 B.n37 585
R1187 B.n735 B.n734 585
R1188 B.n734 B.n733 585
R1189 B.n40 B.n39 585
R1190 B.n732 B.n40 585
R1191 B.n775 B.n774 585
R1192 B.n773 B.n2 585
R1193 B.n103 B.n40 449.257
R1194 B.n730 B.n42 449.257
R1195 B.n634 B.n356 449.257
R1196 B.n630 B.n354 449.257
R1197 B.n100 B.t18 349.998
R1198 B.n98 B.t12 349.998
R1199 B.n415 B.t9 349.998
R1200 B.n413 B.t16 349.998
R1201 B.n99 B.t13 328.082
R1202 B.n416 B.t8 328.082
R1203 B.n101 B.t19 328.082
R1204 B.n414 B.t15 328.082
R1205 B.n731 B.n96 256.663
R1206 B.n731 B.n95 256.663
R1207 B.n731 B.n94 256.663
R1208 B.n731 B.n93 256.663
R1209 B.n731 B.n92 256.663
R1210 B.n731 B.n91 256.663
R1211 B.n731 B.n90 256.663
R1212 B.n731 B.n89 256.663
R1213 B.n731 B.n88 256.663
R1214 B.n731 B.n87 256.663
R1215 B.n731 B.n86 256.663
R1216 B.n731 B.n85 256.663
R1217 B.n731 B.n84 256.663
R1218 B.n731 B.n83 256.663
R1219 B.n731 B.n82 256.663
R1220 B.n731 B.n81 256.663
R1221 B.n731 B.n80 256.663
R1222 B.n731 B.n79 256.663
R1223 B.n731 B.n78 256.663
R1224 B.n731 B.n77 256.663
R1225 B.n731 B.n76 256.663
R1226 B.n731 B.n75 256.663
R1227 B.n731 B.n74 256.663
R1228 B.n731 B.n73 256.663
R1229 B.n731 B.n72 256.663
R1230 B.n731 B.n71 256.663
R1231 B.n731 B.n70 256.663
R1232 B.n731 B.n69 256.663
R1233 B.n731 B.n68 256.663
R1234 B.n731 B.n67 256.663
R1235 B.n731 B.n66 256.663
R1236 B.n731 B.n65 256.663
R1237 B.n731 B.n64 256.663
R1238 B.n731 B.n63 256.663
R1239 B.n731 B.n62 256.663
R1240 B.n731 B.n61 256.663
R1241 B.n731 B.n60 256.663
R1242 B.n731 B.n59 256.663
R1243 B.n731 B.n58 256.663
R1244 B.n731 B.n57 256.663
R1245 B.n731 B.n56 256.663
R1246 B.n731 B.n55 256.663
R1247 B.n731 B.n54 256.663
R1248 B.n731 B.n53 256.663
R1249 B.n731 B.n52 256.663
R1250 B.n731 B.n51 256.663
R1251 B.n731 B.n50 256.663
R1252 B.n731 B.n49 256.663
R1253 B.n731 B.n48 256.663
R1254 B.n731 B.n47 256.663
R1255 B.n731 B.n46 256.663
R1256 B.n731 B.n45 256.663
R1257 B.n731 B.n44 256.663
R1258 B.n731 B.n43 256.663
R1259 B.n632 B.n631 256.663
R1260 B.n632 B.n359 256.663
R1261 B.n632 B.n360 256.663
R1262 B.n632 B.n361 256.663
R1263 B.n632 B.n362 256.663
R1264 B.n632 B.n363 256.663
R1265 B.n632 B.n364 256.663
R1266 B.n632 B.n365 256.663
R1267 B.n632 B.n366 256.663
R1268 B.n632 B.n367 256.663
R1269 B.n632 B.n368 256.663
R1270 B.n632 B.n369 256.663
R1271 B.n632 B.n370 256.663
R1272 B.n632 B.n371 256.663
R1273 B.n632 B.n372 256.663
R1274 B.n632 B.n373 256.663
R1275 B.n632 B.n374 256.663
R1276 B.n632 B.n375 256.663
R1277 B.n632 B.n376 256.663
R1278 B.n632 B.n377 256.663
R1279 B.n632 B.n378 256.663
R1280 B.n632 B.n379 256.663
R1281 B.n632 B.n380 256.663
R1282 B.n632 B.n381 256.663
R1283 B.n632 B.n382 256.663
R1284 B.n632 B.n383 256.663
R1285 B.n632 B.n384 256.663
R1286 B.n632 B.n385 256.663
R1287 B.n632 B.n386 256.663
R1288 B.n632 B.n387 256.663
R1289 B.n632 B.n388 256.663
R1290 B.n632 B.n389 256.663
R1291 B.n632 B.n390 256.663
R1292 B.n632 B.n391 256.663
R1293 B.n632 B.n392 256.663
R1294 B.n632 B.n393 256.663
R1295 B.n632 B.n394 256.663
R1296 B.n632 B.n395 256.663
R1297 B.n632 B.n396 256.663
R1298 B.n632 B.n397 256.663
R1299 B.n632 B.n398 256.663
R1300 B.n632 B.n399 256.663
R1301 B.n632 B.n400 256.663
R1302 B.n632 B.n401 256.663
R1303 B.n632 B.n402 256.663
R1304 B.n632 B.n403 256.663
R1305 B.n632 B.n404 256.663
R1306 B.n632 B.n405 256.663
R1307 B.n632 B.n406 256.663
R1308 B.n632 B.n407 256.663
R1309 B.n632 B.n408 256.663
R1310 B.n632 B.n409 256.663
R1311 B.n632 B.n410 256.663
R1312 B.n633 B.n632 256.663
R1313 B.n777 B.n776 256.663
R1314 B.n107 B.n106 163.367
R1315 B.n111 B.n110 163.367
R1316 B.n115 B.n114 163.367
R1317 B.n119 B.n118 163.367
R1318 B.n123 B.n122 163.367
R1319 B.n127 B.n126 163.367
R1320 B.n131 B.n130 163.367
R1321 B.n135 B.n134 163.367
R1322 B.n139 B.n138 163.367
R1323 B.n143 B.n142 163.367
R1324 B.n147 B.n146 163.367
R1325 B.n151 B.n150 163.367
R1326 B.n155 B.n154 163.367
R1327 B.n159 B.n158 163.367
R1328 B.n163 B.n162 163.367
R1329 B.n167 B.n166 163.367
R1330 B.n171 B.n170 163.367
R1331 B.n175 B.n174 163.367
R1332 B.n179 B.n178 163.367
R1333 B.n183 B.n182 163.367
R1334 B.n187 B.n186 163.367
R1335 B.n191 B.n190 163.367
R1336 B.n195 B.n194 163.367
R1337 B.n199 B.n198 163.367
R1338 B.n203 B.n202 163.367
R1339 B.n207 B.n206 163.367
R1340 B.n211 B.n210 163.367
R1341 B.n215 B.n214 163.367
R1342 B.n219 B.n218 163.367
R1343 B.n224 B.n223 163.367
R1344 B.n228 B.n227 163.367
R1345 B.n232 B.n231 163.367
R1346 B.n236 B.n235 163.367
R1347 B.n240 B.n239 163.367
R1348 B.n244 B.n243 163.367
R1349 B.n248 B.n247 163.367
R1350 B.n252 B.n251 163.367
R1351 B.n256 B.n255 163.367
R1352 B.n260 B.n259 163.367
R1353 B.n264 B.n263 163.367
R1354 B.n268 B.n267 163.367
R1355 B.n272 B.n271 163.367
R1356 B.n276 B.n275 163.367
R1357 B.n280 B.n279 163.367
R1358 B.n284 B.n283 163.367
R1359 B.n288 B.n287 163.367
R1360 B.n292 B.n291 163.367
R1361 B.n296 B.n295 163.367
R1362 B.n300 B.n299 163.367
R1363 B.n304 B.n303 163.367
R1364 B.n308 B.n307 163.367
R1365 B.n312 B.n311 163.367
R1366 B.n316 B.n315 163.367
R1367 B.n730 B.n97 163.367
R1368 B.n638 B.n356 163.367
R1369 B.n638 B.n350 163.367
R1370 B.n646 B.n350 163.367
R1371 B.n646 B.n348 163.367
R1372 B.n650 B.n348 163.367
R1373 B.n650 B.n342 163.367
R1374 B.n658 B.n342 163.367
R1375 B.n658 B.n340 163.367
R1376 B.n662 B.n340 163.367
R1377 B.n662 B.n334 163.367
R1378 B.n670 B.n334 163.367
R1379 B.n670 B.n332 163.367
R1380 B.n674 B.n332 163.367
R1381 B.n674 B.n327 163.367
R1382 B.n683 B.n327 163.367
R1383 B.n683 B.n325 163.367
R1384 B.n688 B.n325 163.367
R1385 B.n688 B.n320 163.367
R1386 B.n697 B.n320 163.367
R1387 B.n698 B.n697 163.367
R1388 B.n698 B.n5 163.367
R1389 B.n6 B.n5 163.367
R1390 B.n7 B.n6 163.367
R1391 B.n704 B.n7 163.367
R1392 B.n705 B.n704 163.367
R1393 B.n705 B.n13 163.367
R1394 B.n14 B.n13 163.367
R1395 B.n15 B.n14 163.367
R1396 B.n710 B.n15 163.367
R1397 B.n710 B.n20 163.367
R1398 B.n21 B.n20 163.367
R1399 B.n22 B.n21 163.367
R1400 B.n715 B.n22 163.367
R1401 B.n715 B.n27 163.367
R1402 B.n28 B.n27 163.367
R1403 B.n29 B.n28 163.367
R1404 B.n720 B.n29 163.367
R1405 B.n720 B.n34 163.367
R1406 B.n35 B.n34 163.367
R1407 B.n36 B.n35 163.367
R1408 B.n725 B.n36 163.367
R1409 B.n725 B.n41 163.367
R1410 B.n42 B.n41 163.367
R1411 B.n412 B.n411 163.367
R1412 B.n625 B.n411 163.367
R1413 B.n623 B.n622 163.367
R1414 B.n619 B.n618 163.367
R1415 B.n615 B.n614 163.367
R1416 B.n611 B.n610 163.367
R1417 B.n607 B.n606 163.367
R1418 B.n603 B.n602 163.367
R1419 B.n599 B.n598 163.367
R1420 B.n595 B.n594 163.367
R1421 B.n591 B.n590 163.367
R1422 B.n587 B.n586 163.367
R1423 B.n583 B.n582 163.367
R1424 B.n579 B.n578 163.367
R1425 B.n575 B.n574 163.367
R1426 B.n571 B.n570 163.367
R1427 B.n567 B.n566 163.367
R1428 B.n563 B.n562 163.367
R1429 B.n559 B.n558 163.367
R1430 B.n555 B.n554 163.367
R1431 B.n551 B.n550 163.367
R1432 B.n547 B.n546 163.367
R1433 B.n543 B.n542 163.367
R1434 B.n539 B.n538 163.367
R1435 B.n535 B.n534 163.367
R1436 B.n530 B.n529 163.367
R1437 B.n526 B.n525 163.367
R1438 B.n522 B.n521 163.367
R1439 B.n518 B.n517 163.367
R1440 B.n514 B.n513 163.367
R1441 B.n510 B.n509 163.367
R1442 B.n506 B.n505 163.367
R1443 B.n502 B.n501 163.367
R1444 B.n498 B.n497 163.367
R1445 B.n494 B.n493 163.367
R1446 B.n490 B.n489 163.367
R1447 B.n486 B.n485 163.367
R1448 B.n482 B.n481 163.367
R1449 B.n478 B.n477 163.367
R1450 B.n474 B.n473 163.367
R1451 B.n470 B.n469 163.367
R1452 B.n466 B.n465 163.367
R1453 B.n462 B.n461 163.367
R1454 B.n458 B.n457 163.367
R1455 B.n454 B.n453 163.367
R1456 B.n450 B.n449 163.367
R1457 B.n446 B.n445 163.367
R1458 B.n442 B.n441 163.367
R1459 B.n438 B.n437 163.367
R1460 B.n434 B.n433 163.367
R1461 B.n430 B.n429 163.367
R1462 B.n426 B.n425 163.367
R1463 B.n422 B.n421 163.367
R1464 B.n418 B.n358 163.367
R1465 B.n640 B.n354 163.367
R1466 B.n640 B.n352 163.367
R1467 B.n644 B.n352 163.367
R1468 B.n644 B.n346 163.367
R1469 B.n652 B.n346 163.367
R1470 B.n652 B.n344 163.367
R1471 B.n656 B.n344 163.367
R1472 B.n656 B.n338 163.367
R1473 B.n664 B.n338 163.367
R1474 B.n664 B.n336 163.367
R1475 B.n668 B.n336 163.367
R1476 B.n668 B.n330 163.367
R1477 B.n677 B.n330 163.367
R1478 B.n677 B.n328 163.367
R1479 B.n681 B.n328 163.367
R1480 B.n681 B.n323 163.367
R1481 B.n691 B.n323 163.367
R1482 B.n691 B.n321 163.367
R1483 B.n695 B.n321 163.367
R1484 B.n695 B.n3 163.367
R1485 B.n775 B.n3 163.367
R1486 B.n771 B.n2 163.367
R1487 B.n771 B.n770 163.367
R1488 B.n770 B.n9 163.367
R1489 B.n766 B.n9 163.367
R1490 B.n766 B.n11 163.367
R1491 B.n762 B.n11 163.367
R1492 B.n762 B.n16 163.367
R1493 B.n758 B.n16 163.367
R1494 B.n758 B.n18 163.367
R1495 B.n754 B.n18 163.367
R1496 B.n754 B.n24 163.367
R1497 B.n750 B.n24 163.367
R1498 B.n750 B.n26 163.367
R1499 B.n746 B.n26 163.367
R1500 B.n746 B.n31 163.367
R1501 B.n742 B.n31 163.367
R1502 B.n742 B.n33 163.367
R1503 B.n738 B.n33 163.367
R1504 B.n738 B.n38 163.367
R1505 B.n734 B.n38 163.367
R1506 B.n734 B.n40 163.367
R1507 B.n103 B.n43 71.676
R1508 B.n107 B.n44 71.676
R1509 B.n111 B.n45 71.676
R1510 B.n115 B.n46 71.676
R1511 B.n119 B.n47 71.676
R1512 B.n123 B.n48 71.676
R1513 B.n127 B.n49 71.676
R1514 B.n131 B.n50 71.676
R1515 B.n135 B.n51 71.676
R1516 B.n139 B.n52 71.676
R1517 B.n143 B.n53 71.676
R1518 B.n147 B.n54 71.676
R1519 B.n151 B.n55 71.676
R1520 B.n155 B.n56 71.676
R1521 B.n159 B.n57 71.676
R1522 B.n163 B.n58 71.676
R1523 B.n167 B.n59 71.676
R1524 B.n171 B.n60 71.676
R1525 B.n175 B.n61 71.676
R1526 B.n179 B.n62 71.676
R1527 B.n183 B.n63 71.676
R1528 B.n187 B.n64 71.676
R1529 B.n191 B.n65 71.676
R1530 B.n195 B.n66 71.676
R1531 B.n199 B.n67 71.676
R1532 B.n203 B.n68 71.676
R1533 B.n207 B.n69 71.676
R1534 B.n211 B.n70 71.676
R1535 B.n215 B.n71 71.676
R1536 B.n219 B.n72 71.676
R1537 B.n224 B.n73 71.676
R1538 B.n228 B.n74 71.676
R1539 B.n232 B.n75 71.676
R1540 B.n236 B.n76 71.676
R1541 B.n240 B.n77 71.676
R1542 B.n244 B.n78 71.676
R1543 B.n248 B.n79 71.676
R1544 B.n252 B.n80 71.676
R1545 B.n256 B.n81 71.676
R1546 B.n260 B.n82 71.676
R1547 B.n264 B.n83 71.676
R1548 B.n268 B.n84 71.676
R1549 B.n272 B.n85 71.676
R1550 B.n276 B.n86 71.676
R1551 B.n280 B.n87 71.676
R1552 B.n284 B.n88 71.676
R1553 B.n288 B.n89 71.676
R1554 B.n292 B.n90 71.676
R1555 B.n296 B.n91 71.676
R1556 B.n300 B.n92 71.676
R1557 B.n304 B.n93 71.676
R1558 B.n308 B.n94 71.676
R1559 B.n312 B.n95 71.676
R1560 B.n316 B.n96 71.676
R1561 B.n97 B.n96 71.676
R1562 B.n315 B.n95 71.676
R1563 B.n311 B.n94 71.676
R1564 B.n307 B.n93 71.676
R1565 B.n303 B.n92 71.676
R1566 B.n299 B.n91 71.676
R1567 B.n295 B.n90 71.676
R1568 B.n291 B.n89 71.676
R1569 B.n287 B.n88 71.676
R1570 B.n283 B.n87 71.676
R1571 B.n279 B.n86 71.676
R1572 B.n275 B.n85 71.676
R1573 B.n271 B.n84 71.676
R1574 B.n267 B.n83 71.676
R1575 B.n263 B.n82 71.676
R1576 B.n259 B.n81 71.676
R1577 B.n255 B.n80 71.676
R1578 B.n251 B.n79 71.676
R1579 B.n247 B.n78 71.676
R1580 B.n243 B.n77 71.676
R1581 B.n239 B.n76 71.676
R1582 B.n235 B.n75 71.676
R1583 B.n231 B.n74 71.676
R1584 B.n227 B.n73 71.676
R1585 B.n223 B.n72 71.676
R1586 B.n218 B.n71 71.676
R1587 B.n214 B.n70 71.676
R1588 B.n210 B.n69 71.676
R1589 B.n206 B.n68 71.676
R1590 B.n202 B.n67 71.676
R1591 B.n198 B.n66 71.676
R1592 B.n194 B.n65 71.676
R1593 B.n190 B.n64 71.676
R1594 B.n186 B.n63 71.676
R1595 B.n182 B.n62 71.676
R1596 B.n178 B.n61 71.676
R1597 B.n174 B.n60 71.676
R1598 B.n170 B.n59 71.676
R1599 B.n166 B.n58 71.676
R1600 B.n162 B.n57 71.676
R1601 B.n158 B.n56 71.676
R1602 B.n154 B.n55 71.676
R1603 B.n150 B.n54 71.676
R1604 B.n146 B.n53 71.676
R1605 B.n142 B.n52 71.676
R1606 B.n138 B.n51 71.676
R1607 B.n134 B.n50 71.676
R1608 B.n130 B.n49 71.676
R1609 B.n126 B.n48 71.676
R1610 B.n122 B.n47 71.676
R1611 B.n118 B.n46 71.676
R1612 B.n114 B.n45 71.676
R1613 B.n110 B.n44 71.676
R1614 B.n106 B.n43 71.676
R1615 B.n631 B.n630 71.676
R1616 B.n625 B.n359 71.676
R1617 B.n622 B.n360 71.676
R1618 B.n618 B.n361 71.676
R1619 B.n614 B.n362 71.676
R1620 B.n610 B.n363 71.676
R1621 B.n606 B.n364 71.676
R1622 B.n602 B.n365 71.676
R1623 B.n598 B.n366 71.676
R1624 B.n594 B.n367 71.676
R1625 B.n590 B.n368 71.676
R1626 B.n586 B.n369 71.676
R1627 B.n582 B.n370 71.676
R1628 B.n578 B.n371 71.676
R1629 B.n574 B.n372 71.676
R1630 B.n570 B.n373 71.676
R1631 B.n566 B.n374 71.676
R1632 B.n562 B.n375 71.676
R1633 B.n558 B.n376 71.676
R1634 B.n554 B.n377 71.676
R1635 B.n550 B.n378 71.676
R1636 B.n546 B.n379 71.676
R1637 B.n542 B.n380 71.676
R1638 B.n538 B.n381 71.676
R1639 B.n534 B.n382 71.676
R1640 B.n529 B.n383 71.676
R1641 B.n525 B.n384 71.676
R1642 B.n521 B.n385 71.676
R1643 B.n517 B.n386 71.676
R1644 B.n513 B.n387 71.676
R1645 B.n509 B.n388 71.676
R1646 B.n505 B.n389 71.676
R1647 B.n501 B.n390 71.676
R1648 B.n497 B.n391 71.676
R1649 B.n493 B.n392 71.676
R1650 B.n489 B.n393 71.676
R1651 B.n485 B.n394 71.676
R1652 B.n481 B.n395 71.676
R1653 B.n477 B.n396 71.676
R1654 B.n473 B.n397 71.676
R1655 B.n469 B.n398 71.676
R1656 B.n465 B.n399 71.676
R1657 B.n461 B.n400 71.676
R1658 B.n457 B.n401 71.676
R1659 B.n453 B.n402 71.676
R1660 B.n449 B.n403 71.676
R1661 B.n445 B.n404 71.676
R1662 B.n441 B.n405 71.676
R1663 B.n437 B.n406 71.676
R1664 B.n433 B.n407 71.676
R1665 B.n429 B.n408 71.676
R1666 B.n425 B.n409 71.676
R1667 B.n421 B.n410 71.676
R1668 B.n633 B.n358 71.676
R1669 B.n631 B.n412 71.676
R1670 B.n623 B.n359 71.676
R1671 B.n619 B.n360 71.676
R1672 B.n615 B.n361 71.676
R1673 B.n611 B.n362 71.676
R1674 B.n607 B.n363 71.676
R1675 B.n603 B.n364 71.676
R1676 B.n599 B.n365 71.676
R1677 B.n595 B.n366 71.676
R1678 B.n591 B.n367 71.676
R1679 B.n587 B.n368 71.676
R1680 B.n583 B.n369 71.676
R1681 B.n579 B.n370 71.676
R1682 B.n575 B.n371 71.676
R1683 B.n571 B.n372 71.676
R1684 B.n567 B.n373 71.676
R1685 B.n563 B.n374 71.676
R1686 B.n559 B.n375 71.676
R1687 B.n555 B.n376 71.676
R1688 B.n551 B.n377 71.676
R1689 B.n547 B.n378 71.676
R1690 B.n543 B.n379 71.676
R1691 B.n539 B.n380 71.676
R1692 B.n535 B.n381 71.676
R1693 B.n530 B.n382 71.676
R1694 B.n526 B.n383 71.676
R1695 B.n522 B.n384 71.676
R1696 B.n518 B.n385 71.676
R1697 B.n514 B.n386 71.676
R1698 B.n510 B.n387 71.676
R1699 B.n506 B.n388 71.676
R1700 B.n502 B.n389 71.676
R1701 B.n498 B.n390 71.676
R1702 B.n494 B.n391 71.676
R1703 B.n490 B.n392 71.676
R1704 B.n486 B.n393 71.676
R1705 B.n482 B.n394 71.676
R1706 B.n478 B.n395 71.676
R1707 B.n474 B.n396 71.676
R1708 B.n470 B.n397 71.676
R1709 B.n466 B.n398 71.676
R1710 B.n462 B.n399 71.676
R1711 B.n458 B.n400 71.676
R1712 B.n454 B.n401 71.676
R1713 B.n450 B.n402 71.676
R1714 B.n446 B.n403 71.676
R1715 B.n442 B.n404 71.676
R1716 B.n438 B.n405 71.676
R1717 B.n434 B.n406 71.676
R1718 B.n430 B.n407 71.676
R1719 B.n426 B.n408 71.676
R1720 B.n422 B.n409 71.676
R1721 B.n418 B.n410 71.676
R1722 B.n634 B.n633 71.676
R1723 B.n776 B.n775 71.676
R1724 B.n776 B.n2 71.676
R1725 B.n632 B.n355 64.4956
R1726 B.n732 B.n731 64.4956
R1727 B.n102 B.n101 59.5399
R1728 B.n221 B.n99 59.5399
R1729 B.n417 B.n416 59.5399
R1730 B.n532 B.n414 59.5399
R1731 B.n639 B.n355 37.4848
R1732 B.n639 B.n351 37.4848
R1733 B.n645 B.n351 37.4848
R1734 B.n645 B.n347 37.4848
R1735 B.n651 B.n347 37.4848
R1736 B.n657 B.n343 37.4848
R1737 B.n657 B.n339 37.4848
R1738 B.n663 B.n339 37.4848
R1739 B.n663 B.n335 37.4848
R1740 B.n669 B.n335 37.4848
R1741 B.n676 B.n331 37.4848
R1742 B.n676 B.n675 37.4848
R1743 B.n682 B.n324 37.4848
R1744 B.n690 B.n324 37.4848
R1745 B.n690 B.n689 37.4848
R1746 B.n696 B.n4 37.4848
R1747 B.n774 B.n4 37.4848
R1748 B.n774 B.n773 37.4848
R1749 B.n773 B.n772 37.4848
R1750 B.n772 B.n8 37.4848
R1751 B.n765 B.n12 37.4848
R1752 B.n765 B.n764 37.4848
R1753 B.n764 B.n763 37.4848
R1754 B.n757 B.n19 37.4848
R1755 B.n757 B.n756 37.4848
R1756 B.n755 B.n23 37.4848
R1757 B.n749 B.n23 37.4848
R1758 B.n749 B.n748 37.4848
R1759 B.n748 B.n747 37.4848
R1760 B.n747 B.n30 37.4848
R1761 B.n741 B.n740 37.4848
R1762 B.n740 B.n739 37.4848
R1763 B.n739 B.n37 37.4848
R1764 B.n733 B.n37 37.4848
R1765 B.n733 B.n732 37.4848
R1766 B.t7 B.n343 35.2799
R1767 B.t11 B.n30 35.2799
R1768 B.n675 B.t4 34.1774
R1769 B.n19 B.t1 34.1774
R1770 B.n729 B.n728 29.1907
R1771 B.n629 B.n353 29.1907
R1772 B.n636 B.n635 29.1907
R1773 B.n104 B.n39 29.1907
R1774 B.n696 B.t2 28.665
R1775 B.t0 B.n8 28.665
R1776 B.n669 B.t5 22.0501
R1777 B.t3 B.n755 22.0501
R1778 B.n101 B.n100 21.9157
R1779 B.n99 B.n98 21.9157
R1780 B.n416 B.n415 21.9157
R1781 B.n414 B.n413 21.9157
R1782 B B.n777 18.0485
R1783 B.t5 B.n331 15.4352
R1784 B.n756 B.t3 15.4352
R1785 B.n641 B.n353 10.6151
R1786 B.n642 B.n641 10.6151
R1787 B.n643 B.n642 10.6151
R1788 B.n643 B.n345 10.6151
R1789 B.n653 B.n345 10.6151
R1790 B.n654 B.n653 10.6151
R1791 B.n655 B.n654 10.6151
R1792 B.n655 B.n337 10.6151
R1793 B.n665 B.n337 10.6151
R1794 B.n666 B.n665 10.6151
R1795 B.n667 B.n666 10.6151
R1796 B.n667 B.n329 10.6151
R1797 B.n678 B.n329 10.6151
R1798 B.n679 B.n678 10.6151
R1799 B.n680 B.n679 10.6151
R1800 B.n680 B.n322 10.6151
R1801 B.n692 B.n322 10.6151
R1802 B.n693 B.n692 10.6151
R1803 B.n694 B.n693 10.6151
R1804 B.n694 B.n0 10.6151
R1805 B.n629 B.n628 10.6151
R1806 B.n628 B.n627 10.6151
R1807 B.n627 B.n626 10.6151
R1808 B.n626 B.n624 10.6151
R1809 B.n624 B.n621 10.6151
R1810 B.n621 B.n620 10.6151
R1811 B.n620 B.n617 10.6151
R1812 B.n617 B.n616 10.6151
R1813 B.n616 B.n613 10.6151
R1814 B.n613 B.n612 10.6151
R1815 B.n612 B.n609 10.6151
R1816 B.n609 B.n608 10.6151
R1817 B.n608 B.n605 10.6151
R1818 B.n605 B.n604 10.6151
R1819 B.n604 B.n601 10.6151
R1820 B.n601 B.n600 10.6151
R1821 B.n600 B.n597 10.6151
R1822 B.n597 B.n596 10.6151
R1823 B.n596 B.n593 10.6151
R1824 B.n593 B.n592 10.6151
R1825 B.n592 B.n589 10.6151
R1826 B.n589 B.n588 10.6151
R1827 B.n588 B.n585 10.6151
R1828 B.n585 B.n584 10.6151
R1829 B.n584 B.n581 10.6151
R1830 B.n581 B.n580 10.6151
R1831 B.n580 B.n577 10.6151
R1832 B.n577 B.n576 10.6151
R1833 B.n576 B.n573 10.6151
R1834 B.n573 B.n572 10.6151
R1835 B.n572 B.n569 10.6151
R1836 B.n569 B.n568 10.6151
R1837 B.n568 B.n565 10.6151
R1838 B.n565 B.n564 10.6151
R1839 B.n564 B.n561 10.6151
R1840 B.n561 B.n560 10.6151
R1841 B.n560 B.n557 10.6151
R1842 B.n557 B.n556 10.6151
R1843 B.n556 B.n553 10.6151
R1844 B.n553 B.n552 10.6151
R1845 B.n552 B.n549 10.6151
R1846 B.n549 B.n548 10.6151
R1847 B.n548 B.n545 10.6151
R1848 B.n545 B.n544 10.6151
R1849 B.n544 B.n541 10.6151
R1850 B.n541 B.n540 10.6151
R1851 B.n540 B.n537 10.6151
R1852 B.n537 B.n536 10.6151
R1853 B.n536 B.n533 10.6151
R1854 B.n531 B.n528 10.6151
R1855 B.n528 B.n527 10.6151
R1856 B.n527 B.n524 10.6151
R1857 B.n524 B.n523 10.6151
R1858 B.n523 B.n520 10.6151
R1859 B.n520 B.n519 10.6151
R1860 B.n519 B.n516 10.6151
R1861 B.n516 B.n515 10.6151
R1862 B.n512 B.n511 10.6151
R1863 B.n511 B.n508 10.6151
R1864 B.n508 B.n507 10.6151
R1865 B.n507 B.n504 10.6151
R1866 B.n504 B.n503 10.6151
R1867 B.n503 B.n500 10.6151
R1868 B.n500 B.n499 10.6151
R1869 B.n499 B.n496 10.6151
R1870 B.n496 B.n495 10.6151
R1871 B.n495 B.n492 10.6151
R1872 B.n492 B.n491 10.6151
R1873 B.n491 B.n488 10.6151
R1874 B.n488 B.n487 10.6151
R1875 B.n487 B.n484 10.6151
R1876 B.n484 B.n483 10.6151
R1877 B.n483 B.n480 10.6151
R1878 B.n480 B.n479 10.6151
R1879 B.n479 B.n476 10.6151
R1880 B.n476 B.n475 10.6151
R1881 B.n475 B.n472 10.6151
R1882 B.n472 B.n471 10.6151
R1883 B.n471 B.n468 10.6151
R1884 B.n468 B.n467 10.6151
R1885 B.n467 B.n464 10.6151
R1886 B.n464 B.n463 10.6151
R1887 B.n463 B.n460 10.6151
R1888 B.n460 B.n459 10.6151
R1889 B.n459 B.n456 10.6151
R1890 B.n456 B.n455 10.6151
R1891 B.n455 B.n452 10.6151
R1892 B.n452 B.n451 10.6151
R1893 B.n451 B.n448 10.6151
R1894 B.n448 B.n447 10.6151
R1895 B.n447 B.n444 10.6151
R1896 B.n444 B.n443 10.6151
R1897 B.n443 B.n440 10.6151
R1898 B.n440 B.n439 10.6151
R1899 B.n439 B.n436 10.6151
R1900 B.n436 B.n435 10.6151
R1901 B.n435 B.n432 10.6151
R1902 B.n432 B.n431 10.6151
R1903 B.n431 B.n428 10.6151
R1904 B.n428 B.n427 10.6151
R1905 B.n427 B.n424 10.6151
R1906 B.n424 B.n423 10.6151
R1907 B.n423 B.n420 10.6151
R1908 B.n420 B.n419 10.6151
R1909 B.n419 B.n357 10.6151
R1910 B.n635 B.n357 10.6151
R1911 B.n637 B.n636 10.6151
R1912 B.n637 B.n349 10.6151
R1913 B.n647 B.n349 10.6151
R1914 B.n648 B.n647 10.6151
R1915 B.n649 B.n648 10.6151
R1916 B.n649 B.n341 10.6151
R1917 B.n659 B.n341 10.6151
R1918 B.n660 B.n659 10.6151
R1919 B.n661 B.n660 10.6151
R1920 B.n661 B.n333 10.6151
R1921 B.n671 B.n333 10.6151
R1922 B.n672 B.n671 10.6151
R1923 B.n673 B.n672 10.6151
R1924 B.n673 B.n326 10.6151
R1925 B.n684 B.n326 10.6151
R1926 B.n685 B.n684 10.6151
R1927 B.n687 B.n685 10.6151
R1928 B.n687 B.n686 10.6151
R1929 B.n686 B.n319 10.6151
R1930 B.n699 B.n319 10.6151
R1931 B.n700 B.n699 10.6151
R1932 B.n701 B.n700 10.6151
R1933 B.n702 B.n701 10.6151
R1934 B.n703 B.n702 10.6151
R1935 B.n706 B.n703 10.6151
R1936 B.n707 B.n706 10.6151
R1937 B.n708 B.n707 10.6151
R1938 B.n709 B.n708 10.6151
R1939 B.n711 B.n709 10.6151
R1940 B.n712 B.n711 10.6151
R1941 B.n713 B.n712 10.6151
R1942 B.n714 B.n713 10.6151
R1943 B.n716 B.n714 10.6151
R1944 B.n717 B.n716 10.6151
R1945 B.n718 B.n717 10.6151
R1946 B.n719 B.n718 10.6151
R1947 B.n721 B.n719 10.6151
R1948 B.n722 B.n721 10.6151
R1949 B.n723 B.n722 10.6151
R1950 B.n724 B.n723 10.6151
R1951 B.n726 B.n724 10.6151
R1952 B.n727 B.n726 10.6151
R1953 B.n728 B.n727 10.6151
R1954 B.n769 B.n1 10.6151
R1955 B.n769 B.n768 10.6151
R1956 B.n768 B.n767 10.6151
R1957 B.n767 B.n10 10.6151
R1958 B.n761 B.n10 10.6151
R1959 B.n761 B.n760 10.6151
R1960 B.n760 B.n759 10.6151
R1961 B.n759 B.n17 10.6151
R1962 B.n753 B.n17 10.6151
R1963 B.n753 B.n752 10.6151
R1964 B.n752 B.n751 10.6151
R1965 B.n751 B.n25 10.6151
R1966 B.n745 B.n25 10.6151
R1967 B.n745 B.n744 10.6151
R1968 B.n744 B.n743 10.6151
R1969 B.n743 B.n32 10.6151
R1970 B.n737 B.n32 10.6151
R1971 B.n737 B.n736 10.6151
R1972 B.n736 B.n735 10.6151
R1973 B.n735 B.n39 10.6151
R1974 B.n105 B.n104 10.6151
R1975 B.n108 B.n105 10.6151
R1976 B.n109 B.n108 10.6151
R1977 B.n112 B.n109 10.6151
R1978 B.n113 B.n112 10.6151
R1979 B.n116 B.n113 10.6151
R1980 B.n117 B.n116 10.6151
R1981 B.n120 B.n117 10.6151
R1982 B.n121 B.n120 10.6151
R1983 B.n124 B.n121 10.6151
R1984 B.n125 B.n124 10.6151
R1985 B.n128 B.n125 10.6151
R1986 B.n129 B.n128 10.6151
R1987 B.n132 B.n129 10.6151
R1988 B.n133 B.n132 10.6151
R1989 B.n136 B.n133 10.6151
R1990 B.n137 B.n136 10.6151
R1991 B.n140 B.n137 10.6151
R1992 B.n141 B.n140 10.6151
R1993 B.n144 B.n141 10.6151
R1994 B.n145 B.n144 10.6151
R1995 B.n148 B.n145 10.6151
R1996 B.n149 B.n148 10.6151
R1997 B.n152 B.n149 10.6151
R1998 B.n153 B.n152 10.6151
R1999 B.n156 B.n153 10.6151
R2000 B.n157 B.n156 10.6151
R2001 B.n160 B.n157 10.6151
R2002 B.n161 B.n160 10.6151
R2003 B.n164 B.n161 10.6151
R2004 B.n165 B.n164 10.6151
R2005 B.n168 B.n165 10.6151
R2006 B.n169 B.n168 10.6151
R2007 B.n172 B.n169 10.6151
R2008 B.n173 B.n172 10.6151
R2009 B.n176 B.n173 10.6151
R2010 B.n177 B.n176 10.6151
R2011 B.n180 B.n177 10.6151
R2012 B.n181 B.n180 10.6151
R2013 B.n184 B.n181 10.6151
R2014 B.n185 B.n184 10.6151
R2015 B.n188 B.n185 10.6151
R2016 B.n189 B.n188 10.6151
R2017 B.n192 B.n189 10.6151
R2018 B.n193 B.n192 10.6151
R2019 B.n196 B.n193 10.6151
R2020 B.n197 B.n196 10.6151
R2021 B.n200 B.n197 10.6151
R2022 B.n201 B.n200 10.6151
R2023 B.n205 B.n204 10.6151
R2024 B.n208 B.n205 10.6151
R2025 B.n209 B.n208 10.6151
R2026 B.n212 B.n209 10.6151
R2027 B.n213 B.n212 10.6151
R2028 B.n216 B.n213 10.6151
R2029 B.n217 B.n216 10.6151
R2030 B.n220 B.n217 10.6151
R2031 B.n225 B.n222 10.6151
R2032 B.n226 B.n225 10.6151
R2033 B.n229 B.n226 10.6151
R2034 B.n230 B.n229 10.6151
R2035 B.n233 B.n230 10.6151
R2036 B.n234 B.n233 10.6151
R2037 B.n237 B.n234 10.6151
R2038 B.n238 B.n237 10.6151
R2039 B.n241 B.n238 10.6151
R2040 B.n242 B.n241 10.6151
R2041 B.n245 B.n242 10.6151
R2042 B.n246 B.n245 10.6151
R2043 B.n249 B.n246 10.6151
R2044 B.n250 B.n249 10.6151
R2045 B.n253 B.n250 10.6151
R2046 B.n254 B.n253 10.6151
R2047 B.n257 B.n254 10.6151
R2048 B.n258 B.n257 10.6151
R2049 B.n261 B.n258 10.6151
R2050 B.n262 B.n261 10.6151
R2051 B.n265 B.n262 10.6151
R2052 B.n266 B.n265 10.6151
R2053 B.n269 B.n266 10.6151
R2054 B.n270 B.n269 10.6151
R2055 B.n273 B.n270 10.6151
R2056 B.n274 B.n273 10.6151
R2057 B.n277 B.n274 10.6151
R2058 B.n278 B.n277 10.6151
R2059 B.n281 B.n278 10.6151
R2060 B.n282 B.n281 10.6151
R2061 B.n285 B.n282 10.6151
R2062 B.n286 B.n285 10.6151
R2063 B.n289 B.n286 10.6151
R2064 B.n290 B.n289 10.6151
R2065 B.n293 B.n290 10.6151
R2066 B.n294 B.n293 10.6151
R2067 B.n297 B.n294 10.6151
R2068 B.n298 B.n297 10.6151
R2069 B.n301 B.n298 10.6151
R2070 B.n302 B.n301 10.6151
R2071 B.n305 B.n302 10.6151
R2072 B.n306 B.n305 10.6151
R2073 B.n309 B.n306 10.6151
R2074 B.n310 B.n309 10.6151
R2075 B.n313 B.n310 10.6151
R2076 B.n314 B.n313 10.6151
R2077 B.n317 B.n314 10.6151
R2078 B.n318 B.n317 10.6151
R2079 B.n729 B.n318 10.6151
R2080 B.n689 B.t2 8.82035
R2081 B.n12 B.t0 8.82035
R2082 B.n777 B.n0 8.11757
R2083 B.n777 B.n1 8.11757
R2084 B.n532 B.n531 6.5566
R2085 B.n515 B.n417 6.5566
R2086 B.n204 B.n102 6.5566
R2087 B.n221 B.n220 6.5566
R2088 B.n533 B.n532 4.05904
R2089 B.n512 B.n417 4.05904
R2090 B.n201 B.n102 4.05904
R2091 B.n222 B.n221 4.05904
R2092 B.n682 B.t4 3.30794
R2093 B.n763 B.t1 3.30794
R2094 B.n651 B.t7 2.20546
R2095 B.n741 B.t11 2.20546
R2096 VN.n1 VN.t5 514.826
R2097 VN.n7 VN.t4 514.826
R2098 VN.n2 VN.t0 491.339
R2099 VN.n4 VN.t1 491.339
R2100 VN.n8 VN.t3 491.339
R2101 VN.n10 VN.t2 491.339
R2102 VN.n5 VN.n4 161.3
R2103 VN.n11 VN.n10 161.3
R2104 VN.n9 VN.n6 161.3
R2105 VN.n3 VN.n0 161.3
R2106 VN.n7 VN.n6 44.8973
R2107 VN.n1 VN.n0 44.8973
R2108 VN VN.n11 44.1047
R2109 VN.n4 VN.n3 33.5944
R2110 VN.n10 VN.n9 33.5944
R2111 VN.n2 VN.n1 18.1882
R2112 VN.n8 VN.n7 18.1882
R2113 VN.n3 VN.n2 14.6066
R2114 VN.n9 VN.n8 14.6066
R2115 VN.n11 VN.n6 0.189894
R2116 VN.n5 VN.n0 0.189894
R2117 VN VN.n5 0.0516364
R2118 VDD2.n159 VDD2.n83 289.615
R2119 VDD2.n76 VDD2.n0 289.615
R2120 VDD2.n160 VDD2.n159 185
R2121 VDD2.n158 VDD2.n157 185
R2122 VDD2.n156 VDD2.n86 185
R2123 VDD2.n90 VDD2.n87 185
R2124 VDD2.n151 VDD2.n150 185
R2125 VDD2.n149 VDD2.n148 185
R2126 VDD2.n92 VDD2.n91 185
R2127 VDD2.n143 VDD2.n142 185
R2128 VDD2.n141 VDD2.n140 185
R2129 VDD2.n96 VDD2.n95 185
R2130 VDD2.n135 VDD2.n134 185
R2131 VDD2.n133 VDD2.n132 185
R2132 VDD2.n100 VDD2.n99 185
R2133 VDD2.n127 VDD2.n126 185
R2134 VDD2.n125 VDD2.n124 185
R2135 VDD2.n104 VDD2.n103 185
R2136 VDD2.n119 VDD2.n118 185
R2137 VDD2.n117 VDD2.n116 185
R2138 VDD2.n108 VDD2.n107 185
R2139 VDD2.n111 VDD2.n110 185
R2140 VDD2.n27 VDD2.n26 185
R2141 VDD2.n24 VDD2.n23 185
R2142 VDD2.n33 VDD2.n32 185
R2143 VDD2.n35 VDD2.n34 185
R2144 VDD2.n20 VDD2.n19 185
R2145 VDD2.n41 VDD2.n40 185
R2146 VDD2.n43 VDD2.n42 185
R2147 VDD2.n16 VDD2.n15 185
R2148 VDD2.n49 VDD2.n48 185
R2149 VDD2.n51 VDD2.n50 185
R2150 VDD2.n12 VDD2.n11 185
R2151 VDD2.n57 VDD2.n56 185
R2152 VDD2.n59 VDD2.n58 185
R2153 VDD2.n8 VDD2.n7 185
R2154 VDD2.n65 VDD2.n64 185
R2155 VDD2.n68 VDD2.n67 185
R2156 VDD2.n66 VDD2.n4 185
R2157 VDD2.n73 VDD2.n3 185
R2158 VDD2.n75 VDD2.n74 185
R2159 VDD2.n77 VDD2.n76 185
R2160 VDD2.t3 VDD2.n109 147.659
R2161 VDD2.t0 VDD2.n25 147.659
R2162 VDD2.n159 VDD2.n158 104.615
R2163 VDD2.n158 VDD2.n86 104.615
R2164 VDD2.n90 VDD2.n86 104.615
R2165 VDD2.n150 VDD2.n90 104.615
R2166 VDD2.n150 VDD2.n149 104.615
R2167 VDD2.n149 VDD2.n91 104.615
R2168 VDD2.n142 VDD2.n91 104.615
R2169 VDD2.n142 VDD2.n141 104.615
R2170 VDD2.n141 VDD2.n95 104.615
R2171 VDD2.n134 VDD2.n95 104.615
R2172 VDD2.n134 VDD2.n133 104.615
R2173 VDD2.n133 VDD2.n99 104.615
R2174 VDD2.n126 VDD2.n99 104.615
R2175 VDD2.n126 VDD2.n125 104.615
R2176 VDD2.n125 VDD2.n103 104.615
R2177 VDD2.n118 VDD2.n103 104.615
R2178 VDD2.n118 VDD2.n117 104.615
R2179 VDD2.n117 VDD2.n107 104.615
R2180 VDD2.n110 VDD2.n107 104.615
R2181 VDD2.n26 VDD2.n23 104.615
R2182 VDD2.n33 VDD2.n23 104.615
R2183 VDD2.n34 VDD2.n33 104.615
R2184 VDD2.n34 VDD2.n19 104.615
R2185 VDD2.n41 VDD2.n19 104.615
R2186 VDD2.n42 VDD2.n41 104.615
R2187 VDD2.n42 VDD2.n15 104.615
R2188 VDD2.n49 VDD2.n15 104.615
R2189 VDD2.n50 VDD2.n49 104.615
R2190 VDD2.n50 VDD2.n11 104.615
R2191 VDD2.n57 VDD2.n11 104.615
R2192 VDD2.n58 VDD2.n57 104.615
R2193 VDD2.n58 VDD2.n7 104.615
R2194 VDD2.n65 VDD2.n7 104.615
R2195 VDD2.n67 VDD2.n65 104.615
R2196 VDD2.n67 VDD2.n66 104.615
R2197 VDD2.n66 VDD2.n3 104.615
R2198 VDD2.n75 VDD2.n3 104.615
R2199 VDD2.n76 VDD2.n75 104.615
R2200 VDD2.n82 VDD2.n81 61.8849
R2201 VDD2 VDD2.n165 61.882
R2202 VDD2.n110 VDD2.t3 52.3082
R2203 VDD2.n26 VDD2.t0 52.3082
R2204 VDD2.n82 VDD2.n80 50.3152
R2205 VDD2.n164 VDD2.n163 49.6399
R2206 VDD2.n164 VDD2.n82 39.5364
R2207 VDD2.n111 VDD2.n109 15.6677
R2208 VDD2.n27 VDD2.n25 15.6677
R2209 VDD2.n157 VDD2.n156 13.1884
R2210 VDD2.n74 VDD2.n73 13.1884
R2211 VDD2.n160 VDD2.n85 12.8005
R2212 VDD2.n155 VDD2.n87 12.8005
R2213 VDD2.n112 VDD2.n108 12.8005
R2214 VDD2.n28 VDD2.n24 12.8005
R2215 VDD2.n72 VDD2.n4 12.8005
R2216 VDD2.n77 VDD2.n2 12.8005
R2217 VDD2.n161 VDD2.n83 12.0247
R2218 VDD2.n152 VDD2.n151 12.0247
R2219 VDD2.n116 VDD2.n115 12.0247
R2220 VDD2.n32 VDD2.n31 12.0247
R2221 VDD2.n69 VDD2.n68 12.0247
R2222 VDD2.n78 VDD2.n0 12.0247
R2223 VDD2.n148 VDD2.n89 11.249
R2224 VDD2.n119 VDD2.n106 11.249
R2225 VDD2.n35 VDD2.n22 11.249
R2226 VDD2.n64 VDD2.n6 11.249
R2227 VDD2.n147 VDD2.n92 10.4732
R2228 VDD2.n120 VDD2.n104 10.4732
R2229 VDD2.n36 VDD2.n20 10.4732
R2230 VDD2.n63 VDD2.n8 10.4732
R2231 VDD2.n144 VDD2.n143 9.69747
R2232 VDD2.n124 VDD2.n123 9.69747
R2233 VDD2.n40 VDD2.n39 9.69747
R2234 VDD2.n60 VDD2.n59 9.69747
R2235 VDD2.n163 VDD2.n162 9.45567
R2236 VDD2.n80 VDD2.n79 9.45567
R2237 VDD2.n137 VDD2.n136 9.3005
R2238 VDD2.n139 VDD2.n138 9.3005
R2239 VDD2.n94 VDD2.n93 9.3005
R2240 VDD2.n145 VDD2.n144 9.3005
R2241 VDD2.n147 VDD2.n146 9.3005
R2242 VDD2.n89 VDD2.n88 9.3005
R2243 VDD2.n153 VDD2.n152 9.3005
R2244 VDD2.n155 VDD2.n154 9.3005
R2245 VDD2.n162 VDD2.n161 9.3005
R2246 VDD2.n85 VDD2.n84 9.3005
R2247 VDD2.n98 VDD2.n97 9.3005
R2248 VDD2.n131 VDD2.n130 9.3005
R2249 VDD2.n129 VDD2.n128 9.3005
R2250 VDD2.n102 VDD2.n101 9.3005
R2251 VDD2.n123 VDD2.n122 9.3005
R2252 VDD2.n121 VDD2.n120 9.3005
R2253 VDD2.n106 VDD2.n105 9.3005
R2254 VDD2.n115 VDD2.n114 9.3005
R2255 VDD2.n113 VDD2.n112 9.3005
R2256 VDD2.n79 VDD2.n78 9.3005
R2257 VDD2.n2 VDD2.n1 9.3005
R2258 VDD2.n47 VDD2.n46 9.3005
R2259 VDD2.n45 VDD2.n44 9.3005
R2260 VDD2.n18 VDD2.n17 9.3005
R2261 VDD2.n39 VDD2.n38 9.3005
R2262 VDD2.n37 VDD2.n36 9.3005
R2263 VDD2.n22 VDD2.n21 9.3005
R2264 VDD2.n31 VDD2.n30 9.3005
R2265 VDD2.n29 VDD2.n28 9.3005
R2266 VDD2.n14 VDD2.n13 9.3005
R2267 VDD2.n53 VDD2.n52 9.3005
R2268 VDD2.n55 VDD2.n54 9.3005
R2269 VDD2.n10 VDD2.n9 9.3005
R2270 VDD2.n61 VDD2.n60 9.3005
R2271 VDD2.n63 VDD2.n62 9.3005
R2272 VDD2.n6 VDD2.n5 9.3005
R2273 VDD2.n70 VDD2.n69 9.3005
R2274 VDD2.n72 VDD2.n71 9.3005
R2275 VDD2.n140 VDD2.n94 8.92171
R2276 VDD2.n127 VDD2.n102 8.92171
R2277 VDD2.n43 VDD2.n18 8.92171
R2278 VDD2.n56 VDD2.n10 8.92171
R2279 VDD2.n139 VDD2.n96 8.14595
R2280 VDD2.n128 VDD2.n100 8.14595
R2281 VDD2.n44 VDD2.n16 8.14595
R2282 VDD2.n55 VDD2.n12 8.14595
R2283 VDD2.n136 VDD2.n135 7.3702
R2284 VDD2.n132 VDD2.n131 7.3702
R2285 VDD2.n48 VDD2.n47 7.3702
R2286 VDD2.n52 VDD2.n51 7.3702
R2287 VDD2.n135 VDD2.n98 6.59444
R2288 VDD2.n132 VDD2.n98 6.59444
R2289 VDD2.n48 VDD2.n14 6.59444
R2290 VDD2.n51 VDD2.n14 6.59444
R2291 VDD2.n136 VDD2.n96 5.81868
R2292 VDD2.n131 VDD2.n100 5.81868
R2293 VDD2.n47 VDD2.n16 5.81868
R2294 VDD2.n52 VDD2.n12 5.81868
R2295 VDD2.n140 VDD2.n139 5.04292
R2296 VDD2.n128 VDD2.n127 5.04292
R2297 VDD2.n44 VDD2.n43 5.04292
R2298 VDD2.n56 VDD2.n55 5.04292
R2299 VDD2.n113 VDD2.n109 4.38563
R2300 VDD2.n29 VDD2.n25 4.38563
R2301 VDD2.n143 VDD2.n94 4.26717
R2302 VDD2.n124 VDD2.n102 4.26717
R2303 VDD2.n40 VDD2.n18 4.26717
R2304 VDD2.n59 VDD2.n10 4.26717
R2305 VDD2.n144 VDD2.n92 3.49141
R2306 VDD2.n123 VDD2.n104 3.49141
R2307 VDD2.n39 VDD2.n20 3.49141
R2308 VDD2.n60 VDD2.n8 3.49141
R2309 VDD2.n148 VDD2.n147 2.71565
R2310 VDD2.n120 VDD2.n119 2.71565
R2311 VDD2.n36 VDD2.n35 2.71565
R2312 VDD2.n64 VDD2.n63 2.71565
R2313 VDD2.n163 VDD2.n83 1.93989
R2314 VDD2.n151 VDD2.n89 1.93989
R2315 VDD2.n116 VDD2.n106 1.93989
R2316 VDD2.n32 VDD2.n22 1.93989
R2317 VDD2.n68 VDD2.n6 1.93989
R2318 VDD2.n80 VDD2.n0 1.93989
R2319 VDD2.n165 VDD2.t2 1.34927
R2320 VDD2.n165 VDD2.t1 1.34927
R2321 VDD2.n81 VDD2.t5 1.34927
R2322 VDD2.n81 VDD2.t4 1.34927
R2323 VDD2.n161 VDD2.n160 1.16414
R2324 VDD2.n152 VDD2.n87 1.16414
R2325 VDD2.n115 VDD2.n108 1.16414
R2326 VDD2.n31 VDD2.n24 1.16414
R2327 VDD2.n69 VDD2.n4 1.16414
R2328 VDD2.n78 VDD2.n77 1.16414
R2329 VDD2 VDD2.n164 0.789293
R2330 VDD2.n157 VDD2.n85 0.388379
R2331 VDD2.n156 VDD2.n155 0.388379
R2332 VDD2.n112 VDD2.n111 0.388379
R2333 VDD2.n28 VDD2.n27 0.388379
R2334 VDD2.n73 VDD2.n72 0.388379
R2335 VDD2.n74 VDD2.n2 0.388379
R2336 VDD2.n162 VDD2.n84 0.155672
R2337 VDD2.n154 VDD2.n84 0.155672
R2338 VDD2.n154 VDD2.n153 0.155672
R2339 VDD2.n153 VDD2.n88 0.155672
R2340 VDD2.n146 VDD2.n88 0.155672
R2341 VDD2.n146 VDD2.n145 0.155672
R2342 VDD2.n145 VDD2.n93 0.155672
R2343 VDD2.n138 VDD2.n93 0.155672
R2344 VDD2.n138 VDD2.n137 0.155672
R2345 VDD2.n137 VDD2.n97 0.155672
R2346 VDD2.n130 VDD2.n97 0.155672
R2347 VDD2.n130 VDD2.n129 0.155672
R2348 VDD2.n129 VDD2.n101 0.155672
R2349 VDD2.n122 VDD2.n101 0.155672
R2350 VDD2.n122 VDD2.n121 0.155672
R2351 VDD2.n121 VDD2.n105 0.155672
R2352 VDD2.n114 VDD2.n105 0.155672
R2353 VDD2.n114 VDD2.n113 0.155672
R2354 VDD2.n30 VDD2.n29 0.155672
R2355 VDD2.n30 VDD2.n21 0.155672
R2356 VDD2.n37 VDD2.n21 0.155672
R2357 VDD2.n38 VDD2.n37 0.155672
R2358 VDD2.n38 VDD2.n17 0.155672
R2359 VDD2.n45 VDD2.n17 0.155672
R2360 VDD2.n46 VDD2.n45 0.155672
R2361 VDD2.n46 VDD2.n13 0.155672
R2362 VDD2.n53 VDD2.n13 0.155672
R2363 VDD2.n54 VDD2.n53 0.155672
R2364 VDD2.n54 VDD2.n9 0.155672
R2365 VDD2.n61 VDD2.n9 0.155672
R2366 VDD2.n62 VDD2.n61 0.155672
R2367 VDD2.n62 VDD2.n5 0.155672
R2368 VDD2.n70 VDD2.n5 0.155672
R2369 VDD2.n71 VDD2.n70 0.155672
R2370 VDD2.n71 VDD2.n1 0.155672
R2371 VDD2.n79 VDD2.n1 0.155672
C0 VDD2 VTAIL 11.180201f
C1 VP VDD2 0.306657f
C2 VDD2 VDD1 0.746866f
C3 VP VTAIL 5.20371f
C4 VTAIL VDD1 11.146501f
C5 VP VDD1 5.73343f
C6 VN VDD2 5.58054f
C7 VN VTAIL 5.18903f
C8 VP VN 5.66769f
C9 VN VDD1 0.148484f
C10 VDD2 B 5.047147f
C11 VDD1 B 5.074131f
C12 VTAIL B 7.473146f
C13 VN B 8.292871f
C14 VP B 6.24226f
C15 VDD2.n0 B 0.02982f
C16 VDD2.n1 B 0.022981f
C17 VDD2.n2 B 0.012349f
C18 VDD2.n3 B 0.029188f
C19 VDD2.n4 B 0.013075f
C20 VDD2.n5 B 0.022981f
C21 VDD2.n6 B 0.012349f
C22 VDD2.n7 B 0.029188f
C23 VDD2.n8 B 0.013075f
C24 VDD2.n9 B 0.022981f
C25 VDD2.n10 B 0.012349f
C26 VDD2.n11 B 0.029188f
C27 VDD2.n12 B 0.013075f
C28 VDD2.n13 B 0.022981f
C29 VDD2.n14 B 0.012349f
C30 VDD2.n15 B 0.029188f
C31 VDD2.n16 B 0.013075f
C32 VDD2.n17 B 0.022981f
C33 VDD2.n18 B 0.012349f
C34 VDD2.n19 B 0.029188f
C35 VDD2.n20 B 0.013075f
C36 VDD2.n21 B 0.022981f
C37 VDD2.n22 B 0.012349f
C38 VDD2.n23 B 0.029188f
C39 VDD2.n24 B 0.013075f
C40 VDD2.n25 B 0.14804f
C41 VDD2.t0 B 0.048102f
C42 VDD2.n26 B 0.021891f
C43 VDD2.n27 B 0.017242f
C44 VDD2.n28 B 0.012349f
C45 VDD2.n29 B 1.46145f
C46 VDD2.n30 B 0.022981f
C47 VDD2.n31 B 0.012349f
C48 VDD2.n32 B 0.013075f
C49 VDD2.n33 B 0.029188f
C50 VDD2.n34 B 0.029188f
C51 VDD2.n35 B 0.013075f
C52 VDD2.n36 B 0.012349f
C53 VDD2.n37 B 0.022981f
C54 VDD2.n38 B 0.022981f
C55 VDD2.n39 B 0.012349f
C56 VDD2.n40 B 0.013075f
C57 VDD2.n41 B 0.029188f
C58 VDD2.n42 B 0.029188f
C59 VDD2.n43 B 0.013075f
C60 VDD2.n44 B 0.012349f
C61 VDD2.n45 B 0.022981f
C62 VDD2.n46 B 0.022981f
C63 VDD2.n47 B 0.012349f
C64 VDD2.n48 B 0.013075f
C65 VDD2.n49 B 0.029188f
C66 VDD2.n50 B 0.029188f
C67 VDD2.n51 B 0.013075f
C68 VDD2.n52 B 0.012349f
C69 VDD2.n53 B 0.022981f
C70 VDD2.n54 B 0.022981f
C71 VDD2.n55 B 0.012349f
C72 VDD2.n56 B 0.013075f
C73 VDD2.n57 B 0.029188f
C74 VDD2.n58 B 0.029188f
C75 VDD2.n59 B 0.013075f
C76 VDD2.n60 B 0.012349f
C77 VDD2.n61 B 0.022981f
C78 VDD2.n62 B 0.022981f
C79 VDD2.n63 B 0.012349f
C80 VDD2.n64 B 0.013075f
C81 VDD2.n65 B 0.029188f
C82 VDD2.n66 B 0.029188f
C83 VDD2.n67 B 0.029188f
C84 VDD2.n68 B 0.013075f
C85 VDD2.n69 B 0.012349f
C86 VDD2.n70 B 0.022981f
C87 VDD2.n71 B 0.022981f
C88 VDD2.n72 B 0.012349f
C89 VDD2.n73 B 0.012712f
C90 VDD2.n74 B 0.012712f
C91 VDD2.n75 B 0.029188f
C92 VDD2.n76 B 0.0588f
C93 VDD2.n77 B 0.013075f
C94 VDD2.n78 B 0.012349f
C95 VDD2.n79 B 0.054374f
C96 VDD2.n80 B 0.049631f
C97 VDD2.t5 B 0.266588f
C98 VDD2.t4 B 0.266588f
C99 VDD2.n81 B 2.4089f
C100 VDD2.n82 B 1.89255f
C101 VDD2.n83 B 0.02982f
C102 VDD2.n84 B 0.022981f
C103 VDD2.n85 B 0.012349f
C104 VDD2.n86 B 0.029188f
C105 VDD2.n87 B 0.013075f
C106 VDD2.n88 B 0.022981f
C107 VDD2.n89 B 0.012349f
C108 VDD2.n90 B 0.029188f
C109 VDD2.n91 B 0.029188f
C110 VDD2.n92 B 0.013075f
C111 VDD2.n93 B 0.022981f
C112 VDD2.n94 B 0.012349f
C113 VDD2.n95 B 0.029188f
C114 VDD2.n96 B 0.013075f
C115 VDD2.n97 B 0.022981f
C116 VDD2.n98 B 0.012349f
C117 VDD2.n99 B 0.029188f
C118 VDD2.n100 B 0.013075f
C119 VDD2.n101 B 0.022981f
C120 VDD2.n102 B 0.012349f
C121 VDD2.n103 B 0.029188f
C122 VDD2.n104 B 0.013075f
C123 VDD2.n105 B 0.022981f
C124 VDD2.n106 B 0.012349f
C125 VDD2.n107 B 0.029188f
C126 VDD2.n108 B 0.013075f
C127 VDD2.n109 B 0.14804f
C128 VDD2.t3 B 0.048102f
C129 VDD2.n110 B 0.021891f
C130 VDD2.n111 B 0.017242f
C131 VDD2.n112 B 0.012349f
C132 VDD2.n113 B 1.46145f
C133 VDD2.n114 B 0.022981f
C134 VDD2.n115 B 0.012349f
C135 VDD2.n116 B 0.013075f
C136 VDD2.n117 B 0.029188f
C137 VDD2.n118 B 0.029188f
C138 VDD2.n119 B 0.013075f
C139 VDD2.n120 B 0.012349f
C140 VDD2.n121 B 0.022981f
C141 VDD2.n122 B 0.022981f
C142 VDD2.n123 B 0.012349f
C143 VDD2.n124 B 0.013075f
C144 VDD2.n125 B 0.029188f
C145 VDD2.n126 B 0.029188f
C146 VDD2.n127 B 0.013075f
C147 VDD2.n128 B 0.012349f
C148 VDD2.n129 B 0.022981f
C149 VDD2.n130 B 0.022981f
C150 VDD2.n131 B 0.012349f
C151 VDD2.n132 B 0.013075f
C152 VDD2.n133 B 0.029188f
C153 VDD2.n134 B 0.029188f
C154 VDD2.n135 B 0.013075f
C155 VDD2.n136 B 0.012349f
C156 VDD2.n137 B 0.022981f
C157 VDD2.n138 B 0.022981f
C158 VDD2.n139 B 0.012349f
C159 VDD2.n140 B 0.013075f
C160 VDD2.n141 B 0.029188f
C161 VDD2.n142 B 0.029188f
C162 VDD2.n143 B 0.013075f
C163 VDD2.n144 B 0.012349f
C164 VDD2.n145 B 0.022981f
C165 VDD2.n146 B 0.022981f
C166 VDD2.n147 B 0.012349f
C167 VDD2.n148 B 0.013075f
C168 VDD2.n149 B 0.029188f
C169 VDD2.n150 B 0.029188f
C170 VDD2.n151 B 0.013075f
C171 VDD2.n152 B 0.012349f
C172 VDD2.n153 B 0.022981f
C173 VDD2.n154 B 0.022981f
C174 VDD2.n155 B 0.012349f
C175 VDD2.n156 B 0.012712f
C176 VDD2.n157 B 0.012712f
C177 VDD2.n158 B 0.029188f
C178 VDD2.n159 B 0.0588f
C179 VDD2.n160 B 0.013075f
C180 VDD2.n161 B 0.012349f
C181 VDD2.n162 B 0.054374f
C182 VDD2.n163 B 0.048346f
C183 VDD2.n164 B 2.09568f
C184 VDD2.t2 B 0.266588f
C185 VDD2.t1 B 0.266588f
C186 VDD2.n165 B 2.40888f
C187 VN.n0 B 0.189041f
C188 VN.t5 B 1.48533f
C189 VN.n1 B 0.541832f
C190 VN.t0 B 1.45962f
C191 VN.n2 B 0.565984f
C192 VN.n3 B 0.009922f
C193 VN.t1 B 1.45962f
C194 VN.n4 B 0.561733f
C195 VN.n5 B 0.033884f
C196 VN.n6 B 0.189041f
C197 VN.t4 B 1.48533f
C198 VN.n7 B 0.541832f
C199 VN.t3 B 1.45962f
C200 VN.n8 B 0.565984f
C201 VN.n9 B 0.009922f
C202 VN.t2 B 1.45962f
C203 VN.n10 B 0.561733f
C204 VN.n11 B 1.95679f
C205 VTAIL.t0 B 0.27377f
C206 VTAIL.t1 B 0.27377f
C207 VTAIL.n0 B 2.4034f
C208 VTAIL.n1 B 0.325247f
C209 VTAIL.n2 B 0.030624f
C210 VTAIL.n3 B 0.0236f
C211 VTAIL.n4 B 0.012681f
C212 VTAIL.n5 B 0.029974f
C213 VTAIL.n6 B 0.013427f
C214 VTAIL.n7 B 0.0236f
C215 VTAIL.n8 B 0.012681f
C216 VTAIL.n9 B 0.029974f
C217 VTAIL.n10 B 0.013427f
C218 VTAIL.n11 B 0.0236f
C219 VTAIL.n12 B 0.012681f
C220 VTAIL.n13 B 0.029974f
C221 VTAIL.n14 B 0.013427f
C222 VTAIL.n15 B 0.0236f
C223 VTAIL.n16 B 0.012681f
C224 VTAIL.n17 B 0.029974f
C225 VTAIL.n18 B 0.013427f
C226 VTAIL.n19 B 0.0236f
C227 VTAIL.n20 B 0.012681f
C228 VTAIL.n21 B 0.029974f
C229 VTAIL.n22 B 0.013427f
C230 VTAIL.n23 B 0.0236f
C231 VTAIL.n24 B 0.012681f
C232 VTAIL.n25 B 0.029974f
C233 VTAIL.n26 B 0.013427f
C234 VTAIL.n27 B 0.152028f
C235 VTAIL.t9 B 0.049398f
C236 VTAIL.n28 B 0.022481f
C237 VTAIL.n29 B 0.017707f
C238 VTAIL.n30 B 0.012681f
C239 VTAIL.n31 B 1.50082f
C240 VTAIL.n32 B 0.0236f
C241 VTAIL.n33 B 0.012681f
C242 VTAIL.n34 B 0.013427f
C243 VTAIL.n35 B 0.029974f
C244 VTAIL.n36 B 0.029974f
C245 VTAIL.n37 B 0.013427f
C246 VTAIL.n38 B 0.012681f
C247 VTAIL.n39 B 0.0236f
C248 VTAIL.n40 B 0.0236f
C249 VTAIL.n41 B 0.012681f
C250 VTAIL.n42 B 0.013427f
C251 VTAIL.n43 B 0.029974f
C252 VTAIL.n44 B 0.029974f
C253 VTAIL.n45 B 0.013427f
C254 VTAIL.n46 B 0.012681f
C255 VTAIL.n47 B 0.0236f
C256 VTAIL.n48 B 0.0236f
C257 VTAIL.n49 B 0.012681f
C258 VTAIL.n50 B 0.013427f
C259 VTAIL.n51 B 0.029974f
C260 VTAIL.n52 B 0.029974f
C261 VTAIL.n53 B 0.013427f
C262 VTAIL.n54 B 0.012681f
C263 VTAIL.n55 B 0.0236f
C264 VTAIL.n56 B 0.0236f
C265 VTAIL.n57 B 0.012681f
C266 VTAIL.n58 B 0.013427f
C267 VTAIL.n59 B 0.029974f
C268 VTAIL.n60 B 0.029974f
C269 VTAIL.n61 B 0.013427f
C270 VTAIL.n62 B 0.012681f
C271 VTAIL.n63 B 0.0236f
C272 VTAIL.n64 B 0.0236f
C273 VTAIL.n65 B 0.012681f
C274 VTAIL.n66 B 0.013427f
C275 VTAIL.n67 B 0.029974f
C276 VTAIL.n68 B 0.029974f
C277 VTAIL.n69 B 0.029974f
C278 VTAIL.n70 B 0.013427f
C279 VTAIL.n71 B 0.012681f
C280 VTAIL.n72 B 0.0236f
C281 VTAIL.n73 B 0.0236f
C282 VTAIL.n74 B 0.012681f
C283 VTAIL.n75 B 0.013054f
C284 VTAIL.n76 B 0.013054f
C285 VTAIL.n77 B 0.029974f
C286 VTAIL.n78 B 0.060384f
C287 VTAIL.n79 B 0.013427f
C288 VTAIL.n80 B 0.012681f
C289 VTAIL.n81 B 0.055839f
C290 VTAIL.n82 B 0.033363f
C291 VTAIL.n83 B 0.167726f
C292 VTAIL.t10 B 0.27377f
C293 VTAIL.t11 B 0.27377f
C294 VTAIL.n84 B 2.4034f
C295 VTAIL.n85 B 1.73468f
C296 VTAIL.t5 B 0.27377f
C297 VTAIL.t4 B 0.27377f
C298 VTAIL.n86 B 2.40341f
C299 VTAIL.n87 B 1.73467f
C300 VTAIL.n88 B 0.030624f
C301 VTAIL.n89 B 0.0236f
C302 VTAIL.n90 B 0.012681f
C303 VTAIL.n91 B 0.029974f
C304 VTAIL.n92 B 0.013427f
C305 VTAIL.n93 B 0.0236f
C306 VTAIL.n94 B 0.012681f
C307 VTAIL.n95 B 0.029974f
C308 VTAIL.n96 B 0.029974f
C309 VTAIL.n97 B 0.013427f
C310 VTAIL.n98 B 0.0236f
C311 VTAIL.n99 B 0.012681f
C312 VTAIL.n100 B 0.029974f
C313 VTAIL.n101 B 0.013427f
C314 VTAIL.n102 B 0.0236f
C315 VTAIL.n103 B 0.012681f
C316 VTAIL.n104 B 0.029974f
C317 VTAIL.n105 B 0.013427f
C318 VTAIL.n106 B 0.0236f
C319 VTAIL.n107 B 0.012681f
C320 VTAIL.n108 B 0.029974f
C321 VTAIL.n109 B 0.013427f
C322 VTAIL.n110 B 0.0236f
C323 VTAIL.n111 B 0.012681f
C324 VTAIL.n112 B 0.029974f
C325 VTAIL.n113 B 0.013427f
C326 VTAIL.n114 B 0.152028f
C327 VTAIL.t2 B 0.049398f
C328 VTAIL.n115 B 0.022481f
C329 VTAIL.n116 B 0.017707f
C330 VTAIL.n117 B 0.012681f
C331 VTAIL.n118 B 1.50082f
C332 VTAIL.n119 B 0.0236f
C333 VTAIL.n120 B 0.012681f
C334 VTAIL.n121 B 0.013427f
C335 VTAIL.n122 B 0.029974f
C336 VTAIL.n123 B 0.029974f
C337 VTAIL.n124 B 0.013427f
C338 VTAIL.n125 B 0.012681f
C339 VTAIL.n126 B 0.0236f
C340 VTAIL.n127 B 0.0236f
C341 VTAIL.n128 B 0.012681f
C342 VTAIL.n129 B 0.013427f
C343 VTAIL.n130 B 0.029974f
C344 VTAIL.n131 B 0.029974f
C345 VTAIL.n132 B 0.013427f
C346 VTAIL.n133 B 0.012681f
C347 VTAIL.n134 B 0.0236f
C348 VTAIL.n135 B 0.0236f
C349 VTAIL.n136 B 0.012681f
C350 VTAIL.n137 B 0.013427f
C351 VTAIL.n138 B 0.029974f
C352 VTAIL.n139 B 0.029974f
C353 VTAIL.n140 B 0.013427f
C354 VTAIL.n141 B 0.012681f
C355 VTAIL.n142 B 0.0236f
C356 VTAIL.n143 B 0.0236f
C357 VTAIL.n144 B 0.012681f
C358 VTAIL.n145 B 0.013427f
C359 VTAIL.n146 B 0.029974f
C360 VTAIL.n147 B 0.029974f
C361 VTAIL.n148 B 0.013427f
C362 VTAIL.n149 B 0.012681f
C363 VTAIL.n150 B 0.0236f
C364 VTAIL.n151 B 0.0236f
C365 VTAIL.n152 B 0.012681f
C366 VTAIL.n153 B 0.013427f
C367 VTAIL.n154 B 0.029974f
C368 VTAIL.n155 B 0.029974f
C369 VTAIL.n156 B 0.013427f
C370 VTAIL.n157 B 0.012681f
C371 VTAIL.n158 B 0.0236f
C372 VTAIL.n159 B 0.0236f
C373 VTAIL.n160 B 0.012681f
C374 VTAIL.n161 B 0.013054f
C375 VTAIL.n162 B 0.013054f
C376 VTAIL.n163 B 0.029974f
C377 VTAIL.n164 B 0.060384f
C378 VTAIL.n165 B 0.013427f
C379 VTAIL.n166 B 0.012681f
C380 VTAIL.n167 B 0.055839f
C381 VTAIL.n168 B 0.033363f
C382 VTAIL.n169 B 0.167726f
C383 VTAIL.t6 B 0.27377f
C384 VTAIL.t7 B 0.27377f
C385 VTAIL.n170 B 2.40341f
C386 VTAIL.n171 B 0.376367f
C387 VTAIL.n172 B 0.030624f
C388 VTAIL.n173 B 0.0236f
C389 VTAIL.n174 B 0.012681f
C390 VTAIL.n175 B 0.029974f
C391 VTAIL.n176 B 0.013427f
C392 VTAIL.n177 B 0.0236f
C393 VTAIL.n178 B 0.012681f
C394 VTAIL.n179 B 0.029974f
C395 VTAIL.n180 B 0.029974f
C396 VTAIL.n181 B 0.013427f
C397 VTAIL.n182 B 0.0236f
C398 VTAIL.n183 B 0.012681f
C399 VTAIL.n184 B 0.029974f
C400 VTAIL.n185 B 0.013427f
C401 VTAIL.n186 B 0.0236f
C402 VTAIL.n187 B 0.012681f
C403 VTAIL.n188 B 0.029974f
C404 VTAIL.n189 B 0.013427f
C405 VTAIL.n190 B 0.0236f
C406 VTAIL.n191 B 0.012681f
C407 VTAIL.n192 B 0.029974f
C408 VTAIL.n193 B 0.013427f
C409 VTAIL.n194 B 0.0236f
C410 VTAIL.n195 B 0.012681f
C411 VTAIL.n196 B 0.029974f
C412 VTAIL.n197 B 0.013427f
C413 VTAIL.n198 B 0.152028f
C414 VTAIL.t8 B 0.049398f
C415 VTAIL.n199 B 0.022481f
C416 VTAIL.n200 B 0.017707f
C417 VTAIL.n201 B 0.012681f
C418 VTAIL.n202 B 1.50082f
C419 VTAIL.n203 B 0.0236f
C420 VTAIL.n204 B 0.012681f
C421 VTAIL.n205 B 0.013427f
C422 VTAIL.n206 B 0.029974f
C423 VTAIL.n207 B 0.029974f
C424 VTAIL.n208 B 0.013427f
C425 VTAIL.n209 B 0.012681f
C426 VTAIL.n210 B 0.0236f
C427 VTAIL.n211 B 0.0236f
C428 VTAIL.n212 B 0.012681f
C429 VTAIL.n213 B 0.013427f
C430 VTAIL.n214 B 0.029974f
C431 VTAIL.n215 B 0.029974f
C432 VTAIL.n216 B 0.013427f
C433 VTAIL.n217 B 0.012681f
C434 VTAIL.n218 B 0.0236f
C435 VTAIL.n219 B 0.0236f
C436 VTAIL.n220 B 0.012681f
C437 VTAIL.n221 B 0.013427f
C438 VTAIL.n222 B 0.029974f
C439 VTAIL.n223 B 0.029974f
C440 VTAIL.n224 B 0.013427f
C441 VTAIL.n225 B 0.012681f
C442 VTAIL.n226 B 0.0236f
C443 VTAIL.n227 B 0.0236f
C444 VTAIL.n228 B 0.012681f
C445 VTAIL.n229 B 0.013427f
C446 VTAIL.n230 B 0.029974f
C447 VTAIL.n231 B 0.029974f
C448 VTAIL.n232 B 0.013427f
C449 VTAIL.n233 B 0.012681f
C450 VTAIL.n234 B 0.0236f
C451 VTAIL.n235 B 0.0236f
C452 VTAIL.n236 B 0.012681f
C453 VTAIL.n237 B 0.013427f
C454 VTAIL.n238 B 0.029974f
C455 VTAIL.n239 B 0.029974f
C456 VTAIL.n240 B 0.013427f
C457 VTAIL.n241 B 0.012681f
C458 VTAIL.n242 B 0.0236f
C459 VTAIL.n243 B 0.0236f
C460 VTAIL.n244 B 0.012681f
C461 VTAIL.n245 B 0.013054f
C462 VTAIL.n246 B 0.013054f
C463 VTAIL.n247 B 0.029974f
C464 VTAIL.n248 B 0.060384f
C465 VTAIL.n249 B 0.013427f
C466 VTAIL.n250 B 0.012681f
C467 VTAIL.n251 B 0.055839f
C468 VTAIL.n252 B 0.033363f
C469 VTAIL.n253 B 1.45195f
C470 VTAIL.n254 B 0.030624f
C471 VTAIL.n255 B 0.0236f
C472 VTAIL.n256 B 0.012681f
C473 VTAIL.n257 B 0.029974f
C474 VTAIL.n258 B 0.013427f
C475 VTAIL.n259 B 0.0236f
C476 VTAIL.n260 B 0.012681f
C477 VTAIL.n261 B 0.029974f
C478 VTAIL.n262 B 0.013427f
C479 VTAIL.n263 B 0.0236f
C480 VTAIL.n264 B 0.012681f
C481 VTAIL.n265 B 0.029974f
C482 VTAIL.n266 B 0.013427f
C483 VTAIL.n267 B 0.0236f
C484 VTAIL.n268 B 0.012681f
C485 VTAIL.n269 B 0.029974f
C486 VTAIL.n270 B 0.013427f
C487 VTAIL.n271 B 0.0236f
C488 VTAIL.n272 B 0.012681f
C489 VTAIL.n273 B 0.029974f
C490 VTAIL.n274 B 0.013427f
C491 VTAIL.n275 B 0.0236f
C492 VTAIL.n276 B 0.012681f
C493 VTAIL.n277 B 0.029974f
C494 VTAIL.n278 B 0.013427f
C495 VTAIL.n279 B 0.152028f
C496 VTAIL.t3 B 0.049398f
C497 VTAIL.n280 B 0.022481f
C498 VTAIL.n281 B 0.017707f
C499 VTAIL.n282 B 0.012681f
C500 VTAIL.n283 B 1.50082f
C501 VTAIL.n284 B 0.0236f
C502 VTAIL.n285 B 0.012681f
C503 VTAIL.n286 B 0.013427f
C504 VTAIL.n287 B 0.029974f
C505 VTAIL.n288 B 0.029974f
C506 VTAIL.n289 B 0.013427f
C507 VTAIL.n290 B 0.012681f
C508 VTAIL.n291 B 0.0236f
C509 VTAIL.n292 B 0.0236f
C510 VTAIL.n293 B 0.012681f
C511 VTAIL.n294 B 0.013427f
C512 VTAIL.n295 B 0.029974f
C513 VTAIL.n296 B 0.029974f
C514 VTAIL.n297 B 0.013427f
C515 VTAIL.n298 B 0.012681f
C516 VTAIL.n299 B 0.0236f
C517 VTAIL.n300 B 0.0236f
C518 VTAIL.n301 B 0.012681f
C519 VTAIL.n302 B 0.013427f
C520 VTAIL.n303 B 0.029974f
C521 VTAIL.n304 B 0.029974f
C522 VTAIL.n305 B 0.013427f
C523 VTAIL.n306 B 0.012681f
C524 VTAIL.n307 B 0.0236f
C525 VTAIL.n308 B 0.0236f
C526 VTAIL.n309 B 0.012681f
C527 VTAIL.n310 B 0.013427f
C528 VTAIL.n311 B 0.029974f
C529 VTAIL.n312 B 0.029974f
C530 VTAIL.n313 B 0.013427f
C531 VTAIL.n314 B 0.012681f
C532 VTAIL.n315 B 0.0236f
C533 VTAIL.n316 B 0.0236f
C534 VTAIL.n317 B 0.012681f
C535 VTAIL.n318 B 0.013427f
C536 VTAIL.n319 B 0.029974f
C537 VTAIL.n320 B 0.029974f
C538 VTAIL.n321 B 0.029974f
C539 VTAIL.n322 B 0.013427f
C540 VTAIL.n323 B 0.012681f
C541 VTAIL.n324 B 0.0236f
C542 VTAIL.n325 B 0.0236f
C543 VTAIL.n326 B 0.012681f
C544 VTAIL.n327 B 0.013054f
C545 VTAIL.n328 B 0.013054f
C546 VTAIL.n329 B 0.029974f
C547 VTAIL.n330 B 0.060384f
C548 VTAIL.n331 B 0.013427f
C549 VTAIL.n332 B 0.012681f
C550 VTAIL.n333 B 0.055839f
C551 VTAIL.n334 B 0.033363f
C552 VTAIL.n335 B 1.42901f
C553 VDD1.n0 B 0.02967f
C554 VDD1.n1 B 0.022865f
C555 VDD1.n2 B 0.012287f
C556 VDD1.n3 B 0.029041f
C557 VDD1.n4 B 0.013009f
C558 VDD1.n5 B 0.022865f
C559 VDD1.n6 B 0.012287f
C560 VDD1.n7 B 0.029041f
C561 VDD1.n8 B 0.029041f
C562 VDD1.n9 B 0.013009f
C563 VDD1.n10 B 0.022865f
C564 VDD1.n11 B 0.012287f
C565 VDD1.n12 B 0.029041f
C566 VDD1.n13 B 0.013009f
C567 VDD1.n14 B 0.022865f
C568 VDD1.n15 B 0.012287f
C569 VDD1.n16 B 0.029041f
C570 VDD1.n17 B 0.013009f
C571 VDD1.n18 B 0.022865f
C572 VDD1.n19 B 0.012287f
C573 VDD1.n20 B 0.029041f
C574 VDD1.n21 B 0.013009f
C575 VDD1.n22 B 0.022865f
C576 VDD1.n23 B 0.012287f
C577 VDD1.n24 B 0.029041f
C578 VDD1.n25 B 0.013009f
C579 VDD1.n26 B 0.147296f
C580 VDD1.t0 B 0.04786f
C581 VDD1.n27 B 0.021781f
C582 VDD1.n28 B 0.017156f
C583 VDD1.n29 B 0.012287f
C584 VDD1.n30 B 1.4541f
C585 VDD1.n31 B 0.022865f
C586 VDD1.n32 B 0.012287f
C587 VDD1.n33 B 0.013009f
C588 VDD1.n34 B 0.029041f
C589 VDD1.n35 B 0.029041f
C590 VDD1.n36 B 0.013009f
C591 VDD1.n37 B 0.012287f
C592 VDD1.n38 B 0.022865f
C593 VDD1.n39 B 0.022865f
C594 VDD1.n40 B 0.012287f
C595 VDD1.n41 B 0.013009f
C596 VDD1.n42 B 0.029041f
C597 VDD1.n43 B 0.029041f
C598 VDD1.n44 B 0.013009f
C599 VDD1.n45 B 0.012287f
C600 VDD1.n46 B 0.022865f
C601 VDD1.n47 B 0.022865f
C602 VDD1.n48 B 0.012287f
C603 VDD1.n49 B 0.013009f
C604 VDD1.n50 B 0.029041f
C605 VDD1.n51 B 0.029041f
C606 VDD1.n52 B 0.013009f
C607 VDD1.n53 B 0.012287f
C608 VDD1.n54 B 0.022865f
C609 VDD1.n55 B 0.022865f
C610 VDD1.n56 B 0.012287f
C611 VDD1.n57 B 0.013009f
C612 VDD1.n58 B 0.029041f
C613 VDD1.n59 B 0.029041f
C614 VDD1.n60 B 0.013009f
C615 VDD1.n61 B 0.012287f
C616 VDD1.n62 B 0.022865f
C617 VDD1.n63 B 0.022865f
C618 VDD1.n64 B 0.012287f
C619 VDD1.n65 B 0.013009f
C620 VDD1.n66 B 0.029041f
C621 VDD1.n67 B 0.029041f
C622 VDD1.n68 B 0.013009f
C623 VDD1.n69 B 0.012287f
C624 VDD1.n70 B 0.022865f
C625 VDD1.n71 B 0.022865f
C626 VDD1.n72 B 0.012287f
C627 VDD1.n73 B 0.012648f
C628 VDD1.n74 B 0.012648f
C629 VDD1.n75 B 0.029041f
C630 VDD1.n76 B 0.058504f
C631 VDD1.n77 B 0.013009f
C632 VDD1.n78 B 0.012287f
C633 VDD1.n79 B 0.054101f
C634 VDD1.n80 B 0.049712f
C635 VDD1.n81 B 0.02967f
C636 VDD1.n82 B 0.022865f
C637 VDD1.n83 B 0.012287f
C638 VDD1.n84 B 0.029041f
C639 VDD1.n85 B 0.013009f
C640 VDD1.n86 B 0.022865f
C641 VDD1.n87 B 0.012287f
C642 VDD1.n88 B 0.029041f
C643 VDD1.n89 B 0.013009f
C644 VDD1.n90 B 0.022865f
C645 VDD1.n91 B 0.012287f
C646 VDD1.n92 B 0.029041f
C647 VDD1.n93 B 0.013009f
C648 VDD1.n94 B 0.022865f
C649 VDD1.n95 B 0.012287f
C650 VDD1.n96 B 0.029041f
C651 VDD1.n97 B 0.013009f
C652 VDD1.n98 B 0.022865f
C653 VDD1.n99 B 0.012287f
C654 VDD1.n100 B 0.029041f
C655 VDD1.n101 B 0.013009f
C656 VDD1.n102 B 0.022865f
C657 VDD1.n103 B 0.012287f
C658 VDD1.n104 B 0.029041f
C659 VDD1.n105 B 0.013009f
C660 VDD1.n106 B 0.147296f
C661 VDD1.t4 B 0.04786f
C662 VDD1.n107 B 0.021781f
C663 VDD1.n108 B 0.017156f
C664 VDD1.n109 B 0.012287f
C665 VDD1.n110 B 1.4541f
C666 VDD1.n111 B 0.022865f
C667 VDD1.n112 B 0.012287f
C668 VDD1.n113 B 0.013009f
C669 VDD1.n114 B 0.029041f
C670 VDD1.n115 B 0.029041f
C671 VDD1.n116 B 0.013009f
C672 VDD1.n117 B 0.012287f
C673 VDD1.n118 B 0.022865f
C674 VDD1.n119 B 0.022865f
C675 VDD1.n120 B 0.012287f
C676 VDD1.n121 B 0.013009f
C677 VDD1.n122 B 0.029041f
C678 VDD1.n123 B 0.029041f
C679 VDD1.n124 B 0.013009f
C680 VDD1.n125 B 0.012287f
C681 VDD1.n126 B 0.022865f
C682 VDD1.n127 B 0.022865f
C683 VDD1.n128 B 0.012287f
C684 VDD1.n129 B 0.013009f
C685 VDD1.n130 B 0.029041f
C686 VDD1.n131 B 0.029041f
C687 VDD1.n132 B 0.013009f
C688 VDD1.n133 B 0.012287f
C689 VDD1.n134 B 0.022865f
C690 VDD1.n135 B 0.022865f
C691 VDD1.n136 B 0.012287f
C692 VDD1.n137 B 0.013009f
C693 VDD1.n138 B 0.029041f
C694 VDD1.n139 B 0.029041f
C695 VDD1.n140 B 0.013009f
C696 VDD1.n141 B 0.012287f
C697 VDD1.n142 B 0.022865f
C698 VDD1.n143 B 0.022865f
C699 VDD1.n144 B 0.012287f
C700 VDD1.n145 B 0.013009f
C701 VDD1.n146 B 0.029041f
C702 VDD1.n147 B 0.029041f
C703 VDD1.n148 B 0.029041f
C704 VDD1.n149 B 0.013009f
C705 VDD1.n150 B 0.012287f
C706 VDD1.n151 B 0.022865f
C707 VDD1.n152 B 0.022865f
C708 VDD1.n153 B 0.012287f
C709 VDD1.n154 B 0.012648f
C710 VDD1.n155 B 0.012648f
C711 VDD1.n156 B 0.029041f
C712 VDD1.n157 B 0.058504f
C713 VDD1.n158 B 0.013009f
C714 VDD1.n159 B 0.012287f
C715 VDD1.n160 B 0.054101f
C716 VDD1.n161 B 0.049382f
C717 VDD1.t2 B 0.265248f
C718 VDD1.t1 B 0.265248f
C719 VDD1.n162 B 2.39679f
C720 VDD1.n163 B 1.95649f
C721 VDD1.t5 B 0.265248f
C722 VDD1.t3 B 0.265248f
C723 VDD1.n164 B 2.39593f
C724 VDD1.n165 B 2.27404f
C725 VP.n0 B 0.044153f
C726 VP.n1 B 0.010019f
C727 VP.n2 B 0.190898f
C728 VP.t3 B 1.47396f
C729 VP.t4 B 1.47396f
C730 VP.t5 B 1.49992f
C731 VP.n3 B 0.547154f
C732 VP.n4 B 0.571544f
C733 VP.n5 B 0.010019f
C734 VP.n6 B 0.56725f
C735 VP.n7 B 1.94709f
C736 VP.t1 B 1.47396f
C737 VP.n8 B 0.56725f
C738 VP.n9 B 1.98349f
C739 VP.n10 B 0.044153f
C740 VP.n11 B 0.044153f
C741 VP.t0 B 1.47396f
C742 VP.n12 B 0.566433f
C743 VP.n13 B 0.010019f
C744 VP.t2 B 1.47396f
C745 VP.n14 B 0.56725f
C746 VP.n15 B 0.034217f
.ends

