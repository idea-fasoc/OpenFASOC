* NGSPICE file created from diff_pair_sample_0813.ext - technology: sky130A

.subckt diff_pair_sample_0813 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.52305 pd=3.5 as=1.2363 ps=7.12 w=3.17 l=3.73
X1 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.52305 pd=3.5 as=1.2363 ps=7.12 w=3.17 l=3.73
X2 VTAIL.t6 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0.52305 ps=3.5 w=3.17 l=3.73
X3 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0.52305 ps=3.5 w=3.17 l=3.73
X4 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0 ps=0 w=3.17 l=3.73
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0 ps=0 w=3.17 l=3.73
X6 VTAIL.t4 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0.52305 ps=3.5 w=3.17 l=3.73
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.52305 pd=3.5 as=1.2363 ps=7.12 w=3.17 l=3.73
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0 ps=0 w=3.17 l=3.73
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0 ps=0 w=3.17 l=3.73
X10 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2363 pd=7.12 as=0.52305 ps=3.5 w=3.17 l=3.73
X11 VDD1.t0 VP.t3 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.52305 pd=3.5 as=1.2363 ps=7.12 w=3.17 l=3.73
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n7 VP.n6 88.5994
R10 VP.n22 VP.n0 88.5994
R11 VP.n5 VP.t2 53.9665
R12 VP.n5 VP.t0 52.6338
R13 VP.n6 VP.n5 45.0006
R14 VP.n14 VP.n13 40.4934
R15 VP.n14 VP.n2 40.4934
R16 VP.n8 VP.n4 24.4675
R17 VP.n12 VP.n4 24.4675
R18 VP.n13 VP.n12 24.4675
R19 VP.n18 VP.n2 24.4675
R20 VP.n19 VP.n18 24.4675
R21 VP.n20 VP.n19 24.4675
R22 VP.n7 VP.t1 20.4823
R23 VP.n0 VP.t3 20.4823
R24 VP.n8 VP.n7 1.46852
R25 VP.n20 VP.n0 1.46852
R26 VP.n9 VP.n6 0.354971
R27 VP.n22 VP.n21 0.354971
R28 VP VP.n22 0.26696
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VTAIL.n122 VTAIL.n112 289.615
R38 VTAIL.n10 VTAIL.n0 289.615
R39 VTAIL.n26 VTAIL.n16 289.615
R40 VTAIL.n42 VTAIL.n32 289.615
R41 VTAIL.n106 VTAIL.n96 289.615
R42 VTAIL.n90 VTAIL.n80 289.615
R43 VTAIL.n74 VTAIL.n64 289.615
R44 VTAIL.n58 VTAIL.n48 289.615
R45 VTAIL.n116 VTAIL.n115 185
R46 VTAIL.n121 VTAIL.n120 185
R47 VTAIL.n123 VTAIL.n122 185
R48 VTAIL.n4 VTAIL.n3 185
R49 VTAIL.n9 VTAIL.n8 185
R50 VTAIL.n11 VTAIL.n10 185
R51 VTAIL.n20 VTAIL.n19 185
R52 VTAIL.n25 VTAIL.n24 185
R53 VTAIL.n27 VTAIL.n26 185
R54 VTAIL.n36 VTAIL.n35 185
R55 VTAIL.n41 VTAIL.n40 185
R56 VTAIL.n43 VTAIL.n42 185
R57 VTAIL.n107 VTAIL.n106 185
R58 VTAIL.n105 VTAIL.n104 185
R59 VTAIL.n100 VTAIL.n99 185
R60 VTAIL.n91 VTAIL.n90 185
R61 VTAIL.n89 VTAIL.n88 185
R62 VTAIL.n84 VTAIL.n83 185
R63 VTAIL.n75 VTAIL.n74 185
R64 VTAIL.n73 VTAIL.n72 185
R65 VTAIL.n68 VTAIL.n67 185
R66 VTAIL.n59 VTAIL.n58 185
R67 VTAIL.n57 VTAIL.n56 185
R68 VTAIL.n52 VTAIL.n51 185
R69 VTAIL.n117 VTAIL.t2 148.606
R70 VTAIL.n5 VTAIL.t1 148.606
R71 VTAIL.n21 VTAIL.t7 148.606
R72 VTAIL.n37 VTAIL.t6 148.606
R73 VTAIL.n101 VTAIL.t5 148.606
R74 VTAIL.n85 VTAIL.t4 148.606
R75 VTAIL.n69 VTAIL.t0 148.606
R76 VTAIL.n53 VTAIL.t3 148.606
R77 VTAIL.n121 VTAIL.n115 104.615
R78 VTAIL.n122 VTAIL.n121 104.615
R79 VTAIL.n9 VTAIL.n3 104.615
R80 VTAIL.n10 VTAIL.n9 104.615
R81 VTAIL.n25 VTAIL.n19 104.615
R82 VTAIL.n26 VTAIL.n25 104.615
R83 VTAIL.n41 VTAIL.n35 104.615
R84 VTAIL.n42 VTAIL.n41 104.615
R85 VTAIL.n106 VTAIL.n105 104.615
R86 VTAIL.n105 VTAIL.n99 104.615
R87 VTAIL.n90 VTAIL.n89 104.615
R88 VTAIL.n89 VTAIL.n83 104.615
R89 VTAIL.n74 VTAIL.n73 104.615
R90 VTAIL.n73 VTAIL.n67 104.615
R91 VTAIL.n58 VTAIL.n57 104.615
R92 VTAIL.n57 VTAIL.n51 104.615
R93 VTAIL.t2 VTAIL.n115 52.3082
R94 VTAIL.t1 VTAIL.n3 52.3082
R95 VTAIL.t7 VTAIL.n19 52.3082
R96 VTAIL.t6 VTAIL.n35 52.3082
R97 VTAIL.t5 VTAIL.n99 52.3082
R98 VTAIL.t4 VTAIL.n83 52.3082
R99 VTAIL.t0 VTAIL.n67 52.3082
R100 VTAIL.t3 VTAIL.n51 52.3082
R101 VTAIL.n127 VTAIL.n126 33.155
R102 VTAIL.n15 VTAIL.n14 33.155
R103 VTAIL.n31 VTAIL.n30 33.155
R104 VTAIL.n47 VTAIL.n46 33.155
R105 VTAIL.n111 VTAIL.n110 33.155
R106 VTAIL.n95 VTAIL.n94 33.155
R107 VTAIL.n79 VTAIL.n78 33.155
R108 VTAIL.n63 VTAIL.n62 33.155
R109 VTAIL.n127 VTAIL.n111 18.5996
R110 VTAIL.n63 VTAIL.n47 18.5996
R111 VTAIL.n117 VTAIL.n116 15.5966
R112 VTAIL.n5 VTAIL.n4 15.5966
R113 VTAIL.n21 VTAIL.n20 15.5966
R114 VTAIL.n37 VTAIL.n36 15.5966
R115 VTAIL.n101 VTAIL.n100 15.5966
R116 VTAIL.n85 VTAIL.n84 15.5966
R117 VTAIL.n69 VTAIL.n68 15.5966
R118 VTAIL.n53 VTAIL.n52 15.5966
R119 VTAIL.n120 VTAIL.n119 12.8005
R120 VTAIL.n8 VTAIL.n7 12.8005
R121 VTAIL.n24 VTAIL.n23 12.8005
R122 VTAIL.n40 VTAIL.n39 12.8005
R123 VTAIL.n104 VTAIL.n103 12.8005
R124 VTAIL.n88 VTAIL.n87 12.8005
R125 VTAIL.n72 VTAIL.n71 12.8005
R126 VTAIL.n56 VTAIL.n55 12.8005
R127 VTAIL.n123 VTAIL.n114 12.0247
R128 VTAIL.n11 VTAIL.n2 12.0247
R129 VTAIL.n27 VTAIL.n18 12.0247
R130 VTAIL.n43 VTAIL.n34 12.0247
R131 VTAIL.n107 VTAIL.n98 12.0247
R132 VTAIL.n91 VTAIL.n82 12.0247
R133 VTAIL.n75 VTAIL.n66 12.0247
R134 VTAIL.n59 VTAIL.n50 12.0247
R135 VTAIL.n124 VTAIL.n112 11.249
R136 VTAIL.n12 VTAIL.n0 11.249
R137 VTAIL.n28 VTAIL.n16 11.249
R138 VTAIL.n44 VTAIL.n32 11.249
R139 VTAIL.n108 VTAIL.n96 11.249
R140 VTAIL.n92 VTAIL.n80 11.249
R141 VTAIL.n76 VTAIL.n64 11.249
R142 VTAIL.n60 VTAIL.n48 11.249
R143 VTAIL.n126 VTAIL.n125 9.45567
R144 VTAIL.n14 VTAIL.n13 9.45567
R145 VTAIL.n30 VTAIL.n29 9.45567
R146 VTAIL.n46 VTAIL.n45 9.45567
R147 VTAIL.n110 VTAIL.n109 9.45567
R148 VTAIL.n94 VTAIL.n93 9.45567
R149 VTAIL.n78 VTAIL.n77 9.45567
R150 VTAIL.n62 VTAIL.n61 9.45567
R151 VTAIL.n125 VTAIL.n124 9.3005
R152 VTAIL.n114 VTAIL.n113 9.3005
R153 VTAIL.n119 VTAIL.n118 9.3005
R154 VTAIL.n13 VTAIL.n12 9.3005
R155 VTAIL.n2 VTAIL.n1 9.3005
R156 VTAIL.n7 VTAIL.n6 9.3005
R157 VTAIL.n29 VTAIL.n28 9.3005
R158 VTAIL.n18 VTAIL.n17 9.3005
R159 VTAIL.n23 VTAIL.n22 9.3005
R160 VTAIL.n45 VTAIL.n44 9.3005
R161 VTAIL.n34 VTAIL.n33 9.3005
R162 VTAIL.n39 VTAIL.n38 9.3005
R163 VTAIL.n109 VTAIL.n108 9.3005
R164 VTAIL.n98 VTAIL.n97 9.3005
R165 VTAIL.n103 VTAIL.n102 9.3005
R166 VTAIL.n93 VTAIL.n92 9.3005
R167 VTAIL.n82 VTAIL.n81 9.3005
R168 VTAIL.n87 VTAIL.n86 9.3005
R169 VTAIL.n77 VTAIL.n76 9.3005
R170 VTAIL.n66 VTAIL.n65 9.3005
R171 VTAIL.n71 VTAIL.n70 9.3005
R172 VTAIL.n61 VTAIL.n60 9.3005
R173 VTAIL.n50 VTAIL.n49 9.3005
R174 VTAIL.n55 VTAIL.n54 9.3005
R175 VTAIL.n118 VTAIL.n117 4.46457
R176 VTAIL.n6 VTAIL.n5 4.46457
R177 VTAIL.n22 VTAIL.n21 4.46457
R178 VTAIL.n38 VTAIL.n37 4.46457
R179 VTAIL.n102 VTAIL.n101 4.46457
R180 VTAIL.n86 VTAIL.n85 4.46457
R181 VTAIL.n70 VTAIL.n69 4.46457
R182 VTAIL.n54 VTAIL.n53 4.46457
R183 VTAIL.n79 VTAIL.n63 3.5005
R184 VTAIL.n111 VTAIL.n95 3.5005
R185 VTAIL.n47 VTAIL.n31 3.5005
R186 VTAIL.n126 VTAIL.n112 2.71565
R187 VTAIL.n14 VTAIL.n0 2.71565
R188 VTAIL.n30 VTAIL.n16 2.71565
R189 VTAIL.n46 VTAIL.n32 2.71565
R190 VTAIL.n110 VTAIL.n96 2.71565
R191 VTAIL.n94 VTAIL.n80 2.71565
R192 VTAIL.n78 VTAIL.n64 2.71565
R193 VTAIL.n62 VTAIL.n48 2.71565
R194 VTAIL.n124 VTAIL.n123 1.93989
R195 VTAIL.n12 VTAIL.n11 1.93989
R196 VTAIL.n28 VTAIL.n27 1.93989
R197 VTAIL.n44 VTAIL.n43 1.93989
R198 VTAIL.n108 VTAIL.n107 1.93989
R199 VTAIL.n92 VTAIL.n91 1.93989
R200 VTAIL.n76 VTAIL.n75 1.93989
R201 VTAIL.n60 VTAIL.n59 1.93989
R202 VTAIL VTAIL.n15 1.80869
R203 VTAIL VTAIL.n127 1.69231
R204 VTAIL.n120 VTAIL.n114 1.16414
R205 VTAIL.n8 VTAIL.n2 1.16414
R206 VTAIL.n24 VTAIL.n18 1.16414
R207 VTAIL.n40 VTAIL.n34 1.16414
R208 VTAIL.n104 VTAIL.n98 1.16414
R209 VTAIL.n88 VTAIL.n82 1.16414
R210 VTAIL.n72 VTAIL.n66 1.16414
R211 VTAIL.n56 VTAIL.n50 1.16414
R212 VTAIL.n95 VTAIL.n79 0.470328
R213 VTAIL.n31 VTAIL.n15 0.470328
R214 VTAIL.n119 VTAIL.n116 0.388379
R215 VTAIL.n7 VTAIL.n4 0.388379
R216 VTAIL.n23 VTAIL.n20 0.388379
R217 VTAIL.n39 VTAIL.n36 0.388379
R218 VTAIL.n103 VTAIL.n100 0.388379
R219 VTAIL.n87 VTAIL.n84 0.388379
R220 VTAIL.n71 VTAIL.n68 0.388379
R221 VTAIL.n55 VTAIL.n52 0.388379
R222 VTAIL.n118 VTAIL.n113 0.155672
R223 VTAIL.n125 VTAIL.n113 0.155672
R224 VTAIL.n6 VTAIL.n1 0.155672
R225 VTAIL.n13 VTAIL.n1 0.155672
R226 VTAIL.n22 VTAIL.n17 0.155672
R227 VTAIL.n29 VTAIL.n17 0.155672
R228 VTAIL.n38 VTAIL.n33 0.155672
R229 VTAIL.n45 VTAIL.n33 0.155672
R230 VTAIL.n109 VTAIL.n97 0.155672
R231 VTAIL.n102 VTAIL.n97 0.155672
R232 VTAIL.n93 VTAIL.n81 0.155672
R233 VTAIL.n86 VTAIL.n81 0.155672
R234 VTAIL.n77 VTAIL.n65 0.155672
R235 VTAIL.n70 VTAIL.n65 0.155672
R236 VTAIL.n61 VTAIL.n49 0.155672
R237 VTAIL.n54 VTAIL.n49 0.155672
R238 VDD1 VDD1.n1 116.192
R239 VDD1 VDD1.n0 78.777
R240 VDD1.n0 VDD1.t1 6.24656
R241 VDD1.n0 VDD1.t3 6.24656
R242 VDD1.n1 VDD1.t2 6.24656
R243 VDD1.n1 VDD1.t0 6.24656
R244 B.n570 B.n569 585
R245 B.n571 B.n570 585
R246 B.n186 B.n103 585
R247 B.n185 B.n184 585
R248 B.n183 B.n182 585
R249 B.n181 B.n180 585
R250 B.n179 B.n178 585
R251 B.n177 B.n176 585
R252 B.n175 B.n174 585
R253 B.n173 B.n172 585
R254 B.n171 B.n170 585
R255 B.n169 B.n168 585
R256 B.n167 B.n166 585
R257 B.n165 B.n164 585
R258 B.n163 B.n162 585
R259 B.n161 B.n160 585
R260 B.n159 B.n158 585
R261 B.n156 B.n155 585
R262 B.n154 B.n153 585
R263 B.n152 B.n151 585
R264 B.n150 B.n149 585
R265 B.n148 B.n147 585
R266 B.n146 B.n145 585
R267 B.n144 B.n143 585
R268 B.n142 B.n141 585
R269 B.n140 B.n139 585
R270 B.n138 B.n137 585
R271 B.n136 B.n135 585
R272 B.n134 B.n133 585
R273 B.n132 B.n131 585
R274 B.n130 B.n129 585
R275 B.n128 B.n127 585
R276 B.n126 B.n125 585
R277 B.n124 B.n123 585
R278 B.n122 B.n121 585
R279 B.n120 B.n119 585
R280 B.n118 B.n117 585
R281 B.n116 B.n115 585
R282 B.n114 B.n113 585
R283 B.n112 B.n111 585
R284 B.n110 B.n109 585
R285 B.n81 B.n80 585
R286 B.n568 B.n82 585
R287 B.n572 B.n82 585
R288 B.n567 B.n566 585
R289 B.n566 B.n78 585
R290 B.n565 B.n77 585
R291 B.n578 B.n77 585
R292 B.n564 B.n76 585
R293 B.n579 B.n76 585
R294 B.n563 B.n75 585
R295 B.n580 B.n75 585
R296 B.n562 B.n561 585
R297 B.n561 B.n71 585
R298 B.n560 B.n70 585
R299 B.n586 B.n70 585
R300 B.n559 B.n69 585
R301 B.n587 B.n69 585
R302 B.n558 B.n68 585
R303 B.n588 B.n68 585
R304 B.n557 B.n556 585
R305 B.n556 B.n67 585
R306 B.n555 B.n63 585
R307 B.n594 B.n63 585
R308 B.n554 B.n62 585
R309 B.n595 B.n62 585
R310 B.n553 B.n61 585
R311 B.n596 B.n61 585
R312 B.n552 B.n551 585
R313 B.n551 B.n57 585
R314 B.n550 B.n56 585
R315 B.n602 B.n56 585
R316 B.n549 B.n55 585
R317 B.n603 B.n55 585
R318 B.n548 B.n54 585
R319 B.n604 B.n54 585
R320 B.n547 B.n546 585
R321 B.n546 B.n50 585
R322 B.n545 B.n49 585
R323 B.n610 B.n49 585
R324 B.n544 B.n48 585
R325 B.n611 B.n48 585
R326 B.n543 B.n47 585
R327 B.n612 B.n47 585
R328 B.n542 B.n541 585
R329 B.n541 B.n43 585
R330 B.n540 B.n42 585
R331 B.n618 B.n42 585
R332 B.n539 B.n41 585
R333 B.n619 B.n41 585
R334 B.n538 B.n40 585
R335 B.n620 B.n40 585
R336 B.n537 B.n536 585
R337 B.n536 B.n36 585
R338 B.n535 B.n35 585
R339 B.n626 B.n35 585
R340 B.n534 B.n34 585
R341 B.n627 B.n34 585
R342 B.n533 B.n33 585
R343 B.n628 B.n33 585
R344 B.n532 B.n531 585
R345 B.n531 B.n29 585
R346 B.n530 B.n28 585
R347 B.n634 B.n28 585
R348 B.n529 B.n27 585
R349 B.n635 B.n27 585
R350 B.n528 B.n26 585
R351 B.n636 B.n26 585
R352 B.n527 B.n526 585
R353 B.n526 B.n22 585
R354 B.n525 B.n21 585
R355 B.n642 B.n21 585
R356 B.n524 B.n20 585
R357 B.n643 B.n20 585
R358 B.n523 B.n19 585
R359 B.n644 B.n19 585
R360 B.n522 B.n521 585
R361 B.n521 B.n15 585
R362 B.n520 B.n14 585
R363 B.n650 B.n14 585
R364 B.n519 B.n13 585
R365 B.n651 B.n13 585
R366 B.n518 B.n12 585
R367 B.n652 B.n12 585
R368 B.n517 B.n516 585
R369 B.n516 B.n8 585
R370 B.n515 B.n7 585
R371 B.n658 B.n7 585
R372 B.n514 B.n6 585
R373 B.n659 B.n6 585
R374 B.n513 B.n5 585
R375 B.n660 B.n5 585
R376 B.n512 B.n511 585
R377 B.n511 B.n4 585
R378 B.n510 B.n187 585
R379 B.n510 B.n509 585
R380 B.n500 B.n188 585
R381 B.n189 B.n188 585
R382 B.n502 B.n501 585
R383 B.n503 B.n502 585
R384 B.n499 B.n194 585
R385 B.n194 B.n193 585
R386 B.n498 B.n497 585
R387 B.n497 B.n496 585
R388 B.n196 B.n195 585
R389 B.n197 B.n196 585
R390 B.n489 B.n488 585
R391 B.n490 B.n489 585
R392 B.n487 B.n202 585
R393 B.n202 B.n201 585
R394 B.n486 B.n485 585
R395 B.n485 B.n484 585
R396 B.n204 B.n203 585
R397 B.n205 B.n204 585
R398 B.n477 B.n476 585
R399 B.n478 B.n477 585
R400 B.n475 B.n210 585
R401 B.n210 B.n209 585
R402 B.n474 B.n473 585
R403 B.n473 B.n472 585
R404 B.n212 B.n211 585
R405 B.n213 B.n212 585
R406 B.n465 B.n464 585
R407 B.n466 B.n465 585
R408 B.n463 B.n218 585
R409 B.n218 B.n217 585
R410 B.n462 B.n461 585
R411 B.n461 B.n460 585
R412 B.n220 B.n219 585
R413 B.n221 B.n220 585
R414 B.n453 B.n452 585
R415 B.n454 B.n453 585
R416 B.n451 B.n226 585
R417 B.n226 B.n225 585
R418 B.n450 B.n449 585
R419 B.n449 B.n448 585
R420 B.n228 B.n227 585
R421 B.n229 B.n228 585
R422 B.n441 B.n440 585
R423 B.n442 B.n441 585
R424 B.n439 B.n234 585
R425 B.n234 B.n233 585
R426 B.n438 B.n437 585
R427 B.n437 B.n436 585
R428 B.n236 B.n235 585
R429 B.n237 B.n236 585
R430 B.n429 B.n428 585
R431 B.n430 B.n429 585
R432 B.n427 B.n242 585
R433 B.n242 B.n241 585
R434 B.n426 B.n425 585
R435 B.n425 B.n424 585
R436 B.n244 B.n243 585
R437 B.n245 B.n244 585
R438 B.n417 B.n416 585
R439 B.n418 B.n417 585
R440 B.n415 B.n250 585
R441 B.n250 B.n249 585
R442 B.n414 B.n413 585
R443 B.n413 B.n412 585
R444 B.n252 B.n251 585
R445 B.n405 B.n252 585
R446 B.n404 B.n403 585
R447 B.n406 B.n404 585
R448 B.n402 B.n257 585
R449 B.n257 B.n256 585
R450 B.n401 B.n400 585
R451 B.n400 B.n399 585
R452 B.n259 B.n258 585
R453 B.n260 B.n259 585
R454 B.n392 B.n391 585
R455 B.n393 B.n392 585
R456 B.n390 B.n265 585
R457 B.n265 B.n264 585
R458 B.n389 B.n388 585
R459 B.n388 B.n387 585
R460 B.n267 B.n266 585
R461 B.n268 B.n267 585
R462 B.n380 B.n379 585
R463 B.n381 B.n380 585
R464 B.n271 B.n270 585
R465 B.n299 B.n297 585
R466 B.n300 B.n296 585
R467 B.n300 B.n272 585
R468 B.n303 B.n302 585
R469 B.n304 B.n295 585
R470 B.n306 B.n305 585
R471 B.n308 B.n294 585
R472 B.n311 B.n310 585
R473 B.n312 B.n293 585
R474 B.n314 B.n313 585
R475 B.n316 B.n292 585
R476 B.n319 B.n318 585
R477 B.n320 B.n291 585
R478 B.n322 B.n321 585
R479 B.n324 B.n290 585
R480 B.n327 B.n326 585
R481 B.n329 B.n287 585
R482 B.n331 B.n330 585
R483 B.n333 B.n286 585
R484 B.n336 B.n335 585
R485 B.n337 B.n285 585
R486 B.n339 B.n338 585
R487 B.n341 B.n284 585
R488 B.n344 B.n343 585
R489 B.n345 B.n281 585
R490 B.n348 B.n347 585
R491 B.n350 B.n280 585
R492 B.n353 B.n352 585
R493 B.n354 B.n279 585
R494 B.n356 B.n355 585
R495 B.n358 B.n278 585
R496 B.n361 B.n360 585
R497 B.n362 B.n277 585
R498 B.n364 B.n363 585
R499 B.n366 B.n276 585
R500 B.n369 B.n368 585
R501 B.n370 B.n275 585
R502 B.n372 B.n371 585
R503 B.n374 B.n274 585
R504 B.n377 B.n376 585
R505 B.n378 B.n273 585
R506 B.n383 B.n382 585
R507 B.n382 B.n381 585
R508 B.n384 B.n269 585
R509 B.n269 B.n268 585
R510 B.n386 B.n385 585
R511 B.n387 B.n386 585
R512 B.n263 B.n262 585
R513 B.n264 B.n263 585
R514 B.n395 B.n394 585
R515 B.n394 B.n393 585
R516 B.n396 B.n261 585
R517 B.n261 B.n260 585
R518 B.n398 B.n397 585
R519 B.n399 B.n398 585
R520 B.n255 B.n254 585
R521 B.n256 B.n255 585
R522 B.n408 B.n407 585
R523 B.n407 B.n406 585
R524 B.n409 B.n253 585
R525 B.n405 B.n253 585
R526 B.n411 B.n410 585
R527 B.n412 B.n411 585
R528 B.n248 B.n247 585
R529 B.n249 B.n248 585
R530 B.n420 B.n419 585
R531 B.n419 B.n418 585
R532 B.n421 B.n246 585
R533 B.n246 B.n245 585
R534 B.n423 B.n422 585
R535 B.n424 B.n423 585
R536 B.n240 B.n239 585
R537 B.n241 B.n240 585
R538 B.n432 B.n431 585
R539 B.n431 B.n430 585
R540 B.n433 B.n238 585
R541 B.n238 B.n237 585
R542 B.n435 B.n434 585
R543 B.n436 B.n435 585
R544 B.n232 B.n231 585
R545 B.n233 B.n232 585
R546 B.n444 B.n443 585
R547 B.n443 B.n442 585
R548 B.n445 B.n230 585
R549 B.n230 B.n229 585
R550 B.n447 B.n446 585
R551 B.n448 B.n447 585
R552 B.n224 B.n223 585
R553 B.n225 B.n224 585
R554 B.n456 B.n455 585
R555 B.n455 B.n454 585
R556 B.n457 B.n222 585
R557 B.n222 B.n221 585
R558 B.n459 B.n458 585
R559 B.n460 B.n459 585
R560 B.n216 B.n215 585
R561 B.n217 B.n216 585
R562 B.n468 B.n467 585
R563 B.n467 B.n466 585
R564 B.n469 B.n214 585
R565 B.n214 B.n213 585
R566 B.n471 B.n470 585
R567 B.n472 B.n471 585
R568 B.n208 B.n207 585
R569 B.n209 B.n208 585
R570 B.n480 B.n479 585
R571 B.n479 B.n478 585
R572 B.n481 B.n206 585
R573 B.n206 B.n205 585
R574 B.n483 B.n482 585
R575 B.n484 B.n483 585
R576 B.n200 B.n199 585
R577 B.n201 B.n200 585
R578 B.n492 B.n491 585
R579 B.n491 B.n490 585
R580 B.n493 B.n198 585
R581 B.n198 B.n197 585
R582 B.n495 B.n494 585
R583 B.n496 B.n495 585
R584 B.n192 B.n191 585
R585 B.n193 B.n192 585
R586 B.n505 B.n504 585
R587 B.n504 B.n503 585
R588 B.n506 B.n190 585
R589 B.n190 B.n189 585
R590 B.n508 B.n507 585
R591 B.n509 B.n508 585
R592 B.n2 B.n0 585
R593 B.n4 B.n2 585
R594 B.n3 B.n1 585
R595 B.n659 B.n3 585
R596 B.n657 B.n656 585
R597 B.n658 B.n657 585
R598 B.n655 B.n9 585
R599 B.n9 B.n8 585
R600 B.n654 B.n653 585
R601 B.n653 B.n652 585
R602 B.n11 B.n10 585
R603 B.n651 B.n11 585
R604 B.n649 B.n648 585
R605 B.n650 B.n649 585
R606 B.n647 B.n16 585
R607 B.n16 B.n15 585
R608 B.n646 B.n645 585
R609 B.n645 B.n644 585
R610 B.n18 B.n17 585
R611 B.n643 B.n18 585
R612 B.n641 B.n640 585
R613 B.n642 B.n641 585
R614 B.n639 B.n23 585
R615 B.n23 B.n22 585
R616 B.n638 B.n637 585
R617 B.n637 B.n636 585
R618 B.n25 B.n24 585
R619 B.n635 B.n25 585
R620 B.n633 B.n632 585
R621 B.n634 B.n633 585
R622 B.n631 B.n30 585
R623 B.n30 B.n29 585
R624 B.n630 B.n629 585
R625 B.n629 B.n628 585
R626 B.n32 B.n31 585
R627 B.n627 B.n32 585
R628 B.n625 B.n624 585
R629 B.n626 B.n625 585
R630 B.n623 B.n37 585
R631 B.n37 B.n36 585
R632 B.n622 B.n621 585
R633 B.n621 B.n620 585
R634 B.n39 B.n38 585
R635 B.n619 B.n39 585
R636 B.n617 B.n616 585
R637 B.n618 B.n617 585
R638 B.n615 B.n44 585
R639 B.n44 B.n43 585
R640 B.n614 B.n613 585
R641 B.n613 B.n612 585
R642 B.n46 B.n45 585
R643 B.n611 B.n46 585
R644 B.n609 B.n608 585
R645 B.n610 B.n609 585
R646 B.n607 B.n51 585
R647 B.n51 B.n50 585
R648 B.n606 B.n605 585
R649 B.n605 B.n604 585
R650 B.n53 B.n52 585
R651 B.n603 B.n53 585
R652 B.n601 B.n600 585
R653 B.n602 B.n601 585
R654 B.n599 B.n58 585
R655 B.n58 B.n57 585
R656 B.n598 B.n597 585
R657 B.n597 B.n596 585
R658 B.n60 B.n59 585
R659 B.n595 B.n60 585
R660 B.n593 B.n592 585
R661 B.n594 B.n593 585
R662 B.n591 B.n64 585
R663 B.n67 B.n64 585
R664 B.n590 B.n589 585
R665 B.n589 B.n588 585
R666 B.n66 B.n65 585
R667 B.n587 B.n66 585
R668 B.n585 B.n584 585
R669 B.n586 B.n585 585
R670 B.n583 B.n72 585
R671 B.n72 B.n71 585
R672 B.n582 B.n581 585
R673 B.n581 B.n580 585
R674 B.n74 B.n73 585
R675 B.n579 B.n74 585
R676 B.n577 B.n576 585
R677 B.n578 B.n577 585
R678 B.n575 B.n79 585
R679 B.n79 B.n78 585
R680 B.n574 B.n573 585
R681 B.n573 B.n572 585
R682 B.n662 B.n661 585
R683 B.n661 B.n660 585
R684 B.n382 B.n271 478.086
R685 B.n573 B.n81 478.086
R686 B.n380 B.n273 478.086
R687 B.n570 B.n82 478.086
R688 B.n571 B.n102 256.663
R689 B.n571 B.n101 256.663
R690 B.n571 B.n100 256.663
R691 B.n571 B.n99 256.663
R692 B.n571 B.n98 256.663
R693 B.n571 B.n97 256.663
R694 B.n571 B.n96 256.663
R695 B.n571 B.n95 256.663
R696 B.n571 B.n94 256.663
R697 B.n571 B.n93 256.663
R698 B.n571 B.n92 256.663
R699 B.n571 B.n91 256.663
R700 B.n571 B.n90 256.663
R701 B.n571 B.n89 256.663
R702 B.n571 B.n88 256.663
R703 B.n571 B.n87 256.663
R704 B.n571 B.n86 256.663
R705 B.n571 B.n85 256.663
R706 B.n571 B.n84 256.663
R707 B.n571 B.n83 256.663
R708 B.n298 B.n272 256.663
R709 B.n301 B.n272 256.663
R710 B.n307 B.n272 256.663
R711 B.n309 B.n272 256.663
R712 B.n315 B.n272 256.663
R713 B.n317 B.n272 256.663
R714 B.n323 B.n272 256.663
R715 B.n325 B.n272 256.663
R716 B.n332 B.n272 256.663
R717 B.n334 B.n272 256.663
R718 B.n340 B.n272 256.663
R719 B.n342 B.n272 256.663
R720 B.n349 B.n272 256.663
R721 B.n351 B.n272 256.663
R722 B.n357 B.n272 256.663
R723 B.n359 B.n272 256.663
R724 B.n365 B.n272 256.663
R725 B.n367 B.n272 256.663
R726 B.n373 B.n272 256.663
R727 B.n375 B.n272 256.663
R728 B.n282 B.t12 229.77
R729 B.n288 B.t8 229.77
R730 B.n106 B.t15 229.77
R731 B.n104 B.t4 229.77
R732 B.n282 B.t14 210.337
R733 B.n104 B.t6 210.337
R734 B.n288 B.t11 210.337
R735 B.n106 B.t16 210.337
R736 B.n382 B.n269 163.367
R737 B.n386 B.n269 163.367
R738 B.n386 B.n263 163.367
R739 B.n394 B.n263 163.367
R740 B.n394 B.n261 163.367
R741 B.n398 B.n261 163.367
R742 B.n398 B.n255 163.367
R743 B.n407 B.n255 163.367
R744 B.n407 B.n253 163.367
R745 B.n411 B.n253 163.367
R746 B.n411 B.n248 163.367
R747 B.n419 B.n248 163.367
R748 B.n419 B.n246 163.367
R749 B.n423 B.n246 163.367
R750 B.n423 B.n240 163.367
R751 B.n431 B.n240 163.367
R752 B.n431 B.n238 163.367
R753 B.n435 B.n238 163.367
R754 B.n435 B.n232 163.367
R755 B.n443 B.n232 163.367
R756 B.n443 B.n230 163.367
R757 B.n447 B.n230 163.367
R758 B.n447 B.n224 163.367
R759 B.n455 B.n224 163.367
R760 B.n455 B.n222 163.367
R761 B.n459 B.n222 163.367
R762 B.n459 B.n216 163.367
R763 B.n467 B.n216 163.367
R764 B.n467 B.n214 163.367
R765 B.n471 B.n214 163.367
R766 B.n471 B.n208 163.367
R767 B.n479 B.n208 163.367
R768 B.n479 B.n206 163.367
R769 B.n483 B.n206 163.367
R770 B.n483 B.n200 163.367
R771 B.n491 B.n200 163.367
R772 B.n491 B.n198 163.367
R773 B.n495 B.n198 163.367
R774 B.n495 B.n192 163.367
R775 B.n504 B.n192 163.367
R776 B.n504 B.n190 163.367
R777 B.n508 B.n190 163.367
R778 B.n508 B.n2 163.367
R779 B.n661 B.n2 163.367
R780 B.n661 B.n3 163.367
R781 B.n657 B.n3 163.367
R782 B.n657 B.n9 163.367
R783 B.n653 B.n9 163.367
R784 B.n653 B.n11 163.367
R785 B.n649 B.n11 163.367
R786 B.n649 B.n16 163.367
R787 B.n645 B.n16 163.367
R788 B.n645 B.n18 163.367
R789 B.n641 B.n18 163.367
R790 B.n641 B.n23 163.367
R791 B.n637 B.n23 163.367
R792 B.n637 B.n25 163.367
R793 B.n633 B.n25 163.367
R794 B.n633 B.n30 163.367
R795 B.n629 B.n30 163.367
R796 B.n629 B.n32 163.367
R797 B.n625 B.n32 163.367
R798 B.n625 B.n37 163.367
R799 B.n621 B.n37 163.367
R800 B.n621 B.n39 163.367
R801 B.n617 B.n39 163.367
R802 B.n617 B.n44 163.367
R803 B.n613 B.n44 163.367
R804 B.n613 B.n46 163.367
R805 B.n609 B.n46 163.367
R806 B.n609 B.n51 163.367
R807 B.n605 B.n51 163.367
R808 B.n605 B.n53 163.367
R809 B.n601 B.n53 163.367
R810 B.n601 B.n58 163.367
R811 B.n597 B.n58 163.367
R812 B.n597 B.n60 163.367
R813 B.n593 B.n60 163.367
R814 B.n593 B.n64 163.367
R815 B.n589 B.n64 163.367
R816 B.n589 B.n66 163.367
R817 B.n585 B.n66 163.367
R818 B.n585 B.n72 163.367
R819 B.n581 B.n72 163.367
R820 B.n581 B.n74 163.367
R821 B.n577 B.n74 163.367
R822 B.n577 B.n79 163.367
R823 B.n573 B.n79 163.367
R824 B.n300 B.n299 163.367
R825 B.n302 B.n300 163.367
R826 B.n306 B.n295 163.367
R827 B.n310 B.n308 163.367
R828 B.n314 B.n293 163.367
R829 B.n318 B.n316 163.367
R830 B.n322 B.n291 163.367
R831 B.n326 B.n324 163.367
R832 B.n331 B.n287 163.367
R833 B.n335 B.n333 163.367
R834 B.n339 B.n285 163.367
R835 B.n343 B.n341 163.367
R836 B.n348 B.n281 163.367
R837 B.n352 B.n350 163.367
R838 B.n356 B.n279 163.367
R839 B.n360 B.n358 163.367
R840 B.n364 B.n277 163.367
R841 B.n368 B.n366 163.367
R842 B.n372 B.n275 163.367
R843 B.n376 B.n374 163.367
R844 B.n380 B.n267 163.367
R845 B.n388 B.n267 163.367
R846 B.n388 B.n265 163.367
R847 B.n392 B.n265 163.367
R848 B.n392 B.n259 163.367
R849 B.n400 B.n259 163.367
R850 B.n400 B.n257 163.367
R851 B.n404 B.n257 163.367
R852 B.n404 B.n252 163.367
R853 B.n413 B.n252 163.367
R854 B.n413 B.n250 163.367
R855 B.n417 B.n250 163.367
R856 B.n417 B.n244 163.367
R857 B.n425 B.n244 163.367
R858 B.n425 B.n242 163.367
R859 B.n429 B.n242 163.367
R860 B.n429 B.n236 163.367
R861 B.n437 B.n236 163.367
R862 B.n437 B.n234 163.367
R863 B.n441 B.n234 163.367
R864 B.n441 B.n228 163.367
R865 B.n449 B.n228 163.367
R866 B.n449 B.n226 163.367
R867 B.n453 B.n226 163.367
R868 B.n453 B.n220 163.367
R869 B.n461 B.n220 163.367
R870 B.n461 B.n218 163.367
R871 B.n465 B.n218 163.367
R872 B.n465 B.n212 163.367
R873 B.n473 B.n212 163.367
R874 B.n473 B.n210 163.367
R875 B.n477 B.n210 163.367
R876 B.n477 B.n204 163.367
R877 B.n485 B.n204 163.367
R878 B.n485 B.n202 163.367
R879 B.n489 B.n202 163.367
R880 B.n489 B.n196 163.367
R881 B.n497 B.n196 163.367
R882 B.n497 B.n194 163.367
R883 B.n502 B.n194 163.367
R884 B.n502 B.n188 163.367
R885 B.n510 B.n188 163.367
R886 B.n511 B.n510 163.367
R887 B.n511 B.n5 163.367
R888 B.n6 B.n5 163.367
R889 B.n7 B.n6 163.367
R890 B.n516 B.n7 163.367
R891 B.n516 B.n12 163.367
R892 B.n13 B.n12 163.367
R893 B.n14 B.n13 163.367
R894 B.n521 B.n14 163.367
R895 B.n521 B.n19 163.367
R896 B.n20 B.n19 163.367
R897 B.n21 B.n20 163.367
R898 B.n526 B.n21 163.367
R899 B.n526 B.n26 163.367
R900 B.n27 B.n26 163.367
R901 B.n28 B.n27 163.367
R902 B.n531 B.n28 163.367
R903 B.n531 B.n33 163.367
R904 B.n34 B.n33 163.367
R905 B.n35 B.n34 163.367
R906 B.n536 B.n35 163.367
R907 B.n536 B.n40 163.367
R908 B.n41 B.n40 163.367
R909 B.n42 B.n41 163.367
R910 B.n541 B.n42 163.367
R911 B.n541 B.n47 163.367
R912 B.n48 B.n47 163.367
R913 B.n49 B.n48 163.367
R914 B.n546 B.n49 163.367
R915 B.n546 B.n54 163.367
R916 B.n55 B.n54 163.367
R917 B.n56 B.n55 163.367
R918 B.n551 B.n56 163.367
R919 B.n551 B.n61 163.367
R920 B.n62 B.n61 163.367
R921 B.n63 B.n62 163.367
R922 B.n556 B.n63 163.367
R923 B.n556 B.n68 163.367
R924 B.n69 B.n68 163.367
R925 B.n70 B.n69 163.367
R926 B.n561 B.n70 163.367
R927 B.n561 B.n75 163.367
R928 B.n76 B.n75 163.367
R929 B.n77 B.n76 163.367
R930 B.n566 B.n77 163.367
R931 B.n566 B.n82 163.367
R932 B.n111 B.n110 163.367
R933 B.n115 B.n114 163.367
R934 B.n119 B.n118 163.367
R935 B.n123 B.n122 163.367
R936 B.n127 B.n126 163.367
R937 B.n131 B.n130 163.367
R938 B.n135 B.n134 163.367
R939 B.n139 B.n138 163.367
R940 B.n143 B.n142 163.367
R941 B.n147 B.n146 163.367
R942 B.n151 B.n150 163.367
R943 B.n155 B.n154 163.367
R944 B.n160 B.n159 163.367
R945 B.n164 B.n163 163.367
R946 B.n168 B.n167 163.367
R947 B.n172 B.n171 163.367
R948 B.n176 B.n175 163.367
R949 B.n180 B.n179 163.367
R950 B.n184 B.n183 163.367
R951 B.n570 B.n103 163.367
R952 B.n381 B.n272 155.004
R953 B.n572 B.n571 155.004
R954 B.n283 B.t13 131.597
R955 B.n105 B.t7 131.597
R956 B.n289 B.t10 131.597
R957 B.n107 B.t17 131.597
R958 B.n381 B.n268 88.5736
R959 B.n387 B.n268 88.5736
R960 B.n387 B.n264 88.5736
R961 B.n393 B.n264 88.5736
R962 B.n393 B.n260 88.5736
R963 B.n399 B.n260 88.5736
R964 B.n399 B.n256 88.5736
R965 B.n406 B.n256 88.5736
R966 B.n406 B.n405 88.5736
R967 B.n412 B.n249 88.5736
R968 B.n418 B.n249 88.5736
R969 B.n418 B.n245 88.5736
R970 B.n424 B.n245 88.5736
R971 B.n424 B.n241 88.5736
R972 B.n430 B.n241 88.5736
R973 B.n430 B.n237 88.5736
R974 B.n436 B.n237 88.5736
R975 B.n436 B.n233 88.5736
R976 B.n442 B.n233 88.5736
R977 B.n442 B.n229 88.5736
R978 B.n448 B.n229 88.5736
R979 B.n448 B.n225 88.5736
R980 B.n454 B.n225 88.5736
R981 B.n460 B.n221 88.5736
R982 B.n460 B.n217 88.5736
R983 B.n466 B.n217 88.5736
R984 B.n466 B.n213 88.5736
R985 B.n472 B.n213 88.5736
R986 B.n472 B.n209 88.5736
R987 B.n478 B.n209 88.5736
R988 B.n478 B.n205 88.5736
R989 B.n484 B.n205 88.5736
R990 B.n484 B.n201 88.5736
R991 B.n490 B.n201 88.5736
R992 B.n496 B.n197 88.5736
R993 B.n496 B.n193 88.5736
R994 B.n503 B.n193 88.5736
R995 B.n503 B.n189 88.5736
R996 B.n509 B.n189 88.5736
R997 B.n509 B.n4 88.5736
R998 B.n660 B.n4 88.5736
R999 B.n660 B.n659 88.5736
R1000 B.n659 B.n658 88.5736
R1001 B.n658 B.n8 88.5736
R1002 B.n652 B.n8 88.5736
R1003 B.n652 B.n651 88.5736
R1004 B.n651 B.n650 88.5736
R1005 B.n650 B.n15 88.5736
R1006 B.n644 B.n643 88.5736
R1007 B.n643 B.n642 88.5736
R1008 B.n642 B.n22 88.5736
R1009 B.n636 B.n22 88.5736
R1010 B.n636 B.n635 88.5736
R1011 B.n635 B.n634 88.5736
R1012 B.n634 B.n29 88.5736
R1013 B.n628 B.n29 88.5736
R1014 B.n628 B.n627 88.5736
R1015 B.n627 B.n626 88.5736
R1016 B.n626 B.n36 88.5736
R1017 B.n620 B.n619 88.5736
R1018 B.n619 B.n618 88.5736
R1019 B.n618 B.n43 88.5736
R1020 B.n612 B.n43 88.5736
R1021 B.n612 B.n611 88.5736
R1022 B.n611 B.n610 88.5736
R1023 B.n610 B.n50 88.5736
R1024 B.n604 B.n50 88.5736
R1025 B.n604 B.n603 88.5736
R1026 B.n603 B.n602 88.5736
R1027 B.n602 B.n57 88.5736
R1028 B.n596 B.n57 88.5736
R1029 B.n596 B.n595 88.5736
R1030 B.n595 B.n594 88.5736
R1031 B.n588 B.n67 88.5736
R1032 B.n588 B.n587 88.5736
R1033 B.n587 B.n586 88.5736
R1034 B.n586 B.n71 88.5736
R1035 B.n580 B.n71 88.5736
R1036 B.n580 B.n579 88.5736
R1037 B.n579 B.n578 88.5736
R1038 B.n578 B.n78 88.5736
R1039 B.n572 B.n78 88.5736
R1040 B.n283 B.n282 78.7399
R1041 B.n289 B.n288 78.7399
R1042 B.n107 B.n106 78.7399
R1043 B.n105 B.n104 78.7399
R1044 B.n298 B.n271 71.676
R1045 B.n302 B.n301 71.676
R1046 B.n307 B.n306 71.676
R1047 B.n310 B.n309 71.676
R1048 B.n315 B.n314 71.676
R1049 B.n318 B.n317 71.676
R1050 B.n323 B.n322 71.676
R1051 B.n326 B.n325 71.676
R1052 B.n332 B.n331 71.676
R1053 B.n335 B.n334 71.676
R1054 B.n340 B.n339 71.676
R1055 B.n343 B.n342 71.676
R1056 B.n349 B.n348 71.676
R1057 B.n352 B.n351 71.676
R1058 B.n357 B.n356 71.676
R1059 B.n360 B.n359 71.676
R1060 B.n365 B.n364 71.676
R1061 B.n368 B.n367 71.676
R1062 B.n373 B.n372 71.676
R1063 B.n376 B.n375 71.676
R1064 B.n83 B.n81 71.676
R1065 B.n111 B.n84 71.676
R1066 B.n115 B.n85 71.676
R1067 B.n119 B.n86 71.676
R1068 B.n123 B.n87 71.676
R1069 B.n127 B.n88 71.676
R1070 B.n131 B.n89 71.676
R1071 B.n135 B.n90 71.676
R1072 B.n139 B.n91 71.676
R1073 B.n143 B.n92 71.676
R1074 B.n147 B.n93 71.676
R1075 B.n151 B.n94 71.676
R1076 B.n155 B.n95 71.676
R1077 B.n160 B.n96 71.676
R1078 B.n164 B.n97 71.676
R1079 B.n168 B.n98 71.676
R1080 B.n172 B.n99 71.676
R1081 B.n176 B.n100 71.676
R1082 B.n180 B.n101 71.676
R1083 B.n184 B.n102 71.676
R1084 B.n103 B.n102 71.676
R1085 B.n183 B.n101 71.676
R1086 B.n179 B.n100 71.676
R1087 B.n175 B.n99 71.676
R1088 B.n171 B.n98 71.676
R1089 B.n167 B.n97 71.676
R1090 B.n163 B.n96 71.676
R1091 B.n159 B.n95 71.676
R1092 B.n154 B.n94 71.676
R1093 B.n150 B.n93 71.676
R1094 B.n146 B.n92 71.676
R1095 B.n142 B.n91 71.676
R1096 B.n138 B.n90 71.676
R1097 B.n134 B.n89 71.676
R1098 B.n130 B.n88 71.676
R1099 B.n126 B.n87 71.676
R1100 B.n122 B.n86 71.676
R1101 B.n118 B.n85 71.676
R1102 B.n114 B.n84 71.676
R1103 B.n110 B.n83 71.676
R1104 B.n299 B.n298 71.676
R1105 B.n301 B.n295 71.676
R1106 B.n308 B.n307 71.676
R1107 B.n309 B.n293 71.676
R1108 B.n316 B.n315 71.676
R1109 B.n317 B.n291 71.676
R1110 B.n324 B.n323 71.676
R1111 B.n325 B.n287 71.676
R1112 B.n333 B.n332 71.676
R1113 B.n334 B.n285 71.676
R1114 B.n341 B.n340 71.676
R1115 B.n342 B.n281 71.676
R1116 B.n350 B.n349 71.676
R1117 B.n351 B.n279 71.676
R1118 B.n358 B.n357 71.676
R1119 B.n359 B.n277 71.676
R1120 B.n366 B.n365 71.676
R1121 B.n367 B.n275 71.676
R1122 B.n374 B.n373 71.676
R1123 B.n375 B.n273 71.676
R1124 B.n346 B.n283 59.5399
R1125 B.n328 B.n289 59.5399
R1126 B.n108 B.n107 59.5399
R1127 B.n157 B.n105 59.5399
R1128 B.n412 B.t9 58.6151
R1129 B.n594 B.t5 58.6151
R1130 B.t0 B.n197 50.7998
R1131 B.t1 B.n15 50.7998
R1132 B.t3 B.n221 45.5896
R1133 B.t2 B.n36 45.5896
R1134 B.n454 B.t3 42.9845
R1135 B.n620 B.t2 42.9845
R1136 B.n490 B.t0 37.7743
R1137 B.n644 B.t1 37.7743
R1138 B.n574 B.n80 31.0639
R1139 B.n569 B.n568 31.0639
R1140 B.n379 B.n378 31.0639
R1141 B.n383 B.n270 31.0639
R1142 B.n405 B.t9 29.9591
R1143 B.n67 B.t5 29.9591
R1144 B B.n662 18.0485
R1145 B.n109 B.n80 10.6151
R1146 B.n112 B.n109 10.6151
R1147 B.n113 B.n112 10.6151
R1148 B.n116 B.n113 10.6151
R1149 B.n117 B.n116 10.6151
R1150 B.n120 B.n117 10.6151
R1151 B.n121 B.n120 10.6151
R1152 B.n124 B.n121 10.6151
R1153 B.n125 B.n124 10.6151
R1154 B.n128 B.n125 10.6151
R1155 B.n129 B.n128 10.6151
R1156 B.n132 B.n129 10.6151
R1157 B.n133 B.n132 10.6151
R1158 B.n136 B.n133 10.6151
R1159 B.n137 B.n136 10.6151
R1160 B.n141 B.n140 10.6151
R1161 B.n144 B.n141 10.6151
R1162 B.n145 B.n144 10.6151
R1163 B.n148 B.n145 10.6151
R1164 B.n149 B.n148 10.6151
R1165 B.n152 B.n149 10.6151
R1166 B.n153 B.n152 10.6151
R1167 B.n156 B.n153 10.6151
R1168 B.n161 B.n158 10.6151
R1169 B.n162 B.n161 10.6151
R1170 B.n165 B.n162 10.6151
R1171 B.n166 B.n165 10.6151
R1172 B.n169 B.n166 10.6151
R1173 B.n170 B.n169 10.6151
R1174 B.n173 B.n170 10.6151
R1175 B.n174 B.n173 10.6151
R1176 B.n177 B.n174 10.6151
R1177 B.n178 B.n177 10.6151
R1178 B.n181 B.n178 10.6151
R1179 B.n182 B.n181 10.6151
R1180 B.n185 B.n182 10.6151
R1181 B.n186 B.n185 10.6151
R1182 B.n569 B.n186 10.6151
R1183 B.n379 B.n266 10.6151
R1184 B.n389 B.n266 10.6151
R1185 B.n390 B.n389 10.6151
R1186 B.n391 B.n390 10.6151
R1187 B.n391 B.n258 10.6151
R1188 B.n401 B.n258 10.6151
R1189 B.n402 B.n401 10.6151
R1190 B.n403 B.n402 10.6151
R1191 B.n403 B.n251 10.6151
R1192 B.n414 B.n251 10.6151
R1193 B.n415 B.n414 10.6151
R1194 B.n416 B.n415 10.6151
R1195 B.n416 B.n243 10.6151
R1196 B.n426 B.n243 10.6151
R1197 B.n427 B.n426 10.6151
R1198 B.n428 B.n427 10.6151
R1199 B.n428 B.n235 10.6151
R1200 B.n438 B.n235 10.6151
R1201 B.n439 B.n438 10.6151
R1202 B.n440 B.n439 10.6151
R1203 B.n440 B.n227 10.6151
R1204 B.n450 B.n227 10.6151
R1205 B.n451 B.n450 10.6151
R1206 B.n452 B.n451 10.6151
R1207 B.n452 B.n219 10.6151
R1208 B.n462 B.n219 10.6151
R1209 B.n463 B.n462 10.6151
R1210 B.n464 B.n463 10.6151
R1211 B.n464 B.n211 10.6151
R1212 B.n474 B.n211 10.6151
R1213 B.n475 B.n474 10.6151
R1214 B.n476 B.n475 10.6151
R1215 B.n476 B.n203 10.6151
R1216 B.n486 B.n203 10.6151
R1217 B.n487 B.n486 10.6151
R1218 B.n488 B.n487 10.6151
R1219 B.n488 B.n195 10.6151
R1220 B.n498 B.n195 10.6151
R1221 B.n499 B.n498 10.6151
R1222 B.n501 B.n499 10.6151
R1223 B.n501 B.n500 10.6151
R1224 B.n500 B.n187 10.6151
R1225 B.n512 B.n187 10.6151
R1226 B.n513 B.n512 10.6151
R1227 B.n514 B.n513 10.6151
R1228 B.n515 B.n514 10.6151
R1229 B.n517 B.n515 10.6151
R1230 B.n518 B.n517 10.6151
R1231 B.n519 B.n518 10.6151
R1232 B.n520 B.n519 10.6151
R1233 B.n522 B.n520 10.6151
R1234 B.n523 B.n522 10.6151
R1235 B.n524 B.n523 10.6151
R1236 B.n525 B.n524 10.6151
R1237 B.n527 B.n525 10.6151
R1238 B.n528 B.n527 10.6151
R1239 B.n529 B.n528 10.6151
R1240 B.n530 B.n529 10.6151
R1241 B.n532 B.n530 10.6151
R1242 B.n533 B.n532 10.6151
R1243 B.n534 B.n533 10.6151
R1244 B.n535 B.n534 10.6151
R1245 B.n537 B.n535 10.6151
R1246 B.n538 B.n537 10.6151
R1247 B.n539 B.n538 10.6151
R1248 B.n540 B.n539 10.6151
R1249 B.n542 B.n540 10.6151
R1250 B.n543 B.n542 10.6151
R1251 B.n544 B.n543 10.6151
R1252 B.n545 B.n544 10.6151
R1253 B.n547 B.n545 10.6151
R1254 B.n548 B.n547 10.6151
R1255 B.n549 B.n548 10.6151
R1256 B.n550 B.n549 10.6151
R1257 B.n552 B.n550 10.6151
R1258 B.n553 B.n552 10.6151
R1259 B.n554 B.n553 10.6151
R1260 B.n555 B.n554 10.6151
R1261 B.n557 B.n555 10.6151
R1262 B.n558 B.n557 10.6151
R1263 B.n559 B.n558 10.6151
R1264 B.n560 B.n559 10.6151
R1265 B.n562 B.n560 10.6151
R1266 B.n563 B.n562 10.6151
R1267 B.n564 B.n563 10.6151
R1268 B.n565 B.n564 10.6151
R1269 B.n567 B.n565 10.6151
R1270 B.n568 B.n567 10.6151
R1271 B.n297 B.n270 10.6151
R1272 B.n297 B.n296 10.6151
R1273 B.n303 B.n296 10.6151
R1274 B.n304 B.n303 10.6151
R1275 B.n305 B.n304 10.6151
R1276 B.n305 B.n294 10.6151
R1277 B.n311 B.n294 10.6151
R1278 B.n312 B.n311 10.6151
R1279 B.n313 B.n312 10.6151
R1280 B.n313 B.n292 10.6151
R1281 B.n319 B.n292 10.6151
R1282 B.n320 B.n319 10.6151
R1283 B.n321 B.n320 10.6151
R1284 B.n321 B.n290 10.6151
R1285 B.n327 B.n290 10.6151
R1286 B.n330 B.n329 10.6151
R1287 B.n330 B.n286 10.6151
R1288 B.n336 B.n286 10.6151
R1289 B.n337 B.n336 10.6151
R1290 B.n338 B.n337 10.6151
R1291 B.n338 B.n284 10.6151
R1292 B.n344 B.n284 10.6151
R1293 B.n345 B.n344 10.6151
R1294 B.n347 B.n280 10.6151
R1295 B.n353 B.n280 10.6151
R1296 B.n354 B.n353 10.6151
R1297 B.n355 B.n354 10.6151
R1298 B.n355 B.n278 10.6151
R1299 B.n361 B.n278 10.6151
R1300 B.n362 B.n361 10.6151
R1301 B.n363 B.n362 10.6151
R1302 B.n363 B.n276 10.6151
R1303 B.n369 B.n276 10.6151
R1304 B.n370 B.n369 10.6151
R1305 B.n371 B.n370 10.6151
R1306 B.n371 B.n274 10.6151
R1307 B.n377 B.n274 10.6151
R1308 B.n378 B.n377 10.6151
R1309 B.n384 B.n383 10.6151
R1310 B.n385 B.n384 10.6151
R1311 B.n385 B.n262 10.6151
R1312 B.n395 B.n262 10.6151
R1313 B.n396 B.n395 10.6151
R1314 B.n397 B.n396 10.6151
R1315 B.n397 B.n254 10.6151
R1316 B.n408 B.n254 10.6151
R1317 B.n409 B.n408 10.6151
R1318 B.n410 B.n409 10.6151
R1319 B.n410 B.n247 10.6151
R1320 B.n420 B.n247 10.6151
R1321 B.n421 B.n420 10.6151
R1322 B.n422 B.n421 10.6151
R1323 B.n422 B.n239 10.6151
R1324 B.n432 B.n239 10.6151
R1325 B.n433 B.n432 10.6151
R1326 B.n434 B.n433 10.6151
R1327 B.n434 B.n231 10.6151
R1328 B.n444 B.n231 10.6151
R1329 B.n445 B.n444 10.6151
R1330 B.n446 B.n445 10.6151
R1331 B.n446 B.n223 10.6151
R1332 B.n456 B.n223 10.6151
R1333 B.n457 B.n456 10.6151
R1334 B.n458 B.n457 10.6151
R1335 B.n458 B.n215 10.6151
R1336 B.n468 B.n215 10.6151
R1337 B.n469 B.n468 10.6151
R1338 B.n470 B.n469 10.6151
R1339 B.n470 B.n207 10.6151
R1340 B.n480 B.n207 10.6151
R1341 B.n481 B.n480 10.6151
R1342 B.n482 B.n481 10.6151
R1343 B.n482 B.n199 10.6151
R1344 B.n492 B.n199 10.6151
R1345 B.n493 B.n492 10.6151
R1346 B.n494 B.n493 10.6151
R1347 B.n494 B.n191 10.6151
R1348 B.n505 B.n191 10.6151
R1349 B.n506 B.n505 10.6151
R1350 B.n507 B.n506 10.6151
R1351 B.n507 B.n0 10.6151
R1352 B.n656 B.n1 10.6151
R1353 B.n656 B.n655 10.6151
R1354 B.n655 B.n654 10.6151
R1355 B.n654 B.n10 10.6151
R1356 B.n648 B.n10 10.6151
R1357 B.n648 B.n647 10.6151
R1358 B.n647 B.n646 10.6151
R1359 B.n646 B.n17 10.6151
R1360 B.n640 B.n17 10.6151
R1361 B.n640 B.n639 10.6151
R1362 B.n639 B.n638 10.6151
R1363 B.n638 B.n24 10.6151
R1364 B.n632 B.n24 10.6151
R1365 B.n632 B.n631 10.6151
R1366 B.n631 B.n630 10.6151
R1367 B.n630 B.n31 10.6151
R1368 B.n624 B.n31 10.6151
R1369 B.n624 B.n623 10.6151
R1370 B.n623 B.n622 10.6151
R1371 B.n622 B.n38 10.6151
R1372 B.n616 B.n38 10.6151
R1373 B.n616 B.n615 10.6151
R1374 B.n615 B.n614 10.6151
R1375 B.n614 B.n45 10.6151
R1376 B.n608 B.n45 10.6151
R1377 B.n608 B.n607 10.6151
R1378 B.n607 B.n606 10.6151
R1379 B.n606 B.n52 10.6151
R1380 B.n600 B.n52 10.6151
R1381 B.n600 B.n599 10.6151
R1382 B.n599 B.n598 10.6151
R1383 B.n598 B.n59 10.6151
R1384 B.n592 B.n59 10.6151
R1385 B.n592 B.n591 10.6151
R1386 B.n591 B.n590 10.6151
R1387 B.n590 B.n65 10.6151
R1388 B.n584 B.n65 10.6151
R1389 B.n584 B.n583 10.6151
R1390 B.n583 B.n582 10.6151
R1391 B.n582 B.n73 10.6151
R1392 B.n576 B.n73 10.6151
R1393 B.n576 B.n575 10.6151
R1394 B.n575 B.n574 10.6151
R1395 B.n140 B.n108 6.5566
R1396 B.n157 B.n156 6.5566
R1397 B.n329 B.n328 6.5566
R1398 B.n346 B.n345 6.5566
R1399 B.n137 B.n108 4.05904
R1400 B.n158 B.n157 4.05904
R1401 B.n328 B.n327 4.05904
R1402 B.n347 B.n346 4.05904
R1403 B.n662 B.n0 2.81026
R1404 B.n662 B.n1 2.81026
R1405 VN.n0 VN.t3 53.9667
R1406 VN.n1 VN.t2 53.9667
R1407 VN.n0 VN.t0 52.6338
R1408 VN.n1 VN.t1 52.6338
R1409 VN VN.n1 45.1659
R1410 VN VN.n0 1.91213
R1411 VDD2.n2 VDD2.n0 115.666
R1412 VDD2.n2 VDD2.n1 78.7188
R1413 VDD2.n1 VDD2.t2 6.24656
R1414 VDD2.n1 VDD2.t1 6.24656
R1415 VDD2.n0 VDD2.t0 6.24656
R1416 VDD2.n0 VDD2.t3 6.24656
R1417 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 2.30105f
C1 VN VP 5.37918f
C2 VDD1 VDD2 1.29942f
C3 VTAIL VDD2 3.93504f
C4 VTAIL VDD1 3.87326f
C5 VN VDD2 1.57823f
C6 VP VDD2 0.471506f
C7 VN VDD1 0.154655f
C8 VTAIL VN 2.28694f
C9 VP VDD1 1.89329f
C10 VDD2 B 3.634738f
C11 VDD1 B 6.3552f
C12 VTAIL B 4.957462f
C13 VN B 12.02205f
C14 VP B 10.511382f
C15 VDD2.t0 B 0.052402f
C16 VDD2.t3 B 0.052402f
C17 VDD2.n0 B 0.679189f
C18 VDD2.t2 B 0.052402f
C19 VDD2.t1 B 0.052402f
C20 VDD2.n1 B 0.394026f
C21 VDD2.n2 B 2.37676f
C22 VN.t0 B 0.955694f
C23 VN.t3 B 0.967485f
C24 VN.n0 B 0.611282f
C25 VN.t1 B 0.955694f
C26 VN.t2 B 0.967485f
C27 VN.n1 B 1.86201f
C28 VDD1.t1 B 0.051383f
C29 VDD1.t3 B 0.051383f
C30 VDD1.n0 B 0.386666f
C31 VDD1.t2 B 0.051383f
C32 VDD1.t0 B 0.051383f
C33 VDD1.n1 B 0.681923f
C34 VTAIL.n0 B 0.033985f
C35 VTAIL.n1 B 0.025527f
C36 VTAIL.n2 B 0.013717f
C37 VTAIL.n3 B 0.024316f
C38 VTAIL.n4 B 0.018905f
C39 VTAIL.t1 B 0.05447f
C40 VTAIL.n5 B 0.09382f
C41 VTAIL.n6 B 0.271976f
C42 VTAIL.n7 B 0.013717f
C43 VTAIL.n8 B 0.014524f
C44 VTAIL.n9 B 0.032422f
C45 VTAIL.n10 B 0.066837f
C46 VTAIL.n11 B 0.014524f
C47 VTAIL.n12 B 0.013717f
C48 VTAIL.n13 B 0.060747f
C49 VTAIL.n14 B 0.037106f
C50 VTAIL.n15 B 0.210158f
C51 VTAIL.n16 B 0.033985f
C52 VTAIL.n17 B 0.025527f
C53 VTAIL.n18 B 0.013717f
C54 VTAIL.n19 B 0.024316f
C55 VTAIL.n20 B 0.018905f
C56 VTAIL.t7 B 0.05447f
C57 VTAIL.n21 B 0.09382f
C58 VTAIL.n22 B 0.271976f
C59 VTAIL.n23 B 0.013717f
C60 VTAIL.n24 B 0.014524f
C61 VTAIL.n25 B 0.032422f
C62 VTAIL.n26 B 0.066837f
C63 VTAIL.n27 B 0.014524f
C64 VTAIL.n28 B 0.013717f
C65 VTAIL.n29 B 0.060747f
C66 VTAIL.n30 B 0.037106f
C67 VTAIL.n31 B 0.349313f
C68 VTAIL.n32 B 0.033985f
C69 VTAIL.n33 B 0.025527f
C70 VTAIL.n34 B 0.013717f
C71 VTAIL.n35 B 0.024316f
C72 VTAIL.n36 B 0.018905f
C73 VTAIL.t6 B 0.05447f
C74 VTAIL.n37 B 0.09382f
C75 VTAIL.n38 B 0.271976f
C76 VTAIL.n39 B 0.013717f
C77 VTAIL.n40 B 0.014524f
C78 VTAIL.n41 B 0.032422f
C79 VTAIL.n42 B 0.066837f
C80 VTAIL.n43 B 0.014524f
C81 VTAIL.n44 B 0.013717f
C82 VTAIL.n45 B 0.060747f
C83 VTAIL.n46 B 0.037106f
C84 VTAIL.n47 B 1.17007f
C85 VTAIL.n48 B 0.033985f
C86 VTAIL.n49 B 0.025527f
C87 VTAIL.n50 B 0.013717f
C88 VTAIL.n51 B 0.024316f
C89 VTAIL.n52 B 0.018905f
C90 VTAIL.t3 B 0.05447f
C91 VTAIL.n53 B 0.09382f
C92 VTAIL.n54 B 0.271976f
C93 VTAIL.n55 B 0.013717f
C94 VTAIL.n56 B 0.014524f
C95 VTAIL.n57 B 0.032422f
C96 VTAIL.n58 B 0.066837f
C97 VTAIL.n59 B 0.014524f
C98 VTAIL.n60 B 0.013717f
C99 VTAIL.n61 B 0.060747f
C100 VTAIL.n62 B 0.037106f
C101 VTAIL.n63 B 1.17007f
C102 VTAIL.n64 B 0.033985f
C103 VTAIL.n65 B 0.025527f
C104 VTAIL.n66 B 0.013717f
C105 VTAIL.n67 B 0.024316f
C106 VTAIL.n68 B 0.018905f
C107 VTAIL.t0 B 0.05447f
C108 VTAIL.n69 B 0.09382f
C109 VTAIL.n70 B 0.271976f
C110 VTAIL.n71 B 0.013717f
C111 VTAIL.n72 B 0.014524f
C112 VTAIL.n73 B 0.032422f
C113 VTAIL.n74 B 0.066837f
C114 VTAIL.n75 B 0.014524f
C115 VTAIL.n76 B 0.013717f
C116 VTAIL.n77 B 0.060747f
C117 VTAIL.n78 B 0.037106f
C118 VTAIL.n79 B 0.349313f
C119 VTAIL.n80 B 0.033985f
C120 VTAIL.n81 B 0.025527f
C121 VTAIL.n82 B 0.013717f
C122 VTAIL.n83 B 0.024316f
C123 VTAIL.n84 B 0.018905f
C124 VTAIL.t4 B 0.05447f
C125 VTAIL.n85 B 0.09382f
C126 VTAIL.n86 B 0.271976f
C127 VTAIL.n87 B 0.013717f
C128 VTAIL.n88 B 0.014524f
C129 VTAIL.n89 B 0.032422f
C130 VTAIL.n90 B 0.066837f
C131 VTAIL.n91 B 0.014524f
C132 VTAIL.n92 B 0.013717f
C133 VTAIL.n93 B 0.060747f
C134 VTAIL.n94 B 0.037106f
C135 VTAIL.n95 B 0.349313f
C136 VTAIL.n96 B 0.033985f
C137 VTAIL.n97 B 0.025527f
C138 VTAIL.n98 B 0.013717f
C139 VTAIL.n99 B 0.024316f
C140 VTAIL.n100 B 0.018905f
C141 VTAIL.t5 B 0.05447f
C142 VTAIL.n101 B 0.09382f
C143 VTAIL.n102 B 0.271976f
C144 VTAIL.n103 B 0.013717f
C145 VTAIL.n104 B 0.014524f
C146 VTAIL.n105 B 0.032422f
C147 VTAIL.n106 B 0.066837f
C148 VTAIL.n107 B 0.014524f
C149 VTAIL.n108 B 0.013717f
C150 VTAIL.n109 B 0.060747f
C151 VTAIL.n110 B 0.037106f
C152 VTAIL.n111 B 1.17007f
C153 VTAIL.n112 B 0.033985f
C154 VTAIL.n113 B 0.025527f
C155 VTAIL.n114 B 0.013717f
C156 VTAIL.n115 B 0.024316f
C157 VTAIL.n116 B 0.018905f
C158 VTAIL.t2 B 0.05447f
C159 VTAIL.n117 B 0.09382f
C160 VTAIL.n118 B 0.271976f
C161 VTAIL.n119 B 0.013717f
C162 VTAIL.n120 B 0.014524f
C163 VTAIL.n121 B 0.032422f
C164 VTAIL.n122 B 0.066837f
C165 VTAIL.n123 B 0.014524f
C166 VTAIL.n124 B 0.013717f
C167 VTAIL.n125 B 0.060747f
C168 VTAIL.n126 B 0.037106f
C169 VTAIL.n127 B 1.02134f
C170 VP.t3 B 0.683599f
C171 VP.n0 B 0.359195f
C172 VP.n1 B 0.023054f
C173 VP.n2 B 0.045819f
C174 VP.n3 B 0.023054f
C175 VP.n4 B 0.042967f
C176 VP.t2 B 0.971556f
C177 VP.t0 B 0.959716f
C178 VP.n5 B 1.86009f
C179 VP.n6 B 1.14334f
C180 VP.t1 B 0.683599f
C181 VP.n7 B 0.359195f
C182 VP.n8 B 0.023027f
C183 VP.n9 B 0.037209f
C184 VP.n10 B 0.023054f
C185 VP.n11 B 0.023054f
C186 VP.n12 B 0.042967f
C187 VP.n13 B 0.045819f
C188 VP.n14 B 0.018637f
C189 VP.n15 B 0.023054f
C190 VP.n16 B 0.023054f
C191 VP.n17 B 0.023054f
C192 VP.n18 B 0.042967f
C193 VP.n19 B 0.042967f
C194 VP.n20 B 0.023027f
C195 VP.n21 B 0.037209f
C196 VP.n22 B 0.070838f
.ends

