* NGSPICE file created from diff_pair_sample_0564.ext - technology: sky130A

.subckt diff_pair_sample_0564 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=2.2542 ps=12.34 w=5.78 l=0.91
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=0 ps=0 w=5.78 l=0.91
X2 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=2.2542 ps=12.34 w=5.78 l=0.91
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=0 ps=0 w=5.78 l=0.91
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=0 ps=0 w=5.78 l=0.91
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=0 ps=0 w=5.78 l=0.91
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=2.2542 ps=12.34 w=5.78 l=0.91
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2542 pd=12.34 as=2.2542 ps=12.34 w=5.78 l=0.91
R0 VN VN.t0 393.401
R1 VN VN.t1 357.594
R2 VTAIL.n118 VTAIL.n117 289.615
R3 VTAIL.n28 VTAIL.n27 289.615
R4 VTAIL.n88 VTAIL.n87 289.615
R5 VTAIL.n58 VTAIL.n57 289.615
R6 VTAIL.n101 VTAIL.n100 185
R7 VTAIL.n103 VTAIL.n102 185
R8 VTAIL.n96 VTAIL.n95 185
R9 VTAIL.n109 VTAIL.n108 185
R10 VTAIL.n111 VTAIL.n110 185
R11 VTAIL.n92 VTAIL.n91 185
R12 VTAIL.n117 VTAIL.n116 185
R13 VTAIL.n11 VTAIL.n10 185
R14 VTAIL.n13 VTAIL.n12 185
R15 VTAIL.n6 VTAIL.n5 185
R16 VTAIL.n19 VTAIL.n18 185
R17 VTAIL.n21 VTAIL.n20 185
R18 VTAIL.n2 VTAIL.n1 185
R19 VTAIL.n27 VTAIL.n26 185
R20 VTAIL.n87 VTAIL.n86 185
R21 VTAIL.n62 VTAIL.n61 185
R22 VTAIL.n81 VTAIL.n80 185
R23 VTAIL.n79 VTAIL.n78 185
R24 VTAIL.n66 VTAIL.n65 185
R25 VTAIL.n73 VTAIL.n72 185
R26 VTAIL.n71 VTAIL.n70 185
R27 VTAIL.n57 VTAIL.n56 185
R28 VTAIL.n32 VTAIL.n31 185
R29 VTAIL.n51 VTAIL.n50 185
R30 VTAIL.n49 VTAIL.n48 185
R31 VTAIL.n36 VTAIL.n35 185
R32 VTAIL.n43 VTAIL.n42 185
R33 VTAIL.n41 VTAIL.n40 185
R34 VTAIL.n99 VTAIL.t2 149.528
R35 VTAIL.n9 VTAIL.t1 149.528
R36 VTAIL.n69 VTAIL.t0 149.528
R37 VTAIL.n39 VTAIL.t3 149.528
R38 VTAIL.n102 VTAIL.n101 104.615
R39 VTAIL.n102 VTAIL.n95 104.615
R40 VTAIL.n109 VTAIL.n95 104.615
R41 VTAIL.n110 VTAIL.n109 104.615
R42 VTAIL.n110 VTAIL.n91 104.615
R43 VTAIL.n117 VTAIL.n91 104.615
R44 VTAIL.n12 VTAIL.n11 104.615
R45 VTAIL.n12 VTAIL.n5 104.615
R46 VTAIL.n19 VTAIL.n5 104.615
R47 VTAIL.n20 VTAIL.n19 104.615
R48 VTAIL.n20 VTAIL.n1 104.615
R49 VTAIL.n27 VTAIL.n1 104.615
R50 VTAIL.n87 VTAIL.n61 104.615
R51 VTAIL.n80 VTAIL.n61 104.615
R52 VTAIL.n80 VTAIL.n79 104.615
R53 VTAIL.n79 VTAIL.n65 104.615
R54 VTAIL.n72 VTAIL.n65 104.615
R55 VTAIL.n72 VTAIL.n71 104.615
R56 VTAIL.n57 VTAIL.n31 104.615
R57 VTAIL.n50 VTAIL.n31 104.615
R58 VTAIL.n50 VTAIL.n49 104.615
R59 VTAIL.n49 VTAIL.n35 104.615
R60 VTAIL.n42 VTAIL.n35 104.615
R61 VTAIL.n42 VTAIL.n41 104.615
R62 VTAIL.n101 VTAIL.t2 52.3082
R63 VTAIL.n11 VTAIL.t1 52.3082
R64 VTAIL.n71 VTAIL.t0 52.3082
R65 VTAIL.n41 VTAIL.t3 52.3082
R66 VTAIL.n119 VTAIL.n118 33.7369
R67 VTAIL.n29 VTAIL.n28 33.7369
R68 VTAIL.n89 VTAIL.n88 33.7369
R69 VTAIL.n59 VTAIL.n58 33.7369
R70 VTAIL.n59 VTAIL.n29 19.5048
R71 VTAIL.n119 VTAIL.n89 18.4358
R72 VTAIL.n116 VTAIL.n90 12.0247
R73 VTAIL.n26 VTAIL.n0 12.0247
R74 VTAIL.n86 VTAIL.n60 12.0247
R75 VTAIL.n56 VTAIL.n30 12.0247
R76 VTAIL.n115 VTAIL.n92 11.249
R77 VTAIL.n25 VTAIL.n2 11.249
R78 VTAIL.n85 VTAIL.n62 11.249
R79 VTAIL.n55 VTAIL.n32 11.249
R80 VTAIL.n112 VTAIL.n111 10.4732
R81 VTAIL.n22 VTAIL.n21 10.4732
R82 VTAIL.n82 VTAIL.n81 10.4732
R83 VTAIL.n52 VTAIL.n51 10.4732
R84 VTAIL.n100 VTAIL.n99 10.2745
R85 VTAIL.n10 VTAIL.n9 10.2745
R86 VTAIL.n70 VTAIL.n69 10.2745
R87 VTAIL.n40 VTAIL.n39 10.2745
R88 VTAIL.n108 VTAIL.n94 9.69747
R89 VTAIL.n18 VTAIL.n4 9.69747
R90 VTAIL.n78 VTAIL.n64 9.69747
R91 VTAIL.n48 VTAIL.n34 9.69747
R92 VTAIL.n114 VTAIL.n90 9.45567
R93 VTAIL.n24 VTAIL.n0 9.45567
R94 VTAIL.n84 VTAIL.n60 9.45567
R95 VTAIL.n54 VTAIL.n30 9.45567
R96 VTAIL.n98 VTAIL.n97 9.3005
R97 VTAIL.n105 VTAIL.n104 9.3005
R98 VTAIL.n107 VTAIL.n106 9.3005
R99 VTAIL.n94 VTAIL.n93 9.3005
R100 VTAIL.n113 VTAIL.n112 9.3005
R101 VTAIL.n115 VTAIL.n114 9.3005
R102 VTAIL.n8 VTAIL.n7 9.3005
R103 VTAIL.n15 VTAIL.n14 9.3005
R104 VTAIL.n17 VTAIL.n16 9.3005
R105 VTAIL.n4 VTAIL.n3 9.3005
R106 VTAIL.n23 VTAIL.n22 9.3005
R107 VTAIL.n25 VTAIL.n24 9.3005
R108 VTAIL.n85 VTAIL.n84 9.3005
R109 VTAIL.n83 VTAIL.n82 9.3005
R110 VTAIL.n64 VTAIL.n63 9.3005
R111 VTAIL.n77 VTAIL.n76 9.3005
R112 VTAIL.n75 VTAIL.n74 9.3005
R113 VTAIL.n68 VTAIL.n67 9.3005
R114 VTAIL.n45 VTAIL.n44 9.3005
R115 VTAIL.n47 VTAIL.n46 9.3005
R116 VTAIL.n34 VTAIL.n33 9.3005
R117 VTAIL.n53 VTAIL.n52 9.3005
R118 VTAIL.n55 VTAIL.n54 9.3005
R119 VTAIL.n38 VTAIL.n37 9.3005
R120 VTAIL.n107 VTAIL.n96 8.92171
R121 VTAIL.n17 VTAIL.n6 8.92171
R122 VTAIL.n77 VTAIL.n66 8.92171
R123 VTAIL.n47 VTAIL.n36 8.92171
R124 VTAIL.n104 VTAIL.n103 8.14595
R125 VTAIL.n14 VTAIL.n13 8.14595
R126 VTAIL.n74 VTAIL.n73 8.14595
R127 VTAIL.n44 VTAIL.n43 8.14595
R128 VTAIL.n100 VTAIL.n98 7.3702
R129 VTAIL.n10 VTAIL.n8 7.3702
R130 VTAIL.n70 VTAIL.n68 7.3702
R131 VTAIL.n40 VTAIL.n38 7.3702
R132 VTAIL.n103 VTAIL.n98 5.81868
R133 VTAIL.n13 VTAIL.n8 5.81868
R134 VTAIL.n73 VTAIL.n68 5.81868
R135 VTAIL.n43 VTAIL.n38 5.81868
R136 VTAIL.n104 VTAIL.n96 5.04292
R137 VTAIL.n14 VTAIL.n6 5.04292
R138 VTAIL.n74 VTAIL.n66 5.04292
R139 VTAIL.n44 VTAIL.n36 5.04292
R140 VTAIL.n108 VTAIL.n107 4.26717
R141 VTAIL.n18 VTAIL.n17 4.26717
R142 VTAIL.n78 VTAIL.n77 4.26717
R143 VTAIL.n48 VTAIL.n47 4.26717
R144 VTAIL.n111 VTAIL.n94 3.49141
R145 VTAIL.n21 VTAIL.n4 3.49141
R146 VTAIL.n81 VTAIL.n64 3.49141
R147 VTAIL.n51 VTAIL.n34 3.49141
R148 VTAIL.n69 VTAIL.n67 2.84323
R149 VTAIL.n39 VTAIL.n37 2.84323
R150 VTAIL.n99 VTAIL.n97 2.84323
R151 VTAIL.n9 VTAIL.n7 2.84323
R152 VTAIL.n112 VTAIL.n92 2.71565
R153 VTAIL.n22 VTAIL.n2 2.71565
R154 VTAIL.n82 VTAIL.n62 2.71565
R155 VTAIL.n52 VTAIL.n32 2.71565
R156 VTAIL.n116 VTAIL.n115 1.93989
R157 VTAIL.n26 VTAIL.n25 1.93989
R158 VTAIL.n86 VTAIL.n85 1.93989
R159 VTAIL.n56 VTAIL.n55 1.93989
R160 VTAIL.n118 VTAIL.n90 1.16414
R161 VTAIL.n28 VTAIL.n0 1.16414
R162 VTAIL.n88 VTAIL.n60 1.16414
R163 VTAIL.n58 VTAIL.n30 1.16414
R164 VTAIL.n89 VTAIL.n59 1.00481
R165 VTAIL VTAIL.n29 0.795759
R166 VTAIL VTAIL.n119 0.209552
R167 VTAIL.n105 VTAIL.n97 0.155672
R168 VTAIL.n106 VTAIL.n105 0.155672
R169 VTAIL.n106 VTAIL.n93 0.155672
R170 VTAIL.n113 VTAIL.n93 0.155672
R171 VTAIL.n114 VTAIL.n113 0.155672
R172 VTAIL.n15 VTAIL.n7 0.155672
R173 VTAIL.n16 VTAIL.n15 0.155672
R174 VTAIL.n16 VTAIL.n3 0.155672
R175 VTAIL.n23 VTAIL.n3 0.155672
R176 VTAIL.n24 VTAIL.n23 0.155672
R177 VTAIL.n84 VTAIL.n83 0.155672
R178 VTAIL.n83 VTAIL.n63 0.155672
R179 VTAIL.n76 VTAIL.n63 0.155672
R180 VTAIL.n76 VTAIL.n75 0.155672
R181 VTAIL.n75 VTAIL.n67 0.155672
R182 VTAIL.n54 VTAIL.n53 0.155672
R183 VTAIL.n53 VTAIL.n33 0.155672
R184 VTAIL.n46 VTAIL.n33 0.155672
R185 VTAIL.n46 VTAIL.n45 0.155672
R186 VTAIL.n45 VTAIL.n37 0.155672
R187 VDD2.n57 VDD2.n56 289.615
R188 VDD2.n28 VDD2.n27 289.615
R189 VDD2.n56 VDD2.n55 185
R190 VDD2.n31 VDD2.n30 185
R191 VDD2.n50 VDD2.n49 185
R192 VDD2.n48 VDD2.n47 185
R193 VDD2.n35 VDD2.n34 185
R194 VDD2.n42 VDD2.n41 185
R195 VDD2.n40 VDD2.n39 185
R196 VDD2.n11 VDD2.n10 185
R197 VDD2.n13 VDD2.n12 185
R198 VDD2.n6 VDD2.n5 185
R199 VDD2.n19 VDD2.n18 185
R200 VDD2.n21 VDD2.n20 185
R201 VDD2.n2 VDD2.n1 185
R202 VDD2.n27 VDD2.n26 185
R203 VDD2.n38 VDD2.t1 149.528
R204 VDD2.n9 VDD2.t0 149.528
R205 VDD2.n56 VDD2.n30 104.615
R206 VDD2.n49 VDD2.n30 104.615
R207 VDD2.n49 VDD2.n48 104.615
R208 VDD2.n48 VDD2.n34 104.615
R209 VDD2.n41 VDD2.n34 104.615
R210 VDD2.n41 VDD2.n40 104.615
R211 VDD2.n12 VDD2.n11 104.615
R212 VDD2.n12 VDD2.n5 104.615
R213 VDD2.n19 VDD2.n5 104.615
R214 VDD2.n20 VDD2.n19 104.615
R215 VDD2.n20 VDD2.n1 104.615
R216 VDD2.n27 VDD2.n1 104.615
R217 VDD2.n58 VDD2.n28 81.213
R218 VDD2.n40 VDD2.t1 52.3082
R219 VDD2.n11 VDD2.t0 52.3082
R220 VDD2.n58 VDD2.n57 50.4157
R221 VDD2.n55 VDD2.n29 12.0247
R222 VDD2.n26 VDD2.n0 12.0247
R223 VDD2.n54 VDD2.n31 11.249
R224 VDD2.n25 VDD2.n2 11.249
R225 VDD2.n51 VDD2.n50 10.4732
R226 VDD2.n22 VDD2.n21 10.4732
R227 VDD2.n39 VDD2.n38 10.2745
R228 VDD2.n10 VDD2.n9 10.2745
R229 VDD2.n47 VDD2.n33 9.69747
R230 VDD2.n18 VDD2.n4 9.69747
R231 VDD2.n53 VDD2.n29 9.45567
R232 VDD2.n24 VDD2.n0 9.45567
R233 VDD2.n54 VDD2.n53 9.3005
R234 VDD2.n52 VDD2.n51 9.3005
R235 VDD2.n33 VDD2.n32 9.3005
R236 VDD2.n46 VDD2.n45 9.3005
R237 VDD2.n44 VDD2.n43 9.3005
R238 VDD2.n37 VDD2.n36 9.3005
R239 VDD2.n8 VDD2.n7 9.3005
R240 VDD2.n15 VDD2.n14 9.3005
R241 VDD2.n17 VDD2.n16 9.3005
R242 VDD2.n4 VDD2.n3 9.3005
R243 VDD2.n23 VDD2.n22 9.3005
R244 VDD2.n25 VDD2.n24 9.3005
R245 VDD2.n46 VDD2.n35 8.92171
R246 VDD2.n17 VDD2.n6 8.92171
R247 VDD2.n43 VDD2.n42 8.14595
R248 VDD2.n14 VDD2.n13 8.14595
R249 VDD2.n39 VDD2.n37 7.3702
R250 VDD2.n10 VDD2.n8 7.3702
R251 VDD2.n42 VDD2.n37 5.81868
R252 VDD2.n13 VDD2.n8 5.81868
R253 VDD2.n43 VDD2.n35 5.04292
R254 VDD2.n14 VDD2.n6 5.04292
R255 VDD2.n47 VDD2.n46 4.26717
R256 VDD2.n18 VDD2.n17 4.26717
R257 VDD2.n50 VDD2.n33 3.49141
R258 VDD2.n21 VDD2.n4 3.49141
R259 VDD2.n38 VDD2.n36 2.84323
R260 VDD2.n9 VDD2.n7 2.84323
R261 VDD2.n51 VDD2.n31 2.71565
R262 VDD2.n22 VDD2.n2 2.71565
R263 VDD2.n55 VDD2.n54 1.93989
R264 VDD2.n26 VDD2.n25 1.93989
R265 VDD2.n57 VDD2.n29 1.16414
R266 VDD2.n28 VDD2.n0 1.16414
R267 VDD2 VDD2.n58 0.325931
R268 VDD2.n53 VDD2.n52 0.155672
R269 VDD2.n52 VDD2.n32 0.155672
R270 VDD2.n45 VDD2.n32 0.155672
R271 VDD2.n45 VDD2.n44 0.155672
R272 VDD2.n44 VDD2.n36 0.155672
R273 VDD2.n15 VDD2.n7 0.155672
R274 VDD2.n16 VDD2.n15 0.155672
R275 VDD2.n16 VDD2.n3 0.155672
R276 VDD2.n23 VDD2.n3 0.155672
R277 VDD2.n24 VDD2.n23 0.155672
R278 B.n413 B.n412 585
R279 B.n172 B.n60 585
R280 B.n171 B.n170 585
R281 B.n169 B.n168 585
R282 B.n167 B.n166 585
R283 B.n165 B.n164 585
R284 B.n163 B.n162 585
R285 B.n161 B.n160 585
R286 B.n159 B.n158 585
R287 B.n157 B.n156 585
R288 B.n155 B.n154 585
R289 B.n153 B.n152 585
R290 B.n151 B.n150 585
R291 B.n149 B.n148 585
R292 B.n147 B.n146 585
R293 B.n145 B.n144 585
R294 B.n143 B.n142 585
R295 B.n141 B.n140 585
R296 B.n139 B.n138 585
R297 B.n137 B.n136 585
R298 B.n135 B.n134 585
R299 B.n133 B.n132 585
R300 B.n131 B.n130 585
R301 B.n128 B.n127 585
R302 B.n126 B.n125 585
R303 B.n124 B.n123 585
R304 B.n122 B.n121 585
R305 B.n120 B.n119 585
R306 B.n118 B.n117 585
R307 B.n116 B.n115 585
R308 B.n114 B.n113 585
R309 B.n112 B.n111 585
R310 B.n110 B.n109 585
R311 B.n107 B.n106 585
R312 B.n105 B.n104 585
R313 B.n103 B.n102 585
R314 B.n101 B.n100 585
R315 B.n99 B.n98 585
R316 B.n97 B.n96 585
R317 B.n95 B.n94 585
R318 B.n93 B.n92 585
R319 B.n91 B.n90 585
R320 B.n89 B.n88 585
R321 B.n87 B.n86 585
R322 B.n85 B.n84 585
R323 B.n83 B.n82 585
R324 B.n81 B.n80 585
R325 B.n79 B.n78 585
R326 B.n77 B.n76 585
R327 B.n75 B.n74 585
R328 B.n73 B.n72 585
R329 B.n71 B.n70 585
R330 B.n69 B.n68 585
R331 B.n67 B.n66 585
R332 B.n33 B.n32 585
R333 B.n418 B.n417 585
R334 B.n411 B.n61 585
R335 B.n61 B.n30 585
R336 B.n410 B.n29 585
R337 B.n422 B.n29 585
R338 B.n409 B.n28 585
R339 B.n423 B.n28 585
R340 B.n408 B.n27 585
R341 B.n424 B.n27 585
R342 B.n407 B.n406 585
R343 B.n406 B.n23 585
R344 B.n405 B.n22 585
R345 B.n430 B.n22 585
R346 B.n404 B.n21 585
R347 B.n431 B.n21 585
R348 B.n403 B.n20 585
R349 B.n432 B.n20 585
R350 B.n402 B.n401 585
R351 B.n401 B.n16 585
R352 B.n400 B.n15 585
R353 B.n438 B.n15 585
R354 B.n399 B.n14 585
R355 B.n439 B.n14 585
R356 B.n398 B.n13 585
R357 B.n440 B.n13 585
R358 B.n397 B.n396 585
R359 B.n396 B.n12 585
R360 B.n395 B.n394 585
R361 B.n395 B.n8 585
R362 B.n393 B.n7 585
R363 B.n447 B.n7 585
R364 B.n392 B.n6 585
R365 B.n448 B.n6 585
R366 B.n391 B.n5 585
R367 B.n449 B.n5 585
R368 B.n390 B.n389 585
R369 B.n389 B.n4 585
R370 B.n388 B.n173 585
R371 B.n388 B.n387 585
R372 B.n377 B.n174 585
R373 B.n380 B.n174 585
R374 B.n379 B.n378 585
R375 B.n381 B.n379 585
R376 B.n376 B.n179 585
R377 B.n179 B.n178 585
R378 B.n375 B.n374 585
R379 B.n374 B.n373 585
R380 B.n181 B.n180 585
R381 B.n182 B.n181 585
R382 B.n366 B.n365 585
R383 B.n367 B.n366 585
R384 B.n364 B.n187 585
R385 B.n187 B.n186 585
R386 B.n363 B.n362 585
R387 B.n362 B.n361 585
R388 B.n189 B.n188 585
R389 B.n190 B.n189 585
R390 B.n354 B.n353 585
R391 B.n355 B.n354 585
R392 B.n352 B.n195 585
R393 B.n195 B.n194 585
R394 B.n351 B.n350 585
R395 B.n350 B.n349 585
R396 B.n197 B.n196 585
R397 B.n198 B.n197 585
R398 B.n345 B.n344 585
R399 B.n201 B.n200 585
R400 B.n341 B.n340 585
R401 B.n342 B.n341 585
R402 B.n339 B.n229 585
R403 B.n338 B.n337 585
R404 B.n336 B.n335 585
R405 B.n334 B.n333 585
R406 B.n332 B.n331 585
R407 B.n330 B.n329 585
R408 B.n328 B.n327 585
R409 B.n326 B.n325 585
R410 B.n324 B.n323 585
R411 B.n322 B.n321 585
R412 B.n320 B.n319 585
R413 B.n318 B.n317 585
R414 B.n316 B.n315 585
R415 B.n314 B.n313 585
R416 B.n312 B.n311 585
R417 B.n310 B.n309 585
R418 B.n308 B.n307 585
R419 B.n306 B.n305 585
R420 B.n304 B.n303 585
R421 B.n302 B.n301 585
R422 B.n300 B.n299 585
R423 B.n298 B.n297 585
R424 B.n296 B.n295 585
R425 B.n294 B.n293 585
R426 B.n292 B.n291 585
R427 B.n290 B.n289 585
R428 B.n288 B.n287 585
R429 B.n286 B.n285 585
R430 B.n284 B.n283 585
R431 B.n282 B.n281 585
R432 B.n280 B.n279 585
R433 B.n278 B.n277 585
R434 B.n276 B.n275 585
R435 B.n274 B.n273 585
R436 B.n272 B.n271 585
R437 B.n270 B.n269 585
R438 B.n268 B.n267 585
R439 B.n266 B.n265 585
R440 B.n264 B.n263 585
R441 B.n262 B.n261 585
R442 B.n260 B.n259 585
R443 B.n258 B.n257 585
R444 B.n256 B.n255 585
R445 B.n254 B.n253 585
R446 B.n252 B.n251 585
R447 B.n250 B.n249 585
R448 B.n248 B.n247 585
R449 B.n246 B.n245 585
R450 B.n244 B.n243 585
R451 B.n242 B.n241 585
R452 B.n240 B.n239 585
R453 B.n238 B.n237 585
R454 B.n236 B.n228 585
R455 B.n342 B.n228 585
R456 B.n346 B.n199 585
R457 B.n199 B.n198 585
R458 B.n348 B.n347 585
R459 B.n349 B.n348 585
R460 B.n193 B.n192 585
R461 B.n194 B.n193 585
R462 B.n357 B.n356 585
R463 B.n356 B.n355 585
R464 B.n358 B.n191 585
R465 B.n191 B.n190 585
R466 B.n360 B.n359 585
R467 B.n361 B.n360 585
R468 B.n185 B.n184 585
R469 B.n186 B.n185 585
R470 B.n369 B.n368 585
R471 B.n368 B.n367 585
R472 B.n370 B.n183 585
R473 B.n183 B.n182 585
R474 B.n372 B.n371 585
R475 B.n373 B.n372 585
R476 B.n177 B.n176 585
R477 B.n178 B.n177 585
R478 B.n383 B.n382 585
R479 B.n382 B.n381 585
R480 B.n384 B.n175 585
R481 B.n380 B.n175 585
R482 B.n386 B.n385 585
R483 B.n387 B.n386 585
R484 B.n3 B.n0 585
R485 B.n4 B.n3 585
R486 B.n446 B.n1 585
R487 B.n447 B.n446 585
R488 B.n445 B.n444 585
R489 B.n445 B.n8 585
R490 B.n443 B.n9 585
R491 B.n12 B.n9 585
R492 B.n442 B.n441 585
R493 B.n441 B.n440 585
R494 B.n11 B.n10 585
R495 B.n439 B.n11 585
R496 B.n437 B.n436 585
R497 B.n438 B.n437 585
R498 B.n435 B.n17 585
R499 B.n17 B.n16 585
R500 B.n434 B.n433 585
R501 B.n433 B.n432 585
R502 B.n19 B.n18 585
R503 B.n431 B.n19 585
R504 B.n429 B.n428 585
R505 B.n430 B.n429 585
R506 B.n427 B.n24 585
R507 B.n24 B.n23 585
R508 B.n426 B.n425 585
R509 B.n425 B.n424 585
R510 B.n26 B.n25 585
R511 B.n423 B.n26 585
R512 B.n421 B.n420 585
R513 B.n422 B.n421 585
R514 B.n419 B.n31 585
R515 B.n31 B.n30 585
R516 B.n450 B.n449 585
R517 B.n448 B.n2 585
R518 B.n417 B.n31 511.721
R519 B.n413 B.n61 511.721
R520 B.n228 B.n197 511.721
R521 B.n344 B.n199 511.721
R522 B.n64 B.t6 355.349
R523 B.n62 B.t13 355.349
R524 B.n233 B.t10 355.349
R525 B.n230 B.t2 355.349
R526 B.n415 B.n414 256.663
R527 B.n415 B.n59 256.663
R528 B.n415 B.n58 256.663
R529 B.n415 B.n57 256.663
R530 B.n415 B.n56 256.663
R531 B.n415 B.n55 256.663
R532 B.n415 B.n54 256.663
R533 B.n415 B.n53 256.663
R534 B.n415 B.n52 256.663
R535 B.n415 B.n51 256.663
R536 B.n415 B.n50 256.663
R537 B.n415 B.n49 256.663
R538 B.n415 B.n48 256.663
R539 B.n415 B.n47 256.663
R540 B.n415 B.n46 256.663
R541 B.n415 B.n45 256.663
R542 B.n415 B.n44 256.663
R543 B.n415 B.n43 256.663
R544 B.n415 B.n42 256.663
R545 B.n415 B.n41 256.663
R546 B.n415 B.n40 256.663
R547 B.n415 B.n39 256.663
R548 B.n415 B.n38 256.663
R549 B.n415 B.n37 256.663
R550 B.n415 B.n36 256.663
R551 B.n415 B.n35 256.663
R552 B.n415 B.n34 256.663
R553 B.n416 B.n415 256.663
R554 B.n343 B.n342 256.663
R555 B.n342 B.n202 256.663
R556 B.n342 B.n203 256.663
R557 B.n342 B.n204 256.663
R558 B.n342 B.n205 256.663
R559 B.n342 B.n206 256.663
R560 B.n342 B.n207 256.663
R561 B.n342 B.n208 256.663
R562 B.n342 B.n209 256.663
R563 B.n342 B.n210 256.663
R564 B.n342 B.n211 256.663
R565 B.n342 B.n212 256.663
R566 B.n342 B.n213 256.663
R567 B.n342 B.n214 256.663
R568 B.n342 B.n215 256.663
R569 B.n342 B.n216 256.663
R570 B.n342 B.n217 256.663
R571 B.n342 B.n218 256.663
R572 B.n342 B.n219 256.663
R573 B.n342 B.n220 256.663
R574 B.n342 B.n221 256.663
R575 B.n342 B.n222 256.663
R576 B.n342 B.n223 256.663
R577 B.n342 B.n224 256.663
R578 B.n342 B.n225 256.663
R579 B.n342 B.n226 256.663
R580 B.n342 B.n227 256.663
R581 B.n452 B.n451 256.663
R582 B.n62 B.t14 198.768
R583 B.n233 B.t12 198.768
R584 B.n64 B.t8 198.768
R585 B.n230 B.t5 198.768
R586 B.n63 B.t15 174.72
R587 B.n234 B.t11 174.72
R588 B.n65 B.t9 174.72
R589 B.n231 B.t4 174.72
R590 B.n66 B.n33 163.367
R591 B.n70 B.n69 163.367
R592 B.n74 B.n73 163.367
R593 B.n78 B.n77 163.367
R594 B.n82 B.n81 163.367
R595 B.n86 B.n85 163.367
R596 B.n90 B.n89 163.367
R597 B.n94 B.n93 163.367
R598 B.n98 B.n97 163.367
R599 B.n102 B.n101 163.367
R600 B.n106 B.n105 163.367
R601 B.n111 B.n110 163.367
R602 B.n115 B.n114 163.367
R603 B.n119 B.n118 163.367
R604 B.n123 B.n122 163.367
R605 B.n127 B.n126 163.367
R606 B.n132 B.n131 163.367
R607 B.n136 B.n135 163.367
R608 B.n140 B.n139 163.367
R609 B.n144 B.n143 163.367
R610 B.n148 B.n147 163.367
R611 B.n152 B.n151 163.367
R612 B.n156 B.n155 163.367
R613 B.n160 B.n159 163.367
R614 B.n164 B.n163 163.367
R615 B.n168 B.n167 163.367
R616 B.n170 B.n60 163.367
R617 B.n350 B.n197 163.367
R618 B.n350 B.n195 163.367
R619 B.n354 B.n195 163.367
R620 B.n354 B.n189 163.367
R621 B.n362 B.n189 163.367
R622 B.n362 B.n187 163.367
R623 B.n366 B.n187 163.367
R624 B.n366 B.n181 163.367
R625 B.n374 B.n181 163.367
R626 B.n374 B.n179 163.367
R627 B.n379 B.n179 163.367
R628 B.n379 B.n174 163.367
R629 B.n388 B.n174 163.367
R630 B.n389 B.n388 163.367
R631 B.n389 B.n5 163.367
R632 B.n6 B.n5 163.367
R633 B.n7 B.n6 163.367
R634 B.n395 B.n7 163.367
R635 B.n396 B.n395 163.367
R636 B.n396 B.n13 163.367
R637 B.n14 B.n13 163.367
R638 B.n15 B.n14 163.367
R639 B.n401 B.n15 163.367
R640 B.n401 B.n20 163.367
R641 B.n21 B.n20 163.367
R642 B.n22 B.n21 163.367
R643 B.n406 B.n22 163.367
R644 B.n406 B.n27 163.367
R645 B.n28 B.n27 163.367
R646 B.n29 B.n28 163.367
R647 B.n61 B.n29 163.367
R648 B.n341 B.n201 163.367
R649 B.n341 B.n229 163.367
R650 B.n337 B.n336 163.367
R651 B.n333 B.n332 163.367
R652 B.n329 B.n328 163.367
R653 B.n325 B.n324 163.367
R654 B.n321 B.n320 163.367
R655 B.n317 B.n316 163.367
R656 B.n313 B.n312 163.367
R657 B.n309 B.n308 163.367
R658 B.n305 B.n304 163.367
R659 B.n301 B.n300 163.367
R660 B.n297 B.n296 163.367
R661 B.n293 B.n292 163.367
R662 B.n289 B.n288 163.367
R663 B.n285 B.n284 163.367
R664 B.n281 B.n280 163.367
R665 B.n277 B.n276 163.367
R666 B.n273 B.n272 163.367
R667 B.n269 B.n268 163.367
R668 B.n265 B.n264 163.367
R669 B.n261 B.n260 163.367
R670 B.n257 B.n256 163.367
R671 B.n253 B.n252 163.367
R672 B.n249 B.n248 163.367
R673 B.n245 B.n244 163.367
R674 B.n241 B.n240 163.367
R675 B.n237 B.n228 163.367
R676 B.n348 B.n199 163.367
R677 B.n348 B.n193 163.367
R678 B.n356 B.n193 163.367
R679 B.n356 B.n191 163.367
R680 B.n360 B.n191 163.367
R681 B.n360 B.n185 163.367
R682 B.n368 B.n185 163.367
R683 B.n368 B.n183 163.367
R684 B.n372 B.n183 163.367
R685 B.n372 B.n177 163.367
R686 B.n382 B.n177 163.367
R687 B.n382 B.n175 163.367
R688 B.n386 B.n175 163.367
R689 B.n386 B.n3 163.367
R690 B.n450 B.n3 163.367
R691 B.n446 B.n2 163.367
R692 B.n446 B.n445 163.367
R693 B.n445 B.n9 163.367
R694 B.n441 B.n9 163.367
R695 B.n441 B.n11 163.367
R696 B.n437 B.n11 163.367
R697 B.n437 B.n17 163.367
R698 B.n433 B.n17 163.367
R699 B.n433 B.n19 163.367
R700 B.n429 B.n19 163.367
R701 B.n429 B.n24 163.367
R702 B.n425 B.n24 163.367
R703 B.n425 B.n26 163.367
R704 B.n421 B.n26 163.367
R705 B.n421 B.n31 163.367
R706 B.n342 B.n198 116.209
R707 B.n415 B.n30 116.209
R708 B.n417 B.n416 71.676
R709 B.n66 B.n34 71.676
R710 B.n70 B.n35 71.676
R711 B.n74 B.n36 71.676
R712 B.n78 B.n37 71.676
R713 B.n82 B.n38 71.676
R714 B.n86 B.n39 71.676
R715 B.n90 B.n40 71.676
R716 B.n94 B.n41 71.676
R717 B.n98 B.n42 71.676
R718 B.n102 B.n43 71.676
R719 B.n106 B.n44 71.676
R720 B.n111 B.n45 71.676
R721 B.n115 B.n46 71.676
R722 B.n119 B.n47 71.676
R723 B.n123 B.n48 71.676
R724 B.n127 B.n49 71.676
R725 B.n132 B.n50 71.676
R726 B.n136 B.n51 71.676
R727 B.n140 B.n52 71.676
R728 B.n144 B.n53 71.676
R729 B.n148 B.n54 71.676
R730 B.n152 B.n55 71.676
R731 B.n156 B.n56 71.676
R732 B.n160 B.n57 71.676
R733 B.n164 B.n58 71.676
R734 B.n168 B.n59 71.676
R735 B.n414 B.n60 71.676
R736 B.n414 B.n413 71.676
R737 B.n170 B.n59 71.676
R738 B.n167 B.n58 71.676
R739 B.n163 B.n57 71.676
R740 B.n159 B.n56 71.676
R741 B.n155 B.n55 71.676
R742 B.n151 B.n54 71.676
R743 B.n147 B.n53 71.676
R744 B.n143 B.n52 71.676
R745 B.n139 B.n51 71.676
R746 B.n135 B.n50 71.676
R747 B.n131 B.n49 71.676
R748 B.n126 B.n48 71.676
R749 B.n122 B.n47 71.676
R750 B.n118 B.n46 71.676
R751 B.n114 B.n45 71.676
R752 B.n110 B.n44 71.676
R753 B.n105 B.n43 71.676
R754 B.n101 B.n42 71.676
R755 B.n97 B.n41 71.676
R756 B.n93 B.n40 71.676
R757 B.n89 B.n39 71.676
R758 B.n85 B.n38 71.676
R759 B.n81 B.n37 71.676
R760 B.n77 B.n36 71.676
R761 B.n73 B.n35 71.676
R762 B.n69 B.n34 71.676
R763 B.n416 B.n33 71.676
R764 B.n344 B.n343 71.676
R765 B.n229 B.n202 71.676
R766 B.n336 B.n203 71.676
R767 B.n332 B.n204 71.676
R768 B.n328 B.n205 71.676
R769 B.n324 B.n206 71.676
R770 B.n320 B.n207 71.676
R771 B.n316 B.n208 71.676
R772 B.n312 B.n209 71.676
R773 B.n308 B.n210 71.676
R774 B.n304 B.n211 71.676
R775 B.n300 B.n212 71.676
R776 B.n296 B.n213 71.676
R777 B.n292 B.n214 71.676
R778 B.n288 B.n215 71.676
R779 B.n284 B.n216 71.676
R780 B.n280 B.n217 71.676
R781 B.n276 B.n218 71.676
R782 B.n272 B.n219 71.676
R783 B.n268 B.n220 71.676
R784 B.n264 B.n221 71.676
R785 B.n260 B.n222 71.676
R786 B.n256 B.n223 71.676
R787 B.n252 B.n224 71.676
R788 B.n248 B.n225 71.676
R789 B.n244 B.n226 71.676
R790 B.n240 B.n227 71.676
R791 B.n343 B.n201 71.676
R792 B.n337 B.n202 71.676
R793 B.n333 B.n203 71.676
R794 B.n329 B.n204 71.676
R795 B.n325 B.n205 71.676
R796 B.n321 B.n206 71.676
R797 B.n317 B.n207 71.676
R798 B.n313 B.n208 71.676
R799 B.n309 B.n209 71.676
R800 B.n305 B.n210 71.676
R801 B.n301 B.n211 71.676
R802 B.n297 B.n212 71.676
R803 B.n293 B.n213 71.676
R804 B.n289 B.n214 71.676
R805 B.n285 B.n215 71.676
R806 B.n281 B.n216 71.676
R807 B.n277 B.n217 71.676
R808 B.n273 B.n218 71.676
R809 B.n269 B.n219 71.676
R810 B.n265 B.n220 71.676
R811 B.n261 B.n221 71.676
R812 B.n257 B.n222 71.676
R813 B.n253 B.n223 71.676
R814 B.n249 B.n224 71.676
R815 B.n245 B.n225 71.676
R816 B.n241 B.n226 71.676
R817 B.n237 B.n227 71.676
R818 B.n451 B.n450 71.676
R819 B.n451 B.n2 71.676
R820 B.n349 B.n198 67.54
R821 B.n349 B.n194 67.54
R822 B.n355 B.n194 67.54
R823 B.n355 B.n190 67.54
R824 B.n361 B.n190 67.54
R825 B.n367 B.n186 67.54
R826 B.n367 B.n182 67.54
R827 B.n373 B.n182 67.54
R828 B.n373 B.n178 67.54
R829 B.n381 B.n178 67.54
R830 B.n381 B.n380 67.54
R831 B.n387 B.n4 67.54
R832 B.n449 B.n4 67.54
R833 B.n449 B.n448 67.54
R834 B.n448 B.n447 67.54
R835 B.n447 B.n8 67.54
R836 B.n440 B.n12 67.54
R837 B.n440 B.n439 67.54
R838 B.n439 B.n438 67.54
R839 B.n438 B.n16 67.54
R840 B.n432 B.n16 67.54
R841 B.n432 B.n431 67.54
R842 B.n430 B.n23 67.54
R843 B.n424 B.n23 67.54
R844 B.n424 B.n423 67.54
R845 B.n423 B.n422 67.54
R846 B.n422 B.n30 67.54
R847 B.n387 B.t1 62.5739
R848 B.t0 B.n8 62.5739
R849 B.n108 B.n65 59.5399
R850 B.n129 B.n63 59.5399
R851 B.n235 B.n234 59.5399
R852 B.n232 B.n231 59.5399
R853 B.t3 B.n186 52.6416
R854 B.n431 B.t7 52.6416
R855 B.n346 B.n345 33.2493
R856 B.n236 B.n196 33.2493
R857 B.n412 B.n411 33.2493
R858 B.n419 B.n418 33.2493
R859 B.n65 B.n64 24.049
R860 B.n63 B.n62 24.049
R861 B.n234 B.n233 24.049
R862 B.n231 B.n230 24.049
R863 B B.n452 18.0485
R864 B.n361 B.t3 14.8989
R865 B.t7 B.n430 14.8989
R866 B.n347 B.n346 10.6151
R867 B.n347 B.n192 10.6151
R868 B.n357 B.n192 10.6151
R869 B.n358 B.n357 10.6151
R870 B.n359 B.n358 10.6151
R871 B.n359 B.n184 10.6151
R872 B.n369 B.n184 10.6151
R873 B.n370 B.n369 10.6151
R874 B.n371 B.n370 10.6151
R875 B.n371 B.n176 10.6151
R876 B.n383 B.n176 10.6151
R877 B.n384 B.n383 10.6151
R878 B.n385 B.n384 10.6151
R879 B.n385 B.n0 10.6151
R880 B.n345 B.n200 10.6151
R881 B.n340 B.n200 10.6151
R882 B.n340 B.n339 10.6151
R883 B.n339 B.n338 10.6151
R884 B.n338 B.n335 10.6151
R885 B.n335 B.n334 10.6151
R886 B.n334 B.n331 10.6151
R887 B.n331 B.n330 10.6151
R888 B.n330 B.n327 10.6151
R889 B.n327 B.n326 10.6151
R890 B.n326 B.n323 10.6151
R891 B.n323 B.n322 10.6151
R892 B.n322 B.n319 10.6151
R893 B.n319 B.n318 10.6151
R894 B.n318 B.n315 10.6151
R895 B.n315 B.n314 10.6151
R896 B.n314 B.n311 10.6151
R897 B.n311 B.n310 10.6151
R898 B.n310 B.n307 10.6151
R899 B.n307 B.n306 10.6151
R900 B.n306 B.n303 10.6151
R901 B.n303 B.n302 10.6151
R902 B.n299 B.n298 10.6151
R903 B.n298 B.n295 10.6151
R904 B.n295 B.n294 10.6151
R905 B.n294 B.n291 10.6151
R906 B.n291 B.n290 10.6151
R907 B.n290 B.n287 10.6151
R908 B.n287 B.n286 10.6151
R909 B.n286 B.n283 10.6151
R910 B.n283 B.n282 10.6151
R911 B.n279 B.n278 10.6151
R912 B.n278 B.n275 10.6151
R913 B.n275 B.n274 10.6151
R914 B.n274 B.n271 10.6151
R915 B.n271 B.n270 10.6151
R916 B.n270 B.n267 10.6151
R917 B.n267 B.n266 10.6151
R918 B.n266 B.n263 10.6151
R919 B.n263 B.n262 10.6151
R920 B.n262 B.n259 10.6151
R921 B.n259 B.n258 10.6151
R922 B.n258 B.n255 10.6151
R923 B.n255 B.n254 10.6151
R924 B.n254 B.n251 10.6151
R925 B.n251 B.n250 10.6151
R926 B.n250 B.n247 10.6151
R927 B.n247 B.n246 10.6151
R928 B.n246 B.n243 10.6151
R929 B.n243 B.n242 10.6151
R930 B.n242 B.n239 10.6151
R931 B.n239 B.n238 10.6151
R932 B.n238 B.n236 10.6151
R933 B.n351 B.n196 10.6151
R934 B.n352 B.n351 10.6151
R935 B.n353 B.n352 10.6151
R936 B.n353 B.n188 10.6151
R937 B.n363 B.n188 10.6151
R938 B.n364 B.n363 10.6151
R939 B.n365 B.n364 10.6151
R940 B.n365 B.n180 10.6151
R941 B.n375 B.n180 10.6151
R942 B.n376 B.n375 10.6151
R943 B.n378 B.n376 10.6151
R944 B.n378 B.n377 10.6151
R945 B.n377 B.n173 10.6151
R946 B.n390 B.n173 10.6151
R947 B.n391 B.n390 10.6151
R948 B.n392 B.n391 10.6151
R949 B.n393 B.n392 10.6151
R950 B.n394 B.n393 10.6151
R951 B.n397 B.n394 10.6151
R952 B.n398 B.n397 10.6151
R953 B.n399 B.n398 10.6151
R954 B.n400 B.n399 10.6151
R955 B.n402 B.n400 10.6151
R956 B.n403 B.n402 10.6151
R957 B.n404 B.n403 10.6151
R958 B.n405 B.n404 10.6151
R959 B.n407 B.n405 10.6151
R960 B.n408 B.n407 10.6151
R961 B.n409 B.n408 10.6151
R962 B.n410 B.n409 10.6151
R963 B.n411 B.n410 10.6151
R964 B.n444 B.n1 10.6151
R965 B.n444 B.n443 10.6151
R966 B.n443 B.n442 10.6151
R967 B.n442 B.n10 10.6151
R968 B.n436 B.n10 10.6151
R969 B.n436 B.n435 10.6151
R970 B.n435 B.n434 10.6151
R971 B.n434 B.n18 10.6151
R972 B.n428 B.n18 10.6151
R973 B.n428 B.n427 10.6151
R974 B.n427 B.n426 10.6151
R975 B.n426 B.n25 10.6151
R976 B.n420 B.n25 10.6151
R977 B.n420 B.n419 10.6151
R978 B.n418 B.n32 10.6151
R979 B.n67 B.n32 10.6151
R980 B.n68 B.n67 10.6151
R981 B.n71 B.n68 10.6151
R982 B.n72 B.n71 10.6151
R983 B.n75 B.n72 10.6151
R984 B.n76 B.n75 10.6151
R985 B.n79 B.n76 10.6151
R986 B.n80 B.n79 10.6151
R987 B.n83 B.n80 10.6151
R988 B.n84 B.n83 10.6151
R989 B.n87 B.n84 10.6151
R990 B.n88 B.n87 10.6151
R991 B.n91 B.n88 10.6151
R992 B.n92 B.n91 10.6151
R993 B.n95 B.n92 10.6151
R994 B.n96 B.n95 10.6151
R995 B.n99 B.n96 10.6151
R996 B.n100 B.n99 10.6151
R997 B.n103 B.n100 10.6151
R998 B.n104 B.n103 10.6151
R999 B.n107 B.n104 10.6151
R1000 B.n112 B.n109 10.6151
R1001 B.n113 B.n112 10.6151
R1002 B.n116 B.n113 10.6151
R1003 B.n117 B.n116 10.6151
R1004 B.n120 B.n117 10.6151
R1005 B.n121 B.n120 10.6151
R1006 B.n124 B.n121 10.6151
R1007 B.n125 B.n124 10.6151
R1008 B.n128 B.n125 10.6151
R1009 B.n133 B.n130 10.6151
R1010 B.n134 B.n133 10.6151
R1011 B.n137 B.n134 10.6151
R1012 B.n138 B.n137 10.6151
R1013 B.n141 B.n138 10.6151
R1014 B.n142 B.n141 10.6151
R1015 B.n145 B.n142 10.6151
R1016 B.n146 B.n145 10.6151
R1017 B.n149 B.n146 10.6151
R1018 B.n150 B.n149 10.6151
R1019 B.n153 B.n150 10.6151
R1020 B.n154 B.n153 10.6151
R1021 B.n157 B.n154 10.6151
R1022 B.n158 B.n157 10.6151
R1023 B.n161 B.n158 10.6151
R1024 B.n162 B.n161 10.6151
R1025 B.n165 B.n162 10.6151
R1026 B.n166 B.n165 10.6151
R1027 B.n169 B.n166 10.6151
R1028 B.n171 B.n169 10.6151
R1029 B.n172 B.n171 10.6151
R1030 B.n412 B.n172 10.6151
R1031 B.n302 B.n232 8.74196
R1032 B.n279 B.n235 8.74196
R1033 B.n108 B.n107 8.74196
R1034 B.n130 B.n129 8.74196
R1035 B.n452 B.n0 8.11757
R1036 B.n452 B.n1 8.11757
R1037 B.n380 B.t1 4.96664
R1038 B.n12 B.t0 4.96664
R1039 B.n299 B.n232 1.87367
R1040 B.n282 B.n235 1.87367
R1041 B.n109 B.n108 1.87367
R1042 B.n129 B.n128 1.87367
R1043 VP.n0 VP.t0 393.021
R1044 VP.n0 VP.t1 357.543
R1045 VP VP.n0 0.0516364
R1046 VDD1.n28 VDD1.n27 289.615
R1047 VDD1.n57 VDD1.n56 289.615
R1048 VDD1.n27 VDD1.n26 185
R1049 VDD1.n2 VDD1.n1 185
R1050 VDD1.n21 VDD1.n20 185
R1051 VDD1.n19 VDD1.n18 185
R1052 VDD1.n6 VDD1.n5 185
R1053 VDD1.n13 VDD1.n12 185
R1054 VDD1.n11 VDD1.n10 185
R1055 VDD1.n40 VDD1.n39 185
R1056 VDD1.n42 VDD1.n41 185
R1057 VDD1.n35 VDD1.n34 185
R1058 VDD1.n48 VDD1.n47 185
R1059 VDD1.n50 VDD1.n49 185
R1060 VDD1.n31 VDD1.n30 185
R1061 VDD1.n56 VDD1.n55 185
R1062 VDD1.n9 VDD1.t1 149.528
R1063 VDD1.n38 VDD1.t0 149.528
R1064 VDD1.n27 VDD1.n1 104.615
R1065 VDD1.n20 VDD1.n1 104.615
R1066 VDD1.n20 VDD1.n19 104.615
R1067 VDD1.n19 VDD1.n5 104.615
R1068 VDD1.n12 VDD1.n5 104.615
R1069 VDD1.n12 VDD1.n11 104.615
R1070 VDD1.n41 VDD1.n40 104.615
R1071 VDD1.n41 VDD1.n34 104.615
R1072 VDD1.n48 VDD1.n34 104.615
R1073 VDD1.n49 VDD1.n48 104.615
R1074 VDD1.n49 VDD1.n30 104.615
R1075 VDD1.n56 VDD1.n30 104.615
R1076 VDD1 VDD1.n57 82.0051
R1077 VDD1.n11 VDD1.t1 52.3082
R1078 VDD1.n40 VDD1.t0 52.3082
R1079 VDD1 VDD1.n28 50.7411
R1080 VDD1.n26 VDD1.n0 12.0247
R1081 VDD1.n55 VDD1.n29 12.0247
R1082 VDD1.n25 VDD1.n2 11.249
R1083 VDD1.n54 VDD1.n31 11.249
R1084 VDD1.n22 VDD1.n21 10.4732
R1085 VDD1.n51 VDD1.n50 10.4732
R1086 VDD1.n10 VDD1.n9 10.2745
R1087 VDD1.n39 VDD1.n38 10.2745
R1088 VDD1.n18 VDD1.n4 9.69747
R1089 VDD1.n47 VDD1.n33 9.69747
R1090 VDD1.n24 VDD1.n0 9.45567
R1091 VDD1.n53 VDD1.n29 9.45567
R1092 VDD1.n25 VDD1.n24 9.3005
R1093 VDD1.n23 VDD1.n22 9.3005
R1094 VDD1.n4 VDD1.n3 9.3005
R1095 VDD1.n17 VDD1.n16 9.3005
R1096 VDD1.n15 VDD1.n14 9.3005
R1097 VDD1.n8 VDD1.n7 9.3005
R1098 VDD1.n37 VDD1.n36 9.3005
R1099 VDD1.n44 VDD1.n43 9.3005
R1100 VDD1.n46 VDD1.n45 9.3005
R1101 VDD1.n33 VDD1.n32 9.3005
R1102 VDD1.n52 VDD1.n51 9.3005
R1103 VDD1.n54 VDD1.n53 9.3005
R1104 VDD1.n17 VDD1.n6 8.92171
R1105 VDD1.n46 VDD1.n35 8.92171
R1106 VDD1.n14 VDD1.n13 8.14595
R1107 VDD1.n43 VDD1.n42 8.14595
R1108 VDD1.n10 VDD1.n8 7.3702
R1109 VDD1.n39 VDD1.n37 7.3702
R1110 VDD1.n13 VDD1.n8 5.81868
R1111 VDD1.n42 VDD1.n37 5.81868
R1112 VDD1.n14 VDD1.n6 5.04292
R1113 VDD1.n43 VDD1.n35 5.04292
R1114 VDD1.n18 VDD1.n17 4.26717
R1115 VDD1.n47 VDD1.n46 4.26717
R1116 VDD1.n21 VDD1.n4 3.49141
R1117 VDD1.n50 VDD1.n33 3.49141
R1118 VDD1.n9 VDD1.n7 2.84323
R1119 VDD1.n38 VDD1.n36 2.84323
R1120 VDD1.n22 VDD1.n2 2.71565
R1121 VDD1.n51 VDD1.n31 2.71565
R1122 VDD1.n26 VDD1.n25 1.93989
R1123 VDD1.n55 VDD1.n54 1.93989
R1124 VDD1.n28 VDD1.n0 1.16414
R1125 VDD1.n57 VDD1.n29 1.16414
R1126 VDD1.n24 VDD1.n23 0.155672
R1127 VDD1.n23 VDD1.n3 0.155672
R1128 VDD1.n16 VDD1.n3 0.155672
R1129 VDD1.n16 VDD1.n15 0.155672
R1130 VDD1.n15 VDD1.n7 0.155672
R1131 VDD1.n44 VDD1.n36 0.155672
R1132 VDD1.n45 VDD1.n44 0.155672
R1133 VDD1.n45 VDD1.n32 0.155672
R1134 VDD1.n52 VDD1.n32 0.155672
R1135 VDD1.n53 VDD1.n52 0.155672
C0 VP VN 3.50258f
C1 VP VDD2 0.263188f
C2 VDD2 VN 1.17078f
C3 VP VDD1 1.2829f
C4 VN VDD1 0.149018f
C5 VDD2 VDD1 0.481334f
C6 VTAIL VP 1.02963f
C7 VTAIL VN 1.01531f
C8 VTAIL VDD2 3.30642f
C9 VTAIL VDD1 3.26732f
C10 VDD2 B 2.692673f
C11 VDD1 B 4.11863f
C12 VTAIL B 3.979858f
C13 VN B 6.08963f
C14 VP B 3.79643f
C15 VDD1.n0 B 0.008529f
C16 VDD1.n1 B 0.019261f
C17 VDD1.n2 B 0.008628f
C18 VDD1.n3 B 0.015165f
C19 VDD1.n4 B 0.008149f
C20 VDD1.n5 B 0.019261f
C21 VDD1.n6 B 0.008628f
C22 VDD1.n7 B 0.345298f
C23 VDD1.n8 B 0.008149f
C24 VDD1.t1 B 0.032094f
C25 VDD1.n9 B 0.07325f
C26 VDD1.n10 B 0.013615f
C27 VDD1.n11 B 0.014446f
C28 VDD1.n12 B 0.019261f
C29 VDD1.n13 B 0.008628f
C30 VDD1.n14 B 0.008149f
C31 VDD1.n15 B 0.015165f
C32 VDD1.n16 B 0.015165f
C33 VDD1.n17 B 0.008149f
C34 VDD1.n18 B 0.008628f
C35 VDD1.n19 B 0.019261f
C36 VDD1.n20 B 0.019261f
C37 VDD1.n21 B 0.008628f
C38 VDD1.n22 B 0.008149f
C39 VDD1.n23 B 0.015165f
C40 VDD1.n24 B 0.037953f
C41 VDD1.n25 B 0.008149f
C42 VDD1.n26 B 0.008628f
C43 VDD1.n27 B 0.037716f
C44 VDD1.n28 B 0.042294f
C45 VDD1.n29 B 0.008529f
C46 VDD1.n30 B 0.019261f
C47 VDD1.n31 B 0.008628f
C48 VDD1.n32 B 0.015165f
C49 VDD1.n33 B 0.008149f
C50 VDD1.n34 B 0.019261f
C51 VDD1.n35 B 0.008628f
C52 VDD1.n36 B 0.345298f
C53 VDD1.n37 B 0.008149f
C54 VDD1.t0 B 0.032094f
C55 VDD1.n38 B 0.07325f
C56 VDD1.n39 B 0.013615f
C57 VDD1.n40 B 0.014446f
C58 VDD1.n41 B 0.019261f
C59 VDD1.n42 B 0.008628f
C60 VDD1.n43 B 0.008149f
C61 VDD1.n44 B 0.015165f
C62 VDD1.n45 B 0.015165f
C63 VDD1.n46 B 0.008149f
C64 VDD1.n47 B 0.008628f
C65 VDD1.n48 B 0.019261f
C66 VDD1.n49 B 0.019261f
C67 VDD1.n50 B 0.008628f
C68 VDD1.n51 B 0.008149f
C69 VDD1.n52 B 0.015165f
C70 VDD1.n53 B 0.037953f
C71 VDD1.n54 B 0.008149f
C72 VDD1.n55 B 0.008628f
C73 VDD1.n56 B 0.037716f
C74 VDD1.n57 B 0.285429f
C75 VP.t0 B 0.703427f
C76 VP.t1 B 0.601248f
C77 VP.n0 B 2.1797f
C78 VDD2.n0 B 0.008676f
C79 VDD2.n1 B 0.019594f
C80 VDD2.n2 B 0.008777f
C81 VDD2.n3 B 0.015427f
C82 VDD2.n4 B 0.00829f
C83 VDD2.n5 B 0.019594f
C84 VDD2.n6 B 0.008777f
C85 VDD2.n7 B 0.351259f
C86 VDD2.n8 B 0.00829f
C87 VDD2.t0 B 0.032648f
C88 VDD2.n9 B 0.074515f
C89 VDD2.n10 B 0.01385f
C90 VDD2.n11 B 0.014695f
C91 VDD2.n12 B 0.019594f
C92 VDD2.n13 B 0.008777f
C93 VDD2.n14 B 0.00829f
C94 VDD2.n15 B 0.015427f
C95 VDD2.n16 B 0.015427f
C96 VDD2.n17 B 0.00829f
C97 VDD2.n18 B 0.008777f
C98 VDD2.n19 B 0.019594f
C99 VDD2.n20 B 0.019594f
C100 VDD2.n21 B 0.008777f
C101 VDD2.n22 B 0.00829f
C102 VDD2.n23 B 0.015427f
C103 VDD2.n24 B 0.038609f
C104 VDD2.n25 B 0.00829f
C105 VDD2.n26 B 0.008777f
C106 VDD2.n27 B 0.038368f
C107 VDD2.n28 B 0.271649f
C108 VDD2.n29 B 0.008676f
C109 VDD2.n30 B 0.019594f
C110 VDD2.n31 B 0.008777f
C111 VDD2.n32 B 0.015427f
C112 VDD2.n33 B 0.00829f
C113 VDD2.n34 B 0.019594f
C114 VDD2.n35 B 0.008777f
C115 VDD2.n36 B 0.351259f
C116 VDD2.n37 B 0.00829f
C117 VDD2.t1 B 0.032648f
C118 VDD2.n38 B 0.074515f
C119 VDD2.n39 B 0.01385f
C120 VDD2.n40 B 0.014695f
C121 VDD2.n41 B 0.019594f
C122 VDD2.n42 B 0.008777f
C123 VDD2.n43 B 0.00829f
C124 VDD2.n44 B 0.015427f
C125 VDD2.n45 B 0.015427f
C126 VDD2.n46 B 0.00829f
C127 VDD2.n47 B 0.008777f
C128 VDD2.n48 B 0.019594f
C129 VDD2.n49 B 0.019594f
C130 VDD2.n50 B 0.008777f
C131 VDD2.n51 B 0.00829f
C132 VDD2.n52 B 0.015427f
C133 VDD2.n53 B 0.038609f
C134 VDD2.n54 B 0.00829f
C135 VDD2.n55 B 0.008777f
C136 VDD2.n56 B 0.038368f
C137 VDD2.n57 B 0.042724f
C138 VDD2.n58 B 1.27306f
C139 VTAIL.n0 B 0.009748f
C140 VTAIL.n1 B 0.022013f
C141 VTAIL.n2 B 0.009861f
C142 VTAIL.n3 B 0.017332f
C143 VTAIL.n4 B 0.009313f
C144 VTAIL.n5 B 0.022013f
C145 VTAIL.n6 B 0.009861f
C146 VTAIL.n7 B 0.394638f
C147 VTAIL.n8 B 0.009313f
C148 VTAIL.t1 B 0.03668f
C149 VTAIL.n9 B 0.083717f
C150 VTAIL.n10 B 0.015561f
C151 VTAIL.n11 B 0.01651f
C152 VTAIL.n12 B 0.022013f
C153 VTAIL.n13 B 0.009861f
C154 VTAIL.n14 B 0.009313f
C155 VTAIL.n15 B 0.017332f
C156 VTAIL.n16 B 0.017332f
C157 VTAIL.n17 B 0.009313f
C158 VTAIL.n18 B 0.009861f
C159 VTAIL.n19 B 0.022013f
C160 VTAIL.n20 B 0.022013f
C161 VTAIL.n21 B 0.009861f
C162 VTAIL.n22 B 0.009313f
C163 VTAIL.n23 B 0.017332f
C164 VTAIL.n24 B 0.043376f
C165 VTAIL.n25 B 0.009313f
C166 VTAIL.n26 B 0.009861f
C167 VTAIL.n27 B 0.043106f
C168 VTAIL.n28 B 0.036047f
C169 VTAIL.n29 B 0.694349f
C170 VTAIL.n30 B 0.009748f
C171 VTAIL.n31 B 0.022013f
C172 VTAIL.n32 B 0.009861f
C173 VTAIL.n33 B 0.017332f
C174 VTAIL.n34 B 0.009313f
C175 VTAIL.n35 B 0.022013f
C176 VTAIL.n36 B 0.009861f
C177 VTAIL.n37 B 0.394638f
C178 VTAIL.n38 B 0.009313f
C179 VTAIL.t3 B 0.03668f
C180 VTAIL.n39 B 0.083717f
C181 VTAIL.n40 B 0.015561f
C182 VTAIL.n41 B 0.01651f
C183 VTAIL.n42 B 0.022013f
C184 VTAIL.n43 B 0.009861f
C185 VTAIL.n44 B 0.009313f
C186 VTAIL.n45 B 0.017332f
C187 VTAIL.n46 B 0.017332f
C188 VTAIL.n47 B 0.009313f
C189 VTAIL.n48 B 0.009861f
C190 VTAIL.n49 B 0.022013f
C191 VTAIL.n50 B 0.022013f
C192 VTAIL.n51 B 0.009861f
C193 VTAIL.n52 B 0.009313f
C194 VTAIL.n53 B 0.017332f
C195 VTAIL.n54 B 0.043376f
C196 VTAIL.n55 B 0.009313f
C197 VTAIL.n56 B 0.009861f
C198 VTAIL.n57 B 0.043106f
C199 VTAIL.n58 B 0.036047f
C200 VTAIL.n59 B 0.706024f
C201 VTAIL.n60 B 0.009748f
C202 VTAIL.n61 B 0.022013f
C203 VTAIL.n62 B 0.009861f
C204 VTAIL.n63 B 0.017332f
C205 VTAIL.n64 B 0.009313f
C206 VTAIL.n65 B 0.022013f
C207 VTAIL.n66 B 0.009861f
C208 VTAIL.n67 B 0.394638f
C209 VTAIL.n68 B 0.009313f
C210 VTAIL.t0 B 0.03668f
C211 VTAIL.n69 B 0.083717f
C212 VTAIL.n70 B 0.015561f
C213 VTAIL.n71 B 0.01651f
C214 VTAIL.n72 B 0.022013f
C215 VTAIL.n73 B 0.009861f
C216 VTAIL.n74 B 0.009313f
C217 VTAIL.n75 B 0.017332f
C218 VTAIL.n76 B 0.017332f
C219 VTAIL.n77 B 0.009313f
C220 VTAIL.n78 B 0.009861f
C221 VTAIL.n79 B 0.022013f
C222 VTAIL.n80 B 0.022013f
C223 VTAIL.n81 B 0.009861f
C224 VTAIL.n82 B 0.009313f
C225 VTAIL.n83 B 0.017332f
C226 VTAIL.n84 B 0.043376f
C227 VTAIL.n85 B 0.009313f
C228 VTAIL.n86 B 0.009861f
C229 VTAIL.n87 B 0.043106f
C230 VTAIL.n88 B 0.036047f
C231 VTAIL.n89 B 0.646326f
C232 VTAIL.n90 B 0.009748f
C233 VTAIL.n91 B 0.022013f
C234 VTAIL.n92 B 0.009861f
C235 VTAIL.n93 B 0.017332f
C236 VTAIL.n94 B 0.009313f
C237 VTAIL.n95 B 0.022013f
C238 VTAIL.n96 B 0.009861f
C239 VTAIL.n97 B 0.394638f
C240 VTAIL.n98 B 0.009313f
C241 VTAIL.t2 B 0.03668f
C242 VTAIL.n99 B 0.083717f
C243 VTAIL.n100 B 0.015561f
C244 VTAIL.n101 B 0.01651f
C245 VTAIL.n102 B 0.022013f
C246 VTAIL.n103 B 0.009861f
C247 VTAIL.n104 B 0.009313f
C248 VTAIL.n105 B 0.017332f
C249 VTAIL.n106 B 0.017332f
C250 VTAIL.n107 B 0.009313f
C251 VTAIL.n108 B 0.009861f
C252 VTAIL.n109 B 0.022013f
C253 VTAIL.n110 B 0.022013f
C254 VTAIL.n111 B 0.009861f
C255 VTAIL.n112 B 0.009313f
C256 VTAIL.n113 B 0.017332f
C257 VTAIL.n114 B 0.043376f
C258 VTAIL.n115 B 0.009313f
C259 VTAIL.n116 B 0.009861f
C260 VTAIL.n117 B 0.043106f
C261 VTAIL.n118 B 0.036047f
C262 VTAIL.n119 B 0.601913f
C263 VN.t1 B 0.593474f
C264 VN.t0 B 0.697243f
.ends

