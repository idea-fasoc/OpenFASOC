* NGSPICE file created from diff_pair_sample_1206.ext - technology: sky130A

.subckt diff_pair_sample_1206 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=0 ps=0 w=6.58 l=2.05
X1 VDD1.t3 VP.t0 VTAIL.t4 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=1.0857 pd=6.91 as=2.5662 ps=13.94 w=6.58 l=2.05
X2 B.t8 B.t6 B.t7 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=0 ps=0 w=6.58 l=2.05
X3 VTAIL.t7 VP.t1 VDD1.t2 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=1.0857 ps=6.91 w=6.58 l=2.05
X4 VDD2.t3 VN.t0 VTAIL.t2 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=1.0857 pd=6.91 as=2.5662 ps=13.94 w=6.58 l=2.05
X5 VTAIL.t0 VN.t1 VDD2.t2 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=1.0857 ps=6.91 w=6.58 l=2.05
X6 B.t5 B.t3 B.t4 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=0 ps=0 w=6.58 l=2.05
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=1.0857 ps=6.91 w=6.58 l=2.05
X8 VDD1.t1 VP.t2 VTAIL.t5 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=1.0857 pd=6.91 as=2.5662 ps=13.94 w=6.58 l=2.05
X9 VTAIL.t6 VP.t3 VDD1.t0 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=1.0857 ps=6.91 w=6.58 l=2.05
X10 VDD2.t0 VN.t3 VTAIL.t3 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=1.0857 pd=6.91 as=2.5662 ps=13.94 w=6.58 l=2.05
X11 B.t2 B.t0 B.t1 w_n2398_n2284# sky130_fd_pr__pfet_01v8 ad=2.5662 pd=13.94 as=0 ps=0 w=6.58 l=2.05
R0 B.n354 B.n51 585
R1 B.n356 B.n355 585
R2 B.n357 B.n50 585
R3 B.n359 B.n358 585
R4 B.n360 B.n49 585
R5 B.n362 B.n361 585
R6 B.n363 B.n48 585
R7 B.n365 B.n364 585
R8 B.n366 B.n47 585
R9 B.n368 B.n367 585
R10 B.n369 B.n46 585
R11 B.n371 B.n370 585
R12 B.n372 B.n45 585
R13 B.n374 B.n373 585
R14 B.n375 B.n44 585
R15 B.n377 B.n376 585
R16 B.n378 B.n43 585
R17 B.n380 B.n379 585
R18 B.n381 B.n42 585
R19 B.n383 B.n382 585
R20 B.n384 B.n41 585
R21 B.n386 B.n385 585
R22 B.n387 B.n40 585
R23 B.n389 B.n388 585
R24 B.n390 B.n39 585
R25 B.n392 B.n391 585
R26 B.n394 B.n393 585
R27 B.n395 B.n35 585
R28 B.n397 B.n396 585
R29 B.n398 B.n34 585
R30 B.n400 B.n399 585
R31 B.n401 B.n33 585
R32 B.n403 B.n402 585
R33 B.n404 B.n32 585
R34 B.n406 B.n405 585
R35 B.n408 B.n29 585
R36 B.n410 B.n409 585
R37 B.n411 B.n28 585
R38 B.n413 B.n412 585
R39 B.n414 B.n27 585
R40 B.n416 B.n415 585
R41 B.n417 B.n26 585
R42 B.n419 B.n418 585
R43 B.n420 B.n25 585
R44 B.n422 B.n421 585
R45 B.n423 B.n24 585
R46 B.n425 B.n424 585
R47 B.n426 B.n23 585
R48 B.n428 B.n427 585
R49 B.n429 B.n22 585
R50 B.n431 B.n430 585
R51 B.n432 B.n21 585
R52 B.n434 B.n433 585
R53 B.n435 B.n20 585
R54 B.n437 B.n436 585
R55 B.n438 B.n19 585
R56 B.n440 B.n439 585
R57 B.n441 B.n18 585
R58 B.n443 B.n442 585
R59 B.n444 B.n17 585
R60 B.n446 B.n445 585
R61 B.n353 B.n352 585
R62 B.n351 B.n52 585
R63 B.n350 B.n349 585
R64 B.n348 B.n53 585
R65 B.n347 B.n346 585
R66 B.n345 B.n54 585
R67 B.n344 B.n343 585
R68 B.n342 B.n55 585
R69 B.n341 B.n340 585
R70 B.n339 B.n56 585
R71 B.n338 B.n337 585
R72 B.n336 B.n57 585
R73 B.n335 B.n334 585
R74 B.n333 B.n58 585
R75 B.n332 B.n331 585
R76 B.n330 B.n59 585
R77 B.n329 B.n328 585
R78 B.n327 B.n60 585
R79 B.n326 B.n325 585
R80 B.n324 B.n61 585
R81 B.n323 B.n322 585
R82 B.n321 B.n62 585
R83 B.n320 B.n319 585
R84 B.n318 B.n63 585
R85 B.n317 B.n316 585
R86 B.n315 B.n64 585
R87 B.n314 B.n313 585
R88 B.n312 B.n65 585
R89 B.n311 B.n310 585
R90 B.n309 B.n66 585
R91 B.n308 B.n307 585
R92 B.n306 B.n67 585
R93 B.n305 B.n304 585
R94 B.n303 B.n68 585
R95 B.n302 B.n301 585
R96 B.n300 B.n69 585
R97 B.n299 B.n298 585
R98 B.n297 B.n70 585
R99 B.n296 B.n295 585
R100 B.n294 B.n71 585
R101 B.n293 B.n292 585
R102 B.n291 B.n72 585
R103 B.n290 B.n289 585
R104 B.n288 B.n73 585
R105 B.n287 B.n286 585
R106 B.n285 B.n74 585
R107 B.n284 B.n283 585
R108 B.n282 B.n75 585
R109 B.n281 B.n280 585
R110 B.n279 B.n76 585
R111 B.n278 B.n277 585
R112 B.n276 B.n77 585
R113 B.n275 B.n274 585
R114 B.n273 B.n78 585
R115 B.n272 B.n271 585
R116 B.n270 B.n79 585
R117 B.n269 B.n268 585
R118 B.n267 B.n80 585
R119 B.n266 B.n265 585
R120 B.n173 B.n172 585
R121 B.n174 B.n115 585
R122 B.n176 B.n175 585
R123 B.n177 B.n114 585
R124 B.n179 B.n178 585
R125 B.n180 B.n113 585
R126 B.n182 B.n181 585
R127 B.n183 B.n112 585
R128 B.n185 B.n184 585
R129 B.n186 B.n111 585
R130 B.n188 B.n187 585
R131 B.n189 B.n110 585
R132 B.n191 B.n190 585
R133 B.n192 B.n109 585
R134 B.n194 B.n193 585
R135 B.n195 B.n108 585
R136 B.n197 B.n196 585
R137 B.n198 B.n107 585
R138 B.n200 B.n199 585
R139 B.n201 B.n106 585
R140 B.n203 B.n202 585
R141 B.n204 B.n105 585
R142 B.n206 B.n205 585
R143 B.n207 B.n104 585
R144 B.n209 B.n208 585
R145 B.n210 B.n101 585
R146 B.n213 B.n212 585
R147 B.n214 B.n100 585
R148 B.n216 B.n215 585
R149 B.n217 B.n99 585
R150 B.n219 B.n218 585
R151 B.n220 B.n98 585
R152 B.n222 B.n221 585
R153 B.n223 B.n97 585
R154 B.n225 B.n224 585
R155 B.n227 B.n226 585
R156 B.n228 B.n93 585
R157 B.n230 B.n229 585
R158 B.n231 B.n92 585
R159 B.n233 B.n232 585
R160 B.n234 B.n91 585
R161 B.n236 B.n235 585
R162 B.n237 B.n90 585
R163 B.n239 B.n238 585
R164 B.n240 B.n89 585
R165 B.n242 B.n241 585
R166 B.n243 B.n88 585
R167 B.n245 B.n244 585
R168 B.n246 B.n87 585
R169 B.n248 B.n247 585
R170 B.n249 B.n86 585
R171 B.n251 B.n250 585
R172 B.n252 B.n85 585
R173 B.n254 B.n253 585
R174 B.n255 B.n84 585
R175 B.n257 B.n256 585
R176 B.n258 B.n83 585
R177 B.n260 B.n259 585
R178 B.n261 B.n82 585
R179 B.n263 B.n262 585
R180 B.n264 B.n81 585
R181 B.n171 B.n116 585
R182 B.n170 B.n169 585
R183 B.n168 B.n117 585
R184 B.n167 B.n166 585
R185 B.n165 B.n118 585
R186 B.n164 B.n163 585
R187 B.n162 B.n119 585
R188 B.n161 B.n160 585
R189 B.n159 B.n120 585
R190 B.n158 B.n157 585
R191 B.n156 B.n121 585
R192 B.n155 B.n154 585
R193 B.n153 B.n122 585
R194 B.n152 B.n151 585
R195 B.n150 B.n123 585
R196 B.n149 B.n148 585
R197 B.n147 B.n124 585
R198 B.n146 B.n145 585
R199 B.n144 B.n125 585
R200 B.n143 B.n142 585
R201 B.n141 B.n126 585
R202 B.n140 B.n139 585
R203 B.n138 B.n127 585
R204 B.n137 B.n136 585
R205 B.n135 B.n128 585
R206 B.n134 B.n133 585
R207 B.n132 B.n129 585
R208 B.n131 B.n130 585
R209 B.n2 B.n0 585
R210 B.n489 B.n1 585
R211 B.n488 B.n487 585
R212 B.n486 B.n3 585
R213 B.n485 B.n484 585
R214 B.n483 B.n4 585
R215 B.n482 B.n481 585
R216 B.n480 B.n5 585
R217 B.n479 B.n478 585
R218 B.n477 B.n6 585
R219 B.n476 B.n475 585
R220 B.n474 B.n7 585
R221 B.n473 B.n472 585
R222 B.n471 B.n8 585
R223 B.n470 B.n469 585
R224 B.n468 B.n9 585
R225 B.n467 B.n466 585
R226 B.n465 B.n10 585
R227 B.n464 B.n463 585
R228 B.n462 B.n11 585
R229 B.n461 B.n460 585
R230 B.n459 B.n12 585
R231 B.n458 B.n457 585
R232 B.n456 B.n13 585
R233 B.n455 B.n454 585
R234 B.n453 B.n14 585
R235 B.n452 B.n451 585
R236 B.n450 B.n15 585
R237 B.n449 B.n448 585
R238 B.n447 B.n16 585
R239 B.n491 B.n490 585
R240 B.n172 B.n171 511.721
R241 B.n447 B.n446 511.721
R242 B.n266 B.n81 511.721
R243 B.n352 B.n51 511.721
R244 B.n94 B.t8 324.404
R245 B.n36 B.t10 324.404
R246 B.n102 B.t5 324.404
R247 B.n30 B.t1 324.404
R248 B.n94 B.t6 284.389
R249 B.n102 B.t3 284.389
R250 B.n30 B.t0 284.389
R251 B.n36 B.t9 284.389
R252 B.n95 B.t7 278.248
R253 B.n37 B.t11 278.248
R254 B.n103 B.t4 278.248
R255 B.n31 B.t2 278.248
R256 B.n171 B.n170 163.367
R257 B.n170 B.n117 163.367
R258 B.n166 B.n117 163.367
R259 B.n166 B.n165 163.367
R260 B.n165 B.n164 163.367
R261 B.n164 B.n119 163.367
R262 B.n160 B.n119 163.367
R263 B.n160 B.n159 163.367
R264 B.n159 B.n158 163.367
R265 B.n158 B.n121 163.367
R266 B.n154 B.n121 163.367
R267 B.n154 B.n153 163.367
R268 B.n153 B.n152 163.367
R269 B.n152 B.n123 163.367
R270 B.n148 B.n123 163.367
R271 B.n148 B.n147 163.367
R272 B.n147 B.n146 163.367
R273 B.n146 B.n125 163.367
R274 B.n142 B.n125 163.367
R275 B.n142 B.n141 163.367
R276 B.n141 B.n140 163.367
R277 B.n140 B.n127 163.367
R278 B.n136 B.n127 163.367
R279 B.n136 B.n135 163.367
R280 B.n135 B.n134 163.367
R281 B.n134 B.n129 163.367
R282 B.n130 B.n129 163.367
R283 B.n130 B.n2 163.367
R284 B.n490 B.n2 163.367
R285 B.n490 B.n489 163.367
R286 B.n489 B.n488 163.367
R287 B.n488 B.n3 163.367
R288 B.n484 B.n3 163.367
R289 B.n484 B.n483 163.367
R290 B.n483 B.n482 163.367
R291 B.n482 B.n5 163.367
R292 B.n478 B.n5 163.367
R293 B.n478 B.n477 163.367
R294 B.n477 B.n476 163.367
R295 B.n476 B.n7 163.367
R296 B.n472 B.n7 163.367
R297 B.n472 B.n471 163.367
R298 B.n471 B.n470 163.367
R299 B.n470 B.n9 163.367
R300 B.n466 B.n9 163.367
R301 B.n466 B.n465 163.367
R302 B.n465 B.n464 163.367
R303 B.n464 B.n11 163.367
R304 B.n460 B.n11 163.367
R305 B.n460 B.n459 163.367
R306 B.n459 B.n458 163.367
R307 B.n458 B.n13 163.367
R308 B.n454 B.n13 163.367
R309 B.n454 B.n453 163.367
R310 B.n453 B.n452 163.367
R311 B.n452 B.n15 163.367
R312 B.n448 B.n15 163.367
R313 B.n448 B.n447 163.367
R314 B.n172 B.n115 163.367
R315 B.n176 B.n115 163.367
R316 B.n177 B.n176 163.367
R317 B.n178 B.n177 163.367
R318 B.n178 B.n113 163.367
R319 B.n182 B.n113 163.367
R320 B.n183 B.n182 163.367
R321 B.n184 B.n183 163.367
R322 B.n184 B.n111 163.367
R323 B.n188 B.n111 163.367
R324 B.n189 B.n188 163.367
R325 B.n190 B.n189 163.367
R326 B.n190 B.n109 163.367
R327 B.n194 B.n109 163.367
R328 B.n195 B.n194 163.367
R329 B.n196 B.n195 163.367
R330 B.n196 B.n107 163.367
R331 B.n200 B.n107 163.367
R332 B.n201 B.n200 163.367
R333 B.n202 B.n201 163.367
R334 B.n202 B.n105 163.367
R335 B.n206 B.n105 163.367
R336 B.n207 B.n206 163.367
R337 B.n208 B.n207 163.367
R338 B.n208 B.n101 163.367
R339 B.n213 B.n101 163.367
R340 B.n214 B.n213 163.367
R341 B.n215 B.n214 163.367
R342 B.n215 B.n99 163.367
R343 B.n219 B.n99 163.367
R344 B.n220 B.n219 163.367
R345 B.n221 B.n220 163.367
R346 B.n221 B.n97 163.367
R347 B.n225 B.n97 163.367
R348 B.n226 B.n225 163.367
R349 B.n226 B.n93 163.367
R350 B.n230 B.n93 163.367
R351 B.n231 B.n230 163.367
R352 B.n232 B.n231 163.367
R353 B.n232 B.n91 163.367
R354 B.n236 B.n91 163.367
R355 B.n237 B.n236 163.367
R356 B.n238 B.n237 163.367
R357 B.n238 B.n89 163.367
R358 B.n242 B.n89 163.367
R359 B.n243 B.n242 163.367
R360 B.n244 B.n243 163.367
R361 B.n244 B.n87 163.367
R362 B.n248 B.n87 163.367
R363 B.n249 B.n248 163.367
R364 B.n250 B.n249 163.367
R365 B.n250 B.n85 163.367
R366 B.n254 B.n85 163.367
R367 B.n255 B.n254 163.367
R368 B.n256 B.n255 163.367
R369 B.n256 B.n83 163.367
R370 B.n260 B.n83 163.367
R371 B.n261 B.n260 163.367
R372 B.n262 B.n261 163.367
R373 B.n262 B.n81 163.367
R374 B.n267 B.n266 163.367
R375 B.n268 B.n267 163.367
R376 B.n268 B.n79 163.367
R377 B.n272 B.n79 163.367
R378 B.n273 B.n272 163.367
R379 B.n274 B.n273 163.367
R380 B.n274 B.n77 163.367
R381 B.n278 B.n77 163.367
R382 B.n279 B.n278 163.367
R383 B.n280 B.n279 163.367
R384 B.n280 B.n75 163.367
R385 B.n284 B.n75 163.367
R386 B.n285 B.n284 163.367
R387 B.n286 B.n285 163.367
R388 B.n286 B.n73 163.367
R389 B.n290 B.n73 163.367
R390 B.n291 B.n290 163.367
R391 B.n292 B.n291 163.367
R392 B.n292 B.n71 163.367
R393 B.n296 B.n71 163.367
R394 B.n297 B.n296 163.367
R395 B.n298 B.n297 163.367
R396 B.n298 B.n69 163.367
R397 B.n302 B.n69 163.367
R398 B.n303 B.n302 163.367
R399 B.n304 B.n303 163.367
R400 B.n304 B.n67 163.367
R401 B.n308 B.n67 163.367
R402 B.n309 B.n308 163.367
R403 B.n310 B.n309 163.367
R404 B.n310 B.n65 163.367
R405 B.n314 B.n65 163.367
R406 B.n315 B.n314 163.367
R407 B.n316 B.n315 163.367
R408 B.n316 B.n63 163.367
R409 B.n320 B.n63 163.367
R410 B.n321 B.n320 163.367
R411 B.n322 B.n321 163.367
R412 B.n322 B.n61 163.367
R413 B.n326 B.n61 163.367
R414 B.n327 B.n326 163.367
R415 B.n328 B.n327 163.367
R416 B.n328 B.n59 163.367
R417 B.n332 B.n59 163.367
R418 B.n333 B.n332 163.367
R419 B.n334 B.n333 163.367
R420 B.n334 B.n57 163.367
R421 B.n338 B.n57 163.367
R422 B.n339 B.n338 163.367
R423 B.n340 B.n339 163.367
R424 B.n340 B.n55 163.367
R425 B.n344 B.n55 163.367
R426 B.n345 B.n344 163.367
R427 B.n346 B.n345 163.367
R428 B.n346 B.n53 163.367
R429 B.n350 B.n53 163.367
R430 B.n351 B.n350 163.367
R431 B.n352 B.n351 163.367
R432 B.n446 B.n17 163.367
R433 B.n442 B.n17 163.367
R434 B.n442 B.n441 163.367
R435 B.n441 B.n440 163.367
R436 B.n440 B.n19 163.367
R437 B.n436 B.n19 163.367
R438 B.n436 B.n435 163.367
R439 B.n435 B.n434 163.367
R440 B.n434 B.n21 163.367
R441 B.n430 B.n21 163.367
R442 B.n430 B.n429 163.367
R443 B.n429 B.n428 163.367
R444 B.n428 B.n23 163.367
R445 B.n424 B.n23 163.367
R446 B.n424 B.n423 163.367
R447 B.n423 B.n422 163.367
R448 B.n422 B.n25 163.367
R449 B.n418 B.n25 163.367
R450 B.n418 B.n417 163.367
R451 B.n417 B.n416 163.367
R452 B.n416 B.n27 163.367
R453 B.n412 B.n27 163.367
R454 B.n412 B.n411 163.367
R455 B.n411 B.n410 163.367
R456 B.n410 B.n29 163.367
R457 B.n405 B.n29 163.367
R458 B.n405 B.n404 163.367
R459 B.n404 B.n403 163.367
R460 B.n403 B.n33 163.367
R461 B.n399 B.n33 163.367
R462 B.n399 B.n398 163.367
R463 B.n398 B.n397 163.367
R464 B.n397 B.n35 163.367
R465 B.n393 B.n35 163.367
R466 B.n393 B.n392 163.367
R467 B.n392 B.n39 163.367
R468 B.n388 B.n39 163.367
R469 B.n388 B.n387 163.367
R470 B.n387 B.n386 163.367
R471 B.n386 B.n41 163.367
R472 B.n382 B.n41 163.367
R473 B.n382 B.n381 163.367
R474 B.n381 B.n380 163.367
R475 B.n380 B.n43 163.367
R476 B.n376 B.n43 163.367
R477 B.n376 B.n375 163.367
R478 B.n375 B.n374 163.367
R479 B.n374 B.n45 163.367
R480 B.n370 B.n45 163.367
R481 B.n370 B.n369 163.367
R482 B.n369 B.n368 163.367
R483 B.n368 B.n47 163.367
R484 B.n364 B.n47 163.367
R485 B.n364 B.n363 163.367
R486 B.n363 B.n362 163.367
R487 B.n362 B.n49 163.367
R488 B.n358 B.n49 163.367
R489 B.n358 B.n357 163.367
R490 B.n357 B.n356 163.367
R491 B.n356 B.n51 163.367
R492 B.n96 B.n95 59.5399
R493 B.n211 B.n103 59.5399
R494 B.n407 B.n31 59.5399
R495 B.n38 B.n37 59.5399
R496 B.n95 B.n94 46.1581
R497 B.n103 B.n102 46.1581
R498 B.n31 B.n30 46.1581
R499 B.n37 B.n36 46.1581
R500 B.n445 B.n16 33.2493
R501 B.n354 B.n353 33.2493
R502 B.n265 B.n264 33.2493
R503 B.n173 B.n116 33.2493
R504 B B.n491 18.0485
R505 B.n445 B.n444 10.6151
R506 B.n444 B.n443 10.6151
R507 B.n443 B.n18 10.6151
R508 B.n439 B.n18 10.6151
R509 B.n439 B.n438 10.6151
R510 B.n438 B.n437 10.6151
R511 B.n437 B.n20 10.6151
R512 B.n433 B.n20 10.6151
R513 B.n433 B.n432 10.6151
R514 B.n432 B.n431 10.6151
R515 B.n431 B.n22 10.6151
R516 B.n427 B.n22 10.6151
R517 B.n427 B.n426 10.6151
R518 B.n426 B.n425 10.6151
R519 B.n425 B.n24 10.6151
R520 B.n421 B.n24 10.6151
R521 B.n421 B.n420 10.6151
R522 B.n420 B.n419 10.6151
R523 B.n419 B.n26 10.6151
R524 B.n415 B.n26 10.6151
R525 B.n415 B.n414 10.6151
R526 B.n414 B.n413 10.6151
R527 B.n413 B.n28 10.6151
R528 B.n409 B.n28 10.6151
R529 B.n409 B.n408 10.6151
R530 B.n406 B.n32 10.6151
R531 B.n402 B.n32 10.6151
R532 B.n402 B.n401 10.6151
R533 B.n401 B.n400 10.6151
R534 B.n400 B.n34 10.6151
R535 B.n396 B.n34 10.6151
R536 B.n396 B.n395 10.6151
R537 B.n395 B.n394 10.6151
R538 B.n391 B.n390 10.6151
R539 B.n390 B.n389 10.6151
R540 B.n389 B.n40 10.6151
R541 B.n385 B.n40 10.6151
R542 B.n385 B.n384 10.6151
R543 B.n384 B.n383 10.6151
R544 B.n383 B.n42 10.6151
R545 B.n379 B.n42 10.6151
R546 B.n379 B.n378 10.6151
R547 B.n378 B.n377 10.6151
R548 B.n377 B.n44 10.6151
R549 B.n373 B.n44 10.6151
R550 B.n373 B.n372 10.6151
R551 B.n372 B.n371 10.6151
R552 B.n371 B.n46 10.6151
R553 B.n367 B.n46 10.6151
R554 B.n367 B.n366 10.6151
R555 B.n366 B.n365 10.6151
R556 B.n365 B.n48 10.6151
R557 B.n361 B.n48 10.6151
R558 B.n361 B.n360 10.6151
R559 B.n360 B.n359 10.6151
R560 B.n359 B.n50 10.6151
R561 B.n355 B.n50 10.6151
R562 B.n355 B.n354 10.6151
R563 B.n265 B.n80 10.6151
R564 B.n269 B.n80 10.6151
R565 B.n270 B.n269 10.6151
R566 B.n271 B.n270 10.6151
R567 B.n271 B.n78 10.6151
R568 B.n275 B.n78 10.6151
R569 B.n276 B.n275 10.6151
R570 B.n277 B.n276 10.6151
R571 B.n277 B.n76 10.6151
R572 B.n281 B.n76 10.6151
R573 B.n282 B.n281 10.6151
R574 B.n283 B.n282 10.6151
R575 B.n283 B.n74 10.6151
R576 B.n287 B.n74 10.6151
R577 B.n288 B.n287 10.6151
R578 B.n289 B.n288 10.6151
R579 B.n289 B.n72 10.6151
R580 B.n293 B.n72 10.6151
R581 B.n294 B.n293 10.6151
R582 B.n295 B.n294 10.6151
R583 B.n295 B.n70 10.6151
R584 B.n299 B.n70 10.6151
R585 B.n300 B.n299 10.6151
R586 B.n301 B.n300 10.6151
R587 B.n301 B.n68 10.6151
R588 B.n305 B.n68 10.6151
R589 B.n306 B.n305 10.6151
R590 B.n307 B.n306 10.6151
R591 B.n307 B.n66 10.6151
R592 B.n311 B.n66 10.6151
R593 B.n312 B.n311 10.6151
R594 B.n313 B.n312 10.6151
R595 B.n313 B.n64 10.6151
R596 B.n317 B.n64 10.6151
R597 B.n318 B.n317 10.6151
R598 B.n319 B.n318 10.6151
R599 B.n319 B.n62 10.6151
R600 B.n323 B.n62 10.6151
R601 B.n324 B.n323 10.6151
R602 B.n325 B.n324 10.6151
R603 B.n325 B.n60 10.6151
R604 B.n329 B.n60 10.6151
R605 B.n330 B.n329 10.6151
R606 B.n331 B.n330 10.6151
R607 B.n331 B.n58 10.6151
R608 B.n335 B.n58 10.6151
R609 B.n336 B.n335 10.6151
R610 B.n337 B.n336 10.6151
R611 B.n337 B.n56 10.6151
R612 B.n341 B.n56 10.6151
R613 B.n342 B.n341 10.6151
R614 B.n343 B.n342 10.6151
R615 B.n343 B.n54 10.6151
R616 B.n347 B.n54 10.6151
R617 B.n348 B.n347 10.6151
R618 B.n349 B.n348 10.6151
R619 B.n349 B.n52 10.6151
R620 B.n353 B.n52 10.6151
R621 B.n174 B.n173 10.6151
R622 B.n175 B.n174 10.6151
R623 B.n175 B.n114 10.6151
R624 B.n179 B.n114 10.6151
R625 B.n180 B.n179 10.6151
R626 B.n181 B.n180 10.6151
R627 B.n181 B.n112 10.6151
R628 B.n185 B.n112 10.6151
R629 B.n186 B.n185 10.6151
R630 B.n187 B.n186 10.6151
R631 B.n187 B.n110 10.6151
R632 B.n191 B.n110 10.6151
R633 B.n192 B.n191 10.6151
R634 B.n193 B.n192 10.6151
R635 B.n193 B.n108 10.6151
R636 B.n197 B.n108 10.6151
R637 B.n198 B.n197 10.6151
R638 B.n199 B.n198 10.6151
R639 B.n199 B.n106 10.6151
R640 B.n203 B.n106 10.6151
R641 B.n204 B.n203 10.6151
R642 B.n205 B.n204 10.6151
R643 B.n205 B.n104 10.6151
R644 B.n209 B.n104 10.6151
R645 B.n210 B.n209 10.6151
R646 B.n212 B.n100 10.6151
R647 B.n216 B.n100 10.6151
R648 B.n217 B.n216 10.6151
R649 B.n218 B.n217 10.6151
R650 B.n218 B.n98 10.6151
R651 B.n222 B.n98 10.6151
R652 B.n223 B.n222 10.6151
R653 B.n224 B.n223 10.6151
R654 B.n228 B.n227 10.6151
R655 B.n229 B.n228 10.6151
R656 B.n229 B.n92 10.6151
R657 B.n233 B.n92 10.6151
R658 B.n234 B.n233 10.6151
R659 B.n235 B.n234 10.6151
R660 B.n235 B.n90 10.6151
R661 B.n239 B.n90 10.6151
R662 B.n240 B.n239 10.6151
R663 B.n241 B.n240 10.6151
R664 B.n241 B.n88 10.6151
R665 B.n245 B.n88 10.6151
R666 B.n246 B.n245 10.6151
R667 B.n247 B.n246 10.6151
R668 B.n247 B.n86 10.6151
R669 B.n251 B.n86 10.6151
R670 B.n252 B.n251 10.6151
R671 B.n253 B.n252 10.6151
R672 B.n253 B.n84 10.6151
R673 B.n257 B.n84 10.6151
R674 B.n258 B.n257 10.6151
R675 B.n259 B.n258 10.6151
R676 B.n259 B.n82 10.6151
R677 B.n263 B.n82 10.6151
R678 B.n264 B.n263 10.6151
R679 B.n169 B.n116 10.6151
R680 B.n169 B.n168 10.6151
R681 B.n168 B.n167 10.6151
R682 B.n167 B.n118 10.6151
R683 B.n163 B.n118 10.6151
R684 B.n163 B.n162 10.6151
R685 B.n162 B.n161 10.6151
R686 B.n161 B.n120 10.6151
R687 B.n157 B.n120 10.6151
R688 B.n157 B.n156 10.6151
R689 B.n156 B.n155 10.6151
R690 B.n155 B.n122 10.6151
R691 B.n151 B.n122 10.6151
R692 B.n151 B.n150 10.6151
R693 B.n150 B.n149 10.6151
R694 B.n149 B.n124 10.6151
R695 B.n145 B.n124 10.6151
R696 B.n145 B.n144 10.6151
R697 B.n144 B.n143 10.6151
R698 B.n143 B.n126 10.6151
R699 B.n139 B.n126 10.6151
R700 B.n139 B.n138 10.6151
R701 B.n138 B.n137 10.6151
R702 B.n137 B.n128 10.6151
R703 B.n133 B.n128 10.6151
R704 B.n133 B.n132 10.6151
R705 B.n132 B.n131 10.6151
R706 B.n131 B.n0 10.6151
R707 B.n487 B.n1 10.6151
R708 B.n487 B.n486 10.6151
R709 B.n486 B.n485 10.6151
R710 B.n485 B.n4 10.6151
R711 B.n481 B.n4 10.6151
R712 B.n481 B.n480 10.6151
R713 B.n480 B.n479 10.6151
R714 B.n479 B.n6 10.6151
R715 B.n475 B.n6 10.6151
R716 B.n475 B.n474 10.6151
R717 B.n474 B.n473 10.6151
R718 B.n473 B.n8 10.6151
R719 B.n469 B.n8 10.6151
R720 B.n469 B.n468 10.6151
R721 B.n468 B.n467 10.6151
R722 B.n467 B.n10 10.6151
R723 B.n463 B.n10 10.6151
R724 B.n463 B.n462 10.6151
R725 B.n462 B.n461 10.6151
R726 B.n461 B.n12 10.6151
R727 B.n457 B.n12 10.6151
R728 B.n457 B.n456 10.6151
R729 B.n456 B.n455 10.6151
R730 B.n455 B.n14 10.6151
R731 B.n451 B.n14 10.6151
R732 B.n451 B.n450 10.6151
R733 B.n450 B.n449 10.6151
R734 B.n449 B.n16 10.6151
R735 B.n407 B.n406 6.5566
R736 B.n394 B.n38 6.5566
R737 B.n212 B.n211 6.5566
R738 B.n224 B.n96 6.5566
R739 B.n408 B.n407 4.05904
R740 B.n391 B.n38 4.05904
R741 B.n211 B.n210 4.05904
R742 B.n227 B.n96 4.05904
R743 B.n491 B.n0 2.81026
R744 B.n491 B.n1 2.81026
R745 VP.n10 VP.n0 161.3
R746 VP.n9 VP.n8 161.3
R747 VP.n7 VP.n1 161.3
R748 VP.n6 VP.n5 161.3
R749 VP.n2 VP.t3 113.29
R750 VP.n2 VP.t0 112.749
R751 VP.n4 VP.n3 89.2674
R752 VP.n12 VP.n11 89.2674
R753 VP.n4 VP.t1 77.3556
R754 VP.n11 VP.t2 77.3556
R755 VP.n9 VP.n1 56.5617
R756 VP.n3 VP.n2 47.5925
R757 VP.n5 VP.n1 24.5923
R758 VP.n10 VP.n9 24.5923
R759 VP.n5 VP.n4 21.6413
R760 VP.n11 VP.n10 21.6413
R761 VP.n6 VP.n3 0.278335
R762 VP.n12 VP.n0 0.278335
R763 VP.n7 VP.n6 0.189894
R764 VP.n8 VP.n7 0.189894
R765 VP.n8 VP.n0 0.189894
R766 VP VP.n12 0.153485
R767 VTAIL.n270 VTAIL.n269 756.745
R768 VTAIL.n32 VTAIL.n31 756.745
R769 VTAIL.n66 VTAIL.n65 756.745
R770 VTAIL.n100 VTAIL.n99 756.745
R771 VTAIL.n236 VTAIL.n235 756.745
R772 VTAIL.n202 VTAIL.n201 756.745
R773 VTAIL.n168 VTAIL.n167 756.745
R774 VTAIL.n134 VTAIL.n133 756.745
R775 VTAIL.n248 VTAIL.n247 585
R776 VTAIL.n253 VTAIL.n252 585
R777 VTAIL.n255 VTAIL.n254 585
R778 VTAIL.n244 VTAIL.n243 585
R779 VTAIL.n261 VTAIL.n260 585
R780 VTAIL.n263 VTAIL.n262 585
R781 VTAIL.n240 VTAIL.n239 585
R782 VTAIL.n269 VTAIL.n268 585
R783 VTAIL.n10 VTAIL.n9 585
R784 VTAIL.n15 VTAIL.n14 585
R785 VTAIL.n17 VTAIL.n16 585
R786 VTAIL.n6 VTAIL.n5 585
R787 VTAIL.n23 VTAIL.n22 585
R788 VTAIL.n25 VTAIL.n24 585
R789 VTAIL.n2 VTAIL.n1 585
R790 VTAIL.n31 VTAIL.n30 585
R791 VTAIL.n44 VTAIL.n43 585
R792 VTAIL.n49 VTAIL.n48 585
R793 VTAIL.n51 VTAIL.n50 585
R794 VTAIL.n40 VTAIL.n39 585
R795 VTAIL.n57 VTAIL.n56 585
R796 VTAIL.n59 VTAIL.n58 585
R797 VTAIL.n36 VTAIL.n35 585
R798 VTAIL.n65 VTAIL.n64 585
R799 VTAIL.n78 VTAIL.n77 585
R800 VTAIL.n83 VTAIL.n82 585
R801 VTAIL.n85 VTAIL.n84 585
R802 VTAIL.n74 VTAIL.n73 585
R803 VTAIL.n91 VTAIL.n90 585
R804 VTAIL.n93 VTAIL.n92 585
R805 VTAIL.n70 VTAIL.n69 585
R806 VTAIL.n99 VTAIL.n98 585
R807 VTAIL.n235 VTAIL.n234 585
R808 VTAIL.n206 VTAIL.n205 585
R809 VTAIL.n229 VTAIL.n228 585
R810 VTAIL.n227 VTAIL.n226 585
R811 VTAIL.n210 VTAIL.n209 585
R812 VTAIL.n221 VTAIL.n220 585
R813 VTAIL.n219 VTAIL.n218 585
R814 VTAIL.n214 VTAIL.n213 585
R815 VTAIL.n201 VTAIL.n200 585
R816 VTAIL.n172 VTAIL.n171 585
R817 VTAIL.n195 VTAIL.n194 585
R818 VTAIL.n193 VTAIL.n192 585
R819 VTAIL.n176 VTAIL.n175 585
R820 VTAIL.n187 VTAIL.n186 585
R821 VTAIL.n185 VTAIL.n184 585
R822 VTAIL.n180 VTAIL.n179 585
R823 VTAIL.n167 VTAIL.n166 585
R824 VTAIL.n138 VTAIL.n137 585
R825 VTAIL.n161 VTAIL.n160 585
R826 VTAIL.n159 VTAIL.n158 585
R827 VTAIL.n142 VTAIL.n141 585
R828 VTAIL.n153 VTAIL.n152 585
R829 VTAIL.n151 VTAIL.n150 585
R830 VTAIL.n146 VTAIL.n145 585
R831 VTAIL.n133 VTAIL.n132 585
R832 VTAIL.n104 VTAIL.n103 585
R833 VTAIL.n127 VTAIL.n126 585
R834 VTAIL.n125 VTAIL.n124 585
R835 VTAIL.n108 VTAIL.n107 585
R836 VTAIL.n119 VTAIL.n118 585
R837 VTAIL.n117 VTAIL.n116 585
R838 VTAIL.n112 VTAIL.n111 585
R839 VTAIL.n249 VTAIL.t3 329.084
R840 VTAIL.n11 VTAIL.t0 329.084
R841 VTAIL.n45 VTAIL.t5 329.084
R842 VTAIL.n79 VTAIL.t7 329.084
R843 VTAIL.n215 VTAIL.t4 329.084
R844 VTAIL.n181 VTAIL.t6 329.084
R845 VTAIL.n147 VTAIL.t2 329.084
R846 VTAIL.n113 VTAIL.t1 329.084
R847 VTAIL.n253 VTAIL.n247 171.744
R848 VTAIL.n254 VTAIL.n253 171.744
R849 VTAIL.n254 VTAIL.n243 171.744
R850 VTAIL.n261 VTAIL.n243 171.744
R851 VTAIL.n262 VTAIL.n261 171.744
R852 VTAIL.n262 VTAIL.n239 171.744
R853 VTAIL.n269 VTAIL.n239 171.744
R854 VTAIL.n15 VTAIL.n9 171.744
R855 VTAIL.n16 VTAIL.n15 171.744
R856 VTAIL.n16 VTAIL.n5 171.744
R857 VTAIL.n23 VTAIL.n5 171.744
R858 VTAIL.n24 VTAIL.n23 171.744
R859 VTAIL.n24 VTAIL.n1 171.744
R860 VTAIL.n31 VTAIL.n1 171.744
R861 VTAIL.n49 VTAIL.n43 171.744
R862 VTAIL.n50 VTAIL.n49 171.744
R863 VTAIL.n50 VTAIL.n39 171.744
R864 VTAIL.n57 VTAIL.n39 171.744
R865 VTAIL.n58 VTAIL.n57 171.744
R866 VTAIL.n58 VTAIL.n35 171.744
R867 VTAIL.n65 VTAIL.n35 171.744
R868 VTAIL.n83 VTAIL.n77 171.744
R869 VTAIL.n84 VTAIL.n83 171.744
R870 VTAIL.n84 VTAIL.n73 171.744
R871 VTAIL.n91 VTAIL.n73 171.744
R872 VTAIL.n92 VTAIL.n91 171.744
R873 VTAIL.n92 VTAIL.n69 171.744
R874 VTAIL.n99 VTAIL.n69 171.744
R875 VTAIL.n235 VTAIL.n205 171.744
R876 VTAIL.n228 VTAIL.n205 171.744
R877 VTAIL.n228 VTAIL.n227 171.744
R878 VTAIL.n227 VTAIL.n209 171.744
R879 VTAIL.n220 VTAIL.n209 171.744
R880 VTAIL.n220 VTAIL.n219 171.744
R881 VTAIL.n219 VTAIL.n213 171.744
R882 VTAIL.n201 VTAIL.n171 171.744
R883 VTAIL.n194 VTAIL.n171 171.744
R884 VTAIL.n194 VTAIL.n193 171.744
R885 VTAIL.n193 VTAIL.n175 171.744
R886 VTAIL.n186 VTAIL.n175 171.744
R887 VTAIL.n186 VTAIL.n185 171.744
R888 VTAIL.n185 VTAIL.n179 171.744
R889 VTAIL.n167 VTAIL.n137 171.744
R890 VTAIL.n160 VTAIL.n137 171.744
R891 VTAIL.n160 VTAIL.n159 171.744
R892 VTAIL.n159 VTAIL.n141 171.744
R893 VTAIL.n152 VTAIL.n141 171.744
R894 VTAIL.n152 VTAIL.n151 171.744
R895 VTAIL.n151 VTAIL.n145 171.744
R896 VTAIL.n133 VTAIL.n103 171.744
R897 VTAIL.n126 VTAIL.n103 171.744
R898 VTAIL.n126 VTAIL.n125 171.744
R899 VTAIL.n125 VTAIL.n107 171.744
R900 VTAIL.n118 VTAIL.n107 171.744
R901 VTAIL.n118 VTAIL.n117 171.744
R902 VTAIL.n117 VTAIL.n111 171.744
R903 VTAIL.t3 VTAIL.n247 85.8723
R904 VTAIL.t0 VTAIL.n9 85.8723
R905 VTAIL.t5 VTAIL.n43 85.8723
R906 VTAIL.t7 VTAIL.n77 85.8723
R907 VTAIL.t4 VTAIL.n213 85.8723
R908 VTAIL.t6 VTAIL.n179 85.8723
R909 VTAIL.t2 VTAIL.n145 85.8723
R910 VTAIL.t1 VTAIL.n111 85.8723
R911 VTAIL.n271 VTAIL.n270 36.0641
R912 VTAIL.n33 VTAIL.n32 36.0641
R913 VTAIL.n67 VTAIL.n66 36.0641
R914 VTAIL.n101 VTAIL.n100 36.0641
R915 VTAIL.n237 VTAIL.n236 36.0641
R916 VTAIL.n203 VTAIL.n202 36.0641
R917 VTAIL.n169 VTAIL.n168 36.0641
R918 VTAIL.n135 VTAIL.n134 36.0641
R919 VTAIL.n271 VTAIL.n237 20.091
R920 VTAIL.n135 VTAIL.n101 20.091
R921 VTAIL.n268 VTAIL.n238 12.8005
R922 VTAIL.n30 VTAIL.n0 12.8005
R923 VTAIL.n64 VTAIL.n34 12.8005
R924 VTAIL.n98 VTAIL.n68 12.8005
R925 VTAIL.n234 VTAIL.n204 12.8005
R926 VTAIL.n200 VTAIL.n170 12.8005
R927 VTAIL.n166 VTAIL.n136 12.8005
R928 VTAIL.n132 VTAIL.n102 12.8005
R929 VTAIL.n267 VTAIL.n240 12.0247
R930 VTAIL.n29 VTAIL.n2 12.0247
R931 VTAIL.n63 VTAIL.n36 12.0247
R932 VTAIL.n97 VTAIL.n70 12.0247
R933 VTAIL.n233 VTAIL.n206 12.0247
R934 VTAIL.n199 VTAIL.n172 12.0247
R935 VTAIL.n165 VTAIL.n138 12.0247
R936 VTAIL.n131 VTAIL.n104 12.0247
R937 VTAIL.n264 VTAIL.n263 11.249
R938 VTAIL.n26 VTAIL.n25 11.249
R939 VTAIL.n60 VTAIL.n59 11.249
R940 VTAIL.n94 VTAIL.n93 11.249
R941 VTAIL.n230 VTAIL.n229 11.249
R942 VTAIL.n196 VTAIL.n195 11.249
R943 VTAIL.n162 VTAIL.n161 11.249
R944 VTAIL.n128 VTAIL.n127 11.249
R945 VTAIL.n249 VTAIL.n248 10.7233
R946 VTAIL.n11 VTAIL.n10 10.7233
R947 VTAIL.n45 VTAIL.n44 10.7233
R948 VTAIL.n79 VTAIL.n78 10.7233
R949 VTAIL.n215 VTAIL.n214 10.7233
R950 VTAIL.n181 VTAIL.n180 10.7233
R951 VTAIL.n147 VTAIL.n146 10.7233
R952 VTAIL.n113 VTAIL.n112 10.7233
R953 VTAIL.n260 VTAIL.n242 10.4732
R954 VTAIL.n22 VTAIL.n4 10.4732
R955 VTAIL.n56 VTAIL.n38 10.4732
R956 VTAIL.n90 VTAIL.n72 10.4732
R957 VTAIL.n226 VTAIL.n208 10.4732
R958 VTAIL.n192 VTAIL.n174 10.4732
R959 VTAIL.n158 VTAIL.n140 10.4732
R960 VTAIL.n124 VTAIL.n106 10.4732
R961 VTAIL.n259 VTAIL.n244 9.69747
R962 VTAIL.n21 VTAIL.n6 9.69747
R963 VTAIL.n55 VTAIL.n40 9.69747
R964 VTAIL.n89 VTAIL.n74 9.69747
R965 VTAIL.n225 VTAIL.n210 9.69747
R966 VTAIL.n191 VTAIL.n176 9.69747
R967 VTAIL.n157 VTAIL.n142 9.69747
R968 VTAIL.n123 VTAIL.n108 9.69747
R969 VTAIL.n266 VTAIL.n238 9.45567
R970 VTAIL.n28 VTAIL.n0 9.45567
R971 VTAIL.n62 VTAIL.n34 9.45567
R972 VTAIL.n96 VTAIL.n68 9.45567
R973 VTAIL.n232 VTAIL.n204 9.45567
R974 VTAIL.n198 VTAIL.n170 9.45567
R975 VTAIL.n164 VTAIL.n136 9.45567
R976 VTAIL.n130 VTAIL.n102 9.45567
R977 VTAIL.n251 VTAIL.n250 9.3005
R978 VTAIL.n246 VTAIL.n245 9.3005
R979 VTAIL.n257 VTAIL.n256 9.3005
R980 VTAIL.n259 VTAIL.n258 9.3005
R981 VTAIL.n242 VTAIL.n241 9.3005
R982 VTAIL.n265 VTAIL.n264 9.3005
R983 VTAIL.n267 VTAIL.n266 9.3005
R984 VTAIL.n13 VTAIL.n12 9.3005
R985 VTAIL.n8 VTAIL.n7 9.3005
R986 VTAIL.n19 VTAIL.n18 9.3005
R987 VTAIL.n21 VTAIL.n20 9.3005
R988 VTAIL.n4 VTAIL.n3 9.3005
R989 VTAIL.n27 VTAIL.n26 9.3005
R990 VTAIL.n29 VTAIL.n28 9.3005
R991 VTAIL.n47 VTAIL.n46 9.3005
R992 VTAIL.n42 VTAIL.n41 9.3005
R993 VTAIL.n53 VTAIL.n52 9.3005
R994 VTAIL.n55 VTAIL.n54 9.3005
R995 VTAIL.n38 VTAIL.n37 9.3005
R996 VTAIL.n61 VTAIL.n60 9.3005
R997 VTAIL.n63 VTAIL.n62 9.3005
R998 VTAIL.n81 VTAIL.n80 9.3005
R999 VTAIL.n76 VTAIL.n75 9.3005
R1000 VTAIL.n87 VTAIL.n86 9.3005
R1001 VTAIL.n89 VTAIL.n88 9.3005
R1002 VTAIL.n72 VTAIL.n71 9.3005
R1003 VTAIL.n95 VTAIL.n94 9.3005
R1004 VTAIL.n97 VTAIL.n96 9.3005
R1005 VTAIL.n233 VTAIL.n232 9.3005
R1006 VTAIL.n231 VTAIL.n230 9.3005
R1007 VTAIL.n208 VTAIL.n207 9.3005
R1008 VTAIL.n225 VTAIL.n224 9.3005
R1009 VTAIL.n223 VTAIL.n222 9.3005
R1010 VTAIL.n212 VTAIL.n211 9.3005
R1011 VTAIL.n217 VTAIL.n216 9.3005
R1012 VTAIL.n178 VTAIL.n177 9.3005
R1013 VTAIL.n189 VTAIL.n188 9.3005
R1014 VTAIL.n191 VTAIL.n190 9.3005
R1015 VTAIL.n174 VTAIL.n173 9.3005
R1016 VTAIL.n197 VTAIL.n196 9.3005
R1017 VTAIL.n199 VTAIL.n198 9.3005
R1018 VTAIL.n183 VTAIL.n182 9.3005
R1019 VTAIL.n144 VTAIL.n143 9.3005
R1020 VTAIL.n155 VTAIL.n154 9.3005
R1021 VTAIL.n157 VTAIL.n156 9.3005
R1022 VTAIL.n140 VTAIL.n139 9.3005
R1023 VTAIL.n163 VTAIL.n162 9.3005
R1024 VTAIL.n165 VTAIL.n164 9.3005
R1025 VTAIL.n149 VTAIL.n148 9.3005
R1026 VTAIL.n110 VTAIL.n109 9.3005
R1027 VTAIL.n121 VTAIL.n120 9.3005
R1028 VTAIL.n123 VTAIL.n122 9.3005
R1029 VTAIL.n106 VTAIL.n105 9.3005
R1030 VTAIL.n129 VTAIL.n128 9.3005
R1031 VTAIL.n131 VTAIL.n130 9.3005
R1032 VTAIL.n115 VTAIL.n114 9.3005
R1033 VTAIL.n256 VTAIL.n255 8.92171
R1034 VTAIL.n18 VTAIL.n17 8.92171
R1035 VTAIL.n52 VTAIL.n51 8.92171
R1036 VTAIL.n86 VTAIL.n85 8.92171
R1037 VTAIL.n222 VTAIL.n221 8.92171
R1038 VTAIL.n188 VTAIL.n187 8.92171
R1039 VTAIL.n154 VTAIL.n153 8.92171
R1040 VTAIL.n120 VTAIL.n119 8.92171
R1041 VTAIL.n252 VTAIL.n246 8.14595
R1042 VTAIL.n14 VTAIL.n8 8.14595
R1043 VTAIL.n48 VTAIL.n42 8.14595
R1044 VTAIL.n82 VTAIL.n76 8.14595
R1045 VTAIL.n218 VTAIL.n212 8.14595
R1046 VTAIL.n184 VTAIL.n178 8.14595
R1047 VTAIL.n150 VTAIL.n144 8.14595
R1048 VTAIL.n116 VTAIL.n110 8.14595
R1049 VTAIL.n251 VTAIL.n248 7.3702
R1050 VTAIL.n13 VTAIL.n10 7.3702
R1051 VTAIL.n47 VTAIL.n44 7.3702
R1052 VTAIL.n81 VTAIL.n78 7.3702
R1053 VTAIL.n217 VTAIL.n214 7.3702
R1054 VTAIL.n183 VTAIL.n180 7.3702
R1055 VTAIL.n149 VTAIL.n146 7.3702
R1056 VTAIL.n115 VTAIL.n112 7.3702
R1057 VTAIL.n252 VTAIL.n251 5.81868
R1058 VTAIL.n14 VTAIL.n13 5.81868
R1059 VTAIL.n48 VTAIL.n47 5.81868
R1060 VTAIL.n82 VTAIL.n81 5.81868
R1061 VTAIL.n218 VTAIL.n217 5.81868
R1062 VTAIL.n184 VTAIL.n183 5.81868
R1063 VTAIL.n150 VTAIL.n149 5.81868
R1064 VTAIL.n116 VTAIL.n115 5.81868
R1065 VTAIL.n255 VTAIL.n246 5.04292
R1066 VTAIL.n17 VTAIL.n8 5.04292
R1067 VTAIL.n51 VTAIL.n42 5.04292
R1068 VTAIL.n85 VTAIL.n76 5.04292
R1069 VTAIL.n221 VTAIL.n212 5.04292
R1070 VTAIL.n187 VTAIL.n178 5.04292
R1071 VTAIL.n153 VTAIL.n144 5.04292
R1072 VTAIL.n119 VTAIL.n110 5.04292
R1073 VTAIL.n256 VTAIL.n244 4.26717
R1074 VTAIL.n18 VTAIL.n6 4.26717
R1075 VTAIL.n52 VTAIL.n40 4.26717
R1076 VTAIL.n86 VTAIL.n74 4.26717
R1077 VTAIL.n222 VTAIL.n210 4.26717
R1078 VTAIL.n188 VTAIL.n176 4.26717
R1079 VTAIL.n154 VTAIL.n142 4.26717
R1080 VTAIL.n120 VTAIL.n108 4.26717
R1081 VTAIL.n260 VTAIL.n259 3.49141
R1082 VTAIL.n22 VTAIL.n21 3.49141
R1083 VTAIL.n56 VTAIL.n55 3.49141
R1084 VTAIL.n90 VTAIL.n89 3.49141
R1085 VTAIL.n226 VTAIL.n225 3.49141
R1086 VTAIL.n192 VTAIL.n191 3.49141
R1087 VTAIL.n158 VTAIL.n157 3.49141
R1088 VTAIL.n124 VTAIL.n123 3.49141
R1089 VTAIL.n263 VTAIL.n242 2.71565
R1090 VTAIL.n25 VTAIL.n4 2.71565
R1091 VTAIL.n59 VTAIL.n38 2.71565
R1092 VTAIL.n93 VTAIL.n72 2.71565
R1093 VTAIL.n229 VTAIL.n208 2.71565
R1094 VTAIL.n195 VTAIL.n174 2.71565
R1095 VTAIL.n161 VTAIL.n140 2.71565
R1096 VTAIL.n127 VTAIL.n106 2.71565
R1097 VTAIL.n182 VTAIL.n181 2.41347
R1098 VTAIL.n148 VTAIL.n147 2.41347
R1099 VTAIL.n114 VTAIL.n113 2.41347
R1100 VTAIL.n250 VTAIL.n249 2.41347
R1101 VTAIL.n12 VTAIL.n11 2.41347
R1102 VTAIL.n46 VTAIL.n45 2.41347
R1103 VTAIL.n80 VTAIL.n79 2.41347
R1104 VTAIL.n216 VTAIL.n215 2.41347
R1105 VTAIL.n169 VTAIL.n135 2.05222
R1106 VTAIL.n237 VTAIL.n203 2.05222
R1107 VTAIL.n101 VTAIL.n67 2.05222
R1108 VTAIL.n264 VTAIL.n240 1.93989
R1109 VTAIL.n26 VTAIL.n2 1.93989
R1110 VTAIL.n60 VTAIL.n36 1.93989
R1111 VTAIL.n94 VTAIL.n70 1.93989
R1112 VTAIL.n230 VTAIL.n206 1.93989
R1113 VTAIL.n196 VTAIL.n172 1.93989
R1114 VTAIL.n162 VTAIL.n138 1.93989
R1115 VTAIL.n128 VTAIL.n104 1.93989
R1116 VTAIL.n268 VTAIL.n267 1.16414
R1117 VTAIL.n30 VTAIL.n29 1.16414
R1118 VTAIL.n64 VTAIL.n63 1.16414
R1119 VTAIL.n98 VTAIL.n97 1.16414
R1120 VTAIL.n234 VTAIL.n233 1.16414
R1121 VTAIL.n200 VTAIL.n199 1.16414
R1122 VTAIL.n166 VTAIL.n165 1.16414
R1123 VTAIL.n132 VTAIL.n131 1.16414
R1124 VTAIL VTAIL.n33 1.08455
R1125 VTAIL VTAIL.n271 0.968172
R1126 VTAIL.n203 VTAIL.n169 0.470328
R1127 VTAIL.n67 VTAIL.n33 0.470328
R1128 VTAIL.n270 VTAIL.n238 0.388379
R1129 VTAIL.n32 VTAIL.n0 0.388379
R1130 VTAIL.n66 VTAIL.n34 0.388379
R1131 VTAIL.n100 VTAIL.n68 0.388379
R1132 VTAIL.n236 VTAIL.n204 0.388379
R1133 VTAIL.n202 VTAIL.n170 0.388379
R1134 VTAIL.n168 VTAIL.n136 0.388379
R1135 VTAIL.n134 VTAIL.n102 0.388379
R1136 VTAIL.n250 VTAIL.n245 0.155672
R1137 VTAIL.n257 VTAIL.n245 0.155672
R1138 VTAIL.n258 VTAIL.n257 0.155672
R1139 VTAIL.n258 VTAIL.n241 0.155672
R1140 VTAIL.n265 VTAIL.n241 0.155672
R1141 VTAIL.n266 VTAIL.n265 0.155672
R1142 VTAIL.n12 VTAIL.n7 0.155672
R1143 VTAIL.n19 VTAIL.n7 0.155672
R1144 VTAIL.n20 VTAIL.n19 0.155672
R1145 VTAIL.n20 VTAIL.n3 0.155672
R1146 VTAIL.n27 VTAIL.n3 0.155672
R1147 VTAIL.n28 VTAIL.n27 0.155672
R1148 VTAIL.n46 VTAIL.n41 0.155672
R1149 VTAIL.n53 VTAIL.n41 0.155672
R1150 VTAIL.n54 VTAIL.n53 0.155672
R1151 VTAIL.n54 VTAIL.n37 0.155672
R1152 VTAIL.n61 VTAIL.n37 0.155672
R1153 VTAIL.n62 VTAIL.n61 0.155672
R1154 VTAIL.n80 VTAIL.n75 0.155672
R1155 VTAIL.n87 VTAIL.n75 0.155672
R1156 VTAIL.n88 VTAIL.n87 0.155672
R1157 VTAIL.n88 VTAIL.n71 0.155672
R1158 VTAIL.n95 VTAIL.n71 0.155672
R1159 VTAIL.n96 VTAIL.n95 0.155672
R1160 VTAIL.n232 VTAIL.n231 0.155672
R1161 VTAIL.n231 VTAIL.n207 0.155672
R1162 VTAIL.n224 VTAIL.n207 0.155672
R1163 VTAIL.n224 VTAIL.n223 0.155672
R1164 VTAIL.n223 VTAIL.n211 0.155672
R1165 VTAIL.n216 VTAIL.n211 0.155672
R1166 VTAIL.n198 VTAIL.n197 0.155672
R1167 VTAIL.n197 VTAIL.n173 0.155672
R1168 VTAIL.n190 VTAIL.n173 0.155672
R1169 VTAIL.n190 VTAIL.n189 0.155672
R1170 VTAIL.n189 VTAIL.n177 0.155672
R1171 VTAIL.n182 VTAIL.n177 0.155672
R1172 VTAIL.n164 VTAIL.n163 0.155672
R1173 VTAIL.n163 VTAIL.n139 0.155672
R1174 VTAIL.n156 VTAIL.n139 0.155672
R1175 VTAIL.n156 VTAIL.n155 0.155672
R1176 VTAIL.n155 VTAIL.n143 0.155672
R1177 VTAIL.n148 VTAIL.n143 0.155672
R1178 VTAIL.n130 VTAIL.n129 0.155672
R1179 VTAIL.n129 VTAIL.n105 0.155672
R1180 VTAIL.n122 VTAIL.n105 0.155672
R1181 VTAIL.n122 VTAIL.n121 0.155672
R1182 VTAIL.n121 VTAIL.n109 0.155672
R1183 VTAIL.n114 VTAIL.n109 0.155672
R1184 VDD1 VDD1.n1 128.19
R1185 VDD1 VDD1.n0 92.1799
R1186 VDD1.n0 VDD1.t0 4.94047
R1187 VDD1.n0 VDD1.t3 4.94047
R1188 VDD1.n1 VDD1.t2 4.94047
R1189 VDD1.n1 VDD1.t1 4.94047
R1190 VN.n0 VN.t1 113.29
R1191 VN.n1 VN.t0 113.29
R1192 VN.n0 VN.t3 112.749
R1193 VN.n1 VN.t2 112.749
R1194 VN VN.n1 47.8714
R1195 VN VN.n0 7.07214
R1196 VDD2.n2 VDD2.n0 127.665
R1197 VDD2.n2 VDD2.n1 92.1217
R1198 VDD2.n1 VDD2.t1 4.94047
R1199 VDD2.n1 VDD2.t3 4.94047
R1200 VDD2.n0 VDD2.t2 4.94047
R1201 VDD2.n0 VDD2.t0 4.94047
R1202 VDD2 VDD2.n2 0.0586897
C0 VDD1 VDD2 0.896309f
C1 VN VTAIL 2.78126f
C2 VDD2 VTAIL 4.00831f
C3 w_n2398_n2284# VP 4.1586f
C4 w_n2398_n2284# B 7.05446f
C5 B VP 1.44889f
C6 VN VDD2 2.62289f
C7 VDD1 w_n2398_n2284# 1.20287f
C8 VDD1 VP 2.83309f
C9 VTAIL w_n2398_n2284# 2.72597f
C10 VDD1 B 1.01996f
C11 VTAIL VP 2.79536f
C12 VTAIL B 2.96366f
C13 VDD1 VTAIL 3.95779f
C14 VN w_n2398_n2284# 3.85172f
C15 VDD2 w_n2398_n2284# 1.24668f
C16 VN VP 4.78702f
C17 VN B 0.942198f
C18 VDD2 VP 0.359768f
C19 VDD2 B 1.06309f
C20 VN VDD1 0.148963f
C21 VDD2 VSUBS 0.720743f
C22 VDD1 VSUBS 4.672505f
C23 VTAIL VSUBS 0.684933f
C24 VN VSUBS 5.0221f
C25 VP VSUBS 1.70479f
C26 B VSUBS 3.340391f
C27 w_n2398_n2284# VSUBS 68.2279f
C28 VDD2.t2 VSUBS 0.140586f
C29 VDD2.t0 VSUBS 0.140586f
C30 VDD2.n0 VSUBS 1.39328f
C31 VDD2.t1 VSUBS 0.140586f
C32 VDD2.t3 VSUBS 0.140586f
C33 VDD2.n1 VSUBS 0.976157f
C34 VDD2.n2 VSUBS 3.48366f
C35 VN.t1 VSUBS 1.84864f
C36 VN.t3 VSUBS 1.8447f
C37 VN.n0 VSUBS 1.25254f
C38 VN.t0 VSUBS 1.84864f
C39 VN.t2 VSUBS 1.8447f
C40 VN.n1 VSUBS 3.02922f
C41 VDD1.t0 VSUBS 0.142687f
C42 VDD1.t3 VSUBS 0.142687f
C43 VDD1.n0 VSUBS 0.991147f
C44 VDD1.t2 VSUBS 0.142687f
C45 VDD1.t1 VSUBS 0.142687f
C46 VDD1.n1 VSUBS 1.43421f
C47 VTAIL.n0 VSUBS 0.014886f
C48 VTAIL.n1 VSUBS 0.033507f
C49 VTAIL.n2 VSUBS 0.01501f
C50 VTAIL.n3 VSUBS 0.026381f
C51 VTAIL.n4 VSUBS 0.014176f
C52 VTAIL.n5 VSUBS 0.033507f
C53 VTAIL.n6 VSUBS 0.01501f
C54 VTAIL.n7 VSUBS 0.026381f
C55 VTAIL.n8 VSUBS 0.014176f
C56 VTAIL.n9 VSUBS 0.025131f
C57 VTAIL.n10 VSUBS 0.025202f
C58 VTAIL.t0 VSUBS 0.07209f
C59 VTAIL.n11 VSUBS 0.143418f
C60 VTAIL.n12 VSUBS 0.66902f
C61 VTAIL.n13 VSUBS 0.014176f
C62 VTAIL.n14 VSUBS 0.01501f
C63 VTAIL.n15 VSUBS 0.033507f
C64 VTAIL.n16 VSUBS 0.033507f
C65 VTAIL.n17 VSUBS 0.01501f
C66 VTAIL.n18 VSUBS 0.014176f
C67 VTAIL.n19 VSUBS 0.026381f
C68 VTAIL.n20 VSUBS 0.026381f
C69 VTAIL.n21 VSUBS 0.014176f
C70 VTAIL.n22 VSUBS 0.01501f
C71 VTAIL.n23 VSUBS 0.033507f
C72 VTAIL.n24 VSUBS 0.033507f
C73 VTAIL.n25 VSUBS 0.01501f
C74 VTAIL.n26 VSUBS 0.014176f
C75 VTAIL.n27 VSUBS 0.026381f
C76 VTAIL.n28 VSUBS 0.068908f
C77 VTAIL.n29 VSUBS 0.014176f
C78 VTAIL.n30 VSUBS 0.01501f
C79 VTAIL.n31 VSUBS 0.076933f
C80 VTAIL.n32 VSUBS 0.051182f
C81 VTAIL.n33 VSUBS 0.158701f
C82 VTAIL.n34 VSUBS 0.014886f
C83 VTAIL.n35 VSUBS 0.033507f
C84 VTAIL.n36 VSUBS 0.01501f
C85 VTAIL.n37 VSUBS 0.026381f
C86 VTAIL.n38 VSUBS 0.014176f
C87 VTAIL.n39 VSUBS 0.033507f
C88 VTAIL.n40 VSUBS 0.01501f
C89 VTAIL.n41 VSUBS 0.026381f
C90 VTAIL.n42 VSUBS 0.014176f
C91 VTAIL.n43 VSUBS 0.025131f
C92 VTAIL.n44 VSUBS 0.025202f
C93 VTAIL.t5 VSUBS 0.07209f
C94 VTAIL.n45 VSUBS 0.143418f
C95 VTAIL.n46 VSUBS 0.66902f
C96 VTAIL.n47 VSUBS 0.014176f
C97 VTAIL.n48 VSUBS 0.01501f
C98 VTAIL.n49 VSUBS 0.033507f
C99 VTAIL.n50 VSUBS 0.033507f
C100 VTAIL.n51 VSUBS 0.01501f
C101 VTAIL.n52 VSUBS 0.014176f
C102 VTAIL.n53 VSUBS 0.026381f
C103 VTAIL.n54 VSUBS 0.026381f
C104 VTAIL.n55 VSUBS 0.014176f
C105 VTAIL.n56 VSUBS 0.01501f
C106 VTAIL.n57 VSUBS 0.033507f
C107 VTAIL.n58 VSUBS 0.033507f
C108 VTAIL.n59 VSUBS 0.01501f
C109 VTAIL.n60 VSUBS 0.014176f
C110 VTAIL.n61 VSUBS 0.026381f
C111 VTAIL.n62 VSUBS 0.068908f
C112 VTAIL.n63 VSUBS 0.014176f
C113 VTAIL.n64 VSUBS 0.01501f
C114 VTAIL.n65 VSUBS 0.076933f
C115 VTAIL.n66 VSUBS 0.051182f
C116 VTAIL.n67 VSUBS 0.24096f
C117 VTAIL.n68 VSUBS 0.014886f
C118 VTAIL.n69 VSUBS 0.033507f
C119 VTAIL.n70 VSUBS 0.01501f
C120 VTAIL.n71 VSUBS 0.026381f
C121 VTAIL.n72 VSUBS 0.014176f
C122 VTAIL.n73 VSUBS 0.033507f
C123 VTAIL.n74 VSUBS 0.01501f
C124 VTAIL.n75 VSUBS 0.026381f
C125 VTAIL.n76 VSUBS 0.014176f
C126 VTAIL.n77 VSUBS 0.025131f
C127 VTAIL.n78 VSUBS 0.025202f
C128 VTAIL.t7 VSUBS 0.07209f
C129 VTAIL.n79 VSUBS 0.143418f
C130 VTAIL.n80 VSUBS 0.66902f
C131 VTAIL.n81 VSUBS 0.014176f
C132 VTAIL.n82 VSUBS 0.01501f
C133 VTAIL.n83 VSUBS 0.033507f
C134 VTAIL.n84 VSUBS 0.033507f
C135 VTAIL.n85 VSUBS 0.01501f
C136 VTAIL.n86 VSUBS 0.014176f
C137 VTAIL.n87 VSUBS 0.026381f
C138 VTAIL.n88 VSUBS 0.026381f
C139 VTAIL.n89 VSUBS 0.014176f
C140 VTAIL.n90 VSUBS 0.01501f
C141 VTAIL.n91 VSUBS 0.033507f
C142 VTAIL.n92 VSUBS 0.033507f
C143 VTAIL.n93 VSUBS 0.01501f
C144 VTAIL.n94 VSUBS 0.014176f
C145 VTAIL.n95 VSUBS 0.026381f
C146 VTAIL.n96 VSUBS 0.068908f
C147 VTAIL.n97 VSUBS 0.014176f
C148 VTAIL.n98 VSUBS 0.01501f
C149 VTAIL.n99 VSUBS 0.076933f
C150 VTAIL.n100 VSUBS 0.051182f
C151 VTAIL.n101 VSUBS 1.21599f
C152 VTAIL.n102 VSUBS 0.014886f
C153 VTAIL.n103 VSUBS 0.033507f
C154 VTAIL.n104 VSUBS 0.01501f
C155 VTAIL.n105 VSUBS 0.026381f
C156 VTAIL.n106 VSUBS 0.014176f
C157 VTAIL.n107 VSUBS 0.033507f
C158 VTAIL.n108 VSUBS 0.01501f
C159 VTAIL.n109 VSUBS 0.026381f
C160 VTAIL.n110 VSUBS 0.014176f
C161 VTAIL.n111 VSUBS 0.025131f
C162 VTAIL.n112 VSUBS 0.025202f
C163 VTAIL.t1 VSUBS 0.07209f
C164 VTAIL.n113 VSUBS 0.143418f
C165 VTAIL.n114 VSUBS 0.66902f
C166 VTAIL.n115 VSUBS 0.014176f
C167 VTAIL.n116 VSUBS 0.01501f
C168 VTAIL.n117 VSUBS 0.033507f
C169 VTAIL.n118 VSUBS 0.033507f
C170 VTAIL.n119 VSUBS 0.01501f
C171 VTAIL.n120 VSUBS 0.014176f
C172 VTAIL.n121 VSUBS 0.026381f
C173 VTAIL.n122 VSUBS 0.026381f
C174 VTAIL.n123 VSUBS 0.014176f
C175 VTAIL.n124 VSUBS 0.01501f
C176 VTAIL.n125 VSUBS 0.033507f
C177 VTAIL.n126 VSUBS 0.033507f
C178 VTAIL.n127 VSUBS 0.01501f
C179 VTAIL.n128 VSUBS 0.014176f
C180 VTAIL.n129 VSUBS 0.026381f
C181 VTAIL.n130 VSUBS 0.068908f
C182 VTAIL.n131 VSUBS 0.014176f
C183 VTAIL.n132 VSUBS 0.01501f
C184 VTAIL.n133 VSUBS 0.076933f
C185 VTAIL.n134 VSUBS 0.051182f
C186 VTAIL.n135 VSUBS 1.21599f
C187 VTAIL.n136 VSUBS 0.014886f
C188 VTAIL.n137 VSUBS 0.033507f
C189 VTAIL.n138 VSUBS 0.01501f
C190 VTAIL.n139 VSUBS 0.026381f
C191 VTAIL.n140 VSUBS 0.014176f
C192 VTAIL.n141 VSUBS 0.033507f
C193 VTAIL.n142 VSUBS 0.01501f
C194 VTAIL.n143 VSUBS 0.026381f
C195 VTAIL.n144 VSUBS 0.014176f
C196 VTAIL.n145 VSUBS 0.025131f
C197 VTAIL.n146 VSUBS 0.025202f
C198 VTAIL.t2 VSUBS 0.07209f
C199 VTAIL.n147 VSUBS 0.143418f
C200 VTAIL.n148 VSUBS 0.66902f
C201 VTAIL.n149 VSUBS 0.014176f
C202 VTAIL.n150 VSUBS 0.01501f
C203 VTAIL.n151 VSUBS 0.033507f
C204 VTAIL.n152 VSUBS 0.033507f
C205 VTAIL.n153 VSUBS 0.01501f
C206 VTAIL.n154 VSUBS 0.014176f
C207 VTAIL.n155 VSUBS 0.026381f
C208 VTAIL.n156 VSUBS 0.026381f
C209 VTAIL.n157 VSUBS 0.014176f
C210 VTAIL.n158 VSUBS 0.01501f
C211 VTAIL.n159 VSUBS 0.033507f
C212 VTAIL.n160 VSUBS 0.033507f
C213 VTAIL.n161 VSUBS 0.01501f
C214 VTAIL.n162 VSUBS 0.014176f
C215 VTAIL.n163 VSUBS 0.026381f
C216 VTAIL.n164 VSUBS 0.068908f
C217 VTAIL.n165 VSUBS 0.014176f
C218 VTAIL.n166 VSUBS 0.01501f
C219 VTAIL.n167 VSUBS 0.076933f
C220 VTAIL.n168 VSUBS 0.051182f
C221 VTAIL.n169 VSUBS 0.24096f
C222 VTAIL.n170 VSUBS 0.014886f
C223 VTAIL.n171 VSUBS 0.033507f
C224 VTAIL.n172 VSUBS 0.01501f
C225 VTAIL.n173 VSUBS 0.026381f
C226 VTAIL.n174 VSUBS 0.014176f
C227 VTAIL.n175 VSUBS 0.033507f
C228 VTAIL.n176 VSUBS 0.01501f
C229 VTAIL.n177 VSUBS 0.026381f
C230 VTAIL.n178 VSUBS 0.014176f
C231 VTAIL.n179 VSUBS 0.025131f
C232 VTAIL.n180 VSUBS 0.025202f
C233 VTAIL.t6 VSUBS 0.07209f
C234 VTAIL.n181 VSUBS 0.143418f
C235 VTAIL.n182 VSUBS 0.66902f
C236 VTAIL.n183 VSUBS 0.014176f
C237 VTAIL.n184 VSUBS 0.01501f
C238 VTAIL.n185 VSUBS 0.033507f
C239 VTAIL.n186 VSUBS 0.033507f
C240 VTAIL.n187 VSUBS 0.01501f
C241 VTAIL.n188 VSUBS 0.014176f
C242 VTAIL.n189 VSUBS 0.026381f
C243 VTAIL.n190 VSUBS 0.026381f
C244 VTAIL.n191 VSUBS 0.014176f
C245 VTAIL.n192 VSUBS 0.01501f
C246 VTAIL.n193 VSUBS 0.033507f
C247 VTAIL.n194 VSUBS 0.033507f
C248 VTAIL.n195 VSUBS 0.01501f
C249 VTAIL.n196 VSUBS 0.014176f
C250 VTAIL.n197 VSUBS 0.026381f
C251 VTAIL.n198 VSUBS 0.068908f
C252 VTAIL.n199 VSUBS 0.014176f
C253 VTAIL.n200 VSUBS 0.01501f
C254 VTAIL.n201 VSUBS 0.076933f
C255 VTAIL.n202 VSUBS 0.051182f
C256 VTAIL.n203 VSUBS 0.24096f
C257 VTAIL.n204 VSUBS 0.014886f
C258 VTAIL.n205 VSUBS 0.033507f
C259 VTAIL.n206 VSUBS 0.01501f
C260 VTAIL.n207 VSUBS 0.026381f
C261 VTAIL.n208 VSUBS 0.014176f
C262 VTAIL.n209 VSUBS 0.033507f
C263 VTAIL.n210 VSUBS 0.01501f
C264 VTAIL.n211 VSUBS 0.026381f
C265 VTAIL.n212 VSUBS 0.014176f
C266 VTAIL.n213 VSUBS 0.025131f
C267 VTAIL.n214 VSUBS 0.025202f
C268 VTAIL.t4 VSUBS 0.07209f
C269 VTAIL.n215 VSUBS 0.143418f
C270 VTAIL.n216 VSUBS 0.66902f
C271 VTAIL.n217 VSUBS 0.014176f
C272 VTAIL.n218 VSUBS 0.01501f
C273 VTAIL.n219 VSUBS 0.033507f
C274 VTAIL.n220 VSUBS 0.033507f
C275 VTAIL.n221 VSUBS 0.01501f
C276 VTAIL.n222 VSUBS 0.014176f
C277 VTAIL.n223 VSUBS 0.026381f
C278 VTAIL.n224 VSUBS 0.026381f
C279 VTAIL.n225 VSUBS 0.014176f
C280 VTAIL.n226 VSUBS 0.01501f
C281 VTAIL.n227 VSUBS 0.033507f
C282 VTAIL.n228 VSUBS 0.033507f
C283 VTAIL.n229 VSUBS 0.01501f
C284 VTAIL.n230 VSUBS 0.014176f
C285 VTAIL.n231 VSUBS 0.026381f
C286 VTAIL.n232 VSUBS 0.068908f
C287 VTAIL.n233 VSUBS 0.014176f
C288 VTAIL.n234 VSUBS 0.01501f
C289 VTAIL.n235 VSUBS 0.076933f
C290 VTAIL.n236 VSUBS 0.051182f
C291 VTAIL.n237 VSUBS 1.21599f
C292 VTAIL.n238 VSUBS 0.014886f
C293 VTAIL.n239 VSUBS 0.033507f
C294 VTAIL.n240 VSUBS 0.01501f
C295 VTAIL.n241 VSUBS 0.026381f
C296 VTAIL.n242 VSUBS 0.014176f
C297 VTAIL.n243 VSUBS 0.033507f
C298 VTAIL.n244 VSUBS 0.01501f
C299 VTAIL.n245 VSUBS 0.026381f
C300 VTAIL.n246 VSUBS 0.014176f
C301 VTAIL.n247 VSUBS 0.025131f
C302 VTAIL.n248 VSUBS 0.025202f
C303 VTAIL.t3 VSUBS 0.07209f
C304 VTAIL.n249 VSUBS 0.143418f
C305 VTAIL.n250 VSUBS 0.66902f
C306 VTAIL.n251 VSUBS 0.014176f
C307 VTAIL.n252 VSUBS 0.01501f
C308 VTAIL.n253 VSUBS 0.033507f
C309 VTAIL.n254 VSUBS 0.033507f
C310 VTAIL.n255 VSUBS 0.01501f
C311 VTAIL.n256 VSUBS 0.014176f
C312 VTAIL.n257 VSUBS 0.026381f
C313 VTAIL.n258 VSUBS 0.026381f
C314 VTAIL.n259 VSUBS 0.014176f
C315 VTAIL.n260 VSUBS 0.01501f
C316 VTAIL.n261 VSUBS 0.033507f
C317 VTAIL.n262 VSUBS 0.033507f
C318 VTAIL.n263 VSUBS 0.01501f
C319 VTAIL.n264 VSUBS 0.014176f
C320 VTAIL.n265 VSUBS 0.026381f
C321 VTAIL.n266 VSUBS 0.068908f
C322 VTAIL.n267 VSUBS 0.014176f
C323 VTAIL.n268 VSUBS 0.01501f
C324 VTAIL.n269 VSUBS 0.076933f
C325 VTAIL.n270 VSUBS 0.051182f
C326 VTAIL.n271 VSUBS 1.12383f
C327 VP.n0 VSUBS 0.060502f
C328 VP.t2 VSUBS 1.64699f
C329 VP.n1 VSUBS 0.066713f
C330 VP.t0 VSUBS 1.91855f
C331 VP.t3 VSUBS 1.92266f
C332 VP.n2 VSUBS 3.12682f
C333 VP.n3 VSUBS 2.18406f
C334 VP.t1 VSUBS 1.64699f
C335 VP.n4 VSUBS 0.768568f
C336 VP.n5 VSUBS 0.080063f
C337 VP.n6 VSUBS 0.060502f
C338 VP.n7 VSUBS 0.045893f
C339 VP.n8 VSUBS 0.045893f
C340 VP.n9 VSUBS 0.066713f
C341 VP.n10 VSUBS 0.080063f
C342 VP.n11 VSUBS 0.768568f
C343 VP.n12 VSUBS 0.053602f
C344 B.n0 VSUBS 0.005282f
C345 B.n1 VSUBS 0.005282f
C346 B.n2 VSUBS 0.008353f
C347 B.n3 VSUBS 0.008353f
C348 B.n4 VSUBS 0.008353f
C349 B.n5 VSUBS 0.008353f
C350 B.n6 VSUBS 0.008353f
C351 B.n7 VSUBS 0.008353f
C352 B.n8 VSUBS 0.008353f
C353 B.n9 VSUBS 0.008353f
C354 B.n10 VSUBS 0.008353f
C355 B.n11 VSUBS 0.008353f
C356 B.n12 VSUBS 0.008353f
C357 B.n13 VSUBS 0.008353f
C358 B.n14 VSUBS 0.008353f
C359 B.n15 VSUBS 0.008353f
C360 B.n16 VSUBS 0.019198f
C361 B.n17 VSUBS 0.008353f
C362 B.n18 VSUBS 0.008353f
C363 B.n19 VSUBS 0.008353f
C364 B.n20 VSUBS 0.008353f
C365 B.n21 VSUBS 0.008353f
C366 B.n22 VSUBS 0.008353f
C367 B.n23 VSUBS 0.008353f
C368 B.n24 VSUBS 0.008353f
C369 B.n25 VSUBS 0.008353f
C370 B.n26 VSUBS 0.008353f
C371 B.n27 VSUBS 0.008353f
C372 B.n28 VSUBS 0.008353f
C373 B.n29 VSUBS 0.008353f
C374 B.t2 VSUBS 0.118883f
C375 B.t1 VSUBS 0.145203f
C376 B.t0 VSUBS 0.748073f
C377 B.n30 VSUBS 0.248941f
C378 B.n31 VSUBS 0.196893f
C379 B.n32 VSUBS 0.008353f
C380 B.n33 VSUBS 0.008353f
C381 B.n34 VSUBS 0.008353f
C382 B.n35 VSUBS 0.008353f
C383 B.t11 VSUBS 0.118886f
C384 B.t10 VSUBS 0.145205f
C385 B.t9 VSUBS 0.748073f
C386 B.n36 VSUBS 0.248939f
C387 B.n37 VSUBS 0.196891f
C388 B.n38 VSUBS 0.019353f
C389 B.n39 VSUBS 0.008353f
C390 B.n40 VSUBS 0.008353f
C391 B.n41 VSUBS 0.008353f
C392 B.n42 VSUBS 0.008353f
C393 B.n43 VSUBS 0.008353f
C394 B.n44 VSUBS 0.008353f
C395 B.n45 VSUBS 0.008353f
C396 B.n46 VSUBS 0.008353f
C397 B.n47 VSUBS 0.008353f
C398 B.n48 VSUBS 0.008353f
C399 B.n49 VSUBS 0.008353f
C400 B.n50 VSUBS 0.008353f
C401 B.n51 VSUBS 0.020357f
C402 B.n52 VSUBS 0.008353f
C403 B.n53 VSUBS 0.008353f
C404 B.n54 VSUBS 0.008353f
C405 B.n55 VSUBS 0.008353f
C406 B.n56 VSUBS 0.008353f
C407 B.n57 VSUBS 0.008353f
C408 B.n58 VSUBS 0.008353f
C409 B.n59 VSUBS 0.008353f
C410 B.n60 VSUBS 0.008353f
C411 B.n61 VSUBS 0.008353f
C412 B.n62 VSUBS 0.008353f
C413 B.n63 VSUBS 0.008353f
C414 B.n64 VSUBS 0.008353f
C415 B.n65 VSUBS 0.008353f
C416 B.n66 VSUBS 0.008353f
C417 B.n67 VSUBS 0.008353f
C418 B.n68 VSUBS 0.008353f
C419 B.n69 VSUBS 0.008353f
C420 B.n70 VSUBS 0.008353f
C421 B.n71 VSUBS 0.008353f
C422 B.n72 VSUBS 0.008353f
C423 B.n73 VSUBS 0.008353f
C424 B.n74 VSUBS 0.008353f
C425 B.n75 VSUBS 0.008353f
C426 B.n76 VSUBS 0.008353f
C427 B.n77 VSUBS 0.008353f
C428 B.n78 VSUBS 0.008353f
C429 B.n79 VSUBS 0.008353f
C430 B.n80 VSUBS 0.008353f
C431 B.n81 VSUBS 0.020357f
C432 B.n82 VSUBS 0.008353f
C433 B.n83 VSUBS 0.008353f
C434 B.n84 VSUBS 0.008353f
C435 B.n85 VSUBS 0.008353f
C436 B.n86 VSUBS 0.008353f
C437 B.n87 VSUBS 0.008353f
C438 B.n88 VSUBS 0.008353f
C439 B.n89 VSUBS 0.008353f
C440 B.n90 VSUBS 0.008353f
C441 B.n91 VSUBS 0.008353f
C442 B.n92 VSUBS 0.008353f
C443 B.n93 VSUBS 0.008353f
C444 B.t7 VSUBS 0.118886f
C445 B.t8 VSUBS 0.145205f
C446 B.t6 VSUBS 0.748073f
C447 B.n94 VSUBS 0.248939f
C448 B.n95 VSUBS 0.196891f
C449 B.n96 VSUBS 0.019353f
C450 B.n97 VSUBS 0.008353f
C451 B.n98 VSUBS 0.008353f
C452 B.n99 VSUBS 0.008353f
C453 B.n100 VSUBS 0.008353f
C454 B.n101 VSUBS 0.008353f
C455 B.t4 VSUBS 0.118883f
C456 B.t5 VSUBS 0.145203f
C457 B.t3 VSUBS 0.748073f
C458 B.n102 VSUBS 0.248941f
C459 B.n103 VSUBS 0.196893f
C460 B.n104 VSUBS 0.008353f
C461 B.n105 VSUBS 0.008353f
C462 B.n106 VSUBS 0.008353f
C463 B.n107 VSUBS 0.008353f
C464 B.n108 VSUBS 0.008353f
C465 B.n109 VSUBS 0.008353f
C466 B.n110 VSUBS 0.008353f
C467 B.n111 VSUBS 0.008353f
C468 B.n112 VSUBS 0.008353f
C469 B.n113 VSUBS 0.008353f
C470 B.n114 VSUBS 0.008353f
C471 B.n115 VSUBS 0.008353f
C472 B.n116 VSUBS 0.019198f
C473 B.n117 VSUBS 0.008353f
C474 B.n118 VSUBS 0.008353f
C475 B.n119 VSUBS 0.008353f
C476 B.n120 VSUBS 0.008353f
C477 B.n121 VSUBS 0.008353f
C478 B.n122 VSUBS 0.008353f
C479 B.n123 VSUBS 0.008353f
C480 B.n124 VSUBS 0.008353f
C481 B.n125 VSUBS 0.008353f
C482 B.n126 VSUBS 0.008353f
C483 B.n127 VSUBS 0.008353f
C484 B.n128 VSUBS 0.008353f
C485 B.n129 VSUBS 0.008353f
C486 B.n130 VSUBS 0.008353f
C487 B.n131 VSUBS 0.008353f
C488 B.n132 VSUBS 0.008353f
C489 B.n133 VSUBS 0.008353f
C490 B.n134 VSUBS 0.008353f
C491 B.n135 VSUBS 0.008353f
C492 B.n136 VSUBS 0.008353f
C493 B.n137 VSUBS 0.008353f
C494 B.n138 VSUBS 0.008353f
C495 B.n139 VSUBS 0.008353f
C496 B.n140 VSUBS 0.008353f
C497 B.n141 VSUBS 0.008353f
C498 B.n142 VSUBS 0.008353f
C499 B.n143 VSUBS 0.008353f
C500 B.n144 VSUBS 0.008353f
C501 B.n145 VSUBS 0.008353f
C502 B.n146 VSUBS 0.008353f
C503 B.n147 VSUBS 0.008353f
C504 B.n148 VSUBS 0.008353f
C505 B.n149 VSUBS 0.008353f
C506 B.n150 VSUBS 0.008353f
C507 B.n151 VSUBS 0.008353f
C508 B.n152 VSUBS 0.008353f
C509 B.n153 VSUBS 0.008353f
C510 B.n154 VSUBS 0.008353f
C511 B.n155 VSUBS 0.008353f
C512 B.n156 VSUBS 0.008353f
C513 B.n157 VSUBS 0.008353f
C514 B.n158 VSUBS 0.008353f
C515 B.n159 VSUBS 0.008353f
C516 B.n160 VSUBS 0.008353f
C517 B.n161 VSUBS 0.008353f
C518 B.n162 VSUBS 0.008353f
C519 B.n163 VSUBS 0.008353f
C520 B.n164 VSUBS 0.008353f
C521 B.n165 VSUBS 0.008353f
C522 B.n166 VSUBS 0.008353f
C523 B.n167 VSUBS 0.008353f
C524 B.n168 VSUBS 0.008353f
C525 B.n169 VSUBS 0.008353f
C526 B.n170 VSUBS 0.008353f
C527 B.n171 VSUBS 0.019198f
C528 B.n172 VSUBS 0.020357f
C529 B.n173 VSUBS 0.020357f
C530 B.n174 VSUBS 0.008353f
C531 B.n175 VSUBS 0.008353f
C532 B.n176 VSUBS 0.008353f
C533 B.n177 VSUBS 0.008353f
C534 B.n178 VSUBS 0.008353f
C535 B.n179 VSUBS 0.008353f
C536 B.n180 VSUBS 0.008353f
C537 B.n181 VSUBS 0.008353f
C538 B.n182 VSUBS 0.008353f
C539 B.n183 VSUBS 0.008353f
C540 B.n184 VSUBS 0.008353f
C541 B.n185 VSUBS 0.008353f
C542 B.n186 VSUBS 0.008353f
C543 B.n187 VSUBS 0.008353f
C544 B.n188 VSUBS 0.008353f
C545 B.n189 VSUBS 0.008353f
C546 B.n190 VSUBS 0.008353f
C547 B.n191 VSUBS 0.008353f
C548 B.n192 VSUBS 0.008353f
C549 B.n193 VSUBS 0.008353f
C550 B.n194 VSUBS 0.008353f
C551 B.n195 VSUBS 0.008353f
C552 B.n196 VSUBS 0.008353f
C553 B.n197 VSUBS 0.008353f
C554 B.n198 VSUBS 0.008353f
C555 B.n199 VSUBS 0.008353f
C556 B.n200 VSUBS 0.008353f
C557 B.n201 VSUBS 0.008353f
C558 B.n202 VSUBS 0.008353f
C559 B.n203 VSUBS 0.008353f
C560 B.n204 VSUBS 0.008353f
C561 B.n205 VSUBS 0.008353f
C562 B.n206 VSUBS 0.008353f
C563 B.n207 VSUBS 0.008353f
C564 B.n208 VSUBS 0.008353f
C565 B.n209 VSUBS 0.008353f
C566 B.n210 VSUBS 0.005774f
C567 B.n211 VSUBS 0.019353f
C568 B.n212 VSUBS 0.006756f
C569 B.n213 VSUBS 0.008353f
C570 B.n214 VSUBS 0.008353f
C571 B.n215 VSUBS 0.008353f
C572 B.n216 VSUBS 0.008353f
C573 B.n217 VSUBS 0.008353f
C574 B.n218 VSUBS 0.008353f
C575 B.n219 VSUBS 0.008353f
C576 B.n220 VSUBS 0.008353f
C577 B.n221 VSUBS 0.008353f
C578 B.n222 VSUBS 0.008353f
C579 B.n223 VSUBS 0.008353f
C580 B.n224 VSUBS 0.006756f
C581 B.n225 VSUBS 0.008353f
C582 B.n226 VSUBS 0.008353f
C583 B.n227 VSUBS 0.005774f
C584 B.n228 VSUBS 0.008353f
C585 B.n229 VSUBS 0.008353f
C586 B.n230 VSUBS 0.008353f
C587 B.n231 VSUBS 0.008353f
C588 B.n232 VSUBS 0.008353f
C589 B.n233 VSUBS 0.008353f
C590 B.n234 VSUBS 0.008353f
C591 B.n235 VSUBS 0.008353f
C592 B.n236 VSUBS 0.008353f
C593 B.n237 VSUBS 0.008353f
C594 B.n238 VSUBS 0.008353f
C595 B.n239 VSUBS 0.008353f
C596 B.n240 VSUBS 0.008353f
C597 B.n241 VSUBS 0.008353f
C598 B.n242 VSUBS 0.008353f
C599 B.n243 VSUBS 0.008353f
C600 B.n244 VSUBS 0.008353f
C601 B.n245 VSUBS 0.008353f
C602 B.n246 VSUBS 0.008353f
C603 B.n247 VSUBS 0.008353f
C604 B.n248 VSUBS 0.008353f
C605 B.n249 VSUBS 0.008353f
C606 B.n250 VSUBS 0.008353f
C607 B.n251 VSUBS 0.008353f
C608 B.n252 VSUBS 0.008353f
C609 B.n253 VSUBS 0.008353f
C610 B.n254 VSUBS 0.008353f
C611 B.n255 VSUBS 0.008353f
C612 B.n256 VSUBS 0.008353f
C613 B.n257 VSUBS 0.008353f
C614 B.n258 VSUBS 0.008353f
C615 B.n259 VSUBS 0.008353f
C616 B.n260 VSUBS 0.008353f
C617 B.n261 VSUBS 0.008353f
C618 B.n262 VSUBS 0.008353f
C619 B.n263 VSUBS 0.008353f
C620 B.n264 VSUBS 0.020357f
C621 B.n265 VSUBS 0.019198f
C622 B.n266 VSUBS 0.019198f
C623 B.n267 VSUBS 0.008353f
C624 B.n268 VSUBS 0.008353f
C625 B.n269 VSUBS 0.008353f
C626 B.n270 VSUBS 0.008353f
C627 B.n271 VSUBS 0.008353f
C628 B.n272 VSUBS 0.008353f
C629 B.n273 VSUBS 0.008353f
C630 B.n274 VSUBS 0.008353f
C631 B.n275 VSUBS 0.008353f
C632 B.n276 VSUBS 0.008353f
C633 B.n277 VSUBS 0.008353f
C634 B.n278 VSUBS 0.008353f
C635 B.n279 VSUBS 0.008353f
C636 B.n280 VSUBS 0.008353f
C637 B.n281 VSUBS 0.008353f
C638 B.n282 VSUBS 0.008353f
C639 B.n283 VSUBS 0.008353f
C640 B.n284 VSUBS 0.008353f
C641 B.n285 VSUBS 0.008353f
C642 B.n286 VSUBS 0.008353f
C643 B.n287 VSUBS 0.008353f
C644 B.n288 VSUBS 0.008353f
C645 B.n289 VSUBS 0.008353f
C646 B.n290 VSUBS 0.008353f
C647 B.n291 VSUBS 0.008353f
C648 B.n292 VSUBS 0.008353f
C649 B.n293 VSUBS 0.008353f
C650 B.n294 VSUBS 0.008353f
C651 B.n295 VSUBS 0.008353f
C652 B.n296 VSUBS 0.008353f
C653 B.n297 VSUBS 0.008353f
C654 B.n298 VSUBS 0.008353f
C655 B.n299 VSUBS 0.008353f
C656 B.n300 VSUBS 0.008353f
C657 B.n301 VSUBS 0.008353f
C658 B.n302 VSUBS 0.008353f
C659 B.n303 VSUBS 0.008353f
C660 B.n304 VSUBS 0.008353f
C661 B.n305 VSUBS 0.008353f
C662 B.n306 VSUBS 0.008353f
C663 B.n307 VSUBS 0.008353f
C664 B.n308 VSUBS 0.008353f
C665 B.n309 VSUBS 0.008353f
C666 B.n310 VSUBS 0.008353f
C667 B.n311 VSUBS 0.008353f
C668 B.n312 VSUBS 0.008353f
C669 B.n313 VSUBS 0.008353f
C670 B.n314 VSUBS 0.008353f
C671 B.n315 VSUBS 0.008353f
C672 B.n316 VSUBS 0.008353f
C673 B.n317 VSUBS 0.008353f
C674 B.n318 VSUBS 0.008353f
C675 B.n319 VSUBS 0.008353f
C676 B.n320 VSUBS 0.008353f
C677 B.n321 VSUBS 0.008353f
C678 B.n322 VSUBS 0.008353f
C679 B.n323 VSUBS 0.008353f
C680 B.n324 VSUBS 0.008353f
C681 B.n325 VSUBS 0.008353f
C682 B.n326 VSUBS 0.008353f
C683 B.n327 VSUBS 0.008353f
C684 B.n328 VSUBS 0.008353f
C685 B.n329 VSUBS 0.008353f
C686 B.n330 VSUBS 0.008353f
C687 B.n331 VSUBS 0.008353f
C688 B.n332 VSUBS 0.008353f
C689 B.n333 VSUBS 0.008353f
C690 B.n334 VSUBS 0.008353f
C691 B.n335 VSUBS 0.008353f
C692 B.n336 VSUBS 0.008353f
C693 B.n337 VSUBS 0.008353f
C694 B.n338 VSUBS 0.008353f
C695 B.n339 VSUBS 0.008353f
C696 B.n340 VSUBS 0.008353f
C697 B.n341 VSUBS 0.008353f
C698 B.n342 VSUBS 0.008353f
C699 B.n343 VSUBS 0.008353f
C700 B.n344 VSUBS 0.008353f
C701 B.n345 VSUBS 0.008353f
C702 B.n346 VSUBS 0.008353f
C703 B.n347 VSUBS 0.008353f
C704 B.n348 VSUBS 0.008353f
C705 B.n349 VSUBS 0.008353f
C706 B.n350 VSUBS 0.008353f
C707 B.n351 VSUBS 0.008353f
C708 B.n352 VSUBS 0.019198f
C709 B.n353 VSUBS 0.020168f
C710 B.n354 VSUBS 0.019387f
C711 B.n355 VSUBS 0.008353f
C712 B.n356 VSUBS 0.008353f
C713 B.n357 VSUBS 0.008353f
C714 B.n358 VSUBS 0.008353f
C715 B.n359 VSUBS 0.008353f
C716 B.n360 VSUBS 0.008353f
C717 B.n361 VSUBS 0.008353f
C718 B.n362 VSUBS 0.008353f
C719 B.n363 VSUBS 0.008353f
C720 B.n364 VSUBS 0.008353f
C721 B.n365 VSUBS 0.008353f
C722 B.n366 VSUBS 0.008353f
C723 B.n367 VSUBS 0.008353f
C724 B.n368 VSUBS 0.008353f
C725 B.n369 VSUBS 0.008353f
C726 B.n370 VSUBS 0.008353f
C727 B.n371 VSUBS 0.008353f
C728 B.n372 VSUBS 0.008353f
C729 B.n373 VSUBS 0.008353f
C730 B.n374 VSUBS 0.008353f
C731 B.n375 VSUBS 0.008353f
C732 B.n376 VSUBS 0.008353f
C733 B.n377 VSUBS 0.008353f
C734 B.n378 VSUBS 0.008353f
C735 B.n379 VSUBS 0.008353f
C736 B.n380 VSUBS 0.008353f
C737 B.n381 VSUBS 0.008353f
C738 B.n382 VSUBS 0.008353f
C739 B.n383 VSUBS 0.008353f
C740 B.n384 VSUBS 0.008353f
C741 B.n385 VSUBS 0.008353f
C742 B.n386 VSUBS 0.008353f
C743 B.n387 VSUBS 0.008353f
C744 B.n388 VSUBS 0.008353f
C745 B.n389 VSUBS 0.008353f
C746 B.n390 VSUBS 0.008353f
C747 B.n391 VSUBS 0.005774f
C748 B.n392 VSUBS 0.008353f
C749 B.n393 VSUBS 0.008353f
C750 B.n394 VSUBS 0.006756f
C751 B.n395 VSUBS 0.008353f
C752 B.n396 VSUBS 0.008353f
C753 B.n397 VSUBS 0.008353f
C754 B.n398 VSUBS 0.008353f
C755 B.n399 VSUBS 0.008353f
C756 B.n400 VSUBS 0.008353f
C757 B.n401 VSUBS 0.008353f
C758 B.n402 VSUBS 0.008353f
C759 B.n403 VSUBS 0.008353f
C760 B.n404 VSUBS 0.008353f
C761 B.n405 VSUBS 0.008353f
C762 B.n406 VSUBS 0.006756f
C763 B.n407 VSUBS 0.019353f
C764 B.n408 VSUBS 0.005774f
C765 B.n409 VSUBS 0.008353f
C766 B.n410 VSUBS 0.008353f
C767 B.n411 VSUBS 0.008353f
C768 B.n412 VSUBS 0.008353f
C769 B.n413 VSUBS 0.008353f
C770 B.n414 VSUBS 0.008353f
C771 B.n415 VSUBS 0.008353f
C772 B.n416 VSUBS 0.008353f
C773 B.n417 VSUBS 0.008353f
C774 B.n418 VSUBS 0.008353f
C775 B.n419 VSUBS 0.008353f
C776 B.n420 VSUBS 0.008353f
C777 B.n421 VSUBS 0.008353f
C778 B.n422 VSUBS 0.008353f
C779 B.n423 VSUBS 0.008353f
C780 B.n424 VSUBS 0.008353f
C781 B.n425 VSUBS 0.008353f
C782 B.n426 VSUBS 0.008353f
C783 B.n427 VSUBS 0.008353f
C784 B.n428 VSUBS 0.008353f
C785 B.n429 VSUBS 0.008353f
C786 B.n430 VSUBS 0.008353f
C787 B.n431 VSUBS 0.008353f
C788 B.n432 VSUBS 0.008353f
C789 B.n433 VSUBS 0.008353f
C790 B.n434 VSUBS 0.008353f
C791 B.n435 VSUBS 0.008353f
C792 B.n436 VSUBS 0.008353f
C793 B.n437 VSUBS 0.008353f
C794 B.n438 VSUBS 0.008353f
C795 B.n439 VSUBS 0.008353f
C796 B.n440 VSUBS 0.008353f
C797 B.n441 VSUBS 0.008353f
C798 B.n442 VSUBS 0.008353f
C799 B.n443 VSUBS 0.008353f
C800 B.n444 VSUBS 0.008353f
C801 B.n445 VSUBS 0.020357f
C802 B.n446 VSUBS 0.020357f
C803 B.n447 VSUBS 0.019198f
C804 B.n448 VSUBS 0.008353f
C805 B.n449 VSUBS 0.008353f
C806 B.n450 VSUBS 0.008353f
C807 B.n451 VSUBS 0.008353f
C808 B.n452 VSUBS 0.008353f
C809 B.n453 VSUBS 0.008353f
C810 B.n454 VSUBS 0.008353f
C811 B.n455 VSUBS 0.008353f
C812 B.n456 VSUBS 0.008353f
C813 B.n457 VSUBS 0.008353f
C814 B.n458 VSUBS 0.008353f
C815 B.n459 VSUBS 0.008353f
C816 B.n460 VSUBS 0.008353f
C817 B.n461 VSUBS 0.008353f
C818 B.n462 VSUBS 0.008353f
C819 B.n463 VSUBS 0.008353f
C820 B.n464 VSUBS 0.008353f
C821 B.n465 VSUBS 0.008353f
C822 B.n466 VSUBS 0.008353f
C823 B.n467 VSUBS 0.008353f
C824 B.n468 VSUBS 0.008353f
C825 B.n469 VSUBS 0.008353f
C826 B.n470 VSUBS 0.008353f
C827 B.n471 VSUBS 0.008353f
C828 B.n472 VSUBS 0.008353f
C829 B.n473 VSUBS 0.008353f
C830 B.n474 VSUBS 0.008353f
C831 B.n475 VSUBS 0.008353f
C832 B.n476 VSUBS 0.008353f
C833 B.n477 VSUBS 0.008353f
C834 B.n478 VSUBS 0.008353f
C835 B.n479 VSUBS 0.008353f
C836 B.n480 VSUBS 0.008353f
C837 B.n481 VSUBS 0.008353f
C838 B.n482 VSUBS 0.008353f
C839 B.n483 VSUBS 0.008353f
C840 B.n484 VSUBS 0.008353f
C841 B.n485 VSUBS 0.008353f
C842 B.n486 VSUBS 0.008353f
C843 B.n487 VSUBS 0.008353f
C844 B.n488 VSUBS 0.008353f
C845 B.n489 VSUBS 0.008353f
C846 B.n490 VSUBS 0.008353f
C847 B.n491 VSUBS 0.018915f
.ends

