* NGSPICE file created from diff_pair_sample_0752.ext - technology: sky130A

.subckt diff_pair_sample_0752 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=2.3199 ps=14.39 w=14.06 l=2.04
X1 VDD1.t1 VP.t1 VTAIL.t14 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=5.4834 ps=28.9 w=14.06 l=2.04
X2 VTAIL.t13 VP.t2 VDD1.t0 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X3 VTAIL.t4 VN.t0 VDD2.t7 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=2.3199 ps=14.39 w=14.06 l=2.04
X4 VTAIL.t6 VN.t1 VDD2.t6 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=2.3199 ps=14.39 w=14.06 l=2.04
X5 VDD2.t5 VN.t2 VTAIL.t0 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X6 B.t11 B.t9 B.t10 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=0 ps=0 w=14.06 l=2.04
X7 VDD1.t7 VP.t3 VTAIL.t12 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X8 VDD2.t4 VN.t3 VTAIL.t5 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=5.4834 ps=28.9 w=14.06 l=2.04
X9 VTAIL.t7 VN.t4 VDD2.t3 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X10 B.t8 B.t6 B.t7 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=0 ps=0 w=14.06 l=2.04
X11 B.t5 B.t3 B.t4 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=0 ps=0 w=14.06 l=2.04
X12 VDD2.t2 VN.t5 VTAIL.t1 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=5.4834 ps=28.9 w=14.06 l=2.04
X13 VTAIL.t11 VP.t4 VDD1.t6 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=2.3199 ps=14.39 w=14.06 l=2.04
X14 VDD1.t2 VP.t5 VTAIL.t10 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=5.4834 ps=28.9 w=14.06 l=2.04
X15 VTAIL.t2 VN.t6 VDD2.t1 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X16 VTAIL.t9 VP.t6 VDD1.t4 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X17 VDD2.t0 VN.t7 VTAIL.t3 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
X18 B.t2 B.t0 B.t1 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=5.4834 pd=28.9 as=0 ps=0 w=14.06 l=2.04
X19 VDD1.t5 VP.t7 VTAIL.t8 w_n3340_n3780# sky130_fd_pr__pfet_01v8 ad=2.3199 pd=14.39 as=2.3199 ps=14.39 w=14.06 l=2.04
R0 VP.n13 VP.t4 199.073
R1 VP.n7 VP.t0 166.101
R2 VP.n40 VP.t7 166.101
R3 VP.n47 VP.t6 166.101
R4 VP.n55 VP.t5 166.101
R5 VP.n29 VP.t1 166.101
R6 VP.n21 VP.t2 166.101
R7 VP.n14 VP.t3 166.101
R8 VP.n15 VP.n12 161.3
R9 VP.n17 VP.n16 161.3
R10 VP.n18 VP.n11 161.3
R11 VP.n20 VP.n19 161.3
R12 VP.n22 VP.n10 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n25 VP.n9 161.3
R15 VP.n27 VP.n26 161.3
R16 VP.n28 VP.n8 161.3
R17 VP.n54 VP.n0 161.3
R18 VP.n53 VP.n52 161.3
R19 VP.n51 VP.n1 161.3
R20 VP.n50 VP.n49 161.3
R21 VP.n48 VP.n2 161.3
R22 VP.n46 VP.n45 161.3
R23 VP.n44 VP.n3 161.3
R24 VP.n43 VP.n42 161.3
R25 VP.n41 VP.n4 161.3
R26 VP.n39 VP.n38 161.3
R27 VP.n37 VP.n5 161.3
R28 VP.n36 VP.n35 161.3
R29 VP.n34 VP.n6 161.3
R30 VP.n33 VP.n32 161.3
R31 VP.n31 VP.n7 95.7567
R32 VP.n56 VP.n55 95.7567
R33 VP.n30 VP.n29 95.7567
R34 VP.n42 VP.n3 56.4773
R35 VP.n16 VP.n11 56.4773
R36 VP.n35 VP.n34 52.0954
R37 VP.n53 VP.n1 52.0954
R38 VP.n27 VP.n9 52.0954
R39 VP.n31 VP.n30 49.795
R40 VP.n14 VP.n13 49.1578
R41 VP.n35 VP.n5 28.7258
R42 VP.n49 VP.n1 28.7258
R43 VP.n23 VP.n9 28.7258
R44 VP.n34 VP.n33 24.3439
R45 VP.n39 VP.n5 24.3439
R46 VP.n42 VP.n41 24.3439
R47 VP.n46 VP.n3 24.3439
R48 VP.n49 VP.n48 24.3439
R49 VP.n54 VP.n53 24.3439
R50 VP.n28 VP.n27 24.3439
R51 VP.n20 VP.n11 24.3439
R52 VP.n23 VP.n22 24.3439
R53 VP.n16 VP.n15 24.3439
R54 VP.n41 VP.n40 21.1793
R55 VP.n47 VP.n46 21.1793
R56 VP.n21 VP.n20 21.1793
R57 VP.n15 VP.n14 21.1793
R58 VP.n33 VP.n7 14.85
R59 VP.n55 VP.n54 14.85
R60 VP.n29 VP.n28 14.85
R61 VP.n13 VP.n12 9.46412
R62 VP.n40 VP.n39 3.16515
R63 VP.n48 VP.n47 3.16515
R64 VP.n22 VP.n21 3.16515
R65 VP.n30 VP.n8 0.278398
R66 VP.n32 VP.n31 0.278398
R67 VP.n56 VP.n0 0.278398
R68 VP.n17 VP.n12 0.189894
R69 VP.n18 VP.n17 0.189894
R70 VP.n19 VP.n18 0.189894
R71 VP.n19 VP.n10 0.189894
R72 VP.n24 VP.n10 0.189894
R73 VP.n25 VP.n24 0.189894
R74 VP.n26 VP.n25 0.189894
R75 VP.n26 VP.n8 0.189894
R76 VP.n32 VP.n6 0.189894
R77 VP.n36 VP.n6 0.189894
R78 VP.n37 VP.n36 0.189894
R79 VP.n38 VP.n37 0.189894
R80 VP.n38 VP.n4 0.189894
R81 VP.n43 VP.n4 0.189894
R82 VP.n44 VP.n43 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n45 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VP VP.n56 0.153422
R90 VDD1 VDD1.n0 75.1292
R91 VDD1.n3 VDD1.n2 75.0155
R92 VDD1.n3 VDD1.n1 75.0155
R93 VDD1.n5 VDD1.n4 74.0493
R94 VDD1.n5 VDD1.n3 45.613
R95 VDD1.n4 VDD1.t0 2.31238
R96 VDD1.n4 VDD1.t1 2.31238
R97 VDD1.n0 VDD1.t6 2.31238
R98 VDD1.n0 VDD1.t7 2.31238
R99 VDD1.n2 VDD1.t4 2.31238
R100 VDD1.n2 VDD1.t2 2.31238
R101 VDD1.n1 VDD1.t3 2.31238
R102 VDD1.n1 VDD1.t5 2.31238
R103 VDD1 VDD1.n5 0.963862
R104 VTAIL.n626 VTAIL.n554 756.745
R105 VTAIL.n74 VTAIL.n2 756.745
R106 VTAIL.n152 VTAIL.n80 756.745
R107 VTAIL.n232 VTAIL.n160 756.745
R108 VTAIL.n548 VTAIL.n476 756.745
R109 VTAIL.n468 VTAIL.n396 756.745
R110 VTAIL.n390 VTAIL.n318 756.745
R111 VTAIL.n310 VTAIL.n238 756.745
R112 VTAIL.n578 VTAIL.n577 585
R113 VTAIL.n583 VTAIL.n582 585
R114 VTAIL.n585 VTAIL.n584 585
R115 VTAIL.n574 VTAIL.n573 585
R116 VTAIL.n591 VTAIL.n590 585
R117 VTAIL.n593 VTAIL.n592 585
R118 VTAIL.n570 VTAIL.n569 585
R119 VTAIL.n599 VTAIL.n598 585
R120 VTAIL.n601 VTAIL.n600 585
R121 VTAIL.n566 VTAIL.n565 585
R122 VTAIL.n607 VTAIL.n606 585
R123 VTAIL.n609 VTAIL.n608 585
R124 VTAIL.n562 VTAIL.n561 585
R125 VTAIL.n615 VTAIL.n614 585
R126 VTAIL.n617 VTAIL.n616 585
R127 VTAIL.n558 VTAIL.n557 585
R128 VTAIL.n624 VTAIL.n623 585
R129 VTAIL.n625 VTAIL.n556 585
R130 VTAIL.n627 VTAIL.n626 585
R131 VTAIL.n26 VTAIL.n25 585
R132 VTAIL.n31 VTAIL.n30 585
R133 VTAIL.n33 VTAIL.n32 585
R134 VTAIL.n22 VTAIL.n21 585
R135 VTAIL.n39 VTAIL.n38 585
R136 VTAIL.n41 VTAIL.n40 585
R137 VTAIL.n18 VTAIL.n17 585
R138 VTAIL.n47 VTAIL.n46 585
R139 VTAIL.n49 VTAIL.n48 585
R140 VTAIL.n14 VTAIL.n13 585
R141 VTAIL.n55 VTAIL.n54 585
R142 VTAIL.n57 VTAIL.n56 585
R143 VTAIL.n10 VTAIL.n9 585
R144 VTAIL.n63 VTAIL.n62 585
R145 VTAIL.n65 VTAIL.n64 585
R146 VTAIL.n6 VTAIL.n5 585
R147 VTAIL.n72 VTAIL.n71 585
R148 VTAIL.n73 VTAIL.n4 585
R149 VTAIL.n75 VTAIL.n74 585
R150 VTAIL.n104 VTAIL.n103 585
R151 VTAIL.n109 VTAIL.n108 585
R152 VTAIL.n111 VTAIL.n110 585
R153 VTAIL.n100 VTAIL.n99 585
R154 VTAIL.n117 VTAIL.n116 585
R155 VTAIL.n119 VTAIL.n118 585
R156 VTAIL.n96 VTAIL.n95 585
R157 VTAIL.n125 VTAIL.n124 585
R158 VTAIL.n127 VTAIL.n126 585
R159 VTAIL.n92 VTAIL.n91 585
R160 VTAIL.n133 VTAIL.n132 585
R161 VTAIL.n135 VTAIL.n134 585
R162 VTAIL.n88 VTAIL.n87 585
R163 VTAIL.n141 VTAIL.n140 585
R164 VTAIL.n143 VTAIL.n142 585
R165 VTAIL.n84 VTAIL.n83 585
R166 VTAIL.n150 VTAIL.n149 585
R167 VTAIL.n151 VTAIL.n82 585
R168 VTAIL.n153 VTAIL.n152 585
R169 VTAIL.n184 VTAIL.n183 585
R170 VTAIL.n189 VTAIL.n188 585
R171 VTAIL.n191 VTAIL.n190 585
R172 VTAIL.n180 VTAIL.n179 585
R173 VTAIL.n197 VTAIL.n196 585
R174 VTAIL.n199 VTAIL.n198 585
R175 VTAIL.n176 VTAIL.n175 585
R176 VTAIL.n205 VTAIL.n204 585
R177 VTAIL.n207 VTAIL.n206 585
R178 VTAIL.n172 VTAIL.n171 585
R179 VTAIL.n213 VTAIL.n212 585
R180 VTAIL.n215 VTAIL.n214 585
R181 VTAIL.n168 VTAIL.n167 585
R182 VTAIL.n221 VTAIL.n220 585
R183 VTAIL.n223 VTAIL.n222 585
R184 VTAIL.n164 VTAIL.n163 585
R185 VTAIL.n230 VTAIL.n229 585
R186 VTAIL.n231 VTAIL.n162 585
R187 VTAIL.n233 VTAIL.n232 585
R188 VTAIL.n549 VTAIL.n548 585
R189 VTAIL.n547 VTAIL.n478 585
R190 VTAIL.n546 VTAIL.n545 585
R191 VTAIL.n481 VTAIL.n479 585
R192 VTAIL.n540 VTAIL.n539 585
R193 VTAIL.n538 VTAIL.n537 585
R194 VTAIL.n485 VTAIL.n484 585
R195 VTAIL.n532 VTAIL.n531 585
R196 VTAIL.n530 VTAIL.n529 585
R197 VTAIL.n489 VTAIL.n488 585
R198 VTAIL.n524 VTAIL.n523 585
R199 VTAIL.n522 VTAIL.n521 585
R200 VTAIL.n493 VTAIL.n492 585
R201 VTAIL.n516 VTAIL.n515 585
R202 VTAIL.n514 VTAIL.n513 585
R203 VTAIL.n497 VTAIL.n496 585
R204 VTAIL.n508 VTAIL.n507 585
R205 VTAIL.n506 VTAIL.n505 585
R206 VTAIL.n501 VTAIL.n500 585
R207 VTAIL.n469 VTAIL.n468 585
R208 VTAIL.n467 VTAIL.n398 585
R209 VTAIL.n466 VTAIL.n465 585
R210 VTAIL.n401 VTAIL.n399 585
R211 VTAIL.n460 VTAIL.n459 585
R212 VTAIL.n458 VTAIL.n457 585
R213 VTAIL.n405 VTAIL.n404 585
R214 VTAIL.n452 VTAIL.n451 585
R215 VTAIL.n450 VTAIL.n449 585
R216 VTAIL.n409 VTAIL.n408 585
R217 VTAIL.n444 VTAIL.n443 585
R218 VTAIL.n442 VTAIL.n441 585
R219 VTAIL.n413 VTAIL.n412 585
R220 VTAIL.n436 VTAIL.n435 585
R221 VTAIL.n434 VTAIL.n433 585
R222 VTAIL.n417 VTAIL.n416 585
R223 VTAIL.n428 VTAIL.n427 585
R224 VTAIL.n426 VTAIL.n425 585
R225 VTAIL.n421 VTAIL.n420 585
R226 VTAIL.n391 VTAIL.n390 585
R227 VTAIL.n389 VTAIL.n320 585
R228 VTAIL.n388 VTAIL.n387 585
R229 VTAIL.n323 VTAIL.n321 585
R230 VTAIL.n382 VTAIL.n381 585
R231 VTAIL.n380 VTAIL.n379 585
R232 VTAIL.n327 VTAIL.n326 585
R233 VTAIL.n374 VTAIL.n373 585
R234 VTAIL.n372 VTAIL.n371 585
R235 VTAIL.n331 VTAIL.n330 585
R236 VTAIL.n366 VTAIL.n365 585
R237 VTAIL.n364 VTAIL.n363 585
R238 VTAIL.n335 VTAIL.n334 585
R239 VTAIL.n358 VTAIL.n357 585
R240 VTAIL.n356 VTAIL.n355 585
R241 VTAIL.n339 VTAIL.n338 585
R242 VTAIL.n350 VTAIL.n349 585
R243 VTAIL.n348 VTAIL.n347 585
R244 VTAIL.n343 VTAIL.n342 585
R245 VTAIL.n311 VTAIL.n310 585
R246 VTAIL.n309 VTAIL.n240 585
R247 VTAIL.n308 VTAIL.n307 585
R248 VTAIL.n243 VTAIL.n241 585
R249 VTAIL.n302 VTAIL.n301 585
R250 VTAIL.n300 VTAIL.n299 585
R251 VTAIL.n247 VTAIL.n246 585
R252 VTAIL.n294 VTAIL.n293 585
R253 VTAIL.n292 VTAIL.n291 585
R254 VTAIL.n251 VTAIL.n250 585
R255 VTAIL.n286 VTAIL.n285 585
R256 VTAIL.n284 VTAIL.n283 585
R257 VTAIL.n255 VTAIL.n254 585
R258 VTAIL.n278 VTAIL.n277 585
R259 VTAIL.n276 VTAIL.n275 585
R260 VTAIL.n259 VTAIL.n258 585
R261 VTAIL.n270 VTAIL.n269 585
R262 VTAIL.n268 VTAIL.n267 585
R263 VTAIL.n263 VTAIL.n262 585
R264 VTAIL.n579 VTAIL.t1 327.466
R265 VTAIL.n27 VTAIL.t4 327.466
R266 VTAIL.n105 VTAIL.t10 327.466
R267 VTAIL.n185 VTAIL.t15 327.466
R268 VTAIL.n502 VTAIL.t14 327.466
R269 VTAIL.n422 VTAIL.t11 327.466
R270 VTAIL.n344 VTAIL.t5 327.466
R271 VTAIL.n264 VTAIL.t6 327.466
R272 VTAIL.n583 VTAIL.n577 171.744
R273 VTAIL.n584 VTAIL.n583 171.744
R274 VTAIL.n584 VTAIL.n573 171.744
R275 VTAIL.n591 VTAIL.n573 171.744
R276 VTAIL.n592 VTAIL.n591 171.744
R277 VTAIL.n592 VTAIL.n569 171.744
R278 VTAIL.n599 VTAIL.n569 171.744
R279 VTAIL.n600 VTAIL.n599 171.744
R280 VTAIL.n600 VTAIL.n565 171.744
R281 VTAIL.n607 VTAIL.n565 171.744
R282 VTAIL.n608 VTAIL.n607 171.744
R283 VTAIL.n608 VTAIL.n561 171.744
R284 VTAIL.n615 VTAIL.n561 171.744
R285 VTAIL.n616 VTAIL.n615 171.744
R286 VTAIL.n616 VTAIL.n557 171.744
R287 VTAIL.n624 VTAIL.n557 171.744
R288 VTAIL.n625 VTAIL.n624 171.744
R289 VTAIL.n626 VTAIL.n625 171.744
R290 VTAIL.n31 VTAIL.n25 171.744
R291 VTAIL.n32 VTAIL.n31 171.744
R292 VTAIL.n32 VTAIL.n21 171.744
R293 VTAIL.n39 VTAIL.n21 171.744
R294 VTAIL.n40 VTAIL.n39 171.744
R295 VTAIL.n40 VTAIL.n17 171.744
R296 VTAIL.n47 VTAIL.n17 171.744
R297 VTAIL.n48 VTAIL.n47 171.744
R298 VTAIL.n48 VTAIL.n13 171.744
R299 VTAIL.n55 VTAIL.n13 171.744
R300 VTAIL.n56 VTAIL.n55 171.744
R301 VTAIL.n56 VTAIL.n9 171.744
R302 VTAIL.n63 VTAIL.n9 171.744
R303 VTAIL.n64 VTAIL.n63 171.744
R304 VTAIL.n64 VTAIL.n5 171.744
R305 VTAIL.n72 VTAIL.n5 171.744
R306 VTAIL.n73 VTAIL.n72 171.744
R307 VTAIL.n74 VTAIL.n73 171.744
R308 VTAIL.n109 VTAIL.n103 171.744
R309 VTAIL.n110 VTAIL.n109 171.744
R310 VTAIL.n110 VTAIL.n99 171.744
R311 VTAIL.n117 VTAIL.n99 171.744
R312 VTAIL.n118 VTAIL.n117 171.744
R313 VTAIL.n118 VTAIL.n95 171.744
R314 VTAIL.n125 VTAIL.n95 171.744
R315 VTAIL.n126 VTAIL.n125 171.744
R316 VTAIL.n126 VTAIL.n91 171.744
R317 VTAIL.n133 VTAIL.n91 171.744
R318 VTAIL.n134 VTAIL.n133 171.744
R319 VTAIL.n134 VTAIL.n87 171.744
R320 VTAIL.n141 VTAIL.n87 171.744
R321 VTAIL.n142 VTAIL.n141 171.744
R322 VTAIL.n142 VTAIL.n83 171.744
R323 VTAIL.n150 VTAIL.n83 171.744
R324 VTAIL.n151 VTAIL.n150 171.744
R325 VTAIL.n152 VTAIL.n151 171.744
R326 VTAIL.n189 VTAIL.n183 171.744
R327 VTAIL.n190 VTAIL.n189 171.744
R328 VTAIL.n190 VTAIL.n179 171.744
R329 VTAIL.n197 VTAIL.n179 171.744
R330 VTAIL.n198 VTAIL.n197 171.744
R331 VTAIL.n198 VTAIL.n175 171.744
R332 VTAIL.n205 VTAIL.n175 171.744
R333 VTAIL.n206 VTAIL.n205 171.744
R334 VTAIL.n206 VTAIL.n171 171.744
R335 VTAIL.n213 VTAIL.n171 171.744
R336 VTAIL.n214 VTAIL.n213 171.744
R337 VTAIL.n214 VTAIL.n167 171.744
R338 VTAIL.n221 VTAIL.n167 171.744
R339 VTAIL.n222 VTAIL.n221 171.744
R340 VTAIL.n222 VTAIL.n163 171.744
R341 VTAIL.n230 VTAIL.n163 171.744
R342 VTAIL.n231 VTAIL.n230 171.744
R343 VTAIL.n232 VTAIL.n231 171.744
R344 VTAIL.n548 VTAIL.n547 171.744
R345 VTAIL.n547 VTAIL.n546 171.744
R346 VTAIL.n546 VTAIL.n479 171.744
R347 VTAIL.n539 VTAIL.n479 171.744
R348 VTAIL.n539 VTAIL.n538 171.744
R349 VTAIL.n538 VTAIL.n484 171.744
R350 VTAIL.n531 VTAIL.n484 171.744
R351 VTAIL.n531 VTAIL.n530 171.744
R352 VTAIL.n530 VTAIL.n488 171.744
R353 VTAIL.n523 VTAIL.n488 171.744
R354 VTAIL.n523 VTAIL.n522 171.744
R355 VTAIL.n522 VTAIL.n492 171.744
R356 VTAIL.n515 VTAIL.n492 171.744
R357 VTAIL.n515 VTAIL.n514 171.744
R358 VTAIL.n514 VTAIL.n496 171.744
R359 VTAIL.n507 VTAIL.n496 171.744
R360 VTAIL.n507 VTAIL.n506 171.744
R361 VTAIL.n506 VTAIL.n500 171.744
R362 VTAIL.n468 VTAIL.n467 171.744
R363 VTAIL.n467 VTAIL.n466 171.744
R364 VTAIL.n466 VTAIL.n399 171.744
R365 VTAIL.n459 VTAIL.n399 171.744
R366 VTAIL.n459 VTAIL.n458 171.744
R367 VTAIL.n458 VTAIL.n404 171.744
R368 VTAIL.n451 VTAIL.n404 171.744
R369 VTAIL.n451 VTAIL.n450 171.744
R370 VTAIL.n450 VTAIL.n408 171.744
R371 VTAIL.n443 VTAIL.n408 171.744
R372 VTAIL.n443 VTAIL.n442 171.744
R373 VTAIL.n442 VTAIL.n412 171.744
R374 VTAIL.n435 VTAIL.n412 171.744
R375 VTAIL.n435 VTAIL.n434 171.744
R376 VTAIL.n434 VTAIL.n416 171.744
R377 VTAIL.n427 VTAIL.n416 171.744
R378 VTAIL.n427 VTAIL.n426 171.744
R379 VTAIL.n426 VTAIL.n420 171.744
R380 VTAIL.n390 VTAIL.n389 171.744
R381 VTAIL.n389 VTAIL.n388 171.744
R382 VTAIL.n388 VTAIL.n321 171.744
R383 VTAIL.n381 VTAIL.n321 171.744
R384 VTAIL.n381 VTAIL.n380 171.744
R385 VTAIL.n380 VTAIL.n326 171.744
R386 VTAIL.n373 VTAIL.n326 171.744
R387 VTAIL.n373 VTAIL.n372 171.744
R388 VTAIL.n372 VTAIL.n330 171.744
R389 VTAIL.n365 VTAIL.n330 171.744
R390 VTAIL.n365 VTAIL.n364 171.744
R391 VTAIL.n364 VTAIL.n334 171.744
R392 VTAIL.n357 VTAIL.n334 171.744
R393 VTAIL.n357 VTAIL.n356 171.744
R394 VTAIL.n356 VTAIL.n338 171.744
R395 VTAIL.n349 VTAIL.n338 171.744
R396 VTAIL.n349 VTAIL.n348 171.744
R397 VTAIL.n348 VTAIL.n342 171.744
R398 VTAIL.n310 VTAIL.n309 171.744
R399 VTAIL.n309 VTAIL.n308 171.744
R400 VTAIL.n308 VTAIL.n241 171.744
R401 VTAIL.n301 VTAIL.n241 171.744
R402 VTAIL.n301 VTAIL.n300 171.744
R403 VTAIL.n300 VTAIL.n246 171.744
R404 VTAIL.n293 VTAIL.n246 171.744
R405 VTAIL.n293 VTAIL.n292 171.744
R406 VTAIL.n292 VTAIL.n250 171.744
R407 VTAIL.n285 VTAIL.n250 171.744
R408 VTAIL.n285 VTAIL.n284 171.744
R409 VTAIL.n284 VTAIL.n254 171.744
R410 VTAIL.n277 VTAIL.n254 171.744
R411 VTAIL.n277 VTAIL.n276 171.744
R412 VTAIL.n276 VTAIL.n258 171.744
R413 VTAIL.n269 VTAIL.n258 171.744
R414 VTAIL.n269 VTAIL.n268 171.744
R415 VTAIL.n268 VTAIL.n262 171.744
R416 VTAIL.t1 VTAIL.n577 85.8723
R417 VTAIL.t4 VTAIL.n25 85.8723
R418 VTAIL.t10 VTAIL.n103 85.8723
R419 VTAIL.t15 VTAIL.n183 85.8723
R420 VTAIL.t14 VTAIL.n500 85.8723
R421 VTAIL.t11 VTAIL.n420 85.8723
R422 VTAIL.t5 VTAIL.n342 85.8723
R423 VTAIL.t6 VTAIL.n262 85.8723
R424 VTAIL.n475 VTAIL.n474 57.3707
R425 VTAIL.n317 VTAIL.n316 57.3707
R426 VTAIL.n1 VTAIL.n0 57.3705
R427 VTAIL.n159 VTAIL.n158 57.3705
R428 VTAIL.n631 VTAIL.n630 34.9005
R429 VTAIL.n79 VTAIL.n78 34.9005
R430 VTAIL.n157 VTAIL.n156 34.9005
R431 VTAIL.n237 VTAIL.n236 34.9005
R432 VTAIL.n553 VTAIL.n552 34.9005
R433 VTAIL.n473 VTAIL.n472 34.9005
R434 VTAIL.n395 VTAIL.n394 34.9005
R435 VTAIL.n315 VTAIL.n314 34.9005
R436 VTAIL.n631 VTAIL.n553 26.5307
R437 VTAIL.n315 VTAIL.n237 26.5307
R438 VTAIL.n579 VTAIL.n578 16.3895
R439 VTAIL.n27 VTAIL.n26 16.3895
R440 VTAIL.n105 VTAIL.n104 16.3895
R441 VTAIL.n185 VTAIL.n184 16.3895
R442 VTAIL.n502 VTAIL.n501 16.3895
R443 VTAIL.n422 VTAIL.n421 16.3895
R444 VTAIL.n344 VTAIL.n343 16.3895
R445 VTAIL.n264 VTAIL.n263 16.3895
R446 VTAIL.n627 VTAIL.n556 13.1884
R447 VTAIL.n75 VTAIL.n4 13.1884
R448 VTAIL.n153 VTAIL.n82 13.1884
R449 VTAIL.n233 VTAIL.n162 13.1884
R450 VTAIL.n549 VTAIL.n478 13.1884
R451 VTAIL.n469 VTAIL.n398 13.1884
R452 VTAIL.n391 VTAIL.n320 13.1884
R453 VTAIL.n311 VTAIL.n240 13.1884
R454 VTAIL.n582 VTAIL.n581 12.8005
R455 VTAIL.n623 VTAIL.n622 12.8005
R456 VTAIL.n628 VTAIL.n554 12.8005
R457 VTAIL.n30 VTAIL.n29 12.8005
R458 VTAIL.n71 VTAIL.n70 12.8005
R459 VTAIL.n76 VTAIL.n2 12.8005
R460 VTAIL.n108 VTAIL.n107 12.8005
R461 VTAIL.n149 VTAIL.n148 12.8005
R462 VTAIL.n154 VTAIL.n80 12.8005
R463 VTAIL.n188 VTAIL.n187 12.8005
R464 VTAIL.n229 VTAIL.n228 12.8005
R465 VTAIL.n234 VTAIL.n160 12.8005
R466 VTAIL.n550 VTAIL.n476 12.8005
R467 VTAIL.n545 VTAIL.n480 12.8005
R468 VTAIL.n505 VTAIL.n504 12.8005
R469 VTAIL.n470 VTAIL.n396 12.8005
R470 VTAIL.n465 VTAIL.n400 12.8005
R471 VTAIL.n425 VTAIL.n424 12.8005
R472 VTAIL.n392 VTAIL.n318 12.8005
R473 VTAIL.n387 VTAIL.n322 12.8005
R474 VTAIL.n347 VTAIL.n346 12.8005
R475 VTAIL.n312 VTAIL.n238 12.8005
R476 VTAIL.n307 VTAIL.n242 12.8005
R477 VTAIL.n267 VTAIL.n266 12.8005
R478 VTAIL.n585 VTAIL.n576 12.0247
R479 VTAIL.n621 VTAIL.n558 12.0247
R480 VTAIL.n33 VTAIL.n24 12.0247
R481 VTAIL.n69 VTAIL.n6 12.0247
R482 VTAIL.n111 VTAIL.n102 12.0247
R483 VTAIL.n147 VTAIL.n84 12.0247
R484 VTAIL.n191 VTAIL.n182 12.0247
R485 VTAIL.n227 VTAIL.n164 12.0247
R486 VTAIL.n544 VTAIL.n481 12.0247
R487 VTAIL.n508 VTAIL.n499 12.0247
R488 VTAIL.n464 VTAIL.n401 12.0247
R489 VTAIL.n428 VTAIL.n419 12.0247
R490 VTAIL.n386 VTAIL.n323 12.0247
R491 VTAIL.n350 VTAIL.n341 12.0247
R492 VTAIL.n306 VTAIL.n243 12.0247
R493 VTAIL.n270 VTAIL.n261 12.0247
R494 VTAIL.n586 VTAIL.n574 11.249
R495 VTAIL.n618 VTAIL.n617 11.249
R496 VTAIL.n34 VTAIL.n22 11.249
R497 VTAIL.n66 VTAIL.n65 11.249
R498 VTAIL.n112 VTAIL.n100 11.249
R499 VTAIL.n144 VTAIL.n143 11.249
R500 VTAIL.n192 VTAIL.n180 11.249
R501 VTAIL.n224 VTAIL.n223 11.249
R502 VTAIL.n541 VTAIL.n540 11.249
R503 VTAIL.n509 VTAIL.n497 11.249
R504 VTAIL.n461 VTAIL.n460 11.249
R505 VTAIL.n429 VTAIL.n417 11.249
R506 VTAIL.n383 VTAIL.n382 11.249
R507 VTAIL.n351 VTAIL.n339 11.249
R508 VTAIL.n303 VTAIL.n302 11.249
R509 VTAIL.n271 VTAIL.n259 11.249
R510 VTAIL.n590 VTAIL.n589 10.4732
R511 VTAIL.n614 VTAIL.n560 10.4732
R512 VTAIL.n38 VTAIL.n37 10.4732
R513 VTAIL.n62 VTAIL.n8 10.4732
R514 VTAIL.n116 VTAIL.n115 10.4732
R515 VTAIL.n140 VTAIL.n86 10.4732
R516 VTAIL.n196 VTAIL.n195 10.4732
R517 VTAIL.n220 VTAIL.n166 10.4732
R518 VTAIL.n537 VTAIL.n483 10.4732
R519 VTAIL.n513 VTAIL.n512 10.4732
R520 VTAIL.n457 VTAIL.n403 10.4732
R521 VTAIL.n433 VTAIL.n432 10.4732
R522 VTAIL.n379 VTAIL.n325 10.4732
R523 VTAIL.n355 VTAIL.n354 10.4732
R524 VTAIL.n299 VTAIL.n245 10.4732
R525 VTAIL.n275 VTAIL.n274 10.4732
R526 VTAIL.n593 VTAIL.n572 9.69747
R527 VTAIL.n613 VTAIL.n562 9.69747
R528 VTAIL.n41 VTAIL.n20 9.69747
R529 VTAIL.n61 VTAIL.n10 9.69747
R530 VTAIL.n119 VTAIL.n98 9.69747
R531 VTAIL.n139 VTAIL.n88 9.69747
R532 VTAIL.n199 VTAIL.n178 9.69747
R533 VTAIL.n219 VTAIL.n168 9.69747
R534 VTAIL.n536 VTAIL.n485 9.69747
R535 VTAIL.n516 VTAIL.n495 9.69747
R536 VTAIL.n456 VTAIL.n405 9.69747
R537 VTAIL.n436 VTAIL.n415 9.69747
R538 VTAIL.n378 VTAIL.n327 9.69747
R539 VTAIL.n358 VTAIL.n337 9.69747
R540 VTAIL.n298 VTAIL.n247 9.69747
R541 VTAIL.n278 VTAIL.n257 9.69747
R542 VTAIL.n630 VTAIL.n629 9.45567
R543 VTAIL.n78 VTAIL.n77 9.45567
R544 VTAIL.n156 VTAIL.n155 9.45567
R545 VTAIL.n236 VTAIL.n235 9.45567
R546 VTAIL.n552 VTAIL.n551 9.45567
R547 VTAIL.n472 VTAIL.n471 9.45567
R548 VTAIL.n394 VTAIL.n393 9.45567
R549 VTAIL.n314 VTAIL.n313 9.45567
R550 VTAIL.n629 VTAIL.n628 9.3005
R551 VTAIL.n568 VTAIL.n567 9.3005
R552 VTAIL.n597 VTAIL.n596 9.3005
R553 VTAIL.n595 VTAIL.n594 9.3005
R554 VTAIL.n572 VTAIL.n571 9.3005
R555 VTAIL.n589 VTAIL.n588 9.3005
R556 VTAIL.n587 VTAIL.n586 9.3005
R557 VTAIL.n576 VTAIL.n575 9.3005
R558 VTAIL.n581 VTAIL.n580 9.3005
R559 VTAIL.n603 VTAIL.n602 9.3005
R560 VTAIL.n605 VTAIL.n604 9.3005
R561 VTAIL.n564 VTAIL.n563 9.3005
R562 VTAIL.n611 VTAIL.n610 9.3005
R563 VTAIL.n613 VTAIL.n612 9.3005
R564 VTAIL.n560 VTAIL.n559 9.3005
R565 VTAIL.n619 VTAIL.n618 9.3005
R566 VTAIL.n621 VTAIL.n620 9.3005
R567 VTAIL.n622 VTAIL.n555 9.3005
R568 VTAIL.n77 VTAIL.n76 9.3005
R569 VTAIL.n16 VTAIL.n15 9.3005
R570 VTAIL.n45 VTAIL.n44 9.3005
R571 VTAIL.n43 VTAIL.n42 9.3005
R572 VTAIL.n20 VTAIL.n19 9.3005
R573 VTAIL.n37 VTAIL.n36 9.3005
R574 VTAIL.n35 VTAIL.n34 9.3005
R575 VTAIL.n24 VTAIL.n23 9.3005
R576 VTAIL.n29 VTAIL.n28 9.3005
R577 VTAIL.n51 VTAIL.n50 9.3005
R578 VTAIL.n53 VTAIL.n52 9.3005
R579 VTAIL.n12 VTAIL.n11 9.3005
R580 VTAIL.n59 VTAIL.n58 9.3005
R581 VTAIL.n61 VTAIL.n60 9.3005
R582 VTAIL.n8 VTAIL.n7 9.3005
R583 VTAIL.n67 VTAIL.n66 9.3005
R584 VTAIL.n69 VTAIL.n68 9.3005
R585 VTAIL.n70 VTAIL.n3 9.3005
R586 VTAIL.n155 VTAIL.n154 9.3005
R587 VTAIL.n94 VTAIL.n93 9.3005
R588 VTAIL.n123 VTAIL.n122 9.3005
R589 VTAIL.n121 VTAIL.n120 9.3005
R590 VTAIL.n98 VTAIL.n97 9.3005
R591 VTAIL.n115 VTAIL.n114 9.3005
R592 VTAIL.n113 VTAIL.n112 9.3005
R593 VTAIL.n102 VTAIL.n101 9.3005
R594 VTAIL.n107 VTAIL.n106 9.3005
R595 VTAIL.n129 VTAIL.n128 9.3005
R596 VTAIL.n131 VTAIL.n130 9.3005
R597 VTAIL.n90 VTAIL.n89 9.3005
R598 VTAIL.n137 VTAIL.n136 9.3005
R599 VTAIL.n139 VTAIL.n138 9.3005
R600 VTAIL.n86 VTAIL.n85 9.3005
R601 VTAIL.n145 VTAIL.n144 9.3005
R602 VTAIL.n147 VTAIL.n146 9.3005
R603 VTAIL.n148 VTAIL.n81 9.3005
R604 VTAIL.n235 VTAIL.n234 9.3005
R605 VTAIL.n174 VTAIL.n173 9.3005
R606 VTAIL.n203 VTAIL.n202 9.3005
R607 VTAIL.n201 VTAIL.n200 9.3005
R608 VTAIL.n178 VTAIL.n177 9.3005
R609 VTAIL.n195 VTAIL.n194 9.3005
R610 VTAIL.n193 VTAIL.n192 9.3005
R611 VTAIL.n182 VTAIL.n181 9.3005
R612 VTAIL.n187 VTAIL.n186 9.3005
R613 VTAIL.n209 VTAIL.n208 9.3005
R614 VTAIL.n211 VTAIL.n210 9.3005
R615 VTAIL.n170 VTAIL.n169 9.3005
R616 VTAIL.n217 VTAIL.n216 9.3005
R617 VTAIL.n219 VTAIL.n218 9.3005
R618 VTAIL.n166 VTAIL.n165 9.3005
R619 VTAIL.n225 VTAIL.n224 9.3005
R620 VTAIL.n227 VTAIL.n226 9.3005
R621 VTAIL.n228 VTAIL.n161 9.3005
R622 VTAIL.n528 VTAIL.n527 9.3005
R623 VTAIL.n487 VTAIL.n486 9.3005
R624 VTAIL.n534 VTAIL.n533 9.3005
R625 VTAIL.n536 VTAIL.n535 9.3005
R626 VTAIL.n483 VTAIL.n482 9.3005
R627 VTAIL.n542 VTAIL.n541 9.3005
R628 VTAIL.n544 VTAIL.n543 9.3005
R629 VTAIL.n480 VTAIL.n477 9.3005
R630 VTAIL.n551 VTAIL.n550 9.3005
R631 VTAIL.n526 VTAIL.n525 9.3005
R632 VTAIL.n491 VTAIL.n490 9.3005
R633 VTAIL.n520 VTAIL.n519 9.3005
R634 VTAIL.n518 VTAIL.n517 9.3005
R635 VTAIL.n495 VTAIL.n494 9.3005
R636 VTAIL.n512 VTAIL.n511 9.3005
R637 VTAIL.n510 VTAIL.n509 9.3005
R638 VTAIL.n499 VTAIL.n498 9.3005
R639 VTAIL.n504 VTAIL.n503 9.3005
R640 VTAIL.n448 VTAIL.n447 9.3005
R641 VTAIL.n407 VTAIL.n406 9.3005
R642 VTAIL.n454 VTAIL.n453 9.3005
R643 VTAIL.n456 VTAIL.n455 9.3005
R644 VTAIL.n403 VTAIL.n402 9.3005
R645 VTAIL.n462 VTAIL.n461 9.3005
R646 VTAIL.n464 VTAIL.n463 9.3005
R647 VTAIL.n400 VTAIL.n397 9.3005
R648 VTAIL.n471 VTAIL.n470 9.3005
R649 VTAIL.n446 VTAIL.n445 9.3005
R650 VTAIL.n411 VTAIL.n410 9.3005
R651 VTAIL.n440 VTAIL.n439 9.3005
R652 VTAIL.n438 VTAIL.n437 9.3005
R653 VTAIL.n415 VTAIL.n414 9.3005
R654 VTAIL.n432 VTAIL.n431 9.3005
R655 VTAIL.n430 VTAIL.n429 9.3005
R656 VTAIL.n419 VTAIL.n418 9.3005
R657 VTAIL.n424 VTAIL.n423 9.3005
R658 VTAIL.n370 VTAIL.n369 9.3005
R659 VTAIL.n329 VTAIL.n328 9.3005
R660 VTAIL.n376 VTAIL.n375 9.3005
R661 VTAIL.n378 VTAIL.n377 9.3005
R662 VTAIL.n325 VTAIL.n324 9.3005
R663 VTAIL.n384 VTAIL.n383 9.3005
R664 VTAIL.n386 VTAIL.n385 9.3005
R665 VTAIL.n322 VTAIL.n319 9.3005
R666 VTAIL.n393 VTAIL.n392 9.3005
R667 VTAIL.n368 VTAIL.n367 9.3005
R668 VTAIL.n333 VTAIL.n332 9.3005
R669 VTAIL.n362 VTAIL.n361 9.3005
R670 VTAIL.n360 VTAIL.n359 9.3005
R671 VTAIL.n337 VTAIL.n336 9.3005
R672 VTAIL.n354 VTAIL.n353 9.3005
R673 VTAIL.n352 VTAIL.n351 9.3005
R674 VTAIL.n341 VTAIL.n340 9.3005
R675 VTAIL.n346 VTAIL.n345 9.3005
R676 VTAIL.n290 VTAIL.n289 9.3005
R677 VTAIL.n249 VTAIL.n248 9.3005
R678 VTAIL.n296 VTAIL.n295 9.3005
R679 VTAIL.n298 VTAIL.n297 9.3005
R680 VTAIL.n245 VTAIL.n244 9.3005
R681 VTAIL.n304 VTAIL.n303 9.3005
R682 VTAIL.n306 VTAIL.n305 9.3005
R683 VTAIL.n242 VTAIL.n239 9.3005
R684 VTAIL.n313 VTAIL.n312 9.3005
R685 VTAIL.n288 VTAIL.n287 9.3005
R686 VTAIL.n253 VTAIL.n252 9.3005
R687 VTAIL.n282 VTAIL.n281 9.3005
R688 VTAIL.n280 VTAIL.n279 9.3005
R689 VTAIL.n257 VTAIL.n256 9.3005
R690 VTAIL.n274 VTAIL.n273 9.3005
R691 VTAIL.n272 VTAIL.n271 9.3005
R692 VTAIL.n261 VTAIL.n260 9.3005
R693 VTAIL.n266 VTAIL.n265 9.3005
R694 VTAIL.n594 VTAIL.n570 8.92171
R695 VTAIL.n610 VTAIL.n609 8.92171
R696 VTAIL.n42 VTAIL.n18 8.92171
R697 VTAIL.n58 VTAIL.n57 8.92171
R698 VTAIL.n120 VTAIL.n96 8.92171
R699 VTAIL.n136 VTAIL.n135 8.92171
R700 VTAIL.n200 VTAIL.n176 8.92171
R701 VTAIL.n216 VTAIL.n215 8.92171
R702 VTAIL.n533 VTAIL.n532 8.92171
R703 VTAIL.n517 VTAIL.n493 8.92171
R704 VTAIL.n453 VTAIL.n452 8.92171
R705 VTAIL.n437 VTAIL.n413 8.92171
R706 VTAIL.n375 VTAIL.n374 8.92171
R707 VTAIL.n359 VTAIL.n335 8.92171
R708 VTAIL.n295 VTAIL.n294 8.92171
R709 VTAIL.n279 VTAIL.n255 8.92171
R710 VTAIL.n598 VTAIL.n597 8.14595
R711 VTAIL.n606 VTAIL.n564 8.14595
R712 VTAIL.n46 VTAIL.n45 8.14595
R713 VTAIL.n54 VTAIL.n12 8.14595
R714 VTAIL.n124 VTAIL.n123 8.14595
R715 VTAIL.n132 VTAIL.n90 8.14595
R716 VTAIL.n204 VTAIL.n203 8.14595
R717 VTAIL.n212 VTAIL.n170 8.14595
R718 VTAIL.n529 VTAIL.n487 8.14595
R719 VTAIL.n521 VTAIL.n520 8.14595
R720 VTAIL.n449 VTAIL.n407 8.14595
R721 VTAIL.n441 VTAIL.n440 8.14595
R722 VTAIL.n371 VTAIL.n329 8.14595
R723 VTAIL.n363 VTAIL.n362 8.14595
R724 VTAIL.n291 VTAIL.n249 8.14595
R725 VTAIL.n283 VTAIL.n282 8.14595
R726 VTAIL.n601 VTAIL.n568 7.3702
R727 VTAIL.n605 VTAIL.n566 7.3702
R728 VTAIL.n49 VTAIL.n16 7.3702
R729 VTAIL.n53 VTAIL.n14 7.3702
R730 VTAIL.n127 VTAIL.n94 7.3702
R731 VTAIL.n131 VTAIL.n92 7.3702
R732 VTAIL.n207 VTAIL.n174 7.3702
R733 VTAIL.n211 VTAIL.n172 7.3702
R734 VTAIL.n528 VTAIL.n489 7.3702
R735 VTAIL.n524 VTAIL.n491 7.3702
R736 VTAIL.n448 VTAIL.n409 7.3702
R737 VTAIL.n444 VTAIL.n411 7.3702
R738 VTAIL.n370 VTAIL.n331 7.3702
R739 VTAIL.n366 VTAIL.n333 7.3702
R740 VTAIL.n290 VTAIL.n251 7.3702
R741 VTAIL.n286 VTAIL.n253 7.3702
R742 VTAIL.n602 VTAIL.n601 6.59444
R743 VTAIL.n602 VTAIL.n566 6.59444
R744 VTAIL.n50 VTAIL.n49 6.59444
R745 VTAIL.n50 VTAIL.n14 6.59444
R746 VTAIL.n128 VTAIL.n127 6.59444
R747 VTAIL.n128 VTAIL.n92 6.59444
R748 VTAIL.n208 VTAIL.n207 6.59444
R749 VTAIL.n208 VTAIL.n172 6.59444
R750 VTAIL.n525 VTAIL.n489 6.59444
R751 VTAIL.n525 VTAIL.n524 6.59444
R752 VTAIL.n445 VTAIL.n409 6.59444
R753 VTAIL.n445 VTAIL.n444 6.59444
R754 VTAIL.n367 VTAIL.n331 6.59444
R755 VTAIL.n367 VTAIL.n366 6.59444
R756 VTAIL.n287 VTAIL.n251 6.59444
R757 VTAIL.n287 VTAIL.n286 6.59444
R758 VTAIL.n598 VTAIL.n568 5.81868
R759 VTAIL.n606 VTAIL.n605 5.81868
R760 VTAIL.n46 VTAIL.n16 5.81868
R761 VTAIL.n54 VTAIL.n53 5.81868
R762 VTAIL.n124 VTAIL.n94 5.81868
R763 VTAIL.n132 VTAIL.n131 5.81868
R764 VTAIL.n204 VTAIL.n174 5.81868
R765 VTAIL.n212 VTAIL.n211 5.81868
R766 VTAIL.n529 VTAIL.n528 5.81868
R767 VTAIL.n521 VTAIL.n491 5.81868
R768 VTAIL.n449 VTAIL.n448 5.81868
R769 VTAIL.n441 VTAIL.n411 5.81868
R770 VTAIL.n371 VTAIL.n370 5.81868
R771 VTAIL.n363 VTAIL.n333 5.81868
R772 VTAIL.n291 VTAIL.n290 5.81868
R773 VTAIL.n283 VTAIL.n253 5.81868
R774 VTAIL.n597 VTAIL.n570 5.04292
R775 VTAIL.n609 VTAIL.n564 5.04292
R776 VTAIL.n45 VTAIL.n18 5.04292
R777 VTAIL.n57 VTAIL.n12 5.04292
R778 VTAIL.n123 VTAIL.n96 5.04292
R779 VTAIL.n135 VTAIL.n90 5.04292
R780 VTAIL.n203 VTAIL.n176 5.04292
R781 VTAIL.n215 VTAIL.n170 5.04292
R782 VTAIL.n532 VTAIL.n487 5.04292
R783 VTAIL.n520 VTAIL.n493 5.04292
R784 VTAIL.n452 VTAIL.n407 5.04292
R785 VTAIL.n440 VTAIL.n413 5.04292
R786 VTAIL.n374 VTAIL.n329 5.04292
R787 VTAIL.n362 VTAIL.n335 5.04292
R788 VTAIL.n294 VTAIL.n249 5.04292
R789 VTAIL.n282 VTAIL.n255 5.04292
R790 VTAIL.n594 VTAIL.n593 4.26717
R791 VTAIL.n610 VTAIL.n562 4.26717
R792 VTAIL.n42 VTAIL.n41 4.26717
R793 VTAIL.n58 VTAIL.n10 4.26717
R794 VTAIL.n120 VTAIL.n119 4.26717
R795 VTAIL.n136 VTAIL.n88 4.26717
R796 VTAIL.n200 VTAIL.n199 4.26717
R797 VTAIL.n216 VTAIL.n168 4.26717
R798 VTAIL.n533 VTAIL.n485 4.26717
R799 VTAIL.n517 VTAIL.n516 4.26717
R800 VTAIL.n453 VTAIL.n405 4.26717
R801 VTAIL.n437 VTAIL.n436 4.26717
R802 VTAIL.n375 VTAIL.n327 4.26717
R803 VTAIL.n359 VTAIL.n358 4.26717
R804 VTAIL.n295 VTAIL.n247 4.26717
R805 VTAIL.n279 VTAIL.n278 4.26717
R806 VTAIL.n580 VTAIL.n579 3.70982
R807 VTAIL.n28 VTAIL.n27 3.70982
R808 VTAIL.n106 VTAIL.n105 3.70982
R809 VTAIL.n186 VTAIL.n185 3.70982
R810 VTAIL.n503 VTAIL.n502 3.70982
R811 VTAIL.n423 VTAIL.n422 3.70982
R812 VTAIL.n345 VTAIL.n344 3.70982
R813 VTAIL.n265 VTAIL.n264 3.70982
R814 VTAIL.n590 VTAIL.n572 3.49141
R815 VTAIL.n614 VTAIL.n613 3.49141
R816 VTAIL.n38 VTAIL.n20 3.49141
R817 VTAIL.n62 VTAIL.n61 3.49141
R818 VTAIL.n116 VTAIL.n98 3.49141
R819 VTAIL.n140 VTAIL.n139 3.49141
R820 VTAIL.n196 VTAIL.n178 3.49141
R821 VTAIL.n220 VTAIL.n219 3.49141
R822 VTAIL.n537 VTAIL.n536 3.49141
R823 VTAIL.n513 VTAIL.n495 3.49141
R824 VTAIL.n457 VTAIL.n456 3.49141
R825 VTAIL.n433 VTAIL.n415 3.49141
R826 VTAIL.n379 VTAIL.n378 3.49141
R827 VTAIL.n355 VTAIL.n337 3.49141
R828 VTAIL.n299 VTAIL.n298 3.49141
R829 VTAIL.n275 VTAIL.n257 3.49141
R830 VTAIL.n589 VTAIL.n574 2.71565
R831 VTAIL.n617 VTAIL.n560 2.71565
R832 VTAIL.n37 VTAIL.n22 2.71565
R833 VTAIL.n65 VTAIL.n8 2.71565
R834 VTAIL.n115 VTAIL.n100 2.71565
R835 VTAIL.n143 VTAIL.n86 2.71565
R836 VTAIL.n195 VTAIL.n180 2.71565
R837 VTAIL.n223 VTAIL.n166 2.71565
R838 VTAIL.n540 VTAIL.n483 2.71565
R839 VTAIL.n512 VTAIL.n497 2.71565
R840 VTAIL.n460 VTAIL.n403 2.71565
R841 VTAIL.n432 VTAIL.n417 2.71565
R842 VTAIL.n382 VTAIL.n325 2.71565
R843 VTAIL.n354 VTAIL.n339 2.71565
R844 VTAIL.n302 VTAIL.n245 2.71565
R845 VTAIL.n274 VTAIL.n259 2.71565
R846 VTAIL.n0 VTAIL.t3 2.31238
R847 VTAIL.n0 VTAIL.t2 2.31238
R848 VTAIL.n158 VTAIL.t8 2.31238
R849 VTAIL.n158 VTAIL.t9 2.31238
R850 VTAIL.n474 VTAIL.t12 2.31238
R851 VTAIL.n474 VTAIL.t13 2.31238
R852 VTAIL.n316 VTAIL.t0 2.31238
R853 VTAIL.n316 VTAIL.t7 2.31238
R854 VTAIL.n317 VTAIL.n315 2.0436
R855 VTAIL.n395 VTAIL.n317 2.0436
R856 VTAIL.n475 VTAIL.n473 2.0436
R857 VTAIL.n553 VTAIL.n475 2.0436
R858 VTAIL.n237 VTAIL.n159 2.0436
R859 VTAIL.n159 VTAIL.n157 2.0436
R860 VTAIL.n79 VTAIL.n1 2.0436
R861 VTAIL VTAIL.n631 1.98541
R862 VTAIL.n586 VTAIL.n585 1.93989
R863 VTAIL.n618 VTAIL.n558 1.93989
R864 VTAIL.n34 VTAIL.n33 1.93989
R865 VTAIL.n66 VTAIL.n6 1.93989
R866 VTAIL.n112 VTAIL.n111 1.93989
R867 VTAIL.n144 VTAIL.n84 1.93989
R868 VTAIL.n192 VTAIL.n191 1.93989
R869 VTAIL.n224 VTAIL.n164 1.93989
R870 VTAIL.n541 VTAIL.n481 1.93989
R871 VTAIL.n509 VTAIL.n508 1.93989
R872 VTAIL.n461 VTAIL.n401 1.93989
R873 VTAIL.n429 VTAIL.n428 1.93989
R874 VTAIL.n383 VTAIL.n323 1.93989
R875 VTAIL.n351 VTAIL.n350 1.93989
R876 VTAIL.n303 VTAIL.n243 1.93989
R877 VTAIL.n271 VTAIL.n270 1.93989
R878 VTAIL.n582 VTAIL.n576 1.16414
R879 VTAIL.n623 VTAIL.n621 1.16414
R880 VTAIL.n630 VTAIL.n554 1.16414
R881 VTAIL.n30 VTAIL.n24 1.16414
R882 VTAIL.n71 VTAIL.n69 1.16414
R883 VTAIL.n78 VTAIL.n2 1.16414
R884 VTAIL.n108 VTAIL.n102 1.16414
R885 VTAIL.n149 VTAIL.n147 1.16414
R886 VTAIL.n156 VTAIL.n80 1.16414
R887 VTAIL.n188 VTAIL.n182 1.16414
R888 VTAIL.n229 VTAIL.n227 1.16414
R889 VTAIL.n236 VTAIL.n160 1.16414
R890 VTAIL.n552 VTAIL.n476 1.16414
R891 VTAIL.n545 VTAIL.n544 1.16414
R892 VTAIL.n505 VTAIL.n499 1.16414
R893 VTAIL.n472 VTAIL.n396 1.16414
R894 VTAIL.n465 VTAIL.n464 1.16414
R895 VTAIL.n425 VTAIL.n419 1.16414
R896 VTAIL.n394 VTAIL.n318 1.16414
R897 VTAIL.n387 VTAIL.n386 1.16414
R898 VTAIL.n347 VTAIL.n341 1.16414
R899 VTAIL.n314 VTAIL.n238 1.16414
R900 VTAIL.n307 VTAIL.n306 1.16414
R901 VTAIL.n267 VTAIL.n261 1.16414
R902 VTAIL.n473 VTAIL.n395 0.470328
R903 VTAIL.n157 VTAIL.n79 0.470328
R904 VTAIL.n581 VTAIL.n578 0.388379
R905 VTAIL.n622 VTAIL.n556 0.388379
R906 VTAIL.n628 VTAIL.n627 0.388379
R907 VTAIL.n29 VTAIL.n26 0.388379
R908 VTAIL.n70 VTAIL.n4 0.388379
R909 VTAIL.n76 VTAIL.n75 0.388379
R910 VTAIL.n107 VTAIL.n104 0.388379
R911 VTAIL.n148 VTAIL.n82 0.388379
R912 VTAIL.n154 VTAIL.n153 0.388379
R913 VTAIL.n187 VTAIL.n184 0.388379
R914 VTAIL.n228 VTAIL.n162 0.388379
R915 VTAIL.n234 VTAIL.n233 0.388379
R916 VTAIL.n550 VTAIL.n549 0.388379
R917 VTAIL.n480 VTAIL.n478 0.388379
R918 VTAIL.n504 VTAIL.n501 0.388379
R919 VTAIL.n470 VTAIL.n469 0.388379
R920 VTAIL.n400 VTAIL.n398 0.388379
R921 VTAIL.n424 VTAIL.n421 0.388379
R922 VTAIL.n392 VTAIL.n391 0.388379
R923 VTAIL.n322 VTAIL.n320 0.388379
R924 VTAIL.n346 VTAIL.n343 0.388379
R925 VTAIL.n312 VTAIL.n311 0.388379
R926 VTAIL.n242 VTAIL.n240 0.388379
R927 VTAIL.n266 VTAIL.n263 0.388379
R928 VTAIL.n580 VTAIL.n575 0.155672
R929 VTAIL.n587 VTAIL.n575 0.155672
R930 VTAIL.n588 VTAIL.n587 0.155672
R931 VTAIL.n588 VTAIL.n571 0.155672
R932 VTAIL.n595 VTAIL.n571 0.155672
R933 VTAIL.n596 VTAIL.n595 0.155672
R934 VTAIL.n596 VTAIL.n567 0.155672
R935 VTAIL.n603 VTAIL.n567 0.155672
R936 VTAIL.n604 VTAIL.n603 0.155672
R937 VTAIL.n604 VTAIL.n563 0.155672
R938 VTAIL.n611 VTAIL.n563 0.155672
R939 VTAIL.n612 VTAIL.n611 0.155672
R940 VTAIL.n612 VTAIL.n559 0.155672
R941 VTAIL.n619 VTAIL.n559 0.155672
R942 VTAIL.n620 VTAIL.n619 0.155672
R943 VTAIL.n620 VTAIL.n555 0.155672
R944 VTAIL.n629 VTAIL.n555 0.155672
R945 VTAIL.n28 VTAIL.n23 0.155672
R946 VTAIL.n35 VTAIL.n23 0.155672
R947 VTAIL.n36 VTAIL.n35 0.155672
R948 VTAIL.n36 VTAIL.n19 0.155672
R949 VTAIL.n43 VTAIL.n19 0.155672
R950 VTAIL.n44 VTAIL.n43 0.155672
R951 VTAIL.n44 VTAIL.n15 0.155672
R952 VTAIL.n51 VTAIL.n15 0.155672
R953 VTAIL.n52 VTAIL.n51 0.155672
R954 VTAIL.n52 VTAIL.n11 0.155672
R955 VTAIL.n59 VTAIL.n11 0.155672
R956 VTAIL.n60 VTAIL.n59 0.155672
R957 VTAIL.n60 VTAIL.n7 0.155672
R958 VTAIL.n67 VTAIL.n7 0.155672
R959 VTAIL.n68 VTAIL.n67 0.155672
R960 VTAIL.n68 VTAIL.n3 0.155672
R961 VTAIL.n77 VTAIL.n3 0.155672
R962 VTAIL.n106 VTAIL.n101 0.155672
R963 VTAIL.n113 VTAIL.n101 0.155672
R964 VTAIL.n114 VTAIL.n113 0.155672
R965 VTAIL.n114 VTAIL.n97 0.155672
R966 VTAIL.n121 VTAIL.n97 0.155672
R967 VTAIL.n122 VTAIL.n121 0.155672
R968 VTAIL.n122 VTAIL.n93 0.155672
R969 VTAIL.n129 VTAIL.n93 0.155672
R970 VTAIL.n130 VTAIL.n129 0.155672
R971 VTAIL.n130 VTAIL.n89 0.155672
R972 VTAIL.n137 VTAIL.n89 0.155672
R973 VTAIL.n138 VTAIL.n137 0.155672
R974 VTAIL.n138 VTAIL.n85 0.155672
R975 VTAIL.n145 VTAIL.n85 0.155672
R976 VTAIL.n146 VTAIL.n145 0.155672
R977 VTAIL.n146 VTAIL.n81 0.155672
R978 VTAIL.n155 VTAIL.n81 0.155672
R979 VTAIL.n186 VTAIL.n181 0.155672
R980 VTAIL.n193 VTAIL.n181 0.155672
R981 VTAIL.n194 VTAIL.n193 0.155672
R982 VTAIL.n194 VTAIL.n177 0.155672
R983 VTAIL.n201 VTAIL.n177 0.155672
R984 VTAIL.n202 VTAIL.n201 0.155672
R985 VTAIL.n202 VTAIL.n173 0.155672
R986 VTAIL.n209 VTAIL.n173 0.155672
R987 VTAIL.n210 VTAIL.n209 0.155672
R988 VTAIL.n210 VTAIL.n169 0.155672
R989 VTAIL.n217 VTAIL.n169 0.155672
R990 VTAIL.n218 VTAIL.n217 0.155672
R991 VTAIL.n218 VTAIL.n165 0.155672
R992 VTAIL.n225 VTAIL.n165 0.155672
R993 VTAIL.n226 VTAIL.n225 0.155672
R994 VTAIL.n226 VTAIL.n161 0.155672
R995 VTAIL.n235 VTAIL.n161 0.155672
R996 VTAIL.n551 VTAIL.n477 0.155672
R997 VTAIL.n543 VTAIL.n477 0.155672
R998 VTAIL.n543 VTAIL.n542 0.155672
R999 VTAIL.n542 VTAIL.n482 0.155672
R1000 VTAIL.n535 VTAIL.n482 0.155672
R1001 VTAIL.n535 VTAIL.n534 0.155672
R1002 VTAIL.n534 VTAIL.n486 0.155672
R1003 VTAIL.n527 VTAIL.n486 0.155672
R1004 VTAIL.n527 VTAIL.n526 0.155672
R1005 VTAIL.n526 VTAIL.n490 0.155672
R1006 VTAIL.n519 VTAIL.n490 0.155672
R1007 VTAIL.n519 VTAIL.n518 0.155672
R1008 VTAIL.n518 VTAIL.n494 0.155672
R1009 VTAIL.n511 VTAIL.n494 0.155672
R1010 VTAIL.n511 VTAIL.n510 0.155672
R1011 VTAIL.n510 VTAIL.n498 0.155672
R1012 VTAIL.n503 VTAIL.n498 0.155672
R1013 VTAIL.n471 VTAIL.n397 0.155672
R1014 VTAIL.n463 VTAIL.n397 0.155672
R1015 VTAIL.n463 VTAIL.n462 0.155672
R1016 VTAIL.n462 VTAIL.n402 0.155672
R1017 VTAIL.n455 VTAIL.n402 0.155672
R1018 VTAIL.n455 VTAIL.n454 0.155672
R1019 VTAIL.n454 VTAIL.n406 0.155672
R1020 VTAIL.n447 VTAIL.n406 0.155672
R1021 VTAIL.n447 VTAIL.n446 0.155672
R1022 VTAIL.n446 VTAIL.n410 0.155672
R1023 VTAIL.n439 VTAIL.n410 0.155672
R1024 VTAIL.n439 VTAIL.n438 0.155672
R1025 VTAIL.n438 VTAIL.n414 0.155672
R1026 VTAIL.n431 VTAIL.n414 0.155672
R1027 VTAIL.n431 VTAIL.n430 0.155672
R1028 VTAIL.n430 VTAIL.n418 0.155672
R1029 VTAIL.n423 VTAIL.n418 0.155672
R1030 VTAIL.n393 VTAIL.n319 0.155672
R1031 VTAIL.n385 VTAIL.n319 0.155672
R1032 VTAIL.n385 VTAIL.n384 0.155672
R1033 VTAIL.n384 VTAIL.n324 0.155672
R1034 VTAIL.n377 VTAIL.n324 0.155672
R1035 VTAIL.n377 VTAIL.n376 0.155672
R1036 VTAIL.n376 VTAIL.n328 0.155672
R1037 VTAIL.n369 VTAIL.n328 0.155672
R1038 VTAIL.n369 VTAIL.n368 0.155672
R1039 VTAIL.n368 VTAIL.n332 0.155672
R1040 VTAIL.n361 VTAIL.n332 0.155672
R1041 VTAIL.n361 VTAIL.n360 0.155672
R1042 VTAIL.n360 VTAIL.n336 0.155672
R1043 VTAIL.n353 VTAIL.n336 0.155672
R1044 VTAIL.n353 VTAIL.n352 0.155672
R1045 VTAIL.n352 VTAIL.n340 0.155672
R1046 VTAIL.n345 VTAIL.n340 0.155672
R1047 VTAIL.n313 VTAIL.n239 0.155672
R1048 VTAIL.n305 VTAIL.n239 0.155672
R1049 VTAIL.n305 VTAIL.n304 0.155672
R1050 VTAIL.n304 VTAIL.n244 0.155672
R1051 VTAIL.n297 VTAIL.n244 0.155672
R1052 VTAIL.n297 VTAIL.n296 0.155672
R1053 VTAIL.n296 VTAIL.n248 0.155672
R1054 VTAIL.n289 VTAIL.n248 0.155672
R1055 VTAIL.n289 VTAIL.n288 0.155672
R1056 VTAIL.n288 VTAIL.n252 0.155672
R1057 VTAIL.n281 VTAIL.n252 0.155672
R1058 VTAIL.n281 VTAIL.n280 0.155672
R1059 VTAIL.n280 VTAIL.n256 0.155672
R1060 VTAIL.n273 VTAIL.n256 0.155672
R1061 VTAIL.n273 VTAIL.n272 0.155672
R1062 VTAIL.n272 VTAIL.n260 0.155672
R1063 VTAIL.n265 VTAIL.n260 0.155672
R1064 VTAIL VTAIL.n1 0.0586897
R1065 VN.n5 VN.t0 199.073
R1066 VN.n28 VN.t3 199.073
R1067 VN.n6 VN.t7 166.101
R1068 VN.n13 VN.t6 166.101
R1069 VN.n21 VN.t5 166.101
R1070 VN.n29 VN.t4 166.101
R1071 VN.n36 VN.t2 166.101
R1072 VN.n44 VN.t1 166.101
R1073 VN.n43 VN.n23 161.3
R1074 VN.n42 VN.n41 161.3
R1075 VN.n40 VN.n24 161.3
R1076 VN.n39 VN.n38 161.3
R1077 VN.n37 VN.n25 161.3
R1078 VN.n35 VN.n34 161.3
R1079 VN.n33 VN.n26 161.3
R1080 VN.n32 VN.n31 161.3
R1081 VN.n30 VN.n27 161.3
R1082 VN.n20 VN.n0 161.3
R1083 VN.n19 VN.n18 161.3
R1084 VN.n17 VN.n1 161.3
R1085 VN.n16 VN.n15 161.3
R1086 VN.n14 VN.n2 161.3
R1087 VN.n12 VN.n11 161.3
R1088 VN.n10 VN.n3 161.3
R1089 VN.n9 VN.n8 161.3
R1090 VN.n7 VN.n4 161.3
R1091 VN.n22 VN.n21 95.7567
R1092 VN.n45 VN.n44 95.7567
R1093 VN.n8 VN.n3 56.4773
R1094 VN.n31 VN.n26 56.4773
R1095 VN.n19 VN.n1 52.0954
R1096 VN.n42 VN.n24 52.0954
R1097 VN VN.n45 50.0739
R1098 VN.n6 VN.n5 49.1578
R1099 VN.n29 VN.n28 49.1578
R1100 VN.n15 VN.n1 28.7258
R1101 VN.n38 VN.n24 28.7258
R1102 VN.n8 VN.n7 24.3439
R1103 VN.n12 VN.n3 24.3439
R1104 VN.n15 VN.n14 24.3439
R1105 VN.n20 VN.n19 24.3439
R1106 VN.n31 VN.n30 24.3439
R1107 VN.n38 VN.n37 24.3439
R1108 VN.n35 VN.n26 24.3439
R1109 VN.n43 VN.n42 24.3439
R1110 VN.n7 VN.n6 21.1793
R1111 VN.n13 VN.n12 21.1793
R1112 VN.n30 VN.n29 21.1793
R1113 VN.n36 VN.n35 21.1793
R1114 VN.n21 VN.n20 14.85
R1115 VN.n44 VN.n43 14.85
R1116 VN.n28 VN.n27 9.46412
R1117 VN.n5 VN.n4 9.46412
R1118 VN.n14 VN.n13 3.16515
R1119 VN.n37 VN.n36 3.16515
R1120 VN.n45 VN.n23 0.278398
R1121 VN.n22 VN.n0 0.278398
R1122 VN.n41 VN.n23 0.189894
R1123 VN.n41 VN.n40 0.189894
R1124 VN.n40 VN.n39 0.189894
R1125 VN.n39 VN.n25 0.189894
R1126 VN.n34 VN.n25 0.189894
R1127 VN.n34 VN.n33 0.189894
R1128 VN.n33 VN.n32 0.189894
R1129 VN.n32 VN.n27 0.189894
R1130 VN.n9 VN.n4 0.189894
R1131 VN.n10 VN.n9 0.189894
R1132 VN.n11 VN.n10 0.189894
R1133 VN.n11 VN.n2 0.189894
R1134 VN.n16 VN.n2 0.189894
R1135 VN.n17 VN.n16 0.189894
R1136 VN.n18 VN.n17 0.189894
R1137 VN.n18 VN.n0 0.189894
R1138 VN VN.n22 0.153422
R1139 VDD2.n2 VDD2.n1 75.0155
R1140 VDD2.n2 VDD2.n0 75.0155
R1141 VDD2 VDD2.n5 75.0126
R1142 VDD2.n4 VDD2.n3 74.0495
R1143 VDD2.n4 VDD2.n2 45.03
R1144 VDD2.n5 VDD2.t3 2.31238
R1145 VDD2.n5 VDD2.t4 2.31238
R1146 VDD2.n3 VDD2.t6 2.31238
R1147 VDD2.n3 VDD2.t5 2.31238
R1148 VDD2.n1 VDD2.t1 2.31238
R1149 VDD2.n1 VDD2.t2 2.31238
R1150 VDD2.n0 VDD2.t7 2.31238
R1151 VDD2.n0 VDD2.t0 2.31238
R1152 VDD2 VDD2.n4 1.08024
R1153 B.n555 B.n80 585
R1154 B.n557 B.n556 585
R1155 B.n558 B.n79 585
R1156 B.n560 B.n559 585
R1157 B.n561 B.n78 585
R1158 B.n563 B.n562 585
R1159 B.n564 B.n77 585
R1160 B.n566 B.n565 585
R1161 B.n567 B.n76 585
R1162 B.n569 B.n568 585
R1163 B.n570 B.n75 585
R1164 B.n572 B.n571 585
R1165 B.n573 B.n74 585
R1166 B.n575 B.n574 585
R1167 B.n576 B.n73 585
R1168 B.n578 B.n577 585
R1169 B.n579 B.n72 585
R1170 B.n581 B.n580 585
R1171 B.n582 B.n71 585
R1172 B.n584 B.n583 585
R1173 B.n585 B.n70 585
R1174 B.n587 B.n586 585
R1175 B.n588 B.n69 585
R1176 B.n590 B.n589 585
R1177 B.n591 B.n68 585
R1178 B.n593 B.n592 585
R1179 B.n594 B.n67 585
R1180 B.n596 B.n595 585
R1181 B.n597 B.n66 585
R1182 B.n599 B.n598 585
R1183 B.n600 B.n65 585
R1184 B.n602 B.n601 585
R1185 B.n603 B.n64 585
R1186 B.n605 B.n604 585
R1187 B.n606 B.n63 585
R1188 B.n608 B.n607 585
R1189 B.n609 B.n62 585
R1190 B.n611 B.n610 585
R1191 B.n612 B.n61 585
R1192 B.n614 B.n613 585
R1193 B.n615 B.n60 585
R1194 B.n617 B.n616 585
R1195 B.n618 B.n59 585
R1196 B.n620 B.n619 585
R1197 B.n621 B.n58 585
R1198 B.n623 B.n622 585
R1199 B.n624 B.n57 585
R1200 B.n626 B.n625 585
R1201 B.n628 B.n627 585
R1202 B.n629 B.n53 585
R1203 B.n631 B.n630 585
R1204 B.n632 B.n52 585
R1205 B.n634 B.n633 585
R1206 B.n635 B.n51 585
R1207 B.n637 B.n636 585
R1208 B.n638 B.n50 585
R1209 B.n640 B.n639 585
R1210 B.n642 B.n47 585
R1211 B.n644 B.n643 585
R1212 B.n645 B.n46 585
R1213 B.n647 B.n646 585
R1214 B.n648 B.n45 585
R1215 B.n650 B.n649 585
R1216 B.n651 B.n44 585
R1217 B.n653 B.n652 585
R1218 B.n654 B.n43 585
R1219 B.n656 B.n655 585
R1220 B.n657 B.n42 585
R1221 B.n659 B.n658 585
R1222 B.n660 B.n41 585
R1223 B.n662 B.n661 585
R1224 B.n663 B.n40 585
R1225 B.n665 B.n664 585
R1226 B.n666 B.n39 585
R1227 B.n668 B.n667 585
R1228 B.n669 B.n38 585
R1229 B.n671 B.n670 585
R1230 B.n672 B.n37 585
R1231 B.n674 B.n673 585
R1232 B.n675 B.n36 585
R1233 B.n677 B.n676 585
R1234 B.n678 B.n35 585
R1235 B.n680 B.n679 585
R1236 B.n681 B.n34 585
R1237 B.n683 B.n682 585
R1238 B.n684 B.n33 585
R1239 B.n686 B.n685 585
R1240 B.n687 B.n32 585
R1241 B.n689 B.n688 585
R1242 B.n690 B.n31 585
R1243 B.n692 B.n691 585
R1244 B.n693 B.n30 585
R1245 B.n695 B.n694 585
R1246 B.n696 B.n29 585
R1247 B.n698 B.n697 585
R1248 B.n699 B.n28 585
R1249 B.n701 B.n700 585
R1250 B.n702 B.n27 585
R1251 B.n704 B.n703 585
R1252 B.n705 B.n26 585
R1253 B.n707 B.n706 585
R1254 B.n708 B.n25 585
R1255 B.n710 B.n709 585
R1256 B.n711 B.n24 585
R1257 B.n713 B.n712 585
R1258 B.n554 B.n553 585
R1259 B.n552 B.n81 585
R1260 B.n551 B.n550 585
R1261 B.n549 B.n82 585
R1262 B.n548 B.n547 585
R1263 B.n546 B.n83 585
R1264 B.n545 B.n544 585
R1265 B.n543 B.n84 585
R1266 B.n542 B.n541 585
R1267 B.n540 B.n85 585
R1268 B.n539 B.n538 585
R1269 B.n537 B.n86 585
R1270 B.n536 B.n535 585
R1271 B.n534 B.n87 585
R1272 B.n533 B.n532 585
R1273 B.n531 B.n88 585
R1274 B.n530 B.n529 585
R1275 B.n528 B.n89 585
R1276 B.n527 B.n526 585
R1277 B.n525 B.n90 585
R1278 B.n524 B.n523 585
R1279 B.n522 B.n91 585
R1280 B.n521 B.n520 585
R1281 B.n519 B.n92 585
R1282 B.n518 B.n517 585
R1283 B.n516 B.n93 585
R1284 B.n515 B.n514 585
R1285 B.n513 B.n94 585
R1286 B.n512 B.n511 585
R1287 B.n510 B.n95 585
R1288 B.n509 B.n508 585
R1289 B.n507 B.n96 585
R1290 B.n506 B.n505 585
R1291 B.n504 B.n97 585
R1292 B.n503 B.n502 585
R1293 B.n501 B.n98 585
R1294 B.n500 B.n499 585
R1295 B.n498 B.n99 585
R1296 B.n497 B.n496 585
R1297 B.n495 B.n100 585
R1298 B.n494 B.n493 585
R1299 B.n492 B.n101 585
R1300 B.n491 B.n490 585
R1301 B.n489 B.n102 585
R1302 B.n488 B.n487 585
R1303 B.n486 B.n103 585
R1304 B.n485 B.n484 585
R1305 B.n483 B.n104 585
R1306 B.n482 B.n481 585
R1307 B.n480 B.n105 585
R1308 B.n479 B.n478 585
R1309 B.n477 B.n106 585
R1310 B.n476 B.n475 585
R1311 B.n474 B.n107 585
R1312 B.n473 B.n472 585
R1313 B.n471 B.n108 585
R1314 B.n470 B.n469 585
R1315 B.n468 B.n109 585
R1316 B.n467 B.n466 585
R1317 B.n465 B.n110 585
R1318 B.n464 B.n463 585
R1319 B.n462 B.n111 585
R1320 B.n461 B.n460 585
R1321 B.n459 B.n112 585
R1322 B.n458 B.n457 585
R1323 B.n456 B.n113 585
R1324 B.n455 B.n454 585
R1325 B.n453 B.n114 585
R1326 B.n452 B.n451 585
R1327 B.n450 B.n115 585
R1328 B.n449 B.n448 585
R1329 B.n447 B.n116 585
R1330 B.n446 B.n445 585
R1331 B.n444 B.n117 585
R1332 B.n443 B.n442 585
R1333 B.n441 B.n118 585
R1334 B.n440 B.n439 585
R1335 B.n438 B.n119 585
R1336 B.n437 B.n436 585
R1337 B.n435 B.n120 585
R1338 B.n434 B.n433 585
R1339 B.n432 B.n121 585
R1340 B.n431 B.n430 585
R1341 B.n429 B.n122 585
R1342 B.n428 B.n427 585
R1343 B.n426 B.n123 585
R1344 B.n425 B.n424 585
R1345 B.n266 B.n265 585
R1346 B.n267 B.n180 585
R1347 B.n269 B.n268 585
R1348 B.n270 B.n179 585
R1349 B.n272 B.n271 585
R1350 B.n273 B.n178 585
R1351 B.n275 B.n274 585
R1352 B.n276 B.n177 585
R1353 B.n278 B.n277 585
R1354 B.n279 B.n176 585
R1355 B.n281 B.n280 585
R1356 B.n282 B.n175 585
R1357 B.n284 B.n283 585
R1358 B.n285 B.n174 585
R1359 B.n287 B.n286 585
R1360 B.n288 B.n173 585
R1361 B.n290 B.n289 585
R1362 B.n291 B.n172 585
R1363 B.n293 B.n292 585
R1364 B.n294 B.n171 585
R1365 B.n296 B.n295 585
R1366 B.n297 B.n170 585
R1367 B.n299 B.n298 585
R1368 B.n300 B.n169 585
R1369 B.n302 B.n301 585
R1370 B.n303 B.n168 585
R1371 B.n305 B.n304 585
R1372 B.n306 B.n167 585
R1373 B.n308 B.n307 585
R1374 B.n309 B.n166 585
R1375 B.n311 B.n310 585
R1376 B.n312 B.n165 585
R1377 B.n314 B.n313 585
R1378 B.n315 B.n164 585
R1379 B.n317 B.n316 585
R1380 B.n318 B.n163 585
R1381 B.n320 B.n319 585
R1382 B.n321 B.n162 585
R1383 B.n323 B.n322 585
R1384 B.n324 B.n161 585
R1385 B.n326 B.n325 585
R1386 B.n327 B.n160 585
R1387 B.n329 B.n328 585
R1388 B.n330 B.n159 585
R1389 B.n332 B.n331 585
R1390 B.n333 B.n158 585
R1391 B.n335 B.n334 585
R1392 B.n336 B.n155 585
R1393 B.n339 B.n338 585
R1394 B.n340 B.n154 585
R1395 B.n342 B.n341 585
R1396 B.n343 B.n153 585
R1397 B.n345 B.n344 585
R1398 B.n346 B.n152 585
R1399 B.n348 B.n347 585
R1400 B.n349 B.n151 585
R1401 B.n351 B.n350 585
R1402 B.n353 B.n352 585
R1403 B.n354 B.n147 585
R1404 B.n356 B.n355 585
R1405 B.n357 B.n146 585
R1406 B.n359 B.n358 585
R1407 B.n360 B.n145 585
R1408 B.n362 B.n361 585
R1409 B.n363 B.n144 585
R1410 B.n365 B.n364 585
R1411 B.n366 B.n143 585
R1412 B.n368 B.n367 585
R1413 B.n369 B.n142 585
R1414 B.n371 B.n370 585
R1415 B.n372 B.n141 585
R1416 B.n374 B.n373 585
R1417 B.n375 B.n140 585
R1418 B.n377 B.n376 585
R1419 B.n378 B.n139 585
R1420 B.n380 B.n379 585
R1421 B.n381 B.n138 585
R1422 B.n383 B.n382 585
R1423 B.n384 B.n137 585
R1424 B.n386 B.n385 585
R1425 B.n387 B.n136 585
R1426 B.n389 B.n388 585
R1427 B.n390 B.n135 585
R1428 B.n392 B.n391 585
R1429 B.n393 B.n134 585
R1430 B.n395 B.n394 585
R1431 B.n396 B.n133 585
R1432 B.n398 B.n397 585
R1433 B.n399 B.n132 585
R1434 B.n401 B.n400 585
R1435 B.n402 B.n131 585
R1436 B.n404 B.n403 585
R1437 B.n405 B.n130 585
R1438 B.n407 B.n406 585
R1439 B.n408 B.n129 585
R1440 B.n410 B.n409 585
R1441 B.n411 B.n128 585
R1442 B.n413 B.n412 585
R1443 B.n414 B.n127 585
R1444 B.n416 B.n415 585
R1445 B.n417 B.n126 585
R1446 B.n419 B.n418 585
R1447 B.n420 B.n125 585
R1448 B.n422 B.n421 585
R1449 B.n423 B.n124 585
R1450 B.n264 B.n181 585
R1451 B.n263 B.n262 585
R1452 B.n261 B.n182 585
R1453 B.n260 B.n259 585
R1454 B.n258 B.n183 585
R1455 B.n257 B.n256 585
R1456 B.n255 B.n184 585
R1457 B.n254 B.n253 585
R1458 B.n252 B.n185 585
R1459 B.n251 B.n250 585
R1460 B.n249 B.n186 585
R1461 B.n248 B.n247 585
R1462 B.n246 B.n187 585
R1463 B.n245 B.n244 585
R1464 B.n243 B.n188 585
R1465 B.n242 B.n241 585
R1466 B.n240 B.n189 585
R1467 B.n239 B.n238 585
R1468 B.n237 B.n190 585
R1469 B.n236 B.n235 585
R1470 B.n234 B.n191 585
R1471 B.n233 B.n232 585
R1472 B.n231 B.n192 585
R1473 B.n230 B.n229 585
R1474 B.n228 B.n193 585
R1475 B.n227 B.n226 585
R1476 B.n225 B.n194 585
R1477 B.n224 B.n223 585
R1478 B.n222 B.n195 585
R1479 B.n221 B.n220 585
R1480 B.n219 B.n196 585
R1481 B.n218 B.n217 585
R1482 B.n216 B.n197 585
R1483 B.n215 B.n214 585
R1484 B.n213 B.n198 585
R1485 B.n212 B.n211 585
R1486 B.n210 B.n199 585
R1487 B.n209 B.n208 585
R1488 B.n207 B.n200 585
R1489 B.n206 B.n205 585
R1490 B.n204 B.n201 585
R1491 B.n203 B.n202 585
R1492 B.n2 B.n0 585
R1493 B.n777 B.n1 585
R1494 B.n776 B.n775 585
R1495 B.n774 B.n3 585
R1496 B.n773 B.n772 585
R1497 B.n771 B.n4 585
R1498 B.n770 B.n769 585
R1499 B.n768 B.n5 585
R1500 B.n767 B.n766 585
R1501 B.n765 B.n6 585
R1502 B.n764 B.n763 585
R1503 B.n762 B.n7 585
R1504 B.n761 B.n760 585
R1505 B.n759 B.n8 585
R1506 B.n758 B.n757 585
R1507 B.n756 B.n9 585
R1508 B.n755 B.n754 585
R1509 B.n753 B.n10 585
R1510 B.n752 B.n751 585
R1511 B.n750 B.n11 585
R1512 B.n749 B.n748 585
R1513 B.n747 B.n12 585
R1514 B.n746 B.n745 585
R1515 B.n744 B.n13 585
R1516 B.n743 B.n742 585
R1517 B.n741 B.n14 585
R1518 B.n740 B.n739 585
R1519 B.n738 B.n15 585
R1520 B.n737 B.n736 585
R1521 B.n735 B.n16 585
R1522 B.n734 B.n733 585
R1523 B.n732 B.n17 585
R1524 B.n731 B.n730 585
R1525 B.n729 B.n18 585
R1526 B.n728 B.n727 585
R1527 B.n726 B.n19 585
R1528 B.n725 B.n724 585
R1529 B.n723 B.n20 585
R1530 B.n722 B.n721 585
R1531 B.n720 B.n21 585
R1532 B.n719 B.n718 585
R1533 B.n717 B.n22 585
R1534 B.n716 B.n715 585
R1535 B.n714 B.n23 585
R1536 B.n779 B.n778 585
R1537 B.n266 B.n181 487.695
R1538 B.n712 B.n23 487.695
R1539 B.n424 B.n423 487.695
R1540 B.n555 B.n554 487.695
R1541 B.n148 B.t2 458.623
R1542 B.n54 B.t7 458.623
R1543 B.n156 B.t5 458.623
R1544 B.n48 B.t10 458.623
R1545 B.n149 B.t1 412.661
R1546 B.n55 B.t8 412.661
R1547 B.n157 B.t4 412.659
R1548 B.n49 B.t11 412.659
R1549 B.n148 B.t0 373.111
R1550 B.n156 B.t3 373.111
R1551 B.n48 B.t9 373.111
R1552 B.n54 B.t6 373.111
R1553 B.n262 B.n181 163.367
R1554 B.n262 B.n261 163.367
R1555 B.n261 B.n260 163.367
R1556 B.n260 B.n183 163.367
R1557 B.n256 B.n183 163.367
R1558 B.n256 B.n255 163.367
R1559 B.n255 B.n254 163.367
R1560 B.n254 B.n185 163.367
R1561 B.n250 B.n185 163.367
R1562 B.n250 B.n249 163.367
R1563 B.n249 B.n248 163.367
R1564 B.n248 B.n187 163.367
R1565 B.n244 B.n187 163.367
R1566 B.n244 B.n243 163.367
R1567 B.n243 B.n242 163.367
R1568 B.n242 B.n189 163.367
R1569 B.n238 B.n189 163.367
R1570 B.n238 B.n237 163.367
R1571 B.n237 B.n236 163.367
R1572 B.n236 B.n191 163.367
R1573 B.n232 B.n191 163.367
R1574 B.n232 B.n231 163.367
R1575 B.n231 B.n230 163.367
R1576 B.n230 B.n193 163.367
R1577 B.n226 B.n193 163.367
R1578 B.n226 B.n225 163.367
R1579 B.n225 B.n224 163.367
R1580 B.n224 B.n195 163.367
R1581 B.n220 B.n195 163.367
R1582 B.n220 B.n219 163.367
R1583 B.n219 B.n218 163.367
R1584 B.n218 B.n197 163.367
R1585 B.n214 B.n197 163.367
R1586 B.n214 B.n213 163.367
R1587 B.n213 B.n212 163.367
R1588 B.n212 B.n199 163.367
R1589 B.n208 B.n199 163.367
R1590 B.n208 B.n207 163.367
R1591 B.n207 B.n206 163.367
R1592 B.n206 B.n201 163.367
R1593 B.n202 B.n201 163.367
R1594 B.n202 B.n2 163.367
R1595 B.n778 B.n2 163.367
R1596 B.n778 B.n777 163.367
R1597 B.n777 B.n776 163.367
R1598 B.n776 B.n3 163.367
R1599 B.n772 B.n3 163.367
R1600 B.n772 B.n771 163.367
R1601 B.n771 B.n770 163.367
R1602 B.n770 B.n5 163.367
R1603 B.n766 B.n5 163.367
R1604 B.n766 B.n765 163.367
R1605 B.n765 B.n764 163.367
R1606 B.n764 B.n7 163.367
R1607 B.n760 B.n7 163.367
R1608 B.n760 B.n759 163.367
R1609 B.n759 B.n758 163.367
R1610 B.n758 B.n9 163.367
R1611 B.n754 B.n9 163.367
R1612 B.n754 B.n753 163.367
R1613 B.n753 B.n752 163.367
R1614 B.n752 B.n11 163.367
R1615 B.n748 B.n11 163.367
R1616 B.n748 B.n747 163.367
R1617 B.n747 B.n746 163.367
R1618 B.n746 B.n13 163.367
R1619 B.n742 B.n13 163.367
R1620 B.n742 B.n741 163.367
R1621 B.n741 B.n740 163.367
R1622 B.n740 B.n15 163.367
R1623 B.n736 B.n15 163.367
R1624 B.n736 B.n735 163.367
R1625 B.n735 B.n734 163.367
R1626 B.n734 B.n17 163.367
R1627 B.n730 B.n17 163.367
R1628 B.n730 B.n729 163.367
R1629 B.n729 B.n728 163.367
R1630 B.n728 B.n19 163.367
R1631 B.n724 B.n19 163.367
R1632 B.n724 B.n723 163.367
R1633 B.n723 B.n722 163.367
R1634 B.n722 B.n21 163.367
R1635 B.n718 B.n21 163.367
R1636 B.n718 B.n717 163.367
R1637 B.n717 B.n716 163.367
R1638 B.n716 B.n23 163.367
R1639 B.n267 B.n266 163.367
R1640 B.n268 B.n267 163.367
R1641 B.n268 B.n179 163.367
R1642 B.n272 B.n179 163.367
R1643 B.n273 B.n272 163.367
R1644 B.n274 B.n273 163.367
R1645 B.n274 B.n177 163.367
R1646 B.n278 B.n177 163.367
R1647 B.n279 B.n278 163.367
R1648 B.n280 B.n279 163.367
R1649 B.n280 B.n175 163.367
R1650 B.n284 B.n175 163.367
R1651 B.n285 B.n284 163.367
R1652 B.n286 B.n285 163.367
R1653 B.n286 B.n173 163.367
R1654 B.n290 B.n173 163.367
R1655 B.n291 B.n290 163.367
R1656 B.n292 B.n291 163.367
R1657 B.n292 B.n171 163.367
R1658 B.n296 B.n171 163.367
R1659 B.n297 B.n296 163.367
R1660 B.n298 B.n297 163.367
R1661 B.n298 B.n169 163.367
R1662 B.n302 B.n169 163.367
R1663 B.n303 B.n302 163.367
R1664 B.n304 B.n303 163.367
R1665 B.n304 B.n167 163.367
R1666 B.n308 B.n167 163.367
R1667 B.n309 B.n308 163.367
R1668 B.n310 B.n309 163.367
R1669 B.n310 B.n165 163.367
R1670 B.n314 B.n165 163.367
R1671 B.n315 B.n314 163.367
R1672 B.n316 B.n315 163.367
R1673 B.n316 B.n163 163.367
R1674 B.n320 B.n163 163.367
R1675 B.n321 B.n320 163.367
R1676 B.n322 B.n321 163.367
R1677 B.n322 B.n161 163.367
R1678 B.n326 B.n161 163.367
R1679 B.n327 B.n326 163.367
R1680 B.n328 B.n327 163.367
R1681 B.n328 B.n159 163.367
R1682 B.n332 B.n159 163.367
R1683 B.n333 B.n332 163.367
R1684 B.n334 B.n333 163.367
R1685 B.n334 B.n155 163.367
R1686 B.n339 B.n155 163.367
R1687 B.n340 B.n339 163.367
R1688 B.n341 B.n340 163.367
R1689 B.n341 B.n153 163.367
R1690 B.n345 B.n153 163.367
R1691 B.n346 B.n345 163.367
R1692 B.n347 B.n346 163.367
R1693 B.n347 B.n151 163.367
R1694 B.n351 B.n151 163.367
R1695 B.n352 B.n351 163.367
R1696 B.n352 B.n147 163.367
R1697 B.n356 B.n147 163.367
R1698 B.n357 B.n356 163.367
R1699 B.n358 B.n357 163.367
R1700 B.n358 B.n145 163.367
R1701 B.n362 B.n145 163.367
R1702 B.n363 B.n362 163.367
R1703 B.n364 B.n363 163.367
R1704 B.n364 B.n143 163.367
R1705 B.n368 B.n143 163.367
R1706 B.n369 B.n368 163.367
R1707 B.n370 B.n369 163.367
R1708 B.n370 B.n141 163.367
R1709 B.n374 B.n141 163.367
R1710 B.n375 B.n374 163.367
R1711 B.n376 B.n375 163.367
R1712 B.n376 B.n139 163.367
R1713 B.n380 B.n139 163.367
R1714 B.n381 B.n380 163.367
R1715 B.n382 B.n381 163.367
R1716 B.n382 B.n137 163.367
R1717 B.n386 B.n137 163.367
R1718 B.n387 B.n386 163.367
R1719 B.n388 B.n387 163.367
R1720 B.n388 B.n135 163.367
R1721 B.n392 B.n135 163.367
R1722 B.n393 B.n392 163.367
R1723 B.n394 B.n393 163.367
R1724 B.n394 B.n133 163.367
R1725 B.n398 B.n133 163.367
R1726 B.n399 B.n398 163.367
R1727 B.n400 B.n399 163.367
R1728 B.n400 B.n131 163.367
R1729 B.n404 B.n131 163.367
R1730 B.n405 B.n404 163.367
R1731 B.n406 B.n405 163.367
R1732 B.n406 B.n129 163.367
R1733 B.n410 B.n129 163.367
R1734 B.n411 B.n410 163.367
R1735 B.n412 B.n411 163.367
R1736 B.n412 B.n127 163.367
R1737 B.n416 B.n127 163.367
R1738 B.n417 B.n416 163.367
R1739 B.n418 B.n417 163.367
R1740 B.n418 B.n125 163.367
R1741 B.n422 B.n125 163.367
R1742 B.n423 B.n422 163.367
R1743 B.n424 B.n123 163.367
R1744 B.n428 B.n123 163.367
R1745 B.n429 B.n428 163.367
R1746 B.n430 B.n429 163.367
R1747 B.n430 B.n121 163.367
R1748 B.n434 B.n121 163.367
R1749 B.n435 B.n434 163.367
R1750 B.n436 B.n435 163.367
R1751 B.n436 B.n119 163.367
R1752 B.n440 B.n119 163.367
R1753 B.n441 B.n440 163.367
R1754 B.n442 B.n441 163.367
R1755 B.n442 B.n117 163.367
R1756 B.n446 B.n117 163.367
R1757 B.n447 B.n446 163.367
R1758 B.n448 B.n447 163.367
R1759 B.n448 B.n115 163.367
R1760 B.n452 B.n115 163.367
R1761 B.n453 B.n452 163.367
R1762 B.n454 B.n453 163.367
R1763 B.n454 B.n113 163.367
R1764 B.n458 B.n113 163.367
R1765 B.n459 B.n458 163.367
R1766 B.n460 B.n459 163.367
R1767 B.n460 B.n111 163.367
R1768 B.n464 B.n111 163.367
R1769 B.n465 B.n464 163.367
R1770 B.n466 B.n465 163.367
R1771 B.n466 B.n109 163.367
R1772 B.n470 B.n109 163.367
R1773 B.n471 B.n470 163.367
R1774 B.n472 B.n471 163.367
R1775 B.n472 B.n107 163.367
R1776 B.n476 B.n107 163.367
R1777 B.n477 B.n476 163.367
R1778 B.n478 B.n477 163.367
R1779 B.n478 B.n105 163.367
R1780 B.n482 B.n105 163.367
R1781 B.n483 B.n482 163.367
R1782 B.n484 B.n483 163.367
R1783 B.n484 B.n103 163.367
R1784 B.n488 B.n103 163.367
R1785 B.n489 B.n488 163.367
R1786 B.n490 B.n489 163.367
R1787 B.n490 B.n101 163.367
R1788 B.n494 B.n101 163.367
R1789 B.n495 B.n494 163.367
R1790 B.n496 B.n495 163.367
R1791 B.n496 B.n99 163.367
R1792 B.n500 B.n99 163.367
R1793 B.n501 B.n500 163.367
R1794 B.n502 B.n501 163.367
R1795 B.n502 B.n97 163.367
R1796 B.n506 B.n97 163.367
R1797 B.n507 B.n506 163.367
R1798 B.n508 B.n507 163.367
R1799 B.n508 B.n95 163.367
R1800 B.n512 B.n95 163.367
R1801 B.n513 B.n512 163.367
R1802 B.n514 B.n513 163.367
R1803 B.n514 B.n93 163.367
R1804 B.n518 B.n93 163.367
R1805 B.n519 B.n518 163.367
R1806 B.n520 B.n519 163.367
R1807 B.n520 B.n91 163.367
R1808 B.n524 B.n91 163.367
R1809 B.n525 B.n524 163.367
R1810 B.n526 B.n525 163.367
R1811 B.n526 B.n89 163.367
R1812 B.n530 B.n89 163.367
R1813 B.n531 B.n530 163.367
R1814 B.n532 B.n531 163.367
R1815 B.n532 B.n87 163.367
R1816 B.n536 B.n87 163.367
R1817 B.n537 B.n536 163.367
R1818 B.n538 B.n537 163.367
R1819 B.n538 B.n85 163.367
R1820 B.n542 B.n85 163.367
R1821 B.n543 B.n542 163.367
R1822 B.n544 B.n543 163.367
R1823 B.n544 B.n83 163.367
R1824 B.n548 B.n83 163.367
R1825 B.n549 B.n548 163.367
R1826 B.n550 B.n549 163.367
R1827 B.n550 B.n81 163.367
R1828 B.n554 B.n81 163.367
R1829 B.n712 B.n711 163.367
R1830 B.n711 B.n710 163.367
R1831 B.n710 B.n25 163.367
R1832 B.n706 B.n25 163.367
R1833 B.n706 B.n705 163.367
R1834 B.n705 B.n704 163.367
R1835 B.n704 B.n27 163.367
R1836 B.n700 B.n27 163.367
R1837 B.n700 B.n699 163.367
R1838 B.n699 B.n698 163.367
R1839 B.n698 B.n29 163.367
R1840 B.n694 B.n29 163.367
R1841 B.n694 B.n693 163.367
R1842 B.n693 B.n692 163.367
R1843 B.n692 B.n31 163.367
R1844 B.n688 B.n31 163.367
R1845 B.n688 B.n687 163.367
R1846 B.n687 B.n686 163.367
R1847 B.n686 B.n33 163.367
R1848 B.n682 B.n33 163.367
R1849 B.n682 B.n681 163.367
R1850 B.n681 B.n680 163.367
R1851 B.n680 B.n35 163.367
R1852 B.n676 B.n35 163.367
R1853 B.n676 B.n675 163.367
R1854 B.n675 B.n674 163.367
R1855 B.n674 B.n37 163.367
R1856 B.n670 B.n37 163.367
R1857 B.n670 B.n669 163.367
R1858 B.n669 B.n668 163.367
R1859 B.n668 B.n39 163.367
R1860 B.n664 B.n39 163.367
R1861 B.n664 B.n663 163.367
R1862 B.n663 B.n662 163.367
R1863 B.n662 B.n41 163.367
R1864 B.n658 B.n41 163.367
R1865 B.n658 B.n657 163.367
R1866 B.n657 B.n656 163.367
R1867 B.n656 B.n43 163.367
R1868 B.n652 B.n43 163.367
R1869 B.n652 B.n651 163.367
R1870 B.n651 B.n650 163.367
R1871 B.n650 B.n45 163.367
R1872 B.n646 B.n45 163.367
R1873 B.n646 B.n645 163.367
R1874 B.n645 B.n644 163.367
R1875 B.n644 B.n47 163.367
R1876 B.n639 B.n47 163.367
R1877 B.n639 B.n638 163.367
R1878 B.n638 B.n637 163.367
R1879 B.n637 B.n51 163.367
R1880 B.n633 B.n51 163.367
R1881 B.n633 B.n632 163.367
R1882 B.n632 B.n631 163.367
R1883 B.n631 B.n53 163.367
R1884 B.n627 B.n53 163.367
R1885 B.n627 B.n626 163.367
R1886 B.n626 B.n57 163.367
R1887 B.n622 B.n57 163.367
R1888 B.n622 B.n621 163.367
R1889 B.n621 B.n620 163.367
R1890 B.n620 B.n59 163.367
R1891 B.n616 B.n59 163.367
R1892 B.n616 B.n615 163.367
R1893 B.n615 B.n614 163.367
R1894 B.n614 B.n61 163.367
R1895 B.n610 B.n61 163.367
R1896 B.n610 B.n609 163.367
R1897 B.n609 B.n608 163.367
R1898 B.n608 B.n63 163.367
R1899 B.n604 B.n63 163.367
R1900 B.n604 B.n603 163.367
R1901 B.n603 B.n602 163.367
R1902 B.n602 B.n65 163.367
R1903 B.n598 B.n65 163.367
R1904 B.n598 B.n597 163.367
R1905 B.n597 B.n596 163.367
R1906 B.n596 B.n67 163.367
R1907 B.n592 B.n67 163.367
R1908 B.n592 B.n591 163.367
R1909 B.n591 B.n590 163.367
R1910 B.n590 B.n69 163.367
R1911 B.n586 B.n69 163.367
R1912 B.n586 B.n585 163.367
R1913 B.n585 B.n584 163.367
R1914 B.n584 B.n71 163.367
R1915 B.n580 B.n71 163.367
R1916 B.n580 B.n579 163.367
R1917 B.n579 B.n578 163.367
R1918 B.n578 B.n73 163.367
R1919 B.n574 B.n73 163.367
R1920 B.n574 B.n573 163.367
R1921 B.n573 B.n572 163.367
R1922 B.n572 B.n75 163.367
R1923 B.n568 B.n75 163.367
R1924 B.n568 B.n567 163.367
R1925 B.n567 B.n566 163.367
R1926 B.n566 B.n77 163.367
R1927 B.n562 B.n77 163.367
R1928 B.n562 B.n561 163.367
R1929 B.n561 B.n560 163.367
R1930 B.n560 B.n79 163.367
R1931 B.n556 B.n79 163.367
R1932 B.n556 B.n555 163.367
R1933 B.n150 B.n149 59.5399
R1934 B.n337 B.n157 59.5399
R1935 B.n641 B.n49 59.5399
R1936 B.n56 B.n55 59.5399
R1937 B.n149 B.n148 45.9641
R1938 B.n157 B.n156 45.9641
R1939 B.n49 B.n48 45.9641
R1940 B.n55 B.n54 45.9641
R1941 B.n714 B.n713 31.6883
R1942 B.n553 B.n80 31.6883
R1943 B.n425 B.n124 31.6883
R1944 B.n265 B.n264 31.6883
R1945 B B.n779 18.0485
R1946 B.n713 B.n24 10.6151
R1947 B.n709 B.n24 10.6151
R1948 B.n709 B.n708 10.6151
R1949 B.n708 B.n707 10.6151
R1950 B.n707 B.n26 10.6151
R1951 B.n703 B.n26 10.6151
R1952 B.n703 B.n702 10.6151
R1953 B.n702 B.n701 10.6151
R1954 B.n701 B.n28 10.6151
R1955 B.n697 B.n28 10.6151
R1956 B.n697 B.n696 10.6151
R1957 B.n696 B.n695 10.6151
R1958 B.n695 B.n30 10.6151
R1959 B.n691 B.n30 10.6151
R1960 B.n691 B.n690 10.6151
R1961 B.n690 B.n689 10.6151
R1962 B.n689 B.n32 10.6151
R1963 B.n685 B.n32 10.6151
R1964 B.n685 B.n684 10.6151
R1965 B.n684 B.n683 10.6151
R1966 B.n683 B.n34 10.6151
R1967 B.n679 B.n34 10.6151
R1968 B.n679 B.n678 10.6151
R1969 B.n678 B.n677 10.6151
R1970 B.n677 B.n36 10.6151
R1971 B.n673 B.n36 10.6151
R1972 B.n673 B.n672 10.6151
R1973 B.n672 B.n671 10.6151
R1974 B.n671 B.n38 10.6151
R1975 B.n667 B.n38 10.6151
R1976 B.n667 B.n666 10.6151
R1977 B.n666 B.n665 10.6151
R1978 B.n665 B.n40 10.6151
R1979 B.n661 B.n40 10.6151
R1980 B.n661 B.n660 10.6151
R1981 B.n660 B.n659 10.6151
R1982 B.n659 B.n42 10.6151
R1983 B.n655 B.n42 10.6151
R1984 B.n655 B.n654 10.6151
R1985 B.n654 B.n653 10.6151
R1986 B.n653 B.n44 10.6151
R1987 B.n649 B.n44 10.6151
R1988 B.n649 B.n648 10.6151
R1989 B.n648 B.n647 10.6151
R1990 B.n647 B.n46 10.6151
R1991 B.n643 B.n46 10.6151
R1992 B.n643 B.n642 10.6151
R1993 B.n640 B.n50 10.6151
R1994 B.n636 B.n50 10.6151
R1995 B.n636 B.n635 10.6151
R1996 B.n635 B.n634 10.6151
R1997 B.n634 B.n52 10.6151
R1998 B.n630 B.n52 10.6151
R1999 B.n630 B.n629 10.6151
R2000 B.n629 B.n628 10.6151
R2001 B.n625 B.n624 10.6151
R2002 B.n624 B.n623 10.6151
R2003 B.n623 B.n58 10.6151
R2004 B.n619 B.n58 10.6151
R2005 B.n619 B.n618 10.6151
R2006 B.n618 B.n617 10.6151
R2007 B.n617 B.n60 10.6151
R2008 B.n613 B.n60 10.6151
R2009 B.n613 B.n612 10.6151
R2010 B.n612 B.n611 10.6151
R2011 B.n611 B.n62 10.6151
R2012 B.n607 B.n62 10.6151
R2013 B.n607 B.n606 10.6151
R2014 B.n606 B.n605 10.6151
R2015 B.n605 B.n64 10.6151
R2016 B.n601 B.n64 10.6151
R2017 B.n601 B.n600 10.6151
R2018 B.n600 B.n599 10.6151
R2019 B.n599 B.n66 10.6151
R2020 B.n595 B.n66 10.6151
R2021 B.n595 B.n594 10.6151
R2022 B.n594 B.n593 10.6151
R2023 B.n593 B.n68 10.6151
R2024 B.n589 B.n68 10.6151
R2025 B.n589 B.n588 10.6151
R2026 B.n588 B.n587 10.6151
R2027 B.n587 B.n70 10.6151
R2028 B.n583 B.n70 10.6151
R2029 B.n583 B.n582 10.6151
R2030 B.n582 B.n581 10.6151
R2031 B.n581 B.n72 10.6151
R2032 B.n577 B.n72 10.6151
R2033 B.n577 B.n576 10.6151
R2034 B.n576 B.n575 10.6151
R2035 B.n575 B.n74 10.6151
R2036 B.n571 B.n74 10.6151
R2037 B.n571 B.n570 10.6151
R2038 B.n570 B.n569 10.6151
R2039 B.n569 B.n76 10.6151
R2040 B.n565 B.n76 10.6151
R2041 B.n565 B.n564 10.6151
R2042 B.n564 B.n563 10.6151
R2043 B.n563 B.n78 10.6151
R2044 B.n559 B.n78 10.6151
R2045 B.n559 B.n558 10.6151
R2046 B.n558 B.n557 10.6151
R2047 B.n557 B.n80 10.6151
R2048 B.n426 B.n425 10.6151
R2049 B.n427 B.n426 10.6151
R2050 B.n427 B.n122 10.6151
R2051 B.n431 B.n122 10.6151
R2052 B.n432 B.n431 10.6151
R2053 B.n433 B.n432 10.6151
R2054 B.n433 B.n120 10.6151
R2055 B.n437 B.n120 10.6151
R2056 B.n438 B.n437 10.6151
R2057 B.n439 B.n438 10.6151
R2058 B.n439 B.n118 10.6151
R2059 B.n443 B.n118 10.6151
R2060 B.n444 B.n443 10.6151
R2061 B.n445 B.n444 10.6151
R2062 B.n445 B.n116 10.6151
R2063 B.n449 B.n116 10.6151
R2064 B.n450 B.n449 10.6151
R2065 B.n451 B.n450 10.6151
R2066 B.n451 B.n114 10.6151
R2067 B.n455 B.n114 10.6151
R2068 B.n456 B.n455 10.6151
R2069 B.n457 B.n456 10.6151
R2070 B.n457 B.n112 10.6151
R2071 B.n461 B.n112 10.6151
R2072 B.n462 B.n461 10.6151
R2073 B.n463 B.n462 10.6151
R2074 B.n463 B.n110 10.6151
R2075 B.n467 B.n110 10.6151
R2076 B.n468 B.n467 10.6151
R2077 B.n469 B.n468 10.6151
R2078 B.n469 B.n108 10.6151
R2079 B.n473 B.n108 10.6151
R2080 B.n474 B.n473 10.6151
R2081 B.n475 B.n474 10.6151
R2082 B.n475 B.n106 10.6151
R2083 B.n479 B.n106 10.6151
R2084 B.n480 B.n479 10.6151
R2085 B.n481 B.n480 10.6151
R2086 B.n481 B.n104 10.6151
R2087 B.n485 B.n104 10.6151
R2088 B.n486 B.n485 10.6151
R2089 B.n487 B.n486 10.6151
R2090 B.n487 B.n102 10.6151
R2091 B.n491 B.n102 10.6151
R2092 B.n492 B.n491 10.6151
R2093 B.n493 B.n492 10.6151
R2094 B.n493 B.n100 10.6151
R2095 B.n497 B.n100 10.6151
R2096 B.n498 B.n497 10.6151
R2097 B.n499 B.n498 10.6151
R2098 B.n499 B.n98 10.6151
R2099 B.n503 B.n98 10.6151
R2100 B.n504 B.n503 10.6151
R2101 B.n505 B.n504 10.6151
R2102 B.n505 B.n96 10.6151
R2103 B.n509 B.n96 10.6151
R2104 B.n510 B.n509 10.6151
R2105 B.n511 B.n510 10.6151
R2106 B.n511 B.n94 10.6151
R2107 B.n515 B.n94 10.6151
R2108 B.n516 B.n515 10.6151
R2109 B.n517 B.n516 10.6151
R2110 B.n517 B.n92 10.6151
R2111 B.n521 B.n92 10.6151
R2112 B.n522 B.n521 10.6151
R2113 B.n523 B.n522 10.6151
R2114 B.n523 B.n90 10.6151
R2115 B.n527 B.n90 10.6151
R2116 B.n528 B.n527 10.6151
R2117 B.n529 B.n528 10.6151
R2118 B.n529 B.n88 10.6151
R2119 B.n533 B.n88 10.6151
R2120 B.n534 B.n533 10.6151
R2121 B.n535 B.n534 10.6151
R2122 B.n535 B.n86 10.6151
R2123 B.n539 B.n86 10.6151
R2124 B.n540 B.n539 10.6151
R2125 B.n541 B.n540 10.6151
R2126 B.n541 B.n84 10.6151
R2127 B.n545 B.n84 10.6151
R2128 B.n546 B.n545 10.6151
R2129 B.n547 B.n546 10.6151
R2130 B.n547 B.n82 10.6151
R2131 B.n551 B.n82 10.6151
R2132 B.n552 B.n551 10.6151
R2133 B.n553 B.n552 10.6151
R2134 B.n265 B.n180 10.6151
R2135 B.n269 B.n180 10.6151
R2136 B.n270 B.n269 10.6151
R2137 B.n271 B.n270 10.6151
R2138 B.n271 B.n178 10.6151
R2139 B.n275 B.n178 10.6151
R2140 B.n276 B.n275 10.6151
R2141 B.n277 B.n276 10.6151
R2142 B.n277 B.n176 10.6151
R2143 B.n281 B.n176 10.6151
R2144 B.n282 B.n281 10.6151
R2145 B.n283 B.n282 10.6151
R2146 B.n283 B.n174 10.6151
R2147 B.n287 B.n174 10.6151
R2148 B.n288 B.n287 10.6151
R2149 B.n289 B.n288 10.6151
R2150 B.n289 B.n172 10.6151
R2151 B.n293 B.n172 10.6151
R2152 B.n294 B.n293 10.6151
R2153 B.n295 B.n294 10.6151
R2154 B.n295 B.n170 10.6151
R2155 B.n299 B.n170 10.6151
R2156 B.n300 B.n299 10.6151
R2157 B.n301 B.n300 10.6151
R2158 B.n301 B.n168 10.6151
R2159 B.n305 B.n168 10.6151
R2160 B.n306 B.n305 10.6151
R2161 B.n307 B.n306 10.6151
R2162 B.n307 B.n166 10.6151
R2163 B.n311 B.n166 10.6151
R2164 B.n312 B.n311 10.6151
R2165 B.n313 B.n312 10.6151
R2166 B.n313 B.n164 10.6151
R2167 B.n317 B.n164 10.6151
R2168 B.n318 B.n317 10.6151
R2169 B.n319 B.n318 10.6151
R2170 B.n319 B.n162 10.6151
R2171 B.n323 B.n162 10.6151
R2172 B.n324 B.n323 10.6151
R2173 B.n325 B.n324 10.6151
R2174 B.n325 B.n160 10.6151
R2175 B.n329 B.n160 10.6151
R2176 B.n330 B.n329 10.6151
R2177 B.n331 B.n330 10.6151
R2178 B.n331 B.n158 10.6151
R2179 B.n335 B.n158 10.6151
R2180 B.n336 B.n335 10.6151
R2181 B.n338 B.n154 10.6151
R2182 B.n342 B.n154 10.6151
R2183 B.n343 B.n342 10.6151
R2184 B.n344 B.n343 10.6151
R2185 B.n344 B.n152 10.6151
R2186 B.n348 B.n152 10.6151
R2187 B.n349 B.n348 10.6151
R2188 B.n350 B.n349 10.6151
R2189 B.n354 B.n353 10.6151
R2190 B.n355 B.n354 10.6151
R2191 B.n355 B.n146 10.6151
R2192 B.n359 B.n146 10.6151
R2193 B.n360 B.n359 10.6151
R2194 B.n361 B.n360 10.6151
R2195 B.n361 B.n144 10.6151
R2196 B.n365 B.n144 10.6151
R2197 B.n366 B.n365 10.6151
R2198 B.n367 B.n366 10.6151
R2199 B.n367 B.n142 10.6151
R2200 B.n371 B.n142 10.6151
R2201 B.n372 B.n371 10.6151
R2202 B.n373 B.n372 10.6151
R2203 B.n373 B.n140 10.6151
R2204 B.n377 B.n140 10.6151
R2205 B.n378 B.n377 10.6151
R2206 B.n379 B.n378 10.6151
R2207 B.n379 B.n138 10.6151
R2208 B.n383 B.n138 10.6151
R2209 B.n384 B.n383 10.6151
R2210 B.n385 B.n384 10.6151
R2211 B.n385 B.n136 10.6151
R2212 B.n389 B.n136 10.6151
R2213 B.n390 B.n389 10.6151
R2214 B.n391 B.n390 10.6151
R2215 B.n391 B.n134 10.6151
R2216 B.n395 B.n134 10.6151
R2217 B.n396 B.n395 10.6151
R2218 B.n397 B.n396 10.6151
R2219 B.n397 B.n132 10.6151
R2220 B.n401 B.n132 10.6151
R2221 B.n402 B.n401 10.6151
R2222 B.n403 B.n402 10.6151
R2223 B.n403 B.n130 10.6151
R2224 B.n407 B.n130 10.6151
R2225 B.n408 B.n407 10.6151
R2226 B.n409 B.n408 10.6151
R2227 B.n409 B.n128 10.6151
R2228 B.n413 B.n128 10.6151
R2229 B.n414 B.n413 10.6151
R2230 B.n415 B.n414 10.6151
R2231 B.n415 B.n126 10.6151
R2232 B.n419 B.n126 10.6151
R2233 B.n420 B.n419 10.6151
R2234 B.n421 B.n420 10.6151
R2235 B.n421 B.n124 10.6151
R2236 B.n264 B.n263 10.6151
R2237 B.n263 B.n182 10.6151
R2238 B.n259 B.n182 10.6151
R2239 B.n259 B.n258 10.6151
R2240 B.n258 B.n257 10.6151
R2241 B.n257 B.n184 10.6151
R2242 B.n253 B.n184 10.6151
R2243 B.n253 B.n252 10.6151
R2244 B.n252 B.n251 10.6151
R2245 B.n251 B.n186 10.6151
R2246 B.n247 B.n186 10.6151
R2247 B.n247 B.n246 10.6151
R2248 B.n246 B.n245 10.6151
R2249 B.n245 B.n188 10.6151
R2250 B.n241 B.n188 10.6151
R2251 B.n241 B.n240 10.6151
R2252 B.n240 B.n239 10.6151
R2253 B.n239 B.n190 10.6151
R2254 B.n235 B.n190 10.6151
R2255 B.n235 B.n234 10.6151
R2256 B.n234 B.n233 10.6151
R2257 B.n233 B.n192 10.6151
R2258 B.n229 B.n192 10.6151
R2259 B.n229 B.n228 10.6151
R2260 B.n228 B.n227 10.6151
R2261 B.n227 B.n194 10.6151
R2262 B.n223 B.n194 10.6151
R2263 B.n223 B.n222 10.6151
R2264 B.n222 B.n221 10.6151
R2265 B.n221 B.n196 10.6151
R2266 B.n217 B.n196 10.6151
R2267 B.n217 B.n216 10.6151
R2268 B.n216 B.n215 10.6151
R2269 B.n215 B.n198 10.6151
R2270 B.n211 B.n198 10.6151
R2271 B.n211 B.n210 10.6151
R2272 B.n210 B.n209 10.6151
R2273 B.n209 B.n200 10.6151
R2274 B.n205 B.n200 10.6151
R2275 B.n205 B.n204 10.6151
R2276 B.n204 B.n203 10.6151
R2277 B.n203 B.n0 10.6151
R2278 B.n775 B.n1 10.6151
R2279 B.n775 B.n774 10.6151
R2280 B.n774 B.n773 10.6151
R2281 B.n773 B.n4 10.6151
R2282 B.n769 B.n4 10.6151
R2283 B.n769 B.n768 10.6151
R2284 B.n768 B.n767 10.6151
R2285 B.n767 B.n6 10.6151
R2286 B.n763 B.n6 10.6151
R2287 B.n763 B.n762 10.6151
R2288 B.n762 B.n761 10.6151
R2289 B.n761 B.n8 10.6151
R2290 B.n757 B.n8 10.6151
R2291 B.n757 B.n756 10.6151
R2292 B.n756 B.n755 10.6151
R2293 B.n755 B.n10 10.6151
R2294 B.n751 B.n10 10.6151
R2295 B.n751 B.n750 10.6151
R2296 B.n750 B.n749 10.6151
R2297 B.n749 B.n12 10.6151
R2298 B.n745 B.n12 10.6151
R2299 B.n745 B.n744 10.6151
R2300 B.n744 B.n743 10.6151
R2301 B.n743 B.n14 10.6151
R2302 B.n739 B.n14 10.6151
R2303 B.n739 B.n738 10.6151
R2304 B.n738 B.n737 10.6151
R2305 B.n737 B.n16 10.6151
R2306 B.n733 B.n16 10.6151
R2307 B.n733 B.n732 10.6151
R2308 B.n732 B.n731 10.6151
R2309 B.n731 B.n18 10.6151
R2310 B.n727 B.n18 10.6151
R2311 B.n727 B.n726 10.6151
R2312 B.n726 B.n725 10.6151
R2313 B.n725 B.n20 10.6151
R2314 B.n721 B.n20 10.6151
R2315 B.n721 B.n720 10.6151
R2316 B.n720 B.n719 10.6151
R2317 B.n719 B.n22 10.6151
R2318 B.n715 B.n22 10.6151
R2319 B.n715 B.n714 10.6151
R2320 B.n641 B.n640 6.5566
R2321 B.n628 B.n56 6.5566
R2322 B.n338 B.n337 6.5566
R2323 B.n350 B.n150 6.5566
R2324 B.n642 B.n641 4.05904
R2325 B.n625 B.n56 4.05904
R2326 B.n337 B.n336 4.05904
R2327 B.n353 B.n150 4.05904
R2328 B.n779 B.n0 2.81026
R2329 B.n779 B.n1 2.81026
C0 VDD2 B 1.61347f
C1 VN B 1.11579f
C2 VDD2 w_n3340_n3780# 1.91796f
C3 VN w_n3340_n3780# 6.69686f
C4 VDD1 VDD2 1.48535f
C5 VN VDD1 0.150292f
C6 VN VDD2 9.58251f
C7 VTAIL B 5.36053f
C8 VTAIL w_n3340_n3780# 4.65182f
C9 VTAIL VDD1 8.88526f
C10 VTAIL VDD2 8.93592f
C11 VN VTAIL 9.708731f
C12 B VP 1.8369f
C13 w_n3340_n3780# VP 7.12881f
C14 VDD1 VP 9.89077f
C15 VDD2 VP 0.459658f
C16 VN VP 7.36867f
C17 w_n3340_n3780# B 9.835589f
C18 VDD1 B 1.53507f
C19 VDD1 w_n3340_n3780# 1.82674f
C20 VTAIL VP 9.722839f
C21 VDD2 VSUBS 1.687866f
C22 VDD1 VSUBS 2.23763f
C23 VTAIL VSUBS 1.335106f
C24 VN VSUBS 6.12546f
C25 VP VSUBS 3.089209f
C26 B VSUBS 4.549396f
C27 w_n3340_n3780# VSUBS 0.154989p
C28 B.n0 VSUBS 0.004289f
C29 B.n1 VSUBS 0.004289f
C30 B.n2 VSUBS 0.006783f
C31 B.n3 VSUBS 0.006783f
C32 B.n4 VSUBS 0.006783f
C33 B.n5 VSUBS 0.006783f
C34 B.n6 VSUBS 0.006783f
C35 B.n7 VSUBS 0.006783f
C36 B.n8 VSUBS 0.006783f
C37 B.n9 VSUBS 0.006783f
C38 B.n10 VSUBS 0.006783f
C39 B.n11 VSUBS 0.006783f
C40 B.n12 VSUBS 0.006783f
C41 B.n13 VSUBS 0.006783f
C42 B.n14 VSUBS 0.006783f
C43 B.n15 VSUBS 0.006783f
C44 B.n16 VSUBS 0.006783f
C45 B.n17 VSUBS 0.006783f
C46 B.n18 VSUBS 0.006783f
C47 B.n19 VSUBS 0.006783f
C48 B.n20 VSUBS 0.006783f
C49 B.n21 VSUBS 0.006783f
C50 B.n22 VSUBS 0.006783f
C51 B.n23 VSUBS 0.015168f
C52 B.n24 VSUBS 0.006783f
C53 B.n25 VSUBS 0.006783f
C54 B.n26 VSUBS 0.006783f
C55 B.n27 VSUBS 0.006783f
C56 B.n28 VSUBS 0.006783f
C57 B.n29 VSUBS 0.006783f
C58 B.n30 VSUBS 0.006783f
C59 B.n31 VSUBS 0.006783f
C60 B.n32 VSUBS 0.006783f
C61 B.n33 VSUBS 0.006783f
C62 B.n34 VSUBS 0.006783f
C63 B.n35 VSUBS 0.006783f
C64 B.n36 VSUBS 0.006783f
C65 B.n37 VSUBS 0.006783f
C66 B.n38 VSUBS 0.006783f
C67 B.n39 VSUBS 0.006783f
C68 B.n40 VSUBS 0.006783f
C69 B.n41 VSUBS 0.006783f
C70 B.n42 VSUBS 0.006783f
C71 B.n43 VSUBS 0.006783f
C72 B.n44 VSUBS 0.006783f
C73 B.n45 VSUBS 0.006783f
C74 B.n46 VSUBS 0.006783f
C75 B.n47 VSUBS 0.006783f
C76 B.t11 VSUBS 0.249701f
C77 B.t10 VSUBS 0.275664f
C78 B.t9 VSUBS 1.23119f
C79 B.n48 VSUBS 0.421884f
C80 B.n49 VSUBS 0.268736f
C81 B.n50 VSUBS 0.006783f
C82 B.n51 VSUBS 0.006783f
C83 B.n52 VSUBS 0.006783f
C84 B.n53 VSUBS 0.006783f
C85 B.t8 VSUBS 0.249704f
C86 B.t7 VSUBS 0.275667f
C87 B.t6 VSUBS 1.23119f
C88 B.n54 VSUBS 0.421881f
C89 B.n55 VSUBS 0.268732f
C90 B.n56 VSUBS 0.015716f
C91 B.n57 VSUBS 0.006783f
C92 B.n58 VSUBS 0.006783f
C93 B.n59 VSUBS 0.006783f
C94 B.n60 VSUBS 0.006783f
C95 B.n61 VSUBS 0.006783f
C96 B.n62 VSUBS 0.006783f
C97 B.n63 VSUBS 0.006783f
C98 B.n64 VSUBS 0.006783f
C99 B.n65 VSUBS 0.006783f
C100 B.n66 VSUBS 0.006783f
C101 B.n67 VSUBS 0.006783f
C102 B.n68 VSUBS 0.006783f
C103 B.n69 VSUBS 0.006783f
C104 B.n70 VSUBS 0.006783f
C105 B.n71 VSUBS 0.006783f
C106 B.n72 VSUBS 0.006783f
C107 B.n73 VSUBS 0.006783f
C108 B.n74 VSUBS 0.006783f
C109 B.n75 VSUBS 0.006783f
C110 B.n76 VSUBS 0.006783f
C111 B.n77 VSUBS 0.006783f
C112 B.n78 VSUBS 0.006783f
C113 B.n79 VSUBS 0.006783f
C114 B.n80 VSUBS 0.015128f
C115 B.n81 VSUBS 0.006783f
C116 B.n82 VSUBS 0.006783f
C117 B.n83 VSUBS 0.006783f
C118 B.n84 VSUBS 0.006783f
C119 B.n85 VSUBS 0.006783f
C120 B.n86 VSUBS 0.006783f
C121 B.n87 VSUBS 0.006783f
C122 B.n88 VSUBS 0.006783f
C123 B.n89 VSUBS 0.006783f
C124 B.n90 VSUBS 0.006783f
C125 B.n91 VSUBS 0.006783f
C126 B.n92 VSUBS 0.006783f
C127 B.n93 VSUBS 0.006783f
C128 B.n94 VSUBS 0.006783f
C129 B.n95 VSUBS 0.006783f
C130 B.n96 VSUBS 0.006783f
C131 B.n97 VSUBS 0.006783f
C132 B.n98 VSUBS 0.006783f
C133 B.n99 VSUBS 0.006783f
C134 B.n100 VSUBS 0.006783f
C135 B.n101 VSUBS 0.006783f
C136 B.n102 VSUBS 0.006783f
C137 B.n103 VSUBS 0.006783f
C138 B.n104 VSUBS 0.006783f
C139 B.n105 VSUBS 0.006783f
C140 B.n106 VSUBS 0.006783f
C141 B.n107 VSUBS 0.006783f
C142 B.n108 VSUBS 0.006783f
C143 B.n109 VSUBS 0.006783f
C144 B.n110 VSUBS 0.006783f
C145 B.n111 VSUBS 0.006783f
C146 B.n112 VSUBS 0.006783f
C147 B.n113 VSUBS 0.006783f
C148 B.n114 VSUBS 0.006783f
C149 B.n115 VSUBS 0.006783f
C150 B.n116 VSUBS 0.006783f
C151 B.n117 VSUBS 0.006783f
C152 B.n118 VSUBS 0.006783f
C153 B.n119 VSUBS 0.006783f
C154 B.n120 VSUBS 0.006783f
C155 B.n121 VSUBS 0.006783f
C156 B.n122 VSUBS 0.006783f
C157 B.n123 VSUBS 0.006783f
C158 B.n124 VSUBS 0.015954f
C159 B.n125 VSUBS 0.006783f
C160 B.n126 VSUBS 0.006783f
C161 B.n127 VSUBS 0.006783f
C162 B.n128 VSUBS 0.006783f
C163 B.n129 VSUBS 0.006783f
C164 B.n130 VSUBS 0.006783f
C165 B.n131 VSUBS 0.006783f
C166 B.n132 VSUBS 0.006783f
C167 B.n133 VSUBS 0.006783f
C168 B.n134 VSUBS 0.006783f
C169 B.n135 VSUBS 0.006783f
C170 B.n136 VSUBS 0.006783f
C171 B.n137 VSUBS 0.006783f
C172 B.n138 VSUBS 0.006783f
C173 B.n139 VSUBS 0.006783f
C174 B.n140 VSUBS 0.006783f
C175 B.n141 VSUBS 0.006783f
C176 B.n142 VSUBS 0.006783f
C177 B.n143 VSUBS 0.006783f
C178 B.n144 VSUBS 0.006783f
C179 B.n145 VSUBS 0.006783f
C180 B.n146 VSUBS 0.006783f
C181 B.n147 VSUBS 0.006783f
C182 B.t1 VSUBS 0.249704f
C183 B.t2 VSUBS 0.275667f
C184 B.t0 VSUBS 1.23119f
C185 B.n148 VSUBS 0.421881f
C186 B.n149 VSUBS 0.268732f
C187 B.n150 VSUBS 0.015716f
C188 B.n151 VSUBS 0.006783f
C189 B.n152 VSUBS 0.006783f
C190 B.n153 VSUBS 0.006783f
C191 B.n154 VSUBS 0.006783f
C192 B.n155 VSUBS 0.006783f
C193 B.t4 VSUBS 0.249701f
C194 B.t5 VSUBS 0.275664f
C195 B.t3 VSUBS 1.23119f
C196 B.n156 VSUBS 0.421884f
C197 B.n157 VSUBS 0.268736f
C198 B.n158 VSUBS 0.006783f
C199 B.n159 VSUBS 0.006783f
C200 B.n160 VSUBS 0.006783f
C201 B.n161 VSUBS 0.006783f
C202 B.n162 VSUBS 0.006783f
C203 B.n163 VSUBS 0.006783f
C204 B.n164 VSUBS 0.006783f
C205 B.n165 VSUBS 0.006783f
C206 B.n166 VSUBS 0.006783f
C207 B.n167 VSUBS 0.006783f
C208 B.n168 VSUBS 0.006783f
C209 B.n169 VSUBS 0.006783f
C210 B.n170 VSUBS 0.006783f
C211 B.n171 VSUBS 0.006783f
C212 B.n172 VSUBS 0.006783f
C213 B.n173 VSUBS 0.006783f
C214 B.n174 VSUBS 0.006783f
C215 B.n175 VSUBS 0.006783f
C216 B.n176 VSUBS 0.006783f
C217 B.n177 VSUBS 0.006783f
C218 B.n178 VSUBS 0.006783f
C219 B.n179 VSUBS 0.006783f
C220 B.n180 VSUBS 0.006783f
C221 B.n181 VSUBS 0.015168f
C222 B.n182 VSUBS 0.006783f
C223 B.n183 VSUBS 0.006783f
C224 B.n184 VSUBS 0.006783f
C225 B.n185 VSUBS 0.006783f
C226 B.n186 VSUBS 0.006783f
C227 B.n187 VSUBS 0.006783f
C228 B.n188 VSUBS 0.006783f
C229 B.n189 VSUBS 0.006783f
C230 B.n190 VSUBS 0.006783f
C231 B.n191 VSUBS 0.006783f
C232 B.n192 VSUBS 0.006783f
C233 B.n193 VSUBS 0.006783f
C234 B.n194 VSUBS 0.006783f
C235 B.n195 VSUBS 0.006783f
C236 B.n196 VSUBS 0.006783f
C237 B.n197 VSUBS 0.006783f
C238 B.n198 VSUBS 0.006783f
C239 B.n199 VSUBS 0.006783f
C240 B.n200 VSUBS 0.006783f
C241 B.n201 VSUBS 0.006783f
C242 B.n202 VSUBS 0.006783f
C243 B.n203 VSUBS 0.006783f
C244 B.n204 VSUBS 0.006783f
C245 B.n205 VSUBS 0.006783f
C246 B.n206 VSUBS 0.006783f
C247 B.n207 VSUBS 0.006783f
C248 B.n208 VSUBS 0.006783f
C249 B.n209 VSUBS 0.006783f
C250 B.n210 VSUBS 0.006783f
C251 B.n211 VSUBS 0.006783f
C252 B.n212 VSUBS 0.006783f
C253 B.n213 VSUBS 0.006783f
C254 B.n214 VSUBS 0.006783f
C255 B.n215 VSUBS 0.006783f
C256 B.n216 VSUBS 0.006783f
C257 B.n217 VSUBS 0.006783f
C258 B.n218 VSUBS 0.006783f
C259 B.n219 VSUBS 0.006783f
C260 B.n220 VSUBS 0.006783f
C261 B.n221 VSUBS 0.006783f
C262 B.n222 VSUBS 0.006783f
C263 B.n223 VSUBS 0.006783f
C264 B.n224 VSUBS 0.006783f
C265 B.n225 VSUBS 0.006783f
C266 B.n226 VSUBS 0.006783f
C267 B.n227 VSUBS 0.006783f
C268 B.n228 VSUBS 0.006783f
C269 B.n229 VSUBS 0.006783f
C270 B.n230 VSUBS 0.006783f
C271 B.n231 VSUBS 0.006783f
C272 B.n232 VSUBS 0.006783f
C273 B.n233 VSUBS 0.006783f
C274 B.n234 VSUBS 0.006783f
C275 B.n235 VSUBS 0.006783f
C276 B.n236 VSUBS 0.006783f
C277 B.n237 VSUBS 0.006783f
C278 B.n238 VSUBS 0.006783f
C279 B.n239 VSUBS 0.006783f
C280 B.n240 VSUBS 0.006783f
C281 B.n241 VSUBS 0.006783f
C282 B.n242 VSUBS 0.006783f
C283 B.n243 VSUBS 0.006783f
C284 B.n244 VSUBS 0.006783f
C285 B.n245 VSUBS 0.006783f
C286 B.n246 VSUBS 0.006783f
C287 B.n247 VSUBS 0.006783f
C288 B.n248 VSUBS 0.006783f
C289 B.n249 VSUBS 0.006783f
C290 B.n250 VSUBS 0.006783f
C291 B.n251 VSUBS 0.006783f
C292 B.n252 VSUBS 0.006783f
C293 B.n253 VSUBS 0.006783f
C294 B.n254 VSUBS 0.006783f
C295 B.n255 VSUBS 0.006783f
C296 B.n256 VSUBS 0.006783f
C297 B.n257 VSUBS 0.006783f
C298 B.n258 VSUBS 0.006783f
C299 B.n259 VSUBS 0.006783f
C300 B.n260 VSUBS 0.006783f
C301 B.n261 VSUBS 0.006783f
C302 B.n262 VSUBS 0.006783f
C303 B.n263 VSUBS 0.006783f
C304 B.n264 VSUBS 0.015168f
C305 B.n265 VSUBS 0.015954f
C306 B.n266 VSUBS 0.015954f
C307 B.n267 VSUBS 0.006783f
C308 B.n268 VSUBS 0.006783f
C309 B.n269 VSUBS 0.006783f
C310 B.n270 VSUBS 0.006783f
C311 B.n271 VSUBS 0.006783f
C312 B.n272 VSUBS 0.006783f
C313 B.n273 VSUBS 0.006783f
C314 B.n274 VSUBS 0.006783f
C315 B.n275 VSUBS 0.006783f
C316 B.n276 VSUBS 0.006783f
C317 B.n277 VSUBS 0.006783f
C318 B.n278 VSUBS 0.006783f
C319 B.n279 VSUBS 0.006783f
C320 B.n280 VSUBS 0.006783f
C321 B.n281 VSUBS 0.006783f
C322 B.n282 VSUBS 0.006783f
C323 B.n283 VSUBS 0.006783f
C324 B.n284 VSUBS 0.006783f
C325 B.n285 VSUBS 0.006783f
C326 B.n286 VSUBS 0.006783f
C327 B.n287 VSUBS 0.006783f
C328 B.n288 VSUBS 0.006783f
C329 B.n289 VSUBS 0.006783f
C330 B.n290 VSUBS 0.006783f
C331 B.n291 VSUBS 0.006783f
C332 B.n292 VSUBS 0.006783f
C333 B.n293 VSUBS 0.006783f
C334 B.n294 VSUBS 0.006783f
C335 B.n295 VSUBS 0.006783f
C336 B.n296 VSUBS 0.006783f
C337 B.n297 VSUBS 0.006783f
C338 B.n298 VSUBS 0.006783f
C339 B.n299 VSUBS 0.006783f
C340 B.n300 VSUBS 0.006783f
C341 B.n301 VSUBS 0.006783f
C342 B.n302 VSUBS 0.006783f
C343 B.n303 VSUBS 0.006783f
C344 B.n304 VSUBS 0.006783f
C345 B.n305 VSUBS 0.006783f
C346 B.n306 VSUBS 0.006783f
C347 B.n307 VSUBS 0.006783f
C348 B.n308 VSUBS 0.006783f
C349 B.n309 VSUBS 0.006783f
C350 B.n310 VSUBS 0.006783f
C351 B.n311 VSUBS 0.006783f
C352 B.n312 VSUBS 0.006783f
C353 B.n313 VSUBS 0.006783f
C354 B.n314 VSUBS 0.006783f
C355 B.n315 VSUBS 0.006783f
C356 B.n316 VSUBS 0.006783f
C357 B.n317 VSUBS 0.006783f
C358 B.n318 VSUBS 0.006783f
C359 B.n319 VSUBS 0.006783f
C360 B.n320 VSUBS 0.006783f
C361 B.n321 VSUBS 0.006783f
C362 B.n322 VSUBS 0.006783f
C363 B.n323 VSUBS 0.006783f
C364 B.n324 VSUBS 0.006783f
C365 B.n325 VSUBS 0.006783f
C366 B.n326 VSUBS 0.006783f
C367 B.n327 VSUBS 0.006783f
C368 B.n328 VSUBS 0.006783f
C369 B.n329 VSUBS 0.006783f
C370 B.n330 VSUBS 0.006783f
C371 B.n331 VSUBS 0.006783f
C372 B.n332 VSUBS 0.006783f
C373 B.n333 VSUBS 0.006783f
C374 B.n334 VSUBS 0.006783f
C375 B.n335 VSUBS 0.006783f
C376 B.n336 VSUBS 0.004688f
C377 B.n337 VSUBS 0.015716f
C378 B.n338 VSUBS 0.005486f
C379 B.n339 VSUBS 0.006783f
C380 B.n340 VSUBS 0.006783f
C381 B.n341 VSUBS 0.006783f
C382 B.n342 VSUBS 0.006783f
C383 B.n343 VSUBS 0.006783f
C384 B.n344 VSUBS 0.006783f
C385 B.n345 VSUBS 0.006783f
C386 B.n346 VSUBS 0.006783f
C387 B.n347 VSUBS 0.006783f
C388 B.n348 VSUBS 0.006783f
C389 B.n349 VSUBS 0.006783f
C390 B.n350 VSUBS 0.005486f
C391 B.n351 VSUBS 0.006783f
C392 B.n352 VSUBS 0.006783f
C393 B.n353 VSUBS 0.004688f
C394 B.n354 VSUBS 0.006783f
C395 B.n355 VSUBS 0.006783f
C396 B.n356 VSUBS 0.006783f
C397 B.n357 VSUBS 0.006783f
C398 B.n358 VSUBS 0.006783f
C399 B.n359 VSUBS 0.006783f
C400 B.n360 VSUBS 0.006783f
C401 B.n361 VSUBS 0.006783f
C402 B.n362 VSUBS 0.006783f
C403 B.n363 VSUBS 0.006783f
C404 B.n364 VSUBS 0.006783f
C405 B.n365 VSUBS 0.006783f
C406 B.n366 VSUBS 0.006783f
C407 B.n367 VSUBS 0.006783f
C408 B.n368 VSUBS 0.006783f
C409 B.n369 VSUBS 0.006783f
C410 B.n370 VSUBS 0.006783f
C411 B.n371 VSUBS 0.006783f
C412 B.n372 VSUBS 0.006783f
C413 B.n373 VSUBS 0.006783f
C414 B.n374 VSUBS 0.006783f
C415 B.n375 VSUBS 0.006783f
C416 B.n376 VSUBS 0.006783f
C417 B.n377 VSUBS 0.006783f
C418 B.n378 VSUBS 0.006783f
C419 B.n379 VSUBS 0.006783f
C420 B.n380 VSUBS 0.006783f
C421 B.n381 VSUBS 0.006783f
C422 B.n382 VSUBS 0.006783f
C423 B.n383 VSUBS 0.006783f
C424 B.n384 VSUBS 0.006783f
C425 B.n385 VSUBS 0.006783f
C426 B.n386 VSUBS 0.006783f
C427 B.n387 VSUBS 0.006783f
C428 B.n388 VSUBS 0.006783f
C429 B.n389 VSUBS 0.006783f
C430 B.n390 VSUBS 0.006783f
C431 B.n391 VSUBS 0.006783f
C432 B.n392 VSUBS 0.006783f
C433 B.n393 VSUBS 0.006783f
C434 B.n394 VSUBS 0.006783f
C435 B.n395 VSUBS 0.006783f
C436 B.n396 VSUBS 0.006783f
C437 B.n397 VSUBS 0.006783f
C438 B.n398 VSUBS 0.006783f
C439 B.n399 VSUBS 0.006783f
C440 B.n400 VSUBS 0.006783f
C441 B.n401 VSUBS 0.006783f
C442 B.n402 VSUBS 0.006783f
C443 B.n403 VSUBS 0.006783f
C444 B.n404 VSUBS 0.006783f
C445 B.n405 VSUBS 0.006783f
C446 B.n406 VSUBS 0.006783f
C447 B.n407 VSUBS 0.006783f
C448 B.n408 VSUBS 0.006783f
C449 B.n409 VSUBS 0.006783f
C450 B.n410 VSUBS 0.006783f
C451 B.n411 VSUBS 0.006783f
C452 B.n412 VSUBS 0.006783f
C453 B.n413 VSUBS 0.006783f
C454 B.n414 VSUBS 0.006783f
C455 B.n415 VSUBS 0.006783f
C456 B.n416 VSUBS 0.006783f
C457 B.n417 VSUBS 0.006783f
C458 B.n418 VSUBS 0.006783f
C459 B.n419 VSUBS 0.006783f
C460 B.n420 VSUBS 0.006783f
C461 B.n421 VSUBS 0.006783f
C462 B.n422 VSUBS 0.006783f
C463 B.n423 VSUBS 0.015954f
C464 B.n424 VSUBS 0.015168f
C465 B.n425 VSUBS 0.015168f
C466 B.n426 VSUBS 0.006783f
C467 B.n427 VSUBS 0.006783f
C468 B.n428 VSUBS 0.006783f
C469 B.n429 VSUBS 0.006783f
C470 B.n430 VSUBS 0.006783f
C471 B.n431 VSUBS 0.006783f
C472 B.n432 VSUBS 0.006783f
C473 B.n433 VSUBS 0.006783f
C474 B.n434 VSUBS 0.006783f
C475 B.n435 VSUBS 0.006783f
C476 B.n436 VSUBS 0.006783f
C477 B.n437 VSUBS 0.006783f
C478 B.n438 VSUBS 0.006783f
C479 B.n439 VSUBS 0.006783f
C480 B.n440 VSUBS 0.006783f
C481 B.n441 VSUBS 0.006783f
C482 B.n442 VSUBS 0.006783f
C483 B.n443 VSUBS 0.006783f
C484 B.n444 VSUBS 0.006783f
C485 B.n445 VSUBS 0.006783f
C486 B.n446 VSUBS 0.006783f
C487 B.n447 VSUBS 0.006783f
C488 B.n448 VSUBS 0.006783f
C489 B.n449 VSUBS 0.006783f
C490 B.n450 VSUBS 0.006783f
C491 B.n451 VSUBS 0.006783f
C492 B.n452 VSUBS 0.006783f
C493 B.n453 VSUBS 0.006783f
C494 B.n454 VSUBS 0.006783f
C495 B.n455 VSUBS 0.006783f
C496 B.n456 VSUBS 0.006783f
C497 B.n457 VSUBS 0.006783f
C498 B.n458 VSUBS 0.006783f
C499 B.n459 VSUBS 0.006783f
C500 B.n460 VSUBS 0.006783f
C501 B.n461 VSUBS 0.006783f
C502 B.n462 VSUBS 0.006783f
C503 B.n463 VSUBS 0.006783f
C504 B.n464 VSUBS 0.006783f
C505 B.n465 VSUBS 0.006783f
C506 B.n466 VSUBS 0.006783f
C507 B.n467 VSUBS 0.006783f
C508 B.n468 VSUBS 0.006783f
C509 B.n469 VSUBS 0.006783f
C510 B.n470 VSUBS 0.006783f
C511 B.n471 VSUBS 0.006783f
C512 B.n472 VSUBS 0.006783f
C513 B.n473 VSUBS 0.006783f
C514 B.n474 VSUBS 0.006783f
C515 B.n475 VSUBS 0.006783f
C516 B.n476 VSUBS 0.006783f
C517 B.n477 VSUBS 0.006783f
C518 B.n478 VSUBS 0.006783f
C519 B.n479 VSUBS 0.006783f
C520 B.n480 VSUBS 0.006783f
C521 B.n481 VSUBS 0.006783f
C522 B.n482 VSUBS 0.006783f
C523 B.n483 VSUBS 0.006783f
C524 B.n484 VSUBS 0.006783f
C525 B.n485 VSUBS 0.006783f
C526 B.n486 VSUBS 0.006783f
C527 B.n487 VSUBS 0.006783f
C528 B.n488 VSUBS 0.006783f
C529 B.n489 VSUBS 0.006783f
C530 B.n490 VSUBS 0.006783f
C531 B.n491 VSUBS 0.006783f
C532 B.n492 VSUBS 0.006783f
C533 B.n493 VSUBS 0.006783f
C534 B.n494 VSUBS 0.006783f
C535 B.n495 VSUBS 0.006783f
C536 B.n496 VSUBS 0.006783f
C537 B.n497 VSUBS 0.006783f
C538 B.n498 VSUBS 0.006783f
C539 B.n499 VSUBS 0.006783f
C540 B.n500 VSUBS 0.006783f
C541 B.n501 VSUBS 0.006783f
C542 B.n502 VSUBS 0.006783f
C543 B.n503 VSUBS 0.006783f
C544 B.n504 VSUBS 0.006783f
C545 B.n505 VSUBS 0.006783f
C546 B.n506 VSUBS 0.006783f
C547 B.n507 VSUBS 0.006783f
C548 B.n508 VSUBS 0.006783f
C549 B.n509 VSUBS 0.006783f
C550 B.n510 VSUBS 0.006783f
C551 B.n511 VSUBS 0.006783f
C552 B.n512 VSUBS 0.006783f
C553 B.n513 VSUBS 0.006783f
C554 B.n514 VSUBS 0.006783f
C555 B.n515 VSUBS 0.006783f
C556 B.n516 VSUBS 0.006783f
C557 B.n517 VSUBS 0.006783f
C558 B.n518 VSUBS 0.006783f
C559 B.n519 VSUBS 0.006783f
C560 B.n520 VSUBS 0.006783f
C561 B.n521 VSUBS 0.006783f
C562 B.n522 VSUBS 0.006783f
C563 B.n523 VSUBS 0.006783f
C564 B.n524 VSUBS 0.006783f
C565 B.n525 VSUBS 0.006783f
C566 B.n526 VSUBS 0.006783f
C567 B.n527 VSUBS 0.006783f
C568 B.n528 VSUBS 0.006783f
C569 B.n529 VSUBS 0.006783f
C570 B.n530 VSUBS 0.006783f
C571 B.n531 VSUBS 0.006783f
C572 B.n532 VSUBS 0.006783f
C573 B.n533 VSUBS 0.006783f
C574 B.n534 VSUBS 0.006783f
C575 B.n535 VSUBS 0.006783f
C576 B.n536 VSUBS 0.006783f
C577 B.n537 VSUBS 0.006783f
C578 B.n538 VSUBS 0.006783f
C579 B.n539 VSUBS 0.006783f
C580 B.n540 VSUBS 0.006783f
C581 B.n541 VSUBS 0.006783f
C582 B.n542 VSUBS 0.006783f
C583 B.n543 VSUBS 0.006783f
C584 B.n544 VSUBS 0.006783f
C585 B.n545 VSUBS 0.006783f
C586 B.n546 VSUBS 0.006783f
C587 B.n547 VSUBS 0.006783f
C588 B.n548 VSUBS 0.006783f
C589 B.n549 VSUBS 0.006783f
C590 B.n550 VSUBS 0.006783f
C591 B.n551 VSUBS 0.006783f
C592 B.n552 VSUBS 0.006783f
C593 B.n553 VSUBS 0.015994f
C594 B.n554 VSUBS 0.015168f
C595 B.n555 VSUBS 0.015954f
C596 B.n556 VSUBS 0.006783f
C597 B.n557 VSUBS 0.006783f
C598 B.n558 VSUBS 0.006783f
C599 B.n559 VSUBS 0.006783f
C600 B.n560 VSUBS 0.006783f
C601 B.n561 VSUBS 0.006783f
C602 B.n562 VSUBS 0.006783f
C603 B.n563 VSUBS 0.006783f
C604 B.n564 VSUBS 0.006783f
C605 B.n565 VSUBS 0.006783f
C606 B.n566 VSUBS 0.006783f
C607 B.n567 VSUBS 0.006783f
C608 B.n568 VSUBS 0.006783f
C609 B.n569 VSUBS 0.006783f
C610 B.n570 VSUBS 0.006783f
C611 B.n571 VSUBS 0.006783f
C612 B.n572 VSUBS 0.006783f
C613 B.n573 VSUBS 0.006783f
C614 B.n574 VSUBS 0.006783f
C615 B.n575 VSUBS 0.006783f
C616 B.n576 VSUBS 0.006783f
C617 B.n577 VSUBS 0.006783f
C618 B.n578 VSUBS 0.006783f
C619 B.n579 VSUBS 0.006783f
C620 B.n580 VSUBS 0.006783f
C621 B.n581 VSUBS 0.006783f
C622 B.n582 VSUBS 0.006783f
C623 B.n583 VSUBS 0.006783f
C624 B.n584 VSUBS 0.006783f
C625 B.n585 VSUBS 0.006783f
C626 B.n586 VSUBS 0.006783f
C627 B.n587 VSUBS 0.006783f
C628 B.n588 VSUBS 0.006783f
C629 B.n589 VSUBS 0.006783f
C630 B.n590 VSUBS 0.006783f
C631 B.n591 VSUBS 0.006783f
C632 B.n592 VSUBS 0.006783f
C633 B.n593 VSUBS 0.006783f
C634 B.n594 VSUBS 0.006783f
C635 B.n595 VSUBS 0.006783f
C636 B.n596 VSUBS 0.006783f
C637 B.n597 VSUBS 0.006783f
C638 B.n598 VSUBS 0.006783f
C639 B.n599 VSUBS 0.006783f
C640 B.n600 VSUBS 0.006783f
C641 B.n601 VSUBS 0.006783f
C642 B.n602 VSUBS 0.006783f
C643 B.n603 VSUBS 0.006783f
C644 B.n604 VSUBS 0.006783f
C645 B.n605 VSUBS 0.006783f
C646 B.n606 VSUBS 0.006783f
C647 B.n607 VSUBS 0.006783f
C648 B.n608 VSUBS 0.006783f
C649 B.n609 VSUBS 0.006783f
C650 B.n610 VSUBS 0.006783f
C651 B.n611 VSUBS 0.006783f
C652 B.n612 VSUBS 0.006783f
C653 B.n613 VSUBS 0.006783f
C654 B.n614 VSUBS 0.006783f
C655 B.n615 VSUBS 0.006783f
C656 B.n616 VSUBS 0.006783f
C657 B.n617 VSUBS 0.006783f
C658 B.n618 VSUBS 0.006783f
C659 B.n619 VSUBS 0.006783f
C660 B.n620 VSUBS 0.006783f
C661 B.n621 VSUBS 0.006783f
C662 B.n622 VSUBS 0.006783f
C663 B.n623 VSUBS 0.006783f
C664 B.n624 VSUBS 0.006783f
C665 B.n625 VSUBS 0.004688f
C666 B.n626 VSUBS 0.006783f
C667 B.n627 VSUBS 0.006783f
C668 B.n628 VSUBS 0.005486f
C669 B.n629 VSUBS 0.006783f
C670 B.n630 VSUBS 0.006783f
C671 B.n631 VSUBS 0.006783f
C672 B.n632 VSUBS 0.006783f
C673 B.n633 VSUBS 0.006783f
C674 B.n634 VSUBS 0.006783f
C675 B.n635 VSUBS 0.006783f
C676 B.n636 VSUBS 0.006783f
C677 B.n637 VSUBS 0.006783f
C678 B.n638 VSUBS 0.006783f
C679 B.n639 VSUBS 0.006783f
C680 B.n640 VSUBS 0.005486f
C681 B.n641 VSUBS 0.015716f
C682 B.n642 VSUBS 0.004688f
C683 B.n643 VSUBS 0.006783f
C684 B.n644 VSUBS 0.006783f
C685 B.n645 VSUBS 0.006783f
C686 B.n646 VSUBS 0.006783f
C687 B.n647 VSUBS 0.006783f
C688 B.n648 VSUBS 0.006783f
C689 B.n649 VSUBS 0.006783f
C690 B.n650 VSUBS 0.006783f
C691 B.n651 VSUBS 0.006783f
C692 B.n652 VSUBS 0.006783f
C693 B.n653 VSUBS 0.006783f
C694 B.n654 VSUBS 0.006783f
C695 B.n655 VSUBS 0.006783f
C696 B.n656 VSUBS 0.006783f
C697 B.n657 VSUBS 0.006783f
C698 B.n658 VSUBS 0.006783f
C699 B.n659 VSUBS 0.006783f
C700 B.n660 VSUBS 0.006783f
C701 B.n661 VSUBS 0.006783f
C702 B.n662 VSUBS 0.006783f
C703 B.n663 VSUBS 0.006783f
C704 B.n664 VSUBS 0.006783f
C705 B.n665 VSUBS 0.006783f
C706 B.n666 VSUBS 0.006783f
C707 B.n667 VSUBS 0.006783f
C708 B.n668 VSUBS 0.006783f
C709 B.n669 VSUBS 0.006783f
C710 B.n670 VSUBS 0.006783f
C711 B.n671 VSUBS 0.006783f
C712 B.n672 VSUBS 0.006783f
C713 B.n673 VSUBS 0.006783f
C714 B.n674 VSUBS 0.006783f
C715 B.n675 VSUBS 0.006783f
C716 B.n676 VSUBS 0.006783f
C717 B.n677 VSUBS 0.006783f
C718 B.n678 VSUBS 0.006783f
C719 B.n679 VSUBS 0.006783f
C720 B.n680 VSUBS 0.006783f
C721 B.n681 VSUBS 0.006783f
C722 B.n682 VSUBS 0.006783f
C723 B.n683 VSUBS 0.006783f
C724 B.n684 VSUBS 0.006783f
C725 B.n685 VSUBS 0.006783f
C726 B.n686 VSUBS 0.006783f
C727 B.n687 VSUBS 0.006783f
C728 B.n688 VSUBS 0.006783f
C729 B.n689 VSUBS 0.006783f
C730 B.n690 VSUBS 0.006783f
C731 B.n691 VSUBS 0.006783f
C732 B.n692 VSUBS 0.006783f
C733 B.n693 VSUBS 0.006783f
C734 B.n694 VSUBS 0.006783f
C735 B.n695 VSUBS 0.006783f
C736 B.n696 VSUBS 0.006783f
C737 B.n697 VSUBS 0.006783f
C738 B.n698 VSUBS 0.006783f
C739 B.n699 VSUBS 0.006783f
C740 B.n700 VSUBS 0.006783f
C741 B.n701 VSUBS 0.006783f
C742 B.n702 VSUBS 0.006783f
C743 B.n703 VSUBS 0.006783f
C744 B.n704 VSUBS 0.006783f
C745 B.n705 VSUBS 0.006783f
C746 B.n706 VSUBS 0.006783f
C747 B.n707 VSUBS 0.006783f
C748 B.n708 VSUBS 0.006783f
C749 B.n709 VSUBS 0.006783f
C750 B.n710 VSUBS 0.006783f
C751 B.n711 VSUBS 0.006783f
C752 B.n712 VSUBS 0.015954f
C753 B.n713 VSUBS 0.015954f
C754 B.n714 VSUBS 0.015168f
C755 B.n715 VSUBS 0.006783f
C756 B.n716 VSUBS 0.006783f
C757 B.n717 VSUBS 0.006783f
C758 B.n718 VSUBS 0.006783f
C759 B.n719 VSUBS 0.006783f
C760 B.n720 VSUBS 0.006783f
C761 B.n721 VSUBS 0.006783f
C762 B.n722 VSUBS 0.006783f
C763 B.n723 VSUBS 0.006783f
C764 B.n724 VSUBS 0.006783f
C765 B.n725 VSUBS 0.006783f
C766 B.n726 VSUBS 0.006783f
C767 B.n727 VSUBS 0.006783f
C768 B.n728 VSUBS 0.006783f
C769 B.n729 VSUBS 0.006783f
C770 B.n730 VSUBS 0.006783f
C771 B.n731 VSUBS 0.006783f
C772 B.n732 VSUBS 0.006783f
C773 B.n733 VSUBS 0.006783f
C774 B.n734 VSUBS 0.006783f
C775 B.n735 VSUBS 0.006783f
C776 B.n736 VSUBS 0.006783f
C777 B.n737 VSUBS 0.006783f
C778 B.n738 VSUBS 0.006783f
C779 B.n739 VSUBS 0.006783f
C780 B.n740 VSUBS 0.006783f
C781 B.n741 VSUBS 0.006783f
C782 B.n742 VSUBS 0.006783f
C783 B.n743 VSUBS 0.006783f
C784 B.n744 VSUBS 0.006783f
C785 B.n745 VSUBS 0.006783f
C786 B.n746 VSUBS 0.006783f
C787 B.n747 VSUBS 0.006783f
C788 B.n748 VSUBS 0.006783f
C789 B.n749 VSUBS 0.006783f
C790 B.n750 VSUBS 0.006783f
C791 B.n751 VSUBS 0.006783f
C792 B.n752 VSUBS 0.006783f
C793 B.n753 VSUBS 0.006783f
C794 B.n754 VSUBS 0.006783f
C795 B.n755 VSUBS 0.006783f
C796 B.n756 VSUBS 0.006783f
C797 B.n757 VSUBS 0.006783f
C798 B.n758 VSUBS 0.006783f
C799 B.n759 VSUBS 0.006783f
C800 B.n760 VSUBS 0.006783f
C801 B.n761 VSUBS 0.006783f
C802 B.n762 VSUBS 0.006783f
C803 B.n763 VSUBS 0.006783f
C804 B.n764 VSUBS 0.006783f
C805 B.n765 VSUBS 0.006783f
C806 B.n766 VSUBS 0.006783f
C807 B.n767 VSUBS 0.006783f
C808 B.n768 VSUBS 0.006783f
C809 B.n769 VSUBS 0.006783f
C810 B.n770 VSUBS 0.006783f
C811 B.n771 VSUBS 0.006783f
C812 B.n772 VSUBS 0.006783f
C813 B.n773 VSUBS 0.006783f
C814 B.n774 VSUBS 0.006783f
C815 B.n775 VSUBS 0.006783f
C816 B.n776 VSUBS 0.006783f
C817 B.n777 VSUBS 0.006783f
C818 B.n778 VSUBS 0.006783f
C819 B.n779 VSUBS 0.015359f
C820 VDD2.t7 VSUBS 0.272513f
C821 VDD2.t0 VSUBS 0.272513f
C822 VDD2.n0 VSUBS 2.20951f
C823 VDD2.t1 VSUBS 0.272513f
C824 VDD2.t2 VSUBS 0.272513f
C825 VDD2.n1 VSUBS 2.20951f
C826 VDD2.n2 VSUBS 3.52506f
C827 VDD2.t6 VSUBS 0.272513f
C828 VDD2.t5 VSUBS 0.272513f
C829 VDD2.n3 VSUBS 2.20046f
C830 VDD2.n4 VSUBS 3.111f
C831 VDD2.t3 VSUBS 0.272513f
C832 VDD2.t4 VSUBS 0.272513f
C833 VDD2.n5 VSUBS 2.20947f
C834 VN.n0 VSUBS 0.041959f
C835 VN.t5 VSUBS 2.4974f
C836 VN.n1 VSUBS 0.032223f
C837 VN.n2 VSUBS 0.031824f
C838 VN.t6 VSUBS 2.4974f
C839 VN.n3 VSUBS 0.046659f
C840 VN.n4 VSUBS 0.266017f
C841 VN.t7 VSUBS 2.4974f
C842 VN.t0 VSUBS 2.67062f
C843 VN.n5 VSUBS 0.955805f
C844 VN.n6 VSUBS 0.971868f
C845 VN.n7 VSUBS 0.055783f
C846 VN.n8 VSUBS 0.046659f
C847 VN.n9 VSUBS 0.031824f
C848 VN.n10 VSUBS 0.031824f
C849 VN.n11 VSUBS 0.031824f
C850 VN.n12 VSUBS 0.055783f
C851 VN.n13 VSUBS 0.882113f
C852 VN.n14 VSUBS 0.034004f
C853 VN.n15 VSUBS 0.06329f
C854 VN.n16 VSUBS 0.031824f
C855 VN.n17 VSUBS 0.031824f
C856 VN.n18 VSUBS 0.031824f
C857 VN.n19 VSUBS 0.057414f
C858 VN.n20 VSUBS 0.048131f
C859 VN.n21 VSUBS 0.973207f
C860 VN.n22 VSUBS 0.042962f
C861 VN.n23 VSUBS 0.041959f
C862 VN.t1 VSUBS 2.4974f
C863 VN.n24 VSUBS 0.032223f
C864 VN.n25 VSUBS 0.031824f
C865 VN.t2 VSUBS 2.4974f
C866 VN.n26 VSUBS 0.046659f
C867 VN.n27 VSUBS 0.266017f
C868 VN.t4 VSUBS 2.4974f
C869 VN.t3 VSUBS 2.67062f
C870 VN.n28 VSUBS 0.955805f
C871 VN.n29 VSUBS 0.971868f
C872 VN.n30 VSUBS 0.055783f
C873 VN.n31 VSUBS 0.046659f
C874 VN.n32 VSUBS 0.031824f
C875 VN.n33 VSUBS 0.031824f
C876 VN.n34 VSUBS 0.031824f
C877 VN.n35 VSUBS 0.055783f
C878 VN.n36 VSUBS 0.882113f
C879 VN.n37 VSUBS 0.034004f
C880 VN.n38 VSUBS 0.06329f
C881 VN.n39 VSUBS 0.031824f
C882 VN.n40 VSUBS 0.031824f
C883 VN.n41 VSUBS 0.031824f
C884 VN.n42 VSUBS 0.057414f
C885 VN.n43 VSUBS 0.048131f
C886 VN.n44 VSUBS 0.973207f
C887 VN.n45 VSUBS 1.76678f
C888 VTAIL.t3 VSUBS 0.267796f
C889 VTAIL.t2 VSUBS 0.267796f
C890 VTAIL.n0 VSUBS 2.03372f
C891 VTAIL.n1 VSUBS 0.706168f
C892 VTAIL.n2 VSUBS 0.025361f
C893 VTAIL.n3 VSUBS 0.024103f
C894 VTAIL.n4 VSUBS 0.013333f
C895 VTAIL.n5 VSUBS 0.030613f
C896 VTAIL.n6 VSUBS 0.013714f
C897 VTAIL.n7 VSUBS 0.024103f
C898 VTAIL.n8 VSUBS 0.012952f
C899 VTAIL.n9 VSUBS 0.030613f
C900 VTAIL.n10 VSUBS 0.013714f
C901 VTAIL.n11 VSUBS 0.024103f
C902 VTAIL.n12 VSUBS 0.012952f
C903 VTAIL.n13 VSUBS 0.030613f
C904 VTAIL.n14 VSUBS 0.013714f
C905 VTAIL.n15 VSUBS 0.024103f
C906 VTAIL.n16 VSUBS 0.012952f
C907 VTAIL.n17 VSUBS 0.030613f
C908 VTAIL.n18 VSUBS 0.013714f
C909 VTAIL.n19 VSUBS 0.024103f
C910 VTAIL.n20 VSUBS 0.012952f
C911 VTAIL.n21 VSUBS 0.030613f
C912 VTAIL.n22 VSUBS 0.013714f
C913 VTAIL.n23 VSUBS 0.024103f
C914 VTAIL.n24 VSUBS 0.012952f
C915 VTAIL.n25 VSUBS 0.02296f
C916 VTAIL.n26 VSUBS 0.019475f
C917 VTAIL.t4 VSUBS 0.065481f
C918 VTAIL.n27 VSUBS 0.163221f
C919 VTAIL.n28 VSUBS 1.43615f
C920 VTAIL.n29 VSUBS 0.012952f
C921 VTAIL.n30 VSUBS 0.013714f
C922 VTAIL.n31 VSUBS 0.030613f
C923 VTAIL.n32 VSUBS 0.030613f
C924 VTAIL.n33 VSUBS 0.013714f
C925 VTAIL.n34 VSUBS 0.012952f
C926 VTAIL.n35 VSUBS 0.024103f
C927 VTAIL.n36 VSUBS 0.024103f
C928 VTAIL.n37 VSUBS 0.012952f
C929 VTAIL.n38 VSUBS 0.013714f
C930 VTAIL.n39 VSUBS 0.030613f
C931 VTAIL.n40 VSUBS 0.030613f
C932 VTAIL.n41 VSUBS 0.013714f
C933 VTAIL.n42 VSUBS 0.012952f
C934 VTAIL.n43 VSUBS 0.024103f
C935 VTAIL.n44 VSUBS 0.024103f
C936 VTAIL.n45 VSUBS 0.012952f
C937 VTAIL.n46 VSUBS 0.013714f
C938 VTAIL.n47 VSUBS 0.030613f
C939 VTAIL.n48 VSUBS 0.030613f
C940 VTAIL.n49 VSUBS 0.013714f
C941 VTAIL.n50 VSUBS 0.012952f
C942 VTAIL.n51 VSUBS 0.024103f
C943 VTAIL.n52 VSUBS 0.024103f
C944 VTAIL.n53 VSUBS 0.012952f
C945 VTAIL.n54 VSUBS 0.013714f
C946 VTAIL.n55 VSUBS 0.030613f
C947 VTAIL.n56 VSUBS 0.030613f
C948 VTAIL.n57 VSUBS 0.013714f
C949 VTAIL.n58 VSUBS 0.012952f
C950 VTAIL.n59 VSUBS 0.024103f
C951 VTAIL.n60 VSUBS 0.024103f
C952 VTAIL.n61 VSUBS 0.012952f
C953 VTAIL.n62 VSUBS 0.013714f
C954 VTAIL.n63 VSUBS 0.030613f
C955 VTAIL.n64 VSUBS 0.030613f
C956 VTAIL.n65 VSUBS 0.013714f
C957 VTAIL.n66 VSUBS 0.012952f
C958 VTAIL.n67 VSUBS 0.024103f
C959 VTAIL.n68 VSUBS 0.024103f
C960 VTAIL.n69 VSUBS 0.012952f
C961 VTAIL.n70 VSUBS 0.012952f
C962 VTAIL.n71 VSUBS 0.013714f
C963 VTAIL.n72 VSUBS 0.030613f
C964 VTAIL.n73 VSUBS 0.030613f
C965 VTAIL.n74 VSUBS 0.070288f
C966 VTAIL.n75 VSUBS 0.013333f
C967 VTAIL.n76 VSUBS 0.012952f
C968 VTAIL.n77 VSUBS 0.060322f
C969 VTAIL.n78 VSUBS 0.035314f
C970 VTAIL.n79 VSUBS 0.218357f
C971 VTAIL.n80 VSUBS 0.025361f
C972 VTAIL.n81 VSUBS 0.024103f
C973 VTAIL.n82 VSUBS 0.013333f
C974 VTAIL.n83 VSUBS 0.030613f
C975 VTAIL.n84 VSUBS 0.013714f
C976 VTAIL.n85 VSUBS 0.024103f
C977 VTAIL.n86 VSUBS 0.012952f
C978 VTAIL.n87 VSUBS 0.030613f
C979 VTAIL.n88 VSUBS 0.013714f
C980 VTAIL.n89 VSUBS 0.024103f
C981 VTAIL.n90 VSUBS 0.012952f
C982 VTAIL.n91 VSUBS 0.030613f
C983 VTAIL.n92 VSUBS 0.013714f
C984 VTAIL.n93 VSUBS 0.024103f
C985 VTAIL.n94 VSUBS 0.012952f
C986 VTAIL.n95 VSUBS 0.030613f
C987 VTAIL.n96 VSUBS 0.013714f
C988 VTAIL.n97 VSUBS 0.024103f
C989 VTAIL.n98 VSUBS 0.012952f
C990 VTAIL.n99 VSUBS 0.030613f
C991 VTAIL.n100 VSUBS 0.013714f
C992 VTAIL.n101 VSUBS 0.024103f
C993 VTAIL.n102 VSUBS 0.012952f
C994 VTAIL.n103 VSUBS 0.02296f
C995 VTAIL.n104 VSUBS 0.019475f
C996 VTAIL.t10 VSUBS 0.065481f
C997 VTAIL.n105 VSUBS 0.163221f
C998 VTAIL.n106 VSUBS 1.43615f
C999 VTAIL.n107 VSUBS 0.012952f
C1000 VTAIL.n108 VSUBS 0.013714f
C1001 VTAIL.n109 VSUBS 0.030613f
C1002 VTAIL.n110 VSUBS 0.030613f
C1003 VTAIL.n111 VSUBS 0.013714f
C1004 VTAIL.n112 VSUBS 0.012952f
C1005 VTAIL.n113 VSUBS 0.024103f
C1006 VTAIL.n114 VSUBS 0.024103f
C1007 VTAIL.n115 VSUBS 0.012952f
C1008 VTAIL.n116 VSUBS 0.013714f
C1009 VTAIL.n117 VSUBS 0.030613f
C1010 VTAIL.n118 VSUBS 0.030613f
C1011 VTAIL.n119 VSUBS 0.013714f
C1012 VTAIL.n120 VSUBS 0.012952f
C1013 VTAIL.n121 VSUBS 0.024103f
C1014 VTAIL.n122 VSUBS 0.024103f
C1015 VTAIL.n123 VSUBS 0.012952f
C1016 VTAIL.n124 VSUBS 0.013714f
C1017 VTAIL.n125 VSUBS 0.030613f
C1018 VTAIL.n126 VSUBS 0.030613f
C1019 VTAIL.n127 VSUBS 0.013714f
C1020 VTAIL.n128 VSUBS 0.012952f
C1021 VTAIL.n129 VSUBS 0.024103f
C1022 VTAIL.n130 VSUBS 0.024103f
C1023 VTAIL.n131 VSUBS 0.012952f
C1024 VTAIL.n132 VSUBS 0.013714f
C1025 VTAIL.n133 VSUBS 0.030613f
C1026 VTAIL.n134 VSUBS 0.030613f
C1027 VTAIL.n135 VSUBS 0.013714f
C1028 VTAIL.n136 VSUBS 0.012952f
C1029 VTAIL.n137 VSUBS 0.024103f
C1030 VTAIL.n138 VSUBS 0.024103f
C1031 VTAIL.n139 VSUBS 0.012952f
C1032 VTAIL.n140 VSUBS 0.013714f
C1033 VTAIL.n141 VSUBS 0.030613f
C1034 VTAIL.n142 VSUBS 0.030613f
C1035 VTAIL.n143 VSUBS 0.013714f
C1036 VTAIL.n144 VSUBS 0.012952f
C1037 VTAIL.n145 VSUBS 0.024103f
C1038 VTAIL.n146 VSUBS 0.024103f
C1039 VTAIL.n147 VSUBS 0.012952f
C1040 VTAIL.n148 VSUBS 0.012952f
C1041 VTAIL.n149 VSUBS 0.013714f
C1042 VTAIL.n150 VSUBS 0.030613f
C1043 VTAIL.n151 VSUBS 0.030613f
C1044 VTAIL.n152 VSUBS 0.070288f
C1045 VTAIL.n153 VSUBS 0.013333f
C1046 VTAIL.n154 VSUBS 0.012952f
C1047 VTAIL.n155 VSUBS 0.060322f
C1048 VTAIL.n156 VSUBS 0.035314f
C1049 VTAIL.n157 VSUBS 0.218357f
C1050 VTAIL.t8 VSUBS 0.267796f
C1051 VTAIL.t9 VSUBS 0.267796f
C1052 VTAIL.n158 VSUBS 2.03372f
C1053 VTAIL.n159 VSUBS 0.860325f
C1054 VTAIL.n160 VSUBS 0.025361f
C1055 VTAIL.n161 VSUBS 0.024103f
C1056 VTAIL.n162 VSUBS 0.013333f
C1057 VTAIL.n163 VSUBS 0.030613f
C1058 VTAIL.n164 VSUBS 0.013714f
C1059 VTAIL.n165 VSUBS 0.024103f
C1060 VTAIL.n166 VSUBS 0.012952f
C1061 VTAIL.n167 VSUBS 0.030613f
C1062 VTAIL.n168 VSUBS 0.013714f
C1063 VTAIL.n169 VSUBS 0.024103f
C1064 VTAIL.n170 VSUBS 0.012952f
C1065 VTAIL.n171 VSUBS 0.030613f
C1066 VTAIL.n172 VSUBS 0.013714f
C1067 VTAIL.n173 VSUBS 0.024103f
C1068 VTAIL.n174 VSUBS 0.012952f
C1069 VTAIL.n175 VSUBS 0.030613f
C1070 VTAIL.n176 VSUBS 0.013714f
C1071 VTAIL.n177 VSUBS 0.024103f
C1072 VTAIL.n178 VSUBS 0.012952f
C1073 VTAIL.n179 VSUBS 0.030613f
C1074 VTAIL.n180 VSUBS 0.013714f
C1075 VTAIL.n181 VSUBS 0.024103f
C1076 VTAIL.n182 VSUBS 0.012952f
C1077 VTAIL.n183 VSUBS 0.02296f
C1078 VTAIL.n184 VSUBS 0.019475f
C1079 VTAIL.t15 VSUBS 0.065481f
C1080 VTAIL.n185 VSUBS 0.163221f
C1081 VTAIL.n186 VSUBS 1.43615f
C1082 VTAIL.n187 VSUBS 0.012952f
C1083 VTAIL.n188 VSUBS 0.013714f
C1084 VTAIL.n189 VSUBS 0.030613f
C1085 VTAIL.n190 VSUBS 0.030613f
C1086 VTAIL.n191 VSUBS 0.013714f
C1087 VTAIL.n192 VSUBS 0.012952f
C1088 VTAIL.n193 VSUBS 0.024103f
C1089 VTAIL.n194 VSUBS 0.024103f
C1090 VTAIL.n195 VSUBS 0.012952f
C1091 VTAIL.n196 VSUBS 0.013714f
C1092 VTAIL.n197 VSUBS 0.030613f
C1093 VTAIL.n198 VSUBS 0.030613f
C1094 VTAIL.n199 VSUBS 0.013714f
C1095 VTAIL.n200 VSUBS 0.012952f
C1096 VTAIL.n201 VSUBS 0.024103f
C1097 VTAIL.n202 VSUBS 0.024103f
C1098 VTAIL.n203 VSUBS 0.012952f
C1099 VTAIL.n204 VSUBS 0.013714f
C1100 VTAIL.n205 VSUBS 0.030613f
C1101 VTAIL.n206 VSUBS 0.030613f
C1102 VTAIL.n207 VSUBS 0.013714f
C1103 VTAIL.n208 VSUBS 0.012952f
C1104 VTAIL.n209 VSUBS 0.024103f
C1105 VTAIL.n210 VSUBS 0.024103f
C1106 VTAIL.n211 VSUBS 0.012952f
C1107 VTAIL.n212 VSUBS 0.013714f
C1108 VTAIL.n213 VSUBS 0.030613f
C1109 VTAIL.n214 VSUBS 0.030613f
C1110 VTAIL.n215 VSUBS 0.013714f
C1111 VTAIL.n216 VSUBS 0.012952f
C1112 VTAIL.n217 VSUBS 0.024103f
C1113 VTAIL.n218 VSUBS 0.024103f
C1114 VTAIL.n219 VSUBS 0.012952f
C1115 VTAIL.n220 VSUBS 0.013714f
C1116 VTAIL.n221 VSUBS 0.030613f
C1117 VTAIL.n222 VSUBS 0.030613f
C1118 VTAIL.n223 VSUBS 0.013714f
C1119 VTAIL.n224 VSUBS 0.012952f
C1120 VTAIL.n225 VSUBS 0.024103f
C1121 VTAIL.n226 VSUBS 0.024103f
C1122 VTAIL.n227 VSUBS 0.012952f
C1123 VTAIL.n228 VSUBS 0.012952f
C1124 VTAIL.n229 VSUBS 0.013714f
C1125 VTAIL.n230 VSUBS 0.030613f
C1126 VTAIL.n231 VSUBS 0.030613f
C1127 VTAIL.n232 VSUBS 0.070288f
C1128 VTAIL.n233 VSUBS 0.013333f
C1129 VTAIL.n234 VSUBS 0.012952f
C1130 VTAIL.n235 VSUBS 0.060322f
C1131 VTAIL.n236 VSUBS 0.035314f
C1132 VTAIL.n237 VSUBS 1.6093f
C1133 VTAIL.n238 VSUBS 0.025361f
C1134 VTAIL.n239 VSUBS 0.024103f
C1135 VTAIL.n240 VSUBS 0.013333f
C1136 VTAIL.n241 VSUBS 0.030613f
C1137 VTAIL.n242 VSUBS 0.012952f
C1138 VTAIL.n243 VSUBS 0.013714f
C1139 VTAIL.n244 VSUBS 0.024103f
C1140 VTAIL.n245 VSUBS 0.012952f
C1141 VTAIL.n246 VSUBS 0.030613f
C1142 VTAIL.n247 VSUBS 0.013714f
C1143 VTAIL.n248 VSUBS 0.024103f
C1144 VTAIL.n249 VSUBS 0.012952f
C1145 VTAIL.n250 VSUBS 0.030613f
C1146 VTAIL.n251 VSUBS 0.013714f
C1147 VTAIL.n252 VSUBS 0.024103f
C1148 VTAIL.n253 VSUBS 0.012952f
C1149 VTAIL.n254 VSUBS 0.030613f
C1150 VTAIL.n255 VSUBS 0.013714f
C1151 VTAIL.n256 VSUBS 0.024103f
C1152 VTAIL.n257 VSUBS 0.012952f
C1153 VTAIL.n258 VSUBS 0.030613f
C1154 VTAIL.n259 VSUBS 0.013714f
C1155 VTAIL.n260 VSUBS 0.024103f
C1156 VTAIL.n261 VSUBS 0.012952f
C1157 VTAIL.n262 VSUBS 0.02296f
C1158 VTAIL.n263 VSUBS 0.019475f
C1159 VTAIL.t6 VSUBS 0.065481f
C1160 VTAIL.n264 VSUBS 0.163221f
C1161 VTAIL.n265 VSUBS 1.43615f
C1162 VTAIL.n266 VSUBS 0.012952f
C1163 VTAIL.n267 VSUBS 0.013714f
C1164 VTAIL.n268 VSUBS 0.030613f
C1165 VTAIL.n269 VSUBS 0.030613f
C1166 VTAIL.n270 VSUBS 0.013714f
C1167 VTAIL.n271 VSUBS 0.012952f
C1168 VTAIL.n272 VSUBS 0.024103f
C1169 VTAIL.n273 VSUBS 0.024103f
C1170 VTAIL.n274 VSUBS 0.012952f
C1171 VTAIL.n275 VSUBS 0.013714f
C1172 VTAIL.n276 VSUBS 0.030613f
C1173 VTAIL.n277 VSUBS 0.030613f
C1174 VTAIL.n278 VSUBS 0.013714f
C1175 VTAIL.n279 VSUBS 0.012952f
C1176 VTAIL.n280 VSUBS 0.024103f
C1177 VTAIL.n281 VSUBS 0.024103f
C1178 VTAIL.n282 VSUBS 0.012952f
C1179 VTAIL.n283 VSUBS 0.013714f
C1180 VTAIL.n284 VSUBS 0.030613f
C1181 VTAIL.n285 VSUBS 0.030613f
C1182 VTAIL.n286 VSUBS 0.013714f
C1183 VTAIL.n287 VSUBS 0.012952f
C1184 VTAIL.n288 VSUBS 0.024103f
C1185 VTAIL.n289 VSUBS 0.024103f
C1186 VTAIL.n290 VSUBS 0.012952f
C1187 VTAIL.n291 VSUBS 0.013714f
C1188 VTAIL.n292 VSUBS 0.030613f
C1189 VTAIL.n293 VSUBS 0.030613f
C1190 VTAIL.n294 VSUBS 0.013714f
C1191 VTAIL.n295 VSUBS 0.012952f
C1192 VTAIL.n296 VSUBS 0.024103f
C1193 VTAIL.n297 VSUBS 0.024103f
C1194 VTAIL.n298 VSUBS 0.012952f
C1195 VTAIL.n299 VSUBS 0.013714f
C1196 VTAIL.n300 VSUBS 0.030613f
C1197 VTAIL.n301 VSUBS 0.030613f
C1198 VTAIL.n302 VSUBS 0.013714f
C1199 VTAIL.n303 VSUBS 0.012952f
C1200 VTAIL.n304 VSUBS 0.024103f
C1201 VTAIL.n305 VSUBS 0.024103f
C1202 VTAIL.n306 VSUBS 0.012952f
C1203 VTAIL.n307 VSUBS 0.013714f
C1204 VTAIL.n308 VSUBS 0.030613f
C1205 VTAIL.n309 VSUBS 0.030613f
C1206 VTAIL.n310 VSUBS 0.070288f
C1207 VTAIL.n311 VSUBS 0.013333f
C1208 VTAIL.n312 VSUBS 0.012952f
C1209 VTAIL.n313 VSUBS 0.060322f
C1210 VTAIL.n314 VSUBS 0.035314f
C1211 VTAIL.n315 VSUBS 1.6093f
C1212 VTAIL.t0 VSUBS 0.267796f
C1213 VTAIL.t7 VSUBS 0.267796f
C1214 VTAIL.n316 VSUBS 2.03373f
C1215 VTAIL.n317 VSUBS 0.860312f
C1216 VTAIL.n318 VSUBS 0.025361f
C1217 VTAIL.n319 VSUBS 0.024103f
C1218 VTAIL.n320 VSUBS 0.013333f
C1219 VTAIL.n321 VSUBS 0.030613f
C1220 VTAIL.n322 VSUBS 0.012952f
C1221 VTAIL.n323 VSUBS 0.013714f
C1222 VTAIL.n324 VSUBS 0.024103f
C1223 VTAIL.n325 VSUBS 0.012952f
C1224 VTAIL.n326 VSUBS 0.030613f
C1225 VTAIL.n327 VSUBS 0.013714f
C1226 VTAIL.n328 VSUBS 0.024103f
C1227 VTAIL.n329 VSUBS 0.012952f
C1228 VTAIL.n330 VSUBS 0.030613f
C1229 VTAIL.n331 VSUBS 0.013714f
C1230 VTAIL.n332 VSUBS 0.024103f
C1231 VTAIL.n333 VSUBS 0.012952f
C1232 VTAIL.n334 VSUBS 0.030613f
C1233 VTAIL.n335 VSUBS 0.013714f
C1234 VTAIL.n336 VSUBS 0.024103f
C1235 VTAIL.n337 VSUBS 0.012952f
C1236 VTAIL.n338 VSUBS 0.030613f
C1237 VTAIL.n339 VSUBS 0.013714f
C1238 VTAIL.n340 VSUBS 0.024103f
C1239 VTAIL.n341 VSUBS 0.012952f
C1240 VTAIL.n342 VSUBS 0.02296f
C1241 VTAIL.n343 VSUBS 0.019475f
C1242 VTAIL.t5 VSUBS 0.065481f
C1243 VTAIL.n344 VSUBS 0.163221f
C1244 VTAIL.n345 VSUBS 1.43615f
C1245 VTAIL.n346 VSUBS 0.012952f
C1246 VTAIL.n347 VSUBS 0.013714f
C1247 VTAIL.n348 VSUBS 0.030613f
C1248 VTAIL.n349 VSUBS 0.030613f
C1249 VTAIL.n350 VSUBS 0.013714f
C1250 VTAIL.n351 VSUBS 0.012952f
C1251 VTAIL.n352 VSUBS 0.024103f
C1252 VTAIL.n353 VSUBS 0.024103f
C1253 VTAIL.n354 VSUBS 0.012952f
C1254 VTAIL.n355 VSUBS 0.013714f
C1255 VTAIL.n356 VSUBS 0.030613f
C1256 VTAIL.n357 VSUBS 0.030613f
C1257 VTAIL.n358 VSUBS 0.013714f
C1258 VTAIL.n359 VSUBS 0.012952f
C1259 VTAIL.n360 VSUBS 0.024103f
C1260 VTAIL.n361 VSUBS 0.024103f
C1261 VTAIL.n362 VSUBS 0.012952f
C1262 VTAIL.n363 VSUBS 0.013714f
C1263 VTAIL.n364 VSUBS 0.030613f
C1264 VTAIL.n365 VSUBS 0.030613f
C1265 VTAIL.n366 VSUBS 0.013714f
C1266 VTAIL.n367 VSUBS 0.012952f
C1267 VTAIL.n368 VSUBS 0.024103f
C1268 VTAIL.n369 VSUBS 0.024103f
C1269 VTAIL.n370 VSUBS 0.012952f
C1270 VTAIL.n371 VSUBS 0.013714f
C1271 VTAIL.n372 VSUBS 0.030613f
C1272 VTAIL.n373 VSUBS 0.030613f
C1273 VTAIL.n374 VSUBS 0.013714f
C1274 VTAIL.n375 VSUBS 0.012952f
C1275 VTAIL.n376 VSUBS 0.024103f
C1276 VTAIL.n377 VSUBS 0.024103f
C1277 VTAIL.n378 VSUBS 0.012952f
C1278 VTAIL.n379 VSUBS 0.013714f
C1279 VTAIL.n380 VSUBS 0.030613f
C1280 VTAIL.n381 VSUBS 0.030613f
C1281 VTAIL.n382 VSUBS 0.013714f
C1282 VTAIL.n383 VSUBS 0.012952f
C1283 VTAIL.n384 VSUBS 0.024103f
C1284 VTAIL.n385 VSUBS 0.024103f
C1285 VTAIL.n386 VSUBS 0.012952f
C1286 VTAIL.n387 VSUBS 0.013714f
C1287 VTAIL.n388 VSUBS 0.030613f
C1288 VTAIL.n389 VSUBS 0.030613f
C1289 VTAIL.n390 VSUBS 0.070288f
C1290 VTAIL.n391 VSUBS 0.013333f
C1291 VTAIL.n392 VSUBS 0.012952f
C1292 VTAIL.n393 VSUBS 0.060322f
C1293 VTAIL.n394 VSUBS 0.035314f
C1294 VTAIL.n395 VSUBS 0.218357f
C1295 VTAIL.n396 VSUBS 0.025361f
C1296 VTAIL.n397 VSUBS 0.024103f
C1297 VTAIL.n398 VSUBS 0.013333f
C1298 VTAIL.n399 VSUBS 0.030613f
C1299 VTAIL.n400 VSUBS 0.012952f
C1300 VTAIL.n401 VSUBS 0.013714f
C1301 VTAIL.n402 VSUBS 0.024103f
C1302 VTAIL.n403 VSUBS 0.012952f
C1303 VTAIL.n404 VSUBS 0.030613f
C1304 VTAIL.n405 VSUBS 0.013714f
C1305 VTAIL.n406 VSUBS 0.024103f
C1306 VTAIL.n407 VSUBS 0.012952f
C1307 VTAIL.n408 VSUBS 0.030613f
C1308 VTAIL.n409 VSUBS 0.013714f
C1309 VTAIL.n410 VSUBS 0.024103f
C1310 VTAIL.n411 VSUBS 0.012952f
C1311 VTAIL.n412 VSUBS 0.030613f
C1312 VTAIL.n413 VSUBS 0.013714f
C1313 VTAIL.n414 VSUBS 0.024103f
C1314 VTAIL.n415 VSUBS 0.012952f
C1315 VTAIL.n416 VSUBS 0.030613f
C1316 VTAIL.n417 VSUBS 0.013714f
C1317 VTAIL.n418 VSUBS 0.024103f
C1318 VTAIL.n419 VSUBS 0.012952f
C1319 VTAIL.n420 VSUBS 0.02296f
C1320 VTAIL.n421 VSUBS 0.019475f
C1321 VTAIL.t11 VSUBS 0.065481f
C1322 VTAIL.n422 VSUBS 0.163221f
C1323 VTAIL.n423 VSUBS 1.43615f
C1324 VTAIL.n424 VSUBS 0.012952f
C1325 VTAIL.n425 VSUBS 0.013714f
C1326 VTAIL.n426 VSUBS 0.030613f
C1327 VTAIL.n427 VSUBS 0.030613f
C1328 VTAIL.n428 VSUBS 0.013714f
C1329 VTAIL.n429 VSUBS 0.012952f
C1330 VTAIL.n430 VSUBS 0.024103f
C1331 VTAIL.n431 VSUBS 0.024103f
C1332 VTAIL.n432 VSUBS 0.012952f
C1333 VTAIL.n433 VSUBS 0.013714f
C1334 VTAIL.n434 VSUBS 0.030613f
C1335 VTAIL.n435 VSUBS 0.030613f
C1336 VTAIL.n436 VSUBS 0.013714f
C1337 VTAIL.n437 VSUBS 0.012952f
C1338 VTAIL.n438 VSUBS 0.024103f
C1339 VTAIL.n439 VSUBS 0.024103f
C1340 VTAIL.n440 VSUBS 0.012952f
C1341 VTAIL.n441 VSUBS 0.013714f
C1342 VTAIL.n442 VSUBS 0.030613f
C1343 VTAIL.n443 VSUBS 0.030613f
C1344 VTAIL.n444 VSUBS 0.013714f
C1345 VTAIL.n445 VSUBS 0.012952f
C1346 VTAIL.n446 VSUBS 0.024103f
C1347 VTAIL.n447 VSUBS 0.024103f
C1348 VTAIL.n448 VSUBS 0.012952f
C1349 VTAIL.n449 VSUBS 0.013714f
C1350 VTAIL.n450 VSUBS 0.030613f
C1351 VTAIL.n451 VSUBS 0.030613f
C1352 VTAIL.n452 VSUBS 0.013714f
C1353 VTAIL.n453 VSUBS 0.012952f
C1354 VTAIL.n454 VSUBS 0.024103f
C1355 VTAIL.n455 VSUBS 0.024103f
C1356 VTAIL.n456 VSUBS 0.012952f
C1357 VTAIL.n457 VSUBS 0.013714f
C1358 VTAIL.n458 VSUBS 0.030613f
C1359 VTAIL.n459 VSUBS 0.030613f
C1360 VTAIL.n460 VSUBS 0.013714f
C1361 VTAIL.n461 VSUBS 0.012952f
C1362 VTAIL.n462 VSUBS 0.024103f
C1363 VTAIL.n463 VSUBS 0.024103f
C1364 VTAIL.n464 VSUBS 0.012952f
C1365 VTAIL.n465 VSUBS 0.013714f
C1366 VTAIL.n466 VSUBS 0.030613f
C1367 VTAIL.n467 VSUBS 0.030613f
C1368 VTAIL.n468 VSUBS 0.070288f
C1369 VTAIL.n469 VSUBS 0.013333f
C1370 VTAIL.n470 VSUBS 0.012952f
C1371 VTAIL.n471 VSUBS 0.060322f
C1372 VTAIL.n472 VSUBS 0.035314f
C1373 VTAIL.n473 VSUBS 0.218357f
C1374 VTAIL.t12 VSUBS 0.267796f
C1375 VTAIL.t13 VSUBS 0.267796f
C1376 VTAIL.n474 VSUBS 2.03373f
C1377 VTAIL.n475 VSUBS 0.860312f
C1378 VTAIL.n476 VSUBS 0.025361f
C1379 VTAIL.n477 VSUBS 0.024103f
C1380 VTAIL.n478 VSUBS 0.013333f
C1381 VTAIL.n479 VSUBS 0.030613f
C1382 VTAIL.n480 VSUBS 0.012952f
C1383 VTAIL.n481 VSUBS 0.013714f
C1384 VTAIL.n482 VSUBS 0.024103f
C1385 VTAIL.n483 VSUBS 0.012952f
C1386 VTAIL.n484 VSUBS 0.030613f
C1387 VTAIL.n485 VSUBS 0.013714f
C1388 VTAIL.n486 VSUBS 0.024103f
C1389 VTAIL.n487 VSUBS 0.012952f
C1390 VTAIL.n488 VSUBS 0.030613f
C1391 VTAIL.n489 VSUBS 0.013714f
C1392 VTAIL.n490 VSUBS 0.024103f
C1393 VTAIL.n491 VSUBS 0.012952f
C1394 VTAIL.n492 VSUBS 0.030613f
C1395 VTAIL.n493 VSUBS 0.013714f
C1396 VTAIL.n494 VSUBS 0.024103f
C1397 VTAIL.n495 VSUBS 0.012952f
C1398 VTAIL.n496 VSUBS 0.030613f
C1399 VTAIL.n497 VSUBS 0.013714f
C1400 VTAIL.n498 VSUBS 0.024103f
C1401 VTAIL.n499 VSUBS 0.012952f
C1402 VTAIL.n500 VSUBS 0.02296f
C1403 VTAIL.n501 VSUBS 0.019475f
C1404 VTAIL.t14 VSUBS 0.065481f
C1405 VTAIL.n502 VSUBS 0.163221f
C1406 VTAIL.n503 VSUBS 1.43615f
C1407 VTAIL.n504 VSUBS 0.012952f
C1408 VTAIL.n505 VSUBS 0.013714f
C1409 VTAIL.n506 VSUBS 0.030613f
C1410 VTAIL.n507 VSUBS 0.030613f
C1411 VTAIL.n508 VSUBS 0.013714f
C1412 VTAIL.n509 VSUBS 0.012952f
C1413 VTAIL.n510 VSUBS 0.024103f
C1414 VTAIL.n511 VSUBS 0.024103f
C1415 VTAIL.n512 VSUBS 0.012952f
C1416 VTAIL.n513 VSUBS 0.013714f
C1417 VTAIL.n514 VSUBS 0.030613f
C1418 VTAIL.n515 VSUBS 0.030613f
C1419 VTAIL.n516 VSUBS 0.013714f
C1420 VTAIL.n517 VSUBS 0.012952f
C1421 VTAIL.n518 VSUBS 0.024103f
C1422 VTAIL.n519 VSUBS 0.024103f
C1423 VTAIL.n520 VSUBS 0.012952f
C1424 VTAIL.n521 VSUBS 0.013714f
C1425 VTAIL.n522 VSUBS 0.030613f
C1426 VTAIL.n523 VSUBS 0.030613f
C1427 VTAIL.n524 VSUBS 0.013714f
C1428 VTAIL.n525 VSUBS 0.012952f
C1429 VTAIL.n526 VSUBS 0.024103f
C1430 VTAIL.n527 VSUBS 0.024103f
C1431 VTAIL.n528 VSUBS 0.012952f
C1432 VTAIL.n529 VSUBS 0.013714f
C1433 VTAIL.n530 VSUBS 0.030613f
C1434 VTAIL.n531 VSUBS 0.030613f
C1435 VTAIL.n532 VSUBS 0.013714f
C1436 VTAIL.n533 VSUBS 0.012952f
C1437 VTAIL.n534 VSUBS 0.024103f
C1438 VTAIL.n535 VSUBS 0.024103f
C1439 VTAIL.n536 VSUBS 0.012952f
C1440 VTAIL.n537 VSUBS 0.013714f
C1441 VTAIL.n538 VSUBS 0.030613f
C1442 VTAIL.n539 VSUBS 0.030613f
C1443 VTAIL.n540 VSUBS 0.013714f
C1444 VTAIL.n541 VSUBS 0.012952f
C1445 VTAIL.n542 VSUBS 0.024103f
C1446 VTAIL.n543 VSUBS 0.024103f
C1447 VTAIL.n544 VSUBS 0.012952f
C1448 VTAIL.n545 VSUBS 0.013714f
C1449 VTAIL.n546 VSUBS 0.030613f
C1450 VTAIL.n547 VSUBS 0.030613f
C1451 VTAIL.n548 VSUBS 0.070288f
C1452 VTAIL.n549 VSUBS 0.013333f
C1453 VTAIL.n550 VSUBS 0.012952f
C1454 VTAIL.n551 VSUBS 0.060322f
C1455 VTAIL.n552 VSUBS 0.035314f
C1456 VTAIL.n553 VSUBS 1.6093f
C1457 VTAIL.n554 VSUBS 0.025361f
C1458 VTAIL.n555 VSUBS 0.024103f
C1459 VTAIL.n556 VSUBS 0.013333f
C1460 VTAIL.n557 VSUBS 0.030613f
C1461 VTAIL.n558 VSUBS 0.013714f
C1462 VTAIL.n559 VSUBS 0.024103f
C1463 VTAIL.n560 VSUBS 0.012952f
C1464 VTAIL.n561 VSUBS 0.030613f
C1465 VTAIL.n562 VSUBS 0.013714f
C1466 VTAIL.n563 VSUBS 0.024103f
C1467 VTAIL.n564 VSUBS 0.012952f
C1468 VTAIL.n565 VSUBS 0.030613f
C1469 VTAIL.n566 VSUBS 0.013714f
C1470 VTAIL.n567 VSUBS 0.024103f
C1471 VTAIL.n568 VSUBS 0.012952f
C1472 VTAIL.n569 VSUBS 0.030613f
C1473 VTAIL.n570 VSUBS 0.013714f
C1474 VTAIL.n571 VSUBS 0.024103f
C1475 VTAIL.n572 VSUBS 0.012952f
C1476 VTAIL.n573 VSUBS 0.030613f
C1477 VTAIL.n574 VSUBS 0.013714f
C1478 VTAIL.n575 VSUBS 0.024103f
C1479 VTAIL.n576 VSUBS 0.012952f
C1480 VTAIL.n577 VSUBS 0.02296f
C1481 VTAIL.n578 VSUBS 0.019475f
C1482 VTAIL.t1 VSUBS 0.065481f
C1483 VTAIL.n579 VSUBS 0.163221f
C1484 VTAIL.n580 VSUBS 1.43615f
C1485 VTAIL.n581 VSUBS 0.012952f
C1486 VTAIL.n582 VSUBS 0.013714f
C1487 VTAIL.n583 VSUBS 0.030613f
C1488 VTAIL.n584 VSUBS 0.030613f
C1489 VTAIL.n585 VSUBS 0.013714f
C1490 VTAIL.n586 VSUBS 0.012952f
C1491 VTAIL.n587 VSUBS 0.024103f
C1492 VTAIL.n588 VSUBS 0.024103f
C1493 VTAIL.n589 VSUBS 0.012952f
C1494 VTAIL.n590 VSUBS 0.013714f
C1495 VTAIL.n591 VSUBS 0.030613f
C1496 VTAIL.n592 VSUBS 0.030613f
C1497 VTAIL.n593 VSUBS 0.013714f
C1498 VTAIL.n594 VSUBS 0.012952f
C1499 VTAIL.n595 VSUBS 0.024103f
C1500 VTAIL.n596 VSUBS 0.024103f
C1501 VTAIL.n597 VSUBS 0.012952f
C1502 VTAIL.n598 VSUBS 0.013714f
C1503 VTAIL.n599 VSUBS 0.030613f
C1504 VTAIL.n600 VSUBS 0.030613f
C1505 VTAIL.n601 VSUBS 0.013714f
C1506 VTAIL.n602 VSUBS 0.012952f
C1507 VTAIL.n603 VSUBS 0.024103f
C1508 VTAIL.n604 VSUBS 0.024103f
C1509 VTAIL.n605 VSUBS 0.012952f
C1510 VTAIL.n606 VSUBS 0.013714f
C1511 VTAIL.n607 VSUBS 0.030613f
C1512 VTAIL.n608 VSUBS 0.030613f
C1513 VTAIL.n609 VSUBS 0.013714f
C1514 VTAIL.n610 VSUBS 0.012952f
C1515 VTAIL.n611 VSUBS 0.024103f
C1516 VTAIL.n612 VSUBS 0.024103f
C1517 VTAIL.n613 VSUBS 0.012952f
C1518 VTAIL.n614 VSUBS 0.013714f
C1519 VTAIL.n615 VSUBS 0.030613f
C1520 VTAIL.n616 VSUBS 0.030613f
C1521 VTAIL.n617 VSUBS 0.013714f
C1522 VTAIL.n618 VSUBS 0.012952f
C1523 VTAIL.n619 VSUBS 0.024103f
C1524 VTAIL.n620 VSUBS 0.024103f
C1525 VTAIL.n621 VSUBS 0.012952f
C1526 VTAIL.n622 VSUBS 0.012952f
C1527 VTAIL.n623 VSUBS 0.013714f
C1528 VTAIL.n624 VSUBS 0.030613f
C1529 VTAIL.n625 VSUBS 0.030613f
C1530 VTAIL.n626 VSUBS 0.070288f
C1531 VTAIL.n627 VSUBS 0.013333f
C1532 VTAIL.n628 VSUBS 0.012952f
C1533 VTAIL.n629 VSUBS 0.060322f
C1534 VTAIL.n630 VSUBS 0.035314f
C1535 VTAIL.n631 VSUBS 1.60478f
C1536 VDD1.t6 VSUBS 0.275582f
C1537 VDD1.t7 VSUBS 0.275582f
C1538 VDD1.n0 VSUBS 2.23559f
C1539 VDD1.t3 VSUBS 0.275582f
C1540 VDD1.t5 VSUBS 0.275582f
C1541 VDD1.n1 VSUBS 2.2344f
C1542 VDD1.t4 VSUBS 0.275582f
C1543 VDD1.t2 VSUBS 0.275582f
C1544 VDD1.n2 VSUBS 2.2344f
C1545 VDD1.n3 VSUBS 3.61667f
C1546 VDD1.t0 VSUBS 0.275582f
C1547 VDD1.t1 VSUBS 0.275582f
C1548 VDD1.n4 VSUBS 2.22524f
C1549 VDD1.n5 VSUBS 3.17646f
C1550 VP.n0 VSUBS 0.042896f
C1551 VP.t5 VSUBS 2.55316f
C1552 VP.n1 VSUBS 0.032942f
C1553 VP.n2 VSUBS 0.032534f
C1554 VP.t6 VSUBS 2.55316f
C1555 VP.n3 VSUBS 0.047701f
C1556 VP.n4 VSUBS 0.032534f
C1557 VP.t7 VSUBS 2.55316f
C1558 VP.n5 VSUBS 0.064703f
C1559 VP.n6 VSUBS 0.032534f
C1560 VP.t0 VSUBS 2.55316f
C1561 VP.n7 VSUBS 0.994936f
C1562 VP.n8 VSUBS 0.042896f
C1563 VP.t1 VSUBS 2.55316f
C1564 VP.n9 VSUBS 0.032942f
C1565 VP.n10 VSUBS 0.032534f
C1566 VP.t2 VSUBS 2.55316f
C1567 VP.n11 VSUBS 0.047701f
C1568 VP.n12 VSUBS 0.271957f
C1569 VP.t3 VSUBS 2.55316f
C1570 VP.t4 VSUBS 2.73025f
C1571 VP.n13 VSUBS 0.977146f
C1572 VP.n14 VSUBS 0.993568f
C1573 VP.n15 VSUBS 0.057028f
C1574 VP.n16 VSUBS 0.047701f
C1575 VP.n17 VSUBS 0.032534f
C1576 VP.n18 VSUBS 0.032534f
C1577 VP.n19 VSUBS 0.032534f
C1578 VP.n20 VSUBS 0.057028f
C1579 VP.n21 VSUBS 0.901808f
C1580 VP.n22 VSUBS 0.034763f
C1581 VP.n23 VSUBS 0.064703f
C1582 VP.n24 VSUBS 0.032534f
C1583 VP.n25 VSUBS 0.032534f
C1584 VP.n26 VSUBS 0.032534f
C1585 VP.n27 VSUBS 0.058696f
C1586 VP.n28 VSUBS 0.049205f
C1587 VP.n29 VSUBS 0.994936f
C1588 VP.n30 VSUBS 1.78873f
C1589 VP.n31 VSUBS 1.81215f
C1590 VP.n32 VSUBS 0.042896f
C1591 VP.n33 VSUBS 0.049205f
C1592 VP.n34 VSUBS 0.058696f
C1593 VP.n35 VSUBS 0.032942f
C1594 VP.n36 VSUBS 0.032534f
C1595 VP.n37 VSUBS 0.032534f
C1596 VP.n38 VSUBS 0.032534f
C1597 VP.n39 VSUBS 0.034763f
C1598 VP.n40 VSUBS 0.901808f
C1599 VP.n41 VSUBS 0.057028f
C1600 VP.n42 VSUBS 0.047701f
C1601 VP.n43 VSUBS 0.032534f
C1602 VP.n44 VSUBS 0.032534f
C1603 VP.n45 VSUBS 0.032534f
C1604 VP.n46 VSUBS 0.057028f
C1605 VP.n47 VSUBS 0.901808f
C1606 VP.n48 VSUBS 0.034763f
C1607 VP.n49 VSUBS 0.064703f
C1608 VP.n50 VSUBS 0.032534f
C1609 VP.n51 VSUBS 0.032534f
C1610 VP.n52 VSUBS 0.032534f
C1611 VP.n53 VSUBS 0.058696f
C1612 VP.n54 VSUBS 0.049205f
C1613 VP.n55 VSUBS 0.994936f
C1614 VP.n56 VSUBS 0.043921f
.ends

