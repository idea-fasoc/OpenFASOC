* NGSPICE file created from diff_pair_sample_0843.ext - technology: sky130A

.subckt diff_pair_sample_0843 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=1.53
X1 VTAIL.t9 VN.t1 VDD2.t4 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=1.61205 ps=10.1 w=9.77 l=1.53
X2 VDD1.t5 VP.t0 VTAIL.t0 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=1.53
X3 VDD2.t3 VN.t2 VTAIL.t6 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=1.53
X4 VDD1.t4 VP.t1 VTAIL.t2 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=1.53
X5 VDD2.t2 VN.t3 VTAIL.t8 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=1.53
X6 VTAIL.t7 VN.t4 VDD2.t1 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=1.61205 ps=10.1 w=9.77 l=1.53
X7 VTAIL.t3 VP.t2 VDD1.t3 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=1.61205 ps=10.1 w=9.77 l=1.53
X8 VDD2.t0 VN.t5 VTAIL.t11 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=1.53
X9 B.t11 B.t9 B.t10 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=1.53
X10 VDD1.t2 VP.t3 VTAIL.t5 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=1.53
X11 B.t8 B.t6 B.t7 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=1.53
X12 B.t5 B.t3 B.t4 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=1.53
X13 VTAIL.t1 VP.t4 VDD1.t1 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=1.61205 ps=10.1 w=9.77 l=1.53
X14 B.t2 B.t0 B.t1 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=1.53
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n2458_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=1.53
R0 VN.n2 VN.t3 185.137
R1 VN.n14 VN.t5 185.137
R2 VN.n11 VN.n10 180.385
R3 VN.n23 VN.n22 180.385
R4 VN.n21 VN.n12 161.3
R5 VN.n20 VN.n19 161.3
R6 VN.n18 VN.n13 161.3
R7 VN.n17 VN.n16 161.3
R8 VN.n9 VN.n0 161.3
R9 VN.n8 VN.n7 161.3
R10 VN.n6 VN.n1 161.3
R11 VN.n5 VN.n4 161.3
R12 VN.n3 VN.t1 153.893
R13 VN.n10 VN.t2 153.893
R14 VN.n15 VN.t4 153.893
R15 VN.n22 VN.t0 153.893
R16 VN.n8 VN.n1 56.5193
R17 VN.n20 VN.n13 56.5193
R18 VN.n3 VN.n2 53.6827
R19 VN.n15 VN.n14 53.6827
R20 VN VN.n23 43.0327
R21 VN.n4 VN.n1 24.4675
R22 VN.n9 VN.n8 24.4675
R23 VN.n16 VN.n13 24.4675
R24 VN.n21 VN.n20 24.4675
R25 VN.n17 VN.n14 18.2406
R26 VN.n5 VN.n2 18.2406
R27 VN.n4 VN.n3 12.234
R28 VN.n16 VN.n15 12.234
R29 VN.n10 VN.n9 5.38324
R30 VN.n22 VN.n21 5.38324
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n7 VTAIL.t11 67.7655
R41 VTAIL.n11 VTAIL.t6 67.7654
R42 VTAIL.n2 VTAIL.t0 67.7654
R43 VTAIL.n10 VTAIL.t4 67.7654
R44 VTAIL.n9 VTAIL.n8 64.4386
R45 VTAIL.n6 VTAIL.n5 64.4386
R46 VTAIL.n1 VTAIL.n0 64.4383
R47 VTAIL.n4 VTAIL.n3 64.4383
R48 VTAIL.n6 VTAIL.n4 23.9962
R49 VTAIL.n11 VTAIL.n10 22.3927
R50 VTAIL.n0 VTAIL.t8 3.32752
R51 VTAIL.n0 VTAIL.t9 3.32752
R52 VTAIL.n3 VTAIL.t2 3.32752
R53 VTAIL.n3 VTAIL.t1 3.32752
R54 VTAIL.n8 VTAIL.t5 3.32752
R55 VTAIL.n8 VTAIL.t3 3.32752
R56 VTAIL.n5 VTAIL.t10 3.32752
R57 VTAIL.n5 VTAIL.t7 3.32752
R58 VTAIL.n7 VTAIL.n6 1.60395
R59 VTAIL.n10 VTAIL.n9 1.60395
R60 VTAIL.n4 VTAIL.n2 1.60395
R61 VTAIL.n9 VTAIL.n7 1.27205
R62 VTAIL.n2 VTAIL.n1 1.27205
R63 VTAIL VTAIL.n11 1.1449
R64 VTAIL VTAIL.n1 0.459552
R65 VDD2.n1 VDD2.t2 85.5914
R66 VDD2.n2 VDD2.t5 84.4443
R67 VDD2.n1 VDD2.n0 81.4626
R68 VDD2 VDD2.n3 81.4598
R69 VDD2.n2 VDD2.n1 37.3489
R70 VDD2.n3 VDD2.t1 3.32752
R71 VDD2.n3 VDD2.t0 3.32752
R72 VDD2.n0 VDD2.t4 3.32752
R73 VDD2.n0 VDD2.t3 3.32752
R74 VDD2 VDD2.n2 1.26128
R75 VP.n6 VP.t3 185.137
R76 VP.n17 VP.n16 180.385
R77 VP.n32 VP.n31 180.385
R78 VP.n15 VP.n14 180.385
R79 VP.n9 VP.n8 161.3
R80 VP.n10 VP.n5 161.3
R81 VP.n12 VP.n11 161.3
R82 VP.n13 VP.n4 161.3
R83 VP.n30 VP.n0 161.3
R84 VP.n29 VP.n28 161.3
R85 VP.n27 VP.n1 161.3
R86 VP.n26 VP.n25 161.3
R87 VP.n23 VP.n2 161.3
R88 VP.n22 VP.n21 161.3
R89 VP.n20 VP.n3 161.3
R90 VP.n19 VP.n18 161.3
R91 VP.n17 VP.t1 153.893
R92 VP.n24 VP.t4 153.893
R93 VP.n31 VP.t0 153.893
R94 VP.n14 VP.t5 153.893
R95 VP.n7 VP.t2 153.893
R96 VP.n29 VP.n1 56.5193
R97 VP.n22 VP.n3 56.5193
R98 VP.n12 VP.n5 56.5193
R99 VP.n7 VP.n6 53.6827
R100 VP.n16 VP.n15 42.652
R101 VP.n18 VP.n3 24.4675
R102 VP.n23 VP.n22 24.4675
R103 VP.n25 VP.n1 24.4675
R104 VP.n30 VP.n29 24.4675
R105 VP.n13 VP.n12 24.4675
R106 VP.n8 VP.n5 24.4675
R107 VP.n9 VP.n6 18.2406
R108 VP.n24 VP.n23 12.234
R109 VP.n25 VP.n24 12.234
R110 VP.n8 VP.n7 12.234
R111 VP.n18 VP.n17 5.38324
R112 VP.n31 VP.n30 5.38324
R113 VP.n14 VP.n13 5.38324
R114 VP.n10 VP.n9 0.189894
R115 VP.n11 VP.n10 0.189894
R116 VP.n11 VP.n4 0.189894
R117 VP.n15 VP.n4 0.189894
R118 VP.n19 VP.n16 0.189894
R119 VP.n20 VP.n19 0.189894
R120 VP.n21 VP.n20 0.189894
R121 VP.n21 VP.n2 0.189894
R122 VP.n26 VP.n2 0.189894
R123 VP.n27 VP.n26 0.189894
R124 VP.n28 VP.n27 0.189894
R125 VP.n28 VP.n0 0.189894
R126 VP.n32 VP.n0 0.189894
R127 VP VP.n32 0.0516364
R128 VDD1 VDD1.t2 85.7051
R129 VDD1.n1 VDD1.t4 85.5914
R130 VDD1.n1 VDD1.n0 81.4626
R131 VDD1.n3 VDD1.n2 81.1172
R132 VDD1.n3 VDD1.n1 38.7337
R133 VDD1.n2 VDD1.t3 3.32752
R134 VDD1.n2 VDD1.t0 3.32752
R135 VDD1.n0 VDD1.t1 3.32752
R136 VDD1.n0 VDD1.t5 3.32752
R137 VDD1 VDD1.n3 0.343172
R138 B.n409 B.n408 585
R139 B.n410 B.n61 585
R140 B.n412 B.n411 585
R141 B.n413 B.n60 585
R142 B.n415 B.n414 585
R143 B.n416 B.n59 585
R144 B.n418 B.n417 585
R145 B.n419 B.n58 585
R146 B.n421 B.n420 585
R147 B.n422 B.n57 585
R148 B.n424 B.n423 585
R149 B.n425 B.n56 585
R150 B.n427 B.n426 585
R151 B.n428 B.n55 585
R152 B.n430 B.n429 585
R153 B.n431 B.n54 585
R154 B.n433 B.n432 585
R155 B.n434 B.n53 585
R156 B.n436 B.n435 585
R157 B.n437 B.n52 585
R158 B.n439 B.n438 585
R159 B.n440 B.n51 585
R160 B.n442 B.n441 585
R161 B.n443 B.n50 585
R162 B.n445 B.n444 585
R163 B.n446 B.n49 585
R164 B.n448 B.n447 585
R165 B.n449 B.n48 585
R166 B.n451 B.n450 585
R167 B.n452 B.n47 585
R168 B.n454 B.n453 585
R169 B.n455 B.n46 585
R170 B.n457 B.n456 585
R171 B.n458 B.n45 585
R172 B.n460 B.n459 585
R173 B.n462 B.n42 585
R174 B.n464 B.n463 585
R175 B.n465 B.n41 585
R176 B.n467 B.n466 585
R177 B.n468 B.n40 585
R178 B.n470 B.n469 585
R179 B.n471 B.n39 585
R180 B.n473 B.n472 585
R181 B.n474 B.n35 585
R182 B.n476 B.n475 585
R183 B.n477 B.n34 585
R184 B.n479 B.n478 585
R185 B.n480 B.n33 585
R186 B.n482 B.n481 585
R187 B.n483 B.n32 585
R188 B.n485 B.n484 585
R189 B.n486 B.n31 585
R190 B.n488 B.n487 585
R191 B.n489 B.n30 585
R192 B.n491 B.n490 585
R193 B.n492 B.n29 585
R194 B.n494 B.n493 585
R195 B.n495 B.n28 585
R196 B.n497 B.n496 585
R197 B.n498 B.n27 585
R198 B.n500 B.n499 585
R199 B.n501 B.n26 585
R200 B.n503 B.n502 585
R201 B.n504 B.n25 585
R202 B.n506 B.n505 585
R203 B.n507 B.n24 585
R204 B.n509 B.n508 585
R205 B.n510 B.n23 585
R206 B.n512 B.n511 585
R207 B.n513 B.n22 585
R208 B.n515 B.n514 585
R209 B.n516 B.n21 585
R210 B.n518 B.n517 585
R211 B.n519 B.n20 585
R212 B.n521 B.n520 585
R213 B.n522 B.n19 585
R214 B.n524 B.n523 585
R215 B.n525 B.n18 585
R216 B.n527 B.n526 585
R217 B.n528 B.n17 585
R218 B.n407 B.n62 585
R219 B.n406 B.n405 585
R220 B.n404 B.n63 585
R221 B.n403 B.n402 585
R222 B.n401 B.n64 585
R223 B.n400 B.n399 585
R224 B.n398 B.n65 585
R225 B.n397 B.n396 585
R226 B.n395 B.n66 585
R227 B.n394 B.n393 585
R228 B.n392 B.n67 585
R229 B.n391 B.n390 585
R230 B.n389 B.n68 585
R231 B.n388 B.n387 585
R232 B.n386 B.n69 585
R233 B.n385 B.n384 585
R234 B.n383 B.n70 585
R235 B.n382 B.n381 585
R236 B.n380 B.n71 585
R237 B.n379 B.n378 585
R238 B.n377 B.n72 585
R239 B.n376 B.n375 585
R240 B.n374 B.n73 585
R241 B.n373 B.n372 585
R242 B.n371 B.n74 585
R243 B.n370 B.n369 585
R244 B.n368 B.n75 585
R245 B.n367 B.n366 585
R246 B.n365 B.n76 585
R247 B.n364 B.n363 585
R248 B.n362 B.n77 585
R249 B.n361 B.n360 585
R250 B.n359 B.n78 585
R251 B.n358 B.n357 585
R252 B.n356 B.n79 585
R253 B.n355 B.n354 585
R254 B.n353 B.n80 585
R255 B.n352 B.n351 585
R256 B.n350 B.n81 585
R257 B.n349 B.n348 585
R258 B.n347 B.n82 585
R259 B.n346 B.n345 585
R260 B.n344 B.n83 585
R261 B.n343 B.n342 585
R262 B.n341 B.n84 585
R263 B.n340 B.n339 585
R264 B.n338 B.n85 585
R265 B.n337 B.n336 585
R266 B.n335 B.n86 585
R267 B.n334 B.n333 585
R268 B.n332 B.n87 585
R269 B.n331 B.n330 585
R270 B.n329 B.n88 585
R271 B.n328 B.n327 585
R272 B.n326 B.n89 585
R273 B.n325 B.n324 585
R274 B.n323 B.n90 585
R275 B.n322 B.n321 585
R276 B.n320 B.n91 585
R277 B.n319 B.n318 585
R278 B.n317 B.n92 585
R279 B.n196 B.n195 585
R280 B.n197 B.n136 585
R281 B.n199 B.n198 585
R282 B.n200 B.n135 585
R283 B.n202 B.n201 585
R284 B.n203 B.n134 585
R285 B.n205 B.n204 585
R286 B.n206 B.n133 585
R287 B.n208 B.n207 585
R288 B.n209 B.n132 585
R289 B.n211 B.n210 585
R290 B.n212 B.n131 585
R291 B.n214 B.n213 585
R292 B.n215 B.n130 585
R293 B.n217 B.n216 585
R294 B.n218 B.n129 585
R295 B.n220 B.n219 585
R296 B.n221 B.n128 585
R297 B.n223 B.n222 585
R298 B.n224 B.n127 585
R299 B.n226 B.n225 585
R300 B.n227 B.n126 585
R301 B.n229 B.n228 585
R302 B.n230 B.n125 585
R303 B.n232 B.n231 585
R304 B.n233 B.n124 585
R305 B.n235 B.n234 585
R306 B.n236 B.n123 585
R307 B.n238 B.n237 585
R308 B.n239 B.n122 585
R309 B.n241 B.n240 585
R310 B.n242 B.n121 585
R311 B.n244 B.n243 585
R312 B.n245 B.n120 585
R313 B.n247 B.n246 585
R314 B.n249 B.n248 585
R315 B.n250 B.n116 585
R316 B.n252 B.n251 585
R317 B.n253 B.n115 585
R318 B.n255 B.n254 585
R319 B.n256 B.n114 585
R320 B.n258 B.n257 585
R321 B.n259 B.n113 585
R322 B.n261 B.n260 585
R323 B.n262 B.n110 585
R324 B.n265 B.n264 585
R325 B.n266 B.n109 585
R326 B.n268 B.n267 585
R327 B.n269 B.n108 585
R328 B.n271 B.n270 585
R329 B.n272 B.n107 585
R330 B.n274 B.n273 585
R331 B.n275 B.n106 585
R332 B.n277 B.n276 585
R333 B.n278 B.n105 585
R334 B.n280 B.n279 585
R335 B.n281 B.n104 585
R336 B.n283 B.n282 585
R337 B.n284 B.n103 585
R338 B.n286 B.n285 585
R339 B.n287 B.n102 585
R340 B.n289 B.n288 585
R341 B.n290 B.n101 585
R342 B.n292 B.n291 585
R343 B.n293 B.n100 585
R344 B.n295 B.n294 585
R345 B.n296 B.n99 585
R346 B.n298 B.n297 585
R347 B.n299 B.n98 585
R348 B.n301 B.n300 585
R349 B.n302 B.n97 585
R350 B.n304 B.n303 585
R351 B.n305 B.n96 585
R352 B.n307 B.n306 585
R353 B.n308 B.n95 585
R354 B.n310 B.n309 585
R355 B.n311 B.n94 585
R356 B.n313 B.n312 585
R357 B.n314 B.n93 585
R358 B.n316 B.n315 585
R359 B.n194 B.n137 585
R360 B.n193 B.n192 585
R361 B.n191 B.n138 585
R362 B.n190 B.n189 585
R363 B.n188 B.n139 585
R364 B.n187 B.n186 585
R365 B.n185 B.n140 585
R366 B.n184 B.n183 585
R367 B.n182 B.n141 585
R368 B.n181 B.n180 585
R369 B.n179 B.n142 585
R370 B.n178 B.n177 585
R371 B.n176 B.n143 585
R372 B.n175 B.n174 585
R373 B.n173 B.n144 585
R374 B.n172 B.n171 585
R375 B.n170 B.n145 585
R376 B.n169 B.n168 585
R377 B.n167 B.n146 585
R378 B.n166 B.n165 585
R379 B.n164 B.n147 585
R380 B.n163 B.n162 585
R381 B.n161 B.n148 585
R382 B.n160 B.n159 585
R383 B.n158 B.n149 585
R384 B.n157 B.n156 585
R385 B.n155 B.n150 585
R386 B.n154 B.n153 585
R387 B.n152 B.n151 585
R388 B.n2 B.n0 585
R389 B.n573 B.n1 585
R390 B.n572 B.n571 585
R391 B.n570 B.n3 585
R392 B.n569 B.n568 585
R393 B.n567 B.n4 585
R394 B.n566 B.n565 585
R395 B.n564 B.n5 585
R396 B.n563 B.n562 585
R397 B.n561 B.n6 585
R398 B.n560 B.n559 585
R399 B.n558 B.n7 585
R400 B.n557 B.n556 585
R401 B.n555 B.n8 585
R402 B.n554 B.n553 585
R403 B.n552 B.n9 585
R404 B.n551 B.n550 585
R405 B.n549 B.n10 585
R406 B.n548 B.n547 585
R407 B.n546 B.n11 585
R408 B.n545 B.n544 585
R409 B.n543 B.n12 585
R410 B.n542 B.n541 585
R411 B.n540 B.n13 585
R412 B.n539 B.n538 585
R413 B.n537 B.n14 585
R414 B.n536 B.n535 585
R415 B.n534 B.n15 585
R416 B.n533 B.n532 585
R417 B.n531 B.n16 585
R418 B.n530 B.n529 585
R419 B.n575 B.n574 585
R420 B.n195 B.n194 473.281
R421 B.n530 B.n17 473.281
R422 B.n315 B.n92 473.281
R423 B.n409 B.n62 473.281
R424 B.n111 B.t3 359.443
R425 B.n117 B.t6 359.443
R426 B.n36 B.t9 359.443
R427 B.n43 B.t0 359.443
R428 B.n194 B.n193 163.367
R429 B.n193 B.n138 163.367
R430 B.n189 B.n138 163.367
R431 B.n189 B.n188 163.367
R432 B.n188 B.n187 163.367
R433 B.n187 B.n140 163.367
R434 B.n183 B.n140 163.367
R435 B.n183 B.n182 163.367
R436 B.n182 B.n181 163.367
R437 B.n181 B.n142 163.367
R438 B.n177 B.n142 163.367
R439 B.n177 B.n176 163.367
R440 B.n176 B.n175 163.367
R441 B.n175 B.n144 163.367
R442 B.n171 B.n144 163.367
R443 B.n171 B.n170 163.367
R444 B.n170 B.n169 163.367
R445 B.n169 B.n146 163.367
R446 B.n165 B.n146 163.367
R447 B.n165 B.n164 163.367
R448 B.n164 B.n163 163.367
R449 B.n163 B.n148 163.367
R450 B.n159 B.n148 163.367
R451 B.n159 B.n158 163.367
R452 B.n158 B.n157 163.367
R453 B.n157 B.n150 163.367
R454 B.n153 B.n150 163.367
R455 B.n153 B.n152 163.367
R456 B.n152 B.n2 163.367
R457 B.n574 B.n2 163.367
R458 B.n574 B.n573 163.367
R459 B.n573 B.n572 163.367
R460 B.n572 B.n3 163.367
R461 B.n568 B.n3 163.367
R462 B.n568 B.n567 163.367
R463 B.n567 B.n566 163.367
R464 B.n566 B.n5 163.367
R465 B.n562 B.n5 163.367
R466 B.n562 B.n561 163.367
R467 B.n561 B.n560 163.367
R468 B.n560 B.n7 163.367
R469 B.n556 B.n7 163.367
R470 B.n556 B.n555 163.367
R471 B.n555 B.n554 163.367
R472 B.n554 B.n9 163.367
R473 B.n550 B.n9 163.367
R474 B.n550 B.n549 163.367
R475 B.n549 B.n548 163.367
R476 B.n548 B.n11 163.367
R477 B.n544 B.n11 163.367
R478 B.n544 B.n543 163.367
R479 B.n543 B.n542 163.367
R480 B.n542 B.n13 163.367
R481 B.n538 B.n13 163.367
R482 B.n538 B.n537 163.367
R483 B.n537 B.n536 163.367
R484 B.n536 B.n15 163.367
R485 B.n532 B.n15 163.367
R486 B.n532 B.n531 163.367
R487 B.n531 B.n530 163.367
R488 B.n195 B.n136 163.367
R489 B.n199 B.n136 163.367
R490 B.n200 B.n199 163.367
R491 B.n201 B.n200 163.367
R492 B.n201 B.n134 163.367
R493 B.n205 B.n134 163.367
R494 B.n206 B.n205 163.367
R495 B.n207 B.n206 163.367
R496 B.n207 B.n132 163.367
R497 B.n211 B.n132 163.367
R498 B.n212 B.n211 163.367
R499 B.n213 B.n212 163.367
R500 B.n213 B.n130 163.367
R501 B.n217 B.n130 163.367
R502 B.n218 B.n217 163.367
R503 B.n219 B.n218 163.367
R504 B.n219 B.n128 163.367
R505 B.n223 B.n128 163.367
R506 B.n224 B.n223 163.367
R507 B.n225 B.n224 163.367
R508 B.n225 B.n126 163.367
R509 B.n229 B.n126 163.367
R510 B.n230 B.n229 163.367
R511 B.n231 B.n230 163.367
R512 B.n231 B.n124 163.367
R513 B.n235 B.n124 163.367
R514 B.n236 B.n235 163.367
R515 B.n237 B.n236 163.367
R516 B.n237 B.n122 163.367
R517 B.n241 B.n122 163.367
R518 B.n242 B.n241 163.367
R519 B.n243 B.n242 163.367
R520 B.n243 B.n120 163.367
R521 B.n247 B.n120 163.367
R522 B.n248 B.n247 163.367
R523 B.n248 B.n116 163.367
R524 B.n252 B.n116 163.367
R525 B.n253 B.n252 163.367
R526 B.n254 B.n253 163.367
R527 B.n254 B.n114 163.367
R528 B.n258 B.n114 163.367
R529 B.n259 B.n258 163.367
R530 B.n260 B.n259 163.367
R531 B.n260 B.n110 163.367
R532 B.n265 B.n110 163.367
R533 B.n266 B.n265 163.367
R534 B.n267 B.n266 163.367
R535 B.n267 B.n108 163.367
R536 B.n271 B.n108 163.367
R537 B.n272 B.n271 163.367
R538 B.n273 B.n272 163.367
R539 B.n273 B.n106 163.367
R540 B.n277 B.n106 163.367
R541 B.n278 B.n277 163.367
R542 B.n279 B.n278 163.367
R543 B.n279 B.n104 163.367
R544 B.n283 B.n104 163.367
R545 B.n284 B.n283 163.367
R546 B.n285 B.n284 163.367
R547 B.n285 B.n102 163.367
R548 B.n289 B.n102 163.367
R549 B.n290 B.n289 163.367
R550 B.n291 B.n290 163.367
R551 B.n291 B.n100 163.367
R552 B.n295 B.n100 163.367
R553 B.n296 B.n295 163.367
R554 B.n297 B.n296 163.367
R555 B.n297 B.n98 163.367
R556 B.n301 B.n98 163.367
R557 B.n302 B.n301 163.367
R558 B.n303 B.n302 163.367
R559 B.n303 B.n96 163.367
R560 B.n307 B.n96 163.367
R561 B.n308 B.n307 163.367
R562 B.n309 B.n308 163.367
R563 B.n309 B.n94 163.367
R564 B.n313 B.n94 163.367
R565 B.n314 B.n313 163.367
R566 B.n315 B.n314 163.367
R567 B.n319 B.n92 163.367
R568 B.n320 B.n319 163.367
R569 B.n321 B.n320 163.367
R570 B.n321 B.n90 163.367
R571 B.n325 B.n90 163.367
R572 B.n326 B.n325 163.367
R573 B.n327 B.n326 163.367
R574 B.n327 B.n88 163.367
R575 B.n331 B.n88 163.367
R576 B.n332 B.n331 163.367
R577 B.n333 B.n332 163.367
R578 B.n333 B.n86 163.367
R579 B.n337 B.n86 163.367
R580 B.n338 B.n337 163.367
R581 B.n339 B.n338 163.367
R582 B.n339 B.n84 163.367
R583 B.n343 B.n84 163.367
R584 B.n344 B.n343 163.367
R585 B.n345 B.n344 163.367
R586 B.n345 B.n82 163.367
R587 B.n349 B.n82 163.367
R588 B.n350 B.n349 163.367
R589 B.n351 B.n350 163.367
R590 B.n351 B.n80 163.367
R591 B.n355 B.n80 163.367
R592 B.n356 B.n355 163.367
R593 B.n357 B.n356 163.367
R594 B.n357 B.n78 163.367
R595 B.n361 B.n78 163.367
R596 B.n362 B.n361 163.367
R597 B.n363 B.n362 163.367
R598 B.n363 B.n76 163.367
R599 B.n367 B.n76 163.367
R600 B.n368 B.n367 163.367
R601 B.n369 B.n368 163.367
R602 B.n369 B.n74 163.367
R603 B.n373 B.n74 163.367
R604 B.n374 B.n373 163.367
R605 B.n375 B.n374 163.367
R606 B.n375 B.n72 163.367
R607 B.n379 B.n72 163.367
R608 B.n380 B.n379 163.367
R609 B.n381 B.n380 163.367
R610 B.n381 B.n70 163.367
R611 B.n385 B.n70 163.367
R612 B.n386 B.n385 163.367
R613 B.n387 B.n386 163.367
R614 B.n387 B.n68 163.367
R615 B.n391 B.n68 163.367
R616 B.n392 B.n391 163.367
R617 B.n393 B.n392 163.367
R618 B.n393 B.n66 163.367
R619 B.n397 B.n66 163.367
R620 B.n398 B.n397 163.367
R621 B.n399 B.n398 163.367
R622 B.n399 B.n64 163.367
R623 B.n403 B.n64 163.367
R624 B.n404 B.n403 163.367
R625 B.n405 B.n404 163.367
R626 B.n405 B.n62 163.367
R627 B.n526 B.n17 163.367
R628 B.n526 B.n525 163.367
R629 B.n525 B.n524 163.367
R630 B.n524 B.n19 163.367
R631 B.n520 B.n19 163.367
R632 B.n520 B.n519 163.367
R633 B.n519 B.n518 163.367
R634 B.n518 B.n21 163.367
R635 B.n514 B.n21 163.367
R636 B.n514 B.n513 163.367
R637 B.n513 B.n512 163.367
R638 B.n512 B.n23 163.367
R639 B.n508 B.n23 163.367
R640 B.n508 B.n507 163.367
R641 B.n507 B.n506 163.367
R642 B.n506 B.n25 163.367
R643 B.n502 B.n25 163.367
R644 B.n502 B.n501 163.367
R645 B.n501 B.n500 163.367
R646 B.n500 B.n27 163.367
R647 B.n496 B.n27 163.367
R648 B.n496 B.n495 163.367
R649 B.n495 B.n494 163.367
R650 B.n494 B.n29 163.367
R651 B.n490 B.n29 163.367
R652 B.n490 B.n489 163.367
R653 B.n489 B.n488 163.367
R654 B.n488 B.n31 163.367
R655 B.n484 B.n31 163.367
R656 B.n484 B.n483 163.367
R657 B.n483 B.n482 163.367
R658 B.n482 B.n33 163.367
R659 B.n478 B.n33 163.367
R660 B.n478 B.n477 163.367
R661 B.n477 B.n476 163.367
R662 B.n476 B.n35 163.367
R663 B.n472 B.n35 163.367
R664 B.n472 B.n471 163.367
R665 B.n471 B.n470 163.367
R666 B.n470 B.n40 163.367
R667 B.n466 B.n40 163.367
R668 B.n466 B.n465 163.367
R669 B.n465 B.n464 163.367
R670 B.n464 B.n42 163.367
R671 B.n459 B.n42 163.367
R672 B.n459 B.n458 163.367
R673 B.n458 B.n457 163.367
R674 B.n457 B.n46 163.367
R675 B.n453 B.n46 163.367
R676 B.n453 B.n452 163.367
R677 B.n452 B.n451 163.367
R678 B.n451 B.n48 163.367
R679 B.n447 B.n48 163.367
R680 B.n447 B.n446 163.367
R681 B.n446 B.n445 163.367
R682 B.n445 B.n50 163.367
R683 B.n441 B.n50 163.367
R684 B.n441 B.n440 163.367
R685 B.n440 B.n439 163.367
R686 B.n439 B.n52 163.367
R687 B.n435 B.n52 163.367
R688 B.n435 B.n434 163.367
R689 B.n434 B.n433 163.367
R690 B.n433 B.n54 163.367
R691 B.n429 B.n54 163.367
R692 B.n429 B.n428 163.367
R693 B.n428 B.n427 163.367
R694 B.n427 B.n56 163.367
R695 B.n423 B.n56 163.367
R696 B.n423 B.n422 163.367
R697 B.n422 B.n421 163.367
R698 B.n421 B.n58 163.367
R699 B.n417 B.n58 163.367
R700 B.n417 B.n416 163.367
R701 B.n416 B.n415 163.367
R702 B.n415 B.n60 163.367
R703 B.n411 B.n60 163.367
R704 B.n411 B.n410 163.367
R705 B.n410 B.n409 163.367
R706 B.n111 B.t5 148.688
R707 B.n43 B.t1 148.688
R708 B.n117 B.t8 148.677
R709 B.n36 B.t10 148.677
R710 B.n112 B.t4 112.615
R711 B.n44 B.t2 112.615
R712 B.n118 B.t7 112.603
R713 B.n37 B.t11 112.603
R714 B.n263 B.n112 59.5399
R715 B.n119 B.n118 59.5399
R716 B.n38 B.n37 59.5399
R717 B.n461 B.n44 59.5399
R718 B.n112 B.n111 36.0732
R719 B.n118 B.n117 36.0732
R720 B.n37 B.n36 36.0732
R721 B.n44 B.n43 36.0732
R722 B.n529 B.n528 30.7517
R723 B.n408 B.n407 30.7517
R724 B.n317 B.n316 30.7517
R725 B.n196 B.n137 30.7517
R726 B B.n575 18.0485
R727 B.n528 B.n527 10.6151
R728 B.n527 B.n18 10.6151
R729 B.n523 B.n18 10.6151
R730 B.n523 B.n522 10.6151
R731 B.n522 B.n521 10.6151
R732 B.n521 B.n20 10.6151
R733 B.n517 B.n20 10.6151
R734 B.n517 B.n516 10.6151
R735 B.n516 B.n515 10.6151
R736 B.n515 B.n22 10.6151
R737 B.n511 B.n22 10.6151
R738 B.n511 B.n510 10.6151
R739 B.n510 B.n509 10.6151
R740 B.n509 B.n24 10.6151
R741 B.n505 B.n24 10.6151
R742 B.n505 B.n504 10.6151
R743 B.n504 B.n503 10.6151
R744 B.n503 B.n26 10.6151
R745 B.n499 B.n26 10.6151
R746 B.n499 B.n498 10.6151
R747 B.n498 B.n497 10.6151
R748 B.n497 B.n28 10.6151
R749 B.n493 B.n28 10.6151
R750 B.n493 B.n492 10.6151
R751 B.n492 B.n491 10.6151
R752 B.n491 B.n30 10.6151
R753 B.n487 B.n30 10.6151
R754 B.n487 B.n486 10.6151
R755 B.n486 B.n485 10.6151
R756 B.n485 B.n32 10.6151
R757 B.n481 B.n32 10.6151
R758 B.n481 B.n480 10.6151
R759 B.n480 B.n479 10.6151
R760 B.n479 B.n34 10.6151
R761 B.n475 B.n474 10.6151
R762 B.n474 B.n473 10.6151
R763 B.n473 B.n39 10.6151
R764 B.n469 B.n39 10.6151
R765 B.n469 B.n468 10.6151
R766 B.n468 B.n467 10.6151
R767 B.n467 B.n41 10.6151
R768 B.n463 B.n41 10.6151
R769 B.n463 B.n462 10.6151
R770 B.n460 B.n45 10.6151
R771 B.n456 B.n45 10.6151
R772 B.n456 B.n455 10.6151
R773 B.n455 B.n454 10.6151
R774 B.n454 B.n47 10.6151
R775 B.n450 B.n47 10.6151
R776 B.n450 B.n449 10.6151
R777 B.n449 B.n448 10.6151
R778 B.n448 B.n49 10.6151
R779 B.n444 B.n49 10.6151
R780 B.n444 B.n443 10.6151
R781 B.n443 B.n442 10.6151
R782 B.n442 B.n51 10.6151
R783 B.n438 B.n51 10.6151
R784 B.n438 B.n437 10.6151
R785 B.n437 B.n436 10.6151
R786 B.n436 B.n53 10.6151
R787 B.n432 B.n53 10.6151
R788 B.n432 B.n431 10.6151
R789 B.n431 B.n430 10.6151
R790 B.n430 B.n55 10.6151
R791 B.n426 B.n55 10.6151
R792 B.n426 B.n425 10.6151
R793 B.n425 B.n424 10.6151
R794 B.n424 B.n57 10.6151
R795 B.n420 B.n57 10.6151
R796 B.n420 B.n419 10.6151
R797 B.n419 B.n418 10.6151
R798 B.n418 B.n59 10.6151
R799 B.n414 B.n59 10.6151
R800 B.n414 B.n413 10.6151
R801 B.n413 B.n412 10.6151
R802 B.n412 B.n61 10.6151
R803 B.n408 B.n61 10.6151
R804 B.n318 B.n317 10.6151
R805 B.n318 B.n91 10.6151
R806 B.n322 B.n91 10.6151
R807 B.n323 B.n322 10.6151
R808 B.n324 B.n323 10.6151
R809 B.n324 B.n89 10.6151
R810 B.n328 B.n89 10.6151
R811 B.n329 B.n328 10.6151
R812 B.n330 B.n329 10.6151
R813 B.n330 B.n87 10.6151
R814 B.n334 B.n87 10.6151
R815 B.n335 B.n334 10.6151
R816 B.n336 B.n335 10.6151
R817 B.n336 B.n85 10.6151
R818 B.n340 B.n85 10.6151
R819 B.n341 B.n340 10.6151
R820 B.n342 B.n341 10.6151
R821 B.n342 B.n83 10.6151
R822 B.n346 B.n83 10.6151
R823 B.n347 B.n346 10.6151
R824 B.n348 B.n347 10.6151
R825 B.n348 B.n81 10.6151
R826 B.n352 B.n81 10.6151
R827 B.n353 B.n352 10.6151
R828 B.n354 B.n353 10.6151
R829 B.n354 B.n79 10.6151
R830 B.n358 B.n79 10.6151
R831 B.n359 B.n358 10.6151
R832 B.n360 B.n359 10.6151
R833 B.n360 B.n77 10.6151
R834 B.n364 B.n77 10.6151
R835 B.n365 B.n364 10.6151
R836 B.n366 B.n365 10.6151
R837 B.n366 B.n75 10.6151
R838 B.n370 B.n75 10.6151
R839 B.n371 B.n370 10.6151
R840 B.n372 B.n371 10.6151
R841 B.n372 B.n73 10.6151
R842 B.n376 B.n73 10.6151
R843 B.n377 B.n376 10.6151
R844 B.n378 B.n377 10.6151
R845 B.n378 B.n71 10.6151
R846 B.n382 B.n71 10.6151
R847 B.n383 B.n382 10.6151
R848 B.n384 B.n383 10.6151
R849 B.n384 B.n69 10.6151
R850 B.n388 B.n69 10.6151
R851 B.n389 B.n388 10.6151
R852 B.n390 B.n389 10.6151
R853 B.n390 B.n67 10.6151
R854 B.n394 B.n67 10.6151
R855 B.n395 B.n394 10.6151
R856 B.n396 B.n395 10.6151
R857 B.n396 B.n65 10.6151
R858 B.n400 B.n65 10.6151
R859 B.n401 B.n400 10.6151
R860 B.n402 B.n401 10.6151
R861 B.n402 B.n63 10.6151
R862 B.n406 B.n63 10.6151
R863 B.n407 B.n406 10.6151
R864 B.n197 B.n196 10.6151
R865 B.n198 B.n197 10.6151
R866 B.n198 B.n135 10.6151
R867 B.n202 B.n135 10.6151
R868 B.n203 B.n202 10.6151
R869 B.n204 B.n203 10.6151
R870 B.n204 B.n133 10.6151
R871 B.n208 B.n133 10.6151
R872 B.n209 B.n208 10.6151
R873 B.n210 B.n209 10.6151
R874 B.n210 B.n131 10.6151
R875 B.n214 B.n131 10.6151
R876 B.n215 B.n214 10.6151
R877 B.n216 B.n215 10.6151
R878 B.n216 B.n129 10.6151
R879 B.n220 B.n129 10.6151
R880 B.n221 B.n220 10.6151
R881 B.n222 B.n221 10.6151
R882 B.n222 B.n127 10.6151
R883 B.n226 B.n127 10.6151
R884 B.n227 B.n226 10.6151
R885 B.n228 B.n227 10.6151
R886 B.n228 B.n125 10.6151
R887 B.n232 B.n125 10.6151
R888 B.n233 B.n232 10.6151
R889 B.n234 B.n233 10.6151
R890 B.n234 B.n123 10.6151
R891 B.n238 B.n123 10.6151
R892 B.n239 B.n238 10.6151
R893 B.n240 B.n239 10.6151
R894 B.n240 B.n121 10.6151
R895 B.n244 B.n121 10.6151
R896 B.n245 B.n244 10.6151
R897 B.n246 B.n245 10.6151
R898 B.n250 B.n249 10.6151
R899 B.n251 B.n250 10.6151
R900 B.n251 B.n115 10.6151
R901 B.n255 B.n115 10.6151
R902 B.n256 B.n255 10.6151
R903 B.n257 B.n256 10.6151
R904 B.n257 B.n113 10.6151
R905 B.n261 B.n113 10.6151
R906 B.n262 B.n261 10.6151
R907 B.n264 B.n109 10.6151
R908 B.n268 B.n109 10.6151
R909 B.n269 B.n268 10.6151
R910 B.n270 B.n269 10.6151
R911 B.n270 B.n107 10.6151
R912 B.n274 B.n107 10.6151
R913 B.n275 B.n274 10.6151
R914 B.n276 B.n275 10.6151
R915 B.n276 B.n105 10.6151
R916 B.n280 B.n105 10.6151
R917 B.n281 B.n280 10.6151
R918 B.n282 B.n281 10.6151
R919 B.n282 B.n103 10.6151
R920 B.n286 B.n103 10.6151
R921 B.n287 B.n286 10.6151
R922 B.n288 B.n287 10.6151
R923 B.n288 B.n101 10.6151
R924 B.n292 B.n101 10.6151
R925 B.n293 B.n292 10.6151
R926 B.n294 B.n293 10.6151
R927 B.n294 B.n99 10.6151
R928 B.n298 B.n99 10.6151
R929 B.n299 B.n298 10.6151
R930 B.n300 B.n299 10.6151
R931 B.n300 B.n97 10.6151
R932 B.n304 B.n97 10.6151
R933 B.n305 B.n304 10.6151
R934 B.n306 B.n305 10.6151
R935 B.n306 B.n95 10.6151
R936 B.n310 B.n95 10.6151
R937 B.n311 B.n310 10.6151
R938 B.n312 B.n311 10.6151
R939 B.n312 B.n93 10.6151
R940 B.n316 B.n93 10.6151
R941 B.n192 B.n137 10.6151
R942 B.n192 B.n191 10.6151
R943 B.n191 B.n190 10.6151
R944 B.n190 B.n139 10.6151
R945 B.n186 B.n139 10.6151
R946 B.n186 B.n185 10.6151
R947 B.n185 B.n184 10.6151
R948 B.n184 B.n141 10.6151
R949 B.n180 B.n141 10.6151
R950 B.n180 B.n179 10.6151
R951 B.n179 B.n178 10.6151
R952 B.n178 B.n143 10.6151
R953 B.n174 B.n143 10.6151
R954 B.n174 B.n173 10.6151
R955 B.n173 B.n172 10.6151
R956 B.n172 B.n145 10.6151
R957 B.n168 B.n145 10.6151
R958 B.n168 B.n167 10.6151
R959 B.n167 B.n166 10.6151
R960 B.n166 B.n147 10.6151
R961 B.n162 B.n147 10.6151
R962 B.n162 B.n161 10.6151
R963 B.n161 B.n160 10.6151
R964 B.n160 B.n149 10.6151
R965 B.n156 B.n149 10.6151
R966 B.n156 B.n155 10.6151
R967 B.n155 B.n154 10.6151
R968 B.n154 B.n151 10.6151
R969 B.n151 B.n0 10.6151
R970 B.n571 B.n1 10.6151
R971 B.n571 B.n570 10.6151
R972 B.n570 B.n569 10.6151
R973 B.n569 B.n4 10.6151
R974 B.n565 B.n4 10.6151
R975 B.n565 B.n564 10.6151
R976 B.n564 B.n563 10.6151
R977 B.n563 B.n6 10.6151
R978 B.n559 B.n6 10.6151
R979 B.n559 B.n558 10.6151
R980 B.n558 B.n557 10.6151
R981 B.n557 B.n8 10.6151
R982 B.n553 B.n8 10.6151
R983 B.n553 B.n552 10.6151
R984 B.n552 B.n551 10.6151
R985 B.n551 B.n10 10.6151
R986 B.n547 B.n10 10.6151
R987 B.n547 B.n546 10.6151
R988 B.n546 B.n545 10.6151
R989 B.n545 B.n12 10.6151
R990 B.n541 B.n12 10.6151
R991 B.n541 B.n540 10.6151
R992 B.n540 B.n539 10.6151
R993 B.n539 B.n14 10.6151
R994 B.n535 B.n14 10.6151
R995 B.n535 B.n534 10.6151
R996 B.n534 B.n533 10.6151
R997 B.n533 B.n16 10.6151
R998 B.n529 B.n16 10.6151
R999 B.n38 B.n34 9.36635
R1000 B.n461 B.n460 9.36635
R1001 B.n246 B.n119 9.36635
R1002 B.n264 B.n263 9.36635
R1003 B.n575 B.n0 2.81026
R1004 B.n575 B.n1 2.81026
R1005 B.n475 B.n38 1.24928
R1006 B.n462 B.n461 1.24928
R1007 B.n249 B.n119 1.24928
R1008 B.n263 B.n262 1.24928
C0 VTAIL VDD1 6.95514f
C1 VN VTAIL 4.87868f
C2 VP B 1.43482f
C3 B VDD2 1.68161f
C4 VP VTAIL 4.89304f
C5 VTAIL VDD2 6.99799f
C6 w_n2458_n2922# B 7.57338f
C7 VTAIL w_n2458_n2922# 2.58475f
C8 VN VDD1 0.149343f
C9 VP VDD1 5.09311f
C10 VDD1 VDD2 1.01852f
C11 VN VP 5.47632f
C12 VN VDD2 4.87804f
C13 VDD1 w_n2458_n2922# 1.87017f
C14 VN w_n2458_n2922# 4.35955f
C15 VTAIL B 2.74809f
C16 VP VDD2 0.367538f
C17 VP w_n2458_n2922# 4.67435f
C18 w_n2458_n2922# VDD2 1.92083f
C19 VDD1 B 1.63307f
C20 VN B 0.914613f
C21 VDD2 VSUBS 1.344276f
C22 VDD1 VSUBS 1.72197f
C23 VTAIL VSUBS 0.897489f
C24 VN VSUBS 4.77906f
C25 VP VSUBS 2.011246f
C26 B VSUBS 3.39075f
C27 w_n2458_n2922# VSUBS 88.7535f
C28 B.n0 VSUBS 0.004461f
C29 B.n1 VSUBS 0.004461f
C30 B.n2 VSUBS 0.007055f
C31 B.n3 VSUBS 0.007055f
C32 B.n4 VSUBS 0.007055f
C33 B.n5 VSUBS 0.007055f
C34 B.n6 VSUBS 0.007055f
C35 B.n7 VSUBS 0.007055f
C36 B.n8 VSUBS 0.007055f
C37 B.n9 VSUBS 0.007055f
C38 B.n10 VSUBS 0.007055f
C39 B.n11 VSUBS 0.007055f
C40 B.n12 VSUBS 0.007055f
C41 B.n13 VSUBS 0.007055f
C42 B.n14 VSUBS 0.007055f
C43 B.n15 VSUBS 0.007055f
C44 B.n16 VSUBS 0.007055f
C45 B.n17 VSUBS 0.016402f
C46 B.n18 VSUBS 0.007055f
C47 B.n19 VSUBS 0.007055f
C48 B.n20 VSUBS 0.007055f
C49 B.n21 VSUBS 0.007055f
C50 B.n22 VSUBS 0.007055f
C51 B.n23 VSUBS 0.007055f
C52 B.n24 VSUBS 0.007055f
C53 B.n25 VSUBS 0.007055f
C54 B.n26 VSUBS 0.007055f
C55 B.n27 VSUBS 0.007055f
C56 B.n28 VSUBS 0.007055f
C57 B.n29 VSUBS 0.007055f
C58 B.n30 VSUBS 0.007055f
C59 B.n31 VSUBS 0.007055f
C60 B.n32 VSUBS 0.007055f
C61 B.n33 VSUBS 0.007055f
C62 B.n34 VSUBS 0.00664f
C63 B.n35 VSUBS 0.007055f
C64 B.t11 VSUBS 0.313045f
C65 B.t10 VSUBS 0.327033f
C66 B.t9 VSUBS 0.669398f
C67 B.n36 VSUBS 0.151816f
C68 B.n37 VSUBS 0.067717f
C69 B.n38 VSUBS 0.016345f
C70 B.n39 VSUBS 0.007055f
C71 B.n40 VSUBS 0.007055f
C72 B.n41 VSUBS 0.007055f
C73 B.n42 VSUBS 0.007055f
C74 B.t2 VSUBS 0.313041f
C75 B.t1 VSUBS 0.327029f
C76 B.t0 VSUBS 0.669398f
C77 B.n43 VSUBS 0.15182f
C78 B.n44 VSUBS 0.067721f
C79 B.n45 VSUBS 0.007055f
C80 B.n46 VSUBS 0.007055f
C81 B.n47 VSUBS 0.007055f
C82 B.n48 VSUBS 0.007055f
C83 B.n49 VSUBS 0.007055f
C84 B.n50 VSUBS 0.007055f
C85 B.n51 VSUBS 0.007055f
C86 B.n52 VSUBS 0.007055f
C87 B.n53 VSUBS 0.007055f
C88 B.n54 VSUBS 0.007055f
C89 B.n55 VSUBS 0.007055f
C90 B.n56 VSUBS 0.007055f
C91 B.n57 VSUBS 0.007055f
C92 B.n58 VSUBS 0.007055f
C93 B.n59 VSUBS 0.007055f
C94 B.n60 VSUBS 0.007055f
C95 B.n61 VSUBS 0.007055f
C96 B.n62 VSUBS 0.015344f
C97 B.n63 VSUBS 0.007055f
C98 B.n64 VSUBS 0.007055f
C99 B.n65 VSUBS 0.007055f
C100 B.n66 VSUBS 0.007055f
C101 B.n67 VSUBS 0.007055f
C102 B.n68 VSUBS 0.007055f
C103 B.n69 VSUBS 0.007055f
C104 B.n70 VSUBS 0.007055f
C105 B.n71 VSUBS 0.007055f
C106 B.n72 VSUBS 0.007055f
C107 B.n73 VSUBS 0.007055f
C108 B.n74 VSUBS 0.007055f
C109 B.n75 VSUBS 0.007055f
C110 B.n76 VSUBS 0.007055f
C111 B.n77 VSUBS 0.007055f
C112 B.n78 VSUBS 0.007055f
C113 B.n79 VSUBS 0.007055f
C114 B.n80 VSUBS 0.007055f
C115 B.n81 VSUBS 0.007055f
C116 B.n82 VSUBS 0.007055f
C117 B.n83 VSUBS 0.007055f
C118 B.n84 VSUBS 0.007055f
C119 B.n85 VSUBS 0.007055f
C120 B.n86 VSUBS 0.007055f
C121 B.n87 VSUBS 0.007055f
C122 B.n88 VSUBS 0.007055f
C123 B.n89 VSUBS 0.007055f
C124 B.n90 VSUBS 0.007055f
C125 B.n91 VSUBS 0.007055f
C126 B.n92 VSUBS 0.015344f
C127 B.n93 VSUBS 0.007055f
C128 B.n94 VSUBS 0.007055f
C129 B.n95 VSUBS 0.007055f
C130 B.n96 VSUBS 0.007055f
C131 B.n97 VSUBS 0.007055f
C132 B.n98 VSUBS 0.007055f
C133 B.n99 VSUBS 0.007055f
C134 B.n100 VSUBS 0.007055f
C135 B.n101 VSUBS 0.007055f
C136 B.n102 VSUBS 0.007055f
C137 B.n103 VSUBS 0.007055f
C138 B.n104 VSUBS 0.007055f
C139 B.n105 VSUBS 0.007055f
C140 B.n106 VSUBS 0.007055f
C141 B.n107 VSUBS 0.007055f
C142 B.n108 VSUBS 0.007055f
C143 B.n109 VSUBS 0.007055f
C144 B.n110 VSUBS 0.007055f
C145 B.t4 VSUBS 0.313041f
C146 B.t5 VSUBS 0.327029f
C147 B.t3 VSUBS 0.669398f
C148 B.n111 VSUBS 0.15182f
C149 B.n112 VSUBS 0.067721f
C150 B.n113 VSUBS 0.007055f
C151 B.n114 VSUBS 0.007055f
C152 B.n115 VSUBS 0.007055f
C153 B.n116 VSUBS 0.007055f
C154 B.t7 VSUBS 0.313045f
C155 B.t8 VSUBS 0.327033f
C156 B.t6 VSUBS 0.669398f
C157 B.n117 VSUBS 0.151816f
C158 B.n118 VSUBS 0.067717f
C159 B.n119 VSUBS 0.016345f
C160 B.n120 VSUBS 0.007055f
C161 B.n121 VSUBS 0.007055f
C162 B.n122 VSUBS 0.007055f
C163 B.n123 VSUBS 0.007055f
C164 B.n124 VSUBS 0.007055f
C165 B.n125 VSUBS 0.007055f
C166 B.n126 VSUBS 0.007055f
C167 B.n127 VSUBS 0.007055f
C168 B.n128 VSUBS 0.007055f
C169 B.n129 VSUBS 0.007055f
C170 B.n130 VSUBS 0.007055f
C171 B.n131 VSUBS 0.007055f
C172 B.n132 VSUBS 0.007055f
C173 B.n133 VSUBS 0.007055f
C174 B.n134 VSUBS 0.007055f
C175 B.n135 VSUBS 0.007055f
C176 B.n136 VSUBS 0.007055f
C177 B.n137 VSUBS 0.015344f
C178 B.n138 VSUBS 0.007055f
C179 B.n139 VSUBS 0.007055f
C180 B.n140 VSUBS 0.007055f
C181 B.n141 VSUBS 0.007055f
C182 B.n142 VSUBS 0.007055f
C183 B.n143 VSUBS 0.007055f
C184 B.n144 VSUBS 0.007055f
C185 B.n145 VSUBS 0.007055f
C186 B.n146 VSUBS 0.007055f
C187 B.n147 VSUBS 0.007055f
C188 B.n148 VSUBS 0.007055f
C189 B.n149 VSUBS 0.007055f
C190 B.n150 VSUBS 0.007055f
C191 B.n151 VSUBS 0.007055f
C192 B.n152 VSUBS 0.007055f
C193 B.n153 VSUBS 0.007055f
C194 B.n154 VSUBS 0.007055f
C195 B.n155 VSUBS 0.007055f
C196 B.n156 VSUBS 0.007055f
C197 B.n157 VSUBS 0.007055f
C198 B.n158 VSUBS 0.007055f
C199 B.n159 VSUBS 0.007055f
C200 B.n160 VSUBS 0.007055f
C201 B.n161 VSUBS 0.007055f
C202 B.n162 VSUBS 0.007055f
C203 B.n163 VSUBS 0.007055f
C204 B.n164 VSUBS 0.007055f
C205 B.n165 VSUBS 0.007055f
C206 B.n166 VSUBS 0.007055f
C207 B.n167 VSUBS 0.007055f
C208 B.n168 VSUBS 0.007055f
C209 B.n169 VSUBS 0.007055f
C210 B.n170 VSUBS 0.007055f
C211 B.n171 VSUBS 0.007055f
C212 B.n172 VSUBS 0.007055f
C213 B.n173 VSUBS 0.007055f
C214 B.n174 VSUBS 0.007055f
C215 B.n175 VSUBS 0.007055f
C216 B.n176 VSUBS 0.007055f
C217 B.n177 VSUBS 0.007055f
C218 B.n178 VSUBS 0.007055f
C219 B.n179 VSUBS 0.007055f
C220 B.n180 VSUBS 0.007055f
C221 B.n181 VSUBS 0.007055f
C222 B.n182 VSUBS 0.007055f
C223 B.n183 VSUBS 0.007055f
C224 B.n184 VSUBS 0.007055f
C225 B.n185 VSUBS 0.007055f
C226 B.n186 VSUBS 0.007055f
C227 B.n187 VSUBS 0.007055f
C228 B.n188 VSUBS 0.007055f
C229 B.n189 VSUBS 0.007055f
C230 B.n190 VSUBS 0.007055f
C231 B.n191 VSUBS 0.007055f
C232 B.n192 VSUBS 0.007055f
C233 B.n193 VSUBS 0.007055f
C234 B.n194 VSUBS 0.015344f
C235 B.n195 VSUBS 0.016402f
C236 B.n196 VSUBS 0.016402f
C237 B.n197 VSUBS 0.007055f
C238 B.n198 VSUBS 0.007055f
C239 B.n199 VSUBS 0.007055f
C240 B.n200 VSUBS 0.007055f
C241 B.n201 VSUBS 0.007055f
C242 B.n202 VSUBS 0.007055f
C243 B.n203 VSUBS 0.007055f
C244 B.n204 VSUBS 0.007055f
C245 B.n205 VSUBS 0.007055f
C246 B.n206 VSUBS 0.007055f
C247 B.n207 VSUBS 0.007055f
C248 B.n208 VSUBS 0.007055f
C249 B.n209 VSUBS 0.007055f
C250 B.n210 VSUBS 0.007055f
C251 B.n211 VSUBS 0.007055f
C252 B.n212 VSUBS 0.007055f
C253 B.n213 VSUBS 0.007055f
C254 B.n214 VSUBS 0.007055f
C255 B.n215 VSUBS 0.007055f
C256 B.n216 VSUBS 0.007055f
C257 B.n217 VSUBS 0.007055f
C258 B.n218 VSUBS 0.007055f
C259 B.n219 VSUBS 0.007055f
C260 B.n220 VSUBS 0.007055f
C261 B.n221 VSUBS 0.007055f
C262 B.n222 VSUBS 0.007055f
C263 B.n223 VSUBS 0.007055f
C264 B.n224 VSUBS 0.007055f
C265 B.n225 VSUBS 0.007055f
C266 B.n226 VSUBS 0.007055f
C267 B.n227 VSUBS 0.007055f
C268 B.n228 VSUBS 0.007055f
C269 B.n229 VSUBS 0.007055f
C270 B.n230 VSUBS 0.007055f
C271 B.n231 VSUBS 0.007055f
C272 B.n232 VSUBS 0.007055f
C273 B.n233 VSUBS 0.007055f
C274 B.n234 VSUBS 0.007055f
C275 B.n235 VSUBS 0.007055f
C276 B.n236 VSUBS 0.007055f
C277 B.n237 VSUBS 0.007055f
C278 B.n238 VSUBS 0.007055f
C279 B.n239 VSUBS 0.007055f
C280 B.n240 VSUBS 0.007055f
C281 B.n241 VSUBS 0.007055f
C282 B.n242 VSUBS 0.007055f
C283 B.n243 VSUBS 0.007055f
C284 B.n244 VSUBS 0.007055f
C285 B.n245 VSUBS 0.007055f
C286 B.n246 VSUBS 0.00664f
C287 B.n247 VSUBS 0.007055f
C288 B.n248 VSUBS 0.007055f
C289 B.n249 VSUBS 0.003942f
C290 B.n250 VSUBS 0.007055f
C291 B.n251 VSUBS 0.007055f
C292 B.n252 VSUBS 0.007055f
C293 B.n253 VSUBS 0.007055f
C294 B.n254 VSUBS 0.007055f
C295 B.n255 VSUBS 0.007055f
C296 B.n256 VSUBS 0.007055f
C297 B.n257 VSUBS 0.007055f
C298 B.n258 VSUBS 0.007055f
C299 B.n259 VSUBS 0.007055f
C300 B.n260 VSUBS 0.007055f
C301 B.n261 VSUBS 0.007055f
C302 B.n262 VSUBS 0.003942f
C303 B.n263 VSUBS 0.016345f
C304 B.n264 VSUBS 0.00664f
C305 B.n265 VSUBS 0.007055f
C306 B.n266 VSUBS 0.007055f
C307 B.n267 VSUBS 0.007055f
C308 B.n268 VSUBS 0.007055f
C309 B.n269 VSUBS 0.007055f
C310 B.n270 VSUBS 0.007055f
C311 B.n271 VSUBS 0.007055f
C312 B.n272 VSUBS 0.007055f
C313 B.n273 VSUBS 0.007055f
C314 B.n274 VSUBS 0.007055f
C315 B.n275 VSUBS 0.007055f
C316 B.n276 VSUBS 0.007055f
C317 B.n277 VSUBS 0.007055f
C318 B.n278 VSUBS 0.007055f
C319 B.n279 VSUBS 0.007055f
C320 B.n280 VSUBS 0.007055f
C321 B.n281 VSUBS 0.007055f
C322 B.n282 VSUBS 0.007055f
C323 B.n283 VSUBS 0.007055f
C324 B.n284 VSUBS 0.007055f
C325 B.n285 VSUBS 0.007055f
C326 B.n286 VSUBS 0.007055f
C327 B.n287 VSUBS 0.007055f
C328 B.n288 VSUBS 0.007055f
C329 B.n289 VSUBS 0.007055f
C330 B.n290 VSUBS 0.007055f
C331 B.n291 VSUBS 0.007055f
C332 B.n292 VSUBS 0.007055f
C333 B.n293 VSUBS 0.007055f
C334 B.n294 VSUBS 0.007055f
C335 B.n295 VSUBS 0.007055f
C336 B.n296 VSUBS 0.007055f
C337 B.n297 VSUBS 0.007055f
C338 B.n298 VSUBS 0.007055f
C339 B.n299 VSUBS 0.007055f
C340 B.n300 VSUBS 0.007055f
C341 B.n301 VSUBS 0.007055f
C342 B.n302 VSUBS 0.007055f
C343 B.n303 VSUBS 0.007055f
C344 B.n304 VSUBS 0.007055f
C345 B.n305 VSUBS 0.007055f
C346 B.n306 VSUBS 0.007055f
C347 B.n307 VSUBS 0.007055f
C348 B.n308 VSUBS 0.007055f
C349 B.n309 VSUBS 0.007055f
C350 B.n310 VSUBS 0.007055f
C351 B.n311 VSUBS 0.007055f
C352 B.n312 VSUBS 0.007055f
C353 B.n313 VSUBS 0.007055f
C354 B.n314 VSUBS 0.007055f
C355 B.n315 VSUBS 0.016402f
C356 B.n316 VSUBS 0.016402f
C357 B.n317 VSUBS 0.015344f
C358 B.n318 VSUBS 0.007055f
C359 B.n319 VSUBS 0.007055f
C360 B.n320 VSUBS 0.007055f
C361 B.n321 VSUBS 0.007055f
C362 B.n322 VSUBS 0.007055f
C363 B.n323 VSUBS 0.007055f
C364 B.n324 VSUBS 0.007055f
C365 B.n325 VSUBS 0.007055f
C366 B.n326 VSUBS 0.007055f
C367 B.n327 VSUBS 0.007055f
C368 B.n328 VSUBS 0.007055f
C369 B.n329 VSUBS 0.007055f
C370 B.n330 VSUBS 0.007055f
C371 B.n331 VSUBS 0.007055f
C372 B.n332 VSUBS 0.007055f
C373 B.n333 VSUBS 0.007055f
C374 B.n334 VSUBS 0.007055f
C375 B.n335 VSUBS 0.007055f
C376 B.n336 VSUBS 0.007055f
C377 B.n337 VSUBS 0.007055f
C378 B.n338 VSUBS 0.007055f
C379 B.n339 VSUBS 0.007055f
C380 B.n340 VSUBS 0.007055f
C381 B.n341 VSUBS 0.007055f
C382 B.n342 VSUBS 0.007055f
C383 B.n343 VSUBS 0.007055f
C384 B.n344 VSUBS 0.007055f
C385 B.n345 VSUBS 0.007055f
C386 B.n346 VSUBS 0.007055f
C387 B.n347 VSUBS 0.007055f
C388 B.n348 VSUBS 0.007055f
C389 B.n349 VSUBS 0.007055f
C390 B.n350 VSUBS 0.007055f
C391 B.n351 VSUBS 0.007055f
C392 B.n352 VSUBS 0.007055f
C393 B.n353 VSUBS 0.007055f
C394 B.n354 VSUBS 0.007055f
C395 B.n355 VSUBS 0.007055f
C396 B.n356 VSUBS 0.007055f
C397 B.n357 VSUBS 0.007055f
C398 B.n358 VSUBS 0.007055f
C399 B.n359 VSUBS 0.007055f
C400 B.n360 VSUBS 0.007055f
C401 B.n361 VSUBS 0.007055f
C402 B.n362 VSUBS 0.007055f
C403 B.n363 VSUBS 0.007055f
C404 B.n364 VSUBS 0.007055f
C405 B.n365 VSUBS 0.007055f
C406 B.n366 VSUBS 0.007055f
C407 B.n367 VSUBS 0.007055f
C408 B.n368 VSUBS 0.007055f
C409 B.n369 VSUBS 0.007055f
C410 B.n370 VSUBS 0.007055f
C411 B.n371 VSUBS 0.007055f
C412 B.n372 VSUBS 0.007055f
C413 B.n373 VSUBS 0.007055f
C414 B.n374 VSUBS 0.007055f
C415 B.n375 VSUBS 0.007055f
C416 B.n376 VSUBS 0.007055f
C417 B.n377 VSUBS 0.007055f
C418 B.n378 VSUBS 0.007055f
C419 B.n379 VSUBS 0.007055f
C420 B.n380 VSUBS 0.007055f
C421 B.n381 VSUBS 0.007055f
C422 B.n382 VSUBS 0.007055f
C423 B.n383 VSUBS 0.007055f
C424 B.n384 VSUBS 0.007055f
C425 B.n385 VSUBS 0.007055f
C426 B.n386 VSUBS 0.007055f
C427 B.n387 VSUBS 0.007055f
C428 B.n388 VSUBS 0.007055f
C429 B.n389 VSUBS 0.007055f
C430 B.n390 VSUBS 0.007055f
C431 B.n391 VSUBS 0.007055f
C432 B.n392 VSUBS 0.007055f
C433 B.n393 VSUBS 0.007055f
C434 B.n394 VSUBS 0.007055f
C435 B.n395 VSUBS 0.007055f
C436 B.n396 VSUBS 0.007055f
C437 B.n397 VSUBS 0.007055f
C438 B.n398 VSUBS 0.007055f
C439 B.n399 VSUBS 0.007055f
C440 B.n400 VSUBS 0.007055f
C441 B.n401 VSUBS 0.007055f
C442 B.n402 VSUBS 0.007055f
C443 B.n403 VSUBS 0.007055f
C444 B.n404 VSUBS 0.007055f
C445 B.n405 VSUBS 0.007055f
C446 B.n406 VSUBS 0.007055f
C447 B.n407 VSUBS 0.01623f
C448 B.n408 VSUBS 0.015517f
C449 B.n409 VSUBS 0.016402f
C450 B.n410 VSUBS 0.007055f
C451 B.n411 VSUBS 0.007055f
C452 B.n412 VSUBS 0.007055f
C453 B.n413 VSUBS 0.007055f
C454 B.n414 VSUBS 0.007055f
C455 B.n415 VSUBS 0.007055f
C456 B.n416 VSUBS 0.007055f
C457 B.n417 VSUBS 0.007055f
C458 B.n418 VSUBS 0.007055f
C459 B.n419 VSUBS 0.007055f
C460 B.n420 VSUBS 0.007055f
C461 B.n421 VSUBS 0.007055f
C462 B.n422 VSUBS 0.007055f
C463 B.n423 VSUBS 0.007055f
C464 B.n424 VSUBS 0.007055f
C465 B.n425 VSUBS 0.007055f
C466 B.n426 VSUBS 0.007055f
C467 B.n427 VSUBS 0.007055f
C468 B.n428 VSUBS 0.007055f
C469 B.n429 VSUBS 0.007055f
C470 B.n430 VSUBS 0.007055f
C471 B.n431 VSUBS 0.007055f
C472 B.n432 VSUBS 0.007055f
C473 B.n433 VSUBS 0.007055f
C474 B.n434 VSUBS 0.007055f
C475 B.n435 VSUBS 0.007055f
C476 B.n436 VSUBS 0.007055f
C477 B.n437 VSUBS 0.007055f
C478 B.n438 VSUBS 0.007055f
C479 B.n439 VSUBS 0.007055f
C480 B.n440 VSUBS 0.007055f
C481 B.n441 VSUBS 0.007055f
C482 B.n442 VSUBS 0.007055f
C483 B.n443 VSUBS 0.007055f
C484 B.n444 VSUBS 0.007055f
C485 B.n445 VSUBS 0.007055f
C486 B.n446 VSUBS 0.007055f
C487 B.n447 VSUBS 0.007055f
C488 B.n448 VSUBS 0.007055f
C489 B.n449 VSUBS 0.007055f
C490 B.n450 VSUBS 0.007055f
C491 B.n451 VSUBS 0.007055f
C492 B.n452 VSUBS 0.007055f
C493 B.n453 VSUBS 0.007055f
C494 B.n454 VSUBS 0.007055f
C495 B.n455 VSUBS 0.007055f
C496 B.n456 VSUBS 0.007055f
C497 B.n457 VSUBS 0.007055f
C498 B.n458 VSUBS 0.007055f
C499 B.n459 VSUBS 0.007055f
C500 B.n460 VSUBS 0.00664f
C501 B.n461 VSUBS 0.016345f
C502 B.n462 VSUBS 0.003942f
C503 B.n463 VSUBS 0.007055f
C504 B.n464 VSUBS 0.007055f
C505 B.n465 VSUBS 0.007055f
C506 B.n466 VSUBS 0.007055f
C507 B.n467 VSUBS 0.007055f
C508 B.n468 VSUBS 0.007055f
C509 B.n469 VSUBS 0.007055f
C510 B.n470 VSUBS 0.007055f
C511 B.n471 VSUBS 0.007055f
C512 B.n472 VSUBS 0.007055f
C513 B.n473 VSUBS 0.007055f
C514 B.n474 VSUBS 0.007055f
C515 B.n475 VSUBS 0.003942f
C516 B.n476 VSUBS 0.007055f
C517 B.n477 VSUBS 0.007055f
C518 B.n478 VSUBS 0.007055f
C519 B.n479 VSUBS 0.007055f
C520 B.n480 VSUBS 0.007055f
C521 B.n481 VSUBS 0.007055f
C522 B.n482 VSUBS 0.007055f
C523 B.n483 VSUBS 0.007055f
C524 B.n484 VSUBS 0.007055f
C525 B.n485 VSUBS 0.007055f
C526 B.n486 VSUBS 0.007055f
C527 B.n487 VSUBS 0.007055f
C528 B.n488 VSUBS 0.007055f
C529 B.n489 VSUBS 0.007055f
C530 B.n490 VSUBS 0.007055f
C531 B.n491 VSUBS 0.007055f
C532 B.n492 VSUBS 0.007055f
C533 B.n493 VSUBS 0.007055f
C534 B.n494 VSUBS 0.007055f
C535 B.n495 VSUBS 0.007055f
C536 B.n496 VSUBS 0.007055f
C537 B.n497 VSUBS 0.007055f
C538 B.n498 VSUBS 0.007055f
C539 B.n499 VSUBS 0.007055f
C540 B.n500 VSUBS 0.007055f
C541 B.n501 VSUBS 0.007055f
C542 B.n502 VSUBS 0.007055f
C543 B.n503 VSUBS 0.007055f
C544 B.n504 VSUBS 0.007055f
C545 B.n505 VSUBS 0.007055f
C546 B.n506 VSUBS 0.007055f
C547 B.n507 VSUBS 0.007055f
C548 B.n508 VSUBS 0.007055f
C549 B.n509 VSUBS 0.007055f
C550 B.n510 VSUBS 0.007055f
C551 B.n511 VSUBS 0.007055f
C552 B.n512 VSUBS 0.007055f
C553 B.n513 VSUBS 0.007055f
C554 B.n514 VSUBS 0.007055f
C555 B.n515 VSUBS 0.007055f
C556 B.n516 VSUBS 0.007055f
C557 B.n517 VSUBS 0.007055f
C558 B.n518 VSUBS 0.007055f
C559 B.n519 VSUBS 0.007055f
C560 B.n520 VSUBS 0.007055f
C561 B.n521 VSUBS 0.007055f
C562 B.n522 VSUBS 0.007055f
C563 B.n523 VSUBS 0.007055f
C564 B.n524 VSUBS 0.007055f
C565 B.n525 VSUBS 0.007055f
C566 B.n526 VSUBS 0.007055f
C567 B.n527 VSUBS 0.007055f
C568 B.n528 VSUBS 0.016402f
C569 B.n529 VSUBS 0.015344f
C570 B.n530 VSUBS 0.015344f
C571 B.n531 VSUBS 0.007055f
C572 B.n532 VSUBS 0.007055f
C573 B.n533 VSUBS 0.007055f
C574 B.n534 VSUBS 0.007055f
C575 B.n535 VSUBS 0.007055f
C576 B.n536 VSUBS 0.007055f
C577 B.n537 VSUBS 0.007055f
C578 B.n538 VSUBS 0.007055f
C579 B.n539 VSUBS 0.007055f
C580 B.n540 VSUBS 0.007055f
C581 B.n541 VSUBS 0.007055f
C582 B.n542 VSUBS 0.007055f
C583 B.n543 VSUBS 0.007055f
C584 B.n544 VSUBS 0.007055f
C585 B.n545 VSUBS 0.007055f
C586 B.n546 VSUBS 0.007055f
C587 B.n547 VSUBS 0.007055f
C588 B.n548 VSUBS 0.007055f
C589 B.n549 VSUBS 0.007055f
C590 B.n550 VSUBS 0.007055f
C591 B.n551 VSUBS 0.007055f
C592 B.n552 VSUBS 0.007055f
C593 B.n553 VSUBS 0.007055f
C594 B.n554 VSUBS 0.007055f
C595 B.n555 VSUBS 0.007055f
C596 B.n556 VSUBS 0.007055f
C597 B.n557 VSUBS 0.007055f
C598 B.n558 VSUBS 0.007055f
C599 B.n559 VSUBS 0.007055f
C600 B.n560 VSUBS 0.007055f
C601 B.n561 VSUBS 0.007055f
C602 B.n562 VSUBS 0.007055f
C603 B.n563 VSUBS 0.007055f
C604 B.n564 VSUBS 0.007055f
C605 B.n565 VSUBS 0.007055f
C606 B.n566 VSUBS 0.007055f
C607 B.n567 VSUBS 0.007055f
C608 B.n568 VSUBS 0.007055f
C609 B.n569 VSUBS 0.007055f
C610 B.n570 VSUBS 0.007055f
C611 B.n571 VSUBS 0.007055f
C612 B.n572 VSUBS 0.007055f
C613 B.n573 VSUBS 0.007055f
C614 B.n574 VSUBS 0.007055f
C615 B.n575 VSUBS 0.015975f
C616 VDD1.t2 VSUBS 1.69842f
C617 VDD1.t4 VSUBS 1.69759f
C618 VDD1.t1 VSUBS 0.17033f
C619 VDD1.t5 VSUBS 0.17033f
C620 VDD1.n0 VSUBS 1.29041f
C621 VDD1.n1 VSUBS 2.53856f
C622 VDD1.t3 VSUBS 0.17033f
C623 VDD1.t0 VSUBS 0.17033f
C624 VDD1.n2 VSUBS 1.28813f
C625 VDD1.n3 VSUBS 2.2501f
C626 VP.n0 VSUBS 0.043322f
C627 VP.t0 VSUBS 1.75289f
C628 VP.n1 VSUBS 0.054791f
C629 VP.n2 VSUBS 0.043322f
C630 VP.t4 VSUBS 1.75289f
C631 VP.n3 VSUBS 0.071692f
C632 VP.n4 VSUBS 0.043322f
C633 VP.t5 VSUBS 1.75289f
C634 VP.n5 VSUBS 0.054791f
C635 VP.t3 VSUBS 1.89017f
C636 VP.n6 VSUBS 0.749492f
C637 VP.t2 VSUBS 1.75289f
C638 VP.n7 VSUBS 0.726437f
C639 VP.n8 VSUBS 0.060809f
C640 VP.n9 VSUBS 0.271833f
C641 VP.n10 VSUBS 0.043322f
C642 VP.n11 VSUBS 0.043322f
C643 VP.n12 VSUBS 0.071692f
C644 VP.n13 VSUBS 0.049648f
C645 VP.n14 VSUBS 0.726976f
C646 VP.n15 VSUBS 1.84416f
C647 VP.n16 VSUBS 1.88067f
C648 VP.t1 VSUBS 1.75289f
C649 VP.n17 VSUBS 0.726976f
C650 VP.n18 VSUBS 0.049648f
C651 VP.n19 VSUBS 0.043322f
C652 VP.n20 VSUBS 0.043322f
C653 VP.n21 VSUBS 0.043322f
C654 VP.n22 VSUBS 0.054791f
C655 VP.n23 VSUBS 0.060809f
C656 VP.n24 VSUBS 0.644797f
C657 VP.n25 VSUBS 0.060809f
C658 VP.n26 VSUBS 0.043322f
C659 VP.n27 VSUBS 0.043322f
C660 VP.n28 VSUBS 0.043322f
C661 VP.n29 VSUBS 0.071692f
C662 VP.n30 VSUBS 0.049648f
C663 VP.n31 VSUBS 0.726976f
C664 VP.n32 VSUBS 0.043295f
C665 VDD2.t2 VSUBS 1.68085f
C666 VDD2.t4 VSUBS 0.168651f
C667 VDD2.t3 VSUBS 0.168651f
C668 VDD2.n0 VSUBS 1.27769f
C669 VDD2.n1 VSUBS 2.42995f
C670 VDD2.t5 VSUBS 1.67366f
C671 VDD2.n2 VSUBS 2.24429f
C672 VDD2.t1 VSUBS 0.168651f
C673 VDD2.t0 VSUBS 0.168651f
C674 VDD2.n3 VSUBS 1.27766f
C675 VTAIL.t8 VSUBS 0.225846f
C676 VTAIL.t9 VSUBS 0.225846f
C677 VTAIL.n0 VSUBS 1.576f
C678 VTAIL.n1 VSUBS 0.770759f
C679 VTAIL.t0 VSUBS 2.09541f
C680 VTAIL.n2 VSUBS 0.975161f
C681 VTAIL.t2 VSUBS 0.225846f
C682 VTAIL.t1 VSUBS 0.225846f
C683 VTAIL.n3 VSUBS 1.576f
C684 VTAIL.n4 VSUBS 2.2523f
C685 VTAIL.t10 VSUBS 0.225846f
C686 VTAIL.t7 VSUBS 0.225846f
C687 VTAIL.n5 VSUBS 1.57601f
C688 VTAIL.n6 VSUBS 2.25229f
C689 VTAIL.t11 VSUBS 2.09543f
C690 VTAIL.n7 VSUBS 0.975147f
C691 VTAIL.t5 VSUBS 0.225846f
C692 VTAIL.t3 VSUBS 0.225846f
C693 VTAIL.n8 VSUBS 1.57601f
C694 VTAIL.n9 VSUBS 0.878623f
C695 VTAIL.t4 VSUBS 2.09541f
C696 VTAIL.n10 VSUBS 2.19769f
C697 VTAIL.t6 VSUBS 2.09541f
C698 VTAIL.n11 VSUBS 2.15442f
C699 VN.n0 VSUBS 0.042122f
C700 VN.t2 VSUBS 1.70436f
C701 VN.n1 VSUBS 0.053274f
C702 VN.t3 VSUBS 1.83784f
C703 VN.n2 VSUBS 0.728743f
C704 VN.t1 VSUBS 1.70436f
C705 VN.n3 VSUBS 0.706326f
C706 VN.n4 VSUBS 0.059126f
C707 VN.n5 VSUBS 0.264308f
C708 VN.n6 VSUBS 0.042122f
C709 VN.n7 VSUBS 0.042122f
C710 VN.n8 VSUBS 0.069707f
C711 VN.n9 VSUBS 0.048274f
C712 VN.n10 VSUBS 0.70685f
C713 VN.n11 VSUBS 0.042097f
C714 VN.n12 VSUBS 0.042122f
C715 VN.t0 VSUBS 1.70436f
C716 VN.n13 VSUBS 0.053274f
C717 VN.t5 VSUBS 1.83784f
C718 VN.n14 VSUBS 0.728743f
C719 VN.t4 VSUBS 1.70436f
C720 VN.n15 VSUBS 0.706326f
C721 VN.n16 VSUBS 0.059126f
C722 VN.n17 VSUBS 0.264308f
C723 VN.n18 VSUBS 0.042122f
C724 VN.n19 VSUBS 0.042122f
C725 VN.n20 VSUBS 0.069707f
C726 VN.n21 VSUBS 0.048274f
C727 VN.n22 VSUBS 0.70685f
C728 VN.n23 VSUBS 1.82073f
.ends

