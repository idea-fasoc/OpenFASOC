* NGSPICE file created from diff_pair_sample_1458.ext - technology: sky130A

.subckt diff_pair_sample_1458 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=0 ps=0 w=19.33 l=3.01
X1 VDD1.t5 VP.t0 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=3.18945 ps=19.66 w=19.33 l=3.01
X2 VDD2.t5 VN.t0 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=3.18945 ps=19.66 w=19.33 l=3.01
X3 VDD1.t4 VP.t1 VTAIL.t9 B.t19 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=3.18945 ps=19.66 w=19.33 l=3.01
X4 VDD2.t4 VN.t1 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=3.18945 ps=19.66 w=19.33 l=3.01
X5 VDD1.t3 VP.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=7.5387 ps=39.44 w=19.33 l=3.01
X6 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=7.5387 ps=39.44 w=19.33 l=3.01
X7 VTAIL.t7 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=3.18945 ps=19.66 w=19.33 l=3.01
X8 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=0 ps=0 w=19.33 l=3.01
X9 VTAIL.t6 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=3.18945 ps=19.66 w=19.33 l=3.01
X10 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=7.5387 ps=39.44 w=19.33 l=3.01
X11 VTAIL.t4 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=3.18945 ps=19.66 w=19.33 l=3.01
X12 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=0 ps=0 w=19.33 l=3.01
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=7.5387 pd=39.44 as=0 ps=0 w=19.33 l=3.01
X14 VDD1.t0 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=7.5387 ps=39.44 w=19.33 l=3.01
X15 VTAIL.t3 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=3.18945 pd=19.66 as=3.18945 ps=19.66 w=19.33 l=3.01
R0 B.n1069 B.n1068 585
R1 B.n428 B.n156 585
R2 B.n427 B.n426 585
R3 B.n425 B.n424 585
R4 B.n423 B.n422 585
R5 B.n421 B.n420 585
R6 B.n419 B.n418 585
R7 B.n417 B.n416 585
R8 B.n415 B.n414 585
R9 B.n413 B.n412 585
R10 B.n411 B.n410 585
R11 B.n409 B.n408 585
R12 B.n407 B.n406 585
R13 B.n405 B.n404 585
R14 B.n403 B.n402 585
R15 B.n401 B.n400 585
R16 B.n399 B.n398 585
R17 B.n397 B.n396 585
R18 B.n395 B.n394 585
R19 B.n393 B.n392 585
R20 B.n391 B.n390 585
R21 B.n389 B.n388 585
R22 B.n387 B.n386 585
R23 B.n385 B.n384 585
R24 B.n383 B.n382 585
R25 B.n381 B.n380 585
R26 B.n379 B.n378 585
R27 B.n377 B.n376 585
R28 B.n375 B.n374 585
R29 B.n373 B.n372 585
R30 B.n371 B.n370 585
R31 B.n369 B.n368 585
R32 B.n367 B.n366 585
R33 B.n365 B.n364 585
R34 B.n363 B.n362 585
R35 B.n361 B.n360 585
R36 B.n359 B.n358 585
R37 B.n357 B.n356 585
R38 B.n355 B.n354 585
R39 B.n353 B.n352 585
R40 B.n351 B.n350 585
R41 B.n349 B.n348 585
R42 B.n347 B.n346 585
R43 B.n345 B.n344 585
R44 B.n343 B.n342 585
R45 B.n341 B.n340 585
R46 B.n339 B.n338 585
R47 B.n337 B.n336 585
R48 B.n335 B.n334 585
R49 B.n333 B.n332 585
R50 B.n331 B.n330 585
R51 B.n329 B.n328 585
R52 B.n327 B.n326 585
R53 B.n325 B.n324 585
R54 B.n323 B.n322 585
R55 B.n321 B.n320 585
R56 B.n319 B.n318 585
R57 B.n317 B.n316 585
R58 B.n315 B.n314 585
R59 B.n313 B.n312 585
R60 B.n311 B.n310 585
R61 B.n309 B.n308 585
R62 B.n307 B.n306 585
R63 B.n304 B.n303 585
R64 B.n302 B.n301 585
R65 B.n300 B.n299 585
R66 B.n298 B.n297 585
R67 B.n296 B.n295 585
R68 B.n294 B.n293 585
R69 B.n292 B.n291 585
R70 B.n290 B.n289 585
R71 B.n288 B.n287 585
R72 B.n286 B.n285 585
R73 B.n283 B.n282 585
R74 B.n281 B.n280 585
R75 B.n279 B.n278 585
R76 B.n277 B.n276 585
R77 B.n275 B.n274 585
R78 B.n273 B.n272 585
R79 B.n271 B.n270 585
R80 B.n269 B.n268 585
R81 B.n267 B.n266 585
R82 B.n265 B.n264 585
R83 B.n263 B.n262 585
R84 B.n261 B.n260 585
R85 B.n259 B.n258 585
R86 B.n257 B.n256 585
R87 B.n255 B.n254 585
R88 B.n253 B.n252 585
R89 B.n251 B.n250 585
R90 B.n249 B.n248 585
R91 B.n247 B.n246 585
R92 B.n245 B.n244 585
R93 B.n243 B.n242 585
R94 B.n241 B.n240 585
R95 B.n239 B.n238 585
R96 B.n237 B.n236 585
R97 B.n235 B.n234 585
R98 B.n233 B.n232 585
R99 B.n231 B.n230 585
R100 B.n229 B.n228 585
R101 B.n227 B.n226 585
R102 B.n225 B.n224 585
R103 B.n223 B.n222 585
R104 B.n221 B.n220 585
R105 B.n219 B.n218 585
R106 B.n217 B.n216 585
R107 B.n215 B.n214 585
R108 B.n213 B.n212 585
R109 B.n211 B.n210 585
R110 B.n209 B.n208 585
R111 B.n207 B.n206 585
R112 B.n205 B.n204 585
R113 B.n203 B.n202 585
R114 B.n201 B.n200 585
R115 B.n199 B.n198 585
R116 B.n197 B.n196 585
R117 B.n195 B.n194 585
R118 B.n193 B.n192 585
R119 B.n191 B.n190 585
R120 B.n189 B.n188 585
R121 B.n187 B.n186 585
R122 B.n185 B.n184 585
R123 B.n183 B.n182 585
R124 B.n181 B.n180 585
R125 B.n179 B.n178 585
R126 B.n177 B.n176 585
R127 B.n175 B.n174 585
R128 B.n173 B.n172 585
R129 B.n171 B.n170 585
R130 B.n169 B.n168 585
R131 B.n167 B.n166 585
R132 B.n165 B.n164 585
R133 B.n163 B.n162 585
R134 B.n89 B.n88 585
R135 B.n1074 B.n1073 585
R136 B.n1067 B.n157 585
R137 B.n157 B.n86 585
R138 B.n1066 B.n85 585
R139 B.n1078 B.n85 585
R140 B.n1065 B.n84 585
R141 B.n1079 B.n84 585
R142 B.n1064 B.n83 585
R143 B.n1080 B.n83 585
R144 B.n1063 B.n1062 585
R145 B.n1062 B.n79 585
R146 B.n1061 B.n78 585
R147 B.n1086 B.n78 585
R148 B.n1060 B.n77 585
R149 B.n1087 B.n77 585
R150 B.n1059 B.n76 585
R151 B.n1088 B.n76 585
R152 B.n1058 B.n1057 585
R153 B.n1057 B.n75 585
R154 B.n1056 B.n71 585
R155 B.n1094 B.n71 585
R156 B.n1055 B.n70 585
R157 B.n1095 B.n70 585
R158 B.n1054 B.n69 585
R159 B.n1096 B.n69 585
R160 B.n1053 B.n1052 585
R161 B.n1052 B.n65 585
R162 B.n1051 B.n64 585
R163 B.n1102 B.n64 585
R164 B.n1050 B.n63 585
R165 B.n1103 B.n63 585
R166 B.n1049 B.n62 585
R167 B.n1104 B.n62 585
R168 B.n1048 B.n1047 585
R169 B.n1047 B.n58 585
R170 B.n1046 B.n57 585
R171 B.n1110 B.n57 585
R172 B.n1045 B.n56 585
R173 B.n1111 B.n56 585
R174 B.n1044 B.n55 585
R175 B.n1112 B.n55 585
R176 B.n1043 B.n1042 585
R177 B.n1042 B.n51 585
R178 B.n1041 B.n50 585
R179 B.n1118 B.n50 585
R180 B.n1040 B.n49 585
R181 B.n1119 B.n49 585
R182 B.n1039 B.n48 585
R183 B.n1120 B.n48 585
R184 B.n1038 B.n1037 585
R185 B.n1037 B.n44 585
R186 B.n1036 B.n43 585
R187 B.n1126 B.n43 585
R188 B.n1035 B.n42 585
R189 B.n1127 B.n42 585
R190 B.n1034 B.n41 585
R191 B.n1128 B.n41 585
R192 B.n1033 B.n1032 585
R193 B.n1032 B.n37 585
R194 B.n1031 B.n36 585
R195 B.n1134 B.n36 585
R196 B.n1030 B.n35 585
R197 B.n1135 B.n35 585
R198 B.n1029 B.n34 585
R199 B.n1136 B.n34 585
R200 B.n1028 B.n1027 585
R201 B.n1027 B.n30 585
R202 B.n1026 B.n29 585
R203 B.n1142 B.n29 585
R204 B.n1025 B.n28 585
R205 B.n1143 B.n28 585
R206 B.n1024 B.n27 585
R207 B.n1144 B.n27 585
R208 B.n1023 B.n1022 585
R209 B.n1022 B.n23 585
R210 B.n1021 B.n22 585
R211 B.n1150 B.n22 585
R212 B.n1020 B.n21 585
R213 B.n1151 B.n21 585
R214 B.n1019 B.n20 585
R215 B.n1152 B.n20 585
R216 B.n1018 B.n1017 585
R217 B.n1017 B.n19 585
R218 B.n1016 B.n15 585
R219 B.n1158 B.n15 585
R220 B.n1015 B.n14 585
R221 B.n1159 B.n14 585
R222 B.n1014 B.n13 585
R223 B.n1160 B.n13 585
R224 B.n1013 B.n1012 585
R225 B.n1012 B.n12 585
R226 B.n1011 B.n1010 585
R227 B.n1011 B.n8 585
R228 B.n1009 B.n7 585
R229 B.n1167 B.n7 585
R230 B.n1008 B.n6 585
R231 B.n1168 B.n6 585
R232 B.n1007 B.n5 585
R233 B.n1169 B.n5 585
R234 B.n1006 B.n1005 585
R235 B.n1005 B.n4 585
R236 B.n1004 B.n429 585
R237 B.n1004 B.n1003 585
R238 B.n994 B.n430 585
R239 B.n431 B.n430 585
R240 B.n996 B.n995 585
R241 B.n997 B.n996 585
R242 B.n993 B.n436 585
R243 B.n436 B.n435 585
R244 B.n992 B.n991 585
R245 B.n991 B.n990 585
R246 B.n438 B.n437 585
R247 B.n983 B.n438 585
R248 B.n982 B.n981 585
R249 B.n984 B.n982 585
R250 B.n980 B.n443 585
R251 B.n443 B.n442 585
R252 B.n979 B.n978 585
R253 B.n978 B.n977 585
R254 B.n445 B.n444 585
R255 B.n446 B.n445 585
R256 B.n970 B.n969 585
R257 B.n971 B.n970 585
R258 B.n968 B.n451 585
R259 B.n451 B.n450 585
R260 B.n967 B.n966 585
R261 B.n966 B.n965 585
R262 B.n453 B.n452 585
R263 B.n454 B.n453 585
R264 B.n958 B.n957 585
R265 B.n959 B.n958 585
R266 B.n956 B.n459 585
R267 B.n459 B.n458 585
R268 B.n955 B.n954 585
R269 B.n954 B.n953 585
R270 B.n461 B.n460 585
R271 B.n462 B.n461 585
R272 B.n946 B.n945 585
R273 B.n947 B.n946 585
R274 B.n944 B.n467 585
R275 B.n467 B.n466 585
R276 B.n943 B.n942 585
R277 B.n942 B.n941 585
R278 B.n469 B.n468 585
R279 B.n470 B.n469 585
R280 B.n934 B.n933 585
R281 B.n935 B.n934 585
R282 B.n932 B.n475 585
R283 B.n475 B.n474 585
R284 B.n931 B.n930 585
R285 B.n930 B.n929 585
R286 B.n477 B.n476 585
R287 B.n478 B.n477 585
R288 B.n922 B.n921 585
R289 B.n923 B.n922 585
R290 B.n920 B.n483 585
R291 B.n483 B.n482 585
R292 B.n919 B.n918 585
R293 B.n918 B.n917 585
R294 B.n485 B.n484 585
R295 B.n486 B.n485 585
R296 B.n910 B.n909 585
R297 B.n911 B.n910 585
R298 B.n908 B.n491 585
R299 B.n491 B.n490 585
R300 B.n907 B.n906 585
R301 B.n906 B.n905 585
R302 B.n493 B.n492 585
R303 B.n494 B.n493 585
R304 B.n898 B.n897 585
R305 B.n899 B.n898 585
R306 B.n896 B.n499 585
R307 B.n499 B.n498 585
R308 B.n895 B.n894 585
R309 B.n894 B.n893 585
R310 B.n501 B.n500 585
R311 B.n886 B.n501 585
R312 B.n885 B.n884 585
R313 B.n887 B.n885 585
R314 B.n883 B.n506 585
R315 B.n506 B.n505 585
R316 B.n882 B.n881 585
R317 B.n881 B.n880 585
R318 B.n508 B.n507 585
R319 B.n509 B.n508 585
R320 B.n873 B.n872 585
R321 B.n874 B.n873 585
R322 B.n871 B.n514 585
R323 B.n514 B.n513 585
R324 B.n870 B.n869 585
R325 B.n869 B.n868 585
R326 B.n516 B.n515 585
R327 B.n517 B.n516 585
R328 B.n864 B.n863 585
R329 B.n520 B.n519 585
R330 B.n860 B.n859 585
R331 B.n861 B.n860 585
R332 B.n858 B.n588 585
R333 B.n857 B.n856 585
R334 B.n855 B.n854 585
R335 B.n853 B.n852 585
R336 B.n851 B.n850 585
R337 B.n849 B.n848 585
R338 B.n847 B.n846 585
R339 B.n845 B.n844 585
R340 B.n843 B.n842 585
R341 B.n841 B.n840 585
R342 B.n839 B.n838 585
R343 B.n837 B.n836 585
R344 B.n835 B.n834 585
R345 B.n833 B.n832 585
R346 B.n831 B.n830 585
R347 B.n829 B.n828 585
R348 B.n827 B.n826 585
R349 B.n825 B.n824 585
R350 B.n823 B.n822 585
R351 B.n821 B.n820 585
R352 B.n819 B.n818 585
R353 B.n817 B.n816 585
R354 B.n815 B.n814 585
R355 B.n813 B.n812 585
R356 B.n811 B.n810 585
R357 B.n809 B.n808 585
R358 B.n807 B.n806 585
R359 B.n805 B.n804 585
R360 B.n803 B.n802 585
R361 B.n801 B.n800 585
R362 B.n799 B.n798 585
R363 B.n797 B.n796 585
R364 B.n795 B.n794 585
R365 B.n793 B.n792 585
R366 B.n791 B.n790 585
R367 B.n789 B.n788 585
R368 B.n787 B.n786 585
R369 B.n785 B.n784 585
R370 B.n783 B.n782 585
R371 B.n781 B.n780 585
R372 B.n779 B.n778 585
R373 B.n777 B.n776 585
R374 B.n775 B.n774 585
R375 B.n773 B.n772 585
R376 B.n771 B.n770 585
R377 B.n769 B.n768 585
R378 B.n767 B.n766 585
R379 B.n765 B.n764 585
R380 B.n763 B.n762 585
R381 B.n761 B.n760 585
R382 B.n759 B.n758 585
R383 B.n757 B.n756 585
R384 B.n755 B.n754 585
R385 B.n753 B.n752 585
R386 B.n751 B.n750 585
R387 B.n749 B.n748 585
R388 B.n747 B.n746 585
R389 B.n745 B.n744 585
R390 B.n743 B.n742 585
R391 B.n741 B.n740 585
R392 B.n739 B.n738 585
R393 B.n737 B.n736 585
R394 B.n735 B.n734 585
R395 B.n733 B.n732 585
R396 B.n731 B.n730 585
R397 B.n729 B.n728 585
R398 B.n727 B.n726 585
R399 B.n725 B.n724 585
R400 B.n723 B.n722 585
R401 B.n721 B.n720 585
R402 B.n719 B.n718 585
R403 B.n717 B.n716 585
R404 B.n715 B.n714 585
R405 B.n713 B.n712 585
R406 B.n711 B.n710 585
R407 B.n709 B.n708 585
R408 B.n707 B.n706 585
R409 B.n705 B.n704 585
R410 B.n703 B.n702 585
R411 B.n701 B.n700 585
R412 B.n699 B.n698 585
R413 B.n697 B.n696 585
R414 B.n695 B.n694 585
R415 B.n693 B.n692 585
R416 B.n691 B.n690 585
R417 B.n689 B.n688 585
R418 B.n687 B.n686 585
R419 B.n685 B.n684 585
R420 B.n683 B.n682 585
R421 B.n681 B.n680 585
R422 B.n679 B.n678 585
R423 B.n677 B.n676 585
R424 B.n675 B.n674 585
R425 B.n673 B.n672 585
R426 B.n671 B.n670 585
R427 B.n669 B.n668 585
R428 B.n667 B.n666 585
R429 B.n665 B.n664 585
R430 B.n663 B.n662 585
R431 B.n661 B.n660 585
R432 B.n659 B.n658 585
R433 B.n657 B.n656 585
R434 B.n655 B.n654 585
R435 B.n653 B.n652 585
R436 B.n651 B.n650 585
R437 B.n649 B.n648 585
R438 B.n647 B.n646 585
R439 B.n645 B.n644 585
R440 B.n643 B.n642 585
R441 B.n641 B.n640 585
R442 B.n639 B.n638 585
R443 B.n637 B.n636 585
R444 B.n635 B.n634 585
R445 B.n633 B.n632 585
R446 B.n631 B.n630 585
R447 B.n629 B.n628 585
R448 B.n627 B.n626 585
R449 B.n625 B.n624 585
R450 B.n623 B.n622 585
R451 B.n621 B.n620 585
R452 B.n619 B.n618 585
R453 B.n617 B.n616 585
R454 B.n615 B.n614 585
R455 B.n613 B.n612 585
R456 B.n611 B.n610 585
R457 B.n609 B.n608 585
R458 B.n607 B.n606 585
R459 B.n605 B.n604 585
R460 B.n603 B.n602 585
R461 B.n601 B.n600 585
R462 B.n599 B.n598 585
R463 B.n597 B.n596 585
R464 B.n595 B.n587 585
R465 B.n861 B.n587 585
R466 B.n865 B.n518 585
R467 B.n518 B.n517 585
R468 B.n867 B.n866 585
R469 B.n868 B.n867 585
R470 B.n512 B.n511 585
R471 B.n513 B.n512 585
R472 B.n876 B.n875 585
R473 B.n875 B.n874 585
R474 B.n877 B.n510 585
R475 B.n510 B.n509 585
R476 B.n879 B.n878 585
R477 B.n880 B.n879 585
R478 B.n504 B.n503 585
R479 B.n505 B.n504 585
R480 B.n889 B.n888 585
R481 B.n888 B.n887 585
R482 B.n890 B.n502 585
R483 B.n886 B.n502 585
R484 B.n892 B.n891 585
R485 B.n893 B.n892 585
R486 B.n497 B.n496 585
R487 B.n498 B.n497 585
R488 B.n901 B.n900 585
R489 B.n900 B.n899 585
R490 B.n902 B.n495 585
R491 B.n495 B.n494 585
R492 B.n904 B.n903 585
R493 B.n905 B.n904 585
R494 B.n489 B.n488 585
R495 B.n490 B.n489 585
R496 B.n913 B.n912 585
R497 B.n912 B.n911 585
R498 B.n914 B.n487 585
R499 B.n487 B.n486 585
R500 B.n916 B.n915 585
R501 B.n917 B.n916 585
R502 B.n481 B.n480 585
R503 B.n482 B.n481 585
R504 B.n925 B.n924 585
R505 B.n924 B.n923 585
R506 B.n926 B.n479 585
R507 B.n479 B.n478 585
R508 B.n928 B.n927 585
R509 B.n929 B.n928 585
R510 B.n473 B.n472 585
R511 B.n474 B.n473 585
R512 B.n937 B.n936 585
R513 B.n936 B.n935 585
R514 B.n938 B.n471 585
R515 B.n471 B.n470 585
R516 B.n940 B.n939 585
R517 B.n941 B.n940 585
R518 B.n465 B.n464 585
R519 B.n466 B.n465 585
R520 B.n949 B.n948 585
R521 B.n948 B.n947 585
R522 B.n950 B.n463 585
R523 B.n463 B.n462 585
R524 B.n952 B.n951 585
R525 B.n953 B.n952 585
R526 B.n457 B.n456 585
R527 B.n458 B.n457 585
R528 B.n961 B.n960 585
R529 B.n960 B.n959 585
R530 B.n962 B.n455 585
R531 B.n455 B.n454 585
R532 B.n964 B.n963 585
R533 B.n965 B.n964 585
R534 B.n449 B.n448 585
R535 B.n450 B.n449 585
R536 B.n973 B.n972 585
R537 B.n972 B.n971 585
R538 B.n974 B.n447 585
R539 B.n447 B.n446 585
R540 B.n976 B.n975 585
R541 B.n977 B.n976 585
R542 B.n441 B.n440 585
R543 B.n442 B.n441 585
R544 B.n986 B.n985 585
R545 B.n985 B.n984 585
R546 B.n987 B.n439 585
R547 B.n983 B.n439 585
R548 B.n989 B.n988 585
R549 B.n990 B.n989 585
R550 B.n434 B.n433 585
R551 B.n435 B.n434 585
R552 B.n999 B.n998 585
R553 B.n998 B.n997 585
R554 B.n1000 B.n432 585
R555 B.n432 B.n431 585
R556 B.n1002 B.n1001 585
R557 B.n1003 B.n1002 585
R558 B.n3 B.n0 585
R559 B.n4 B.n3 585
R560 B.n1166 B.n1 585
R561 B.n1167 B.n1166 585
R562 B.n1165 B.n1164 585
R563 B.n1165 B.n8 585
R564 B.n1163 B.n9 585
R565 B.n12 B.n9 585
R566 B.n1162 B.n1161 585
R567 B.n1161 B.n1160 585
R568 B.n11 B.n10 585
R569 B.n1159 B.n11 585
R570 B.n1157 B.n1156 585
R571 B.n1158 B.n1157 585
R572 B.n1155 B.n16 585
R573 B.n19 B.n16 585
R574 B.n1154 B.n1153 585
R575 B.n1153 B.n1152 585
R576 B.n18 B.n17 585
R577 B.n1151 B.n18 585
R578 B.n1149 B.n1148 585
R579 B.n1150 B.n1149 585
R580 B.n1147 B.n24 585
R581 B.n24 B.n23 585
R582 B.n1146 B.n1145 585
R583 B.n1145 B.n1144 585
R584 B.n26 B.n25 585
R585 B.n1143 B.n26 585
R586 B.n1141 B.n1140 585
R587 B.n1142 B.n1141 585
R588 B.n1139 B.n31 585
R589 B.n31 B.n30 585
R590 B.n1138 B.n1137 585
R591 B.n1137 B.n1136 585
R592 B.n33 B.n32 585
R593 B.n1135 B.n33 585
R594 B.n1133 B.n1132 585
R595 B.n1134 B.n1133 585
R596 B.n1131 B.n38 585
R597 B.n38 B.n37 585
R598 B.n1130 B.n1129 585
R599 B.n1129 B.n1128 585
R600 B.n40 B.n39 585
R601 B.n1127 B.n40 585
R602 B.n1125 B.n1124 585
R603 B.n1126 B.n1125 585
R604 B.n1123 B.n45 585
R605 B.n45 B.n44 585
R606 B.n1122 B.n1121 585
R607 B.n1121 B.n1120 585
R608 B.n47 B.n46 585
R609 B.n1119 B.n47 585
R610 B.n1117 B.n1116 585
R611 B.n1118 B.n1117 585
R612 B.n1115 B.n52 585
R613 B.n52 B.n51 585
R614 B.n1114 B.n1113 585
R615 B.n1113 B.n1112 585
R616 B.n54 B.n53 585
R617 B.n1111 B.n54 585
R618 B.n1109 B.n1108 585
R619 B.n1110 B.n1109 585
R620 B.n1107 B.n59 585
R621 B.n59 B.n58 585
R622 B.n1106 B.n1105 585
R623 B.n1105 B.n1104 585
R624 B.n61 B.n60 585
R625 B.n1103 B.n61 585
R626 B.n1101 B.n1100 585
R627 B.n1102 B.n1101 585
R628 B.n1099 B.n66 585
R629 B.n66 B.n65 585
R630 B.n1098 B.n1097 585
R631 B.n1097 B.n1096 585
R632 B.n68 B.n67 585
R633 B.n1095 B.n68 585
R634 B.n1093 B.n1092 585
R635 B.n1094 B.n1093 585
R636 B.n1091 B.n72 585
R637 B.n75 B.n72 585
R638 B.n1090 B.n1089 585
R639 B.n1089 B.n1088 585
R640 B.n74 B.n73 585
R641 B.n1087 B.n74 585
R642 B.n1085 B.n1084 585
R643 B.n1086 B.n1085 585
R644 B.n1083 B.n80 585
R645 B.n80 B.n79 585
R646 B.n1082 B.n1081 585
R647 B.n1081 B.n1080 585
R648 B.n82 B.n81 585
R649 B.n1079 B.n82 585
R650 B.n1077 B.n1076 585
R651 B.n1078 B.n1077 585
R652 B.n1075 B.n87 585
R653 B.n87 B.n86 585
R654 B.n1170 B.n1169 585
R655 B.n1168 B.n2 585
R656 B.n1073 B.n87 478.086
R657 B.n1069 B.n157 478.086
R658 B.n587 B.n516 478.086
R659 B.n863 B.n518 478.086
R660 B.n160 B.t16 363.361
R661 B.n158 B.t5 363.361
R662 B.n592 B.t13 363.361
R663 B.n589 B.t9 363.361
R664 B.n1071 B.n1070 256.663
R665 B.n1071 B.n155 256.663
R666 B.n1071 B.n154 256.663
R667 B.n1071 B.n153 256.663
R668 B.n1071 B.n152 256.663
R669 B.n1071 B.n151 256.663
R670 B.n1071 B.n150 256.663
R671 B.n1071 B.n149 256.663
R672 B.n1071 B.n148 256.663
R673 B.n1071 B.n147 256.663
R674 B.n1071 B.n146 256.663
R675 B.n1071 B.n145 256.663
R676 B.n1071 B.n144 256.663
R677 B.n1071 B.n143 256.663
R678 B.n1071 B.n142 256.663
R679 B.n1071 B.n141 256.663
R680 B.n1071 B.n140 256.663
R681 B.n1071 B.n139 256.663
R682 B.n1071 B.n138 256.663
R683 B.n1071 B.n137 256.663
R684 B.n1071 B.n136 256.663
R685 B.n1071 B.n135 256.663
R686 B.n1071 B.n134 256.663
R687 B.n1071 B.n133 256.663
R688 B.n1071 B.n132 256.663
R689 B.n1071 B.n131 256.663
R690 B.n1071 B.n130 256.663
R691 B.n1071 B.n129 256.663
R692 B.n1071 B.n128 256.663
R693 B.n1071 B.n127 256.663
R694 B.n1071 B.n126 256.663
R695 B.n1071 B.n125 256.663
R696 B.n1071 B.n124 256.663
R697 B.n1071 B.n123 256.663
R698 B.n1071 B.n122 256.663
R699 B.n1071 B.n121 256.663
R700 B.n1071 B.n120 256.663
R701 B.n1071 B.n119 256.663
R702 B.n1071 B.n118 256.663
R703 B.n1071 B.n117 256.663
R704 B.n1071 B.n116 256.663
R705 B.n1071 B.n115 256.663
R706 B.n1071 B.n114 256.663
R707 B.n1071 B.n113 256.663
R708 B.n1071 B.n112 256.663
R709 B.n1071 B.n111 256.663
R710 B.n1071 B.n110 256.663
R711 B.n1071 B.n109 256.663
R712 B.n1071 B.n108 256.663
R713 B.n1071 B.n107 256.663
R714 B.n1071 B.n106 256.663
R715 B.n1071 B.n105 256.663
R716 B.n1071 B.n104 256.663
R717 B.n1071 B.n103 256.663
R718 B.n1071 B.n102 256.663
R719 B.n1071 B.n101 256.663
R720 B.n1071 B.n100 256.663
R721 B.n1071 B.n99 256.663
R722 B.n1071 B.n98 256.663
R723 B.n1071 B.n97 256.663
R724 B.n1071 B.n96 256.663
R725 B.n1071 B.n95 256.663
R726 B.n1071 B.n94 256.663
R727 B.n1071 B.n93 256.663
R728 B.n1071 B.n92 256.663
R729 B.n1071 B.n91 256.663
R730 B.n1071 B.n90 256.663
R731 B.n1072 B.n1071 256.663
R732 B.n862 B.n861 256.663
R733 B.n861 B.n521 256.663
R734 B.n861 B.n522 256.663
R735 B.n861 B.n523 256.663
R736 B.n861 B.n524 256.663
R737 B.n861 B.n525 256.663
R738 B.n861 B.n526 256.663
R739 B.n861 B.n527 256.663
R740 B.n861 B.n528 256.663
R741 B.n861 B.n529 256.663
R742 B.n861 B.n530 256.663
R743 B.n861 B.n531 256.663
R744 B.n861 B.n532 256.663
R745 B.n861 B.n533 256.663
R746 B.n861 B.n534 256.663
R747 B.n861 B.n535 256.663
R748 B.n861 B.n536 256.663
R749 B.n861 B.n537 256.663
R750 B.n861 B.n538 256.663
R751 B.n861 B.n539 256.663
R752 B.n861 B.n540 256.663
R753 B.n861 B.n541 256.663
R754 B.n861 B.n542 256.663
R755 B.n861 B.n543 256.663
R756 B.n861 B.n544 256.663
R757 B.n861 B.n545 256.663
R758 B.n861 B.n546 256.663
R759 B.n861 B.n547 256.663
R760 B.n861 B.n548 256.663
R761 B.n861 B.n549 256.663
R762 B.n861 B.n550 256.663
R763 B.n861 B.n551 256.663
R764 B.n861 B.n552 256.663
R765 B.n861 B.n553 256.663
R766 B.n861 B.n554 256.663
R767 B.n861 B.n555 256.663
R768 B.n861 B.n556 256.663
R769 B.n861 B.n557 256.663
R770 B.n861 B.n558 256.663
R771 B.n861 B.n559 256.663
R772 B.n861 B.n560 256.663
R773 B.n861 B.n561 256.663
R774 B.n861 B.n562 256.663
R775 B.n861 B.n563 256.663
R776 B.n861 B.n564 256.663
R777 B.n861 B.n565 256.663
R778 B.n861 B.n566 256.663
R779 B.n861 B.n567 256.663
R780 B.n861 B.n568 256.663
R781 B.n861 B.n569 256.663
R782 B.n861 B.n570 256.663
R783 B.n861 B.n571 256.663
R784 B.n861 B.n572 256.663
R785 B.n861 B.n573 256.663
R786 B.n861 B.n574 256.663
R787 B.n861 B.n575 256.663
R788 B.n861 B.n576 256.663
R789 B.n861 B.n577 256.663
R790 B.n861 B.n578 256.663
R791 B.n861 B.n579 256.663
R792 B.n861 B.n580 256.663
R793 B.n861 B.n581 256.663
R794 B.n861 B.n582 256.663
R795 B.n861 B.n583 256.663
R796 B.n861 B.n584 256.663
R797 B.n861 B.n585 256.663
R798 B.n861 B.n586 256.663
R799 B.n1172 B.n1171 256.663
R800 B.n162 B.n89 163.367
R801 B.n166 B.n165 163.367
R802 B.n170 B.n169 163.367
R803 B.n174 B.n173 163.367
R804 B.n178 B.n177 163.367
R805 B.n182 B.n181 163.367
R806 B.n186 B.n185 163.367
R807 B.n190 B.n189 163.367
R808 B.n194 B.n193 163.367
R809 B.n198 B.n197 163.367
R810 B.n202 B.n201 163.367
R811 B.n206 B.n205 163.367
R812 B.n210 B.n209 163.367
R813 B.n214 B.n213 163.367
R814 B.n218 B.n217 163.367
R815 B.n222 B.n221 163.367
R816 B.n226 B.n225 163.367
R817 B.n230 B.n229 163.367
R818 B.n234 B.n233 163.367
R819 B.n238 B.n237 163.367
R820 B.n242 B.n241 163.367
R821 B.n246 B.n245 163.367
R822 B.n250 B.n249 163.367
R823 B.n254 B.n253 163.367
R824 B.n258 B.n257 163.367
R825 B.n262 B.n261 163.367
R826 B.n266 B.n265 163.367
R827 B.n270 B.n269 163.367
R828 B.n274 B.n273 163.367
R829 B.n278 B.n277 163.367
R830 B.n282 B.n281 163.367
R831 B.n287 B.n286 163.367
R832 B.n291 B.n290 163.367
R833 B.n295 B.n294 163.367
R834 B.n299 B.n298 163.367
R835 B.n303 B.n302 163.367
R836 B.n308 B.n307 163.367
R837 B.n312 B.n311 163.367
R838 B.n316 B.n315 163.367
R839 B.n320 B.n319 163.367
R840 B.n324 B.n323 163.367
R841 B.n328 B.n327 163.367
R842 B.n332 B.n331 163.367
R843 B.n336 B.n335 163.367
R844 B.n340 B.n339 163.367
R845 B.n344 B.n343 163.367
R846 B.n348 B.n347 163.367
R847 B.n352 B.n351 163.367
R848 B.n356 B.n355 163.367
R849 B.n360 B.n359 163.367
R850 B.n364 B.n363 163.367
R851 B.n368 B.n367 163.367
R852 B.n372 B.n371 163.367
R853 B.n376 B.n375 163.367
R854 B.n380 B.n379 163.367
R855 B.n384 B.n383 163.367
R856 B.n388 B.n387 163.367
R857 B.n392 B.n391 163.367
R858 B.n396 B.n395 163.367
R859 B.n400 B.n399 163.367
R860 B.n404 B.n403 163.367
R861 B.n408 B.n407 163.367
R862 B.n412 B.n411 163.367
R863 B.n416 B.n415 163.367
R864 B.n420 B.n419 163.367
R865 B.n424 B.n423 163.367
R866 B.n426 B.n156 163.367
R867 B.n869 B.n516 163.367
R868 B.n869 B.n514 163.367
R869 B.n873 B.n514 163.367
R870 B.n873 B.n508 163.367
R871 B.n881 B.n508 163.367
R872 B.n881 B.n506 163.367
R873 B.n885 B.n506 163.367
R874 B.n885 B.n501 163.367
R875 B.n894 B.n501 163.367
R876 B.n894 B.n499 163.367
R877 B.n898 B.n499 163.367
R878 B.n898 B.n493 163.367
R879 B.n906 B.n493 163.367
R880 B.n906 B.n491 163.367
R881 B.n910 B.n491 163.367
R882 B.n910 B.n485 163.367
R883 B.n918 B.n485 163.367
R884 B.n918 B.n483 163.367
R885 B.n922 B.n483 163.367
R886 B.n922 B.n477 163.367
R887 B.n930 B.n477 163.367
R888 B.n930 B.n475 163.367
R889 B.n934 B.n475 163.367
R890 B.n934 B.n469 163.367
R891 B.n942 B.n469 163.367
R892 B.n942 B.n467 163.367
R893 B.n946 B.n467 163.367
R894 B.n946 B.n461 163.367
R895 B.n954 B.n461 163.367
R896 B.n954 B.n459 163.367
R897 B.n958 B.n459 163.367
R898 B.n958 B.n453 163.367
R899 B.n966 B.n453 163.367
R900 B.n966 B.n451 163.367
R901 B.n970 B.n451 163.367
R902 B.n970 B.n445 163.367
R903 B.n978 B.n445 163.367
R904 B.n978 B.n443 163.367
R905 B.n982 B.n443 163.367
R906 B.n982 B.n438 163.367
R907 B.n991 B.n438 163.367
R908 B.n991 B.n436 163.367
R909 B.n996 B.n436 163.367
R910 B.n996 B.n430 163.367
R911 B.n1004 B.n430 163.367
R912 B.n1005 B.n1004 163.367
R913 B.n1005 B.n5 163.367
R914 B.n6 B.n5 163.367
R915 B.n7 B.n6 163.367
R916 B.n1011 B.n7 163.367
R917 B.n1012 B.n1011 163.367
R918 B.n1012 B.n13 163.367
R919 B.n14 B.n13 163.367
R920 B.n15 B.n14 163.367
R921 B.n1017 B.n15 163.367
R922 B.n1017 B.n20 163.367
R923 B.n21 B.n20 163.367
R924 B.n22 B.n21 163.367
R925 B.n1022 B.n22 163.367
R926 B.n1022 B.n27 163.367
R927 B.n28 B.n27 163.367
R928 B.n29 B.n28 163.367
R929 B.n1027 B.n29 163.367
R930 B.n1027 B.n34 163.367
R931 B.n35 B.n34 163.367
R932 B.n36 B.n35 163.367
R933 B.n1032 B.n36 163.367
R934 B.n1032 B.n41 163.367
R935 B.n42 B.n41 163.367
R936 B.n43 B.n42 163.367
R937 B.n1037 B.n43 163.367
R938 B.n1037 B.n48 163.367
R939 B.n49 B.n48 163.367
R940 B.n50 B.n49 163.367
R941 B.n1042 B.n50 163.367
R942 B.n1042 B.n55 163.367
R943 B.n56 B.n55 163.367
R944 B.n57 B.n56 163.367
R945 B.n1047 B.n57 163.367
R946 B.n1047 B.n62 163.367
R947 B.n63 B.n62 163.367
R948 B.n64 B.n63 163.367
R949 B.n1052 B.n64 163.367
R950 B.n1052 B.n69 163.367
R951 B.n70 B.n69 163.367
R952 B.n71 B.n70 163.367
R953 B.n1057 B.n71 163.367
R954 B.n1057 B.n76 163.367
R955 B.n77 B.n76 163.367
R956 B.n78 B.n77 163.367
R957 B.n1062 B.n78 163.367
R958 B.n1062 B.n83 163.367
R959 B.n84 B.n83 163.367
R960 B.n85 B.n84 163.367
R961 B.n157 B.n85 163.367
R962 B.n860 B.n520 163.367
R963 B.n860 B.n588 163.367
R964 B.n856 B.n855 163.367
R965 B.n852 B.n851 163.367
R966 B.n848 B.n847 163.367
R967 B.n844 B.n843 163.367
R968 B.n840 B.n839 163.367
R969 B.n836 B.n835 163.367
R970 B.n832 B.n831 163.367
R971 B.n828 B.n827 163.367
R972 B.n824 B.n823 163.367
R973 B.n820 B.n819 163.367
R974 B.n816 B.n815 163.367
R975 B.n812 B.n811 163.367
R976 B.n808 B.n807 163.367
R977 B.n804 B.n803 163.367
R978 B.n800 B.n799 163.367
R979 B.n796 B.n795 163.367
R980 B.n792 B.n791 163.367
R981 B.n788 B.n787 163.367
R982 B.n784 B.n783 163.367
R983 B.n780 B.n779 163.367
R984 B.n776 B.n775 163.367
R985 B.n772 B.n771 163.367
R986 B.n768 B.n767 163.367
R987 B.n764 B.n763 163.367
R988 B.n760 B.n759 163.367
R989 B.n756 B.n755 163.367
R990 B.n752 B.n751 163.367
R991 B.n748 B.n747 163.367
R992 B.n744 B.n743 163.367
R993 B.n740 B.n739 163.367
R994 B.n736 B.n735 163.367
R995 B.n732 B.n731 163.367
R996 B.n728 B.n727 163.367
R997 B.n724 B.n723 163.367
R998 B.n720 B.n719 163.367
R999 B.n716 B.n715 163.367
R1000 B.n712 B.n711 163.367
R1001 B.n708 B.n707 163.367
R1002 B.n704 B.n703 163.367
R1003 B.n700 B.n699 163.367
R1004 B.n696 B.n695 163.367
R1005 B.n692 B.n691 163.367
R1006 B.n688 B.n687 163.367
R1007 B.n684 B.n683 163.367
R1008 B.n680 B.n679 163.367
R1009 B.n676 B.n675 163.367
R1010 B.n672 B.n671 163.367
R1011 B.n668 B.n667 163.367
R1012 B.n664 B.n663 163.367
R1013 B.n660 B.n659 163.367
R1014 B.n656 B.n655 163.367
R1015 B.n652 B.n651 163.367
R1016 B.n648 B.n647 163.367
R1017 B.n644 B.n643 163.367
R1018 B.n640 B.n639 163.367
R1019 B.n636 B.n635 163.367
R1020 B.n632 B.n631 163.367
R1021 B.n628 B.n627 163.367
R1022 B.n624 B.n623 163.367
R1023 B.n620 B.n619 163.367
R1024 B.n616 B.n615 163.367
R1025 B.n612 B.n611 163.367
R1026 B.n608 B.n607 163.367
R1027 B.n604 B.n603 163.367
R1028 B.n600 B.n599 163.367
R1029 B.n596 B.n587 163.367
R1030 B.n867 B.n518 163.367
R1031 B.n867 B.n512 163.367
R1032 B.n875 B.n512 163.367
R1033 B.n875 B.n510 163.367
R1034 B.n879 B.n510 163.367
R1035 B.n879 B.n504 163.367
R1036 B.n888 B.n504 163.367
R1037 B.n888 B.n502 163.367
R1038 B.n892 B.n502 163.367
R1039 B.n892 B.n497 163.367
R1040 B.n900 B.n497 163.367
R1041 B.n900 B.n495 163.367
R1042 B.n904 B.n495 163.367
R1043 B.n904 B.n489 163.367
R1044 B.n912 B.n489 163.367
R1045 B.n912 B.n487 163.367
R1046 B.n916 B.n487 163.367
R1047 B.n916 B.n481 163.367
R1048 B.n924 B.n481 163.367
R1049 B.n924 B.n479 163.367
R1050 B.n928 B.n479 163.367
R1051 B.n928 B.n473 163.367
R1052 B.n936 B.n473 163.367
R1053 B.n936 B.n471 163.367
R1054 B.n940 B.n471 163.367
R1055 B.n940 B.n465 163.367
R1056 B.n948 B.n465 163.367
R1057 B.n948 B.n463 163.367
R1058 B.n952 B.n463 163.367
R1059 B.n952 B.n457 163.367
R1060 B.n960 B.n457 163.367
R1061 B.n960 B.n455 163.367
R1062 B.n964 B.n455 163.367
R1063 B.n964 B.n449 163.367
R1064 B.n972 B.n449 163.367
R1065 B.n972 B.n447 163.367
R1066 B.n976 B.n447 163.367
R1067 B.n976 B.n441 163.367
R1068 B.n985 B.n441 163.367
R1069 B.n985 B.n439 163.367
R1070 B.n989 B.n439 163.367
R1071 B.n989 B.n434 163.367
R1072 B.n998 B.n434 163.367
R1073 B.n998 B.n432 163.367
R1074 B.n1002 B.n432 163.367
R1075 B.n1002 B.n3 163.367
R1076 B.n1170 B.n3 163.367
R1077 B.n1166 B.n2 163.367
R1078 B.n1166 B.n1165 163.367
R1079 B.n1165 B.n9 163.367
R1080 B.n1161 B.n9 163.367
R1081 B.n1161 B.n11 163.367
R1082 B.n1157 B.n11 163.367
R1083 B.n1157 B.n16 163.367
R1084 B.n1153 B.n16 163.367
R1085 B.n1153 B.n18 163.367
R1086 B.n1149 B.n18 163.367
R1087 B.n1149 B.n24 163.367
R1088 B.n1145 B.n24 163.367
R1089 B.n1145 B.n26 163.367
R1090 B.n1141 B.n26 163.367
R1091 B.n1141 B.n31 163.367
R1092 B.n1137 B.n31 163.367
R1093 B.n1137 B.n33 163.367
R1094 B.n1133 B.n33 163.367
R1095 B.n1133 B.n38 163.367
R1096 B.n1129 B.n38 163.367
R1097 B.n1129 B.n40 163.367
R1098 B.n1125 B.n40 163.367
R1099 B.n1125 B.n45 163.367
R1100 B.n1121 B.n45 163.367
R1101 B.n1121 B.n47 163.367
R1102 B.n1117 B.n47 163.367
R1103 B.n1117 B.n52 163.367
R1104 B.n1113 B.n52 163.367
R1105 B.n1113 B.n54 163.367
R1106 B.n1109 B.n54 163.367
R1107 B.n1109 B.n59 163.367
R1108 B.n1105 B.n59 163.367
R1109 B.n1105 B.n61 163.367
R1110 B.n1101 B.n61 163.367
R1111 B.n1101 B.n66 163.367
R1112 B.n1097 B.n66 163.367
R1113 B.n1097 B.n68 163.367
R1114 B.n1093 B.n68 163.367
R1115 B.n1093 B.n72 163.367
R1116 B.n1089 B.n72 163.367
R1117 B.n1089 B.n74 163.367
R1118 B.n1085 B.n74 163.367
R1119 B.n1085 B.n80 163.367
R1120 B.n1081 B.n80 163.367
R1121 B.n1081 B.n82 163.367
R1122 B.n1077 B.n82 163.367
R1123 B.n1077 B.n87 163.367
R1124 B.n158 B.t7 137.575
R1125 B.n592 B.t15 137.575
R1126 B.n160 B.t17 137.548
R1127 B.n589 B.t12 137.548
R1128 B.n159 B.t8 72.7989
R1129 B.n593 B.t14 72.7989
R1130 B.n161 B.t18 72.7732
R1131 B.n590 B.t11 72.7732
R1132 B.n1073 B.n1072 71.676
R1133 B.n162 B.n90 71.676
R1134 B.n166 B.n91 71.676
R1135 B.n170 B.n92 71.676
R1136 B.n174 B.n93 71.676
R1137 B.n178 B.n94 71.676
R1138 B.n182 B.n95 71.676
R1139 B.n186 B.n96 71.676
R1140 B.n190 B.n97 71.676
R1141 B.n194 B.n98 71.676
R1142 B.n198 B.n99 71.676
R1143 B.n202 B.n100 71.676
R1144 B.n206 B.n101 71.676
R1145 B.n210 B.n102 71.676
R1146 B.n214 B.n103 71.676
R1147 B.n218 B.n104 71.676
R1148 B.n222 B.n105 71.676
R1149 B.n226 B.n106 71.676
R1150 B.n230 B.n107 71.676
R1151 B.n234 B.n108 71.676
R1152 B.n238 B.n109 71.676
R1153 B.n242 B.n110 71.676
R1154 B.n246 B.n111 71.676
R1155 B.n250 B.n112 71.676
R1156 B.n254 B.n113 71.676
R1157 B.n258 B.n114 71.676
R1158 B.n262 B.n115 71.676
R1159 B.n266 B.n116 71.676
R1160 B.n270 B.n117 71.676
R1161 B.n274 B.n118 71.676
R1162 B.n278 B.n119 71.676
R1163 B.n282 B.n120 71.676
R1164 B.n287 B.n121 71.676
R1165 B.n291 B.n122 71.676
R1166 B.n295 B.n123 71.676
R1167 B.n299 B.n124 71.676
R1168 B.n303 B.n125 71.676
R1169 B.n308 B.n126 71.676
R1170 B.n312 B.n127 71.676
R1171 B.n316 B.n128 71.676
R1172 B.n320 B.n129 71.676
R1173 B.n324 B.n130 71.676
R1174 B.n328 B.n131 71.676
R1175 B.n332 B.n132 71.676
R1176 B.n336 B.n133 71.676
R1177 B.n340 B.n134 71.676
R1178 B.n344 B.n135 71.676
R1179 B.n348 B.n136 71.676
R1180 B.n352 B.n137 71.676
R1181 B.n356 B.n138 71.676
R1182 B.n360 B.n139 71.676
R1183 B.n364 B.n140 71.676
R1184 B.n368 B.n141 71.676
R1185 B.n372 B.n142 71.676
R1186 B.n376 B.n143 71.676
R1187 B.n380 B.n144 71.676
R1188 B.n384 B.n145 71.676
R1189 B.n388 B.n146 71.676
R1190 B.n392 B.n147 71.676
R1191 B.n396 B.n148 71.676
R1192 B.n400 B.n149 71.676
R1193 B.n404 B.n150 71.676
R1194 B.n408 B.n151 71.676
R1195 B.n412 B.n152 71.676
R1196 B.n416 B.n153 71.676
R1197 B.n420 B.n154 71.676
R1198 B.n424 B.n155 71.676
R1199 B.n1070 B.n156 71.676
R1200 B.n1070 B.n1069 71.676
R1201 B.n426 B.n155 71.676
R1202 B.n423 B.n154 71.676
R1203 B.n419 B.n153 71.676
R1204 B.n415 B.n152 71.676
R1205 B.n411 B.n151 71.676
R1206 B.n407 B.n150 71.676
R1207 B.n403 B.n149 71.676
R1208 B.n399 B.n148 71.676
R1209 B.n395 B.n147 71.676
R1210 B.n391 B.n146 71.676
R1211 B.n387 B.n145 71.676
R1212 B.n383 B.n144 71.676
R1213 B.n379 B.n143 71.676
R1214 B.n375 B.n142 71.676
R1215 B.n371 B.n141 71.676
R1216 B.n367 B.n140 71.676
R1217 B.n363 B.n139 71.676
R1218 B.n359 B.n138 71.676
R1219 B.n355 B.n137 71.676
R1220 B.n351 B.n136 71.676
R1221 B.n347 B.n135 71.676
R1222 B.n343 B.n134 71.676
R1223 B.n339 B.n133 71.676
R1224 B.n335 B.n132 71.676
R1225 B.n331 B.n131 71.676
R1226 B.n327 B.n130 71.676
R1227 B.n323 B.n129 71.676
R1228 B.n319 B.n128 71.676
R1229 B.n315 B.n127 71.676
R1230 B.n311 B.n126 71.676
R1231 B.n307 B.n125 71.676
R1232 B.n302 B.n124 71.676
R1233 B.n298 B.n123 71.676
R1234 B.n294 B.n122 71.676
R1235 B.n290 B.n121 71.676
R1236 B.n286 B.n120 71.676
R1237 B.n281 B.n119 71.676
R1238 B.n277 B.n118 71.676
R1239 B.n273 B.n117 71.676
R1240 B.n269 B.n116 71.676
R1241 B.n265 B.n115 71.676
R1242 B.n261 B.n114 71.676
R1243 B.n257 B.n113 71.676
R1244 B.n253 B.n112 71.676
R1245 B.n249 B.n111 71.676
R1246 B.n245 B.n110 71.676
R1247 B.n241 B.n109 71.676
R1248 B.n237 B.n108 71.676
R1249 B.n233 B.n107 71.676
R1250 B.n229 B.n106 71.676
R1251 B.n225 B.n105 71.676
R1252 B.n221 B.n104 71.676
R1253 B.n217 B.n103 71.676
R1254 B.n213 B.n102 71.676
R1255 B.n209 B.n101 71.676
R1256 B.n205 B.n100 71.676
R1257 B.n201 B.n99 71.676
R1258 B.n197 B.n98 71.676
R1259 B.n193 B.n97 71.676
R1260 B.n189 B.n96 71.676
R1261 B.n185 B.n95 71.676
R1262 B.n181 B.n94 71.676
R1263 B.n177 B.n93 71.676
R1264 B.n173 B.n92 71.676
R1265 B.n169 B.n91 71.676
R1266 B.n165 B.n90 71.676
R1267 B.n1072 B.n89 71.676
R1268 B.n863 B.n862 71.676
R1269 B.n588 B.n521 71.676
R1270 B.n855 B.n522 71.676
R1271 B.n851 B.n523 71.676
R1272 B.n847 B.n524 71.676
R1273 B.n843 B.n525 71.676
R1274 B.n839 B.n526 71.676
R1275 B.n835 B.n527 71.676
R1276 B.n831 B.n528 71.676
R1277 B.n827 B.n529 71.676
R1278 B.n823 B.n530 71.676
R1279 B.n819 B.n531 71.676
R1280 B.n815 B.n532 71.676
R1281 B.n811 B.n533 71.676
R1282 B.n807 B.n534 71.676
R1283 B.n803 B.n535 71.676
R1284 B.n799 B.n536 71.676
R1285 B.n795 B.n537 71.676
R1286 B.n791 B.n538 71.676
R1287 B.n787 B.n539 71.676
R1288 B.n783 B.n540 71.676
R1289 B.n779 B.n541 71.676
R1290 B.n775 B.n542 71.676
R1291 B.n771 B.n543 71.676
R1292 B.n767 B.n544 71.676
R1293 B.n763 B.n545 71.676
R1294 B.n759 B.n546 71.676
R1295 B.n755 B.n547 71.676
R1296 B.n751 B.n548 71.676
R1297 B.n747 B.n549 71.676
R1298 B.n743 B.n550 71.676
R1299 B.n739 B.n551 71.676
R1300 B.n735 B.n552 71.676
R1301 B.n731 B.n553 71.676
R1302 B.n727 B.n554 71.676
R1303 B.n723 B.n555 71.676
R1304 B.n719 B.n556 71.676
R1305 B.n715 B.n557 71.676
R1306 B.n711 B.n558 71.676
R1307 B.n707 B.n559 71.676
R1308 B.n703 B.n560 71.676
R1309 B.n699 B.n561 71.676
R1310 B.n695 B.n562 71.676
R1311 B.n691 B.n563 71.676
R1312 B.n687 B.n564 71.676
R1313 B.n683 B.n565 71.676
R1314 B.n679 B.n566 71.676
R1315 B.n675 B.n567 71.676
R1316 B.n671 B.n568 71.676
R1317 B.n667 B.n569 71.676
R1318 B.n663 B.n570 71.676
R1319 B.n659 B.n571 71.676
R1320 B.n655 B.n572 71.676
R1321 B.n651 B.n573 71.676
R1322 B.n647 B.n574 71.676
R1323 B.n643 B.n575 71.676
R1324 B.n639 B.n576 71.676
R1325 B.n635 B.n577 71.676
R1326 B.n631 B.n578 71.676
R1327 B.n627 B.n579 71.676
R1328 B.n623 B.n580 71.676
R1329 B.n619 B.n581 71.676
R1330 B.n615 B.n582 71.676
R1331 B.n611 B.n583 71.676
R1332 B.n607 B.n584 71.676
R1333 B.n603 B.n585 71.676
R1334 B.n599 B.n586 71.676
R1335 B.n862 B.n520 71.676
R1336 B.n856 B.n521 71.676
R1337 B.n852 B.n522 71.676
R1338 B.n848 B.n523 71.676
R1339 B.n844 B.n524 71.676
R1340 B.n840 B.n525 71.676
R1341 B.n836 B.n526 71.676
R1342 B.n832 B.n527 71.676
R1343 B.n828 B.n528 71.676
R1344 B.n824 B.n529 71.676
R1345 B.n820 B.n530 71.676
R1346 B.n816 B.n531 71.676
R1347 B.n812 B.n532 71.676
R1348 B.n808 B.n533 71.676
R1349 B.n804 B.n534 71.676
R1350 B.n800 B.n535 71.676
R1351 B.n796 B.n536 71.676
R1352 B.n792 B.n537 71.676
R1353 B.n788 B.n538 71.676
R1354 B.n784 B.n539 71.676
R1355 B.n780 B.n540 71.676
R1356 B.n776 B.n541 71.676
R1357 B.n772 B.n542 71.676
R1358 B.n768 B.n543 71.676
R1359 B.n764 B.n544 71.676
R1360 B.n760 B.n545 71.676
R1361 B.n756 B.n546 71.676
R1362 B.n752 B.n547 71.676
R1363 B.n748 B.n548 71.676
R1364 B.n744 B.n549 71.676
R1365 B.n740 B.n550 71.676
R1366 B.n736 B.n551 71.676
R1367 B.n732 B.n552 71.676
R1368 B.n728 B.n553 71.676
R1369 B.n724 B.n554 71.676
R1370 B.n720 B.n555 71.676
R1371 B.n716 B.n556 71.676
R1372 B.n712 B.n557 71.676
R1373 B.n708 B.n558 71.676
R1374 B.n704 B.n559 71.676
R1375 B.n700 B.n560 71.676
R1376 B.n696 B.n561 71.676
R1377 B.n692 B.n562 71.676
R1378 B.n688 B.n563 71.676
R1379 B.n684 B.n564 71.676
R1380 B.n680 B.n565 71.676
R1381 B.n676 B.n566 71.676
R1382 B.n672 B.n567 71.676
R1383 B.n668 B.n568 71.676
R1384 B.n664 B.n569 71.676
R1385 B.n660 B.n570 71.676
R1386 B.n656 B.n571 71.676
R1387 B.n652 B.n572 71.676
R1388 B.n648 B.n573 71.676
R1389 B.n644 B.n574 71.676
R1390 B.n640 B.n575 71.676
R1391 B.n636 B.n576 71.676
R1392 B.n632 B.n577 71.676
R1393 B.n628 B.n578 71.676
R1394 B.n624 B.n579 71.676
R1395 B.n620 B.n580 71.676
R1396 B.n616 B.n581 71.676
R1397 B.n612 B.n582 71.676
R1398 B.n608 B.n583 71.676
R1399 B.n604 B.n584 71.676
R1400 B.n600 B.n585 71.676
R1401 B.n596 B.n586 71.676
R1402 B.n1171 B.n1170 71.676
R1403 B.n1171 B.n2 71.676
R1404 B.n161 B.n160 64.7763
R1405 B.n159 B.n158 64.7763
R1406 B.n593 B.n592 64.7763
R1407 B.n590 B.n589 64.7763
R1408 B.n284 B.n161 59.5399
R1409 B.n305 B.n159 59.5399
R1410 B.n594 B.n593 59.5399
R1411 B.n591 B.n590 59.5399
R1412 B.n861 B.n517 52.3069
R1413 B.n1071 B.n86 52.3069
R1414 B.n865 B.n864 31.0639
R1415 B.n595 B.n515 31.0639
R1416 B.n1068 B.n1067 31.0639
R1417 B.n1075 B.n1074 31.0639
R1418 B.n868 B.n517 30.4008
R1419 B.n868 B.n513 30.4008
R1420 B.n874 B.n513 30.4008
R1421 B.n874 B.n509 30.4008
R1422 B.n880 B.n509 30.4008
R1423 B.n880 B.n505 30.4008
R1424 B.n887 B.n505 30.4008
R1425 B.n887 B.n886 30.4008
R1426 B.n893 B.n498 30.4008
R1427 B.n899 B.n498 30.4008
R1428 B.n899 B.n494 30.4008
R1429 B.n905 B.n494 30.4008
R1430 B.n905 B.n490 30.4008
R1431 B.n911 B.n490 30.4008
R1432 B.n911 B.n486 30.4008
R1433 B.n917 B.n486 30.4008
R1434 B.n917 B.n482 30.4008
R1435 B.n923 B.n482 30.4008
R1436 B.n923 B.n478 30.4008
R1437 B.n929 B.n478 30.4008
R1438 B.n935 B.n474 30.4008
R1439 B.n935 B.n470 30.4008
R1440 B.n941 B.n470 30.4008
R1441 B.n941 B.n466 30.4008
R1442 B.n947 B.n466 30.4008
R1443 B.n947 B.n462 30.4008
R1444 B.n953 B.n462 30.4008
R1445 B.n953 B.n458 30.4008
R1446 B.n959 B.n458 30.4008
R1447 B.n965 B.n454 30.4008
R1448 B.n965 B.n450 30.4008
R1449 B.n971 B.n450 30.4008
R1450 B.n971 B.n446 30.4008
R1451 B.n977 B.n446 30.4008
R1452 B.n977 B.n442 30.4008
R1453 B.n984 B.n442 30.4008
R1454 B.n984 B.n983 30.4008
R1455 B.n990 B.n435 30.4008
R1456 B.n997 B.n435 30.4008
R1457 B.n997 B.n431 30.4008
R1458 B.n1003 B.n431 30.4008
R1459 B.n1003 B.n4 30.4008
R1460 B.n1169 B.n4 30.4008
R1461 B.n1169 B.n1168 30.4008
R1462 B.n1168 B.n1167 30.4008
R1463 B.n1167 B.n8 30.4008
R1464 B.n12 B.n8 30.4008
R1465 B.n1160 B.n12 30.4008
R1466 B.n1160 B.n1159 30.4008
R1467 B.n1159 B.n1158 30.4008
R1468 B.n1152 B.n19 30.4008
R1469 B.n1152 B.n1151 30.4008
R1470 B.n1151 B.n1150 30.4008
R1471 B.n1150 B.n23 30.4008
R1472 B.n1144 B.n23 30.4008
R1473 B.n1144 B.n1143 30.4008
R1474 B.n1143 B.n1142 30.4008
R1475 B.n1142 B.n30 30.4008
R1476 B.n1136 B.n1135 30.4008
R1477 B.n1135 B.n1134 30.4008
R1478 B.n1134 B.n37 30.4008
R1479 B.n1128 B.n37 30.4008
R1480 B.n1128 B.n1127 30.4008
R1481 B.n1127 B.n1126 30.4008
R1482 B.n1126 B.n44 30.4008
R1483 B.n1120 B.n44 30.4008
R1484 B.n1120 B.n1119 30.4008
R1485 B.n1118 B.n51 30.4008
R1486 B.n1112 B.n51 30.4008
R1487 B.n1112 B.n1111 30.4008
R1488 B.n1111 B.n1110 30.4008
R1489 B.n1110 B.n58 30.4008
R1490 B.n1104 B.n58 30.4008
R1491 B.n1104 B.n1103 30.4008
R1492 B.n1103 B.n1102 30.4008
R1493 B.n1102 B.n65 30.4008
R1494 B.n1096 B.n65 30.4008
R1495 B.n1096 B.n1095 30.4008
R1496 B.n1095 B.n1094 30.4008
R1497 B.n1088 B.n75 30.4008
R1498 B.n1088 B.n1087 30.4008
R1499 B.n1087 B.n1086 30.4008
R1500 B.n1086 B.n79 30.4008
R1501 B.n1080 B.n79 30.4008
R1502 B.n1080 B.n1079 30.4008
R1503 B.n1079 B.n1078 30.4008
R1504 B.n1078 B.n86 30.4008
R1505 B.n983 B.t1 29.9538
R1506 B.n19 B.t19 29.9538
R1507 B.t4 B.n454 25.4831
R1508 B.t2 B.n30 25.4831
R1509 B.n893 B.t10 21.0125
R1510 B.n1094 B.t6 21.0125
R1511 B.t3 B.n474 20.1184
R1512 B.n1119 B.t0 20.1184
R1513 B B.n1172 18.0485
R1514 B.n866 B.n865 10.6151
R1515 B.n866 B.n511 10.6151
R1516 B.n876 B.n511 10.6151
R1517 B.n877 B.n876 10.6151
R1518 B.n878 B.n877 10.6151
R1519 B.n878 B.n503 10.6151
R1520 B.n889 B.n503 10.6151
R1521 B.n890 B.n889 10.6151
R1522 B.n891 B.n890 10.6151
R1523 B.n891 B.n496 10.6151
R1524 B.n901 B.n496 10.6151
R1525 B.n902 B.n901 10.6151
R1526 B.n903 B.n902 10.6151
R1527 B.n903 B.n488 10.6151
R1528 B.n913 B.n488 10.6151
R1529 B.n914 B.n913 10.6151
R1530 B.n915 B.n914 10.6151
R1531 B.n915 B.n480 10.6151
R1532 B.n925 B.n480 10.6151
R1533 B.n926 B.n925 10.6151
R1534 B.n927 B.n926 10.6151
R1535 B.n927 B.n472 10.6151
R1536 B.n937 B.n472 10.6151
R1537 B.n938 B.n937 10.6151
R1538 B.n939 B.n938 10.6151
R1539 B.n939 B.n464 10.6151
R1540 B.n949 B.n464 10.6151
R1541 B.n950 B.n949 10.6151
R1542 B.n951 B.n950 10.6151
R1543 B.n951 B.n456 10.6151
R1544 B.n961 B.n456 10.6151
R1545 B.n962 B.n961 10.6151
R1546 B.n963 B.n962 10.6151
R1547 B.n963 B.n448 10.6151
R1548 B.n973 B.n448 10.6151
R1549 B.n974 B.n973 10.6151
R1550 B.n975 B.n974 10.6151
R1551 B.n975 B.n440 10.6151
R1552 B.n986 B.n440 10.6151
R1553 B.n987 B.n986 10.6151
R1554 B.n988 B.n987 10.6151
R1555 B.n988 B.n433 10.6151
R1556 B.n999 B.n433 10.6151
R1557 B.n1000 B.n999 10.6151
R1558 B.n1001 B.n1000 10.6151
R1559 B.n1001 B.n0 10.6151
R1560 B.n864 B.n519 10.6151
R1561 B.n859 B.n519 10.6151
R1562 B.n859 B.n858 10.6151
R1563 B.n858 B.n857 10.6151
R1564 B.n857 B.n854 10.6151
R1565 B.n854 B.n853 10.6151
R1566 B.n853 B.n850 10.6151
R1567 B.n850 B.n849 10.6151
R1568 B.n849 B.n846 10.6151
R1569 B.n846 B.n845 10.6151
R1570 B.n845 B.n842 10.6151
R1571 B.n842 B.n841 10.6151
R1572 B.n841 B.n838 10.6151
R1573 B.n838 B.n837 10.6151
R1574 B.n837 B.n834 10.6151
R1575 B.n834 B.n833 10.6151
R1576 B.n833 B.n830 10.6151
R1577 B.n830 B.n829 10.6151
R1578 B.n829 B.n826 10.6151
R1579 B.n826 B.n825 10.6151
R1580 B.n825 B.n822 10.6151
R1581 B.n822 B.n821 10.6151
R1582 B.n821 B.n818 10.6151
R1583 B.n818 B.n817 10.6151
R1584 B.n817 B.n814 10.6151
R1585 B.n814 B.n813 10.6151
R1586 B.n813 B.n810 10.6151
R1587 B.n810 B.n809 10.6151
R1588 B.n809 B.n806 10.6151
R1589 B.n806 B.n805 10.6151
R1590 B.n805 B.n802 10.6151
R1591 B.n802 B.n801 10.6151
R1592 B.n801 B.n798 10.6151
R1593 B.n798 B.n797 10.6151
R1594 B.n797 B.n794 10.6151
R1595 B.n794 B.n793 10.6151
R1596 B.n793 B.n790 10.6151
R1597 B.n790 B.n789 10.6151
R1598 B.n789 B.n786 10.6151
R1599 B.n786 B.n785 10.6151
R1600 B.n785 B.n782 10.6151
R1601 B.n782 B.n781 10.6151
R1602 B.n781 B.n778 10.6151
R1603 B.n778 B.n777 10.6151
R1604 B.n777 B.n774 10.6151
R1605 B.n774 B.n773 10.6151
R1606 B.n773 B.n770 10.6151
R1607 B.n770 B.n769 10.6151
R1608 B.n769 B.n766 10.6151
R1609 B.n766 B.n765 10.6151
R1610 B.n765 B.n762 10.6151
R1611 B.n762 B.n761 10.6151
R1612 B.n761 B.n758 10.6151
R1613 B.n758 B.n757 10.6151
R1614 B.n757 B.n754 10.6151
R1615 B.n754 B.n753 10.6151
R1616 B.n753 B.n750 10.6151
R1617 B.n750 B.n749 10.6151
R1618 B.n749 B.n746 10.6151
R1619 B.n746 B.n745 10.6151
R1620 B.n745 B.n742 10.6151
R1621 B.n742 B.n741 10.6151
R1622 B.n738 B.n737 10.6151
R1623 B.n737 B.n734 10.6151
R1624 B.n734 B.n733 10.6151
R1625 B.n733 B.n730 10.6151
R1626 B.n730 B.n729 10.6151
R1627 B.n729 B.n726 10.6151
R1628 B.n726 B.n725 10.6151
R1629 B.n725 B.n722 10.6151
R1630 B.n722 B.n721 10.6151
R1631 B.n718 B.n717 10.6151
R1632 B.n717 B.n714 10.6151
R1633 B.n714 B.n713 10.6151
R1634 B.n713 B.n710 10.6151
R1635 B.n710 B.n709 10.6151
R1636 B.n709 B.n706 10.6151
R1637 B.n706 B.n705 10.6151
R1638 B.n705 B.n702 10.6151
R1639 B.n702 B.n701 10.6151
R1640 B.n701 B.n698 10.6151
R1641 B.n698 B.n697 10.6151
R1642 B.n697 B.n694 10.6151
R1643 B.n694 B.n693 10.6151
R1644 B.n693 B.n690 10.6151
R1645 B.n690 B.n689 10.6151
R1646 B.n689 B.n686 10.6151
R1647 B.n686 B.n685 10.6151
R1648 B.n685 B.n682 10.6151
R1649 B.n682 B.n681 10.6151
R1650 B.n681 B.n678 10.6151
R1651 B.n678 B.n677 10.6151
R1652 B.n677 B.n674 10.6151
R1653 B.n674 B.n673 10.6151
R1654 B.n673 B.n670 10.6151
R1655 B.n670 B.n669 10.6151
R1656 B.n669 B.n666 10.6151
R1657 B.n666 B.n665 10.6151
R1658 B.n665 B.n662 10.6151
R1659 B.n662 B.n661 10.6151
R1660 B.n661 B.n658 10.6151
R1661 B.n658 B.n657 10.6151
R1662 B.n657 B.n654 10.6151
R1663 B.n654 B.n653 10.6151
R1664 B.n653 B.n650 10.6151
R1665 B.n650 B.n649 10.6151
R1666 B.n649 B.n646 10.6151
R1667 B.n646 B.n645 10.6151
R1668 B.n645 B.n642 10.6151
R1669 B.n642 B.n641 10.6151
R1670 B.n641 B.n638 10.6151
R1671 B.n638 B.n637 10.6151
R1672 B.n637 B.n634 10.6151
R1673 B.n634 B.n633 10.6151
R1674 B.n633 B.n630 10.6151
R1675 B.n630 B.n629 10.6151
R1676 B.n629 B.n626 10.6151
R1677 B.n626 B.n625 10.6151
R1678 B.n625 B.n622 10.6151
R1679 B.n622 B.n621 10.6151
R1680 B.n621 B.n618 10.6151
R1681 B.n618 B.n617 10.6151
R1682 B.n617 B.n614 10.6151
R1683 B.n614 B.n613 10.6151
R1684 B.n613 B.n610 10.6151
R1685 B.n610 B.n609 10.6151
R1686 B.n609 B.n606 10.6151
R1687 B.n606 B.n605 10.6151
R1688 B.n605 B.n602 10.6151
R1689 B.n602 B.n601 10.6151
R1690 B.n601 B.n598 10.6151
R1691 B.n598 B.n597 10.6151
R1692 B.n597 B.n595 10.6151
R1693 B.n870 B.n515 10.6151
R1694 B.n871 B.n870 10.6151
R1695 B.n872 B.n871 10.6151
R1696 B.n872 B.n507 10.6151
R1697 B.n882 B.n507 10.6151
R1698 B.n883 B.n882 10.6151
R1699 B.n884 B.n883 10.6151
R1700 B.n884 B.n500 10.6151
R1701 B.n895 B.n500 10.6151
R1702 B.n896 B.n895 10.6151
R1703 B.n897 B.n896 10.6151
R1704 B.n897 B.n492 10.6151
R1705 B.n907 B.n492 10.6151
R1706 B.n908 B.n907 10.6151
R1707 B.n909 B.n908 10.6151
R1708 B.n909 B.n484 10.6151
R1709 B.n919 B.n484 10.6151
R1710 B.n920 B.n919 10.6151
R1711 B.n921 B.n920 10.6151
R1712 B.n921 B.n476 10.6151
R1713 B.n931 B.n476 10.6151
R1714 B.n932 B.n931 10.6151
R1715 B.n933 B.n932 10.6151
R1716 B.n933 B.n468 10.6151
R1717 B.n943 B.n468 10.6151
R1718 B.n944 B.n943 10.6151
R1719 B.n945 B.n944 10.6151
R1720 B.n945 B.n460 10.6151
R1721 B.n955 B.n460 10.6151
R1722 B.n956 B.n955 10.6151
R1723 B.n957 B.n956 10.6151
R1724 B.n957 B.n452 10.6151
R1725 B.n967 B.n452 10.6151
R1726 B.n968 B.n967 10.6151
R1727 B.n969 B.n968 10.6151
R1728 B.n969 B.n444 10.6151
R1729 B.n979 B.n444 10.6151
R1730 B.n980 B.n979 10.6151
R1731 B.n981 B.n980 10.6151
R1732 B.n981 B.n437 10.6151
R1733 B.n992 B.n437 10.6151
R1734 B.n993 B.n992 10.6151
R1735 B.n995 B.n993 10.6151
R1736 B.n995 B.n994 10.6151
R1737 B.n994 B.n429 10.6151
R1738 B.n1006 B.n429 10.6151
R1739 B.n1007 B.n1006 10.6151
R1740 B.n1008 B.n1007 10.6151
R1741 B.n1009 B.n1008 10.6151
R1742 B.n1010 B.n1009 10.6151
R1743 B.n1013 B.n1010 10.6151
R1744 B.n1014 B.n1013 10.6151
R1745 B.n1015 B.n1014 10.6151
R1746 B.n1016 B.n1015 10.6151
R1747 B.n1018 B.n1016 10.6151
R1748 B.n1019 B.n1018 10.6151
R1749 B.n1020 B.n1019 10.6151
R1750 B.n1021 B.n1020 10.6151
R1751 B.n1023 B.n1021 10.6151
R1752 B.n1024 B.n1023 10.6151
R1753 B.n1025 B.n1024 10.6151
R1754 B.n1026 B.n1025 10.6151
R1755 B.n1028 B.n1026 10.6151
R1756 B.n1029 B.n1028 10.6151
R1757 B.n1030 B.n1029 10.6151
R1758 B.n1031 B.n1030 10.6151
R1759 B.n1033 B.n1031 10.6151
R1760 B.n1034 B.n1033 10.6151
R1761 B.n1035 B.n1034 10.6151
R1762 B.n1036 B.n1035 10.6151
R1763 B.n1038 B.n1036 10.6151
R1764 B.n1039 B.n1038 10.6151
R1765 B.n1040 B.n1039 10.6151
R1766 B.n1041 B.n1040 10.6151
R1767 B.n1043 B.n1041 10.6151
R1768 B.n1044 B.n1043 10.6151
R1769 B.n1045 B.n1044 10.6151
R1770 B.n1046 B.n1045 10.6151
R1771 B.n1048 B.n1046 10.6151
R1772 B.n1049 B.n1048 10.6151
R1773 B.n1050 B.n1049 10.6151
R1774 B.n1051 B.n1050 10.6151
R1775 B.n1053 B.n1051 10.6151
R1776 B.n1054 B.n1053 10.6151
R1777 B.n1055 B.n1054 10.6151
R1778 B.n1056 B.n1055 10.6151
R1779 B.n1058 B.n1056 10.6151
R1780 B.n1059 B.n1058 10.6151
R1781 B.n1060 B.n1059 10.6151
R1782 B.n1061 B.n1060 10.6151
R1783 B.n1063 B.n1061 10.6151
R1784 B.n1064 B.n1063 10.6151
R1785 B.n1065 B.n1064 10.6151
R1786 B.n1066 B.n1065 10.6151
R1787 B.n1067 B.n1066 10.6151
R1788 B.n1164 B.n1 10.6151
R1789 B.n1164 B.n1163 10.6151
R1790 B.n1163 B.n1162 10.6151
R1791 B.n1162 B.n10 10.6151
R1792 B.n1156 B.n10 10.6151
R1793 B.n1156 B.n1155 10.6151
R1794 B.n1155 B.n1154 10.6151
R1795 B.n1154 B.n17 10.6151
R1796 B.n1148 B.n17 10.6151
R1797 B.n1148 B.n1147 10.6151
R1798 B.n1147 B.n1146 10.6151
R1799 B.n1146 B.n25 10.6151
R1800 B.n1140 B.n25 10.6151
R1801 B.n1140 B.n1139 10.6151
R1802 B.n1139 B.n1138 10.6151
R1803 B.n1138 B.n32 10.6151
R1804 B.n1132 B.n32 10.6151
R1805 B.n1132 B.n1131 10.6151
R1806 B.n1131 B.n1130 10.6151
R1807 B.n1130 B.n39 10.6151
R1808 B.n1124 B.n39 10.6151
R1809 B.n1124 B.n1123 10.6151
R1810 B.n1123 B.n1122 10.6151
R1811 B.n1122 B.n46 10.6151
R1812 B.n1116 B.n46 10.6151
R1813 B.n1116 B.n1115 10.6151
R1814 B.n1115 B.n1114 10.6151
R1815 B.n1114 B.n53 10.6151
R1816 B.n1108 B.n53 10.6151
R1817 B.n1108 B.n1107 10.6151
R1818 B.n1107 B.n1106 10.6151
R1819 B.n1106 B.n60 10.6151
R1820 B.n1100 B.n60 10.6151
R1821 B.n1100 B.n1099 10.6151
R1822 B.n1099 B.n1098 10.6151
R1823 B.n1098 B.n67 10.6151
R1824 B.n1092 B.n67 10.6151
R1825 B.n1092 B.n1091 10.6151
R1826 B.n1091 B.n1090 10.6151
R1827 B.n1090 B.n73 10.6151
R1828 B.n1084 B.n73 10.6151
R1829 B.n1084 B.n1083 10.6151
R1830 B.n1083 B.n1082 10.6151
R1831 B.n1082 B.n81 10.6151
R1832 B.n1076 B.n81 10.6151
R1833 B.n1076 B.n1075 10.6151
R1834 B.n1074 B.n88 10.6151
R1835 B.n163 B.n88 10.6151
R1836 B.n164 B.n163 10.6151
R1837 B.n167 B.n164 10.6151
R1838 B.n168 B.n167 10.6151
R1839 B.n171 B.n168 10.6151
R1840 B.n172 B.n171 10.6151
R1841 B.n175 B.n172 10.6151
R1842 B.n176 B.n175 10.6151
R1843 B.n179 B.n176 10.6151
R1844 B.n180 B.n179 10.6151
R1845 B.n183 B.n180 10.6151
R1846 B.n184 B.n183 10.6151
R1847 B.n187 B.n184 10.6151
R1848 B.n188 B.n187 10.6151
R1849 B.n191 B.n188 10.6151
R1850 B.n192 B.n191 10.6151
R1851 B.n195 B.n192 10.6151
R1852 B.n196 B.n195 10.6151
R1853 B.n199 B.n196 10.6151
R1854 B.n200 B.n199 10.6151
R1855 B.n203 B.n200 10.6151
R1856 B.n204 B.n203 10.6151
R1857 B.n207 B.n204 10.6151
R1858 B.n208 B.n207 10.6151
R1859 B.n211 B.n208 10.6151
R1860 B.n212 B.n211 10.6151
R1861 B.n215 B.n212 10.6151
R1862 B.n216 B.n215 10.6151
R1863 B.n219 B.n216 10.6151
R1864 B.n220 B.n219 10.6151
R1865 B.n223 B.n220 10.6151
R1866 B.n224 B.n223 10.6151
R1867 B.n227 B.n224 10.6151
R1868 B.n228 B.n227 10.6151
R1869 B.n231 B.n228 10.6151
R1870 B.n232 B.n231 10.6151
R1871 B.n235 B.n232 10.6151
R1872 B.n236 B.n235 10.6151
R1873 B.n239 B.n236 10.6151
R1874 B.n240 B.n239 10.6151
R1875 B.n243 B.n240 10.6151
R1876 B.n244 B.n243 10.6151
R1877 B.n247 B.n244 10.6151
R1878 B.n248 B.n247 10.6151
R1879 B.n251 B.n248 10.6151
R1880 B.n252 B.n251 10.6151
R1881 B.n255 B.n252 10.6151
R1882 B.n256 B.n255 10.6151
R1883 B.n259 B.n256 10.6151
R1884 B.n260 B.n259 10.6151
R1885 B.n263 B.n260 10.6151
R1886 B.n264 B.n263 10.6151
R1887 B.n267 B.n264 10.6151
R1888 B.n268 B.n267 10.6151
R1889 B.n271 B.n268 10.6151
R1890 B.n272 B.n271 10.6151
R1891 B.n275 B.n272 10.6151
R1892 B.n276 B.n275 10.6151
R1893 B.n279 B.n276 10.6151
R1894 B.n280 B.n279 10.6151
R1895 B.n283 B.n280 10.6151
R1896 B.n288 B.n285 10.6151
R1897 B.n289 B.n288 10.6151
R1898 B.n292 B.n289 10.6151
R1899 B.n293 B.n292 10.6151
R1900 B.n296 B.n293 10.6151
R1901 B.n297 B.n296 10.6151
R1902 B.n300 B.n297 10.6151
R1903 B.n301 B.n300 10.6151
R1904 B.n304 B.n301 10.6151
R1905 B.n309 B.n306 10.6151
R1906 B.n310 B.n309 10.6151
R1907 B.n313 B.n310 10.6151
R1908 B.n314 B.n313 10.6151
R1909 B.n317 B.n314 10.6151
R1910 B.n318 B.n317 10.6151
R1911 B.n321 B.n318 10.6151
R1912 B.n322 B.n321 10.6151
R1913 B.n325 B.n322 10.6151
R1914 B.n326 B.n325 10.6151
R1915 B.n329 B.n326 10.6151
R1916 B.n330 B.n329 10.6151
R1917 B.n333 B.n330 10.6151
R1918 B.n334 B.n333 10.6151
R1919 B.n337 B.n334 10.6151
R1920 B.n338 B.n337 10.6151
R1921 B.n341 B.n338 10.6151
R1922 B.n342 B.n341 10.6151
R1923 B.n345 B.n342 10.6151
R1924 B.n346 B.n345 10.6151
R1925 B.n349 B.n346 10.6151
R1926 B.n350 B.n349 10.6151
R1927 B.n353 B.n350 10.6151
R1928 B.n354 B.n353 10.6151
R1929 B.n357 B.n354 10.6151
R1930 B.n358 B.n357 10.6151
R1931 B.n361 B.n358 10.6151
R1932 B.n362 B.n361 10.6151
R1933 B.n365 B.n362 10.6151
R1934 B.n366 B.n365 10.6151
R1935 B.n369 B.n366 10.6151
R1936 B.n370 B.n369 10.6151
R1937 B.n373 B.n370 10.6151
R1938 B.n374 B.n373 10.6151
R1939 B.n377 B.n374 10.6151
R1940 B.n378 B.n377 10.6151
R1941 B.n381 B.n378 10.6151
R1942 B.n382 B.n381 10.6151
R1943 B.n385 B.n382 10.6151
R1944 B.n386 B.n385 10.6151
R1945 B.n389 B.n386 10.6151
R1946 B.n390 B.n389 10.6151
R1947 B.n393 B.n390 10.6151
R1948 B.n394 B.n393 10.6151
R1949 B.n397 B.n394 10.6151
R1950 B.n398 B.n397 10.6151
R1951 B.n401 B.n398 10.6151
R1952 B.n402 B.n401 10.6151
R1953 B.n405 B.n402 10.6151
R1954 B.n406 B.n405 10.6151
R1955 B.n409 B.n406 10.6151
R1956 B.n410 B.n409 10.6151
R1957 B.n413 B.n410 10.6151
R1958 B.n414 B.n413 10.6151
R1959 B.n417 B.n414 10.6151
R1960 B.n418 B.n417 10.6151
R1961 B.n421 B.n418 10.6151
R1962 B.n422 B.n421 10.6151
R1963 B.n425 B.n422 10.6151
R1964 B.n427 B.n425 10.6151
R1965 B.n428 B.n427 10.6151
R1966 B.n1068 B.n428 10.6151
R1967 B.n929 B.t3 10.283
R1968 B.t0 B.n1118 10.283
R1969 B.n886 B.t10 9.38884
R1970 B.n75 B.t6 9.38884
R1971 B.n741 B.n591 9.36635
R1972 B.n718 B.n594 9.36635
R1973 B.n284 B.n283 9.36635
R1974 B.n306 B.n305 9.36635
R1975 B.n1172 B.n0 8.11757
R1976 B.n1172 B.n1 8.11757
R1977 B.n959 B.t4 4.9182
R1978 B.n1136 B.t2 4.9182
R1979 B.n738 B.n591 1.24928
R1980 B.n721 B.n594 1.24928
R1981 B.n285 B.n284 1.24928
R1982 B.n305 B.n304 1.24928
R1983 B.n990 B.t1 0.447564
R1984 B.n1158 B.t19 0.447564
R1985 VP.n11 VP.t1 188.018
R1986 VP.n13 VP.n10 161.3
R1987 VP.n15 VP.n14 161.3
R1988 VP.n16 VP.n9 161.3
R1989 VP.n18 VP.n17 161.3
R1990 VP.n19 VP.n8 161.3
R1991 VP.n21 VP.n20 161.3
R1992 VP.n44 VP.n43 161.3
R1993 VP.n42 VP.n1 161.3
R1994 VP.n41 VP.n40 161.3
R1995 VP.n39 VP.n2 161.3
R1996 VP.n38 VP.n37 161.3
R1997 VP.n36 VP.n3 161.3
R1998 VP.n35 VP.n34 161.3
R1999 VP.n33 VP.n4 161.3
R2000 VP.n32 VP.n31 161.3
R2001 VP.n30 VP.n5 161.3
R2002 VP.n29 VP.n28 161.3
R2003 VP.n27 VP.n6 161.3
R2004 VP.n26 VP.n25 161.3
R2005 VP.n35 VP.t4 154.768
R2006 VP.n24 VP.t0 154.768
R2007 VP.n0 VP.t5 154.768
R2008 VP.n12 VP.t3 154.768
R2009 VP.n7 VP.t2 154.768
R2010 VP.n24 VP.n23 73.4298
R2011 VP.n45 VP.n0 73.4298
R2012 VP.n22 VP.n7 73.4298
R2013 VP.n30 VP.n29 56.5193
R2014 VP.n41 VP.n2 56.5193
R2015 VP.n18 VP.n9 56.5193
R2016 VP.n23 VP.n22 55.9084
R2017 VP.n12 VP.n11 49.2372
R2018 VP.n25 VP.n6 24.4675
R2019 VP.n29 VP.n6 24.4675
R2020 VP.n31 VP.n30 24.4675
R2021 VP.n31 VP.n4 24.4675
R2022 VP.n35 VP.n4 24.4675
R2023 VP.n36 VP.n35 24.4675
R2024 VP.n37 VP.n36 24.4675
R2025 VP.n37 VP.n2 24.4675
R2026 VP.n42 VP.n41 24.4675
R2027 VP.n43 VP.n42 24.4675
R2028 VP.n19 VP.n18 24.4675
R2029 VP.n20 VP.n19 24.4675
R2030 VP.n13 VP.n12 24.4675
R2031 VP.n14 VP.n13 24.4675
R2032 VP.n14 VP.n9 24.4675
R2033 VP.n25 VP.n24 16.6381
R2034 VP.n43 VP.n0 16.6381
R2035 VP.n20 VP.n7 16.6381
R2036 VP.n11 VP.n10 4.07657
R2037 VP.n22 VP.n21 0.354971
R2038 VP.n26 VP.n23 0.354971
R2039 VP.n45 VP.n44 0.354971
R2040 VP VP.n45 0.26696
R2041 VP.n15 VP.n10 0.189894
R2042 VP.n16 VP.n15 0.189894
R2043 VP.n17 VP.n16 0.189894
R2044 VP.n17 VP.n8 0.189894
R2045 VP.n21 VP.n8 0.189894
R2046 VP.n27 VP.n26 0.189894
R2047 VP.n28 VP.n27 0.189894
R2048 VP.n28 VP.n5 0.189894
R2049 VP.n32 VP.n5 0.189894
R2050 VP.n33 VP.n32 0.189894
R2051 VP.n34 VP.n33 0.189894
R2052 VP.n34 VP.n3 0.189894
R2053 VP.n38 VP.n3 0.189894
R2054 VP.n39 VP.n38 0.189894
R2055 VP.n40 VP.n39 0.189894
R2056 VP.n40 VP.n1 0.189894
R2057 VP.n44 VP.n1 0.189894
R2058 VTAIL.n7 VTAIL.t1 45.1506
R2059 VTAIL.n11 VTAIL.t0 45.1504
R2060 VTAIL.n2 VTAIL.t10 45.1504
R2061 VTAIL.n10 VTAIL.t5 45.1504
R2062 VTAIL.n9 VTAIL.n8 44.1263
R2063 VTAIL.n6 VTAIL.n5 44.1263
R2064 VTAIL.n1 VTAIL.n0 44.1262
R2065 VTAIL.n4 VTAIL.n3 44.1262
R2066 VTAIL.n6 VTAIL.n4 34.7893
R2067 VTAIL.n11 VTAIL.n10 31.91
R2068 VTAIL.n7 VTAIL.n6 2.87981
R2069 VTAIL.n10 VTAIL.n9 2.87981
R2070 VTAIL.n4 VTAIL.n2 2.87981
R2071 VTAIL VTAIL.n11 2.10179
R2072 VTAIL.n9 VTAIL.n7 1.90998
R2073 VTAIL.n2 VTAIL.n1 1.90998
R2074 VTAIL.n0 VTAIL.t11 1.02481
R2075 VTAIL.n0 VTAIL.t4 1.02481
R2076 VTAIL.n3 VTAIL.t8 1.02481
R2077 VTAIL.n3 VTAIL.t6 1.02481
R2078 VTAIL.n8 VTAIL.t9 1.02481
R2079 VTAIL.n8 VTAIL.t7 1.02481
R2080 VTAIL.n5 VTAIL.t2 1.02481
R2081 VTAIL.n5 VTAIL.t3 1.02481
R2082 VTAIL VTAIL.n1 0.778517
R2083 VDD1 VDD1.t4 64.0471
R2084 VDD1.n1 VDD1.t5 63.9333
R2085 VDD1.n1 VDD1.n0 61.4695
R2086 VDD1.n3 VDD1.n2 60.8049
R2087 VDD1.n3 VDD1.n1 51.7595
R2088 VDD1.n2 VDD1.t2 1.02481
R2089 VDD1.n2 VDD1.t3 1.02481
R2090 VDD1.n0 VDD1.t1 1.02481
R2091 VDD1.n0 VDD1.t0 1.02481
R2092 VDD1 VDD1.n3 0.662138
R2093 VN.n20 VN.t3 188.018
R2094 VN.n4 VN.t0 188.018
R2095 VN.n30 VN.n29 161.3
R2096 VN.n28 VN.n17 161.3
R2097 VN.n27 VN.n26 161.3
R2098 VN.n25 VN.n18 161.3
R2099 VN.n24 VN.n23 161.3
R2100 VN.n22 VN.n19 161.3
R2101 VN.n14 VN.n13 161.3
R2102 VN.n12 VN.n1 161.3
R2103 VN.n11 VN.n10 161.3
R2104 VN.n9 VN.n2 161.3
R2105 VN.n8 VN.n7 161.3
R2106 VN.n6 VN.n3 161.3
R2107 VN.n5 VN.t4 154.768
R2108 VN.n0 VN.t2 154.768
R2109 VN.n21 VN.t5 154.768
R2110 VN.n16 VN.t1 154.768
R2111 VN.n15 VN.n0 73.4298
R2112 VN.n31 VN.n16 73.4298
R2113 VN.n11 VN.n2 56.5193
R2114 VN.n27 VN.n18 56.5193
R2115 VN VN.n31 56.0738
R2116 VN.n5 VN.n4 49.2372
R2117 VN.n21 VN.n20 49.2372
R2118 VN.n6 VN.n5 24.4675
R2119 VN.n7 VN.n6 24.4675
R2120 VN.n7 VN.n2 24.4675
R2121 VN.n12 VN.n11 24.4675
R2122 VN.n13 VN.n12 24.4675
R2123 VN.n23 VN.n18 24.4675
R2124 VN.n23 VN.n22 24.4675
R2125 VN.n22 VN.n21 24.4675
R2126 VN.n29 VN.n28 24.4675
R2127 VN.n28 VN.n27 24.4675
R2128 VN.n13 VN.n0 16.6381
R2129 VN.n29 VN.n16 16.6381
R2130 VN.n20 VN.n19 4.07659
R2131 VN.n4 VN.n3 4.07659
R2132 VN.n31 VN.n30 0.354971
R2133 VN.n15 VN.n14 0.354971
R2134 VN VN.n15 0.26696
R2135 VN.n30 VN.n17 0.189894
R2136 VN.n26 VN.n17 0.189894
R2137 VN.n26 VN.n25 0.189894
R2138 VN.n25 VN.n24 0.189894
R2139 VN.n24 VN.n19 0.189894
R2140 VN.n8 VN.n3 0.189894
R2141 VN.n9 VN.n8 0.189894
R2142 VN.n10 VN.n9 0.189894
R2143 VN.n10 VN.n1 0.189894
R2144 VN.n14 VN.n1 0.189894
R2145 VDD2.n1 VDD2.t5 63.9333
R2146 VDD2.n2 VDD2.t4 61.8294
R2147 VDD2.n1 VDD2.n0 61.4695
R2148 VDD2 VDD2.n3 61.4665
R2149 VDD2.n2 VDD2.n1 49.7368
R2150 VDD2 VDD2.n2 2.21817
R2151 VDD2.n3 VDD2.t0 1.02481
R2152 VDD2.n3 VDD2.t2 1.02481
R2153 VDD2.n0 VDD2.t1 1.02481
R2154 VDD2.n0 VDD2.t3 1.02481
C0 VDD1 VN 0.151387f
C1 VN VTAIL 10.8028f
C2 VN VP 8.686861f
C3 VDD1 VDD2 1.56821f
C4 VTAIL VDD2 10.4033f
C5 VP VDD2 0.493688f
C6 VN VDD2 10.8779f
C7 VDD1 VTAIL 10.350801f
C8 VDD1 VP 11.216001f
C9 VP VTAIL 10.817201f
C10 VDD2 B 7.604861f
C11 VDD1 B 7.949708f
C12 VTAIL B 11.058321f
C13 VN B 14.70707f
C14 VP B 13.262875f
C15 VDD2.t5 B 3.78251f
C16 VDD2.t1 B 0.322708f
C17 VDD2.t3 B 0.322708f
C18 VDD2.n0 B 2.95237f
C19 VDD2.n1 B 3.00148f
C20 VDD2.t4 B 3.76979f
C21 VDD2.n2 B 2.93309f
C22 VDD2.t0 B 0.322708f
C23 VDD2.t2 B 0.322708f
C24 VDD2.n3 B 2.95232f
C25 VN.t2 B 3.20174f
C26 VN.n0 B 1.1791f
C27 VN.n1 B 0.01998f
C28 VN.n2 B 0.024713f
C29 VN.n3 B 0.227119f
C30 VN.t4 B 3.20174f
C31 VN.t0 B 3.42124f
C32 VN.n4 B 1.1323f
C33 VN.n5 B 1.17839f
C34 VN.n6 B 0.037238f
C35 VN.n7 B 0.037238f
C36 VN.n8 B 0.01998f
C37 VN.n9 B 0.01998f
C38 VN.n10 B 0.01998f
C39 VN.n11 B 0.033622f
C40 VN.n12 B 0.037238f
C41 VN.n13 B 0.031355f
C42 VN.n14 B 0.032248f
C43 VN.n15 B 0.044494f
C44 VN.t1 B 3.20174f
C45 VN.n16 B 1.1791f
C46 VN.n17 B 0.01998f
C47 VN.n18 B 0.024713f
C48 VN.n19 B 0.227119f
C49 VN.t5 B 3.20174f
C50 VN.t3 B 3.42124f
C51 VN.n20 B 1.1323f
C52 VN.n21 B 1.17839f
C53 VN.n22 B 0.037238f
C54 VN.n23 B 0.037238f
C55 VN.n24 B 0.01998f
C56 VN.n25 B 0.01998f
C57 VN.n26 B 0.01998f
C58 VN.n27 B 0.033622f
C59 VN.n28 B 0.037238f
C60 VN.n29 B 0.031355f
C61 VN.n30 B 0.032248f
C62 VN.n31 B 1.3322f
C63 VDD1.t4 B 3.82272f
C64 VDD1.t5 B 3.82179f
C65 VDD1.t1 B 0.326059f
C66 VDD1.t0 B 0.326059f
C67 VDD1.n0 B 2.98302f
C68 VDD1.n1 B 3.15222f
C69 VDD1.t2 B 0.326059f
C70 VDD1.t3 B 0.326059f
C71 VDD1.n2 B 2.97834f
C72 VDD1.n3 B 2.95516f
C73 VTAIL.t11 B 0.343645f
C74 VTAIL.t4 B 0.343645f
C75 VTAIL.n0 B 3.06952f
C76 VTAIL.n1 B 0.421797f
C77 VTAIL.t10 B 3.92362f
C78 VTAIL.n2 B 0.657235f
C79 VTAIL.t8 B 0.343645f
C80 VTAIL.t6 B 0.343645f
C81 VTAIL.n3 B 3.06952f
C82 VTAIL.n4 B 2.3667f
C83 VTAIL.t2 B 0.343645f
C84 VTAIL.t3 B 0.343645f
C85 VTAIL.n5 B 3.06951f
C86 VTAIL.n6 B 2.36671f
C87 VTAIL.t1 B 3.92362f
C88 VTAIL.n7 B 0.657231f
C89 VTAIL.t9 B 0.343645f
C90 VTAIL.t7 B 0.343645f
C91 VTAIL.n8 B 3.06951f
C92 VTAIL.n9 B 0.574127f
C93 VTAIL.t5 B 3.92361f
C94 VTAIL.n10 B 2.2411f
C95 VTAIL.t0 B 3.92362f
C96 VTAIL.n11 B 2.1847f
C97 VP.t5 B 3.23633f
C98 VP.n0 B 1.19184f
C99 VP.n1 B 0.020196f
C100 VP.n2 B 0.02498f
C101 VP.n3 B 0.020196f
C102 VP.t4 B 3.23633f
C103 VP.n4 B 0.037641f
C104 VP.n5 B 0.020196f
C105 VP.n6 B 0.037641f
C106 VP.t2 B 3.23633f
C107 VP.n7 B 1.19184f
C108 VP.n8 B 0.020196f
C109 VP.n9 B 0.02498f
C110 VP.n10 B 0.229572f
C111 VP.t3 B 3.23633f
C112 VP.t1 B 3.4582f
C113 VP.n11 B 1.14453f
C114 VP.n12 B 1.19112f
C115 VP.n13 B 0.037641f
C116 VP.n14 B 0.037641f
C117 VP.n15 B 0.020196f
C118 VP.n16 B 0.020196f
C119 VP.n17 B 0.020196f
C120 VP.n18 B 0.033985f
C121 VP.n19 B 0.037641f
C122 VP.n20 B 0.031694f
C123 VP.n21 B 0.032596f
C124 VP.n22 B 1.33862f
C125 VP.n23 B 1.35161f
C126 VP.t0 B 3.23633f
C127 VP.n24 B 1.19184f
C128 VP.n25 B 0.031694f
C129 VP.n26 B 0.032596f
C130 VP.n27 B 0.020196f
C131 VP.n28 B 0.020196f
C132 VP.n29 B 0.033985f
C133 VP.n30 B 0.02498f
C134 VP.n31 B 0.037641f
C135 VP.n32 B 0.020196f
C136 VP.n33 B 0.020196f
C137 VP.n34 B 0.020196f
C138 VP.n35 B 1.13535f
C139 VP.n36 B 0.037641f
C140 VP.n37 B 0.037641f
C141 VP.n38 B 0.020196f
C142 VP.n39 B 0.020196f
C143 VP.n40 B 0.020196f
C144 VP.n41 B 0.033985f
C145 VP.n42 B 0.037641f
C146 VP.n43 B 0.031694f
C147 VP.n44 B 0.032596f
C148 VP.n45 B 0.044974f
.ends

