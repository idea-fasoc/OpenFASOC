* NGSPICE file created from diff_pair_sample_1796.ext - technology: sky130A

.subckt diff_pair_sample_1796 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X1 VTAIL.t12 VN.t1 VDD2.t6 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=2.08065 ps=12.94 w=12.61 l=1.88
X2 VDD1.t7 VP.t0 VTAIL.t6 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X3 VDD2.t5 VN.t2 VTAIL.t8 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X4 B.t11 B.t9 B.t10 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=0 ps=0 w=12.61 l=1.88
X5 VTAIL.t15 VN.t3 VDD2.t4 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=2.08065 ps=12.94 w=12.61 l=1.88
X6 VDD1.t6 VP.t1 VTAIL.t1 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=4.9179 ps=26 w=12.61 l=1.88
X7 VTAIL.t14 VN.t4 VDD2.t3 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X8 VTAIL.t5 VP.t2 VDD1.t5 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X9 VDD2.t2 VN.t5 VTAIL.t13 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=4.9179 ps=26 w=12.61 l=1.88
X10 VTAIL.t7 VP.t3 VDD1.t4 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X11 VDD2.t1 VN.t6 VTAIL.t9 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=4.9179 ps=26 w=12.61 l=1.88
X12 VDD1.t3 VP.t4 VTAIL.t4 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X13 VDD1.t2 VP.t5 VTAIL.t3 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=4.9179 ps=26 w=12.61 l=1.88
X14 B.t8 B.t6 B.t7 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=0 ps=0 w=12.61 l=1.88
X15 VTAIL.t0 VP.t6 VDD1.t1 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=2.08065 ps=12.94 w=12.61 l=1.88
X16 VTAIL.t10 VN.t7 VDD2.t0 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=2.08065 pd=12.94 as=2.08065 ps=12.94 w=12.61 l=1.88
X17 B.t5 B.t3 B.t4 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=0 ps=0 w=12.61 l=1.88
X18 B.t2 B.t0 B.t1 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=0 ps=0 w=12.61 l=1.88
X19 VTAIL.t2 VP.t7 VDD1.t0 w_n3180_n3490# sky130_fd_pr__pfet_01v8 ad=4.9179 pd=26 as=2.08065 ps=12.94 w=12.61 l=1.88
R0 VN.n5 VN.t1 195.512
R1 VN.n28 VN.t6 195.512
R2 VN.n22 VN.n21 182.587
R3 VN.n45 VN.n44 182.587
R4 VN.n6 VN.t2 161.649
R5 VN.n13 VN.t4 161.649
R6 VN.n21 VN.t5 161.649
R7 VN.n29 VN.t7 161.649
R8 VN.n36 VN.t0 161.649
R9 VN.n44 VN.t3 161.649
R10 VN.n43 VN.n23 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n24 161.3
R13 VN.n39 VN.n38 161.3
R14 VN.n37 VN.n25 161.3
R15 VN.n35 VN.n34 161.3
R16 VN.n33 VN.n26 161.3
R17 VN.n32 VN.n31 161.3
R18 VN.n30 VN.n27 161.3
R19 VN.n20 VN.n0 161.3
R20 VN.n19 VN.n18 161.3
R21 VN.n17 VN.n1 161.3
R22 VN.n16 VN.n15 161.3
R23 VN.n14 VN.n2 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n3 161.3
R26 VN.n9 VN.n8 161.3
R27 VN.n7 VN.n4 161.3
R28 VN.n8 VN.n3 56.5193
R29 VN.n31 VN.n26 56.5193
R30 VN.n6 VN.n5 52.3231
R31 VN.n29 VN.n28 52.3231
R32 VN VN.n45 48.2827
R33 VN.n15 VN.n1 44.3785
R34 VN.n38 VN.n24 44.3785
R35 VN.n19 VN.n1 36.6083
R36 VN.n42 VN.n24 36.6083
R37 VN.n8 VN.n7 24.4675
R38 VN.n12 VN.n3 24.4675
R39 VN.n15 VN.n14 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n37 24.4675
R43 VN.n35 VN.n26 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n7 VN.n6 17.3721
R46 VN.n13 VN.n12 17.3721
R47 VN.n30 VN.n29 17.3721
R48 VN.n36 VN.n35 17.3721
R49 VN.n28 VN.n27 12.3513
R50 VN.n5 VN.n4 12.3513
R51 VN.n14 VN.n13 7.09593
R52 VN.n37 VN.n36 7.09593
R53 VN.n21 VN.n20 3.18121
R54 VN.n44 VN.n43 3.18121
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VTAIL.n566 VTAIL.n565 756.745
R75 VTAIL.n70 VTAIL.n69 756.745
R76 VTAIL.n140 VTAIL.n139 756.745
R77 VTAIL.n212 VTAIL.n211 756.745
R78 VTAIL.n496 VTAIL.n495 756.745
R79 VTAIL.n424 VTAIL.n423 756.745
R80 VTAIL.n354 VTAIL.n353 756.745
R81 VTAIL.n282 VTAIL.n281 756.745
R82 VTAIL.n520 VTAIL.n519 585
R83 VTAIL.n525 VTAIL.n524 585
R84 VTAIL.n527 VTAIL.n526 585
R85 VTAIL.n516 VTAIL.n515 585
R86 VTAIL.n533 VTAIL.n532 585
R87 VTAIL.n535 VTAIL.n534 585
R88 VTAIL.n512 VTAIL.n511 585
R89 VTAIL.n541 VTAIL.n540 585
R90 VTAIL.n543 VTAIL.n542 585
R91 VTAIL.n508 VTAIL.n507 585
R92 VTAIL.n549 VTAIL.n548 585
R93 VTAIL.n551 VTAIL.n550 585
R94 VTAIL.n504 VTAIL.n503 585
R95 VTAIL.n557 VTAIL.n556 585
R96 VTAIL.n559 VTAIL.n558 585
R97 VTAIL.n500 VTAIL.n499 585
R98 VTAIL.n565 VTAIL.n564 585
R99 VTAIL.n24 VTAIL.n23 585
R100 VTAIL.n29 VTAIL.n28 585
R101 VTAIL.n31 VTAIL.n30 585
R102 VTAIL.n20 VTAIL.n19 585
R103 VTAIL.n37 VTAIL.n36 585
R104 VTAIL.n39 VTAIL.n38 585
R105 VTAIL.n16 VTAIL.n15 585
R106 VTAIL.n45 VTAIL.n44 585
R107 VTAIL.n47 VTAIL.n46 585
R108 VTAIL.n12 VTAIL.n11 585
R109 VTAIL.n53 VTAIL.n52 585
R110 VTAIL.n55 VTAIL.n54 585
R111 VTAIL.n8 VTAIL.n7 585
R112 VTAIL.n61 VTAIL.n60 585
R113 VTAIL.n63 VTAIL.n62 585
R114 VTAIL.n4 VTAIL.n3 585
R115 VTAIL.n69 VTAIL.n68 585
R116 VTAIL.n94 VTAIL.n93 585
R117 VTAIL.n99 VTAIL.n98 585
R118 VTAIL.n101 VTAIL.n100 585
R119 VTAIL.n90 VTAIL.n89 585
R120 VTAIL.n107 VTAIL.n106 585
R121 VTAIL.n109 VTAIL.n108 585
R122 VTAIL.n86 VTAIL.n85 585
R123 VTAIL.n115 VTAIL.n114 585
R124 VTAIL.n117 VTAIL.n116 585
R125 VTAIL.n82 VTAIL.n81 585
R126 VTAIL.n123 VTAIL.n122 585
R127 VTAIL.n125 VTAIL.n124 585
R128 VTAIL.n78 VTAIL.n77 585
R129 VTAIL.n131 VTAIL.n130 585
R130 VTAIL.n133 VTAIL.n132 585
R131 VTAIL.n74 VTAIL.n73 585
R132 VTAIL.n139 VTAIL.n138 585
R133 VTAIL.n166 VTAIL.n165 585
R134 VTAIL.n171 VTAIL.n170 585
R135 VTAIL.n173 VTAIL.n172 585
R136 VTAIL.n162 VTAIL.n161 585
R137 VTAIL.n179 VTAIL.n178 585
R138 VTAIL.n181 VTAIL.n180 585
R139 VTAIL.n158 VTAIL.n157 585
R140 VTAIL.n187 VTAIL.n186 585
R141 VTAIL.n189 VTAIL.n188 585
R142 VTAIL.n154 VTAIL.n153 585
R143 VTAIL.n195 VTAIL.n194 585
R144 VTAIL.n197 VTAIL.n196 585
R145 VTAIL.n150 VTAIL.n149 585
R146 VTAIL.n203 VTAIL.n202 585
R147 VTAIL.n205 VTAIL.n204 585
R148 VTAIL.n146 VTAIL.n145 585
R149 VTAIL.n211 VTAIL.n210 585
R150 VTAIL.n495 VTAIL.n494 585
R151 VTAIL.n430 VTAIL.n429 585
R152 VTAIL.n489 VTAIL.n488 585
R153 VTAIL.n487 VTAIL.n486 585
R154 VTAIL.n434 VTAIL.n433 585
R155 VTAIL.n481 VTAIL.n480 585
R156 VTAIL.n479 VTAIL.n478 585
R157 VTAIL.n438 VTAIL.n437 585
R158 VTAIL.n473 VTAIL.n472 585
R159 VTAIL.n471 VTAIL.n470 585
R160 VTAIL.n442 VTAIL.n441 585
R161 VTAIL.n465 VTAIL.n464 585
R162 VTAIL.n463 VTAIL.n462 585
R163 VTAIL.n446 VTAIL.n445 585
R164 VTAIL.n457 VTAIL.n456 585
R165 VTAIL.n455 VTAIL.n454 585
R166 VTAIL.n450 VTAIL.n449 585
R167 VTAIL.n423 VTAIL.n422 585
R168 VTAIL.n358 VTAIL.n357 585
R169 VTAIL.n417 VTAIL.n416 585
R170 VTAIL.n415 VTAIL.n414 585
R171 VTAIL.n362 VTAIL.n361 585
R172 VTAIL.n409 VTAIL.n408 585
R173 VTAIL.n407 VTAIL.n406 585
R174 VTAIL.n366 VTAIL.n365 585
R175 VTAIL.n401 VTAIL.n400 585
R176 VTAIL.n399 VTAIL.n398 585
R177 VTAIL.n370 VTAIL.n369 585
R178 VTAIL.n393 VTAIL.n392 585
R179 VTAIL.n391 VTAIL.n390 585
R180 VTAIL.n374 VTAIL.n373 585
R181 VTAIL.n385 VTAIL.n384 585
R182 VTAIL.n383 VTAIL.n382 585
R183 VTAIL.n378 VTAIL.n377 585
R184 VTAIL.n353 VTAIL.n352 585
R185 VTAIL.n288 VTAIL.n287 585
R186 VTAIL.n347 VTAIL.n346 585
R187 VTAIL.n345 VTAIL.n344 585
R188 VTAIL.n292 VTAIL.n291 585
R189 VTAIL.n339 VTAIL.n338 585
R190 VTAIL.n337 VTAIL.n336 585
R191 VTAIL.n296 VTAIL.n295 585
R192 VTAIL.n331 VTAIL.n330 585
R193 VTAIL.n329 VTAIL.n328 585
R194 VTAIL.n300 VTAIL.n299 585
R195 VTAIL.n323 VTAIL.n322 585
R196 VTAIL.n321 VTAIL.n320 585
R197 VTAIL.n304 VTAIL.n303 585
R198 VTAIL.n315 VTAIL.n314 585
R199 VTAIL.n313 VTAIL.n312 585
R200 VTAIL.n308 VTAIL.n307 585
R201 VTAIL.n281 VTAIL.n280 585
R202 VTAIL.n216 VTAIL.n215 585
R203 VTAIL.n275 VTAIL.n274 585
R204 VTAIL.n273 VTAIL.n272 585
R205 VTAIL.n220 VTAIL.n219 585
R206 VTAIL.n267 VTAIL.n266 585
R207 VTAIL.n265 VTAIL.n264 585
R208 VTAIL.n224 VTAIL.n223 585
R209 VTAIL.n259 VTAIL.n258 585
R210 VTAIL.n257 VTAIL.n256 585
R211 VTAIL.n228 VTAIL.n227 585
R212 VTAIL.n251 VTAIL.n250 585
R213 VTAIL.n249 VTAIL.n248 585
R214 VTAIL.n232 VTAIL.n231 585
R215 VTAIL.n243 VTAIL.n242 585
R216 VTAIL.n241 VTAIL.n240 585
R217 VTAIL.n236 VTAIL.n235 585
R218 VTAIL.n521 VTAIL.t13 327.466
R219 VTAIL.n25 VTAIL.t12 327.466
R220 VTAIL.n95 VTAIL.t1 327.466
R221 VTAIL.n167 VTAIL.t0 327.466
R222 VTAIL.n451 VTAIL.t3 327.466
R223 VTAIL.n379 VTAIL.t2 327.466
R224 VTAIL.n309 VTAIL.t9 327.466
R225 VTAIL.n237 VTAIL.t15 327.466
R226 VTAIL.n525 VTAIL.n519 171.744
R227 VTAIL.n526 VTAIL.n525 171.744
R228 VTAIL.n526 VTAIL.n515 171.744
R229 VTAIL.n533 VTAIL.n515 171.744
R230 VTAIL.n534 VTAIL.n533 171.744
R231 VTAIL.n534 VTAIL.n511 171.744
R232 VTAIL.n541 VTAIL.n511 171.744
R233 VTAIL.n542 VTAIL.n541 171.744
R234 VTAIL.n542 VTAIL.n507 171.744
R235 VTAIL.n549 VTAIL.n507 171.744
R236 VTAIL.n550 VTAIL.n549 171.744
R237 VTAIL.n550 VTAIL.n503 171.744
R238 VTAIL.n557 VTAIL.n503 171.744
R239 VTAIL.n558 VTAIL.n557 171.744
R240 VTAIL.n558 VTAIL.n499 171.744
R241 VTAIL.n565 VTAIL.n499 171.744
R242 VTAIL.n29 VTAIL.n23 171.744
R243 VTAIL.n30 VTAIL.n29 171.744
R244 VTAIL.n30 VTAIL.n19 171.744
R245 VTAIL.n37 VTAIL.n19 171.744
R246 VTAIL.n38 VTAIL.n37 171.744
R247 VTAIL.n38 VTAIL.n15 171.744
R248 VTAIL.n45 VTAIL.n15 171.744
R249 VTAIL.n46 VTAIL.n45 171.744
R250 VTAIL.n46 VTAIL.n11 171.744
R251 VTAIL.n53 VTAIL.n11 171.744
R252 VTAIL.n54 VTAIL.n53 171.744
R253 VTAIL.n54 VTAIL.n7 171.744
R254 VTAIL.n61 VTAIL.n7 171.744
R255 VTAIL.n62 VTAIL.n61 171.744
R256 VTAIL.n62 VTAIL.n3 171.744
R257 VTAIL.n69 VTAIL.n3 171.744
R258 VTAIL.n99 VTAIL.n93 171.744
R259 VTAIL.n100 VTAIL.n99 171.744
R260 VTAIL.n100 VTAIL.n89 171.744
R261 VTAIL.n107 VTAIL.n89 171.744
R262 VTAIL.n108 VTAIL.n107 171.744
R263 VTAIL.n108 VTAIL.n85 171.744
R264 VTAIL.n115 VTAIL.n85 171.744
R265 VTAIL.n116 VTAIL.n115 171.744
R266 VTAIL.n116 VTAIL.n81 171.744
R267 VTAIL.n123 VTAIL.n81 171.744
R268 VTAIL.n124 VTAIL.n123 171.744
R269 VTAIL.n124 VTAIL.n77 171.744
R270 VTAIL.n131 VTAIL.n77 171.744
R271 VTAIL.n132 VTAIL.n131 171.744
R272 VTAIL.n132 VTAIL.n73 171.744
R273 VTAIL.n139 VTAIL.n73 171.744
R274 VTAIL.n171 VTAIL.n165 171.744
R275 VTAIL.n172 VTAIL.n171 171.744
R276 VTAIL.n172 VTAIL.n161 171.744
R277 VTAIL.n179 VTAIL.n161 171.744
R278 VTAIL.n180 VTAIL.n179 171.744
R279 VTAIL.n180 VTAIL.n157 171.744
R280 VTAIL.n187 VTAIL.n157 171.744
R281 VTAIL.n188 VTAIL.n187 171.744
R282 VTAIL.n188 VTAIL.n153 171.744
R283 VTAIL.n195 VTAIL.n153 171.744
R284 VTAIL.n196 VTAIL.n195 171.744
R285 VTAIL.n196 VTAIL.n149 171.744
R286 VTAIL.n203 VTAIL.n149 171.744
R287 VTAIL.n204 VTAIL.n203 171.744
R288 VTAIL.n204 VTAIL.n145 171.744
R289 VTAIL.n211 VTAIL.n145 171.744
R290 VTAIL.n495 VTAIL.n429 171.744
R291 VTAIL.n488 VTAIL.n429 171.744
R292 VTAIL.n488 VTAIL.n487 171.744
R293 VTAIL.n487 VTAIL.n433 171.744
R294 VTAIL.n480 VTAIL.n433 171.744
R295 VTAIL.n480 VTAIL.n479 171.744
R296 VTAIL.n479 VTAIL.n437 171.744
R297 VTAIL.n472 VTAIL.n437 171.744
R298 VTAIL.n472 VTAIL.n471 171.744
R299 VTAIL.n471 VTAIL.n441 171.744
R300 VTAIL.n464 VTAIL.n441 171.744
R301 VTAIL.n464 VTAIL.n463 171.744
R302 VTAIL.n463 VTAIL.n445 171.744
R303 VTAIL.n456 VTAIL.n445 171.744
R304 VTAIL.n456 VTAIL.n455 171.744
R305 VTAIL.n455 VTAIL.n449 171.744
R306 VTAIL.n423 VTAIL.n357 171.744
R307 VTAIL.n416 VTAIL.n357 171.744
R308 VTAIL.n416 VTAIL.n415 171.744
R309 VTAIL.n415 VTAIL.n361 171.744
R310 VTAIL.n408 VTAIL.n361 171.744
R311 VTAIL.n408 VTAIL.n407 171.744
R312 VTAIL.n407 VTAIL.n365 171.744
R313 VTAIL.n400 VTAIL.n365 171.744
R314 VTAIL.n400 VTAIL.n399 171.744
R315 VTAIL.n399 VTAIL.n369 171.744
R316 VTAIL.n392 VTAIL.n369 171.744
R317 VTAIL.n392 VTAIL.n391 171.744
R318 VTAIL.n391 VTAIL.n373 171.744
R319 VTAIL.n384 VTAIL.n373 171.744
R320 VTAIL.n384 VTAIL.n383 171.744
R321 VTAIL.n383 VTAIL.n377 171.744
R322 VTAIL.n353 VTAIL.n287 171.744
R323 VTAIL.n346 VTAIL.n287 171.744
R324 VTAIL.n346 VTAIL.n345 171.744
R325 VTAIL.n345 VTAIL.n291 171.744
R326 VTAIL.n338 VTAIL.n291 171.744
R327 VTAIL.n338 VTAIL.n337 171.744
R328 VTAIL.n337 VTAIL.n295 171.744
R329 VTAIL.n330 VTAIL.n295 171.744
R330 VTAIL.n330 VTAIL.n329 171.744
R331 VTAIL.n329 VTAIL.n299 171.744
R332 VTAIL.n322 VTAIL.n299 171.744
R333 VTAIL.n322 VTAIL.n321 171.744
R334 VTAIL.n321 VTAIL.n303 171.744
R335 VTAIL.n314 VTAIL.n303 171.744
R336 VTAIL.n314 VTAIL.n313 171.744
R337 VTAIL.n313 VTAIL.n307 171.744
R338 VTAIL.n281 VTAIL.n215 171.744
R339 VTAIL.n274 VTAIL.n215 171.744
R340 VTAIL.n274 VTAIL.n273 171.744
R341 VTAIL.n273 VTAIL.n219 171.744
R342 VTAIL.n266 VTAIL.n219 171.744
R343 VTAIL.n266 VTAIL.n265 171.744
R344 VTAIL.n265 VTAIL.n223 171.744
R345 VTAIL.n258 VTAIL.n223 171.744
R346 VTAIL.n258 VTAIL.n257 171.744
R347 VTAIL.n257 VTAIL.n227 171.744
R348 VTAIL.n250 VTAIL.n227 171.744
R349 VTAIL.n250 VTAIL.n249 171.744
R350 VTAIL.n249 VTAIL.n231 171.744
R351 VTAIL.n242 VTAIL.n231 171.744
R352 VTAIL.n242 VTAIL.n241 171.744
R353 VTAIL.n241 VTAIL.n235 171.744
R354 VTAIL.t13 VTAIL.n519 85.8723
R355 VTAIL.t12 VTAIL.n23 85.8723
R356 VTAIL.t1 VTAIL.n93 85.8723
R357 VTAIL.t0 VTAIL.n165 85.8723
R358 VTAIL.t3 VTAIL.n449 85.8723
R359 VTAIL.t2 VTAIL.n377 85.8723
R360 VTAIL.t9 VTAIL.n307 85.8723
R361 VTAIL.t15 VTAIL.n235 85.8723
R362 VTAIL.n427 VTAIL.n426 58.4982
R363 VTAIL.n285 VTAIL.n284 58.4982
R364 VTAIL.n1 VTAIL.n0 58.4972
R365 VTAIL.n143 VTAIL.n142 58.4972
R366 VTAIL.n567 VTAIL.n566 34.3187
R367 VTAIL.n71 VTAIL.n70 34.3187
R368 VTAIL.n141 VTAIL.n140 34.3187
R369 VTAIL.n213 VTAIL.n212 34.3187
R370 VTAIL.n497 VTAIL.n496 34.3187
R371 VTAIL.n425 VTAIL.n424 34.3187
R372 VTAIL.n355 VTAIL.n354 34.3187
R373 VTAIL.n283 VTAIL.n282 34.3187
R374 VTAIL.n567 VTAIL.n497 25.1427
R375 VTAIL.n283 VTAIL.n213 25.1427
R376 VTAIL.n521 VTAIL.n520 16.3895
R377 VTAIL.n25 VTAIL.n24 16.3895
R378 VTAIL.n95 VTAIL.n94 16.3895
R379 VTAIL.n167 VTAIL.n166 16.3895
R380 VTAIL.n451 VTAIL.n450 16.3895
R381 VTAIL.n379 VTAIL.n378 16.3895
R382 VTAIL.n309 VTAIL.n308 16.3895
R383 VTAIL.n237 VTAIL.n236 16.3895
R384 VTAIL.n524 VTAIL.n523 12.8005
R385 VTAIL.n564 VTAIL.n498 12.8005
R386 VTAIL.n28 VTAIL.n27 12.8005
R387 VTAIL.n68 VTAIL.n2 12.8005
R388 VTAIL.n98 VTAIL.n97 12.8005
R389 VTAIL.n138 VTAIL.n72 12.8005
R390 VTAIL.n170 VTAIL.n169 12.8005
R391 VTAIL.n210 VTAIL.n144 12.8005
R392 VTAIL.n494 VTAIL.n428 12.8005
R393 VTAIL.n454 VTAIL.n453 12.8005
R394 VTAIL.n422 VTAIL.n356 12.8005
R395 VTAIL.n382 VTAIL.n381 12.8005
R396 VTAIL.n352 VTAIL.n286 12.8005
R397 VTAIL.n312 VTAIL.n311 12.8005
R398 VTAIL.n280 VTAIL.n214 12.8005
R399 VTAIL.n240 VTAIL.n239 12.8005
R400 VTAIL.n527 VTAIL.n518 12.0247
R401 VTAIL.n563 VTAIL.n500 12.0247
R402 VTAIL.n31 VTAIL.n22 12.0247
R403 VTAIL.n67 VTAIL.n4 12.0247
R404 VTAIL.n101 VTAIL.n92 12.0247
R405 VTAIL.n137 VTAIL.n74 12.0247
R406 VTAIL.n173 VTAIL.n164 12.0247
R407 VTAIL.n209 VTAIL.n146 12.0247
R408 VTAIL.n493 VTAIL.n430 12.0247
R409 VTAIL.n457 VTAIL.n448 12.0247
R410 VTAIL.n421 VTAIL.n358 12.0247
R411 VTAIL.n385 VTAIL.n376 12.0247
R412 VTAIL.n351 VTAIL.n288 12.0247
R413 VTAIL.n315 VTAIL.n306 12.0247
R414 VTAIL.n279 VTAIL.n216 12.0247
R415 VTAIL.n243 VTAIL.n234 12.0247
R416 VTAIL.n528 VTAIL.n516 11.249
R417 VTAIL.n560 VTAIL.n559 11.249
R418 VTAIL.n32 VTAIL.n20 11.249
R419 VTAIL.n64 VTAIL.n63 11.249
R420 VTAIL.n102 VTAIL.n90 11.249
R421 VTAIL.n134 VTAIL.n133 11.249
R422 VTAIL.n174 VTAIL.n162 11.249
R423 VTAIL.n206 VTAIL.n205 11.249
R424 VTAIL.n490 VTAIL.n489 11.249
R425 VTAIL.n458 VTAIL.n446 11.249
R426 VTAIL.n418 VTAIL.n417 11.249
R427 VTAIL.n386 VTAIL.n374 11.249
R428 VTAIL.n348 VTAIL.n347 11.249
R429 VTAIL.n316 VTAIL.n304 11.249
R430 VTAIL.n276 VTAIL.n275 11.249
R431 VTAIL.n244 VTAIL.n232 11.249
R432 VTAIL.n532 VTAIL.n531 10.4732
R433 VTAIL.n556 VTAIL.n502 10.4732
R434 VTAIL.n36 VTAIL.n35 10.4732
R435 VTAIL.n60 VTAIL.n6 10.4732
R436 VTAIL.n106 VTAIL.n105 10.4732
R437 VTAIL.n130 VTAIL.n76 10.4732
R438 VTAIL.n178 VTAIL.n177 10.4732
R439 VTAIL.n202 VTAIL.n148 10.4732
R440 VTAIL.n486 VTAIL.n432 10.4732
R441 VTAIL.n462 VTAIL.n461 10.4732
R442 VTAIL.n414 VTAIL.n360 10.4732
R443 VTAIL.n390 VTAIL.n389 10.4732
R444 VTAIL.n344 VTAIL.n290 10.4732
R445 VTAIL.n320 VTAIL.n319 10.4732
R446 VTAIL.n272 VTAIL.n218 10.4732
R447 VTAIL.n248 VTAIL.n247 10.4732
R448 VTAIL.n535 VTAIL.n514 9.69747
R449 VTAIL.n555 VTAIL.n504 9.69747
R450 VTAIL.n39 VTAIL.n18 9.69747
R451 VTAIL.n59 VTAIL.n8 9.69747
R452 VTAIL.n109 VTAIL.n88 9.69747
R453 VTAIL.n129 VTAIL.n78 9.69747
R454 VTAIL.n181 VTAIL.n160 9.69747
R455 VTAIL.n201 VTAIL.n150 9.69747
R456 VTAIL.n485 VTAIL.n434 9.69747
R457 VTAIL.n465 VTAIL.n444 9.69747
R458 VTAIL.n413 VTAIL.n362 9.69747
R459 VTAIL.n393 VTAIL.n372 9.69747
R460 VTAIL.n343 VTAIL.n292 9.69747
R461 VTAIL.n323 VTAIL.n302 9.69747
R462 VTAIL.n271 VTAIL.n220 9.69747
R463 VTAIL.n251 VTAIL.n230 9.69747
R464 VTAIL.n562 VTAIL.n498 9.45567
R465 VTAIL.n66 VTAIL.n2 9.45567
R466 VTAIL.n136 VTAIL.n72 9.45567
R467 VTAIL.n208 VTAIL.n144 9.45567
R468 VTAIL.n492 VTAIL.n428 9.45567
R469 VTAIL.n420 VTAIL.n356 9.45567
R470 VTAIL.n350 VTAIL.n286 9.45567
R471 VTAIL.n278 VTAIL.n214 9.45567
R472 VTAIL.n545 VTAIL.n544 9.3005
R473 VTAIL.n547 VTAIL.n546 9.3005
R474 VTAIL.n506 VTAIL.n505 9.3005
R475 VTAIL.n553 VTAIL.n552 9.3005
R476 VTAIL.n555 VTAIL.n554 9.3005
R477 VTAIL.n502 VTAIL.n501 9.3005
R478 VTAIL.n561 VTAIL.n560 9.3005
R479 VTAIL.n563 VTAIL.n562 9.3005
R480 VTAIL.n539 VTAIL.n538 9.3005
R481 VTAIL.n537 VTAIL.n536 9.3005
R482 VTAIL.n514 VTAIL.n513 9.3005
R483 VTAIL.n531 VTAIL.n530 9.3005
R484 VTAIL.n529 VTAIL.n528 9.3005
R485 VTAIL.n518 VTAIL.n517 9.3005
R486 VTAIL.n523 VTAIL.n522 9.3005
R487 VTAIL.n510 VTAIL.n509 9.3005
R488 VTAIL.n49 VTAIL.n48 9.3005
R489 VTAIL.n51 VTAIL.n50 9.3005
R490 VTAIL.n10 VTAIL.n9 9.3005
R491 VTAIL.n57 VTAIL.n56 9.3005
R492 VTAIL.n59 VTAIL.n58 9.3005
R493 VTAIL.n6 VTAIL.n5 9.3005
R494 VTAIL.n65 VTAIL.n64 9.3005
R495 VTAIL.n67 VTAIL.n66 9.3005
R496 VTAIL.n43 VTAIL.n42 9.3005
R497 VTAIL.n41 VTAIL.n40 9.3005
R498 VTAIL.n18 VTAIL.n17 9.3005
R499 VTAIL.n35 VTAIL.n34 9.3005
R500 VTAIL.n33 VTAIL.n32 9.3005
R501 VTAIL.n22 VTAIL.n21 9.3005
R502 VTAIL.n27 VTAIL.n26 9.3005
R503 VTAIL.n14 VTAIL.n13 9.3005
R504 VTAIL.n119 VTAIL.n118 9.3005
R505 VTAIL.n121 VTAIL.n120 9.3005
R506 VTAIL.n80 VTAIL.n79 9.3005
R507 VTAIL.n127 VTAIL.n126 9.3005
R508 VTAIL.n129 VTAIL.n128 9.3005
R509 VTAIL.n76 VTAIL.n75 9.3005
R510 VTAIL.n135 VTAIL.n134 9.3005
R511 VTAIL.n137 VTAIL.n136 9.3005
R512 VTAIL.n113 VTAIL.n112 9.3005
R513 VTAIL.n111 VTAIL.n110 9.3005
R514 VTAIL.n88 VTAIL.n87 9.3005
R515 VTAIL.n105 VTAIL.n104 9.3005
R516 VTAIL.n103 VTAIL.n102 9.3005
R517 VTAIL.n92 VTAIL.n91 9.3005
R518 VTAIL.n97 VTAIL.n96 9.3005
R519 VTAIL.n84 VTAIL.n83 9.3005
R520 VTAIL.n191 VTAIL.n190 9.3005
R521 VTAIL.n193 VTAIL.n192 9.3005
R522 VTAIL.n152 VTAIL.n151 9.3005
R523 VTAIL.n199 VTAIL.n198 9.3005
R524 VTAIL.n201 VTAIL.n200 9.3005
R525 VTAIL.n148 VTAIL.n147 9.3005
R526 VTAIL.n207 VTAIL.n206 9.3005
R527 VTAIL.n209 VTAIL.n208 9.3005
R528 VTAIL.n185 VTAIL.n184 9.3005
R529 VTAIL.n183 VTAIL.n182 9.3005
R530 VTAIL.n160 VTAIL.n159 9.3005
R531 VTAIL.n177 VTAIL.n176 9.3005
R532 VTAIL.n175 VTAIL.n174 9.3005
R533 VTAIL.n164 VTAIL.n163 9.3005
R534 VTAIL.n169 VTAIL.n168 9.3005
R535 VTAIL.n156 VTAIL.n155 9.3005
R536 VTAIL.n493 VTAIL.n492 9.3005
R537 VTAIL.n491 VTAIL.n490 9.3005
R538 VTAIL.n432 VTAIL.n431 9.3005
R539 VTAIL.n485 VTAIL.n484 9.3005
R540 VTAIL.n483 VTAIL.n482 9.3005
R541 VTAIL.n436 VTAIL.n435 9.3005
R542 VTAIL.n477 VTAIL.n476 9.3005
R543 VTAIL.n475 VTAIL.n474 9.3005
R544 VTAIL.n440 VTAIL.n439 9.3005
R545 VTAIL.n469 VTAIL.n468 9.3005
R546 VTAIL.n467 VTAIL.n466 9.3005
R547 VTAIL.n444 VTAIL.n443 9.3005
R548 VTAIL.n461 VTAIL.n460 9.3005
R549 VTAIL.n459 VTAIL.n458 9.3005
R550 VTAIL.n448 VTAIL.n447 9.3005
R551 VTAIL.n453 VTAIL.n452 9.3005
R552 VTAIL.n405 VTAIL.n404 9.3005
R553 VTAIL.n364 VTAIL.n363 9.3005
R554 VTAIL.n411 VTAIL.n410 9.3005
R555 VTAIL.n413 VTAIL.n412 9.3005
R556 VTAIL.n360 VTAIL.n359 9.3005
R557 VTAIL.n419 VTAIL.n418 9.3005
R558 VTAIL.n421 VTAIL.n420 9.3005
R559 VTAIL.n403 VTAIL.n402 9.3005
R560 VTAIL.n368 VTAIL.n367 9.3005
R561 VTAIL.n397 VTAIL.n396 9.3005
R562 VTAIL.n395 VTAIL.n394 9.3005
R563 VTAIL.n372 VTAIL.n371 9.3005
R564 VTAIL.n389 VTAIL.n388 9.3005
R565 VTAIL.n387 VTAIL.n386 9.3005
R566 VTAIL.n376 VTAIL.n375 9.3005
R567 VTAIL.n381 VTAIL.n380 9.3005
R568 VTAIL.n335 VTAIL.n334 9.3005
R569 VTAIL.n294 VTAIL.n293 9.3005
R570 VTAIL.n341 VTAIL.n340 9.3005
R571 VTAIL.n343 VTAIL.n342 9.3005
R572 VTAIL.n290 VTAIL.n289 9.3005
R573 VTAIL.n349 VTAIL.n348 9.3005
R574 VTAIL.n351 VTAIL.n350 9.3005
R575 VTAIL.n333 VTAIL.n332 9.3005
R576 VTAIL.n298 VTAIL.n297 9.3005
R577 VTAIL.n327 VTAIL.n326 9.3005
R578 VTAIL.n325 VTAIL.n324 9.3005
R579 VTAIL.n302 VTAIL.n301 9.3005
R580 VTAIL.n319 VTAIL.n318 9.3005
R581 VTAIL.n317 VTAIL.n316 9.3005
R582 VTAIL.n306 VTAIL.n305 9.3005
R583 VTAIL.n311 VTAIL.n310 9.3005
R584 VTAIL.n263 VTAIL.n262 9.3005
R585 VTAIL.n222 VTAIL.n221 9.3005
R586 VTAIL.n269 VTAIL.n268 9.3005
R587 VTAIL.n271 VTAIL.n270 9.3005
R588 VTAIL.n218 VTAIL.n217 9.3005
R589 VTAIL.n277 VTAIL.n276 9.3005
R590 VTAIL.n279 VTAIL.n278 9.3005
R591 VTAIL.n261 VTAIL.n260 9.3005
R592 VTAIL.n226 VTAIL.n225 9.3005
R593 VTAIL.n255 VTAIL.n254 9.3005
R594 VTAIL.n253 VTAIL.n252 9.3005
R595 VTAIL.n230 VTAIL.n229 9.3005
R596 VTAIL.n247 VTAIL.n246 9.3005
R597 VTAIL.n245 VTAIL.n244 9.3005
R598 VTAIL.n234 VTAIL.n233 9.3005
R599 VTAIL.n239 VTAIL.n238 9.3005
R600 VTAIL.n536 VTAIL.n512 8.92171
R601 VTAIL.n552 VTAIL.n551 8.92171
R602 VTAIL.n40 VTAIL.n16 8.92171
R603 VTAIL.n56 VTAIL.n55 8.92171
R604 VTAIL.n110 VTAIL.n86 8.92171
R605 VTAIL.n126 VTAIL.n125 8.92171
R606 VTAIL.n182 VTAIL.n158 8.92171
R607 VTAIL.n198 VTAIL.n197 8.92171
R608 VTAIL.n482 VTAIL.n481 8.92171
R609 VTAIL.n466 VTAIL.n442 8.92171
R610 VTAIL.n410 VTAIL.n409 8.92171
R611 VTAIL.n394 VTAIL.n370 8.92171
R612 VTAIL.n340 VTAIL.n339 8.92171
R613 VTAIL.n324 VTAIL.n300 8.92171
R614 VTAIL.n268 VTAIL.n267 8.92171
R615 VTAIL.n252 VTAIL.n228 8.92171
R616 VTAIL.n540 VTAIL.n539 8.14595
R617 VTAIL.n548 VTAIL.n506 8.14595
R618 VTAIL.n44 VTAIL.n43 8.14595
R619 VTAIL.n52 VTAIL.n10 8.14595
R620 VTAIL.n114 VTAIL.n113 8.14595
R621 VTAIL.n122 VTAIL.n80 8.14595
R622 VTAIL.n186 VTAIL.n185 8.14595
R623 VTAIL.n194 VTAIL.n152 8.14595
R624 VTAIL.n478 VTAIL.n436 8.14595
R625 VTAIL.n470 VTAIL.n469 8.14595
R626 VTAIL.n406 VTAIL.n364 8.14595
R627 VTAIL.n398 VTAIL.n397 8.14595
R628 VTAIL.n336 VTAIL.n294 8.14595
R629 VTAIL.n328 VTAIL.n327 8.14595
R630 VTAIL.n264 VTAIL.n222 8.14595
R631 VTAIL.n256 VTAIL.n255 8.14595
R632 VTAIL.n543 VTAIL.n510 7.3702
R633 VTAIL.n547 VTAIL.n508 7.3702
R634 VTAIL.n47 VTAIL.n14 7.3702
R635 VTAIL.n51 VTAIL.n12 7.3702
R636 VTAIL.n117 VTAIL.n84 7.3702
R637 VTAIL.n121 VTAIL.n82 7.3702
R638 VTAIL.n189 VTAIL.n156 7.3702
R639 VTAIL.n193 VTAIL.n154 7.3702
R640 VTAIL.n477 VTAIL.n438 7.3702
R641 VTAIL.n473 VTAIL.n440 7.3702
R642 VTAIL.n405 VTAIL.n366 7.3702
R643 VTAIL.n401 VTAIL.n368 7.3702
R644 VTAIL.n335 VTAIL.n296 7.3702
R645 VTAIL.n331 VTAIL.n298 7.3702
R646 VTAIL.n263 VTAIL.n224 7.3702
R647 VTAIL.n259 VTAIL.n226 7.3702
R648 VTAIL.n544 VTAIL.n543 6.59444
R649 VTAIL.n544 VTAIL.n508 6.59444
R650 VTAIL.n48 VTAIL.n47 6.59444
R651 VTAIL.n48 VTAIL.n12 6.59444
R652 VTAIL.n118 VTAIL.n117 6.59444
R653 VTAIL.n118 VTAIL.n82 6.59444
R654 VTAIL.n190 VTAIL.n189 6.59444
R655 VTAIL.n190 VTAIL.n154 6.59444
R656 VTAIL.n474 VTAIL.n438 6.59444
R657 VTAIL.n474 VTAIL.n473 6.59444
R658 VTAIL.n402 VTAIL.n366 6.59444
R659 VTAIL.n402 VTAIL.n401 6.59444
R660 VTAIL.n332 VTAIL.n296 6.59444
R661 VTAIL.n332 VTAIL.n331 6.59444
R662 VTAIL.n260 VTAIL.n224 6.59444
R663 VTAIL.n260 VTAIL.n259 6.59444
R664 VTAIL.n540 VTAIL.n510 5.81868
R665 VTAIL.n548 VTAIL.n547 5.81868
R666 VTAIL.n44 VTAIL.n14 5.81868
R667 VTAIL.n52 VTAIL.n51 5.81868
R668 VTAIL.n114 VTAIL.n84 5.81868
R669 VTAIL.n122 VTAIL.n121 5.81868
R670 VTAIL.n186 VTAIL.n156 5.81868
R671 VTAIL.n194 VTAIL.n193 5.81868
R672 VTAIL.n478 VTAIL.n477 5.81868
R673 VTAIL.n470 VTAIL.n440 5.81868
R674 VTAIL.n406 VTAIL.n405 5.81868
R675 VTAIL.n398 VTAIL.n368 5.81868
R676 VTAIL.n336 VTAIL.n335 5.81868
R677 VTAIL.n328 VTAIL.n298 5.81868
R678 VTAIL.n264 VTAIL.n263 5.81868
R679 VTAIL.n256 VTAIL.n226 5.81868
R680 VTAIL.n539 VTAIL.n512 5.04292
R681 VTAIL.n551 VTAIL.n506 5.04292
R682 VTAIL.n43 VTAIL.n16 5.04292
R683 VTAIL.n55 VTAIL.n10 5.04292
R684 VTAIL.n113 VTAIL.n86 5.04292
R685 VTAIL.n125 VTAIL.n80 5.04292
R686 VTAIL.n185 VTAIL.n158 5.04292
R687 VTAIL.n197 VTAIL.n152 5.04292
R688 VTAIL.n481 VTAIL.n436 5.04292
R689 VTAIL.n469 VTAIL.n442 5.04292
R690 VTAIL.n409 VTAIL.n364 5.04292
R691 VTAIL.n397 VTAIL.n370 5.04292
R692 VTAIL.n339 VTAIL.n294 5.04292
R693 VTAIL.n327 VTAIL.n300 5.04292
R694 VTAIL.n267 VTAIL.n222 5.04292
R695 VTAIL.n255 VTAIL.n228 5.04292
R696 VTAIL.n536 VTAIL.n535 4.26717
R697 VTAIL.n552 VTAIL.n504 4.26717
R698 VTAIL.n40 VTAIL.n39 4.26717
R699 VTAIL.n56 VTAIL.n8 4.26717
R700 VTAIL.n110 VTAIL.n109 4.26717
R701 VTAIL.n126 VTAIL.n78 4.26717
R702 VTAIL.n182 VTAIL.n181 4.26717
R703 VTAIL.n198 VTAIL.n150 4.26717
R704 VTAIL.n482 VTAIL.n434 4.26717
R705 VTAIL.n466 VTAIL.n465 4.26717
R706 VTAIL.n410 VTAIL.n362 4.26717
R707 VTAIL.n394 VTAIL.n393 4.26717
R708 VTAIL.n340 VTAIL.n292 4.26717
R709 VTAIL.n324 VTAIL.n323 4.26717
R710 VTAIL.n268 VTAIL.n220 4.26717
R711 VTAIL.n252 VTAIL.n251 4.26717
R712 VTAIL.n522 VTAIL.n521 3.70982
R713 VTAIL.n26 VTAIL.n25 3.70982
R714 VTAIL.n96 VTAIL.n95 3.70982
R715 VTAIL.n168 VTAIL.n167 3.70982
R716 VTAIL.n452 VTAIL.n451 3.70982
R717 VTAIL.n380 VTAIL.n379 3.70982
R718 VTAIL.n310 VTAIL.n309 3.70982
R719 VTAIL.n238 VTAIL.n237 3.70982
R720 VTAIL.n532 VTAIL.n514 3.49141
R721 VTAIL.n556 VTAIL.n555 3.49141
R722 VTAIL.n36 VTAIL.n18 3.49141
R723 VTAIL.n60 VTAIL.n59 3.49141
R724 VTAIL.n106 VTAIL.n88 3.49141
R725 VTAIL.n130 VTAIL.n129 3.49141
R726 VTAIL.n178 VTAIL.n160 3.49141
R727 VTAIL.n202 VTAIL.n201 3.49141
R728 VTAIL.n486 VTAIL.n485 3.49141
R729 VTAIL.n462 VTAIL.n444 3.49141
R730 VTAIL.n414 VTAIL.n413 3.49141
R731 VTAIL.n390 VTAIL.n372 3.49141
R732 VTAIL.n344 VTAIL.n343 3.49141
R733 VTAIL.n320 VTAIL.n302 3.49141
R734 VTAIL.n272 VTAIL.n271 3.49141
R735 VTAIL.n248 VTAIL.n230 3.49141
R736 VTAIL.n531 VTAIL.n516 2.71565
R737 VTAIL.n559 VTAIL.n502 2.71565
R738 VTAIL.n35 VTAIL.n20 2.71565
R739 VTAIL.n63 VTAIL.n6 2.71565
R740 VTAIL.n105 VTAIL.n90 2.71565
R741 VTAIL.n133 VTAIL.n76 2.71565
R742 VTAIL.n177 VTAIL.n162 2.71565
R743 VTAIL.n205 VTAIL.n148 2.71565
R744 VTAIL.n489 VTAIL.n432 2.71565
R745 VTAIL.n461 VTAIL.n446 2.71565
R746 VTAIL.n417 VTAIL.n360 2.71565
R747 VTAIL.n389 VTAIL.n374 2.71565
R748 VTAIL.n347 VTAIL.n290 2.71565
R749 VTAIL.n319 VTAIL.n304 2.71565
R750 VTAIL.n275 VTAIL.n218 2.71565
R751 VTAIL.n247 VTAIL.n232 2.71565
R752 VTAIL.n0 VTAIL.t8 2.57822
R753 VTAIL.n0 VTAIL.t14 2.57822
R754 VTAIL.n142 VTAIL.t4 2.57822
R755 VTAIL.n142 VTAIL.t5 2.57822
R756 VTAIL.n426 VTAIL.t6 2.57822
R757 VTAIL.n426 VTAIL.t7 2.57822
R758 VTAIL.n284 VTAIL.t11 2.57822
R759 VTAIL.n284 VTAIL.t10 2.57822
R760 VTAIL.n528 VTAIL.n527 1.93989
R761 VTAIL.n560 VTAIL.n500 1.93989
R762 VTAIL.n32 VTAIL.n31 1.93989
R763 VTAIL.n64 VTAIL.n4 1.93989
R764 VTAIL.n102 VTAIL.n101 1.93989
R765 VTAIL.n134 VTAIL.n74 1.93989
R766 VTAIL.n174 VTAIL.n173 1.93989
R767 VTAIL.n206 VTAIL.n146 1.93989
R768 VTAIL.n490 VTAIL.n430 1.93989
R769 VTAIL.n458 VTAIL.n457 1.93989
R770 VTAIL.n418 VTAIL.n358 1.93989
R771 VTAIL.n386 VTAIL.n385 1.93989
R772 VTAIL.n348 VTAIL.n288 1.93989
R773 VTAIL.n316 VTAIL.n315 1.93989
R774 VTAIL.n276 VTAIL.n216 1.93989
R775 VTAIL.n244 VTAIL.n243 1.93989
R776 VTAIL.n285 VTAIL.n283 1.90567
R777 VTAIL.n355 VTAIL.n285 1.90567
R778 VTAIL.n427 VTAIL.n425 1.90567
R779 VTAIL.n497 VTAIL.n427 1.90567
R780 VTAIL.n213 VTAIL.n143 1.90567
R781 VTAIL.n143 VTAIL.n141 1.90567
R782 VTAIL.n71 VTAIL.n1 1.90567
R783 VTAIL VTAIL.n567 1.84748
R784 VTAIL.n524 VTAIL.n518 1.16414
R785 VTAIL.n564 VTAIL.n563 1.16414
R786 VTAIL.n28 VTAIL.n22 1.16414
R787 VTAIL.n68 VTAIL.n67 1.16414
R788 VTAIL.n98 VTAIL.n92 1.16414
R789 VTAIL.n138 VTAIL.n137 1.16414
R790 VTAIL.n170 VTAIL.n164 1.16414
R791 VTAIL.n210 VTAIL.n209 1.16414
R792 VTAIL.n494 VTAIL.n493 1.16414
R793 VTAIL.n454 VTAIL.n448 1.16414
R794 VTAIL.n422 VTAIL.n421 1.16414
R795 VTAIL.n382 VTAIL.n376 1.16414
R796 VTAIL.n352 VTAIL.n351 1.16414
R797 VTAIL.n312 VTAIL.n306 1.16414
R798 VTAIL.n280 VTAIL.n279 1.16414
R799 VTAIL.n240 VTAIL.n234 1.16414
R800 VTAIL.n425 VTAIL.n355 0.470328
R801 VTAIL.n141 VTAIL.n71 0.470328
R802 VTAIL.n523 VTAIL.n520 0.388379
R803 VTAIL.n566 VTAIL.n498 0.388379
R804 VTAIL.n27 VTAIL.n24 0.388379
R805 VTAIL.n70 VTAIL.n2 0.388379
R806 VTAIL.n97 VTAIL.n94 0.388379
R807 VTAIL.n140 VTAIL.n72 0.388379
R808 VTAIL.n169 VTAIL.n166 0.388379
R809 VTAIL.n212 VTAIL.n144 0.388379
R810 VTAIL.n496 VTAIL.n428 0.388379
R811 VTAIL.n453 VTAIL.n450 0.388379
R812 VTAIL.n424 VTAIL.n356 0.388379
R813 VTAIL.n381 VTAIL.n378 0.388379
R814 VTAIL.n354 VTAIL.n286 0.388379
R815 VTAIL.n311 VTAIL.n308 0.388379
R816 VTAIL.n282 VTAIL.n214 0.388379
R817 VTAIL.n239 VTAIL.n236 0.388379
R818 VTAIL.n522 VTAIL.n517 0.155672
R819 VTAIL.n529 VTAIL.n517 0.155672
R820 VTAIL.n530 VTAIL.n529 0.155672
R821 VTAIL.n530 VTAIL.n513 0.155672
R822 VTAIL.n537 VTAIL.n513 0.155672
R823 VTAIL.n538 VTAIL.n537 0.155672
R824 VTAIL.n538 VTAIL.n509 0.155672
R825 VTAIL.n545 VTAIL.n509 0.155672
R826 VTAIL.n546 VTAIL.n545 0.155672
R827 VTAIL.n546 VTAIL.n505 0.155672
R828 VTAIL.n553 VTAIL.n505 0.155672
R829 VTAIL.n554 VTAIL.n553 0.155672
R830 VTAIL.n554 VTAIL.n501 0.155672
R831 VTAIL.n561 VTAIL.n501 0.155672
R832 VTAIL.n562 VTAIL.n561 0.155672
R833 VTAIL.n26 VTAIL.n21 0.155672
R834 VTAIL.n33 VTAIL.n21 0.155672
R835 VTAIL.n34 VTAIL.n33 0.155672
R836 VTAIL.n34 VTAIL.n17 0.155672
R837 VTAIL.n41 VTAIL.n17 0.155672
R838 VTAIL.n42 VTAIL.n41 0.155672
R839 VTAIL.n42 VTAIL.n13 0.155672
R840 VTAIL.n49 VTAIL.n13 0.155672
R841 VTAIL.n50 VTAIL.n49 0.155672
R842 VTAIL.n50 VTAIL.n9 0.155672
R843 VTAIL.n57 VTAIL.n9 0.155672
R844 VTAIL.n58 VTAIL.n57 0.155672
R845 VTAIL.n58 VTAIL.n5 0.155672
R846 VTAIL.n65 VTAIL.n5 0.155672
R847 VTAIL.n66 VTAIL.n65 0.155672
R848 VTAIL.n96 VTAIL.n91 0.155672
R849 VTAIL.n103 VTAIL.n91 0.155672
R850 VTAIL.n104 VTAIL.n103 0.155672
R851 VTAIL.n104 VTAIL.n87 0.155672
R852 VTAIL.n111 VTAIL.n87 0.155672
R853 VTAIL.n112 VTAIL.n111 0.155672
R854 VTAIL.n112 VTAIL.n83 0.155672
R855 VTAIL.n119 VTAIL.n83 0.155672
R856 VTAIL.n120 VTAIL.n119 0.155672
R857 VTAIL.n120 VTAIL.n79 0.155672
R858 VTAIL.n127 VTAIL.n79 0.155672
R859 VTAIL.n128 VTAIL.n127 0.155672
R860 VTAIL.n128 VTAIL.n75 0.155672
R861 VTAIL.n135 VTAIL.n75 0.155672
R862 VTAIL.n136 VTAIL.n135 0.155672
R863 VTAIL.n168 VTAIL.n163 0.155672
R864 VTAIL.n175 VTAIL.n163 0.155672
R865 VTAIL.n176 VTAIL.n175 0.155672
R866 VTAIL.n176 VTAIL.n159 0.155672
R867 VTAIL.n183 VTAIL.n159 0.155672
R868 VTAIL.n184 VTAIL.n183 0.155672
R869 VTAIL.n184 VTAIL.n155 0.155672
R870 VTAIL.n191 VTAIL.n155 0.155672
R871 VTAIL.n192 VTAIL.n191 0.155672
R872 VTAIL.n192 VTAIL.n151 0.155672
R873 VTAIL.n199 VTAIL.n151 0.155672
R874 VTAIL.n200 VTAIL.n199 0.155672
R875 VTAIL.n200 VTAIL.n147 0.155672
R876 VTAIL.n207 VTAIL.n147 0.155672
R877 VTAIL.n208 VTAIL.n207 0.155672
R878 VTAIL.n492 VTAIL.n491 0.155672
R879 VTAIL.n491 VTAIL.n431 0.155672
R880 VTAIL.n484 VTAIL.n431 0.155672
R881 VTAIL.n484 VTAIL.n483 0.155672
R882 VTAIL.n483 VTAIL.n435 0.155672
R883 VTAIL.n476 VTAIL.n435 0.155672
R884 VTAIL.n476 VTAIL.n475 0.155672
R885 VTAIL.n475 VTAIL.n439 0.155672
R886 VTAIL.n468 VTAIL.n439 0.155672
R887 VTAIL.n468 VTAIL.n467 0.155672
R888 VTAIL.n467 VTAIL.n443 0.155672
R889 VTAIL.n460 VTAIL.n443 0.155672
R890 VTAIL.n460 VTAIL.n459 0.155672
R891 VTAIL.n459 VTAIL.n447 0.155672
R892 VTAIL.n452 VTAIL.n447 0.155672
R893 VTAIL.n420 VTAIL.n419 0.155672
R894 VTAIL.n419 VTAIL.n359 0.155672
R895 VTAIL.n412 VTAIL.n359 0.155672
R896 VTAIL.n412 VTAIL.n411 0.155672
R897 VTAIL.n411 VTAIL.n363 0.155672
R898 VTAIL.n404 VTAIL.n363 0.155672
R899 VTAIL.n404 VTAIL.n403 0.155672
R900 VTAIL.n403 VTAIL.n367 0.155672
R901 VTAIL.n396 VTAIL.n367 0.155672
R902 VTAIL.n396 VTAIL.n395 0.155672
R903 VTAIL.n395 VTAIL.n371 0.155672
R904 VTAIL.n388 VTAIL.n371 0.155672
R905 VTAIL.n388 VTAIL.n387 0.155672
R906 VTAIL.n387 VTAIL.n375 0.155672
R907 VTAIL.n380 VTAIL.n375 0.155672
R908 VTAIL.n350 VTAIL.n349 0.155672
R909 VTAIL.n349 VTAIL.n289 0.155672
R910 VTAIL.n342 VTAIL.n289 0.155672
R911 VTAIL.n342 VTAIL.n341 0.155672
R912 VTAIL.n341 VTAIL.n293 0.155672
R913 VTAIL.n334 VTAIL.n293 0.155672
R914 VTAIL.n334 VTAIL.n333 0.155672
R915 VTAIL.n333 VTAIL.n297 0.155672
R916 VTAIL.n326 VTAIL.n297 0.155672
R917 VTAIL.n326 VTAIL.n325 0.155672
R918 VTAIL.n325 VTAIL.n301 0.155672
R919 VTAIL.n318 VTAIL.n301 0.155672
R920 VTAIL.n318 VTAIL.n317 0.155672
R921 VTAIL.n317 VTAIL.n305 0.155672
R922 VTAIL.n310 VTAIL.n305 0.155672
R923 VTAIL.n278 VTAIL.n277 0.155672
R924 VTAIL.n277 VTAIL.n217 0.155672
R925 VTAIL.n270 VTAIL.n217 0.155672
R926 VTAIL.n270 VTAIL.n269 0.155672
R927 VTAIL.n269 VTAIL.n221 0.155672
R928 VTAIL.n262 VTAIL.n221 0.155672
R929 VTAIL.n262 VTAIL.n261 0.155672
R930 VTAIL.n261 VTAIL.n225 0.155672
R931 VTAIL.n254 VTAIL.n225 0.155672
R932 VTAIL.n254 VTAIL.n253 0.155672
R933 VTAIL.n253 VTAIL.n229 0.155672
R934 VTAIL.n246 VTAIL.n229 0.155672
R935 VTAIL.n246 VTAIL.n245 0.155672
R936 VTAIL.n245 VTAIL.n233 0.155672
R937 VTAIL.n238 VTAIL.n233 0.155672
R938 VTAIL VTAIL.n1 0.0586897
R939 VDD2.n2 VDD2.n1 76.0732
R940 VDD2.n2 VDD2.n0 76.0732
R941 VDD2 VDD2.n5 76.0703
R942 VDD2.n4 VDD2.n3 75.177
R943 VDD2.n4 VDD2.n2 43.1593
R944 VDD2.n5 VDD2.t0 2.57822
R945 VDD2.n5 VDD2.t1 2.57822
R946 VDD2.n3 VDD2.t4 2.57822
R947 VDD2.n3 VDD2.t7 2.57822
R948 VDD2.n1 VDD2.t3 2.57822
R949 VDD2.n1 VDD2.t2 2.57822
R950 VDD2.n0 VDD2.t6 2.57822
R951 VDD2.n0 VDD2.t5 2.57822
R952 VDD2 VDD2.n4 1.01128
R953 VP.n13 VP.t7 195.512
R954 VP.n31 VP.n7 182.587
R955 VP.n56 VP.n55 182.587
R956 VP.n30 VP.n29 182.587
R957 VP.n7 VP.t6 161.649
R958 VP.n40 VP.t4 161.649
R959 VP.n47 VP.t2 161.649
R960 VP.n55 VP.t1 161.649
R961 VP.n29 VP.t5 161.649
R962 VP.n21 VP.t3 161.649
R963 VP.n14 VP.t0 161.649
R964 VP.n15 VP.n12 161.3
R965 VP.n17 VP.n16 161.3
R966 VP.n18 VP.n11 161.3
R967 VP.n20 VP.n19 161.3
R968 VP.n22 VP.n10 161.3
R969 VP.n24 VP.n23 161.3
R970 VP.n25 VP.n9 161.3
R971 VP.n27 VP.n26 161.3
R972 VP.n28 VP.n8 161.3
R973 VP.n54 VP.n0 161.3
R974 VP.n53 VP.n52 161.3
R975 VP.n51 VP.n1 161.3
R976 VP.n50 VP.n49 161.3
R977 VP.n48 VP.n2 161.3
R978 VP.n46 VP.n45 161.3
R979 VP.n44 VP.n3 161.3
R980 VP.n43 VP.n42 161.3
R981 VP.n41 VP.n4 161.3
R982 VP.n39 VP.n38 161.3
R983 VP.n37 VP.n5 161.3
R984 VP.n36 VP.n35 161.3
R985 VP.n34 VP.n6 161.3
R986 VP.n33 VP.n32 161.3
R987 VP.n42 VP.n3 56.5193
R988 VP.n16 VP.n11 56.5193
R989 VP.n14 VP.n13 52.3231
R990 VP.n31 VP.n30 47.902
R991 VP.n35 VP.n5 44.3785
R992 VP.n49 VP.n1 44.3785
R993 VP.n23 VP.n9 44.3785
R994 VP.n35 VP.n34 36.6083
R995 VP.n53 VP.n1 36.6083
R996 VP.n27 VP.n9 36.6083
R997 VP.n34 VP.n33 24.4675
R998 VP.n39 VP.n5 24.4675
R999 VP.n42 VP.n41 24.4675
R1000 VP.n46 VP.n3 24.4675
R1001 VP.n49 VP.n48 24.4675
R1002 VP.n54 VP.n53 24.4675
R1003 VP.n28 VP.n27 24.4675
R1004 VP.n20 VP.n11 24.4675
R1005 VP.n23 VP.n22 24.4675
R1006 VP.n16 VP.n15 24.4675
R1007 VP.n41 VP.n40 17.3721
R1008 VP.n47 VP.n46 17.3721
R1009 VP.n21 VP.n20 17.3721
R1010 VP.n15 VP.n14 17.3721
R1011 VP.n13 VP.n12 12.3512
R1012 VP.n40 VP.n39 7.09593
R1013 VP.n48 VP.n47 7.09593
R1014 VP.n22 VP.n21 7.09593
R1015 VP.n33 VP.n7 3.18121
R1016 VP.n55 VP.n54 3.18121
R1017 VP.n29 VP.n28 3.18121
R1018 VP.n17 VP.n12 0.189894
R1019 VP.n18 VP.n17 0.189894
R1020 VP.n19 VP.n18 0.189894
R1021 VP.n19 VP.n10 0.189894
R1022 VP.n24 VP.n10 0.189894
R1023 VP.n25 VP.n24 0.189894
R1024 VP.n26 VP.n25 0.189894
R1025 VP.n26 VP.n8 0.189894
R1026 VP.n30 VP.n8 0.189894
R1027 VP.n32 VP.n31 0.189894
R1028 VP.n32 VP.n6 0.189894
R1029 VP.n36 VP.n6 0.189894
R1030 VP.n37 VP.n36 0.189894
R1031 VP.n38 VP.n37 0.189894
R1032 VP.n38 VP.n4 0.189894
R1033 VP.n43 VP.n4 0.189894
R1034 VP.n44 VP.n43 0.189894
R1035 VP.n45 VP.n44 0.189894
R1036 VP.n45 VP.n2 0.189894
R1037 VP.n50 VP.n2 0.189894
R1038 VP.n51 VP.n50 0.189894
R1039 VP.n52 VP.n51 0.189894
R1040 VP.n52 VP.n0 0.189894
R1041 VP.n56 VP.n0 0.189894
R1042 VP VP.n56 0.0516364
R1043 VDD1 VDD1.n0 76.1878
R1044 VDD1.n3 VDD1.n2 76.0732
R1045 VDD1.n3 VDD1.n1 76.0732
R1046 VDD1.n5 VDD1.n4 75.1759
R1047 VDD1.n5 VDD1.n3 43.7423
R1048 VDD1.n4 VDD1.t4 2.57822
R1049 VDD1.n4 VDD1.t2 2.57822
R1050 VDD1.n0 VDD1.t0 2.57822
R1051 VDD1.n0 VDD1.t7 2.57822
R1052 VDD1.n2 VDD1.t5 2.57822
R1053 VDD1.n2 VDD1.t6 2.57822
R1054 VDD1.n1 VDD1.t1 2.57822
R1055 VDD1.n1 VDD1.t3 2.57822
R1056 VDD1 VDD1.n5 0.894897
R1057 B.n391 B.n116 585
R1058 B.n390 B.n389 585
R1059 B.n388 B.n117 585
R1060 B.n387 B.n386 585
R1061 B.n385 B.n118 585
R1062 B.n384 B.n383 585
R1063 B.n382 B.n119 585
R1064 B.n381 B.n380 585
R1065 B.n379 B.n120 585
R1066 B.n378 B.n377 585
R1067 B.n376 B.n121 585
R1068 B.n375 B.n374 585
R1069 B.n373 B.n122 585
R1070 B.n372 B.n371 585
R1071 B.n370 B.n123 585
R1072 B.n369 B.n368 585
R1073 B.n367 B.n124 585
R1074 B.n366 B.n365 585
R1075 B.n364 B.n125 585
R1076 B.n363 B.n362 585
R1077 B.n361 B.n126 585
R1078 B.n360 B.n359 585
R1079 B.n358 B.n127 585
R1080 B.n357 B.n356 585
R1081 B.n355 B.n128 585
R1082 B.n354 B.n353 585
R1083 B.n352 B.n129 585
R1084 B.n351 B.n350 585
R1085 B.n349 B.n130 585
R1086 B.n348 B.n347 585
R1087 B.n346 B.n131 585
R1088 B.n345 B.n344 585
R1089 B.n343 B.n132 585
R1090 B.n342 B.n341 585
R1091 B.n340 B.n133 585
R1092 B.n339 B.n338 585
R1093 B.n337 B.n134 585
R1094 B.n336 B.n335 585
R1095 B.n334 B.n135 585
R1096 B.n333 B.n332 585
R1097 B.n331 B.n136 585
R1098 B.n330 B.n329 585
R1099 B.n328 B.n137 585
R1100 B.n327 B.n326 585
R1101 B.n322 B.n138 585
R1102 B.n321 B.n320 585
R1103 B.n319 B.n139 585
R1104 B.n318 B.n317 585
R1105 B.n316 B.n140 585
R1106 B.n315 B.n314 585
R1107 B.n313 B.n141 585
R1108 B.n312 B.n311 585
R1109 B.n310 B.n142 585
R1110 B.n308 B.n307 585
R1111 B.n306 B.n145 585
R1112 B.n305 B.n304 585
R1113 B.n303 B.n146 585
R1114 B.n302 B.n301 585
R1115 B.n300 B.n147 585
R1116 B.n299 B.n298 585
R1117 B.n297 B.n148 585
R1118 B.n296 B.n295 585
R1119 B.n294 B.n149 585
R1120 B.n293 B.n292 585
R1121 B.n291 B.n150 585
R1122 B.n290 B.n289 585
R1123 B.n288 B.n151 585
R1124 B.n287 B.n286 585
R1125 B.n285 B.n152 585
R1126 B.n284 B.n283 585
R1127 B.n282 B.n153 585
R1128 B.n281 B.n280 585
R1129 B.n279 B.n154 585
R1130 B.n278 B.n277 585
R1131 B.n276 B.n155 585
R1132 B.n275 B.n274 585
R1133 B.n273 B.n156 585
R1134 B.n272 B.n271 585
R1135 B.n270 B.n157 585
R1136 B.n269 B.n268 585
R1137 B.n267 B.n158 585
R1138 B.n266 B.n265 585
R1139 B.n264 B.n159 585
R1140 B.n263 B.n262 585
R1141 B.n261 B.n160 585
R1142 B.n260 B.n259 585
R1143 B.n258 B.n161 585
R1144 B.n257 B.n256 585
R1145 B.n255 B.n162 585
R1146 B.n254 B.n253 585
R1147 B.n252 B.n163 585
R1148 B.n251 B.n250 585
R1149 B.n249 B.n164 585
R1150 B.n248 B.n247 585
R1151 B.n246 B.n165 585
R1152 B.n245 B.n244 585
R1153 B.n393 B.n392 585
R1154 B.n394 B.n115 585
R1155 B.n396 B.n395 585
R1156 B.n397 B.n114 585
R1157 B.n399 B.n398 585
R1158 B.n400 B.n113 585
R1159 B.n402 B.n401 585
R1160 B.n403 B.n112 585
R1161 B.n405 B.n404 585
R1162 B.n406 B.n111 585
R1163 B.n408 B.n407 585
R1164 B.n409 B.n110 585
R1165 B.n411 B.n410 585
R1166 B.n412 B.n109 585
R1167 B.n414 B.n413 585
R1168 B.n415 B.n108 585
R1169 B.n417 B.n416 585
R1170 B.n418 B.n107 585
R1171 B.n420 B.n419 585
R1172 B.n421 B.n106 585
R1173 B.n423 B.n422 585
R1174 B.n424 B.n105 585
R1175 B.n426 B.n425 585
R1176 B.n427 B.n104 585
R1177 B.n429 B.n428 585
R1178 B.n430 B.n103 585
R1179 B.n432 B.n431 585
R1180 B.n433 B.n102 585
R1181 B.n435 B.n434 585
R1182 B.n436 B.n101 585
R1183 B.n438 B.n437 585
R1184 B.n439 B.n100 585
R1185 B.n441 B.n440 585
R1186 B.n442 B.n99 585
R1187 B.n444 B.n443 585
R1188 B.n445 B.n98 585
R1189 B.n447 B.n446 585
R1190 B.n448 B.n97 585
R1191 B.n450 B.n449 585
R1192 B.n451 B.n96 585
R1193 B.n453 B.n452 585
R1194 B.n454 B.n95 585
R1195 B.n456 B.n455 585
R1196 B.n457 B.n94 585
R1197 B.n459 B.n458 585
R1198 B.n460 B.n93 585
R1199 B.n462 B.n461 585
R1200 B.n463 B.n92 585
R1201 B.n465 B.n464 585
R1202 B.n466 B.n91 585
R1203 B.n468 B.n467 585
R1204 B.n469 B.n90 585
R1205 B.n471 B.n470 585
R1206 B.n472 B.n89 585
R1207 B.n474 B.n473 585
R1208 B.n475 B.n88 585
R1209 B.n477 B.n476 585
R1210 B.n478 B.n87 585
R1211 B.n480 B.n479 585
R1212 B.n481 B.n86 585
R1213 B.n483 B.n482 585
R1214 B.n484 B.n85 585
R1215 B.n486 B.n485 585
R1216 B.n487 B.n84 585
R1217 B.n489 B.n488 585
R1218 B.n490 B.n83 585
R1219 B.n492 B.n491 585
R1220 B.n493 B.n82 585
R1221 B.n495 B.n494 585
R1222 B.n496 B.n81 585
R1223 B.n498 B.n497 585
R1224 B.n499 B.n80 585
R1225 B.n501 B.n500 585
R1226 B.n502 B.n79 585
R1227 B.n504 B.n503 585
R1228 B.n505 B.n78 585
R1229 B.n507 B.n506 585
R1230 B.n508 B.n77 585
R1231 B.n510 B.n509 585
R1232 B.n511 B.n76 585
R1233 B.n513 B.n512 585
R1234 B.n514 B.n75 585
R1235 B.n659 B.n22 585
R1236 B.n658 B.n657 585
R1237 B.n656 B.n23 585
R1238 B.n655 B.n654 585
R1239 B.n653 B.n24 585
R1240 B.n652 B.n651 585
R1241 B.n650 B.n25 585
R1242 B.n649 B.n648 585
R1243 B.n647 B.n26 585
R1244 B.n646 B.n645 585
R1245 B.n644 B.n27 585
R1246 B.n643 B.n642 585
R1247 B.n641 B.n28 585
R1248 B.n640 B.n639 585
R1249 B.n638 B.n29 585
R1250 B.n637 B.n636 585
R1251 B.n635 B.n30 585
R1252 B.n634 B.n633 585
R1253 B.n632 B.n31 585
R1254 B.n631 B.n630 585
R1255 B.n629 B.n32 585
R1256 B.n628 B.n627 585
R1257 B.n626 B.n33 585
R1258 B.n625 B.n624 585
R1259 B.n623 B.n34 585
R1260 B.n622 B.n621 585
R1261 B.n620 B.n35 585
R1262 B.n619 B.n618 585
R1263 B.n617 B.n36 585
R1264 B.n616 B.n615 585
R1265 B.n614 B.n37 585
R1266 B.n613 B.n612 585
R1267 B.n611 B.n38 585
R1268 B.n610 B.n609 585
R1269 B.n608 B.n39 585
R1270 B.n607 B.n606 585
R1271 B.n605 B.n40 585
R1272 B.n604 B.n603 585
R1273 B.n602 B.n41 585
R1274 B.n601 B.n600 585
R1275 B.n599 B.n42 585
R1276 B.n598 B.n597 585
R1277 B.n596 B.n43 585
R1278 B.n594 B.n593 585
R1279 B.n592 B.n46 585
R1280 B.n591 B.n590 585
R1281 B.n589 B.n47 585
R1282 B.n588 B.n587 585
R1283 B.n586 B.n48 585
R1284 B.n585 B.n584 585
R1285 B.n583 B.n49 585
R1286 B.n582 B.n581 585
R1287 B.n580 B.n50 585
R1288 B.n579 B.n578 585
R1289 B.n577 B.n51 585
R1290 B.n576 B.n575 585
R1291 B.n574 B.n55 585
R1292 B.n573 B.n572 585
R1293 B.n571 B.n56 585
R1294 B.n570 B.n569 585
R1295 B.n568 B.n57 585
R1296 B.n567 B.n566 585
R1297 B.n565 B.n58 585
R1298 B.n564 B.n563 585
R1299 B.n562 B.n59 585
R1300 B.n561 B.n560 585
R1301 B.n559 B.n60 585
R1302 B.n558 B.n557 585
R1303 B.n556 B.n61 585
R1304 B.n555 B.n554 585
R1305 B.n553 B.n62 585
R1306 B.n552 B.n551 585
R1307 B.n550 B.n63 585
R1308 B.n549 B.n548 585
R1309 B.n547 B.n64 585
R1310 B.n546 B.n545 585
R1311 B.n544 B.n65 585
R1312 B.n543 B.n542 585
R1313 B.n541 B.n66 585
R1314 B.n540 B.n539 585
R1315 B.n538 B.n67 585
R1316 B.n537 B.n536 585
R1317 B.n535 B.n68 585
R1318 B.n534 B.n533 585
R1319 B.n532 B.n69 585
R1320 B.n531 B.n530 585
R1321 B.n529 B.n70 585
R1322 B.n528 B.n527 585
R1323 B.n526 B.n71 585
R1324 B.n525 B.n524 585
R1325 B.n523 B.n72 585
R1326 B.n522 B.n521 585
R1327 B.n520 B.n73 585
R1328 B.n519 B.n518 585
R1329 B.n517 B.n74 585
R1330 B.n516 B.n515 585
R1331 B.n661 B.n660 585
R1332 B.n662 B.n21 585
R1333 B.n664 B.n663 585
R1334 B.n665 B.n20 585
R1335 B.n667 B.n666 585
R1336 B.n668 B.n19 585
R1337 B.n670 B.n669 585
R1338 B.n671 B.n18 585
R1339 B.n673 B.n672 585
R1340 B.n674 B.n17 585
R1341 B.n676 B.n675 585
R1342 B.n677 B.n16 585
R1343 B.n679 B.n678 585
R1344 B.n680 B.n15 585
R1345 B.n682 B.n681 585
R1346 B.n683 B.n14 585
R1347 B.n685 B.n684 585
R1348 B.n686 B.n13 585
R1349 B.n688 B.n687 585
R1350 B.n689 B.n12 585
R1351 B.n691 B.n690 585
R1352 B.n692 B.n11 585
R1353 B.n694 B.n693 585
R1354 B.n695 B.n10 585
R1355 B.n697 B.n696 585
R1356 B.n698 B.n9 585
R1357 B.n700 B.n699 585
R1358 B.n701 B.n8 585
R1359 B.n703 B.n702 585
R1360 B.n704 B.n7 585
R1361 B.n706 B.n705 585
R1362 B.n707 B.n6 585
R1363 B.n709 B.n708 585
R1364 B.n710 B.n5 585
R1365 B.n712 B.n711 585
R1366 B.n713 B.n4 585
R1367 B.n715 B.n714 585
R1368 B.n716 B.n3 585
R1369 B.n718 B.n717 585
R1370 B.n719 B.n0 585
R1371 B.n2 B.n1 585
R1372 B.n186 B.n185 585
R1373 B.n188 B.n187 585
R1374 B.n189 B.n184 585
R1375 B.n191 B.n190 585
R1376 B.n192 B.n183 585
R1377 B.n194 B.n193 585
R1378 B.n195 B.n182 585
R1379 B.n197 B.n196 585
R1380 B.n198 B.n181 585
R1381 B.n200 B.n199 585
R1382 B.n201 B.n180 585
R1383 B.n203 B.n202 585
R1384 B.n204 B.n179 585
R1385 B.n206 B.n205 585
R1386 B.n207 B.n178 585
R1387 B.n209 B.n208 585
R1388 B.n210 B.n177 585
R1389 B.n212 B.n211 585
R1390 B.n213 B.n176 585
R1391 B.n215 B.n214 585
R1392 B.n216 B.n175 585
R1393 B.n218 B.n217 585
R1394 B.n219 B.n174 585
R1395 B.n221 B.n220 585
R1396 B.n222 B.n173 585
R1397 B.n224 B.n223 585
R1398 B.n225 B.n172 585
R1399 B.n227 B.n226 585
R1400 B.n228 B.n171 585
R1401 B.n230 B.n229 585
R1402 B.n231 B.n170 585
R1403 B.n233 B.n232 585
R1404 B.n234 B.n169 585
R1405 B.n236 B.n235 585
R1406 B.n237 B.n168 585
R1407 B.n239 B.n238 585
R1408 B.n240 B.n167 585
R1409 B.n242 B.n241 585
R1410 B.n243 B.n166 585
R1411 B.n245 B.n166 550.159
R1412 B.n393 B.n116 550.159
R1413 B.n515 B.n514 550.159
R1414 B.n660 B.n659 550.159
R1415 B.n323 B.t7 429.279
R1416 B.n52 B.t5 429.279
R1417 B.n143 B.t10 429.279
R1418 B.n44 B.t2 429.279
R1419 B.n324 B.t8 386.42
R1420 B.n53 B.t4 386.42
R1421 B.n144 B.t11 386.42
R1422 B.n45 B.t1 386.42
R1423 B.n143 B.t9 368.272
R1424 B.n323 B.t6 368.272
R1425 B.n52 B.t3 368.272
R1426 B.n44 B.t0 368.272
R1427 B.n721 B.n720 256.663
R1428 B.n720 B.n719 235.042
R1429 B.n720 B.n2 235.042
R1430 B.n246 B.n245 163.367
R1431 B.n247 B.n246 163.367
R1432 B.n247 B.n164 163.367
R1433 B.n251 B.n164 163.367
R1434 B.n252 B.n251 163.367
R1435 B.n253 B.n252 163.367
R1436 B.n253 B.n162 163.367
R1437 B.n257 B.n162 163.367
R1438 B.n258 B.n257 163.367
R1439 B.n259 B.n258 163.367
R1440 B.n259 B.n160 163.367
R1441 B.n263 B.n160 163.367
R1442 B.n264 B.n263 163.367
R1443 B.n265 B.n264 163.367
R1444 B.n265 B.n158 163.367
R1445 B.n269 B.n158 163.367
R1446 B.n270 B.n269 163.367
R1447 B.n271 B.n270 163.367
R1448 B.n271 B.n156 163.367
R1449 B.n275 B.n156 163.367
R1450 B.n276 B.n275 163.367
R1451 B.n277 B.n276 163.367
R1452 B.n277 B.n154 163.367
R1453 B.n281 B.n154 163.367
R1454 B.n282 B.n281 163.367
R1455 B.n283 B.n282 163.367
R1456 B.n283 B.n152 163.367
R1457 B.n287 B.n152 163.367
R1458 B.n288 B.n287 163.367
R1459 B.n289 B.n288 163.367
R1460 B.n289 B.n150 163.367
R1461 B.n293 B.n150 163.367
R1462 B.n294 B.n293 163.367
R1463 B.n295 B.n294 163.367
R1464 B.n295 B.n148 163.367
R1465 B.n299 B.n148 163.367
R1466 B.n300 B.n299 163.367
R1467 B.n301 B.n300 163.367
R1468 B.n301 B.n146 163.367
R1469 B.n305 B.n146 163.367
R1470 B.n306 B.n305 163.367
R1471 B.n307 B.n306 163.367
R1472 B.n307 B.n142 163.367
R1473 B.n312 B.n142 163.367
R1474 B.n313 B.n312 163.367
R1475 B.n314 B.n313 163.367
R1476 B.n314 B.n140 163.367
R1477 B.n318 B.n140 163.367
R1478 B.n319 B.n318 163.367
R1479 B.n320 B.n319 163.367
R1480 B.n320 B.n138 163.367
R1481 B.n327 B.n138 163.367
R1482 B.n328 B.n327 163.367
R1483 B.n329 B.n328 163.367
R1484 B.n329 B.n136 163.367
R1485 B.n333 B.n136 163.367
R1486 B.n334 B.n333 163.367
R1487 B.n335 B.n334 163.367
R1488 B.n335 B.n134 163.367
R1489 B.n339 B.n134 163.367
R1490 B.n340 B.n339 163.367
R1491 B.n341 B.n340 163.367
R1492 B.n341 B.n132 163.367
R1493 B.n345 B.n132 163.367
R1494 B.n346 B.n345 163.367
R1495 B.n347 B.n346 163.367
R1496 B.n347 B.n130 163.367
R1497 B.n351 B.n130 163.367
R1498 B.n352 B.n351 163.367
R1499 B.n353 B.n352 163.367
R1500 B.n353 B.n128 163.367
R1501 B.n357 B.n128 163.367
R1502 B.n358 B.n357 163.367
R1503 B.n359 B.n358 163.367
R1504 B.n359 B.n126 163.367
R1505 B.n363 B.n126 163.367
R1506 B.n364 B.n363 163.367
R1507 B.n365 B.n364 163.367
R1508 B.n365 B.n124 163.367
R1509 B.n369 B.n124 163.367
R1510 B.n370 B.n369 163.367
R1511 B.n371 B.n370 163.367
R1512 B.n371 B.n122 163.367
R1513 B.n375 B.n122 163.367
R1514 B.n376 B.n375 163.367
R1515 B.n377 B.n376 163.367
R1516 B.n377 B.n120 163.367
R1517 B.n381 B.n120 163.367
R1518 B.n382 B.n381 163.367
R1519 B.n383 B.n382 163.367
R1520 B.n383 B.n118 163.367
R1521 B.n387 B.n118 163.367
R1522 B.n388 B.n387 163.367
R1523 B.n389 B.n388 163.367
R1524 B.n389 B.n116 163.367
R1525 B.n514 B.n513 163.367
R1526 B.n513 B.n76 163.367
R1527 B.n509 B.n76 163.367
R1528 B.n509 B.n508 163.367
R1529 B.n508 B.n507 163.367
R1530 B.n507 B.n78 163.367
R1531 B.n503 B.n78 163.367
R1532 B.n503 B.n502 163.367
R1533 B.n502 B.n501 163.367
R1534 B.n501 B.n80 163.367
R1535 B.n497 B.n80 163.367
R1536 B.n497 B.n496 163.367
R1537 B.n496 B.n495 163.367
R1538 B.n495 B.n82 163.367
R1539 B.n491 B.n82 163.367
R1540 B.n491 B.n490 163.367
R1541 B.n490 B.n489 163.367
R1542 B.n489 B.n84 163.367
R1543 B.n485 B.n84 163.367
R1544 B.n485 B.n484 163.367
R1545 B.n484 B.n483 163.367
R1546 B.n483 B.n86 163.367
R1547 B.n479 B.n86 163.367
R1548 B.n479 B.n478 163.367
R1549 B.n478 B.n477 163.367
R1550 B.n477 B.n88 163.367
R1551 B.n473 B.n88 163.367
R1552 B.n473 B.n472 163.367
R1553 B.n472 B.n471 163.367
R1554 B.n471 B.n90 163.367
R1555 B.n467 B.n90 163.367
R1556 B.n467 B.n466 163.367
R1557 B.n466 B.n465 163.367
R1558 B.n465 B.n92 163.367
R1559 B.n461 B.n92 163.367
R1560 B.n461 B.n460 163.367
R1561 B.n460 B.n459 163.367
R1562 B.n459 B.n94 163.367
R1563 B.n455 B.n94 163.367
R1564 B.n455 B.n454 163.367
R1565 B.n454 B.n453 163.367
R1566 B.n453 B.n96 163.367
R1567 B.n449 B.n96 163.367
R1568 B.n449 B.n448 163.367
R1569 B.n448 B.n447 163.367
R1570 B.n447 B.n98 163.367
R1571 B.n443 B.n98 163.367
R1572 B.n443 B.n442 163.367
R1573 B.n442 B.n441 163.367
R1574 B.n441 B.n100 163.367
R1575 B.n437 B.n100 163.367
R1576 B.n437 B.n436 163.367
R1577 B.n436 B.n435 163.367
R1578 B.n435 B.n102 163.367
R1579 B.n431 B.n102 163.367
R1580 B.n431 B.n430 163.367
R1581 B.n430 B.n429 163.367
R1582 B.n429 B.n104 163.367
R1583 B.n425 B.n104 163.367
R1584 B.n425 B.n424 163.367
R1585 B.n424 B.n423 163.367
R1586 B.n423 B.n106 163.367
R1587 B.n419 B.n106 163.367
R1588 B.n419 B.n418 163.367
R1589 B.n418 B.n417 163.367
R1590 B.n417 B.n108 163.367
R1591 B.n413 B.n108 163.367
R1592 B.n413 B.n412 163.367
R1593 B.n412 B.n411 163.367
R1594 B.n411 B.n110 163.367
R1595 B.n407 B.n110 163.367
R1596 B.n407 B.n406 163.367
R1597 B.n406 B.n405 163.367
R1598 B.n405 B.n112 163.367
R1599 B.n401 B.n112 163.367
R1600 B.n401 B.n400 163.367
R1601 B.n400 B.n399 163.367
R1602 B.n399 B.n114 163.367
R1603 B.n395 B.n114 163.367
R1604 B.n395 B.n394 163.367
R1605 B.n394 B.n393 163.367
R1606 B.n659 B.n658 163.367
R1607 B.n658 B.n23 163.367
R1608 B.n654 B.n23 163.367
R1609 B.n654 B.n653 163.367
R1610 B.n653 B.n652 163.367
R1611 B.n652 B.n25 163.367
R1612 B.n648 B.n25 163.367
R1613 B.n648 B.n647 163.367
R1614 B.n647 B.n646 163.367
R1615 B.n646 B.n27 163.367
R1616 B.n642 B.n27 163.367
R1617 B.n642 B.n641 163.367
R1618 B.n641 B.n640 163.367
R1619 B.n640 B.n29 163.367
R1620 B.n636 B.n29 163.367
R1621 B.n636 B.n635 163.367
R1622 B.n635 B.n634 163.367
R1623 B.n634 B.n31 163.367
R1624 B.n630 B.n31 163.367
R1625 B.n630 B.n629 163.367
R1626 B.n629 B.n628 163.367
R1627 B.n628 B.n33 163.367
R1628 B.n624 B.n33 163.367
R1629 B.n624 B.n623 163.367
R1630 B.n623 B.n622 163.367
R1631 B.n622 B.n35 163.367
R1632 B.n618 B.n35 163.367
R1633 B.n618 B.n617 163.367
R1634 B.n617 B.n616 163.367
R1635 B.n616 B.n37 163.367
R1636 B.n612 B.n37 163.367
R1637 B.n612 B.n611 163.367
R1638 B.n611 B.n610 163.367
R1639 B.n610 B.n39 163.367
R1640 B.n606 B.n39 163.367
R1641 B.n606 B.n605 163.367
R1642 B.n605 B.n604 163.367
R1643 B.n604 B.n41 163.367
R1644 B.n600 B.n41 163.367
R1645 B.n600 B.n599 163.367
R1646 B.n599 B.n598 163.367
R1647 B.n598 B.n43 163.367
R1648 B.n593 B.n43 163.367
R1649 B.n593 B.n592 163.367
R1650 B.n592 B.n591 163.367
R1651 B.n591 B.n47 163.367
R1652 B.n587 B.n47 163.367
R1653 B.n587 B.n586 163.367
R1654 B.n586 B.n585 163.367
R1655 B.n585 B.n49 163.367
R1656 B.n581 B.n49 163.367
R1657 B.n581 B.n580 163.367
R1658 B.n580 B.n579 163.367
R1659 B.n579 B.n51 163.367
R1660 B.n575 B.n51 163.367
R1661 B.n575 B.n574 163.367
R1662 B.n574 B.n573 163.367
R1663 B.n573 B.n56 163.367
R1664 B.n569 B.n56 163.367
R1665 B.n569 B.n568 163.367
R1666 B.n568 B.n567 163.367
R1667 B.n567 B.n58 163.367
R1668 B.n563 B.n58 163.367
R1669 B.n563 B.n562 163.367
R1670 B.n562 B.n561 163.367
R1671 B.n561 B.n60 163.367
R1672 B.n557 B.n60 163.367
R1673 B.n557 B.n556 163.367
R1674 B.n556 B.n555 163.367
R1675 B.n555 B.n62 163.367
R1676 B.n551 B.n62 163.367
R1677 B.n551 B.n550 163.367
R1678 B.n550 B.n549 163.367
R1679 B.n549 B.n64 163.367
R1680 B.n545 B.n64 163.367
R1681 B.n545 B.n544 163.367
R1682 B.n544 B.n543 163.367
R1683 B.n543 B.n66 163.367
R1684 B.n539 B.n66 163.367
R1685 B.n539 B.n538 163.367
R1686 B.n538 B.n537 163.367
R1687 B.n537 B.n68 163.367
R1688 B.n533 B.n68 163.367
R1689 B.n533 B.n532 163.367
R1690 B.n532 B.n531 163.367
R1691 B.n531 B.n70 163.367
R1692 B.n527 B.n70 163.367
R1693 B.n527 B.n526 163.367
R1694 B.n526 B.n525 163.367
R1695 B.n525 B.n72 163.367
R1696 B.n521 B.n72 163.367
R1697 B.n521 B.n520 163.367
R1698 B.n520 B.n519 163.367
R1699 B.n519 B.n74 163.367
R1700 B.n515 B.n74 163.367
R1701 B.n660 B.n21 163.367
R1702 B.n664 B.n21 163.367
R1703 B.n665 B.n664 163.367
R1704 B.n666 B.n665 163.367
R1705 B.n666 B.n19 163.367
R1706 B.n670 B.n19 163.367
R1707 B.n671 B.n670 163.367
R1708 B.n672 B.n671 163.367
R1709 B.n672 B.n17 163.367
R1710 B.n676 B.n17 163.367
R1711 B.n677 B.n676 163.367
R1712 B.n678 B.n677 163.367
R1713 B.n678 B.n15 163.367
R1714 B.n682 B.n15 163.367
R1715 B.n683 B.n682 163.367
R1716 B.n684 B.n683 163.367
R1717 B.n684 B.n13 163.367
R1718 B.n688 B.n13 163.367
R1719 B.n689 B.n688 163.367
R1720 B.n690 B.n689 163.367
R1721 B.n690 B.n11 163.367
R1722 B.n694 B.n11 163.367
R1723 B.n695 B.n694 163.367
R1724 B.n696 B.n695 163.367
R1725 B.n696 B.n9 163.367
R1726 B.n700 B.n9 163.367
R1727 B.n701 B.n700 163.367
R1728 B.n702 B.n701 163.367
R1729 B.n702 B.n7 163.367
R1730 B.n706 B.n7 163.367
R1731 B.n707 B.n706 163.367
R1732 B.n708 B.n707 163.367
R1733 B.n708 B.n5 163.367
R1734 B.n712 B.n5 163.367
R1735 B.n713 B.n712 163.367
R1736 B.n714 B.n713 163.367
R1737 B.n714 B.n3 163.367
R1738 B.n718 B.n3 163.367
R1739 B.n719 B.n718 163.367
R1740 B.n186 B.n2 163.367
R1741 B.n187 B.n186 163.367
R1742 B.n187 B.n184 163.367
R1743 B.n191 B.n184 163.367
R1744 B.n192 B.n191 163.367
R1745 B.n193 B.n192 163.367
R1746 B.n193 B.n182 163.367
R1747 B.n197 B.n182 163.367
R1748 B.n198 B.n197 163.367
R1749 B.n199 B.n198 163.367
R1750 B.n199 B.n180 163.367
R1751 B.n203 B.n180 163.367
R1752 B.n204 B.n203 163.367
R1753 B.n205 B.n204 163.367
R1754 B.n205 B.n178 163.367
R1755 B.n209 B.n178 163.367
R1756 B.n210 B.n209 163.367
R1757 B.n211 B.n210 163.367
R1758 B.n211 B.n176 163.367
R1759 B.n215 B.n176 163.367
R1760 B.n216 B.n215 163.367
R1761 B.n217 B.n216 163.367
R1762 B.n217 B.n174 163.367
R1763 B.n221 B.n174 163.367
R1764 B.n222 B.n221 163.367
R1765 B.n223 B.n222 163.367
R1766 B.n223 B.n172 163.367
R1767 B.n227 B.n172 163.367
R1768 B.n228 B.n227 163.367
R1769 B.n229 B.n228 163.367
R1770 B.n229 B.n170 163.367
R1771 B.n233 B.n170 163.367
R1772 B.n234 B.n233 163.367
R1773 B.n235 B.n234 163.367
R1774 B.n235 B.n168 163.367
R1775 B.n239 B.n168 163.367
R1776 B.n240 B.n239 163.367
R1777 B.n241 B.n240 163.367
R1778 B.n241 B.n166 163.367
R1779 B.n309 B.n144 59.5399
R1780 B.n325 B.n324 59.5399
R1781 B.n54 B.n53 59.5399
R1782 B.n595 B.n45 59.5399
R1783 B.n144 B.n143 42.8611
R1784 B.n324 B.n323 42.8611
R1785 B.n53 B.n52 42.8611
R1786 B.n45 B.n44 42.8611
R1787 B.n661 B.n22 35.7468
R1788 B.n516 B.n75 35.7468
R1789 B.n244 B.n243 35.7468
R1790 B.n392 B.n391 35.7468
R1791 B B.n721 18.0485
R1792 B.n662 B.n661 10.6151
R1793 B.n663 B.n662 10.6151
R1794 B.n663 B.n20 10.6151
R1795 B.n667 B.n20 10.6151
R1796 B.n668 B.n667 10.6151
R1797 B.n669 B.n668 10.6151
R1798 B.n669 B.n18 10.6151
R1799 B.n673 B.n18 10.6151
R1800 B.n674 B.n673 10.6151
R1801 B.n675 B.n674 10.6151
R1802 B.n675 B.n16 10.6151
R1803 B.n679 B.n16 10.6151
R1804 B.n680 B.n679 10.6151
R1805 B.n681 B.n680 10.6151
R1806 B.n681 B.n14 10.6151
R1807 B.n685 B.n14 10.6151
R1808 B.n686 B.n685 10.6151
R1809 B.n687 B.n686 10.6151
R1810 B.n687 B.n12 10.6151
R1811 B.n691 B.n12 10.6151
R1812 B.n692 B.n691 10.6151
R1813 B.n693 B.n692 10.6151
R1814 B.n693 B.n10 10.6151
R1815 B.n697 B.n10 10.6151
R1816 B.n698 B.n697 10.6151
R1817 B.n699 B.n698 10.6151
R1818 B.n699 B.n8 10.6151
R1819 B.n703 B.n8 10.6151
R1820 B.n704 B.n703 10.6151
R1821 B.n705 B.n704 10.6151
R1822 B.n705 B.n6 10.6151
R1823 B.n709 B.n6 10.6151
R1824 B.n710 B.n709 10.6151
R1825 B.n711 B.n710 10.6151
R1826 B.n711 B.n4 10.6151
R1827 B.n715 B.n4 10.6151
R1828 B.n716 B.n715 10.6151
R1829 B.n717 B.n716 10.6151
R1830 B.n717 B.n0 10.6151
R1831 B.n657 B.n22 10.6151
R1832 B.n657 B.n656 10.6151
R1833 B.n656 B.n655 10.6151
R1834 B.n655 B.n24 10.6151
R1835 B.n651 B.n24 10.6151
R1836 B.n651 B.n650 10.6151
R1837 B.n650 B.n649 10.6151
R1838 B.n649 B.n26 10.6151
R1839 B.n645 B.n26 10.6151
R1840 B.n645 B.n644 10.6151
R1841 B.n644 B.n643 10.6151
R1842 B.n643 B.n28 10.6151
R1843 B.n639 B.n28 10.6151
R1844 B.n639 B.n638 10.6151
R1845 B.n638 B.n637 10.6151
R1846 B.n637 B.n30 10.6151
R1847 B.n633 B.n30 10.6151
R1848 B.n633 B.n632 10.6151
R1849 B.n632 B.n631 10.6151
R1850 B.n631 B.n32 10.6151
R1851 B.n627 B.n32 10.6151
R1852 B.n627 B.n626 10.6151
R1853 B.n626 B.n625 10.6151
R1854 B.n625 B.n34 10.6151
R1855 B.n621 B.n34 10.6151
R1856 B.n621 B.n620 10.6151
R1857 B.n620 B.n619 10.6151
R1858 B.n619 B.n36 10.6151
R1859 B.n615 B.n36 10.6151
R1860 B.n615 B.n614 10.6151
R1861 B.n614 B.n613 10.6151
R1862 B.n613 B.n38 10.6151
R1863 B.n609 B.n38 10.6151
R1864 B.n609 B.n608 10.6151
R1865 B.n608 B.n607 10.6151
R1866 B.n607 B.n40 10.6151
R1867 B.n603 B.n40 10.6151
R1868 B.n603 B.n602 10.6151
R1869 B.n602 B.n601 10.6151
R1870 B.n601 B.n42 10.6151
R1871 B.n597 B.n42 10.6151
R1872 B.n597 B.n596 10.6151
R1873 B.n594 B.n46 10.6151
R1874 B.n590 B.n46 10.6151
R1875 B.n590 B.n589 10.6151
R1876 B.n589 B.n588 10.6151
R1877 B.n588 B.n48 10.6151
R1878 B.n584 B.n48 10.6151
R1879 B.n584 B.n583 10.6151
R1880 B.n583 B.n582 10.6151
R1881 B.n582 B.n50 10.6151
R1882 B.n578 B.n577 10.6151
R1883 B.n577 B.n576 10.6151
R1884 B.n576 B.n55 10.6151
R1885 B.n572 B.n55 10.6151
R1886 B.n572 B.n571 10.6151
R1887 B.n571 B.n570 10.6151
R1888 B.n570 B.n57 10.6151
R1889 B.n566 B.n57 10.6151
R1890 B.n566 B.n565 10.6151
R1891 B.n565 B.n564 10.6151
R1892 B.n564 B.n59 10.6151
R1893 B.n560 B.n59 10.6151
R1894 B.n560 B.n559 10.6151
R1895 B.n559 B.n558 10.6151
R1896 B.n558 B.n61 10.6151
R1897 B.n554 B.n61 10.6151
R1898 B.n554 B.n553 10.6151
R1899 B.n553 B.n552 10.6151
R1900 B.n552 B.n63 10.6151
R1901 B.n548 B.n63 10.6151
R1902 B.n548 B.n547 10.6151
R1903 B.n547 B.n546 10.6151
R1904 B.n546 B.n65 10.6151
R1905 B.n542 B.n65 10.6151
R1906 B.n542 B.n541 10.6151
R1907 B.n541 B.n540 10.6151
R1908 B.n540 B.n67 10.6151
R1909 B.n536 B.n67 10.6151
R1910 B.n536 B.n535 10.6151
R1911 B.n535 B.n534 10.6151
R1912 B.n534 B.n69 10.6151
R1913 B.n530 B.n69 10.6151
R1914 B.n530 B.n529 10.6151
R1915 B.n529 B.n528 10.6151
R1916 B.n528 B.n71 10.6151
R1917 B.n524 B.n71 10.6151
R1918 B.n524 B.n523 10.6151
R1919 B.n523 B.n522 10.6151
R1920 B.n522 B.n73 10.6151
R1921 B.n518 B.n73 10.6151
R1922 B.n518 B.n517 10.6151
R1923 B.n517 B.n516 10.6151
R1924 B.n512 B.n75 10.6151
R1925 B.n512 B.n511 10.6151
R1926 B.n511 B.n510 10.6151
R1927 B.n510 B.n77 10.6151
R1928 B.n506 B.n77 10.6151
R1929 B.n506 B.n505 10.6151
R1930 B.n505 B.n504 10.6151
R1931 B.n504 B.n79 10.6151
R1932 B.n500 B.n79 10.6151
R1933 B.n500 B.n499 10.6151
R1934 B.n499 B.n498 10.6151
R1935 B.n498 B.n81 10.6151
R1936 B.n494 B.n81 10.6151
R1937 B.n494 B.n493 10.6151
R1938 B.n493 B.n492 10.6151
R1939 B.n492 B.n83 10.6151
R1940 B.n488 B.n83 10.6151
R1941 B.n488 B.n487 10.6151
R1942 B.n487 B.n486 10.6151
R1943 B.n486 B.n85 10.6151
R1944 B.n482 B.n85 10.6151
R1945 B.n482 B.n481 10.6151
R1946 B.n481 B.n480 10.6151
R1947 B.n480 B.n87 10.6151
R1948 B.n476 B.n87 10.6151
R1949 B.n476 B.n475 10.6151
R1950 B.n475 B.n474 10.6151
R1951 B.n474 B.n89 10.6151
R1952 B.n470 B.n89 10.6151
R1953 B.n470 B.n469 10.6151
R1954 B.n469 B.n468 10.6151
R1955 B.n468 B.n91 10.6151
R1956 B.n464 B.n91 10.6151
R1957 B.n464 B.n463 10.6151
R1958 B.n463 B.n462 10.6151
R1959 B.n462 B.n93 10.6151
R1960 B.n458 B.n93 10.6151
R1961 B.n458 B.n457 10.6151
R1962 B.n457 B.n456 10.6151
R1963 B.n456 B.n95 10.6151
R1964 B.n452 B.n95 10.6151
R1965 B.n452 B.n451 10.6151
R1966 B.n451 B.n450 10.6151
R1967 B.n450 B.n97 10.6151
R1968 B.n446 B.n97 10.6151
R1969 B.n446 B.n445 10.6151
R1970 B.n445 B.n444 10.6151
R1971 B.n444 B.n99 10.6151
R1972 B.n440 B.n99 10.6151
R1973 B.n440 B.n439 10.6151
R1974 B.n439 B.n438 10.6151
R1975 B.n438 B.n101 10.6151
R1976 B.n434 B.n101 10.6151
R1977 B.n434 B.n433 10.6151
R1978 B.n433 B.n432 10.6151
R1979 B.n432 B.n103 10.6151
R1980 B.n428 B.n103 10.6151
R1981 B.n428 B.n427 10.6151
R1982 B.n427 B.n426 10.6151
R1983 B.n426 B.n105 10.6151
R1984 B.n422 B.n105 10.6151
R1985 B.n422 B.n421 10.6151
R1986 B.n421 B.n420 10.6151
R1987 B.n420 B.n107 10.6151
R1988 B.n416 B.n107 10.6151
R1989 B.n416 B.n415 10.6151
R1990 B.n415 B.n414 10.6151
R1991 B.n414 B.n109 10.6151
R1992 B.n410 B.n109 10.6151
R1993 B.n410 B.n409 10.6151
R1994 B.n409 B.n408 10.6151
R1995 B.n408 B.n111 10.6151
R1996 B.n404 B.n111 10.6151
R1997 B.n404 B.n403 10.6151
R1998 B.n403 B.n402 10.6151
R1999 B.n402 B.n113 10.6151
R2000 B.n398 B.n113 10.6151
R2001 B.n398 B.n397 10.6151
R2002 B.n397 B.n396 10.6151
R2003 B.n396 B.n115 10.6151
R2004 B.n392 B.n115 10.6151
R2005 B.n185 B.n1 10.6151
R2006 B.n188 B.n185 10.6151
R2007 B.n189 B.n188 10.6151
R2008 B.n190 B.n189 10.6151
R2009 B.n190 B.n183 10.6151
R2010 B.n194 B.n183 10.6151
R2011 B.n195 B.n194 10.6151
R2012 B.n196 B.n195 10.6151
R2013 B.n196 B.n181 10.6151
R2014 B.n200 B.n181 10.6151
R2015 B.n201 B.n200 10.6151
R2016 B.n202 B.n201 10.6151
R2017 B.n202 B.n179 10.6151
R2018 B.n206 B.n179 10.6151
R2019 B.n207 B.n206 10.6151
R2020 B.n208 B.n207 10.6151
R2021 B.n208 B.n177 10.6151
R2022 B.n212 B.n177 10.6151
R2023 B.n213 B.n212 10.6151
R2024 B.n214 B.n213 10.6151
R2025 B.n214 B.n175 10.6151
R2026 B.n218 B.n175 10.6151
R2027 B.n219 B.n218 10.6151
R2028 B.n220 B.n219 10.6151
R2029 B.n220 B.n173 10.6151
R2030 B.n224 B.n173 10.6151
R2031 B.n225 B.n224 10.6151
R2032 B.n226 B.n225 10.6151
R2033 B.n226 B.n171 10.6151
R2034 B.n230 B.n171 10.6151
R2035 B.n231 B.n230 10.6151
R2036 B.n232 B.n231 10.6151
R2037 B.n232 B.n169 10.6151
R2038 B.n236 B.n169 10.6151
R2039 B.n237 B.n236 10.6151
R2040 B.n238 B.n237 10.6151
R2041 B.n238 B.n167 10.6151
R2042 B.n242 B.n167 10.6151
R2043 B.n243 B.n242 10.6151
R2044 B.n244 B.n165 10.6151
R2045 B.n248 B.n165 10.6151
R2046 B.n249 B.n248 10.6151
R2047 B.n250 B.n249 10.6151
R2048 B.n250 B.n163 10.6151
R2049 B.n254 B.n163 10.6151
R2050 B.n255 B.n254 10.6151
R2051 B.n256 B.n255 10.6151
R2052 B.n256 B.n161 10.6151
R2053 B.n260 B.n161 10.6151
R2054 B.n261 B.n260 10.6151
R2055 B.n262 B.n261 10.6151
R2056 B.n262 B.n159 10.6151
R2057 B.n266 B.n159 10.6151
R2058 B.n267 B.n266 10.6151
R2059 B.n268 B.n267 10.6151
R2060 B.n268 B.n157 10.6151
R2061 B.n272 B.n157 10.6151
R2062 B.n273 B.n272 10.6151
R2063 B.n274 B.n273 10.6151
R2064 B.n274 B.n155 10.6151
R2065 B.n278 B.n155 10.6151
R2066 B.n279 B.n278 10.6151
R2067 B.n280 B.n279 10.6151
R2068 B.n280 B.n153 10.6151
R2069 B.n284 B.n153 10.6151
R2070 B.n285 B.n284 10.6151
R2071 B.n286 B.n285 10.6151
R2072 B.n286 B.n151 10.6151
R2073 B.n290 B.n151 10.6151
R2074 B.n291 B.n290 10.6151
R2075 B.n292 B.n291 10.6151
R2076 B.n292 B.n149 10.6151
R2077 B.n296 B.n149 10.6151
R2078 B.n297 B.n296 10.6151
R2079 B.n298 B.n297 10.6151
R2080 B.n298 B.n147 10.6151
R2081 B.n302 B.n147 10.6151
R2082 B.n303 B.n302 10.6151
R2083 B.n304 B.n303 10.6151
R2084 B.n304 B.n145 10.6151
R2085 B.n308 B.n145 10.6151
R2086 B.n311 B.n310 10.6151
R2087 B.n311 B.n141 10.6151
R2088 B.n315 B.n141 10.6151
R2089 B.n316 B.n315 10.6151
R2090 B.n317 B.n316 10.6151
R2091 B.n317 B.n139 10.6151
R2092 B.n321 B.n139 10.6151
R2093 B.n322 B.n321 10.6151
R2094 B.n326 B.n322 10.6151
R2095 B.n330 B.n137 10.6151
R2096 B.n331 B.n330 10.6151
R2097 B.n332 B.n331 10.6151
R2098 B.n332 B.n135 10.6151
R2099 B.n336 B.n135 10.6151
R2100 B.n337 B.n336 10.6151
R2101 B.n338 B.n337 10.6151
R2102 B.n338 B.n133 10.6151
R2103 B.n342 B.n133 10.6151
R2104 B.n343 B.n342 10.6151
R2105 B.n344 B.n343 10.6151
R2106 B.n344 B.n131 10.6151
R2107 B.n348 B.n131 10.6151
R2108 B.n349 B.n348 10.6151
R2109 B.n350 B.n349 10.6151
R2110 B.n350 B.n129 10.6151
R2111 B.n354 B.n129 10.6151
R2112 B.n355 B.n354 10.6151
R2113 B.n356 B.n355 10.6151
R2114 B.n356 B.n127 10.6151
R2115 B.n360 B.n127 10.6151
R2116 B.n361 B.n360 10.6151
R2117 B.n362 B.n361 10.6151
R2118 B.n362 B.n125 10.6151
R2119 B.n366 B.n125 10.6151
R2120 B.n367 B.n366 10.6151
R2121 B.n368 B.n367 10.6151
R2122 B.n368 B.n123 10.6151
R2123 B.n372 B.n123 10.6151
R2124 B.n373 B.n372 10.6151
R2125 B.n374 B.n373 10.6151
R2126 B.n374 B.n121 10.6151
R2127 B.n378 B.n121 10.6151
R2128 B.n379 B.n378 10.6151
R2129 B.n380 B.n379 10.6151
R2130 B.n380 B.n119 10.6151
R2131 B.n384 B.n119 10.6151
R2132 B.n385 B.n384 10.6151
R2133 B.n386 B.n385 10.6151
R2134 B.n386 B.n117 10.6151
R2135 B.n390 B.n117 10.6151
R2136 B.n391 B.n390 10.6151
R2137 B.n596 B.n595 9.36635
R2138 B.n578 B.n54 9.36635
R2139 B.n309 B.n308 9.36635
R2140 B.n325 B.n137 9.36635
R2141 B.n721 B.n0 8.11757
R2142 B.n721 B.n1 8.11757
R2143 B.n595 B.n594 1.24928
R2144 B.n54 B.n50 1.24928
R2145 B.n310 B.n309 1.24928
R2146 B.n326 B.n325 1.24928
C0 VN w_n3180_n3490# 6.27946f
C1 VP VTAIL 8.613831f
C2 B w_n3180_n3490# 9.184091f
C3 VDD1 VN 0.150048f
C4 VDD2 VN 8.469f
C5 VDD1 B 1.44708f
C6 VDD2 B 1.52046f
C7 VN VTAIL 8.59973f
C8 VN VP 6.89328f
C9 B VTAIL 4.81408f
C10 VDD1 w_n3180_n3490# 1.73008f
C11 B VP 1.74944f
C12 VDD2 w_n3180_n3490# 1.81458f
C13 VTAIL w_n3180_n3490# 4.31258f
C14 VDD2 VDD1 1.40012f
C15 VP w_n3180_n3490# 6.69017f
C16 B VN 1.06479f
C17 VDD1 VTAIL 8.40004f
C18 VDD1 VP 8.76059f
C19 VDD2 VTAIL 8.44963f
C20 VDD2 VP 0.442677f
C21 VDD2 VSUBS 1.607506f
C22 VDD1 VSUBS 2.129638f
C23 VTAIL VSUBS 1.239678f
C24 VN VSUBS 5.84929f
C25 VP VSUBS 2.855427f
C26 B VSUBS 4.249143f
C27 w_n3180_n3490# VSUBS 0.136498p
C28 B.n0 VSUBS 0.006227f
C29 B.n1 VSUBS 0.006227f
C30 B.n2 VSUBS 0.00921f
C31 B.n3 VSUBS 0.007057f
C32 B.n4 VSUBS 0.007057f
C33 B.n5 VSUBS 0.007057f
C34 B.n6 VSUBS 0.007057f
C35 B.n7 VSUBS 0.007057f
C36 B.n8 VSUBS 0.007057f
C37 B.n9 VSUBS 0.007057f
C38 B.n10 VSUBS 0.007057f
C39 B.n11 VSUBS 0.007057f
C40 B.n12 VSUBS 0.007057f
C41 B.n13 VSUBS 0.007057f
C42 B.n14 VSUBS 0.007057f
C43 B.n15 VSUBS 0.007057f
C44 B.n16 VSUBS 0.007057f
C45 B.n17 VSUBS 0.007057f
C46 B.n18 VSUBS 0.007057f
C47 B.n19 VSUBS 0.007057f
C48 B.n20 VSUBS 0.007057f
C49 B.n21 VSUBS 0.007057f
C50 B.n22 VSUBS 0.017846f
C51 B.n23 VSUBS 0.007057f
C52 B.n24 VSUBS 0.007057f
C53 B.n25 VSUBS 0.007057f
C54 B.n26 VSUBS 0.007057f
C55 B.n27 VSUBS 0.007057f
C56 B.n28 VSUBS 0.007057f
C57 B.n29 VSUBS 0.007057f
C58 B.n30 VSUBS 0.007057f
C59 B.n31 VSUBS 0.007057f
C60 B.n32 VSUBS 0.007057f
C61 B.n33 VSUBS 0.007057f
C62 B.n34 VSUBS 0.007057f
C63 B.n35 VSUBS 0.007057f
C64 B.n36 VSUBS 0.007057f
C65 B.n37 VSUBS 0.007057f
C66 B.n38 VSUBS 0.007057f
C67 B.n39 VSUBS 0.007057f
C68 B.n40 VSUBS 0.007057f
C69 B.n41 VSUBS 0.007057f
C70 B.n42 VSUBS 0.007057f
C71 B.n43 VSUBS 0.007057f
C72 B.t1 VSUBS 0.226299f
C73 B.t2 VSUBS 0.251211f
C74 B.t0 VSUBS 1.0601f
C75 B.n44 VSUBS 0.388681f
C76 B.n45 VSUBS 0.259582f
C77 B.n46 VSUBS 0.007057f
C78 B.n47 VSUBS 0.007057f
C79 B.n48 VSUBS 0.007057f
C80 B.n49 VSUBS 0.007057f
C81 B.n50 VSUBS 0.003944f
C82 B.n51 VSUBS 0.007057f
C83 B.t4 VSUBS 0.226302f
C84 B.t5 VSUBS 0.251214f
C85 B.t3 VSUBS 1.0601f
C86 B.n52 VSUBS 0.388678f
C87 B.n53 VSUBS 0.259579f
C88 B.n54 VSUBS 0.016351f
C89 B.n55 VSUBS 0.007057f
C90 B.n56 VSUBS 0.007057f
C91 B.n57 VSUBS 0.007057f
C92 B.n58 VSUBS 0.007057f
C93 B.n59 VSUBS 0.007057f
C94 B.n60 VSUBS 0.007057f
C95 B.n61 VSUBS 0.007057f
C96 B.n62 VSUBS 0.007057f
C97 B.n63 VSUBS 0.007057f
C98 B.n64 VSUBS 0.007057f
C99 B.n65 VSUBS 0.007057f
C100 B.n66 VSUBS 0.007057f
C101 B.n67 VSUBS 0.007057f
C102 B.n68 VSUBS 0.007057f
C103 B.n69 VSUBS 0.007057f
C104 B.n70 VSUBS 0.007057f
C105 B.n71 VSUBS 0.007057f
C106 B.n72 VSUBS 0.007057f
C107 B.n73 VSUBS 0.007057f
C108 B.n74 VSUBS 0.007057f
C109 B.n75 VSUBS 0.017233f
C110 B.n76 VSUBS 0.007057f
C111 B.n77 VSUBS 0.007057f
C112 B.n78 VSUBS 0.007057f
C113 B.n79 VSUBS 0.007057f
C114 B.n80 VSUBS 0.007057f
C115 B.n81 VSUBS 0.007057f
C116 B.n82 VSUBS 0.007057f
C117 B.n83 VSUBS 0.007057f
C118 B.n84 VSUBS 0.007057f
C119 B.n85 VSUBS 0.007057f
C120 B.n86 VSUBS 0.007057f
C121 B.n87 VSUBS 0.007057f
C122 B.n88 VSUBS 0.007057f
C123 B.n89 VSUBS 0.007057f
C124 B.n90 VSUBS 0.007057f
C125 B.n91 VSUBS 0.007057f
C126 B.n92 VSUBS 0.007057f
C127 B.n93 VSUBS 0.007057f
C128 B.n94 VSUBS 0.007057f
C129 B.n95 VSUBS 0.007057f
C130 B.n96 VSUBS 0.007057f
C131 B.n97 VSUBS 0.007057f
C132 B.n98 VSUBS 0.007057f
C133 B.n99 VSUBS 0.007057f
C134 B.n100 VSUBS 0.007057f
C135 B.n101 VSUBS 0.007057f
C136 B.n102 VSUBS 0.007057f
C137 B.n103 VSUBS 0.007057f
C138 B.n104 VSUBS 0.007057f
C139 B.n105 VSUBS 0.007057f
C140 B.n106 VSUBS 0.007057f
C141 B.n107 VSUBS 0.007057f
C142 B.n108 VSUBS 0.007057f
C143 B.n109 VSUBS 0.007057f
C144 B.n110 VSUBS 0.007057f
C145 B.n111 VSUBS 0.007057f
C146 B.n112 VSUBS 0.007057f
C147 B.n113 VSUBS 0.007057f
C148 B.n114 VSUBS 0.007057f
C149 B.n115 VSUBS 0.007057f
C150 B.n116 VSUBS 0.017846f
C151 B.n117 VSUBS 0.007057f
C152 B.n118 VSUBS 0.007057f
C153 B.n119 VSUBS 0.007057f
C154 B.n120 VSUBS 0.007057f
C155 B.n121 VSUBS 0.007057f
C156 B.n122 VSUBS 0.007057f
C157 B.n123 VSUBS 0.007057f
C158 B.n124 VSUBS 0.007057f
C159 B.n125 VSUBS 0.007057f
C160 B.n126 VSUBS 0.007057f
C161 B.n127 VSUBS 0.007057f
C162 B.n128 VSUBS 0.007057f
C163 B.n129 VSUBS 0.007057f
C164 B.n130 VSUBS 0.007057f
C165 B.n131 VSUBS 0.007057f
C166 B.n132 VSUBS 0.007057f
C167 B.n133 VSUBS 0.007057f
C168 B.n134 VSUBS 0.007057f
C169 B.n135 VSUBS 0.007057f
C170 B.n136 VSUBS 0.007057f
C171 B.n137 VSUBS 0.006642f
C172 B.n138 VSUBS 0.007057f
C173 B.n139 VSUBS 0.007057f
C174 B.n140 VSUBS 0.007057f
C175 B.n141 VSUBS 0.007057f
C176 B.n142 VSUBS 0.007057f
C177 B.t11 VSUBS 0.226299f
C178 B.t10 VSUBS 0.251211f
C179 B.t9 VSUBS 1.0601f
C180 B.n143 VSUBS 0.388681f
C181 B.n144 VSUBS 0.259582f
C182 B.n145 VSUBS 0.007057f
C183 B.n146 VSUBS 0.007057f
C184 B.n147 VSUBS 0.007057f
C185 B.n148 VSUBS 0.007057f
C186 B.n149 VSUBS 0.007057f
C187 B.n150 VSUBS 0.007057f
C188 B.n151 VSUBS 0.007057f
C189 B.n152 VSUBS 0.007057f
C190 B.n153 VSUBS 0.007057f
C191 B.n154 VSUBS 0.007057f
C192 B.n155 VSUBS 0.007057f
C193 B.n156 VSUBS 0.007057f
C194 B.n157 VSUBS 0.007057f
C195 B.n158 VSUBS 0.007057f
C196 B.n159 VSUBS 0.007057f
C197 B.n160 VSUBS 0.007057f
C198 B.n161 VSUBS 0.007057f
C199 B.n162 VSUBS 0.007057f
C200 B.n163 VSUBS 0.007057f
C201 B.n164 VSUBS 0.007057f
C202 B.n165 VSUBS 0.007057f
C203 B.n166 VSUBS 0.017233f
C204 B.n167 VSUBS 0.007057f
C205 B.n168 VSUBS 0.007057f
C206 B.n169 VSUBS 0.007057f
C207 B.n170 VSUBS 0.007057f
C208 B.n171 VSUBS 0.007057f
C209 B.n172 VSUBS 0.007057f
C210 B.n173 VSUBS 0.007057f
C211 B.n174 VSUBS 0.007057f
C212 B.n175 VSUBS 0.007057f
C213 B.n176 VSUBS 0.007057f
C214 B.n177 VSUBS 0.007057f
C215 B.n178 VSUBS 0.007057f
C216 B.n179 VSUBS 0.007057f
C217 B.n180 VSUBS 0.007057f
C218 B.n181 VSUBS 0.007057f
C219 B.n182 VSUBS 0.007057f
C220 B.n183 VSUBS 0.007057f
C221 B.n184 VSUBS 0.007057f
C222 B.n185 VSUBS 0.007057f
C223 B.n186 VSUBS 0.007057f
C224 B.n187 VSUBS 0.007057f
C225 B.n188 VSUBS 0.007057f
C226 B.n189 VSUBS 0.007057f
C227 B.n190 VSUBS 0.007057f
C228 B.n191 VSUBS 0.007057f
C229 B.n192 VSUBS 0.007057f
C230 B.n193 VSUBS 0.007057f
C231 B.n194 VSUBS 0.007057f
C232 B.n195 VSUBS 0.007057f
C233 B.n196 VSUBS 0.007057f
C234 B.n197 VSUBS 0.007057f
C235 B.n198 VSUBS 0.007057f
C236 B.n199 VSUBS 0.007057f
C237 B.n200 VSUBS 0.007057f
C238 B.n201 VSUBS 0.007057f
C239 B.n202 VSUBS 0.007057f
C240 B.n203 VSUBS 0.007057f
C241 B.n204 VSUBS 0.007057f
C242 B.n205 VSUBS 0.007057f
C243 B.n206 VSUBS 0.007057f
C244 B.n207 VSUBS 0.007057f
C245 B.n208 VSUBS 0.007057f
C246 B.n209 VSUBS 0.007057f
C247 B.n210 VSUBS 0.007057f
C248 B.n211 VSUBS 0.007057f
C249 B.n212 VSUBS 0.007057f
C250 B.n213 VSUBS 0.007057f
C251 B.n214 VSUBS 0.007057f
C252 B.n215 VSUBS 0.007057f
C253 B.n216 VSUBS 0.007057f
C254 B.n217 VSUBS 0.007057f
C255 B.n218 VSUBS 0.007057f
C256 B.n219 VSUBS 0.007057f
C257 B.n220 VSUBS 0.007057f
C258 B.n221 VSUBS 0.007057f
C259 B.n222 VSUBS 0.007057f
C260 B.n223 VSUBS 0.007057f
C261 B.n224 VSUBS 0.007057f
C262 B.n225 VSUBS 0.007057f
C263 B.n226 VSUBS 0.007057f
C264 B.n227 VSUBS 0.007057f
C265 B.n228 VSUBS 0.007057f
C266 B.n229 VSUBS 0.007057f
C267 B.n230 VSUBS 0.007057f
C268 B.n231 VSUBS 0.007057f
C269 B.n232 VSUBS 0.007057f
C270 B.n233 VSUBS 0.007057f
C271 B.n234 VSUBS 0.007057f
C272 B.n235 VSUBS 0.007057f
C273 B.n236 VSUBS 0.007057f
C274 B.n237 VSUBS 0.007057f
C275 B.n238 VSUBS 0.007057f
C276 B.n239 VSUBS 0.007057f
C277 B.n240 VSUBS 0.007057f
C278 B.n241 VSUBS 0.007057f
C279 B.n242 VSUBS 0.007057f
C280 B.n243 VSUBS 0.017233f
C281 B.n244 VSUBS 0.017846f
C282 B.n245 VSUBS 0.017846f
C283 B.n246 VSUBS 0.007057f
C284 B.n247 VSUBS 0.007057f
C285 B.n248 VSUBS 0.007057f
C286 B.n249 VSUBS 0.007057f
C287 B.n250 VSUBS 0.007057f
C288 B.n251 VSUBS 0.007057f
C289 B.n252 VSUBS 0.007057f
C290 B.n253 VSUBS 0.007057f
C291 B.n254 VSUBS 0.007057f
C292 B.n255 VSUBS 0.007057f
C293 B.n256 VSUBS 0.007057f
C294 B.n257 VSUBS 0.007057f
C295 B.n258 VSUBS 0.007057f
C296 B.n259 VSUBS 0.007057f
C297 B.n260 VSUBS 0.007057f
C298 B.n261 VSUBS 0.007057f
C299 B.n262 VSUBS 0.007057f
C300 B.n263 VSUBS 0.007057f
C301 B.n264 VSUBS 0.007057f
C302 B.n265 VSUBS 0.007057f
C303 B.n266 VSUBS 0.007057f
C304 B.n267 VSUBS 0.007057f
C305 B.n268 VSUBS 0.007057f
C306 B.n269 VSUBS 0.007057f
C307 B.n270 VSUBS 0.007057f
C308 B.n271 VSUBS 0.007057f
C309 B.n272 VSUBS 0.007057f
C310 B.n273 VSUBS 0.007057f
C311 B.n274 VSUBS 0.007057f
C312 B.n275 VSUBS 0.007057f
C313 B.n276 VSUBS 0.007057f
C314 B.n277 VSUBS 0.007057f
C315 B.n278 VSUBS 0.007057f
C316 B.n279 VSUBS 0.007057f
C317 B.n280 VSUBS 0.007057f
C318 B.n281 VSUBS 0.007057f
C319 B.n282 VSUBS 0.007057f
C320 B.n283 VSUBS 0.007057f
C321 B.n284 VSUBS 0.007057f
C322 B.n285 VSUBS 0.007057f
C323 B.n286 VSUBS 0.007057f
C324 B.n287 VSUBS 0.007057f
C325 B.n288 VSUBS 0.007057f
C326 B.n289 VSUBS 0.007057f
C327 B.n290 VSUBS 0.007057f
C328 B.n291 VSUBS 0.007057f
C329 B.n292 VSUBS 0.007057f
C330 B.n293 VSUBS 0.007057f
C331 B.n294 VSUBS 0.007057f
C332 B.n295 VSUBS 0.007057f
C333 B.n296 VSUBS 0.007057f
C334 B.n297 VSUBS 0.007057f
C335 B.n298 VSUBS 0.007057f
C336 B.n299 VSUBS 0.007057f
C337 B.n300 VSUBS 0.007057f
C338 B.n301 VSUBS 0.007057f
C339 B.n302 VSUBS 0.007057f
C340 B.n303 VSUBS 0.007057f
C341 B.n304 VSUBS 0.007057f
C342 B.n305 VSUBS 0.007057f
C343 B.n306 VSUBS 0.007057f
C344 B.n307 VSUBS 0.007057f
C345 B.n308 VSUBS 0.006642f
C346 B.n309 VSUBS 0.016351f
C347 B.n310 VSUBS 0.003944f
C348 B.n311 VSUBS 0.007057f
C349 B.n312 VSUBS 0.007057f
C350 B.n313 VSUBS 0.007057f
C351 B.n314 VSUBS 0.007057f
C352 B.n315 VSUBS 0.007057f
C353 B.n316 VSUBS 0.007057f
C354 B.n317 VSUBS 0.007057f
C355 B.n318 VSUBS 0.007057f
C356 B.n319 VSUBS 0.007057f
C357 B.n320 VSUBS 0.007057f
C358 B.n321 VSUBS 0.007057f
C359 B.n322 VSUBS 0.007057f
C360 B.t8 VSUBS 0.226302f
C361 B.t7 VSUBS 0.251214f
C362 B.t6 VSUBS 1.0601f
C363 B.n323 VSUBS 0.388678f
C364 B.n324 VSUBS 0.259579f
C365 B.n325 VSUBS 0.016351f
C366 B.n326 VSUBS 0.003944f
C367 B.n327 VSUBS 0.007057f
C368 B.n328 VSUBS 0.007057f
C369 B.n329 VSUBS 0.007057f
C370 B.n330 VSUBS 0.007057f
C371 B.n331 VSUBS 0.007057f
C372 B.n332 VSUBS 0.007057f
C373 B.n333 VSUBS 0.007057f
C374 B.n334 VSUBS 0.007057f
C375 B.n335 VSUBS 0.007057f
C376 B.n336 VSUBS 0.007057f
C377 B.n337 VSUBS 0.007057f
C378 B.n338 VSUBS 0.007057f
C379 B.n339 VSUBS 0.007057f
C380 B.n340 VSUBS 0.007057f
C381 B.n341 VSUBS 0.007057f
C382 B.n342 VSUBS 0.007057f
C383 B.n343 VSUBS 0.007057f
C384 B.n344 VSUBS 0.007057f
C385 B.n345 VSUBS 0.007057f
C386 B.n346 VSUBS 0.007057f
C387 B.n347 VSUBS 0.007057f
C388 B.n348 VSUBS 0.007057f
C389 B.n349 VSUBS 0.007057f
C390 B.n350 VSUBS 0.007057f
C391 B.n351 VSUBS 0.007057f
C392 B.n352 VSUBS 0.007057f
C393 B.n353 VSUBS 0.007057f
C394 B.n354 VSUBS 0.007057f
C395 B.n355 VSUBS 0.007057f
C396 B.n356 VSUBS 0.007057f
C397 B.n357 VSUBS 0.007057f
C398 B.n358 VSUBS 0.007057f
C399 B.n359 VSUBS 0.007057f
C400 B.n360 VSUBS 0.007057f
C401 B.n361 VSUBS 0.007057f
C402 B.n362 VSUBS 0.007057f
C403 B.n363 VSUBS 0.007057f
C404 B.n364 VSUBS 0.007057f
C405 B.n365 VSUBS 0.007057f
C406 B.n366 VSUBS 0.007057f
C407 B.n367 VSUBS 0.007057f
C408 B.n368 VSUBS 0.007057f
C409 B.n369 VSUBS 0.007057f
C410 B.n370 VSUBS 0.007057f
C411 B.n371 VSUBS 0.007057f
C412 B.n372 VSUBS 0.007057f
C413 B.n373 VSUBS 0.007057f
C414 B.n374 VSUBS 0.007057f
C415 B.n375 VSUBS 0.007057f
C416 B.n376 VSUBS 0.007057f
C417 B.n377 VSUBS 0.007057f
C418 B.n378 VSUBS 0.007057f
C419 B.n379 VSUBS 0.007057f
C420 B.n380 VSUBS 0.007057f
C421 B.n381 VSUBS 0.007057f
C422 B.n382 VSUBS 0.007057f
C423 B.n383 VSUBS 0.007057f
C424 B.n384 VSUBS 0.007057f
C425 B.n385 VSUBS 0.007057f
C426 B.n386 VSUBS 0.007057f
C427 B.n387 VSUBS 0.007057f
C428 B.n388 VSUBS 0.007057f
C429 B.n389 VSUBS 0.007057f
C430 B.n390 VSUBS 0.007057f
C431 B.n391 VSUBS 0.017084f
C432 B.n392 VSUBS 0.017995f
C433 B.n393 VSUBS 0.017233f
C434 B.n394 VSUBS 0.007057f
C435 B.n395 VSUBS 0.007057f
C436 B.n396 VSUBS 0.007057f
C437 B.n397 VSUBS 0.007057f
C438 B.n398 VSUBS 0.007057f
C439 B.n399 VSUBS 0.007057f
C440 B.n400 VSUBS 0.007057f
C441 B.n401 VSUBS 0.007057f
C442 B.n402 VSUBS 0.007057f
C443 B.n403 VSUBS 0.007057f
C444 B.n404 VSUBS 0.007057f
C445 B.n405 VSUBS 0.007057f
C446 B.n406 VSUBS 0.007057f
C447 B.n407 VSUBS 0.007057f
C448 B.n408 VSUBS 0.007057f
C449 B.n409 VSUBS 0.007057f
C450 B.n410 VSUBS 0.007057f
C451 B.n411 VSUBS 0.007057f
C452 B.n412 VSUBS 0.007057f
C453 B.n413 VSUBS 0.007057f
C454 B.n414 VSUBS 0.007057f
C455 B.n415 VSUBS 0.007057f
C456 B.n416 VSUBS 0.007057f
C457 B.n417 VSUBS 0.007057f
C458 B.n418 VSUBS 0.007057f
C459 B.n419 VSUBS 0.007057f
C460 B.n420 VSUBS 0.007057f
C461 B.n421 VSUBS 0.007057f
C462 B.n422 VSUBS 0.007057f
C463 B.n423 VSUBS 0.007057f
C464 B.n424 VSUBS 0.007057f
C465 B.n425 VSUBS 0.007057f
C466 B.n426 VSUBS 0.007057f
C467 B.n427 VSUBS 0.007057f
C468 B.n428 VSUBS 0.007057f
C469 B.n429 VSUBS 0.007057f
C470 B.n430 VSUBS 0.007057f
C471 B.n431 VSUBS 0.007057f
C472 B.n432 VSUBS 0.007057f
C473 B.n433 VSUBS 0.007057f
C474 B.n434 VSUBS 0.007057f
C475 B.n435 VSUBS 0.007057f
C476 B.n436 VSUBS 0.007057f
C477 B.n437 VSUBS 0.007057f
C478 B.n438 VSUBS 0.007057f
C479 B.n439 VSUBS 0.007057f
C480 B.n440 VSUBS 0.007057f
C481 B.n441 VSUBS 0.007057f
C482 B.n442 VSUBS 0.007057f
C483 B.n443 VSUBS 0.007057f
C484 B.n444 VSUBS 0.007057f
C485 B.n445 VSUBS 0.007057f
C486 B.n446 VSUBS 0.007057f
C487 B.n447 VSUBS 0.007057f
C488 B.n448 VSUBS 0.007057f
C489 B.n449 VSUBS 0.007057f
C490 B.n450 VSUBS 0.007057f
C491 B.n451 VSUBS 0.007057f
C492 B.n452 VSUBS 0.007057f
C493 B.n453 VSUBS 0.007057f
C494 B.n454 VSUBS 0.007057f
C495 B.n455 VSUBS 0.007057f
C496 B.n456 VSUBS 0.007057f
C497 B.n457 VSUBS 0.007057f
C498 B.n458 VSUBS 0.007057f
C499 B.n459 VSUBS 0.007057f
C500 B.n460 VSUBS 0.007057f
C501 B.n461 VSUBS 0.007057f
C502 B.n462 VSUBS 0.007057f
C503 B.n463 VSUBS 0.007057f
C504 B.n464 VSUBS 0.007057f
C505 B.n465 VSUBS 0.007057f
C506 B.n466 VSUBS 0.007057f
C507 B.n467 VSUBS 0.007057f
C508 B.n468 VSUBS 0.007057f
C509 B.n469 VSUBS 0.007057f
C510 B.n470 VSUBS 0.007057f
C511 B.n471 VSUBS 0.007057f
C512 B.n472 VSUBS 0.007057f
C513 B.n473 VSUBS 0.007057f
C514 B.n474 VSUBS 0.007057f
C515 B.n475 VSUBS 0.007057f
C516 B.n476 VSUBS 0.007057f
C517 B.n477 VSUBS 0.007057f
C518 B.n478 VSUBS 0.007057f
C519 B.n479 VSUBS 0.007057f
C520 B.n480 VSUBS 0.007057f
C521 B.n481 VSUBS 0.007057f
C522 B.n482 VSUBS 0.007057f
C523 B.n483 VSUBS 0.007057f
C524 B.n484 VSUBS 0.007057f
C525 B.n485 VSUBS 0.007057f
C526 B.n486 VSUBS 0.007057f
C527 B.n487 VSUBS 0.007057f
C528 B.n488 VSUBS 0.007057f
C529 B.n489 VSUBS 0.007057f
C530 B.n490 VSUBS 0.007057f
C531 B.n491 VSUBS 0.007057f
C532 B.n492 VSUBS 0.007057f
C533 B.n493 VSUBS 0.007057f
C534 B.n494 VSUBS 0.007057f
C535 B.n495 VSUBS 0.007057f
C536 B.n496 VSUBS 0.007057f
C537 B.n497 VSUBS 0.007057f
C538 B.n498 VSUBS 0.007057f
C539 B.n499 VSUBS 0.007057f
C540 B.n500 VSUBS 0.007057f
C541 B.n501 VSUBS 0.007057f
C542 B.n502 VSUBS 0.007057f
C543 B.n503 VSUBS 0.007057f
C544 B.n504 VSUBS 0.007057f
C545 B.n505 VSUBS 0.007057f
C546 B.n506 VSUBS 0.007057f
C547 B.n507 VSUBS 0.007057f
C548 B.n508 VSUBS 0.007057f
C549 B.n509 VSUBS 0.007057f
C550 B.n510 VSUBS 0.007057f
C551 B.n511 VSUBS 0.007057f
C552 B.n512 VSUBS 0.007057f
C553 B.n513 VSUBS 0.007057f
C554 B.n514 VSUBS 0.017233f
C555 B.n515 VSUBS 0.017846f
C556 B.n516 VSUBS 0.017846f
C557 B.n517 VSUBS 0.007057f
C558 B.n518 VSUBS 0.007057f
C559 B.n519 VSUBS 0.007057f
C560 B.n520 VSUBS 0.007057f
C561 B.n521 VSUBS 0.007057f
C562 B.n522 VSUBS 0.007057f
C563 B.n523 VSUBS 0.007057f
C564 B.n524 VSUBS 0.007057f
C565 B.n525 VSUBS 0.007057f
C566 B.n526 VSUBS 0.007057f
C567 B.n527 VSUBS 0.007057f
C568 B.n528 VSUBS 0.007057f
C569 B.n529 VSUBS 0.007057f
C570 B.n530 VSUBS 0.007057f
C571 B.n531 VSUBS 0.007057f
C572 B.n532 VSUBS 0.007057f
C573 B.n533 VSUBS 0.007057f
C574 B.n534 VSUBS 0.007057f
C575 B.n535 VSUBS 0.007057f
C576 B.n536 VSUBS 0.007057f
C577 B.n537 VSUBS 0.007057f
C578 B.n538 VSUBS 0.007057f
C579 B.n539 VSUBS 0.007057f
C580 B.n540 VSUBS 0.007057f
C581 B.n541 VSUBS 0.007057f
C582 B.n542 VSUBS 0.007057f
C583 B.n543 VSUBS 0.007057f
C584 B.n544 VSUBS 0.007057f
C585 B.n545 VSUBS 0.007057f
C586 B.n546 VSUBS 0.007057f
C587 B.n547 VSUBS 0.007057f
C588 B.n548 VSUBS 0.007057f
C589 B.n549 VSUBS 0.007057f
C590 B.n550 VSUBS 0.007057f
C591 B.n551 VSUBS 0.007057f
C592 B.n552 VSUBS 0.007057f
C593 B.n553 VSUBS 0.007057f
C594 B.n554 VSUBS 0.007057f
C595 B.n555 VSUBS 0.007057f
C596 B.n556 VSUBS 0.007057f
C597 B.n557 VSUBS 0.007057f
C598 B.n558 VSUBS 0.007057f
C599 B.n559 VSUBS 0.007057f
C600 B.n560 VSUBS 0.007057f
C601 B.n561 VSUBS 0.007057f
C602 B.n562 VSUBS 0.007057f
C603 B.n563 VSUBS 0.007057f
C604 B.n564 VSUBS 0.007057f
C605 B.n565 VSUBS 0.007057f
C606 B.n566 VSUBS 0.007057f
C607 B.n567 VSUBS 0.007057f
C608 B.n568 VSUBS 0.007057f
C609 B.n569 VSUBS 0.007057f
C610 B.n570 VSUBS 0.007057f
C611 B.n571 VSUBS 0.007057f
C612 B.n572 VSUBS 0.007057f
C613 B.n573 VSUBS 0.007057f
C614 B.n574 VSUBS 0.007057f
C615 B.n575 VSUBS 0.007057f
C616 B.n576 VSUBS 0.007057f
C617 B.n577 VSUBS 0.007057f
C618 B.n578 VSUBS 0.006642f
C619 B.n579 VSUBS 0.007057f
C620 B.n580 VSUBS 0.007057f
C621 B.n581 VSUBS 0.007057f
C622 B.n582 VSUBS 0.007057f
C623 B.n583 VSUBS 0.007057f
C624 B.n584 VSUBS 0.007057f
C625 B.n585 VSUBS 0.007057f
C626 B.n586 VSUBS 0.007057f
C627 B.n587 VSUBS 0.007057f
C628 B.n588 VSUBS 0.007057f
C629 B.n589 VSUBS 0.007057f
C630 B.n590 VSUBS 0.007057f
C631 B.n591 VSUBS 0.007057f
C632 B.n592 VSUBS 0.007057f
C633 B.n593 VSUBS 0.007057f
C634 B.n594 VSUBS 0.003944f
C635 B.n595 VSUBS 0.016351f
C636 B.n596 VSUBS 0.006642f
C637 B.n597 VSUBS 0.007057f
C638 B.n598 VSUBS 0.007057f
C639 B.n599 VSUBS 0.007057f
C640 B.n600 VSUBS 0.007057f
C641 B.n601 VSUBS 0.007057f
C642 B.n602 VSUBS 0.007057f
C643 B.n603 VSUBS 0.007057f
C644 B.n604 VSUBS 0.007057f
C645 B.n605 VSUBS 0.007057f
C646 B.n606 VSUBS 0.007057f
C647 B.n607 VSUBS 0.007057f
C648 B.n608 VSUBS 0.007057f
C649 B.n609 VSUBS 0.007057f
C650 B.n610 VSUBS 0.007057f
C651 B.n611 VSUBS 0.007057f
C652 B.n612 VSUBS 0.007057f
C653 B.n613 VSUBS 0.007057f
C654 B.n614 VSUBS 0.007057f
C655 B.n615 VSUBS 0.007057f
C656 B.n616 VSUBS 0.007057f
C657 B.n617 VSUBS 0.007057f
C658 B.n618 VSUBS 0.007057f
C659 B.n619 VSUBS 0.007057f
C660 B.n620 VSUBS 0.007057f
C661 B.n621 VSUBS 0.007057f
C662 B.n622 VSUBS 0.007057f
C663 B.n623 VSUBS 0.007057f
C664 B.n624 VSUBS 0.007057f
C665 B.n625 VSUBS 0.007057f
C666 B.n626 VSUBS 0.007057f
C667 B.n627 VSUBS 0.007057f
C668 B.n628 VSUBS 0.007057f
C669 B.n629 VSUBS 0.007057f
C670 B.n630 VSUBS 0.007057f
C671 B.n631 VSUBS 0.007057f
C672 B.n632 VSUBS 0.007057f
C673 B.n633 VSUBS 0.007057f
C674 B.n634 VSUBS 0.007057f
C675 B.n635 VSUBS 0.007057f
C676 B.n636 VSUBS 0.007057f
C677 B.n637 VSUBS 0.007057f
C678 B.n638 VSUBS 0.007057f
C679 B.n639 VSUBS 0.007057f
C680 B.n640 VSUBS 0.007057f
C681 B.n641 VSUBS 0.007057f
C682 B.n642 VSUBS 0.007057f
C683 B.n643 VSUBS 0.007057f
C684 B.n644 VSUBS 0.007057f
C685 B.n645 VSUBS 0.007057f
C686 B.n646 VSUBS 0.007057f
C687 B.n647 VSUBS 0.007057f
C688 B.n648 VSUBS 0.007057f
C689 B.n649 VSUBS 0.007057f
C690 B.n650 VSUBS 0.007057f
C691 B.n651 VSUBS 0.007057f
C692 B.n652 VSUBS 0.007057f
C693 B.n653 VSUBS 0.007057f
C694 B.n654 VSUBS 0.007057f
C695 B.n655 VSUBS 0.007057f
C696 B.n656 VSUBS 0.007057f
C697 B.n657 VSUBS 0.007057f
C698 B.n658 VSUBS 0.007057f
C699 B.n659 VSUBS 0.017846f
C700 B.n660 VSUBS 0.017233f
C701 B.n661 VSUBS 0.017233f
C702 B.n662 VSUBS 0.007057f
C703 B.n663 VSUBS 0.007057f
C704 B.n664 VSUBS 0.007057f
C705 B.n665 VSUBS 0.007057f
C706 B.n666 VSUBS 0.007057f
C707 B.n667 VSUBS 0.007057f
C708 B.n668 VSUBS 0.007057f
C709 B.n669 VSUBS 0.007057f
C710 B.n670 VSUBS 0.007057f
C711 B.n671 VSUBS 0.007057f
C712 B.n672 VSUBS 0.007057f
C713 B.n673 VSUBS 0.007057f
C714 B.n674 VSUBS 0.007057f
C715 B.n675 VSUBS 0.007057f
C716 B.n676 VSUBS 0.007057f
C717 B.n677 VSUBS 0.007057f
C718 B.n678 VSUBS 0.007057f
C719 B.n679 VSUBS 0.007057f
C720 B.n680 VSUBS 0.007057f
C721 B.n681 VSUBS 0.007057f
C722 B.n682 VSUBS 0.007057f
C723 B.n683 VSUBS 0.007057f
C724 B.n684 VSUBS 0.007057f
C725 B.n685 VSUBS 0.007057f
C726 B.n686 VSUBS 0.007057f
C727 B.n687 VSUBS 0.007057f
C728 B.n688 VSUBS 0.007057f
C729 B.n689 VSUBS 0.007057f
C730 B.n690 VSUBS 0.007057f
C731 B.n691 VSUBS 0.007057f
C732 B.n692 VSUBS 0.007057f
C733 B.n693 VSUBS 0.007057f
C734 B.n694 VSUBS 0.007057f
C735 B.n695 VSUBS 0.007057f
C736 B.n696 VSUBS 0.007057f
C737 B.n697 VSUBS 0.007057f
C738 B.n698 VSUBS 0.007057f
C739 B.n699 VSUBS 0.007057f
C740 B.n700 VSUBS 0.007057f
C741 B.n701 VSUBS 0.007057f
C742 B.n702 VSUBS 0.007057f
C743 B.n703 VSUBS 0.007057f
C744 B.n704 VSUBS 0.007057f
C745 B.n705 VSUBS 0.007057f
C746 B.n706 VSUBS 0.007057f
C747 B.n707 VSUBS 0.007057f
C748 B.n708 VSUBS 0.007057f
C749 B.n709 VSUBS 0.007057f
C750 B.n710 VSUBS 0.007057f
C751 B.n711 VSUBS 0.007057f
C752 B.n712 VSUBS 0.007057f
C753 B.n713 VSUBS 0.007057f
C754 B.n714 VSUBS 0.007057f
C755 B.n715 VSUBS 0.007057f
C756 B.n716 VSUBS 0.007057f
C757 B.n717 VSUBS 0.007057f
C758 B.n718 VSUBS 0.007057f
C759 B.n719 VSUBS 0.00921f
C760 B.n720 VSUBS 0.00981f
C761 B.n721 VSUBS 0.019509f
C762 VDD1.t0 VSUBS 0.248393f
C763 VDD1.t7 VSUBS 0.248393f
C764 VDD1.n0 VSUBS 1.98237f
C765 VDD1.t1 VSUBS 0.248393f
C766 VDD1.t3 VSUBS 0.248393f
C767 VDD1.n1 VSUBS 1.98124f
C768 VDD1.t5 VSUBS 0.248393f
C769 VDD1.t6 VSUBS 0.248393f
C770 VDD1.n2 VSUBS 1.98124f
C771 VDD1.n3 VSUBS 3.43522f
C772 VDD1.t4 VSUBS 0.248393f
C773 VDD1.t2 VSUBS 0.248393f
C774 VDD1.n4 VSUBS 1.9731f
C775 VDD1.n5 VSUBS 3.01785f
C776 VP.n0 VSUBS 0.034972f
C777 VP.t1 VSUBS 2.26206f
C778 VP.n1 VSUBS 0.028997f
C779 VP.n2 VSUBS 0.034972f
C780 VP.t2 VSUBS 2.26206f
C781 VP.n3 VSUBS 0.051053f
C782 VP.n4 VSUBS 0.034972f
C783 VP.t4 VSUBS 2.26206f
C784 VP.n5 VSUBS 0.067776f
C785 VP.n6 VSUBS 0.034972f
C786 VP.t6 VSUBS 2.26206f
C787 VP.n7 VSUBS 0.889549f
C788 VP.n8 VSUBS 0.034972f
C789 VP.t5 VSUBS 2.26206f
C790 VP.n9 VSUBS 0.028997f
C791 VP.n10 VSUBS 0.034972f
C792 VP.t3 VSUBS 2.26206f
C793 VP.n11 VSUBS 0.051053f
C794 VP.n12 VSUBS 0.259568f
C795 VP.t0 VSUBS 2.26206f
C796 VP.t7 VSUBS 2.43139f
C797 VP.n13 VSUBS 0.887573f
C798 VP.n14 VSUBS 0.893285f
C799 VP.n15 VSUBS 0.055846f
C800 VP.n16 VSUBS 0.051053f
C801 VP.n17 VSUBS 0.034972f
C802 VP.n18 VSUBS 0.034972f
C803 VP.n19 VSUBS 0.034972f
C804 VP.n20 VSUBS 0.055846f
C805 VP.n21 VSUBS 0.806669f
C806 VP.n22 VSUBS 0.04233f
C807 VP.n23 VSUBS 0.067776f
C808 VP.n24 VSUBS 0.034972f
C809 VP.n25 VSUBS 0.034972f
C810 VP.n26 VSUBS 0.034972f
C811 VP.n27 VSUBS 0.070513f
C812 VP.n28 VSUBS 0.037182f
C813 VP.n29 VSUBS 0.889549f
C814 VP.n30 VSUBS 1.7923f
C815 VP.n31 VSUBS 1.81854f
C816 VP.n32 VSUBS 0.034972f
C817 VP.n33 VSUBS 0.037182f
C818 VP.n34 VSUBS 0.070513f
C819 VP.n35 VSUBS 0.028997f
C820 VP.n36 VSUBS 0.034972f
C821 VP.n37 VSUBS 0.034972f
C822 VP.n38 VSUBS 0.034972f
C823 VP.n39 VSUBS 0.04233f
C824 VP.n40 VSUBS 0.806669f
C825 VP.n41 VSUBS 0.055846f
C826 VP.n42 VSUBS 0.051053f
C827 VP.n43 VSUBS 0.034972f
C828 VP.n44 VSUBS 0.034972f
C829 VP.n45 VSUBS 0.034972f
C830 VP.n46 VSUBS 0.055846f
C831 VP.n47 VSUBS 0.806669f
C832 VP.n48 VSUBS 0.04233f
C833 VP.n49 VSUBS 0.067776f
C834 VP.n50 VSUBS 0.034972f
C835 VP.n51 VSUBS 0.034972f
C836 VP.n52 VSUBS 0.034972f
C837 VP.n53 VSUBS 0.070513f
C838 VP.n54 VSUBS 0.037182f
C839 VP.n55 VSUBS 0.889549f
C840 VP.n56 VSUBS 0.03804f
C841 VDD2.t6 VSUBS 0.245374f
C842 VDD2.t5 VSUBS 0.245374f
C843 VDD2.n0 VSUBS 1.95716f
C844 VDD2.t3 VSUBS 0.245374f
C845 VDD2.t2 VSUBS 0.245374f
C846 VDD2.n1 VSUBS 1.95716f
C847 VDD2.n2 VSUBS 3.34178f
C848 VDD2.t4 VSUBS 0.245374f
C849 VDD2.t7 VSUBS 0.245374f
C850 VDD2.n3 VSUBS 1.94913f
C851 VDD2.n4 VSUBS 2.95114f
C852 VDD2.t0 VSUBS 0.245374f
C853 VDD2.t1 VSUBS 0.245374f
C854 VDD2.n5 VSUBS 1.95712f
C855 VTAIL.t8 VSUBS 0.242312f
C856 VTAIL.t14 VSUBS 0.242312f
C857 VTAIL.n0 VSUBS 1.7999f
C858 VTAIL.n1 VSUBS 0.688398f
C859 VTAIL.n2 VSUBS 0.013671f
C860 VTAIL.n3 VSUBS 0.030885f
C861 VTAIL.n4 VSUBS 0.013835f
C862 VTAIL.n5 VSUBS 0.024317f
C863 VTAIL.n6 VSUBS 0.013067f
C864 VTAIL.n7 VSUBS 0.030885f
C865 VTAIL.n8 VSUBS 0.013835f
C866 VTAIL.n9 VSUBS 0.024317f
C867 VTAIL.n10 VSUBS 0.013067f
C868 VTAIL.n11 VSUBS 0.030885f
C869 VTAIL.n12 VSUBS 0.013835f
C870 VTAIL.n13 VSUBS 0.024317f
C871 VTAIL.n14 VSUBS 0.013067f
C872 VTAIL.n15 VSUBS 0.030885f
C873 VTAIL.n16 VSUBS 0.013835f
C874 VTAIL.n17 VSUBS 0.024317f
C875 VTAIL.n18 VSUBS 0.013067f
C876 VTAIL.n19 VSUBS 0.030885f
C877 VTAIL.n20 VSUBS 0.013835f
C878 VTAIL.n21 VSUBS 0.024317f
C879 VTAIL.n22 VSUBS 0.013067f
C880 VTAIL.n23 VSUBS 0.023164f
C881 VTAIL.n24 VSUBS 0.019648f
C882 VTAIL.t12 VSUBS 0.065976f
C883 VTAIL.n25 VSUBS 0.154272f
C884 VTAIL.n26 VSUBS 1.28884f
C885 VTAIL.n27 VSUBS 0.013067f
C886 VTAIL.n28 VSUBS 0.013835f
C887 VTAIL.n29 VSUBS 0.030885f
C888 VTAIL.n30 VSUBS 0.030885f
C889 VTAIL.n31 VSUBS 0.013835f
C890 VTAIL.n32 VSUBS 0.013067f
C891 VTAIL.n33 VSUBS 0.024317f
C892 VTAIL.n34 VSUBS 0.024317f
C893 VTAIL.n35 VSUBS 0.013067f
C894 VTAIL.n36 VSUBS 0.013835f
C895 VTAIL.n37 VSUBS 0.030885f
C896 VTAIL.n38 VSUBS 0.030885f
C897 VTAIL.n39 VSUBS 0.013835f
C898 VTAIL.n40 VSUBS 0.013067f
C899 VTAIL.n41 VSUBS 0.024317f
C900 VTAIL.n42 VSUBS 0.024317f
C901 VTAIL.n43 VSUBS 0.013067f
C902 VTAIL.n44 VSUBS 0.013835f
C903 VTAIL.n45 VSUBS 0.030885f
C904 VTAIL.n46 VSUBS 0.030885f
C905 VTAIL.n47 VSUBS 0.013835f
C906 VTAIL.n48 VSUBS 0.013067f
C907 VTAIL.n49 VSUBS 0.024317f
C908 VTAIL.n50 VSUBS 0.024317f
C909 VTAIL.n51 VSUBS 0.013067f
C910 VTAIL.n52 VSUBS 0.013835f
C911 VTAIL.n53 VSUBS 0.030885f
C912 VTAIL.n54 VSUBS 0.030885f
C913 VTAIL.n55 VSUBS 0.013835f
C914 VTAIL.n56 VSUBS 0.013067f
C915 VTAIL.n57 VSUBS 0.024317f
C916 VTAIL.n58 VSUBS 0.024317f
C917 VTAIL.n59 VSUBS 0.013067f
C918 VTAIL.n60 VSUBS 0.013835f
C919 VTAIL.n61 VSUBS 0.030885f
C920 VTAIL.n62 VSUBS 0.030885f
C921 VTAIL.n63 VSUBS 0.013835f
C922 VTAIL.n64 VSUBS 0.013067f
C923 VTAIL.n65 VSUBS 0.024317f
C924 VTAIL.n66 VSUBS 0.060526f
C925 VTAIL.n67 VSUBS 0.013067f
C926 VTAIL.n68 VSUBS 0.013835f
C927 VTAIL.n69 VSUBS 0.067752f
C928 VTAIL.n70 VSUBS 0.044484f
C929 VTAIL.n71 VSUBS 0.208925f
C930 VTAIL.n72 VSUBS 0.013671f
C931 VTAIL.n73 VSUBS 0.030885f
C932 VTAIL.n74 VSUBS 0.013835f
C933 VTAIL.n75 VSUBS 0.024317f
C934 VTAIL.n76 VSUBS 0.013067f
C935 VTAIL.n77 VSUBS 0.030885f
C936 VTAIL.n78 VSUBS 0.013835f
C937 VTAIL.n79 VSUBS 0.024317f
C938 VTAIL.n80 VSUBS 0.013067f
C939 VTAIL.n81 VSUBS 0.030885f
C940 VTAIL.n82 VSUBS 0.013835f
C941 VTAIL.n83 VSUBS 0.024317f
C942 VTAIL.n84 VSUBS 0.013067f
C943 VTAIL.n85 VSUBS 0.030885f
C944 VTAIL.n86 VSUBS 0.013835f
C945 VTAIL.n87 VSUBS 0.024317f
C946 VTAIL.n88 VSUBS 0.013067f
C947 VTAIL.n89 VSUBS 0.030885f
C948 VTAIL.n90 VSUBS 0.013835f
C949 VTAIL.n91 VSUBS 0.024317f
C950 VTAIL.n92 VSUBS 0.013067f
C951 VTAIL.n93 VSUBS 0.023164f
C952 VTAIL.n94 VSUBS 0.019648f
C953 VTAIL.t1 VSUBS 0.065976f
C954 VTAIL.n95 VSUBS 0.154272f
C955 VTAIL.n96 VSUBS 1.28884f
C956 VTAIL.n97 VSUBS 0.013067f
C957 VTAIL.n98 VSUBS 0.013835f
C958 VTAIL.n99 VSUBS 0.030885f
C959 VTAIL.n100 VSUBS 0.030885f
C960 VTAIL.n101 VSUBS 0.013835f
C961 VTAIL.n102 VSUBS 0.013067f
C962 VTAIL.n103 VSUBS 0.024317f
C963 VTAIL.n104 VSUBS 0.024317f
C964 VTAIL.n105 VSUBS 0.013067f
C965 VTAIL.n106 VSUBS 0.013835f
C966 VTAIL.n107 VSUBS 0.030885f
C967 VTAIL.n108 VSUBS 0.030885f
C968 VTAIL.n109 VSUBS 0.013835f
C969 VTAIL.n110 VSUBS 0.013067f
C970 VTAIL.n111 VSUBS 0.024317f
C971 VTAIL.n112 VSUBS 0.024317f
C972 VTAIL.n113 VSUBS 0.013067f
C973 VTAIL.n114 VSUBS 0.013835f
C974 VTAIL.n115 VSUBS 0.030885f
C975 VTAIL.n116 VSUBS 0.030885f
C976 VTAIL.n117 VSUBS 0.013835f
C977 VTAIL.n118 VSUBS 0.013067f
C978 VTAIL.n119 VSUBS 0.024317f
C979 VTAIL.n120 VSUBS 0.024317f
C980 VTAIL.n121 VSUBS 0.013067f
C981 VTAIL.n122 VSUBS 0.013835f
C982 VTAIL.n123 VSUBS 0.030885f
C983 VTAIL.n124 VSUBS 0.030885f
C984 VTAIL.n125 VSUBS 0.013835f
C985 VTAIL.n126 VSUBS 0.013067f
C986 VTAIL.n127 VSUBS 0.024317f
C987 VTAIL.n128 VSUBS 0.024317f
C988 VTAIL.n129 VSUBS 0.013067f
C989 VTAIL.n130 VSUBS 0.013835f
C990 VTAIL.n131 VSUBS 0.030885f
C991 VTAIL.n132 VSUBS 0.030885f
C992 VTAIL.n133 VSUBS 0.013835f
C993 VTAIL.n134 VSUBS 0.013067f
C994 VTAIL.n135 VSUBS 0.024317f
C995 VTAIL.n136 VSUBS 0.060526f
C996 VTAIL.n137 VSUBS 0.013067f
C997 VTAIL.n138 VSUBS 0.013835f
C998 VTAIL.n139 VSUBS 0.067752f
C999 VTAIL.n140 VSUBS 0.044484f
C1000 VTAIL.n141 VSUBS 0.208925f
C1001 VTAIL.t4 VSUBS 0.242312f
C1002 VTAIL.t5 VSUBS 0.242312f
C1003 VTAIL.n142 VSUBS 1.7999f
C1004 VTAIL.n143 VSUBS 0.833117f
C1005 VTAIL.n144 VSUBS 0.013671f
C1006 VTAIL.n145 VSUBS 0.030885f
C1007 VTAIL.n146 VSUBS 0.013835f
C1008 VTAIL.n147 VSUBS 0.024317f
C1009 VTAIL.n148 VSUBS 0.013067f
C1010 VTAIL.n149 VSUBS 0.030885f
C1011 VTAIL.n150 VSUBS 0.013835f
C1012 VTAIL.n151 VSUBS 0.024317f
C1013 VTAIL.n152 VSUBS 0.013067f
C1014 VTAIL.n153 VSUBS 0.030885f
C1015 VTAIL.n154 VSUBS 0.013835f
C1016 VTAIL.n155 VSUBS 0.024317f
C1017 VTAIL.n156 VSUBS 0.013067f
C1018 VTAIL.n157 VSUBS 0.030885f
C1019 VTAIL.n158 VSUBS 0.013835f
C1020 VTAIL.n159 VSUBS 0.024317f
C1021 VTAIL.n160 VSUBS 0.013067f
C1022 VTAIL.n161 VSUBS 0.030885f
C1023 VTAIL.n162 VSUBS 0.013835f
C1024 VTAIL.n163 VSUBS 0.024317f
C1025 VTAIL.n164 VSUBS 0.013067f
C1026 VTAIL.n165 VSUBS 0.023164f
C1027 VTAIL.n166 VSUBS 0.019648f
C1028 VTAIL.t0 VSUBS 0.065976f
C1029 VTAIL.n167 VSUBS 0.154272f
C1030 VTAIL.n168 VSUBS 1.28884f
C1031 VTAIL.n169 VSUBS 0.013067f
C1032 VTAIL.n170 VSUBS 0.013835f
C1033 VTAIL.n171 VSUBS 0.030885f
C1034 VTAIL.n172 VSUBS 0.030885f
C1035 VTAIL.n173 VSUBS 0.013835f
C1036 VTAIL.n174 VSUBS 0.013067f
C1037 VTAIL.n175 VSUBS 0.024317f
C1038 VTAIL.n176 VSUBS 0.024317f
C1039 VTAIL.n177 VSUBS 0.013067f
C1040 VTAIL.n178 VSUBS 0.013835f
C1041 VTAIL.n179 VSUBS 0.030885f
C1042 VTAIL.n180 VSUBS 0.030885f
C1043 VTAIL.n181 VSUBS 0.013835f
C1044 VTAIL.n182 VSUBS 0.013067f
C1045 VTAIL.n183 VSUBS 0.024317f
C1046 VTAIL.n184 VSUBS 0.024317f
C1047 VTAIL.n185 VSUBS 0.013067f
C1048 VTAIL.n186 VSUBS 0.013835f
C1049 VTAIL.n187 VSUBS 0.030885f
C1050 VTAIL.n188 VSUBS 0.030885f
C1051 VTAIL.n189 VSUBS 0.013835f
C1052 VTAIL.n190 VSUBS 0.013067f
C1053 VTAIL.n191 VSUBS 0.024317f
C1054 VTAIL.n192 VSUBS 0.024317f
C1055 VTAIL.n193 VSUBS 0.013067f
C1056 VTAIL.n194 VSUBS 0.013835f
C1057 VTAIL.n195 VSUBS 0.030885f
C1058 VTAIL.n196 VSUBS 0.030885f
C1059 VTAIL.n197 VSUBS 0.013835f
C1060 VTAIL.n198 VSUBS 0.013067f
C1061 VTAIL.n199 VSUBS 0.024317f
C1062 VTAIL.n200 VSUBS 0.024317f
C1063 VTAIL.n201 VSUBS 0.013067f
C1064 VTAIL.n202 VSUBS 0.013835f
C1065 VTAIL.n203 VSUBS 0.030885f
C1066 VTAIL.n204 VSUBS 0.030885f
C1067 VTAIL.n205 VSUBS 0.013835f
C1068 VTAIL.n206 VSUBS 0.013067f
C1069 VTAIL.n207 VSUBS 0.024317f
C1070 VTAIL.n208 VSUBS 0.060526f
C1071 VTAIL.n209 VSUBS 0.013067f
C1072 VTAIL.n210 VSUBS 0.013835f
C1073 VTAIL.n211 VSUBS 0.067752f
C1074 VTAIL.n212 VSUBS 0.044484f
C1075 VTAIL.n213 VSUBS 1.50347f
C1076 VTAIL.n214 VSUBS 0.013671f
C1077 VTAIL.n215 VSUBS 0.030885f
C1078 VTAIL.n216 VSUBS 0.013835f
C1079 VTAIL.n217 VSUBS 0.024317f
C1080 VTAIL.n218 VSUBS 0.013067f
C1081 VTAIL.n219 VSUBS 0.030885f
C1082 VTAIL.n220 VSUBS 0.013835f
C1083 VTAIL.n221 VSUBS 0.024317f
C1084 VTAIL.n222 VSUBS 0.013067f
C1085 VTAIL.n223 VSUBS 0.030885f
C1086 VTAIL.n224 VSUBS 0.013835f
C1087 VTAIL.n225 VSUBS 0.024317f
C1088 VTAIL.n226 VSUBS 0.013067f
C1089 VTAIL.n227 VSUBS 0.030885f
C1090 VTAIL.n228 VSUBS 0.013835f
C1091 VTAIL.n229 VSUBS 0.024317f
C1092 VTAIL.n230 VSUBS 0.013067f
C1093 VTAIL.n231 VSUBS 0.030885f
C1094 VTAIL.n232 VSUBS 0.013835f
C1095 VTAIL.n233 VSUBS 0.024317f
C1096 VTAIL.n234 VSUBS 0.013067f
C1097 VTAIL.n235 VSUBS 0.023164f
C1098 VTAIL.n236 VSUBS 0.019648f
C1099 VTAIL.t15 VSUBS 0.065976f
C1100 VTAIL.n237 VSUBS 0.154272f
C1101 VTAIL.n238 VSUBS 1.28884f
C1102 VTAIL.n239 VSUBS 0.013067f
C1103 VTAIL.n240 VSUBS 0.013835f
C1104 VTAIL.n241 VSUBS 0.030885f
C1105 VTAIL.n242 VSUBS 0.030885f
C1106 VTAIL.n243 VSUBS 0.013835f
C1107 VTAIL.n244 VSUBS 0.013067f
C1108 VTAIL.n245 VSUBS 0.024317f
C1109 VTAIL.n246 VSUBS 0.024317f
C1110 VTAIL.n247 VSUBS 0.013067f
C1111 VTAIL.n248 VSUBS 0.013835f
C1112 VTAIL.n249 VSUBS 0.030885f
C1113 VTAIL.n250 VSUBS 0.030885f
C1114 VTAIL.n251 VSUBS 0.013835f
C1115 VTAIL.n252 VSUBS 0.013067f
C1116 VTAIL.n253 VSUBS 0.024317f
C1117 VTAIL.n254 VSUBS 0.024317f
C1118 VTAIL.n255 VSUBS 0.013067f
C1119 VTAIL.n256 VSUBS 0.013835f
C1120 VTAIL.n257 VSUBS 0.030885f
C1121 VTAIL.n258 VSUBS 0.030885f
C1122 VTAIL.n259 VSUBS 0.013835f
C1123 VTAIL.n260 VSUBS 0.013067f
C1124 VTAIL.n261 VSUBS 0.024317f
C1125 VTAIL.n262 VSUBS 0.024317f
C1126 VTAIL.n263 VSUBS 0.013067f
C1127 VTAIL.n264 VSUBS 0.013835f
C1128 VTAIL.n265 VSUBS 0.030885f
C1129 VTAIL.n266 VSUBS 0.030885f
C1130 VTAIL.n267 VSUBS 0.013835f
C1131 VTAIL.n268 VSUBS 0.013067f
C1132 VTAIL.n269 VSUBS 0.024317f
C1133 VTAIL.n270 VSUBS 0.024317f
C1134 VTAIL.n271 VSUBS 0.013067f
C1135 VTAIL.n272 VSUBS 0.013835f
C1136 VTAIL.n273 VSUBS 0.030885f
C1137 VTAIL.n274 VSUBS 0.030885f
C1138 VTAIL.n275 VSUBS 0.013835f
C1139 VTAIL.n276 VSUBS 0.013067f
C1140 VTAIL.n277 VSUBS 0.024317f
C1141 VTAIL.n278 VSUBS 0.060526f
C1142 VTAIL.n279 VSUBS 0.013067f
C1143 VTAIL.n280 VSUBS 0.013835f
C1144 VTAIL.n281 VSUBS 0.067752f
C1145 VTAIL.n282 VSUBS 0.044484f
C1146 VTAIL.n283 VSUBS 1.50347f
C1147 VTAIL.t11 VSUBS 0.242312f
C1148 VTAIL.t10 VSUBS 0.242312f
C1149 VTAIL.n284 VSUBS 1.7999f
C1150 VTAIL.n285 VSUBS 0.833114f
C1151 VTAIL.n286 VSUBS 0.013671f
C1152 VTAIL.n287 VSUBS 0.030885f
C1153 VTAIL.n288 VSUBS 0.013835f
C1154 VTAIL.n289 VSUBS 0.024317f
C1155 VTAIL.n290 VSUBS 0.013067f
C1156 VTAIL.n291 VSUBS 0.030885f
C1157 VTAIL.n292 VSUBS 0.013835f
C1158 VTAIL.n293 VSUBS 0.024317f
C1159 VTAIL.n294 VSUBS 0.013067f
C1160 VTAIL.n295 VSUBS 0.030885f
C1161 VTAIL.n296 VSUBS 0.013835f
C1162 VTAIL.n297 VSUBS 0.024317f
C1163 VTAIL.n298 VSUBS 0.013067f
C1164 VTAIL.n299 VSUBS 0.030885f
C1165 VTAIL.n300 VSUBS 0.013835f
C1166 VTAIL.n301 VSUBS 0.024317f
C1167 VTAIL.n302 VSUBS 0.013067f
C1168 VTAIL.n303 VSUBS 0.030885f
C1169 VTAIL.n304 VSUBS 0.013835f
C1170 VTAIL.n305 VSUBS 0.024317f
C1171 VTAIL.n306 VSUBS 0.013067f
C1172 VTAIL.n307 VSUBS 0.023164f
C1173 VTAIL.n308 VSUBS 0.019648f
C1174 VTAIL.t9 VSUBS 0.065976f
C1175 VTAIL.n309 VSUBS 0.154272f
C1176 VTAIL.n310 VSUBS 1.28884f
C1177 VTAIL.n311 VSUBS 0.013067f
C1178 VTAIL.n312 VSUBS 0.013835f
C1179 VTAIL.n313 VSUBS 0.030885f
C1180 VTAIL.n314 VSUBS 0.030885f
C1181 VTAIL.n315 VSUBS 0.013835f
C1182 VTAIL.n316 VSUBS 0.013067f
C1183 VTAIL.n317 VSUBS 0.024317f
C1184 VTAIL.n318 VSUBS 0.024317f
C1185 VTAIL.n319 VSUBS 0.013067f
C1186 VTAIL.n320 VSUBS 0.013835f
C1187 VTAIL.n321 VSUBS 0.030885f
C1188 VTAIL.n322 VSUBS 0.030885f
C1189 VTAIL.n323 VSUBS 0.013835f
C1190 VTAIL.n324 VSUBS 0.013067f
C1191 VTAIL.n325 VSUBS 0.024317f
C1192 VTAIL.n326 VSUBS 0.024317f
C1193 VTAIL.n327 VSUBS 0.013067f
C1194 VTAIL.n328 VSUBS 0.013835f
C1195 VTAIL.n329 VSUBS 0.030885f
C1196 VTAIL.n330 VSUBS 0.030885f
C1197 VTAIL.n331 VSUBS 0.013835f
C1198 VTAIL.n332 VSUBS 0.013067f
C1199 VTAIL.n333 VSUBS 0.024317f
C1200 VTAIL.n334 VSUBS 0.024317f
C1201 VTAIL.n335 VSUBS 0.013067f
C1202 VTAIL.n336 VSUBS 0.013835f
C1203 VTAIL.n337 VSUBS 0.030885f
C1204 VTAIL.n338 VSUBS 0.030885f
C1205 VTAIL.n339 VSUBS 0.013835f
C1206 VTAIL.n340 VSUBS 0.013067f
C1207 VTAIL.n341 VSUBS 0.024317f
C1208 VTAIL.n342 VSUBS 0.024317f
C1209 VTAIL.n343 VSUBS 0.013067f
C1210 VTAIL.n344 VSUBS 0.013835f
C1211 VTAIL.n345 VSUBS 0.030885f
C1212 VTAIL.n346 VSUBS 0.030885f
C1213 VTAIL.n347 VSUBS 0.013835f
C1214 VTAIL.n348 VSUBS 0.013067f
C1215 VTAIL.n349 VSUBS 0.024317f
C1216 VTAIL.n350 VSUBS 0.060526f
C1217 VTAIL.n351 VSUBS 0.013067f
C1218 VTAIL.n352 VSUBS 0.013835f
C1219 VTAIL.n353 VSUBS 0.067752f
C1220 VTAIL.n354 VSUBS 0.044484f
C1221 VTAIL.n355 VSUBS 0.208925f
C1222 VTAIL.n356 VSUBS 0.013671f
C1223 VTAIL.n357 VSUBS 0.030885f
C1224 VTAIL.n358 VSUBS 0.013835f
C1225 VTAIL.n359 VSUBS 0.024317f
C1226 VTAIL.n360 VSUBS 0.013067f
C1227 VTAIL.n361 VSUBS 0.030885f
C1228 VTAIL.n362 VSUBS 0.013835f
C1229 VTAIL.n363 VSUBS 0.024317f
C1230 VTAIL.n364 VSUBS 0.013067f
C1231 VTAIL.n365 VSUBS 0.030885f
C1232 VTAIL.n366 VSUBS 0.013835f
C1233 VTAIL.n367 VSUBS 0.024317f
C1234 VTAIL.n368 VSUBS 0.013067f
C1235 VTAIL.n369 VSUBS 0.030885f
C1236 VTAIL.n370 VSUBS 0.013835f
C1237 VTAIL.n371 VSUBS 0.024317f
C1238 VTAIL.n372 VSUBS 0.013067f
C1239 VTAIL.n373 VSUBS 0.030885f
C1240 VTAIL.n374 VSUBS 0.013835f
C1241 VTAIL.n375 VSUBS 0.024317f
C1242 VTAIL.n376 VSUBS 0.013067f
C1243 VTAIL.n377 VSUBS 0.023164f
C1244 VTAIL.n378 VSUBS 0.019648f
C1245 VTAIL.t2 VSUBS 0.065976f
C1246 VTAIL.n379 VSUBS 0.154272f
C1247 VTAIL.n380 VSUBS 1.28884f
C1248 VTAIL.n381 VSUBS 0.013067f
C1249 VTAIL.n382 VSUBS 0.013835f
C1250 VTAIL.n383 VSUBS 0.030885f
C1251 VTAIL.n384 VSUBS 0.030885f
C1252 VTAIL.n385 VSUBS 0.013835f
C1253 VTAIL.n386 VSUBS 0.013067f
C1254 VTAIL.n387 VSUBS 0.024317f
C1255 VTAIL.n388 VSUBS 0.024317f
C1256 VTAIL.n389 VSUBS 0.013067f
C1257 VTAIL.n390 VSUBS 0.013835f
C1258 VTAIL.n391 VSUBS 0.030885f
C1259 VTAIL.n392 VSUBS 0.030885f
C1260 VTAIL.n393 VSUBS 0.013835f
C1261 VTAIL.n394 VSUBS 0.013067f
C1262 VTAIL.n395 VSUBS 0.024317f
C1263 VTAIL.n396 VSUBS 0.024317f
C1264 VTAIL.n397 VSUBS 0.013067f
C1265 VTAIL.n398 VSUBS 0.013835f
C1266 VTAIL.n399 VSUBS 0.030885f
C1267 VTAIL.n400 VSUBS 0.030885f
C1268 VTAIL.n401 VSUBS 0.013835f
C1269 VTAIL.n402 VSUBS 0.013067f
C1270 VTAIL.n403 VSUBS 0.024317f
C1271 VTAIL.n404 VSUBS 0.024317f
C1272 VTAIL.n405 VSUBS 0.013067f
C1273 VTAIL.n406 VSUBS 0.013835f
C1274 VTAIL.n407 VSUBS 0.030885f
C1275 VTAIL.n408 VSUBS 0.030885f
C1276 VTAIL.n409 VSUBS 0.013835f
C1277 VTAIL.n410 VSUBS 0.013067f
C1278 VTAIL.n411 VSUBS 0.024317f
C1279 VTAIL.n412 VSUBS 0.024317f
C1280 VTAIL.n413 VSUBS 0.013067f
C1281 VTAIL.n414 VSUBS 0.013835f
C1282 VTAIL.n415 VSUBS 0.030885f
C1283 VTAIL.n416 VSUBS 0.030885f
C1284 VTAIL.n417 VSUBS 0.013835f
C1285 VTAIL.n418 VSUBS 0.013067f
C1286 VTAIL.n419 VSUBS 0.024317f
C1287 VTAIL.n420 VSUBS 0.060526f
C1288 VTAIL.n421 VSUBS 0.013067f
C1289 VTAIL.n422 VSUBS 0.013835f
C1290 VTAIL.n423 VSUBS 0.067752f
C1291 VTAIL.n424 VSUBS 0.044484f
C1292 VTAIL.n425 VSUBS 0.208925f
C1293 VTAIL.t6 VSUBS 0.242312f
C1294 VTAIL.t7 VSUBS 0.242312f
C1295 VTAIL.n426 VSUBS 1.7999f
C1296 VTAIL.n427 VSUBS 0.833114f
C1297 VTAIL.n428 VSUBS 0.013671f
C1298 VTAIL.n429 VSUBS 0.030885f
C1299 VTAIL.n430 VSUBS 0.013835f
C1300 VTAIL.n431 VSUBS 0.024317f
C1301 VTAIL.n432 VSUBS 0.013067f
C1302 VTAIL.n433 VSUBS 0.030885f
C1303 VTAIL.n434 VSUBS 0.013835f
C1304 VTAIL.n435 VSUBS 0.024317f
C1305 VTAIL.n436 VSUBS 0.013067f
C1306 VTAIL.n437 VSUBS 0.030885f
C1307 VTAIL.n438 VSUBS 0.013835f
C1308 VTAIL.n439 VSUBS 0.024317f
C1309 VTAIL.n440 VSUBS 0.013067f
C1310 VTAIL.n441 VSUBS 0.030885f
C1311 VTAIL.n442 VSUBS 0.013835f
C1312 VTAIL.n443 VSUBS 0.024317f
C1313 VTAIL.n444 VSUBS 0.013067f
C1314 VTAIL.n445 VSUBS 0.030885f
C1315 VTAIL.n446 VSUBS 0.013835f
C1316 VTAIL.n447 VSUBS 0.024317f
C1317 VTAIL.n448 VSUBS 0.013067f
C1318 VTAIL.n449 VSUBS 0.023164f
C1319 VTAIL.n450 VSUBS 0.019648f
C1320 VTAIL.t3 VSUBS 0.065976f
C1321 VTAIL.n451 VSUBS 0.154272f
C1322 VTAIL.n452 VSUBS 1.28884f
C1323 VTAIL.n453 VSUBS 0.013067f
C1324 VTAIL.n454 VSUBS 0.013835f
C1325 VTAIL.n455 VSUBS 0.030885f
C1326 VTAIL.n456 VSUBS 0.030885f
C1327 VTAIL.n457 VSUBS 0.013835f
C1328 VTAIL.n458 VSUBS 0.013067f
C1329 VTAIL.n459 VSUBS 0.024317f
C1330 VTAIL.n460 VSUBS 0.024317f
C1331 VTAIL.n461 VSUBS 0.013067f
C1332 VTAIL.n462 VSUBS 0.013835f
C1333 VTAIL.n463 VSUBS 0.030885f
C1334 VTAIL.n464 VSUBS 0.030885f
C1335 VTAIL.n465 VSUBS 0.013835f
C1336 VTAIL.n466 VSUBS 0.013067f
C1337 VTAIL.n467 VSUBS 0.024317f
C1338 VTAIL.n468 VSUBS 0.024317f
C1339 VTAIL.n469 VSUBS 0.013067f
C1340 VTAIL.n470 VSUBS 0.013835f
C1341 VTAIL.n471 VSUBS 0.030885f
C1342 VTAIL.n472 VSUBS 0.030885f
C1343 VTAIL.n473 VSUBS 0.013835f
C1344 VTAIL.n474 VSUBS 0.013067f
C1345 VTAIL.n475 VSUBS 0.024317f
C1346 VTAIL.n476 VSUBS 0.024317f
C1347 VTAIL.n477 VSUBS 0.013067f
C1348 VTAIL.n478 VSUBS 0.013835f
C1349 VTAIL.n479 VSUBS 0.030885f
C1350 VTAIL.n480 VSUBS 0.030885f
C1351 VTAIL.n481 VSUBS 0.013835f
C1352 VTAIL.n482 VSUBS 0.013067f
C1353 VTAIL.n483 VSUBS 0.024317f
C1354 VTAIL.n484 VSUBS 0.024317f
C1355 VTAIL.n485 VSUBS 0.013067f
C1356 VTAIL.n486 VSUBS 0.013835f
C1357 VTAIL.n487 VSUBS 0.030885f
C1358 VTAIL.n488 VSUBS 0.030885f
C1359 VTAIL.n489 VSUBS 0.013835f
C1360 VTAIL.n490 VSUBS 0.013067f
C1361 VTAIL.n491 VSUBS 0.024317f
C1362 VTAIL.n492 VSUBS 0.060526f
C1363 VTAIL.n493 VSUBS 0.013067f
C1364 VTAIL.n494 VSUBS 0.013835f
C1365 VTAIL.n495 VSUBS 0.067752f
C1366 VTAIL.n496 VSUBS 0.044484f
C1367 VTAIL.n497 VSUBS 1.50347f
C1368 VTAIL.n498 VSUBS 0.013671f
C1369 VTAIL.n499 VSUBS 0.030885f
C1370 VTAIL.n500 VSUBS 0.013835f
C1371 VTAIL.n501 VSUBS 0.024317f
C1372 VTAIL.n502 VSUBS 0.013067f
C1373 VTAIL.n503 VSUBS 0.030885f
C1374 VTAIL.n504 VSUBS 0.013835f
C1375 VTAIL.n505 VSUBS 0.024317f
C1376 VTAIL.n506 VSUBS 0.013067f
C1377 VTAIL.n507 VSUBS 0.030885f
C1378 VTAIL.n508 VSUBS 0.013835f
C1379 VTAIL.n509 VSUBS 0.024317f
C1380 VTAIL.n510 VSUBS 0.013067f
C1381 VTAIL.n511 VSUBS 0.030885f
C1382 VTAIL.n512 VSUBS 0.013835f
C1383 VTAIL.n513 VSUBS 0.024317f
C1384 VTAIL.n514 VSUBS 0.013067f
C1385 VTAIL.n515 VSUBS 0.030885f
C1386 VTAIL.n516 VSUBS 0.013835f
C1387 VTAIL.n517 VSUBS 0.024317f
C1388 VTAIL.n518 VSUBS 0.013067f
C1389 VTAIL.n519 VSUBS 0.023164f
C1390 VTAIL.n520 VSUBS 0.019648f
C1391 VTAIL.t13 VSUBS 0.065976f
C1392 VTAIL.n521 VSUBS 0.154272f
C1393 VTAIL.n522 VSUBS 1.28884f
C1394 VTAIL.n523 VSUBS 0.013067f
C1395 VTAIL.n524 VSUBS 0.013835f
C1396 VTAIL.n525 VSUBS 0.030885f
C1397 VTAIL.n526 VSUBS 0.030885f
C1398 VTAIL.n527 VSUBS 0.013835f
C1399 VTAIL.n528 VSUBS 0.013067f
C1400 VTAIL.n529 VSUBS 0.024317f
C1401 VTAIL.n530 VSUBS 0.024317f
C1402 VTAIL.n531 VSUBS 0.013067f
C1403 VTAIL.n532 VSUBS 0.013835f
C1404 VTAIL.n533 VSUBS 0.030885f
C1405 VTAIL.n534 VSUBS 0.030885f
C1406 VTAIL.n535 VSUBS 0.013835f
C1407 VTAIL.n536 VSUBS 0.013067f
C1408 VTAIL.n537 VSUBS 0.024317f
C1409 VTAIL.n538 VSUBS 0.024317f
C1410 VTAIL.n539 VSUBS 0.013067f
C1411 VTAIL.n540 VSUBS 0.013835f
C1412 VTAIL.n541 VSUBS 0.030885f
C1413 VTAIL.n542 VSUBS 0.030885f
C1414 VTAIL.n543 VSUBS 0.013835f
C1415 VTAIL.n544 VSUBS 0.013067f
C1416 VTAIL.n545 VSUBS 0.024317f
C1417 VTAIL.n546 VSUBS 0.024317f
C1418 VTAIL.n547 VSUBS 0.013067f
C1419 VTAIL.n548 VSUBS 0.013835f
C1420 VTAIL.n549 VSUBS 0.030885f
C1421 VTAIL.n550 VSUBS 0.030885f
C1422 VTAIL.n551 VSUBS 0.013835f
C1423 VTAIL.n552 VSUBS 0.013067f
C1424 VTAIL.n553 VSUBS 0.024317f
C1425 VTAIL.n554 VSUBS 0.024317f
C1426 VTAIL.n555 VSUBS 0.013067f
C1427 VTAIL.n556 VSUBS 0.013835f
C1428 VTAIL.n557 VSUBS 0.030885f
C1429 VTAIL.n558 VSUBS 0.030885f
C1430 VTAIL.n559 VSUBS 0.013835f
C1431 VTAIL.n560 VSUBS 0.013067f
C1432 VTAIL.n561 VSUBS 0.024317f
C1433 VTAIL.n562 VSUBS 0.060526f
C1434 VTAIL.n563 VSUBS 0.013067f
C1435 VTAIL.n564 VSUBS 0.013835f
C1436 VTAIL.n565 VSUBS 0.067752f
C1437 VTAIL.n566 VSUBS 0.044484f
C1438 VTAIL.n567 VSUBS 1.49891f
C1439 VN.n0 VSUBS 0.034129f
C1440 VN.t5 VSUBS 2.20748f
C1441 VN.n1 VSUBS 0.028298f
C1442 VN.n2 VSUBS 0.034129f
C1443 VN.t4 VSUBS 2.20748f
C1444 VN.n3 VSUBS 0.049821f
C1445 VN.n4 VSUBS 0.253305f
C1446 VN.t2 VSUBS 2.20748f
C1447 VN.t1 VSUBS 2.37272f
C1448 VN.n5 VSUBS 0.866157f
C1449 VN.n6 VSUBS 0.871731f
C1450 VN.n7 VSUBS 0.054499f
C1451 VN.n8 VSUBS 0.049821f
C1452 VN.n9 VSUBS 0.034129f
C1453 VN.n10 VSUBS 0.034129f
C1454 VN.n11 VSUBS 0.034129f
C1455 VN.n12 VSUBS 0.054499f
C1456 VN.n13 VSUBS 0.787205f
C1457 VN.n14 VSUBS 0.041309f
C1458 VN.n15 VSUBS 0.06614f
C1459 VN.n16 VSUBS 0.034129f
C1460 VN.n17 VSUBS 0.034129f
C1461 VN.n18 VSUBS 0.034129f
C1462 VN.n19 VSUBS 0.068812f
C1463 VN.n20 VSUBS 0.036285f
C1464 VN.n21 VSUBS 0.868086f
C1465 VN.n22 VSUBS 0.037122f
C1466 VN.n23 VSUBS 0.034129f
C1467 VN.t3 VSUBS 2.20748f
C1468 VN.n24 VSUBS 0.028298f
C1469 VN.n25 VSUBS 0.034129f
C1470 VN.t0 VSUBS 2.20748f
C1471 VN.n26 VSUBS 0.049821f
C1472 VN.n27 VSUBS 0.253305f
C1473 VN.t7 VSUBS 2.20748f
C1474 VN.t6 VSUBS 2.37272f
C1475 VN.n28 VSUBS 0.866157f
C1476 VN.n29 VSUBS 0.871731f
C1477 VN.n30 VSUBS 0.054499f
C1478 VN.n31 VSUBS 0.049821f
C1479 VN.n32 VSUBS 0.034129f
C1480 VN.n33 VSUBS 0.034129f
C1481 VN.n34 VSUBS 0.034129f
C1482 VN.n35 VSUBS 0.054499f
C1483 VN.n36 VSUBS 0.787205f
C1484 VN.n37 VSUBS 0.041309f
C1485 VN.n38 VSUBS 0.06614f
C1486 VN.n39 VSUBS 0.034129f
C1487 VN.n40 VSUBS 0.034129f
C1488 VN.n41 VSUBS 0.034129f
C1489 VN.n42 VSUBS 0.068812f
C1490 VN.n43 VSUBS 0.036285f
C1491 VN.n44 VSUBS 0.868086f
C1492 VN.n45 VSUBS 1.77129f
.ends

