* NGSPICE file created from diff_pair_sample_1326.ext - technology: sky130A

.subckt diff_pair_sample_1326 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=4.9374 ps=26.1 w=12.66 l=0.95
X1 B.t22 B.t20 B.t21 B.t14 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=0.95
X2 VDD2.t9 VN.t0 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X3 VDD1.t8 VP.t1 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=2.0889 ps=12.99 w=12.66 l=0.95
X4 VDD2.t8 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X5 VTAIL.t5 VN.t2 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X6 B.t19 B.t17 B.t18 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=0.95
X7 VDD1.t7 VP.t2 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=4.9374 ps=26.1 w=12.66 l=0.95
X8 VDD1.t6 VP.t3 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=2.0889 ps=12.99 w=12.66 l=0.95
X9 VTAIL.t17 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X10 VDD2.t6 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=2.0889 ps=12.99 w=12.66 l=0.95
X11 VDD2.t5 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=4.9374 ps=26.1 w=12.66 l=0.95
X12 VTAIL.t19 VN.t5 VDD2.t4 B.t23 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X13 VTAIL.t11 VP.t5 VDD1.t4 B.t23 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X14 VDD1.t3 VP.t6 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X15 VDD1.t2 VP.t7 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X16 VTAIL.t2 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X17 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=4.9374 ps=26.1 w=12.66 l=0.95
X18 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=0.95
X19 VTAIL.t14 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X20 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=0.95
X21 VTAIL.t15 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
X22 VDD2.t1 VN.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9374 pd=26.1 as=2.0889 ps=12.99 w=12.66 l=0.95
X23 VTAIL.t1 VN.t9 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0889 pd=12.99 as=2.0889 ps=12.99 w=12.66 l=0.95
R0 VP.n10 VP.t1 382.909
R1 VP.n5 VP.t3 362.515
R2 VP.n41 VP.t0 362.515
R3 VP.n23 VP.t2 362.515
R4 VP.n34 VP.t7 321.164
R5 VP.n29 VP.t5 321.164
R6 VP.n1 VP.t9 321.164
R7 VP.n16 VP.t6 321.164
R8 VP.n7 VP.t8 321.164
R9 VP.n11 VP.t4 321.164
R10 VP.n42 VP.n41 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n9 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n8 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n40 VP.n0 161.3
R20 VP.n39 VP.n38 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n25 VP.n5 161.3
R29 VP.n30 VP.n3 54.1398
R30 VP.n36 VP.n35 54.1398
R31 VP.n18 VP.n17 54.1398
R32 VP.n12 VP.n9 54.1398
R33 VP.n28 VP.n27 48.3272
R34 VP.n40 VP.n39 48.3272
R35 VP.n22 VP.n21 48.3272
R36 VP.n25 VP.n24 44.705
R37 VP.n13 VP.n10 43.0014
R38 VP.n11 VP.n10 40.664
R39 VP.n34 VP.n3 27.0143
R40 VP.n35 VP.n34 27.0143
R41 VP.n17 VP.n16 27.0143
R42 VP.n16 VP.n9 27.0143
R43 VP.n30 VP.n29 13.7719
R44 VP.n36 VP.n1 13.7719
R45 VP.n18 VP.n7 13.7719
R46 VP.n12 VP.n11 13.7719
R47 VP.n27 VP.n5 12.4157
R48 VP.n41 VP.n40 12.4157
R49 VP.n23 VP.n22 12.4157
R50 VP.n29 VP.n28 10.8209
R51 VP.n39 VP.n1 10.8209
R52 VP.n21 VP.n7 10.8209
R53 VP.n14 VP.n13 0.189894
R54 VP.n15 VP.n14 0.189894
R55 VP.n15 VP.n8 0.189894
R56 VP.n19 VP.n8 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n37 VP.n2 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n38 VP.n0 0.189894
R69 VP.n42 VP.n0 0.189894
R70 VP VP.n42 0.0516364
R71 VTAIL.n292 VTAIL.n291 289.615
R72 VTAIL.n70 VTAIL.n69 289.615
R73 VTAIL.n222 VTAIL.n221 289.615
R74 VTAIL.n148 VTAIL.n147 289.615
R75 VTAIL.n246 VTAIL.n245 185
R76 VTAIL.n251 VTAIL.n250 185
R77 VTAIL.n253 VTAIL.n252 185
R78 VTAIL.n242 VTAIL.n241 185
R79 VTAIL.n259 VTAIL.n258 185
R80 VTAIL.n261 VTAIL.n260 185
R81 VTAIL.n238 VTAIL.n237 185
R82 VTAIL.n267 VTAIL.n266 185
R83 VTAIL.n269 VTAIL.n268 185
R84 VTAIL.n234 VTAIL.n233 185
R85 VTAIL.n275 VTAIL.n274 185
R86 VTAIL.n277 VTAIL.n276 185
R87 VTAIL.n230 VTAIL.n229 185
R88 VTAIL.n283 VTAIL.n282 185
R89 VTAIL.n285 VTAIL.n284 185
R90 VTAIL.n226 VTAIL.n225 185
R91 VTAIL.n291 VTAIL.n290 185
R92 VTAIL.n24 VTAIL.n23 185
R93 VTAIL.n29 VTAIL.n28 185
R94 VTAIL.n31 VTAIL.n30 185
R95 VTAIL.n20 VTAIL.n19 185
R96 VTAIL.n37 VTAIL.n36 185
R97 VTAIL.n39 VTAIL.n38 185
R98 VTAIL.n16 VTAIL.n15 185
R99 VTAIL.n45 VTAIL.n44 185
R100 VTAIL.n47 VTAIL.n46 185
R101 VTAIL.n12 VTAIL.n11 185
R102 VTAIL.n53 VTAIL.n52 185
R103 VTAIL.n55 VTAIL.n54 185
R104 VTAIL.n8 VTAIL.n7 185
R105 VTAIL.n61 VTAIL.n60 185
R106 VTAIL.n63 VTAIL.n62 185
R107 VTAIL.n4 VTAIL.n3 185
R108 VTAIL.n69 VTAIL.n68 185
R109 VTAIL.n221 VTAIL.n220 185
R110 VTAIL.n156 VTAIL.n155 185
R111 VTAIL.n215 VTAIL.n214 185
R112 VTAIL.n213 VTAIL.n212 185
R113 VTAIL.n160 VTAIL.n159 185
R114 VTAIL.n207 VTAIL.n206 185
R115 VTAIL.n205 VTAIL.n204 185
R116 VTAIL.n164 VTAIL.n163 185
R117 VTAIL.n199 VTAIL.n198 185
R118 VTAIL.n197 VTAIL.n196 185
R119 VTAIL.n168 VTAIL.n167 185
R120 VTAIL.n191 VTAIL.n190 185
R121 VTAIL.n189 VTAIL.n188 185
R122 VTAIL.n172 VTAIL.n171 185
R123 VTAIL.n183 VTAIL.n182 185
R124 VTAIL.n181 VTAIL.n180 185
R125 VTAIL.n176 VTAIL.n175 185
R126 VTAIL.n147 VTAIL.n146 185
R127 VTAIL.n82 VTAIL.n81 185
R128 VTAIL.n141 VTAIL.n140 185
R129 VTAIL.n139 VTAIL.n138 185
R130 VTAIL.n86 VTAIL.n85 185
R131 VTAIL.n133 VTAIL.n132 185
R132 VTAIL.n131 VTAIL.n130 185
R133 VTAIL.n90 VTAIL.n89 185
R134 VTAIL.n125 VTAIL.n124 185
R135 VTAIL.n123 VTAIL.n122 185
R136 VTAIL.n94 VTAIL.n93 185
R137 VTAIL.n117 VTAIL.n116 185
R138 VTAIL.n115 VTAIL.n114 185
R139 VTAIL.n98 VTAIL.n97 185
R140 VTAIL.n109 VTAIL.n108 185
R141 VTAIL.n107 VTAIL.n106 185
R142 VTAIL.n102 VTAIL.n101 185
R143 VTAIL.n247 VTAIL.t6 147.659
R144 VTAIL.n25 VTAIL.t18 147.659
R145 VTAIL.n177 VTAIL.t16 147.659
R146 VTAIL.n103 VTAIL.t3 147.659
R147 VTAIL.n251 VTAIL.n245 104.615
R148 VTAIL.n252 VTAIL.n251 104.615
R149 VTAIL.n252 VTAIL.n241 104.615
R150 VTAIL.n259 VTAIL.n241 104.615
R151 VTAIL.n260 VTAIL.n259 104.615
R152 VTAIL.n260 VTAIL.n237 104.615
R153 VTAIL.n267 VTAIL.n237 104.615
R154 VTAIL.n268 VTAIL.n267 104.615
R155 VTAIL.n268 VTAIL.n233 104.615
R156 VTAIL.n275 VTAIL.n233 104.615
R157 VTAIL.n276 VTAIL.n275 104.615
R158 VTAIL.n276 VTAIL.n229 104.615
R159 VTAIL.n283 VTAIL.n229 104.615
R160 VTAIL.n284 VTAIL.n283 104.615
R161 VTAIL.n284 VTAIL.n225 104.615
R162 VTAIL.n291 VTAIL.n225 104.615
R163 VTAIL.n29 VTAIL.n23 104.615
R164 VTAIL.n30 VTAIL.n29 104.615
R165 VTAIL.n30 VTAIL.n19 104.615
R166 VTAIL.n37 VTAIL.n19 104.615
R167 VTAIL.n38 VTAIL.n37 104.615
R168 VTAIL.n38 VTAIL.n15 104.615
R169 VTAIL.n45 VTAIL.n15 104.615
R170 VTAIL.n46 VTAIL.n45 104.615
R171 VTAIL.n46 VTAIL.n11 104.615
R172 VTAIL.n53 VTAIL.n11 104.615
R173 VTAIL.n54 VTAIL.n53 104.615
R174 VTAIL.n54 VTAIL.n7 104.615
R175 VTAIL.n61 VTAIL.n7 104.615
R176 VTAIL.n62 VTAIL.n61 104.615
R177 VTAIL.n62 VTAIL.n3 104.615
R178 VTAIL.n69 VTAIL.n3 104.615
R179 VTAIL.n221 VTAIL.n155 104.615
R180 VTAIL.n214 VTAIL.n155 104.615
R181 VTAIL.n214 VTAIL.n213 104.615
R182 VTAIL.n213 VTAIL.n159 104.615
R183 VTAIL.n206 VTAIL.n159 104.615
R184 VTAIL.n206 VTAIL.n205 104.615
R185 VTAIL.n205 VTAIL.n163 104.615
R186 VTAIL.n198 VTAIL.n163 104.615
R187 VTAIL.n198 VTAIL.n197 104.615
R188 VTAIL.n197 VTAIL.n167 104.615
R189 VTAIL.n190 VTAIL.n167 104.615
R190 VTAIL.n190 VTAIL.n189 104.615
R191 VTAIL.n189 VTAIL.n171 104.615
R192 VTAIL.n182 VTAIL.n171 104.615
R193 VTAIL.n182 VTAIL.n181 104.615
R194 VTAIL.n181 VTAIL.n175 104.615
R195 VTAIL.n147 VTAIL.n81 104.615
R196 VTAIL.n140 VTAIL.n81 104.615
R197 VTAIL.n140 VTAIL.n139 104.615
R198 VTAIL.n139 VTAIL.n85 104.615
R199 VTAIL.n132 VTAIL.n85 104.615
R200 VTAIL.n132 VTAIL.n131 104.615
R201 VTAIL.n131 VTAIL.n89 104.615
R202 VTAIL.n124 VTAIL.n89 104.615
R203 VTAIL.n124 VTAIL.n123 104.615
R204 VTAIL.n123 VTAIL.n93 104.615
R205 VTAIL.n116 VTAIL.n93 104.615
R206 VTAIL.n116 VTAIL.n115 104.615
R207 VTAIL.n115 VTAIL.n97 104.615
R208 VTAIL.n108 VTAIL.n97 104.615
R209 VTAIL.n108 VTAIL.n107 104.615
R210 VTAIL.n107 VTAIL.n101 104.615
R211 VTAIL.t6 VTAIL.n245 52.3082
R212 VTAIL.t18 VTAIL.n23 52.3082
R213 VTAIL.t16 VTAIL.n175 52.3082
R214 VTAIL.t3 VTAIL.n101 52.3082
R215 VTAIL.n153 VTAIL.n152 48.0206
R216 VTAIL.n151 VTAIL.n150 48.0206
R217 VTAIL.n79 VTAIL.n78 48.0206
R218 VTAIL.n77 VTAIL.n76 48.0206
R219 VTAIL.n295 VTAIL.n294 48.0196
R220 VTAIL.n1 VTAIL.n0 48.0196
R221 VTAIL.n73 VTAIL.n72 48.0196
R222 VTAIL.n75 VTAIL.n74 48.0196
R223 VTAIL.n293 VTAIL.n292 35.2884
R224 VTAIL.n71 VTAIL.n70 35.2884
R225 VTAIL.n223 VTAIL.n222 35.2884
R226 VTAIL.n149 VTAIL.n148 35.2884
R227 VTAIL.n77 VTAIL.n75 25.4876
R228 VTAIL.n293 VTAIL.n223 24.3841
R229 VTAIL.n247 VTAIL.n246 15.6677
R230 VTAIL.n25 VTAIL.n24 15.6677
R231 VTAIL.n177 VTAIL.n176 15.6677
R232 VTAIL.n103 VTAIL.n102 15.6677
R233 VTAIL.n250 VTAIL.n249 12.8005
R234 VTAIL.n290 VTAIL.n224 12.8005
R235 VTAIL.n28 VTAIL.n27 12.8005
R236 VTAIL.n68 VTAIL.n2 12.8005
R237 VTAIL.n220 VTAIL.n154 12.8005
R238 VTAIL.n180 VTAIL.n179 12.8005
R239 VTAIL.n146 VTAIL.n80 12.8005
R240 VTAIL.n106 VTAIL.n105 12.8005
R241 VTAIL.n253 VTAIL.n244 12.0247
R242 VTAIL.n289 VTAIL.n226 12.0247
R243 VTAIL.n31 VTAIL.n22 12.0247
R244 VTAIL.n67 VTAIL.n4 12.0247
R245 VTAIL.n219 VTAIL.n156 12.0247
R246 VTAIL.n183 VTAIL.n174 12.0247
R247 VTAIL.n145 VTAIL.n82 12.0247
R248 VTAIL.n109 VTAIL.n100 12.0247
R249 VTAIL.n254 VTAIL.n242 11.249
R250 VTAIL.n286 VTAIL.n285 11.249
R251 VTAIL.n32 VTAIL.n20 11.249
R252 VTAIL.n64 VTAIL.n63 11.249
R253 VTAIL.n216 VTAIL.n215 11.249
R254 VTAIL.n184 VTAIL.n172 11.249
R255 VTAIL.n142 VTAIL.n141 11.249
R256 VTAIL.n110 VTAIL.n98 11.249
R257 VTAIL.n258 VTAIL.n257 10.4732
R258 VTAIL.n282 VTAIL.n228 10.4732
R259 VTAIL.n36 VTAIL.n35 10.4732
R260 VTAIL.n60 VTAIL.n6 10.4732
R261 VTAIL.n212 VTAIL.n158 10.4732
R262 VTAIL.n188 VTAIL.n187 10.4732
R263 VTAIL.n138 VTAIL.n84 10.4732
R264 VTAIL.n114 VTAIL.n113 10.4732
R265 VTAIL.n261 VTAIL.n240 9.69747
R266 VTAIL.n281 VTAIL.n230 9.69747
R267 VTAIL.n39 VTAIL.n18 9.69747
R268 VTAIL.n59 VTAIL.n8 9.69747
R269 VTAIL.n211 VTAIL.n160 9.69747
R270 VTAIL.n191 VTAIL.n170 9.69747
R271 VTAIL.n137 VTAIL.n86 9.69747
R272 VTAIL.n117 VTAIL.n96 9.69747
R273 VTAIL.n288 VTAIL.n224 9.45567
R274 VTAIL.n66 VTAIL.n2 9.45567
R275 VTAIL.n218 VTAIL.n154 9.45567
R276 VTAIL.n144 VTAIL.n80 9.45567
R277 VTAIL.n271 VTAIL.n270 9.3005
R278 VTAIL.n273 VTAIL.n272 9.3005
R279 VTAIL.n232 VTAIL.n231 9.3005
R280 VTAIL.n279 VTAIL.n278 9.3005
R281 VTAIL.n281 VTAIL.n280 9.3005
R282 VTAIL.n228 VTAIL.n227 9.3005
R283 VTAIL.n287 VTAIL.n286 9.3005
R284 VTAIL.n289 VTAIL.n288 9.3005
R285 VTAIL.n265 VTAIL.n264 9.3005
R286 VTAIL.n263 VTAIL.n262 9.3005
R287 VTAIL.n240 VTAIL.n239 9.3005
R288 VTAIL.n257 VTAIL.n256 9.3005
R289 VTAIL.n255 VTAIL.n254 9.3005
R290 VTAIL.n244 VTAIL.n243 9.3005
R291 VTAIL.n249 VTAIL.n248 9.3005
R292 VTAIL.n236 VTAIL.n235 9.3005
R293 VTAIL.n49 VTAIL.n48 9.3005
R294 VTAIL.n51 VTAIL.n50 9.3005
R295 VTAIL.n10 VTAIL.n9 9.3005
R296 VTAIL.n57 VTAIL.n56 9.3005
R297 VTAIL.n59 VTAIL.n58 9.3005
R298 VTAIL.n6 VTAIL.n5 9.3005
R299 VTAIL.n65 VTAIL.n64 9.3005
R300 VTAIL.n67 VTAIL.n66 9.3005
R301 VTAIL.n43 VTAIL.n42 9.3005
R302 VTAIL.n41 VTAIL.n40 9.3005
R303 VTAIL.n18 VTAIL.n17 9.3005
R304 VTAIL.n35 VTAIL.n34 9.3005
R305 VTAIL.n33 VTAIL.n32 9.3005
R306 VTAIL.n22 VTAIL.n21 9.3005
R307 VTAIL.n27 VTAIL.n26 9.3005
R308 VTAIL.n14 VTAIL.n13 9.3005
R309 VTAIL.n219 VTAIL.n218 9.3005
R310 VTAIL.n217 VTAIL.n216 9.3005
R311 VTAIL.n158 VTAIL.n157 9.3005
R312 VTAIL.n211 VTAIL.n210 9.3005
R313 VTAIL.n209 VTAIL.n208 9.3005
R314 VTAIL.n162 VTAIL.n161 9.3005
R315 VTAIL.n203 VTAIL.n202 9.3005
R316 VTAIL.n201 VTAIL.n200 9.3005
R317 VTAIL.n166 VTAIL.n165 9.3005
R318 VTAIL.n195 VTAIL.n194 9.3005
R319 VTAIL.n193 VTAIL.n192 9.3005
R320 VTAIL.n170 VTAIL.n169 9.3005
R321 VTAIL.n187 VTAIL.n186 9.3005
R322 VTAIL.n185 VTAIL.n184 9.3005
R323 VTAIL.n174 VTAIL.n173 9.3005
R324 VTAIL.n179 VTAIL.n178 9.3005
R325 VTAIL.n129 VTAIL.n128 9.3005
R326 VTAIL.n88 VTAIL.n87 9.3005
R327 VTAIL.n135 VTAIL.n134 9.3005
R328 VTAIL.n137 VTAIL.n136 9.3005
R329 VTAIL.n84 VTAIL.n83 9.3005
R330 VTAIL.n143 VTAIL.n142 9.3005
R331 VTAIL.n145 VTAIL.n144 9.3005
R332 VTAIL.n127 VTAIL.n126 9.3005
R333 VTAIL.n92 VTAIL.n91 9.3005
R334 VTAIL.n121 VTAIL.n120 9.3005
R335 VTAIL.n119 VTAIL.n118 9.3005
R336 VTAIL.n96 VTAIL.n95 9.3005
R337 VTAIL.n113 VTAIL.n112 9.3005
R338 VTAIL.n111 VTAIL.n110 9.3005
R339 VTAIL.n100 VTAIL.n99 9.3005
R340 VTAIL.n105 VTAIL.n104 9.3005
R341 VTAIL.n262 VTAIL.n238 8.92171
R342 VTAIL.n278 VTAIL.n277 8.92171
R343 VTAIL.n40 VTAIL.n16 8.92171
R344 VTAIL.n56 VTAIL.n55 8.92171
R345 VTAIL.n208 VTAIL.n207 8.92171
R346 VTAIL.n192 VTAIL.n168 8.92171
R347 VTAIL.n134 VTAIL.n133 8.92171
R348 VTAIL.n118 VTAIL.n94 8.92171
R349 VTAIL.n266 VTAIL.n265 8.14595
R350 VTAIL.n274 VTAIL.n232 8.14595
R351 VTAIL.n44 VTAIL.n43 8.14595
R352 VTAIL.n52 VTAIL.n10 8.14595
R353 VTAIL.n204 VTAIL.n162 8.14595
R354 VTAIL.n196 VTAIL.n195 8.14595
R355 VTAIL.n130 VTAIL.n88 8.14595
R356 VTAIL.n122 VTAIL.n121 8.14595
R357 VTAIL.n269 VTAIL.n236 7.3702
R358 VTAIL.n273 VTAIL.n234 7.3702
R359 VTAIL.n47 VTAIL.n14 7.3702
R360 VTAIL.n51 VTAIL.n12 7.3702
R361 VTAIL.n203 VTAIL.n164 7.3702
R362 VTAIL.n199 VTAIL.n166 7.3702
R363 VTAIL.n129 VTAIL.n90 7.3702
R364 VTAIL.n125 VTAIL.n92 7.3702
R365 VTAIL.n270 VTAIL.n269 6.59444
R366 VTAIL.n270 VTAIL.n234 6.59444
R367 VTAIL.n48 VTAIL.n47 6.59444
R368 VTAIL.n48 VTAIL.n12 6.59444
R369 VTAIL.n200 VTAIL.n164 6.59444
R370 VTAIL.n200 VTAIL.n199 6.59444
R371 VTAIL.n126 VTAIL.n90 6.59444
R372 VTAIL.n126 VTAIL.n125 6.59444
R373 VTAIL.n266 VTAIL.n236 5.81868
R374 VTAIL.n274 VTAIL.n273 5.81868
R375 VTAIL.n44 VTAIL.n14 5.81868
R376 VTAIL.n52 VTAIL.n51 5.81868
R377 VTAIL.n204 VTAIL.n203 5.81868
R378 VTAIL.n196 VTAIL.n166 5.81868
R379 VTAIL.n130 VTAIL.n129 5.81868
R380 VTAIL.n122 VTAIL.n92 5.81868
R381 VTAIL.n265 VTAIL.n238 5.04292
R382 VTAIL.n277 VTAIL.n232 5.04292
R383 VTAIL.n43 VTAIL.n16 5.04292
R384 VTAIL.n55 VTAIL.n10 5.04292
R385 VTAIL.n207 VTAIL.n162 5.04292
R386 VTAIL.n195 VTAIL.n168 5.04292
R387 VTAIL.n133 VTAIL.n88 5.04292
R388 VTAIL.n121 VTAIL.n94 5.04292
R389 VTAIL.n248 VTAIL.n247 4.38563
R390 VTAIL.n26 VTAIL.n25 4.38563
R391 VTAIL.n178 VTAIL.n177 4.38563
R392 VTAIL.n104 VTAIL.n103 4.38563
R393 VTAIL.n262 VTAIL.n261 4.26717
R394 VTAIL.n278 VTAIL.n230 4.26717
R395 VTAIL.n40 VTAIL.n39 4.26717
R396 VTAIL.n56 VTAIL.n8 4.26717
R397 VTAIL.n208 VTAIL.n160 4.26717
R398 VTAIL.n192 VTAIL.n191 4.26717
R399 VTAIL.n134 VTAIL.n86 4.26717
R400 VTAIL.n118 VTAIL.n117 4.26717
R401 VTAIL.n258 VTAIL.n240 3.49141
R402 VTAIL.n282 VTAIL.n281 3.49141
R403 VTAIL.n36 VTAIL.n18 3.49141
R404 VTAIL.n60 VTAIL.n59 3.49141
R405 VTAIL.n212 VTAIL.n211 3.49141
R406 VTAIL.n188 VTAIL.n170 3.49141
R407 VTAIL.n138 VTAIL.n137 3.49141
R408 VTAIL.n114 VTAIL.n96 3.49141
R409 VTAIL.n257 VTAIL.n242 2.71565
R410 VTAIL.n285 VTAIL.n228 2.71565
R411 VTAIL.n35 VTAIL.n20 2.71565
R412 VTAIL.n63 VTAIL.n6 2.71565
R413 VTAIL.n215 VTAIL.n158 2.71565
R414 VTAIL.n187 VTAIL.n172 2.71565
R415 VTAIL.n141 VTAIL.n84 2.71565
R416 VTAIL.n113 VTAIL.n98 2.71565
R417 VTAIL.n254 VTAIL.n253 1.93989
R418 VTAIL.n286 VTAIL.n226 1.93989
R419 VTAIL.n32 VTAIL.n31 1.93989
R420 VTAIL.n64 VTAIL.n4 1.93989
R421 VTAIL.n216 VTAIL.n156 1.93989
R422 VTAIL.n184 VTAIL.n183 1.93989
R423 VTAIL.n142 VTAIL.n82 1.93989
R424 VTAIL.n110 VTAIL.n109 1.93989
R425 VTAIL.n294 VTAIL.t8 1.56448
R426 VTAIL.n294 VTAIL.t1 1.56448
R427 VTAIL.n0 VTAIL.t7 1.56448
R428 VTAIL.n0 VTAIL.t5 1.56448
R429 VTAIL.n72 VTAIL.t12 1.56448
R430 VTAIL.n72 VTAIL.t15 1.56448
R431 VTAIL.n74 VTAIL.t9 1.56448
R432 VTAIL.n74 VTAIL.t11 1.56448
R433 VTAIL.n152 VTAIL.t10 1.56448
R434 VTAIL.n152 VTAIL.t14 1.56448
R435 VTAIL.n150 VTAIL.t13 1.56448
R436 VTAIL.n150 VTAIL.t17 1.56448
R437 VTAIL.n78 VTAIL.t4 1.56448
R438 VTAIL.n78 VTAIL.t2 1.56448
R439 VTAIL.n76 VTAIL.t0 1.56448
R440 VTAIL.n76 VTAIL.t19 1.56448
R441 VTAIL.n250 VTAIL.n244 1.16414
R442 VTAIL.n290 VTAIL.n289 1.16414
R443 VTAIL.n28 VTAIL.n22 1.16414
R444 VTAIL.n68 VTAIL.n67 1.16414
R445 VTAIL.n220 VTAIL.n219 1.16414
R446 VTAIL.n180 VTAIL.n174 1.16414
R447 VTAIL.n146 VTAIL.n145 1.16414
R448 VTAIL.n106 VTAIL.n100 1.16414
R449 VTAIL.n79 VTAIL.n77 1.10395
R450 VTAIL.n149 VTAIL.n79 1.10395
R451 VTAIL.n153 VTAIL.n151 1.10395
R452 VTAIL.n223 VTAIL.n153 1.10395
R453 VTAIL.n75 VTAIL.n73 1.10395
R454 VTAIL.n73 VTAIL.n71 1.10395
R455 VTAIL.n295 VTAIL.n293 1.10395
R456 VTAIL.n151 VTAIL.n149 1.02205
R457 VTAIL.n71 VTAIL.n1 1.02205
R458 VTAIL VTAIL.n1 0.886276
R459 VTAIL.n249 VTAIL.n246 0.388379
R460 VTAIL.n292 VTAIL.n224 0.388379
R461 VTAIL.n27 VTAIL.n24 0.388379
R462 VTAIL.n70 VTAIL.n2 0.388379
R463 VTAIL.n222 VTAIL.n154 0.388379
R464 VTAIL.n179 VTAIL.n176 0.388379
R465 VTAIL.n148 VTAIL.n80 0.388379
R466 VTAIL.n105 VTAIL.n102 0.388379
R467 VTAIL VTAIL.n295 0.218172
R468 VTAIL.n248 VTAIL.n243 0.155672
R469 VTAIL.n255 VTAIL.n243 0.155672
R470 VTAIL.n256 VTAIL.n255 0.155672
R471 VTAIL.n256 VTAIL.n239 0.155672
R472 VTAIL.n263 VTAIL.n239 0.155672
R473 VTAIL.n264 VTAIL.n263 0.155672
R474 VTAIL.n264 VTAIL.n235 0.155672
R475 VTAIL.n271 VTAIL.n235 0.155672
R476 VTAIL.n272 VTAIL.n271 0.155672
R477 VTAIL.n272 VTAIL.n231 0.155672
R478 VTAIL.n279 VTAIL.n231 0.155672
R479 VTAIL.n280 VTAIL.n279 0.155672
R480 VTAIL.n280 VTAIL.n227 0.155672
R481 VTAIL.n287 VTAIL.n227 0.155672
R482 VTAIL.n288 VTAIL.n287 0.155672
R483 VTAIL.n26 VTAIL.n21 0.155672
R484 VTAIL.n33 VTAIL.n21 0.155672
R485 VTAIL.n34 VTAIL.n33 0.155672
R486 VTAIL.n34 VTAIL.n17 0.155672
R487 VTAIL.n41 VTAIL.n17 0.155672
R488 VTAIL.n42 VTAIL.n41 0.155672
R489 VTAIL.n42 VTAIL.n13 0.155672
R490 VTAIL.n49 VTAIL.n13 0.155672
R491 VTAIL.n50 VTAIL.n49 0.155672
R492 VTAIL.n50 VTAIL.n9 0.155672
R493 VTAIL.n57 VTAIL.n9 0.155672
R494 VTAIL.n58 VTAIL.n57 0.155672
R495 VTAIL.n58 VTAIL.n5 0.155672
R496 VTAIL.n65 VTAIL.n5 0.155672
R497 VTAIL.n66 VTAIL.n65 0.155672
R498 VTAIL.n218 VTAIL.n217 0.155672
R499 VTAIL.n217 VTAIL.n157 0.155672
R500 VTAIL.n210 VTAIL.n157 0.155672
R501 VTAIL.n210 VTAIL.n209 0.155672
R502 VTAIL.n209 VTAIL.n161 0.155672
R503 VTAIL.n202 VTAIL.n161 0.155672
R504 VTAIL.n202 VTAIL.n201 0.155672
R505 VTAIL.n201 VTAIL.n165 0.155672
R506 VTAIL.n194 VTAIL.n165 0.155672
R507 VTAIL.n194 VTAIL.n193 0.155672
R508 VTAIL.n193 VTAIL.n169 0.155672
R509 VTAIL.n186 VTAIL.n169 0.155672
R510 VTAIL.n186 VTAIL.n185 0.155672
R511 VTAIL.n185 VTAIL.n173 0.155672
R512 VTAIL.n178 VTAIL.n173 0.155672
R513 VTAIL.n144 VTAIL.n143 0.155672
R514 VTAIL.n143 VTAIL.n83 0.155672
R515 VTAIL.n136 VTAIL.n83 0.155672
R516 VTAIL.n136 VTAIL.n135 0.155672
R517 VTAIL.n135 VTAIL.n87 0.155672
R518 VTAIL.n128 VTAIL.n87 0.155672
R519 VTAIL.n128 VTAIL.n127 0.155672
R520 VTAIL.n127 VTAIL.n91 0.155672
R521 VTAIL.n120 VTAIL.n91 0.155672
R522 VTAIL.n120 VTAIL.n119 0.155672
R523 VTAIL.n119 VTAIL.n95 0.155672
R524 VTAIL.n112 VTAIL.n95 0.155672
R525 VTAIL.n112 VTAIL.n111 0.155672
R526 VTAIL.n111 VTAIL.n99 0.155672
R527 VTAIL.n104 VTAIL.n99 0.155672
R528 VDD1.n68 VDD1.n67 289.615
R529 VDD1.n139 VDD1.n138 289.615
R530 VDD1.n67 VDD1.n66 185
R531 VDD1.n2 VDD1.n1 185
R532 VDD1.n61 VDD1.n60 185
R533 VDD1.n59 VDD1.n58 185
R534 VDD1.n6 VDD1.n5 185
R535 VDD1.n53 VDD1.n52 185
R536 VDD1.n51 VDD1.n50 185
R537 VDD1.n10 VDD1.n9 185
R538 VDD1.n45 VDD1.n44 185
R539 VDD1.n43 VDD1.n42 185
R540 VDD1.n14 VDD1.n13 185
R541 VDD1.n37 VDD1.n36 185
R542 VDD1.n35 VDD1.n34 185
R543 VDD1.n18 VDD1.n17 185
R544 VDD1.n29 VDD1.n28 185
R545 VDD1.n27 VDD1.n26 185
R546 VDD1.n22 VDD1.n21 185
R547 VDD1.n93 VDD1.n92 185
R548 VDD1.n98 VDD1.n97 185
R549 VDD1.n100 VDD1.n99 185
R550 VDD1.n89 VDD1.n88 185
R551 VDD1.n106 VDD1.n105 185
R552 VDD1.n108 VDD1.n107 185
R553 VDD1.n85 VDD1.n84 185
R554 VDD1.n114 VDD1.n113 185
R555 VDD1.n116 VDD1.n115 185
R556 VDD1.n81 VDD1.n80 185
R557 VDD1.n122 VDD1.n121 185
R558 VDD1.n124 VDD1.n123 185
R559 VDD1.n77 VDD1.n76 185
R560 VDD1.n130 VDD1.n129 185
R561 VDD1.n132 VDD1.n131 185
R562 VDD1.n73 VDD1.n72 185
R563 VDD1.n138 VDD1.n137 185
R564 VDD1.n94 VDD1.t6 147.659
R565 VDD1.n23 VDD1.t8 147.659
R566 VDD1.n67 VDD1.n1 104.615
R567 VDD1.n60 VDD1.n1 104.615
R568 VDD1.n60 VDD1.n59 104.615
R569 VDD1.n59 VDD1.n5 104.615
R570 VDD1.n52 VDD1.n5 104.615
R571 VDD1.n52 VDD1.n51 104.615
R572 VDD1.n51 VDD1.n9 104.615
R573 VDD1.n44 VDD1.n9 104.615
R574 VDD1.n44 VDD1.n43 104.615
R575 VDD1.n43 VDD1.n13 104.615
R576 VDD1.n36 VDD1.n13 104.615
R577 VDD1.n36 VDD1.n35 104.615
R578 VDD1.n35 VDD1.n17 104.615
R579 VDD1.n28 VDD1.n17 104.615
R580 VDD1.n28 VDD1.n27 104.615
R581 VDD1.n27 VDD1.n21 104.615
R582 VDD1.n98 VDD1.n92 104.615
R583 VDD1.n99 VDD1.n98 104.615
R584 VDD1.n99 VDD1.n88 104.615
R585 VDD1.n106 VDD1.n88 104.615
R586 VDD1.n107 VDD1.n106 104.615
R587 VDD1.n107 VDD1.n84 104.615
R588 VDD1.n114 VDD1.n84 104.615
R589 VDD1.n115 VDD1.n114 104.615
R590 VDD1.n115 VDD1.n80 104.615
R591 VDD1.n122 VDD1.n80 104.615
R592 VDD1.n123 VDD1.n122 104.615
R593 VDD1.n123 VDD1.n76 104.615
R594 VDD1.n130 VDD1.n76 104.615
R595 VDD1.n131 VDD1.n130 104.615
R596 VDD1.n131 VDD1.n72 104.615
R597 VDD1.n138 VDD1.n72 104.615
R598 VDD1.n143 VDD1.n142 65.4706
R599 VDD1.n70 VDD1.n69 64.6993
R600 VDD1.n141 VDD1.n140 64.6983
R601 VDD1.n145 VDD1.n144 64.6983
R602 VDD1.n70 VDD1.n68 53.0706
R603 VDD1.n141 VDD1.n139 53.0706
R604 VDD1.t8 VDD1.n21 52.3082
R605 VDD1.t6 VDD1.n92 52.3082
R606 VDD1.n145 VDD1.n143 41.0052
R607 VDD1.n23 VDD1.n22 15.6677
R608 VDD1.n94 VDD1.n93 15.6677
R609 VDD1.n66 VDD1.n0 12.8005
R610 VDD1.n26 VDD1.n25 12.8005
R611 VDD1.n97 VDD1.n96 12.8005
R612 VDD1.n137 VDD1.n71 12.8005
R613 VDD1.n65 VDD1.n2 12.0247
R614 VDD1.n29 VDD1.n20 12.0247
R615 VDD1.n100 VDD1.n91 12.0247
R616 VDD1.n136 VDD1.n73 12.0247
R617 VDD1.n62 VDD1.n61 11.249
R618 VDD1.n30 VDD1.n18 11.249
R619 VDD1.n101 VDD1.n89 11.249
R620 VDD1.n133 VDD1.n132 11.249
R621 VDD1.n58 VDD1.n4 10.4732
R622 VDD1.n34 VDD1.n33 10.4732
R623 VDD1.n105 VDD1.n104 10.4732
R624 VDD1.n129 VDD1.n75 10.4732
R625 VDD1.n57 VDD1.n6 9.69747
R626 VDD1.n37 VDD1.n16 9.69747
R627 VDD1.n108 VDD1.n87 9.69747
R628 VDD1.n128 VDD1.n77 9.69747
R629 VDD1.n64 VDD1.n0 9.45567
R630 VDD1.n135 VDD1.n71 9.45567
R631 VDD1.n49 VDD1.n48 9.3005
R632 VDD1.n8 VDD1.n7 9.3005
R633 VDD1.n55 VDD1.n54 9.3005
R634 VDD1.n57 VDD1.n56 9.3005
R635 VDD1.n4 VDD1.n3 9.3005
R636 VDD1.n63 VDD1.n62 9.3005
R637 VDD1.n65 VDD1.n64 9.3005
R638 VDD1.n47 VDD1.n46 9.3005
R639 VDD1.n12 VDD1.n11 9.3005
R640 VDD1.n41 VDD1.n40 9.3005
R641 VDD1.n39 VDD1.n38 9.3005
R642 VDD1.n16 VDD1.n15 9.3005
R643 VDD1.n33 VDD1.n32 9.3005
R644 VDD1.n31 VDD1.n30 9.3005
R645 VDD1.n20 VDD1.n19 9.3005
R646 VDD1.n25 VDD1.n24 9.3005
R647 VDD1.n118 VDD1.n117 9.3005
R648 VDD1.n120 VDD1.n119 9.3005
R649 VDD1.n79 VDD1.n78 9.3005
R650 VDD1.n126 VDD1.n125 9.3005
R651 VDD1.n128 VDD1.n127 9.3005
R652 VDD1.n75 VDD1.n74 9.3005
R653 VDD1.n134 VDD1.n133 9.3005
R654 VDD1.n136 VDD1.n135 9.3005
R655 VDD1.n112 VDD1.n111 9.3005
R656 VDD1.n110 VDD1.n109 9.3005
R657 VDD1.n87 VDD1.n86 9.3005
R658 VDD1.n104 VDD1.n103 9.3005
R659 VDD1.n102 VDD1.n101 9.3005
R660 VDD1.n91 VDD1.n90 9.3005
R661 VDD1.n96 VDD1.n95 9.3005
R662 VDD1.n83 VDD1.n82 9.3005
R663 VDD1.n54 VDD1.n53 8.92171
R664 VDD1.n38 VDD1.n14 8.92171
R665 VDD1.n109 VDD1.n85 8.92171
R666 VDD1.n125 VDD1.n124 8.92171
R667 VDD1.n50 VDD1.n8 8.14595
R668 VDD1.n42 VDD1.n41 8.14595
R669 VDD1.n113 VDD1.n112 8.14595
R670 VDD1.n121 VDD1.n79 8.14595
R671 VDD1.n49 VDD1.n10 7.3702
R672 VDD1.n45 VDD1.n12 7.3702
R673 VDD1.n116 VDD1.n83 7.3702
R674 VDD1.n120 VDD1.n81 7.3702
R675 VDD1.n46 VDD1.n10 6.59444
R676 VDD1.n46 VDD1.n45 6.59444
R677 VDD1.n117 VDD1.n116 6.59444
R678 VDD1.n117 VDD1.n81 6.59444
R679 VDD1.n50 VDD1.n49 5.81868
R680 VDD1.n42 VDD1.n12 5.81868
R681 VDD1.n113 VDD1.n83 5.81868
R682 VDD1.n121 VDD1.n120 5.81868
R683 VDD1.n53 VDD1.n8 5.04292
R684 VDD1.n41 VDD1.n14 5.04292
R685 VDD1.n112 VDD1.n85 5.04292
R686 VDD1.n124 VDD1.n79 5.04292
R687 VDD1.n95 VDD1.n94 4.38563
R688 VDD1.n24 VDD1.n23 4.38563
R689 VDD1.n54 VDD1.n6 4.26717
R690 VDD1.n38 VDD1.n37 4.26717
R691 VDD1.n109 VDD1.n108 4.26717
R692 VDD1.n125 VDD1.n77 4.26717
R693 VDD1.n58 VDD1.n57 3.49141
R694 VDD1.n34 VDD1.n16 3.49141
R695 VDD1.n105 VDD1.n87 3.49141
R696 VDD1.n129 VDD1.n128 3.49141
R697 VDD1.n61 VDD1.n4 2.71565
R698 VDD1.n33 VDD1.n18 2.71565
R699 VDD1.n104 VDD1.n89 2.71565
R700 VDD1.n132 VDD1.n75 2.71565
R701 VDD1.n62 VDD1.n2 1.93989
R702 VDD1.n30 VDD1.n29 1.93989
R703 VDD1.n101 VDD1.n100 1.93989
R704 VDD1.n133 VDD1.n73 1.93989
R705 VDD1.n144 VDD1.t1 1.56448
R706 VDD1.n144 VDD1.t7 1.56448
R707 VDD1.n69 VDD1.t5 1.56448
R708 VDD1.n69 VDD1.t3 1.56448
R709 VDD1.n142 VDD1.t0 1.56448
R710 VDD1.n142 VDD1.t9 1.56448
R711 VDD1.n140 VDD1.t4 1.56448
R712 VDD1.n140 VDD1.t2 1.56448
R713 VDD1.n66 VDD1.n65 1.16414
R714 VDD1.n26 VDD1.n20 1.16414
R715 VDD1.n97 VDD1.n91 1.16414
R716 VDD1.n137 VDD1.n136 1.16414
R717 VDD1 VDD1.n145 0.769897
R718 VDD1.n68 VDD1.n0 0.388379
R719 VDD1.n25 VDD1.n22 0.388379
R720 VDD1.n96 VDD1.n93 0.388379
R721 VDD1.n139 VDD1.n71 0.388379
R722 VDD1 VDD1.n70 0.334552
R723 VDD1.n143 VDD1.n141 0.221016
R724 VDD1.n64 VDD1.n63 0.155672
R725 VDD1.n63 VDD1.n3 0.155672
R726 VDD1.n56 VDD1.n3 0.155672
R727 VDD1.n56 VDD1.n55 0.155672
R728 VDD1.n55 VDD1.n7 0.155672
R729 VDD1.n48 VDD1.n7 0.155672
R730 VDD1.n48 VDD1.n47 0.155672
R731 VDD1.n47 VDD1.n11 0.155672
R732 VDD1.n40 VDD1.n11 0.155672
R733 VDD1.n40 VDD1.n39 0.155672
R734 VDD1.n39 VDD1.n15 0.155672
R735 VDD1.n32 VDD1.n15 0.155672
R736 VDD1.n32 VDD1.n31 0.155672
R737 VDD1.n31 VDD1.n19 0.155672
R738 VDD1.n24 VDD1.n19 0.155672
R739 VDD1.n95 VDD1.n90 0.155672
R740 VDD1.n102 VDD1.n90 0.155672
R741 VDD1.n103 VDD1.n102 0.155672
R742 VDD1.n103 VDD1.n86 0.155672
R743 VDD1.n110 VDD1.n86 0.155672
R744 VDD1.n111 VDD1.n110 0.155672
R745 VDD1.n111 VDD1.n82 0.155672
R746 VDD1.n118 VDD1.n82 0.155672
R747 VDD1.n119 VDD1.n118 0.155672
R748 VDD1.n119 VDD1.n78 0.155672
R749 VDD1.n126 VDD1.n78 0.155672
R750 VDD1.n127 VDD1.n126 0.155672
R751 VDD1.n127 VDD1.n74 0.155672
R752 VDD1.n134 VDD1.n74 0.155672
R753 VDD1.n135 VDD1.n134 0.155672
R754 B.n548 B.n111 585
R755 B.n111 B.n58 585
R756 B.n550 B.n549 585
R757 B.n552 B.n110 585
R758 B.n555 B.n554 585
R759 B.n556 B.n109 585
R760 B.n558 B.n557 585
R761 B.n560 B.n108 585
R762 B.n563 B.n562 585
R763 B.n564 B.n107 585
R764 B.n566 B.n565 585
R765 B.n568 B.n106 585
R766 B.n571 B.n570 585
R767 B.n572 B.n105 585
R768 B.n574 B.n573 585
R769 B.n576 B.n104 585
R770 B.n579 B.n578 585
R771 B.n580 B.n103 585
R772 B.n582 B.n581 585
R773 B.n584 B.n102 585
R774 B.n587 B.n586 585
R775 B.n588 B.n101 585
R776 B.n590 B.n589 585
R777 B.n592 B.n100 585
R778 B.n595 B.n594 585
R779 B.n596 B.n99 585
R780 B.n598 B.n597 585
R781 B.n600 B.n98 585
R782 B.n603 B.n602 585
R783 B.n604 B.n97 585
R784 B.n606 B.n605 585
R785 B.n608 B.n96 585
R786 B.n611 B.n610 585
R787 B.n612 B.n95 585
R788 B.n614 B.n613 585
R789 B.n616 B.n94 585
R790 B.n619 B.n618 585
R791 B.n620 B.n93 585
R792 B.n622 B.n621 585
R793 B.n624 B.n92 585
R794 B.n627 B.n626 585
R795 B.n628 B.n91 585
R796 B.n630 B.n629 585
R797 B.n632 B.n90 585
R798 B.n635 B.n634 585
R799 B.n637 B.n87 585
R800 B.n639 B.n638 585
R801 B.n641 B.n86 585
R802 B.n644 B.n643 585
R803 B.n645 B.n85 585
R804 B.n647 B.n646 585
R805 B.n649 B.n84 585
R806 B.n652 B.n651 585
R807 B.n653 B.n81 585
R808 B.n656 B.n655 585
R809 B.n658 B.n80 585
R810 B.n661 B.n660 585
R811 B.n662 B.n79 585
R812 B.n664 B.n663 585
R813 B.n666 B.n78 585
R814 B.n669 B.n668 585
R815 B.n670 B.n77 585
R816 B.n672 B.n671 585
R817 B.n674 B.n76 585
R818 B.n677 B.n676 585
R819 B.n678 B.n75 585
R820 B.n680 B.n679 585
R821 B.n682 B.n74 585
R822 B.n685 B.n684 585
R823 B.n686 B.n73 585
R824 B.n688 B.n687 585
R825 B.n690 B.n72 585
R826 B.n693 B.n692 585
R827 B.n694 B.n71 585
R828 B.n696 B.n695 585
R829 B.n698 B.n70 585
R830 B.n701 B.n700 585
R831 B.n702 B.n69 585
R832 B.n704 B.n703 585
R833 B.n706 B.n68 585
R834 B.n709 B.n708 585
R835 B.n710 B.n67 585
R836 B.n712 B.n711 585
R837 B.n714 B.n66 585
R838 B.n717 B.n716 585
R839 B.n718 B.n65 585
R840 B.n720 B.n719 585
R841 B.n722 B.n64 585
R842 B.n725 B.n724 585
R843 B.n726 B.n63 585
R844 B.n728 B.n727 585
R845 B.n730 B.n62 585
R846 B.n733 B.n732 585
R847 B.n734 B.n61 585
R848 B.n736 B.n735 585
R849 B.n738 B.n60 585
R850 B.n741 B.n740 585
R851 B.n742 B.n59 585
R852 B.n547 B.n57 585
R853 B.n745 B.n57 585
R854 B.n546 B.n56 585
R855 B.n746 B.n56 585
R856 B.n545 B.n55 585
R857 B.n747 B.n55 585
R858 B.n544 B.n543 585
R859 B.n543 B.n51 585
R860 B.n542 B.n50 585
R861 B.n753 B.n50 585
R862 B.n541 B.n49 585
R863 B.n754 B.n49 585
R864 B.n540 B.n48 585
R865 B.n755 B.n48 585
R866 B.n539 B.n538 585
R867 B.n538 B.n44 585
R868 B.n537 B.n43 585
R869 B.n761 B.n43 585
R870 B.n536 B.n42 585
R871 B.n762 B.n42 585
R872 B.n535 B.n41 585
R873 B.n763 B.n41 585
R874 B.n534 B.n533 585
R875 B.n533 B.n40 585
R876 B.n532 B.n36 585
R877 B.n769 B.n36 585
R878 B.n531 B.n35 585
R879 B.n770 B.n35 585
R880 B.n530 B.n34 585
R881 B.n771 B.n34 585
R882 B.n529 B.n528 585
R883 B.n528 B.n33 585
R884 B.n527 B.n29 585
R885 B.n777 B.n29 585
R886 B.n526 B.n28 585
R887 B.n778 B.n28 585
R888 B.n525 B.n27 585
R889 B.n779 B.n27 585
R890 B.n524 B.n523 585
R891 B.n523 B.n26 585
R892 B.n522 B.n22 585
R893 B.n785 B.n22 585
R894 B.n521 B.n21 585
R895 B.n786 B.n21 585
R896 B.n520 B.n20 585
R897 B.n787 B.n20 585
R898 B.n519 B.n518 585
R899 B.n518 B.n19 585
R900 B.n517 B.n15 585
R901 B.n793 B.n15 585
R902 B.n516 B.n14 585
R903 B.n794 B.n14 585
R904 B.n515 B.n13 585
R905 B.n795 B.n13 585
R906 B.n514 B.n513 585
R907 B.n513 B.n12 585
R908 B.n512 B.n511 585
R909 B.n512 B.n8 585
R910 B.n510 B.n7 585
R911 B.n802 B.n7 585
R912 B.n509 B.n6 585
R913 B.n803 B.n6 585
R914 B.n508 B.n5 585
R915 B.n804 B.n5 585
R916 B.n507 B.n506 585
R917 B.n506 B.n4 585
R918 B.n505 B.n112 585
R919 B.n505 B.n504 585
R920 B.n494 B.n113 585
R921 B.n497 B.n113 585
R922 B.n496 B.n495 585
R923 B.n498 B.n496 585
R924 B.n493 B.n118 585
R925 B.n118 B.n117 585
R926 B.n492 B.n491 585
R927 B.n491 B.n490 585
R928 B.n120 B.n119 585
R929 B.n483 B.n120 585
R930 B.n482 B.n481 585
R931 B.n484 B.n482 585
R932 B.n480 B.n125 585
R933 B.n125 B.n124 585
R934 B.n479 B.n478 585
R935 B.n478 B.n477 585
R936 B.n127 B.n126 585
R937 B.n470 B.n127 585
R938 B.n469 B.n468 585
R939 B.n471 B.n469 585
R940 B.n467 B.n132 585
R941 B.n132 B.n131 585
R942 B.n466 B.n465 585
R943 B.n465 B.n464 585
R944 B.n134 B.n133 585
R945 B.n457 B.n134 585
R946 B.n456 B.n455 585
R947 B.n458 B.n456 585
R948 B.n454 B.n139 585
R949 B.n139 B.n138 585
R950 B.n453 B.n452 585
R951 B.n452 B.n451 585
R952 B.n141 B.n140 585
R953 B.n444 B.n141 585
R954 B.n443 B.n442 585
R955 B.n445 B.n443 585
R956 B.n441 B.n146 585
R957 B.n146 B.n145 585
R958 B.n440 B.n439 585
R959 B.n439 B.n438 585
R960 B.n148 B.n147 585
R961 B.n149 B.n148 585
R962 B.n431 B.n430 585
R963 B.n432 B.n431 585
R964 B.n429 B.n154 585
R965 B.n154 B.n153 585
R966 B.n428 B.n427 585
R967 B.n427 B.n426 585
R968 B.n156 B.n155 585
R969 B.n157 B.n156 585
R970 B.n419 B.n418 585
R971 B.n420 B.n419 585
R972 B.n417 B.n162 585
R973 B.n162 B.n161 585
R974 B.n416 B.n415 585
R975 B.n415 B.n414 585
R976 B.n411 B.n166 585
R977 B.n410 B.n409 585
R978 B.n407 B.n167 585
R979 B.n407 B.n165 585
R980 B.n406 B.n405 585
R981 B.n404 B.n403 585
R982 B.n402 B.n169 585
R983 B.n400 B.n399 585
R984 B.n398 B.n170 585
R985 B.n397 B.n396 585
R986 B.n394 B.n171 585
R987 B.n392 B.n391 585
R988 B.n390 B.n172 585
R989 B.n389 B.n388 585
R990 B.n386 B.n173 585
R991 B.n384 B.n383 585
R992 B.n382 B.n174 585
R993 B.n381 B.n380 585
R994 B.n378 B.n175 585
R995 B.n376 B.n375 585
R996 B.n374 B.n176 585
R997 B.n373 B.n372 585
R998 B.n370 B.n177 585
R999 B.n368 B.n367 585
R1000 B.n366 B.n178 585
R1001 B.n365 B.n364 585
R1002 B.n362 B.n179 585
R1003 B.n360 B.n359 585
R1004 B.n358 B.n180 585
R1005 B.n357 B.n356 585
R1006 B.n354 B.n181 585
R1007 B.n352 B.n351 585
R1008 B.n350 B.n182 585
R1009 B.n349 B.n348 585
R1010 B.n346 B.n183 585
R1011 B.n344 B.n343 585
R1012 B.n342 B.n184 585
R1013 B.n341 B.n340 585
R1014 B.n338 B.n185 585
R1015 B.n336 B.n335 585
R1016 B.n334 B.n186 585
R1017 B.n333 B.n332 585
R1018 B.n330 B.n187 585
R1019 B.n328 B.n327 585
R1020 B.n326 B.n188 585
R1021 B.n324 B.n323 585
R1022 B.n321 B.n191 585
R1023 B.n319 B.n318 585
R1024 B.n317 B.n192 585
R1025 B.n316 B.n315 585
R1026 B.n313 B.n193 585
R1027 B.n311 B.n310 585
R1028 B.n309 B.n194 585
R1029 B.n308 B.n307 585
R1030 B.n305 B.n304 585
R1031 B.n303 B.n302 585
R1032 B.n301 B.n199 585
R1033 B.n299 B.n298 585
R1034 B.n297 B.n200 585
R1035 B.n296 B.n295 585
R1036 B.n293 B.n201 585
R1037 B.n291 B.n290 585
R1038 B.n289 B.n202 585
R1039 B.n288 B.n287 585
R1040 B.n285 B.n203 585
R1041 B.n283 B.n282 585
R1042 B.n281 B.n204 585
R1043 B.n280 B.n279 585
R1044 B.n277 B.n205 585
R1045 B.n275 B.n274 585
R1046 B.n273 B.n206 585
R1047 B.n272 B.n271 585
R1048 B.n269 B.n207 585
R1049 B.n267 B.n266 585
R1050 B.n265 B.n208 585
R1051 B.n264 B.n263 585
R1052 B.n261 B.n209 585
R1053 B.n259 B.n258 585
R1054 B.n257 B.n210 585
R1055 B.n256 B.n255 585
R1056 B.n253 B.n211 585
R1057 B.n251 B.n250 585
R1058 B.n249 B.n212 585
R1059 B.n248 B.n247 585
R1060 B.n245 B.n213 585
R1061 B.n243 B.n242 585
R1062 B.n241 B.n214 585
R1063 B.n240 B.n239 585
R1064 B.n237 B.n215 585
R1065 B.n235 B.n234 585
R1066 B.n233 B.n216 585
R1067 B.n232 B.n231 585
R1068 B.n229 B.n217 585
R1069 B.n227 B.n226 585
R1070 B.n225 B.n218 585
R1071 B.n224 B.n223 585
R1072 B.n221 B.n219 585
R1073 B.n164 B.n163 585
R1074 B.n413 B.n412 585
R1075 B.n414 B.n413 585
R1076 B.n160 B.n159 585
R1077 B.n161 B.n160 585
R1078 B.n422 B.n421 585
R1079 B.n421 B.n420 585
R1080 B.n423 B.n158 585
R1081 B.n158 B.n157 585
R1082 B.n425 B.n424 585
R1083 B.n426 B.n425 585
R1084 B.n152 B.n151 585
R1085 B.n153 B.n152 585
R1086 B.n434 B.n433 585
R1087 B.n433 B.n432 585
R1088 B.n435 B.n150 585
R1089 B.n150 B.n149 585
R1090 B.n437 B.n436 585
R1091 B.n438 B.n437 585
R1092 B.n144 B.n143 585
R1093 B.n145 B.n144 585
R1094 B.n447 B.n446 585
R1095 B.n446 B.n445 585
R1096 B.n448 B.n142 585
R1097 B.n444 B.n142 585
R1098 B.n450 B.n449 585
R1099 B.n451 B.n450 585
R1100 B.n137 B.n136 585
R1101 B.n138 B.n137 585
R1102 B.n460 B.n459 585
R1103 B.n459 B.n458 585
R1104 B.n461 B.n135 585
R1105 B.n457 B.n135 585
R1106 B.n463 B.n462 585
R1107 B.n464 B.n463 585
R1108 B.n130 B.n129 585
R1109 B.n131 B.n130 585
R1110 B.n473 B.n472 585
R1111 B.n472 B.n471 585
R1112 B.n474 B.n128 585
R1113 B.n470 B.n128 585
R1114 B.n476 B.n475 585
R1115 B.n477 B.n476 585
R1116 B.n123 B.n122 585
R1117 B.n124 B.n123 585
R1118 B.n486 B.n485 585
R1119 B.n485 B.n484 585
R1120 B.n487 B.n121 585
R1121 B.n483 B.n121 585
R1122 B.n489 B.n488 585
R1123 B.n490 B.n489 585
R1124 B.n116 B.n115 585
R1125 B.n117 B.n116 585
R1126 B.n500 B.n499 585
R1127 B.n499 B.n498 585
R1128 B.n501 B.n114 585
R1129 B.n497 B.n114 585
R1130 B.n503 B.n502 585
R1131 B.n504 B.n503 585
R1132 B.n3 B.n0 585
R1133 B.n4 B.n3 585
R1134 B.n801 B.n1 585
R1135 B.n802 B.n801 585
R1136 B.n800 B.n799 585
R1137 B.n800 B.n8 585
R1138 B.n798 B.n9 585
R1139 B.n12 B.n9 585
R1140 B.n797 B.n796 585
R1141 B.n796 B.n795 585
R1142 B.n11 B.n10 585
R1143 B.n794 B.n11 585
R1144 B.n792 B.n791 585
R1145 B.n793 B.n792 585
R1146 B.n790 B.n16 585
R1147 B.n19 B.n16 585
R1148 B.n789 B.n788 585
R1149 B.n788 B.n787 585
R1150 B.n18 B.n17 585
R1151 B.n786 B.n18 585
R1152 B.n784 B.n783 585
R1153 B.n785 B.n784 585
R1154 B.n782 B.n23 585
R1155 B.n26 B.n23 585
R1156 B.n781 B.n780 585
R1157 B.n780 B.n779 585
R1158 B.n25 B.n24 585
R1159 B.n778 B.n25 585
R1160 B.n776 B.n775 585
R1161 B.n777 B.n776 585
R1162 B.n774 B.n30 585
R1163 B.n33 B.n30 585
R1164 B.n773 B.n772 585
R1165 B.n772 B.n771 585
R1166 B.n32 B.n31 585
R1167 B.n770 B.n32 585
R1168 B.n768 B.n767 585
R1169 B.n769 B.n768 585
R1170 B.n766 B.n37 585
R1171 B.n40 B.n37 585
R1172 B.n765 B.n764 585
R1173 B.n764 B.n763 585
R1174 B.n39 B.n38 585
R1175 B.n762 B.n39 585
R1176 B.n760 B.n759 585
R1177 B.n761 B.n760 585
R1178 B.n758 B.n45 585
R1179 B.n45 B.n44 585
R1180 B.n757 B.n756 585
R1181 B.n756 B.n755 585
R1182 B.n47 B.n46 585
R1183 B.n754 B.n47 585
R1184 B.n752 B.n751 585
R1185 B.n753 B.n752 585
R1186 B.n750 B.n52 585
R1187 B.n52 B.n51 585
R1188 B.n749 B.n748 585
R1189 B.n748 B.n747 585
R1190 B.n54 B.n53 585
R1191 B.n746 B.n54 585
R1192 B.n744 B.n743 585
R1193 B.n745 B.n744 585
R1194 B.n805 B.n804 585
R1195 B.n803 B.n2 585
R1196 B.n82 B.t17 523.74
R1197 B.n88 B.t9 523.74
R1198 B.n195 B.t20 523.74
R1199 B.n189 B.t13 523.74
R1200 B.n744 B.n59 506.916
R1201 B.n111 B.n57 506.916
R1202 B.n415 B.n164 506.916
R1203 B.n413 B.n166 506.916
R1204 B.n88 B.t11 318.156
R1205 B.n195 B.t22 318.156
R1206 B.n82 B.t18 318.156
R1207 B.n189 B.t16 318.156
R1208 B.n89 B.t12 293.332
R1209 B.n196 B.t21 293.332
R1210 B.n83 B.t19 293.332
R1211 B.n190 B.t15 293.332
R1212 B.n551 B.n58 256.663
R1213 B.n553 B.n58 256.663
R1214 B.n559 B.n58 256.663
R1215 B.n561 B.n58 256.663
R1216 B.n567 B.n58 256.663
R1217 B.n569 B.n58 256.663
R1218 B.n575 B.n58 256.663
R1219 B.n577 B.n58 256.663
R1220 B.n583 B.n58 256.663
R1221 B.n585 B.n58 256.663
R1222 B.n591 B.n58 256.663
R1223 B.n593 B.n58 256.663
R1224 B.n599 B.n58 256.663
R1225 B.n601 B.n58 256.663
R1226 B.n607 B.n58 256.663
R1227 B.n609 B.n58 256.663
R1228 B.n615 B.n58 256.663
R1229 B.n617 B.n58 256.663
R1230 B.n623 B.n58 256.663
R1231 B.n625 B.n58 256.663
R1232 B.n631 B.n58 256.663
R1233 B.n633 B.n58 256.663
R1234 B.n640 B.n58 256.663
R1235 B.n642 B.n58 256.663
R1236 B.n648 B.n58 256.663
R1237 B.n650 B.n58 256.663
R1238 B.n657 B.n58 256.663
R1239 B.n659 B.n58 256.663
R1240 B.n665 B.n58 256.663
R1241 B.n667 B.n58 256.663
R1242 B.n673 B.n58 256.663
R1243 B.n675 B.n58 256.663
R1244 B.n681 B.n58 256.663
R1245 B.n683 B.n58 256.663
R1246 B.n689 B.n58 256.663
R1247 B.n691 B.n58 256.663
R1248 B.n697 B.n58 256.663
R1249 B.n699 B.n58 256.663
R1250 B.n705 B.n58 256.663
R1251 B.n707 B.n58 256.663
R1252 B.n713 B.n58 256.663
R1253 B.n715 B.n58 256.663
R1254 B.n721 B.n58 256.663
R1255 B.n723 B.n58 256.663
R1256 B.n729 B.n58 256.663
R1257 B.n731 B.n58 256.663
R1258 B.n737 B.n58 256.663
R1259 B.n739 B.n58 256.663
R1260 B.n408 B.n165 256.663
R1261 B.n168 B.n165 256.663
R1262 B.n401 B.n165 256.663
R1263 B.n395 B.n165 256.663
R1264 B.n393 B.n165 256.663
R1265 B.n387 B.n165 256.663
R1266 B.n385 B.n165 256.663
R1267 B.n379 B.n165 256.663
R1268 B.n377 B.n165 256.663
R1269 B.n371 B.n165 256.663
R1270 B.n369 B.n165 256.663
R1271 B.n363 B.n165 256.663
R1272 B.n361 B.n165 256.663
R1273 B.n355 B.n165 256.663
R1274 B.n353 B.n165 256.663
R1275 B.n347 B.n165 256.663
R1276 B.n345 B.n165 256.663
R1277 B.n339 B.n165 256.663
R1278 B.n337 B.n165 256.663
R1279 B.n331 B.n165 256.663
R1280 B.n329 B.n165 256.663
R1281 B.n322 B.n165 256.663
R1282 B.n320 B.n165 256.663
R1283 B.n314 B.n165 256.663
R1284 B.n312 B.n165 256.663
R1285 B.n306 B.n165 256.663
R1286 B.n198 B.n165 256.663
R1287 B.n300 B.n165 256.663
R1288 B.n294 B.n165 256.663
R1289 B.n292 B.n165 256.663
R1290 B.n286 B.n165 256.663
R1291 B.n284 B.n165 256.663
R1292 B.n278 B.n165 256.663
R1293 B.n276 B.n165 256.663
R1294 B.n270 B.n165 256.663
R1295 B.n268 B.n165 256.663
R1296 B.n262 B.n165 256.663
R1297 B.n260 B.n165 256.663
R1298 B.n254 B.n165 256.663
R1299 B.n252 B.n165 256.663
R1300 B.n246 B.n165 256.663
R1301 B.n244 B.n165 256.663
R1302 B.n238 B.n165 256.663
R1303 B.n236 B.n165 256.663
R1304 B.n230 B.n165 256.663
R1305 B.n228 B.n165 256.663
R1306 B.n222 B.n165 256.663
R1307 B.n220 B.n165 256.663
R1308 B.n807 B.n806 256.663
R1309 B.n740 B.n738 163.367
R1310 B.n736 B.n61 163.367
R1311 B.n732 B.n730 163.367
R1312 B.n728 B.n63 163.367
R1313 B.n724 B.n722 163.367
R1314 B.n720 B.n65 163.367
R1315 B.n716 B.n714 163.367
R1316 B.n712 B.n67 163.367
R1317 B.n708 B.n706 163.367
R1318 B.n704 B.n69 163.367
R1319 B.n700 B.n698 163.367
R1320 B.n696 B.n71 163.367
R1321 B.n692 B.n690 163.367
R1322 B.n688 B.n73 163.367
R1323 B.n684 B.n682 163.367
R1324 B.n680 B.n75 163.367
R1325 B.n676 B.n674 163.367
R1326 B.n672 B.n77 163.367
R1327 B.n668 B.n666 163.367
R1328 B.n664 B.n79 163.367
R1329 B.n660 B.n658 163.367
R1330 B.n656 B.n81 163.367
R1331 B.n651 B.n649 163.367
R1332 B.n647 B.n85 163.367
R1333 B.n643 B.n641 163.367
R1334 B.n639 B.n87 163.367
R1335 B.n634 B.n632 163.367
R1336 B.n630 B.n91 163.367
R1337 B.n626 B.n624 163.367
R1338 B.n622 B.n93 163.367
R1339 B.n618 B.n616 163.367
R1340 B.n614 B.n95 163.367
R1341 B.n610 B.n608 163.367
R1342 B.n606 B.n97 163.367
R1343 B.n602 B.n600 163.367
R1344 B.n598 B.n99 163.367
R1345 B.n594 B.n592 163.367
R1346 B.n590 B.n101 163.367
R1347 B.n586 B.n584 163.367
R1348 B.n582 B.n103 163.367
R1349 B.n578 B.n576 163.367
R1350 B.n574 B.n105 163.367
R1351 B.n570 B.n568 163.367
R1352 B.n566 B.n107 163.367
R1353 B.n562 B.n560 163.367
R1354 B.n558 B.n109 163.367
R1355 B.n554 B.n552 163.367
R1356 B.n550 B.n111 163.367
R1357 B.n415 B.n162 163.367
R1358 B.n419 B.n162 163.367
R1359 B.n419 B.n156 163.367
R1360 B.n427 B.n156 163.367
R1361 B.n427 B.n154 163.367
R1362 B.n431 B.n154 163.367
R1363 B.n431 B.n148 163.367
R1364 B.n439 B.n148 163.367
R1365 B.n439 B.n146 163.367
R1366 B.n443 B.n146 163.367
R1367 B.n443 B.n141 163.367
R1368 B.n452 B.n141 163.367
R1369 B.n452 B.n139 163.367
R1370 B.n456 B.n139 163.367
R1371 B.n456 B.n134 163.367
R1372 B.n465 B.n134 163.367
R1373 B.n465 B.n132 163.367
R1374 B.n469 B.n132 163.367
R1375 B.n469 B.n127 163.367
R1376 B.n478 B.n127 163.367
R1377 B.n478 B.n125 163.367
R1378 B.n482 B.n125 163.367
R1379 B.n482 B.n120 163.367
R1380 B.n491 B.n120 163.367
R1381 B.n491 B.n118 163.367
R1382 B.n496 B.n118 163.367
R1383 B.n496 B.n113 163.367
R1384 B.n505 B.n113 163.367
R1385 B.n506 B.n505 163.367
R1386 B.n506 B.n5 163.367
R1387 B.n6 B.n5 163.367
R1388 B.n7 B.n6 163.367
R1389 B.n512 B.n7 163.367
R1390 B.n513 B.n512 163.367
R1391 B.n513 B.n13 163.367
R1392 B.n14 B.n13 163.367
R1393 B.n15 B.n14 163.367
R1394 B.n518 B.n15 163.367
R1395 B.n518 B.n20 163.367
R1396 B.n21 B.n20 163.367
R1397 B.n22 B.n21 163.367
R1398 B.n523 B.n22 163.367
R1399 B.n523 B.n27 163.367
R1400 B.n28 B.n27 163.367
R1401 B.n29 B.n28 163.367
R1402 B.n528 B.n29 163.367
R1403 B.n528 B.n34 163.367
R1404 B.n35 B.n34 163.367
R1405 B.n36 B.n35 163.367
R1406 B.n533 B.n36 163.367
R1407 B.n533 B.n41 163.367
R1408 B.n42 B.n41 163.367
R1409 B.n43 B.n42 163.367
R1410 B.n538 B.n43 163.367
R1411 B.n538 B.n48 163.367
R1412 B.n49 B.n48 163.367
R1413 B.n50 B.n49 163.367
R1414 B.n543 B.n50 163.367
R1415 B.n543 B.n55 163.367
R1416 B.n56 B.n55 163.367
R1417 B.n57 B.n56 163.367
R1418 B.n409 B.n407 163.367
R1419 B.n407 B.n406 163.367
R1420 B.n403 B.n402 163.367
R1421 B.n400 B.n170 163.367
R1422 B.n396 B.n394 163.367
R1423 B.n392 B.n172 163.367
R1424 B.n388 B.n386 163.367
R1425 B.n384 B.n174 163.367
R1426 B.n380 B.n378 163.367
R1427 B.n376 B.n176 163.367
R1428 B.n372 B.n370 163.367
R1429 B.n368 B.n178 163.367
R1430 B.n364 B.n362 163.367
R1431 B.n360 B.n180 163.367
R1432 B.n356 B.n354 163.367
R1433 B.n352 B.n182 163.367
R1434 B.n348 B.n346 163.367
R1435 B.n344 B.n184 163.367
R1436 B.n340 B.n338 163.367
R1437 B.n336 B.n186 163.367
R1438 B.n332 B.n330 163.367
R1439 B.n328 B.n188 163.367
R1440 B.n323 B.n321 163.367
R1441 B.n319 B.n192 163.367
R1442 B.n315 B.n313 163.367
R1443 B.n311 B.n194 163.367
R1444 B.n307 B.n305 163.367
R1445 B.n302 B.n301 163.367
R1446 B.n299 B.n200 163.367
R1447 B.n295 B.n293 163.367
R1448 B.n291 B.n202 163.367
R1449 B.n287 B.n285 163.367
R1450 B.n283 B.n204 163.367
R1451 B.n279 B.n277 163.367
R1452 B.n275 B.n206 163.367
R1453 B.n271 B.n269 163.367
R1454 B.n267 B.n208 163.367
R1455 B.n263 B.n261 163.367
R1456 B.n259 B.n210 163.367
R1457 B.n255 B.n253 163.367
R1458 B.n251 B.n212 163.367
R1459 B.n247 B.n245 163.367
R1460 B.n243 B.n214 163.367
R1461 B.n239 B.n237 163.367
R1462 B.n235 B.n216 163.367
R1463 B.n231 B.n229 163.367
R1464 B.n227 B.n218 163.367
R1465 B.n223 B.n221 163.367
R1466 B.n413 B.n160 163.367
R1467 B.n421 B.n160 163.367
R1468 B.n421 B.n158 163.367
R1469 B.n425 B.n158 163.367
R1470 B.n425 B.n152 163.367
R1471 B.n433 B.n152 163.367
R1472 B.n433 B.n150 163.367
R1473 B.n437 B.n150 163.367
R1474 B.n437 B.n144 163.367
R1475 B.n446 B.n144 163.367
R1476 B.n446 B.n142 163.367
R1477 B.n450 B.n142 163.367
R1478 B.n450 B.n137 163.367
R1479 B.n459 B.n137 163.367
R1480 B.n459 B.n135 163.367
R1481 B.n463 B.n135 163.367
R1482 B.n463 B.n130 163.367
R1483 B.n472 B.n130 163.367
R1484 B.n472 B.n128 163.367
R1485 B.n476 B.n128 163.367
R1486 B.n476 B.n123 163.367
R1487 B.n485 B.n123 163.367
R1488 B.n485 B.n121 163.367
R1489 B.n489 B.n121 163.367
R1490 B.n489 B.n116 163.367
R1491 B.n499 B.n116 163.367
R1492 B.n499 B.n114 163.367
R1493 B.n503 B.n114 163.367
R1494 B.n503 B.n3 163.367
R1495 B.n805 B.n3 163.367
R1496 B.n801 B.n2 163.367
R1497 B.n801 B.n800 163.367
R1498 B.n800 B.n9 163.367
R1499 B.n796 B.n9 163.367
R1500 B.n796 B.n11 163.367
R1501 B.n792 B.n11 163.367
R1502 B.n792 B.n16 163.367
R1503 B.n788 B.n16 163.367
R1504 B.n788 B.n18 163.367
R1505 B.n784 B.n18 163.367
R1506 B.n784 B.n23 163.367
R1507 B.n780 B.n23 163.367
R1508 B.n780 B.n25 163.367
R1509 B.n776 B.n25 163.367
R1510 B.n776 B.n30 163.367
R1511 B.n772 B.n30 163.367
R1512 B.n772 B.n32 163.367
R1513 B.n768 B.n32 163.367
R1514 B.n768 B.n37 163.367
R1515 B.n764 B.n37 163.367
R1516 B.n764 B.n39 163.367
R1517 B.n760 B.n39 163.367
R1518 B.n760 B.n45 163.367
R1519 B.n756 B.n45 163.367
R1520 B.n756 B.n47 163.367
R1521 B.n752 B.n47 163.367
R1522 B.n752 B.n52 163.367
R1523 B.n748 B.n52 163.367
R1524 B.n748 B.n54 163.367
R1525 B.n744 B.n54 163.367
R1526 B.n414 B.n165 84.0262
R1527 B.n745 B.n58 84.0262
R1528 B.n739 B.n59 71.676
R1529 B.n738 B.n737 71.676
R1530 B.n731 B.n61 71.676
R1531 B.n730 B.n729 71.676
R1532 B.n723 B.n63 71.676
R1533 B.n722 B.n721 71.676
R1534 B.n715 B.n65 71.676
R1535 B.n714 B.n713 71.676
R1536 B.n707 B.n67 71.676
R1537 B.n706 B.n705 71.676
R1538 B.n699 B.n69 71.676
R1539 B.n698 B.n697 71.676
R1540 B.n691 B.n71 71.676
R1541 B.n690 B.n689 71.676
R1542 B.n683 B.n73 71.676
R1543 B.n682 B.n681 71.676
R1544 B.n675 B.n75 71.676
R1545 B.n674 B.n673 71.676
R1546 B.n667 B.n77 71.676
R1547 B.n666 B.n665 71.676
R1548 B.n659 B.n79 71.676
R1549 B.n658 B.n657 71.676
R1550 B.n650 B.n81 71.676
R1551 B.n649 B.n648 71.676
R1552 B.n642 B.n85 71.676
R1553 B.n641 B.n640 71.676
R1554 B.n633 B.n87 71.676
R1555 B.n632 B.n631 71.676
R1556 B.n625 B.n91 71.676
R1557 B.n624 B.n623 71.676
R1558 B.n617 B.n93 71.676
R1559 B.n616 B.n615 71.676
R1560 B.n609 B.n95 71.676
R1561 B.n608 B.n607 71.676
R1562 B.n601 B.n97 71.676
R1563 B.n600 B.n599 71.676
R1564 B.n593 B.n99 71.676
R1565 B.n592 B.n591 71.676
R1566 B.n585 B.n101 71.676
R1567 B.n584 B.n583 71.676
R1568 B.n577 B.n103 71.676
R1569 B.n576 B.n575 71.676
R1570 B.n569 B.n105 71.676
R1571 B.n568 B.n567 71.676
R1572 B.n561 B.n107 71.676
R1573 B.n560 B.n559 71.676
R1574 B.n553 B.n109 71.676
R1575 B.n552 B.n551 71.676
R1576 B.n551 B.n550 71.676
R1577 B.n554 B.n553 71.676
R1578 B.n559 B.n558 71.676
R1579 B.n562 B.n561 71.676
R1580 B.n567 B.n566 71.676
R1581 B.n570 B.n569 71.676
R1582 B.n575 B.n574 71.676
R1583 B.n578 B.n577 71.676
R1584 B.n583 B.n582 71.676
R1585 B.n586 B.n585 71.676
R1586 B.n591 B.n590 71.676
R1587 B.n594 B.n593 71.676
R1588 B.n599 B.n598 71.676
R1589 B.n602 B.n601 71.676
R1590 B.n607 B.n606 71.676
R1591 B.n610 B.n609 71.676
R1592 B.n615 B.n614 71.676
R1593 B.n618 B.n617 71.676
R1594 B.n623 B.n622 71.676
R1595 B.n626 B.n625 71.676
R1596 B.n631 B.n630 71.676
R1597 B.n634 B.n633 71.676
R1598 B.n640 B.n639 71.676
R1599 B.n643 B.n642 71.676
R1600 B.n648 B.n647 71.676
R1601 B.n651 B.n650 71.676
R1602 B.n657 B.n656 71.676
R1603 B.n660 B.n659 71.676
R1604 B.n665 B.n664 71.676
R1605 B.n668 B.n667 71.676
R1606 B.n673 B.n672 71.676
R1607 B.n676 B.n675 71.676
R1608 B.n681 B.n680 71.676
R1609 B.n684 B.n683 71.676
R1610 B.n689 B.n688 71.676
R1611 B.n692 B.n691 71.676
R1612 B.n697 B.n696 71.676
R1613 B.n700 B.n699 71.676
R1614 B.n705 B.n704 71.676
R1615 B.n708 B.n707 71.676
R1616 B.n713 B.n712 71.676
R1617 B.n716 B.n715 71.676
R1618 B.n721 B.n720 71.676
R1619 B.n724 B.n723 71.676
R1620 B.n729 B.n728 71.676
R1621 B.n732 B.n731 71.676
R1622 B.n737 B.n736 71.676
R1623 B.n740 B.n739 71.676
R1624 B.n408 B.n166 71.676
R1625 B.n406 B.n168 71.676
R1626 B.n402 B.n401 71.676
R1627 B.n395 B.n170 71.676
R1628 B.n394 B.n393 71.676
R1629 B.n387 B.n172 71.676
R1630 B.n386 B.n385 71.676
R1631 B.n379 B.n174 71.676
R1632 B.n378 B.n377 71.676
R1633 B.n371 B.n176 71.676
R1634 B.n370 B.n369 71.676
R1635 B.n363 B.n178 71.676
R1636 B.n362 B.n361 71.676
R1637 B.n355 B.n180 71.676
R1638 B.n354 B.n353 71.676
R1639 B.n347 B.n182 71.676
R1640 B.n346 B.n345 71.676
R1641 B.n339 B.n184 71.676
R1642 B.n338 B.n337 71.676
R1643 B.n331 B.n186 71.676
R1644 B.n330 B.n329 71.676
R1645 B.n322 B.n188 71.676
R1646 B.n321 B.n320 71.676
R1647 B.n314 B.n192 71.676
R1648 B.n313 B.n312 71.676
R1649 B.n306 B.n194 71.676
R1650 B.n305 B.n198 71.676
R1651 B.n301 B.n300 71.676
R1652 B.n294 B.n200 71.676
R1653 B.n293 B.n292 71.676
R1654 B.n286 B.n202 71.676
R1655 B.n285 B.n284 71.676
R1656 B.n278 B.n204 71.676
R1657 B.n277 B.n276 71.676
R1658 B.n270 B.n206 71.676
R1659 B.n269 B.n268 71.676
R1660 B.n262 B.n208 71.676
R1661 B.n261 B.n260 71.676
R1662 B.n254 B.n210 71.676
R1663 B.n253 B.n252 71.676
R1664 B.n246 B.n212 71.676
R1665 B.n245 B.n244 71.676
R1666 B.n238 B.n214 71.676
R1667 B.n237 B.n236 71.676
R1668 B.n230 B.n216 71.676
R1669 B.n229 B.n228 71.676
R1670 B.n222 B.n218 71.676
R1671 B.n221 B.n220 71.676
R1672 B.n409 B.n408 71.676
R1673 B.n403 B.n168 71.676
R1674 B.n401 B.n400 71.676
R1675 B.n396 B.n395 71.676
R1676 B.n393 B.n392 71.676
R1677 B.n388 B.n387 71.676
R1678 B.n385 B.n384 71.676
R1679 B.n380 B.n379 71.676
R1680 B.n377 B.n376 71.676
R1681 B.n372 B.n371 71.676
R1682 B.n369 B.n368 71.676
R1683 B.n364 B.n363 71.676
R1684 B.n361 B.n360 71.676
R1685 B.n356 B.n355 71.676
R1686 B.n353 B.n352 71.676
R1687 B.n348 B.n347 71.676
R1688 B.n345 B.n344 71.676
R1689 B.n340 B.n339 71.676
R1690 B.n337 B.n336 71.676
R1691 B.n332 B.n331 71.676
R1692 B.n329 B.n328 71.676
R1693 B.n323 B.n322 71.676
R1694 B.n320 B.n319 71.676
R1695 B.n315 B.n314 71.676
R1696 B.n312 B.n311 71.676
R1697 B.n307 B.n306 71.676
R1698 B.n302 B.n198 71.676
R1699 B.n300 B.n299 71.676
R1700 B.n295 B.n294 71.676
R1701 B.n292 B.n291 71.676
R1702 B.n287 B.n286 71.676
R1703 B.n284 B.n283 71.676
R1704 B.n279 B.n278 71.676
R1705 B.n276 B.n275 71.676
R1706 B.n271 B.n270 71.676
R1707 B.n268 B.n267 71.676
R1708 B.n263 B.n262 71.676
R1709 B.n260 B.n259 71.676
R1710 B.n255 B.n254 71.676
R1711 B.n252 B.n251 71.676
R1712 B.n247 B.n246 71.676
R1713 B.n244 B.n243 71.676
R1714 B.n239 B.n238 71.676
R1715 B.n236 B.n235 71.676
R1716 B.n231 B.n230 71.676
R1717 B.n228 B.n227 71.676
R1718 B.n223 B.n222 71.676
R1719 B.n220 B.n164 71.676
R1720 B.n806 B.n805 71.676
R1721 B.n806 B.n2 71.676
R1722 B.n654 B.n83 59.5399
R1723 B.n636 B.n89 59.5399
R1724 B.n197 B.n196 59.5399
R1725 B.n325 B.n190 59.5399
R1726 B.n414 B.n161 41.7067
R1727 B.n420 B.n161 41.7067
R1728 B.n420 B.n157 41.7067
R1729 B.n426 B.n157 41.7067
R1730 B.n432 B.n153 41.7067
R1731 B.n432 B.n149 41.7067
R1732 B.n438 B.n149 41.7067
R1733 B.n438 B.n145 41.7067
R1734 B.n445 B.n145 41.7067
R1735 B.n445 B.n444 41.7067
R1736 B.n451 B.n138 41.7067
R1737 B.n458 B.n138 41.7067
R1738 B.n458 B.n457 41.7067
R1739 B.n464 B.n131 41.7067
R1740 B.n471 B.n131 41.7067
R1741 B.n471 B.n470 41.7067
R1742 B.n477 B.n124 41.7067
R1743 B.n484 B.n124 41.7067
R1744 B.n484 B.n483 41.7067
R1745 B.n490 B.n117 41.7067
R1746 B.n498 B.n117 41.7067
R1747 B.n498 B.n497 41.7067
R1748 B.n504 B.n4 41.7067
R1749 B.n804 B.n4 41.7067
R1750 B.n804 B.n803 41.7067
R1751 B.n803 B.n802 41.7067
R1752 B.n802 B.n8 41.7067
R1753 B.n795 B.n12 41.7067
R1754 B.n795 B.n794 41.7067
R1755 B.n794 B.n793 41.7067
R1756 B.n787 B.n19 41.7067
R1757 B.n787 B.n786 41.7067
R1758 B.n786 B.n785 41.7067
R1759 B.n779 B.n26 41.7067
R1760 B.n779 B.n778 41.7067
R1761 B.n778 B.n777 41.7067
R1762 B.n771 B.n33 41.7067
R1763 B.n771 B.n770 41.7067
R1764 B.n770 B.n769 41.7067
R1765 B.n763 B.n40 41.7067
R1766 B.n763 B.n762 41.7067
R1767 B.n762 B.n761 41.7067
R1768 B.n761 B.n44 41.7067
R1769 B.n755 B.n44 41.7067
R1770 B.n755 B.n754 41.7067
R1771 B.n753 B.n51 41.7067
R1772 B.n747 B.n51 41.7067
R1773 B.n747 B.n746 41.7067
R1774 B.n746 B.n745 41.7067
R1775 B.n426 B.t14 41.0933
R1776 B.n504 B.t3 41.0933
R1777 B.t7 B.n8 41.0933
R1778 B.t10 B.n753 41.0933
R1779 B.n444 B.t0 39.8667
R1780 B.n40 B.t6 39.8667
R1781 B.n412 B.n411 32.9371
R1782 B.n416 B.n163 32.9371
R1783 B.n548 B.n547 32.9371
R1784 B.n743 B.n742 32.9371
R1785 B.n490 B.t2 31.2801
R1786 B.n793 B.t5 31.2801
R1787 B.n457 B.t23 30.0535
R1788 B.n33 B.t1 30.0535
R1789 B.n83 B.n82 24.8247
R1790 B.n89 B.n88 24.8247
R1791 B.n196 B.n195 24.8247
R1792 B.n190 B.n189 24.8247
R1793 B.n477 B.t4 21.4669
R1794 B.n785 B.t8 21.4669
R1795 B.n470 B.t4 20.2403
R1796 B.n26 B.t8 20.2403
R1797 B B.n807 18.0485
R1798 B.n464 B.t23 11.6537
R1799 B.n777 B.t1 11.6537
R1800 B.n412 B.n159 10.6151
R1801 B.n422 B.n159 10.6151
R1802 B.n423 B.n422 10.6151
R1803 B.n424 B.n423 10.6151
R1804 B.n424 B.n151 10.6151
R1805 B.n434 B.n151 10.6151
R1806 B.n435 B.n434 10.6151
R1807 B.n436 B.n435 10.6151
R1808 B.n436 B.n143 10.6151
R1809 B.n447 B.n143 10.6151
R1810 B.n448 B.n447 10.6151
R1811 B.n449 B.n448 10.6151
R1812 B.n449 B.n136 10.6151
R1813 B.n460 B.n136 10.6151
R1814 B.n461 B.n460 10.6151
R1815 B.n462 B.n461 10.6151
R1816 B.n462 B.n129 10.6151
R1817 B.n473 B.n129 10.6151
R1818 B.n474 B.n473 10.6151
R1819 B.n475 B.n474 10.6151
R1820 B.n475 B.n122 10.6151
R1821 B.n486 B.n122 10.6151
R1822 B.n487 B.n486 10.6151
R1823 B.n488 B.n487 10.6151
R1824 B.n488 B.n115 10.6151
R1825 B.n500 B.n115 10.6151
R1826 B.n501 B.n500 10.6151
R1827 B.n502 B.n501 10.6151
R1828 B.n502 B.n0 10.6151
R1829 B.n411 B.n410 10.6151
R1830 B.n410 B.n167 10.6151
R1831 B.n405 B.n167 10.6151
R1832 B.n405 B.n404 10.6151
R1833 B.n404 B.n169 10.6151
R1834 B.n399 B.n169 10.6151
R1835 B.n399 B.n398 10.6151
R1836 B.n398 B.n397 10.6151
R1837 B.n397 B.n171 10.6151
R1838 B.n391 B.n171 10.6151
R1839 B.n391 B.n390 10.6151
R1840 B.n390 B.n389 10.6151
R1841 B.n389 B.n173 10.6151
R1842 B.n383 B.n173 10.6151
R1843 B.n383 B.n382 10.6151
R1844 B.n382 B.n381 10.6151
R1845 B.n381 B.n175 10.6151
R1846 B.n375 B.n175 10.6151
R1847 B.n375 B.n374 10.6151
R1848 B.n374 B.n373 10.6151
R1849 B.n373 B.n177 10.6151
R1850 B.n367 B.n177 10.6151
R1851 B.n367 B.n366 10.6151
R1852 B.n366 B.n365 10.6151
R1853 B.n365 B.n179 10.6151
R1854 B.n359 B.n179 10.6151
R1855 B.n359 B.n358 10.6151
R1856 B.n358 B.n357 10.6151
R1857 B.n357 B.n181 10.6151
R1858 B.n351 B.n181 10.6151
R1859 B.n351 B.n350 10.6151
R1860 B.n350 B.n349 10.6151
R1861 B.n349 B.n183 10.6151
R1862 B.n343 B.n183 10.6151
R1863 B.n343 B.n342 10.6151
R1864 B.n342 B.n341 10.6151
R1865 B.n341 B.n185 10.6151
R1866 B.n335 B.n185 10.6151
R1867 B.n335 B.n334 10.6151
R1868 B.n334 B.n333 10.6151
R1869 B.n333 B.n187 10.6151
R1870 B.n327 B.n187 10.6151
R1871 B.n327 B.n326 10.6151
R1872 B.n324 B.n191 10.6151
R1873 B.n318 B.n191 10.6151
R1874 B.n318 B.n317 10.6151
R1875 B.n317 B.n316 10.6151
R1876 B.n316 B.n193 10.6151
R1877 B.n310 B.n193 10.6151
R1878 B.n310 B.n309 10.6151
R1879 B.n309 B.n308 10.6151
R1880 B.n304 B.n303 10.6151
R1881 B.n303 B.n199 10.6151
R1882 B.n298 B.n199 10.6151
R1883 B.n298 B.n297 10.6151
R1884 B.n297 B.n296 10.6151
R1885 B.n296 B.n201 10.6151
R1886 B.n290 B.n201 10.6151
R1887 B.n290 B.n289 10.6151
R1888 B.n289 B.n288 10.6151
R1889 B.n288 B.n203 10.6151
R1890 B.n282 B.n203 10.6151
R1891 B.n282 B.n281 10.6151
R1892 B.n281 B.n280 10.6151
R1893 B.n280 B.n205 10.6151
R1894 B.n274 B.n205 10.6151
R1895 B.n274 B.n273 10.6151
R1896 B.n273 B.n272 10.6151
R1897 B.n272 B.n207 10.6151
R1898 B.n266 B.n207 10.6151
R1899 B.n266 B.n265 10.6151
R1900 B.n265 B.n264 10.6151
R1901 B.n264 B.n209 10.6151
R1902 B.n258 B.n209 10.6151
R1903 B.n258 B.n257 10.6151
R1904 B.n257 B.n256 10.6151
R1905 B.n256 B.n211 10.6151
R1906 B.n250 B.n211 10.6151
R1907 B.n250 B.n249 10.6151
R1908 B.n249 B.n248 10.6151
R1909 B.n248 B.n213 10.6151
R1910 B.n242 B.n213 10.6151
R1911 B.n242 B.n241 10.6151
R1912 B.n241 B.n240 10.6151
R1913 B.n240 B.n215 10.6151
R1914 B.n234 B.n215 10.6151
R1915 B.n234 B.n233 10.6151
R1916 B.n233 B.n232 10.6151
R1917 B.n232 B.n217 10.6151
R1918 B.n226 B.n217 10.6151
R1919 B.n226 B.n225 10.6151
R1920 B.n225 B.n224 10.6151
R1921 B.n224 B.n219 10.6151
R1922 B.n219 B.n163 10.6151
R1923 B.n417 B.n416 10.6151
R1924 B.n418 B.n417 10.6151
R1925 B.n418 B.n155 10.6151
R1926 B.n428 B.n155 10.6151
R1927 B.n429 B.n428 10.6151
R1928 B.n430 B.n429 10.6151
R1929 B.n430 B.n147 10.6151
R1930 B.n440 B.n147 10.6151
R1931 B.n441 B.n440 10.6151
R1932 B.n442 B.n441 10.6151
R1933 B.n442 B.n140 10.6151
R1934 B.n453 B.n140 10.6151
R1935 B.n454 B.n453 10.6151
R1936 B.n455 B.n454 10.6151
R1937 B.n455 B.n133 10.6151
R1938 B.n466 B.n133 10.6151
R1939 B.n467 B.n466 10.6151
R1940 B.n468 B.n467 10.6151
R1941 B.n468 B.n126 10.6151
R1942 B.n479 B.n126 10.6151
R1943 B.n480 B.n479 10.6151
R1944 B.n481 B.n480 10.6151
R1945 B.n481 B.n119 10.6151
R1946 B.n492 B.n119 10.6151
R1947 B.n493 B.n492 10.6151
R1948 B.n495 B.n493 10.6151
R1949 B.n495 B.n494 10.6151
R1950 B.n494 B.n112 10.6151
R1951 B.n507 B.n112 10.6151
R1952 B.n508 B.n507 10.6151
R1953 B.n509 B.n508 10.6151
R1954 B.n510 B.n509 10.6151
R1955 B.n511 B.n510 10.6151
R1956 B.n514 B.n511 10.6151
R1957 B.n515 B.n514 10.6151
R1958 B.n516 B.n515 10.6151
R1959 B.n517 B.n516 10.6151
R1960 B.n519 B.n517 10.6151
R1961 B.n520 B.n519 10.6151
R1962 B.n521 B.n520 10.6151
R1963 B.n522 B.n521 10.6151
R1964 B.n524 B.n522 10.6151
R1965 B.n525 B.n524 10.6151
R1966 B.n526 B.n525 10.6151
R1967 B.n527 B.n526 10.6151
R1968 B.n529 B.n527 10.6151
R1969 B.n530 B.n529 10.6151
R1970 B.n531 B.n530 10.6151
R1971 B.n532 B.n531 10.6151
R1972 B.n534 B.n532 10.6151
R1973 B.n535 B.n534 10.6151
R1974 B.n536 B.n535 10.6151
R1975 B.n537 B.n536 10.6151
R1976 B.n539 B.n537 10.6151
R1977 B.n540 B.n539 10.6151
R1978 B.n541 B.n540 10.6151
R1979 B.n542 B.n541 10.6151
R1980 B.n544 B.n542 10.6151
R1981 B.n545 B.n544 10.6151
R1982 B.n546 B.n545 10.6151
R1983 B.n547 B.n546 10.6151
R1984 B.n799 B.n1 10.6151
R1985 B.n799 B.n798 10.6151
R1986 B.n798 B.n797 10.6151
R1987 B.n797 B.n10 10.6151
R1988 B.n791 B.n10 10.6151
R1989 B.n791 B.n790 10.6151
R1990 B.n790 B.n789 10.6151
R1991 B.n789 B.n17 10.6151
R1992 B.n783 B.n17 10.6151
R1993 B.n783 B.n782 10.6151
R1994 B.n782 B.n781 10.6151
R1995 B.n781 B.n24 10.6151
R1996 B.n775 B.n24 10.6151
R1997 B.n775 B.n774 10.6151
R1998 B.n774 B.n773 10.6151
R1999 B.n773 B.n31 10.6151
R2000 B.n767 B.n31 10.6151
R2001 B.n767 B.n766 10.6151
R2002 B.n766 B.n765 10.6151
R2003 B.n765 B.n38 10.6151
R2004 B.n759 B.n38 10.6151
R2005 B.n759 B.n758 10.6151
R2006 B.n758 B.n757 10.6151
R2007 B.n757 B.n46 10.6151
R2008 B.n751 B.n46 10.6151
R2009 B.n751 B.n750 10.6151
R2010 B.n750 B.n749 10.6151
R2011 B.n749 B.n53 10.6151
R2012 B.n743 B.n53 10.6151
R2013 B.n742 B.n741 10.6151
R2014 B.n741 B.n60 10.6151
R2015 B.n735 B.n60 10.6151
R2016 B.n735 B.n734 10.6151
R2017 B.n734 B.n733 10.6151
R2018 B.n733 B.n62 10.6151
R2019 B.n727 B.n62 10.6151
R2020 B.n727 B.n726 10.6151
R2021 B.n726 B.n725 10.6151
R2022 B.n725 B.n64 10.6151
R2023 B.n719 B.n64 10.6151
R2024 B.n719 B.n718 10.6151
R2025 B.n718 B.n717 10.6151
R2026 B.n717 B.n66 10.6151
R2027 B.n711 B.n66 10.6151
R2028 B.n711 B.n710 10.6151
R2029 B.n710 B.n709 10.6151
R2030 B.n709 B.n68 10.6151
R2031 B.n703 B.n68 10.6151
R2032 B.n703 B.n702 10.6151
R2033 B.n702 B.n701 10.6151
R2034 B.n701 B.n70 10.6151
R2035 B.n695 B.n70 10.6151
R2036 B.n695 B.n694 10.6151
R2037 B.n694 B.n693 10.6151
R2038 B.n693 B.n72 10.6151
R2039 B.n687 B.n72 10.6151
R2040 B.n687 B.n686 10.6151
R2041 B.n686 B.n685 10.6151
R2042 B.n685 B.n74 10.6151
R2043 B.n679 B.n74 10.6151
R2044 B.n679 B.n678 10.6151
R2045 B.n678 B.n677 10.6151
R2046 B.n677 B.n76 10.6151
R2047 B.n671 B.n76 10.6151
R2048 B.n671 B.n670 10.6151
R2049 B.n670 B.n669 10.6151
R2050 B.n669 B.n78 10.6151
R2051 B.n663 B.n78 10.6151
R2052 B.n663 B.n662 10.6151
R2053 B.n662 B.n661 10.6151
R2054 B.n661 B.n80 10.6151
R2055 B.n655 B.n80 10.6151
R2056 B.n653 B.n652 10.6151
R2057 B.n652 B.n84 10.6151
R2058 B.n646 B.n84 10.6151
R2059 B.n646 B.n645 10.6151
R2060 B.n645 B.n644 10.6151
R2061 B.n644 B.n86 10.6151
R2062 B.n638 B.n86 10.6151
R2063 B.n638 B.n637 10.6151
R2064 B.n635 B.n90 10.6151
R2065 B.n629 B.n90 10.6151
R2066 B.n629 B.n628 10.6151
R2067 B.n628 B.n627 10.6151
R2068 B.n627 B.n92 10.6151
R2069 B.n621 B.n92 10.6151
R2070 B.n621 B.n620 10.6151
R2071 B.n620 B.n619 10.6151
R2072 B.n619 B.n94 10.6151
R2073 B.n613 B.n94 10.6151
R2074 B.n613 B.n612 10.6151
R2075 B.n612 B.n611 10.6151
R2076 B.n611 B.n96 10.6151
R2077 B.n605 B.n96 10.6151
R2078 B.n605 B.n604 10.6151
R2079 B.n604 B.n603 10.6151
R2080 B.n603 B.n98 10.6151
R2081 B.n597 B.n98 10.6151
R2082 B.n597 B.n596 10.6151
R2083 B.n596 B.n595 10.6151
R2084 B.n595 B.n100 10.6151
R2085 B.n589 B.n100 10.6151
R2086 B.n589 B.n588 10.6151
R2087 B.n588 B.n587 10.6151
R2088 B.n587 B.n102 10.6151
R2089 B.n581 B.n102 10.6151
R2090 B.n581 B.n580 10.6151
R2091 B.n580 B.n579 10.6151
R2092 B.n579 B.n104 10.6151
R2093 B.n573 B.n104 10.6151
R2094 B.n573 B.n572 10.6151
R2095 B.n572 B.n571 10.6151
R2096 B.n571 B.n106 10.6151
R2097 B.n565 B.n106 10.6151
R2098 B.n565 B.n564 10.6151
R2099 B.n564 B.n563 10.6151
R2100 B.n563 B.n108 10.6151
R2101 B.n557 B.n108 10.6151
R2102 B.n557 B.n556 10.6151
R2103 B.n556 B.n555 10.6151
R2104 B.n555 B.n110 10.6151
R2105 B.n549 B.n110 10.6151
R2106 B.n549 B.n548 10.6151
R2107 B.n483 B.t2 10.427
R2108 B.n19 B.t5 10.427
R2109 B.n807 B.n0 8.11757
R2110 B.n807 B.n1 8.11757
R2111 B.n325 B.n324 6.5566
R2112 B.n308 B.n197 6.5566
R2113 B.n654 B.n653 6.5566
R2114 B.n637 B.n636 6.5566
R2115 B.n326 B.n325 4.05904
R2116 B.n304 B.n197 4.05904
R2117 B.n655 B.n654 4.05904
R2118 B.n636 B.n635 4.05904
R2119 B.n451 B.t0 1.84048
R2120 B.n769 B.t6 1.84048
R2121 B.t14 B.n153 0.613826
R2122 B.n497 B.t3 0.613826
R2123 B.n12 B.t7 0.613826
R2124 B.n754 B.t10 0.613826
R2125 VN.n4 VN.t3 382.909
R2126 VN.n23 VN.t4 382.909
R2127 VN.n17 VN.t7 362.515
R2128 VN.n36 VN.t8 362.515
R2129 VN.n10 VN.t0 321.164
R2130 VN.n5 VN.t2 321.164
R2131 VN.n1 VN.t9 321.164
R2132 VN.n29 VN.t1 321.164
R2133 VN.n24 VN.t6 321.164
R2134 VN.n20 VN.t5 321.164
R2135 VN.n18 VN.n17 161.3
R2136 VN.n37 VN.n36 161.3
R2137 VN.n35 VN.n19 161.3
R2138 VN.n34 VN.n33 161.3
R2139 VN.n32 VN.n31 161.3
R2140 VN.n30 VN.n21 161.3
R2141 VN.n29 VN.n28 161.3
R2142 VN.n27 VN.n22 161.3
R2143 VN.n26 VN.n25 161.3
R2144 VN.n16 VN.n0 161.3
R2145 VN.n15 VN.n14 161.3
R2146 VN.n13 VN.n12 161.3
R2147 VN.n11 VN.n2 161.3
R2148 VN.n10 VN.n9 161.3
R2149 VN.n8 VN.n3 161.3
R2150 VN.n7 VN.n6 161.3
R2151 VN.n6 VN.n3 54.1398
R2152 VN.n12 VN.n11 54.1398
R2153 VN.n25 VN.n22 54.1398
R2154 VN.n31 VN.n30 54.1398
R2155 VN.n16 VN.n15 48.3272
R2156 VN.n35 VN.n34 48.3272
R2157 VN VN.n37 45.0857
R2158 VN.n26 VN.n23 43.0014
R2159 VN.n7 VN.n4 43.0014
R2160 VN.n5 VN.n4 40.664
R2161 VN.n24 VN.n23 40.664
R2162 VN.n10 VN.n3 27.0143
R2163 VN.n11 VN.n10 27.0143
R2164 VN.n29 VN.n22 27.0143
R2165 VN.n30 VN.n29 27.0143
R2166 VN.n6 VN.n5 13.7719
R2167 VN.n12 VN.n1 13.7719
R2168 VN.n25 VN.n24 13.7719
R2169 VN.n31 VN.n20 13.7719
R2170 VN.n17 VN.n16 12.4157
R2171 VN.n36 VN.n35 12.4157
R2172 VN.n15 VN.n1 10.8209
R2173 VN.n34 VN.n20 10.8209
R2174 VN.n37 VN.n19 0.189894
R2175 VN.n33 VN.n19 0.189894
R2176 VN.n33 VN.n32 0.189894
R2177 VN.n32 VN.n21 0.189894
R2178 VN.n28 VN.n21 0.189894
R2179 VN.n28 VN.n27 0.189894
R2180 VN.n27 VN.n26 0.189894
R2181 VN.n8 VN.n7 0.189894
R2182 VN.n9 VN.n8 0.189894
R2183 VN.n9 VN.n2 0.189894
R2184 VN.n13 VN.n2 0.189894
R2185 VN.n14 VN.n13 0.189894
R2186 VN.n14 VN.n0 0.189894
R2187 VN.n18 VN.n0 0.189894
R2188 VN VN.n18 0.0516364
R2189 VDD2.n141 VDD2.n140 289.615
R2190 VDD2.n68 VDD2.n67 289.615
R2191 VDD2.n140 VDD2.n139 185
R2192 VDD2.n75 VDD2.n74 185
R2193 VDD2.n134 VDD2.n133 185
R2194 VDD2.n132 VDD2.n131 185
R2195 VDD2.n79 VDD2.n78 185
R2196 VDD2.n126 VDD2.n125 185
R2197 VDD2.n124 VDD2.n123 185
R2198 VDD2.n83 VDD2.n82 185
R2199 VDD2.n118 VDD2.n117 185
R2200 VDD2.n116 VDD2.n115 185
R2201 VDD2.n87 VDD2.n86 185
R2202 VDD2.n110 VDD2.n109 185
R2203 VDD2.n108 VDD2.n107 185
R2204 VDD2.n91 VDD2.n90 185
R2205 VDD2.n102 VDD2.n101 185
R2206 VDD2.n100 VDD2.n99 185
R2207 VDD2.n95 VDD2.n94 185
R2208 VDD2.n22 VDD2.n21 185
R2209 VDD2.n27 VDD2.n26 185
R2210 VDD2.n29 VDD2.n28 185
R2211 VDD2.n18 VDD2.n17 185
R2212 VDD2.n35 VDD2.n34 185
R2213 VDD2.n37 VDD2.n36 185
R2214 VDD2.n14 VDD2.n13 185
R2215 VDD2.n43 VDD2.n42 185
R2216 VDD2.n45 VDD2.n44 185
R2217 VDD2.n10 VDD2.n9 185
R2218 VDD2.n51 VDD2.n50 185
R2219 VDD2.n53 VDD2.n52 185
R2220 VDD2.n6 VDD2.n5 185
R2221 VDD2.n59 VDD2.n58 185
R2222 VDD2.n61 VDD2.n60 185
R2223 VDD2.n2 VDD2.n1 185
R2224 VDD2.n67 VDD2.n66 185
R2225 VDD2.n23 VDD2.t6 147.659
R2226 VDD2.n96 VDD2.t1 147.659
R2227 VDD2.n140 VDD2.n74 104.615
R2228 VDD2.n133 VDD2.n74 104.615
R2229 VDD2.n133 VDD2.n132 104.615
R2230 VDD2.n132 VDD2.n78 104.615
R2231 VDD2.n125 VDD2.n78 104.615
R2232 VDD2.n125 VDD2.n124 104.615
R2233 VDD2.n124 VDD2.n82 104.615
R2234 VDD2.n117 VDD2.n82 104.615
R2235 VDD2.n117 VDD2.n116 104.615
R2236 VDD2.n116 VDD2.n86 104.615
R2237 VDD2.n109 VDD2.n86 104.615
R2238 VDD2.n109 VDD2.n108 104.615
R2239 VDD2.n108 VDD2.n90 104.615
R2240 VDD2.n101 VDD2.n90 104.615
R2241 VDD2.n101 VDD2.n100 104.615
R2242 VDD2.n100 VDD2.n94 104.615
R2243 VDD2.n27 VDD2.n21 104.615
R2244 VDD2.n28 VDD2.n27 104.615
R2245 VDD2.n28 VDD2.n17 104.615
R2246 VDD2.n35 VDD2.n17 104.615
R2247 VDD2.n36 VDD2.n35 104.615
R2248 VDD2.n36 VDD2.n13 104.615
R2249 VDD2.n43 VDD2.n13 104.615
R2250 VDD2.n44 VDD2.n43 104.615
R2251 VDD2.n44 VDD2.n9 104.615
R2252 VDD2.n51 VDD2.n9 104.615
R2253 VDD2.n52 VDD2.n51 104.615
R2254 VDD2.n52 VDD2.n5 104.615
R2255 VDD2.n59 VDD2.n5 104.615
R2256 VDD2.n60 VDD2.n59 104.615
R2257 VDD2.n60 VDD2.n1 104.615
R2258 VDD2.n67 VDD2.n1 104.615
R2259 VDD2.n72 VDD2.n71 65.4706
R2260 VDD2 VDD2.n145 65.4677
R2261 VDD2.n144 VDD2.n143 64.6993
R2262 VDD2.n70 VDD2.n69 64.6983
R2263 VDD2.n70 VDD2.n68 53.0706
R2264 VDD2.t1 VDD2.n94 52.3082
R2265 VDD2.t6 VDD2.n21 52.3082
R2266 VDD2.n142 VDD2.n141 51.9672
R2267 VDD2.n142 VDD2.n72 39.8705
R2268 VDD2.n96 VDD2.n95 15.6677
R2269 VDD2.n23 VDD2.n22 15.6677
R2270 VDD2.n139 VDD2.n73 12.8005
R2271 VDD2.n99 VDD2.n98 12.8005
R2272 VDD2.n26 VDD2.n25 12.8005
R2273 VDD2.n66 VDD2.n0 12.8005
R2274 VDD2.n138 VDD2.n75 12.0247
R2275 VDD2.n102 VDD2.n93 12.0247
R2276 VDD2.n29 VDD2.n20 12.0247
R2277 VDD2.n65 VDD2.n2 12.0247
R2278 VDD2.n135 VDD2.n134 11.249
R2279 VDD2.n103 VDD2.n91 11.249
R2280 VDD2.n30 VDD2.n18 11.249
R2281 VDD2.n62 VDD2.n61 11.249
R2282 VDD2.n131 VDD2.n77 10.4732
R2283 VDD2.n107 VDD2.n106 10.4732
R2284 VDD2.n34 VDD2.n33 10.4732
R2285 VDD2.n58 VDD2.n4 10.4732
R2286 VDD2.n130 VDD2.n79 9.69747
R2287 VDD2.n110 VDD2.n89 9.69747
R2288 VDD2.n37 VDD2.n16 9.69747
R2289 VDD2.n57 VDD2.n6 9.69747
R2290 VDD2.n137 VDD2.n73 9.45567
R2291 VDD2.n64 VDD2.n0 9.45567
R2292 VDD2.n122 VDD2.n121 9.3005
R2293 VDD2.n81 VDD2.n80 9.3005
R2294 VDD2.n128 VDD2.n127 9.3005
R2295 VDD2.n130 VDD2.n129 9.3005
R2296 VDD2.n77 VDD2.n76 9.3005
R2297 VDD2.n136 VDD2.n135 9.3005
R2298 VDD2.n138 VDD2.n137 9.3005
R2299 VDD2.n120 VDD2.n119 9.3005
R2300 VDD2.n85 VDD2.n84 9.3005
R2301 VDD2.n114 VDD2.n113 9.3005
R2302 VDD2.n112 VDD2.n111 9.3005
R2303 VDD2.n89 VDD2.n88 9.3005
R2304 VDD2.n106 VDD2.n105 9.3005
R2305 VDD2.n104 VDD2.n103 9.3005
R2306 VDD2.n93 VDD2.n92 9.3005
R2307 VDD2.n98 VDD2.n97 9.3005
R2308 VDD2.n47 VDD2.n46 9.3005
R2309 VDD2.n49 VDD2.n48 9.3005
R2310 VDD2.n8 VDD2.n7 9.3005
R2311 VDD2.n55 VDD2.n54 9.3005
R2312 VDD2.n57 VDD2.n56 9.3005
R2313 VDD2.n4 VDD2.n3 9.3005
R2314 VDD2.n63 VDD2.n62 9.3005
R2315 VDD2.n65 VDD2.n64 9.3005
R2316 VDD2.n41 VDD2.n40 9.3005
R2317 VDD2.n39 VDD2.n38 9.3005
R2318 VDD2.n16 VDD2.n15 9.3005
R2319 VDD2.n33 VDD2.n32 9.3005
R2320 VDD2.n31 VDD2.n30 9.3005
R2321 VDD2.n20 VDD2.n19 9.3005
R2322 VDD2.n25 VDD2.n24 9.3005
R2323 VDD2.n12 VDD2.n11 9.3005
R2324 VDD2.n127 VDD2.n126 8.92171
R2325 VDD2.n111 VDD2.n87 8.92171
R2326 VDD2.n38 VDD2.n14 8.92171
R2327 VDD2.n54 VDD2.n53 8.92171
R2328 VDD2.n123 VDD2.n81 8.14595
R2329 VDD2.n115 VDD2.n114 8.14595
R2330 VDD2.n42 VDD2.n41 8.14595
R2331 VDD2.n50 VDD2.n8 8.14595
R2332 VDD2.n122 VDD2.n83 7.3702
R2333 VDD2.n118 VDD2.n85 7.3702
R2334 VDD2.n45 VDD2.n12 7.3702
R2335 VDD2.n49 VDD2.n10 7.3702
R2336 VDD2.n119 VDD2.n83 6.59444
R2337 VDD2.n119 VDD2.n118 6.59444
R2338 VDD2.n46 VDD2.n45 6.59444
R2339 VDD2.n46 VDD2.n10 6.59444
R2340 VDD2.n123 VDD2.n122 5.81868
R2341 VDD2.n115 VDD2.n85 5.81868
R2342 VDD2.n42 VDD2.n12 5.81868
R2343 VDD2.n50 VDD2.n49 5.81868
R2344 VDD2.n126 VDD2.n81 5.04292
R2345 VDD2.n114 VDD2.n87 5.04292
R2346 VDD2.n41 VDD2.n14 5.04292
R2347 VDD2.n53 VDD2.n8 5.04292
R2348 VDD2.n24 VDD2.n23 4.38563
R2349 VDD2.n97 VDD2.n96 4.38563
R2350 VDD2.n127 VDD2.n79 4.26717
R2351 VDD2.n111 VDD2.n110 4.26717
R2352 VDD2.n38 VDD2.n37 4.26717
R2353 VDD2.n54 VDD2.n6 4.26717
R2354 VDD2.n131 VDD2.n130 3.49141
R2355 VDD2.n107 VDD2.n89 3.49141
R2356 VDD2.n34 VDD2.n16 3.49141
R2357 VDD2.n58 VDD2.n57 3.49141
R2358 VDD2.n134 VDD2.n77 2.71565
R2359 VDD2.n106 VDD2.n91 2.71565
R2360 VDD2.n33 VDD2.n18 2.71565
R2361 VDD2.n61 VDD2.n4 2.71565
R2362 VDD2.n135 VDD2.n75 1.93989
R2363 VDD2.n103 VDD2.n102 1.93989
R2364 VDD2.n30 VDD2.n29 1.93989
R2365 VDD2.n62 VDD2.n2 1.93989
R2366 VDD2.n145 VDD2.t3 1.56448
R2367 VDD2.n145 VDD2.t5 1.56448
R2368 VDD2.n143 VDD2.t4 1.56448
R2369 VDD2.n143 VDD2.t8 1.56448
R2370 VDD2.n71 VDD2.t0 1.56448
R2371 VDD2.n71 VDD2.t2 1.56448
R2372 VDD2.n69 VDD2.t7 1.56448
R2373 VDD2.n69 VDD2.t9 1.56448
R2374 VDD2.n139 VDD2.n138 1.16414
R2375 VDD2.n99 VDD2.n93 1.16414
R2376 VDD2.n26 VDD2.n20 1.16414
R2377 VDD2.n66 VDD2.n65 1.16414
R2378 VDD2.n144 VDD2.n142 1.10395
R2379 VDD2.n141 VDD2.n73 0.388379
R2380 VDD2.n98 VDD2.n95 0.388379
R2381 VDD2.n25 VDD2.n22 0.388379
R2382 VDD2.n68 VDD2.n0 0.388379
R2383 VDD2 VDD2.n144 0.334552
R2384 VDD2.n72 VDD2.n70 0.221016
R2385 VDD2.n137 VDD2.n136 0.155672
R2386 VDD2.n136 VDD2.n76 0.155672
R2387 VDD2.n129 VDD2.n76 0.155672
R2388 VDD2.n129 VDD2.n128 0.155672
R2389 VDD2.n128 VDD2.n80 0.155672
R2390 VDD2.n121 VDD2.n80 0.155672
R2391 VDD2.n121 VDD2.n120 0.155672
R2392 VDD2.n120 VDD2.n84 0.155672
R2393 VDD2.n113 VDD2.n84 0.155672
R2394 VDD2.n113 VDD2.n112 0.155672
R2395 VDD2.n112 VDD2.n88 0.155672
R2396 VDD2.n105 VDD2.n88 0.155672
R2397 VDD2.n105 VDD2.n104 0.155672
R2398 VDD2.n104 VDD2.n92 0.155672
R2399 VDD2.n97 VDD2.n92 0.155672
R2400 VDD2.n24 VDD2.n19 0.155672
R2401 VDD2.n31 VDD2.n19 0.155672
R2402 VDD2.n32 VDD2.n31 0.155672
R2403 VDD2.n32 VDD2.n15 0.155672
R2404 VDD2.n39 VDD2.n15 0.155672
R2405 VDD2.n40 VDD2.n39 0.155672
R2406 VDD2.n40 VDD2.n11 0.155672
R2407 VDD2.n47 VDD2.n11 0.155672
R2408 VDD2.n48 VDD2.n47 0.155672
R2409 VDD2.n48 VDD2.n7 0.155672
R2410 VDD2.n55 VDD2.n7 0.155672
R2411 VDD2.n56 VDD2.n55 0.155672
R2412 VDD2.n56 VDD2.n3 0.155672
R2413 VDD2.n63 VDD2.n3 0.155672
R2414 VDD2.n64 VDD2.n63 0.155672
C0 VP VTAIL 8.1123f
C1 VP VN 6.08096f
C2 VN VTAIL 8.09774f
C3 VP VDD1 8.38896f
C4 VTAIL VDD1 13.0845f
C5 VN VDD1 0.14984f
C6 VP VDD2 0.373707f
C7 VTAIL VDD2 13.1209f
C8 VN VDD2 8.169741f
C9 VDD1 VDD2 1.12929f
C10 VDD2 B 5.372115f
C11 VDD1 B 5.322545f
C12 VTAIL B 7.020792f
C13 VN B 10.60577f
C14 VP B 8.740136f
C15 VDD2.n0 B 0.013192f
C16 VDD2.n1 B 0.029743f
C17 VDD2.n2 B 0.013324f
C18 VDD2.n3 B 0.023418f
C19 VDD2.n4 B 0.012584f
C20 VDD2.n5 B 0.029743f
C21 VDD2.n6 B 0.013324f
C22 VDD2.n7 B 0.023418f
C23 VDD2.n8 B 0.012584f
C24 VDD2.n9 B 0.029743f
C25 VDD2.n10 B 0.013324f
C26 VDD2.n11 B 0.023418f
C27 VDD2.n12 B 0.012584f
C28 VDD2.n13 B 0.029743f
C29 VDD2.n14 B 0.013324f
C30 VDD2.n15 B 0.023418f
C31 VDD2.n16 B 0.012584f
C32 VDD2.n17 B 0.029743f
C33 VDD2.n18 B 0.013324f
C34 VDD2.n19 B 0.023418f
C35 VDD2.n20 B 0.012584f
C36 VDD2.n21 B 0.022307f
C37 VDD2.n22 B 0.01757f
C38 VDD2.t6 B 0.048855f
C39 VDD2.n23 B 0.138996f
C40 VDD2.n24 B 1.27245f
C41 VDD2.n25 B 0.012584f
C42 VDD2.n26 B 0.013324f
C43 VDD2.n27 B 0.029743f
C44 VDD2.n28 B 0.029743f
C45 VDD2.n29 B 0.013324f
C46 VDD2.n30 B 0.012584f
C47 VDD2.n31 B 0.023418f
C48 VDD2.n32 B 0.023418f
C49 VDD2.n33 B 0.012584f
C50 VDD2.n34 B 0.013324f
C51 VDD2.n35 B 0.029743f
C52 VDD2.n36 B 0.029743f
C53 VDD2.n37 B 0.013324f
C54 VDD2.n38 B 0.012584f
C55 VDD2.n39 B 0.023418f
C56 VDD2.n40 B 0.023418f
C57 VDD2.n41 B 0.012584f
C58 VDD2.n42 B 0.013324f
C59 VDD2.n43 B 0.029743f
C60 VDD2.n44 B 0.029743f
C61 VDD2.n45 B 0.013324f
C62 VDD2.n46 B 0.012584f
C63 VDD2.n47 B 0.023418f
C64 VDD2.n48 B 0.023418f
C65 VDD2.n49 B 0.012584f
C66 VDD2.n50 B 0.013324f
C67 VDD2.n51 B 0.029743f
C68 VDD2.n52 B 0.029743f
C69 VDD2.n53 B 0.013324f
C70 VDD2.n54 B 0.012584f
C71 VDD2.n55 B 0.023418f
C72 VDD2.n56 B 0.023418f
C73 VDD2.n57 B 0.012584f
C74 VDD2.n58 B 0.013324f
C75 VDD2.n59 B 0.029743f
C76 VDD2.n60 B 0.029743f
C77 VDD2.n61 B 0.013324f
C78 VDD2.n62 B 0.012584f
C79 VDD2.n63 B 0.023418f
C80 VDD2.n64 B 0.059887f
C81 VDD2.n65 B 0.012584f
C82 VDD2.n66 B 0.013324f
C83 VDD2.n67 B 0.060477f
C84 VDD2.n68 B 0.069603f
C85 VDD2.t7 B 0.234277f
C86 VDD2.t9 B 0.234277f
C87 VDD2.n69 B 2.1032f
C88 VDD2.n70 B 0.416487f
C89 VDD2.t0 B 0.234277f
C90 VDD2.t2 B 0.234277f
C91 VDD2.n71 B 2.10718f
C92 VDD2.n72 B 1.93852f
C93 VDD2.n73 B 0.013192f
C94 VDD2.n74 B 0.029743f
C95 VDD2.n75 B 0.013324f
C96 VDD2.n76 B 0.023418f
C97 VDD2.n77 B 0.012584f
C98 VDD2.n78 B 0.029743f
C99 VDD2.n79 B 0.013324f
C100 VDD2.n80 B 0.023418f
C101 VDD2.n81 B 0.012584f
C102 VDD2.n82 B 0.029743f
C103 VDD2.n83 B 0.013324f
C104 VDD2.n84 B 0.023418f
C105 VDD2.n85 B 0.012584f
C106 VDD2.n86 B 0.029743f
C107 VDD2.n87 B 0.013324f
C108 VDD2.n88 B 0.023418f
C109 VDD2.n89 B 0.012584f
C110 VDD2.n90 B 0.029743f
C111 VDD2.n91 B 0.013324f
C112 VDD2.n92 B 0.023418f
C113 VDD2.n93 B 0.012584f
C114 VDD2.n94 B 0.022307f
C115 VDD2.n95 B 0.01757f
C116 VDD2.t1 B 0.048855f
C117 VDD2.n96 B 0.138996f
C118 VDD2.n97 B 1.27245f
C119 VDD2.n98 B 0.012584f
C120 VDD2.n99 B 0.013324f
C121 VDD2.n100 B 0.029743f
C122 VDD2.n101 B 0.029743f
C123 VDD2.n102 B 0.013324f
C124 VDD2.n103 B 0.012584f
C125 VDD2.n104 B 0.023418f
C126 VDD2.n105 B 0.023418f
C127 VDD2.n106 B 0.012584f
C128 VDD2.n107 B 0.013324f
C129 VDD2.n108 B 0.029743f
C130 VDD2.n109 B 0.029743f
C131 VDD2.n110 B 0.013324f
C132 VDD2.n111 B 0.012584f
C133 VDD2.n112 B 0.023418f
C134 VDD2.n113 B 0.023418f
C135 VDD2.n114 B 0.012584f
C136 VDD2.n115 B 0.013324f
C137 VDD2.n116 B 0.029743f
C138 VDD2.n117 B 0.029743f
C139 VDD2.n118 B 0.013324f
C140 VDD2.n119 B 0.012584f
C141 VDD2.n120 B 0.023418f
C142 VDD2.n121 B 0.023418f
C143 VDD2.n122 B 0.012584f
C144 VDD2.n123 B 0.013324f
C145 VDD2.n124 B 0.029743f
C146 VDD2.n125 B 0.029743f
C147 VDD2.n126 B 0.013324f
C148 VDD2.n127 B 0.012584f
C149 VDD2.n128 B 0.023418f
C150 VDD2.n129 B 0.023418f
C151 VDD2.n130 B 0.012584f
C152 VDD2.n131 B 0.013324f
C153 VDD2.n132 B 0.029743f
C154 VDD2.n133 B 0.029743f
C155 VDD2.n134 B 0.013324f
C156 VDD2.n135 B 0.012584f
C157 VDD2.n136 B 0.023418f
C158 VDD2.n137 B 0.059887f
C159 VDD2.n138 B 0.012584f
C160 VDD2.n139 B 0.013324f
C161 VDD2.n140 B 0.060477f
C162 VDD2.n141 B 0.066873f
C163 VDD2.n142 B 2.15942f
C164 VDD2.t4 B 0.234277f
C165 VDD2.t8 B 0.234277f
C166 VDD2.n143 B 2.1032f
C167 VDD2.n144 B 0.294041f
C168 VDD2.t3 B 0.234277f
C169 VDD2.t5 B 0.234277f
C170 VDD2.n145 B 2.10715f
C171 VN.n0 B 0.037748f
C172 VN.t9 B 1.2388f
C173 VN.n1 B 0.458657f
C174 VN.n2 B 0.037748f
C175 VN.t0 B 1.2388f
C176 VN.n3 B 0.041106f
C177 VN.t3 B 1.32073f
C178 VN.n4 B 0.504187f
C179 VN.t2 B 1.2388f
C180 VN.n5 B 0.497257f
C181 VN.n6 B 0.050645f
C182 VN.n7 B 0.163425f
C183 VN.n8 B 0.037748f
C184 VN.n9 B 0.037748f
C185 VN.n10 B 0.499676f
C186 VN.n11 B 0.041106f
C187 VN.n12 B 0.050645f
C188 VN.n13 B 0.037748f
C189 VN.n14 B 0.037748f
C190 VN.n15 B 0.050987f
C191 VN.n16 B 0.014619f
C192 VN.t7 B 1.2934f
C193 VN.n17 B 0.503676f
C194 VN.n18 B 0.029253f
C195 VN.n19 B 0.037748f
C196 VN.t5 B 1.2388f
C197 VN.n20 B 0.458657f
C198 VN.n21 B 0.037748f
C199 VN.t1 B 1.2388f
C200 VN.n22 B 0.041106f
C201 VN.t4 B 1.32073f
C202 VN.n23 B 0.504187f
C203 VN.t6 B 1.2388f
C204 VN.n24 B 0.497257f
C205 VN.n25 B 0.050645f
C206 VN.n26 B 0.163425f
C207 VN.n27 B 0.037748f
C208 VN.n28 B 0.037748f
C209 VN.n29 B 0.499676f
C210 VN.n30 B 0.041106f
C211 VN.n31 B 0.050645f
C212 VN.n32 B 0.037748f
C213 VN.n33 B 0.037748f
C214 VN.n34 B 0.050987f
C215 VN.n35 B 0.014619f
C216 VN.t8 B 1.2934f
C217 VN.n36 B 0.503676f
C218 VN.n37 B 1.74993f
C219 VDD1.n0 B 0.013262f
C220 VDD1.n1 B 0.029901f
C221 VDD1.n2 B 0.013395f
C222 VDD1.n3 B 0.023542f
C223 VDD1.n4 B 0.01265f
C224 VDD1.n5 B 0.029901f
C225 VDD1.n6 B 0.013395f
C226 VDD1.n7 B 0.023542f
C227 VDD1.n8 B 0.01265f
C228 VDD1.n9 B 0.029901f
C229 VDD1.n10 B 0.013395f
C230 VDD1.n11 B 0.023542f
C231 VDD1.n12 B 0.01265f
C232 VDD1.n13 B 0.029901f
C233 VDD1.n14 B 0.013395f
C234 VDD1.n15 B 0.023542f
C235 VDD1.n16 B 0.01265f
C236 VDD1.n17 B 0.029901f
C237 VDD1.n18 B 0.013395f
C238 VDD1.n19 B 0.023542f
C239 VDD1.n20 B 0.01265f
C240 VDD1.n21 B 0.022426f
C241 VDD1.n22 B 0.017663f
C242 VDD1.t8 B 0.049114f
C243 VDD1.n23 B 0.139734f
C244 VDD1.n24 B 1.2792f
C245 VDD1.n25 B 0.01265f
C246 VDD1.n26 B 0.013395f
C247 VDD1.n27 B 0.029901f
C248 VDD1.n28 B 0.029901f
C249 VDD1.n29 B 0.013395f
C250 VDD1.n30 B 0.01265f
C251 VDD1.n31 B 0.023542f
C252 VDD1.n32 B 0.023542f
C253 VDD1.n33 B 0.01265f
C254 VDD1.n34 B 0.013395f
C255 VDD1.n35 B 0.029901f
C256 VDD1.n36 B 0.029901f
C257 VDD1.n37 B 0.013395f
C258 VDD1.n38 B 0.01265f
C259 VDD1.n39 B 0.023542f
C260 VDD1.n40 B 0.023542f
C261 VDD1.n41 B 0.01265f
C262 VDD1.n42 B 0.013395f
C263 VDD1.n43 B 0.029901f
C264 VDD1.n44 B 0.029901f
C265 VDD1.n45 B 0.013395f
C266 VDD1.n46 B 0.01265f
C267 VDD1.n47 B 0.023542f
C268 VDD1.n48 B 0.023542f
C269 VDD1.n49 B 0.01265f
C270 VDD1.n50 B 0.013395f
C271 VDD1.n51 B 0.029901f
C272 VDD1.n52 B 0.029901f
C273 VDD1.n53 B 0.013395f
C274 VDD1.n54 B 0.01265f
C275 VDD1.n55 B 0.023542f
C276 VDD1.n56 B 0.023542f
C277 VDD1.n57 B 0.01265f
C278 VDD1.n58 B 0.013395f
C279 VDD1.n59 B 0.029901f
C280 VDD1.n60 B 0.029901f
C281 VDD1.n61 B 0.013395f
C282 VDD1.n62 B 0.01265f
C283 VDD1.n63 B 0.023542f
C284 VDD1.n64 B 0.060205f
C285 VDD1.n65 B 0.01265f
C286 VDD1.n66 B 0.013395f
C287 VDD1.n67 B 0.060798f
C288 VDD1.n68 B 0.069972f
C289 VDD1.t5 B 0.23552f
C290 VDD1.t3 B 0.23552f
C291 VDD1.n69 B 2.11436f
C292 VDD1.n70 B 0.42484f
C293 VDD1.n71 B 0.013262f
C294 VDD1.n72 B 0.029901f
C295 VDD1.n73 B 0.013395f
C296 VDD1.n74 B 0.023542f
C297 VDD1.n75 B 0.01265f
C298 VDD1.n76 B 0.029901f
C299 VDD1.n77 B 0.013395f
C300 VDD1.n78 B 0.023542f
C301 VDD1.n79 B 0.01265f
C302 VDD1.n80 B 0.029901f
C303 VDD1.n81 B 0.013395f
C304 VDD1.n82 B 0.023542f
C305 VDD1.n83 B 0.01265f
C306 VDD1.n84 B 0.029901f
C307 VDD1.n85 B 0.013395f
C308 VDD1.n86 B 0.023542f
C309 VDD1.n87 B 0.01265f
C310 VDD1.n88 B 0.029901f
C311 VDD1.n89 B 0.013395f
C312 VDD1.n90 B 0.023542f
C313 VDD1.n91 B 0.01265f
C314 VDD1.n92 B 0.022426f
C315 VDD1.n93 B 0.017663f
C316 VDD1.t6 B 0.049114f
C317 VDD1.n94 B 0.139733f
C318 VDD1.n95 B 1.2792f
C319 VDD1.n96 B 0.01265f
C320 VDD1.n97 B 0.013395f
C321 VDD1.n98 B 0.029901f
C322 VDD1.n99 B 0.029901f
C323 VDD1.n100 B 0.013395f
C324 VDD1.n101 B 0.01265f
C325 VDD1.n102 B 0.023542f
C326 VDD1.n103 B 0.023542f
C327 VDD1.n104 B 0.01265f
C328 VDD1.n105 B 0.013395f
C329 VDD1.n106 B 0.029901f
C330 VDD1.n107 B 0.029901f
C331 VDD1.n108 B 0.013395f
C332 VDD1.n109 B 0.01265f
C333 VDD1.n110 B 0.023542f
C334 VDD1.n111 B 0.023542f
C335 VDD1.n112 B 0.01265f
C336 VDD1.n113 B 0.013395f
C337 VDD1.n114 B 0.029901f
C338 VDD1.n115 B 0.029901f
C339 VDD1.n116 B 0.013395f
C340 VDD1.n117 B 0.01265f
C341 VDD1.n118 B 0.023542f
C342 VDD1.n119 B 0.023542f
C343 VDD1.n120 B 0.01265f
C344 VDD1.n121 B 0.013395f
C345 VDD1.n122 B 0.029901f
C346 VDD1.n123 B 0.029901f
C347 VDD1.n124 B 0.013395f
C348 VDD1.n125 B 0.01265f
C349 VDD1.n126 B 0.023542f
C350 VDD1.n127 B 0.023542f
C351 VDD1.n128 B 0.01265f
C352 VDD1.n129 B 0.013395f
C353 VDD1.n130 B 0.029901f
C354 VDD1.n131 B 0.029901f
C355 VDD1.n132 B 0.013395f
C356 VDD1.n133 B 0.01265f
C357 VDD1.n134 B 0.023542f
C358 VDD1.n135 B 0.060205f
C359 VDD1.n136 B 0.01265f
C360 VDD1.n137 B 0.013395f
C361 VDD1.n138 B 0.060798f
C362 VDD1.n139 B 0.069972f
C363 VDD1.t4 B 0.23552f
C364 VDD1.t2 B 0.23552f
C365 VDD1.n140 B 2.11436f
C366 VDD1.n141 B 0.418698f
C367 VDD1.t0 B 0.23552f
C368 VDD1.t9 B 0.23552f
C369 VDD1.n142 B 2.11836f
C370 VDD1.n143 B 2.02713f
C371 VDD1.t1 B 0.23552f
C372 VDD1.t7 B 0.23552f
C373 VDD1.n144 B 2.11436f
C374 VDD1.n145 B 2.38564f
C375 VTAIL.t7 B 0.247751f
C376 VTAIL.t5 B 0.247751f
C377 VTAIL.n0 B 2.15764f
C378 VTAIL.n1 B 0.381301f
C379 VTAIL.n2 B 0.013951f
C380 VTAIL.n3 B 0.031454f
C381 VTAIL.n4 B 0.01409f
C382 VTAIL.n5 B 0.024764f
C383 VTAIL.n6 B 0.013307f
C384 VTAIL.n7 B 0.031454f
C385 VTAIL.n8 B 0.01409f
C386 VTAIL.n9 B 0.024764f
C387 VTAIL.n10 B 0.013307f
C388 VTAIL.n11 B 0.031454f
C389 VTAIL.n12 B 0.01409f
C390 VTAIL.n13 B 0.024764f
C391 VTAIL.n14 B 0.013307f
C392 VTAIL.n15 B 0.031454f
C393 VTAIL.n16 B 0.01409f
C394 VTAIL.n17 B 0.024764f
C395 VTAIL.n18 B 0.013307f
C396 VTAIL.n19 B 0.031454f
C397 VTAIL.n20 B 0.01409f
C398 VTAIL.n21 B 0.024764f
C399 VTAIL.n22 B 0.013307f
C400 VTAIL.n23 B 0.02359f
C401 VTAIL.n24 B 0.018581f
C402 VTAIL.t18 B 0.051665f
C403 VTAIL.n25 B 0.14699f
C404 VTAIL.n26 B 1.34563f
C405 VTAIL.n27 B 0.013307f
C406 VTAIL.n28 B 0.01409f
C407 VTAIL.n29 B 0.031454f
C408 VTAIL.n30 B 0.031454f
C409 VTAIL.n31 B 0.01409f
C410 VTAIL.n32 B 0.013307f
C411 VTAIL.n33 B 0.024764f
C412 VTAIL.n34 B 0.024764f
C413 VTAIL.n35 B 0.013307f
C414 VTAIL.n36 B 0.01409f
C415 VTAIL.n37 B 0.031454f
C416 VTAIL.n38 B 0.031454f
C417 VTAIL.n39 B 0.01409f
C418 VTAIL.n40 B 0.013307f
C419 VTAIL.n41 B 0.024764f
C420 VTAIL.n42 B 0.024764f
C421 VTAIL.n43 B 0.013307f
C422 VTAIL.n44 B 0.01409f
C423 VTAIL.n45 B 0.031454f
C424 VTAIL.n46 B 0.031454f
C425 VTAIL.n47 B 0.01409f
C426 VTAIL.n48 B 0.013307f
C427 VTAIL.n49 B 0.024764f
C428 VTAIL.n50 B 0.024764f
C429 VTAIL.n51 B 0.013307f
C430 VTAIL.n52 B 0.01409f
C431 VTAIL.n53 B 0.031454f
C432 VTAIL.n54 B 0.031454f
C433 VTAIL.n55 B 0.01409f
C434 VTAIL.n56 B 0.013307f
C435 VTAIL.n57 B 0.024764f
C436 VTAIL.n58 B 0.024764f
C437 VTAIL.n59 B 0.013307f
C438 VTAIL.n60 B 0.01409f
C439 VTAIL.n61 B 0.031454f
C440 VTAIL.n62 B 0.031454f
C441 VTAIL.n63 B 0.01409f
C442 VTAIL.n64 B 0.013307f
C443 VTAIL.n65 B 0.024764f
C444 VTAIL.n66 B 0.063331f
C445 VTAIL.n67 B 0.013307f
C446 VTAIL.n68 B 0.01409f
C447 VTAIL.n69 B 0.063955f
C448 VTAIL.n70 B 0.053659f
C449 VTAIL.n71 B 0.19378f
C450 VTAIL.t12 B 0.247751f
C451 VTAIL.t15 B 0.247751f
C452 VTAIL.n72 B 2.15764f
C453 VTAIL.n73 B 0.405206f
C454 VTAIL.t9 B 0.247751f
C455 VTAIL.t11 B 0.247751f
C456 VTAIL.n74 B 2.15764f
C457 VTAIL.n75 B 1.70054f
C458 VTAIL.t0 B 0.247751f
C459 VTAIL.t19 B 0.247751f
C460 VTAIL.n76 B 2.15764f
C461 VTAIL.n77 B 1.70054f
C462 VTAIL.t4 B 0.247751f
C463 VTAIL.t2 B 0.247751f
C464 VTAIL.n78 B 2.15764f
C465 VTAIL.n79 B 0.405211f
C466 VTAIL.n80 B 0.013951f
C467 VTAIL.n81 B 0.031454f
C468 VTAIL.n82 B 0.01409f
C469 VTAIL.n83 B 0.024764f
C470 VTAIL.n84 B 0.013307f
C471 VTAIL.n85 B 0.031454f
C472 VTAIL.n86 B 0.01409f
C473 VTAIL.n87 B 0.024764f
C474 VTAIL.n88 B 0.013307f
C475 VTAIL.n89 B 0.031454f
C476 VTAIL.n90 B 0.01409f
C477 VTAIL.n91 B 0.024764f
C478 VTAIL.n92 B 0.013307f
C479 VTAIL.n93 B 0.031454f
C480 VTAIL.n94 B 0.01409f
C481 VTAIL.n95 B 0.024764f
C482 VTAIL.n96 B 0.013307f
C483 VTAIL.n97 B 0.031454f
C484 VTAIL.n98 B 0.01409f
C485 VTAIL.n99 B 0.024764f
C486 VTAIL.n100 B 0.013307f
C487 VTAIL.n101 B 0.02359f
C488 VTAIL.n102 B 0.018581f
C489 VTAIL.t3 B 0.051665f
C490 VTAIL.n103 B 0.14699f
C491 VTAIL.n104 B 1.34563f
C492 VTAIL.n105 B 0.013307f
C493 VTAIL.n106 B 0.01409f
C494 VTAIL.n107 B 0.031454f
C495 VTAIL.n108 B 0.031454f
C496 VTAIL.n109 B 0.01409f
C497 VTAIL.n110 B 0.013307f
C498 VTAIL.n111 B 0.024764f
C499 VTAIL.n112 B 0.024764f
C500 VTAIL.n113 B 0.013307f
C501 VTAIL.n114 B 0.01409f
C502 VTAIL.n115 B 0.031454f
C503 VTAIL.n116 B 0.031454f
C504 VTAIL.n117 B 0.01409f
C505 VTAIL.n118 B 0.013307f
C506 VTAIL.n119 B 0.024764f
C507 VTAIL.n120 B 0.024764f
C508 VTAIL.n121 B 0.013307f
C509 VTAIL.n122 B 0.01409f
C510 VTAIL.n123 B 0.031454f
C511 VTAIL.n124 B 0.031454f
C512 VTAIL.n125 B 0.01409f
C513 VTAIL.n126 B 0.013307f
C514 VTAIL.n127 B 0.024764f
C515 VTAIL.n128 B 0.024764f
C516 VTAIL.n129 B 0.013307f
C517 VTAIL.n130 B 0.01409f
C518 VTAIL.n131 B 0.031454f
C519 VTAIL.n132 B 0.031454f
C520 VTAIL.n133 B 0.01409f
C521 VTAIL.n134 B 0.013307f
C522 VTAIL.n135 B 0.024764f
C523 VTAIL.n136 B 0.024764f
C524 VTAIL.n137 B 0.013307f
C525 VTAIL.n138 B 0.01409f
C526 VTAIL.n139 B 0.031454f
C527 VTAIL.n140 B 0.031454f
C528 VTAIL.n141 B 0.01409f
C529 VTAIL.n142 B 0.013307f
C530 VTAIL.n143 B 0.024764f
C531 VTAIL.n144 B 0.063331f
C532 VTAIL.n145 B 0.013307f
C533 VTAIL.n146 B 0.01409f
C534 VTAIL.n147 B 0.063955f
C535 VTAIL.n148 B 0.053659f
C536 VTAIL.n149 B 0.19378f
C537 VTAIL.t13 B 0.247751f
C538 VTAIL.t17 B 0.247751f
C539 VTAIL.n150 B 2.15764f
C540 VTAIL.n151 B 0.398676f
C541 VTAIL.t10 B 0.247751f
C542 VTAIL.t14 B 0.247751f
C543 VTAIL.n152 B 2.15764f
C544 VTAIL.n153 B 0.405211f
C545 VTAIL.n154 B 0.013951f
C546 VTAIL.n155 B 0.031454f
C547 VTAIL.n156 B 0.01409f
C548 VTAIL.n157 B 0.024764f
C549 VTAIL.n158 B 0.013307f
C550 VTAIL.n159 B 0.031454f
C551 VTAIL.n160 B 0.01409f
C552 VTAIL.n161 B 0.024764f
C553 VTAIL.n162 B 0.013307f
C554 VTAIL.n163 B 0.031454f
C555 VTAIL.n164 B 0.01409f
C556 VTAIL.n165 B 0.024764f
C557 VTAIL.n166 B 0.013307f
C558 VTAIL.n167 B 0.031454f
C559 VTAIL.n168 B 0.01409f
C560 VTAIL.n169 B 0.024764f
C561 VTAIL.n170 B 0.013307f
C562 VTAIL.n171 B 0.031454f
C563 VTAIL.n172 B 0.01409f
C564 VTAIL.n173 B 0.024764f
C565 VTAIL.n174 B 0.013307f
C566 VTAIL.n175 B 0.02359f
C567 VTAIL.n176 B 0.018581f
C568 VTAIL.t16 B 0.051665f
C569 VTAIL.n177 B 0.14699f
C570 VTAIL.n178 B 1.34563f
C571 VTAIL.n179 B 0.013307f
C572 VTAIL.n180 B 0.01409f
C573 VTAIL.n181 B 0.031454f
C574 VTAIL.n182 B 0.031454f
C575 VTAIL.n183 B 0.01409f
C576 VTAIL.n184 B 0.013307f
C577 VTAIL.n185 B 0.024764f
C578 VTAIL.n186 B 0.024764f
C579 VTAIL.n187 B 0.013307f
C580 VTAIL.n188 B 0.01409f
C581 VTAIL.n189 B 0.031454f
C582 VTAIL.n190 B 0.031454f
C583 VTAIL.n191 B 0.01409f
C584 VTAIL.n192 B 0.013307f
C585 VTAIL.n193 B 0.024764f
C586 VTAIL.n194 B 0.024764f
C587 VTAIL.n195 B 0.013307f
C588 VTAIL.n196 B 0.01409f
C589 VTAIL.n197 B 0.031454f
C590 VTAIL.n198 B 0.031454f
C591 VTAIL.n199 B 0.01409f
C592 VTAIL.n200 B 0.013307f
C593 VTAIL.n201 B 0.024764f
C594 VTAIL.n202 B 0.024764f
C595 VTAIL.n203 B 0.013307f
C596 VTAIL.n204 B 0.01409f
C597 VTAIL.n205 B 0.031454f
C598 VTAIL.n206 B 0.031454f
C599 VTAIL.n207 B 0.01409f
C600 VTAIL.n208 B 0.013307f
C601 VTAIL.n209 B 0.024764f
C602 VTAIL.n210 B 0.024764f
C603 VTAIL.n211 B 0.013307f
C604 VTAIL.n212 B 0.01409f
C605 VTAIL.n213 B 0.031454f
C606 VTAIL.n214 B 0.031454f
C607 VTAIL.n215 B 0.01409f
C608 VTAIL.n216 B 0.013307f
C609 VTAIL.n217 B 0.024764f
C610 VTAIL.n218 B 0.063331f
C611 VTAIL.n219 B 0.013307f
C612 VTAIL.n220 B 0.01409f
C613 VTAIL.n221 B 0.063955f
C614 VTAIL.n222 B 0.053659f
C615 VTAIL.n223 B 1.40759f
C616 VTAIL.n224 B 0.013951f
C617 VTAIL.n225 B 0.031454f
C618 VTAIL.n226 B 0.01409f
C619 VTAIL.n227 B 0.024764f
C620 VTAIL.n228 B 0.013307f
C621 VTAIL.n229 B 0.031454f
C622 VTAIL.n230 B 0.01409f
C623 VTAIL.n231 B 0.024764f
C624 VTAIL.n232 B 0.013307f
C625 VTAIL.n233 B 0.031454f
C626 VTAIL.n234 B 0.01409f
C627 VTAIL.n235 B 0.024764f
C628 VTAIL.n236 B 0.013307f
C629 VTAIL.n237 B 0.031454f
C630 VTAIL.n238 B 0.01409f
C631 VTAIL.n239 B 0.024764f
C632 VTAIL.n240 B 0.013307f
C633 VTAIL.n241 B 0.031454f
C634 VTAIL.n242 B 0.01409f
C635 VTAIL.n243 B 0.024764f
C636 VTAIL.n244 B 0.013307f
C637 VTAIL.n245 B 0.02359f
C638 VTAIL.n246 B 0.018581f
C639 VTAIL.t6 B 0.051665f
C640 VTAIL.n247 B 0.14699f
C641 VTAIL.n248 B 1.34563f
C642 VTAIL.n249 B 0.013307f
C643 VTAIL.n250 B 0.01409f
C644 VTAIL.n251 B 0.031454f
C645 VTAIL.n252 B 0.031454f
C646 VTAIL.n253 B 0.01409f
C647 VTAIL.n254 B 0.013307f
C648 VTAIL.n255 B 0.024764f
C649 VTAIL.n256 B 0.024764f
C650 VTAIL.n257 B 0.013307f
C651 VTAIL.n258 B 0.01409f
C652 VTAIL.n259 B 0.031454f
C653 VTAIL.n260 B 0.031454f
C654 VTAIL.n261 B 0.01409f
C655 VTAIL.n262 B 0.013307f
C656 VTAIL.n263 B 0.024764f
C657 VTAIL.n264 B 0.024764f
C658 VTAIL.n265 B 0.013307f
C659 VTAIL.n266 B 0.01409f
C660 VTAIL.n267 B 0.031454f
C661 VTAIL.n268 B 0.031454f
C662 VTAIL.n269 B 0.01409f
C663 VTAIL.n270 B 0.013307f
C664 VTAIL.n271 B 0.024764f
C665 VTAIL.n272 B 0.024764f
C666 VTAIL.n273 B 0.013307f
C667 VTAIL.n274 B 0.01409f
C668 VTAIL.n275 B 0.031454f
C669 VTAIL.n276 B 0.031454f
C670 VTAIL.n277 B 0.01409f
C671 VTAIL.n278 B 0.013307f
C672 VTAIL.n279 B 0.024764f
C673 VTAIL.n280 B 0.024764f
C674 VTAIL.n281 B 0.013307f
C675 VTAIL.n282 B 0.01409f
C676 VTAIL.n283 B 0.031454f
C677 VTAIL.n284 B 0.031454f
C678 VTAIL.n285 B 0.01409f
C679 VTAIL.n286 B 0.013307f
C680 VTAIL.n287 B 0.024764f
C681 VTAIL.n288 B 0.063331f
C682 VTAIL.n289 B 0.013307f
C683 VTAIL.n290 B 0.01409f
C684 VTAIL.n291 B 0.063955f
C685 VTAIL.n292 B 0.053659f
C686 VTAIL.n293 B 1.40759f
C687 VTAIL.t8 B 0.247751f
C688 VTAIL.t1 B 0.247751f
C689 VTAIL.n294 B 2.15764f
C690 VTAIL.n295 B 0.334524f
C691 VP.n0 B 0.038175f
C692 VP.t9 B 1.25283f
C693 VP.n1 B 0.463851f
C694 VP.n2 B 0.038175f
C695 VP.t7 B 1.25283f
C696 VP.n3 B 0.041571f
C697 VP.n4 B 0.038175f
C698 VP.t5 B 1.25283f
C699 VP.t3 B 1.30805f
C700 VP.n5 B 0.50938f
C701 VP.n6 B 0.038175f
C702 VP.t2 B 1.30805f
C703 VP.t8 B 1.25283f
C704 VP.n7 B 0.463851f
C705 VP.n8 B 0.038175f
C706 VP.t6 B 1.25283f
C707 VP.n9 B 0.041571f
C708 VP.t1 B 1.33569f
C709 VP.n10 B 0.509896f
C710 VP.t4 B 1.25283f
C711 VP.n11 B 0.502888f
C712 VP.n12 B 0.051219f
C713 VP.n13 B 0.165276f
C714 VP.n14 B 0.038175f
C715 VP.n15 B 0.038175f
C716 VP.n16 B 0.505335f
C717 VP.n17 B 0.041571f
C718 VP.n18 B 0.051219f
C719 VP.n19 B 0.038175f
C720 VP.n20 B 0.038175f
C721 VP.n21 B 0.051565f
C722 VP.n22 B 0.014785f
C723 VP.n23 B 0.50938f
C724 VP.n24 B 1.74478f
C725 VP.n25 B 1.77557f
C726 VP.n26 B 0.038175f
C727 VP.n27 B 0.014785f
C728 VP.n28 B 0.051565f
C729 VP.n29 B 0.463851f
C730 VP.n30 B 0.051219f
C731 VP.n31 B 0.038175f
C732 VP.n32 B 0.038175f
C733 VP.n33 B 0.038175f
C734 VP.n34 B 0.505335f
C735 VP.n35 B 0.041571f
C736 VP.n36 B 0.051219f
C737 VP.n37 B 0.038175f
C738 VP.n38 B 0.038175f
C739 VP.n39 B 0.051565f
C740 VP.n40 B 0.014785f
C741 VP.t0 B 1.30805f
C742 VP.n41 B 0.50938f
C743 VP.n42 B 0.029584f
.ends

