* NGSPICE file created from diff_pair_sample_1465.ext - technology: sky130A

.subckt diff_pair_sample_1465 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X1 VTAIL.t12 VN.t1 VDD2.t6 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X2 B.t11 B.t9 B.t10 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=0 ps=0 w=17.37 l=1.13
X3 VTAIL.t8 VN.t2 VDD2.t5 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X4 VTAIL.t7 VP.t0 VDD1.t7 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X5 VTAIL.t5 VP.t1 VDD1.t6 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=2.86605 ps=17.7 w=17.37 l=1.13
X6 VDD1.t5 VP.t2 VTAIL.t6 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=6.7743 ps=35.52 w=17.37 l=1.13
X7 VDD2.t4 VN.t3 VTAIL.t9 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=6.7743 ps=35.52 w=17.37 l=1.13
X8 B.t8 B.t6 B.t7 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=0 ps=0 w=17.37 l=1.13
X9 VDD2.t3 VN.t4 VTAIL.t14 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=6.7743 ps=35.52 w=17.37 l=1.13
X10 VDD1.t4 VP.t3 VTAIL.t0 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X11 VTAIL.t2 VP.t4 VDD1.t3 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X12 VTAIL.t13 VN.t5 VDD2.t2 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=2.86605 ps=17.7 w=17.37 l=1.13
X13 VTAIL.t10 VN.t6 VDD2.t1 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=2.86605 ps=17.7 w=17.37 l=1.13
X14 VTAIL.t4 VP.t5 VDD1.t2 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=2.86605 ps=17.7 w=17.37 l=1.13
X15 VDD2.t0 VN.t7 VTAIL.t15 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
X16 B.t5 B.t3 B.t4 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=0 ps=0 w=17.37 l=1.13
X17 VDD1.t1 VP.t6 VTAIL.t1 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=6.7743 ps=35.52 w=17.37 l=1.13
X18 B.t2 B.t0 B.t1 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=6.7743 pd=35.52 as=0 ps=0 w=17.37 l=1.13
X19 VDD1.t0 VP.t7 VTAIL.t3 w_n2430_n4442# sky130_fd_pr__pfet_01v8 ad=2.86605 pd=17.7 as=2.86605 ps=17.7 w=17.37 l=1.13
R0 VN.n3 VN.t6 428.428
R1 VN.n16 VN.t3 428.428
R2 VN.n11 VN.t4 405.435
R3 VN.n24 VN.t5 405.435
R4 VN.n4 VN.t0 370.459
R5 VN.n1 VN.t2 370.459
R6 VN.n17 VN.t1 370.459
R7 VN.n14 VN.t7 370.459
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN.n11 VN.n10 50.4025
R21 VN.n24 VN.n23 50.4025
R22 VN VN.n25 48.5748
R23 VN.n4 VN.n3 33.6057
R24 VN.n17 VN.n16 33.6057
R25 VN.n16 VN.n15 28.1515
R26 VN.n3 VN.n2 28.1515
R27 VN.n10 VN.n9 24.4675
R28 VN.n23 VN.n22 24.4675
R29 VN.n5 VN.n4 23.4888
R30 VN.n6 VN.n1 23.4888
R31 VN.n18 VN.n17 23.4888
R32 VN.n19 VN.n14 23.4888
R33 VN.n9 VN.n1 0.97918
R34 VN.n22 VN.n14 0.97918
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VTAIL.n774 VTAIL.n773 756.745
R45 VTAIL.n96 VTAIL.n95 756.745
R46 VTAIL.n192 VTAIL.n191 756.745
R47 VTAIL.n290 VTAIL.n289 756.745
R48 VTAIL.n678 VTAIL.n677 756.745
R49 VTAIL.n580 VTAIL.n579 756.745
R50 VTAIL.n484 VTAIL.n483 756.745
R51 VTAIL.n386 VTAIL.n385 756.745
R52 VTAIL.n710 VTAIL.n709 585
R53 VTAIL.n715 VTAIL.n714 585
R54 VTAIL.n717 VTAIL.n716 585
R55 VTAIL.n706 VTAIL.n705 585
R56 VTAIL.n723 VTAIL.n722 585
R57 VTAIL.n725 VTAIL.n724 585
R58 VTAIL.n702 VTAIL.n701 585
R59 VTAIL.n732 VTAIL.n731 585
R60 VTAIL.n733 VTAIL.n700 585
R61 VTAIL.n735 VTAIL.n734 585
R62 VTAIL.n698 VTAIL.n697 585
R63 VTAIL.n741 VTAIL.n740 585
R64 VTAIL.n743 VTAIL.n742 585
R65 VTAIL.n694 VTAIL.n693 585
R66 VTAIL.n749 VTAIL.n748 585
R67 VTAIL.n751 VTAIL.n750 585
R68 VTAIL.n690 VTAIL.n689 585
R69 VTAIL.n757 VTAIL.n756 585
R70 VTAIL.n759 VTAIL.n758 585
R71 VTAIL.n686 VTAIL.n685 585
R72 VTAIL.n765 VTAIL.n764 585
R73 VTAIL.n767 VTAIL.n766 585
R74 VTAIL.n682 VTAIL.n681 585
R75 VTAIL.n773 VTAIL.n772 585
R76 VTAIL.n32 VTAIL.n31 585
R77 VTAIL.n37 VTAIL.n36 585
R78 VTAIL.n39 VTAIL.n38 585
R79 VTAIL.n28 VTAIL.n27 585
R80 VTAIL.n45 VTAIL.n44 585
R81 VTAIL.n47 VTAIL.n46 585
R82 VTAIL.n24 VTAIL.n23 585
R83 VTAIL.n54 VTAIL.n53 585
R84 VTAIL.n55 VTAIL.n22 585
R85 VTAIL.n57 VTAIL.n56 585
R86 VTAIL.n20 VTAIL.n19 585
R87 VTAIL.n63 VTAIL.n62 585
R88 VTAIL.n65 VTAIL.n64 585
R89 VTAIL.n16 VTAIL.n15 585
R90 VTAIL.n71 VTAIL.n70 585
R91 VTAIL.n73 VTAIL.n72 585
R92 VTAIL.n12 VTAIL.n11 585
R93 VTAIL.n79 VTAIL.n78 585
R94 VTAIL.n81 VTAIL.n80 585
R95 VTAIL.n8 VTAIL.n7 585
R96 VTAIL.n87 VTAIL.n86 585
R97 VTAIL.n89 VTAIL.n88 585
R98 VTAIL.n4 VTAIL.n3 585
R99 VTAIL.n95 VTAIL.n94 585
R100 VTAIL.n128 VTAIL.n127 585
R101 VTAIL.n133 VTAIL.n132 585
R102 VTAIL.n135 VTAIL.n134 585
R103 VTAIL.n124 VTAIL.n123 585
R104 VTAIL.n141 VTAIL.n140 585
R105 VTAIL.n143 VTAIL.n142 585
R106 VTAIL.n120 VTAIL.n119 585
R107 VTAIL.n150 VTAIL.n149 585
R108 VTAIL.n151 VTAIL.n118 585
R109 VTAIL.n153 VTAIL.n152 585
R110 VTAIL.n116 VTAIL.n115 585
R111 VTAIL.n159 VTAIL.n158 585
R112 VTAIL.n161 VTAIL.n160 585
R113 VTAIL.n112 VTAIL.n111 585
R114 VTAIL.n167 VTAIL.n166 585
R115 VTAIL.n169 VTAIL.n168 585
R116 VTAIL.n108 VTAIL.n107 585
R117 VTAIL.n175 VTAIL.n174 585
R118 VTAIL.n177 VTAIL.n176 585
R119 VTAIL.n104 VTAIL.n103 585
R120 VTAIL.n183 VTAIL.n182 585
R121 VTAIL.n185 VTAIL.n184 585
R122 VTAIL.n100 VTAIL.n99 585
R123 VTAIL.n191 VTAIL.n190 585
R124 VTAIL.n226 VTAIL.n225 585
R125 VTAIL.n231 VTAIL.n230 585
R126 VTAIL.n233 VTAIL.n232 585
R127 VTAIL.n222 VTAIL.n221 585
R128 VTAIL.n239 VTAIL.n238 585
R129 VTAIL.n241 VTAIL.n240 585
R130 VTAIL.n218 VTAIL.n217 585
R131 VTAIL.n248 VTAIL.n247 585
R132 VTAIL.n249 VTAIL.n216 585
R133 VTAIL.n251 VTAIL.n250 585
R134 VTAIL.n214 VTAIL.n213 585
R135 VTAIL.n257 VTAIL.n256 585
R136 VTAIL.n259 VTAIL.n258 585
R137 VTAIL.n210 VTAIL.n209 585
R138 VTAIL.n265 VTAIL.n264 585
R139 VTAIL.n267 VTAIL.n266 585
R140 VTAIL.n206 VTAIL.n205 585
R141 VTAIL.n273 VTAIL.n272 585
R142 VTAIL.n275 VTAIL.n274 585
R143 VTAIL.n202 VTAIL.n201 585
R144 VTAIL.n281 VTAIL.n280 585
R145 VTAIL.n283 VTAIL.n282 585
R146 VTAIL.n198 VTAIL.n197 585
R147 VTAIL.n289 VTAIL.n288 585
R148 VTAIL.n677 VTAIL.n676 585
R149 VTAIL.n586 VTAIL.n585 585
R150 VTAIL.n671 VTAIL.n670 585
R151 VTAIL.n669 VTAIL.n668 585
R152 VTAIL.n590 VTAIL.n589 585
R153 VTAIL.n663 VTAIL.n662 585
R154 VTAIL.n661 VTAIL.n660 585
R155 VTAIL.n594 VTAIL.n593 585
R156 VTAIL.n655 VTAIL.n654 585
R157 VTAIL.n653 VTAIL.n652 585
R158 VTAIL.n598 VTAIL.n597 585
R159 VTAIL.n647 VTAIL.n646 585
R160 VTAIL.n645 VTAIL.n644 585
R161 VTAIL.n602 VTAIL.n601 585
R162 VTAIL.n639 VTAIL.n638 585
R163 VTAIL.n637 VTAIL.n604 585
R164 VTAIL.n636 VTAIL.n635 585
R165 VTAIL.n607 VTAIL.n605 585
R166 VTAIL.n630 VTAIL.n629 585
R167 VTAIL.n628 VTAIL.n627 585
R168 VTAIL.n611 VTAIL.n610 585
R169 VTAIL.n622 VTAIL.n621 585
R170 VTAIL.n620 VTAIL.n619 585
R171 VTAIL.n615 VTAIL.n614 585
R172 VTAIL.n579 VTAIL.n578 585
R173 VTAIL.n488 VTAIL.n487 585
R174 VTAIL.n573 VTAIL.n572 585
R175 VTAIL.n571 VTAIL.n570 585
R176 VTAIL.n492 VTAIL.n491 585
R177 VTAIL.n565 VTAIL.n564 585
R178 VTAIL.n563 VTAIL.n562 585
R179 VTAIL.n496 VTAIL.n495 585
R180 VTAIL.n557 VTAIL.n556 585
R181 VTAIL.n555 VTAIL.n554 585
R182 VTAIL.n500 VTAIL.n499 585
R183 VTAIL.n549 VTAIL.n548 585
R184 VTAIL.n547 VTAIL.n546 585
R185 VTAIL.n504 VTAIL.n503 585
R186 VTAIL.n541 VTAIL.n540 585
R187 VTAIL.n539 VTAIL.n506 585
R188 VTAIL.n538 VTAIL.n537 585
R189 VTAIL.n509 VTAIL.n507 585
R190 VTAIL.n532 VTAIL.n531 585
R191 VTAIL.n530 VTAIL.n529 585
R192 VTAIL.n513 VTAIL.n512 585
R193 VTAIL.n524 VTAIL.n523 585
R194 VTAIL.n522 VTAIL.n521 585
R195 VTAIL.n517 VTAIL.n516 585
R196 VTAIL.n483 VTAIL.n482 585
R197 VTAIL.n392 VTAIL.n391 585
R198 VTAIL.n477 VTAIL.n476 585
R199 VTAIL.n475 VTAIL.n474 585
R200 VTAIL.n396 VTAIL.n395 585
R201 VTAIL.n469 VTAIL.n468 585
R202 VTAIL.n467 VTAIL.n466 585
R203 VTAIL.n400 VTAIL.n399 585
R204 VTAIL.n461 VTAIL.n460 585
R205 VTAIL.n459 VTAIL.n458 585
R206 VTAIL.n404 VTAIL.n403 585
R207 VTAIL.n453 VTAIL.n452 585
R208 VTAIL.n451 VTAIL.n450 585
R209 VTAIL.n408 VTAIL.n407 585
R210 VTAIL.n445 VTAIL.n444 585
R211 VTAIL.n443 VTAIL.n410 585
R212 VTAIL.n442 VTAIL.n441 585
R213 VTAIL.n413 VTAIL.n411 585
R214 VTAIL.n436 VTAIL.n435 585
R215 VTAIL.n434 VTAIL.n433 585
R216 VTAIL.n417 VTAIL.n416 585
R217 VTAIL.n428 VTAIL.n427 585
R218 VTAIL.n426 VTAIL.n425 585
R219 VTAIL.n421 VTAIL.n420 585
R220 VTAIL.n385 VTAIL.n384 585
R221 VTAIL.n294 VTAIL.n293 585
R222 VTAIL.n379 VTAIL.n378 585
R223 VTAIL.n377 VTAIL.n376 585
R224 VTAIL.n298 VTAIL.n297 585
R225 VTAIL.n371 VTAIL.n370 585
R226 VTAIL.n369 VTAIL.n368 585
R227 VTAIL.n302 VTAIL.n301 585
R228 VTAIL.n363 VTAIL.n362 585
R229 VTAIL.n361 VTAIL.n360 585
R230 VTAIL.n306 VTAIL.n305 585
R231 VTAIL.n355 VTAIL.n354 585
R232 VTAIL.n353 VTAIL.n352 585
R233 VTAIL.n310 VTAIL.n309 585
R234 VTAIL.n347 VTAIL.n346 585
R235 VTAIL.n345 VTAIL.n312 585
R236 VTAIL.n344 VTAIL.n343 585
R237 VTAIL.n315 VTAIL.n313 585
R238 VTAIL.n338 VTAIL.n337 585
R239 VTAIL.n336 VTAIL.n335 585
R240 VTAIL.n319 VTAIL.n318 585
R241 VTAIL.n330 VTAIL.n329 585
R242 VTAIL.n328 VTAIL.n327 585
R243 VTAIL.n323 VTAIL.n322 585
R244 VTAIL.n711 VTAIL.t14 329.036
R245 VTAIL.n33 VTAIL.t10 329.036
R246 VTAIL.n129 VTAIL.t1 329.036
R247 VTAIL.n227 VTAIL.t4 329.036
R248 VTAIL.n616 VTAIL.t6 329.036
R249 VTAIL.n518 VTAIL.t5 329.036
R250 VTAIL.n422 VTAIL.t9 329.036
R251 VTAIL.n324 VTAIL.t13 329.036
R252 VTAIL.n715 VTAIL.n709 171.744
R253 VTAIL.n716 VTAIL.n715 171.744
R254 VTAIL.n716 VTAIL.n705 171.744
R255 VTAIL.n723 VTAIL.n705 171.744
R256 VTAIL.n724 VTAIL.n723 171.744
R257 VTAIL.n724 VTAIL.n701 171.744
R258 VTAIL.n732 VTAIL.n701 171.744
R259 VTAIL.n733 VTAIL.n732 171.744
R260 VTAIL.n734 VTAIL.n733 171.744
R261 VTAIL.n734 VTAIL.n697 171.744
R262 VTAIL.n741 VTAIL.n697 171.744
R263 VTAIL.n742 VTAIL.n741 171.744
R264 VTAIL.n742 VTAIL.n693 171.744
R265 VTAIL.n749 VTAIL.n693 171.744
R266 VTAIL.n750 VTAIL.n749 171.744
R267 VTAIL.n750 VTAIL.n689 171.744
R268 VTAIL.n757 VTAIL.n689 171.744
R269 VTAIL.n758 VTAIL.n757 171.744
R270 VTAIL.n758 VTAIL.n685 171.744
R271 VTAIL.n765 VTAIL.n685 171.744
R272 VTAIL.n766 VTAIL.n765 171.744
R273 VTAIL.n766 VTAIL.n681 171.744
R274 VTAIL.n773 VTAIL.n681 171.744
R275 VTAIL.n37 VTAIL.n31 171.744
R276 VTAIL.n38 VTAIL.n37 171.744
R277 VTAIL.n38 VTAIL.n27 171.744
R278 VTAIL.n45 VTAIL.n27 171.744
R279 VTAIL.n46 VTAIL.n45 171.744
R280 VTAIL.n46 VTAIL.n23 171.744
R281 VTAIL.n54 VTAIL.n23 171.744
R282 VTAIL.n55 VTAIL.n54 171.744
R283 VTAIL.n56 VTAIL.n55 171.744
R284 VTAIL.n56 VTAIL.n19 171.744
R285 VTAIL.n63 VTAIL.n19 171.744
R286 VTAIL.n64 VTAIL.n63 171.744
R287 VTAIL.n64 VTAIL.n15 171.744
R288 VTAIL.n71 VTAIL.n15 171.744
R289 VTAIL.n72 VTAIL.n71 171.744
R290 VTAIL.n72 VTAIL.n11 171.744
R291 VTAIL.n79 VTAIL.n11 171.744
R292 VTAIL.n80 VTAIL.n79 171.744
R293 VTAIL.n80 VTAIL.n7 171.744
R294 VTAIL.n87 VTAIL.n7 171.744
R295 VTAIL.n88 VTAIL.n87 171.744
R296 VTAIL.n88 VTAIL.n3 171.744
R297 VTAIL.n95 VTAIL.n3 171.744
R298 VTAIL.n133 VTAIL.n127 171.744
R299 VTAIL.n134 VTAIL.n133 171.744
R300 VTAIL.n134 VTAIL.n123 171.744
R301 VTAIL.n141 VTAIL.n123 171.744
R302 VTAIL.n142 VTAIL.n141 171.744
R303 VTAIL.n142 VTAIL.n119 171.744
R304 VTAIL.n150 VTAIL.n119 171.744
R305 VTAIL.n151 VTAIL.n150 171.744
R306 VTAIL.n152 VTAIL.n151 171.744
R307 VTAIL.n152 VTAIL.n115 171.744
R308 VTAIL.n159 VTAIL.n115 171.744
R309 VTAIL.n160 VTAIL.n159 171.744
R310 VTAIL.n160 VTAIL.n111 171.744
R311 VTAIL.n167 VTAIL.n111 171.744
R312 VTAIL.n168 VTAIL.n167 171.744
R313 VTAIL.n168 VTAIL.n107 171.744
R314 VTAIL.n175 VTAIL.n107 171.744
R315 VTAIL.n176 VTAIL.n175 171.744
R316 VTAIL.n176 VTAIL.n103 171.744
R317 VTAIL.n183 VTAIL.n103 171.744
R318 VTAIL.n184 VTAIL.n183 171.744
R319 VTAIL.n184 VTAIL.n99 171.744
R320 VTAIL.n191 VTAIL.n99 171.744
R321 VTAIL.n231 VTAIL.n225 171.744
R322 VTAIL.n232 VTAIL.n231 171.744
R323 VTAIL.n232 VTAIL.n221 171.744
R324 VTAIL.n239 VTAIL.n221 171.744
R325 VTAIL.n240 VTAIL.n239 171.744
R326 VTAIL.n240 VTAIL.n217 171.744
R327 VTAIL.n248 VTAIL.n217 171.744
R328 VTAIL.n249 VTAIL.n248 171.744
R329 VTAIL.n250 VTAIL.n249 171.744
R330 VTAIL.n250 VTAIL.n213 171.744
R331 VTAIL.n257 VTAIL.n213 171.744
R332 VTAIL.n258 VTAIL.n257 171.744
R333 VTAIL.n258 VTAIL.n209 171.744
R334 VTAIL.n265 VTAIL.n209 171.744
R335 VTAIL.n266 VTAIL.n265 171.744
R336 VTAIL.n266 VTAIL.n205 171.744
R337 VTAIL.n273 VTAIL.n205 171.744
R338 VTAIL.n274 VTAIL.n273 171.744
R339 VTAIL.n274 VTAIL.n201 171.744
R340 VTAIL.n281 VTAIL.n201 171.744
R341 VTAIL.n282 VTAIL.n281 171.744
R342 VTAIL.n282 VTAIL.n197 171.744
R343 VTAIL.n289 VTAIL.n197 171.744
R344 VTAIL.n677 VTAIL.n585 171.744
R345 VTAIL.n670 VTAIL.n585 171.744
R346 VTAIL.n670 VTAIL.n669 171.744
R347 VTAIL.n669 VTAIL.n589 171.744
R348 VTAIL.n662 VTAIL.n589 171.744
R349 VTAIL.n662 VTAIL.n661 171.744
R350 VTAIL.n661 VTAIL.n593 171.744
R351 VTAIL.n654 VTAIL.n593 171.744
R352 VTAIL.n654 VTAIL.n653 171.744
R353 VTAIL.n653 VTAIL.n597 171.744
R354 VTAIL.n646 VTAIL.n597 171.744
R355 VTAIL.n646 VTAIL.n645 171.744
R356 VTAIL.n645 VTAIL.n601 171.744
R357 VTAIL.n638 VTAIL.n601 171.744
R358 VTAIL.n638 VTAIL.n637 171.744
R359 VTAIL.n637 VTAIL.n636 171.744
R360 VTAIL.n636 VTAIL.n605 171.744
R361 VTAIL.n629 VTAIL.n605 171.744
R362 VTAIL.n629 VTAIL.n628 171.744
R363 VTAIL.n628 VTAIL.n610 171.744
R364 VTAIL.n621 VTAIL.n610 171.744
R365 VTAIL.n621 VTAIL.n620 171.744
R366 VTAIL.n620 VTAIL.n614 171.744
R367 VTAIL.n579 VTAIL.n487 171.744
R368 VTAIL.n572 VTAIL.n487 171.744
R369 VTAIL.n572 VTAIL.n571 171.744
R370 VTAIL.n571 VTAIL.n491 171.744
R371 VTAIL.n564 VTAIL.n491 171.744
R372 VTAIL.n564 VTAIL.n563 171.744
R373 VTAIL.n563 VTAIL.n495 171.744
R374 VTAIL.n556 VTAIL.n495 171.744
R375 VTAIL.n556 VTAIL.n555 171.744
R376 VTAIL.n555 VTAIL.n499 171.744
R377 VTAIL.n548 VTAIL.n499 171.744
R378 VTAIL.n548 VTAIL.n547 171.744
R379 VTAIL.n547 VTAIL.n503 171.744
R380 VTAIL.n540 VTAIL.n503 171.744
R381 VTAIL.n540 VTAIL.n539 171.744
R382 VTAIL.n539 VTAIL.n538 171.744
R383 VTAIL.n538 VTAIL.n507 171.744
R384 VTAIL.n531 VTAIL.n507 171.744
R385 VTAIL.n531 VTAIL.n530 171.744
R386 VTAIL.n530 VTAIL.n512 171.744
R387 VTAIL.n523 VTAIL.n512 171.744
R388 VTAIL.n523 VTAIL.n522 171.744
R389 VTAIL.n522 VTAIL.n516 171.744
R390 VTAIL.n483 VTAIL.n391 171.744
R391 VTAIL.n476 VTAIL.n391 171.744
R392 VTAIL.n476 VTAIL.n475 171.744
R393 VTAIL.n475 VTAIL.n395 171.744
R394 VTAIL.n468 VTAIL.n395 171.744
R395 VTAIL.n468 VTAIL.n467 171.744
R396 VTAIL.n467 VTAIL.n399 171.744
R397 VTAIL.n460 VTAIL.n399 171.744
R398 VTAIL.n460 VTAIL.n459 171.744
R399 VTAIL.n459 VTAIL.n403 171.744
R400 VTAIL.n452 VTAIL.n403 171.744
R401 VTAIL.n452 VTAIL.n451 171.744
R402 VTAIL.n451 VTAIL.n407 171.744
R403 VTAIL.n444 VTAIL.n407 171.744
R404 VTAIL.n444 VTAIL.n443 171.744
R405 VTAIL.n443 VTAIL.n442 171.744
R406 VTAIL.n442 VTAIL.n411 171.744
R407 VTAIL.n435 VTAIL.n411 171.744
R408 VTAIL.n435 VTAIL.n434 171.744
R409 VTAIL.n434 VTAIL.n416 171.744
R410 VTAIL.n427 VTAIL.n416 171.744
R411 VTAIL.n427 VTAIL.n426 171.744
R412 VTAIL.n426 VTAIL.n420 171.744
R413 VTAIL.n385 VTAIL.n293 171.744
R414 VTAIL.n378 VTAIL.n293 171.744
R415 VTAIL.n378 VTAIL.n377 171.744
R416 VTAIL.n377 VTAIL.n297 171.744
R417 VTAIL.n370 VTAIL.n297 171.744
R418 VTAIL.n370 VTAIL.n369 171.744
R419 VTAIL.n369 VTAIL.n301 171.744
R420 VTAIL.n362 VTAIL.n301 171.744
R421 VTAIL.n362 VTAIL.n361 171.744
R422 VTAIL.n361 VTAIL.n305 171.744
R423 VTAIL.n354 VTAIL.n305 171.744
R424 VTAIL.n354 VTAIL.n353 171.744
R425 VTAIL.n353 VTAIL.n309 171.744
R426 VTAIL.n346 VTAIL.n309 171.744
R427 VTAIL.n346 VTAIL.n345 171.744
R428 VTAIL.n345 VTAIL.n344 171.744
R429 VTAIL.n344 VTAIL.n313 171.744
R430 VTAIL.n337 VTAIL.n313 171.744
R431 VTAIL.n337 VTAIL.n336 171.744
R432 VTAIL.n336 VTAIL.n318 171.744
R433 VTAIL.n329 VTAIL.n318 171.744
R434 VTAIL.n329 VTAIL.n328 171.744
R435 VTAIL.n328 VTAIL.n322 171.744
R436 VTAIL.t14 VTAIL.n709 85.8723
R437 VTAIL.t10 VTAIL.n31 85.8723
R438 VTAIL.t1 VTAIL.n127 85.8723
R439 VTAIL.t4 VTAIL.n225 85.8723
R440 VTAIL.t6 VTAIL.n614 85.8723
R441 VTAIL.t5 VTAIL.n516 85.8723
R442 VTAIL.t9 VTAIL.n420 85.8723
R443 VTAIL.t13 VTAIL.n322 85.8723
R444 VTAIL.n583 VTAIL.n582 56.0114
R445 VTAIL.n389 VTAIL.n388 56.0114
R446 VTAIL.n1 VTAIL.n0 56.0105
R447 VTAIL.n195 VTAIL.n194 56.0105
R448 VTAIL.n775 VTAIL.n774 34.3187
R449 VTAIL.n97 VTAIL.n96 34.3187
R450 VTAIL.n193 VTAIL.n192 34.3187
R451 VTAIL.n291 VTAIL.n290 34.3187
R452 VTAIL.n679 VTAIL.n678 34.3187
R453 VTAIL.n581 VTAIL.n580 34.3187
R454 VTAIL.n485 VTAIL.n484 34.3187
R455 VTAIL.n387 VTAIL.n386 34.3187
R456 VTAIL.n775 VTAIL.n679 28.5996
R457 VTAIL.n387 VTAIL.n291 28.5996
R458 VTAIL.n735 VTAIL.n700 13.1884
R459 VTAIL.n57 VTAIL.n22 13.1884
R460 VTAIL.n153 VTAIL.n118 13.1884
R461 VTAIL.n251 VTAIL.n216 13.1884
R462 VTAIL.n639 VTAIL.n604 13.1884
R463 VTAIL.n541 VTAIL.n506 13.1884
R464 VTAIL.n445 VTAIL.n410 13.1884
R465 VTAIL.n347 VTAIL.n312 13.1884
R466 VTAIL.n731 VTAIL.n730 12.8005
R467 VTAIL.n736 VTAIL.n698 12.8005
R468 VTAIL.n53 VTAIL.n52 12.8005
R469 VTAIL.n58 VTAIL.n20 12.8005
R470 VTAIL.n149 VTAIL.n148 12.8005
R471 VTAIL.n154 VTAIL.n116 12.8005
R472 VTAIL.n247 VTAIL.n246 12.8005
R473 VTAIL.n252 VTAIL.n214 12.8005
R474 VTAIL.n640 VTAIL.n602 12.8005
R475 VTAIL.n635 VTAIL.n606 12.8005
R476 VTAIL.n542 VTAIL.n504 12.8005
R477 VTAIL.n537 VTAIL.n508 12.8005
R478 VTAIL.n446 VTAIL.n408 12.8005
R479 VTAIL.n441 VTAIL.n412 12.8005
R480 VTAIL.n348 VTAIL.n310 12.8005
R481 VTAIL.n343 VTAIL.n314 12.8005
R482 VTAIL.n729 VTAIL.n702 12.0247
R483 VTAIL.n740 VTAIL.n739 12.0247
R484 VTAIL.n51 VTAIL.n24 12.0247
R485 VTAIL.n62 VTAIL.n61 12.0247
R486 VTAIL.n147 VTAIL.n120 12.0247
R487 VTAIL.n158 VTAIL.n157 12.0247
R488 VTAIL.n245 VTAIL.n218 12.0247
R489 VTAIL.n256 VTAIL.n255 12.0247
R490 VTAIL.n644 VTAIL.n643 12.0247
R491 VTAIL.n634 VTAIL.n607 12.0247
R492 VTAIL.n546 VTAIL.n545 12.0247
R493 VTAIL.n536 VTAIL.n509 12.0247
R494 VTAIL.n450 VTAIL.n449 12.0247
R495 VTAIL.n440 VTAIL.n413 12.0247
R496 VTAIL.n352 VTAIL.n351 12.0247
R497 VTAIL.n342 VTAIL.n315 12.0247
R498 VTAIL.n726 VTAIL.n725 11.249
R499 VTAIL.n743 VTAIL.n696 11.249
R500 VTAIL.n772 VTAIL.n680 11.249
R501 VTAIL.n48 VTAIL.n47 11.249
R502 VTAIL.n65 VTAIL.n18 11.249
R503 VTAIL.n94 VTAIL.n2 11.249
R504 VTAIL.n144 VTAIL.n143 11.249
R505 VTAIL.n161 VTAIL.n114 11.249
R506 VTAIL.n190 VTAIL.n98 11.249
R507 VTAIL.n242 VTAIL.n241 11.249
R508 VTAIL.n259 VTAIL.n212 11.249
R509 VTAIL.n288 VTAIL.n196 11.249
R510 VTAIL.n676 VTAIL.n584 11.249
R511 VTAIL.n647 VTAIL.n600 11.249
R512 VTAIL.n631 VTAIL.n630 11.249
R513 VTAIL.n578 VTAIL.n486 11.249
R514 VTAIL.n549 VTAIL.n502 11.249
R515 VTAIL.n533 VTAIL.n532 11.249
R516 VTAIL.n482 VTAIL.n390 11.249
R517 VTAIL.n453 VTAIL.n406 11.249
R518 VTAIL.n437 VTAIL.n436 11.249
R519 VTAIL.n384 VTAIL.n292 11.249
R520 VTAIL.n355 VTAIL.n308 11.249
R521 VTAIL.n339 VTAIL.n338 11.249
R522 VTAIL.n711 VTAIL.n710 10.7239
R523 VTAIL.n33 VTAIL.n32 10.7239
R524 VTAIL.n129 VTAIL.n128 10.7239
R525 VTAIL.n227 VTAIL.n226 10.7239
R526 VTAIL.n616 VTAIL.n615 10.7239
R527 VTAIL.n518 VTAIL.n517 10.7239
R528 VTAIL.n422 VTAIL.n421 10.7239
R529 VTAIL.n324 VTAIL.n323 10.7239
R530 VTAIL.n722 VTAIL.n704 10.4732
R531 VTAIL.n744 VTAIL.n694 10.4732
R532 VTAIL.n771 VTAIL.n682 10.4732
R533 VTAIL.n44 VTAIL.n26 10.4732
R534 VTAIL.n66 VTAIL.n16 10.4732
R535 VTAIL.n93 VTAIL.n4 10.4732
R536 VTAIL.n140 VTAIL.n122 10.4732
R537 VTAIL.n162 VTAIL.n112 10.4732
R538 VTAIL.n189 VTAIL.n100 10.4732
R539 VTAIL.n238 VTAIL.n220 10.4732
R540 VTAIL.n260 VTAIL.n210 10.4732
R541 VTAIL.n287 VTAIL.n198 10.4732
R542 VTAIL.n675 VTAIL.n586 10.4732
R543 VTAIL.n648 VTAIL.n598 10.4732
R544 VTAIL.n627 VTAIL.n609 10.4732
R545 VTAIL.n577 VTAIL.n488 10.4732
R546 VTAIL.n550 VTAIL.n500 10.4732
R547 VTAIL.n529 VTAIL.n511 10.4732
R548 VTAIL.n481 VTAIL.n392 10.4732
R549 VTAIL.n454 VTAIL.n404 10.4732
R550 VTAIL.n433 VTAIL.n415 10.4732
R551 VTAIL.n383 VTAIL.n294 10.4732
R552 VTAIL.n356 VTAIL.n306 10.4732
R553 VTAIL.n335 VTAIL.n317 10.4732
R554 VTAIL.n721 VTAIL.n706 9.69747
R555 VTAIL.n748 VTAIL.n747 9.69747
R556 VTAIL.n768 VTAIL.n767 9.69747
R557 VTAIL.n43 VTAIL.n28 9.69747
R558 VTAIL.n70 VTAIL.n69 9.69747
R559 VTAIL.n90 VTAIL.n89 9.69747
R560 VTAIL.n139 VTAIL.n124 9.69747
R561 VTAIL.n166 VTAIL.n165 9.69747
R562 VTAIL.n186 VTAIL.n185 9.69747
R563 VTAIL.n237 VTAIL.n222 9.69747
R564 VTAIL.n264 VTAIL.n263 9.69747
R565 VTAIL.n284 VTAIL.n283 9.69747
R566 VTAIL.n672 VTAIL.n671 9.69747
R567 VTAIL.n652 VTAIL.n651 9.69747
R568 VTAIL.n626 VTAIL.n611 9.69747
R569 VTAIL.n574 VTAIL.n573 9.69747
R570 VTAIL.n554 VTAIL.n553 9.69747
R571 VTAIL.n528 VTAIL.n513 9.69747
R572 VTAIL.n478 VTAIL.n477 9.69747
R573 VTAIL.n458 VTAIL.n457 9.69747
R574 VTAIL.n432 VTAIL.n417 9.69747
R575 VTAIL.n380 VTAIL.n379 9.69747
R576 VTAIL.n360 VTAIL.n359 9.69747
R577 VTAIL.n334 VTAIL.n319 9.69747
R578 VTAIL.n770 VTAIL.n680 9.45567
R579 VTAIL.n92 VTAIL.n2 9.45567
R580 VTAIL.n188 VTAIL.n98 9.45567
R581 VTAIL.n286 VTAIL.n196 9.45567
R582 VTAIL.n674 VTAIL.n584 9.45567
R583 VTAIL.n576 VTAIL.n486 9.45567
R584 VTAIL.n480 VTAIL.n390 9.45567
R585 VTAIL.n382 VTAIL.n292 9.45567
R586 VTAIL.n688 VTAIL.n687 9.3005
R587 VTAIL.n761 VTAIL.n760 9.3005
R588 VTAIL.n763 VTAIL.n762 9.3005
R589 VTAIL.n684 VTAIL.n683 9.3005
R590 VTAIL.n769 VTAIL.n768 9.3005
R591 VTAIL.n771 VTAIL.n770 9.3005
R592 VTAIL.n753 VTAIL.n752 9.3005
R593 VTAIL.n692 VTAIL.n691 9.3005
R594 VTAIL.n747 VTAIL.n746 9.3005
R595 VTAIL.n745 VTAIL.n744 9.3005
R596 VTAIL.n696 VTAIL.n695 9.3005
R597 VTAIL.n739 VTAIL.n738 9.3005
R598 VTAIL.n737 VTAIL.n736 9.3005
R599 VTAIL.n713 VTAIL.n712 9.3005
R600 VTAIL.n708 VTAIL.n707 9.3005
R601 VTAIL.n719 VTAIL.n718 9.3005
R602 VTAIL.n721 VTAIL.n720 9.3005
R603 VTAIL.n704 VTAIL.n703 9.3005
R604 VTAIL.n727 VTAIL.n726 9.3005
R605 VTAIL.n729 VTAIL.n728 9.3005
R606 VTAIL.n730 VTAIL.n699 9.3005
R607 VTAIL.n755 VTAIL.n754 9.3005
R608 VTAIL.n10 VTAIL.n9 9.3005
R609 VTAIL.n83 VTAIL.n82 9.3005
R610 VTAIL.n85 VTAIL.n84 9.3005
R611 VTAIL.n6 VTAIL.n5 9.3005
R612 VTAIL.n91 VTAIL.n90 9.3005
R613 VTAIL.n93 VTAIL.n92 9.3005
R614 VTAIL.n75 VTAIL.n74 9.3005
R615 VTAIL.n14 VTAIL.n13 9.3005
R616 VTAIL.n69 VTAIL.n68 9.3005
R617 VTAIL.n67 VTAIL.n66 9.3005
R618 VTAIL.n18 VTAIL.n17 9.3005
R619 VTAIL.n61 VTAIL.n60 9.3005
R620 VTAIL.n59 VTAIL.n58 9.3005
R621 VTAIL.n35 VTAIL.n34 9.3005
R622 VTAIL.n30 VTAIL.n29 9.3005
R623 VTAIL.n41 VTAIL.n40 9.3005
R624 VTAIL.n43 VTAIL.n42 9.3005
R625 VTAIL.n26 VTAIL.n25 9.3005
R626 VTAIL.n49 VTAIL.n48 9.3005
R627 VTAIL.n51 VTAIL.n50 9.3005
R628 VTAIL.n52 VTAIL.n21 9.3005
R629 VTAIL.n77 VTAIL.n76 9.3005
R630 VTAIL.n106 VTAIL.n105 9.3005
R631 VTAIL.n179 VTAIL.n178 9.3005
R632 VTAIL.n181 VTAIL.n180 9.3005
R633 VTAIL.n102 VTAIL.n101 9.3005
R634 VTAIL.n187 VTAIL.n186 9.3005
R635 VTAIL.n189 VTAIL.n188 9.3005
R636 VTAIL.n171 VTAIL.n170 9.3005
R637 VTAIL.n110 VTAIL.n109 9.3005
R638 VTAIL.n165 VTAIL.n164 9.3005
R639 VTAIL.n163 VTAIL.n162 9.3005
R640 VTAIL.n114 VTAIL.n113 9.3005
R641 VTAIL.n157 VTAIL.n156 9.3005
R642 VTAIL.n155 VTAIL.n154 9.3005
R643 VTAIL.n131 VTAIL.n130 9.3005
R644 VTAIL.n126 VTAIL.n125 9.3005
R645 VTAIL.n137 VTAIL.n136 9.3005
R646 VTAIL.n139 VTAIL.n138 9.3005
R647 VTAIL.n122 VTAIL.n121 9.3005
R648 VTAIL.n145 VTAIL.n144 9.3005
R649 VTAIL.n147 VTAIL.n146 9.3005
R650 VTAIL.n148 VTAIL.n117 9.3005
R651 VTAIL.n173 VTAIL.n172 9.3005
R652 VTAIL.n204 VTAIL.n203 9.3005
R653 VTAIL.n277 VTAIL.n276 9.3005
R654 VTAIL.n279 VTAIL.n278 9.3005
R655 VTAIL.n200 VTAIL.n199 9.3005
R656 VTAIL.n285 VTAIL.n284 9.3005
R657 VTAIL.n287 VTAIL.n286 9.3005
R658 VTAIL.n269 VTAIL.n268 9.3005
R659 VTAIL.n208 VTAIL.n207 9.3005
R660 VTAIL.n263 VTAIL.n262 9.3005
R661 VTAIL.n261 VTAIL.n260 9.3005
R662 VTAIL.n212 VTAIL.n211 9.3005
R663 VTAIL.n255 VTAIL.n254 9.3005
R664 VTAIL.n253 VTAIL.n252 9.3005
R665 VTAIL.n229 VTAIL.n228 9.3005
R666 VTAIL.n224 VTAIL.n223 9.3005
R667 VTAIL.n235 VTAIL.n234 9.3005
R668 VTAIL.n237 VTAIL.n236 9.3005
R669 VTAIL.n220 VTAIL.n219 9.3005
R670 VTAIL.n243 VTAIL.n242 9.3005
R671 VTAIL.n245 VTAIL.n244 9.3005
R672 VTAIL.n246 VTAIL.n215 9.3005
R673 VTAIL.n271 VTAIL.n270 9.3005
R674 VTAIL.n675 VTAIL.n674 9.3005
R675 VTAIL.n673 VTAIL.n672 9.3005
R676 VTAIL.n588 VTAIL.n587 9.3005
R677 VTAIL.n667 VTAIL.n666 9.3005
R678 VTAIL.n665 VTAIL.n664 9.3005
R679 VTAIL.n592 VTAIL.n591 9.3005
R680 VTAIL.n659 VTAIL.n658 9.3005
R681 VTAIL.n657 VTAIL.n656 9.3005
R682 VTAIL.n596 VTAIL.n595 9.3005
R683 VTAIL.n651 VTAIL.n650 9.3005
R684 VTAIL.n649 VTAIL.n648 9.3005
R685 VTAIL.n600 VTAIL.n599 9.3005
R686 VTAIL.n643 VTAIL.n642 9.3005
R687 VTAIL.n641 VTAIL.n640 9.3005
R688 VTAIL.n606 VTAIL.n603 9.3005
R689 VTAIL.n634 VTAIL.n633 9.3005
R690 VTAIL.n632 VTAIL.n631 9.3005
R691 VTAIL.n609 VTAIL.n608 9.3005
R692 VTAIL.n626 VTAIL.n625 9.3005
R693 VTAIL.n624 VTAIL.n623 9.3005
R694 VTAIL.n613 VTAIL.n612 9.3005
R695 VTAIL.n618 VTAIL.n617 9.3005
R696 VTAIL.n520 VTAIL.n519 9.3005
R697 VTAIL.n515 VTAIL.n514 9.3005
R698 VTAIL.n526 VTAIL.n525 9.3005
R699 VTAIL.n528 VTAIL.n527 9.3005
R700 VTAIL.n511 VTAIL.n510 9.3005
R701 VTAIL.n534 VTAIL.n533 9.3005
R702 VTAIL.n536 VTAIL.n535 9.3005
R703 VTAIL.n508 VTAIL.n505 9.3005
R704 VTAIL.n567 VTAIL.n566 9.3005
R705 VTAIL.n569 VTAIL.n568 9.3005
R706 VTAIL.n490 VTAIL.n489 9.3005
R707 VTAIL.n575 VTAIL.n574 9.3005
R708 VTAIL.n577 VTAIL.n576 9.3005
R709 VTAIL.n494 VTAIL.n493 9.3005
R710 VTAIL.n561 VTAIL.n560 9.3005
R711 VTAIL.n559 VTAIL.n558 9.3005
R712 VTAIL.n498 VTAIL.n497 9.3005
R713 VTAIL.n553 VTAIL.n552 9.3005
R714 VTAIL.n551 VTAIL.n550 9.3005
R715 VTAIL.n502 VTAIL.n501 9.3005
R716 VTAIL.n545 VTAIL.n544 9.3005
R717 VTAIL.n543 VTAIL.n542 9.3005
R718 VTAIL.n424 VTAIL.n423 9.3005
R719 VTAIL.n419 VTAIL.n418 9.3005
R720 VTAIL.n430 VTAIL.n429 9.3005
R721 VTAIL.n432 VTAIL.n431 9.3005
R722 VTAIL.n415 VTAIL.n414 9.3005
R723 VTAIL.n438 VTAIL.n437 9.3005
R724 VTAIL.n440 VTAIL.n439 9.3005
R725 VTAIL.n412 VTAIL.n409 9.3005
R726 VTAIL.n471 VTAIL.n470 9.3005
R727 VTAIL.n473 VTAIL.n472 9.3005
R728 VTAIL.n394 VTAIL.n393 9.3005
R729 VTAIL.n479 VTAIL.n478 9.3005
R730 VTAIL.n481 VTAIL.n480 9.3005
R731 VTAIL.n398 VTAIL.n397 9.3005
R732 VTAIL.n465 VTAIL.n464 9.3005
R733 VTAIL.n463 VTAIL.n462 9.3005
R734 VTAIL.n402 VTAIL.n401 9.3005
R735 VTAIL.n457 VTAIL.n456 9.3005
R736 VTAIL.n455 VTAIL.n454 9.3005
R737 VTAIL.n406 VTAIL.n405 9.3005
R738 VTAIL.n449 VTAIL.n448 9.3005
R739 VTAIL.n447 VTAIL.n446 9.3005
R740 VTAIL.n326 VTAIL.n325 9.3005
R741 VTAIL.n321 VTAIL.n320 9.3005
R742 VTAIL.n332 VTAIL.n331 9.3005
R743 VTAIL.n334 VTAIL.n333 9.3005
R744 VTAIL.n317 VTAIL.n316 9.3005
R745 VTAIL.n340 VTAIL.n339 9.3005
R746 VTAIL.n342 VTAIL.n341 9.3005
R747 VTAIL.n314 VTAIL.n311 9.3005
R748 VTAIL.n373 VTAIL.n372 9.3005
R749 VTAIL.n375 VTAIL.n374 9.3005
R750 VTAIL.n296 VTAIL.n295 9.3005
R751 VTAIL.n381 VTAIL.n380 9.3005
R752 VTAIL.n383 VTAIL.n382 9.3005
R753 VTAIL.n300 VTAIL.n299 9.3005
R754 VTAIL.n367 VTAIL.n366 9.3005
R755 VTAIL.n365 VTAIL.n364 9.3005
R756 VTAIL.n304 VTAIL.n303 9.3005
R757 VTAIL.n359 VTAIL.n358 9.3005
R758 VTAIL.n357 VTAIL.n356 9.3005
R759 VTAIL.n308 VTAIL.n307 9.3005
R760 VTAIL.n351 VTAIL.n350 9.3005
R761 VTAIL.n349 VTAIL.n348 9.3005
R762 VTAIL.n718 VTAIL.n717 8.92171
R763 VTAIL.n751 VTAIL.n692 8.92171
R764 VTAIL.n764 VTAIL.n684 8.92171
R765 VTAIL.n40 VTAIL.n39 8.92171
R766 VTAIL.n73 VTAIL.n14 8.92171
R767 VTAIL.n86 VTAIL.n6 8.92171
R768 VTAIL.n136 VTAIL.n135 8.92171
R769 VTAIL.n169 VTAIL.n110 8.92171
R770 VTAIL.n182 VTAIL.n102 8.92171
R771 VTAIL.n234 VTAIL.n233 8.92171
R772 VTAIL.n267 VTAIL.n208 8.92171
R773 VTAIL.n280 VTAIL.n200 8.92171
R774 VTAIL.n668 VTAIL.n588 8.92171
R775 VTAIL.n655 VTAIL.n596 8.92171
R776 VTAIL.n623 VTAIL.n622 8.92171
R777 VTAIL.n570 VTAIL.n490 8.92171
R778 VTAIL.n557 VTAIL.n498 8.92171
R779 VTAIL.n525 VTAIL.n524 8.92171
R780 VTAIL.n474 VTAIL.n394 8.92171
R781 VTAIL.n461 VTAIL.n402 8.92171
R782 VTAIL.n429 VTAIL.n428 8.92171
R783 VTAIL.n376 VTAIL.n296 8.92171
R784 VTAIL.n363 VTAIL.n304 8.92171
R785 VTAIL.n331 VTAIL.n330 8.92171
R786 VTAIL.n714 VTAIL.n708 8.14595
R787 VTAIL.n752 VTAIL.n690 8.14595
R788 VTAIL.n763 VTAIL.n686 8.14595
R789 VTAIL.n36 VTAIL.n30 8.14595
R790 VTAIL.n74 VTAIL.n12 8.14595
R791 VTAIL.n85 VTAIL.n8 8.14595
R792 VTAIL.n132 VTAIL.n126 8.14595
R793 VTAIL.n170 VTAIL.n108 8.14595
R794 VTAIL.n181 VTAIL.n104 8.14595
R795 VTAIL.n230 VTAIL.n224 8.14595
R796 VTAIL.n268 VTAIL.n206 8.14595
R797 VTAIL.n279 VTAIL.n202 8.14595
R798 VTAIL.n667 VTAIL.n590 8.14595
R799 VTAIL.n656 VTAIL.n594 8.14595
R800 VTAIL.n619 VTAIL.n613 8.14595
R801 VTAIL.n569 VTAIL.n492 8.14595
R802 VTAIL.n558 VTAIL.n496 8.14595
R803 VTAIL.n521 VTAIL.n515 8.14595
R804 VTAIL.n473 VTAIL.n396 8.14595
R805 VTAIL.n462 VTAIL.n400 8.14595
R806 VTAIL.n425 VTAIL.n419 8.14595
R807 VTAIL.n375 VTAIL.n298 8.14595
R808 VTAIL.n364 VTAIL.n302 8.14595
R809 VTAIL.n327 VTAIL.n321 8.14595
R810 VTAIL.n713 VTAIL.n710 7.3702
R811 VTAIL.n756 VTAIL.n755 7.3702
R812 VTAIL.n760 VTAIL.n759 7.3702
R813 VTAIL.n35 VTAIL.n32 7.3702
R814 VTAIL.n78 VTAIL.n77 7.3702
R815 VTAIL.n82 VTAIL.n81 7.3702
R816 VTAIL.n131 VTAIL.n128 7.3702
R817 VTAIL.n174 VTAIL.n173 7.3702
R818 VTAIL.n178 VTAIL.n177 7.3702
R819 VTAIL.n229 VTAIL.n226 7.3702
R820 VTAIL.n272 VTAIL.n271 7.3702
R821 VTAIL.n276 VTAIL.n275 7.3702
R822 VTAIL.n664 VTAIL.n663 7.3702
R823 VTAIL.n660 VTAIL.n659 7.3702
R824 VTAIL.n618 VTAIL.n615 7.3702
R825 VTAIL.n566 VTAIL.n565 7.3702
R826 VTAIL.n562 VTAIL.n561 7.3702
R827 VTAIL.n520 VTAIL.n517 7.3702
R828 VTAIL.n470 VTAIL.n469 7.3702
R829 VTAIL.n466 VTAIL.n465 7.3702
R830 VTAIL.n424 VTAIL.n421 7.3702
R831 VTAIL.n372 VTAIL.n371 7.3702
R832 VTAIL.n368 VTAIL.n367 7.3702
R833 VTAIL.n326 VTAIL.n323 7.3702
R834 VTAIL.n756 VTAIL.n688 6.59444
R835 VTAIL.n759 VTAIL.n688 6.59444
R836 VTAIL.n78 VTAIL.n10 6.59444
R837 VTAIL.n81 VTAIL.n10 6.59444
R838 VTAIL.n174 VTAIL.n106 6.59444
R839 VTAIL.n177 VTAIL.n106 6.59444
R840 VTAIL.n272 VTAIL.n204 6.59444
R841 VTAIL.n275 VTAIL.n204 6.59444
R842 VTAIL.n663 VTAIL.n592 6.59444
R843 VTAIL.n660 VTAIL.n592 6.59444
R844 VTAIL.n565 VTAIL.n494 6.59444
R845 VTAIL.n562 VTAIL.n494 6.59444
R846 VTAIL.n469 VTAIL.n398 6.59444
R847 VTAIL.n466 VTAIL.n398 6.59444
R848 VTAIL.n371 VTAIL.n300 6.59444
R849 VTAIL.n368 VTAIL.n300 6.59444
R850 VTAIL.n714 VTAIL.n713 5.81868
R851 VTAIL.n755 VTAIL.n690 5.81868
R852 VTAIL.n760 VTAIL.n686 5.81868
R853 VTAIL.n36 VTAIL.n35 5.81868
R854 VTAIL.n77 VTAIL.n12 5.81868
R855 VTAIL.n82 VTAIL.n8 5.81868
R856 VTAIL.n132 VTAIL.n131 5.81868
R857 VTAIL.n173 VTAIL.n108 5.81868
R858 VTAIL.n178 VTAIL.n104 5.81868
R859 VTAIL.n230 VTAIL.n229 5.81868
R860 VTAIL.n271 VTAIL.n206 5.81868
R861 VTAIL.n276 VTAIL.n202 5.81868
R862 VTAIL.n664 VTAIL.n590 5.81868
R863 VTAIL.n659 VTAIL.n594 5.81868
R864 VTAIL.n619 VTAIL.n618 5.81868
R865 VTAIL.n566 VTAIL.n492 5.81868
R866 VTAIL.n561 VTAIL.n496 5.81868
R867 VTAIL.n521 VTAIL.n520 5.81868
R868 VTAIL.n470 VTAIL.n396 5.81868
R869 VTAIL.n465 VTAIL.n400 5.81868
R870 VTAIL.n425 VTAIL.n424 5.81868
R871 VTAIL.n372 VTAIL.n298 5.81868
R872 VTAIL.n367 VTAIL.n302 5.81868
R873 VTAIL.n327 VTAIL.n326 5.81868
R874 VTAIL.n717 VTAIL.n708 5.04292
R875 VTAIL.n752 VTAIL.n751 5.04292
R876 VTAIL.n764 VTAIL.n763 5.04292
R877 VTAIL.n39 VTAIL.n30 5.04292
R878 VTAIL.n74 VTAIL.n73 5.04292
R879 VTAIL.n86 VTAIL.n85 5.04292
R880 VTAIL.n135 VTAIL.n126 5.04292
R881 VTAIL.n170 VTAIL.n169 5.04292
R882 VTAIL.n182 VTAIL.n181 5.04292
R883 VTAIL.n233 VTAIL.n224 5.04292
R884 VTAIL.n268 VTAIL.n267 5.04292
R885 VTAIL.n280 VTAIL.n279 5.04292
R886 VTAIL.n668 VTAIL.n667 5.04292
R887 VTAIL.n656 VTAIL.n655 5.04292
R888 VTAIL.n622 VTAIL.n613 5.04292
R889 VTAIL.n570 VTAIL.n569 5.04292
R890 VTAIL.n558 VTAIL.n557 5.04292
R891 VTAIL.n524 VTAIL.n515 5.04292
R892 VTAIL.n474 VTAIL.n473 5.04292
R893 VTAIL.n462 VTAIL.n461 5.04292
R894 VTAIL.n428 VTAIL.n419 5.04292
R895 VTAIL.n376 VTAIL.n375 5.04292
R896 VTAIL.n364 VTAIL.n363 5.04292
R897 VTAIL.n330 VTAIL.n321 5.04292
R898 VTAIL.n718 VTAIL.n706 4.26717
R899 VTAIL.n748 VTAIL.n692 4.26717
R900 VTAIL.n767 VTAIL.n684 4.26717
R901 VTAIL.n40 VTAIL.n28 4.26717
R902 VTAIL.n70 VTAIL.n14 4.26717
R903 VTAIL.n89 VTAIL.n6 4.26717
R904 VTAIL.n136 VTAIL.n124 4.26717
R905 VTAIL.n166 VTAIL.n110 4.26717
R906 VTAIL.n185 VTAIL.n102 4.26717
R907 VTAIL.n234 VTAIL.n222 4.26717
R908 VTAIL.n264 VTAIL.n208 4.26717
R909 VTAIL.n283 VTAIL.n200 4.26717
R910 VTAIL.n671 VTAIL.n588 4.26717
R911 VTAIL.n652 VTAIL.n596 4.26717
R912 VTAIL.n623 VTAIL.n611 4.26717
R913 VTAIL.n573 VTAIL.n490 4.26717
R914 VTAIL.n554 VTAIL.n498 4.26717
R915 VTAIL.n525 VTAIL.n513 4.26717
R916 VTAIL.n477 VTAIL.n394 4.26717
R917 VTAIL.n458 VTAIL.n402 4.26717
R918 VTAIL.n429 VTAIL.n417 4.26717
R919 VTAIL.n379 VTAIL.n296 4.26717
R920 VTAIL.n360 VTAIL.n304 4.26717
R921 VTAIL.n331 VTAIL.n319 4.26717
R922 VTAIL.n722 VTAIL.n721 3.49141
R923 VTAIL.n747 VTAIL.n694 3.49141
R924 VTAIL.n768 VTAIL.n682 3.49141
R925 VTAIL.n44 VTAIL.n43 3.49141
R926 VTAIL.n69 VTAIL.n16 3.49141
R927 VTAIL.n90 VTAIL.n4 3.49141
R928 VTAIL.n140 VTAIL.n139 3.49141
R929 VTAIL.n165 VTAIL.n112 3.49141
R930 VTAIL.n186 VTAIL.n100 3.49141
R931 VTAIL.n238 VTAIL.n237 3.49141
R932 VTAIL.n263 VTAIL.n210 3.49141
R933 VTAIL.n284 VTAIL.n198 3.49141
R934 VTAIL.n672 VTAIL.n586 3.49141
R935 VTAIL.n651 VTAIL.n598 3.49141
R936 VTAIL.n627 VTAIL.n626 3.49141
R937 VTAIL.n574 VTAIL.n488 3.49141
R938 VTAIL.n553 VTAIL.n500 3.49141
R939 VTAIL.n529 VTAIL.n528 3.49141
R940 VTAIL.n478 VTAIL.n392 3.49141
R941 VTAIL.n457 VTAIL.n404 3.49141
R942 VTAIL.n433 VTAIL.n432 3.49141
R943 VTAIL.n380 VTAIL.n294 3.49141
R944 VTAIL.n359 VTAIL.n306 3.49141
R945 VTAIL.n335 VTAIL.n334 3.49141
R946 VTAIL.n725 VTAIL.n704 2.71565
R947 VTAIL.n744 VTAIL.n743 2.71565
R948 VTAIL.n772 VTAIL.n771 2.71565
R949 VTAIL.n47 VTAIL.n26 2.71565
R950 VTAIL.n66 VTAIL.n65 2.71565
R951 VTAIL.n94 VTAIL.n93 2.71565
R952 VTAIL.n143 VTAIL.n122 2.71565
R953 VTAIL.n162 VTAIL.n161 2.71565
R954 VTAIL.n190 VTAIL.n189 2.71565
R955 VTAIL.n241 VTAIL.n220 2.71565
R956 VTAIL.n260 VTAIL.n259 2.71565
R957 VTAIL.n288 VTAIL.n287 2.71565
R958 VTAIL.n676 VTAIL.n675 2.71565
R959 VTAIL.n648 VTAIL.n647 2.71565
R960 VTAIL.n630 VTAIL.n609 2.71565
R961 VTAIL.n578 VTAIL.n577 2.71565
R962 VTAIL.n550 VTAIL.n549 2.71565
R963 VTAIL.n532 VTAIL.n511 2.71565
R964 VTAIL.n482 VTAIL.n481 2.71565
R965 VTAIL.n454 VTAIL.n453 2.71565
R966 VTAIL.n436 VTAIL.n415 2.71565
R967 VTAIL.n384 VTAIL.n383 2.71565
R968 VTAIL.n356 VTAIL.n355 2.71565
R969 VTAIL.n338 VTAIL.n317 2.71565
R970 VTAIL.n617 VTAIL.n616 2.41282
R971 VTAIL.n519 VTAIL.n518 2.41282
R972 VTAIL.n423 VTAIL.n422 2.41282
R973 VTAIL.n325 VTAIL.n324 2.41282
R974 VTAIL.n712 VTAIL.n711 2.41282
R975 VTAIL.n34 VTAIL.n33 2.41282
R976 VTAIL.n130 VTAIL.n129 2.41282
R977 VTAIL.n228 VTAIL.n227 2.41282
R978 VTAIL.n726 VTAIL.n702 1.93989
R979 VTAIL.n740 VTAIL.n696 1.93989
R980 VTAIL.n774 VTAIL.n680 1.93989
R981 VTAIL.n48 VTAIL.n24 1.93989
R982 VTAIL.n62 VTAIL.n18 1.93989
R983 VTAIL.n96 VTAIL.n2 1.93989
R984 VTAIL.n144 VTAIL.n120 1.93989
R985 VTAIL.n158 VTAIL.n114 1.93989
R986 VTAIL.n192 VTAIL.n98 1.93989
R987 VTAIL.n242 VTAIL.n218 1.93989
R988 VTAIL.n256 VTAIL.n212 1.93989
R989 VTAIL.n290 VTAIL.n196 1.93989
R990 VTAIL.n678 VTAIL.n584 1.93989
R991 VTAIL.n644 VTAIL.n600 1.93989
R992 VTAIL.n631 VTAIL.n607 1.93989
R993 VTAIL.n580 VTAIL.n486 1.93989
R994 VTAIL.n546 VTAIL.n502 1.93989
R995 VTAIL.n533 VTAIL.n509 1.93989
R996 VTAIL.n484 VTAIL.n390 1.93989
R997 VTAIL.n450 VTAIL.n406 1.93989
R998 VTAIL.n437 VTAIL.n413 1.93989
R999 VTAIL.n386 VTAIL.n292 1.93989
R1000 VTAIL.n352 VTAIL.n308 1.93989
R1001 VTAIL.n339 VTAIL.n315 1.93989
R1002 VTAIL.n0 VTAIL.t11 1.87183
R1003 VTAIL.n0 VTAIL.t8 1.87183
R1004 VTAIL.n194 VTAIL.t0 1.87183
R1005 VTAIL.n194 VTAIL.t7 1.87183
R1006 VTAIL.n582 VTAIL.t3 1.87183
R1007 VTAIL.n582 VTAIL.t2 1.87183
R1008 VTAIL.n388 VTAIL.t15 1.87183
R1009 VTAIL.n388 VTAIL.t12 1.87183
R1010 VTAIL.n389 VTAIL.n387 1.25912
R1011 VTAIL.n485 VTAIL.n389 1.25912
R1012 VTAIL.n583 VTAIL.n581 1.25912
R1013 VTAIL.n679 VTAIL.n583 1.25912
R1014 VTAIL.n291 VTAIL.n195 1.25912
R1015 VTAIL.n195 VTAIL.n193 1.25912
R1016 VTAIL.n97 VTAIL.n1 1.25912
R1017 VTAIL VTAIL.n775 1.20093
R1018 VTAIL.n731 VTAIL.n729 1.16414
R1019 VTAIL.n739 VTAIL.n698 1.16414
R1020 VTAIL.n53 VTAIL.n51 1.16414
R1021 VTAIL.n61 VTAIL.n20 1.16414
R1022 VTAIL.n149 VTAIL.n147 1.16414
R1023 VTAIL.n157 VTAIL.n116 1.16414
R1024 VTAIL.n247 VTAIL.n245 1.16414
R1025 VTAIL.n255 VTAIL.n214 1.16414
R1026 VTAIL.n643 VTAIL.n602 1.16414
R1027 VTAIL.n635 VTAIL.n634 1.16414
R1028 VTAIL.n545 VTAIL.n504 1.16414
R1029 VTAIL.n537 VTAIL.n536 1.16414
R1030 VTAIL.n449 VTAIL.n408 1.16414
R1031 VTAIL.n441 VTAIL.n440 1.16414
R1032 VTAIL.n351 VTAIL.n310 1.16414
R1033 VTAIL.n343 VTAIL.n342 1.16414
R1034 VTAIL.n581 VTAIL.n485 0.470328
R1035 VTAIL.n193 VTAIL.n97 0.470328
R1036 VTAIL.n730 VTAIL.n700 0.388379
R1037 VTAIL.n736 VTAIL.n735 0.388379
R1038 VTAIL.n52 VTAIL.n22 0.388379
R1039 VTAIL.n58 VTAIL.n57 0.388379
R1040 VTAIL.n148 VTAIL.n118 0.388379
R1041 VTAIL.n154 VTAIL.n153 0.388379
R1042 VTAIL.n246 VTAIL.n216 0.388379
R1043 VTAIL.n252 VTAIL.n251 0.388379
R1044 VTAIL.n640 VTAIL.n639 0.388379
R1045 VTAIL.n606 VTAIL.n604 0.388379
R1046 VTAIL.n542 VTAIL.n541 0.388379
R1047 VTAIL.n508 VTAIL.n506 0.388379
R1048 VTAIL.n446 VTAIL.n445 0.388379
R1049 VTAIL.n412 VTAIL.n410 0.388379
R1050 VTAIL.n348 VTAIL.n347 0.388379
R1051 VTAIL.n314 VTAIL.n312 0.388379
R1052 VTAIL.n712 VTAIL.n707 0.155672
R1053 VTAIL.n719 VTAIL.n707 0.155672
R1054 VTAIL.n720 VTAIL.n719 0.155672
R1055 VTAIL.n720 VTAIL.n703 0.155672
R1056 VTAIL.n727 VTAIL.n703 0.155672
R1057 VTAIL.n728 VTAIL.n727 0.155672
R1058 VTAIL.n728 VTAIL.n699 0.155672
R1059 VTAIL.n737 VTAIL.n699 0.155672
R1060 VTAIL.n738 VTAIL.n737 0.155672
R1061 VTAIL.n738 VTAIL.n695 0.155672
R1062 VTAIL.n745 VTAIL.n695 0.155672
R1063 VTAIL.n746 VTAIL.n745 0.155672
R1064 VTAIL.n746 VTAIL.n691 0.155672
R1065 VTAIL.n753 VTAIL.n691 0.155672
R1066 VTAIL.n754 VTAIL.n753 0.155672
R1067 VTAIL.n754 VTAIL.n687 0.155672
R1068 VTAIL.n761 VTAIL.n687 0.155672
R1069 VTAIL.n762 VTAIL.n761 0.155672
R1070 VTAIL.n762 VTAIL.n683 0.155672
R1071 VTAIL.n769 VTAIL.n683 0.155672
R1072 VTAIL.n770 VTAIL.n769 0.155672
R1073 VTAIL.n34 VTAIL.n29 0.155672
R1074 VTAIL.n41 VTAIL.n29 0.155672
R1075 VTAIL.n42 VTAIL.n41 0.155672
R1076 VTAIL.n42 VTAIL.n25 0.155672
R1077 VTAIL.n49 VTAIL.n25 0.155672
R1078 VTAIL.n50 VTAIL.n49 0.155672
R1079 VTAIL.n50 VTAIL.n21 0.155672
R1080 VTAIL.n59 VTAIL.n21 0.155672
R1081 VTAIL.n60 VTAIL.n59 0.155672
R1082 VTAIL.n60 VTAIL.n17 0.155672
R1083 VTAIL.n67 VTAIL.n17 0.155672
R1084 VTAIL.n68 VTAIL.n67 0.155672
R1085 VTAIL.n68 VTAIL.n13 0.155672
R1086 VTAIL.n75 VTAIL.n13 0.155672
R1087 VTAIL.n76 VTAIL.n75 0.155672
R1088 VTAIL.n76 VTAIL.n9 0.155672
R1089 VTAIL.n83 VTAIL.n9 0.155672
R1090 VTAIL.n84 VTAIL.n83 0.155672
R1091 VTAIL.n84 VTAIL.n5 0.155672
R1092 VTAIL.n91 VTAIL.n5 0.155672
R1093 VTAIL.n92 VTAIL.n91 0.155672
R1094 VTAIL.n130 VTAIL.n125 0.155672
R1095 VTAIL.n137 VTAIL.n125 0.155672
R1096 VTAIL.n138 VTAIL.n137 0.155672
R1097 VTAIL.n138 VTAIL.n121 0.155672
R1098 VTAIL.n145 VTAIL.n121 0.155672
R1099 VTAIL.n146 VTAIL.n145 0.155672
R1100 VTAIL.n146 VTAIL.n117 0.155672
R1101 VTAIL.n155 VTAIL.n117 0.155672
R1102 VTAIL.n156 VTAIL.n155 0.155672
R1103 VTAIL.n156 VTAIL.n113 0.155672
R1104 VTAIL.n163 VTAIL.n113 0.155672
R1105 VTAIL.n164 VTAIL.n163 0.155672
R1106 VTAIL.n164 VTAIL.n109 0.155672
R1107 VTAIL.n171 VTAIL.n109 0.155672
R1108 VTAIL.n172 VTAIL.n171 0.155672
R1109 VTAIL.n172 VTAIL.n105 0.155672
R1110 VTAIL.n179 VTAIL.n105 0.155672
R1111 VTAIL.n180 VTAIL.n179 0.155672
R1112 VTAIL.n180 VTAIL.n101 0.155672
R1113 VTAIL.n187 VTAIL.n101 0.155672
R1114 VTAIL.n188 VTAIL.n187 0.155672
R1115 VTAIL.n228 VTAIL.n223 0.155672
R1116 VTAIL.n235 VTAIL.n223 0.155672
R1117 VTAIL.n236 VTAIL.n235 0.155672
R1118 VTAIL.n236 VTAIL.n219 0.155672
R1119 VTAIL.n243 VTAIL.n219 0.155672
R1120 VTAIL.n244 VTAIL.n243 0.155672
R1121 VTAIL.n244 VTAIL.n215 0.155672
R1122 VTAIL.n253 VTAIL.n215 0.155672
R1123 VTAIL.n254 VTAIL.n253 0.155672
R1124 VTAIL.n254 VTAIL.n211 0.155672
R1125 VTAIL.n261 VTAIL.n211 0.155672
R1126 VTAIL.n262 VTAIL.n261 0.155672
R1127 VTAIL.n262 VTAIL.n207 0.155672
R1128 VTAIL.n269 VTAIL.n207 0.155672
R1129 VTAIL.n270 VTAIL.n269 0.155672
R1130 VTAIL.n270 VTAIL.n203 0.155672
R1131 VTAIL.n277 VTAIL.n203 0.155672
R1132 VTAIL.n278 VTAIL.n277 0.155672
R1133 VTAIL.n278 VTAIL.n199 0.155672
R1134 VTAIL.n285 VTAIL.n199 0.155672
R1135 VTAIL.n286 VTAIL.n285 0.155672
R1136 VTAIL.n674 VTAIL.n673 0.155672
R1137 VTAIL.n673 VTAIL.n587 0.155672
R1138 VTAIL.n666 VTAIL.n587 0.155672
R1139 VTAIL.n666 VTAIL.n665 0.155672
R1140 VTAIL.n665 VTAIL.n591 0.155672
R1141 VTAIL.n658 VTAIL.n591 0.155672
R1142 VTAIL.n658 VTAIL.n657 0.155672
R1143 VTAIL.n657 VTAIL.n595 0.155672
R1144 VTAIL.n650 VTAIL.n595 0.155672
R1145 VTAIL.n650 VTAIL.n649 0.155672
R1146 VTAIL.n649 VTAIL.n599 0.155672
R1147 VTAIL.n642 VTAIL.n599 0.155672
R1148 VTAIL.n642 VTAIL.n641 0.155672
R1149 VTAIL.n641 VTAIL.n603 0.155672
R1150 VTAIL.n633 VTAIL.n603 0.155672
R1151 VTAIL.n633 VTAIL.n632 0.155672
R1152 VTAIL.n632 VTAIL.n608 0.155672
R1153 VTAIL.n625 VTAIL.n608 0.155672
R1154 VTAIL.n625 VTAIL.n624 0.155672
R1155 VTAIL.n624 VTAIL.n612 0.155672
R1156 VTAIL.n617 VTAIL.n612 0.155672
R1157 VTAIL.n576 VTAIL.n575 0.155672
R1158 VTAIL.n575 VTAIL.n489 0.155672
R1159 VTAIL.n568 VTAIL.n489 0.155672
R1160 VTAIL.n568 VTAIL.n567 0.155672
R1161 VTAIL.n567 VTAIL.n493 0.155672
R1162 VTAIL.n560 VTAIL.n493 0.155672
R1163 VTAIL.n560 VTAIL.n559 0.155672
R1164 VTAIL.n559 VTAIL.n497 0.155672
R1165 VTAIL.n552 VTAIL.n497 0.155672
R1166 VTAIL.n552 VTAIL.n551 0.155672
R1167 VTAIL.n551 VTAIL.n501 0.155672
R1168 VTAIL.n544 VTAIL.n501 0.155672
R1169 VTAIL.n544 VTAIL.n543 0.155672
R1170 VTAIL.n543 VTAIL.n505 0.155672
R1171 VTAIL.n535 VTAIL.n505 0.155672
R1172 VTAIL.n535 VTAIL.n534 0.155672
R1173 VTAIL.n534 VTAIL.n510 0.155672
R1174 VTAIL.n527 VTAIL.n510 0.155672
R1175 VTAIL.n527 VTAIL.n526 0.155672
R1176 VTAIL.n526 VTAIL.n514 0.155672
R1177 VTAIL.n519 VTAIL.n514 0.155672
R1178 VTAIL.n480 VTAIL.n479 0.155672
R1179 VTAIL.n479 VTAIL.n393 0.155672
R1180 VTAIL.n472 VTAIL.n393 0.155672
R1181 VTAIL.n472 VTAIL.n471 0.155672
R1182 VTAIL.n471 VTAIL.n397 0.155672
R1183 VTAIL.n464 VTAIL.n397 0.155672
R1184 VTAIL.n464 VTAIL.n463 0.155672
R1185 VTAIL.n463 VTAIL.n401 0.155672
R1186 VTAIL.n456 VTAIL.n401 0.155672
R1187 VTAIL.n456 VTAIL.n455 0.155672
R1188 VTAIL.n455 VTAIL.n405 0.155672
R1189 VTAIL.n448 VTAIL.n405 0.155672
R1190 VTAIL.n448 VTAIL.n447 0.155672
R1191 VTAIL.n447 VTAIL.n409 0.155672
R1192 VTAIL.n439 VTAIL.n409 0.155672
R1193 VTAIL.n439 VTAIL.n438 0.155672
R1194 VTAIL.n438 VTAIL.n414 0.155672
R1195 VTAIL.n431 VTAIL.n414 0.155672
R1196 VTAIL.n431 VTAIL.n430 0.155672
R1197 VTAIL.n430 VTAIL.n418 0.155672
R1198 VTAIL.n423 VTAIL.n418 0.155672
R1199 VTAIL.n382 VTAIL.n381 0.155672
R1200 VTAIL.n381 VTAIL.n295 0.155672
R1201 VTAIL.n374 VTAIL.n295 0.155672
R1202 VTAIL.n374 VTAIL.n373 0.155672
R1203 VTAIL.n373 VTAIL.n299 0.155672
R1204 VTAIL.n366 VTAIL.n299 0.155672
R1205 VTAIL.n366 VTAIL.n365 0.155672
R1206 VTAIL.n365 VTAIL.n303 0.155672
R1207 VTAIL.n358 VTAIL.n303 0.155672
R1208 VTAIL.n358 VTAIL.n357 0.155672
R1209 VTAIL.n357 VTAIL.n307 0.155672
R1210 VTAIL.n350 VTAIL.n307 0.155672
R1211 VTAIL.n350 VTAIL.n349 0.155672
R1212 VTAIL.n349 VTAIL.n311 0.155672
R1213 VTAIL.n341 VTAIL.n311 0.155672
R1214 VTAIL.n341 VTAIL.n340 0.155672
R1215 VTAIL.n340 VTAIL.n316 0.155672
R1216 VTAIL.n333 VTAIL.n316 0.155672
R1217 VTAIL.n333 VTAIL.n332 0.155672
R1218 VTAIL.n332 VTAIL.n320 0.155672
R1219 VTAIL.n325 VTAIL.n320 0.155672
R1220 VTAIL VTAIL.n1 0.0586897
R1221 VDD2.n2 VDD2.n1 73.2632
R1222 VDD2.n2 VDD2.n0 73.2632
R1223 VDD2 VDD2.n5 73.2602
R1224 VDD2.n4 VDD2.n3 72.6902
R1225 VDD2.n4 VDD2.n2 44.3532
R1226 VDD2.n5 VDD2.t6 1.87183
R1227 VDD2.n5 VDD2.t4 1.87183
R1228 VDD2.n3 VDD2.t2 1.87183
R1229 VDD2.n3 VDD2.t0 1.87183
R1230 VDD2.n1 VDD2.t5 1.87183
R1231 VDD2.n1 VDD2.t3 1.87183
R1232 VDD2.n0 VDD2.t1 1.87183
R1233 VDD2.n0 VDD2.t7 1.87183
R1234 VDD2 VDD2.n4 0.688
R1235 B.n422 B.n113 585
R1236 B.n421 B.n420 585
R1237 B.n419 B.n114 585
R1238 B.n418 B.n417 585
R1239 B.n416 B.n115 585
R1240 B.n415 B.n414 585
R1241 B.n413 B.n116 585
R1242 B.n412 B.n411 585
R1243 B.n410 B.n117 585
R1244 B.n409 B.n408 585
R1245 B.n407 B.n118 585
R1246 B.n406 B.n405 585
R1247 B.n404 B.n119 585
R1248 B.n403 B.n402 585
R1249 B.n401 B.n120 585
R1250 B.n400 B.n399 585
R1251 B.n398 B.n121 585
R1252 B.n397 B.n396 585
R1253 B.n395 B.n122 585
R1254 B.n394 B.n393 585
R1255 B.n392 B.n123 585
R1256 B.n391 B.n390 585
R1257 B.n389 B.n124 585
R1258 B.n388 B.n387 585
R1259 B.n386 B.n125 585
R1260 B.n385 B.n384 585
R1261 B.n383 B.n126 585
R1262 B.n382 B.n381 585
R1263 B.n380 B.n127 585
R1264 B.n379 B.n378 585
R1265 B.n377 B.n128 585
R1266 B.n376 B.n375 585
R1267 B.n374 B.n129 585
R1268 B.n373 B.n372 585
R1269 B.n371 B.n130 585
R1270 B.n370 B.n369 585
R1271 B.n368 B.n131 585
R1272 B.n367 B.n366 585
R1273 B.n365 B.n132 585
R1274 B.n364 B.n363 585
R1275 B.n362 B.n133 585
R1276 B.n361 B.n360 585
R1277 B.n359 B.n134 585
R1278 B.n358 B.n357 585
R1279 B.n356 B.n135 585
R1280 B.n355 B.n354 585
R1281 B.n353 B.n136 585
R1282 B.n352 B.n351 585
R1283 B.n350 B.n137 585
R1284 B.n349 B.n348 585
R1285 B.n347 B.n138 585
R1286 B.n346 B.n345 585
R1287 B.n344 B.n139 585
R1288 B.n343 B.n342 585
R1289 B.n341 B.n140 585
R1290 B.n340 B.n339 585
R1291 B.n338 B.n141 585
R1292 B.n336 B.n335 585
R1293 B.n334 B.n144 585
R1294 B.n333 B.n332 585
R1295 B.n331 B.n145 585
R1296 B.n330 B.n329 585
R1297 B.n328 B.n146 585
R1298 B.n327 B.n326 585
R1299 B.n325 B.n147 585
R1300 B.n324 B.n323 585
R1301 B.n322 B.n148 585
R1302 B.n321 B.n320 585
R1303 B.n316 B.n149 585
R1304 B.n315 B.n314 585
R1305 B.n313 B.n150 585
R1306 B.n312 B.n311 585
R1307 B.n310 B.n151 585
R1308 B.n309 B.n308 585
R1309 B.n307 B.n152 585
R1310 B.n306 B.n305 585
R1311 B.n304 B.n153 585
R1312 B.n303 B.n302 585
R1313 B.n301 B.n154 585
R1314 B.n300 B.n299 585
R1315 B.n298 B.n155 585
R1316 B.n297 B.n296 585
R1317 B.n295 B.n156 585
R1318 B.n294 B.n293 585
R1319 B.n292 B.n157 585
R1320 B.n291 B.n290 585
R1321 B.n289 B.n158 585
R1322 B.n288 B.n287 585
R1323 B.n286 B.n159 585
R1324 B.n285 B.n284 585
R1325 B.n283 B.n160 585
R1326 B.n282 B.n281 585
R1327 B.n280 B.n161 585
R1328 B.n279 B.n278 585
R1329 B.n277 B.n162 585
R1330 B.n276 B.n275 585
R1331 B.n274 B.n163 585
R1332 B.n273 B.n272 585
R1333 B.n271 B.n164 585
R1334 B.n270 B.n269 585
R1335 B.n268 B.n165 585
R1336 B.n267 B.n266 585
R1337 B.n265 B.n166 585
R1338 B.n264 B.n263 585
R1339 B.n262 B.n167 585
R1340 B.n261 B.n260 585
R1341 B.n259 B.n168 585
R1342 B.n258 B.n257 585
R1343 B.n256 B.n169 585
R1344 B.n255 B.n254 585
R1345 B.n253 B.n170 585
R1346 B.n252 B.n251 585
R1347 B.n250 B.n171 585
R1348 B.n249 B.n248 585
R1349 B.n247 B.n172 585
R1350 B.n246 B.n245 585
R1351 B.n244 B.n173 585
R1352 B.n243 B.n242 585
R1353 B.n241 B.n174 585
R1354 B.n240 B.n239 585
R1355 B.n238 B.n175 585
R1356 B.n237 B.n236 585
R1357 B.n235 B.n176 585
R1358 B.n234 B.n233 585
R1359 B.n424 B.n423 585
R1360 B.n425 B.n112 585
R1361 B.n427 B.n426 585
R1362 B.n428 B.n111 585
R1363 B.n430 B.n429 585
R1364 B.n431 B.n110 585
R1365 B.n433 B.n432 585
R1366 B.n434 B.n109 585
R1367 B.n436 B.n435 585
R1368 B.n437 B.n108 585
R1369 B.n439 B.n438 585
R1370 B.n440 B.n107 585
R1371 B.n442 B.n441 585
R1372 B.n443 B.n106 585
R1373 B.n445 B.n444 585
R1374 B.n446 B.n105 585
R1375 B.n448 B.n447 585
R1376 B.n449 B.n104 585
R1377 B.n451 B.n450 585
R1378 B.n452 B.n103 585
R1379 B.n454 B.n453 585
R1380 B.n455 B.n102 585
R1381 B.n457 B.n456 585
R1382 B.n458 B.n101 585
R1383 B.n460 B.n459 585
R1384 B.n461 B.n100 585
R1385 B.n463 B.n462 585
R1386 B.n464 B.n99 585
R1387 B.n466 B.n465 585
R1388 B.n467 B.n98 585
R1389 B.n469 B.n468 585
R1390 B.n470 B.n97 585
R1391 B.n472 B.n471 585
R1392 B.n473 B.n96 585
R1393 B.n475 B.n474 585
R1394 B.n476 B.n95 585
R1395 B.n478 B.n477 585
R1396 B.n479 B.n94 585
R1397 B.n481 B.n480 585
R1398 B.n482 B.n93 585
R1399 B.n484 B.n483 585
R1400 B.n485 B.n92 585
R1401 B.n487 B.n486 585
R1402 B.n488 B.n91 585
R1403 B.n490 B.n489 585
R1404 B.n491 B.n90 585
R1405 B.n493 B.n492 585
R1406 B.n494 B.n89 585
R1407 B.n496 B.n495 585
R1408 B.n497 B.n88 585
R1409 B.n499 B.n498 585
R1410 B.n500 B.n87 585
R1411 B.n502 B.n501 585
R1412 B.n503 B.n86 585
R1413 B.n505 B.n504 585
R1414 B.n506 B.n85 585
R1415 B.n508 B.n507 585
R1416 B.n509 B.n84 585
R1417 B.n511 B.n510 585
R1418 B.n512 B.n83 585
R1419 B.n700 B.n699 585
R1420 B.n698 B.n17 585
R1421 B.n697 B.n696 585
R1422 B.n695 B.n18 585
R1423 B.n694 B.n693 585
R1424 B.n692 B.n19 585
R1425 B.n691 B.n690 585
R1426 B.n689 B.n20 585
R1427 B.n688 B.n687 585
R1428 B.n686 B.n21 585
R1429 B.n685 B.n684 585
R1430 B.n683 B.n22 585
R1431 B.n682 B.n681 585
R1432 B.n680 B.n23 585
R1433 B.n679 B.n678 585
R1434 B.n677 B.n24 585
R1435 B.n676 B.n675 585
R1436 B.n674 B.n25 585
R1437 B.n673 B.n672 585
R1438 B.n671 B.n26 585
R1439 B.n670 B.n669 585
R1440 B.n668 B.n27 585
R1441 B.n667 B.n666 585
R1442 B.n665 B.n28 585
R1443 B.n664 B.n663 585
R1444 B.n662 B.n29 585
R1445 B.n661 B.n660 585
R1446 B.n659 B.n30 585
R1447 B.n658 B.n657 585
R1448 B.n656 B.n31 585
R1449 B.n655 B.n654 585
R1450 B.n653 B.n32 585
R1451 B.n652 B.n651 585
R1452 B.n650 B.n33 585
R1453 B.n649 B.n648 585
R1454 B.n647 B.n34 585
R1455 B.n646 B.n645 585
R1456 B.n644 B.n35 585
R1457 B.n643 B.n642 585
R1458 B.n641 B.n36 585
R1459 B.n640 B.n639 585
R1460 B.n638 B.n37 585
R1461 B.n637 B.n636 585
R1462 B.n635 B.n38 585
R1463 B.n634 B.n633 585
R1464 B.n632 B.n39 585
R1465 B.n631 B.n630 585
R1466 B.n629 B.n40 585
R1467 B.n628 B.n627 585
R1468 B.n626 B.n41 585
R1469 B.n625 B.n624 585
R1470 B.n623 B.n42 585
R1471 B.n622 B.n621 585
R1472 B.n620 B.n43 585
R1473 B.n619 B.n618 585
R1474 B.n617 B.n44 585
R1475 B.n616 B.n615 585
R1476 B.n613 B.n45 585
R1477 B.n612 B.n611 585
R1478 B.n610 B.n48 585
R1479 B.n609 B.n608 585
R1480 B.n607 B.n49 585
R1481 B.n606 B.n605 585
R1482 B.n604 B.n50 585
R1483 B.n603 B.n602 585
R1484 B.n601 B.n51 585
R1485 B.n600 B.n599 585
R1486 B.n598 B.n597 585
R1487 B.n596 B.n55 585
R1488 B.n595 B.n594 585
R1489 B.n593 B.n56 585
R1490 B.n592 B.n591 585
R1491 B.n590 B.n57 585
R1492 B.n589 B.n588 585
R1493 B.n587 B.n58 585
R1494 B.n586 B.n585 585
R1495 B.n584 B.n59 585
R1496 B.n583 B.n582 585
R1497 B.n581 B.n60 585
R1498 B.n580 B.n579 585
R1499 B.n578 B.n61 585
R1500 B.n577 B.n576 585
R1501 B.n575 B.n62 585
R1502 B.n574 B.n573 585
R1503 B.n572 B.n63 585
R1504 B.n571 B.n570 585
R1505 B.n569 B.n64 585
R1506 B.n568 B.n567 585
R1507 B.n566 B.n65 585
R1508 B.n565 B.n564 585
R1509 B.n563 B.n66 585
R1510 B.n562 B.n561 585
R1511 B.n560 B.n67 585
R1512 B.n559 B.n558 585
R1513 B.n557 B.n68 585
R1514 B.n556 B.n555 585
R1515 B.n554 B.n69 585
R1516 B.n553 B.n552 585
R1517 B.n551 B.n70 585
R1518 B.n550 B.n549 585
R1519 B.n548 B.n71 585
R1520 B.n547 B.n546 585
R1521 B.n545 B.n72 585
R1522 B.n544 B.n543 585
R1523 B.n542 B.n73 585
R1524 B.n541 B.n540 585
R1525 B.n539 B.n74 585
R1526 B.n538 B.n537 585
R1527 B.n536 B.n75 585
R1528 B.n535 B.n534 585
R1529 B.n533 B.n76 585
R1530 B.n532 B.n531 585
R1531 B.n530 B.n77 585
R1532 B.n529 B.n528 585
R1533 B.n527 B.n78 585
R1534 B.n526 B.n525 585
R1535 B.n524 B.n79 585
R1536 B.n523 B.n522 585
R1537 B.n521 B.n80 585
R1538 B.n520 B.n519 585
R1539 B.n518 B.n81 585
R1540 B.n517 B.n516 585
R1541 B.n515 B.n82 585
R1542 B.n514 B.n513 585
R1543 B.n701 B.n16 585
R1544 B.n703 B.n702 585
R1545 B.n704 B.n15 585
R1546 B.n706 B.n705 585
R1547 B.n707 B.n14 585
R1548 B.n709 B.n708 585
R1549 B.n710 B.n13 585
R1550 B.n712 B.n711 585
R1551 B.n713 B.n12 585
R1552 B.n715 B.n714 585
R1553 B.n716 B.n11 585
R1554 B.n718 B.n717 585
R1555 B.n719 B.n10 585
R1556 B.n721 B.n720 585
R1557 B.n722 B.n9 585
R1558 B.n724 B.n723 585
R1559 B.n725 B.n8 585
R1560 B.n727 B.n726 585
R1561 B.n728 B.n7 585
R1562 B.n730 B.n729 585
R1563 B.n731 B.n6 585
R1564 B.n733 B.n732 585
R1565 B.n734 B.n5 585
R1566 B.n736 B.n735 585
R1567 B.n737 B.n4 585
R1568 B.n739 B.n738 585
R1569 B.n740 B.n3 585
R1570 B.n742 B.n741 585
R1571 B.n743 B.n0 585
R1572 B.n2 B.n1 585
R1573 B.n192 B.n191 585
R1574 B.n193 B.n190 585
R1575 B.n195 B.n194 585
R1576 B.n196 B.n189 585
R1577 B.n198 B.n197 585
R1578 B.n199 B.n188 585
R1579 B.n201 B.n200 585
R1580 B.n202 B.n187 585
R1581 B.n204 B.n203 585
R1582 B.n205 B.n186 585
R1583 B.n207 B.n206 585
R1584 B.n208 B.n185 585
R1585 B.n210 B.n209 585
R1586 B.n211 B.n184 585
R1587 B.n213 B.n212 585
R1588 B.n214 B.n183 585
R1589 B.n216 B.n215 585
R1590 B.n217 B.n182 585
R1591 B.n219 B.n218 585
R1592 B.n220 B.n181 585
R1593 B.n222 B.n221 585
R1594 B.n223 B.n180 585
R1595 B.n225 B.n224 585
R1596 B.n226 B.n179 585
R1597 B.n228 B.n227 585
R1598 B.n229 B.n178 585
R1599 B.n231 B.n230 585
R1600 B.n232 B.n177 585
R1601 B.n317 B.t6 574.193
R1602 B.n142 B.t3 574.193
R1603 B.n52 B.t9 574.193
R1604 B.n46 B.t0 574.193
R1605 B.n234 B.n177 545.355
R1606 B.n424 B.n113 545.355
R1607 B.n514 B.n83 545.355
R1608 B.n701 B.n700 545.355
R1609 B.n142 B.t4 500.471
R1610 B.n52 B.t11 500.471
R1611 B.n317 B.t7 500.471
R1612 B.n46 B.t2 500.471
R1613 B.n143 B.t5 472.156
R1614 B.n53 B.t10 472.156
R1615 B.n318 B.t8 472.156
R1616 B.n47 B.t1 472.156
R1617 B.n745 B.n744 256.663
R1618 B.n744 B.n743 235.042
R1619 B.n744 B.n2 235.042
R1620 B.n235 B.n234 163.367
R1621 B.n236 B.n235 163.367
R1622 B.n236 B.n175 163.367
R1623 B.n240 B.n175 163.367
R1624 B.n241 B.n240 163.367
R1625 B.n242 B.n241 163.367
R1626 B.n242 B.n173 163.367
R1627 B.n246 B.n173 163.367
R1628 B.n247 B.n246 163.367
R1629 B.n248 B.n247 163.367
R1630 B.n248 B.n171 163.367
R1631 B.n252 B.n171 163.367
R1632 B.n253 B.n252 163.367
R1633 B.n254 B.n253 163.367
R1634 B.n254 B.n169 163.367
R1635 B.n258 B.n169 163.367
R1636 B.n259 B.n258 163.367
R1637 B.n260 B.n259 163.367
R1638 B.n260 B.n167 163.367
R1639 B.n264 B.n167 163.367
R1640 B.n265 B.n264 163.367
R1641 B.n266 B.n265 163.367
R1642 B.n266 B.n165 163.367
R1643 B.n270 B.n165 163.367
R1644 B.n271 B.n270 163.367
R1645 B.n272 B.n271 163.367
R1646 B.n272 B.n163 163.367
R1647 B.n276 B.n163 163.367
R1648 B.n277 B.n276 163.367
R1649 B.n278 B.n277 163.367
R1650 B.n278 B.n161 163.367
R1651 B.n282 B.n161 163.367
R1652 B.n283 B.n282 163.367
R1653 B.n284 B.n283 163.367
R1654 B.n284 B.n159 163.367
R1655 B.n288 B.n159 163.367
R1656 B.n289 B.n288 163.367
R1657 B.n290 B.n289 163.367
R1658 B.n290 B.n157 163.367
R1659 B.n294 B.n157 163.367
R1660 B.n295 B.n294 163.367
R1661 B.n296 B.n295 163.367
R1662 B.n296 B.n155 163.367
R1663 B.n300 B.n155 163.367
R1664 B.n301 B.n300 163.367
R1665 B.n302 B.n301 163.367
R1666 B.n302 B.n153 163.367
R1667 B.n306 B.n153 163.367
R1668 B.n307 B.n306 163.367
R1669 B.n308 B.n307 163.367
R1670 B.n308 B.n151 163.367
R1671 B.n312 B.n151 163.367
R1672 B.n313 B.n312 163.367
R1673 B.n314 B.n313 163.367
R1674 B.n314 B.n149 163.367
R1675 B.n321 B.n149 163.367
R1676 B.n322 B.n321 163.367
R1677 B.n323 B.n322 163.367
R1678 B.n323 B.n147 163.367
R1679 B.n327 B.n147 163.367
R1680 B.n328 B.n327 163.367
R1681 B.n329 B.n328 163.367
R1682 B.n329 B.n145 163.367
R1683 B.n333 B.n145 163.367
R1684 B.n334 B.n333 163.367
R1685 B.n335 B.n334 163.367
R1686 B.n335 B.n141 163.367
R1687 B.n340 B.n141 163.367
R1688 B.n341 B.n340 163.367
R1689 B.n342 B.n341 163.367
R1690 B.n342 B.n139 163.367
R1691 B.n346 B.n139 163.367
R1692 B.n347 B.n346 163.367
R1693 B.n348 B.n347 163.367
R1694 B.n348 B.n137 163.367
R1695 B.n352 B.n137 163.367
R1696 B.n353 B.n352 163.367
R1697 B.n354 B.n353 163.367
R1698 B.n354 B.n135 163.367
R1699 B.n358 B.n135 163.367
R1700 B.n359 B.n358 163.367
R1701 B.n360 B.n359 163.367
R1702 B.n360 B.n133 163.367
R1703 B.n364 B.n133 163.367
R1704 B.n365 B.n364 163.367
R1705 B.n366 B.n365 163.367
R1706 B.n366 B.n131 163.367
R1707 B.n370 B.n131 163.367
R1708 B.n371 B.n370 163.367
R1709 B.n372 B.n371 163.367
R1710 B.n372 B.n129 163.367
R1711 B.n376 B.n129 163.367
R1712 B.n377 B.n376 163.367
R1713 B.n378 B.n377 163.367
R1714 B.n378 B.n127 163.367
R1715 B.n382 B.n127 163.367
R1716 B.n383 B.n382 163.367
R1717 B.n384 B.n383 163.367
R1718 B.n384 B.n125 163.367
R1719 B.n388 B.n125 163.367
R1720 B.n389 B.n388 163.367
R1721 B.n390 B.n389 163.367
R1722 B.n390 B.n123 163.367
R1723 B.n394 B.n123 163.367
R1724 B.n395 B.n394 163.367
R1725 B.n396 B.n395 163.367
R1726 B.n396 B.n121 163.367
R1727 B.n400 B.n121 163.367
R1728 B.n401 B.n400 163.367
R1729 B.n402 B.n401 163.367
R1730 B.n402 B.n119 163.367
R1731 B.n406 B.n119 163.367
R1732 B.n407 B.n406 163.367
R1733 B.n408 B.n407 163.367
R1734 B.n408 B.n117 163.367
R1735 B.n412 B.n117 163.367
R1736 B.n413 B.n412 163.367
R1737 B.n414 B.n413 163.367
R1738 B.n414 B.n115 163.367
R1739 B.n418 B.n115 163.367
R1740 B.n419 B.n418 163.367
R1741 B.n420 B.n419 163.367
R1742 B.n420 B.n113 163.367
R1743 B.n510 B.n83 163.367
R1744 B.n510 B.n509 163.367
R1745 B.n509 B.n508 163.367
R1746 B.n508 B.n85 163.367
R1747 B.n504 B.n85 163.367
R1748 B.n504 B.n503 163.367
R1749 B.n503 B.n502 163.367
R1750 B.n502 B.n87 163.367
R1751 B.n498 B.n87 163.367
R1752 B.n498 B.n497 163.367
R1753 B.n497 B.n496 163.367
R1754 B.n496 B.n89 163.367
R1755 B.n492 B.n89 163.367
R1756 B.n492 B.n491 163.367
R1757 B.n491 B.n490 163.367
R1758 B.n490 B.n91 163.367
R1759 B.n486 B.n91 163.367
R1760 B.n486 B.n485 163.367
R1761 B.n485 B.n484 163.367
R1762 B.n484 B.n93 163.367
R1763 B.n480 B.n93 163.367
R1764 B.n480 B.n479 163.367
R1765 B.n479 B.n478 163.367
R1766 B.n478 B.n95 163.367
R1767 B.n474 B.n95 163.367
R1768 B.n474 B.n473 163.367
R1769 B.n473 B.n472 163.367
R1770 B.n472 B.n97 163.367
R1771 B.n468 B.n97 163.367
R1772 B.n468 B.n467 163.367
R1773 B.n467 B.n466 163.367
R1774 B.n466 B.n99 163.367
R1775 B.n462 B.n99 163.367
R1776 B.n462 B.n461 163.367
R1777 B.n461 B.n460 163.367
R1778 B.n460 B.n101 163.367
R1779 B.n456 B.n101 163.367
R1780 B.n456 B.n455 163.367
R1781 B.n455 B.n454 163.367
R1782 B.n454 B.n103 163.367
R1783 B.n450 B.n103 163.367
R1784 B.n450 B.n449 163.367
R1785 B.n449 B.n448 163.367
R1786 B.n448 B.n105 163.367
R1787 B.n444 B.n105 163.367
R1788 B.n444 B.n443 163.367
R1789 B.n443 B.n442 163.367
R1790 B.n442 B.n107 163.367
R1791 B.n438 B.n107 163.367
R1792 B.n438 B.n437 163.367
R1793 B.n437 B.n436 163.367
R1794 B.n436 B.n109 163.367
R1795 B.n432 B.n109 163.367
R1796 B.n432 B.n431 163.367
R1797 B.n431 B.n430 163.367
R1798 B.n430 B.n111 163.367
R1799 B.n426 B.n111 163.367
R1800 B.n426 B.n425 163.367
R1801 B.n425 B.n424 163.367
R1802 B.n700 B.n17 163.367
R1803 B.n696 B.n17 163.367
R1804 B.n696 B.n695 163.367
R1805 B.n695 B.n694 163.367
R1806 B.n694 B.n19 163.367
R1807 B.n690 B.n19 163.367
R1808 B.n690 B.n689 163.367
R1809 B.n689 B.n688 163.367
R1810 B.n688 B.n21 163.367
R1811 B.n684 B.n21 163.367
R1812 B.n684 B.n683 163.367
R1813 B.n683 B.n682 163.367
R1814 B.n682 B.n23 163.367
R1815 B.n678 B.n23 163.367
R1816 B.n678 B.n677 163.367
R1817 B.n677 B.n676 163.367
R1818 B.n676 B.n25 163.367
R1819 B.n672 B.n25 163.367
R1820 B.n672 B.n671 163.367
R1821 B.n671 B.n670 163.367
R1822 B.n670 B.n27 163.367
R1823 B.n666 B.n27 163.367
R1824 B.n666 B.n665 163.367
R1825 B.n665 B.n664 163.367
R1826 B.n664 B.n29 163.367
R1827 B.n660 B.n29 163.367
R1828 B.n660 B.n659 163.367
R1829 B.n659 B.n658 163.367
R1830 B.n658 B.n31 163.367
R1831 B.n654 B.n31 163.367
R1832 B.n654 B.n653 163.367
R1833 B.n653 B.n652 163.367
R1834 B.n652 B.n33 163.367
R1835 B.n648 B.n33 163.367
R1836 B.n648 B.n647 163.367
R1837 B.n647 B.n646 163.367
R1838 B.n646 B.n35 163.367
R1839 B.n642 B.n35 163.367
R1840 B.n642 B.n641 163.367
R1841 B.n641 B.n640 163.367
R1842 B.n640 B.n37 163.367
R1843 B.n636 B.n37 163.367
R1844 B.n636 B.n635 163.367
R1845 B.n635 B.n634 163.367
R1846 B.n634 B.n39 163.367
R1847 B.n630 B.n39 163.367
R1848 B.n630 B.n629 163.367
R1849 B.n629 B.n628 163.367
R1850 B.n628 B.n41 163.367
R1851 B.n624 B.n41 163.367
R1852 B.n624 B.n623 163.367
R1853 B.n623 B.n622 163.367
R1854 B.n622 B.n43 163.367
R1855 B.n618 B.n43 163.367
R1856 B.n618 B.n617 163.367
R1857 B.n617 B.n616 163.367
R1858 B.n616 B.n45 163.367
R1859 B.n611 B.n45 163.367
R1860 B.n611 B.n610 163.367
R1861 B.n610 B.n609 163.367
R1862 B.n609 B.n49 163.367
R1863 B.n605 B.n49 163.367
R1864 B.n605 B.n604 163.367
R1865 B.n604 B.n603 163.367
R1866 B.n603 B.n51 163.367
R1867 B.n599 B.n51 163.367
R1868 B.n599 B.n598 163.367
R1869 B.n598 B.n55 163.367
R1870 B.n594 B.n55 163.367
R1871 B.n594 B.n593 163.367
R1872 B.n593 B.n592 163.367
R1873 B.n592 B.n57 163.367
R1874 B.n588 B.n57 163.367
R1875 B.n588 B.n587 163.367
R1876 B.n587 B.n586 163.367
R1877 B.n586 B.n59 163.367
R1878 B.n582 B.n59 163.367
R1879 B.n582 B.n581 163.367
R1880 B.n581 B.n580 163.367
R1881 B.n580 B.n61 163.367
R1882 B.n576 B.n61 163.367
R1883 B.n576 B.n575 163.367
R1884 B.n575 B.n574 163.367
R1885 B.n574 B.n63 163.367
R1886 B.n570 B.n63 163.367
R1887 B.n570 B.n569 163.367
R1888 B.n569 B.n568 163.367
R1889 B.n568 B.n65 163.367
R1890 B.n564 B.n65 163.367
R1891 B.n564 B.n563 163.367
R1892 B.n563 B.n562 163.367
R1893 B.n562 B.n67 163.367
R1894 B.n558 B.n67 163.367
R1895 B.n558 B.n557 163.367
R1896 B.n557 B.n556 163.367
R1897 B.n556 B.n69 163.367
R1898 B.n552 B.n69 163.367
R1899 B.n552 B.n551 163.367
R1900 B.n551 B.n550 163.367
R1901 B.n550 B.n71 163.367
R1902 B.n546 B.n71 163.367
R1903 B.n546 B.n545 163.367
R1904 B.n545 B.n544 163.367
R1905 B.n544 B.n73 163.367
R1906 B.n540 B.n73 163.367
R1907 B.n540 B.n539 163.367
R1908 B.n539 B.n538 163.367
R1909 B.n538 B.n75 163.367
R1910 B.n534 B.n75 163.367
R1911 B.n534 B.n533 163.367
R1912 B.n533 B.n532 163.367
R1913 B.n532 B.n77 163.367
R1914 B.n528 B.n77 163.367
R1915 B.n528 B.n527 163.367
R1916 B.n527 B.n526 163.367
R1917 B.n526 B.n79 163.367
R1918 B.n522 B.n79 163.367
R1919 B.n522 B.n521 163.367
R1920 B.n521 B.n520 163.367
R1921 B.n520 B.n81 163.367
R1922 B.n516 B.n81 163.367
R1923 B.n516 B.n515 163.367
R1924 B.n515 B.n514 163.367
R1925 B.n702 B.n701 163.367
R1926 B.n702 B.n15 163.367
R1927 B.n706 B.n15 163.367
R1928 B.n707 B.n706 163.367
R1929 B.n708 B.n707 163.367
R1930 B.n708 B.n13 163.367
R1931 B.n712 B.n13 163.367
R1932 B.n713 B.n712 163.367
R1933 B.n714 B.n713 163.367
R1934 B.n714 B.n11 163.367
R1935 B.n718 B.n11 163.367
R1936 B.n719 B.n718 163.367
R1937 B.n720 B.n719 163.367
R1938 B.n720 B.n9 163.367
R1939 B.n724 B.n9 163.367
R1940 B.n725 B.n724 163.367
R1941 B.n726 B.n725 163.367
R1942 B.n726 B.n7 163.367
R1943 B.n730 B.n7 163.367
R1944 B.n731 B.n730 163.367
R1945 B.n732 B.n731 163.367
R1946 B.n732 B.n5 163.367
R1947 B.n736 B.n5 163.367
R1948 B.n737 B.n736 163.367
R1949 B.n738 B.n737 163.367
R1950 B.n738 B.n3 163.367
R1951 B.n742 B.n3 163.367
R1952 B.n743 B.n742 163.367
R1953 B.n192 B.n2 163.367
R1954 B.n193 B.n192 163.367
R1955 B.n194 B.n193 163.367
R1956 B.n194 B.n189 163.367
R1957 B.n198 B.n189 163.367
R1958 B.n199 B.n198 163.367
R1959 B.n200 B.n199 163.367
R1960 B.n200 B.n187 163.367
R1961 B.n204 B.n187 163.367
R1962 B.n205 B.n204 163.367
R1963 B.n206 B.n205 163.367
R1964 B.n206 B.n185 163.367
R1965 B.n210 B.n185 163.367
R1966 B.n211 B.n210 163.367
R1967 B.n212 B.n211 163.367
R1968 B.n212 B.n183 163.367
R1969 B.n216 B.n183 163.367
R1970 B.n217 B.n216 163.367
R1971 B.n218 B.n217 163.367
R1972 B.n218 B.n181 163.367
R1973 B.n222 B.n181 163.367
R1974 B.n223 B.n222 163.367
R1975 B.n224 B.n223 163.367
R1976 B.n224 B.n179 163.367
R1977 B.n228 B.n179 163.367
R1978 B.n229 B.n228 163.367
R1979 B.n230 B.n229 163.367
R1980 B.n230 B.n177 163.367
R1981 B.n319 B.n318 59.5399
R1982 B.n337 B.n143 59.5399
R1983 B.n54 B.n53 59.5399
R1984 B.n614 B.n47 59.5399
R1985 B.n699 B.n16 35.4346
R1986 B.n513 B.n512 35.4346
R1987 B.n233 B.n232 35.4346
R1988 B.n423 B.n422 35.4346
R1989 B.n318 B.n317 28.3157
R1990 B.n143 B.n142 28.3157
R1991 B.n53 B.n52 28.3157
R1992 B.n47 B.n46 28.3157
R1993 B B.n745 18.0485
R1994 B.n703 B.n16 10.6151
R1995 B.n704 B.n703 10.6151
R1996 B.n705 B.n704 10.6151
R1997 B.n705 B.n14 10.6151
R1998 B.n709 B.n14 10.6151
R1999 B.n710 B.n709 10.6151
R2000 B.n711 B.n710 10.6151
R2001 B.n711 B.n12 10.6151
R2002 B.n715 B.n12 10.6151
R2003 B.n716 B.n715 10.6151
R2004 B.n717 B.n716 10.6151
R2005 B.n717 B.n10 10.6151
R2006 B.n721 B.n10 10.6151
R2007 B.n722 B.n721 10.6151
R2008 B.n723 B.n722 10.6151
R2009 B.n723 B.n8 10.6151
R2010 B.n727 B.n8 10.6151
R2011 B.n728 B.n727 10.6151
R2012 B.n729 B.n728 10.6151
R2013 B.n729 B.n6 10.6151
R2014 B.n733 B.n6 10.6151
R2015 B.n734 B.n733 10.6151
R2016 B.n735 B.n734 10.6151
R2017 B.n735 B.n4 10.6151
R2018 B.n739 B.n4 10.6151
R2019 B.n740 B.n739 10.6151
R2020 B.n741 B.n740 10.6151
R2021 B.n741 B.n0 10.6151
R2022 B.n699 B.n698 10.6151
R2023 B.n698 B.n697 10.6151
R2024 B.n697 B.n18 10.6151
R2025 B.n693 B.n18 10.6151
R2026 B.n693 B.n692 10.6151
R2027 B.n692 B.n691 10.6151
R2028 B.n691 B.n20 10.6151
R2029 B.n687 B.n20 10.6151
R2030 B.n687 B.n686 10.6151
R2031 B.n686 B.n685 10.6151
R2032 B.n685 B.n22 10.6151
R2033 B.n681 B.n22 10.6151
R2034 B.n681 B.n680 10.6151
R2035 B.n680 B.n679 10.6151
R2036 B.n679 B.n24 10.6151
R2037 B.n675 B.n24 10.6151
R2038 B.n675 B.n674 10.6151
R2039 B.n674 B.n673 10.6151
R2040 B.n673 B.n26 10.6151
R2041 B.n669 B.n26 10.6151
R2042 B.n669 B.n668 10.6151
R2043 B.n668 B.n667 10.6151
R2044 B.n667 B.n28 10.6151
R2045 B.n663 B.n28 10.6151
R2046 B.n663 B.n662 10.6151
R2047 B.n662 B.n661 10.6151
R2048 B.n661 B.n30 10.6151
R2049 B.n657 B.n30 10.6151
R2050 B.n657 B.n656 10.6151
R2051 B.n656 B.n655 10.6151
R2052 B.n655 B.n32 10.6151
R2053 B.n651 B.n32 10.6151
R2054 B.n651 B.n650 10.6151
R2055 B.n650 B.n649 10.6151
R2056 B.n649 B.n34 10.6151
R2057 B.n645 B.n34 10.6151
R2058 B.n645 B.n644 10.6151
R2059 B.n644 B.n643 10.6151
R2060 B.n643 B.n36 10.6151
R2061 B.n639 B.n36 10.6151
R2062 B.n639 B.n638 10.6151
R2063 B.n638 B.n637 10.6151
R2064 B.n637 B.n38 10.6151
R2065 B.n633 B.n38 10.6151
R2066 B.n633 B.n632 10.6151
R2067 B.n632 B.n631 10.6151
R2068 B.n631 B.n40 10.6151
R2069 B.n627 B.n40 10.6151
R2070 B.n627 B.n626 10.6151
R2071 B.n626 B.n625 10.6151
R2072 B.n625 B.n42 10.6151
R2073 B.n621 B.n42 10.6151
R2074 B.n621 B.n620 10.6151
R2075 B.n620 B.n619 10.6151
R2076 B.n619 B.n44 10.6151
R2077 B.n615 B.n44 10.6151
R2078 B.n613 B.n612 10.6151
R2079 B.n612 B.n48 10.6151
R2080 B.n608 B.n48 10.6151
R2081 B.n608 B.n607 10.6151
R2082 B.n607 B.n606 10.6151
R2083 B.n606 B.n50 10.6151
R2084 B.n602 B.n50 10.6151
R2085 B.n602 B.n601 10.6151
R2086 B.n601 B.n600 10.6151
R2087 B.n597 B.n596 10.6151
R2088 B.n596 B.n595 10.6151
R2089 B.n595 B.n56 10.6151
R2090 B.n591 B.n56 10.6151
R2091 B.n591 B.n590 10.6151
R2092 B.n590 B.n589 10.6151
R2093 B.n589 B.n58 10.6151
R2094 B.n585 B.n58 10.6151
R2095 B.n585 B.n584 10.6151
R2096 B.n584 B.n583 10.6151
R2097 B.n583 B.n60 10.6151
R2098 B.n579 B.n60 10.6151
R2099 B.n579 B.n578 10.6151
R2100 B.n578 B.n577 10.6151
R2101 B.n577 B.n62 10.6151
R2102 B.n573 B.n62 10.6151
R2103 B.n573 B.n572 10.6151
R2104 B.n572 B.n571 10.6151
R2105 B.n571 B.n64 10.6151
R2106 B.n567 B.n64 10.6151
R2107 B.n567 B.n566 10.6151
R2108 B.n566 B.n565 10.6151
R2109 B.n565 B.n66 10.6151
R2110 B.n561 B.n66 10.6151
R2111 B.n561 B.n560 10.6151
R2112 B.n560 B.n559 10.6151
R2113 B.n559 B.n68 10.6151
R2114 B.n555 B.n68 10.6151
R2115 B.n555 B.n554 10.6151
R2116 B.n554 B.n553 10.6151
R2117 B.n553 B.n70 10.6151
R2118 B.n549 B.n70 10.6151
R2119 B.n549 B.n548 10.6151
R2120 B.n548 B.n547 10.6151
R2121 B.n547 B.n72 10.6151
R2122 B.n543 B.n72 10.6151
R2123 B.n543 B.n542 10.6151
R2124 B.n542 B.n541 10.6151
R2125 B.n541 B.n74 10.6151
R2126 B.n537 B.n74 10.6151
R2127 B.n537 B.n536 10.6151
R2128 B.n536 B.n535 10.6151
R2129 B.n535 B.n76 10.6151
R2130 B.n531 B.n76 10.6151
R2131 B.n531 B.n530 10.6151
R2132 B.n530 B.n529 10.6151
R2133 B.n529 B.n78 10.6151
R2134 B.n525 B.n78 10.6151
R2135 B.n525 B.n524 10.6151
R2136 B.n524 B.n523 10.6151
R2137 B.n523 B.n80 10.6151
R2138 B.n519 B.n80 10.6151
R2139 B.n519 B.n518 10.6151
R2140 B.n518 B.n517 10.6151
R2141 B.n517 B.n82 10.6151
R2142 B.n513 B.n82 10.6151
R2143 B.n512 B.n511 10.6151
R2144 B.n511 B.n84 10.6151
R2145 B.n507 B.n84 10.6151
R2146 B.n507 B.n506 10.6151
R2147 B.n506 B.n505 10.6151
R2148 B.n505 B.n86 10.6151
R2149 B.n501 B.n86 10.6151
R2150 B.n501 B.n500 10.6151
R2151 B.n500 B.n499 10.6151
R2152 B.n499 B.n88 10.6151
R2153 B.n495 B.n88 10.6151
R2154 B.n495 B.n494 10.6151
R2155 B.n494 B.n493 10.6151
R2156 B.n493 B.n90 10.6151
R2157 B.n489 B.n90 10.6151
R2158 B.n489 B.n488 10.6151
R2159 B.n488 B.n487 10.6151
R2160 B.n487 B.n92 10.6151
R2161 B.n483 B.n92 10.6151
R2162 B.n483 B.n482 10.6151
R2163 B.n482 B.n481 10.6151
R2164 B.n481 B.n94 10.6151
R2165 B.n477 B.n94 10.6151
R2166 B.n477 B.n476 10.6151
R2167 B.n476 B.n475 10.6151
R2168 B.n475 B.n96 10.6151
R2169 B.n471 B.n96 10.6151
R2170 B.n471 B.n470 10.6151
R2171 B.n470 B.n469 10.6151
R2172 B.n469 B.n98 10.6151
R2173 B.n465 B.n98 10.6151
R2174 B.n465 B.n464 10.6151
R2175 B.n464 B.n463 10.6151
R2176 B.n463 B.n100 10.6151
R2177 B.n459 B.n100 10.6151
R2178 B.n459 B.n458 10.6151
R2179 B.n458 B.n457 10.6151
R2180 B.n457 B.n102 10.6151
R2181 B.n453 B.n102 10.6151
R2182 B.n453 B.n452 10.6151
R2183 B.n452 B.n451 10.6151
R2184 B.n451 B.n104 10.6151
R2185 B.n447 B.n104 10.6151
R2186 B.n447 B.n446 10.6151
R2187 B.n446 B.n445 10.6151
R2188 B.n445 B.n106 10.6151
R2189 B.n441 B.n106 10.6151
R2190 B.n441 B.n440 10.6151
R2191 B.n440 B.n439 10.6151
R2192 B.n439 B.n108 10.6151
R2193 B.n435 B.n108 10.6151
R2194 B.n435 B.n434 10.6151
R2195 B.n434 B.n433 10.6151
R2196 B.n433 B.n110 10.6151
R2197 B.n429 B.n110 10.6151
R2198 B.n429 B.n428 10.6151
R2199 B.n428 B.n427 10.6151
R2200 B.n427 B.n112 10.6151
R2201 B.n423 B.n112 10.6151
R2202 B.n191 B.n1 10.6151
R2203 B.n191 B.n190 10.6151
R2204 B.n195 B.n190 10.6151
R2205 B.n196 B.n195 10.6151
R2206 B.n197 B.n196 10.6151
R2207 B.n197 B.n188 10.6151
R2208 B.n201 B.n188 10.6151
R2209 B.n202 B.n201 10.6151
R2210 B.n203 B.n202 10.6151
R2211 B.n203 B.n186 10.6151
R2212 B.n207 B.n186 10.6151
R2213 B.n208 B.n207 10.6151
R2214 B.n209 B.n208 10.6151
R2215 B.n209 B.n184 10.6151
R2216 B.n213 B.n184 10.6151
R2217 B.n214 B.n213 10.6151
R2218 B.n215 B.n214 10.6151
R2219 B.n215 B.n182 10.6151
R2220 B.n219 B.n182 10.6151
R2221 B.n220 B.n219 10.6151
R2222 B.n221 B.n220 10.6151
R2223 B.n221 B.n180 10.6151
R2224 B.n225 B.n180 10.6151
R2225 B.n226 B.n225 10.6151
R2226 B.n227 B.n226 10.6151
R2227 B.n227 B.n178 10.6151
R2228 B.n231 B.n178 10.6151
R2229 B.n232 B.n231 10.6151
R2230 B.n233 B.n176 10.6151
R2231 B.n237 B.n176 10.6151
R2232 B.n238 B.n237 10.6151
R2233 B.n239 B.n238 10.6151
R2234 B.n239 B.n174 10.6151
R2235 B.n243 B.n174 10.6151
R2236 B.n244 B.n243 10.6151
R2237 B.n245 B.n244 10.6151
R2238 B.n245 B.n172 10.6151
R2239 B.n249 B.n172 10.6151
R2240 B.n250 B.n249 10.6151
R2241 B.n251 B.n250 10.6151
R2242 B.n251 B.n170 10.6151
R2243 B.n255 B.n170 10.6151
R2244 B.n256 B.n255 10.6151
R2245 B.n257 B.n256 10.6151
R2246 B.n257 B.n168 10.6151
R2247 B.n261 B.n168 10.6151
R2248 B.n262 B.n261 10.6151
R2249 B.n263 B.n262 10.6151
R2250 B.n263 B.n166 10.6151
R2251 B.n267 B.n166 10.6151
R2252 B.n268 B.n267 10.6151
R2253 B.n269 B.n268 10.6151
R2254 B.n269 B.n164 10.6151
R2255 B.n273 B.n164 10.6151
R2256 B.n274 B.n273 10.6151
R2257 B.n275 B.n274 10.6151
R2258 B.n275 B.n162 10.6151
R2259 B.n279 B.n162 10.6151
R2260 B.n280 B.n279 10.6151
R2261 B.n281 B.n280 10.6151
R2262 B.n281 B.n160 10.6151
R2263 B.n285 B.n160 10.6151
R2264 B.n286 B.n285 10.6151
R2265 B.n287 B.n286 10.6151
R2266 B.n287 B.n158 10.6151
R2267 B.n291 B.n158 10.6151
R2268 B.n292 B.n291 10.6151
R2269 B.n293 B.n292 10.6151
R2270 B.n293 B.n156 10.6151
R2271 B.n297 B.n156 10.6151
R2272 B.n298 B.n297 10.6151
R2273 B.n299 B.n298 10.6151
R2274 B.n299 B.n154 10.6151
R2275 B.n303 B.n154 10.6151
R2276 B.n304 B.n303 10.6151
R2277 B.n305 B.n304 10.6151
R2278 B.n305 B.n152 10.6151
R2279 B.n309 B.n152 10.6151
R2280 B.n310 B.n309 10.6151
R2281 B.n311 B.n310 10.6151
R2282 B.n311 B.n150 10.6151
R2283 B.n315 B.n150 10.6151
R2284 B.n316 B.n315 10.6151
R2285 B.n320 B.n316 10.6151
R2286 B.n324 B.n148 10.6151
R2287 B.n325 B.n324 10.6151
R2288 B.n326 B.n325 10.6151
R2289 B.n326 B.n146 10.6151
R2290 B.n330 B.n146 10.6151
R2291 B.n331 B.n330 10.6151
R2292 B.n332 B.n331 10.6151
R2293 B.n332 B.n144 10.6151
R2294 B.n336 B.n144 10.6151
R2295 B.n339 B.n338 10.6151
R2296 B.n339 B.n140 10.6151
R2297 B.n343 B.n140 10.6151
R2298 B.n344 B.n343 10.6151
R2299 B.n345 B.n344 10.6151
R2300 B.n345 B.n138 10.6151
R2301 B.n349 B.n138 10.6151
R2302 B.n350 B.n349 10.6151
R2303 B.n351 B.n350 10.6151
R2304 B.n351 B.n136 10.6151
R2305 B.n355 B.n136 10.6151
R2306 B.n356 B.n355 10.6151
R2307 B.n357 B.n356 10.6151
R2308 B.n357 B.n134 10.6151
R2309 B.n361 B.n134 10.6151
R2310 B.n362 B.n361 10.6151
R2311 B.n363 B.n362 10.6151
R2312 B.n363 B.n132 10.6151
R2313 B.n367 B.n132 10.6151
R2314 B.n368 B.n367 10.6151
R2315 B.n369 B.n368 10.6151
R2316 B.n369 B.n130 10.6151
R2317 B.n373 B.n130 10.6151
R2318 B.n374 B.n373 10.6151
R2319 B.n375 B.n374 10.6151
R2320 B.n375 B.n128 10.6151
R2321 B.n379 B.n128 10.6151
R2322 B.n380 B.n379 10.6151
R2323 B.n381 B.n380 10.6151
R2324 B.n381 B.n126 10.6151
R2325 B.n385 B.n126 10.6151
R2326 B.n386 B.n385 10.6151
R2327 B.n387 B.n386 10.6151
R2328 B.n387 B.n124 10.6151
R2329 B.n391 B.n124 10.6151
R2330 B.n392 B.n391 10.6151
R2331 B.n393 B.n392 10.6151
R2332 B.n393 B.n122 10.6151
R2333 B.n397 B.n122 10.6151
R2334 B.n398 B.n397 10.6151
R2335 B.n399 B.n398 10.6151
R2336 B.n399 B.n120 10.6151
R2337 B.n403 B.n120 10.6151
R2338 B.n404 B.n403 10.6151
R2339 B.n405 B.n404 10.6151
R2340 B.n405 B.n118 10.6151
R2341 B.n409 B.n118 10.6151
R2342 B.n410 B.n409 10.6151
R2343 B.n411 B.n410 10.6151
R2344 B.n411 B.n116 10.6151
R2345 B.n415 B.n116 10.6151
R2346 B.n416 B.n415 10.6151
R2347 B.n417 B.n416 10.6151
R2348 B.n417 B.n114 10.6151
R2349 B.n421 B.n114 10.6151
R2350 B.n422 B.n421 10.6151
R2351 B.n615 B.n614 9.36635
R2352 B.n597 B.n54 9.36635
R2353 B.n320 B.n319 9.36635
R2354 B.n338 B.n337 9.36635
R2355 B.n745 B.n0 8.11757
R2356 B.n745 B.n1 8.11757
R2357 B.n614 B.n613 1.24928
R2358 B.n600 B.n54 1.24928
R2359 B.n319 B.n148 1.24928
R2360 B.n337 B.n336 1.24928
R2361 VP.n7 VP.t1 428.428
R2362 VP.n17 VP.t5 405.435
R2363 VP.n29 VP.t6 405.435
R2364 VP.n15 VP.t2 405.435
R2365 VP.n22 VP.t3 370.459
R2366 VP.n1 VP.t0 370.459
R2367 VP.n5 VP.t4 370.459
R2368 VP.n8 VP.t7 370.459
R2369 VP.n9 VP.n6 161.3
R2370 VP.n11 VP.n10 161.3
R2371 VP.n13 VP.n12 161.3
R2372 VP.n14 VP.n4 161.3
R2373 VP.n28 VP.n0 161.3
R2374 VP.n27 VP.n26 161.3
R2375 VP.n25 VP.n24 161.3
R2376 VP.n23 VP.n2 161.3
R2377 VP.n21 VP.n20 161.3
R2378 VP.n19 VP.n3 161.3
R2379 VP.n16 VP.n15 80.6037
R2380 VP.n30 VP.n29 80.6037
R2381 VP.n18 VP.n17 80.6037
R2382 VP.n24 VP.n23 56.5193
R2383 VP.n10 VP.n9 56.5193
R2384 VP.n17 VP.n3 50.4025
R2385 VP.n29 VP.n28 50.4025
R2386 VP.n15 VP.n14 50.4025
R2387 VP.n18 VP.n16 48.2893
R2388 VP.n8 VP.n7 33.6057
R2389 VP.n7 VP.n6 28.1515
R2390 VP.n21 VP.n3 24.4675
R2391 VP.n28 VP.n27 24.4675
R2392 VP.n14 VP.n13 24.4675
R2393 VP.n23 VP.n22 23.4888
R2394 VP.n24 VP.n1 23.4888
R2395 VP.n10 VP.n5 23.4888
R2396 VP.n9 VP.n8 23.4888
R2397 VP.n22 VP.n21 0.97918
R2398 VP.n27 VP.n1 0.97918
R2399 VP.n13 VP.n5 0.97918
R2400 VP.n16 VP.n4 0.285035
R2401 VP.n19 VP.n18 0.285035
R2402 VP.n30 VP.n0 0.285035
R2403 VP.n11 VP.n6 0.189894
R2404 VP.n12 VP.n11 0.189894
R2405 VP.n12 VP.n4 0.189894
R2406 VP.n20 VP.n19 0.189894
R2407 VP.n20 VP.n2 0.189894
R2408 VP.n25 VP.n2 0.189894
R2409 VP.n26 VP.n25 0.189894
R2410 VP.n26 VP.n0 0.189894
R2411 VP VP.n30 0.146778
R2412 VDD1 VDD1.n0 73.3777
R2413 VDD1.n3 VDD1.n2 73.2632
R2414 VDD1.n3 VDD1.n1 73.2632
R2415 VDD1.n5 VDD1.n4 72.6891
R2416 VDD1.n5 VDD1.n3 44.9362
R2417 VDD1.n4 VDD1.t3 1.87183
R2418 VDD1.n4 VDD1.t5 1.87183
R2419 VDD1.n0 VDD1.t6 1.87183
R2420 VDD1.n0 VDD1.t0 1.87183
R2421 VDD1.n2 VDD1.t7 1.87183
R2422 VDD1.n2 VDD1.t1 1.87183
R2423 VDD1.n1 VDD1.t2 1.87183
R2424 VDD1.n1 VDD1.t4 1.87183
R2425 VDD1 VDD1.n5 0.571621
C0 VTAIL VDD1 12.134099f
C1 B VDD1 1.34611f
C2 w_n2430_n4442# VP 4.93664f
C3 VDD1 VDD2 1.04164f
C4 VP VN 6.85701f
C5 w_n2430_n4442# VTAIL 5.4551f
C6 w_n2430_n4442# B 9.37088f
C7 VTAIL VN 9.43763f
C8 B VN 0.945473f
C9 w_n2430_n4442# VDD2 1.65949f
C10 VDD2 VN 9.7241f
C11 w_n2430_n4442# VDD1 1.60662f
C12 VDD1 VN 0.149127f
C13 VTAIL VP 9.451731f
C14 B VP 1.4592f
C15 VDD2 VP 0.363304f
C16 VDD1 VP 9.93762f
C17 w_n2430_n4442# VN 4.62551f
C18 B VTAIL 5.7087f
C19 VTAIL VDD2 12.1786f
C20 B VDD2 1.39608f
C21 VDD2 VSUBS 1.531752f
C22 VDD1 VSUBS 1.911954f
C23 VTAIL VSUBS 1.288669f
C24 VN VSUBS 5.39359f
C25 VP VSUBS 2.301394f
C26 B VSUBS 3.818469f
C27 w_n2430_n4442# VSUBS 0.132066p
C28 VDD1.t6 VSUBS 0.352622f
C29 VDD1.t0 VSUBS 0.352622f
C30 VDD1.n0 VSUBS 2.9489f
C31 VDD1.t2 VSUBS 0.352622f
C32 VDD1.t4 VSUBS 0.352622f
C33 VDD1.n1 VSUBS 2.94784f
C34 VDD1.t7 VSUBS 0.352622f
C35 VDD1.t1 VSUBS 0.352622f
C36 VDD1.n2 VSUBS 2.94784f
C37 VDD1.n3 VSUBS 3.41767f
C38 VDD1.t3 VSUBS 0.352622f
C39 VDD1.t5 VSUBS 0.352622f
C40 VDD1.n4 VSUBS 2.94281f
C41 VDD1.n5 VSUBS 3.22664f
C42 VP.n0 VSUBS 0.056537f
C43 VP.t0 VSUBS 2.28592f
C44 VP.n1 VSUBS 0.815867f
C45 VP.n2 VSUBS 0.04237f
C46 VP.t3 VSUBS 2.28592f
C47 VP.n3 VSUBS 0.055085f
C48 VP.n4 VSUBS 0.056537f
C49 VP.t2 VSUBS 2.35927f
C50 VP.t4 VSUBS 2.28592f
C51 VP.n5 VSUBS 0.815867f
C52 VP.n6 VSUBS 0.22306f
C53 VP.t7 VSUBS 2.28592f
C54 VP.t1 VSUBS 2.40765f
C55 VP.n7 VSUBS 0.872469f
C56 VP.n8 VSUBS 0.884636f
C57 VP.n9 VSUBS 0.060293f
C58 VP.n10 VSUBS 0.060293f
C59 VP.n11 VSUBS 0.04237f
C60 VP.n12 VSUBS 0.04237f
C61 VP.n13 VSUBS 0.04154f
C62 VP.n14 VSUBS 0.055085f
C63 VP.n15 VSUBS 0.890888f
C64 VP.n16 VSUBS 2.20007f
C65 VP.t5 VSUBS 2.35927f
C66 VP.n17 VSUBS 0.890888f
C67 VP.n18 VSUBS 2.23161f
C68 VP.n19 VSUBS 0.056537f
C69 VP.n20 VSUBS 0.04237f
C70 VP.n21 VSUBS 0.04154f
C71 VP.n22 VSUBS 0.815867f
C72 VP.n23 VSUBS 0.060293f
C73 VP.n24 VSUBS 0.060293f
C74 VP.n25 VSUBS 0.04237f
C75 VP.n26 VSUBS 0.04237f
C76 VP.n27 VSUBS 0.04154f
C77 VP.n28 VSUBS 0.055085f
C78 VP.t6 VSUBS 2.35927f
C79 VP.n29 VSUBS 0.890888f
C80 VP.n30 VSUBS 0.039681f
C81 B.n0 VSUBS 0.006405f
C82 B.n1 VSUBS 0.006405f
C83 B.n2 VSUBS 0.009473f
C84 B.n3 VSUBS 0.007259f
C85 B.n4 VSUBS 0.007259f
C86 B.n5 VSUBS 0.007259f
C87 B.n6 VSUBS 0.007259f
C88 B.n7 VSUBS 0.007259f
C89 B.n8 VSUBS 0.007259f
C90 B.n9 VSUBS 0.007259f
C91 B.n10 VSUBS 0.007259f
C92 B.n11 VSUBS 0.007259f
C93 B.n12 VSUBS 0.007259f
C94 B.n13 VSUBS 0.007259f
C95 B.n14 VSUBS 0.007259f
C96 B.n15 VSUBS 0.007259f
C97 B.n16 VSUBS 0.017636f
C98 B.n17 VSUBS 0.007259f
C99 B.n18 VSUBS 0.007259f
C100 B.n19 VSUBS 0.007259f
C101 B.n20 VSUBS 0.007259f
C102 B.n21 VSUBS 0.007259f
C103 B.n22 VSUBS 0.007259f
C104 B.n23 VSUBS 0.007259f
C105 B.n24 VSUBS 0.007259f
C106 B.n25 VSUBS 0.007259f
C107 B.n26 VSUBS 0.007259f
C108 B.n27 VSUBS 0.007259f
C109 B.n28 VSUBS 0.007259f
C110 B.n29 VSUBS 0.007259f
C111 B.n30 VSUBS 0.007259f
C112 B.n31 VSUBS 0.007259f
C113 B.n32 VSUBS 0.007259f
C114 B.n33 VSUBS 0.007259f
C115 B.n34 VSUBS 0.007259f
C116 B.n35 VSUBS 0.007259f
C117 B.n36 VSUBS 0.007259f
C118 B.n37 VSUBS 0.007259f
C119 B.n38 VSUBS 0.007259f
C120 B.n39 VSUBS 0.007259f
C121 B.n40 VSUBS 0.007259f
C122 B.n41 VSUBS 0.007259f
C123 B.n42 VSUBS 0.007259f
C124 B.n43 VSUBS 0.007259f
C125 B.n44 VSUBS 0.007259f
C126 B.n45 VSUBS 0.007259f
C127 B.t1 VSUBS 0.348116f
C128 B.t2 VSUBS 0.366027f
C129 B.t0 VSUBS 0.849231f
C130 B.n46 VSUBS 0.489811f
C131 B.n47 VSUBS 0.32693f
C132 B.n48 VSUBS 0.007259f
C133 B.n49 VSUBS 0.007259f
C134 B.n50 VSUBS 0.007259f
C135 B.n51 VSUBS 0.007259f
C136 B.t10 VSUBS 0.34812f
C137 B.t11 VSUBS 0.36603f
C138 B.t9 VSUBS 0.849231f
C139 B.n52 VSUBS 0.489808f
C140 B.n53 VSUBS 0.326927f
C141 B.n54 VSUBS 0.016819f
C142 B.n55 VSUBS 0.007259f
C143 B.n56 VSUBS 0.007259f
C144 B.n57 VSUBS 0.007259f
C145 B.n58 VSUBS 0.007259f
C146 B.n59 VSUBS 0.007259f
C147 B.n60 VSUBS 0.007259f
C148 B.n61 VSUBS 0.007259f
C149 B.n62 VSUBS 0.007259f
C150 B.n63 VSUBS 0.007259f
C151 B.n64 VSUBS 0.007259f
C152 B.n65 VSUBS 0.007259f
C153 B.n66 VSUBS 0.007259f
C154 B.n67 VSUBS 0.007259f
C155 B.n68 VSUBS 0.007259f
C156 B.n69 VSUBS 0.007259f
C157 B.n70 VSUBS 0.007259f
C158 B.n71 VSUBS 0.007259f
C159 B.n72 VSUBS 0.007259f
C160 B.n73 VSUBS 0.007259f
C161 B.n74 VSUBS 0.007259f
C162 B.n75 VSUBS 0.007259f
C163 B.n76 VSUBS 0.007259f
C164 B.n77 VSUBS 0.007259f
C165 B.n78 VSUBS 0.007259f
C166 B.n79 VSUBS 0.007259f
C167 B.n80 VSUBS 0.007259f
C168 B.n81 VSUBS 0.007259f
C169 B.n82 VSUBS 0.007259f
C170 B.n83 VSUBS 0.017636f
C171 B.n84 VSUBS 0.007259f
C172 B.n85 VSUBS 0.007259f
C173 B.n86 VSUBS 0.007259f
C174 B.n87 VSUBS 0.007259f
C175 B.n88 VSUBS 0.007259f
C176 B.n89 VSUBS 0.007259f
C177 B.n90 VSUBS 0.007259f
C178 B.n91 VSUBS 0.007259f
C179 B.n92 VSUBS 0.007259f
C180 B.n93 VSUBS 0.007259f
C181 B.n94 VSUBS 0.007259f
C182 B.n95 VSUBS 0.007259f
C183 B.n96 VSUBS 0.007259f
C184 B.n97 VSUBS 0.007259f
C185 B.n98 VSUBS 0.007259f
C186 B.n99 VSUBS 0.007259f
C187 B.n100 VSUBS 0.007259f
C188 B.n101 VSUBS 0.007259f
C189 B.n102 VSUBS 0.007259f
C190 B.n103 VSUBS 0.007259f
C191 B.n104 VSUBS 0.007259f
C192 B.n105 VSUBS 0.007259f
C193 B.n106 VSUBS 0.007259f
C194 B.n107 VSUBS 0.007259f
C195 B.n108 VSUBS 0.007259f
C196 B.n109 VSUBS 0.007259f
C197 B.n110 VSUBS 0.007259f
C198 B.n111 VSUBS 0.007259f
C199 B.n112 VSUBS 0.007259f
C200 B.n113 VSUBS 0.018234f
C201 B.n114 VSUBS 0.007259f
C202 B.n115 VSUBS 0.007259f
C203 B.n116 VSUBS 0.007259f
C204 B.n117 VSUBS 0.007259f
C205 B.n118 VSUBS 0.007259f
C206 B.n119 VSUBS 0.007259f
C207 B.n120 VSUBS 0.007259f
C208 B.n121 VSUBS 0.007259f
C209 B.n122 VSUBS 0.007259f
C210 B.n123 VSUBS 0.007259f
C211 B.n124 VSUBS 0.007259f
C212 B.n125 VSUBS 0.007259f
C213 B.n126 VSUBS 0.007259f
C214 B.n127 VSUBS 0.007259f
C215 B.n128 VSUBS 0.007259f
C216 B.n129 VSUBS 0.007259f
C217 B.n130 VSUBS 0.007259f
C218 B.n131 VSUBS 0.007259f
C219 B.n132 VSUBS 0.007259f
C220 B.n133 VSUBS 0.007259f
C221 B.n134 VSUBS 0.007259f
C222 B.n135 VSUBS 0.007259f
C223 B.n136 VSUBS 0.007259f
C224 B.n137 VSUBS 0.007259f
C225 B.n138 VSUBS 0.007259f
C226 B.n139 VSUBS 0.007259f
C227 B.n140 VSUBS 0.007259f
C228 B.n141 VSUBS 0.007259f
C229 B.t5 VSUBS 0.34812f
C230 B.t4 VSUBS 0.36603f
C231 B.t3 VSUBS 0.849231f
C232 B.n142 VSUBS 0.489808f
C233 B.n143 VSUBS 0.326927f
C234 B.n144 VSUBS 0.007259f
C235 B.n145 VSUBS 0.007259f
C236 B.n146 VSUBS 0.007259f
C237 B.n147 VSUBS 0.007259f
C238 B.n148 VSUBS 0.004057f
C239 B.n149 VSUBS 0.007259f
C240 B.n150 VSUBS 0.007259f
C241 B.n151 VSUBS 0.007259f
C242 B.n152 VSUBS 0.007259f
C243 B.n153 VSUBS 0.007259f
C244 B.n154 VSUBS 0.007259f
C245 B.n155 VSUBS 0.007259f
C246 B.n156 VSUBS 0.007259f
C247 B.n157 VSUBS 0.007259f
C248 B.n158 VSUBS 0.007259f
C249 B.n159 VSUBS 0.007259f
C250 B.n160 VSUBS 0.007259f
C251 B.n161 VSUBS 0.007259f
C252 B.n162 VSUBS 0.007259f
C253 B.n163 VSUBS 0.007259f
C254 B.n164 VSUBS 0.007259f
C255 B.n165 VSUBS 0.007259f
C256 B.n166 VSUBS 0.007259f
C257 B.n167 VSUBS 0.007259f
C258 B.n168 VSUBS 0.007259f
C259 B.n169 VSUBS 0.007259f
C260 B.n170 VSUBS 0.007259f
C261 B.n171 VSUBS 0.007259f
C262 B.n172 VSUBS 0.007259f
C263 B.n173 VSUBS 0.007259f
C264 B.n174 VSUBS 0.007259f
C265 B.n175 VSUBS 0.007259f
C266 B.n176 VSUBS 0.007259f
C267 B.n177 VSUBS 0.017636f
C268 B.n178 VSUBS 0.007259f
C269 B.n179 VSUBS 0.007259f
C270 B.n180 VSUBS 0.007259f
C271 B.n181 VSUBS 0.007259f
C272 B.n182 VSUBS 0.007259f
C273 B.n183 VSUBS 0.007259f
C274 B.n184 VSUBS 0.007259f
C275 B.n185 VSUBS 0.007259f
C276 B.n186 VSUBS 0.007259f
C277 B.n187 VSUBS 0.007259f
C278 B.n188 VSUBS 0.007259f
C279 B.n189 VSUBS 0.007259f
C280 B.n190 VSUBS 0.007259f
C281 B.n191 VSUBS 0.007259f
C282 B.n192 VSUBS 0.007259f
C283 B.n193 VSUBS 0.007259f
C284 B.n194 VSUBS 0.007259f
C285 B.n195 VSUBS 0.007259f
C286 B.n196 VSUBS 0.007259f
C287 B.n197 VSUBS 0.007259f
C288 B.n198 VSUBS 0.007259f
C289 B.n199 VSUBS 0.007259f
C290 B.n200 VSUBS 0.007259f
C291 B.n201 VSUBS 0.007259f
C292 B.n202 VSUBS 0.007259f
C293 B.n203 VSUBS 0.007259f
C294 B.n204 VSUBS 0.007259f
C295 B.n205 VSUBS 0.007259f
C296 B.n206 VSUBS 0.007259f
C297 B.n207 VSUBS 0.007259f
C298 B.n208 VSUBS 0.007259f
C299 B.n209 VSUBS 0.007259f
C300 B.n210 VSUBS 0.007259f
C301 B.n211 VSUBS 0.007259f
C302 B.n212 VSUBS 0.007259f
C303 B.n213 VSUBS 0.007259f
C304 B.n214 VSUBS 0.007259f
C305 B.n215 VSUBS 0.007259f
C306 B.n216 VSUBS 0.007259f
C307 B.n217 VSUBS 0.007259f
C308 B.n218 VSUBS 0.007259f
C309 B.n219 VSUBS 0.007259f
C310 B.n220 VSUBS 0.007259f
C311 B.n221 VSUBS 0.007259f
C312 B.n222 VSUBS 0.007259f
C313 B.n223 VSUBS 0.007259f
C314 B.n224 VSUBS 0.007259f
C315 B.n225 VSUBS 0.007259f
C316 B.n226 VSUBS 0.007259f
C317 B.n227 VSUBS 0.007259f
C318 B.n228 VSUBS 0.007259f
C319 B.n229 VSUBS 0.007259f
C320 B.n230 VSUBS 0.007259f
C321 B.n231 VSUBS 0.007259f
C322 B.n232 VSUBS 0.017636f
C323 B.n233 VSUBS 0.018234f
C324 B.n234 VSUBS 0.018234f
C325 B.n235 VSUBS 0.007259f
C326 B.n236 VSUBS 0.007259f
C327 B.n237 VSUBS 0.007259f
C328 B.n238 VSUBS 0.007259f
C329 B.n239 VSUBS 0.007259f
C330 B.n240 VSUBS 0.007259f
C331 B.n241 VSUBS 0.007259f
C332 B.n242 VSUBS 0.007259f
C333 B.n243 VSUBS 0.007259f
C334 B.n244 VSUBS 0.007259f
C335 B.n245 VSUBS 0.007259f
C336 B.n246 VSUBS 0.007259f
C337 B.n247 VSUBS 0.007259f
C338 B.n248 VSUBS 0.007259f
C339 B.n249 VSUBS 0.007259f
C340 B.n250 VSUBS 0.007259f
C341 B.n251 VSUBS 0.007259f
C342 B.n252 VSUBS 0.007259f
C343 B.n253 VSUBS 0.007259f
C344 B.n254 VSUBS 0.007259f
C345 B.n255 VSUBS 0.007259f
C346 B.n256 VSUBS 0.007259f
C347 B.n257 VSUBS 0.007259f
C348 B.n258 VSUBS 0.007259f
C349 B.n259 VSUBS 0.007259f
C350 B.n260 VSUBS 0.007259f
C351 B.n261 VSUBS 0.007259f
C352 B.n262 VSUBS 0.007259f
C353 B.n263 VSUBS 0.007259f
C354 B.n264 VSUBS 0.007259f
C355 B.n265 VSUBS 0.007259f
C356 B.n266 VSUBS 0.007259f
C357 B.n267 VSUBS 0.007259f
C358 B.n268 VSUBS 0.007259f
C359 B.n269 VSUBS 0.007259f
C360 B.n270 VSUBS 0.007259f
C361 B.n271 VSUBS 0.007259f
C362 B.n272 VSUBS 0.007259f
C363 B.n273 VSUBS 0.007259f
C364 B.n274 VSUBS 0.007259f
C365 B.n275 VSUBS 0.007259f
C366 B.n276 VSUBS 0.007259f
C367 B.n277 VSUBS 0.007259f
C368 B.n278 VSUBS 0.007259f
C369 B.n279 VSUBS 0.007259f
C370 B.n280 VSUBS 0.007259f
C371 B.n281 VSUBS 0.007259f
C372 B.n282 VSUBS 0.007259f
C373 B.n283 VSUBS 0.007259f
C374 B.n284 VSUBS 0.007259f
C375 B.n285 VSUBS 0.007259f
C376 B.n286 VSUBS 0.007259f
C377 B.n287 VSUBS 0.007259f
C378 B.n288 VSUBS 0.007259f
C379 B.n289 VSUBS 0.007259f
C380 B.n290 VSUBS 0.007259f
C381 B.n291 VSUBS 0.007259f
C382 B.n292 VSUBS 0.007259f
C383 B.n293 VSUBS 0.007259f
C384 B.n294 VSUBS 0.007259f
C385 B.n295 VSUBS 0.007259f
C386 B.n296 VSUBS 0.007259f
C387 B.n297 VSUBS 0.007259f
C388 B.n298 VSUBS 0.007259f
C389 B.n299 VSUBS 0.007259f
C390 B.n300 VSUBS 0.007259f
C391 B.n301 VSUBS 0.007259f
C392 B.n302 VSUBS 0.007259f
C393 B.n303 VSUBS 0.007259f
C394 B.n304 VSUBS 0.007259f
C395 B.n305 VSUBS 0.007259f
C396 B.n306 VSUBS 0.007259f
C397 B.n307 VSUBS 0.007259f
C398 B.n308 VSUBS 0.007259f
C399 B.n309 VSUBS 0.007259f
C400 B.n310 VSUBS 0.007259f
C401 B.n311 VSUBS 0.007259f
C402 B.n312 VSUBS 0.007259f
C403 B.n313 VSUBS 0.007259f
C404 B.n314 VSUBS 0.007259f
C405 B.n315 VSUBS 0.007259f
C406 B.n316 VSUBS 0.007259f
C407 B.t8 VSUBS 0.348116f
C408 B.t7 VSUBS 0.366027f
C409 B.t6 VSUBS 0.849231f
C410 B.n317 VSUBS 0.489811f
C411 B.n318 VSUBS 0.32693f
C412 B.n319 VSUBS 0.016819f
C413 B.n320 VSUBS 0.006832f
C414 B.n321 VSUBS 0.007259f
C415 B.n322 VSUBS 0.007259f
C416 B.n323 VSUBS 0.007259f
C417 B.n324 VSUBS 0.007259f
C418 B.n325 VSUBS 0.007259f
C419 B.n326 VSUBS 0.007259f
C420 B.n327 VSUBS 0.007259f
C421 B.n328 VSUBS 0.007259f
C422 B.n329 VSUBS 0.007259f
C423 B.n330 VSUBS 0.007259f
C424 B.n331 VSUBS 0.007259f
C425 B.n332 VSUBS 0.007259f
C426 B.n333 VSUBS 0.007259f
C427 B.n334 VSUBS 0.007259f
C428 B.n335 VSUBS 0.007259f
C429 B.n336 VSUBS 0.004057f
C430 B.n337 VSUBS 0.016819f
C431 B.n338 VSUBS 0.006832f
C432 B.n339 VSUBS 0.007259f
C433 B.n340 VSUBS 0.007259f
C434 B.n341 VSUBS 0.007259f
C435 B.n342 VSUBS 0.007259f
C436 B.n343 VSUBS 0.007259f
C437 B.n344 VSUBS 0.007259f
C438 B.n345 VSUBS 0.007259f
C439 B.n346 VSUBS 0.007259f
C440 B.n347 VSUBS 0.007259f
C441 B.n348 VSUBS 0.007259f
C442 B.n349 VSUBS 0.007259f
C443 B.n350 VSUBS 0.007259f
C444 B.n351 VSUBS 0.007259f
C445 B.n352 VSUBS 0.007259f
C446 B.n353 VSUBS 0.007259f
C447 B.n354 VSUBS 0.007259f
C448 B.n355 VSUBS 0.007259f
C449 B.n356 VSUBS 0.007259f
C450 B.n357 VSUBS 0.007259f
C451 B.n358 VSUBS 0.007259f
C452 B.n359 VSUBS 0.007259f
C453 B.n360 VSUBS 0.007259f
C454 B.n361 VSUBS 0.007259f
C455 B.n362 VSUBS 0.007259f
C456 B.n363 VSUBS 0.007259f
C457 B.n364 VSUBS 0.007259f
C458 B.n365 VSUBS 0.007259f
C459 B.n366 VSUBS 0.007259f
C460 B.n367 VSUBS 0.007259f
C461 B.n368 VSUBS 0.007259f
C462 B.n369 VSUBS 0.007259f
C463 B.n370 VSUBS 0.007259f
C464 B.n371 VSUBS 0.007259f
C465 B.n372 VSUBS 0.007259f
C466 B.n373 VSUBS 0.007259f
C467 B.n374 VSUBS 0.007259f
C468 B.n375 VSUBS 0.007259f
C469 B.n376 VSUBS 0.007259f
C470 B.n377 VSUBS 0.007259f
C471 B.n378 VSUBS 0.007259f
C472 B.n379 VSUBS 0.007259f
C473 B.n380 VSUBS 0.007259f
C474 B.n381 VSUBS 0.007259f
C475 B.n382 VSUBS 0.007259f
C476 B.n383 VSUBS 0.007259f
C477 B.n384 VSUBS 0.007259f
C478 B.n385 VSUBS 0.007259f
C479 B.n386 VSUBS 0.007259f
C480 B.n387 VSUBS 0.007259f
C481 B.n388 VSUBS 0.007259f
C482 B.n389 VSUBS 0.007259f
C483 B.n390 VSUBS 0.007259f
C484 B.n391 VSUBS 0.007259f
C485 B.n392 VSUBS 0.007259f
C486 B.n393 VSUBS 0.007259f
C487 B.n394 VSUBS 0.007259f
C488 B.n395 VSUBS 0.007259f
C489 B.n396 VSUBS 0.007259f
C490 B.n397 VSUBS 0.007259f
C491 B.n398 VSUBS 0.007259f
C492 B.n399 VSUBS 0.007259f
C493 B.n400 VSUBS 0.007259f
C494 B.n401 VSUBS 0.007259f
C495 B.n402 VSUBS 0.007259f
C496 B.n403 VSUBS 0.007259f
C497 B.n404 VSUBS 0.007259f
C498 B.n405 VSUBS 0.007259f
C499 B.n406 VSUBS 0.007259f
C500 B.n407 VSUBS 0.007259f
C501 B.n408 VSUBS 0.007259f
C502 B.n409 VSUBS 0.007259f
C503 B.n410 VSUBS 0.007259f
C504 B.n411 VSUBS 0.007259f
C505 B.n412 VSUBS 0.007259f
C506 B.n413 VSUBS 0.007259f
C507 B.n414 VSUBS 0.007259f
C508 B.n415 VSUBS 0.007259f
C509 B.n416 VSUBS 0.007259f
C510 B.n417 VSUBS 0.007259f
C511 B.n418 VSUBS 0.007259f
C512 B.n419 VSUBS 0.007259f
C513 B.n420 VSUBS 0.007259f
C514 B.n421 VSUBS 0.007259f
C515 B.n422 VSUBS 0.017443f
C516 B.n423 VSUBS 0.018427f
C517 B.n424 VSUBS 0.017636f
C518 B.n425 VSUBS 0.007259f
C519 B.n426 VSUBS 0.007259f
C520 B.n427 VSUBS 0.007259f
C521 B.n428 VSUBS 0.007259f
C522 B.n429 VSUBS 0.007259f
C523 B.n430 VSUBS 0.007259f
C524 B.n431 VSUBS 0.007259f
C525 B.n432 VSUBS 0.007259f
C526 B.n433 VSUBS 0.007259f
C527 B.n434 VSUBS 0.007259f
C528 B.n435 VSUBS 0.007259f
C529 B.n436 VSUBS 0.007259f
C530 B.n437 VSUBS 0.007259f
C531 B.n438 VSUBS 0.007259f
C532 B.n439 VSUBS 0.007259f
C533 B.n440 VSUBS 0.007259f
C534 B.n441 VSUBS 0.007259f
C535 B.n442 VSUBS 0.007259f
C536 B.n443 VSUBS 0.007259f
C537 B.n444 VSUBS 0.007259f
C538 B.n445 VSUBS 0.007259f
C539 B.n446 VSUBS 0.007259f
C540 B.n447 VSUBS 0.007259f
C541 B.n448 VSUBS 0.007259f
C542 B.n449 VSUBS 0.007259f
C543 B.n450 VSUBS 0.007259f
C544 B.n451 VSUBS 0.007259f
C545 B.n452 VSUBS 0.007259f
C546 B.n453 VSUBS 0.007259f
C547 B.n454 VSUBS 0.007259f
C548 B.n455 VSUBS 0.007259f
C549 B.n456 VSUBS 0.007259f
C550 B.n457 VSUBS 0.007259f
C551 B.n458 VSUBS 0.007259f
C552 B.n459 VSUBS 0.007259f
C553 B.n460 VSUBS 0.007259f
C554 B.n461 VSUBS 0.007259f
C555 B.n462 VSUBS 0.007259f
C556 B.n463 VSUBS 0.007259f
C557 B.n464 VSUBS 0.007259f
C558 B.n465 VSUBS 0.007259f
C559 B.n466 VSUBS 0.007259f
C560 B.n467 VSUBS 0.007259f
C561 B.n468 VSUBS 0.007259f
C562 B.n469 VSUBS 0.007259f
C563 B.n470 VSUBS 0.007259f
C564 B.n471 VSUBS 0.007259f
C565 B.n472 VSUBS 0.007259f
C566 B.n473 VSUBS 0.007259f
C567 B.n474 VSUBS 0.007259f
C568 B.n475 VSUBS 0.007259f
C569 B.n476 VSUBS 0.007259f
C570 B.n477 VSUBS 0.007259f
C571 B.n478 VSUBS 0.007259f
C572 B.n479 VSUBS 0.007259f
C573 B.n480 VSUBS 0.007259f
C574 B.n481 VSUBS 0.007259f
C575 B.n482 VSUBS 0.007259f
C576 B.n483 VSUBS 0.007259f
C577 B.n484 VSUBS 0.007259f
C578 B.n485 VSUBS 0.007259f
C579 B.n486 VSUBS 0.007259f
C580 B.n487 VSUBS 0.007259f
C581 B.n488 VSUBS 0.007259f
C582 B.n489 VSUBS 0.007259f
C583 B.n490 VSUBS 0.007259f
C584 B.n491 VSUBS 0.007259f
C585 B.n492 VSUBS 0.007259f
C586 B.n493 VSUBS 0.007259f
C587 B.n494 VSUBS 0.007259f
C588 B.n495 VSUBS 0.007259f
C589 B.n496 VSUBS 0.007259f
C590 B.n497 VSUBS 0.007259f
C591 B.n498 VSUBS 0.007259f
C592 B.n499 VSUBS 0.007259f
C593 B.n500 VSUBS 0.007259f
C594 B.n501 VSUBS 0.007259f
C595 B.n502 VSUBS 0.007259f
C596 B.n503 VSUBS 0.007259f
C597 B.n504 VSUBS 0.007259f
C598 B.n505 VSUBS 0.007259f
C599 B.n506 VSUBS 0.007259f
C600 B.n507 VSUBS 0.007259f
C601 B.n508 VSUBS 0.007259f
C602 B.n509 VSUBS 0.007259f
C603 B.n510 VSUBS 0.007259f
C604 B.n511 VSUBS 0.007259f
C605 B.n512 VSUBS 0.017636f
C606 B.n513 VSUBS 0.018234f
C607 B.n514 VSUBS 0.018234f
C608 B.n515 VSUBS 0.007259f
C609 B.n516 VSUBS 0.007259f
C610 B.n517 VSUBS 0.007259f
C611 B.n518 VSUBS 0.007259f
C612 B.n519 VSUBS 0.007259f
C613 B.n520 VSUBS 0.007259f
C614 B.n521 VSUBS 0.007259f
C615 B.n522 VSUBS 0.007259f
C616 B.n523 VSUBS 0.007259f
C617 B.n524 VSUBS 0.007259f
C618 B.n525 VSUBS 0.007259f
C619 B.n526 VSUBS 0.007259f
C620 B.n527 VSUBS 0.007259f
C621 B.n528 VSUBS 0.007259f
C622 B.n529 VSUBS 0.007259f
C623 B.n530 VSUBS 0.007259f
C624 B.n531 VSUBS 0.007259f
C625 B.n532 VSUBS 0.007259f
C626 B.n533 VSUBS 0.007259f
C627 B.n534 VSUBS 0.007259f
C628 B.n535 VSUBS 0.007259f
C629 B.n536 VSUBS 0.007259f
C630 B.n537 VSUBS 0.007259f
C631 B.n538 VSUBS 0.007259f
C632 B.n539 VSUBS 0.007259f
C633 B.n540 VSUBS 0.007259f
C634 B.n541 VSUBS 0.007259f
C635 B.n542 VSUBS 0.007259f
C636 B.n543 VSUBS 0.007259f
C637 B.n544 VSUBS 0.007259f
C638 B.n545 VSUBS 0.007259f
C639 B.n546 VSUBS 0.007259f
C640 B.n547 VSUBS 0.007259f
C641 B.n548 VSUBS 0.007259f
C642 B.n549 VSUBS 0.007259f
C643 B.n550 VSUBS 0.007259f
C644 B.n551 VSUBS 0.007259f
C645 B.n552 VSUBS 0.007259f
C646 B.n553 VSUBS 0.007259f
C647 B.n554 VSUBS 0.007259f
C648 B.n555 VSUBS 0.007259f
C649 B.n556 VSUBS 0.007259f
C650 B.n557 VSUBS 0.007259f
C651 B.n558 VSUBS 0.007259f
C652 B.n559 VSUBS 0.007259f
C653 B.n560 VSUBS 0.007259f
C654 B.n561 VSUBS 0.007259f
C655 B.n562 VSUBS 0.007259f
C656 B.n563 VSUBS 0.007259f
C657 B.n564 VSUBS 0.007259f
C658 B.n565 VSUBS 0.007259f
C659 B.n566 VSUBS 0.007259f
C660 B.n567 VSUBS 0.007259f
C661 B.n568 VSUBS 0.007259f
C662 B.n569 VSUBS 0.007259f
C663 B.n570 VSUBS 0.007259f
C664 B.n571 VSUBS 0.007259f
C665 B.n572 VSUBS 0.007259f
C666 B.n573 VSUBS 0.007259f
C667 B.n574 VSUBS 0.007259f
C668 B.n575 VSUBS 0.007259f
C669 B.n576 VSUBS 0.007259f
C670 B.n577 VSUBS 0.007259f
C671 B.n578 VSUBS 0.007259f
C672 B.n579 VSUBS 0.007259f
C673 B.n580 VSUBS 0.007259f
C674 B.n581 VSUBS 0.007259f
C675 B.n582 VSUBS 0.007259f
C676 B.n583 VSUBS 0.007259f
C677 B.n584 VSUBS 0.007259f
C678 B.n585 VSUBS 0.007259f
C679 B.n586 VSUBS 0.007259f
C680 B.n587 VSUBS 0.007259f
C681 B.n588 VSUBS 0.007259f
C682 B.n589 VSUBS 0.007259f
C683 B.n590 VSUBS 0.007259f
C684 B.n591 VSUBS 0.007259f
C685 B.n592 VSUBS 0.007259f
C686 B.n593 VSUBS 0.007259f
C687 B.n594 VSUBS 0.007259f
C688 B.n595 VSUBS 0.007259f
C689 B.n596 VSUBS 0.007259f
C690 B.n597 VSUBS 0.006832f
C691 B.n598 VSUBS 0.007259f
C692 B.n599 VSUBS 0.007259f
C693 B.n600 VSUBS 0.004057f
C694 B.n601 VSUBS 0.007259f
C695 B.n602 VSUBS 0.007259f
C696 B.n603 VSUBS 0.007259f
C697 B.n604 VSUBS 0.007259f
C698 B.n605 VSUBS 0.007259f
C699 B.n606 VSUBS 0.007259f
C700 B.n607 VSUBS 0.007259f
C701 B.n608 VSUBS 0.007259f
C702 B.n609 VSUBS 0.007259f
C703 B.n610 VSUBS 0.007259f
C704 B.n611 VSUBS 0.007259f
C705 B.n612 VSUBS 0.007259f
C706 B.n613 VSUBS 0.004057f
C707 B.n614 VSUBS 0.016819f
C708 B.n615 VSUBS 0.006832f
C709 B.n616 VSUBS 0.007259f
C710 B.n617 VSUBS 0.007259f
C711 B.n618 VSUBS 0.007259f
C712 B.n619 VSUBS 0.007259f
C713 B.n620 VSUBS 0.007259f
C714 B.n621 VSUBS 0.007259f
C715 B.n622 VSUBS 0.007259f
C716 B.n623 VSUBS 0.007259f
C717 B.n624 VSUBS 0.007259f
C718 B.n625 VSUBS 0.007259f
C719 B.n626 VSUBS 0.007259f
C720 B.n627 VSUBS 0.007259f
C721 B.n628 VSUBS 0.007259f
C722 B.n629 VSUBS 0.007259f
C723 B.n630 VSUBS 0.007259f
C724 B.n631 VSUBS 0.007259f
C725 B.n632 VSUBS 0.007259f
C726 B.n633 VSUBS 0.007259f
C727 B.n634 VSUBS 0.007259f
C728 B.n635 VSUBS 0.007259f
C729 B.n636 VSUBS 0.007259f
C730 B.n637 VSUBS 0.007259f
C731 B.n638 VSUBS 0.007259f
C732 B.n639 VSUBS 0.007259f
C733 B.n640 VSUBS 0.007259f
C734 B.n641 VSUBS 0.007259f
C735 B.n642 VSUBS 0.007259f
C736 B.n643 VSUBS 0.007259f
C737 B.n644 VSUBS 0.007259f
C738 B.n645 VSUBS 0.007259f
C739 B.n646 VSUBS 0.007259f
C740 B.n647 VSUBS 0.007259f
C741 B.n648 VSUBS 0.007259f
C742 B.n649 VSUBS 0.007259f
C743 B.n650 VSUBS 0.007259f
C744 B.n651 VSUBS 0.007259f
C745 B.n652 VSUBS 0.007259f
C746 B.n653 VSUBS 0.007259f
C747 B.n654 VSUBS 0.007259f
C748 B.n655 VSUBS 0.007259f
C749 B.n656 VSUBS 0.007259f
C750 B.n657 VSUBS 0.007259f
C751 B.n658 VSUBS 0.007259f
C752 B.n659 VSUBS 0.007259f
C753 B.n660 VSUBS 0.007259f
C754 B.n661 VSUBS 0.007259f
C755 B.n662 VSUBS 0.007259f
C756 B.n663 VSUBS 0.007259f
C757 B.n664 VSUBS 0.007259f
C758 B.n665 VSUBS 0.007259f
C759 B.n666 VSUBS 0.007259f
C760 B.n667 VSUBS 0.007259f
C761 B.n668 VSUBS 0.007259f
C762 B.n669 VSUBS 0.007259f
C763 B.n670 VSUBS 0.007259f
C764 B.n671 VSUBS 0.007259f
C765 B.n672 VSUBS 0.007259f
C766 B.n673 VSUBS 0.007259f
C767 B.n674 VSUBS 0.007259f
C768 B.n675 VSUBS 0.007259f
C769 B.n676 VSUBS 0.007259f
C770 B.n677 VSUBS 0.007259f
C771 B.n678 VSUBS 0.007259f
C772 B.n679 VSUBS 0.007259f
C773 B.n680 VSUBS 0.007259f
C774 B.n681 VSUBS 0.007259f
C775 B.n682 VSUBS 0.007259f
C776 B.n683 VSUBS 0.007259f
C777 B.n684 VSUBS 0.007259f
C778 B.n685 VSUBS 0.007259f
C779 B.n686 VSUBS 0.007259f
C780 B.n687 VSUBS 0.007259f
C781 B.n688 VSUBS 0.007259f
C782 B.n689 VSUBS 0.007259f
C783 B.n690 VSUBS 0.007259f
C784 B.n691 VSUBS 0.007259f
C785 B.n692 VSUBS 0.007259f
C786 B.n693 VSUBS 0.007259f
C787 B.n694 VSUBS 0.007259f
C788 B.n695 VSUBS 0.007259f
C789 B.n696 VSUBS 0.007259f
C790 B.n697 VSUBS 0.007259f
C791 B.n698 VSUBS 0.007259f
C792 B.n699 VSUBS 0.018234f
C793 B.n700 VSUBS 0.018234f
C794 B.n701 VSUBS 0.017636f
C795 B.n702 VSUBS 0.007259f
C796 B.n703 VSUBS 0.007259f
C797 B.n704 VSUBS 0.007259f
C798 B.n705 VSUBS 0.007259f
C799 B.n706 VSUBS 0.007259f
C800 B.n707 VSUBS 0.007259f
C801 B.n708 VSUBS 0.007259f
C802 B.n709 VSUBS 0.007259f
C803 B.n710 VSUBS 0.007259f
C804 B.n711 VSUBS 0.007259f
C805 B.n712 VSUBS 0.007259f
C806 B.n713 VSUBS 0.007259f
C807 B.n714 VSUBS 0.007259f
C808 B.n715 VSUBS 0.007259f
C809 B.n716 VSUBS 0.007259f
C810 B.n717 VSUBS 0.007259f
C811 B.n718 VSUBS 0.007259f
C812 B.n719 VSUBS 0.007259f
C813 B.n720 VSUBS 0.007259f
C814 B.n721 VSUBS 0.007259f
C815 B.n722 VSUBS 0.007259f
C816 B.n723 VSUBS 0.007259f
C817 B.n724 VSUBS 0.007259f
C818 B.n725 VSUBS 0.007259f
C819 B.n726 VSUBS 0.007259f
C820 B.n727 VSUBS 0.007259f
C821 B.n728 VSUBS 0.007259f
C822 B.n729 VSUBS 0.007259f
C823 B.n730 VSUBS 0.007259f
C824 B.n731 VSUBS 0.007259f
C825 B.n732 VSUBS 0.007259f
C826 B.n733 VSUBS 0.007259f
C827 B.n734 VSUBS 0.007259f
C828 B.n735 VSUBS 0.007259f
C829 B.n736 VSUBS 0.007259f
C830 B.n737 VSUBS 0.007259f
C831 B.n738 VSUBS 0.007259f
C832 B.n739 VSUBS 0.007259f
C833 B.n740 VSUBS 0.007259f
C834 B.n741 VSUBS 0.007259f
C835 B.n742 VSUBS 0.007259f
C836 B.n743 VSUBS 0.009473f
C837 B.n744 VSUBS 0.010091f
C838 B.n745 VSUBS 0.020068f
C839 VDD2.t1 VSUBS 0.352539f
C840 VDD2.t7 VSUBS 0.352539f
C841 VDD2.n0 VSUBS 2.94715f
C842 VDD2.t5 VSUBS 0.352539f
C843 VDD2.t3 VSUBS 0.352539f
C844 VDD2.n1 VSUBS 2.94715f
C845 VDD2.n2 VSUBS 3.3627f
C846 VDD2.t2 VSUBS 0.352539f
C847 VDD2.t0 VSUBS 0.352539f
C848 VDD2.n3 VSUBS 2.94213f
C849 VDD2.n4 VSUBS 3.19481f
C850 VDD2.t6 VSUBS 0.352539f
C851 VDD2.t4 VSUBS 0.352539f
C852 VDD2.n5 VSUBS 2.9471f
C853 VTAIL.t11 VSUBS 0.321123f
C854 VTAIL.t8 VSUBS 0.321123f
C855 VTAIL.n0 VSUBS 2.5517f
C856 VTAIL.n1 VSUBS 0.63083f
C857 VTAIL.n2 VSUBS 0.013195f
C858 VTAIL.n3 VSUBS 0.029714f
C859 VTAIL.n4 VSUBS 0.013311f
C860 VTAIL.n5 VSUBS 0.023395f
C861 VTAIL.n6 VSUBS 0.012571f
C862 VTAIL.n7 VSUBS 0.029714f
C863 VTAIL.n8 VSUBS 0.013311f
C864 VTAIL.n9 VSUBS 0.023395f
C865 VTAIL.n10 VSUBS 0.012571f
C866 VTAIL.n11 VSUBS 0.029714f
C867 VTAIL.n12 VSUBS 0.013311f
C868 VTAIL.n13 VSUBS 0.023395f
C869 VTAIL.n14 VSUBS 0.012571f
C870 VTAIL.n15 VSUBS 0.029714f
C871 VTAIL.n16 VSUBS 0.013311f
C872 VTAIL.n17 VSUBS 0.023395f
C873 VTAIL.n18 VSUBS 0.012571f
C874 VTAIL.n19 VSUBS 0.029714f
C875 VTAIL.n20 VSUBS 0.013311f
C876 VTAIL.n21 VSUBS 0.023395f
C877 VTAIL.n22 VSUBS 0.012941f
C878 VTAIL.n23 VSUBS 0.029714f
C879 VTAIL.n24 VSUBS 0.013311f
C880 VTAIL.n25 VSUBS 0.023395f
C881 VTAIL.n26 VSUBS 0.012571f
C882 VTAIL.n27 VSUBS 0.029714f
C883 VTAIL.n28 VSUBS 0.013311f
C884 VTAIL.n29 VSUBS 0.023395f
C885 VTAIL.n30 VSUBS 0.012571f
C886 VTAIL.n31 VSUBS 0.022286f
C887 VTAIL.n32 VSUBS 0.022352f
C888 VTAIL.t10 VSUBS 0.064453f
C889 VTAIL.n33 VSUBS 0.24105f
C890 VTAIL.n34 VSUBS 1.69992f
C891 VTAIL.n35 VSUBS 0.012571f
C892 VTAIL.n36 VSUBS 0.013311f
C893 VTAIL.n37 VSUBS 0.029714f
C894 VTAIL.n38 VSUBS 0.029714f
C895 VTAIL.n39 VSUBS 0.013311f
C896 VTAIL.n40 VSUBS 0.012571f
C897 VTAIL.n41 VSUBS 0.023395f
C898 VTAIL.n42 VSUBS 0.023395f
C899 VTAIL.n43 VSUBS 0.012571f
C900 VTAIL.n44 VSUBS 0.013311f
C901 VTAIL.n45 VSUBS 0.029714f
C902 VTAIL.n46 VSUBS 0.029714f
C903 VTAIL.n47 VSUBS 0.013311f
C904 VTAIL.n48 VSUBS 0.012571f
C905 VTAIL.n49 VSUBS 0.023395f
C906 VTAIL.n50 VSUBS 0.023395f
C907 VTAIL.n51 VSUBS 0.012571f
C908 VTAIL.n52 VSUBS 0.012571f
C909 VTAIL.n53 VSUBS 0.013311f
C910 VTAIL.n54 VSUBS 0.029714f
C911 VTAIL.n55 VSUBS 0.029714f
C912 VTAIL.n56 VSUBS 0.029714f
C913 VTAIL.n57 VSUBS 0.012941f
C914 VTAIL.n58 VSUBS 0.012571f
C915 VTAIL.n59 VSUBS 0.023395f
C916 VTAIL.n60 VSUBS 0.023395f
C917 VTAIL.n61 VSUBS 0.012571f
C918 VTAIL.n62 VSUBS 0.013311f
C919 VTAIL.n63 VSUBS 0.029714f
C920 VTAIL.n64 VSUBS 0.029714f
C921 VTAIL.n65 VSUBS 0.013311f
C922 VTAIL.n66 VSUBS 0.012571f
C923 VTAIL.n67 VSUBS 0.023395f
C924 VTAIL.n68 VSUBS 0.023395f
C925 VTAIL.n69 VSUBS 0.012571f
C926 VTAIL.n70 VSUBS 0.013311f
C927 VTAIL.n71 VSUBS 0.029714f
C928 VTAIL.n72 VSUBS 0.029714f
C929 VTAIL.n73 VSUBS 0.013311f
C930 VTAIL.n74 VSUBS 0.012571f
C931 VTAIL.n75 VSUBS 0.023395f
C932 VTAIL.n76 VSUBS 0.023395f
C933 VTAIL.n77 VSUBS 0.012571f
C934 VTAIL.n78 VSUBS 0.013311f
C935 VTAIL.n79 VSUBS 0.029714f
C936 VTAIL.n80 VSUBS 0.029714f
C937 VTAIL.n81 VSUBS 0.013311f
C938 VTAIL.n82 VSUBS 0.012571f
C939 VTAIL.n83 VSUBS 0.023395f
C940 VTAIL.n84 VSUBS 0.023395f
C941 VTAIL.n85 VSUBS 0.012571f
C942 VTAIL.n86 VSUBS 0.013311f
C943 VTAIL.n87 VSUBS 0.029714f
C944 VTAIL.n88 VSUBS 0.029714f
C945 VTAIL.n89 VSUBS 0.013311f
C946 VTAIL.n90 VSUBS 0.012571f
C947 VTAIL.n91 VSUBS 0.023395f
C948 VTAIL.n92 VSUBS 0.060787f
C949 VTAIL.n93 VSUBS 0.012571f
C950 VTAIL.n94 VSUBS 0.013311f
C951 VTAIL.n95 VSUBS 0.065183f
C952 VTAIL.n96 VSUBS 0.044276f
C953 VTAIL.n97 VSUBS 0.152264f
C954 VTAIL.n98 VSUBS 0.013195f
C955 VTAIL.n99 VSUBS 0.029714f
C956 VTAIL.n100 VSUBS 0.013311f
C957 VTAIL.n101 VSUBS 0.023395f
C958 VTAIL.n102 VSUBS 0.012571f
C959 VTAIL.n103 VSUBS 0.029714f
C960 VTAIL.n104 VSUBS 0.013311f
C961 VTAIL.n105 VSUBS 0.023395f
C962 VTAIL.n106 VSUBS 0.012571f
C963 VTAIL.n107 VSUBS 0.029714f
C964 VTAIL.n108 VSUBS 0.013311f
C965 VTAIL.n109 VSUBS 0.023395f
C966 VTAIL.n110 VSUBS 0.012571f
C967 VTAIL.n111 VSUBS 0.029714f
C968 VTAIL.n112 VSUBS 0.013311f
C969 VTAIL.n113 VSUBS 0.023395f
C970 VTAIL.n114 VSUBS 0.012571f
C971 VTAIL.n115 VSUBS 0.029714f
C972 VTAIL.n116 VSUBS 0.013311f
C973 VTAIL.n117 VSUBS 0.023395f
C974 VTAIL.n118 VSUBS 0.012941f
C975 VTAIL.n119 VSUBS 0.029714f
C976 VTAIL.n120 VSUBS 0.013311f
C977 VTAIL.n121 VSUBS 0.023395f
C978 VTAIL.n122 VSUBS 0.012571f
C979 VTAIL.n123 VSUBS 0.029714f
C980 VTAIL.n124 VSUBS 0.013311f
C981 VTAIL.n125 VSUBS 0.023395f
C982 VTAIL.n126 VSUBS 0.012571f
C983 VTAIL.n127 VSUBS 0.022286f
C984 VTAIL.n128 VSUBS 0.022352f
C985 VTAIL.t1 VSUBS 0.064453f
C986 VTAIL.n129 VSUBS 0.24105f
C987 VTAIL.n130 VSUBS 1.69992f
C988 VTAIL.n131 VSUBS 0.012571f
C989 VTAIL.n132 VSUBS 0.013311f
C990 VTAIL.n133 VSUBS 0.029714f
C991 VTAIL.n134 VSUBS 0.029714f
C992 VTAIL.n135 VSUBS 0.013311f
C993 VTAIL.n136 VSUBS 0.012571f
C994 VTAIL.n137 VSUBS 0.023395f
C995 VTAIL.n138 VSUBS 0.023395f
C996 VTAIL.n139 VSUBS 0.012571f
C997 VTAIL.n140 VSUBS 0.013311f
C998 VTAIL.n141 VSUBS 0.029714f
C999 VTAIL.n142 VSUBS 0.029714f
C1000 VTAIL.n143 VSUBS 0.013311f
C1001 VTAIL.n144 VSUBS 0.012571f
C1002 VTAIL.n145 VSUBS 0.023395f
C1003 VTAIL.n146 VSUBS 0.023395f
C1004 VTAIL.n147 VSUBS 0.012571f
C1005 VTAIL.n148 VSUBS 0.012571f
C1006 VTAIL.n149 VSUBS 0.013311f
C1007 VTAIL.n150 VSUBS 0.029714f
C1008 VTAIL.n151 VSUBS 0.029714f
C1009 VTAIL.n152 VSUBS 0.029714f
C1010 VTAIL.n153 VSUBS 0.012941f
C1011 VTAIL.n154 VSUBS 0.012571f
C1012 VTAIL.n155 VSUBS 0.023395f
C1013 VTAIL.n156 VSUBS 0.023395f
C1014 VTAIL.n157 VSUBS 0.012571f
C1015 VTAIL.n158 VSUBS 0.013311f
C1016 VTAIL.n159 VSUBS 0.029714f
C1017 VTAIL.n160 VSUBS 0.029714f
C1018 VTAIL.n161 VSUBS 0.013311f
C1019 VTAIL.n162 VSUBS 0.012571f
C1020 VTAIL.n163 VSUBS 0.023395f
C1021 VTAIL.n164 VSUBS 0.023395f
C1022 VTAIL.n165 VSUBS 0.012571f
C1023 VTAIL.n166 VSUBS 0.013311f
C1024 VTAIL.n167 VSUBS 0.029714f
C1025 VTAIL.n168 VSUBS 0.029714f
C1026 VTAIL.n169 VSUBS 0.013311f
C1027 VTAIL.n170 VSUBS 0.012571f
C1028 VTAIL.n171 VSUBS 0.023395f
C1029 VTAIL.n172 VSUBS 0.023395f
C1030 VTAIL.n173 VSUBS 0.012571f
C1031 VTAIL.n174 VSUBS 0.013311f
C1032 VTAIL.n175 VSUBS 0.029714f
C1033 VTAIL.n176 VSUBS 0.029714f
C1034 VTAIL.n177 VSUBS 0.013311f
C1035 VTAIL.n178 VSUBS 0.012571f
C1036 VTAIL.n179 VSUBS 0.023395f
C1037 VTAIL.n180 VSUBS 0.023395f
C1038 VTAIL.n181 VSUBS 0.012571f
C1039 VTAIL.n182 VSUBS 0.013311f
C1040 VTAIL.n183 VSUBS 0.029714f
C1041 VTAIL.n184 VSUBS 0.029714f
C1042 VTAIL.n185 VSUBS 0.013311f
C1043 VTAIL.n186 VSUBS 0.012571f
C1044 VTAIL.n187 VSUBS 0.023395f
C1045 VTAIL.n188 VSUBS 0.060787f
C1046 VTAIL.n189 VSUBS 0.012571f
C1047 VTAIL.n190 VSUBS 0.013311f
C1048 VTAIL.n191 VSUBS 0.065183f
C1049 VTAIL.n192 VSUBS 0.044276f
C1050 VTAIL.n193 VSUBS 0.152264f
C1051 VTAIL.t0 VSUBS 0.321123f
C1052 VTAIL.t7 VSUBS 0.321123f
C1053 VTAIL.n194 VSUBS 2.5517f
C1054 VTAIL.n195 VSUBS 0.721322f
C1055 VTAIL.n196 VSUBS 0.013195f
C1056 VTAIL.n197 VSUBS 0.029714f
C1057 VTAIL.n198 VSUBS 0.013311f
C1058 VTAIL.n199 VSUBS 0.023395f
C1059 VTAIL.n200 VSUBS 0.012571f
C1060 VTAIL.n201 VSUBS 0.029714f
C1061 VTAIL.n202 VSUBS 0.013311f
C1062 VTAIL.n203 VSUBS 0.023395f
C1063 VTAIL.n204 VSUBS 0.012571f
C1064 VTAIL.n205 VSUBS 0.029714f
C1065 VTAIL.n206 VSUBS 0.013311f
C1066 VTAIL.n207 VSUBS 0.023395f
C1067 VTAIL.n208 VSUBS 0.012571f
C1068 VTAIL.n209 VSUBS 0.029714f
C1069 VTAIL.n210 VSUBS 0.013311f
C1070 VTAIL.n211 VSUBS 0.023395f
C1071 VTAIL.n212 VSUBS 0.012571f
C1072 VTAIL.n213 VSUBS 0.029714f
C1073 VTAIL.n214 VSUBS 0.013311f
C1074 VTAIL.n215 VSUBS 0.023395f
C1075 VTAIL.n216 VSUBS 0.012941f
C1076 VTAIL.n217 VSUBS 0.029714f
C1077 VTAIL.n218 VSUBS 0.013311f
C1078 VTAIL.n219 VSUBS 0.023395f
C1079 VTAIL.n220 VSUBS 0.012571f
C1080 VTAIL.n221 VSUBS 0.029714f
C1081 VTAIL.n222 VSUBS 0.013311f
C1082 VTAIL.n223 VSUBS 0.023395f
C1083 VTAIL.n224 VSUBS 0.012571f
C1084 VTAIL.n225 VSUBS 0.022286f
C1085 VTAIL.n226 VSUBS 0.022352f
C1086 VTAIL.t4 VSUBS 0.064453f
C1087 VTAIL.n227 VSUBS 0.24105f
C1088 VTAIL.n228 VSUBS 1.69992f
C1089 VTAIL.n229 VSUBS 0.012571f
C1090 VTAIL.n230 VSUBS 0.013311f
C1091 VTAIL.n231 VSUBS 0.029714f
C1092 VTAIL.n232 VSUBS 0.029714f
C1093 VTAIL.n233 VSUBS 0.013311f
C1094 VTAIL.n234 VSUBS 0.012571f
C1095 VTAIL.n235 VSUBS 0.023395f
C1096 VTAIL.n236 VSUBS 0.023395f
C1097 VTAIL.n237 VSUBS 0.012571f
C1098 VTAIL.n238 VSUBS 0.013311f
C1099 VTAIL.n239 VSUBS 0.029714f
C1100 VTAIL.n240 VSUBS 0.029714f
C1101 VTAIL.n241 VSUBS 0.013311f
C1102 VTAIL.n242 VSUBS 0.012571f
C1103 VTAIL.n243 VSUBS 0.023395f
C1104 VTAIL.n244 VSUBS 0.023395f
C1105 VTAIL.n245 VSUBS 0.012571f
C1106 VTAIL.n246 VSUBS 0.012571f
C1107 VTAIL.n247 VSUBS 0.013311f
C1108 VTAIL.n248 VSUBS 0.029714f
C1109 VTAIL.n249 VSUBS 0.029714f
C1110 VTAIL.n250 VSUBS 0.029714f
C1111 VTAIL.n251 VSUBS 0.012941f
C1112 VTAIL.n252 VSUBS 0.012571f
C1113 VTAIL.n253 VSUBS 0.023395f
C1114 VTAIL.n254 VSUBS 0.023395f
C1115 VTAIL.n255 VSUBS 0.012571f
C1116 VTAIL.n256 VSUBS 0.013311f
C1117 VTAIL.n257 VSUBS 0.029714f
C1118 VTAIL.n258 VSUBS 0.029714f
C1119 VTAIL.n259 VSUBS 0.013311f
C1120 VTAIL.n260 VSUBS 0.012571f
C1121 VTAIL.n261 VSUBS 0.023395f
C1122 VTAIL.n262 VSUBS 0.023395f
C1123 VTAIL.n263 VSUBS 0.012571f
C1124 VTAIL.n264 VSUBS 0.013311f
C1125 VTAIL.n265 VSUBS 0.029714f
C1126 VTAIL.n266 VSUBS 0.029714f
C1127 VTAIL.n267 VSUBS 0.013311f
C1128 VTAIL.n268 VSUBS 0.012571f
C1129 VTAIL.n269 VSUBS 0.023395f
C1130 VTAIL.n270 VSUBS 0.023395f
C1131 VTAIL.n271 VSUBS 0.012571f
C1132 VTAIL.n272 VSUBS 0.013311f
C1133 VTAIL.n273 VSUBS 0.029714f
C1134 VTAIL.n274 VSUBS 0.029714f
C1135 VTAIL.n275 VSUBS 0.013311f
C1136 VTAIL.n276 VSUBS 0.012571f
C1137 VTAIL.n277 VSUBS 0.023395f
C1138 VTAIL.n278 VSUBS 0.023395f
C1139 VTAIL.n279 VSUBS 0.012571f
C1140 VTAIL.n280 VSUBS 0.013311f
C1141 VTAIL.n281 VSUBS 0.029714f
C1142 VTAIL.n282 VSUBS 0.029714f
C1143 VTAIL.n283 VSUBS 0.013311f
C1144 VTAIL.n284 VSUBS 0.012571f
C1145 VTAIL.n285 VSUBS 0.023395f
C1146 VTAIL.n286 VSUBS 0.060787f
C1147 VTAIL.n287 VSUBS 0.012571f
C1148 VTAIL.n288 VSUBS 0.013311f
C1149 VTAIL.n289 VSUBS 0.065183f
C1150 VTAIL.n290 VSUBS 0.044276f
C1151 VTAIL.n291 VSUBS 1.65831f
C1152 VTAIL.n292 VSUBS 0.013195f
C1153 VTAIL.n293 VSUBS 0.029714f
C1154 VTAIL.n294 VSUBS 0.013311f
C1155 VTAIL.n295 VSUBS 0.023395f
C1156 VTAIL.n296 VSUBS 0.012571f
C1157 VTAIL.n297 VSUBS 0.029714f
C1158 VTAIL.n298 VSUBS 0.013311f
C1159 VTAIL.n299 VSUBS 0.023395f
C1160 VTAIL.n300 VSUBS 0.012571f
C1161 VTAIL.n301 VSUBS 0.029714f
C1162 VTAIL.n302 VSUBS 0.013311f
C1163 VTAIL.n303 VSUBS 0.023395f
C1164 VTAIL.n304 VSUBS 0.012571f
C1165 VTAIL.n305 VSUBS 0.029714f
C1166 VTAIL.n306 VSUBS 0.013311f
C1167 VTAIL.n307 VSUBS 0.023395f
C1168 VTAIL.n308 VSUBS 0.012571f
C1169 VTAIL.n309 VSUBS 0.029714f
C1170 VTAIL.n310 VSUBS 0.013311f
C1171 VTAIL.n311 VSUBS 0.023395f
C1172 VTAIL.n312 VSUBS 0.012941f
C1173 VTAIL.n313 VSUBS 0.029714f
C1174 VTAIL.n314 VSUBS 0.012571f
C1175 VTAIL.n315 VSUBS 0.013311f
C1176 VTAIL.n316 VSUBS 0.023395f
C1177 VTAIL.n317 VSUBS 0.012571f
C1178 VTAIL.n318 VSUBS 0.029714f
C1179 VTAIL.n319 VSUBS 0.013311f
C1180 VTAIL.n320 VSUBS 0.023395f
C1181 VTAIL.n321 VSUBS 0.012571f
C1182 VTAIL.n322 VSUBS 0.022286f
C1183 VTAIL.n323 VSUBS 0.022352f
C1184 VTAIL.t13 VSUBS 0.064453f
C1185 VTAIL.n324 VSUBS 0.24105f
C1186 VTAIL.n325 VSUBS 1.69992f
C1187 VTAIL.n326 VSUBS 0.012571f
C1188 VTAIL.n327 VSUBS 0.013311f
C1189 VTAIL.n328 VSUBS 0.029714f
C1190 VTAIL.n329 VSUBS 0.029714f
C1191 VTAIL.n330 VSUBS 0.013311f
C1192 VTAIL.n331 VSUBS 0.012571f
C1193 VTAIL.n332 VSUBS 0.023395f
C1194 VTAIL.n333 VSUBS 0.023395f
C1195 VTAIL.n334 VSUBS 0.012571f
C1196 VTAIL.n335 VSUBS 0.013311f
C1197 VTAIL.n336 VSUBS 0.029714f
C1198 VTAIL.n337 VSUBS 0.029714f
C1199 VTAIL.n338 VSUBS 0.013311f
C1200 VTAIL.n339 VSUBS 0.012571f
C1201 VTAIL.n340 VSUBS 0.023395f
C1202 VTAIL.n341 VSUBS 0.023395f
C1203 VTAIL.n342 VSUBS 0.012571f
C1204 VTAIL.n343 VSUBS 0.013311f
C1205 VTAIL.n344 VSUBS 0.029714f
C1206 VTAIL.n345 VSUBS 0.029714f
C1207 VTAIL.n346 VSUBS 0.029714f
C1208 VTAIL.n347 VSUBS 0.012941f
C1209 VTAIL.n348 VSUBS 0.012571f
C1210 VTAIL.n349 VSUBS 0.023395f
C1211 VTAIL.n350 VSUBS 0.023395f
C1212 VTAIL.n351 VSUBS 0.012571f
C1213 VTAIL.n352 VSUBS 0.013311f
C1214 VTAIL.n353 VSUBS 0.029714f
C1215 VTAIL.n354 VSUBS 0.029714f
C1216 VTAIL.n355 VSUBS 0.013311f
C1217 VTAIL.n356 VSUBS 0.012571f
C1218 VTAIL.n357 VSUBS 0.023395f
C1219 VTAIL.n358 VSUBS 0.023395f
C1220 VTAIL.n359 VSUBS 0.012571f
C1221 VTAIL.n360 VSUBS 0.013311f
C1222 VTAIL.n361 VSUBS 0.029714f
C1223 VTAIL.n362 VSUBS 0.029714f
C1224 VTAIL.n363 VSUBS 0.013311f
C1225 VTAIL.n364 VSUBS 0.012571f
C1226 VTAIL.n365 VSUBS 0.023395f
C1227 VTAIL.n366 VSUBS 0.023395f
C1228 VTAIL.n367 VSUBS 0.012571f
C1229 VTAIL.n368 VSUBS 0.013311f
C1230 VTAIL.n369 VSUBS 0.029714f
C1231 VTAIL.n370 VSUBS 0.029714f
C1232 VTAIL.n371 VSUBS 0.013311f
C1233 VTAIL.n372 VSUBS 0.012571f
C1234 VTAIL.n373 VSUBS 0.023395f
C1235 VTAIL.n374 VSUBS 0.023395f
C1236 VTAIL.n375 VSUBS 0.012571f
C1237 VTAIL.n376 VSUBS 0.013311f
C1238 VTAIL.n377 VSUBS 0.029714f
C1239 VTAIL.n378 VSUBS 0.029714f
C1240 VTAIL.n379 VSUBS 0.013311f
C1241 VTAIL.n380 VSUBS 0.012571f
C1242 VTAIL.n381 VSUBS 0.023395f
C1243 VTAIL.n382 VSUBS 0.060787f
C1244 VTAIL.n383 VSUBS 0.012571f
C1245 VTAIL.n384 VSUBS 0.013311f
C1246 VTAIL.n385 VSUBS 0.065183f
C1247 VTAIL.n386 VSUBS 0.044276f
C1248 VTAIL.n387 VSUBS 1.65831f
C1249 VTAIL.t15 VSUBS 0.321123f
C1250 VTAIL.t12 VSUBS 0.321123f
C1251 VTAIL.n388 VSUBS 2.5517f
C1252 VTAIL.n389 VSUBS 0.721321f
C1253 VTAIL.n390 VSUBS 0.013195f
C1254 VTAIL.n391 VSUBS 0.029714f
C1255 VTAIL.n392 VSUBS 0.013311f
C1256 VTAIL.n393 VSUBS 0.023395f
C1257 VTAIL.n394 VSUBS 0.012571f
C1258 VTAIL.n395 VSUBS 0.029714f
C1259 VTAIL.n396 VSUBS 0.013311f
C1260 VTAIL.n397 VSUBS 0.023395f
C1261 VTAIL.n398 VSUBS 0.012571f
C1262 VTAIL.n399 VSUBS 0.029714f
C1263 VTAIL.n400 VSUBS 0.013311f
C1264 VTAIL.n401 VSUBS 0.023395f
C1265 VTAIL.n402 VSUBS 0.012571f
C1266 VTAIL.n403 VSUBS 0.029714f
C1267 VTAIL.n404 VSUBS 0.013311f
C1268 VTAIL.n405 VSUBS 0.023395f
C1269 VTAIL.n406 VSUBS 0.012571f
C1270 VTAIL.n407 VSUBS 0.029714f
C1271 VTAIL.n408 VSUBS 0.013311f
C1272 VTAIL.n409 VSUBS 0.023395f
C1273 VTAIL.n410 VSUBS 0.012941f
C1274 VTAIL.n411 VSUBS 0.029714f
C1275 VTAIL.n412 VSUBS 0.012571f
C1276 VTAIL.n413 VSUBS 0.013311f
C1277 VTAIL.n414 VSUBS 0.023395f
C1278 VTAIL.n415 VSUBS 0.012571f
C1279 VTAIL.n416 VSUBS 0.029714f
C1280 VTAIL.n417 VSUBS 0.013311f
C1281 VTAIL.n418 VSUBS 0.023395f
C1282 VTAIL.n419 VSUBS 0.012571f
C1283 VTAIL.n420 VSUBS 0.022286f
C1284 VTAIL.n421 VSUBS 0.022352f
C1285 VTAIL.t9 VSUBS 0.064453f
C1286 VTAIL.n422 VSUBS 0.24105f
C1287 VTAIL.n423 VSUBS 1.69992f
C1288 VTAIL.n424 VSUBS 0.012571f
C1289 VTAIL.n425 VSUBS 0.013311f
C1290 VTAIL.n426 VSUBS 0.029714f
C1291 VTAIL.n427 VSUBS 0.029714f
C1292 VTAIL.n428 VSUBS 0.013311f
C1293 VTAIL.n429 VSUBS 0.012571f
C1294 VTAIL.n430 VSUBS 0.023395f
C1295 VTAIL.n431 VSUBS 0.023395f
C1296 VTAIL.n432 VSUBS 0.012571f
C1297 VTAIL.n433 VSUBS 0.013311f
C1298 VTAIL.n434 VSUBS 0.029714f
C1299 VTAIL.n435 VSUBS 0.029714f
C1300 VTAIL.n436 VSUBS 0.013311f
C1301 VTAIL.n437 VSUBS 0.012571f
C1302 VTAIL.n438 VSUBS 0.023395f
C1303 VTAIL.n439 VSUBS 0.023395f
C1304 VTAIL.n440 VSUBS 0.012571f
C1305 VTAIL.n441 VSUBS 0.013311f
C1306 VTAIL.n442 VSUBS 0.029714f
C1307 VTAIL.n443 VSUBS 0.029714f
C1308 VTAIL.n444 VSUBS 0.029714f
C1309 VTAIL.n445 VSUBS 0.012941f
C1310 VTAIL.n446 VSUBS 0.012571f
C1311 VTAIL.n447 VSUBS 0.023395f
C1312 VTAIL.n448 VSUBS 0.023395f
C1313 VTAIL.n449 VSUBS 0.012571f
C1314 VTAIL.n450 VSUBS 0.013311f
C1315 VTAIL.n451 VSUBS 0.029714f
C1316 VTAIL.n452 VSUBS 0.029714f
C1317 VTAIL.n453 VSUBS 0.013311f
C1318 VTAIL.n454 VSUBS 0.012571f
C1319 VTAIL.n455 VSUBS 0.023395f
C1320 VTAIL.n456 VSUBS 0.023395f
C1321 VTAIL.n457 VSUBS 0.012571f
C1322 VTAIL.n458 VSUBS 0.013311f
C1323 VTAIL.n459 VSUBS 0.029714f
C1324 VTAIL.n460 VSUBS 0.029714f
C1325 VTAIL.n461 VSUBS 0.013311f
C1326 VTAIL.n462 VSUBS 0.012571f
C1327 VTAIL.n463 VSUBS 0.023395f
C1328 VTAIL.n464 VSUBS 0.023395f
C1329 VTAIL.n465 VSUBS 0.012571f
C1330 VTAIL.n466 VSUBS 0.013311f
C1331 VTAIL.n467 VSUBS 0.029714f
C1332 VTAIL.n468 VSUBS 0.029714f
C1333 VTAIL.n469 VSUBS 0.013311f
C1334 VTAIL.n470 VSUBS 0.012571f
C1335 VTAIL.n471 VSUBS 0.023395f
C1336 VTAIL.n472 VSUBS 0.023395f
C1337 VTAIL.n473 VSUBS 0.012571f
C1338 VTAIL.n474 VSUBS 0.013311f
C1339 VTAIL.n475 VSUBS 0.029714f
C1340 VTAIL.n476 VSUBS 0.029714f
C1341 VTAIL.n477 VSUBS 0.013311f
C1342 VTAIL.n478 VSUBS 0.012571f
C1343 VTAIL.n479 VSUBS 0.023395f
C1344 VTAIL.n480 VSUBS 0.060787f
C1345 VTAIL.n481 VSUBS 0.012571f
C1346 VTAIL.n482 VSUBS 0.013311f
C1347 VTAIL.n483 VSUBS 0.065183f
C1348 VTAIL.n484 VSUBS 0.044276f
C1349 VTAIL.n485 VSUBS 0.152264f
C1350 VTAIL.n486 VSUBS 0.013195f
C1351 VTAIL.n487 VSUBS 0.029714f
C1352 VTAIL.n488 VSUBS 0.013311f
C1353 VTAIL.n489 VSUBS 0.023395f
C1354 VTAIL.n490 VSUBS 0.012571f
C1355 VTAIL.n491 VSUBS 0.029714f
C1356 VTAIL.n492 VSUBS 0.013311f
C1357 VTAIL.n493 VSUBS 0.023395f
C1358 VTAIL.n494 VSUBS 0.012571f
C1359 VTAIL.n495 VSUBS 0.029714f
C1360 VTAIL.n496 VSUBS 0.013311f
C1361 VTAIL.n497 VSUBS 0.023395f
C1362 VTAIL.n498 VSUBS 0.012571f
C1363 VTAIL.n499 VSUBS 0.029714f
C1364 VTAIL.n500 VSUBS 0.013311f
C1365 VTAIL.n501 VSUBS 0.023395f
C1366 VTAIL.n502 VSUBS 0.012571f
C1367 VTAIL.n503 VSUBS 0.029714f
C1368 VTAIL.n504 VSUBS 0.013311f
C1369 VTAIL.n505 VSUBS 0.023395f
C1370 VTAIL.n506 VSUBS 0.012941f
C1371 VTAIL.n507 VSUBS 0.029714f
C1372 VTAIL.n508 VSUBS 0.012571f
C1373 VTAIL.n509 VSUBS 0.013311f
C1374 VTAIL.n510 VSUBS 0.023395f
C1375 VTAIL.n511 VSUBS 0.012571f
C1376 VTAIL.n512 VSUBS 0.029714f
C1377 VTAIL.n513 VSUBS 0.013311f
C1378 VTAIL.n514 VSUBS 0.023395f
C1379 VTAIL.n515 VSUBS 0.012571f
C1380 VTAIL.n516 VSUBS 0.022286f
C1381 VTAIL.n517 VSUBS 0.022352f
C1382 VTAIL.t5 VSUBS 0.064453f
C1383 VTAIL.n518 VSUBS 0.24105f
C1384 VTAIL.n519 VSUBS 1.69992f
C1385 VTAIL.n520 VSUBS 0.012571f
C1386 VTAIL.n521 VSUBS 0.013311f
C1387 VTAIL.n522 VSUBS 0.029714f
C1388 VTAIL.n523 VSUBS 0.029714f
C1389 VTAIL.n524 VSUBS 0.013311f
C1390 VTAIL.n525 VSUBS 0.012571f
C1391 VTAIL.n526 VSUBS 0.023395f
C1392 VTAIL.n527 VSUBS 0.023395f
C1393 VTAIL.n528 VSUBS 0.012571f
C1394 VTAIL.n529 VSUBS 0.013311f
C1395 VTAIL.n530 VSUBS 0.029714f
C1396 VTAIL.n531 VSUBS 0.029714f
C1397 VTAIL.n532 VSUBS 0.013311f
C1398 VTAIL.n533 VSUBS 0.012571f
C1399 VTAIL.n534 VSUBS 0.023395f
C1400 VTAIL.n535 VSUBS 0.023395f
C1401 VTAIL.n536 VSUBS 0.012571f
C1402 VTAIL.n537 VSUBS 0.013311f
C1403 VTAIL.n538 VSUBS 0.029714f
C1404 VTAIL.n539 VSUBS 0.029714f
C1405 VTAIL.n540 VSUBS 0.029714f
C1406 VTAIL.n541 VSUBS 0.012941f
C1407 VTAIL.n542 VSUBS 0.012571f
C1408 VTAIL.n543 VSUBS 0.023395f
C1409 VTAIL.n544 VSUBS 0.023395f
C1410 VTAIL.n545 VSUBS 0.012571f
C1411 VTAIL.n546 VSUBS 0.013311f
C1412 VTAIL.n547 VSUBS 0.029714f
C1413 VTAIL.n548 VSUBS 0.029714f
C1414 VTAIL.n549 VSUBS 0.013311f
C1415 VTAIL.n550 VSUBS 0.012571f
C1416 VTAIL.n551 VSUBS 0.023395f
C1417 VTAIL.n552 VSUBS 0.023395f
C1418 VTAIL.n553 VSUBS 0.012571f
C1419 VTAIL.n554 VSUBS 0.013311f
C1420 VTAIL.n555 VSUBS 0.029714f
C1421 VTAIL.n556 VSUBS 0.029714f
C1422 VTAIL.n557 VSUBS 0.013311f
C1423 VTAIL.n558 VSUBS 0.012571f
C1424 VTAIL.n559 VSUBS 0.023395f
C1425 VTAIL.n560 VSUBS 0.023395f
C1426 VTAIL.n561 VSUBS 0.012571f
C1427 VTAIL.n562 VSUBS 0.013311f
C1428 VTAIL.n563 VSUBS 0.029714f
C1429 VTAIL.n564 VSUBS 0.029714f
C1430 VTAIL.n565 VSUBS 0.013311f
C1431 VTAIL.n566 VSUBS 0.012571f
C1432 VTAIL.n567 VSUBS 0.023395f
C1433 VTAIL.n568 VSUBS 0.023395f
C1434 VTAIL.n569 VSUBS 0.012571f
C1435 VTAIL.n570 VSUBS 0.013311f
C1436 VTAIL.n571 VSUBS 0.029714f
C1437 VTAIL.n572 VSUBS 0.029714f
C1438 VTAIL.n573 VSUBS 0.013311f
C1439 VTAIL.n574 VSUBS 0.012571f
C1440 VTAIL.n575 VSUBS 0.023395f
C1441 VTAIL.n576 VSUBS 0.060787f
C1442 VTAIL.n577 VSUBS 0.012571f
C1443 VTAIL.n578 VSUBS 0.013311f
C1444 VTAIL.n579 VSUBS 0.065183f
C1445 VTAIL.n580 VSUBS 0.044276f
C1446 VTAIL.n581 VSUBS 0.152264f
C1447 VTAIL.t3 VSUBS 0.321123f
C1448 VTAIL.t2 VSUBS 0.321123f
C1449 VTAIL.n582 VSUBS 2.5517f
C1450 VTAIL.n583 VSUBS 0.721321f
C1451 VTAIL.n584 VSUBS 0.013195f
C1452 VTAIL.n585 VSUBS 0.029714f
C1453 VTAIL.n586 VSUBS 0.013311f
C1454 VTAIL.n587 VSUBS 0.023395f
C1455 VTAIL.n588 VSUBS 0.012571f
C1456 VTAIL.n589 VSUBS 0.029714f
C1457 VTAIL.n590 VSUBS 0.013311f
C1458 VTAIL.n591 VSUBS 0.023395f
C1459 VTAIL.n592 VSUBS 0.012571f
C1460 VTAIL.n593 VSUBS 0.029714f
C1461 VTAIL.n594 VSUBS 0.013311f
C1462 VTAIL.n595 VSUBS 0.023395f
C1463 VTAIL.n596 VSUBS 0.012571f
C1464 VTAIL.n597 VSUBS 0.029714f
C1465 VTAIL.n598 VSUBS 0.013311f
C1466 VTAIL.n599 VSUBS 0.023395f
C1467 VTAIL.n600 VSUBS 0.012571f
C1468 VTAIL.n601 VSUBS 0.029714f
C1469 VTAIL.n602 VSUBS 0.013311f
C1470 VTAIL.n603 VSUBS 0.023395f
C1471 VTAIL.n604 VSUBS 0.012941f
C1472 VTAIL.n605 VSUBS 0.029714f
C1473 VTAIL.n606 VSUBS 0.012571f
C1474 VTAIL.n607 VSUBS 0.013311f
C1475 VTAIL.n608 VSUBS 0.023395f
C1476 VTAIL.n609 VSUBS 0.012571f
C1477 VTAIL.n610 VSUBS 0.029714f
C1478 VTAIL.n611 VSUBS 0.013311f
C1479 VTAIL.n612 VSUBS 0.023395f
C1480 VTAIL.n613 VSUBS 0.012571f
C1481 VTAIL.n614 VSUBS 0.022286f
C1482 VTAIL.n615 VSUBS 0.022352f
C1483 VTAIL.t6 VSUBS 0.064453f
C1484 VTAIL.n616 VSUBS 0.24105f
C1485 VTAIL.n617 VSUBS 1.69992f
C1486 VTAIL.n618 VSUBS 0.012571f
C1487 VTAIL.n619 VSUBS 0.013311f
C1488 VTAIL.n620 VSUBS 0.029714f
C1489 VTAIL.n621 VSUBS 0.029714f
C1490 VTAIL.n622 VSUBS 0.013311f
C1491 VTAIL.n623 VSUBS 0.012571f
C1492 VTAIL.n624 VSUBS 0.023395f
C1493 VTAIL.n625 VSUBS 0.023395f
C1494 VTAIL.n626 VSUBS 0.012571f
C1495 VTAIL.n627 VSUBS 0.013311f
C1496 VTAIL.n628 VSUBS 0.029714f
C1497 VTAIL.n629 VSUBS 0.029714f
C1498 VTAIL.n630 VSUBS 0.013311f
C1499 VTAIL.n631 VSUBS 0.012571f
C1500 VTAIL.n632 VSUBS 0.023395f
C1501 VTAIL.n633 VSUBS 0.023395f
C1502 VTAIL.n634 VSUBS 0.012571f
C1503 VTAIL.n635 VSUBS 0.013311f
C1504 VTAIL.n636 VSUBS 0.029714f
C1505 VTAIL.n637 VSUBS 0.029714f
C1506 VTAIL.n638 VSUBS 0.029714f
C1507 VTAIL.n639 VSUBS 0.012941f
C1508 VTAIL.n640 VSUBS 0.012571f
C1509 VTAIL.n641 VSUBS 0.023395f
C1510 VTAIL.n642 VSUBS 0.023395f
C1511 VTAIL.n643 VSUBS 0.012571f
C1512 VTAIL.n644 VSUBS 0.013311f
C1513 VTAIL.n645 VSUBS 0.029714f
C1514 VTAIL.n646 VSUBS 0.029714f
C1515 VTAIL.n647 VSUBS 0.013311f
C1516 VTAIL.n648 VSUBS 0.012571f
C1517 VTAIL.n649 VSUBS 0.023395f
C1518 VTAIL.n650 VSUBS 0.023395f
C1519 VTAIL.n651 VSUBS 0.012571f
C1520 VTAIL.n652 VSUBS 0.013311f
C1521 VTAIL.n653 VSUBS 0.029714f
C1522 VTAIL.n654 VSUBS 0.029714f
C1523 VTAIL.n655 VSUBS 0.013311f
C1524 VTAIL.n656 VSUBS 0.012571f
C1525 VTAIL.n657 VSUBS 0.023395f
C1526 VTAIL.n658 VSUBS 0.023395f
C1527 VTAIL.n659 VSUBS 0.012571f
C1528 VTAIL.n660 VSUBS 0.013311f
C1529 VTAIL.n661 VSUBS 0.029714f
C1530 VTAIL.n662 VSUBS 0.029714f
C1531 VTAIL.n663 VSUBS 0.013311f
C1532 VTAIL.n664 VSUBS 0.012571f
C1533 VTAIL.n665 VSUBS 0.023395f
C1534 VTAIL.n666 VSUBS 0.023395f
C1535 VTAIL.n667 VSUBS 0.012571f
C1536 VTAIL.n668 VSUBS 0.013311f
C1537 VTAIL.n669 VSUBS 0.029714f
C1538 VTAIL.n670 VSUBS 0.029714f
C1539 VTAIL.n671 VSUBS 0.013311f
C1540 VTAIL.n672 VSUBS 0.012571f
C1541 VTAIL.n673 VSUBS 0.023395f
C1542 VTAIL.n674 VSUBS 0.060787f
C1543 VTAIL.n675 VSUBS 0.012571f
C1544 VTAIL.n676 VSUBS 0.013311f
C1545 VTAIL.n677 VSUBS 0.065183f
C1546 VTAIL.n678 VSUBS 0.044276f
C1547 VTAIL.n679 VSUBS 1.65831f
C1548 VTAIL.n680 VSUBS 0.013195f
C1549 VTAIL.n681 VSUBS 0.029714f
C1550 VTAIL.n682 VSUBS 0.013311f
C1551 VTAIL.n683 VSUBS 0.023395f
C1552 VTAIL.n684 VSUBS 0.012571f
C1553 VTAIL.n685 VSUBS 0.029714f
C1554 VTAIL.n686 VSUBS 0.013311f
C1555 VTAIL.n687 VSUBS 0.023395f
C1556 VTAIL.n688 VSUBS 0.012571f
C1557 VTAIL.n689 VSUBS 0.029714f
C1558 VTAIL.n690 VSUBS 0.013311f
C1559 VTAIL.n691 VSUBS 0.023395f
C1560 VTAIL.n692 VSUBS 0.012571f
C1561 VTAIL.n693 VSUBS 0.029714f
C1562 VTAIL.n694 VSUBS 0.013311f
C1563 VTAIL.n695 VSUBS 0.023395f
C1564 VTAIL.n696 VSUBS 0.012571f
C1565 VTAIL.n697 VSUBS 0.029714f
C1566 VTAIL.n698 VSUBS 0.013311f
C1567 VTAIL.n699 VSUBS 0.023395f
C1568 VTAIL.n700 VSUBS 0.012941f
C1569 VTAIL.n701 VSUBS 0.029714f
C1570 VTAIL.n702 VSUBS 0.013311f
C1571 VTAIL.n703 VSUBS 0.023395f
C1572 VTAIL.n704 VSUBS 0.012571f
C1573 VTAIL.n705 VSUBS 0.029714f
C1574 VTAIL.n706 VSUBS 0.013311f
C1575 VTAIL.n707 VSUBS 0.023395f
C1576 VTAIL.n708 VSUBS 0.012571f
C1577 VTAIL.n709 VSUBS 0.022286f
C1578 VTAIL.n710 VSUBS 0.022352f
C1579 VTAIL.t14 VSUBS 0.064453f
C1580 VTAIL.n711 VSUBS 0.24105f
C1581 VTAIL.n712 VSUBS 1.69992f
C1582 VTAIL.n713 VSUBS 0.012571f
C1583 VTAIL.n714 VSUBS 0.013311f
C1584 VTAIL.n715 VSUBS 0.029714f
C1585 VTAIL.n716 VSUBS 0.029714f
C1586 VTAIL.n717 VSUBS 0.013311f
C1587 VTAIL.n718 VSUBS 0.012571f
C1588 VTAIL.n719 VSUBS 0.023395f
C1589 VTAIL.n720 VSUBS 0.023395f
C1590 VTAIL.n721 VSUBS 0.012571f
C1591 VTAIL.n722 VSUBS 0.013311f
C1592 VTAIL.n723 VSUBS 0.029714f
C1593 VTAIL.n724 VSUBS 0.029714f
C1594 VTAIL.n725 VSUBS 0.013311f
C1595 VTAIL.n726 VSUBS 0.012571f
C1596 VTAIL.n727 VSUBS 0.023395f
C1597 VTAIL.n728 VSUBS 0.023395f
C1598 VTAIL.n729 VSUBS 0.012571f
C1599 VTAIL.n730 VSUBS 0.012571f
C1600 VTAIL.n731 VSUBS 0.013311f
C1601 VTAIL.n732 VSUBS 0.029714f
C1602 VTAIL.n733 VSUBS 0.029714f
C1603 VTAIL.n734 VSUBS 0.029714f
C1604 VTAIL.n735 VSUBS 0.012941f
C1605 VTAIL.n736 VSUBS 0.012571f
C1606 VTAIL.n737 VSUBS 0.023395f
C1607 VTAIL.n738 VSUBS 0.023395f
C1608 VTAIL.n739 VSUBS 0.012571f
C1609 VTAIL.n740 VSUBS 0.013311f
C1610 VTAIL.n741 VSUBS 0.029714f
C1611 VTAIL.n742 VSUBS 0.029714f
C1612 VTAIL.n743 VSUBS 0.013311f
C1613 VTAIL.n744 VSUBS 0.012571f
C1614 VTAIL.n745 VSUBS 0.023395f
C1615 VTAIL.n746 VSUBS 0.023395f
C1616 VTAIL.n747 VSUBS 0.012571f
C1617 VTAIL.n748 VSUBS 0.013311f
C1618 VTAIL.n749 VSUBS 0.029714f
C1619 VTAIL.n750 VSUBS 0.029714f
C1620 VTAIL.n751 VSUBS 0.013311f
C1621 VTAIL.n752 VSUBS 0.012571f
C1622 VTAIL.n753 VSUBS 0.023395f
C1623 VTAIL.n754 VSUBS 0.023395f
C1624 VTAIL.n755 VSUBS 0.012571f
C1625 VTAIL.n756 VSUBS 0.013311f
C1626 VTAIL.n757 VSUBS 0.029714f
C1627 VTAIL.n758 VSUBS 0.029714f
C1628 VTAIL.n759 VSUBS 0.013311f
C1629 VTAIL.n760 VSUBS 0.012571f
C1630 VTAIL.n761 VSUBS 0.023395f
C1631 VTAIL.n762 VSUBS 0.023395f
C1632 VTAIL.n763 VSUBS 0.012571f
C1633 VTAIL.n764 VSUBS 0.013311f
C1634 VTAIL.n765 VSUBS 0.029714f
C1635 VTAIL.n766 VSUBS 0.029714f
C1636 VTAIL.n767 VSUBS 0.013311f
C1637 VTAIL.n768 VSUBS 0.012571f
C1638 VTAIL.n769 VSUBS 0.023395f
C1639 VTAIL.n770 VSUBS 0.060787f
C1640 VTAIL.n771 VSUBS 0.012571f
C1641 VTAIL.n772 VSUBS 0.013311f
C1642 VTAIL.n773 VSUBS 0.065183f
C1643 VTAIL.n774 VSUBS 0.044276f
C1644 VTAIL.n775 VSUBS 1.65392f
C1645 VN.n0 VSUBS 0.055344f
C1646 VN.t2 VSUBS 2.23769f
C1647 VN.n1 VSUBS 0.798653f
C1648 VN.n2 VSUBS 0.218354f
C1649 VN.t0 VSUBS 2.23769f
C1650 VN.t6 VSUBS 2.35685f
C1651 VN.n3 VSUBS 0.85406f
C1652 VN.n4 VSUBS 0.865971f
C1653 VN.n5 VSUBS 0.059021f
C1654 VN.n6 VSUBS 0.059021f
C1655 VN.n7 VSUBS 0.041476f
C1656 VN.n8 VSUBS 0.041476f
C1657 VN.n9 VSUBS 0.040663f
C1658 VN.n10 VSUBS 0.053922f
C1659 VN.t4 VSUBS 2.30949f
C1660 VN.n11 VSUBS 0.87209f
C1661 VN.n12 VSUBS 0.038844f
C1662 VN.n13 VSUBS 0.055344f
C1663 VN.t7 VSUBS 2.23769f
C1664 VN.n14 VSUBS 0.798653f
C1665 VN.n15 VSUBS 0.218354f
C1666 VN.t1 VSUBS 2.23769f
C1667 VN.t3 VSUBS 2.35685f
C1668 VN.n16 VSUBS 0.85406f
C1669 VN.n17 VSUBS 0.865971f
C1670 VN.n18 VSUBS 0.059021f
C1671 VN.n19 VSUBS 0.059021f
C1672 VN.n20 VSUBS 0.041476f
C1673 VN.n21 VSUBS 0.041476f
C1674 VN.n22 VSUBS 0.040663f
C1675 VN.n23 VSUBS 0.053922f
C1676 VN.t5 VSUBS 2.30949f
C1677 VN.n24 VSUBS 0.87209f
C1678 VN.n25 VSUBS 2.17639f
.ends

