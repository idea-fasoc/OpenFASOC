* NGSPICE file created from diff_pair_sample_0609.ext - technology: sky130A

.subckt diff_pair_sample_0609 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=1.4547 ps=8.24 w=3.73 l=2.96
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=1.4547 ps=8.24 w=3.73 l=2.96
X2 B.t11 B.t9 B.t10 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=0 ps=0 w=3.73 l=2.96
X3 B.t8 B.t6 B.t7 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=0 ps=0 w=3.73 l=2.96
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=1.4547 ps=8.24 w=3.73 l=2.96
X5 B.t5 B.t3 B.t4 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=0 ps=0 w=3.73 l=2.96
X6 B.t2 B.t0 B.t1 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=0 ps=0 w=3.73 l=2.96
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n2286_n1714# sky130_fd_pr__pfet_01v8 ad=1.4547 pd=8.24 as=1.4547 ps=8.24 w=3.73 l=2.96
R0 VN VN.t1 110.814
R1 VN VN.t0 71.8968
R2 VTAIL.n2 VTAIL.t1 110.761
R3 VTAIL.n1 VTAIL.t2 110.761
R4 VTAIL.n3 VTAIL.t3 110.761
R5 VTAIL.n0 VTAIL.t0 110.761
R6 VTAIL.n1 VTAIL.n0 21.2548
R7 VTAIL.n3 VTAIL.n2 18.4186
R8 VTAIL.n2 VTAIL.n1 1.88843
R9 VTAIL VTAIL.n0 1.23757
R10 VTAIL VTAIL.n3 0.651362
R11 VDD2.n0 VDD2.t1 159.988
R12 VDD2.n0 VDD2.t0 127.441
R13 VDD2 VDD2.n0 0.767741
R14 VP.n0 VP.t0 110.811
R15 VP.n0 VP.t1 71.4654
R16 VP VP.n0 0.431811
R17 VDD1 VDD1.t0 161.221
R18 VDD1 VDD1.t1 128.208
R19 B.n215 B.n70 585
R20 B.n214 B.n213 585
R21 B.n212 B.n71 585
R22 B.n211 B.n210 585
R23 B.n209 B.n72 585
R24 B.n208 B.n207 585
R25 B.n206 B.n73 585
R26 B.n205 B.n204 585
R27 B.n203 B.n74 585
R28 B.n202 B.n201 585
R29 B.n200 B.n75 585
R30 B.n199 B.n198 585
R31 B.n197 B.n76 585
R32 B.n196 B.n195 585
R33 B.n194 B.n77 585
R34 B.n193 B.n192 585
R35 B.n191 B.n78 585
R36 B.n190 B.n189 585
R37 B.n185 B.n79 585
R38 B.n184 B.n183 585
R39 B.n182 B.n80 585
R40 B.n181 B.n180 585
R41 B.n179 B.n81 585
R42 B.n178 B.n177 585
R43 B.n176 B.n82 585
R44 B.n175 B.n174 585
R45 B.n173 B.n83 585
R46 B.n171 B.n170 585
R47 B.n169 B.n86 585
R48 B.n168 B.n167 585
R49 B.n166 B.n87 585
R50 B.n165 B.n164 585
R51 B.n163 B.n88 585
R52 B.n162 B.n161 585
R53 B.n160 B.n89 585
R54 B.n159 B.n158 585
R55 B.n157 B.n90 585
R56 B.n156 B.n155 585
R57 B.n154 B.n91 585
R58 B.n153 B.n152 585
R59 B.n151 B.n92 585
R60 B.n150 B.n149 585
R61 B.n148 B.n93 585
R62 B.n147 B.n146 585
R63 B.n217 B.n216 585
R64 B.n218 B.n69 585
R65 B.n220 B.n219 585
R66 B.n221 B.n68 585
R67 B.n223 B.n222 585
R68 B.n224 B.n67 585
R69 B.n226 B.n225 585
R70 B.n227 B.n66 585
R71 B.n229 B.n228 585
R72 B.n230 B.n65 585
R73 B.n232 B.n231 585
R74 B.n233 B.n64 585
R75 B.n235 B.n234 585
R76 B.n236 B.n63 585
R77 B.n238 B.n237 585
R78 B.n239 B.n62 585
R79 B.n241 B.n240 585
R80 B.n242 B.n61 585
R81 B.n244 B.n243 585
R82 B.n245 B.n60 585
R83 B.n247 B.n246 585
R84 B.n248 B.n59 585
R85 B.n250 B.n249 585
R86 B.n251 B.n58 585
R87 B.n253 B.n252 585
R88 B.n254 B.n57 585
R89 B.n256 B.n255 585
R90 B.n257 B.n56 585
R91 B.n259 B.n258 585
R92 B.n260 B.n55 585
R93 B.n262 B.n261 585
R94 B.n263 B.n54 585
R95 B.n265 B.n264 585
R96 B.n266 B.n53 585
R97 B.n268 B.n267 585
R98 B.n269 B.n52 585
R99 B.n271 B.n270 585
R100 B.n272 B.n51 585
R101 B.n274 B.n273 585
R102 B.n275 B.n50 585
R103 B.n277 B.n276 585
R104 B.n278 B.n49 585
R105 B.n280 B.n279 585
R106 B.n281 B.n48 585
R107 B.n283 B.n282 585
R108 B.n284 B.n47 585
R109 B.n286 B.n285 585
R110 B.n287 B.n46 585
R111 B.n289 B.n288 585
R112 B.n290 B.n45 585
R113 B.n292 B.n291 585
R114 B.n293 B.n44 585
R115 B.n295 B.n294 585
R116 B.n296 B.n43 585
R117 B.n298 B.n297 585
R118 B.n299 B.n42 585
R119 B.n367 B.n366 585
R120 B.n365 B.n16 585
R121 B.n364 B.n363 585
R122 B.n362 B.n17 585
R123 B.n361 B.n360 585
R124 B.n359 B.n18 585
R125 B.n358 B.n357 585
R126 B.n356 B.n19 585
R127 B.n355 B.n354 585
R128 B.n353 B.n20 585
R129 B.n352 B.n351 585
R130 B.n350 B.n21 585
R131 B.n349 B.n348 585
R132 B.n347 B.n22 585
R133 B.n346 B.n345 585
R134 B.n344 B.n23 585
R135 B.n343 B.n342 585
R136 B.n341 B.n340 585
R137 B.n339 B.n27 585
R138 B.n338 B.n337 585
R139 B.n336 B.n28 585
R140 B.n335 B.n334 585
R141 B.n333 B.n29 585
R142 B.n332 B.n331 585
R143 B.n330 B.n30 585
R144 B.n329 B.n328 585
R145 B.n327 B.n31 585
R146 B.n325 B.n324 585
R147 B.n323 B.n34 585
R148 B.n322 B.n321 585
R149 B.n320 B.n35 585
R150 B.n319 B.n318 585
R151 B.n317 B.n36 585
R152 B.n316 B.n315 585
R153 B.n314 B.n37 585
R154 B.n313 B.n312 585
R155 B.n311 B.n38 585
R156 B.n310 B.n309 585
R157 B.n308 B.n39 585
R158 B.n307 B.n306 585
R159 B.n305 B.n40 585
R160 B.n304 B.n303 585
R161 B.n302 B.n41 585
R162 B.n301 B.n300 585
R163 B.n368 B.n15 585
R164 B.n370 B.n369 585
R165 B.n371 B.n14 585
R166 B.n373 B.n372 585
R167 B.n374 B.n13 585
R168 B.n376 B.n375 585
R169 B.n377 B.n12 585
R170 B.n379 B.n378 585
R171 B.n380 B.n11 585
R172 B.n382 B.n381 585
R173 B.n383 B.n10 585
R174 B.n385 B.n384 585
R175 B.n386 B.n9 585
R176 B.n388 B.n387 585
R177 B.n389 B.n8 585
R178 B.n391 B.n390 585
R179 B.n392 B.n7 585
R180 B.n394 B.n393 585
R181 B.n395 B.n6 585
R182 B.n397 B.n396 585
R183 B.n398 B.n5 585
R184 B.n400 B.n399 585
R185 B.n401 B.n4 585
R186 B.n403 B.n402 585
R187 B.n404 B.n3 585
R188 B.n406 B.n405 585
R189 B.n407 B.n0 585
R190 B.n2 B.n1 585
R191 B.n108 B.n107 585
R192 B.n109 B.n106 585
R193 B.n111 B.n110 585
R194 B.n112 B.n105 585
R195 B.n114 B.n113 585
R196 B.n115 B.n104 585
R197 B.n117 B.n116 585
R198 B.n118 B.n103 585
R199 B.n120 B.n119 585
R200 B.n121 B.n102 585
R201 B.n123 B.n122 585
R202 B.n124 B.n101 585
R203 B.n126 B.n125 585
R204 B.n127 B.n100 585
R205 B.n129 B.n128 585
R206 B.n130 B.n99 585
R207 B.n132 B.n131 585
R208 B.n133 B.n98 585
R209 B.n135 B.n134 585
R210 B.n136 B.n97 585
R211 B.n138 B.n137 585
R212 B.n139 B.n96 585
R213 B.n141 B.n140 585
R214 B.n142 B.n95 585
R215 B.n144 B.n143 585
R216 B.n145 B.n94 585
R217 B.n146 B.n145 506.916
R218 B.n216 B.n215 506.916
R219 B.n300 B.n299 506.916
R220 B.n366 B.n15 506.916
R221 B.n409 B.n408 256.663
R222 B.n84 B.t9 238.901
R223 B.n186 B.t6 238.901
R224 B.n32 B.t0 238.901
R225 B.n24 B.t3 238.901
R226 B.n408 B.n407 235.042
R227 B.n408 B.n2 235.042
R228 B.n186 B.t7 195.989
R229 B.n32 B.t2 195.989
R230 B.n84 B.t10 195.987
R231 B.n24 B.t5 195.987
R232 B.n146 B.n93 163.367
R233 B.n150 B.n93 163.367
R234 B.n151 B.n150 163.367
R235 B.n152 B.n151 163.367
R236 B.n152 B.n91 163.367
R237 B.n156 B.n91 163.367
R238 B.n157 B.n156 163.367
R239 B.n158 B.n157 163.367
R240 B.n158 B.n89 163.367
R241 B.n162 B.n89 163.367
R242 B.n163 B.n162 163.367
R243 B.n164 B.n163 163.367
R244 B.n164 B.n87 163.367
R245 B.n168 B.n87 163.367
R246 B.n169 B.n168 163.367
R247 B.n170 B.n169 163.367
R248 B.n170 B.n83 163.367
R249 B.n175 B.n83 163.367
R250 B.n176 B.n175 163.367
R251 B.n177 B.n176 163.367
R252 B.n177 B.n81 163.367
R253 B.n181 B.n81 163.367
R254 B.n182 B.n181 163.367
R255 B.n183 B.n182 163.367
R256 B.n183 B.n79 163.367
R257 B.n190 B.n79 163.367
R258 B.n191 B.n190 163.367
R259 B.n192 B.n191 163.367
R260 B.n192 B.n77 163.367
R261 B.n196 B.n77 163.367
R262 B.n197 B.n196 163.367
R263 B.n198 B.n197 163.367
R264 B.n198 B.n75 163.367
R265 B.n202 B.n75 163.367
R266 B.n203 B.n202 163.367
R267 B.n204 B.n203 163.367
R268 B.n204 B.n73 163.367
R269 B.n208 B.n73 163.367
R270 B.n209 B.n208 163.367
R271 B.n210 B.n209 163.367
R272 B.n210 B.n71 163.367
R273 B.n214 B.n71 163.367
R274 B.n215 B.n214 163.367
R275 B.n299 B.n298 163.367
R276 B.n298 B.n43 163.367
R277 B.n294 B.n43 163.367
R278 B.n294 B.n293 163.367
R279 B.n293 B.n292 163.367
R280 B.n292 B.n45 163.367
R281 B.n288 B.n45 163.367
R282 B.n288 B.n287 163.367
R283 B.n287 B.n286 163.367
R284 B.n286 B.n47 163.367
R285 B.n282 B.n47 163.367
R286 B.n282 B.n281 163.367
R287 B.n281 B.n280 163.367
R288 B.n280 B.n49 163.367
R289 B.n276 B.n49 163.367
R290 B.n276 B.n275 163.367
R291 B.n275 B.n274 163.367
R292 B.n274 B.n51 163.367
R293 B.n270 B.n51 163.367
R294 B.n270 B.n269 163.367
R295 B.n269 B.n268 163.367
R296 B.n268 B.n53 163.367
R297 B.n264 B.n53 163.367
R298 B.n264 B.n263 163.367
R299 B.n263 B.n262 163.367
R300 B.n262 B.n55 163.367
R301 B.n258 B.n55 163.367
R302 B.n258 B.n257 163.367
R303 B.n257 B.n256 163.367
R304 B.n256 B.n57 163.367
R305 B.n252 B.n57 163.367
R306 B.n252 B.n251 163.367
R307 B.n251 B.n250 163.367
R308 B.n250 B.n59 163.367
R309 B.n246 B.n59 163.367
R310 B.n246 B.n245 163.367
R311 B.n245 B.n244 163.367
R312 B.n244 B.n61 163.367
R313 B.n240 B.n61 163.367
R314 B.n240 B.n239 163.367
R315 B.n239 B.n238 163.367
R316 B.n238 B.n63 163.367
R317 B.n234 B.n63 163.367
R318 B.n234 B.n233 163.367
R319 B.n233 B.n232 163.367
R320 B.n232 B.n65 163.367
R321 B.n228 B.n65 163.367
R322 B.n228 B.n227 163.367
R323 B.n227 B.n226 163.367
R324 B.n226 B.n67 163.367
R325 B.n222 B.n67 163.367
R326 B.n222 B.n221 163.367
R327 B.n221 B.n220 163.367
R328 B.n220 B.n69 163.367
R329 B.n216 B.n69 163.367
R330 B.n366 B.n365 163.367
R331 B.n365 B.n364 163.367
R332 B.n364 B.n17 163.367
R333 B.n360 B.n17 163.367
R334 B.n360 B.n359 163.367
R335 B.n359 B.n358 163.367
R336 B.n358 B.n19 163.367
R337 B.n354 B.n19 163.367
R338 B.n354 B.n353 163.367
R339 B.n353 B.n352 163.367
R340 B.n352 B.n21 163.367
R341 B.n348 B.n21 163.367
R342 B.n348 B.n347 163.367
R343 B.n347 B.n346 163.367
R344 B.n346 B.n23 163.367
R345 B.n342 B.n23 163.367
R346 B.n342 B.n341 163.367
R347 B.n341 B.n27 163.367
R348 B.n337 B.n27 163.367
R349 B.n337 B.n336 163.367
R350 B.n336 B.n335 163.367
R351 B.n335 B.n29 163.367
R352 B.n331 B.n29 163.367
R353 B.n331 B.n330 163.367
R354 B.n330 B.n329 163.367
R355 B.n329 B.n31 163.367
R356 B.n324 B.n31 163.367
R357 B.n324 B.n323 163.367
R358 B.n323 B.n322 163.367
R359 B.n322 B.n35 163.367
R360 B.n318 B.n35 163.367
R361 B.n318 B.n317 163.367
R362 B.n317 B.n316 163.367
R363 B.n316 B.n37 163.367
R364 B.n312 B.n37 163.367
R365 B.n312 B.n311 163.367
R366 B.n311 B.n310 163.367
R367 B.n310 B.n39 163.367
R368 B.n306 B.n39 163.367
R369 B.n306 B.n305 163.367
R370 B.n305 B.n304 163.367
R371 B.n304 B.n41 163.367
R372 B.n300 B.n41 163.367
R373 B.n370 B.n15 163.367
R374 B.n371 B.n370 163.367
R375 B.n372 B.n371 163.367
R376 B.n372 B.n13 163.367
R377 B.n376 B.n13 163.367
R378 B.n377 B.n376 163.367
R379 B.n378 B.n377 163.367
R380 B.n378 B.n11 163.367
R381 B.n382 B.n11 163.367
R382 B.n383 B.n382 163.367
R383 B.n384 B.n383 163.367
R384 B.n384 B.n9 163.367
R385 B.n388 B.n9 163.367
R386 B.n389 B.n388 163.367
R387 B.n390 B.n389 163.367
R388 B.n390 B.n7 163.367
R389 B.n394 B.n7 163.367
R390 B.n395 B.n394 163.367
R391 B.n396 B.n395 163.367
R392 B.n396 B.n5 163.367
R393 B.n400 B.n5 163.367
R394 B.n401 B.n400 163.367
R395 B.n402 B.n401 163.367
R396 B.n402 B.n3 163.367
R397 B.n406 B.n3 163.367
R398 B.n407 B.n406 163.367
R399 B.n108 B.n2 163.367
R400 B.n109 B.n108 163.367
R401 B.n110 B.n109 163.367
R402 B.n110 B.n105 163.367
R403 B.n114 B.n105 163.367
R404 B.n115 B.n114 163.367
R405 B.n116 B.n115 163.367
R406 B.n116 B.n103 163.367
R407 B.n120 B.n103 163.367
R408 B.n121 B.n120 163.367
R409 B.n122 B.n121 163.367
R410 B.n122 B.n101 163.367
R411 B.n126 B.n101 163.367
R412 B.n127 B.n126 163.367
R413 B.n128 B.n127 163.367
R414 B.n128 B.n99 163.367
R415 B.n132 B.n99 163.367
R416 B.n133 B.n132 163.367
R417 B.n134 B.n133 163.367
R418 B.n134 B.n97 163.367
R419 B.n138 B.n97 163.367
R420 B.n139 B.n138 163.367
R421 B.n140 B.n139 163.367
R422 B.n140 B.n95 163.367
R423 B.n144 B.n95 163.367
R424 B.n145 B.n144 163.367
R425 B.n187 B.t8 132.184
R426 B.n33 B.t1 132.184
R427 B.n85 B.t11 132.18
R428 B.n25 B.t4 132.18
R429 B.n85 B.n84 63.8066
R430 B.n187 B.n186 63.8066
R431 B.n33 B.n32 63.8066
R432 B.n25 B.n24 63.8066
R433 B.n172 B.n85 59.5399
R434 B.n188 B.n187 59.5399
R435 B.n326 B.n33 59.5399
R436 B.n26 B.n25 59.5399
R437 B.n368 B.n367 32.9371
R438 B.n301 B.n42 32.9371
R439 B.n217 B.n70 32.9371
R440 B.n147 B.n94 32.9371
R441 B B.n409 18.0485
R442 B.n369 B.n368 10.6151
R443 B.n369 B.n14 10.6151
R444 B.n373 B.n14 10.6151
R445 B.n374 B.n373 10.6151
R446 B.n375 B.n374 10.6151
R447 B.n375 B.n12 10.6151
R448 B.n379 B.n12 10.6151
R449 B.n380 B.n379 10.6151
R450 B.n381 B.n380 10.6151
R451 B.n381 B.n10 10.6151
R452 B.n385 B.n10 10.6151
R453 B.n386 B.n385 10.6151
R454 B.n387 B.n386 10.6151
R455 B.n387 B.n8 10.6151
R456 B.n391 B.n8 10.6151
R457 B.n392 B.n391 10.6151
R458 B.n393 B.n392 10.6151
R459 B.n393 B.n6 10.6151
R460 B.n397 B.n6 10.6151
R461 B.n398 B.n397 10.6151
R462 B.n399 B.n398 10.6151
R463 B.n399 B.n4 10.6151
R464 B.n403 B.n4 10.6151
R465 B.n404 B.n403 10.6151
R466 B.n405 B.n404 10.6151
R467 B.n405 B.n0 10.6151
R468 B.n367 B.n16 10.6151
R469 B.n363 B.n16 10.6151
R470 B.n363 B.n362 10.6151
R471 B.n362 B.n361 10.6151
R472 B.n361 B.n18 10.6151
R473 B.n357 B.n18 10.6151
R474 B.n357 B.n356 10.6151
R475 B.n356 B.n355 10.6151
R476 B.n355 B.n20 10.6151
R477 B.n351 B.n20 10.6151
R478 B.n351 B.n350 10.6151
R479 B.n350 B.n349 10.6151
R480 B.n349 B.n22 10.6151
R481 B.n345 B.n22 10.6151
R482 B.n345 B.n344 10.6151
R483 B.n344 B.n343 10.6151
R484 B.n340 B.n339 10.6151
R485 B.n339 B.n338 10.6151
R486 B.n338 B.n28 10.6151
R487 B.n334 B.n28 10.6151
R488 B.n334 B.n333 10.6151
R489 B.n333 B.n332 10.6151
R490 B.n332 B.n30 10.6151
R491 B.n328 B.n30 10.6151
R492 B.n328 B.n327 10.6151
R493 B.n325 B.n34 10.6151
R494 B.n321 B.n34 10.6151
R495 B.n321 B.n320 10.6151
R496 B.n320 B.n319 10.6151
R497 B.n319 B.n36 10.6151
R498 B.n315 B.n36 10.6151
R499 B.n315 B.n314 10.6151
R500 B.n314 B.n313 10.6151
R501 B.n313 B.n38 10.6151
R502 B.n309 B.n38 10.6151
R503 B.n309 B.n308 10.6151
R504 B.n308 B.n307 10.6151
R505 B.n307 B.n40 10.6151
R506 B.n303 B.n40 10.6151
R507 B.n303 B.n302 10.6151
R508 B.n302 B.n301 10.6151
R509 B.n297 B.n42 10.6151
R510 B.n297 B.n296 10.6151
R511 B.n296 B.n295 10.6151
R512 B.n295 B.n44 10.6151
R513 B.n291 B.n44 10.6151
R514 B.n291 B.n290 10.6151
R515 B.n290 B.n289 10.6151
R516 B.n289 B.n46 10.6151
R517 B.n285 B.n46 10.6151
R518 B.n285 B.n284 10.6151
R519 B.n284 B.n283 10.6151
R520 B.n283 B.n48 10.6151
R521 B.n279 B.n48 10.6151
R522 B.n279 B.n278 10.6151
R523 B.n278 B.n277 10.6151
R524 B.n277 B.n50 10.6151
R525 B.n273 B.n50 10.6151
R526 B.n273 B.n272 10.6151
R527 B.n272 B.n271 10.6151
R528 B.n271 B.n52 10.6151
R529 B.n267 B.n52 10.6151
R530 B.n267 B.n266 10.6151
R531 B.n266 B.n265 10.6151
R532 B.n265 B.n54 10.6151
R533 B.n261 B.n54 10.6151
R534 B.n261 B.n260 10.6151
R535 B.n260 B.n259 10.6151
R536 B.n259 B.n56 10.6151
R537 B.n255 B.n56 10.6151
R538 B.n255 B.n254 10.6151
R539 B.n254 B.n253 10.6151
R540 B.n253 B.n58 10.6151
R541 B.n249 B.n58 10.6151
R542 B.n249 B.n248 10.6151
R543 B.n248 B.n247 10.6151
R544 B.n247 B.n60 10.6151
R545 B.n243 B.n60 10.6151
R546 B.n243 B.n242 10.6151
R547 B.n242 B.n241 10.6151
R548 B.n241 B.n62 10.6151
R549 B.n237 B.n62 10.6151
R550 B.n237 B.n236 10.6151
R551 B.n236 B.n235 10.6151
R552 B.n235 B.n64 10.6151
R553 B.n231 B.n64 10.6151
R554 B.n231 B.n230 10.6151
R555 B.n230 B.n229 10.6151
R556 B.n229 B.n66 10.6151
R557 B.n225 B.n66 10.6151
R558 B.n225 B.n224 10.6151
R559 B.n224 B.n223 10.6151
R560 B.n223 B.n68 10.6151
R561 B.n219 B.n68 10.6151
R562 B.n219 B.n218 10.6151
R563 B.n218 B.n217 10.6151
R564 B.n107 B.n1 10.6151
R565 B.n107 B.n106 10.6151
R566 B.n111 B.n106 10.6151
R567 B.n112 B.n111 10.6151
R568 B.n113 B.n112 10.6151
R569 B.n113 B.n104 10.6151
R570 B.n117 B.n104 10.6151
R571 B.n118 B.n117 10.6151
R572 B.n119 B.n118 10.6151
R573 B.n119 B.n102 10.6151
R574 B.n123 B.n102 10.6151
R575 B.n124 B.n123 10.6151
R576 B.n125 B.n124 10.6151
R577 B.n125 B.n100 10.6151
R578 B.n129 B.n100 10.6151
R579 B.n130 B.n129 10.6151
R580 B.n131 B.n130 10.6151
R581 B.n131 B.n98 10.6151
R582 B.n135 B.n98 10.6151
R583 B.n136 B.n135 10.6151
R584 B.n137 B.n136 10.6151
R585 B.n137 B.n96 10.6151
R586 B.n141 B.n96 10.6151
R587 B.n142 B.n141 10.6151
R588 B.n143 B.n142 10.6151
R589 B.n143 B.n94 10.6151
R590 B.n148 B.n147 10.6151
R591 B.n149 B.n148 10.6151
R592 B.n149 B.n92 10.6151
R593 B.n153 B.n92 10.6151
R594 B.n154 B.n153 10.6151
R595 B.n155 B.n154 10.6151
R596 B.n155 B.n90 10.6151
R597 B.n159 B.n90 10.6151
R598 B.n160 B.n159 10.6151
R599 B.n161 B.n160 10.6151
R600 B.n161 B.n88 10.6151
R601 B.n165 B.n88 10.6151
R602 B.n166 B.n165 10.6151
R603 B.n167 B.n166 10.6151
R604 B.n167 B.n86 10.6151
R605 B.n171 B.n86 10.6151
R606 B.n174 B.n173 10.6151
R607 B.n174 B.n82 10.6151
R608 B.n178 B.n82 10.6151
R609 B.n179 B.n178 10.6151
R610 B.n180 B.n179 10.6151
R611 B.n180 B.n80 10.6151
R612 B.n184 B.n80 10.6151
R613 B.n185 B.n184 10.6151
R614 B.n189 B.n185 10.6151
R615 B.n193 B.n78 10.6151
R616 B.n194 B.n193 10.6151
R617 B.n195 B.n194 10.6151
R618 B.n195 B.n76 10.6151
R619 B.n199 B.n76 10.6151
R620 B.n200 B.n199 10.6151
R621 B.n201 B.n200 10.6151
R622 B.n201 B.n74 10.6151
R623 B.n205 B.n74 10.6151
R624 B.n206 B.n205 10.6151
R625 B.n207 B.n206 10.6151
R626 B.n207 B.n72 10.6151
R627 B.n211 B.n72 10.6151
R628 B.n212 B.n211 10.6151
R629 B.n213 B.n212 10.6151
R630 B.n213 B.n70 10.6151
R631 B.n343 B.n26 9.36635
R632 B.n326 B.n325 9.36635
R633 B.n172 B.n171 9.36635
R634 B.n188 B.n78 9.36635
R635 B.n409 B.n0 8.11757
R636 B.n409 B.n1 8.11757
R637 B.n340 B.n26 1.24928
R638 B.n327 B.n326 1.24928
R639 B.n173 B.n172 1.24928
R640 B.n189 B.n188 1.24928
C0 VN B 1.00203f
C1 VTAIL w_n2286_n1714# 1.58632f
C2 VDD1 VP 1.25608f
C3 VDD2 B 1.12838f
C4 VTAIL VN 1.25611f
C5 VDD2 VTAIL 3.04285f
C6 VP w_n2286_n1714# 3.3185f
C7 VDD1 w_n2286_n1714# 1.24846f
C8 VN VP 4.09798f
C9 VTAIL B 1.85404f
C10 VDD1 VN 0.152707f
C11 VDD2 VP 0.352429f
C12 VDD2 VDD1 0.717413f
C13 VN w_n2286_n1714# 3.02777f
C14 VP B 1.48323f
C15 VDD1 B 1.09491f
C16 VDD2 w_n2286_n1714# 1.27839f
C17 VTAIL VP 1.27026f
C18 VDD1 VTAIL 2.98779f
C19 VDD2 VN 1.05787f
C20 B w_n2286_n1714# 6.89773f
C21 VDD2 VSUBS 0.621493f
C22 VDD1 VSUBS 2.873214f
C23 VTAIL VSUBS 0.437711f
C24 VN VSUBS 5.48041f
C25 VP VSUBS 1.35207f
C26 B VSUBS 3.295468f
C27 w_n2286_n1714# VSUBS 49.405f
C28 B.n0 VSUBS 0.006412f
C29 B.n1 VSUBS 0.006412f
C30 B.n2 VSUBS 0.009483f
C31 B.n3 VSUBS 0.007267f
C32 B.n4 VSUBS 0.007267f
C33 B.n5 VSUBS 0.007267f
C34 B.n6 VSUBS 0.007267f
C35 B.n7 VSUBS 0.007267f
C36 B.n8 VSUBS 0.007267f
C37 B.n9 VSUBS 0.007267f
C38 B.n10 VSUBS 0.007267f
C39 B.n11 VSUBS 0.007267f
C40 B.n12 VSUBS 0.007267f
C41 B.n13 VSUBS 0.007267f
C42 B.n14 VSUBS 0.007267f
C43 B.n15 VSUBS 0.016777f
C44 B.n16 VSUBS 0.007267f
C45 B.n17 VSUBS 0.007267f
C46 B.n18 VSUBS 0.007267f
C47 B.n19 VSUBS 0.007267f
C48 B.n20 VSUBS 0.007267f
C49 B.n21 VSUBS 0.007267f
C50 B.n22 VSUBS 0.007267f
C51 B.n23 VSUBS 0.007267f
C52 B.t4 VSUBS 0.099217f
C53 B.t5 VSUBS 0.119427f
C54 B.t3 VSUBS 0.555349f
C55 B.n24 VSUBS 0.096065f
C56 B.n25 VSUBS 0.072441f
C57 B.n26 VSUBS 0.016837f
C58 B.n27 VSUBS 0.007267f
C59 B.n28 VSUBS 0.007267f
C60 B.n29 VSUBS 0.007267f
C61 B.n30 VSUBS 0.007267f
C62 B.n31 VSUBS 0.007267f
C63 B.t1 VSUBS 0.099217f
C64 B.t2 VSUBS 0.119427f
C65 B.t0 VSUBS 0.555349f
C66 B.n32 VSUBS 0.096065f
C67 B.n33 VSUBS 0.072441f
C68 B.n34 VSUBS 0.007267f
C69 B.n35 VSUBS 0.007267f
C70 B.n36 VSUBS 0.007267f
C71 B.n37 VSUBS 0.007267f
C72 B.n38 VSUBS 0.007267f
C73 B.n39 VSUBS 0.007267f
C74 B.n40 VSUBS 0.007267f
C75 B.n41 VSUBS 0.007267f
C76 B.n42 VSUBS 0.016777f
C77 B.n43 VSUBS 0.007267f
C78 B.n44 VSUBS 0.007267f
C79 B.n45 VSUBS 0.007267f
C80 B.n46 VSUBS 0.007267f
C81 B.n47 VSUBS 0.007267f
C82 B.n48 VSUBS 0.007267f
C83 B.n49 VSUBS 0.007267f
C84 B.n50 VSUBS 0.007267f
C85 B.n51 VSUBS 0.007267f
C86 B.n52 VSUBS 0.007267f
C87 B.n53 VSUBS 0.007267f
C88 B.n54 VSUBS 0.007267f
C89 B.n55 VSUBS 0.007267f
C90 B.n56 VSUBS 0.007267f
C91 B.n57 VSUBS 0.007267f
C92 B.n58 VSUBS 0.007267f
C93 B.n59 VSUBS 0.007267f
C94 B.n60 VSUBS 0.007267f
C95 B.n61 VSUBS 0.007267f
C96 B.n62 VSUBS 0.007267f
C97 B.n63 VSUBS 0.007267f
C98 B.n64 VSUBS 0.007267f
C99 B.n65 VSUBS 0.007267f
C100 B.n66 VSUBS 0.007267f
C101 B.n67 VSUBS 0.007267f
C102 B.n68 VSUBS 0.007267f
C103 B.n69 VSUBS 0.007267f
C104 B.n70 VSUBS 0.016569f
C105 B.n71 VSUBS 0.007267f
C106 B.n72 VSUBS 0.007267f
C107 B.n73 VSUBS 0.007267f
C108 B.n74 VSUBS 0.007267f
C109 B.n75 VSUBS 0.007267f
C110 B.n76 VSUBS 0.007267f
C111 B.n77 VSUBS 0.007267f
C112 B.n78 VSUBS 0.00684f
C113 B.n79 VSUBS 0.007267f
C114 B.n80 VSUBS 0.007267f
C115 B.n81 VSUBS 0.007267f
C116 B.n82 VSUBS 0.007267f
C117 B.n83 VSUBS 0.007267f
C118 B.t11 VSUBS 0.099217f
C119 B.t10 VSUBS 0.119427f
C120 B.t9 VSUBS 0.555349f
C121 B.n84 VSUBS 0.096065f
C122 B.n85 VSUBS 0.072441f
C123 B.n86 VSUBS 0.007267f
C124 B.n87 VSUBS 0.007267f
C125 B.n88 VSUBS 0.007267f
C126 B.n89 VSUBS 0.007267f
C127 B.n90 VSUBS 0.007267f
C128 B.n91 VSUBS 0.007267f
C129 B.n92 VSUBS 0.007267f
C130 B.n93 VSUBS 0.007267f
C131 B.n94 VSUBS 0.016777f
C132 B.n95 VSUBS 0.007267f
C133 B.n96 VSUBS 0.007267f
C134 B.n97 VSUBS 0.007267f
C135 B.n98 VSUBS 0.007267f
C136 B.n99 VSUBS 0.007267f
C137 B.n100 VSUBS 0.007267f
C138 B.n101 VSUBS 0.007267f
C139 B.n102 VSUBS 0.007267f
C140 B.n103 VSUBS 0.007267f
C141 B.n104 VSUBS 0.007267f
C142 B.n105 VSUBS 0.007267f
C143 B.n106 VSUBS 0.007267f
C144 B.n107 VSUBS 0.007267f
C145 B.n108 VSUBS 0.007267f
C146 B.n109 VSUBS 0.007267f
C147 B.n110 VSUBS 0.007267f
C148 B.n111 VSUBS 0.007267f
C149 B.n112 VSUBS 0.007267f
C150 B.n113 VSUBS 0.007267f
C151 B.n114 VSUBS 0.007267f
C152 B.n115 VSUBS 0.007267f
C153 B.n116 VSUBS 0.007267f
C154 B.n117 VSUBS 0.007267f
C155 B.n118 VSUBS 0.007267f
C156 B.n119 VSUBS 0.007267f
C157 B.n120 VSUBS 0.007267f
C158 B.n121 VSUBS 0.007267f
C159 B.n122 VSUBS 0.007267f
C160 B.n123 VSUBS 0.007267f
C161 B.n124 VSUBS 0.007267f
C162 B.n125 VSUBS 0.007267f
C163 B.n126 VSUBS 0.007267f
C164 B.n127 VSUBS 0.007267f
C165 B.n128 VSUBS 0.007267f
C166 B.n129 VSUBS 0.007267f
C167 B.n130 VSUBS 0.007267f
C168 B.n131 VSUBS 0.007267f
C169 B.n132 VSUBS 0.007267f
C170 B.n133 VSUBS 0.007267f
C171 B.n134 VSUBS 0.007267f
C172 B.n135 VSUBS 0.007267f
C173 B.n136 VSUBS 0.007267f
C174 B.n137 VSUBS 0.007267f
C175 B.n138 VSUBS 0.007267f
C176 B.n139 VSUBS 0.007267f
C177 B.n140 VSUBS 0.007267f
C178 B.n141 VSUBS 0.007267f
C179 B.n142 VSUBS 0.007267f
C180 B.n143 VSUBS 0.007267f
C181 B.n144 VSUBS 0.007267f
C182 B.n145 VSUBS 0.016777f
C183 B.n146 VSUBS 0.017421f
C184 B.n147 VSUBS 0.017421f
C185 B.n148 VSUBS 0.007267f
C186 B.n149 VSUBS 0.007267f
C187 B.n150 VSUBS 0.007267f
C188 B.n151 VSUBS 0.007267f
C189 B.n152 VSUBS 0.007267f
C190 B.n153 VSUBS 0.007267f
C191 B.n154 VSUBS 0.007267f
C192 B.n155 VSUBS 0.007267f
C193 B.n156 VSUBS 0.007267f
C194 B.n157 VSUBS 0.007267f
C195 B.n158 VSUBS 0.007267f
C196 B.n159 VSUBS 0.007267f
C197 B.n160 VSUBS 0.007267f
C198 B.n161 VSUBS 0.007267f
C199 B.n162 VSUBS 0.007267f
C200 B.n163 VSUBS 0.007267f
C201 B.n164 VSUBS 0.007267f
C202 B.n165 VSUBS 0.007267f
C203 B.n166 VSUBS 0.007267f
C204 B.n167 VSUBS 0.007267f
C205 B.n168 VSUBS 0.007267f
C206 B.n169 VSUBS 0.007267f
C207 B.n170 VSUBS 0.007267f
C208 B.n171 VSUBS 0.00684f
C209 B.n172 VSUBS 0.016837f
C210 B.n173 VSUBS 0.004061f
C211 B.n174 VSUBS 0.007267f
C212 B.n175 VSUBS 0.007267f
C213 B.n176 VSUBS 0.007267f
C214 B.n177 VSUBS 0.007267f
C215 B.n178 VSUBS 0.007267f
C216 B.n179 VSUBS 0.007267f
C217 B.n180 VSUBS 0.007267f
C218 B.n181 VSUBS 0.007267f
C219 B.n182 VSUBS 0.007267f
C220 B.n183 VSUBS 0.007267f
C221 B.n184 VSUBS 0.007267f
C222 B.n185 VSUBS 0.007267f
C223 B.t8 VSUBS 0.099217f
C224 B.t7 VSUBS 0.119427f
C225 B.t6 VSUBS 0.555349f
C226 B.n186 VSUBS 0.096065f
C227 B.n187 VSUBS 0.072441f
C228 B.n188 VSUBS 0.016837f
C229 B.n189 VSUBS 0.004061f
C230 B.n190 VSUBS 0.007267f
C231 B.n191 VSUBS 0.007267f
C232 B.n192 VSUBS 0.007267f
C233 B.n193 VSUBS 0.007267f
C234 B.n194 VSUBS 0.007267f
C235 B.n195 VSUBS 0.007267f
C236 B.n196 VSUBS 0.007267f
C237 B.n197 VSUBS 0.007267f
C238 B.n198 VSUBS 0.007267f
C239 B.n199 VSUBS 0.007267f
C240 B.n200 VSUBS 0.007267f
C241 B.n201 VSUBS 0.007267f
C242 B.n202 VSUBS 0.007267f
C243 B.n203 VSUBS 0.007267f
C244 B.n204 VSUBS 0.007267f
C245 B.n205 VSUBS 0.007267f
C246 B.n206 VSUBS 0.007267f
C247 B.n207 VSUBS 0.007267f
C248 B.n208 VSUBS 0.007267f
C249 B.n209 VSUBS 0.007267f
C250 B.n210 VSUBS 0.007267f
C251 B.n211 VSUBS 0.007267f
C252 B.n212 VSUBS 0.007267f
C253 B.n213 VSUBS 0.007267f
C254 B.n214 VSUBS 0.007267f
C255 B.n215 VSUBS 0.017421f
C256 B.n216 VSUBS 0.016777f
C257 B.n217 VSUBS 0.017629f
C258 B.n218 VSUBS 0.007267f
C259 B.n219 VSUBS 0.007267f
C260 B.n220 VSUBS 0.007267f
C261 B.n221 VSUBS 0.007267f
C262 B.n222 VSUBS 0.007267f
C263 B.n223 VSUBS 0.007267f
C264 B.n224 VSUBS 0.007267f
C265 B.n225 VSUBS 0.007267f
C266 B.n226 VSUBS 0.007267f
C267 B.n227 VSUBS 0.007267f
C268 B.n228 VSUBS 0.007267f
C269 B.n229 VSUBS 0.007267f
C270 B.n230 VSUBS 0.007267f
C271 B.n231 VSUBS 0.007267f
C272 B.n232 VSUBS 0.007267f
C273 B.n233 VSUBS 0.007267f
C274 B.n234 VSUBS 0.007267f
C275 B.n235 VSUBS 0.007267f
C276 B.n236 VSUBS 0.007267f
C277 B.n237 VSUBS 0.007267f
C278 B.n238 VSUBS 0.007267f
C279 B.n239 VSUBS 0.007267f
C280 B.n240 VSUBS 0.007267f
C281 B.n241 VSUBS 0.007267f
C282 B.n242 VSUBS 0.007267f
C283 B.n243 VSUBS 0.007267f
C284 B.n244 VSUBS 0.007267f
C285 B.n245 VSUBS 0.007267f
C286 B.n246 VSUBS 0.007267f
C287 B.n247 VSUBS 0.007267f
C288 B.n248 VSUBS 0.007267f
C289 B.n249 VSUBS 0.007267f
C290 B.n250 VSUBS 0.007267f
C291 B.n251 VSUBS 0.007267f
C292 B.n252 VSUBS 0.007267f
C293 B.n253 VSUBS 0.007267f
C294 B.n254 VSUBS 0.007267f
C295 B.n255 VSUBS 0.007267f
C296 B.n256 VSUBS 0.007267f
C297 B.n257 VSUBS 0.007267f
C298 B.n258 VSUBS 0.007267f
C299 B.n259 VSUBS 0.007267f
C300 B.n260 VSUBS 0.007267f
C301 B.n261 VSUBS 0.007267f
C302 B.n262 VSUBS 0.007267f
C303 B.n263 VSUBS 0.007267f
C304 B.n264 VSUBS 0.007267f
C305 B.n265 VSUBS 0.007267f
C306 B.n266 VSUBS 0.007267f
C307 B.n267 VSUBS 0.007267f
C308 B.n268 VSUBS 0.007267f
C309 B.n269 VSUBS 0.007267f
C310 B.n270 VSUBS 0.007267f
C311 B.n271 VSUBS 0.007267f
C312 B.n272 VSUBS 0.007267f
C313 B.n273 VSUBS 0.007267f
C314 B.n274 VSUBS 0.007267f
C315 B.n275 VSUBS 0.007267f
C316 B.n276 VSUBS 0.007267f
C317 B.n277 VSUBS 0.007267f
C318 B.n278 VSUBS 0.007267f
C319 B.n279 VSUBS 0.007267f
C320 B.n280 VSUBS 0.007267f
C321 B.n281 VSUBS 0.007267f
C322 B.n282 VSUBS 0.007267f
C323 B.n283 VSUBS 0.007267f
C324 B.n284 VSUBS 0.007267f
C325 B.n285 VSUBS 0.007267f
C326 B.n286 VSUBS 0.007267f
C327 B.n287 VSUBS 0.007267f
C328 B.n288 VSUBS 0.007267f
C329 B.n289 VSUBS 0.007267f
C330 B.n290 VSUBS 0.007267f
C331 B.n291 VSUBS 0.007267f
C332 B.n292 VSUBS 0.007267f
C333 B.n293 VSUBS 0.007267f
C334 B.n294 VSUBS 0.007267f
C335 B.n295 VSUBS 0.007267f
C336 B.n296 VSUBS 0.007267f
C337 B.n297 VSUBS 0.007267f
C338 B.n298 VSUBS 0.007267f
C339 B.n299 VSUBS 0.016777f
C340 B.n300 VSUBS 0.017421f
C341 B.n301 VSUBS 0.017421f
C342 B.n302 VSUBS 0.007267f
C343 B.n303 VSUBS 0.007267f
C344 B.n304 VSUBS 0.007267f
C345 B.n305 VSUBS 0.007267f
C346 B.n306 VSUBS 0.007267f
C347 B.n307 VSUBS 0.007267f
C348 B.n308 VSUBS 0.007267f
C349 B.n309 VSUBS 0.007267f
C350 B.n310 VSUBS 0.007267f
C351 B.n311 VSUBS 0.007267f
C352 B.n312 VSUBS 0.007267f
C353 B.n313 VSUBS 0.007267f
C354 B.n314 VSUBS 0.007267f
C355 B.n315 VSUBS 0.007267f
C356 B.n316 VSUBS 0.007267f
C357 B.n317 VSUBS 0.007267f
C358 B.n318 VSUBS 0.007267f
C359 B.n319 VSUBS 0.007267f
C360 B.n320 VSUBS 0.007267f
C361 B.n321 VSUBS 0.007267f
C362 B.n322 VSUBS 0.007267f
C363 B.n323 VSUBS 0.007267f
C364 B.n324 VSUBS 0.007267f
C365 B.n325 VSUBS 0.00684f
C366 B.n326 VSUBS 0.016837f
C367 B.n327 VSUBS 0.004061f
C368 B.n328 VSUBS 0.007267f
C369 B.n329 VSUBS 0.007267f
C370 B.n330 VSUBS 0.007267f
C371 B.n331 VSUBS 0.007267f
C372 B.n332 VSUBS 0.007267f
C373 B.n333 VSUBS 0.007267f
C374 B.n334 VSUBS 0.007267f
C375 B.n335 VSUBS 0.007267f
C376 B.n336 VSUBS 0.007267f
C377 B.n337 VSUBS 0.007267f
C378 B.n338 VSUBS 0.007267f
C379 B.n339 VSUBS 0.007267f
C380 B.n340 VSUBS 0.004061f
C381 B.n341 VSUBS 0.007267f
C382 B.n342 VSUBS 0.007267f
C383 B.n343 VSUBS 0.00684f
C384 B.n344 VSUBS 0.007267f
C385 B.n345 VSUBS 0.007267f
C386 B.n346 VSUBS 0.007267f
C387 B.n347 VSUBS 0.007267f
C388 B.n348 VSUBS 0.007267f
C389 B.n349 VSUBS 0.007267f
C390 B.n350 VSUBS 0.007267f
C391 B.n351 VSUBS 0.007267f
C392 B.n352 VSUBS 0.007267f
C393 B.n353 VSUBS 0.007267f
C394 B.n354 VSUBS 0.007267f
C395 B.n355 VSUBS 0.007267f
C396 B.n356 VSUBS 0.007267f
C397 B.n357 VSUBS 0.007267f
C398 B.n358 VSUBS 0.007267f
C399 B.n359 VSUBS 0.007267f
C400 B.n360 VSUBS 0.007267f
C401 B.n361 VSUBS 0.007267f
C402 B.n362 VSUBS 0.007267f
C403 B.n363 VSUBS 0.007267f
C404 B.n364 VSUBS 0.007267f
C405 B.n365 VSUBS 0.007267f
C406 B.n366 VSUBS 0.017421f
C407 B.n367 VSUBS 0.017421f
C408 B.n368 VSUBS 0.016777f
C409 B.n369 VSUBS 0.007267f
C410 B.n370 VSUBS 0.007267f
C411 B.n371 VSUBS 0.007267f
C412 B.n372 VSUBS 0.007267f
C413 B.n373 VSUBS 0.007267f
C414 B.n374 VSUBS 0.007267f
C415 B.n375 VSUBS 0.007267f
C416 B.n376 VSUBS 0.007267f
C417 B.n377 VSUBS 0.007267f
C418 B.n378 VSUBS 0.007267f
C419 B.n379 VSUBS 0.007267f
C420 B.n380 VSUBS 0.007267f
C421 B.n381 VSUBS 0.007267f
C422 B.n382 VSUBS 0.007267f
C423 B.n383 VSUBS 0.007267f
C424 B.n384 VSUBS 0.007267f
C425 B.n385 VSUBS 0.007267f
C426 B.n386 VSUBS 0.007267f
C427 B.n387 VSUBS 0.007267f
C428 B.n388 VSUBS 0.007267f
C429 B.n389 VSUBS 0.007267f
C430 B.n390 VSUBS 0.007267f
C431 B.n391 VSUBS 0.007267f
C432 B.n392 VSUBS 0.007267f
C433 B.n393 VSUBS 0.007267f
C434 B.n394 VSUBS 0.007267f
C435 B.n395 VSUBS 0.007267f
C436 B.n396 VSUBS 0.007267f
C437 B.n397 VSUBS 0.007267f
C438 B.n398 VSUBS 0.007267f
C439 B.n399 VSUBS 0.007267f
C440 B.n400 VSUBS 0.007267f
C441 B.n401 VSUBS 0.007267f
C442 B.n402 VSUBS 0.007267f
C443 B.n403 VSUBS 0.007267f
C444 B.n404 VSUBS 0.007267f
C445 B.n405 VSUBS 0.007267f
C446 B.n406 VSUBS 0.007267f
C447 B.n407 VSUBS 0.009483f
C448 B.n408 VSUBS 0.010102f
C449 B.n409 VSUBS 0.020089f
C450 VDD1.t1 VSUBS 0.357696f
C451 VDD1.t0 VSUBS 0.55491f
C452 VP.t1 VSUBS 1.60273f
C453 VP.t0 VSUBS 2.34075f
C454 VP.n0 VSUBS 3.33557f
C455 VDD2.t1 VSUBS 0.549057f
C456 VDD2.t0 VSUBS 0.362926f
C457 VDD2.n0 VSUBS 1.97543f
C458 VTAIL.t0 VSUBS 0.378335f
C459 VTAIL.n0 VSUBS 1.16744f
C460 VTAIL.t2 VSUBS 0.378337f
C461 VTAIL.n1 VSUBS 1.20628f
C462 VTAIL.t1 VSUBS 0.378337f
C463 VTAIL.n2 VSUBS 1.03705f
C464 VTAIL.t3 VSUBS 0.378335f
C465 VTAIL.n3 VSUBS 0.963243f
C466 VN.t0 VSUBS 1.52892f
C467 VN.t1 VSUBS 2.23236f
.ends

