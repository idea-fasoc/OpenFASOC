* NGSPICE file created from diff_pair_sample_0185.ext - technology: sky130A

.subckt diff_pair_sample_0185 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=2.63835 ps=16.32 w=15.99 l=2.33
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=0 ps=0 w=15.99 l=2.33
X2 VDD1.t3 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.63835 pd=16.32 as=6.2361 ps=32.76 w=15.99 l=2.33
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=0 ps=0 w=15.99 l=2.33
X4 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.63835 pd=16.32 as=6.2361 ps=32.76 w=15.99 l=2.33
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=0 ps=0 w=15.99 l=2.33
X6 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=2.63835 ps=16.32 w=15.99 l=2.33
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=0 ps=0 w=15.99 l=2.33
X8 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=2.63835 ps=16.32 w=15.99 l=2.33
X9 VDD1.t0 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.63835 pd=16.32 as=6.2361 ps=32.76 w=15.99 l=2.33
X10 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.63835 pd=16.32 as=6.2361 ps=32.76 w=15.99 l=2.33
X11 VTAIL.t4 VP.t3 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2361 pd=32.76 as=2.63835 ps=16.32 w=15.99 l=2.33
R0 VP.n3 VP.t0 201.917
R1 VP.n3 VP.t1 201.258
R2 VP.n5 VP.t3 165.391
R3 VP.n13 VP.t2 165.391
R4 VP.n12 VP.n0 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n1 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n6 VP.n2 161.3
R9 VP.n5 VP.n4 94.6082
R10 VP.n14 VP.n13 94.6082
R11 VP.n4 VP.n3 54.0078
R12 VP.n7 VP.n1 40.4934
R13 VP.n11 VP.n1 40.4934
R14 VP.n7 VP.n6 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 16.1487
R17 VP.n13 VP.n12 16.1487
R18 VP.n4 VP.n2 0.278367
R19 VP.n14 VP.n0 0.278367
R20 VP.n8 VP.n2 0.189894
R21 VP.n9 VP.n8 0.189894
R22 VP.n10 VP.n9 0.189894
R23 VP.n10 VP.n0 0.189894
R24 VP VP.n14 0.153454
R25 VDD1 VDD1.n1 103.936
R26 VDD1 VDD1.n0 59.0903
R27 VDD1.n0 VDD1.t2 1.23877
R28 VDD1.n0 VDD1.t3 1.23877
R29 VDD1.n1 VDD1.t1 1.23877
R30 VDD1.n1 VDD1.t0 1.23877
R31 VTAIL.n714 VTAIL.n630 289.615
R32 VTAIL.n84 VTAIL.n0 289.615
R33 VTAIL.n174 VTAIL.n90 289.615
R34 VTAIL.n264 VTAIL.n180 289.615
R35 VTAIL.n624 VTAIL.n540 289.615
R36 VTAIL.n534 VTAIL.n450 289.615
R37 VTAIL.n444 VTAIL.n360 289.615
R38 VTAIL.n354 VTAIL.n270 289.615
R39 VTAIL.n658 VTAIL.n657 185
R40 VTAIL.n663 VTAIL.n662 185
R41 VTAIL.n665 VTAIL.n664 185
R42 VTAIL.n654 VTAIL.n653 185
R43 VTAIL.n671 VTAIL.n670 185
R44 VTAIL.n673 VTAIL.n672 185
R45 VTAIL.n650 VTAIL.n649 185
R46 VTAIL.n679 VTAIL.n678 185
R47 VTAIL.n681 VTAIL.n680 185
R48 VTAIL.n646 VTAIL.n645 185
R49 VTAIL.n687 VTAIL.n686 185
R50 VTAIL.n689 VTAIL.n688 185
R51 VTAIL.n642 VTAIL.n641 185
R52 VTAIL.n695 VTAIL.n694 185
R53 VTAIL.n697 VTAIL.n696 185
R54 VTAIL.n638 VTAIL.n637 185
R55 VTAIL.n704 VTAIL.n703 185
R56 VTAIL.n705 VTAIL.n636 185
R57 VTAIL.n707 VTAIL.n706 185
R58 VTAIL.n634 VTAIL.n633 185
R59 VTAIL.n713 VTAIL.n712 185
R60 VTAIL.n715 VTAIL.n714 185
R61 VTAIL.n28 VTAIL.n27 185
R62 VTAIL.n33 VTAIL.n32 185
R63 VTAIL.n35 VTAIL.n34 185
R64 VTAIL.n24 VTAIL.n23 185
R65 VTAIL.n41 VTAIL.n40 185
R66 VTAIL.n43 VTAIL.n42 185
R67 VTAIL.n20 VTAIL.n19 185
R68 VTAIL.n49 VTAIL.n48 185
R69 VTAIL.n51 VTAIL.n50 185
R70 VTAIL.n16 VTAIL.n15 185
R71 VTAIL.n57 VTAIL.n56 185
R72 VTAIL.n59 VTAIL.n58 185
R73 VTAIL.n12 VTAIL.n11 185
R74 VTAIL.n65 VTAIL.n64 185
R75 VTAIL.n67 VTAIL.n66 185
R76 VTAIL.n8 VTAIL.n7 185
R77 VTAIL.n74 VTAIL.n73 185
R78 VTAIL.n75 VTAIL.n6 185
R79 VTAIL.n77 VTAIL.n76 185
R80 VTAIL.n4 VTAIL.n3 185
R81 VTAIL.n83 VTAIL.n82 185
R82 VTAIL.n85 VTAIL.n84 185
R83 VTAIL.n118 VTAIL.n117 185
R84 VTAIL.n123 VTAIL.n122 185
R85 VTAIL.n125 VTAIL.n124 185
R86 VTAIL.n114 VTAIL.n113 185
R87 VTAIL.n131 VTAIL.n130 185
R88 VTAIL.n133 VTAIL.n132 185
R89 VTAIL.n110 VTAIL.n109 185
R90 VTAIL.n139 VTAIL.n138 185
R91 VTAIL.n141 VTAIL.n140 185
R92 VTAIL.n106 VTAIL.n105 185
R93 VTAIL.n147 VTAIL.n146 185
R94 VTAIL.n149 VTAIL.n148 185
R95 VTAIL.n102 VTAIL.n101 185
R96 VTAIL.n155 VTAIL.n154 185
R97 VTAIL.n157 VTAIL.n156 185
R98 VTAIL.n98 VTAIL.n97 185
R99 VTAIL.n164 VTAIL.n163 185
R100 VTAIL.n165 VTAIL.n96 185
R101 VTAIL.n167 VTAIL.n166 185
R102 VTAIL.n94 VTAIL.n93 185
R103 VTAIL.n173 VTAIL.n172 185
R104 VTAIL.n175 VTAIL.n174 185
R105 VTAIL.n208 VTAIL.n207 185
R106 VTAIL.n213 VTAIL.n212 185
R107 VTAIL.n215 VTAIL.n214 185
R108 VTAIL.n204 VTAIL.n203 185
R109 VTAIL.n221 VTAIL.n220 185
R110 VTAIL.n223 VTAIL.n222 185
R111 VTAIL.n200 VTAIL.n199 185
R112 VTAIL.n229 VTAIL.n228 185
R113 VTAIL.n231 VTAIL.n230 185
R114 VTAIL.n196 VTAIL.n195 185
R115 VTAIL.n237 VTAIL.n236 185
R116 VTAIL.n239 VTAIL.n238 185
R117 VTAIL.n192 VTAIL.n191 185
R118 VTAIL.n245 VTAIL.n244 185
R119 VTAIL.n247 VTAIL.n246 185
R120 VTAIL.n188 VTAIL.n187 185
R121 VTAIL.n254 VTAIL.n253 185
R122 VTAIL.n255 VTAIL.n186 185
R123 VTAIL.n257 VTAIL.n256 185
R124 VTAIL.n184 VTAIL.n183 185
R125 VTAIL.n263 VTAIL.n262 185
R126 VTAIL.n265 VTAIL.n264 185
R127 VTAIL.n625 VTAIL.n624 185
R128 VTAIL.n623 VTAIL.n622 185
R129 VTAIL.n544 VTAIL.n543 185
R130 VTAIL.n617 VTAIL.n616 185
R131 VTAIL.n615 VTAIL.n546 185
R132 VTAIL.n614 VTAIL.n613 185
R133 VTAIL.n549 VTAIL.n547 185
R134 VTAIL.n608 VTAIL.n607 185
R135 VTAIL.n606 VTAIL.n605 185
R136 VTAIL.n553 VTAIL.n552 185
R137 VTAIL.n600 VTAIL.n599 185
R138 VTAIL.n598 VTAIL.n597 185
R139 VTAIL.n557 VTAIL.n556 185
R140 VTAIL.n592 VTAIL.n591 185
R141 VTAIL.n590 VTAIL.n589 185
R142 VTAIL.n561 VTAIL.n560 185
R143 VTAIL.n584 VTAIL.n583 185
R144 VTAIL.n582 VTAIL.n581 185
R145 VTAIL.n565 VTAIL.n564 185
R146 VTAIL.n576 VTAIL.n575 185
R147 VTAIL.n574 VTAIL.n573 185
R148 VTAIL.n569 VTAIL.n568 185
R149 VTAIL.n535 VTAIL.n534 185
R150 VTAIL.n533 VTAIL.n532 185
R151 VTAIL.n454 VTAIL.n453 185
R152 VTAIL.n527 VTAIL.n526 185
R153 VTAIL.n525 VTAIL.n456 185
R154 VTAIL.n524 VTAIL.n523 185
R155 VTAIL.n459 VTAIL.n457 185
R156 VTAIL.n518 VTAIL.n517 185
R157 VTAIL.n516 VTAIL.n515 185
R158 VTAIL.n463 VTAIL.n462 185
R159 VTAIL.n510 VTAIL.n509 185
R160 VTAIL.n508 VTAIL.n507 185
R161 VTAIL.n467 VTAIL.n466 185
R162 VTAIL.n502 VTAIL.n501 185
R163 VTAIL.n500 VTAIL.n499 185
R164 VTAIL.n471 VTAIL.n470 185
R165 VTAIL.n494 VTAIL.n493 185
R166 VTAIL.n492 VTAIL.n491 185
R167 VTAIL.n475 VTAIL.n474 185
R168 VTAIL.n486 VTAIL.n485 185
R169 VTAIL.n484 VTAIL.n483 185
R170 VTAIL.n479 VTAIL.n478 185
R171 VTAIL.n445 VTAIL.n444 185
R172 VTAIL.n443 VTAIL.n442 185
R173 VTAIL.n364 VTAIL.n363 185
R174 VTAIL.n437 VTAIL.n436 185
R175 VTAIL.n435 VTAIL.n366 185
R176 VTAIL.n434 VTAIL.n433 185
R177 VTAIL.n369 VTAIL.n367 185
R178 VTAIL.n428 VTAIL.n427 185
R179 VTAIL.n426 VTAIL.n425 185
R180 VTAIL.n373 VTAIL.n372 185
R181 VTAIL.n420 VTAIL.n419 185
R182 VTAIL.n418 VTAIL.n417 185
R183 VTAIL.n377 VTAIL.n376 185
R184 VTAIL.n412 VTAIL.n411 185
R185 VTAIL.n410 VTAIL.n409 185
R186 VTAIL.n381 VTAIL.n380 185
R187 VTAIL.n404 VTAIL.n403 185
R188 VTAIL.n402 VTAIL.n401 185
R189 VTAIL.n385 VTAIL.n384 185
R190 VTAIL.n396 VTAIL.n395 185
R191 VTAIL.n394 VTAIL.n393 185
R192 VTAIL.n389 VTAIL.n388 185
R193 VTAIL.n355 VTAIL.n354 185
R194 VTAIL.n353 VTAIL.n352 185
R195 VTAIL.n274 VTAIL.n273 185
R196 VTAIL.n347 VTAIL.n346 185
R197 VTAIL.n345 VTAIL.n276 185
R198 VTAIL.n344 VTAIL.n343 185
R199 VTAIL.n279 VTAIL.n277 185
R200 VTAIL.n338 VTAIL.n337 185
R201 VTAIL.n336 VTAIL.n335 185
R202 VTAIL.n283 VTAIL.n282 185
R203 VTAIL.n330 VTAIL.n329 185
R204 VTAIL.n328 VTAIL.n327 185
R205 VTAIL.n287 VTAIL.n286 185
R206 VTAIL.n322 VTAIL.n321 185
R207 VTAIL.n320 VTAIL.n319 185
R208 VTAIL.n291 VTAIL.n290 185
R209 VTAIL.n314 VTAIL.n313 185
R210 VTAIL.n312 VTAIL.n311 185
R211 VTAIL.n295 VTAIL.n294 185
R212 VTAIL.n306 VTAIL.n305 185
R213 VTAIL.n304 VTAIL.n303 185
R214 VTAIL.n299 VTAIL.n298 185
R215 VTAIL.n659 VTAIL.t1 147.659
R216 VTAIL.n29 VTAIL.t0 147.659
R217 VTAIL.n119 VTAIL.t5 147.659
R218 VTAIL.n209 VTAIL.t4 147.659
R219 VTAIL.n570 VTAIL.t6 147.659
R220 VTAIL.n480 VTAIL.t7 147.659
R221 VTAIL.n390 VTAIL.t3 147.659
R222 VTAIL.n300 VTAIL.t2 147.659
R223 VTAIL.n663 VTAIL.n657 104.615
R224 VTAIL.n664 VTAIL.n663 104.615
R225 VTAIL.n664 VTAIL.n653 104.615
R226 VTAIL.n671 VTAIL.n653 104.615
R227 VTAIL.n672 VTAIL.n671 104.615
R228 VTAIL.n672 VTAIL.n649 104.615
R229 VTAIL.n679 VTAIL.n649 104.615
R230 VTAIL.n680 VTAIL.n679 104.615
R231 VTAIL.n680 VTAIL.n645 104.615
R232 VTAIL.n687 VTAIL.n645 104.615
R233 VTAIL.n688 VTAIL.n687 104.615
R234 VTAIL.n688 VTAIL.n641 104.615
R235 VTAIL.n695 VTAIL.n641 104.615
R236 VTAIL.n696 VTAIL.n695 104.615
R237 VTAIL.n696 VTAIL.n637 104.615
R238 VTAIL.n704 VTAIL.n637 104.615
R239 VTAIL.n705 VTAIL.n704 104.615
R240 VTAIL.n706 VTAIL.n705 104.615
R241 VTAIL.n706 VTAIL.n633 104.615
R242 VTAIL.n713 VTAIL.n633 104.615
R243 VTAIL.n714 VTAIL.n713 104.615
R244 VTAIL.n33 VTAIL.n27 104.615
R245 VTAIL.n34 VTAIL.n33 104.615
R246 VTAIL.n34 VTAIL.n23 104.615
R247 VTAIL.n41 VTAIL.n23 104.615
R248 VTAIL.n42 VTAIL.n41 104.615
R249 VTAIL.n42 VTAIL.n19 104.615
R250 VTAIL.n49 VTAIL.n19 104.615
R251 VTAIL.n50 VTAIL.n49 104.615
R252 VTAIL.n50 VTAIL.n15 104.615
R253 VTAIL.n57 VTAIL.n15 104.615
R254 VTAIL.n58 VTAIL.n57 104.615
R255 VTAIL.n58 VTAIL.n11 104.615
R256 VTAIL.n65 VTAIL.n11 104.615
R257 VTAIL.n66 VTAIL.n65 104.615
R258 VTAIL.n66 VTAIL.n7 104.615
R259 VTAIL.n74 VTAIL.n7 104.615
R260 VTAIL.n75 VTAIL.n74 104.615
R261 VTAIL.n76 VTAIL.n75 104.615
R262 VTAIL.n76 VTAIL.n3 104.615
R263 VTAIL.n83 VTAIL.n3 104.615
R264 VTAIL.n84 VTAIL.n83 104.615
R265 VTAIL.n123 VTAIL.n117 104.615
R266 VTAIL.n124 VTAIL.n123 104.615
R267 VTAIL.n124 VTAIL.n113 104.615
R268 VTAIL.n131 VTAIL.n113 104.615
R269 VTAIL.n132 VTAIL.n131 104.615
R270 VTAIL.n132 VTAIL.n109 104.615
R271 VTAIL.n139 VTAIL.n109 104.615
R272 VTAIL.n140 VTAIL.n139 104.615
R273 VTAIL.n140 VTAIL.n105 104.615
R274 VTAIL.n147 VTAIL.n105 104.615
R275 VTAIL.n148 VTAIL.n147 104.615
R276 VTAIL.n148 VTAIL.n101 104.615
R277 VTAIL.n155 VTAIL.n101 104.615
R278 VTAIL.n156 VTAIL.n155 104.615
R279 VTAIL.n156 VTAIL.n97 104.615
R280 VTAIL.n164 VTAIL.n97 104.615
R281 VTAIL.n165 VTAIL.n164 104.615
R282 VTAIL.n166 VTAIL.n165 104.615
R283 VTAIL.n166 VTAIL.n93 104.615
R284 VTAIL.n173 VTAIL.n93 104.615
R285 VTAIL.n174 VTAIL.n173 104.615
R286 VTAIL.n213 VTAIL.n207 104.615
R287 VTAIL.n214 VTAIL.n213 104.615
R288 VTAIL.n214 VTAIL.n203 104.615
R289 VTAIL.n221 VTAIL.n203 104.615
R290 VTAIL.n222 VTAIL.n221 104.615
R291 VTAIL.n222 VTAIL.n199 104.615
R292 VTAIL.n229 VTAIL.n199 104.615
R293 VTAIL.n230 VTAIL.n229 104.615
R294 VTAIL.n230 VTAIL.n195 104.615
R295 VTAIL.n237 VTAIL.n195 104.615
R296 VTAIL.n238 VTAIL.n237 104.615
R297 VTAIL.n238 VTAIL.n191 104.615
R298 VTAIL.n245 VTAIL.n191 104.615
R299 VTAIL.n246 VTAIL.n245 104.615
R300 VTAIL.n246 VTAIL.n187 104.615
R301 VTAIL.n254 VTAIL.n187 104.615
R302 VTAIL.n255 VTAIL.n254 104.615
R303 VTAIL.n256 VTAIL.n255 104.615
R304 VTAIL.n256 VTAIL.n183 104.615
R305 VTAIL.n263 VTAIL.n183 104.615
R306 VTAIL.n264 VTAIL.n263 104.615
R307 VTAIL.n624 VTAIL.n623 104.615
R308 VTAIL.n623 VTAIL.n543 104.615
R309 VTAIL.n616 VTAIL.n543 104.615
R310 VTAIL.n616 VTAIL.n615 104.615
R311 VTAIL.n615 VTAIL.n614 104.615
R312 VTAIL.n614 VTAIL.n547 104.615
R313 VTAIL.n607 VTAIL.n547 104.615
R314 VTAIL.n607 VTAIL.n606 104.615
R315 VTAIL.n606 VTAIL.n552 104.615
R316 VTAIL.n599 VTAIL.n552 104.615
R317 VTAIL.n599 VTAIL.n598 104.615
R318 VTAIL.n598 VTAIL.n556 104.615
R319 VTAIL.n591 VTAIL.n556 104.615
R320 VTAIL.n591 VTAIL.n590 104.615
R321 VTAIL.n590 VTAIL.n560 104.615
R322 VTAIL.n583 VTAIL.n560 104.615
R323 VTAIL.n583 VTAIL.n582 104.615
R324 VTAIL.n582 VTAIL.n564 104.615
R325 VTAIL.n575 VTAIL.n564 104.615
R326 VTAIL.n575 VTAIL.n574 104.615
R327 VTAIL.n574 VTAIL.n568 104.615
R328 VTAIL.n534 VTAIL.n533 104.615
R329 VTAIL.n533 VTAIL.n453 104.615
R330 VTAIL.n526 VTAIL.n453 104.615
R331 VTAIL.n526 VTAIL.n525 104.615
R332 VTAIL.n525 VTAIL.n524 104.615
R333 VTAIL.n524 VTAIL.n457 104.615
R334 VTAIL.n517 VTAIL.n457 104.615
R335 VTAIL.n517 VTAIL.n516 104.615
R336 VTAIL.n516 VTAIL.n462 104.615
R337 VTAIL.n509 VTAIL.n462 104.615
R338 VTAIL.n509 VTAIL.n508 104.615
R339 VTAIL.n508 VTAIL.n466 104.615
R340 VTAIL.n501 VTAIL.n466 104.615
R341 VTAIL.n501 VTAIL.n500 104.615
R342 VTAIL.n500 VTAIL.n470 104.615
R343 VTAIL.n493 VTAIL.n470 104.615
R344 VTAIL.n493 VTAIL.n492 104.615
R345 VTAIL.n492 VTAIL.n474 104.615
R346 VTAIL.n485 VTAIL.n474 104.615
R347 VTAIL.n485 VTAIL.n484 104.615
R348 VTAIL.n484 VTAIL.n478 104.615
R349 VTAIL.n444 VTAIL.n443 104.615
R350 VTAIL.n443 VTAIL.n363 104.615
R351 VTAIL.n436 VTAIL.n363 104.615
R352 VTAIL.n436 VTAIL.n435 104.615
R353 VTAIL.n435 VTAIL.n434 104.615
R354 VTAIL.n434 VTAIL.n367 104.615
R355 VTAIL.n427 VTAIL.n367 104.615
R356 VTAIL.n427 VTAIL.n426 104.615
R357 VTAIL.n426 VTAIL.n372 104.615
R358 VTAIL.n419 VTAIL.n372 104.615
R359 VTAIL.n419 VTAIL.n418 104.615
R360 VTAIL.n418 VTAIL.n376 104.615
R361 VTAIL.n411 VTAIL.n376 104.615
R362 VTAIL.n411 VTAIL.n410 104.615
R363 VTAIL.n410 VTAIL.n380 104.615
R364 VTAIL.n403 VTAIL.n380 104.615
R365 VTAIL.n403 VTAIL.n402 104.615
R366 VTAIL.n402 VTAIL.n384 104.615
R367 VTAIL.n395 VTAIL.n384 104.615
R368 VTAIL.n395 VTAIL.n394 104.615
R369 VTAIL.n394 VTAIL.n388 104.615
R370 VTAIL.n354 VTAIL.n353 104.615
R371 VTAIL.n353 VTAIL.n273 104.615
R372 VTAIL.n346 VTAIL.n273 104.615
R373 VTAIL.n346 VTAIL.n345 104.615
R374 VTAIL.n345 VTAIL.n344 104.615
R375 VTAIL.n344 VTAIL.n277 104.615
R376 VTAIL.n337 VTAIL.n277 104.615
R377 VTAIL.n337 VTAIL.n336 104.615
R378 VTAIL.n336 VTAIL.n282 104.615
R379 VTAIL.n329 VTAIL.n282 104.615
R380 VTAIL.n329 VTAIL.n328 104.615
R381 VTAIL.n328 VTAIL.n286 104.615
R382 VTAIL.n321 VTAIL.n286 104.615
R383 VTAIL.n321 VTAIL.n320 104.615
R384 VTAIL.n320 VTAIL.n290 104.615
R385 VTAIL.n313 VTAIL.n290 104.615
R386 VTAIL.n313 VTAIL.n312 104.615
R387 VTAIL.n312 VTAIL.n294 104.615
R388 VTAIL.n305 VTAIL.n294 104.615
R389 VTAIL.n305 VTAIL.n304 104.615
R390 VTAIL.n304 VTAIL.n298 104.615
R391 VTAIL.t1 VTAIL.n657 52.3082
R392 VTAIL.t0 VTAIL.n27 52.3082
R393 VTAIL.t5 VTAIL.n117 52.3082
R394 VTAIL.t4 VTAIL.n207 52.3082
R395 VTAIL.t6 VTAIL.n568 52.3082
R396 VTAIL.t7 VTAIL.n478 52.3082
R397 VTAIL.t3 VTAIL.n388 52.3082
R398 VTAIL.t2 VTAIL.n298 52.3082
R399 VTAIL.n719 VTAIL.n718 30.4399
R400 VTAIL.n89 VTAIL.n88 30.4399
R401 VTAIL.n179 VTAIL.n178 30.4399
R402 VTAIL.n269 VTAIL.n268 30.4399
R403 VTAIL.n629 VTAIL.n628 30.4399
R404 VTAIL.n539 VTAIL.n538 30.4399
R405 VTAIL.n449 VTAIL.n448 30.4399
R406 VTAIL.n359 VTAIL.n358 30.4399
R407 VTAIL.n719 VTAIL.n629 28.4445
R408 VTAIL.n359 VTAIL.n269 28.4445
R409 VTAIL.n659 VTAIL.n658 15.6677
R410 VTAIL.n29 VTAIL.n28 15.6677
R411 VTAIL.n119 VTAIL.n118 15.6677
R412 VTAIL.n209 VTAIL.n208 15.6677
R413 VTAIL.n570 VTAIL.n569 15.6677
R414 VTAIL.n480 VTAIL.n479 15.6677
R415 VTAIL.n390 VTAIL.n389 15.6677
R416 VTAIL.n300 VTAIL.n299 15.6677
R417 VTAIL.n707 VTAIL.n636 13.1884
R418 VTAIL.n77 VTAIL.n6 13.1884
R419 VTAIL.n167 VTAIL.n96 13.1884
R420 VTAIL.n257 VTAIL.n186 13.1884
R421 VTAIL.n617 VTAIL.n546 13.1884
R422 VTAIL.n527 VTAIL.n456 13.1884
R423 VTAIL.n437 VTAIL.n366 13.1884
R424 VTAIL.n347 VTAIL.n276 13.1884
R425 VTAIL.n662 VTAIL.n661 12.8005
R426 VTAIL.n703 VTAIL.n702 12.8005
R427 VTAIL.n708 VTAIL.n634 12.8005
R428 VTAIL.n32 VTAIL.n31 12.8005
R429 VTAIL.n73 VTAIL.n72 12.8005
R430 VTAIL.n78 VTAIL.n4 12.8005
R431 VTAIL.n122 VTAIL.n121 12.8005
R432 VTAIL.n163 VTAIL.n162 12.8005
R433 VTAIL.n168 VTAIL.n94 12.8005
R434 VTAIL.n212 VTAIL.n211 12.8005
R435 VTAIL.n253 VTAIL.n252 12.8005
R436 VTAIL.n258 VTAIL.n184 12.8005
R437 VTAIL.n618 VTAIL.n544 12.8005
R438 VTAIL.n613 VTAIL.n548 12.8005
R439 VTAIL.n573 VTAIL.n572 12.8005
R440 VTAIL.n528 VTAIL.n454 12.8005
R441 VTAIL.n523 VTAIL.n458 12.8005
R442 VTAIL.n483 VTAIL.n482 12.8005
R443 VTAIL.n438 VTAIL.n364 12.8005
R444 VTAIL.n433 VTAIL.n368 12.8005
R445 VTAIL.n393 VTAIL.n392 12.8005
R446 VTAIL.n348 VTAIL.n274 12.8005
R447 VTAIL.n343 VTAIL.n278 12.8005
R448 VTAIL.n303 VTAIL.n302 12.8005
R449 VTAIL.n665 VTAIL.n656 12.0247
R450 VTAIL.n701 VTAIL.n638 12.0247
R451 VTAIL.n712 VTAIL.n711 12.0247
R452 VTAIL.n35 VTAIL.n26 12.0247
R453 VTAIL.n71 VTAIL.n8 12.0247
R454 VTAIL.n82 VTAIL.n81 12.0247
R455 VTAIL.n125 VTAIL.n116 12.0247
R456 VTAIL.n161 VTAIL.n98 12.0247
R457 VTAIL.n172 VTAIL.n171 12.0247
R458 VTAIL.n215 VTAIL.n206 12.0247
R459 VTAIL.n251 VTAIL.n188 12.0247
R460 VTAIL.n262 VTAIL.n261 12.0247
R461 VTAIL.n622 VTAIL.n621 12.0247
R462 VTAIL.n612 VTAIL.n549 12.0247
R463 VTAIL.n576 VTAIL.n567 12.0247
R464 VTAIL.n532 VTAIL.n531 12.0247
R465 VTAIL.n522 VTAIL.n459 12.0247
R466 VTAIL.n486 VTAIL.n477 12.0247
R467 VTAIL.n442 VTAIL.n441 12.0247
R468 VTAIL.n432 VTAIL.n369 12.0247
R469 VTAIL.n396 VTAIL.n387 12.0247
R470 VTAIL.n352 VTAIL.n351 12.0247
R471 VTAIL.n342 VTAIL.n279 12.0247
R472 VTAIL.n306 VTAIL.n297 12.0247
R473 VTAIL.n666 VTAIL.n654 11.249
R474 VTAIL.n698 VTAIL.n697 11.249
R475 VTAIL.n715 VTAIL.n632 11.249
R476 VTAIL.n36 VTAIL.n24 11.249
R477 VTAIL.n68 VTAIL.n67 11.249
R478 VTAIL.n85 VTAIL.n2 11.249
R479 VTAIL.n126 VTAIL.n114 11.249
R480 VTAIL.n158 VTAIL.n157 11.249
R481 VTAIL.n175 VTAIL.n92 11.249
R482 VTAIL.n216 VTAIL.n204 11.249
R483 VTAIL.n248 VTAIL.n247 11.249
R484 VTAIL.n265 VTAIL.n182 11.249
R485 VTAIL.n625 VTAIL.n542 11.249
R486 VTAIL.n609 VTAIL.n608 11.249
R487 VTAIL.n577 VTAIL.n565 11.249
R488 VTAIL.n535 VTAIL.n452 11.249
R489 VTAIL.n519 VTAIL.n518 11.249
R490 VTAIL.n487 VTAIL.n475 11.249
R491 VTAIL.n445 VTAIL.n362 11.249
R492 VTAIL.n429 VTAIL.n428 11.249
R493 VTAIL.n397 VTAIL.n385 11.249
R494 VTAIL.n355 VTAIL.n272 11.249
R495 VTAIL.n339 VTAIL.n338 11.249
R496 VTAIL.n307 VTAIL.n295 11.249
R497 VTAIL.n670 VTAIL.n669 10.4732
R498 VTAIL.n694 VTAIL.n640 10.4732
R499 VTAIL.n716 VTAIL.n630 10.4732
R500 VTAIL.n40 VTAIL.n39 10.4732
R501 VTAIL.n64 VTAIL.n10 10.4732
R502 VTAIL.n86 VTAIL.n0 10.4732
R503 VTAIL.n130 VTAIL.n129 10.4732
R504 VTAIL.n154 VTAIL.n100 10.4732
R505 VTAIL.n176 VTAIL.n90 10.4732
R506 VTAIL.n220 VTAIL.n219 10.4732
R507 VTAIL.n244 VTAIL.n190 10.4732
R508 VTAIL.n266 VTAIL.n180 10.4732
R509 VTAIL.n626 VTAIL.n540 10.4732
R510 VTAIL.n605 VTAIL.n551 10.4732
R511 VTAIL.n581 VTAIL.n580 10.4732
R512 VTAIL.n536 VTAIL.n450 10.4732
R513 VTAIL.n515 VTAIL.n461 10.4732
R514 VTAIL.n491 VTAIL.n490 10.4732
R515 VTAIL.n446 VTAIL.n360 10.4732
R516 VTAIL.n425 VTAIL.n371 10.4732
R517 VTAIL.n401 VTAIL.n400 10.4732
R518 VTAIL.n356 VTAIL.n270 10.4732
R519 VTAIL.n335 VTAIL.n281 10.4732
R520 VTAIL.n311 VTAIL.n310 10.4732
R521 VTAIL.n673 VTAIL.n652 9.69747
R522 VTAIL.n693 VTAIL.n642 9.69747
R523 VTAIL.n43 VTAIL.n22 9.69747
R524 VTAIL.n63 VTAIL.n12 9.69747
R525 VTAIL.n133 VTAIL.n112 9.69747
R526 VTAIL.n153 VTAIL.n102 9.69747
R527 VTAIL.n223 VTAIL.n202 9.69747
R528 VTAIL.n243 VTAIL.n192 9.69747
R529 VTAIL.n604 VTAIL.n553 9.69747
R530 VTAIL.n584 VTAIL.n563 9.69747
R531 VTAIL.n514 VTAIL.n463 9.69747
R532 VTAIL.n494 VTAIL.n473 9.69747
R533 VTAIL.n424 VTAIL.n373 9.69747
R534 VTAIL.n404 VTAIL.n383 9.69747
R535 VTAIL.n334 VTAIL.n283 9.69747
R536 VTAIL.n314 VTAIL.n293 9.69747
R537 VTAIL.n718 VTAIL.n717 9.45567
R538 VTAIL.n88 VTAIL.n87 9.45567
R539 VTAIL.n178 VTAIL.n177 9.45567
R540 VTAIL.n268 VTAIL.n267 9.45567
R541 VTAIL.n628 VTAIL.n627 9.45567
R542 VTAIL.n538 VTAIL.n537 9.45567
R543 VTAIL.n448 VTAIL.n447 9.45567
R544 VTAIL.n358 VTAIL.n357 9.45567
R545 VTAIL.n717 VTAIL.n716 9.3005
R546 VTAIL.n632 VTAIL.n631 9.3005
R547 VTAIL.n711 VTAIL.n710 9.3005
R548 VTAIL.n709 VTAIL.n708 9.3005
R549 VTAIL.n648 VTAIL.n647 9.3005
R550 VTAIL.n677 VTAIL.n676 9.3005
R551 VTAIL.n675 VTAIL.n674 9.3005
R552 VTAIL.n652 VTAIL.n651 9.3005
R553 VTAIL.n669 VTAIL.n668 9.3005
R554 VTAIL.n667 VTAIL.n666 9.3005
R555 VTAIL.n656 VTAIL.n655 9.3005
R556 VTAIL.n661 VTAIL.n660 9.3005
R557 VTAIL.n683 VTAIL.n682 9.3005
R558 VTAIL.n685 VTAIL.n684 9.3005
R559 VTAIL.n644 VTAIL.n643 9.3005
R560 VTAIL.n691 VTAIL.n690 9.3005
R561 VTAIL.n693 VTAIL.n692 9.3005
R562 VTAIL.n640 VTAIL.n639 9.3005
R563 VTAIL.n699 VTAIL.n698 9.3005
R564 VTAIL.n701 VTAIL.n700 9.3005
R565 VTAIL.n702 VTAIL.n635 9.3005
R566 VTAIL.n87 VTAIL.n86 9.3005
R567 VTAIL.n2 VTAIL.n1 9.3005
R568 VTAIL.n81 VTAIL.n80 9.3005
R569 VTAIL.n79 VTAIL.n78 9.3005
R570 VTAIL.n18 VTAIL.n17 9.3005
R571 VTAIL.n47 VTAIL.n46 9.3005
R572 VTAIL.n45 VTAIL.n44 9.3005
R573 VTAIL.n22 VTAIL.n21 9.3005
R574 VTAIL.n39 VTAIL.n38 9.3005
R575 VTAIL.n37 VTAIL.n36 9.3005
R576 VTAIL.n26 VTAIL.n25 9.3005
R577 VTAIL.n31 VTAIL.n30 9.3005
R578 VTAIL.n53 VTAIL.n52 9.3005
R579 VTAIL.n55 VTAIL.n54 9.3005
R580 VTAIL.n14 VTAIL.n13 9.3005
R581 VTAIL.n61 VTAIL.n60 9.3005
R582 VTAIL.n63 VTAIL.n62 9.3005
R583 VTAIL.n10 VTAIL.n9 9.3005
R584 VTAIL.n69 VTAIL.n68 9.3005
R585 VTAIL.n71 VTAIL.n70 9.3005
R586 VTAIL.n72 VTAIL.n5 9.3005
R587 VTAIL.n177 VTAIL.n176 9.3005
R588 VTAIL.n92 VTAIL.n91 9.3005
R589 VTAIL.n171 VTAIL.n170 9.3005
R590 VTAIL.n169 VTAIL.n168 9.3005
R591 VTAIL.n108 VTAIL.n107 9.3005
R592 VTAIL.n137 VTAIL.n136 9.3005
R593 VTAIL.n135 VTAIL.n134 9.3005
R594 VTAIL.n112 VTAIL.n111 9.3005
R595 VTAIL.n129 VTAIL.n128 9.3005
R596 VTAIL.n127 VTAIL.n126 9.3005
R597 VTAIL.n116 VTAIL.n115 9.3005
R598 VTAIL.n121 VTAIL.n120 9.3005
R599 VTAIL.n143 VTAIL.n142 9.3005
R600 VTAIL.n145 VTAIL.n144 9.3005
R601 VTAIL.n104 VTAIL.n103 9.3005
R602 VTAIL.n151 VTAIL.n150 9.3005
R603 VTAIL.n153 VTAIL.n152 9.3005
R604 VTAIL.n100 VTAIL.n99 9.3005
R605 VTAIL.n159 VTAIL.n158 9.3005
R606 VTAIL.n161 VTAIL.n160 9.3005
R607 VTAIL.n162 VTAIL.n95 9.3005
R608 VTAIL.n267 VTAIL.n266 9.3005
R609 VTAIL.n182 VTAIL.n181 9.3005
R610 VTAIL.n261 VTAIL.n260 9.3005
R611 VTAIL.n259 VTAIL.n258 9.3005
R612 VTAIL.n198 VTAIL.n197 9.3005
R613 VTAIL.n227 VTAIL.n226 9.3005
R614 VTAIL.n225 VTAIL.n224 9.3005
R615 VTAIL.n202 VTAIL.n201 9.3005
R616 VTAIL.n219 VTAIL.n218 9.3005
R617 VTAIL.n217 VTAIL.n216 9.3005
R618 VTAIL.n206 VTAIL.n205 9.3005
R619 VTAIL.n211 VTAIL.n210 9.3005
R620 VTAIL.n233 VTAIL.n232 9.3005
R621 VTAIL.n235 VTAIL.n234 9.3005
R622 VTAIL.n194 VTAIL.n193 9.3005
R623 VTAIL.n241 VTAIL.n240 9.3005
R624 VTAIL.n243 VTAIL.n242 9.3005
R625 VTAIL.n190 VTAIL.n189 9.3005
R626 VTAIL.n249 VTAIL.n248 9.3005
R627 VTAIL.n251 VTAIL.n250 9.3005
R628 VTAIL.n252 VTAIL.n185 9.3005
R629 VTAIL.n596 VTAIL.n595 9.3005
R630 VTAIL.n555 VTAIL.n554 9.3005
R631 VTAIL.n602 VTAIL.n601 9.3005
R632 VTAIL.n604 VTAIL.n603 9.3005
R633 VTAIL.n551 VTAIL.n550 9.3005
R634 VTAIL.n610 VTAIL.n609 9.3005
R635 VTAIL.n612 VTAIL.n611 9.3005
R636 VTAIL.n548 VTAIL.n545 9.3005
R637 VTAIL.n627 VTAIL.n626 9.3005
R638 VTAIL.n542 VTAIL.n541 9.3005
R639 VTAIL.n621 VTAIL.n620 9.3005
R640 VTAIL.n619 VTAIL.n618 9.3005
R641 VTAIL.n594 VTAIL.n593 9.3005
R642 VTAIL.n559 VTAIL.n558 9.3005
R643 VTAIL.n588 VTAIL.n587 9.3005
R644 VTAIL.n586 VTAIL.n585 9.3005
R645 VTAIL.n563 VTAIL.n562 9.3005
R646 VTAIL.n580 VTAIL.n579 9.3005
R647 VTAIL.n578 VTAIL.n577 9.3005
R648 VTAIL.n567 VTAIL.n566 9.3005
R649 VTAIL.n572 VTAIL.n571 9.3005
R650 VTAIL.n506 VTAIL.n505 9.3005
R651 VTAIL.n465 VTAIL.n464 9.3005
R652 VTAIL.n512 VTAIL.n511 9.3005
R653 VTAIL.n514 VTAIL.n513 9.3005
R654 VTAIL.n461 VTAIL.n460 9.3005
R655 VTAIL.n520 VTAIL.n519 9.3005
R656 VTAIL.n522 VTAIL.n521 9.3005
R657 VTAIL.n458 VTAIL.n455 9.3005
R658 VTAIL.n537 VTAIL.n536 9.3005
R659 VTAIL.n452 VTAIL.n451 9.3005
R660 VTAIL.n531 VTAIL.n530 9.3005
R661 VTAIL.n529 VTAIL.n528 9.3005
R662 VTAIL.n504 VTAIL.n503 9.3005
R663 VTAIL.n469 VTAIL.n468 9.3005
R664 VTAIL.n498 VTAIL.n497 9.3005
R665 VTAIL.n496 VTAIL.n495 9.3005
R666 VTAIL.n473 VTAIL.n472 9.3005
R667 VTAIL.n490 VTAIL.n489 9.3005
R668 VTAIL.n488 VTAIL.n487 9.3005
R669 VTAIL.n477 VTAIL.n476 9.3005
R670 VTAIL.n482 VTAIL.n481 9.3005
R671 VTAIL.n416 VTAIL.n415 9.3005
R672 VTAIL.n375 VTAIL.n374 9.3005
R673 VTAIL.n422 VTAIL.n421 9.3005
R674 VTAIL.n424 VTAIL.n423 9.3005
R675 VTAIL.n371 VTAIL.n370 9.3005
R676 VTAIL.n430 VTAIL.n429 9.3005
R677 VTAIL.n432 VTAIL.n431 9.3005
R678 VTAIL.n368 VTAIL.n365 9.3005
R679 VTAIL.n447 VTAIL.n446 9.3005
R680 VTAIL.n362 VTAIL.n361 9.3005
R681 VTAIL.n441 VTAIL.n440 9.3005
R682 VTAIL.n439 VTAIL.n438 9.3005
R683 VTAIL.n414 VTAIL.n413 9.3005
R684 VTAIL.n379 VTAIL.n378 9.3005
R685 VTAIL.n408 VTAIL.n407 9.3005
R686 VTAIL.n406 VTAIL.n405 9.3005
R687 VTAIL.n383 VTAIL.n382 9.3005
R688 VTAIL.n400 VTAIL.n399 9.3005
R689 VTAIL.n398 VTAIL.n397 9.3005
R690 VTAIL.n387 VTAIL.n386 9.3005
R691 VTAIL.n392 VTAIL.n391 9.3005
R692 VTAIL.n326 VTAIL.n325 9.3005
R693 VTAIL.n285 VTAIL.n284 9.3005
R694 VTAIL.n332 VTAIL.n331 9.3005
R695 VTAIL.n334 VTAIL.n333 9.3005
R696 VTAIL.n281 VTAIL.n280 9.3005
R697 VTAIL.n340 VTAIL.n339 9.3005
R698 VTAIL.n342 VTAIL.n341 9.3005
R699 VTAIL.n278 VTAIL.n275 9.3005
R700 VTAIL.n357 VTAIL.n356 9.3005
R701 VTAIL.n272 VTAIL.n271 9.3005
R702 VTAIL.n351 VTAIL.n350 9.3005
R703 VTAIL.n349 VTAIL.n348 9.3005
R704 VTAIL.n324 VTAIL.n323 9.3005
R705 VTAIL.n289 VTAIL.n288 9.3005
R706 VTAIL.n318 VTAIL.n317 9.3005
R707 VTAIL.n316 VTAIL.n315 9.3005
R708 VTAIL.n293 VTAIL.n292 9.3005
R709 VTAIL.n310 VTAIL.n309 9.3005
R710 VTAIL.n308 VTAIL.n307 9.3005
R711 VTAIL.n297 VTAIL.n296 9.3005
R712 VTAIL.n302 VTAIL.n301 9.3005
R713 VTAIL.n674 VTAIL.n650 8.92171
R714 VTAIL.n690 VTAIL.n689 8.92171
R715 VTAIL.n44 VTAIL.n20 8.92171
R716 VTAIL.n60 VTAIL.n59 8.92171
R717 VTAIL.n134 VTAIL.n110 8.92171
R718 VTAIL.n150 VTAIL.n149 8.92171
R719 VTAIL.n224 VTAIL.n200 8.92171
R720 VTAIL.n240 VTAIL.n239 8.92171
R721 VTAIL.n601 VTAIL.n600 8.92171
R722 VTAIL.n585 VTAIL.n561 8.92171
R723 VTAIL.n511 VTAIL.n510 8.92171
R724 VTAIL.n495 VTAIL.n471 8.92171
R725 VTAIL.n421 VTAIL.n420 8.92171
R726 VTAIL.n405 VTAIL.n381 8.92171
R727 VTAIL.n331 VTAIL.n330 8.92171
R728 VTAIL.n315 VTAIL.n291 8.92171
R729 VTAIL.n678 VTAIL.n677 8.14595
R730 VTAIL.n686 VTAIL.n644 8.14595
R731 VTAIL.n48 VTAIL.n47 8.14595
R732 VTAIL.n56 VTAIL.n14 8.14595
R733 VTAIL.n138 VTAIL.n137 8.14595
R734 VTAIL.n146 VTAIL.n104 8.14595
R735 VTAIL.n228 VTAIL.n227 8.14595
R736 VTAIL.n236 VTAIL.n194 8.14595
R737 VTAIL.n597 VTAIL.n555 8.14595
R738 VTAIL.n589 VTAIL.n588 8.14595
R739 VTAIL.n507 VTAIL.n465 8.14595
R740 VTAIL.n499 VTAIL.n498 8.14595
R741 VTAIL.n417 VTAIL.n375 8.14595
R742 VTAIL.n409 VTAIL.n408 8.14595
R743 VTAIL.n327 VTAIL.n285 8.14595
R744 VTAIL.n319 VTAIL.n318 8.14595
R745 VTAIL.n681 VTAIL.n648 7.3702
R746 VTAIL.n685 VTAIL.n646 7.3702
R747 VTAIL.n51 VTAIL.n18 7.3702
R748 VTAIL.n55 VTAIL.n16 7.3702
R749 VTAIL.n141 VTAIL.n108 7.3702
R750 VTAIL.n145 VTAIL.n106 7.3702
R751 VTAIL.n231 VTAIL.n198 7.3702
R752 VTAIL.n235 VTAIL.n196 7.3702
R753 VTAIL.n596 VTAIL.n557 7.3702
R754 VTAIL.n592 VTAIL.n559 7.3702
R755 VTAIL.n506 VTAIL.n467 7.3702
R756 VTAIL.n502 VTAIL.n469 7.3702
R757 VTAIL.n416 VTAIL.n377 7.3702
R758 VTAIL.n412 VTAIL.n379 7.3702
R759 VTAIL.n326 VTAIL.n287 7.3702
R760 VTAIL.n322 VTAIL.n289 7.3702
R761 VTAIL.n682 VTAIL.n681 6.59444
R762 VTAIL.n682 VTAIL.n646 6.59444
R763 VTAIL.n52 VTAIL.n51 6.59444
R764 VTAIL.n52 VTAIL.n16 6.59444
R765 VTAIL.n142 VTAIL.n141 6.59444
R766 VTAIL.n142 VTAIL.n106 6.59444
R767 VTAIL.n232 VTAIL.n231 6.59444
R768 VTAIL.n232 VTAIL.n196 6.59444
R769 VTAIL.n593 VTAIL.n557 6.59444
R770 VTAIL.n593 VTAIL.n592 6.59444
R771 VTAIL.n503 VTAIL.n467 6.59444
R772 VTAIL.n503 VTAIL.n502 6.59444
R773 VTAIL.n413 VTAIL.n377 6.59444
R774 VTAIL.n413 VTAIL.n412 6.59444
R775 VTAIL.n323 VTAIL.n287 6.59444
R776 VTAIL.n323 VTAIL.n322 6.59444
R777 VTAIL.n678 VTAIL.n648 5.81868
R778 VTAIL.n686 VTAIL.n685 5.81868
R779 VTAIL.n48 VTAIL.n18 5.81868
R780 VTAIL.n56 VTAIL.n55 5.81868
R781 VTAIL.n138 VTAIL.n108 5.81868
R782 VTAIL.n146 VTAIL.n145 5.81868
R783 VTAIL.n228 VTAIL.n198 5.81868
R784 VTAIL.n236 VTAIL.n235 5.81868
R785 VTAIL.n597 VTAIL.n596 5.81868
R786 VTAIL.n589 VTAIL.n559 5.81868
R787 VTAIL.n507 VTAIL.n506 5.81868
R788 VTAIL.n499 VTAIL.n469 5.81868
R789 VTAIL.n417 VTAIL.n416 5.81868
R790 VTAIL.n409 VTAIL.n379 5.81868
R791 VTAIL.n327 VTAIL.n326 5.81868
R792 VTAIL.n319 VTAIL.n289 5.81868
R793 VTAIL.n677 VTAIL.n650 5.04292
R794 VTAIL.n689 VTAIL.n644 5.04292
R795 VTAIL.n47 VTAIL.n20 5.04292
R796 VTAIL.n59 VTAIL.n14 5.04292
R797 VTAIL.n137 VTAIL.n110 5.04292
R798 VTAIL.n149 VTAIL.n104 5.04292
R799 VTAIL.n227 VTAIL.n200 5.04292
R800 VTAIL.n239 VTAIL.n194 5.04292
R801 VTAIL.n600 VTAIL.n555 5.04292
R802 VTAIL.n588 VTAIL.n561 5.04292
R803 VTAIL.n510 VTAIL.n465 5.04292
R804 VTAIL.n498 VTAIL.n471 5.04292
R805 VTAIL.n420 VTAIL.n375 5.04292
R806 VTAIL.n408 VTAIL.n381 5.04292
R807 VTAIL.n330 VTAIL.n285 5.04292
R808 VTAIL.n318 VTAIL.n291 5.04292
R809 VTAIL.n660 VTAIL.n659 4.38563
R810 VTAIL.n30 VTAIL.n29 4.38563
R811 VTAIL.n120 VTAIL.n119 4.38563
R812 VTAIL.n210 VTAIL.n209 4.38563
R813 VTAIL.n571 VTAIL.n570 4.38563
R814 VTAIL.n481 VTAIL.n480 4.38563
R815 VTAIL.n391 VTAIL.n390 4.38563
R816 VTAIL.n301 VTAIL.n300 4.38563
R817 VTAIL.n674 VTAIL.n673 4.26717
R818 VTAIL.n690 VTAIL.n642 4.26717
R819 VTAIL.n44 VTAIL.n43 4.26717
R820 VTAIL.n60 VTAIL.n12 4.26717
R821 VTAIL.n134 VTAIL.n133 4.26717
R822 VTAIL.n150 VTAIL.n102 4.26717
R823 VTAIL.n224 VTAIL.n223 4.26717
R824 VTAIL.n240 VTAIL.n192 4.26717
R825 VTAIL.n601 VTAIL.n553 4.26717
R826 VTAIL.n585 VTAIL.n584 4.26717
R827 VTAIL.n511 VTAIL.n463 4.26717
R828 VTAIL.n495 VTAIL.n494 4.26717
R829 VTAIL.n421 VTAIL.n373 4.26717
R830 VTAIL.n405 VTAIL.n404 4.26717
R831 VTAIL.n331 VTAIL.n283 4.26717
R832 VTAIL.n315 VTAIL.n314 4.26717
R833 VTAIL.n670 VTAIL.n652 3.49141
R834 VTAIL.n694 VTAIL.n693 3.49141
R835 VTAIL.n718 VTAIL.n630 3.49141
R836 VTAIL.n40 VTAIL.n22 3.49141
R837 VTAIL.n64 VTAIL.n63 3.49141
R838 VTAIL.n88 VTAIL.n0 3.49141
R839 VTAIL.n130 VTAIL.n112 3.49141
R840 VTAIL.n154 VTAIL.n153 3.49141
R841 VTAIL.n178 VTAIL.n90 3.49141
R842 VTAIL.n220 VTAIL.n202 3.49141
R843 VTAIL.n244 VTAIL.n243 3.49141
R844 VTAIL.n268 VTAIL.n180 3.49141
R845 VTAIL.n628 VTAIL.n540 3.49141
R846 VTAIL.n605 VTAIL.n604 3.49141
R847 VTAIL.n581 VTAIL.n563 3.49141
R848 VTAIL.n538 VTAIL.n450 3.49141
R849 VTAIL.n515 VTAIL.n514 3.49141
R850 VTAIL.n491 VTAIL.n473 3.49141
R851 VTAIL.n448 VTAIL.n360 3.49141
R852 VTAIL.n425 VTAIL.n424 3.49141
R853 VTAIL.n401 VTAIL.n383 3.49141
R854 VTAIL.n358 VTAIL.n270 3.49141
R855 VTAIL.n335 VTAIL.n334 3.49141
R856 VTAIL.n311 VTAIL.n293 3.49141
R857 VTAIL.n669 VTAIL.n654 2.71565
R858 VTAIL.n697 VTAIL.n640 2.71565
R859 VTAIL.n716 VTAIL.n715 2.71565
R860 VTAIL.n39 VTAIL.n24 2.71565
R861 VTAIL.n67 VTAIL.n10 2.71565
R862 VTAIL.n86 VTAIL.n85 2.71565
R863 VTAIL.n129 VTAIL.n114 2.71565
R864 VTAIL.n157 VTAIL.n100 2.71565
R865 VTAIL.n176 VTAIL.n175 2.71565
R866 VTAIL.n219 VTAIL.n204 2.71565
R867 VTAIL.n247 VTAIL.n190 2.71565
R868 VTAIL.n266 VTAIL.n265 2.71565
R869 VTAIL.n626 VTAIL.n625 2.71565
R870 VTAIL.n608 VTAIL.n551 2.71565
R871 VTAIL.n580 VTAIL.n565 2.71565
R872 VTAIL.n536 VTAIL.n535 2.71565
R873 VTAIL.n518 VTAIL.n461 2.71565
R874 VTAIL.n490 VTAIL.n475 2.71565
R875 VTAIL.n446 VTAIL.n445 2.71565
R876 VTAIL.n428 VTAIL.n371 2.71565
R877 VTAIL.n400 VTAIL.n385 2.71565
R878 VTAIL.n356 VTAIL.n355 2.71565
R879 VTAIL.n338 VTAIL.n281 2.71565
R880 VTAIL.n310 VTAIL.n295 2.71565
R881 VTAIL.n449 VTAIL.n359 2.2936
R882 VTAIL.n629 VTAIL.n539 2.2936
R883 VTAIL.n269 VTAIL.n179 2.2936
R884 VTAIL.n666 VTAIL.n665 1.93989
R885 VTAIL.n698 VTAIL.n638 1.93989
R886 VTAIL.n712 VTAIL.n632 1.93989
R887 VTAIL.n36 VTAIL.n35 1.93989
R888 VTAIL.n68 VTAIL.n8 1.93989
R889 VTAIL.n82 VTAIL.n2 1.93989
R890 VTAIL.n126 VTAIL.n125 1.93989
R891 VTAIL.n158 VTAIL.n98 1.93989
R892 VTAIL.n172 VTAIL.n92 1.93989
R893 VTAIL.n216 VTAIL.n215 1.93989
R894 VTAIL.n248 VTAIL.n188 1.93989
R895 VTAIL.n262 VTAIL.n182 1.93989
R896 VTAIL.n622 VTAIL.n542 1.93989
R897 VTAIL.n609 VTAIL.n549 1.93989
R898 VTAIL.n577 VTAIL.n576 1.93989
R899 VTAIL.n532 VTAIL.n452 1.93989
R900 VTAIL.n519 VTAIL.n459 1.93989
R901 VTAIL.n487 VTAIL.n486 1.93989
R902 VTAIL.n442 VTAIL.n362 1.93989
R903 VTAIL.n429 VTAIL.n369 1.93989
R904 VTAIL.n397 VTAIL.n396 1.93989
R905 VTAIL.n352 VTAIL.n272 1.93989
R906 VTAIL.n339 VTAIL.n279 1.93989
R907 VTAIL.n307 VTAIL.n306 1.93989
R908 VTAIL VTAIL.n89 1.20524
R909 VTAIL.n662 VTAIL.n656 1.16414
R910 VTAIL.n703 VTAIL.n701 1.16414
R911 VTAIL.n711 VTAIL.n634 1.16414
R912 VTAIL.n32 VTAIL.n26 1.16414
R913 VTAIL.n73 VTAIL.n71 1.16414
R914 VTAIL.n81 VTAIL.n4 1.16414
R915 VTAIL.n122 VTAIL.n116 1.16414
R916 VTAIL.n163 VTAIL.n161 1.16414
R917 VTAIL.n171 VTAIL.n94 1.16414
R918 VTAIL.n212 VTAIL.n206 1.16414
R919 VTAIL.n253 VTAIL.n251 1.16414
R920 VTAIL.n261 VTAIL.n184 1.16414
R921 VTAIL.n621 VTAIL.n544 1.16414
R922 VTAIL.n613 VTAIL.n612 1.16414
R923 VTAIL.n573 VTAIL.n567 1.16414
R924 VTAIL.n531 VTAIL.n454 1.16414
R925 VTAIL.n523 VTAIL.n522 1.16414
R926 VTAIL.n483 VTAIL.n477 1.16414
R927 VTAIL.n441 VTAIL.n364 1.16414
R928 VTAIL.n433 VTAIL.n432 1.16414
R929 VTAIL.n393 VTAIL.n387 1.16414
R930 VTAIL.n351 VTAIL.n274 1.16414
R931 VTAIL.n343 VTAIL.n342 1.16414
R932 VTAIL.n303 VTAIL.n297 1.16414
R933 VTAIL VTAIL.n719 1.08886
R934 VTAIL.n539 VTAIL.n449 0.470328
R935 VTAIL.n179 VTAIL.n89 0.470328
R936 VTAIL.n661 VTAIL.n658 0.388379
R937 VTAIL.n702 VTAIL.n636 0.388379
R938 VTAIL.n708 VTAIL.n707 0.388379
R939 VTAIL.n31 VTAIL.n28 0.388379
R940 VTAIL.n72 VTAIL.n6 0.388379
R941 VTAIL.n78 VTAIL.n77 0.388379
R942 VTAIL.n121 VTAIL.n118 0.388379
R943 VTAIL.n162 VTAIL.n96 0.388379
R944 VTAIL.n168 VTAIL.n167 0.388379
R945 VTAIL.n211 VTAIL.n208 0.388379
R946 VTAIL.n252 VTAIL.n186 0.388379
R947 VTAIL.n258 VTAIL.n257 0.388379
R948 VTAIL.n618 VTAIL.n617 0.388379
R949 VTAIL.n548 VTAIL.n546 0.388379
R950 VTAIL.n572 VTAIL.n569 0.388379
R951 VTAIL.n528 VTAIL.n527 0.388379
R952 VTAIL.n458 VTAIL.n456 0.388379
R953 VTAIL.n482 VTAIL.n479 0.388379
R954 VTAIL.n438 VTAIL.n437 0.388379
R955 VTAIL.n368 VTAIL.n366 0.388379
R956 VTAIL.n392 VTAIL.n389 0.388379
R957 VTAIL.n348 VTAIL.n347 0.388379
R958 VTAIL.n278 VTAIL.n276 0.388379
R959 VTAIL.n302 VTAIL.n299 0.388379
R960 VTAIL.n660 VTAIL.n655 0.155672
R961 VTAIL.n667 VTAIL.n655 0.155672
R962 VTAIL.n668 VTAIL.n667 0.155672
R963 VTAIL.n668 VTAIL.n651 0.155672
R964 VTAIL.n675 VTAIL.n651 0.155672
R965 VTAIL.n676 VTAIL.n675 0.155672
R966 VTAIL.n676 VTAIL.n647 0.155672
R967 VTAIL.n683 VTAIL.n647 0.155672
R968 VTAIL.n684 VTAIL.n683 0.155672
R969 VTAIL.n684 VTAIL.n643 0.155672
R970 VTAIL.n691 VTAIL.n643 0.155672
R971 VTAIL.n692 VTAIL.n691 0.155672
R972 VTAIL.n692 VTAIL.n639 0.155672
R973 VTAIL.n699 VTAIL.n639 0.155672
R974 VTAIL.n700 VTAIL.n699 0.155672
R975 VTAIL.n700 VTAIL.n635 0.155672
R976 VTAIL.n709 VTAIL.n635 0.155672
R977 VTAIL.n710 VTAIL.n709 0.155672
R978 VTAIL.n710 VTAIL.n631 0.155672
R979 VTAIL.n717 VTAIL.n631 0.155672
R980 VTAIL.n30 VTAIL.n25 0.155672
R981 VTAIL.n37 VTAIL.n25 0.155672
R982 VTAIL.n38 VTAIL.n37 0.155672
R983 VTAIL.n38 VTAIL.n21 0.155672
R984 VTAIL.n45 VTAIL.n21 0.155672
R985 VTAIL.n46 VTAIL.n45 0.155672
R986 VTAIL.n46 VTAIL.n17 0.155672
R987 VTAIL.n53 VTAIL.n17 0.155672
R988 VTAIL.n54 VTAIL.n53 0.155672
R989 VTAIL.n54 VTAIL.n13 0.155672
R990 VTAIL.n61 VTAIL.n13 0.155672
R991 VTAIL.n62 VTAIL.n61 0.155672
R992 VTAIL.n62 VTAIL.n9 0.155672
R993 VTAIL.n69 VTAIL.n9 0.155672
R994 VTAIL.n70 VTAIL.n69 0.155672
R995 VTAIL.n70 VTAIL.n5 0.155672
R996 VTAIL.n79 VTAIL.n5 0.155672
R997 VTAIL.n80 VTAIL.n79 0.155672
R998 VTAIL.n80 VTAIL.n1 0.155672
R999 VTAIL.n87 VTAIL.n1 0.155672
R1000 VTAIL.n120 VTAIL.n115 0.155672
R1001 VTAIL.n127 VTAIL.n115 0.155672
R1002 VTAIL.n128 VTAIL.n127 0.155672
R1003 VTAIL.n128 VTAIL.n111 0.155672
R1004 VTAIL.n135 VTAIL.n111 0.155672
R1005 VTAIL.n136 VTAIL.n135 0.155672
R1006 VTAIL.n136 VTAIL.n107 0.155672
R1007 VTAIL.n143 VTAIL.n107 0.155672
R1008 VTAIL.n144 VTAIL.n143 0.155672
R1009 VTAIL.n144 VTAIL.n103 0.155672
R1010 VTAIL.n151 VTAIL.n103 0.155672
R1011 VTAIL.n152 VTAIL.n151 0.155672
R1012 VTAIL.n152 VTAIL.n99 0.155672
R1013 VTAIL.n159 VTAIL.n99 0.155672
R1014 VTAIL.n160 VTAIL.n159 0.155672
R1015 VTAIL.n160 VTAIL.n95 0.155672
R1016 VTAIL.n169 VTAIL.n95 0.155672
R1017 VTAIL.n170 VTAIL.n169 0.155672
R1018 VTAIL.n170 VTAIL.n91 0.155672
R1019 VTAIL.n177 VTAIL.n91 0.155672
R1020 VTAIL.n210 VTAIL.n205 0.155672
R1021 VTAIL.n217 VTAIL.n205 0.155672
R1022 VTAIL.n218 VTAIL.n217 0.155672
R1023 VTAIL.n218 VTAIL.n201 0.155672
R1024 VTAIL.n225 VTAIL.n201 0.155672
R1025 VTAIL.n226 VTAIL.n225 0.155672
R1026 VTAIL.n226 VTAIL.n197 0.155672
R1027 VTAIL.n233 VTAIL.n197 0.155672
R1028 VTAIL.n234 VTAIL.n233 0.155672
R1029 VTAIL.n234 VTAIL.n193 0.155672
R1030 VTAIL.n241 VTAIL.n193 0.155672
R1031 VTAIL.n242 VTAIL.n241 0.155672
R1032 VTAIL.n242 VTAIL.n189 0.155672
R1033 VTAIL.n249 VTAIL.n189 0.155672
R1034 VTAIL.n250 VTAIL.n249 0.155672
R1035 VTAIL.n250 VTAIL.n185 0.155672
R1036 VTAIL.n259 VTAIL.n185 0.155672
R1037 VTAIL.n260 VTAIL.n259 0.155672
R1038 VTAIL.n260 VTAIL.n181 0.155672
R1039 VTAIL.n267 VTAIL.n181 0.155672
R1040 VTAIL.n627 VTAIL.n541 0.155672
R1041 VTAIL.n620 VTAIL.n541 0.155672
R1042 VTAIL.n620 VTAIL.n619 0.155672
R1043 VTAIL.n619 VTAIL.n545 0.155672
R1044 VTAIL.n611 VTAIL.n545 0.155672
R1045 VTAIL.n611 VTAIL.n610 0.155672
R1046 VTAIL.n610 VTAIL.n550 0.155672
R1047 VTAIL.n603 VTAIL.n550 0.155672
R1048 VTAIL.n603 VTAIL.n602 0.155672
R1049 VTAIL.n602 VTAIL.n554 0.155672
R1050 VTAIL.n595 VTAIL.n554 0.155672
R1051 VTAIL.n595 VTAIL.n594 0.155672
R1052 VTAIL.n594 VTAIL.n558 0.155672
R1053 VTAIL.n587 VTAIL.n558 0.155672
R1054 VTAIL.n587 VTAIL.n586 0.155672
R1055 VTAIL.n586 VTAIL.n562 0.155672
R1056 VTAIL.n579 VTAIL.n562 0.155672
R1057 VTAIL.n579 VTAIL.n578 0.155672
R1058 VTAIL.n578 VTAIL.n566 0.155672
R1059 VTAIL.n571 VTAIL.n566 0.155672
R1060 VTAIL.n537 VTAIL.n451 0.155672
R1061 VTAIL.n530 VTAIL.n451 0.155672
R1062 VTAIL.n530 VTAIL.n529 0.155672
R1063 VTAIL.n529 VTAIL.n455 0.155672
R1064 VTAIL.n521 VTAIL.n455 0.155672
R1065 VTAIL.n521 VTAIL.n520 0.155672
R1066 VTAIL.n520 VTAIL.n460 0.155672
R1067 VTAIL.n513 VTAIL.n460 0.155672
R1068 VTAIL.n513 VTAIL.n512 0.155672
R1069 VTAIL.n512 VTAIL.n464 0.155672
R1070 VTAIL.n505 VTAIL.n464 0.155672
R1071 VTAIL.n505 VTAIL.n504 0.155672
R1072 VTAIL.n504 VTAIL.n468 0.155672
R1073 VTAIL.n497 VTAIL.n468 0.155672
R1074 VTAIL.n497 VTAIL.n496 0.155672
R1075 VTAIL.n496 VTAIL.n472 0.155672
R1076 VTAIL.n489 VTAIL.n472 0.155672
R1077 VTAIL.n489 VTAIL.n488 0.155672
R1078 VTAIL.n488 VTAIL.n476 0.155672
R1079 VTAIL.n481 VTAIL.n476 0.155672
R1080 VTAIL.n447 VTAIL.n361 0.155672
R1081 VTAIL.n440 VTAIL.n361 0.155672
R1082 VTAIL.n440 VTAIL.n439 0.155672
R1083 VTAIL.n439 VTAIL.n365 0.155672
R1084 VTAIL.n431 VTAIL.n365 0.155672
R1085 VTAIL.n431 VTAIL.n430 0.155672
R1086 VTAIL.n430 VTAIL.n370 0.155672
R1087 VTAIL.n423 VTAIL.n370 0.155672
R1088 VTAIL.n423 VTAIL.n422 0.155672
R1089 VTAIL.n422 VTAIL.n374 0.155672
R1090 VTAIL.n415 VTAIL.n374 0.155672
R1091 VTAIL.n415 VTAIL.n414 0.155672
R1092 VTAIL.n414 VTAIL.n378 0.155672
R1093 VTAIL.n407 VTAIL.n378 0.155672
R1094 VTAIL.n407 VTAIL.n406 0.155672
R1095 VTAIL.n406 VTAIL.n382 0.155672
R1096 VTAIL.n399 VTAIL.n382 0.155672
R1097 VTAIL.n399 VTAIL.n398 0.155672
R1098 VTAIL.n398 VTAIL.n386 0.155672
R1099 VTAIL.n391 VTAIL.n386 0.155672
R1100 VTAIL.n357 VTAIL.n271 0.155672
R1101 VTAIL.n350 VTAIL.n271 0.155672
R1102 VTAIL.n350 VTAIL.n349 0.155672
R1103 VTAIL.n349 VTAIL.n275 0.155672
R1104 VTAIL.n341 VTAIL.n275 0.155672
R1105 VTAIL.n341 VTAIL.n340 0.155672
R1106 VTAIL.n340 VTAIL.n280 0.155672
R1107 VTAIL.n333 VTAIL.n280 0.155672
R1108 VTAIL.n333 VTAIL.n332 0.155672
R1109 VTAIL.n332 VTAIL.n284 0.155672
R1110 VTAIL.n325 VTAIL.n284 0.155672
R1111 VTAIL.n325 VTAIL.n324 0.155672
R1112 VTAIL.n324 VTAIL.n288 0.155672
R1113 VTAIL.n317 VTAIL.n288 0.155672
R1114 VTAIL.n317 VTAIL.n316 0.155672
R1115 VTAIL.n316 VTAIL.n292 0.155672
R1116 VTAIL.n309 VTAIL.n292 0.155672
R1117 VTAIL.n309 VTAIL.n308 0.155672
R1118 VTAIL.n308 VTAIL.n296 0.155672
R1119 VTAIL.n301 VTAIL.n296 0.155672
R1120 B.n841 B.n840 585
R1121 B.n350 B.n118 585
R1122 B.n349 B.n348 585
R1123 B.n347 B.n346 585
R1124 B.n345 B.n344 585
R1125 B.n343 B.n342 585
R1126 B.n341 B.n340 585
R1127 B.n339 B.n338 585
R1128 B.n337 B.n336 585
R1129 B.n335 B.n334 585
R1130 B.n333 B.n332 585
R1131 B.n331 B.n330 585
R1132 B.n329 B.n328 585
R1133 B.n327 B.n326 585
R1134 B.n325 B.n324 585
R1135 B.n323 B.n322 585
R1136 B.n321 B.n320 585
R1137 B.n319 B.n318 585
R1138 B.n317 B.n316 585
R1139 B.n315 B.n314 585
R1140 B.n313 B.n312 585
R1141 B.n311 B.n310 585
R1142 B.n309 B.n308 585
R1143 B.n307 B.n306 585
R1144 B.n305 B.n304 585
R1145 B.n303 B.n302 585
R1146 B.n301 B.n300 585
R1147 B.n299 B.n298 585
R1148 B.n297 B.n296 585
R1149 B.n295 B.n294 585
R1150 B.n293 B.n292 585
R1151 B.n291 B.n290 585
R1152 B.n289 B.n288 585
R1153 B.n287 B.n286 585
R1154 B.n285 B.n284 585
R1155 B.n283 B.n282 585
R1156 B.n281 B.n280 585
R1157 B.n279 B.n278 585
R1158 B.n277 B.n276 585
R1159 B.n275 B.n274 585
R1160 B.n273 B.n272 585
R1161 B.n271 B.n270 585
R1162 B.n269 B.n268 585
R1163 B.n267 B.n266 585
R1164 B.n265 B.n264 585
R1165 B.n263 B.n262 585
R1166 B.n261 B.n260 585
R1167 B.n259 B.n258 585
R1168 B.n257 B.n256 585
R1169 B.n255 B.n254 585
R1170 B.n253 B.n252 585
R1171 B.n251 B.n250 585
R1172 B.n249 B.n248 585
R1173 B.n246 B.n245 585
R1174 B.n244 B.n243 585
R1175 B.n242 B.n241 585
R1176 B.n240 B.n239 585
R1177 B.n238 B.n237 585
R1178 B.n236 B.n235 585
R1179 B.n234 B.n233 585
R1180 B.n232 B.n231 585
R1181 B.n230 B.n229 585
R1182 B.n228 B.n227 585
R1183 B.n225 B.n224 585
R1184 B.n223 B.n222 585
R1185 B.n221 B.n220 585
R1186 B.n219 B.n218 585
R1187 B.n217 B.n216 585
R1188 B.n215 B.n214 585
R1189 B.n213 B.n212 585
R1190 B.n211 B.n210 585
R1191 B.n209 B.n208 585
R1192 B.n207 B.n206 585
R1193 B.n205 B.n204 585
R1194 B.n203 B.n202 585
R1195 B.n201 B.n200 585
R1196 B.n199 B.n198 585
R1197 B.n197 B.n196 585
R1198 B.n195 B.n194 585
R1199 B.n193 B.n192 585
R1200 B.n191 B.n190 585
R1201 B.n189 B.n188 585
R1202 B.n187 B.n186 585
R1203 B.n185 B.n184 585
R1204 B.n183 B.n182 585
R1205 B.n181 B.n180 585
R1206 B.n179 B.n178 585
R1207 B.n177 B.n176 585
R1208 B.n175 B.n174 585
R1209 B.n173 B.n172 585
R1210 B.n171 B.n170 585
R1211 B.n169 B.n168 585
R1212 B.n167 B.n166 585
R1213 B.n165 B.n164 585
R1214 B.n163 B.n162 585
R1215 B.n161 B.n160 585
R1216 B.n159 B.n158 585
R1217 B.n157 B.n156 585
R1218 B.n155 B.n154 585
R1219 B.n153 B.n152 585
R1220 B.n151 B.n150 585
R1221 B.n149 B.n148 585
R1222 B.n147 B.n146 585
R1223 B.n145 B.n144 585
R1224 B.n143 B.n142 585
R1225 B.n141 B.n140 585
R1226 B.n139 B.n138 585
R1227 B.n137 B.n136 585
R1228 B.n135 B.n134 585
R1229 B.n133 B.n132 585
R1230 B.n131 B.n130 585
R1231 B.n129 B.n128 585
R1232 B.n127 B.n126 585
R1233 B.n125 B.n124 585
R1234 B.n61 B.n60 585
R1235 B.n846 B.n845 585
R1236 B.n839 B.n119 585
R1237 B.n119 B.n58 585
R1238 B.n838 B.n57 585
R1239 B.n850 B.n57 585
R1240 B.n837 B.n56 585
R1241 B.n851 B.n56 585
R1242 B.n836 B.n55 585
R1243 B.n852 B.n55 585
R1244 B.n835 B.n834 585
R1245 B.n834 B.n51 585
R1246 B.n833 B.n50 585
R1247 B.n858 B.n50 585
R1248 B.n832 B.n49 585
R1249 B.n859 B.n49 585
R1250 B.n831 B.n48 585
R1251 B.n860 B.n48 585
R1252 B.n830 B.n829 585
R1253 B.n829 B.n44 585
R1254 B.n828 B.n43 585
R1255 B.n866 B.n43 585
R1256 B.n827 B.n42 585
R1257 B.n867 B.n42 585
R1258 B.n826 B.n41 585
R1259 B.n868 B.n41 585
R1260 B.n825 B.n824 585
R1261 B.n824 B.n37 585
R1262 B.n823 B.n36 585
R1263 B.n874 B.n36 585
R1264 B.n822 B.n35 585
R1265 B.n875 B.n35 585
R1266 B.n821 B.n34 585
R1267 B.n876 B.n34 585
R1268 B.n820 B.n819 585
R1269 B.n819 B.n30 585
R1270 B.n818 B.n29 585
R1271 B.n882 B.n29 585
R1272 B.n817 B.n28 585
R1273 B.n883 B.n28 585
R1274 B.n816 B.n27 585
R1275 B.n884 B.n27 585
R1276 B.n815 B.n814 585
R1277 B.n814 B.n23 585
R1278 B.n813 B.n22 585
R1279 B.n890 B.n22 585
R1280 B.n812 B.n21 585
R1281 B.n891 B.n21 585
R1282 B.n811 B.n20 585
R1283 B.n892 B.n20 585
R1284 B.n810 B.n809 585
R1285 B.n809 B.n16 585
R1286 B.n808 B.n15 585
R1287 B.n898 B.n15 585
R1288 B.n807 B.n14 585
R1289 B.n899 B.n14 585
R1290 B.n806 B.n13 585
R1291 B.n900 B.n13 585
R1292 B.n805 B.n804 585
R1293 B.n804 B.n12 585
R1294 B.n803 B.n802 585
R1295 B.n803 B.n8 585
R1296 B.n801 B.n7 585
R1297 B.n907 B.n7 585
R1298 B.n800 B.n6 585
R1299 B.n908 B.n6 585
R1300 B.n799 B.n5 585
R1301 B.n909 B.n5 585
R1302 B.n798 B.n797 585
R1303 B.n797 B.n4 585
R1304 B.n796 B.n351 585
R1305 B.n796 B.n795 585
R1306 B.n786 B.n352 585
R1307 B.n353 B.n352 585
R1308 B.n788 B.n787 585
R1309 B.n789 B.n788 585
R1310 B.n785 B.n358 585
R1311 B.n358 B.n357 585
R1312 B.n784 B.n783 585
R1313 B.n783 B.n782 585
R1314 B.n360 B.n359 585
R1315 B.n361 B.n360 585
R1316 B.n775 B.n774 585
R1317 B.n776 B.n775 585
R1318 B.n773 B.n366 585
R1319 B.n366 B.n365 585
R1320 B.n772 B.n771 585
R1321 B.n771 B.n770 585
R1322 B.n368 B.n367 585
R1323 B.n369 B.n368 585
R1324 B.n763 B.n762 585
R1325 B.n764 B.n763 585
R1326 B.n761 B.n373 585
R1327 B.n377 B.n373 585
R1328 B.n760 B.n759 585
R1329 B.n759 B.n758 585
R1330 B.n375 B.n374 585
R1331 B.n376 B.n375 585
R1332 B.n751 B.n750 585
R1333 B.n752 B.n751 585
R1334 B.n749 B.n382 585
R1335 B.n382 B.n381 585
R1336 B.n748 B.n747 585
R1337 B.n747 B.n746 585
R1338 B.n384 B.n383 585
R1339 B.n385 B.n384 585
R1340 B.n739 B.n738 585
R1341 B.n740 B.n739 585
R1342 B.n737 B.n390 585
R1343 B.n390 B.n389 585
R1344 B.n736 B.n735 585
R1345 B.n735 B.n734 585
R1346 B.n392 B.n391 585
R1347 B.n393 B.n392 585
R1348 B.n727 B.n726 585
R1349 B.n728 B.n727 585
R1350 B.n725 B.n398 585
R1351 B.n398 B.n397 585
R1352 B.n724 B.n723 585
R1353 B.n723 B.n722 585
R1354 B.n400 B.n399 585
R1355 B.n401 B.n400 585
R1356 B.n715 B.n714 585
R1357 B.n716 B.n715 585
R1358 B.n713 B.n406 585
R1359 B.n406 B.n405 585
R1360 B.n712 B.n711 585
R1361 B.n711 B.n710 585
R1362 B.n408 B.n407 585
R1363 B.n409 B.n408 585
R1364 B.n706 B.n705 585
R1365 B.n412 B.n411 585
R1366 B.n702 B.n701 585
R1367 B.n703 B.n702 585
R1368 B.n700 B.n470 585
R1369 B.n699 B.n698 585
R1370 B.n697 B.n696 585
R1371 B.n695 B.n694 585
R1372 B.n693 B.n692 585
R1373 B.n691 B.n690 585
R1374 B.n689 B.n688 585
R1375 B.n687 B.n686 585
R1376 B.n685 B.n684 585
R1377 B.n683 B.n682 585
R1378 B.n681 B.n680 585
R1379 B.n679 B.n678 585
R1380 B.n677 B.n676 585
R1381 B.n675 B.n674 585
R1382 B.n673 B.n672 585
R1383 B.n671 B.n670 585
R1384 B.n669 B.n668 585
R1385 B.n667 B.n666 585
R1386 B.n665 B.n664 585
R1387 B.n663 B.n662 585
R1388 B.n661 B.n660 585
R1389 B.n659 B.n658 585
R1390 B.n657 B.n656 585
R1391 B.n655 B.n654 585
R1392 B.n653 B.n652 585
R1393 B.n651 B.n650 585
R1394 B.n649 B.n648 585
R1395 B.n647 B.n646 585
R1396 B.n645 B.n644 585
R1397 B.n643 B.n642 585
R1398 B.n641 B.n640 585
R1399 B.n639 B.n638 585
R1400 B.n637 B.n636 585
R1401 B.n635 B.n634 585
R1402 B.n633 B.n632 585
R1403 B.n631 B.n630 585
R1404 B.n629 B.n628 585
R1405 B.n627 B.n626 585
R1406 B.n625 B.n624 585
R1407 B.n623 B.n622 585
R1408 B.n621 B.n620 585
R1409 B.n619 B.n618 585
R1410 B.n617 B.n616 585
R1411 B.n615 B.n614 585
R1412 B.n613 B.n612 585
R1413 B.n611 B.n610 585
R1414 B.n609 B.n608 585
R1415 B.n607 B.n606 585
R1416 B.n605 B.n604 585
R1417 B.n603 B.n602 585
R1418 B.n601 B.n600 585
R1419 B.n599 B.n598 585
R1420 B.n597 B.n596 585
R1421 B.n595 B.n594 585
R1422 B.n593 B.n592 585
R1423 B.n591 B.n590 585
R1424 B.n589 B.n588 585
R1425 B.n587 B.n586 585
R1426 B.n585 B.n584 585
R1427 B.n583 B.n582 585
R1428 B.n581 B.n580 585
R1429 B.n579 B.n578 585
R1430 B.n577 B.n576 585
R1431 B.n575 B.n574 585
R1432 B.n573 B.n572 585
R1433 B.n571 B.n570 585
R1434 B.n569 B.n568 585
R1435 B.n567 B.n566 585
R1436 B.n565 B.n564 585
R1437 B.n563 B.n562 585
R1438 B.n561 B.n560 585
R1439 B.n559 B.n558 585
R1440 B.n557 B.n556 585
R1441 B.n555 B.n554 585
R1442 B.n553 B.n552 585
R1443 B.n551 B.n550 585
R1444 B.n549 B.n548 585
R1445 B.n547 B.n546 585
R1446 B.n545 B.n544 585
R1447 B.n543 B.n542 585
R1448 B.n541 B.n540 585
R1449 B.n539 B.n538 585
R1450 B.n537 B.n536 585
R1451 B.n535 B.n534 585
R1452 B.n533 B.n532 585
R1453 B.n531 B.n530 585
R1454 B.n529 B.n528 585
R1455 B.n527 B.n526 585
R1456 B.n525 B.n524 585
R1457 B.n523 B.n522 585
R1458 B.n521 B.n520 585
R1459 B.n519 B.n518 585
R1460 B.n517 B.n516 585
R1461 B.n515 B.n514 585
R1462 B.n513 B.n512 585
R1463 B.n511 B.n510 585
R1464 B.n509 B.n508 585
R1465 B.n507 B.n506 585
R1466 B.n505 B.n504 585
R1467 B.n503 B.n502 585
R1468 B.n501 B.n500 585
R1469 B.n499 B.n498 585
R1470 B.n497 B.n496 585
R1471 B.n495 B.n494 585
R1472 B.n493 B.n492 585
R1473 B.n491 B.n490 585
R1474 B.n489 B.n488 585
R1475 B.n487 B.n486 585
R1476 B.n485 B.n484 585
R1477 B.n483 B.n482 585
R1478 B.n481 B.n480 585
R1479 B.n479 B.n478 585
R1480 B.n477 B.n469 585
R1481 B.n703 B.n469 585
R1482 B.n707 B.n410 585
R1483 B.n410 B.n409 585
R1484 B.n709 B.n708 585
R1485 B.n710 B.n709 585
R1486 B.n404 B.n403 585
R1487 B.n405 B.n404 585
R1488 B.n718 B.n717 585
R1489 B.n717 B.n716 585
R1490 B.n719 B.n402 585
R1491 B.n402 B.n401 585
R1492 B.n721 B.n720 585
R1493 B.n722 B.n721 585
R1494 B.n396 B.n395 585
R1495 B.n397 B.n396 585
R1496 B.n730 B.n729 585
R1497 B.n729 B.n728 585
R1498 B.n731 B.n394 585
R1499 B.n394 B.n393 585
R1500 B.n733 B.n732 585
R1501 B.n734 B.n733 585
R1502 B.n388 B.n387 585
R1503 B.n389 B.n388 585
R1504 B.n742 B.n741 585
R1505 B.n741 B.n740 585
R1506 B.n743 B.n386 585
R1507 B.n386 B.n385 585
R1508 B.n745 B.n744 585
R1509 B.n746 B.n745 585
R1510 B.n380 B.n379 585
R1511 B.n381 B.n380 585
R1512 B.n754 B.n753 585
R1513 B.n753 B.n752 585
R1514 B.n755 B.n378 585
R1515 B.n378 B.n376 585
R1516 B.n757 B.n756 585
R1517 B.n758 B.n757 585
R1518 B.n372 B.n371 585
R1519 B.n377 B.n372 585
R1520 B.n766 B.n765 585
R1521 B.n765 B.n764 585
R1522 B.n767 B.n370 585
R1523 B.n370 B.n369 585
R1524 B.n769 B.n768 585
R1525 B.n770 B.n769 585
R1526 B.n364 B.n363 585
R1527 B.n365 B.n364 585
R1528 B.n778 B.n777 585
R1529 B.n777 B.n776 585
R1530 B.n779 B.n362 585
R1531 B.n362 B.n361 585
R1532 B.n781 B.n780 585
R1533 B.n782 B.n781 585
R1534 B.n356 B.n355 585
R1535 B.n357 B.n356 585
R1536 B.n791 B.n790 585
R1537 B.n790 B.n789 585
R1538 B.n792 B.n354 585
R1539 B.n354 B.n353 585
R1540 B.n794 B.n793 585
R1541 B.n795 B.n794 585
R1542 B.n3 B.n0 585
R1543 B.n4 B.n3 585
R1544 B.n906 B.n1 585
R1545 B.n907 B.n906 585
R1546 B.n905 B.n904 585
R1547 B.n905 B.n8 585
R1548 B.n903 B.n9 585
R1549 B.n12 B.n9 585
R1550 B.n902 B.n901 585
R1551 B.n901 B.n900 585
R1552 B.n11 B.n10 585
R1553 B.n899 B.n11 585
R1554 B.n897 B.n896 585
R1555 B.n898 B.n897 585
R1556 B.n895 B.n17 585
R1557 B.n17 B.n16 585
R1558 B.n894 B.n893 585
R1559 B.n893 B.n892 585
R1560 B.n19 B.n18 585
R1561 B.n891 B.n19 585
R1562 B.n889 B.n888 585
R1563 B.n890 B.n889 585
R1564 B.n887 B.n24 585
R1565 B.n24 B.n23 585
R1566 B.n886 B.n885 585
R1567 B.n885 B.n884 585
R1568 B.n26 B.n25 585
R1569 B.n883 B.n26 585
R1570 B.n881 B.n880 585
R1571 B.n882 B.n881 585
R1572 B.n879 B.n31 585
R1573 B.n31 B.n30 585
R1574 B.n878 B.n877 585
R1575 B.n877 B.n876 585
R1576 B.n33 B.n32 585
R1577 B.n875 B.n33 585
R1578 B.n873 B.n872 585
R1579 B.n874 B.n873 585
R1580 B.n871 B.n38 585
R1581 B.n38 B.n37 585
R1582 B.n870 B.n869 585
R1583 B.n869 B.n868 585
R1584 B.n40 B.n39 585
R1585 B.n867 B.n40 585
R1586 B.n865 B.n864 585
R1587 B.n866 B.n865 585
R1588 B.n863 B.n45 585
R1589 B.n45 B.n44 585
R1590 B.n862 B.n861 585
R1591 B.n861 B.n860 585
R1592 B.n47 B.n46 585
R1593 B.n859 B.n47 585
R1594 B.n857 B.n856 585
R1595 B.n858 B.n857 585
R1596 B.n855 B.n52 585
R1597 B.n52 B.n51 585
R1598 B.n854 B.n853 585
R1599 B.n853 B.n852 585
R1600 B.n54 B.n53 585
R1601 B.n851 B.n54 585
R1602 B.n849 B.n848 585
R1603 B.n850 B.n849 585
R1604 B.n847 B.n59 585
R1605 B.n59 B.n58 585
R1606 B.n910 B.n909 585
R1607 B.n908 B.n2 585
R1608 B.n845 B.n59 535.745
R1609 B.n841 B.n119 535.745
R1610 B.n469 B.n408 535.745
R1611 B.n705 B.n410 535.745
R1612 B.n122 B.t6 402.318
R1613 B.n120 B.t16 402.318
R1614 B.n474 B.t14 402.318
R1615 B.n471 B.t11 402.318
R1616 B.n120 B.t15 373.647
R1617 B.n474 B.t12 373.647
R1618 B.n122 B.t4 373.293
R1619 B.n471 B.t8 373.293
R1620 B.n121 B.t17 350.731
R1621 B.n475 B.t13 350.731
R1622 B.n123 B.t7 350.731
R1623 B.n472 B.t10 350.731
R1624 B.n843 B.n842 256.663
R1625 B.n843 B.n117 256.663
R1626 B.n843 B.n116 256.663
R1627 B.n843 B.n115 256.663
R1628 B.n843 B.n114 256.663
R1629 B.n843 B.n113 256.663
R1630 B.n843 B.n112 256.663
R1631 B.n843 B.n111 256.663
R1632 B.n843 B.n110 256.663
R1633 B.n843 B.n109 256.663
R1634 B.n843 B.n108 256.663
R1635 B.n843 B.n107 256.663
R1636 B.n843 B.n106 256.663
R1637 B.n843 B.n105 256.663
R1638 B.n843 B.n104 256.663
R1639 B.n843 B.n103 256.663
R1640 B.n843 B.n102 256.663
R1641 B.n843 B.n101 256.663
R1642 B.n843 B.n100 256.663
R1643 B.n843 B.n99 256.663
R1644 B.n843 B.n98 256.663
R1645 B.n843 B.n97 256.663
R1646 B.n843 B.n96 256.663
R1647 B.n843 B.n95 256.663
R1648 B.n843 B.n94 256.663
R1649 B.n843 B.n93 256.663
R1650 B.n843 B.n92 256.663
R1651 B.n843 B.n91 256.663
R1652 B.n843 B.n90 256.663
R1653 B.n843 B.n89 256.663
R1654 B.n843 B.n88 256.663
R1655 B.n843 B.n87 256.663
R1656 B.n843 B.n86 256.663
R1657 B.n843 B.n85 256.663
R1658 B.n843 B.n84 256.663
R1659 B.n843 B.n83 256.663
R1660 B.n843 B.n82 256.663
R1661 B.n843 B.n81 256.663
R1662 B.n843 B.n80 256.663
R1663 B.n843 B.n79 256.663
R1664 B.n843 B.n78 256.663
R1665 B.n843 B.n77 256.663
R1666 B.n843 B.n76 256.663
R1667 B.n843 B.n75 256.663
R1668 B.n843 B.n74 256.663
R1669 B.n843 B.n73 256.663
R1670 B.n843 B.n72 256.663
R1671 B.n843 B.n71 256.663
R1672 B.n843 B.n70 256.663
R1673 B.n843 B.n69 256.663
R1674 B.n843 B.n68 256.663
R1675 B.n843 B.n67 256.663
R1676 B.n843 B.n66 256.663
R1677 B.n843 B.n65 256.663
R1678 B.n843 B.n64 256.663
R1679 B.n843 B.n63 256.663
R1680 B.n843 B.n62 256.663
R1681 B.n844 B.n843 256.663
R1682 B.n704 B.n703 256.663
R1683 B.n703 B.n413 256.663
R1684 B.n703 B.n414 256.663
R1685 B.n703 B.n415 256.663
R1686 B.n703 B.n416 256.663
R1687 B.n703 B.n417 256.663
R1688 B.n703 B.n418 256.663
R1689 B.n703 B.n419 256.663
R1690 B.n703 B.n420 256.663
R1691 B.n703 B.n421 256.663
R1692 B.n703 B.n422 256.663
R1693 B.n703 B.n423 256.663
R1694 B.n703 B.n424 256.663
R1695 B.n703 B.n425 256.663
R1696 B.n703 B.n426 256.663
R1697 B.n703 B.n427 256.663
R1698 B.n703 B.n428 256.663
R1699 B.n703 B.n429 256.663
R1700 B.n703 B.n430 256.663
R1701 B.n703 B.n431 256.663
R1702 B.n703 B.n432 256.663
R1703 B.n703 B.n433 256.663
R1704 B.n703 B.n434 256.663
R1705 B.n703 B.n435 256.663
R1706 B.n703 B.n436 256.663
R1707 B.n703 B.n437 256.663
R1708 B.n703 B.n438 256.663
R1709 B.n703 B.n439 256.663
R1710 B.n703 B.n440 256.663
R1711 B.n703 B.n441 256.663
R1712 B.n703 B.n442 256.663
R1713 B.n703 B.n443 256.663
R1714 B.n703 B.n444 256.663
R1715 B.n703 B.n445 256.663
R1716 B.n703 B.n446 256.663
R1717 B.n703 B.n447 256.663
R1718 B.n703 B.n448 256.663
R1719 B.n703 B.n449 256.663
R1720 B.n703 B.n450 256.663
R1721 B.n703 B.n451 256.663
R1722 B.n703 B.n452 256.663
R1723 B.n703 B.n453 256.663
R1724 B.n703 B.n454 256.663
R1725 B.n703 B.n455 256.663
R1726 B.n703 B.n456 256.663
R1727 B.n703 B.n457 256.663
R1728 B.n703 B.n458 256.663
R1729 B.n703 B.n459 256.663
R1730 B.n703 B.n460 256.663
R1731 B.n703 B.n461 256.663
R1732 B.n703 B.n462 256.663
R1733 B.n703 B.n463 256.663
R1734 B.n703 B.n464 256.663
R1735 B.n703 B.n465 256.663
R1736 B.n703 B.n466 256.663
R1737 B.n703 B.n467 256.663
R1738 B.n703 B.n468 256.663
R1739 B.n912 B.n911 256.663
R1740 B.n124 B.n61 163.367
R1741 B.n128 B.n127 163.367
R1742 B.n132 B.n131 163.367
R1743 B.n136 B.n135 163.367
R1744 B.n140 B.n139 163.367
R1745 B.n144 B.n143 163.367
R1746 B.n148 B.n147 163.367
R1747 B.n152 B.n151 163.367
R1748 B.n156 B.n155 163.367
R1749 B.n160 B.n159 163.367
R1750 B.n164 B.n163 163.367
R1751 B.n168 B.n167 163.367
R1752 B.n172 B.n171 163.367
R1753 B.n176 B.n175 163.367
R1754 B.n180 B.n179 163.367
R1755 B.n184 B.n183 163.367
R1756 B.n188 B.n187 163.367
R1757 B.n192 B.n191 163.367
R1758 B.n196 B.n195 163.367
R1759 B.n200 B.n199 163.367
R1760 B.n204 B.n203 163.367
R1761 B.n208 B.n207 163.367
R1762 B.n212 B.n211 163.367
R1763 B.n216 B.n215 163.367
R1764 B.n220 B.n219 163.367
R1765 B.n224 B.n223 163.367
R1766 B.n229 B.n228 163.367
R1767 B.n233 B.n232 163.367
R1768 B.n237 B.n236 163.367
R1769 B.n241 B.n240 163.367
R1770 B.n245 B.n244 163.367
R1771 B.n250 B.n249 163.367
R1772 B.n254 B.n253 163.367
R1773 B.n258 B.n257 163.367
R1774 B.n262 B.n261 163.367
R1775 B.n266 B.n265 163.367
R1776 B.n270 B.n269 163.367
R1777 B.n274 B.n273 163.367
R1778 B.n278 B.n277 163.367
R1779 B.n282 B.n281 163.367
R1780 B.n286 B.n285 163.367
R1781 B.n290 B.n289 163.367
R1782 B.n294 B.n293 163.367
R1783 B.n298 B.n297 163.367
R1784 B.n302 B.n301 163.367
R1785 B.n306 B.n305 163.367
R1786 B.n310 B.n309 163.367
R1787 B.n314 B.n313 163.367
R1788 B.n318 B.n317 163.367
R1789 B.n322 B.n321 163.367
R1790 B.n326 B.n325 163.367
R1791 B.n330 B.n329 163.367
R1792 B.n334 B.n333 163.367
R1793 B.n338 B.n337 163.367
R1794 B.n342 B.n341 163.367
R1795 B.n346 B.n345 163.367
R1796 B.n348 B.n118 163.367
R1797 B.n711 B.n408 163.367
R1798 B.n711 B.n406 163.367
R1799 B.n715 B.n406 163.367
R1800 B.n715 B.n400 163.367
R1801 B.n723 B.n400 163.367
R1802 B.n723 B.n398 163.367
R1803 B.n727 B.n398 163.367
R1804 B.n727 B.n392 163.367
R1805 B.n735 B.n392 163.367
R1806 B.n735 B.n390 163.367
R1807 B.n739 B.n390 163.367
R1808 B.n739 B.n384 163.367
R1809 B.n747 B.n384 163.367
R1810 B.n747 B.n382 163.367
R1811 B.n751 B.n382 163.367
R1812 B.n751 B.n375 163.367
R1813 B.n759 B.n375 163.367
R1814 B.n759 B.n373 163.367
R1815 B.n763 B.n373 163.367
R1816 B.n763 B.n368 163.367
R1817 B.n771 B.n368 163.367
R1818 B.n771 B.n366 163.367
R1819 B.n775 B.n366 163.367
R1820 B.n775 B.n360 163.367
R1821 B.n783 B.n360 163.367
R1822 B.n783 B.n358 163.367
R1823 B.n788 B.n358 163.367
R1824 B.n788 B.n352 163.367
R1825 B.n796 B.n352 163.367
R1826 B.n797 B.n796 163.367
R1827 B.n797 B.n5 163.367
R1828 B.n6 B.n5 163.367
R1829 B.n7 B.n6 163.367
R1830 B.n803 B.n7 163.367
R1831 B.n804 B.n803 163.367
R1832 B.n804 B.n13 163.367
R1833 B.n14 B.n13 163.367
R1834 B.n15 B.n14 163.367
R1835 B.n809 B.n15 163.367
R1836 B.n809 B.n20 163.367
R1837 B.n21 B.n20 163.367
R1838 B.n22 B.n21 163.367
R1839 B.n814 B.n22 163.367
R1840 B.n814 B.n27 163.367
R1841 B.n28 B.n27 163.367
R1842 B.n29 B.n28 163.367
R1843 B.n819 B.n29 163.367
R1844 B.n819 B.n34 163.367
R1845 B.n35 B.n34 163.367
R1846 B.n36 B.n35 163.367
R1847 B.n824 B.n36 163.367
R1848 B.n824 B.n41 163.367
R1849 B.n42 B.n41 163.367
R1850 B.n43 B.n42 163.367
R1851 B.n829 B.n43 163.367
R1852 B.n829 B.n48 163.367
R1853 B.n49 B.n48 163.367
R1854 B.n50 B.n49 163.367
R1855 B.n834 B.n50 163.367
R1856 B.n834 B.n55 163.367
R1857 B.n56 B.n55 163.367
R1858 B.n57 B.n56 163.367
R1859 B.n119 B.n57 163.367
R1860 B.n702 B.n412 163.367
R1861 B.n702 B.n470 163.367
R1862 B.n698 B.n697 163.367
R1863 B.n694 B.n693 163.367
R1864 B.n690 B.n689 163.367
R1865 B.n686 B.n685 163.367
R1866 B.n682 B.n681 163.367
R1867 B.n678 B.n677 163.367
R1868 B.n674 B.n673 163.367
R1869 B.n670 B.n669 163.367
R1870 B.n666 B.n665 163.367
R1871 B.n662 B.n661 163.367
R1872 B.n658 B.n657 163.367
R1873 B.n654 B.n653 163.367
R1874 B.n650 B.n649 163.367
R1875 B.n646 B.n645 163.367
R1876 B.n642 B.n641 163.367
R1877 B.n638 B.n637 163.367
R1878 B.n634 B.n633 163.367
R1879 B.n630 B.n629 163.367
R1880 B.n626 B.n625 163.367
R1881 B.n622 B.n621 163.367
R1882 B.n618 B.n617 163.367
R1883 B.n614 B.n613 163.367
R1884 B.n610 B.n609 163.367
R1885 B.n606 B.n605 163.367
R1886 B.n602 B.n601 163.367
R1887 B.n598 B.n597 163.367
R1888 B.n594 B.n593 163.367
R1889 B.n590 B.n589 163.367
R1890 B.n586 B.n585 163.367
R1891 B.n582 B.n581 163.367
R1892 B.n578 B.n577 163.367
R1893 B.n574 B.n573 163.367
R1894 B.n570 B.n569 163.367
R1895 B.n566 B.n565 163.367
R1896 B.n562 B.n561 163.367
R1897 B.n558 B.n557 163.367
R1898 B.n554 B.n553 163.367
R1899 B.n550 B.n549 163.367
R1900 B.n546 B.n545 163.367
R1901 B.n542 B.n541 163.367
R1902 B.n538 B.n537 163.367
R1903 B.n534 B.n533 163.367
R1904 B.n530 B.n529 163.367
R1905 B.n526 B.n525 163.367
R1906 B.n522 B.n521 163.367
R1907 B.n518 B.n517 163.367
R1908 B.n514 B.n513 163.367
R1909 B.n510 B.n509 163.367
R1910 B.n506 B.n505 163.367
R1911 B.n502 B.n501 163.367
R1912 B.n498 B.n497 163.367
R1913 B.n494 B.n493 163.367
R1914 B.n490 B.n489 163.367
R1915 B.n486 B.n485 163.367
R1916 B.n482 B.n481 163.367
R1917 B.n478 B.n469 163.367
R1918 B.n709 B.n410 163.367
R1919 B.n709 B.n404 163.367
R1920 B.n717 B.n404 163.367
R1921 B.n717 B.n402 163.367
R1922 B.n721 B.n402 163.367
R1923 B.n721 B.n396 163.367
R1924 B.n729 B.n396 163.367
R1925 B.n729 B.n394 163.367
R1926 B.n733 B.n394 163.367
R1927 B.n733 B.n388 163.367
R1928 B.n741 B.n388 163.367
R1929 B.n741 B.n386 163.367
R1930 B.n745 B.n386 163.367
R1931 B.n745 B.n380 163.367
R1932 B.n753 B.n380 163.367
R1933 B.n753 B.n378 163.367
R1934 B.n757 B.n378 163.367
R1935 B.n757 B.n372 163.367
R1936 B.n765 B.n372 163.367
R1937 B.n765 B.n370 163.367
R1938 B.n769 B.n370 163.367
R1939 B.n769 B.n364 163.367
R1940 B.n777 B.n364 163.367
R1941 B.n777 B.n362 163.367
R1942 B.n781 B.n362 163.367
R1943 B.n781 B.n356 163.367
R1944 B.n790 B.n356 163.367
R1945 B.n790 B.n354 163.367
R1946 B.n794 B.n354 163.367
R1947 B.n794 B.n3 163.367
R1948 B.n910 B.n3 163.367
R1949 B.n906 B.n2 163.367
R1950 B.n906 B.n905 163.367
R1951 B.n905 B.n9 163.367
R1952 B.n901 B.n9 163.367
R1953 B.n901 B.n11 163.367
R1954 B.n897 B.n11 163.367
R1955 B.n897 B.n17 163.367
R1956 B.n893 B.n17 163.367
R1957 B.n893 B.n19 163.367
R1958 B.n889 B.n19 163.367
R1959 B.n889 B.n24 163.367
R1960 B.n885 B.n24 163.367
R1961 B.n885 B.n26 163.367
R1962 B.n881 B.n26 163.367
R1963 B.n881 B.n31 163.367
R1964 B.n877 B.n31 163.367
R1965 B.n877 B.n33 163.367
R1966 B.n873 B.n33 163.367
R1967 B.n873 B.n38 163.367
R1968 B.n869 B.n38 163.367
R1969 B.n869 B.n40 163.367
R1970 B.n865 B.n40 163.367
R1971 B.n865 B.n45 163.367
R1972 B.n861 B.n45 163.367
R1973 B.n861 B.n47 163.367
R1974 B.n857 B.n47 163.367
R1975 B.n857 B.n52 163.367
R1976 B.n853 B.n52 163.367
R1977 B.n853 B.n54 163.367
R1978 B.n849 B.n54 163.367
R1979 B.n849 B.n59 163.367
R1980 B.n845 B.n844 71.676
R1981 B.n124 B.n62 71.676
R1982 B.n128 B.n63 71.676
R1983 B.n132 B.n64 71.676
R1984 B.n136 B.n65 71.676
R1985 B.n140 B.n66 71.676
R1986 B.n144 B.n67 71.676
R1987 B.n148 B.n68 71.676
R1988 B.n152 B.n69 71.676
R1989 B.n156 B.n70 71.676
R1990 B.n160 B.n71 71.676
R1991 B.n164 B.n72 71.676
R1992 B.n168 B.n73 71.676
R1993 B.n172 B.n74 71.676
R1994 B.n176 B.n75 71.676
R1995 B.n180 B.n76 71.676
R1996 B.n184 B.n77 71.676
R1997 B.n188 B.n78 71.676
R1998 B.n192 B.n79 71.676
R1999 B.n196 B.n80 71.676
R2000 B.n200 B.n81 71.676
R2001 B.n204 B.n82 71.676
R2002 B.n208 B.n83 71.676
R2003 B.n212 B.n84 71.676
R2004 B.n216 B.n85 71.676
R2005 B.n220 B.n86 71.676
R2006 B.n224 B.n87 71.676
R2007 B.n229 B.n88 71.676
R2008 B.n233 B.n89 71.676
R2009 B.n237 B.n90 71.676
R2010 B.n241 B.n91 71.676
R2011 B.n245 B.n92 71.676
R2012 B.n250 B.n93 71.676
R2013 B.n254 B.n94 71.676
R2014 B.n258 B.n95 71.676
R2015 B.n262 B.n96 71.676
R2016 B.n266 B.n97 71.676
R2017 B.n270 B.n98 71.676
R2018 B.n274 B.n99 71.676
R2019 B.n278 B.n100 71.676
R2020 B.n282 B.n101 71.676
R2021 B.n286 B.n102 71.676
R2022 B.n290 B.n103 71.676
R2023 B.n294 B.n104 71.676
R2024 B.n298 B.n105 71.676
R2025 B.n302 B.n106 71.676
R2026 B.n306 B.n107 71.676
R2027 B.n310 B.n108 71.676
R2028 B.n314 B.n109 71.676
R2029 B.n318 B.n110 71.676
R2030 B.n322 B.n111 71.676
R2031 B.n326 B.n112 71.676
R2032 B.n330 B.n113 71.676
R2033 B.n334 B.n114 71.676
R2034 B.n338 B.n115 71.676
R2035 B.n342 B.n116 71.676
R2036 B.n346 B.n117 71.676
R2037 B.n842 B.n118 71.676
R2038 B.n842 B.n841 71.676
R2039 B.n348 B.n117 71.676
R2040 B.n345 B.n116 71.676
R2041 B.n341 B.n115 71.676
R2042 B.n337 B.n114 71.676
R2043 B.n333 B.n113 71.676
R2044 B.n329 B.n112 71.676
R2045 B.n325 B.n111 71.676
R2046 B.n321 B.n110 71.676
R2047 B.n317 B.n109 71.676
R2048 B.n313 B.n108 71.676
R2049 B.n309 B.n107 71.676
R2050 B.n305 B.n106 71.676
R2051 B.n301 B.n105 71.676
R2052 B.n297 B.n104 71.676
R2053 B.n293 B.n103 71.676
R2054 B.n289 B.n102 71.676
R2055 B.n285 B.n101 71.676
R2056 B.n281 B.n100 71.676
R2057 B.n277 B.n99 71.676
R2058 B.n273 B.n98 71.676
R2059 B.n269 B.n97 71.676
R2060 B.n265 B.n96 71.676
R2061 B.n261 B.n95 71.676
R2062 B.n257 B.n94 71.676
R2063 B.n253 B.n93 71.676
R2064 B.n249 B.n92 71.676
R2065 B.n244 B.n91 71.676
R2066 B.n240 B.n90 71.676
R2067 B.n236 B.n89 71.676
R2068 B.n232 B.n88 71.676
R2069 B.n228 B.n87 71.676
R2070 B.n223 B.n86 71.676
R2071 B.n219 B.n85 71.676
R2072 B.n215 B.n84 71.676
R2073 B.n211 B.n83 71.676
R2074 B.n207 B.n82 71.676
R2075 B.n203 B.n81 71.676
R2076 B.n199 B.n80 71.676
R2077 B.n195 B.n79 71.676
R2078 B.n191 B.n78 71.676
R2079 B.n187 B.n77 71.676
R2080 B.n183 B.n76 71.676
R2081 B.n179 B.n75 71.676
R2082 B.n175 B.n74 71.676
R2083 B.n171 B.n73 71.676
R2084 B.n167 B.n72 71.676
R2085 B.n163 B.n71 71.676
R2086 B.n159 B.n70 71.676
R2087 B.n155 B.n69 71.676
R2088 B.n151 B.n68 71.676
R2089 B.n147 B.n67 71.676
R2090 B.n143 B.n66 71.676
R2091 B.n139 B.n65 71.676
R2092 B.n135 B.n64 71.676
R2093 B.n131 B.n63 71.676
R2094 B.n127 B.n62 71.676
R2095 B.n844 B.n61 71.676
R2096 B.n705 B.n704 71.676
R2097 B.n470 B.n413 71.676
R2098 B.n697 B.n414 71.676
R2099 B.n693 B.n415 71.676
R2100 B.n689 B.n416 71.676
R2101 B.n685 B.n417 71.676
R2102 B.n681 B.n418 71.676
R2103 B.n677 B.n419 71.676
R2104 B.n673 B.n420 71.676
R2105 B.n669 B.n421 71.676
R2106 B.n665 B.n422 71.676
R2107 B.n661 B.n423 71.676
R2108 B.n657 B.n424 71.676
R2109 B.n653 B.n425 71.676
R2110 B.n649 B.n426 71.676
R2111 B.n645 B.n427 71.676
R2112 B.n641 B.n428 71.676
R2113 B.n637 B.n429 71.676
R2114 B.n633 B.n430 71.676
R2115 B.n629 B.n431 71.676
R2116 B.n625 B.n432 71.676
R2117 B.n621 B.n433 71.676
R2118 B.n617 B.n434 71.676
R2119 B.n613 B.n435 71.676
R2120 B.n609 B.n436 71.676
R2121 B.n605 B.n437 71.676
R2122 B.n601 B.n438 71.676
R2123 B.n597 B.n439 71.676
R2124 B.n593 B.n440 71.676
R2125 B.n589 B.n441 71.676
R2126 B.n585 B.n442 71.676
R2127 B.n581 B.n443 71.676
R2128 B.n577 B.n444 71.676
R2129 B.n573 B.n445 71.676
R2130 B.n569 B.n446 71.676
R2131 B.n565 B.n447 71.676
R2132 B.n561 B.n448 71.676
R2133 B.n557 B.n449 71.676
R2134 B.n553 B.n450 71.676
R2135 B.n549 B.n451 71.676
R2136 B.n545 B.n452 71.676
R2137 B.n541 B.n453 71.676
R2138 B.n537 B.n454 71.676
R2139 B.n533 B.n455 71.676
R2140 B.n529 B.n456 71.676
R2141 B.n525 B.n457 71.676
R2142 B.n521 B.n458 71.676
R2143 B.n517 B.n459 71.676
R2144 B.n513 B.n460 71.676
R2145 B.n509 B.n461 71.676
R2146 B.n505 B.n462 71.676
R2147 B.n501 B.n463 71.676
R2148 B.n497 B.n464 71.676
R2149 B.n493 B.n465 71.676
R2150 B.n489 B.n466 71.676
R2151 B.n485 B.n467 71.676
R2152 B.n481 B.n468 71.676
R2153 B.n704 B.n412 71.676
R2154 B.n698 B.n413 71.676
R2155 B.n694 B.n414 71.676
R2156 B.n690 B.n415 71.676
R2157 B.n686 B.n416 71.676
R2158 B.n682 B.n417 71.676
R2159 B.n678 B.n418 71.676
R2160 B.n674 B.n419 71.676
R2161 B.n670 B.n420 71.676
R2162 B.n666 B.n421 71.676
R2163 B.n662 B.n422 71.676
R2164 B.n658 B.n423 71.676
R2165 B.n654 B.n424 71.676
R2166 B.n650 B.n425 71.676
R2167 B.n646 B.n426 71.676
R2168 B.n642 B.n427 71.676
R2169 B.n638 B.n428 71.676
R2170 B.n634 B.n429 71.676
R2171 B.n630 B.n430 71.676
R2172 B.n626 B.n431 71.676
R2173 B.n622 B.n432 71.676
R2174 B.n618 B.n433 71.676
R2175 B.n614 B.n434 71.676
R2176 B.n610 B.n435 71.676
R2177 B.n606 B.n436 71.676
R2178 B.n602 B.n437 71.676
R2179 B.n598 B.n438 71.676
R2180 B.n594 B.n439 71.676
R2181 B.n590 B.n440 71.676
R2182 B.n586 B.n441 71.676
R2183 B.n582 B.n442 71.676
R2184 B.n578 B.n443 71.676
R2185 B.n574 B.n444 71.676
R2186 B.n570 B.n445 71.676
R2187 B.n566 B.n446 71.676
R2188 B.n562 B.n447 71.676
R2189 B.n558 B.n448 71.676
R2190 B.n554 B.n449 71.676
R2191 B.n550 B.n450 71.676
R2192 B.n546 B.n451 71.676
R2193 B.n542 B.n452 71.676
R2194 B.n538 B.n453 71.676
R2195 B.n534 B.n454 71.676
R2196 B.n530 B.n455 71.676
R2197 B.n526 B.n456 71.676
R2198 B.n522 B.n457 71.676
R2199 B.n518 B.n458 71.676
R2200 B.n514 B.n459 71.676
R2201 B.n510 B.n460 71.676
R2202 B.n506 B.n461 71.676
R2203 B.n502 B.n462 71.676
R2204 B.n498 B.n463 71.676
R2205 B.n494 B.n464 71.676
R2206 B.n490 B.n465 71.676
R2207 B.n486 B.n466 71.676
R2208 B.n482 B.n467 71.676
R2209 B.n478 B.n468 71.676
R2210 B.n911 B.n910 71.676
R2211 B.n911 B.n2 71.676
R2212 B.n703 B.n409 66.7299
R2213 B.n843 B.n58 66.7299
R2214 B.n226 B.n123 59.5399
R2215 B.n247 B.n121 59.5399
R2216 B.n476 B.n475 59.5399
R2217 B.n473 B.n472 59.5399
R2218 B.n123 B.n122 51.5884
R2219 B.n121 B.n120 51.5884
R2220 B.n475 B.n474 51.5884
R2221 B.n472 B.n471 51.5884
R2222 B.n710 B.n409 35.1757
R2223 B.n710 B.n405 35.1757
R2224 B.n716 B.n405 35.1757
R2225 B.n716 B.n401 35.1757
R2226 B.n722 B.n401 35.1757
R2227 B.n722 B.n397 35.1757
R2228 B.n728 B.n397 35.1757
R2229 B.n734 B.n393 35.1757
R2230 B.n734 B.n389 35.1757
R2231 B.n740 B.n389 35.1757
R2232 B.n740 B.n385 35.1757
R2233 B.n746 B.n385 35.1757
R2234 B.n746 B.n381 35.1757
R2235 B.n752 B.n381 35.1757
R2236 B.n752 B.n376 35.1757
R2237 B.n758 B.n376 35.1757
R2238 B.n758 B.n377 35.1757
R2239 B.n764 B.n369 35.1757
R2240 B.n770 B.n369 35.1757
R2241 B.n770 B.n365 35.1757
R2242 B.n776 B.n365 35.1757
R2243 B.n776 B.n361 35.1757
R2244 B.n782 B.n361 35.1757
R2245 B.n789 B.n357 35.1757
R2246 B.n789 B.n353 35.1757
R2247 B.n795 B.n353 35.1757
R2248 B.n795 B.n4 35.1757
R2249 B.n909 B.n4 35.1757
R2250 B.n909 B.n908 35.1757
R2251 B.n908 B.n907 35.1757
R2252 B.n907 B.n8 35.1757
R2253 B.n12 B.n8 35.1757
R2254 B.n900 B.n12 35.1757
R2255 B.n900 B.n899 35.1757
R2256 B.n898 B.n16 35.1757
R2257 B.n892 B.n16 35.1757
R2258 B.n892 B.n891 35.1757
R2259 B.n891 B.n890 35.1757
R2260 B.n890 B.n23 35.1757
R2261 B.n884 B.n23 35.1757
R2262 B.n883 B.n882 35.1757
R2263 B.n882 B.n30 35.1757
R2264 B.n876 B.n30 35.1757
R2265 B.n876 B.n875 35.1757
R2266 B.n875 B.n874 35.1757
R2267 B.n874 B.n37 35.1757
R2268 B.n868 B.n37 35.1757
R2269 B.n868 B.n867 35.1757
R2270 B.n867 B.n866 35.1757
R2271 B.n866 B.n44 35.1757
R2272 B.n860 B.n859 35.1757
R2273 B.n859 B.n858 35.1757
R2274 B.n858 B.n51 35.1757
R2275 B.n852 B.n51 35.1757
R2276 B.n852 B.n851 35.1757
R2277 B.n851 B.n850 35.1757
R2278 B.n850 B.n58 35.1757
R2279 B.n707 B.n706 34.8103
R2280 B.n477 B.n407 34.8103
R2281 B.n847 B.n846 34.8103
R2282 B.n840 B.n839 34.8103
R2283 B.n782 B.t3 34.6584
R2284 B.t0 B.n898 34.6584
R2285 B.t9 B.n393 30.5201
R2286 B.t5 B.n44 30.5201
R2287 B.n764 B.t2 29.4856
R2288 B.n884 B.t1 29.4856
R2289 B B.n912 18.0485
R2290 B.n708 B.n707 10.6151
R2291 B.n708 B.n403 10.6151
R2292 B.n718 B.n403 10.6151
R2293 B.n719 B.n718 10.6151
R2294 B.n720 B.n719 10.6151
R2295 B.n720 B.n395 10.6151
R2296 B.n730 B.n395 10.6151
R2297 B.n731 B.n730 10.6151
R2298 B.n732 B.n731 10.6151
R2299 B.n732 B.n387 10.6151
R2300 B.n742 B.n387 10.6151
R2301 B.n743 B.n742 10.6151
R2302 B.n744 B.n743 10.6151
R2303 B.n744 B.n379 10.6151
R2304 B.n754 B.n379 10.6151
R2305 B.n755 B.n754 10.6151
R2306 B.n756 B.n755 10.6151
R2307 B.n756 B.n371 10.6151
R2308 B.n766 B.n371 10.6151
R2309 B.n767 B.n766 10.6151
R2310 B.n768 B.n767 10.6151
R2311 B.n768 B.n363 10.6151
R2312 B.n778 B.n363 10.6151
R2313 B.n779 B.n778 10.6151
R2314 B.n780 B.n779 10.6151
R2315 B.n780 B.n355 10.6151
R2316 B.n791 B.n355 10.6151
R2317 B.n792 B.n791 10.6151
R2318 B.n793 B.n792 10.6151
R2319 B.n793 B.n0 10.6151
R2320 B.n706 B.n411 10.6151
R2321 B.n701 B.n411 10.6151
R2322 B.n701 B.n700 10.6151
R2323 B.n700 B.n699 10.6151
R2324 B.n699 B.n696 10.6151
R2325 B.n696 B.n695 10.6151
R2326 B.n695 B.n692 10.6151
R2327 B.n692 B.n691 10.6151
R2328 B.n691 B.n688 10.6151
R2329 B.n688 B.n687 10.6151
R2330 B.n687 B.n684 10.6151
R2331 B.n684 B.n683 10.6151
R2332 B.n683 B.n680 10.6151
R2333 B.n680 B.n679 10.6151
R2334 B.n679 B.n676 10.6151
R2335 B.n676 B.n675 10.6151
R2336 B.n675 B.n672 10.6151
R2337 B.n672 B.n671 10.6151
R2338 B.n671 B.n668 10.6151
R2339 B.n668 B.n667 10.6151
R2340 B.n667 B.n664 10.6151
R2341 B.n664 B.n663 10.6151
R2342 B.n663 B.n660 10.6151
R2343 B.n660 B.n659 10.6151
R2344 B.n659 B.n656 10.6151
R2345 B.n656 B.n655 10.6151
R2346 B.n655 B.n652 10.6151
R2347 B.n652 B.n651 10.6151
R2348 B.n651 B.n648 10.6151
R2349 B.n648 B.n647 10.6151
R2350 B.n647 B.n644 10.6151
R2351 B.n644 B.n643 10.6151
R2352 B.n643 B.n640 10.6151
R2353 B.n640 B.n639 10.6151
R2354 B.n639 B.n636 10.6151
R2355 B.n636 B.n635 10.6151
R2356 B.n635 B.n632 10.6151
R2357 B.n632 B.n631 10.6151
R2358 B.n631 B.n628 10.6151
R2359 B.n628 B.n627 10.6151
R2360 B.n627 B.n624 10.6151
R2361 B.n624 B.n623 10.6151
R2362 B.n623 B.n620 10.6151
R2363 B.n620 B.n619 10.6151
R2364 B.n619 B.n616 10.6151
R2365 B.n616 B.n615 10.6151
R2366 B.n615 B.n612 10.6151
R2367 B.n612 B.n611 10.6151
R2368 B.n611 B.n608 10.6151
R2369 B.n608 B.n607 10.6151
R2370 B.n607 B.n604 10.6151
R2371 B.n604 B.n603 10.6151
R2372 B.n600 B.n599 10.6151
R2373 B.n599 B.n596 10.6151
R2374 B.n596 B.n595 10.6151
R2375 B.n595 B.n592 10.6151
R2376 B.n592 B.n591 10.6151
R2377 B.n591 B.n588 10.6151
R2378 B.n588 B.n587 10.6151
R2379 B.n587 B.n584 10.6151
R2380 B.n584 B.n583 10.6151
R2381 B.n580 B.n579 10.6151
R2382 B.n579 B.n576 10.6151
R2383 B.n576 B.n575 10.6151
R2384 B.n575 B.n572 10.6151
R2385 B.n572 B.n571 10.6151
R2386 B.n571 B.n568 10.6151
R2387 B.n568 B.n567 10.6151
R2388 B.n567 B.n564 10.6151
R2389 B.n564 B.n563 10.6151
R2390 B.n563 B.n560 10.6151
R2391 B.n560 B.n559 10.6151
R2392 B.n559 B.n556 10.6151
R2393 B.n556 B.n555 10.6151
R2394 B.n555 B.n552 10.6151
R2395 B.n552 B.n551 10.6151
R2396 B.n551 B.n548 10.6151
R2397 B.n548 B.n547 10.6151
R2398 B.n547 B.n544 10.6151
R2399 B.n544 B.n543 10.6151
R2400 B.n543 B.n540 10.6151
R2401 B.n540 B.n539 10.6151
R2402 B.n539 B.n536 10.6151
R2403 B.n536 B.n535 10.6151
R2404 B.n535 B.n532 10.6151
R2405 B.n532 B.n531 10.6151
R2406 B.n531 B.n528 10.6151
R2407 B.n528 B.n527 10.6151
R2408 B.n527 B.n524 10.6151
R2409 B.n524 B.n523 10.6151
R2410 B.n523 B.n520 10.6151
R2411 B.n520 B.n519 10.6151
R2412 B.n519 B.n516 10.6151
R2413 B.n516 B.n515 10.6151
R2414 B.n515 B.n512 10.6151
R2415 B.n512 B.n511 10.6151
R2416 B.n511 B.n508 10.6151
R2417 B.n508 B.n507 10.6151
R2418 B.n507 B.n504 10.6151
R2419 B.n504 B.n503 10.6151
R2420 B.n503 B.n500 10.6151
R2421 B.n500 B.n499 10.6151
R2422 B.n499 B.n496 10.6151
R2423 B.n496 B.n495 10.6151
R2424 B.n495 B.n492 10.6151
R2425 B.n492 B.n491 10.6151
R2426 B.n491 B.n488 10.6151
R2427 B.n488 B.n487 10.6151
R2428 B.n487 B.n484 10.6151
R2429 B.n484 B.n483 10.6151
R2430 B.n483 B.n480 10.6151
R2431 B.n480 B.n479 10.6151
R2432 B.n479 B.n477 10.6151
R2433 B.n712 B.n407 10.6151
R2434 B.n713 B.n712 10.6151
R2435 B.n714 B.n713 10.6151
R2436 B.n714 B.n399 10.6151
R2437 B.n724 B.n399 10.6151
R2438 B.n725 B.n724 10.6151
R2439 B.n726 B.n725 10.6151
R2440 B.n726 B.n391 10.6151
R2441 B.n736 B.n391 10.6151
R2442 B.n737 B.n736 10.6151
R2443 B.n738 B.n737 10.6151
R2444 B.n738 B.n383 10.6151
R2445 B.n748 B.n383 10.6151
R2446 B.n749 B.n748 10.6151
R2447 B.n750 B.n749 10.6151
R2448 B.n750 B.n374 10.6151
R2449 B.n760 B.n374 10.6151
R2450 B.n761 B.n760 10.6151
R2451 B.n762 B.n761 10.6151
R2452 B.n762 B.n367 10.6151
R2453 B.n772 B.n367 10.6151
R2454 B.n773 B.n772 10.6151
R2455 B.n774 B.n773 10.6151
R2456 B.n774 B.n359 10.6151
R2457 B.n784 B.n359 10.6151
R2458 B.n785 B.n784 10.6151
R2459 B.n787 B.n785 10.6151
R2460 B.n787 B.n786 10.6151
R2461 B.n786 B.n351 10.6151
R2462 B.n798 B.n351 10.6151
R2463 B.n799 B.n798 10.6151
R2464 B.n800 B.n799 10.6151
R2465 B.n801 B.n800 10.6151
R2466 B.n802 B.n801 10.6151
R2467 B.n805 B.n802 10.6151
R2468 B.n806 B.n805 10.6151
R2469 B.n807 B.n806 10.6151
R2470 B.n808 B.n807 10.6151
R2471 B.n810 B.n808 10.6151
R2472 B.n811 B.n810 10.6151
R2473 B.n812 B.n811 10.6151
R2474 B.n813 B.n812 10.6151
R2475 B.n815 B.n813 10.6151
R2476 B.n816 B.n815 10.6151
R2477 B.n817 B.n816 10.6151
R2478 B.n818 B.n817 10.6151
R2479 B.n820 B.n818 10.6151
R2480 B.n821 B.n820 10.6151
R2481 B.n822 B.n821 10.6151
R2482 B.n823 B.n822 10.6151
R2483 B.n825 B.n823 10.6151
R2484 B.n826 B.n825 10.6151
R2485 B.n827 B.n826 10.6151
R2486 B.n828 B.n827 10.6151
R2487 B.n830 B.n828 10.6151
R2488 B.n831 B.n830 10.6151
R2489 B.n832 B.n831 10.6151
R2490 B.n833 B.n832 10.6151
R2491 B.n835 B.n833 10.6151
R2492 B.n836 B.n835 10.6151
R2493 B.n837 B.n836 10.6151
R2494 B.n838 B.n837 10.6151
R2495 B.n839 B.n838 10.6151
R2496 B.n904 B.n1 10.6151
R2497 B.n904 B.n903 10.6151
R2498 B.n903 B.n902 10.6151
R2499 B.n902 B.n10 10.6151
R2500 B.n896 B.n10 10.6151
R2501 B.n896 B.n895 10.6151
R2502 B.n895 B.n894 10.6151
R2503 B.n894 B.n18 10.6151
R2504 B.n888 B.n18 10.6151
R2505 B.n888 B.n887 10.6151
R2506 B.n887 B.n886 10.6151
R2507 B.n886 B.n25 10.6151
R2508 B.n880 B.n25 10.6151
R2509 B.n880 B.n879 10.6151
R2510 B.n879 B.n878 10.6151
R2511 B.n878 B.n32 10.6151
R2512 B.n872 B.n32 10.6151
R2513 B.n872 B.n871 10.6151
R2514 B.n871 B.n870 10.6151
R2515 B.n870 B.n39 10.6151
R2516 B.n864 B.n39 10.6151
R2517 B.n864 B.n863 10.6151
R2518 B.n863 B.n862 10.6151
R2519 B.n862 B.n46 10.6151
R2520 B.n856 B.n46 10.6151
R2521 B.n856 B.n855 10.6151
R2522 B.n855 B.n854 10.6151
R2523 B.n854 B.n53 10.6151
R2524 B.n848 B.n53 10.6151
R2525 B.n848 B.n847 10.6151
R2526 B.n846 B.n60 10.6151
R2527 B.n125 B.n60 10.6151
R2528 B.n126 B.n125 10.6151
R2529 B.n129 B.n126 10.6151
R2530 B.n130 B.n129 10.6151
R2531 B.n133 B.n130 10.6151
R2532 B.n134 B.n133 10.6151
R2533 B.n137 B.n134 10.6151
R2534 B.n138 B.n137 10.6151
R2535 B.n141 B.n138 10.6151
R2536 B.n142 B.n141 10.6151
R2537 B.n145 B.n142 10.6151
R2538 B.n146 B.n145 10.6151
R2539 B.n149 B.n146 10.6151
R2540 B.n150 B.n149 10.6151
R2541 B.n153 B.n150 10.6151
R2542 B.n154 B.n153 10.6151
R2543 B.n157 B.n154 10.6151
R2544 B.n158 B.n157 10.6151
R2545 B.n161 B.n158 10.6151
R2546 B.n162 B.n161 10.6151
R2547 B.n165 B.n162 10.6151
R2548 B.n166 B.n165 10.6151
R2549 B.n169 B.n166 10.6151
R2550 B.n170 B.n169 10.6151
R2551 B.n173 B.n170 10.6151
R2552 B.n174 B.n173 10.6151
R2553 B.n177 B.n174 10.6151
R2554 B.n178 B.n177 10.6151
R2555 B.n181 B.n178 10.6151
R2556 B.n182 B.n181 10.6151
R2557 B.n185 B.n182 10.6151
R2558 B.n186 B.n185 10.6151
R2559 B.n189 B.n186 10.6151
R2560 B.n190 B.n189 10.6151
R2561 B.n193 B.n190 10.6151
R2562 B.n194 B.n193 10.6151
R2563 B.n197 B.n194 10.6151
R2564 B.n198 B.n197 10.6151
R2565 B.n201 B.n198 10.6151
R2566 B.n202 B.n201 10.6151
R2567 B.n205 B.n202 10.6151
R2568 B.n206 B.n205 10.6151
R2569 B.n209 B.n206 10.6151
R2570 B.n210 B.n209 10.6151
R2571 B.n213 B.n210 10.6151
R2572 B.n214 B.n213 10.6151
R2573 B.n217 B.n214 10.6151
R2574 B.n218 B.n217 10.6151
R2575 B.n221 B.n218 10.6151
R2576 B.n222 B.n221 10.6151
R2577 B.n225 B.n222 10.6151
R2578 B.n230 B.n227 10.6151
R2579 B.n231 B.n230 10.6151
R2580 B.n234 B.n231 10.6151
R2581 B.n235 B.n234 10.6151
R2582 B.n238 B.n235 10.6151
R2583 B.n239 B.n238 10.6151
R2584 B.n242 B.n239 10.6151
R2585 B.n243 B.n242 10.6151
R2586 B.n246 B.n243 10.6151
R2587 B.n251 B.n248 10.6151
R2588 B.n252 B.n251 10.6151
R2589 B.n255 B.n252 10.6151
R2590 B.n256 B.n255 10.6151
R2591 B.n259 B.n256 10.6151
R2592 B.n260 B.n259 10.6151
R2593 B.n263 B.n260 10.6151
R2594 B.n264 B.n263 10.6151
R2595 B.n267 B.n264 10.6151
R2596 B.n268 B.n267 10.6151
R2597 B.n271 B.n268 10.6151
R2598 B.n272 B.n271 10.6151
R2599 B.n275 B.n272 10.6151
R2600 B.n276 B.n275 10.6151
R2601 B.n279 B.n276 10.6151
R2602 B.n280 B.n279 10.6151
R2603 B.n283 B.n280 10.6151
R2604 B.n284 B.n283 10.6151
R2605 B.n287 B.n284 10.6151
R2606 B.n288 B.n287 10.6151
R2607 B.n291 B.n288 10.6151
R2608 B.n292 B.n291 10.6151
R2609 B.n295 B.n292 10.6151
R2610 B.n296 B.n295 10.6151
R2611 B.n299 B.n296 10.6151
R2612 B.n300 B.n299 10.6151
R2613 B.n303 B.n300 10.6151
R2614 B.n304 B.n303 10.6151
R2615 B.n307 B.n304 10.6151
R2616 B.n308 B.n307 10.6151
R2617 B.n311 B.n308 10.6151
R2618 B.n312 B.n311 10.6151
R2619 B.n315 B.n312 10.6151
R2620 B.n316 B.n315 10.6151
R2621 B.n319 B.n316 10.6151
R2622 B.n320 B.n319 10.6151
R2623 B.n323 B.n320 10.6151
R2624 B.n324 B.n323 10.6151
R2625 B.n327 B.n324 10.6151
R2626 B.n328 B.n327 10.6151
R2627 B.n331 B.n328 10.6151
R2628 B.n332 B.n331 10.6151
R2629 B.n335 B.n332 10.6151
R2630 B.n336 B.n335 10.6151
R2631 B.n339 B.n336 10.6151
R2632 B.n340 B.n339 10.6151
R2633 B.n343 B.n340 10.6151
R2634 B.n344 B.n343 10.6151
R2635 B.n347 B.n344 10.6151
R2636 B.n349 B.n347 10.6151
R2637 B.n350 B.n349 10.6151
R2638 B.n840 B.n350 10.6151
R2639 B.n603 B.n473 9.52245
R2640 B.n580 B.n476 9.52245
R2641 B.n226 B.n225 9.52245
R2642 B.n248 B.n247 9.52245
R2643 B.n912 B.n0 8.11757
R2644 B.n912 B.n1 8.11757
R2645 B.n377 B.t2 5.6906
R2646 B.t1 B.n883 5.6906
R2647 B.n728 B.t9 4.65604
R2648 B.n860 B.t5 4.65604
R2649 B.n600 B.n473 1.09318
R2650 B.n583 B.n476 1.09318
R2651 B.n227 B.n226 1.09318
R2652 B.n247 B.n246 1.09318
R2653 B.t3 B.n357 0.517782
R2654 B.n899 B.t0 0.517782
R2655 VN.n0 VN.t2 201.917
R2656 VN.n1 VN.t0 201.917
R2657 VN.n0 VN.t3 201.258
R2658 VN.n1 VN.t1 201.258
R2659 VN VN.n1 54.2866
R2660 VN VN.n0 5.4874
R2661 VDD2.n2 VDD2.n0 103.41
R2662 VDD2.n2 VDD2.n1 59.0321
R2663 VDD2.n1 VDD2.t2 1.23877
R2664 VDD2.n1 VDD2.t3 1.23877
R2665 VDD2.n0 VDD2.t1 1.23877
R2666 VDD2.n0 VDD2.t0 1.23877
R2667 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 6.1022f
C1 VDD2 VTAIL 6.41999f
C2 VN VTAIL 5.79853f
C3 VDD1 VP 6.3299f
C4 VDD2 VP 0.376965f
C5 VP VN 6.73422f
C6 VP VTAIL 5.81264f
C7 VDD1 VDD2 0.964595f
C8 VDD1 VN 0.148593f
C9 VDD1 VTAIL 6.367589f
C10 VDD2 B 3.914462f
C11 VDD1 B 8.35315f
C12 VTAIL B 12.30466f
C13 VN B 10.546339f
C14 VP B 8.641189f
C15 VDD2.t1 B 0.334968f
C16 VDD2.t0 B 0.334968f
C17 VDD2.n0 B 3.85078f
C18 VDD2.t2 B 0.334968f
C19 VDD2.t3 B 0.334968f
C20 VDD2.n1 B 3.03398f
C21 VDD2.n2 B 4.07379f
C22 VN.t2 B 2.89115f
C23 VN.t3 B 2.88762f
C24 VN.n0 B 1.88972f
C25 VN.t0 B 2.89115f
C26 VN.t1 B 2.88762f
C27 VN.n1 B 3.34761f
C28 VTAIL.n0 B 0.019596f
C29 VTAIL.n1 B 0.015504f
C30 VTAIL.n2 B 0.008331f
C31 VTAIL.n3 B 0.019692f
C32 VTAIL.n4 B 0.008821f
C33 VTAIL.n5 B 0.015504f
C34 VTAIL.n6 B 0.008576f
C35 VTAIL.n7 B 0.019692f
C36 VTAIL.n8 B 0.008821f
C37 VTAIL.n9 B 0.015504f
C38 VTAIL.n10 B 0.008331f
C39 VTAIL.n11 B 0.019692f
C40 VTAIL.n12 B 0.008821f
C41 VTAIL.n13 B 0.015504f
C42 VTAIL.n14 B 0.008331f
C43 VTAIL.n15 B 0.019692f
C44 VTAIL.n16 B 0.008821f
C45 VTAIL.n17 B 0.015504f
C46 VTAIL.n18 B 0.008331f
C47 VTAIL.n19 B 0.019692f
C48 VTAIL.n20 B 0.008821f
C49 VTAIL.n21 B 0.015504f
C50 VTAIL.n22 B 0.008331f
C51 VTAIL.n23 B 0.019692f
C52 VTAIL.n24 B 0.008821f
C53 VTAIL.n25 B 0.015504f
C54 VTAIL.n26 B 0.008331f
C55 VTAIL.n27 B 0.014769f
C56 VTAIL.n28 B 0.011633f
C57 VTAIL.t0 B 0.032523f
C58 VTAIL.n29 B 0.104971f
C59 VTAIL.n30 B 1.07908f
C60 VTAIL.n31 B 0.008331f
C61 VTAIL.n32 B 0.008821f
C62 VTAIL.n33 B 0.019692f
C63 VTAIL.n34 B 0.019692f
C64 VTAIL.n35 B 0.008821f
C65 VTAIL.n36 B 0.008331f
C66 VTAIL.n37 B 0.015504f
C67 VTAIL.n38 B 0.015504f
C68 VTAIL.n39 B 0.008331f
C69 VTAIL.n40 B 0.008821f
C70 VTAIL.n41 B 0.019692f
C71 VTAIL.n42 B 0.019692f
C72 VTAIL.n43 B 0.008821f
C73 VTAIL.n44 B 0.008331f
C74 VTAIL.n45 B 0.015504f
C75 VTAIL.n46 B 0.015504f
C76 VTAIL.n47 B 0.008331f
C77 VTAIL.n48 B 0.008821f
C78 VTAIL.n49 B 0.019692f
C79 VTAIL.n50 B 0.019692f
C80 VTAIL.n51 B 0.008821f
C81 VTAIL.n52 B 0.008331f
C82 VTAIL.n53 B 0.015504f
C83 VTAIL.n54 B 0.015504f
C84 VTAIL.n55 B 0.008331f
C85 VTAIL.n56 B 0.008821f
C86 VTAIL.n57 B 0.019692f
C87 VTAIL.n58 B 0.019692f
C88 VTAIL.n59 B 0.008821f
C89 VTAIL.n60 B 0.008331f
C90 VTAIL.n61 B 0.015504f
C91 VTAIL.n62 B 0.015504f
C92 VTAIL.n63 B 0.008331f
C93 VTAIL.n64 B 0.008821f
C94 VTAIL.n65 B 0.019692f
C95 VTAIL.n66 B 0.019692f
C96 VTAIL.n67 B 0.008821f
C97 VTAIL.n68 B 0.008331f
C98 VTAIL.n69 B 0.015504f
C99 VTAIL.n70 B 0.015504f
C100 VTAIL.n71 B 0.008331f
C101 VTAIL.n72 B 0.008331f
C102 VTAIL.n73 B 0.008821f
C103 VTAIL.n74 B 0.019692f
C104 VTAIL.n75 B 0.019692f
C105 VTAIL.n76 B 0.019692f
C106 VTAIL.n77 B 0.008576f
C107 VTAIL.n78 B 0.008331f
C108 VTAIL.n79 B 0.015504f
C109 VTAIL.n80 B 0.015504f
C110 VTAIL.n81 B 0.008331f
C111 VTAIL.n82 B 0.008821f
C112 VTAIL.n83 B 0.019692f
C113 VTAIL.n84 B 0.038746f
C114 VTAIL.n85 B 0.008821f
C115 VTAIL.n86 B 0.008331f
C116 VTAIL.n87 B 0.033931f
C117 VTAIL.n88 B 0.021221f
C118 VTAIL.n89 B 0.095827f
C119 VTAIL.n90 B 0.019596f
C120 VTAIL.n91 B 0.015504f
C121 VTAIL.n92 B 0.008331f
C122 VTAIL.n93 B 0.019692f
C123 VTAIL.n94 B 0.008821f
C124 VTAIL.n95 B 0.015504f
C125 VTAIL.n96 B 0.008576f
C126 VTAIL.n97 B 0.019692f
C127 VTAIL.n98 B 0.008821f
C128 VTAIL.n99 B 0.015504f
C129 VTAIL.n100 B 0.008331f
C130 VTAIL.n101 B 0.019692f
C131 VTAIL.n102 B 0.008821f
C132 VTAIL.n103 B 0.015504f
C133 VTAIL.n104 B 0.008331f
C134 VTAIL.n105 B 0.019692f
C135 VTAIL.n106 B 0.008821f
C136 VTAIL.n107 B 0.015504f
C137 VTAIL.n108 B 0.008331f
C138 VTAIL.n109 B 0.019692f
C139 VTAIL.n110 B 0.008821f
C140 VTAIL.n111 B 0.015504f
C141 VTAIL.n112 B 0.008331f
C142 VTAIL.n113 B 0.019692f
C143 VTAIL.n114 B 0.008821f
C144 VTAIL.n115 B 0.015504f
C145 VTAIL.n116 B 0.008331f
C146 VTAIL.n117 B 0.014769f
C147 VTAIL.n118 B 0.011633f
C148 VTAIL.t5 B 0.032523f
C149 VTAIL.n119 B 0.104971f
C150 VTAIL.n120 B 1.07908f
C151 VTAIL.n121 B 0.008331f
C152 VTAIL.n122 B 0.008821f
C153 VTAIL.n123 B 0.019692f
C154 VTAIL.n124 B 0.019692f
C155 VTAIL.n125 B 0.008821f
C156 VTAIL.n126 B 0.008331f
C157 VTAIL.n127 B 0.015504f
C158 VTAIL.n128 B 0.015504f
C159 VTAIL.n129 B 0.008331f
C160 VTAIL.n130 B 0.008821f
C161 VTAIL.n131 B 0.019692f
C162 VTAIL.n132 B 0.019692f
C163 VTAIL.n133 B 0.008821f
C164 VTAIL.n134 B 0.008331f
C165 VTAIL.n135 B 0.015504f
C166 VTAIL.n136 B 0.015504f
C167 VTAIL.n137 B 0.008331f
C168 VTAIL.n138 B 0.008821f
C169 VTAIL.n139 B 0.019692f
C170 VTAIL.n140 B 0.019692f
C171 VTAIL.n141 B 0.008821f
C172 VTAIL.n142 B 0.008331f
C173 VTAIL.n143 B 0.015504f
C174 VTAIL.n144 B 0.015504f
C175 VTAIL.n145 B 0.008331f
C176 VTAIL.n146 B 0.008821f
C177 VTAIL.n147 B 0.019692f
C178 VTAIL.n148 B 0.019692f
C179 VTAIL.n149 B 0.008821f
C180 VTAIL.n150 B 0.008331f
C181 VTAIL.n151 B 0.015504f
C182 VTAIL.n152 B 0.015504f
C183 VTAIL.n153 B 0.008331f
C184 VTAIL.n154 B 0.008821f
C185 VTAIL.n155 B 0.019692f
C186 VTAIL.n156 B 0.019692f
C187 VTAIL.n157 B 0.008821f
C188 VTAIL.n158 B 0.008331f
C189 VTAIL.n159 B 0.015504f
C190 VTAIL.n160 B 0.015504f
C191 VTAIL.n161 B 0.008331f
C192 VTAIL.n162 B 0.008331f
C193 VTAIL.n163 B 0.008821f
C194 VTAIL.n164 B 0.019692f
C195 VTAIL.n165 B 0.019692f
C196 VTAIL.n166 B 0.019692f
C197 VTAIL.n167 B 0.008576f
C198 VTAIL.n168 B 0.008331f
C199 VTAIL.n169 B 0.015504f
C200 VTAIL.n170 B 0.015504f
C201 VTAIL.n171 B 0.008331f
C202 VTAIL.n172 B 0.008821f
C203 VTAIL.n173 B 0.019692f
C204 VTAIL.n174 B 0.038746f
C205 VTAIL.n175 B 0.008821f
C206 VTAIL.n176 B 0.008331f
C207 VTAIL.n177 B 0.033931f
C208 VTAIL.n178 B 0.021221f
C209 VTAIL.n179 B 0.1502f
C210 VTAIL.n180 B 0.019596f
C211 VTAIL.n181 B 0.015504f
C212 VTAIL.n182 B 0.008331f
C213 VTAIL.n183 B 0.019692f
C214 VTAIL.n184 B 0.008821f
C215 VTAIL.n185 B 0.015504f
C216 VTAIL.n186 B 0.008576f
C217 VTAIL.n187 B 0.019692f
C218 VTAIL.n188 B 0.008821f
C219 VTAIL.n189 B 0.015504f
C220 VTAIL.n190 B 0.008331f
C221 VTAIL.n191 B 0.019692f
C222 VTAIL.n192 B 0.008821f
C223 VTAIL.n193 B 0.015504f
C224 VTAIL.n194 B 0.008331f
C225 VTAIL.n195 B 0.019692f
C226 VTAIL.n196 B 0.008821f
C227 VTAIL.n197 B 0.015504f
C228 VTAIL.n198 B 0.008331f
C229 VTAIL.n199 B 0.019692f
C230 VTAIL.n200 B 0.008821f
C231 VTAIL.n201 B 0.015504f
C232 VTAIL.n202 B 0.008331f
C233 VTAIL.n203 B 0.019692f
C234 VTAIL.n204 B 0.008821f
C235 VTAIL.n205 B 0.015504f
C236 VTAIL.n206 B 0.008331f
C237 VTAIL.n207 B 0.014769f
C238 VTAIL.n208 B 0.011633f
C239 VTAIL.t4 B 0.032523f
C240 VTAIL.n209 B 0.104971f
C241 VTAIL.n210 B 1.07908f
C242 VTAIL.n211 B 0.008331f
C243 VTAIL.n212 B 0.008821f
C244 VTAIL.n213 B 0.019692f
C245 VTAIL.n214 B 0.019692f
C246 VTAIL.n215 B 0.008821f
C247 VTAIL.n216 B 0.008331f
C248 VTAIL.n217 B 0.015504f
C249 VTAIL.n218 B 0.015504f
C250 VTAIL.n219 B 0.008331f
C251 VTAIL.n220 B 0.008821f
C252 VTAIL.n221 B 0.019692f
C253 VTAIL.n222 B 0.019692f
C254 VTAIL.n223 B 0.008821f
C255 VTAIL.n224 B 0.008331f
C256 VTAIL.n225 B 0.015504f
C257 VTAIL.n226 B 0.015504f
C258 VTAIL.n227 B 0.008331f
C259 VTAIL.n228 B 0.008821f
C260 VTAIL.n229 B 0.019692f
C261 VTAIL.n230 B 0.019692f
C262 VTAIL.n231 B 0.008821f
C263 VTAIL.n232 B 0.008331f
C264 VTAIL.n233 B 0.015504f
C265 VTAIL.n234 B 0.015504f
C266 VTAIL.n235 B 0.008331f
C267 VTAIL.n236 B 0.008821f
C268 VTAIL.n237 B 0.019692f
C269 VTAIL.n238 B 0.019692f
C270 VTAIL.n239 B 0.008821f
C271 VTAIL.n240 B 0.008331f
C272 VTAIL.n241 B 0.015504f
C273 VTAIL.n242 B 0.015504f
C274 VTAIL.n243 B 0.008331f
C275 VTAIL.n244 B 0.008821f
C276 VTAIL.n245 B 0.019692f
C277 VTAIL.n246 B 0.019692f
C278 VTAIL.n247 B 0.008821f
C279 VTAIL.n248 B 0.008331f
C280 VTAIL.n249 B 0.015504f
C281 VTAIL.n250 B 0.015504f
C282 VTAIL.n251 B 0.008331f
C283 VTAIL.n252 B 0.008331f
C284 VTAIL.n253 B 0.008821f
C285 VTAIL.n254 B 0.019692f
C286 VTAIL.n255 B 0.019692f
C287 VTAIL.n256 B 0.019692f
C288 VTAIL.n257 B 0.008576f
C289 VTAIL.n258 B 0.008331f
C290 VTAIL.n259 B 0.015504f
C291 VTAIL.n260 B 0.015504f
C292 VTAIL.n261 B 0.008331f
C293 VTAIL.n262 B 0.008821f
C294 VTAIL.n263 B 0.019692f
C295 VTAIL.n264 B 0.038746f
C296 VTAIL.n265 B 0.008821f
C297 VTAIL.n266 B 0.008331f
C298 VTAIL.n267 B 0.033931f
C299 VTAIL.n268 B 0.021221f
C300 VTAIL.n269 B 1.14055f
C301 VTAIL.n270 B 0.019596f
C302 VTAIL.n271 B 0.015504f
C303 VTAIL.n272 B 0.008331f
C304 VTAIL.n273 B 0.019692f
C305 VTAIL.n274 B 0.008821f
C306 VTAIL.n275 B 0.015504f
C307 VTAIL.n276 B 0.008576f
C308 VTAIL.n277 B 0.019692f
C309 VTAIL.n278 B 0.008331f
C310 VTAIL.n279 B 0.008821f
C311 VTAIL.n280 B 0.015504f
C312 VTAIL.n281 B 0.008331f
C313 VTAIL.n282 B 0.019692f
C314 VTAIL.n283 B 0.008821f
C315 VTAIL.n284 B 0.015504f
C316 VTAIL.n285 B 0.008331f
C317 VTAIL.n286 B 0.019692f
C318 VTAIL.n287 B 0.008821f
C319 VTAIL.n288 B 0.015504f
C320 VTAIL.n289 B 0.008331f
C321 VTAIL.n290 B 0.019692f
C322 VTAIL.n291 B 0.008821f
C323 VTAIL.n292 B 0.015504f
C324 VTAIL.n293 B 0.008331f
C325 VTAIL.n294 B 0.019692f
C326 VTAIL.n295 B 0.008821f
C327 VTAIL.n296 B 0.015504f
C328 VTAIL.n297 B 0.008331f
C329 VTAIL.n298 B 0.014769f
C330 VTAIL.n299 B 0.011633f
C331 VTAIL.t2 B 0.032523f
C332 VTAIL.n300 B 0.104971f
C333 VTAIL.n301 B 1.07908f
C334 VTAIL.n302 B 0.008331f
C335 VTAIL.n303 B 0.008821f
C336 VTAIL.n304 B 0.019692f
C337 VTAIL.n305 B 0.019692f
C338 VTAIL.n306 B 0.008821f
C339 VTAIL.n307 B 0.008331f
C340 VTAIL.n308 B 0.015504f
C341 VTAIL.n309 B 0.015504f
C342 VTAIL.n310 B 0.008331f
C343 VTAIL.n311 B 0.008821f
C344 VTAIL.n312 B 0.019692f
C345 VTAIL.n313 B 0.019692f
C346 VTAIL.n314 B 0.008821f
C347 VTAIL.n315 B 0.008331f
C348 VTAIL.n316 B 0.015504f
C349 VTAIL.n317 B 0.015504f
C350 VTAIL.n318 B 0.008331f
C351 VTAIL.n319 B 0.008821f
C352 VTAIL.n320 B 0.019692f
C353 VTAIL.n321 B 0.019692f
C354 VTAIL.n322 B 0.008821f
C355 VTAIL.n323 B 0.008331f
C356 VTAIL.n324 B 0.015504f
C357 VTAIL.n325 B 0.015504f
C358 VTAIL.n326 B 0.008331f
C359 VTAIL.n327 B 0.008821f
C360 VTAIL.n328 B 0.019692f
C361 VTAIL.n329 B 0.019692f
C362 VTAIL.n330 B 0.008821f
C363 VTAIL.n331 B 0.008331f
C364 VTAIL.n332 B 0.015504f
C365 VTAIL.n333 B 0.015504f
C366 VTAIL.n334 B 0.008331f
C367 VTAIL.n335 B 0.008821f
C368 VTAIL.n336 B 0.019692f
C369 VTAIL.n337 B 0.019692f
C370 VTAIL.n338 B 0.008821f
C371 VTAIL.n339 B 0.008331f
C372 VTAIL.n340 B 0.015504f
C373 VTAIL.n341 B 0.015504f
C374 VTAIL.n342 B 0.008331f
C375 VTAIL.n343 B 0.008821f
C376 VTAIL.n344 B 0.019692f
C377 VTAIL.n345 B 0.019692f
C378 VTAIL.n346 B 0.019692f
C379 VTAIL.n347 B 0.008576f
C380 VTAIL.n348 B 0.008331f
C381 VTAIL.n349 B 0.015504f
C382 VTAIL.n350 B 0.015504f
C383 VTAIL.n351 B 0.008331f
C384 VTAIL.n352 B 0.008821f
C385 VTAIL.n353 B 0.019692f
C386 VTAIL.n354 B 0.038746f
C387 VTAIL.n355 B 0.008821f
C388 VTAIL.n356 B 0.008331f
C389 VTAIL.n357 B 0.033931f
C390 VTAIL.n358 B 0.021221f
C391 VTAIL.n359 B 1.14055f
C392 VTAIL.n360 B 0.019596f
C393 VTAIL.n361 B 0.015504f
C394 VTAIL.n362 B 0.008331f
C395 VTAIL.n363 B 0.019692f
C396 VTAIL.n364 B 0.008821f
C397 VTAIL.n365 B 0.015504f
C398 VTAIL.n366 B 0.008576f
C399 VTAIL.n367 B 0.019692f
C400 VTAIL.n368 B 0.008331f
C401 VTAIL.n369 B 0.008821f
C402 VTAIL.n370 B 0.015504f
C403 VTAIL.n371 B 0.008331f
C404 VTAIL.n372 B 0.019692f
C405 VTAIL.n373 B 0.008821f
C406 VTAIL.n374 B 0.015504f
C407 VTAIL.n375 B 0.008331f
C408 VTAIL.n376 B 0.019692f
C409 VTAIL.n377 B 0.008821f
C410 VTAIL.n378 B 0.015504f
C411 VTAIL.n379 B 0.008331f
C412 VTAIL.n380 B 0.019692f
C413 VTAIL.n381 B 0.008821f
C414 VTAIL.n382 B 0.015504f
C415 VTAIL.n383 B 0.008331f
C416 VTAIL.n384 B 0.019692f
C417 VTAIL.n385 B 0.008821f
C418 VTAIL.n386 B 0.015504f
C419 VTAIL.n387 B 0.008331f
C420 VTAIL.n388 B 0.014769f
C421 VTAIL.n389 B 0.011633f
C422 VTAIL.t3 B 0.032523f
C423 VTAIL.n390 B 0.104971f
C424 VTAIL.n391 B 1.07908f
C425 VTAIL.n392 B 0.008331f
C426 VTAIL.n393 B 0.008821f
C427 VTAIL.n394 B 0.019692f
C428 VTAIL.n395 B 0.019692f
C429 VTAIL.n396 B 0.008821f
C430 VTAIL.n397 B 0.008331f
C431 VTAIL.n398 B 0.015504f
C432 VTAIL.n399 B 0.015504f
C433 VTAIL.n400 B 0.008331f
C434 VTAIL.n401 B 0.008821f
C435 VTAIL.n402 B 0.019692f
C436 VTAIL.n403 B 0.019692f
C437 VTAIL.n404 B 0.008821f
C438 VTAIL.n405 B 0.008331f
C439 VTAIL.n406 B 0.015504f
C440 VTAIL.n407 B 0.015504f
C441 VTAIL.n408 B 0.008331f
C442 VTAIL.n409 B 0.008821f
C443 VTAIL.n410 B 0.019692f
C444 VTAIL.n411 B 0.019692f
C445 VTAIL.n412 B 0.008821f
C446 VTAIL.n413 B 0.008331f
C447 VTAIL.n414 B 0.015504f
C448 VTAIL.n415 B 0.015504f
C449 VTAIL.n416 B 0.008331f
C450 VTAIL.n417 B 0.008821f
C451 VTAIL.n418 B 0.019692f
C452 VTAIL.n419 B 0.019692f
C453 VTAIL.n420 B 0.008821f
C454 VTAIL.n421 B 0.008331f
C455 VTAIL.n422 B 0.015504f
C456 VTAIL.n423 B 0.015504f
C457 VTAIL.n424 B 0.008331f
C458 VTAIL.n425 B 0.008821f
C459 VTAIL.n426 B 0.019692f
C460 VTAIL.n427 B 0.019692f
C461 VTAIL.n428 B 0.008821f
C462 VTAIL.n429 B 0.008331f
C463 VTAIL.n430 B 0.015504f
C464 VTAIL.n431 B 0.015504f
C465 VTAIL.n432 B 0.008331f
C466 VTAIL.n433 B 0.008821f
C467 VTAIL.n434 B 0.019692f
C468 VTAIL.n435 B 0.019692f
C469 VTAIL.n436 B 0.019692f
C470 VTAIL.n437 B 0.008576f
C471 VTAIL.n438 B 0.008331f
C472 VTAIL.n439 B 0.015504f
C473 VTAIL.n440 B 0.015504f
C474 VTAIL.n441 B 0.008331f
C475 VTAIL.n442 B 0.008821f
C476 VTAIL.n443 B 0.019692f
C477 VTAIL.n444 B 0.038746f
C478 VTAIL.n445 B 0.008821f
C479 VTAIL.n446 B 0.008331f
C480 VTAIL.n447 B 0.033931f
C481 VTAIL.n448 B 0.021221f
C482 VTAIL.n449 B 0.1502f
C483 VTAIL.n450 B 0.019596f
C484 VTAIL.n451 B 0.015504f
C485 VTAIL.n452 B 0.008331f
C486 VTAIL.n453 B 0.019692f
C487 VTAIL.n454 B 0.008821f
C488 VTAIL.n455 B 0.015504f
C489 VTAIL.n456 B 0.008576f
C490 VTAIL.n457 B 0.019692f
C491 VTAIL.n458 B 0.008331f
C492 VTAIL.n459 B 0.008821f
C493 VTAIL.n460 B 0.015504f
C494 VTAIL.n461 B 0.008331f
C495 VTAIL.n462 B 0.019692f
C496 VTAIL.n463 B 0.008821f
C497 VTAIL.n464 B 0.015504f
C498 VTAIL.n465 B 0.008331f
C499 VTAIL.n466 B 0.019692f
C500 VTAIL.n467 B 0.008821f
C501 VTAIL.n468 B 0.015504f
C502 VTAIL.n469 B 0.008331f
C503 VTAIL.n470 B 0.019692f
C504 VTAIL.n471 B 0.008821f
C505 VTAIL.n472 B 0.015504f
C506 VTAIL.n473 B 0.008331f
C507 VTAIL.n474 B 0.019692f
C508 VTAIL.n475 B 0.008821f
C509 VTAIL.n476 B 0.015504f
C510 VTAIL.n477 B 0.008331f
C511 VTAIL.n478 B 0.014769f
C512 VTAIL.n479 B 0.011633f
C513 VTAIL.t7 B 0.032523f
C514 VTAIL.n480 B 0.104971f
C515 VTAIL.n481 B 1.07908f
C516 VTAIL.n482 B 0.008331f
C517 VTAIL.n483 B 0.008821f
C518 VTAIL.n484 B 0.019692f
C519 VTAIL.n485 B 0.019692f
C520 VTAIL.n486 B 0.008821f
C521 VTAIL.n487 B 0.008331f
C522 VTAIL.n488 B 0.015504f
C523 VTAIL.n489 B 0.015504f
C524 VTAIL.n490 B 0.008331f
C525 VTAIL.n491 B 0.008821f
C526 VTAIL.n492 B 0.019692f
C527 VTAIL.n493 B 0.019692f
C528 VTAIL.n494 B 0.008821f
C529 VTAIL.n495 B 0.008331f
C530 VTAIL.n496 B 0.015504f
C531 VTAIL.n497 B 0.015504f
C532 VTAIL.n498 B 0.008331f
C533 VTAIL.n499 B 0.008821f
C534 VTAIL.n500 B 0.019692f
C535 VTAIL.n501 B 0.019692f
C536 VTAIL.n502 B 0.008821f
C537 VTAIL.n503 B 0.008331f
C538 VTAIL.n504 B 0.015504f
C539 VTAIL.n505 B 0.015504f
C540 VTAIL.n506 B 0.008331f
C541 VTAIL.n507 B 0.008821f
C542 VTAIL.n508 B 0.019692f
C543 VTAIL.n509 B 0.019692f
C544 VTAIL.n510 B 0.008821f
C545 VTAIL.n511 B 0.008331f
C546 VTAIL.n512 B 0.015504f
C547 VTAIL.n513 B 0.015504f
C548 VTAIL.n514 B 0.008331f
C549 VTAIL.n515 B 0.008821f
C550 VTAIL.n516 B 0.019692f
C551 VTAIL.n517 B 0.019692f
C552 VTAIL.n518 B 0.008821f
C553 VTAIL.n519 B 0.008331f
C554 VTAIL.n520 B 0.015504f
C555 VTAIL.n521 B 0.015504f
C556 VTAIL.n522 B 0.008331f
C557 VTAIL.n523 B 0.008821f
C558 VTAIL.n524 B 0.019692f
C559 VTAIL.n525 B 0.019692f
C560 VTAIL.n526 B 0.019692f
C561 VTAIL.n527 B 0.008576f
C562 VTAIL.n528 B 0.008331f
C563 VTAIL.n529 B 0.015504f
C564 VTAIL.n530 B 0.015504f
C565 VTAIL.n531 B 0.008331f
C566 VTAIL.n532 B 0.008821f
C567 VTAIL.n533 B 0.019692f
C568 VTAIL.n534 B 0.038746f
C569 VTAIL.n535 B 0.008821f
C570 VTAIL.n536 B 0.008331f
C571 VTAIL.n537 B 0.033931f
C572 VTAIL.n538 B 0.021221f
C573 VTAIL.n539 B 0.1502f
C574 VTAIL.n540 B 0.019596f
C575 VTAIL.n541 B 0.015504f
C576 VTAIL.n542 B 0.008331f
C577 VTAIL.n543 B 0.019692f
C578 VTAIL.n544 B 0.008821f
C579 VTAIL.n545 B 0.015504f
C580 VTAIL.n546 B 0.008576f
C581 VTAIL.n547 B 0.019692f
C582 VTAIL.n548 B 0.008331f
C583 VTAIL.n549 B 0.008821f
C584 VTAIL.n550 B 0.015504f
C585 VTAIL.n551 B 0.008331f
C586 VTAIL.n552 B 0.019692f
C587 VTAIL.n553 B 0.008821f
C588 VTAIL.n554 B 0.015504f
C589 VTAIL.n555 B 0.008331f
C590 VTAIL.n556 B 0.019692f
C591 VTAIL.n557 B 0.008821f
C592 VTAIL.n558 B 0.015504f
C593 VTAIL.n559 B 0.008331f
C594 VTAIL.n560 B 0.019692f
C595 VTAIL.n561 B 0.008821f
C596 VTAIL.n562 B 0.015504f
C597 VTAIL.n563 B 0.008331f
C598 VTAIL.n564 B 0.019692f
C599 VTAIL.n565 B 0.008821f
C600 VTAIL.n566 B 0.015504f
C601 VTAIL.n567 B 0.008331f
C602 VTAIL.n568 B 0.014769f
C603 VTAIL.n569 B 0.011633f
C604 VTAIL.t6 B 0.032523f
C605 VTAIL.n570 B 0.104971f
C606 VTAIL.n571 B 1.07908f
C607 VTAIL.n572 B 0.008331f
C608 VTAIL.n573 B 0.008821f
C609 VTAIL.n574 B 0.019692f
C610 VTAIL.n575 B 0.019692f
C611 VTAIL.n576 B 0.008821f
C612 VTAIL.n577 B 0.008331f
C613 VTAIL.n578 B 0.015504f
C614 VTAIL.n579 B 0.015504f
C615 VTAIL.n580 B 0.008331f
C616 VTAIL.n581 B 0.008821f
C617 VTAIL.n582 B 0.019692f
C618 VTAIL.n583 B 0.019692f
C619 VTAIL.n584 B 0.008821f
C620 VTAIL.n585 B 0.008331f
C621 VTAIL.n586 B 0.015504f
C622 VTAIL.n587 B 0.015504f
C623 VTAIL.n588 B 0.008331f
C624 VTAIL.n589 B 0.008821f
C625 VTAIL.n590 B 0.019692f
C626 VTAIL.n591 B 0.019692f
C627 VTAIL.n592 B 0.008821f
C628 VTAIL.n593 B 0.008331f
C629 VTAIL.n594 B 0.015504f
C630 VTAIL.n595 B 0.015504f
C631 VTAIL.n596 B 0.008331f
C632 VTAIL.n597 B 0.008821f
C633 VTAIL.n598 B 0.019692f
C634 VTAIL.n599 B 0.019692f
C635 VTAIL.n600 B 0.008821f
C636 VTAIL.n601 B 0.008331f
C637 VTAIL.n602 B 0.015504f
C638 VTAIL.n603 B 0.015504f
C639 VTAIL.n604 B 0.008331f
C640 VTAIL.n605 B 0.008821f
C641 VTAIL.n606 B 0.019692f
C642 VTAIL.n607 B 0.019692f
C643 VTAIL.n608 B 0.008821f
C644 VTAIL.n609 B 0.008331f
C645 VTAIL.n610 B 0.015504f
C646 VTAIL.n611 B 0.015504f
C647 VTAIL.n612 B 0.008331f
C648 VTAIL.n613 B 0.008821f
C649 VTAIL.n614 B 0.019692f
C650 VTAIL.n615 B 0.019692f
C651 VTAIL.n616 B 0.019692f
C652 VTAIL.n617 B 0.008576f
C653 VTAIL.n618 B 0.008331f
C654 VTAIL.n619 B 0.015504f
C655 VTAIL.n620 B 0.015504f
C656 VTAIL.n621 B 0.008331f
C657 VTAIL.n622 B 0.008821f
C658 VTAIL.n623 B 0.019692f
C659 VTAIL.n624 B 0.038746f
C660 VTAIL.n625 B 0.008821f
C661 VTAIL.n626 B 0.008331f
C662 VTAIL.n627 B 0.033931f
C663 VTAIL.n628 B 0.021221f
C664 VTAIL.n629 B 1.14055f
C665 VTAIL.n630 B 0.019596f
C666 VTAIL.n631 B 0.015504f
C667 VTAIL.n632 B 0.008331f
C668 VTAIL.n633 B 0.019692f
C669 VTAIL.n634 B 0.008821f
C670 VTAIL.n635 B 0.015504f
C671 VTAIL.n636 B 0.008576f
C672 VTAIL.n637 B 0.019692f
C673 VTAIL.n638 B 0.008821f
C674 VTAIL.n639 B 0.015504f
C675 VTAIL.n640 B 0.008331f
C676 VTAIL.n641 B 0.019692f
C677 VTAIL.n642 B 0.008821f
C678 VTAIL.n643 B 0.015504f
C679 VTAIL.n644 B 0.008331f
C680 VTAIL.n645 B 0.019692f
C681 VTAIL.n646 B 0.008821f
C682 VTAIL.n647 B 0.015504f
C683 VTAIL.n648 B 0.008331f
C684 VTAIL.n649 B 0.019692f
C685 VTAIL.n650 B 0.008821f
C686 VTAIL.n651 B 0.015504f
C687 VTAIL.n652 B 0.008331f
C688 VTAIL.n653 B 0.019692f
C689 VTAIL.n654 B 0.008821f
C690 VTAIL.n655 B 0.015504f
C691 VTAIL.n656 B 0.008331f
C692 VTAIL.n657 B 0.014769f
C693 VTAIL.n658 B 0.011633f
C694 VTAIL.t1 B 0.032523f
C695 VTAIL.n659 B 0.104971f
C696 VTAIL.n660 B 1.07908f
C697 VTAIL.n661 B 0.008331f
C698 VTAIL.n662 B 0.008821f
C699 VTAIL.n663 B 0.019692f
C700 VTAIL.n664 B 0.019692f
C701 VTAIL.n665 B 0.008821f
C702 VTAIL.n666 B 0.008331f
C703 VTAIL.n667 B 0.015504f
C704 VTAIL.n668 B 0.015504f
C705 VTAIL.n669 B 0.008331f
C706 VTAIL.n670 B 0.008821f
C707 VTAIL.n671 B 0.019692f
C708 VTAIL.n672 B 0.019692f
C709 VTAIL.n673 B 0.008821f
C710 VTAIL.n674 B 0.008331f
C711 VTAIL.n675 B 0.015504f
C712 VTAIL.n676 B 0.015504f
C713 VTAIL.n677 B 0.008331f
C714 VTAIL.n678 B 0.008821f
C715 VTAIL.n679 B 0.019692f
C716 VTAIL.n680 B 0.019692f
C717 VTAIL.n681 B 0.008821f
C718 VTAIL.n682 B 0.008331f
C719 VTAIL.n683 B 0.015504f
C720 VTAIL.n684 B 0.015504f
C721 VTAIL.n685 B 0.008331f
C722 VTAIL.n686 B 0.008821f
C723 VTAIL.n687 B 0.019692f
C724 VTAIL.n688 B 0.019692f
C725 VTAIL.n689 B 0.008821f
C726 VTAIL.n690 B 0.008331f
C727 VTAIL.n691 B 0.015504f
C728 VTAIL.n692 B 0.015504f
C729 VTAIL.n693 B 0.008331f
C730 VTAIL.n694 B 0.008821f
C731 VTAIL.n695 B 0.019692f
C732 VTAIL.n696 B 0.019692f
C733 VTAIL.n697 B 0.008821f
C734 VTAIL.n698 B 0.008331f
C735 VTAIL.n699 B 0.015504f
C736 VTAIL.n700 B 0.015504f
C737 VTAIL.n701 B 0.008331f
C738 VTAIL.n702 B 0.008331f
C739 VTAIL.n703 B 0.008821f
C740 VTAIL.n704 B 0.019692f
C741 VTAIL.n705 B 0.019692f
C742 VTAIL.n706 B 0.019692f
C743 VTAIL.n707 B 0.008576f
C744 VTAIL.n708 B 0.008331f
C745 VTAIL.n709 B 0.015504f
C746 VTAIL.n710 B 0.015504f
C747 VTAIL.n711 B 0.008331f
C748 VTAIL.n712 B 0.008821f
C749 VTAIL.n713 B 0.019692f
C750 VTAIL.n714 B 0.038746f
C751 VTAIL.n715 B 0.008821f
C752 VTAIL.n716 B 0.008331f
C753 VTAIL.n717 B 0.033931f
C754 VTAIL.n718 B 0.021221f
C755 VTAIL.n719 B 1.08036f
C756 VDD1.t2 B 0.337682f
C757 VDD1.t3 B 0.337682f
C758 VDD1.n0 B 3.05899f
C759 VDD1.t1 B 0.337682f
C760 VDD1.t0 B 0.337682f
C761 VDD1.n1 B 3.91036f
C762 VP.n0 B 0.035178f
C763 VP.t2 B 2.72666f
C764 VP.n1 B 0.02157f
C765 VP.n2 B 0.035178f
C766 VP.t3 B 2.72666f
C767 VP.t1 B 2.9245f
C768 VP.t0 B 2.92806f
C769 VP.n3 B 3.37654f
C770 VP.n4 B 1.60116f
C771 VP.n5 B 1.0422f
C772 VP.n6 B 0.041381f
C773 VP.n7 B 0.05303f
C774 VP.n8 B 0.026682f
C775 VP.n9 B 0.026682f
C776 VP.n10 B 0.026682f
C777 VP.n11 B 0.05303f
C778 VP.n12 B 0.041381f
C779 VP.n13 B 1.0422f
C780 VP.n14 B 0.03693f
.ends

