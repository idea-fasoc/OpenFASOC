* NGSPICE file created from diff_pair_sample_0278.ext - technology: sky130A

.subckt diff_pair_sample_0278 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=0.21
X1 VDD2.t2 VN.t1 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=0.21
X2 VTAIL.t7 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=0.21
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=0.21
X4 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=0.21
X5 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=0.21
X6 VDD1.t1 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94195 pd=18.16 as=6.9537 ps=36.44 w=17.83 l=0.21
X7 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=0.21
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=0.21
X9 VTAIL.t5 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=2.94195 ps=18.16 w=17.83 l=0.21
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=0.21
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.9537 pd=36.44 as=0 ps=0 w=17.83 l=0.21
R0 VN.n0 VN.t1 2235.98
R1 VN.n0 VN.t3 2235.98
R2 VN.n1 VN.t2 2235.98
R3 VN.n1 VN.t0 2235.98
R4 VN VN.n1 205.044
R5 VN VN.n0 161.351
R6 VTAIL.n5 VTAIL.t1 44.126
R7 VTAIL.n4 VTAIL.t6 44.126
R8 VTAIL.n3 VTAIL.t7 44.126
R9 VTAIL.n7 VTAIL.t4 44.1258
R10 VTAIL.n0 VTAIL.t5 44.1258
R11 VTAIL.n1 VTAIL.t2 44.1258
R12 VTAIL.n2 VTAIL.t3 44.1258
R13 VTAIL.n6 VTAIL.t0 44.1258
R14 VTAIL.n7 VTAIL.n6 28.2203
R15 VTAIL.n3 VTAIL.n2 28.2203
R16 VTAIL.n5 VTAIL.n4 0.470328
R17 VTAIL.n1 VTAIL.n0 0.470328
R18 VTAIL.n4 VTAIL.n3 0.466017
R19 VTAIL.n6 VTAIL.n5 0.466017
R20 VTAIL.n2 VTAIL.n1 0.466017
R21 VTAIL VTAIL.n0 0.291448
R22 VTAIL VTAIL.n7 0.175069
R23 VDD2.n2 VDD2.n0 100.194
R24 VDD2.n2 VDD2.n1 59.6941
R25 VDD2.n1 VDD2.t1 1.11099
R26 VDD2.n1 VDD2.t3 1.11099
R27 VDD2.n0 VDD2.t0 1.11099
R28 VDD2.n0 VDD2.t2 1.11099
R29 VDD2 VDD2.n2 0.0586897
R30 B.n439 B.t8 2279.69
R31 B.n436 B.t12 2279.69
R32 B.n94 B.t15 2279.69
R33 B.n91 B.t4 2279.69
R34 B.n753 B.n752 585
R35 B.n754 B.n753 585
R36 B.n347 B.n90 585
R37 B.n346 B.n345 585
R38 B.n344 B.n343 585
R39 B.n342 B.n341 585
R40 B.n340 B.n339 585
R41 B.n338 B.n337 585
R42 B.n336 B.n335 585
R43 B.n334 B.n333 585
R44 B.n332 B.n331 585
R45 B.n330 B.n329 585
R46 B.n328 B.n327 585
R47 B.n326 B.n325 585
R48 B.n324 B.n323 585
R49 B.n322 B.n321 585
R50 B.n320 B.n319 585
R51 B.n318 B.n317 585
R52 B.n316 B.n315 585
R53 B.n314 B.n313 585
R54 B.n312 B.n311 585
R55 B.n310 B.n309 585
R56 B.n308 B.n307 585
R57 B.n306 B.n305 585
R58 B.n304 B.n303 585
R59 B.n302 B.n301 585
R60 B.n300 B.n299 585
R61 B.n298 B.n297 585
R62 B.n296 B.n295 585
R63 B.n294 B.n293 585
R64 B.n292 B.n291 585
R65 B.n290 B.n289 585
R66 B.n288 B.n287 585
R67 B.n286 B.n285 585
R68 B.n284 B.n283 585
R69 B.n282 B.n281 585
R70 B.n280 B.n279 585
R71 B.n278 B.n277 585
R72 B.n276 B.n275 585
R73 B.n274 B.n273 585
R74 B.n272 B.n271 585
R75 B.n270 B.n269 585
R76 B.n268 B.n267 585
R77 B.n266 B.n265 585
R78 B.n264 B.n263 585
R79 B.n262 B.n261 585
R80 B.n260 B.n259 585
R81 B.n258 B.n257 585
R82 B.n256 B.n255 585
R83 B.n254 B.n253 585
R84 B.n252 B.n251 585
R85 B.n250 B.n249 585
R86 B.n248 B.n247 585
R87 B.n246 B.n245 585
R88 B.n244 B.n243 585
R89 B.n242 B.n241 585
R90 B.n240 B.n239 585
R91 B.n238 B.n237 585
R92 B.n236 B.n235 585
R93 B.n234 B.n233 585
R94 B.n232 B.n231 585
R95 B.n230 B.n229 585
R96 B.n228 B.n227 585
R97 B.n226 B.n225 585
R98 B.n224 B.n223 585
R99 B.n222 B.n221 585
R100 B.n220 B.n219 585
R101 B.n218 B.n217 585
R102 B.n216 B.n215 585
R103 B.n213 B.n212 585
R104 B.n211 B.n210 585
R105 B.n209 B.n208 585
R106 B.n207 B.n206 585
R107 B.n205 B.n204 585
R108 B.n203 B.n202 585
R109 B.n201 B.n200 585
R110 B.n199 B.n198 585
R111 B.n197 B.n196 585
R112 B.n195 B.n194 585
R113 B.n193 B.n192 585
R114 B.n191 B.n190 585
R115 B.n189 B.n188 585
R116 B.n187 B.n186 585
R117 B.n185 B.n184 585
R118 B.n183 B.n182 585
R119 B.n181 B.n180 585
R120 B.n179 B.n178 585
R121 B.n177 B.n176 585
R122 B.n175 B.n174 585
R123 B.n173 B.n172 585
R124 B.n171 B.n170 585
R125 B.n169 B.n168 585
R126 B.n167 B.n166 585
R127 B.n165 B.n164 585
R128 B.n163 B.n162 585
R129 B.n161 B.n160 585
R130 B.n159 B.n158 585
R131 B.n157 B.n156 585
R132 B.n155 B.n154 585
R133 B.n153 B.n152 585
R134 B.n151 B.n150 585
R135 B.n149 B.n148 585
R136 B.n147 B.n146 585
R137 B.n145 B.n144 585
R138 B.n143 B.n142 585
R139 B.n141 B.n140 585
R140 B.n139 B.n138 585
R141 B.n137 B.n136 585
R142 B.n135 B.n134 585
R143 B.n133 B.n132 585
R144 B.n131 B.n130 585
R145 B.n129 B.n128 585
R146 B.n127 B.n126 585
R147 B.n125 B.n124 585
R148 B.n123 B.n122 585
R149 B.n121 B.n120 585
R150 B.n119 B.n118 585
R151 B.n117 B.n116 585
R152 B.n115 B.n114 585
R153 B.n113 B.n112 585
R154 B.n111 B.n110 585
R155 B.n109 B.n108 585
R156 B.n107 B.n106 585
R157 B.n105 B.n104 585
R158 B.n103 B.n102 585
R159 B.n101 B.n100 585
R160 B.n99 B.n98 585
R161 B.n97 B.n96 585
R162 B.n751 B.n26 585
R163 B.n755 B.n26 585
R164 B.n750 B.n25 585
R165 B.n756 B.n25 585
R166 B.n749 B.n748 585
R167 B.n748 B.n21 585
R168 B.n747 B.n20 585
R169 B.n762 B.n20 585
R170 B.n746 B.n19 585
R171 B.n763 B.n19 585
R172 B.n745 B.n18 585
R173 B.n764 B.n18 585
R174 B.n744 B.n743 585
R175 B.n743 B.n14 585
R176 B.n742 B.n13 585
R177 B.n770 B.n13 585
R178 B.n741 B.n12 585
R179 B.n771 B.n12 585
R180 B.n740 B.n11 585
R181 B.n772 B.n11 585
R182 B.n739 B.n738 585
R183 B.n738 B.n737 585
R184 B.n736 B.n7 585
R185 B.n778 B.n7 585
R186 B.n735 B.n6 585
R187 B.n779 B.n6 585
R188 B.n734 B.n5 585
R189 B.n780 B.n5 585
R190 B.n733 B.n732 585
R191 B.n732 B.n4 585
R192 B.n731 B.n348 585
R193 B.n731 B.n730 585
R194 B.n720 B.n349 585
R195 B.n723 B.n349 585
R196 B.n722 B.n721 585
R197 B.n724 B.n722 585
R198 B.n719 B.n354 585
R199 B.n354 B.n353 585
R200 B.n718 B.n717 585
R201 B.n717 B.n716 585
R202 B.n356 B.n355 585
R203 B.n357 B.n356 585
R204 B.n709 B.n708 585
R205 B.n710 B.n709 585
R206 B.n707 B.n361 585
R207 B.n365 B.n361 585
R208 B.n706 B.n705 585
R209 B.n705 B.n704 585
R210 B.n363 B.n362 585
R211 B.n364 B.n363 585
R212 B.n697 B.n696 585
R213 B.n698 B.n697 585
R214 B.n695 B.n370 585
R215 B.n370 B.n369 585
R216 B.n689 B.n688 585
R217 B.n687 B.n435 585
R218 B.n686 B.n434 585
R219 B.n691 B.n434 585
R220 B.n685 B.n684 585
R221 B.n683 B.n682 585
R222 B.n681 B.n680 585
R223 B.n679 B.n678 585
R224 B.n677 B.n676 585
R225 B.n675 B.n674 585
R226 B.n673 B.n672 585
R227 B.n671 B.n670 585
R228 B.n669 B.n668 585
R229 B.n667 B.n666 585
R230 B.n665 B.n664 585
R231 B.n663 B.n662 585
R232 B.n661 B.n660 585
R233 B.n659 B.n658 585
R234 B.n657 B.n656 585
R235 B.n655 B.n654 585
R236 B.n653 B.n652 585
R237 B.n651 B.n650 585
R238 B.n649 B.n648 585
R239 B.n647 B.n646 585
R240 B.n645 B.n644 585
R241 B.n643 B.n642 585
R242 B.n641 B.n640 585
R243 B.n639 B.n638 585
R244 B.n637 B.n636 585
R245 B.n635 B.n634 585
R246 B.n633 B.n632 585
R247 B.n631 B.n630 585
R248 B.n629 B.n628 585
R249 B.n627 B.n626 585
R250 B.n625 B.n624 585
R251 B.n623 B.n622 585
R252 B.n621 B.n620 585
R253 B.n619 B.n618 585
R254 B.n617 B.n616 585
R255 B.n615 B.n614 585
R256 B.n613 B.n612 585
R257 B.n611 B.n610 585
R258 B.n609 B.n608 585
R259 B.n607 B.n606 585
R260 B.n605 B.n604 585
R261 B.n603 B.n602 585
R262 B.n601 B.n600 585
R263 B.n599 B.n598 585
R264 B.n597 B.n596 585
R265 B.n595 B.n594 585
R266 B.n593 B.n592 585
R267 B.n591 B.n590 585
R268 B.n589 B.n588 585
R269 B.n587 B.n586 585
R270 B.n585 B.n584 585
R271 B.n583 B.n582 585
R272 B.n581 B.n580 585
R273 B.n579 B.n578 585
R274 B.n577 B.n576 585
R275 B.n575 B.n574 585
R276 B.n573 B.n572 585
R277 B.n571 B.n570 585
R278 B.n569 B.n568 585
R279 B.n567 B.n566 585
R280 B.n565 B.n564 585
R281 B.n563 B.n562 585
R282 B.n561 B.n560 585
R283 B.n559 B.n558 585
R284 B.n557 B.n556 585
R285 B.n554 B.n553 585
R286 B.n552 B.n551 585
R287 B.n550 B.n549 585
R288 B.n548 B.n547 585
R289 B.n546 B.n545 585
R290 B.n544 B.n543 585
R291 B.n542 B.n541 585
R292 B.n540 B.n539 585
R293 B.n538 B.n537 585
R294 B.n536 B.n535 585
R295 B.n534 B.n533 585
R296 B.n532 B.n531 585
R297 B.n530 B.n529 585
R298 B.n528 B.n527 585
R299 B.n526 B.n525 585
R300 B.n524 B.n523 585
R301 B.n522 B.n521 585
R302 B.n520 B.n519 585
R303 B.n518 B.n517 585
R304 B.n516 B.n515 585
R305 B.n514 B.n513 585
R306 B.n512 B.n511 585
R307 B.n510 B.n509 585
R308 B.n508 B.n507 585
R309 B.n506 B.n505 585
R310 B.n504 B.n503 585
R311 B.n502 B.n501 585
R312 B.n500 B.n499 585
R313 B.n498 B.n497 585
R314 B.n496 B.n495 585
R315 B.n494 B.n493 585
R316 B.n492 B.n491 585
R317 B.n490 B.n489 585
R318 B.n488 B.n487 585
R319 B.n486 B.n485 585
R320 B.n484 B.n483 585
R321 B.n482 B.n481 585
R322 B.n480 B.n479 585
R323 B.n478 B.n477 585
R324 B.n476 B.n475 585
R325 B.n474 B.n473 585
R326 B.n472 B.n471 585
R327 B.n470 B.n469 585
R328 B.n468 B.n467 585
R329 B.n466 B.n465 585
R330 B.n464 B.n463 585
R331 B.n462 B.n461 585
R332 B.n460 B.n459 585
R333 B.n458 B.n457 585
R334 B.n456 B.n455 585
R335 B.n454 B.n453 585
R336 B.n452 B.n451 585
R337 B.n450 B.n449 585
R338 B.n448 B.n447 585
R339 B.n446 B.n445 585
R340 B.n444 B.n443 585
R341 B.n442 B.n441 585
R342 B.n372 B.n371 585
R343 B.n694 B.n693 585
R344 B.n368 B.n367 585
R345 B.n369 B.n368 585
R346 B.n700 B.n699 585
R347 B.n699 B.n698 585
R348 B.n701 B.n366 585
R349 B.n366 B.n364 585
R350 B.n703 B.n702 585
R351 B.n704 B.n703 585
R352 B.n360 B.n359 585
R353 B.n365 B.n360 585
R354 B.n712 B.n711 585
R355 B.n711 B.n710 585
R356 B.n713 B.n358 585
R357 B.n358 B.n357 585
R358 B.n715 B.n714 585
R359 B.n716 B.n715 585
R360 B.n352 B.n351 585
R361 B.n353 B.n352 585
R362 B.n726 B.n725 585
R363 B.n725 B.n724 585
R364 B.n727 B.n350 585
R365 B.n723 B.n350 585
R366 B.n729 B.n728 585
R367 B.n730 B.n729 585
R368 B.n2 B.n0 585
R369 B.n4 B.n2 585
R370 B.n3 B.n1 585
R371 B.n779 B.n3 585
R372 B.n777 B.n776 585
R373 B.n778 B.n777 585
R374 B.n775 B.n8 585
R375 B.n737 B.n8 585
R376 B.n774 B.n773 585
R377 B.n773 B.n772 585
R378 B.n10 B.n9 585
R379 B.n771 B.n10 585
R380 B.n769 B.n768 585
R381 B.n770 B.n769 585
R382 B.n767 B.n15 585
R383 B.n15 B.n14 585
R384 B.n766 B.n765 585
R385 B.n765 B.n764 585
R386 B.n17 B.n16 585
R387 B.n763 B.n17 585
R388 B.n761 B.n760 585
R389 B.n762 B.n761 585
R390 B.n759 B.n22 585
R391 B.n22 B.n21 585
R392 B.n758 B.n757 585
R393 B.n757 B.n756 585
R394 B.n24 B.n23 585
R395 B.n755 B.n24 585
R396 B.n782 B.n781 585
R397 B.n781 B.n780 585
R398 B.n689 B.n368 497.305
R399 B.n96 B.n24 497.305
R400 B.n693 B.n370 497.305
R401 B.n753 B.n26 497.305
R402 B.n754 B.n89 256.663
R403 B.n754 B.n88 256.663
R404 B.n754 B.n87 256.663
R405 B.n754 B.n86 256.663
R406 B.n754 B.n85 256.663
R407 B.n754 B.n84 256.663
R408 B.n754 B.n83 256.663
R409 B.n754 B.n82 256.663
R410 B.n754 B.n81 256.663
R411 B.n754 B.n80 256.663
R412 B.n754 B.n79 256.663
R413 B.n754 B.n78 256.663
R414 B.n754 B.n77 256.663
R415 B.n754 B.n76 256.663
R416 B.n754 B.n75 256.663
R417 B.n754 B.n74 256.663
R418 B.n754 B.n73 256.663
R419 B.n754 B.n72 256.663
R420 B.n754 B.n71 256.663
R421 B.n754 B.n70 256.663
R422 B.n754 B.n69 256.663
R423 B.n754 B.n68 256.663
R424 B.n754 B.n67 256.663
R425 B.n754 B.n66 256.663
R426 B.n754 B.n65 256.663
R427 B.n754 B.n64 256.663
R428 B.n754 B.n63 256.663
R429 B.n754 B.n62 256.663
R430 B.n754 B.n61 256.663
R431 B.n754 B.n60 256.663
R432 B.n754 B.n59 256.663
R433 B.n754 B.n58 256.663
R434 B.n754 B.n57 256.663
R435 B.n754 B.n56 256.663
R436 B.n754 B.n55 256.663
R437 B.n754 B.n54 256.663
R438 B.n754 B.n53 256.663
R439 B.n754 B.n52 256.663
R440 B.n754 B.n51 256.663
R441 B.n754 B.n50 256.663
R442 B.n754 B.n49 256.663
R443 B.n754 B.n48 256.663
R444 B.n754 B.n47 256.663
R445 B.n754 B.n46 256.663
R446 B.n754 B.n45 256.663
R447 B.n754 B.n44 256.663
R448 B.n754 B.n43 256.663
R449 B.n754 B.n42 256.663
R450 B.n754 B.n41 256.663
R451 B.n754 B.n40 256.663
R452 B.n754 B.n39 256.663
R453 B.n754 B.n38 256.663
R454 B.n754 B.n37 256.663
R455 B.n754 B.n36 256.663
R456 B.n754 B.n35 256.663
R457 B.n754 B.n34 256.663
R458 B.n754 B.n33 256.663
R459 B.n754 B.n32 256.663
R460 B.n754 B.n31 256.663
R461 B.n754 B.n30 256.663
R462 B.n754 B.n29 256.663
R463 B.n754 B.n28 256.663
R464 B.n754 B.n27 256.663
R465 B.n691 B.n690 256.663
R466 B.n691 B.n373 256.663
R467 B.n691 B.n374 256.663
R468 B.n691 B.n375 256.663
R469 B.n691 B.n376 256.663
R470 B.n691 B.n377 256.663
R471 B.n691 B.n378 256.663
R472 B.n691 B.n379 256.663
R473 B.n691 B.n380 256.663
R474 B.n691 B.n381 256.663
R475 B.n691 B.n382 256.663
R476 B.n691 B.n383 256.663
R477 B.n691 B.n384 256.663
R478 B.n691 B.n385 256.663
R479 B.n691 B.n386 256.663
R480 B.n691 B.n387 256.663
R481 B.n691 B.n388 256.663
R482 B.n691 B.n389 256.663
R483 B.n691 B.n390 256.663
R484 B.n691 B.n391 256.663
R485 B.n691 B.n392 256.663
R486 B.n691 B.n393 256.663
R487 B.n691 B.n394 256.663
R488 B.n691 B.n395 256.663
R489 B.n691 B.n396 256.663
R490 B.n691 B.n397 256.663
R491 B.n691 B.n398 256.663
R492 B.n691 B.n399 256.663
R493 B.n691 B.n400 256.663
R494 B.n691 B.n401 256.663
R495 B.n691 B.n402 256.663
R496 B.n691 B.n403 256.663
R497 B.n691 B.n404 256.663
R498 B.n691 B.n405 256.663
R499 B.n691 B.n406 256.663
R500 B.n691 B.n407 256.663
R501 B.n691 B.n408 256.663
R502 B.n691 B.n409 256.663
R503 B.n691 B.n410 256.663
R504 B.n691 B.n411 256.663
R505 B.n691 B.n412 256.663
R506 B.n691 B.n413 256.663
R507 B.n691 B.n414 256.663
R508 B.n691 B.n415 256.663
R509 B.n691 B.n416 256.663
R510 B.n691 B.n417 256.663
R511 B.n691 B.n418 256.663
R512 B.n691 B.n419 256.663
R513 B.n691 B.n420 256.663
R514 B.n691 B.n421 256.663
R515 B.n691 B.n422 256.663
R516 B.n691 B.n423 256.663
R517 B.n691 B.n424 256.663
R518 B.n691 B.n425 256.663
R519 B.n691 B.n426 256.663
R520 B.n691 B.n427 256.663
R521 B.n691 B.n428 256.663
R522 B.n691 B.n429 256.663
R523 B.n691 B.n430 256.663
R524 B.n691 B.n431 256.663
R525 B.n691 B.n432 256.663
R526 B.n691 B.n433 256.663
R527 B.n692 B.n691 256.663
R528 B.n699 B.n368 163.367
R529 B.n699 B.n366 163.367
R530 B.n703 B.n366 163.367
R531 B.n703 B.n360 163.367
R532 B.n711 B.n360 163.367
R533 B.n711 B.n358 163.367
R534 B.n715 B.n358 163.367
R535 B.n715 B.n352 163.367
R536 B.n725 B.n352 163.367
R537 B.n725 B.n350 163.367
R538 B.n729 B.n350 163.367
R539 B.n729 B.n2 163.367
R540 B.n781 B.n2 163.367
R541 B.n781 B.n3 163.367
R542 B.n777 B.n3 163.367
R543 B.n777 B.n8 163.367
R544 B.n773 B.n8 163.367
R545 B.n773 B.n10 163.367
R546 B.n769 B.n10 163.367
R547 B.n769 B.n15 163.367
R548 B.n765 B.n15 163.367
R549 B.n765 B.n17 163.367
R550 B.n761 B.n17 163.367
R551 B.n761 B.n22 163.367
R552 B.n757 B.n22 163.367
R553 B.n757 B.n24 163.367
R554 B.n435 B.n434 163.367
R555 B.n684 B.n434 163.367
R556 B.n682 B.n681 163.367
R557 B.n678 B.n677 163.367
R558 B.n674 B.n673 163.367
R559 B.n670 B.n669 163.367
R560 B.n666 B.n665 163.367
R561 B.n662 B.n661 163.367
R562 B.n658 B.n657 163.367
R563 B.n654 B.n653 163.367
R564 B.n650 B.n649 163.367
R565 B.n646 B.n645 163.367
R566 B.n642 B.n641 163.367
R567 B.n638 B.n637 163.367
R568 B.n634 B.n633 163.367
R569 B.n630 B.n629 163.367
R570 B.n626 B.n625 163.367
R571 B.n622 B.n621 163.367
R572 B.n618 B.n617 163.367
R573 B.n614 B.n613 163.367
R574 B.n610 B.n609 163.367
R575 B.n606 B.n605 163.367
R576 B.n602 B.n601 163.367
R577 B.n598 B.n597 163.367
R578 B.n594 B.n593 163.367
R579 B.n590 B.n589 163.367
R580 B.n586 B.n585 163.367
R581 B.n582 B.n581 163.367
R582 B.n578 B.n577 163.367
R583 B.n574 B.n573 163.367
R584 B.n570 B.n569 163.367
R585 B.n566 B.n565 163.367
R586 B.n562 B.n561 163.367
R587 B.n558 B.n557 163.367
R588 B.n553 B.n552 163.367
R589 B.n549 B.n548 163.367
R590 B.n545 B.n544 163.367
R591 B.n541 B.n540 163.367
R592 B.n537 B.n536 163.367
R593 B.n533 B.n532 163.367
R594 B.n529 B.n528 163.367
R595 B.n525 B.n524 163.367
R596 B.n521 B.n520 163.367
R597 B.n517 B.n516 163.367
R598 B.n513 B.n512 163.367
R599 B.n509 B.n508 163.367
R600 B.n505 B.n504 163.367
R601 B.n501 B.n500 163.367
R602 B.n497 B.n496 163.367
R603 B.n493 B.n492 163.367
R604 B.n489 B.n488 163.367
R605 B.n485 B.n484 163.367
R606 B.n481 B.n480 163.367
R607 B.n477 B.n476 163.367
R608 B.n473 B.n472 163.367
R609 B.n469 B.n468 163.367
R610 B.n465 B.n464 163.367
R611 B.n461 B.n460 163.367
R612 B.n457 B.n456 163.367
R613 B.n453 B.n452 163.367
R614 B.n449 B.n448 163.367
R615 B.n445 B.n444 163.367
R616 B.n441 B.n372 163.367
R617 B.n697 B.n370 163.367
R618 B.n697 B.n363 163.367
R619 B.n705 B.n363 163.367
R620 B.n705 B.n361 163.367
R621 B.n709 B.n361 163.367
R622 B.n709 B.n356 163.367
R623 B.n717 B.n356 163.367
R624 B.n717 B.n354 163.367
R625 B.n722 B.n354 163.367
R626 B.n722 B.n349 163.367
R627 B.n731 B.n349 163.367
R628 B.n732 B.n731 163.367
R629 B.n732 B.n5 163.367
R630 B.n6 B.n5 163.367
R631 B.n7 B.n6 163.367
R632 B.n738 B.n7 163.367
R633 B.n738 B.n11 163.367
R634 B.n12 B.n11 163.367
R635 B.n13 B.n12 163.367
R636 B.n743 B.n13 163.367
R637 B.n743 B.n18 163.367
R638 B.n19 B.n18 163.367
R639 B.n20 B.n19 163.367
R640 B.n748 B.n20 163.367
R641 B.n748 B.n25 163.367
R642 B.n26 B.n25 163.367
R643 B.n100 B.n99 163.367
R644 B.n104 B.n103 163.367
R645 B.n108 B.n107 163.367
R646 B.n112 B.n111 163.367
R647 B.n116 B.n115 163.367
R648 B.n120 B.n119 163.367
R649 B.n124 B.n123 163.367
R650 B.n128 B.n127 163.367
R651 B.n132 B.n131 163.367
R652 B.n136 B.n135 163.367
R653 B.n140 B.n139 163.367
R654 B.n144 B.n143 163.367
R655 B.n148 B.n147 163.367
R656 B.n152 B.n151 163.367
R657 B.n156 B.n155 163.367
R658 B.n160 B.n159 163.367
R659 B.n164 B.n163 163.367
R660 B.n168 B.n167 163.367
R661 B.n172 B.n171 163.367
R662 B.n176 B.n175 163.367
R663 B.n180 B.n179 163.367
R664 B.n184 B.n183 163.367
R665 B.n188 B.n187 163.367
R666 B.n192 B.n191 163.367
R667 B.n196 B.n195 163.367
R668 B.n200 B.n199 163.367
R669 B.n204 B.n203 163.367
R670 B.n208 B.n207 163.367
R671 B.n212 B.n211 163.367
R672 B.n217 B.n216 163.367
R673 B.n221 B.n220 163.367
R674 B.n225 B.n224 163.367
R675 B.n229 B.n228 163.367
R676 B.n233 B.n232 163.367
R677 B.n237 B.n236 163.367
R678 B.n241 B.n240 163.367
R679 B.n245 B.n244 163.367
R680 B.n249 B.n248 163.367
R681 B.n253 B.n252 163.367
R682 B.n257 B.n256 163.367
R683 B.n261 B.n260 163.367
R684 B.n265 B.n264 163.367
R685 B.n269 B.n268 163.367
R686 B.n273 B.n272 163.367
R687 B.n277 B.n276 163.367
R688 B.n281 B.n280 163.367
R689 B.n285 B.n284 163.367
R690 B.n289 B.n288 163.367
R691 B.n293 B.n292 163.367
R692 B.n297 B.n296 163.367
R693 B.n301 B.n300 163.367
R694 B.n305 B.n304 163.367
R695 B.n309 B.n308 163.367
R696 B.n313 B.n312 163.367
R697 B.n317 B.n316 163.367
R698 B.n321 B.n320 163.367
R699 B.n325 B.n324 163.367
R700 B.n329 B.n328 163.367
R701 B.n333 B.n332 163.367
R702 B.n337 B.n336 163.367
R703 B.n341 B.n340 163.367
R704 B.n345 B.n344 163.367
R705 B.n753 B.n90 163.367
R706 B.n439 B.t11 80.6407
R707 B.n91 B.t6 80.6407
R708 B.n436 B.t14 80.617
R709 B.n94 B.t16 80.617
R710 B.n690 B.n689 71.676
R711 B.n684 B.n373 71.676
R712 B.n681 B.n374 71.676
R713 B.n677 B.n375 71.676
R714 B.n673 B.n376 71.676
R715 B.n669 B.n377 71.676
R716 B.n665 B.n378 71.676
R717 B.n661 B.n379 71.676
R718 B.n657 B.n380 71.676
R719 B.n653 B.n381 71.676
R720 B.n649 B.n382 71.676
R721 B.n645 B.n383 71.676
R722 B.n641 B.n384 71.676
R723 B.n637 B.n385 71.676
R724 B.n633 B.n386 71.676
R725 B.n629 B.n387 71.676
R726 B.n625 B.n388 71.676
R727 B.n621 B.n389 71.676
R728 B.n617 B.n390 71.676
R729 B.n613 B.n391 71.676
R730 B.n609 B.n392 71.676
R731 B.n605 B.n393 71.676
R732 B.n601 B.n394 71.676
R733 B.n597 B.n395 71.676
R734 B.n593 B.n396 71.676
R735 B.n589 B.n397 71.676
R736 B.n585 B.n398 71.676
R737 B.n581 B.n399 71.676
R738 B.n577 B.n400 71.676
R739 B.n573 B.n401 71.676
R740 B.n569 B.n402 71.676
R741 B.n565 B.n403 71.676
R742 B.n561 B.n404 71.676
R743 B.n557 B.n405 71.676
R744 B.n552 B.n406 71.676
R745 B.n548 B.n407 71.676
R746 B.n544 B.n408 71.676
R747 B.n540 B.n409 71.676
R748 B.n536 B.n410 71.676
R749 B.n532 B.n411 71.676
R750 B.n528 B.n412 71.676
R751 B.n524 B.n413 71.676
R752 B.n520 B.n414 71.676
R753 B.n516 B.n415 71.676
R754 B.n512 B.n416 71.676
R755 B.n508 B.n417 71.676
R756 B.n504 B.n418 71.676
R757 B.n500 B.n419 71.676
R758 B.n496 B.n420 71.676
R759 B.n492 B.n421 71.676
R760 B.n488 B.n422 71.676
R761 B.n484 B.n423 71.676
R762 B.n480 B.n424 71.676
R763 B.n476 B.n425 71.676
R764 B.n472 B.n426 71.676
R765 B.n468 B.n427 71.676
R766 B.n464 B.n428 71.676
R767 B.n460 B.n429 71.676
R768 B.n456 B.n430 71.676
R769 B.n452 B.n431 71.676
R770 B.n448 B.n432 71.676
R771 B.n444 B.n433 71.676
R772 B.n692 B.n372 71.676
R773 B.n96 B.n27 71.676
R774 B.n100 B.n28 71.676
R775 B.n104 B.n29 71.676
R776 B.n108 B.n30 71.676
R777 B.n112 B.n31 71.676
R778 B.n116 B.n32 71.676
R779 B.n120 B.n33 71.676
R780 B.n124 B.n34 71.676
R781 B.n128 B.n35 71.676
R782 B.n132 B.n36 71.676
R783 B.n136 B.n37 71.676
R784 B.n140 B.n38 71.676
R785 B.n144 B.n39 71.676
R786 B.n148 B.n40 71.676
R787 B.n152 B.n41 71.676
R788 B.n156 B.n42 71.676
R789 B.n160 B.n43 71.676
R790 B.n164 B.n44 71.676
R791 B.n168 B.n45 71.676
R792 B.n172 B.n46 71.676
R793 B.n176 B.n47 71.676
R794 B.n180 B.n48 71.676
R795 B.n184 B.n49 71.676
R796 B.n188 B.n50 71.676
R797 B.n192 B.n51 71.676
R798 B.n196 B.n52 71.676
R799 B.n200 B.n53 71.676
R800 B.n204 B.n54 71.676
R801 B.n208 B.n55 71.676
R802 B.n212 B.n56 71.676
R803 B.n217 B.n57 71.676
R804 B.n221 B.n58 71.676
R805 B.n225 B.n59 71.676
R806 B.n229 B.n60 71.676
R807 B.n233 B.n61 71.676
R808 B.n237 B.n62 71.676
R809 B.n241 B.n63 71.676
R810 B.n245 B.n64 71.676
R811 B.n249 B.n65 71.676
R812 B.n253 B.n66 71.676
R813 B.n257 B.n67 71.676
R814 B.n261 B.n68 71.676
R815 B.n265 B.n69 71.676
R816 B.n269 B.n70 71.676
R817 B.n273 B.n71 71.676
R818 B.n277 B.n72 71.676
R819 B.n281 B.n73 71.676
R820 B.n285 B.n74 71.676
R821 B.n289 B.n75 71.676
R822 B.n293 B.n76 71.676
R823 B.n297 B.n77 71.676
R824 B.n301 B.n78 71.676
R825 B.n305 B.n79 71.676
R826 B.n309 B.n80 71.676
R827 B.n313 B.n81 71.676
R828 B.n317 B.n82 71.676
R829 B.n321 B.n83 71.676
R830 B.n325 B.n84 71.676
R831 B.n329 B.n85 71.676
R832 B.n333 B.n86 71.676
R833 B.n337 B.n87 71.676
R834 B.n341 B.n88 71.676
R835 B.n345 B.n89 71.676
R836 B.n90 B.n89 71.676
R837 B.n344 B.n88 71.676
R838 B.n340 B.n87 71.676
R839 B.n336 B.n86 71.676
R840 B.n332 B.n85 71.676
R841 B.n328 B.n84 71.676
R842 B.n324 B.n83 71.676
R843 B.n320 B.n82 71.676
R844 B.n316 B.n81 71.676
R845 B.n312 B.n80 71.676
R846 B.n308 B.n79 71.676
R847 B.n304 B.n78 71.676
R848 B.n300 B.n77 71.676
R849 B.n296 B.n76 71.676
R850 B.n292 B.n75 71.676
R851 B.n288 B.n74 71.676
R852 B.n284 B.n73 71.676
R853 B.n280 B.n72 71.676
R854 B.n276 B.n71 71.676
R855 B.n272 B.n70 71.676
R856 B.n268 B.n69 71.676
R857 B.n264 B.n68 71.676
R858 B.n260 B.n67 71.676
R859 B.n256 B.n66 71.676
R860 B.n252 B.n65 71.676
R861 B.n248 B.n64 71.676
R862 B.n244 B.n63 71.676
R863 B.n240 B.n62 71.676
R864 B.n236 B.n61 71.676
R865 B.n232 B.n60 71.676
R866 B.n228 B.n59 71.676
R867 B.n224 B.n58 71.676
R868 B.n220 B.n57 71.676
R869 B.n216 B.n56 71.676
R870 B.n211 B.n55 71.676
R871 B.n207 B.n54 71.676
R872 B.n203 B.n53 71.676
R873 B.n199 B.n52 71.676
R874 B.n195 B.n51 71.676
R875 B.n191 B.n50 71.676
R876 B.n187 B.n49 71.676
R877 B.n183 B.n48 71.676
R878 B.n179 B.n47 71.676
R879 B.n175 B.n46 71.676
R880 B.n171 B.n45 71.676
R881 B.n167 B.n44 71.676
R882 B.n163 B.n43 71.676
R883 B.n159 B.n42 71.676
R884 B.n155 B.n41 71.676
R885 B.n151 B.n40 71.676
R886 B.n147 B.n39 71.676
R887 B.n143 B.n38 71.676
R888 B.n139 B.n37 71.676
R889 B.n135 B.n36 71.676
R890 B.n131 B.n35 71.676
R891 B.n127 B.n34 71.676
R892 B.n123 B.n33 71.676
R893 B.n119 B.n32 71.676
R894 B.n115 B.n31 71.676
R895 B.n111 B.n30 71.676
R896 B.n107 B.n29 71.676
R897 B.n103 B.n28 71.676
R898 B.n99 B.n27 71.676
R899 B.n690 B.n435 71.676
R900 B.n682 B.n373 71.676
R901 B.n678 B.n374 71.676
R902 B.n674 B.n375 71.676
R903 B.n670 B.n376 71.676
R904 B.n666 B.n377 71.676
R905 B.n662 B.n378 71.676
R906 B.n658 B.n379 71.676
R907 B.n654 B.n380 71.676
R908 B.n650 B.n381 71.676
R909 B.n646 B.n382 71.676
R910 B.n642 B.n383 71.676
R911 B.n638 B.n384 71.676
R912 B.n634 B.n385 71.676
R913 B.n630 B.n386 71.676
R914 B.n626 B.n387 71.676
R915 B.n622 B.n388 71.676
R916 B.n618 B.n389 71.676
R917 B.n614 B.n390 71.676
R918 B.n610 B.n391 71.676
R919 B.n606 B.n392 71.676
R920 B.n602 B.n393 71.676
R921 B.n598 B.n394 71.676
R922 B.n594 B.n395 71.676
R923 B.n590 B.n396 71.676
R924 B.n586 B.n397 71.676
R925 B.n582 B.n398 71.676
R926 B.n578 B.n399 71.676
R927 B.n574 B.n400 71.676
R928 B.n570 B.n401 71.676
R929 B.n566 B.n402 71.676
R930 B.n562 B.n403 71.676
R931 B.n558 B.n404 71.676
R932 B.n553 B.n405 71.676
R933 B.n549 B.n406 71.676
R934 B.n545 B.n407 71.676
R935 B.n541 B.n408 71.676
R936 B.n537 B.n409 71.676
R937 B.n533 B.n410 71.676
R938 B.n529 B.n411 71.676
R939 B.n525 B.n412 71.676
R940 B.n521 B.n413 71.676
R941 B.n517 B.n414 71.676
R942 B.n513 B.n415 71.676
R943 B.n509 B.n416 71.676
R944 B.n505 B.n417 71.676
R945 B.n501 B.n418 71.676
R946 B.n497 B.n419 71.676
R947 B.n493 B.n420 71.676
R948 B.n489 B.n421 71.676
R949 B.n485 B.n422 71.676
R950 B.n481 B.n423 71.676
R951 B.n477 B.n424 71.676
R952 B.n473 B.n425 71.676
R953 B.n469 B.n426 71.676
R954 B.n465 B.n427 71.676
R955 B.n461 B.n428 71.676
R956 B.n457 B.n429 71.676
R957 B.n453 B.n430 71.676
R958 B.n449 B.n431 71.676
R959 B.n445 B.n432 71.676
R960 B.n441 B.n433 71.676
R961 B.n693 B.n692 71.676
R962 B.n440 B.t10 70.168
R963 B.n92 B.t7 70.168
R964 B.n437 B.t13 70.1442
R965 B.n95 B.t17 70.1442
R966 B.n555 B.n440 59.5399
R967 B.n438 B.n437 59.5399
R968 B.n214 B.n95 59.5399
R969 B.n93 B.n92 59.5399
R970 B.n691 B.n369 54.7032
R971 B.n755 B.n754 54.7032
R972 B.n698 B.n369 32.3464
R973 B.n698 B.n364 32.3464
R974 B.n704 B.n364 32.3464
R975 B.n704 B.n365 32.3464
R976 B.n710 B.n357 32.3464
R977 B.n716 B.n357 32.3464
R978 B.n716 B.n353 32.3464
R979 B.n724 B.n353 32.3464
R980 B.n730 B.n4 32.3464
R981 B.n780 B.n4 32.3464
R982 B.n780 B.n779 32.3464
R983 B.n779 B.n778 32.3464
R984 B.n772 B.n771 32.3464
R985 B.n771 B.n770 32.3464
R986 B.n770 B.n14 32.3464
R987 B.n764 B.n14 32.3464
R988 B.n763 B.n762 32.3464
R989 B.n762 B.n21 32.3464
R990 B.n756 B.n21 32.3464
R991 B.n756 B.n755 32.3464
R992 B.n97 B.n23 32.3127
R993 B.n752 B.n751 32.3127
R994 B.n695 B.n694 32.3127
R995 B.n688 B.n367 32.3127
R996 B.t3 B.n723 31.8708
R997 B.n737 B.t0 31.8708
R998 B.n710 B.t9 25.2113
R999 B.n764 B.t5 25.2113
R1000 B.n723 B.t2 19.5032
R1001 B.n737 B.t1 19.5032
R1002 B B.n782 18.0485
R1003 B.n730 B.t2 12.8437
R1004 B.n778 B.t1 12.8437
R1005 B.n98 B.n97 10.6151
R1006 B.n101 B.n98 10.6151
R1007 B.n102 B.n101 10.6151
R1008 B.n105 B.n102 10.6151
R1009 B.n106 B.n105 10.6151
R1010 B.n109 B.n106 10.6151
R1011 B.n110 B.n109 10.6151
R1012 B.n113 B.n110 10.6151
R1013 B.n114 B.n113 10.6151
R1014 B.n117 B.n114 10.6151
R1015 B.n118 B.n117 10.6151
R1016 B.n121 B.n118 10.6151
R1017 B.n122 B.n121 10.6151
R1018 B.n125 B.n122 10.6151
R1019 B.n126 B.n125 10.6151
R1020 B.n129 B.n126 10.6151
R1021 B.n130 B.n129 10.6151
R1022 B.n133 B.n130 10.6151
R1023 B.n134 B.n133 10.6151
R1024 B.n137 B.n134 10.6151
R1025 B.n138 B.n137 10.6151
R1026 B.n141 B.n138 10.6151
R1027 B.n142 B.n141 10.6151
R1028 B.n145 B.n142 10.6151
R1029 B.n146 B.n145 10.6151
R1030 B.n149 B.n146 10.6151
R1031 B.n150 B.n149 10.6151
R1032 B.n153 B.n150 10.6151
R1033 B.n154 B.n153 10.6151
R1034 B.n157 B.n154 10.6151
R1035 B.n158 B.n157 10.6151
R1036 B.n161 B.n158 10.6151
R1037 B.n162 B.n161 10.6151
R1038 B.n165 B.n162 10.6151
R1039 B.n166 B.n165 10.6151
R1040 B.n169 B.n166 10.6151
R1041 B.n170 B.n169 10.6151
R1042 B.n173 B.n170 10.6151
R1043 B.n174 B.n173 10.6151
R1044 B.n177 B.n174 10.6151
R1045 B.n178 B.n177 10.6151
R1046 B.n181 B.n178 10.6151
R1047 B.n182 B.n181 10.6151
R1048 B.n185 B.n182 10.6151
R1049 B.n186 B.n185 10.6151
R1050 B.n189 B.n186 10.6151
R1051 B.n190 B.n189 10.6151
R1052 B.n193 B.n190 10.6151
R1053 B.n194 B.n193 10.6151
R1054 B.n197 B.n194 10.6151
R1055 B.n198 B.n197 10.6151
R1056 B.n201 B.n198 10.6151
R1057 B.n202 B.n201 10.6151
R1058 B.n205 B.n202 10.6151
R1059 B.n206 B.n205 10.6151
R1060 B.n209 B.n206 10.6151
R1061 B.n210 B.n209 10.6151
R1062 B.n213 B.n210 10.6151
R1063 B.n218 B.n215 10.6151
R1064 B.n219 B.n218 10.6151
R1065 B.n222 B.n219 10.6151
R1066 B.n223 B.n222 10.6151
R1067 B.n226 B.n223 10.6151
R1068 B.n227 B.n226 10.6151
R1069 B.n230 B.n227 10.6151
R1070 B.n231 B.n230 10.6151
R1071 B.n235 B.n234 10.6151
R1072 B.n238 B.n235 10.6151
R1073 B.n239 B.n238 10.6151
R1074 B.n242 B.n239 10.6151
R1075 B.n243 B.n242 10.6151
R1076 B.n246 B.n243 10.6151
R1077 B.n247 B.n246 10.6151
R1078 B.n250 B.n247 10.6151
R1079 B.n251 B.n250 10.6151
R1080 B.n254 B.n251 10.6151
R1081 B.n255 B.n254 10.6151
R1082 B.n258 B.n255 10.6151
R1083 B.n259 B.n258 10.6151
R1084 B.n262 B.n259 10.6151
R1085 B.n263 B.n262 10.6151
R1086 B.n266 B.n263 10.6151
R1087 B.n267 B.n266 10.6151
R1088 B.n270 B.n267 10.6151
R1089 B.n271 B.n270 10.6151
R1090 B.n274 B.n271 10.6151
R1091 B.n275 B.n274 10.6151
R1092 B.n278 B.n275 10.6151
R1093 B.n279 B.n278 10.6151
R1094 B.n282 B.n279 10.6151
R1095 B.n283 B.n282 10.6151
R1096 B.n286 B.n283 10.6151
R1097 B.n287 B.n286 10.6151
R1098 B.n290 B.n287 10.6151
R1099 B.n291 B.n290 10.6151
R1100 B.n294 B.n291 10.6151
R1101 B.n295 B.n294 10.6151
R1102 B.n298 B.n295 10.6151
R1103 B.n299 B.n298 10.6151
R1104 B.n302 B.n299 10.6151
R1105 B.n303 B.n302 10.6151
R1106 B.n306 B.n303 10.6151
R1107 B.n307 B.n306 10.6151
R1108 B.n310 B.n307 10.6151
R1109 B.n311 B.n310 10.6151
R1110 B.n314 B.n311 10.6151
R1111 B.n315 B.n314 10.6151
R1112 B.n318 B.n315 10.6151
R1113 B.n319 B.n318 10.6151
R1114 B.n322 B.n319 10.6151
R1115 B.n323 B.n322 10.6151
R1116 B.n326 B.n323 10.6151
R1117 B.n327 B.n326 10.6151
R1118 B.n330 B.n327 10.6151
R1119 B.n331 B.n330 10.6151
R1120 B.n334 B.n331 10.6151
R1121 B.n335 B.n334 10.6151
R1122 B.n338 B.n335 10.6151
R1123 B.n339 B.n338 10.6151
R1124 B.n342 B.n339 10.6151
R1125 B.n343 B.n342 10.6151
R1126 B.n346 B.n343 10.6151
R1127 B.n347 B.n346 10.6151
R1128 B.n752 B.n347 10.6151
R1129 B.n696 B.n695 10.6151
R1130 B.n696 B.n362 10.6151
R1131 B.n706 B.n362 10.6151
R1132 B.n707 B.n706 10.6151
R1133 B.n708 B.n707 10.6151
R1134 B.n708 B.n355 10.6151
R1135 B.n718 B.n355 10.6151
R1136 B.n719 B.n718 10.6151
R1137 B.n721 B.n719 10.6151
R1138 B.n721 B.n720 10.6151
R1139 B.n720 B.n348 10.6151
R1140 B.n733 B.n348 10.6151
R1141 B.n734 B.n733 10.6151
R1142 B.n735 B.n734 10.6151
R1143 B.n736 B.n735 10.6151
R1144 B.n739 B.n736 10.6151
R1145 B.n740 B.n739 10.6151
R1146 B.n741 B.n740 10.6151
R1147 B.n742 B.n741 10.6151
R1148 B.n744 B.n742 10.6151
R1149 B.n745 B.n744 10.6151
R1150 B.n746 B.n745 10.6151
R1151 B.n747 B.n746 10.6151
R1152 B.n749 B.n747 10.6151
R1153 B.n750 B.n749 10.6151
R1154 B.n751 B.n750 10.6151
R1155 B.n688 B.n687 10.6151
R1156 B.n687 B.n686 10.6151
R1157 B.n686 B.n685 10.6151
R1158 B.n685 B.n683 10.6151
R1159 B.n683 B.n680 10.6151
R1160 B.n680 B.n679 10.6151
R1161 B.n679 B.n676 10.6151
R1162 B.n676 B.n675 10.6151
R1163 B.n675 B.n672 10.6151
R1164 B.n672 B.n671 10.6151
R1165 B.n671 B.n668 10.6151
R1166 B.n668 B.n667 10.6151
R1167 B.n667 B.n664 10.6151
R1168 B.n664 B.n663 10.6151
R1169 B.n663 B.n660 10.6151
R1170 B.n660 B.n659 10.6151
R1171 B.n659 B.n656 10.6151
R1172 B.n656 B.n655 10.6151
R1173 B.n655 B.n652 10.6151
R1174 B.n652 B.n651 10.6151
R1175 B.n651 B.n648 10.6151
R1176 B.n648 B.n647 10.6151
R1177 B.n647 B.n644 10.6151
R1178 B.n644 B.n643 10.6151
R1179 B.n643 B.n640 10.6151
R1180 B.n640 B.n639 10.6151
R1181 B.n639 B.n636 10.6151
R1182 B.n636 B.n635 10.6151
R1183 B.n635 B.n632 10.6151
R1184 B.n632 B.n631 10.6151
R1185 B.n631 B.n628 10.6151
R1186 B.n628 B.n627 10.6151
R1187 B.n627 B.n624 10.6151
R1188 B.n624 B.n623 10.6151
R1189 B.n623 B.n620 10.6151
R1190 B.n620 B.n619 10.6151
R1191 B.n619 B.n616 10.6151
R1192 B.n616 B.n615 10.6151
R1193 B.n615 B.n612 10.6151
R1194 B.n612 B.n611 10.6151
R1195 B.n611 B.n608 10.6151
R1196 B.n608 B.n607 10.6151
R1197 B.n607 B.n604 10.6151
R1198 B.n604 B.n603 10.6151
R1199 B.n603 B.n600 10.6151
R1200 B.n600 B.n599 10.6151
R1201 B.n599 B.n596 10.6151
R1202 B.n596 B.n595 10.6151
R1203 B.n595 B.n592 10.6151
R1204 B.n592 B.n591 10.6151
R1205 B.n591 B.n588 10.6151
R1206 B.n588 B.n587 10.6151
R1207 B.n587 B.n584 10.6151
R1208 B.n584 B.n583 10.6151
R1209 B.n583 B.n580 10.6151
R1210 B.n580 B.n579 10.6151
R1211 B.n579 B.n576 10.6151
R1212 B.n576 B.n575 10.6151
R1213 B.n572 B.n571 10.6151
R1214 B.n571 B.n568 10.6151
R1215 B.n568 B.n567 10.6151
R1216 B.n567 B.n564 10.6151
R1217 B.n564 B.n563 10.6151
R1218 B.n563 B.n560 10.6151
R1219 B.n560 B.n559 10.6151
R1220 B.n559 B.n556 10.6151
R1221 B.n554 B.n551 10.6151
R1222 B.n551 B.n550 10.6151
R1223 B.n550 B.n547 10.6151
R1224 B.n547 B.n546 10.6151
R1225 B.n546 B.n543 10.6151
R1226 B.n543 B.n542 10.6151
R1227 B.n542 B.n539 10.6151
R1228 B.n539 B.n538 10.6151
R1229 B.n538 B.n535 10.6151
R1230 B.n535 B.n534 10.6151
R1231 B.n534 B.n531 10.6151
R1232 B.n531 B.n530 10.6151
R1233 B.n530 B.n527 10.6151
R1234 B.n527 B.n526 10.6151
R1235 B.n526 B.n523 10.6151
R1236 B.n523 B.n522 10.6151
R1237 B.n522 B.n519 10.6151
R1238 B.n519 B.n518 10.6151
R1239 B.n518 B.n515 10.6151
R1240 B.n515 B.n514 10.6151
R1241 B.n514 B.n511 10.6151
R1242 B.n511 B.n510 10.6151
R1243 B.n510 B.n507 10.6151
R1244 B.n507 B.n506 10.6151
R1245 B.n506 B.n503 10.6151
R1246 B.n503 B.n502 10.6151
R1247 B.n502 B.n499 10.6151
R1248 B.n499 B.n498 10.6151
R1249 B.n498 B.n495 10.6151
R1250 B.n495 B.n494 10.6151
R1251 B.n494 B.n491 10.6151
R1252 B.n491 B.n490 10.6151
R1253 B.n490 B.n487 10.6151
R1254 B.n487 B.n486 10.6151
R1255 B.n486 B.n483 10.6151
R1256 B.n483 B.n482 10.6151
R1257 B.n482 B.n479 10.6151
R1258 B.n479 B.n478 10.6151
R1259 B.n478 B.n475 10.6151
R1260 B.n475 B.n474 10.6151
R1261 B.n474 B.n471 10.6151
R1262 B.n471 B.n470 10.6151
R1263 B.n470 B.n467 10.6151
R1264 B.n467 B.n466 10.6151
R1265 B.n466 B.n463 10.6151
R1266 B.n463 B.n462 10.6151
R1267 B.n462 B.n459 10.6151
R1268 B.n459 B.n458 10.6151
R1269 B.n458 B.n455 10.6151
R1270 B.n455 B.n454 10.6151
R1271 B.n454 B.n451 10.6151
R1272 B.n451 B.n450 10.6151
R1273 B.n450 B.n447 10.6151
R1274 B.n447 B.n446 10.6151
R1275 B.n446 B.n443 10.6151
R1276 B.n443 B.n442 10.6151
R1277 B.n442 B.n371 10.6151
R1278 B.n694 B.n371 10.6151
R1279 B.n700 B.n367 10.6151
R1280 B.n701 B.n700 10.6151
R1281 B.n702 B.n701 10.6151
R1282 B.n702 B.n359 10.6151
R1283 B.n712 B.n359 10.6151
R1284 B.n713 B.n712 10.6151
R1285 B.n714 B.n713 10.6151
R1286 B.n714 B.n351 10.6151
R1287 B.n726 B.n351 10.6151
R1288 B.n727 B.n726 10.6151
R1289 B.n728 B.n727 10.6151
R1290 B.n728 B.n0 10.6151
R1291 B.n776 B.n1 10.6151
R1292 B.n776 B.n775 10.6151
R1293 B.n775 B.n774 10.6151
R1294 B.n774 B.n9 10.6151
R1295 B.n768 B.n9 10.6151
R1296 B.n768 B.n767 10.6151
R1297 B.n767 B.n766 10.6151
R1298 B.n766 B.n16 10.6151
R1299 B.n760 B.n16 10.6151
R1300 B.n760 B.n759 10.6151
R1301 B.n759 B.n758 10.6151
R1302 B.n758 B.n23 10.6151
R1303 B.n440 B.n439 10.4732
R1304 B.n437 B.n436 10.4732
R1305 B.n95 B.n94 10.4732
R1306 B.n92 B.n91 10.4732
R1307 B.n215 B.n214 7.18099
R1308 B.n231 B.n93 7.18099
R1309 B.n572 B.n438 7.18099
R1310 B.n556 B.n555 7.18099
R1311 B.n365 B.t9 7.13564
R1312 B.t5 B.n763 7.13564
R1313 B.n214 B.n213 3.43465
R1314 B.n234 B.n93 3.43465
R1315 B.n575 B.n438 3.43465
R1316 B.n555 B.n554 3.43465
R1317 B.n782 B.n0 2.81026
R1318 B.n782 B.n1 2.81026
R1319 B.n724 B.t3 0.476176
R1320 B.n772 B.t0 0.476176
R1321 VP.n1 VP.t0 2235.98
R1322 VP.n1 VP.t3 2235.98
R1323 VP.n0 VP.t1 2235.98
R1324 VP.n0 VP.t2 2235.98
R1325 VP.n2 VP.n0 204.665
R1326 VP.n2 VP.n1 161.3
R1327 VP VP.n2 0.0516364
R1328 VDD1 VDD1.n1 100.719
R1329 VDD1 VDD1.n0 59.7523
R1330 VDD1.n0 VDD1.t2 1.11099
R1331 VDD1.n0 VDD1.t1 1.11099
R1332 VDD1.n1 VDD1.t0 1.11099
R1333 VDD1.n1 VDD1.t3 1.11099
C0 VDD2 VP 0.243364f
C1 VDD1 VN 0.147979f
C2 VDD2 VN 2.46973f
C3 VDD1 VTAIL 15.4249f
C4 VDD2 VTAIL 15.463099f
C5 VN VP 5.54599f
C6 VDD2 VDD1 0.460209f
C7 VTAIL VP 1.64946f
C8 VTAIL VN 1.63535f
C9 VDD1 VP 2.56499f
C10 VDD2 B 2.884251f
C11 VDD1 B 8.35233f
C12 VTAIL B 11.014419f
C13 VN B 8.640161f
C14 VP B 4.256843f
C15 VDD1.t2 B 0.518009f
C16 VDD1.t1 B 0.518009f
C17 VDD1.n0 B 4.71531f
C18 VDD1.t0 B 0.518009f
C19 VDD1.t3 B 0.518009f
C20 VDD1.n1 B 5.81025f
C21 VP.t1 B 0.584334f
C22 VP.t2 B 0.584334f
C23 VP.n0 B 0.965984f
C24 VP.t3 B 0.584334f
C25 VP.t0 B 0.584334f
C26 VP.n1 B 0.457263f
C27 VP.n2 B 4.31857f
C28 VDD2.t0 B 0.521946f
C29 VDD2.t2 B 0.521946f
C30 VDD2.n0 B 5.81588f
C31 VDD2.t1 B 0.521946f
C32 VDD2.t3 B 0.521946f
C33 VDD2.n1 B 4.75077f
C34 VDD2.n2 B 5.28203f
C35 VTAIL.t5 B 2.96255f
C36 VTAIL.n0 B 0.303912f
C37 VTAIL.t2 B 2.96255f
C38 VTAIL.n1 B 0.314344f
C39 VTAIL.t3 B 2.96255f
C40 VTAIL.n2 B 1.48557f
C41 VTAIL.t7 B 2.96255f
C42 VTAIL.n3 B 1.48556f
C43 VTAIL.t6 B 2.96255f
C44 VTAIL.n4 B 0.31434f
C45 VTAIL.t1 B 2.96255f
C46 VTAIL.n5 B 0.31434f
C47 VTAIL.t0 B 2.96255f
C48 VTAIL.n6 B 1.48557f
C49 VTAIL.t4 B 2.96255f
C50 VTAIL.n7 B 1.46818f
C51 VN.t3 B 0.571664f
C52 VN.t1 B 0.571664f
C53 VN.n0 B 0.447364f
C54 VN.t2 B 0.571664f
C55 VN.t0 B 0.571664f
C56 VN.n1 B 0.955997f
.ends

