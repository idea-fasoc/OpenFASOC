* NGSPICE file created from diff_pair_sample_1041.ext - technology: sky130A

.subckt diff_pair_sample_1041 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X1 VTAIL.t4 VP.t0 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X2 VTAIL.t6 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X3 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=0 ps=0 w=6.56 l=0.17
X4 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X5 VDD1.t6 VP.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=2.5584 ps=13.9 w=6.56 l=0.17
X6 VTAIL.t8 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X7 VTAIL.t18 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X8 VDD2.t7 VN.t2 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=2.5584 ps=13.9 w=6.56 l=0.17
X9 VDD1.t4 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=2.5584 ps=13.9 w=6.56 l=0.17
X10 VDD2.t6 VN.t3 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=1.0824 ps=6.89 w=6.56 l=0.17
X11 VTAIL.t19 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X12 VDD1.t3 VP.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=1.0824 ps=6.89 w=6.56 l=0.17
X13 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=0 ps=0 w=6.56 l=0.17
X14 VDD2.t4 VN.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X15 VTAIL.t7 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X16 VTAIL.t11 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X17 VDD2.t2 VN.t7 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=2.5584 ps=13.9 w=6.56 l=0.17
X18 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=0 ps=0 w=6.56 l=0.17
X19 VDD2.t1 VN.t8 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=1.0824 ps=6.89 w=6.56 l=0.17
X20 VTAIL.t10 VN.t9 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=0 ps=0 w=6.56 l=0.17
X22 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0824 pd=6.89 as=1.0824 ps=6.89 w=6.56 l=0.17
X23 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5584 pd=13.9 as=1.0824 ps=6.89 w=6.56 l=0.17
R0 VN.n8 VN.t2 1150.79
R1 VN.n2 VN.t8 1150.79
R2 VN.n18 VN.t3 1150.79
R3 VN.n12 VN.t7 1150.79
R4 VN.n7 VN.t4 1114.27
R5 VN.n5 VN.t5 1114.27
R6 VN.n1 VN.t6 1114.27
R7 VN.n17 VN.t9 1114.27
R8 VN.n15 VN.t0 1114.27
R9 VN.n11 VN.t1 1114.27
R10 VN.n13 VN.n12 161.489
R11 VN.n3 VN.n2 161.489
R12 VN.n9 VN.n8 161.3
R13 VN.n19 VN.n18 161.3
R14 VN.n16 VN.n10 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n6 VN.n0 161.3
R17 VN.n4 VN.n3 161.3
R18 VN.n2 VN.n1 36.5157
R19 VN.n4 VN.n1 36.5157
R20 VN.n5 VN.n4 36.5157
R21 VN.n6 VN.n5 36.5157
R22 VN.n7 VN.n6 36.5157
R23 VN.n8 VN.n7 36.5157
R24 VN.n18 VN.n17 36.5157
R25 VN.n17 VN.n16 36.5157
R26 VN.n16 VN.n15 36.5157
R27 VN.n15 VN.n14 36.5157
R28 VN.n14 VN.n11 36.5157
R29 VN.n12 VN.n11 36.5157
R30 VN VN.n19 36.1766
R31 VN.n19 VN.n10 0.189894
R32 VN.n13 VN.n10 0.189894
R33 VN.n3 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VTAIL.n148 VTAIL.n147 289.615
R37 VTAIL.n34 VTAIL.n33 289.615
R38 VTAIL.n114 VTAIL.n113 289.615
R39 VTAIL.n76 VTAIL.n75 289.615
R40 VTAIL.n126 VTAIL.n125 185
R41 VTAIL.n131 VTAIL.n130 185
R42 VTAIL.n133 VTAIL.n132 185
R43 VTAIL.n122 VTAIL.n121 185
R44 VTAIL.n139 VTAIL.n138 185
R45 VTAIL.n141 VTAIL.n140 185
R46 VTAIL.n118 VTAIL.n117 185
R47 VTAIL.n147 VTAIL.n146 185
R48 VTAIL.n12 VTAIL.n11 185
R49 VTAIL.n17 VTAIL.n16 185
R50 VTAIL.n19 VTAIL.n18 185
R51 VTAIL.n8 VTAIL.n7 185
R52 VTAIL.n25 VTAIL.n24 185
R53 VTAIL.n27 VTAIL.n26 185
R54 VTAIL.n4 VTAIL.n3 185
R55 VTAIL.n33 VTAIL.n32 185
R56 VTAIL.n113 VTAIL.n112 185
R57 VTAIL.n84 VTAIL.n83 185
R58 VTAIL.n107 VTAIL.n106 185
R59 VTAIL.n105 VTAIL.n104 185
R60 VTAIL.n88 VTAIL.n87 185
R61 VTAIL.n99 VTAIL.n98 185
R62 VTAIL.n97 VTAIL.n96 185
R63 VTAIL.n92 VTAIL.n91 185
R64 VTAIL.n75 VTAIL.n74 185
R65 VTAIL.n46 VTAIL.n45 185
R66 VTAIL.n69 VTAIL.n68 185
R67 VTAIL.n67 VTAIL.n66 185
R68 VTAIL.n50 VTAIL.n49 185
R69 VTAIL.n61 VTAIL.n60 185
R70 VTAIL.n59 VTAIL.n58 185
R71 VTAIL.n54 VTAIL.n53 185
R72 VTAIL.n55 VTAIL.t15 149.525
R73 VTAIL.n127 VTAIL.t13 149.525
R74 VTAIL.n13 VTAIL.t3 149.525
R75 VTAIL.n93 VTAIL.t9 149.525
R76 VTAIL.n131 VTAIL.n125 104.615
R77 VTAIL.n132 VTAIL.n131 104.615
R78 VTAIL.n132 VTAIL.n121 104.615
R79 VTAIL.n139 VTAIL.n121 104.615
R80 VTAIL.n140 VTAIL.n139 104.615
R81 VTAIL.n140 VTAIL.n117 104.615
R82 VTAIL.n147 VTAIL.n117 104.615
R83 VTAIL.n17 VTAIL.n11 104.615
R84 VTAIL.n18 VTAIL.n17 104.615
R85 VTAIL.n18 VTAIL.n7 104.615
R86 VTAIL.n25 VTAIL.n7 104.615
R87 VTAIL.n26 VTAIL.n25 104.615
R88 VTAIL.n26 VTAIL.n3 104.615
R89 VTAIL.n33 VTAIL.n3 104.615
R90 VTAIL.n113 VTAIL.n83 104.615
R91 VTAIL.n106 VTAIL.n83 104.615
R92 VTAIL.n106 VTAIL.n105 104.615
R93 VTAIL.n105 VTAIL.n87 104.615
R94 VTAIL.n98 VTAIL.n87 104.615
R95 VTAIL.n98 VTAIL.n97 104.615
R96 VTAIL.n97 VTAIL.n91 104.615
R97 VTAIL.n75 VTAIL.n45 104.615
R98 VTAIL.n68 VTAIL.n45 104.615
R99 VTAIL.n68 VTAIL.n67 104.615
R100 VTAIL.n67 VTAIL.n49 104.615
R101 VTAIL.n60 VTAIL.n49 104.615
R102 VTAIL.n60 VTAIL.n59 104.615
R103 VTAIL.n59 VTAIL.n53 104.615
R104 VTAIL.n81 VTAIL.n80 52.614
R105 VTAIL.n79 VTAIL.n78 52.614
R106 VTAIL.n43 VTAIL.n42 52.614
R107 VTAIL.n41 VTAIL.n40 52.614
R108 VTAIL.n151 VTAIL.n150 52.613
R109 VTAIL.n1 VTAIL.n0 52.613
R110 VTAIL.n37 VTAIL.n36 52.613
R111 VTAIL.n39 VTAIL.n38 52.613
R112 VTAIL.t13 VTAIL.n125 52.3082
R113 VTAIL.t3 VTAIL.n11 52.3082
R114 VTAIL.t9 VTAIL.n91 52.3082
R115 VTAIL.t15 VTAIL.n53 52.3082
R116 VTAIL.n149 VTAIL.n148 35.6763
R117 VTAIL.n35 VTAIL.n34 35.6763
R118 VTAIL.n115 VTAIL.n114 35.6763
R119 VTAIL.n77 VTAIL.n76 35.6763
R120 VTAIL.n41 VTAIL.n39 18.8841
R121 VTAIL.n149 VTAIL.n115 18.4531
R122 VTAIL.n146 VTAIL.n116 12.8005
R123 VTAIL.n32 VTAIL.n2 12.8005
R124 VTAIL.n112 VTAIL.n82 12.8005
R125 VTAIL.n74 VTAIL.n44 12.8005
R126 VTAIL.n145 VTAIL.n118 12.0247
R127 VTAIL.n31 VTAIL.n4 12.0247
R128 VTAIL.n111 VTAIL.n84 12.0247
R129 VTAIL.n73 VTAIL.n46 12.0247
R130 VTAIL.n142 VTAIL.n141 11.249
R131 VTAIL.n28 VTAIL.n27 11.249
R132 VTAIL.n108 VTAIL.n107 11.249
R133 VTAIL.n70 VTAIL.n69 11.249
R134 VTAIL.n138 VTAIL.n120 10.4732
R135 VTAIL.n24 VTAIL.n6 10.4732
R136 VTAIL.n104 VTAIL.n86 10.4732
R137 VTAIL.n66 VTAIL.n48 10.4732
R138 VTAIL.n127 VTAIL.n126 10.2746
R139 VTAIL.n13 VTAIL.n12 10.2746
R140 VTAIL.n93 VTAIL.n92 10.2746
R141 VTAIL.n55 VTAIL.n54 10.2746
R142 VTAIL.n137 VTAIL.n122 9.69747
R143 VTAIL.n23 VTAIL.n8 9.69747
R144 VTAIL.n103 VTAIL.n88 9.69747
R145 VTAIL.n65 VTAIL.n50 9.69747
R146 VTAIL.n144 VTAIL.n116 9.45567
R147 VTAIL.n30 VTAIL.n2 9.45567
R148 VTAIL.n110 VTAIL.n82 9.45567
R149 VTAIL.n72 VTAIL.n44 9.45567
R150 VTAIL.n129 VTAIL.n128 9.3005
R151 VTAIL.n124 VTAIL.n123 9.3005
R152 VTAIL.n135 VTAIL.n134 9.3005
R153 VTAIL.n137 VTAIL.n136 9.3005
R154 VTAIL.n120 VTAIL.n119 9.3005
R155 VTAIL.n143 VTAIL.n142 9.3005
R156 VTAIL.n145 VTAIL.n144 9.3005
R157 VTAIL.n15 VTAIL.n14 9.3005
R158 VTAIL.n10 VTAIL.n9 9.3005
R159 VTAIL.n21 VTAIL.n20 9.3005
R160 VTAIL.n23 VTAIL.n22 9.3005
R161 VTAIL.n6 VTAIL.n5 9.3005
R162 VTAIL.n29 VTAIL.n28 9.3005
R163 VTAIL.n31 VTAIL.n30 9.3005
R164 VTAIL.n111 VTAIL.n110 9.3005
R165 VTAIL.n109 VTAIL.n108 9.3005
R166 VTAIL.n86 VTAIL.n85 9.3005
R167 VTAIL.n103 VTAIL.n102 9.3005
R168 VTAIL.n101 VTAIL.n100 9.3005
R169 VTAIL.n90 VTAIL.n89 9.3005
R170 VTAIL.n95 VTAIL.n94 9.3005
R171 VTAIL.n52 VTAIL.n51 9.3005
R172 VTAIL.n63 VTAIL.n62 9.3005
R173 VTAIL.n65 VTAIL.n64 9.3005
R174 VTAIL.n48 VTAIL.n47 9.3005
R175 VTAIL.n71 VTAIL.n70 9.3005
R176 VTAIL.n73 VTAIL.n72 9.3005
R177 VTAIL.n57 VTAIL.n56 9.3005
R178 VTAIL.n134 VTAIL.n133 8.92171
R179 VTAIL.n20 VTAIL.n19 8.92171
R180 VTAIL.n100 VTAIL.n99 8.92171
R181 VTAIL.n62 VTAIL.n61 8.92171
R182 VTAIL.n130 VTAIL.n124 8.14595
R183 VTAIL.n16 VTAIL.n10 8.14595
R184 VTAIL.n96 VTAIL.n90 8.14595
R185 VTAIL.n58 VTAIL.n52 8.14595
R186 VTAIL.n129 VTAIL.n126 7.3702
R187 VTAIL.n15 VTAIL.n12 7.3702
R188 VTAIL.n95 VTAIL.n92 7.3702
R189 VTAIL.n57 VTAIL.n54 7.3702
R190 VTAIL.n130 VTAIL.n129 5.81868
R191 VTAIL.n16 VTAIL.n15 5.81868
R192 VTAIL.n96 VTAIL.n95 5.81868
R193 VTAIL.n58 VTAIL.n57 5.81868
R194 VTAIL.n133 VTAIL.n124 5.04292
R195 VTAIL.n19 VTAIL.n10 5.04292
R196 VTAIL.n99 VTAIL.n90 5.04292
R197 VTAIL.n61 VTAIL.n52 5.04292
R198 VTAIL.n134 VTAIL.n122 4.26717
R199 VTAIL.n20 VTAIL.n8 4.26717
R200 VTAIL.n100 VTAIL.n88 4.26717
R201 VTAIL.n62 VTAIL.n50 4.26717
R202 VTAIL.n138 VTAIL.n137 3.49141
R203 VTAIL.n24 VTAIL.n23 3.49141
R204 VTAIL.n104 VTAIL.n103 3.49141
R205 VTAIL.n66 VTAIL.n65 3.49141
R206 VTAIL.n150 VTAIL.t14 3.01879
R207 VTAIL.n150 VTAIL.t19 3.01879
R208 VTAIL.n0 VTAIL.t12 3.01879
R209 VTAIL.n0 VTAIL.t11 3.01879
R210 VTAIL.n36 VTAIL.t2 3.01879
R211 VTAIL.n36 VTAIL.t8 3.01879
R212 VTAIL.n38 VTAIL.t1 3.01879
R213 VTAIL.n38 VTAIL.t4 3.01879
R214 VTAIL.n80 VTAIL.t0 3.01879
R215 VTAIL.n80 VTAIL.t7 3.01879
R216 VTAIL.n78 VTAIL.t5 3.01879
R217 VTAIL.n78 VTAIL.t6 3.01879
R218 VTAIL.n42 VTAIL.t16 3.01879
R219 VTAIL.n42 VTAIL.t18 3.01879
R220 VTAIL.n40 VTAIL.t17 3.01879
R221 VTAIL.n40 VTAIL.t10 3.01879
R222 VTAIL.n56 VTAIL.n55 2.84308
R223 VTAIL.n128 VTAIL.n127 2.84308
R224 VTAIL.n14 VTAIL.n13 2.84308
R225 VTAIL.n94 VTAIL.n93 2.84308
R226 VTAIL.n141 VTAIL.n120 2.71565
R227 VTAIL.n27 VTAIL.n6 2.71565
R228 VTAIL.n107 VTAIL.n86 2.71565
R229 VTAIL.n69 VTAIL.n48 2.71565
R230 VTAIL.n142 VTAIL.n118 1.93989
R231 VTAIL.n28 VTAIL.n4 1.93989
R232 VTAIL.n108 VTAIL.n84 1.93989
R233 VTAIL.n70 VTAIL.n46 1.93989
R234 VTAIL.n146 VTAIL.n145 1.16414
R235 VTAIL.n32 VTAIL.n31 1.16414
R236 VTAIL.n112 VTAIL.n111 1.16414
R237 VTAIL.n74 VTAIL.n73 1.16414
R238 VTAIL.n79 VTAIL.n77 0.685845
R239 VTAIL.n35 VTAIL.n1 0.685845
R240 VTAIL.n43 VTAIL.n41 0.431534
R241 VTAIL.n77 VTAIL.n43 0.431534
R242 VTAIL.n81 VTAIL.n79 0.431534
R243 VTAIL.n115 VTAIL.n81 0.431534
R244 VTAIL.n39 VTAIL.n37 0.431534
R245 VTAIL.n37 VTAIL.n35 0.431534
R246 VTAIL.n151 VTAIL.n149 0.431534
R247 VTAIL.n148 VTAIL.n116 0.388379
R248 VTAIL.n34 VTAIL.n2 0.388379
R249 VTAIL.n114 VTAIL.n82 0.388379
R250 VTAIL.n76 VTAIL.n44 0.388379
R251 VTAIL VTAIL.n1 0.381966
R252 VTAIL.n128 VTAIL.n123 0.155672
R253 VTAIL.n135 VTAIL.n123 0.155672
R254 VTAIL.n136 VTAIL.n135 0.155672
R255 VTAIL.n136 VTAIL.n119 0.155672
R256 VTAIL.n143 VTAIL.n119 0.155672
R257 VTAIL.n144 VTAIL.n143 0.155672
R258 VTAIL.n14 VTAIL.n9 0.155672
R259 VTAIL.n21 VTAIL.n9 0.155672
R260 VTAIL.n22 VTAIL.n21 0.155672
R261 VTAIL.n22 VTAIL.n5 0.155672
R262 VTAIL.n29 VTAIL.n5 0.155672
R263 VTAIL.n30 VTAIL.n29 0.155672
R264 VTAIL.n110 VTAIL.n109 0.155672
R265 VTAIL.n109 VTAIL.n85 0.155672
R266 VTAIL.n102 VTAIL.n85 0.155672
R267 VTAIL.n102 VTAIL.n101 0.155672
R268 VTAIL.n101 VTAIL.n89 0.155672
R269 VTAIL.n94 VTAIL.n89 0.155672
R270 VTAIL.n72 VTAIL.n71 0.155672
R271 VTAIL.n71 VTAIL.n47 0.155672
R272 VTAIL.n64 VTAIL.n47 0.155672
R273 VTAIL.n64 VTAIL.n63 0.155672
R274 VTAIL.n63 VTAIL.n51 0.155672
R275 VTAIL.n56 VTAIL.n51 0.155672
R276 VTAIL VTAIL.n151 0.050069
R277 VDD2.n69 VDD2.n68 289.615
R278 VDD2.n32 VDD2.n31 289.615
R279 VDD2.n68 VDD2.n67 185
R280 VDD2.n39 VDD2.n38 185
R281 VDD2.n62 VDD2.n61 185
R282 VDD2.n60 VDD2.n59 185
R283 VDD2.n43 VDD2.n42 185
R284 VDD2.n54 VDD2.n53 185
R285 VDD2.n52 VDD2.n51 185
R286 VDD2.n47 VDD2.n46 185
R287 VDD2.n10 VDD2.n9 185
R288 VDD2.n15 VDD2.n14 185
R289 VDD2.n17 VDD2.n16 185
R290 VDD2.n6 VDD2.n5 185
R291 VDD2.n23 VDD2.n22 185
R292 VDD2.n25 VDD2.n24 185
R293 VDD2.n2 VDD2.n1 185
R294 VDD2.n31 VDD2.n30 185
R295 VDD2.n48 VDD2.t6 149.525
R296 VDD2.n11 VDD2.t1 149.525
R297 VDD2.n68 VDD2.n38 104.615
R298 VDD2.n61 VDD2.n38 104.615
R299 VDD2.n61 VDD2.n60 104.615
R300 VDD2.n60 VDD2.n42 104.615
R301 VDD2.n53 VDD2.n42 104.615
R302 VDD2.n53 VDD2.n52 104.615
R303 VDD2.n52 VDD2.n46 104.615
R304 VDD2.n15 VDD2.n9 104.615
R305 VDD2.n16 VDD2.n15 104.615
R306 VDD2.n16 VDD2.n5 104.615
R307 VDD2.n23 VDD2.n5 104.615
R308 VDD2.n24 VDD2.n23 104.615
R309 VDD2.n24 VDD2.n1 104.615
R310 VDD2.n31 VDD2.n1 104.615
R311 VDD2.n36 VDD2.n35 69.5597
R312 VDD2 VDD2.n73 69.5568
R313 VDD2.n72 VDD2.n71 69.2928
R314 VDD2.n34 VDD2.n33 69.2918
R315 VDD2.n34 VDD2.n32 52.7861
R316 VDD2.n70 VDD2.n69 52.355
R317 VDD2.t6 VDD2.n46 52.3082
R318 VDD2.t1 VDD2.n9 52.3082
R319 VDD2.n70 VDD2.n36 31.4179
R320 VDD2.n67 VDD2.n37 12.8005
R321 VDD2.n30 VDD2.n0 12.8005
R322 VDD2.n66 VDD2.n39 12.0247
R323 VDD2.n29 VDD2.n2 12.0247
R324 VDD2.n63 VDD2.n62 11.249
R325 VDD2.n26 VDD2.n25 11.249
R326 VDD2.n59 VDD2.n41 10.4732
R327 VDD2.n22 VDD2.n4 10.4732
R328 VDD2.n48 VDD2.n47 10.2746
R329 VDD2.n11 VDD2.n10 10.2746
R330 VDD2.n58 VDD2.n43 9.69747
R331 VDD2.n21 VDD2.n6 9.69747
R332 VDD2.n65 VDD2.n37 9.45567
R333 VDD2.n28 VDD2.n0 9.45567
R334 VDD2.n45 VDD2.n44 9.3005
R335 VDD2.n56 VDD2.n55 9.3005
R336 VDD2.n58 VDD2.n57 9.3005
R337 VDD2.n41 VDD2.n40 9.3005
R338 VDD2.n64 VDD2.n63 9.3005
R339 VDD2.n66 VDD2.n65 9.3005
R340 VDD2.n50 VDD2.n49 9.3005
R341 VDD2.n13 VDD2.n12 9.3005
R342 VDD2.n8 VDD2.n7 9.3005
R343 VDD2.n19 VDD2.n18 9.3005
R344 VDD2.n21 VDD2.n20 9.3005
R345 VDD2.n4 VDD2.n3 9.3005
R346 VDD2.n27 VDD2.n26 9.3005
R347 VDD2.n29 VDD2.n28 9.3005
R348 VDD2.n55 VDD2.n54 8.92171
R349 VDD2.n18 VDD2.n17 8.92171
R350 VDD2.n51 VDD2.n45 8.14595
R351 VDD2.n14 VDD2.n8 8.14595
R352 VDD2.n50 VDD2.n47 7.3702
R353 VDD2.n13 VDD2.n10 7.3702
R354 VDD2.n51 VDD2.n50 5.81868
R355 VDD2.n14 VDD2.n13 5.81868
R356 VDD2.n54 VDD2.n45 5.04292
R357 VDD2.n17 VDD2.n8 5.04292
R358 VDD2.n55 VDD2.n43 4.26717
R359 VDD2.n18 VDD2.n6 4.26717
R360 VDD2.n59 VDD2.n58 3.49141
R361 VDD2.n22 VDD2.n21 3.49141
R362 VDD2.n73 VDD2.t8 3.01879
R363 VDD2.n73 VDD2.t2 3.01879
R364 VDD2.n71 VDD2.t0 3.01879
R365 VDD2.n71 VDD2.t9 3.01879
R366 VDD2.n35 VDD2.t5 3.01879
R367 VDD2.n35 VDD2.t7 3.01879
R368 VDD2.n33 VDD2.t3 3.01879
R369 VDD2.n33 VDD2.t4 3.01879
R370 VDD2.n49 VDD2.n48 2.84308
R371 VDD2.n12 VDD2.n11 2.84308
R372 VDD2.n62 VDD2.n41 2.71565
R373 VDD2.n25 VDD2.n4 2.71565
R374 VDD2.n63 VDD2.n39 1.93989
R375 VDD2.n26 VDD2.n2 1.93989
R376 VDD2.n67 VDD2.n66 1.16414
R377 VDD2.n30 VDD2.n29 1.16414
R378 VDD2.n72 VDD2.n70 0.431534
R379 VDD2.n69 VDD2.n37 0.388379
R380 VDD2.n32 VDD2.n0 0.388379
R381 VDD2 VDD2.n72 0.166448
R382 VDD2.n65 VDD2.n64 0.155672
R383 VDD2.n64 VDD2.n40 0.155672
R384 VDD2.n57 VDD2.n40 0.155672
R385 VDD2.n57 VDD2.n56 0.155672
R386 VDD2.n56 VDD2.n44 0.155672
R387 VDD2.n49 VDD2.n44 0.155672
R388 VDD2.n12 VDD2.n7 0.155672
R389 VDD2.n19 VDD2.n7 0.155672
R390 VDD2.n20 VDD2.n19 0.155672
R391 VDD2.n20 VDD2.n3 0.155672
R392 VDD2.n27 VDD2.n3 0.155672
R393 VDD2.n28 VDD2.n27 0.155672
R394 VDD2.n36 VDD2.n34 0.0529126
R395 B.n254 B.t10 1176.96
R396 B.n252 B.t14 1176.96
R397 B.n67 B.t17 1176.96
R398 B.n65 B.t21 1176.96
R399 B.n455 B.n454 585
R400 B.n456 B.n455 585
R401 B.n189 B.n64 585
R402 B.n188 B.n187 585
R403 B.n186 B.n185 585
R404 B.n184 B.n183 585
R405 B.n182 B.n181 585
R406 B.n180 B.n179 585
R407 B.n178 B.n177 585
R408 B.n176 B.n175 585
R409 B.n174 B.n173 585
R410 B.n172 B.n171 585
R411 B.n170 B.n169 585
R412 B.n168 B.n167 585
R413 B.n166 B.n165 585
R414 B.n164 B.n163 585
R415 B.n162 B.n161 585
R416 B.n160 B.n159 585
R417 B.n158 B.n157 585
R418 B.n156 B.n155 585
R419 B.n154 B.n153 585
R420 B.n152 B.n151 585
R421 B.n150 B.n149 585
R422 B.n148 B.n147 585
R423 B.n146 B.n145 585
R424 B.n144 B.n143 585
R425 B.n142 B.n141 585
R426 B.n139 B.n138 585
R427 B.n137 B.n136 585
R428 B.n135 B.n134 585
R429 B.n133 B.n132 585
R430 B.n131 B.n130 585
R431 B.n129 B.n128 585
R432 B.n127 B.n126 585
R433 B.n125 B.n124 585
R434 B.n123 B.n122 585
R435 B.n121 B.n120 585
R436 B.n119 B.n118 585
R437 B.n117 B.n116 585
R438 B.n115 B.n114 585
R439 B.n113 B.n112 585
R440 B.n111 B.n110 585
R441 B.n109 B.n108 585
R442 B.n107 B.n106 585
R443 B.n105 B.n104 585
R444 B.n103 B.n102 585
R445 B.n101 B.n100 585
R446 B.n99 B.n98 585
R447 B.n97 B.n96 585
R448 B.n95 B.n94 585
R449 B.n93 B.n92 585
R450 B.n91 B.n90 585
R451 B.n89 B.n88 585
R452 B.n87 B.n86 585
R453 B.n85 B.n84 585
R454 B.n83 B.n82 585
R455 B.n81 B.n80 585
R456 B.n79 B.n78 585
R457 B.n77 B.n76 585
R458 B.n75 B.n74 585
R459 B.n73 B.n72 585
R460 B.n71 B.n70 585
R461 B.n453 B.n33 585
R462 B.n457 B.n33 585
R463 B.n452 B.n32 585
R464 B.n458 B.n32 585
R465 B.n451 B.n450 585
R466 B.n450 B.n28 585
R467 B.n449 B.n27 585
R468 B.n464 B.n27 585
R469 B.n448 B.n26 585
R470 B.n465 B.n26 585
R471 B.n447 B.n25 585
R472 B.n466 B.n25 585
R473 B.n446 B.n445 585
R474 B.n445 B.n21 585
R475 B.n444 B.n20 585
R476 B.n472 B.n20 585
R477 B.n443 B.n19 585
R478 B.n473 B.n19 585
R479 B.n442 B.n18 585
R480 B.n474 B.n18 585
R481 B.n441 B.n440 585
R482 B.n440 B.n17 585
R483 B.n439 B.n13 585
R484 B.n480 B.n13 585
R485 B.n438 B.n12 585
R486 B.n481 B.n12 585
R487 B.n437 B.n11 585
R488 B.n482 B.n11 585
R489 B.n436 B.n435 585
R490 B.n435 B.n434 585
R491 B.n433 B.n7 585
R492 B.n488 B.n7 585
R493 B.n432 B.n6 585
R494 B.n489 B.n6 585
R495 B.n431 B.n5 585
R496 B.n490 B.n5 585
R497 B.n430 B.n429 585
R498 B.n429 B.n4 585
R499 B.n428 B.n190 585
R500 B.n428 B.n427 585
R501 B.n417 B.n191 585
R502 B.n420 B.n191 585
R503 B.n419 B.n418 585
R504 B.n421 B.n419 585
R505 B.n416 B.n196 585
R506 B.n196 B.n195 585
R507 B.n415 B.n414 585
R508 B.n414 B.n413 585
R509 B.n198 B.n197 585
R510 B.n406 B.n198 585
R511 B.n405 B.n404 585
R512 B.n407 B.n405 585
R513 B.n403 B.n202 585
R514 B.n206 B.n202 585
R515 B.n402 B.n401 585
R516 B.n401 B.n400 585
R517 B.n204 B.n203 585
R518 B.n205 B.n204 585
R519 B.n393 B.n392 585
R520 B.n394 B.n393 585
R521 B.n391 B.n210 585
R522 B.n214 B.n210 585
R523 B.n390 B.n389 585
R524 B.n389 B.n388 585
R525 B.n212 B.n211 585
R526 B.n213 B.n212 585
R527 B.n381 B.n380 585
R528 B.n382 B.n381 585
R529 B.n379 B.n219 585
R530 B.n219 B.n218 585
R531 B.n373 B.n372 585
R532 B.n371 B.n251 585
R533 B.n370 B.n250 585
R534 B.n375 B.n250 585
R535 B.n369 B.n368 585
R536 B.n367 B.n366 585
R537 B.n365 B.n364 585
R538 B.n363 B.n362 585
R539 B.n361 B.n360 585
R540 B.n359 B.n358 585
R541 B.n357 B.n356 585
R542 B.n355 B.n354 585
R543 B.n353 B.n352 585
R544 B.n351 B.n350 585
R545 B.n349 B.n348 585
R546 B.n347 B.n346 585
R547 B.n345 B.n344 585
R548 B.n343 B.n342 585
R549 B.n341 B.n340 585
R550 B.n339 B.n338 585
R551 B.n337 B.n336 585
R552 B.n335 B.n334 585
R553 B.n333 B.n332 585
R554 B.n331 B.n330 585
R555 B.n329 B.n328 585
R556 B.n327 B.n326 585
R557 B.n325 B.n324 585
R558 B.n322 B.n321 585
R559 B.n320 B.n319 585
R560 B.n318 B.n317 585
R561 B.n316 B.n315 585
R562 B.n314 B.n313 585
R563 B.n312 B.n311 585
R564 B.n310 B.n309 585
R565 B.n308 B.n307 585
R566 B.n306 B.n305 585
R567 B.n304 B.n303 585
R568 B.n302 B.n301 585
R569 B.n300 B.n299 585
R570 B.n298 B.n297 585
R571 B.n296 B.n295 585
R572 B.n294 B.n293 585
R573 B.n292 B.n291 585
R574 B.n290 B.n289 585
R575 B.n288 B.n287 585
R576 B.n286 B.n285 585
R577 B.n284 B.n283 585
R578 B.n282 B.n281 585
R579 B.n280 B.n279 585
R580 B.n278 B.n277 585
R581 B.n276 B.n275 585
R582 B.n274 B.n273 585
R583 B.n272 B.n271 585
R584 B.n270 B.n269 585
R585 B.n268 B.n267 585
R586 B.n266 B.n265 585
R587 B.n264 B.n263 585
R588 B.n262 B.n261 585
R589 B.n260 B.n259 585
R590 B.n258 B.n257 585
R591 B.n221 B.n220 585
R592 B.n378 B.n377 585
R593 B.n217 B.n216 585
R594 B.n218 B.n217 585
R595 B.n384 B.n383 585
R596 B.n383 B.n382 585
R597 B.n385 B.n215 585
R598 B.n215 B.n213 585
R599 B.n387 B.n386 585
R600 B.n388 B.n387 585
R601 B.n209 B.n208 585
R602 B.n214 B.n209 585
R603 B.n396 B.n395 585
R604 B.n395 B.n394 585
R605 B.n397 B.n207 585
R606 B.n207 B.n205 585
R607 B.n399 B.n398 585
R608 B.n400 B.n399 585
R609 B.n201 B.n200 585
R610 B.n206 B.n201 585
R611 B.n409 B.n408 585
R612 B.n408 B.n407 585
R613 B.n410 B.n199 585
R614 B.n406 B.n199 585
R615 B.n412 B.n411 585
R616 B.n413 B.n412 585
R617 B.n194 B.n193 585
R618 B.n195 B.n194 585
R619 B.n423 B.n422 585
R620 B.n422 B.n421 585
R621 B.n424 B.n192 585
R622 B.n420 B.n192 585
R623 B.n426 B.n425 585
R624 B.n427 B.n426 585
R625 B.n2 B.n0 585
R626 B.n4 B.n2 585
R627 B.n3 B.n1 585
R628 B.n489 B.n3 585
R629 B.n487 B.n486 585
R630 B.n488 B.n487 585
R631 B.n485 B.n8 585
R632 B.n434 B.n8 585
R633 B.n484 B.n483 585
R634 B.n483 B.n482 585
R635 B.n10 B.n9 585
R636 B.n481 B.n10 585
R637 B.n479 B.n478 585
R638 B.n480 B.n479 585
R639 B.n477 B.n14 585
R640 B.n17 B.n14 585
R641 B.n476 B.n475 585
R642 B.n475 B.n474 585
R643 B.n16 B.n15 585
R644 B.n473 B.n16 585
R645 B.n471 B.n470 585
R646 B.n472 B.n471 585
R647 B.n469 B.n22 585
R648 B.n22 B.n21 585
R649 B.n468 B.n467 585
R650 B.n467 B.n466 585
R651 B.n24 B.n23 585
R652 B.n465 B.n24 585
R653 B.n463 B.n462 585
R654 B.n464 B.n463 585
R655 B.n461 B.n29 585
R656 B.n29 B.n28 585
R657 B.n460 B.n459 585
R658 B.n459 B.n458 585
R659 B.n31 B.n30 585
R660 B.n457 B.n31 585
R661 B.n492 B.n491 585
R662 B.n491 B.n490 585
R663 B.n373 B.n217 473.281
R664 B.n70 B.n31 473.281
R665 B.n377 B.n219 473.281
R666 B.n455 B.n33 473.281
R667 B.n456 B.n63 256.663
R668 B.n456 B.n62 256.663
R669 B.n456 B.n61 256.663
R670 B.n456 B.n60 256.663
R671 B.n456 B.n59 256.663
R672 B.n456 B.n58 256.663
R673 B.n456 B.n57 256.663
R674 B.n456 B.n56 256.663
R675 B.n456 B.n55 256.663
R676 B.n456 B.n54 256.663
R677 B.n456 B.n53 256.663
R678 B.n456 B.n52 256.663
R679 B.n456 B.n51 256.663
R680 B.n456 B.n50 256.663
R681 B.n456 B.n49 256.663
R682 B.n456 B.n48 256.663
R683 B.n456 B.n47 256.663
R684 B.n456 B.n46 256.663
R685 B.n456 B.n45 256.663
R686 B.n456 B.n44 256.663
R687 B.n456 B.n43 256.663
R688 B.n456 B.n42 256.663
R689 B.n456 B.n41 256.663
R690 B.n456 B.n40 256.663
R691 B.n456 B.n39 256.663
R692 B.n456 B.n38 256.663
R693 B.n456 B.n37 256.663
R694 B.n456 B.n36 256.663
R695 B.n456 B.n35 256.663
R696 B.n456 B.n34 256.663
R697 B.n375 B.n374 256.663
R698 B.n375 B.n222 256.663
R699 B.n375 B.n223 256.663
R700 B.n375 B.n224 256.663
R701 B.n375 B.n225 256.663
R702 B.n375 B.n226 256.663
R703 B.n375 B.n227 256.663
R704 B.n375 B.n228 256.663
R705 B.n375 B.n229 256.663
R706 B.n375 B.n230 256.663
R707 B.n375 B.n231 256.663
R708 B.n375 B.n232 256.663
R709 B.n375 B.n233 256.663
R710 B.n375 B.n234 256.663
R711 B.n375 B.n235 256.663
R712 B.n375 B.n236 256.663
R713 B.n375 B.n237 256.663
R714 B.n375 B.n238 256.663
R715 B.n375 B.n239 256.663
R716 B.n375 B.n240 256.663
R717 B.n375 B.n241 256.663
R718 B.n375 B.n242 256.663
R719 B.n375 B.n243 256.663
R720 B.n375 B.n244 256.663
R721 B.n375 B.n245 256.663
R722 B.n375 B.n246 256.663
R723 B.n375 B.n247 256.663
R724 B.n375 B.n248 256.663
R725 B.n375 B.n249 256.663
R726 B.n376 B.n375 256.663
R727 B.n254 B.t13 198.035
R728 B.n65 B.t22 198.035
R729 B.n252 B.t16 198.035
R730 B.n67 B.t19 198.035
R731 B.n255 B.t12 188.338
R732 B.n66 B.t23 188.338
R733 B.n253 B.t15 188.338
R734 B.n68 B.t20 188.338
R735 B.n383 B.n217 163.367
R736 B.n383 B.n215 163.367
R737 B.n387 B.n215 163.367
R738 B.n387 B.n209 163.367
R739 B.n395 B.n209 163.367
R740 B.n395 B.n207 163.367
R741 B.n399 B.n207 163.367
R742 B.n399 B.n201 163.367
R743 B.n408 B.n201 163.367
R744 B.n408 B.n199 163.367
R745 B.n412 B.n199 163.367
R746 B.n412 B.n194 163.367
R747 B.n422 B.n194 163.367
R748 B.n422 B.n192 163.367
R749 B.n426 B.n192 163.367
R750 B.n426 B.n2 163.367
R751 B.n491 B.n2 163.367
R752 B.n491 B.n3 163.367
R753 B.n487 B.n3 163.367
R754 B.n487 B.n8 163.367
R755 B.n483 B.n8 163.367
R756 B.n483 B.n10 163.367
R757 B.n479 B.n10 163.367
R758 B.n479 B.n14 163.367
R759 B.n475 B.n14 163.367
R760 B.n475 B.n16 163.367
R761 B.n471 B.n16 163.367
R762 B.n471 B.n22 163.367
R763 B.n467 B.n22 163.367
R764 B.n467 B.n24 163.367
R765 B.n463 B.n24 163.367
R766 B.n463 B.n29 163.367
R767 B.n459 B.n29 163.367
R768 B.n459 B.n31 163.367
R769 B.n251 B.n250 163.367
R770 B.n368 B.n250 163.367
R771 B.n366 B.n365 163.367
R772 B.n362 B.n361 163.367
R773 B.n358 B.n357 163.367
R774 B.n354 B.n353 163.367
R775 B.n350 B.n349 163.367
R776 B.n346 B.n345 163.367
R777 B.n342 B.n341 163.367
R778 B.n338 B.n337 163.367
R779 B.n334 B.n333 163.367
R780 B.n330 B.n329 163.367
R781 B.n326 B.n325 163.367
R782 B.n321 B.n320 163.367
R783 B.n317 B.n316 163.367
R784 B.n313 B.n312 163.367
R785 B.n309 B.n308 163.367
R786 B.n305 B.n304 163.367
R787 B.n301 B.n300 163.367
R788 B.n297 B.n296 163.367
R789 B.n293 B.n292 163.367
R790 B.n289 B.n288 163.367
R791 B.n285 B.n284 163.367
R792 B.n281 B.n280 163.367
R793 B.n277 B.n276 163.367
R794 B.n273 B.n272 163.367
R795 B.n269 B.n268 163.367
R796 B.n265 B.n264 163.367
R797 B.n261 B.n260 163.367
R798 B.n257 B.n221 163.367
R799 B.n381 B.n219 163.367
R800 B.n381 B.n212 163.367
R801 B.n389 B.n212 163.367
R802 B.n389 B.n210 163.367
R803 B.n393 B.n210 163.367
R804 B.n393 B.n204 163.367
R805 B.n401 B.n204 163.367
R806 B.n401 B.n202 163.367
R807 B.n405 B.n202 163.367
R808 B.n405 B.n198 163.367
R809 B.n414 B.n198 163.367
R810 B.n414 B.n196 163.367
R811 B.n419 B.n196 163.367
R812 B.n419 B.n191 163.367
R813 B.n428 B.n191 163.367
R814 B.n429 B.n428 163.367
R815 B.n429 B.n5 163.367
R816 B.n6 B.n5 163.367
R817 B.n7 B.n6 163.367
R818 B.n435 B.n7 163.367
R819 B.n435 B.n11 163.367
R820 B.n12 B.n11 163.367
R821 B.n13 B.n12 163.367
R822 B.n440 B.n13 163.367
R823 B.n440 B.n18 163.367
R824 B.n19 B.n18 163.367
R825 B.n20 B.n19 163.367
R826 B.n445 B.n20 163.367
R827 B.n445 B.n25 163.367
R828 B.n26 B.n25 163.367
R829 B.n27 B.n26 163.367
R830 B.n450 B.n27 163.367
R831 B.n450 B.n32 163.367
R832 B.n33 B.n32 163.367
R833 B.n74 B.n73 163.367
R834 B.n78 B.n77 163.367
R835 B.n82 B.n81 163.367
R836 B.n86 B.n85 163.367
R837 B.n90 B.n89 163.367
R838 B.n94 B.n93 163.367
R839 B.n98 B.n97 163.367
R840 B.n102 B.n101 163.367
R841 B.n106 B.n105 163.367
R842 B.n110 B.n109 163.367
R843 B.n114 B.n113 163.367
R844 B.n118 B.n117 163.367
R845 B.n122 B.n121 163.367
R846 B.n126 B.n125 163.367
R847 B.n130 B.n129 163.367
R848 B.n134 B.n133 163.367
R849 B.n138 B.n137 163.367
R850 B.n143 B.n142 163.367
R851 B.n147 B.n146 163.367
R852 B.n151 B.n150 163.367
R853 B.n155 B.n154 163.367
R854 B.n159 B.n158 163.367
R855 B.n163 B.n162 163.367
R856 B.n167 B.n166 163.367
R857 B.n171 B.n170 163.367
R858 B.n175 B.n174 163.367
R859 B.n179 B.n178 163.367
R860 B.n183 B.n182 163.367
R861 B.n187 B.n186 163.367
R862 B.n455 B.n64 163.367
R863 B.n375 B.n218 110.605
R864 B.n457 B.n456 110.605
R865 B.n374 B.n373 71.676
R866 B.n368 B.n222 71.676
R867 B.n365 B.n223 71.676
R868 B.n361 B.n224 71.676
R869 B.n357 B.n225 71.676
R870 B.n353 B.n226 71.676
R871 B.n349 B.n227 71.676
R872 B.n345 B.n228 71.676
R873 B.n341 B.n229 71.676
R874 B.n337 B.n230 71.676
R875 B.n333 B.n231 71.676
R876 B.n329 B.n232 71.676
R877 B.n325 B.n233 71.676
R878 B.n320 B.n234 71.676
R879 B.n316 B.n235 71.676
R880 B.n312 B.n236 71.676
R881 B.n308 B.n237 71.676
R882 B.n304 B.n238 71.676
R883 B.n300 B.n239 71.676
R884 B.n296 B.n240 71.676
R885 B.n292 B.n241 71.676
R886 B.n288 B.n242 71.676
R887 B.n284 B.n243 71.676
R888 B.n280 B.n244 71.676
R889 B.n276 B.n245 71.676
R890 B.n272 B.n246 71.676
R891 B.n268 B.n247 71.676
R892 B.n264 B.n248 71.676
R893 B.n260 B.n249 71.676
R894 B.n376 B.n221 71.676
R895 B.n70 B.n34 71.676
R896 B.n74 B.n35 71.676
R897 B.n78 B.n36 71.676
R898 B.n82 B.n37 71.676
R899 B.n86 B.n38 71.676
R900 B.n90 B.n39 71.676
R901 B.n94 B.n40 71.676
R902 B.n98 B.n41 71.676
R903 B.n102 B.n42 71.676
R904 B.n106 B.n43 71.676
R905 B.n110 B.n44 71.676
R906 B.n114 B.n45 71.676
R907 B.n118 B.n46 71.676
R908 B.n122 B.n47 71.676
R909 B.n126 B.n48 71.676
R910 B.n130 B.n49 71.676
R911 B.n134 B.n50 71.676
R912 B.n138 B.n51 71.676
R913 B.n143 B.n52 71.676
R914 B.n147 B.n53 71.676
R915 B.n151 B.n54 71.676
R916 B.n155 B.n55 71.676
R917 B.n159 B.n56 71.676
R918 B.n163 B.n57 71.676
R919 B.n167 B.n58 71.676
R920 B.n171 B.n59 71.676
R921 B.n175 B.n60 71.676
R922 B.n179 B.n61 71.676
R923 B.n183 B.n62 71.676
R924 B.n187 B.n63 71.676
R925 B.n64 B.n63 71.676
R926 B.n186 B.n62 71.676
R927 B.n182 B.n61 71.676
R928 B.n178 B.n60 71.676
R929 B.n174 B.n59 71.676
R930 B.n170 B.n58 71.676
R931 B.n166 B.n57 71.676
R932 B.n162 B.n56 71.676
R933 B.n158 B.n55 71.676
R934 B.n154 B.n54 71.676
R935 B.n150 B.n53 71.676
R936 B.n146 B.n52 71.676
R937 B.n142 B.n51 71.676
R938 B.n137 B.n50 71.676
R939 B.n133 B.n49 71.676
R940 B.n129 B.n48 71.676
R941 B.n125 B.n47 71.676
R942 B.n121 B.n46 71.676
R943 B.n117 B.n45 71.676
R944 B.n113 B.n44 71.676
R945 B.n109 B.n43 71.676
R946 B.n105 B.n42 71.676
R947 B.n101 B.n41 71.676
R948 B.n97 B.n40 71.676
R949 B.n93 B.n39 71.676
R950 B.n89 B.n38 71.676
R951 B.n85 B.n37 71.676
R952 B.n81 B.n36 71.676
R953 B.n77 B.n35 71.676
R954 B.n73 B.n34 71.676
R955 B.n374 B.n251 71.676
R956 B.n366 B.n222 71.676
R957 B.n362 B.n223 71.676
R958 B.n358 B.n224 71.676
R959 B.n354 B.n225 71.676
R960 B.n350 B.n226 71.676
R961 B.n346 B.n227 71.676
R962 B.n342 B.n228 71.676
R963 B.n338 B.n229 71.676
R964 B.n334 B.n230 71.676
R965 B.n330 B.n231 71.676
R966 B.n326 B.n232 71.676
R967 B.n321 B.n233 71.676
R968 B.n317 B.n234 71.676
R969 B.n313 B.n235 71.676
R970 B.n309 B.n236 71.676
R971 B.n305 B.n237 71.676
R972 B.n301 B.n238 71.676
R973 B.n297 B.n239 71.676
R974 B.n293 B.n240 71.676
R975 B.n289 B.n241 71.676
R976 B.n285 B.n242 71.676
R977 B.n281 B.n243 71.676
R978 B.n277 B.n244 71.676
R979 B.n273 B.n245 71.676
R980 B.n269 B.n246 71.676
R981 B.n265 B.n247 71.676
R982 B.n261 B.n248 71.676
R983 B.n257 B.n249 71.676
R984 B.n377 B.n376 71.676
R985 B.n382 B.n218 63.2029
R986 B.n382 B.n213 63.2029
R987 B.n388 B.n213 63.2029
R988 B.n388 B.n214 63.2029
R989 B.n394 B.n205 63.2029
R990 B.n400 B.n205 63.2029
R991 B.n400 B.n206 63.2029
R992 B.n407 B.n406 63.2029
R993 B.n421 B.n195 63.2029
R994 B.n427 B.n4 63.2029
R995 B.n490 B.n4 63.2029
R996 B.n490 B.n489 63.2029
R997 B.n489 B.n488 63.2029
R998 B.n482 B.n481 63.2029
R999 B.n474 B.n17 63.2029
R1000 B.n473 B.n472 63.2029
R1001 B.n472 B.n21 63.2029
R1002 B.n466 B.n21 63.2029
R1003 B.n465 B.n464 63.2029
R1004 B.n464 B.n28 63.2029
R1005 B.n458 B.n28 63.2029
R1006 B.n458 B.n457 63.2029
R1007 B.n256 B.n255 59.5399
R1008 B.n323 B.n253 59.5399
R1009 B.n69 B.n68 59.5399
R1010 B.n140 B.n66 59.5399
R1011 B.n394 B.t11 56.6967
R1012 B.n466 B.t18 56.6967
R1013 B.t8 B.n420 51.1201
R1014 B.n434 B.t6 51.1201
R1015 B.n206 B.t1 49.2612
R1016 B.t9 B.n473 49.2612
R1017 B.n413 B.t4 47.4023
R1018 B.n480 B.t7 47.4023
R1019 B.n413 B.t2 45.5434
R1020 B.t0 B.n480 45.5434
R1021 B.n420 B.t3 41.8256
R1022 B.n434 B.t5 41.8256
R1023 B.n71 B.n30 30.7517
R1024 B.n454 B.n453 30.7517
R1025 B.n379 B.n378 30.7517
R1026 B.n372 B.n216 30.7517
R1027 B.n427 B.t3 21.3778
R1028 B.n488 B.t5 21.3778
R1029 B B.n492 18.0485
R1030 B.t2 B.n195 17.66
R1031 B.n481 B.t0 17.66
R1032 B.n406 B.t4 15.8011
R1033 B.n17 B.t7 15.8011
R1034 B.n407 B.t1 13.9422
R1035 B.n474 B.t9 13.9422
R1036 B.n421 B.t8 12.0833
R1037 B.n482 B.t6 12.0833
R1038 B.n72 B.n71 10.6151
R1039 B.n75 B.n72 10.6151
R1040 B.n76 B.n75 10.6151
R1041 B.n79 B.n76 10.6151
R1042 B.n80 B.n79 10.6151
R1043 B.n83 B.n80 10.6151
R1044 B.n84 B.n83 10.6151
R1045 B.n87 B.n84 10.6151
R1046 B.n88 B.n87 10.6151
R1047 B.n91 B.n88 10.6151
R1048 B.n92 B.n91 10.6151
R1049 B.n95 B.n92 10.6151
R1050 B.n96 B.n95 10.6151
R1051 B.n99 B.n96 10.6151
R1052 B.n100 B.n99 10.6151
R1053 B.n103 B.n100 10.6151
R1054 B.n104 B.n103 10.6151
R1055 B.n107 B.n104 10.6151
R1056 B.n108 B.n107 10.6151
R1057 B.n111 B.n108 10.6151
R1058 B.n112 B.n111 10.6151
R1059 B.n115 B.n112 10.6151
R1060 B.n116 B.n115 10.6151
R1061 B.n119 B.n116 10.6151
R1062 B.n120 B.n119 10.6151
R1063 B.n124 B.n123 10.6151
R1064 B.n127 B.n124 10.6151
R1065 B.n128 B.n127 10.6151
R1066 B.n131 B.n128 10.6151
R1067 B.n132 B.n131 10.6151
R1068 B.n135 B.n132 10.6151
R1069 B.n136 B.n135 10.6151
R1070 B.n139 B.n136 10.6151
R1071 B.n144 B.n141 10.6151
R1072 B.n145 B.n144 10.6151
R1073 B.n148 B.n145 10.6151
R1074 B.n149 B.n148 10.6151
R1075 B.n152 B.n149 10.6151
R1076 B.n153 B.n152 10.6151
R1077 B.n156 B.n153 10.6151
R1078 B.n157 B.n156 10.6151
R1079 B.n160 B.n157 10.6151
R1080 B.n161 B.n160 10.6151
R1081 B.n164 B.n161 10.6151
R1082 B.n165 B.n164 10.6151
R1083 B.n168 B.n165 10.6151
R1084 B.n169 B.n168 10.6151
R1085 B.n172 B.n169 10.6151
R1086 B.n173 B.n172 10.6151
R1087 B.n176 B.n173 10.6151
R1088 B.n177 B.n176 10.6151
R1089 B.n180 B.n177 10.6151
R1090 B.n181 B.n180 10.6151
R1091 B.n184 B.n181 10.6151
R1092 B.n185 B.n184 10.6151
R1093 B.n188 B.n185 10.6151
R1094 B.n189 B.n188 10.6151
R1095 B.n454 B.n189 10.6151
R1096 B.n380 B.n379 10.6151
R1097 B.n380 B.n211 10.6151
R1098 B.n390 B.n211 10.6151
R1099 B.n391 B.n390 10.6151
R1100 B.n392 B.n391 10.6151
R1101 B.n392 B.n203 10.6151
R1102 B.n402 B.n203 10.6151
R1103 B.n403 B.n402 10.6151
R1104 B.n404 B.n403 10.6151
R1105 B.n404 B.n197 10.6151
R1106 B.n415 B.n197 10.6151
R1107 B.n416 B.n415 10.6151
R1108 B.n418 B.n416 10.6151
R1109 B.n418 B.n417 10.6151
R1110 B.n417 B.n190 10.6151
R1111 B.n430 B.n190 10.6151
R1112 B.n431 B.n430 10.6151
R1113 B.n432 B.n431 10.6151
R1114 B.n433 B.n432 10.6151
R1115 B.n436 B.n433 10.6151
R1116 B.n437 B.n436 10.6151
R1117 B.n438 B.n437 10.6151
R1118 B.n439 B.n438 10.6151
R1119 B.n441 B.n439 10.6151
R1120 B.n442 B.n441 10.6151
R1121 B.n443 B.n442 10.6151
R1122 B.n444 B.n443 10.6151
R1123 B.n446 B.n444 10.6151
R1124 B.n447 B.n446 10.6151
R1125 B.n448 B.n447 10.6151
R1126 B.n449 B.n448 10.6151
R1127 B.n451 B.n449 10.6151
R1128 B.n452 B.n451 10.6151
R1129 B.n453 B.n452 10.6151
R1130 B.n372 B.n371 10.6151
R1131 B.n371 B.n370 10.6151
R1132 B.n370 B.n369 10.6151
R1133 B.n369 B.n367 10.6151
R1134 B.n367 B.n364 10.6151
R1135 B.n364 B.n363 10.6151
R1136 B.n363 B.n360 10.6151
R1137 B.n360 B.n359 10.6151
R1138 B.n359 B.n356 10.6151
R1139 B.n356 B.n355 10.6151
R1140 B.n355 B.n352 10.6151
R1141 B.n352 B.n351 10.6151
R1142 B.n351 B.n348 10.6151
R1143 B.n348 B.n347 10.6151
R1144 B.n347 B.n344 10.6151
R1145 B.n344 B.n343 10.6151
R1146 B.n343 B.n340 10.6151
R1147 B.n340 B.n339 10.6151
R1148 B.n339 B.n336 10.6151
R1149 B.n336 B.n335 10.6151
R1150 B.n335 B.n332 10.6151
R1151 B.n332 B.n331 10.6151
R1152 B.n331 B.n328 10.6151
R1153 B.n328 B.n327 10.6151
R1154 B.n327 B.n324 10.6151
R1155 B.n322 B.n319 10.6151
R1156 B.n319 B.n318 10.6151
R1157 B.n318 B.n315 10.6151
R1158 B.n315 B.n314 10.6151
R1159 B.n314 B.n311 10.6151
R1160 B.n311 B.n310 10.6151
R1161 B.n310 B.n307 10.6151
R1162 B.n307 B.n306 10.6151
R1163 B.n303 B.n302 10.6151
R1164 B.n302 B.n299 10.6151
R1165 B.n299 B.n298 10.6151
R1166 B.n298 B.n295 10.6151
R1167 B.n295 B.n294 10.6151
R1168 B.n294 B.n291 10.6151
R1169 B.n291 B.n290 10.6151
R1170 B.n290 B.n287 10.6151
R1171 B.n287 B.n286 10.6151
R1172 B.n286 B.n283 10.6151
R1173 B.n283 B.n282 10.6151
R1174 B.n282 B.n279 10.6151
R1175 B.n279 B.n278 10.6151
R1176 B.n278 B.n275 10.6151
R1177 B.n275 B.n274 10.6151
R1178 B.n274 B.n271 10.6151
R1179 B.n271 B.n270 10.6151
R1180 B.n270 B.n267 10.6151
R1181 B.n267 B.n266 10.6151
R1182 B.n266 B.n263 10.6151
R1183 B.n263 B.n262 10.6151
R1184 B.n262 B.n259 10.6151
R1185 B.n259 B.n258 10.6151
R1186 B.n258 B.n220 10.6151
R1187 B.n378 B.n220 10.6151
R1188 B.n384 B.n216 10.6151
R1189 B.n385 B.n384 10.6151
R1190 B.n386 B.n385 10.6151
R1191 B.n386 B.n208 10.6151
R1192 B.n396 B.n208 10.6151
R1193 B.n397 B.n396 10.6151
R1194 B.n398 B.n397 10.6151
R1195 B.n398 B.n200 10.6151
R1196 B.n409 B.n200 10.6151
R1197 B.n410 B.n409 10.6151
R1198 B.n411 B.n410 10.6151
R1199 B.n411 B.n193 10.6151
R1200 B.n423 B.n193 10.6151
R1201 B.n424 B.n423 10.6151
R1202 B.n425 B.n424 10.6151
R1203 B.n425 B.n0 10.6151
R1204 B.n486 B.n1 10.6151
R1205 B.n486 B.n485 10.6151
R1206 B.n485 B.n484 10.6151
R1207 B.n484 B.n9 10.6151
R1208 B.n478 B.n9 10.6151
R1209 B.n478 B.n477 10.6151
R1210 B.n477 B.n476 10.6151
R1211 B.n476 B.n15 10.6151
R1212 B.n470 B.n15 10.6151
R1213 B.n470 B.n469 10.6151
R1214 B.n469 B.n468 10.6151
R1215 B.n468 B.n23 10.6151
R1216 B.n462 B.n23 10.6151
R1217 B.n462 B.n461 10.6151
R1218 B.n461 B.n460 10.6151
R1219 B.n460 B.n30 10.6151
R1220 B.n255 B.n254 9.69747
R1221 B.n253 B.n252 9.69747
R1222 B.n68 B.n67 9.69747
R1223 B.n66 B.n65 9.69747
R1224 B.n123 B.n69 6.5566
R1225 B.n140 B.n139 6.5566
R1226 B.n323 B.n322 6.5566
R1227 B.n306 B.n256 6.5566
R1228 B.n214 B.t11 6.50663
R1229 B.t18 B.n465 6.50663
R1230 B.n120 B.n69 4.05904
R1231 B.n141 B.n140 4.05904
R1232 B.n324 B.n323 4.05904
R1233 B.n303 B.n256 4.05904
R1234 B.n492 B.n0 2.81026
R1235 B.n492 B.n1 2.81026
R1236 VP.n19 VP.t5 1150.79
R1237 VP.n12 VP.t9 1150.79
R1238 VP.n4 VP.t6 1150.79
R1239 VP.n10 VP.t3 1150.79
R1240 VP.n18 VP.t4 1114.27
R1241 VP.n16 VP.t2 1114.27
R1242 VP.n1 VP.t0 1114.27
R1243 VP.n3 VP.t1 1114.27
R1244 VP.n7 VP.t8 1114.27
R1245 VP.n9 VP.t7 1114.27
R1246 VP.n5 VP.n4 161.489
R1247 VP.n20 VP.n19 161.3
R1248 VP.n6 VP.n5 161.3
R1249 VP.n8 VP.n2 161.3
R1250 VP.n11 VP.n10 161.3
R1251 VP.n17 VP.n0 161.3
R1252 VP.n15 VP.n14 161.3
R1253 VP.n13 VP.n12 161.3
R1254 VP.n12 VP.n1 36.5157
R1255 VP.n15 VP.n1 36.5157
R1256 VP.n16 VP.n15 36.5157
R1257 VP.n17 VP.n16 36.5157
R1258 VP.n18 VP.n17 36.5157
R1259 VP.n19 VP.n18 36.5157
R1260 VP.n4 VP.n3 36.5157
R1261 VP.n6 VP.n3 36.5157
R1262 VP.n7 VP.n6 36.5157
R1263 VP.n8 VP.n7 36.5157
R1264 VP.n9 VP.n8 36.5157
R1265 VP.n10 VP.n9 36.5157
R1266 VP.n13 VP.n11 35.796
R1267 VP.n5 VP.n2 0.189894
R1268 VP.n11 VP.n2 0.189894
R1269 VP.n14 VP.n13 0.189894
R1270 VP.n14 VP.n0 0.189894
R1271 VP.n20 VP.n0 0.189894
R1272 VP VP.n20 0.0516364
R1273 VDD1.n32 VDD1.n31 289.615
R1274 VDD1.n67 VDD1.n66 289.615
R1275 VDD1.n31 VDD1.n30 185
R1276 VDD1.n2 VDD1.n1 185
R1277 VDD1.n25 VDD1.n24 185
R1278 VDD1.n23 VDD1.n22 185
R1279 VDD1.n6 VDD1.n5 185
R1280 VDD1.n17 VDD1.n16 185
R1281 VDD1.n15 VDD1.n14 185
R1282 VDD1.n10 VDD1.n9 185
R1283 VDD1.n45 VDD1.n44 185
R1284 VDD1.n50 VDD1.n49 185
R1285 VDD1.n52 VDD1.n51 185
R1286 VDD1.n41 VDD1.n40 185
R1287 VDD1.n58 VDD1.n57 185
R1288 VDD1.n60 VDD1.n59 185
R1289 VDD1.n37 VDD1.n36 185
R1290 VDD1.n66 VDD1.n65 185
R1291 VDD1.n11 VDD1.t3 149.525
R1292 VDD1.n46 VDD1.t0 149.525
R1293 VDD1.n31 VDD1.n1 104.615
R1294 VDD1.n24 VDD1.n1 104.615
R1295 VDD1.n24 VDD1.n23 104.615
R1296 VDD1.n23 VDD1.n5 104.615
R1297 VDD1.n16 VDD1.n5 104.615
R1298 VDD1.n16 VDD1.n15 104.615
R1299 VDD1.n15 VDD1.n9 104.615
R1300 VDD1.n50 VDD1.n44 104.615
R1301 VDD1.n51 VDD1.n50 104.615
R1302 VDD1.n51 VDD1.n40 104.615
R1303 VDD1.n58 VDD1.n40 104.615
R1304 VDD1.n59 VDD1.n58 104.615
R1305 VDD1.n59 VDD1.n36 104.615
R1306 VDD1.n66 VDD1.n36 104.615
R1307 VDD1.n71 VDD1.n70 69.5597
R1308 VDD1.n34 VDD1.n33 69.2928
R1309 VDD1.n69 VDD1.n68 69.2918
R1310 VDD1.n73 VDD1.n72 69.2917
R1311 VDD1.n34 VDD1.n32 52.7861
R1312 VDD1.n69 VDD1.n67 52.7861
R1313 VDD1.t3 VDD1.n9 52.3082
R1314 VDD1.t0 VDD1.n44 52.3082
R1315 VDD1.n73 VDD1.n71 32.2164
R1316 VDD1.n30 VDD1.n0 12.8005
R1317 VDD1.n65 VDD1.n35 12.8005
R1318 VDD1.n29 VDD1.n2 12.0247
R1319 VDD1.n64 VDD1.n37 12.0247
R1320 VDD1.n26 VDD1.n25 11.249
R1321 VDD1.n61 VDD1.n60 11.249
R1322 VDD1.n22 VDD1.n4 10.4732
R1323 VDD1.n57 VDD1.n39 10.4732
R1324 VDD1.n11 VDD1.n10 10.2746
R1325 VDD1.n46 VDD1.n45 10.2746
R1326 VDD1.n21 VDD1.n6 9.69747
R1327 VDD1.n56 VDD1.n41 9.69747
R1328 VDD1.n28 VDD1.n0 9.45567
R1329 VDD1.n63 VDD1.n35 9.45567
R1330 VDD1.n8 VDD1.n7 9.3005
R1331 VDD1.n19 VDD1.n18 9.3005
R1332 VDD1.n21 VDD1.n20 9.3005
R1333 VDD1.n4 VDD1.n3 9.3005
R1334 VDD1.n27 VDD1.n26 9.3005
R1335 VDD1.n29 VDD1.n28 9.3005
R1336 VDD1.n13 VDD1.n12 9.3005
R1337 VDD1.n48 VDD1.n47 9.3005
R1338 VDD1.n43 VDD1.n42 9.3005
R1339 VDD1.n54 VDD1.n53 9.3005
R1340 VDD1.n56 VDD1.n55 9.3005
R1341 VDD1.n39 VDD1.n38 9.3005
R1342 VDD1.n62 VDD1.n61 9.3005
R1343 VDD1.n64 VDD1.n63 9.3005
R1344 VDD1.n18 VDD1.n17 8.92171
R1345 VDD1.n53 VDD1.n52 8.92171
R1346 VDD1.n14 VDD1.n8 8.14595
R1347 VDD1.n49 VDD1.n43 8.14595
R1348 VDD1.n13 VDD1.n10 7.3702
R1349 VDD1.n48 VDD1.n45 7.3702
R1350 VDD1.n14 VDD1.n13 5.81868
R1351 VDD1.n49 VDD1.n48 5.81868
R1352 VDD1.n17 VDD1.n8 5.04292
R1353 VDD1.n52 VDD1.n43 5.04292
R1354 VDD1.n18 VDD1.n6 4.26717
R1355 VDD1.n53 VDD1.n41 4.26717
R1356 VDD1.n22 VDD1.n21 3.49141
R1357 VDD1.n57 VDD1.n56 3.49141
R1358 VDD1.n72 VDD1.t2 3.01879
R1359 VDD1.n72 VDD1.t6 3.01879
R1360 VDD1.n33 VDD1.t8 3.01879
R1361 VDD1.n33 VDD1.t1 3.01879
R1362 VDD1.n70 VDD1.t5 3.01879
R1363 VDD1.n70 VDD1.t4 3.01879
R1364 VDD1.n68 VDD1.t9 3.01879
R1365 VDD1.n68 VDD1.t7 3.01879
R1366 VDD1.n12 VDD1.n11 2.84308
R1367 VDD1.n47 VDD1.n46 2.84308
R1368 VDD1.n25 VDD1.n4 2.71565
R1369 VDD1.n60 VDD1.n39 2.71565
R1370 VDD1.n26 VDD1.n2 1.93989
R1371 VDD1.n61 VDD1.n37 1.93989
R1372 VDD1.n30 VDD1.n29 1.16414
R1373 VDD1.n65 VDD1.n64 1.16414
R1374 VDD1.n32 VDD1.n0 0.388379
R1375 VDD1.n67 VDD1.n35 0.388379
R1376 VDD1 VDD1.n73 0.265586
R1377 VDD1 VDD1.n34 0.166448
R1378 VDD1.n28 VDD1.n27 0.155672
R1379 VDD1.n27 VDD1.n3 0.155672
R1380 VDD1.n20 VDD1.n3 0.155672
R1381 VDD1.n20 VDD1.n19 0.155672
R1382 VDD1.n19 VDD1.n7 0.155672
R1383 VDD1.n12 VDD1.n7 0.155672
R1384 VDD1.n47 VDD1.n42 0.155672
R1385 VDD1.n54 VDD1.n42 0.155672
R1386 VDD1.n55 VDD1.n54 0.155672
R1387 VDD1.n55 VDD1.n38 0.155672
R1388 VDD1.n62 VDD1.n38 0.155672
R1389 VDD1.n63 VDD1.n62 0.155672
R1390 VDD1.n71 VDD1.n69 0.0529126
C0 VDD1 VN 0.147658f
C1 VDD1 VTAIL 15.318401f
C2 VDD2 VN 1.68255f
C3 VDD1 VP 1.805f
C4 VDD2 VTAIL 15.3506f
C5 VDD2 VP 0.273106f
C6 VN VTAIL 1.47515f
C7 VP VN 3.80889f
C8 VDD2 VDD1 0.643228f
C9 VP VTAIL 1.48965f
C10 VDD2 B 3.383593f
C11 VDD1 B 3.226351f
C12 VTAIL B 3.927841f
C13 VN B 5.63111f
C14 VP B 4.527647f
C15 VDD1.n0 B 0.017354f
C16 VDD1.n1 B 0.039095f
C17 VDD1.n2 B 0.017513f
C18 VDD1.n3 B 0.03078f
C19 VDD1.n4 B 0.01654f
C20 VDD1.n5 B 0.039095f
C21 VDD1.n6 B 0.017513f
C22 VDD1.n7 B 0.03078f
C23 VDD1.n8 B 0.01654f
C24 VDD1.n9 B 0.029321f
C25 VDD1.n10 B 0.027637f
C26 VDD1.t3 B 0.065216f
C27 VDD1.n11 B 0.157796f
C28 VDD1.n12 B 0.807798f
C29 VDD1.n13 B 0.01654f
C30 VDD1.n14 B 0.017513f
C31 VDD1.n15 B 0.039095f
C32 VDD1.n16 B 0.039095f
C33 VDD1.n17 B 0.017513f
C34 VDD1.n18 B 0.01654f
C35 VDD1.n19 B 0.03078f
C36 VDD1.n20 B 0.03078f
C37 VDD1.n21 B 0.01654f
C38 VDD1.n22 B 0.017513f
C39 VDD1.n23 B 0.039095f
C40 VDD1.n24 B 0.039095f
C41 VDD1.n25 B 0.017513f
C42 VDD1.n26 B 0.01654f
C43 VDD1.n27 B 0.03078f
C44 VDD1.n28 B 0.079557f
C45 VDD1.n29 B 0.01654f
C46 VDD1.n30 B 0.017513f
C47 VDD1.n31 B 0.080226f
C48 VDD1.n32 B 0.089674f
C49 VDD1.t8 B 0.159563f
C50 VDD1.t1 B 0.159563f
C51 VDD1.n33 B 1.35777f
C52 VDD1.n34 B 0.403516f
C53 VDD1.n35 B 0.017354f
C54 VDD1.n36 B 0.039095f
C55 VDD1.n37 B 0.017513f
C56 VDD1.n38 B 0.03078f
C57 VDD1.n39 B 0.01654f
C58 VDD1.n40 B 0.039095f
C59 VDD1.n41 B 0.017513f
C60 VDD1.n42 B 0.03078f
C61 VDD1.n43 B 0.01654f
C62 VDD1.n44 B 0.029321f
C63 VDD1.n45 B 0.027637f
C64 VDD1.t0 B 0.065216f
C65 VDD1.n46 B 0.157796f
C66 VDD1.n47 B 0.807798f
C67 VDD1.n48 B 0.01654f
C68 VDD1.n49 B 0.017513f
C69 VDD1.n50 B 0.039095f
C70 VDD1.n51 B 0.039095f
C71 VDD1.n52 B 0.017513f
C72 VDD1.n53 B 0.01654f
C73 VDD1.n54 B 0.03078f
C74 VDD1.n55 B 0.03078f
C75 VDD1.n56 B 0.01654f
C76 VDD1.n57 B 0.017513f
C77 VDD1.n58 B 0.039095f
C78 VDD1.n59 B 0.039095f
C79 VDD1.n60 B 0.017513f
C80 VDD1.n61 B 0.01654f
C81 VDD1.n62 B 0.03078f
C82 VDD1.n63 B 0.079557f
C83 VDD1.n64 B 0.01654f
C84 VDD1.n65 B 0.017513f
C85 VDD1.n66 B 0.080226f
C86 VDD1.n67 B 0.089674f
C87 VDD1.t9 B 0.159563f
C88 VDD1.t7 B 0.159563f
C89 VDD1.n68 B 1.35777f
C90 VDD1.n69 B 0.405868f
C91 VDD1.t5 B 0.159563f
C92 VDD1.t4 B 0.159563f
C93 VDD1.n70 B 1.35902f
C94 VDD1.n71 B 1.65438f
C95 VDD1.t2 B 0.159563f
C96 VDD1.t6 B 0.159563f
C97 VDD1.n72 B 1.35777f
C98 VDD1.n73 B 2.12182f
C99 VP.n0 B 0.031886f
C100 VP.t4 B 0.101173f
C101 VP.t2 B 0.101173f
C102 VP.t0 B 0.101173f
C103 VP.n1 B 0.049631f
C104 VP.n2 B 0.031886f
C105 VP.t7 B 0.101173f
C106 VP.t8 B 0.101173f
C107 VP.t1 B 0.101173f
C108 VP.n3 B 0.049631f
C109 VP.t6 B 0.102698f
C110 VP.n4 B 0.057152f
C111 VP.n5 B 0.067073f
C112 VP.n6 B 0.010578f
C113 VP.n7 B 0.049631f
C114 VP.n8 B 0.010578f
C115 VP.n9 B 0.049631f
C116 VP.t3 B 0.102698f
C117 VP.n10 B 0.057111f
C118 VP.n11 B 0.991759f
C119 VP.t9 B 0.102698f
C120 VP.n12 B 0.057111f
C121 VP.n13 B 1.02387f
C122 VP.n14 B 0.031886f
C123 VP.n15 B 0.010578f
C124 VP.n16 B 0.049631f
C125 VP.n17 B 0.010578f
C126 VP.n18 B 0.049631f
C127 VP.t5 B 0.102698f
C128 VP.n19 B 0.057111f
C129 VP.n20 B 0.024711f
C130 VDD2.n0 B 0.017598f
C131 VDD2.n1 B 0.039645f
C132 VDD2.n2 B 0.017759f
C133 VDD2.n3 B 0.031213f
C134 VDD2.n4 B 0.016773f
C135 VDD2.n5 B 0.039645f
C136 VDD2.n6 B 0.017759f
C137 VDD2.n7 B 0.031213f
C138 VDD2.n8 B 0.016773f
C139 VDD2.n9 B 0.029734f
C140 VDD2.n10 B 0.028025f
C141 VDD2.t1 B 0.066133f
C142 VDD2.n11 B 0.160016f
C143 VDD2.n12 B 0.819165f
C144 VDD2.n13 B 0.016773f
C145 VDD2.n14 B 0.017759f
C146 VDD2.n15 B 0.039645f
C147 VDD2.n16 B 0.039645f
C148 VDD2.n17 B 0.017759f
C149 VDD2.n18 B 0.016773f
C150 VDD2.n19 B 0.031213f
C151 VDD2.n20 B 0.031213f
C152 VDD2.n21 B 0.016773f
C153 VDD2.n22 B 0.017759f
C154 VDD2.n23 B 0.039645f
C155 VDD2.n24 B 0.039645f
C156 VDD2.n25 B 0.017759f
C157 VDD2.n26 B 0.016773f
C158 VDD2.n27 B 0.031213f
C159 VDD2.n28 B 0.080677f
C160 VDD2.n29 B 0.016773f
C161 VDD2.n30 B 0.017759f
C162 VDD2.n31 B 0.081355f
C163 VDD2.n32 B 0.090936f
C164 VDD2.t3 B 0.161808f
C165 VDD2.t4 B 0.161808f
C166 VDD2.n33 B 1.37688f
C167 VDD2.n34 B 0.411579f
C168 VDD2.t5 B 0.161808f
C169 VDD2.t7 B 0.161808f
C170 VDD2.n35 B 1.37814f
C171 VDD2.n36 B 1.59792f
C172 VDD2.n37 B 0.017598f
C173 VDD2.n38 B 0.039645f
C174 VDD2.n39 B 0.017759f
C175 VDD2.n40 B 0.031213f
C176 VDD2.n41 B 0.016773f
C177 VDD2.n42 B 0.039645f
C178 VDD2.n43 B 0.017759f
C179 VDD2.n44 B 0.031213f
C180 VDD2.n45 B 0.016773f
C181 VDD2.n46 B 0.029734f
C182 VDD2.n47 B 0.028025f
C183 VDD2.t6 B 0.066133f
C184 VDD2.n48 B 0.160016f
C185 VDD2.n49 B 0.819165f
C186 VDD2.n50 B 0.016773f
C187 VDD2.n51 B 0.017759f
C188 VDD2.n52 B 0.039645f
C189 VDD2.n53 B 0.039645f
C190 VDD2.n54 B 0.017759f
C191 VDD2.n55 B 0.016773f
C192 VDD2.n56 B 0.031213f
C193 VDD2.n57 B 0.031213f
C194 VDD2.n58 B 0.016773f
C195 VDD2.n59 B 0.017759f
C196 VDD2.n60 B 0.039645f
C197 VDD2.n61 B 0.039645f
C198 VDD2.n62 B 0.017759f
C199 VDD2.n63 B 0.016773f
C200 VDD2.n64 B 0.031213f
C201 VDD2.n65 B 0.080677f
C202 VDD2.n66 B 0.016773f
C203 VDD2.n67 B 0.017759f
C204 VDD2.n68 B 0.081355f
C205 VDD2.n69 B 0.090055f
C206 VDD2.n70 B 1.89921f
C207 VDD2.t0 B 0.161808f
C208 VDD2.t9 B 0.161808f
C209 VDD2.n71 B 1.37687f
C210 VDD2.n72 B 0.302222f
C211 VDD2.t8 B 0.161808f
C212 VDD2.t2 B 0.161808f
C213 VDD2.n73 B 1.37811f
C214 VTAIL.t12 B 0.174456f
C215 VTAIL.t11 B 0.174456f
C216 VTAIL.n0 B 1.40376f
C217 VTAIL.n1 B 0.411793f
C218 VTAIL.n2 B 0.018974f
C219 VTAIL.n3 B 0.042744f
C220 VTAIL.n4 B 0.019148f
C221 VTAIL.n5 B 0.033653f
C222 VTAIL.n6 B 0.018084f
C223 VTAIL.n7 B 0.042744f
C224 VTAIL.n8 B 0.019148f
C225 VTAIL.n9 B 0.033653f
C226 VTAIL.n10 B 0.018084f
C227 VTAIL.n11 B 0.032058f
C228 VTAIL.n12 B 0.030216f
C229 VTAIL.t3 B 0.071303f
C230 VTAIL.n13 B 0.172524f
C231 VTAIL.n14 B 0.883197f
C232 VTAIL.n15 B 0.018084f
C233 VTAIL.n16 B 0.019148f
C234 VTAIL.n17 B 0.042744f
C235 VTAIL.n18 B 0.042744f
C236 VTAIL.n19 B 0.019148f
C237 VTAIL.n20 B 0.018084f
C238 VTAIL.n21 B 0.033653f
C239 VTAIL.n22 B 0.033653f
C240 VTAIL.n23 B 0.018084f
C241 VTAIL.n24 B 0.019148f
C242 VTAIL.n25 B 0.042744f
C243 VTAIL.n26 B 0.042744f
C244 VTAIL.n27 B 0.019148f
C245 VTAIL.n28 B 0.018084f
C246 VTAIL.n29 B 0.033653f
C247 VTAIL.n30 B 0.086983f
C248 VTAIL.n31 B 0.018084f
C249 VTAIL.n32 B 0.019148f
C250 VTAIL.n33 B 0.087715f
C251 VTAIL.n34 B 0.073915f
C252 VTAIL.n35 B 0.154483f
C253 VTAIL.t2 B 0.174456f
C254 VTAIL.t8 B 0.174456f
C255 VTAIL.n36 B 1.40376f
C256 VTAIL.n37 B 0.389591f
C257 VTAIL.t1 B 0.174456f
C258 VTAIL.t4 B 0.174456f
C259 VTAIL.n38 B 1.40376f
C260 VTAIL.n39 B 1.50671f
C261 VTAIL.t17 B 0.174456f
C262 VTAIL.t10 B 0.174456f
C263 VTAIL.n40 B 1.40376f
C264 VTAIL.n41 B 1.50672f
C265 VTAIL.t16 B 0.174456f
C266 VTAIL.t18 B 0.174456f
C267 VTAIL.n42 B 1.40376f
C268 VTAIL.n43 B 0.389592f
C269 VTAIL.n44 B 0.018974f
C270 VTAIL.n45 B 0.042744f
C271 VTAIL.n46 B 0.019148f
C272 VTAIL.n47 B 0.033653f
C273 VTAIL.n48 B 0.018084f
C274 VTAIL.n49 B 0.042744f
C275 VTAIL.n50 B 0.019148f
C276 VTAIL.n51 B 0.033653f
C277 VTAIL.n52 B 0.018084f
C278 VTAIL.n53 B 0.032058f
C279 VTAIL.n54 B 0.030216f
C280 VTAIL.t15 B 0.071303f
C281 VTAIL.n55 B 0.172524f
C282 VTAIL.n56 B 0.883197f
C283 VTAIL.n57 B 0.018084f
C284 VTAIL.n58 B 0.019148f
C285 VTAIL.n59 B 0.042744f
C286 VTAIL.n60 B 0.042744f
C287 VTAIL.n61 B 0.019148f
C288 VTAIL.n62 B 0.018084f
C289 VTAIL.n63 B 0.033653f
C290 VTAIL.n64 B 0.033653f
C291 VTAIL.n65 B 0.018084f
C292 VTAIL.n66 B 0.019148f
C293 VTAIL.n67 B 0.042744f
C294 VTAIL.n68 B 0.042744f
C295 VTAIL.n69 B 0.019148f
C296 VTAIL.n70 B 0.018084f
C297 VTAIL.n71 B 0.033653f
C298 VTAIL.n72 B 0.086983f
C299 VTAIL.n73 B 0.018084f
C300 VTAIL.n74 B 0.019148f
C301 VTAIL.n75 B 0.087715f
C302 VTAIL.n76 B 0.073915f
C303 VTAIL.n77 B 0.154483f
C304 VTAIL.t5 B 0.174456f
C305 VTAIL.t6 B 0.174456f
C306 VTAIL.n78 B 1.40376f
C307 VTAIL.n79 B 0.417169f
C308 VTAIL.t0 B 0.174456f
C309 VTAIL.t7 B 0.174456f
C310 VTAIL.n80 B 1.40376f
C311 VTAIL.n81 B 0.389592f
C312 VTAIL.n82 B 0.018974f
C313 VTAIL.n83 B 0.042744f
C314 VTAIL.n84 B 0.019148f
C315 VTAIL.n85 B 0.033653f
C316 VTAIL.n86 B 0.018084f
C317 VTAIL.n87 B 0.042744f
C318 VTAIL.n88 B 0.019148f
C319 VTAIL.n89 B 0.033653f
C320 VTAIL.n90 B 0.018084f
C321 VTAIL.n91 B 0.032058f
C322 VTAIL.n92 B 0.030216f
C323 VTAIL.t9 B 0.071303f
C324 VTAIL.n93 B 0.172524f
C325 VTAIL.n94 B 0.883197f
C326 VTAIL.n95 B 0.018084f
C327 VTAIL.n96 B 0.019148f
C328 VTAIL.n97 B 0.042744f
C329 VTAIL.n98 B 0.042744f
C330 VTAIL.n99 B 0.019148f
C331 VTAIL.n100 B 0.018084f
C332 VTAIL.n101 B 0.033653f
C333 VTAIL.n102 B 0.033653f
C334 VTAIL.n103 B 0.018084f
C335 VTAIL.n104 B 0.019148f
C336 VTAIL.n105 B 0.042744f
C337 VTAIL.n106 B 0.042744f
C338 VTAIL.n107 B 0.019148f
C339 VTAIL.n108 B 0.018084f
C340 VTAIL.n109 B 0.033653f
C341 VTAIL.n110 B 0.086983f
C342 VTAIL.n111 B 0.018084f
C343 VTAIL.n112 B 0.019148f
C344 VTAIL.n113 B 0.087715f
C345 VTAIL.n114 B 0.073915f
C346 VTAIL.n115 B 1.19729f
C347 VTAIL.n116 B 0.018974f
C348 VTAIL.n117 B 0.042744f
C349 VTAIL.n118 B 0.019148f
C350 VTAIL.n119 B 0.033653f
C351 VTAIL.n120 B 0.018084f
C352 VTAIL.n121 B 0.042744f
C353 VTAIL.n122 B 0.019148f
C354 VTAIL.n123 B 0.033653f
C355 VTAIL.n124 B 0.018084f
C356 VTAIL.n125 B 0.032058f
C357 VTAIL.n126 B 0.030216f
C358 VTAIL.t13 B 0.071303f
C359 VTAIL.n127 B 0.172524f
C360 VTAIL.n128 B 0.883197f
C361 VTAIL.n129 B 0.018084f
C362 VTAIL.n130 B 0.019148f
C363 VTAIL.n131 B 0.042744f
C364 VTAIL.n132 B 0.042744f
C365 VTAIL.n133 B 0.019148f
C366 VTAIL.n134 B 0.018084f
C367 VTAIL.n135 B 0.033653f
C368 VTAIL.n136 B 0.033653f
C369 VTAIL.n137 B 0.018084f
C370 VTAIL.n138 B 0.019148f
C371 VTAIL.n139 B 0.042744f
C372 VTAIL.n140 B 0.042744f
C373 VTAIL.n141 B 0.019148f
C374 VTAIL.n142 B 0.018084f
C375 VTAIL.n143 B 0.033653f
C376 VTAIL.n144 B 0.086983f
C377 VTAIL.n145 B 0.018084f
C378 VTAIL.n146 B 0.019148f
C379 VTAIL.n147 B 0.087715f
C380 VTAIL.n148 B 0.073915f
C381 VTAIL.n149 B 1.19729f
C382 VTAIL.t14 B 0.174456f
C383 VTAIL.t19 B 0.174456f
C384 VTAIL.n150 B 1.40376f
C385 VTAIL.n151 B 0.348225f
C386 VN.n0 B 0.031514f
C387 VN.t4 B 0.099994f
C388 VN.t5 B 0.099994f
C389 VN.t6 B 0.099994f
C390 VN.n1 B 0.049052f
C391 VN.t8 B 0.101501f
C392 VN.n2 B 0.056486f
C393 VN.n3 B 0.066291f
C394 VN.n4 B 0.010454f
C395 VN.n5 B 0.049052f
C396 VN.n6 B 0.010454f
C397 VN.n7 B 0.049052f
C398 VN.t2 B 0.101501f
C399 VN.n8 B 0.056445f
C400 VN.n9 B 0.024423f
C401 VN.n10 B 0.031514f
C402 VN.t3 B 0.101501f
C403 VN.t9 B 0.099994f
C404 VN.t0 B 0.099994f
C405 VN.t1 B 0.099994f
C406 VN.n11 B 0.049052f
C407 VN.t7 B 0.101501f
C408 VN.n12 B 0.056486f
C409 VN.n13 B 0.066291f
C410 VN.n14 B 0.010454f
C411 VN.n15 B 0.049052f
C412 VN.n16 B 0.010454f
C413 VN.n17 B 0.049052f
C414 VN.n18 B 0.056445f
C415 VN.n19 B 1.00111f
.ends

