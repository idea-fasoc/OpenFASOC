* NGSPICE file created from diff_pair_sample_1247.ext - technology: sky130A

.subckt diff_pair_sample_1247 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X1 VTAIL.t12 VN.t0 VDD2.t7 B.t20 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=1.73415 ps=10.84 w=10.51 l=0.18
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=0 ps=0 w=10.51 l=0.18
X3 VTAIL.t11 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=1.73415 ps=10.84 w=10.51 l=0.18
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=0 ps=0 w=10.51 l=0.18
X5 VDD1.t5 VP.t2 VTAIL.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=4.0989 ps=21.8 w=10.51 l=0.18
X6 VDD2.t6 VN.t1 VTAIL.t13 B.t18 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X7 VTAIL.t14 VN.t2 VDD2.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X8 VDD2.t4 VN.t3 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=4.0989 ps=21.8 w=10.51 l=0.18
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=0 ps=0 w=10.51 l=0.18
X10 VTAIL.t1 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X11 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X12 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=0 ps=0 w=10.51 l=0.18
X13 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=1.73415 ps=10.84 w=10.51 l=0.18
X14 VTAIL.t9 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X15 VTAIL.t6 VP.t4 VDD1.t3 B.t20 sky130_fd_pr__nfet_01v8 ad=4.0989 pd=21.8 as=1.73415 ps=10.84 w=10.51 l=0.18
X16 VTAIL.t10 VP.t5 VDD1.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X17 VDD1.t1 VP.t6 VTAIL.t4 B.t18 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=1.73415 ps=10.84 w=10.51 l=0.18
X18 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=4.0989 ps=21.8 w=10.51 l=0.18
X19 VDD1.t0 VP.t7 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.73415 pd=10.84 as=4.0989 ps=21.8 w=10.51 l=0.18
R0 VP.n13 VP.t2 1621.27
R1 VP.n9 VP.t1 1621.27
R2 VP.n2 VP.t4 1621.27
R3 VP.n6 VP.t7 1621.27
R4 VP.n12 VP.t3 1582.57
R5 VP.n10 VP.t0 1582.57
R6 VP.n3 VP.t6 1582.57
R7 VP.n5 VP.t5 1582.57
R8 VP.n2 VP.n1 161.489
R9 VP.n14 VP.n13 161.3
R10 VP.n4 VP.n1 161.3
R11 VP.n7 VP.n6 161.3
R12 VP.n11 VP.n0 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n8 VP.n7 38.4702
R15 VP.n11 VP.n10 37.246
R16 VP.n12 VP.n11 37.246
R17 VP.n4 VP.n3 37.246
R18 VP.n5 VP.n4 37.246
R19 VP.n10 VP.n9 35.7853
R20 VP.n13 VP.n12 35.7853
R21 VP.n3 VP.n2 35.7853
R22 VP.n6 VP.n5 35.7853
R23 VP.n7 VP.n1 0.189894
R24 VP.n8 VP.n0 0.189894
R25 VP.n14 VP.n0 0.189894
R26 VP VP.n14 0.0516364
R27 VTAIL.n11 VTAIL.t6 51.373
R28 VTAIL.n10 VTAIL.t15 51.373
R29 VTAIL.n7 VTAIL.t2 51.373
R30 VTAIL.n14 VTAIL.t7 51.3727
R31 VTAIL.n15 VTAIL.t3 51.3727
R32 VTAIL.n2 VTAIL.t12 51.3727
R33 VTAIL.n3 VTAIL.t8 51.3727
R34 VTAIL.n6 VTAIL.t11 51.3727
R35 VTAIL.n13 VTAIL.n12 49.4891
R36 VTAIL.n9 VTAIL.n8 49.4891
R37 VTAIL.n1 VTAIL.n0 49.4888
R38 VTAIL.n5 VTAIL.n4 49.4888
R39 VTAIL.n15 VTAIL.n14 21.8669
R40 VTAIL.n7 VTAIL.n6 21.8669
R41 VTAIL.n0 VTAIL.t13 1.88442
R42 VTAIL.n0 VTAIL.t14 1.88442
R43 VTAIL.n4 VTAIL.t5 1.88442
R44 VTAIL.n4 VTAIL.t9 1.88442
R45 VTAIL.n12 VTAIL.t4 1.88442
R46 VTAIL.n12 VTAIL.t10 1.88442
R47 VTAIL.n8 VTAIL.t0 1.88442
R48 VTAIL.n8 VTAIL.t1 1.88442
R49 VTAIL.n11 VTAIL.n10 0.470328
R50 VTAIL.n3 VTAIL.n2 0.470328
R51 VTAIL.n9 VTAIL.n7 0.440155
R52 VTAIL.n10 VTAIL.n9 0.440155
R53 VTAIL.n13 VTAIL.n11 0.440155
R54 VTAIL.n14 VTAIL.n13 0.440155
R55 VTAIL.n6 VTAIL.n5 0.440155
R56 VTAIL.n5 VTAIL.n3 0.440155
R57 VTAIL.n2 VTAIL.n1 0.440155
R58 VTAIL VTAIL.n15 0.381966
R59 VTAIL VTAIL.n1 0.0586897
R60 VDD1 VDD1.n0 66.4459
R61 VDD1.n3 VDD1.n2 66.3321
R62 VDD1.n3 VDD1.n1 66.3321
R63 VDD1.n5 VDD1.n4 66.1677
R64 VDD1.n5 VDD1.n3 35.3371
R65 VDD1.n4 VDD1.t2 1.88442
R66 VDD1.n4 VDD1.t0 1.88442
R67 VDD1.n0 VDD1.t3 1.88442
R68 VDD1.n0 VDD1.t1 1.88442
R69 VDD1.n2 VDD1.t4 1.88442
R70 VDD1.n2 VDD1.t5 1.88442
R71 VDD1.n1 VDD1.t6 1.88442
R72 VDD1.n1 VDD1.t7 1.88442
R73 VDD1 VDD1.n5 0.162138
R74 B.n78 B.t4 1650.22
R75 B.n76 B.t12 1650.22
R76 B.n321 B.t8 1650.22
R77 B.n318 B.t15 1650.22
R78 B.n556 B.n555 585
R79 B.n246 B.n75 585
R80 B.n245 B.n244 585
R81 B.n243 B.n242 585
R82 B.n241 B.n240 585
R83 B.n239 B.n238 585
R84 B.n237 B.n236 585
R85 B.n235 B.n234 585
R86 B.n233 B.n232 585
R87 B.n231 B.n230 585
R88 B.n229 B.n228 585
R89 B.n227 B.n226 585
R90 B.n225 B.n224 585
R91 B.n223 B.n222 585
R92 B.n221 B.n220 585
R93 B.n219 B.n218 585
R94 B.n217 B.n216 585
R95 B.n215 B.n214 585
R96 B.n213 B.n212 585
R97 B.n211 B.n210 585
R98 B.n209 B.n208 585
R99 B.n207 B.n206 585
R100 B.n205 B.n204 585
R101 B.n203 B.n202 585
R102 B.n201 B.n200 585
R103 B.n199 B.n198 585
R104 B.n197 B.n196 585
R105 B.n195 B.n194 585
R106 B.n193 B.n192 585
R107 B.n191 B.n190 585
R108 B.n189 B.n188 585
R109 B.n187 B.n186 585
R110 B.n185 B.n184 585
R111 B.n183 B.n182 585
R112 B.n181 B.n180 585
R113 B.n179 B.n178 585
R114 B.n177 B.n176 585
R115 B.n174 B.n173 585
R116 B.n172 B.n171 585
R117 B.n170 B.n169 585
R118 B.n168 B.n167 585
R119 B.n166 B.n165 585
R120 B.n164 B.n163 585
R121 B.n162 B.n161 585
R122 B.n160 B.n159 585
R123 B.n158 B.n157 585
R124 B.n156 B.n155 585
R125 B.n153 B.n152 585
R126 B.n151 B.n150 585
R127 B.n149 B.n148 585
R128 B.n147 B.n146 585
R129 B.n145 B.n144 585
R130 B.n143 B.n142 585
R131 B.n141 B.n140 585
R132 B.n139 B.n138 585
R133 B.n137 B.n136 585
R134 B.n135 B.n134 585
R135 B.n133 B.n132 585
R136 B.n131 B.n130 585
R137 B.n129 B.n128 585
R138 B.n127 B.n126 585
R139 B.n125 B.n124 585
R140 B.n123 B.n122 585
R141 B.n121 B.n120 585
R142 B.n119 B.n118 585
R143 B.n117 B.n116 585
R144 B.n115 B.n114 585
R145 B.n113 B.n112 585
R146 B.n111 B.n110 585
R147 B.n109 B.n108 585
R148 B.n107 B.n106 585
R149 B.n105 B.n104 585
R150 B.n103 B.n102 585
R151 B.n101 B.n100 585
R152 B.n99 B.n98 585
R153 B.n97 B.n96 585
R154 B.n95 B.n94 585
R155 B.n93 B.n92 585
R156 B.n91 B.n90 585
R157 B.n89 B.n88 585
R158 B.n87 B.n86 585
R159 B.n85 B.n84 585
R160 B.n83 B.n82 585
R161 B.n81 B.n80 585
R162 B.n554 B.n33 585
R163 B.n559 B.n33 585
R164 B.n553 B.n32 585
R165 B.n560 B.n32 585
R166 B.n552 B.n551 585
R167 B.n551 B.n28 585
R168 B.n550 B.n27 585
R169 B.n566 B.n27 585
R170 B.n549 B.n26 585
R171 B.n567 B.n26 585
R172 B.n548 B.n25 585
R173 B.n568 B.n25 585
R174 B.n547 B.n546 585
R175 B.n546 B.n21 585
R176 B.n545 B.n20 585
R177 B.n574 B.n20 585
R178 B.n544 B.n19 585
R179 B.n575 B.n19 585
R180 B.n543 B.n18 585
R181 B.n576 B.n18 585
R182 B.n542 B.n541 585
R183 B.n541 B.n17 585
R184 B.n540 B.n12 585
R185 B.n582 B.n12 585
R186 B.n539 B.n11 585
R187 B.n583 B.n11 585
R188 B.n538 B.n10 585
R189 B.n584 B.n10 585
R190 B.n537 B.n7 585
R191 B.n587 B.n7 585
R192 B.n536 B.n6 585
R193 B.n588 B.n6 585
R194 B.n535 B.n5 585
R195 B.n589 B.n5 585
R196 B.n534 B.n533 585
R197 B.n533 B.n4 585
R198 B.n532 B.n247 585
R199 B.n532 B.n531 585
R200 B.n522 B.n248 585
R201 B.n249 B.n248 585
R202 B.n524 B.n523 585
R203 B.n525 B.n524 585
R204 B.n521 B.n253 585
R205 B.n256 B.n253 585
R206 B.n520 B.n519 585
R207 B.n519 B.n518 585
R208 B.n255 B.n254 585
R209 B.n511 B.n255 585
R210 B.n510 B.n509 585
R211 B.n512 B.n510 585
R212 B.n508 B.n261 585
R213 B.n261 B.n260 585
R214 B.n507 B.n506 585
R215 B.n506 B.n505 585
R216 B.n263 B.n262 585
R217 B.n264 B.n263 585
R218 B.n498 B.n497 585
R219 B.n499 B.n498 585
R220 B.n496 B.n269 585
R221 B.n269 B.n268 585
R222 B.n495 B.n494 585
R223 B.n494 B.n493 585
R224 B.n271 B.n270 585
R225 B.n272 B.n271 585
R226 B.n489 B.n488 585
R227 B.n275 B.n274 585
R228 B.n485 B.n484 585
R229 B.n486 B.n485 585
R230 B.n483 B.n317 585
R231 B.n482 B.n481 585
R232 B.n480 B.n479 585
R233 B.n478 B.n477 585
R234 B.n476 B.n475 585
R235 B.n474 B.n473 585
R236 B.n472 B.n471 585
R237 B.n470 B.n469 585
R238 B.n468 B.n467 585
R239 B.n466 B.n465 585
R240 B.n464 B.n463 585
R241 B.n462 B.n461 585
R242 B.n460 B.n459 585
R243 B.n458 B.n457 585
R244 B.n456 B.n455 585
R245 B.n454 B.n453 585
R246 B.n452 B.n451 585
R247 B.n450 B.n449 585
R248 B.n448 B.n447 585
R249 B.n446 B.n445 585
R250 B.n444 B.n443 585
R251 B.n442 B.n441 585
R252 B.n440 B.n439 585
R253 B.n438 B.n437 585
R254 B.n436 B.n435 585
R255 B.n434 B.n433 585
R256 B.n432 B.n431 585
R257 B.n430 B.n429 585
R258 B.n428 B.n427 585
R259 B.n426 B.n425 585
R260 B.n424 B.n423 585
R261 B.n422 B.n421 585
R262 B.n420 B.n419 585
R263 B.n418 B.n417 585
R264 B.n416 B.n415 585
R265 B.n414 B.n413 585
R266 B.n412 B.n411 585
R267 B.n410 B.n409 585
R268 B.n408 B.n407 585
R269 B.n406 B.n405 585
R270 B.n404 B.n403 585
R271 B.n402 B.n401 585
R272 B.n400 B.n399 585
R273 B.n398 B.n397 585
R274 B.n396 B.n395 585
R275 B.n394 B.n393 585
R276 B.n392 B.n391 585
R277 B.n390 B.n389 585
R278 B.n388 B.n387 585
R279 B.n386 B.n385 585
R280 B.n384 B.n383 585
R281 B.n382 B.n381 585
R282 B.n380 B.n379 585
R283 B.n378 B.n377 585
R284 B.n376 B.n375 585
R285 B.n374 B.n373 585
R286 B.n372 B.n371 585
R287 B.n370 B.n369 585
R288 B.n368 B.n367 585
R289 B.n366 B.n365 585
R290 B.n364 B.n363 585
R291 B.n362 B.n361 585
R292 B.n360 B.n359 585
R293 B.n358 B.n357 585
R294 B.n356 B.n355 585
R295 B.n354 B.n353 585
R296 B.n352 B.n351 585
R297 B.n350 B.n349 585
R298 B.n348 B.n347 585
R299 B.n346 B.n345 585
R300 B.n344 B.n343 585
R301 B.n342 B.n341 585
R302 B.n340 B.n339 585
R303 B.n338 B.n337 585
R304 B.n336 B.n335 585
R305 B.n334 B.n333 585
R306 B.n332 B.n331 585
R307 B.n330 B.n329 585
R308 B.n328 B.n327 585
R309 B.n326 B.n325 585
R310 B.n324 B.n316 585
R311 B.n486 B.n316 585
R312 B.n490 B.n273 585
R313 B.n273 B.n272 585
R314 B.n492 B.n491 585
R315 B.n493 B.n492 585
R316 B.n267 B.n266 585
R317 B.n268 B.n267 585
R318 B.n501 B.n500 585
R319 B.n500 B.n499 585
R320 B.n502 B.n265 585
R321 B.n265 B.n264 585
R322 B.n504 B.n503 585
R323 B.n505 B.n504 585
R324 B.n259 B.n258 585
R325 B.n260 B.n259 585
R326 B.n514 B.n513 585
R327 B.n513 B.n512 585
R328 B.n515 B.n257 585
R329 B.n511 B.n257 585
R330 B.n517 B.n516 585
R331 B.n518 B.n517 585
R332 B.n252 B.n251 585
R333 B.n256 B.n252 585
R334 B.n527 B.n526 585
R335 B.n526 B.n525 585
R336 B.n528 B.n250 585
R337 B.n250 B.n249 585
R338 B.n530 B.n529 585
R339 B.n531 B.n530 585
R340 B.n3 B.n0 585
R341 B.n4 B.n3 585
R342 B.n586 B.n1 585
R343 B.n587 B.n586 585
R344 B.n585 B.n9 585
R345 B.n585 B.n584 585
R346 B.n14 B.n8 585
R347 B.n583 B.n8 585
R348 B.n581 B.n580 585
R349 B.n582 B.n581 585
R350 B.n579 B.n13 585
R351 B.n17 B.n13 585
R352 B.n578 B.n577 585
R353 B.n577 B.n576 585
R354 B.n16 B.n15 585
R355 B.n575 B.n16 585
R356 B.n573 B.n572 585
R357 B.n574 B.n573 585
R358 B.n571 B.n22 585
R359 B.n22 B.n21 585
R360 B.n570 B.n569 585
R361 B.n569 B.n568 585
R362 B.n24 B.n23 585
R363 B.n567 B.n24 585
R364 B.n565 B.n564 585
R365 B.n566 B.n565 585
R366 B.n563 B.n29 585
R367 B.n29 B.n28 585
R368 B.n562 B.n561 585
R369 B.n561 B.n560 585
R370 B.n31 B.n30 585
R371 B.n559 B.n31 585
R372 B.n590 B.n589 585
R373 B.n588 B.n2 585
R374 B.n80 B.n31 521.33
R375 B.n556 B.n33 521.33
R376 B.n316 B.n271 521.33
R377 B.n488 B.n273 521.33
R378 B.n558 B.n557 256.663
R379 B.n558 B.n74 256.663
R380 B.n558 B.n73 256.663
R381 B.n558 B.n72 256.663
R382 B.n558 B.n71 256.663
R383 B.n558 B.n70 256.663
R384 B.n558 B.n69 256.663
R385 B.n558 B.n68 256.663
R386 B.n558 B.n67 256.663
R387 B.n558 B.n66 256.663
R388 B.n558 B.n65 256.663
R389 B.n558 B.n64 256.663
R390 B.n558 B.n63 256.663
R391 B.n558 B.n62 256.663
R392 B.n558 B.n61 256.663
R393 B.n558 B.n60 256.663
R394 B.n558 B.n59 256.663
R395 B.n558 B.n58 256.663
R396 B.n558 B.n57 256.663
R397 B.n558 B.n56 256.663
R398 B.n558 B.n55 256.663
R399 B.n558 B.n54 256.663
R400 B.n558 B.n53 256.663
R401 B.n558 B.n52 256.663
R402 B.n558 B.n51 256.663
R403 B.n558 B.n50 256.663
R404 B.n558 B.n49 256.663
R405 B.n558 B.n48 256.663
R406 B.n558 B.n47 256.663
R407 B.n558 B.n46 256.663
R408 B.n558 B.n45 256.663
R409 B.n558 B.n44 256.663
R410 B.n558 B.n43 256.663
R411 B.n558 B.n42 256.663
R412 B.n558 B.n41 256.663
R413 B.n558 B.n40 256.663
R414 B.n558 B.n39 256.663
R415 B.n558 B.n38 256.663
R416 B.n558 B.n37 256.663
R417 B.n558 B.n36 256.663
R418 B.n558 B.n35 256.663
R419 B.n558 B.n34 256.663
R420 B.n487 B.n486 256.663
R421 B.n486 B.n276 256.663
R422 B.n486 B.n277 256.663
R423 B.n486 B.n278 256.663
R424 B.n486 B.n279 256.663
R425 B.n486 B.n280 256.663
R426 B.n486 B.n281 256.663
R427 B.n486 B.n282 256.663
R428 B.n486 B.n283 256.663
R429 B.n486 B.n284 256.663
R430 B.n486 B.n285 256.663
R431 B.n486 B.n286 256.663
R432 B.n486 B.n287 256.663
R433 B.n486 B.n288 256.663
R434 B.n486 B.n289 256.663
R435 B.n486 B.n290 256.663
R436 B.n486 B.n291 256.663
R437 B.n486 B.n292 256.663
R438 B.n486 B.n293 256.663
R439 B.n486 B.n294 256.663
R440 B.n486 B.n295 256.663
R441 B.n486 B.n296 256.663
R442 B.n486 B.n297 256.663
R443 B.n486 B.n298 256.663
R444 B.n486 B.n299 256.663
R445 B.n486 B.n300 256.663
R446 B.n486 B.n301 256.663
R447 B.n486 B.n302 256.663
R448 B.n486 B.n303 256.663
R449 B.n486 B.n304 256.663
R450 B.n486 B.n305 256.663
R451 B.n486 B.n306 256.663
R452 B.n486 B.n307 256.663
R453 B.n486 B.n308 256.663
R454 B.n486 B.n309 256.663
R455 B.n486 B.n310 256.663
R456 B.n486 B.n311 256.663
R457 B.n486 B.n312 256.663
R458 B.n486 B.n313 256.663
R459 B.n486 B.n314 256.663
R460 B.n486 B.n315 256.663
R461 B.n592 B.n591 256.663
R462 B.n84 B.n83 163.367
R463 B.n88 B.n87 163.367
R464 B.n92 B.n91 163.367
R465 B.n96 B.n95 163.367
R466 B.n100 B.n99 163.367
R467 B.n104 B.n103 163.367
R468 B.n108 B.n107 163.367
R469 B.n112 B.n111 163.367
R470 B.n116 B.n115 163.367
R471 B.n120 B.n119 163.367
R472 B.n124 B.n123 163.367
R473 B.n128 B.n127 163.367
R474 B.n132 B.n131 163.367
R475 B.n136 B.n135 163.367
R476 B.n140 B.n139 163.367
R477 B.n144 B.n143 163.367
R478 B.n148 B.n147 163.367
R479 B.n152 B.n151 163.367
R480 B.n157 B.n156 163.367
R481 B.n161 B.n160 163.367
R482 B.n165 B.n164 163.367
R483 B.n169 B.n168 163.367
R484 B.n173 B.n172 163.367
R485 B.n178 B.n177 163.367
R486 B.n182 B.n181 163.367
R487 B.n186 B.n185 163.367
R488 B.n190 B.n189 163.367
R489 B.n194 B.n193 163.367
R490 B.n198 B.n197 163.367
R491 B.n202 B.n201 163.367
R492 B.n206 B.n205 163.367
R493 B.n210 B.n209 163.367
R494 B.n214 B.n213 163.367
R495 B.n218 B.n217 163.367
R496 B.n222 B.n221 163.367
R497 B.n226 B.n225 163.367
R498 B.n230 B.n229 163.367
R499 B.n234 B.n233 163.367
R500 B.n238 B.n237 163.367
R501 B.n242 B.n241 163.367
R502 B.n244 B.n75 163.367
R503 B.n494 B.n271 163.367
R504 B.n494 B.n269 163.367
R505 B.n498 B.n269 163.367
R506 B.n498 B.n263 163.367
R507 B.n506 B.n263 163.367
R508 B.n506 B.n261 163.367
R509 B.n510 B.n261 163.367
R510 B.n510 B.n255 163.367
R511 B.n519 B.n255 163.367
R512 B.n519 B.n253 163.367
R513 B.n524 B.n253 163.367
R514 B.n524 B.n248 163.367
R515 B.n532 B.n248 163.367
R516 B.n533 B.n532 163.367
R517 B.n533 B.n5 163.367
R518 B.n6 B.n5 163.367
R519 B.n7 B.n6 163.367
R520 B.n10 B.n7 163.367
R521 B.n11 B.n10 163.367
R522 B.n12 B.n11 163.367
R523 B.n541 B.n12 163.367
R524 B.n541 B.n18 163.367
R525 B.n19 B.n18 163.367
R526 B.n20 B.n19 163.367
R527 B.n546 B.n20 163.367
R528 B.n546 B.n25 163.367
R529 B.n26 B.n25 163.367
R530 B.n27 B.n26 163.367
R531 B.n551 B.n27 163.367
R532 B.n551 B.n32 163.367
R533 B.n33 B.n32 163.367
R534 B.n485 B.n275 163.367
R535 B.n485 B.n317 163.367
R536 B.n481 B.n480 163.367
R537 B.n477 B.n476 163.367
R538 B.n473 B.n472 163.367
R539 B.n469 B.n468 163.367
R540 B.n465 B.n464 163.367
R541 B.n461 B.n460 163.367
R542 B.n457 B.n456 163.367
R543 B.n453 B.n452 163.367
R544 B.n449 B.n448 163.367
R545 B.n445 B.n444 163.367
R546 B.n441 B.n440 163.367
R547 B.n437 B.n436 163.367
R548 B.n433 B.n432 163.367
R549 B.n429 B.n428 163.367
R550 B.n425 B.n424 163.367
R551 B.n421 B.n420 163.367
R552 B.n417 B.n416 163.367
R553 B.n413 B.n412 163.367
R554 B.n409 B.n408 163.367
R555 B.n405 B.n404 163.367
R556 B.n401 B.n400 163.367
R557 B.n397 B.n396 163.367
R558 B.n393 B.n392 163.367
R559 B.n389 B.n388 163.367
R560 B.n385 B.n384 163.367
R561 B.n381 B.n380 163.367
R562 B.n377 B.n376 163.367
R563 B.n373 B.n372 163.367
R564 B.n369 B.n368 163.367
R565 B.n365 B.n364 163.367
R566 B.n361 B.n360 163.367
R567 B.n357 B.n356 163.367
R568 B.n353 B.n352 163.367
R569 B.n349 B.n348 163.367
R570 B.n345 B.n344 163.367
R571 B.n341 B.n340 163.367
R572 B.n337 B.n336 163.367
R573 B.n333 B.n332 163.367
R574 B.n329 B.n328 163.367
R575 B.n325 B.n316 163.367
R576 B.n492 B.n273 163.367
R577 B.n492 B.n267 163.367
R578 B.n500 B.n267 163.367
R579 B.n500 B.n265 163.367
R580 B.n504 B.n265 163.367
R581 B.n504 B.n259 163.367
R582 B.n513 B.n259 163.367
R583 B.n513 B.n257 163.367
R584 B.n517 B.n257 163.367
R585 B.n517 B.n252 163.367
R586 B.n526 B.n252 163.367
R587 B.n526 B.n250 163.367
R588 B.n530 B.n250 163.367
R589 B.n530 B.n3 163.367
R590 B.n590 B.n3 163.367
R591 B.n586 B.n2 163.367
R592 B.n586 B.n585 163.367
R593 B.n585 B.n8 163.367
R594 B.n581 B.n8 163.367
R595 B.n581 B.n13 163.367
R596 B.n577 B.n13 163.367
R597 B.n577 B.n16 163.367
R598 B.n573 B.n16 163.367
R599 B.n573 B.n22 163.367
R600 B.n569 B.n22 163.367
R601 B.n569 B.n24 163.367
R602 B.n565 B.n24 163.367
R603 B.n565 B.n29 163.367
R604 B.n561 B.n29 163.367
R605 B.n561 B.n31 163.367
R606 B.n486 B.n272 91.2897
R607 B.n559 B.n558 91.2897
R608 B.n76 B.t13 83.9244
R609 B.n321 B.t11 83.9244
R610 B.n78 B.t6 83.9116
R611 B.n318 B.t17 83.9116
R612 B.n77 B.t14 74.0335
R613 B.n322 B.t10 74.0335
R614 B.n79 B.t7 74.0207
R615 B.n319 B.t16 74.0207
R616 B.n80 B.n34 71.676
R617 B.n84 B.n35 71.676
R618 B.n88 B.n36 71.676
R619 B.n92 B.n37 71.676
R620 B.n96 B.n38 71.676
R621 B.n100 B.n39 71.676
R622 B.n104 B.n40 71.676
R623 B.n108 B.n41 71.676
R624 B.n112 B.n42 71.676
R625 B.n116 B.n43 71.676
R626 B.n120 B.n44 71.676
R627 B.n124 B.n45 71.676
R628 B.n128 B.n46 71.676
R629 B.n132 B.n47 71.676
R630 B.n136 B.n48 71.676
R631 B.n140 B.n49 71.676
R632 B.n144 B.n50 71.676
R633 B.n148 B.n51 71.676
R634 B.n152 B.n52 71.676
R635 B.n157 B.n53 71.676
R636 B.n161 B.n54 71.676
R637 B.n165 B.n55 71.676
R638 B.n169 B.n56 71.676
R639 B.n173 B.n57 71.676
R640 B.n178 B.n58 71.676
R641 B.n182 B.n59 71.676
R642 B.n186 B.n60 71.676
R643 B.n190 B.n61 71.676
R644 B.n194 B.n62 71.676
R645 B.n198 B.n63 71.676
R646 B.n202 B.n64 71.676
R647 B.n206 B.n65 71.676
R648 B.n210 B.n66 71.676
R649 B.n214 B.n67 71.676
R650 B.n218 B.n68 71.676
R651 B.n222 B.n69 71.676
R652 B.n226 B.n70 71.676
R653 B.n230 B.n71 71.676
R654 B.n234 B.n72 71.676
R655 B.n238 B.n73 71.676
R656 B.n242 B.n74 71.676
R657 B.n557 B.n75 71.676
R658 B.n557 B.n556 71.676
R659 B.n244 B.n74 71.676
R660 B.n241 B.n73 71.676
R661 B.n237 B.n72 71.676
R662 B.n233 B.n71 71.676
R663 B.n229 B.n70 71.676
R664 B.n225 B.n69 71.676
R665 B.n221 B.n68 71.676
R666 B.n217 B.n67 71.676
R667 B.n213 B.n66 71.676
R668 B.n209 B.n65 71.676
R669 B.n205 B.n64 71.676
R670 B.n201 B.n63 71.676
R671 B.n197 B.n62 71.676
R672 B.n193 B.n61 71.676
R673 B.n189 B.n60 71.676
R674 B.n185 B.n59 71.676
R675 B.n181 B.n58 71.676
R676 B.n177 B.n57 71.676
R677 B.n172 B.n56 71.676
R678 B.n168 B.n55 71.676
R679 B.n164 B.n54 71.676
R680 B.n160 B.n53 71.676
R681 B.n156 B.n52 71.676
R682 B.n151 B.n51 71.676
R683 B.n147 B.n50 71.676
R684 B.n143 B.n49 71.676
R685 B.n139 B.n48 71.676
R686 B.n135 B.n47 71.676
R687 B.n131 B.n46 71.676
R688 B.n127 B.n45 71.676
R689 B.n123 B.n44 71.676
R690 B.n119 B.n43 71.676
R691 B.n115 B.n42 71.676
R692 B.n111 B.n41 71.676
R693 B.n107 B.n40 71.676
R694 B.n103 B.n39 71.676
R695 B.n99 B.n38 71.676
R696 B.n95 B.n37 71.676
R697 B.n91 B.n36 71.676
R698 B.n87 B.n35 71.676
R699 B.n83 B.n34 71.676
R700 B.n488 B.n487 71.676
R701 B.n317 B.n276 71.676
R702 B.n480 B.n277 71.676
R703 B.n476 B.n278 71.676
R704 B.n472 B.n279 71.676
R705 B.n468 B.n280 71.676
R706 B.n464 B.n281 71.676
R707 B.n460 B.n282 71.676
R708 B.n456 B.n283 71.676
R709 B.n452 B.n284 71.676
R710 B.n448 B.n285 71.676
R711 B.n444 B.n286 71.676
R712 B.n440 B.n287 71.676
R713 B.n436 B.n288 71.676
R714 B.n432 B.n289 71.676
R715 B.n428 B.n290 71.676
R716 B.n424 B.n291 71.676
R717 B.n420 B.n292 71.676
R718 B.n416 B.n293 71.676
R719 B.n412 B.n294 71.676
R720 B.n408 B.n295 71.676
R721 B.n404 B.n296 71.676
R722 B.n400 B.n297 71.676
R723 B.n396 B.n298 71.676
R724 B.n392 B.n299 71.676
R725 B.n388 B.n300 71.676
R726 B.n384 B.n301 71.676
R727 B.n380 B.n302 71.676
R728 B.n376 B.n303 71.676
R729 B.n372 B.n304 71.676
R730 B.n368 B.n305 71.676
R731 B.n364 B.n306 71.676
R732 B.n360 B.n307 71.676
R733 B.n356 B.n308 71.676
R734 B.n352 B.n309 71.676
R735 B.n348 B.n310 71.676
R736 B.n344 B.n311 71.676
R737 B.n340 B.n312 71.676
R738 B.n336 B.n313 71.676
R739 B.n332 B.n314 71.676
R740 B.n328 B.n315 71.676
R741 B.n487 B.n275 71.676
R742 B.n481 B.n276 71.676
R743 B.n477 B.n277 71.676
R744 B.n473 B.n278 71.676
R745 B.n469 B.n279 71.676
R746 B.n465 B.n280 71.676
R747 B.n461 B.n281 71.676
R748 B.n457 B.n282 71.676
R749 B.n453 B.n283 71.676
R750 B.n449 B.n284 71.676
R751 B.n445 B.n285 71.676
R752 B.n441 B.n286 71.676
R753 B.n437 B.n287 71.676
R754 B.n433 B.n288 71.676
R755 B.n429 B.n289 71.676
R756 B.n425 B.n290 71.676
R757 B.n421 B.n291 71.676
R758 B.n417 B.n292 71.676
R759 B.n413 B.n293 71.676
R760 B.n409 B.n294 71.676
R761 B.n405 B.n295 71.676
R762 B.n401 B.n296 71.676
R763 B.n397 B.n297 71.676
R764 B.n393 B.n298 71.676
R765 B.n389 B.n299 71.676
R766 B.n385 B.n300 71.676
R767 B.n381 B.n301 71.676
R768 B.n377 B.n302 71.676
R769 B.n373 B.n303 71.676
R770 B.n369 B.n304 71.676
R771 B.n365 B.n305 71.676
R772 B.n361 B.n306 71.676
R773 B.n357 B.n307 71.676
R774 B.n353 B.n308 71.676
R775 B.n349 B.n309 71.676
R776 B.n345 B.n310 71.676
R777 B.n341 B.n311 71.676
R778 B.n337 B.n312 71.676
R779 B.n333 B.n313 71.676
R780 B.n329 B.n314 71.676
R781 B.n325 B.n315 71.676
R782 B.n591 B.n590 71.676
R783 B.n591 B.n2 71.676
R784 B.n154 B.n79 59.5399
R785 B.n175 B.n77 59.5399
R786 B.n323 B.n322 59.5399
R787 B.n320 B.n319 59.5399
R788 B.n493 B.n272 47.3873
R789 B.n493 B.n268 47.3873
R790 B.n499 B.n268 47.3873
R791 B.n505 B.n264 47.3873
R792 B.n505 B.n260 47.3873
R793 B.n512 B.n260 47.3873
R794 B.n512 B.n511 47.3873
R795 B.n518 B.n256 47.3873
R796 B.n531 B.n249 47.3873
R797 B.n589 B.n4 47.3873
R798 B.n589 B.n588 47.3873
R799 B.n588 B.n587 47.3873
R800 B.n584 B.n583 47.3873
R801 B.n576 B.n17 47.3873
R802 B.n575 B.n574 47.3873
R803 B.n574 B.n21 47.3873
R804 B.n568 B.n21 47.3873
R805 B.n568 B.n567 47.3873
R806 B.n566 B.n28 47.3873
R807 B.n560 B.n28 47.3873
R808 B.n560 B.n559 47.3873
R809 B.n499 B.t9 44.5998
R810 B.t5 B.n566 44.5998
R811 B.n525 B.t0 40.4186
R812 B.t21 B.n4 40.4186
R813 B.n587 B.t20 40.4186
R814 B.n582 B.t19 40.4186
R815 B.n490 B.n489 33.8737
R816 B.n324 B.n270 33.8737
R817 B.n555 B.n554 33.8737
R818 B.n81 B.n30 33.8737
R819 B.n511 B.t2 30.6625
R820 B.n525 B.t1 30.6625
R821 B.t18 B.n582 30.6625
R822 B.t3 B.n575 30.6625
R823 B B.n592 18.0485
R824 B.n518 B.t2 16.7252
R825 B.t1 B.n249 16.7252
R826 B.n583 B.t18 16.7252
R827 B.n576 B.t3 16.7252
R828 B.n491 B.n490 10.6151
R829 B.n491 B.n266 10.6151
R830 B.n501 B.n266 10.6151
R831 B.n502 B.n501 10.6151
R832 B.n503 B.n502 10.6151
R833 B.n503 B.n258 10.6151
R834 B.n514 B.n258 10.6151
R835 B.n515 B.n514 10.6151
R836 B.n516 B.n515 10.6151
R837 B.n516 B.n251 10.6151
R838 B.n527 B.n251 10.6151
R839 B.n528 B.n527 10.6151
R840 B.n529 B.n528 10.6151
R841 B.n529 B.n0 10.6151
R842 B.n489 B.n274 10.6151
R843 B.n484 B.n274 10.6151
R844 B.n484 B.n483 10.6151
R845 B.n483 B.n482 10.6151
R846 B.n482 B.n479 10.6151
R847 B.n479 B.n478 10.6151
R848 B.n478 B.n475 10.6151
R849 B.n475 B.n474 10.6151
R850 B.n474 B.n471 10.6151
R851 B.n471 B.n470 10.6151
R852 B.n470 B.n467 10.6151
R853 B.n467 B.n466 10.6151
R854 B.n466 B.n463 10.6151
R855 B.n463 B.n462 10.6151
R856 B.n462 B.n459 10.6151
R857 B.n459 B.n458 10.6151
R858 B.n458 B.n455 10.6151
R859 B.n455 B.n454 10.6151
R860 B.n454 B.n451 10.6151
R861 B.n451 B.n450 10.6151
R862 B.n450 B.n447 10.6151
R863 B.n447 B.n446 10.6151
R864 B.n446 B.n443 10.6151
R865 B.n443 B.n442 10.6151
R866 B.n442 B.n439 10.6151
R867 B.n439 B.n438 10.6151
R868 B.n438 B.n435 10.6151
R869 B.n435 B.n434 10.6151
R870 B.n434 B.n431 10.6151
R871 B.n431 B.n430 10.6151
R872 B.n430 B.n427 10.6151
R873 B.n427 B.n426 10.6151
R874 B.n426 B.n423 10.6151
R875 B.n423 B.n422 10.6151
R876 B.n422 B.n419 10.6151
R877 B.n419 B.n418 10.6151
R878 B.n415 B.n414 10.6151
R879 B.n414 B.n411 10.6151
R880 B.n411 B.n410 10.6151
R881 B.n410 B.n407 10.6151
R882 B.n407 B.n406 10.6151
R883 B.n406 B.n403 10.6151
R884 B.n403 B.n402 10.6151
R885 B.n402 B.n399 10.6151
R886 B.n399 B.n398 10.6151
R887 B.n395 B.n394 10.6151
R888 B.n394 B.n391 10.6151
R889 B.n391 B.n390 10.6151
R890 B.n390 B.n387 10.6151
R891 B.n387 B.n386 10.6151
R892 B.n386 B.n383 10.6151
R893 B.n383 B.n382 10.6151
R894 B.n382 B.n379 10.6151
R895 B.n379 B.n378 10.6151
R896 B.n378 B.n375 10.6151
R897 B.n375 B.n374 10.6151
R898 B.n374 B.n371 10.6151
R899 B.n371 B.n370 10.6151
R900 B.n370 B.n367 10.6151
R901 B.n367 B.n366 10.6151
R902 B.n366 B.n363 10.6151
R903 B.n363 B.n362 10.6151
R904 B.n362 B.n359 10.6151
R905 B.n359 B.n358 10.6151
R906 B.n358 B.n355 10.6151
R907 B.n355 B.n354 10.6151
R908 B.n354 B.n351 10.6151
R909 B.n351 B.n350 10.6151
R910 B.n350 B.n347 10.6151
R911 B.n347 B.n346 10.6151
R912 B.n346 B.n343 10.6151
R913 B.n343 B.n342 10.6151
R914 B.n342 B.n339 10.6151
R915 B.n339 B.n338 10.6151
R916 B.n338 B.n335 10.6151
R917 B.n335 B.n334 10.6151
R918 B.n334 B.n331 10.6151
R919 B.n331 B.n330 10.6151
R920 B.n330 B.n327 10.6151
R921 B.n327 B.n326 10.6151
R922 B.n326 B.n324 10.6151
R923 B.n495 B.n270 10.6151
R924 B.n496 B.n495 10.6151
R925 B.n497 B.n496 10.6151
R926 B.n497 B.n262 10.6151
R927 B.n507 B.n262 10.6151
R928 B.n508 B.n507 10.6151
R929 B.n509 B.n508 10.6151
R930 B.n509 B.n254 10.6151
R931 B.n520 B.n254 10.6151
R932 B.n521 B.n520 10.6151
R933 B.n523 B.n521 10.6151
R934 B.n523 B.n522 10.6151
R935 B.n522 B.n247 10.6151
R936 B.n534 B.n247 10.6151
R937 B.n535 B.n534 10.6151
R938 B.n536 B.n535 10.6151
R939 B.n537 B.n536 10.6151
R940 B.n538 B.n537 10.6151
R941 B.n539 B.n538 10.6151
R942 B.n540 B.n539 10.6151
R943 B.n542 B.n540 10.6151
R944 B.n543 B.n542 10.6151
R945 B.n544 B.n543 10.6151
R946 B.n545 B.n544 10.6151
R947 B.n547 B.n545 10.6151
R948 B.n548 B.n547 10.6151
R949 B.n549 B.n548 10.6151
R950 B.n550 B.n549 10.6151
R951 B.n552 B.n550 10.6151
R952 B.n553 B.n552 10.6151
R953 B.n554 B.n553 10.6151
R954 B.n9 B.n1 10.6151
R955 B.n14 B.n9 10.6151
R956 B.n580 B.n14 10.6151
R957 B.n580 B.n579 10.6151
R958 B.n579 B.n578 10.6151
R959 B.n578 B.n15 10.6151
R960 B.n572 B.n15 10.6151
R961 B.n572 B.n571 10.6151
R962 B.n571 B.n570 10.6151
R963 B.n570 B.n23 10.6151
R964 B.n564 B.n23 10.6151
R965 B.n564 B.n563 10.6151
R966 B.n563 B.n562 10.6151
R967 B.n562 B.n30 10.6151
R968 B.n82 B.n81 10.6151
R969 B.n85 B.n82 10.6151
R970 B.n86 B.n85 10.6151
R971 B.n89 B.n86 10.6151
R972 B.n90 B.n89 10.6151
R973 B.n93 B.n90 10.6151
R974 B.n94 B.n93 10.6151
R975 B.n97 B.n94 10.6151
R976 B.n98 B.n97 10.6151
R977 B.n101 B.n98 10.6151
R978 B.n102 B.n101 10.6151
R979 B.n105 B.n102 10.6151
R980 B.n106 B.n105 10.6151
R981 B.n109 B.n106 10.6151
R982 B.n110 B.n109 10.6151
R983 B.n113 B.n110 10.6151
R984 B.n114 B.n113 10.6151
R985 B.n117 B.n114 10.6151
R986 B.n118 B.n117 10.6151
R987 B.n121 B.n118 10.6151
R988 B.n122 B.n121 10.6151
R989 B.n125 B.n122 10.6151
R990 B.n126 B.n125 10.6151
R991 B.n129 B.n126 10.6151
R992 B.n130 B.n129 10.6151
R993 B.n133 B.n130 10.6151
R994 B.n134 B.n133 10.6151
R995 B.n137 B.n134 10.6151
R996 B.n138 B.n137 10.6151
R997 B.n141 B.n138 10.6151
R998 B.n142 B.n141 10.6151
R999 B.n145 B.n142 10.6151
R1000 B.n146 B.n145 10.6151
R1001 B.n149 B.n146 10.6151
R1002 B.n150 B.n149 10.6151
R1003 B.n153 B.n150 10.6151
R1004 B.n158 B.n155 10.6151
R1005 B.n159 B.n158 10.6151
R1006 B.n162 B.n159 10.6151
R1007 B.n163 B.n162 10.6151
R1008 B.n166 B.n163 10.6151
R1009 B.n167 B.n166 10.6151
R1010 B.n170 B.n167 10.6151
R1011 B.n171 B.n170 10.6151
R1012 B.n174 B.n171 10.6151
R1013 B.n179 B.n176 10.6151
R1014 B.n180 B.n179 10.6151
R1015 B.n183 B.n180 10.6151
R1016 B.n184 B.n183 10.6151
R1017 B.n187 B.n184 10.6151
R1018 B.n188 B.n187 10.6151
R1019 B.n191 B.n188 10.6151
R1020 B.n192 B.n191 10.6151
R1021 B.n195 B.n192 10.6151
R1022 B.n196 B.n195 10.6151
R1023 B.n199 B.n196 10.6151
R1024 B.n200 B.n199 10.6151
R1025 B.n203 B.n200 10.6151
R1026 B.n204 B.n203 10.6151
R1027 B.n207 B.n204 10.6151
R1028 B.n208 B.n207 10.6151
R1029 B.n211 B.n208 10.6151
R1030 B.n212 B.n211 10.6151
R1031 B.n215 B.n212 10.6151
R1032 B.n216 B.n215 10.6151
R1033 B.n219 B.n216 10.6151
R1034 B.n220 B.n219 10.6151
R1035 B.n223 B.n220 10.6151
R1036 B.n224 B.n223 10.6151
R1037 B.n227 B.n224 10.6151
R1038 B.n228 B.n227 10.6151
R1039 B.n231 B.n228 10.6151
R1040 B.n232 B.n231 10.6151
R1041 B.n235 B.n232 10.6151
R1042 B.n236 B.n235 10.6151
R1043 B.n239 B.n236 10.6151
R1044 B.n240 B.n239 10.6151
R1045 B.n243 B.n240 10.6151
R1046 B.n245 B.n243 10.6151
R1047 B.n246 B.n245 10.6151
R1048 B.n555 B.n246 10.6151
R1049 B.n79 B.n78 9.89141
R1050 B.n77 B.n76 9.89141
R1051 B.n322 B.n321 9.89141
R1052 B.n319 B.n318 9.89141
R1053 B.n418 B.n320 9.36635
R1054 B.n395 B.n323 9.36635
R1055 B.n154 B.n153 9.36635
R1056 B.n176 B.n175 9.36635
R1057 B.n592 B.n0 8.11757
R1058 B.n592 B.n1 8.11757
R1059 B.n256 B.t0 6.96914
R1060 B.n531 B.t21 6.96914
R1061 B.n584 B.t20 6.96914
R1062 B.n17 B.t19 6.96914
R1063 B.t9 B.n264 2.78796
R1064 B.n567 B.t5 2.78796
R1065 B.n415 B.n320 1.24928
R1066 B.n398 B.n323 1.24928
R1067 B.n155 B.n154 1.24928
R1068 B.n175 B.n174 1.24928
R1069 VN.n5 VN.t7 1621.27
R1070 VN.n1 VN.t0 1621.27
R1071 VN.n12 VN.t6 1621.27
R1072 VN.n8 VN.t3 1621.27
R1073 VN.n4 VN.t2 1582.57
R1074 VN.n2 VN.t1 1582.57
R1075 VN.n11 VN.t5 1582.57
R1076 VN.n9 VN.t4 1582.57
R1077 VN.n8 VN.n7 161.489
R1078 VN.n1 VN.n0 161.489
R1079 VN.n6 VN.n5 161.3
R1080 VN.n13 VN.n12 161.3
R1081 VN.n10 VN.n7 161.3
R1082 VN.n3 VN.n0 161.3
R1083 VN VN.n13 38.8509
R1084 VN.n3 VN.n2 37.246
R1085 VN.n4 VN.n3 37.246
R1086 VN.n11 VN.n10 37.246
R1087 VN.n10 VN.n9 37.246
R1088 VN.n2 VN.n1 35.7853
R1089 VN.n5 VN.n4 35.7853
R1090 VN.n12 VN.n11 35.7853
R1091 VN.n9 VN.n8 35.7853
R1092 VN.n13 VN.n7 0.189894
R1093 VN.n6 VN.n0 0.189894
R1094 VN VN.n6 0.0516364
R1095 VDD2.n2 VDD2.n1 66.3321
R1096 VDD2.n2 VDD2.n0 66.3321
R1097 VDD2 VDD2.n5 66.3293
R1098 VDD2.n4 VDD2.n3 66.1678
R1099 VDD2.n4 VDD2.n2 34.7541
R1100 VDD2.n5 VDD2.t3 1.88442
R1101 VDD2.n5 VDD2.t4 1.88442
R1102 VDD2.n3 VDD2.t1 1.88442
R1103 VDD2.n3 VDD2.t2 1.88442
R1104 VDD2.n1 VDD2.t5 1.88442
R1105 VDD2.n1 VDD2.t0 1.88442
R1106 VDD2.n0 VDD2.t7 1.88442
R1107 VDD2.n0 VDD2.t6 1.88442
R1108 VDD2 VDD2.n4 0.278517
C0 VP VTAIL 1.7594f
C1 VP VN 4.42914f
C2 VP VDD1 2.3052f
C3 VP VDD2 0.261618f
C4 VTAIL VN 1.7453f
C5 VTAIL VDD1 18.0133f
C6 VDD1 VN 0.146814f
C7 VDD2 VTAIL 18.0515f
C8 VDD2 VN 2.19057f
C9 VDD2 VDD1 0.572911f
C10 VDD2 B 2.944451f
C11 VDD1 B 3.109275f
C12 VTAIL B 7.512165f
C13 VN B 6.28599f
C14 VP B 4.495215f
C15 VDD2.t7 B 0.322576f
C16 VDD2.t6 B 0.322576f
C17 VDD2.n0 B 2.85584f
C18 VDD2.t5 B 0.322576f
C19 VDD2.t0 B 0.322576f
C20 VDD2.n1 B 2.85584f
C21 VDD2.n2 B 2.74921f
C22 VDD2.t1 B 0.322576f
C23 VDD2.t2 B 0.322576f
C24 VDD2.n3 B 2.85482f
C25 VDD2.n4 B 3.08959f
C26 VDD2.t3 B 0.322576f
C27 VDD2.t4 B 0.322576f
C28 VDD2.n5 B 2.8558f
C29 VN.n0 B 0.099848f
C30 VN.t2 B 0.251189f
C31 VN.t1 B 0.251189f
C32 VN.t0 B 0.253722f
C33 VN.n1 B 0.119503f
C34 VN.n2 B 0.107712f
C35 VN.n3 B 0.015853f
C36 VN.n4 B 0.107712f
C37 VN.t7 B 0.253722f
C38 VN.n5 B 0.119441f
C39 VN.n6 B 0.036359f
C40 VN.n7 B 0.099848f
C41 VN.t6 B 0.253722f
C42 VN.t5 B 0.251189f
C43 VN.t4 B 0.251189f
C44 VN.t3 B 0.253722f
C45 VN.n8 B 0.119503f
C46 VN.n9 B 0.107712f
C47 VN.n10 B 0.015853f
C48 VN.n11 B 0.107712f
C49 VN.n12 B 0.119441f
C50 VN.n13 B 1.69619f
C51 VDD1.t3 B 0.320313f
C52 VDD1.t1 B 0.320313f
C53 VDD1.n0 B 2.83653f
C54 VDD1.t6 B 0.320313f
C55 VDD1.t7 B 0.320313f
C56 VDD1.n1 B 2.8358f
C57 VDD1.t4 B 0.320313f
C58 VDD1.t5 B 0.320313f
C59 VDD1.n2 B 2.8358f
C60 VDD1.n3 B 2.81302f
C61 VDD1.t2 B 0.320313f
C62 VDD1.t0 B 0.320313f
C63 VDD1.n4 B 2.83478f
C64 VDD1.n5 B 3.11279f
C65 VTAIL.t13 B 0.211785f
C66 VTAIL.t14 B 0.211785f
C67 VTAIL.n0 B 1.8066f
C68 VTAIL.n1 B 0.279692f
C69 VTAIL.t12 B 2.30453f
C70 VTAIL.n2 B 0.393182f
C71 VTAIL.t8 B 2.30453f
C72 VTAIL.n3 B 0.393182f
C73 VTAIL.t5 B 0.211785f
C74 VTAIL.t9 B 0.211785f
C75 VTAIL.n4 B 1.8066f
C76 VTAIL.n5 B 0.311036f
C77 VTAIL.t11 B 2.30453f
C78 VTAIL.n6 B 1.48154f
C79 VTAIL.t2 B 2.30454f
C80 VTAIL.n7 B 1.48154f
C81 VTAIL.t0 B 0.211785f
C82 VTAIL.t1 B 0.211785f
C83 VTAIL.n8 B 1.80661f
C84 VTAIL.n9 B 0.311031f
C85 VTAIL.t15 B 2.30454f
C86 VTAIL.n10 B 0.393176f
C87 VTAIL.t6 B 2.30454f
C88 VTAIL.n11 B 0.393176f
C89 VTAIL.t4 B 0.211785f
C90 VTAIL.t10 B 0.211785f
C91 VTAIL.n12 B 1.80661f
C92 VTAIL.n13 B 0.311031f
C93 VTAIL.t7 B 2.30453f
C94 VTAIL.n14 B 1.48154f
C95 VTAIL.t3 B 2.30453f
C96 VTAIL.n15 B 1.47676f
C97 VP.n0 B 0.048109f
C98 VP.t3 B 0.257569f
C99 VP.t0 B 0.257569f
C100 VP.t1 B 0.260166f
C101 VP.n1 B 0.102383f
C102 VP.t5 B 0.257569f
C103 VP.t6 B 0.257569f
C104 VP.t4 B 0.260166f
C105 VP.n2 B 0.122539f
C106 VP.n3 B 0.110448f
C107 VP.n4 B 0.016256f
C108 VP.n5 B 0.110448f
C109 VP.t7 B 0.260166f
C110 VP.n6 B 0.122475f
C111 VP.n7 B 1.7075f
C112 VP.n8 B 1.75246f
C113 VP.n9 B 0.122475f
C114 VP.n10 B 0.110448f
C115 VP.n11 B 0.016256f
C116 VP.n12 B 0.110448f
C117 VP.t2 B 0.260166f
C118 VP.n13 B 0.122475f
C119 VP.n14 B 0.037283f
.ends

