* NGSPICE file created from diff_pair_sample_1275.ext - technology: sky130A

.subckt diff_pair_sample_1275 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=0 ps=0 w=9.03 l=1.39
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=3.5217 ps=18.84 w=9.03 l=1.39
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=0 ps=0 w=9.03 l=1.39
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=0 ps=0 w=9.03 l=1.39
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=3.5217 ps=18.84 w=9.03 l=1.39
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=0 ps=0 w=9.03 l=1.39
X6 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=3.5217 ps=18.84 w=9.03 l=1.39
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5217 pd=18.84 as=3.5217 ps=18.84 w=9.03 l=1.39
R0 B.n384 B.n79 585
R1 B.n79 B.n36 585
R2 B.n386 B.n385 585
R3 B.n388 B.n78 585
R4 B.n391 B.n390 585
R5 B.n392 B.n77 585
R6 B.n394 B.n393 585
R7 B.n396 B.n76 585
R8 B.n399 B.n398 585
R9 B.n400 B.n75 585
R10 B.n402 B.n401 585
R11 B.n404 B.n74 585
R12 B.n407 B.n406 585
R13 B.n408 B.n73 585
R14 B.n410 B.n409 585
R15 B.n412 B.n72 585
R16 B.n415 B.n414 585
R17 B.n416 B.n71 585
R18 B.n418 B.n417 585
R19 B.n420 B.n70 585
R20 B.n423 B.n422 585
R21 B.n424 B.n69 585
R22 B.n426 B.n425 585
R23 B.n428 B.n68 585
R24 B.n431 B.n430 585
R25 B.n432 B.n67 585
R26 B.n434 B.n433 585
R27 B.n436 B.n66 585
R28 B.n439 B.n438 585
R29 B.n440 B.n65 585
R30 B.n442 B.n441 585
R31 B.n444 B.n64 585
R32 B.n446 B.n445 585
R33 B.n448 B.n447 585
R34 B.n451 B.n450 585
R35 B.n452 B.n59 585
R36 B.n454 B.n453 585
R37 B.n456 B.n58 585
R38 B.n459 B.n458 585
R39 B.n460 B.n57 585
R40 B.n462 B.n461 585
R41 B.n464 B.n56 585
R42 B.n467 B.n466 585
R43 B.n469 B.n53 585
R44 B.n471 B.n470 585
R45 B.n473 B.n52 585
R46 B.n476 B.n475 585
R47 B.n477 B.n51 585
R48 B.n479 B.n478 585
R49 B.n481 B.n50 585
R50 B.n484 B.n483 585
R51 B.n485 B.n49 585
R52 B.n487 B.n486 585
R53 B.n489 B.n48 585
R54 B.n492 B.n491 585
R55 B.n493 B.n47 585
R56 B.n495 B.n494 585
R57 B.n497 B.n46 585
R58 B.n500 B.n499 585
R59 B.n501 B.n45 585
R60 B.n503 B.n502 585
R61 B.n505 B.n44 585
R62 B.n508 B.n507 585
R63 B.n509 B.n43 585
R64 B.n511 B.n510 585
R65 B.n513 B.n42 585
R66 B.n516 B.n515 585
R67 B.n517 B.n41 585
R68 B.n519 B.n518 585
R69 B.n521 B.n40 585
R70 B.n524 B.n523 585
R71 B.n525 B.n39 585
R72 B.n527 B.n526 585
R73 B.n529 B.n38 585
R74 B.n532 B.n531 585
R75 B.n533 B.n37 585
R76 B.n383 B.n35 585
R77 B.n536 B.n35 585
R78 B.n382 B.n34 585
R79 B.n537 B.n34 585
R80 B.n381 B.n33 585
R81 B.n538 B.n33 585
R82 B.n380 B.n379 585
R83 B.n379 B.n29 585
R84 B.n378 B.n28 585
R85 B.n544 B.n28 585
R86 B.n377 B.n27 585
R87 B.n545 B.n27 585
R88 B.n376 B.n26 585
R89 B.n546 B.n26 585
R90 B.n375 B.n374 585
R91 B.n374 B.n22 585
R92 B.n373 B.n21 585
R93 B.n552 B.n21 585
R94 B.n372 B.n20 585
R95 B.n553 B.n20 585
R96 B.n371 B.n19 585
R97 B.n554 B.n19 585
R98 B.n370 B.n369 585
R99 B.n369 B.n15 585
R100 B.n368 B.n14 585
R101 B.n560 B.n14 585
R102 B.n367 B.n13 585
R103 B.n561 B.n13 585
R104 B.n366 B.n12 585
R105 B.n562 B.n12 585
R106 B.n365 B.n364 585
R107 B.n364 B.n8 585
R108 B.n363 B.n7 585
R109 B.n568 B.n7 585
R110 B.n362 B.n6 585
R111 B.n569 B.n6 585
R112 B.n361 B.n5 585
R113 B.n570 B.n5 585
R114 B.n360 B.n359 585
R115 B.n359 B.n4 585
R116 B.n358 B.n80 585
R117 B.n358 B.n357 585
R118 B.n348 B.n81 585
R119 B.n82 B.n81 585
R120 B.n350 B.n349 585
R121 B.n351 B.n350 585
R122 B.n347 B.n86 585
R123 B.n90 B.n86 585
R124 B.n346 B.n345 585
R125 B.n345 B.n344 585
R126 B.n88 B.n87 585
R127 B.n89 B.n88 585
R128 B.n337 B.n336 585
R129 B.n338 B.n337 585
R130 B.n335 B.n95 585
R131 B.n95 B.n94 585
R132 B.n334 B.n333 585
R133 B.n333 B.n332 585
R134 B.n97 B.n96 585
R135 B.n98 B.n97 585
R136 B.n325 B.n324 585
R137 B.n326 B.n325 585
R138 B.n323 B.n102 585
R139 B.n106 B.n102 585
R140 B.n322 B.n321 585
R141 B.n321 B.n320 585
R142 B.n104 B.n103 585
R143 B.n105 B.n104 585
R144 B.n313 B.n312 585
R145 B.n314 B.n313 585
R146 B.n311 B.n111 585
R147 B.n111 B.n110 585
R148 B.n310 B.n309 585
R149 B.n309 B.n308 585
R150 B.n305 B.n115 585
R151 B.n304 B.n303 585
R152 B.n301 B.n116 585
R153 B.n301 B.n114 585
R154 B.n300 B.n299 585
R155 B.n298 B.n297 585
R156 B.n296 B.n118 585
R157 B.n294 B.n293 585
R158 B.n292 B.n119 585
R159 B.n291 B.n290 585
R160 B.n288 B.n120 585
R161 B.n286 B.n285 585
R162 B.n284 B.n121 585
R163 B.n283 B.n282 585
R164 B.n280 B.n122 585
R165 B.n278 B.n277 585
R166 B.n276 B.n123 585
R167 B.n275 B.n274 585
R168 B.n272 B.n124 585
R169 B.n270 B.n269 585
R170 B.n268 B.n125 585
R171 B.n267 B.n266 585
R172 B.n264 B.n126 585
R173 B.n262 B.n261 585
R174 B.n260 B.n127 585
R175 B.n259 B.n258 585
R176 B.n256 B.n128 585
R177 B.n254 B.n253 585
R178 B.n252 B.n129 585
R179 B.n251 B.n250 585
R180 B.n248 B.n130 585
R181 B.n246 B.n245 585
R182 B.n244 B.n131 585
R183 B.n243 B.n242 585
R184 B.n240 B.n239 585
R185 B.n238 B.n237 585
R186 B.n236 B.n136 585
R187 B.n234 B.n233 585
R188 B.n232 B.n137 585
R189 B.n231 B.n230 585
R190 B.n228 B.n138 585
R191 B.n226 B.n225 585
R192 B.n224 B.n139 585
R193 B.n222 B.n221 585
R194 B.n219 B.n142 585
R195 B.n217 B.n216 585
R196 B.n215 B.n143 585
R197 B.n214 B.n213 585
R198 B.n211 B.n144 585
R199 B.n209 B.n208 585
R200 B.n207 B.n145 585
R201 B.n206 B.n205 585
R202 B.n203 B.n146 585
R203 B.n201 B.n200 585
R204 B.n199 B.n147 585
R205 B.n198 B.n197 585
R206 B.n195 B.n148 585
R207 B.n193 B.n192 585
R208 B.n191 B.n149 585
R209 B.n190 B.n189 585
R210 B.n187 B.n150 585
R211 B.n185 B.n184 585
R212 B.n183 B.n151 585
R213 B.n182 B.n181 585
R214 B.n179 B.n152 585
R215 B.n177 B.n176 585
R216 B.n175 B.n153 585
R217 B.n174 B.n173 585
R218 B.n171 B.n154 585
R219 B.n169 B.n168 585
R220 B.n167 B.n155 585
R221 B.n166 B.n165 585
R222 B.n163 B.n156 585
R223 B.n161 B.n160 585
R224 B.n159 B.n158 585
R225 B.n113 B.n112 585
R226 B.n307 B.n306 585
R227 B.n308 B.n307 585
R228 B.n109 B.n108 585
R229 B.n110 B.n109 585
R230 B.n316 B.n315 585
R231 B.n315 B.n314 585
R232 B.n317 B.n107 585
R233 B.n107 B.n105 585
R234 B.n319 B.n318 585
R235 B.n320 B.n319 585
R236 B.n101 B.n100 585
R237 B.n106 B.n101 585
R238 B.n328 B.n327 585
R239 B.n327 B.n326 585
R240 B.n329 B.n99 585
R241 B.n99 B.n98 585
R242 B.n331 B.n330 585
R243 B.n332 B.n331 585
R244 B.n93 B.n92 585
R245 B.n94 B.n93 585
R246 B.n340 B.n339 585
R247 B.n339 B.n338 585
R248 B.n341 B.n91 585
R249 B.n91 B.n89 585
R250 B.n343 B.n342 585
R251 B.n344 B.n343 585
R252 B.n85 B.n84 585
R253 B.n90 B.n85 585
R254 B.n353 B.n352 585
R255 B.n352 B.n351 585
R256 B.n354 B.n83 585
R257 B.n83 B.n82 585
R258 B.n356 B.n355 585
R259 B.n357 B.n356 585
R260 B.n2 B.n0 585
R261 B.n4 B.n2 585
R262 B.n3 B.n1 585
R263 B.n569 B.n3 585
R264 B.n567 B.n566 585
R265 B.n568 B.n567 585
R266 B.n565 B.n9 585
R267 B.n9 B.n8 585
R268 B.n564 B.n563 585
R269 B.n563 B.n562 585
R270 B.n11 B.n10 585
R271 B.n561 B.n11 585
R272 B.n559 B.n558 585
R273 B.n560 B.n559 585
R274 B.n557 B.n16 585
R275 B.n16 B.n15 585
R276 B.n556 B.n555 585
R277 B.n555 B.n554 585
R278 B.n18 B.n17 585
R279 B.n553 B.n18 585
R280 B.n551 B.n550 585
R281 B.n552 B.n551 585
R282 B.n549 B.n23 585
R283 B.n23 B.n22 585
R284 B.n548 B.n547 585
R285 B.n547 B.n546 585
R286 B.n25 B.n24 585
R287 B.n545 B.n25 585
R288 B.n543 B.n542 585
R289 B.n544 B.n543 585
R290 B.n541 B.n30 585
R291 B.n30 B.n29 585
R292 B.n540 B.n539 585
R293 B.n539 B.n538 585
R294 B.n32 B.n31 585
R295 B.n537 B.n32 585
R296 B.n535 B.n534 585
R297 B.n536 B.n535 585
R298 B.n572 B.n571 585
R299 B.n571 B.n570 585
R300 B.n307 B.n115 564.573
R301 B.n535 B.n37 564.573
R302 B.n309 B.n113 564.573
R303 B.n79 B.n35 564.573
R304 B.n140 B.t2 361.57
R305 B.n132 B.t10 361.57
R306 B.n54 B.t13 361.57
R307 B.n60 B.t6 361.57
R308 B.n387 B.n36 256.663
R309 B.n389 B.n36 256.663
R310 B.n395 B.n36 256.663
R311 B.n397 B.n36 256.663
R312 B.n403 B.n36 256.663
R313 B.n405 B.n36 256.663
R314 B.n411 B.n36 256.663
R315 B.n413 B.n36 256.663
R316 B.n419 B.n36 256.663
R317 B.n421 B.n36 256.663
R318 B.n427 B.n36 256.663
R319 B.n429 B.n36 256.663
R320 B.n435 B.n36 256.663
R321 B.n437 B.n36 256.663
R322 B.n443 B.n36 256.663
R323 B.n63 B.n36 256.663
R324 B.n449 B.n36 256.663
R325 B.n455 B.n36 256.663
R326 B.n457 B.n36 256.663
R327 B.n463 B.n36 256.663
R328 B.n465 B.n36 256.663
R329 B.n472 B.n36 256.663
R330 B.n474 B.n36 256.663
R331 B.n480 B.n36 256.663
R332 B.n482 B.n36 256.663
R333 B.n488 B.n36 256.663
R334 B.n490 B.n36 256.663
R335 B.n496 B.n36 256.663
R336 B.n498 B.n36 256.663
R337 B.n504 B.n36 256.663
R338 B.n506 B.n36 256.663
R339 B.n512 B.n36 256.663
R340 B.n514 B.n36 256.663
R341 B.n520 B.n36 256.663
R342 B.n522 B.n36 256.663
R343 B.n528 B.n36 256.663
R344 B.n530 B.n36 256.663
R345 B.n302 B.n114 256.663
R346 B.n117 B.n114 256.663
R347 B.n295 B.n114 256.663
R348 B.n289 B.n114 256.663
R349 B.n287 B.n114 256.663
R350 B.n281 B.n114 256.663
R351 B.n279 B.n114 256.663
R352 B.n273 B.n114 256.663
R353 B.n271 B.n114 256.663
R354 B.n265 B.n114 256.663
R355 B.n263 B.n114 256.663
R356 B.n257 B.n114 256.663
R357 B.n255 B.n114 256.663
R358 B.n249 B.n114 256.663
R359 B.n247 B.n114 256.663
R360 B.n241 B.n114 256.663
R361 B.n135 B.n114 256.663
R362 B.n235 B.n114 256.663
R363 B.n229 B.n114 256.663
R364 B.n227 B.n114 256.663
R365 B.n220 B.n114 256.663
R366 B.n218 B.n114 256.663
R367 B.n212 B.n114 256.663
R368 B.n210 B.n114 256.663
R369 B.n204 B.n114 256.663
R370 B.n202 B.n114 256.663
R371 B.n196 B.n114 256.663
R372 B.n194 B.n114 256.663
R373 B.n188 B.n114 256.663
R374 B.n186 B.n114 256.663
R375 B.n180 B.n114 256.663
R376 B.n178 B.n114 256.663
R377 B.n172 B.n114 256.663
R378 B.n170 B.n114 256.663
R379 B.n164 B.n114 256.663
R380 B.n162 B.n114 256.663
R381 B.n157 B.n114 256.663
R382 B.n307 B.n109 163.367
R383 B.n315 B.n109 163.367
R384 B.n315 B.n107 163.367
R385 B.n319 B.n107 163.367
R386 B.n319 B.n101 163.367
R387 B.n327 B.n101 163.367
R388 B.n327 B.n99 163.367
R389 B.n331 B.n99 163.367
R390 B.n331 B.n93 163.367
R391 B.n339 B.n93 163.367
R392 B.n339 B.n91 163.367
R393 B.n343 B.n91 163.367
R394 B.n343 B.n85 163.367
R395 B.n352 B.n85 163.367
R396 B.n352 B.n83 163.367
R397 B.n356 B.n83 163.367
R398 B.n356 B.n2 163.367
R399 B.n571 B.n2 163.367
R400 B.n571 B.n3 163.367
R401 B.n567 B.n3 163.367
R402 B.n567 B.n9 163.367
R403 B.n563 B.n9 163.367
R404 B.n563 B.n11 163.367
R405 B.n559 B.n11 163.367
R406 B.n559 B.n16 163.367
R407 B.n555 B.n16 163.367
R408 B.n555 B.n18 163.367
R409 B.n551 B.n18 163.367
R410 B.n551 B.n23 163.367
R411 B.n547 B.n23 163.367
R412 B.n547 B.n25 163.367
R413 B.n543 B.n25 163.367
R414 B.n543 B.n30 163.367
R415 B.n539 B.n30 163.367
R416 B.n539 B.n32 163.367
R417 B.n535 B.n32 163.367
R418 B.n303 B.n301 163.367
R419 B.n301 B.n300 163.367
R420 B.n297 B.n296 163.367
R421 B.n294 B.n119 163.367
R422 B.n290 B.n288 163.367
R423 B.n286 B.n121 163.367
R424 B.n282 B.n280 163.367
R425 B.n278 B.n123 163.367
R426 B.n274 B.n272 163.367
R427 B.n270 B.n125 163.367
R428 B.n266 B.n264 163.367
R429 B.n262 B.n127 163.367
R430 B.n258 B.n256 163.367
R431 B.n254 B.n129 163.367
R432 B.n250 B.n248 163.367
R433 B.n246 B.n131 163.367
R434 B.n242 B.n240 163.367
R435 B.n237 B.n236 163.367
R436 B.n234 B.n137 163.367
R437 B.n230 B.n228 163.367
R438 B.n226 B.n139 163.367
R439 B.n221 B.n219 163.367
R440 B.n217 B.n143 163.367
R441 B.n213 B.n211 163.367
R442 B.n209 B.n145 163.367
R443 B.n205 B.n203 163.367
R444 B.n201 B.n147 163.367
R445 B.n197 B.n195 163.367
R446 B.n193 B.n149 163.367
R447 B.n189 B.n187 163.367
R448 B.n185 B.n151 163.367
R449 B.n181 B.n179 163.367
R450 B.n177 B.n153 163.367
R451 B.n173 B.n171 163.367
R452 B.n169 B.n155 163.367
R453 B.n165 B.n163 163.367
R454 B.n161 B.n158 163.367
R455 B.n309 B.n111 163.367
R456 B.n313 B.n111 163.367
R457 B.n313 B.n104 163.367
R458 B.n321 B.n104 163.367
R459 B.n321 B.n102 163.367
R460 B.n325 B.n102 163.367
R461 B.n325 B.n97 163.367
R462 B.n333 B.n97 163.367
R463 B.n333 B.n95 163.367
R464 B.n337 B.n95 163.367
R465 B.n337 B.n88 163.367
R466 B.n345 B.n88 163.367
R467 B.n345 B.n86 163.367
R468 B.n350 B.n86 163.367
R469 B.n350 B.n81 163.367
R470 B.n358 B.n81 163.367
R471 B.n359 B.n358 163.367
R472 B.n359 B.n5 163.367
R473 B.n6 B.n5 163.367
R474 B.n7 B.n6 163.367
R475 B.n364 B.n7 163.367
R476 B.n364 B.n12 163.367
R477 B.n13 B.n12 163.367
R478 B.n14 B.n13 163.367
R479 B.n369 B.n14 163.367
R480 B.n369 B.n19 163.367
R481 B.n20 B.n19 163.367
R482 B.n21 B.n20 163.367
R483 B.n374 B.n21 163.367
R484 B.n374 B.n26 163.367
R485 B.n27 B.n26 163.367
R486 B.n28 B.n27 163.367
R487 B.n379 B.n28 163.367
R488 B.n379 B.n33 163.367
R489 B.n34 B.n33 163.367
R490 B.n35 B.n34 163.367
R491 B.n531 B.n529 163.367
R492 B.n527 B.n39 163.367
R493 B.n523 B.n521 163.367
R494 B.n519 B.n41 163.367
R495 B.n515 B.n513 163.367
R496 B.n511 B.n43 163.367
R497 B.n507 B.n505 163.367
R498 B.n503 B.n45 163.367
R499 B.n499 B.n497 163.367
R500 B.n495 B.n47 163.367
R501 B.n491 B.n489 163.367
R502 B.n487 B.n49 163.367
R503 B.n483 B.n481 163.367
R504 B.n479 B.n51 163.367
R505 B.n475 B.n473 163.367
R506 B.n471 B.n53 163.367
R507 B.n466 B.n464 163.367
R508 B.n462 B.n57 163.367
R509 B.n458 B.n456 163.367
R510 B.n454 B.n59 163.367
R511 B.n450 B.n448 163.367
R512 B.n445 B.n444 163.367
R513 B.n442 B.n65 163.367
R514 B.n438 B.n436 163.367
R515 B.n434 B.n67 163.367
R516 B.n430 B.n428 163.367
R517 B.n426 B.n69 163.367
R518 B.n422 B.n420 163.367
R519 B.n418 B.n71 163.367
R520 B.n414 B.n412 163.367
R521 B.n410 B.n73 163.367
R522 B.n406 B.n404 163.367
R523 B.n402 B.n75 163.367
R524 B.n398 B.n396 163.367
R525 B.n394 B.n77 163.367
R526 B.n390 B.n388 163.367
R527 B.n386 B.n79 163.367
R528 B.n308 B.n114 106.886
R529 B.n536 B.n36 106.886
R530 B.n140 B.t5 105.371
R531 B.n60 B.t8 105.371
R532 B.n132 B.t12 105.359
R533 B.n54 B.t14 105.359
R534 B.n141 B.t4 72.0131
R535 B.n61 B.t9 72.0131
R536 B.n133 B.t11 72.0024
R537 B.n55 B.t15 72.0024
R538 B.n302 B.n115 71.676
R539 B.n300 B.n117 71.676
R540 B.n296 B.n295 71.676
R541 B.n289 B.n119 71.676
R542 B.n288 B.n287 71.676
R543 B.n281 B.n121 71.676
R544 B.n280 B.n279 71.676
R545 B.n273 B.n123 71.676
R546 B.n272 B.n271 71.676
R547 B.n265 B.n125 71.676
R548 B.n264 B.n263 71.676
R549 B.n257 B.n127 71.676
R550 B.n256 B.n255 71.676
R551 B.n249 B.n129 71.676
R552 B.n248 B.n247 71.676
R553 B.n241 B.n131 71.676
R554 B.n240 B.n135 71.676
R555 B.n236 B.n235 71.676
R556 B.n229 B.n137 71.676
R557 B.n228 B.n227 71.676
R558 B.n220 B.n139 71.676
R559 B.n219 B.n218 71.676
R560 B.n212 B.n143 71.676
R561 B.n211 B.n210 71.676
R562 B.n204 B.n145 71.676
R563 B.n203 B.n202 71.676
R564 B.n196 B.n147 71.676
R565 B.n195 B.n194 71.676
R566 B.n188 B.n149 71.676
R567 B.n187 B.n186 71.676
R568 B.n180 B.n151 71.676
R569 B.n179 B.n178 71.676
R570 B.n172 B.n153 71.676
R571 B.n171 B.n170 71.676
R572 B.n164 B.n155 71.676
R573 B.n163 B.n162 71.676
R574 B.n158 B.n157 71.676
R575 B.n530 B.n37 71.676
R576 B.n529 B.n528 71.676
R577 B.n522 B.n39 71.676
R578 B.n521 B.n520 71.676
R579 B.n514 B.n41 71.676
R580 B.n513 B.n512 71.676
R581 B.n506 B.n43 71.676
R582 B.n505 B.n504 71.676
R583 B.n498 B.n45 71.676
R584 B.n497 B.n496 71.676
R585 B.n490 B.n47 71.676
R586 B.n489 B.n488 71.676
R587 B.n482 B.n49 71.676
R588 B.n481 B.n480 71.676
R589 B.n474 B.n51 71.676
R590 B.n473 B.n472 71.676
R591 B.n465 B.n53 71.676
R592 B.n464 B.n463 71.676
R593 B.n457 B.n57 71.676
R594 B.n456 B.n455 71.676
R595 B.n449 B.n59 71.676
R596 B.n448 B.n63 71.676
R597 B.n444 B.n443 71.676
R598 B.n437 B.n65 71.676
R599 B.n436 B.n435 71.676
R600 B.n429 B.n67 71.676
R601 B.n428 B.n427 71.676
R602 B.n421 B.n69 71.676
R603 B.n420 B.n419 71.676
R604 B.n413 B.n71 71.676
R605 B.n412 B.n411 71.676
R606 B.n405 B.n73 71.676
R607 B.n404 B.n403 71.676
R608 B.n397 B.n75 71.676
R609 B.n396 B.n395 71.676
R610 B.n389 B.n77 71.676
R611 B.n388 B.n387 71.676
R612 B.n387 B.n386 71.676
R613 B.n390 B.n389 71.676
R614 B.n395 B.n394 71.676
R615 B.n398 B.n397 71.676
R616 B.n403 B.n402 71.676
R617 B.n406 B.n405 71.676
R618 B.n411 B.n410 71.676
R619 B.n414 B.n413 71.676
R620 B.n419 B.n418 71.676
R621 B.n422 B.n421 71.676
R622 B.n427 B.n426 71.676
R623 B.n430 B.n429 71.676
R624 B.n435 B.n434 71.676
R625 B.n438 B.n437 71.676
R626 B.n443 B.n442 71.676
R627 B.n445 B.n63 71.676
R628 B.n450 B.n449 71.676
R629 B.n455 B.n454 71.676
R630 B.n458 B.n457 71.676
R631 B.n463 B.n462 71.676
R632 B.n466 B.n465 71.676
R633 B.n472 B.n471 71.676
R634 B.n475 B.n474 71.676
R635 B.n480 B.n479 71.676
R636 B.n483 B.n482 71.676
R637 B.n488 B.n487 71.676
R638 B.n491 B.n490 71.676
R639 B.n496 B.n495 71.676
R640 B.n499 B.n498 71.676
R641 B.n504 B.n503 71.676
R642 B.n507 B.n506 71.676
R643 B.n512 B.n511 71.676
R644 B.n515 B.n514 71.676
R645 B.n520 B.n519 71.676
R646 B.n523 B.n522 71.676
R647 B.n528 B.n527 71.676
R648 B.n531 B.n530 71.676
R649 B.n303 B.n302 71.676
R650 B.n297 B.n117 71.676
R651 B.n295 B.n294 71.676
R652 B.n290 B.n289 71.676
R653 B.n287 B.n286 71.676
R654 B.n282 B.n281 71.676
R655 B.n279 B.n278 71.676
R656 B.n274 B.n273 71.676
R657 B.n271 B.n270 71.676
R658 B.n266 B.n265 71.676
R659 B.n263 B.n262 71.676
R660 B.n258 B.n257 71.676
R661 B.n255 B.n254 71.676
R662 B.n250 B.n249 71.676
R663 B.n247 B.n246 71.676
R664 B.n242 B.n241 71.676
R665 B.n237 B.n135 71.676
R666 B.n235 B.n234 71.676
R667 B.n230 B.n229 71.676
R668 B.n227 B.n226 71.676
R669 B.n221 B.n220 71.676
R670 B.n218 B.n217 71.676
R671 B.n213 B.n212 71.676
R672 B.n210 B.n209 71.676
R673 B.n205 B.n204 71.676
R674 B.n202 B.n201 71.676
R675 B.n197 B.n196 71.676
R676 B.n194 B.n193 71.676
R677 B.n189 B.n188 71.676
R678 B.n186 B.n185 71.676
R679 B.n181 B.n180 71.676
R680 B.n178 B.n177 71.676
R681 B.n173 B.n172 71.676
R682 B.n170 B.n169 71.676
R683 B.n165 B.n164 71.676
R684 B.n162 B.n161 71.676
R685 B.n157 B.n113 71.676
R686 B.n223 B.n141 59.5399
R687 B.n134 B.n133 59.5399
R688 B.n468 B.n55 59.5399
R689 B.n62 B.n61 59.5399
R690 B.n308 B.n110 52.2899
R691 B.n314 B.n110 52.2899
R692 B.n314 B.n105 52.2899
R693 B.n320 B.n105 52.2899
R694 B.n320 B.n106 52.2899
R695 B.n326 B.n98 52.2899
R696 B.n332 B.n98 52.2899
R697 B.n332 B.n94 52.2899
R698 B.n338 B.n94 52.2899
R699 B.n338 B.n89 52.2899
R700 B.n344 B.n89 52.2899
R701 B.n344 B.n90 52.2899
R702 B.n351 B.n82 52.2899
R703 B.n357 B.n82 52.2899
R704 B.n357 B.n4 52.2899
R705 B.n570 B.n4 52.2899
R706 B.n570 B.n569 52.2899
R707 B.n569 B.n568 52.2899
R708 B.n568 B.n8 52.2899
R709 B.n562 B.n8 52.2899
R710 B.n561 B.n560 52.2899
R711 B.n560 B.n15 52.2899
R712 B.n554 B.n15 52.2899
R713 B.n554 B.n553 52.2899
R714 B.n553 B.n552 52.2899
R715 B.n552 B.n22 52.2899
R716 B.n546 B.n22 52.2899
R717 B.n545 B.n544 52.2899
R718 B.n544 B.n29 52.2899
R719 B.n538 B.n29 52.2899
R720 B.n538 B.n537 52.2899
R721 B.n537 B.n536 52.2899
R722 B.n90 B.t0 45.3693
R723 B.t1 B.n561 45.3693
R724 B.n534 B.n533 36.6834
R725 B.n384 B.n383 36.6834
R726 B.n310 B.n112 36.6834
R727 B.n306 B.n305 36.6834
R728 B.n141 B.n140 33.3581
R729 B.n133 B.n132 33.3581
R730 B.n55 B.n54 33.3581
R731 B.n61 B.n60 33.3581
R732 B.n106 B.t3 31.5279
R733 B.t7 B.n545 31.5279
R734 B.n326 B.t3 20.7625
R735 B.n546 B.t7 20.7625
R736 B B.n572 18.0485
R737 B.n533 B.n532 10.6151
R738 B.n532 B.n38 10.6151
R739 B.n526 B.n38 10.6151
R740 B.n526 B.n525 10.6151
R741 B.n525 B.n524 10.6151
R742 B.n524 B.n40 10.6151
R743 B.n518 B.n40 10.6151
R744 B.n518 B.n517 10.6151
R745 B.n517 B.n516 10.6151
R746 B.n516 B.n42 10.6151
R747 B.n510 B.n42 10.6151
R748 B.n510 B.n509 10.6151
R749 B.n509 B.n508 10.6151
R750 B.n508 B.n44 10.6151
R751 B.n502 B.n44 10.6151
R752 B.n502 B.n501 10.6151
R753 B.n501 B.n500 10.6151
R754 B.n500 B.n46 10.6151
R755 B.n494 B.n46 10.6151
R756 B.n494 B.n493 10.6151
R757 B.n493 B.n492 10.6151
R758 B.n492 B.n48 10.6151
R759 B.n486 B.n48 10.6151
R760 B.n486 B.n485 10.6151
R761 B.n485 B.n484 10.6151
R762 B.n484 B.n50 10.6151
R763 B.n478 B.n50 10.6151
R764 B.n478 B.n477 10.6151
R765 B.n477 B.n476 10.6151
R766 B.n476 B.n52 10.6151
R767 B.n470 B.n52 10.6151
R768 B.n470 B.n469 10.6151
R769 B.n467 B.n56 10.6151
R770 B.n461 B.n56 10.6151
R771 B.n461 B.n460 10.6151
R772 B.n460 B.n459 10.6151
R773 B.n459 B.n58 10.6151
R774 B.n453 B.n58 10.6151
R775 B.n453 B.n452 10.6151
R776 B.n452 B.n451 10.6151
R777 B.n447 B.n446 10.6151
R778 B.n446 B.n64 10.6151
R779 B.n441 B.n64 10.6151
R780 B.n441 B.n440 10.6151
R781 B.n440 B.n439 10.6151
R782 B.n439 B.n66 10.6151
R783 B.n433 B.n66 10.6151
R784 B.n433 B.n432 10.6151
R785 B.n432 B.n431 10.6151
R786 B.n431 B.n68 10.6151
R787 B.n425 B.n68 10.6151
R788 B.n425 B.n424 10.6151
R789 B.n424 B.n423 10.6151
R790 B.n423 B.n70 10.6151
R791 B.n417 B.n70 10.6151
R792 B.n417 B.n416 10.6151
R793 B.n416 B.n415 10.6151
R794 B.n415 B.n72 10.6151
R795 B.n409 B.n72 10.6151
R796 B.n409 B.n408 10.6151
R797 B.n408 B.n407 10.6151
R798 B.n407 B.n74 10.6151
R799 B.n401 B.n74 10.6151
R800 B.n401 B.n400 10.6151
R801 B.n400 B.n399 10.6151
R802 B.n399 B.n76 10.6151
R803 B.n393 B.n76 10.6151
R804 B.n393 B.n392 10.6151
R805 B.n392 B.n391 10.6151
R806 B.n391 B.n78 10.6151
R807 B.n385 B.n78 10.6151
R808 B.n385 B.n384 10.6151
R809 B.n311 B.n310 10.6151
R810 B.n312 B.n311 10.6151
R811 B.n312 B.n103 10.6151
R812 B.n322 B.n103 10.6151
R813 B.n323 B.n322 10.6151
R814 B.n324 B.n323 10.6151
R815 B.n324 B.n96 10.6151
R816 B.n334 B.n96 10.6151
R817 B.n335 B.n334 10.6151
R818 B.n336 B.n335 10.6151
R819 B.n336 B.n87 10.6151
R820 B.n346 B.n87 10.6151
R821 B.n347 B.n346 10.6151
R822 B.n349 B.n347 10.6151
R823 B.n349 B.n348 10.6151
R824 B.n348 B.n80 10.6151
R825 B.n360 B.n80 10.6151
R826 B.n361 B.n360 10.6151
R827 B.n362 B.n361 10.6151
R828 B.n363 B.n362 10.6151
R829 B.n365 B.n363 10.6151
R830 B.n366 B.n365 10.6151
R831 B.n367 B.n366 10.6151
R832 B.n368 B.n367 10.6151
R833 B.n370 B.n368 10.6151
R834 B.n371 B.n370 10.6151
R835 B.n372 B.n371 10.6151
R836 B.n373 B.n372 10.6151
R837 B.n375 B.n373 10.6151
R838 B.n376 B.n375 10.6151
R839 B.n377 B.n376 10.6151
R840 B.n378 B.n377 10.6151
R841 B.n380 B.n378 10.6151
R842 B.n381 B.n380 10.6151
R843 B.n382 B.n381 10.6151
R844 B.n383 B.n382 10.6151
R845 B.n305 B.n304 10.6151
R846 B.n304 B.n116 10.6151
R847 B.n299 B.n116 10.6151
R848 B.n299 B.n298 10.6151
R849 B.n298 B.n118 10.6151
R850 B.n293 B.n118 10.6151
R851 B.n293 B.n292 10.6151
R852 B.n292 B.n291 10.6151
R853 B.n291 B.n120 10.6151
R854 B.n285 B.n120 10.6151
R855 B.n285 B.n284 10.6151
R856 B.n284 B.n283 10.6151
R857 B.n283 B.n122 10.6151
R858 B.n277 B.n122 10.6151
R859 B.n277 B.n276 10.6151
R860 B.n276 B.n275 10.6151
R861 B.n275 B.n124 10.6151
R862 B.n269 B.n124 10.6151
R863 B.n269 B.n268 10.6151
R864 B.n268 B.n267 10.6151
R865 B.n267 B.n126 10.6151
R866 B.n261 B.n126 10.6151
R867 B.n261 B.n260 10.6151
R868 B.n260 B.n259 10.6151
R869 B.n259 B.n128 10.6151
R870 B.n253 B.n128 10.6151
R871 B.n253 B.n252 10.6151
R872 B.n252 B.n251 10.6151
R873 B.n251 B.n130 10.6151
R874 B.n245 B.n130 10.6151
R875 B.n245 B.n244 10.6151
R876 B.n244 B.n243 10.6151
R877 B.n239 B.n238 10.6151
R878 B.n238 B.n136 10.6151
R879 B.n233 B.n136 10.6151
R880 B.n233 B.n232 10.6151
R881 B.n232 B.n231 10.6151
R882 B.n231 B.n138 10.6151
R883 B.n225 B.n138 10.6151
R884 B.n225 B.n224 10.6151
R885 B.n222 B.n142 10.6151
R886 B.n216 B.n142 10.6151
R887 B.n216 B.n215 10.6151
R888 B.n215 B.n214 10.6151
R889 B.n214 B.n144 10.6151
R890 B.n208 B.n144 10.6151
R891 B.n208 B.n207 10.6151
R892 B.n207 B.n206 10.6151
R893 B.n206 B.n146 10.6151
R894 B.n200 B.n146 10.6151
R895 B.n200 B.n199 10.6151
R896 B.n199 B.n198 10.6151
R897 B.n198 B.n148 10.6151
R898 B.n192 B.n148 10.6151
R899 B.n192 B.n191 10.6151
R900 B.n191 B.n190 10.6151
R901 B.n190 B.n150 10.6151
R902 B.n184 B.n150 10.6151
R903 B.n184 B.n183 10.6151
R904 B.n183 B.n182 10.6151
R905 B.n182 B.n152 10.6151
R906 B.n176 B.n152 10.6151
R907 B.n176 B.n175 10.6151
R908 B.n175 B.n174 10.6151
R909 B.n174 B.n154 10.6151
R910 B.n168 B.n154 10.6151
R911 B.n168 B.n167 10.6151
R912 B.n167 B.n166 10.6151
R913 B.n166 B.n156 10.6151
R914 B.n160 B.n156 10.6151
R915 B.n160 B.n159 10.6151
R916 B.n159 B.n112 10.6151
R917 B.n306 B.n108 10.6151
R918 B.n316 B.n108 10.6151
R919 B.n317 B.n316 10.6151
R920 B.n318 B.n317 10.6151
R921 B.n318 B.n100 10.6151
R922 B.n328 B.n100 10.6151
R923 B.n329 B.n328 10.6151
R924 B.n330 B.n329 10.6151
R925 B.n330 B.n92 10.6151
R926 B.n340 B.n92 10.6151
R927 B.n341 B.n340 10.6151
R928 B.n342 B.n341 10.6151
R929 B.n342 B.n84 10.6151
R930 B.n353 B.n84 10.6151
R931 B.n354 B.n353 10.6151
R932 B.n355 B.n354 10.6151
R933 B.n355 B.n0 10.6151
R934 B.n566 B.n1 10.6151
R935 B.n566 B.n565 10.6151
R936 B.n565 B.n564 10.6151
R937 B.n564 B.n10 10.6151
R938 B.n558 B.n10 10.6151
R939 B.n558 B.n557 10.6151
R940 B.n557 B.n556 10.6151
R941 B.n556 B.n17 10.6151
R942 B.n550 B.n17 10.6151
R943 B.n550 B.n549 10.6151
R944 B.n549 B.n548 10.6151
R945 B.n548 B.n24 10.6151
R946 B.n542 B.n24 10.6151
R947 B.n542 B.n541 10.6151
R948 B.n541 B.n540 10.6151
R949 B.n540 B.n31 10.6151
R950 B.n534 B.n31 10.6151
R951 B.n351 B.t0 6.92116
R952 B.n562 B.t1 6.92116
R953 B.n468 B.n467 6.5566
R954 B.n451 B.n62 6.5566
R955 B.n239 B.n134 6.5566
R956 B.n224 B.n223 6.5566
R957 B.n469 B.n468 4.05904
R958 B.n447 B.n62 4.05904
R959 B.n243 B.n134 4.05904
R960 B.n223 B.n222 4.05904
R961 B.n572 B.n0 2.81026
R962 B.n572 B.n1 2.81026
R963 VN VN.t1 305.084
R964 VN VN.t0 265.748
R965 VTAIL.n1 VTAIL.t3 51.6333
R966 VTAIL.n3 VTAIL.t2 51.6331
R967 VTAIL.n0 VTAIL.t1 51.6331
R968 VTAIL.n2 VTAIL.t0 51.6331
R969 VTAIL.n1 VTAIL.n0 23.1169
R970 VTAIL.n3 VTAIL.n2 21.6341
R971 VTAIL.n2 VTAIL.n1 1.21171
R972 VTAIL VTAIL.n0 0.899207
R973 VTAIL VTAIL.n3 0.313
R974 VDD2.n0 VDD2.t1 102.722
R975 VDD2.n0 VDD2.t0 68.3118
R976 VDD2 VDD2.n0 0.429379
R977 VP.n0 VP.t1 304.8
R978 VP.n0 VP.t0 265.601
R979 VP VP.n0 0.146778
R980 VDD1 VDD1.t1 103.617
R981 VDD1 VDD1.t0 68.7407
C0 VDD1 VP 2.03608f
C1 VDD1 VN 0.147567f
C2 VN VP 4.33709f
C3 VTAIL VDD2 4.23916f
C4 VDD1 VDD2 0.53339f
C5 VDD1 VTAIL 4.19744f
C6 VDD2 VP 0.282048f
C7 VDD2 VN 1.90426f
C8 VTAIL VP 1.6301f
C9 VTAIL VN 1.61574f
C10 VDD2 B 3.445639f
C11 VDD1 B 6.08676f
C12 VTAIL B 5.54719f
C13 VN B 6.95344f
C14 VP B 4.677186f
C15 VDD1.t0 B 1.62074f
C16 VDD1.t1 B 2.03795f
C17 VP.t1 B 1.65389f
C18 VP.t0 B 1.43549f
C19 VP.n0 B 3.17625f
C20 VDD2.t1 B 1.37968f
C21 VDD2.t0 B 1.11034f
C22 VDD2.n0 B 1.65692f
C23 VTAIL.t1 B 1.15735f
C24 VTAIL.n0 B 0.963635f
C25 VTAIL.t3 B 1.15736f
C26 VTAIL.n1 B 0.978924f
C27 VTAIL.t0 B 1.15735f
C28 VTAIL.n2 B 0.906369f
C29 VTAIL.t2 B 1.15735f
C30 VTAIL.n3 B 0.862392f
C31 VN.t0 B 0.972241f
C32 VN.t1 B 1.12269f
.ends

