* NGSPICE file created from diff_pair_sample_0719.ext - technology: sky130A

.subckt diff_pair_sample_0719 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.24
X1 VTAIL.t8 VP.t1 VDD1.t4 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=3.0492 ps=18.81 w=18.48 l=0.24
X2 VDD1.t3 VP.t2 VTAIL.t10 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.24
X3 VDD2.t5 VN.t0 VTAIL.t2 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.24
X4 VDD2.t4 VN.t1 VTAIL.t1 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.24
X5 VDD1.t2 VP.t3 VTAIL.t6 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.24
X6 VDD2.t3 VN.t2 VTAIL.t0 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=7.2072 ps=37.74 w=18.48 l=0.24
X7 VTAIL.t5 VN.t3 VDD2.t2 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=3.0492 ps=18.81 w=18.48 l=0.24
X8 B.t11 B.t9 B.t10 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.24
X9 VDD2.t1 VN.t4 VTAIL.t4 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.24
X10 VDD1.t1 VP.t4 VTAIL.t7 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=3.0492 ps=18.81 w=18.48 l=0.24
X11 B.t8 B.t6 B.t7 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.24
X12 B.t5 B.t3 B.t4 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.24
X13 VTAIL.t11 VP.t5 VDD1.t0 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=3.0492 ps=18.81 w=18.48 l=0.24
X14 VTAIL.t3 VN.t5 VDD2.t0 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=3.0492 pd=18.81 as=3.0492 ps=18.81 w=18.48 l=0.24
X15 B.t2 B.t0 B.t1 w_n1426_n4664# sky130_fd_pr__pfet_01v8 ad=7.2072 pd=37.74 as=0 ps=0 w=18.48 l=0.24
R0 VP.n7 VP.t3 2032.98
R1 VP.n5 VP.t0 2032.98
R2 VP.n0 VP.t4 2032.98
R3 VP.n2 VP.t2 2032.98
R4 VP.n6 VP.t5 1986.24
R5 VP.n1 VP.t1 1986.24
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n4 VP.n3 44.4134
R11 VP.n6 VP.n5 36.5157
R12 VP.n7 VP.n6 36.5157
R13 VP.n1 VP.n0 36.5157
R14 VP.n2 VP.n1 36.5157
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VTAIL.n7 VTAIL.t0 51.2853
R18 VTAIL.n11 VTAIL.t1 51.2852
R19 VTAIL.n2 VTAIL.t6 51.2852
R20 VTAIL.n10 VTAIL.t10 51.2852
R21 VTAIL.n9 VTAIL.n8 49.5265
R22 VTAIL.n6 VTAIL.n5 49.5265
R23 VTAIL.n1 VTAIL.n0 49.5262
R24 VTAIL.n4 VTAIL.n3 49.5262
R25 VTAIL.n6 VTAIL.n4 29.2807
R26 VTAIL.n11 VTAIL.n10 28.7893
R27 VTAIL.n0 VTAIL.t2 1.75943
R28 VTAIL.n0 VTAIL.t3 1.75943
R29 VTAIL.n3 VTAIL.t9 1.75943
R30 VTAIL.n3 VTAIL.t11 1.75943
R31 VTAIL.n8 VTAIL.t7 1.75943
R32 VTAIL.n8 VTAIL.t8 1.75943
R33 VTAIL.n5 VTAIL.t4 1.75943
R34 VTAIL.n5 VTAIL.t5 1.75943
R35 VTAIL.n9 VTAIL.n7 0.716017
R36 VTAIL.n2 VTAIL.n1 0.716017
R37 VTAIL.n7 VTAIL.n6 0.491879
R38 VTAIL.n10 VTAIL.n9 0.491879
R39 VTAIL.n4 VTAIL.n2 0.491879
R40 VTAIL VTAIL.n11 0.310845
R41 VTAIL VTAIL.n1 0.181534
R42 VDD1 VDD1.t1 68.3909
R43 VDD1.n1 VDD1.t5 68.2772
R44 VDD1.n1 VDD1.n0 66.2725
R45 VDD1.n3 VDD1.n2 66.2051
R46 VDD1.n3 VDD1.n1 42.072
R47 VDD1.n2 VDD1.t4 1.75943
R48 VDD1.n2 VDD1.t3 1.75943
R49 VDD1.n0 VDD1.t0 1.75943
R50 VDD1.n0 VDD1.t2 1.75943
R51 VDD1 VDD1.n3 0.0651552
R52 VN.n2 VN.t1 2032.98
R53 VN.n0 VN.t0 2032.98
R54 VN.n6 VN.t4 2032.98
R55 VN.n4 VN.t2 2032.98
R56 VN.n1 VN.t5 1986.24
R57 VN.n5 VN.t3 1986.24
R58 VN.n7 VN.n4 161.489
R59 VN.n3 VN.n0 161.489
R60 VN.n3 VN.n2 161.3
R61 VN.n7 VN.n6 161.3
R62 VN VN.n7 44.7941
R63 VN.n1 VN.n0 36.5157
R64 VN.n2 VN.n1 36.5157
R65 VN.n6 VN.n5 36.5157
R66 VN.n5 VN.n4 36.5157
R67 VN VN.n3 0.0516364
R68 VDD2.n1 VDD2.t5 68.2772
R69 VDD2.n2 VDD2.t1 67.9641
R70 VDD2.n1 VDD2.n0 66.2725
R71 VDD2 VDD2.n3 66.2697
R72 VDD2.n2 VDD2.n1 41.2433
R73 VDD2.n3 VDD2.t2 1.75943
R74 VDD2.n3 VDD2.t3 1.75943
R75 VDD2.n0 VDD2.t0 1.75943
R76 VDD2.n0 VDD2.t4 1.75943
R77 VDD2 VDD2.n2 0.427224
R78 B.n126 B.t3 2082.01
R79 B.n132 B.t9 2082.01
R80 B.n40 B.t0 2082.01
R81 B.n48 B.t6 2082.01
R82 B.n438 B.n79 585
R83 B.n440 B.n439 585
R84 B.n441 B.n78 585
R85 B.n443 B.n442 585
R86 B.n444 B.n77 585
R87 B.n446 B.n445 585
R88 B.n447 B.n76 585
R89 B.n449 B.n448 585
R90 B.n450 B.n75 585
R91 B.n452 B.n451 585
R92 B.n453 B.n74 585
R93 B.n455 B.n454 585
R94 B.n456 B.n73 585
R95 B.n458 B.n457 585
R96 B.n459 B.n72 585
R97 B.n461 B.n460 585
R98 B.n462 B.n71 585
R99 B.n464 B.n463 585
R100 B.n465 B.n70 585
R101 B.n467 B.n466 585
R102 B.n468 B.n69 585
R103 B.n470 B.n469 585
R104 B.n471 B.n68 585
R105 B.n473 B.n472 585
R106 B.n474 B.n67 585
R107 B.n476 B.n475 585
R108 B.n477 B.n66 585
R109 B.n479 B.n478 585
R110 B.n480 B.n65 585
R111 B.n482 B.n481 585
R112 B.n483 B.n64 585
R113 B.n485 B.n484 585
R114 B.n486 B.n63 585
R115 B.n488 B.n487 585
R116 B.n489 B.n62 585
R117 B.n491 B.n490 585
R118 B.n492 B.n61 585
R119 B.n494 B.n493 585
R120 B.n495 B.n60 585
R121 B.n497 B.n496 585
R122 B.n498 B.n59 585
R123 B.n500 B.n499 585
R124 B.n501 B.n58 585
R125 B.n503 B.n502 585
R126 B.n504 B.n57 585
R127 B.n506 B.n505 585
R128 B.n507 B.n56 585
R129 B.n509 B.n508 585
R130 B.n510 B.n55 585
R131 B.n512 B.n511 585
R132 B.n513 B.n54 585
R133 B.n515 B.n514 585
R134 B.n516 B.n53 585
R135 B.n518 B.n517 585
R136 B.n519 B.n52 585
R137 B.n521 B.n520 585
R138 B.n522 B.n51 585
R139 B.n524 B.n523 585
R140 B.n525 B.n50 585
R141 B.n527 B.n526 585
R142 B.n528 B.n47 585
R143 B.n531 B.n530 585
R144 B.n532 B.n46 585
R145 B.n534 B.n533 585
R146 B.n535 B.n45 585
R147 B.n537 B.n536 585
R148 B.n538 B.n44 585
R149 B.n540 B.n539 585
R150 B.n541 B.n43 585
R151 B.n543 B.n542 585
R152 B.n545 B.n544 585
R153 B.n546 B.n39 585
R154 B.n548 B.n547 585
R155 B.n549 B.n38 585
R156 B.n551 B.n550 585
R157 B.n552 B.n37 585
R158 B.n554 B.n553 585
R159 B.n555 B.n36 585
R160 B.n557 B.n556 585
R161 B.n558 B.n35 585
R162 B.n560 B.n559 585
R163 B.n561 B.n34 585
R164 B.n563 B.n562 585
R165 B.n564 B.n33 585
R166 B.n566 B.n565 585
R167 B.n567 B.n32 585
R168 B.n569 B.n568 585
R169 B.n570 B.n31 585
R170 B.n572 B.n571 585
R171 B.n573 B.n30 585
R172 B.n575 B.n574 585
R173 B.n576 B.n29 585
R174 B.n578 B.n577 585
R175 B.n579 B.n28 585
R176 B.n581 B.n580 585
R177 B.n582 B.n27 585
R178 B.n584 B.n583 585
R179 B.n585 B.n26 585
R180 B.n587 B.n586 585
R181 B.n588 B.n25 585
R182 B.n590 B.n589 585
R183 B.n591 B.n24 585
R184 B.n593 B.n592 585
R185 B.n594 B.n23 585
R186 B.n596 B.n595 585
R187 B.n597 B.n22 585
R188 B.n599 B.n598 585
R189 B.n600 B.n21 585
R190 B.n602 B.n601 585
R191 B.n603 B.n20 585
R192 B.n605 B.n604 585
R193 B.n606 B.n19 585
R194 B.n608 B.n607 585
R195 B.n609 B.n18 585
R196 B.n611 B.n610 585
R197 B.n612 B.n17 585
R198 B.n614 B.n613 585
R199 B.n615 B.n16 585
R200 B.n617 B.n616 585
R201 B.n618 B.n15 585
R202 B.n620 B.n619 585
R203 B.n621 B.n14 585
R204 B.n623 B.n622 585
R205 B.n624 B.n13 585
R206 B.n626 B.n625 585
R207 B.n627 B.n12 585
R208 B.n629 B.n628 585
R209 B.n630 B.n11 585
R210 B.n632 B.n631 585
R211 B.n633 B.n10 585
R212 B.n635 B.n634 585
R213 B.n437 B.n436 585
R214 B.n435 B.n80 585
R215 B.n434 B.n433 585
R216 B.n432 B.n81 585
R217 B.n431 B.n430 585
R218 B.n429 B.n82 585
R219 B.n428 B.n427 585
R220 B.n426 B.n83 585
R221 B.n425 B.n424 585
R222 B.n423 B.n84 585
R223 B.n422 B.n421 585
R224 B.n420 B.n85 585
R225 B.n419 B.n418 585
R226 B.n417 B.n86 585
R227 B.n416 B.n415 585
R228 B.n414 B.n87 585
R229 B.n413 B.n412 585
R230 B.n411 B.n88 585
R231 B.n410 B.n409 585
R232 B.n408 B.n89 585
R233 B.n407 B.n406 585
R234 B.n405 B.n90 585
R235 B.n404 B.n403 585
R236 B.n402 B.n91 585
R237 B.n401 B.n400 585
R238 B.n399 B.n92 585
R239 B.n398 B.n397 585
R240 B.n396 B.n93 585
R241 B.n395 B.n394 585
R242 B.n393 B.n94 585
R243 B.n392 B.n391 585
R244 B.n194 B.n193 585
R245 B.n195 B.n164 585
R246 B.n197 B.n196 585
R247 B.n198 B.n163 585
R248 B.n200 B.n199 585
R249 B.n201 B.n162 585
R250 B.n203 B.n202 585
R251 B.n204 B.n161 585
R252 B.n206 B.n205 585
R253 B.n207 B.n160 585
R254 B.n209 B.n208 585
R255 B.n210 B.n159 585
R256 B.n212 B.n211 585
R257 B.n213 B.n158 585
R258 B.n215 B.n214 585
R259 B.n216 B.n157 585
R260 B.n218 B.n217 585
R261 B.n219 B.n156 585
R262 B.n221 B.n220 585
R263 B.n222 B.n155 585
R264 B.n224 B.n223 585
R265 B.n225 B.n154 585
R266 B.n227 B.n226 585
R267 B.n228 B.n153 585
R268 B.n230 B.n229 585
R269 B.n231 B.n152 585
R270 B.n233 B.n232 585
R271 B.n234 B.n151 585
R272 B.n236 B.n235 585
R273 B.n237 B.n150 585
R274 B.n239 B.n238 585
R275 B.n240 B.n149 585
R276 B.n242 B.n241 585
R277 B.n243 B.n148 585
R278 B.n245 B.n244 585
R279 B.n246 B.n147 585
R280 B.n248 B.n247 585
R281 B.n249 B.n146 585
R282 B.n251 B.n250 585
R283 B.n252 B.n145 585
R284 B.n254 B.n253 585
R285 B.n255 B.n144 585
R286 B.n257 B.n256 585
R287 B.n258 B.n143 585
R288 B.n260 B.n259 585
R289 B.n261 B.n142 585
R290 B.n263 B.n262 585
R291 B.n264 B.n141 585
R292 B.n266 B.n265 585
R293 B.n267 B.n140 585
R294 B.n269 B.n268 585
R295 B.n270 B.n139 585
R296 B.n272 B.n271 585
R297 B.n273 B.n138 585
R298 B.n275 B.n274 585
R299 B.n276 B.n137 585
R300 B.n278 B.n277 585
R301 B.n279 B.n136 585
R302 B.n281 B.n280 585
R303 B.n282 B.n135 585
R304 B.n284 B.n283 585
R305 B.n286 B.n285 585
R306 B.n287 B.n131 585
R307 B.n289 B.n288 585
R308 B.n290 B.n130 585
R309 B.n292 B.n291 585
R310 B.n293 B.n129 585
R311 B.n295 B.n294 585
R312 B.n296 B.n128 585
R313 B.n298 B.n297 585
R314 B.n300 B.n125 585
R315 B.n302 B.n301 585
R316 B.n303 B.n124 585
R317 B.n305 B.n304 585
R318 B.n306 B.n123 585
R319 B.n308 B.n307 585
R320 B.n309 B.n122 585
R321 B.n311 B.n310 585
R322 B.n312 B.n121 585
R323 B.n314 B.n313 585
R324 B.n315 B.n120 585
R325 B.n317 B.n316 585
R326 B.n318 B.n119 585
R327 B.n320 B.n319 585
R328 B.n321 B.n118 585
R329 B.n323 B.n322 585
R330 B.n324 B.n117 585
R331 B.n326 B.n325 585
R332 B.n327 B.n116 585
R333 B.n329 B.n328 585
R334 B.n330 B.n115 585
R335 B.n332 B.n331 585
R336 B.n333 B.n114 585
R337 B.n335 B.n334 585
R338 B.n336 B.n113 585
R339 B.n338 B.n337 585
R340 B.n339 B.n112 585
R341 B.n341 B.n340 585
R342 B.n342 B.n111 585
R343 B.n344 B.n343 585
R344 B.n345 B.n110 585
R345 B.n347 B.n346 585
R346 B.n348 B.n109 585
R347 B.n350 B.n349 585
R348 B.n351 B.n108 585
R349 B.n353 B.n352 585
R350 B.n354 B.n107 585
R351 B.n356 B.n355 585
R352 B.n357 B.n106 585
R353 B.n359 B.n358 585
R354 B.n360 B.n105 585
R355 B.n362 B.n361 585
R356 B.n363 B.n104 585
R357 B.n365 B.n364 585
R358 B.n366 B.n103 585
R359 B.n368 B.n367 585
R360 B.n369 B.n102 585
R361 B.n371 B.n370 585
R362 B.n372 B.n101 585
R363 B.n374 B.n373 585
R364 B.n375 B.n100 585
R365 B.n377 B.n376 585
R366 B.n378 B.n99 585
R367 B.n380 B.n379 585
R368 B.n381 B.n98 585
R369 B.n383 B.n382 585
R370 B.n384 B.n97 585
R371 B.n386 B.n385 585
R372 B.n387 B.n96 585
R373 B.n389 B.n388 585
R374 B.n390 B.n95 585
R375 B.n192 B.n165 585
R376 B.n191 B.n190 585
R377 B.n189 B.n166 585
R378 B.n188 B.n187 585
R379 B.n186 B.n167 585
R380 B.n185 B.n184 585
R381 B.n183 B.n168 585
R382 B.n182 B.n181 585
R383 B.n180 B.n169 585
R384 B.n179 B.n178 585
R385 B.n177 B.n170 585
R386 B.n176 B.n175 585
R387 B.n174 B.n171 585
R388 B.n173 B.n172 585
R389 B.n2 B.n0 585
R390 B.n657 B.n1 585
R391 B.n656 B.n655 585
R392 B.n654 B.n3 585
R393 B.n653 B.n652 585
R394 B.n651 B.n4 585
R395 B.n650 B.n649 585
R396 B.n648 B.n5 585
R397 B.n647 B.n646 585
R398 B.n645 B.n6 585
R399 B.n644 B.n643 585
R400 B.n642 B.n7 585
R401 B.n641 B.n640 585
R402 B.n639 B.n8 585
R403 B.n638 B.n637 585
R404 B.n636 B.n9 585
R405 B.n659 B.n658 585
R406 B.n194 B.n165 463.671
R407 B.n634 B.n9 463.671
R408 B.n392 B.n95 463.671
R409 B.n436 B.n79 463.671
R410 B.n190 B.n165 163.367
R411 B.n190 B.n189 163.367
R412 B.n189 B.n188 163.367
R413 B.n188 B.n167 163.367
R414 B.n184 B.n167 163.367
R415 B.n184 B.n183 163.367
R416 B.n183 B.n182 163.367
R417 B.n182 B.n169 163.367
R418 B.n178 B.n169 163.367
R419 B.n178 B.n177 163.367
R420 B.n177 B.n176 163.367
R421 B.n176 B.n171 163.367
R422 B.n172 B.n171 163.367
R423 B.n172 B.n2 163.367
R424 B.n658 B.n2 163.367
R425 B.n658 B.n657 163.367
R426 B.n657 B.n656 163.367
R427 B.n656 B.n3 163.367
R428 B.n652 B.n3 163.367
R429 B.n652 B.n651 163.367
R430 B.n651 B.n650 163.367
R431 B.n650 B.n5 163.367
R432 B.n646 B.n5 163.367
R433 B.n646 B.n645 163.367
R434 B.n645 B.n644 163.367
R435 B.n644 B.n7 163.367
R436 B.n640 B.n7 163.367
R437 B.n640 B.n639 163.367
R438 B.n639 B.n638 163.367
R439 B.n638 B.n9 163.367
R440 B.n195 B.n194 163.367
R441 B.n196 B.n195 163.367
R442 B.n196 B.n163 163.367
R443 B.n200 B.n163 163.367
R444 B.n201 B.n200 163.367
R445 B.n202 B.n201 163.367
R446 B.n202 B.n161 163.367
R447 B.n206 B.n161 163.367
R448 B.n207 B.n206 163.367
R449 B.n208 B.n207 163.367
R450 B.n208 B.n159 163.367
R451 B.n212 B.n159 163.367
R452 B.n213 B.n212 163.367
R453 B.n214 B.n213 163.367
R454 B.n214 B.n157 163.367
R455 B.n218 B.n157 163.367
R456 B.n219 B.n218 163.367
R457 B.n220 B.n219 163.367
R458 B.n220 B.n155 163.367
R459 B.n224 B.n155 163.367
R460 B.n225 B.n224 163.367
R461 B.n226 B.n225 163.367
R462 B.n226 B.n153 163.367
R463 B.n230 B.n153 163.367
R464 B.n231 B.n230 163.367
R465 B.n232 B.n231 163.367
R466 B.n232 B.n151 163.367
R467 B.n236 B.n151 163.367
R468 B.n237 B.n236 163.367
R469 B.n238 B.n237 163.367
R470 B.n238 B.n149 163.367
R471 B.n242 B.n149 163.367
R472 B.n243 B.n242 163.367
R473 B.n244 B.n243 163.367
R474 B.n244 B.n147 163.367
R475 B.n248 B.n147 163.367
R476 B.n249 B.n248 163.367
R477 B.n250 B.n249 163.367
R478 B.n250 B.n145 163.367
R479 B.n254 B.n145 163.367
R480 B.n255 B.n254 163.367
R481 B.n256 B.n255 163.367
R482 B.n256 B.n143 163.367
R483 B.n260 B.n143 163.367
R484 B.n261 B.n260 163.367
R485 B.n262 B.n261 163.367
R486 B.n262 B.n141 163.367
R487 B.n266 B.n141 163.367
R488 B.n267 B.n266 163.367
R489 B.n268 B.n267 163.367
R490 B.n268 B.n139 163.367
R491 B.n272 B.n139 163.367
R492 B.n273 B.n272 163.367
R493 B.n274 B.n273 163.367
R494 B.n274 B.n137 163.367
R495 B.n278 B.n137 163.367
R496 B.n279 B.n278 163.367
R497 B.n280 B.n279 163.367
R498 B.n280 B.n135 163.367
R499 B.n284 B.n135 163.367
R500 B.n285 B.n284 163.367
R501 B.n285 B.n131 163.367
R502 B.n289 B.n131 163.367
R503 B.n290 B.n289 163.367
R504 B.n291 B.n290 163.367
R505 B.n291 B.n129 163.367
R506 B.n295 B.n129 163.367
R507 B.n296 B.n295 163.367
R508 B.n297 B.n296 163.367
R509 B.n297 B.n125 163.367
R510 B.n302 B.n125 163.367
R511 B.n303 B.n302 163.367
R512 B.n304 B.n303 163.367
R513 B.n304 B.n123 163.367
R514 B.n308 B.n123 163.367
R515 B.n309 B.n308 163.367
R516 B.n310 B.n309 163.367
R517 B.n310 B.n121 163.367
R518 B.n314 B.n121 163.367
R519 B.n315 B.n314 163.367
R520 B.n316 B.n315 163.367
R521 B.n316 B.n119 163.367
R522 B.n320 B.n119 163.367
R523 B.n321 B.n320 163.367
R524 B.n322 B.n321 163.367
R525 B.n322 B.n117 163.367
R526 B.n326 B.n117 163.367
R527 B.n327 B.n326 163.367
R528 B.n328 B.n327 163.367
R529 B.n328 B.n115 163.367
R530 B.n332 B.n115 163.367
R531 B.n333 B.n332 163.367
R532 B.n334 B.n333 163.367
R533 B.n334 B.n113 163.367
R534 B.n338 B.n113 163.367
R535 B.n339 B.n338 163.367
R536 B.n340 B.n339 163.367
R537 B.n340 B.n111 163.367
R538 B.n344 B.n111 163.367
R539 B.n345 B.n344 163.367
R540 B.n346 B.n345 163.367
R541 B.n346 B.n109 163.367
R542 B.n350 B.n109 163.367
R543 B.n351 B.n350 163.367
R544 B.n352 B.n351 163.367
R545 B.n352 B.n107 163.367
R546 B.n356 B.n107 163.367
R547 B.n357 B.n356 163.367
R548 B.n358 B.n357 163.367
R549 B.n358 B.n105 163.367
R550 B.n362 B.n105 163.367
R551 B.n363 B.n362 163.367
R552 B.n364 B.n363 163.367
R553 B.n364 B.n103 163.367
R554 B.n368 B.n103 163.367
R555 B.n369 B.n368 163.367
R556 B.n370 B.n369 163.367
R557 B.n370 B.n101 163.367
R558 B.n374 B.n101 163.367
R559 B.n375 B.n374 163.367
R560 B.n376 B.n375 163.367
R561 B.n376 B.n99 163.367
R562 B.n380 B.n99 163.367
R563 B.n381 B.n380 163.367
R564 B.n382 B.n381 163.367
R565 B.n382 B.n97 163.367
R566 B.n386 B.n97 163.367
R567 B.n387 B.n386 163.367
R568 B.n388 B.n387 163.367
R569 B.n388 B.n95 163.367
R570 B.n393 B.n392 163.367
R571 B.n394 B.n393 163.367
R572 B.n394 B.n93 163.367
R573 B.n398 B.n93 163.367
R574 B.n399 B.n398 163.367
R575 B.n400 B.n399 163.367
R576 B.n400 B.n91 163.367
R577 B.n404 B.n91 163.367
R578 B.n405 B.n404 163.367
R579 B.n406 B.n405 163.367
R580 B.n406 B.n89 163.367
R581 B.n410 B.n89 163.367
R582 B.n411 B.n410 163.367
R583 B.n412 B.n411 163.367
R584 B.n412 B.n87 163.367
R585 B.n416 B.n87 163.367
R586 B.n417 B.n416 163.367
R587 B.n418 B.n417 163.367
R588 B.n418 B.n85 163.367
R589 B.n422 B.n85 163.367
R590 B.n423 B.n422 163.367
R591 B.n424 B.n423 163.367
R592 B.n424 B.n83 163.367
R593 B.n428 B.n83 163.367
R594 B.n429 B.n428 163.367
R595 B.n430 B.n429 163.367
R596 B.n430 B.n81 163.367
R597 B.n434 B.n81 163.367
R598 B.n435 B.n434 163.367
R599 B.n436 B.n435 163.367
R600 B.n634 B.n633 163.367
R601 B.n633 B.n632 163.367
R602 B.n632 B.n11 163.367
R603 B.n628 B.n11 163.367
R604 B.n628 B.n627 163.367
R605 B.n627 B.n626 163.367
R606 B.n626 B.n13 163.367
R607 B.n622 B.n13 163.367
R608 B.n622 B.n621 163.367
R609 B.n621 B.n620 163.367
R610 B.n620 B.n15 163.367
R611 B.n616 B.n15 163.367
R612 B.n616 B.n615 163.367
R613 B.n615 B.n614 163.367
R614 B.n614 B.n17 163.367
R615 B.n610 B.n17 163.367
R616 B.n610 B.n609 163.367
R617 B.n609 B.n608 163.367
R618 B.n608 B.n19 163.367
R619 B.n604 B.n19 163.367
R620 B.n604 B.n603 163.367
R621 B.n603 B.n602 163.367
R622 B.n602 B.n21 163.367
R623 B.n598 B.n21 163.367
R624 B.n598 B.n597 163.367
R625 B.n597 B.n596 163.367
R626 B.n596 B.n23 163.367
R627 B.n592 B.n23 163.367
R628 B.n592 B.n591 163.367
R629 B.n591 B.n590 163.367
R630 B.n590 B.n25 163.367
R631 B.n586 B.n25 163.367
R632 B.n586 B.n585 163.367
R633 B.n585 B.n584 163.367
R634 B.n584 B.n27 163.367
R635 B.n580 B.n27 163.367
R636 B.n580 B.n579 163.367
R637 B.n579 B.n578 163.367
R638 B.n578 B.n29 163.367
R639 B.n574 B.n29 163.367
R640 B.n574 B.n573 163.367
R641 B.n573 B.n572 163.367
R642 B.n572 B.n31 163.367
R643 B.n568 B.n31 163.367
R644 B.n568 B.n567 163.367
R645 B.n567 B.n566 163.367
R646 B.n566 B.n33 163.367
R647 B.n562 B.n33 163.367
R648 B.n562 B.n561 163.367
R649 B.n561 B.n560 163.367
R650 B.n560 B.n35 163.367
R651 B.n556 B.n35 163.367
R652 B.n556 B.n555 163.367
R653 B.n555 B.n554 163.367
R654 B.n554 B.n37 163.367
R655 B.n550 B.n37 163.367
R656 B.n550 B.n549 163.367
R657 B.n549 B.n548 163.367
R658 B.n548 B.n39 163.367
R659 B.n544 B.n39 163.367
R660 B.n544 B.n543 163.367
R661 B.n543 B.n43 163.367
R662 B.n539 B.n43 163.367
R663 B.n539 B.n538 163.367
R664 B.n538 B.n537 163.367
R665 B.n537 B.n45 163.367
R666 B.n533 B.n45 163.367
R667 B.n533 B.n532 163.367
R668 B.n532 B.n531 163.367
R669 B.n531 B.n47 163.367
R670 B.n526 B.n47 163.367
R671 B.n526 B.n525 163.367
R672 B.n525 B.n524 163.367
R673 B.n524 B.n51 163.367
R674 B.n520 B.n51 163.367
R675 B.n520 B.n519 163.367
R676 B.n519 B.n518 163.367
R677 B.n518 B.n53 163.367
R678 B.n514 B.n53 163.367
R679 B.n514 B.n513 163.367
R680 B.n513 B.n512 163.367
R681 B.n512 B.n55 163.367
R682 B.n508 B.n55 163.367
R683 B.n508 B.n507 163.367
R684 B.n507 B.n506 163.367
R685 B.n506 B.n57 163.367
R686 B.n502 B.n57 163.367
R687 B.n502 B.n501 163.367
R688 B.n501 B.n500 163.367
R689 B.n500 B.n59 163.367
R690 B.n496 B.n59 163.367
R691 B.n496 B.n495 163.367
R692 B.n495 B.n494 163.367
R693 B.n494 B.n61 163.367
R694 B.n490 B.n61 163.367
R695 B.n490 B.n489 163.367
R696 B.n489 B.n488 163.367
R697 B.n488 B.n63 163.367
R698 B.n484 B.n63 163.367
R699 B.n484 B.n483 163.367
R700 B.n483 B.n482 163.367
R701 B.n482 B.n65 163.367
R702 B.n478 B.n65 163.367
R703 B.n478 B.n477 163.367
R704 B.n477 B.n476 163.367
R705 B.n476 B.n67 163.367
R706 B.n472 B.n67 163.367
R707 B.n472 B.n471 163.367
R708 B.n471 B.n470 163.367
R709 B.n470 B.n69 163.367
R710 B.n466 B.n69 163.367
R711 B.n466 B.n465 163.367
R712 B.n465 B.n464 163.367
R713 B.n464 B.n71 163.367
R714 B.n460 B.n71 163.367
R715 B.n460 B.n459 163.367
R716 B.n459 B.n458 163.367
R717 B.n458 B.n73 163.367
R718 B.n454 B.n73 163.367
R719 B.n454 B.n453 163.367
R720 B.n453 B.n452 163.367
R721 B.n452 B.n75 163.367
R722 B.n448 B.n75 163.367
R723 B.n448 B.n447 163.367
R724 B.n447 B.n446 163.367
R725 B.n446 B.n77 163.367
R726 B.n442 B.n77 163.367
R727 B.n442 B.n441 163.367
R728 B.n441 B.n440 163.367
R729 B.n440 B.n79 163.367
R730 B.n126 B.t5 119.54
R731 B.n48 B.t7 119.54
R732 B.n132 B.t11 119.516
R733 B.n40 B.t1 119.516
R734 B.n127 B.t4 108.486
R735 B.n49 B.t8 108.486
R736 B.n133 B.t10 108.462
R737 B.n41 B.t2 108.462
R738 B.n299 B.n127 59.5399
R739 B.n134 B.n133 59.5399
R740 B.n42 B.n41 59.5399
R741 B.n529 B.n49 59.5399
R742 B.n636 B.n635 30.1273
R743 B.n391 B.n390 30.1273
R744 B.n193 B.n192 30.1273
R745 B.n438 B.n437 30.1273
R746 B B.n659 18.0485
R747 B.n127 B.n126 11.055
R748 B.n133 B.n132 11.055
R749 B.n41 B.n40 11.055
R750 B.n49 B.n48 11.055
R751 B.n635 B.n10 10.6151
R752 B.n631 B.n10 10.6151
R753 B.n631 B.n630 10.6151
R754 B.n630 B.n629 10.6151
R755 B.n629 B.n12 10.6151
R756 B.n625 B.n12 10.6151
R757 B.n625 B.n624 10.6151
R758 B.n624 B.n623 10.6151
R759 B.n623 B.n14 10.6151
R760 B.n619 B.n14 10.6151
R761 B.n619 B.n618 10.6151
R762 B.n618 B.n617 10.6151
R763 B.n617 B.n16 10.6151
R764 B.n613 B.n16 10.6151
R765 B.n613 B.n612 10.6151
R766 B.n612 B.n611 10.6151
R767 B.n611 B.n18 10.6151
R768 B.n607 B.n18 10.6151
R769 B.n607 B.n606 10.6151
R770 B.n606 B.n605 10.6151
R771 B.n605 B.n20 10.6151
R772 B.n601 B.n20 10.6151
R773 B.n601 B.n600 10.6151
R774 B.n600 B.n599 10.6151
R775 B.n599 B.n22 10.6151
R776 B.n595 B.n22 10.6151
R777 B.n595 B.n594 10.6151
R778 B.n594 B.n593 10.6151
R779 B.n593 B.n24 10.6151
R780 B.n589 B.n24 10.6151
R781 B.n589 B.n588 10.6151
R782 B.n588 B.n587 10.6151
R783 B.n587 B.n26 10.6151
R784 B.n583 B.n26 10.6151
R785 B.n583 B.n582 10.6151
R786 B.n582 B.n581 10.6151
R787 B.n581 B.n28 10.6151
R788 B.n577 B.n28 10.6151
R789 B.n577 B.n576 10.6151
R790 B.n576 B.n575 10.6151
R791 B.n575 B.n30 10.6151
R792 B.n571 B.n30 10.6151
R793 B.n571 B.n570 10.6151
R794 B.n570 B.n569 10.6151
R795 B.n569 B.n32 10.6151
R796 B.n565 B.n32 10.6151
R797 B.n565 B.n564 10.6151
R798 B.n564 B.n563 10.6151
R799 B.n563 B.n34 10.6151
R800 B.n559 B.n34 10.6151
R801 B.n559 B.n558 10.6151
R802 B.n558 B.n557 10.6151
R803 B.n557 B.n36 10.6151
R804 B.n553 B.n36 10.6151
R805 B.n553 B.n552 10.6151
R806 B.n552 B.n551 10.6151
R807 B.n551 B.n38 10.6151
R808 B.n547 B.n38 10.6151
R809 B.n547 B.n546 10.6151
R810 B.n546 B.n545 10.6151
R811 B.n542 B.n541 10.6151
R812 B.n541 B.n540 10.6151
R813 B.n540 B.n44 10.6151
R814 B.n536 B.n44 10.6151
R815 B.n536 B.n535 10.6151
R816 B.n535 B.n534 10.6151
R817 B.n534 B.n46 10.6151
R818 B.n530 B.n46 10.6151
R819 B.n528 B.n527 10.6151
R820 B.n527 B.n50 10.6151
R821 B.n523 B.n50 10.6151
R822 B.n523 B.n522 10.6151
R823 B.n522 B.n521 10.6151
R824 B.n521 B.n52 10.6151
R825 B.n517 B.n52 10.6151
R826 B.n517 B.n516 10.6151
R827 B.n516 B.n515 10.6151
R828 B.n515 B.n54 10.6151
R829 B.n511 B.n54 10.6151
R830 B.n511 B.n510 10.6151
R831 B.n510 B.n509 10.6151
R832 B.n509 B.n56 10.6151
R833 B.n505 B.n56 10.6151
R834 B.n505 B.n504 10.6151
R835 B.n504 B.n503 10.6151
R836 B.n503 B.n58 10.6151
R837 B.n499 B.n58 10.6151
R838 B.n499 B.n498 10.6151
R839 B.n498 B.n497 10.6151
R840 B.n497 B.n60 10.6151
R841 B.n493 B.n60 10.6151
R842 B.n493 B.n492 10.6151
R843 B.n492 B.n491 10.6151
R844 B.n491 B.n62 10.6151
R845 B.n487 B.n62 10.6151
R846 B.n487 B.n486 10.6151
R847 B.n486 B.n485 10.6151
R848 B.n485 B.n64 10.6151
R849 B.n481 B.n64 10.6151
R850 B.n481 B.n480 10.6151
R851 B.n480 B.n479 10.6151
R852 B.n479 B.n66 10.6151
R853 B.n475 B.n66 10.6151
R854 B.n475 B.n474 10.6151
R855 B.n474 B.n473 10.6151
R856 B.n473 B.n68 10.6151
R857 B.n469 B.n68 10.6151
R858 B.n469 B.n468 10.6151
R859 B.n468 B.n467 10.6151
R860 B.n467 B.n70 10.6151
R861 B.n463 B.n70 10.6151
R862 B.n463 B.n462 10.6151
R863 B.n462 B.n461 10.6151
R864 B.n461 B.n72 10.6151
R865 B.n457 B.n72 10.6151
R866 B.n457 B.n456 10.6151
R867 B.n456 B.n455 10.6151
R868 B.n455 B.n74 10.6151
R869 B.n451 B.n74 10.6151
R870 B.n451 B.n450 10.6151
R871 B.n450 B.n449 10.6151
R872 B.n449 B.n76 10.6151
R873 B.n445 B.n76 10.6151
R874 B.n445 B.n444 10.6151
R875 B.n444 B.n443 10.6151
R876 B.n443 B.n78 10.6151
R877 B.n439 B.n78 10.6151
R878 B.n439 B.n438 10.6151
R879 B.n391 B.n94 10.6151
R880 B.n395 B.n94 10.6151
R881 B.n396 B.n395 10.6151
R882 B.n397 B.n396 10.6151
R883 B.n397 B.n92 10.6151
R884 B.n401 B.n92 10.6151
R885 B.n402 B.n401 10.6151
R886 B.n403 B.n402 10.6151
R887 B.n403 B.n90 10.6151
R888 B.n407 B.n90 10.6151
R889 B.n408 B.n407 10.6151
R890 B.n409 B.n408 10.6151
R891 B.n409 B.n88 10.6151
R892 B.n413 B.n88 10.6151
R893 B.n414 B.n413 10.6151
R894 B.n415 B.n414 10.6151
R895 B.n415 B.n86 10.6151
R896 B.n419 B.n86 10.6151
R897 B.n420 B.n419 10.6151
R898 B.n421 B.n420 10.6151
R899 B.n421 B.n84 10.6151
R900 B.n425 B.n84 10.6151
R901 B.n426 B.n425 10.6151
R902 B.n427 B.n426 10.6151
R903 B.n427 B.n82 10.6151
R904 B.n431 B.n82 10.6151
R905 B.n432 B.n431 10.6151
R906 B.n433 B.n432 10.6151
R907 B.n433 B.n80 10.6151
R908 B.n437 B.n80 10.6151
R909 B.n193 B.n164 10.6151
R910 B.n197 B.n164 10.6151
R911 B.n198 B.n197 10.6151
R912 B.n199 B.n198 10.6151
R913 B.n199 B.n162 10.6151
R914 B.n203 B.n162 10.6151
R915 B.n204 B.n203 10.6151
R916 B.n205 B.n204 10.6151
R917 B.n205 B.n160 10.6151
R918 B.n209 B.n160 10.6151
R919 B.n210 B.n209 10.6151
R920 B.n211 B.n210 10.6151
R921 B.n211 B.n158 10.6151
R922 B.n215 B.n158 10.6151
R923 B.n216 B.n215 10.6151
R924 B.n217 B.n216 10.6151
R925 B.n217 B.n156 10.6151
R926 B.n221 B.n156 10.6151
R927 B.n222 B.n221 10.6151
R928 B.n223 B.n222 10.6151
R929 B.n223 B.n154 10.6151
R930 B.n227 B.n154 10.6151
R931 B.n228 B.n227 10.6151
R932 B.n229 B.n228 10.6151
R933 B.n229 B.n152 10.6151
R934 B.n233 B.n152 10.6151
R935 B.n234 B.n233 10.6151
R936 B.n235 B.n234 10.6151
R937 B.n235 B.n150 10.6151
R938 B.n239 B.n150 10.6151
R939 B.n240 B.n239 10.6151
R940 B.n241 B.n240 10.6151
R941 B.n241 B.n148 10.6151
R942 B.n245 B.n148 10.6151
R943 B.n246 B.n245 10.6151
R944 B.n247 B.n246 10.6151
R945 B.n247 B.n146 10.6151
R946 B.n251 B.n146 10.6151
R947 B.n252 B.n251 10.6151
R948 B.n253 B.n252 10.6151
R949 B.n253 B.n144 10.6151
R950 B.n257 B.n144 10.6151
R951 B.n258 B.n257 10.6151
R952 B.n259 B.n258 10.6151
R953 B.n259 B.n142 10.6151
R954 B.n263 B.n142 10.6151
R955 B.n264 B.n263 10.6151
R956 B.n265 B.n264 10.6151
R957 B.n265 B.n140 10.6151
R958 B.n269 B.n140 10.6151
R959 B.n270 B.n269 10.6151
R960 B.n271 B.n270 10.6151
R961 B.n271 B.n138 10.6151
R962 B.n275 B.n138 10.6151
R963 B.n276 B.n275 10.6151
R964 B.n277 B.n276 10.6151
R965 B.n277 B.n136 10.6151
R966 B.n281 B.n136 10.6151
R967 B.n282 B.n281 10.6151
R968 B.n283 B.n282 10.6151
R969 B.n287 B.n286 10.6151
R970 B.n288 B.n287 10.6151
R971 B.n288 B.n130 10.6151
R972 B.n292 B.n130 10.6151
R973 B.n293 B.n292 10.6151
R974 B.n294 B.n293 10.6151
R975 B.n294 B.n128 10.6151
R976 B.n298 B.n128 10.6151
R977 B.n301 B.n300 10.6151
R978 B.n301 B.n124 10.6151
R979 B.n305 B.n124 10.6151
R980 B.n306 B.n305 10.6151
R981 B.n307 B.n306 10.6151
R982 B.n307 B.n122 10.6151
R983 B.n311 B.n122 10.6151
R984 B.n312 B.n311 10.6151
R985 B.n313 B.n312 10.6151
R986 B.n313 B.n120 10.6151
R987 B.n317 B.n120 10.6151
R988 B.n318 B.n317 10.6151
R989 B.n319 B.n318 10.6151
R990 B.n319 B.n118 10.6151
R991 B.n323 B.n118 10.6151
R992 B.n324 B.n323 10.6151
R993 B.n325 B.n324 10.6151
R994 B.n325 B.n116 10.6151
R995 B.n329 B.n116 10.6151
R996 B.n330 B.n329 10.6151
R997 B.n331 B.n330 10.6151
R998 B.n331 B.n114 10.6151
R999 B.n335 B.n114 10.6151
R1000 B.n336 B.n335 10.6151
R1001 B.n337 B.n336 10.6151
R1002 B.n337 B.n112 10.6151
R1003 B.n341 B.n112 10.6151
R1004 B.n342 B.n341 10.6151
R1005 B.n343 B.n342 10.6151
R1006 B.n343 B.n110 10.6151
R1007 B.n347 B.n110 10.6151
R1008 B.n348 B.n347 10.6151
R1009 B.n349 B.n348 10.6151
R1010 B.n349 B.n108 10.6151
R1011 B.n353 B.n108 10.6151
R1012 B.n354 B.n353 10.6151
R1013 B.n355 B.n354 10.6151
R1014 B.n355 B.n106 10.6151
R1015 B.n359 B.n106 10.6151
R1016 B.n360 B.n359 10.6151
R1017 B.n361 B.n360 10.6151
R1018 B.n361 B.n104 10.6151
R1019 B.n365 B.n104 10.6151
R1020 B.n366 B.n365 10.6151
R1021 B.n367 B.n366 10.6151
R1022 B.n367 B.n102 10.6151
R1023 B.n371 B.n102 10.6151
R1024 B.n372 B.n371 10.6151
R1025 B.n373 B.n372 10.6151
R1026 B.n373 B.n100 10.6151
R1027 B.n377 B.n100 10.6151
R1028 B.n378 B.n377 10.6151
R1029 B.n379 B.n378 10.6151
R1030 B.n379 B.n98 10.6151
R1031 B.n383 B.n98 10.6151
R1032 B.n384 B.n383 10.6151
R1033 B.n385 B.n384 10.6151
R1034 B.n385 B.n96 10.6151
R1035 B.n389 B.n96 10.6151
R1036 B.n390 B.n389 10.6151
R1037 B.n192 B.n191 10.6151
R1038 B.n191 B.n166 10.6151
R1039 B.n187 B.n166 10.6151
R1040 B.n187 B.n186 10.6151
R1041 B.n186 B.n185 10.6151
R1042 B.n185 B.n168 10.6151
R1043 B.n181 B.n168 10.6151
R1044 B.n181 B.n180 10.6151
R1045 B.n180 B.n179 10.6151
R1046 B.n179 B.n170 10.6151
R1047 B.n175 B.n170 10.6151
R1048 B.n175 B.n174 10.6151
R1049 B.n174 B.n173 10.6151
R1050 B.n173 B.n0 10.6151
R1051 B.n655 B.n1 10.6151
R1052 B.n655 B.n654 10.6151
R1053 B.n654 B.n653 10.6151
R1054 B.n653 B.n4 10.6151
R1055 B.n649 B.n4 10.6151
R1056 B.n649 B.n648 10.6151
R1057 B.n648 B.n647 10.6151
R1058 B.n647 B.n6 10.6151
R1059 B.n643 B.n6 10.6151
R1060 B.n643 B.n642 10.6151
R1061 B.n642 B.n641 10.6151
R1062 B.n641 B.n8 10.6151
R1063 B.n637 B.n8 10.6151
R1064 B.n637 B.n636 10.6151
R1065 B.n542 B.n42 6.5566
R1066 B.n530 B.n529 6.5566
R1067 B.n286 B.n134 6.5566
R1068 B.n299 B.n298 6.5566
R1069 B.n545 B.n42 4.05904
R1070 B.n529 B.n528 4.05904
R1071 B.n283 B.n134 4.05904
R1072 B.n300 B.n299 4.05904
R1073 B.n659 B.n0 2.81026
R1074 B.n659 B.n1 2.81026
C0 VDD2 VP 0.260243f
C1 VDD2 VN 3.5154f
C2 B VTAIL 3.43298f
C3 B VDD1 1.86435f
C4 VTAIL VDD1 22.5502f
C5 B VP 1.02645f
C6 VN B 0.741506f
C7 VTAIL VP 2.74477f
C8 VN VTAIL 2.72961f
C9 VDD1 VP 3.62001f
C10 VN VDD1 0.14766f
C11 VDD2 w_n1426_n4664# 2.17524f
C12 VN VP 5.83051f
C13 w_n1426_n4664# B 8.27645f
C14 w_n1426_n4664# VTAIL 4.11691f
C15 w_n1426_n4664# VDD1 2.16475f
C16 VDD2 B 1.8833f
C17 VDD2 VTAIL 22.5742f
C18 VDD2 VDD1 0.551537f
C19 w_n1426_n4664# VP 2.42823f
C20 w_n1426_n4664# VN 2.25045f
C21 VDD2 VSUBS 1.689416f
C22 VDD1 VSUBS 1.969345f
C23 VTAIL VSUBS 0.701877f
C24 VN VSUBS 5.18136f
C25 VP VSUBS 1.367279f
C26 B VSUBS 2.839097f
C27 w_n1426_n4664# VSUBS 81.2991f
C28 B.n0 VSUBS 0.004655f
C29 B.n1 VSUBS 0.004655f
C30 B.n2 VSUBS 0.007361f
C31 B.n3 VSUBS 0.007361f
C32 B.n4 VSUBS 0.007361f
C33 B.n5 VSUBS 0.007361f
C34 B.n6 VSUBS 0.007361f
C35 B.n7 VSUBS 0.007361f
C36 B.n8 VSUBS 0.007361f
C37 B.n9 VSUBS 0.016012f
C38 B.n10 VSUBS 0.007361f
C39 B.n11 VSUBS 0.007361f
C40 B.n12 VSUBS 0.007361f
C41 B.n13 VSUBS 0.007361f
C42 B.n14 VSUBS 0.007361f
C43 B.n15 VSUBS 0.007361f
C44 B.n16 VSUBS 0.007361f
C45 B.n17 VSUBS 0.007361f
C46 B.n18 VSUBS 0.007361f
C47 B.n19 VSUBS 0.007361f
C48 B.n20 VSUBS 0.007361f
C49 B.n21 VSUBS 0.007361f
C50 B.n22 VSUBS 0.007361f
C51 B.n23 VSUBS 0.007361f
C52 B.n24 VSUBS 0.007361f
C53 B.n25 VSUBS 0.007361f
C54 B.n26 VSUBS 0.007361f
C55 B.n27 VSUBS 0.007361f
C56 B.n28 VSUBS 0.007361f
C57 B.n29 VSUBS 0.007361f
C58 B.n30 VSUBS 0.007361f
C59 B.n31 VSUBS 0.007361f
C60 B.n32 VSUBS 0.007361f
C61 B.n33 VSUBS 0.007361f
C62 B.n34 VSUBS 0.007361f
C63 B.n35 VSUBS 0.007361f
C64 B.n36 VSUBS 0.007361f
C65 B.n37 VSUBS 0.007361f
C66 B.n38 VSUBS 0.007361f
C67 B.n39 VSUBS 0.007361f
C68 B.t2 VSUBS 0.657207f
C69 B.t1 VSUBS 0.662301f
C70 B.t0 VSUBS 0.17958f
C71 B.n40 VSUBS 0.115305f
C72 B.n41 VSUBS 0.065572f
C73 B.n42 VSUBS 0.017054f
C74 B.n43 VSUBS 0.007361f
C75 B.n44 VSUBS 0.007361f
C76 B.n45 VSUBS 0.007361f
C77 B.n46 VSUBS 0.007361f
C78 B.n47 VSUBS 0.007361f
C79 B.t8 VSUBS 0.657181f
C80 B.t7 VSUBS 0.662277f
C81 B.t6 VSUBS 0.17958f
C82 B.n48 VSUBS 0.115329f
C83 B.n49 VSUBS 0.065598f
C84 B.n50 VSUBS 0.007361f
C85 B.n51 VSUBS 0.007361f
C86 B.n52 VSUBS 0.007361f
C87 B.n53 VSUBS 0.007361f
C88 B.n54 VSUBS 0.007361f
C89 B.n55 VSUBS 0.007361f
C90 B.n56 VSUBS 0.007361f
C91 B.n57 VSUBS 0.007361f
C92 B.n58 VSUBS 0.007361f
C93 B.n59 VSUBS 0.007361f
C94 B.n60 VSUBS 0.007361f
C95 B.n61 VSUBS 0.007361f
C96 B.n62 VSUBS 0.007361f
C97 B.n63 VSUBS 0.007361f
C98 B.n64 VSUBS 0.007361f
C99 B.n65 VSUBS 0.007361f
C100 B.n66 VSUBS 0.007361f
C101 B.n67 VSUBS 0.007361f
C102 B.n68 VSUBS 0.007361f
C103 B.n69 VSUBS 0.007361f
C104 B.n70 VSUBS 0.007361f
C105 B.n71 VSUBS 0.007361f
C106 B.n72 VSUBS 0.007361f
C107 B.n73 VSUBS 0.007361f
C108 B.n74 VSUBS 0.007361f
C109 B.n75 VSUBS 0.007361f
C110 B.n76 VSUBS 0.007361f
C111 B.n77 VSUBS 0.007361f
C112 B.n78 VSUBS 0.007361f
C113 B.n79 VSUBS 0.016678f
C114 B.n80 VSUBS 0.007361f
C115 B.n81 VSUBS 0.007361f
C116 B.n82 VSUBS 0.007361f
C117 B.n83 VSUBS 0.007361f
C118 B.n84 VSUBS 0.007361f
C119 B.n85 VSUBS 0.007361f
C120 B.n86 VSUBS 0.007361f
C121 B.n87 VSUBS 0.007361f
C122 B.n88 VSUBS 0.007361f
C123 B.n89 VSUBS 0.007361f
C124 B.n90 VSUBS 0.007361f
C125 B.n91 VSUBS 0.007361f
C126 B.n92 VSUBS 0.007361f
C127 B.n93 VSUBS 0.007361f
C128 B.n94 VSUBS 0.007361f
C129 B.n95 VSUBS 0.016678f
C130 B.n96 VSUBS 0.007361f
C131 B.n97 VSUBS 0.007361f
C132 B.n98 VSUBS 0.007361f
C133 B.n99 VSUBS 0.007361f
C134 B.n100 VSUBS 0.007361f
C135 B.n101 VSUBS 0.007361f
C136 B.n102 VSUBS 0.007361f
C137 B.n103 VSUBS 0.007361f
C138 B.n104 VSUBS 0.007361f
C139 B.n105 VSUBS 0.007361f
C140 B.n106 VSUBS 0.007361f
C141 B.n107 VSUBS 0.007361f
C142 B.n108 VSUBS 0.007361f
C143 B.n109 VSUBS 0.007361f
C144 B.n110 VSUBS 0.007361f
C145 B.n111 VSUBS 0.007361f
C146 B.n112 VSUBS 0.007361f
C147 B.n113 VSUBS 0.007361f
C148 B.n114 VSUBS 0.007361f
C149 B.n115 VSUBS 0.007361f
C150 B.n116 VSUBS 0.007361f
C151 B.n117 VSUBS 0.007361f
C152 B.n118 VSUBS 0.007361f
C153 B.n119 VSUBS 0.007361f
C154 B.n120 VSUBS 0.007361f
C155 B.n121 VSUBS 0.007361f
C156 B.n122 VSUBS 0.007361f
C157 B.n123 VSUBS 0.007361f
C158 B.n124 VSUBS 0.007361f
C159 B.n125 VSUBS 0.007361f
C160 B.t4 VSUBS 0.657181f
C161 B.t5 VSUBS 0.662277f
C162 B.t3 VSUBS 0.17958f
C163 B.n126 VSUBS 0.115329f
C164 B.n127 VSUBS 0.065598f
C165 B.n128 VSUBS 0.007361f
C166 B.n129 VSUBS 0.007361f
C167 B.n130 VSUBS 0.007361f
C168 B.n131 VSUBS 0.007361f
C169 B.t10 VSUBS 0.657207f
C170 B.t11 VSUBS 0.662301f
C171 B.t9 VSUBS 0.17958f
C172 B.n132 VSUBS 0.115305f
C173 B.n133 VSUBS 0.065572f
C174 B.n134 VSUBS 0.017054f
C175 B.n135 VSUBS 0.007361f
C176 B.n136 VSUBS 0.007361f
C177 B.n137 VSUBS 0.007361f
C178 B.n138 VSUBS 0.007361f
C179 B.n139 VSUBS 0.007361f
C180 B.n140 VSUBS 0.007361f
C181 B.n141 VSUBS 0.007361f
C182 B.n142 VSUBS 0.007361f
C183 B.n143 VSUBS 0.007361f
C184 B.n144 VSUBS 0.007361f
C185 B.n145 VSUBS 0.007361f
C186 B.n146 VSUBS 0.007361f
C187 B.n147 VSUBS 0.007361f
C188 B.n148 VSUBS 0.007361f
C189 B.n149 VSUBS 0.007361f
C190 B.n150 VSUBS 0.007361f
C191 B.n151 VSUBS 0.007361f
C192 B.n152 VSUBS 0.007361f
C193 B.n153 VSUBS 0.007361f
C194 B.n154 VSUBS 0.007361f
C195 B.n155 VSUBS 0.007361f
C196 B.n156 VSUBS 0.007361f
C197 B.n157 VSUBS 0.007361f
C198 B.n158 VSUBS 0.007361f
C199 B.n159 VSUBS 0.007361f
C200 B.n160 VSUBS 0.007361f
C201 B.n161 VSUBS 0.007361f
C202 B.n162 VSUBS 0.007361f
C203 B.n163 VSUBS 0.007361f
C204 B.n164 VSUBS 0.007361f
C205 B.n165 VSUBS 0.016012f
C206 B.n166 VSUBS 0.007361f
C207 B.n167 VSUBS 0.007361f
C208 B.n168 VSUBS 0.007361f
C209 B.n169 VSUBS 0.007361f
C210 B.n170 VSUBS 0.007361f
C211 B.n171 VSUBS 0.007361f
C212 B.n172 VSUBS 0.007361f
C213 B.n173 VSUBS 0.007361f
C214 B.n174 VSUBS 0.007361f
C215 B.n175 VSUBS 0.007361f
C216 B.n176 VSUBS 0.007361f
C217 B.n177 VSUBS 0.007361f
C218 B.n178 VSUBS 0.007361f
C219 B.n179 VSUBS 0.007361f
C220 B.n180 VSUBS 0.007361f
C221 B.n181 VSUBS 0.007361f
C222 B.n182 VSUBS 0.007361f
C223 B.n183 VSUBS 0.007361f
C224 B.n184 VSUBS 0.007361f
C225 B.n185 VSUBS 0.007361f
C226 B.n186 VSUBS 0.007361f
C227 B.n187 VSUBS 0.007361f
C228 B.n188 VSUBS 0.007361f
C229 B.n189 VSUBS 0.007361f
C230 B.n190 VSUBS 0.007361f
C231 B.n191 VSUBS 0.007361f
C232 B.n192 VSUBS 0.016012f
C233 B.n193 VSUBS 0.016678f
C234 B.n194 VSUBS 0.016678f
C235 B.n195 VSUBS 0.007361f
C236 B.n196 VSUBS 0.007361f
C237 B.n197 VSUBS 0.007361f
C238 B.n198 VSUBS 0.007361f
C239 B.n199 VSUBS 0.007361f
C240 B.n200 VSUBS 0.007361f
C241 B.n201 VSUBS 0.007361f
C242 B.n202 VSUBS 0.007361f
C243 B.n203 VSUBS 0.007361f
C244 B.n204 VSUBS 0.007361f
C245 B.n205 VSUBS 0.007361f
C246 B.n206 VSUBS 0.007361f
C247 B.n207 VSUBS 0.007361f
C248 B.n208 VSUBS 0.007361f
C249 B.n209 VSUBS 0.007361f
C250 B.n210 VSUBS 0.007361f
C251 B.n211 VSUBS 0.007361f
C252 B.n212 VSUBS 0.007361f
C253 B.n213 VSUBS 0.007361f
C254 B.n214 VSUBS 0.007361f
C255 B.n215 VSUBS 0.007361f
C256 B.n216 VSUBS 0.007361f
C257 B.n217 VSUBS 0.007361f
C258 B.n218 VSUBS 0.007361f
C259 B.n219 VSUBS 0.007361f
C260 B.n220 VSUBS 0.007361f
C261 B.n221 VSUBS 0.007361f
C262 B.n222 VSUBS 0.007361f
C263 B.n223 VSUBS 0.007361f
C264 B.n224 VSUBS 0.007361f
C265 B.n225 VSUBS 0.007361f
C266 B.n226 VSUBS 0.007361f
C267 B.n227 VSUBS 0.007361f
C268 B.n228 VSUBS 0.007361f
C269 B.n229 VSUBS 0.007361f
C270 B.n230 VSUBS 0.007361f
C271 B.n231 VSUBS 0.007361f
C272 B.n232 VSUBS 0.007361f
C273 B.n233 VSUBS 0.007361f
C274 B.n234 VSUBS 0.007361f
C275 B.n235 VSUBS 0.007361f
C276 B.n236 VSUBS 0.007361f
C277 B.n237 VSUBS 0.007361f
C278 B.n238 VSUBS 0.007361f
C279 B.n239 VSUBS 0.007361f
C280 B.n240 VSUBS 0.007361f
C281 B.n241 VSUBS 0.007361f
C282 B.n242 VSUBS 0.007361f
C283 B.n243 VSUBS 0.007361f
C284 B.n244 VSUBS 0.007361f
C285 B.n245 VSUBS 0.007361f
C286 B.n246 VSUBS 0.007361f
C287 B.n247 VSUBS 0.007361f
C288 B.n248 VSUBS 0.007361f
C289 B.n249 VSUBS 0.007361f
C290 B.n250 VSUBS 0.007361f
C291 B.n251 VSUBS 0.007361f
C292 B.n252 VSUBS 0.007361f
C293 B.n253 VSUBS 0.007361f
C294 B.n254 VSUBS 0.007361f
C295 B.n255 VSUBS 0.007361f
C296 B.n256 VSUBS 0.007361f
C297 B.n257 VSUBS 0.007361f
C298 B.n258 VSUBS 0.007361f
C299 B.n259 VSUBS 0.007361f
C300 B.n260 VSUBS 0.007361f
C301 B.n261 VSUBS 0.007361f
C302 B.n262 VSUBS 0.007361f
C303 B.n263 VSUBS 0.007361f
C304 B.n264 VSUBS 0.007361f
C305 B.n265 VSUBS 0.007361f
C306 B.n266 VSUBS 0.007361f
C307 B.n267 VSUBS 0.007361f
C308 B.n268 VSUBS 0.007361f
C309 B.n269 VSUBS 0.007361f
C310 B.n270 VSUBS 0.007361f
C311 B.n271 VSUBS 0.007361f
C312 B.n272 VSUBS 0.007361f
C313 B.n273 VSUBS 0.007361f
C314 B.n274 VSUBS 0.007361f
C315 B.n275 VSUBS 0.007361f
C316 B.n276 VSUBS 0.007361f
C317 B.n277 VSUBS 0.007361f
C318 B.n278 VSUBS 0.007361f
C319 B.n279 VSUBS 0.007361f
C320 B.n280 VSUBS 0.007361f
C321 B.n281 VSUBS 0.007361f
C322 B.n282 VSUBS 0.007361f
C323 B.n283 VSUBS 0.005087f
C324 B.n284 VSUBS 0.007361f
C325 B.n285 VSUBS 0.007361f
C326 B.n286 VSUBS 0.005953f
C327 B.n287 VSUBS 0.007361f
C328 B.n288 VSUBS 0.007361f
C329 B.n289 VSUBS 0.007361f
C330 B.n290 VSUBS 0.007361f
C331 B.n291 VSUBS 0.007361f
C332 B.n292 VSUBS 0.007361f
C333 B.n293 VSUBS 0.007361f
C334 B.n294 VSUBS 0.007361f
C335 B.n295 VSUBS 0.007361f
C336 B.n296 VSUBS 0.007361f
C337 B.n297 VSUBS 0.007361f
C338 B.n298 VSUBS 0.005953f
C339 B.n299 VSUBS 0.017054f
C340 B.n300 VSUBS 0.005087f
C341 B.n301 VSUBS 0.007361f
C342 B.n302 VSUBS 0.007361f
C343 B.n303 VSUBS 0.007361f
C344 B.n304 VSUBS 0.007361f
C345 B.n305 VSUBS 0.007361f
C346 B.n306 VSUBS 0.007361f
C347 B.n307 VSUBS 0.007361f
C348 B.n308 VSUBS 0.007361f
C349 B.n309 VSUBS 0.007361f
C350 B.n310 VSUBS 0.007361f
C351 B.n311 VSUBS 0.007361f
C352 B.n312 VSUBS 0.007361f
C353 B.n313 VSUBS 0.007361f
C354 B.n314 VSUBS 0.007361f
C355 B.n315 VSUBS 0.007361f
C356 B.n316 VSUBS 0.007361f
C357 B.n317 VSUBS 0.007361f
C358 B.n318 VSUBS 0.007361f
C359 B.n319 VSUBS 0.007361f
C360 B.n320 VSUBS 0.007361f
C361 B.n321 VSUBS 0.007361f
C362 B.n322 VSUBS 0.007361f
C363 B.n323 VSUBS 0.007361f
C364 B.n324 VSUBS 0.007361f
C365 B.n325 VSUBS 0.007361f
C366 B.n326 VSUBS 0.007361f
C367 B.n327 VSUBS 0.007361f
C368 B.n328 VSUBS 0.007361f
C369 B.n329 VSUBS 0.007361f
C370 B.n330 VSUBS 0.007361f
C371 B.n331 VSUBS 0.007361f
C372 B.n332 VSUBS 0.007361f
C373 B.n333 VSUBS 0.007361f
C374 B.n334 VSUBS 0.007361f
C375 B.n335 VSUBS 0.007361f
C376 B.n336 VSUBS 0.007361f
C377 B.n337 VSUBS 0.007361f
C378 B.n338 VSUBS 0.007361f
C379 B.n339 VSUBS 0.007361f
C380 B.n340 VSUBS 0.007361f
C381 B.n341 VSUBS 0.007361f
C382 B.n342 VSUBS 0.007361f
C383 B.n343 VSUBS 0.007361f
C384 B.n344 VSUBS 0.007361f
C385 B.n345 VSUBS 0.007361f
C386 B.n346 VSUBS 0.007361f
C387 B.n347 VSUBS 0.007361f
C388 B.n348 VSUBS 0.007361f
C389 B.n349 VSUBS 0.007361f
C390 B.n350 VSUBS 0.007361f
C391 B.n351 VSUBS 0.007361f
C392 B.n352 VSUBS 0.007361f
C393 B.n353 VSUBS 0.007361f
C394 B.n354 VSUBS 0.007361f
C395 B.n355 VSUBS 0.007361f
C396 B.n356 VSUBS 0.007361f
C397 B.n357 VSUBS 0.007361f
C398 B.n358 VSUBS 0.007361f
C399 B.n359 VSUBS 0.007361f
C400 B.n360 VSUBS 0.007361f
C401 B.n361 VSUBS 0.007361f
C402 B.n362 VSUBS 0.007361f
C403 B.n363 VSUBS 0.007361f
C404 B.n364 VSUBS 0.007361f
C405 B.n365 VSUBS 0.007361f
C406 B.n366 VSUBS 0.007361f
C407 B.n367 VSUBS 0.007361f
C408 B.n368 VSUBS 0.007361f
C409 B.n369 VSUBS 0.007361f
C410 B.n370 VSUBS 0.007361f
C411 B.n371 VSUBS 0.007361f
C412 B.n372 VSUBS 0.007361f
C413 B.n373 VSUBS 0.007361f
C414 B.n374 VSUBS 0.007361f
C415 B.n375 VSUBS 0.007361f
C416 B.n376 VSUBS 0.007361f
C417 B.n377 VSUBS 0.007361f
C418 B.n378 VSUBS 0.007361f
C419 B.n379 VSUBS 0.007361f
C420 B.n380 VSUBS 0.007361f
C421 B.n381 VSUBS 0.007361f
C422 B.n382 VSUBS 0.007361f
C423 B.n383 VSUBS 0.007361f
C424 B.n384 VSUBS 0.007361f
C425 B.n385 VSUBS 0.007361f
C426 B.n386 VSUBS 0.007361f
C427 B.n387 VSUBS 0.007361f
C428 B.n388 VSUBS 0.007361f
C429 B.n389 VSUBS 0.007361f
C430 B.n390 VSUBS 0.016678f
C431 B.n391 VSUBS 0.016012f
C432 B.n392 VSUBS 0.016012f
C433 B.n393 VSUBS 0.007361f
C434 B.n394 VSUBS 0.007361f
C435 B.n395 VSUBS 0.007361f
C436 B.n396 VSUBS 0.007361f
C437 B.n397 VSUBS 0.007361f
C438 B.n398 VSUBS 0.007361f
C439 B.n399 VSUBS 0.007361f
C440 B.n400 VSUBS 0.007361f
C441 B.n401 VSUBS 0.007361f
C442 B.n402 VSUBS 0.007361f
C443 B.n403 VSUBS 0.007361f
C444 B.n404 VSUBS 0.007361f
C445 B.n405 VSUBS 0.007361f
C446 B.n406 VSUBS 0.007361f
C447 B.n407 VSUBS 0.007361f
C448 B.n408 VSUBS 0.007361f
C449 B.n409 VSUBS 0.007361f
C450 B.n410 VSUBS 0.007361f
C451 B.n411 VSUBS 0.007361f
C452 B.n412 VSUBS 0.007361f
C453 B.n413 VSUBS 0.007361f
C454 B.n414 VSUBS 0.007361f
C455 B.n415 VSUBS 0.007361f
C456 B.n416 VSUBS 0.007361f
C457 B.n417 VSUBS 0.007361f
C458 B.n418 VSUBS 0.007361f
C459 B.n419 VSUBS 0.007361f
C460 B.n420 VSUBS 0.007361f
C461 B.n421 VSUBS 0.007361f
C462 B.n422 VSUBS 0.007361f
C463 B.n423 VSUBS 0.007361f
C464 B.n424 VSUBS 0.007361f
C465 B.n425 VSUBS 0.007361f
C466 B.n426 VSUBS 0.007361f
C467 B.n427 VSUBS 0.007361f
C468 B.n428 VSUBS 0.007361f
C469 B.n429 VSUBS 0.007361f
C470 B.n430 VSUBS 0.007361f
C471 B.n431 VSUBS 0.007361f
C472 B.n432 VSUBS 0.007361f
C473 B.n433 VSUBS 0.007361f
C474 B.n434 VSUBS 0.007361f
C475 B.n435 VSUBS 0.007361f
C476 B.n436 VSUBS 0.016012f
C477 B.n437 VSUBS 0.016954f
C478 B.n438 VSUBS 0.015736f
C479 B.n439 VSUBS 0.007361f
C480 B.n440 VSUBS 0.007361f
C481 B.n441 VSUBS 0.007361f
C482 B.n442 VSUBS 0.007361f
C483 B.n443 VSUBS 0.007361f
C484 B.n444 VSUBS 0.007361f
C485 B.n445 VSUBS 0.007361f
C486 B.n446 VSUBS 0.007361f
C487 B.n447 VSUBS 0.007361f
C488 B.n448 VSUBS 0.007361f
C489 B.n449 VSUBS 0.007361f
C490 B.n450 VSUBS 0.007361f
C491 B.n451 VSUBS 0.007361f
C492 B.n452 VSUBS 0.007361f
C493 B.n453 VSUBS 0.007361f
C494 B.n454 VSUBS 0.007361f
C495 B.n455 VSUBS 0.007361f
C496 B.n456 VSUBS 0.007361f
C497 B.n457 VSUBS 0.007361f
C498 B.n458 VSUBS 0.007361f
C499 B.n459 VSUBS 0.007361f
C500 B.n460 VSUBS 0.007361f
C501 B.n461 VSUBS 0.007361f
C502 B.n462 VSUBS 0.007361f
C503 B.n463 VSUBS 0.007361f
C504 B.n464 VSUBS 0.007361f
C505 B.n465 VSUBS 0.007361f
C506 B.n466 VSUBS 0.007361f
C507 B.n467 VSUBS 0.007361f
C508 B.n468 VSUBS 0.007361f
C509 B.n469 VSUBS 0.007361f
C510 B.n470 VSUBS 0.007361f
C511 B.n471 VSUBS 0.007361f
C512 B.n472 VSUBS 0.007361f
C513 B.n473 VSUBS 0.007361f
C514 B.n474 VSUBS 0.007361f
C515 B.n475 VSUBS 0.007361f
C516 B.n476 VSUBS 0.007361f
C517 B.n477 VSUBS 0.007361f
C518 B.n478 VSUBS 0.007361f
C519 B.n479 VSUBS 0.007361f
C520 B.n480 VSUBS 0.007361f
C521 B.n481 VSUBS 0.007361f
C522 B.n482 VSUBS 0.007361f
C523 B.n483 VSUBS 0.007361f
C524 B.n484 VSUBS 0.007361f
C525 B.n485 VSUBS 0.007361f
C526 B.n486 VSUBS 0.007361f
C527 B.n487 VSUBS 0.007361f
C528 B.n488 VSUBS 0.007361f
C529 B.n489 VSUBS 0.007361f
C530 B.n490 VSUBS 0.007361f
C531 B.n491 VSUBS 0.007361f
C532 B.n492 VSUBS 0.007361f
C533 B.n493 VSUBS 0.007361f
C534 B.n494 VSUBS 0.007361f
C535 B.n495 VSUBS 0.007361f
C536 B.n496 VSUBS 0.007361f
C537 B.n497 VSUBS 0.007361f
C538 B.n498 VSUBS 0.007361f
C539 B.n499 VSUBS 0.007361f
C540 B.n500 VSUBS 0.007361f
C541 B.n501 VSUBS 0.007361f
C542 B.n502 VSUBS 0.007361f
C543 B.n503 VSUBS 0.007361f
C544 B.n504 VSUBS 0.007361f
C545 B.n505 VSUBS 0.007361f
C546 B.n506 VSUBS 0.007361f
C547 B.n507 VSUBS 0.007361f
C548 B.n508 VSUBS 0.007361f
C549 B.n509 VSUBS 0.007361f
C550 B.n510 VSUBS 0.007361f
C551 B.n511 VSUBS 0.007361f
C552 B.n512 VSUBS 0.007361f
C553 B.n513 VSUBS 0.007361f
C554 B.n514 VSUBS 0.007361f
C555 B.n515 VSUBS 0.007361f
C556 B.n516 VSUBS 0.007361f
C557 B.n517 VSUBS 0.007361f
C558 B.n518 VSUBS 0.007361f
C559 B.n519 VSUBS 0.007361f
C560 B.n520 VSUBS 0.007361f
C561 B.n521 VSUBS 0.007361f
C562 B.n522 VSUBS 0.007361f
C563 B.n523 VSUBS 0.007361f
C564 B.n524 VSUBS 0.007361f
C565 B.n525 VSUBS 0.007361f
C566 B.n526 VSUBS 0.007361f
C567 B.n527 VSUBS 0.007361f
C568 B.n528 VSUBS 0.005087f
C569 B.n529 VSUBS 0.017054f
C570 B.n530 VSUBS 0.005953f
C571 B.n531 VSUBS 0.007361f
C572 B.n532 VSUBS 0.007361f
C573 B.n533 VSUBS 0.007361f
C574 B.n534 VSUBS 0.007361f
C575 B.n535 VSUBS 0.007361f
C576 B.n536 VSUBS 0.007361f
C577 B.n537 VSUBS 0.007361f
C578 B.n538 VSUBS 0.007361f
C579 B.n539 VSUBS 0.007361f
C580 B.n540 VSUBS 0.007361f
C581 B.n541 VSUBS 0.007361f
C582 B.n542 VSUBS 0.005953f
C583 B.n543 VSUBS 0.007361f
C584 B.n544 VSUBS 0.007361f
C585 B.n545 VSUBS 0.005087f
C586 B.n546 VSUBS 0.007361f
C587 B.n547 VSUBS 0.007361f
C588 B.n548 VSUBS 0.007361f
C589 B.n549 VSUBS 0.007361f
C590 B.n550 VSUBS 0.007361f
C591 B.n551 VSUBS 0.007361f
C592 B.n552 VSUBS 0.007361f
C593 B.n553 VSUBS 0.007361f
C594 B.n554 VSUBS 0.007361f
C595 B.n555 VSUBS 0.007361f
C596 B.n556 VSUBS 0.007361f
C597 B.n557 VSUBS 0.007361f
C598 B.n558 VSUBS 0.007361f
C599 B.n559 VSUBS 0.007361f
C600 B.n560 VSUBS 0.007361f
C601 B.n561 VSUBS 0.007361f
C602 B.n562 VSUBS 0.007361f
C603 B.n563 VSUBS 0.007361f
C604 B.n564 VSUBS 0.007361f
C605 B.n565 VSUBS 0.007361f
C606 B.n566 VSUBS 0.007361f
C607 B.n567 VSUBS 0.007361f
C608 B.n568 VSUBS 0.007361f
C609 B.n569 VSUBS 0.007361f
C610 B.n570 VSUBS 0.007361f
C611 B.n571 VSUBS 0.007361f
C612 B.n572 VSUBS 0.007361f
C613 B.n573 VSUBS 0.007361f
C614 B.n574 VSUBS 0.007361f
C615 B.n575 VSUBS 0.007361f
C616 B.n576 VSUBS 0.007361f
C617 B.n577 VSUBS 0.007361f
C618 B.n578 VSUBS 0.007361f
C619 B.n579 VSUBS 0.007361f
C620 B.n580 VSUBS 0.007361f
C621 B.n581 VSUBS 0.007361f
C622 B.n582 VSUBS 0.007361f
C623 B.n583 VSUBS 0.007361f
C624 B.n584 VSUBS 0.007361f
C625 B.n585 VSUBS 0.007361f
C626 B.n586 VSUBS 0.007361f
C627 B.n587 VSUBS 0.007361f
C628 B.n588 VSUBS 0.007361f
C629 B.n589 VSUBS 0.007361f
C630 B.n590 VSUBS 0.007361f
C631 B.n591 VSUBS 0.007361f
C632 B.n592 VSUBS 0.007361f
C633 B.n593 VSUBS 0.007361f
C634 B.n594 VSUBS 0.007361f
C635 B.n595 VSUBS 0.007361f
C636 B.n596 VSUBS 0.007361f
C637 B.n597 VSUBS 0.007361f
C638 B.n598 VSUBS 0.007361f
C639 B.n599 VSUBS 0.007361f
C640 B.n600 VSUBS 0.007361f
C641 B.n601 VSUBS 0.007361f
C642 B.n602 VSUBS 0.007361f
C643 B.n603 VSUBS 0.007361f
C644 B.n604 VSUBS 0.007361f
C645 B.n605 VSUBS 0.007361f
C646 B.n606 VSUBS 0.007361f
C647 B.n607 VSUBS 0.007361f
C648 B.n608 VSUBS 0.007361f
C649 B.n609 VSUBS 0.007361f
C650 B.n610 VSUBS 0.007361f
C651 B.n611 VSUBS 0.007361f
C652 B.n612 VSUBS 0.007361f
C653 B.n613 VSUBS 0.007361f
C654 B.n614 VSUBS 0.007361f
C655 B.n615 VSUBS 0.007361f
C656 B.n616 VSUBS 0.007361f
C657 B.n617 VSUBS 0.007361f
C658 B.n618 VSUBS 0.007361f
C659 B.n619 VSUBS 0.007361f
C660 B.n620 VSUBS 0.007361f
C661 B.n621 VSUBS 0.007361f
C662 B.n622 VSUBS 0.007361f
C663 B.n623 VSUBS 0.007361f
C664 B.n624 VSUBS 0.007361f
C665 B.n625 VSUBS 0.007361f
C666 B.n626 VSUBS 0.007361f
C667 B.n627 VSUBS 0.007361f
C668 B.n628 VSUBS 0.007361f
C669 B.n629 VSUBS 0.007361f
C670 B.n630 VSUBS 0.007361f
C671 B.n631 VSUBS 0.007361f
C672 B.n632 VSUBS 0.007361f
C673 B.n633 VSUBS 0.007361f
C674 B.n634 VSUBS 0.016678f
C675 B.n635 VSUBS 0.016678f
C676 B.n636 VSUBS 0.016012f
C677 B.n637 VSUBS 0.007361f
C678 B.n638 VSUBS 0.007361f
C679 B.n639 VSUBS 0.007361f
C680 B.n640 VSUBS 0.007361f
C681 B.n641 VSUBS 0.007361f
C682 B.n642 VSUBS 0.007361f
C683 B.n643 VSUBS 0.007361f
C684 B.n644 VSUBS 0.007361f
C685 B.n645 VSUBS 0.007361f
C686 B.n646 VSUBS 0.007361f
C687 B.n647 VSUBS 0.007361f
C688 B.n648 VSUBS 0.007361f
C689 B.n649 VSUBS 0.007361f
C690 B.n650 VSUBS 0.007361f
C691 B.n651 VSUBS 0.007361f
C692 B.n652 VSUBS 0.007361f
C693 B.n653 VSUBS 0.007361f
C694 B.n654 VSUBS 0.007361f
C695 B.n655 VSUBS 0.007361f
C696 B.n656 VSUBS 0.007361f
C697 B.n657 VSUBS 0.007361f
C698 B.n658 VSUBS 0.007361f
C699 B.n659 VSUBS 0.016667f
C700 VDD2.t5 VSUBS 5.08737f
C701 VDD2.t0 VSUBS 0.472101f
C702 VDD2.t4 VSUBS 0.472101f
C703 VDD2.n0 VSUBS 3.91931f
C704 VDD2.n1 VSUBS 3.7674f
C705 VDD2.t1 VSUBS 5.08361f
C706 VDD2.n2 VSUBS 3.85741f
C707 VDD2.t2 VSUBS 0.472101f
C708 VDD2.t3 VSUBS 0.472101f
C709 VDD2.n3 VSUBS 3.91926f
C710 VN.t0 VSUBS 0.900359f
C711 VN.n0 VSUBS 0.360406f
C712 VN.t5 VSUBS 0.892511f
C713 VN.n1 VSUBS 0.338735f
C714 VN.t1 VSUBS 0.900359f
C715 VN.n2 VSUBS 0.360303f
C716 VN.n3 VSUBS 0.143396f
C717 VN.t2 VSUBS 0.900359f
C718 VN.n4 VSUBS 0.360406f
C719 VN.t4 VSUBS 0.900359f
C720 VN.t3 VSUBS 0.892511f
C721 VN.n5 VSUBS 0.338735f
C722 VN.n6 VSUBS 0.360303f
C723 VN.n7 VSUBS 3.36487f
C724 VDD1.t1 VSUBS 5.08535f
C725 VDD1.t5 VSUBS 5.0839f
C726 VDD1.t0 VSUBS 0.471779f
C727 VDD1.t2 VSUBS 0.471779f
C728 VDD1.n0 VSUBS 3.91664f
C729 VDD1.n1 VSUBS 3.85196f
C730 VDD1.t4 VSUBS 0.471779f
C731 VDD1.t3 VSUBS 0.471779f
C732 VDD1.n2 VSUBS 3.91587f
C733 VDD1.n3 VSUBS 3.77802f
C734 VTAIL.t2 VSUBS 0.50255f
C735 VTAIL.t3 VSUBS 0.50255f
C736 VTAIL.n0 VSUBS 3.9384f
C737 VTAIL.n1 VSUBS 0.983647f
C738 VTAIL.t6 VSUBS 5.14413f
C739 VTAIL.n2 VSUBS 1.18292f
C740 VTAIL.t9 VSUBS 0.50255f
C741 VTAIL.t11 VSUBS 0.50255f
C742 VTAIL.n3 VSUBS 3.9384f
C743 VTAIL.n4 VSUBS 3.28169f
C744 VTAIL.t4 VSUBS 0.50255f
C745 VTAIL.t5 VSUBS 0.50255f
C746 VTAIL.n5 VSUBS 3.93841f
C747 VTAIL.n6 VSUBS 3.28169f
C748 VTAIL.t0 VSUBS 5.14417f
C749 VTAIL.n7 VSUBS 1.18288f
C750 VTAIL.t7 VSUBS 0.50255f
C751 VTAIL.t8 VSUBS 0.50255f
C752 VTAIL.n8 VSUBS 3.93841f
C753 VTAIL.n9 VSUBS 1.01805f
C754 VTAIL.t10 VSUBS 5.14413f
C755 VTAIL.n10 VSUBS 3.39207f
C756 VTAIL.t1 VSUBS 5.14413f
C757 VTAIL.n11 VSUBS 3.372f
C758 VP.t4 VSUBS 0.919406f
C759 VP.n0 VSUBS 0.36803f
C760 VP.t1 VSUBS 0.911392f
C761 VP.n1 VSUBS 0.345901f
C762 VP.t2 VSUBS 0.919406f
C763 VP.n2 VSUBS 0.367925f
C764 VP.n3 VSUBS 3.38834f
C765 VP.n4 VSUBS 3.35763f
C766 VP.t5 VSUBS 0.911392f
C767 VP.t0 VSUBS 0.919406f
C768 VP.n5 VSUBS 0.367925f
C769 VP.n6 VSUBS 0.345901f
C770 VP.t3 VSUBS 0.919406f
C771 VP.n7 VSUBS 0.367925f
C772 VP.n8 VSUBS 0.056518f
.ends

