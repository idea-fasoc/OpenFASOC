* NGSPICE file created from diff_pair_sample_0137.ext - technology: sky130A

.subckt diff_pair_sample_0137 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=3.29505 ps=20.3 w=19.97 l=3.55
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=0 ps=0 w=19.97 l=3.55
X2 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=3.29505 ps=20.3 w=19.97 l=3.55
X3 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=3.29505 ps=20.3 w=19.97 l=3.55
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=0 ps=0 w=19.97 l=3.55
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=0 ps=0 w=19.97 l=3.55
X6 VTAIL.t6 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=3.29505 ps=20.3 w=19.97 l=3.55
X7 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.29505 pd=20.3 as=7.7883 ps=40.72 w=19.97 l=3.55
X8 VDD2.t1 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.29505 pd=20.3 as=7.7883 ps=40.72 w=19.97 l=3.55
X9 VDD2.t0 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29505 pd=20.3 as=7.7883 ps=40.72 w=19.97 l=3.55
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7883 pd=40.72 as=0 ps=0 w=19.97 l=3.55
X11 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29505 pd=20.3 as=7.7883 ps=40.72 w=19.97 l=3.55
R0 VN.n1 VN.t3 170.238
R1 VN.n0 VN.t1 170.238
R2 VN.n0 VN.t2 169.006
R3 VN.n1 VN.t0 169.006
R4 VN VN.n1 57.6382
R5 VN VN.n0 2.14959
R6 VDD2.n2 VDD2.n0 110.201
R7 VDD2.n2 VDD2.n1 59.2366
R8 VDD2.n1 VDD2.t3 0.991987
R9 VDD2.n1 VDD2.t0 0.991987
R10 VDD2.n0 VDD2.t2 0.991987
R11 VDD2.n0 VDD2.t1 0.991987
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n6 VTAIL.t1 43.5493
R14 VTAIL.n5 VTAIL.t3 43.5493
R15 VTAIL.n4 VTAIL.t4 43.5493
R16 VTAIL.n3 VTAIL.t7 43.5493
R17 VTAIL.n7 VTAIL.t5 43.5492
R18 VTAIL.n0 VTAIL.t6 43.5492
R19 VTAIL.n1 VTAIL.t0 43.5492
R20 VTAIL.n2 VTAIL.t2 43.5492
R21 VTAIL.n7 VTAIL.n6 32.9272
R22 VTAIL.n3 VTAIL.n2 32.9272
R23 VTAIL.n4 VTAIL.n3 3.34533
R24 VTAIL.n6 VTAIL.n5 3.34533
R25 VTAIL.n2 VTAIL.n1 3.34533
R26 VTAIL VTAIL.n0 1.7311
R27 VTAIL VTAIL.n7 1.61472
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n774 B.n773 585
R31 B.n776 B.n154 585
R32 B.n779 B.n778 585
R33 B.n780 B.n153 585
R34 B.n782 B.n781 585
R35 B.n784 B.n152 585
R36 B.n787 B.n786 585
R37 B.n788 B.n151 585
R38 B.n790 B.n789 585
R39 B.n792 B.n150 585
R40 B.n795 B.n794 585
R41 B.n796 B.n149 585
R42 B.n798 B.n797 585
R43 B.n800 B.n148 585
R44 B.n803 B.n802 585
R45 B.n804 B.n147 585
R46 B.n806 B.n805 585
R47 B.n808 B.n146 585
R48 B.n811 B.n810 585
R49 B.n812 B.n145 585
R50 B.n814 B.n813 585
R51 B.n816 B.n144 585
R52 B.n819 B.n818 585
R53 B.n820 B.n143 585
R54 B.n822 B.n821 585
R55 B.n824 B.n142 585
R56 B.n827 B.n826 585
R57 B.n828 B.n141 585
R58 B.n830 B.n829 585
R59 B.n832 B.n140 585
R60 B.n835 B.n834 585
R61 B.n836 B.n139 585
R62 B.n838 B.n837 585
R63 B.n840 B.n138 585
R64 B.n843 B.n842 585
R65 B.n844 B.n137 585
R66 B.n846 B.n845 585
R67 B.n848 B.n136 585
R68 B.n851 B.n850 585
R69 B.n852 B.n135 585
R70 B.n854 B.n853 585
R71 B.n856 B.n134 585
R72 B.n859 B.n858 585
R73 B.n860 B.n133 585
R74 B.n862 B.n861 585
R75 B.n864 B.n132 585
R76 B.n867 B.n866 585
R77 B.n868 B.n131 585
R78 B.n870 B.n869 585
R79 B.n872 B.n130 585
R80 B.n875 B.n874 585
R81 B.n876 B.n129 585
R82 B.n878 B.n877 585
R83 B.n880 B.n128 585
R84 B.n883 B.n882 585
R85 B.n884 B.n127 585
R86 B.n886 B.n885 585
R87 B.n888 B.n126 585
R88 B.n891 B.n890 585
R89 B.n892 B.n125 585
R90 B.n894 B.n893 585
R91 B.n896 B.n124 585
R92 B.n899 B.n898 585
R93 B.n900 B.n120 585
R94 B.n902 B.n901 585
R95 B.n904 B.n119 585
R96 B.n907 B.n906 585
R97 B.n908 B.n118 585
R98 B.n910 B.n909 585
R99 B.n912 B.n117 585
R100 B.n915 B.n914 585
R101 B.n916 B.n116 585
R102 B.n918 B.n917 585
R103 B.n920 B.n115 585
R104 B.n923 B.n922 585
R105 B.n925 B.n112 585
R106 B.n927 B.n926 585
R107 B.n929 B.n111 585
R108 B.n932 B.n931 585
R109 B.n933 B.n110 585
R110 B.n935 B.n934 585
R111 B.n937 B.n109 585
R112 B.n940 B.n939 585
R113 B.n941 B.n108 585
R114 B.n943 B.n942 585
R115 B.n945 B.n107 585
R116 B.n948 B.n947 585
R117 B.n949 B.n106 585
R118 B.n951 B.n950 585
R119 B.n953 B.n105 585
R120 B.n956 B.n955 585
R121 B.n957 B.n104 585
R122 B.n959 B.n958 585
R123 B.n961 B.n103 585
R124 B.n964 B.n963 585
R125 B.n965 B.n102 585
R126 B.n967 B.n966 585
R127 B.n969 B.n101 585
R128 B.n972 B.n971 585
R129 B.n973 B.n100 585
R130 B.n975 B.n974 585
R131 B.n977 B.n99 585
R132 B.n980 B.n979 585
R133 B.n981 B.n98 585
R134 B.n983 B.n982 585
R135 B.n985 B.n97 585
R136 B.n988 B.n987 585
R137 B.n989 B.n96 585
R138 B.n991 B.n990 585
R139 B.n993 B.n95 585
R140 B.n996 B.n995 585
R141 B.n997 B.n94 585
R142 B.n999 B.n998 585
R143 B.n1001 B.n93 585
R144 B.n1004 B.n1003 585
R145 B.n1005 B.n92 585
R146 B.n1007 B.n1006 585
R147 B.n1009 B.n91 585
R148 B.n1012 B.n1011 585
R149 B.n1013 B.n90 585
R150 B.n1015 B.n1014 585
R151 B.n1017 B.n89 585
R152 B.n1020 B.n1019 585
R153 B.n1021 B.n88 585
R154 B.n1023 B.n1022 585
R155 B.n1025 B.n87 585
R156 B.n1028 B.n1027 585
R157 B.n1029 B.n86 585
R158 B.n1031 B.n1030 585
R159 B.n1033 B.n85 585
R160 B.n1036 B.n1035 585
R161 B.n1037 B.n84 585
R162 B.n1039 B.n1038 585
R163 B.n1041 B.n83 585
R164 B.n1044 B.n1043 585
R165 B.n1045 B.n82 585
R166 B.n1047 B.n1046 585
R167 B.n1049 B.n81 585
R168 B.n1052 B.n1051 585
R169 B.n1053 B.n80 585
R170 B.n772 B.n78 585
R171 B.n1056 B.n78 585
R172 B.n771 B.n77 585
R173 B.n1057 B.n77 585
R174 B.n770 B.n76 585
R175 B.n1058 B.n76 585
R176 B.n769 B.n768 585
R177 B.n768 B.n72 585
R178 B.n767 B.n71 585
R179 B.n1064 B.n71 585
R180 B.n766 B.n70 585
R181 B.n1065 B.n70 585
R182 B.n765 B.n69 585
R183 B.n1066 B.n69 585
R184 B.n764 B.n763 585
R185 B.n763 B.n65 585
R186 B.n762 B.n64 585
R187 B.n1072 B.n64 585
R188 B.n761 B.n63 585
R189 B.n1073 B.n63 585
R190 B.n760 B.n62 585
R191 B.n1074 B.n62 585
R192 B.n759 B.n758 585
R193 B.n758 B.n58 585
R194 B.n757 B.n57 585
R195 B.n1080 B.n57 585
R196 B.n756 B.n56 585
R197 B.n1081 B.n56 585
R198 B.n755 B.n55 585
R199 B.n1082 B.n55 585
R200 B.n754 B.n753 585
R201 B.n753 B.n51 585
R202 B.n752 B.n50 585
R203 B.n1088 B.n50 585
R204 B.n751 B.n49 585
R205 B.n1089 B.n49 585
R206 B.n750 B.n48 585
R207 B.n1090 B.n48 585
R208 B.n749 B.n748 585
R209 B.n748 B.n44 585
R210 B.n747 B.n43 585
R211 B.n1096 B.n43 585
R212 B.n746 B.n42 585
R213 B.n1097 B.n42 585
R214 B.n745 B.n41 585
R215 B.n1098 B.n41 585
R216 B.n744 B.n743 585
R217 B.n743 B.n40 585
R218 B.n742 B.n36 585
R219 B.n1104 B.n36 585
R220 B.n741 B.n35 585
R221 B.n1105 B.n35 585
R222 B.n740 B.n34 585
R223 B.n1106 B.n34 585
R224 B.n739 B.n738 585
R225 B.n738 B.n30 585
R226 B.n737 B.n29 585
R227 B.n1112 B.n29 585
R228 B.n736 B.n28 585
R229 B.n1113 B.n28 585
R230 B.n735 B.n27 585
R231 B.n1114 B.n27 585
R232 B.n734 B.n733 585
R233 B.n733 B.n23 585
R234 B.n732 B.n22 585
R235 B.n1120 B.n22 585
R236 B.n731 B.n21 585
R237 B.n1121 B.n21 585
R238 B.n730 B.n20 585
R239 B.n1122 B.n20 585
R240 B.n729 B.n728 585
R241 B.n728 B.n19 585
R242 B.n727 B.n15 585
R243 B.n1128 B.n15 585
R244 B.n726 B.n14 585
R245 B.n1129 B.n14 585
R246 B.n725 B.n13 585
R247 B.n1130 B.n13 585
R248 B.n724 B.n723 585
R249 B.n723 B.n12 585
R250 B.n722 B.n721 585
R251 B.n722 B.n8 585
R252 B.n720 B.n7 585
R253 B.n1137 B.n7 585
R254 B.n719 B.n6 585
R255 B.n1138 B.n6 585
R256 B.n718 B.n5 585
R257 B.n1139 B.n5 585
R258 B.n717 B.n716 585
R259 B.n716 B.n4 585
R260 B.n715 B.n155 585
R261 B.n715 B.n714 585
R262 B.n705 B.n156 585
R263 B.n157 B.n156 585
R264 B.n707 B.n706 585
R265 B.n708 B.n707 585
R266 B.n704 B.n162 585
R267 B.n162 B.n161 585
R268 B.n703 B.n702 585
R269 B.n702 B.n701 585
R270 B.n164 B.n163 585
R271 B.n694 B.n164 585
R272 B.n693 B.n692 585
R273 B.n695 B.n693 585
R274 B.n691 B.n169 585
R275 B.n169 B.n168 585
R276 B.n690 B.n689 585
R277 B.n689 B.n688 585
R278 B.n171 B.n170 585
R279 B.n172 B.n171 585
R280 B.n681 B.n680 585
R281 B.n682 B.n681 585
R282 B.n679 B.n177 585
R283 B.n177 B.n176 585
R284 B.n678 B.n677 585
R285 B.n677 B.n676 585
R286 B.n179 B.n178 585
R287 B.n180 B.n179 585
R288 B.n669 B.n668 585
R289 B.n670 B.n669 585
R290 B.n667 B.n185 585
R291 B.n185 B.n184 585
R292 B.n666 B.n665 585
R293 B.n665 B.n664 585
R294 B.n187 B.n186 585
R295 B.n657 B.n187 585
R296 B.n656 B.n655 585
R297 B.n658 B.n656 585
R298 B.n654 B.n192 585
R299 B.n192 B.n191 585
R300 B.n653 B.n652 585
R301 B.n652 B.n651 585
R302 B.n194 B.n193 585
R303 B.n195 B.n194 585
R304 B.n644 B.n643 585
R305 B.n645 B.n644 585
R306 B.n642 B.n200 585
R307 B.n200 B.n199 585
R308 B.n641 B.n640 585
R309 B.n640 B.n639 585
R310 B.n202 B.n201 585
R311 B.n203 B.n202 585
R312 B.n632 B.n631 585
R313 B.n633 B.n632 585
R314 B.n630 B.n208 585
R315 B.n208 B.n207 585
R316 B.n629 B.n628 585
R317 B.n628 B.n627 585
R318 B.n210 B.n209 585
R319 B.n211 B.n210 585
R320 B.n620 B.n619 585
R321 B.n621 B.n620 585
R322 B.n618 B.n215 585
R323 B.n219 B.n215 585
R324 B.n617 B.n616 585
R325 B.n616 B.n615 585
R326 B.n217 B.n216 585
R327 B.n218 B.n217 585
R328 B.n608 B.n607 585
R329 B.n609 B.n608 585
R330 B.n606 B.n224 585
R331 B.n224 B.n223 585
R332 B.n605 B.n604 585
R333 B.n604 B.n603 585
R334 B.n226 B.n225 585
R335 B.n227 B.n226 585
R336 B.n596 B.n595 585
R337 B.n597 B.n596 585
R338 B.n594 B.n232 585
R339 B.n232 B.n231 585
R340 B.n593 B.n592 585
R341 B.n592 B.n591 585
R342 B.n588 B.n236 585
R343 B.n587 B.n586 585
R344 B.n584 B.n237 585
R345 B.n584 B.n235 585
R346 B.n583 B.n582 585
R347 B.n581 B.n580 585
R348 B.n579 B.n239 585
R349 B.n577 B.n576 585
R350 B.n575 B.n240 585
R351 B.n574 B.n573 585
R352 B.n571 B.n241 585
R353 B.n569 B.n568 585
R354 B.n567 B.n242 585
R355 B.n566 B.n565 585
R356 B.n563 B.n243 585
R357 B.n561 B.n560 585
R358 B.n559 B.n244 585
R359 B.n558 B.n557 585
R360 B.n555 B.n245 585
R361 B.n553 B.n552 585
R362 B.n551 B.n246 585
R363 B.n550 B.n549 585
R364 B.n547 B.n247 585
R365 B.n545 B.n544 585
R366 B.n543 B.n248 585
R367 B.n542 B.n541 585
R368 B.n539 B.n249 585
R369 B.n537 B.n536 585
R370 B.n535 B.n250 585
R371 B.n534 B.n533 585
R372 B.n531 B.n251 585
R373 B.n529 B.n528 585
R374 B.n527 B.n252 585
R375 B.n526 B.n525 585
R376 B.n523 B.n253 585
R377 B.n521 B.n520 585
R378 B.n519 B.n254 585
R379 B.n518 B.n517 585
R380 B.n515 B.n255 585
R381 B.n513 B.n512 585
R382 B.n511 B.n256 585
R383 B.n510 B.n509 585
R384 B.n507 B.n257 585
R385 B.n505 B.n504 585
R386 B.n503 B.n258 585
R387 B.n502 B.n501 585
R388 B.n499 B.n259 585
R389 B.n497 B.n496 585
R390 B.n495 B.n260 585
R391 B.n494 B.n493 585
R392 B.n491 B.n261 585
R393 B.n489 B.n488 585
R394 B.n487 B.n262 585
R395 B.n486 B.n485 585
R396 B.n483 B.n263 585
R397 B.n481 B.n480 585
R398 B.n479 B.n264 585
R399 B.n478 B.n477 585
R400 B.n475 B.n265 585
R401 B.n473 B.n472 585
R402 B.n471 B.n266 585
R403 B.n470 B.n469 585
R404 B.n467 B.n267 585
R405 B.n465 B.n464 585
R406 B.n463 B.n268 585
R407 B.n462 B.n461 585
R408 B.n459 B.n458 585
R409 B.n457 B.n456 585
R410 B.n455 B.n273 585
R411 B.n453 B.n452 585
R412 B.n451 B.n274 585
R413 B.n450 B.n449 585
R414 B.n447 B.n275 585
R415 B.n445 B.n444 585
R416 B.n443 B.n276 585
R417 B.n442 B.n441 585
R418 B.n439 B.n438 585
R419 B.n437 B.n436 585
R420 B.n435 B.n281 585
R421 B.n433 B.n432 585
R422 B.n431 B.n282 585
R423 B.n430 B.n429 585
R424 B.n427 B.n283 585
R425 B.n425 B.n424 585
R426 B.n423 B.n284 585
R427 B.n422 B.n421 585
R428 B.n419 B.n285 585
R429 B.n417 B.n416 585
R430 B.n415 B.n286 585
R431 B.n414 B.n413 585
R432 B.n411 B.n287 585
R433 B.n409 B.n408 585
R434 B.n407 B.n288 585
R435 B.n406 B.n405 585
R436 B.n403 B.n289 585
R437 B.n401 B.n400 585
R438 B.n399 B.n290 585
R439 B.n398 B.n397 585
R440 B.n395 B.n291 585
R441 B.n393 B.n392 585
R442 B.n391 B.n292 585
R443 B.n390 B.n389 585
R444 B.n387 B.n293 585
R445 B.n385 B.n384 585
R446 B.n383 B.n294 585
R447 B.n382 B.n381 585
R448 B.n379 B.n295 585
R449 B.n377 B.n376 585
R450 B.n375 B.n296 585
R451 B.n374 B.n373 585
R452 B.n371 B.n297 585
R453 B.n369 B.n368 585
R454 B.n367 B.n298 585
R455 B.n366 B.n365 585
R456 B.n363 B.n299 585
R457 B.n361 B.n360 585
R458 B.n359 B.n300 585
R459 B.n358 B.n357 585
R460 B.n355 B.n301 585
R461 B.n353 B.n352 585
R462 B.n351 B.n302 585
R463 B.n350 B.n349 585
R464 B.n347 B.n303 585
R465 B.n345 B.n344 585
R466 B.n343 B.n304 585
R467 B.n342 B.n341 585
R468 B.n339 B.n305 585
R469 B.n337 B.n336 585
R470 B.n335 B.n306 585
R471 B.n334 B.n333 585
R472 B.n331 B.n307 585
R473 B.n329 B.n328 585
R474 B.n327 B.n308 585
R475 B.n326 B.n325 585
R476 B.n323 B.n309 585
R477 B.n321 B.n320 585
R478 B.n319 B.n310 585
R479 B.n318 B.n317 585
R480 B.n315 B.n311 585
R481 B.n313 B.n312 585
R482 B.n234 B.n233 585
R483 B.n235 B.n234 585
R484 B.n590 B.n589 585
R485 B.n591 B.n590 585
R486 B.n230 B.n229 585
R487 B.n231 B.n230 585
R488 B.n599 B.n598 585
R489 B.n598 B.n597 585
R490 B.n600 B.n228 585
R491 B.n228 B.n227 585
R492 B.n602 B.n601 585
R493 B.n603 B.n602 585
R494 B.n222 B.n221 585
R495 B.n223 B.n222 585
R496 B.n611 B.n610 585
R497 B.n610 B.n609 585
R498 B.n612 B.n220 585
R499 B.n220 B.n218 585
R500 B.n614 B.n613 585
R501 B.n615 B.n614 585
R502 B.n214 B.n213 585
R503 B.n219 B.n214 585
R504 B.n623 B.n622 585
R505 B.n622 B.n621 585
R506 B.n624 B.n212 585
R507 B.n212 B.n211 585
R508 B.n626 B.n625 585
R509 B.n627 B.n626 585
R510 B.n206 B.n205 585
R511 B.n207 B.n206 585
R512 B.n635 B.n634 585
R513 B.n634 B.n633 585
R514 B.n636 B.n204 585
R515 B.n204 B.n203 585
R516 B.n638 B.n637 585
R517 B.n639 B.n638 585
R518 B.n198 B.n197 585
R519 B.n199 B.n198 585
R520 B.n647 B.n646 585
R521 B.n646 B.n645 585
R522 B.n648 B.n196 585
R523 B.n196 B.n195 585
R524 B.n650 B.n649 585
R525 B.n651 B.n650 585
R526 B.n190 B.n189 585
R527 B.n191 B.n190 585
R528 B.n660 B.n659 585
R529 B.n659 B.n658 585
R530 B.n661 B.n188 585
R531 B.n657 B.n188 585
R532 B.n663 B.n662 585
R533 B.n664 B.n663 585
R534 B.n183 B.n182 585
R535 B.n184 B.n183 585
R536 B.n672 B.n671 585
R537 B.n671 B.n670 585
R538 B.n673 B.n181 585
R539 B.n181 B.n180 585
R540 B.n675 B.n674 585
R541 B.n676 B.n675 585
R542 B.n175 B.n174 585
R543 B.n176 B.n175 585
R544 B.n684 B.n683 585
R545 B.n683 B.n682 585
R546 B.n685 B.n173 585
R547 B.n173 B.n172 585
R548 B.n687 B.n686 585
R549 B.n688 B.n687 585
R550 B.n167 B.n166 585
R551 B.n168 B.n167 585
R552 B.n697 B.n696 585
R553 B.n696 B.n695 585
R554 B.n698 B.n165 585
R555 B.n694 B.n165 585
R556 B.n700 B.n699 585
R557 B.n701 B.n700 585
R558 B.n160 B.n159 585
R559 B.n161 B.n160 585
R560 B.n710 B.n709 585
R561 B.n709 B.n708 585
R562 B.n711 B.n158 585
R563 B.n158 B.n157 585
R564 B.n713 B.n712 585
R565 B.n714 B.n713 585
R566 B.n3 B.n0 585
R567 B.n4 B.n3 585
R568 B.n1136 B.n1 585
R569 B.n1137 B.n1136 585
R570 B.n1135 B.n1134 585
R571 B.n1135 B.n8 585
R572 B.n1133 B.n9 585
R573 B.n12 B.n9 585
R574 B.n1132 B.n1131 585
R575 B.n1131 B.n1130 585
R576 B.n11 B.n10 585
R577 B.n1129 B.n11 585
R578 B.n1127 B.n1126 585
R579 B.n1128 B.n1127 585
R580 B.n1125 B.n16 585
R581 B.n19 B.n16 585
R582 B.n1124 B.n1123 585
R583 B.n1123 B.n1122 585
R584 B.n18 B.n17 585
R585 B.n1121 B.n18 585
R586 B.n1119 B.n1118 585
R587 B.n1120 B.n1119 585
R588 B.n1117 B.n24 585
R589 B.n24 B.n23 585
R590 B.n1116 B.n1115 585
R591 B.n1115 B.n1114 585
R592 B.n26 B.n25 585
R593 B.n1113 B.n26 585
R594 B.n1111 B.n1110 585
R595 B.n1112 B.n1111 585
R596 B.n1109 B.n31 585
R597 B.n31 B.n30 585
R598 B.n1108 B.n1107 585
R599 B.n1107 B.n1106 585
R600 B.n33 B.n32 585
R601 B.n1105 B.n33 585
R602 B.n1103 B.n1102 585
R603 B.n1104 B.n1103 585
R604 B.n1101 B.n37 585
R605 B.n40 B.n37 585
R606 B.n1100 B.n1099 585
R607 B.n1099 B.n1098 585
R608 B.n39 B.n38 585
R609 B.n1097 B.n39 585
R610 B.n1095 B.n1094 585
R611 B.n1096 B.n1095 585
R612 B.n1093 B.n45 585
R613 B.n45 B.n44 585
R614 B.n1092 B.n1091 585
R615 B.n1091 B.n1090 585
R616 B.n47 B.n46 585
R617 B.n1089 B.n47 585
R618 B.n1087 B.n1086 585
R619 B.n1088 B.n1087 585
R620 B.n1085 B.n52 585
R621 B.n52 B.n51 585
R622 B.n1084 B.n1083 585
R623 B.n1083 B.n1082 585
R624 B.n54 B.n53 585
R625 B.n1081 B.n54 585
R626 B.n1079 B.n1078 585
R627 B.n1080 B.n1079 585
R628 B.n1077 B.n59 585
R629 B.n59 B.n58 585
R630 B.n1076 B.n1075 585
R631 B.n1075 B.n1074 585
R632 B.n61 B.n60 585
R633 B.n1073 B.n61 585
R634 B.n1071 B.n1070 585
R635 B.n1072 B.n1071 585
R636 B.n1069 B.n66 585
R637 B.n66 B.n65 585
R638 B.n1068 B.n1067 585
R639 B.n1067 B.n1066 585
R640 B.n68 B.n67 585
R641 B.n1065 B.n68 585
R642 B.n1063 B.n1062 585
R643 B.n1064 B.n1063 585
R644 B.n1061 B.n73 585
R645 B.n73 B.n72 585
R646 B.n1060 B.n1059 585
R647 B.n1059 B.n1058 585
R648 B.n75 B.n74 585
R649 B.n1057 B.n75 585
R650 B.n1055 B.n1054 585
R651 B.n1056 B.n1055 585
R652 B.n1140 B.n1139 585
R653 B.n1138 B.n2 585
R654 B.n1055 B.n80 449.257
R655 B.n774 B.n78 449.257
R656 B.n592 B.n234 449.257
R657 B.n590 B.n236 449.257
R658 B.n113 B.t12 344.709
R659 B.n121 B.t8 344.709
R660 B.n277 B.t4 344.709
R661 B.n269 B.t15 344.709
R662 B.n775 B.n79 256.663
R663 B.n777 B.n79 256.663
R664 B.n783 B.n79 256.663
R665 B.n785 B.n79 256.663
R666 B.n791 B.n79 256.663
R667 B.n793 B.n79 256.663
R668 B.n799 B.n79 256.663
R669 B.n801 B.n79 256.663
R670 B.n807 B.n79 256.663
R671 B.n809 B.n79 256.663
R672 B.n815 B.n79 256.663
R673 B.n817 B.n79 256.663
R674 B.n823 B.n79 256.663
R675 B.n825 B.n79 256.663
R676 B.n831 B.n79 256.663
R677 B.n833 B.n79 256.663
R678 B.n839 B.n79 256.663
R679 B.n841 B.n79 256.663
R680 B.n847 B.n79 256.663
R681 B.n849 B.n79 256.663
R682 B.n855 B.n79 256.663
R683 B.n857 B.n79 256.663
R684 B.n863 B.n79 256.663
R685 B.n865 B.n79 256.663
R686 B.n871 B.n79 256.663
R687 B.n873 B.n79 256.663
R688 B.n879 B.n79 256.663
R689 B.n881 B.n79 256.663
R690 B.n887 B.n79 256.663
R691 B.n889 B.n79 256.663
R692 B.n895 B.n79 256.663
R693 B.n897 B.n79 256.663
R694 B.n903 B.n79 256.663
R695 B.n905 B.n79 256.663
R696 B.n911 B.n79 256.663
R697 B.n913 B.n79 256.663
R698 B.n919 B.n79 256.663
R699 B.n921 B.n79 256.663
R700 B.n928 B.n79 256.663
R701 B.n930 B.n79 256.663
R702 B.n936 B.n79 256.663
R703 B.n938 B.n79 256.663
R704 B.n944 B.n79 256.663
R705 B.n946 B.n79 256.663
R706 B.n952 B.n79 256.663
R707 B.n954 B.n79 256.663
R708 B.n960 B.n79 256.663
R709 B.n962 B.n79 256.663
R710 B.n968 B.n79 256.663
R711 B.n970 B.n79 256.663
R712 B.n976 B.n79 256.663
R713 B.n978 B.n79 256.663
R714 B.n984 B.n79 256.663
R715 B.n986 B.n79 256.663
R716 B.n992 B.n79 256.663
R717 B.n994 B.n79 256.663
R718 B.n1000 B.n79 256.663
R719 B.n1002 B.n79 256.663
R720 B.n1008 B.n79 256.663
R721 B.n1010 B.n79 256.663
R722 B.n1016 B.n79 256.663
R723 B.n1018 B.n79 256.663
R724 B.n1024 B.n79 256.663
R725 B.n1026 B.n79 256.663
R726 B.n1032 B.n79 256.663
R727 B.n1034 B.n79 256.663
R728 B.n1040 B.n79 256.663
R729 B.n1042 B.n79 256.663
R730 B.n1048 B.n79 256.663
R731 B.n1050 B.n79 256.663
R732 B.n585 B.n235 256.663
R733 B.n238 B.n235 256.663
R734 B.n578 B.n235 256.663
R735 B.n572 B.n235 256.663
R736 B.n570 B.n235 256.663
R737 B.n564 B.n235 256.663
R738 B.n562 B.n235 256.663
R739 B.n556 B.n235 256.663
R740 B.n554 B.n235 256.663
R741 B.n548 B.n235 256.663
R742 B.n546 B.n235 256.663
R743 B.n540 B.n235 256.663
R744 B.n538 B.n235 256.663
R745 B.n532 B.n235 256.663
R746 B.n530 B.n235 256.663
R747 B.n524 B.n235 256.663
R748 B.n522 B.n235 256.663
R749 B.n516 B.n235 256.663
R750 B.n514 B.n235 256.663
R751 B.n508 B.n235 256.663
R752 B.n506 B.n235 256.663
R753 B.n500 B.n235 256.663
R754 B.n498 B.n235 256.663
R755 B.n492 B.n235 256.663
R756 B.n490 B.n235 256.663
R757 B.n484 B.n235 256.663
R758 B.n482 B.n235 256.663
R759 B.n476 B.n235 256.663
R760 B.n474 B.n235 256.663
R761 B.n468 B.n235 256.663
R762 B.n466 B.n235 256.663
R763 B.n460 B.n235 256.663
R764 B.n272 B.n235 256.663
R765 B.n454 B.n235 256.663
R766 B.n448 B.n235 256.663
R767 B.n446 B.n235 256.663
R768 B.n440 B.n235 256.663
R769 B.n280 B.n235 256.663
R770 B.n434 B.n235 256.663
R771 B.n428 B.n235 256.663
R772 B.n426 B.n235 256.663
R773 B.n420 B.n235 256.663
R774 B.n418 B.n235 256.663
R775 B.n412 B.n235 256.663
R776 B.n410 B.n235 256.663
R777 B.n404 B.n235 256.663
R778 B.n402 B.n235 256.663
R779 B.n396 B.n235 256.663
R780 B.n394 B.n235 256.663
R781 B.n388 B.n235 256.663
R782 B.n386 B.n235 256.663
R783 B.n380 B.n235 256.663
R784 B.n378 B.n235 256.663
R785 B.n372 B.n235 256.663
R786 B.n370 B.n235 256.663
R787 B.n364 B.n235 256.663
R788 B.n362 B.n235 256.663
R789 B.n356 B.n235 256.663
R790 B.n354 B.n235 256.663
R791 B.n348 B.n235 256.663
R792 B.n346 B.n235 256.663
R793 B.n340 B.n235 256.663
R794 B.n338 B.n235 256.663
R795 B.n332 B.n235 256.663
R796 B.n330 B.n235 256.663
R797 B.n324 B.n235 256.663
R798 B.n322 B.n235 256.663
R799 B.n316 B.n235 256.663
R800 B.n314 B.n235 256.663
R801 B.n1142 B.n1141 256.663
R802 B.n1051 B.n1049 163.367
R803 B.n1047 B.n82 163.367
R804 B.n1043 B.n1041 163.367
R805 B.n1039 B.n84 163.367
R806 B.n1035 B.n1033 163.367
R807 B.n1031 B.n86 163.367
R808 B.n1027 B.n1025 163.367
R809 B.n1023 B.n88 163.367
R810 B.n1019 B.n1017 163.367
R811 B.n1015 B.n90 163.367
R812 B.n1011 B.n1009 163.367
R813 B.n1007 B.n92 163.367
R814 B.n1003 B.n1001 163.367
R815 B.n999 B.n94 163.367
R816 B.n995 B.n993 163.367
R817 B.n991 B.n96 163.367
R818 B.n987 B.n985 163.367
R819 B.n983 B.n98 163.367
R820 B.n979 B.n977 163.367
R821 B.n975 B.n100 163.367
R822 B.n971 B.n969 163.367
R823 B.n967 B.n102 163.367
R824 B.n963 B.n961 163.367
R825 B.n959 B.n104 163.367
R826 B.n955 B.n953 163.367
R827 B.n951 B.n106 163.367
R828 B.n947 B.n945 163.367
R829 B.n943 B.n108 163.367
R830 B.n939 B.n937 163.367
R831 B.n935 B.n110 163.367
R832 B.n931 B.n929 163.367
R833 B.n927 B.n112 163.367
R834 B.n922 B.n920 163.367
R835 B.n918 B.n116 163.367
R836 B.n914 B.n912 163.367
R837 B.n910 B.n118 163.367
R838 B.n906 B.n904 163.367
R839 B.n902 B.n120 163.367
R840 B.n898 B.n896 163.367
R841 B.n894 B.n125 163.367
R842 B.n890 B.n888 163.367
R843 B.n886 B.n127 163.367
R844 B.n882 B.n880 163.367
R845 B.n878 B.n129 163.367
R846 B.n874 B.n872 163.367
R847 B.n870 B.n131 163.367
R848 B.n866 B.n864 163.367
R849 B.n862 B.n133 163.367
R850 B.n858 B.n856 163.367
R851 B.n854 B.n135 163.367
R852 B.n850 B.n848 163.367
R853 B.n846 B.n137 163.367
R854 B.n842 B.n840 163.367
R855 B.n838 B.n139 163.367
R856 B.n834 B.n832 163.367
R857 B.n830 B.n141 163.367
R858 B.n826 B.n824 163.367
R859 B.n822 B.n143 163.367
R860 B.n818 B.n816 163.367
R861 B.n814 B.n145 163.367
R862 B.n810 B.n808 163.367
R863 B.n806 B.n147 163.367
R864 B.n802 B.n800 163.367
R865 B.n798 B.n149 163.367
R866 B.n794 B.n792 163.367
R867 B.n790 B.n151 163.367
R868 B.n786 B.n784 163.367
R869 B.n782 B.n153 163.367
R870 B.n778 B.n776 163.367
R871 B.n592 B.n232 163.367
R872 B.n596 B.n232 163.367
R873 B.n596 B.n226 163.367
R874 B.n604 B.n226 163.367
R875 B.n604 B.n224 163.367
R876 B.n608 B.n224 163.367
R877 B.n608 B.n217 163.367
R878 B.n616 B.n217 163.367
R879 B.n616 B.n215 163.367
R880 B.n620 B.n215 163.367
R881 B.n620 B.n210 163.367
R882 B.n628 B.n210 163.367
R883 B.n628 B.n208 163.367
R884 B.n632 B.n208 163.367
R885 B.n632 B.n202 163.367
R886 B.n640 B.n202 163.367
R887 B.n640 B.n200 163.367
R888 B.n644 B.n200 163.367
R889 B.n644 B.n194 163.367
R890 B.n652 B.n194 163.367
R891 B.n652 B.n192 163.367
R892 B.n656 B.n192 163.367
R893 B.n656 B.n187 163.367
R894 B.n665 B.n187 163.367
R895 B.n665 B.n185 163.367
R896 B.n669 B.n185 163.367
R897 B.n669 B.n179 163.367
R898 B.n677 B.n179 163.367
R899 B.n677 B.n177 163.367
R900 B.n681 B.n177 163.367
R901 B.n681 B.n171 163.367
R902 B.n689 B.n171 163.367
R903 B.n689 B.n169 163.367
R904 B.n693 B.n169 163.367
R905 B.n693 B.n164 163.367
R906 B.n702 B.n164 163.367
R907 B.n702 B.n162 163.367
R908 B.n707 B.n162 163.367
R909 B.n707 B.n156 163.367
R910 B.n715 B.n156 163.367
R911 B.n716 B.n715 163.367
R912 B.n716 B.n5 163.367
R913 B.n6 B.n5 163.367
R914 B.n7 B.n6 163.367
R915 B.n722 B.n7 163.367
R916 B.n723 B.n722 163.367
R917 B.n723 B.n13 163.367
R918 B.n14 B.n13 163.367
R919 B.n15 B.n14 163.367
R920 B.n728 B.n15 163.367
R921 B.n728 B.n20 163.367
R922 B.n21 B.n20 163.367
R923 B.n22 B.n21 163.367
R924 B.n733 B.n22 163.367
R925 B.n733 B.n27 163.367
R926 B.n28 B.n27 163.367
R927 B.n29 B.n28 163.367
R928 B.n738 B.n29 163.367
R929 B.n738 B.n34 163.367
R930 B.n35 B.n34 163.367
R931 B.n36 B.n35 163.367
R932 B.n743 B.n36 163.367
R933 B.n743 B.n41 163.367
R934 B.n42 B.n41 163.367
R935 B.n43 B.n42 163.367
R936 B.n748 B.n43 163.367
R937 B.n748 B.n48 163.367
R938 B.n49 B.n48 163.367
R939 B.n50 B.n49 163.367
R940 B.n753 B.n50 163.367
R941 B.n753 B.n55 163.367
R942 B.n56 B.n55 163.367
R943 B.n57 B.n56 163.367
R944 B.n758 B.n57 163.367
R945 B.n758 B.n62 163.367
R946 B.n63 B.n62 163.367
R947 B.n64 B.n63 163.367
R948 B.n763 B.n64 163.367
R949 B.n763 B.n69 163.367
R950 B.n70 B.n69 163.367
R951 B.n71 B.n70 163.367
R952 B.n768 B.n71 163.367
R953 B.n768 B.n76 163.367
R954 B.n77 B.n76 163.367
R955 B.n78 B.n77 163.367
R956 B.n586 B.n584 163.367
R957 B.n584 B.n583 163.367
R958 B.n580 B.n579 163.367
R959 B.n577 B.n240 163.367
R960 B.n573 B.n571 163.367
R961 B.n569 B.n242 163.367
R962 B.n565 B.n563 163.367
R963 B.n561 B.n244 163.367
R964 B.n557 B.n555 163.367
R965 B.n553 B.n246 163.367
R966 B.n549 B.n547 163.367
R967 B.n545 B.n248 163.367
R968 B.n541 B.n539 163.367
R969 B.n537 B.n250 163.367
R970 B.n533 B.n531 163.367
R971 B.n529 B.n252 163.367
R972 B.n525 B.n523 163.367
R973 B.n521 B.n254 163.367
R974 B.n517 B.n515 163.367
R975 B.n513 B.n256 163.367
R976 B.n509 B.n507 163.367
R977 B.n505 B.n258 163.367
R978 B.n501 B.n499 163.367
R979 B.n497 B.n260 163.367
R980 B.n493 B.n491 163.367
R981 B.n489 B.n262 163.367
R982 B.n485 B.n483 163.367
R983 B.n481 B.n264 163.367
R984 B.n477 B.n475 163.367
R985 B.n473 B.n266 163.367
R986 B.n469 B.n467 163.367
R987 B.n465 B.n268 163.367
R988 B.n461 B.n459 163.367
R989 B.n456 B.n455 163.367
R990 B.n453 B.n274 163.367
R991 B.n449 B.n447 163.367
R992 B.n445 B.n276 163.367
R993 B.n441 B.n439 163.367
R994 B.n436 B.n435 163.367
R995 B.n433 B.n282 163.367
R996 B.n429 B.n427 163.367
R997 B.n425 B.n284 163.367
R998 B.n421 B.n419 163.367
R999 B.n417 B.n286 163.367
R1000 B.n413 B.n411 163.367
R1001 B.n409 B.n288 163.367
R1002 B.n405 B.n403 163.367
R1003 B.n401 B.n290 163.367
R1004 B.n397 B.n395 163.367
R1005 B.n393 B.n292 163.367
R1006 B.n389 B.n387 163.367
R1007 B.n385 B.n294 163.367
R1008 B.n381 B.n379 163.367
R1009 B.n377 B.n296 163.367
R1010 B.n373 B.n371 163.367
R1011 B.n369 B.n298 163.367
R1012 B.n365 B.n363 163.367
R1013 B.n361 B.n300 163.367
R1014 B.n357 B.n355 163.367
R1015 B.n353 B.n302 163.367
R1016 B.n349 B.n347 163.367
R1017 B.n345 B.n304 163.367
R1018 B.n341 B.n339 163.367
R1019 B.n337 B.n306 163.367
R1020 B.n333 B.n331 163.367
R1021 B.n329 B.n308 163.367
R1022 B.n325 B.n323 163.367
R1023 B.n321 B.n310 163.367
R1024 B.n317 B.n315 163.367
R1025 B.n313 B.n234 163.367
R1026 B.n590 B.n230 163.367
R1027 B.n598 B.n230 163.367
R1028 B.n598 B.n228 163.367
R1029 B.n602 B.n228 163.367
R1030 B.n602 B.n222 163.367
R1031 B.n610 B.n222 163.367
R1032 B.n610 B.n220 163.367
R1033 B.n614 B.n220 163.367
R1034 B.n614 B.n214 163.367
R1035 B.n622 B.n214 163.367
R1036 B.n622 B.n212 163.367
R1037 B.n626 B.n212 163.367
R1038 B.n626 B.n206 163.367
R1039 B.n634 B.n206 163.367
R1040 B.n634 B.n204 163.367
R1041 B.n638 B.n204 163.367
R1042 B.n638 B.n198 163.367
R1043 B.n646 B.n198 163.367
R1044 B.n646 B.n196 163.367
R1045 B.n650 B.n196 163.367
R1046 B.n650 B.n190 163.367
R1047 B.n659 B.n190 163.367
R1048 B.n659 B.n188 163.367
R1049 B.n663 B.n188 163.367
R1050 B.n663 B.n183 163.367
R1051 B.n671 B.n183 163.367
R1052 B.n671 B.n181 163.367
R1053 B.n675 B.n181 163.367
R1054 B.n675 B.n175 163.367
R1055 B.n683 B.n175 163.367
R1056 B.n683 B.n173 163.367
R1057 B.n687 B.n173 163.367
R1058 B.n687 B.n167 163.367
R1059 B.n696 B.n167 163.367
R1060 B.n696 B.n165 163.367
R1061 B.n700 B.n165 163.367
R1062 B.n700 B.n160 163.367
R1063 B.n709 B.n160 163.367
R1064 B.n709 B.n158 163.367
R1065 B.n713 B.n158 163.367
R1066 B.n713 B.n3 163.367
R1067 B.n1140 B.n3 163.367
R1068 B.n1136 B.n2 163.367
R1069 B.n1136 B.n1135 163.367
R1070 B.n1135 B.n9 163.367
R1071 B.n1131 B.n9 163.367
R1072 B.n1131 B.n11 163.367
R1073 B.n1127 B.n11 163.367
R1074 B.n1127 B.n16 163.367
R1075 B.n1123 B.n16 163.367
R1076 B.n1123 B.n18 163.367
R1077 B.n1119 B.n18 163.367
R1078 B.n1119 B.n24 163.367
R1079 B.n1115 B.n24 163.367
R1080 B.n1115 B.n26 163.367
R1081 B.n1111 B.n26 163.367
R1082 B.n1111 B.n31 163.367
R1083 B.n1107 B.n31 163.367
R1084 B.n1107 B.n33 163.367
R1085 B.n1103 B.n33 163.367
R1086 B.n1103 B.n37 163.367
R1087 B.n1099 B.n37 163.367
R1088 B.n1099 B.n39 163.367
R1089 B.n1095 B.n39 163.367
R1090 B.n1095 B.n45 163.367
R1091 B.n1091 B.n45 163.367
R1092 B.n1091 B.n47 163.367
R1093 B.n1087 B.n47 163.367
R1094 B.n1087 B.n52 163.367
R1095 B.n1083 B.n52 163.367
R1096 B.n1083 B.n54 163.367
R1097 B.n1079 B.n54 163.367
R1098 B.n1079 B.n59 163.367
R1099 B.n1075 B.n59 163.367
R1100 B.n1075 B.n61 163.367
R1101 B.n1071 B.n61 163.367
R1102 B.n1071 B.n66 163.367
R1103 B.n1067 B.n66 163.367
R1104 B.n1067 B.n68 163.367
R1105 B.n1063 B.n68 163.367
R1106 B.n1063 B.n73 163.367
R1107 B.n1059 B.n73 163.367
R1108 B.n1059 B.n75 163.367
R1109 B.n1055 B.n75 163.367
R1110 B.n121 B.t10 147.239
R1111 B.n277 B.t7 147.239
R1112 B.n113 B.t13 147.214
R1113 B.n269 B.t17 147.214
R1114 B.n114 B.n113 75.249
R1115 B.n122 B.n121 75.249
R1116 B.n278 B.n277 75.249
R1117 B.n270 B.n269 75.249
R1118 B.n122 B.t11 71.9914
R1119 B.n278 B.t6 71.9914
R1120 B.n114 B.t14 71.9646
R1121 B.n270 B.t16 71.9646
R1122 B.n1050 B.n80 71.676
R1123 B.n1049 B.n1048 71.676
R1124 B.n1042 B.n82 71.676
R1125 B.n1041 B.n1040 71.676
R1126 B.n1034 B.n84 71.676
R1127 B.n1033 B.n1032 71.676
R1128 B.n1026 B.n86 71.676
R1129 B.n1025 B.n1024 71.676
R1130 B.n1018 B.n88 71.676
R1131 B.n1017 B.n1016 71.676
R1132 B.n1010 B.n90 71.676
R1133 B.n1009 B.n1008 71.676
R1134 B.n1002 B.n92 71.676
R1135 B.n1001 B.n1000 71.676
R1136 B.n994 B.n94 71.676
R1137 B.n993 B.n992 71.676
R1138 B.n986 B.n96 71.676
R1139 B.n985 B.n984 71.676
R1140 B.n978 B.n98 71.676
R1141 B.n977 B.n976 71.676
R1142 B.n970 B.n100 71.676
R1143 B.n969 B.n968 71.676
R1144 B.n962 B.n102 71.676
R1145 B.n961 B.n960 71.676
R1146 B.n954 B.n104 71.676
R1147 B.n953 B.n952 71.676
R1148 B.n946 B.n106 71.676
R1149 B.n945 B.n944 71.676
R1150 B.n938 B.n108 71.676
R1151 B.n937 B.n936 71.676
R1152 B.n930 B.n110 71.676
R1153 B.n929 B.n928 71.676
R1154 B.n921 B.n112 71.676
R1155 B.n920 B.n919 71.676
R1156 B.n913 B.n116 71.676
R1157 B.n912 B.n911 71.676
R1158 B.n905 B.n118 71.676
R1159 B.n904 B.n903 71.676
R1160 B.n897 B.n120 71.676
R1161 B.n896 B.n895 71.676
R1162 B.n889 B.n125 71.676
R1163 B.n888 B.n887 71.676
R1164 B.n881 B.n127 71.676
R1165 B.n880 B.n879 71.676
R1166 B.n873 B.n129 71.676
R1167 B.n872 B.n871 71.676
R1168 B.n865 B.n131 71.676
R1169 B.n864 B.n863 71.676
R1170 B.n857 B.n133 71.676
R1171 B.n856 B.n855 71.676
R1172 B.n849 B.n135 71.676
R1173 B.n848 B.n847 71.676
R1174 B.n841 B.n137 71.676
R1175 B.n840 B.n839 71.676
R1176 B.n833 B.n139 71.676
R1177 B.n832 B.n831 71.676
R1178 B.n825 B.n141 71.676
R1179 B.n824 B.n823 71.676
R1180 B.n817 B.n143 71.676
R1181 B.n816 B.n815 71.676
R1182 B.n809 B.n145 71.676
R1183 B.n808 B.n807 71.676
R1184 B.n801 B.n147 71.676
R1185 B.n800 B.n799 71.676
R1186 B.n793 B.n149 71.676
R1187 B.n792 B.n791 71.676
R1188 B.n785 B.n151 71.676
R1189 B.n784 B.n783 71.676
R1190 B.n777 B.n153 71.676
R1191 B.n776 B.n775 71.676
R1192 B.n775 B.n774 71.676
R1193 B.n778 B.n777 71.676
R1194 B.n783 B.n782 71.676
R1195 B.n786 B.n785 71.676
R1196 B.n791 B.n790 71.676
R1197 B.n794 B.n793 71.676
R1198 B.n799 B.n798 71.676
R1199 B.n802 B.n801 71.676
R1200 B.n807 B.n806 71.676
R1201 B.n810 B.n809 71.676
R1202 B.n815 B.n814 71.676
R1203 B.n818 B.n817 71.676
R1204 B.n823 B.n822 71.676
R1205 B.n826 B.n825 71.676
R1206 B.n831 B.n830 71.676
R1207 B.n834 B.n833 71.676
R1208 B.n839 B.n838 71.676
R1209 B.n842 B.n841 71.676
R1210 B.n847 B.n846 71.676
R1211 B.n850 B.n849 71.676
R1212 B.n855 B.n854 71.676
R1213 B.n858 B.n857 71.676
R1214 B.n863 B.n862 71.676
R1215 B.n866 B.n865 71.676
R1216 B.n871 B.n870 71.676
R1217 B.n874 B.n873 71.676
R1218 B.n879 B.n878 71.676
R1219 B.n882 B.n881 71.676
R1220 B.n887 B.n886 71.676
R1221 B.n890 B.n889 71.676
R1222 B.n895 B.n894 71.676
R1223 B.n898 B.n897 71.676
R1224 B.n903 B.n902 71.676
R1225 B.n906 B.n905 71.676
R1226 B.n911 B.n910 71.676
R1227 B.n914 B.n913 71.676
R1228 B.n919 B.n918 71.676
R1229 B.n922 B.n921 71.676
R1230 B.n928 B.n927 71.676
R1231 B.n931 B.n930 71.676
R1232 B.n936 B.n935 71.676
R1233 B.n939 B.n938 71.676
R1234 B.n944 B.n943 71.676
R1235 B.n947 B.n946 71.676
R1236 B.n952 B.n951 71.676
R1237 B.n955 B.n954 71.676
R1238 B.n960 B.n959 71.676
R1239 B.n963 B.n962 71.676
R1240 B.n968 B.n967 71.676
R1241 B.n971 B.n970 71.676
R1242 B.n976 B.n975 71.676
R1243 B.n979 B.n978 71.676
R1244 B.n984 B.n983 71.676
R1245 B.n987 B.n986 71.676
R1246 B.n992 B.n991 71.676
R1247 B.n995 B.n994 71.676
R1248 B.n1000 B.n999 71.676
R1249 B.n1003 B.n1002 71.676
R1250 B.n1008 B.n1007 71.676
R1251 B.n1011 B.n1010 71.676
R1252 B.n1016 B.n1015 71.676
R1253 B.n1019 B.n1018 71.676
R1254 B.n1024 B.n1023 71.676
R1255 B.n1027 B.n1026 71.676
R1256 B.n1032 B.n1031 71.676
R1257 B.n1035 B.n1034 71.676
R1258 B.n1040 B.n1039 71.676
R1259 B.n1043 B.n1042 71.676
R1260 B.n1048 B.n1047 71.676
R1261 B.n1051 B.n1050 71.676
R1262 B.n585 B.n236 71.676
R1263 B.n583 B.n238 71.676
R1264 B.n579 B.n578 71.676
R1265 B.n572 B.n240 71.676
R1266 B.n571 B.n570 71.676
R1267 B.n564 B.n242 71.676
R1268 B.n563 B.n562 71.676
R1269 B.n556 B.n244 71.676
R1270 B.n555 B.n554 71.676
R1271 B.n548 B.n246 71.676
R1272 B.n547 B.n546 71.676
R1273 B.n540 B.n248 71.676
R1274 B.n539 B.n538 71.676
R1275 B.n532 B.n250 71.676
R1276 B.n531 B.n530 71.676
R1277 B.n524 B.n252 71.676
R1278 B.n523 B.n522 71.676
R1279 B.n516 B.n254 71.676
R1280 B.n515 B.n514 71.676
R1281 B.n508 B.n256 71.676
R1282 B.n507 B.n506 71.676
R1283 B.n500 B.n258 71.676
R1284 B.n499 B.n498 71.676
R1285 B.n492 B.n260 71.676
R1286 B.n491 B.n490 71.676
R1287 B.n484 B.n262 71.676
R1288 B.n483 B.n482 71.676
R1289 B.n476 B.n264 71.676
R1290 B.n475 B.n474 71.676
R1291 B.n468 B.n266 71.676
R1292 B.n467 B.n466 71.676
R1293 B.n460 B.n268 71.676
R1294 B.n459 B.n272 71.676
R1295 B.n455 B.n454 71.676
R1296 B.n448 B.n274 71.676
R1297 B.n447 B.n446 71.676
R1298 B.n440 B.n276 71.676
R1299 B.n439 B.n280 71.676
R1300 B.n435 B.n434 71.676
R1301 B.n428 B.n282 71.676
R1302 B.n427 B.n426 71.676
R1303 B.n420 B.n284 71.676
R1304 B.n419 B.n418 71.676
R1305 B.n412 B.n286 71.676
R1306 B.n411 B.n410 71.676
R1307 B.n404 B.n288 71.676
R1308 B.n403 B.n402 71.676
R1309 B.n396 B.n290 71.676
R1310 B.n395 B.n394 71.676
R1311 B.n388 B.n292 71.676
R1312 B.n387 B.n386 71.676
R1313 B.n380 B.n294 71.676
R1314 B.n379 B.n378 71.676
R1315 B.n372 B.n296 71.676
R1316 B.n371 B.n370 71.676
R1317 B.n364 B.n298 71.676
R1318 B.n363 B.n362 71.676
R1319 B.n356 B.n300 71.676
R1320 B.n355 B.n354 71.676
R1321 B.n348 B.n302 71.676
R1322 B.n347 B.n346 71.676
R1323 B.n340 B.n304 71.676
R1324 B.n339 B.n338 71.676
R1325 B.n332 B.n306 71.676
R1326 B.n331 B.n330 71.676
R1327 B.n324 B.n308 71.676
R1328 B.n323 B.n322 71.676
R1329 B.n316 B.n310 71.676
R1330 B.n315 B.n314 71.676
R1331 B.n586 B.n585 71.676
R1332 B.n580 B.n238 71.676
R1333 B.n578 B.n577 71.676
R1334 B.n573 B.n572 71.676
R1335 B.n570 B.n569 71.676
R1336 B.n565 B.n564 71.676
R1337 B.n562 B.n561 71.676
R1338 B.n557 B.n556 71.676
R1339 B.n554 B.n553 71.676
R1340 B.n549 B.n548 71.676
R1341 B.n546 B.n545 71.676
R1342 B.n541 B.n540 71.676
R1343 B.n538 B.n537 71.676
R1344 B.n533 B.n532 71.676
R1345 B.n530 B.n529 71.676
R1346 B.n525 B.n524 71.676
R1347 B.n522 B.n521 71.676
R1348 B.n517 B.n516 71.676
R1349 B.n514 B.n513 71.676
R1350 B.n509 B.n508 71.676
R1351 B.n506 B.n505 71.676
R1352 B.n501 B.n500 71.676
R1353 B.n498 B.n497 71.676
R1354 B.n493 B.n492 71.676
R1355 B.n490 B.n489 71.676
R1356 B.n485 B.n484 71.676
R1357 B.n482 B.n481 71.676
R1358 B.n477 B.n476 71.676
R1359 B.n474 B.n473 71.676
R1360 B.n469 B.n468 71.676
R1361 B.n466 B.n465 71.676
R1362 B.n461 B.n460 71.676
R1363 B.n456 B.n272 71.676
R1364 B.n454 B.n453 71.676
R1365 B.n449 B.n448 71.676
R1366 B.n446 B.n445 71.676
R1367 B.n441 B.n440 71.676
R1368 B.n436 B.n280 71.676
R1369 B.n434 B.n433 71.676
R1370 B.n429 B.n428 71.676
R1371 B.n426 B.n425 71.676
R1372 B.n421 B.n420 71.676
R1373 B.n418 B.n417 71.676
R1374 B.n413 B.n412 71.676
R1375 B.n410 B.n409 71.676
R1376 B.n405 B.n404 71.676
R1377 B.n402 B.n401 71.676
R1378 B.n397 B.n396 71.676
R1379 B.n394 B.n393 71.676
R1380 B.n389 B.n388 71.676
R1381 B.n386 B.n385 71.676
R1382 B.n381 B.n380 71.676
R1383 B.n378 B.n377 71.676
R1384 B.n373 B.n372 71.676
R1385 B.n370 B.n369 71.676
R1386 B.n365 B.n364 71.676
R1387 B.n362 B.n361 71.676
R1388 B.n357 B.n356 71.676
R1389 B.n354 B.n353 71.676
R1390 B.n349 B.n348 71.676
R1391 B.n346 B.n345 71.676
R1392 B.n341 B.n340 71.676
R1393 B.n338 B.n337 71.676
R1394 B.n333 B.n332 71.676
R1395 B.n330 B.n329 71.676
R1396 B.n325 B.n324 71.676
R1397 B.n322 B.n321 71.676
R1398 B.n317 B.n316 71.676
R1399 B.n314 B.n313 71.676
R1400 B.n1141 B.n1140 71.676
R1401 B.n1141 B.n2 71.676
R1402 B.n924 B.n114 59.5399
R1403 B.n123 B.n122 59.5399
R1404 B.n279 B.n278 59.5399
R1405 B.n271 B.n270 59.5399
R1406 B.n591 B.n235 49.238
R1407 B.n1056 B.n79 49.238
R1408 B.n591 B.n231 29.6301
R1409 B.n597 B.n231 29.6301
R1410 B.n597 B.n227 29.6301
R1411 B.n603 B.n227 29.6301
R1412 B.n603 B.n223 29.6301
R1413 B.n609 B.n223 29.6301
R1414 B.n609 B.n218 29.6301
R1415 B.n615 B.n218 29.6301
R1416 B.n615 B.n219 29.6301
R1417 B.n621 B.n211 29.6301
R1418 B.n627 B.n211 29.6301
R1419 B.n627 B.n207 29.6301
R1420 B.n633 B.n207 29.6301
R1421 B.n633 B.n203 29.6301
R1422 B.n639 B.n203 29.6301
R1423 B.n639 B.n199 29.6301
R1424 B.n645 B.n199 29.6301
R1425 B.n645 B.n195 29.6301
R1426 B.n651 B.n195 29.6301
R1427 B.n651 B.n191 29.6301
R1428 B.n658 B.n191 29.6301
R1429 B.n658 B.n657 29.6301
R1430 B.n664 B.n184 29.6301
R1431 B.n670 B.n184 29.6301
R1432 B.n670 B.n180 29.6301
R1433 B.n676 B.n180 29.6301
R1434 B.n676 B.n176 29.6301
R1435 B.n682 B.n176 29.6301
R1436 B.n682 B.n172 29.6301
R1437 B.n688 B.n172 29.6301
R1438 B.n688 B.n168 29.6301
R1439 B.n695 B.n168 29.6301
R1440 B.n695 B.n694 29.6301
R1441 B.n701 B.n161 29.6301
R1442 B.n708 B.n161 29.6301
R1443 B.n708 B.n157 29.6301
R1444 B.n714 B.n157 29.6301
R1445 B.n714 B.n4 29.6301
R1446 B.n1139 B.n4 29.6301
R1447 B.n1139 B.n1138 29.6301
R1448 B.n1138 B.n1137 29.6301
R1449 B.n1137 B.n8 29.6301
R1450 B.n12 B.n8 29.6301
R1451 B.n1130 B.n12 29.6301
R1452 B.n1130 B.n1129 29.6301
R1453 B.n1129 B.n1128 29.6301
R1454 B.n1122 B.n19 29.6301
R1455 B.n1122 B.n1121 29.6301
R1456 B.n1121 B.n1120 29.6301
R1457 B.n1120 B.n23 29.6301
R1458 B.n1114 B.n23 29.6301
R1459 B.n1114 B.n1113 29.6301
R1460 B.n1113 B.n1112 29.6301
R1461 B.n1112 B.n30 29.6301
R1462 B.n1106 B.n30 29.6301
R1463 B.n1106 B.n1105 29.6301
R1464 B.n1105 B.n1104 29.6301
R1465 B.n1098 B.n40 29.6301
R1466 B.n1098 B.n1097 29.6301
R1467 B.n1097 B.n1096 29.6301
R1468 B.n1096 B.n44 29.6301
R1469 B.n1090 B.n44 29.6301
R1470 B.n1090 B.n1089 29.6301
R1471 B.n1089 B.n1088 29.6301
R1472 B.n1088 B.n51 29.6301
R1473 B.n1082 B.n51 29.6301
R1474 B.n1082 B.n1081 29.6301
R1475 B.n1081 B.n1080 29.6301
R1476 B.n1080 B.n58 29.6301
R1477 B.n1074 B.n58 29.6301
R1478 B.n1073 B.n1072 29.6301
R1479 B.n1072 B.n65 29.6301
R1480 B.n1066 B.n65 29.6301
R1481 B.n1066 B.n1065 29.6301
R1482 B.n1065 B.n1064 29.6301
R1483 B.n1064 B.n72 29.6301
R1484 B.n1058 B.n72 29.6301
R1485 B.n1058 B.n1057 29.6301
R1486 B.n1057 B.n1056 29.6301
R1487 B.n589 B.n588 29.1907
R1488 B.n593 B.n233 29.1907
R1489 B.n773 B.n772 29.1907
R1490 B.n1054 B.n1053 29.1907
R1491 B.n621 B.t5 24.8371
R1492 B.n1074 B.t9 24.8371
R1493 B.n701 B.t0 23.9656
R1494 B.n1128 B.t3 23.9656
R1495 B.n657 B.t2 23.0942
R1496 B.n40 B.t1 23.0942
R1497 B B.n1142 18.0485
R1498 B.n589 B.n229 10.6151
R1499 B.n599 B.n229 10.6151
R1500 B.n600 B.n599 10.6151
R1501 B.n601 B.n600 10.6151
R1502 B.n601 B.n221 10.6151
R1503 B.n611 B.n221 10.6151
R1504 B.n612 B.n611 10.6151
R1505 B.n613 B.n612 10.6151
R1506 B.n613 B.n213 10.6151
R1507 B.n623 B.n213 10.6151
R1508 B.n624 B.n623 10.6151
R1509 B.n625 B.n624 10.6151
R1510 B.n625 B.n205 10.6151
R1511 B.n635 B.n205 10.6151
R1512 B.n636 B.n635 10.6151
R1513 B.n637 B.n636 10.6151
R1514 B.n637 B.n197 10.6151
R1515 B.n647 B.n197 10.6151
R1516 B.n648 B.n647 10.6151
R1517 B.n649 B.n648 10.6151
R1518 B.n649 B.n189 10.6151
R1519 B.n660 B.n189 10.6151
R1520 B.n661 B.n660 10.6151
R1521 B.n662 B.n661 10.6151
R1522 B.n662 B.n182 10.6151
R1523 B.n672 B.n182 10.6151
R1524 B.n673 B.n672 10.6151
R1525 B.n674 B.n673 10.6151
R1526 B.n674 B.n174 10.6151
R1527 B.n684 B.n174 10.6151
R1528 B.n685 B.n684 10.6151
R1529 B.n686 B.n685 10.6151
R1530 B.n686 B.n166 10.6151
R1531 B.n697 B.n166 10.6151
R1532 B.n698 B.n697 10.6151
R1533 B.n699 B.n698 10.6151
R1534 B.n699 B.n159 10.6151
R1535 B.n710 B.n159 10.6151
R1536 B.n711 B.n710 10.6151
R1537 B.n712 B.n711 10.6151
R1538 B.n712 B.n0 10.6151
R1539 B.n588 B.n587 10.6151
R1540 B.n587 B.n237 10.6151
R1541 B.n582 B.n237 10.6151
R1542 B.n582 B.n581 10.6151
R1543 B.n581 B.n239 10.6151
R1544 B.n576 B.n239 10.6151
R1545 B.n576 B.n575 10.6151
R1546 B.n575 B.n574 10.6151
R1547 B.n574 B.n241 10.6151
R1548 B.n568 B.n241 10.6151
R1549 B.n568 B.n567 10.6151
R1550 B.n567 B.n566 10.6151
R1551 B.n566 B.n243 10.6151
R1552 B.n560 B.n243 10.6151
R1553 B.n560 B.n559 10.6151
R1554 B.n559 B.n558 10.6151
R1555 B.n558 B.n245 10.6151
R1556 B.n552 B.n245 10.6151
R1557 B.n552 B.n551 10.6151
R1558 B.n551 B.n550 10.6151
R1559 B.n550 B.n247 10.6151
R1560 B.n544 B.n247 10.6151
R1561 B.n544 B.n543 10.6151
R1562 B.n543 B.n542 10.6151
R1563 B.n542 B.n249 10.6151
R1564 B.n536 B.n249 10.6151
R1565 B.n536 B.n535 10.6151
R1566 B.n535 B.n534 10.6151
R1567 B.n534 B.n251 10.6151
R1568 B.n528 B.n251 10.6151
R1569 B.n528 B.n527 10.6151
R1570 B.n527 B.n526 10.6151
R1571 B.n526 B.n253 10.6151
R1572 B.n520 B.n253 10.6151
R1573 B.n520 B.n519 10.6151
R1574 B.n519 B.n518 10.6151
R1575 B.n518 B.n255 10.6151
R1576 B.n512 B.n255 10.6151
R1577 B.n512 B.n511 10.6151
R1578 B.n511 B.n510 10.6151
R1579 B.n510 B.n257 10.6151
R1580 B.n504 B.n257 10.6151
R1581 B.n504 B.n503 10.6151
R1582 B.n503 B.n502 10.6151
R1583 B.n502 B.n259 10.6151
R1584 B.n496 B.n259 10.6151
R1585 B.n496 B.n495 10.6151
R1586 B.n495 B.n494 10.6151
R1587 B.n494 B.n261 10.6151
R1588 B.n488 B.n261 10.6151
R1589 B.n488 B.n487 10.6151
R1590 B.n487 B.n486 10.6151
R1591 B.n486 B.n263 10.6151
R1592 B.n480 B.n263 10.6151
R1593 B.n480 B.n479 10.6151
R1594 B.n479 B.n478 10.6151
R1595 B.n478 B.n265 10.6151
R1596 B.n472 B.n265 10.6151
R1597 B.n472 B.n471 10.6151
R1598 B.n471 B.n470 10.6151
R1599 B.n470 B.n267 10.6151
R1600 B.n464 B.n267 10.6151
R1601 B.n464 B.n463 10.6151
R1602 B.n463 B.n462 10.6151
R1603 B.n458 B.n457 10.6151
R1604 B.n457 B.n273 10.6151
R1605 B.n452 B.n273 10.6151
R1606 B.n452 B.n451 10.6151
R1607 B.n451 B.n450 10.6151
R1608 B.n450 B.n275 10.6151
R1609 B.n444 B.n275 10.6151
R1610 B.n444 B.n443 10.6151
R1611 B.n443 B.n442 10.6151
R1612 B.n438 B.n437 10.6151
R1613 B.n437 B.n281 10.6151
R1614 B.n432 B.n281 10.6151
R1615 B.n432 B.n431 10.6151
R1616 B.n431 B.n430 10.6151
R1617 B.n430 B.n283 10.6151
R1618 B.n424 B.n283 10.6151
R1619 B.n424 B.n423 10.6151
R1620 B.n423 B.n422 10.6151
R1621 B.n422 B.n285 10.6151
R1622 B.n416 B.n285 10.6151
R1623 B.n416 B.n415 10.6151
R1624 B.n415 B.n414 10.6151
R1625 B.n414 B.n287 10.6151
R1626 B.n408 B.n287 10.6151
R1627 B.n408 B.n407 10.6151
R1628 B.n407 B.n406 10.6151
R1629 B.n406 B.n289 10.6151
R1630 B.n400 B.n289 10.6151
R1631 B.n400 B.n399 10.6151
R1632 B.n399 B.n398 10.6151
R1633 B.n398 B.n291 10.6151
R1634 B.n392 B.n291 10.6151
R1635 B.n392 B.n391 10.6151
R1636 B.n391 B.n390 10.6151
R1637 B.n390 B.n293 10.6151
R1638 B.n384 B.n293 10.6151
R1639 B.n384 B.n383 10.6151
R1640 B.n383 B.n382 10.6151
R1641 B.n382 B.n295 10.6151
R1642 B.n376 B.n295 10.6151
R1643 B.n376 B.n375 10.6151
R1644 B.n375 B.n374 10.6151
R1645 B.n374 B.n297 10.6151
R1646 B.n368 B.n297 10.6151
R1647 B.n368 B.n367 10.6151
R1648 B.n367 B.n366 10.6151
R1649 B.n366 B.n299 10.6151
R1650 B.n360 B.n299 10.6151
R1651 B.n360 B.n359 10.6151
R1652 B.n359 B.n358 10.6151
R1653 B.n358 B.n301 10.6151
R1654 B.n352 B.n301 10.6151
R1655 B.n352 B.n351 10.6151
R1656 B.n351 B.n350 10.6151
R1657 B.n350 B.n303 10.6151
R1658 B.n344 B.n303 10.6151
R1659 B.n344 B.n343 10.6151
R1660 B.n343 B.n342 10.6151
R1661 B.n342 B.n305 10.6151
R1662 B.n336 B.n305 10.6151
R1663 B.n336 B.n335 10.6151
R1664 B.n335 B.n334 10.6151
R1665 B.n334 B.n307 10.6151
R1666 B.n328 B.n307 10.6151
R1667 B.n328 B.n327 10.6151
R1668 B.n327 B.n326 10.6151
R1669 B.n326 B.n309 10.6151
R1670 B.n320 B.n309 10.6151
R1671 B.n320 B.n319 10.6151
R1672 B.n319 B.n318 10.6151
R1673 B.n318 B.n311 10.6151
R1674 B.n312 B.n311 10.6151
R1675 B.n312 B.n233 10.6151
R1676 B.n594 B.n593 10.6151
R1677 B.n595 B.n594 10.6151
R1678 B.n595 B.n225 10.6151
R1679 B.n605 B.n225 10.6151
R1680 B.n606 B.n605 10.6151
R1681 B.n607 B.n606 10.6151
R1682 B.n607 B.n216 10.6151
R1683 B.n617 B.n216 10.6151
R1684 B.n618 B.n617 10.6151
R1685 B.n619 B.n618 10.6151
R1686 B.n619 B.n209 10.6151
R1687 B.n629 B.n209 10.6151
R1688 B.n630 B.n629 10.6151
R1689 B.n631 B.n630 10.6151
R1690 B.n631 B.n201 10.6151
R1691 B.n641 B.n201 10.6151
R1692 B.n642 B.n641 10.6151
R1693 B.n643 B.n642 10.6151
R1694 B.n643 B.n193 10.6151
R1695 B.n653 B.n193 10.6151
R1696 B.n654 B.n653 10.6151
R1697 B.n655 B.n654 10.6151
R1698 B.n655 B.n186 10.6151
R1699 B.n666 B.n186 10.6151
R1700 B.n667 B.n666 10.6151
R1701 B.n668 B.n667 10.6151
R1702 B.n668 B.n178 10.6151
R1703 B.n678 B.n178 10.6151
R1704 B.n679 B.n678 10.6151
R1705 B.n680 B.n679 10.6151
R1706 B.n680 B.n170 10.6151
R1707 B.n690 B.n170 10.6151
R1708 B.n691 B.n690 10.6151
R1709 B.n692 B.n691 10.6151
R1710 B.n692 B.n163 10.6151
R1711 B.n703 B.n163 10.6151
R1712 B.n704 B.n703 10.6151
R1713 B.n706 B.n704 10.6151
R1714 B.n706 B.n705 10.6151
R1715 B.n705 B.n155 10.6151
R1716 B.n717 B.n155 10.6151
R1717 B.n718 B.n717 10.6151
R1718 B.n719 B.n718 10.6151
R1719 B.n720 B.n719 10.6151
R1720 B.n721 B.n720 10.6151
R1721 B.n724 B.n721 10.6151
R1722 B.n725 B.n724 10.6151
R1723 B.n726 B.n725 10.6151
R1724 B.n727 B.n726 10.6151
R1725 B.n729 B.n727 10.6151
R1726 B.n730 B.n729 10.6151
R1727 B.n731 B.n730 10.6151
R1728 B.n732 B.n731 10.6151
R1729 B.n734 B.n732 10.6151
R1730 B.n735 B.n734 10.6151
R1731 B.n736 B.n735 10.6151
R1732 B.n737 B.n736 10.6151
R1733 B.n739 B.n737 10.6151
R1734 B.n740 B.n739 10.6151
R1735 B.n741 B.n740 10.6151
R1736 B.n742 B.n741 10.6151
R1737 B.n744 B.n742 10.6151
R1738 B.n745 B.n744 10.6151
R1739 B.n746 B.n745 10.6151
R1740 B.n747 B.n746 10.6151
R1741 B.n749 B.n747 10.6151
R1742 B.n750 B.n749 10.6151
R1743 B.n751 B.n750 10.6151
R1744 B.n752 B.n751 10.6151
R1745 B.n754 B.n752 10.6151
R1746 B.n755 B.n754 10.6151
R1747 B.n756 B.n755 10.6151
R1748 B.n757 B.n756 10.6151
R1749 B.n759 B.n757 10.6151
R1750 B.n760 B.n759 10.6151
R1751 B.n761 B.n760 10.6151
R1752 B.n762 B.n761 10.6151
R1753 B.n764 B.n762 10.6151
R1754 B.n765 B.n764 10.6151
R1755 B.n766 B.n765 10.6151
R1756 B.n767 B.n766 10.6151
R1757 B.n769 B.n767 10.6151
R1758 B.n770 B.n769 10.6151
R1759 B.n771 B.n770 10.6151
R1760 B.n772 B.n771 10.6151
R1761 B.n1134 B.n1 10.6151
R1762 B.n1134 B.n1133 10.6151
R1763 B.n1133 B.n1132 10.6151
R1764 B.n1132 B.n10 10.6151
R1765 B.n1126 B.n10 10.6151
R1766 B.n1126 B.n1125 10.6151
R1767 B.n1125 B.n1124 10.6151
R1768 B.n1124 B.n17 10.6151
R1769 B.n1118 B.n17 10.6151
R1770 B.n1118 B.n1117 10.6151
R1771 B.n1117 B.n1116 10.6151
R1772 B.n1116 B.n25 10.6151
R1773 B.n1110 B.n25 10.6151
R1774 B.n1110 B.n1109 10.6151
R1775 B.n1109 B.n1108 10.6151
R1776 B.n1108 B.n32 10.6151
R1777 B.n1102 B.n32 10.6151
R1778 B.n1102 B.n1101 10.6151
R1779 B.n1101 B.n1100 10.6151
R1780 B.n1100 B.n38 10.6151
R1781 B.n1094 B.n38 10.6151
R1782 B.n1094 B.n1093 10.6151
R1783 B.n1093 B.n1092 10.6151
R1784 B.n1092 B.n46 10.6151
R1785 B.n1086 B.n46 10.6151
R1786 B.n1086 B.n1085 10.6151
R1787 B.n1085 B.n1084 10.6151
R1788 B.n1084 B.n53 10.6151
R1789 B.n1078 B.n53 10.6151
R1790 B.n1078 B.n1077 10.6151
R1791 B.n1077 B.n1076 10.6151
R1792 B.n1076 B.n60 10.6151
R1793 B.n1070 B.n60 10.6151
R1794 B.n1070 B.n1069 10.6151
R1795 B.n1069 B.n1068 10.6151
R1796 B.n1068 B.n67 10.6151
R1797 B.n1062 B.n67 10.6151
R1798 B.n1062 B.n1061 10.6151
R1799 B.n1061 B.n1060 10.6151
R1800 B.n1060 B.n74 10.6151
R1801 B.n1054 B.n74 10.6151
R1802 B.n1053 B.n1052 10.6151
R1803 B.n1052 B.n81 10.6151
R1804 B.n1046 B.n81 10.6151
R1805 B.n1046 B.n1045 10.6151
R1806 B.n1045 B.n1044 10.6151
R1807 B.n1044 B.n83 10.6151
R1808 B.n1038 B.n83 10.6151
R1809 B.n1038 B.n1037 10.6151
R1810 B.n1037 B.n1036 10.6151
R1811 B.n1036 B.n85 10.6151
R1812 B.n1030 B.n85 10.6151
R1813 B.n1030 B.n1029 10.6151
R1814 B.n1029 B.n1028 10.6151
R1815 B.n1028 B.n87 10.6151
R1816 B.n1022 B.n87 10.6151
R1817 B.n1022 B.n1021 10.6151
R1818 B.n1021 B.n1020 10.6151
R1819 B.n1020 B.n89 10.6151
R1820 B.n1014 B.n89 10.6151
R1821 B.n1014 B.n1013 10.6151
R1822 B.n1013 B.n1012 10.6151
R1823 B.n1012 B.n91 10.6151
R1824 B.n1006 B.n91 10.6151
R1825 B.n1006 B.n1005 10.6151
R1826 B.n1005 B.n1004 10.6151
R1827 B.n1004 B.n93 10.6151
R1828 B.n998 B.n93 10.6151
R1829 B.n998 B.n997 10.6151
R1830 B.n997 B.n996 10.6151
R1831 B.n996 B.n95 10.6151
R1832 B.n990 B.n95 10.6151
R1833 B.n990 B.n989 10.6151
R1834 B.n989 B.n988 10.6151
R1835 B.n988 B.n97 10.6151
R1836 B.n982 B.n97 10.6151
R1837 B.n982 B.n981 10.6151
R1838 B.n981 B.n980 10.6151
R1839 B.n980 B.n99 10.6151
R1840 B.n974 B.n99 10.6151
R1841 B.n974 B.n973 10.6151
R1842 B.n973 B.n972 10.6151
R1843 B.n972 B.n101 10.6151
R1844 B.n966 B.n101 10.6151
R1845 B.n966 B.n965 10.6151
R1846 B.n965 B.n964 10.6151
R1847 B.n964 B.n103 10.6151
R1848 B.n958 B.n103 10.6151
R1849 B.n958 B.n957 10.6151
R1850 B.n957 B.n956 10.6151
R1851 B.n956 B.n105 10.6151
R1852 B.n950 B.n105 10.6151
R1853 B.n950 B.n949 10.6151
R1854 B.n949 B.n948 10.6151
R1855 B.n948 B.n107 10.6151
R1856 B.n942 B.n107 10.6151
R1857 B.n942 B.n941 10.6151
R1858 B.n941 B.n940 10.6151
R1859 B.n940 B.n109 10.6151
R1860 B.n934 B.n109 10.6151
R1861 B.n934 B.n933 10.6151
R1862 B.n933 B.n932 10.6151
R1863 B.n932 B.n111 10.6151
R1864 B.n926 B.n111 10.6151
R1865 B.n926 B.n925 10.6151
R1866 B.n923 B.n115 10.6151
R1867 B.n917 B.n115 10.6151
R1868 B.n917 B.n916 10.6151
R1869 B.n916 B.n915 10.6151
R1870 B.n915 B.n117 10.6151
R1871 B.n909 B.n117 10.6151
R1872 B.n909 B.n908 10.6151
R1873 B.n908 B.n907 10.6151
R1874 B.n907 B.n119 10.6151
R1875 B.n901 B.n900 10.6151
R1876 B.n900 B.n899 10.6151
R1877 B.n899 B.n124 10.6151
R1878 B.n893 B.n124 10.6151
R1879 B.n893 B.n892 10.6151
R1880 B.n892 B.n891 10.6151
R1881 B.n891 B.n126 10.6151
R1882 B.n885 B.n126 10.6151
R1883 B.n885 B.n884 10.6151
R1884 B.n884 B.n883 10.6151
R1885 B.n883 B.n128 10.6151
R1886 B.n877 B.n128 10.6151
R1887 B.n877 B.n876 10.6151
R1888 B.n876 B.n875 10.6151
R1889 B.n875 B.n130 10.6151
R1890 B.n869 B.n130 10.6151
R1891 B.n869 B.n868 10.6151
R1892 B.n868 B.n867 10.6151
R1893 B.n867 B.n132 10.6151
R1894 B.n861 B.n132 10.6151
R1895 B.n861 B.n860 10.6151
R1896 B.n860 B.n859 10.6151
R1897 B.n859 B.n134 10.6151
R1898 B.n853 B.n134 10.6151
R1899 B.n853 B.n852 10.6151
R1900 B.n852 B.n851 10.6151
R1901 B.n851 B.n136 10.6151
R1902 B.n845 B.n136 10.6151
R1903 B.n845 B.n844 10.6151
R1904 B.n844 B.n843 10.6151
R1905 B.n843 B.n138 10.6151
R1906 B.n837 B.n138 10.6151
R1907 B.n837 B.n836 10.6151
R1908 B.n836 B.n835 10.6151
R1909 B.n835 B.n140 10.6151
R1910 B.n829 B.n140 10.6151
R1911 B.n829 B.n828 10.6151
R1912 B.n828 B.n827 10.6151
R1913 B.n827 B.n142 10.6151
R1914 B.n821 B.n142 10.6151
R1915 B.n821 B.n820 10.6151
R1916 B.n820 B.n819 10.6151
R1917 B.n819 B.n144 10.6151
R1918 B.n813 B.n144 10.6151
R1919 B.n813 B.n812 10.6151
R1920 B.n812 B.n811 10.6151
R1921 B.n811 B.n146 10.6151
R1922 B.n805 B.n146 10.6151
R1923 B.n805 B.n804 10.6151
R1924 B.n804 B.n803 10.6151
R1925 B.n803 B.n148 10.6151
R1926 B.n797 B.n148 10.6151
R1927 B.n797 B.n796 10.6151
R1928 B.n796 B.n795 10.6151
R1929 B.n795 B.n150 10.6151
R1930 B.n789 B.n150 10.6151
R1931 B.n789 B.n788 10.6151
R1932 B.n788 B.n787 10.6151
R1933 B.n787 B.n152 10.6151
R1934 B.n781 B.n152 10.6151
R1935 B.n781 B.n780 10.6151
R1936 B.n780 B.n779 10.6151
R1937 B.n779 B.n154 10.6151
R1938 B.n773 B.n154 10.6151
R1939 B.n462 B.n271 9.36635
R1940 B.n438 B.n279 9.36635
R1941 B.n925 B.n924 9.36635
R1942 B.n901 B.n123 9.36635
R1943 B.n1142 B.n0 8.11757
R1944 B.n1142 B.n1 8.11757
R1945 B.n664 B.t2 6.53645
R1946 B.n1104 B.t1 6.53645
R1947 B.n694 B.t0 5.66499
R1948 B.n19 B.t3 5.66499
R1949 B.n219 B.t5 4.79353
R1950 B.t9 B.n1073 4.79353
R1951 B.n458 B.n271 1.24928
R1952 B.n442 B.n279 1.24928
R1953 B.n924 B.n923 1.24928
R1954 B.n123 B.n119 1.24928
R1955 VP.n5 VP.t0 170.238
R1956 VP.n5 VP.t2 169.006
R1957 VP.n19 VP.n18 161.3
R1958 VP.n17 VP.n1 161.3
R1959 VP.n16 VP.n15 161.3
R1960 VP.n14 VP.n2 161.3
R1961 VP.n13 VP.n12 161.3
R1962 VP.n11 VP.n3 161.3
R1963 VP.n10 VP.n9 161.3
R1964 VP.n8 VP.n4 161.3
R1965 VP.n6 VP.t1 135.571
R1966 VP.n0 VP.t3 135.571
R1967 VP.n7 VP.n6 80.7699
R1968 VP.n20 VP.n0 80.7699
R1969 VP.n7 VP.n5 57.4729
R1970 VP.n12 VP.n2 56.5193
R1971 VP.n10 VP.n4 24.4675
R1972 VP.n11 VP.n10 24.4675
R1973 VP.n12 VP.n11 24.4675
R1974 VP.n16 VP.n2 24.4675
R1975 VP.n17 VP.n16 24.4675
R1976 VP.n18 VP.n17 24.4675
R1977 VP.n6 VP.n4 9.29796
R1978 VP.n18 VP.n0 9.29796
R1979 VP.n8 VP.n7 0.354971
R1980 VP.n20 VP.n19 0.354971
R1981 VP VP.n20 0.26696
R1982 VP.n9 VP.n8 0.189894
R1983 VP.n9 VP.n3 0.189894
R1984 VP.n13 VP.n3 0.189894
R1985 VP.n14 VP.n13 0.189894
R1986 VP.n15 VP.n14 0.189894
R1987 VP.n15 VP.n1 0.189894
R1988 VP.n19 VP.n1 0.189894
R1989 VDD1 VDD1.n1 110.727
R1990 VDD1 VDD1.n0 59.2948
R1991 VDD1.n0 VDD1.t3 0.991987
R1992 VDD1.n0 VDD1.t1 0.991987
R1993 VDD1.n1 VDD1.t2 0.991987
R1994 VDD1.n1 VDD1.t0 0.991987
C0 VTAIL VP 7.77432f
C1 VDD1 VN 0.15001f
C2 VDD1 VDD2 1.25461f
C3 VDD1 VP 8.38517f
C4 VTAIL VDD1 7.35342f
C5 VDD2 VN 8.08125f
C6 VP VN 8.35193f
C7 VDD2 VP 0.454907f
C8 VTAIL VN 7.76022f
C9 VTAIL VDD2 7.414f
C10 VDD2 B 4.928629f
C11 VDD1 B 10.20035f
C12 VTAIL B 15.443799f
C13 VN B 13.16512f
C14 VP B 11.494373f
C15 VDD1.t3 B 0.424975f
C16 VDD1.t1 B 0.424975f
C17 VDD1.n0 B 3.88462f
C18 VDD1.t2 B 0.424975f
C19 VDD1.t0 B 0.424975f
C20 VDD1.n1 B 4.97671f
C21 VP.t3 B 3.83592f
C22 VP.n0 B 1.39436f
C23 VP.n1 B 0.019635f
C24 VP.n2 B 0.028664f
C25 VP.n3 B 0.019635f
C26 VP.n4 B 0.025393f
C27 VP.t0 B 4.13589f
C28 VP.t2 B 4.12564f
C29 VP.n5 B 3.98211f
C30 VP.t1 B 3.83592f
C31 VP.n6 B 1.39436f
C32 VP.n7 B 1.36555f
C33 VP.n8 B 0.031691f
C34 VP.n9 B 0.019635f
C35 VP.n10 B 0.036595f
C36 VP.n11 B 0.036595f
C37 VP.n12 B 0.028664f
C38 VP.n13 B 0.019635f
C39 VP.n14 B 0.019635f
C40 VP.n15 B 0.019635f
C41 VP.n16 B 0.036595f
C42 VP.n17 B 0.036595f
C43 VP.n18 B 0.025393f
C44 VP.n19 B 0.031691f
C45 VP.n20 B 0.053694f
C46 VTAIL.t6 B 2.78536f
C47 VTAIL.n0 B 0.328922f
C48 VTAIL.t0 B 2.78536f
C49 VTAIL.n1 B 0.409323f
C50 VTAIL.t2 B 2.78536f
C51 VTAIL.n2 B 1.61996f
C52 VTAIL.t7 B 2.78537f
C53 VTAIL.n3 B 1.61995f
C54 VTAIL.t4 B 2.78537f
C55 VTAIL.n4 B 0.409308f
C56 VTAIL.t3 B 2.78537f
C57 VTAIL.n5 B 0.409308f
C58 VTAIL.t1 B 2.78537f
C59 VTAIL.n6 B 1.61995f
C60 VTAIL.t5 B 2.78536f
C61 VTAIL.n7 B 1.53377f
C62 VDD2.t2 B 0.419547f
C63 VDD2.t1 B 0.419547f
C64 VDD2.n0 B 4.88332f
C65 VDD2.t3 B 0.419547f
C66 VDD2.t0 B 0.419547f
C67 VDD2.n1 B 3.83449f
C68 VDD2.n2 B 4.81174f
C69 VN.t2 B 4.07076f
C70 VN.t1 B 4.08087f
C71 VN.n0 B 2.50584f
C72 VN.t3 B 4.08087f
C73 VN.t0 B 4.07076f
C74 VN.n1 B 3.93668f
.ends

