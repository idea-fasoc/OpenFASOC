* NGSPICE file created from diff_pair_sample_1272.ext - technology: sky130A

.subckt diff_pair_sample_1272 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=0 ps=0 w=18.12 l=1.77
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=7.0668 ps=37.02 w=18.12 l=1.77
X2 VDD2.t0 VN.t1 VTAIL.t3 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=7.0668 ps=37.02 w=18.12 l=1.77
X3 B.t8 B.t6 B.t7 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=0 ps=0 w=18.12 l=1.77
X4 VDD1.t1 VP.t0 VTAIL.t1 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=7.0668 ps=37.02 w=18.12 l=1.77
X5 B.t5 B.t3 B.t4 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=0 ps=0 w=18.12 l=1.77
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=7.0668 ps=37.02 w=18.12 l=1.77
X7 B.t2 B.t0 B.t1 w_n1810_n4592# sky130_fd_pr__pfet_01v8 ad=7.0668 pd=37.02 as=0 ps=0 w=18.12 l=1.77
R0 B.n403 B.n102 585
R1 B.n402 B.n401 585
R2 B.n400 B.n103 585
R3 B.n399 B.n398 585
R4 B.n397 B.n104 585
R5 B.n396 B.n395 585
R6 B.n394 B.n105 585
R7 B.n393 B.n392 585
R8 B.n391 B.n106 585
R9 B.n390 B.n389 585
R10 B.n388 B.n107 585
R11 B.n387 B.n386 585
R12 B.n385 B.n108 585
R13 B.n384 B.n383 585
R14 B.n382 B.n109 585
R15 B.n381 B.n380 585
R16 B.n379 B.n110 585
R17 B.n378 B.n377 585
R18 B.n376 B.n111 585
R19 B.n375 B.n374 585
R20 B.n373 B.n112 585
R21 B.n372 B.n371 585
R22 B.n370 B.n113 585
R23 B.n369 B.n368 585
R24 B.n367 B.n114 585
R25 B.n366 B.n365 585
R26 B.n364 B.n115 585
R27 B.n363 B.n362 585
R28 B.n361 B.n116 585
R29 B.n360 B.n359 585
R30 B.n358 B.n117 585
R31 B.n357 B.n356 585
R32 B.n355 B.n118 585
R33 B.n354 B.n353 585
R34 B.n352 B.n119 585
R35 B.n351 B.n350 585
R36 B.n349 B.n120 585
R37 B.n348 B.n347 585
R38 B.n346 B.n121 585
R39 B.n345 B.n344 585
R40 B.n343 B.n122 585
R41 B.n342 B.n341 585
R42 B.n340 B.n123 585
R43 B.n339 B.n338 585
R44 B.n337 B.n124 585
R45 B.n336 B.n335 585
R46 B.n334 B.n125 585
R47 B.n333 B.n332 585
R48 B.n331 B.n126 585
R49 B.n330 B.n329 585
R50 B.n328 B.n127 585
R51 B.n327 B.n326 585
R52 B.n325 B.n128 585
R53 B.n324 B.n323 585
R54 B.n322 B.n129 585
R55 B.n321 B.n320 585
R56 B.n319 B.n130 585
R57 B.n318 B.n317 585
R58 B.n316 B.n131 585
R59 B.n315 B.n314 585
R60 B.n313 B.n312 585
R61 B.n311 B.n135 585
R62 B.n310 B.n309 585
R63 B.n308 B.n136 585
R64 B.n307 B.n306 585
R65 B.n305 B.n137 585
R66 B.n304 B.n303 585
R67 B.n302 B.n138 585
R68 B.n301 B.n300 585
R69 B.n298 B.n139 585
R70 B.n297 B.n296 585
R71 B.n295 B.n142 585
R72 B.n294 B.n293 585
R73 B.n292 B.n143 585
R74 B.n291 B.n290 585
R75 B.n289 B.n144 585
R76 B.n288 B.n287 585
R77 B.n286 B.n145 585
R78 B.n285 B.n284 585
R79 B.n283 B.n146 585
R80 B.n282 B.n281 585
R81 B.n280 B.n147 585
R82 B.n279 B.n278 585
R83 B.n277 B.n148 585
R84 B.n276 B.n275 585
R85 B.n274 B.n149 585
R86 B.n273 B.n272 585
R87 B.n271 B.n150 585
R88 B.n270 B.n269 585
R89 B.n268 B.n151 585
R90 B.n267 B.n266 585
R91 B.n265 B.n152 585
R92 B.n264 B.n263 585
R93 B.n262 B.n153 585
R94 B.n261 B.n260 585
R95 B.n259 B.n154 585
R96 B.n258 B.n257 585
R97 B.n256 B.n155 585
R98 B.n255 B.n254 585
R99 B.n253 B.n156 585
R100 B.n252 B.n251 585
R101 B.n250 B.n157 585
R102 B.n249 B.n248 585
R103 B.n247 B.n158 585
R104 B.n246 B.n245 585
R105 B.n244 B.n159 585
R106 B.n243 B.n242 585
R107 B.n241 B.n160 585
R108 B.n240 B.n239 585
R109 B.n238 B.n161 585
R110 B.n237 B.n236 585
R111 B.n235 B.n162 585
R112 B.n234 B.n233 585
R113 B.n232 B.n163 585
R114 B.n231 B.n230 585
R115 B.n229 B.n164 585
R116 B.n228 B.n227 585
R117 B.n226 B.n165 585
R118 B.n225 B.n224 585
R119 B.n223 B.n166 585
R120 B.n222 B.n221 585
R121 B.n220 B.n167 585
R122 B.n219 B.n218 585
R123 B.n217 B.n168 585
R124 B.n216 B.n215 585
R125 B.n214 B.n169 585
R126 B.n213 B.n212 585
R127 B.n211 B.n170 585
R128 B.n210 B.n209 585
R129 B.n405 B.n404 585
R130 B.n406 B.n101 585
R131 B.n408 B.n407 585
R132 B.n409 B.n100 585
R133 B.n411 B.n410 585
R134 B.n412 B.n99 585
R135 B.n414 B.n413 585
R136 B.n415 B.n98 585
R137 B.n417 B.n416 585
R138 B.n418 B.n97 585
R139 B.n420 B.n419 585
R140 B.n421 B.n96 585
R141 B.n423 B.n422 585
R142 B.n424 B.n95 585
R143 B.n426 B.n425 585
R144 B.n427 B.n94 585
R145 B.n429 B.n428 585
R146 B.n430 B.n93 585
R147 B.n432 B.n431 585
R148 B.n433 B.n92 585
R149 B.n435 B.n434 585
R150 B.n436 B.n91 585
R151 B.n438 B.n437 585
R152 B.n439 B.n90 585
R153 B.n441 B.n440 585
R154 B.n442 B.n89 585
R155 B.n444 B.n443 585
R156 B.n445 B.n88 585
R157 B.n447 B.n446 585
R158 B.n448 B.n87 585
R159 B.n450 B.n449 585
R160 B.n451 B.n86 585
R161 B.n453 B.n452 585
R162 B.n454 B.n85 585
R163 B.n456 B.n455 585
R164 B.n457 B.n84 585
R165 B.n459 B.n458 585
R166 B.n460 B.n83 585
R167 B.n462 B.n461 585
R168 B.n463 B.n82 585
R169 B.n465 B.n464 585
R170 B.n466 B.n81 585
R171 B.n661 B.n12 585
R172 B.n660 B.n659 585
R173 B.n658 B.n13 585
R174 B.n657 B.n656 585
R175 B.n655 B.n14 585
R176 B.n654 B.n653 585
R177 B.n652 B.n15 585
R178 B.n651 B.n650 585
R179 B.n649 B.n16 585
R180 B.n648 B.n647 585
R181 B.n646 B.n17 585
R182 B.n645 B.n644 585
R183 B.n643 B.n18 585
R184 B.n642 B.n641 585
R185 B.n640 B.n19 585
R186 B.n639 B.n638 585
R187 B.n637 B.n20 585
R188 B.n636 B.n635 585
R189 B.n634 B.n21 585
R190 B.n633 B.n632 585
R191 B.n631 B.n22 585
R192 B.n630 B.n629 585
R193 B.n628 B.n23 585
R194 B.n627 B.n626 585
R195 B.n625 B.n24 585
R196 B.n624 B.n623 585
R197 B.n622 B.n25 585
R198 B.n621 B.n620 585
R199 B.n619 B.n26 585
R200 B.n618 B.n617 585
R201 B.n616 B.n27 585
R202 B.n615 B.n614 585
R203 B.n613 B.n28 585
R204 B.n612 B.n611 585
R205 B.n610 B.n29 585
R206 B.n609 B.n608 585
R207 B.n607 B.n30 585
R208 B.n606 B.n605 585
R209 B.n604 B.n31 585
R210 B.n603 B.n602 585
R211 B.n601 B.n32 585
R212 B.n600 B.n599 585
R213 B.n598 B.n33 585
R214 B.n597 B.n596 585
R215 B.n595 B.n34 585
R216 B.n594 B.n593 585
R217 B.n592 B.n35 585
R218 B.n591 B.n590 585
R219 B.n589 B.n36 585
R220 B.n588 B.n587 585
R221 B.n586 B.n37 585
R222 B.n585 B.n584 585
R223 B.n583 B.n38 585
R224 B.n582 B.n581 585
R225 B.n580 B.n39 585
R226 B.n579 B.n578 585
R227 B.n577 B.n40 585
R228 B.n576 B.n575 585
R229 B.n574 B.n41 585
R230 B.n573 B.n572 585
R231 B.n571 B.n570 585
R232 B.n569 B.n45 585
R233 B.n568 B.n567 585
R234 B.n566 B.n46 585
R235 B.n565 B.n564 585
R236 B.n563 B.n47 585
R237 B.n562 B.n561 585
R238 B.n560 B.n48 585
R239 B.n559 B.n558 585
R240 B.n556 B.n49 585
R241 B.n555 B.n554 585
R242 B.n553 B.n52 585
R243 B.n552 B.n551 585
R244 B.n550 B.n53 585
R245 B.n549 B.n548 585
R246 B.n547 B.n54 585
R247 B.n546 B.n545 585
R248 B.n544 B.n55 585
R249 B.n543 B.n542 585
R250 B.n541 B.n56 585
R251 B.n540 B.n539 585
R252 B.n538 B.n57 585
R253 B.n537 B.n536 585
R254 B.n535 B.n58 585
R255 B.n534 B.n533 585
R256 B.n532 B.n59 585
R257 B.n531 B.n530 585
R258 B.n529 B.n60 585
R259 B.n528 B.n527 585
R260 B.n526 B.n61 585
R261 B.n525 B.n524 585
R262 B.n523 B.n62 585
R263 B.n522 B.n521 585
R264 B.n520 B.n63 585
R265 B.n519 B.n518 585
R266 B.n517 B.n64 585
R267 B.n516 B.n515 585
R268 B.n514 B.n65 585
R269 B.n513 B.n512 585
R270 B.n511 B.n66 585
R271 B.n510 B.n509 585
R272 B.n508 B.n67 585
R273 B.n507 B.n506 585
R274 B.n505 B.n68 585
R275 B.n504 B.n503 585
R276 B.n502 B.n69 585
R277 B.n501 B.n500 585
R278 B.n499 B.n70 585
R279 B.n498 B.n497 585
R280 B.n496 B.n71 585
R281 B.n495 B.n494 585
R282 B.n493 B.n72 585
R283 B.n492 B.n491 585
R284 B.n490 B.n73 585
R285 B.n489 B.n488 585
R286 B.n487 B.n74 585
R287 B.n486 B.n485 585
R288 B.n484 B.n75 585
R289 B.n483 B.n482 585
R290 B.n481 B.n76 585
R291 B.n480 B.n479 585
R292 B.n478 B.n77 585
R293 B.n477 B.n476 585
R294 B.n475 B.n78 585
R295 B.n474 B.n473 585
R296 B.n472 B.n79 585
R297 B.n471 B.n470 585
R298 B.n469 B.n80 585
R299 B.n468 B.n467 585
R300 B.n663 B.n662 585
R301 B.n664 B.n11 585
R302 B.n666 B.n665 585
R303 B.n667 B.n10 585
R304 B.n669 B.n668 585
R305 B.n670 B.n9 585
R306 B.n672 B.n671 585
R307 B.n673 B.n8 585
R308 B.n675 B.n674 585
R309 B.n676 B.n7 585
R310 B.n678 B.n677 585
R311 B.n679 B.n6 585
R312 B.n681 B.n680 585
R313 B.n682 B.n5 585
R314 B.n684 B.n683 585
R315 B.n685 B.n4 585
R316 B.n687 B.n686 585
R317 B.n688 B.n3 585
R318 B.n690 B.n689 585
R319 B.n691 B.n0 585
R320 B.n2 B.n1 585
R321 B.n181 B.n180 585
R322 B.n183 B.n182 585
R323 B.n184 B.n179 585
R324 B.n186 B.n185 585
R325 B.n187 B.n178 585
R326 B.n189 B.n188 585
R327 B.n190 B.n177 585
R328 B.n192 B.n191 585
R329 B.n193 B.n176 585
R330 B.n195 B.n194 585
R331 B.n196 B.n175 585
R332 B.n198 B.n197 585
R333 B.n199 B.n174 585
R334 B.n201 B.n200 585
R335 B.n202 B.n173 585
R336 B.n204 B.n203 585
R337 B.n205 B.n172 585
R338 B.n207 B.n206 585
R339 B.n208 B.n171 585
R340 B.n132 B.t4 526.489
R341 B.n50 B.t2 526.489
R342 B.n140 B.t7 526.489
R343 B.n42 B.t11 526.489
R344 B.n133 B.t5 485.762
R345 B.n51 B.t1 485.762
R346 B.n141 B.t8 485.762
R347 B.n43 B.t10 485.762
R348 B.n210 B.n171 478.086
R349 B.n404 B.n403 478.086
R350 B.n468 B.n81 478.086
R351 B.n662 B.n661 478.086
R352 B.n140 B.t6 453.041
R353 B.n132 B.t3 453.041
R354 B.n50 B.t0 453.041
R355 B.n42 B.t9 453.041
R356 B.n693 B.n692 256.663
R357 B.n692 B.n691 235.042
R358 B.n692 B.n2 235.042
R359 B.n211 B.n210 163.367
R360 B.n212 B.n211 163.367
R361 B.n212 B.n169 163.367
R362 B.n216 B.n169 163.367
R363 B.n217 B.n216 163.367
R364 B.n218 B.n217 163.367
R365 B.n218 B.n167 163.367
R366 B.n222 B.n167 163.367
R367 B.n223 B.n222 163.367
R368 B.n224 B.n223 163.367
R369 B.n224 B.n165 163.367
R370 B.n228 B.n165 163.367
R371 B.n229 B.n228 163.367
R372 B.n230 B.n229 163.367
R373 B.n230 B.n163 163.367
R374 B.n234 B.n163 163.367
R375 B.n235 B.n234 163.367
R376 B.n236 B.n235 163.367
R377 B.n236 B.n161 163.367
R378 B.n240 B.n161 163.367
R379 B.n241 B.n240 163.367
R380 B.n242 B.n241 163.367
R381 B.n242 B.n159 163.367
R382 B.n246 B.n159 163.367
R383 B.n247 B.n246 163.367
R384 B.n248 B.n247 163.367
R385 B.n248 B.n157 163.367
R386 B.n252 B.n157 163.367
R387 B.n253 B.n252 163.367
R388 B.n254 B.n253 163.367
R389 B.n254 B.n155 163.367
R390 B.n258 B.n155 163.367
R391 B.n259 B.n258 163.367
R392 B.n260 B.n259 163.367
R393 B.n260 B.n153 163.367
R394 B.n264 B.n153 163.367
R395 B.n265 B.n264 163.367
R396 B.n266 B.n265 163.367
R397 B.n266 B.n151 163.367
R398 B.n270 B.n151 163.367
R399 B.n271 B.n270 163.367
R400 B.n272 B.n271 163.367
R401 B.n272 B.n149 163.367
R402 B.n276 B.n149 163.367
R403 B.n277 B.n276 163.367
R404 B.n278 B.n277 163.367
R405 B.n278 B.n147 163.367
R406 B.n282 B.n147 163.367
R407 B.n283 B.n282 163.367
R408 B.n284 B.n283 163.367
R409 B.n284 B.n145 163.367
R410 B.n288 B.n145 163.367
R411 B.n289 B.n288 163.367
R412 B.n290 B.n289 163.367
R413 B.n290 B.n143 163.367
R414 B.n294 B.n143 163.367
R415 B.n295 B.n294 163.367
R416 B.n296 B.n295 163.367
R417 B.n296 B.n139 163.367
R418 B.n301 B.n139 163.367
R419 B.n302 B.n301 163.367
R420 B.n303 B.n302 163.367
R421 B.n303 B.n137 163.367
R422 B.n307 B.n137 163.367
R423 B.n308 B.n307 163.367
R424 B.n309 B.n308 163.367
R425 B.n309 B.n135 163.367
R426 B.n313 B.n135 163.367
R427 B.n314 B.n313 163.367
R428 B.n314 B.n131 163.367
R429 B.n318 B.n131 163.367
R430 B.n319 B.n318 163.367
R431 B.n320 B.n319 163.367
R432 B.n320 B.n129 163.367
R433 B.n324 B.n129 163.367
R434 B.n325 B.n324 163.367
R435 B.n326 B.n325 163.367
R436 B.n326 B.n127 163.367
R437 B.n330 B.n127 163.367
R438 B.n331 B.n330 163.367
R439 B.n332 B.n331 163.367
R440 B.n332 B.n125 163.367
R441 B.n336 B.n125 163.367
R442 B.n337 B.n336 163.367
R443 B.n338 B.n337 163.367
R444 B.n338 B.n123 163.367
R445 B.n342 B.n123 163.367
R446 B.n343 B.n342 163.367
R447 B.n344 B.n343 163.367
R448 B.n344 B.n121 163.367
R449 B.n348 B.n121 163.367
R450 B.n349 B.n348 163.367
R451 B.n350 B.n349 163.367
R452 B.n350 B.n119 163.367
R453 B.n354 B.n119 163.367
R454 B.n355 B.n354 163.367
R455 B.n356 B.n355 163.367
R456 B.n356 B.n117 163.367
R457 B.n360 B.n117 163.367
R458 B.n361 B.n360 163.367
R459 B.n362 B.n361 163.367
R460 B.n362 B.n115 163.367
R461 B.n366 B.n115 163.367
R462 B.n367 B.n366 163.367
R463 B.n368 B.n367 163.367
R464 B.n368 B.n113 163.367
R465 B.n372 B.n113 163.367
R466 B.n373 B.n372 163.367
R467 B.n374 B.n373 163.367
R468 B.n374 B.n111 163.367
R469 B.n378 B.n111 163.367
R470 B.n379 B.n378 163.367
R471 B.n380 B.n379 163.367
R472 B.n380 B.n109 163.367
R473 B.n384 B.n109 163.367
R474 B.n385 B.n384 163.367
R475 B.n386 B.n385 163.367
R476 B.n386 B.n107 163.367
R477 B.n390 B.n107 163.367
R478 B.n391 B.n390 163.367
R479 B.n392 B.n391 163.367
R480 B.n392 B.n105 163.367
R481 B.n396 B.n105 163.367
R482 B.n397 B.n396 163.367
R483 B.n398 B.n397 163.367
R484 B.n398 B.n103 163.367
R485 B.n402 B.n103 163.367
R486 B.n403 B.n402 163.367
R487 B.n464 B.n81 163.367
R488 B.n464 B.n463 163.367
R489 B.n463 B.n462 163.367
R490 B.n462 B.n83 163.367
R491 B.n458 B.n83 163.367
R492 B.n458 B.n457 163.367
R493 B.n457 B.n456 163.367
R494 B.n456 B.n85 163.367
R495 B.n452 B.n85 163.367
R496 B.n452 B.n451 163.367
R497 B.n451 B.n450 163.367
R498 B.n450 B.n87 163.367
R499 B.n446 B.n87 163.367
R500 B.n446 B.n445 163.367
R501 B.n445 B.n444 163.367
R502 B.n444 B.n89 163.367
R503 B.n440 B.n89 163.367
R504 B.n440 B.n439 163.367
R505 B.n439 B.n438 163.367
R506 B.n438 B.n91 163.367
R507 B.n434 B.n91 163.367
R508 B.n434 B.n433 163.367
R509 B.n433 B.n432 163.367
R510 B.n432 B.n93 163.367
R511 B.n428 B.n93 163.367
R512 B.n428 B.n427 163.367
R513 B.n427 B.n426 163.367
R514 B.n426 B.n95 163.367
R515 B.n422 B.n95 163.367
R516 B.n422 B.n421 163.367
R517 B.n421 B.n420 163.367
R518 B.n420 B.n97 163.367
R519 B.n416 B.n97 163.367
R520 B.n416 B.n415 163.367
R521 B.n415 B.n414 163.367
R522 B.n414 B.n99 163.367
R523 B.n410 B.n99 163.367
R524 B.n410 B.n409 163.367
R525 B.n409 B.n408 163.367
R526 B.n408 B.n101 163.367
R527 B.n404 B.n101 163.367
R528 B.n661 B.n660 163.367
R529 B.n660 B.n13 163.367
R530 B.n656 B.n13 163.367
R531 B.n656 B.n655 163.367
R532 B.n655 B.n654 163.367
R533 B.n654 B.n15 163.367
R534 B.n650 B.n15 163.367
R535 B.n650 B.n649 163.367
R536 B.n649 B.n648 163.367
R537 B.n648 B.n17 163.367
R538 B.n644 B.n17 163.367
R539 B.n644 B.n643 163.367
R540 B.n643 B.n642 163.367
R541 B.n642 B.n19 163.367
R542 B.n638 B.n19 163.367
R543 B.n638 B.n637 163.367
R544 B.n637 B.n636 163.367
R545 B.n636 B.n21 163.367
R546 B.n632 B.n21 163.367
R547 B.n632 B.n631 163.367
R548 B.n631 B.n630 163.367
R549 B.n630 B.n23 163.367
R550 B.n626 B.n23 163.367
R551 B.n626 B.n625 163.367
R552 B.n625 B.n624 163.367
R553 B.n624 B.n25 163.367
R554 B.n620 B.n25 163.367
R555 B.n620 B.n619 163.367
R556 B.n619 B.n618 163.367
R557 B.n618 B.n27 163.367
R558 B.n614 B.n27 163.367
R559 B.n614 B.n613 163.367
R560 B.n613 B.n612 163.367
R561 B.n612 B.n29 163.367
R562 B.n608 B.n29 163.367
R563 B.n608 B.n607 163.367
R564 B.n607 B.n606 163.367
R565 B.n606 B.n31 163.367
R566 B.n602 B.n31 163.367
R567 B.n602 B.n601 163.367
R568 B.n601 B.n600 163.367
R569 B.n600 B.n33 163.367
R570 B.n596 B.n33 163.367
R571 B.n596 B.n595 163.367
R572 B.n595 B.n594 163.367
R573 B.n594 B.n35 163.367
R574 B.n590 B.n35 163.367
R575 B.n590 B.n589 163.367
R576 B.n589 B.n588 163.367
R577 B.n588 B.n37 163.367
R578 B.n584 B.n37 163.367
R579 B.n584 B.n583 163.367
R580 B.n583 B.n582 163.367
R581 B.n582 B.n39 163.367
R582 B.n578 B.n39 163.367
R583 B.n578 B.n577 163.367
R584 B.n577 B.n576 163.367
R585 B.n576 B.n41 163.367
R586 B.n572 B.n41 163.367
R587 B.n572 B.n571 163.367
R588 B.n571 B.n45 163.367
R589 B.n567 B.n45 163.367
R590 B.n567 B.n566 163.367
R591 B.n566 B.n565 163.367
R592 B.n565 B.n47 163.367
R593 B.n561 B.n47 163.367
R594 B.n561 B.n560 163.367
R595 B.n560 B.n559 163.367
R596 B.n559 B.n49 163.367
R597 B.n554 B.n49 163.367
R598 B.n554 B.n553 163.367
R599 B.n553 B.n552 163.367
R600 B.n552 B.n53 163.367
R601 B.n548 B.n53 163.367
R602 B.n548 B.n547 163.367
R603 B.n547 B.n546 163.367
R604 B.n546 B.n55 163.367
R605 B.n542 B.n55 163.367
R606 B.n542 B.n541 163.367
R607 B.n541 B.n540 163.367
R608 B.n540 B.n57 163.367
R609 B.n536 B.n57 163.367
R610 B.n536 B.n535 163.367
R611 B.n535 B.n534 163.367
R612 B.n534 B.n59 163.367
R613 B.n530 B.n59 163.367
R614 B.n530 B.n529 163.367
R615 B.n529 B.n528 163.367
R616 B.n528 B.n61 163.367
R617 B.n524 B.n61 163.367
R618 B.n524 B.n523 163.367
R619 B.n523 B.n522 163.367
R620 B.n522 B.n63 163.367
R621 B.n518 B.n63 163.367
R622 B.n518 B.n517 163.367
R623 B.n517 B.n516 163.367
R624 B.n516 B.n65 163.367
R625 B.n512 B.n65 163.367
R626 B.n512 B.n511 163.367
R627 B.n511 B.n510 163.367
R628 B.n510 B.n67 163.367
R629 B.n506 B.n67 163.367
R630 B.n506 B.n505 163.367
R631 B.n505 B.n504 163.367
R632 B.n504 B.n69 163.367
R633 B.n500 B.n69 163.367
R634 B.n500 B.n499 163.367
R635 B.n499 B.n498 163.367
R636 B.n498 B.n71 163.367
R637 B.n494 B.n71 163.367
R638 B.n494 B.n493 163.367
R639 B.n493 B.n492 163.367
R640 B.n492 B.n73 163.367
R641 B.n488 B.n73 163.367
R642 B.n488 B.n487 163.367
R643 B.n487 B.n486 163.367
R644 B.n486 B.n75 163.367
R645 B.n482 B.n75 163.367
R646 B.n482 B.n481 163.367
R647 B.n481 B.n480 163.367
R648 B.n480 B.n77 163.367
R649 B.n476 B.n77 163.367
R650 B.n476 B.n475 163.367
R651 B.n475 B.n474 163.367
R652 B.n474 B.n79 163.367
R653 B.n470 B.n79 163.367
R654 B.n470 B.n469 163.367
R655 B.n469 B.n468 163.367
R656 B.n662 B.n11 163.367
R657 B.n666 B.n11 163.367
R658 B.n667 B.n666 163.367
R659 B.n668 B.n667 163.367
R660 B.n668 B.n9 163.367
R661 B.n672 B.n9 163.367
R662 B.n673 B.n672 163.367
R663 B.n674 B.n673 163.367
R664 B.n674 B.n7 163.367
R665 B.n678 B.n7 163.367
R666 B.n679 B.n678 163.367
R667 B.n680 B.n679 163.367
R668 B.n680 B.n5 163.367
R669 B.n684 B.n5 163.367
R670 B.n685 B.n684 163.367
R671 B.n686 B.n685 163.367
R672 B.n686 B.n3 163.367
R673 B.n690 B.n3 163.367
R674 B.n691 B.n690 163.367
R675 B.n181 B.n2 163.367
R676 B.n182 B.n181 163.367
R677 B.n182 B.n179 163.367
R678 B.n186 B.n179 163.367
R679 B.n187 B.n186 163.367
R680 B.n188 B.n187 163.367
R681 B.n188 B.n177 163.367
R682 B.n192 B.n177 163.367
R683 B.n193 B.n192 163.367
R684 B.n194 B.n193 163.367
R685 B.n194 B.n175 163.367
R686 B.n198 B.n175 163.367
R687 B.n199 B.n198 163.367
R688 B.n200 B.n199 163.367
R689 B.n200 B.n173 163.367
R690 B.n204 B.n173 163.367
R691 B.n205 B.n204 163.367
R692 B.n206 B.n205 163.367
R693 B.n206 B.n171 163.367
R694 B.n299 B.n141 59.5399
R695 B.n134 B.n133 59.5399
R696 B.n557 B.n51 59.5399
R697 B.n44 B.n43 59.5399
R698 B.n141 B.n140 40.7278
R699 B.n133 B.n132 40.7278
R700 B.n51 B.n50 40.7278
R701 B.n43 B.n42 40.7278
R702 B.n663 B.n12 31.0639
R703 B.n467 B.n466 31.0639
R704 B.n405 B.n102 31.0639
R705 B.n209 B.n208 31.0639
R706 B B.n693 18.0485
R707 B.n664 B.n663 10.6151
R708 B.n665 B.n664 10.6151
R709 B.n665 B.n10 10.6151
R710 B.n669 B.n10 10.6151
R711 B.n670 B.n669 10.6151
R712 B.n671 B.n670 10.6151
R713 B.n671 B.n8 10.6151
R714 B.n675 B.n8 10.6151
R715 B.n676 B.n675 10.6151
R716 B.n677 B.n676 10.6151
R717 B.n677 B.n6 10.6151
R718 B.n681 B.n6 10.6151
R719 B.n682 B.n681 10.6151
R720 B.n683 B.n682 10.6151
R721 B.n683 B.n4 10.6151
R722 B.n687 B.n4 10.6151
R723 B.n688 B.n687 10.6151
R724 B.n689 B.n688 10.6151
R725 B.n689 B.n0 10.6151
R726 B.n659 B.n12 10.6151
R727 B.n659 B.n658 10.6151
R728 B.n658 B.n657 10.6151
R729 B.n657 B.n14 10.6151
R730 B.n653 B.n14 10.6151
R731 B.n653 B.n652 10.6151
R732 B.n652 B.n651 10.6151
R733 B.n651 B.n16 10.6151
R734 B.n647 B.n16 10.6151
R735 B.n647 B.n646 10.6151
R736 B.n646 B.n645 10.6151
R737 B.n645 B.n18 10.6151
R738 B.n641 B.n18 10.6151
R739 B.n641 B.n640 10.6151
R740 B.n640 B.n639 10.6151
R741 B.n639 B.n20 10.6151
R742 B.n635 B.n20 10.6151
R743 B.n635 B.n634 10.6151
R744 B.n634 B.n633 10.6151
R745 B.n633 B.n22 10.6151
R746 B.n629 B.n22 10.6151
R747 B.n629 B.n628 10.6151
R748 B.n628 B.n627 10.6151
R749 B.n627 B.n24 10.6151
R750 B.n623 B.n24 10.6151
R751 B.n623 B.n622 10.6151
R752 B.n622 B.n621 10.6151
R753 B.n621 B.n26 10.6151
R754 B.n617 B.n26 10.6151
R755 B.n617 B.n616 10.6151
R756 B.n616 B.n615 10.6151
R757 B.n615 B.n28 10.6151
R758 B.n611 B.n28 10.6151
R759 B.n611 B.n610 10.6151
R760 B.n610 B.n609 10.6151
R761 B.n609 B.n30 10.6151
R762 B.n605 B.n30 10.6151
R763 B.n605 B.n604 10.6151
R764 B.n604 B.n603 10.6151
R765 B.n603 B.n32 10.6151
R766 B.n599 B.n32 10.6151
R767 B.n599 B.n598 10.6151
R768 B.n598 B.n597 10.6151
R769 B.n597 B.n34 10.6151
R770 B.n593 B.n34 10.6151
R771 B.n593 B.n592 10.6151
R772 B.n592 B.n591 10.6151
R773 B.n591 B.n36 10.6151
R774 B.n587 B.n36 10.6151
R775 B.n587 B.n586 10.6151
R776 B.n586 B.n585 10.6151
R777 B.n585 B.n38 10.6151
R778 B.n581 B.n38 10.6151
R779 B.n581 B.n580 10.6151
R780 B.n580 B.n579 10.6151
R781 B.n579 B.n40 10.6151
R782 B.n575 B.n40 10.6151
R783 B.n575 B.n574 10.6151
R784 B.n574 B.n573 10.6151
R785 B.n570 B.n569 10.6151
R786 B.n569 B.n568 10.6151
R787 B.n568 B.n46 10.6151
R788 B.n564 B.n46 10.6151
R789 B.n564 B.n563 10.6151
R790 B.n563 B.n562 10.6151
R791 B.n562 B.n48 10.6151
R792 B.n558 B.n48 10.6151
R793 B.n556 B.n555 10.6151
R794 B.n555 B.n52 10.6151
R795 B.n551 B.n52 10.6151
R796 B.n551 B.n550 10.6151
R797 B.n550 B.n549 10.6151
R798 B.n549 B.n54 10.6151
R799 B.n545 B.n54 10.6151
R800 B.n545 B.n544 10.6151
R801 B.n544 B.n543 10.6151
R802 B.n543 B.n56 10.6151
R803 B.n539 B.n56 10.6151
R804 B.n539 B.n538 10.6151
R805 B.n538 B.n537 10.6151
R806 B.n537 B.n58 10.6151
R807 B.n533 B.n58 10.6151
R808 B.n533 B.n532 10.6151
R809 B.n532 B.n531 10.6151
R810 B.n531 B.n60 10.6151
R811 B.n527 B.n60 10.6151
R812 B.n527 B.n526 10.6151
R813 B.n526 B.n525 10.6151
R814 B.n525 B.n62 10.6151
R815 B.n521 B.n62 10.6151
R816 B.n521 B.n520 10.6151
R817 B.n520 B.n519 10.6151
R818 B.n519 B.n64 10.6151
R819 B.n515 B.n64 10.6151
R820 B.n515 B.n514 10.6151
R821 B.n514 B.n513 10.6151
R822 B.n513 B.n66 10.6151
R823 B.n509 B.n66 10.6151
R824 B.n509 B.n508 10.6151
R825 B.n508 B.n507 10.6151
R826 B.n507 B.n68 10.6151
R827 B.n503 B.n68 10.6151
R828 B.n503 B.n502 10.6151
R829 B.n502 B.n501 10.6151
R830 B.n501 B.n70 10.6151
R831 B.n497 B.n70 10.6151
R832 B.n497 B.n496 10.6151
R833 B.n496 B.n495 10.6151
R834 B.n495 B.n72 10.6151
R835 B.n491 B.n72 10.6151
R836 B.n491 B.n490 10.6151
R837 B.n490 B.n489 10.6151
R838 B.n489 B.n74 10.6151
R839 B.n485 B.n74 10.6151
R840 B.n485 B.n484 10.6151
R841 B.n484 B.n483 10.6151
R842 B.n483 B.n76 10.6151
R843 B.n479 B.n76 10.6151
R844 B.n479 B.n478 10.6151
R845 B.n478 B.n477 10.6151
R846 B.n477 B.n78 10.6151
R847 B.n473 B.n78 10.6151
R848 B.n473 B.n472 10.6151
R849 B.n472 B.n471 10.6151
R850 B.n471 B.n80 10.6151
R851 B.n467 B.n80 10.6151
R852 B.n466 B.n465 10.6151
R853 B.n465 B.n82 10.6151
R854 B.n461 B.n82 10.6151
R855 B.n461 B.n460 10.6151
R856 B.n460 B.n459 10.6151
R857 B.n459 B.n84 10.6151
R858 B.n455 B.n84 10.6151
R859 B.n455 B.n454 10.6151
R860 B.n454 B.n453 10.6151
R861 B.n453 B.n86 10.6151
R862 B.n449 B.n86 10.6151
R863 B.n449 B.n448 10.6151
R864 B.n448 B.n447 10.6151
R865 B.n447 B.n88 10.6151
R866 B.n443 B.n88 10.6151
R867 B.n443 B.n442 10.6151
R868 B.n442 B.n441 10.6151
R869 B.n441 B.n90 10.6151
R870 B.n437 B.n90 10.6151
R871 B.n437 B.n436 10.6151
R872 B.n436 B.n435 10.6151
R873 B.n435 B.n92 10.6151
R874 B.n431 B.n92 10.6151
R875 B.n431 B.n430 10.6151
R876 B.n430 B.n429 10.6151
R877 B.n429 B.n94 10.6151
R878 B.n425 B.n94 10.6151
R879 B.n425 B.n424 10.6151
R880 B.n424 B.n423 10.6151
R881 B.n423 B.n96 10.6151
R882 B.n419 B.n96 10.6151
R883 B.n419 B.n418 10.6151
R884 B.n418 B.n417 10.6151
R885 B.n417 B.n98 10.6151
R886 B.n413 B.n98 10.6151
R887 B.n413 B.n412 10.6151
R888 B.n412 B.n411 10.6151
R889 B.n411 B.n100 10.6151
R890 B.n407 B.n100 10.6151
R891 B.n407 B.n406 10.6151
R892 B.n406 B.n405 10.6151
R893 B.n180 B.n1 10.6151
R894 B.n183 B.n180 10.6151
R895 B.n184 B.n183 10.6151
R896 B.n185 B.n184 10.6151
R897 B.n185 B.n178 10.6151
R898 B.n189 B.n178 10.6151
R899 B.n190 B.n189 10.6151
R900 B.n191 B.n190 10.6151
R901 B.n191 B.n176 10.6151
R902 B.n195 B.n176 10.6151
R903 B.n196 B.n195 10.6151
R904 B.n197 B.n196 10.6151
R905 B.n197 B.n174 10.6151
R906 B.n201 B.n174 10.6151
R907 B.n202 B.n201 10.6151
R908 B.n203 B.n202 10.6151
R909 B.n203 B.n172 10.6151
R910 B.n207 B.n172 10.6151
R911 B.n208 B.n207 10.6151
R912 B.n209 B.n170 10.6151
R913 B.n213 B.n170 10.6151
R914 B.n214 B.n213 10.6151
R915 B.n215 B.n214 10.6151
R916 B.n215 B.n168 10.6151
R917 B.n219 B.n168 10.6151
R918 B.n220 B.n219 10.6151
R919 B.n221 B.n220 10.6151
R920 B.n221 B.n166 10.6151
R921 B.n225 B.n166 10.6151
R922 B.n226 B.n225 10.6151
R923 B.n227 B.n226 10.6151
R924 B.n227 B.n164 10.6151
R925 B.n231 B.n164 10.6151
R926 B.n232 B.n231 10.6151
R927 B.n233 B.n232 10.6151
R928 B.n233 B.n162 10.6151
R929 B.n237 B.n162 10.6151
R930 B.n238 B.n237 10.6151
R931 B.n239 B.n238 10.6151
R932 B.n239 B.n160 10.6151
R933 B.n243 B.n160 10.6151
R934 B.n244 B.n243 10.6151
R935 B.n245 B.n244 10.6151
R936 B.n245 B.n158 10.6151
R937 B.n249 B.n158 10.6151
R938 B.n250 B.n249 10.6151
R939 B.n251 B.n250 10.6151
R940 B.n251 B.n156 10.6151
R941 B.n255 B.n156 10.6151
R942 B.n256 B.n255 10.6151
R943 B.n257 B.n256 10.6151
R944 B.n257 B.n154 10.6151
R945 B.n261 B.n154 10.6151
R946 B.n262 B.n261 10.6151
R947 B.n263 B.n262 10.6151
R948 B.n263 B.n152 10.6151
R949 B.n267 B.n152 10.6151
R950 B.n268 B.n267 10.6151
R951 B.n269 B.n268 10.6151
R952 B.n269 B.n150 10.6151
R953 B.n273 B.n150 10.6151
R954 B.n274 B.n273 10.6151
R955 B.n275 B.n274 10.6151
R956 B.n275 B.n148 10.6151
R957 B.n279 B.n148 10.6151
R958 B.n280 B.n279 10.6151
R959 B.n281 B.n280 10.6151
R960 B.n281 B.n146 10.6151
R961 B.n285 B.n146 10.6151
R962 B.n286 B.n285 10.6151
R963 B.n287 B.n286 10.6151
R964 B.n287 B.n144 10.6151
R965 B.n291 B.n144 10.6151
R966 B.n292 B.n291 10.6151
R967 B.n293 B.n292 10.6151
R968 B.n293 B.n142 10.6151
R969 B.n297 B.n142 10.6151
R970 B.n298 B.n297 10.6151
R971 B.n300 B.n138 10.6151
R972 B.n304 B.n138 10.6151
R973 B.n305 B.n304 10.6151
R974 B.n306 B.n305 10.6151
R975 B.n306 B.n136 10.6151
R976 B.n310 B.n136 10.6151
R977 B.n311 B.n310 10.6151
R978 B.n312 B.n311 10.6151
R979 B.n316 B.n315 10.6151
R980 B.n317 B.n316 10.6151
R981 B.n317 B.n130 10.6151
R982 B.n321 B.n130 10.6151
R983 B.n322 B.n321 10.6151
R984 B.n323 B.n322 10.6151
R985 B.n323 B.n128 10.6151
R986 B.n327 B.n128 10.6151
R987 B.n328 B.n327 10.6151
R988 B.n329 B.n328 10.6151
R989 B.n329 B.n126 10.6151
R990 B.n333 B.n126 10.6151
R991 B.n334 B.n333 10.6151
R992 B.n335 B.n334 10.6151
R993 B.n335 B.n124 10.6151
R994 B.n339 B.n124 10.6151
R995 B.n340 B.n339 10.6151
R996 B.n341 B.n340 10.6151
R997 B.n341 B.n122 10.6151
R998 B.n345 B.n122 10.6151
R999 B.n346 B.n345 10.6151
R1000 B.n347 B.n346 10.6151
R1001 B.n347 B.n120 10.6151
R1002 B.n351 B.n120 10.6151
R1003 B.n352 B.n351 10.6151
R1004 B.n353 B.n352 10.6151
R1005 B.n353 B.n118 10.6151
R1006 B.n357 B.n118 10.6151
R1007 B.n358 B.n357 10.6151
R1008 B.n359 B.n358 10.6151
R1009 B.n359 B.n116 10.6151
R1010 B.n363 B.n116 10.6151
R1011 B.n364 B.n363 10.6151
R1012 B.n365 B.n364 10.6151
R1013 B.n365 B.n114 10.6151
R1014 B.n369 B.n114 10.6151
R1015 B.n370 B.n369 10.6151
R1016 B.n371 B.n370 10.6151
R1017 B.n371 B.n112 10.6151
R1018 B.n375 B.n112 10.6151
R1019 B.n376 B.n375 10.6151
R1020 B.n377 B.n376 10.6151
R1021 B.n377 B.n110 10.6151
R1022 B.n381 B.n110 10.6151
R1023 B.n382 B.n381 10.6151
R1024 B.n383 B.n382 10.6151
R1025 B.n383 B.n108 10.6151
R1026 B.n387 B.n108 10.6151
R1027 B.n388 B.n387 10.6151
R1028 B.n389 B.n388 10.6151
R1029 B.n389 B.n106 10.6151
R1030 B.n393 B.n106 10.6151
R1031 B.n394 B.n393 10.6151
R1032 B.n395 B.n394 10.6151
R1033 B.n395 B.n104 10.6151
R1034 B.n399 B.n104 10.6151
R1035 B.n400 B.n399 10.6151
R1036 B.n401 B.n400 10.6151
R1037 B.n401 B.n102 10.6151
R1038 B.n693 B.n0 8.11757
R1039 B.n693 B.n1 8.11757
R1040 B.n570 B.n44 6.5566
R1041 B.n558 B.n557 6.5566
R1042 B.n300 B.n299 6.5566
R1043 B.n312 B.n134 6.5566
R1044 B.n573 B.n44 4.05904
R1045 B.n557 B.n556 4.05904
R1046 B.n299 B.n298 4.05904
R1047 B.n315 B.n134 4.05904
R1048 VN VN.t0 352.887
R1049 VN VN.t1 305.846
R1050 VTAIL.n402 VTAIL.n306 756.745
R1051 VTAIL.n96 VTAIL.n0 756.745
R1052 VTAIL.n300 VTAIL.n204 756.745
R1053 VTAIL.n198 VTAIL.n102 756.745
R1054 VTAIL.n338 VTAIL.n337 585
R1055 VTAIL.n343 VTAIL.n342 585
R1056 VTAIL.n345 VTAIL.n344 585
R1057 VTAIL.n334 VTAIL.n333 585
R1058 VTAIL.n351 VTAIL.n350 585
R1059 VTAIL.n353 VTAIL.n352 585
R1060 VTAIL.n330 VTAIL.n329 585
R1061 VTAIL.n359 VTAIL.n358 585
R1062 VTAIL.n361 VTAIL.n360 585
R1063 VTAIL.n326 VTAIL.n325 585
R1064 VTAIL.n367 VTAIL.n366 585
R1065 VTAIL.n369 VTAIL.n368 585
R1066 VTAIL.n322 VTAIL.n321 585
R1067 VTAIL.n375 VTAIL.n374 585
R1068 VTAIL.n377 VTAIL.n376 585
R1069 VTAIL.n318 VTAIL.n317 585
R1070 VTAIL.n384 VTAIL.n383 585
R1071 VTAIL.n385 VTAIL.n316 585
R1072 VTAIL.n387 VTAIL.n386 585
R1073 VTAIL.n314 VTAIL.n313 585
R1074 VTAIL.n393 VTAIL.n392 585
R1075 VTAIL.n395 VTAIL.n394 585
R1076 VTAIL.n310 VTAIL.n309 585
R1077 VTAIL.n401 VTAIL.n400 585
R1078 VTAIL.n403 VTAIL.n402 585
R1079 VTAIL.n32 VTAIL.n31 585
R1080 VTAIL.n37 VTAIL.n36 585
R1081 VTAIL.n39 VTAIL.n38 585
R1082 VTAIL.n28 VTAIL.n27 585
R1083 VTAIL.n45 VTAIL.n44 585
R1084 VTAIL.n47 VTAIL.n46 585
R1085 VTAIL.n24 VTAIL.n23 585
R1086 VTAIL.n53 VTAIL.n52 585
R1087 VTAIL.n55 VTAIL.n54 585
R1088 VTAIL.n20 VTAIL.n19 585
R1089 VTAIL.n61 VTAIL.n60 585
R1090 VTAIL.n63 VTAIL.n62 585
R1091 VTAIL.n16 VTAIL.n15 585
R1092 VTAIL.n69 VTAIL.n68 585
R1093 VTAIL.n71 VTAIL.n70 585
R1094 VTAIL.n12 VTAIL.n11 585
R1095 VTAIL.n78 VTAIL.n77 585
R1096 VTAIL.n79 VTAIL.n10 585
R1097 VTAIL.n81 VTAIL.n80 585
R1098 VTAIL.n8 VTAIL.n7 585
R1099 VTAIL.n87 VTAIL.n86 585
R1100 VTAIL.n89 VTAIL.n88 585
R1101 VTAIL.n4 VTAIL.n3 585
R1102 VTAIL.n95 VTAIL.n94 585
R1103 VTAIL.n97 VTAIL.n96 585
R1104 VTAIL.n301 VTAIL.n300 585
R1105 VTAIL.n299 VTAIL.n298 585
R1106 VTAIL.n208 VTAIL.n207 585
R1107 VTAIL.n293 VTAIL.n292 585
R1108 VTAIL.n291 VTAIL.n290 585
R1109 VTAIL.n212 VTAIL.n211 585
R1110 VTAIL.n285 VTAIL.n284 585
R1111 VTAIL.n283 VTAIL.n214 585
R1112 VTAIL.n282 VTAIL.n281 585
R1113 VTAIL.n217 VTAIL.n215 585
R1114 VTAIL.n276 VTAIL.n275 585
R1115 VTAIL.n274 VTAIL.n273 585
R1116 VTAIL.n221 VTAIL.n220 585
R1117 VTAIL.n268 VTAIL.n267 585
R1118 VTAIL.n266 VTAIL.n265 585
R1119 VTAIL.n225 VTAIL.n224 585
R1120 VTAIL.n260 VTAIL.n259 585
R1121 VTAIL.n258 VTAIL.n257 585
R1122 VTAIL.n229 VTAIL.n228 585
R1123 VTAIL.n252 VTAIL.n251 585
R1124 VTAIL.n250 VTAIL.n249 585
R1125 VTAIL.n233 VTAIL.n232 585
R1126 VTAIL.n244 VTAIL.n243 585
R1127 VTAIL.n242 VTAIL.n241 585
R1128 VTAIL.n237 VTAIL.n236 585
R1129 VTAIL.n199 VTAIL.n198 585
R1130 VTAIL.n197 VTAIL.n196 585
R1131 VTAIL.n106 VTAIL.n105 585
R1132 VTAIL.n191 VTAIL.n190 585
R1133 VTAIL.n189 VTAIL.n188 585
R1134 VTAIL.n110 VTAIL.n109 585
R1135 VTAIL.n183 VTAIL.n182 585
R1136 VTAIL.n181 VTAIL.n112 585
R1137 VTAIL.n180 VTAIL.n179 585
R1138 VTAIL.n115 VTAIL.n113 585
R1139 VTAIL.n174 VTAIL.n173 585
R1140 VTAIL.n172 VTAIL.n171 585
R1141 VTAIL.n119 VTAIL.n118 585
R1142 VTAIL.n166 VTAIL.n165 585
R1143 VTAIL.n164 VTAIL.n163 585
R1144 VTAIL.n123 VTAIL.n122 585
R1145 VTAIL.n158 VTAIL.n157 585
R1146 VTAIL.n156 VTAIL.n155 585
R1147 VTAIL.n127 VTAIL.n126 585
R1148 VTAIL.n150 VTAIL.n149 585
R1149 VTAIL.n148 VTAIL.n147 585
R1150 VTAIL.n131 VTAIL.n130 585
R1151 VTAIL.n142 VTAIL.n141 585
R1152 VTAIL.n140 VTAIL.n139 585
R1153 VTAIL.n135 VTAIL.n134 585
R1154 VTAIL.n339 VTAIL.t3 327.466
R1155 VTAIL.n33 VTAIL.t0 327.466
R1156 VTAIL.n238 VTAIL.t1 327.466
R1157 VTAIL.n136 VTAIL.t2 327.466
R1158 VTAIL.n343 VTAIL.n337 171.744
R1159 VTAIL.n344 VTAIL.n343 171.744
R1160 VTAIL.n344 VTAIL.n333 171.744
R1161 VTAIL.n351 VTAIL.n333 171.744
R1162 VTAIL.n352 VTAIL.n351 171.744
R1163 VTAIL.n352 VTAIL.n329 171.744
R1164 VTAIL.n359 VTAIL.n329 171.744
R1165 VTAIL.n360 VTAIL.n359 171.744
R1166 VTAIL.n360 VTAIL.n325 171.744
R1167 VTAIL.n367 VTAIL.n325 171.744
R1168 VTAIL.n368 VTAIL.n367 171.744
R1169 VTAIL.n368 VTAIL.n321 171.744
R1170 VTAIL.n375 VTAIL.n321 171.744
R1171 VTAIL.n376 VTAIL.n375 171.744
R1172 VTAIL.n376 VTAIL.n317 171.744
R1173 VTAIL.n384 VTAIL.n317 171.744
R1174 VTAIL.n385 VTAIL.n384 171.744
R1175 VTAIL.n386 VTAIL.n385 171.744
R1176 VTAIL.n386 VTAIL.n313 171.744
R1177 VTAIL.n393 VTAIL.n313 171.744
R1178 VTAIL.n394 VTAIL.n393 171.744
R1179 VTAIL.n394 VTAIL.n309 171.744
R1180 VTAIL.n401 VTAIL.n309 171.744
R1181 VTAIL.n402 VTAIL.n401 171.744
R1182 VTAIL.n37 VTAIL.n31 171.744
R1183 VTAIL.n38 VTAIL.n37 171.744
R1184 VTAIL.n38 VTAIL.n27 171.744
R1185 VTAIL.n45 VTAIL.n27 171.744
R1186 VTAIL.n46 VTAIL.n45 171.744
R1187 VTAIL.n46 VTAIL.n23 171.744
R1188 VTAIL.n53 VTAIL.n23 171.744
R1189 VTAIL.n54 VTAIL.n53 171.744
R1190 VTAIL.n54 VTAIL.n19 171.744
R1191 VTAIL.n61 VTAIL.n19 171.744
R1192 VTAIL.n62 VTAIL.n61 171.744
R1193 VTAIL.n62 VTAIL.n15 171.744
R1194 VTAIL.n69 VTAIL.n15 171.744
R1195 VTAIL.n70 VTAIL.n69 171.744
R1196 VTAIL.n70 VTAIL.n11 171.744
R1197 VTAIL.n78 VTAIL.n11 171.744
R1198 VTAIL.n79 VTAIL.n78 171.744
R1199 VTAIL.n80 VTAIL.n79 171.744
R1200 VTAIL.n80 VTAIL.n7 171.744
R1201 VTAIL.n87 VTAIL.n7 171.744
R1202 VTAIL.n88 VTAIL.n87 171.744
R1203 VTAIL.n88 VTAIL.n3 171.744
R1204 VTAIL.n95 VTAIL.n3 171.744
R1205 VTAIL.n96 VTAIL.n95 171.744
R1206 VTAIL.n300 VTAIL.n299 171.744
R1207 VTAIL.n299 VTAIL.n207 171.744
R1208 VTAIL.n292 VTAIL.n207 171.744
R1209 VTAIL.n292 VTAIL.n291 171.744
R1210 VTAIL.n291 VTAIL.n211 171.744
R1211 VTAIL.n284 VTAIL.n211 171.744
R1212 VTAIL.n284 VTAIL.n283 171.744
R1213 VTAIL.n283 VTAIL.n282 171.744
R1214 VTAIL.n282 VTAIL.n215 171.744
R1215 VTAIL.n275 VTAIL.n215 171.744
R1216 VTAIL.n275 VTAIL.n274 171.744
R1217 VTAIL.n274 VTAIL.n220 171.744
R1218 VTAIL.n267 VTAIL.n220 171.744
R1219 VTAIL.n267 VTAIL.n266 171.744
R1220 VTAIL.n266 VTAIL.n224 171.744
R1221 VTAIL.n259 VTAIL.n224 171.744
R1222 VTAIL.n259 VTAIL.n258 171.744
R1223 VTAIL.n258 VTAIL.n228 171.744
R1224 VTAIL.n251 VTAIL.n228 171.744
R1225 VTAIL.n251 VTAIL.n250 171.744
R1226 VTAIL.n250 VTAIL.n232 171.744
R1227 VTAIL.n243 VTAIL.n232 171.744
R1228 VTAIL.n243 VTAIL.n242 171.744
R1229 VTAIL.n242 VTAIL.n236 171.744
R1230 VTAIL.n198 VTAIL.n197 171.744
R1231 VTAIL.n197 VTAIL.n105 171.744
R1232 VTAIL.n190 VTAIL.n105 171.744
R1233 VTAIL.n190 VTAIL.n189 171.744
R1234 VTAIL.n189 VTAIL.n109 171.744
R1235 VTAIL.n182 VTAIL.n109 171.744
R1236 VTAIL.n182 VTAIL.n181 171.744
R1237 VTAIL.n181 VTAIL.n180 171.744
R1238 VTAIL.n180 VTAIL.n113 171.744
R1239 VTAIL.n173 VTAIL.n113 171.744
R1240 VTAIL.n173 VTAIL.n172 171.744
R1241 VTAIL.n172 VTAIL.n118 171.744
R1242 VTAIL.n165 VTAIL.n118 171.744
R1243 VTAIL.n165 VTAIL.n164 171.744
R1244 VTAIL.n164 VTAIL.n122 171.744
R1245 VTAIL.n157 VTAIL.n122 171.744
R1246 VTAIL.n157 VTAIL.n156 171.744
R1247 VTAIL.n156 VTAIL.n126 171.744
R1248 VTAIL.n149 VTAIL.n126 171.744
R1249 VTAIL.n149 VTAIL.n148 171.744
R1250 VTAIL.n148 VTAIL.n130 171.744
R1251 VTAIL.n141 VTAIL.n130 171.744
R1252 VTAIL.n141 VTAIL.n140 171.744
R1253 VTAIL.n140 VTAIL.n134 171.744
R1254 VTAIL.t3 VTAIL.n337 85.8723
R1255 VTAIL.t0 VTAIL.n31 85.8723
R1256 VTAIL.t1 VTAIL.n236 85.8723
R1257 VTAIL.t2 VTAIL.n134 85.8723
R1258 VTAIL.n203 VTAIL.n101 31.6083
R1259 VTAIL.n407 VTAIL.n406 29.8581
R1260 VTAIL.n101 VTAIL.n100 29.8581
R1261 VTAIL.n305 VTAIL.n304 29.8581
R1262 VTAIL.n203 VTAIL.n202 29.8581
R1263 VTAIL.n407 VTAIL.n305 29.7979
R1264 VTAIL.n339 VTAIL.n338 16.3895
R1265 VTAIL.n33 VTAIL.n32 16.3895
R1266 VTAIL.n238 VTAIL.n237 16.3895
R1267 VTAIL.n136 VTAIL.n135 16.3895
R1268 VTAIL.n387 VTAIL.n316 13.1884
R1269 VTAIL.n81 VTAIL.n10 13.1884
R1270 VTAIL.n285 VTAIL.n214 13.1884
R1271 VTAIL.n183 VTAIL.n112 13.1884
R1272 VTAIL.n342 VTAIL.n341 12.8005
R1273 VTAIL.n383 VTAIL.n382 12.8005
R1274 VTAIL.n388 VTAIL.n314 12.8005
R1275 VTAIL.n36 VTAIL.n35 12.8005
R1276 VTAIL.n77 VTAIL.n76 12.8005
R1277 VTAIL.n82 VTAIL.n8 12.8005
R1278 VTAIL.n286 VTAIL.n212 12.8005
R1279 VTAIL.n281 VTAIL.n216 12.8005
R1280 VTAIL.n241 VTAIL.n240 12.8005
R1281 VTAIL.n184 VTAIL.n110 12.8005
R1282 VTAIL.n179 VTAIL.n114 12.8005
R1283 VTAIL.n139 VTAIL.n138 12.8005
R1284 VTAIL.n345 VTAIL.n336 12.0247
R1285 VTAIL.n381 VTAIL.n318 12.0247
R1286 VTAIL.n392 VTAIL.n391 12.0247
R1287 VTAIL.n39 VTAIL.n30 12.0247
R1288 VTAIL.n75 VTAIL.n12 12.0247
R1289 VTAIL.n86 VTAIL.n85 12.0247
R1290 VTAIL.n290 VTAIL.n289 12.0247
R1291 VTAIL.n280 VTAIL.n217 12.0247
R1292 VTAIL.n244 VTAIL.n235 12.0247
R1293 VTAIL.n188 VTAIL.n187 12.0247
R1294 VTAIL.n178 VTAIL.n115 12.0247
R1295 VTAIL.n142 VTAIL.n133 12.0247
R1296 VTAIL.n346 VTAIL.n334 11.249
R1297 VTAIL.n378 VTAIL.n377 11.249
R1298 VTAIL.n395 VTAIL.n312 11.249
R1299 VTAIL.n40 VTAIL.n28 11.249
R1300 VTAIL.n72 VTAIL.n71 11.249
R1301 VTAIL.n89 VTAIL.n6 11.249
R1302 VTAIL.n293 VTAIL.n210 11.249
R1303 VTAIL.n277 VTAIL.n276 11.249
R1304 VTAIL.n245 VTAIL.n233 11.249
R1305 VTAIL.n191 VTAIL.n108 11.249
R1306 VTAIL.n175 VTAIL.n174 11.249
R1307 VTAIL.n143 VTAIL.n131 11.249
R1308 VTAIL.n350 VTAIL.n349 10.4732
R1309 VTAIL.n374 VTAIL.n320 10.4732
R1310 VTAIL.n396 VTAIL.n310 10.4732
R1311 VTAIL.n44 VTAIL.n43 10.4732
R1312 VTAIL.n68 VTAIL.n14 10.4732
R1313 VTAIL.n90 VTAIL.n4 10.4732
R1314 VTAIL.n294 VTAIL.n208 10.4732
R1315 VTAIL.n273 VTAIL.n219 10.4732
R1316 VTAIL.n249 VTAIL.n248 10.4732
R1317 VTAIL.n192 VTAIL.n106 10.4732
R1318 VTAIL.n171 VTAIL.n117 10.4732
R1319 VTAIL.n147 VTAIL.n146 10.4732
R1320 VTAIL.n353 VTAIL.n332 9.69747
R1321 VTAIL.n373 VTAIL.n322 9.69747
R1322 VTAIL.n400 VTAIL.n399 9.69747
R1323 VTAIL.n47 VTAIL.n26 9.69747
R1324 VTAIL.n67 VTAIL.n16 9.69747
R1325 VTAIL.n94 VTAIL.n93 9.69747
R1326 VTAIL.n298 VTAIL.n297 9.69747
R1327 VTAIL.n272 VTAIL.n221 9.69747
R1328 VTAIL.n252 VTAIL.n231 9.69747
R1329 VTAIL.n196 VTAIL.n195 9.69747
R1330 VTAIL.n170 VTAIL.n119 9.69747
R1331 VTAIL.n150 VTAIL.n129 9.69747
R1332 VTAIL.n406 VTAIL.n405 9.45567
R1333 VTAIL.n100 VTAIL.n99 9.45567
R1334 VTAIL.n304 VTAIL.n303 9.45567
R1335 VTAIL.n202 VTAIL.n201 9.45567
R1336 VTAIL.n405 VTAIL.n404 9.3005
R1337 VTAIL.n308 VTAIL.n307 9.3005
R1338 VTAIL.n399 VTAIL.n398 9.3005
R1339 VTAIL.n397 VTAIL.n396 9.3005
R1340 VTAIL.n312 VTAIL.n311 9.3005
R1341 VTAIL.n391 VTAIL.n390 9.3005
R1342 VTAIL.n389 VTAIL.n388 9.3005
R1343 VTAIL.n328 VTAIL.n327 9.3005
R1344 VTAIL.n357 VTAIL.n356 9.3005
R1345 VTAIL.n355 VTAIL.n354 9.3005
R1346 VTAIL.n332 VTAIL.n331 9.3005
R1347 VTAIL.n349 VTAIL.n348 9.3005
R1348 VTAIL.n347 VTAIL.n346 9.3005
R1349 VTAIL.n336 VTAIL.n335 9.3005
R1350 VTAIL.n341 VTAIL.n340 9.3005
R1351 VTAIL.n363 VTAIL.n362 9.3005
R1352 VTAIL.n365 VTAIL.n364 9.3005
R1353 VTAIL.n324 VTAIL.n323 9.3005
R1354 VTAIL.n371 VTAIL.n370 9.3005
R1355 VTAIL.n373 VTAIL.n372 9.3005
R1356 VTAIL.n320 VTAIL.n319 9.3005
R1357 VTAIL.n379 VTAIL.n378 9.3005
R1358 VTAIL.n381 VTAIL.n380 9.3005
R1359 VTAIL.n382 VTAIL.n315 9.3005
R1360 VTAIL.n99 VTAIL.n98 9.3005
R1361 VTAIL.n2 VTAIL.n1 9.3005
R1362 VTAIL.n93 VTAIL.n92 9.3005
R1363 VTAIL.n91 VTAIL.n90 9.3005
R1364 VTAIL.n6 VTAIL.n5 9.3005
R1365 VTAIL.n85 VTAIL.n84 9.3005
R1366 VTAIL.n83 VTAIL.n82 9.3005
R1367 VTAIL.n22 VTAIL.n21 9.3005
R1368 VTAIL.n51 VTAIL.n50 9.3005
R1369 VTAIL.n49 VTAIL.n48 9.3005
R1370 VTAIL.n26 VTAIL.n25 9.3005
R1371 VTAIL.n43 VTAIL.n42 9.3005
R1372 VTAIL.n41 VTAIL.n40 9.3005
R1373 VTAIL.n30 VTAIL.n29 9.3005
R1374 VTAIL.n35 VTAIL.n34 9.3005
R1375 VTAIL.n57 VTAIL.n56 9.3005
R1376 VTAIL.n59 VTAIL.n58 9.3005
R1377 VTAIL.n18 VTAIL.n17 9.3005
R1378 VTAIL.n65 VTAIL.n64 9.3005
R1379 VTAIL.n67 VTAIL.n66 9.3005
R1380 VTAIL.n14 VTAIL.n13 9.3005
R1381 VTAIL.n73 VTAIL.n72 9.3005
R1382 VTAIL.n75 VTAIL.n74 9.3005
R1383 VTAIL.n76 VTAIL.n9 9.3005
R1384 VTAIL.n264 VTAIL.n263 9.3005
R1385 VTAIL.n223 VTAIL.n222 9.3005
R1386 VTAIL.n270 VTAIL.n269 9.3005
R1387 VTAIL.n272 VTAIL.n271 9.3005
R1388 VTAIL.n219 VTAIL.n218 9.3005
R1389 VTAIL.n278 VTAIL.n277 9.3005
R1390 VTAIL.n280 VTAIL.n279 9.3005
R1391 VTAIL.n216 VTAIL.n213 9.3005
R1392 VTAIL.n303 VTAIL.n302 9.3005
R1393 VTAIL.n206 VTAIL.n205 9.3005
R1394 VTAIL.n297 VTAIL.n296 9.3005
R1395 VTAIL.n295 VTAIL.n294 9.3005
R1396 VTAIL.n210 VTAIL.n209 9.3005
R1397 VTAIL.n289 VTAIL.n288 9.3005
R1398 VTAIL.n287 VTAIL.n286 9.3005
R1399 VTAIL.n262 VTAIL.n261 9.3005
R1400 VTAIL.n227 VTAIL.n226 9.3005
R1401 VTAIL.n256 VTAIL.n255 9.3005
R1402 VTAIL.n254 VTAIL.n253 9.3005
R1403 VTAIL.n231 VTAIL.n230 9.3005
R1404 VTAIL.n248 VTAIL.n247 9.3005
R1405 VTAIL.n246 VTAIL.n245 9.3005
R1406 VTAIL.n235 VTAIL.n234 9.3005
R1407 VTAIL.n240 VTAIL.n239 9.3005
R1408 VTAIL.n162 VTAIL.n161 9.3005
R1409 VTAIL.n121 VTAIL.n120 9.3005
R1410 VTAIL.n168 VTAIL.n167 9.3005
R1411 VTAIL.n170 VTAIL.n169 9.3005
R1412 VTAIL.n117 VTAIL.n116 9.3005
R1413 VTAIL.n176 VTAIL.n175 9.3005
R1414 VTAIL.n178 VTAIL.n177 9.3005
R1415 VTAIL.n114 VTAIL.n111 9.3005
R1416 VTAIL.n201 VTAIL.n200 9.3005
R1417 VTAIL.n104 VTAIL.n103 9.3005
R1418 VTAIL.n195 VTAIL.n194 9.3005
R1419 VTAIL.n193 VTAIL.n192 9.3005
R1420 VTAIL.n108 VTAIL.n107 9.3005
R1421 VTAIL.n187 VTAIL.n186 9.3005
R1422 VTAIL.n185 VTAIL.n184 9.3005
R1423 VTAIL.n160 VTAIL.n159 9.3005
R1424 VTAIL.n125 VTAIL.n124 9.3005
R1425 VTAIL.n154 VTAIL.n153 9.3005
R1426 VTAIL.n152 VTAIL.n151 9.3005
R1427 VTAIL.n129 VTAIL.n128 9.3005
R1428 VTAIL.n146 VTAIL.n145 9.3005
R1429 VTAIL.n144 VTAIL.n143 9.3005
R1430 VTAIL.n133 VTAIL.n132 9.3005
R1431 VTAIL.n138 VTAIL.n137 9.3005
R1432 VTAIL.n354 VTAIL.n330 8.92171
R1433 VTAIL.n370 VTAIL.n369 8.92171
R1434 VTAIL.n403 VTAIL.n308 8.92171
R1435 VTAIL.n48 VTAIL.n24 8.92171
R1436 VTAIL.n64 VTAIL.n63 8.92171
R1437 VTAIL.n97 VTAIL.n2 8.92171
R1438 VTAIL.n301 VTAIL.n206 8.92171
R1439 VTAIL.n269 VTAIL.n268 8.92171
R1440 VTAIL.n253 VTAIL.n229 8.92171
R1441 VTAIL.n199 VTAIL.n104 8.92171
R1442 VTAIL.n167 VTAIL.n166 8.92171
R1443 VTAIL.n151 VTAIL.n127 8.92171
R1444 VTAIL.n358 VTAIL.n357 8.14595
R1445 VTAIL.n366 VTAIL.n324 8.14595
R1446 VTAIL.n404 VTAIL.n306 8.14595
R1447 VTAIL.n52 VTAIL.n51 8.14595
R1448 VTAIL.n60 VTAIL.n18 8.14595
R1449 VTAIL.n98 VTAIL.n0 8.14595
R1450 VTAIL.n302 VTAIL.n204 8.14595
R1451 VTAIL.n265 VTAIL.n223 8.14595
R1452 VTAIL.n257 VTAIL.n256 8.14595
R1453 VTAIL.n200 VTAIL.n102 8.14595
R1454 VTAIL.n163 VTAIL.n121 8.14595
R1455 VTAIL.n155 VTAIL.n154 8.14595
R1456 VTAIL.n361 VTAIL.n328 7.3702
R1457 VTAIL.n365 VTAIL.n326 7.3702
R1458 VTAIL.n55 VTAIL.n22 7.3702
R1459 VTAIL.n59 VTAIL.n20 7.3702
R1460 VTAIL.n264 VTAIL.n225 7.3702
R1461 VTAIL.n260 VTAIL.n227 7.3702
R1462 VTAIL.n162 VTAIL.n123 7.3702
R1463 VTAIL.n158 VTAIL.n125 7.3702
R1464 VTAIL.n362 VTAIL.n361 6.59444
R1465 VTAIL.n362 VTAIL.n326 6.59444
R1466 VTAIL.n56 VTAIL.n55 6.59444
R1467 VTAIL.n56 VTAIL.n20 6.59444
R1468 VTAIL.n261 VTAIL.n225 6.59444
R1469 VTAIL.n261 VTAIL.n260 6.59444
R1470 VTAIL.n159 VTAIL.n123 6.59444
R1471 VTAIL.n159 VTAIL.n158 6.59444
R1472 VTAIL.n358 VTAIL.n328 5.81868
R1473 VTAIL.n366 VTAIL.n365 5.81868
R1474 VTAIL.n406 VTAIL.n306 5.81868
R1475 VTAIL.n52 VTAIL.n22 5.81868
R1476 VTAIL.n60 VTAIL.n59 5.81868
R1477 VTAIL.n100 VTAIL.n0 5.81868
R1478 VTAIL.n304 VTAIL.n204 5.81868
R1479 VTAIL.n265 VTAIL.n264 5.81868
R1480 VTAIL.n257 VTAIL.n227 5.81868
R1481 VTAIL.n202 VTAIL.n102 5.81868
R1482 VTAIL.n163 VTAIL.n162 5.81868
R1483 VTAIL.n155 VTAIL.n125 5.81868
R1484 VTAIL.n357 VTAIL.n330 5.04292
R1485 VTAIL.n369 VTAIL.n324 5.04292
R1486 VTAIL.n404 VTAIL.n403 5.04292
R1487 VTAIL.n51 VTAIL.n24 5.04292
R1488 VTAIL.n63 VTAIL.n18 5.04292
R1489 VTAIL.n98 VTAIL.n97 5.04292
R1490 VTAIL.n302 VTAIL.n301 5.04292
R1491 VTAIL.n268 VTAIL.n223 5.04292
R1492 VTAIL.n256 VTAIL.n229 5.04292
R1493 VTAIL.n200 VTAIL.n199 5.04292
R1494 VTAIL.n166 VTAIL.n121 5.04292
R1495 VTAIL.n154 VTAIL.n127 5.04292
R1496 VTAIL.n354 VTAIL.n353 4.26717
R1497 VTAIL.n370 VTAIL.n322 4.26717
R1498 VTAIL.n400 VTAIL.n308 4.26717
R1499 VTAIL.n48 VTAIL.n47 4.26717
R1500 VTAIL.n64 VTAIL.n16 4.26717
R1501 VTAIL.n94 VTAIL.n2 4.26717
R1502 VTAIL.n298 VTAIL.n206 4.26717
R1503 VTAIL.n269 VTAIL.n221 4.26717
R1504 VTAIL.n253 VTAIL.n252 4.26717
R1505 VTAIL.n196 VTAIL.n104 4.26717
R1506 VTAIL.n167 VTAIL.n119 4.26717
R1507 VTAIL.n151 VTAIL.n150 4.26717
R1508 VTAIL.n340 VTAIL.n339 3.70982
R1509 VTAIL.n34 VTAIL.n33 3.70982
R1510 VTAIL.n239 VTAIL.n238 3.70982
R1511 VTAIL.n137 VTAIL.n136 3.70982
R1512 VTAIL.n350 VTAIL.n332 3.49141
R1513 VTAIL.n374 VTAIL.n373 3.49141
R1514 VTAIL.n399 VTAIL.n310 3.49141
R1515 VTAIL.n44 VTAIL.n26 3.49141
R1516 VTAIL.n68 VTAIL.n67 3.49141
R1517 VTAIL.n93 VTAIL.n4 3.49141
R1518 VTAIL.n297 VTAIL.n208 3.49141
R1519 VTAIL.n273 VTAIL.n272 3.49141
R1520 VTAIL.n249 VTAIL.n231 3.49141
R1521 VTAIL.n195 VTAIL.n106 3.49141
R1522 VTAIL.n171 VTAIL.n170 3.49141
R1523 VTAIL.n147 VTAIL.n129 3.49141
R1524 VTAIL.n349 VTAIL.n334 2.71565
R1525 VTAIL.n377 VTAIL.n320 2.71565
R1526 VTAIL.n396 VTAIL.n395 2.71565
R1527 VTAIL.n43 VTAIL.n28 2.71565
R1528 VTAIL.n71 VTAIL.n14 2.71565
R1529 VTAIL.n90 VTAIL.n89 2.71565
R1530 VTAIL.n294 VTAIL.n293 2.71565
R1531 VTAIL.n276 VTAIL.n219 2.71565
R1532 VTAIL.n248 VTAIL.n233 2.71565
R1533 VTAIL.n192 VTAIL.n191 2.71565
R1534 VTAIL.n174 VTAIL.n117 2.71565
R1535 VTAIL.n146 VTAIL.n131 2.71565
R1536 VTAIL.n346 VTAIL.n345 1.93989
R1537 VTAIL.n378 VTAIL.n318 1.93989
R1538 VTAIL.n392 VTAIL.n312 1.93989
R1539 VTAIL.n40 VTAIL.n39 1.93989
R1540 VTAIL.n72 VTAIL.n12 1.93989
R1541 VTAIL.n86 VTAIL.n6 1.93989
R1542 VTAIL.n290 VTAIL.n210 1.93989
R1543 VTAIL.n277 VTAIL.n217 1.93989
R1544 VTAIL.n245 VTAIL.n244 1.93989
R1545 VTAIL.n188 VTAIL.n108 1.93989
R1546 VTAIL.n175 VTAIL.n115 1.93989
R1547 VTAIL.n143 VTAIL.n142 1.93989
R1548 VTAIL.n305 VTAIL.n203 1.3755
R1549 VTAIL.n342 VTAIL.n336 1.16414
R1550 VTAIL.n383 VTAIL.n381 1.16414
R1551 VTAIL.n391 VTAIL.n314 1.16414
R1552 VTAIL.n36 VTAIL.n30 1.16414
R1553 VTAIL.n77 VTAIL.n75 1.16414
R1554 VTAIL.n85 VTAIL.n8 1.16414
R1555 VTAIL.n289 VTAIL.n212 1.16414
R1556 VTAIL.n281 VTAIL.n280 1.16414
R1557 VTAIL.n241 VTAIL.n235 1.16414
R1558 VTAIL.n187 VTAIL.n110 1.16414
R1559 VTAIL.n179 VTAIL.n178 1.16414
R1560 VTAIL.n139 VTAIL.n133 1.16414
R1561 VTAIL VTAIL.n101 0.981103
R1562 VTAIL VTAIL.n407 0.394897
R1563 VTAIL.n341 VTAIL.n338 0.388379
R1564 VTAIL.n382 VTAIL.n316 0.388379
R1565 VTAIL.n388 VTAIL.n387 0.388379
R1566 VTAIL.n35 VTAIL.n32 0.388379
R1567 VTAIL.n76 VTAIL.n10 0.388379
R1568 VTAIL.n82 VTAIL.n81 0.388379
R1569 VTAIL.n286 VTAIL.n285 0.388379
R1570 VTAIL.n216 VTAIL.n214 0.388379
R1571 VTAIL.n240 VTAIL.n237 0.388379
R1572 VTAIL.n184 VTAIL.n183 0.388379
R1573 VTAIL.n114 VTAIL.n112 0.388379
R1574 VTAIL.n138 VTAIL.n135 0.388379
R1575 VTAIL.n340 VTAIL.n335 0.155672
R1576 VTAIL.n347 VTAIL.n335 0.155672
R1577 VTAIL.n348 VTAIL.n347 0.155672
R1578 VTAIL.n348 VTAIL.n331 0.155672
R1579 VTAIL.n355 VTAIL.n331 0.155672
R1580 VTAIL.n356 VTAIL.n355 0.155672
R1581 VTAIL.n356 VTAIL.n327 0.155672
R1582 VTAIL.n363 VTAIL.n327 0.155672
R1583 VTAIL.n364 VTAIL.n363 0.155672
R1584 VTAIL.n364 VTAIL.n323 0.155672
R1585 VTAIL.n371 VTAIL.n323 0.155672
R1586 VTAIL.n372 VTAIL.n371 0.155672
R1587 VTAIL.n372 VTAIL.n319 0.155672
R1588 VTAIL.n379 VTAIL.n319 0.155672
R1589 VTAIL.n380 VTAIL.n379 0.155672
R1590 VTAIL.n380 VTAIL.n315 0.155672
R1591 VTAIL.n389 VTAIL.n315 0.155672
R1592 VTAIL.n390 VTAIL.n389 0.155672
R1593 VTAIL.n390 VTAIL.n311 0.155672
R1594 VTAIL.n397 VTAIL.n311 0.155672
R1595 VTAIL.n398 VTAIL.n397 0.155672
R1596 VTAIL.n398 VTAIL.n307 0.155672
R1597 VTAIL.n405 VTAIL.n307 0.155672
R1598 VTAIL.n34 VTAIL.n29 0.155672
R1599 VTAIL.n41 VTAIL.n29 0.155672
R1600 VTAIL.n42 VTAIL.n41 0.155672
R1601 VTAIL.n42 VTAIL.n25 0.155672
R1602 VTAIL.n49 VTAIL.n25 0.155672
R1603 VTAIL.n50 VTAIL.n49 0.155672
R1604 VTAIL.n50 VTAIL.n21 0.155672
R1605 VTAIL.n57 VTAIL.n21 0.155672
R1606 VTAIL.n58 VTAIL.n57 0.155672
R1607 VTAIL.n58 VTAIL.n17 0.155672
R1608 VTAIL.n65 VTAIL.n17 0.155672
R1609 VTAIL.n66 VTAIL.n65 0.155672
R1610 VTAIL.n66 VTAIL.n13 0.155672
R1611 VTAIL.n73 VTAIL.n13 0.155672
R1612 VTAIL.n74 VTAIL.n73 0.155672
R1613 VTAIL.n74 VTAIL.n9 0.155672
R1614 VTAIL.n83 VTAIL.n9 0.155672
R1615 VTAIL.n84 VTAIL.n83 0.155672
R1616 VTAIL.n84 VTAIL.n5 0.155672
R1617 VTAIL.n91 VTAIL.n5 0.155672
R1618 VTAIL.n92 VTAIL.n91 0.155672
R1619 VTAIL.n92 VTAIL.n1 0.155672
R1620 VTAIL.n99 VTAIL.n1 0.155672
R1621 VTAIL.n303 VTAIL.n205 0.155672
R1622 VTAIL.n296 VTAIL.n205 0.155672
R1623 VTAIL.n296 VTAIL.n295 0.155672
R1624 VTAIL.n295 VTAIL.n209 0.155672
R1625 VTAIL.n288 VTAIL.n209 0.155672
R1626 VTAIL.n288 VTAIL.n287 0.155672
R1627 VTAIL.n287 VTAIL.n213 0.155672
R1628 VTAIL.n279 VTAIL.n213 0.155672
R1629 VTAIL.n279 VTAIL.n278 0.155672
R1630 VTAIL.n278 VTAIL.n218 0.155672
R1631 VTAIL.n271 VTAIL.n218 0.155672
R1632 VTAIL.n271 VTAIL.n270 0.155672
R1633 VTAIL.n270 VTAIL.n222 0.155672
R1634 VTAIL.n263 VTAIL.n222 0.155672
R1635 VTAIL.n263 VTAIL.n262 0.155672
R1636 VTAIL.n262 VTAIL.n226 0.155672
R1637 VTAIL.n255 VTAIL.n226 0.155672
R1638 VTAIL.n255 VTAIL.n254 0.155672
R1639 VTAIL.n254 VTAIL.n230 0.155672
R1640 VTAIL.n247 VTAIL.n230 0.155672
R1641 VTAIL.n247 VTAIL.n246 0.155672
R1642 VTAIL.n246 VTAIL.n234 0.155672
R1643 VTAIL.n239 VTAIL.n234 0.155672
R1644 VTAIL.n201 VTAIL.n103 0.155672
R1645 VTAIL.n194 VTAIL.n103 0.155672
R1646 VTAIL.n194 VTAIL.n193 0.155672
R1647 VTAIL.n193 VTAIL.n107 0.155672
R1648 VTAIL.n186 VTAIL.n107 0.155672
R1649 VTAIL.n186 VTAIL.n185 0.155672
R1650 VTAIL.n185 VTAIL.n111 0.155672
R1651 VTAIL.n177 VTAIL.n111 0.155672
R1652 VTAIL.n177 VTAIL.n176 0.155672
R1653 VTAIL.n176 VTAIL.n116 0.155672
R1654 VTAIL.n169 VTAIL.n116 0.155672
R1655 VTAIL.n169 VTAIL.n168 0.155672
R1656 VTAIL.n168 VTAIL.n120 0.155672
R1657 VTAIL.n161 VTAIL.n120 0.155672
R1658 VTAIL.n161 VTAIL.n160 0.155672
R1659 VTAIL.n160 VTAIL.n124 0.155672
R1660 VTAIL.n153 VTAIL.n124 0.155672
R1661 VTAIL.n153 VTAIL.n152 0.155672
R1662 VTAIL.n152 VTAIL.n128 0.155672
R1663 VTAIL.n145 VTAIL.n128 0.155672
R1664 VTAIL.n145 VTAIL.n144 0.155672
R1665 VTAIL.n144 VTAIL.n132 0.155672
R1666 VTAIL.n137 VTAIL.n132 0.155672
R1667 VDD2.n197 VDD2.n101 756.745
R1668 VDD2.n96 VDD2.n0 756.745
R1669 VDD2.n198 VDD2.n197 585
R1670 VDD2.n196 VDD2.n195 585
R1671 VDD2.n105 VDD2.n104 585
R1672 VDD2.n190 VDD2.n189 585
R1673 VDD2.n188 VDD2.n187 585
R1674 VDD2.n109 VDD2.n108 585
R1675 VDD2.n182 VDD2.n181 585
R1676 VDD2.n180 VDD2.n111 585
R1677 VDD2.n179 VDD2.n178 585
R1678 VDD2.n114 VDD2.n112 585
R1679 VDD2.n173 VDD2.n172 585
R1680 VDD2.n171 VDD2.n170 585
R1681 VDD2.n118 VDD2.n117 585
R1682 VDD2.n165 VDD2.n164 585
R1683 VDD2.n163 VDD2.n162 585
R1684 VDD2.n122 VDD2.n121 585
R1685 VDD2.n157 VDD2.n156 585
R1686 VDD2.n155 VDD2.n154 585
R1687 VDD2.n126 VDD2.n125 585
R1688 VDD2.n149 VDD2.n148 585
R1689 VDD2.n147 VDD2.n146 585
R1690 VDD2.n130 VDD2.n129 585
R1691 VDD2.n141 VDD2.n140 585
R1692 VDD2.n139 VDD2.n138 585
R1693 VDD2.n134 VDD2.n133 585
R1694 VDD2.n32 VDD2.n31 585
R1695 VDD2.n37 VDD2.n36 585
R1696 VDD2.n39 VDD2.n38 585
R1697 VDD2.n28 VDD2.n27 585
R1698 VDD2.n45 VDD2.n44 585
R1699 VDD2.n47 VDD2.n46 585
R1700 VDD2.n24 VDD2.n23 585
R1701 VDD2.n53 VDD2.n52 585
R1702 VDD2.n55 VDD2.n54 585
R1703 VDD2.n20 VDD2.n19 585
R1704 VDD2.n61 VDD2.n60 585
R1705 VDD2.n63 VDD2.n62 585
R1706 VDD2.n16 VDD2.n15 585
R1707 VDD2.n69 VDD2.n68 585
R1708 VDD2.n71 VDD2.n70 585
R1709 VDD2.n12 VDD2.n11 585
R1710 VDD2.n78 VDD2.n77 585
R1711 VDD2.n79 VDD2.n10 585
R1712 VDD2.n81 VDD2.n80 585
R1713 VDD2.n8 VDD2.n7 585
R1714 VDD2.n87 VDD2.n86 585
R1715 VDD2.n89 VDD2.n88 585
R1716 VDD2.n4 VDD2.n3 585
R1717 VDD2.n95 VDD2.n94 585
R1718 VDD2.n97 VDD2.n96 585
R1719 VDD2.n135 VDD2.t1 327.466
R1720 VDD2.n33 VDD2.t0 327.466
R1721 VDD2.n197 VDD2.n196 171.744
R1722 VDD2.n196 VDD2.n104 171.744
R1723 VDD2.n189 VDD2.n104 171.744
R1724 VDD2.n189 VDD2.n188 171.744
R1725 VDD2.n188 VDD2.n108 171.744
R1726 VDD2.n181 VDD2.n108 171.744
R1727 VDD2.n181 VDD2.n180 171.744
R1728 VDD2.n180 VDD2.n179 171.744
R1729 VDD2.n179 VDD2.n112 171.744
R1730 VDD2.n172 VDD2.n112 171.744
R1731 VDD2.n172 VDD2.n171 171.744
R1732 VDD2.n171 VDD2.n117 171.744
R1733 VDD2.n164 VDD2.n117 171.744
R1734 VDD2.n164 VDD2.n163 171.744
R1735 VDD2.n163 VDD2.n121 171.744
R1736 VDD2.n156 VDD2.n121 171.744
R1737 VDD2.n156 VDD2.n155 171.744
R1738 VDD2.n155 VDD2.n125 171.744
R1739 VDD2.n148 VDD2.n125 171.744
R1740 VDD2.n148 VDD2.n147 171.744
R1741 VDD2.n147 VDD2.n129 171.744
R1742 VDD2.n140 VDD2.n129 171.744
R1743 VDD2.n140 VDD2.n139 171.744
R1744 VDD2.n139 VDD2.n133 171.744
R1745 VDD2.n37 VDD2.n31 171.744
R1746 VDD2.n38 VDD2.n37 171.744
R1747 VDD2.n38 VDD2.n27 171.744
R1748 VDD2.n45 VDD2.n27 171.744
R1749 VDD2.n46 VDD2.n45 171.744
R1750 VDD2.n46 VDD2.n23 171.744
R1751 VDD2.n53 VDD2.n23 171.744
R1752 VDD2.n54 VDD2.n53 171.744
R1753 VDD2.n54 VDD2.n19 171.744
R1754 VDD2.n61 VDD2.n19 171.744
R1755 VDD2.n62 VDD2.n61 171.744
R1756 VDD2.n62 VDD2.n15 171.744
R1757 VDD2.n69 VDD2.n15 171.744
R1758 VDD2.n70 VDD2.n69 171.744
R1759 VDD2.n70 VDD2.n11 171.744
R1760 VDD2.n78 VDD2.n11 171.744
R1761 VDD2.n79 VDD2.n78 171.744
R1762 VDD2.n80 VDD2.n79 171.744
R1763 VDD2.n80 VDD2.n7 171.744
R1764 VDD2.n87 VDD2.n7 171.744
R1765 VDD2.n88 VDD2.n87 171.744
R1766 VDD2.n88 VDD2.n3 171.744
R1767 VDD2.n95 VDD2.n3 171.744
R1768 VDD2.n96 VDD2.n95 171.744
R1769 VDD2.n202 VDD2.n100 89.4377
R1770 VDD2.t1 VDD2.n133 85.8723
R1771 VDD2.t0 VDD2.n31 85.8723
R1772 VDD2.n202 VDD2.n201 46.5369
R1773 VDD2.n135 VDD2.n134 16.3895
R1774 VDD2.n33 VDD2.n32 16.3895
R1775 VDD2.n182 VDD2.n111 13.1884
R1776 VDD2.n81 VDD2.n10 13.1884
R1777 VDD2.n183 VDD2.n109 12.8005
R1778 VDD2.n178 VDD2.n113 12.8005
R1779 VDD2.n138 VDD2.n137 12.8005
R1780 VDD2.n36 VDD2.n35 12.8005
R1781 VDD2.n77 VDD2.n76 12.8005
R1782 VDD2.n82 VDD2.n8 12.8005
R1783 VDD2.n187 VDD2.n186 12.0247
R1784 VDD2.n177 VDD2.n114 12.0247
R1785 VDD2.n141 VDD2.n132 12.0247
R1786 VDD2.n39 VDD2.n30 12.0247
R1787 VDD2.n75 VDD2.n12 12.0247
R1788 VDD2.n86 VDD2.n85 12.0247
R1789 VDD2.n190 VDD2.n107 11.249
R1790 VDD2.n174 VDD2.n173 11.249
R1791 VDD2.n142 VDD2.n130 11.249
R1792 VDD2.n40 VDD2.n28 11.249
R1793 VDD2.n72 VDD2.n71 11.249
R1794 VDD2.n89 VDD2.n6 11.249
R1795 VDD2.n191 VDD2.n105 10.4732
R1796 VDD2.n170 VDD2.n116 10.4732
R1797 VDD2.n146 VDD2.n145 10.4732
R1798 VDD2.n44 VDD2.n43 10.4732
R1799 VDD2.n68 VDD2.n14 10.4732
R1800 VDD2.n90 VDD2.n4 10.4732
R1801 VDD2.n195 VDD2.n194 9.69747
R1802 VDD2.n169 VDD2.n118 9.69747
R1803 VDD2.n149 VDD2.n128 9.69747
R1804 VDD2.n47 VDD2.n26 9.69747
R1805 VDD2.n67 VDD2.n16 9.69747
R1806 VDD2.n94 VDD2.n93 9.69747
R1807 VDD2.n201 VDD2.n200 9.45567
R1808 VDD2.n100 VDD2.n99 9.45567
R1809 VDD2.n161 VDD2.n160 9.3005
R1810 VDD2.n120 VDD2.n119 9.3005
R1811 VDD2.n167 VDD2.n166 9.3005
R1812 VDD2.n169 VDD2.n168 9.3005
R1813 VDD2.n116 VDD2.n115 9.3005
R1814 VDD2.n175 VDD2.n174 9.3005
R1815 VDD2.n177 VDD2.n176 9.3005
R1816 VDD2.n113 VDD2.n110 9.3005
R1817 VDD2.n200 VDD2.n199 9.3005
R1818 VDD2.n103 VDD2.n102 9.3005
R1819 VDD2.n194 VDD2.n193 9.3005
R1820 VDD2.n192 VDD2.n191 9.3005
R1821 VDD2.n107 VDD2.n106 9.3005
R1822 VDD2.n186 VDD2.n185 9.3005
R1823 VDD2.n184 VDD2.n183 9.3005
R1824 VDD2.n159 VDD2.n158 9.3005
R1825 VDD2.n124 VDD2.n123 9.3005
R1826 VDD2.n153 VDD2.n152 9.3005
R1827 VDD2.n151 VDD2.n150 9.3005
R1828 VDD2.n128 VDD2.n127 9.3005
R1829 VDD2.n145 VDD2.n144 9.3005
R1830 VDD2.n143 VDD2.n142 9.3005
R1831 VDD2.n132 VDD2.n131 9.3005
R1832 VDD2.n137 VDD2.n136 9.3005
R1833 VDD2.n99 VDD2.n98 9.3005
R1834 VDD2.n2 VDD2.n1 9.3005
R1835 VDD2.n93 VDD2.n92 9.3005
R1836 VDD2.n91 VDD2.n90 9.3005
R1837 VDD2.n6 VDD2.n5 9.3005
R1838 VDD2.n85 VDD2.n84 9.3005
R1839 VDD2.n83 VDD2.n82 9.3005
R1840 VDD2.n22 VDD2.n21 9.3005
R1841 VDD2.n51 VDD2.n50 9.3005
R1842 VDD2.n49 VDD2.n48 9.3005
R1843 VDD2.n26 VDD2.n25 9.3005
R1844 VDD2.n43 VDD2.n42 9.3005
R1845 VDD2.n41 VDD2.n40 9.3005
R1846 VDD2.n30 VDD2.n29 9.3005
R1847 VDD2.n35 VDD2.n34 9.3005
R1848 VDD2.n57 VDD2.n56 9.3005
R1849 VDD2.n59 VDD2.n58 9.3005
R1850 VDD2.n18 VDD2.n17 9.3005
R1851 VDD2.n65 VDD2.n64 9.3005
R1852 VDD2.n67 VDD2.n66 9.3005
R1853 VDD2.n14 VDD2.n13 9.3005
R1854 VDD2.n73 VDD2.n72 9.3005
R1855 VDD2.n75 VDD2.n74 9.3005
R1856 VDD2.n76 VDD2.n9 9.3005
R1857 VDD2.n198 VDD2.n103 8.92171
R1858 VDD2.n166 VDD2.n165 8.92171
R1859 VDD2.n150 VDD2.n126 8.92171
R1860 VDD2.n48 VDD2.n24 8.92171
R1861 VDD2.n64 VDD2.n63 8.92171
R1862 VDD2.n97 VDD2.n2 8.92171
R1863 VDD2.n199 VDD2.n101 8.14595
R1864 VDD2.n162 VDD2.n120 8.14595
R1865 VDD2.n154 VDD2.n153 8.14595
R1866 VDD2.n52 VDD2.n51 8.14595
R1867 VDD2.n60 VDD2.n18 8.14595
R1868 VDD2.n98 VDD2.n0 8.14595
R1869 VDD2.n161 VDD2.n122 7.3702
R1870 VDD2.n157 VDD2.n124 7.3702
R1871 VDD2.n55 VDD2.n22 7.3702
R1872 VDD2.n59 VDD2.n20 7.3702
R1873 VDD2.n158 VDD2.n122 6.59444
R1874 VDD2.n158 VDD2.n157 6.59444
R1875 VDD2.n56 VDD2.n55 6.59444
R1876 VDD2.n56 VDD2.n20 6.59444
R1877 VDD2.n201 VDD2.n101 5.81868
R1878 VDD2.n162 VDD2.n161 5.81868
R1879 VDD2.n154 VDD2.n124 5.81868
R1880 VDD2.n52 VDD2.n22 5.81868
R1881 VDD2.n60 VDD2.n59 5.81868
R1882 VDD2.n100 VDD2.n0 5.81868
R1883 VDD2.n199 VDD2.n198 5.04292
R1884 VDD2.n165 VDD2.n120 5.04292
R1885 VDD2.n153 VDD2.n126 5.04292
R1886 VDD2.n51 VDD2.n24 5.04292
R1887 VDD2.n63 VDD2.n18 5.04292
R1888 VDD2.n98 VDD2.n97 5.04292
R1889 VDD2.n195 VDD2.n103 4.26717
R1890 VDD2.n166 VDD2.n118 4.26717
R1891 VDD2.n150 VDD2.n149 4.26717
R1892 VDD2.n48 VDD2.n47 4.26717
R1893 VDD2.n64 VDD2.n16 4.26717
R1894 VDD2.n94 VDD2.n2 4.26717
R1895 VDD2.n136 VDD2.n135 3.70982
R1896 VDD2.n34 VDD2.n33 3.70982
R1897 VDD2.n194 VDD2.n105 3.49141
R1898 VDD2.n170 VDD2.n169 3.49141
R1899 VDD2.n146 VDD2.n128 3.49141
R1900 VDD2.n44 VDD2.n26 3.49141
R1901 VDD2.n68 VDD2.n67 3.49141
R1902 VDD2.n93 VDD2.n4 3.49141
R1903 VDD2.n191 VDD2.n190 2.71565
R1904 VDD2.n173 VDD2.n116 2.71565
R1905 VDD2.n145 VDD2.n130 2.71565
R1906 VDD2.n43 VDD2.n28 2.71565
R1907 VDD2.n71 VDD2.n14 2.71565
R1908 VDD2.n90 VDD2.n89 2.71565
R1909 VDD2.n187 VDD2.n107 1.93989
R1910 VDD2.n174 VDD2.n114 1.93989
R1911 VDD2.n142 VDD2.n141 1.93989
R1912 VDD2.n40 VDD2.n39 1.93989
R1913 VDD2.n72 VDD2.n12 1.93989
R1914 VDD2.n86 VDD2.n6 1.93989
R1915 VDD2.n186 VDD2.n109 1.16414
R1916 VDD2.n178 VDD2.n177 1.16414
R1917 VDD2.n138 VDD2.n132 1.16414
R1918 VDD2.n36 VDD2.n30 1.16414
R1919 VDD2.n77 VDD2.n75 1.16414
R1920 VDD2.n85 VDD2.n8 1.16414
R1921 VDD2 VDD2.n202 0.511276
R1922 VDD2.n183 VDD2.n182 0.388379
R1923 VDD2.n113 VDD2.n111 0.388379
R1924 VDD2.n137 VDD2.n134 0.388379
R1925 VDD2.n35 VDD2.n32 0.388379
R1926 VDD2.n76 VDD2.n10 0.388379
R1927 VDD2.n82 VDD2.n81 0.388379
R1928 VDD2.n200 VDD2.n102 0.155672
R1929 VDD2.n193 VDD2.n102 0.155672
R1930 VDD2.n193 VDD2.n192 0.155672
R1931 VDD2.n192 VDD2.n106 0.155672
R1932 VDD2.n185 VDD2.n106 0.155672
R1933 VDD2.n185 VDD2.n184 0.155672
R1934 VDD2.n184 VDD2.n110 0.155672
R1935 VDD2.n176 VDD2.n110 0.155672
R1936 VDD2.n176 VDD2.n175 0.155672
R1937 VDD2.n175 VDD2.n115 0.155672
R1938 VDD2.n168 VDD2.n115 0.155672
R1939 VDD2.n168 VDD2.n167 0.155672
R1940 VDD2.n167 VDD2.n119 0.155672
R1941 VDD2.n160 VDD2.n119 0.155672
R1942 VDD2.n160 VDD2.n159 0.155672
R1943 VDD2.n159 VDD2.n123 0.155672
R1944 VDD2.n152 VDD2.n123 0.155672
R1945 VDD2.n152 VDD2.n151 0.155672
R1946 VDD2.n151 VDD2.n127 0.155672
R1947 VDD2.n144 VDD2.n127 0.155672
R1948 VDD2.n144 VDD2.n143 0.155672
R1949 VDD2.n143 VDD2.n131 0.155672
R1950 VDD2.n136 VDD2.n131 0.155672
R1951 VDD2.n34 VDD2.n29 0.155672
R1952 VDD2.n41 VDD2.n29 0.155672
R1953 VDD2.n42 VDD2.n41 0.155672
R1954 VDD2.n42 VDD2.n25 0.155672
R1955 VDD2.n49 VDD2.n25 0.155672
R1956 VDD2.n50 VDD2.n49 0.155672
R1957 VDD2.n50 VDD2.n21 0.155672
R1958 VDD2.n57 VDD2.n21 0.155672
R1959 VDD2.n58 VDD2.n57 0.155672
R1960 VDD2.n58 VDD2.n17 0.155672
R1961 VDD2.n65 VDD2.n17 0.155672
R1962 VDD2.n66 VDD2.n65 0.155672
R1963 VDD2.n66 VDD2.n13 0.155672
R1964 VDD2.n73 VDD2.n13 0.155672
R1965 VDD2.n74 VDD2.n73 0.155672
R1966 VDD2.n74 VDD2.n9 0.155672
R1967 VDD2.n83 VDD2.n9 0.155672
R1968 VDD2.n84 VDD2.n83 0.155672
R1969 VDD2.n84 VDD2.n5 0.155672
R1970 VDD2.n91 VDD2.n5 0.155672
R1971 VDD2.n92 VDD2.n91 0.155672
R1972 VDD2.n92 VDD2.n1 0.155672
R1973 VDD2.n99 VDD2.n1 0.155672
R1974 VP.n0 VP.t0 352.697
R1975 VP.n0 VP.t1 305.606
R1976 VP VP.n0 0.241678
R1977 VDD1.n96 VDD1.n0 756.745
R1978 VDD1.n197 VDD1.n101 756.745
R1979 VDD1.n97 VDD1.n96 585
R1980 VDD1.n95 VDD1.n94 585
R1981 VDD1.n4 VDD1.n3 585
R1982 VDD1.n89 VDD1.n88 585
R1983 VDD1.n87 VDD1.n86 585
R1984 VDD1.n8 VDD1.n7 585
R1985 VDD1.n81 VDD1.n80 585
R1986 VDD1.n79 VDD1.n10 585
R1987 VDD1.n78 VDD1.n77 585
R1988 VDD1.n13 VDD1.n11 585
R1989 VDD1.n72 VDD1.n71 585
R1990 VDD1.n70 VDD1.n69 585
R1991 VDD1.n17 VDD1.n16 585
R1992 VDD1.n64 VDD1.n63 585
R1993 VDD1.n62 VDD1.n61 585
R1994 VDD1.n21 VDD1.n20 585
R1995 VDD1.n56 VDD1.n55 585
R1996 VDD1.n54 VDD1.n53 585
R1997 VDD1.n25 VDD1.n24 585
R1998 VDD1.n48 VDD1.n47 585
R1999 VDD1.n46 VDD1.n45 585
R2000 VDD1.n29 VDD1.n28 585
R2001 VDD1.n40 VDD1.n39 585
R2002 VDD1.n38 VDD1.n37 585
R2003 VDD1.n33 VDD1.n32 585
R2004 VDD1.n133 VDD1.n132 585
R2005 VDD1.n138 VDD1.n137 585
R2006 VDD1.n140 VDD1.n139 585
R2007 VDD1.n129 VDD1.n128 585
R2008 VDD1.n146 VDD1.n145 585
R2009 VDD1.n148 VDD1.n147 585
R2010 VDD1.n125 VDD1.n124 585
R2011 VDD1.n154 VDD1.n153 585
R2012 VDD1.n156 VDD1.n155 585
R2013 VDD1.n121 VDD1.n120 585
R2014 VDD1.n162 VDD1.n161 585
R2015 VDD1.n164 VDD1.n163 585
R2016 VDD1.n117 VDD1.n116 585
R2017 VDD1.n170 VDD1.n169 585
R2018 VDD1.n172 VDD1.n171 585
R2019 VDD1.n113 VDD1.n112 585
R2020 VDD1.n179 VDD1.n178 585
R2021 VDD1.n180 VDD1.n111 585
R2022 VDD1.n182 VDD1.n181 585
R2023 VDD1.n109 VDD1.n108 585
R2024 VDD1.n188 VDD1.n187 585
R2025 VDD1.n190 VDD1.n189 585
R2026 VDD1.n105 VDD1.n104 585
R2027 VDD1.n196 VDD1.n195 585
R2028 VDD1.n198 VDD1.n197 585
R2029 VDD1.n34 VDD1.t1 327.466
R2030 VDD1.n134 VDD1.t0 327.466
R2031 VDD1.n96 VDD1.n95 171.744
R2032 VDD1.n95 VDD1.n3 171.744
R2033 VDD1.n88 VDD1.n3 171.744
R2034 VDD1.n88 VDD1.n87 171.744
R2035 VDD1.n87 VDD1.n7 171.744
R2036 VDD1.n80 VDD1.n7 171.744
R2037 VDD1.n80 VDD1.n79 171.744
R2038 VDD1.n79 VDD1.n78 171.744
R2039 VDD1.n78 VDD1.n11 171.744
R2040 VDD1.n71 VDD1.n11 171.744
R2041 VDD1.n71 VDD1.n70 171.744
R2042 VDD1.n70 VDD1.n16 171.744
R2043 VDD1.n63 VDD1.n16 171.744
R2044 VDD1.n63 VDD1.n62 171.744
R2045 VDD1.n62 VDD1.n20 171.744
R2046 VDD1.n55 VDD1.n20 171.744
R2047 VDD1.n55 VDD1.n54 171.744
R2048 VDD1.n54 VDD1.n24 171.744
R2049 VDD1.n47 VDD1.n24 171.744
R2050 VDD1.n47 VDD1.n46 171.744
R2051 VDD1.n46 VDD1.n28 171.744
R2052 VDD1.n39 VDD1.n28 171.744
R2053 VDD1.n39 VDD1.n38 171.744
R2054 VDD1.n38 VDD1.n32 171.744
R2055 VDD1.n138 VDD1.n132 171.744
R2056 VDD1.n139 VDD1.n138 171.744
R2057 VDD1.n139 VDD1.n128 171.744
R2058 VDD1.n146 VDD1.n128 171.744
R2059 VDD1.n147 VDD1.n146 171.744
R2060 VDD1.n147 VDD1.n124 171.744
R2061 VDD1.n154 VDD1.n124 171.744
R2062 VDD1.n155 VDD1.n154 171.744
R2063 VDD1.n155 VDD1.n120 171.744
R2064 VDD1.n162 VDD1.n120 171.744
R2065 VDD1.n163 VDD1.n162 171.744
R2066 VDD1.n163 VDD1.n116 171.744
R2067 VDD1.n170 VDD1.n116 171.744
R2068 VDD1.n171 VDD1.n170 171.744
R2069 VDD1.n171 VDD1.n112 171.744
R2070 VDD1.n179 VDD1.n112 171.744
R2071 VDD1.n180 VDD1.n179 171.744
R2072 VDD1.n181 VDD1.n180 171.744
R2073 VDD1.n181 VDD1.n108 171.744
R2074 VDD1.n188 VDD1.n108 171.744
R2075 VDD1.n189 VDD1.n188 171.744
R2076 VDD1.n189 VDD1.n104 171.744
R2077 VDD1.n196 VDD1.n104 171.744
R2078 VDD1.n197 VDD1.n196 171.744
R2079 VDD1 VDD1.n201 90.4151
R2080 VDD1.t1 VDD1.n32 85.8723
R2081 VDD1.t0 VDD1.n132 85.8723
R2082 VDD1 VDD1.n100 47.0476
R2083 VDD1.n34 VDD1.n33 16.3895
R2084 VDD1.n134 VDD1.n133 16.3895
R2085 VDD1.n81 VDD1.n10 13.1884
R2086 VDD1.n182 VDD1.n111 13.1884
R2087 VDD1.n82 VDD1.n8 12.8005
R2088 VDD1.n77 VDD1.n12 12.8005
R2089 VDD1.n37 VDD1.n36 12.8005
R2090 VDD1.n137 VDD1.n136 12.8005
R2091 VDD1.n178 VDD1.n177 12.8005
R2092 VDD1.n183 VDD1.n109 12.8005
R2093 VDD1.n86 VDD1.n85 12.0247
R2094 VDD1.n76 VDD1.n13 12.0247
R2095 VDD1.n40 VDD1.n31 12.0247
R2096 VDD1.n140 VDD1.n131 12.0247
R2097 VDD1.n176 VDD1.n113 12.0247
R2098 VDD1.n187 VDD1.n186 12.0247
R2099 VDD1.n89 VDD1.n6 11.249
R2100 VDD1.n73 VDD1.n72 11.249
R2101 VDD1.n41 VDD1.n29 11.249
R2102 VDD1.n141 VDD1.n129 11.249
R2103 VDD1.n173 VDD1.n172 11.249
R2104 VDD1.n190 VDD1.n107 11.249
R2105 VDD1.n90 VDD1.n4 10.4732
R2106 VDD1.n69 VDD1.n15 10.4732
R2107 VDD1.n45 VDD1.n44 10.4732
R2108 VDD1.n145 VDD1.n144 10.4732
R2109 VDD1.n169 VDD1.n115 10.4732
R2110 VDD1.n191 VDD1.n105 10.4732
R2111 VDD1.n94 VDD1.n93 9.69747
R2112 VDD1.n68 VDD1.n17 9.69747
R2113 VDD1.n48 VDD1.n27 9.69747
R2114 VDD1.n148 VDD1.n127 9.69747
R2115 VDD1.n168 VDD1.n117 9.69747
R2116 VDD1.n195 VDD1.n194 9.69747
R2117 VDD1.n100 VDD1.n99 9.45567
R2118 VDD1.n201 VDD1.n200 9.45567
R2119 VDD1.n60 VDD1.n59 9.3005
R2120 VDD1.n19 VDD1.n18 9.3005
R2121 VDD1.n66 VDD1.n65 9.3005
R2122 VDD1.n68 VDD1.n67 9.3005
R2123 VDD1.n15 VDD1.n14 9.3005
R2124 VDD1.n74 VDD1.n73 9.3005
R2125 VDD1.n76 VDD1.n75 9.3005
R2126 VDD1.n12 VDD1.n9 9.3005
R2127 VDD1.n99 VDD1.n98 9.3005
R2128 VDD1.n2 VDD1.n1 9.3005
R2129 VDD1.n93 VDD1.n92 9.3005
R2130 VDD1.n91 VDD1.n90 9.3005
R2131 VDD1.n6 VDD1.n5 9.3005
R2132 VDD1.n85 VDD1.n84 9.3005
R2133 VDD1.n83 VDD1.n82 9.3005
R2134 VDD1.n58 VDD1.n57 9.3005
R2135 VDD1.n23 VDD1.n22 9.3005
R2136 VDD1.n52 VDD1.n51 9.3005
R2137 VDD1.n50 VDD1.n49 9.3005
R2138 VDD1.n27 VDD1.n26 9.3005
R2139 VDD1.n44 VDD1.n43 9.3005
R2140 VDD1.n42 VDD1.n41 9.3005
R2141 VDD1.n31 VDD1.n30 9.3005
R2142 VDD1.n36 VDD1.n35 9.3005
R2143 VDD1.n200 VDD1.n199 9.3005
R2144 VDD1.n103 VDD1.n102 9.3005
R2145 VDD1.n194 VDD1.n193 9.3005
R2146 VDD1.n192 VDD1.n191 9.3005
R2147 VDD1.n107 VDD1.n106 9.3005
R2148 VDD1.n186 VDD1.n185 9.3005
R2149 VDD1.n184 VDD1.n183 9.3005
R2150 VDD1.n123 VDD1.n122 9.3005
R2151 VDD1.n152 VDD1.n151 9.3005
R2152 VDD1.n150 VDD1.n149 9.3005
R2153 VDD1.n127 VDD1.n126 9.3005
R2154 VDD1.n144 VDD1.n143 9.3005
R2155 VDD1.n142 VDD1.n141 9.3005
R2156 VDD1.n131 VDD1.n130 9.3005
R2157 VDD1.n136 VDD1.n135 9.3005
R2158 VDD1.n158 VDD1.n157 9.3005
R2159 VDD1.n160 VDD1.n159 9.3005
R2160 VDD1.n119 VDD1.n118 9.3005
R2161 VDD1.n166 VDD1.n165 9.3005
R2162 VDD1.n168 VDD1.n167 9.3005
R2163 VDD1.n115 VDD1.n114 9.3005
R2164 VDD1.n174 VDD1.n173 9.3005
R2165 VDD1.n176 VDD1.n175 9.3005
R2166 VDD1.n177 VDD1.n110 9.3005
R2167 VDD1.n97 VDD1.n2 8.92171
R2168 VDD1.n65 VDD1.n64 8.92171
R2169 VDD1.n49 VDD1.n25 8.92171
R2170 VDD1.n149 VDD1.n125 8.92171
R2171 VDD1.n165 VDD1.n164 8.92171
R2172 VDD1.n198 VDD1.n103 8.92171
R2173 VDD1.n98 VDD1.n0 8.14595
R2174 VDD1.n61 VDD1.n19 8.14595
R2175 VDD1.n53 VDD1.n52 8.14595
R2176 VDD1.n153 VDD1.n152 8.14595
R2177 VDD1.n161 VDD1.n119 8.14595
R2178 VDD1.n199 VDD1.n101 8.14595
R2179 VDD1.n60 VDD1.n21 7.3702
R2180 VDD1.n56 VDD1.n23 7.3702
R2181 VDD1.n156 VDD1.n123 7.3702
R2182 VDD1.n160 VDD1.n121 7.3702
R2183 VDD1.n57 VDD1.n21 6.59444
R2184 VDD1.n57 VDD1.n56 6.59444
R2185 VDD1.n157 VDD1.n156 6.59444
R2186 VDD1.n157 VDD1.n121 6.59444
R2187 VDD1.n100 VDD1.n0 5.81868
R2188 VDD1.n61 VDD1.n60 5.81868
R2189 VDD1.n53 VDD1.n23 5.81868
R2190 VDD1.n153 VDD1.n123 5.81868
R2191 VDD1.n161 VDD1.n160 5.81868
R2192 VDD1.n201 VDD1.n101 5.81868
R2193 VDD1.n98 VDD1.n97 5.04292
R2194 VDD1.n64 VDD1.n19 5.04292
R2195 VDD1.n52 VDD1.n25 5.04292
R2196 VDD1.n152 VDD1.n125 5.04292
R2197 VDD1.n164 VDD1.n119 5.04292
R2198 VDD1.n199 VDD1.n198 5.04292
R2199 VDD1.n94 VDD1.n2 4.26717
R2200 VDD1.n65 VDD1.n17 4.26717
R2201 VDD1.n49 VDD1.n48 4.26717
R2202 VDD1.n149 VDD1.n148 4.26717
R2203 VDD1.n165 VDD1.n117 4.26717
R2204 VDD1.n195 VDD1.n103 4.26717
R2205 VDD1.n35 VDD1.n34 3.70982
R2206 VDD1.n135 VDD1.n134 3.70982
R2207 VDD1.n93 VDD1.n4 3.49141
R2208 VDD1.n69 VDD1.n68 3.49141
R2209 VDD1.n45 VDD1.n27 3.49141
R2210 VDD1.n145 VDD1.n127 3.49141
R2211 VDD1.n169 VDD1.n168 3.49141
R2212 VDD1.n194 VDD1.n105 3.49141
R2213 VDD1.n90 VDD1.n89 2.71565
R2214 VDD1.n72 VDD1.n15 2.71565
R2215 VDD1.n44 VDD1.n29 2.71565
R2216 VDD1.n144 VDD1.n129 2.71565
R2217 VDD1.n172 VDD1.n115 2.71565
R2218 VDD1.n191 VDD1.n190 2.71565
R2219 VDD1.n86 VDD1.n6 1.93989
R2220 VDD1.n73 VDD1.n13 1.93989
R2221 VDD1.n41 VDD1.n40 1.93989
R2222 VDD1.n141 VDD1.n140 1.93989
R2223 VDD1.n173 VDD1.n113 1.93989
R2224 VDD1.n187 VDD1.n107 1.93989
R2225 VDD1.n85 VDD1.n8 1.16414
R2226 VDD1.n77 VDD1.n76 1.16414
R2227 VDD1.n37 VDD1.n31 1.16414
R2228 VDD1.n137 VDD1.n131 1.16414
R2229 VDD1.n178 VDD1.n176 1.16414
R2230 VDD1.n186 VDD1.n109 1.16414
R2231 VDD1.n82 VDD1.n81 0.388379
R2232 VDD1.n12 VDD1.n10 0.388379
R2233 VDD1.n36 VDD1.n33 0.388379
R2234 VDD1.n136 VDD1.n133 0.388379
R2235 VDD1.n177 VDD1.n111 0.388379
R2236 VDD1.n183 VDD1.n182 0.388379
R2237 VDD1.n99 VDD1.n1 0.155672
R2238 VDD1.n92 VDD1.n1 0.155672
R2239 VDD1.n92 VDD1.n91 0.155672
R2240 VDD1.n91 VDD1.n5 0.155672
R2241 VDD1.n84 VDD1.n5 0.155672
R2242 VDD1.n84 VDD1.n83 0.155672
R2243 VDD1.n83 VDD1.n9 0.155672
R2244 VDD1.n75 VDD1.n9 0.155672
R2245 VDD1.n75 VDD1.n74 0.155672
R2246 VDD1.n74 VDD1.n14 0.155672
R2247 VDD1.n67 VDD1.n14 0.155672
R2248 VDD1.n67 VDD1.n66 0.155672
R2249 VDD1.n66 VDD1.n18 0.155672
R2250 VDD1.n59 VDD1.n18 0.155672
R2251 VDD1.n59 VDD1.n58 0.155672
R2252 VDD1.n58 VDD1.n22 0.155672
R2253 VDD1.n51 VDD1.n22 0.155672
R2254 VDD1.n51 VDD1.n50 0.155672
R2255 VDD1.n50 VDD1.n26 0.155672
R2256 VDD1.n43 VDD1.n26 0.155672
R2257 VDD1.n43 VDD1.n42 0.155672
R2258 VDD1.n42 VDD1.n30 0.155672
R2259 VDD1.n35 VDD1.n30 0.155672
R2260 VDD1.n135 VDD1.n130 0.155672
R2261 VDD1.n142 VDD1.n130 0.155672
R2262 VDD1.n143 VDD1.n142 0.155672
R2263 VDD1.n143 VDD1.n126 0.155672
R2264 VDD1.n150 VDD1.n126 0.155672
R2265 VDD1.n151 VDD1.n150 0.155672
R2266 VDD1.n151 VDD1.n122 0.155672
R2267 VDD1.n158 VDD1.n122 0.155672
R2268 VDD1.n159 VDD1.n158 0.155672
R2269 VDD1.n159 VDD1.n118 0.155672
R2270 VDD1.n166 VDD1.n118 0.155672
R2271 VDD1.n167 VDD1.n166 0.155672
R2272 VDD1.n167 VDD1.n114 0.155672
R2273 VDD1.n174 VDD1.n114 0.155672
R2274 VDD1.n175 VDD1.n174 0.155672
R2275 VDD1.n175 VDD1.n110 0.155672
R2276 VDD1.n184 VDD1.n110 0.155672
R2277 VDD1.n185 VDD1.n184 0.155672
R2278 VDD1.n185 VDD1.n106 0.155672
R2279 VDD1.n192 VDD1.n106 0.155672
R2280 VDD1.n193 VDD1.n192 0.155672
R2281 VDD1.n193 VDD1.n102 0.155672
R2282 VDD1.n200 VDD1.n102 0.155672
C0 w_n1810_n4592# VN 2.54456f
C1 VTAIL VDD1 6.77297f
C2 VTAIL VDD2 6.81487f
C3 VN VTAIL 3.13244f
C4 B VP 1.35734f
C5 w_n1810_n4592# VTAIL 3.68712f
C6 VDD1 VP 3.93821f
C7 VDD2 VP 0.299245f
C8 VN VP 6.19832f
C9 w_n1810_n4592# VP 2.77332f
C10 VDD1 B 2.06091f
C11 VDD2 B 2.08365f
C12 VTAIL VP 3.14695f
C13 VN B 0.984563f
C14 VDD1 VDD2 0.577762f
C15 w_n1810_n4592# B 9.62801f
C16 VN VDD1 0.148075f
C17 w_n1810_n4592# VDD1 2.12181f
C18 VN VDD2 3.79152f
C19 VTAIL B 4.56869f
C20 w_n1810_n4592# VDD2 2.13771f
C21 VDD2 VSUBS 1.054582f
C22 VDD1 VSUBS 5.207261f
C23 VTAIL VSUBS 1.14316f
C24 VN VSUBS 9.04443f
C25 VP VSUBS 1.667394f
C26 B VSUBS 3.797498f
C27 w_n1810_n4592# VSUBS 0.101628p
C28 VDD1.n0 VSUBS 0.029038f
C29 VDD1.n1 VSUBS 0.027821f
C30 VDD1.n2 VSUBS 0.01495f
C31 VDD1.n3 VSUBS 0.035336f
C32 VDD1.n4 VSUBS 0.015829f
C33 VDD1.n5 VSUBS 0.027821f
C34 VDD1.n6 VSUBS 0.01495f
C35 VDD1.n7 VSUBS 0.035336f
C36 VDD1.n8 VSUBS 0.015829f
C37 VDD1.n9 VSUBS 0.027821f
C38 VDD1.n10 VSUBS 0.01539f
C39 VDD1.n11 VSUBS 0.035336f
C40 VDD1.n12 VSUBS 0.01495f
C41 VDD1.n13 VSUBS 0.015829f
C42 VDD1.n14 VSUBS 0.027821f
C43 VDD1.n15 VSUBS 0.01495f
C44 VDD1.n16 VSUBS 0.035336f
C45 VDD1.n17 VSUBS 0.015829f
C46 VDD1.n18 VSUBS 0.027821f
C47 VDD1.n19 VSUBS 0.01495f
C48 VDD1.n20 VSUBS 0.035336f
C49 VDD1.n21 VSUBS 0.015829f
C50 VDD1.n22 VSUBS 0.027821f
C51 VDD1.n23 VSUBS 0.01495f
C52 VDD1.n24 VSUBS 0.035336f
C53 VDD1.n25 VSUBS 0.015829f
C54 VDD1.n26 VSUBS 0.027821f
C55 VDD1.n27 VSUBS 0.01495f
C56 VDD1.n28 VSUBS 0.035336f
C57 VDD1.n29 VSUBS 0.015829f
C58 VDD1.n30 VSUBS 0.027821f
C59 VDD1.n31 VSUBS 0.01495f
C60 VDD1.n32 VSUBS 0.026502f
C61 VDD1.n33 VSUBS 0.022479f
C62 VDD1.t1 VSUBS 0.075863f
C63 VDD1.n34 VSUBS 0.221717f
C64 VDD1.n35 VSUBS 2.17049f
C65 VDD1.n36 VSUBS 0.01495f
C66 VDD1.n37 VSUBS 0.015829f
C67 VDD1.n38 VSUBS 0.035336f
C68 VDD1.n39 VSUBS 0.035336f
C69 VDD1.n40 VSUBS 0.015829f
C70 VDD1.n41 VSUBS 0.01495f
C71 VDD1.n42 VSUBS 0.027821f
C72 VDD1.n43 VSUBS 0.027821f
C73 VDD1.n44 VSUBS 0.01495f
C74 VDD1.n45 VSUBS 0.015829f
C75 VDD1.n46 VSUBS 0.035336f
C76 VDD1.n47 VSUBS 0.035336f
C77 VDD1.n48 VSUBS 0.015829f
C78 VDD1.n49 VSUBS 0.01495f
C79 VDD1.n50 VSUBS 0.027821f
C80 VDD1.n51 VSUBS 0.027821f
C81 VDD1.n52 VSUBS 0.01495f
C82 VDD1.n53 VSUBS 0.015829f
C83 VDD1.n54 VSUBS 0.035336f
C84 VDD1.n55 VSUBS 0.035336f
C85 VDD1.n56 VSUBS 0.015829f
C86 VDD1.n57 VSUBS 0.01495f
C87 VDD1.n58 VSUBS 0.027821f
C88 VDD1.n59 VSUBS 0.027821f
C89 VDD1.n60 VSUBS 0.01495f
C90 VDD1.n61 VSUBS 0.015829f
C91 VDD1.n62 VSUBS 0.035336f
C92 VDD1.n63 VSUBS 0.035336f
C93 VDD1.n64 VSUBS 0.015829f
C94 VDD1.n65 VSUBS 0.01495f
C95 VDD1.n66 VSUBS 0.027821f
C96 VDD1.n67 VSUBS 0.027821f
C97 VDD1.n68 VSUBS 0.01495f
C98 VDD1.n69 VSUBS 0.015829f
C99 VDD1.n70 VSUBS 0.035336f
C100 VDD1.n71 VSUBS 0.035336f
C101 VDD1.n72 VSUBS 0.015829f
C102 VDD1.n73 VSUBS 0.01495f
C103 VDD1.n74 VSUBS 0.027821f
C104 VDD1.n75 VSUBS 0.027821f
C105 VDD1.n76 VSUBS 0.01495f
C106 VDD1.n77 VSUBS 0.015829f
C107 VDD1.n78 VSUBS 0.035336f
C108 VDD1.n79 VSUBS 0.035336f
C109 VDD1.n80 VSUBS 0.035336f
C110 VDD1.n81 VSUBS 0.01539f
C111 VDD1.n82 VSUBS 0.01495f
C112 VDD1.n83 VSUBS 0.027821f
C113 VDD1.n84 VSUBS 0.027821f
C114 VDD1.n85 VSUBS 0.01495f
C115 VDD1.n86 VSUBS 0.015829f
C116 VDD1.n87 VSUBS 0.035336f
C117 VDD1.n88 VSUBS 0.035336f
C118 VDD1.n89 VSUBS 0.015829f
C119 VDD1.n90 VSUBS 0.01495f
C120 VDD1.n91 VSUBS 0.027821f
C121 VDD1.n92 VSUBS 0.027821f
C122 VDD1.n93 VSUBS 0.01495f
C123 VDD1.n94 VSUBS 0.015829f
C124 VDD1.n95 VSUBS 0.035336f
C125 VDD1.n96 VSUBS 0.080328f
C126 VDD1.n97 VSUBS 0.015829f
C127 VDD1.n98 VSUBS 0.01495f
C128 VDD1.n99 VSUBS 0.059746f
C129 VDD1.n100 VSUBS 0.060319f
C130 VDD1.n101 VSUBS 0.029038f
C131 VDD1.n102 VSUBS 0.027821f
C132 VDD1.n103 VSUBS 0.01495f
C133 VDD1.n104 VSUBS 0.035336f
C134 VDD1.n105 VSUBS 0.015829f
C135 VDD1.n106 VSUBS 0.027821f
C136 VDD1.n107 VSUBS 0.01495f
C137 VDD1.n108 VSUBS 0.035336f
C138 VDD1.n109 VSUBS 0.015829f
C139 VDD1.n110 VSUBS 0.027821f
C140 VDD1.n111 VSUBS 0.01539f
C141 VDD1.n112 VSUBS 0.035336f
C142 VDD1.n113 VSUBS 0.015829f
C143 VDD1.n114 VSUBS 0.027821f
C144 VDD1.n115 VSUBS 0.01495f
C145 VDD1.n116 VSUBS 0.035336f
C146 VDD1.n117 VSUBS 0.015829f
C147 VDD1.n118 VSUBS 0.027821f
C148 VDD1.n119 VSUBS 0.01495f
C149 VDD1.n120 VSUBS 0.035336f
C150 VDD1.n121 VSUBS 0.015829f
C151 VDD1.n122 VSUBS 0.027821f
C152 VDD1.n123 VSUBS 0.01495f
C153 VDD1.n124 VSUBS 0.035336f
C154 VDD1.n125 VSUBS 0.015829f
C155 VDD1.n126 VSUBS 0.027821f
C156 VDD1.n127 VSUBS 0.01495f
C157 VDD1.n128 VSUBS 0.035336f
C158 VDD1.n129 VSUBS 0.015829f
C159 VDD1.n130 VSUBS 0.027821f
C160 VDD1.n131 VSUBS 0.01495f
C161 VDD1.n132 VSUBS 0.026502f
C162 VDD1.n133 VSUBS 0.022479f
C163 VDD1.t0 VSUBS 0.075863f
C164 VDD1.n134 VSUBS 0.221717f
C165 VDD1.n135 VSUBS 2.17049f
C166 VDD1.n136 VSUBS 0.01495f
C167 VDD1.n137 VSUBS 0.015829f
C168 VDD1.n138 VSUBS 0.035336f
C169 VDD1.n139 VSUBS 0.035336f
C170 VDD1.n140 VSUBS 0.015829f
C171 VDD1.n141 VSUBS 0.01495f
C172 VDD1.n142 VSUBS 0.027821f
C173 VDD1.n143 VSUBS 0.027821f
C174 VDD1.n144 VSUBS 0.01495f
C175 VDD1.n145 VSUBS 0.015829f
C176 VDD1.n146 VSUBS 0.035336f
C177 VDD1.n147 VSUBS 0.035336f
C178 VDD1.n148 VSUBS 0.015829f
C179 VDD1.n149 VSUBS 0.01495f
C180 VDD1.n150 VSUBS 0.027821f
C181 VDD1.n151 VSUBS 0.027821f
C182 VDD1.n152 VSUBS 0.01495f
C183 VDD1.n153 VSUBS 0.015829f
C184 VDD1.n154 VSUBS 0.035336f
C185 VDD1.n155 VSUBS 0.035336f
C186 VDD1.n156 VSUBS 0.015829f
C187 VDD1.n157 VSUBS 0.01495f
C188 VDD1.n158 VSUBS 0.027821f
C189 VDD1.n159 VSUBS 0.027821f
C190 VDD1.n160 VSUBS 0.01495f
C191 VDD1.n161 VSUBS 0.015829f
C192 VDD1.n162 VSUBS 0.035336f
C193 VDD1.n163 VSUBS 0.035336f
C194 VDD1.n164 VSUBS 0.015829f
C195 VDD1.n165 VSUBS 0.01495f
C196 VDD1.n166 VSUBS 0.027821f
C197 VDD1.n167 VSUBS 0.027821f
C198 VDD1.n168 VSUBS 0.01495f
C199 VDD1.n169 VSUBS 0.015829f
C200 VDD1.n170 VSUBS 0.035336f
C201 VDD1.n171 VSUBS 0.035336f
C202 VDD1.n172 VSUBS 0.015829f
C203 VDD1.n173 VSUBS 0.01495f
C204 VDD1.n174 VSUBS 0.027821f
C205 VDD1.n175 VSUBS 0.027821f
C206 VDD1.n176 VSUBS 0.01495f
C207 VDD1.n177 VSUBS 0.01495f
C208 VDD1.n178 VSUBS 0.015829f
C209 VDD1.n179 VSUBS 0.035336f
C210 VDD1.n180 VSUBS 0.035336f
C211 VDD1.n181 VSUBS 0.035336f
C212 VDD1.n182 VSUBS 0.01539f
C213 VDD1.n183 VSUBS 0.01495f
C214 VDD1.n184 VSUBS 0.027821f
C215 VDD1.n185 VSUBS 0.027821f
C216 VDD1.n186 VSUBS 0.01495f
C217 VDD1.n187 VSUBS 0.015829f
C218 VDD1.n188 VSUBS 0.035336f
C219 VDD1.n189 VSUBS 0.035336f
C220 VDD1.n190 VSUBS 0.015829f
C221 VDD1.n191 VSUBS 0.01495f
C222 VDD1.n192 VSUBS 0.027821f
C223 VDD1.n193 VSUBS 0.027821f
C224 VDD1.n194 VSUBS 0.01495f
C225 VDD1.n195 VSUBS 0.015829f
C226 VDD1.n196 VSUBS 0.035336f
C227 VDD1.n197 VSUBS 0.080328f
C228 VDD1.n198 VSUBS 0.015829f
C229 VDD1.n199 VSUBS 0.01495f
C230 VDD1.n200 VSUBS 0.059746f
C231 VDD1.n201 VSUBS 1.08006f
C232 VP.t0 VSUBS 4.80713f
C233 VP.t1 VSUBS 4.31779f
C234 VP.n0 VSUBS 6.80711f
C235 VDD2.n0 VSUBS 0.029043f
C236 VDD2.n1 VSUBS 0.027826f
C237 VDD2.n2 VSUBS 0.014953f
C238 VDD2.n3 VSUBS 0.035343f
C239 VDD2.n4 VSUBS 0.015832f
C240 VDD2.n5 VSUBS 0.027826f
C241 VDD2.n6 VSUBS 0.014953f
C242 VDD2.n7 VSUBS 0.035343f
C243 VDD2.n8 VSUBS 0.015832f
C244 VDD2.n9 VSUBS 0.027826f
C245 VDD2.n10 VSUBS 0.015392f
C246 VDD2.n11 VSUBS 0.035343f
C247 VDD2.n12 VSUBS 0.015832f
C248 VDD2.n13 VSUBS 0.027826f
C249 VDD2.n14 VSUBS 0.014953f
C250 VDD2.n15 VSUBS 0.035343f
C251 VDD2.n16 VSUBS 0.015832f
C252 VDD2.n17 VSUBS 0.027826f
C253 VDD2.n18 VSUBS 0.014953f
C254 VDD2.n19 VSUBS 0.035343f
C255 VDD2.n20 VSUBS 0.015832f
C256 VDD2.n21 VSUBS 0.027826f
C257 VDD2.n22 VSUBS 0.014953f
C258 VDD2.n23 VSUBS 0.035343f
C259 VDD2.n24 VSUBS 0.015832f
C260 VDD2.n25 VSUBS 0.027826f
C261 VDD2.n26 VSUBS 0.014953f
C262 VDD2.n27 VSUBS 0.035343f
C263 VDD2.n28 VSUBS 0.015832f
C264 VDD2.n29 VSUBS 0.027826f
C265 VDD2.n30 VSUBS 0.014953f
C266 VDD2.n31 VSUBS 0.026507f
C267 VDD2.n32 VSUBS 0.022483f
C268 VDD2.t0 VSUBS 0.075877f
C269 VDD2.n33 VSUBS 0.221758f
C270 VDD2.n34 VSUBS 2.17089f
C271 VDD2.n35 VSUBS 0.014953f
C272 VDD2.n36 VSUBS 0.015832f
C273 VDD2.n37 VSUBS 0.035343f
C274 VDD2.n38 VSUBS 0.035343f
C275 VDD2.n39 VSUBS 0.015832f
C276 VDD2.n40 VSUBS 0.014953f
C277 VDD2.n41 VSUBS 0.027826f
C278 VDD2.n42 VSUBS 0.027826f
C279 VDD2.n43 VSUBS 0.014953f
C280 VDD2.n44 VSUBS 0.015832f
C281 VDD2.n45 VSUBS 0.035343f
C282 VDD2.n46 VSUBS 0.035343f
C283 VDD2.n47 VSUBS 0.015832f
C284 VDD2.n48 VSUBS 0.014953f
C285 VDD2.n49 VSUBS 0.027826f
C286 VDD2.n50 VSUBS 0.027826f
C287 VDD2.n51 VSUBS 0.014953f
C288 VDD2.n52 VSUBS 0.015832f
C289 VDD2.n53 VSUBS 0.035343f
C290 VDD2.n54 VSUBS 0.035343f
C291 VDD2.n55 VSUBS 0.015832f
C292 VDD2.n56 VSUBS 0.014953f
C293 VDD2.n57 VSUBS 0.027826f
C294 VDD2.n58 VSUBS 0.027826f
C295 VDD2.n59 VSUBS 0.014953f
C296 VDD2.n60 VSUBS 0.015832f
C297 VDD2.n61 VSUBS 0.035343f
C298 VDD2.n62 VSUBS 0.035343f
C299 VDD2.n63 VSUBS 0.015832f
C300 VDD2.n64 VSUBS 0.014953f
C301 VDD2.n65 VSUBS 0.027826f
C302 VDD2.n66 VSUBS 0.027826f
C303 VDD2.n67 VSUBS 0.014953f
C304 VDD2.n68 VSUBS 0.015832f
C305 VDD2.n69 VSUBS 0.035343f
C306 VDD2.n70 VSUBS 0.035343f
C307 VDD2.n71 VSUBS 0.015832f
C308 VDD2.n72 VSUBS 0.014953f
C309 VDD2.n73 VSUBS 0.027826f
C310 VDD2.n74 VSUBS 0.027826f
C311 VDD2.n75 VSUBS 0.014953f
C312 VDD2.n76 VSUBS 0.014953f
C313 VDD2.n77 VSUBS 0.015832f
C314 VDD2.n78 VSUBS 0.035343f
C315 VDD2.n79 VSUBS 0.035343f
C316 VDD2.n80 VSUBS 0.035343f
C317 VDD2.n81 VSUBS 0.015392f
C318 VDD2.n82 VSUBS 0.014953f
C319 VDD2.n83 VSUBS 0.027826f
C320 VDD2.n84 VSUBS 0.027826f
C321 VDD2.n85 VSUBS 0.014953f
C322 VDD2.n86 VSUBS 0.015832f
C323 VDD2.n87 VSUBS 0.035343f
C324 VDD2.n88 VSUBS 0.035343f
C325 VDD2.n89 VSUBS 0.015832f
C326 VDD2.n90 VSUBS 0.014953f
C327 VDD2.n91 VSUBS 0.027826f
C328 VDD2.n92 VSUBS 0.027826f
C329 VDD2.n93 VSUBS 0.014953f
C330 VDD2.n94 VSUBS 0.015832f
C331 VDD2.n95 VSUBS 0.035343f
C332 VDD2.n96 VSUBS 0.080343f
C333 VDD2.n97 VSUBS 0.015832f
C334 VDD2.n98 VSUBS 0.014953f
C335 VDD2.n99 VSUBS 0.059758f
C336 VDD2.n100 VSUBS 1.02796f
C337 VDD2.n101 VSUBS 0.029043f
C338 VDD2.n102 VSUBS 0.027826f
C339 VDD2.n103 VSUBS 0.014953f
C340 VDD2.n104 VSUBS 0.035343f
C341 VDD2.n105 VSUBS 0.015832f
C342 VDD2.n106 VSUBS 0.027826f
C343 VDD2.n107 VSUBS 0.014953f
C344 VDD2.n108 VSUBS 0.035343f
C345 VDD2.n109 VSUBS 0.015832f
C346 VDD2.n110 VSUBS 0.027826f
C347 VDD2.n111 VSUBS 0.015392f
C348 VDD2.n112 VSUBS 0.035343f
C349 VDD2.n113 VSUBS 0.014953f
C350 VDD2.n114 VSUBS 0.015832f
C351 VDD2.n115 VSUBS 0.027826f
C352 VDD2.n116 VSUBS 0.014953f
C353 VDD2.n117 VSUBS 0.035343f
C354 VDD2.n118 VSUBS 0.015832f
C355 VDD2.n119 VSUBS 0.027826f
C356 VDD2.n120 VSUBS 0.014953f
C357 VDD2.n121 VSUBS 0.035343f
C358 VDD2.n122 VSUBS 0.015832f
C359 VDD2.n123 VSUBS 0.027826f
C360 VDD2.n124 VSUBS 0.014953f
C361 VDD2.n125 VSUBS 0.035343f
C362 VDD2.n126 VSUBS 0.015832f
C363 VDD2.n127 VSUBS 0.027826f
C364 VDD2.n128 VSUBS 0.014953f
C365 VDD2.n129 VSUBS 0.035343f
C366 VDD2.n130 VSUBS 0.015832f
C367 VDD2.n131 VSUBS 0.027826f
C368 VDD2.n132 VSUBS 0.014953f
C369 VDD2.n133 VSUBS 0.026507f
C370 VDD2.n134 VSUBS 0.022483f
C371 VDD2.t1 VSUBS 0.075877f
C372 VDD2.n135 VSUBS 0.221758f
C373 VDD2.n136 VSUBS 2.17089f
C374 VDD2.n137 VSUBS 0.014953f
C375 VDD2.n138 VSUBS 0.015832f
C376 VDD2.n139 VSUBS 0.035343f
C377 VDD2.n140 VSUBS 0.035343f
C378 VDD2.n141 VSUBS 0.015832f
C379 VDD2.n142 VSUBS 0.014953f
C380 VDD2.n143 VSUBS 0.027826f
C381 VDD2.n144 VSUBS 0.027826f
C382 VDD2.n145 VSUBS 0.014953f
C383 VDD2.n146 VSUBS 0.015832f
C384 VDD2.n147 VSUBS 0.035343f
C385 VDD2.n148 VSUBS 0.035343f
C386 VDD2.n149 VSUBS 0.015832f
C387 VDD2.n150 VSUBS 0.014953f
C388 VDD2.n151 VSUBS 0.027826f
C389 VDD2.n152 VSUBS 0.027826f
C390 VDD2.n153 VSUBS 0.014953f
C391 VDD2.n154 VSUBS 0.015832f
C392 VDD2.n155 VSUBS 0.035343f
C393 VDD2.n156 VSUBS 0.035343f
C394 VDD2.n157 VSUBS 0.015832f
C395 VDD2.n158 VSUBS 0.014953f
C396 VDD2.n159 VSUBS 0.027826f
C397 VDD2.n160 VSUBS 0.027826f
C398 VDD2.n161 VSUBS 0.014953f
C399 VDD2.n162 VSUBS 0.015832f
C400 VDD2.n163 VSUBS 0.035343f
C401 VDD2.n164 VSUBS 0.035343f
C402 VDD2.n165 VSUBS 0.015832f
C403 VDD2.n166 VSUBS 0.014953f
C404 VDD2.n167 VSUBS 0.027826f
C405 VDD2.n168 VSUBS 0.027826f
C406 VDD2.n169 VSUBS 0.014953f
C407 VDD2.n170 VSUBS 0.015832f
C408 VDD2.n171 VSUBS 0.035343f
C409 VDD2.n172 VSUBS 0.035343f
C410 VDD2.n173 VSUBS 0.015832f
C411 VDD2.n174 VSUBS 0.014953f
C412 VDD2.n175 VSUBS 0.027826f
C413 VDD2.n176 VSUBS 0.027826f
C414 VDD2.n177 VSUBS 0.014953f
C415 VDD2.n178 VSUBS 0.015832f
C416 VDD2.n179 VSUBS 0.035343f
C417 VDD2.n180 VSUBS 0.035343f
C418 VDD2.n181 VSUBS 0.035343f
C419 VDD2.n182 VSUBS 0.015392f
C420 VDD2.n183 VSUBS 0.014953f
C421 VDD2.n184 VSUBS 0.027826f
C422 VDD2.n185 VSUBS 0.027826f
C423 VDD2.n186 VSUBS 0.014953f
C424 VDD2.n187 VSUBS 0.015832f
C425 VDD2.n188 VSUBS 0.035343f
C426 VDD2.n189 VSUBS 0.035343f
C427 VDD2.n190 VSUBS 0.015832f
C428 VDD2.n191 VSUBS 0.014953f
C429 VDD2.n192 VSUBS 0.027826f
C430 VDD2.n193 VSUBS 0.027826f
C431 VDD2.n194 VSUBS 0.014953f
C432 VDD2.n195 VSUBS 0.015832f
C433 VDD2.n196 VSUBS 0.035343f
C434 VDD2.n197 VSUBS 0.080343f
C435 VDD2.n198 VSUBS 0.015832f
C436 VDD2.n199 VSUBS 0.014953f
C437 VDD2.n200 VSUBS 0.059758f
C438 VDD2.n201 VSUBS 0.05928f
C439 VDD2.n202 VSUBS 3.88568f
C440 VTAIL.n0 VSUBS 0.028915f
C441 VTAIL.n1 VSUBS 0.027703f
C442 VTAIL.n2 VSUBS 0.014886f
C443 VTAIL.n3 VSUBS 0.035186f
C444 VTAIL.n4 VSUBS 0.015762f
C445 VTAIL.n5 VSUBS 0.027703f
C446 VTAIL.n6 VSUBS 0.014886f
C447 VTAIL.n7 VSUBS 0.035186f
C448 VTAIL.n8 VSUBS 0.015762f
C449 VTAIL.n9 VSUBS 0.027703f
C450 VTAIL.n10 VSUBS 0.015324f
C451 VTAIL.n11 VSUBS 0.035186f
C452 VTAIL.n12 VSUBS 0.015762f
C453 VTAIL.n13 VSUBS 0.027703f
C454 VTAIL.n14 VSUBS 0.014886f
C455 VTAIL.n15 VSUBS 0.035186f
C456 VTAIL.n16 VSUBS 0.015762f
C457 VTAIL.n17 VSUBS 0.027703f
C458 VTAIL.n18 VSUBS 0.014886f
C459 VTAIL.n19 VSUBS 0.035186f
C460 VTAIL.n20 VSUBS 0.015762f
C461 VTAIL.n21 VSUBS 0.027703f
C462 VTAIL.n22 VSUBS 0.014886f
C463 VTAIL.n23 VSUBS 0.035186f
C464 VTAIL.n24 VSUBS 0.015762f
C465 VTAIL.n25 VSUBS 0.027703f
C466 VTAIL.n26 VSUBS 0.014886f
C467 VTAIL.n27 VSUBS 0.035186f
C468 VTAIL.n28 VSUBS 0.015762f
C469 VTAIL.n29 VSUBS 0.027703f
C470 VTAIL.n30 VSUBS 0.014886f
C471 VTAIL.n31 VSUBS 0.02639f
C472 VTAIL.n32 VSUBS 0.022384f
C473 VTAIL.t0 VSUBS 0.075541f
C474 VTAIL.n33 VSUBS 0.220777f
C475 VTAIL.n34 VSUBS 2.16128f
C476 VTAIL.n35 VSUBS 0.014886f
C477 VTAIL.n36 VSUBS 0.015762f
C478 VTAIL.n37 VSUBS 0.035186f
C479 VTAIL.n38 VSUBS 0.035186f
C480 VTAIL.n39 VSUBS 0.015762f
C481 VTAIL.n40 VSUBS 0.014886f
C482 VTAIL.n41 VSUBS 0.027703f
C483 VTAIL.n42 VSUBS 0.027703f
C484 VTAIL.n43 VSUBS 0.014886f
C485 VTAIL.n44 VSUBS 0.015762f
C486 VTAIL.n45 VSUBS 0.035186f
C487 VTAIL.n46 VSUBS 0.035186f
C488 VTAIL.n47 VSUBS 0.015762f
C489 VTAIL.n48 VSUBS 0.014886f
C490 VTAIL.n49 VSUBS 0.027703f
C491 VTAIL.n50 VSUBS 0.027703f
C492 VTAIL.n51 VSUBS 0.014886f
C493 VTAIL.n52 VSUBS 0.015762f
C494 VTAIL.n53 VSUBS 0.035186f
C495 VTAIL.n54 VSUBS 0.035186f
C496 VTAIL.n55 VSUBS 0.015762f
C497 VTAIL.n56 VSUBS 0.014886f
C498 VTAIL.n57 VSUBS 0.027703f
C499 VTAIL.n58 VSUBS 0.027703f
C500 VTAIL.n59 VSUBS 0.014886f
C501 VTAIL.n60 VSUBS 0.015762f
C502 VTAIL.n61 VSUBS 0.035186f
C503 VTAIL.n62 VSUBS 0.035186f
C504 VTAIL.n63 VSUBS 0.015762f
C505 VTAIL.n64 VSUBS 0.014886f
C506 VTAIL.n65 VSUBS 0.027703f
C507 VTAIL.n66 VSUBS 0.027703f
C508 VTAIL.n67 VSUBS 0.014886f
C509 VTAIL.n68 VSUBS 0.015762f
C510 VTAIL.n69 VSUBS 0.035186f
C511 VTAIL.n70 VSUBS 0.035186f
C512 VTAIL.n71 VSUBS 0.015762f
C513 VTAIL.n72 VSUBS 0.014886f
C514 VTAIL.n73 VSUBS 0.027703f
C515 VTAIL.n74 VSUBS 0.027703f
C516 VTAIL.n75 VSUBS 0.014886f
C517 VTAIL.n76 VSUBS 0.014886f
C518 VTAIL.n77 VSUBS 0.015762f
C519 VTAIL.n78 VSUBS 0.035186f
C520 VTAIL.n79 VSUBS 0.035186f
C521 VTAIL.n80 VSUBS 0.035186f
C522 VTAIL.n81 VSUBS 0.015324f
C523 VTAIL.n82 VSUBS 0.014886f
C524 VTAIL.n83 VSUBS 0.027703f
C525 VTAIL.n84 VSUBS 0.027703f
C526 VTAIL.n85 VSUBS 0.014886f
C527 VTAIL.n86 VSUBS 0.015762f
C528 VTAIL.n87 VSUBS 0.035186f
C529 VTAIL.n88 VSUBS 0.035186f
C530 VTAIL.n89 VSUBS 0.015762f
C531 VTAIL.n90 VSUBS 0.014886f
C532 VTAIL.n91 VSUBS 0.027703f
C533 VTAIL.n92 VSUBS 0.027703f
C534 VTAIL.n93 VSUBS 0.014886f
C535 VTAIL.n94 VSUBS 0.015762f
C536 VTAIL.n95 VSUBS 0.035186f
C537 VTAIL.n96 VSUBS 0.079987f
C538 VTAIL.n97 VSUBS 0.015762f
C539 VTAIL.n98 VSUBS 0.014886f
C540 VTAIL.n99 VSUBS 0.059493f
C541 VTAIL.n100 VSUBS 0.03985f
C542 VTAIL.n101 VSUBS 2.20254f
C543 VTAIL.n102 VSUBS 0.028915f
C544 VTAIL.n103 VSUBS 0.027703f
C545 VTAIL.n104 VSUBS 0.014886f
C546 VTAIL.n105 VSUBS 0.035186f
C547 VTAIL.n106 VSUBS 0.015762f
C548 VTAIL.n107 VSUBS 0.027703f
C549 VTAIL.n108 VSUBS 0.014886f
C550 VTAIL.n109 VSUBS 0.035186f
C551 VTAIL.n110 VSUBS 0.015762f
C552 VTAIL.n111 VSUBS 0.027703f
C553 VTAIL.n112 VSUBS 0.015324f
C554 VTAIL.n113 VSUBS 0.035186f
C555 VTAIL.n114 VSUBS 0.014886f
C556 VTAIL.n115 VSUBS 0.015762f
C557 VTAIL.n116 VSUBS 0.027703f
C558 VTAIL.n117 VSUBS 0.014886f
C559 VTAIL.n118 VSUBS 0.035186f
C560 VTAIL.n119 VSUBS 0.015762f
C561 VTAIL.n120 VSUBS 0.027703f
C562 VTAIL.n121 VSUBS 0.014886f
C563 VTAIL.n122 VSUBS 0.035186f
C564 VTAIL.n123 VSUBS 0.015762f
C565 VTAIL.n124 VSUBS 0.027703f
C566 VTAIL.n125 VSUBS 0.014886f
C567 VTAIL.n126 VSUBS 0.035186f
C568 VTAIL.n127 VSUBS 0.015762f
C569 VTAIL.n128 VSUBS 0.027703f
C570 VTAIL.n129 VSUBS 0.014886f
C571 VTAIL.n130 VSUBS 0.035186f
C572 VTAIL.n131 VSUBS 0.015762f
C573 VTAIL.n132 VSUBS 0.027703f
C574 VTAIL.n133 VSUBS 0.014886f
C575 VTAIL.n134 VSUBS 0.02639f
C576 VTAIL.n135 VSUBS 0.022384f
C577 VTAIL.t2 VSUBS 0.075541f
C578 VTAIL.n136 VSUBS 0.220777f
C579 VTAIL.n137 VSUBS 2.16128f
C580 VTAIL.n138 VSUBS 0.014886f
C581 VTAIL.n139 VSUBS 0.015762f
C582 VTAIL.n140 VSUBS 0.035186f
C583 VTAIL.n141 VSUBS 0.035186f
C584 VTAIL.n142 VSUBS 0.015762f
C585 VTAIL.n143 VSUBS 0.014886f
C586 VTAIL.n144 VSUBS 0.027703f
C587 VTAIL.n145 VSUBS 0.027703f
C588 VTAIL.n146 VSUBS 0.014886f
C589 VTAIL.n147 VSUBS 0.015762f
C590 VTAIL.n148 VSUBS 0.035186f
C591 VTAIL.n149 VSUBS 0.035186f
C592 VTAIL.n150 VSUBS 0.015762f
C593 VTAIL.n151 VSUBS 0.014886f
C594 VTAIL.n152 VSUBS 0.027703f
C595 VTAIL.n153 VSUBS 0.027703f
C596 VTAIL.n154 VSUBS 0.014886f
C597 VTAIL.n155 VSUBS 0.015762f
C598 VTAIL.n156 VSUBS 0.035186f
C599 VTAIL.n157 VSUBS 0.035186f
C600 VTAIL.n158 VSUBS 0.015762f
C601 VTAIL.n159 VSUBS 0.014886f
C602 VTAIL.n160 VSUBS 0.027703f
C603 VTAIL.n161 VSUBS 0.027703f
C604 VTAIL.n162 VSUBS 0.014886f
C605 VTAIL.n163 VSUBS 0.015762f
C606 VTAIL.n164 VSUBS 0.035186f
C607 VTAIL.n165 VSUBS 0.035186f
C608 VTAIL.n166 VSUBS 0.015762f
C609 VTAIL.n167 VSUBS 0.014886f
C610 VTAIL.n168 VSUBS 0.027703f
C611 VTAIL.n169 VSUBS 0.027703f
C612 VTAIL.n170 VSUBS 0.014886f
C613 VTAIL.n171 VSUBS 0.015762f
C614 VTAIL.n172 VSUBS 0.035186f
C615 VTAIL.n173 VSUBS 0.035186f
C616 VTAIL.n174 VSUBS 0.015762f
C617 VTAIL.n175 VSUBS 0.014886f
C618 VTAIL.n176 VSUBS 0.027703f
C619 VTAIL.n177 VSUBS 0.027703f
C620 VTAIL.n178 VSUBS 0.014886f
C621 VTAIL.n179 VSUBS 0.015762f
C622 VTAIL.n180 VSUBS 0.035186f
C623 VTAIL.n181 VSUBS 0.035186f
C624 VTAIL.n182 VSUBS 0.035186f
C625 VTAIL.n183 VSUBS 0.015324f
C626 VTAIL.n184 VSUBS 0.014886f
C627 VTAIL.n185 VSUBS 0.027703f
C628 VTAIL.n186 VSUBS 0.027703f
C629 VTAIL.n187 VSUBS 0.014886f
C630 VTAIL.n188 VSUBS 0.015762f
C631 VTAIL.n189 VSUBS 0.035186f
C632 VTAIL.n190 VSUBS 0.035186f
C633 VTAIL.n191 VSUBS 0.015762f
C634 VTAIL.n192 VSUBS 0.014886f
C635 VTAIL.n193 VSUBS 0.027703f
C636 VTAIL.n194 VSUBS 0.027703f
C637 VTAIL.n195 VSUBS 0.014886f
C638 VTAIL.n196 VSUBS 0.015762f
C639 VTAIL.n197 VSUBS 0.035186f
C640 VTAIL.n198 VSUBS 0.079987f
C641 VTAIL.n199 VSUBS 0.015762f
C642 VTAIL.n200 VSUBS 0.014886f
C643 VTAIL.n201 VSUBS 0.059493f
C644 VTAIL.n202 VSUBS 0.03985f
C645 VTAIL.n203 VSUBS 2.23775f
C646 VTAIL.n204 VSUBS 0.028915f
C647 VTAIL.n205 VSUBS 0.027703f
C648 VTAIL.n206 VSUBS 0.014886f
C649 VTAIL.n207 VSUBS 0.035186f
C650 VTAIL.n208 VSUBS 0.015762f
C651 VTAIL.n209 VSUBS 0.027703f
C652 VTAIL.n210 VSUBS 0.014886f
C653 VTAIL.n211 VSUBS 0.035186f
C654 VTAIL.n212 VSUBS 0.015762f
C655 VTAIL.n213 VSUBS 0.027703f
C656 VTAIL.n214 VSUBS 0.015324f
C657 VTAIL.n215 VSUBS 0.035186f
C658 VTAIL.n216 VSUBS 0.014886f
C659 VTAIL.n217 VSUBS 0.015762f
C660 VTAIL.n218 VSUBS 0.027703f
C661 VTAIL.n219 VSUBS 0.014886f
C662 VTAIL.n220 VSUBS 0.035186f
C663 VTAIL.n221 VSUBS 0.015762f
C664 VTAIL.n222 VSUBS 0.027703f
C665 VTAIL.n223 VSUBS 0.014886f
C666 VTAIL.n224 VSUBS 0.035186f
C667 VTAIL.n225 VSUBS 0.015762f
C668 VTAIL.n226 VSUBS 0.027703f
C669 VTAIL.n227 VSUBS 0.014886f
C670 VTAIL.n228 VSUBS 0.035186f
C671 VTAIL.n229 VSUBS 0.015762f
C672 VTAIL.n230 VSUBS 0.027703f
C673 VTAIL.n231 VSUBS 0.014886f
C674 VTAIL.n232 VSUBS 0.035186f
C675 VTAIL.n233 VSUBS 0.015762f
C676 VTAIL.n234 VSUBS 0.027703f
C677 VTAIL.n235 VSUBS 0.014886f
C678 VTAIL.n236 VSUBS 0.02639f
C679 VTAIL.n237 VSUBS 0.022384f
C680 VTAIL.t1 VSUBS 0.075541f
C681 VTAIL.n238 VSUBS 0.220777f
C682 VTAIL.n239 VSUBS 2.16128f
C683 VTAIL.n240 VSUBS 0.014886f
C684 VTAIL.n241 VSUBS 0.015762f
C685 VTAIL.n242 VSUBS 0.035186f
C686 VTAIL.n243 VSUBS 0.035186f
C687 VTAIL.n244 VSUBS 0.015762f
C688 VTAIL.n245 VSUBS 0.014886f
C689 VTAIL.n246 VSUBS 0.027703f
C690 VTAIL.n247 VSUBS 0.027703f
C691 VTAIL.n248 VSUBS 0.014886f
C692 VTAIL.n249 VSUBS 0.015762f
C693 VTAIL.n250 VSUBS 0.035186f
C694 VTAIL.n251 VSUBS 0.035186f
C695 VTAIL.n252 VSUBS 0.015762f
C696 VTAIL.n253 VSUBS 0.014886f
C697 VTAIL.n254 VSUBS 0.027703f
C698 VTAIL.n255 VSUBS 0.027703f
C699 VTAIL.n256 VSUBS 0.014886f
C700 VTAIL.n257 VSUBS 0.015762f
C701 VTAIL.n258 VSUBS 0.035186f
C702 VTAIL.n259 VSUBS 0.035186f
C703 VTAIL.n260 VSUBS 0.015762f
C704 VTAIL.n261 VSUBS 0.014886f
C705 VTAIL.n262 VSUBS 0.027703f
C706 VTAIL.n263 VSUBS 0.027703f
C707 VTAIL.n264 VSUBS 0.014886f
C708 VTAIL.n265 VSUBS 0.015762f
C709 VTAIL.n266 VSUBS 0.035186f
C710 VTAIL.n267 VSUBS 0.035186f
C711 VTAIL.n268 VSUBS 0.015762f
C712 VTAIL.n269 VSUBS 0.014886f
C713 VTAIL.n270 VSUBS 0.027703f
C714 VTAIL.n271 VSUBS 0.027703f
C715 VTAIL.n272 VSUBS 0.014886f
C716 VTAIL.n273 VSUBS 0.015762f
C717 VTAIL.n274 VSUBS 0.035186f
C718 VTAIL.n275 VSUBS 0.035186f
C719 VTAIL.n276 VSUBS 0.015762f
C720 VTAIL.n277 VSUBS 0.014886f
C721 VTAIL.n278 VSUBS 0.027703f
C722 VTAIL.n279 VSUBS 0.027703f
C723 VTAIL.n280 VSUBS 0.014886f
C724 VTAIL.n281 VSUBS 0.015762f
C725 VTAIL.n282 VSUBS 0.035186f
C726 VTAIL.n283 VSUBS 0.035186f
C727 VTAIL.n284 VSUBS 0.035186f
C728 VTAIL.n285 VSUBS 0.015324f
C729 VTAIL.n286 VSUBS 0.014886f
C730 VTAIL.n287 VSUBS 0.027703f
C731 VTAIL.n288 VSUBS 0.027703f
C732 VTAIL.n289 VSUBS 0.014886f
C733 VTAIL.n290 VSUBS 0.015762f
C734 VTAIL.n291 VSUBS 0.035186f
C735 VTAIL.n292 VSUBS 0.035186f
C736 VTAIL.n293 VSUBS 0.015762f
C737 VTAIL.n294 VSUBS 0.014886f
C738 VTAIL.n295 VSUBS 0.027703f
C739 VTAIL.n296 VSUBS 0.027703f
C740 VTAIL.n297 VSUBS 0.014886f
C741 VTAIL.n298 VSUBS 0.015762f
C742 VTAIL.n299 VSUBS 0.035186f
C743 VTAIL.n300 VSUBS 0.079987f
C744 VTAIL.n301 VSUBS 0.015762f
C745 VTAIL.n302 VSUBS 0.014886f
C746 VTAIL.n303 VSUBS 0.059493f
C747 VTAIL.n304 VSUBS 0.03985f
C748 VTAIL.n305 VSUBS 2.07615f
C749 VTAIL.n306 VSUBS 0.028915f
C750 VTAIL.n307 VSUBS 0.027703f
C751 VTAIL.n308 VSUBS 0.014886f
C752 VTAIL.n309 VSUBS 0.035186f
C753 VTAIL.n310 VSUBS 0.015762f
C754 VTAIL.n311 VSUBS 0.027703f
C755 VTAIL.n312 VSUBS 0.014886f
C756 VTAIL.n313 VSUBS 0.035186f
C757 VTAIL.n314 VSUBS 0.015762f
C758 VTAIL.n315 VSUBS 0.027703f
C759 VTAIL.n316 VSUBS 0.015324f
C760 VTAIL.n317 VSUBS 0.035186f
C761 VTAIL.n318 VSUBS 0.015762f
C762 VTAIL.n319 VSUBS 0.027703f
C763 VTAIL.n320 VSUBS 0.014886f
C764 VTAIL.n321 VSUBS 0.035186f
C765 VTAIL.n322 VSUBS 0.015762f
C766 VTAIL.n323 VSUBS 0.027703f
C767 VTAIL.n324 VSUBS 0.014886f
C768 VTAIL.n325 VSUBS 0.035186f
C769 VTAIL.n326 VSUBS 0.015762f
C770 VTAIL.n327 VSUBS 0.027703f
C771 VTAIL.n328 VSUBS 0.014886f
C772 VTAIL.n329 VSUBS 0.035186f
C773 VTAIL.n330 VSUBS 0.015762f
C774 VTAIL.n331 VSUBS 0.027703f
C775 VTAIL.n332 VSUBS 0.014886f
C776 VTAIL.n333 VSUBS 0.035186f
C777 VTAIL.n334 VSUBS 0.015762f
C778 VTAIL.n335 VSUBS 0.027703f
C779 VTAIL.n336 VSUBS 0.014886f
C780 VTAIL.n337 VSUBS 0.02639f
C781 VTAIL.n338 VSUBS 0.022384f
C782 VTAIL.t3 VSUBS 0.075541f
C783 VTAIL.n339 VSUBS 0.220777f
C784 VTAIL.n340 VSUBS 2.16128f
C785 VTAIL.n341 VSUBS 0.014886f
C786 VTAIL.n342 VSUBS 0.015762f
C787 VTAIL.n343 VSUBS 0.035186f
C788 VTAIL.n344 VSUBS 0.035186f
C789 VTAIL.n345 VSUBS 0.015762f
C790 VTAIL.n346 VSUBS 0.014886f
C791 VTAIL.n347 VSUBS 0.027703f
C792 VTAIL.n348 VSUBS 0.027703f
C793 VTAIL.n349 VSUBS 0.014886f
C794 VTAIL.n350 VSUBS 0.015762f
C795 VTAIL.n351 VSUBS 0.035186f
C796 VTAIL.n352 VSUBS 0.035186f
C797 VTAIL.n353 VSUBS 0.015762f
C798 VTAIL.n354 VSUBS 0.014886f
C799 VTAIL.n355 VSUBS 0.027703f
C800 VTAIL.n356 VSUBS 0.027703f
C801 VTAIL.n357 VSUBS 0.014886f
C802 VTAIL.n358 VSUBS 0.015762f
C803 VTAIL.n359 VSUBS 0.035186f
C804 VTAIL.n360 VSUBS 0.035186f
C805 VTAIL.n361 VSUBS 0.015762f
C806 VTAIL.n362 VSUBS 0.014886f
C807 VTAIL.n363 VSUBS 0.027703f
C808 VTAIL.n364 VSUBS 0.027703f
C809 VTAIL.n365 VSUBS 0.014886f
C810 VTAIL.n366 VSUBS 0.015762f
C811 VTAIL.n367 VSUBS 0.035186f
C812 VTAIL.n368 VSUBS 0.035186f
C813 VTAIL.n369 VSUBS 0.015762f
C814 VTAIL.n370 VSUBS 0.014886f
C815 VTAIL.n371 VSUBS 0.027703f
C816 VTAIL.n372 VSUBS 0.027703f
C817 VTAIL.n373 VSUBS 0.014886f
C818 VTAIL.n374 VSUBS 0.015762f
C819 VTAIL.n375 VSUBS 0.035186f
C820 VTAIL.n376 VSUBS 0.035186f
C821 VTAIL.n377 VSUBS 0.015762f
C822 VTAIL.n378 VSUBS 0.014886f
C823 VTAIL.n379 VSUBS 0.027703f
C824 VTAIL.n380 VSUBS 0.027703f
C825 VTAIL.n381 VSUBS 0.014886f
C826 VTAIL.n382 VSUBS 0.014886f
C827 VTAIL.n383 VSUBS 0.015762f
C828 VTAIL.n384 VSUBS 0.035186f
C829 VTAIL.n385 VSUBS 0.035186f
C830 VTAIL.n386 VSUBS 0.035186f
C831 VTAIL.n387 VSUBS 0.015324f
C832 VTAIL.n388 VSUBS 0.014886f
C833 VTAIL.n389 VSUBS 0.027703f
C834 VTAIL.n390 VSUBS 0.027703f
C835 VTAIL.n391 VSUBS 0.014886f
C836 VTAIL.n392 VSUBS 0.015762f
C837 VTAIL.n393 VSUBS 0.035186f
C838 VTAIL.n394 VSUBS 0.035186f
C839 VTAIL.n395 VSUBS 0.015762f
C840 VTAIL.n396 VSUBS 0.014886f
C841 VTAIL.n397 VSUBS 0.027703f
C842 VTAIL.n398 VSUBS 0.027703f
C843 VTAIL.n399 VSUBS 0.014886f
C844 VTAIL.n400 VSUBS 0.015762f
C845 VTAIL.n401 VSUBS 0.035186f
C846 VTAIL.n402 VSUBS 0.079987f
C847 VTAIL.n403 VSUBS 0.015762f
C848 VTAIL.n404 VSUBS 0.014886f
C849 VTAIL.n405 VSUBS 0.059493f
C850 VTAIL.n406 VSUBS 0.03985f
C851 VTAIL.n407 VSUBS 1.98861f
C852 VN.t1 VSUBS 4.19422f
C853 VN.t0 VSUBS 4.67264f
C854 B.n0 VSUBS 0.006712f
C855 B.n1 VSUBS 0.006712f
C856 B.n2 VSUBS 0.009926f
C857 B.n3 VSUBS 0.007607f
C858 B.n4 VSUBS 0.007607f
C859 B.n5 VSUBS 0.007607f
C860 B.n6 VSUBS 0.007607f
C861 B.n7 VSUBS 0.007607f
C862 B.n8 VSUBS 0.007607f
C863 B.n9 VSUBS 0.007607f
C864 B.n10 VSUBS 0.007607f
C865 B.n11 VSUBS 0.007607f
C866 B.n12 VSUBS 0.017723f
C867 B.n13 VSUBS 0.007607f
C868 B.n14 VSUBS 0.007607f
C869 B.n15 VSUBS 0.007607f
C870 B.n16 VSUBS 0.007607f
C871 B.n17 VSUBS 0.007607f
C872 B.n18 VSUBS 0.007607f
C873 B.n19 VSUBS 0.007607f
C874 B.n20 VSUBS 0.007607f
C875 B.n21 VSUBS 0.007607f
C876 B.n22 VSUBS 0.007607f
C877 B.n23 VSUBS 0.007607f
C878 B.n24 VSUBS 0.007607f
C879 B.n25 VSUBS 0.007607f
C880 B.n26 VSUBS 0.007607f
C881 B.n27 VSUBS 0.007607f
C882 B.n28 VSUBS 0.007607f
C883 B.n29 VSUBS 0.007607f
C884 B.n30 VSUBS 0.007607f
C885 B.n31 VSUBS 0.007607f
C886 B.n32 VSUBS 0.007607f
C887 B.n33 VSUBS 0.007607f
C888 B.n34 VSUBS 0.007607f
C889 B.n35 VSUBS 0.007607f
C890 B.n36 VSUBS 0.007607f
C891 B.n37 VSUBS 0.007607f
C892 B.n38 VSUBS 0.007607f
C893 B.n39 VSUBS 0.007607f
C894 B.n40 VSUBS 0.007607f
C895 B.n41 VSUBS 0.007607f
C896 B.t10 VSUBS 0.384549f
C897 B.t11 VSUBS 0.411182f
C898 B.t9 VSUBS 1.50052f
C899 B.n42 VSUBS 0.592129f
C900 B.n43 VSUBS 0.355146f
C901 B.n44 VSUBS 0.017624f
C902 B.n45 VSUBS 0.007607f
C903 B.n46 VSUBS 0.007607f
C904 B.n47 VSUBS 0.007607f
C905 B.n48 VSUBS 0.007607f
C906 B.n49 VSUBS 0.007607f
C907 B.t1 VSUBS 0.384552f
C908 B.t2 VSUBS 0.411186f
C909 B.t0 VSUBS 1.50052f
C910 B.n50 VSUBS 0.592125f
C911 B.n51 VSUBS 0.355143f
C912 B.n52 VSUBS 0.007607f
C913 B.n53 VSUBS 0.007607f
C914 B.n54 VSUBS 0.007607f
C915 B.n55 VSUBS 0.007607f
C916 B.n56 VSUBS 0.007607f
C917 B.n57 VSUBS 0.007607f
C918 B.n58 VSUBS 0.007607f
C919 B.n59 VSUBS 0.007607f
C920 B.n60 VSUBS 0.007607f
C921 B.n61 VSUBS 0.007607f
C922 B.n62 VSUBS 0.007607f
C923 B.n63 VSUBS 0.007607f
C924 B.n64 VSUBS 0.007607f
C925 B.n65 VSUBS 0.007607f
C926 B.n66 VSUBS 0.007607f
C927 B.n67 VSUBS 0.007607f
C928 B.n68 VSUBS 0.007607f
C929 B.n69 VSUBS 0.007607f
C930 B.n70 VSUBS 0.007607f
C931 B.n71 VSUBS 0.007607f
C932 B.n72 VSUBS 0.007607f
C933 B.n73 VSUBS 0.007607f
C934 B.n74 VSUBS 0.007607f
C935 B.n75 VSUBS 0.007607f
C936 B.n76 VSUBS 0.007607f
C937 B.n77 VSUBS 0.007607f
C938 B.n78 VSUBS 0.007607f
C939 B.n79 VSUBS 0.007607f
C940 B.n80 VSUBS 0.007607f
C941 B.n81 VSUBS 0.016732f
C942 B.n82 VSUBS 0.007607f
C943 B.n83 VSUBS 0.007607f
C944 B.n84 VSUBS 0.007607f
C945 B.n85 VSUBS 0.007607f
C946 B.n86 VSUBS 0.007607f
C947 B.n87 VSUBS 0.007607f
C948 B.n88 VSUBS 0.007607f
C949 B.n89 VSUBS 0.007607f
C950 B.n90 VSUBS 0.007607f
C951 B.n91 VSUBS 0.007607f
C952 B.n92 VSUBS 0.007607f
C953 B.n93 VSUBS 0.007607f
C954 B.n94 VSUBS 0.007607f
C955 B.n95 VSUBS 0.007607f
C956 B.n96 VSUBS 0.007607f
C957 B.n97 VSUBS 0.007607f
C958 B.n98 VSUBS 0.007607f
C959 B.n99 VSUBS 0.007607f
C960 B.n100 VSUBS 0.007607f
C961 B.n101 VSUBS 0.007607f
C962 B.n102 VSUBS 0.016778f
C963 B.n103 VSUBS 0.007607f
C964 B.n104 VSUBS 0.007607f
C965 B.n105 VSUBS 0.007607f
C966 B.n106 VSUBS 0.007607f
C967 B.n107 VSUBS 0.007607f
C968 B.n108 VSUBS 0.007607f
C969 B.n109 VSUBS 0.007607f
C970 B.n110 VSUBS 0.007607f
C971 B.n111 VSUBS 0.007607f
C972 B.n112 VSUBS 0.007607f
C973 B.n113 VSUBS 0.007607f
C974 B.n114 VSUBS 0.007607f
C975 B.n115 VSUBS 0.007607f
C976 B.n116 VSUBS 0.007607f
C977 B.n117 VSUBS 0.007607f
C978 B.n118 VSUBS 0.007607f
C979 B.n119 VSUBS 0.007607f
C980 B.n120 VSUBS 0.007607f
C981 B.n121 VSUBS 0.007607f
C982 B.n122 VSUBS 0.007607f
C983 B.n123 VSUBS 0.007607f
C984 B.n124 VSUBS 0.007607f
C985 B.n125 VSUBS 0.007607f
C986 B.n126 VSUBS 0.007607f
C987 B.n127 VSUBS 0.007607f
C988 B.n128 VSUBS 0.007607f
C989 B.n129 VSUBS 0.007607f
C990 B.n130 VSUBS 0.007607f
C991 B.n131 VSUBS 0.007607f
C992 B.t5 VSUBS 0.384552f
C993 B.t4 VSUBS 0.411186f
C994 B.t3 VSUBS 1.50052f
C995 B.n132 VSUBS 0.592125f
C996 B.n133 VSUBS 0.355143f
C997 B.n134 VSUBS 0.017624f
C998 B.n135 VSUBS 0.007607f
C999 B.n136 VSUBS 0.007607f
C1000 B.n137 VSUBS 0.007607f
C1001 B.n138 VSUBS 0.007607f
C1002 B.n139 VSUBS 0.007607f
C1003 B.t8 VSUBS 0.384549f
C1004 B.t7 VSUBS 0.411182f
C1005 B.t6 VSUBS 1.50052f
C1006 B.n140 VSUBS 0.592129f
C1007 B.n141 VSUBS 0.355146f
C1008 B.n142 VSUBS 0.007607f
C1009 B.n143 VSUBS 0.007607f
C1010 B.n144 VSUBS 0.007607f
C1011 B.n145 VSUBS 0.007607f
C1012 B.n146 VSUBS 0.007607f
C1013 B.n147 VSUBS 0.007607f
C1014 B.n148 VSUBS 0.007607f
C1015 B.n149 VSUBS 0.007607f
C1016 B.n150 VSUBS 0.007607f
C1017 B.n151 VSUBS 0.007607f
C1018 B.n152 VSUBS 0.007607f
C1019 B.n153 VSUBS 0.007607f
C1020 B.n154 VSUBS 0.007607f
C1021 B.n155 VSUBS 0.007607f
C1022 B.n156 VSUBS 0.007607f
C1023 B.n157 VSUBS 0.007607f
C1024 B.n158 VSUBS 0.007607f
C1025 B.n159 VSUBS 0.007607f
C1026 B.n160 VSUBS 0.007607f
C1027 B.n161 VSUBS 0.007607f
C1028 B.n162 VSUBS 0.007607f
C1029 B.n163 VSUBS 0.007607f
C1030 B.n164 VSUBS 0.007607f
C1031 B.n165 VSUBS 0.007607f
C1032 B.n166 VSUBS 0.007607f
C1033 B.n167 VSUBS 0.007607f
C1034 B.n168 VSUBS 0.007607f
C1035 B.n169 VSUBS 0.007607f
C1036 B.n170 VSUBS 0.007607f
C1037 B.n171 VSUBS 0.016732f
C1038 B.n172 VSUBS 0.007607f
C1039 B.n173 VSUBS 0.007607f
C1040 B.n174 VSUBS 0.007607f
C1041 B.n175 VSUBS 0.007607f
C1042 B.n176 VSUBS 0.007607f
C1043 B.n177 VSUBS 0.007607f
C1044 B.n178 VSUBS 0.007607f
C1045 B.n179 VSUBS 0.007607f
C1046 B.n180 VSUBS 0.007607f
C1047 B.n181 VSUBS 0.007607f
C1048 B.n182 VSUBS 0.007607f
C1049 B.n183 VSUBS 0.007607f
C1050 B.n184 VSUBS 0.007607f
C1051 B.n185 VSUBS 0.007607f
C1052 B.n186 VSUBS 0.007607f
C1053 B.n187 VSUBS 0.007607f
C1054 B.n188 VSUBS 0.007607f
C1055 B.n189 VSUBS 0.007607f
C1056 B.n190 VSUBS 0.007607f
C1057 B.n191 VSUBS 0.007607f
C1058 B.n192 VSUBS 0.007607f
C1059 B.n193 VSUBS 0.007607f
C1060 B.n194 VSUBS 0.007607f
C1061 B.n195 VSUBS 0.007607f
C1062 B.n196 VSUBS 0.007607f
C1063 B.n197 VSUBS 0.007607f
C1064 B.n198 VSUBS 0.007607f
C1065 B.n199 VSUBS 0.007607f
C1066 B.n200 VSUBS 0.007607f
C1067 B.n201 VSUBS 0.007607f
C1068 B.n202 VSUBS 0.007607f
C1069 B.n203 VSUBS 0.007607f
C1070 B.n204 VSUBS 0.007607f
C1071 B.n205 VSUBS 0.007607f
C1072 B.n206 VSUBS 0.007607f
C1073 B.n207 VSUBS 0.007607f
C1074 B.n208 VSUBS 0.016732f
C1075 B.n209 VSUBS 0.017723f
C1076 B.n210 VSUBS 0.017723f
C1077 B.n211 VSUBS 0.007607f
C1078 B.n212 VSUBS 0.007607f
C1079 B.n213 VSUBS 0.007607f
C1080 B.n214 VSUBS 0.007607f
C1081 B.n215 VSUBS 0.007607f
C1082 B.n216 VSUBS 0.007607f
C1083 B.n217 VSUBS 0.007607f
C1084 B.n218 VSUBS 0.007607f
C1085 B.n219 VSUBS 0.007607f
C1086 B.n220 VSUBS 0.007607f
C1087 B.n221 VSUBS 0.007607f
C1088 B.n222 VSUBS 0.007607f
C1089 B.n223 VSUBS 0.007607f
C1090 B.n224 VSUBS 0.007607f
C1091 B.n225 VSUBS 0.007607f
C1092 B.n226 VSUBS 0.007607f
C1093 B.n227 VSUBS 0.007607f
C1094 B.n228 VSUBS 0.007607f
C1095 B.n229 VSUBS 0.007607f
C1096 B.n230 VSUBS 0.007607f
C1097 B.n231 VSUBS 0.007607f
C1098 B.n232 VSUBS 0.007607f
C1099 B.n233 VSUBS 0.007607f
C1100 B.n234 VSUBS 0.007607f
C1101 B.n235 VSUBS 0.007607f
C1102 B.n236 VSUBS 0.007607f
C1103 B.n237 VSUBS 0.007607f
C1104 B.n238 VSUBS 0.007607f
C1105 B.n239 VSUBS 0.007607f
C1106 B.n240 VSUBS 0.007607f
C1107 B.n241 VSUBS 0.007607f
C1108 B.n242 VSUBS 0.007607f
C1109 B.n243 VSUBS 0.007607f
C1110 B.n244 VSUBS 0.007607f
C1111 B.n245 VSUBS 0.007607f
C1112 B.n246 VSUBS 0.007607f
C1113 B.n247 VSUBS 0.007607f
C1114 B.n248 VSUBS 0.007607f
C1115 B.n249 VSUBS 0.007607f
C1116 B.n250 VSUBS 0.007607f
C1117 B.n251 VSUBS 0.007607f
C1118 B.n252 VSUBS 0.007607f
C1119 B.n253 VSUBS 0.007607f
C1120 B.n254 VSUBS 0.007607f
C1121 B.n255 VSUBS 0.007607f
C1122 B.n256 VSUBS 0.007607f
C1123 B.n257 VSUBS 0.007607f
C1124 B.n258 VSUBS 0.007607f
C1125 B.n259 VSUBS 0.007607f
C1126 B.n260 VSUBS 0.007607f
C1127 B.n261 VSUBS 0.007607f
C1128 B.n262 VSUBS 0.007607f
C1129 B.n263 VSUBS 0.007607f
C1130 B.n264 VSUBS 0.007607f
C1131 B.n265 VSUBS 0.007607f
C1132 B.n266 VSUBS 0.007607f
C1133 B.n267 VSUBS 0.007607f
C1134 B.n268 VSUBS 0.007607f
C1135 B.n269 VSUBS 0.007607f
C1136 B.n270 VSUBS 0.007607f
C1137 B.n271 VSUBS 0.007607f
C1138 B.n272 VSUBS 0.007607f
C1139 B.n273 VSUBS 0.007607f
C1140 B.n274 VSUBS 0.007607f
C1141 B.n275 VSUBS 0.007607f
C1142 B.n276 VSUBS 0.007607f
C1143 B.n277 VSUBS 0.007607f
C1144 B.n278 VSUBS 0.007607f
C1145 B.n279 VSUBS 0.007607f
C1146 B.n280 VSUBS 0.007607f
C1147 B.n281 VSUBS 0.007607f
C1148 B.n282 VSUBS 0.007607f
C1149 B.n283 VSUBS 0.007607f
C1150 B.n284 VSUBS 0.007607f
C1151 B.n285 VSUBS 0.007607f
C1152 B.n286 VSUBS 0.007607f
C1153 B.n287 VSUBS 0.007607f
C1154 B.n288 VSUBS 0.007607f
C1155 B.n289 VSUBS 0.007607f
C1156 B.n290 VSUBS 0.007607f
C1157 B.n291 VSUBS 0.007607f
C1158 B.n292 VSUBS 0.007607f
C1159 B.n293 VSUBS 0.007607f
C1160 B.n294 VSUBS 0.007607f
C1161 B.n295 VSUBS 0.007607f
C1162 B.n296 VSUBS 0.007607f
C1163 B.n297 VSUBS 0.007607f
C1164 B.n298 VSUBS 0.005258f
C1165 B.n299 VSUBS 0.017624f
C1166 B.n300 VSUBS 0.006153f
C1167 B.n301 VSUBS 0.007607f
C1168 B.n302 VSUBS 0.007607f
C1169 B.n303 VSUBS 0.007607f
C1170 B.n304 VSUBS 0.007607f
C1171 B.n305 VSUBS 0.007607f
C1172 B.n306 VSUBS 0.007607f
C1173 B.n307 VSUBS 0.007607f
C1174 B.n308 VSUBS 0.007607f
C1175 B.n309 VSUBS 0.007607f
C1176 B.n310 VSUBS 0.007607f
C1177 B.n311 VSUBS 0.007607f
C1178 B.n312 VSUBS 0.006153f
C1179 B.n313 VSUBS 0.007607f
C1180 B.n314 VSUBS 0.007607f
C1181 B.n315 VSUBS 0.005258f
C1182 B.n316 VSUBS 0.007607f
C1183 B.n317 VSUBS 0.007607f
C1184 B.n318 VSUBS 0.007607f
C1185 B.n319 VSUBS 0.007607f
C1186 B.n320 VSUBS 0.007607f
C1187 B.n321 VSUBS 0.007607f
C1188 B.n322 VSUBS 0.007607f
C1189 B.n323 VSUBS 0.007607f
C1190 B.n324 VSUBS 0.007607f
C1191 B.n325 VSUBS 0.007607f
C1192 B.n326 VSUBS 0.007607f
C1193 B.n327 VSUBS 0.007607f
C1194 B.n328 VSUBS 0.007607f
C1195 B.n329 VSUBS 0.007607f
C1196 B.n330 VSUBS 0.007607f
C1197 B.n331 VSUBS 0.007607f
C1198 B.n332 VSUBS 0.007607f
C1199 B.n333 VSUBS 0.007607f
C1200 B.n334 VSUBS 0.007607f
C1201 B.n335 VSUBS 0.007607f
C1202 B.n336 VSUBS 0.007607f
C1203 B.n337 VSUBS 0.007607f
C1204 B.n338 VSUBS 0.007607f
C1205 B.n339 VSUBS 0.007607f
C1206 B.n340 VSUBS 0.007607f
C1207 B.n341 VSUBS 0.007607f
C1208 B.n342 VSUBS 0.007607f
C1209 B.n343 VSUBS 0.007607f
C1210 B.n344 VSUBS 0.007607f
C1211 B.n345 VSUBS 0.007607f
C1212 B.n346 VSUBS 0.007607f
C1213 B.n347 VSUBS 0.007607f
C1214 B.n348 VSUBS 0.007607f
C1215 B.n349 VSUBS 0.007607f
C1216 B.n350 VSUBS 0.007607f
C1217 B.n351 VSUBS 0.007607f
C1218 B.n352 VSUBS 0.007607f
C1219 B.n353 VSUBS 0.007607f
C1220 B.n354 VSUBS 0.007607f
C1221 B.n355 VSUBS 0.007607f
C1222 B.n356 VSUBS 0.007607f
C1223 B.n357 VSUBS 0.007607f
C1224 B.n358 VSUBS 0.007607f
C1225 B.n359 VSUBS 0.007607f
C1226 B.n360 VSUBS 0.007607f
C1227 B.n361 VSUBS 0.007607f
C1228 B.n362 VSUBS 0.007607f
C1229 B.n363 VSUBS 0.007607f
C1230 B.n364 VSUBS 0.007607f
C1231 B.n365 VSUBS 0.007607f
C1232 B.n366 VSUBS 0.007607f
C1233 B.n367 VSUBS 0.007607f
C1234 B.n368 VSUBS 0.007607f
C1235 B.n369 VSUBS 0.007607f
C1236 B.n370 VSUBS 0.007607f
C1237 B.n371 VSUBS 0.007607f
C1238 B.n372 VSUBS 0.007607f
C1239 B.n373 VSUBS 0.007607f
C1240 B.n374 VSUBS 0.007607f
C1241 B.n375 VSUBS 0.007607f
C1242 B.n376 VSUBS 0.007607f
C1243 B.n377 VSUBS 0.007607f
C1244 B.n378 VSUBS 0.007607f
C1245 B.n379 VSUBS 0.007607f
C1246 B.n380 VSUBS 0.007607f
C1247 B.n381 VSUBS 0.007607f
C1248 B.n382 VSUBS 0.007607f
C1249 B.n383 VSUBS 0.007607f
C1250 B.n384 VSUBS 0.007607f
C1251 B.n385 VSUBS 0.007607f
C1252 B.n386 VSUBS 0.007607f
C1253 B.n387 VSUBS 0.007607f
C1254 B.n388 VSUBS 0.007607f
C1255 B.n389 VSUBS 0.007607f
C1256 B.n390 VSUBS 0.007607f
C1257 B.n391 VSUBS 0.007607f
C1258 B.n392 VSUBS 0.007607f
C1259 B.n393 VSUBS 0.007607f
C1260 B.n394 VSUBS 0.007607f
C1261 B.n395 VSUBS 0.007607f
C1262 B.n396 VSUBS 0.007607f
C1263 B.n397 VSUBS 0.007607f
C1264 B.n398 VSUBS 0.007607f
C1265 B.n399 VSUBS 0.007607f
C1266 B.n400 VSUBS 0.007607f
C1267 B.n401 VSUBS 0.007607f
C1268 B.n402 VSUBS 0.007607f
C1269 B.n403 VSUBS 0.017723f
C1270 B.n404 VSUBS 0.016732f
C1271 B.n405 VSUBS 0.017677f
C1272 B.n406 VSUBS 0.007607f
C1273 B.n407 VSUBS 0.007607f
C1274 B.n408 VSUBS 0.007607f
C1275 B.n409 VSUBS 0.007607f
C1276 B.n410 VSUBS 0.007607f
C1277 B.n411 VSUBS 0.007607f
C1278 B.n412 VSUBS 0.007607f
C1279 B.n413 VSUBS 0.007607f
C1280 B.n414 VSUBS 0.007607f
C1281 B.n415 VSUBS 0.007607f
C1282 B.n416 VSUBS 0.007607f
C1283 B.n417 VSUBS 0.007607f
C1284 B.n418 VSUBS 0.007607f
C1285 B.n419 VSUBS 0.007607f
C1286 B.n420 VSUBS 0.007607f
C1287 B.n421 VSUBS 0.007607f
C1288 B.n422 VSUBS 0.007607f
C1289 B.n423 VSUBS 0.007607f
C1290 B.n424 VSUBS 0.007607f
C1291 B.n425 VSUBS 0.007607f
C1292 B.n426 VSUBS 0.007607f
C1293 B.n427 VSUBS 0.007607f
C1294 B.n428 VSUBS 0.007607f
C1295 B.n429 VSUBS 0.007607f
C1296 B.n430 VSUBS 0.007607f
C1297 B.n431 VSUBS 0.007607f
C1298 B.n432 VSUBS 0.007607f
C1299 B.n433 VSUBS 0.007607f
C1300 B.n434 VSUBS 0.007607f
C1301 B.n435 VSUBS 0.007607f
C1302 B.n436 VSUBS 0.007607f
C1303 B.n437 VSUBS 0.007607f
C1304 B.n438 VSUBS 0.007607f
C1305 B.n439 VSUBS 0.007607f
C1306 B.n440 VSUBS 0.007607f
C1307 B.n441 VSUBS 0.007607f
C1308 B.n442 VSUBS 0.007607f
C1309 B.n443 VSUBS 0.007607f
C1310 B.n444 VSUBS 0.007607f
C1311 B.n445 VSUBS 0.007607f
C1312 B.n446 VSUBS 0.007607f
C1313 B.n447 VSUBS 0.007607f
C1314 B.n448 VSUBS 0.007607f
C1315 B.n449 VSUBS 0.007607f
C1316 B.n450 VSUBS 0.007607f
C1317 B.n451 VSUBS 0.007607f
C1318 B.n452 VSUBS 0.007607f
C1319 B.n453 VSUBS 0.007607f
C1320 B.n454 VSUBS 0.007607f
C1321 B.n455 VSUBS 0.007607f
C1322 B.n456 VSUBS 0.007607f
C1323 B.n457 VSUBS 0.007607f
C1324 B.n458 VSUBS 0.007607f
C1325 B.n459 VSUBS 0.007607f
C1326 B.n460 VSUBS 0.007607f
C1327 B.n461 VSUBS 0.007607f
C1328 B.n462 VSUBS 0.007607f
C1329 B.n463 VSUBS 0.007607f
C1330 B.n464 VSUBS 0.007607f
C1331 B.n465 VSUBS 0.007607f
C1332 B.n466 VSUBS 0.016732f
C1333 B.n467 VSUBS 0.017723f
C1334 B.n468 VSUBS 0.017723f
C1335 B.n469 VSUBS 0.007607f
C1336 B.n470 VSUBS 0.007607f
C1337 B.n471 VSUBS 0.007607f
C1338 B.n472 VSUBS 0.007607f
C1339 B.n473 VSUBS 0.007607f
C1340 B.n474 VSUBS 0.007607f
C1341 B.n475 VSUBS 0.007607f
C1342 B.n476 VSUBS 0.007607f
C1343 B.n477 VSUBS 0.007607f
C1344 B.n478 VSUBS 0.007607f
C1345 B.n479 VSUBS 0.007607f
C1346 B.n480 VSUBS 0.007607f
C1347 B.n481 VSUBS 0.007607f
C1348 B.n482 VSUBS 0.007607f
C1349 B.n483 VSUBS 0.007607f
C1350 B.n484 VSUBS 0.007607f
C1351 B.n485 VSUBS 0.007607f
C1352 B.n486 VSUBS 0.007607f
C1353 B.n487 VSUBS 0.007607f
C1354 B.n488 VSUBS 0.007607f
C1355 B.n489 VSUBS 0.007607f
C1356 B.n490 VSUBS 0.007607f
C1357 B.n491 VSUBS 0.007607f
C1358 B.n492 VSUBS 0.007607f
C1359 B.n493 VSUBS 0.007607f
C1360 B.n494 VSUBS 0.007607f
C1361 B.n495 VSUBS 0.007607f
C1362 B.n496 VSUBS 0.007607f
C1363 B.n497 VSUBS 0.007607f
C1364 B.n498 VSUBS 0.007607f
C1365 B.n499 VSUBS 0.007607f
C1366 B.n500 VSUBS 0.007607f
C1367 B.n501 VSUBS 0.007607f
C1368 B.n502 VSUBS 0.007607f
C1369 B.n503 VSUBS 0.007607f
C1370 B.n504 VSUBS 0.007607f
C1371 B.n505 VSUBS 0.007607f
C1372 B.n506 VSUBS 0.007607f
C1373 B.n507 VSUBS 0.007607f
C1374 B.n508 VSUBS 0.007607f
C1375 B.n509 VSUBS 0.007607f
C1376 B.n510 VSUBS 0.007607f
C1377 B.n511 VSUBS 0.007607f
C1378 B.n512 VSUBS 0.007607f
C1379 B.n513 VSUBS 0.007607f
C1380 B.n514 VSUBS 0.007607f
C1381 B.n515 VSUBS 0.007607f
C1382 B.n516 VSUBS 0.007607f
C1383 B.n517 VSUBS 0.007607f
C1384 B.n518 VSUBS 0.007607f
C1385 B.n519 VSUBS 0.007607f
C1386 B.n520 VSUBS 0.007607f
C1387 B.n521 VSUBS 0.007607f
C1388 B.n522 VSUBS 0.007607f
C1389 B.n523 VSUBS 0.007607f
C1390 B.n524 VSUBS 0.007607f
C1391 B.n525 VSUBS 0.007607f
C1392 B.n526 VSUBS 0.007607f
C1393 B.n527 VSUBS 0.007607f
C1394 B.n528 VSUBS 0.007607f
C1395 B.n529 VSUBS 0.007607f
C1396 B.n530 VSUBS 0.007607f
C1397 B.n531 VSUBS 0.007607f
C1398 B.n532 VSUBS 0.007607f
C1399 B.n533 VSUBS 0.007607f
C1400 B.n534 VSUBS 0.007607f
C1401 B.n535 VSUBS 0.007607f
C1402 B.n536 VSUBS 0.007607f
C1403 B.n537 VSUBS 0.007607f
C1404 B.n538 VSUBS 0.007607f
C1405 B.n539 VSUBS 0.007607f
C1406 B.n540 VSUBS 0.007607f
C1407 B.n541 VSUBS 0.007607f
C1408 B.n542 VSUBS 0.007607f
C1409 B.n543 VSUBS 0.007607f
C1410 B.n544 VSUBS 0.007607f
C1411 B.n545 VSUBS 0.007607f
C1412 B.n546 VSUBS 0.007607f
C1413 B.n547 VSUBS 0.007607f
C1414 B.n548 VSUBS 0.007607f
C1415 B.n549 VSUBS 0.007607f
C1416 B.n550 VSUBS 0.007607f
C1417 B.n551 VSUBS 0.007607f
C1418 B.n552 VSUBS 0.007607f
C1419 B.n553 VSUBS 0.007607f
C1420 B.n554 VSUBS 0.007607f
C1421 B.n555 VSUBS 0.007607f
C1422 B.n556 VSUBS 0.005258f
C1423 B.n557 VSUBS 0.017624f
C1424 B.n558 VSUBS 0.006153f
C1425 B.n559 VSUBS 0.007607f
C1426 B.n560 VSUBS 0.007607f
C1427 B.n561 VSUBS 0.007607f
C1428 B.n562 VSUBS 0.007607f
C1429 B.n563 VSUBS 0.007607f
C1430 B.n564 VSUBS 0.007607f
C1431 B.n565 VSUBS 0.007607f
C1432 B.n566 VSUBS 0.007607f
C1433 B.n567 VSUBS 0.007607f
C1434 B.n568 VSUBS 0.007607f
C1435 B.n569 VSUBS 0.007607f
C1436 B.n570 VSUBS 0.006153f
C1437 B.n571 VSUBS 0.007607f
C1438 B.n572 VSUBS 0.007607f
C1439 B.n573 VSUBS 0.005258f
C1440 B.n574 VSUBS 0.007607f
C1441 B.n575 VSUBS 0.007607f
C1442 B.n576 VSUBS 0.007607f
C1443 B.n577 VSUBS 0.007607f
C1444 B.n578 VSUBS 0.007607f
C1445 B.n579 VSUBS 0.007607f
C1446 B.n580 VSUBS 0.007607f
C1447 B.n581 VSUBS 0.007607f
C1448 B.n582 VSUBS 0.007607f
C1449 B.n583 VSUBS 0.007607f
C1450 B.n584 VSUBS 0.007607f
C1451 B.n585 VSUBS 0.007607f
C1452 B.n586 VSUBS 0.007607f
C1453 B.n587 VSUBS 0.007607f
C1454 B.n588 VSUBS 0.007607f
C1455 B.n589 VSUBS 0.007607f
C1456 B.n590 VSUBS 0.007607f
C1457 B.n591 VSUBS 0.007607f
C1458 B.n592 VSUBS 0.007607f
C1459 B.n593 VSUBS 0.007607f
C1460 B.n594 VSUBS 0.007607f
C1461 B.n595 VSUBS 0.007607f
C1462 B.n596 VSUBS 0.007607f
C1463 B.n597 VSUBS 0.007607f
C1464 B.n598 VSUBS 0.007607f
C1465 B.n599 VSUBS 0.007607f
C1466 B.n600 VSUBS 0.007607f
C1467 B.n601 VSUBS 0.007607f
C1468 B.n602 VSUBS 0.007607f
C1469 B.n603 VSUBS 0.007607f
C1470 B.n604 VSUBS 0.007607f
C1471 B.n605 VSUBS 0.007607f
C1472 B.n606 VSUBS 0.007607f
C1473 B.n607 VSUBS 0.007607f
C1474 B.n608 VSUBS 0.007607f
C1475 B.n609 VSUBS 0.007607f
C1476 B.n610 VSUBS 0.007607f
C1477 B.n611 VSUBS 0.007607f
C1478 B.n612 VSUBS 0.007607f
C1479 B.n613 VSUBS 0.007607f
C1480 B.n614 VSUBS 0.007607f
C1481 B.n615 VSUBS 0.007607f
C1482 B.n616 VSUBS 0.007607f
C1483 B.n617 VSUBS 0.007607f
C1484 B.n618 VSUBS 0.007607f
C1485 B.n619 VSUBS 0.007607f
C1486 B.n620 VSUBS 0.007607f
C1487 B.n621 VSUBS 0.007607f
C1488 B.n622 VSUBS 0.007607f
C1489 B.n623 VSUBS 0.007607f
C1490 B.n624 VSUBS 0.007607f
C1491 B.n625 VSUBS 0.007607f
C1492 B.n626 VSUBS 0.007607f
C1493 B.n627 VSUBS 0.007607f
C1494 B.n628 VSUBS 0.007607f
C1495 B.n629 VSUBS 0.007607f
C1496 B.n630 VSUBS 0.007607f
C1497 B.n631 VSUBS 0.007607f
C1498 B.n632 VSUBS 0.007607f
C1499 B.n633 VSUBS 0.007607f
C1500 B.n634 VSUBS 0.007607f
C1501 B.n635 VSUBS 0.007607f
C1502 B.n636 VSUBS 0.007607f
C1503 B.n637 VSUBS 0.007607f
C1504 B.n638 VSUBS 0.007607f
C1505 B.n639 VSUBS 0.007607f
C1506 B.n640 VSUBS 0.007607f
C1507 B.n641 VSUBS 0.007607f
C1508 B.n642 VSUBS 0.007607f
C1509 B.n643 VSUBS 0.007607f
C1510 B.n644 VSUBS 0.007607f
C1511 B.n645 VSUBS 0.007607f
C1512 B.n646 VSUBS 0.007607f
C1513 B.n647 VSUBS 0.007607f
C1514 B.n648 VSUBS 0.007607f
C1515 B.n649 VSUBS 0.007607f
C1516 B.n650 VSUBS 0.007607f
C1517 B.n651 VSUBS 0.007607f
C1518 B.n652 VSUBS 0.007607f
C1519 B.n653 VSUBS 0.007607f
C1520 B.n654 VSUBS 0.007607f
C1521 B.n655 VSUBS 0.007607f
C1522 B.n656 VSUBS 0.007607f
C1523 B.n657 VSUBS 0.007607f
C1524 B.n658 VSUBS 0.007607f
C1525 B.n659 VSUBS 0.007607f
C1526 B.n660 VSUBS 0.007607f
C1527 B.n661 VSUBS 0.017723f
C1528 B.n662 VSUBS 0.016732f
C1529 B.n663 VSUBS 0.016732f
C1530 B.n664 VSUBS 0.007607f
C1531 B.n665 VSUBS 0.007607f
C1532 B.n666 VSUBS 0.007607f
C1533 B.n667 VSUBS 0.007607f
C1534 B.n668 VSUBS 0.007607f
C1535 B.n669 VSUBS 0.007607f
C1536 B.n670 VSUBS 0.007607f
C1537 B.n671 VSUBS 0.007607f
C1538 B.n672 VSUBS 0.007607f
C1539 B.n673 VSUBS 0.007607f
C1540 B.n674 VSUBS 0.007607f
C1541 B.n675 VSUBS 0.007607f
C1542 B.n676 VSUBS 0.007607f
C1543 B.n677 VSUBS 0.007607f
C1544 B.n678 VSUBS 0.007607f
C1545 B.n679 VSUBS 0.007607f
C1546 B.n680 VSUBS 0.007607f
C1547 B.n681 VSUBS 0.007607f
C1548 B.n682 VSUBS 0.007607f
C1549 B.n683 VSUBS 0.007607f
C1550 B.n684 VSUBS 0.007607f
C1551 B.n685 VSUBS 0.007607f
C1552 B.n686 VSUBS 0.007607f
C1553 B.n687 VSUBS 0.007607f
C1554 B.n688 VSUBS 0.007607f
C1555 B.n689 VSUBS 0.007607f
C1556 B.n690 VSUBS 0.007607f
C1557 B.n691 VSUBS 0.009926f
C1558 B.n692 VSUBS 0.010574f
C1559 B.n693 VSUBS 0.021028f
.ends

