* NGSPICE file created from diff_pair_sample_0841.ext - technology: sky130A

.subckt diff_pair_sample_0841 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=0 ps=0 w=2.57 l=3.88
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=0 ps=0 w=2.57 l=3.88
X2 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=1.0023 ps=5.92 w=2.57 l=3.88
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=0 ps=0 w=2.57 l=3.88
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=0 ps=0 w=2.57 l=3.88
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=1.0023 ps=5.92 w=2.57 l=3.88
X6 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=1.0023 ps=5.92 w=2.57 l=3.88
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0023 pd=5.92 as=1.0023 ps=5.92 w=2.57 l=3.88
R0 B.n463 B.n462 585
R1 B.n464 B.n463 585
R2 B.n158 B.n81 585
R3 B.n157 B.n156 585
R4 B.n155 B.n154 585
R5 B.n153 B.n152 585
R6 B.n151 B.n150 585
R7 B.n149 B.n148 585
R8 B.n147 B.n146 585
R9 B.n145 B.n144 585
R10 B.n143 B.n142 585
R11 B.n141 B.n140 585
R12 B.n139 B.n138 585
R13 B.n137 B.n136 585
R14 B.n135 B.n134 585
R15 B.n132 B.n131 585
R16 B.n130 B.n129 585
R17 B.n128 B.n127 585
R18 B.n126 B.n125 585
R19 B.n124 B.n123 585
R20 B.n122 B.n121 585
R21 B.n120 B.n119 585
R22 B.n118 B.n117 585
R23 B.n116 B.n115 585
R24 B.n114 B.n113 585
R25 B.n112 B.n111 585
R26 B.n110 B.n109 585
R27 B.n108 B.n107 585
R28 B.n106 B.n105 585
R29 B.n104 B.n103 585
R30 B.n102 B.n101 585
R31 B.n100 B.n99 585
R32 B.n98 B.n97 585
R33 B.n96 B.n95 585
R34 B.n94 B.n93 585
R35 B.n92 B.n91 585
R36 B.n90 B.n89 585
R37 B.n88 B.n87 585
R38 B.n461 B.n62 585
R39 B.n465 B.n62 585
R40 B.n460 B.n61 585
R41 B.n466 B.n61 585
R42 B.n459 B.n458 585
R43 B.n458 B.n57 585
R44 B.n457 B.n56 585
R45 B.n472 B.n56 585
R46 B.n456 B.n55 585
R47 B.n473 B.n55 585
R48 B.n455 B.n54 585
R49 B.n474 B.n54 585
R50 B.n454 B.n453 585
R51 B.n453 B.n50 585
R52 B.n452 B.n49 585
R53 B.n480 B.n49 585
R54 B.n451 B.n48 585
R55 B.n481 B.n48 585
R56 B.n450 B.n47 585
R57 B.n482 B.n47 585
R58 B.n449 B.n448 585
R59 B.n448 B.n43 585
R60 B.n447 B.n42 585
R61 B.n488 B.n42 585
R62 B.n446 B.n41 585
R63 B.n489 B.n41 585
R64 B.n445 B.n40 585
R65 B.n490 B.n40 585
R66 B.n444 B.n443 585
R67 B.n443 B.n36 585
R68 B.n442 B.n35 585
R69 B.n496 B.n35 585
R70 B.n441 B.n34 585
R71 B.n497 B.n34 585
R72 B.n440 B.n33 585
R73 B.n498 B.n33 585
R74 B.n439 B.n438 585
R75 B.n438 B.n29 585
R76 B.n437 B.n28 585
R77 B.n504 B.n28 585
R78 B.n436 B.n27 585
R79 B.n505 B.n27 585
R80 B.n435 B.n26 585
R81 B.n506 B.n26 585
R82 B.n434 B.n433 585
R83 B.n433 B.n22 585
R84 B.n432 B.n21 585
R85 B.n512 B.n21 585
R86 B.n431 B.n20 585
R87 B.n513 B.n20 585
R88 B.n430 B.n19 585
R89 B.n514 B.n19 585
R90 B.n429 B.n428 585
R91 B.n428 B.n15 585
R92 B.n427 B.n14 585
R93 B.n520 B.n14 585
R94 B.n426 B.n13 585
R95 B.n521 B.n13 585
R96 B.n425 B.n12 585
R97 B.n522 B.n12 585
R98 B.n424 B.n423 585
R99 B.n423 B.n8 585
R100 B.n422 B.n7 585
R101 B.n528 B.n7 585
R102 B.n421 B.n6 585
R103 B.n529 B.n6 585
R104 B.n420 B.n5 585
R105 B.n530 B.n5 585
R106 B.n419 B.n418 585
R107 B.n418 B.n4 585
R108 B.n417 B.n159 585
R109 B.n417 B.n416 585
R110 B.n407 B.n160 585
R111 B.n161 B.n160 585
R112 B.n409 B.n408 585
R113 B.n410 B.n409 585
R114 B.n406 B.n166 585
R115 B.n166 B.n165 585
R116 B.n405 B.n404 585
R117 B.n404 B.n403 585
R118 B.n168 B.n167 585
R119 B.n169 B.n168 585
R120 B.n396 B.n395 585
R121 B.n397 B.n396 585
R122 B.n394 B.n174 585
R123 B.n174 B.n173 585
R124 B.n393 B.n392 585
R125 B.n392 B.n391 585
R126 B.n176 B.n175 585
R127 B.n177 B.n176 585
R128 B.n384 B.n383 585
R129 B.n385 B.n384 585
R130 B.n382 B.n182 585
R131 B.n182 B.n181 585
R132 B.n381 B.n380 585
R133 B.n380 B.n379 585
R134 B.n184 B.n183 585
R135 B.n185 B.n184 585
R136 B.n372 B.n371 585
R137 B.n373 B.n372 585
R138 B.n370 B.n190 585
R139 B.n190 B.n189 585
R140 B.n369 B.n368 585
R141 B.n368 B.n367 585
R142 B.n192 B.n191 585
R143 B.n193 B.n192 585
R144 B.n360 B.n359 585
R145 B.n361 B.n360 585
R146 B.n358 B.n198 585
R147 B.n198 B.n197 585
R148 B.n357 B.n356 585
R149 B.n356 B.n355 585
R150 B.n200 B.n199 585
R151 B.n201 B.n200 585
R152 B.n348 B.n347 585
R153 B.n349 B.n348 585
R154 B.n346 B.n206 585
R155 B.n206 B.n205 585
R156 B.n345 B.n344 585
R157 B.n344 B.n343 585
R158 B.n208 B.n207 585
R159 B.n209 B.n208 585
R160 B.n336 B.n335 585
R161 B.n337 B.n336 585
R162 B.n334 B.n214 585
R163 B.n214 B.n213 585
R164 B.n333 B.n332 585
R165 B.n332 B.n331 585
R166 B.n216 B.n215 585
R167 B.n217 B.n216 585
R168 B.n324 B.n323 585
R169 B.n325 B.n324 585
R170 B.n322 B.n222 585
R171 B.n222 B.n221 585
R172 B.n316 B.n315 585
R173 B.n314 B.n242 585
R174 B.n313 B.n241 585
R175 B.n318 B.n241 585
R176 B.n312 B.n311 585
R177 B.n310 B.n309 585
R178 B.n308 B.n307 585
R179 B.n306 B.n305 585
R180 B.n304 B.n303 585
R181 B.n302 B.n301 585
R182 B.n300 B.n299 585
R183 B.n298 B.n297 585
R184 B.n296 B.n295 585
R185 B.n294 B.n293 585
R186 B.n292 B.n291 585
R187 B.n289 B.n288 585
R188 B.n287 B.n286 585
R189 B.n285 B.n284 585
R190 B.n283 B.n282 585
R191 B.n281 B.n280 585
R192 B.n279 B.n278 585
R193 B.n277 B.n276 585
R194 B.n275 B.n274 585
R195 B.n273 B.n272 585
R196 B.n271 B.n270 585
R197 B.n269 B.n268 585
R198 B.n267 B.n266 585
R199 B.n265 B.n264 585
R200 B.n263 B.n262 585
R201 B.n261 B.n260 585
R202 B.n259 B.n258 585
R203 B.n257 B.n256 585
R204 B.n255 B.n254 585
R205 B.n253 B.n252 585
R206 B.n251 B.n250 585
R207 B.n249 B.n248 585
R208 B.n224 B.n223 585
R209 B.n321 B.n320 585
R210 B.n220 B.n219 585
R211 B.n221 B.n220 585
R212 B.n327 B.n326 585
R213 B.n326 B.n325 585
R214 B.n328 B.n218 585
R215 B.n218 B.n217 585
R216 B.n330 B.n329 585
R217 B.n331 B.n330 585
R218 B.n212 B.n211 585
R219 B.n213 B.n212 585
R220 B.n339 B.n338 585
R221 B.n338 B.n337 585
R222 B.n340 B.n210 585
R223 B.n210 B.n209 585
R224 B.n342 B.n341 585
R225 B.n343 B.n342 585
R226 B.n204 B.n203 585
R227 B.n205 B.n204 585
R228 B.n351 B.n350 585
R229 B.n350 B.n349 585
R230 B.n352 B.n202 585
R231 B.n202 B.n201 585
R232 B.n354 B.n353 585
R233 B.n355 B.n354 585
R234 B.n196 B.n195 585
R235 B.n197 B.n196 585
R236 B.n363 B.n362 585
R237 B.n362 B.n361 585
R238 B.n364 B.n194 585
R239 B.n194 B.n193 585
R240 B.n366 B.n365 585
R241 B.n367 B.n366 585
R242 B.n188 B.n187 585
R243 B.n189 B.n188 585
R244 B.n375 B.n374 585
R245 B.n374 B.n373 585
R246 B.n376 B.n186 585
R247 B.n186 B.n185 585
R248 B.n378 B.n377 585
R249 B.n379 B.n378 585
R250 B.n180 B.n179 585
R251 B.n181 B.n180 585
R252 B.n387 B.n386 585
R253 B.n386 B.n385 585
R254 B.n388 B.n178 585
R255 B.n178 B.n177 585
R256 B.n390 B.n389 585
R257 B.n391 B.n390 585
R258 B.n172 B.n171 585
R259 B.n173 B.n172 585
R260 B.n399 B.n398 585
R261 B.n398 B.n397 585
R262 B.n400 B.n170 585
R263 B.n170 B.n169 585
R264 B.n402 B.n401 585
R265 B.n403 B.n402 585
R266 B.n164 B.n163 585
R267 B.n165 B.n164 585
R268 B.n412 B.n411 585
R269 B.n411 B.n410 585
R270 B.n413 B.n162 585
R271 B.n162 B.n161 585
R272 B.n415 B.n414 585
R273 B.n416 B.n415 585
R274 B.n2 B.n0 585
R275 B.n4 B.n2 585
R276 B.n3 B.n1 585
R277 B.n529 B.n3 585
R278 B.n527 B.n526 585
R279 B.n528 B.n527 585
R280 B.n525 B.n9 585
R281 B.n9 B.n8 585
R282 B.n524 B.n523 585
R283 B.n523 B.n522 585
R284 B.n11 B.n10 585
R285 B.n521 B.n11 585
R286 B.n519 B.n518 585
R287 B.n520 B.n519 585
R288 B.n517 B.n16 585
R289 B.n16 B.n15 585
R290 B.n516 B.n515 585
R291 B.n515 B.n514 585
R292 B.n18 B.n17 585
R293 B.n513 B.n18 585
R294 B.n511 B.n510 585
R295 B.n512 B.n511 585
R296 B.n509 B.n23 585
R297 B.n23 B.n22 585
R298 B.n508 B.n507 585
R299 B.n507 B.n506 585
R300 B.n25 B.n24 585
R301 B.n505 B.n25 585
R302 B.n503 B.n502 585
R303 B.n504 B.n503 585
R304 B.n501 B.n30 585
R305 B.n30 B.n29 585
R306 B.n500 B.n499 585
R307 B.n499 B.n498 585
R308 B.n32 B.n31 585
R309 B.n497 B.n32 585
R310 B.n495 B.n494 585
R311 B.n496 B.n495 585
R312 B.n493 B.n37 585
R313 B.n37 B.n36 585
R314 B.n492 B.n491 585
R315 B.n491 B.n490 585
R316 B.n39 B.n38 585
R317 B.n489 B.n39 585
R318 B.n487 B.n486 585
R319 B.n488 B.n487 585
R320 B.n485 B.n44 585
R321 B.n44 B.n43 585
R322 B.n484 B.n483 585
R323 B.n483 B.n482 585
R324 B.n46 B.n45 585
R325 B.n481 B.n46 585
R326 B.n479 B.n478 585
R327 B.n480 B.n479 585
R328 B.n477 B.n51 585
R329 B.n51 B.n50 585
R330 B.n476 B.n475 585
R331 B.n475 B.n474 585
R332 B.n53 B.n52 585
R333 B.n473 B.n53 585
R334 B.n471 B.n470 585
R335 B.n472 B.n471 585
R336 B.n469 B.n58 585
R337 B.n58 B.n57 585
R338 B.n468 B.n467 585
R339 B.n467 B.n466 585
R340 B.n60 B.n59 585
R341 B.n465 B.n60 585
R342 B.n532 B.n531 585
R343 B.n531 B.n530 585
R344 B.n316 B.n220 506.916
R345 B.n87 B.n60 506.916
R346 B.n320 B.n222 506.916
R347 B.n463 B.n62 506.916
R348 B.n464 B.n80 256.663
R349 B.n464 B.n79 256.663
R350 B.n464 B.n78 256.663
R351 B.n464 B.n77 256.663
R352 B.n464 B.n76 256.663
R353 B.n464 B.n75 256.663
R354 B.n464 B.n74 256.663
R355 B.n464 B.n73 256.663
R356 B.n464 B.n72 256.663
R357 B.n464 B.n71 256.663
R358 B.n464 B.n70 256.663
R359 B.n464 B.n69 256.663
R360 B.n464 B.n68 256.663
R361 B.n464 B.n67 256.663
R362 B.n464 B.n66 256.663
R363 B.n464 B.n65 256.663
R364 B.n464 B.n64 256.663
R365 B.n464 B.n63 256.663
R366 B.n318 B.n317 256.663
R367 B.n318 B.n225 256.663
R368 B.n318 B.n226 256.663
R369 B.n318 B.n227 256.663
R370 B.n318 B.n228 256.663
R371 B.n318 B.n229 256.663
R372 B.n318 B.n230 256.663
R373 B.n318 B.n231 256.663
R374 B.n318 B.n232 256.663
R375 B.n318 B.n233 256.663
R376 B.n318 B.n234 256.663
R377 B.n318 B.n235 256.663
R378 B.n318 B.n236 256.663
R379 B.n318 B.n237 256.663
R380 B.n318 B.n238 256.663
R381 B.n318 B.n239 256.663
R382 B.n318 B.n240 256.663
R383 B.n319 B.n318 256.663
R384 B.n245 B.t10 225.368
R385 B.n243 B.t2 225.368
R386 B.n84 B.t6 225.368
R387 B.n82 B.t13 225.368
R388 B.n245 B.t12 205.706
R389 B.n82 B.t14 205.706
R390 B.n243 B.t5 205.706
R391 B.n84 B.t8 205.706
R392 B.n326 B.n220 163.367
R393 B.n326 B.n218 163.367
R394 B.n330 B.n218 163.367
R395 B.n330 B.n212 163.367
R396 B.n338 B.n212 163.367
R397 B.n338 B.n210 163.367
R398 B.n342 B.n210 163.367
R399 B.n342 B.n204 163.367
R400 B.n350 B.n204 163.367
R401 B.n350 B.n202 163.367
R402 B.n354 B.n202 163.367
R403 B.n354 B.n196 163.367
R404 B.n362 B.n196 163.367
R405 B.n362 B.n194 163.367
R406 B.n366 B.n194 163.367
R407 B.n366 B.n188 163.367
R408 B.n374 B.n188 163.367
R409 B.n374 B.n186 163.367
R410 B.n378 B.n186 163.367
R411 B.n378 B.n180 163.367
R412 B.n386 B.n180 163.367
R413 B.n386 B.n178 163.367
R414 B.n390 B.n178 163.367
R415 B.n390 B.n172 163.367
R416 B.n398 B.n172 163.367
R417 B.n398 B.n170 163.367
R418 B.n402 B.n170 163.367
R419 B.n402 B.n164 163.367
R420 B.n411 B.n164 163.367
R421 B.n411 B.n162 163.367
R422 B.n415 B.n162 163.367
R423 B.n415 B.n2 163.367
R424 B.n531 B.n2 163.367
R425 B.n531 B.n3 163.367
R426 B.n527 B.n3 163.367
R427 B.n527 B.n9 163.367
R428 B.n523 B.n9 163.367
R429 B.n523 B.n11 163.367
R430 B.n519 B.n11 163.367
R431 B.n519 B.n16 163.367
R432 B.n515 B.n16 163.367
R433 B.n515 B.n18 163.367
R434 B.n511 B.n18 163.367
R435 B.n511 B.n23 163.367
R436 B.n507 B.n23 163.367
R437 B.n507 B.n25 163.367
R438 B.n503 B.n25 163.367
R439 B.n503 B.n30 163.367
R440 B.n499 B.n30 163.367
R441 B.n499 B.n32 163.367
R442 B.n495 B.n32 163.367
R443 B.n495 B.n37 163.367
R444 B.n491 B.n37 163.367
R445 B.n491 B.n39 163.367
R446 B.n487 B.n39 163.367
R447 B.n487 B.n44 163.367
R448 B.n483 B.n44 163.367
R449 B.n483 B.n46 163.367
R450 B.n479 B.n46 163.367
R451 B.n479 B.n51 163.367
R452 B.n475 B.n51 163.367
R453 B.n475 B.n53 163.367
R454 B.n471 B.n53 163.367
R455 B.n471 B.n58 163.367
R456 B.n467 B.n58 163.367
R457 B.n467 B.n60 163.367
R458 B.n242 B.n241 163.367
R459 B.n311 B.n241 163.367
R460 B.n309 B.n308 163.367
R461 B.n305 B.n304 163.367
R462 B.n301 B.n300 163.367
R463 B.n297 B.n296 163.367
R464 B.n293 B.n292 163.367
R465 B.n288 B.n287 163.367
R466 B.n284 B.n283 163.367
R467 B.n280 B.n279 163.367
R468 B.n276 B.n275 163.367
R469 B.n272 B.n271 163.367
R470 B.n268 B.n267 163.367
R471 B.n264 B.n263 163.367
R472 B.n260 B.n259 163.367
R473 B.n256 B.n255 163.367
R474 B.n252 B.n251 163.367
R475 B.n248 B.n224 163.367
R476 B.n324 B.n222 163.367
R477 B.n324 B.n216 163.367
R478 B.n332 B.n216 163.367
R479 B.n332 B.n214 163.367
R480 B.n336 B.n214 163.367
R481 B.n336 B.n208 163.367
R482 B.n344 B.n208 163.367
R483 B.n344 B.n206 163.367
R484 B.n348 B.n206 163.367
R485 B.n348 B.n200 163.367
R486 B.n356 B.n200 163.367
R487 B.n356 B.n198 163.367
R488 B.n360 B.n198 163.367
R489 B.n360 B.n192 163.367
R490 B.n368 B.n192 163.367
R491 B.n368 B.n190 163.367
R492 B.n372 B.n190 163.367
R493 B.n372 B.n184 163.367
R494 B.n380 B.n184 163.367
R495 B.n380 B.n182 163.367
R496 B.n384 B.n182 163.367
R497 B.n384 B.n176 163.367
R498 B.n392 B.n176 163.367
R499 B.n392 B.n174 163.367
R500 B.n396 B.n174 163.367
R501 B.n396 B.n168 163.367
R502 B.n404 B.n168 163.367
R503 B.n404 B.n166 163.367
R504 B.n409 B.n166 163.367
R505 B.n409 B.n160 163.367
R506 B.n417 B.n160 163.367
R507 B.n418 B.n417 163.367
R508 B.n418 B.n5 163.367
R509 B.n6 B.n5 163.367
R510 B.n7 B.n6 163.367
R511 B.n423 B.n7 163.367
R512 B.n423 B.n12 163.367
R513 B.n13 B.n12 163.367
R514 B.n14 B.n13 163.367
R515 B.n428 B.n14 163.367
R516 B.n428 B.n19 163.367
R517 B.n20 B.n19 163.367
R518 B.n21 B.n20 163.367
R519 B.n433 B.n21 163.367
R520 B.n433 B.n26 163.367
R521 B.n27 B.n26 163.367
R522 B.n28 B.n27 163.367
R523 B.n438 B.n28 163.367
R524 B.n438 B.n33 163.367
R525 B.n34 B.n33 163.367
R526 B.n35 B.n34 163.367
R527 B.n443 B.n35 163.367
R528 B.n443 B.n40 163.367
R529 B.n41 B.n40 163.367
R530 B.n42 B.n41 163.367
R531 B.n448 B.n42 163.367
R532 B.n448 B.n47 163.367
R533 B.n48 B.n47 163.367
R534 B.n49 B.n48 163.367
R535 B.n453 B.n49 163.367
R536 B.n453 B.n54 163.367
R537 B.n55 B.n54 163.367
R538 B.n56 B.n55 163.367
R539 B.n458 B.n56 163.367
R540 B.n458 B.n61 163.367
R541 B.n62 B.n61 163.367
R542 B.n91 B.n90 163.367
R543 B.n95 B.n94 163.367
R544 B.n99 B.n98 163.367
R545 B.n103 B.n102 163.367
R546 B.n107 B.n106 163.367
R547 B.n111 B.n110 163.367
R548 B.n115 B.n114 163.367
R549 B.n119 B.n118 163.367
R550 B.n123 B.n122 163.367
R551 B.n127 B.n126 163.367
R552 B.n131 B.n130 163.367
R553 B.n136 B.n135 163.367
R554 B.n140 B.n139 163.367
R555 B.n144 B.n143 163.367
R556 B.n148 B.n147 163.367
R557 B.n152 B.n151 163.367
R558 B.n156 B.n155 163.367
R559 B.n463 B.n81 163.367
R560 B.n318 B.n221 161.25
R561 B.n465 B.n464 161.25
R562 B.n246 B.t11 124.056
R563 B.n83 B.t15 124.056
R564 B.n244 B.t4 124.056
R565 B.n85 B.t9 124.056
R566 B.n325 B.n221 95.3479
R567 B.n325 B.n217 95.3479
R568 B.n331 B.n217 95.3479
R569 B.n331 B.n213 95.3479
R570 B.n337 B.n213 95.3479
R571 B.n337 B.n209 95.3479
R572 B.n343 B.n209 95.3479
R573 B.n343 B.n205 95.3479
R574 B.n349 B.n205 95.3479
R575 B.n355 B.n201 95.3479
R576 B.n355 B.n197 95.3479
R577 B.n361 B.n197 95.3479
R578 B.n361 B.n193 95.3479
R579 B.n367 B.n193 95.3479
R580 B.n367 B.n189 95.3479
R581 B.n373 B.n189 95.3479
R582 B.n373 B.n185 95.3479
R583 B.n379 B.n185 95.3479
R584 B.n379 B.n181 95.3479
R585 B.n385 B.n181 95.3479
R586 B.n385 B.n177 95.3479
R587 B.n391 B.n177 95.3479
R588 B.n391 B.n173 95.3479
R589 B.n397 B.n173 95.3479
R590 B.n403 B.n169 95.3479
R591 B.n403 B.n165 95.3479
R592 B.n410 B.n165 95.3479
R593 B.n410 B.n161 95.3479
R594 B.n416 B.n161 95.3479
R595 B.n416 B.n4 95.3479
R596 B.n530 B.n4 95.3479
R597 B.n530 B.n529 95.3479
R598 B.n529 B.n528 95.3479
R599 B.n528 B.n8 95.3479
R600 B.n522 B.n8 95.3479
R601 B.n522 B.n521 95.3479
R602 B.n521 B.n520 95.3479
R603 B.n520 B.n15 95.3479
R604 B.n514 B.n513 95.3479
R605 B.n513 B.n512 95.3479
R606 B.n512 B.n22 95.3479
R607 B.n506 B.n22 95.3479
R608 B.n506 B.n505 95.3479
R609 B.n505 B.n504 95.3479
R610 B.n504 B.n29 95.3479
R611 B.n498 B.n29 95.3479
R612 B.n498 B.n497 95.3479
R613 B.n497 B.n496 95.3479
R614 B.n496 B.n36 95.3479
R615 B.n490 B.n36 95.3479
R616 B.n490 B.n489 95.3479
R617 B.n489 B.n488 95.3479
R618 B.n488 B.n43 95.3479
R619 B.n482 B.n481 95.3479
R620 B.n481 B.n480 95.3479
R621 B.n480 B.n50 95.3479
R622 B.n474 B.n50 95.3479
R623 B.n474 B.n473 95.3479
R624 B.n473 B.n472 95.3479
R625 B.n472 B.n57 95.3479
R626 B.n466 B.n57 95.3479
R627 B.n466 B.n465 95.3479
R628 B.n246 B.n245 81.649
R629 B.n244 B.n243 81.649
R630 B.n85 B.n84 81.649
R631 B.n83 B.n82 81.649
R632 B.t1 B.n169 75.7175
R633 B.t0 B.n15 75.7175
R634 B.n317 B.n316 71.676
R635 B.n311 B.n225 71.676
R636 B.n308 B.n226 71.676
R637 B.n304 B.n227 71.676
R638 B.n300 B.n228 71.676
R639 B.n296 B.n229 71.676
R640 B.n292 B.n230 71.676
R641 B.n287 B.n231 71.676
R642 B.n283 B.n232 71.676
R643 B.n279 B.n233 71.676
R644 B.n275 B.n234 71.676
R645 B.n271 B.n235 71.676
R646 B.n267 B.n236 71.676
R647 B.n263 B.n237 71.676
R648 B.n259 B.n238 71.676
R649 B.n255 B.n239 71.676
R650 B.n251 B.n240 71.676
R651 B.n319 B.n224 71.676
R652 B.n87 B.n63 71.676
R653 B.n91 B.n64 71.676
R654 B.n95 B.n65 71.676
R655 B.n99 B.n66 71.676
R656 B.n103 B.n67 71.676
R657 B.n107 B.n68 71.676
R658 B.n111 B.n69 71.676
R659 B.n115 B.n70 71.676
R660 B.n119 B.n71 71.676
R661 B.n123 B.n72 71.676
R662 B.n127 B.n73 71.676
R663 B.n131 B.n74 71.676
R664 B.n136 B.n75 71.676
R665 B.n140 B.n76 71.676
R666 B.n144 B.n77 71.676
R667 B.n148 B.n78 71.676
R668 B.n152 B.n79 71.676
R669 B.n156 B.n80 71.676
R670 B.n81 B.n80 71.676
R671 B.n155 B.n79 71.676
R672 B.n151 B.n78 71.676
R673 B.n147 B.n77 71.676
R674 B.n143 B.n76 71.676
R675 B.n139 B.n75 71.676
R676 B.n135 B.n74 71.676
R677 B.n130 B.n73 71.676
R678 B.n126 B.n72 71.676
R679 B.n122 B.n71 71.676
R680 B.n118 B.n70 71.676
R681 B.n114 B.n69 71.676
R682 B.n110 B.n68 71.676
R683 B.n106 B.n67 71.676
R684 B.n102 B.n66 71.676
R685 B.n98 B.n65 71.676
R686 B.n94 B.n64 71.676
R687 B.n90 B.n63 71.676
R688 B.n317 B.n242 71.676
R689 B.n309 B.n225 71.676
R690 B.n305 B.n226 71.676
R691 B.n301 B.n227 71.676
R692 B.n297 B.n228 71.676
R693 B.n293 B.n229 71.676
R694 B.n288 B.n230 71.676
R695 B.n284 B.n231 71.676
R696 B.n280 B.n232 71.676
R697 B.n276 B.n233 71.676
R698 B.n272 B.n234 71.676
R699 B.n268 B.n235 71.676
R700 B.n264 B.n236 71.676
R701 B.n260 B.n237 71.676
R702 B.n256 B.n238 71.676
R703 B.n252 B.n239 71.676
R704 B.n248 B.n240 71.676
R705 B.n320 B.n319 71.676
R706 B.n247 B.n246 59.5399
R707 B.n290 B.n244 59.5399
R708 B.n86 B.n85 59.5399
R709 B.n133 B.n83 59.5399
R710 B.n349 B.t3 58.8915
R711 B.n482 B.t7 58.8915
R712 B.t3 B.n201 36.4568
R713 B.t7 B.n43 36.4568
R714 B.n88 B.n59 32.9371
R715 B.n462 B.n461 32.9371
R716 B.n322 B.n321 32.9371
R717 B.n315 B.n219 32.9371
R718 B.n397 B.t1 19.6308
R719 B.n514 B.t0 19.6308
R720 B B.n532 18.0485
R721 B.n89 B.n88 10.6151
R722 B.n92 B.n89 10.6151
R723 B.n93 B.n92 10.6151
R724 B.n96 B.n93 10.6151
R725 B.n97 B.n96 10.6151
R726 B.n100 B.n97 10.6151
R727 B.n101 B.n100 10.6151
R728 B.n104 B.n101 10.6151
R729 B.n105 B.n104 10.6151
R730 B.n108 B.n105 10.6151
R731 B.n109 B.n108 10.6151
R732 B.n112 B.n109 10.6151
R733 B.n113 B.n112 10.6151
R734 B.n117 B.n116 10.6151
R735 B.n120 B.n117 10.6151
R736 B.n121 B.n120 10.6151
R737 B.n124 B.n121 10.6151
R738 B.n125 B.n124 10.6151
R739 B.n128 B.n125 10.6151
R740 B.n129 B.n128 10.6151
R741 B.n132 B.n129 10.6151
R742 B.n137 B.n134 10.6151
R743 B.n138 B.n137 10.6151
R744 B.n141 B.n138 10.6151
R745 B.n142 B.n141 10.6151
R746 B.n145 B.n142 10.6151
R747 B.n146 B.n145 10.6151
R748 B.n149 B.n146 10.6151
R749 B.n150 B.n149 10.6151
R750 B.n153 B.n150 10.6151
R751 B.n154 B.n153 10.6151
R752 B.n157 B.n154 10.6151
R753 B.n158 B.n157 10.6151
R754 B.n462 B.n158 10.6151
R755 B.n323 B.n322 10.6151
R756 B.n323 B.n215 10.6151
R757 B.n333 B.n215 10.6151
R758 B.n334 B.n333 10.6151
R759 B.n335 B.n334 10.6151
R760 B.n335 B.n207 10.6151
R761 B.n345 B.n207 10.6151
R762 B.n346 B.n345 10.6151
R763 B.n347 B.n346 10.6151
R764 B.n347 B.n199 10.6151
R765 B.n357 B.n199 10.6151
R766 B.n358 B.n357 10.6151
R767 B.n359 B.n358 10.6151
R768 B.n359 B.n191 10.6151
R769 B.n369 B.n191 10.6151
R770 B.n370 B.n369 10.6151
R771 B.n371 B.n370 10.6151
R772 B.n371 B.n183 10.6151
R773 B.n381 B.n183 10.6151
R774 B.n382 B.n381 10.6151
R775 B.n383 B.n382 10.6151
R776 B.n383 B.n175 10.6151
R777 B.n393 B.n175 10.6151
R778 B.n394 B.n393 10.6151
R779 B.n395 B.n394 10.6151
R780 B.n395 B.n167 10.6151
R781 B.n405 B.n167 10.6151
R782 B.n406 B.n405 10.6151
R783 B.n408 B.n406 10.6151
R784 B.n408 B.n407 10.6151
R785 B.n407 B.n159 10.6151
R786 B.n419 B.n159 10.6151
R787 B.n420 B.n419 10.6151
R788 B.n421 B.n420 10.6151
R789 B.n422 B.n421 10.6151
R790 B.n424 B.n422 10.6151
R791 B.n425 B.n424 10.6151
R792 B.n426 B.n425 10.6151
R793 B.n427 B.n426 10.6151
R794 B.n429 B.n427 10.6151
R795 B.n430 B.n429 10.6151
R796 B.n431 B.n430 10.6151
R797 B.n432 B.n431 10.6151
R798 B.n434 B.n432 10.6151
R799 B.n435 B.n434 10.6151
R800 B.n436 B.n435 10.6151
R801 B.n437 B.n436 10.6151
R802 B.n439 B.n437 10.6151
R803 B.n440 B.n439 10.6151
R804 B.n441 B.n440 10.6151
R805 B.n442 B.n441 10.6151
R806 B.n444 B.n442 10.6151
R807 B.n445 B.n444 10.6151
R808 B.n446 B.n445 10.6151
R809 B.n447 B.n446 10.6151
R810 B.n449 B.n447 10.6151
R811 B.n450 B.n449 10.6151
R812 B.n451 B.n450 10.6151
R813 B.n452 B.n451 10.6151
R814 B.n454 B.n452 10.6151
R815 B.n455 B.n454 10.6151
R816 B.n456 B.n455 10.6151
R817 B.n457 B.n456 10.6151
R818 B.n459 B.n457 10.6151
R819 B.n460 B.n459 10.6151
R820 B.n461 B.n460 10.6151
R821 B.n315 B.n314 10.6151
R822 B.n314 B.n313 10.6151
R823 B.n313 B.n312 10.6151
R824 B.n312 B.n310 10.6151
R825 B.n310 B.n307 10.6151
R826 B.n307 B.n306 10.6151
R827 B.n306 B.n303 10.6151
R828 B.n303 B.n302 10.6151
R829 B.n302 B.n299 10.6151
R830 B.n299 B.n298 10.6151
R831 B.n298 B.n295 10.6151
R832 B.n295 B.n294 10.6151
R833 B.n294 B.n291 10.6151
R834 B.n289 B.n286 10.6151
R835 B.n286 B.n285 10.6151
R836 B.n285 B.n282 10.6151
R837 B.n282 B.n281 10.6151
R838 B.n281 B.n278 10.6151
R839 B.n278 B.n277 10.6151
R840 B.n277 B.n274 10.6151
R841 B.n274 B.n273 10.6151
R842 B.n270 B.n269 10.6151
R843 B.n269 B.n266 10.6151
R844 B.n266 B.n265 10.6151
R845 B.n265 B.n262 10.6151
R846 B.n262 B.n261 10.6151
R847 B.n261 B.n258 10.6151
R848 B.n258 B.n257 10.6151
R849 B.n257 B.n254 10.6151
R850 B.n254 B.n253 10.6151
R851 B.n253 B.n250 10.6151
R852 B.n250 B.n249 10.6151
R853 B.n249 B.n223 10.6151
R854 B.n321 B.n223 10.6151
R855 B.n327 B.n219 10.6151
R856 B.n328 B.n327 10.6151
R857 B.n329 B.n328 10.6151
R858 B.n329 B.n211 10.6151
R859 B.n339 B.n211 10.6151
R860 B.n340 B.n339 10.6151
R861 B.n341 B.n340 10.6151
R862 B.n341 B.n203 10.6151
R863 B.n351 B.n203 10.6151
R864 B.n352 B.n351 10.6151
R865 B.n353 B.n352 10.6151
R866 B.n353 B.n195 10.6151
R867 B.n363 B.n195 10.6151
R868 B.n364 B.n363 10.6151
R869 B.n365 B.n364 10.6151
R870 B.n365 B.n187 10.6151
R871 B.n375 B.n187 10.6151
R872 B.n376 B.n375 10.6151
R873 B.n377 B.n376 10.6151
R874 B.n377 B.n179 10.6151
R875 B.n387 B.n179 10.6151
R876 B.n388 B.n387 10.6151
R877 B.n389 B.n388 10.6151
R878 B.n389 B.n171 10.6151
R879 B.n399 B.n171 10.6151
R880 B.n400 B.n399 10.6151
R881 B.n401 B.n400 10.6151
R882 B.n401 B.n163 10.6151
R883 B.n412 B.n163 10.6151
R884 B.n413 B.n412 10.6151
R885 B.n414 B.n413 10.6151
R886 B.n414 B.n0 10.6151
R887 B.n526 B.n1 10.6151
R888 B.n526 B.n525 10.6151
R889 B.n525 B.n524 10.6151
R890 B.n524 B.n10 10.6151
R891 B.n518 B.n10 10.6151
R892 B.n518 B.n517 10.6151
R893 B.n517 B.n516 10.6151
R894 B.n516 B.n17 10.6151
R895 B.n510 B.n17 10.6151
R896 B.n510 B.n509 10.6151
R897 B.n509 B.n508 10.6151
R898 B.n508 B.n24 10.6151
R899 B.n502 B.n24 10.6151
R900 B.n502 B.n501 10.6151
R901 B.n501 B.n500 10.6151
R902 B.n500 B.n31 10.6151
R903 B.n494 B.n31 10.6151
R904 B.n494 B.n493 10.6151
R905 B.n493 B.n492 10.6151
R906 B.n492 B.n38 10.6151
R907 B.n486 B.n38 10.6151
R908 B.n486 B.n485 10.6151
R909 B.n485 B.n484 10.6151
R910 B.n484 B.n45 10.6151
R911 B.n478 B.n45 10.6151
R912 B.n478 B.n477 10.6151
R913 B.n477 B.n476 10.6151
R914 B.n476 B.n52 10.6151
R915 B.n470 B.n52 10.6151
R916 B.n470 B.n469 10.6151
R917 B.n469 B.n468 10.6151
R918 B.n468 B.n59 10.6151
R919 B.n116 B.n86 6.5566
R920 B.n133 B.n132 6.5566
R921 B.n290 B.n289 6.5566
R922 B.n273 B.n247 6.5566
R923 B.n113 B.n86 4.05904
R924 B.n134 B.n133 4.05904
R925 B.n291 B.n290 4.05904
R926 B.n270 B.n247 4.05904
R927 B.n532 B.n0 2.81026
R928 B.n532 B.n1 2.81026
R929 VN VN.t1 91.72
R930 VN VN.t0 51.6215
R931 VTAIL.n42 VTAIL.n36 289.615
R932 VTAIL.n6 VTAIL.n0 289.615
R933 VTAIL.n30 VTAIL.n24 289.615
R934 VTAIL.n18 VTAIL.n12 289.615
R935 VTAIL.n41 VTAIL.n40 185
R936 VTAIL.n43 VTAIL.n42 185
R937 VTAIL.n5 VTAIL.n4 185
R938 VTAIL.n7 VTAIL.n6 185
R939 VTAIL.n31 VTAIL.n30 185
R940 VTAIL.n29 VTAIL.n28 185
R941 VTAIL.n19 VTAIL.n18 185
R942 VTAIL.n17 VTAIL.n16 185
R943 VTAIL.n39 VTAIL.t2 151.613
R944 VTAIL.n3 VTAIL.t1 151.613
R945 VTAIL.n27 VTAIL.t0 151.613
R946 VTAIL.n15 VTAIL.t3 151.613
R947 VTAIL.n42 VTAIL.n41 104.615
R948 VTAIL.n6 VTAIL.n5 104.615
R949 VTAIL.n30 VTAIL.n29 104.615
R950 VTAIL.n18 VTAIL.n17 104.615
R951 VTAIL.n41 VTAIL.t2 52.3082
R952 VTAIL.n5 VTAIL.t1 52.3082
R953 VTAIL.n29 VTAIL.t0 52.3082
R954 VTAIL.n17 VTAIL.t3 52.3082
R955 VTAIL.n47 VTAIL.n46 35.4823
R956 VTAIL.n11 VTAIL.n10 35.4823
R957 VTAIL.n35 VTAIL.n34 35.4823
R958 VTAIL.n23 VTAIL.n22 35.4823
R959 VTAIL.n23 VTAIL.n11 21.841
R960 VTAIL.n47 VTAIL.n35 18.2117
R961 VTAIL.n40 VTAIL.n39 15.3979
R962 VTAIL.n4 VTAIL.n3 15.3979
R963 VTAIL.n28 VTAIL.n27 15.3979
R964 VTAIL.n16 VTAIL.n15 15.3979
R965 VTAIL.n43 VTAIL.n38 12.8005
R966 VTAIL.n7 VTAIL.n2 12.8005
R967 VTAIL.n31 VTAIL.n26 12.8005
R968 VTAIL.n19 VTAIL.n14 12.8005
R969 VTAIL.n44 VTAIL.n36 12.0247
R970 VTAIL.n8 VTAIL.n0 12.0247
R971 VTAIL.n32 VTAIL.n24 12.0247
R972 VTAIL.n20 VTAIL.n12 12.0247
R973 VTAIL.n46 VTAIL.n45 9.45567
R974 VTAIL.n10 VTAIL.n9 9.45567
R975 VTAIL.n34 VTAIL.n33 9.45567
R976 VTAIL.n22 VTAIL.n21 9.45567
R977 VTAIL.n45 VTAIL.n44 9.3005
R978 VTAIL.n38 VTAIL.n37 9.3005
R979 VTAIL.n9 VTAIL.n8 9.3005
R980 VTAIL.n2 VTAIL.n1 9.3005
R981 VTAIL.n33 VTAIL.n32 9.3005
R982 VTAIL.n26 VTAIL.n25 9.3005
R983 VTAIL.n21 VTAIL.n20 9.3005
R984 VTAIL.n14 VTAIL.n13 9.3005
R985 VTAIL.n39 VTAIL.n37 4.69785
R986 VTAIL.n3 VTAIL.n1 4.69785
R987 VTAIL.n27 VTAIL.n25 4.69785
R988 VTAIL.n15 VTAIL.n13 4.69785
R989 VTAIL.n35 VTAIL.n23 2.28498
R990 VTAIL.n46 VTAIL.n36 1.93989
R991 VTAIL.n10 VTAIL.n0 1.93989
R992 VTAIL.n34 VTAIL.n24 1.93989
R993 VTAIL.n22 VTAIL.n12 1.93989
R994 VTAIL VTAIL.n11 1.43584
R995 VTAIL.n44 VTAIL.n43 1.16414
R996 VTAIL.n8 VTAIL.n7 1.16414
R997 VTAIL.n32 VTAIL.n31 1.16414
R998 VTAIL.n20 VTAIL.n19 1.16414
R999 VTAIL VTAIL.n47 0.849638
R1000 VTAIL.n40 VTAIL.n38 0.388379
R1001 VTAIL.n4 VTAIL.n2 0.388379
R1002 VTAIL.n28 VTAIL.n26 0.388379
R1003 VTAIL.n16 VTAIL.n14 0.388379
R1004 VTAIL.n45 VTAIL.n37 0.155672
R1005 VTAIL.n9 VTAIL.n1 0.155672
R1006 VTAIL.n33 VTAIL.n25 0.155672
R1007 VTAIL.n21 VTAIL.n13 0.155672
R1008 VDD2.n17 VDD2.n11 289.615
R1009 VDD2.n6 VDD2.n0 289.615
R1010 VDD2.n18 VDD2.n17 185
R1011 VDD2.n16 VDD2.n15 185
R1012 VDD2.n5 VDD2.n4 185
R1013 VDD2.n7 VDD2.n6 185
R1014 VDD2.n14 VDD2.t0 151.613
R1015 VDD2.n3 VDD2.t1 151.613
R1016 VDD2.n17 VDD2.n16 104.615
R1017 VDD2.n6 VDD2.n5 104.615
R1018 VDD2.n22 VDD2.n10 85.2947
R1019 VDD2.n16 VDD2.t0 52.3082
R1020 VDD2.n5 VDD2.t1 52.3082
R1021 VDD2.n22 VDD2.n21 52.1611
R1022 VDD2.n15 VDD2.n14 15.3979
R1023 VDD2.n4 VDD2.n3 15.3979
R1024 VDD2.n18 VDD2.n13 12.8005
R1025 VDD2.n7 VDD2.n2 12.8005
R1026 VDD2.n19 VDD2.n11 12.0247
R1027 VDD2.n8 VDD2.n0 12.0247
R1028 VDD2.n21 VDD2.n20 9.45567
R1029 VDD2.n10 VDD2.n9 9.45567
R1030 VDD2.n20 VDD2.n19 9.3005
R1031 VDD2.n13 VDD2.n12 9.3005
R1032 VDD2.n9 VDD2.n8 9.3005
R1033 VDD2.n2 VDD2.n1 9.3005
R1034 VDD2.n14 VDD2.n12 4.69785
R1035 VDD2.n3 VDD2.n1 4.69785
R1036 VDD2.n21 VDD2.n11 1.93989
R1037 VDD2.n10 VDD2.n0 1.93989
R1038 VDD2.n19 VDD2.n18 1.16414
R1039 VDD2.n8 VDD2.n7 1.16414
R1040 VDD2 VDD2.n22 0.966017
R1041 VDD2.n15 VDD2.n13 0.388379
R1042 VDD2.n4 VDD2.n2 0.388379
R1043 VDD2.n20 VDD2.n12 0.155672
R1044 VDD2.n9 VDD2.n1 0.155672
R1045 VP.n0 VP.t1 91.9076
R1046 VP.n0 VP.t0 51.0008
R1047 VP VP.n0 0.621237
R1048 VDD1.n6 VDD1.n0 289.615
R1049 VDD1.n17 VDD1.n11 289.615
R1050 VDD1.n7 VDD1.n6 185
R1051 VDD1.n5 VDD1.n4 185
R1052 VDD1.n16 VDD1.n15 185
R1053 VDD1.n18 VDD1.n17 185
R1054 VDD1.n3 VDD1.t0 151.613
R1055 VDD1.n14 VDD1.t1 151.613
R1056 VDD1.n6 VDD1.n5 104.615
R1057 VDD1.n17 VDD1.n16 104.615
R1058 VDD1 VDD1.n21 86.7268
R1059 VDD1 VDD1.n10 53.1266
R1060 VDD1.n5 VDD1.t0 52.3082
R1061 VDD1.n16 VDD1.t1 52.3082
R1062 VDD1.n4 VDD1.n3 15.3979
R1063 VDD1.n15 VDD1.n14 15.3979
R1064 VDD1.n7 VDD1.n2 12.8005
R1065 VDD1.n18 VDD1.n13 12.8005
R1066 VDD1.n8 VDD1.n0 12.0247
R1067 VDD1.n19 VDD1.n11 12.0247
R1068 VDD1.n10 VDD1.n9 9.45567
R1069 VDD1.n21 VDD1.n20 9.45567
R1070 VDD1.n9 VDD1.n8 9.3005
R1071 VDD1.n2 VDD1.n1 9.3005
R1072 VDD1.n20 VDD1.n19 9.3005
R1073 VDD1.n13 VDD1.n12 9.3005
R1074 VDD1.n3 VDD1.n1 4.69785
R1075 VDD1.n14 VDD1.n12 4.69785
R1076 VDD1.n10 VDD1.n0 1.93989
R1077 VDD1.n21 VDD1.n11 1.93989
R1078 VDD1.n8 VDD1.n7 1.16414
R1079 VDD1.n19 VDD1.n18 1.16414
R1080 VDD1.n4 VDD1.n2 0.388379
R1081 VDD1.n15 VDD1.n13 0.388379
R1082 VDD1.n9 VDD1.n1 0.155672
R1083 VDD1.n20 VDD1.n12 0.155672
C0 VTAIL VN 1.22886f
C1 VP VDD2 0.39242f
C2 VDD1 VN 0.154274f
C3 VTAIL VP 1.24313f
C4 VP VDD1 1.07043f
C5 VP VN 4.31777f
C6 VTAIL VDD2 3.052f
C7 VDD1 VDD2 0.817405f
C8 VN VDD2 0.833792f
C9 VTAIL VDD1 2.99037f
C10 VDD2 B 3.168209f
C11 VDD1 B 5.02831f
C12 VTAIL B 3.665312f
C13 VN B 9.196779f
C14 VP B 7.124809f
C15 VDD1.n0 B 0.023792f
C16 VDD1.n1 B 0.133189f
C17 VDD1.n2 B 0.009229f
C18 VDD1.t0 B 0.038204f
C19 VDD1.n3 B 0.061889f
C20 VDD1.n4 B 0.012348f
C21 VDD1.n5 B 0.01636f
C22 VDD1.n6 B 0.046607f
C23 VDD1.n7 B 0.009772f
C24 VDD1.n8 B 0.009229f
C25 VDD1.n9 B 0.043686f
C26 VDD1.n10 B 0.039577f
C27 VDD1.n11 B 0.023792f
C28 VDD1.n12 B 0.133189f
C29 VDD1.n13 B 0.009229f
C30 VDD1.t1 B 0.038204f
C31 VDD1.n14 B 0.061889f
C32 VDD1.n15 B 0.012348f
C33 VDD1.n16 B 0.01636f
C34 VDD1.n17 B 0.046607f
C35 VDD1.n18 B 0.009772f
C36 VDD1.n19 B 0.009229f
C37 VDD1.n20 B 0.043686f
C38 VDD1.n21 B 0.368257f
C39 VP.t1 B 1.43089f
C40 VP.t0 B 0.862285f
C41 VP.n0 B 1.90547f
C42 VDD2.n0 B 0.025117f
C43 VDD2.n1 B 0.140602f
C44 VDD2.n2 B 0.009742f
C45 VDD2.t1 B 0.04033f
C46 VDD2.n3 B 0.065333f
C47 VDD2.n4 B 0.013035f
C48 VDD2.n5 B 0.01727f
C49 VDD2.n6 B 0.049201f
C50 VDD2.n7 B 0.010315f
C51 VDD2.n8 B 0.009742f
C52 VDD2.n9 B 0.046117f
C53 VDD2.n10 B 0.353788f
C54 VDD2.n11 B 0.025117f
C55 VDD2.n12 B 0.140602f
C56 VDD2.n13 B 0.009742f
C57 VDD2.t0 B 0.04033f
C58 VDD2.n14 B 0.065333f
C59 VDD2.n15 B 0.013035f
C60 VDD2.n16 B 0.01727f
C61 VDD2.n17 B 0.049201f
C62 VDD2.n18 B 0.010315f
C63 VDD2.n19 B 0.009742f
C64 VDD2.n20 B 0.046117f
C65 VDD2.n21 B 0.040076f
C66 VDD2.n22 B 1.6896f
C67 VTAIL.n0 B 0.029476f
C68 VTAIL.n1 B 0.165006f
C69 VTAIL.n2 B 0.011433f
C70 VTAIL.t1 B 0.04733f
C71 VTAIL.n3 B 0.076673f
C72 VTAIL.n4 B 0.015298f
C73 VTAIL.n5 B 0.020268f
C74 VTAIL.n6 B 0.057741f
C75 VTAIL.n7 B 0.012106f
C76 VTAIL.n8 B 0.011433f
C77 VTAIL.n9 B 0.054122f
C78 VTAIL.n10 B 0.032376f
C79 VTAIL.n11 B 1.05793f
C80 VTAIL.n12 B 0.029476f
C81 VTAIL.n13 B 0.165006f
C82 VTAIL.n14 B 0.011433f
C83 VTAIL.t3 B 0.04733f
C84 VTAIL.n15 B 0.076673f
C85 VTAIL.n16 B 0.015298f
C86 VTAIL.n17 B 0.020268f
C87 VTAIL.n18 B 0.057741f
C88 VTAIL.n19 B 0.012106f
C89 VTAIL.n20 B 0.011433f
C90 VTAIL.n21 B 0.054122f
C91 VTAIL.n22 B 0.032376f
C92 VTAIL.n23 B 1.11615f
C93 VTAIL.n24 B 0.029476f
C94 VTAIL.n25 B 0.165006f
C95 VTAIL.n26 B 0.011433f
C96 VTAIL.t0 B 0.04733f
C97 VTAIL.n27 B 0.076673f
C98 VTAIL.n28 B 0.015298f
C99 VTAIL.n29 B 0.020268f
C100 VTAIL.n30 B 0.057741f
C101 VTAIL.n31 B 0.012106f
C102 VTAIL.n32 B 0.011433f
C103 VTAIL.n33 B 0.054122f
C104 VTAIL.n34 B 0.032376f
C105 VTAIL.n35 B 0.867327f
C106 VTAIL.n36 B 0.029476f
C107 VTAIL.n37 B 0.165006f
C108 VTAIL.n38 B 0.011433f
C109 VTAIL.t2 B 0.04733f
C110 VTAIL.n39 B 0.076673f
C111 VTAIL.n40 B 0.015298f
C112 VTAIL.n41 B 0.020268f
C113 VTAIL.n42 B 0.057741f
C114 VTAIL.n43 B 0.012106f
C115 VTAIL.n44 B 0.011433f
C116 VTAIL.n45 B 0.054122f
C117 VTAIL.n46 B 0.032376f
C118 VTAIL.n47 B 0.768921f
C119 VN.t0 B 0.859701f
C120 VN.t1 B 1.41928f
.ends

