* NGSPICE file created from diff_pair_sample_0636.ext - technology: sky130A

.subckt diff_pair_sample_0636 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=3.93
X1 VTAIL.t8 VN.t0 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=3.93
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=3.93
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=3.93
X4 VTAIL.t10 VP.t0 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=3.93
X5 VTAIL.t7 VN.t1 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=3.93
X6 VDD2.t2 VN.t2 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=3.93
X7 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=3.93
X8 VDD1.t3 VP.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=3.93
X9 VDD2.t3 VN.t3 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=3.93
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=0 ps=0 w=9.39 l=3.93
X11 VDD2.t4 VN.t4 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=3.93
X12 VDD2.t5 VN.t5 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=3.93
X13 VDD1.t2 VP.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6621 pd=19.56 as=1.54935 ps=9.72 w=9.39 l=3.93
X14 VTAIL.t9 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=1.54935 ps=9.72 w=9.39 l=3.93
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.54935 pd=9.72 as=3.6621 ps=19.56 w=9.39 l=3.93
R0 B.n710 B.n709 585
R1 B.n710 B.n106 585
R2 B.n713 B.n712 585
R3 B.n714 B.n149 585
R4 B.n716 B.n715 585
R5 B.n718 B.n148 585
R6 B.n721 B.n720 585
R7 B.n722 B.n147 585
R8 B.n724 B.n723 585
R9 B.n726 B.n146 585
R10 B.n729 B.n728 585
R11 B.n730 B.n145 585
R12 B.n732 B.n731 585
R13 B.n734 B.n144 585
R14 B.n737 B.n736 585
R15 B.n738 B.n143 585
R16 B.n740 B.n739 585
R17 B.n742 B.n142 585
R18 B.n745 B.n744 585
R19 B.n746 B.n141 585
R20 B.n748 B.n747 585
R21 B.n750 B.n140 585
R22 B.n753 B.n752 585
R23 B.n754 B.n139 585
R24 B.n756 B.n755 585
R25 B.n758 B.n138 585
R26 B.n761 B.n760 585
R27 B.n762 B.n137 585
R28 B.n764 B.n763 585
R29 B.n766 B.n136 585
R30 B.n769 B.n768 585
R31 B.n770 B.n135 585
R32 B.n772 B.n771 585
R33 B.n774 B.n134 585
R34 B.n777 B.n776 585
R35 B.n779 B.n131 585
R36 B.n781 B.n780 585
R37 B.n783 B.n130 585
R38 B.n786 B.n785 585
R39 B.n787 B.n129 585
R40 B.n789 B.n788 585
R41 B.n791 B.n128 585
R42 B.n793 B.n792 585
R43 B.n795 B.n794 585
R44 B.n798 B.n797 585
R45 B.n799 B.n123 585
R46 B.n801 B.n800 585
R47 B.n803 B.n122 585
R48 B.n806 B.n805 585
R49 B.n807 B.n121 585
R50 B.n809 B.n808 585
R51 B.n811 B.n120 585
R52 B.n814 B.n813 585
R53 B.n815 B.n119 585
R54 B.n817 B.n816 585
R55 B.n819 B.n118 585
R56 B.n822 B.n821 585
R57 B.n823 B.n117 585
R58 B.n825 B.n824 585
R59 B.n827 B.n116 585
R60 B.n830 B.n829 585
R61 B.n831 B.n115 585
R62 B.n833 B.n832 585
R63 B.n835 B.n114 585
R64 B.n838 B.n837 585
R65 B.n839 B.n113 585
R66 B.n841 B.n840 585
R67 B.n843 B.n112 585
R68 B.n846 B.n845 585
R69 B.n847 B.n111 585
R70 B.n849 B.n848 585
R71 B.n851 B.n110 585
R72 B.n854 B.n853 585
R73 B.n855 B.n109 585
R74 B.n857 B.n856 585
R75 B.n859 B.n108 585
R76 B.n862 B.n861 585
R77 B.n863 B.n107 585
R78 B.n708 B.n105 585
R79 B.n866 B.n105 585
R80 B.n707 B.n104 585
R81 B.n867 B.n104 585
R82 B.n706 B.n103 585
R83 B.n868 B.n103 585
R84 B.n705 B.n704 585
R85 B.n704 B.n99 585
R86 B.n703 B.n98 585
R87 B.n874 B.n98 585
R88 B.n702 B.n97 585
R89 B.n875 B.n97 585
R90 B.n701 B.n96 585
R91 B.n876 B.n96 585
R92 B.n700 B.n699 585
R93 B.n699 B.n92 585
R94 B.n698 B.n91 585
R95 B.n882 B.n91 585
R96 B.n697 B.n90 585
R97 B.n883 B.n90 585
R98 B.n696 B.n89 585
R99 B.n884 B.n89 585
R100 B.n695 B.n694 585
R101 B.n694 B.n85 585
R102 B.n693 B.n84 585
R103 B.n890 B.n84 585
R104 B.n692 B.n83 585
R105 B.n891 B.n83 585
R106 B.n691 B.n82 585
R107 B.n892 B.n82 585
R108 B.n690 B.n689 585
R109 B.n689 B.n78 585
R110 B.n688 B.n77 585
R111 B.n898 B.n77 585
R112 B.n687 B.n76 585
R113 B.n899 B.n76 585
R114 B.n686 B.n75 585
R115 B.n900 B.n75 585
R116 B.n685 B.n684 585
R117 B.n684 B.n71 585
R118 B.n683 B.n70 585
R119 B.n906 B.n70 585
R120 B.n682 B.n69 585
R121 B.n907 B.n69 585
R122 B.n681 B.n68 585
R123 B.n908 B.n68 585
R124 B.n680 B.n679 585
R125 B.n679 B.n64 585
R126 B.n678 B.n63 585
R127 B.n914 B.n63 585
R128 B.n677 B.n62 585
R129 B.n915 B.n62 585
R130 B.n676 B.n61 585
R131 B.n916 B.n61 585
R132 B.n675 B.n674 585
R133 B.n674 B.n57 585
R134 B.n673 B.n56 585
R135 B.n922 B.n56 585
R136 B.n672 B.n55 585
R137 B.n923 B.n55 585
R138 B.n671 B.n54 585
R139 B.n924 B.n54 585
R140 B.n670 B.n669 585
R141 B.n669 B.n50 585
R142 B.n668 B.n49 585
R143 B.n930 B.n49 585
R144 B.n667 B.n48 585
R145 B.n931 B.n48 585
R146 B.n666 B.n47 585
R147 B.n932 B.n47 585
R148 B.n665 B.n664 585
R149 B.n664 B.n43 585
R150 B.n663 B.n42 585
R151 B.n938 B.n42 585
R152 B.n662 B.n41 585
R153 B.n939 B.n41 585
R154 B.n661 B.n40 585
R155 B.n940 B.n40 585
R156 B.n660 B.n659 585
R157 B.n659 B.n36 585
R158 B.n658 B.n35 585
R159 B.n946 B.n35 585
R160 B.n657 B.n34 585
R161 B.n947 B.n34 585
R162 B.n656 B.n33 585
R163 B.n948 B.n33 585
R164 B.n655 B.n654 585
R165 B.n654 B.n29 585
R166 B.n653 B.n28 585
R167 B.n954 B.n28 585
R168 B.n652 B.n27 585
R169 B.n955 B.n27 585
R170 B.n651 B.n26 585
R171 B.n956 B.n26 585
R172 B.n650 B.n649 585
R173 B.n649 B.n22 585
R174 B.n648 B.n21 585
R175 B.n962 B.n21 585
R176 B.n647 B.n20 585
R177 B.n963 B.n20 585
R178 B.n646 B.n19 585
R179 B.n964 B.n19 585
R180 B.n645 B.n644 585
R181 B.n644 B.n15 585
R182 B.n643 B.n14 585
R183 B.n970 B.n14 585
R184 B.n642 B.n13 585
R185 B.n971 B.n13 585
R186 B.n641 B.n12 585
R187 B.n972 B.n12 585
R188 B.n640 B.n639 585
R189 B.n639 B.n8 585
R190 B.n638 B.n7 585
R191 B.n978 B.n7 585
R192 B.n637 B.n6 585
R193 B.n979 B.n6 585
R194 B.n636 B.n5 585
R195 B.n980 B.n5 585
R196 B.n635 B.n634 585
R197 B.n634 B.n4 585
R198 B.n633 B.n150 585
R199 B.n633 B.n632 585
R200 B.n623 B.n151 585
R201 B.n152 B.n151 585
R202 B.n625 B.n624 585
R203 B.n626 B.n625 585
R204 B.n622 B.n157 585
R205 B.n157 B.n156 585
R206 B.n621 B.n620 585
R207 B.n620 B.n619 585
R208 B.n159 B.n158 585
R209 B.n160 B.n159 585
R210 B.n612 B.n611 585
R211 B.n613 B.n612 585
R212 B.n610 B.n165 585
R213 B.n165 B.n164 585
R214 B.n609 B.n608 585
R215 B.n608 B.n607 585
R216 B.n167 B.n166 585
R217 B.n168 B.n167 585
R218 B.n600 B.n599 585
R219 B.n601 B.n600 585
R220 B.n598 B.n173 585
R221 B.n173 B.n172 585
R222 B.n597 B.n596 585
R223 B.n596 B.n595 585
R224 B.n175 B.n174 585
R225 B.n176 B.n175 585
R226 B.n588 B.n587 585
R227 B.n589 B.n588 585
R228 B.n586 B.n181 585
R229 B.n181 B.n180 585
R230 B.n585 B.n584 585
R231 B.n584 B.n583 585
R232 B.n183 B.n182 585
R233 B.n184 B.n183 585
R234 B.n576 B.n575 585
R235 B.n577 B.n576 585
R236 B.n574 B.n188 585
R237 B.n192 B.n188 585
R238 B.n573 B.n572 585
R239 B.n572 B.n571 585
R240 B.n190 B.n189 585
R241 B.n191 B.n190 585
R242 B.n564 B.n563 585
R243 B.n565 B.n564 585
R244 B.n562 B.n197 585
R245 B.n197 B.n196 585
R246 B.n561 B.n560 585
R247 B.n560 B.n559 585
R248 B.n199 B.n198 585
R249 B.n200 B.n199 585
R250 B.n552 B.n551 585
R251 B.n553 B.n552 585
R252 B.n550 B.n205 585
R253 B.n205 B.n204 585
R254 B.n549 B.n548 585
R255 B.n548 B.n547 585
R256 B.n207 B.n206 585
R257 B.n208 B.n207 585
R258 B.n540 B.n539 585
R259 B.n541 B.n540 585
R260 B.n538 B.n212 585
R261 B.n216 B.n212 585
R262 B.n537 B.n536 585
R263 B.n536 B.n535 585
R264 B.n214 B.n213 585
R265 B.n215 B.n214 585
R266 B.n528 B.n527 585
R267 B.n529 B.n528 585
R268 B.n526 B.n221 585
R269 B.n221 B.n220 585
R270 B.n525 B.n524 585
R271 B.n524 B.n523 585
R272 B.n223 B.n222 585
R273 B.n224 B.n223 585
R274 B.n516 B.n515 585
R275 B.n517 B.n516 585
R276 B.n514 B.n229 585
R277 B.n229 B.n228 585
R278 B.n513 B.n512 585
R279 B.n512 B.n511 585
R280 B.n231 B.n230 585
R281 B.n232 B.n231 585
R282 B.n504 B.n503 585
R283 B.n505 B.n504 585
R284 B.n502 B.n237 585
R285 B.n237 B.n236 585
R286 B.n501 B.n500 585
R287 B.n500 B.n499 585
R288 B.n239 B.n238 585
R289 B.n240 B.n239 585
R290 B.n492 B.n491 585
R291 B.n493 B.n492 585
R292 B.n490 B.n244 585
R293 B.n248 B.n244 585
R294 B.n489 B.n488 585
R295 B.n488 B.n487 585
R296 B.n246 B.n245 585
R297 B.n247 B.n246 585
R298 B.n480 B.n479 585
R299 B.n481 B.n480 585
R300 B.n478 B.n253 585
R301 B.n253 B.n252 585
R302 B.n477 B.n476 585
R303 B.n476 B.n475 585
R304 B.n255 B.n254 585
R305 B.n256 B.n255 585
R306 B.n468 B.n467 585
R307 B.n469 B.n468 585
R308 B.n466 B.n261 585
R309 B.n261 B.n260 585
R310 B.n465 B.n464 585
R311 B.n464 B.n463 585
R312 B.n460 B.n265 585
R313 B.n459 B.n458 585
R314 B.n456 B.n266 585
R315 B.n456 B.n264 585
R316 B.n455 B.n454 585
R317 B.n453 B.n452 585
R318 B.n451 B.n268 585
R319 B.n449 B.n448 585
R320 B.n447 B.n269 585
R321 B.n446 B.n445 585
R322 B.n443 B.n270 585
R323 B.n441 B.n440 585
R324 B.n439 B.n271 585
R325 B.n438 B.n437 585
R326 B.n435 B.n272 585
R327 B.n433 B.n432 585
R328 B.n431 B.n273 585
R329 B.n430 B.n429 585
R330 B.n427 B.n274 585
R331 B.n425 B.n424 585
R332 B.n423 B.n275 585
R333 B.n422 B.n421 585
R334 B.n419 B.n276 585
R335 B.n417 B.n416 585
R336 B.n415 B.n277 585
R337 B.n414 B.n413 585
R338 B.n411 B.n278 585
R339 B.n409 B.n408 585
R340 B.n407 B.n279 585
R341 B.n406 B.n405 585
R342 B.n403 B.n280 585
R343 B.n401 B.n400 585
R344 B.n399 B.n281 585
R345 B.n398 B.n397 585
R346 B.n395 B.n282 585
R347 B.n393 B.n392 585
R348 B.n391 B.n283 585
R349 B.n390 B.n389 585
R350 B.n387 B.n287 585
R351 B.n385 B.n384 585
R352 B.n383 B.n288 585
R353 B.n382 B.n381 585
R354 B.n379 B.n289 585
R355 B.n377 B.n376 585
R356 B.n374 B.n290 585
R357 B.n373 B.n372 585
R358 B.n370 B.n293 585
R359 B.n368 B.n367 585
R360 B.n366 B.n294 585
R361 B.n365 B.n364 585
R362 B.n362 B.n295 585
R363 B.n360 B.n359 585
R364 B.n358 B.n296 585
R365 B.n357 B.n356 585
R366 B.n354 B.n297 585
R367 B.n352 B.n351 585
R368 B.n350 B.n298 585
R369 B.n349 B.n348 585
R370 B.n346 B.n299 585
R371 B.n344 B.n343 585
R372 B.n342 B.n300 585
R373 B.n341 B.n340 585
R374 B.n338 B.n301 585
R375 B.n336 B.n335 585
R376 B.n334 B.n302 585
R377 B.n333 B.n332 585
R378 B.n330 B.n303 585
R379 B.n328 B.n327 585
R380 B.n326 B.n304 585
R381 B.n325 B.n324 585
R382 B.n322 B.n305 585
R383 B.n320 B.n319 585
R384 B.n318 B.n306 585
R385 B.n317 B.n316 585
R386 B.n314 B.n307 585
R387 B.n312 B.n311 585
R388 B.n310 B.n309 585
R389 B.n263 B.n262 585
R390 B.n462 B.n461 585
R391 B.n463 B.n462 585
R392 B.n259 B.n258 585
R393 B.n260 B.n259 585
R394 B.n471 B.n470 585
R395 B.n470 B.n469 585
R396 B.n472 B.n257 585
R397 B.n257 B.n256 585
R398 B.n474 B.n473 585
R399 B.n475 B.n474 585
R400 B.n251 B.n250 585
R401 B.n252 B.n251 585
R402 B.n483 B.n482 585
R403 B.n482 B.n481 585
R404 B.n484 B.n249 585
R405 B.n249 B.n247 585
R406 B.n486 B.n485 585
R407 B.n487 B.n486 585
R408 B.n243 B.n242 585
R409 B.n248 B.n243 585
R410 B.n495 B.n494 585
R411 B.n494 B.n493 585
R412 B.n496 B.n241 585
R413 B.n241 B.n240 585
R414 B.n498 B.n497 585
R415 B.n499 B.n498 585
R416 B.n235 B.n234 585
R417 B.n236 B.n235 585
R418 B.n507 B.n506 585
R419 B.n506 B.n505 585
R420 B.n508 B.n233 585
R421 B.n233 B.n232 585
R422 B.n510 B.n509 585
R423 B.n511 B.n510 585
R424 B.n227 B.n226 585
R425 B.n228 B.n227 585
R426 B.n519 B.n518 585
R427 B.n518 B.n517 585
R428 B.n520 B.n225 585
R429 B.n225 B.n224 585
R430 B.n522 B.n521 585
R431 B.n523 B.n522 585
R432 B.n219 B.n218 585
R433 B.n220 B.n219 585
R434 B.n531 B.n530 585
R435 B.n530 B.n529 585
R436 B.n532 B.n217 585
R437 B.n217 B.n215 585
R438 B.n534 B.n533 585
R439 B.n535 B.n534 585
R440 B.n211 B.n210 585
R441 B.n216 B.n211 585
R442 B.n543 B.n542 585
R443 B.n542 B.n541 585
R444 B.n544 B.n209 585
R445 B.n209 B.n208 585
R446 B.n546 B.n545 585
R447 B.n547 B.n546 585
R448 B.n203 B.n202 585
R449 B.n204 B.n203 585
R450 B.n555 B.n554 585
R451 B.n554 B.n553 585
R452 B.n556 B.n201 585
R453 B.n201 B.n200 585
R454 B.n558 B.n557 585
R455 B.n559 B.n558 585
R456 B.n195 B.n194 585
R457 B.n196 B.n195 585
R458 B.n567 B.n566 585
R459 B.n566 B.n565 585
R460 B.n568 B.n193 585
R461 B.n193 B.n191 585
R462 B.n570 B.n569 585
R463 B.n571 B.n570 585
R464 B.n187 B.n186 585
R465 B.n192 B.n187 585
R466 B.n579 B.n578 585
R467 B.n578 B.n577 585
R468 B.n580 B.n185 585
R469 B.n185 B.n184 585
R470 B.n582 B.n581 585
R471 B.n583 B.n582 585
R472 B.n179 B.n178 585
R473 B.n180 B.n179 585
R474 B.n591 B.n590 585
R475 B.n590 B.n589 585
R476 B.n592 B.n177 585
R477 B.n177 B.n176 585
R478 B.n594 B.n593 585
R479 B.n595 B.n594 585
R480 B.n171 B.n170 585
R481 B.n172 B.n171 585
R482 B.n603 B.n602 585
R483 B.n602 B.n601 585
R484 B.n604 B.n169 585
R485 B.n169 B.n168 585
R486 B.n606 B.n605 585
R487 B.n607 B.n606 585
R488 B.n163 B.n162 585
R489 B.n164 B.n163 585
R490 B.n615 B.n614 585
R491 B.n614 B.n613 585
R492 B.n616 B.n161 585
R493 B.n161 B.n160 585
R494 B.n618 B.n617 585
R495 B.n619 B.n618 585
R496 B.n155 B.n154 585
R497 B.n156 B.n155 585
R498 B.n628 B.n627 585
R499 B.n627 B.n626 585
R500 B.n629 B.n153 585
R501 B.n153 B.n152 585
R502 B.n631 B.n630 585
R503 B.n632 B.n631 585
R504 B.n2 B.n0 585
R505 B.n4 B.n2 585
R506 B.n3 B.n1 585
R507 B.n979 B.n3 585
R508 B.n977 B.n976 585
R509 B.n978 B.n977 585
R510 B.n975 B.n9 585
R511 B.n9 B.n8 585
R512 B.n974 B.n973 585
R513 B.n973 B.n972 585
R514 B.n11 B.n10 585
R515 B.n971 B.n11 585
R516 B.n969 B.n968 585
R517 B.n970 B.n969 585
R518 B.n967 B.n16 585
R519 B.n16 B.n15 585
R520 B.n966 B.n965 585
R521 B.n965 B.n964 585
R522 B.n18 B.n17 585
R523 B.n963 B.n18 585
R524 B.n961 B.n960 585
R525 B.n962 B.n961 585
R526 B.n959 B.n23 585
R527 B.n23 B.n22 585
R528 B.n958 B.n957 585
R529 B.n957 B.n956 585
R530 B.n25 B.n24 585
R531 B.n955 B.n25 585
R532 B.n953 B.n952 585
R533 B.n954 B.n953 585
R534 B.n951 B.n30 585
R535 B.n30 B.n29 585
R536 B.n950 B.n949 585
R537 B.n949 B.n948 585
R538 B.n32 B.n31 585
R539 B.n947 B.n32 585
R540 B.n945 B.n944 585
R541 B.n946 B.n945 585
R542 B.n943 B.n37 585
R543 B.n37 B.n36 585
R544 B.n942 B.n941 585
R545 B.n941 B.n940 585
R546 B.n39 B.n38 585
R547 B.n939 B.n39 585
R548 B.n937 B.n936 585
R549 B.n938 B.n937 585
R550 B.n935 B.n44 585
R551 B.n44 B.n43 585
R552 B.n934 B.n933 585
R553 B.n933 B.n932 585
R554 B.n46 B.n45 585
R555 B.n931 B.n46 585
R556 B.n929 B.n928 585
R557 B.n930 B.n929 585
R558 B.n927 B.n51 585
R559 B.n51 B.n50 585
R560 B.n926 B.n925 585
R561 B.n925 B.n924 585
R562 B.n53 B.n52 585
R563 B.n923 B.n53 585
R564 B.n921 B.n920 585
R565 B.n922 B.n921 585
R566 B.n919 B.n58 585
R567 B.n58 B.n57 585
R568 B.n918 B.n917 585
R569 B.n917 B.n916 585
R570 B.n60 B.n59 585
R571 B.n915 B.n60 585
R572 B.n913 B.n912 585
R573 B.n914 B.n913 585
R574 B.n911 B.n65 585
R575 B.n65 B.n64 585
R576 B.n910 B.n909 585
R577 B.n909 B.n908 585
R578 B.n67 B.n66 585
R579 B.n907 B.n67 585
R580 B.n905 B.n904 585
R581 B.n906 B.n905 585
R582 B.n903 B.n72 585
R583 B.n72 B.n71 585
R584 B.n902 B.n901 585
R585 B.n901 B.n900 585
R586 B.n74 B.n73 585
R587 B.n899 B.n74 585
R588 B.n897 B.n896 585
R589 B.n898 B.n897 585
R590 B.n895 B.n79 585
R591 B.n79 B.n78 585
R592 B.n894 B.n893 585
R593 B.n893 B.n892 585
R594 B.n81 B.n80 585
R595 B.n891 B.n81 585
R596 B.n889 B.n888 585
R597 B.n890 B.n889 585
R598 B.n887 B.n86 585
R599 B.n86 B.n85 585
R600 B.n886 B.n885 585
R601 B.n885 B.n884 585
R602 B.n88 B.n87 585
R603 B.n883 B.n88 585
R604 B.n881 B.n880 585
R605 B.n882 B.n881 585
R606 B.n879 B.n93 585
R607 B.n93 B.n92 585
R608 B.n878 B.n877 585
R609 B.n877 B.n876 585
R610 B.n95 B.n94 585
R611 B.n875 B.n95 585
R612 B.n873 B.n872 585
R613 B.n874 B.n873 585
R614 B.n871 B.n100 585
R615 B.n100 B.n99 585
R616 B.n870 B.n869 585
R617 B.n869 B.n868 585
R618 B.n102 B.n101 585
R619 B.n867 B.n102 585
R620 B.n865 B.n864 585
R621 B.n866 B.n865 585
R622 B.n982 B.n981 585
R623 B.n981 B.n980 585
R624 B.n462 B.n265 574.183
R625 B.n865 B.n107 574.183
R626 B.n464 B.n263 574.183
R627 B.n710 B.n105 574.183
R628 B.n291 B.t19 319.911
R629 B.n132 B.t15 319.911
R630 B.n284 B.t9 319.911
R631 B.n124 B.t12 319.911
R632 B.n291 B.t17 267.024
R633 B.n284 B.t6 267.024
R634 B.n124 B.t10 267.024
R635 B.n132 B.t14 267.024
R636 B.n711 B.n106 256.663
R637 B.n717 B.n106 256.663
R638 B.n719 B.n106 256.663
R639 B.n725 B.n106 256.663
R640 B.n727 B.n106 256.663
R641 B.n733 B.n106 256.663
R642 B.n735 B.n106 256.663
R643 B.n741 B.n106 256.663
R644 B.n743 B.n106 256.663
R645 B.n749 B.n106 256.663
R646 B.n751 B.n106 256.663
R647 B.n757 B.n106 256.663
R648 B.n759 B.n106 256.663
R649 B.n765 B.n106 256.663
R650 B.n767 B.n106 256.663
R651 B.n773 B.n106 256.663
R652 B.n775 B.n106 256.663
R653 B.n782 B.n106 256.663
R654 B.n784 B.n106 256.663
R655 B.n790 B.n106 256.663
R656 B.n127 B.n106 256.663
R657 B.n796 B.n106 256.663
R658 B.n802 B.n106 256.663
R659 B.n804 B.n106 256.663
R660 B.n810 B.n106 256.663
R661 B.n812 B.n106 256.663
R662 B.n818 B.n106 256.663
R663 B.n820 B.n106 256.663
R664 B.n826 B.n106 256.663
R665 B.n828 B.n106 256.663
R666 B.n834 B.n106 256.663
R667 B.n836 B.n106 256.663
R668 B.n842 B.n106 256.663
R669 B.n844 B.n106 256.663
R670 B.n850 B.n106 256.663
R671 B.n852 B.n106 256.663
R672 B.n858 B.n106 256.663
R673 B.n860 B.n106 256.663
R674 B.n457 B.n264 256.663
R675 B.n267 B.n264 256.663
R676 B.n450 B.n264 256.663
R677 B.n444 B.n264 256.663
R678 B.n442 B.n264 256.663
R679 B.n436 B.n264 256.663
R680 B.n434 B.n264 256.663
R681 B.n428 B.n264 256.663
R682 B.n426 B.n264 256.663
R683 B.n420 B.n264 256.663
R684 B.n418 B.n264 256.663
R685 B.n412 B.n264 256.663
R686 B.n410 B.n264 256.663
R687 B.n404 B.n264 256.663
R688 B.n402 B.n264 256.663
R689 B.n396 B.n264 256.663
R690 B.n394 B.n264 256.663
R691 B.n388 B.n264 256.663
R692 B.n386 B.n264 256.663
R693 B.n380 B.n264 256.663
R694 B.n378 B.n264 256.663
R695 B.n371 B.n264 256.663
R696 B.n369 B.n264 256.663
R697 B.n363 B.n264 256.663
R698 B.n361 B.n264 256.663
R699 B.n355 B.n264 256.663
R700 B.n353 B.n264 256.663
R701 B.n347 B.n264 256.663
R702 B.n345 B.n264 256.663
R703 B.n339 B.n264 256.663
R704 B.n337 B.n264 256.663
R705 B.n331 B.n264 256.663
R706 B.n329 B.n264 256.663
R707 B.n323 B.n264 256.663
R708 B.n321 B.n264 256.663
R709 B.n315 B.n264 256.663
R710 B.n313 B.n264 256.663
R711 B.n308 B.n264 256.663
R712 B.n292 B.t18 237.293
R713 B.n133 B.t16 237.293
R714 B.n285 B.t8 237.292
R715 B.n125 B.t13 237.292
R716 B.n462 B.n259 163.367
R717 B.n470 B.n259 163.367
R718 B.n470 B.n257 163.367
R719 B.n474 B.n257 163.367
R720 B.n474 B.n251 163.367
R721 B.n482 B.n251 163.367
R722 B.n482 B.n249 163.367
R723 B.n486 B.n249 163.367
R724 B.n486 B.n243 163.367
R725 B.n494 B.n243 163.367
R726 B.n494 B.n241 163.367
R727 B.n498 B.n241 163.367
R728 B.n498 B.n235 163.367
R729 B.n506 B.n235 163.367
R730 B.n506 B.n233 163.367
R731 B.n510 B.n233 163.367
R732 B.n510 B.n227 163.367
R733 B.n518 B.n227 163.367
R734 B.n518 B.n225 163.367
R735 B.n522 B.n225 163.367
R736 B.n522 B.n219 163.367
R737 B.n530 B.n219 163.367
R738 B.n530 B.n217 163.367
R739 B.n534 B.n217 163.367
R740 B.n534 B.n211 163.367
R741 B.n542 B.n211 163.367
R742 B.n542 B.n209 163.367
R743 B.n546 B.n209 163.367
R744 B.n546 B.n203 163.367
R745 B.n554 B.n203 163.367
R746 B.n554 B.n201 163.367
R747 B.n558 B.n201 163.367
R748 B.n558 B.n195 163.367
R749 B.n566 B.n195 163.367
R750 B.n566 B.n193 163.367
R751 B.n570 B.n193 163.367
R752 B.n570 B.n187 163.367
R753 B.n578 B.n187 163.367
R754 B.n578 B.n185 163.367
R755 B.n582 B.n185 163.367
R756 B.n582 B.n179 163.367
R757 B.n590 B.n179 163.367
R758 B.n590 B.n177 163.367
R759 B.n594 B.n177 163.367
R760 B.n594 B.n171 163.367
R761 B.n602 B.n171 163.367
R762 B.n602 B.n169 163.367
R763 B.n606 B.n169 163.367
R764 B.n606 B.n163 163.367
R765 B.n614 B.n163 163.367
R766 B.n614 B.n161 163.367
R767 B.n618 B.n161 163.367
R768 B.n618 B.n155 163.367
R769 B.n627 B.n155 163.367
R770 B.n627 B.n153 163.367
R771 B.n631 B.n153 163.367
R772 B.n631 B.n2 163.367
R773 B.n981 B.n2 163.367
R774 B.n981 B.n3 163.367
R775 B.n977 B.n3 163.367
R776 B.n977 B.n9 163.367
R777 B.n973 B.n9 163.367
R778 B.n973 B.n11 163.367
R779 B.n969 B.n11 163.367
R780 B.n969 B.n16 163.367
R781 B.n965 B.n16 163.367
R782 B.n965 B.n18 163.367
R783 B.n961 B.n18 163.367
R784 B.n961 B.n23 163.367
R785 B.n957 B.n23 163.367
R786 B.n957 B.n25 163.367
R787 B.n953 B.n25 163.367
R788 B.n953 B.n30 163.367
R789 B.n949 B.n30 163.367
R790 B.n949 B.n32 163.367
R791 B.n945 B.n32 163.367
R792 B.n945 B.n37 163.367
R793 B.n941 B.n37 163.367
R794 B.n941 B.n39 163.367
R795 B.n937 B.n39 163.367
R796 B.n937 B.n44 163.367
R797 B.n933 B.n44 163.367
R798 B.n933 B.n46 163.367
R799 B.n929 B.n46 163.367
R800 B.n929 B.n51 163.367
R801 B.n925 B.n51 163.367
R802 B.n925 B.n53 163.367
R803 B.n921 B.n53 163.367
R804 B.n921 B.n58 163.367
R805 B.n917 B.n58 163.367
R806 B.n917 B.n60 163.367
R807 B.n913 B.n60 163.367
R808 B.n913 B.n65 163.367
R809 B.n909 B.n65 163.367
R810 B.n909 B.n67 163.367
R811 B.n905 B.n67 163.367
R812 B.n905 B.n72 163.367
R813 B.n901 B.n72 163.367
R814 B.n901 B.n74 163.367
R815 B.n897 B.n74 163.367
R816 B.n897 B.n79 163.367
R817 B.n893 B.n79 163.367
R818 B.n893 B.n81 163.367
R819 B.n889 B.n81 163.367
R820 B.n889 B.n86 163.367
R821 B.n885 B.n86 163.367
R822 B.n885 B.n88 163.367
R823 B.n881 B.n88 163.367
R824 B.n881 B.n93 163.367
R825 B.n877 B.n93 163.367
R826 B.n877 B.n95 163.367
R827 B.n873 B.n95 163.367
R828 B.n873 B.n100 163.367
R829 B.n869 B.n100 163.367
R830 B.n869 B.n102 163.367
R831 B.n865 B.n102 163.367
R832 B.n458 B.n456 163.367
R833 B.n456 B.n455 163.367
R834 B.n452 B.n451 163.367
R835 B.n449 B.n269 163.367
R836 B.n445 B.n443 163.367
R837 B.n441 B.n271 163.367
R838 B.n437 B.n435 163.367
R839 B.n433 B.n273 163.367
R840 B.n429 B.n427 163.367
R841 B.n425 B.n275 163.367
R842 B.n421 B.n419 163.367
R843 B.n417 B.n277 163.367
R844 B.n413 B.n411 163.367
R845 B.n409 B.n279 163.367
R846 B.n405 B.n403 163.367
R847 B.n401 B.n281 163.367
R848 B.n397 B.n395 163.367
R849 B.n393 B.n283 163.367
R850 B.n389 B.n387 163.367
R851 B.n385 B.n288 163.367
R852 B.n381 B.n379 163.367
R853 B.n377 B.n290 163.367
R854 B.n372 B.n370 163.367
R855 B.n368 B.n294 163.367
R856 B.n364 B.n362 163.367
R857 B.n360 B.n296 163.367
R858 B.n356 B.n354 163.367
R859 B.n352 B.n298 163.367
R860 B.n348 B.n346 163.367
R861 B.n344 B.n300 163.367
R862 B.n340 B.n338 163.367
R863 B.n336 B.n302 163.367
R864 B.n332 B.n330 163.367
R865 B.n328 B.n304 163.367
R866 B.n324 B.n322 163.367
R867 B.n320 B.n306 163.367
R868 B.n316 B.n314 163.367
R869 B.n312 B.n309 163.367
R870 B.n464 B.n261 163.367
R871 B.n468 B.n261 163.367
R872 B.n468 B.n255 163.367
R873 B.n476 B.n255 163.367
R874 B.n476 B.n253 163.367
R875 B.n480 B.n253 163.367
R876 B.n480 B.n246 163.367
R877 B.n488 B.n246 163.367
R878 B.n488 B.n244 163.367
R879 B.n492 B.n244 163.367
R880 B.n492 B.n239 163.367
R881 B.n500 B.n239 163.367
R882 B.n500 B.n237 163.367
R883 B.n504 B.n237 163.367
R884 B.n504 B.n231 163.367
R885 B.n512 B.n231 163.367
R886 B.n512 B.n229 163.367
R887 B.n516 B.n229 163.367
R888 B.n516 B.n223 163.367
R889 B.n524 B.n223 163.367
R890 B.n524 B.n221 163.367
R891 B.n528 B.n221 163.367
R892 B.n528 B.n214 163.367
R893 B.n536 B.n214 163.367
R894 B.n536 B.n212 163.367
R895 B.n540 B.n212 163.367
R896 B.n540 B.n207 163.367
R897 B.n548 B.n207 163.367
R898 B.n548 B.n205 163.367
R899 B.n552 B.n205 163.367
R900 B.n552 B.n199 163.367
R901 B.n560 B.n199 163.367
R902 B.n560 B.n197 163.367
R903 B.n564 B.n197 163.367
R904 B.n564 B.n190 163.367
R905 B.n572 B.n190 163.367
R906 B.n572 B.n188 163.367
R907 B.n576 B.n188 163.367
R908 B.n576 B.n183 163.367
R909 B.n584 B.n183 163.367
R910 B.n584 B.n181 163.367
R911 B.n588 B.n181 163.367
R912 B.n588 B.n175 163.367
R913 B.n596 B.n175 163.367
R914 B.n596 B.n173 163.367
R915 B.n600 B.n173 163.367
R916 B.n600 B.n167 163.367
R917 B.n608 B.n167 163.367
R918 B.n608 B.n165 163.367
R919 B.n612 B.n165 163.367
R920 B.n612 B.n159 163.367
R921 B.n620 B.n159 163.367
R922 B.n620 B.n157 163.367
R923 B.n625 B.n157 163.367
R924 B.n625 B.n151 163.367
R925 B.n633 B.n151 163.367
R926 B.n634 B.n633 163.367
R927 B.n634 B.n5 163.367
R928 B.n6 B.n5 163.367
R929 B.n7 B.n6 163.367
R930 B.n639 B.n7 163.367
R931 B.n639 B.n12 163.367
R932 B.n13 B.n12 163.367
R933 B.n14 B.n13 163.367
R934 B.n644 B.n14 163.367
R935 B.n644 B.n19 163.367
R936 B.n20 B.n19 163.367
R937 B.n21 B.n20 163.367
R938 B.n649 B.n21 163.367
R939 B.n649 B.n26 163.367
R940 B.n27 B.n26 163.367
R941 B.n28 B.n27 163.367
R942 B.n654 B.n28 163.367
R943 B.n654 B.n33 163.367
R944 B.n34 B.n33 163.367
R945 B.n35 B.n34 163.367
R946 B.n659 B.n35 163.367
R947 B.n659 B.n40 163.367
R948 B.n41 B.n40 163.367
R949 B.n42 B.n41 163.367
R950 B.n664 B.n42 163.367
R951 B.n664 B.n47 163.367
R952 B.n48 B.n47 163.367
R953 B.n49 B.n48 163.367
R954 B.n669 B.n49 163.367
R955 B.n669 B.n54 163.367
R956 B.n55 B.n54 163.367
R957 B.n56 B.n55 163.367
R958 B.n674 B.n56 163.367
R959 B.n674 B.n61 163.367
R960 B.n62 B.n61 163.367
R961 B.n63 B.n62 163.367
R962 B.n679 B.n63 163.367
R963 B.n679 B.n68 163.367
R964 B.n69 B.n68 163.367
R965 B.n70 B.n69 163.367
R966 B.n684 B.n70 163.367
R967 B.n684 B.n75 163.367
R968 B.n76 B.n75 163.367
R969 B.n77 B.n76 163.367
R970 B.n689 B.n77 163.367
R971 B.n689 B.n82 163.367
R972 B.n83 B.n82 163.367
R973 B.n84 B.n83 163.367
R974 B.n694 B.n84 163.367
R975 B.n694 B.n89 163.367
R976 B.n90 B.n89 163.367
R977 B.n91 B.n90 163.367
R978 B.n699 B.n91 163.367
R979 B.n699 B.n96 163.367
R980 B.n97 B.n96 163.367
R981 B.n98 B.n97 163.367
R982 B.n704 B.n98 163.367
R983 B.n704 B.n103 163.367
R984 B.n104 B.n103 163.367
R985 B.n105 B.n104 163.367
R986 B.n861 B.n859 163.367
R987 B.n857 B.n109 163.367
R988 B.n853 B.n851 163.367
R989 B.n849 B.n111 163.367
R990 B.n845 B.n843 163.367
R991 B.n841 B.n113 163.367
R992 B.n837 B.n835 163.367
R993 B.n833 B.n115 163.367
R994 B.n829 B.n827 163.367
R995 B.n825 B.n117 163.367
R996 B.n821 B.n819 163.367
R997 B.n817 B.n119 163.367
R998 B.n813 B.n811 163.367
R999 B.n809 B.n121 163.367
R1000 B.n805 B.n803 163.367
R1001 B.n801 B.n123 163.367
R1002 B.n797 B.n795 163.367
R1003 B.n792 B.n791 163.367
R1004 B.n789 B.n129 163.367
R1005 B.n785 B.n783 163.367
R1006 B.n781 B.n131 163.367
R1007 B.n776 B.n774 163.367
R1008 B.n772 B.n135 163.367
R1009 B.n768 B.n766 163.367
R1010 B.n764 B.n137 163.367
R1011 B.n760 B.n758 163.367
R1012 B.n756 B.n139 163.367
R1013 B.n752 B.n750 163.367
R1014 B.n748 B.n141 163.367
R1015 B.n744 B.n742 163.367
R1016 B.n740 B.n143 163.367
R1017 B.n736 B.n734 163.367
R1018 B.n732 B.n145 163.367
R1019 B.n728 B.n726 163.367
R1020 B.n724 B.n147 163.367
R1021 B.n720 B.n718 163.367
R1022 B.n716 B.n149 163.367
R1023 B.n712 B.n710 163.367
R1024 B.n463 B.n264 104.263
R1025 B.n866 B.n106 104.263
R1026 B.n292 B.n291 82.6187
R1027 B.n285 B.n284 82.6187
R1028 B.n125 B.n124 82.6187
R1029 B.n133 B.n132 82.6187
R1030 B.n457 B.n265 71.676
R1031 B.n455 B.n267 71.676
R1032 B.n451 B.n450 71.676
R1033 B.n444 B.n269 71.676
R1034 B.n443 B.n442 71.676
R1035 B.n436 B.n271 71.676
R1036 B.n435 B.n434 71.676
R1037 B.n428 B.n273 71.676
R1038 B.n427 B.n426 71.676
R1039 B.n420 B.n275 71.676
R1040 B.n419 B.n418 71.676
R1041 B.n412 B.n277 71.676
R1042 B.n411 B.n410 71.676
R1043 B.n404 B.n279 71.676
R1044 B.n403 B.n402 71.676
R1045 B.n396 B.n281 71.676
R1046 B.n395 B.n394 71.676
R1047 B.n388 B.n283 71.676
R1048 B.n387 B.n386 71.676
R1049 B.n380 B.n288 71.676
R1050 B.n379 B.n378 71.676
R1051 B.n371 B.n290 71.676
R1052 B.n370 B.n369 71.676
R1053 B.n363 B.n294 71.676
R1054 B.n362 B.n361 71.676
R1055 B.n355 B.n296 71.676
R1056 B.n354 B.n353 71.676
R1057 B.n347 B.n298 71.676
R1058 B.n346 B.n345 71.676
R1059 B.n339 B.n300 71.676
R1060 B.n338 B.n337 71.676
R1061 B.n331 B.n302 71.676
R1062 B.n330 B.n329 71.676
R1063 B.n323 B.n304 71.676
R1064 B.n322 B.n321 71.676
R1065 B.n315 B.n306 71.676
R1066 B.n314 B.n313 71.676
R1067 B.n309 B.n308 71.676
R1068 B.n860 B.n107 71.676
R1069 B.n859 B.n858 71.676
R1070 B.n852 B.n109 71.676
R1071 B.n851 B.n850 71.676
R1072 B.n844 B.n111 71.676
R1073 B.n843 B.n842 71.676
R1074 B.n836 B.n113 71.676
R1075 B.n835 B.n834 71.676
R1076 B.n828 B.n115 71.676
R1077 B.n827 B.n826 71.676
R1078 B.n820 B.n117 71.676
R1079 B.n819 B.n818 71.676
R1080 B.n812 B.n119 71.676
R1081 B.n811 B.n810 71.676
R1082 B.n804 B.n121 71.676
R1083 B.n803 B.n802 71.676
R1084 B.n796 B.n123 71.676
R1085 B.n795 B.n127 71.676
R1086 B.n791 B.n790 71.676
R1087 B.n784 B.n129 71.676
R1088 B.n783 B.n782 71.676
R1089 B.n775 B.n131 71.676
R1090 B.n774 B.n773 71.676
R1091 B.n767 B.n135 71.676
R1092 B.n766 B.n765 71.676
R1093 B.n759 B.n137 71.676
R1094 B.n758 B.n757 71.676
R1095 B.n751 B.n139 71.676
R1096 B.n750 B.n749 71.676
R1097 B.n743 B.n141 71.676
R1098 B.n742 B.n741 71.676
R1099 B.n735 B.n143 71.676
R1100 B.n734 B.n733 71.676
R1101 B.n727 B.n145 71.676
R1102 B.n726 B.n725 71.676
R1103 B.n719 B.n147 71.676
R1104 B.n718 B.n717 71.676
R1105 B.n711 B.n149 71.676
R1106 B.n712 B.n711 71.676
R1107 B.n717 B.n716 71.676
R1108 B.n720 B.n719 71.676
R1109 B.n725 B.n724 71.676
R1110 B.n728 B.n727 71.676
R1111 B.n733 B.n732 71.676
R1112 B.n736 B.n735 71.676
R1113 B.n741 B.n740 71.676
R1114 B.n744 B.n743 71.676
R1115 B.n749 B.n748 71.676
R1116 B.n752 B.n751 71.676
R1117 B.n757 B.n756 71.676
R1118 B.n760 B.n759 71.676
R1119 B.n765 B.n764 71.676
R1120 B.n768 B.n767 71.676
R1121 B.n773 B.n772 71.676
R1122 B.n776 B.n775 71.676
R1123 B.n782 B.n781 71.676
R1124 B.n785 B.n784 71.676
R1125 B.n790 B.n789 71.676
R1126 B.n792 B.n127 71.676
R1127 B.n797 B.n796 71.676
R1128 B.n802 B.n801 71.676
R1129 B.n805 B.n804 71.676
R1130 B.n810 B.n809 71.676
R1131 B.n813 B.n812 71.676
R1132 B.n818 B.n817 71.676
R1133 B.n821 B.n820 71.676
R1134 B.n826 B.n825 71.676
R1135 B.n829 B.n828 71.676
R1136 B.n834 B.n833 71.676
R1137 B.n837 B.n836 71.676
R1138 B.n842 B.n841 71.676
R1139 B.n845 B.n844 71.676
R1140 B.n850 B.n849 71.676
R1141 B.n853 B.n852 71.676
R1142 B.n858 B.n857 71.676
R1143 B.n861 B.n860 71.676
R1144 B.n458 B.n457 71.676
R1145 B.n452 B.n267 71.676
R1146 B.n450 B.n449 71.676
R1147 B.n445 B.n444 71.676
R1148 B.n442 B.n441 71.676
R1149 B.n437 B.n436 71.676
R1150 B.n434 B.n433 71.676
R1151 B.n429 B.n428 71.676
R1152 B.n426 B.n425 71.676
R1153 B.n421 B.n420 71.676
R1154 B.n418 B.n417 71.676
R1155 B.n413 B.n412 71.676
R1156 B.n410 B.n409 71.676
R1157 B.n405 B.n404 71.676
R1158 B.n402 B.n401 71.676
R1159 B.n397 B.n396 71.676
R1160 B.n394 B.n393 71.676
R1161 B.n389 B.n388 71.676
R1162 B.n386 B.n385 71.676
R1163 B.n381 B.n380 71.676
R1164 B.n378 B.n377 71.676
R1165 B.n372 B.n371 71.676
R1166 B.n369 B.n368 71.676
R1167 B.n364 B.n363 71.676
R1168 B.n361 B.n360 71.676
R1169 B.n356 B.n355 71.676
R1170 B.n353 B.n352 71.676
R1171 B.n348 B.n347 71.676
R1172 B.n345 B.n344 71.676
R1173 B.n340 B.n339 71.676
R1174 B.n337 B.n336 71.676
R1175 B.n332 B.n331 71.676
R1176 B.n329 B.n328 71.676
R1177 B.n324 B.n323 71.676
R1178 B.n321 B.n320 71.676
R1179 B.n316 B.n315 71.676
R1180 B.n313 B.n312 71.676
R1181 B.n308 B.n263 71.676
R1182 B.n375 B.n292 59.5399
R1183 B.n286 B.n285 59.5399
R1184 B.n126 B.n125 59.5399
R1185 B.n778 B.n133 59.5399
R1186 B.n463 B.n260 51.0063
R1187 B.n469 B.n260 51.0063
R1188 B.n469 B.n256 51.0063
R1189 B.n475 B.n256 51.0063
R1190 B.n475 B.n252 51.0063
R1191 B.n481 B.n252 51.0063
R1192 B.n481 B.n247 51.0063
R1193 B.n487 B.n247 51.0063
R1194 B.n487 B.n248 51.0063
R1195 B.n493 B.n240 51.0063
R1196 B.n499 B.n240 51.0063
R1197 B.n499 B.n236 51.0063
R1198 B.n505 B.n236 51.0063
R1199 B.n505 B.n232 51.0063
R1200 B.n511 B.n232 51.0063
R1201 B.n511 B.n228 51.0063
R1202 B.n517 B.n228 51.0063
R1203 B.n517 B.n224 51.0063
R1204 B.n523 B.n224 51.0063
R1205 B.n523 B.n220 51.0063
R1206 B.n529 B.n220 51.0063
R1207 B.n529 B.n215 51.0063
R1208 B.n535 B.n215 51.0063
R1209 B.n535 B.n216 51.0063
R1210 B.n541 B.n208 51.0063
R1211 B.n547 B.n208 51.0063
R1212 B.n547 B.n204 51.0063
R1213 B.n553 B.n204 51.0063
R1214 B.n553 B.n200 51.0063
R1215 B.n559 B.n200 51.0063
R1216 B.n559 B.n196 51.0063
R1217 B.n565 B.n196 51.0063
R1218 B.n565 B.n191 51.0063
R1219 B.n571 B.n191 51.0063
R1220 B.n571 B.n192 51.0063
R1221 B.n577 B.n184 51.0063
R1222 B.n583 B.n184 51.0063
R1223 B.n583 B.n180 51.0063
R1224 B.n589 B.n180 51.0063
R1225 B.n589 B.n176 51.0063
R1226 B.n595 B.n176 51.0063
R1227 B.n595 B.n172 51.0063
R1228 B.n601 B.n172 51.0063
R1229 B.n601 B.n168 51.0063
R1230 B.n607 B.n168 51.0063
R1231 B.n607 B.n164 51.0063
R1232 B.n613 B.n164 51.0063
R1233 B.n619 B.n160 51.0063
R1234 B.n619 B.n156 51.0063
R1235 B.n626 B.n156 51.0063
R1236 B.n626 B.n152 51.0063
R1237 B.n632 B.n152 51.0063
R1238 B.n632 B.n4 51.0063
R1239 B.n980 B.n4 51.0063
R1240 B.n980 B.n979 51.0063
R1241 B.n979 B.n978 51.0063
R1242 B.n978 B.n8 51.0063
R1243 B.n972 B.n8 51.0063
R1244 B.n972 B.n971 51.0063
R1245 B.n971 B.n970 51.0063
R1246 B.n970 B.n15 51.0063
R1247 B.n964 B.n963 51.0063
R1248 B.n963 B.n962 51.0063
R1249 B.n962 B.n22 51.0063
R1250 B.n956 B.n22 51.0063
R1251 B.n956 B.n955 51.0063
R1252 B.n955 B.n954 51.0063
R1253 B.n954 B.n29 51.0063
R1254 B.n948 B.n29 51.0063
R1255 B.n948 B.n947 51.0063
R1256 B.n947 B.n946 51.0063
R1257 B.n946 B.n36 51.0063
R1258 B.n940 B.n36 51.0063
R1259 B.n939 B.n938 51.0063
R1260 B.n938 B.n43 51.0063
R1261 B.n932 B.n43 51.0063
R1262 B.n932 B.n931 51.0063
R1263 B.n931 B.n930 51.0063
R1264 B.n930 B.n50 51.0063
R1265 B.n924 B.n50 51.0063
R1266 B.n924 B.n923 51.0063
R1267 B.n923 B.n922 51.0063
R1268 B.n922 B.n57 51.0063
R1269 B.n916 B.n57 51.0063
R1270 B.n915 B.n914 51.0063
R1271 B.n914 B.n64 51.0063
R1272 B.n908 B.n64 51.0063
R1273 B.n908 B.n907 51.0063
R1274 B.n907 B.n906 51.0063
R1275 B.n906 B.n71 51.0063
R1276 B.n900 B.n71 51.0063
R1277 B.n900 B.n899 51.0063
R1278 B.n899 B.n898 51.0063
R1279 B.n898 B.n78 51.0063
R1280 B.n892 B.n78 51.0063
R1281 B.n892 B.n891 51.0063
R1282 B.n891 B.n890 51.0063
R1283 B.n890 B.n85 51.0063
R1284 B.n884 B.n85 51.0063
R1285 B.n883 B.n882 51.0063
R1286 B.n882 B.n92 51.0063
R1287 B.n876 B.n92 51.0063
R1288 B.n876 B.n875 51.0063
R1289 B.n875 B.n874 51.0063
R1290 B.n874 B.n99 51.0063
R1291 B.n868 B.n99 51.0063
R1292 B.n868 B.n867 51.0063
R1293 B.n867 B.n866 51.0063
R1294 B.n541 B.t3 47.2559
R1295 B.n916 B.t1 47.2559
R1296 B.t2 B.n160 44.2555
R1297 B.t0 B.n15 44.2555
R1298 B.n864 B.n863 37.3078
R1299 B.n709 B.n708 37.3078
R1300 B.n465 B.n262 37.3078
R1301 B.n461 B.n460 37.3078
R1302 B.n493 B.t7 33.7543
R1303 B.n884 B.t11 33.7543
R1304 B.n192 B.t5 30.754
R1305 B.t4 B.n939 30.754
R1306 B.n577 B.t5 20.2528
R1307 B.n940 B.t4 20.2528
R1308 B B.n982 18.0485
R1309 B.n248 B.t7 17.2525
R1310 B.t11 B.n883 17.2525
R1311 B.n863 B.n862 10.6151
R1312 B.n862 B.n108 10.6151
R1313 B.n856 B.n108 10.6151
R1314 B.n856 B.n855 10.6151
R1315 B.n855 B.n854 10.6151
R1316 B.n854 B.n110 10.6151
R1317 B.n848 B.n110 10.6151
R1318 B.n848 B.n847 10.6151
R1319 B.n847 B.n846 10.6151
R1320 B.n846 B.n112 10.6151
R1321 B.n840 B.n112 10.6151
R1322 B.n840 B.n839 10.6151
R1323 B.n839 B.n838 10.6151
R1324 B.n838 B.n114 10.6151
R1325 B.n832 B.n114 10.6151
R1326 B.n832 B.n831 10.6151
R1327 B.n831 B.n830 10.6151
R1328 B.n830 B.n116 10.6151
R1329 B.n824 B.n116 10.6151
R1330 B.n824 B.n823 10.6151
R1331 B.n823 B.n822 10.6151
R1332 B.n822 B.n118 10.6151
R1333 B.n816 B.n118 10.6151
R1334 B.n816 B.n815 10.6151
R1335 B.n815 B.n814 10.6151
R1336 B.n814 B.n120 10.6151
R1337 B.n808 B.n120 10.6151
R1338 B.n808 B.n807 10.6151
R1339 B.n807 B.n806 10.6151
R1340 B.n806 B.n122 10.6151
R1341 B.n800 B.n122 10.6151
R1342 B.n800 B.n799 10.6151
R1343 B.n799 B.n798 10.6151
R1344 B.n794 B.n793 10.6151
R1345 B.n793 B.n128 10.6151
R1346 B.n788 B.n128 10.6151
R1347 B.n788 B.n787 10.6151
R1348 B.n787 B.n786 10.6151
R1349 B.n786 B.n130 10.6151
R1350 B.n780 B.n130 10.6151
R1351 B.n780 B.n779 10.6151
R1352 B.n777 B.n134 10.6151
R1353 B.n771 B.n134 10.6151
R1354 B.n771 B.n770 10.6151
R1355 B.n770 B.n769 10.6151
R1356 B.n769 B.n136 10.6151
R1357 B.n763 B.n136 10.6151
R1358 B.n763 B.n762 10.6151
R1359 B.n762 B.n761 10.6151
R1360 B.n761 B.n138 10.6151
R1361 B.n755 B.n138 10.6151
R1362 B.n755 B.n754 10.6151
R1363 B.n754 B.n753 10.6151
R1364 B.n753 B.n140 10.6151
R1365 B.n747 B.n140 10.6151
R1366 B.n747 B.n746 10.6151
R1367 B.n746 B.n745 10.6151
R1368 B.n745 B.n142 10.6151
R1369 B.n739 B.n142 10.6151
R1370 B.n739 B.n738 10.6151
R1371 B.n738 B.n737 10.6151
R1372 B.n737 B.n144 10.6151
R1373 B.n731 B.n144 10.6151
R1374 B.n731 B.n730 10.6151
R1375 B.n730 B.n729 10.6151
R1376 B.n729 B.n146 10.6151
R1377 B.n723 B.n146 10.6151
R1378 B.n723 B.n722 10.6151
R1379 B.n722 B.n721 10.6151
R1380 B.n721 B.n148 10.6151
R1381 B.n715 B.n148 10.6151
R1382 B.n715 B.n714 10.6151
R1383 B.n714 B.n713 10.6151
R1384 B.n713 B.n709 10.6151
R1385 B.n466 B.n465 10.6151
R1386 B.n467 B.n466 10.6151
R1387 B.n467 B.n254 10.6151
R1388 B.n477 B.n254 10.6151
R1389 B.n478 B.n477 10.6151
R1390 B.n479 B.n478 10.6151
R1391 B.n479 B.n245 10.6151
R1392 B.n489 B.n245 10.6151
R1393 B.n490 B.n489 10.6151
R1394 B.n491 B.n490 10.6151
R1395 B.n491 B.n238 10.6151
R1396 B.n501 B.n238 10.6151
R1397 B.n502 B.n501 10.6151
R1398 B.n503 B.n502 10.6151
R1399 B.n503 B.n230 10.6151
R1400 B.n513 B.n230 10.6151
R1401 B.n514 B.n513 10.6151
R1402 B.n515 B.n514 10.6151
R1403 B.n515 B.n222 10.6151
R1404 B.n525 B.n222 10.6151
R1405 B.n526 B.n525 10.6151
R1406 B.n527 B.n526 10.6151
R1407 B.n527 B.n213 10.6151
R1408 B.n537 B.n213 10.6151
R1409 B.n538 B.n537 10.6151
R1410 B.n539 B.n538 10.6151
R1411 B.n539 B.n206 10.6151
R1412 B.n549 B.n206 10.6151
R1413 B.n550 B.n549 10.6151
R1414 B.n551 B.n550 10.6151
R1415 B.n551 B.n198 10.6151
R1416 B.n561 B.n198 10.6151
R1417 B.n562 B.n561 10.6151
R1418 B.n563 B.n562 10.6151
R1419 B.n563 B.n189 10.6151
R1420 B.n573 B.n189 10.6151
R1421 B.n574 B.n573 10.6151
R1422 B.n575 B.n574 10.6151
R1423 B.n575 B.n182 10.6151
R1424 B.n585 B.n182 10.6151
R1425 B.n586 B.n585 10.6151
R1426 B.n587 B.n586 10.6151
R1427 B.n587 B.n174 10.6151
R1428 B.n597 B.n174 10.6151
R1429 B.n598 B.n597 10.6151
R1430 B.n599 B.n598 10.6151
R1431 B.n599 B.n166 10.6151
R1432 B.n609 B.n166 10.6151
R1433 B.n610 B.n609 10.6151
R1434 B.n611 B.n610 10.6151
R1435 B.n611 B.n158 10.6151
R1436 B.n621 B.n158 10.6151
R1437 B.n622 B.n621 10.6151
R1438 B.n624 B.n622 10.6151
R1439 B.n624 B.n623 10.6151
R1440 B.n623 B.n150 10.6151
R1441 B.n635 B.n150 10.6151
R1442 B.n636 B.n635 10.6151
R1443 B.n637 B.n636 10.6151
R1444 B.n638 B.n637 10.6151
R1445 B.n640 B.n638 10.6151
R1446 B.n641 B.n640 10.6151
R1447 B.n642 B.n641 10.6151
R1448 B.n643 B.n642 10.6151
R1449 B.n645 B.n643 10.6151
R1450 B.n646 B.n645 10.6151
R1451 B.n647 B.n646 10.6151
R1452 B.n648 B.n647 10.6151
R1453 B.n650 B.n648 10.6151
R1454 B.n651 B.n650 10.6151
R1455 B.n652 B.n651 10.6151
R1456 B.n653 B.n652 10.6151
R1457 B.n655 B.n653 10.6151
R1458 B.n656 B.n655 10.6151
R1459 B.n657 B.n656 10.6151
R1460 B.n658 B.n657 10.6151
R1461 B.n660 B.n658 10.6151
R1462 B.n661 B.n660 10.6151
R1463 B.n662 B.n661 10.6151
R1464 B.n663 B.n662 10.6151
R1465 B.n665 B.n663 10.6151
R1466 B.n666 B.n665 10.6151
R1467 B.n667 B.n666 10.6151
R1468 B.n668 B.n667 10.6151
R1469 B.n670 B.n668 10.6151
R1470 B.n671 B.n670 10.6151
R1471 B.n672 B.n671 10.6151
R1472 B.n673 B.n672 10.6151
R1473 B.n675 B.n673 10.6151
R1474 B.n676 B.n675 10.6151
R1475 B.n677 B.n676 10.6151
R1476 B.n678 B.n677 10.6151
R1477 B.n680 B.n678 10.6151
R1478 B.n681 B.n680 10.6151
R1479 B.n682 B.n681 10.6151
R1480 B.n683 B.n682 10.6151
R1481 B.n685 B.n683 10.6151
R1482 B.n686 B.n685 10.6151
R1483 B.n687 B.n686 10.6151
R1484 B.n688 B.n687 10.6151
R1485 B.n690 B.n688 10.6151
R1486 B.n691 B.n690 10.6151
R1487 B.n692 B.n691 10.6151
R1488 B.n693 B.n692 10.6151
R1489 B.n695 B.n693 10.6151
R1490 B.n696 B.n695 10.6151
R1491 B.n697 B.n696 10.6151
R1492 B.n698 B.n697 10.6151
R1493 B.n700 B.n698 10.6151
R1494 B.n701 B.n700 10.6151
R1495 B.n702 B.n701 10.6151
R1496 B.n703 B.n702 10.6151
R1497 B.n705 B.n703 10.6151
R1498 B.n706 B.n705 10.6151
R1499 B.n707 B.n706 10.6151
R1500 B.n708 B.n707 10.6151
R1501 B.n460 B.n459 10.6151
R1502 B.n459 B.n266 10.6151
R1503 B.n454 B.n266 10.6151
R1504 B.n454 B.n453 10.6151
R1505 B.n453 B.n268 10.6151
R1506 B.n448 B.n268 10.6151
R1507 B.n448 B.n447 10.6151
R1508 B.n447 B.n446 10.6151
R1509 B.n446 B.n270 10.6151
R1510 B.n440 B.n270 10.6151
R1511 B.n440 B.n439 10.6151
R1512 B.n439 B.n438 10.6151
R1513 B.n438 B.n272 10.6151
R1514 B.n432 B.n272 10.6151
R1515 B.n432 B.n431 10.6151
R1516 B.n431 B.n430 10.6151
R1517 B.n430 B.n274 10.6151
R1518 B.n424 B.n274 10.6151
R1519 B.n424 B.n423 10.6151
R1520 B.n423 B.n422 10.6151
R1521 B.n422 B.n276 10.6151
R1522 B.n416 B.n276 10.6151
R1523 B.n416 B.n415 10.6151
R1524 B.n415 B.n414 10.6151
R1525 B.n414 B.n278 10.6151
R1526 B.n408 B.n278 10.6151
R1527 B.n408 B.n407 10.6151
R1528 B.n407 B.n406 10.6151
R1529 B.n406 B.n280 10.6151
R1530 B.n400 B.n280 10.6151
R1531 B.n400 B.n399 10.6151
R1532 B.n399 B.n398 10.6151
R1533 B.n398 B.n282 10.6151
R1534 B.n392 B.n391 10.6151
R1535 B.n391 B.n390 10.6151
R1536 B.n390 B.n287 10.6151
R1537 B.n384 B.n287 10.6151
R1538 B.n384 B.n383 10.6151
R1539 B.n383 B.n382 10.6151
R1540 B.n382 B.n289 10.6151
R1541 B.n376 B.n289 10.6151
R1542 B.n374 B.n373 10.6151
R1543 B.n373 B.n293 10.6151
R1544 B.n367 B.n293 10.6151
R1545 B.n367 B.n366 10.6151
R1546 B.n366 B.n365 10.6151
R1547 B.n365 B.n295 10.6151
R1548 B.n359 B.n295 10.6151
R1549 B.n359 B.n358 10.6151
R1550 B.n358 B.n357 10.6151
R1551 B.n357 B.n297 10.6151
R1552 B.n351 B.n297 10.6151
R1553 B.n351 B.n350 10.6151
R1554 B.n350 B.n349 10.6151
R1555 B.n349 B.n299 10.6151
R1556 B.n343 B.n299 10.6151
R1557 B.n343 B.n342 10.6151
R1558 B.n342 B.n341 10.6151
R1559 B.n341 B.n301 10.6151
R1560 B.n335 B.n301 10.6151
R1561 B.n335 B.n334 10.6151
R1562 B.n334 B.n333 10.6151
R1563 B.n333 B.n303 10.6151
R1564 B.n327 B.n303 10.6151
R1565 B.n327 B.n326 10.6151
R1566 B.n326 B.n325 10.6151
R1567 B.n325 B.n305 10.6151
R1568 B.n319 B.n305 10.6151
R1569 B.n319 B.n318 10.6151
R1570 B.n318 B.n317 10.6151
R1571 B.n317 B.n307 10.6151
R1572 B.n311 B.n307 10.6151
R1573 B.n311 B.n310 10.6151
R1574 B.n310 B.n262 10.6151
R1575 B.n461 B.n258 10.6151
R1576 B.n471 B.n258 10.6151
R1577 B.n472 B.n471 10.6151
R1578 B.n473 B.n472 10.6151
R1579 B.n473 B.n250 10.6151
R1580 B.n483 B.n250 10.6151
R1581 B.n484 B.n483 10.6151
R1582 B.n485 B.n484 10.6151
R1583 B.n485 B.n242 10.6151
R1584 B.n495 B.n242 10.6151
R1585 B.n496 B.n495 10.6151
R1586 B.n497 B.n496 10.6151
R1587 B.n497 B.n234 10.6151
R1588 B.n507 B.n234 10.6151
R1589 B.n508 B.n507 10.6151
R1590 B.n509 B.n508 10.6151
R1591 B.n509 B.n226 10.6151
R1592 B.n519 B.n226 10.6151
R1593 B.n520 B.n519 10.6151
R1594 B.n521 B.n520 10.6151
R1595 B.n521 B.n218 10.6151
R1596 B.n531 B.n218 10.6151
R1597 B.n532 B.n531 10.6151
R1598 B.n533 B.n532 10.6151
R1599 B.n533 B.n210 10.6151
R1600 B.n543 B.n210 10.6151
R1601 B.n544 B.n543 10.6151
R1602 B.n545 B.n544 10.6151
R1603 B.n545 B.n202 10.6151
R1604 B.n555 B.n202 10.6151
R1605 B.n556 B.n555 10.6151
R1606 B.n557 B.n556 10.6151
R1607 B.n557 B.n194 10.6151
R1608 B.n567 B.n194 10.6151
R1609 B.n568 B.n567 10.6151
R1610 B.n569 B.n568 10.6151
R1611 B.n569 B.n186 10.6151
R1612 B.n579 B.n186 10.6151
R1613 B.n580 B.n579 10.6151
R1614 B.n581 B.n580 10.6151
R1615 B.n581 B.n178 10.6151
R1616 B.n591 B.n178 10.6151
R1617 B.n592 B.n591 10.6151
R1618 B.n593 B.n592 10.6151
R1619 B.n593 B.n170 10.6151
R1620 B.n603 B.n170 10.6151
R1621 B.n604 B.n603 10.6151
R1622 B.n605 B.n604 10.6151
R1623 B.n605 B.n162 10.6151
R1624 B.n615 B.n162 10.6151
R1625 B.n616 B.n615 10.6151
R1626 B.n617 B.n616 10.6151
R1627 B.n617 B.n154 10.6151
R1628 B.n628 B.n154 10.6151
R1629 B.n629 B.n628 10.6151
R1630 B.n630 B.n629 10.6151
R1631 B.n630 B.n0 10.6151
R1632 B.n976 B.n1 10.6151
R1633 B.n976 B.n975 10.6151
R1634 B.n975 B.n974 10.6151
R1635 B.n974 B.n10 10.6151
R1636 B.n968 B.n10 10.6151
R1637 B.n968 B.n967 10.6151
R1638 B.n967 B.n966 10.6151
R1639 B.n966 B.n17 10.6151
R1640 B.n960 B.n17 10.6151
R1641 B.n960 B.n959 10.6151
R1642 B.n959 B.n958 10.6151
R1643 B.n958 B.n24 10.6151
R1644 B.n952 B.n24 10.6151
R1645 B.n952 B.n951 10.6151
R1646 B.n951 B.n950 10.6151
R1647 B.n950 B.n31 10.6151
R1648 B.n944 B.n31 10.6151
R1649 B.n944 B.n943 10.6151
R1650 B.n943 B.n942 10.6151
R1651 B.n942 B.n38 10.6151
R1652 B.n936 B.n38 10.6151
R1653 B.n936 B.n935 10.6151
R1654 B.n935 B.n934 10.6151
R1655 B.n934 B.n45 10.6151
R1656 B.n928 B.n45 10.6151
R1657 B.n928 B.n927 10.6151
R1658 B.n927 B.n926 10.6151
R1659 B.n926 B.n52 10.6151
R1660 B.n920 B.n52 10.6151
R1661 B.n920 B.n919 10.6151
R1662 B.n919 B.n918 10.6151
R1663 B.n918 B.n59 10.6151
R1664 B.n912 B.n59 10.6151
R1665 B.n912 B.n911 10.6151
R1666 B.n911 B.n910 10.6151
R1667 B.n910 B.n66 10.6151
R1668 B.n904 B.n66 10.6151
R1669 B.n904 B.n903 10.6151
R1670 B.n903 B.n902 10.6151
R1671 B.n902 B.n73 10.6151
R1672 B.n896 B.n73 10.6151
R1673 B.n896 B.n895 10.6151
R1674 B.n895 B.n894 10.6151
R1675 B.n894 B.n80 10.6151
R1676 B.n888 B.n80 10.6151
R1677 B.n888 B.n887 10.6151
R1678 B.n887 B.n886 10.6151
R1679 B.n886 B.n87 10.6151
R1680 B.n880 B.n87 10.6151
R1681 B.n880 B.n879 10.6151
R1682 B.n879 B.n878 10.6151
R1683 B.n878 B.n94 10.6151
R1684 B.n872 B.n94 10.6151
R1685 B.n872 B.n871 10.6151
R1686 B.n871 B.n870 10.6151
R1687 B.n870 B.n101 10.6151
R1688 B.n864 B.n101 10.6151
R1689 B.n613 B.t2 6.75127
R1690 B.n964 B.t0 6.75127
R1691 B.n794 B.n126 6.5566
R1692 B.n779 B.n778 6.5566
R1693 B.n392 B.n286 6.5566
R1694 B.n376 B.n375 6.5566
R1695 B.n798 B.n126 4.05904
R1696 B.n778 B.n777 4.05904
R1697 B.n286 B.n282 4.05904
R1698 B.n375 B.n374 4.05904
R1699 B.n216 B.t3 3.75093
R1700 B.t1 B.n915 3.75093
R1701 B.n982 B.n0 2.81026
R1702 B.n982 B.n1 2.81026
R1703 VN.n42 VN.n41 161.3
R1704 VN.n40 VN.n23 161.3
R1705 VN.n39 VN.n38 161.3
R1706 VN.n37 VN.n24 161.3
R1707 VN.n36 VN.n35 161.3
R1708 VN.n34 VN.n25 161.3
R1709 VN.n33 VN.n32 161.3
R1710 VN.n31 VN.n26 161.3
R1711 VN.n30 VN.n29 161.3
R1712 VN.n20 VN.n19 161.3
R1713 VN.n18 VN.n1 161.3
R1714 VN.n17 VN.n16 161.3
R1715 VN.n15 VN.n2 161.3
R1716 VN.n14 VN.n13 161.3
R1717 VN.n12 VN.n3 161.3
R1718 VN.n11 VN.n10 161.3
R1719 VN.n9 VN.n4 161.3
R1720 VN.n8 VN.n7 161.3
R1721 VN.n27 VN.t5 89.7239
R1722 VN.n5 VN.t4 89.7239
R1723 VN.n21 VN.n0 89.5781
R1724 VN.n43 VN.n22 89.5781
R1725 VN.n6 VN.n5 62.9256
R1726 VN.n28 VN.n27 62.9256
R1727 VN.n6 VN.t0 57.5829
R1728 VN.n0 VN.t3 57.5829
R1729 VN.n28 VN.t1 57.5829
R1730 VN.n22 VN.t2 57.5829
R1731 VN.n13 VN.n12 52.1486
R1732 VN.n35 VN.n34 52.1486
R1733 VN VN.n43 52.1268
R1734 VN.n13 VN.n2 28.8382
R1735 VN.n35 VN.n24 28.8382
R1736 VN.n7 VN.n4 24.4675
R1737 VN.n11 VN.n4 24.4675
R1738 VN.n12 VN.n11 24.4675
R1739 VN.n17 VN.n2 24.4675
R1740 VN.n18 VN.n17 24.4675
R1741 VN.n19 VN.n18 24.4675
R1742 VN.n34 VN.n33 24.4675
R1743 VN.n33 VN.n26 24.4675
R1744 VN.n29 VN.n26 24.4675
R1745 VN.n41 VN.n40 24.4675
R1746 VN.n40 VN.n39 24.4675
R1747 VN.n39 VN.n24 24.4675
R1748 VN.n7 VN.n6 12.234
R1749 VN.n29 VN.n28 12.234
R1750 VN.n30 VN.n27 2.52278
R1751 VN.n8 VN.n5 2.52278
R1752 VN.n19 VN.n0 0.48984
R1753 VN.n41 VN.n22 0.48984
R1754 VN.n43 VN.n42 0.354971
R1755 VN.n21 VN.n20 0.354971
R1756 VN VN.n21 0.26696
R1757 VN.n42 VN.n23 0.189894
R1758 VN.n38 VN.n23 0.189894
R1759 VN.n38 VN.n37 0.189894
R1760 VN.n37 VN.n36 0.189894
R1761 VN.n36 VN.n25 0.189894
R1762 VN.n32 VN.n25 0.189894
R1763 VN.n32 VN.n31 0.189894
R1764 VN.n31 VN.n30 0.189894
R1765 VN.n9 VN.n8 0.189894
R1766 VN.n10 VN.n9 0.189894
R1767 VN.n10 VN.n3 0.189894
R1768 VN.n14 VN.n3 0.189894
R1769 VN.n15 VN.n14 0.189894
R1770 VN.n16 VN.n15 0.189894
R1771 VN.n16 VN.n1 0.189894
R1772 VN.n20 VN.n1 0.189894
R1773 VDD2.n95 VDD2.n51 289.615
R1774 VDD2.n44 VDD2.n0 289.615
R1775 VDD2.n96 VDD2.n95 185
R1776 VDD2.n94 VDD2.n93 185
R1777 VDD2.n55 VDD2.n54 185
R1778 VDD2.n59 VDD2.n57 185
R1779 VDD2.n88 VDD2.n87 185
R1780 VDD2.n86 VDD2.n85 185
R1781 VDD2.n61 VDD2.n60 185
R1782 VDD2.n80 VDD2.n79 185
R1783 VDD2.n78 VDD2.n77 185
R1784 VDD2.n65 VDD2.n64 185
R1785 VDD2.n72 VDD2.n71 185
R1786 VDD2.n70 VDD2.n69 185
R1787 VDD2.n17 VDD2.n16 185
R1788 VDD2.n19 VDD2.n18 185
R1789 VDD2.n12 VDD2.n11 185
R1790 VDD2.n25 VDD2.n24 185
R1791 VDD2.n27 VDD2.n26 185
R1792 VDD2.n8 VDD2.n7 185
R1793 VDD2.n34 VDD2.n33 185
R1794 VDD2.n35 VDD2.n6 185
R1795 VDD2.n37 VDD2.n36 185
R1796 VDD2.n4 VDD2.n3 185
R1797 VDD2.n43 VDD2.n42 185
R1798 VDD2.n45 VDD2.n44 185
R1799 VDD2.n68 VDD2.t2 149.524
R1800 VDD2.n15 VDD2.t4 149.524
R1801 VDD2.n95 VDD2.n94 104.615
R1802 VDD2.n94 VDD2.n54 104.615
R1803 VDD2.n59 VDD2.n54 104.615
R1804 VDD2.n87 VDD2.n59 104.615
R1805 VDD2.n87 VDD2.n86 104.615
R1806 VDD2.n86 VDD2.n60 104.615
R1807 VDD2.n79 VDD2.n60 104.615
R1808 VDD2.n79 VDD2.n78 104.615
R1809 VDD2.n78 VDD2.n64 104.615
R1810 VDD2.n71 VDD2.n64 104.615
R1811 VDD2.n71 VDD2.n70 104.615
R1812 VDD2.n18 VDD2.n17 104.615
R1813 VDD2.n18 VDD2.n11 104.615
R1814 VDD2.n25 VDD2.n11 104.615
R1815 VDD2.n26 VDD2.n25 104.615
R1816 VDD2.n26 VDD2.n7 104.615
R1817 VDD2.n34 VDD2.n7 104.615
R1818 VDD2.n35 VDD2.n34 104.615
R1819 VDD2.n36 VDD2.n35 104.615
R1820 VDD2.n36 VDD2.n3 104.615
R1821 VDD2.n43 VDD2.n3 104.615
R1822 VDD2.n44 VDD2.n43 104.615
R1823 VDD2.n50 VDD2.n49 66.7737
R1824 VDD2 VDD2.n101 66.7709
R1825 VDD2.n50 VDD2.n48 54.4722
R1826 VDD2.n70 VDD2.t2 52.3082
R1827 VDD2.n17 VDD2.t4 52.3082
R1828 VDD2.n100 VDD2.n99 51.7732
R1829 VDD2.n100 VDD2.n50 43.7455
R1830 VDD2.n57 VDD2.n55 13.1884
R1831 VDD2.n37 VDD2.n4 13.1884
R1832 VDD2.n93 VDD2.n92 12.8005
R1833 VDD2.n89 VDD2.n88 12.8005
R1834 VDD2.n38 VDD2.n6 12.8005
R1835 VDD2.n42 VDD2.n41 12.8005
R1836 VDD2.n96 VDD2.n53 12.0247
R1837 VDD2.n85 VDD2.n58 12.0247
R1838 VDD2.n33 VDD2.n32 12.0247
R1839 VDD2.n45 VDD2.n2 12.0247
R1840 VDD2.n97 VDD2.n51 11.249
R1841 VDD2.n84 VDD2.n61 11.249
R1842 VDD2.n31 VDD2.n8 11.249
R1843 VDD2.n46 VDD2.n0 11.249
R1844 VDD2.n81 VDD2.n80 10.4732
R1845 VDD2.n28 VDD2.n27 10.4732
R1846 VDD2.n69 VDD2.n68 10.2747
R1847 VDD2.n16 VDD2.n15 10.2747
R1848 VDD2.n77 VDD2.n63 9.69747
R1849 VDD2.n24 VDD2.n10 9.69747
R1850 VDD2.n99 VDD2.n98 9.45567
R1851 VDD2.n48 VDD2.n47 9.45567
R1852 VDD2.n67 VDD2.n66 9.3005
R1853 VDD2.n74 VDD2.n73 9.3005
R1854 VDD2.n76 VDD2.n75 9.3005
R1855 VDD2.n63 VDD2.n62 9.3005
R1856 VDD2.n82 VDD2.n81 9.3005
R1857 VDD2.n84 VDD2.n83 9.3005
R1858 VDD2.n58 VDD2.n56 9.3005
R1859 VDD2.n90 VDD2.n89 9.3005
R1860 VDD2.n98 VDD2.n97 9.3005
R1861 VDD2.n53 VDD2.n52 9.3005
R1862 VDD2.n92 VDD2.n91 9.3005
R1863 VDD2.n47 VDD2.n46 9.3005
R1864 VDD2.n2 VDD2.n1 9.3005
R1865 VDD2.n41 VDD2.n40 9.3005
R1866 VDD2.n14 VDD2.n13 9.3005
R1867 VDD2.n21 VDD2.n20 9.3005
R1868 VDD2.n23 VDD2.n22 9.3005
R1869 VDD2.n10 VDD2.n9 9.3005
R1870 VDD2.n29 VDD2.n28 9.3005
R1871 VDD2.n31 VDD2.n30 9.3005
R1872 VDD2.n32 VDD2.n5 9.3005
R1873 VDD2.n39 VDD2.n38 9.3005
R1874 VDD2.n76 VDD2.n65 8.92171
R1875 VDD2.n23 VDD2.n12 8.92171
R1876 VDD2.n73 VDD2.n72 8.14595
R1877 VDD2.n20 VDD2.n19 8.14595
R1878 VDD2.n69 VDD2.n67 7.3702
R1879 VDD2.n16 VDD2.n14 7.3702
R1880 VDD2.n72 VDD2.n67 5.81868
R1881 VDD2.n19 VDD2.n14 5.81868
R1882 VDD2.n73 VDD2.n65 5.04292
R1883 VDD2.n20 VDD2.n12 5.04292
R1884 VDD2.n77 VDD2.n76 4.26717
R1885 VDD2.n24 VDD2.n23 4.26717
R1886 VDD2.n80 VDD2.n63 3.49141
R1887 VDD2.n27 VDD2.n10 3.49141
R1888 VDD2.n68 VDD2.n66 2.84303
R1889 VDD2.n15 VDD2.n13 2.84303
R1890 VDD2 VDD2.n100 2.813
R1891 VDD2.n99 VDD2.n51 2.71565
R1892 VDD2.n81 VDD2.n61 2.71565
R1893 VDD2.n28 VDD2.n8 2.71565
R1894 VDD2.n48 VDD2.n0 2.71565
R1895 VDD2.n101 VDD2.t1 2.10913
R1896 VDD2.n101 VDD2.t5 2.10913
R1897 VDD2.n49 VDD2.t0 2.10913
R1898 VDD2.n49 VDD2.t3 2.10913
R1899 VDD2.n97 VDD2.n96 1.93989
R1900 VDD2.n85 VDD2.n84 1.93989
R1901 VDD2.n33 VDD2.n31 1.93989
R1902 VDD2.n46 VDD2.n45 1.93989
R1903 VDD2.n93 VDD2.n53 1.16414
R1904 VDD2.n88 VDD2.n58 1.16414
R1905 VDD2.n32 VDD2.n6 1.16414
R1906 VDD2.n42 VDD2.n2 1.16414
R1907 VDD2.n92 VDD2.n55 0.388379
R1908 VDD2.n89 VDD2.n57 0.388379
R1909 VDD2.n38 VDD2.n37 0.388379
R1910 VDD2.n41 VDD2.n4 0.388379
R1911 VDD2.n98 VDD2.n52 0.155672
R1912 VDD2.n91 VDD2.n52 0.155672
R1913 VDD2.n91 VDD2.n90 0.155672
R1914 VDD2.n90 VDD2.n56 0.155672
R1915 VDD2.n83 VDD2.n56 0.155672
R1916 VDD2.n83 VDD2.n82 0.155672
R1917 VDD2.n82 VDD2.n62 0.155672
R1918 VDD2.n75 VDD2.n62 0.155672
R1919 VDD2.n75 VDD2.n74 0.155672
R1920 VDD2.n74 VDD2.n66 0.155672
R1921 VDD2.n21 VDD2.n13 0.155672
R1922 VDD2.n22 VDD2.n21 0.155672
R1923 VDD2.n22 VDD2.n9 0.155672
R1924 VDD2.n29 VDD2.n9 0.155672
R1925 VDD2.n30 VDD2.n29 0.155672
R1926 VDD2.n30 VDD2.n5 0.155672
R1927 VDD2.n39 VDD2.n5 0.155672
R1928 VDD2.n40 VDD2.n39 0.155672
R1929 VDD2.n40 VDD2.n1 0.155672
R1930 VDD2.n47 VDD2.n1 0.155672
R1931 VTAIL.n202 VTAIL.n158 289.615
R1932 VTAIL.n46 VTAIL.n2 289.615
R1933 VTAIL.n152 VTAIL.n108 289.615
R1934 VTAIL.n100 VTAIL.n56 289.615
R1935 VTAIL.n175 VTAIL.n174 185
R1936 VTAIL.n177 VTAIL.n176 185
R1937 VTAIL.n170 VTAIL.n169 185
R1938 VTAIL.n183 VTAIL.n182 185
R1939 VTAIL.n185 VTAIL.n184 185
R1940 VTAIL.n166 VTAIL.n165 185
R1941 VTAIL.n192 VTAIL.n191 185
R1942 VTAIL.n193 VTAIL.n164 185
R1943 VTAIL.n195 VTAIL.n194 185
R1944 VTAIL.n162 VTAIL.n161 185
R1945 VTAIL.n201 VTAIL.n200 185
R1946 VTAIL.n203 VTAIL.n202 185
R1947 VTAIL.n19 VTAIL.n18 185
R1948 VTAIL.n21 VTAIL.n20 185
R1949 VTAIL.n14 VTAIL.n13 185
R1950 VTAIL.n27 VTAIL.n26 185
R1951 VTAIL.n29 VTAIL.n28 185
R1952 VTAIL.n10 VTAIL.n9 185
R1953 VTAIL.n36 VTAIL.n35 185
R1954 VTAIL.n37 VTAIL.n8 185
R1955 VTAIL.n39 VTAIL.n38 185
R1956 VTAIL.n6 VTAIL.n5 185
R1957 VTAIL.n45 VTAIL.n44 185
R1958 VTAIL.n47 VTAIL.n46 185
R1959 VTAIL.n153 VTAIL.n152 185
R1960 VTAIL.n151 VTAIL.n150 185
R1961 VTAIL.n112 VTAIL.n111 185
R1962 VTAIL.n116 VTAIL.n114 185
R1963 VTAIL.n145 VTAIL.n144 185
R1964 VTAIL.n143 VTAIL.n142 185
R1965 VTAIL.n118 VTAIL.n117 185
R1966 VTAIL.n137 VTAIL.n136 185
R1967 VTAIL.n135 VTAIL.n134 185
R1968 VTAIL.n122 VTAIL.n121 185
R1969 VTAIL.n129 VTAIL.n128 185
R1970 VTAIL.n127 VTAIL.n126 185
R1971 VTAIL.n101 VTAIL.n100 185
R1972 VTAIL.n99 VTAIL.n98 185
R1973 VTAIL.n60 VTAIL.n59 185
R1974 VTAIL.n64 VTAIL.n62 185
R1975 VTAIL.n93 VTAIL.n92 185
R1976 VTAIL.n91 VTAIL.n90 185
R1977 VTAIL.n66 VTAIL.n65 185
R1978 VTAIL.n85 VTAIL.n84 185
R1979 VTAIL.n83 VTAIL.n82 185
R1980 VTAIL.n70 VTAIL.n69 185
R1981 VTAIL.n77 VTAIL.n76 185
R1982 VTAIL.n75 VTAIL.n74 185
R1983 VTAIL.n173 VTAIL.t5 149.524
R1984 VTAIL.n17 VTAIL.t2 149.524
R1985 VTAIL.n125 VTAIL.t0 149.524
R1986 VTAIL.n73 VTAIL.t3 149.524
R1987 VTAIL.n176 VTAIL.n175 104.615
R1988 VTAIL.n176 VTAIL.n169 104.615
R1989 VTAIL.n183 VTAIL.n169 104.615
R1990 VTAIL.n184 VTAIL.n183 104.615
R1991 VTAIL.n184 VTAIL.n165 104.615
R1992 VTAIL.n192 VTAIL.n165 104.615
R1993 VTAIL.n193 VTAIL.n192 104.615
R1994 VTAIL.n194 VTAIL.n193 104.615
R1995 VTAIL.n194 VTAIL.n161 104.615
R1996 VTAIL.n201 VTAIL.n161 104.615
R1997 VTAIL.n202 VTAIL.n201 104.615
R1998 VTAIL.n20 VTAIL.n19 104.615
R1999 VTAIL.n20 VTAIL.n13 104.615
R2000 VTAIL.n27 VTAIL.n13 104.615
R2001 VTAIL.n28 VTAIL.n27 104.615
R2002 VTAIL.n28 VTAIL.n9 104.615
R2003 VTAIL.n36 VTAIL.n9 104.615
R2004 VTAIL.n37 VTAIL.n36 104.615
R2005 VTAIL.n38 VTAIL.n37 104.615
R2006 VTAIL.n38 VTAIL.n5 104.615
R2007 VTAIL.n45 VTAIL.n5 104.615
R2008 VTAIL.n46 VTAIL.n45 104.615
R2009 VTAIL.n152 VTAIL.n151 104.615
R2010 VTAIL.n151 VTAIL.n111 104.615
R2011 VTAIL.n116 VTAIL.n111 104.615
R2012 VTAIL.n144 VTAIL.n116 104.615
R2013 VTAIL.n144 VTAIL.n143 104.615
R2014 VTAIL.n143 VTAIL.n117 104.615
R2015 VTAIL.n136 VTAIL.n117 104.615
R2016 VTAIL.n136 VTAIL.n135 104.615
R2017 VTAIL.n135 VTAIL.n121 104.615
R2018 VTAIL.n128 VTAIL.n121 104.615
R2019 VTAIL.n128 VTAIL.n127 104.615
R2020 VTAIL.n100 VTAIL.n99 104.615
R2021 VTAIL.n99 VTAIL.n59 104.615
R2022 VTAIL.n64 VTAIL.n59 104.615
R2023 VTAIL.n92 VTAIL.n64 104.615
R2024 VTAIL.n92 VTAIL.n91 104.615
R2025 VTAIL.n91 VTAIL.n65 104.615
R2026 VTAIL.n84 VTAIL.n65 104.615
R2027 VTAIL.n84 VTAIL.n83 104.615
R2028 VTAIL.n83 VTAIL.n69 104.615
R2029 VTAIL.n76 VTAIL.n69 104.615
R2030 VTAIL.n76 VTAIL.n75 104.615
R2031 VTAIL.n175 VTAIL.t5 52.3082
R2032 VTAIL.n19 VTAIL.t2 52.3082
R2033 VTAIL.n127 VTAIL.t0 52.3082
R2034 VTAIL.n75 VTAIL.t3 52.3082
R2035 VTAIL.n107 VTAIL.n106 49.2323
R2036 VTAIL.n55 VTAIL.n54 49.2323
R2037 VTAIL.n1 VTAIL.n0 49.2322
R2038 VTAIL.n53 VTAIL.n52 49.2322
R2039 VTAIL.n207 VTAIL.n206 35.0944
R2040 VTAIL.n51 VTAIL.n50 35.0944
R2041 VTAIL.n157 VTAIL.n156 35.0944
R2042 VTAIL.n105 VTAIL.n104 35.0944
R2043 VTAIL.n55 VTAIL.n53 27.8065
R2044 VTAIL.n207 VTAIL.n157 24.1341
R2045 VTAIL.n195 VTAIL.n162 13.1884
R2046 VTAIL.n39 VTAIL.n6 13.1884
R2047 VTAIL.n114 VTAIL.n112 13.1884
R2048 VTAIL.n62 VTAIL.n60 13.1884
R2049 VTAIL.n196 VTAIL.n164 12.8005
R2050 VTAIL.n200 VTAIL.n199 12.8005
R2051 VTAIL.n40 VTAIL.n8 12.8005
R2052 VTAIL.n44 VTAIL.n43 12.8005
R2053 VTAIL.n150 VTAIL.n149 12.8005
R2054 VTAIL.n146 VTAIL.n145 12.8005
R2055 VTAIL.n98 VTAIL.n97 12.8005
R2056 VTAIL.n94 VTAIL.n93 12.8005
R2057 VTAIL.n191 VTAIL.n190 12.0247
R2058 VTAIL.n203 VTAIL.n160 12.0247
R2059 VTAIL.n35 VTAIL.n34 12.0247
R2060 VTAIL.n47 VTAIL.n4 12.0247
R2061 VTAIL.n153 VTAIL.n110 12.0247
R2062 VTAIL.n142 VTAIL.n115 12.0247
R2063 VTAIL.n101 VTAIL.n58 12.0247
R2064 VTAIL.n90 VTAIL.n63 12.0247
R2065 VTAIL.n189 VTAIL.n166 11.249
R2066 VTAIL.n204 VTAIL.n158 11.249
R2067 VTAIL.n33 VTAIL.n10 11.249
R2068 VTAIL.n48 VTAIL.n2 11.249
R2069 VTAIL.n154 VTAIL.n108 11.249
R2070 VTAIL.n141 VTAIL.n118 11.249
R2071 VTAIL.n102 VTAIL.n56 11.249
R2072 VTAIL.n89 VTAIL.n66 11.249
R2073 VTAIL.n186 VTAIL.n185 10.4732
R2074 VTAIL.n30 VTAIL.n29 10.4732
R2075 VTAIL.n138 VTAIL.n137 10.4732
R2076 VTAIL.n86 VTAIL.n85 10.4732
R2077 VTAIL.n174 VTAIL.n173 10.2747
R2078 VTAIL.n18 VTAIL.n17 10.2747
R2079 VTAIL.n126 VTAIL.n125 10.2747
R2080 VTAIL.n74 VTAIL.n73 10.2747
R2081 VTAIL.n182 VTAIL.n168 9.69747
R2082 VTAIL.n26 VTAIL.n12 9.69747
R2083 VTAIL.n134 VTAIL.n120 9.69747
R2084 VTAIL.n82 VTAIL.n68 9.69747
R2085 VTAIL.n206 VTAIL.n205 9.45567
R2086 VTAIL.n50 VTAIL.n49 9.45567
R2087 VTAIL.n156 VTAIL.n155 9.45567
R2088 VTAIL.n104 VTAIL.n103 9.45567
R2089 VTAIL.n205 VTAIL.n204 9.3005
R2090 VTAIL.n160 VTAIL.n159 9.3005
R2091 VTAIL.n199 VTAIL.n198 9.3005
R2092 VTAIL.n172 VTAIL.n171 9.3005
R2093 VTAIL.n179 VTAIL.n178 9.3005
R2094 VTAIL.n181 VTAIL.n180 9.3005
R2095 VTAIL.n168 VTAIL.n167 9.3005
R2096 VTAIL.n187 VTAIL.n186 9.3005
R2097 VTAIL.n189 VTAIL.n188 9.3005
R2098 VTAIL.n190 VTAIL.n163 9.3005
R2099 VTAIL.n197 VTAIL.n196 9.3005
R2100 VTAIL.n49 VTAIL.n48 9.3005
R2101 VTAIL.n4 VTAIL.n3 9.3005
R2102 VTAIL.n43 VTAIL.n42 9.3005
R2103 VTAIL.n16 VTAIL.n15 9.3005
R2104 VTAIL.n23 VTAIL.n22 9.3005
R2105 VTAIL.n25 VTAIL.n24 9.3005
R2106 VTAIL.n12 VTAIL.n11 9.3005
R2107 VTAIL.n31 VTAIL.n30 9.3005
R2108 VTAIL.n33 VTAIL.n32 9.3005
R2109 VTAIL.n34 VTAIL.n7 9.3005
R2110 VTAIL.n41 VTAIL.n40 9.3005
R2111 VTAIL.n124 VTAIL.n123 9.3005
R2112 VTAIL.n131 VTAIL.n130 9.3005
R2113 VTAIL.n133 VTAIL.n132 9.3005
R2114 VTAIL.n120 VTAIL.n119 9.3005
R2115 VTAIL.n139 VTAIL.n138 9.3005
R2116 VTAIL.n141 VTAIL.n140 9.3005
R2117 VTAIL.n115 VTAIL.n113 9.3005
R2118 VTAIL.n147 VTAIL.n146 9.3005
R2119 VTAIL.n155 VTAIL.n154 9.3005
R2120 VTAIL.n110 VTAIL.n109 9.3005
R2121 VTAIL.n149 VTAIL.n148 9.3005
R2122 VTAIL.n72 VTAIL.n71 9.3005
R2123 VTAIL.n79 VTAIL.n78 9.3005
R2124 VTAIL.n81 VTAIL.n80 9.3005
R2125 VTAIL.n68 VTAIL.n67 9.3005
R2126 VTAIL.n87 VTAIL.n86 9.3005
R2127 VTAIL.n89 VTAIL.n88 9.3005
R2128 VTAIL.n63 VTAIL.n61 9.3005
R2129 VTAIL.n95 VTAIL.n94 9.3005
R2130 VTAIL.n103 VTAIL.n102 9.3005
R2131 VTAIL.n58 VTAIL.n57 9.3005
R2132 VTAIL.n97 VTAIL.n96 9.3005
R2133 VTAIL.n181 VTAIL.n170 8.92171
R2134 VTAIL.n25 VTAIL.n14 8.92171
R2135 VTAIL.n133 VTAIL.n122 8.92171
R2136 VTAIL.n81 VTAIL.n70 8.92171
R2137 VTAIL.n178 VTAIL.n177 8.14595
R2138 VTAIL.n22 VTAIL.n21 8.14595
R2139 VTAIL.n130 VTAIL.n129 8.14595
R2140 VTAIL.n78 VTAIL.n77 8.14595
R2141 VTAIL.n174 VTAIL.n172 7.3702
R2142 VTAIL.n18 VTAIL.n16 7.3702
R2143 VTAIL.n126 VTAIL.n124 7.3702
R2144 VTAIL.n74 VTAIL.n72 7.3702
R2145 VTAIL.n177 VTAIL.n172 5.81868
R2146 VTAIL.n21 VTAIL.n16 5.81868
R2147 VTAIL.n129 VTAIL.n124 5.81868
R2148 VTAIL.n77 VTAIL.n72 5.81868
R2149 VTAIL.n178 VTAIL.n170 5.04292
R2150 VTAIL.n22 VTAIL.n14 5.04292
R2151 VTAIL.n130 VTAIL.n122 5.04292
R2152 VTAIL.n78 VTAIL.n70 5.04292
R2153 VTAIL.n182 VTAIL.n181 4.26717
R2154 VTAIL.n26 VTAIL.n25 4.26717
R2155 VTAIL.n134 VTAIL.n133 4.26717
R2156 VTAIL.n82 VTAIL.n81 4.26717
R2157 VTAIL.n105 VTAIL.n55 3.67291
R2158 VTAIL.n157 VTAIL.n107 3.67291
R2159 VTAIL.n53 VTAIL.n51 3.67291
R2160 VTAIL.n185 VTAIL.n168 3.49141
R2161 VTAIL.n29 VTAIL.n12 3.49141
R2162 VTAIL.n137 VTAIL.n120 3.49141
R2163 VTAIL.n85 VTAIL.n68 3.49141
R2164 VTAIL.n173 VTAIL.n171 2.84303
R2165 VTAIL.n17 VTAIL.n15 2.84303
R2166 VTAIL.n125 VTAIL.n123 2.84303
R2167 VTAIL.n73 VTAIL.n71 2.84303
R2168 VTAIL.n186 VTAIL.n166 2.71565
R2169 VTAIL.n206 VTAIL.n158 2.71565
R2170 VTAIL.n30 VTAIL.n10 2.71565
R2171 VTAIL.n50 VTAIL.n2 2.71565
R2172 VTAIL.n156 VTAIL.n108 2.71565
R2173 VTAIL.n138 VTAIL.n118 2.71565
R2174 VTAIL.n104 VTAIL.n56 2.71565
R2175 VTAIL.n86 VTAIL.n66 2.71565
R2176 VTAIL VTAIL.n207 2.69662
R2177 VTAIL.n107 VTAIL.n105 2.30653
R2178 VTAIL.n51 VTAIL.n1 2.30653
R2179 VTAIL.n0 VTAIL.t4 2.10913
R2180 VTAIL.n0 VTAIL.t8 2.10913
R2181 VTAIL.n52 VTAIL.t11 2.10913
R2182 VTAIL.n52 VTAIL.t9 2.10913
R2183 VTAIL.n106 VTAIL.t1 2.10913
R2184 VTAIL.n106 VTAIL.t10 2.10913
R2185 VTAIL.n54 VTAIL.t6 2.10913
R2186 VTAIL.n54 VTAIL.t7 2.10913
R2187 VTAIL.n191 VTAIL.n189 1.93989
R2188 VTAIL.n204 VTAIL.n203 1.93989
R2189 VTAIL.n35 VTAIL.n33 1.93989
R2190 VTAIL.n48 VTAIL.n47 1.93989
R2191 VTAIL.n154 VTAIL.n153 1.93989
R2192 VTAIL.n142 VTAIL.n141 1.93989
R2193 VTAIL.n102 VTAIL.n101 1.93989
R2194 VTAIL.n90 VTAIL.n89 1.93989
R2195 VTAIL.n190 VTAIL.n164 1.16414
R2196 VTAIL.n200 VTAIL.n160 1.16414
R2197 VTAIL.n34 VTAIL.n8 1.16414
R2198 VTAIL.n44 VTAIL.n4 1.16414
R2199 VTAIL.n150 VTAIL.n110 1.16414
R2200 VTAIL.n145 VTAIL.n115 1.16414
R2201 VTAIL.n98 VTAIL.n58 1.16414
R2202 VTAIL.n93 VTAIL.n63 1.16414
R2203 VTAIL VTAIL.n1 0.976793
R2204 VTAIL.n196 VTAIL.n195 0.388379
R2205 VTAIL.n199 VTAIL.n162 0.388379
R2206 VTAIL.n40 VTAIL.n39 0.388379
R2207 VTAIL.n43 VTAIL.n6 0.388379
R2208 VTAIL.n149 VTAIL.n112 0.388379
R2209 VTAIL.n146 VTAIL.n114 0.388379
R2210 VTAIL.n97 VTAIL.n60 0.388379
R2211 VTAIL.n94 VTAIL.n62 0.388379
R2212 VTAIL.n179 VTAIL.n171 0.155672
R2213 VTAIL.n180 VTAIL.n179 0.155672
R2214 VTAIL.n180 VTAIL.n167 0.155672
R2215 VTAIL.n187 VTAIL.n167 0.155672
R2216 VTAIL.n188 VTAIL.n187 0.155672
R2217 VTAIL.n188 VTAIL.n163 0.155672
R2218 VTAIL.n197 VTAIL.n163 0.155672
R2219 VTAIL.n198 VTAIL.n197 0.155672
R2220 VTAIL.n198 VTAIL.n159 0.155672
R2221 VTAIL.n205 VTAIL.n159 0.155672
R2222 VTAIL.n23 VTAIL.n15 0.155672
R2223 VTAIL.n24 VTAIL.n23 0.155672
R2224 VTAIL.n24 VTAIL.n11 0.155672
R2225 VTAIL.n31 VTAIL.n11 0.155672
R2226 VTAIL.n32 VTAIL.n31 0.155672
R2227 VTAIL.n32 VTAIL.n7 0.155672
R2228 VTAIL.n41 VTAIL.n7 0.155672
R2229 VTAIL.n42 VTAIL.n41 0.155672
R2230 VTAIL.n42 VTAIL.n3 0.155672
R2231 VTAIL.n49 VTAIL.n3 0.155672
R2232 VTAIL.n155 VTAIL.n109 0.155672
R2233 VTAIL.n148 VTAIL.n109 0.155672
R2234 VTAIL.n148 VTAIL.n147 0.155672
R2235 VTAIL.n147 VTAIL.n113 0.155672
R2236 VTAIL.n140 VTAIL.n113 0.155672
R2237 VTAIL.n140 VTAIL.n139 0.155672
R2238 VTAIL.n139 VTAIL.n119 0.155672
R2239 VTAIL.n132 VTAIL.n119 0.155672
R2240 VTAIL.n132 VTAIL.n131 0.155672
R2241 VTAIL.n131 VTAIL.n123 0.155672
R2242 VTAIL.n103 VTAIL.n57 0.155672
R2243 VTAIL.n96 VTAIL.n57 0.155672
R2244 VTAIL.n96 VTAIL.n95 0.155672
R2245 VTAIL.n95 VTAIL.n61 0.155672
R2246 VTAIL.n88 VTAIL.n61 0.155672
R2247 VTAIL.n88 VTAIL.n87 0.155672
R2248 VTAIL.n87 VTAIL.n67 0.155672
R2249 VTAIL.n80 VTAIL.n67 0.155672
R2250 VTAIL.n80 VTAIL.n79 0.155672
R2251 VTAIL.n79 VTAIL.n71 0.155672
R2252 VP.n18 VP.n17 161.3
R2253 VP.n19 VP.n14 161.3
R2254 VP.n21 VP.n20 161.3
R2255 VP.n22 VP.n13 161.3
R2256 VP.n24 VP.n23 161.3
R2257 VP.n25 VP.n12 161.3
R2258 VP.n27 VP.n26 161.3
R2259 VP.n28 VP.n11 161.3
R2260 VP.n30 VP.n29 161.3
R2261 VP.n61 VP.n60 161.3
R2262 VP.n59 VP.n1 161.3
R2263 VP.n58 VP.n57 161.3
R2264 VP.n56 VP.n2 161.3
R2265 VP.n55 VP.n54 161.3
R2266 VP.n53 VP.n3 161.3
R2267 VP.n52 VP.n51 161.3
R2268 VP.n50 VP.n4 161.3
R2269 VP.n49 VP.n48 161.3
R2270 VP.n46 VP.n5 161.3
R2271 VP.n45 VP.n44 161.3
R2272 VP.n43 VP.n6 161.3
R2273 VP.n42 VP.n41 161.3
R2274 VP.n40 VP.n7 161.3
R2275 VP.n39 VP.n38 161.3
R2276 VP.n37 VP.n8 161.3
R2277 VP.n36 VP.n35 161.3
R2278 VP.n34 VP.n9 161.3
R2279 VP.n15 VP.t3 89.7238
R2280 VP.n33 VP.n32 89.5781
R2281 VP.n62 VP.n0 89.5781
R2282 VP.n31 VP.n10 89.5781
R2283 VP.n16 VP.n15 62.9256
R2284 VP.n33 VP.t2 57.5829
R2285 VP.n47 VP.t4 57.5829
R2286 VP.n0 VP.t1 57.5829
R2287 VP.n10 VP.t5 57.5829
R2288 VP.n16 VP.t0 57.5829
R2289 VP.n41 VP.n40 52.1486
R2290 VP.n54 VP.n53 52.1486
R2291 VP.n23 VP.n22 52.1486
R2292 VP.n32 VP.n31 51.9615
R2293 VP.n40 VP.n39 28.8382
R2294 VP.n54 VP.n2 28.8382
R2295 VP.n23 VP.n12 28.8382
R2296 VP.n35 VP.n34 24.4675
R2297 VP.n35 VP.n8 24.4675
R2298 VP.n39 VP.n8 24.4675
R2299 VP.n41 VP.n6 24.4675
R2300 VP.n45 VP.n6 24.4675
R2301 VP.n46 VP.n45 24.4675
R2302 VP.n48 VP.n4 24.4675
R2303 VP.n52 VP.n4 24.4675
R2304 VP.n53 VP.n52 24.4675
R2305 VP.n58 VP.n2 24.4675
R2306 VP.n59 VP.n58 24.4675
R2307 VP.n60 VP.n59 24.4675
R2308 VP.n27 VP.n12 24.4675
R2309 VP.n28 VP.n27 24.4675
R2310 VP.n29 VP.n28 24.4675
R2311 VP.n17 VP.n14 24.4675
R2312 VP.n21 VP.n14 24.4675
R2313 VP.n22 VP.n21 24.4675
R2314 VP.n47 VP.n46 12.234
R2315 VP.n48 VP.n47 12.234
R2316 VP.n17 VP.n16 12.234
R2317 VP.n18 VP.n15 2.52277
R2318 VP.n34 VP.n33 0.48984
R2319 VP.n60 VP.n0 0.48984
R2320 VP.n29 VP.n10 0.48984
R2321 VP.n31 VP.n30 0.354971
R2322 VP.n32 VP.n9 0.354971
R2323 VP.n62 VP.n61 0.354971
R2324 VP VP.n62 0.26696
R2325 VP.n19 VP.n18 0.189894
R2326 VP.n20 VP.n19 0.189894
R2327 VP.n20 VP.n13 0.189894
R2328 VP.n24 VP.n13 0.189894
R2329 VP.n25 VP.n24 0.189894
R2330 VP.n26 VP.n25 0.189894
R2331 VP.n26 VP.n11 0.189894
R2332 VP.n30 VP.n11 0.189894
R2333 VP.n36 VP.n9 0.189894
R2334 VP.n37 VP.n36 0.189894
R2335 VP.n38 VP.n37 0.189894
R2336 VP.n38 VP.n7 0.189894
R2337 VP.n42 VP.n7 0.189894
R2338 VP.n43 VP.n42 0.189894
R2339 VP.n44 VP.n43 0.189894
R2340 VP.n44 VP.n5 0.189894
R2341 VP.n49 VP.n5 0.189894
R2342 VP.n50 VP.n49 0.189894
R2343 VP.n51 VP.n50 0.189894
R2344 VP.n51 VP.n3 0.189894
R2345 VP.n55 VP.n3 0.189894
R2346 VP.n56 VP.n55 0.189894
R2347 VP.n57 VP.n56 0.189894
R2348 VP.n57 VP.n1 0.189894
R2349 VP.n61 VP.n1 0.189894
R2350 VDD1.n44 VDD1.n0 289.615
R2351 VDD1.n93 VDD1.n49 289.615
R2352 VDD1.n45 VDD1.n44 185
R2353 VDD1.n43 VDD1.n42 185
R2354 VDD1.n4 VDD1.n3 185
R2355 VDD1.n8 VDD1.n6 185
R2356 VDD1.n37 VDD1.n36 185
R2357 VDD1.n35 VDD1.n34 185
R2358 VDD1.n10 VDD1.n9 185
R2359 VDD1.n29 VDD1.n28 185
R2360 VDD1.n27 VDD1.n26 185
R2361 VDD1.n14 VDD1.n13 185
R2362 VDD1.n21 VDD1.n20 185
R2363 VDD1.n19 VDD1.n18 185
R2364 VDD1.n66 VDD1.n65 185
R2365 VDD1.n68 VDD1.n67 185
R2366 VDD1.n61 VDD1.n60 185
R2367 VDD1.n74 VDD1.n73 185
R2368 VDD1.n76 VDD1.n75 185
R2369 VDD1.n57 VDD1.n56 185
R2370 VDD1.n83 VDD1.n82 185
R2371 VDD1.n84 VDD1.n55 185
R2372 VDD1.n86 VDD1.n85 185
R2373 VDD1.n53 VDD1.n52 185
R2374 VDD1.n92 VDD1.n91 185
R2375 VDD1.n94 VDD1.n93 185
R2376 VDD1.n17 VDD1.t2 149.524
R2377 VDD1.n64 VDD1.t3 149.524
R2378 VDD1.n44 VDD1.n43 104.615
R2379 VDD1.n43 VDD1.n3 104.615
R2380 VDD1.n8 VDD1.n3 104.615
R2381 VDD1.n36 VDD1.n8 104.615
R2382 VDD1.n36 VDD1.n35 104.615
R2383 VDD1.n35 VDD1.n9 104.615
R2384 VDD1.n28 VDD1.n9 104.615
R2385 VDD1.n28 VDD1.n27 104.615
R2386 VDD1.n27 VDD1.n13 104.615
R2387 VDD1.n20 VDD1.n13 104.615
R2388 VDD1.n20 VDD1.n19 104.615
R2389 VDD1.n67 VDD1.n66 104.615
R2390 VDD1.n67 VDD1.n60 104.615
R2391 VDD1.n74 VDD1.n60 104.615
R2392 VDD1.n75 VDD1.n74 104.615
R2393 VDD1.n75 VDD1.n56 104.615
R2394 VDD1.n83 VDD1.n56 104.615
R2395 VDD1.n84 VDD1.n83 104.615
R2396 VDD1.n85 VDD1.n84 104.615
R2397 VDD1.n85 VDD1.n52 104.615
R2398 VDD1.n92 VDD1.n52 104.615
R2399 VDD1.n93 VDD1.n92 104.615
R2400 VDD1.n99 VDD1.n98 66.7737
R2401 VDD1.n101 VDD1.n100 65.911
R2402 VDD1 VDD1.n48 54.5857
R2403 VDD1.n99 VDD1.n97 54.4722
R2404 VDD1.n19 VDD1.t2 52.3082
R2405 VDD1.n66 VDD1.t3 52.3082
R2406 VDD1.n101 VDD1.n99 46.1647
R2407 VDD1.n6 VDD1.n4 13.1884
R2408 VDD1.n86 VDD1.n53 13.1884
R2409 VDD1.n42 VDD1.n41 12.8005
R2410 VDD1.n38 VDD1.n37 12.8005
R2411 VDD1.n87 VDD1.n55 12.8005
R2412 VDD1.n91 VDD1.n90 12.8005
R2413 VDD1.n45 VDD1.n2 12.0247
R2414 VDD1.n34 VDD1.n7 12.0247
R2415 VDD1.n82 VDD1.n81 12.0247
R2416 VDD1.n94 VDD1.n51 12.0247
R2417 VDD1.n46 VDD1.n0 11.249
R2418 VDD1.n33 VDD1.n10 11.249
R2419 VDD1.n80 VDD1.n57 11.249
R2420 VDD1.n95 VDD1.n49 11.249
R2421 VDD1.n30 VDD1.n29 10.4732
R2422 VDD1.n77 VDD1.n76 10.4732
R2423 VDD1.n18 VDD1.n17 10.2747
R2424 VDD1.n65 VDD1.n64 10.2747
R2425 VDD1.n26 VDD1.n12 9.69747
R2426 VDD1.n73 VDD1.n59 9.69747
R2427 VDD1.n48 VDD1.n47 9.45567
R2428 VDD1.n97 VDD1.n96 9.45567
R2429 VDD1.n16 VDD1.n15 9.3005
R2430 VDD1.n23 VDD1.n22 9.3005
R2431 VDD1.n25 VDD1.n24 9.3005
R2432 VDD1.n12 VDD1.n11 9.3005
R2433 VDD1.n31 VDD1.n30 9.3005
R2434 VDD1.n33 VDD1.n32 9.3005
R2435 VDD1.n7 VDD1.n5 9.3005
R2436 VDD1.n39 VDD1.n38 9.3005
R2437 VDD1.n47 VDD1.n46 9.3005
R2438 VDD1.n2 VDD1.n1 9.3005
R2439 VDD1.n41 VDD1.n40 9.3005
R2440 VDD1.n96 VDD1.n95 9.3005
R2441 VDD1.n51 VDD1.n50 9.3005
R2442 VDD1.n90 VDD1.n89 9.3005
R2443 VDD1.n63 VDD1.n62 9.3005
R2444 VDD1.n70 VDD1.n69 9.3005
R2445 VDD1.n72 VDD1.n71 9.3005
R2446 VDD1.n59 VDD1.n58 9.3005
R2447 VDD1.n78 VDD1.n77 9.3005
R2448 VDD1.n80 VDD1.n79 9.3005
R2449 VDD1.n81 VDD1.n54 9.3005
R2450 VDD1.n88 VDD1.n87 9.3005
R2451 VDD1.n25 VDD1.n14 8.92171
R2452 VDD1.n72 VDD1.n61 8.92171
R2453 VDD1.n22 VDD1.n21 8.14595
R2454 VDD1.n69 VDD1.n68 8.14595
R2455 VDD1.n18 VDD1.n16 7.3702
R2456 VDD1.n65 VDD1.n63 7.3702
R2457 VDD1.n21 VDD1.n16 5.81868
R2458 VDD1.n68 VDD1.n63 5.81868
R2459 VDD1.n22 VDD1.n14 5.04292
R2460 VDD1.n69 VDD1.n61 5.04292
R2461 VDD1.n26 VDD1.n25 4.26717
R2462 VDD1.n73 VDD1.n72 4.26717
R2463 VDD1.n29 VDD1.n12 3.49141
R2464 VDD1.n76 VDD1.n59 3.49141
R2465 VDD1.n17 VDD1.n15 2.84303
R2466 VDD1.n64 VDD1.n62 2.84303
R2467 VDD1.n48 VDD1.n0 2.71565
R2468 VDD1.n30 VDD1.n10 2.71565
R2469 VDD1.n77 VDD1.n57 2.71565
R2470 VDD1.n97 VDD1.n49 2.71565
R2471 VDD1.n100 VDD1.t5 2.10913
R2472 VDD1.n100 VDD1.t0 2.10913
R2473 VDD1.n98 VDD1.t1 2.10913
R2474 VDD1.n98 VDD1.t4 2.10913
R2475 VDD1.n46 VDD1.n45 1.93989
R2476 VDD1.n34 VDD1.n33 1.93989
R2477 VDD1.n82 VDD1.n80 1.93989
R2478 VDD1.n95 VDD1.n94 1.93989
R2479 VDD1.n42 VDD1.n2 1.16414
R2480 VDD1.n37 VDD1.n7 1.16414
R2481 VDD1.n81 VDD1.n55 1.16414
R2482 VDD1.n91 VDD1.n51 1.16414
R2483 VDD1 VDD1.n101 0.860414
R2484 VDD1.n41 VDD1.n4 0.388379
R2485 VDD1.n38 VDD1.n6 0.388379
R2486 VDD1.n87 VDD1.n86 0.388379
R2487 VDD1.n90 VDD1.n53 0.388379
R2488 VDD1.n47 VDD1.n1 0.155672
R2489 VDD1.n40 VDD1.n1 0.155672
R2490 VDD1.n40 VDD1.n39 0.155672
R2491 VDD1.n39 VDD1.n5 0.155672
R2492 VDD1.n32 VDD1.n5 0.155672
R2493 VDD1.n32 VDD1.n31 0.155672
R2494 VDD1.n31 VDD1.n11 0.155672
R2495 VDD1.n24 VDD1.n11 0.155672
R2496 VDD1.n24 VDD1.n23 0.155672
R2497 VDD1.n23 VDD1.n15 0.155672
R2498 VDD1.n70 VDD1.n62 0.155672
R2499 VDD1.n71 VDD1.n70 0.155672
R2500 VDD1.n71 VDD1.n58 0.155672
R2501 VDD1.n78 VDD1.n58 0.155672
R2502 VDD1.n79 VDD1.n78 0.155672
R2503 VDD1.n79 VDD1.n54 0.155672
R2504 VDD1.n88 VDD1.n54 0.155672
R2505 VDD1.n89 VDD1.n88 0.155672
R2506 VDD1.n89 VDD1.n50 0.155672
R2507 VDD1.n96 VDD1.n50 0.155672
C0 VTAIL VDD1 7.40626f
C1 VDD2 VP 0.570469f
C2 VP VN 7.73644f
C3 VDD2 VN 5.70488f
C4 VTAIL VP 6.32585f
C5 VDD1 VP 6.12058f
C6 VTAIL VDD2 7.46744f
C7 VTAIL VN 6.31113f
C8 VDD1 VDD2 1.92596f
C9 VDD1 VN 0.15257f
C10 VDD2 B 6.542317f
C11 VDD1 B 6.738877f
C12 VTAIL B 7.587101f
C13 VN B 16.617708f
C14 VP B 15.359194f
C15 VDD1.n0 B 0.030686f
C16 VDD1.n1 B 0.021937f
C17 VDD1.n2 B 0.011788f
C18 VDD1.n3 B 0.027862f
C19 VDD1.n4 B 0.012134f
C20 VDD1.n5 B 0.021937f
C21 VDD1.n6 B 0.012134f
C22 VDD1.n7 B 0.011788f
C23 VDD1.n8 B 0.027862f
C24 VDD1.n9 B 0.027862f
C25 VDD1.n10 B 0.012481f
C26 VDD1.n11 B 0.021937f
C27 VDD1.n12 B 0.011788f
C28 VDD1.n13 B 0.027862f
C29 VDD1.n14 B 0.012481f
C30 VDD1.n15 B 0.851993f
C31 VDD1.n16 B 0.011788f
C32 VDD1.t2 B 0.046753f
C33 VDD1.n17 B 0.136187f
C34 VDD1.n18 B 0.019696f
C35 VDD1.n19 B 0.020896f
C36 VDD1.n20 B 0.027862f
C37 VDD1.n21 B 0.012481f
C38 VDD1.n22 B 0.011788f
C39 VDD1.n23 B 0.021937f
C40 VDD1.n24 B 0.021937f
C41 VDD1.n25 B 0.011788f
C42 VDD1.n26 B 0.012481f
C43 VDD1.n27 B 0.027862f
C44 VDD1.n28 B 0.027862f
C45 VDD1.n29 B 0.012481f
C46 VDD1.n30 B 0.011788f
C47 VDD1.n31 B 0.021937f
C48 VDD1.n32 B 0.021937f
C49 VDD1.n33 B 0.011788f
C50 VDD1.n34 B 0.012481f
C51 VDD1.n35 B 0.027862f
C52 VDD1.n36 B 0.027862f
C53 VDD1.n37 B 0.012481f
C54 VDD1.n38 B 0.011788f
C55 VDD1.n39 B 0.021937f
C56 VDD1.n40 B 0.021937f
C57 VDD1.n41 B 0.011788f
C58 VDD1.n42 B 0.012481f
C59 VDD1.n43 B 0.027862f
C60 VDD1.n44 B 0.060055f
C61 VDD1.n45 B 0.012481f
C62 VDD1.n46 B 0.011788f
C63 VDD1.n47 B 0.055201f
C64 VDD1.n48 B 0.061376f
C65 VDD1.n49 B 0.030686f
C66 VDD1.n50 B 0.021937f
C67 VDD1.n51 B 0.011788f
C68 VDD1.n52 B 0.027862f
C69 VDD1.n53 B 0.012134f
C70 VDD1.n54 B 0.021937f
C71 VDD1.n55 B 0.012481f
C72 VDD1.n56 B 0.027862f
C73 VDD1.n57 B 0.012481f
C74 VDD1.n58 B 0.021937f
C75 VDD1.n59 B 0.011788f
C76 VDD1.n60 B 0.027862f
C77 VDD1.n61 B 0.012481f
C78 VDD1.n62 B 0.851993f
C79 VDD1.n63 B 0.011788f
C80 VDD1.t3 B 0.046753f
C81 VDD1.n64 B 0.136187f
C82 VDD1.n65 B 0.019696f
C83 VDD1.n66 B 0.020896f
C84 VDD1.n67 B 0.027862f
C85 VDD1.n68 B 0.012481f
C86 VDD1.n69 B 0.011788f
C87 VDD1.n70 B 0.021937f
C88 VDD1.n71 B 0.021937f
C89 VDD1.n72 B 0.011788f
C90 VDD1.n73 B 0.012481f
C91 VDD1.n74 B 0.027862f
C92 VDD1.n75 B 0.027862f
C93 VDD1.n76 B 0.012481f
C94 VDD1.n77 B 0.011788f
C95 VDD1.n78 B 0.021937f
C96 VDD1.n79 B 0.021937f
C97 VDD1.n80 B 0.011788f
C98 VDD1.n81 B 0.011788f
C99 VDD1.n82 B 0.012481f
C100 VDD1.n83 B 0.027862f
C101 VDD1.n84 B 0.027862f
C102 VDD1.n85 B 0.027862f
C103 VDD1.n86 B 0.012134f
C104 VDD1.n87 B 0.011788f
C105 VDD1.n88 B 0.021937f
C106 VDD1.n89 B 0.021937f
C107 VDD1.n90 B 0.011788f
C108 VDD1.n91 B 0.012481f
C109 VDD1.n92 B 0.027862f
C110 VDD1.n93 B 0.060055f
C111 VDD1.n94 B 0.012481f
C112 VDD1.n95 B 0.011788f
C113 VDD1.n96 B 0.055201f
C114 VDD1.n97 B 0.060506f
C115 VDD1.t1 B 0.162775f
C116 VDD1.t4 B 0.162775f
C117 VDD1.n98 B 1.43521f
C118 VDD1.n99 B 2.84757f
C119 VDD1.t5 B 0.162775f
C120 VDD1.t0 B 0.162775f
C121 VDD1.n100 B 1.42867f
C122 VDD1.n101 B 2.59736f
C123 VP.t1 B 1.89886f
C124 VP.n0 B 0.745123f
C125 VP.n1 B 0.019037f
C126 VP.n2 B 0.037656f
C127 VP.n3 B 0.019037f
C128 VP.n4 B 0.03548f
C129 VP.n5 B 0.019037f
C130 VP.t4 B 1.89886f
C131 VP.n6 B 0.03548f
C132 VP.n7 B 0.019037f
C133 VP.n8 B 0.03548f
C134 VP.n9 B 0.030725f
C135 VP.t2 B 1.89886f
C136 VP.t5 B 1.89886f
C137 VP.n10 B 0.745123f
C138 VP.n11 B 0.019037f
C139 VP.n12 B 0.037656f
C140 VP.n13 B 0.019037f
C141 VP.n14 B 0.03548f
C142 VP.t3 B 2.19538f
C143 VP.n15 B 0.711797f
C144 VP.t0 B 1.89886f
C145 VP.n16 B 0.743001f
C146 VP.n17 B 0.026721f
C147 VP.n18 B 0.248849f
C148 VP.n19 B 0.019037f
C149 VP.n20 B 0.019037f
C150 VP.n21 B 0.03548f
C151 VP.n22 B 0.034176f
C152 VP.n23 B 0.019228f
C153 VP.n24 B 0.019037f
C154 VP.n25 B 0.019037f
C155 VP.n26 B 0.019037f
C156 VP.n27 B 0.03548f
C157 VP.n28 B 0.03548f
C158 VP.n29 B 0.018313f
C159 VP.n30 B 0.030725f
C160 VP.n31 B 1.15954f
C161 VP.n32 B 1.17271f
C162 VP.n33 B 0.745123f
C163 VP.n34 B 0.018313f
C164 VP.n35 B 0.03548f
C165 VP.n36 B 0.019037f
C166 VP.n37 B 0.019037f
C167 VP.n38 B 0.019037f
C168 VP.n39 B 0.037656f
C169 VP.n40 B 0.019228f
C170 VP.n41 B 0.034176f
C171 VP.n42 B 0.019037f
C172 VP.n43 B 0.019037f
C173 VP.n44 B 0.019037f
C174 VP.n45 B 0.03548f
C175 VP.n46 B 0.026721f
C176 VP.n47 B 0.673767f
C177 VP.n48 B 0.026721f
C178 VP.n49 B 0.019037f
C179 VP.n50 B 0.019037f
C180 VP.n51 B 0.019037f
C181 VP.n52 B 0.03548f
C182 VP.n53 B 0.034176f
C183 VP.n54 B 0.019228f
C184 VP.n55 B 0.019037f
C185 VP.n56 B 0.019037f
C186 VP.n57 B 0.019037f
C187 VP.n58 B 0.03548f
C188 VP.n59 B 0.03548f
C189 VP.n60 B 0.018313f
C190 VP.n61 B 0.030725f
C191 VP.n62 B 0.061207f
C192 VTAIL.t4 B 0.190941f
C193 VTAIL.t8 B 0.190941f
C194 VTAIL.n0 B 1.60761f
C195 VTAIL.n1 B 0.511889f
C196 VTAIL.n2 B 0.035996f
C197 VTAIL.n3 B 0.025732f
C198 VTAIL.n4 B 0.013827f
C199 VTAIL.n5 B 0.032683f
C200 VTAIL.n6 B 0.014234f
C201 VTAIL.n7 B 0.025732f
C202 VTAIL.n8 B 0.014641f
C203 VTAIL.n9 B 0.032683f
C204 VTAIL.n10 B 0.014641f
C205 VTAIL.n11 B 0.025732f
C206 VTAIL.n12 B 0.013827f
C207 VTAIL.n13 B 0.032683f
C208 VTAIL.n14 B 0.014641f
C209 VTAIL.n15 B 0.999418f
C210 VTAIL.n16 B 0.013827f
C211 VTAIL.t2 B 0.054843f
C212 VTAIL.n17 B 0.159752f
C213 VTAIL.n18 B 0.023105f
C214 VTAIL.n19 B 0.024512f
C215 VTAIL.n20 B 0.032683f
C216 VTAIL.n21 B 0.014641f
C217 VTAIL.n22 B 0.013827f
C218 VTAIL.n23 B 0.025732f
C219 VTAIL.n24 B 0.025732f
C220 VTAIL.n25 B 0.013827f
C221 VTAIL.n26 B 0.014641f
C222 VTAIL.n27 B 0.032683f
C223 VTAIL.n28 B 0.032683f
C224 VTAIL.n29 B 0.014641f
C225 VTAIL.n30 B 0.013827f
C226 VTAIL.n31 B 0.025732f
C227 VTAIL.n32 B 0.025732f
C228 VTAIL.n33 B 0.013827f
C229 VTAIL.n34 B 0.013827f
C230 VTAIL.n35 B 0.014641f
C231 VTAIL.n36 B 0.032683f
C232 VTAIL.n37 B 0.032683f
C233 VTAIL.n38 B 0.032683f
C234 VTAIL.n39 B 0.014234f
C235 VTAIL.n40 B 0.013827f
C236 VTAIL.n41 B 0.025732f
C237 VTAIL.n42 B 0.025732f
C238 VTAIL.n43 B 0.013827f
C239 VTAIL.n44 B 0.014641f
C240 VTAIL.n45 B 0.032683f
C241 VTAIL.n46 B 0.070446f
C242 VTAIL.n47 B 0.014641f
C243 VTAIL.n48 B 0.013827f
C244 VTAIL.n49 B 0.064752f
C245 VTAIL.n50 B 0.039542f
C246 VTAIL.n51 B 0.520667f
C247 VTAIL.t11 B 0.190941f
C248 VTAIL.t9 B 0.190941f
C249 VTAIL.n52 B 1.60761f
C250 VTAIL.n53 B 2.17397f
C251 VTAIL.t6 B 0.190941f
C252 VTAIL.t7 B 0.190941f
C253 VTAIL.n54 B 1.60762f
C254 VTAIL.n55 B 2.17396f
C255 VTAIL.n56 B 0.035996f
C256 VTAIL.n57 B 0.025732f
C257 VTAIL.n58 B 0.013827f
C258 VTAIL.n59 B 0.032683f
C259 VTAIL.n60 B 0.014234f
C260 VTAIL.n61 B 0.025732f
C261 VTAIL.n62 B 0.014234f
C262 VTAIL.n63 B 0.013827f
C263 VTAIL.n64 B 0.032683f
C264 VTAIL.n65 B 0.032683f
C265 VTAIL.n66 B 0.014641f
C266 VTAIL.n67 B 0.025732f
C267 VTAIL.n68 B 0.013827f
C268 VTAIL.n69 B 0.032683f
C269 VTAIL.n70 B 0.014641f
C270 VTAIL.n71 B 0.999418f
C271 VTAIL.n72 B 0.013827f
C272 VTAIL.t3 B 0.054843f
C273 VTAIL.n73 B 0.159752f
C274 VTAIL.n74 B 0.023105f
C275 VTAIL.n75 B 0.024512f
C276 VTAIL.n76 B 0.032683f
C277 VTAIL.n77 B 0.014641f
C278 VTAIL.n78 B 0.013827f
C279 VTAIL.n79 B 0.025732f
C280 VTAIL.n80 B 0.025732f
C281 VTAIL.n81 B 0.013827f
C282 VTAIL.n82 B 0.014641f
C283 VTAIL.n83 B 0.032683f
C284 VTAIL.n84 B 0.032683f
C285 VTAIL.n85 B 0.014641f
C286 VTAIL.n86 B 0.013827f
C287 VTAIL.n87 B 0.025732f
C288 VTAIL.n88 B 0.025732f
C289 VTAIL.n89 B 0.013827f
C290 VTAIL.n90 B 0.014641f
C291 VTAIL.n91 B 0.032683f
C292 VTAIL.n92 B 0.032683f
C293 VTAIL.n93 B 0.014641f
C294 VTAIL.n94 B 0.013827f
C295 VTAIL.n95 B 0.025732f
C296 VTAIL.n96 B 0.025732f
C297 VTAIL.n97 B 0.013827f
C298 VTAIL.n98 B 0.014641f
C299 VTAIL.n99 B 0.032683f
C300 VTAIL.n100 B 0.070446f
C301 VTAIL.n101 B 0.014641f
C302 VTAIL.n102 B 0.013827f
C303 VTAIL.n103 B 0.064752f
C304 VTAIL.n104 B 0.039542f
C305 VTAIL.n105 B 0.520667f
C306 VTAIL.t1 B 0.190941f
C307 VTAIL.t10 B 0.190941f
C308 VTAIL.n106 B 1.60762f
C309 VTAIL.n107 B 0.73543f
C310 VTAIL.n108 B 0.035996f
C311 VTAIL.n109 B 0.025732f
C312 VTAIL.n110 B 0.013827f
C313 VTAIL.n111 B 0.032683f
C314 VTAIL.n112 B 0.014234f
C315 VTAIL.n113 B 0.025732f
C316 VTAIL.n114 B 0.014234f
C317 VTAIL.n115 B 0.013827f
C318 VTAIL.n116 B 0.032683f
C319 VTAIL.n117 B 0.032683f
C320 VTAIL.n118 B 0.014641f
C321 VTAIL.n119 B 0.025732f
C322 VTAIL.n120 B 0.013827f
C323 VTAIL.n121 B 0.032683f
C324 VTAIL.n122 B 0.014641f
C325 VTAIL.n123 B 0.999418f
C326 VTAIL.n124 B 0.013827f
C327 VTAIL.t0 B 0.054843f
C328 VTAIL.n125 B 0.159752f
C329 VTAIL.n126 B 0.023105f
C330 VTAIL.n127 B 0.024512f
C331 VTAIL.n128 B 0.032683f
C332 VTAIL.n129 B 0.014641f
C333 VTAIL.n130 B 0.013827f
C334 VTAIL.n131 B 0.025732f
C335 VTAIL.n132 B 0.025732f
C336 VTAIL.n133 B 0.013827f
C337 VTAIL.n134 B 0.014641f
C338 VTAIL.n135 B 0.032683f
C339 VTAIL.n136 B 0.032683f
C340 VTAIL.n137 B 0.014641f
C341 VTAIL.n138 B 0.013827f
C342 VTAIL.n139 B 0.025732f
C343 VTAIL.n140 B 0.025732f
C344 VTAIL.n141 B 0.013827f
C345 VTAIL.n142 B 0.014641f
C346 VTAIL.n143 B 0.032683f
C347 VTAIL.n144 B 0.032683f
C348 VTAIL.n145 B 0.014641f
C349 VTAIL.n146 B 0.013827f
C350 VTAIL.n147 B 0.025732f
C351 VTAIL.n148 B 0.025732f
C352 VTAIL.n149 B 0.013827f
C353 VTAIL.n150 B 0.014641f
C354 VTAIL.n151 B 0.032683f
C355 VTAIL.n152 B 0.070446f
C356 VTAIL.n153 B 0.014641f
C357 VTAIL.n154 B 0.013827f
C358 VTAIL.n155 B 0.064752f
C359 VTAIL.n156 B 0.039542f
C360 VTAIL.n157 B 1.65469f
C361 VTAIL.n158 B 0.035996f
C362 VTAIL.n159 B 0.025732f
C363 VTAIL.n160 B 0.013827f
C364 VTAIL.n161 B 0.032683f
C365 VTAIL.n162 B 0.014234f
C366 VTAIL.n163 B 0.025732f
C367 VTAIL.n164 B 0.014641f
C368 VTAIL.n165 B 0.032683f
C369 VTAIL.n166 B 0.014641f
C370 VTAIL.n167 B 0.025732f
C371 VTAIL.n168 B 0.013827f
C372 VTAIL.n169 B 0.032683f
C373 VTAIL.n170 B 0.014641f
C374 VTAIL.n171 B 0.999418f
C375 VTAIL.n172 B 0.013827f
C376 VTAIL.t5 B 0.054843f
C377 VTAIL.n173 B 0.159752f
C378 VTAIL.n174 B 0.023105f
C379 VTAIL.n175 B 0.024512f
C380 VTAIL.n176 B 0.032683f
C381 VTAIL.n177 B 0.014641f
C382 VTAIL.n178 B 0.013827f
C383 VTAIL.n179 B 0.025732f
C384 VTAIL.n180 B 0.025732f
C385 VTAIL.n181 B 0.013827f
C386 VTAIL.n182 B 0.014641f
C387 VTAIL.n183 B 0.032683f
C388 VTAIL.n184 B 0.032683f
C389 VTAIL.n185 B 0.014641f
C390 VTAIL.n186 B 0.013827f
C391 VTAIL.n187 B 0.025732f
C392 VTAIL.n188 B 0.025732f
C393 VTAIL.n189 B 0.013827f
C394 VTAIL.n190 B 0.013827f
C395 VTAIL.n191 B 0.014641f
C396 VTAIL.n192 B 0.032683f
C397 VTAIL.n193 B 0.032683f
C398 VTAIL.n194 B 0.032683f
C399 VTAIL.n195 B 0.014234f
C400 VTAIL.n196 B 0.013827f
C401 VTAIL.n197 B 0.025732f
C402 VTAIL.n198 B 0.025732f
C403 VTAIL.n199 B 0.013827f
C404 VTAIL.n200 B 0.014641f
C405 VTAIL.n201 B 0.032683f
C406 VTAIL.n202 B 0.070446f
C407 VTAIL.n203 B 0.014641f
C408 VTAIL.n204 B 0.013827f
C409 VTAIL.n205 B 0.064752f
C410 VTAIL.n206 B 0.039542f
C411 VTAIL.n207 B 1.57374f
C412 VDD2.n0 B 0.030185f
C413 VDD2.n1 B 0.021579f
C414 VDD2.n2 B 0.011595f
C415 VDD2.n3 B 0.027407f
C416 VDD2.n4 B 0.011936f
C417 VDD2.n5 B 0.021579f
C418 VDD2.n6 B 0.012277f
C419 VDD2.n7 B 0.027407f
C420 VDD2.n8 B 0.012277f
C421 VDD2.n9 B 0.021579f
C422 VDD2.n10 B 0.011595f
C423 VDD2.n11 B 0.027407f
C424 VDD2.n12 B 0.012277f
C425 VDD2.n13 B 0.838089f
C426 VDD2.n14 B 0.011595f
C427 VDD2.t4 B 0.04599f
C428 VDD2.n15 B 0.133964f
C429 VDD2.n16 B 0.019375f
C430 VDD2.n17 B 0.020555f
C431 VDD2.n18 B 0.027407f
C432 VDD2.n19 B 0.012277f
C433 VDD2.n20 B 0.011595f
C434 VDD2.n21 B 0.021579f
C435 VDD2.n22 B 0.021579f
C436 VDD2.n23 B 0.011595f
C437 VDD2.n24 B 0.012277f
C438 VDD2.n25 B 0.027407f
C439 VDD2.n26 B 0.027407f
C440 VDD2.n27 B 0.012277f
C441 VDD2.n28 B 0.011595f
C442 VDD2.n29 B 0.021579f
C443 VDD2.n30 B 0.021579f
C444 VDD2.n31 B 0.011595f
C445 VDD2.n32 B 0.011595f
C446 VDD2.n33 B 0.012277f
C447 VDD2.n34 B 0.027407f
C448 VDD2.n35 B 0.027407f
C449 VDD2.n36 B 0.027407f
C450 VDD2.n37 B 0.011936f
C451 VDD2.n38 B 0.011595f
C452 VDD2.n39 B 0.021579f
C453 VDD2.n40 B 0.021579f
C454 VDD2.n41 B 0.011595f
C455 VDD2.n42 B 0.012277f
C456 VDD2.n43 B 0.027407f
C457 VDD2.n44 B 0.059075f
C458 VDD2.n45 B 0.012277f
C459 VDD2.n46 B 0.011595f
C460 VDD2.n47 B 0.0543f
C461 VDD2.n48 B 0.059519f
C462 VDD2.t0 B 0.160119f
C463 VDD2.t3 B 0.160119f
C464 VDD2.n49 B 1.41179f
C465 VDD2.n50 B 2.66553f
C466 VDD2.n51 B 0.030185f
C467 VDD2.n52 B 0.021579f
C468 VDD2.n53 B 0.011595f
C469 VDD2.n54 B 0.027407f
C470 VDD2.n55 B 0.011936f
C471 VDD2.n56 B 0.021579f
C472 VDD2.n57 B 0.011936f
C473 VDD2.n58 B 0.011595f
C474 VDD2.n59 B 0.027407f
C475 VDD2.n60 B 0.027407f
C476 VDD2.n61 B 0.012277f
C477 VDD2.n62 B 0.021579f
C478 VDD2.n63 B 0.011595f
C479 VDD2.n64 B 0.027407f
C480 VDD2.n65 B 0.012277f
C481 VDD2.n66 B 0.838089f
C482 VDD2.n67 B 0.011595f
C483 VDD2.t2 B 0.04599f
C484 VDD2.n68 B 0.133964f
C485 VDD2.n69 B 0.019375f
C486 VDD2.n70 B 0.020555f
C487 VDD2.n71 B 0.027407f
C488 VDD2.n72 B 0.012277f
C489 VDD2.n73 B 0.011595f
C490 VDD2.n74 B 0.021579f
C491 VDD2.n75 B 0.021579f
C492 VDD2.n76 B 0.011595f
C493 VDD2.n77 B 0.012277f
C494 VDD2.n78 B 0.027407f
C495 VDD2.n79 B 0.027407f
C496 VDD2.n80 B 0.012277f
C497 VDD2.n81 B 0.011595f
C498 VDD2.n82 B 0.021579f
C499 VDD2.n83 B 0.021579f
C500 VDD2.n84 B 0.011595f
C501 VDD2.n85 B 0.012277f
C502 VDD2.n86 B 0.027407f
C503 VDD2.n87 B 0.027407f
C504 VDD2.n88 B 0.012277f
C505 VDD2.n89 B 0.011595f
C506 VDD2.n90 B 0.021579f
C507 VDD2.n91 B 0.021579f
C508 VDD2.n92 B 0.011595f
C509 VDD2.n93 B 0.012277f
C510 VDD2.n94 B 0.027407f
C511 VDD2.n95 B 0.059075f
C512 VDD2.n96 B 0.012277f
C513 VDD2.n97 B 0.011595f
C514 VDD2.n98 B 0.0543f
C515 VDD2.n99 B 0.048027f
C516 VDD2.n100 B 2.35355f
C517 VDD2.t1 B 0.160119f
C518 VDD2.t5 B 0.160119f
C519 VDD2.n101 B 1.41176f
C520 VN.t3 B 1.8586f
C521 VN.n0 B 0.729324f
C522 VN.n1 B 0.018633f
C523 VN.n2 B 0.036857f
C524 VN.n3 B 0.018633f
C525 VN.n4 B 0.034727f
C526 VN.t4 B 2.14883f
C527 VN.n5 B 0.696704f
C528 VN.t0 B 1.8586f
C529 VN.n6 B 0.727247f
C530 VN.n7 B 0.026155f
C531 VN.n8 B 0.243572f
C532 VN.n9 B 0.018633f
C533 VN.n10 B 0.018633f
C534 VN.n11 B 0.034727f
C535 VN.n12 B 0.033452f
C536 VN.n13 B 0.018821f
C537 VN.n14 B 0.018633f
C538 VN.n15 B 0.018633f
C539 VN.n16 B 0.018633f
C540 VN.n17 B 0.034727f
C541 VN.n18 B 0.034727f
C542 VN.n19 B 0.017925f
C543 VN.n20 B 0.030073f
C544 VN.n21 B 0.05991f
C545 VN.t2 B 1.8586f
C546 VN.n22 B 0.729324f
C547 VN.n23 B 0.018633f
C548 VN.n24 B 0.036857f
C549 VN.n25 B 0.018633f
C550 VN.n26 B 0.034727f
C551 VN.t5 B 2.14883f
C552 VN.n27 B 0.696704f
C553 VN.t1 B 1.8586f
C554 VN.n28 B 0.727247f
C555 VN.n29 B 0.026155f
C556 VN.n30 B 0.243572f
C557 VN.n31 B 0.018633f
C558 VN.n32 B 0.018633f
C559 VN.n33 B 0.034727f
C560 VN.n34 B 0.033452f
C561 VN.n35 B 0.018821f
C562 VN.n36 B 0.018633f
C563 VN.n37 B 0.018633f
C564 VN.n38 B 0.018633f
C565 VN.n39 B 0.034727f
C566 VN.n40 B 0.034727f
C567 VN.n41 B 0.017925f
C568 VN.n42 B 0.030073f
C569 VN.n43 B 1.14248f
.ends

