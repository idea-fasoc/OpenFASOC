* NGSPICE file created from diff_pair_sample_1581.ext - technology: sky130A

.subckt diff_pair_sample_1581 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=1.17
X1 VTAIL.t7 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X2 VDD1.t6 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X3 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=1.17
X4 VTAIL.t14 VN.t1 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X5 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=1.17
X6 VTAIL.t2 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X7 VDD2.t0 VN.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=1.17
X9 VTAIL.t4 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=1.17
X10 VDD2.t2 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=1.17
X11 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=1.17
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=1.17
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=0 ps=0 w=8.36 l=1.17
X14 VTAIL.t11 VN.t4 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X15 VTAIL.t10 VN.t5 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=1.17
X16 VDD2.t4 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X17 VTAIL.t6 VP.t6 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2604 pd=17.5 as=1.3794 ps=8.69 w=8.36 l=1.17
X18 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=1.3794 ps=8.69 w=8.36 l=1.17
X19 VDD2.t7 VN.t7 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3794 pd=8.69 as=3.2604 ps=17.5 w=8.36 l=1.17
R0 VN.n4 VN.t5 202.382
R1 VN.n22 VN.t3 202.382
R2 VN.n16 VN.n15 173.596
R3 VN.n33 VN.n32 173.596
R4 VN.n3 VN.t2 172.202
R5 VN.n8 VN.t1 172.202
R6 VN.n15 VN.t7 172.202
R7 VN.n21 VN.t4 172.202
R8 VN.n20 VN.t6 172.202
R9 VN.n32 VN.t0 172.202
R10 VN.n31 VN.n17 161.3
R11 VN.n30 VN.n29 161.3
R12 VN.n28 VN.n18 161.3
R13 VN.n27 VN.n26 161.3
R14 VN.n25 VN.n19 161.3
R15 VN.n24 VN.n23 161.3
R16 VN.n14 VN.n0 161.3
R17 VN.n13 VN.n12 161.3
R18 VN.n11 VN.n1 161.3
R19 VN.n10 VN.n9 161.3
R20 VN.n7 VN.n2 161.3
R21 VN.n6 VN.n5 161.3
R22 VN.n4 VN.n3 51.5382
R23 VN.n22 VN.n21 51.5382
R24 VN VN.n33 41.7069
R25 VN.n7 VN.n6 40.577
R26 VN.n9 VN.n7 40.577
R27 VN.n13 VN.n1 40.577
R28 VN.n14 VN.n13 40.577
R29 VN.n25 VN.n24 40.577
R30 VN.n26 VN.n25 40.577
R31 VN.n30 VN.n18 40.577
R32 VN.n31 VN.n30 40.577
R33 VN.n23 VN.n22 27.0073
R34 VN.n5 VN.n4 27.0073
R35 VN.n6 VN.n3 12.2964
R36 VN.n9 VN.n8 12.2964
R37 VN.n8 VN.n1 12.2964
R38 VN.n15 VN.n14 12.2964
R39 VN.n24 VN.n21 12.2964
R40 VN.n20 VN.n18 12.2964
R41 VN.n26 VN.n20 12.2964
R42 VN.n32 VN.n31 12.2964
R43 VN.n33 VN.n17 0.189894
R44 VN.n29 VN.n17 0.189894
R45 VN.n29 VN.n28 0.189894
R46 VN.n28 VN.n27 0.189894
R47 VN.n27 VN.n19 0.189894
R48 VN.n23 VN.n19 0.189894
R49 VN.n5 VN.n2 0.189894
R50 VN.n10 VN.n2 0.189894
R51 VN.n11 VN.n10 0.189894
R52 VN.n12 VN.n11 0.189894
R53 VN.n12 VN.n0 0.189894
R54 VN.n16 VN.n0 0.189894
R55 VN VN.n16 0.0516364
R56 VDD2.n2 VDD2.n1 68.1655
R57 VDD2.n2 VDD2.n0 68.1655
R58 VDD2 VDD2.n5 68.1627
R59 VDD2.n4 VDD2.n3 67.5745
R60 VDD2.n4 VDD2.n2 36.7412
R61 VDD2.n5 VDD2.t6 2.36892
R62 VDD2.n5 VDD2.t2 2.36892
R63 VDD2.n3 VDD2.t3 2.36892
R64 VDD2.n3 VDD2.t4 2.36892
R65 VDD2.n1 VDD2.t1 2.36892
R66 VDD2.n1 VDD2.t7 2.36892
R67 VDD2.n0 VDD2.t5 2.36892
R68 VDD2.n0 VDD2.t0 2.36892
R69 VDD2 VDD2.n4 0.705241
R70 VTAIL.n11 VTAIL.t6 53.2641
R71 VTAIL.n10 VTAIL.t12 53.2641
R72 VTAIL.n7 VTAIL.t15 53.2641
R73 VTAIL.n14 VTAIL.t1 53.264
R74 VTAIL.n15 VTAIL.t8 53.264
R75 VTAIL.n2 VTAIL.t10 53.264
R76 VTAIL.n3 VTAIL.t5 53.264
R77 VTAIL.n6 VTAIL.t4 53.264
R78 VTAIL.n13 VTAIL.n12 50.8957
R79 VTAIL.n9 VTAIL.n8 50.8957
R80 VTAIL.n1 VTAIL.n0 50.8955
R81 VTAIL.n5 VTAIL.n4 50.8955
R82 VTAIL.n15 VTAIL.n14 20.8669
R83 VTAIL.n7 VTAIL.n6 20.8669
R84 VTAIL.n0 VTAIL.t13 2.36892
R85 VTAIL.n0 VTAIL.t14 2.36892
R86 VTAIL.n4 VTAIL.t3 2.36892
R87 VTAIL.n4 VTAIL.t2 2.36892
R88 VTAIL.n12 VTAIL.t0 2.36892
R89 VTAIL.n12 VTAIL.t7 2.36892
R90 VTAIL.n8 VTAIL.t9 2.36892
R91 VTAIL.n8 VTAIL.t11 2.36892
R92 VTAIL.n9 VTAIL.n7 1.2936
R93 VTAIL.n10 VTAIL.n9 1.2936
R94 VTAIL.n13 VTAIL.n11 1.2936
R95 VTAIL.n14 VTAIL.n13 1.2936
R96 VTAIL.n6 VTAIL.n5 1.2936
R97 VTAIL.n5 VTAIL.n3 1.2936
R98 VTAIL.n2 VTAIL.n1 1.2936
R99 VTAIL VTAIL.n15 1.23541
R100 VTAIL.n11 VTAIL.n10 0.470328
R101 VTAIL.n3 VTAIL.n2 0.470328
R102 VTAIL VTAIL.n1 0.0586897
R103 B.n468 B.n467 585
R104 B.n468 B.n57 585
R105 B.n471 B.n470 585
R106 B.n472 B.n97 585
R107 B.n474 B.n473 585
R108 B.n476 B.n96 585
R109 B.n479 B.n478 585
R110 B.n480 B.n95 585
R111 B.n482 B.n481 585
R112 B.n484 B.n94 585
R113 B.n487 B.n486 585
R114 B.n488 B.n93 585
R115 B.n490 B.n489 585
R116 B.n492 B.n92 585
R117 B.n495 B.n494 585
R118 B.n496 B.n91 585
R119 B.n498 B.n497 585
R120 B.n500 B.n90 585
R121 B.n503 B.n502 585
R122 B.n504 B.n89 585
R123 B.n506 B.n505 585
R124 B.n508 B.n88 585
R125 B.n511 B.n510 585
R126 B.n512 B.n87 585
R127 B.n514 B.n513 585
R128 B.n516 B.n86 585
R129 B.n519 B.n518 585
R130 B.n520 B.n85 585
R131 B.n522 B.n521 585
R132 B.n524 B.n84 585
R133 B.n527 B.n526 585
R134 B.n528 B.n81 585
R135 B.n531 B.n530 585
R136 B.n533 B.n80 585
R137 B.n536 B.n535 585
R138 B.n537 B.n79 585
R139 B.n539 B.n538 585
R140 B.n541 B.n78 585
R141 B.n544 B.n543 585
R142 B.n545 B.n74 585
R143 B.n547 B.n546 585
R144 B.n549 B.n73 585
R145 B.n552 B.n551 585
R146 B.n553 B.n72 585
R147 B.n555 B.n554 585
R148 B.n557 B.n71 585
R149 B.n560 B.n559 585
R150 B.n561 B.n70 585
R151 B.n563 B.n562 585
R152 B.n565 B.n69 585
R153 B.n568 B.n567 585
R154 B.n569 B.n68 585
R155 B.n571 B.n570 585
R156 B.n573 B.n67 585
R157 B.n576 B.n575 585
R158 B.n577 B.n66 585
R159 B.n579 B.n578 585
R160 B.n581 B.n65 585
R161 B.n584 B.n583 585
R162 B.n585 B.n64 585
R163 B.n587 B.n586 585
R164 B.n589 B.n63 585
R165 B.n592 B.n591 585
R166 B.n593 B.n62 585
R167 B.n595 B.n594 585
R168 B.n597 B.n61 585
R169 B.n600 B.n599 585
R170 B.n601 B.n60 585
R171 B.n603 B.n602 585
R172 B.n605 B.n59 585
R173 B.n608 B.n607 585
R174 B.n609 B.n58 585
R175 B.n466 B.n56 585
R176 B.n612 B.n56 585
R177 B.n465 B.n55 585
R178 B.n613 B.n55 585
R179 B.n464 B.n54 585
R180 B.n614 B.n54 585
R181 B.n463 B.n462 585
R182 B.n462 B.n50 585
R183 B.n461 B.n49 585
R184 B.n620 B.n49 585
R185 B.n460 B.n48 585
R186 B.n621 B.n48 585
R187 B.n459 B.n47 585
R188 B.n622 B.n47 585
R189 B.n458 B.n457 585
R190 B.n457 B.n43 585
R191 B.n456 B.n42 585
R192 B.n628 B.n42 585
R193 B.n455 B.n41 585
R194 B.n629 B.n41 585
R195 B.n454 B.n40 585
R196 B.n630 B.n40 585
R197 B.n453 B.n452 585
R198 B.n452 B.n36 585
R199 B.n451 B.n35 585
R200 B.n636 B.n35 585
R201 B.n450 B.n34 585
R202 B.n637 B.n34 585
R203 B.n449 B.n33 585
R204 B.n638 B.n33 585
R205 B.n448 B.n447 585
R206 B.n447 B.n29 585
R207 B.n446 B.n28 585
R208 B.n644 B.n28 585
R209 B.n445 B.n27 585
R210 B.n645 B.n27 585
R211 B.n444 B.n26 585
R212 B.n646 B.n26 585
R213 B.n443 B.n442 585
R214 B.n442 B.n22 585
R215 B.n441 B.n21 585
R216 B.n652 B.n21 585
R217 B.n440 B.n20 585
R218 B.n653 B.n20 585
R219 B.n439 B.n19 585
R220 B.n654 B.n19 585
R221 B.n438 B.n437 585
R222 B.n437 B.n15 585
R223 B.n436 B.n14 585
R224 B.n660 B.n14 585
R225 B.n435 B.n13 585
R226 B.n661 B.n13 585
R227 B.n434 B.n12 585
R228 B.n662 B.n12 585
R229 B.n433 B.n432 585
R230 B.n432 B.n8 585
R231 B.n431 B.n7 585
R232 B.n668 B.n7 585
R233 B.n430 B.n6 585
R234 B.n669 B.n6 585
R235 B.n429 B.n5 585
R236 B.n670 B.n5 585
R237 B.n428 B.n427 585
R238 B.n427 B.n4 585
R239 B.n426 B.n98 585
R240 B.n426 B.n425 585
R241 B.n416 B.n99 585
R242 B.n100 B.n99 585
R243 B.n418 B.n417 585
R244 B.n419 B.n418 585
R245 B.n415 B.n105 585
R246 B.n105 B.n104 585
R247 B.n414 B.n413 585
R248 B.n413 B.n412 585
R249 B.n107 B.n106 585
R250 B.n108 B.n107 585
R251 B.n405 B.n404 585
R252 B.n406 B.n405 585
R253 B.n403 B.n112 585
R254 B.n116 B.n112 585
R255 B.n402 B.n401 585
R256 B.n401 B.n400 585
R257 B.n114 B.n113 585
R258 B.n115 B.n114 585
R259 B.n393 B.n392 585
R260 B.n394 B.n393 585
R261 B.n391 B.n120 585
R262 B.n124 B.n120 585
R263 B.n390 B.n389 585
R264 B.n389 B.n388 585
R265 B.n122 B.n121 585
R266 B.n123 B.n122 585
R267 B.n381 B.n380 585
R268 B.n382 B.n381 585
R269 B.n379 B.n129 585
R270 B.n129 B.n128 585
R271 B.n378 B.n377 585
R272 B.n377 B.n376 585
R273 B.n131 B.n130 585
R274 B.n132 B.n131 585
R275 B.n369 B.n368 585
R276 B.n370 B.n369 585
R277 B.n367 B.n137 585
R278 B.n137 B.n136 585
R279 B.n366 B.n365 585
R280 B.n365 B.n364 585
R281 B.n139 B.n138 585
R282 B.n140 B.n139 585
R283 B.n357 B.n356 585
R284 B.n358 B.n357 585
R285 B.n355 B.n144 585
R286 B.n148 B.n144 585
R287 B.n354 B.n353 585
R288 B.n353 B.n352 585
R289 B.n146 B.n145 585
R290 B.n147 B.n146 585
R291 B.n345 B.n344 585
R292 B.n346 B.n345 585
R293 B.n343 B.n153 585
R294 B.n153 B.n152 585
R295 B.n342 B.n341 585
R296 B.n341 B.n340 585
R297 B.n337 B.n157 585
R298 B.n336 B.n335 585
R299 B.n333 B.n158 585
R300 B.n333 B.n156 585
R301 B.n332 B.n331 585
R302 B.n330 B.n329 585
R303 B.n328 B.n160 585
R304 B.n326 B.n325 585
R305 B.n324 B.n161 585
R306 B.n323 B.n322 585
R307 B.n320 B.n162 585
R308 B.n318 B.n317 585
R309 B.n316 B.n163 585
R310 B.n315 B.n314 585
R311 B.n312 B.n164 585
R312 B.n310 B.n309 585
R313 B.n308 B.n165 585
R314 B.n307 B.n306 585
R315 B.n304 B.n166 585
R316 B.n302 B.n301 585
R317 B.n300 B.n167 585
R318 B.n299 B.n298 585
R319 B.n296 B.n168 585
R320 B.n294 B.n293 585
R321 B.n292 B.n169 585
R322 B.n291 B.n290 585
R323 B.n288 B.n170 585
R324 B.n286 B.n285 585
R325 B.n284 B.n171 585
R326 B.n283 B.n282 585
R327 B.n280 B.n172 585
R328 B.n278 B.n277 585
R329 B.n275 B.n173 585
R330 B.n274 B.n273 585
R331 B.n271 B.n176 585
R332 B.n269 B.n268 585
R333 B.n267 B.n177 585
R334 B.n266 B.n265 585
R335 B.n263 B.n178 585
R336 B.n261 B.n260 585
R337 B.n259 B.n179 585
R338 B.n257 B.n256 585
R339 B.n254 B.n182 585
R340 B.n252 B.n251 585
R341 B.n250 B.n183 585
R342 B.n249 B.n248 585
R343 B.n246 B.n184 585
R344 B.n244 B.n243 585
R345 B.n242 B.n185 585
R346 B.n241 B.n240 585
R347 B.n238 B.n186 585
R348 B.n236 B.n235 585
R349 B.n234 B.n187 585
R350 B.n233 B.n232 585
R351 B.n230 B.n188 585
R352 B.n228 B.n227 585
R353 B.n226 B.n189 585
R354 B.n225 B.n224 585
R355 B.n222 B.n190 585
R356 B.n220 B.n219 585
R357 B.n218 B.n191 585
R358 B.n217 B.n216 585
R359 B.n214 B.n192 585
R360 B.n212 B.n211 585
R361 B.n210 B.n193 585
R362 B.n209 B.n208 585
R363 B.n206 B.n194 585
R364 B.n204 B.n203 585
R365 B.n202 B.n195 585
R366 B.n201 B.n200 585
R367 B.n198 B.n196 585
R368 B.n155 B.n154 585
R369 B.n339 B.n338 585
R370 B.n340 B.n339 585
R371 B.n151 B.n150 585
R372 B.n152 B.n151 585
R373 B.n348 B.n347 585
R374 B.n347 B.n346 585
R375 B.n349 B.n149 585
R376 B.n149 B.n147 585
R377 B.n351 B.n350 585
R378 B.n352 B.n351 585
R379 B.n143 B.n142 585
R380 B.n148 B.n143 585
R381 B.n360 B.n359 585
R382 B.n359 B.n358 585
R383 B.n361 B.n141 585
R384 B.n141 B.n140 585
R385 B.n363 B.n362 585
R386 B.n364 B.n363 585
R387 B.n135 B.n134 585
R388 B.n136 B.n135 585
R389 B.n372 B.n371 585
R390 B.n371 B.n370 585
R391 B.n373 B.n133 585
R392 B.n133 B.n132 585
R393 B.n375 B.n374 585
R394 B.n376 B.n375 585
R395 B.n127 B.n126 585
R396 B.n128 B.n127 585
R397 B.n384 B.n383 585
R398 B.n383 B.n382 585
R399 B.n385 B.n125 585
R400 B.n125 B.n123 585
R401 B.n387 B.n386 585
R402 B.n388 B.n387 585
R403 B.n119 B.n118 585
R404 B.n124 B.n119 585
R405 B.n396 B.n395 585
R406 B.n395 B.n394 585
R407 B.n397 B.n117 585
R408 B.n117 B.n115 585
R409 B.n399 B.n398 585
R410 B.n400 B.n399 585
R411 B.n111 B.n110 585
R412 B.n116 B.n111 585
R413 B.n408 B.n407 585
R414 B.n407 B.n406 585
R415 B.n409 B.n109 585
R416 B.n109 B.n108 585
R417 B.n411 B.n410 585
R418 B.n412 B.n411 585
R419 B.n103 B.n102 585
R420 B.n104 B.n103 585
R421 B.n421 B.n420 585
R422 B.n420 B.n419 585
R423 B.n422 B.n101 585
R424 B.n101 B.n100 585
R425 B.n424 B.n423 585
R426 B.n425 B.n424 585
R427 B.n2 B.n0 585
R428 B.n4 B.n2 585
R429 B.n3 B.n1 585
R430 B.n669 B.n3 585
R431 B.n667 B.n666 585
R432 B.n668 B.n667 585
R433 B.n665 B.n9 585
R434 B.n9 B.n8 585
R435 B.n664 B.n663 585
R436 B.n663 B.n662 585
R437 B.n11 B.n10 585
R438 B.n661 B.n11 585
R439 B.n659 B.n658 585
R440 B.n660 B.n659 585
R441 B.n657 B.n16 585
R442 B.n16 B.n15 585
R443 B.n656 B.n655 585
R444 B.n655 B.n654 585
R445 B.n18 B.n17 585
R446 B.n653 B.n18 585
R447 B.n651 B.n650 585
R448 B.n652 B.n651 585
R449 B.n649 B.n23 585
R450 B.n23 B.n22 585
R451 B.n648 B.n647 585
R452 B.n647 B.n646 585
R453 B.n25 B.n24 585
R454 B.n645 B.n25 585
R455 B.n643 B.n642 585
R456 B.n644 B.n643 585
R457 B.n641 B.n30 585
R458 B.n30 B.n29 585
R459 B.n640 B.n639 585
R460 B.n639 B.n638 585
R461 B.n32 B.n31 585
R462 B.n637 B.n32 585
R463 B.n635 B.n634 585
R464 B.n636 B.n635 585
R465 B.n633 B.n37 585
R466 B.n37 B.n36 585
R467 B.n632 B.n631 585
R468 B.n631 B.n630 585
R469 B.n39 B.n38 585
R470 B.n629 B.n39 585
R471 B.n627 B.n626 585
R472 B.n628 B.n627 585
R473 B.n625 B.n44 585
R474 B.n44 B.n43 585
R475 B.n624 B.n623 585
R476 B.n623 B.n622 585
R477 B.n46 B.n45 585
R478 B.n621 B.n46 585
R479 B.n619 B.n618 585
R480 B.n620 B.n619 585
R481 B.n617 B.n51 585
R482 B.n51 B.n50 585
R483 B.n616 B.n615 585
R484 B.n615 B.n614 585
R485 B.n53 B.n52 585
R486 B.n613 B.n53 585
R487 B.n611 B.n610 585
R488 B.n612 B.n611 585
R489 B.n672 B.n671 585
R490 B.n671 B.n670 585
R491 B.n339 B.n157 559.769
R492 B.n611 B.n58 559.769
R493 B.n341 B.n155 559.769
R494 B.n468 B.n56 559.769
R495 B.n180 B.t19 376.159
R496 B.n174 B.t12 376.159
R497 B.n75 B.t8 376.159
R498 B.n82 B.t16 376.159
R499 B.n469 B.n57 256.663
R500 B.n475 B.n57 256.663
R501 B.n477 B.n57 256.663
R502 B.n483 B.n57 256.663
R503 B.n485 B.n57 256.663
R504 B.n491 B.n57 256.663
R505 B.n493 B.n57 256.663
R506 B.n499 B.n57 256.663
R507 B.n501 B.n57 256.663
R508 B.n507 B.n57 256.663
R509 B.n509 B.n57 256.663
R510 B.n515 B.n57 256.663
R511 B.n517 B.n57 256.663
R512 B.n523 B.n57 256.663
R513 B.n525 B.n57 256.663
R514 B.n532 B.n57 256.663
R515 B.n534 B.n57 256.663
R516 B.n540 B.n57 256.663
R517 B.n542 B.n57 256.663
R518 B.n548 B.n57 256.663
R519 B.n550 B.n57 256.663
R520 B.n556 B.n57 256.663
R521 B.n558 B.n57 256.663
R522 B.n564 B.n57 256.663
R523 B.n566 B.n57 256.663
R524 B.n572 B.n57 256.663
R525 B.n574 B.n57 256.663
R526 B.n580 B.n57 256.663
R527 B.n582 B.n57 256.663
R528 B.n588 B.n57 256.663
R529 B.n590 B.n57 256.663
R530 B.n596 B.n57 256.663
R531 B.n598 B.n57 256.663
R532 B.n604 B.n57 256.663
R533 B.n606 B.n57 256.663
R534 B.n334 B.n156 256.663
R535 B.n159 B.n156 256.663
R536 B.n327 B.n156 256.663
R537 B.n321 B.n156 256.663
R538 B.n319 B.n156 256.663
R539 B.n313 B.n156 256.663
R540 B.n311 B.n156 256.663
R541 B.n305 B.n156 256.663
R542 B.n303 B.n156 256.663
R543 B.n297 B.n156 256.663
R544 B.n295 B.n156 256.663
R545 B.n289 B.n156 256.663
R546 B.n287 B.n156 256.663
R547 B.n281 B.n156 256.663
R548 B.n279 B.n156 256.663
R549 B.n272 B.n156 256.663
R550 B.n270 B.n156 256.663
R551 B.n264 B.n156 256.663
R552 B.n262 B.n156 256.663
R553 B.n255 B.n156 256.663
R554 B.n253 B.n156 256.663
R555 B.n247 B.n156 256.663
R556 B.n245 B.n156 256.663
R557 B.n239 B.n156 256.663
R558 B.n237 B.n156 256.663
R559 B.n231 B.n156 256.663
R560 B.n229 B.n156 256.663
R561 B.n223 B.n156 256.663
R562 B.n221 B.n156 256.663
R563 B.n215 B.n156 256.663
R564 B.n213 B.n156 256.663
R565 B.n207 B.n156 256.663
R566 B.n205 B.n156 256.663
R567 B.n199 B.n156 256.663
R568 B.n197 B.n156 256.663
R569 B.n339 B.n151 163.367
R570 B.n347 B.n151 163.367
R571 B.n347 B.n149 163.367
R572 B.n351 B.n149 163.367
R573 B.n351 B.n143 163.367
R574 B.n359 B.n143 163.367
R575 B.n359 B.n141 163.367
R576 B.n363 B.n141 163.367
R577 B.n363 B.n135 163.367
R578 B.n371 B.n135 163.367
R579 B.n371 B.n133 163.367
R580 B.n375 B.n133 163.367
R581 B.n375 B.n127 163.367
R582 B.n383 B.n127 163.367
R583 B.n383 B.n125 163.367
R584 B.n387 B.n125 163.367
R585 B.n387 B.n119 163.367
R586 B.n395 B.n119 163.367
R587 B.n395 B.n117 163.367
R588 B.n399 B.n117 163.367
R589 B.n399 B.n111 163.367
R590 B.n407 B.n111 163.367
R591 B.n407 B.n109 163.367
R592 B.n411 B.n109 163.367
R593 B.n411 B.n103 163.367
R594 B.n420 B.n103 163.367
R595 B.n420 B.n101 163.367
R596 B.n424 B.n101 163.367
R597 B.n424 B.n2 163.367
R598 B.n671 B.n2 163.367
R599 B.n671 B.n3 163.367
R600 B.n667 B.n3 163.367
R601 B.n667 B.n9 163.367
R602 B.n663 B.n9 163.367
R603 B.n663 B.n11 163.367
R604 B.n659 B.n11 163.367
R605 B.n659 B.n16 163.367
R606 B.n655 B.n16 163.367
R607 B.n655 B.n18 163.367
R608 B.n651 B.n18 163.367
R609 B.n651 B.n23 163.367
R610 B.n647 B.n23 163.367
R611 B.n647 B.n25 163.367
R612 B.n643 B.n25 163.367
R613 B.n643 B.n30 163.367
R614 B.n639 B.n30 163.367
R615 B.n639 B.n32 163.367
R616 B.n635 B.n32 163.367
R617 B.n635 B.n37 163.367
R618 B.n631 B.n37 163.367
R619 B.n631 B.n39 163.367
R620 B.n627 B.n39 163.367
R621 B.n627 B.n44 163.367
R622 B.n623 B.n44 163.367
R623 B.n623 B.n46 163.367
R624 B.n619 B.n46 163.367
R625 B.n619 B.n51 163.367
R626 B.n615 B.n51 163.367
R627 B.n615 B.n53 163.367
R628 B.n611 B.n53 163.367
R629 B.n335 B.n333 163.367
R630 B.n333 B.n332 163.367
R631 B.n329 B.n328 163.367
R632 B.n326 B.n161 163.367
R633 B.n322 B.n320 163.367
R634 B.n318 B.n163 163.367
R635 B.n314 B.n312 163.367
R636 B.n310 B.n165 163.367
R637 B.n306 B.n304 163.367
R638 B.n302 B.n167 163.367
R639 B.n298 B.n296 163.367
R640 B.n294 B.n169 163.367
R641 B.n290 B.n288 163.367
R642 B.n286 B.n171 163.367
R643 B.n282 B.n280 163.367
R644 B.n278 B.n173 163.367
R645 B.n273 B.n271 163.367
R646 B.n269 B.n177 163.367
R647 B.n265 B.n263 163.367
R648 B.n261 B.n179 163.367
R649 B.n256 B.n254 163.367
R650 B.n252 B.n183 163.367
R651 B.n248 B.n246 163.367
R652 B.n244 B.n185 163.367
R653 B.n240 B.n238 163.367
R654 B.n236 B.n187 163.367
R655 B.n232 B.n230 163.367
R656 B.n228 B.n189 163.367
R657 B.n224 B.n222 163.367
R658 B.n220 B.n191 163.367
R659 B.n216 B.n214 163.367
R660 B.n212 B.n193 163.367
R661 B.n208 B.n206 163.367
R662 B.n204 B.n195 163.367
R663 B.n200 B.n198 163.367
R664 B.n341 B.n153 163.367
R665 B.n345 B.n153 163.367
R666 B.n345 B.n146 163.367
R667 B.n353 B.n146 163.367
R668 B.n353 B.n144 163.367
R669 B.n357 B.n144 163.367
R670 B.n357 B.n139 163.367
R671 B.n365 B.n139 163.367
R672 B.n365 B.n137 163.367
R673 B.n369 B.n137 163.367
R674 B.n369 B.n131 163.367
R675 B.n377 B.n131 163.367
R676 B.n377 B.n129 163.367
R677 B.n381 B.n129 163.367
R678 B.n381 B.n122 163.367
R679 B.n389 B.n122 163.367
R680 B.n389 B.n120 163.367
R681 B.n393 B.n120 163.367
R682 B.n393 B.n114 163.367
R683 B.n401 B.n114 163.367
R684 B.n401 B.n112 163.367
R685 B.n405 B.n112 163.367
R686 B.n405 B.n107 163.367
R687 B.n413 B.n107 163.367
R688 B.n413 B.n105 163.367
R689 B.n418 B.n105 163.367
R690 B.n418 B.n99 163.367
R691 B.n426 B.n99 163.367
R692 B.n427 B.n426 163.367
R693 B.n427 B.n5 163.367
R694 B.n6 B.n5 163.367
R695 B.n7 B.n6 163.367
R696 B.n432 B.n7 163.367
R697 B.n432 B.n12 163.367
R698 B.n13 B.n12 163.367
R699 B.n14 B.n13 163.367
R700 B.n437 B.n14 163.367
R701 B.n437 B.n19 163.367
R702 B.n20 B.n19 163.367
R703 B.n21 B.n20 163.367
R704 B.n442 B.n21 163.367
R705 B.n442 B.n26 163.367
R706 B.n27 B.n26 163.367
R707 B.n28 B.n27 163.367
R708 B.n447 B.n28 163.367
R709 B.n447 B.n33 163.367
R710 B.n34 B.n33 163.367
R711 B.n35 B.n34 163.367
R712 B.n452 B.n35 163.367
R713 B.n452 B.n40 163.367
R714 B.n41 B.n40 163.367
R715 B.n42 B.n41 163.367
R716 B.n457 B.n42 163.367
R717 B.n457 B.n47 163.367
R718 B.n48 B.n47 163.367
R719 B.n49 B.n48 163.367
R720 B.n462 B.n49 163.367
R721 B.n462 B.n54 163.367
R722 B.n55 B.n54 163.367
R723 B.n56 B.n55 163.367
R724 B.n607 B.n605 163.367
R725 B.n603 B.n60 163.367
R726 B.n599 B.n597 163.367
R727 B.n595 B.n62 163.367
R728 B.n591 B.n589 163.367
R729 B.n587 B.n64 163.367
R730 B.n583 B.n581 163.367
R731 B.n579 B.n66 163.367
R732 B.n575 B.n573 163.367
R733 B.n571 B.n68 163.367
R734 B.n567 B.n565 163.367
R735 B.n563 B.n70 163.367
R736 B.n559 B.n557 163.367
R737 B.n555 B.n72 163.367
R738 B.n551 B.n549 163.367
R739 B.n547 B.n74 163.367
R740 B.n543 B.n541 163.367
R741 B.n539 B.n79 163.367
R742 B.n535 B.n533 163.367
R743 B.n531 B.n81 163.367
R744 B.n526 B.n524 163.367
R745 B.n522 B.n85 163.367
R746 B.n518 B.n516 163.367
R747 B.n514 B.n87 163.367
R748 B.n510 B.n508 163.367
R749 B.n506 B.n89 163.367
R750 B.n502 B.n500 163.367
R751 B.n498 B.n91 163.367
R752 B.n494 B.n492 163.367
R753 B.n490 B.n93 163.367
R754 B.n486 B.n484 163.367
R755 B.n482 B.n95 163.367
R756 B.n478 B.n476 163.367
R757 B.n474 B.n97 163.367
R758 B.n470 B.n468 163.367
R759 B.n340 B.n156 108.912
R760 B.n612 B.n57 108.912
R761 B.n180 B.t21 101.474
R762 B.n82 B.t17 101.474
R763 B.n174 B.t15 101.463
R764 B.n75 B.t10 101.463
R765 B.n181 B.t20 72.3821
R766 B.n83 B.t18 72.3821
R767 B.n175 B.t14 72.3723
R768 B.n76 B.t11 72.3723
R769 B.n334 B.n157 71.676
R770 B.n332 B.n159 71.676
R771 B.n328 B.n327 71.676
R772 B.n321 B.n161 71.676
R773 B.n320 B.n319 71.676
R774 B.n313 B.n163 71.676
R775 B.n312 B.n311 71.676
R776 B.n305 B.n165 71.676
R777 B.n304 B.n303 71.676
R778 B.n297 B.n167 71.676
R779 B.n296 B.n295 71.676
R780 B.n289 B.n169 71.676
R781 B.n288 B.n287 71.676
R782 B.n281 B.n171 71.676
R783 B.n280 B.n279 71.676
R784 B.n272 B.n173 71.676
R785 B.n271 B.n270 71.676
R786 B.n264 B.n177 71.676
R787 B.n263 B.n262 71.676
R788 B.n255 B.n179 71.676
R789 B.n254 B.n253 71.676
R790 B.n247 B.n183 71.676
R791 B.n246 B.n245 71.676
R792 B.n239 B.n185 71.676
R793 B.n238 B.n237 71.676
R794 B.n231 B.n187 71.676
R795 B.n230 B.n229 71.676
R796 B.n223 B.n189 71.676
R797 B.n222 B.n221 71.676
R798 B.n215 B.n191 71.676
R799 B.n214 B.n213 71.676
R800 B.n207 B.n193 71.676
R801 B.n206 B.n205 71.676
R802 B.n199 B.n195 71.676
R803 B.n198 B.n197 71.676
R804 B.n606 B.n58 71.676
R805 B.n605 B.n604 71.676
R806 B.n598 B.n60 71.676
R807 B.n597 B.n596 71.676
R808 B.n590 B.n62 71.676
R809 B.n589 B.n588 71.676
R810 B.n582 B.n64 71.676
R811 B.n581 B.n580 71.676
R812 B.n574 B.n66 71.676
R813 B.n573 B.n572 71.676
R814 B.n566 B.n68 71.676
R815 B.n565 B.n564 71.676
R816 B.n558 B.n70 71.676
R817 B.n557 B.n556 71.676
R818 B.n550 B.n72 71.676
R819 B.n549 B.n548 71.676
R820 B.n542 B.n74 71.676
R821 B.n541 B.n540 71.676
R822 B.n534 B.n79 71.676
R823 B.n533 B.n532 71.676
R824 B.n525 B.n81 71.676
R825 B.n524 B.n523 71.676
R826 B.n517 B.n85 71.676
R827 B.n516 B.n515 71.676
R828 B.n509 B.n87 71.676
R829 B.n508 B.n507 71.676
R830 B.n501 B.n89 71.676
R831 B.n500 B.n499 71.676
R832 B.n493 B.n91 71.676
R833 B.n492 B.n491 71.676
R834 B.n485 B.n93 71.676
R835 B.n484 B.n483 71.676
R836 B.n477 B.n95 71.676
R837 B.n476 B.n475 71.676
R838 B.n469 B.n97 71.676
R839 B.n470 B.n469 71.676
R840 B.n475 B.n474 71.676
R841 B.n478 B.n477 71.676
R842 B.n483 B.n482 71.676
R843 B.n486 B.n485 71.676
R844 B.n491 B.n490 71.676
R845 B.n494 B.n493 71.676
R846 B.n499 B.n498 71.676
R847 B.n502 B.n501 71.676
R848 B.n507 B.n506 71.676
R849 B.n510 B.n509 71.676
R850 B.n515 B.n514 71.676
R851 B.n518 B.n517 71.676
R852 B.n523 B.n522 71.676
R853 B.n526 B.n525 71.676
R854 B.n532 B.n531 71.676
R855 B.n535 B.n534 71.676
R856 B.n540 B.n539 71.676
R857 B.n543 B.n542 71.676
R858 B.n548 B.n547 71.676
R859 B.n551 B.n550 71.676
R860 B.n556 B.n555 71.676
R861 B.n559 B.n558 71.676
R862 B.n564 B.n563 71.676
R863 B.n567 B.n566 71.676
R864 B.n572 B.n571 71.676
R865 B.n575 B.n574 71.676
R866 B.n580 B.n579 71.676
R867 B.n583 B.n582 71.676
R868 B.n588 B.n587 71.676
R869 B.n591 B.n590 71.676
R870 B.n596 B.n595 71.676
R871 B.n599 B.n598 71.676
R872 B.n604 B.n603 71.676
R873 B.n607 B.n606 71.676
R874 B.n335 B.n334 71.676
R875 B.n329 B.n159 71.676
R876 B.n327 B.n326 71.676
R877 B.n322 B.n321 71.676
R878 B.n319 B.n318 71.676
R879 B.n314 B.n313 71.676
R880 B.n311 B.n310 71.676
R881 B.n306 B.n305 71.676
R882 B.n303 B.n302 71.676
R883 B.n298 B.n297 71.676
R884 B.n295 B.n294 71.676
R885 B.n290 B.n289 71.676
R886 B.n287 B.n286 71.676
R887 B.n282 B.n281 71.676
R888 B.n279 B.n278 71.676
R889 B.n273 B.n272 71.676
R890 B.n270 B.n269 71.676
R891 B.n265 B.n264 71.676
R892 B.n262 B.n261 71.676
R893 B.n256 B.n255 71.676
R894 B.n253 B.n252 71.676
R895 B.n248 B.n247 71.676
R896 B.n245 B.n244 71.676
R897 B.n240 B.n239 71.676
R898 B.n237 B.n236 71.676
R899 B.n232 B.n231 71.676
R900 B.n229 B.n228 71.676
R901 B.n224 B.n223 71.676
R902 B.n221 B.n220 71.676
R903 B.n216 B.n215 71.676
R904 B.n213 B.n212 71.676
R905 B.n208 B.n207 71.676
R906 B.n205 B.n204 71.676
R907 B.n200 B.n199 71.676
R908 B.n197 B.n155 71.676
R909 B.n258 B.n181 59.5399
R910 B.n276 B.n175 59.5399
R911 B.n77 B.n76 59.5399
R912 B.n529 B.n83 59.5399
R913 B.n340 B.n152 54.8593
R914 B.n346 B.n152 54.8593
R915 B.n346 B.n147 54.8593
R916 B.n352 B.n147 54.8593
R917 B.n352 B.n148 54.8593
R918 B.n358 B.n140 54.8593
R919 B.n364 B.n140 54.8593
R920 B.n364 B.n136 54.8593
R921 B.n370 B.n136 54.8593
R922 B.n370 B.n132 54.8593
R923 B.n376 B.n132 54.8593
R924 B.n382 B.n128 54.8593
R925 B.n382 B.n123 54.8593
R926 B.n388 B.n123 54.8593
R927 B.n388 B.n124 54.8593
R928 B.n394 B.n115 54.8593
R929 B.n400 B.n115 54.8593
R930 B.n400 B.n116 54.8593
R931 B.n406 B.n108 54.8593
R932 B.n412 B.n108 54.8593
R933 B.n412 B.n104 54.8593
R934 B.n419 B.n104 54.8593
R935 B.n425 B.n100 54.8593
R936 B.n425 B.n4 54.8593
R937 B.n670 B.n4 54.8593
R938 B.n670 B.n669 54.8593
R939 B.n669 B.n668 54.8593
R940 B.n668 B.n8 54.8593
R941 B.n662 B.n661 54.8593
R942 B.n661 B.n660 54.8593
R943 B.n660 B.n15 54.8593
R944 B.n654 B.n15 54.8593
R945 B.n653 B.n652 54.8593
R946 B.n652 B.n22 54.8593
R947 B.n646 B.n22 54.8593
R948 B.n645 B.n644 54.8593
R949 B.n644 B.n29 54.8593
R950 B.n638 B.n29 54.8593
R951 B.n638 B.n637 54.8593
R952 B.n636 B.n36 54.8593
R953 B.n630 B.n36 54.8593
R954 B.n630 B.n629 54.8593
R955 B.n629 B.n628 54.8593
R956 B.n628 B.n43 54.8593
R957 B.n622 B.n43 54.8593
R958 B.n621 B.n620 54.8593
R959 B.n620 B.n50 54.8593
R960 B.n614 B.n50 54.8593
R961 B.n614 B.n613 54.8593
R962 B.n613 B.n612 54.8593
R963 B.n376 B.t4 52.4391
R964 B.t1 B.n636 52.4391
R965 B.t5 B.n100 44.3716
R966 B.t6 B.n8 44.3716
R967 B.n116 B.t2 42.7581
R968 B.t0 B.n653 42.7581
R969 B.n610 B.n609 36.3712
R970 B.n467 B.n466 36.3712
R971 B.n342 B.n154 36.3712
R972 B.n338 B.n337 36.3712
R973 B.n358 B.t13 36.3041
R974 B.n622 B.t9 36.3041
R975 B.n394 B.t3 34.6906
R976 B.n646 B.t7 34.6906
R977 B.n181 B.n180 29.0914
R978 B.n175 B.n174 29.0914
R979 B.n76 B.n75 29.0914
R980 B.n83 B.n82 29.0914
R981 B.n124 B.t3 20.1692
R982 B.t7 B.n645 20.1692
R983 B.n148 B.t13 18.5557
R984 B.t9 B.n621 18.5557
R985 B B.n672 18.0485
R986 B.n406 B.t2 12.1017
R987 B.n654 B.t0 12.1017
R988 B.n609 B.n608 10.6151
R989 B.n608 B.n59 10.6151
R990 B.n602 B.n59 10.6151
R991 B.n602 B.n601 10.6151
R992 B.n601 B.n600 10.6151
R993 B.n600 B.n61 10.6151
R994 B.n594 B.n61 10.6151
R995 B.n594 B.n593 10.6151
R996 B.n593 B.n592 10.6151
R997 B.n592 B.n63 10.6151
R998 B.n586 B.n63 10.6151
R999 B.n586 B.n585 10.6151
R1000 B.n585 B.n584 10.6151
R1001 B.n584 B.n65 10.6151
R1002 B.n578 B.n65 10.6151
R1003 B.n578 B.n577 10.6151
R1004 B.n577 B.n576 10.6151
R1005 B.n576 B.n67 10.6151
R1006 B.n570 B.n67 10.6151
R1007 B.n570 B.n569 10.6151
R1008 B.n569 B.n568 10.6151
R1009 B.n568 B.n69 10.6151
R1010 B.n562 B.n69 10.6151
R1011 B.n562 B.n561 10.6151
R1012 B.n561 B.n560 10.6151
R1013 B.n560 B.n71 10.6151
R1014 B.n554 B.n71 10.6151
R1015 B.n554 B.n553 10.6151
R1016 B.n553 B.n552 10.6151
R1017 B.n552 B.n73 10.6151
R1018 B.n546 B.n545 10.6151
R1019 B.n545 B.n544 10.6151
R1020 B.n544 B.n78 10.6151
R1021 B.n538 B.n78 10.6151
R1022 B.n538 B.n537 10.6151
R1023 B.n537 B.n536 10.6151
R1024 B.n536 B.n80 10.6151
R1025 B.n530 B.n80 10.6151
R1026 B.n528 B.n527 10.6151
R1027 B.n527 B.n84 10.6151
R1028 B.n521 B.n84 10.6151
R1029 B.n521 B.n520 10.6151
R1030 B.n520 B.n519 10.6151
R1031 B.n519 B.n86 10.6151
R1032 B.n513 B.n86 10.6151
R1033 B.n513 B.n512 10.6151
R1034 B.n512 B.n511 10.6151
R1035 B.n511 B.n88 10.6151
R1036 B.n505 B.n88 10.6151
R1037 B.n505 B.n504 10.6151
R1038 B.n504 B.n503 10.6151
R1039 B.n503 B.n90 10.6151
R1040 B.n497 B.n90 10.6151
R1041 B.n497 B.n496 10.6151
R1042 B.n496 B.n495 10.6151
R1043 B.n495 B.n92 10.6151
R1044 B.n489 B.n92 10.6151
R1045 B.n489 B.n488 10.6151
R1046 B.n488 B.n487 10.6151
R1047 B.n487 B.n94 10.6151
R1048 B.n481 B.n94 10.6151
R1049 B.n481 B.n480 10.6151
R1050 B.n480 B.n479 10.6151
R1051 B.n479 B.n96 10.6151
R1052 B.n473 B.n96 10.6151
R1053 B.n473 B.n472 10.6151
R1054 B.n472 B.n471 10.6151
R1055 B.n471 B.n467 10.6151
R1056 B.n343 B.n342 10.6151
R1057 B.n344 B.n343 10.6151
R1058 B.n344 B.n145 10.6151
R1059 B.n354 B.n145 10.6151
R1060 B.n355 B.n354 10.6151
R1061 B.n356 B.n355 10.6151
R1062 B.n356 B.n138 10.6151
R1063 B.n366 B.n138 10.6151
R1064 B.n367 B.n366 10.6151
R1065 B.n368 B.n367 10.6151
R1066 B.n368 B.n130 10.6151
R1067 B.n378 B.n130 10.6151
R1068 B.n379 B.n378 10.6151
R1069 B.n380 B.n379 10.6151
R1070 B.n380 B.n121 10.6151
R1071 B.n390 B.n121 10.6151
R1072 B.n391 B.n390 10.6151
R1073 B.n392 B.n391 10.6151
R1074 B.n392 B.n113 10.6151
R1075 B.n402 B.n113 10.6151
R1076 B.n403 B.n402 10.6151
R1077 B.n404 B.n403 10.6151
R1078 B.n404 B.n106 10.6151
R1079 B.n414 B.n106 10.6151
R1080 B.n415 B.n414 10.6151
R1081 B.n417 B.n415 10.6151
R1082 B.n417 B.n416 10.6151
R1083 B.n416 B.n98 10.6151
R1084 B.n428 B.n98 10.6151
R1085 B.n429 B.n428 10.6151
R1086 B.n430 B.n429 10.6151
R1087 B.n431 B.n430 10.6151
R1088 B.n433 B.n431 10.6151
R1089 B.n434 B.n433 10.6151
R1090 B.n435 B.n434 10.6151
R1091 B.n436 B.n435 10.6151
R1092 B.n438 B.n436 10.6151
R1093 B.n439 B.n438 10.6151
R1094 B.n440 B.n439 10.6151
R1095 B.n441 B.n440 10.6151
R1096 B.n443 B.n441 10.6151
R1097 B.n444 B.n443 10.6151
R1098 B.n445 B.n444 10.6151
R1099 B.n446 B.n445 10.6151
R1100 B.n448 B.n446 10.6151
R1101 B.n449 B.n448 10.6151
R1102 B.n450 B.n449 10.6151
R1103 B.n451 B.n450 10.6151
R1104 B.n453 B.n451 10.6151
R1105 B.n454 B.n453 10.6151
R1106 B.n455 B.n454 10.6151
R1107 B.n456 B.n455 10.6151
R1108 B.n458 B.n456 10.6151
R1109 B.n459 B.n458 10.6151
R1110 B.n460 B.n459 10.6151
R1111 B.n461 B.n460 10.6151
R1112 B.n463 B.n461 10.6151
R1113 B.n464 B.n463 10.6151
R1114 B.n465 B.n464 10.6151
R1115 B.n466 B.n465 10.6151
R1116 B.n337 B.n336 10.6151
R1117 B.n336 B.n158 10.6151
R1118 B.n331 B.n158 10.6151
R1119 B.n331 B.n330 10.6151
R1120 B.n330 B.n160 10.6151
R1121 B.n325 B.n160 10.6151
R1122 B.n325 B.n324 10.6151
R1123 B.n324 B.n323 10.6151
R1124 B.n323 B.n162 10.6151
R1125 B.n317 B.n162 10.6151
R1126 B.n317 B.n316 10.6151
R1127 B.n316 B.n315 10.6151
R1128 B.n315 B.n164 10.6151
R1129 B.n309 B.n164 10.6151
R1130 B.n309 B.n308 10.6151
R1131 B.n308 B.n307 10.6151
R1132 B.n307 B.n166 10.6151
R1133 B.n301 B.n166 10.6151
R1134 B.n301 B.n300 10.6151
R1135 B.n300 B.n299 10.6151
R1136 B.n299 B.n168 10.6151
R1137 B.n293 B.n168 10.6151
R1138 B.n293 B.n292 10.6151
R1139 B.n292 B.n291 10.6151
R1140 B.n291 B.n170 10.6151
R1141 B.n285 B.n170 10.6151
R1142 B.n285 B.n284 10.6151
R1143 B.n284 B.n283 10.6151
R1144 B.n283 B.n172 10.6151
R1145 B.n277 B.n172 10.6151
R1146 B.n275 B.n274 10.6151
R1147 B.n274 B.n176 10.6151
R1148 B.n268 B.n176 10.6151
R1149 B.n268 B.n267 10.6151
R1150 B.n267 B.n266 10.6151
R1151 B.n266 B.n178 10.6151
R1152 B.n260 B.n178 10.6151
R1153 B.n260 B.n259 10.6151
R1154 B.n257 B.n182 10.6151
R1155 B.n251 B.n182 10.6151
R1156 B.n251 B.n250 10.6151
R1157 B.n250 B.n249 10.6151
R1158 B.n249 B.n184 10.6151
R1159 B.n243 B.n184 10.6151
R1160 B.n243 B.n242 10.6151
R1161 B.n242 B.n241 10.6151
R1162 B.n241 B.n186 10.6151
R1163 B.n235 B.n186 10.6151
R1164 B.n235 B.n234 10.6151
R1165 B.n234 B.n233 10.6151
R1166 B.n233 B.n188 10.6151
R1167 B.n227 B.n188 10.6151
R1168 B.n227 B.n226 10.6151
R1169 B.n226 B.n225 10.6151
R1170 B.n225 B.n190 10.6151
R1171 B.n219 B.n190 10.6151
R1172 B.n219 B.n218 10.6151
R1173 B.n218 B.n217 10.6151
R1174 B.n217 B.n192 10.6151
R1175 B.n211 B.n192 10.6151
R1176 B.n211 B.n210 10.6151
R1177 B.n210 B.n209 10.6151
R1178 B.n209 B.n194 10.6151
R1179 B.n203 B.n194 10.6151
R1180 B.n203 B.n202 10.6151
R1181 B.n202 B.n201 10.6151
R1182 B.n201 B.n196 10.6151
R1183 B.n196 B.n154 10.6151
R1184 B.n338 B.n150 10.6151
R1185 B.n348 B.n150 10.6151
R1186 B.n349 B.n348 10.6151
R1187 B.n350 B.n349 10.6151
R1188 B.n350 B.n142 10.6151
R1189 B.n360 B.n142 10.6151
R1190 B.n361 B.n360 10.6151
R1191 B.n362 B.n361 10.6151
R1192 B.n362 B.n134 10.6151
R1193 B.n372 B.n134 10.6151
R1194 B.n373 B.n372 10.6151
R1195 B.n374 B.n373 10.6151
R1196 B.n374 B.n126 10.6151
R1197 B.n384 B.n126 10.6151
R1198 B.n385 B.n384 10.6151
R1199 B.n386 B.n385 10.6151
R1200 B.n386 B.n118 10.6151
R1201 B.n396 B.n118 10.6151
R1202 B.n397 B.n396 10.6151
R1203 B.n398 B.n397 10.6151
R1204 B.n398 B.n110 10.6151
R1205 B.n408 B.n110 10.6151
R1206 B.n409 B.n408 10.6151
R1207 B.n410 B.n409 10.6151
R1208 B.n410 B.n102 10.6151
R1209 B.n421 B.n102 10.6151
R1210 B.n422 B.n421 10.6151
R1211 B.n423 B.n422 10.6151
R1212 B.n423 B.n0 10.6151
R1213 B.n666 B.n1 10.6151
R1214 B.n666 B.n665 10.6151
R1215 B.n665 B.n664 10.6151
R1216 B.n664 B.n10 10.6151
R1217 B.n658 B.n10 10.6151
R1218 B.n658 B.n657 10.6151
R1219 B.n657 B.n656 10.6151
R1220 B.n656 B.n17 10.6151
R1221 B.n650 B.n17 10.6151
R1222 B.n650 B.n649 10.6151
R1223 B.n649 B.n648 10.6151
R1224 B.n648 B.n24 10.6151
R1225 B.n642 B.n24 10.6151
R1226 B.n642 B.n641 10.6151
R1227 B.n641 B.n640 10.6151
R1228 B.n640 B.n31 10.6151
R1229 B.n634 B.n31 10.6151
R1230 B.n634 B.n633 10.6151
R1231 B.n633 B.n632 10.6151
R1232 B.n632 B.n38 10.6151
R1233 B.n626 B.n38 10.6151
R1234 B.n626 B.n625 10.6151
R1235 B.n625 B.n624 10.6151
R1236 B.n624 B.n45 10.6151
R1237 B.n618 B.n45 10.6151
R1238 B.n618 B.n617 10.6151
R1239 B.n617 B.n616 10.6151
R1240 B.n616 B.n52 10.6151
R1241 B.n610 B.n52 10.6151
R1242 B.n419 B.t5 10.4882
R1243 B.n662 B.t6 10.4882
R1244 B.n546 B.n77 6.5566
R1245 B.n530 B.n529 6.5566
R1246 B.n276 B.n275 6.5566
R1247 B.n259 B.n258 6.5566
R1248 B.n77 B.n73 4.05904
R1249 B.n529 B.n528 4.05904
R1250 B.n277 B.n276 4.05904
R1251 B.n258 B.n257 4.05904
R1252 B.n672 B.n0 2.81026
R1253 B.n672 B.n1 2.81026
R1254 B.t4 B.n128 2.42074
R1255 B.n637 B.t1 2.42074
R1256 VP.n10 VP.t6 202.382
R1257 VP.n23 VP.n5 173.596
R1258 VP.n40 VP.n39 173.596
R1259 VP.n22 VP.n21 173.596
R1260 VP.n5 VP.t4 172.202
R1261 VP.n3 VP.t1 172.202
R1262 VP.n32 VP.t3 172.202
R1263 VP.n39 VP.t5 172.202
R1264 VP.n21 VP.t2 172.202
R1265 VP.n14 VP.t0 172.202
R1266 VP.n9 VP.t7 172.202
R1267 VP.n12 VP.n11 161.3
R1268 VP.n13 VP.n8 161.3
R1269 VP.n16 VP.n15 161.3
R1270 VP.n17 VP.n7 161.3
R1271 VP.n19 VP.n18 161.3
R1272 VP.n20 VP.n6 161.3
R1273 VP.n38 VP.n0 161.3
R1274 VP.n37 VP.n36 161.3
R1275 VP.n35 VP.n1 161.3
R1276 VP.n34 VP.n33 161.3
R1277 VP.n31 VP.n2 161.3
R1278 VP.n30 VP.n29 161.3
R1279 VP.n28 VP.n27 161.3
R1280 VP.n26 VP.n4 161.3
R1281 VP.n25 VP.n24 161.3
R1282 VP.n10 VP.n9 51.5382
R1283 VP.n23 VP.n22 41.3263
R1284 VP.n26 VP.n25 40.577
R1285 VP.n27 VP.n26 40.577
R1286 VP.n31 VP.n30 40.577
R1287 VP.n33 VP.n31 40.577
R1288 VP.n37 VP.n1 40.577
R1289 VP.n38 VP.n37 40.577
R1290 VP.n20 VP.n19 40.577
R1291 VP.n19 VP.n7 40.577
R1292 VP.n15 VP.n13 40.577
R1293 VP.n13 VP.n12 40.577
R1294 VP.n11 VP.n10 27.0073
R1295 VP.n25 VP.n5 12.2964
R1296 VP.n27 VP.n3 12.2964
R1297 VP.n30 VP.n3 12.2964
R1298 VP.n33 VP.n32 12.2964
R1299 VP.n32 VP.n1 12.2964
R1300 VP.n39 VP.n38 12.2964
R1301 VP.n21 VP.n20 12.2964
R1302 VP.n15 VP.n14 12.2964
R1303 VP.n14 VP.n7 12.2964
R1304 VP.n12 VP.n9 12.2964
R1305 VP.n11 VP.n8 0.189894
R1306 VP.n16 VP.n8 0.189894
R1307 VP.n17 VP.n16 0.189894
R1308 VP.n18 VP.n17 0.189894
R1309 VP.n18 VP.n6 0.189894
R1310 VP.n22 VP.n6 0.189894
R1311 VP.n24 VP.n23 0.189894
R1312 VP.n24 VP.n4 0.189894
R1313 VP.n28 VP.n4 0.189894
R1314 VP.n29 VP.n28 0.189894
R1315 VP.n29 VP.n2 0.189894
R1316 VP.n34 VP.n2 0.189894
R1317 VP.n35 VP.n34 0.189894
R1318 VP.n36 VP.n35 0.189894
R1319 VP.n36 VP.n0 0.189894
R1320 VP.n40 VP.n0 0.189894
R1321 VP VP.n40 0.0516364
R1322 VDD1 VDD1.n0 68.2793
R1323 VDD1.n3 VDD1.n2 68.1655
R1324 VDD1.n3 VDD1.n1 68.1655
R1325 VDD1.n5 VDD1.n4 67.5743
R1326 VDD1.n5 VDD1.n3 37.3242
R1327 VDD1.n4 VDD1.t7 2.36892
R1328 VDD1.n4 VDD1.t5 2.36892
R1329 VDD1.n0 VDD1.t1 2.36892
R1330 VDD1.n0 VDD1.t0 2.36892
R1331 VDD1.n2 VDD1.t4 2.36892
R1332 VDD1.n2 VDD1.t2 2.36892
R1333 VDD1.n1 VDD1.t3 2.36892
R1334 VDD1.n1 VDD1.t6 2.36892
R1335 VDD1 VDD1.n5 0.588862
C0 VDD2 VTAIL 7.14491f
C1 VN VP 5.23922f
C2 VDD2 VDD1 1.05764f
C3 VTAIL VP 5.0481f
C4 VDD1 VP 5.18315f
C5 VTAIL VN 5.03399f
C6 VDD1 VN 0.148933f
C7 VDD2 VP 0.367294f
C8 VDD2 VN 4.96546f
C9 VDD1 VTAIL 7.10008f
C10 VDD2 B 3.645532f
C11 VDD1 B 3.931257f
C12 VTAIL B 7.272138f
C13 VN B 9.82354f
C14 VP B 8.232537f
C15 VDD1.t1 B 0.169233f
C16 VDD1.t0 B 0.169233f
C17 VDD1.n0 B 1.47632f
C18 VDD1.t3 B 0.169233f
C19 VDD1.t6 B 0.169233f
C20 VDD1.n1 B 1.47562f
C21 VDD1.t4 B 0.169233f
C22 VDD1.t2 B 0.169233f
C23 VDD1.n2 B 1.47562f
C24 VDD1.n3 B 2.31926f
C25 VDD1.t7 B 0.169233f
C26 VDD1.t5 B 0.169233f
C27 VDD1.n4 B 1.47241f
C28 VDD1.n5 B 2.24582f
C29 VP.n0 B 0.036467f
C30 VP.t5 B 0.959747f
C31 VP.n1 B 0.055403f
C32 VP.n2 B 0.036467f
C33 VP.t1 B 0.959747f
C34 VP.n3 B 0.366585f
C35 VP.n4 B 0.036467f
C36 VP.t4 B 0.959747f
C37 VP.n5 B 0.424456f
C38 VP.n6 B 0.036467f
C39 VP.t2 B 0.959747f
C40 VP.n7 B 0.055403f
C41 VP.n8 B 0.036467f
C42 VP.t7 B 0.959747f
C43 VP.n9 B 0.419531f
C44 VP.t6 B 1.03008f
C45 VP.n10 B 0.443245f
C46 VP.n11 B 0.188763f
C47 VP.n12 B 0.055403f
C48 VP.n13 B 0.029453f
C49 VP.t0 B 0.959747f
C50 VP.n14 B 0.366585f
C51 VP.n15 B 0.055403f
C52 VP.n16 B 0.036467f
C53 VP.n17 B 0.036467f
C54 VP.n18 B 0.036467f
C55 VP.n19 B 0.029453f
C56 VP.n20 B 0.055403f
C57 VP.n21 B 0.424456f
C58 VP.n22 B 1.46935f
C59 VP.n23 B 1.50116f
C60 VP.n24 B 0.036467f
C61 VP.n25 B 0.055403f
C62 VP.n26 B 0.029453f
C63 VP.n27 B 0.055403f
C64 VP.n28 B 0.036467f
C65 VP.n29 B 0.036467f
C66 VP.n30 B 0.055403f
C67 VP.n31 B 0.029453f
C68 VP.t3 B 0.959747f
C69 VP.n32 B 0.366585f
C70 VP.n33 B 0.055403f
C71 VP.n34 B 0.036467f
C72 VP.n35 B 0.036467f
C73 VP.n36 B 0.036467f
C74 VP.n37 B 0.029453f
C75 VP.n38 B 0.055403f
C76 VP.n39 B 0.424456f
C77 VP.n40 B 0.032672f
C78 VTAIL.t13 B 0.132989f
C79 VTAIL.t14 B 0.132989f
C80 VTAIL.n0 B 1.10604f
C81 VTAIL.n1 B 0.270891f
C82 VTAIL.t10 B 1.40934f
C83 VTAIL.n2 B 0.356991f
C84 VTAIL.t5 B 1.40934f
C85 VTAIL.n3 B 0.356991f
C86 VTAIL.t3 B 0.132989f
C87 VTAIL.t2 B 0.132989f
C88 VTAIL.n4 B 1.10604f
C89 VTAIL.n5 B 0.350994f
C90 VTAIL.t4 B 1.40934f
C91 VTAIL.n6 B 1.15132f
C92 VTAIL.t15 B 1.40935f
C93 VTAIL.n7 B 1.15131f
C94 VTAIL.t9 B 0.132989f
C95 VTAIL.t11 B 0.132989f
C96 VTAIL.n8 B 1.10604f
C97 VTAIL.n9 B 0.350991f
C98 VTAIL.t12 B 1.40935f
C99 VTAIL.n10 B 0.356981f
C100 VTAIL.t6 B 1.40935f
C101 VTAIL.n11 B 0.356981f
C102 VTAIL.t0 B 0.132989f
C103 VTAIL.t7 B 0.132989f
C104 VTAIL.n12 B 1.10604f
C105 VTAIL.n13 B 0.350991f
C106 VTAIL.t1 B 1.40934f
C107 VTAIL.n14 B 1.15132f
C108 VTAIL.t8 B 1.40934f
C109 VTAIL.n15 B 1.14755f
C110 VDD2.t5 B 0.167772f
C111 VDD2.t0 B 0.167772f
C112 VDD2.n0 B 1.46288f
C113 VDD2.t1 B 0.167772f
C114 VDD2.t7 B 0.167772f
C115 VDD2.n1 B 1.46288f
C116 VDD2.n2 B 2.24525f
C117 VDD2.t3 B 0.167772f
C118 VDD2.t4 B 0.167772f
C119 VDD2.n3 B 1.4597f
C120 VDD2.n4 B 2.19613f
C121 VDD2.t6 B 0.167772f
C122 VDD2.t2 B 0.167772f
C123 VDD2.n5 B 1.46285f
C124 VN.n0 B 0.035874f
C125 VN.t7 B 0.94414f
C126 VN.n1 B 0.054502f
C127 VN.n2 B 0.035874f
C128 VN.t2 B 0.94414f
C129 VN.n3 B 0.412708f
C130 VN.t5 B 1.01333f
C131 VN.n4 B 0.436037f
C132 VN.n5 B 0.185693f
C133 VN.n6 B 0.054502f
C134 VN.n7 B 0.028974f
C135 VN.t1 B 0.94414f
C136 VN.n8 B 0.360624f
C137 VN.n9 B 0.054502f
C138 VN.n10 B 0.035874f
C139 VN.n11 B 0.035874f
C140 VN.n12 B 0.035874f
C141 VN.n13 B 0.028974f
C142 VN.n14 B 0.054502f
C143 VN.n15 B 0.417554f
C144 VN.n16 B 0.03214f
C145 VN.n17 B 0.035874f
C146 VN.t0 B 0.94414f
C147 VN.n18 B 0.054502f
C148 VN.n19 B 0.035874f
C149 VN.t6 B 0.94414f
C150 VN.n20 B 0.360624f
C151 VN.t4 B 0.94414f
C152 VN.n21 B 0.412708f
C153 VN.t3 B 1.01333f
C154 VN.n22 B 0.436037f
C155 VN.n23 B 0.185693f
C156 VN.n24 B 0.054502f
C157 VN.n25 B 0.028974f
C158 VN.n26 B 0.054502f
C159 VN.n27 B 0.035874f
C160 VN.n28 B 0.035874f
C161 VN.n29 B 0.035874f
C162 VN.n30 B 0.028974f
C163 VN.n31 B 0.054502f
C164 VN.n32 B 0.417554f
C165 VN.n33 B 1.46903f
.ends

