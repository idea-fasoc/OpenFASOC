* NGSPICE file created from diff_pair_sample_1209.ext - technology: sky130A

.subckt diff_pair_sample_1209 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X1 VTAIL.t4 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=2.7027 ps=16.71 w=16.38 l=2.31
X2 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X3 VTAIL.t14 VN.t1 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=2.7027 ps=16.71 w=16.38 l=2.31
X4 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=6.3882 ps=33.54 w=16.38 l=2.31
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=0 ps=0 w=16.38 l=2.31
X6 VDD1.t4 VP.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X7 VTAIL.t0 VP.t4 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=2.7027 ps=16.71 w=16.38 l=2.31
X8 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=6.3882 ps=33.54 w=16.38 l=2.31
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=0 ps=0 w=16.38 l=2.31
X10 VDD2.t3 VN.t2 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X11 VTAIL.t12 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=2.7027 ps=16.71 w=16.38 l=2.31
X12 VDD2.t7 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=6.3882 ps=33.54 w=16.38 l=2.31
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=0 ps=0 w=16.38 l=2.31
X14 VTAIL.t10 VN.t5 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X15 VDD1.t1 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X16 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.3882 pd=33.54 as=0 ps=0 w=16.38 l=2.31
X18 VDD2.t5 VN.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=6.3882 ps=33.54 w=16.38 l=2.31
X19 VDD2.t4 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7027 pd=16.71 as=2.7027 ps=16.71 w=16.38 l=2.31
R0 VN.n7 VN.t3 201.946
R1 VN.n34 VN.t4 201.946
R2 VN.n6 VN.t7 170.892
R3 VN.n17 VN.t5 170.892
R4 VN.n25 VN.t6 170.892
R5 VN.n33 VN.t0 170.892
R6 VN.n44 VN.t2 170.892
R7 VN.n52 VN.t1 170.892
R8 VN.n51 VN.n27 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n28 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n29 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n41 VN.n30 161.3
R15 VN.n40 VN.n39 161.3
R16 VN.n38 VN.n31 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n32 161.3
R19 VN.n24 VN.n0 161.3
R20 VN.n23 VN.n22 161.3
R21 VN.n21 VN.n1 161.3
R22 VN.n20 VN.n19 161.3
R23 VN.n18 VN.n2 161.3
R24 VN.n16 VN.n15 161.3
R25 VN.n14 VN.n3 161.3
R26 VN.n13 VN.n12 161.3
R27 VN.n11 VN.n4 161.3
R28 VN.n10 VN.n9 161.3
R29 VN.n8 VN.n5 161.3
R30 VN.n26 VN.n25 100.579
R31 VN.n53 VN.n52 100.579
R32 VN.n7 VN.n6 68.9827
R33 VN.n34 VN.n33 68.9827
R34 VN.n12 VN.n11 56.5617
R35 VN.n39 VN.n38 56.5617
R36 VN VN.n53 53.0891
R37 VN.n19 VN.n1 51.2335
R38 VN.n46 VN.n28 51.2335
R39 VN.n23 VN.n1 29.9206
R40 VN.n50 VN.n28 29.9206
R41 VN.n10 VN.n5 24.5923
R42 VN.n11 VN.n10 24.5923
R43 VN.n12 VN.n3 24.5923
R44 VN.n16 VN.n3 24.5923
R45 VN.n19 VN.n18 24.5923
R46 VN.n24 VN.n23 24.5923
R47 VN.n38 VN.n37 24.5923
R48 VN.n37 VN.n32 24.5923
R49 VN.n46 VN.n45 24.5923
R50 VN.n43 VN.n30 24.5923
R51 VN.n39 VN.n30 24.5923
R52 VN.n51 VN.n50 24.5923
R53 VN.n18 VN.n17 21.1495
R54 VN.n45 VN.n44 21.1495
R55 VN.n25 VN.n24 10.3291
R56 VN.n52 VN.n51 10.3291
R57 VN.n35 VN.n34 9.96756
R58 VN.n8 VN.n7 9.96756
R59 VN.n6 VN.n5 3.44336
R60 VN.n17 VN.n16 3.44336
R61 VN.n33 VN.n32 3.44336
R62 VN.n44 VN.n43 3.44336
R63 VN.n53 VN.n27 0.278335
R64 VN.n26 VN.n0 0.278335
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n42 VN.n29 0.189894
R70 VN.n42 VN.n41 0.189894
R71 VN.n41 VN.n40 0.189894
R72 VN.n40 VN.n31 0.189894
R73 VN.n36 VN.n31 0.189894
R74 VN.n36 VN.n35 0.189894
R75 VN.n9 VN.n8 0.189894
R76 VN.n9 VN.n4 0.189894
R77 VN.n13 VN.n4 0.189894
R78 VN.n14 VN.n13 0.189894
R79 VN.n15 VN.n14 0.189894
R80 VN.n15 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153485
R86 VDD2.n2 VDD2.n1 60.6684
R87 VDD2.n2 VDD2.n0 60.6684
R88 VDD2 VDD2.n5 60.6656
R89 VDD2.n4 VDD2.n3 59.586
R90 VDD2.n4 VDD2.n2 48.0774
R91 VDD2.n5 VDD2.t1 1.20929
R92 VDD2.n5 VDD2.t7 1.20929
R93 VDD2.n3 VDD2.t0 1.20929
R94 VDD2.n3 VDD2.t3 1.20929
R95 VDD2.n1 VDD2.t6 1.20929
R96 VDD2.n1 VDD2.t5 1.20929
R97 VDD2.n0 VDD2.t2 1.20929
R98 VDD2.n0 VDD2.t4 1.20929
R99 VDD2 VDD2.n4 1.19662
R100 VTAIL.n11 VTAIL.t0 44.116
R101 VTAIL.n10 VTAIL.t11 44.116
R102 VTAIL.n7 VTAIL.t14 44.116
R103 VTAIL.n14 VTAIL.t2 44.1158
R104 VTAIL.n15 VTAIL.t9 44.1158
R105 VTAIL.n2 VTAIL.t12 44.1158
R106 VTAIL.n3 VTAIL.t5 44.1158
R107 VTAIL.n6 VTAIL.t4 44.1158
R108 VTAIL.n13 VTAIL.n12 42.9072
R109 VTAIL.n9 VTAIL.n8 42.9072
R110 VTAIL.n1 VTAIL.n0 42.907
R111 VTAIL.n5 VTAIL.n4 42.907
R112 VTAIL.n15 VTAIL.n14 28.7634
R113 VTAIL.n7 VTAIL.n6 28.7634
R114 VTAIL.n9 VTAIL.n7 2.27636
R115 VTAIL.n10 VTAIL.n9 2.27636
R116 VTAIL.n13 VTAIL.n11 2.27636
R117 VTAIL.n14 VTAIL.n13 2.27636
R118 VTAIL.n6 VTAIL.n5 2.27636
R119 VTAIL.n5 VTAIL.n3 2.27636
R120 VTAIL.n2 VTAIL.n1 2.27636
R121 VTAIL VTAIL.n15 2.21817
R122 VTAIL.n0 VTAIL.t8 1.20929
R123 VTAIL.n0 VTAIL.t10 1.20929
R124 VTAIL.n4 VTAIL.t7 1.20929
R125 VTAIL.n4 VTAIL.t3 1.20929
R126 VTAIL.n12 VTAIL.t6 1.20929
R127 VTAIL.n12 VTAIL.t1 1.20929
R128 VTAIL.n8 VTAIL.t13 1.20929
R129 VTAIL.n8 VTAIL.t15 1.20929
R130 VTAIL.n11 VTAIL.n10 0.470328
R131 VTAIL.n3 VTAIL.n2 0.470328
R132 VTAIL VTAIL.n1 0.0586897
R133 B.n982 B.n981 585
R134 B.n983 B.n982 585
R135 B.n385 B.n147 585
R136 B.n384 B.n383 585
R137 B.n382 B.n381 585
R138 B.n380 B.n379 585
R139 B.n378 B.n377 585
R140 B.n376 B.n375 585
R141 B.n374 B.n373 585
R142 B.n372 B.n371 585
R143 B.n370 B.n369 585
R144 B.n368 B.n367 585
R145 B.n366 B.n365 585
R146 B.n364 B.n363 585
R147 B.n362 B.n361 585
R148 B.n360 B.n359 585
R149 B.n358 B.n357 585
R150 B.n356 B.n355 585
R151 B.n354 B.n353 585
R152 B.n352 B.n351 585
R153 B.n350 B.n349 585
R154 B.n348 B.n347 585
R155 B.n346 B.n345 585
R156 B.n344 B.n343 585
R157 B.n342 B.n341 585
R158 B.n340 B.n339 585
R159 B.n338 B.n337 585
R160 B.n336 B.n335 585
R161 B.n334 B.n333 585
R162 B.n332 B.n331 585
R163 B.n330 B.n329 585
R164 B.n328 B.n327 585
R165 B.n326 B.n325 585
R166 B.n324 B.n323 585
R167 B.n322 B.n321 585
R168 B.n320 B.n319 585
R169 B.n318 B.n317 585
R170 B.n316 B.n315 585
R171 B.n314 B.n313 585
R172 B.n312 B.n311 585
R173 B.n310 B.n309 585
R174 B.n308 B.n307 585
R175 B.n306 B.n305 585
R176 B.n304 B.n303 585
R177 B.n302 B.n301 585
R178 B.n300 B.n299 585
R179 B.n298 B.n297 585
R180 B.n296 B.n295 585
R181 B.n294 B.n293 585
R182 B.n292 B.n291 585
R183 B.n290 B.n289 585
R184 B.n288 B.n287 585
R185 B.n286 B.n285 585
R186 B.n284 B.n283 585
R187 B.n282 B.n281 585
R188 B.n280 B.n279 585
R189 B.n278 B.n277 585
R190 B.n276 B.n275 585
R191 B.n274 B.n273 585
R192 B.n272 B.n271 585
R193 B.n270 B.n269 585
R194 B.n268 B.n267 585
R195 B.n266 B.n265 585
R196 B.n264 B.n263 585
R197 B.n262 B.n261 585
R198 B.n259 B.n258 585
R199 B.n257 B.n256 585
R200 B.n255 B.n254 585
R201 B.n253 B.n252 585
R202 B.n251 B.n250 585
R203 B.n249 B.n248 585
R204 B.n247 B.n246 585
R205 B.n245 B.n244 585
R206 B.n243 B.n242 585
R207 B.n241 B.n240 585
R208 B.n239 B.n238 585
R209 B.n237 B.n236 585
R210 B.n235 B.n234 585
R211 B.n233 B.n232 585
R212 B.n231 B.n230 585
R213 B.n229 B.n228 585
R214 B.n227 B.n226 585
R215 B.n225 B.n224 585
R216 B.n223 B.n222 585
R217 B.n221 B.n220 585
R218 B.n219 B.n218 585
R219 B.n217 B.n216 585
R220 B.n215 B.n214 585
R221 B.n213 B.n212 585
R222 B.n211 B.n210 585
R223 B.n209 B.n208 585
R224 B.n207 B.n206 585
R225 B.n205 B.n204 585
R226 B.n203 B.n202 585
R227 B.n201 B.n200 585
R228 B.n199 B.n198 585
R229 B.n197 B.n196 585
R230 B.n195 B.n194 585
R231 B.n193 B.n192 585
R232 B.n191 B.n190 585
R233 B.n189 B.n188 585
R234 B.n187 B.n186 585
R235 B.n185 B.n184 585
R236 B.n183 B.n182 585
R237 B.n181 B.n180 585
R238 B.n179 B.n178 585
R239 B.n177 B.n176 585
R240 B.n175 B.n174 585
R241 B.n173 B.n172 585
R242 B.n171 B.n170 585
R243 B.n169 B.n168 585
R244 B.n167 B.n166 585
R245 B.n165 B.n164 585
R246 B.n163 B.n162 585
R247 B.n161 B.n160 585
R248 B.n159 B.n158 585
R249 B.n157 B.n156 585
R250 B.n155 B.n154 585
R251 B.n88 B.n87 585
R252 B.n986 B.n985 585
R253 B.n980 B.n148 585
R254 B.n148 B.n85 585
R255 B.n979 B.n84 585
R256 B.n990 B.n84 585
R257 B.n978 B.n83 585
R258 B.n991 B.n83 585
R259 B.n977 B.n82 585
R260 B.n992 B.n82 585
R261 B.n976 B.n975 585
R262 B.n975 B.n78 585
R263 B.n974 B.n77 585
R264 B.n998 B.n77 585
R265 B.n973 B.n76 585
R266 B.n999 B.n76 585
R267 B.n972 B.n75 585
R268 B.n1000 B.n75 585
R269 B.n971 B.n970 585
R270 B.n970 B.n71 585
R271 B.n969 B.n70 585
R272 B.n1006 B.n70 585
R273 B.n968 B.n69 585
R274 B.n1007 B.n69 585
R275 B.n967 B.n68 585
R276 B.n1008 B.n68 585
R277 B.n966 B.n965 585
R278 B.n965 B.n64 585
R279 B.n964 B.n63 585
R280 B.n1014 B.n63 585
R281 B.n963 B.n62 585
R282 B.n1015 B.n62 585
R283 B.n962 B.n61 585
R284 B.n1016 B.n61 585
R285 B.n961 B.n960 585
R286 B.n960 B.n57 585
R287 B.n959 B.n56 585
R288 B.n1022 B.n56 585
R289 B.n958 B.n55 585
R290 B.n1023 B.n55 585
R291 B.n957 B.n54 585
R292 B.n1024 B.n54 585
R293 B.n956 B.n955 585
R294 B.n955 B.n50 585
R295 B.n954 B.n49 585
R296 B.n1030 B.n49 585
R297 B.n953 B.n48 585
R298 B.n1031 B.n48 585
R299 B.n952 B.n47 585
R300 B.n1032 B.n47 585
R301 B.n951 B.n950 585
R302 B.n950 B.n43 585
R303 B.n949 B.n42 585
R304 B.n1038 B.n42 585
R305 B.n948 B.n41 585
R306 B.n1039 B.n41 585
R307 B.n947 B.n40 585
R308 B.n1040 B.n40 585
R309 B.n946 B.n945 585
R310 B.n945 B.n36 585
R311 B.n944 B.n35 585
R312 B.n1046 B.n35 585
R313 B.n943 B.n34 585
R314 B.n1047 B.n34 585
R315 B.n942 B.n33 585
R316 B.n1048 B.n33 585
R317 B.n941 B.n940 585
R318 B.n940 B.n29 585
R319 B.n939 B.n28 585
R320 B.n1054 B.n28 585
R321 B.n938 B.n27 585
R322 B.n1055 B.n27 585
R323 B.n937 B.n26 585
R324 B.n1056 B.n26 585
R325 B.n936 B.n935 585
R326 B.n935 B.n22 585
R327 B.n934 B.n21 585
R328 B.n1062 B.n21 585
R329 B.n933 B.n20 585
R330 B.n1063 B.n20 585
R331 B.n932 B.n19 585
R332 B.n1064 B.n19 585
R333 B.n931 B.n930 585
R334 B.n930 B.n15 585
R335 B.n929 B.n14 585
R336 B.n1070 B.n14 585
R337 B.n928 B.n13 585
R338 B.n1071 B.n13 585
R339 B.n927 B.n12 585
R340 B.n1072 B.n12 585
R341 B.n926 B.n925 585
R342 B.n925 B.n8 585
R343 B.n924 B.n7 585
R344 B.n1078 B.n7 585
R345 B.n923 B.n6 585
R346 B.n1079 B.n6 585
R347 B.n922 B.n5 585
R348 B.n1080 B.n5 585
R349 B.n921 B.n920 585
R350 B.n920 B.n4 585
R351 B.n919 B.n386 585
R352 B.n919 B.n918 585
R353 B.n909 B.n387 585
R354 B.n388 B.n387 585
R355 B.n911 B.n910 585
R356 B.n912 B.n911 585
R357 B.n908 B.n393 585
R358 B.n393 B.n392 585
R359 B.n907 B.n906 585
R360 B.n906 B.n905 585
R361 B.n395 B.n394 585
R362 B.n396 B.n395 585
R363 B.n898 B.n897 585
R364 B.n899 B.n898 585
R365 B.n896 B.n401 585
R366 B.n401 B.n400 585
R367 B.n895 B.n894 585
R368 B.n894 B.n893 585
R369 B.n403 B.n402 585
R370 B.n404 B.n403 585
R371 B.n886 B.n885 585
R372 B.n887 B.n886 585
R373 B.n884 B.n409 585
R374 B.n409 B.n408 585
R375 B.n883 B.n882 585
R376 B.n882 B.n881 585
R377 B.n411 B.n410 585
R378 B.n412 B.n411 585
R379 B.n874 B.n873 585
R380 B.n875 B.n874 585
R381 B.n872 B.n417 585
R382 B.n417 B.n416 585
R383 B.n871 B.n870 585
R384 B.n870 B.n869 585
R385 B.n419 B.n418 585
R386 B.n420 B.n419 585
R387 B.n862 B.n861 585
R388 B.n863 B.n862 585
R389 B.n860 B.n425 585
R390 B.n425 B.n424 585
R391 B.n859 B.n858 585
R392 B.n858 B.n857 585
R393 B.n427 B.n426 585
R394 B.n428 B.n427 585
R395 B.n850 B.n849 585
R396 B.n851 B.n850 585
R397 B.n848 B.n433 585
R398 B.n433 B.n432 585
R399 B.n847 B.n846 585
R400 B.n846 B.n845 585
R401 B.n435 B.n434 585
R402 B.n436 B.n435 585
R403 B.n838 B.n837 585
R404 B.n839 B.n838 585
R405 B.n836 B.n440 585
R406 B.n444 B.n440 585
R407 B.n835 B.n834 585
R408 B.n834 B.n833 585
R409 B.n442 B.n441 585
R410 B.n443 B.n442 585
R411 B.n826 B.n825 585
R412 B.n827 B.n826 585
R413 B.n824 B.n449 585
R414 B.n449 B.n448 585
R415 B.n823 B.n822 585
R416 B.n822 B.n821 585
R417 B.n451 B.n450 585
R418 B.n452 B.n451 585
R419 B.n814 B.n813 585
R420 B.n815 B.n814 585
R421 B.n812 B.n457 585
R422 B.n457 B.n456 585
R423 B.n811 B.n810 585
R424 B.n810 B.n809 585
R425 B.n459 B.n458 585
R426 B.n460 B.n459 585
R427 B.n802 B.n801 585
R428 B.n803 B.n802 585
R429 B.n800 B.n465 585
R430 B.n465 B.n464 585
R431 B.n799 B.n798 585
R432 B.n798 B.n797 585
R433 B.n467 B.n466 585
R434 B.n468 B.n467 585
R435 B.n790 B.n789 585
R436 B.n791 B.n790 585
R437 B.n788 B.n473 585
R438 B.n473 B.n472 585
R439 B.n787 B.n786 585
R440 B.n786 B.n785 585
R441 B.n475 B.n474 585
R442 B.n476 B.n475 585
R443 B.n781 B.n780 585
R444 B.n479 B.n478 585
R445 B.n777 B.n776 585
R446 B.n778 B.n777 585
R447 B.n775 B.n538 585
R448 B.n774 B.n773 585
R449 B.n772 B.n771 585
R450 B.n770 B.n769 585
R451 B.n768 B.n767 585
R452 B.n766 B.n765 585
R453 B.n764 B.n763 585
R454 B.n762 B.n761 585
R455 B.n760 B.n759 585
R456 B.n758 B.n757 585
R457 B.n756 B.n755 585
R458 B.n754 B.n753 585
R459 B.n752 B.n751 585
R460 B.n750 B.n749 585
R461 B.n748 B.n747 585
R462 B.n746 B.n745 585
R463 B.n744 B.n743 585
R464 B.n742 B.n741 585
R465 B.n740 B.n739 585
R466 B.n738 B.n737 585
R467 B.n736 B.n735 585
R468 B.n734 B.n733 585
R469 B.n732 B.n731 585
R470 B.n730 B.n729 585
R471 B.n728 B.n727 585
R472 B.n726 B.n725 585
R473 B.n724 B.n723 585
R474 B.n722 B.n721 585
R475 B.n720 B.n719 585
R476 B.n718 B.n717 585
R477 B.n716 B.n715 585
R478 B.n714 B.n713 585
R479 B.n712 B.n711 585
R480 B.n710 B.n709 585
R481 B.n708 B.n707 585
R482 B.n706 B.n705 585
R483 B.n704 B.n703 585
R484 B.n702 B.n701 585
R485 B.n700 B.n699 585
R486 B.n698 B.n697 585
R487 B.n696 B.n695 585
R488 B.n694 B.n693 585
R489 B.n692 B.n691 585
R490 B.n690 B.n689 585
R491 B.n688 B.n687 585
R492 B.n686 B.n685 585
R493 B.n684 B.n683 585
R494 B.n682 B.n681 585
R495 B.n680 B.n679 585
R496 B.n678 B.n677 585
R497 B.n676 B.n675 585
R498 B.n674 B.n673 585
R499 B.n672 B.n671 585
R500 B.n670 B.n669 585
R501 B.n668 B.n667 585
R502 B.n666 B.n665 585
R503 B.n664 B.n663 585
R504 B.n662 B.n661 585
R505 B.n660 B.n659 585
R506 B.n658 B.n657 585
R507 B.n656 B.n655 585
R508 B.n653 B.n652 585
R509 B.n651 B.n650 585
R510 B.n649 B.n648 585
R511 B.n647 B.n646 585
R512 B.n645 B.n644 585
R513 B.n643 B.n642 585
R514 B.n641 B.n640 585
R515 B.n639 B.n638 585
R516 B.n637 B.n636 585
R517 B.n635 B.n634 585
R518 B.n633 B.n632 585
R519 B.n631 B.n630 585
R520 B.n629 B.n628 585
R521 B.n627 B.n626 585
R522 B.n625 B.n624 585
R523 B.n623 B.n622 585
R524 B.n621 B.n620 585
R525 B.n619 B.n618 585
R526 B.n617 B.n616 585
R527 B.n615 B.n614 585
R528 B.n613 B.n612 585
R529 B.n611 B.n610 585
R530 B.n609 B.n608 585
R531 B.n607 B.n606 585
R532 B.n605 B.n604 585
R533 B.n603 B.n602 585
R534 B.n601 B.n600 585
R535 B.n599 B.n598 585
R536 B.n597 B.n596 585
R537 B.n595 B.n594 585
R538 B.n593 B.n592 585
R539 B.n591 B.n590 585
R540 B.n589 B.n588 585
R541 B.n587 B.n586 585
R542 B.n585 B.n584 585
R543 B.n583 B.n582 585
R544 B.n581 B.n580 585
R545 B.n579 B.n578 585
R546 B.n577 B.n576 585
R547 B.n575 B.n574 585
R548 B.n573 B.n572 585
R549 B.n571 B.n570 585
R550 B.n569 B.n568 585
R551 B.n567 B.n566 585
R552 B.n565 B.n564 585
R553 B.n563 B.n562 585
R554 B.n561 B.n560 585
R555 B.n559 B.n558 585
R556 B.n557 B.n556 585
R557 B.n555 B.n554 585
R558 B.n553 B.n552 585
R559 B.n551 B.n550 585
R560 B.n549 B.n548 585
R561 B.n547 B.n546 585
R562 B.n545 B.n544 585
R563 B.n782 B.n477 585
R564 B.n477 B.n476 585
R565 B.n784 B.n783 585
R566 B.n785 B.n784 585
R567 B.n471 B.n470 585
R568 B.n472 B.n471 585
R569 B.n793 B.n792 585
R570 B.n792 B.n791 585
R571 B.n794 B.n469 585
R572 B.n469 B.n468 585
R573 B.n796 B.n795 585
R574 B.n797 B.n796 585
R575 B.n463 B.n462 585
R576 B.n464 B.n463 585
R577 B.n805 B.n804 585
R578 B.n804 B.n803 585
R579 B.n806 B.n461 585
R580 B.n461 B.n460 585
R581 B.n808 B.n807 585
R582 B.n809 B.n808 585
R583 B.n455 B.n454 585
R584 B.n456 B.n455 585
R585 B.n817 B.n816 585
R586 B.n816 B.n815 585
R587 B.n818 B.n453 585
R588 B.n453 B.n452 585
R589 B.n820 B.n819 585
R590 B.n821 B.n820 585
R591 B.n447 B.n446 585
R592 B.n448 B.n447 585
R593 B.n829 B.n828 585
R594 B.n828 B.n827 585
R595 B.n830 B.n445 585
R596 B.n445 B.n443 585
R597 B.n832 B.n831 585
R598 B.n833 B.n832 585
R599 B.n439 B.n438 585
R600 B.n444 B.n439 585
R601 B.n841 B.n840 585
R602 B.n840 B.n839 585
R603 B.n842 B.n437 585
R604 B.n437 B.n436 585
R605 B.n844 B.n843 585
R606 B.n845 B.n844 585
R607 B.n431 B.n430 585
R608 B.n432 B.n431 585
R609 B.n853 B.n852 585
R610 B.n852 B.n851 585
R611 B.n854 B.n429 585
R612 B.n429 B.n428 585
R613 B.n856 B.n855 585
R614 B.n857 B.n856 585
R615 B.n423 B.n422 585
R616 B.n424 B.n423 585
R617 B.n865 B.n864 585
R618 B.n864 B.n863 585
R619 B.n866 B.n421 585
R620 B.n421 B.n420 585
R621 B.n868 B.n867 585
R622 B.n869 B.n868 585
R623 B.n415 B.n414 585
R624 B.n416 B.n415 585
R625 B.n877 B.n876 585
R626 B.n876 B.n875 585
R627 B.n878 B.n413 585
R628 B.n413 B.n412 585
R629 B.n880 B.n879 585
R630 B.n881 B.n880 585
R631 B.n407 B.n406 585
R632 B.n408 B.n407 585
R633 B.n889 B.n888 585
R634 B.n888 B.n887 585
R635 B.n890 B.n405 585
R636 B.n405 B.n404 585
R637 B.n892 B.n891 585
R638 B.n893 B.n892 585
R639 B.n399 B.n398 585
R640 B.n400 B.n399 585
R641 B.n901 B.n900 585
R642 B.n900 B.n899 585
R643 B.n902 B.n397 585
R644 B.n397 B.n396 585
R645 B.n904 B.n903 585
R646 B.n905 B.n904 585
R647 B.n391 B.n390 585
R648 B.n392 B.n391 585
R649 B.n914 B.n913 585
R650 B.n913 B.n912 585
R651 B.n915 B.n389 585
R652 B.n389 B.n388 585
R653 B.n917 B.n916 585
R654 B.n918 B.n917 585
R655 B.n2 B.n0 585
R656 B.n4 B.n2 585
R657 B.n3 B.n1 585
R658 B.n1079 B.n3 585
R659 B.n1077 B.n1076 585
R660 B.n1078 B.n1077 585
R661 B.n1075 B.n9 585
R662 B.n9 B.n8 585
R663 B.n1074 B.n1073 585
R664 B.n1073 B.n1072 585
R665 B.n11 B.n10 585
R666 B.n1071 B.n11 585
R667 B.n1069 B.n1068 585
R668 B.n1070 B.n1069 585
R669 B.n1067 B.n16 585
R670 B.n16 B.n15 585
R671 B.n1066 B.n1065 585
R672 B.n1065 B.n1064 585
R673 B.n18 B.n17 585
R674 B.n1063 B.n18 585
R675 B.n1061 B.n1060 585
R676 B.n1062 B.n1061 585
R677 B.n1059 B.n23 585
R678 B.n23 B.n22 585
R679 B.n1058 B.n1057 585
R680 B.n1057 B.n1056 585
R681 B.n25 B.n24 585
R682 B.n1055 B.n25 585
R683 B.n1053 B.n1052 585
R684 B.n1054 B.n1053 585
R685 B.n1051 B.n30 585
R686 B.n30 B.n29 585
R687 B.n1050 B.n1049 585
R688 B.n1049 B.n1048 585
R689 B.n32 B.n31 585
R690 B.n1047 B.n32 585
R691 B.n1045 B.n1044 585
R692 B.n1046 B.n1045 585
R693 B.n1043 B.n37 585
R694 B.n37 B.n36 585
R695 B.n1042 B.n1041 585
R696 B.n1041 B.n1040 585
R697 B.n39 B.n38 585
R698 B.n1039 B.n39 585
R699 B.n1037 B.n1036 585
R700 B.n1038 B.n1037 585
R701 B.n1035 B.n44 585
R702 B.n44 B.n43 585
R703 B.n1034 B.n1033 585
R704 B.n1033 B.n1032 585
R705 B.n46 B.n45 585
R706 B.n1031 B.n46 585
R707 B.n1029 B.n1028 585
R708 B.n1030 B.n1029 585
R709 B.n1027 B.n51 585
R710 B.n51 B.n50 585
R711 B.n1026 B.n1025 585
R712 B.n1025 B.n1024 585
R713 B.n53 B.n52 585
R714 B.n1023 B.n53 585
R715 B.n1021 B.n1020 585
R716 B.n1022 B.n1021 585
R717 B.n1019 B.n58 585
R718 B.n58 B.n57 585
R719 B.n1018 B.n1017 585
R720 B.n1017 B.n1016 585
R721 B.n60 B.n59 585
R722 B.n1015 B.n60 585
R723 B.n1013 B.n1012 585
R724 B.n1014 B.n1013 585
R725 B.n1011 B.n65 585
R726 B.n65 B.n64 585
R727 B.n1010 B.n1009 585
R728 B.n1009 B.n1008 585
R729 B.n67 B.n66 585
R730 B.n1007 B.n67 585
R731 B.n1005 B.n1004 585
R732 B.n1006 B.n1005 585
R733 B.n1003 B.n72 585
R734 B.n72 B.n71 585
R735 B.n1002 B.n1001 585
R736 B.n1001 B.n1000 585
R737 B.n74 B.n73 585
R738 B.n999 B.n74 585
R739 B.n997 B.n996 585
R740 B.n998 B.n997 585
R741 B.n995 B.n79 585
R742 B.n79 B.n78 585
R743 B.n994 B.n993 585
R744 B.n993 B.n992 585
R745 B.n81 B.n80 585
R746 B.n991 B.n81 585
R747 B.n989 B.n988 585
R748 B.n990 B.n989 585
R749 B.n987 B.n86 585
R750 B.n86 B.n85 585
R751 B.n1082 B.n1081 585
R752 B.n1081 B.n1080 585
R753 B.n780 B.n477 454.062
R754 B.n985 B.n86 454.062
R755 B.n544 B.n475 454.062
R756 B.n982 B.n148 454.062
R757 B.n542 B.t19 378.454
R758 B.n539 B.t8 378.454
R759 B.n152 B.t16 378.454
R760 B.n149 B.t12 378.454
R761 B.n983 B.n146 256.663
R762 B.n983 B.n145 256.663
R763 B.n983 B.n144 256.663
R764 B.n983 B.n143 256.663
R765 B.n983 B.n142 256.663
R766 B.n983 B.n141 256.663
R767 B.n983 B.n140 256.663
R768 B.n983 B.n139 256.663
R769 B.n983 B.n138 256.663
R770 B.n983 B.n137 256.663
R771 B.n983 B.n136 256.663
R772 B.n983 B.n135 256.663
R773 B.n983 B.n134 256.663
R774 B.n983 B.n133 256.663
R775 B.n983 B.n132 256.663
R776 B.n983 B.n131 256.663
R777 B.n983 B.n130 256.663
R778 B.n983 B.n129 256.663
R779 B.n983 B.n128 256.663
R780 B.n983 B.n127 256.663
R781 B.n983 B.n126 256.663
R782 B.n983 B.n125 256.663
R783 B.n983 B.n124 256.663
R784 B.n983 B.n123 256.663
R785 B.n983 B.n122 256.663
R786 B.n983 B.n121 256.663
R787 B.n983 B.n120 256.663
R788 B.n983 B.n119 256.663
R789 B.n983 B.n118 256.663
R790 B.n983 B.n117 256.663
R791 B.n983 B.n116 256.663
R792 B.n983 B.n115 256.663
R793 B.n983 B.n114 256.663
R794 B.n983 B.n113 256.663
R795 B.n983 B.n112 256.663
R796 B.n983 B.n111 256.663
R797 B.n983 B.n110 256.663
R798 B.n983 B.n109 256.663
R799 B.n983 B.n108 256.663
R800 B.n983 B.n107 256.663
R801 B.n983 B.n106 256.663
R802 B.n983 B.n105 256.663
R803 B.n983 B.n104 256.663
R804 B.n983 B.n103 256.663
R805 B.n983 B.n102 256.663
R806 B.n983 B.n101 256.663
R807 B.n983 B.n100 256.663
R808 B.n983 B.n99 256.663
R809 B.n983 B.n98 256.663
R810 B.n983 B.n97 256.663
R811 B.n983 B.n96 256.663
R812 B.n983 B.n95 256.663
R813 B.n983 B.n94 256.663
R814 B.n983 B.n93 256.663
R815 B.n983 B.n92 256.663
R816 B.n983 B.n91 256.663
R817 B.n983 B.n90 256.663
R818 B.n983 B.n89 256.663
R819 B.n984 B.n983 256.663
R820 B.n779 B.n778 256.663
R821 B.n778 B.n480 256.663
R822 B.n778 B.n481 256.663
R823 B.n778 B.n482 256.663
R824 B.n778 B.n483 256.663
R825 B.n778 B.n484 256.663
R826 B.n778 B.n485 256.663
R827 B.n778 B.n486 256.663
R828 B.n778 B.n487 256.663
R829 B.n778 B.n488 256.663
R830 B.n778 B.n489 256.663
R831 B.n778 B.n490 256.663
R832 B.n778 B.n491 256.663
R833 B.n778 B.n492 256.663
R834 B.n778 B.n493 256.663
R835 B.n778 B.n494 256.663
R836 B.n778 B.n495 256.663
R837 B.n778 B.n496 256.663
R838 B.n778 B.n497 256.663
R839 B.n778 B.n498 256.663
R840 B.n778 B.n499 256.663
R841 B.n778 B.n500 256.663
R842 B.n778 B.n501 256.663
R843 B.n778 B.n502 256.663
R844 B.n778 B.n503 256.663
R845 B.n778 B.n504 256.663
R846 B.n778 B.n505 256.663
R847 B.n778 B.n506 256.663
R848 B.n778 B.n507 256.663
R849 B.n778 B.n508 256.663
R850 B.n778 B.n509 256.663
R851 B.n778 B.n510 256.663
R852 B.n778 B.n511 256.663
R853 B.n778 B.n512 256.663
R854 B.n778 B.n513 256.663
R855 B.n778 B.n514 256.663
R856 B.n778 B.n515 256.663
R857 B.n778 B.n516 256.663
R858 B.n778 B.n517 256.663
R859 B.n778 B.n518 256.663
R860 B.n778 B.n519 256.663
R861 B.n778 B.n520 256.663
R862 B.n778 B.n521 256.663
R863 B.n778 B.n522 256.663
R864 B.n778 B.n523 256.663
R865 B.n778 B.n524 256.663
R866 B.n778 B.n525 256.663
R867 B.n778 B.n526 256.663
R868 B.n778 B.n527 256.663
R869 B.n778 B.n528 256.663
R870 B.n778 B.n529 256.663
R871 B.n778 B.n530 256.663
R872 B.n778 B.n531 256.663
R873 B.n778 B.n532 256.663
R874 B.n778 B.n533 256.663
R875 B.n778 B.n534 256.663
R876 B.n778 B.n535 256.663
R877 B.n778 B.n536 256.663
R878 B.n778 B.n537 256.663
R879 B.n784 B.n477 163.367
R880 B.n784 B.n471 163.367
R881 B.n792 B.n471 163.367
R882 B.n792 B.n469 163.367
R883 B.n796 B.n469 163.367
R884 B.n796 B.n463 163.367
R885 B.n804 B.n463 163.367
R886 B.n804 B.n461 163.367
R887 B.n808 B.n461 163.367
R888 B.n808 B.n455 163.367
R889 B.n816 B.n455 163.367
R890 B.n816 B.n453 163.367
R891 B.n820 B.n453 163.367
R892 B.n820 B.n447 163.367
R893 B.n828 B.n447 163.367
R894 B.n828 B.n445 163.367
R895 B.n832 B.n445 163.367
R896 B.n832 B.n439 163.367
R897 B.n840 B.n439 163.367
R898 B.n840 B.n437 163.367
R899 B.n844 B.n437 163.367
R900 B.n844 B.n431 163.367
R901 B.n852 B.n431 163.367
R902 B.n852 B.n429 163.367
R903 B.n856 B.n429 163.367
R904 B.n856 B.n423 163.367
R905 B.n864 B.n423 163.367
R906 B.n864 B.n421 163.367
R907 B.n868 B.n421 163.367
R908 B.n868 B.n415 163.367
R909 B.n876 B.n415 163.367
R910 B.n876 B.n413 163.367
R911 B.n880 B.n413 163.367
R912 B.n880 B.n407 163.367
R913 B.n888 B.n407 163.367
R914 B.n888 B.n405 163.367
R915 B.n892 B.n405 163.367
R916 B.n892 B.n399 163.367
R917 B.n900 B.n399 163.367
R918 B.n900 B.n397 163.367
R919 B.n904 B.n397 163.367
R920 B.n904 B.n391 163.367
R921 B.n913 B.n391 163.367
R922 B.n913 B.n389 163.367
R923 B.n917 B.n389 163.367
R924 B.n917 B.n2 163.367
R925 B.n1081 B.n2 163.367
R926 B.n1081 B.n3 163.367
R927 B.n1077 B.n3 163.367
R928 B.n1077 B.n9 163.367
R929 B.n1073 B.n9 163.367
R930 B.n1073 B.n11 163.367
R931 B.n1069 B.n11 163.367
R932 B.n1069 B.n16 163.367
R933 B.n1065 B.n16 163.367
R934 B.n1065 B.n18 163.367
R935 B.n1061 B.n18 163.367
R936 B.n1061 B.n23 163.367
R937 B.n1057 B.n23 163.367
R938 B.n1057 B.n25 163.367
R939 B.n1053 B.n25 163.367
R940 B.n1053 B.n30 163.367
R941 B.n1049 B.n30 163.367
R942 B.n1049 B.n32 163.367
R943 B.n1045 B.n32 163.367
R944 B.n1045 B.n37 163.367
R945 B.n1041 B.n37 163.367
R946 B.n1041 B.n39 163.367
R947 B.n1037 B.n39 163.367
R948 B.n1037 B.n44 163.367
R949 B.n1033 B.n44 163.367
R950 B.n1033 B.n46 163.367
R951 B.n1029 B.n46 163.367
R952 B.n1029 B.n51 163.367
R953 B.n1025 B.n51 163.367
R954 B.n1025 B.n53 163.367
R955 B.n1021 B.n53 163.367
R956 B.n1021 B.n58 163.367
R957 B.n1017 B.n58 163.367
R958 B.n1017 B.n60 163.367
R959 B.n1013 B.n60 163.367
R960 B.n1013 B.n65 163.367
R961 B.n1009 B.n65 163.367
R962 B.n1009 B.n67 163.367
R963 B.n1005 B.n67 163.367
R964 B.n1005 B.n72 163.367
R965 B.n1001 B.n72 163.367
R966 B.n1001 B.n74 163.367
R967 B.n997 B.n74 163.367
R968 B.n997 B.n79 163.367
R969 B.n993 B.n79 163.367
R970 B.n993 B.n81 163.367
R971 B.n989 B.n81 163.367
R972 B.n989 B.n86 163.367
R973 B.n777 B.n479 163.367
R974 B.n777 B.n538 163.367
R975 B.n773 B.n772 163.367
R976 B.n769 B.n768 163.367
R977 B.n765 B.n764 163.367
R978 B.n761 B.n760 163.367
R979 B.n757 B.n756 163.367
R980 B.n753 B.n752 163.367
R981 B.n749 B.n748 163.367
R982 B.n745 B.n744 163.367
R983 B.n741 B.n740 163.367
R984 B.n737 B.n736 163.367
R985 B.n733 B.n732 163.367
R986 B.n729 B.n728 163.367
R987 B.n725 B.n724 163.367
R988 B.n721 B.n720 163.367
R989 B.n717 B.n716 163.367
R990 B.n713 B.n712 163.367
R991 B.n709 B.n708 163.367
R992 B.n705 B.n704 163.367
R993 B.n701 B.n700 163.367
R994 B.n697 B.n696 163.367
R995 B.n693 B.n692 163.367
R996 B.n689 B.n688 163.367
R997 B.n685 B.n684 163.367
R998 B.n681 B.n680 163.367
R999 B.n677 B.n676 163.367
R1000 B.n673 B.n672 163.367
R1001 B.n669 B.n668 163.367
R1002 B.n665 B.n664 163.367
R1003 B.n661 B.n660 163.367
R1004 B.n657 B.n656 163.367
R1005 B.n652 B.n651 163.367
R1006 B.n648 B.n647 163.367
R1007 B.n644 B.n643 163.367
R1008 B.n640 B.n639 163.367
R1009 B.n636 B.n635 163.367
R1010 B.n632 B.n631 163.367
R1011 B.n628 B.n627 163.367
R1012 B.n624 B.n623 163.367
R1013 B.n620 B.n619 163.367
R1014 B.n616 B.n615 163.367
R1015 B.n612 B.n611 163.367
R1016 B.n608 B.n607 163.367
R1017 B.n604 B.n603 163.367
R1018 B.n600 B.n599 163.367
R1019 B.n596 B.n595 163.367
R1020 B.n592 B.n591 163.367
R1021 B.n588 B.n587 163.367
R1022 B.n584 B.n583 163.367
R1023 B.n580 B.n579 163.367
R1024 B.n576 B.n575 163.367
R1025 B.n572 B.n571 163.367
R1026 B.n568 B.n567 163.367
R1027 B.n564 B.n563 163.367
R1028 B.n560 B.n559 163.367
R1029 B.n556 B.n555 163.367
R1030 B.n552 B.n551 163.367
R1031 B.n548 B.n547 163.367
R1032 B.n786 B.n475 163.367
R1033 B.n786 B.n473 163.367
R1034 B.n790 B.n473 163.367
R1035 B.n790 B.n467 163.367
R1036 B.n798 B.n467 163.367
R1037 B.n798 B.n465 163.367
R1038 B.n802 B.n465 163.367
R1039 B.n802 B.n459 163.367
R1040 B.n810 B.n459 163.367
R1041 B.n810 B.n457 163.367
R1042 B.n814 B.n457 163.367
R1043 B.n814 B.n451 163.367
R1044 B.n822 B.n451 163.367
R1045 B.n822 B.n449 163.367
R1046 B.n826 B.n449 163.367
R1047 B.n826 B.n442 163.367
R1048 B.n834 B.n442 163.367
R1049 B.n834 B.n440 163.367
R1050 B.n838 B.n440 163.367
R1051 B.n838 B.n435 163.367
R1052 B.n846 B.n435 163.367
R1053 B.n846 B.n433 163.367
R1054 B.n850 B.n433 163.367
R1055 B.n850 B.n427 163.367
R1056 B.n858 B.n427 163.367
R1057 B.n858 B.n425 163.367
R1058 B.n862 B.n425 163.367
R1059 B.n862 B.n419 163.367
R1060 B.n870 B.n419 163.367
R1061 B.n870 B.n417 163.367
R1062 B.n874 B.n417 163.367
R1063 B.n874 B.n411 163.367
R1064 B.n882 B.n411 163.367
R1065 B.n882 B.n409 163.367
R1066 B.n886 B.n409 163.367
R1067 B.n886 B.n403 163.367
R1068 B.n894 B.n403 163.367
R1069 B.n894 B.n401 163.367
R1070 B.n898 B.n401 163.367
R1071 B.n898 B.n395 163.367
R1072 B.n906 B.n395 163.367
R1073 B.n906 B.n393 163.367
R1074 B.n911 B.n393 163.367
R1075 B.n911 B.n387 163.367
R1076 B.n919 B.n387 163.367
R1077 B.n920 B.n919 163.367
R1078 B.n920 B.n5 163.367
R1079 B.n6 B.n5 163.367
R1080 B.n7 B.n6 163.367
R1081 B.n925 B.n7 163.367
R1082 B.n925 B.n12 163.367
R1083 B.n13 B.n12 163.367
R1084 B.n14 B.n13 163.367
R1085 B.n930 B.n14 163.367
R1086 B.n930 B.n19 163.367
R1087 B.n20 B.n19 163.367
R1088 B.n21 B.n20 163.367
R1089 B.n935 B.n21 163.367
R1090 B.n935 B.n26 163.367
R1091 B.n27 B.n26 163.367
R1092 B.n28 B.n27 163.367
R1093 B.n940 B.n28 163.367
R1094 B.n940 B.n33 163.367
R1095 B.n34 B.n33 163.367
R1096 B.n35 B.n34 163.367
R1097 B.n945 B.n35 163.367
R1098 B.n945 B.n40 163.367
R1099 B.n41 B.n40 163.367
R1100 B.n42 B.n41 163.367
R1101 B.n950 B.n42 163.367
R1102 B.n950 B.n47 163.367
R1103 B.n48 B.n47 163.367
R1104 B.n49 B.n48 163.367
R1105 B.n955 B.n49 163.367
R1106 B.n955 B.n54 163.367
R1107 B.n55 B.n54 163.367
R1108 B.n56 B.n55 163.367
R1109 B.n960 B.n56 163.367
R1110 B.n960 B.n61 163.367
R1111 B.n62 B.n61 163.367
R1112 B.n63 B.n62 163.367
R1113 B.n965 B.n63 163.367
R1114 B.n965 B.n68 163.367
R1115 B.n69 B.n68 163.367
R1116 B.n70 B.n69 163.367
R1117 B.n970 B.n70 163.367
R1118 B.n970 B.n75 163.367
R1119 B.n76 B.n75 163.367
R1120 B.n77 B.n76 163.367
R1121 B.n975 B.n77 163.367
R1122 B.n975 B.n82 163.367
R1123 B.n83 B.n82 163.367
R1124 B.n84 B.n83 163.367
R1125 B.n148 B.n84 163.367
R1126 B.n154 B.n88 163.367
R1127 B.n158 B.n157 163.367
R1128 B.n162 B.n161 163.367
R1129 B.n166 B.n165 163.367
R1130 B.n170 B.n169 163.367
R1131 B.n174 B.n173 163.367
R1132 B.n178 B.n177 163.367
R1133 B.n182 B.n181 163.367
R1134 B.n186 B.n185 163.367
R1135 B.n190 B.n189 163.367
R1136 B.n194 B.n193 163.367
R1137 B.n198 B.n197 163.367
R1138 B.n202 B.n201 163.367
R1139 B.n206 B.n205 163.367
R1140 B.n210 B.n209 163.367
R1141 B.n214 B.n213 163.367
R1142 B.n218 B.n217 163.367
R1143 B.n222 B.n221 163.367
R1144 B.n226 B.n225 163.367
R1145 B.n230 B.n229 163.367
R1146 B.n234 B.n233 163.367
R1147 B.n238 B.n237 163.367
R1148 B.n242 B.n241 163.367
R1149 B.n246 B.n245 163.367
R1150 B.n250 B.n249 163.367
R1151 B.n254 B.n253 163.367
R1152 B.n258 B.n257 163.367
R1153 B.n263 B.n262 163.367
R1154 B.n267 B.n266 163.367
R1155 B.n271 B.n270 163.367
R1156 B.n275 B.n274 163.367
R1157 B.n279 B.n278 163.367
R1158 B.n283 B.n282 163.367
R1159 B.n287 B.n286 163.367
R1160 B.n291 B.n290 163.367
R1161 B.n295 B.n294 163.367
R1162 B.n299 B.n298 163.367
R1163 B.n303 B.n302 163.367
R1164 B.n307 B.n306 163.367
R1165 B.n311 B.n310 163.367
R1166 B.n315 B.n314 163.367
R1167 B.n319 B.n318 163.367
R1168 B.n323 B.n322 163.367
R1169 B.n327 B.n326 163.367
R1170 B.n331 B.n330 163.367
R1171 B.n335 B.n334 163.367
R1172 B.n339 B.n338 163.367
R1173 B.n343 B.n342 163.367
R1174 B.n347 B.n346 163.367
R1175 B.n351 B.n350 163.367
R1176 B.n355 B.n354 163.367
R1177 B.n359 B.n358 163.367
R1178 B.n363 B.n362 163.367
R1179 B.n367 B.n366 163.367
R1180 B.n371 B.n370 163.367
R1181 B.n375 B.n374 163.367
R1182 B.n379 B.n378 163.367
R1183 B.n383 B.n382 163.367
R1184 B.n982 B.n147 163.367
R1185 B.n542 B.t21 119.719
R1186 B.n149 B.t14 119.719
R1187 B.n539 B.t11 119.698
R1188 B.n152 B.t17 119.698
R1189 B.n780 B.n779 71.676
R1190 B.n538 B.n480 71.676
R1191 B.n772 B.n481 71.676
R1192 B.n768 B.n482 71.676
R1193 B.n764 B.n483 71.676
R1194 B.n760 B.n484 71.676
R1195 B.n756 B.n485 71.676
R1196 B.n752 B.n486 71.676
R1197 B.n748 B.n487 71.676
R1198 B.n744 B.n488 71.676
R1199 B.n740 B.n489 71.676
R1200 B.n736 B.n490 71.676
R1201 B.n732 B.n491 71.676
R1202 B.n728 B.n492 71.676
R1203 B.n724 B.n493 71.676
R1204 B.n720 B.n494 71.676
R1205 B.n716 B.n495 71.676
R1206 B.n712 B.n496 71.676
R1207 B.n708 B.n497 71.676
R1208 B.n704 B.n498 71.676
R1209 B.n700 B.n499 71.676
R1210 B.n696 B.n500 71.676
R1211 B.n692 B.n501 71.676
R1212 B.n688 B.n502 71.676
R1213 B.n684 B.n503 71.676
R1214 B.n680 B.n504 71.676
R1215 B.n676 B.n505 71.676
R1216 B.n672 B.n506 71.676
R1217 B.n668 B.n507 71.676
R1218 B.n664 B.n508 71.676
R1219 B.n660 B.n509 71.676
R1220 B.n656 B.n510 71.676
R1221 B.n651 B.n511 71.676
R1222 B.n647 B.n512 71.676
R1223 B.n643 B.n513 71.676
R1224 B.n639 B.n514 71.676
R1225 B.n635 B.n515 71.676
R1226 B.n631 B.n516 71.676
R1227 B.n627 B.n517 71.676
R1228 B.n623 B.n518 71.676
R1229 B.n619 B.n519 71.676
R1230 B.n615 B.n520 71.676
R1231 B.n611 B.n521 71.676
R1232 B.n607 B.n522 71.676
R1233 B.n603 B.n523 71.676
R1234 B.n599 B.n524 71.676
R1235 B.n595 B.n525 71.676
R1236 B.n591 B.n526 71.676
R1237 B.n587 B.n527 71.676
R1238 B.n583 B.n528 71.676
R1239 B.n579 B.n529 71.676
R1240 B.n575 B.n530 71.676
R1241 B.n571 B.n531 71.676
R1242 B.n567 B.n532 71.676
R1243 B.n563 B.n533 71.676
R1244 B.n559 B.n534 71.676
R1245 B.n555 B.n535 71.676
R1246 B.n551 B.n536 71.676
R1247 B.n547 B.n537 71.676
R1248 B.n985 B.n984 71.676
R1249 B.n154 B.n89 71.676
R1250 B.n158 B.n90 71.676
R1251 B.n162 B.n91 71.676
R1252 B.n166 B.n92 71.676
R1253 B.n170 B.n93 71.676
R1254 B.n174 B.n94 71.676
R1255 B.n178 B.n95 71.676
R1256 B.n182 B.n96 71.676
R1257 B.n186 B.n97 71.676
R1258 B.n190 B.n98 71.676
R1259 B.n194 B.n99 71.676
R1260 B.n198 B.n100 71.676
R1261 B.n202 B.n101 71.676
R1262 B.n206 B.n102 71.676
R1263 B.n210 B.n103 71.676
R1264 B.n214 B.n104 71.676
R1265 B.n218 B.n105 71.676
R1266 B.n222 B.n106 71.676
R1267 B.n226 B.n107 71.676
R1268 B.n230 B.n108 71.676
R1269 B.n234 B.n109 71.676
R1270 B.n238 B.n110 71.676
R1271 B.n242 B.n111 71.676
R1272 B.n246 B.n112 71.676
R1273 B.n250 B.n113 71.676
R1274 B.n254 B.n114 71.676
R1275 B.n258 B.n115 71.676
R1276 B.n263 B.n116 71.676
R1277 B.n267 B.n117 71.676
R1278 B.n271 B.n118 71.676
R1279 B.n275 B.n119 71.676
R1280 B.n279 B.n120 71.676
R1281 B.n283 B.n121 71.676
R1282 B.n287 B.n122 71.676
R1283 B.n291 B.n123 71.676
R1284 B.n295 B.n124 71.676
R1285 B.n299 B.n125 71.676
R1286 B.n303 B.n126 71.676
R1287 B.n307 B.n127 71.676
R1288 B.n311 B.n128 71.676
R1289 B.n315 B.n129 71.676
R1290 B.n319 B.n130 71.676
R1291 B.n323 B.n131 71.676
R1292 B.n327 B.n132 71.676
R1293 B.n331 B.n133 71.676
R1294 B.n335 B.n134 71.676
R1295 B.n339 B.n135 71.676
R1296 B.n343 B.n136 71.676
R1297 B.n347 B.n137 71.676
R1298 B.n351 B.n138 71.676
R1299 B.n355 B.n139 71.676
R1300 B.n359 B.n140 71.676
R1301 B.n363 B.n141 71.676
R1302 B.n367 B.n142 71.676
R1303 B.n371 B.n143 71.676
R1304 B.n375 B.n144 71.676
R1305 B.n379 B.n145 71.676
R1306 B.n383 B.n146 71.676
R1307 B.n147 B.n146 71.676
R1308 B.n382 B.n145 71.676
R1309 B.n378 B.n144 71.676
R1310 B.n374 B.n143 71.676
R1311 B.n370 B.n142 71.676
R1312 B.n366 B.n141 71.676
R1313 B.n362 B.n140 71.676
R1314 B.n358 B.n139 71.676
R1315 B.n354 B.n138 71.676
R1316 B.n350 B.n137 71.676
R1317 B.n346 B.n136 71.676
R1318 B.n342 B.n135 71.676
R1319 B.n338 B.n134 71.676
R1320 B.n334 B.n133 71.676
R1321 B.n330 B.n132 71.676
R1322 B.n326 B.n131 71.676
R1323 B.n322 B.n130 71.676
R1324 B.n318 B.n129 71.676
R1325 B.n314 B.n128 71.676
R1326 B.n310 B.n127 71.676
R1327 B.n306 B.n126 71.676
R1328 B.n302 B.n125 71.676
R1329 B.n298 B.n124 71.676
R1330 B.n294 B.n123 71.676
R1331 B.n290 B.n122 71.676
R1332 B.n286 B.n121 71.676
R1333 B.n282 B.n120 71.676
R1334 B.n278 B.n119 71.676
R1335 B.n274 B.n118 71.676
R1336 B.n270 B.n117 71.676
R1337 B.n266 B.n116 71.676
R1338 B.n262 B.n115 71.676
R1339 B.n257 B.n114 71.676
R1340 B.n253 B.n113 71.676
R1341 B.n249 B.n112 71.676
R1342 B.n245 B.n111 71.676
R1343 B.n241 B.n110 71.676
R1344 B.n237 B.n109 71.676
R1345 B.n233 B.n108 71.676
R1346 B.n229 B.n107 71.676
R1347 B.n225 B.n106 71.676
R1348 B.n221 B.n105 71.676
R1349 B.n217 B.n104 71.676
R1350 B.n213 B.n103 71.676
R1351 B.n209 B.n102 71.676
R1352 B.n205 B.n101 71.676
R1353 B.n201 B.n100 71.676
R1354 B.n197 B.n99 71.676
R1355 B.n193 B.n98 71.676
R1356 B.n189 B.n97 71.676
R1357 B.n185 B.n96 71.676
R1358 B.n181 B.n95 71.676
R1359 B.n177 B.n94 71.676
R1360 B.n173 B.n93 71.676
R1361 B.n169 B.n92 71.676
R1362 B.n165 B.n91 71.676
R1363 B.n161 B.n90 71.676
R1364 B.n157 B.n89 71.676
R1365 B.n984 B.n88 71.676
R1366 B.n779 B.n479 71.676
R1367 B.n773 B.n480 71.676
R1368 B.n769 B.n481 71.676
R1369 B.n765 B.n482 71.676
R1370 B.n761 B.n483 71.676
R1371 B.n757 B.n484 71.676
R1372 B.n753 B.n485 71.676
R1373 B.n749 B.n486 71.676
R1374 B.n745 B.n487 71.676
R1375 B.n741 B.n488 71.676
R1376 B.n737 B.n489 71.676
R1377 B.n733 B.n490 71.676
R1378 B.n729 B.n491 71.676
R1379 B.n725 B.n492 71.676
R1380 B.n721 B.n493 71.676
R1381 B.n717 B.n494 71.676
R1382 B.n713 B.n495 71.676
R1383 B.n709 B.n496 71.676
R1384 B.n705 B.n497 71.676
R1385 B.n701 B.n498 71.676
R1386 B.n697 B.n499 71.676
R1387 B.n693 B.n500 71.676
R1388 B.n689 B.n501 71.676
R1389 B.n685 B.n502 71.676
R1390 B.n681 B.n503 71.676
R1391 B.n677 B.n504 71.676
R1392 B.n673 B.n505 71.676
R1393 B.n669 B.n506 71.676
R1394 B.n665 B.n507 71.676
R1395 B.n661 B.n508 71.676
R1396 B.n657 B.n509 71.676
R1397 B.n652 B.n510 71.676
R1398 B.n648 B.n511 71.676
R1399 B.n644 B.n512 71.676
R1400 B.n640 B.n513 71.676
R1401 B.n636 B.n514 71.676
R1402 B.n632 B.n515 71.676
R1403 B.n628 B.n516 71.676
R1404 B.n624 B.n517 71.676
R1405 B.n620 B.n518 71.676
R1406 B.n616 B.n519 71.676
R1407 B.n612 B.n520 71.676
R1408 B.n608 B.n521 71.676
R1409 B.n604 B.n522 71.676
R1410 B.n600 B.n523 71.676
R1411 B.n596 B.n524 71.676
R1412 B.n592 B.n525 71.676
R1413 B.n588 B.n526 71.676
R1414 B.n584 B.n527 71.676
R1415 B.n580 B.n528 71.676
R1416 B.n576 B.n529 71.676
R1417 B.n572 B.n530 71.676
R1418 B.n568 B.n531 71.676
R1419 B.n564 B.n532 71.676
R1420 B.n560 B.n533 71.676
R1421 B.n556 B.n534 71.676
R1422 B.n552 B.n535 71.676
R1423 B.n548 B.n536 71.676
R1424 B.n544 B.n537 71.676
R1425 B.n543 B.t20 68.5188
R1426 B.n150 B.t15 68.5188
R1427 B.n540 B.t10 68.4971
R1428 B.n153 B.t18 68.4971
R1429 B.n778 B.n476 60.4484
R1430 B.n983 B.n85 60.4484
R1431 B.n654 B.n543 59.5399
R1432 B.n541 B.n540 59.5399
R1433 B.n260 B.n153 59.5399
R1434 B.n151 B.n150 59.5399
R1435 B.n543 B.n542 51.2005
R1436 B.n540 B.n539 51.2005
R1437 B.n153 B.n152 51.2005
R1438 B.n150 B.n149 51.2005
R1439 B.n785 B.n476 34.5422
R1440 B.n785 B.n472 34.5422
R1441 B.n791 B.n472 34.5422
R1442 B.n791 B.n468 34.5422
R1443 B.n797 B.n468 34.5422
R1444 B.n797 B.n464 34.5422
R1445 B.n803 B.n464 34.5422
R1446 B.n809 B.n460 34.5422
R1447 B.n809 B.n456 34.5422
R1448 B.n815 B.n456 34.5422
R1449 B.n815 B.n452 34.5422
R1450 B.n821 B.n452 34.5422
R1451 B.n821 B.n448 34.5422
R1452 B.n827 B.n448 34.5422
R1453 B.n827 B.n443 34.5422
R1454 B.n833 B.n443 34.5422
R1455 B.n833 B.n444 34.5422
R1456 B.n839 B.n436 34.5422
R1457 B.n845 B.n436 34.5422
R1458 B.n845 B.n432 34.5422
R1459 B.n851 B.n432 34.5422
R1460 B.n851 B.n428 34.5422
R1461 B.n857 B.n428 34.5422
R1462 B.n863 B.n424 34.5422
R1463 B.n863 B.n420 34.5422
R1464 B.n869 B.n420 34.5422
R1465 B.n869 B.n416 34.5422
R1466 B.n875 B.n416 34.5422
R1467 B.n875 B.n412 34.5422
R1468 B.n881 B.n412 34.5422
R1469 B.n887 B.n408 34.5422
R1470 B.n887 B.n404 34.5422
R1471 B.n893 B.n404 34.5422
R1472 B.n893 B.n400 34.5422
R1473 B.n899 B.n400 34.5422
R1474 B.n899 B.n396 34.5422
R1475 B.n905 B.n396 34.5422
R1476 B.n912 B.n392 34.5422
R1477 B.n912 B.n388 34.5422
R1478 B.n918 B.n388 34.5422
R1479 B.n918 B.n4 34.5422
R1480 B.n1080 B.n4 34.5422
R1481 B.n1080 B.n1079 34.5422
R1482 B.n1079 B.n1078 34.5422
R1483 B.n1078 B.n8 34.5422
R1484 B.n1072 B.n8 34.5422
R1485 B.n1072 B.n1071 34.5422
R1486 B.n1070 B.n15 34.5422
R1487 B.n1064 B.n15 34.5422
R1488 B.n1064 B.n1063 34.5422
R1489 B.n1063 B.n1062 34.5422
R1490 B.n1062 B.n22 34.5422
R1491 B.n1056 B.n22 34.5422
R1492 B.n1056 B.n1055 34.5422
R1493 B.n1054 B.n29 34.5422
R1494 B.n1048 B.n29 34.5422
R1495 B.n1048 B.n1047 34.5422
R1496 B.n1047 B.n1046 34.5422
R1497 B.n1046 B.n36 34.5422
R1498 B.n1040 B.n36 34.5422
R1499 B.n1040 B.n1039 34.5422
R1500 B.n1038 B.n43 34.5422
R1501 B.n1032 B.n43 34.5422
R1502 B.n1032 B.n1031 34.5422
R1503 B.n1031 B.n1030 34.5422
R1504 B.n1030 B.n50 34.5422
R1505 B.n1024 B.n50 34.5422
R1506 B.n1023 B.n1022 34.5422
R1507 B.n1022 B.n57 34.5422
R1508 B.n1016 B.n57 34.5422
R1509 B.n1016 B.n1015 34.5422
R1510 B.n1015 B.n1014 34.5422
R1511 B.n1014 B.n64 34.5422
R1512 B.n1008 B.n64 34.5422
R1513 B.n1008 B.n1007 34.5422
R1514 B.n1007 B.n1006 34.5422
R1515 B.n1006 B.n71 34.5422
R1516 B.n1000 B.n999 34.5422
R1517 B.n999 B.n998 34.5422
R1518 B.n998 B.n78 34.5422
R1519 B.n992 B.n78 34.5422
R1520 B.n992 B.n991 34.5422
R1521 B.n991 B.n990 34.5422
R1522 B.n990 B.n85 34.5422
R1523 B.n857 B.t7 34.0342
R1524 B.t1 B.n1038 34.0342
R1525 B.n981 B.n980 29.5029
R1526 B.n987 B.n986 29.5029
R1527 B.n545 B.n474 29.5029
R1528 B.n782 B.n781 29.5029
R1529 B.n839 B.t4 26.9227
R1530 B.n1024 B.t2 26.9227
R1531 B.t9 B.n460 25.9068
R1532 B.n881 B.t3 25.9068
R1533 B.t6 B.n1054 25.9068
R1534 B.t13 B.n71 25.9068
R1535 B B.n1082 18.0485
R1536 B.n905 B.t5 17.7793
R1537 B.t0 B.n1070 17.7793
R1538 B.t5 B.n392 16.7634
R1539 B.n1071 B.t0 16.7634
R1540 B.n986 B.n87 10.6151
R1541 B.n155 B.n87 10.6151
R1542 B.n156 B.n155 10.6151
R1543 B.n159 B.n156 10.6151
R1544 B.n160 B.n159 10.6151
R1545 B.n163 B.n160 10.6151
R1546 B.n164 B.n163 10.6151
R1547 B.n167 B.n164 10.6151
R1548 B.n168 B.n167 10.6151
R1549 B.n171 B.n168 10.6151
R1550 B.n172 B.n171 10.6151
R1551 B.n175 B.n172 10.6151
R1552 B.n176 B.n175 10.6151
R1553 B.n179 B.n176 10.6151
R1554 B.n180 B.n179 10.6151
R1555 B.n183 B.n180 10.6151
R1556 B.n184 B.n183 10.6151
R1557 B.n187 B.n184 10.6151
R1558 B.n188 B.n187 10.6151
R1559 B.n191 B.n188 10.6151
R1560 B.n192 B.n191 10.6151
R1561 B.n195 B.n192 10.6151
R1562 B.n196 B.n195 10.6151
R1563 B.n199 B.n196 10.6151
R1564 B.n200 B.n199 10.6151
R1565 B.n203 B.n200 10.6151
R1566 B.n204 B.n203 10.6151
R1567 B.n207 B.n204 10.6151
R1568 B.n208 B.n207 10.6151
R1569 B.n211 B.n208 10.6151
R1570 B.n212 B.n211 10.6151
R1571 B.n215 B.n212 10.6151
R1572 B.n216 B.n215 10.6151
R1573 B.n219 B.n216 10.6151
R1574 B.n220 B.n219 10.6151
R1575 B.n223 B.n220 10.6151
R1576 B.n224 B.n223 10.6151
R1577 B.n227 B.n224 10.6151
R1578 B.n228 B.n227 10.6151
R1579 B.n231 B.n228 10.6151
R1580 B.n232 B.n231 10.6151
R1581 B.n235 B.n232 10.6151
R1582 B.n236 B.n235 10.6151
R1583 B.n239 B.n236 10.6151
R1584 B.n240 B.n239 10.6151
R1585 B.n243 B.n240 10.6151
R1586 B.n244 B.n243 10.6151
R1587 B.n247 B.n244 10.6151
R1588 B.n248 B.n247 10.6151
R1589 B.n251 B.n248 10.6151
R1590 B.n252 B.n251 10.6151
R1591 B.n255 B.n252 10.6151
R1592 B.n256 B.n255 10.6151
R1593 B.n259 B.n256 10.6151
R1594 B.n264 B.n261 10.6151
R1595 B.n265 B.n264 10.6151
R1596 B.n268 B.n265 10.6151
R1597 B.n269 B.n268 10.6151
R1598 B.n272 B.n269 10.6151
R1599 B.n273 B.n272 10.6151
R1600 B.n276 B.n273 10.6151
R1601 B.n277 B.n276 10.6151
R1602 B.n281 B.n280 10.6151
R1603 B.n284 B.n281 10.6151
R1604 B.n285 B.n284 10.6151
R1605 B.n288 B.n285 10.6151
R1606 B.n289 B.n288 10.6151
R1607 B.n292 B.n289 10.6151
R1608 B.n293 B.n292 10.6151
R1609 B.n296 B.n293 10.6151
R1610 B.n297 B.n296 10.6151
R1611 B.n300 B.n297 10.6151
R1612 B.n301 B.n300 10.6151
R1613 B.n304 B.n301 10.6151
R1614 B.n305 B.n304 10.6151
R1615 B.n308 B.n305 10.6151
R1616 B.n309 B.n308 10.6151
R1617 B.n312 B.n309 10.6151
R1618 B.n313 B.n312 10.6151
R1619 B.n316 B.n313 10.6151
R1620 B.n317 B.n316 10.6151
R1621 B.n320 B.n317 10.6151
R1622 B.n321 B.n320 10.6151
R1623 B.n324 B.n321 10.6151
R1624 B.n325 B.n324 10.6151
R1625 B.n328 B.n325 10.6151
R1626 B.n329 B.n328 10.6151
R1627 B.n332 B.n329 10.6151
R1628 B.n333 B.n332 10.6151
R1629 B.n336 B.n333 10.6151
R1630 B.n337 B.n336 10.6151
R1631 B.n340 B.n337 10.6151
R1632 B.n341 B.n340 10.6151
R1633 B.n344 B.n341 10.6151
R1634 B.n345 B.n344 10.6151
R1635 B.n348 B.n345 10.6151
R1636 B.n349 B.n348 10.6151
R1637 B.n352 B.n349 10.6151
R1638 B.n353 B.n352 10.6151
R1639 B.n356 B.n353 10.6151
R1640 B.n357 B.n356 10.6151
R1641 B.n360 B.n357 10.6151
R1642 B.n361 B.n360 10.6151
R1643 B.n364 B.n361 10.6151
R1644 B.n365 B.n364 10.6151
R1645 B.n368 B.n365 10.6151
R1646 B.n369 B.n368 10.6151
R1647 B.n372 B.n369 10.6151
R1648 B.n373 B.n372 10.6151
R1649 B.n376 B.n373 10.6151
R1650 B.n377 B.n376 10.6151
R1651 B.n380 B.n377 10.6151
R1652 B.n381 B.n380 10.6151
R1653 B.n384 B.n381 10.6151
R1654 B.n385 B.n384 10.6151
R1655 B.n981 B.n385 10.6151
R1656 B.n787 B.n474 10.6151
R1657 B.n788 B.n787 10.6151
R1658 B.n789 B.n788 10.6151
R1659 B.n789 B.n466 10.6151
R1660 B.n799 B.n466 10.6151
R1661 B.n800 B.n799 10.6151
R1662 B.n801 B.n800 10.6151
R1663 B.n801 B.n458 10.6151
R1664 B.n811 B.n458 10.6151
R1665 B.n812 B.n811 10.6151
R1666 B.n813 B.n812 10.6151
R1667 B.n813 B.n450 10.6151
R1668 B.n823 B.n450 10.6151
R1669 B.n824 B.n823 10.6151
R1670 B.n825 B.n824 10.6151
R1671 B.n825 B.n441 10.6151
R1672 B.n835 B.n441 10.6151
R1673 B.n836 B.n835 10.6151
R1674 B.n837 B.n836 10.6151
R1675 B.n837 B.n434 10.6151
R1676 B.n847 B.n434 10.6151
R1677 B.n848 B.n847 10.6151
R1678 B.n849 B.n848 10.6151
R1679 B.n849 B.n426 10.6151
R1680 B.n859 B.n426 10.6151
R1681 B.n860 B.n859 10.6151
R1682 B.n861 B.n860 10.6151
R1683 B.n861 B.n418 10.6151
R1684 B.n871 B.n418 10.6151
R1685 B.n872 B.n871 10.6151
R1686 B.n873 B.n872 10.6151
R1687 B.n873 B.n410 10.6151
R1688 B.n883 B.n410 10.6151
R1689 B.n884 B.n883 10.6151
R1690 B.n885 B.n884 10.6151
R1691 B.n885 B.n402 10.6151
R1692 B.n895 B.n402 10.6151
R1693 B.n896 B.n895 10.6151
R1694 B.n897 B.n896 10.6151
R1695 B.n897 B.n394 10.6151
R1696 B.n907 B.n394 10.6151
R1697 B.n908 B.n907 10.6151
R1698 B.n910 B.n908 10.6151
R1699 B.n910 B.n909 10.6151
R1700 B.n909 B.n386 10.6151
R1701 B.n921 B.n386 10.6151
R1702 B.n922 B.n921 10.6151
R1703 B.n923 B.n922 10.6151
R1704 B.n924 B.n923 10.6151
R1705 B.n926 B.n924 10.6151
R1706 B.n927 B.n926 10.6151
R1707 B.n928 B.n927 10.6151
R1708 B.n929 B.n928 10.6151
R1709 B.n931 B.n929 10.6151
R1710 B.n932 B.n931 10.6151
R1711 B.n933 B.n932 10.6151
R1712 B.n934 B.n933 10.6151
R1713 B.n936 B.n934 10.6151
R1714 B.n937 B.n936 10.6151
R1715 B.n938 B.n937 10.6151
R1716 B.n939 B.n938 10.6151
R1717 B.n941 B.n939 10.6151
R1718 B.n942 B.n941 10.6151
R1719 B.n943 B.n942 10.6151
R1720 B.n944 B.n943 10.6151
R1721 B.n946 B.n944 10.6151
R1722 B.n947 B.n946 10.6151
R1723 B.n948 B.n947 10.6151
R1724 B.n949 B.n948 10.6151
R1725 B.n951 B.n949 10.6151
R1726 B.n952 B.n951 10.6151
R1727 B.n953 B.n952 10.6151
R1728 B.n954 B.n953 10.6151
R1729 B.n956 B.n954 10.6151
R1730 B.n957 B.n956 10.6151
R1731 B.n958 B.n957 10.6151
R1732 B.n959 B.n958 10.6151
R1733 B.n961 B.n959 10.6151
R1734 B.n962 B.n961 10.6151
R1735 B.n963 B.n962 10.6151
R1736 B.n964 B.n963 10.6151
R1737 B.n966 B.n964 10.6151
R1738 B.n967 B.n966 10.6151
R1739 B.n968 B.n967 10.6151
R1740 B.n969 B.n968 10.6151
R1741 B.n971 B.n969 10.6151
R1742 B.n972 B.n971 10.6151
R1743 B.n973 B.n972 10.6151
R1744 B.n974 B.n973 10.6151
R1745 B.n976 B.n974 10.6151
R1746 B.n977 B.n976 10.6151
R1747 B.n978 B.n977 10.6151
R1748 B.n979 B.n978 10.6151
R1749 B.n980 B.n979 10.6151
R1750 B.n781 B.n478 10.6151
R1751 B.n776 B.n478 10.6151
R1752 B.n776 B.n775 10.6151
R1753 B.n775 B.n774 10.6151
R1754 B.n774 B.n771 10.6151
R1755 B.n771 B.n770 10.6151
R1756 B.n770 B.n767 10.6151
R1757 B.n767 B.n766 10.6151
R1758 B.n766 B.n763 10.6151
R1759 B.n763 B.n762 10.6151
R1760 B.n762 B.n759 10.6151
R1761 B.n759 B.n758 10.6151
R1762 B.n758 B.n755 10.6151
R1763 B.n755 B.n754 10.6151
R1764 B.n754 B.n751 10.6151
R1765 B.n751 B.n750 10.6151
R1766 B.n750 B.n747 10.6151
R1767 B.n747 B.n746 10.6151
R1768 B.n746 B.n743 10.6151
R1769 B.n743 B.n742 10.6151
R1770 B.n742 B.n739 10.6151
R1771 B.n739 B.n738 10.6151
R1772 B.n738 B.n735 10.6151
R1773 B.n735 B.n734 10.6151
R1774 B.n734 B.n731 10.6151
R1775 B.n731 B.n730 10.6151
R1776 B.n730 B.n727 10.6151
R1777 B.n727 B.n726 10.6151
R1778 B.n726 B.n723 10.6151
R1779 B.n723 B.n722 10.6151
R1780 B.n722 B.n719 10.6151
R1781 B.n719 B.n718 10.6151
R1782 B.n718 B.n715 10.6151
R1783 B.n715 B.n714 10.6151
R1784 B.n714 B.n711 10.6151
R1785 B.n711 B.n710 10.6151
R1786 B.n710 B.n707 10.6151
R1787 B.n707 B.n706 10.6151
R1788 B.n706 B.n703 10.6151
R1789 B.n703 B.n702 10.6151
R1790 B.n702 B.n699 10.6151
R1791 B.n699 B.n698 10.6151
R1792 B.n698 B.n695 10.6151
R1793 B.n695 B.n694 10.6151
R1794 B.n694 B.n691 10.6151
R1795 B.n691 B.n690 10.6151
R1796 B.n690 B.n687 10.6151
R1797 B.n687 B.n686 10.6151
R1798 B.n686 B.n683 10.6151
R1799 B.n683 B.n682 10.6151
R1800 B.n682 B.n679 10.6151
R1801 B.n679 B.n678 10.6151
R1802 B.n678 B.n675 10.6151
R1803 B.n675 B.n674 10.6151
R1804 B.n671 B.n670 10.6151
R1805 B.n670 B.n667 10.6151
R1806 B.n667 B.n666 10.6151
R1807 B.n666 B.n663 10.6151
R1808 B.n663 B.n662 10.6151
R1809 B.n662 B.n659 10.6151
R1810 B.n659 B.n658 10.6151
R1811 B.n658 B.n655 10.6151
R1812 B.n653 B.n650 10.6151
R1813 B.n650 B.n649 10.6151
R1814 B.n649 B.n646 10.6151
R1815 B.n646 B.n645 10.6151
R1816 B.n645 B.n642 10.6151
R1817 B.n642 B.n641 10.6151
R1818 B.n641 B.n638 10.6151
R1819 B.n638 B.n637 10.6151
R1820 B.n637 B.n634 10.6151
R1821 B.n634 B.n633 10.6151
R1822 B.n633 B.n630 10.6151
R1823 B.n630 B.n629 10.6151
R1824 B.n629 B.n626 10.6151
R1825 B.n626 B.n625 10.6151
R1826 B.n625 B.n622 10.6151
R1827 B.n622 B.n621 10.6151
R1828 B.n621 B.n618 10.6151
R1829 B.n618 B.n617 10.6151
R1830 B.n617 B.n614 10.6151
R1831 B.n614 B.n613 10.6151
R1832 B.n613 B.n610 10.6151
R1833 B.n610 B.n609 10.6151
R1834 B.n609 B.n606 10.6151
R1835 B.n606 B.n605 10.6151
R1836 B.n605 B.n602 10.6151
R1837 B.n602 B.n601 10.6151
R1838 B.n601 B.n598 10.6151
R1839 B.n598 B.n597 10.6151
R1840 B.n597 B.n594 10.6151
R1841 B.n594 B.n593 10.6151
R1842 B.n593 B.n590 10.6151
R1843 B.n590 B.n589 10.6151
R1844 B.n589 B.n586 10.6151
R1845 B.n586 B.n585 10.6151
R1846 B.n585 B.n582 10.6151
R1847 B.n582 B.n581 10.6151
R1848 B.n581 B.n578 10.6151
R1849 B.n578 B.n577 10.6151
R1850 B.n577 B.n574 10.6151
R1851 B.n574 B.n573 10.6151
R1852 B.n573 B.n570 10.6151
R1853 B.n570 B.n569 10.6151
R1854 B.n569 B.n566 10.6151
R1855 B.n566 B.n565 10.6151
R1856 B.n565 B.n562 10.6151
R1857 B.n562 B.n561 10.6151
R1858 B.n561 B.n558 10.6151
R1859 B.n558 B.n557 10.6151
R1860 B.n557 B.n554 10.6151
R1861 B.n554 B.n553 10.6151
R1862 B.n553 B.n550 10.6151
R1863 B.n550 B.n549 10.6151
R1864 B.n549 B.n546 10.6151
R1865 B.n546 B.n545 10.6151
R1866 B.n783 B.n782 10.6151
R1867 B.n783 B.n470 10.6151
R1868 B.n793 B.n470 10.6151
R1869 B.n794 B.n793 10.6151
R1870 B.n795 B.n794 10.6151
R1871 B.n795 B.n462 10.6151
R1872 B.n805 B.n462 10.6151
R1873 B.n806 B.n805 10.6151
R1874 B.n807 B.n806 10.6151
R1875 B.n807 B.n454 10.6151
R1876 B.n817 B.n454 10.6151
R1877 B.n818 B.n817 10.6151
R1878 B.n819 B.n818 10.6151
R1879 B.n819 B.n446 10.6151
R1880 B.n829 B.n446 10.6151
R1881 B.n830 B.n829 10.6151
R1882 B.n831 B.n830 10.6151
R1883 B.n831 B.n438 10.6151
R1884 B.n841 B.n438 10.6151
R1885 B.n842 B.n841 10.6151
R1886 B.n843 B.n842 10.6151
R1887 B.n843 B.n430 10.6151
R1888 B.n853 B.n430 10.6151
R1889 B.n854 B.n853 10.6151
R1890 B.n855 B.n854 10.6151
R1891 B.n855 B.n422 10.6151
R1892 B.n865 B.n422 10.6151
R1893 B.n866 B.n865 10.6151
R1894 B.n867 B.n866 10.6151
R1895 B.n867 B.n414 10.6151
R1896 B.n877 B.n414 10.6151
R1897 B.n878 B.n877 10.6151
R1898 B.n879 B.n878 10.6151
R1899 B.n879 B.n406 10.6151
R1900 B.n889 B.n406 10.6151
R1901 B.n890 B.n889 10.6151
R1902 B.n891 B.n890 10.6151
R1903 B.n891 B.n398 10.6151
R1904 B.n901 B.n398 10.6151
R1905 B.n902 B.n901 10.6151
R1906 B.n903 B.n902 10.6151
R1907 B.n903 B.n390 10.6151
R1908 B.n914 B.n390 10.6151
R1909 B.n915 B.n914 10.6151
R1910 B.n916 B.n915 10.6151
R1911 B.n916 B.n0 10.6151
R1912 B.n1076 B.n1 10.6151
R1913 B.n1076 B.n1075 10.6151
R1914 B.n1075 B.n1074 10.6151
R1915 B.n1074 B.n10 10.6151
R1916 B.n1068 B.n10 10.6151
R1917 B.n1068 B.n1067 10.6151
R1918 B.n1067 B.n1066 10.6151
R1919 B.n1066 B.n17 10.6151
R1920 B.n1060 B.n17 10.6151
R1921 B.n1060 B.n1059 10.6151
R1922 B.n1059 B.n1058 10.6151
R1923 B.n1058 B.n24 10.6151
R1924 B.n1052 B.n24 10.6151
R1925 B.n1052 B.n1051 10.6151
R1926 B.n1051 B.n1050 10.6151
R1927 B.n1050 B.n31 10.6151
R1928 B.n1044 B.n31 10.6151
R1929 B.n1044 B.n1043 10.6151
R1930 B.n1043 B.n1042 10.6151
R1931 B.n1042 B.n38 10.6151
R1932 B.n1036 B.n38 10.6151
R1933 B.n1036 B.n1035 10.6151
R1934 B.n1035 B.n1034 10.6151
R1935 B.n1034 B.n45 10.6151
R1936 B.n1028 B.n45 10.6151
R1937 B.n1028 B.n1027 10.6151
R1938 B.n1027 B.n1026 10.6151
R1939 B.n1026 B.n52 10.6151
R1940 B.n1020 B.n52 10.6151
R1941 B.n1020 B.n1019 10.6151
R1942 B.n1019 B.n1018 10.6151
R1943 B.n1018 B.n59 10.6151
R1944 B.n1012 B.n59 10.6151
R1945 B.n1012 B.n1011 10.6151
R1946 B.n1011 B.n1010 10.6151
R1947 B.n1010 B.n66 10.6151
R1948 B.n1004 B.n66 10.6151
R1949 B.n1004 B.n1003 10.6151
R1950 B.n1003 B.n1002 10.6151
R1951 B.n1002 B.n73 10.6151
R1952 B.n996 B.n73 10.6151
R1953 B.n996 B.n995 10.6151
R1954 B.n995 B.n994 10.6151
R1955 B.n994 B.n80 10.6151
R1956 B.n988 B.n80 10.6151
R1957 B.n988 B.n987 10.6151
R1958 B.n803 B.t9 8.63592
R1959 B.t3 B.n408 8.63592
R1960 B.n1055 B.t6 8.63592
R1961 B.n1000 B.t13 8.63592
R1962 B.n444 B.t4 7.61999
R1963 B.t2 B.n1023 7.61999
R1964 B.n261 B.n260 6.5566
R1965 B.n277 B.n151 6.5566
R1966 B.n671 B.n541 6.5566
R1967 B.n655 B.n654 6.5566
R1968 B.n260 B.n259 4.05904
R1969 B.n280 B.n151 4.05904
R1970 B.n674 B.n541 4.05904
R1971 B.n654 B.n653 4.05904
R1972 B.n1082 B.n0 2.81026
R1973 B.n1082 B.n1 2.81026
R1974 B.t7 B.n424 0.508466
R1975 B.n1039 B.t1 0.508466
R1976 VP.n15 VP.t4 201.946
R1977 VP.n36 VP.t0 170.892
R1978 VP.n43 VP.t3 170.892
R1979 VP.n55 VP.t7 170.892
R1980 VP.n63 VP.t5 170.892
R1981 VP.n33 VP.t2 170.892
R1982 VP.n25 VP.t1 170.892
R1983 VP.n14 VP.t6 170.892
R1984 VP.n16 VP.n13 161.3
R1985 VP.n18 VP.n17 161.3
R1986 VP.n19 VP.n12 161.3
R1987 VP.n21 VP.n20 161.3
R1988 VP.n22 VP.n11 161.3
R1989 VP.n24 VP.n23 161.3
R1990 VP.n26 VP.n10 161.3
R1991 VP.n28 VP.n27 161.3
R1992 VP.n29 VP.n9 161.3
R1993 VP.n31 VP.n30 161.3
R1994 VP.n32 VP.n8 161.3
R1995 VP.n62 VP.n0 161.3
R1996 VP.n61 VP.n60 161.3
R1997 VP.n59 VP.n1 161.3
R1998 VP.n58 VP.n57 161.3
R1999 VP.n56 VP.n2 161.3
R2000 VP.n54 VP.n53 161.3
R2001 VP.n52 VP.n3 161.3
R2002 VP.n51 VP.n50 161.3
R2003 VP.n49 VP.n4 161.3
R2004 VP.n48 VP.n47 161.3
R2005 VP.n46 VP.n5 161.3
R2006 VP.n45 VP.n44 161.3
R2007 VP.n42 VP.n6 161.3
R2008 VP.n41 VP.n40 161.3
R2009 VP.n39 VP.n7 161.3
R2010 VP.n38 VP.n37 161.3
R2011 VP.n36 VP.n35 100.579
R2012 VP.n64 VP.n63 100.579
R2013 VP.n34 VP.n33 100.579
R2014 VP.n15 VP.n14 68.9827
R2015 VP.n50 VP.n49 56.5617
R2016 VP.n20 VP.n19 56.5617
R2017 VP.n35 VP.n34 52.8103
R2018 VP.n42 VP.n41 51.2335
R2019 VP.n57 VP.n1 51.2335
R2020 VP.n27 VP.n9 51.2335
R2021 VP.n41 VP.n7 29.9206
R2022 VP.n61 VP.n1 29.9206
R2023 VP.n31 VP.n9 29.9206
R2024 VP.n37 VP.n7 24.5923
R2025 VP.n44 VP.n42 24.5923
R2026 VP.n48 VP.n5 24.5923
R2027 VP.n49 VP.n48 24.5923
R2028 VP.n50 VP.n3 24.5923
R2029 VP.n54 VP.n3 24.5923
R2030 VP.n57 VP.n56 24.5923
R2031 VP.n62 VP.n61 24.5923
R2032 VP.n32 VP.n31 24.5923
R2033 VP.n20 VP.n11 24.5923
R2034 VP.n24 VP.n11 24.5923
R2035 VP.n27 VP.n26 24.5923
R2036 VP.n18 VP.n13 24.5923
R2037 VP.n19 VP.n18 24.5923
R2038 VP.n44 VP.n43 21.1495
R2039 VP.n56 VP.n55 21.1495
R2040 VP.n26 VP.n25 21.1495
R2041 VP.n37 VP.n36 10.3291
R2042 VP.n63 VP.n62 10.3291
R2043 VP.n33 VP.n32 10.3291
R2044 VP.n16 VP.n15 9.96756
R2045 VP.n43 VP.n5 3.44336
R2046 VP.n55 VP.n54 3.44336
R2047 VP.n25 VP.n24 3.44336
R2048 VP.n14 VP.n13 3.44336
R2049 VP.n34 VP.n8 0.278335
R2050 VP.n38 VP.n35 0.278335
R2051 VP.n64 VP.n0 0.278335
R2052 VP.n17 VP.n16 0.189894
R2053 VP.n17 VP.n12 0.189894
R2054 VP.n21 VP.n12 0.189894
R2055 VP.n22 VP.n21 0.189894
R2056 VP.n23 VP.n22 0.189894
R2057 VP.n23 VP.n10 0.189894
R2058 VP.n28 VP.n10 0.189894
R2059 VP.n29 VP.n28 0.189894
R2060 VP.n30 VP.n29 0.189894
R2061 VP.n30 VP.n8 0.189894
R2062 VP.n39 VP.n38 0.189894
R2063 VP.n40 VP.n39 0.189894
R2064 VP.n40 VP.n6 0.189894
R2065 VP.n45 VP.n6 0.189894
R2066 VP.n46 VP.n45 0.189894
R2067 VP.n47 VP.n46 0.189894
R2068 VP.n47 VP.n4 0.189894
R2069 VP.n51 VP.n4 0.189894
R2070 VP.n52 VP.n51 0.189894
R2071 VP.n53 VP.n52 0.189894
R2072 VP.n53 VP.n2 0.189894
R2073 VP.n58 VP.n2 0.189894
R2074 VP.n59 VP.n58 0.189894
R2075 VP.n60 VP.n59 0.189894
R2076 VP.n60 VP.n0 0.189894
R2077 VP VP.n64 0.153485
R2078 VDD1 VDD1.n0 60.7821
R2079 VDD1.n3 VDD1.n2 60.6684
R2080 VDD1.n3 VDD1.n1 60.6684
R2081 VDD1.n5 VDD1.n4 59.5858
R2082 VDD1.n5 VDD1.n3 48.6604
R2083 VDD1.n4 VDD1.t6 1.20929
R2084 VDD1.n4 VDD1.t5 1.20929
R2085 VDD1.n0 VDD1.t3 1.20929
R2086 VDD1.n0 VDD1.t1 1.20929
R2087 VDD1.n2 VDD1.t0 1.20929
R2088 VDD1.n2 VDD1.t2 1.20929
R2089 VDD1.n1 VDD1.t7 1.20929
R2090 VDD1.n1 VDD1.t4 1.20929
R2091 VDD1 VDD1.n5 1.08024
C0 VDD1 VN 0.15142f
C1 VDD2 VN 11.419901f
C2 VDD1 VDD2 1.62566f
C3 VTAIL VN 11.5282f
C4 VTAIL VDD1 9.62462f
C5 VTAIL VDD2 9.67709f
C6 VP VN 8.11674f
C7 VDD1 VP 11.7563f
C8 VDD2 VP 0.489028f
C9 VTAIL VP 11.542299f
C10 VDD2 B 5.406326f
C11 VDD1 B 5.811144f
C12 VTAIL B 12.89672f
C13 VN B 14.780049f
C14 VP B 13.249262f
C15 VDD1.t3 B 0.319386f
C16 VDD1.t1 B 0.319386f
C17 VDD1.n0 B 2.90634f
C18 VDD1.t7 B 0.319386f
C19 VDD1.t4 B 0.319386f
C20 VDD1.n1 B 2.90529f
C21 VDD1.t0 B 0.319386f
C22 VDD1.t2 B 0.319386f
C23 VDD1.n2 B 2.90529f
C24 VDD1.n3 B 3.39568f
C25 VDD1.t6 B 0.319386f
C26 VDD1.t5 B 0.319386f
C27 VDD1.n4 B 2.89667f
C28 VDD1.n5 B 3.17326f
C29 VP.n0 B 0.030867f
C30 VP.t5 B 2.43225f
C31 VP.n1 B 0.02279f
C32 VP.n2 B 0.023414f
C33 VP.t7 B 2.43225f
C34 VP.n3 B 0.043418f
C35 VP.n4 B 0.023414f
C36 VP.n5 B 0.024985f
C37 VP.n6 B 0.023414f
C38 VP.n7 B 0.046396f
C39 VP.n8 B 0.030867f
C40 VP.t2 B 2.43225f
C41 VP.n9 B 0.02279f
C42 VP.n10 B 0.023414f
C43 VP.t1 B 2.43225f
C44 VP.n11 B 0.043418f
C45 VP.n12 B 0.023414f
C46 VP.n13 B 0.024985f
C47 VP.t4 B 2.58222f
C48 VP.t6 B 2.43225f
C49 VP.n14 B 0.904488f
C50 VP.n15 B 0.9032f
C51 VP.n16 B 0.201604f
C52 VP.n17 B 0.023414f
C53 VP.n18 B 0.043418f
C54 VP.n19 B 0.034035f
C55 VP.n20 B 0.034035f
C56 VP.n21 B 0.023414f
C57 VP.n22 B 0.023414f
C58 VP.n23 B 0.023414f
C59 VP.n24 B 0.024985f
C60 VP.n25 B 0.849025f
C61 VP.n26 B 0.040418f
C62 VP.n27 B 0.042304f
C63 VP.n28 B 0.023414f
C64 VP.n29 B 0.023414f
C65 VP.n30 B 0.023414f
C66 VP.n31 B 0.046396f
C67 VP.n32 B 0.030987f
C68 VP.n33 B 0.918235f
C69 VP.n34 B 1.40713f
C70 VP.n35 B 1.42312f
C71 VP.t0 B 2.43225f
C72 VP.n36 B 0.918235f
C73 VP.n37 B 0.030987f
C74 VP.n38 B 0.030867f
C75 VP.n39 B 0.023414f
C76 VP.n40 B 0.023414f
C77 VP.n41 B 0.02279f
C78 VP.n42 B 0.042304f
C79 VP.t3 B 2.43225f
C80 VP.n43 B 0.849025f
C81 VP.n44 B 0.040418f
C82 VP.n45 B 0.023414f
C83 VP.n46 B 0.023414f
C84 VP.n47 B 0.023414f
C85 VP.n48 B 0.043418f
C86 VP.n49 B 0.034035f
C87 VP.n50 B 0.034035f
C88 VP.n51 B 0.023414f
C89 VP.n52 B 0.023414f
C90 VP.n53 B 0.023414f
C91 VP.n54 B 0.024985f
C92 VP.n55 B 0.849025f
C93 VP.n56 B 0.040418f
C94 VP.n57 B 0.042304f
C95 VP.n58 B 0.023414f
C96 VP.n59 B 0.023414f
C97 VP.n60 B 0.023414f
C98 VP.n61 B 0.046396f
C99 VP.n62 B 0.030987f
C100 VP.n63 B 0.918235f
C101 VP.n64 B 0.035818f
C102 VTAIL.t8 B 0.241499f
C103 VTAIL.t10 B 0.241499f
C104 VTAIL.n0 B 2.13137f
C105 VTAIL.n1 B 0.328967f
C106 VTAIL.t12 B 2.72017f
C107 VTAIL.n2 B 0.423544f
C108 VTAIL.t5 B 2.72017f
C109 VTAIL.n3 B 0.423544f
C110 VTAIL.t7 B 0.241499f
C111 VTAIL.t3 B 0.241499f
C112 VTAIL.n4 B 2.13137f
C113 VTAIL.n5 B 0.462288f
C114 VTAIL.t4 B 2.72017f
C115 VTAIL.n6 B 1.63446f
C116 VTAIL.t14 B 2.72017f
C117 VTAIL.n7 B 1.63446f
C118 VTAIL.t13 B 0.241499f
C119 VTAIL.t15 B 0.241499f
C120 VTAIL.n8 B 2.13137f
C121 VTAIL.n9 B 0.462286f
C122 VTAIL.t11 B 2.72017f
C123 VTAIL.n10 B 0.423541f
C124 VTAIL.t0 B 2.72017f
C125 VTAIL.n11 B 0.423541f
C126 VTAIL.t6 B 0.241499f
C127 VTAIL.t1 B 0.241499f
C128 VTAIL.n12 B 2.13137f
C129 VTAIL.n13 B 0.462286f
C130 VTAIL.t2 B 2.72017f
C131 VTAIL.n14 B 1.63446f
C132 VTAIL.t9 B 2.72017f
C133 VTAIL.n15 B 1.63096f
C134 VDD2.t2 B 0.316256f
C135 VDD2.t4 B 0.316256f
C136 VDD2.n0 B 2.87681f
C137 VDD2.t6 B 0.316256f
C138 VDD2.t5 B 0.316256f
C139 VDD2.n1 B 2.87681f
C140 VDD2.n2 B 3.31153f
C141 VDD2.t0 B 0.316256f
C142 VDD2.t3 B 0.316256f
C143 VDD2.n3 B 2.86828f
C144 VDD2.n4 B 3.11194f
C145 VDD2.t1 B 0.316256f
C146 VDD2.t7 B 0.316256f
C147 VDD2.n5 B 2.87677f
C148 VN.n0 B 0.030442f
C149 VN.t6 B 2.39875f
C150 VN.n1 B 0.022476f
C151 VN.n2 B 0.023091f
C152 VN.t5 B 2.39875f
C153 VN.n3 B 0.042821f
C154 VN.n4 B 0.023091f
C155 VN.n5 B 0.024641f
C156 VN.t3 B 2.54666f
C157 VN.t7 B 2.39875f
C158 VN.n6 B 0.892031f
C159 VN.n7 B 0.89076f
C160 VN.n8 B 0.198827f
C161 VN.n9 B 0.023091f
C162 VN.n10 B 0.042821f
C163 VN.n11 B 0.033567f
C164 VN.n12 B 0.033567f
C165 VN.n13 B 0.023091f
C166 VN.n14 B 0.023091f
C167 VN.n15 B 0.023091f
C168 VN.n16 B 0.024641f
C169 VN.n17 B 0.837332f
C170 VN.n18 B 0.039861f
C171 VN.n19 B 0.041721f
C172 VN.n20 B 0.023091f
C173 VN.n21 B 0.023091f
C174 VN.n22 B 0.023091f
C175 VN.n23 B 0.045757f
C176 VN.n24 B 0.03056f
C177 VN.n25 B 0.905588f
C178 VN.n26 B 0.035325f
C179 VN.n27 B 0.030442f
C180 VN.t1 B 2.39875f
C181 VN.n28 B 0.022476f
C182 VN.n29 B 0.023091f
C183 VN.t2 B 2.39875f
C184 VN.n30 B 0.042821f
C185 VN.n31 B 0.023091f
C186 VN.n32 B 0.024641f
C187 VN.t4 B 2.54666f
C188 VN.t0 B 2.39875f
C189 VN.n33 B 0.892031f
C190 VN.n34 B 0.89076f
C191 VN.n35 B 0.198827f
C192 VN.n36 B 0.023091f
C193 VN.n37 B 0.042821f
C194 VN.n38 B 0.033567f
C195 VN.n39 B 0.033567f
C196 VN.n40 B 0.023091f
C197 VN.n41 B 0.023091f
C198 VN.n42 B 0.023091f
C199 VN.n43 B 0.024641f
C200 VN.n44 B 0.837332f
C201 VN.n45 B 0.039861f
C202 VN.n46 B 0.041721f
C203 VN.n47 B 0.023091f
C204 VN.n48 B 0.023091f
C205 VN.n49 B 0.023091f
C206 VN.n50 B 0.045757f
C207 VN.n51 B 0.03056f
C208 VN.n52 B 0.905588f
C209 VN.n53 B 1.40006f
.ends

