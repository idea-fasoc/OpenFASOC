* NGSPICE file created from diff_pair_sample_1665.ext - technology: sky130A

.subckt diff_pair_sample_1665 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X1 B.t11 B.t9 B.t10 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=0 ps=0 w=13.64 l=3.98
X2 VTAIL.t3 VN.t0 VDD2.t7 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=2.2506 ps=13.97 w=13.64 l=3.98
X3 B.t8 B.t6 B.t7 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=0 ps=0 w=13.64 l=3.98
X4 VDD2.t6 VN.t1 VTAIL.t2 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X5 VTAIL.t5 VN.t2 VDD2.t5 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X6 VTAIL.t14 VP.t1 VDD1.t0 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=2.2506 ps=13.97 w=13.64 l=3.98
X7 VTAIL.t13 VP.t2 VDD1.t5 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X8 VTAIL.t1 VN.t3 VDD2.t4 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X9 B.t5 B.t3 B.t4 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=0 ps=0 w=13.64 l=3.98
X10 B.t2 B.t0 B.t1 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=0 ps=0 w=13.64 l=3.98
X11 VDD2.t3 VN.t4 VTAIL.t4 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=5.3196 ps=28.06 w=13.64 l=3.98
X12 VDD1.t4 VP.t3 VTAIL.t12 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=5.3196 ps=28.06 w=13.64 l=3.98
X13 VDD1.t7 VP.t4 VTAIL.t11 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X14 VDD1.t6 VP.t5 VTAIL.t10 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X15 VDD2.t2 VN.t5 VTAIL.t7 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=2.2506 ps=13.97 w=13.64 l=3.98
X16 VDD2.t1 VN.t6 VTAIL.t0 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=5.3196 ps=28.06 w=13.64 l=3.98
X17 VTAIL.t6 VN.t7 VDD2.t0 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=2.2506 ps=13.97 w=13.64 l=3.98
X18 VDD1.t3 VP.t6 VTAIL.t9 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=2.2506 pd=13.97 as=5.3196 ps=28.06 w=13.64 l=3.98
X19 VTAIL.t8 VP.t7 VDD1.t2 w_n5280_n3696# sky130_fd_pr__pfet_01v8 ad=5.3196 pd=28.06 as=2.2506 ps=13.97 w=13.64 l=3.98
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n92 VP.n0 161.3
R18 VP.n91 VP.n90 161.3
R19 VP.n89 VP.n1 161.3
R20 VP.n88 VP.n87 161.3
R21 VP.n86 VP.n2 161.3
R22 VP.n85 VP.n84 161.3
R23 VP.n83 VP.n3 161.3
R24 VP.n82 VP.n81 161.3
R25 VP.n79 VP.n4 161.3
R26 VP.n78 VP.n77 161.3
R27 VP.n76 VP.n5 161.3
R28 VP.n75 VP.n74 161.3
R29 VP.n73 VP.n6 161.3
R30 VP.n72 VP.n71 161.3
R31 VP.n70 VP.n7 161.3
R32 VP.n69 VP.n68 161.3
R33 VP.n67 VP.n8 161.3
R34 VP.n65 VP.n64 161.3
R35 VP.n63 VP.n9 161.3
R36 VP.n62 VP.n61 161.3
R37 VP.n60 VP.n10 161.3
R38 VP.n59 VP.n58 161.3
R39 VP.n57 VP.n11 161.3
R40 VP.n56 VP.n55 161.3
R41 VP.n54 VP.n12 161.3
R42 VP.n22 VP.t1 114.624
R43 VP.n53 VP.t7 82.5945
R44 VP.n66 VP.t4 82.5945
R45 VP.n80 VP.t2 82.5945
R46 VP.n93 VP.t6 82.5945
R47 VP.n50 VP.t3 82.5945
R48 VP.n37 VP.t0 82.5945
R49 VP.n23 VP.t5 82.5945
R50 VP.n23 VP.n22 67.3782
R51 VP.n53 VP.n52 59.3461
R52 VP.n94 VP.n93 59.3461
R53 VP.n51 VP.n50 59.3461
R54 VP.n52 VP.n51 58.8747
R55 VP.n60 VP.n59 56.4773
R56 VP.n87 VP.n86 56.4773
R57 VP.n44 VP.n43 56.4773
R58 VP.n73 VP.n72 40.4106
R59 VP.n74 VP.n73 40.4106
R60 VP.n31 VP.n30 40.4106
R61 VP.n30 VP.n29 40.4106
R62 VP.n55 VP.n54 24.3439
R63 VP.n55 VP.n11 24.3439
R64 VP.n59 VP.n11 24.3439
R65 VP.n61 VP.n60 24.3439
R66 VP.n61 VP.n9 24.3439
R67 VP.n65 VP.n9 24.3439
R68 VP.n68 VP.n67 24.3439
R69 VP.n68 VP.n7 24.3439
R70 VP.n72 VP.n7 24.3439
R71 VP.n74 VP.n5 24.3439
R72 VP.n78 VP.n5 24.3439
R73 VP.n79 VP.n78 24.3439
R74 VP.n81 VP.n3 24.3439
R75 VP.n85 VP.n3 24.3439
R76 VP.n86 VP.n85 24.3439
R77 VP.n87 VP.n1 24.3439
R78 VP.n91 VP.n1 24.3439
R79 VP.n92 VP.n91 24.3439
R80 VP.n44 VP.n14 24.3439
R81 VP.n48 VP.n14 24.3439
R82 VP.n49 VP.n48 24.3439
R83 VP.n31 VP.n18 24.3439
R84 VP.n35 VP.n18 24.3439
R85 VP.n36 VP.n35 24.3439
R86 VP.n38 VP.n16 24.3439
R87 VP.n42 VP.n16 24.3439
R88 VP.n43 VP.n42 24.3439
R89 VP.n25 VP.n24 24.3439
R90 VP.n25 VP.n20 24.3439
R91 VP.n29 VP.n20 24.3439
R92 VP.n54 VP.n53 22.6399
R93 VP.n93 VP.n92 22.6399
R94 VP.n50 VP.n49 22.6399
R95 VP.n66 VP.n65 16.7975
R96 VP.n81 VP.n80 16.7975
R97 VP.n38 VP.n37 16.7975
R98 VP.n67 VP.n66 7.54696
R99 VP.n80 VP.n79 7.54696
R100 VP.n37 VP.n36 7.54696
R101 VP.n24 VP.n23 7.54696
R102 VP.n22 VP.n21 2.61018
R103 VP.n51 VP.n13 0.417764
R104 VP.n52 VP.n12 0.417764
R105 VP.n94 VP.n0 0.417764
R106 VP VP.n94 0.394061
R107 VP.n26 VP.n21 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n28 VP.n27 0.189894
R110 VP.n28 VP.n19 0.189894
R111 VP.n32 VP.n19 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n34 VP.n33 0.189894
R114 VP.n34 VP.n17 0.189894
R115 VP.n39 VP.n17 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n41 VP.n40 0.189894
R118 VP.n41 VP.n15 0.189894
R119 VP.n45 VP.n15 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n47 VP.n46 0.189894
R122 VP.n47 VP.n13 0.189894
R123 VP.n56 VP.n12 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n58 VP.n57 0.189894
R126 VP.n58 VP.n10 0.189894
R127 VP.n62 VP.n10 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n64 VP.n63 0.189894
R130 VP.n64 VP.n8 0.189894
R131 VP.n69 VP.n8 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n71 VP.n70 0.189894
R134 VP.n71 VP.n6 0.189894
R135 VP.n75 VP.n6 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n77 VP.n76 0.189894
R138 VP.n77 VP.n4 0.189894
R139 VP.n82 VP.n4 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n84 VP.n83 0.189894
R142 VP.n84 VP.n2 0.189894
R143 VP.n88 VP.n2 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n90 VP.n89 0.189894
R146 VP.n90 VP.n0 0.189894
R147 VDD1 VDD1.n0 75.1105
R148 VDD1.n3 VDD1.n2 74.9967
R149 VDD1.n3 VDD1.n1 74.9967
R150 VDD1.n5 VDD1.n4 73.1944
R151 VDD1.n5 VDD1.n3 52.7768
R152 VDD1.n4 VDD1.t1 2.38356
R153 VDD1.n4 VDD1.t4 2.38356
R154 VDD1.n0 VDD1.t0 2.38356
R155 VDD1.n0 VDD1.t6 2.38356
R156 VDD1.n2 VDD1.t5 2.38356
R157 VDD1.n2 VDD1.t3 2.38356
R158 VDD1.n1 VDD1.t2 2.38356
R159 VDD1.n1 VDD1.t7 2.38356
R160 VDD1 VDD1.n5 1.80007
R161 VTAIL.n11 VTAIL.t14 58.8988
R162 VTAIL.n10 VTAIL.t4 58.8988
R163 VTAIL.n7 VTAIL.t3 58.8988
R164 VTAIL.n15 VTAIL.t0 58.8986
R165 VTAIL.n2 VTAIL.t6 58.8986
R166 VTAIL.n3 VTAIL.t9 58.8986
R167 VTAIL.n6 VTAIL.t8 58.8986
R168 VTAIL.n14 VTAIL.t12 58.8986
R169 VTAIL.n13 VTAIL.n12 56.5158
R170 VTAIL.n9 VTAIL.n8 56.5158
R171 VTAIL.n1 VTAIL.n0 56.5155
R172 VTAIL.n5 VTAIL.n4 56.5155
R173 VTAIL.n15 VTAIL.n14 27.841
R174 VTAIL.n7 VTAIL.n6 27.841
R175 VTAIL.n9 VTAIL.n7 3.71602
R176 VTAIL.n10 VTAIL.n9 3.71602
R177 VTAIL.n13 VTAIL.n11 3.71602
R178 VTAIL.n14 VTAIL.n13 3.71602
R179 VTAIL.n6 VTAIL.n5 3.71602
R180 VTAIL.n5 VTAIL.n3 3.71602
R181 VTAIL.n2 VTAIL.n1 3.71602
R182 VTAIL VTAIL.n15 3.65783
R183 VTAIL.n0 VTAIL.t2 2.38356
R184 VTAIL.n0 VTAIL.t1 2.38356
R185 VTAIL.n4 VTAIL.t11 2.38356
R186 VTAIL.n4 VTAIL.t13 2.38356
R187 VTAIL.n12 VTAIL.t10 2.38356
R188 VTAIL.n12 VTAIL.t15 2.38356
R189 VTAIL.n8 VTAIL.t7 2.38356
R190 VTAIL.n8 VTAIL.t5 2.38356
R191 VTAIL.n11 VTAIL.n10 0.470328
R192 VTAIL.n3 VTAIL.n2 0.470328
R193 VTAIL VTAIL.n1 0.0586897
R194 B.n515 B.n514 585
R195 B.n513 B.n166 585
R196 B.n512 B.n511 585
R197 B.n510 B.n167 585
R198 B.n509 B.n508 585
R199 B.n507 B.n168 585
R200 B.n506 B.n505 585
R201 B.n504 B.n169 585
R202 B.n503 B.n502 585
R203 B.n501 B.n170 585
R204 B.n500 B.n499 585
R205 B.n498 B.n171 585
R206 B.n497 B.n496 585
R207 B.n495 B.n172 585
R208 B.n494 B.n493 585
R209 B.n492 B.n173 585
R210 B.n491 B.n490 585
R211 B.n489 B.n174 585
R212 B.n488 B.n487 585
R213 B.n486 B.n175 585
R214 B.n485 B.n484 585
R215 B.n483 B.n176 585
R216 B.n482 B.n481 585
R217 B.n480 B.n177 585
R218 B.n479 B.n478 585
R219 B.n477 B.n178 585
R220 B.n476 B.n475 585
R221 B.n474 B.n179 585
R222 B.n473 B.n472 585
R223 B.n471 B.n180 585
R224 B.n470 B.n469 585
R225 B.n468 B.n181 585
R226 B.n467 B.n466 585
R227 B.n465 B.n182 585
R228 B.n464 B.n463 585
R229 B.n462 B.n183 585
R230 B.n461 B.n460 585
R231 B.n459 B.n184 585
R232 B.n458 B.n457 585
R233 B.n456 B.n185 585
R234 B.n455 B.n454 585
R235 B.n453 B.n186 585
R236 B.n452 B.n451 585
R237 B.n450 B.n187 585
R238 B.n449 B.n448 585
R239 B.n447 B.n188 585
R240 B.n445 B.n444 585
R241 B.n443 B.n191 585
R242 B.n442 B.n441 585
R243 B.n440 B.n192 585
R244 B.n439 B.n438 585
R245 B.n437 B.n193 585
R246 B.n436 B.n435 585
R247 B.n434 B.n194 585
R248 B.n433 B.n432 585
R249 B.n431 B.n195 585
R250 B.n430 B.n429 585
R251 B.n425 B.n196 585
R252 B.n424 B.n423 585
R253 B.n422 B.n197 585
R254 B.n421 B.n420 585
R255 B.n419 B.n198 585
R256 B.n418 B.n417 585
R257 B.n416 B.n199 585
R258 B.n415 B.n414 585
R259 B.n413 B.n200 585
R260 B.n412 B.n411 585
R261 B.n410 B.n201 585
R262 B.n409 B.n408 585
R263 B.n407 B.n202 585
R264 B.n406 B.n405 585
R265 B.n404 B.n203 585
R266 B.n403 B.n402 585
R267 B.n401 B.n204 585
R268 B.n400 B.n399 585
R269 B.n398 B.n205 585
R270 B.n397 B.n396 585
R271 B.n395 B.n206 585
R272 B.n394 B.n393 585
R273 B.n392 B.n207 585
R274 B.n391 B.n390 585
R275 B.n389 B.n208 585
R276 B.n388 B.n387 585
R277 B.n386 B.n209 585
R278 B.n385 B.n384 585
R279 B.n383 B.n210 585
R280 B.n382 B.n381 585
R281 B.n380 B.n211 585
R282 B.n379 B.n378 585
R283 B.n377 B.n212 585
R284 B.n376 B.n375 585
R285 B.n374 B.n213 585
R286 B.n373 B.n372 585
R287 B.n371 B.n214 585
R288 B.n370 B.n369 585
R289 B.n368 B.n215 585
R290 B.n367 B.n366 585
R291 B.n365 B.n216 585
R292 B.n364 B.n363 585
R293 B.n362 B.n217 585
R294 B.n361 B.n360 585
R295 B.n359 B.n218 585
R296 B.n516 B.n165 585
R297 B.n518 B.n517 585
R298 B.n519 B.n164 585
R299 B.n521 B.n520 585
R300 B.n522 B.n163 585
R301 B.n524 B.n523 585
R302 B.n525 B.n162 585
R303 B.n527 B.n526 585
R304 B.n528 B.n161 585
R305 B.n530 B.n529 585
R306 B.n531 B.n160 585
R307 B.n533 B.n532 585
R308 B.n534 B.n159 585
R309 B.n536 B.n535 585
R310 B.n537 B.n158 585
R311 B.n539 B.n538 585
R312 B.n540 B.n157 585
R313 B.n542 B.n541 585
R314 B.n543 B.n156 585
R315 B.n545 B.n544 585
R316 B.n546 B.n155 585
R317 B.n548 B.n547 585
R318 B.n549 B.n154 585
R319 B.n551 B.n550 585
R320 B.n552 B.n153 585
R321 B.n554 B.n553 585
R322 B.n555 B.n152 585
R323 B.n557 B.n556 585
R324 B.n558 B.n151 585
R325 B.n560 B.n559 585
R326 B.n561 B.n150 585
R327 B.n563 B.n562 585
R328 B.n564 B.n149 585
R329 B.n566 B.n565 585
R330 B.n567 B.n148 585
R331 B.n569 B.n568 585
R332 B.n570 B.n147 585
R333 B.n572 B.n571 585
R334 B.n573 B.n146 585
R335 B.n575 B.n574 585
R336 B.n576 B.n145 585
R337 B.n578 B.n577 585
R338 B.n579 B.n144 585
R339 B.n581 B.n580 585
R340 B.n582 B.n143 585
R341 B.n584 B.n583 585
R342 B.n585 B.n142 585
R343 B.n587 B.n586 585
R344 B.n588 B.n141 585
R345 B.n590 B.n589 585
R346 B.n591 B.n140 585
R347 B.n593 B.n592 585
R348 B.n594 B.n139 585
R349 B.n596 B.n595 585
R350 B.n597 B.n138 585
R351 B.n599 B.n598 585
R352 B.n600 B.n137 585
R353 B.n602 B.n601 585
R354 B.n603 B.n136 585
R355 B.n605 B.n604 585
R356 B.n606 B.n135 585
R357 B.n608 B.n607 585
R358 B.n609 B.n134 585
R359 B.n611 B.n610 585
R360 B.n612 B.n133 585
R361 B.n614 B.n613 585
R362 B.n615 B.n132 585
R363 B.n617 B.n616 585
R364 B.n618 B.n131 585
R365 B.n620 B.n619 585
R366 B.n621 B.n130 585
R367 B.n623 B.n622 585
R368 B.n624 B.n129 585
R369 B.n626 B.n625 585
R370 B.n627 B.n128 585
R371 B.n629 B.n628 585
R372 B.n630 B.n127 585
R373 B.n632 B.n631 585
R374 B.n633 B.n126 585
R375 B.n635 B.n634 585
R376 B.n636 B.n125 585
R377 B.n638 B.n637 585
R378 B.n639 B.n124 585
R379 B.n641 B.n640 585
R380 B.n642 B.n123 585
R381 B.n644 B.n643 585
R382 B.n645 B.n122 585
R383 B.n647 B.n646 585
R384 B.n648 B.n121 585
R385 B.n650 B.n649 585
R386 B.n651 B.n120 585
R387 B.n653 B.n652 585
R388 B.n654 B.n119 585
R389 B.n656 B.n655 585
R390 B.n657 B.n118 585
R391 B.n659 B.n658 585
R392 B.n660 B.n117 585
R393 B.n662 B.n661 585
R394 B.n663 B.n116 585
R395 B.n665 B.n664 585
R396 B.n666 B.n115 585
R397 B.n668 B.n667 585
R398 B.n669 B.n114 585
R399 B.n671 B.n670 585
R400 B.n672 B.n113 585
R401 B.n674 B.n673 585
R402 B.n675 B.n112 585
R403 B.n677 B.n676 585
R404 B.n678 B.n111 585
R405 B.n680 B.n679 585
R406 B.n681 B.n110 585
R407 B.n683 B.n682 585
R408 B.n684 B.n109 585
R409 B.n686 B.n685 585
R410 B.n687 B.n108 585
R411 B.n689 B.n688 585
R412 B.n690 B.n107 585
R413 B.n692 B.n691 585
R414 B.n693 B.n106 585
R415 B.n695 B.n694 585
R416 B.n696 B.n105 585
R417 B.n698 B.n697 585
R418 B.n699 B.n104 585
R419 B.n701 B.n700 585
R420 B.n702 B.n103 585
R421 B.n704 B.n703 585
R422 B.n705 B.n102 585
R423 B.n707 B.n706 585
R424 B.n708 B.n101 585
R425 B.n710 B.n709 585
R426 B.n711 B.n100 585
R427 B.n713 B.n712 585
R428 B.n714 B.n99 585
R429 B.n716 B.n715 585
R430 B.n717 B.n98 585
R431 B.n719 B.n718 585
R432 B.n720 B.n97 585
R433 B.n722 B.n721 585
R434 B.n723 B.n96 585
R435 B.n725 B.n724 585
R436 B.n726 B.n95 585
R437 B.n728 B.n727 585
R438 B.n729 B.n94 585
R439 B.n731 B.n730 585
R440 B.n885 B.n884 585
R441 B.n883 B.n38 585
R442 B.n882 B.n881 585
R443 B.n880 B.n39 585
R444 B.n879 B.n878 585
R445 B.n877 B.n40 585
R446 B.n876 B.n875 585
R447 B.n874 B.n41 585
R448 B.n873 B.n872 585
R449 B.n871 B.n42 585
R450 B.n870 B.n869 585
R451 B.n868 B.n43 585
R452 B.n867 B.n866 585
R453 B.n865 B.n44 585
R454 B.n864 B.n863 585
R455 B.n862 B.n45 585
R456 B.n861 B.n860 585
R457 B.n859 B.n46 585
R458 B.n858 B.n857 585
R459 B.n856 B.n47 585
R460 B.n855 B.n854 585
R461 B.n853 B.n48 585
R462 B.n852 B.n851 585
R463 B.n850 B.n49 585
R464 B.n849 B.n848 585
R465 B.n847 B.n50 585
R466 B.n846 B.n845 585
R467 B.n844 B.n51 585
R468 B.n843 B.n842 585
R469 B.n841 B.n52 585
R470 B.n840 B.n839 585
R471 B.n838 B.n53 585
R472 B.n837 B.n836 585
R473 B.n835 B.n54 585
R474 B.n834 B.n833 585
R475 B.n832 B.n55 585
R476 B.n831 B.n830 585
R477 B.n829 B.n56 585
R478 B.n828 B.n827 585
R479 B.n826 B.n57 585
R480 B.n825 B.n824 585
R481 B.n823 B.n58 585
R482 B.n822 B.n821 585
R483 B.n820 B.n59 585
R484 B.n819 B.n818 585
R485 B.n817 B.n60 585
R486 B.n816 B.n815 585
R487 B.n814 B.n61 585
R488 B.n813 B.n812 585
R489 B.n811 B.n65 585
R490 B.n810 B.n809 585
R491 B.n808 B.n66 585
R492 B.n807 B.n806 585
R493 B.n805 B.n67 585
R494 B.n804 B.n803 585
R495 B.n802 B.n68 585
R496 B.n800 B.n799 585
R497 B.n798 B.n71 585
R498 B.n797 B.n796 585
R499 B.n795 B.n72 585
R500 B.n794 B.n793 585
R501 B.n792 B.n73 585
R502 B.n791 B.n790 585
R503 B.n789 B.n74 585
R504 B.n788 B.n787 585
R505 B.n786 B.n75 585
R506 B.n785 B.n784 585
R507 B.n783 B.n76 585
R508 B.n782 B.n781 585
R509 B.n780 B.n77 585
R510 B.n779 B.n778 585
R511 B.n777 B.n78 585
R512 B.n776 B.n775 585
R513 B.n774 B.n79 585
R514 B.n773 B.n772 585
R515 B.n771 B.n80 585
R516 B.n770 B.n769 585
R517 B.n768 B.n81 585
R518 B.n767 B.n766 585
R519 B.n765 B.n82 585
R520 B.n764 B.n763 585
R521 B.n762 B.n83 585
R522 B.n761 B.n760 585
R523 B.n759 B.n84 585
R524 B.n758 B.n757 585
R525 B.n756 B.n85 585
R526 B.n755 B.n754 585
R527 B.n753 B.n86 585
R528 B.n752 B.n751 585
R529 B.n750 B.n87 585
R530 B.n749 B.n748 585
R531 B.n747 B.n88 585
R532 B.n746 B.n745 585
R533 B.n744 B.n89 585
R534 B.n743 B.n742 585
R535 B.n741 B.n90 585
R536 B.n740 B.n739 585
R537 B.n738 B.n91 585
R538 B.n737 B.n736 585
R539 B.n735 B.n92 585
R540 B.n734 B.n733 585
R541 B.n732 B.n93 585
R542 B.n886 B.n37 585
R543 B.n888 B.n887 585
R544 B.n889 B.n36 585
R545 B.n891 B.n890 585
R546 B.n892 B.n35 585
R547 B.n894 B.n893 585
R548 B.n895 B.n34 585
R549 B.n897 B.n896 585
R550 B.n898 B.n33 585
R551 B.n900 B.n899 585
R552 B.n901 B.n32 585
R553 B.n903 B.n902 585
R554 B.n904 B.n31 585
R555 B.n906 B.n905 585
R556 B.n907 B.n30 585
R557 B.n909 B.n908 585
R558 B.n910 B.n29 585
R559 B.n912 B.n911 585
R560 B.n913 B.n28 585
R561 B.n915 B.n914 585
R562 B.n916 B.n27 585
R563 B.n918 B.n917 585
R564 B.n919 B.n26 585
R565 B.n921 B.n920 585
R566 B.n922 B.n25 585
R567 B.n924 B.n923 585
R568 B.n925 B.n24 585
R569 B.n927 B.n926 585
R570 B.n928 B.n23 585
R571 B.n930 B.n929 585
R572 B.n931 B.n22 585
R573 B.n933 B.n932 585
R574 B.n934 B.n21 585
R575 B.n936 B.n935 585
R576 B.n937 B.n20 585
R577 B.n939 B.n938 585
R578 B.n940 B.n19 585
R579 B.n942 B.n941 585
R580 B.n943 B.n18 585
R581 B.n945 B.n944 585
R582 B.n946 B.n17 585
R583 B.n948 B.n947 585
R584 B.n949 B.n16 585
R585 B.n951 B.n950 585
R586 B.n952 B.n15 585
R587 B.n954 B.n953 585
R588 B.n955 B.n14 585
R589 B.n957 B.n956 585
R590 B.n958 B.n13 585
R591 B.n960 B.n959 585
R592 B.n961 B.n12 585
R593 B.n963 B.n962 585
R594 B.n964 B.n11 585
R595 B.n966 B.n965 585
R596 B.n967 B.n10 585
R597 B.n969 B.n968 585
R598 B.n970 B.n9 585
R599 B.n972 B.n971 585
R600 B.n973 B.n8 585
R601 B.n975 B.n974 585
R602 B.n976 B.n7 585
R603 B.n978 B.n977 585
R604 B.n979 B.n6 585
R605 B.n981 B.n980 585
R606 B.n982 B.n5 585
R607 B.n984 B.n983 585
R608 B.n985 B.n4 585
R609 B.n987 B.n986 585
R610 B.n988 B.n3 585
R611 B.n990 B.n989 585
R612 B.n991 B.n0 585
R613 B.n2 B.n1 585
R614 B.n254 B.n253 585
R615 B.n256 B.n255 585
R616 B.n257 B.n252 585
R617 B.n259 B.n258 585
R618 B.n260 B.n251 585
R619 B.n262 B.n261 585
R620 B.n263 B.n250 585
R621 B.n265 B.n264 585
R622 B.n266 B.n249 585
R623 B.n268 B.n267 585
R624 B.n269 B.n248 585
R625 B.n271 B.n270 585
R626 B.n272 B.n247 585
R627 B.n274 B.n273 585
R628 B.n275 B.n246 585
R629 B.n277 B.n276 585
R630 B.n278 B.n245 585
R631 B.n280 B.n279 585
R632 B.n281 B.n244 585
R633 B.n283 B.n282 585
R634 B.n284 B.n243 585
R635 B.n286 B.n285 585
R636 B.n287 B.n242 585
R637 B.n289 B.n288 585
R638 B.n290 B.n241 585
R639 B.n292 B.n291 585
R640 B.n293 B.n240 585
R641 B.n295 B.n294 585
R642 B.n296 B.n239 585
R643 B.n298 B.n297 585
R644 B.n299 B.n238 585
R645 B.n301 B.n300 585
R646 B.n302 B.n237 585
R647 B.n304 B.n303 585
R648 B.n305 B.n236 585
R649 B.n307 B.n306 585
R650 B.n308 B.n235 585
R651 B.n310 B.n309 585
R652 B.n311 B.n234 585
R653 B.n313 B.n312 585
R654 B.n314 B.n233 585
R655 B.n316 B.n315 585
R656 B.n317 B.n232 585
R657 B.n319 B.n318 585
R658 B.n320 B.n231 585
R659 B.n322 B.n321 585
R660 B.n323 B.n230 585
R661 B.n325 B.n324 585
R662 B.n326 B.n229 585
R663 B.n328 B.n327 585
R664 B.n329 B.n228 585
R665 B.n331 B.n330 585
R666 B.n332 B.n227 585
R667 B.n334 B.n333 585
R668 B.n335 B.n226 585
R669 B.n337 B.n336 585
R670 B.n338 B.n225 585
R671 B.n340 B.n339 585
R672 B.n341 B.n224 585
R673 B.n343 B.n342 585
R674 B.n344 B.n223 585
R675 B.n346 B.n345 585
R676 B.n347 B.n222 585
R677 B.n349 B.n348 585
R678 B.n350 B.n221 585
R679 B.n352 B.n351 585
R680 B.n353 B.n220 585
R681 B.n355 B.n354 585
R682 B.n356 B.n219 585
R683 B.n358 B.n357 585
R684 B.n357 B.n218 535.745
R685 B.n516 B.n515 535.745
R686 B.n732 B.n731 535.745
R687 B.n884 B.n37 535.745
R688 B.n426 B.t0 292.072
R689 B.n189 B.t6 292.072
R690 B.n69 B.t3 292.072
R691 B.n62 B.t9 292.072
R692 B.n993 B.n992 256.663
R693 B.n992 B.n991 235.042
R694 B.n992 B.n2 235.042
R695 B.n189 B.t7 191.141
R696 B.n69 B.t5 191.141
R697 B.n426 B.t1 191.124
R698 B.n62 B.t11 191.124
R699 B.n361 B.n218 163.367
R700 B.n362 B.n361 163.367
R701 B.n363 B.n362 163.367
R702 B.n363 B.n216 163.367
R703 B.n367 B.n216 163.367
R704 B.n368 B.n367 163.367
R705 B.n369 B.n368 163.367
R706 B.n369 B.n214 163.367
R707 B.n373 B.n214 163.367
R708 B.n374 B.n373 163.367
R709 B.n375 B.n374 163.367
R710 B.n375 B.n212 163.367
R711 B.n379 B.n212 163.367
R712 B.n380 B.n379 163.367
R713 B.n381 B.n380 163.367
R714 B.n381 B.n210 163.367
R715 B.n385 B.n210 163.367
R716 B.n386 B.n385 163.367
R717 B.n387 B.n386 163.367
R718 B.n387 B.n208 163.367
R719 B.n391 B.n208 163.367
R720 B.n392 B.n391 163.367
R721 B.n393 B.n392 163.367
R722 B.n393 B.n206 163.367
R723 B.n397 B.n206 163.367
R724 B.n398 B.n397 163.367
R725 B.n399 B.n398 163.367
R726 B.n399 B.n204 163.367
R727 B.n403 B.n204 163.367
R728 B.n404 B.n403 163.367
R729 B.n405 B.n404 163.367
R730 B.n405 B.n202 163.367
R731 B.n409 B.n202 163.367
R732 B.n410 B.n409 163.367
R733 B.n411 B.n410 163.367
R734 B.n411 B.n200 163.367
R735 B.n415 B.n200 163.367
R736 B.n416 B.n415 163.367
R737 B.n417 B.n416 163.367
R738 B.n417 B.n198 163.367
R739 B.n421 B.n198 163.367
R740 B.n422 B.n421 163.367
R741 B.n423 B.n422 163.367
R742 B.n423 B.n196 163.367
R743 B.n430 B.n196 163.367
R744 B.n431 B.n430 163.367
R745 B.n432 B.n431 163.367
R746 B.n432 B.n194 163.367
R747 B.n436 B.n194 163.367
R748 B.n437 B.n436 163.367
R749 B.n438 B.n437 163.367
R750 B.n438 B.n192 163.367
R751 B.n442 B.n192 163.367
R752 B.n443 B.n442 163.367
R753 B.n444 B.n443 163.367
R754 B.n444 B.n188 163.367
R755 B.n449 B.n188 163.367
R756 B.n450 B.n449 163.367
R757 B.n451 B.n450 163.367
R758 B.n451 B.n186 163.367
R759 B.n455 B.n186 163.367
R760 B.n456 B.n455 163.367
R761 B.n457 B.n456 163.367
R762 B.n457 B.n184 163.367
R763 B.n461 B.n184 163.367
R764 B.n462 B.n461 163.367
R765 B.n463 B.n462 163.367
R766 B.n463 B.n182 163.367
R767 B.n467 B.n182 163.367
R768 B.n468 B.n467 163.367
R769 B.n469 B.n468 163.367
R770 B.n469 B.n180 163.367
R771 B.n473 B.n180 163.367
R772 B.n474 B.n473 163.367
R773 B.n475 B.n474 163.367
R774 B.n475 B.n178 163.367
R775 B.n479 B.n178 163.367
R776 B.n480 B.n479 163.367
R777 B.n481 B.n480 163.367
R778 B.n481 B.n176 163.367
R779 B.n485 B.n176 163.367
R780 B.n486 B.n485 163.367
R781 B.n487 B.n486 163.367
R782 B.n487 B.n174 163.367
R783 B.n491 B.n174 163.367
R784 B.n492 B.n491 163.367
R785 B.n493 B.n492 163.367
R786 B.n493 B.n172 163.367
R787 B.n497 B.n172 163.367
R788 B.n498 B.n497 163.367
R789 B.n499 B.n498 163.367
R790 B.n499 B.n170 163.367
R791 B.n503 B.n170 163.367
R792 B.n504 B.n503 163.367
R793 B.n505 B.n504 163.367
R794 B.n505 B.n168 163.367
R795 B.n509 B.n168 163.367
R796 B.n510 B.n509 163.367
R797 B.n511 B.n510 163.367
R798 B.n511 B.n166 163.367
R799 B.n515 B.n166 163.367
R800 B.n731 B.n94 163.367
R801 B.n727 B.n94 163.367
R802 B.n727 B.n726 163.367
R803 B.n726 B.n725 163.367
R804 B.n725 B.n96 163.367
R805 B.n721 B.n96 163.367
R806 B.n721 B.n720 163.367
R807 B.n720 B.n719 163.367
R808 B.n719 B.n98 163.367
R809 B.n715 B.n98 163.367
R810 B.n715 B.n714 163.367
R811 B.n714 B.n713 163.367
R812 B.n713 B.n100 163.367
R813 B.n709 B.n100 163.367
R814 B.n709 B.n708 163.367
R815 B.n708 B.n707 163.367
R816 B.n707 B.n102 163.367
R817 B.n703 B.n102 163.367
R818 B.n703 B.n702 163.367
R819 B.n702 B.n701 163.367
R820 B.n701 B.n104 163.367
R821 B.n697 B.n104 163.367
R822 B.n697 B.n696 163.367
R823 B.n696 B.n695 163.367
R824 B.n695 B.n106 163.367
R825 B.n691 B.n106 163.367
R826 B.n691 B.n690 163.367
R827 B.n690 B.n689 163.367
R828 B.n689 B.n108 163.367
R829 B.n685 B.n108 163.367
R830 B.n685 B.n684 163.367
R831 B.n684 B.n683 163.367
R832 B.n683 B.n110 163.367
R833 B.n679 B.n110 163.367
R834 B.n679 B.n678 163.367
R835 B.n678 B.n677 163.367
R836 B.n677 B.n112 163.367
R837 B.n673 B.n112 163.367
R838 B.n673 B.n672 163.367
R839 B.n672 B.n671 163.367
R840 B.n671 B.n114 163.367
R841 B.n667 B.n114 163.367
R842 B.n667 B.n666 163.367
R843 B.n666 B.n665 163.367
R844 B.n665 B.n116 163.367
R845 B.n661 B.n116 163.367
R846 B.n661 B.n660 163.367
R847 B.n660 B.n659 163.367
R848 B.n659 B.n118 163.367
R849 B.n655 B.n118 163.367
R850 B.n655 B.n654 163.367
R851 B.n654 B.n653 163.367
R852 B.n653 B.n120 163.367
R853 B.n649 B.n120 163.367
R854 B.n649 B.n648 163.367
R855 B.n648 B.n647 163.367
R856 B.n647 B.n122 163.367
R857 B.n643 B.n122 163.367
R858 B.n643 B.n642 163.367
R859 B.n642 B.n641 163.367
R860 B.n641 B.n124 163.367
R861 B.n637 B.n124 163.367
R862 B.n637 B.n636 163.367
R863 B.n636 B.n635 163.367
R864 B.n635 B.n126 163.367
R865 B.n631 B.n126 163.367
R866 B.n631 B.n630 163.367
R867 B.n630 B.n629 163.367
R868 B.n629 B.n128 163.367
R869 B.n625 B.n128 163.367
R870 B.n625 B.n624 163.367
R871 B.n624 B.n623 163.367
R872 B.n623 B.n130 163.367
R873 B.n619 B.n130 163.367
R874 B.n619 B.n618 163.367
R875 B.n618 B.n617 163.367
R876 B.n617 B.n132 163.367
R877 B.n613 B.n132 163.367
R878 B.n613 B.n612 163.367
R879 B.n612 B.n611 163.367
R880 B.n611 B.n134 163.367
R881 B.n607 B.n134 163.367
R882 B.n607 B.n606 163.367
R883 B.n606 B.n605 163.367
R884 B.n605 B.n136 163.367
R885 B.n601 B.n136 163.367
R886 B.n601 B.n600 163.367
R887 B.n600 B.n599 163.367
R888 B.n599 B.n138 163.367
R889 B.n595 B.n138 163.367
R890 B.n595 B.n594 163.367
R891 B.n594 B.n593 163.367
R892 B.n593 B.n140 163.367
R893 B.n589 B.n140 163.367
R894 B.n589 B.n588 163.367
R895 B.n588 B.n587 163.367
R896 B.n587 B.n142 163.367
R897 B.n583 B.n142 163.367
R898 B.n583 B.n582 163.367
R899 B.n582 B.n581 163.367
R900 B.n581 B.n144 163.367
R901 B.n577 B.n144 163.367
R902 B.n577 B.n576 163.367
R903 B.n576 B.n575 163.367
R904 B.n575 B.n146 163.367
R905 B.n571 B.n146 163.367
R906 B.n571 B.n570 163.367
R907 B.n570 B.n569 163.367
R908 B.n569 B.n148 163.367
R909 B.n565 B.n148 163.367
R910 B.n565 B.n564 163.367
R911 B.n564 B.n563 163.367
R912 B.n563 B.n150 163.367
R913 B.n559 B.n150 163.367
R914 B.n559 B.n558 163.367
R915 B.n558 B.n557 163.367
R916 B.n557 B.n152 163.367
R917 B.n553 B.n152 163.367
R918 B.n553 B.n552 163.367
R919 B.n552 B.n551 163.367
R920 B.n551 B.n154 163.367
R921 B.n547 B.n154 163.367
R922 B.n547 B.n546 163.367
R923 B.n546 B.n545 163.367
R924 B.n545 B.n156 163.367
R925 B.n541 B.n156 163.367
R926 B.n541 B.n540 163.367
R927 B.n540 B.n539 163.367
R928 B.n539 B.n158 163.367
R929 B.n535 B.n158 163.367
R930 B.n535 B.n534 163.367
R931 B.n534 B.n533 163.367
R932 B.n533 B.n160 163.367
R933 B.n529 B.n160 163.367
R934 B.n529 B.n528 163.367
R935 B.n528 B.n527 163.367
R936 B.n527 B.n162 163.367
R937 B.n523 B.n162 163.367
R938 B.n523 B.n522 163.367
R939 B.n522 B.n521 163.367
R940 B.n521 B.n164 163.367
R941 B.n517 B.n164 163.367
R942 B.n517 B.n516 163.367
R943 B.n884 B.n883 163.367
R944 B.n883 B.n882 163.367
R945 B.n882 B.n39 163.367
R946 B.n878 B.n39 163.367
R947 B.n878 B.n877 163.367
R948 B.n877 B.n876 163.367
R949 B.n876 B.n41 163.367
R950 B.n872 B.n41 163.367
R951 B.n872 B.n871 163.367
R952 B.n871 B.n870 163.367
R953 B.n870 B.n43 163.367
R954 B.n866 B.n43 163.367
R955 B.n866 B.n865 163.367
R956 B.n865 B.n864 163.367
R957 B.n864 B.n45 163.367
R958 B.n860 B.n45 163.367
R959 B.n860 B.n859 163.367
R960 B.n859 B.n858 163.367
R961 B.n858 B.n47 163.367
R962 B.n854 B.n47 163.367
R963 B.n854 B.n853 163.367
R964 B.n853 B.n852 163.367
R965 B.n852 B.n49 163.367
R966 B.n848 B.n49 163.367
R967 B.n848 B.n847 163.367
R968 B.n847 B.n846 163.367
R969 B.n846 B.n51 163.367
R970 B.n842 B.n51 163.367
R971 B.n842 B.n841 163.367
R972 B.n841 B.n840 163.367
R973 B.n840 B.n53 163.367
R974 B.n836 B.n53 163.367
R975 B.n836 B.n835 163.367
R976 B.n835 B.n834 163.367
R977 B.n834 B.n55 163.367
R978 B.n830 B.n55 163.367
R979 B.n830 B.n829 163.367
R980 B.n829 B.n828 163.367
R981 B.n828 B.n57 163.367
R982 B.n824 B.n57 163.367
R983 B.n824 B.n823 163.367
R984 B.n823 B.n822 163.367
R985 B.n822 B.n59 163.367
R986 B.n818 B.n59 163.367
R987 B.n818 B.n817 163.367
R988 B.n817 B.n816 163.367
R989 B.n816 B.n61 163.367
R990 B.n812 B.n61 163.367
R991 B.n812 B.n811 163.367
R992 B.n811 B.n810 163.367
R993 B.n810 B.n66 163.367
R994 B.n806 B.n66 163.367
R995 B.n806 B.n805 163.367
R996 B.n805 B.n804 163.367
R997 B.n804 B.n68 163.367
R998 B.n799 B.n68 163.367
R999 B.n799 B.n798 163.367
R1000 B.n798 B.n797 163.367
R1001 B.n797 B.n72 163.367
R1002 B.n793 B.n72 163.367
R1003 B.n793 B.n792 163.367
R1004 B.n792 B.n791 163.367
R1005 B.n791 B.n74 163.367
R1006 B.n787 B.n74 163.367
R1007 B.n787 B.n786 163.367
R1008 B.n786 B.n785 163.367
R1009 B.n785 B.n76 163.367
R1010 B.n781 B.n76 163.367
R1011 B.n781 B.n780 163.367
R1012 B.n780 B.n779 163.367
R1013 B.n779 B.n78 163.367
R1014 B.n775 B.n78 163.367
R1015 B.n775 B.n774 163.367
R1016 B.n774 B.n773 163.367
R1017 B.n773 B.n80 163.367
R1018 B.n769 B.n80 163.367
R1019 B.n769 B.n768 163.367
R1020 B.n768 B.n767 163.367
R1021 B.n767 B.n82 163.367
R1022 B.n763 B.n82 163.367
R1023 B.n763 B.n762 163.367
R1024 B.n762 B.n761 163.367
R1025 B.n761 B.n84 163.367
R1026 B.n757 B.n84 163.367
R1027 B.n757 B.n756 163.367
R1028 B.n756 B.n755 163.367
R1029 B.n755 B.n86 163.367
R1030 B.n751 B.n86 163.367
R1031 B.n751 B.n750 163.367
R1032 B.n750 B.n749 163.367
R1033 B.n749 B.n88 163.367
R1034 B.n745 B.n88 163.367
R1035 B.n745 B.n744 163.367
R1036 B.n744 B.n743 163.367
R1037 B.n743 B.n90 163.367
R1038 B.n739 B.n90 163.367
R1039 B.n739 B.n738 163.367
R1040 B.n738 B.n737 163.367
R1041 B.n737 B.n92 163.367
R1042 B.n733 B.n92 163.367
R1043 B.n733 B.n732 163.367
R1044 B.n888 B.n37 163.367
R1045 B.n889 B.n888 163.367
R1046 B.n890 B.n889 163.367
R1047 B.n890 B.n35 163.367
R1048 B.n894 B.n35 163.367
R1049 B.n895 B.n894 163.367
R1050 B.n896 B.n895 163.367
R1051 B.n896 B.n33 163.367
R1052 B.n900 B.n33 163.367
R1053 B.n901 B.n900 163.367
R1054 B.n902 B.n901 163.367
R1055 B.n902 B.n31 163.367
R1056 B.n906 B.n31 163.367
R1057 B.n907 B.n906 163.367
R1058 B.n908 B.n907 163.367
R1059 B.n908 B.n29 163.367
R1060 B.n912 B.n29 163.367
R1061 B.n913 B.n912 163.367
R1062 B.n914 B.n913 163.367
R1063 B.n914 B.n27 163.367
R1064 B.n918 B.n27 163.367
R1065 B.n919 B.n918 163.367
R1066 B.n920 B.n919 163.367
R1067 B.n920 B.n25 163.367
R1068 B.n924 B.n25 163.367
R1069 B.n925 B.n924 163.367
R1070 B.n926 B.n925 163.367
R1071 B.n926 B.n23 163.367
R1072 B.n930 B.n23 163.367
R1073 B.n931 B.n930 163.367
R1074 B.n932 B.n931 163.367
R1075 B.n932 B.n21 163.367
R1076 B.n936 B.n21 163.367
R1077 B.n937 B.n936 163.367
R1078 B.n938 B.n937 163.367
R1079 B.n938 B.n19 163.367
R1080 B.n942 B.n19 163.367
R1081 B.n943 B.n942 163.367
R1082 B.n944 B.n943 163.367
R1083 B.n944 B.n17 163.367
R1084 B.n948 B.n17 163.367
R1085 B.n949 B.n948 163.367
R1086 B.n950 B.n949 163.367
R1087 B.n950 B.n15 163.367
R1088 B.n954 B.n15 163.367
R1089 B.n955 B.n954 163.367
R1090 B.n956 B.n955 163.367
R1091 B.n956 B.n13 163.367
R1092 B.n960 B.n13 163.367
R1093 B.n961 B.n960 163.367
R1094 B.n962 B.n961 163.367
R1095 B.n962 B.n11 163.367
R1096 B.n966 B.n11 163.367
R1097 B.n967 B.n966 163.367
R1098 B.n968 B.n967 163.367
R1099 B.n968 B.n9 163.367
R1100 B.n972 B.n9 163.367
R1101 B.n973 B.n972 163.367
R1102 B.n974 B.n973 163.367
R1103 B.n974 B.n7 163.367
R1104 B.n978 B.n7 163.367
R1105 B.n979 B.n978 163.367
R1106 B.n980 B.n979 163.367
R1107 B.n980 B.n5 163.367
R1108 B.n984 B.n5 163.367
R1109 B.n985 B.n984 163.367
R1110 B.n986 B.n985 163.367
R1111 B.n986 B.n3 163.367
R1112 B.n990 B.n3 163.367
R1113 B.n991 B.n990 163.367
R1114 B.n254 B.n2 163.367
R1115 B.n255 B.n254 163.367
R1116 B.n255 B.n252 163.367
R1117 B.n259 B.n252 163.367
R1118 B.n260 B.n259 163.367
R1119 B.n261 B.n260 163.367
R1120 B.n261 B.n250 163.367
R1121 B.n265 B.n250 163.367
R1122 B.n266 B.n265 163.367
R1123 B.n267 B.n266 163.367
R1124 B.n267 B.n248 163.367
R1125 B.n271 B.n248 163.367
R1126 B.n272 B.n271 163.367
R1127 B.n273 B.n272 163.367
R1128 B.n273 B.n246 163.367
R1129 B.n277 B.n246 163.367
R1130 B.n278 B.n277 163.367
R1131 B.n279 B.n278 163.367
R1132 B.n279 B.n244 163.367
R1133 B.n283 B.n244 163.367
R1134 B.n284 B.n283 163.367
R1135 B.n285 B.n284 163.367
R1136 B.n285 B.n242 163.367
R1137 B.n289 B.n242 163.367
R1138 B.n290 B.n289 163.367
R1139 B.n291 B.n290 163.367
R1140 B.n291 B.n240 163.367
R1141 B.n295 B.n240 163.367
R1142 B.n296 B.n295 163.367
R1143 B.n297 B.n296 163.367
R1144 B.n297 B.n238 163.367
R1145 B.n301 B.n238 163.367
R1146 B.n302 B.n301 163.367
R1147 B.n303 B.n302 163.367
R1148 B.n303 B.n236 163.367
R1149 B.n307 B.n236 163.367
R1150 B.n308 B.n307 163.367
R1151 B.n309 B.n308 163.367
R1152 B.n309 B.n234 163.367
R1153 B.n313 B.n234 163.367
R1154 B.n314 B.n313 163.367
R1155 B.n315 B.n314 163.367
R1156 B.n315 B.n232 163.367
R1157 B.n319 B.n232 163.367
R1158 B.n320 B.n319 163.367
R1159 B.n321 B.n320 163.367
R1160 B.n321 B.n230 163.367
R1161 B.n325 B.n230 163.367
R1162 B.n326 B.n325 163.367
R1163 B.n327 B.n326 163.367
R1164 B.n327 B.n228 163.367
R1165 B.n331 B.n228 163.367
R1166 B.n332 B.n331 163.367
R1167 B.n333 B.n332 163.367
R1168 B.n333 B.n226 163.367
R1169 B.n337 B.n226 163.367
R1170 B.n338 B.n337 163.367
R1171 B.n339 B.n338 163.367
R1172 B.n339 B.n224 163.367
R1173 B.n343 B.n224 163.367
R1174 B.n344 B.n343 163.367
R1175 B.n345 B.n344 163.367
R1176 B.n345 B.n222 163.367
R1177 B.n349 B.n222 163.367
R1178 B.n350 B.n349 163.367
R1179 B.n351 B.n350 163.367
R1180 B.n351 B.n220 163.367
R1181 B.n355 B.n220 163.367
R1182 B.n356 B.n355 163.367
R1183 B.n357 B.n356 163.367
R1184 B.n190 B.t8 107.552
R1185 B.n70 B.t4 107.552
R1186 B.n427 B.t2 107.535
R1187 B.n63 B.t10 107.535
R1188 B.n427 B.n426 83.5884
R1189 B.n190 B.n189 83.5884
R1190 B.n70 B.n69 83.5884
R1191 B.n63 B.n62 83.5884
R1192 B.n428 B.n427 59.5399
R1193 B.n446 B.n190 59.5399
R1194 B.n801 B.n70 59.5399
R1195 B.n64 B.n63 59.5399
R1196 B.n886 B.n885 34.8103
R1197 B.n730 B.n93 34.8103
R1198 B.n514 B.n165 34.8103
R1199 B.n359 B.n358 34.8103
R1200 B B.n993 18.0485
R1201 B.n887 B.n886 10.6151
R1202 B.n887 B.n36 10.6151
R1203 B.n891 B.n36 10.6151
R1204 B.n892 B.n891 10.6151
R1205 B.n893 B.n892 10.6151
R1206 B.n893 B.n34 10.6151
R1207 B.n897 B.n34 10.6151
R1208 B.n898 B.n897 10.6151
R1209 B.n899 B.n898 10.6151
R1210 B.n899 B.n32 10.6151
R1211 B.n903 B.n32 10.6151
R1212 B.n904 B.n903 10.6151
R1213 B.n905 B.n904 10.6151
R1214 B.n905 B.n30 10.6151
R1215 B.n909 B.n30 10.6151
R1216 B.n910 B.n909 10.6151
R1217 B.n911 B.n910 10.6151
R1218 B.n911 B.n28 10.6151
R1219 B.n915 B.n28 10.6151
R1220 B.n916 B.n915 10.6151
R1221 B.n917 B.n916 10.6151
R1222 B.n917 B.n26 10.6151
R1223 B.n921 B.n26 10.6151
R1224 B.n922 B.n921 10.6151
R1225 B.n923 B.n922 10.6151
R1226 B.n923 B.n24 10.6151
R1227 B.n927 B.n24 10.6151
R1228 B.n928 B.n927 10.6151
R1229 B.n929 B.n928 10.6151
R1230 B.n929 B.n22 10.6151
R1231 B.n933 B.n22 10.6151
R1232 B.n934 B.n933 10.6151
R1233 B.n935 B.n934 10.6151
R1234 B.n935 B.n20 10.6151
R1235 B.n939 B.n20 10.6151
R1236 B.n940 B.n939 10.6151
R1237 B.n941 B.n940 10.6151
R1238 B.n941 B.n18 10.6151
R1239 B.n945 B.n18 10.6151
R1240 B.n946 B.n945 10.6151
R1241 B.n947 B.n946 10.6151
R1242 B.n947 B.n16 10.6151
R1243 B.n951 B.n16 10.6151
R1244 B.n952 B.n951 10.6151
R1245 B.n953 B.n952 10.6151
R1246 B.n953 B.n14 10.6151
R1247 B.n957 B.n14 10.6151
R1248 B.n958 B.n957 10.6151
R1249 B.n959 B.n958 10.6151
R1250 B.n959 B.n12 10.6151
R1251 B.n963 B.n12 10.6151
R1252 B.n964 B.n963 10.6151
R1253 B.n965 B.n964 10.6151
R1254 B.n965 B.n10 10.6151
R1255 B.n969 B.n10 10.6151
R1256 B.n970 B.n969 10.6151
R1257 B.n971 B.n970 10.6151
R1258 B.n971 B.n8 10.6151
R1259 B.n975 B.n8 10.6151
R1260 B.n976 B.n975 10.6151
R1261 B.n977 B.n976 10.6151
R1262 B.n977 B.n6 10.6151
R1263 B.n981 B.n6 10.6151
R1264 B.n982 B.n981 10.6151
R1265 B.n983 B.n982 10.6151
R1266 B.n983 B.n4 10.6151
R1267 B.n987 B.n4 10.6151
R1268 B.n988 B.n987 10.6151
R1269 B.n989 B.n988 10.6151
R1270 B.n989 B.n0 10.6151
R1271 B.n885 B.n38 10.6151
R1272 B.n881 B.n38 10.6151
R1273 B.n881 B.n880 10.6151
R1274 B.n880 B.n879 10.6151
R1275 B.n879 B.n40 10.6151
R1276 B.n875 B.n40 10.6151
R1277 B.n875 B.n874 10.6151
R1278 B.n874 B.n873 10.6151
R1279 B.n873 B.n42 10.6151
R1280 B.n869 B.n42 10.6151
R1281 B.n869 B.n868 10.6151
R1282 B.n868 B.n867 10.6151
R1283 B.n867 B.n44 10.6151
R1284 B.n863 B.n44 10.6151
R1285 B.n863 B.n862 10.6151
R1286 B.n862 B.n861 10.6151
R1287 B.n861 B.n46 10.6151
R1288 B.n857 B.n46 10.6151
R1289 B.n857 B.n856 10.6151
R1290 B.n856 B.n855 10.6151
R1291 B.n855 B.n48 10.6151
R1292 B.n851 B.n48 10.6151
R1293 B.n851 B.n850 10.6151
R1294 B.n850 B.n849 10.6151
R1295 B.n849 B.n50 10.6151
R1296 B.n845 B.n50 10.6151
R1297 B.n845 B.n844 10.6151
R1298 B.n844 B.n843 10.6151
R1299 B.n843 B.n52 10.6151
R1300 B.n839 B.n52 10.6151
R1301 B.n839 B.n838 10.6151
R1302 B.n838 B.n837 10.6151
R1303 B.n837 B.n54 10.6151
R1304 B.n833 B.n54 10.6151
R1305 B.n833 B.n832 10.6151
R1306 B.n832 B.n831 10.6151
R1307 B.n831 B.n56 10.6151
R1308 B.n827 B.n56 10.6151
R1309 B.n827 B.n826 10.6151
R1310 B.n826 B.n825 10.6151
R1311 B.n825 B.n58 10.6151
R1312 B.n821 B.n58 10.6151
R1313 B.n821 B.n820 10.6151
R1314 B.n820 B.n819 10.6151
R1315 B.n819 B.n60 10.6151
R1316 B.n815 B.n814 10.6151
R1317 B.n814 B.n813 10.6151
R1318 B.n813 B.n65 10.6151
R1319 B.n809 B.n65 10.6151
R1320 B.n809 B.n808 10.6151
R1321 B.n808 B.n807 10.6151
R1322 B.n807 B.n67 10.6151
R1323 B.n803 B.n67 10.6151
R1324 B.n803 B.n802 10.6151
R1325 B.n800 B.n71 10.6151
R1326 B.n796 B.n71 10.6151
R1327 B.n796 B.n795 10.6151
R1328 B.n795 B.n794 10.6151
R1329 B.n794 B.n73 10.6151
R1330 B.n790 B.n73 10.6151
R1331 B.n790 B.n789 10.6151
R1332 B.n789 B.n788 10.6151
R1333 B.n788 B.n75 10.6151
R1334 B.n784 B.n75 10.6151
R1335 B.n784 B.n783 10.6151
R1336 B.n783 B.n782 10.6151
R1337 B.n782 B.n77 10.6151
R1338 B.n778 B.n77 10.6151
R1339 B.n778 B.n777 10.6151
R1340 B.n777 B.n776 10.6151
R1341 B.n776 B.n79 10.6151
R1342 B.n772 B.n79 10.6151
R1343 B.n772 B.n771 10.6151
R1344 B.n771 B.n770 10.6151
R1345 B.n770 B.n81 10.6151
R1346 B.n766 B.n81 10.6151
R1347 B.n766 B.n765 10.6151
R1348 B.n765 B.n764 10.6151
R1349 B.n764 B.n83 10.6151
R1350 B.n760 B.n83 10.6151
R1351 B.n760 B.n759 10.6151
R1352 B.n759 B.n758 10.6151
R1353 B.n758 B.n85 10.6151
R1354 B.n754 B.n85 10.6151
R1355 B.n754 B.n753 10.6151
R1356 B.n753 B.n752 10.6151
R1357 B.n752 B.n87 10.6151
R1358 B.n748 B.n87 10.6151
R1359 B.n748 B.n747 10.6151
R1360 B.n747 B.n746 10.6151
R1361 B.n746 B.n89 10.6151
R1362 B.n742 B.n89 10.6151
R1363 B.n742 B.n741 10.6151
R1364 B.n741 B.n740 10.6151
R1365 B.n740 B.n91 10.6151
R1366 B.n736 B.n91 10.6151
R1367 B.n736 B.n735 10.6151
R1368 B.n735 B.n734 10.6151
R1369 B.n734 B.n93 10.6151
R1370 B.n730 B.n729 10.6151
R1371 B.n729 B.n728 10.6151
R1372 B.n728 B.n95 10.6151
R1373 B.n724 B.n95 10.6151
R1374 B.n724 B.n723 10.6151
R1375 B.n723 B.n722 10.6151
R1376 B.n722 B.n97 10.6151
R1377 B.n718 B.n97 10.6151
R1378 B.n718 B.n717 10.6151
R1379 B.n717 B.n716 10.6151
R1380 B.n716 B.n99 10.6151
R1381 B.n712 B.n99 10.6151
R1382 B.n712 B.n711 10.6151
R1383 B.n711 B.n710 10.6151
R1384 B.n710 B.n101 10.6151
R1385 B.n706 B.n101 10.6151
R1386 B.n706 B.n705 10.6151
R1387 B.n705 B.n704 10.6151
R1388 B.n704 B.n103 10.6151
R1389 B.n700 B.n103 10.6151
R1390 B.n700 B.n699 10.6151
R1391 B.n699 B.n698 10.6151
R1392 B.n698 B.n105 10.6151
R1393 B.n694 B.n105 10.6151
R1394 B.n694 B.n693 10.6151
R1395 B.n693 B.n692 10.6151
R1396 B.n692 B.n107 10.6151
R1397 B.n688 B.n107 10.6151
R1398 B.n688 B.n687 10.6151
R1399 B.n687 B.n686 10.6151
R1400 B.n686 B.n109 10.6151
R1401 B.n682 B.n109 10.6151
R1402 B.n682 B.n681 10.6151
R1403 B.n681 B.n680 10.6151
R1404 B.n680 B.n111 10.6151
R1405 B.n676 B.n111 10.6151
R1406 B.n676 B.n675 10.6151
R1407 B.n675 B.n674 10.6151
R1408 B.n674 B.n113 10.6151
R1409 B.n670 B.n113 10.6151
R1410 B.n670 B.n669 10.6151
R1411 B.n669 B.n668 10.6151
R1412 B.n668 B.n115 10.6151
R1413 B.n664 B.n115 10.6151
R1414 B.n664 B.n663 10.6151
R1415 B.n663 B.n662 10.6151
R1416 B.n662 B.n117 10.6151
R1417 B.n658 B.n117 10.6151
R1418 B.n658 B.n657 10.6151
R1419 B.n657 B.n656 10.6151
R1420 B.n656 B.n119 10.6151
R1421 B.n652 B.n119 10.6151
R1422 B.n652 B.n651 10.6151
R1423 B.n651 B.n650 10.6151
R1424 B.n650 B.n121 10.6151
R1425 B.n646 B.n121 10.6151
R1426 B.n646 B.n645 10.6151
R1427 B.n645 B.n644 10.6151
R1428 B.n644 B.n123 10.6151
R1429 B.n640 B.n123 10.6151
R1430 B.n640 B.n639 10.6151
R1431 B.n639 B.n638 10.6151
R1432 B.n638 B.n125 10.6151
R1433 B.n634 B.n125 10.6151
R1434 B.n634 B.n633 10.6151
R1435 B.n633 B.n632 10.6151
R1436 B.n632 B.n127 10.6151
R1437 B.n628 B.n127 10.6151
R1438 B.n628 B.n627 10.6151
R1439 B.n627 B.n626 10.6151
R1440 B.n626 B.n129 10.6151
R1441 B.n622 B.n129 10.6151
R1442 B.n622 B.n621 10.6151
R1443 B.n621 B.n620 10.6151
R1444 B.n620 B.n131 10.6151
R1445 B.n616 B.n131 10.6151
R1446 B.n616 B.n615 10.6151
R1447 B.n615 B.n614 10.6151
R1448 B.n614 B.n133 10.6151
R1449 B.n610 B.n133 10.6151
R1450 B.n610 B.n609 10.6151
R1451 B.n609 B.n608 10.6151
R1452 B.n608 B.n135 10.6151
R1453 B.n604 B.n135 10.6151
R1454 B.n604 B.n603 10.6151
R1455 B.n603 B.n602 10.6151
R1456 B.n602 B.n137 10.6151
R1457 B.n598 B.n137 10.6151
R1458 B.n598 B.n597 10.6151
R1459 B.n597 B.n596 10.6151
R1460 B.n596 B.n139 10.6151
R1461 B.n592 B.n139 10.6151
R1462 B.n592 B.n591 10.6151
R1463 B.n591 B.n590 10.6151
R1464 B.n590 B.n141 10.6151
R1465 B.n586 B.n141 10.6151
R1466 B.n586 B.n585 10.6151
R1467 B.n585 B.n584 10.6151
R1468 B.n584 B.n143 10.6151
R1469 B.n580 B.n143 10.6151
R1470 B.n580 B.n579 10.6151
R1471 B.n579 B.n578 10.6151
R1472 B.n578 B.n145 10.6151
R1473 B.n574 B.n145 10.6151
R1474 B.n574 B.n573 10.6151
R1475 B.n573 B.n572 10.6151
R1476 B.n572 B.n147 10.6151
R1477 B.n568 B.n147 10.6151
R1478 B.n568 B.n567 10.6151
R1479 B.n567 B.n566 10.6151
R1480 B.n566 B.n149 10.6151
R1481 B.n562 B.n149 10.6151
R1482 B.n562 B.n561 10.6151
R1483 B.n561 B.n560 10.6151
R1484 B.n560 B.n151 10.6151
R1485 B.n556 B.n151 10.6151
R1486 B.n556 B.n555 10.6151
R1487 B.n555 B.n554 10.6151
R1488 B.n554 B.n153 10.6151
R1489 B.n550 B.n153 10.6151
R1490 B.n550 B.n549 10.6151
R1491 B.n549 B.n548 10.6151
R1492 B.n548 B.n155 10.6151
R1493 B.n544 B.n155 10.6151
R1494 B.n544 B.n543 10.6151
R1495 B.n543 B.n542 10.6151
R1496 B.n542 B.n157 10.6151
R1497 B.n538 B.n157 10.6151
R1498 B.n538 B.n537 10.6151
R1499 B.n537 B.n536 10.6151
R1500 B.n536 B.n159 10.6151
R1501 B.n532 B.n159 10.6151
R1502 B.n532 B.n531 10.6151
R1503 B.n531 B.n530 10.6151
R1504 B.n530 B.n161 10.6151
R1505 B.n526 B.n161 10.6151
R1506 B.n526 B.n525 10.6151
R1507 B.n525 B.n524 10.6151
R1508 B.n524 B.n163 10.6151
R1509 B.n520 B.n163 10.6151
R1510 B.n520 B.n519 10.6151
R1511 B.n519 B.n518 10.6151
R1512 B.n518 B.n165 10.6151
R1513 B.n253 B.n1 10.6151
R1514 B.n256 B.n253 10.6151
R1515 B.n257 B.n256 10.6151
R1516 B.n258 B.n257 10.6151
R1517 B.n258 B.n251 10.6151
R1518 B.n262 B.n251 10.6151
R1519 B.n263 B.n262 10.6151
R1520 B.n264 B.n263 10.6151
R1521 B.n264 B.n249 10.6151
R1522 B.n268 B.n249 10.6151
R1523 B.n269 B.n268 10.6151
R1524 B.n270 B.n269 10.6151
R1525 B.n270 B.n247 10.6151
R1526 B.n274 B.n247 10.6151
R1527 B.n275 B.n274 10.6151
R1528 B.n276 B.n275 10.6151
R1529 B.n276 B.n245 10.6151
R1530 B.n280 B.n245 10.6151
R1531 B.n281 B.n280 10.6151
R1532 B.n282 B.n281 10.6151
R1533 B.n282 B.n243 10.6151
R1534 B.n286 B.n243 10.6151
R1535 B.n287 B.n286 10.6151
R1536 B.n288 B.n287 10.6151
R1537 B.n288 B.n241 10.6151
R1538 B.n292 B.n241 10.6151
R1539 B.n293 B.n292 10.6151
R1540 B.n294 B.n293 10.6151
R1541 B.n294 B.n239 10.6151
R1542 B.n298 B.n239 10.6151
R1543 B.n299 B.n298 10.6151
R1544 B.n300 B.n299 10.6151
R1545 B.n300 B.n237 10.6151
R1546 B.n304 B.n237 10.6151
R1547 B.n305 B.n304 10.6151
R1548 B.n306 B.n305 10.6151
R1549 B.n306 B.n235 10.6151
R1550 B.n310 B.n235 10.6151
R1551 B.n311 B.n310 10.6151
R1552 B.n312 B.n311 10.6151
R1553 B.n312 B.n233 10.6151
R1554 B.n316 B.n233 10.6151
R1555 B.n317 B.n316 10.6151
R1556 B.n318 B.n317 10.6151
R1557 B.n318 B.n231 10.6151
R1558 B.n322 B.n231 10.6151
R1559 B.n323 B.n322 10.6151
R1560 B.n324 B.n323 10.6151
R1561 B.n324 B.n229 10.6151
R1562 B.n328 B.n229 10.6151
R1563 B.n329 B.n328 10.6151
R1564 B.n330 B.n329 10.6151
R1565 B.n330 B.n227 10.6151
R1566 B.n334 B.n227 10.6151
R1567 B.n335 B.n334 10.6151
R1568 B.n336 B.n335 10.6151
R1569 B.n336 B.n225 10.6151
R1570 B.n340 B.n225 10.6151
R1571 B.n341 B.n340 10.6151
R1572 B.n342 B.n341 10.6151
R1573 B.n342 B.n223 10.6151
R1574 B.n346 B.n223 10.6151
R1575 B.n347 B.n346 10.6151
R1576 B.n348 B.n347 10.6151
R1577 B.n348 B.n221 10.6151
R1578 B.n352 B.n221 10.6151
R1579 B.n353 B.n352 10.6151
R1580 B.n354 B.n353 10.6151
R1581 B.n354 B.n219 10.6151
R1582 B.n358 B.n219 10.6151
R1583 B.n360 B.n359 10.6151
R1584 B.n360 B.n217 10.6151
R1585 B.n364 B.n217 10.6151
R1586 B.n365 B.n364 10.6151
R1587 B.n366 B.n365 10.6151
R1588 B.n366 B.n215 10.6151
R1589 B.n370 B.n215 10.6151
R1590 B.n371 B.n370 10.6151
R1591 B.n372 B.n371 10.6151
R1592 B.n372 B.n213 10.6151
R1593 B.n376 B.n213 10.6151
R1594 B.n377 B.n376 10.6151
R1595 B.n378 B.n377 10.6151
R1596 B.n378 B.n211 10.6151
R1597 B.n382 B.n211 10.6151
R1598 B.n383 B.n382 10.6151
R1599 B.n384 B.n383 10.6151
R1600 B.n384 B.n209 10.6151
R1601 B.n388 B.n209 10.6151
R1602 B.n389 B.n388 10.6151
R1603 B.n390 B.n389 10.6151
R1604 B.n390 B.n207 10.6151
R1605 B.n394 B.n207 10.6151
R1606 B.n395 B.n394 10.6151
R1607 B.n396 B.n395 10.6151
R1608 B.n396 B.n205 10.6151
R1609 B.n400 B.n205 10.6151
R1610 B.n401 B.n400 10.6151
R1611 B.n402 B.n401 10.6151
R1612 B.n402 B.n203 10.6151
R1613 B.n406 B.n203 10.6151
R1614 B.n407 B.n406 10.6151
R1615 B.n408 B.n407 10.6151
R1616 B.n408 B.n201 10.6151
R1617 B.n412 B.n201 10.6151
R1618 B.n413 B.n412 10.6151
R1619 B.n414 B.n413 10.6151
R1620 B.n414 B.n199 10.6151
R1621 B.n418 B.n199 10.6151
R1622 B.n419 B.n418 10.6151
R1623 B.n420 B.n419 10.6151
R1624 B.n420 B.n197 10.6151
R1625 B.n424 B.n197 10.6151
R1626 B.n425 B.n424 10.6151
R1627 B.n429 B.n425 10.6151
R1628 B.n433 B.n195 10.6151
R1629 B.n434 B.n433 10.6151
R1630 B.n435 B.n434 10.6151
R1631 B.n435 B.n193 10.6151
R1632 B.n439 B.n193 10.6151
R1633 B.n440 B.n439 10.6151
R1634 B.n441 B.n440 10.6151
R1635 B.n441 B.n191 10.6151
R1636 B.n445 B.n191 10.6151
R1637 B.n448 B.n447 10.6151
R1638 B.n448 B.n187 10.6151
R1639 B.n452 B.n187 10.6151
R1640 B.n453 B.n452 10.6151
R1641 B.n454 B.n453 10.6151
R1642 B.n454 B.n185 10.6151
R1643 B.n458 B.n185 10.6151
R1644 B.n459 B.n458 10.6151
R1645 B.n460 B.n459 10.6151
R1646 B.n460 B.n183 10.6151
R1647 B.n464 B.n183 10.6151
R1648 B.n465 B.n464 10.6151
R1649 B.n466 B.n465 10.6151
R1650 B.n466 B.n181 10.6151
R1651 B.n470 B.n181 10.6151
R1652 B.n471 B.n470 10.6151
R1653 B.n472 B.n471 10.6151
R1654 B.n472 B.n179 10.6151
R1655 B.n476 B.n179 10.6151
R1656 B.n477 B.n476 10.6151
R1657 B.n478 B.n477 10.6151
R1658 B.n478 B.n177 10.6151
R1659 B.n482 B.n177 10.6151
R1660 B.n483 B.n482 10.6151
R1661 B.n484 B.n483 10.6151
R1662 B.n484 B.n175 10.6151
R1663 B.n488 B.n175 10.6151
R1664 B.n489 B.n488 10.6151
R1665 B.n490 B.n489 10.6151
R1666 B.n490 B.n173 10.6151
R1667 B.n494 B.n173 10.6151
R1668 B.n495 B.n494 10.6151
R1669 B.n496 B.n495 10.6151
R1670 B.n496 B.n171 10.6151
R1671 B.n500 B.n171 10.6151
R1672 B.n501 B.n500 10.6151
R1673 B.n502 B.n501 10.6151
R1674 B.n502 B.n169 10.6151
R1675 B.n506 B.n169 10.6151
R1676 B.n507 B.n506 10.6151
R1677 B.n508 B.n507 10.6151
R1678 B.n508 B.n167 10.6151
R1679 B.n512 B.n167 10.6151
R1680 B.n513 B.n512 10.6151
R1681 B.n514 B.n513 10.6151
R1682 B.n64 B.n60 9.36635
R1683 B.n801 B.n800 9.36635
R1684 B.n429 B.n428 9.36635
R1685 B.n447 B.n446 9.36635
R1686 B.n993 B.n0 8.11757
R1687 B.n993 B.n1 8.11757
R1688 B.n815 B.n64 1.24928
R1689 B.n802 B.n801 1.24928
R1690 B.n428 B.n195 1.24928
R1691 B.n446 B.n445 1.24928
R1692 VN.n75 VN.n39 161.3
R1693 VN.n74 VN.n73 161.3
R1694 VN.n72 VN.n40 161.3
R1695 VN.n71 VN.n70 161.3
R1696 VN.n69 VN.n41 161.3
R1697 VN.n68 VN.n67 161.3
R1698 VN.n66 VN.n42 161.3
R1699 VN.n65 VN.n64 161.3
R1700 VN.n62 VN.n43 161.3
R1701 VN.n61 VN.n60 161.3
R1702 VN.n59 VN.n44 161.3
R1703 VN.n58 VN.n57 161.3
R1704 VN.n56 VN.n45 161.3
R1705 VN.n55 VN.n54 161.3
R1706 VN.n53 VN.n46 161.3
R1707 VN.n52 VN.n51 161.3
R1708 VN.n50 VN.n47 161.3
R1709 VN.n36 VN.n0 161.3
R1710 VN.n35 VN.n34 161.3
R1711 VN.n33 VN.n1 161.3
R1712 VN.n32 VN.n31 161.3
R1713 VN.n30 VN.n2 161.3
R1714 VN.n29 VN.n28 161.3
R1715 VN.n27 VN.n3 161.3
R1716 VN.n26 VN.n25 161.3
R1717 VN.n23 VN.n4 161.3
R1718 VN.n22 VN.n21 161.3
R1719 VN.n20 VN.n5 161.3
R1720 VN.n19 VN.n18 161.3
R1721 VN.n17 VN.n6 161.3
R1722 VN.n16 VN.n15 161.3
R1723 VN.n14 VN.n7 161.3
R1724 VN.n13 VN.n12 161.3
R1725 VN.n11 VN.n8 161.3
R1726 VN.n9 VN.t7 114.626
R1727 VN.n48 VN.t4 114.626
R1728 VN.n10 VN.t1 82.5945
R1729 VN.n24 VN.t3 82.5945
R1730 VN.n37 VN.t6 82.5945
R1731 VN.n49 VN.t2 82.5945
R1732 VN.n63 VN.t5 82.5945
R1733 VN.n76 VN.t0 82.5945
R1734 VN.n10 VN.n9 67.3782
R1735 VN.n49 VN.n48 67.3782
R1736 VN.n38 VN.n37 59.3461
R1737 VN.n77 VN.n76 59.3461
R1738 VN VN.n77 58.913
R1739 VN.n31 VN.n30 56.4773
R1740 VN.n70 VN.n69 56.4773
R1741 VN.n17 VN.n16 40.4106
R1742 VN.n18 VN.n17 40.4106
R1743 VN.n56 VN.n55 40.4106
R1744 VN.n57 VN.n56 40.4106
R1745 VN.n12 VN.n11 24.3439
R1746 VN.n12 VN.n7 24.3439
R1747 VN.n16 VN.n7 24.3439
R1748 VN.n18 VN.n5 24.3439
R1749 VN.n22 VN.n5 24.3439
R1750 VN.n23 VN.n22 24.3439
R1751 VN.n25 VN.n3 24.3439
R1752 VN.n29 VN.n3 24.3439
R1753 VN.n30 VN.n29 24.3439
R1754 VN.n31 VN.n1 24.3439
R1755 VN.n35 VN.n1 24.3439
R1756 VN.n36 VN.n35 24.3439
R1757 VN.n55 VN.n46 24.3439
R1758 VN.n51 VN.n46 24.3439
R1759 VN.n51 VN.n50 24.3439
R1760 VN.n69 VN.n68 24.3439
R1761 VN.n68 VN.n42 24.3439
R1762 VN.n64 VN.n42 24.3439
R1763 VN.n62 VN.n61 24.3439
R1764 VN.n61 VN.n44 24.3439
R1765 VN.n57 VN.n44 24.3439
R1766 VN.n75 VN.n74 24.3439
R1767 VN.n74 VN.n40 24.3439
R1768 VN.n70 VN.n40 24.3439
R1769 VN.n37 VN.n36 22.6399
R1770 VN.n76 VN.n75 22.6399
R1771 VN.n25 VN.n24 16.7975
R1772 VN.n64 VN.n63 16.7975
R1773 VN.n11 VN.n10 7.54696
R1774 VN.n24 VN.n23 7.54696
R1775 VN.n50 VN.n49 7.54696
R1776 VN.n63 VN.n62 7.54696
R1777 VN.n48 VN.n47 2.61021
R1778 VN.n9 VN.n8 2.61021
R1779 VN.n77 VN.n39 0.417764
R1780 VN.n38 VN.n0 0.417764
R1781 VN VN.n38 0.394061
R1782 VN.n73 VN.n39 0.189894
R1783 VN.n73 VN.n72 0.189894
R1784 VN.n72 VN.n71 0.189894
R1785 VN.n71 VN.n41 0.189894
R1786 VN.n67 VN.n41 0.189894
R1787 VN.n67 VN.n66 0.189894
R1788 VN.n66 VN.n65 0.189894
R1789 VN.n65 VN.n43 0.189894
R1790 VN.n60 VN.n43 0.189894
R1791 VN.n60 VN.n59 0.189894
R1792 VN.n59 VN.n58 0.189894
R1793 VN.n58 VN.n45 0.189894
R1794 VN.n54 VN.n45 0.189894
R1795 VN.n54 VN.n53 0.189894
R1796 VN.n53 VN.n52 0.189894
R1797 VN.n52 VN.n47 0.189894
R1798 VN.n13 VN.n8 0.189894
R1799 VN.n14 VN.n13 0.189894
R1800 VN.n15 VN.n14 0.189894
R1801 VN.n15 VN.n6 0.189894
R1802 VN.n19 VN.n6 0.189894
R1803 VN.n20 VN.n19 0.189894
R1804 VN.n21 VN.n20 0.189894
R1805 VN.n21 VN.n4 0.189894
R1806 VN.n26 VN.n4 0.189894
R1807 VN.n27 VN.n26 0.189894
R1808 VN.n28 VN.n27 0.189894
R1809 VN.n28 VN.n2 0.189894
R1810 VN.n32 VN.n2 0.189894
R1811 VN.n33 VN.n32 0.189894
R1812 VN.n34 VN.n33 0.189894
R1813 VN.n34 VN.n0 0.189894
R1814 VDD2.n2 VDD2.n1 74.9967
R1815 VDD2.n2 VDD2.n0 74.9967
R1816 VDD2 VDD2.n5 74.9939
R1817 VDD2.n4 VDD2.n3 73.1945
R1818 VDD2.n4 VDD2.n2 52.1937
R1819 VDD2.n5 VDD2.t5 2.38356
R1820 VDD2.n5 VDD2.t3 2.38356
R1821 VDD2.n3 VDD2.t7 2.38356
R1822 VDD2.n3 VDD2.t2 2.38356
R1823 VDD2.n1 VDD2.t4 2.38356
R1824 VDD2.n1 VDD2.t1 2.38356
R1825 VDD2.n0 VDD2.t0 2.38356
R1826 VDD2.n0 VDD2.t6 2.38356
R1827 VDD2 VDD2.n4 1.91645
C0 VP VN 9.663401f
C1 VDD2 B 2.2548f
C2 w_n5280_n3696# VDD1 2.44366f
C3 VP w_n5280_n3696# 11.8655f
C4 VDD2 VDD1 2.49528f
C5 B VDD1 2.11535f
C6 VDD2 VP 0.666339f
C7 B VP 2.72393f
C8 VN VTAIL 11.307099f
C9 VTAIL w_n5280_n3696# 4.67645f
C10 VP VDD1 11.0291f
C11 VN w_n5280_n3696# 11.176f
C12 VDD2 VTAIL 9.22787f
C13 B VTAIL 6.10976f
C14 VDD2 VN 10.518901f
C15 B VN 1.5607f
C16 VDD2 w_n5280_n3696# 2.61626f
C17 VTAIL VDD1 9.1642f
C18 B w_n5280_n3696# 12.6873f
C19 VP VTAIL 11.3212f
C20 VN VDD1 0.154044f
C21 VDD2 VSUBS 2.59805f
C22 VDD1 VSUBS 3.48134f
C23 VTAIL VSUBS 1.672062f
C24 VN VSUBS 8.66651f
C25 VP VSUBS 5.078333f
C26 B VSUBS 6.680069f
C27 w_n5280_n3696# VSUBS 0.239691p
C28 VDD2.t0 VSUBS 0.354983f
C29 VDD2.t6 VSUBS 0.354983f
C30 VDD2.n0 VSUBS 2.87754f
C31 VDD2.t4 VSUBS 0.354983f
C32 VDD2.t1 VSUBS 0.354983f
C33 VDD2.n1 VSUBS 2.87754f
C34 VDD2.n2 VSUBS 6.17978f
C35 VDD2.t7 VSUBS 0.354983f
C36 VDD2.t2 VSUBS 0.354983f
C37 VDD2.n3 VSUBS 2.8484f
C38 VDD2.n4 VSUBS 5.02254f
C39 VDD2.t5 VSUBS 0.354983f
C40 VDD2.t3 VSUBS 0.354983f
C41 VDD2.n5 VSUBS 2.87747f
C42 VN.n0 VSUBS 0.041913f
C43 VN.t6 VSUBS 3.30621f
C44 VN.n1 VSUBS 0.041725f
C45 VN.n2 VSUBS 0.022276f
C46 VN.n3 VSUBS 0.041725f
C47 VN.n4 VSUBS 0.022276f
C48 VN.t3 VSUBS 3.30621f
C49 VN.n5 VSUBS 0.041725f
C50 VN.n6 VSUBS 0.022276f
C51 VN.n7 VSUBS 0.041725f
C52 VN.n8 VSUBS 0.295192f
C53 VN.t1 VSUBS 3.30621f
C54 VN.t7 VSUBS 3.67796f
C55 VN.n9 VSUBS 1.17281f
C56 VN.n10 VSUBS 1.2285f
C57 VN.n11 VSUBS 0.02751f
C58 VN.n12 VSUBS 0.041725f
C59 VN.n13 VSUBS 0.022276f
C60 VN.n14 VSUBS 0.022276f
C61 VN.n15 VSUBS 0.022276f
C62 VN.n16 VSUBS 0.04451f
C63 VN.n17 VSUBS 0.018026f
C64 VN.n18 VSUBS 0.04451f
C65 VN.n19 VSUBS 0.022276f
C66 VN.n20 VSUBS 0.022276f
C67 VN.n21 VSUBS 0.022276f
C68 VN.n22 VSUBS 0.041725f
C69 VN.n23 VSUBS 0.02751f
C70 VN.n24 VSUBS 1.15028f
C71 VN.n25 VSUBS 0.035339f
C72 VN.n26 VSUBS 0.022276f
C73 VN.n27 VSUBS 0.022276f
C74 VN.n28 VSUBS 0.022276f
C75 VN.n29 VSUBS 0.041725f
C76 VN.n30 VSUBS 0.036411f
C77 VN.n31 VSUBS 0.02891f
C78 VN.n32 VSUBS 0.022276f
C79 VN.n33 VSUBS 0.022276f
C80 VN.n34 VSUBS 0.022276f
C81 VN.n35 VSUBS 0.041725f
C82 VN.n36 VSUBS 0.040283f
C83 VN.n37 VSUBS 1.25293f
C84 VN.n38 VSUBS 0.067929f
C85 VN.n39 VSUBS 0.041913f
C86 VN.t0 VSUBS 3.30621f
C87 VN.n40 VSUBS 0.041725f
C88 VN.n41 VSUBS 0.022276f
C89 VN.n42 VSUBS 0.041725f
C90 VN.n43 VSUBS 0.022276f
C91 VN.t5 VSUBS 3.30621f
C92 VN.n44 VSUBS 0.041725f
C93 VN.n45 VSUBS 0.022276f
C94 VN.n46 VSUBS 0.041725f
C95 VN.n47 VSUBS 0.295192f
C96 VN.t2 VSUBS 3.30621f
C97 VN.t4 VSUBS 3.67796f
C98 VN.n48 VSUBS 1.17281f
C99 VN.n49 VSUBS 1.2285f
C100 VN.n50 VSUBS 0.02751f
C101 VN.n51 VSUBS 0.041725f
C102 VN.n52 VSUBS 0.022276f
C103 VN.n53 VSUBS 0.022276f
C104 VN.n54 VSUBS 0.022276f
C105 VN.n55 VSUBS 0.04451f
C106 VN.n56 VSUBS 0.018026f
C107 VN.n57 VSUBS 0.04451f
C108 VN.n58 VSUBS 0.022276f
C109 VN.n59 VSUBS 0.022276f
C110 VN.n60 VSUBS 0.022276f
C111 VN.n61 VSUBS 0.041725f
C112 VN.n62 VSUBS 0.02751f
C113 VN.n63 VSUBS 1.15028f
C114 VN.n64 VSUBS 0.035339f
C115 VN.n65 VSUBS 0.022276f
C116 VN.n66 VSUBS 0.022276f
C117 VN.n67 VSUBS 0.022276f
C118 VN.n68 VSUBS 0.041725f
C119 VN.n69 VSUBS 0.036411f
C120 VN.n70 VSUBS 0.02891f
C121 VN.n71 VSUBS 0.022276f
C122 VN.n72 VSUBS 0.022276f
C123 VN.n73 VSUBS 0.022276f
C124 VN.n74 VSUBS 0.041725f
C125 VN.n75 VSUBS 0.040283f
C126 VN.n76 VSUBS 1.25293f
C127 VN.n77 VSUBS 1.62358f
C128 B.n0 VSUBS 0.007153f
C129 B.n1 VSUBS 0.007153f
C130 B.n2 VSUBS 0.010579f
C131 B.n3 VSUBS 0.008107f
C132 B.n4 VSUBS 0.008107f
C133 B.n5 VSUBS 0.008107f
C134 B.n6 VSUBS 0.008107f
C135 B.n7 VSUBS 0.008107f
C136 B.n8 VSUBS 0.008107f
C137 B.n9 VSUBS 0.008107f
C138 B.n10 VSUBS 0.008107f
C139 B.n11 VSUBS 0.008107f
C140 B.n12 VSUBS 0.008107f
C141 B.n13 VSUBS 0.008107f
C142 B.n14 VSUBS 0.008107f
C143 B.n15 VSUBS 0.008107f
C144 B.n16 VSUBS 0.008107f
C145 B.n17 VSUBS 0.008107f
C146 B.n18 VSUBS 0.008107f
C147 B.n19 VSUBS 0.008107f
C148 B.n20 VSUBS 0.008107f
C149 B.n21 VSUBS 0.008107f
C150 B.n22 VSUBS 0.008107f
C151 B.n23 VSUBS 0.008107f
C152 B.n24 VSUBS 0.008107f
C153 B.n25 VSUBS 0.008107f
C154 B.n26 VSUBS 0.008107f
C155 B.n27 VSUBS 0.008107f
C156 B.n28 VSUBS 0.008107f
C157 B.n29 VSUBS 0.008107f
C158 B.n30 VSUBS 0.008107f
C159 B.n31 VSUBS 0.008107f
C160 B.n32 VSUBS 0.008107f
C161 B.n33 VSUBS 0.008107f
C162 B.n34 VSUBS 0.008107f
C163 B.n35 VSUBS 0.008107f
C164 B.n36 VSUBS 0.008107f
C165 B.n37 VSUBS 0.019537f
C166 B.n38 VSUBS 0.008107f
C167 B.n39 VSUBS 0.008107f
C168 B.n40 VSUBS 0.008107f
C169 B.n41 VSUBS 0.008107f
C170 B.n42 VSUBS 0.008107f
C171 B.n43 VSUBS 0.008107f
C172 B.n44 VSUBS 0.008107f
C173 B.n45 VSUBS 0.008107f
C174 B.n46 VSUBS 0.008107f
C175 B.n47 VSUBS 0.008107f
C176 B.n48 VSUBS 0.008107f
C177 B.n49 VSUBS 0.008107f
C178 B.n50 VSUBS 0.008107f
C179 B.n51 VSUBS 0.008107f
C180 B.n52 VSUBS 0.008107f
C181 B.n53 VSUBS 0.008107f
C182 B.n54 VSUBS 0.008107f
C183 B.n55 VSUBS 0.008107f
C184 B.n56 VSUBS 0.008107f
C185 B.n57 VSUBS 0.008107f
C186 B.n58 VSUBS 0.008107f
C187 B.n59 VSUBS 0.008107f
C188 B.n60 VSUBS 0.00763f
C189 B.n61 VSUBS 0.008107f
C190 B.t10 VSUBS 0.521393f
C191 B.t11 VSUBS 0.555662f
C192 B.t9 VSUBS 2.91988f
C193 B.n62 VSUBS 0.328846f
C194 B.n63 VSUBS 0.089918f
C195 B.n64 VSUBS 0.018782f
C196 B.n65 VSUBS 0.008107f
C197 B.n66 VSUBS 0.008107f
C198 B.n67 VSUBS 0.008107f
C199 B.n68 VSUBS 0.008107f
C200 B.t4 VSUBS 0.521381f
C201 B.t5 VSUBS 0.555652f
C202 B.t3 VSUBS 2.91988f
C203 B.n69 VSUBS 0.328856f
C204 B.n70 VSUBS 0.089931f
C205 B.n71 VSUBS 0.008107f
C206 B.n72 VSUBS 0.008107f
C207 B.n73 VSUBS 0.008107f
C208 B.n74 VSUBS 0.008107f
C209 B.n75 VSUBS 0.008107f
C210 B.n76 VSUBS 0.008107f
C211 B.n77 VSUBS 0.008107f
C212 B.n78 VSUBS 0.008107f
C213 B.n79 VSUBS 0.008107f
C214 B.n80 VSUBS 0.008107f
C215 B.n81 VSUBS 0.008107f
C216 B.n82 VSUBS 0.008107f
C217 B.n83 VSUBS 0.008107f
C218 B.n84 VSUBS 0.008107f
C219 B.n85 VSUBS 0.008107f
C220 B.n86 VSUBS 0.008107f
C221 B.n87 VSUBS 0.008107f
C222 B.n88 VSUBS 0.008107f
C223 B.n89 VSUBS 0.008107f
C224 B.n90 VSUBS 0.008107f
C225 B.n91 VSUBS 0.008107f
C226 B.n92 VSUBS 0.008107f
C227 B.n93 VSUBS 0.020041f
C228 B.n94 VSUBS 0.008107f
C229 B.n95 VSUBS 0.008107f
C230 B.n96 VSUBS 0.008107f
C231 B.n97 VSUBS 0.008107f
C232 B.n98 VSUBS 0.008107f
C233 B.n99 VSUBS 0.008107f
C234 B.n100 VSUBS 0.008107f
C235 B.n101 VSUBS 0.008107f
C236 B.n102 VSUBS 0.008107f
C237 B.n103 VSUBS 0.008107f
C238 B.n104 VSUBS 0.008107f
C239 B.n105 VSUBS 0.008107f
C240 B.n106 VSUBS 0.008107f
C241 B.n107 VSUBS 0.008107f
C242 B.n108 VSUBS 0.008107f
C243 B.n109 VSUBS 0.008107f
C244 B.n110 VSUBS 0.008107f
C245 B.n111 VSUBS 0.008107f
C246 B.n112 VSUBS 0.008107f
C247 B.n113 VSUBS 0.008107f
C248 B.n114 VSUBS 0.008107f
C249 B.n115 VSUBS 0.008107f
C250 B.n116 VSUBS 0.008107f
C251 B.n117 VSUBS 0.008107f
C252 B.n118 VSUBS 0.008107f
C253 B.n119 VSUBS 0.008107f
C254 B.n120 VSUBS 0.008107f
C255 B.n121 VSUBS 0.008107f
C256 B.n122 VSUBS 0.008107f
C257 B.n123 VSUBS 0.008107f
C258 B.n124 VSUBS 0.008107f
C259 B.n125 VSUBS 0.008107f
C260 B.n126 VSUBS 0.008107f
C261 B.n127 VSUBS 0.008107f
C262 B.n128 VSUBS 0.008107f
C263 B.n129 VSUBS 0.008107f
C264 B.n130 VSUBS 0.008107f
C265 B.n131 VSUBS 0.008107f
C266 B.n132 VSUBS 0.008107f
C267 B.n133 VSUBS 0.008107f
C268 B.n134 VSUBS 0.008107f
C269 B.n135 VSUBS 0.008107f
C270 B.n136 VSUBS 0.008107f
C271 B.n137 VSUBS 0.008107f
C272 B.n138 VSUBS 0.008107f
C273 B.n139 VSUBS 0.008107f
C274 B.n140 VSUBS 0.008107f
C275 B.n141 VSUBS 0.008107f
C276 B.n142 VSUBS 0.008107f
C277 B.n143 VSUBS 0.008107f
C278 B.n144 VSUBS 0.008107f
C279 B.n145 VSUBS 0.008107f
C280 B.n146 VSUBS 0.008107f
C281 B.n147 VSUBS 0.008107f
C282 B.n148 VSUBS 0.008107f
C283 B.n149 VSUBS 0.008107f
C284 B.n150 VSUBS 0.008107f
C285 B.n151 VSUBS 0.008107f
C286 B.n152 VSUBS 0.008107f
C287 B.n153 VSUBS 0.008107f
C288 B.n154 VSUBS 0.008107f
C289 B.n155 VSUBS 0.008107f
C290 B.n156 VSUBS 0.008107f
C291 B.n157 VSUBS 0.008107f
C292 B.n158 VSUBS 0.008107f
C293 B.n159 VSUBS 0.008107f
C294 B.n160 VSUBS 0.008107f
C295 B.n161 VSUBS 0.008107f
C296 B.n162 VSUBS 0.008107f
C297 B.n163 VSUBS 0.008107f
C298 B.n164 VSUBS 0.008107f
C299 B.n165 VSUBS 0.020436f
C300 B.n166 VSUBS 0.008107f
C301 B.n167 VSUBS 0.008107f
C302 B.n168 VSUBS 0.008107f
C303 B.n169 VSUBS 0.008107f
C304 B.n170 VSUBS 0.008107f
C305 B.n171 VSUBS 0.008107f
C306 B.n172 VSUBS 0.008107f
C307 B.n173 VSUBS 0.008107f
C308 B.n174 VSUBS 0.008107f
C309 B.n175 VSUBS 0.008107f
C310 B.n176 VSUBS 0.008107f
C311 B.n177 VSUBS 0.008107f
C312 B.n178 VSUBS 0.008107f
C313 B.n179 VSUBS 0.008107f
C314 B.n180 VSUBS 0.008107f
C315 B.n181 VSUBS 0.008107f
C316 B.n182 VSUBS 0.008107f
C317 B.n183 VSUBS 0.008107f
C318 B.n184 VSUBS 0.008107f
C319 B.n185 VSUBS 0.008107f
C320 B.n186 VSUBS 0.008107f
C321 B.n187 VSUBS 0.008107f
C322 B.n188 VSUBS 0.008107f
C323 B.t8 VSUBS 0.521381f
C324 B.t7 VSUBS 0.555652f
C325 B.t6 VSUBS 2.91988f
C326 B.n189 VSUBS 0.328856f
C327 B.n190 VSUBS 0.089931f
C328 B.n191 VSUBS 0.008107f
C329 B.n192 VSUBS 0.008107f
C330 B.n193 VSUBS 0.008107f
C331 B.n194 VSUBS 0.008107f
C332 B.n195 VSUBS 0.00453f
C333 B.n196 VSUBS 0.008107f
C334 B.n197 VSUBS 0.008107f
C335 B.n198 VSUBS 0.008107f
C336 B.n199 VSUBS 0.008107f
C337 B.n200 VSUBS 0.008107f
C338 B.n201 VSUBS 0.008107f
C339 B.n202 VSUBS 0.008107f
C340 B.n203 VSUBS 0.008107f
C341 B.n204 VSUBS 0.008107f
C342 B.n205 VSUBS 0.008107f
C343 B.n206 VSUBS 0.008107f
C344 B.n207 VSUBS 0.008107f
C345 B.n208 VSUBS 0.008107f
C346 B.n209 VSUBS 0.008107f
C347 B.n210 VSUBS 0.008107f
C348 B.n211 VSUBS 0.008107f
C349 B.n212 VSUBS 0.008107f
C350 B.n213 VSUBS 0.008107f
C351 B.n214 VSUBS 0.008107f
C352 B.n215 VSUBS 0.008107f
C353 B.n216 VSUBS 0.008107f
C354 B.n217 VSUBS 0.008107f
C355 B.n218 VSUBS 0.020041f
C356 B.n219 VSUBS 0.008107f
C357 B.n220 VSUBS 0.008107f
C358 B.n221 VSUBS 0.008107f
C359 B.n222 VSUBS 0.008107f
C360 B.n223 VSUBS 0.008107f
C361 B.n224 VSUBS 0.008107f
C362 B.n225 VSUBS 0.008107f
C363 B.n226 VSUBS 0.008107f
C364 B.n227 VSUBS 0.008107f
C365 B.n228 VSUBS 0.008107f
C366 B.n229 VSUBS 0.008107f
C367 B.n230 VSUBS 0.008107f
C368 B.n231 VSUBS 0.008107f
C369 B.n232 VSUBS 0.008107f
C370 B.n233 VSUBS 0.008107f
C371 B.n234 VSUBS 0.008107f
C372 B.n235 VSUBS 0.008107f
C373 B.n236 VSUBS 0.008107f
C374 B.n237 VSUBS 0.008107f
C375 B.n238 VSUBS 0.008107f
C376 B.n239 VSUBS 0.008107f
C377 B.n240 VSUBS 0.008107f
C378 B.n241 VSUBS 0.008107f
C379 B.n242 VSUBS 0.008107f
C380 B.n243 VSUBS 0.008107f
C381 B.n244 VSUBS 0.008107f
C382 B.n245 VSUBS 0.008107f
C383 B.n246 VSUBS 0.008107f
C384 B.n247 VSUBS 0.008107f
C385 B.n248 VSUBS 0.008107f
C386 B.n249 VSUBS 0.008107f
C387 B.n250 VSUBS 0.008107f
C388 B.n251 VSUBS 0.008107f
C389 B.n252 VSUBS 0.008107f
C390 B.n253 VSUBS 0.008107f
C391 B.n254 VSUBS 0.008107f
C392 B.n255 VSUBS 0.008107f
C393 B.n256 VSUBS 0.008107f
C394 B.n257 VSUBS 0.008107f
C395 B.n258 VSUBS 0.008107f
C396 B.n259 VSUBS 0.008107f
C397 B.n260 VSUBS 0.008107f
C398 B.n261 VSUBS 0.008107f
C399 B.n262 VSUBS 0.008107f
C400 B.n263 VSUBS 0.008107f
C401 B.n264 VSUBS 0.008107f
C402 B.n265 VSUBS 0.008107f
C403 B.n266 VSUBS 0.008107f
C404 B.n267 VSUBS 0.008107f
C405 B.n268 VSUBS 0.008107f
C406 B.n269 VSUBS 0.008107f
C407 B.n270 VSUBS 0.008107f
C408 B.n271 VSUBS 0.008107f
C409 B.n272 VSUBS 0.008107f
C410 B.n273 VSUBS 0.008107f
C411 B.n274 VSUBS 0.008107f
C412 B.n275 VSUBS 0.008107f
C413 B.n276 VSUBS 0.008107f
C414 B.n277 VSUBS 0.008107f
C415 B.n278 VSUBS 0.008107f
C416 B.n279 VSUBS 0.008107f
C417 B.n280 VSUBS 0.008107f
C418 B.n281 VSUBS 0.008107f
C419 B.n282 VSUBS 0.008107f
C420 B.n283 VSUBS 0.008107f
C421 B.n284 VSUBS 0.008107f
C422 B.n285 VSUBS 0.008107f
C423 B.n286 VSUBS 0.008107f
C424 B.n287 VSUBS 0.008107f
C425 B.n288 VSUBS 0.008107f
C426 B.n289 VSUBS 0.008107f
C427 B.n290 VSUBS 0.008107f
C428 B.n291 VSUBS 0.008107f
C429 B.n292 VSUBS 0.008107f
C430 B.n293 VSUBS 0.008107f
C431 B.n294 VSUBS 0.008107f
C432 B.n295 VSUBS 0.008107f
C433 B.n296 VSUBS 0.008107f
C434 B.n297 VSUBS 0.008107f
C435 B.n298 VSUBS 0.008107f
C436 B.n299 VSUBS 0.008107f
C437 B.n300 VSUBS 0.008107f
C438 B.n301 VSUBS 0.008107f
C439 B.n302 VSUBS 0.008107f
C440 B.n303 VSUBS 0.008107f
C441 B.n304 VSUBS 0.008107f
C442 B.n305 VSUBS 0.008107f
C443 B.n306 VSUBS 0.008107f
C444 B.n307 VSUBS 0.008107f
C445 B.n308 VSUBS 0.008107f
C446 B.n309 VSUBS 0.008107f
C447 B.n310 VSUBS 0.008107f
C448 B.n311 VSUBS 0.008107f
C449 B.n312 VSUBS 0.008107f
C450 B.n313 VSUBS 0.008107f
C451 B.n314 VSUBS 0.008107f
C452 B.n315 VSUBS 0.008107f
C453 B.n316 VSUBS 0.008107f
C454 B.n317 VSUBS 0.008107f
C455 B.n318 VSUBS 0.008107f
C456 B.n319 VSUBS 0.008107f
C457 B.n320 VSUBS 0.008107f
C458 B.n321 VSUBS 0.008107f
C459 B.n322 VSUBS 0.008107f
C460 B.n323 VSUBS 0.008107f
C461 B.n324 VSUBS 0.008107f
C462 B.n325 VSUBS 0.008107f
C463 B.n326 VSUBS 0.008107f
C464 B.n327 VSUBS 0.008107f
C465 B.n328 VSUBS 0.008107f
C466 B.n329 VSUBS 0.008107f
C467 B.n330 VSUBS 0.008107f
C468 B.n331 VSUBS 0.008107f
C469 B.n332 VSUBS 0.008107f
C470 B.n333 VSUBS 0.008107f
C471 B.n334 VSUBS 0.008107f
C472 B.n335 VSUBS 0.008107f
C473 B.n336 VSUBS 0.008107f
C474 B.n337 VSUBS 0.008107f
C475 B.n338 VSUBS 0.008107f
C476 B.n339 VSUBS 0.008107f
C477 B.n340 VSUBS 0.008107f
C478 B.n341 VSUBS 0.008107f
C479 B.n342 VSUBS 0.008107f
C480 B.n343 VSUBS 0.008107f
C481 B.n344 VSUBS 0.008107f
C482 B.n345 VSUBS 0.008107f
C483 B.n346 VSUBS 0.008107f
C484 B.n347 VSUBS 0.008107f
C485 B.n348 VSUBS 0.008107f
C486 B.n349 VSUBS 0.008107f
C487 B.n350 VSUBS 0.008107f
C488 B.n351 VSUBS 0.008107f
C489 B.n352 VSUBS 0.008107f
C490 B.n353 VSUBS 0.008107f
C491 B.n354 VSUBS 0.008107f
C492 B.n355 VSUBS 0.008107f
C493 B.n356 VSUBS 0.008107f
C494 B.n357 VSUBS 0.019537f
C495 B.n358 VSUBS 0.019537f
C496 B.n359 VSUBS 0.020041f
C497 B.n360 VSUBS 0.008107f
C498 B.n361 VSUBS 0.008107f
C499 B.n362 VSUBS 0.008107f
C500 B.n363 VSUBS 0.008107f
C501 B.n364 VSUBS 0.008107f
C502 B.n365 VSUBS 0.008107f
C503 B.n366 VSUBS 0.008107f
C504 B.n367 VSUBS 0.008107f
C505 B.n368 VSUBS 0.008107f
C506 B.n369 VSUBS 0.008107f
C507 B.n370 VSUBS 0.008107f
C508 B.n371 VSUBS 0.008107f
C509 B.n372 VSUBS 0.008107f
C510 B.n373 VSUBS 0.008107f
C511 B.n374 VSUBS 0.008107f
C512 B.n375 VSUBS 0.008107f
C513 B.n376 VSUBS 0.008107f
C514 B.n377 VSUBS 0.008107f
C515 B.n378 VSUBS 0.008107f
C516 B.n379 VSUBS 0.008107f
C517 B.n380 VSUBS 0.008107f
C518 B.n381 VSUBS 0.008107f
C519 B.n382 VSUBS 0.008107f
C520 B.n383 VSUBS 0.008107f
C521 B.n384 VSUBS 0.008107f
C522 B.n385 VSUBS 0.008107f
C523 B.n386 VSUBS 0.008107f
C524 B.n387 VSUBS 0.008107f
C525 B.n388 VSUBS 0.008107f
C526 B.n389 VSUBS 0.008107f
C527 B.n390 VSUBS 0.008107f
C528 B.n391 VSUBS 0.008107f
C529 B.n392 VSUBS 0.008107f
C530 B.n393 VSUBS 0.008107f
C531 B.n394 VSUBS 0.008107f
C532 B.n395 VSUBS 0.008107f
C533 B.n396 VSUBS 0.008107f
C534 B.n397 VSUBS 0.008107f
C535 B.n398 VSUBS 0.008107f
C536 B.n399 VSUBS 0.008107f
C537 B.n400 VSUBS 0.008107f
C538 B.n401 VSUBS 0.008107f
C539 B.n402 VSUBS 0.008107f
C540 B.n403 VSUBS 0.008107f
C541 B.n404 VSUBS 0.008107f
C542 B.n405 VSUBS 0.008107f
C543 B.n406 VSUBS 0.008107f
C544 B.n407 VSUBS 0.008107f
C545 B.n408 VSUBS 0.008107f
C546 B.n409 VSUBS 0.008107f
C547 B.n410 VSUBS 0.008107f
C548 B.n411 VSUBS 0.008107f
C549 B.n412 VSUBS 0.008107f
C550 B.n413 VSUBS 0.008107f
C551 B.n414 VSUBS 0.008107f
C552 B.n415 VSUBS 0.008107f
C553 B.n416 VSUBS 0.008107f
C554 B.n417 VSUBS 0.008107f
C555 B.n418 VSUBS 0.008107f
C556 B.n419 VSUBS 0.008107f
C557 B.n420 VSUBS 0.008107f
C558 B.n421 VSUBS 0.008107f
C559 B.n422 VSUBS 0.008107f
C560 B.n423 VSUBS 0.008107f
C561 B.n424 VSUBS 0.008107f
C562 B.n425 VSUBS 0.008107f
C563 B.t2 VSUBS 0.521393f
C564 B.t1 VSUBS 0.555662f
C565 B.t0 VSUBS 2.91988f
C566 B.n426 VSUBS 0.328846f
C567 B.n427 VSUBS 0.089918f
C568 B.n428 VSUBS 0.018782f
C569 B.n429 VSUBS 0.00763f
C570 B.n430 VSUBS 0.008107f
C571 B.n431 VSUBS 0.008107f
C572 B.n432 VSUBS 0.008107f
C573 B.n433 VSUBS 0.008107f
C574 B.n434 VSUBS 0.008107f
C575 B.n435 VSUBS 0.008107f
C576 B.n436 VSUBS 0.008107f
C577 B.n437 VSUBS 0.008107f
C578 B.n438 VSUBS 0.008107f
C579 B.n439 VSUBS 0.008107f
C580 B.n440 VSUBS 0.008107f
C581 B.n441 VSUBS 0.008107f
C582 B.n442 VSUBS 0.008107f
C583 B.n443 VSUBS 0.008107f
C584 B.n444 VSUBS 0.008107f
C585 B.n445 VSUBS 0.00453f
C586 B.n446 VSUBS 0.018782f
C587 B.n447 VSUBS 0.00763f
C588 B.n448 VSUBS 0.008107f
C589 B.n449 VSUBS 0.008107f
C590 B.n450 VSUBS 0.008107f
C591 B.n451 VSUBS 0.008107f
C592 B.n452 VSUBS 0.008107f
C593 B.n453 VSUBS 0.008107f
C594 B.n454 VSUBS 0.008107f
C595 B.n455 VSUBS 0.008107f
C596 B.n456 VSUBS 0.008107f
C597 B.n457 VSUBS 0.008107f
C598 B.n458 VSUBS 0.008107f
C599 B.n459 VSUBS 0.008107f
C600 B.n460 VSUBS 0.008107f
C601 B.n461 VSUBS 0.008107f
C602 B.n462 VSUBS 0.008107f
C603 B.n463 VSUBS 0.008107f
C604 B.n464 VSUBS 0.008107f
C605 B.n465 VSUBS 0.008107f
C606 B.n466 VSUBS 0.008107f
C607 B.n467 VSUBS 0.008107f
C608 B.n468 VSUBS 0.008107f
C609 B.n469 VSUBS 0.008107f
C610 B.n470 VSUBS 0.008107f
C611 B.n471 VSUBS 0.008107f
C612 B.n472 VSUBS 0.008107f
C613 B.n473 VSUBS 0.008107f
C614 B.n474 VSUBS 0.008107f
C615 B.n475 VSUBS 0.008107f
C616 B.n476 VSUBS 0.008107f
C617 B.n477 VSUBS 0.008107f
C618 B.n478 VSUBS 0.008107f
C619 B.n479 VSUBS 0.008107f
C620 B.n480 VSUBS 0.008107f
C621 B.n481 VSUBS 0.008107f
C622 B.n482 VSUBS 0.008107f
C623 B.n483 VSUBS 0.008107f
C624 B.n484 VSUBS 0.008107f
C625 B.n485 VSUBS 0.008107f
C626 B.n486 VSUBS 0.008107f
C627 B.n487 VSUBS 0.008107f
C628 B.n488 VSUBS 0.008107f
C629 B.n489 VSUBS 0.008107f
C630 B.n490 VSUBS 0.008107f
C631 B.n491 VSUBS 0.008107f
C632 B.n492 VSUBS 0.008107f
C633 B.n493 VSUBS 0.008107f
C634 B.n494 VSUBS 0.008107f
C635 B.n495 VSUBS 0.008107f
C636 B.n496 VSUBS 0.008107f
C637 B.n497 VSUBS 0.008107f
C638 B.n498 VSUBS 0.008107f
C639 B.n499 VSUBS 0.008107f
C640 B.n500 VSUBS 0.008107f
C641 B.n501 VSUBS 0.008107f
C642 B.n502 VSUBS 0.008107f
C643 B.n503 VSUBS 0.008107f
C644 B.n504 VSUBS 0.008107f
C645 B.n505 VSUBS 0.008107f
C646 B.n506 VSUBS 0.008107f
C647 B.n507 VSUBS 0.008107f
C648 B.n508 VSUBS 0.008107f
C649 B.n509 VSUBS 0.008107f
C650 B.n510 VSUBS 0.008107f
C651 B.n511 VSUBS 0.008107f
C652 B.n512 VSUBS 0.008107f
C653 B.n513 VSUBS 0.008107f
C654 B.n514 VSUBS 0.019143f
C655 B.n515 VSUBS 0.020041f
C656 B.n516 VSUBS 0.019537f
C657 B.n517 VSUBS 0.008107f
C658 B.n518 VSUBS 0.008107f
C659 B.n519 VSUBS 0.008107f
C660 B.n520 VSUBS 0.008107f
C661 B.n521 VSUBS 0.008107f
C662 B.n522 VSUBS 0.008107f
C663 B.n523 VSUBS 0.008107f
C664 B.n524 VSUBS 0.008107f
C665 B.n525 VSUBS 0.008107f
C666 B.n526 VSUBS 0.008107f
C667 B.n527 VSUBS 0.008107f
C668 B.n528 VSUBS 0.008107f
C669 B.n529 VSUBS 0.008107f
C670 B.n530 VSUBS 0.008107f
C671 B.n531 VSUBS 0.008107f
C672 B.n532 VSUBS 0.008107f
C673 B.n533 VSUBS 0.008107f
C674 B.n534 VSUBS 0.008107f
C675 B.n535 VSUBS 0.008107f
C676 B.n536 VSUBS 0.008107f
C677 B.n537 VSUBS 0.008107f
C678 B.n538 VSUBS 0.008107f
C679 B.n539 VSUBS 0.008107f
C680 B.n540 VSUBS 0.008107f
C681 B.n541 VSUBS 0.008107f
C682 B.n542 VSUBS 0.008107f
C683 B.n543 VSUBS 0.008107f
C684 B.n544 VSUBS 0.008107f
C685 B.n545 VSUBS 0.008107f
C686 B.n546 VSUBS 0.008107f
C687 B.n547 VSUBS 0.008107f
C688 B.n548 VSUBS 0.008107f
C689 B.n549 VSUBS 0.008107f
C690 B.n550 VSUBS 0.008107f
C691 B.n551 VSUBS 0.008107f
C692 B.n552 VSUBS 0.008107f
C693 B.n553 VSUBS 0.008107f
C694 B.n554 VSUBS 0.008107f
C695 B.n555 VSUBS 0.008107f
C696 B.n556 VSUBS 0.008107f
C697 B.n557 VSUBS 0.008107f
C698 B.n558 VSUBS 0.008107f
C699 B.n559 VSUBS 0.008107f
C700 B.n560 VSUBS 0.008107f
C701 B.n561 VSUBS 0.008107f
C702 B.n562 VSUBS 0.008107f
C703 B.n563 VSUBS 0.008107f
C704 B.n564 VSUBS 0.008107f
C705 B.n565 VSUBS 0.008107f
C706 B.n566 VSUBS 0.008107f
C707 B.n567 VSUBS 0.008107f
C708 B.n568 VSUBS 0.008107f
C709 B.n569 VSUBS 0.008107f
C710 B.n570 VSUBS 0.008107f
C711 B.n571 VSUBS 0.008107f
C712 B.n572 VSUBS 0.008107f
C713 B.n573 VSUBS 0.008107f
C714 B.n574 VSUBS 0.008107f
C715 B.n575 VSUBS 0.008107f
C716 B.n576 VSUBS 0.008107f
C717 B.n577 VSUBS 0.008107f
C718 B.n578 VSUBS 0.008107f
C719 B.n579 VSUBS 0.008107f
C720 B.n580 VSUBS 0.008107f
C721 B.n581 VSUBS 0.008107f
C722 B.n582 VSUBS 0.008107f
C723 B.n583 VSUBS 0.008107f
C724 B.n584 VSUBS 0.008107f
C725 B.n585 VSUBS 0.008107f
C726 B.n586 VSUBS 0.008107f
C727 B.n587 VSUBS 0.008107f
C728 B.n588 VSUBS 0.008107f
C729 B.n589 VSUBS 0.008107f
C730 B.n590 VSUBS 0.008107f
C731 B.n591 VSUBS 0.008107f
C732 B.n592 VSUBS 0.008107f
C733 B.n593 VSUBS 0.008107f
C734 B.n594 VSUBS 0.008107f
C735 B.n595 VSUBS 0.008107f
C736 B.n596 VSUBS 0.008107f
C737 B.n597 VSUBS 0.008107f
C738 B.n598 VSUBS 0.008107f
C739 B.n599 VSUBS 0.008107f
C740 B.n600 VSUBS 0.008107f
C741 B.n601 VSUBS 0.008107f
C742 B.n602 VSUBS 0.008107f
C743 B.n603 VSUBS 0.008107f
C744 B.n604 VSUBS 0.008107f
C745 B.n605 VSUBS 0.008107f
C746 B.n606 VSUBS 0.008107f
C747 B.n607 VSUBS 0.008107f
C748 B.n608 VSUBS 0.008107f
C749 B.n609 VSUBS 0.008107f
C750 B.n610 VSUBS 0.008107f
C751 B.n611 VSUBS 0.008107f
C752 B.n612 VSUBS 0.008107f
C753 B.n613 VSUBS 0.008107f
C754 B.n614 VSUBS 0.008107f
C755 B.n615 VSUBS 0.008107f
C756 B.n616 VSUBS 0.008107f
C757 B.n617 VSUBS 0.008107f
C758 B.n618 VSUBS 0.008107f
C759 B.n619 VSUBS 0.008107f
C760 B.n620 VSUBS 0.008107f
C761 B.n621 VSUBS 0.008107f
C762 B.n622 VSUBS 0.008107f
C763 B.n623 VSUBS 0.008107f
C764 B.n624 VSUBS 0.008107f
C765 B.n625 VSUBS 0.008107f
C766 B.n626 VSUBS 0.008107f
C767 B.n627 VSUBS 0.008107f
C768 B.n628 VSUBS 0.008107f
C769 B.n629 VSUBS 0.008107f
C770 B.n630 VSUBS 0.008107f
C771 B.n631 VSUBS 0.008107f
C772 B.n632 VSUBS 0.008107f
C773 B.n633 VSUBS 0.008107f
C774 B.n634 VSUBS 0.008107f
C775 B.n635 VSUBS 0.008107f
C776 B.n636 VSUBS 0.008107f
C777 B.n637 VSUBS 0.008107f
C778 B.n638 VSUBS 0.008107f
C779 B.n639 VSUBS 0.008107f
C780 B.n640 VSUBS 0.008107f
C781 B.n641 VSUBS 0.008107f
C782 B.n642 VSUBS 0.008107f
C783 B.n643 VSUBS 0.008107f
C784 B.n644 VSUBS 0.008107f
C785 B.n645 VSUBS 0.008107f
C786 B.n646 VSUBS 0.008107f
C787 B.n647 VSUBS 0.008107f
C788 B.n648 VSUBS 0.008107f
C789 B.n649 VSUBS 0.008107f
C790 B.n650 VSUBS 0.008107f
C791 B.n651 VSUBS 0.008107f
C792 B.n652 VSUBS 0.008107f
C793 B.n653 VSUBS 0.008107f
C794 B.n654 VSUBS 0.008107f
C795 B.n655 VSUBS 0.008107f
C796 B.n656 VSUBS 0.008107f
C797 B.n657 VSUBS 0.008107f
C798 B.n658 VSUBS 0.008107f
C799 B.n659 VSUBS 0.008107f
C800 B.n660 VSUBS 0.008107f
C801 B.n661 VSUBS 0.008107f
C802 B.n662 VSUBS 0.008107f
C803 B.n663 VSUBS 0.008107f
C804 B.n664 VSUBS 0.008107f
C805 B.n665 VSUBS 0.008107f
C806 B.n666 VSUBS 0.008107f
C807 B.n667 VSUBS 0.008107f
C808 B.n668 VSUBS 0.008107f
C809 B.n669 VSUBS 0.008107f
C810 B.n670 VSUBS 0.008107f
C811 B.n671 VSUBS 0.008107f
C812 B.n672 VSUBS 0.008107f
C813 B.n673 VSUBS 0.008107f
C814 B.n674 VSUBS 0.008107f
C815 B.n675 VSUBS 0.008107f
C816 B.n676 VSUBS 0.008107f
C817 B.n677 VSUBS 0.008107f
C818 B.n678 VSUBS 0.008107f
C819 B.n679 VSUBS 0.008107f
C820 B.n680 VSUBS 0.008107f
C821 B.n681 VSUBS 0.008107f
C822 B.n682 VSUBS 0.008107f
C823 B.n683 VSUBS 0.008107f
C824 B.n684 VSUBS 0.008107f
C825 B.n685 VSUBS 0.008107f
C826 B.n686 VSUBS 0.008107f
C827 B.n687 VSUBS 0.008107f
C828 B.n688 VSUBS 0.008107f
C829 B.n689 VSUBS 0.008107f
C830 B.n690 VSUBS 0.008107f
C831 B.n691 VSUBS 0.008107f
C832 B.n692 VSUBS 0.008107f
C833 B.n693 VSUBS 0.008107f
C834 B.n694 VSUBS 0.008107f
C835 B.n695 VSUBS 0.008107f
C836 B.n696 VSUBS 0.008107f
C837 B.n697 VSUBS 0.008107f
C838 B.n698 VSUBS 0.008107f
C839 B.n699 VSUBS 0.008107f
C840 B.n700 VSUBS 0.008107f
C841 B.n701 VSUBS 0.008107f
C842 B.n702 VSUBS 0.008107f
C843 B.n703 VSUBS 0.008107f
C844 B.n704 VSUBS 0.008107f
C845 B.n705 VSUBS 0.008107f
C846 B.n706 VSUBS 0.008107f
C847 B.n707 VSUBS 0.008107f
C848 B.n708 VSUBS 0.008107f
C849 B.n709 VSUBS 0.008107f
C850 B.n710 VSUBS 0.008107f
C851 B.n711 VSUBS 0.008107f
C852 B.n712 VSUBS 0.008107f
C853 B.n713 VSUBS 0.008107f
C854 B.n714 VSUBS 0.008107f
C855 B.n715 VSUBS 0.008107f
C856 B.n716 VSUBS 0.008107f
C857 B.n717 VSUBS 0.008107f
C858 B.n718 VSUBS 0.008107f
C859 B.n719 VSUBS 0.008107f
C860 B.n720 VSUBS 0.008107f
C861 B.n721 VSUBS 0.008107f
C862 B.n722 VSUBS 0.008107f
C863 B.n723 VSUBS 0.008107f
C864 B.n724 VSUBS 0.008107f
C865 B.n725 VSUBS 0.008107f
C866 B.n726 VSUBS 0.008107f
C867 B.n727 VSUBS 0.008107f
C868 B.n728 VSUBS 0.008107f
C869 B.n729 VSUBS 0.008107f
C870 B.n730 VSUBS 0.019537f
C871 B.n731 VSUBS 0.019537f
C872 B.n732 VSUBS 0.020041f
C873 B.n733 VSUBS 0.008107f
C874 B.n734 VSUBS 0.008107f
C875 B.n735 VSUBS 0.008107f
C876 B.n736 VSUBS 0.008107f
C877 B.n737 VSUBS 0.008107f
C878 B.n738 VSUBS 0.008107f
C879 B.n739 VSUBS 0.008107f
C880 B.n740 VSUBS 0.008107f
C881 B.n741 VSUBS 0.008107f
C882 B.n742 VSUBS 0.008107f
C883 B.n743 VSUBS 0.008107f
C884 B.n744 VSUBS 0.008107f
C885 B.n745 VSUBS 0.008107f
C886 B.n746 VSUBS 0.008107f
C887 B.n747 VSUBS 0.008107f
C888 B.n748 VSUBS 0.008107f
C889 B.n749 VSUBS 0.008107f
C890 B.n750 VSUBS 0.008107f
C891 B.n751 VSUBS 0.008107f
C892 B.n752 VSUBS 0.008107f
C893 B.n753 VSUBS 0.008107f
C894 B.n754 VSUBS 0.008107f
C895 B.n755 VSUBS 0.008107f
C896 B.n756 VSUBS 0.008107f
C897 B.n757 VSUBS 0.008107f
C898 B.n758 VSUBS 0.008107f
C899 B.n759 VSUBS 0.008107f
C900 B.n760 VSUBS 0.008107f
C901 B.n761 VSUBS 0.008107f
C902 B.n762 VSUBS 0.008107f
C903 B.n763 VSUBS 0.008107f
C904 B.n764 VSUBS 0.008107f
C905 B.n765 VSUBS 0.008107f
C906 B.n766 VSUBS 0.008107f
C907 B.n767 VSUBS 0.008107f
C908 B.n768 VSUBS 0.008107f
C909 B.n769 VSUBS 0.008107f
C910 B.n770 VSUBS 0.008107f
C911 B.n771 VSUBS 0.008107f
C912 B.n772 VSUBS 0.008107f
C913 B.n773 VSUBS 0.008107f
C914 B.n774 VSUBS 0.008107f
C915 B.n775 VSUBS 0.008107f
C916 B.n776 VSUBS 0.008107f
C917 B.n777 VSUBS 0.008107f
C918 B.n778 VSUBS 0.008107f
C919 B.n779 VSUBS 0.008107f
C920 B.n780 VSUBS 0.008107f
C921 B.n781 VSUBS 0.008107f
C922 B.n782 VSUBS 0.008107f
C923 B.n783 VSUBS 0.008107f
C924 B.n784 VSUBS 0.008107f
C925 B.n785 VSUBS 0.008107f
C926 B.n786 VSUBS 0.008107f
C927 B.n787 VSUBS 0.008107f
C928 B.n788 VSUBS 0.008107f
C929 B.n789 VSUBS 0.008107f
C930 B.n790 VSUBS 0.008107f
C931 B.n791 VSUBS 0.008107f
C932 B.n792 VSUBS 0.008107f
C933 B.n793 VSUBS 0.008107f
C934 B.n794 VSUBS 0.008107f
C935 B.n795 VSUBS 0.008107f
C936 B.n796 VSUBS 0.008107f
C937 B.n797 VSUBS 0.008107f
C938 B.n798 VSUBS 0.008107f
C939 B.n799 VSUBS 0.008107f
C940 B.n800 VSUBS 0.00763f
C941 B.n801 VSUBS 0.018782f
C942 B.n802 VSUBS 0.00453f
C943 B.n803 VSUBS 0.008107f
C944 B.n804 VSUBS 0.008107f
C945 B.n805 VSUBS 0.008107f
C946 B.n806 VSUBS 0.008107f
C947 B.n807 VSUBS 0.008107f
C948 B.n808 VSUBS 0.008107f
C949 B.n809 VSUBS 0.008107f
C950 B.n810 VSUBS 0.008107f
C951 B.n811 VSUBS 0.008107f
C952 B.n812 VSUBS 0.008107f
C953 B.n813 VSUBS 0.008107f
C954 B.n814 VSUBS 0.008107f
C955 B.n815 VSUBS 0.00453f
C956 B.n816 VSUBS 0.008107f
C957 B.n817 VSUBS 0.008107f
C958 B.n818 VSUBS 0.008107f
C959 B.n819 VSUBS 0.008107f
C960 B.n820 VSUBS 0.008107f
C961 B.n821 VSUBS 0.008107f
C962 B.n822 VSUBS 0.008107f
C963 B.n823 VSUBS 0.008107f
C964 B.n824 VSUBS 0.008107f
C965 B.n825 VSUBS 0.008107f
C966 B.n826 VSUBS 0.008107f
C967 B.n827 VSUBS 0.008107f
C968 B.n828 VSUBS 0.008107f
C969 B.n829 VSUBS 0.008107f
C970 B.n830 VSUBS 0.008107f
C971 B.n831 VSUBS 0.008107f
C972 B.n832 VSUBS 0.008107f
C973 B.n833 VSUBS 0.008107f
C974 B.n834 VSUBS 0.008107f
C975 B.n835 VSUBS 0.008107f
C976 B.n836 VSUBS 0.008107f
C977 B.n837 VSUBS 0.008107f
C978 B.n838 VSUBS 0.008107f
C979 B.n839 VSUBS 0.008107f
C980 B.n840 VSUBS 0.008107f
C981 B.n841 VSUBS 0.008107f
C982 B.n842 VSUBS 0.008107f
C983 B.n843 VSUBS 0.008107f
C984 B.n844 VSUBS 0.008107f
C985 B.n845 VSUBS 0.008107f
C986 B.n846 VSUBS 0.008107f
C987 B.n847 VSUBS 0.008107f
C988 B.n848 VSUBS 0.008107f
C989 B.n849 VSUBS 0.008107f
C990 B.n850 VSUBS 0.008107f
C991 B.n851 VSUBS 0.008107f
C992 B.n852 VSUBS 0.008107f
C993 B.n853 VSUBS 0.008107f
C994 B.n854 VSUBS 0.008107f
C995 B.n855 VSUBS 0.008107f
C996 B.n856 VSUBS 0.008107f
C997 B.n857 VSUBS 0.008107f
C998 B.n858 VSUBS 0.008107f
C999 B.n859 VSUBS 0.008107f
C1000 B.n860 VSUBS 0.008107f
C1001 B.n861 VSUBS 0.008107f
C1002 B.n862 VSUBS 0.008107f
C1003 B.n863 VSUBS 0.008107f
C1004 B.n864 VSUBS 0.008107f
C1005 B.n865 VSUBS 0.008107f
C1006 B.n866 VSUBS 0.008107f
C1007 B.n867 VSUBS 0.008107f
C1008 B.n868 VSUBS 0.008107f
C1009 B.n869 VSUBS 0.008107f
C1010 B.n870 VSUBS 0.008107f
C1011 B.n871 VSUBS 0.008107f
C1012 B.n872 VSUBS 0.008107f
C1013 B.n873 VSUBS 0.008107f
C1014 B.n874 VSUBS 0.008107f
C1015 B.n875 VSUBS 0.008107f
C1016 B.n876 VSUBS 0.008107f
C1017 B.n877 VSUBS 0.008107f
C1018 B.n878 VSUBS 0.008107f
C1019 B.n879 VSUBS 0.008107f
C1020 B.n880 VSUBS 0.008107f
C1021 B.n881 VSUBS 0.008107f
C1022 B.n882 VSUBS 0.008107f
C1023 B.n883 VSUBS 0.008107f
C1024 B.n884 VSUBS 0.020041f
C1025 B.n885 VSUBS 0.020041f
C1026 B.n886 VSUBS 0.019537f
C1027 B.n887 VSUBS 0.008107f
C1028 B.n888 VSUBS 0.008107f
C1029 B.n889 VSUBS 0.008107f
C1030 B.n890 VSUBS 0.008107f
C1031 B.n891 VSUBS 0.008107f
C1032 B.n892 VSUBS 0.008107f
C1033 B.n893 VSUBS 0.008107f
C1034 B.n894 VSUBS 0.008107f
C1035 B.n895 VSUBS 0.008107f
C1036 B.n896 VSUBS 0.008107f
C1037 B.n897 VSUBS 0.008107f
C1038 B.n898 VSUBS 0.008107f
C1039 B.n899 VSUBS 0.008107f
C1040 B.n900 VSUBS 0.008107f
C1041 B.n901 VSUBS 0.008107f
C1042 B.n902 VSUBS 0.008107f
C1043 B.n903 VSUBS 0.008107f
C1044 B.n904 VSUBS 0.008107f
C1045 B.n905 VSUBS 0.008107f
C1046 B.n906 VSUBS 0.008107f
C1047 B.n907 VSUBS 0.008107f
C1048 B.n908 VSUBS 0.008107f
C1049 B.n909 VSUBS 0.008107f
C1050 B.n910 VSUBS 0.008107f
C1051 B.n911 VSUBS 0.008107f
C1052 B.n912 VSUBS 0.008107f
C1053 B.n913 VSUBS 0.008107f
C1054 B.n914 VSUBS 0.008107f
C1055 B.n915 VSUBS 0.008107f
C1056 B.n916 VSUBS 0.008107f
C1057 B.n917 VSUBS 0.008107f
C1058 B.n918 VSUBS 0.008107f
C1059 B.n919 VSUBS 0.008107f
C1060 B.n920 VSUBS 0.008107f
C1061 B.n921 VSUBS 0.008107f
C1062 B.n922 VSUBS 0.008107f
C1063 B.n923 VSUBS 0.008107f
C1064 B.n924 VSUBS 0.008107f
C1065 B.n925 VSUBS 0.008107f
C1066 B.n926 VSUBS 0.008107f
C1067 B.n927 VSUBS 0.008107f
C1068 B.n928 VSUBS 0.008107f
C1069 B.n929 VSUBS 0.008107f
C1070 B.n930 VSUBS 0.008107f
C1071 B.n931 VSUBS 0.008107f
C1072 B.n932 VSUBS 0.008107f
C1073 B.n933 VSUBS 0.008107f
C1074 B.n934 VSUBS 0.008107f
C1075 B.n935 VSUBS 0.008107f
C1076 B.n936 VSUBS 0.008107f
C1077 B.n937 VSUBS 0.008107f
C1078 B.n938 VSUBS 0.008107f
C1079 B.n939 VSUBS 0.008107f
C1080 B.n940 VSUBS 0.008107f
C1081 B.n941 VSUBS 0.008107f
C1082 B.n942 VSUBS 0.008107f
C1083 B.n943 VSUBS 0.008107f
C1084 B.n944 VSUBS 0.008107f
C1085 B.n945 VSUBS 0.008107f
C1086 B.n946 VSUBS 0.008107f
C1087 B.n947 VSUBS 0.008107f
C1088 B.n948 VSUBS 0.008107f
C1089 B.n949 VSUBS 0.008107f
C1090 B.n950 VSUBS 0.008107f
C1091 B.n951 VSUBS 0.008107f
C1092 B.n952 VSUBS 0.008107f
C1093 B.n953 VSUBS 0.008107f
C1094 B.n954 VSUBS 0.008107f
C1095 B.n955 VSUBS 0.008107f
C1096 B.n956 VSUBS 0.008107f
C1097 B.n957 VSUBS 0.008107f
C1098 B.n958 VSUBS 0.008107f
C1099 B.n959 VSUBS 0.008107f
C1100 B.n960 VSUBS 0.008107f
C1101 B.n961 VSUBS 0.008107f
C1102 B.n962 VSUBS 0.008107f
C1103 B.n963 VSUBS 0.008107f
C1104 B.n964 VSUBS 0.008107f
C1105 B.n965 VSUBS 0.008107f
C1106 B.n966 VSUBS 0.008107f
C1107 B.n967 VSUBS 0.008107f
C1108 B.n968 VSUBS 0.008107f
C1109 B.n969 VSUBS 0.008107f
C1110 B.n970 VSUBS 0.008107f
C1111 B.n971 VSUBS 0.008107f
C1112 B.n972 VSUBS 0.008107f
C1113 B.n973 VSUBS 0.008107f
C1114 B.n974 VSUBS 0.008107f
C1115 B.n975 VSUBS 0.008107f
C1116 B.n976 VSUBS 0.008107f
C1117 B.n977 VSUBS 0.008107f
C1118 B.n978 VSUBS 0.008107f
C1119 B.n979 VSUBS 0.008107f
C1120 B.n980 VSUBS 0.008107f
C1121 B.n981 VSUBS 0.008107f
C1122 B.n982 VSUBS 0.008107f
C1123 B.n983 VSUBS 0.008107f
C1124 B.n984 VSUBS 0.008107f
C1125 B.n985 VSUBS 0.008107f
C1126 B.n986 VSUBS 0.008107f
C1127 B.n987 VSUBS 0.008107f
C1128 B.n988 VSUBS 0.008107f
C1129 B.n989 VSUBS 0.008107f
C1130 B.n990 VSUBS 0.008107f
C1131 B.n991 VSUBS 0.010579f
C1132 B.n992 VSUBS 0.011269f
C1133 B.n993 VSUBS 0.022409f
C1134 VTAIL.t2 VSUBS 0.276713f
C1135 VTAIL.t1 VSUBS 0.276713f
C1136 VTAIL.n0 VSUBS 2.08075f
C1137 VTAIL.n1 VSUBS 0.894813f
C1138 VTAIL.t6 VSUBS 2.73189f
C1139 VTAIL.n2 VSUBS 1.03239f
C1140 VTAIL.t9 VSUBS 2.73189f
C1141 VTAIL.n3 VSUBS 1.03239f
C1142 VTAIL.t11 VSUBS 0.276713f
C1143 VTAIL.t13 VSUBS 0.276713f
C1144 VTAIL.n4 VSUBS 2.08075f
C1145 VTAIL.n5 VSUBS 1.19735f
C1146 VTAIL.t8 VSUBS 2.73189f
C1147 VTAIL.n6 VSUBS 2.62229f
C1148 VTAIL.t3 VSUBS 2.7319f
C1149 VTAIL.n7 VSUBS 2.62229f
C1150 VTAIL.t7 VSUBS 0.276713f
C1151 VTAIL.t5 VSUBS 0.276713f
C1152 VTAIL.n8 VSUBS 2.08075f
C1153 VTAIL.n9 VSUBS 1.19735f
C1154 VTAIL.t4 VSUBS 2.7319f
C1155 VTAIL.n10 VSUBS 1.03239f
C1156 VTAIL.t14 VSUBS 2.7319f
C1157 VTAIL.n11 VSUBS 1.03239f
C1158 VTAIL.t10 VSUBS 0.276713f
C1159 VTAIL.t15 VSUBS 0.276713f
C1160 VTAIL.n12 VSUBS 2.08075f
C1161 VTAIL.n13 VSUBS 1.19735f
C1162 VTAIL.t12 VSUBS 2.7319f
C1163 VTAIL.n14 VSUBS 2.62229f
C1164 VTAIL.t0 VSUBS 2.73189f
C1165 VTAIL.n15 VSUBS 2.61748f
C1166 VDD1.t0 VSUBS 0.354701f
C1167 VDD1.t6 VSUBS 0.354701f
C1168 VDD1.n0 VSUBS 2.87734f
C1169 VDD1.t2 VSUBS 0.354701f
C1170 VDD1.t7 VSUBS 0.354701f
C1171 VDD1.n1 VSUBS 2.87525f
C1172 VDD1.t5 VSUBS 0.354701f
C1173 VDD1.t3 VSUBS 0.354701f
C1174 VDD1.n2 VSUBS 2.87525f
C1175 VDD1.n3 VSUBS 6.24242f
C1176 VDD1.t1 VSUBS 0.354701f
C1177 VDD1.t4 VSUBS 0.354701f
C1178 VDD1.n4 VSUBS 2.84613f
C1179 VDD1.n5 VSUBS 5.0602f
C1180 VP.n0 VSUBS 0.045775f
C1181 VP.t6 VSUBS 3.61083f
C1182 VP.n1 VSUBS 0.045569f
C1183 VP.n2 VSUBS 0.024328f
C1184 VP.n3 VSUBS 0.045569f
C1185 VP.n4 VSUBS 0.024328f
C1186 VP.t2 VSUBS 3.61083f
C1187 VP.n5 VSUBS 0.045569f
C1188 VP.n6 VSUBS 0.024328f
C1189 VP.n7 VSUBS 0.045569f
C1190 VP.n8 VSUBS 0.024328f
C1191 VP.t4 VSUBS 3.61083f
C1192 VP.n9 VSUBS 0.045569f
C1193 VP.n10 VSUBS 0.024328f
C1194 VP.n11 VSUBS 0.045569f
C1195 VP.n12 VSUBS 0.045775f
C1196 VP.t7 VSUBS 3.61083f
C1197 VP.n13 VSUBS 0.045775f
C1198 VP.t3 VSUBS 3.61083f
C1199 VP.n14 VSUBS 0.045569f
C1200 VP.n15 VSUBS 0.024328f
C1201 VP.n16 VSUBS 0.045569f
C1202 VP.n17 VSUBS 0.024328f
C1203 VP.t0 VSUBS 3.61083f
C1204 VP.n18 VSUBS 0.045569f
C1205 VP.n19 VSUBS 0.024328f
C1206 VP.n20 VSUBS 0.045569f
C1207 VP.n21 VSUBS 0.322391f
C1208 VP.t5 VSUBS 3.61083f
C1209 VP.t1 VSUBS 4.01683f
C1210 VP.n22 VSUBS 1.28087f
C1211 VP.n23 VSUBS 1.34168f
C1212 VP.n24 VSUBS 0.030045f
C1213 VP.n25 VSUBS 0.045569f
C1214 VP.n26 VSUBS 0.024328f
C1215 VP.n27 VSUBS 0.024328f
C1216 VP.n28 VSUBS 0.024328f
C1217 VP.n29 VSUBS 0.048611f
C1218 VP.n30 VSUBS 0.019687f
C1219 VP.n31 VSUBS 0.048611f
C1220 VP.n32 VSUBS 0.024328f
C1221 VP.n33 VSUBS 0.024328f
C1222 VP.n34 VSUBS 0.024328f
C1223 VP.n35 VSUBS 0.045569f
C1224 VP.n36 VSUBS 0.030045f
C1225 VP.n37 VSUBS 1.25626f
C1226 VP.n38 VSUBS 0.038594f
C1227 VP.n39 VSUBS 0.024328f
C1228 VP.n40 VSUBS 0.024328f
C1229 VP.n41 VSUBS 0.024328f
C1230 VP.n42 VSUBS 0.045569f
C1231 VP.n43 VSUBS 0.039766f
C1232 VP.n44 VSUBS 0.031573f
C1233 VP.n45 VSUBS 0.024328f
C1234 VP.n46 VSUBS 0.024328f
C1235 VP.n47 VSUBS 0.024328f
C1236 VP.n48 VSUBS 0.045569f
C1237 VP.n49 VSUBS 0.043994f
C1238 VP.n50 VSUBS 1.36837f
C1239 VP.n51 VSUBS 1.76754f
C1240 VP.n52 VSUBS 1.78235f
C1241 VP.n53 VSUBS 1.36837f
C1242 VP.n54 VSUBS 0.043994f
C1243 VP.n55 VSUBS 0.045569f
C1244 VP.n56 VSUBS 0.024328f
C1245 VP.n57 VSUBS 0.024328f
C1246 VP.n58 VSUBS 0.024328f
C1247 VP.n59 VSUBS 0.031573f
C1248 VP.n60 VSUBS 0.039766f
C1249 VP.n61 VSUBS 0.045569f
C1250 VP.n62 VSUBS 0.024328f
C1251 VP.n63 VSUBS 0.024328f
C1252 VP.n64 VSUBS 0.024328f
C1253 VP.n65 VSUBS 0.038594f
C1254 VP.n66 VSUBS 1.25626f
C1255 VP.n67 VSUBS 0.030045f
C1256 VP.n68 VSUBS 0.045569f
C1257 VP.n69 VSUBS 0.024328f
C1258 VP.n70 VSUBS 0.024328f
C1259 VP.n71 VSUBS 0.024328f
C1260 VP.n72 VSUBS 0.048611f
C1261 VP.n73 VSUBS 0.019687f
C1262 VP.n74 VSUBS 0.048611f
C1263 VP.n75 VSUBS 0.024328f
C1264 VP.n76 VSUBS 0.024328f
C1265 VP.n77 VSUBS 0.024328f
C1266 VP.n78 VSUBS 0.045569f
C1267 VP.n79 VSUBS 0.030045f
C1268 VP.n80 VSUBS 1.25626f
C1269 VP.n81 VSUBS 0.038594f
C1270 VP.n82 VSUBS 0.024328f
C1271 VP.n83 VSUBS 0.024328f
C1272 VP.n84 VSUBS 0.024328f
C1273 VP.n85 VSUBS 0.045569f
C1274 VP.n86 VSUBS 0.039766f
C1275 VP.n87 VSUBS 0.031573f
C1276 VP.n88 VSUBS 0.024328f
C1277 VP.n89 VSUBS 0.024328f
C1278 VP.n90 VSUBS 0.024328f
C1279 VP.n91 VSUBS 0.045569f
C1280 VP.n92 VSUBS 0.043994f
C1281 VP.n93 VSUBS 1.36837f
C1282 VP.n94 VSUBS 0.074188f
.ends

