* NGSPICE file created from diff_pair_sample_0826.ext - technology: sky130A

.subckt diff_pair_sample_0826 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=2.5467 ps=13.84 w=6.53 l=2.28
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=2.5467 ps=13.84 w=6.53 l=2.28
X2 B.t11 B.t9 B.t10 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=2.28
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=2.5467 ps=13.84 w=6.53 l=2.28
X4 B.t8 B.t6 B.t7 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=2.28
X5 B.t5 B.t3 B.t4 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=2.28
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=2.5467 ps=13.84 w=6.53 l=2.28
X7 B.t2 B.t0 B.t1 w_n2014_n2274# sky130_fd_pr__pfet_01v8 ad=2.5467 pd=13.84 as=0 ps=0 w=6.53 l=2.28
R0 VN VN.t1 157.954
R1 VN VN.t0 118.531
R2 VTAIL.n134 VTAIL.n133 756.745
R3 VTAIL.n32 VTAIL.n31 756.745
R4 VTAIL.n100 VTAIL.n99 756.745
R5 VTAIL.n66 VTAIL.n65 756.745
R6 VTAIL.n112 VTAIL.n111 585
R7 VTAIL.n117 VTAIL.n116 585
R8 VTAIL.n119 VTAIL.n118 585
R9 VTAIL.n108 VTAIL.n107 585
R10 VTAIL.n125 VTAIL.n124 585
R11 VTAIL.n127 VTAIL.n126 585
R12 VTAIL.n104 VTAIL.n103 585
R13 VTAIL.n133 VTAIL.n132 585
R14 VTAIL.n10 VTAIL.n9 585
R15 VTAIL.n15 VTAIL.n14 585
R16 VTAIL.n17 VTAIL.n16 585
R17 VTAIL.n6 VTAIL.n5 585
R18 VTAIL.n23 VTAIL.n22 585
R19 VTAIL.n25 VTAIL.n24 585
R20 VTAIL.n2 VTAIL.n1 585
R21 VTAIL.n31 VTAIL.n30 585
R22 VTAIL.n99 VTAIL.n98 585
R23 VTAIL.n70 VTAIL.n69 585
R24 VTAIL.n93 VTAIL.n92 585
R25 VTAIL.n91 VTAIL.n90 585
R26 VTAIL.n74 VTAIL.n73 585
R27 VTAIL.n85 VTAIL.n84 585
R28 VTAIL.n83 VTAIL.n82 585
R29 VTAIL.n78 VTAIL.n77 585
R30 VTAIL.n65 VTAIL.n64 585
R31 VTAIL.n36 VTAIL.n35 585
R32 VTAIL.n59 VTAIL.n58 585
R33 VTAIL.n57 VTAIL.n56 585
R34 VTAIL.n40 VTAIL.n39 585
R35 VTAIL.n51 VTAIL.n50 585
R36 VTAIL.n49 VTAIL.n48 585
R37 VTAIL.n44 VTAIL.n43 585
R38 VTAIL.n113 VTAIL.t3 329.084
R39 VTAIL.n11 VTAIL.t1 329.084
R40 VTAIL.n79 VTAIL.t0 329.084
R41 VTAIL.n45 VTAIL.t2 329.084
R42 VTAIL.n117 VTAIL.n111 171.744
R43 VTAIL.n118 VTAIL.n117 171.744
R44 VTAIL.n118 VTAIL.n107 171.744
R45 VTAIL.n125 VTAIL.n107 171.744
R46 VTAIL.n126 VTAIL.n125 171.744
R47 VTAIL.n126 VTAIL.n103 171.744
R48 VTAIL.n133 VTAIL.n103 171.744
R49 VTAIL.n15 VTAIL.n9 171.744
R50 VTAIL.n16 VTAIL.n15 171.744
R51 VTAIL.n16 VTAIL.n5 171.744
R52 VTAIL.n23 VTAIL.n5 171.744
R53 VTAIL.n24 VTAIL.n23 171.744
R54 VTAIL.n24 VTAIL.n1 171.744
R55 VTAIL.n31 VTAIL.n1 171.744
R56 VTAIL.n99 VTAIL.n69 171.744
R57 VTAIL.n92 VTAIL.n69 171.744
R58 VTAIL.n92 VTAIL.n91 171.744
R59 VTAIL.n91 VTAIL.n73 171.744
R60 VTAIL.n84 VTAIL.n73 171.744
R61 VTAIL.n84 VTAIL.n83 171.744
R62 VTAIL.n83 VTAIL.n77 171.744
R63 VTAIL.n65 VTAIL.n35 171.744
R64 VTAIL.n58 VTAIL.n35 171.744
R65 VTAIL.n58 VTAIL.n57 171.744
R66 VTAIL.n57 VTAIL.n39 171.744
R67 VTAIL.n50 VTAIL.n39 171.744
R68 VTAIL.n50 VTAIL.n49 171.744
R69 VTAIL.n49 VTAIL.n43 171.744
R70 VTAIL.t3 VTAIL.n111 85.8723
R71 VTAIL.t1 VTAIL.n9 85.8723
R72 VTAIL.t0 VTAIL.n77 85.8723
R73 VTAIL.t2 VTAIL.n43 85.8723
R74 VTAIL.n135 VTAIL.n134 35.0944
R75 VTAIL.n33 VTAIL.n32 35.0944
R76 VTAIL.n101 VTAIL.n100 35.0944
R77 VTAIL.n67 VTAIL.n66 35.0944
R78 VTAIL.n67 VTAIL.n33 22.4962
R79 VTAIL.n135 VTAIL.n101 20.2462
R80 VTAIL.n132 VTAIL.n102 12.8005
R81 VTAIL.n30 VTAIL.n0 12.8005
R82 VTAIL.n98 VTAIL.n68 12.8005
R83 VTAIL.n64 VTAIL.n34 12.8005
R84 VTAIL.n131 VTAIL.n104 12.0247
R85 VTAIL.n29 VTAIL.n2 12.0247
R86 VTAIL.n97 VTAIL.n70 12.0247
R87 VTAIL.n63 VTAIL.n36 12.0247
R88 VTAIL.n128 VTAIL.n127 11.249
R89 VTAIL.n26 VTAIL.n25 11.249
R90 VTAIL.n94 VTAIL.n93 11.249
R91 VTAIL.n60 VTAIL.n59 11.249
R92 VTAIL.n113 VTAIL.n112 10.7233
R93 VTAIL.n11 VTAIL.n10 10.7233
R94 VTAIL.n79 VTAIL.n78 10.7233
R95 VTAIL.n45 VTAIL.n44 10.7233
R96 VTAIL.n124 VTAIL.n106 10.4732
R97 VTAIL.n22 VTAIL.n4 10.4732
R98 VTAIL.n90 VTAIL.n72 10.4732
R99 VTAIL.n56 VTAIL.n38 10.4732
R100 VTAIL.n123 VTAIL.n108 9.69747
R101 VTAIL.n21 VTAIL.n6 9.69747
R102 VTAIL.n89 VTAIL.n74 9.69747
R103 VTAIL.n55 VTAIL.n40 9.69747
R104 VTAIL.n130 VTAIL.n102 9.45567
R105 VTAIL.n28 VTAIL.n0 9.45567
R106 VTAIL.n96 VTAIL.n68 9.45567
R107 VTAIL.n62 VTAIL.n34 9.45567
R108 VTAIL.n115 VTAIL.n114 9.3005
R109 VTAIL.n110 VTAIL.n109 9.3005
R110 VTAIL.n121 VTAIL.n120 9.3005
R111 VTAIL.n123 VTAIL.n122 9.3005
R112 VTAIL.n106 VTAIL.n105 9.3005
R113 VTAIL.n129 VTAIL.n128 9.3005
R114 VTAIL.n131 VTAIL.n130 9.3005
R115 VTAIL.n13 VTAIL.n12 9.3005
R116 VTAIL.n8 VTAIL.n7 9.3005
R117 VTAIL.n19 VTAIL.n18 9.3005
R118 VTAIL.n21 VTAIL.n20 9.3005
R119 VTAIL.n4 VTAIL.n3 9.3005
R120 VTAIL.n27 VTAIL.n26 9.3005
R121 VTAIL.n29 VTAIL.n28 9.3005
R122 VTAIL.n97 VTAIL.n96 9.3005
R123 VTAIL.n95 VTAIL.n94 9.3005
R124 VTAIL.n72 VTAIL.n71 9.3005
R125 VTAIL.n89 VTAIL.n88 9.3005
R126 VTAIL.n87 VTAIL.n86 9.3005
R127 VTAIL.n76 VTAIL.n75 9.3005
R128 VTAIL.n81 VTAIL.n80 9.3005
R129 VTAIL.n42 VTAIL.n41 9.3005
R130 VTAIL.n53 VTAIL.n52 9.3005
R131 VTAIL.n55 VTAIL.n54 9.3005
R132 VTAIL.n38 VTAIL.n37 9.3005
R133 VTAIL.n61 VTAIL.n60 9.3005
R134 VTAIL.n63 VTAIL.n62 9.3005
R135 VTAIL.n47 VTAIL.n46 9.3005
R136 VTAIL.n120 VTAIL.n119 8.92171
R137 VTAIL.n18 VTAIL.n17 8.92171
R138 VTAIL.n86 VTAIL.n85 8.92171
R139 VTAIL.n52 VTAIL.n51 8.92171
R140 VTAIL.n116 VTAIL.n110 8.14595
R141 VTAIL.n14 VTAIL.n8 8.14595
R142 VTAIL.n82 VTAIL.n76 8.14595
R143 VTAIL.n48 VTAIL.n42 8.14595
R144 VTAIL.n115 VTAIL.n112 7.3702
R145 VTAIL.n13 VTAIL.n10 7.3702
R146 VTAIL.n81 VTAIL.n78 7.3702
R147 VTAIL.n47 VTAIL.n44 7.3702
R148 VTAIL.n116 VTAIL.n115 5.81868
R149 VTAIL.n14 VTAIL.n13 5.81868
R150 VTAIL.n82 VTAIL.n81 5.81868
R151 VTAIL.n48 VTAIL.n47 5.81868
R152 VTAIL.n119 VTAIL.n110 5.04292
R153 VTAIL.n17 VTAIL.n8 5.04292
R154 VTAIL.n85 VTAIL.n76 5.04292
R155 VTAIL.n51 VTAIL.n42 5.04292
R156 VTAIL.n120 VTAIL.n108 4.26717
R157 VTAIL.n18 VTAIL.n6 4.26717
R158 VTAIL.n86 VTAIL.n74 4.26717
R159 VTAIL.n52 VTAIL.n40 4.26717
R160 VTAIL.n124 VTAIL.n123 3.49141
R161 VTAIL.n22 VTAIL.n21 3.49141
R162 VTAIL.n90 VTAIL.n89 3.49141
R163 VTAIL.n56 VTAIL.n55 3.49141
R164 VTAIL.n127 VTAIL.n106 2.71565
R165 VTAIL.n25 VTAIL.n4 2.71565
R166 VTAIL.n93 VTAIL.n72 2.71565
R167 VTAIL.n59 VTAIL.n38 2.71565
R168 VTAIL.n46 VTAIL.n45 2.41347
R169 VTAIL.n114 VTAIL.n113 2.41347
R170 VTAIL.n12 VTAIL.n11 2.41347
R171 VTAIL.n80 VTAIL.n79 2.41347
R172 VTAIL.n128 VTAIL.n104 1.93989
R173 VTAIL.n26 VTAIL.n2 1.93989
R174 VTAIL.n94 VTAIL.n70 1.93989
R175 VTAIL.n60 VTAIL.n36 1.93989
R176 VTAIL.n101 VTAIL.n67 1.59533
R177 VTAIL.n132 VTAIL.n131 1.16414
R178 VTAIL.n30 VTAIL.n29 1.16414
R179 VTAIL.n98 VTAIL.n97 1.16414
R180 VTAIL.n64 VTAIL.n63 1.16414
R181 VTAIL VTAIL.n33 1.09102
R182 VTAIL VTAIL.n135 0.50481
R183 VTAIL.n134 VTAIL.n102 0.388379
R184 VTAIL.n32 VTAIL.n0 0.388379
R185 VTAIL.n100 VTAIL.n68 0.388379
R186 VTAIL.n66 VTAIL.n34 0.388379
R187 VTAIL.n114 VTAIL.n109 0.155672
R188 VTAIL.n121 VTAIL.n109 0.155672
R189 VTAIL.n122 VTAIL.n121 0.155672
R190 VTAIL.n122 VTAIL.n105 0.155672
R191 VTAIL.n129 VTAIL.n105 0.155672
R192 VTAIL.n130 VTAIL.n129 0.155672
R193 VTAIL.n12 VTAIL.n7 0.155672
R194 VTAIL.n19 VTAIL.n7 0.155672
R195 VTAIL.n20 VTAIL.n19 0.155672
R196 VTAIL.n20 VTAIL.n3 0.155672
R197 VTAIL.n27 VTAIL.n3 0.155672
R198 VTAIL.n28 VTAIL.n27 0.155672
R199 VTAIL.n96 VTAIL.n95 0.155672
R200 VTAIL.n95 VTAIL.n71 0.155672
R201 VTAIL.n88 VTAIL.n71 0.155672
R202 VTAIL.n88 VTAIL.n87 0.155672
R203 VTAIL.n87 VTAIL.n75 0.155672
R204 VTAIL.n80 VTAIL.n75 0.155672
R205 VTAIL.n62 VTAIL.n61 0.155672
R206 VTAIL.n61 VTAIL.n37 0.155672
R207 VTAIL.n54 VTAIL.n37 0.155672
R208 VTAIL.n54 VTAIL.n53 0.155672
R209 VTAIL.n53 VTAIL.n41 0.155672
R210 VTAIL.n46 VTAIL.n41 0.155672
R211 VDD2.n65 VDD2.n64 756.745
R212 VDD2.n32 VDD2.n31 756.745
R213 VDD2.n64 VDD2.n63 585
R214 VDD2.n35 VDD2.n34 585
R215 VDD2.n58 VDD2.n57 585
R216 VDD2.n56 VDD2.n55 585
R217 VDD2.n39 VDD2.n38 585
R218 VDD2.n50 VDD2.n49 585
R219 VDD2.n48 VDD2.n47 585
R220 VDD2.n43 VDD2.n42 585
R221 VDD2.n10 VDD2.n9 585
R222 VDD2.n15 VDD2.n14 585
R223 VDD2.n17 VDD2.n16 585
R224 VDD2.n6 VDD2.n5 585
R225 VDD2.n23 VDD2.n22 585
R226 VDD2.n25 VDD2.n24 585
R227 VDD2.n2 VDD2.n1 585
R228 VDD2.n31 VDD2.n30 585
R229 VDD2.n44 VDD2.t0 329.084
R230 VDD2.n11 VDD2.t1 329.084
R231 VDD2.n64 VDD2.n34 171.744
R232 VDD2.n57 VDD2.n34 171.744
R233 VDD2.n57 VDD2.n56 171.744
R234 VDD2.n56 VDD2.n38 171.744
R235 VDD2.n49 VDD2.n38 171.744
R236 VDD2.n49 VDD2.n48 171.744
R237 VDD2.n48 VDD2.n42 171.744
R238 VDD2.n15 VDD2.n9 171.744
R239 VDD2.n16 VDD2.n15 171.744
R240 VDD2.n16 VDD2.n5 171.744
R241 VDD2.n23 VDD2.n5 171.744
R242 VDD2.n24 VDD2.n23 171.744
R243 VDD2.n24 VDD2.n1 171.744
R244 VDD2.n31 VDD2.n1 171.744
R245 VDD2.t0 VDD2.n42 85.8723
R246 VDD2.t1 VDD2.n9 85.8723
R247 VDD2.n66 VDD2.n32 85.562
R248 VDD2.n66 VDD2.n65 51.7732
R249 VDD2.n63 VDD2.n33 12.8005
R250 VDD2.n30 VDD2.n0 12.8005
R251 VDD2.n62 VDD2.n35 12.0247
R252 VDD2.n29 VDD2.n2 12.0247
R253 VDD2.n59 VDD2.n58 11.249
R254 VDD2.n26 VDD2.n25 11.249
R255 VDD2.n44 VDD2.n43 10.7233
R256 VDD2.n11 VDD2.n10 10.7233
R257 VDD2.n55 VDD2.n37 10.4732
R258 VDD2.n22 VDD2.n4 10.4732
R259 VDD2.n54 VDD2.n39 9.69747
R260 VDD2.n21 VDD2.n6 9.69747
R261 VDD2.n61 VDD2.n33 9.45567
R262 VDD2.n28 VDD2.n0 9.45567
R263 VDD2.n62 VDD2.n61 9.3005
R264 VDD2.n60 VDD2.n59 9.3005
R265 VDD2.n37 VDD2.n36 9.3005
R266 VDD2.n54 VDD2.n53 9.3005
R267 VDD2.n52 VDD2.n51 9.3005
R268 VDD2.n41 VDD2.n40 9.3005
R269 VDD2.n46 VDD2.n45 9.3005
R270 VDD2.n13 VDD2.n12 9.3005
R271 VDD2.n8 VDD2.n7 9.3005
R272 VDD2.n19 VDD2.n18 9.3005
R273 VDD2.n21 VDD2.n20 9.3005
R274 VDD2.n4 VDD2.n3 9.3005
R275 VDD2.n27 VDD2.n26 9.3005
R276 VDD2.n29 VDD2.n28 9.3005
R277 VDD2.n51 VDD2.n50 8.92171
R278 VDD2.n18 VDD2.n17 8.92171
R279 VDD2.n47 VDD2.n41 8.14595
R280 VDD2.n14 VDD2.n8 8.14595
R281 VDD2.n46 VDD2.n43 7.3702
R282 VDD2.n13 VDD2.n10 7.3702
R283 VDD2.n47 VDD2.n46 5.81868
R284 VDD2.n14 VDD2.n13 5.81868
R285 VDD2.n50 VDD2.n41 5.04292
R286 VDD2.n17 VDD2.n8 5.04292
R287 VDD2.n51 VDD2.n39 4.26717
R288 VDD2.n18 VDD2.n6 4.26717
R289 VDD2.n55 VDD2.n54 3.49141
R290 VDD2.n22 VDD2.n21 3.49141
R291 VDD2.n58 VDD2.n37 2.71565
R292 VDD2.n25 VDD2.n4 2.71565
R293 VDD2.n45 VDD2.n44 2.41347
R294 VDD2.n12 VDD2.n11 2.41347
R295 VDD2.n59 VDD2.n35 1.93989
R296 VDD2.n26 VDD2.n2 1.93989
R297 VDD2.n63 VDD2.n62 1.16414
R298 VDD2.n30 VDD2.n29 1.16414
R299 VDD2 VDD2.n66 0.62119
R300 VDD2.n65 VDD2.n33 0.388379
R301 VDD2.n32 VDD2.n0 0.388379
R302 VDD2.n61 VDD2.n60 0.155672
R303 VDD2.n60 VDD2.n36 0.155672
R304 VDD2.n53 VDD2.n36 0.155672
R305 VDD2.n53 VDD2.n52 0.155672
R306 VDD2.n52 VDD2.n40 0.155672
R307 VDD2.n45 VDD2.n40 0.155672
R308 VDD2.n12 VDD2.n7 0.155672
R309 VDD2.n19 VDD2.n7 0.155672
R310 VDD2.n20 VDD2.n19 0.155672
R311 VDD2.n20 VDD2.n3 0.155672
R312 VDD2.n27 VDD2.n3 0.155672
R313 VDD2.n28 VDD2.n27 0.155672
R314 VP.n0 VP.t1 157.858
R315 VP.n0 VP.t0 118.195
R316 VP VP.n0 0.336784
R317 VDD1.n32 VDD1.n31 756.745
R318 VDD1.n65 VDD1.n64 756.745
R319 VDD1.n31 VDD1.n30 585
R320 VDD1.n2 VDD1.n1 585
R321 VDD1.n25 VDD1.n24 585
R322 VDD1.n23 VDD1.n22 585
R323 VDD1.n6 VDD1.n5 585
R324 VDD1.n17 VDD1.n16 585
R325 VDD1.n15 VDD1.n14 585
R326 VDD1.n10 VDD1.n9 585
R327 VDD1.n43 VDD1.n42 585
R328 VDD1.n48 VDD1.n47 585
R329 VDD1.n50 VDD1.n49 585
R330 VDD1.n39 VDD1.n38 585
R331 VDD1.n56 VDD1.n55 585
R332 VDD1.n58 VDD1.n57 585
R333 VDD1.n35 VDD1.n34 585
R334 VDD1.n64 VDD1.n63 585
R335 VDD1.n11 VDD1.t0 329.084
R336 VDD1.n44 VDD1.t1 329.084
R337 VDD1.n31 VDD1.n1 171.744
R338 VDD1.n24 VDD1.n1 171.744
R339 VDD1.n24 VDD1.n23 171.744
R340 VDD1.n23 VDD1.n5 171.744
R341 VDD1.n16 VDD1.n5 171.744
R342 VDD1.n16 VDD1.n15 171.744
R343 VDD1.n15 VDD1.n9 171.744
R344 VDD1.n48 VDD1.n42 171.744
R345 VDD1.n49 VDD1.n48 171.744
R346 VDD1.n49 VDD1.n38 171.744
R347 VDD1.n56 VDD1.n38 171.744
R348 VDD1.n57 VDD1.n56 171.744
R349 VDD1.n57 VDD1.n34 171.744
R350 VDD1.n64 VDD1.n34 171.744
R351 VDD1 VDD1.n65 86.6493
R352 VDD1.t0 VDD1.n9 85.8723
R353 VDD1.t1 VDD1.n42 85.8723
R354 VDD1 VDD1.n32 52.3939
R355 VDD1.n30 VDD1.n0 12.8005
R356 VDD1.n63 VDD1.n33 12.8005
R357 VDD1.n29 VDD1.n2 12.0247
R358 VDD1.n62 VDD1.n35 12.0247
R359 VDD1.n26 VDD1.n25 11.249
R360 VDD1.n59 VDD1.n58 11.249
R361 VDD1.n11 VDD1.n10 10.7233
R362 VDD1.n44 VDD1.n43 10.7233
R363 VDD1.n22 VDD1.n4 10.4732
R364 VDD1.n55 VDD1.n37 10.4732
R365 VDD1.n21 VDD1.n6 9.69747
R366 VDD1.n54 VDD1.n39 9.69747
R367 VDD1.n28 VDD1.n0 9.45567
R368 VDD1.n61 VDD1.n33 9.45567
R369 VDD1.n29 VDD1.n28 9.3005
R370 VDD1.n27 VDD1.n26 9.3005
R371 VDD1.n4 VDD1.n3 9.3005
R372 VDD1.n21 VDD1.n20 9.3005
R373 VDD1.n19 VDD1.n18 9.3005
R374 VDD1.n8 VDD1.n7 9.3005
R375 VDD1.n13 VDD1.n12 9.3005
R376 VDD1.n46 VDD1.n45 9.3005
R377 VDD1.n41 VDD1.n40 9.3005
R378 VDD1.n52 VDD1.n51 9.3005
R379 VDD1.n54 VDD1.n53 9.3005
R380 VDD1.n37 VDD1.n36 9.3005
R381 VDD1.n60 VDD1.n59 9.3005
R382 VDD1.n62 VDD1.n61 9.3005
R383 VDD1.n18 VDD1.n17 8.92171
R384 VDD1.n51 VDD1.n50 8.92171
R385 VDD1.n14 VDD1.n8 8.14595
R386 VDD1.n47 VDD1.n41 8.14595
R387 VDD1.n13 VDD1.n10 7.3702
R388 VDD1.n46 VDD1.n43 7.3702
R389 VDD1.n14 VDD1.n13 5.81868
R390 VDD1.n47 VDD1.n46 5.81868
R391 VDD1.n17 VDD1.n8 5.04292
R392 VDD1.n50 VDD1.n41 5.04292
R393 VDD1.n18 VDD1.n6 4.26717
R394 VDD1.n51 VDD1.n39 4.26717
R395 VDD1.n22 VDD1.n21 3.49141
R396 VDD1.n55 VDD1.n54 3.49141
R397 VDD1.n25 VDD1.n4 2.71565
R398 VDD1.n58 VDD1.n37 2.71565
R399 VDD1.n12 VDD1.n11 2.41347
R400 VDD1.n45 VDD1.n44 2.41347
R401 VDD1.n26 VDD1.n2 1.93989
R402 VDD1.n59 VDD1.n35 1.93989
R403 VDD1.n30 VDD1.n29 1.16414
R404 VDD1.n63 VDD1.n62 1.16414
R405 VDD1.n32 VDD1.n0 0.388379
R406 VDD1.n65 VDD1.n33 0.388379
R407 VDD1.n28 VDD1.n27 0.155672
R408 VDD1.n27 VDD1.n3 0.155672
R409 VDD1.n20 VDD1.n3 0.155672
R410 VDD1.n20 VDD1.n19 0.155672
R411 VDD1.n19 VDD1.n7 0.155672
R412 VDD1.n12 VDD1.n7 0.155672
R413 VDD1.n45 VDD1.n40 0.155672
R414 VDD1.n52 VDD1.n40 0.155672
R415 VDD1.n53 VDD1.n52 0.155672
R416 VDD1.n53 VDD1.n36 0.155672
R417 VDD1.n60 VDD1.n36 0.155672
R418 VDD1.n61 VDD1.n60 0.155672
R419 B.n244 B.n73 585
R420 B.n243 B.n242 585
R421 B.n241 B.n74 585
R422 B.n240 B.n239 585
R423 B.n238 B.n75 585
R424 B.n237 B.n236 585
R425 B.n235 B.n76 585
R426 B.n234 B.n233 585
R427 B.n232 B.n77 585
R428 B.n231 B.n230 585
R429 B.n229 B.n78 585
R430 B.n228 B.n227 585
R431 B.n226 B.n79 585
R432 B.n225 B.n224 585
R433 B.n223 B.n80 585
R434 B.n222 B.n221 585
R435 B.n220 B.n81 585
R436 B.n219 B.n218 585
R437 B.n217 B.n82 585
R438 B.n216 B.n215 585
R439 B.n214 B.n83 585
R440 B.n213 B.n212 585
R441 B.n211 B.n84 585
R442 B.n210 B.n209 585
R443 B.n208 B.n85 585
R444 B.n207 B.n206 585
R445 B.n204 B.n86 585
R446 B.n203 B.n202 585
R447 B.n201 B.n89 585
R448 B.n200 B.n199 585
R449 B.n198 B.n90 585
R450 B.n197 B.n196 585
R451 B.n195 B.n91 585
R452 B.n194 B.n193 585
R453 B.n192 B.n92 585
R454 B.n190 B.n189 585
R455 B.n188 B.n95 585
R456 B.n187 B.n186 585
R457 B.n185 B.n96 585
R458 B.n184 B.n183 585
R459 B.n182 B.n97 585
R460 B.n181 B.n180 585
R461 B.n179 B.n98 585
R462 B.n178 B.n177 585
R463 B.n176 B.n99 585
R464 B.n175 B.n174 585
R465 B.n173 B.n100 585
R466 B.n172 B.n171 585
R467 B.n170 B.n101 585
R468 B.n169 B.n168 585
R469 B.n167 B.n102 585
R470 B.n166 B.n165 585
R471 B.n164 B.n103 585
R472 B.n163 B.n162 585
R473 B.n161 B.n104 585
R474 B.n160 B.n159 585
R475 B.n158 B.n105 585
R476 B.n157 B.n156 585
R477 B.n155 B.n106 585
R478 B.n154 B.n153 585
R479 B.n152 B.n107 585
R480 B.n246 B.n245 585
R481 B.n247 B.n72 585
R482 B.n249 B.n248 585
R483 B.n250 B.n71 585
R484 B.n252 B.n251 585
R485 B.n253 B.n70 585
R486 B.n255 B.n254 585
R487 B.n256 B.n69 585
R488 B.n258 B.n257 585
R489 B.n259 B.n68 585
R490 B.n261 B.n260 585
R491 B.n262 B.n67 585
R492 B.n264 B.n263 585
R493 B.n265 B.n66 585
R494 B.n267 B.n266 585
R495 B.n268 B.n65 585
R496 B.n270 B.n269 585
R497 B.n271 B.n64 585
R498 B.n273 B.n272 585
R499 B.n274 B.n63 585
R500 B.n276 B.n275 585
R501 B.n277 B.n62 585
R502 B.n279 B.n278 585
R503 B.n280 B.n61 585
R504 B.n282 B.n281 585
R505 B.n283 B.n60 585
R506 B.n285 B.n284 585
R507 B.n286 B.n59 585
R508 B.n288 B.n287 585
R509 B.n289 B.n58 585
R510 B.n291 B.n290 585
R511 B.n292 B.n57 585
R512 B.n294 B.n293 585
R513 B.n295 B.n56 585
R514 B.n297 B.n296 585
R515 B.n298 B.n55 585
R516 B.n300 B.n299 585
R517 B.n301 B.n54 585
R518 B.n303 B.n302 585
R519 B.n304 B.n53 585
R520 B.n306 B.n305 585
R521 B.n307 B.n52 585
R522 B.n309 B.n308 585
R523 B.n310 B.n51 585
R524 B.n312 B.n311 585
R525 B.n313 B.n50 585
R526 B.n315 B.n314 585
R527 B.n316 B.n49 585
R528 B.n409 B.n408 585
R529 B.n407 B.n14 585
R530 B.n406 B.n405 585
R531 B.n404 B.n15 585
R532 B.n403 B.n402 585
R533 B.n401 B.n16 585
R534 B.n400 B.n399 585
R535 B.n398 B.n17 585
R536 B.n397 B.n396 585
R537 B.n395 B.n18 585
R538 B.n394 B.n393 585
R539 B.n392 B.n19 585
R540 B.n391 B.n390 585
R541 B.n389 B.n20 585
R542 B.n388 B.n387 585
R543 B.n386 B.n21 585
R544 B.n385 B.n384 585
R545 B.n383 B.n22 585
R546 B.n382 B.n381 585
R547 B.n380 B.n23 585
R548 B.n379 B.n378 585
R549 B.n377 B.n24 585
R550 B.n376 B.n375 585
R551 B.n374 B.n25 585
R552 B.n373 B.n372 585
R553 B.n371 B.n26 585
R554 B.n370 B.n369 585
R555 B.n368 B.n27 585
R556 B.n367 B.n366 585
R557 B.n365 B.n31 585
R558 B.n364 B.n363 585
R559 B.n362 B.n32 585
R560 B.n361 B.n360 585
R561 B.n359 B.n33 585
R562 B.n358 B.n357 585
R563 B.n355 B.n34 585
R564 B.n354 B.n353 585
R565 B.n352 B.n37 585
R566 B.n351 B.n350 585
R567 B.n349 B.n38 585
R568 B.n348 B.n347 585
R569 B.n346 B.n39 585
R570 B.n345 B.n344 585
R571 B.n343 B.n40 585
R572 B.n342 B.n341 585
R573 B.n340 B.n41 585
R574 B.n339 B.n338 585
R575 B.n337 B.n42 585
R576 B.n336 B.n335 585
R577 B.n334 B.n43 585
R578 B.n333 B.n332 585
R579 B.n331 B.n44 585
R580 B.n330 B.n329 585
R581 B.n328 B.n45 585
R582 B.n327 B.n326 585
R583 B.n325 B.n46 585
R584 B.n324 B.n323 585
R585 B.n322 B.n47 585
R586 B.n321 B.n320 585
R587 B.n319 B.n48 585
R588 B.n318 B.n317 585
R589 B.n410 B.n13 585
R590 B.n412 B.n411 585
R591 B.n413 B.n12 585
R592 B.n415 B.n414 585
R593 B.n416 B.n11 585
R594 B.n418 B.n417 585
R595 B.n419 B.n10 585
R596 B.n421 B.n420 585
R597 B.n422 B.n9 585
R598 B.n424 B.n423 585
R599 B.n425 B.n8 585
R600 B.n427 B.n426 585
R601 B.n428 B.n7 585
R602 B.n430 B.n429 585
R603 B.n431 B.n6 585
R604 B.n433 B.n432 585
R605 B.n434 B.n5 585
R606 B.n436 B.n435 585
R607 B.n437 B.n4 585
R608 B.n439 B.n438 585
R609 B.n440 B.n3 585
R610 B.n442 B.n441 585
R611 B.n443 B.n0 585
R612 B.n2 B.n1 585
R613 B.n119 B.n118 585
R614 B.n121 B.n120 585
R615 B.n122 B.n117 585
R616 B.n124 B.n123 585
R617 B.n125 B.n116 585
R618 B.n127 B.n126 585
R619 B.n128 B.n115 585
R620 B.n130 B.n129 585
R621 B.n131 B.n114 585
R622 B.n133 B.n132 585
R623 B.n134 B.n113 585
R624 B.n136 B.n135 585
R625 B.n137 B.n112 585
R626 B.n139 B.n138 585
R627 B.n140 B.n111 585
R628 B.n142 B.n141 585
R629 B.n143 B.n110 585
R630 B.n145 B.n144 585
R631 B.n146 B.n109 585
R632 B.n148 B.n147 585
R633 B.n149 B.n108 585
R634 B.n151 B.n150 585
R635 B.n152 B.n151 463.671
R636 B.n245 B.n244 463.671
R637 B.n317 B.n316 463.671
R638 B.n408 B.n13 463.671
R639 B.n87 B.t4 327.896
R640 B.n35 B.t8 327.896
R641 B.n93 B.t1 327.896
R642 B.n28 B.t11 327.896
R643 B.n88 B.t5 277.277
R644 B.n36 B.t7 277.277
R645 B.n94 B.t2 277.277
R646 B.n29 B.t10 277.277
R647 B.n93 B.t0 276.531
R648 B.n87 B.t3 276.531
R649 B.n35 B.t6 276.531
R650 B.n28 B.t9 276.531
R651 B.n445 B.n444 256.663
R652 B.n444 B.n443 235.042
R653 B.n444 B.n2 235.042
R654 B.n153 B.n152 163.367
R655 B.n153 B.n106 163.367
R656 B.n157 B.n106 163.367
R657 B.n158 B.n157 163.367
R658 B.n159 B.n158 163.367
R659 B.n159 B.n104 163.367
R660 B.n163 B.n104 163.367
R661 B.n164 B.n163 163.367
R662 B.n165 B.n164 163.367
R663 B.n165 B.n102 163.367
R664 B.n169 B.n102 163.367
R665 B.n170 B.n169 163.367
R666 B.n171 B.n170 163.367
R667 B.n171 B.n100 163.367
R668 B.n175 B.n100 163.367
R669 B.n176 B.n175 163.367
R670 B.n177 B.n176 163.367
R671 B.n177 B.n98 163.367
R672 B.n181 B.n98 163.367
R673 B.n182 B.n181 163.367
R674 B.n183 B.n182 163.367
R675 B.n183 B.n96 163.367
R676 B.n187 B.n96 163.367
R677 B.n188 B.n187 163.367
R678 B.n189 B.n188 163.367
R679 B.n189 B.n92 163.367
R680 B.n194 B.n92 163.367
R681 B.n195 B.n194 163.367
R682 B.n196 B.n195 163.367
R683 B.n196 B.n90 163.367
R684 B.n200 B.n90 163.367
R685 B.n201 B.n200 163.367
R686 B.n202 B.n201 163.367
R687 B.n202 B.n86 163.367
R688 B.n207 B.n86 163.367
R689 B.n208 B.n207 163.367
R690 B.n209 B.n208 163.367
R691 B.n209 B.n84 163.367
R692 B.n213 B.n84 163.367
R693 B.n214 B.n213 163.367
R694 B.n215 B.n214 163.367
R695 B.n215 B.n82 163.367
R696 B.n219 B.n82 163.367
R697 B.n220 B.n219 163.367
R698 B.n221 B.n220 163.367
R699 B.n221 B.n80 163.367
R700 B.n225 B.n80 163.367
R701 B.n226 B.n225 163.367
R702 B.n227 B.n226 163.367
R703 B.n227 B.n78 163.367
R704 B.n231 B.n78 163.367
R705 B.n232 B.n231 163.367
R706 B.n233 B.n232 163.367
R707 B.n233 B.n76 163.367
R708 B.n237 B.n76 163.367
R709 B.n238 B.n237 163.367
R710 B.n239 B.n238 163.367
R711 B.n239 B.n74 163.367
R712 B.n243 B.n74 163.367
R713 B.n244 B.n243 163.367
R714 B.n316 B.n315 163.367
R715 B.n315 B.n50 163.367
R716 B.n311 B.n50 163.367
R717 B.n311 B.n310 163.367
R718 B.n310 B.n309 163.367
R719 B.n309 B.n52 163.367
R720 B.n305 B.n52 163.367
R721 B.n305 B.n304 163.367
R722 B.n304 B.n303 163.367
R723 B.n303 B.n54 163.367
R724 B.n299 B.n54 163.367
R725 B.n299 B.n298 163.367
R726 B.n298 B.n297 163.367
R727 B.n297 B.n56 163.367
R728 B.n293 B.n56 163.367
R729 B.n293 B.n292 163.367
R730 B.n292 B.n291 163.367
R731 B.n291 B.n58 163.367
R732 B.n287 B.n58 163.367
R733 B.n287 B.n286 163.367
R734 B.n286 B.n285 163.367
R735 B.n285 B.n60 163.367
R736 B.n281 B.n60 163.367
R737 B.n281 B.n280 163.367
R738 B.n280 B.n279 163.367
R739 B.n279 B.n62 163.367
R740 B.n275 B.n62 163.367
R741 B.n275 B.n274 163.367
R742 B.n274 B.n273 163.367
R743 B.n273 B.n64 163.367
R744 B.n269 B.n64 163.367
R745 B.n269 B.n268 163.367
R746 B.n268 B.n267 163.367
R747 B.n267 B.n66 163.367
R748 B.n263 B.n66 163.367
R749 B.n263 B.n262 163.367
R750 B.n262 B.n261 163.367
R751 B.n261 B.n68 163.367
R752 B.n257 B.n68 163.367
R753 B.n257 B.n256 163.367
R754 B.n256 B.n255 163.367
R755 B.n255 B.n70 163.367
R756 B.n251 B.n70 163.367
R757 B.n251 B.n250 163.367
R758 B.n250 B.n249 163.367
R759 B.n249 B.n72 163.367
R760 B.n245 B.n72 163.367
R761 B.n408 B.n407 163.367
R762 B.n407 B.n406 163.367
R763 B.n406 B.n15 163.367
R764 B.n402 B.n15 163.367
R765 B.n402 B.n401 163.367
R766 B.n401 B.n400 163.367
R767 B.n400 B.n17 163.367
R768 B.n396 B.n17 163.367
R769 B.n396 B.n395 163.367
R770 B.n395 B.n394 163.367
R771 B.n394 B.n19 163.367
R772 B.n390 B.n19 163.367
R773 B.n390 B.n389 163.367
R774 B.n389 B.n388 163.367
R775 B.n388 B.n21 163.367
R776 B.n384 B.n21 163.367
R777 B.n384 B.n383 163.367
R778 B.n383 B.n382 163.367
R779 B.n382 B.n23 163.367
R780 B.n378 B.n23 163.367
R781 B.n378 B.n377 163.367
R782 B.n377 B.n376 163.367
R783 B.n376 B.n25 163.367
R784 B.n372 B.n25 163.367
R785 B.n372 B.n371 163.367
R786 B.n371 B.n370 163.367
R787 B.n370 B.n27 163.367
R788 B.n366 B.n27 163.367
R789 B.n366 B.n365 163.367
R790 B.n365 B.n364 163.367
R791 B.n364 B.n32 163.367
R792 B.n360 B.n32 163.367
R793 B.n360 B.n359 163.367
R794 B.n359 B.n358 163.367
R795 B.n358 B.n34 163.367
R796 B.n353 B.n34 163.367
R797 B.n353 B.n352 163.367
R798 B.n352 B.n351 163.367
R799 B.n351 B.n38 163.367
R800 B.n347 B.n38 163.367
R801 B.n347 B.n346 163.367
R802 B.n346 B.n345 163.367
R803 B.n345 B.n40 163.367
R804 B.n341 B.n40 163.367
R805 B.n341 B.n340 163.367
R806 B.n340 B.n339 163.367
R807 B.n339 B.n42 163.367
R808 B.n335 B.n42 163.367
R809 B.n335 B.n334 163.367
R810 B.n334 B.n333 163.367
R811 B.n333 B.n44 163.367
R812 B.n329 B.n44 163.367
R813 B.n329 B.n328 163.367
R814 B.n328 B.n327 163.367
R815 B.n327 B.n46 163.367
R816 B.n323 B.n46 163.367
R817 B.n323 B.n322 163.367
R818 B.n322 B.n321 163.367
R819 B.n321 B.n48 163.367
R820 B.n317 B.n48 163.367
R821 B.n412 B.n13 163.367
R822 B.n413 B.n412 163.367
R823 B.n414 B.n413 163.367
R824 B.n414 B.n11 163.367
R825 B.n418 B.n11 163.367
R826 B.n419 B.n418 163.367
R827 B.n420 B.n419 163.367
R828 B.n420 B.n9 163.367
R829 B.n424 B.n9 163.367
R830 B.n425 B.n424 163.367
R831 B.n426 B.n425 163.367
R832 B.n426 B.n7 163.367
R833 B.n430 B.n7 163.367
R834 B.n431 B.n430 163.367
R835 B.n432 B.n431 163.367
R836 B.n432 B.n5 163.367
R837 B.n436 B.n5 163.367
R838 B.n437 B.n436 163.367
R839 B.n438 B.n437 163.367
R840 B.n438 B.n3 163.367
R841 B.n442 B.n3 163.367
R842 B.n443 B.n442 163.367
R843 B.n118 B.n2 163.367
R844 B.n121 B.n118 163.367
R845 B.n122 B.n121 163.367
R846 B.n123 B.n122 163.367
R847 B.n123 B.n116 163.367
R848 B.n127 B.n116 163.367
R849 B.n128 B.n127 163.367
R850 B.n129 B.n128 163.367
R851 B.n129 B.n114 163.367
R852 B.n133 B.n114 163.367
R853 B.n134 B.n133 163.367
R854 B.n135 B.n134 163.367
R855 B.n135 B.n112 163.367
R856 B.n139 B.n112 163.367
R857 B.n140 B.n139 163.367
R858 B.n141 B.n140 163.367
R859 B.n141 B.n110 163.367
R860 B.n145 B.n110 163.367
R861 B.n146 B.n145 163.367
R862 B.n147 B.n146 163.367
R863 B.n147 B.n108 163.367
R864 B.n151 B.n108 163.367
R865 B.n191 B.n94 59.5399
R866 B.n205 B.n88 59.5399
R867 B.n356 B.n36 59.5399
R868 B.n30 B.n29 59.5399
R869 B.n94 B.n93 50.6187
R870 B.n88 B.n87 50.6187
R871 B.n36 B.n35 50.6187
R872 B.n29 B.n28 50.6187
R873 B.n410 B.n409 30.1273
R874 B.n318 B.n49 30.1273
R875 B.n246 B.n73 30.1273
R876 B.n150 B.n107 30.1273
R877 B B.n445 18.0485
R878 B.n411 B.n410 10.6151
R879 B.n411 B.n12 10.6151
R880 B.n415 B.n12 10.6151
R881 B.n416 B.n415 10.6151
R882 B.n417 B.n416 10.6151
R883 B.n417 B.n10 10.6151
R884 B.n421 B.n10 10.6151
R885 B.n422 B.n421 10.6151
R886 B.n423 B.n422 10.6151
R887 B.n423 B.n8 10.6151
R888 B.n427 B.n8 10.6151
R889 B.n428 B.n427 10.6151
R890 B.n429 B.n428 10.6151
R891 B.n429 B.n6 10.6151
R892 B.n433 B.n6 10.6151
R893 B.n434 B.n433 10.6151
R894 B.n435 B.n434 10.6151
R895 B.n435 B.n4 10.6151
R896 B.n439 B.n4 10.6151
R897 B.n440 B.n439 10.6151
R898 B.n441 B.n440 10.6151
R899 B.n441 B.n0 10.6151
R900 B.n409 B.n14 10.6151
R901 B.n405 B.n14 10.6151
R902 B.n405 B.n404 10.6151
R903 B.n404 B.n403 10.6151
R904 B.n403 B.n16 10.6151
R905 B.n399 B.n16 10.6151
R906 B.n399 B.n398 10.6151
R907 B.n398 B.n397 10.6151
R908 B.n397 B.n18 10.6151
R909 B.n393 B.n18 10.6151
R910 B.n393 B.n392 10.6151
R911 B.n392 B.n391 10.6151
R912 B.n391 B.n20 10.6151
R913 B.n387 B.n20 10.6151
R914 B.n387 B.n386 10.6151
R915 B.n386 B.n385 10.6151
R916 B.n385 B.n22 10.6151
R917 B.n381 B.n22 10.6151
R918 B.n381 B.n380 10.6151
R919 B.n380 B.n379 10.6151
R920 B.n379 B.n24 10.6151
R921 B.n375 B.n24 10.6151
R922 B.n375 B.n374 10.6151
R923 B.n374 B.n373 10.6151
R924 B.n373 B.n26 10.6151
R925 B.n369 B.n368 10.6151
R926 B.n368 B.n367 10.6151
R927 B.n367 B.n31 10.6151
R928 B.n363 B.n31 10.6151
R929 B.n363 B.n362 10.6151
R930 B.n362 B.n361 10.6151
R931 B.n361 B.n33 10.6151
R932 B.n357 B.n33 10.6151
R933 B.n355 B.n354 10.6151
R934 B.n354 B.n37 10.6151
R935 B.n350 B.n37 10.6151
R936 B.n350 B.n349 10.6151
R937 B.n349 B.n348 10.6151
R938 B.n348 B.n39 10.6151
R939 B.n344 B.n39 10.6151
R940 B.n344 B.n343 10.6151
R941 B.n343 B.n342 10.6151
R942 B.n342 B.n41 10.6151
R943 B.n338 B.n41 10.6151
R944 B.n338 B.n337 10.6151
R945 B.n337 B.n336 10.6151
R946 B.n336 B.n43 10.6151
R947 B.n332 B.n43 10.6151
R948 B.n332 B.n331 10.6151
R949 B.n331 B.n330 10.6151
R950 B.n330 B.n45 10.6151
R951 B.n326 B.n45 10.6151
R952 B.n326 B.n325 10.6151
R953 B.n325 B.n324 10.6151
R954 B.n324 B.n47 10.6151
R955 B.n320 B.n47 10.6151
R956 B.n320 B.n319 10.6151
R957 B.n319 B.n318 10.6151
R958 B.n314 B.n49 10.6151
R959 B.n314 B.n313 10.6151
R960 B.n313 B.n312 10.6151
R961 B.n312 B.n51 10.6151
R962 B.n308 B.n51 10.6151
R963 B.n308 B.n307 10.6151
R964 B.n307 B.n306 10.6151
R965 B.n306 B.n53 10.6151
R966 B.n302 B.n53 10.6151
R967 B.n302 B.n301 10.6151
R968 B.n301 B.n300 10.6151
R969 B.n300 B.n55 10.6151
R970 B.n296 B.n55 10.6151
R971 B.n296 B.n295 10.6151
R972 B.n295 B.n294 10.6151
R973 B.n294 B.n57 10.6151
R974 B.n290 B.n57 10.6151
R975 B.n290 B.n289 10.6151
R976 B.n289 B.n288 10.6151
R977 B.n288 B.n59 10.6151
R978 B.n284 B.n59 10.6151
R979 B.n284 B.n283 10.6151
R980 B.n283 B.n282 10.6151
R981 B.n282 B.n61 10.6151
R982 B.n278 B.n61 10.6151
R983 B.n278 B.n277 10.6151
R984 B.n277 B.n276 10.6151
R985 B.n276 B.n63 10.6151
R986 B.n272 B.n63 10.6151
R987 B.n272 B.n271 10.6151
R988 B.n271 B.n270 10.6151
R989 B.n270 B.n65 10.6151
R990 B.n266 B.n65 10.6151
R991 B.n266 B.n265 10.6151
R992 B.n265 B.n264 10.6151
R993 B.n264 B.n67 10.6151
R994 B.n260 B.n67 10.6151
R995 B.n260 B.n259 10.6151
R996 B.n259 B.n258 10.6151
R997 B.n258 B.n69 10.6151
R998 B.n254 B.n69 10.6151
R999 B.n254 B.n253 10.6151
R1000 B.n253 B.n252 10.6151
R1001 B.n252 B.n71 10.6151
R1002 B.n248 B.n71 10.6151
R1003 B.n248 B.n247 10.6151
R1004 B.n247 B.n246 10.6151
R1005 B.n119 B.n1 10.6151
R1006 B.n120 B.n119 10.6151
R1007 B.n120 B.n117 10.6151
R1008 B.n124 B.n117 10.6151
R1009 B.n125 B.n124 10.6151
R1010 B.n126 B.n125 10.6151
R1011 B.n126 B.n115 10.6151
R1012 B.n130 B.n115 10.6151
R1013 B.n131 B.n130 10.6151
R1014 B.n132 B.n131 10.6151
R1015 B.n132 B.n113 10.6151
R1016 B.n136 B.n113 10.6151
R1017 B.n137 B.n136 10.6151
R1018 B.n138 B.n137 10.6151
R1019 B.n138 B.n111 10.6151
R1020 B.n142 B.n111 10.6151
R1021 B.n143 B.n142 10.6151
R1022 B.n144 B.n143 10.6151
R1023 B.n144 B.n109 10.6151
R1024 B.n148 B.n109 10.6151
R1025 B.n149 B.n148 10.6151
R1026 B.n150 B.n149 10.6151
R1027 B.n154 B.n107 10.6151
R1028 B.n155 B.n154 10.6151
R1029 B.n156 B.n155 10.6151
R1030 B.n156 B.n105 10.6151
R1031 B.n160 B.n105 10.6151
R1032 B.n161 B.n160 10.6151
R1033 B.n162 B.n161 10.6151
R1034 B.n162 B.n103 10.6151
R1035 B.n166 B.n103 10.6151
R1036 B.n167 B.n166 10.6151
R1037 B.n168 B.n167 10.6151
R1038 B.n168 B.n101 10.6151
R1039 B.n172 B.n101 10.6151
R1040 B.n173 B.n172 10.6151
R1041 B.n174 B.n173 10.6151
R1042 B.n174 B.n99 10.6151
R1043 B.n178 B.n99 10.6151
R1044 B.n179 B.n178 10.6151
R1045 B.n180 B.n179 10.6151
R1046 B.n180 B.n97 10.6151
R1047 B.n184 B.n97 10.6151
R1048 B.n185 B.n184 10.6151
R1049 B.n186 B.n185 10.6151
R1050 B.n186 B.n95 10.6151
R1051 B.n190 B.n95 10.6151
R1052 B.n193 B.n192 10.6151
R1053 B.n193 B.n91 10.6151
R1054 B.n197 B.n91 10.6151
R1055 B.n198 B.n197 10.6151
R1056 B.n199 B.n198 10.6151
R1057 B.n199 B.n89 10.6151
R1058 B.n203 B.n89 10.6151
R1059 B.n204 B.n203 10.6151
R1060 B.n206 B.n85 10.6151
R1061 B.n210 B.n85 10.6151
R1062 B.n211 B.n210 10.6151
R1063 B.n212 B.n211 10.6151
R1064 B.n212 B.n83 10.6151
R1065 B.n216 B.n83 10.6151
R1066 B.n217 B.n216 10.6151
R1067 B.n218 B.n217 10.6151
R1068 B.n218 B.n81 10.6151
R1069 B.n222 B.n81 10.6151
R1070 B.n223 B.n222 10.6151
R1071 B.n224 B.n223 10.6151
R1072 B.n224 B.n79 10.6151
R1073 B.n228 B.n79 10.6151
R1074 B.n229 B.n228 10.6151
R1075 B.n230 B.n229 10.6151
R1076 B.n230 B.n77 10.6151
R1077 B.n234 B.n77 10.6151
R1078 B.n235 B.n234 10.6151
R1079 B.n236 B.n235 10.6151
R1080 B.n236 B.n75 10.6151
R1081 B.n240 B.n75 10.6151
R1082 B.n241 B.n240 10.6151
R1083 B.n242 B.n241 10.6151
R1084 B.n242 B.n73 10.6151
R1085 B.n445 B.n0 8.11757
R1086 B.n445 B.n1 8.11757
R1087 B.n369 B.n30 6.5566
R1088 B.n357 B.n356 6.5566
R1089 B.n192 B.n191 6.5566
R1090 B.n205 B.n204 6.5566
R1091 B.n30 B.n26 4.05904
R1092 B.n356 B.n355 4.05904
R1093 B.n191 B.n190 4.05904
R1094 B.n206 B.n205 4.05904
C0 VDD2 VP 0.319162f
C1 VP VN 4.29417f
C2 w_n2014_n2274# VP 2.91405f
C3 VDD1 VDD2 0.635655f
C4 VDD1 VN 0.147975f
C5 w_n2014_n2274# VDD1 1.36274f
C6 VTAIL VP 1.56783f
C7 VDD2 B 1.26137f
C8 VDD1 VTAIL 3.55052f
C9 VN B 0.929499f
C10 w_n2014_n2274# B 6.93594f
C11 VTAIL B 2.32319f
C12 VDD1 VP 1.76642f
C13 VP B 1.34885f
C14 VDD2 VN 1.59689f
C15 VDD1 B 1.23413f
C16 w_n2014_n2274# VDD2 1.38477f
C17 w_n2014_n2274# VN 2.6582f
C18 VTAIL VDD2 3.60005f
C19 VTAIL VN 1.5536f
C20 w_n2014_n2274# VTAIL 1.98164f
C21 VDD2 VSUBS 0.65168f
C22 VDD1 VSUBS 2.305734f
C23 VTAIL VSUBS 0.539338f
C24 VN VSUBS 5.25466f
C25 VP VSUBS 1.285995f
C26 B VSUBS 3.209399f
C27 w_n2014_n2274# VSUBS 57.060604f
C28 B.n0 VSUBS 0.006748f
C29 B.n1 VSUBS 0.006748f
C30 B.n2 VSUBS 0.009979f
C31 B.n3 VSUBS 0.007647f
C32 B.n4 VSUBS 0.007647f
C33 B.n5 VSUBS 0.007647f
C34 B.n6 VSUBS 0.007647f
C35 B.n7 VSUBS 0.007647f
C36 B.n8 VSUBS 0.007647f
C37 B.n9 VSUBS 0.007647f
C38 B.n10 VSUBS 0.007647f
C39 B.n11 VSUBS 0.007647f
C40 B.n12 VSUBS 0.007647f
C41 B.n13 VSUBS 0.016396f
C42 B.n14 VSUBS 0.007647f
C43 B.n15 VSUBS 0.007647f
C44 B.n16 VSUBS 0.007647f
C45 B.n17 VSUBS 0.007647f
C46 B.n18 VSUBS 0.007647f
C47 B.n19 VSUBS 0.007647f
C48 B.n20 VSUBS 0.007647f
C49 B.n21 VSUBS 0.007647f
C50 B.n22 VSUBS 0.007647f
C51 B.n23 VSUBS 0.007647f
C52 B.n24 VSUBS 0.007647f
C53 B.n25 VSUBS 0.007647f
C54 B.n26 VSUBS 0.005286f
C55 B.n27 VSUBS 0.007647f
C56 B.t10 VSUBS 0.107743f
C57 B.t11 VSUBS 0.133911f
C58 B.t9 VSUBS 0.760854f
C59 B.n28 VSUBS 0.228853f
C60 B.n29 VSUBS 0.180416f
C61 B.n30 VSUBS 0.017718f
C62 B.n31 VSUBS 0.007647f
C63 B.n32 VSUBS 0.007647f
C64 B.n33 VSUBS 0.007647f
C65 B.n34 VSUBS 0.007647f
C66 B.t7 VSUBS 0.107745f
C67 B.t8 VSUBS 0.133913f
C68 B.t6 VSUBS 0.760854f
C69 B.n35 VSUBS 0.228851f
C70 B.n36 VSUBS 0.180414f
C71 B.n37 VSUBS 0.007647f
C72 B.n38 VSUBS 0.007647f
C73 B.n39 VSUBS 0.007647f
C74 B.n40 VSUBS 0.007647f
C75 B.n41 VSUBS 0.007647f
C76 B.n42 VSUBS 0.007647f
C77 B.n43 VSUBS 0.007647f
C78 B.n44 VSUBS 0.007647f
C79 B.n45 VSUBS 0.007647f
C80 B.n46 VSUBS 0.007647f
C81 B.n47 VSUBS 0.007647f
C82 B.n48 VSUBS 0.007647f
C83 B.n49 VSUBS 0.016396f
C84 B.n50 VSUBS 0.007647f
C85 B.n51 VSUBS 0.007647f
C86 B.n52 VSUBS 0.007647f
C87 B.n53 VSUBS 0.007647f
C88 B.n54 VSUBS 0.007647f
C89 B.n55 VSUBS 0.007647f
C90 B.n56 VSUBS 0.007647f
C91 B.n57 VSUBS 0.007647f
C92 B.n58 VSUBS 0.007647f
C93 B.n59 VSUBS 0.007647f
C94 B.n60 VSUBS 0.007647f
C95 B.n61 VSUBS 0.007647f
C96 B.n62 VSUBS 0.007647f
C97 B.n63 VSUBS 0.007647f
C98 B.n64 VSUBS 0.007647f
C99 B.n65 VSUBS 0.007647f
C100 B.n66 VSUBS 0.007647f
C101 B.n67 VSUBS 0.007647f
C102 B.n68 VSUBS 0.007647f
C103 B.n69 VSUBS 0.007647f
C104 B.n70 VSUBS 0.007647f
C105 B.n71 VSUBS 0.007647f
C106 B.n72 VSUBS 0.007647f
C107 B.n73 VSUBS 0.016587f
C108 B.n74 VSUBS 0.007647f
C109 B.n75 VSUBS 0.007647f
C110 B.n76 VSUBS 0.007647f
C111 B.n77 VSUBS 0.007647f
C112 B.n78 VSUBS 0.007647f
C113 B.n79 VSUBS 0.007647f
C114 B.n80 VSUBS 0.007647f
C115 B.n81 VSUBS 0.007647f
C116 B.n82 VSUBS 0.007647f
C117 B.n83 VSUBS 0.007647f
C118 B.n84 VSUBS 0.007647f
C119 B.n85 VSUBS 0.007647f
C120 B.n86 VSUBS 0.007647f
C121 B.t5 VSUBS 0.107745f
C122 B.t4 VSUBS 0.133913f
C123 B.t3 VSUBS 0.760854f
C124 B.n87 VSUBS 0.228851f
C125 B.n88 VSUBS 0.180414f
C126 B.n89 VSUBS 0.007647f
C127 B.n90 VSUBS 0.007647f
C128 B.n91 VSUBS 0.007647f
C129 B.n92 VSUBS 0.007647f
C130 B.t2 VSUBS 0.107743f
C131 B.t1 VSUBS 0.133911f
C132 B.t0 VSUBS 0.760854f
C133 B.n93 VSUBS 0.228853f
C134 B.n94 VSUBS 0.180416f
C135 B.n95 VSUBS 0.007647f
C136 B.n96 VSUBS 0.007647f
C137 B.n97 VSUBS 0.007647f
C138 B.n98 VSUBS 0.007647f
C139 B.n99 VSUBS 0.007647f
C140 B.n100 VSUBS 0.007647f
C141 B.n101 VSUBS 0.007647f
C142 B.n102 VSUBS 0.007647f
C143 B.n103 VSUBS 0.007647f
C144 B.n104 VSUBS 0.007647f
C145 B.n105 VSUBS 0.007647f
C146 B.n106 VSUBS 0.007647f
C147 B.n107 VSUBS 0.017567f
C148 B.n108 VSUBS 0.007647f
C149 B.n109 VSUBS 0.007647f
C150 B.n110 VSUBS 0.007647f
C151 B.n111 VSUBS 0.007647f
C152 B.n112 VSUBS 0.007647f
C153 B.n113 VSUBS 0.007647f
C154 B.n114 VSUBS 0.007647f
C155 B.n115 VSUBS 0.007647f
C156 B.n116 VSUBS 0.007647f
C157 B.n117 VSUBS 0.007647f
C158 B.n118 VSUBS 0.007647f
C159 B.n119 VSUBS 0.007647f
C160 B.n120 VSUBS 0.007647f
C161 B.n121 VSUBS 0.007647f
C162 B.n122 VSUBS 0.007647f
C163 B.n123 VSUBS 0.007647f
C164 B.n124 VSUBS 0.007647f
C165 B.n125 VSUBS 0.007647f
C166 B.n126 VSUBS 0.007647f
C167 B.n127 VSUBS 0.007647f
C168 B.n128 VSUBS 0.007647f
C169 B.n129 VSUBS 0.007647f
C170 B.n130 VSUBS 0.007647f
C171 B.n131 VSUBS 0.007647f
C172 B.n132 VSUBS 0.007647f
C173 B.n133 VSUBS 0.007647f
C174 B.n134 VSUBS 0.007647f
C175 B.n135 VSUBS 0.007647f
C176 B.n136 VSUBS 0.007647f
C177 B.n137 VSUBS 0.007647f
C178 B.n138 VSUBS 0.007647f
C179 B.n139 VSUBS 0.007647f
C180 B.n140 VSUBS 0.007647f
C181 B.n141 VSUBS 0.007647f
C182 B.n142 VSUBS 0.007647f
C183 B.n143 VSUBS 0.007647f
C184 B.n144 VSUBS 0.007647f
C185 B.n145 VSUBS 0.007647f
C186 B.n146 VSUBS 0.007647f
C187 B.n147 VSUBS 0.007647f
C188 B.n148 VSUBS 0.007647f
C189 B.n149 VSUBS 0.007647f
C190 B.n150 VSUBS 0.016396f
C191 B.n151 VSUBS 0.016396f
C192 B.n152 VSUBS 0.017567f
C193 B.n153 VSUBS 0.007647f
C194 B.n154 VSUBS 0.007647f
C195 B.n155 VSUBS 0.007647f
C196 B.n156 VSUBS 0.007647f
C197 B.n157 VSUBS 0.007647f
C198 B.n158 VSUBS 0.007647f
C199 B.n159 VSUBS 0.007647f
C200 B.n160 VSUBS 0.007647f
C201 B.n161 VSUBS 0.007647f
C202 B.n162 VSUBS 0.007647f
C203 B.n163 VSUBS 0.007647f
C204 B.n164 VSUBS 0.007647f
C205 B.n165 VSUBS 0.007647f
C206 B.n166 VSUBS 0.007647f
C207 B.n167 VSUBS 0.007647f
C208 B.n168 VSUBS 0.007647f
C209 B.n169 VSUBS 0.007647f
C210 B.n170 VSUBS 0.007647f
C211 B.n171 VSUBS 0.007647f
C212 B.n172 VSUBS 0.007647f
C213 B.n173 VSUBS 0.007647f
C214 B.n174 VSUBS 0.007647f
C215 B.n175 VSUBS 0.007647f
C216 B.n176 VSUBS 0.007647f
C217 B.n177 VSUBS 0.007647f
C218 B.n178 VSUBS 0.007647f
C219 B.n179 VSUBS 0.007647f
C220 B.n180 VSUBS 0.007647f
C221 B.n181 VSUBS 0.007647f
C222 B.n182 VSUBS 0.007647f
C223 B.n183 VSUBS 0.007647f
C224 B.n184 VSUBS 0.007647f
C225 B.n185 VSUBS 0.007647f
C226 B.n186 VSUBS 0.007647f
C227 B.n187 VSUBS 0.007647f
C228 B.n188 VSUBS 0.007647f
C229 B.n189 VSUBS 0.007647f
C230 B.n190 VSUBS 0.005286f
C231 B.n191 VSUBS 0.017718f
C232 B.n192 VSUBS 0.006185f
C233 B.n193 VSUBS 0.007647f
C234 B.n194 VSUBS 0.007647f
C235 B.n195 VSUBS 0.007647f
C236 B.n196 VSUBS 0.007647f
C237 B.n197 VSUBS 0.007647f
C238 B.n198 VSUBS 0.007647f
C239 B.n199 VSUBS 0.007647f
C240 B.n200 VSUBS 0.007647f
C241 B.n201 VSUBS 0.007647f
C242 B.n202 VSUBS 0.007647f
C243 B.n203 VSUBS 0.007647f
C244 B.n204 VSUBS 0.006185f
C245 B.n205 VSUBS 0.017718f
C246 B.n206 VSUBS 0.005286f
C247 B.n207 VSUBS 0.007647f
C248 B.n208 VSUBS 0.007647f
C249 B.n209 VSUBS 0.007647f
C250 B.n210 VSUBS 0.007647f
C251 B.n211 VSUBS 0.007647f
C252 B.n212 VSUBS 0.007647f
C253 B.n213 VSUBS 0.007647f
C254 B.n214 VSUBS 0.007647f
C255 B.n215 VSUBS 0.007647f
C256 B.n216 VSUBS 0.007647f
C257 B.n217 VSUBS 0.007647f
C258 B.n218 VSUBS 0.007647f
C259 B.n219 VSUBS 0.007647f
C260 B.n220 VSUBS 0.007647f
C261 B.n221 VSUBS 0.007647f
C262 B.n222 VSUBS 0.007647f
C263 B.n223 VSUBS 0.007647f
C264 B.n224 VSUBS 0.007647f
C265 B.n225 VSUBS 0.007647f
C266 B.n226 VSUBS 0.007647f
C267 B.n227 VSUBS 0.007647f
C268 B.n228 VSUBS 0.007647f
C269 B.n229 VSUBS 0.007647f
C270 B.n230 VSUBS 0.007647f
C271 B.n231 VSUBS 0.007647f
C272 B.n232 VSUBS 0.007647f
C273 B.n233 VSUBS 0.007647f
C274 B.n234 VSUBS 0.007647f
C275 B.n235 VSUBS 0.007647f
C276 B.n236 VSUBS 0.007647f
C277 B.n237 VSUBS 0.007647f
C278 B.n238 VSUBS 0.007647f
C279 B.n239 VSUBS 0.007647f
C280 B.n240 VSUBS 0.007647f
C281 B.n241 VSUBS 0.007647f
C282 B.n242 VSUBS 0.007647f
C283 B.n243 VSUBS 0.007647f
C284 B.n244 VSUBS 0.017567f
C285 B.n245 VSUBS 0.016396f
C286 B.n246 VSUBS 0.017376f
C287 B.n247 VSUBS 0.007647f
C288 B.n248 VSUBS 0.007647f
C289 B.n249 VSUBS 0.007647f
C290 B.n250 VSUBS 0.007647f
C291 B.n251 VSUBS 0.007647f
C292 B.n252 VSUBS 0.007647f
C293 B.n253 VSUBS 0.007647f
C294 B.n254 VSUBS 0.007647f
C295 B.n255 VSUBS 0.007647f
C296 B.n256 VSUBS 0.007647f
C297 B.n257 VSUBS 0.007647f
C298 B.n258 VSUBS 0.007647f
C299 B.n259 VSUBS 0.007647f
C300 B.n260 VSUBS 0.007647f
C301 B.n261 VSUBS 0.007647f
C302 B.n262 VSUBS 0.007647f
C303 B.n263 VSUBS 0.007647f
C304 B.n264 VSUBS 0.007647f
C305 B.n265 VSUBS 0.007647f
C306 B.n266 VSUBS 0.007647f
C307 B.n267 VSUBS 0.007647f
C308 B.n268 VSUBS 0.007647f
C309 B.n269 VSUBS 0.007647f
C310 B.n270 VSUBS 0.007647f
C311 B.n271 VSUBS 0.007647f
C312 B.n272 VSUBS 0.007647f
C313 B.n273 VSUBS 0.007647f
C314 B.n274 VSUBS 0.007647f
C315 B.n275 VSUBS 0.007647f
C316 B.n276 VSUBS 0.007647f
C317 B.n277 VSUBS 0.007647f
C318 B.n278 VSUBS 0.007647f
C319 B.n279 VSUBS 0.007647f
C320 B.n280 VSUBS 0.007647f
C321 B.n281 VSUBS 0.007647f
C322 B.n282 VSUBS 0.007647f
C323 B.n283 VSUBS 0.007647f
C324 B.n284 VSUBS 0.007647f
C325 B.n285 VSUBS 0.007647f
C326 B.n286 VSUBS 0.007647f
C327 B.n287 VSUBS 0.007647f
C328 B.n288 VSUBS 0.007647f
C329 B.n289 VSUBS 0.007647f
C330 B.n290 VSUBS 0.007647f
C331 B.n291 VSUBS 0.007647f
C332 B.n292 VSUBS 0.007647f
C333 B.n293 VSUBS 0.007647f
C334 B.n294 VSUBS 0.007647f
C335 B.n295 VSUBS 0.007647f
C336 B.n296 VSUBS 0.007647f
C337 B.n297 VSUBS 0.007647f
C338 B.n298 VSUBS 0.007647f
C339 B.n299 VSUBS 0.007647f
C340 B.n300 VSUBS 0.007647f
C341 B.n301 VSUBS 0.007647f
C342 B.n302 VSUBS 0.007647f
C343 B.n303 VSUBS 0.007647f
C344 B.n304 VSUBS 0.007647f
C345 B.n305 VSUBS 0.007647f
C346 B.n306 VSUBS 0.007647f
C347 B.n307 VSUBS 0.007647f
C348 B.n308 VSUBS 0.007647f
C349 B.n309 VSUBS 0.007647f
C350 B.n310 VSUBS 0.007647f
C351 B.n311 VSUBS 0.007647f
C352 B.n312 VSUBS 0.007647f
C353 B.n313 VSUBS 0.007647f
C354 B.n314 VSUBS 0.007647f
C355 B.n315 VSUBS 0.007647f
C356 B.n316 VSUBS 0.016396f
C357 B.n317 VSUBS 0.017567f
C358 B.n318 VSUBS 0.017567f
C359 B.n319 VSUBS 0.007647f
C360 B.n320 VSUBS 0.007647f
C361 B.n321 VSUBS 0.007647f
C362 B.n322 VSUBS 0.007647f
C363 B.n323 VSUBS 0.007647f
C364 B.n324 VSUBS 0.007647f
C365 B.n325 VSUBS 0.007647f
C366 B.n326 VSUBS 0.007647f
C367 B.n327 VSUBS 0.007647f
C368 B.n328 VSUBS 0.007647f
C369 B.n329 VSUBS 0.007647f
C370 B.n330 VSUBS 0.007647f
C371 B.n331 VSUBS 0.007647f
C372 B.n332 VSUBS 0.007647f
C373 B.n333 VSUBS 0.007647f
C374 B.n334 VSUBS 0.007647f
C375 B.n335 VSUBS 0.007647f
C376 B.n336 VSUBS 0.007647f
C377 B.n337 VSUBS 0.007647f
C378 B.n338 VSUBS 0.007647f
C379 B.n339 VSUBS 0.007647f
C380 B.n340 VSUBS 0.007647f
C381 B.n341 VSUBS 0.007647f
C382 B.n342 VSUBS 0.007647f
C383 B.n343 VSUBS 0.007647f
C384 B.n344 VSUBS 0.007647f
C385 B.n345 VSUBS 0.007647f
C386 B.n346 VSUBS 0.007647f
C387 B.n347 VSUBS 0.007647f
C388 B.n348 VSUBS 0.007647f
C389 B.n349 VSUBS 0.007647f
C390 B.n350 VSUBS 0.007647f
C391 B.n351 VSUBS 0.007647f
C392 B.n352 VSUBS 0.007647f
C393 B.n353 VSUBS 0.007647f
C394 B.n354 VSUBS 0.007647f
C395 B.n355 VSUBS 0.005286f
C396 B.n356 VSUBS 0.017718f
C397 B.n357 VSUBS 0.006185f
C398 B.n358 VSUBS 0.007647f
C399 B.n359 VSUBS 0.007647f
C400 B.n360 VSUBS 0.007647f
C401 B.n361 VSUBS 0.007647f
C402 B.n362 VSUBS 0.007647f
C403 B.n363 VSUBS 0.007647f
C404 B.n364 VSUBS 0.007647f
C405 B.n365 VSUBS 0.007647f
C406 B.n366 VSUBS 0.007647f
C407 B.n367 VSUBS 0.007647f
C408 B.n368 VSUBS 0.007647f
C409 B.n369 VSUBS 0.006185f
C410 B.n370 VSUBS 0.007647f
C411 B.n371 VSUBS 0.007647f
C412 B.n372 VSUBS 0.007647f
C413 B.n373 VSUBS 0.007647f
C414 B.n374 VSUBS 0.007647f
C415 B.n375 VSUBS 0.007647f
C416 B.n376 VSUBS 0.007647f
C417 B.n377 VSUBS 0.007647f
C418 B.n378 VSUBS 0.007647f
C419 B.n379 VSUBS 0.007647f
C420 B.n380 VSUBS 0.007647f
C421 B.n381 VSUBS 0.007647f
C422 B.n382 VSUBS 0.007647f
C423 B.n383 VSUBS 0.007647f
C424 B.n384 VSUBS 0.007647f
C425 B.n385 VSUBS 0.007647f
C426 B.n386 VSUBS 0.007647f
C427 B.n387 VSUBS 0.007647f
C428 B.n388 VSUBS 0.007647f
C429 B.n389 VSUBS 0.007647f
C430 B.n390 VSUBS 0.007647f
C431 B.n391 VSUBS 0.007647f
C432 B.n392 VSUBS 0.007647f
C433 B.n393 VSUBS 0.007647f
C434 B.n394 VSUBS 0.007647f
C435 B.n395 VSUBS 0.007647f
C436 B.n396 VSUBS 0.007647f
C437 B.n397 VSUBS 0.007647f
C438 B.n398 VSUBS 0.007647f
C439 B.n399 VSUBS 0.007647f
C440 B.n400 VSUBS 0.007647f
C441 B.n401 VSUBS 0.007647f
C442 B.n402 VSUBS 0.007647f
C443 B.n403 VSUBS 0.007647f
C444 B.n404 VSUBS 0.007647f
C445 B.n405 VSUBS 0.007647f
C446 B.n406 VSUBS 0.007647f
C447 B.n407 VSUBS 0.007647f
C448 B.n408 VSUBS 0.017567f
C449 B.n409 VSUBS 0.017567f
C450 B.n410 VSUBS 0.016396f
C451 B.n411 VSUBS 0.007647f
C452 B.n412 VSUBS 0.007647f
C453 B.n413 VSUBS 0.007647f
C454 B.n414 VSUBS 0.007647f
C455 B.n415 VSUBS 0.007647f
C456 B.n416 VSUBS 0.007647f
C457 B.n417 VSUBS 0.007647f
C458 B.n418 VSUBS 0.007647f
C459 B.n419 VSUBS 0.007647f
C460 B.n420 VSUBS 0.007647f
C461 B.n421 VSUBS 0.007647f
C462 B.n422 VSUBS 0.007647f
C463 B.n423 VSUBS 0.007647f
C464 B.n424 VSUBS 0.007647f
C465 B.n425 VSUBS 0.007647f
C466 B.n426 VSUBS 0.007647f
C467 B.n427 VSUBS 0.007647f
C468 B.n428 VSUBS 0.007647f
C469 B.n429 VSUBS 0.007647f
C470 B.n430 VSUBS 0.007647f
C471 B.n431 VSUBS 0.007647f
C472 B.n432 VSUBS 0.007647f
C473 B.n433 VSUBS 0.007647f
C474 B.n434 VSUBS 0.007647f
C475 B.n435 VSUBS 0.007647f
C476 B.n436 VSUBS 0.007647f
C477 B.n437 VSUBS 0.007647f
C478 B.n438 VSUBS 0.007647f
C479 B.n439 VSUBS 0.007647f
C480 B.n440 VSUBS 0.007647f
C481 B.n441 VSUBS 0.007647f
C482 B.n442 VSUBS 0.007647f
C483 B.n443 VSUBS 0.009979f
C484 B.n444 VSUBS 0.010631f
C485 B.n445 VSUBS 0.02114f
C486 VDD1.n0 VSUBS 0.008003f
C487 VDD1.n1 VSUBS 0.018051f
C488 VDD1.n2 VSUBS 0.008086f
C489 VDD1.n3 VSUBS 0.014212f
C490 VDD1.n4 VSUBS 0.007637f
C491 VDD1.n5 VSUBS 0.018051f
C492 VDD1.n6 VSUBS 0.008086f
C493 VDD1.n7 VSUBS 0.014212f
C494 VDD1.n8 VSUBS 0.007637f
C495 VDD1.n9 VSUBS 0.013538f
C496 VDD1.n10 VSUBS 0.013577f
C497 VDD1.t0 VSUBS 0.038812f
C498 VDD1.n11 VSUBS 0.076922f
C499 VDD1.n12 VSUBS 0.357347f
C500 VDD1.n13 VSUBS 0.007637f
C501 VDD1.n14 VSUBS 0.008086f
C502 VDD1.n15 VSUBS 0.018051f
C503 VDD1.n16 VSUBS 0.018051f
C504 VDD1.n17 VSUBS 0.008086f
C505 VDD1.n18 VSUBS 0.007637f
C506 VDD1.n19 VSUBS 0.014212f
C507 VDD1.n20 VSUBS 0.014212f
C508 VDD1.n21 VSUBS 0.007637f
C509 VDD1.n22 VSUBS 0.008086f
C510 VDD1.n23 VSUBS 0.018051f
C511 VDD1.n24 VSUBS 0.018051f
C512 VDD1.n25 VSUBS 0.008086f
C513 VDD1.n26 VSUBS 0.007637f
C514 VDD1.n27 VSUBS 0.014212f
C515 VDD1.n28 VSUBS 0.036152f
C516 VDD1.n29 VSUBS 0.007637f
C517 VDD1.n30 VSUBS 0.008086f
C518 VDD1.n31 VSUBS 0.04042f
C519 VDD1.n32 VSUBS 0.037172f
C520 VDD1.n33 VSUBS 0.008003f
C521 VDD1.n34 VSUBS 0.018051f
C522 VDD1.n35 VSUBS 0.008086f
C523 VDD1.n36 VSUBS 0.014212f
C524 VDD1.n37 VSUBS 0.007637f
C525 VDD1.n38 VSUBS 0.018051f
C526 VDD1.n39 VSUBS 0.008086f
C527 VDD1.n40 VSUBS 0.014212f
C528 VDD1.n41 VSUBS 0.007637f
C529 VDD1.n42 VSUBS 0.013538f
C530 VDD1.n43 VSUBS 0.013577f
C531 VDD1.t1 VSUBS 0.038812f
C532 VDD1.n44 VSUBS 0.076922f
C533 VDD1.n45 VSUBS 0.357347f
C534 VDD1.n46 VSUBS 0.007637f
C535 VDD1.n47 VSUBS 0.008086f
C536 VDD1.n48 VSUBS 0.018051f
C537 VDD1.n49 VSUBS 0.018051f
C538 VDD1.n50 VSUBS 0.008086f
C539 VDD1.n51 VSUBS 0.007637f
C540 VDD1.n52 VSUBS 0.014212f
C541 VDD1.n53 VSUBS 0.014212f
C542 VDD1.n54 VSUBS 0.007637f
C543 VDD1.n55 VSUBS 0.008086f
C544 VDD1.n56 VSUBS 0.018051f
C545 VDD1.n57 VSUBS 0.018051f
C546 VDD1.n58 VSUBS 0.008086f
C547 VDD1.n59 VSUBS 0.007637f
C548 VDD1.n60 VSUBS 0.014212f
C549 VDD1.n61 VSUBS 0.036152f
C550 VDD1.n62 VSUBS 0.007637f
C551 VDD1.n63 VSUBS 0.008086f
C552 VDD1.n64 VSUBS 0.04042f
C553 VDD1.n65 VSUBS 0.322038f
C554 VP.t1 VSUBS 2.17498f
C555 VP.t0 VSUBS 1.70211f
C556 VP.n0 VSUBS 3.24888f
C557 VDD2.n0 VSUBS 0.008122f
C558 VDD2.n1 VSUBS 0.018319f
C559 VDD2.n2 VSUBS 0.008206f
C560 VDD2.n3 VSUBS 0.014423f
C561 VDD2.n4 VSUBS 0.00775f
C562 VDD2.n5 VSUBS 0.018319f
C563 VDD2.n6 VSUBS 0.008206f
C564 VDD2.n7 VSUBS 0.014423f
C565 VDD2.n8 VSUBS 0.00775f
C566 VDD2.n9 VSUBS 0.013739f
C567 VDD2.n10 VSUBS 0.013778f
C568 VDD2.t1 VSUBS 0.039386f
C569 VDD2.n11 VSUBS 0.07806f
C570 VDD2.n12 VSUBS 0.362635f
C571 VDD2.n13 VSUBS 0.00775f
C572 VDD2.n14 VSUBS 0.008206f
C573 VDD2.n15 VSUBS 0.018319f
C574 VDD2.n16 VSUBS 0.018319f
C575 VDD2.n17 VSUBS 0.008206f
C576 VDD2.n18 VSUBS 0.00775f
C577 VDD2.n19 VSUBS 0.014423f
C578 VDD2.n20 VSUBS 0.014423f
C579 VDD2.n21 VSUBS 0.00775f
C580 VDD2.n22 VSUBS 0.008206f
C581 VDD2.n23 VSUBS 0.018319f
C582 VDD2.n24 VSUBS 0.018319f
C583 VDD2.n25 VSUBS 0.008206f
C584 VDD2.n26 VSUBS 0.00775f
C585 VDD2.n27 VSUBS 0.014423f
C586 VDD2.n28 VSUBS 0.036687f
C587 VDD2.n29 VSUBS 0.00775f
C588 VDD2.n30 VSUBS 0.008206f
C589 VDD2.n31 VSUBS 0.041018f
C590 VDD2.n32 VSUBS 0.303562f
C591 VDD2.n33 VSUBS 0.008122f
C592 VDD2.n34 VSUBS 0.018319f
C593 VDD2.n35 VSUBS 0.008206f
C594 VDD2.n36 VSUBS 0.014423f
C595 VDD2.n37 VSUBS 0.00775f
C596 VDD2.n38 VSUBS 0.018319f
C597 VDD2.n39 VSUBS 0.008206f
C598 VDD2.n40 VSUBS 0.014423f
C599 VDD2.n41 VSUBS 0.00775f
C600 VDD2.n42 VSUBS 0.013739f
C601 VDD2.n43 VSUBS 0.013778f
C602 VDD2.t0 VSUBS 0.039386f
C603 VDD2.n44 VSUBS 0.07806f
C604 VDD2.n45 VSUBS 0.362635f
C605 VDD2.n46 VSUBS 0.00775f
C606 VDD2.n47 VSUBS 0.008206f
C607 VDD2.n48 VSUBS 0.018319f
C608 VDD2.n49 VSUBS 0.018319f
C609 VDD2.n50 VSUBS 0.008206f
C610 VDD2.n51 VSUBS 0.00775f
C611 VDD2.n52 VSUBS 0.014423f
C612 VDD2.n53 VSUBS 0.014423f
C613 VDD2.n54 VSUBS 0.00775f
C614 VDD2.n55 VSUBS 0.008206f
C615 VDD2.n56 VSUBS 0.018319f
C616 VDD2.n57 VSUBS 0.018319f
C617 VDD2.n58 VSUBS 0.008206f
C618 VDD2.n59 VSUBS 0.00775f
C619 VDD2.n60 VSUBS 0.014423f
C620 VDD2.n61 VSUBS 0.036687f
C621 VDD2.n62 VSUBS 0.00775f
C622 VDD2.n63 VSUBS 0.008206f
C623 VDD2.n64 VSUBS 0.041018f
C624 VDD2.n65 VSUBS 0.037032f
C625 VDD2.n66 VSUBS 1.40359f
C626 VTAIL.n0 VSUBS 0.011931f
C627 VTAIL.n1 VSUBS 0.02691f
C628 VTAIL.n2 VSUBS 0.012055f
C629 VTAIL.n3 VSUBS 0.021187f
C630 VTAIL.n4 VSUBS 0.011385f
C631 VTAIL.n5 VSUBS 0.02691f
C632 VTAIL.n6 VSUBS 0.012055f
C633 VTAIL.n7 VSUBS 0.021187f
C634 VTAIL.n8 VSUBS 0.011385f
C635 VTAIL.n9 VSUBS 0.020183f
C636 VTAIL.n10 VSUBS 0.02024f
C637 VTAIL.t1 VSUBS 0.057859f
C638 VTAIL.n11 VSUBS 0.114673f
C639 VTAIL.n12 VSUBS 0.532721f
C640 VTAIL.n13 VSUBS 0.011385f
C641 VTAIL.n14 VSUBS 0.012055f
C642 VTAIL.n15 VSUBS 0.02691f
C643 VTAIL.n16 VSUBS 0.02691f
C644 VTAIL.n17 VSUBS 0.012055f
C645 VTAIL.n18 VSUBS 0.011385f
C646 VTAIL.n19 VSUBS 0.021187f
C647 VTAIL.n20 VSUBS 0.021187f
C648 VTAIL.n21 VSUBS 0.011385f
C649 VTAIL.n22 VSUBS 0.012055f
C650 VTAIL.n23 VSUBS 0.02691f
C651 VTAIL.n24 VSUBS 0.02691f
C652 VTAIL.n25 VSUBS 0.012055f
C653 VTAIL.n26 VSUBS 0.011385f
C654 VTAIL.n27 VSUBS 0.021187f
C655 VTAIL.n28 VSUBS 0.053894f
C656 VTAIL.n29 VSUBS 0.011385f
C657 VTAIL.n30 VSUBS 0.012055f
C658 VTAIL.n31 VSUBS 0.060256f
C659 VTAIL.n32 VSUBS 0.039802f
C660 VTAIL.n33 VSUBS 1.07434f
C661 VTAIL.n34 VSUBS 0.011931f
C662 VTAIL.n35 VSUBS 0.02691f
C663 VTAIL.n36 VSUBS 0.012055f
C664 VTAIL.n37 VSUBS 0.021187f
C665 VTAIL.n38 VSUBS 0.011385f
C666 VTAIL.n39 VSUBS 0.02691f
C667 VTAIL.n40 VSUBS 0.012055f
C668 VTAIL.n41 VSUBS 0.021187f
C669 VTAIL.n42 VSUBS 0.011385f
C670 VTAIL.n43 VSUBS 0.020183f
C671 VTAIL.n44 VSUBS 0.02024f
C672 VTAIL.t2 VSUBS 0.057859f
C673 VTAIL.n45 VSUBS 0.114673f
C674 VTAIL.n46 VSUBS 0.532721f
C675 VTAIL.n47 VSUBS 0.011385f
C676 VTAIL.n48 VSUBS 0.012055f
C677 VTAIL.n49 VSUBS 0.02691f
C678 VTAIL.n50 VSUBS 0.02691f
C679 VTAIL.n51 VSUBS 0.012055f
C680 VTAIL.n52 VSUBS 0.011385f
C681 VTAIL.n53 VSUBS 0.021187f
C682 VTAIL.n54 VSUBS 0.021187f
C683 VTAIL.n55 VSUBS 0.011385f
C684 VTAIL.n56 VSUBS 0.012055f
C685 VTAIL.n57 VSUBS 0.02691f
C686 VTAIL.n58 VSUBS 0.02691f
C687 VTAIL.n59 VSUBS 0.012055f
C688 VTAIL.n60 VSUBS 0.011385f
C689 VTAIL.n61 VSUBS 0.021187f
C690 VTAIL.n62 VSUBS 0.053894f
C691 VTAIL.n63 VSUBS 0.011385f
C692 VTAIL.n64 VSUBS 0.012055f
C693 VTAIL.n65 VSUBS 0.060256f
C694 VTAIL.n66 VSUBS 0.039802f
C695 VTAIL.n67 VSUBS 1.10877f
C696 VTAIL.n68 VSUBS 0.011931f
C697 VTAIL.n69 VSUBS 0.02691f
C698 VTAIL.n70 VSUBS 0.012055f
C699 VTAIL.n71 VSUBS 0.021187f
C700 VTAIL.n72 VSUBS 0.011385f
C701 VTAIL.n73 VSUBS 0.02691f
C702 VTAIL.n74 VSUBS 0.012055f
C703 VTAIL.n75 VSUBS 0.021187f
C704 VTAIL.n76 VSUBS 0.011385f
C705 VTAIL.n77 VSUBS 0.020183f
C706 VTAIL.n78 VSUBS 0.02024f
C707 VTAIL.t0 VSUBS 0.057859f
C708 VTAIL.n79 VSUBS 0.114673f
C709 VTAIL.n80 VSUBS 0.532721f
C710 VTAIL.n81 VSUBS 0.011385f
C711 VTAIL.n82 VSUBS 0.012055f
C712 VTAIL.n83 VSUBS 0.02691f
C713 VTAIL.n84 VSUBS 0.02691f
C714 VTAIL.n85 VSUBS 0.012055f
C715 VTAIL.n86 VSUBS 0.011385f
C716 VTAIL.n87 VSUBS 0.021187f
C717 VTAIL.n88 VSUBS 0.021187f
C718 VTAIL.n89 VSUBS 0.011385f
C719 VTAIL.n90 VSUBS 0.012055f
C720 VTAIL.n91 VSUBS 0.02691f
C721 VTAIL.n92 VSUBS 0.02691f
C722 VTAIL.n93 VSUBS 0.012055f
C723 VTAIL.n94 VSUBS 0.011385f
C724 VTAIL.n95 VSUBS 0.021187f
C725 VTAIL.n96 VSUBS 0.053894f
C726 VTAIL.n97 VSUBS 0.011385f
C727 VTAIL.n98 VSUBS 0.012055f
C728 VTAIL.n99 VSUBS 0.060256f
C729 VTAIL.n100 VSUBS 0.039802f
C730 VTAIL.n101 VSUBS 0.955157f
C731 VTAIL.n102 VSUBS 0.011931f
C732 VTAIL.n103 VSUBS 0.02691f
C733 VTAIL.n104 VSUBS 0.012055f
C734 VTAIL.n105 VSUBS 0.021187f
C735 VTAIL.n106 VSUBS 0.011385f
C736 VTAIL.n107 VSUBS 0.02691f
C737 VTAIL.n108 VSUBS 0.012055f
C738 VTAIL.n109 VSUBS 0.021187f
C739 VTAIL.n110 VSUBS 0.011385f
C740 VTAIL.n111 VSUBS 0.020183f
C741 VTAIL.n112 VSUBS 0.02024f
C742 VTAIL.t3 VSUBS 0.057859f
C743 VTAIL.n113 VSUBS 0.114673f
C744 VTAIL.n114 VSUBS 0.532721f
C745 VTAIL.n115 VSUBS 0.011385f
C746 VTAIL.n116 VSUBS 0.012055f
C747 VTAIL.n117 VSUBS 0.02691f
C748 VTAIL.n118 VSUBS 0.02691f
C749 VTAIL.n119 VSUBS 0.012055f
C750 VTAIL.n120 VSUBS 0.011385f
C751 VTAIL.n121 VSUBS 0.021187f
C752 VTAIL.n122 VSUBS 0.021187f
C753 VTAIL.n123 VSUBS 0.011385f
C754 VTAIL.n124 VSUBS 0.012055f
C755 VTAIL.n125 VSUBS 0.02691f
C756 VTAIL.n126 VSUBS 0.02691f
C757 VTAIL.n127 VSUBS 0.012055f
C758 VTAIL.n128 VSUBS 0.011385f
C759 VTAIL.n129 VSUBS 0.021187f
C760 VTAIL.n130 VSUBS 0.053894f
C761 VTAIL.n131 VSUBS 0.011385f
C762 VTAIL.n132 VSUBS 0.012055f
C763 VTAIL.n133 VSUBS 0.060256f
C764 VTAIL.n134 VSUBS 0.039802f
C765 VTAIL.n135 VSUBS 0.880707f
C766 VN.t0 VSUBS 1.64506f
C767 VN.t1 VSUBS 2.10416f
.ends

