* NGSPICE file created from diff_pair_sample_1765.ext - technology: sky130A

.subckt diff_pair_sample_1765 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=2.0163 ps=11.12 w=5.17 l=0.34
X1 VDD2.t4 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0.85305 ps=5.5 w=5.17 l=0.34
X2 VTAIL.t7 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=0.85305 ps=5.5 w=5.17 l=0.34
X3 VTAIL.t5 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=0.85305 ps=5.5 w=5.17 l=0.34
X4 VTAIL.t10 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=0.85305 ps=5.5 w=5.17 l=0.34
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0 ps=0 w=5.17 l=0.34
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0 ps=0 w=5.17 l=0.34
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0 ps=0 w=5.17 l=0.34
X8 VDD2.t1 VN.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0.85305 ps=5.5 w=5.17 l=0.34
X9 VTAIL.t0 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=0.85305 ps=5.5 w=5.17 l=0.34
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0 ps=0 w=5.17 l=0.34
X11 VDD2.t0 VN.t5 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=2.0163 ps=11.12 w=5.17 l=0.34
X12 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=2.0163 ps=11.12 w=5.17 l=0.34
X13 VDD1.t2 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0.85305 ps=5.5 w=5.17 l=0.34
X14 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=11.12 as=0.85305 ps=5.5 w=5.17 l=0.34
X15 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85305 pd=5.5 as=2.0163 ps=11.12 w=5.17 l=0.34
R0 VN.n0 VN.t4 503.69
R1 VN.n4 VN.t5 503.69
R2 VN.n2 VN.t0 482.709
R3 VN.n1 VN.t2 482.709
R4 VN.n5 VN.t3 482.709
R5 VN.n6 VN.t1 482.709
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 70.4033
R9 VN.n3 VN.n0 70.4033
R10 VN.n2 VN.n1 48.2005
R11 VN.n6 VN.n5 48.2005
R12 VN VN.n7 35.0138
R13 VN.n5 VN.n4 20.9576
R14 VN.n1 VN.n0 20.9576
R15 VN VN.n3 0.0516364
R16 VTAIL.n114 VTAIL.n92 289.615
R17 VTAIL.n24 VTAIL.n2 289.615
R18 VTAIL.n86 VTAIL.n64 289.615
R19 VTAIL.n56 VTAIL.n34 289.615
R20 VTAIL.n100 VTAIL.n99 185
R21 VTAIL.n105 VTAIL.n104 185
R22 VTAIL.n107 VTAIL.n106 185
R23 VTAIL.n96 VTAIL.n95 185
R24 VTAIL.n113 VTAIL.n112 185
R25 VTAIL.n115 VTAIL.n114 185
R26 VTAIL.n10 VTAIL.n9 185
R27 VTAIL.n15 VTAIL.n14 185
R28 VTAIL.n17 VTAIL.n16 185
R29 VTAIL.n6 VTAIL.n5 185
R30 VTAIL.n23 VTAIL.n22 185
R31 VTAIL.n25 VTAIL.n24 185
R32 VTAIL.n87 VTAIL.n86 185
R33 VTAIL.n85 VTAIL.n84 185
R34 VTAIL.n68 VTAIL.n67 185
R35 VTAIL.n79 VTAIL.n78 185
R36 VTAIL.n77 VTAIL.n76 185
R37 VTAIL.n72 VTAIL.n71 185
R38 VTAIL.n57 VTAIL.n56 185
R39 VTAIL.n55 VTAIL.n54 185
R40 VTAIL.n38 VTAIL.n37 185
R41 VTAIL.n49 VTAIL.n48 185
R42 VTAIL.n47 VTAIL.n46 185
R43 VTAIL.n42 VTAIL.n41 185
R44 VTAIL.n101 VTAIL.t9 147.672
R45 VTAIL.n11 VTAIL.t4 147.672
R46 VTAIL.n73 VTAIL.t2 147.672
R47 VTAIL.n43 VTAIL.t8 147.672
R48 VTAIL.n105 VTAIL.n99 104.615
R49 VTAIL.n106 VTAIL.n105 104.615
R50 VTAIL.n106 VTAIL.n95 104.615
R51 VTAIL.n113 VTAIL.n95 104.615
R52 VTAIL.n114 VTAIL.n113 104.615
R53 VTAIL.n15 VTAIL.n9 104.615
R54 VTAIL.n16 VTAIL.n15 104.615
R55 VTAIL.n16 VTAIL.n5 104.615
R56 VTAIL.n23 VTAIL.n5 104.615
R57 VTAIL.n24 VTAIL.n23 104.615
R58 VTAIL.n86 VTAIL.n85 104.615
R59 VTAIL.n85 VTAIL.n67 104.615
R60 VTAIL.n78 VTAIL.n67 104.615
R61 VTAIL.n78 VTAIL.n77 104.615
R62 VTAIL.n77 VTAIL.n71 104.615
R63 VTAIL.n56 VTAIL.n55 104.615
R64 VTAIL.n55 VTAIL.n37 104.615
R65 VTAIL.n48 VTAIL.n37 104.615
R66 VTAIL.n48 VTAIL.n47 104.615
R67 VTAIL.n47 VTAIL.n41 104.615
R68 VTAIL.t9 VTAIL.n99 52.3082
R69 VTAIL.t4 VTAIL.n9 52.3082
R70 VTAIL.t2 VTAIL.n71 52.3082
R71 VTAIL.t8 VTAIL.n41 52.3082
R72 VTAIL.n63 VTAIL.n62 49.8431
R73 VTAIL.n33 VTAIL.n32 49.8431
R74 VTAIL.n1 VTAIL.n0 49.843
R75 VTAIL.n31 VTAIL.n30 49.843
R76 VTAIL.n119 VTAIL.n118 30.052
R77 VTAIL.n29 VTAIL.n28 30.052
R78 VTAIL.n91 VTAIL.n90 30.052
R79 VTAIL.n61 VTAIL.n60 30.052
R80 VTAIL.n33 VTAIL.n31 17.9789
R81 VTAIL.n119 VTAIL.n91 17.4014
R82 VTAIL.n101 VTAIL.n100 15.6666
R83 VTAIL.n11 VTAIL.n10 15.6666
R84 VTAIL.n73 VTAIL.n72 15.6666
R85 VTAIL.n43 VTAIL.n42 15.6666
R86 VTAIL.n104 VTAIL.n103 12.8005
R87 VTAIL.n14 VTAIL.n13 12.8005
R88 VTAIL.n76 VTAIL.n75 12.8005
R89 VTAIL.n46 VTAIL.n45 12.8005
R90 VTAIL.n107 VTAIL.n98 12.0247
R91 VTAIL.n17 VTAIL.n8 12.0247
R92 VTAIL.n79 VTAIL.n70 12.0247
R93 VTAIL.n49 VTAIL.n40 12.0247
R94 VTAIL.n108 VTAIL.n96 11.249
R95 VTAIL.n18 VTAIL.n6 11.249
R96 VTAIL.n80 VTAIL.n68 11.249
R97 VTAIL.n50 VTAIL.n38 11.249
R98 VTAIL.n112 VTAIL.n111 10.4732
R99 VTAIL.n22 VTAIL.n21 10.4732
R100 VTAIL.n84 VTAIL.n83 10.4732
R101 VTAIL.n54 VTAIL.n53 10.4732
R102 VTAIL.n115 VTAIL.n94 9.69747
R103 VTAIL.n25 VTAIL.n4 9.69747
R104 VTAIL.n87 VTAIL.n66 9.69747
R105 VTAIL.n57 VTAIL.n36 9.69747
R106 VTAIL.n118 VTAIL.n117 9.45567
R107 VTAIL.n28 VTAIL.n27 9.45567
R108 VTAIL.n90 VTAIL.n89 9.45567
R109 VTAIL.n60 VTAIL.n59 9.45567
R110 VTAIL.n117 VTAIL.n116 9.3005
R111 VTAIL.n94 VTAIL.n93 9.3005
R112 VTAIL.n111 VTAIL.n110 9.3005
R113 VTAIL.n109 VTAIL.n108 9.3005
R114 VTAIL.n98 VTAIL.n97 9.3005
R115 VTAIL.n103 VTAIL.n102 9.3005
R116 VTAIL.n27 VTAIL.n26 9.3005
R117 VTAIL.n4 VTAIL.n3 9.3005
R118 VTAIL.n21 VTAIL.n20 9.3005
R119 VTAIL.n19 VTAIL.n18 9.3005
R120 VTAIL.n8 VTAIL.n7 9.3005
R121 VTAIL.n13 VTAIL.n12 9.3005
R122 VTAIL.n89 VTAIL.n88 9.3005
R123 VTAIL.n66 VTAIL.n65 9.3005
R124 VTAIL.n83 VTAIL.n82 9.3005
R125 VTAIL.n81 VTAIL.n80 9.3005
R126 VTAIL.n70 VTAIL.n69 9.3005
R127 VTAIL.n75 VTAIL.n74 9.3005
R128 VTAIL.n59 VTAIL.n58 9.3005
R129 VTAIL.n36 VTAIL.n35 9.3005
R130 VTAIL.n53 VTAIL.n52 9.3005
R131 VTAIL.n51 VTAIL.n50 9.3005
R132 VTAIL.n40 VTAIL.n39 9.3005
R133 VTAIL.n45 VTAIL.n44 9.3005
R134 VTAIL.n116 VTAIL.n92 8.92171
R135 VTAIL.n26 VTAIL.n2 8.92171
R136 VTAIL.n88 VTAIL.n64 8.92171
R137 VTAIL.n58 VTAIL.n34 8.92171
R138 VTAIL.n118 VTAIL.n92 5.04292
R139 VTAIL.n28 VTAIL.n2 5.04292
R140 VTAIL.n90 VTAIL.n64 5.04292
R141 VTAIL.n60 VTAIL.n34 5.04292
R142 VTAIL.n102 VTAIL.n101 4.38687
R143 VTAIL.n12 VTAIL.n11 4.38687
R144 VTAIL.n74 VTAIL.n73 4.38687
R145 VTAIL.n44 VTAIL.n43 4.38687
R146 VTAIL.n116 VTAIL.n115 4.26717
R147 VTAIL.n26 VTAIL.n25 4.26717
R148 VTAIL.n88 VTAIL.n87 4.26717
R149 VTAIL.n58 VTAIL.n57 4.26717
R150 VTAIL.n0 VTAIL.t11 3.83029
R151 VTAIL.n0 VTAIL.t7 3.83029
R152 VTAIL.n30 VTAIL.t1 3.83029
R153 VTAIL.n30 VTAIL.t0 3.83029
R154 VTAIL.n62 VTAIL.t3 3.83029
R155 VTAIL.n62 VTAIL.t5 3.83029
R156 VTAIL.n32 VTAIL.t6 3.83029
R157 VTAIL.n32 VTAIL.t10 3.83029
R158 VTAIL.n112 VTAIL.n94 3.49141
R159 VTAIL.n22 VTAIL.n4 3.49141
R160 VTAIL.n84 VTAIL.n66 3.49141
R161 VTAIL.n54 VTAIL.n36 3.49141
R162 VTAIL.n111 VTAIL.n96 2.71565
R163 VTAIL.n21 VTAIL.n6 2.71565
R164 VTAIL.n83 VTAIL.n68 2.71565
R165 VTAIL.n53 VTAIL.n38 2.71565
R166 VTAIL.n108 VTAIL.n107 1.93989
R167 VTAIL.n18 VTAIL.n17 1.93989
R168 VTAIL.n80 VTAIL.n79 1.93989
R169 VTAIL.n50 VTAIL.n49 1.93989
R170 VTAIL.n104 VTAIL.n98 1.16414
R171 VTAIL.n14 VTAIL.n8 1.16414
R172 VTAIL.n76 VTAIL.n70 1.16414
R173 VTAIL.n46 VTAIL.n40 1.16414
R174 VTAIL.n63 VTAIL.n61 0.759121
R175 VTAIL.n29 VTAIL.n1 0.759121
R176 VTAIL.n61 VTAIL.n33 0.578086
R177 VTAIL.n91 VTAIL.n63 0.578086
R178 VTAIL.n31 VTAIL.n29 0.578086
R179 VTAIL.n103 VTAIL.n100 0.388379
R180 VTAIL.n13 VTAIL.n10 0.388379
R181 VTAIL.n75 VTAIL.n72 0.388379
R182 VTAIL.n45 VTAIL.n42 0.388379
R183 VTAIL VTAIL.n119 0.3755
R184 VTAIL VTAIL.n1 0.203086
R185 VTAIL.n102 VTAIL.n97 0.155672
R186 VTAIL.n109 VTAIL.n97 0.155672
R187 VTAIL.n110 VTAIL.n109 0.155672
R188 VTAIL.n110 VTAIL.n93 0.155672
R189 VTAIL.n117 VTAIL.n93 0.155672
R190 VTAIL.n12 VTAIL.n7 0.155672
R191 VTAIL.n19 VTAIL.n7 0.155672
R192 VTAIL.n20 VTAIL.n19 0.155672
R193 VTAIL.n20 VTAIL.n3 0.155672
R194 VTAIL.n27 VTAIL.n3 0.155672
R195 VTAIL.n89 VTAIL.n65 0.155672
R196 VTAIL.n82 VTAIL.n65 0.155672
R197 VTAIL.n82 VTAIL.n81 0.155672
R198 VTAIL.n81 VTAIL.n69 0.155672
R199 VTAIL.n74 VTAIL.n69 0.155672
R200 VTAIL.n59 VTAIL.n35 0.155672
R201 VTAIL.n52 VTAIL.n35 0.155672
R202 VTAIL.n52 VTAIL.n51 0.155672
R203 VTAIL.n51 VTAIL.n39 0.155672
R204 VTAIL.n44 VTAIL.n39 0.155672
R205 VDD2.n51 VDD2.n29 289.615
R206 VDD2.n22 VDD2.n0 289.615
R207 VDD2.n52 VDD2.n51 185
R208 VDD2.n50 VDD2.n49 185
R209 VDD2.n33 VDD2.n32 185
R210 VDD2.n44 VDD2.n43 185
R211 VDD2.n42 VDD2.n41 185
R212 VDD2.n37 VDD2.n36 185
R213 VDD2.n8 VDD2.n7 185
R214 VDD2.n13 VDD2.n12 185
R215 VDD2.n15 VDD2.n14 185
R216 VDD2.n4 VDD2.n3 185
R217 VDD2.n21 VDD2.n20 185
R218 VDD2.n23 VDD2.n22 185
R219 VDD2.n38 VDD2.t4 147.672
R220 VDD2.n9 VDD2.t1 147.672
R221 VDD2.n51 VDD2.n50 104.615
R222 VDD2.n50 VDD2.n32 104.615
R223 VDD2.n43 VDD2.n32 104.615
R224 VDD2.n43 VDD2.n42 104.615
R225 VDD2.n42 VDD2.n36 104.615
R226 VDD2.n13 VDD2.n7 104.615
R227 VDD2.n14 VDD2.n13 104.615
R228 VDD2.n14 VDD2.n3 104.615
R229 VDD2.n21 VDD2.n3 104.615
R230 VDD2.n22 VDD2.n21 104.615
R231 VDD2.n28 VDD2.n27 66.6108
R232 VDD2 VDD2.n57 66.608
R233 VDD2.t4 VDD2.n36 52.3082
R234 VDD2.t1 VDD2.n7 52.3082
R235 VDD2.n28 VDD2.n26 47.1086
R236 VDD2.n56 VDD2.n55 46.7308
R237 VDD2.n56 VDD2.n28 30.0493
R238 VDD2.n38 VDD2.n37 15.6666
R239 VDD2.n9 VDD2.n8 15.6666
R240 VDD2.n41 VDD2.n40 12.8005
R241 VDD2.n12 VDD2.n11 12.8005
R242 VDD2.n44 VDD2.n35 12.0247
R243 VDD2.n15 VDD2.n6 12.0247
R244 VDD2.n45 VDD2.n33 11.249
R245 VDD2.n16 VDD2.n4 11.249
R246 VDD2.n49 VDD2.n48 10.4732
R247 VDD2.n20 VDD2.n19 10.4732
R248 VDD2.n52 VDD2.n31 9.69747
R249 VDD2.n23 VDD2.n2 9.69747
R250 VDD2.n55 VDD2.n54 9.45567
R251 VDD2.n26 VDD2.n25 9.45567
R252 VDD2.n54 VDD2.n53 9.3005
R253 VDD2.n31 VDD2.n30 9.3005
R254 VDD2.n48 VDD2.n47 9.3005
R255 VDD2.n46 VDD2.n45 9.3005
R256 VDD2.n35 VDD2.n34 9.3005
R257 VDD2.n40 VDD2.n39 9.3005
R258 VDD2.n25 VDD2.n24 9.3005
R259 VDD2.n2 VDD2.n1 9.3005
R260 VDD2.n19 VDD2.n18 9.3005
R261 VDD2.n17 VDD2.n16 9.3005
R262 VDD2.n6 VDD2.n5 9.3005
R263 VDD2.n11 VDD2.n10 9.3005
R264 VDD2.n53 VDD2.n29 8.92171
R265 VDD2.n24 VDD2.n0 8.92171
R266 VDD2.n55 VDD2.n29 5.04292
R267 VDD2.n26 VDD2.n0 5.04292
R268 VDD2.n39 VDD2.n38 4.38687
R269 VDD2.n10 VDD2.n9 4.38687
R270 VDD2.n53 VDD2.n52 4.26717
R271 VDD2.n24 VDD2.n23 4.26717
R272 VDD2.n57 VDD2.t2 3.83029
R273 VDD2.n57 VDD2.t0 3.83029
R274 VDD2.n27 VDD2.t3 3.83029
R275 VDD2.n27 VDD2.t5 3.83029
R276 VDD2.n49 VDD2.n31 3.49141
R277 VDD2.n20 VDD2.n2 3.49141
R278 VDD2.n48 VDD2.n33 2.71565
R279 VDD2.n19 VDD2.n4 2.71565
R280 VDD2.n45 VDD2.n44 1.93989
R281 VDD2.n16 VDD2.n15 1.93989
R282 VDD2.n41 VDD2.n35 1.16414
R283 VDD2.n12 VDD2.n6 1.16414
R284 VDD2 VDD2.n56 0.491879
R285 VDD2.n40 VDD2.n37 0.388379
R286 VDD2.n11 VDD2.n8 0.388379
R287 VDD2.n54 VDD2.n30 0.155672
R288 VDD2.n47 VDD2.n30 0.155672
R289 VDD2.n47 VDD2.n46 0.155672
R290 VDD2.n46 VDD2.n34 0.155672
R291 VDD2.n39 VDD2.n34 0.155672
R292 VDD2.n10 VDD2.n5 0.155672
R293 VDD2.n17 VDD2.n5 0.155672
R294 VDD2.n18 VDD2.n17 0.155672
R295 VDD2.n18 VDD2.n1 0.155672
R296 VDD2.n25 VDD2.n1 0.155672
R297 B.n406 B.n405 585
R298 B.n407 B.n406 585
R299 B.n167 B.n60 585
R300 B.n166 B.n165 585
R301 B.n164 B.n163 585
R302 B.n162 B.n161 585
R303 B.n160 B.n159 585
R304 B.n158 B.n157 585
R305 B.n156 B.n155 585
R306 B.n154 B.n153 585
R307 B.n152 B.n151 585
R308 B.n150 B.n149 585
R309 B.n148 B.n147 585
R310 B.n146 B.n145 585
R311 B.n144 B.n143 585
R312 B.n142 B.n141 585
R313 B.n140 B.n139 585
R314 B.n138 B.n137 585
R315 B.n136 B.n135 585
R316 B.n134 B.n133 585
R317 B.n132 B.n131 585
R318 B.n130 B.n129 585
R319 B.n128 B.n127 585
R320 B.n125 B.n124 585
R321 B.n123 B.n122 585
R322 B.n121 B.n120 585
R323 B.n119 B.n118 585
R324 B.n117 B.n116 585
R325 B.n115 B.n114 585
R326 B.n113 B.n112 585
R327 B.n111 B.n110 585
R328 B.n109 B.n108 585
R329 B.n107 B.n106 585
R330 B.n105 B.n104 585
R331 B.n103 B.n102 585
R332 B.n101 B.n100 585
R333 B.n99 B.n98 585
R334 B.n97 B.n96 585
R335 B.n95 B.n94 585
R336 B.n93 B.n92 585
R337 B.n91 B.n90 585
R338 B.n89 B.n88 585
R339 B.n87 B.n86 585
R340 B.n85 B.n84 585
R341 B.n83 B.n82 585
R342 B.n81 B.n80 585
R343 B.n79 B.n78 585
R344 B.n77 B.n76 585
R345 B.n75 B.n74 585
R346 B.n73 B.n72 585
R347 B.n71 B.n70 585
R348 B.n69 B.n68 585
R349 B.n67 B.n66 585
R350 B.n32 B.n31 585
R351 B.n404 B.n33 585
R352 B.n408 B.n33 585
R353 B.n403 B.n402 585
R354 B.n402 B.n29 585
R355 B.n401 B.n28 585
R356 B.n414 B.n28 585
R357 B.n400 B.n27 585
R358 B.n415 B.n27 585
R359 B.n399 B.n26 585
R360 B.n416 B.n26 585
R361 B.n398 B.n397 585
R362 B.n397 B.n22 585
R363 B.n396 B.n21 585
R364 B.n422 B.n21 585
R365 B.n395 B.n20 585
R366 B.n423 B.n20 585
R367 B.n394 B.n19 585
R368 B.n424 B.n19 585
R369 B.n393 B.n392 585
R370 B.n392 B.n18 585
R371 B.n391 B.n14 585
R372 B.n430 B.n14 585
R373 B.n390 B.n13 585
R374 B.n431 B.n13 585
R375 B.n389 B.n12 585
R376 B.n432 B.n12 585
R377 B.n388 B.n387 585
R378 B.n387 B.n11 585
R379 B.n386 B.n7 585
R380 B.n438 B.n7 585
R381 B.n385 B.n6 585
R382 B.n439 B.n6 585
R383 B.n384 B.n5 585
R384 B.n440 B.n5 585
R385 B.n383 B.n382 585
R386 B.n382 B.n4 585
R387 B.n381 B.n168 585
R388 B.n381 B.n380 585
R389 B.n370 B.n169 585
R390 B.n373 B.n169 585
R391 B.n372 B.n371 585
R392 B.n374 B.n372 585
R393 B.n369 B.n173 585
R394 B.n176 B.n173 585
R395 B.n368 B.n367 585
R396 B.n367 B.n366 585
R397 B.n175 B.n174 585
R398 B.n359 B.n175 585
R399 B.n358 B.n357 585
R400 B.n360 B.n358 585
R401 B.n356 B.n181 585
R402 B.n181 B.n180 585
R403 B.n355 B.n354 585
R404 B.n354 B.n353 585
R405 B.n183 B.n182 585
R406 B.n184 B.n183 585
R407 B.n346 B.n345 585
R408 B.n347 B.n346 585
R409 B.n344 B.n189 585
R410 B.n189 B.n188 585
R411 B.n343 B.n342 585
R412 B.n342 B.n341 585
R413 B.n191 B.n190 585
R414 B.n192 B.n191 585
R415 B.n334 B.n333 585
R416 B.n335 B.n334 585
R417 B.n195 B.n194 585
R418 B.n228 B.n226 585
R419 B.n229 B.n225 585
R420 B.n229 B.n196 585
R421 B.n232 B.n231 585
R422 B.n233 B.n224 585
R423 B.n235 B.n234 585
R424 B.n237 B.n223 585
R425 B.n240 B.n239 585
R426 B.n241 B.n222 585
R427 B.n243 B.n242 585
R428 B.n245 B.n221 585
R429 B.n248 B.n247 585
R430 B.n249 B.n220 585
R431 B.n251 B.n250 585
R432 B.n253 B.n219 585
R433 B.n256 B.n255 585
R434 B.n257 B.n218 585
R435 B.n259 B.n258 585
R436 B.n261 B.n217 585
R437 B.n264 B.n263 585
R438 B.n265 B.n216 585
R439 B.n270 B.n269 585
R440 B.n272 B.n215 585
R441 B.n275 B.n274 585
R442 B.n276 B.n214 585
R443 B.n278 B.n277 585
R444 B.n280 B.n213 585
R445 B.n283 B.n282 585
R446 B.n284 B.n212 585
R447 B.n286 B.n285 585
R448 B.n288 B.n211 585
R449 B.n291 B.n290 585
R450 B.n292 B.n207 585
R451 B.n294 B.n293 585
R452 B.n296 B.n206 585
R453 B.n299 B.n298 585
R454 B.n300 B.n205 585
R455 B.n302 B.n301 585
R456 B.n304 B.n204 585
R457 B.n307 B.n306 585
R458 B.n308 B.n203 585
R459 B.n310 B.n309 585
R460 B.n312 B.n202 585
R461 B.n315 B.n314 585
R462 B.n316 B.n201 585
R463 B.n318 B.n317 585
R464 B.n320 B.n200 585
R465 B.n323 B.n322 585
R466 B.n324 B.n199 585
R467 B.n326 B.n325 585
R468 B.n328 B.n198 585
R469 B.n331 B.n330 585
R470 B.n332 B.n197 585
R471 B.n337 B.n336 585
R472 B.n336 B.n335 585
R473 B.n338 B.n193 585
R474 B.n193 B.n192 585
R475 B.n340 B.n339 585
R476 B.n341 B.n340 585
R477 B.n187 B.n186 585
R478 B.n188 B.n187 585
R479 B.n349 B.n348 585
R480 B.n348 B.n347 585
R481 B.n350 B.n185 585
R482 B.n185 B.n184 585
R483 B.n352 B.n351 585
R484 B.n353 B.n352 585
R485 B.n179 B.n178 585
R486 B.n180 B.n179 585
R487 B.n362 B.n361 585
R488 B.n361 B.n360 585
R489 B.n363 B.n177 585
R490 B.n359 B.n177 585
R491 B.n365 B.n364 585
R492 B.n366 B.n365 585
R493 B.n172 B.n171 585
R494 B.n176 B.n172 585
R495 B.n376 B.n375 585
R496 B.n375 B.n374 585
R497 B.n377 B.n170 585
R498 B.n373 B.n170 585
R499 B.n379 B.n378 585
R500 B.n380 B.n379 585
R501 B.n2 B.n0 585
R502 B.n4 B.n2 585
R503 B.n3 B.n1 585
R504 B.n439 B.n3 585
R505 B.n437 B.n436 585
R506 B.n438 B.n437 585
R507 B.n435 B.n8 585
R508 B.n11 B.n8 585
R509 B.n434 B.n433 585
R510 B.n433 B.n432 585
R511 B.n10 B.n9 585
R512 B.n431 B.n10 585
R513 B.n429 B.n428 585
R514 B.n430 B.n429 585
R515 B.n427 B.n15 585
R516 B.n18 B.n15 585
R517 B.n426 B.n425 585
R518 B.n425 B.n424 585
R519 B.n17 B.n16 585
R520 B.n423 B.n17 585
R521 B.n421 B.n420 585
R522 B.n422 B.n421 585
R523 B.n419 B.n23 585
R524 B.n23 B.n22 585
R525 B.n418 B.n417 585
R526 B.n417 B.n416 585
R527 B.n25 B.n24 585
R528 B.n415 B.n25 585
R529 B.n413 B.n412 585
R530 B.n414 B.n413 585
R531 B.n411 B.n30 585
R532 B.n30 B.n29 585
R533 B.n410 B.n409 585
R534 B.n409 B.n408 585
R535 B.n442 B.n441 585
R536 B.n441 B.n440 585
R537 B.n208 B.t6 578.54
R538 B.n266 B.t17 578.54
R539 B.n63 B.t14 578.54
R540 B.n61 B.t10 578.54
R541 B.n336 B.n195 468.476
R542 B.n409 B.n32 468.476
R543 B.n334 B.n197 468.476
R544 B.n406 B.n33 468.476
R545 B.n407 B.n59 256.663
R546 B.n407 B.n58 256.663
R547 B.n407 B.n57 256.663
R548 B.n407 B.n56 256.663
R549 B.n407 B.n55 256.663
R550 B.n407 B.n54 256.663
R551 B.n407 B.n53 256.663
R552 B.n407 B.n52 256.663
R553 B.n407 B.n51 256.663
R554 B.n407 B.n50 256.663
R555 B.n407 B.n49 256.663
R556 B.n407 B.n48 256.663
R557 B.n407 B.n47 256.663
R558 B.n407 B.n46 256.663
R559 B.n407 B.n45 256.663
R560 B.n407 B.n44 256.663
R561 B.n407 B.n43 256.663
R562 B.n407 B.n42 256.663
R563 B.n407 B.n41 256.663
R564 B.n407 B.n40 256.663
R565 B.n407 B.n39 256.663
R566 B.n407 B.n38 256.663
R567 B.n407 B.n37 256.663
R568 B.n407 B.n36 256.663
R569 B.n407 B.n35 256.663
R570 B.n407 B.n34 256.663
R571 B.n227 B.n196 256.663
R572 B.n230 B.n196 256.663
R573 B.n236 B.n196 256.663
R574 B.n238 B.n196 256.663
R575 B.n244 B.n196 256.663
R576 B.n246 B.n196 256.663
R577 B.n252 B.n196 256.663
R578 B.n254 B.n196 256.663
R579 B.n260 B.n196 256.663
R580 B.n262 B.n196 256.663
R581 B.n271 B.n196 256.663
R582 B.n273 B.n196 256.663
R583 B.n279 B.n196 256.663
R584 B.n281 B.n196 256.663
R585 B.n287 B.n196 256.663
R586 B.n289 B.n196 256.663
R587 B.n295 B.n196 256.663
R588 B.n297 B.n196 256.663
R589 B.n303 B.n196 256.663
R590 B.n305 B.n196 256.663
R591 B.n311 B.n196 256.663
R592 B.n313 B.n196 256.663
R593 B.n319 B.n196 256.663
R594 B.n321 B.n196 256.663
R595 B.n327 B.n196 256.663
R596 B.n329 B.n196 256.663
R597 B.n208 B.t9 177.435
R598 B.n61 B.t12 177.435
R599 B.n266 B.t19 177.435
R600 B.n63 B.t15 177.435
R601 B.n209 B.t8 164.44
R602 B.n62 B.t13 164.44
R603 B.n267 B.t18 164.44
R604 B.n64 B.t16 164.44
R605 B.n336 B.n193 163.367
R606 B.n340 B.n193 163.367
R607 B.n340 B.n187 163.367
R608 B.n348 B.n187 163.367
R609 B.n348 B.n185 163.367
R610 B.n352 B.n185 163.367
R611 B.n352 B.n179 163.367
R612 B.n361 B.n179 163.367
R613 B.n361 B.n177 163.367
R614 B.n365 B.n177 163.367
R615 B.n365 B.n172 163.367
R616 B.n375 B.n172 163.367
R617 B.n375 B.n170 163.367
R618 B.n379 B.n170 163.367
R619 B.n379 B.n2 163.367
R620 B.n441 B.n2 163.367
R621 B.n441 B.n3 163.367
R622 B.n437 B.n3 163.367
R623 B.n437 B.n8 163.367
R624 B.n433 B.n8 163.367
R625 B.n433 B.n10 163.367
R626 B.n429 B.n10 163.367
R627 B.n429 B.n15 163.367
R628 B.n425 B.n15 163.367
R629 B.n425 B.n17 163.367
R630 B.n421 B.n17 163.367
R631 B.n421 B.n23 163.367
R632 B.n417 B.n23 163.367
R633 B.n417 B.n25 163.367
R634 B.n413 B.n25 163.367
R635 B.n413 B.n30 163.367
R636 B.n409 B.n30 163.367
R637 B.n229 B.n228 163.367
R638 B.n231 B.n229 163.367
R639 B.n235 B.n224 163.367
R640 B.n239 B.n237 163.367
R641 B.n243 B.n222 163.367
R642 B.n247 B.n245 163.367
R643 B.n251 B.n220 163.367
R644 B.n255 B.n253 163.367
R645 B.n259 B.n218 163.367
R646 B.n263 B.n261 163.367
R647 B.n270 B.n216 163.367
R648 B.n274 B.n272 163.367
R649 B.n278 B.n214 163.367
R650 B.n282 B.n280 163.367
R651 B.n286 B.n212 163.367
R652 B.n290 B.n288 163.367
R653 B.n294 B.n207 163.367
R654 B.n298 B.n296 163.367
R655 B.n302 B.n205 163.367
R656 B.n306 B.n304 163.367
R657 B.n310 B.n203 163.367
R658 B.n314 B.n312 163.367
R659 B.n318 B.n201 163.367
R660 B.n322 B.n320 163.367
R661 B.n326 B.n199 163.367
R662 B.n330 B.n328 163.367
R663 B.n334 B.n191 163.367
R664 B.n342 B.n191 163.367
R665 B.n342 B.n189 163.367
R666 B.n346 B.n189 163.367
R667 B.n346 B.n183 163.367
R668 B.n354 B.n183 163.367
R669 B.n354 B.n181 163.367
R670 B.n358 B.n181 163.367
R671 B.n358 B.n175 163.367
R672 B.n367 B.n175 163.367
R673 B.n367 B.n173 163.367
R674 B.n372 B.n173 163.367
R675 B.n372 B.n169 163.367
R676 B.n381 B.n169 163.367
R677 B.n382 B.n381 163.367
R678 B.n382 B.n5 163.367
R679 B.n6 B.n5 163.367
R680 B.n7 B.n6 163.367
R681 B.n387 B.n7 163.367
R682 B.n387 B.n12 163.367
R683 B.n13 B.n12 163.367
R684 B.n14 B.n13 163.367
R685 B.n392 B.n14 163.367
R686 B.n392 B.n19 163.367
R687 B.n20 B.n19 163.367
R688 B.n21 B.n20 163.367
R689 B.n397 B.n21 163.367
R690 B.n397 B.n26 163.367
R691 B.n27 B.n26 163.367
R692 B.n28 B.n27 163.367
R693 B.n402 B.n28 163.367
R694 B.n402 B.n33 163.367
R695 B.n68 B.n67 163.367
R696 B.n72 B.n71 163.367
R697 B.n76 B.n75 163.367
R698 B.n80 B.n79 163.367
R699 B.n84 B.n83 163.367
R700 B.n88 B.n87 163.367
R701 B.n92 B.n91 163.367
R702 B.n96 B.n95 163.367
R703 B.n100 B.n99 163.367
R704 B.n104 B.n103 163.367
R705 B.n108 B.n107 163.367
R706 B.n112 B.n111 163.367
R707 B.n116 B.n115 163.367
R708 B.n120 B.n119 163.367
R709 B.n124 B.n123 163.367
R710 B.n129 B.n128 163.367
R711 B.n133 B.n132 163.367
R712 B.n137 B.n136 163.367
R713 B.n141 B.n140 163.367
R714 B.n145 B.n144 163.367
R715 B.n149 B.n148 163.367
R716 B.n153 B.n152 163.367
R717 B.n157 B.n156 163.367
R718 B.n161 B.n160 163.367
R719 B.n165 B.n164 163.367
R720 B.n406 B.n60 163.367
R721 B.n335 B.n196 129.536
R722 B.n408 B.n407 129.536
R723 B.n227 B.n195 71.676
R724 B.n231 B.n230 71.676
R725 B.n236 B.n235 71.676
R726 B.n239 B.n238 71.676
R727 B.n244 B.n243 71.676
R728 B.n247 B.n246 71.676
R729 B.n252 B.n251 71.676
R730 B.n255 B.n254 71.676
R731 B.n260 B.n259 71.676
R732 B.n263 B.n262 71.676
R733 B.n271 B.n270 71.676
R734 B.n274 B.n273 71.676
R735 B.n279 B.n278 71.676
R736 B.n282 B.n281 71.676
R737 B.n287 B.n286 71.676
R738 B.n290 B.n289 71.676
R739 B.n295 B.n294 71.676
R740 B.n298 B.n297 71.676
R741 B.n303 B.n302 71.676
R742 B.n306 B.n305 71.676
R743 B.n311 B.n310 71.676
R744 B.n314 B.n313 71.676
R745 B.n319 B.n318 71.676
R746 B.n322 B.n321 71.676
R747 B.n327 B.n326 71.676
R748 B.n330 B.n329 71.676
R749 B.n34 B.n32 71.676
R750 B.n68 B.n35 71.676
R751 B.n72 B.n36 71.676
R752 B.n76 B.n37 71.676
R753 B.n80 B.n38 71.676
R754 B.n84 B.n39 71.676
R755 B.n88 B.n40 71.676
R756 B.n92 B.n41 71.676
R757 B.n96 B.n42 71.676
R758 B.n100 B.n43 71.676
R759 B.n104 B.n44 71.676
R760 B.n108 B.n45 71.676
R761 B.n112 B.n46 71.676
R762 B.n116 B.n47 71.676
R763 B.n120 B.n48 71.676
R764 B.n124 B.n49 71.676
R765 B.n129 B.n50 71.676
R766 B.n133 B.n51 71.676
R767 B.n137 B.n52 71.676
R768 B.n141 B.n53 71.676
R769 B.n145 B.n54 71.676
R770 B.n149 B.n55 71.676
R771 B.n153 B.n56 71.676
R772 B.n157 B.n57 71.676
R773 B.n161 B.n58 71.676
R774 B.n165 B.n59 71.676
R775 B.n60 B.n59 71.676
R776 B.n164 B.n58 71.676
R777 B.n160 B.n57 71.676
R778 B.n156 B.n56 71.676
R779 B.n152 B.n55 71.676
R780 B.n148 B.n54 71.676
R781 B.n144 B.n53 71.676
R782 B.n140 B.n52 71.676
R783 B.n136 B.n51 71.676
R784 B.n132 B.n50 71.676
R785 B.n128 B.n49 71.676
R786 B.n123 B.n48 71.676
R787 B.n119 B.n47 71.676
R788 B.n115 B.n46 71.676
R789 B.n111 B.n45 71.676
R790 B.n107 B.n44 71.676
R791 B.n103 B.n43 71.676
R792 B.n99 B.n42 71.676
R793 B.n95 B.n41 71.676
R794 B.n91 B.n40 71.676
R795 B.n87 B.n39 71.676
R796 B.n83 B.n38 71.676
R797 B.n79 B.n37 71.676
R798 B.n75 B.n36 71.676
R799 B.n71 B.n35 71.676
R800 B.n67 B.n34 71.676
R801 B.n228 B.n227 71.676
R802 B.n230 B.n224 71.676
R803 B.n237 B.n236 71.676
R804 B.n238 B.n222 71.676
R805 B.n245 B.n244 71.676
R806 B.n246 B.n220 71.676
R807 B.n253 B.n252 71.676
R808 B.n254 B.n218 71.676
R809 B.n261 B.n260 71.676
R810 B.n262 B.n216 71.676
R811 B.n272 B.n271 71.676
R812 B.n273 B.n214 71.676
R813 B.n280 B.n279 71.676
R814 B.n281 B.n212 71.676
R815 B.n288 B.n287 71.676
R816 B.n289 B.n207 71.676
R817 B.n296 B.n295 71.676
R818 B.n297 B.n205 71.676
R819 B.n304 B.n303 71.676
R820 B.n305 B.n203 71.676
R821 B.n312 B.n311 71.676
R822 B.n313 B.n201 71.676
R823 B.n320 B.n319 71.676
R824 B.n321 B.n199 71.676
R825 B.n328 B.n327 71.676
R826 B.n329 B.n197 71.676
R827 B.n335 B.n192 71.6137
R828 B.n341 B.n192 71.6137
R829 B.n341 B.n188 71.6137
R830 B.n347 B.n188 71.6137
R831 B.n353 B.n184 71.6137
R832 B.n353 B.n180 71.6137
R833 B.n360 B.n180 71.6137
R834 B.n360 B.n359 71.6137
R835 B.n366 B.n176 71.6137
R836 B.n374 B.n373 71.6137
R837 B.n380 B.n4 71.6137
R838 B.n440 B.n4 71.6137
R839 B.n440 B.n439 71.6137
R840 B.n439 B.n438 71.6137
R841 B.n432 B.n11 71.6137
R842 B.n431 B.n430 71.6137
R843 B.n424 B.n18 71.6137
R844 B.n424 B.n423 71.6137
R845 B.n423 B.n422 71.6137
R846 B.n422 B.n22 71.6137
R847 B.n416 B.n415 71.6137
R848 B.n415 B.n414 71.6137
R849 B.n414 B.n29 71.6137
R850 B.n408 B.n29 71.6137
R851 B.n210 B.n209 59.5399
R852 B.n268 B.n267 59.5399
R853 B.n65 B.n64 59.5399
R854 B.n126 B.n62 59.5399
R855 B.t7 B.n184 50.551
R856 B.t11 B.n22 50.551
R857 B.n380 B.t4 42.1259
R858 B.n438 B.t3 42.1259
R859 B.n374 B.t0 40.0196
R860 B.n432 B.t5 40.0196
R861 B.n366 B.t1 37.9134
R862 B.n430 B.t2 37.9134
R863 B.n359 B.t1 33.7008
R864 B.n18 B.t2 33.7008
R865 B.n176 B.t0 31.5946
R866 B.t5 B.n431 31.5946
R867 B.n410 B.n31 30.4395
R868 B.n405 B.n404 30.4395
R869 B.n333 B.n332 30.4395
R870 B.n337 B.n194 30.4395
R871 B.n373 B.t4 29.4883
R872 B.n11 B.t3 29.4883
R873 B.n347 B.t7 21.0632
R874 B.n416 B.t11 21.0632
R875 B B.n442 18.0485
R876 B.n209 B.n208 12.9944
R877 B.n267 B.n266 12.9944
R878 B.n64 B.n63 12.9944
R879 B.n62 B.n61 12.9944
R880 B.n66 B.n31 10.6151
R881 B.n69 B.n66 10.6151
R882 B.n70 B.n69 10.6151
R883 B.n73 B.n70 10.6151
R884 B.n74 B.n73 10.6151
R885 B.n77 B.n74 10.6151
R886 B.n78 B.n77 10.6151
R887 B.n81 B.n78 10.6151
R888 B.n82 B.n81 10.6151
R889 B.n85 B.n82 10.6151
R890 B.n86 B.n85 10.6151
R891 B.n89 B.n86 10.6151
R892 B.n90 B.n89 10.6151
R893 B.n93 B.n90 10.6151
R894 B.n94 B.n93 10.6151
R895 B.n97 B.n94 10.6151
R896 B.n98 B.n97 10.6151
R897 B.n101 B.n98 10.6151
R898 B.n102 B.n101 10.6151
R899 B.n105 B.n102 10.6151
R900 B.n106 B.n105 10.6151
R901 B.n110 B.n109 10.6151
R902 B.n113 B.n110 10.6151
R903 B.n114 B.n113 10.6151
R904 B.n117 B.n114 10.6151
R905 B.n118 B.n117 10.6151
R906 B.n121 B.n118 10.6151
R907 B.n122 B.n121 10.6151
R908 B.n125 B.n122 10.6151
R909 B.n130 B.n127 10.6151
R910 B.n131 B.n130 10.6151
R911 B.n134 B.n131 10.6151
R912 B.n135 B.n134 10.6151
R913 B.n138 B.n135 10.6151
R914 B.n139 B.n138 10.6151
R915 B.n142 B.n139 10.6151
R916 B.n143 B.n142 10.6151
R917 B.n146 B.n143 10.6151
R918 B.n147 B.n146 10.6151
R919 B.n150 B.n147 10.6151
R920 B.n151 B.n150 10.6151
R921 B.n154 B.n151 10.6151
R922 B.n155 B.n154 10.6151
R923 B.n158 B.n155 10.6151
R924 B.n159 B.n158 10.6151
R925 B.n162 B.n159 10.6151
R926 B.n163 B.n162 10.6151
R927 B.n166 B.n163 10.6151
R928 B.n167 B.n166 10.6151
R929 B.n405 B.n167 10.6151
R930 B.n333 B.n190 10.6151
R931 B.n343 B.n190 10.6151
R932 B.n344 B.n343 10.6151
R933 B.n345 B.n344 10.6151
R934 B.n345 B.n182 10.6151
R935 B.n355 B.n182 10.6151
R936 B.n356 B.n355 10.6151
R937 B.n357 B.n356 10.6151
R938 B.n357 B.n174 10.6151
R939 B.n368 B.n174 10.6151
R940 B.n369 B.n368 10.6151
R941 B.n371 B.n369 10.6151
R942 B.n371 B.n370 10.6151
R943 B.n370 B.n168 10.6151
R944 B.n383 B.n168 10.6151
R945 B.n384 B.n383 10.6151
R946 B.n385 B.n384 10.6151
R947 B.n386 B.n385 10.6151
R948 B.n388 B.n386 10.6151
R949 B.n389 B.n388 10.6151
R950 B.n390 B.n389 10.6151
R951 B.n391 B.n390 10.6151
R952 B.n393 B.n391 10.6151
R953 B.n394 B.n393 10.6151
R954 B.n395 B.n394 10.6151
R955 B.n396 B.n395 10.6151
R956 B.n398 B.n396 10.6151
R957 B.n399 B.n398 10.6151
R958 B.n400 B.n399 10.6151
R959 B.n401 B.n400 10.6151
R960 B.n403 B.n401 10.6151
R961 B.n404 B.n403 10.6151
R962 B.n226 B.n194 10.6151
R963 B.n226 B.n225 10.6151
R964 B.n232 B.n225 10.6151
R965 B.n233 B.n232 10.6151
R966 B.n234 B.n233 10.6151
R967 B.n234 B.n223 10.6151
R968 B.n240 B.n223 10.6151
R969 B.n241 B.n240 10.6151
R970 B.n242 B.n241 10.6151
R971 B.n242 B.n221 10.6151
R972 B.n248 B.n221 10.6151
R973 B.n249 B.n248 10.6151
R974 B.n250 B.n249 10.6151
R975 B.n250 B.n219 10.6151
R976 B.n256 B.n219 10.6151
R977 B.n257 B.n256 10.6151
R978 B.n258 B.n257 10.6151
R979 B.n258 B.n217 10.6151
R980 B.n264 B.n217 10.6151
R981 B.n265 B.n264 10.6151
R982 B.n269 B.n265 10.6151
R983 B.n275 B.n215 10.6151
R984 B.n276 B.n275 10.6151
R985 B.n277 B.n276 10.6151
R986 B.n277 B.n213 10.6151
R987 B.n283 B.n213 10.6151
R988 B.n284 B.n283 10.6151
R989 B.n285 B.n284 10.6151
R990 B.n285 B.n211 10.6151
R991 B.n292 B.n291 10.6151
R992 B.n293 B.n292 10.6151
R993 B.n293 B.n206 10.6151
R994 B.n299 B.n206 10.6151
R995 B.n300 B.n299 10.6151
R996 B.n301 B.n300 10.6151
R997 B.n301 B.n204 10.6151
R998 B.n307 B.n204 10.6151
R999 B.n308 B.n307 10.6151
R1000 B.n309 B.n308 10.6151
R1001 B.n309 B.n202 10.6151
R1002 B.n315 B.n202 10.6151
R1003 B.n316 B.n315 10.6151
R1004 B.n317 B.n316 10.6151
R1005 B.n317 B.n200 10.6151
R1006 B.n323 B.n200 10.6151
R1007 B.n324 B.n323 10.6151
R1008 B.n325 B.n324 10.6151
R1009 B.n325 B.n198 10.6151
R1010 B.n331 B.n198 10.6151
R1011 B.n332 B.n331 10.6151
R1012 B.n338 B.n337 10.6151
R1013 B.n339 B.n338 10.6151
R1014 B.n339 B.n186 10.6151
R1015 B.n349 B.n186 10.6151
R1016 B.n350 B.n349 10.6151
R1017 B.n351 B.n350 10.6151
R1018 B.n351 B.n178 10.6151
R1019 B.n362 B.n178 10.6151
R1020 B.n363 B.n362 10.6151
R1021 B.n364 B.n363 10.6151
R1022 B.n364 B.n171 10.6151
R1023 B.n376 B.n171 10.6151
R1024 B.n377 B.n376 10.6151
R1025 B.n378 B.n377 10.6151
R1026 B.n378 B.n0 10.6151
R1027 B.n436 B.n1 10.6151
R1028 B.n436 B.n435 10.6151
R1029 B.n435 B.n434 10.6151
R1030 B.n434 B.n9 10.6151
R1031 B.n428 B.n9 10.6151
R1032 B.n428 B.n427 10.6151
R1033 B.n427 B.n426 10.6151
R1034 B.n426 B.n16 10.6151
R1035 B.n420 B.n16 10.6151
R1036 B.n420 B.n419 10.6151
R1037 B.n419 B.n418 10.6151
R1038 B.n418 B.n24 10.6151
R1039 B.n412 B.n24 10.6151
R1040 B.n412 B.n411 10.6151
R1041 B.n411 B.n410 10.6151
R1042 B.n109 B.n65 6.5566
R1043 B.n126 B.n125 6.5566
R1044 B.n268 B.n215 6.5566
R1045 B.n211 B.n210 6.5566
R1046 B.n106 B.n65 4.05904
R1047 B.n127 B.n126 4.05904
R1048 B.n269 B.n268 4.05904
R1049 B.n291 B.n210 4.05904
R1050 B.n442 B.n0 2.81026
R1051 B.n442 B.n1 2.81026
R1052 VP.n1 VP.t3 503.69
R1053 VP.n8 VP.t2 482.709
R1054 VP.n6 VP.t4 482.709
R1055 VP.n7 VP.t1 482.709
R1056 VP.n3 VP.t5 482.709
R1057 VP.n2 VP.t0 482.709
R1058 VP.n9 VP.n8 161.3
R1059 VP.n4 VP.n3 161.3
R1060 VP.n7 VP.n0 161.3
R1061 VP.n6 VP.n5 161.3
R1062 VP.n4 VP.n1 70.4033
R1063 VP.n7 VP.n6 48.2005
R1064 VP.n8 VP.n7 48.2005
R1065 VP.n3 VP.n2 48.2005
R1066 VP.n5 VP.n4 34.6331
R1067 VP.n2 VP.n1 20.9576
R1068 VP.n5 VP.n0 0.189894
R1069 VP.n9 VP.n0 0.189894
R1070 VP VP.n9 0.0516364
R1071 VDD1.n22 VDD1.n0 289.615
R1072 VDD1.n49 VDD1.n27 289.615
R1073 VDD1.n23 VDD1.n22 185
R1074 VDD1.n21 VDD1.n20 185
R1075 VDD1.n4 VDD1.n3 185
R1076 VDD1.n15 VDD1.n14 185
R1077 VDD1.n13 VDD1.n12 185
R1078 VDD1.n8 VDD1.n7 185
R1079 VDD1.n35 VDD1.n34 185
R1080 VDD1.n40 VDD1.n39 185
R1081 VDD1.n42 VDD1.n41 185
R1082 VDD1.n31 VDD1.n30 185
R1083 VDD1.n48 VDD1.n47 185
R1084 VDD1.n50 VDD1.n49 185
R1085 VDD1.n9 VDD1.t2 147.672
R1086 VDD1.n36 VDD1.t1 147.672
R1087 VDD1.n22 VDD1.n21 104.615
R1088 VDD1.n21 VDD1.n3 104.615
R1089 VDD1.n14 VDD1.n3 104.615
R1090 VDD1.n14 VDD1.n13 104.615
R1091 VDD1.n13 VDD1.n7 104.615
R1092 VDD1.n40 VDD1.n34 104.615
R1093 VDD1.n41 VDD1.n40 104.615
R1094 VDD1.n41 VDD1.n30 104.615
R1095 VDD1.n48 VDD1.n30 104.615
R1096 VDD1.n49 VDD1.n48 104.615
R1097 VDD1.n55 VDD1.n54 66.6108
R1098 VDD1.n57 VDD1.n56 66.5218
R1099 VDD1.t2 VDD1.n7 52.3082
R1100 VDD1.t1 VDD1.n34 52.3082
R1101 VDD1 VDD1.n26 47.2222
R1102 VDD1.n55 VDD1.n53 47.1086
R1103 VDD1.n57 VDD1.n55 30.9211
R1104 VDD1.n9 VDD1.n8 15.6666
R1105 VDD1.n36 VDD1.n35 15.6666
R1106 VDD1.n12 VDD1.n11 12.8005
R1107 VDD1.n39 VDD1.n38 12.8005
R1108 VDD1.n15 VDD1.n6 12.0247
R1109 VDD1.n42 VDD1.n33 12.0247
R1110 VDD1.n16 VDD1.n4 11.249
R1111 VDD1.n43 VDD1.n31 11.249
R1112 VDD1.n20 VDD1.n19 10.4732
R1113 VDD1.n47 VDD1.n46 10.4732
R1114 VDD1.n23 VDD1.n2 9.69747
R1115 VDD1.n50 VDD1.n29 9.69747
R1116 VDD1.n26 VDD1.n25 9.45567
R1117 VDD1.n53 VDD1.n52 9.45567
R1118 VDD1.n25 VDD1.n24 9.3005
R1119 VDD1.n2 VDD1.n1 9.3005
R1120 VDD1.n19 VDD1.n18 9.3005
R1121 VDD1.n17 VDD1.n16 9.3005
R1122 VDD1.n6 VDD1.n5 9.3005
R1123 VDD1.n11 VDD1.n10 9.3005
R1124 VDD1.n52 VDD1.n51 9.3005
R1125 VDD1.n29 VDD1.n28 9.3005
R1126 VDD1.n46 VDD1.n45 9.3005
R1127 VDD1.n44 VDD1.n43 9.3005
R1128 VDD1.n33 VDD1.n32 9.3005
R1129 VDD1.n38 VDD1.n37 9.3005
R1130 VDD1.n24 VDD1.n0 8.92171
R1131 VDD1.n51 VDD1.n27 8.92171
R1132 VDD1.n26 VDD1.n0 5.04292
R1133 VDD1.n53 VDD1.n27 5.04292
R1134 VDD1.n10 VDD1.n9 4.38687
R1135 VDD1.n37 VDD1.n36 4.38687
R1136 VDD1.n24 VDD1.n23 4.26717
R1137 VDD1.n51 VDD1.n50 4.26717
R1138 VDD1.n56 VDD1.t5 3.83029
R1139 VDD1.n56 VDD1.t0 3.83029
R1140 VDD1.n54 VDD1.t4 3.83029
R1141 VDD1.n54 VDD1.t3 3.83029
R1142 VDD1.n20 VDD1.n2 3.49141
R1143 VDD1.n47 VDD1.n29 3.49141
R1144 VDD1.n19 VDD1.n4 2.71565
R1145 VDD1.n46 VDD1.n31 2.71565
R1146 VDD1.n16 VDD1.n15 1.93989
R1147 VDD1.n43 VDD1.n42 1.93989
R1148 VDD1.n12 VDD1.n6 1.16414
R1149 VDD1.n39 VDD1.n33 1.16414
R1150 VDD1.n11 VDD1.n8 0.388379
R1151 VDD1.n38 VDD1.n35 0.388379
R1152 VDD1.n25 VDD1.n1 0.155672
R1153 VDD1.n18 VDD1.n1 0.155672
R1154 VDD1.n18 VDD1.n17 0.155672
R1155 VDD1.n17 VDD1.n5 0.155672
R1156 VDD1.n10 VDD1.n5 0.155672
R1157 VDD1.n37 VDD1.n32 0.155672
R1158 VDD1.n44 VDD1.n32 0.155672
R1159 VDD1.n45 VDD1.n44 0.155672
R1160 VDD1.n45 VDD1.n28 0.155672
R1161 VDD1.n52 VDD1.n28 0.155672
R1162 VDD1 VDD1.n57 0.0867069
C0 VTAIL VDD2 6.66663f
C1 VN VDD1 0.147694f
C2 VP VTAIL 1.33627f
C3 VN VDD2 1.43364f
C4 VN VP 3.46846f
C5 VDD2 VDD1 0.582072f
C6 VN VTAIL 1.32189f
C7 VP VDD1 1.54981f
C8 VTAIL VDD1 6.63186f
C9 VP VDD2 0.270126f
C10 VDD2 B 2.931709f
C11 VDD1 B 2.931263f
C12 VTAIL B 3.51318f
C13 VN B 5.183354f
C14 VP B 4.14345f
C15 VDD1.n0 B 0.027873f
C16 VDD1.n1 B 0.021369f
C17 VDD1.n2 B 0.011483f
C18 VDD1.n3 B 0.027141f
C19 VDD1.n4 B 0.012158f
C20 VDD1.n5 B 0.021369f
C21 VDD1.n6 B 0.011483f
C22 VDD1.n7 B 0.020356f
C23 VDD1.n8 B 0.016029f
C24 VDD1.t2 B 0.044239f
C25 VDD1.n9 B 0.087106f
C26 VDD1.n10 B 0.426998f
C27 VDD1.n11 B 0.011483f
C28 VDD1.n12 B 0.012158f
C29 VDD1.n13 B 0.027141f
C30 VDD1.n14 B 0.027141f
C31 VDD1.n15 B 0.012158f
C32 VDD1.n16 B 0.011483f
C33 VDD1.n17 B 0.021369f
C34 VDD1.n18 B 0.021369f
C35 VDD1.n19 B 0.011483f
C36 VDD1.n20 B 0.012158f
C37 VDD1.n21 B 0.027141f
C38 VDD1.n22 B 0.054931f
C39 VDD1.n23 B 0.012158f
C40 VDD1.n24 B 0.011483f
C41 VDD1.n25 B 0.046182f
C42 VDD1.n26 B 0.045785f
C43 VDD1.n27 B 0.027873f
C44 VDD1.n28 B 0.021369f
C45 VDD1.n29 B 0.011483f
C46 VDD1.n30 B 0.027141f
C47 VDD1.n31 B 0.012158f
C48 VDD1.n32 B 0.021369f
C49 VDD1.n33 B 0.011483f
C50 VDD1.n34 B 0.020356f
C51 VDD1.n35 B 0.016029f
C52 VDD1.t1 B 0.044239f
C53 VDD1.n36 B 0.087106f
C54 VDD1.n37 B 0.426998f
C55 VDD1.n38 B 0.011483f
C56 VDD1.n39 B 0.012158f
C57 VDD1.n40 B 0.027141f
C58 VDD1.n41 B 0.027141f
C59 VDD1.n42 B 0.012158f
C60 VDD1.n43 B 0.011483f
C61 VDD1.n44 B 0.021369f
C62 VDD1.n45 B 0.021369f
C63 VDD1.n46 B 0.011483f
C64 VDD1.n47 B 0.012158f
C65 VDD1.n48 B 0.027141f
C66 VDD1.n49 B 0.054931f
C67 VDD1.n50 B 0.012158f
C68 VDD1.n51 B 0.011483f
C69 VDD1.n52 B 0.046182f
C70 VDD1.n53 B 0.045558f
C71 VDD1.t4 B 0.087302f
C72 VDD1.t3 B 0.087302f
C73 VDD1.n54 B 0.714154f
C74 VDD1.n55 B 1.15578f
C75 VDD1.t5 B 0.087302f
C76 VDD1.t0 B 0.087302f
C77 VDD1.n56 B 0.713845f
C78 VDD1.n57 B 1.36863f
C79 VP.n0 B 0.031694f
C80 VP.t2 B 0.162574f
C81 VP.t3 B 0.166008f
C82 VP.n1 B 0.079176f
C83 VP.t5 B 0.162574f
C84 VP.t0 B 0.162574f
C85 VP.n2 B 0.088837f
C86 VP.n3 B 0.082389f
C87 VP.n4 B 0.991994f
C88 VP.n5 B 0.958206f
C89 VP.t4 B 0.162574f
C90 VP.n6 B 0.082389f
C91 VP.t1 B 0.162574f
C92 VP.n7 B 0.088837f
C93 VP.n8 B 0.082389f
C94 VP.n9 B 0.024562f
C95 VDD2.n0 B 0.028638f
C96 VDD2.n1 B 0.021955f
C97 VDD2.n2 B 0.011798f
C98 VDD2.n3 B 0.027886f
C99 VDD2.n4 B 0.012492f
C100 VDD2.n5 B 0.021955f
C101 VDD2.n6 B 0.011798f
C102 VDD2.n7 B 0.020914f
C103 VDD2.n8 B 0.016469f
C104 VDD2.t1 B 0.045453f
C105 VDD2.n9 B 0.089496f
C106 VDD2.n10 B 0.438714f
C107 VDD2.n11 B 0.011798f
C108 VDD2.n12 B 0.012492f
C109 VDD2.n13 B 0.027886f
C110 VDD2.n14 B 0.027886f
C111 VDD2.n15 B 0.012492f
C112 VDD2.n16 B 0.011798f
C113 VDD2.n17 B 0.021955f
C114 VDD2.n18 B 0.021955f
C115 VDD2.n19 B 0.011798f
C116 VDD2.n20 B 0.012492f
C117 VDD2.n21 B 0.027886f
C118 VDD2.n22 B 0.056439f
C119 VDD2.n23 B 0.012492f
C120 VDD2.n24 B 0.011798f
C121 VDD2.n25 B 0.047449f
C122 VDD2.n26 B 0.046808f
C123 VDD2.t3 B 0.089698f
C124 VDD2.t5 B 0.089698f
C125 VDD2.n27 B 0.733749f
C126 VDD2.n28 B 1.12875f
C127 VDD2.n29 B 0.028638f
C128 VDD2.n30 B 0.021955f
C129 VDD2.n31 B 0.011798f
C130 VDD2.n32 B 0.027886f
C131 VDD2.n33 B 0.012492f
C132 VDD2.n34 B 0.021955f
C133 VDD2.n35 B 0.011798f
C134 VDD2.n36 B 0.020914f
C135 VDD2.n37 B 0.016469f
C136 VDD2.t4 B 0.045453f
C137 VDD2.n38 B 0.089496f
C138 VDD2.n39 B 0.438714f
C139 VDD2.n40 B 0.011798f
C140 VDD2.n41 B 0.012492f
C141 VDD2.n42 B 0.027886f
C142 VDD2.n43 B 0.027886f
C143 VDD2.n44 B 0.012492f
C144 VDD2.n45 B 0.011798f
C145 VDD2.n46 B 0.021955f
C146 VDD2.n47 B 0.021955f
C147 VDD2.n48 B 0.011798f
C148 VDD2.n49 B 0.012492f
C149 VDD2.n50 B 0.027886f
C150 VDD2.n51 B 0.056439f
C151 VDD2.n52 B 0.012492f
C152 VDD2.n53 B 0.011798f
C153 VDD2.n54 B 0.047449f
C154 VDD2.n55 B 0.046259f
C155 VDD2.n56 B 1.22726f
C156 VDD2.t2 B 0.089698f
C157 VDD2.t0 B 0.089698f
C158 VDD2.n57 B 0.733731f
C159 VTAIL.t11 B 0.099639f
C160 VTAIL.t7 B 0.099639f
C161 VTAIL.n0 B 0.750872f
C162 VTAIL.n1 B 0.301648f
C163 VTAIL.n2 B 0.031812f
C164 VTAIL.n3 B 0.024388f
C165 VTAIL.n4 B 0.013105f
C166 VTAIL.n5 B 0.030976f
C167 VTAIL.n6 B 0.013876f
C168 VTAIL.n7 B 0.024388f
C169 VTAIL.n8 B 0.013105f
C170 VTAIL.n9 B 0.023232f
C171 VTAIL.n10 B 0.018294f
C172 VTAIL.t4 B 0.05049f
C173 VTAIL.n11 B 0.099414f
C174 VTAIL.n12 B 0.487334f
C175 VTAIL.n13 B 0.013105f
C176 VTAIL.n14 B 0.013876f
C177 VTAIL.n15 B 0.030976f
C178 VTAIL.n16 B 0.030976f
C179 VTAIL.n17 B 0.013876f
C180 VTAIL.n18 B 0.013105f
C181 VTAIL.n19 B 0.024388f
C182 VTAIL.n20 B 0.024388f
C183 VTAIL.n21 B 0.013105f
C184 VTAIL.n22 B 0.013876f
C185 VTAIL.n23 B 0.030976f
C186 VTAIL.n24 B 0.062693f
C187 VTAIL.n25 B 0.013876f
C188 VTAIL.n26 B 0.013105f
C189 VTAIL.n27 B 0.052708f
C190 VTAIL.n28 B 0.034514f
C191 VTAIL.n29 B 0.12377f
C192 VTAIL.t1 B 0.099639f
C193 VTAIL.t0 B 0.099639f
C194 VTAIL.n30 B 0.750872f
C195 VTAIL.n31 B 1.04381f
C196 VTAIL.t6 B 0.099639f
C197 VTAIL.t10 B 0.099639f
C198 VTAIL.n32 B 0.750878f
C199 VTAIL.n33 B 1.04381f
C200 VTAIL.n34 B 0.031812f
C201 VTAIL.n35 B 0.024388f
C202 VTAIL.n36 B 0.013105f
C203 VTAIL.n37 B 0.030976f
C204 VTAIL.n38 B 0.013876f
C205 VTAIL.n39 B 0.024388f
C206 VTAIL.n40 B 0.013105f
C207 VTAIL.n41 B 0.023232f
C208 VTAIL.n42 B 0.018294f
C209 VTAIL.t8 B 0.05049f
C210 VTAIL.n43 B 0.099414f
C211 VTAIL.n44 B 0.487334f
C212 VTAIL.n45 B 0.013105f
C213 VTAIL.n46 B 0.013876f
C214 VTAIL.n47 B 0.030976f
C215 VTAIL.n48 B 0.030976f
C216 VTAIL.n49 B 0.013876f
C217 VTAIL.n50 B 0.013105f
C218 VTAIL.n51 B 0.024388f
C219 VTAIL.n52 B 0.024388f
C220 VTAIL.n53 B 0.013105f
C221 VTAIL.n54 B 0.013876f
C222 VTAIL.n55 B 0.030976f
C223 VTAIL.n56 B 0.062693f
C224 VTAIL.n57 B 0.013876f
C225 VTAIL.n58 B 0.013105f
C226 VTAIL.n59 B 0.052708f
C227 VTAIL.n60 B 0.034514f
C228 VTAIL.n61 B 0.12377f
C229 VTAIL.t3 B 0.099639f
C230 VTAIL.t5 B 0.099639f
C231 VTAIL.n62 B 0.750878f
C232 VTAIL.n63 B 0.331112f
C233 VTAIL.n64 B 0.031812f
C234 VTAIL.n65 B 0.024388f
C235 VTAIL.n66 B 0.013105f
C236 VTAIL.n67 B 0.030976f
C237 VTAIL.n68 B 0.013876f
C238 VTAIL.n69 B 0.024388f
C239 VTAIL.n70 B 0.013105f
C240 VTAIL.n71 B 0.023232f
C241 VTAIL.n72 B 0.018294f
C242 VTAIL.t2 B 0.05049f
C243 VTAIL.n73 B 0.099414f
C244 VTAIL.n74 B 0.487334f
C245 VTAIL.n75 B 0.013105f
C246 VTAIL.n76 B 0.013876f
C247 VTAIL.n77 B 0.030976f
C248 VTAIL.n78 B 0.030976f
C249 VTAIL.n79 B 0.013876f
C250 VTAIL.n80 B 0.013105f
C251 VTAIL.n81 B 0.024388f
C252 VTAIL.n82 B 0.024388f
C253 VTAIL.n83 B 0.013105f
C254 VTAIL.n84 B 0.013876f
C255 VTAIL.n85 B 0.030976f
C256 VTAIL.n86 B 0.062693f
C257 VTAIL.n87 B 0.013876f
C258 VTAIL.n88 B 0.013105f
C259 VTAIL.n89 B 0.052708f
C260 VTAIL.n90 B 0.034514f
C261 VTAIL.n91 B 0.791076f
C262 VTAIL.n92 B 0.031812f
C263 VTAIL.n93 B 0.024388f
C264 VTAIL.n94 B 0.013105f
C265 VTAIL.n95 B 0.030976f
C266 VTAIL.n96 B 0.013876f
C267 VTAIL.n97 B 0.024388f
C268 VTAIL.n98 B 0.013105f
C269 VTAIL.n99 B 0.023232f
C270 VTAIL.n100 B 0.018294f
C271 VTAIL.t9 B 0.05049f
C272 VTAIL.n101 B 0.099414f
C273 VTAIL.n102 B 0.487334f
C274 VTAIL.n103 B 0.013105f
C275 VTAIL.n104 B 0.013876f
C276 VTAIL.n105 B 0.030976f
C277 VTAIL.n106 B 0.030976f
C278 VTAIL.n107 B 0.013876f
C279 VTAIL.n108 B 0.013105f
C280 VTAIL.n109 B 0.024388f
C281 VTAIL.n110 B 0.024388f
C282 VTAIL.n111 B 0.013105f
C283 VTAIL.n112 B 0.013876f
C284 VTAIL.n113 B 0.030976f
C285 VTAIL.n114 B 0.062693f
C286 VTAIL.n115 B 0.013876f
C287 VTAIL.n116 B 0.013105f
C288 VTAIL.n117 B 0.052708f
C289 VTAIL.n118 B 0.034514f
C290 VTAIL.n119 B 0.775156f
C291 VN.t4 B 0.163921f
C292 VN.n0 B 0.078181f
C293 VN.t0 B 0.16053f
C294 VN.t2 B 0.16053f
C295 VN.n1 B 0.087721f
C296 VN.n2 B 0.081353f
C297 VN.n3 B 0.090099f
C298 VN.t5 B 0.163921f
C299 VN.n4 B 0.078181f
C300 VN.t3 B 0.16053f
C301 VN.n5 B 0.087721f
C302 VN.t1 B 0.16053f
C303 VN.n6 B 0.081353f
C304 VN.n7 B 1.00034f
.ends

