* NGSPICE file created from diff_pair_sample_0337.ext - technology: sky130A

.subckt diff_pair_sample_0337 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=0 ps=0 w=6.54 l=1.96
X1 B.t8 B.t6 B.t7 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=0 ps=0 w=6.54 l=1.96
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=2.5506 ps=13.86 w=6.54 l=1.96
X3 B.t5 B.t3 B.t4 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=0 ps=0 w=6.54 l=1.96
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=2.5506 ps=13.86 w=6.54 l=1.96
X5 B.t2 B.t0 B.t1 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=0 ps=0 w=6.54 l=1.96
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=2.5506 ps=13.86 w=6.54 l=1.96
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1886_n2276# sky130_fd_pr__pfet_01v8 ad=2.5506 pd=13.86 as=2.5506 ps=13.86 w=6.54 l=1.96
R0 B.n237 B.n236 585
R1 B.n235 B.n70 585
R2 B.n234 B.n233 585
R3 B.n232 B.n71 585
R4 B.n231 B.n230 585
R5 B.n229 B.n72 585
R6 B.n228 B.n227 585
R7 B.n226 B.n73 585
R8 B.n225 B.n224 585
R9 B.n223 B.n74 585
R10 B.n222 B.n221 585
R11 B.n220 B.n75 585
R12 B.n219 B.n218 585
R13 B.n217 B.n76 585
R14 B.n216 B.n215 585
R15 B.n214 B.n77 585
R16 B.n213 B.n212 585
R17 B.n211 B.n78 585
R18 B.n210 B.n209 585
R19 B.n208 B.n79 585
R20 B.n207 B.n206 585
R21 B.n205 B.n80 585
R22 B.n204 B.n203 585
R23 B.n202 B.n81 585
R24 B.n201 B.n200 585
R25 B.n199 B.n82 585
R26 B.n198 B.n197 585
R27 B.n193 B.n83 585
R28 B.n192 B.n191 585
R29 B.n190 B.n84 585
R30 B.n189 B.n188 585
R31 B.n187 B.n85 585
R32 B.n186 B.n185 585
R33 B.n184 B.n86 585
R34 B.n183 B.n182 585
R35 B.n180 B.n87 585
R36 B.n179 B.n178 585
R37 B.n177 B.n90 585
R38 B.n176 B.n175 585
R39 B.n174 B.n91 585
R40 B.n173 B.n172 585
R41 B.n171 B.n92 585
R42 B.n170 B.n169 585
R43 B.n168 B.n93 585
R44 B.n167 B.n166 585
R45 B.n165 B.n94 585
R46 B.n164 B.n163 585
R47 B.n162 B.n95 585
R48 B.n161 B.n160 585
R49 B.n159 B.n96 585
R50 B.n158 B.n157 585
R51 B.n156 B.n97 585
R52 B.n155 B.n154 585
R53 B.n153 B.n98 585
R54 B.n152 B.n151 585
R55 B.n150 B.n99 585
R56 B.n149 B.n148 585
R57 B.n147 B.n100 585
R58 B.n146 B.n145 585
R59 B.n144 B.n101 585
R60 B.n143 B.n142 585
R61 B.n238 B.n69 585
R62 B.n240 B.n239 585
R63 B.n241 B.n68 585
R64 B.n243 B.n242 585
R65 B.n244 B.n67 585
R66 B.n246 B.n245 585
R67 B.n247 B.n66 585
R68 B.n249 B.n248 585
R69 B.n250 B.n65 585
R70 B.n252 B.n251 585
R71 B.n253 B.n64 585
R72 B.n255 B.n254 585
R73 B.n256 B.n63 585
R74 B.n258 B.n257 585
R75 B.n259 B.n62 585
R76 B.n261 B.n260 585
R77 B.n262 B.n61 585
R78 B.n264 B.n263 585
R79 B.n265 B.n60 585
R80 B.n267 B.n266 585
R81 B.n268 B.n59 585
R82 B.n270 B.n269 585
R83 B.n271 B.n58 585
R84 B.n273 B.n272 585
R85 B.n274 B.n57 585
R86 B.n276 B.n275 585
R87 B.n277 B.n56 585
R88 B.n279 B.n278 585
R89 B.n280 B.n55 585
R90 B.n282 B.n281 585
R91 B.n283 B.n54 585
R92 B.n285 B.n284 585
R93 B.n286 B.n53 585
R94 B.n288 B.n287 585
R95 B.n289 B.n52 585
R96 B.n291 B.n290 585
R97 B.n292 B.n51 585
R98 B.n294 B.n293 585
R99 B.n295 B.n50 585
R100 B.n297 B.n296 585
R101 B.n298 B.n49 585
R102 B.n300 B.n299 585
R103 B.n301 B.n48 585
R104 B.n303 B.n302 585
R105 B.n396 B.n395 585
R106 B.n394 B.n13 585
R107 B.n393 B.n392 585
R108 B.n391 B.n14 585
R109 B.n390 B.n389 585
R110 B.n388 B.n15 585
R111 B.n387 B.n386 585
R112 B.n385 B.n16 585
R113 B.n384 B.n383 585
R114 B.n382 B.n17 585
R115 B.n381 B.n380 585
R116 B.n379 B.n18 585
R117 B.n378 B.n377 585
R118 B.n376 B.n19 585
R119 B.n375 B.n374 585
R120 B.n373 B.n20 585
R121 B.n372 B.n371 585
R122 B.n370 B.n21 585
R123 B.n369 B.n368 585
R124 B.n367 B.n22 585
R125 B.n366 B.n365 585
R126 B.n364 B.n23 585
R127 B.n363 B.n362 585
R128 B.n361 B.n24 585
R129 B.n360 B.n359 585
R130 B.n358 B.n25 585
R131 B.n356 B.n355 585
R132 B.n354 B.n28 585
R133 B.n353 B.n352 585
R134 B.n351 B.n29 585
R135 B.n350 B.n349 585
R136 B.n348 B.n30 585
R137 B.n347 B.n346 585
R138 B.n345 B.n31 585
R139 B.n344 B.n343 585
R140 B.n342 B.n341 585
R141 B.n340 B.n35 585
R142 B.n339 B.n338 585
R143 B.n337 B.n36 585
R144 B.n336 B.n335 585
R145 B.n334 B.n37 585
R146 B.n333 B.n332 585
R147 B.n331 B.n38 585
R148 B.n330 B.n329 585
R149 B.n328 B.n39 585
R150 B.n327 B.n326 585
R151 B.n325 B.n40 585
R152 B.n324 B.n323 585
R153 B.n322 B.n41 585
R154 B.n321 B.n320 585
R155 B.n319 B.n42 585
R156 B.n318 B.n317 585
R157 B.n316 B.n43 585
R158 B.n315 B.n314 585
R159 B.n313 B.n44 585
R160 B.n312 B.n311 585
R161 B.n310 B.n45 585
R162 B.n309 B.n308 585
R163 B.n307 B.n46 585
R164 B.n306 B.n305 585
R165 B.n304 B.n47 585
R166 B.n397 B.n12 585
R167 B.n399 B.n398 585
R168 B.n400 B.n11 585
R169 B.n402 B.n401 585
R170 B.n403 B.n10 585
R171 B.n405 B.n404 585
R172 B.n406 B.n9 585
R173 B.n408 B.n407 585
R174 B.n409 B.n8 585
R175 B.n411 B.n410 585
R176 B.n412 B.n7 585
R177 B.n414 B.n413 585
R178 B.n415 B.n6 585
R179 B.n417 B.n416 585
R180 B.n418 B.n5 585
R181 B.n420 B.n419 585
R182 B.n421 B.n4 585
R183 B.n423 B.n422 585
R184 B.n424 B.n3 585
R185 B.n426 B.n425 585
R186 B.n427 B.n0 585
R187 B.n2 B.n1 585
R188 B.n113 B.n112 585
R189 B.n114 B.n111 585
R190 B.n116 B.n115 585
R191 B.n117 B.n110 585
R192 B.n119 B.n118 585
R193 B.n120 B.n109 585
R194 B.n122 B.n121 585
R195 B.n123 B.n108 585
R196 B.n125 B.n124 585
R197 B.n126 B.n107 585
R198 B.n128 B.n127 585
R199 B.n129 B.n106 585
R200 B.n131 B.n130 585
R201 B.n132 B.n105 585
R202 B.n134 B.n133 585
R203 B.n135 B.n104 585
R204 B.n137 B.n136 585
R205 B.n138 B.n103 585
R206 B.n140 B.n139 585
R207 B.n141 B.n102 585
R208 B.n142 B.n141 487.695
R209 B.n236 B.n69 487.695
R210 B.n302 B.n47 487.695
R211 B.n397 B.n396 487.695
R212 B.n194 B.t1 321.884
R213 B.n32 B.t11 321.884
R214 B.n88 B.t4 321.884
R215 B.n26 B.t8 321.884
R216 B.n88 B.t3 287.238
R217 B.n194 B.t0 287.238
R218 B.n32 B.t9 287.238
R219 B.n26 B.t6 287.238
R220 B.n195 B.t2 277.471
R221 B.n33 B.t10 277.471
R222 B.n89 B.t5 277.471
R223 B.n27 B.t7 277.471
R224 B.n429 B.n428 256.663
R225 B.n428 B.n427 235.042
R226 B.n428 B.n2 235.042
R227 B.n142 B.n101 163.367
R228 B.n146 B.n101 163.367
R229 B.n147 B.n146 163.367
R230 B.n148 B.n147 163.367
R231 B.n148 B.n99 163.367
R232 B.n152 B.n99 163.367
R233 B.n153 B.n152 163.367
R234 B.n154 B.n153 163.367
R235 B.n154 B.n97 163.367
R236 B.n158 B.n97 163.367
R237 B.n159 B.n158 163.367
R238 B.n160 B.n159 163.367
R239 B.n160 B.n95 163.367
R240 B.n164 B.n95 163.367
R241 B.n165 B.n164 163.367
R242 B.n166 B.n165 163.367
R243 B.n166 B.n93 163.367
R244 B.n170 B.n93 163.367
R245 B.n171 B.n170 163.367
R246 B.n172 B.n171 163.367
R247 B.n172 B.n91 163.367
R248 B.n176 B.n91 163.367
R249 B.n177 B.n176 163.367
R250 B.n178 B.n177 163.367
R251 B.n178 B.n87 163.367
R252 B.n183 B.n87 163.367
R253 B.n184 B.n183 163.367
R254 B.n185 B.n184 163.367
R255 B.n185 B.n85 163.367
R256 B.n189 B.n85 163.367
R257 B.n190 B.n189 163.367
R258 B.n191 B.n190 163.367
R259 B.n191 B.n83 163.367
R260 B.n198 B.n83 163.367
R261 B.n199 B.n198 163.367
R262 B.n200 B.n199 163.367
R263 B.n200 B.n81 163.367
R264 B.n204 B.n81 163.367
R265 B.n205 B.n204 163.367
R266 B.n206 B.n205 163.367
R267 B.n206 B.n79 163.367
R268 B.n210 B.n79 163.367
R269 B.n211 B.n210 163.367
R270 B.n212 B.n211 163.367
R271 B.n212 B.n77 163.367
R272 B.n216 B.n77 163.367
R273 B.n217 B.n216 163.367
R274 B.n218 B.n217 163.367
R275 B.n218 B.n75 163.367
R276 B.n222 B.n75 163.367
R277 B.n223 B.n222 163.367
R278 B.n224 B.n223 163.367
R279 B.n224 B.n73 163.367
R280 B.n228 B.n73 163.367
R281 B.n229 B.n228 163.367
R282 B.n230 B.n229 163.367
R283 B.n230 B.n71 163.367
R284 B.n234 B.n71 163.367
R285 B.n235 B.n234 163.367
R286 B.n236 B.n235 163.367
R287 B.n302 B.n301 163.367
R288 B.n301 B.n300 163.367
R289 B.n300 B.n49 163.367
R290 B.n296 B.n49 163.367
R291 B.n296 B.n295 163.367
R292 B.n295 B.n294 163.367
R293 B.n294 B.n51 163.367
R294 B.n290 B.n51 163.367
R295 B.n290 B.n289 163.367
R296 B.n289 B.n288 163.367
R297 B.n288 B.n53 163.367
R298 B.n284 B.n53 163.367
R299 B.n284 B.n283 163.367
R300 B.n283 B.n282 163.367
R301 B.n282 B.n55 163.367
R302 B.n278 B.n55 163.367
R303 B.n278 B.n277 163.367
R304 B.n277 B.n276 163.367
R305 B.n276 B.n57 163.367
R306 B.n272 B.n57 163.367
R307 B.n272 B.n271 163.367
R308 B.n271 B.n270 163.367
R309 B.n270 B.n59 163.367
R310 B.n266 B.n59 163.367
R311 B.n266 B.n265 163.367
R312 B.n265 B.n264 163.367
R313 B.n264 B.n61 163.367
R314 B.n260 B.n61 163.367
R315 B.n260 B.n259 163.367
R316 B.n259 B.n258 163.367
R317 B.n258 B.n63 163.367
R318 B.n254 B.n63 163.367
R319 B.n254 B.n253 163.367
R320 B.n253 B.n252 163.367
R321 B.n252 B.n65 163.367
R322 B.n248 B.n65 163.367
R323 B.n248 B.n247 163.367
R324 B.n247 B.n246 163.367
R325 B.n246 B.n67 163.367
R326 B.n242 B.n67 163.367
R327 B.n242 B.n241 163.367
R328 B.n241 B.n240 163.367
R329 B.n240 B.n69 163.367
R330 B.n396 B.n13 163.367
R331 B.n392 B.n13 163.367
R332 B.n392 B.n391 163.367
R333 B.n391 B.n390 163.367
R334 B.n390 B.n15 163.367
R335 B.n386 B.n15 163.367
R336 B.n386 B.n385 163.367
R337 B.n385 B.n384 163.367
R338 B.n384 B.n17 163.367
R339 B.n380 B.n17 163.367
R340 B.n380 B.n379 163.367
R341 B.n379 B.n378 163.367
R342 B.n378 B.n19 163.367
R343 B.n374 B.n19 163.367
R344 B.n374 B.n373 163.367
R345 B.n373 B.n372 163.367
R346 B.n372 B.n21 163.367
R347 B.n368 B.n21 163.367
R348 B.n368 B.n367 163.367
R349 B.n367 B.n366 163.367
R350 B.n366 B.n23 163.367
R351 B.n362 B.n23 163.367
R352 B.n362 B.n361 163.367
R353 B.n361 B.n360 163.367
R354 B.n360 B.n25 163.367
R355 B.n355 B.n25 163.367
R356 B.n355 B.n354 163.367
R357 B.n354 B.n353 163.367
R358 B.n353 B.n29 163.367
R359 B.n349 B.n29 163.367
R360 B.n349 B.n348 163.367
R361 B.n348 B.n347 163.367
R362 B.n347 B.n31 163.367
R363 B.n343 B.n31 163.367
R364 B.n343 B.n342 163.367
R365 B.n342 B.n35 163.367
R366 B.n338 B.n35 163.367
R367 B.n338 B.n337 163.367
R368 B.n337 B.n336 163.367
R369 B.n336 B.n37 163.367
R370 B.n332 B.n37 163.367
R371 B.n332 B.n331 163.367
R372 B.n331 B.n330 163.367
R373 B.n330 B.n39 163.367
R374 B.n326 B.n39 163.367
R375 B.n326 B.n325 163.367
R376 B.n325 B.n324 163.367
R377 B.n324 B.n41 163.367
R378 B.n320 B.n41 163.367
R379 B.n320 B.n319 163.367
R380 B.n319 B.n318 163.367
R381 B.n318 B.n43 163.367
R382 B.n314 B.n43 163.367
R383 B.n314 B.n313 163.367
R384 B.n313 B.n312 163.367
R385 B.n312 B.n45 163.367
R386 B.n308 B.n45 163.367
R387 B.n308 B.n307 163.367
R388 B.n307 B.n306 163.367
R389 B.n306 B.n47 163.367
R390 B.n398 B.n397 163.367
R391 B.n398 B.n11 163.367
R392 B.n402 B.n11 163.367
R393 B.n403 B.n402 163.367
R394 B.n404 B.n403 163.367
R395 B.n404 B.n9 163.367
R396 B.n408 B.n9 163.367
R397 B.n409 B.n408 163.367
R398 B.n410 B.n409 163.367
R399 B.n410 B.n7 163.367
R400 B.n414 B.n7 163.367
R401 B.n415 B.n414 163.367
R402 B.n416 B.n415 163.367
R403 B.n416 B.n5 163.367
R404 B.n420 B.n5 163.367
R405 B.n421 B.n420 163.367
R406 B.n422 B.n421 163.367
R407 B.n422 B.n3 163.367
R408 B.n426 B.n3 163.367
R409 B.n427 B.n426 163.367
R410 B.n112 B.n2 163.367
R411 B.n112 B.n111 163.367
R412 B.n116 B.n111 163.367
R413 B.n117 B.n116 163.367
R414 B.n118 B.n117 163.367
R415 B.n118 B.n109 163.367
R416 B.n122 B.n109 163.367
R417 B.n123 B.n122 163.367
R418 B.n124 B.n123 163.367
R419 B.n124 B.n107 163.367
R420 B.n128 B.n107 163.367
R421 B.n129 B.n128 163.367
R422 B.n130 B.n129 163.367
R423 B.n130 B.n105 163.367
R424 B.n134 B.n105 163.367
R425 B.n135 B.n134 163.367
R426 B.n136 B.n135 163.367
R427 B.n136 B.n103 163.367
R428 B.n140 B.n103 163.367
R429 B.n141 B.n140 163.367
R430 B.n181 B.n89 59.5399
R431 B.n196 B.n195 59.5399
R432 B.n34 B.n33 59.5399
R433 B.n357 B.n27 59.5399
R434 B.n89 B.n88 44.4126
R435 B.n195 B.n194 44.4126
R436 B.n33 B.n32 44.4126
R437 B.n27 B.n26 44.4126
R438 B.n395 B.n12 31.6883
R439 B.n304 B.n303 31.6883
R440 B.n238 B.n237 31.6883
R441 B.n143 B.n102 31.6883
R442 B B.n429 18.0485
R443 B.n399 B.n12 10.6151
R444 B.n400 B.n399 10.6151
R445 B.n401 B.n400 10.6151
R446 B.n401 B.n10 10.6151
R447 B.n405 B.n10 10.6151
R448 B.n406 B.n405 10.6151
R449 B.n407 B.n406 10.6151
R450 B.n407 B.n8 10.6151
R451 B.n411 B.n8 10.6151
R452 B.n412 B.n411 10.6151
R453 B.n413 B.n412 10.6151
R454 B.n413 B.n6 10.6151
R455 B.n417 B.n6 10.6151
R456 B.n418 B.n417 10.6151
R457 B.n419 B.n418 10.6151
R458 B.n419 B.n4 10.6151
R459 B.n423 B.n4 10.6151
R460 B.n424 B.n423 10.6151
R461 B.n425 B.n424 10.6151
R462 B.n425 B.n0 10.6151
R463 B.n395 B.n394 10.6151
R464 B.n394 B.n393 10.6151
R465 B.n393 B.n14 10.6151
R466 B.n389 B.n14 10.6151
R467 B.n389 B.n388 10.6151
R468 B.n388 B.n387 10.6151
R469 B.n387 B.n16 10.6151
R470 B.n383 B.n16 10.6151
R471 B.n383 B.n382 10.6151
R472 B.n382 B.n381 10.6151
R473 B.n381 B.n18 10.6151
R474 B.n377 B.n18 10.6151
R475 B.n377 B.n376 10.6151
R476 B.n376 B.n375 10.6151
R477 B.n375 B.n20 10.6151
R478 B.n371 B.n20 10.6151
R479 B.n371 B.n370 10.6151
R480 B.n370 B.n369 10.6151
R481 B.n369 B.n22 10.6151
R482 B.n365 B.n22 10.6151
R483 B.n365 B.n364 10.6151
R484 B.n364 B.n363 10.6151
R485 B.n363 B.n24 10.6151
R486 B.n359 B.n24 10.6151
R487 B.n359 B.n358 10.6151
R488 B.n356 B.n28 10.6151
R489 B.n352 B.n28 10.6151
R490 B.n352 B.n351 10.6151
R491 B.n351 B.n350 10.6151
R492 B.n350 B.n30 10.6151
R493 B.n346 B.n30 10.6151
R494 B.n346 B.n345 10.6151
R495 B.n345 B.n344 10.6151
R496 B.n341 B.n340 10.6151
R497 B.n340 B.n339 10.6151
R498 B.n339 B.n36 10.6151
R499 B.n335 B.n36 10.6151
R500 B.n335 B.n334 10.6151
R501 B.n334 B.n333 10.6151
R502 B.n333 B.n38 10.6151
R503 B.n329 B.n38 10.6151
R504 B.n329 B.n328 10.6151
R505 B.n328 B.n327 10.6151
R506 B.n327 B.n40 10.6151
R507 B.n323 B.n40 10.6151
R508 B.n323 B.n322 10.6151
R509 B.n322 B.n321 10.6151
R510 B.n321 B.n42 10.6151
R511 B.n317 B.n42 10.6151
R512 B.n317 B.n316 10.6151
R513 B.n316 B.n315 10.6151
R514 B.n315 B.n44 10.6151
R515 B.n311 B.n44 10.6151
R516 B.n311 B.n310 10.6151
R517 B.n310 B.n309 10.6151
R518 B.n309 B.n46 10.6151
R519 B.n305 B.n46 10.6151
R520 B.n305 B.n304 10.6151
R521 B.n303 B.n48 10.6151
R522 B.n299 B.n48 10.6151
R523 B.n299 B.n298 10.6151
R524 B.n298 B.n297 10.6151
R525 B.n297 B.n50 10.6151
R526 B.n293 B.n50 10.6151
R527 B.n293 B.n292 10.6151
R528 B.n292 B.n291 10.6151
R529 B.n291 B.n52 10.6151
R530 B.n287 B.n52 10.6151
R531 B.n287 B.n286 10.6151
R532 B.n286 B.n285 10.6151
R533 B.n285 B.n54 10.6151
R534 B.n281 B.n54 10.6151
R535 B.n281 B.n280 10.6151
R536 B.n280 B.n279 10.6151
R537 B.n279 B.n56 10.6151
R538 B.n275 B.n56 10.6151
R539 B.n275 B.n274 10.6151
R540 B.n274 B.n273 10.6151
R541 B.n273 B.n58 10.6151
R542 B.n269 B.n58 10.6151
R543 B.n269 B.n268 10.6151
R544 B.n268 B.n267 10.6151
R545 B.n267 B.n60 10.6151
R546 B.n263 B.n60 10.6151
R547 B.n263 B.n262 10.6151
R548 B.n262 B.n261 10.6151
R549 B.n261 B.n62 10.6151
R550 B.n257 B.n62 10.6151
R551 B.n257 B.n256 10.6151
R552 B.n256 B.n255 10.6151
R553 B.n255 B.n64 10.6151
R554 B.n251 B.n64 10.6151
R555 B.n251 B.n250 10.6151
R556 B.n250 B.n249 10.6151
R557 B.n249 B.n66 10.6151
R558 B.n245 B.n66 10.6151
R559 B.n245 B.n244 10.6151
R560 B.n244 B.n243 10.6151
R561 B.n243 B.n68 10.6151
R562 B.n239 B.n68 10.6151
R563 B.n239 B.n238 10.6151
R564 B.n113 B.n1 10.6151
R565 B.n114 B.n113 10.6151
R566 B.n115 B.n114 10.6151
R567 B.n115 B.n110 10.6151
R568 B.n119 B.n110 10.6151
R569 B.n120 B.n119 10.6151
R570 B.n121 B.n120 10.6151
R571 B.n121 B.n108 10.6151
R572 B.n125 B.n108 10.6151
R573 B.n126 B.n125 10.6151
R574 B.n127 B.n126 10.6151
R575 B.n127 B.n106 10.6151
R576 B.n131 B.n106 10.6151
R577 B.n132 B.n131 10.6151
R578 B.n133 B.n132 10.6151
R579 B.n133 B.n104 10.6151
R580 B.n137 B.n104 10.6151
R581 B.n138 B.n137 10.6151
R582 B.n139 B.n138 10.6151
R583 B.n139 B.n102 10.6151
R584 B.n144 B.n143 10.6151
R585 B.n145 B.n144 10.6151
R586 B.n145 B.n100 10.6151
R587 B.n149 B.n100 10.6151
R588 B.n150 B.n149 10.6151
R589 B.n151 B.n150 10.6151
R590 B.n151 B.n98 10.6151
R591 B.n155 B.n98 10.6151
R592 B.n156 B.n155 10.6151
R593 B.n157 B.n156 10.6151
R594 B.n157 B.n96 10.6151
R595 B.n161 B.n96 10.6151
R596 B.n162 B.n161 10.6151
R597 B.n163 B.n162 10.6151
R598 B.n163 B.n94 10.6151
R599 B.n167 B.n94 10.6151
R600 B.n168 B.n167 10.6151
R601 B.n169 B.n168 10.6151
R602 B.n169 B.n92 10.6151
R603 B.n173 B.n92 10.6151
R604 B.n174 B.n173 10.6151
R605 B.n175 B.n174 10.6151
R606 B.n175 B.n90 10.6151
R607 B.n179 B.n90 10.6151
R608 B.n180 B.n179 10.6151
R609 B.n182 B.n86 10.6151
R610 B.n186 B.n86 10.6151
R611 B.n187 B.n186 10.6151
R612 B.n188 B.n187 10.6151
R613 B.n188 B.n84 10.6151
R614 B.n192 B.n84 10.6151
R615 B.n193 B.n192 10.6151
R616 B.n197 B.n193 10.6151
R617 B.n201 B.n82 10.6151
R618 B.n202 B.n201 10.6151
R619 B.n203 B.n202 10.6151
R620 B.n203 B.n80 10.6151
R621 B.n207 B.n80 10.6151
R622 B.n208 B.n207 10.6151
R623 B.n209 B.n208 10.6151
R624 B.n209 B.n78 10.6151
R625 B.n213 B.n78 10.6151
R626 B.n214 B.n213 10.6151
R627 B.n215 B.n214 10.6151
R628 B.n215 B.n76 10.6151
R629 B.n219 B.n76 10.6151
R630 B.n220 B.n219 10.6151
R631 B.n221 B.n220 10.6151
R632 B.n221 B.n74 10.6151
R633 B.n225 B.n74 10.6151
R634 B.n226 B.n225 10.6151
R635 B.n227 B.n226 10.6151
R636 B.n227 B.n72 10.6151
R637 B.n231 B.n72 10.6151
R638 B.n232 B.n231 10.6151
R639 B.n233 B.n232 10.6151
R640 B.n233 B.n70 10.6151
R641 B.n237 B.n70 10.6151
R642 B.n429 B.n0 8.11757
R643 B.n429 B.n1 8.11757
R644 B.n357 B.n356 6.5566
R645 B.n344 B.n34 6.5566
R646 B.n182 B.n181 6.5566
R647 B.n197 B.n196 6.5566
R648 B.n358 B.n357 4.05904
R649 B.n341 B.n34 4.05904
R650 B.n181 B.n180 4.05904
R651 B.n196 B.n82 4.05904
R652 VN VN.t1 178.315
R653 VN VN.t0 139.542
R654 VTAIL.n134 VTAIL.n133 756.745
R655 VTAIL.n32 VTAIL.n31 756.745
R656 VTAIL.n100 VTAIL.n99 756.745
R657 VTAIL.n66 VTAIL.n65 756.745
R658 VTAIL.n112 VTAIL.n111 585
R659 VTAIL.n117 VTAIL.n116 585
R660 VTAIL.n119 VTAIL.n118 585
R661 VTAIL.n108 VTAIL.n107 585
R662 VTAIL.n125 VTAIL.n124 585
R663 VTAIL.n127 VTAIL.n126 585
R664 VTAIL.n104 VTAIL.n103 585
R665 VTAIL.n133 VTAIL.n132 585
R666 VTAIL.n10 VTAIL.n9 585
R667 VTAIL.n15 VTAIL.n14 585
R668 VTAIL.n17 VTAIL.n16 585
R669 VTAIL.n6 VTAIL.n5 585
R670 VTAIL.n23 VTAIL.n22 585
R671 VTAIL.n25 VTAIL.n24 585
R672 VTAIL.n2 VTAIL.n1 585
R673 VTAIL.n31 VTAIL.n30 585
R674 VTAIL.n99 VTAIL.n98 585
R675 VTAIL.n70 VTAIL.n69 585
R676 VTAIL.n93 VTAIL.n92 585
R677 VTAIL.n91 VTAIL.n90 585
R678 VTAIL.n74 VTAIL.n73 585
R679 VTAIL.n85 VTAIL.n84 585
R680 VTAIL.n83 VTAIL.n82 585
R681 VTAIL.n78 VTAIL.n77 585
R682 VTAIL.n65 VTAIL.n64 585
R683 VTAIL.n36 VTAIL.n35 585
R684 VTAIL.n59 VTAIL.n58 585
R685 VTAIL.n57 VTAIL.n56 585
R686 VTAIL.n40 VTAIL.n39 585
R687 VTAIL.n51 VTAIL.n50 585
R688 VTAIL.n49 VTAIL.n48 585
R689 VTAIL.n44 VTAIL.n43 585
R690 VTAIL.n113 VTAIL.t3 329.084
R691 VTAIL.n11 VTAIL.t0 329.084
R692 VTAIL.n79 VTAIL.t1 329.084
R693 VTAIL.n45 VTAIL.t2 329.084
R694 VTAIL.n117 VTAIL.n111 171.744
R695 VTAIL.n118 VTAIL.n117 171.744
R696 VTAIL.n118 VTAIL.n107 171.744
R697 VTAIL.n125 VTAIL.n107 171.744
R698 VTAIL.n126 VTAIL.n125 171.744
R699 VTAIL.n126 VTAIL.n103 171.744
R700 VTAIL.n133 VTAIL.n103 171.744
R701 VTAIL.n15 VTAIL.n9 171.744
R702 VTAIL.n16 VTAIL.n15 171.744
R703 VTAIL.n16 VTAIL.n5 171.744
R704 VTAIL.n23 VTAIL.n5 171.744
R705 VTAIL.n24 VTAIL.n23 171.744
R706 VTAIL.n24 VTAIL.n1 171.744
R707 VTAIL.n31 VTAIL.n1 171.744
R708 VTAIL.n99 VTAIL.n69 171.744
R709 VTAIL.n92 VTAIL.n69 171.744
R710 VTAIL.n92 VTAIL.n91 171.744
R711 VTAIL.n91 VTAIL.n73 171.744
R712 VTAIL.n84 VTAIL.n73 171.744
R713 VTAIL.n84 VTAIL.n83 171.744
R714 VTAIL.n83 VTAIL.n77 171.744
R715 VTAIL.n65 VTAIL.n35 171.744
R716 VTAIL.n58 VTAIL.n35 171.744
R717 VTAIL.n58 VTAIL.n57 171.744
R718 VTAIL.n57 VTAIL.n39 171.744
R719 VTAIL.n50 VTAIL.n39 171.744
R720 VTAIL.n50 VTAIL.n49 171.744
R721 VTAIL.n49 VTAIL.n43 171.744
R722 VTAIL.t3 VTAIL.n111 85.8723
R723 VTAIL.t0 VTAIL.n9 85.8723
R724 VTAIL.t1 VTAIL.n77 85.8723
R725 VTAIL.t2 VTAIL.n43 85.8723
R726 VTAIL.n135 VTAIL.n134 35.2884
R727 VTAIL.n33 VTAIL.n32 35.2884
R728 VTAIL.n101 VTAIL.n100 35.2884
R729 VTAIL.n67 VTAIL.n66 35.2884
R730 VTAIL.n67 VTAIL.n33 21.9531
R731 VTAIL.n135 VTAIL.n101 19.9789
R732 VTAIL.n132 VTAIL.n102 12.8005
R733 VTAIL.n30 VTAIL.n0 12.8005
R734 VTAIL.n98 VTAIL.n68 12.8005
R735 VTAIL.n64 VTAIL.n34 12.8005
R736 VTAIL.n131 VTAIL.n104 12.0247
R737 VTAIL.n29 VTAIL.n2 12.0247
R738 VTAIL.n97 VTAIL.n70 12.0247
R739 VTAIL.n63 VTAIL.n36 12.0247
R740 VTAIL.n128 VTAIL.n127 11.249
R741 VTAIL.n26 VTAIL.n25 11.249
R742 VTAIL.n94 VTAIL.n93 11.249
R743 VTAIL.n60 VTAIL.n59 11.249
R744 VTAIL.n113 VTAIL.n112 10.7233
R745 VTAIL.n11 VTAIL.n10 10.7233
R746 VTAIL.n79 VTAIL.n78 10.7233
R747 VTAIL.n45 VTAIL.n44 10.7233
R748 VTAIL.n124 VTAIL.n106 10.4732
R749 VTAIL.n22 VTAIL.n4 10.4732
R750 VTAIL.n90 VTAIL.n72 10.4732
R751 VTAIL.n56 VTAIL.n38 10.4732
R752 VTAIL.n123 VTAIL.n108 9.69747
R753 VTAIL.n21 VTAIL.n6 9.69747
R754 VTAIL.n89 VTAIL.n74 9.69747
R755 VTAIL.n55 VTAIL.n40 9.69747
R756 VTAIL.n130 VTAIL.n102 9.45567
R757 VTAIL.n28 VTAIL.n0 9.45567
R758 VTAIL.n96 VTAIL.n68 9.45567
R759 VTAIL.n62 VTAIL.n34 9.45567
R760 VTAIL.n115 VTAIL.n114 9.3005
R761 VTAIL.n110 VTAIL.n109 9.3005
R762 VTAIL.n121 VTAIL.n120 9.3005
R763 VTAIL.n123 VTAIL.n122 9.3005
R764 VTAIL.n106 VTAIL.n105 9.3005
R765 VTAIL.n129 VTAIL.n128 9.3005
R766 VTAIL.n131 VTAIL.n130 9.3005
R767 VTAIL.n13 VTAIL.n12 9.3005
R768 VTAIL.n8 VTAIL.n7 9.3005
R769 VTAIL.n19 VTAIL.n18 9.3005
R770 VTAIL.n21 VTAIL.n20 9.3005
R771 VTAIL.n4 VTAIL.n3 9.3005
R772 VTAIL.n27 VTAIL.n26 9.3005
R773 VTAIL.n29 VTAIL.n28 9.3005
R774 VTAIL.n97 VTAIL.n96 9.3005
R775 VTAIL.n95 VTAIL.n94 9.3005
R776 VTAIL.n72 VTAIL.n71 9.3005
R777 VTAIL.n89 VTAIL.n88 9.3005
R778 VTAIL.n87 VTAIL.n86 9.3005
R779 VTAIL.n76 VTAIL.n75 9.3005
R780 VTAIL.n81 VTAIL.n80 9.3005
R781 VTAIL.n42 VTAIL.n41 9.3005
R782 VTAIL.n53 VTAIL.n52 9.3005
R783 VTAIL.n55 VTAIL.n54 9.3005
R784 VTAIL.n38 VTAIL.n37 9.3005
R785 VTAIL.n61 VTAIL.n60 9.3005
R786 VTAIL.n63 VTAIL.n62 9.3005
R787 VTAIL.n47 VTAIL.n46 9.3005
R788 VTAIL.n120 VTAIL.n119 8.92171
R789 VTAIL.n18 VTAIL.n17 8.92171
R790 VTAIL.n86 VTAIL.n85 8.92171
R791 VTAIL.n52 VTAIL.n51 8.92171
R792 VTAIL.n116 VTAIL.n110 8.14595
R793 VTAIL.n14 VTAIL.n8 8.14595
R794 VTAIL.n82 VTAIL.n76 8.14595
R795 VTAIL.n48 VTAIL.n42 8.14595
R796 VTAIL.n115 VTAIL.n112 7.3702
R797 VTAIL.n13 VTAIL.n10 7.3702
R798 VTAIL.n81 VTAIL.n78 7.3702
R799 VTAIL.n47 VTAIL.n44 7.3702
R800 VTAIL.n116 VTAIL.n115 5.81868
R801 VTAIL.n14 VTAIL.n13 5.81868
R802 VTAIL.n82 VTAIL.n81 5.81868
R803 VTAIL.n48 VTAIL.n47 5.81868
R804 VTAIL.n119 VTAIL.n110 5.04292
R805 VTAIL.n17 VTAIL.n8 5.04292
R806 VTAIL.n85 VTAIL.n76 5.04292
R807 VTAIL.n51 VTAIL.n42 5.04292
R808 VTAIL.n120 VTAIL.n108 4.26717
R809 VTAIL.n18 VTAIL.n6 4.26717
R810 VTAIL.n86 VTAIL.n74 4.26717
R811 VTAIL.n52 VTAIL.n40 4.26717
R812 VTAIL.n124 VTAIL.n123 3.49141
R813 VTAIL.n22 VTAIL.n21 3.49141
R814 VTAIL.n90 VTAIL.n89 3.49141
R815 VTAIL.n56 VTAIL.n55 3.49141
R816 VTAIL.n127 VTAIL.n106 2.71565
R817 VTAIL.n25 VTAIL.n4 2.71565
R818 VTAIL.n93 VTAIL.n72 2.71565
R819 VTAIL.n59 VTAIL.n38 2.71565
R820 VTAIL.n46 VTAIL.n45 2.41347
R821 VTAIL.n114 VTAIL.n113 2.41347
R822 VTAIL.n12 VTAIL.n11 2.41347
R823 VTAIL.n80 VTAIL.n79 2.41347
R824 VTAIL.n128 VTAIL.n104 1.93989
R825 VTAIL.n26 VTAIL.n2 1.93989
R826 VTAIL.n94 VTAIL.n70 1.93989
R827 VTAIL.n60 VTAIL.n36 1.93989
R828 VTAIL.n101 VTAIL.n67 1.4574
R829 VTAIL.n132 VTAIL.n131 1.16414
R830 VTAIL.n30 VTAIL.n29 1.16414
R831 VTAIL.n98 VTAIL.n97 1.16414
R832 VTAIL.n64 VTAIL.n63 1.16414
R833 VTAIL VTAIL.n33 1.02205
R834 VTAIL VTAIL.n135 0.435845
R835 VTAIL.n134 VTAIL.n102 0.388379
R836 VTAIL.n32 VTAIL.n0 0.388379
R837 VTAIL.n100 VTAIL.n68 0.388379
R838 VTAIL.n66 VTAIL.n34 0.388379
R839 VTAIL.n114 VTAIL.n109 0.155672
R840 VTAIL.n121 VTAIL.n109 0.155672
R841 VTAIL.n122 VTAIL.n121 0.155672
R842 VTAIL.n122 VTAIL.n105 0.155672
R843 VTAIL.n129 VTAIL.n105 0.155672
R844 VTAIL.n130 VTAIL.n129 0.155672
R845 VTAIL.n12 VTAIL.n7 0.155672
R846 VTAIL.n19 VTAIL.n7 0.155672
R847 VTAIL.n20 VTAIL.n19 0.155672
R848 VTAIL.n20 VTAIL.n3 0.155672
R849 VTAIL.n27 VTAIL.n3 0.155672
R850 VTAIL.n28 VTAIL.n27 0.155672
R851 VTAIL.n96 VTAIL.n95 0.155672
R852 VTAIL.n95 VTAIL.n71 0.155672
R853 VTAIL.n88 VTAIL.n71 0.155672
R854 VTAIL.n88 VTAIL.n87 0.155672
R855 VTAIL.n87 VTAIL.n75 0.155672
R856 VTAIL.n80 VTAIL.n75 0.155672
R857 VTAIL.n62 VTAIL.n61 0.155672
R858 VTAIL.n61 VTAIL.n37 0.155672
R859 VTAIL.n54 VTAIL.n37 0.155672
R860 VTAIL.n54 VTAIL.n53 0.155672
R861 VTAIL.n53 VTAIL.n41 0.155672
R862 VTAIL.n46 VTAIL.n41 0.155672
R863 VDD2.n65 VDD2.n64 756.745
R864 VDD2.n32 VDD2.n31 756.745
R865 VDD2.n64 VDD2.n63 585
R866 VDD2.n35 VDD2.n34 585
R867 VDD2.n58 VDD2.n57 585
R868 VDD2.n56 VDD2.n55 585
R869 VDD2.n39 VDD2.n38 585
R870 VDD2.n50 VDD2.n49 585
R871 VDD2.n48 VDD2.n47 585
R872 VDD2.n43 VDD2.n42 585
R873 VDD2.n10 VDD2.n9 585
R874 VDD2.n15 VDD2.n14 585
R875 VDD2.n17 VDD2.n16 585
R876 VDD2.n6 VDD2.n5 585
R877 VDD2.n23 VDD2.n22 585
R878 VDD2.n25 VDD2.n24 585
R879 VDD2.n2 VDD2.n1 585
R880 VDD2.n31 VDD2.n30 585
R881 VDD2.n44 VDD2.t0 329.084
R882 VDD2.n11 VDD2.t1 329.084
R883 VDD2.n64 VDD2.n34 171.744
R884 VDD2.n57 VDD2.n34 171.744
R885 VDD2.n57 VDD2.n56 171.744
R886 VDD2.n56 VDD2.n38 171.744
R887 VDD2.n49 VDD2.n38 171.744
R888 VDD2.n49 VDD2.n48 171.744
R889 VDD2.n48 VDD2.n42 171.744
R890 VDD2.n15 VDD2.n9 171.744
R891 VDD2.n16 VDD2.n15 171.744
R892 VDD2.n16 VDD2.n5 171.744
R893 VDD2.n23 VDD2.n5 171.744
R894 VDD2.n24 VDD2.n23 171.744
R895 VDD2.n24 VDD2.n1 171.744
R896 VDD2.n31 VDD2.n1 171.744
R897 VDD2.t0 VDD2.n42 85.8723
R898 VDD2.t1 VDD2.n9 85.8723
R899 VDD2.n66 VDD2.n32 85.2128
R900 VDD2.n66 VDD2.n65 51.9672
R901 VDD2.n63 VDD2.n33 12.8005
R902 VDD2.n30 VDD2.n0 12.8005
R903 VDD2.n62 VDD2.n35 12.0247
R904 VDD2.n29 VDD2.n2 12.0247
R905 VDD2.n59 VDD2.n58 11.249
R906 VDD2.n26 VDD2.n25 11.249
R907 VDD2.n44 VDD2.n43 10.7233
R908 VDD2.n11 VDD2.n10 10.7233
R909 VDD2.n55 VDD2.n37 10.4732
R910 VDD2.n22 VDD2.n4 10.4732
R911 VDD2.n54 VDD2.n39 9.69747
R912 VDD2.n21 VDD2.n6 9.69747
R913 VDD2.n61 VDD2.n33 9.45567
R914 VDD2.n28 VDD2.n0 9.45567
R915 VDD2.n62 VDD2.n61 9.3005
R916 VDD2.n60 VDD2.n59 9.3005
R917 VDD2.n37 VDD2.n36 9.3005
R918 VDD2.n54 VDD2.n53 9.3005
R919 VDD2.n52 VDD2.n51 9.3005
R920 VDD2.n41 VDD2.n40 9.3005
R921 VDD2.n46 VDD2.n45 9.3005
R922 VDD2.n13 VDD2.n12 9.3005
R923 VDD2.n8 VDD2.n7 9.3005
R924 VDD2.n19 VDD2.n18 9.3005
R925 VDD2.n21 VDD2.n20 9.3005
R926 VDD2.n4 VDD2.n3 9.3005
R927 VDD2.n27 VDD2.n26 9.3005
R928 VDD2.n29 VDD2.n28 9.3005
R929 VDD2.n51 VDD2.n50 8.92171
R930 VDD2.n18 VDD2.n17 8.92171
R931 VDD2.n47 VDD2.n41 8.14595
R932 VDD2.n14 VDD2.n8 8.14595
R933 VDD2.n46 VDD2.n43 7.3702
R934 VDD2.n13 VDD2.n10 7.3702
R935 VDD2.n47 VDD2.n46 5.81868
R936 VDD2.n14 VDD2.n13 5.81868
R937 VDD2.n50 VDD2.n41 5.04292
R938 VDD2.n17 VDD2.n8 5.04292
R939 VDD2.n51 VDD2.n39 4.26717
R940 VDD2.n18 VDD2.n6 4.26717
R941 VDD2.n55 VDD2.n54 3.49141
R942 VDD2.n22 VDD2.n21 3.49141
R943 VDD2.n58 VDD2.n37 2.71565
R944 VDD2.n25 VDD2.n4 2.71565
R945 VDD2.n45 VDD2.n44 2.41347
R946 VDD2.n12 VDD2.n11 2.41347
R947 VDD2.n59 VDD2.n35 1.93989
R948 VDD2.n26 VDD2.n2 1.93989
R949 VDD2.n63 VDD2.n62 1.16414
R950 VDD2.n30 VDD2.n29 1.16414
R951 VDD2 VDD2.n66 0.552224
R952 VDD2.n65 VDD2.n33 0.388379
R953 VDD2.n32 VDD2.n0 0.388379
R954 VDD2.n61 VDD2.n60 0.155672
R955 VDD2.n60 VDD2.n36 0.155672
R956 VDD2.n53 VDD2.n36 0.155672
R957 VDD2.n53 VDD2.n52 0.155672
R958 VDD2.n52 VDD2.n40 0.155672
R959 VDD2.n45 VDD2.n40 0.155672
R960 VDD2.n12 VDD2.n7 0.155672
R961 VDD2.n19 VDD2.n7 0.155672
R962 VDD2.n20 VDD2.n19 0.155672
R963 VDD2.n20 VDD2.n3 0.155672
R964 VDD2.n27 VDD2.n3 0.155672
R965 VDD2.n28 VDD2.n27 0.155672
R966 VP.n0 VP.t0 178.125
R967 VP.n0 VP.t1 139.302
R968 VP VP.n0 0.241678
R969 VDD1.n32 VDD1.n31 756.745
R970 VDD1.n65 VDD1.n64 756.745
R971 VDD1.n31 VDD1.n30 585
R972 VDD1.n2 VDD1.n1 585
R973 VDD1.n25 VDD1.n24 585
R974 VDD1.n23 VDD1.n22 585
R975 VDD1.n6 VDD1.n5 585
R976 VDD1.n17 VDD1.n16 585
R977 VDD1.n15 VDD1.n14 585
R978 VDD1.n10 VDD1.n9 585
R979 VDD1.n43 VDD1.n42 585
R980 VDD1.n48 VDD1.n47 585
R981 VDD1.n50 VDD1.n49 585
R982 VDD1.n39 VDD1.n38 585
R983 VDD1.n56 VDD1.n55 585
R984 VDD1.n58 VDD1.n57 585
R985 VDD1.n35 VDD1.n34 585
R986 VDD1.n64 VDD1.n63 585
R987 VDD1.n11 VDD1.t1 329.084
R988 VDD1.n44 VDD1.t0 329.084
R989 VDD1.n31 VDD1.n1 171.744
R990 VDD1.n24 VDD1.n1 171.744
R991 VDD1.n24 VDD1.n23 171.744
R992 VDD1.n23 VDD1.n5 171.744
R993 VDD1.n16 VDD1.n5 171.744
R994 VDD1.n16 VDD1.n15 171.744
R995 VDD1.n15 VDD1.n9 171.744
R996 VDD1.n48 VDD1.n42 171.744
R997 VDD1.n49 VDD1.n48 171.744
R998 VDD1.n49 VDD1.n38 171.744
R999 VDD1.n56 VDD1.n38 171.744
R1000 VDD1.n57 VDD1.n56 171.744
R1001 VDD1.n57 VDD1.n34 171.744
R1002 VDD1.n64 VDD1.n34 171.744
R1003 VDD1 VDD1.n65 86.2312
R1004 VDD1.t1 VDD1.n9 85.8723
R1005 VDD1.t0 VDD1.n42 85.8723
R1006 VDD1 VDD1.n32 52.5189
R1007 VDD1.n30 VDD1.n0 12.8005
R1008 VDD1.n63 VDD1.n33 12.8005
R1009 VDD1.n29 VDD1.n2 12.0247
R1010 VDD1.n62 VDD1.n35 12.0247
R1011 VDD1.n26 VDD1.n25 11.249
R1012 VDD1.n59 VDD1.n58 11.249
R1013 VDD1.n11 VDD1.n10 10.7233
R1014 VDD1.n44 VDD1.n43 10.7233
R1015 VDD1.n22 VDD1.n4 10.4732
R1016 VDD1.n55 VDD1.n37 10.4732
R1017 VDD1.n21 VDD1.n6 9.69747
R1018 VDD1.n54 VDD1.n39 9.69747
R1019 VDD1.n28 VDD1.n0 9.45567
R1020 VDD1.n61 VDD1.n33 9.45567
R1021 VDD1.n29 VDD1.n28 9.3005
R1022 VDD1.n27 VDD1.n26 9.3005
R1023 VDD1.n4 VDD1.n3 9.3005
R1024 VDD1.n21 VDD1.n20 9.3005
R1025 VDD1.n19 VDD1.n18 9.3005
R1026 VDD1.n8 VDD1.n7 9.3005
R1027 VDD1.n13 VDD1.n12 9.3005
R1028 VDD1.n46 VDD1.n45 9.3005
R1029 VDD1.n41 VDD1.n40 9.3005
R1030 VDD1.n52 VDD1.n51 9.3005
R1031 VDD1.n54 VDD1.n53 9.3005
R1032 VDD1.n37 VDD1.n36 9.3005
R1033 VDD1.n60 VDD1.n59 9.3005
R1034 VDD1.n62 VDD1.n61 9.3005
R1035 VDD1.n18 VDD1.n17 8.92171
R1036 VDD1.n51 VDD1.n50 8.92171
R1037 VDD1.n14 VDD1.n8 8.14595
R1038 VDD1.n47 VDD1.n41 8.14595
R1039 VDD1.n13 VDD1.n10 7.3702
R1040 VDD1.n46 VDD1.n43 7.3702
R1041 VDD1.n14 VDD1.n13 5.81868
R1042 VDD1.n47 VDD1.n46 5.81868
R1043 VDD1.n17 VDD1.n8 5.04292
R1044 VDD1.n50 VDD1.n41 5.04292
R1045 VDD1.n18 VDD1.n6 4.26717
R1046 VDD1.n51 VDD1.n39 4.26717
R1047 VDD1.n22 VDD1.n21 3.49141
R1048 VDD1.n55 VDD1.n54 3.49141
R1049 VDD1.n25 VDD1.n4 2.71565
R1050 VDD1.n58 VDD1.n37 2.71565
R1051 VDD1.n12 VDD1.n11 2.41347
R1052 VDD1.n45 VDD1.n44 2.41347
R1053 VDD1.n26 VDD1.n2 1.93989
R1054 VDD1.n59 VDD1.n35 1.93989
R1055 VDD1.n30 VDD1.n29 1.16414
R1056 VDD1.n63 VDD1.n62 1.16414
R1057 VDD1.n32 VDD1.n0 0.388379
R1058 VDD1.n65 VDD1.n33 0.388379
R1059 VDD1.n28 VDD1.n27 0.155672
R1060 VDD1.n27 VDD1.n3 0.155672
R1061 VDD1.n20 VDD1.n3 0.155672
R1062 VDD1.n20 VDD1.n19 0.155672
R1063 VDD1.n19 VDD1.n7 0.155672
R1064 VDD1.n12 VDD1.n7 0.155672
R1065 VDD1.n45 VDD1.n40 0.155672
R1066 VDD1.n52 VDD1.n40 0.155672
R1067 VDD1.n53 VDD1.n52 0.155672
R1068 VDD1.n53 VDD1.n36 0.155672
R1069 VDD1.n60 VDD1.n36 0.155672
R1070 VDD1.n61 VDD1.n60 0.155672
C0 w_n1886_n2276# B 6.59186f
C1 VP VDD2 0.306037f
C2 VDD1 VN 0.148162f
C3 VTAIL B 2.21654f
C4 VTAIL w_n1886_n2276# 1.97449f
C5 VP B 1.26913f
C6 VDD1 VDD2 0.597878f
C7 w_n1886_n2276# VP 2.68067f
C8 VN VDD2 1.55732f
C9 VTAIL VP 1.49676f
C10 VDD1 B 1.19352f
C11 w_n1886_n2276# VDD1 1.3248f
C12 B VN 0.878996f
C13 w_n1886_n2276# VN 2.44181f
C14 VTAIL VDD1 3.49454f
C15 VTAIL VN 1.48252f
C16 B VDD2 1.21794f
C17 w_n1886_n2276# VDD2 1.34301f
C18 VDD1 VP 1.71344f
C19 VP VN 4.13994f
C20 VTAIL VDD2 3.54166f
C21 VDD2 VSUBS 0.628847f
C22 VDD1 VSUBS 2.215071f
C23 VTAIL VSUBS 0.523695f
C24 VN VSUBS 5.03928f
C25 VP VSUBS 1.196788f
C26 B VSUBS 2.95705f
C27 w_n1886_n2276# VSUBS 53.479397f
C28 VDD1.n0 VSUBS 0.007901f
C29 VDD1.n1 VSUBS 0.017814f
C30 VDD1.n2 VSUBS 0.00798f
C31 VDD1.n3 VSUBS 0.014025f
C32 VDD1.n4 VSUBS 0.007537f
C33 VDD1.n5 VSUBS 0.017814f
C34 VDD1.n6 VSUBS 0.00798f
C35 VDD1.n7 VSUBS 0.014025f
C36 VDD1.n8 VSUBS 0.007537f
C37 VDD1.n9 VSUBS 0.01336f
C38 VDD1.n10 VSUBS 0.013399f
C39 VDD1.t1 VSUBS 0.038306f
C40 VDD1.n11 VSUBS 0.075977f
C41 VDD1.n12 VSUBS 0.353249f
C42 VDD1.n13 VSUBS 0.007537f
C43 VDD1.n14 VSUBS 0.00798f
C44 VDD1.n15 VSUBS 0.017814f
C45 VDD1.n16 VSUBS 0.017814f
C46 VDD1.n17 VSUBS 0.00798f
C47 VDD1.n18 VSUBS 0.007537f
C48 VDD1.n19 VSUBS 0.014025f
C49 VDD1.n20 VSUBS 0.014025f
C50 VDD1.n21 VSUBS 0.007537f
C51 VDD1.n22 VSUBS 0.00798f
C52 VDD1.n23 VSUBS 0.017814f
C53 VDD1.n24 VSUBS 0.017814f
C54 VDD1.n25 VSUBS 0.00798f
C55 VDD1.n26 VSUBS 0.007537f
C56 VDD1.n27 VSUBS 0.014025f
C57 VDD1.n28 VSUBS 0.035868f
C58 VDD1.n29 VSUBS 0.007537f
C59 VDD1.n30 VSUBS 0.00798f
C60 VDD1.n31 VSUBS 0.04009f
C61 VDD1.n32 VSUBS 0.036747f
C62 VDD1.n33 VSUBS 0.007901f
C63 VDD1.n34 VSUBS 0.017814f
C64 VDD1.n35 VSUBS 0.00798f
C65 VDD1.n36 VSUBS 0.014025f
C66 VDD1.n37 VSUBS 0.007537f
C67 VDD1.n38 VSUBS 0.017814f
C68 VDD1.n39 VSUBS 0.00798f
C69 VDD1.n40 VSUBS 0.014025f
C70 VDD1.n41 VSUBS 0.007537f
C71 VDD1.n42 VSUBS 0.01336f
C72 VDD1.n43 VSUBS 0.013399f
C73 VDD1.t0 VSUBS 0.038306f
C74 VDD1.n44 VSUBS 0.075977f
C75 VDD1.n45 VSUBS 0.353249f
C76 VDD1.n46 VSUBS 0.007537f
C77 VDD1.n47 VSUBS 0.00798f
C78 VDD1.n48 VSUBS 0.017814f
C79 VDD1.n49 VSUBS 0.017814f
C80 VDD1.n50 VSUBS 0.00798f
C81 VDD1.n51 VSUBS 0.007537f
C82 VDD1.n52 VSUBS 0.014025f
C83 VDD1.n53 VSUBS 0.014025f
C84 VDD1.n54 VSUBS 0.007537f
C85 VDD1.n55 VSUBS 0.00798f
C86 VDD1.n56 VSUBS 0.017814f
C87 VDD1.n57 VSUBS 0.017814f
C88 VDD1.n58 VSUBS 0.00798f
C89 VDD1.n59 VSUBS 0.007537f
C90 VDD1.n60 VSUBS 0.014025f
C91 VDD1.n61 VSUBS 0.035868f
C92 VDD1.n62 VSUBS 0.007537f
C93 VDD1.n63 VSUBS 0.00798f
C94 VDD1.n64 VSUBS 0.04009f
C95 VDD1.n65 VSUBS 0.306047f
C96 VP.t0 VSUBS 1.95517f
C97 VP.t1 VSUBS 1.5573f
C98 VP.n0 VSUBS 3.22618f
C99 VDD2.n0 VSUBS 0.00802f
C100 VDD2.n1 VSUBS 0.018081f
C101 VDD2.n2 VSUBS 0.0081f
C102 VDD2.n3 VSUBS 0.014236f
C103 VDD2.n4 VSUBS 0.00765f
C104 VDD2.n5 VSUBS 0.018081f
C105 VDD2.n6 VSUBS 0.0081f
C106 VDD2.n7 VSUBS 0.014236f
C107 VDD2.n8 VSUBS 0.00765f
C108 VDD2.n9 VSUBS 0.013561f
C109 VDD2.n10 VSUBS 0.0136f
C110 VDD2.t1 VSUBS 0.038881f
C111 VDD2.n11 VSUBS 0.077118f
C112 VDD2.n12 VSUBS 0.358556f
C113 VDD2.n13 VSUBS 0.00765f
C114 VDD2.n14 VSUBS 0.0081f
C115 VDD2.n15 VSUBS 0.018081f
C116 VDD2.n16 VSUBS 0.018081f
C117 VDD2.n17 VSUBS 0.0081f
C118 VDD2.n18 VSUBS 0.00765f
C119 VDD2.n19 VSUBS 0.014236f
C120 VDD2.n20 VSUBS 0.014236f
C121 VDD2.n21 VSUBS 0.00765f
C122 VDD2.n22 VSUBS 0.0081f
C123 VDD2.n23 VSUBS 0.018081f
C124 VDD2.n24 VSUBS 0.018081f
C125 VDD2.n25 VSUBS 0.0081f
C126 VDD2.n26 VSUBS 0.00765f
C127 VDD2.n27 VSUBS 0.014236f
C128 VDD2.n28 VSUBS 0.036406f
C129 VDD2.n29 VSUBS 0.00765f
C130 VDD2.n30 VSUBS 0.0081f
C131 VDD2.n31 VSUBS 0.040692f
C132 VDD2.n32 VSUBS 0.289118f
C133 VDD2.n33 VSUBS 0.00802f
C134 VDD2.n34 VSUBS 0.018081f
C135 VDD2.n35 VSUBS 0.0081f
C136 VDD2.n36 VSUBS 0.014236f
C137 VDD2.n37 VSUBS 0.00765f
C138 VDD2.n38 VSUBS 0.018081f
C139 VDD2.n39 VSUBS 0.0081f
C140 VDD2.n40 VSUBS 0.014236f
C141 VDD2.n41 VSUBS 0.00765f
C142 VDD2.n42 VSUBS 0.013561f
C143 VDD2.n43 VSUBS 0.0136f
C144 VDD2.t0 VSUBS 0.038881f
C145 VDD2.n44 VSUBS 0.077118f
C146 VDD2.n45 VSUBS 0.358556f
C147 VDD2.n46 VSUBS 0.00765f
C148 VDD2.n47 VSUBS 0.0081f
C149 VDD2.n48 VSUBS 0.018081f
C150 VDD2.n49 VSUBS 0.018081f
C151 VDD2.n50 VSUBS 0.0081f
C152 VDD2.n51 VSUBS 0.00765f
C153 VDD2.n52 VSUBS 0.014236f
C154 VDD2.n53 VSUBS 0.014236f
C155 VDD2.n54 VSUBS 0.00765f
C156 VDD2.n55 VSUBS 0.0081f
C157 VDD2.n56 VSUBS 0.018081f
C158 VDD2.n57 VSUBS 0.018081f
C159 VDD2.n58 VSUBS 0.0081f
C160 VDD2.n59 VSUBS 0.00765f
C161 VDD2.n60 VSUBS 0.014236f
C162 VDD2.n61 VSUBS 0.036406f
C163 VDD2.n62 VSUBS 0.00765f
C164 VDD2.n63 VSUBS 0.0081f
C165 VDD2.n64 VSUBS 0.040692f
C166 VDD2.n65 VSUBS 0.036726f
C167 VDD2.n66 VSUBS 1.34967f
C168 VTAIL.n0 VSUBS 0.011732f
C169 VTAIL.n1 VSUBS 0.026451f
C170 VTAIL.n2 VSUBS 0.011849f
C171 VTAIL.n3 VSUBS 0.020825f
C172 VTAIL.n4 VSUBS 0.011191f
C173 VTAIL.n5 VSUBS 0.026451f
C174 VTAIL.n6 VSUBS 0.011849f
C175 VTAIL.n7 VSUBS 0.020825f
C176 VTAIL.n8 VSUBS 0.011191f
C177 VTAIL.n9 VSUBS 0.019838f
C178 VTAIL.n10 VSUBS 0.019895f
C179 VTAIL.t0 VSUBS 0.056878f
C180 VTAIL.n11 VSUBS 0.112814f
C181 VTAIL.n12 VSUBS 0.524521f
C182 VTAIL.n13 VSUBS 0.011191f
C183 VTAIL.n14 VSUBS 0.011849f
C184 VTAIL.n15 VSUBS 0.026451f
C185 VTAIL.n16 VSUBS 0.026451f
C186 VTAIL.n17 VSUBS 0.011849f
C187 VTAIL.n18 VSUBS 0.011191f
C188 VTAIL.n19 VSUBS 0.020825f
C189 VTAIL.n20 VSUBS 0.020825f
C190 VTAIL.n21 VSUBS 0.011191f
C191 VTAIL.n22 VSUBS 0.011849f
C192 VTAIL.n23 VSUBS 0.026451f
C193 VTAIL.n24 VSUBS 0.026451f
C194 VTAIL.n25 VSUBS 0.011849f
C195 VTAIL.n26 VSUBS 0.011191f
C196 VTAIL.n27 VSUBS 0.020825f
C197 VTAIL.n28 VSUBS 0.053258f
C198 VTAIL.n29 VSUBS 0.011191f
C199 VTAIL.n30 VSUBS 0.011849f
C200 VTAIL.n31 VSUBS 0.059528f
C201 VTAIL.n32 VSUBS 0.039379f
C202 VTAIL.n33 VSUBS 1.01507f
C203 VTAIL.n34 VSUBS 0.011732f
C204 VTAIL.n35 VSUBS 0.026451f
C205 VTAIL.n36 VSUBS 0.011849f
C206 VTAIL.n37 VSUBS 0.020825f
C207 VTAIL.n38 VSUBS 0.011191f
C208 VTAIL.n39 VSUBS 0.026451f
C209 VTAIL.n40 VSUBS 0.011849f
C210 VTAIL.n41 VSUBS 0.020825f
C211 VTAIL.n42 VSUBS 0.011191f
C212 VTAIL.n43 VSUBS 0.019838f
C213 VTAIL.n44 VSUBS 0.019895f
C214 VTAIL.t2 VSUBS 0.056878f
C215 VTAIL.n45 VSUBS 0.112814f
C216 VTAIL.n46 VSUBS 0.524521f
C217 VTAIL.n47 VSUBS 0.011191f
C218 VTAIL.n48 VSUBS 0.011849f
C219 VTAIL.n49 VSUBS 0.026451f
C220 VTAIL.n50 VSUBS 0.026451f
C221 VTAIL.n51 VSUBS 0.011849f
C222 VTAIL.n52 VSUBS 0.011191f
C223 VTAIL.n53 VSUBS 0.020825f
C224 VTAIL.n54 VSUBS 0.020825f
C225 VTAIL.n55 VSUBS 0.011191f
C226 VTAIL.n56 VSUBS 0.011849f
C227 VTAIL.n57 VSUBS 0.026451f
C228 VTAIL.n58 VSUBS 0.026451f
C229 VTAIL.n59 VSUBS 0.011849f
C230 VTAIL.n60 VSUBS 0.011191f
C231 VTAIL.n61 VSUBS 0.020825f
C232 VTAIL.n62 VSUBS 0.053258f
C233 VTAIL.n63 VSUBS 0.011191f
C234 VTAIL.n64 VSUBS 0.011849f
C235 VTAIL.n65 VSUBS 0.059528f
C236 VTAIL.n66 VSUBS 0.039379f
C237 VTAIL.n67 VSUBS 1.04429f
C238 VTAIL.n68 VSUBS 0.011732f
C239 VTAIL.n69 VSUBS 0.026451f
C240 VTAIL.n70 VSUBS 0.011849f
C241 VTAIL.n71 VSUBS 0.020825f
C242 VTAIL.n72 VSUBS 0.011191f
C243 VTAIL.n73 VSUBS 0.026451f
C244 VTAIL.n74 VSUBS 0.011849f
C245 VTAIL.n75 VSUBS 0.020825f
C246 VTAIL.n76 VSUBS 0.011191f
C247 VTAIL.n77 VSUBS 0.019838f
C248 VTAIL.n78 VSUBS 0.019895f
C249 VTAIL.t1 VSUBS 0.056878f
C250 VTAIL.n79 VSUBS 0.112814f
C251 VTAIL.n80 VSUBS 0.524521f
C252 VTAIL.n81 VSUBS 0.011191f
C253 VTAIL.n82 VSUBS 0.011849f
C254 VTAIL.n83 VSUBS 0.026451f
C255 VTAIL.n84 VSUBS 0.026451f
C256 VTAIL.n85 VSUBS 0.011849f
C257 VTAIL.n86 VSUBS 0.011191f
C258 VTAIL.n87 VSUBS 0.020825f
C259 VTAIL.n88 VSUBS 0.020825f
C260 VTAIL.n89 VSUBS 0.011191f
C261 VTAIL.n90 VSUBS 0.011849f
C262 VTAIL.n91 VSUBS 0.026451f
C263 VTAIL.n92 VSUBS 0.026451f
C264 VTAIL.n93 VSUBS 0.011849f
C265 VTAIL.n94 VSUBS 0.011191f
C266 VTAIL.n95 VSUBS 0.020825f
C267 VTAIL.n96 VSUBS 0.053258f
C268 VTAIL.n97 VSUBS 0.011191f
C269 VTAIL.n98 VSUBS 0.011849f
C270 VTAIL.n99 VSUBS 0.059528f
C271 VTAIL.n100 VSUBS 0.039379f
C272 VTAIL.n101 VSUBS 0.911814f
C273 VTAIL.n102 VSUBS 0.011732f
C274 VTAIL.n103 VSUBS 0.026451f
C275 VTAIL.n104 VSUBS 0.011849f
C276 VTAIL.n105 VSUBS 0.020825f
C277 VTAIL.n106 VSUBS 0.011191f
C278 VTAIL.n107 VSUBS 0.026451f
C279 VTAIL.n108 VSUBS 0.011849f
C280 VTAIL.n109 VSUBS 0.020825f
C281 VTAIL.n110 VSUBS 0.011191f
C282 VTAIL.n111 VSUBS 0.019838f
C283 VTAIL.n112 VSUBS 0.019895f
C284 VTAIL.t3 VSUBS 0.056878f
C285 VTAIL.n113 VSUBS 0.112814f
C286 VTAIL.n114 VSUBS 0.524521f
C287 VTAIL.n115 VSUBS 0.011191f
C288 VTAIL.n116 VSUBS 0.011849f
C289 VTAIL.n117 VSUBS 0.026451f
C290 VTAIL.n118 VSUBS 0.026451f
C291 VTAIL.n119 VSUBS 0.011849f
C292 VTAIL.n120 VSUBS 0.011191f
C293 VTAIL.n121 VSUBS 0.020825f
C294 VTAIL.n122 VSUBS 0.020825f
C295 VTAIL.n123 VSUBS 0.011191f
C296 VTAIL.n124 VSUBS 0.011849f
C297 VTAIL.n125 VSUBS 0.026451f
C298 VTAIL.n126 VSUBS 0.026451f
C299 VTAIL.n127 VSUBS 0.011849f
C300 VTAIL.n128 VSUBS 0.011191f
C301 VTAIL.n129 VSUBS 0.020825f
C302 VTAIL.n130 VSUBS 0.053258f
C303 VTAIL.n131 VSUBS 0.011191f
C304 VTAIL.n132 VSUBS 0.011849f
C305 VTAIL.n133 VSUBS 0.059528f
C306 VTAIL.n134 VSUBS 0.039379f
C307 VTAIL.n135 VSUBS 0.843264f
C308 VN.t0 VSUBS 1.47806f
C309 VN.t1 VSUBS 1.85979f
C310 B.n0 VSUBS 0.006895f
C311 B.n1 VSUBS 0.006895f
C312 B.n2 VSUBS 0.010197f
C313 B.n3 VSUBS 0.007814f
C314 B.n4 VSUBS 0.007814f
C315 B.n5 VSUBS 0.007814f
C316 B.n6 VSUBS 0.007814f
C317 B.n7 VSUBS 0.007814f
C318 B.n8 VSUBS 0.007814f
C319 B.n9 VSUBS 0.007814f
C320 B.n10 VSUBS 0.007814f
C321 B.n11 VSUBS 0.007814f
C322 B.n12 VSUBS 0.017288f
C323 B.n13 VSUBS 0.007814f
C324 B.n14 VSUBS 0.007814f
C325 B.n15 VSUBS 0.007814f
C326 B.n16 VSUBS 0.007814f
C327 B.n17 VSUBS 0.007814f
C328 B.n18 VSUBS 0.007814f
C329 B.n19 VSUBS 0.007814f
C330 B.n20 VSUBS 0.007814f
C331 B.n21 VSUBS 0.007814f
C332 B.n22 VSUBS 0.007814f
C333 B.n23 VSUBS 0.007814f
C334 B.n24 VSUBS 0.007814f
C335 B.n25 VSUBS 0.007814f
C336 B.t7 VSUBS 0.110313f
C337 B.t8 VSUBS 0.134032f
C338 B.t6 VSUBS 0.663433f
C339 B.n26 VSUBS 0.23056f
C340 B.n27 VSUBS 0.183046f
C341 B.n28 VSUBS 0.007814f
C342 B.n29 VSUBS 0.007814f
C343 B.n30 VSUBS 0.007814f
C344 B.n31 VSUBS 0.007814f
C345 B.t10 VSUBS 0.110316f
C346 B.t11 VSUBS 0.134034f
C347 B.t9 VSUBS 0.663433f
C348 B.n32 VSUBS 0.230559f
C349 B.n33 VSUBS 0.183044f
C350 B.n34 VSUBS 0.018104f
C351 B.n35 VSUBS 0.007814f
C352 B.n36 VSUBS 0.007814f
C353 B.n37 VSUBS 0.007814f
C354 B.n38 VSUBS 0.007814f
C355 B.n39 VSUBS 0.007814f
C356 B.n40 VSUBS 0.007814f
C357 B.n41 VSUBS 0.007814f
C358 B.n42 VSUBS 0.007814f
C359 B.n43 VSUBS 0.007814f
C360 B.n44 VSUBS 0.007814f
C361 B.n45 VSUBS 0.007814f
C362 B.n46 VSUBS 0.007814f
C363 B.n47 VSUBS 0.018564f
C364 B.n48 VSUBS 0.007814f
C365 B.n49 VSUBS 0.007814f
C366 B.n50 VSUBS 0.007814f
C367 B.n51 VSUBS 0.007814f
C368 B.n52 VSUBS 0.007814f
C369 B.n53 VSUBS 0.007814f
C370 B.n54 VSUBS 0.007814f
C371 B.n55 VSUBS 0.007814f
C372 B.n56 VSUBS 0.007814f
C373 B.n57 VSUBS 0.007814f
C374 B.n58 VSUBS 0.007814f
C375 B.n59 VSUBS 0.007814f
C376 B.n60 VSUBS 0.007814f
C377 B.n61 VSUBS 0.007814f
C378 B.n62 VSUBS 0.007814f
C379 B.n63 VSUBS 0.007814f
C380 B.n64 VSUBS 0.007814f
C381 B.n65 VSUBS 0.007814f
C382 B.n66 VSUBS 0.007814f
C383 B.n67 VSUBS 0.007814f
C384 B.n68 VSUBS 0.007814f
C385 B.n69 VSUBS 0.017288f
C386 B.n70 VSUBS 0.007814f
C387 B.n71 VSUBS 0.007814f
C388 B.n72 VSUBS 0.007814f
C389 B.n73 VSUBS 0.007814f
C390 B.n74 VSUBS 0.007814f
C391 B.n75 VSUBS 0.007814f
C392 B.n76 VSUBS 0.007814f
C393 B.n77 VSUBS 0.007814f
C394 B.n78 VSUBS 0.007814f
C395 B.n79 VSUBS 0.007814f
C396 B.n80 VSUBS 0.007814f
C397 B.n81 VSUBS 0.007814f
C398 B.n82 VSUBS 0.005401f
C399 B.n83 VSUBS 0.007814f
C400 B.n84 VSUBS 0.007814f
C401 B.n85 VSUBS 0.007814f
C402 B.n86 VSUBS 0.007814f
C403 B.n87 VSUBS 0.007814f
C404 B.t5 VSUBS 0.110313f
C405 B.t4 VSUBS 0.134032f
C406 B.t3 VSUBS 0.663433f
C407 B.n88 VSUBS 0.23056f
C408 B.n89 VSUBS 0.183046f
C409 B.n90 VSUBS 0.007814f
C410 B.n91 VSUBS 0.007814f
C411 B.n92 VSUBS 0.007814f
C412 B.n93 VSUBS 0.007814f
C413 B.n94 VSUBS 0.007814f
C414 B.n95 VSUBS 0.007814f
C415 B.n96 VSUBS 0.007814f
C416 B.n97 VSUBS 0.007814f
C417 B.n98 VSUBS 0.007814f
C418 B.n99 VSUBS 0.007814f
C419 B.n100 VSUBS 0.007814f
C420 B.n101 VSUBS 0.007814f
C421 B.n102 VSUBS 0.017288f
C422 B.n103 VSUBS 0.007814f
C423 B.n104 VSUBS 0.007814f
C424 B.n105 VSUBS 0.007814f
C425 B.n106 VSUBS 0.007814f
C426 B.n107 VSUBS 0.007814f
C427 B.n108 VSUBS 0.007814f
C428 B.n109 VSUBS 0.007814f
C429 B.n110 VSUBS 0.007814f
C430 B.n111 VSUBS 0.007814f
C431 B.n112 VSUBS 0.007814f
C432 B.n113 VSUBS 0.007814f
C433 B.n114 VSUBS 0.007814f
C434 B.n115 VSUBS 0.007814f
C435 B.n116 VSUBS 0.007814f
C436 B.n117 VSUBS 0.007814f
C437 B.n118 VSUBS 0.007814f
C438 B.n119 VSUBS 0.007814f
C439 B.n120 VSUBS 0.007814f
C440 B.n121 VSUBS 0.007814f
C441 B.n122 VSUBS 0.007814f
C442 B.n123 VSUBS 0.007814f
C443 B.n124 VSUBS 0.007814f
C444 B.n125 VSUBS 0.007814f
C445 B.n126 VSUBS 0.007814f
C446 B.n127 VSUBS 0.007814f
C447 B.n128 VSUBS 0.007814f
C448 B.n129 VSUBS 0.007814f
C449 B.n130 VSUBS 0.007814f
C450 B.n131 VSUBS 0.007814f
C451 B.n132 VSUBS 0.007814f
C452 B.n133 VSUBS 0.007814f
C453 B.n134 VSUBS 0.007814f
C454 B.n135 VSUBS 0.007814f
C455 B.n136 VSUBS 0.007814f
C456 B.n137 VSUBS 0.007814f
C457 B.n138 VSUBS 0.007814f
C458 B.n139 VSUBS 0.007814f
C459 B.n140 VSUBS 0.007814f
C460 B.n141 VSUBS 0.017288f
C461 B.n142 VSUBS 0.018564f
C462 B.n143 VSUBS 0.018564f
C463 B.n144 VSUBS 0.007814f
C464 B.n145 VSUBS 0.007814f
C465 B.n146 VSUBS 0.007814f
C466 B.n147 VSUBS 0.007814f
C467 B.n148 VSUBS 0.007814f
C468 B.n149 VSUBS 0.007814f
C469 B.n150 VSUBS 0.007814f
C470 B.n151 VSUBS 0.007814f
C471 B.n152 VSUBS 0.007814f
C472 B.n153 VSUBS 0.007814f
C473 B.n154 VSUBS 0.007814f
C474 B.n155 VSUBS 0.007814f
C475 B.n156 VSUBS 0.007814f
C476 B.n157 VSUBS 0.007814f
C477 B.n158 VSUBS 0.007814f
C478 B.n159 VSUBS 0.007814f
C479 B.n160 VSUBS 0.007814f
C480 B.n161 VSUBS 0.007814f
C481 B.n162 VSUBS 0.007814f
C482 B.n163 VSUBS 0.007814f
C483 B.n164 VSUBS 0.007814f
C484 B.n165 VSUBS 0.007814f
C485 B.n166 VSUBS 0.007814f
C486 B.n167 VSUBS 0.007814f
C487 B.n168 VSUBS 0.007814f
C488 B.n169 VSUBS 0.007814f
C489 B.n170 VSUBS 0.007814f
C490 B.n171 VSUBS 0.007814f
C491 B.n172 VSUBS 0.007814f
C492 B.n173 VSUBS 0.007814f
C493 B.n174 VSUBS 0.007814f
C494 B.n175 VSUBS 0.007814f
C495 B.n176 VSUBS 0.007814f
C496 B.n177 VSUBS 0.007814f
C497 B.n178 VSUBS 0.007814f
C498 B.n179 VSUBS 0.007814f
C499 B.n180 VSUBS 0.005401f
C500 B.n181 VSUBS 0.018104f
C501 B.n182 VSUBS 0.00632f
C502 B.n183 VSUBS 0.007814f
C503 B.n184 VSUBS 0.007814f
C504 B.n185 VSUBS 0.007814f
C505 B.n186 VSUBS 0.007814f
C506 B.n187 VSUBS 0.007814f
C507 B.n188 VSUBS 0.007814f
C508 B.n189 VSUBS 0.007814f
C509 B.n190 VSUBS 0.007814f
C510 B.n191 VSUBS 0.007814f
C511 B.n192 VSUBS 0.007814f
C512 B.n193 VSUBS 0.007814f
C513 B.t2 VSUBS 0.110316f
C514 B.t1 VSUBS 0.134034f
C515 B.t0 VSUBS 0.663433f
C516 B.n194 VSUBS 0.230559f
C517 B.n195 VSUBS 0.183044f
C518 B.n196 VSUBS 0.018104f
C519 B.n197 VSUBS 0.00632f
C520 B.n198 VSUBS 0.007814f
C521 B.n199 VSUBS 0.007814f
C522 B.n200 VSUBS 0.007814f
C523 B.n201 VSUBS 0.007814f
C524 B.n202 VSUBS 0.007814f
C525 B.n203 VSUBS 0.007814f
C526 B.n204 VSUBS 0.007814f
C527 B.n205 VSUBS 0.007814f
C528 B.n206 VSUBS 0.007814f
C529 B.n207 VSUBS 0.007814f
C530 B.n208 VSUBS 0.007814f
C531 B.n209 VSUBS 0.007814f
C532 B.n210 VSUBS 0.007814f
C533 B.n211 VSUBS 0.007814f
C534 B.n212 VSUBS 0.007814f
C535 B.n213 VSUBS 0.007814f
C536 B.n214 VSUBS 0.007814f
C537 B.n215 VSUBS 0.007814f
C538 B.n216 VSUBS 0.007814f
C539 B.n217 VSUBS 0.007814f
C540 B.n218 VSUBS 0.007814f
C541 B.n219 VSUBS 0.007814f
C542 B.n220 VSUBS 0.007814f
C543 B.n221 VSUBS 0.007814f
C544 B.n222 VSUBS 0.007814f
C545 B.n223 VSUBS 0.007814f
C546 B.n224 VSUBS 0.007814f
C547 B.n225 VSUBS 0.007814f
C548 B.n226 VSUBS 0.007814f
C549 B.n227 VSUBS 0.007814f
C550 B.n228 VSUBS 0.007814f
C551 B.n229 VSUBS 0.007814f
C552 B.n230 VSUBS 0.007814f
C553 B.n231 VSUBS 0.007814f
C554 B.n232 VSUBS 0.007814f
C555 B.n233 VSUBS 0.007814f
C556 B.n234 VSUBS 0.007814f
C557 B.n235 VSUBS 0.007814f
C558 B.n236 VSUBS 0.018564f
C559 B.n237 VSUBS 0.017613f
C560 B.n238 VSUBS 0.01824f
C561 B.n239 VSUBS 0.007814f
C562 B.n240 VSUBS 0.007814f
C563 B.n241 VSUBS 0.007814f
C564 B.n242 VSUBS 0.007814f
C565 B.n243 VSUBS 0.007814f
C566 B.n244 VSUBS 0.007814f
C567 B.n245 VSUBS 0.007814f
C568 B.n246 VSUBS 0.007814f
C569 B.n247 VSUBS 0.007814f
C570 B.n248 VSUBS 0.007814f
C571 B.n249 VSUBS 0.007814f
C572 B.n250 VSUBS 0.007814f
C573 B.n251 VSUBS 0.007814f
C574 B.n252 VSUBS 0.007814f
C575 B.n253 VSUBS 0.007814f
C576 B.n254 VSUBS 0.007814f
C577 B.n255 VSUBS 0.007814f
C578 B.n256 VSUBS 0.007814f
C579 B.n257 VSUBS 0.007814f
C580 B.n258 VSUBS 0.007814f
C581 B.n259 VSUBS 0.007814f
C582 B.n260 VSUBS 0.007814f
C583 B.n261 VSUBS 0.007814f
C584 B.n262 VSUBS 0.007814f
C585 B.n263 VSUBS 0.007814f
C586 B.n264 VSUBS 0.007814f
C587 B.n265 VSUBS 0.007814f
C588 B.n266 VSUBS 0.007814f
C589 B.n267 VSUBS 0.007814f
C590 B.n268 VSUBS 0.007814f
C591 B.n269 VSUBS 0.007814f
C592 B.n270 VSUBS 0.007814f
C593 B.n271 VSUBS 0.007814f
C594 B.n272 VSUBS 0.007814f
C595 B.n273 VSUBS 0.007814f
C596 B.n274 VSUBS 0.007814f
C597 B.n275 VSUBS 0.007814f
C598 B.n276 VSUBS 0.007814f
C599 B.n277 VSUBS 0.007814f
C600 B.n278 VSUBS 0.007814f
C601 B.n279 VSUBS 0.007814f
C602 B.n280 VSUBS 0.007814f
C603 B.n281 VSUBS 0.007814f
C604 B.n282 VSUBS 0.007814f
C605 B.n283 VSUBS 0.007814f
C606 B.n284 VSUBS 0.007814f
C607 B.n285 VSUBS 0.007814f
C608 B.n286 VSUBS 0.007814f
C609 B.n287 VSUBS 0.007814f
C610 B.n288 VSUBS 0.007814f
C611 B.n289 VSUBS 0.007814f
C612 B.n290 VSUBS 0.007814f
C613 B.n291 VSUBS 0.007814f
C614 B.n292 VSUBS 0.007814f
C615 B.n293 VSUBS 0.007814f
C616 B.n294 VSUBS 0.007814f
C617 B.n295 VSUBS 0.007814f
C618 B.n296 VSUBS 0.007814f
C619 B.n297 VSUBS 0.007814f
C620 B.n298 VSUBS 0.007814f
C621 B.n299 VSUBS 0.007814f
C622 B.n300 VSUBS 0.007814f
C623 B.n301 VSUBS 0.007814f
C624 B.n302 VSUBS 0.017288f
C625 B.n303 VSUBS 0.017288f
C626 B.n304 VSUBS 0.018564f
C627 B.n305 VSUBS 0.007814f
C628 B.n306 VSUBS 0.007814f
C629 B.n307 VSUBS 0.007814f
C630 B.n308 VSUBS 0.007814f
C631 B.n309 VSUBS 0.007814f
C632 B.n310 VSUBS 0.007814f
C633 B.n311 VSUBS 0.007814f
C634 B.n312 VSUBS 0.007814f
C635 B.n313 VSUBS 0.007814f
C636 B.n314 VSUBS 0.007814f
C637 B.n315 VSUBS 0.007814f
C638 B.n316 VSUBS 0.007814f
C639 B.n317 VSUBS 0.007814f
C640 B.n318 VSUBS 0.007814f
C641 B.n319 VSUBS 0.007814f
C642 B.n320 VSUBS 0.007814f
C643 B.n321 VSUBS 0.007814f
C644 B.n322 VSUBS 0.007814f
C645 B.n323 VSUBS 0.007814f
C646 B.n324 VSUBS 0.007814f
C647 B.n325 VSUBS 0.007814f
C648 B.n326 VSUBS 0.007814f
C649 B.n327 VSUBS 0.007814f
C650 B.n328 VSUBS 0.007814f
C651 B.n329 VSUBS 0.007814f
C652 B.n330 VSUBS 0.007814f
C653 B.n331 VSUBS 0.007814f
C654 B.n332 VSUBS 0.007814f
C655 B.n333 VSUBS 0.007814f
C656 B.n334 VSUBS 0.007814f
C657 B.n335 VSUBS 0.007814f
C658 B.n336 VSUBS 0.007814f
C659 B.n337 VSUBS 0.007814f
C660 B.n338 VSUBS 0.007814f
C661 B.n339 VSUBS 0.007814f
C662 B.n340 VSUBS 0.007814f
C663 B.n341 VSUBS 0.005401f
C664 B.n342 VSUBS 0.007814f
C665 B.n343 VSUBS 0.007814f
C666 B.n344 VSUBS 0.00632f
C667 B.n345 VSUBS 0.007814f
C668 B.n346 VSUBS 0.007814f
C669 B.n347 VSUBS 0.007814f
C670 B.n348 VSUBS 0.007814f
C671 B.n349 VSUBS 0.007814f
C672 B.n350 VSUBS 0.007814f
C673 B.n351 VSUBS 0.007814f
C674 B.n352 VSUBS 0.007814f
C675 B.n353 VSUBS 0.007814f
C676 B.n354 VSUBS 0.007814f
C677 B.n355 VSUBS 0.007814f
C678 B.n356 VSUBS 0.00632f
C679 B.n357 VSUBS 0.018104f
C680 B.n358 VSUBS 0.005401f
C681 B.n359 VSUBS 0.007814f
C682 B.n360 VSUBS 0.007814f
C683 B.n361 VSUBS 0.007814f
C684 B.n362 VSUBS 0.007814f
C685 B.n363 VSUBS 0.007814f
C686 B.n364 VSUBS 0.007814f
C687 B.n365 VSUBS 0.007814f
C688 B.n366 VSUBS 0.007814f
C689 B.n367 VSUBS 0.007814f
C690 B.n368 VSUBS 0.007814f
C691 B.n369 VSUBS 0.007814f
C692 B.n370 VSUBS 0.007814f
C693 B.n371 VSUBS 0.007814f
C694 B.n372 VSUBS 0.007814f
C695 B.n373 VSUBS 0.007814f
C696 B.n374 VSUBS 0.007814f
C697 B.n375 VSUBS 0.007814f
C698 B.n376 VSUBS 0.007814f
C699 B.n377 VSUBS 0.007814f
C700 B.n378 VSUBS 0.007814f
C701 B.n379 VSUBS 0.007814f
C702 B.n380 VSUBS 0.007814f
C703 B.n381 VSUBS 0.007814f
C704 B.n382 VSUBS 0.007814f
C705 B.n383 VSUBS 0.007814f
C706 B.n384 VSUBS 0.007814f
C707 B.n385 VSUBS 0.007814f
C708 B.n386 VSUBS 0.007814f
C709 B.n387 VSUBS 0.007814f
C710 B.n388 VSUBS 0.007814f
C711 B.n389 VSUBS 0.007814f
C712 B.n390 VSUBS 0.007814f
C713 B.n391 VSUBS 0.007814f
C714 B.n392 VSUBS 0.007814f
C715 B.n393 VSUBS 0.007814f
C716 B.n394 VSUBS 0.007814f
C717 B.n395 VSUBS 0.018564f
C718 B.n396 VSUBS 0.018564f
C719 B.n397 VSUBS 0.017288f
C720 B.n398 VSUBS 0.007814f
C721 B.n399 VSUBS 0.007814f
C722 B.n400 VSUBS 0.007814f
C723 B.n401 VSUBS 0.007814f
C724 B.n402 VSUBS 0.007814f
C725 B.n403 VSUBS 0.007814f
C726 B.n404 VSUBS 0.007814f
C727 B.n405 VSUBS 0.007814f
C728 B.n406 VSUBS 0.007814f
C729 B.n407 VSUBS 0.007814f
C730 B.n408 VSUBS 0.007814f
C731 B.n409 VSUBS 0.007814f
C732 B.n410 VSUBS 0.007814f
C733 B.n411 VSUBS 0.007814f
C734 B.n412 VSUBS 0.007814f
C735 B.n413 VSUBS 0.007814f
C736 B.n414 VSUBS 0.007814f
C737 B.n415 VSUBS 0.007814f
C738 B.n416 VSUBS 0.007814f
C739 B.n417 VSUBS 0.007814f
C740 B.n418 VSUBS 0.007814f
C741 B.n419 VSUBS 0.007814f
C742 B.n420 VSUBS 0.007814f
C743 B.n421 VSUBS 0.007814f
C744 B.n422 VSUBS 0.007814f
C745 B.n423 VSUBS 0.007814f
C746 B.n424 VSUBS 0.007814f
C747 B.n425 VSUBS 0.007814f
C748 B.n426 VSUBS 0.007814f
C749 B.n427 VSUBS 0.010197f
C750 B.n428 VSUBS 0.010862f
C751 B.n429 VSUBS 0.0216f
.ends

