* NGSPICE file created from diff_pair_sample_0095.ext - technology: sky130A

.subckt diff_pair_sample_0095 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=0 ps=0 w=7.59 l=2.75
X1 B.t8 B.t6 B.t7 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=0 ps=0 w=7.59 l=2.75
X2 VDD1.t9 VP.t0 VTAIL.t10 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=1.25235 ps=7.92 w=7.59 l=2.75
X3 VDD1.t8 VP.t1 VTAIL.t12 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=2.9601 ps=15.96 w=7.59 l=2.75
X4 VTAIL.t6 VN.t0 VDD2.t9 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X5 VDD1.t7 VP.t2 VTAIL.t19 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X6 VTAIL.t13 VP.t3 VDD1.t6 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X7 VDD2.t8 VN.t1 VTAIL.t1 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X8 VDD2.t7 VN.t2 VTAIL.t5 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=2.9601 ps=15.96 w=7.59 l=2.75
X9 VTAIL.t14 VP.t4 VDD1.t5 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X10 VTAIL.t9 VN.t3 VDD2.t6 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X11 VTAIL.t0 VN.t4 VDD2.t5 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X12 VDD2.t4 VN.t5 VTAIL.t4 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=1.25235 ps=7.92 w=7.59 l=2.75
X13 VTAIL.t15 VP.t5 VDD1.t4 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X14 VDD2.t3 VN.t6 VTAIL.t7 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X15 VDD2.t2 VN.t7 VTAIL.t2 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=1.25235 ps=7.92 w=7.59 l=2.75
X16 VDD1.t3 VP.t6 VTAIL.t16 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=1.25235 ps=7.92 w=7.59 l=2.75
X17 VTAIL.t8 VN.t8 VDD2.t1 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X18 VDD1.t2 VP.t7 VTAIL.t11 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X19 VDD2.t0 VN.t9 VTAIL.t3 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=2.9601 ps=15.96 w=7.59 l=2.75
X20 VTAIL.t17 VP.t8 VDD1.t1 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=1.25235 ps=7.92 w=7.59 l=2.75
X21 B.t5 B.t3 B.t4 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=0 ps=0 w=7.59 l=2.75
X22 B.t2 B.t0 B.t1 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=2.9601 pd=15.96 as=0 ps=0 w=7.59 l=2.75
X23 VDD1.t0 VP.t9 VTAIL.t18 w_n4666_n2486# sky130_fd_pr__pfet_01v8 ad=1.25235 pd=7.92 as=2.9601 ps=15.96 w=7.59 l=2.75
R0 B.n395 B.n134 585
R1 B.n394 B.n393 585
R2 B.n392 B.n135 585
R3 B.n391 B.n390 585
R4 B.n389 B.n136 585
R5 B.n388 B.n387 585
R6 B.n386 B.n137 585
R7 B.n385 B.n384 585
R8 B.n383 B.n138 585
R9 B.n382 B.n381 585
R10 B.n380 B.n139 585
R11 B.n379 B.n378 585
R12 B.n377 B.n140 585
R13 B.n376 B.n375 585
R14 B.n374 B.n141 585
R15 B.n373 B.n372 585
R16 B.n371 B.n142 585
R17 B.n370 B.n369 585
R18 B.n368 B.n143 585
R19 B.n367 B.n366 585
R20 B.n365 B.n144 585
R21 B.n364 B.n363 585
R22 B.n362 B.n145 585
R23 B.n361 B.n360 585
R24 B.n359 B.n146 585
R25 B.n358 B.n357 585
R26 B.n356 B.n147 585
R27 B.n355 B.n354 585
R28 B.n353 B.n148 585
R29 B.n352 B.n351 585
R30 B.n347 B.n149 585
R31 B.n346 B.n345 585
R32 B.n344 B.n150 585
R33 B.n343 B.n342 585
R34 B.n341 B.n151 585
R35 B.n340 B.n339 585
R36 B.n338 B.n152 585
R37 B.n337 B.n336 585
R38 B.n334 B.n153 585
R39 B.n333 B.n332 585
R40 B.n331 B.n156 585
R41 B.n330 B.n329 585
R42 B.n328 B.n157 585
R43 B.n327 B.n326 585
R44 B.n325 B.n158 585
R45 B.n324 B.n323 585
R46 B.n322 B.n159 585
R47 B.n321 B.n320 585
R48 B.n319 B.n160 585
R49 B.n318 B.n317 585
R50 B.n316 B.n161 585
R51 B.n315 B.n314 585
R52 B.n313 B.n162 585
R53 B.n312 B.n311 585
R54 B.n310 B.n163 585
R55 B.n309 B.n308 585
R56 B.n307 B.n164 585
R57 B.n306 B.n305 585
R58 B.n304 B.n165 585
R59 B.n303 B.n302 585
R60 B.n301 B.n166 585
R61 B.n300 B.n299 585
R62 B.n298 B.n167 585
R63 B.n297 B.n296 585
R64 B.n295 B.n168 585
R65 B.n294 B.n293 585
R66 B.n292 B.n169 585
R67 B.n397 B.n396 585
R68 B.n398 B.n133 585
R69 B.n400 B.n399 585
R70 B.n401 B.n132 585
R71 B.n403 B.n402 585
R72 B.n404 B.n131 585
R73 B.n406 B.n405 585
R74 B.n407 B.n130 585
R75 B.n409 B.n408 585
R76 B.n410 B.n129 585
R77 B.n412 B.n411 585
R78 B.n413 B.n128 585
R79 B.n415 B.n414 585
R80 B.n416 B.n127 585
R81 B.n418 B.n417 585
R82 B.n419 B.n126 585
R83 B.n421 B.n420 585
R84 B.n422 B.n125 585
R85 B.n424 B.n423 585
R86 B.n425 B.n124 585
R87 B.n427 B.n426 585
R88 B.n428 B.n123 585
R89 B.n430 B.n429 585
R90 B.n431 B.n122 585
R91 B.n433 B.n432 585
R92 B.n434 B.n121 585
R93 B.n436 B.n435 585
R94 B.n437 B.n120 585
R95 B.n439 B.n438 585
R96 B.n440 B.n119 585
R97 B.n442 B.n441 585
R98 B.n443 B.n118 585
R99 B.n445 B.n444 585
R100 B.n446 B.n117 585
R101 B.n448 B.n447 585
R102 B.n449 B.n116 585
R103 B.n451 B.n450 585
R104 B.n452 B.n115 585
R105 B.n454 B.n453 585
R106 B.n455 B.n114 585
R107 B.n457 B.n456 585
R108 B.n458 B.n113 585
R109 B.n460 B.n459 585
R110 B.n461 B.n112 585
R111 B.n463 B.n462 585
R112 B.n464 B.n111 585
R113 B.n466 B.n465 585
R114 B.n467 B.n110 585
R115 B.n469 B.n468 585
R116 B.n470 B.n109 585
R117 B.n472 B.n471 585
R118 B.n473 B.n108 585
R119 B.n475 B.n474 585
R120 B.n476 B.n107 585
R121 B.n478 B.n477 585
R122 B.n479 B.n106 585
R123 B.n481 B.n480 585
R124 B.n482 B.n105 585
R125 B.n484 B.n483 585
R126 B.n485 B.n104 585
R127 B.n487 B.n486 585
R128 B.n488 B.n103 585
R129 B.n490 B.n489 585
R130 B.n491 B.n102 585
R131 B.n493 B.n492 585
R132 B.n494 B.n101 585
R133 B.n496 B.n495 585
R134 B.n497 B.n100 585
R135 B.n499 B.n498 585
R136 B.n500 B.n99 585
R137 B.n502 B.n501 585
R138 B.n503 B.n98 585
R139 B.n505 B.n504 585
R140 B.n506 B.n97 585
R141 B.n508 B.n507 585
R142 B.n509 B.n96 585
R143 B.n511 B.n510 585
R144 B.n512 B.n95 585
R145 B.n514 B.n513 585
R146 B.n515 B.n94 585
R147 B.n517 B.n516 585
R148 B.n518 B.n93 585
R149 B.n520 B.n519 585
R150 B.n521 B.n92 585
R151 B.n523 B.n522 585
R152 B.n524 B.n91 585
R153 B.n526 B.n525 585
R154 B.n527 B.n90 585
R155 B.n529 B.n528 585
R156 B.n530 B.n89 585
R157 B.n532 B.n531 585
R158 B.n533 B.n88 585
R159 B.n535 B.n534 585
R160 B.n536 B.n87 585
R161 B.n538 B.n537 585
R162 B.n539 B.n86 585
R163 B.n541 B.n540 585
R164 B.n542 B.n85 585
R165 B.n544 B.n543 585
R166 B.n545 B.n84 585
R167 B.n547 B.n546 585
R168 B.n548 B.n83 585
R169 B.n550 B.n549 585
R170 B.n551 B.n82 585
R171 B.n553 B.n552 585
R172 B.n554 B.n81 585
R173 B.n556 B.n555 585
R174 B.n557 B.n80 585
R175 B.n559 B.n558 585
R176 B.n560 B.n79 585
R177 B.n562 B.n561 585
R178 B.n563 B.n78 585
R179 B.n565 B.n564 585
R180 B.n566 B.n77 585
R181 B.n568 B.n567 585
R182 B.n569 B.n76 585
R183 B.n571 B.n570 585
R184 B.n572 B.n75 585
R185 B.n574 B.n573 585
R186 B.n575 B.n74 585
R187 B.n577 B.n576 585
R188 B.n578 B.n73 585
R189 B.n580 B.n579 585
R190 B.n581 B.n72 585
R191 B.n583 B.n582 585
R192 B.n584 B.n71 585
R193 B.n686 B.n33 585
R194 B.n685 B.n684 585
R195 B.n683 B.n34 585
R196 B.n682 B.n681 585
R197 B.n680 B.n35 585
R198 B.n679 B.n678 585
R199 B.n677 B.n36 585
R200 B.n676 B.n675 585
R201 B.n674 B.n37 585
R202 B.n673 B.n672 585
R203 B.n671 B.n38 585
R204 B.n670 B.n669 585
R205 B.n668 B.n39 585
R206 B.n667 B.n666 585
R207 B.n665 B.n40 585
R208 B.n664 B.n663 585
R209 B.n662 B.n41 585
R210 B.n661 B.n660 585
R211 B.n659 B.n42 585
R212 B.n658 B.n657 585
R213 B.n656 B.n43 585
R214 B.n655 B.n654 585
R215 B.n653 B.n44 585
R216 B.n652 B.n651 585
R217 B.n650 B.n45 585
R218 B.n649 B.n648 585
R219 B.n647 B.n46 585
R220 B.n646 B.n645 585
R221 B.n644 B.n47 585
R222 B.n642 B.n641 585
R223 B.n640 B.n50 585
R224 B.n639 B.n638 585
R225 B.n637 B.n51 585
R226 B.n636 B.n635 585
R227 B.n634 B.n52 585
R228 B.n633 B.n632 585
R229 B.n631 B.n53 585
R230 B.n630 B.n629 585
R231 B.n628 B.n627 585
R232 B.n626 B.n57 585
R233 B.n625 B.n624 585
R234 B.n623 B.n58 585
R235 B.n622 B.n621 585
R236 B.n620 B.n59 585
R237 B.n619 B.n618 585
R238 B.n617 B.n60 585
R239 B.n616 B.n615 585
R240 B.n614 B.n61 585
R241 B.n613 B.n612 585
R242 B.n611 B.n62 585
R243 B.n610 B.n609 585
R244 B.n608 B.n63 585
R245 B.n607 B.n606 585
R246 B.n605 B.n64 585
R247 B.n604 B.n603 585
R248 B.n602 B.n65 585
R249 B.n601 B.n600 585
R250 B.n599 B.n66 585
R251 B.n598 B.n597 585
R252 B.n596 B.n67 585
R253 B.n595 B.n594 585
R254 B.n593 B.n68 585
R255 B.n592 B.n591 585
R256 B.n590 B.n69 585
R257 B.n589 B.n588 585
R258 B.n587 B.n70 585
R259 B.n586 B.n585 585
R260 B.n688 B.n687 585
R261 B.n689 B.n32 585
R262 B.n691 B.n690 585
R263 B.n692 B.n31 585
R264 B.n694 B.n693 585
R265 B.n695 B.n30 585
R266 B.n697 B.n696 585
R267 B.n698 B.n29 585
R268 B.n700 B.n699 585
R269 B.n701 B.n28 585
R270 B.n703 B.n702 585
R271 B.n704 B.n27 585
R272 B.n706 B.n705 585
R273 B.n707 B.n26 585
R274 B.n709 B.n708 585
R275 B.n710 B.n25 585
R276 B.n712 B.n711 585
R277 B.n713 B.n24 585
R278 B.n715 B.n714 585
R279 B.n716 B.n23 585
R280 B.n718 B.n717 585
R281 B.n719 B.n22 585
R282 B.n721 B.n720 585
R283 B.n722 B.n21 585
R284 B.n724 B.n723 585
R285 B.n725 B.n20 585
R286 B.n727 B.n726 585
R287 B.n728 B.n19 585
R288 B.n730 B.n729 585
R289 B.n731 B.n18 585
R290 B.n733 B.n732 585
R291 B.n734 B.n17 585
R292 B.n736 B.n735 585
R293 B.n737 B.n16 585
R294 B.n739 B.n738 585
R295 B.n740 B.n15 585
R296 B.n742 B.n741 585
R297 B.n743 B.n14 585
R298 B.n745 B.n744 585
R299 B.n746 B.n13 585
R300 B.n748 B.n747 585
R301 B.n749 B.n12 585
R302 B.n751 B.n750 585
R303 B.n752 B.n11 585
R304 B.n754 B.n753 585
R305 B.n755 B.n10 585
R306 B.n757 B.n756 585
R307 B.n758 B.n9 585
R308 B.n760 B.n759 585
R309 B.n761 B.n8 585
R310 B.n763 B.n762 585
R311 B.n764 B.n7 585
R312 B.n766 B.n765 585
R313 B.n767 B.n6 585
R314 B.n769 B.n768 585
R315 B.n770 B.n5 585
R316 B.n772 B.n771 585
R317 B.n773 B.n4 585
R318 B.n775 B.n774 585
R319 B.n776 B.n3 585
R320 B.n778 B.n777 585
R321 B.n779 B.n0 585
R322 B.n2 B.n1 585
R323 B.n201 B.n200 585
R324 B.n202 B.n199 585
R325 B.n204 B.n203 585
R326 B.n205 B.n198 585
R327 B.n207 B.n206 585
R328 B.n208 B.n197 585
R329 B.n210 B.n209 585
R330 B.n211 B.n196 585
R331 B.n213 B.n212 585
R332 B.n214 B.n195 585
R333 B.n216 B.n215 585
R334 B.n217 B.n194 585
R335 B.n219 B.n218 585
R336 B.n220 B.n193 585
R337 B.n222 B.n221 585
R338 B.n223 B.n192 585
R339 B.n225 B.n224 585
R340 B.n226 B.n191 585
R341 B.n228 B.n227 585
R342 B.n229 B.n190 585
R343 B.n231 B.n230 585
R344 B.n232 B.n189 585
R345 B.n234 B.n233 585
R346 B.n235 B.n188 585
R347 B.n237 B.n236 585
R348 B.n238 B.n187 585
R349 B.n240 B.n239 585
R350 B.n241 B.n186 585
R351 B.n243 B.n242 585
R352 B.n244 B.n185 585
R353 B.n246 B.n245 585
R354 B.n247 B.n184 585
R355 B.n249 B.n248 585
R356 B.n250 B.n183 585
R357 B.n252 B.n251 585
R358 B.n253 B.n182 585
R359 B.n255 B.n254 585
R360 B.n256 B.n181 585
R361 B.n258 B.n257 585
R362 B.n259 B.n180 585
R363 B.n261 B.n260 585
R364 B.n262 B.n179 585
R365 B.n264 B.n263 585
R366 B.n265 B.n178 585
R367 B.n267 B.n266 585
R368 B.n268 B.n177 585
R369 B.n270 B.n269 585
R370 B.n271 B.n176 585
R371 B.n273 B.n272 585
R372 B.n274 B.n175 585
R373 B.n276 B.n275 585
R374 B.n277 B.n174 585
R375 B.n279 B.n278 585
R376 B.n280 B.n173 585
R377 B.n282 B.n281 585
R378 B.n283 B.n172 585
R379 B.n285 B.n284 585
R380 B.n286 B.n171 585
R381 B.n288 B.n287 585
R382 B.n289 B.n170 585
R383 B.n291 B.n290 585
R384 B.n290 B.n169 482.89
R385 B.n396 B.n395 482.89
R386 B.n586 B.n71 482.89
R387 B.n688 B.n33 482.89
R388 B.n154 B.t3 274.779
R389 B.n348 B.t6 274.779
R390 B.n54 B.t9 274.779
R391 B.n48 B.t0 274.779
R392 B.n781 B.n780 256.663
R393 B.n780 B.n779 235.042
R394 B.n780 B.n2 235.042
R395 B.n348 B.t7 170.857
R396 B.n54 B.t11 170.857
R397 B.n154 B.t4 170.849
R398 B.n48 B.t2 170.849
R399 B.n294 B.n169 163.367
R400 B.n295 B.n294 163.367
R401 B.n296 B.n295 163.367
R402 B.n296 B.n167 163.367
R403 B.n300 B.n167 163.367
R404 B.n301 B.n300 163.367
R405 B.n302 B.n301 163.367
R406 B.n302 B.n165 163.367
R407 B.n306 B.n165 163.367
R408 B.n307 B.n306 163.367
R409 B.n308 B.n307 163.367
R410 B.n308 B.n163 163.367
R411 B.n312 B.n163 163.367
R412 B.n313 B.n312 163.367
R413 B.n314 B.n313 163.367
R414 B.n314 B.n161 163.367
R415 B.n318 B.n161 163.367
R416 B.n319 B.n318 163.367
R417 B.n320 B.n319 163.367
R418 B.n320 B.n159 163.367
R419 B.n324 B.n159 163.367
R420 B.n325 B.n324 163.367
R421 B.n326 B.n325 163.367
R422 B.n326 B.n157 163.367
R423 B.n330 B.n157 163.367
R424 B.n331 B.n330 163.367
R425 B.n332 B.n331 163.367
R426 B.n332 B.n153 163.367
R427 B.n337 B.n153 163.367
R428 B.n338 B.n337 163.367
R429 B.n339 B.n338 163.367
R430 B.n339 B.n151 163.367
R431 B.n343 B.n151 163.367
R432 B.n344 B.n343 163.367
R433 B.n345 B.n344 163.367
R434 B.n345 B.n149 163.367
R435 B.n352 B.n149 163.367
R436 B.n353 B.n352 163.367
R437 B.n354 B.n353 163.367
R438 B.n354 B.n147 163.367
R439 B.n358 B.n147 163.367
R440 B.n359 B.n358 163.367
R441 B.n360 B.n359 163.367
R442 B.n360 B.n145 163.367
R443 B.n364 B.n145 163.367
R444 B.n365 B.n364 163.367
R445 B.n366 B.n365 163.367
R446 B.n366 B.n143 163.367
R447 B.n370 B.n143 163.367
R448 B.n371 B.n370 163.367
R449 B.n372 B.n371 163.367
R450 B.n372 B.n141 163.367
R451 B.n376 B.n141 163.367
R452 B.n377 B.n376 163.367
R453 B.n378 B.n377 163.367
R454 B.n378 B.n139 163.367
R455 B.n382 B.n139 163.367
R456 B.n383 B.n382 163.367
R457 B.n384 B.n383 163.367
R458 B.n384 B.n137 163.367
R459 B.n388 B.n137 163.367
R460 B.n389 B.n388 163.367
R461 B.n390 B.n389 163.367
R462 B.n390 B.n135 163.367
R463 B.n394 B.n135 163.367
R464 B.n395 B.n394 163.367
R465 B.n582 B.n71 163.367
R466 B.n582 B.n581 163.367
R467 B.n581 B.n580 163.367
R468 B.n580 B.n73 163.367
R469 B.n576 B.n73 163.367
R470 B.n576 B.n575 163.367
R471 B.n575 B.n574 163.367
R472 B.n574 B.n75 163.367
R473 B.n570 B.n75 163.367
R474 B.n570 B.n569 163.367
R475 B.n569 B.n568 163.367
R476 B.n568 B.n77 163.367
R477 B.n564 B.n77 163.367
R478 B.n564 B.n563 163.367
R479 B.n563 B.n562 163.367
R480 B.n562 B.n79 163.367
R481 B.n558 B.n79 163.367
R482 B.n558 B.n557 163.367
R483 B.n557 B.n556 163.367
R484 B.n556 B.n81 163.367
R485 B.n552 B.n81 163.367
R486 B.n552 B.n551 163.367
R487 B.n551 B.n550 163.367
R488 B.n550 B.n83 163.367
R489 B.n546 B.n83 163.367
R490 B.n546 B.n545 163.367
R491 B.n545 B.n544 163.367
R492 B.n544 B.n85 163.367
R493 B.n540 B.n85 163.367
R494 B.n540 B.n539 163.367
R495 B.n539 B.n538 163.367
R496 B.n538 B.n87 163.367
R497 B.n534 B.n87 163.367
R498 B.n534 B.n533 163.367
R499 B.n533 B.n532 163.367
R500 B.n532 B.n89 163.367
R501 B.n528 B.n89 163.367
R502 B.n528 B.n527 163.367
R503 B.n527 B.n526 163.367
R504 B.n526 B.n91 163.367
R505 B.n522 B.n91 163.367
R506 B.n522 B.n521 163.367
R507 B.n521 B.n520 163.367
R508 B.n520 B.n93 163.367
R509 B.n516 B.n93 163.367
R510 B.n516 B.n515 163.367
R511 B.n515 B.n514 163.367
R512 B.n514 B.n95 163.367
R513 B.n510 B.n95 163.367
R514 B.n510 B.n509 163.367
R515 B.n509 B.n508 163.367
R516 B.n508 B.n97 163.367
R517 B.n504 B.n97 163.367
R518 B.n504 B.n503 163.367
R519 B.n503 B.n502 163.367
R520 B.n502 B.n99 163.367
R521 B.n498 B.n99 163.367
R522 B.n498 B.n497 163.367
R523 B.n497 B.n496 163.367
R524 B.n496 B.n101 163.367
R525 B.n492 B.n101 163.367
R526 B.n492 B.n491 163.367
R527 B.n491 B.n490 163.367
R528 B.n490 B.n103 163.367
R529 B.n486 B.n103 163.367
R530 B.n486 B.n485 163.367
R531 B.n485 B.n484 163.367
R532 B.n484 B.n105 163.367
R533 B.n480 B.n105 163.367
R534 B.n480 B.n479 163.367
R535 B.n479 B.n478 163.367
R536 B.n478 B.n107 163.367
R537 B.n474 B.n107 163.367
R538 B.n474 B.n473 163.367
R539 B.n473 B.n472 163.367
R540 B.n472 B.n109 163.367
R541 B.n468 B.n109 163.367
R542 B.n468 B.n467 163.367
R543 B.n467 B.n466 163.367
R544 B.n466 B.n111 163.367
R545 B.n462 B.n111 163.367
R546 B.n462 B.n461 163.367
R547 B.n461 B.n460 163.367
R548 B.n460 B.n113 163.367
R549 B.n456 B.n113 163.367
R550 B.n456 B.n455 163.367
R551 B.n455 B.n454 163.367
R552 B.n454 B.n115 163.367
R553 B.n450 B.n115 163.367
R554 B.n450 B.n449 163.367
R555 B.n449 B.n448 163.367
R556 B.n448 B.n117 163.367
R557 B.n444 B.n117 163.367
R558 B.n444 B.n443 163.367
R559 B.n443 B.n442 163.367
R560 B.n442 B.n119 163.367
R561 B.n438 B.n119 163.367
R562 B.n438 B.n437 163.367
R563 B.n437 B.n436 163.367
R564 B.n436 B.n121 163.367
R565 B.n432 B.n121 163.367
R566 B.n432 B.n431 163.367
R567 B.n431 B.n430 163.367
R568 B.n430 B.n123 163.367
R569 B.n426 B.n123 163.367
R570 B.n426 B.n425 163.367
R571 B.n425 B.n424 163.367
R572 B.n424 B.n125 163.367
R573 B.n420 B.n125 163.367
R574 B.n420 B.n419 163.367
R575 B.n419 B.n418 163.367
R576 B.n418 B.n127 163.367
R577 B.n414 B.n127 163.367
R578 B.n414 B.n413 163.367
R579 B.n413 B.n412 163.367
R580 B.n412 B.n129 163.367
R581 B.n408 B.n129 163.367
R582 B.n408 B.n407 163.367
R583 B.n407 B.n406 163.367
R584 B.n406 B.n131 163.367
R585 B.n402 B.n131 163.367
R586 B.n402 B.n401 163.367
R587 B.n401 B.n400 163.367
R588 B.n400 B.n133 163.367
R589 B.n396 B.n133 163.367
R590 B.n684 B.n33 163.367
R591 B.n684 B.n683 163.367
R592 B.n683 B.n682 163.367
R593 B.n682 B.n35 163.367
R594 B.n678 B.n35 163.367
R595 B.n678 B.n677 163.367
R596 B.n677 B.n676 163.367
R597 B.n676 B.n37 163.367
R598 B.n672 B.n37 163.367
R599 B.n672 B.n671 163.367
R600 B.n671 B.n670 163.367
R601 B.n670 B.n39 163.367
R602 B.n666 B.n39 163.367
R603 B.n666 B.n665 163.367
R604 B.n665 B.n664 163.367
R605 B.n664 B.n41 163.367
R606 B.n660 B.n41 163.367
R607 B.n660 B.n659 163.367
R608 B.n659 B.n658 163.367
R609 B.n658 B.n43 163.367
R610 B.n654 B.n43 163.367
R611 B.n654 B.n653 163.367
R612 B.n653 B.n652 163.367
R613 B.n652 B.n45 163.367
R614 B.n648 B.n45 163.367
R615 B.n648 B.n647 163.367
R616 B.n647 B.n646 163.367
R617 B.n646 B.n47 163.367
R618 B.n641 B.n47 163.367
R619 B.n641 B.n640 163.367
R620 B.n640 B.n639 163.367
R621 B.n639 B.n51 163.367
R622 B.n635 B.n51 163.367
R623 B.n635 B.n634 163.367
R624 B.n634 B.n633 163.367
R625 B.n633 B.n53 163.367
R626 B.n629 B.n53 163.367
R627 B.n629 B.n628 163.367
R628 B.n628 B.n57 163.367
R629 B.n624 B.n57 163.367
R630 B.n624 B.n623 163.367
R631 B.n623 B.n622 163.367
R632 B.n622 B.n59 163.367
R633 B.n618 B.n59 163.367
R634 B.n618 B.n617 163.367
R635 B.n617 B.n616 163.367
R636 B.n616 B.n61 163.367
R637 B.n612 B.n61 163.367
R638 B.n612 B.n611 163.367
R639 B.n611 B.n610 163.367
R640 B.n610 B.n63 163.367
R641 B.n606 B.n63 163.367
R642 B.n606 B.n605 163.367
R643 B.n605 B.n604 163.367
R644 B.n604 B.n65 163.367
R645 B.n600 B.n65 163.367
R646 B.n600 B.n599 163.367
R647 B.n599 B.n598 163.367
R648 B.n598 B.n67 163.367
R649 B.n594 B.n67 163.367
R650 B.n594 B.n593 163.367
R651 B.n593 B.n592 163.367
R652 B.n592 B.n69 163.367
R653 B.n588 B.n69 163.367
R654 B.n588 B.n587 163.367
R655 B.n587 B.n586 163.367
R656 B.n689 B.n688 163.367
R657 B.n690 B.n689 163.367
R658 B.n690 B.n31 163.367
R659 B.n694 B.n31 163.367
R660 B.n695 B.n694 163.367
R661 B.n696 B.n695 163.367
R662 B.n696 B.n29 163.367
R663 B.n700 B.n29 163.367
R664 B.n701 B.n700 163.367
R665 B.n702 B.n701 163.367
R666 B.n702 B.n27 163.367
R667 B.n706 B.n27 163.367
R668 B.n707 B.n706 163.367
R669 B.n708 B.n707 163.367
R670 B.n708 B.n25 163.367
R671 B.n712 B.n25 163.367
R672 B.n713 B.n712 163.367
R673 B.n714 B.n713 163.367
R674 B.n714 B.n23 163.367
R675 B.n718 B.n23 163.367
R676 B.n719 B.n718 163.367
R677 B.n720 B.n719 163.367
R678 B.n720 B.n21 163.367
R679 B.n724 B.n21 163.367
R680 B.n725 B.n724 163.367
R681 B.n726 B.n725 163.367
R682 B.n726 B.n19 163.367
R683 B.n730 B.n19 163.367
R684 B.n731 B.n730 163.367
R685 B.n732 B.n731 163.367
R686 B.n732 B.n17 163.367
R687 B.n736 B.n17 163.367
R688 B.n737 B.n736 163.367
R689 B.n738 B.n737 163.367
R690 B.n738 B.n15 163.367
R691 B.n742 B.n15 163.367
R692 B.n743 B.n742 163.367
R693 B.n744 B.n743 163.367
R694 B.n744 B.n13 163.367
R695 B.n748 B.n13 163.367
R696 B.n749 B.n748 163.367
R697 B.n750 B.n749 163.367
R698 B.n750 B.n11 163.367
R699 B.n754 B.n11 163.367
R700 B.n755 B.n754 163.367
R701 B.n756 B.n755 163.367
R702 B.n756 B.n9 163.367
R703 B.n760 B.n9 163.367
R704 B.n761 B.n760 163.367
R705 B.n762 B.n761 163.367
R706 B.n762 B.n7 163.367
R707 B.n766 B.n7 163.367
R708 B.n767 B.n766 163.367
R709 B.n768 B.n767 163.367
R710 B.n768 B.n5 163.367
R711 B.n772 B.n5 163.367
R712 B.n773 B.n772 163.367
R713 B.n774 B.n773 163.367
R714 B.n774 B.n3 163.367
R715 B.n778 B.n3 163.367
R716 B.n779 B.n778 163.367
R717 B.n200 B.n2 163.367
R718 B.n200 B.n199 163.367
R719 B.n204 B.n199 163.367
R720 B.n205 B.n204 163.367
R721 B.n206 B.n205 163.367
R722 B.n206 B.n197 163.367
R723 B.n210 B.n197 163.367
R724 B.n211 B.n210 163.367
R725 B.n212 B.n211 163.367
R726 B.n212 B.n195 163.367
R727 B.n216 B.n195 163.367
R728 B.n217 B.n216 163.367
R729 B.n218 B.n217 163.367
R730 B.n218 B.n193 163.367
R731 B.n222 B.n193 163.367
R732 B.n223 B.n222 163.367
R733 B.n224 B.n223 163.367
R734 B.n224 B.n191 163.367
R735 B.n228 B.n191 163.367
R736 B.n229 B.n228 163.367
R737 B.n230 B.n229 163.367
R738 B.n230 B.n189 163.367
R739 B.n234 B.n189 163.367
R740 B.n235 B.n234 163.367
R741 B.n236 B.n235 163.367
R742 B.n236 B.n187 163.367
R743 B.n240 B.n187 163.367
R744 B.n241 B.n240 163.367
R745 B.n242 B.n241 163.367
R746 B.n242 B.n185 163.367
R747 B.n246 B.n185 163.367
R748 B.n247 B.n246 163.367
R749 B.n248 B.n247 163.367
R750 B.n248 B.n183 163.367
R751 B.n252 B.n183 163.367
R752 B.n253 B.n252 163.367
R753 B.n254 B.n253 163.367
R754 B.n254 B.n181 163.367
R755 B.n258 B.n181 163.367
R756 B.n259 B.n258 163.367
R757 B.n260 B.n259 163.367
R758 B.n260 B.n179 163.367
R759 B.n264 B.n179 163.367
R760 B.n265 B.n264 163.367
R761 B.n266 B.n265 163.367
R762 B.n266 B.n177 163.367
R763 B.n270 B.n177 163.367
R764 B.n271 B.n270 163.367
R765 B.n272 B.n271 163.367
R766 B.n272 B.n175 163.367
R767 B.n276 B.n175 163.367
R768 B.n277 B.n276 163.367
R769 B.n278 B.n277 163.367
R770 B.n278 B.n173 163.367
R771 B.n282 B.n173 163.367
R772 B.n283 B.n282 163.367
R773 B.n284 B.n283 163.367
R774 B.n284 B.n171 163.367
R775 B.n288 B.n171 163.367
R776 B.n289 B.n288 163.367
R777 B.n290 B.n289 163.367
R778 B.n349 B.t8 111.124
R779 B.n55 B.t10 111.124
R780 B.n155 B.t5 111.115
R781 B.n49 B.t1 111.115
R782 B.n155 B.n154 59.7338
R783 B.n349 B.n348 59.7338
R784 B.n55 B.n54 59.7338
R785 B.n49 B.n48 59.7338
R786 B.n335 B.n155 59.5399
R787 B.n350 B.n349 59.5399
R788 B.n56 B.n55 59.5399
R789 B.n643 B.n49 59.5399
R790 B.n687 B.n686 31.3761
R791 B.n585 B.n584 31.3761
R792 B.n397 B.n134 31.3761
R793 B.n292 B.n291 31.3761
R794 B B.n781 18.0485
R795 B.n687 B.n32 10.6151
R796 B.n691 B.n32 10.6151
R797 B.n692 B.n691 10.6151
R798 B.n693 B.n692 10.6151
R799 B.n693 B.n30 10.6151
R800 B.n697 B.n30 10.6151
R801 B.n698 B.n697 10.6151
R802 B.n699 B.n698 10.6151
R803 B.n699 B.n28 10.6151
R804 B.n703 B.n28 10.6151
R805 B.n704 B.n703 10.6151
R806 B.n705 B.n704 10.6151
R807 B.n705 B.n26 10.6151
R808 B.n709 B.n26 10.6151
R809 B.n710 B.n709 10.6151
R810 B.n711 B.n710 10.6151
R811 B.n711 B.n24 10.6151
R812 B.n715 B.n24 10.6151
R813 B.n716 B.n715 10.6151
R814 B.n717 B.n716 10.6151
R815 B.n717 B.n22 10.6151
R816 B.n721 B.n22 10.6151
R817 B.n722 B.n721 10.6151
R818 B.n723 B.n722 10.6151
R819 B.n723 B.n20 10.6151
R820 B.n727 B.n20 10.6151
R821 B.n728 B.n727 10.6151
R822 B.n729 B.n728 10.6151
R823 B.n729 B.n18 10.6151
R824 B.n733 B.n18 10.6151
R825 B.n734 B.n733 10.6151
R826 B.n735 B.n734 10.6151
R827 B.n735 B.n16 10.6151
R828 B.n739 B.n16 10.6151
R829 B.n740 B.n739 10.6151
R830 B.n741 B.n740 10.6151
R831 B.n741 B.n14 10.6151
R832 B.n745 B.n14 10.6151
R833 B.n746 B.n745 10.6151
R834 B.n747 B.n746 10.6151
R835 B.n747 B.n12 10.6151
R836 B.n751 B.n12 10.6151
R837 B.n752 B.n751 10.6151
R838 B.n753 B.n752 10.6151
R839 B.n753 B.n10 10.6151
R840 B.n757 B.n10 10.6151
R841 B.n758 B.n757 10.6151
R842 B.n759 B.n758 10.6151
R843 B.n759 B.n8 10.6151
R844 B.n763 B.n8 10.6151
R845 B.n764 B.n763 10.6151
R846 B.n765 B.n764 10.6151
R847 B.n765 B.n6 10.6151
R848 B.n769 B.n6 10.6151
R849 B.n770 B.n769 10.6151
R850 B.n771 B.n770 10.6151
R851 B.n771 B.n4 10.6151
R852 B.n775 B.n4 10.6151
R853 B.n776 B.n775 10.6151
R854 B.n777 B.n776 10.6151
R855 B.n777 B.n0 10.6151
R856 B.n686 B.n685 10.6151
R857 B.n685 B.n34 10.6151
R858 B.n681 B.n34 10.6151
R859 B.n681 B.n680 10.6151
R860 B.n680 B.n679 10.6151
R861 B.n679 B.n36 10.6151
R862 B.n675 B.n36 10.6151
R863 B.n675 B.n674 10.6151
R864 B.n674 B.n673 10.6151
R865 B.n673 B.n38 10.6151
R866 B.n669 B.n38 10.6151
R867 B.n669 B.n668 10.6151
R868 B.n668 B.n667 10.6151
R869 B.n667 B.n40 10.6151
R870 B.n663 B.n40 10.6151
R871 B.n663 B.n662 10.6151
R872 B.n662 B.n661 10.6151
R873 B.n661 B.n42 10.6151
R874 B.n657 B.n42 10.6151
R875 B.n657 B.n656 10.6151
R876 B.n656 B.n655 10.6151
R877 B.n655 B.n44 10.6151
R878 B.n651 B.n44 10.6151
R879 B.n651 B.n650 10.6151
R880 B.n650 B.n649 10.6151
R881 B.n649 B.n46 10.6151
R882 B.n645 B.n46 10.6151
R883 B.n645 B.n644 10.6151
R884 B.n642 B.n50 10.6151
R885 B.n638 B.n50 10.6151
R886 B.n638 B.n637 10.6151
R887 B.n637 B.n636 10.6151
R888 B.n636 B.n52 10.6151
R889 B.n632 B.n52 10.6151
R890 B.n632 B.n631 10.6151
R891 B.n631 B.n630 10.6151
R892 B.n627 B.n626 10.6151
R893 B.n626 B.n625 10.6151
R894 B.n625 B.n58 10.6151
R895 B.n621 B.n58 10.6151
R896 B.n621 B.n620 10.6151
R897 B.n620 B.n619 10.6151
R898 B.n619 B.n60 10.6151
R899 B.n615 B.n60 10.6151
R900 B.n615 B.n614 10.6151
R901 B.n614 B.n613 10.6151
R902 B.n613 B.n62 10.6151
R903 B.n609 B.n62 10.6151
R904 B.n609 B.n608 10.6151
R905 B.n608 B.n607 10.6151
R906 B.n607 B.n64 10.6151
R907 B.n603 B.n64 10.6151
R908 B.n603 B.n602 10.6151
R909 B.n602 B.n601 10.6151
R910 B.n601 B.n66 10.6151
R911 B.n597 B.n66 10.6151
R912 B.n597 B.n596 10.6151
R913 B.n596 B.n595 10.6151
R914 B.n595 B.n68 10.6151
R915 B.n591 B.n68 10.6151
R916 B.n591 B.n590 10.6151
R917 B.n590 B.n589 10.6151
R918 B.n589 B.n70 10.6151
R919 B.n585 B.n70 10.6151
R920 B.n584 B.n583 10.6151
R921 B.n583 B.n72 10.6151
R922 B.n579 B.n72 10.6151
R923 B.n579 B.n578 10.6151
R924 B.n578 B.n577 10.6151
R925 B.n577 B.n74 10.6151
R926 B.n573 B.n74 10.6151
R927 B.n573 B.n572 10.6151
R928 B.n572 B.n571 10.6151
R929 B.n571 B.n76 10.6151
R930 B.n567 B.n76 10.6151
R931 B.n567 B.n566 10.6151
R932 B.n566 B.n565 10.6151
R933 B.n565 B.n78 10.6151
R934 B.n561 B.n78 10.6151
R935 B.n561 B.n560 10.6151
R936 B.n560 B.n559 10.6151
R937 B.n559 B.n80 10.6151
R938 B.n555 B.n80 10.6151
R939 B.n555 B.n554 10.6151
R940 B.n554 B.n553 10.6151
R941 B.n553 B.n82 10.6151
R942 B.n549 B.n82 10.6151
R943 B.n549 B.n548 10.6151
R944 B.n548 B.n547 10.6151
R945 B.n547 B.n84 10.6151
R946 B.n543 B.n84 10.6151
R947 B.n543 B.n542 10.6151
R948 B.n542 B.n541 10.6151
R949 B.n541 B.n86 10.6151
R950 B.n537 B.n86 10.6151
R951 B.n537 B.n536 10.6151
R952 B.n536 B.n535 10.6151
R953 B.n535 B.n88 10.6151
R954 B.n531 B.n88 10.6151
R955 B.n531 B.n530 10.6151
R956 B.n530 B.n529 10.6151
R957 B.n529 B.n90 10.6151
R958 B.n525 B.n90 10.6151
R959 B.n525 B.n524 10.6151
R960 B.n524 B.n523 10.6151
R961 B.n523 B.n92 10.6151
R962 B.n519 B.n92 10.6151
R963 B.n519 B.n518 10.6151
R964 B.n518 B.n517 10.6151
R965 B.n517 B.n94 10.6151
R966 B.n513 B.n94 10.6151
R967 B.n513 B.n512 10.6151
R968 B.n512 B.n511 10.6151
R969 B.n511 B.n96 10.6151
R970 B.n507 B.n96 10.6151
R971 B.n507 B.n506 10.6151
R972 B.n506 B.n505 10.6151
R973 B.n505 B.n98 10.6151
R974 B.n501 B.n98 10.6151
R975 B.n501 B.n500 10.6151
R976 B.n500 B.n499 10.6151
R977 B.n499 B.n100 10.6151
R978 B.n495 B.n100 10.6151
R979 B.n495 B.n494 10.6151
R980 B.n494 B.n493 10.6151
R981 B.n493 B.n102 10.6151
R982 B.n489 B.n102 10.6151
R983 B.n489 B.n488 10.6151
R984 B.n488 B.n487 10.6151
R985 B.n487 B.n104 10.6151
R986 B.n483 B.n104 10.6151
R987 B.n483 B.n482 10.6151
R988 B.n482 B.n481 10.6151
R989 B.n481 B.n106 10.6151
R990 B.n477 B.n106 10.6151
R991 B.n477 B.n476 10.6151
R992 B.n476 B.n475 10.6151
R993 B.n475 B.n108 10.6151
R994 B.n471 B.n108 10.6151
R995 B.n471 B.n470 10.6151
R996 B.n470 B.n469 10.6151
R997 B.n469 B.n110 10.6151
R998 B.n465 B.n110 10.6151
R999 B.n465 B.n464 10.6151
R1000 B.n464 B.n463 10.6151
R1001 B.n463 B.n112 10.6151
R1002 B.n459 B.n112 10.6151
R1003 B.n459 B.n458 10.6151
R1004 B.n458 B.n457 10.6151
R1005 B.n457 B.n114 10.6151
R1006 B.n453 B.n114 10.6151
R1007 B.n453 B.n452 10.6151
R1008 B.n452 B.n451 10.6151
R1009 B.n451 B.n116 10.6151
R1010 B.n447 B.n116 10.6151
R1011 B.n447 B.n446 10.6151
R1012 B.n446 B.n445 10.6151
R1013 B.n445 B.n118 10.6151
R1014 B.n441 B.n118 10.6151
R1015 B.n441 B.n440 10.6151
R1016 B.n440 B.n439 10.6151
R1017 B.n439 B.n120 10.6151
R1018 B.n435 B.n120 10.6151
R1019 B.n435 B.n434 10.6151
R1020 B.n434 B.n433 10.6151
R1021 B.n433 B.n122 10.6151
R1022 B.n429 B.n122 10.6151
R1023 B.n429 B.n428 10.6151
R1024 B.n428 B.n427 10.6151
R1025 B.n427 B.n124 10.6151
R1026 B.n423 B.n124 10.6151
R1027 B.n423 B.n422 10.6151
R1028 B.n422 B.n421 10.6151
R1029 B.n421 B.n126 10.6151
R1030 B.n417 B.n126 10.6151
R1031 B.n417 B.n416 10.6151
R1032 B.n416 B.n415 10.6151
R1033 B.n415 B.n128 10.6151
R1034 B.n411 B.n128 10.6151
R1035 B.n411 B.n410 10.6151
R1036 B.n410 B.n409 10.6151
R1037 B.n409 B.n130 10.6151
R1038 B.n405 B.n130 10.6151
R1039 B.n405 B.n404 10.6151
R1040 B.n404 B.n403 10.6151
R1041 B.n403 B.n132 10.6151
R1042 B.n399 B.n132 10.6151
R1043 B.n399 B.n398 10.6151
R1044 B.n398 B.n397 10.6151
R1045 B.n201 B.n1 10.6151
R1046 B.n202 B.n201 10.6151
R1047 B.n203 B.n202 10.6151
R1048 B.n203 B.n198 10.6151
R1049 B.n207 B.n198 10.6151
R1050 B.n208 B.n207 10.6151
R1051 B.n209 B.n208 10.6151
R1052 B.n209 B.n196 10.6151
R1053 B.n213 B.n196 10.6151
R1054 B.n214 B.n213 10.6151
R1055 B.n215 B.n214 10.6151
R1056 B.n215 B.n194 10.6151
R1057 B.n219 B.n194 10.6151
R1058 B.n220 B.n219 10.6151
R1059 B.n221 B.n220 10.6151
R1060 B.n221 B.n192 10.6151
R1061 B.n225 B.n192 10.6151
R1062 B.n226 B.n225 10.6151
R1063 B.n227 B.n226 10.6151
R1064 B.n227 B.n190 10.6151
R1065 B.n231 B.n190 10.6151
R1066 B.n232 B.n231 10.6151
R1067 B.n233 B.n232 10.6151
R1068 B.n233 B.n188 10.6151
R1069 B.n237 B.n188 10.6151
R1070 B.n238 B.n237 10.6151
R1071 B.n239 B.n238 10.6151
R1072 B.n239 B.n186 10.6151
R1073 B.n243 B.n186 10.6151
R1074 B.n244 B.n243 10.6151
R1075 B.n245 B.n244 10.6151
R1076 B.n245 B.n184 10.6151
R1077 B.n249 B.n184 10.6151
R1078 B.n250 B.n249 10.6151
R1079 B.n251 B.n250 10.6151
R1080 B.n251 B.n182 10.6151
R1081 B.n255 B.n182 10.6151
R1082 B.n256 B.n255 10.6151
R1083 B.n257 B.n256 10.6151
R1084 B.n257 B.n180 10.6151
R1085 B.n261 B.n180 10.6151
R1086 B.n262 B.n261 10.6151
R1087 B.n263 B.n262 10.6151
R1088 B.n263 B.n178 10.6151
R1089 B.n267 B.n178 10.6151
R1090 B.n268 B.n267 10.6151
R1091 B.n269 B.n268 10.6151
R1092 B.n269 B.n176 10.6151
R1093 B.n273 B.n176 10.6151
R1094 B.n274 B.n273 10.6151
R1095 B.n275 B.n274 10.6151
R1096 B.n275 B.n174 10.6151
R1097 B.n279 B.n174 10.6151
R1098 B.n280 B.n279 10.6151
R1099 B.n281 B.n280 10.6151
R1100 B.n281 B.n172 10.6151
R1101 B.n285 B.n172 10.6151
R1102 B.n286 B.n285 10.6151
R1103 B.n287 B.n286 10.6151
R1104 B.n287 B.n170 10.6151
R1105 B.n291 B.n170 10.6151
R1106 B.n293 B.n292 10.6151
R1107 B.n293 B.n168 10.6151
R1108 B.n297 B.n168 10.6151
R1109 B.n298 B.n297 10.6151
R1110 B.n299 B.n298 10.6151
R1111 B.n299 B.n166 10.6151
R1112 B.n303 B.n166 10.6151
R1113 B.n304 B.n303 10.6151
R1114 B.n305 B.n304 10.6151
R1115 B.n305 B.n164 10.6151
R1116 B.n309 B.n164 10.6151
R1117 B.n310 B.n309 10.6151
R1118 B.n311 B.n310 10.6151
R1119 B.n311 B.n162 10.6151
R1120 B.n315 B.n162 10.6151
R1121 B.n316 B.n315 10.6151
R1122 B.n317 B.n316 10.6151
R1123 B.n317 B.n160 10.6151
R1124 B.n321 B.n160 10.6151
R1125 B.n322 B.n321 10.6151
R1126 B.n323 B.n322 10.6151
R1127 B.n323 B.n158 10.6151
R1128 B.n327 B.n158 10.6151
R1129 B.n328 B.n327 10.6151
R1130 B.n329 B.n328 10.6151
R1131 B.n329 B.n156 10.6151
R1132 B.n333 B.n156 10.6151
R1133 B.n334 B.n333 10.6151
R1134 B.n336 B.n152 10.6151
R1135 B.n340 B.n152 10.6151
R1136 B.n341 B.n340 10.6151
R1137 B.n342 B.n341 10.6151
R1138 B.n342 B.n150 10.6151
R1139 B.n346 B.n150 10.6151
R1140 B.n347 B.n346 10.6151
R1141 B.n351 B.n347 10.6151
R1142 B.n355 B.n148 10.6151
R1143 B.n356 B.n355 10.6151
R1144 B.n357 B.n356 10.6151
R1145 B.n357 B.n146 10.6151
R1146 B.n361 B.n146 10.6151
R1147 B.n362 B.n361 10.6151
R1148 B.n363 B.n362 10.6151
R1149 B.n363 B.n144 10.6151
R1150 B.n367 B.n144 10.6151
R1151 B.n368 B.n367 10.6151
R1152 B.n369 B.n368 10.6151
R1153 B.n369 B.n142 10.6151
R1154 B.n373 B.n142 10.6151
R1155 B.n374 B.n373 10.6151
R1156 B.n375 B.n374 10.6151
R1157 B.n375 B.n140 10.6151
R1158 B.n379 B.n140 10.6151
R1159 B.n380 B.n379 10.6151
R1160 B.n381 B.n380 10.6151
R1161 B.n381 B.n138 10.6151
R1162 B.n385 B.n138 10.6151
R1163 B.n386 B.n385 10.6151
R1164 B.n387 B.n386 10.6151
R1165 B.n387 B.n136 10.6151
R1166 B.n391 B.n136 10.6151
R1167 B.n392 B.n391 10.6151
R1168 B.n393 B.n392 10.6151
R1169 B.n393 B.n134 10.6151
R1170 B.n781 B.n0 8.11757
R1171 B.n781 B.n1 8.11757
R1172 B.n643 B.n642 6.5566
R1173 B.n630 B.n56 6.5566
R1174 B.n336 B.n335 6.5566
R1175 B.n351 B.n350 6.5566
R1176 B.n644 B.n643 4.05904
R1177 B.n627 B.n56 4.05904
R1178 B.n335 B.n334 4.05904
R1179 B.n350 B.n148 4.05904
R1180 VP.n27 VP.n26 161.3
R1181 VP.n28 VP.n23 161.3
R1182 VP.n30 VP.n29 161.3
R1183 VP.n31 VP.n22 161.3
R1184 VP.n33 VP.n32 161.3
R1185 VP.n34 VP.n21 161.3
R1186 VP.n36 VP.n35 161.3
R1187 VP.n37 VP.n20 161.3
R1188 VP.n39 VP.n38 161.3
R1189 VP.n40 VP.n19 161.3
R1190 VP.n42 VP.n41 161.3
R1191 VP.n43 VP.n18 161.3
R1192 VP.n45 VP.n44 161.3
R1193 VP.n47 VP.n46 161.3
R1194 VP.n48 VP.n16 161.3
R1195 VP.n50 VP.n49 161.3
R1196 VP.n51 VP.n15 161.3
R1197 VP.n53 VP.n52 161.3
R1198 VP.n54 VP.n14 161.3
R1199 VP.n96 VP.n0 161.3
R1200 VP.n95 VP.n94 161.3
R1201 VP.n93 VP.n1 161.3
R1202 VP.n92 VP.n91 161.3
R1203 VP.n90 VP.n2 161.3
R1204 VP.n89 VP.n88 161.3
R1205 VP.n87 VP.n86 161.3
R1206 VP.n85 VP.n4 161.3
R1207 VP.n84 VP.n83 161.3
R1208 VP.n82 VP.n5 161.3
R1209 VP.n81 VP.n80 161.3
R1210 VP.n79 VP.n6 161.3
R1211 VP.n78 VP.n77 161.3
R1212 VP.n76 VP.n7 161.3
R1213 VP.n75 VP.n74 161.3
R1214 VP.n73 VP.n8 161.3
R1215 VP.n72 VP.n71 161.3
R1216 VP.n70 VP.n9 161.3
R1217 VP.n69 VP.n68 161.3
R1218 VP.n66 VP.n10 161.3
R1219 VP.n65 VP.n64 161.3
R1220 VP.n63 VP.n11 161.3
R1221 VP.n62 VP.n61 161.3
R1222 VP.n60 VP.n12 161.3
R1223 VP.n59 VP.n58 161.3
R1224 VP.n57 VP.n13 102.927
R1225 VP.n98 VP.n97 102.927
R1226 VP.n56 VP.n55 102.927
R1227 VP.n24 VP.t6 99.4197
R1228 VP.n25 VP.n24 68.8984
R1229 VP.n78 VP.t2 66.5165
R1230 VP.n13 VP.t0 66.5165
R1231 VP.n67 VP.t4 66.5165
R1232 VP.n3 VP.t3 66.5165
R1233 VP.n97 VP.t9 66.5165
R1234 VP.n36 VP.t7 66.5165
R1235 VP.n55 VP.t1 66.5165
R1236 VP.n17 VP.t5 66.5165
R1237 VP.n25 VP.t8 66.5165
R1238 VP.n61 VP.n11 52.1486
R1239 VP.n91 VP.n1 52.1486
R1240 VP.n49 VP.n15 52.1486
R1241 VP.n57 VP.n56 50.6132
R1242 VP.n73 VP.n72 44.3785
R1243 VP.n84 VP.n5 44.3785
R1244 VP.n42 VP.n19 44.3785
R1245 VP.n31 VP.n30 44.3785
R1246 VP.n74 VP.n73 36.6083
R1247 VP.n80 VP.n5 36.6083
R1248 VP.n38 VP.n19 36.6083
R1249 VP.n32 VP.n31 36.6083
R1250 VP.n65 VP.n11 28.8382
R1251 VP.n91 VP.n90 28.8382
R1252 VP.n49 VP.n48 28.8382
R1253 VP.n60 VP.n59 24.4675
R1254 VP.n61 VP.n60 24.4675
R1255 VP.n66 VP.n65 24.4675
R1256 VP.n68 VP.n9 24.4675
R1257 VP.n72 VP.n9 24.4675
R1258 VP.n74 VP.n7 24.4675
R1259 VP.n78 VP.n7 24.4675
R1260 VP.n79 VP.n78 24.4675
R1261 VP.n80 VP.n79 24.4675
R1262 VP.n85 VP.n84 24.4675
R1263 VP.n86 VP.n85 24.4675
R1264 VP.n90 VP.n89 24.4675
R1265 VP.n95 VP.n1 24.4675
R1266 VP.n96 VP.n95 24.4675
R1267 VP.n53 VP.n15 24.4675
R1268 VP.n54 VP.n53 24.4675
R1269 VP.n43 VP.n42 24.4675
R1270 VP.n44 VP.n43 24.4675
R1271 VP.n48 VP.n47 24.4675
R1272 VP.n32 VP.n21 24.4675
R1273 VP.n36 VP.n21 24.4675
R1274 VP.n37 VP.n36 24.4675
R1275 VP.n38 VP.n37 24.4675
R1276 VP.n26 VP.n23 24.4675
R1277 VP.n30 VP.n23 24.4675
R1278 VP.n67 VP.n66 20.5528
R1279 VP.n89 VP.n3 20.5528
R1280 VP.n47 VP.n17 20.5528
R1281 VP.n59 VP.n13 7.82994
R1282 VP.n97 VP.n96 7.82994
R1283 VP.n55 VP.n54 7.82994
R1284 VP.n27 VP.n24 6.98708
R1285 VP.n68 VP.n67 3.91522
R1286 VP.n86 VP.n3 3.91522
R1287 VP.n44 VP.n17 3.91522
R1288 VP.n26 VP.n25 3.91522
R1289 VP.n56 VP.n14 0.278367
R1290 VP.n58 VP.n57 0.278367
R1291 VP.n98 VP.n0 0.278367
R1292 VP.n28 VP.n27 0.189894
R1293 VP.n29 VP.n28 0.189894
R1294 VP.n29 VP.n22 0.189894
R1295 VP.n33 VP.n22 0.189894
R1296 VP.n34 VP.n33 0.189894
R1297 VP.n35 VP.n34 0.189894
R1298 VP.n35 VP.n20 0.189894
R1299 VP.n39 VP.n20 0.189894
R1300 VP.n40 VP.n39 0.189894
R1301 VP.n41 VP.n40 0.189894
R1302 VP.n41 VP.n18 0.189894
R1303 VP.n45 VP.n18 0.189894
R1304 VP.n46 VP.n45 0.189894
R1305 VP.n46 VP.n16 0.189894
R1306 VP.n50 VP.n16 0.189894
R1307 VP.n51 VP.n50 0.189894
R1308 VP.n52 VP.n51 0.189894
R1309 VP.n52 VP.n14 0.189894
R1310 VP.n58 VP.n12 0.189894
R1311 VP.n62 VP.n12 0.189894
R1312 VP.n63 VP.n62 0.189894
R1313 VP.n64 VP.n63 0.189894
R1314 VP.n64 VP.n10 0.189894
R1315 VP.n69 VP.n10 0.189894
R1316 VP.n70 VP.n69 0.189894
R1317 VP.n71 VP.n70 0.189894
R1318 VP.n71 VP.n8 0.189894
R1319 VP.n75 VP.n8 0.189894
R1320 VP.n76 VP.n75 0.189894
R1321 VP.n77 VP.n76 0.189894
R1322 VP.n77 VP.n6 0.189894
R1323 VP.n81 VP.n6 0.189894
R1324 VP.n82 VP.n81 0.189894
R1325 VP.n83 VP.n82 0.189894
R1326 VP.n83 VP.n4 0.189894
R1327 VP.n87 VP.n4 0.189894
R1328 VP.n88 VP.n87 0.189894
R1329 VP.n88 VP.n2 0.189894
R1330 VP.n92 VP.n2 0.189894
R1331 VP.n93 VP.n92 0.189894
R1332 VP.n94 VP.n93 0.189894
R1333 VP.n94 VP.n0 0.189894
R1334 VP VP.n98 0.153454
R1335 VTAIL.n11 VTAIL.t5 74.0531
R1336 VTAIL.n17 VTAIL.t3 74.0529
R1337 VTAIL.n2 VTAIL.t18 74.0529
R1338 VTAIL.n16 VTAIL.t12 74.0529
R1339 VTAIL.n15 VTAIL.n14 69.7705
R1340 VTAIL.n13 VTAIL.n12 69.7705
R1341 VTAIL.n10 VTAIL.n9 69.7705
R1342 VTAIL.n8 VTAIL.n7 69.7705
R1343 VTAIL.n19 VTAIL.n18 69.7703
R1344 VTAIL.n1 VTAIL.n0 69.7703
R1345 VTAIL.n4 VTAIL.n3 69.7703
R1346 VTAIL.n6 VTAIL.n5 69.7703
R1347 VTAIL.n8 VTAIL.n6 24.2203
R1348 VTAIL.n17 VTAIL.n16 21.5652
R1349 VTAIL.n18 VTAIL.t1 4.28311
R1350 VTAIL.n18 VTAIL.t8 4.28311
R1351 VTAIL.n0 VTAIL.t4 4.28311
R1352 VTAIL.n0 VTAIL.t6 4.28311
R1353 VTAIL.n3 VTAIL.t19 4.28311
R1354 VTAIL.n3 VTAIL.t13 4.28311
R1355 VTAIL.n5 VTAIL.t10 4.28311
R1356 VTAIL.n5 VTAIL.t14 4.28311
R1357 VTAIL.n14 VTAIL.t11 4.28311
R1358 VTAIL.n14 VTAIL.t15 4.28311
R1359 VTAIL.n12 VTAIL.t16 4.28311
R1360 VTAIL.n12 VTAIL.t17 4.28311
R1361 VTAIL.n9 VTAIL.t7 4.28311
R1362 VTAIL.n9 VTAIL.t9 4.28311
R1363 VTAIL.n7 VTAIL.t2 4.28311
R1364 VTAIL.n7 VTAIL.t0 4.28311
R1365 VTAIL.n10 VTAIL.n8 2.65567
R1366 VTAIL.n11 VTAIL.n10 2.65567
R1367 VTAIL.n15 VTAIL.n13 2.65567
R1368 VTAIL.n16 VTAIL.n15 2.65567
R1369 VTAIL.n6 VTAIL.n4 2.65567
R1370 VTAIL.n4 VTAIL.n2 2.65567
R1371 VTAIL.n19 VTAIL.n17 2.65567
R1372 VTAIL VTAIL.n1 2.05007
R1373 VTAIL.n13 VTAIL.n11 1.79791
R1374 VTAIL.n2 VTAIL.n1 1.79791
R1375 VTAIL VTAIL.n19 0.606103
R1376 VDD1.n1 VDD1.t3 93.387
R1377 VDD1.n3 VDD1.t9 93.3868
R1378 VDD1.n5 VDD1.n4 88.3851
R1379 VDD1.n1 VDD1.n0 86.4493
R1380 VDD1.n7 VDD1.n6 86.449
R1381 VDD1.n3 VDD1.n2 86.449
R1382 VDD1.n7 VDD1.n5 44.7811
R1383 VDD1.n6 VDD1.t4 4.28311
R1384 VDD1.n6 VDD1.t8 4.28311
R1385 VDD1.n0 VDD1.t1 4.28311
R1386 VDD1.n0 VDD1.t2 4.28311
R1387 VDD1.n4 VDD1.t6 4.28311
R1388 VDD1.n4 VDD1.t0 4.28311
R1389 VDD1.n2 VDD1.t5 4.28311
R1390 VDD1.n2 VDD1.t7 4.28311
R1391 VDD1 VDD1.n7 1.93369
R1392 VDD1 VDD1.n1 0.722483
R1393 VDD1.n5 VDD1.n3 0.608947
R1394 VN.n83 VN.n43 161.3
R1395 VN.n82 VN.n81 161.3
R1396 VN.n80 VN.n44 161.3
R1397 VN.n79 VN.n78 161.3
R1398 VN.n77 VN.n45 161.3
R1399 VN.n76 VN.n75 161.3
R1400 VN.n74 VN.n73 161.3
R1401 VN.n72 VN.n47 161.3
R1402 VN.n71 VN.n70 161.3
R1403 VN.n69 VN.n48 161.3
R1404 VN.n68 VN.n67 161.3
R1405 VN.n66 VN.n49 161.3
R1406 VN.n65 VN.n64 161.3
R1407 VN.n63 VN.n50 161.3
R1408 VN.n62 VN.n61 161.3
R1409 VN.n60 VN.n51 161.3
R1410 VN.n59 VN.n58 161.3
R1411 VN.n57 VN.n52 161.3
R1412 VN.n56 VN.n55 161.3
R1413 VN.n40 VN.n0 161.3
R1414 VN.n39 VN.n38 161.3
R1415 VN.n37 VN.n1 161.3
R1416 VN.n36 VN.n35 161.3
R1417 VN.n34 VN.n2 161.3
R1418 VN.n33 VN.n32 161.3
R1419 VN.n31 VN.n30 161.3
R1420 VN.n29 VN.n4 161.3
R1421 VN.n28 VN.n27 161.3
R1422 VN.n26 VN.n5 161.3
R1423 VN.n25 VN.n24 161.3
R1424 VN.n23 VN.n6 161.3
R1425 VN.n22 VN.n21 161.3
R1426 VN.n20 VN.n7 161.3
R1427 VN.n19 VN.n18 161.3
R1428 VN.n17 VN.n8 161.3
R1429 VN.n16 VN.n15 161.3
R1430 VN.n14 VN.n9 161.3
R1431 VN.n13 VN.n12 161.3
R1432 VN.n42 VN.n41 102.927
R1433 VN.n85 VN.n84 102.927
R1434 VN.n10 VN.t5 99.4197
R1435 VN.n53 VN.t2 99.4197
R1436 VN.n11 VN.n10 68.8984
R1437 VN.n54 VN.n53 68.8984
R1438 VN.n22 VN.t1 66.5165
R1439 VN.n11 VN.t0 66.5165
R1440 VN.n3 VN.t8 66.5165
R1441 VN.n41 VN.t9 66.5165
R1442 VN.n65 VN.t6 66.5165
R1443 VN.n54 VN.t3 66.5165
R1444 VN.n46 VN.t4 66.5165
R1445 VN.n84 VN.t7 66.5165
R1446 VN.n35 VN.n1 52.1486
R1447 VN.n78 VN.n44 52.1486
R1448 VN VN.n85 50.8921
R1449 VN.n17 VN.n16 44.3785
R1450 VN.n28 VN.n5 44.3785
R1451 VN.n60 VN.n59 44.3785
R1452 VN.n71 VN.n48 44.3785
R1453 VN.n18 VN.n17 36.6083
R1454 VN.n24 VN.n5 36.6083
R1455 VN.n61 VN.n60 36.6083
R1456 VN.n67 VN.n48 36.6083
R1457 VN.n35 VN.n34 28.8382
R1458 VN.n78 VN.n77 28.8382
R1459 VN.n12 VN.n9 24.4675
R1460 VN.n16 VN.n9 24.4675
R1461 VN.n18 VN.n7 24.4675
R1462 VN.n22 VN.n7 24.4675
R1463 VN.n23 VN.n22 24.4675
R1464 VN.n24 VN.n23 24.4675
R1465 VN.n29 VN.n28 24.4675
R1466 VN.n30 VN.n29 24.4675
R1467 VN.n34 VN.n33 24.4675
R1468 VN.n39 VN.n1 24.4675
R1469 VN.n40 VN.n39 24.4675
R1470 VN.n59 VN.n52 24.4675
R1471 VN.n55 VN.n52 24.4675
R1472 VN.n67 VN.n66 24.4675
R1473 VN.n66 VN.n65 24.4675
R1474 VN.n65 VN.n50 24.4675
R1475 VN.n61 VN.n50 24.4675
R1476 VN.n77 VN.n76 24.4675
R1477 VN.n73 VN.n72 24.4675
R1478 VN.n72 VN.n71 24.4675
R1479 VN.n83 VN.n82 24.4675
R1480 VN.n82 VN.n44 24.4675
R1481 VN.n33 VN.n3 20.5528
R1482 VN.n76 VN.n46 20.5528
R1483 VN.n41 VN.n40 7.82994
R1484 VN.n84 VN.n83 7.82994
R1485 VN.n56 VN.n53 6.98708
R1486 VN.n13 VN.n10 6.98708
R1487 VN.n12 VN.n11 3.91522
R1488 VN.n30 VN.n3 3.91522
R1489 VN.n55 VN.n54 3.91522
R1490 VN.n73 VN.n46 3.91522
R1491 VN.n85 VN.n43 0.278367
R1492 VN.n42 VN.n0 0.278367
R1493 VN.n81 VN.n43 0.189894
R1494 VN.n81 VN.n80 0.189894
R1495 VN.n80 VN.n79 0.189894
R1496 VN.n79 VN.n45 0.189894
R1497 VN.n75 VN.n45 0.189894
R1498 VN.n75 VN.n74 0.189894
R1499 VN.n74 VN.n47 0.189894
R1500 VN.n70 VN.n47 0.189894
R1501 VN.n70 VN.n69 0.189894
R1502 VN.n69 VN.n68 0.189894
R1503 VN.n68 VN.n49 0.189894
R1504 VN.n64 VN.n49 0.189894
R1505 VN.n64 VN.n63 0.189894
R1506 VN.n63 VN.n62 0.189894
R1507 VN.n62 VN.n51 0.189894
R1508 VN.n58 VN.n51 0.189894
R1509 VN.n58 VN.n57 0.189894
R1510 VN.n57 VN.n56 0.189894
R1511 VN.n14 VN.n13 0.189894
R1512 VN.n15 VN.n14 0.189894
R1513 VN.n15 VN.n8 0.189894
R1514 VN.n19 VN.n8 0.189894
R1515 VN.n20 VN.n19 0.189894
R1516 VN.n21 VN.n20 0.189894
R1517 VN.n21 VN.n6 0.189894
R1518 VN.n25 VN.n6 0.189894
R1519 VN.n26 VN.n25 0.189894
R1520 VN.n27 VN.n26 0.189894
R1521 VN.n27 VN.n4 0.189894
R1522 VN.n31 VN.n4 0.189894
R1523 VN.n32 VN.n31 0.189894
R1524 VN.n32 VN.n2 0.189894
R1525 VN.n36 VN.n2 0.189894
R1526 VN.n37 VN.n36 0.189894
R1527 VN.n38 VN.n37 0.189894
R1528 VN.n38 VN.n0 0.189894
R1529 VN VN.n42 0.153454
R1530 VDD2.n1 VDD2.t4 93.3868
R1531 VDD2.n4 VDD2.t2 90.7319
R1532 VDD2.n3 VDD2.n2 88.3851
R1533 VDD2 VDD2.n7 88.3822
R1534 VDD2.n6 VDD2.n5 86.4493
R1535 VDD2.n1 VDD2.n0 86.449
R1536 VDD2.n4 VDD2.n3 42.8705
R1537 VDD2.n7 VDD2.t6 4.28311
R1538 VDD2.n7 VDD2.t7 4.28311
R1539 VDD2.n5 VDD2.t5 4.28311
R1540 VDD2.n5 VDD2.t3 4.28311
R1541 VDD2.n2 VDD2.t1 4.28311
R1542 VDD2.n2 VDD2.t0 4.28311
R1543 VDD2.n0 VDD2.t9 4.28311
R1544 VDD2.n0 VDD2.t8 4.28311
R1545 VDD2.n6 VDD2.n4 2.65567
R1546 VDD2 VDD2.n6 0.722483
R1547 VDD2.n3 VDD2.n1 0.608947
C0 VDD2 VN 7.0146f
C1 VN B 1.26971f
C2 VDD2 VTAIL 8.50537f
C3 VTAIL B 2.79453f
C4 VP w_n4666_n2486# 10.548201f
C5 VDD2 VDD1 2.27048f
C6 VDD1 B 2.18941f
C7 VTAIL VN 7.91777f
C8 VDD2 VP 0.602219f
C9 VDD1 VN 0.153546f
C10 VP B 2.29284f
C11 VTAIL VDD1 8.452291f
C12 VP VN 7.80083f
C13 VTAIL VP 7.93198f
C14 VDD2 w_n4666_n2486# 2.68951f
C15 w_n4666_n2486# B 9.56293f
C16 VP VDD1 7.460161f
C17 w_n4666_n2486# VN 9.9402f
C18 VDD2 B 2.31317f
C19 VTAIL w_n4666_n2486# 2.61538f
C20 w_n4666_n2486# VDD1 2.53816f
C21 VDD2 VSUBS 2.146841f
C22 VDD1 VSUBS 1.916557f
C23 VTAIL VSUBS 1.193877f
C24 VN VSUBS 7.84527f
C25 VP VSUBS 4.266276f
C26 B VSUBS 5.183023f
C27 w_n4666_n2486# VSUBS 0.144067p
C28 VDD2.t4 VSUBS 1.88702f
C29 VDD2.t9 VSUBS 0.196406f
C30 VDD2.t8 VSUBS 0.196406f
C31 VDD2.n0 VSUBS 1.40766f
C32 VDD2.n1 VSUBS 1.78423f
C33 VDD2.t1 VSUBS 0.196406f
C34 VDD2.t0 VSUBS 0.196406f
C35 VDD2.n2 VSUBS 1.4305f
C36 VDD2.n3 VSUBS 3.82937f
C37 VDD2.t2 VSUBS 1.86086f
C38 VDD2.n4 VSUBS 3.99097f
C39 VDD2.t5 VSUBS 0.196406f
C40 VDD2.t3 VSUBS 0.196406f
C41 VDD2.n5 VSUBS 1.40766f
C42 VDD2.n6 VSUBS 0.900829f
C43 VDD2.t6 VSUBS 0.196406f
C44 VDD2.t7 VSUBS 0.196406f
C45 VDD2.n7 VSUBS 1.43045f
C46 VN.n0 VSUBS 0.04177f
C47 VN.t9 VSUBS 1.77186f
C48 VN.n1 VSUBS 0.056879f
C49 VN.n2 VSUBS 0.031682f
C50 VN.t8 VSUBS 1.77186f
C51 VN.n3 VSUBS 0.646901f
C52 VN.n4 VSUBS 0.031682f
C53 VN.n5 VSUBS 0.026269f
C54 VN.n6 VSUBS 0.031682f
C55 VN.t1 VSUBS 1.77186f
C56 VN.n7 VSUBS 0.059048f
C57 VN.n8 VSUBS 0.031682f
C58 VN.n9 VSUBS 0.059048f
C59 VN.t5 VSUBS 2.05311f
C60 VN.n10 VSUBS 0.711254f
C61 VN.t0 VSUBS 1.77186f
C62 VN.n11 VSUBS 0.732613f
C63 VN.n12 VSUBS 0.03456f
C64 VN.n13 VSUBS 0.31116f
C65 VN.n14 VSUBS 0.031682f
C66 VN.n15 VSUBS 0.031682f
C67 VN.n16 VSUBS 0.0614f
C68 VN.n17 VSUBS 0.026269f
C69 VN.n18 VSUBS 0.06388f
C70 VN.n19 VSUBS 0.031682f
C71 VN.n20 VSUBS 0.031682f
C72 VN.n21 VSUBS 0.031682f
C73 VN.n22 VSUBS 0.676797f
C74 VN.n23 VSUBS 0.059048f
C75 VN.n24 VSUBS 0.06388f
C76 VN.n25 VSUBS 0.031682f
C77 VN.n26 VSUBS 0.031682f
C78 VN.n27 VSUBS 0.031682f
C79 VN.n28 VSUBS 0.0614f
C80 VN.n29 VSUBS 0.059048f
C81 VN.n30 VSUBS 0.03456f
C82 VN.n31 VSUBS 0.031682f
C83 VN.n32 VSUBS 0.031682f
C84 VN.n33 VSUBS 0.054384f
C85 VN.n34 VSUBS 0.062669f
C86 VN.n35 VSUBS 0.032001f
C87 VN.n36 VSUBS 0.031682f
C88 VN.n37 VSUBS 0.031682f
C89 VN.n38 VSUBS 0.031682f
C90 VN.n39 VSUBS 0.059048f
C91 VN.n40 VSUBS 0.039224f
C92 VN.n41 VSUBS 0.755759f
C93 VN.n42 VSUBS 0.054856f
C94 VN.n43 VSUBS 0.04177f
C95 VN.t7 VSUBS 1.77186f
C96 VN.n44 VSUBS 0.056879f
C97 VN.n45 VSUBS 0.031682f
C98 VN.t4 VSUBS 1.77186f
C99 VN.n46 VSUBS 0.646901f
C100 VN.n47 VSUBS 0.031682f
C101 VN.n48 VSUBS 0.026269f
C102 VN.n49 VSUBS 0.031682f
C103 VN.t6 VSUBS 1.77186f
C104 VN.n50 VSUBS 0.059048f
C105 VN.n51 VSUBS 0.031682f
C106 VN.n52 VSUBS 0.059048f
C107 VN.t2 VSUBS 2.05311f
C108 VN.n53 VSUBS 0.711254f
C109 VN.t3 VSUBS 1.77186f
C110 VN.n54 VSUBS 0.732613f
C111 VN.n55 VSUBS 0.03456f
C112 VN.n56 VSUBS 0.31116f
C113 VN.n57 VSUBS 0.031682f
C114 VN.n58 VSUBS 0.031682f
C115 VN.n59 VSUBS 0.0614f
C116 VN.n60 VSUBS 0.026269f
C117 VN.n61 VSUBS 0.06388f
C118 VN.n62 VSUBS 0.031682f
C119 VN.n63 VSUBS 0.031682f
C120 VN.n64 VSUBS 0.031682f
C121 VN.n65 VSUBS 0.676797f
C122 VN.n66 VSUBS 0.059048f
C123 VN.n67 VSUBS 0.06388f
C124 VN.n68 VSUBS 0.031682f
C125 VN.n69 VSUBS 0.031682f
C126 VN.n70 VSUBS 0.031682f
C127 VN.n71 VSUBS 0.0614f
C128 VN.n72 VSUBS 0.059048f
C129 VN.n73 VSUBS 0.03456f
C130 VN.n74 VSUBS 0.031682f
C131 VN.n75 VSUBS 0.031682f
C132 VN.n76 VSUBS 0.054384f
C133 VN.n77 VSUBS 0.062669f
C134 VN.n78 VSUBS 0.032001f
C135 VN.n79 VSUBS 0.031682f
C136 VN.n80 VSUBS 0.031682f
C137 VN.n81 VSUBS 0.031682f
C138 VN.n82 VSUBS 0.059048f
C139 VN.n83 VSUBS 0.039224f
C140 VN.n84 VSUBS 0.755759f
C141 VN.n85 VSUBS 1.81546f
C142 VDD1.t3 VSUBS 1.89353f
C143 VDD1.t1 VSUBS 0.197083f
C144 VDD1.t2 VSUBS 0.197083f
C145 VDD1.n0 VSUBS 1.41252f
C146 VDD1.n1 VSUBS 1.80115f
C147 VDD1.t9 VSUBS 1.89353f
C148 VDD1.t5 VSUBS 0.197083f
C149 VDD1.t7 VSUBS 0.197083f
C150 VDD1.n2 VSUBS 1.41252f
C151 VDD1.n3 VSUBS 1.79039f
C152 VDD1.t6 VSUBS 0.197083f
C153 VDD1.t0 VSUBS 0.197083f
C154 VDD1.n4 VSUBS 1.43543f
C155 VDD1.n5 VSUBS 4.00767f
C156 VDD1.t4 VSUBS 0.197083f
C157 VDD1.t8 VSUBS 0.197083f
C158 VDD1.n6 VSUBS 1.41252f
C159 VDD1.n7 VSUBS 4.08295f
C160 VTAIL.t4 VSUBS 0.189272f
C161 VTAIL.t6 VSUBS 0.189272f
C162 VTAIL.n0 VSUBS 1.23253f
C163 VTAIL.n1 VSUBS 0.996992f
C164 VTAIL.t18 VSUBS 1.65854f
C165 VTAIL.n2 VSUBS 1.14876f
C166 VTAIL.t19 VSUBS 0.189272f
C167 VTAIL.t13 VSUBS 0.189272f
C168 VTAIL.n3 VSUBS 1.23253f
C169 VTAIL.n4 VSUBS 1.14579f
C170 VTAIL.t10 VSUBS 0.189272f
C171 VTAIL.t14 VSUBS 0.189272f
C172 VTAIL.n5 VSUBS 1.23253f
C173 VTAIL.n6 VSUBS 2.50975f
C174 VTAIL.t2 VSUBS 0.189272f
C175 VTAIL.t0 VSUBS 0.189272f
C176 VTAIL.n7 VSUBS 1.23254f
C177 VTAIL.n8 VSUBS 2.50975f
C178 VTAIL.t7 VSUBS 0.189272f
C179 VTAIL.t9 VSUBS 0.189272f
C180 VTAIL.n9 VSUBS 1.23254f
C181 VTAIL.n10 VSUBS 1.14579f
C182 VTAIL.t5 VSUBS 1.65854f
C183 VTAIL.n11 VSUBS 1.14875f
C184 VTAIL.t16 VSUBS 0.189272f
C185 VTAIL.t17 VSUBS 0.189272f
C186 VTAIL.n12 VSUBS 1.23254f
C187 VTAIL.n13 VSUBS 1.05857f
C188 VTAIL.t11 VSUBS 0.189272f
C189 VTAIL.t15 VSUBS 0.189272f
C190 VTAIL.n14 VSUBS 1.23254f
C191 VTAIL.n15 VSUBS 1.14579f
C192 VTAIL.t12 VSUBS 1.65854f
C193 VTAIL.n16 VSUBS 2.32995f
C194 VTAIL.t3 VSUBS 1.65854f
C195 VTAIL.n17 VSUBS 2.32995f
C196 VTAIL.t1 VSUBS 0.189272f
C197 VTAIL.t8 VSUBS 0.189272f
C198 VTAIL.n18 VSUBS 1.23253f
C199 VTAIL.n19 VSUBS 0.937385f
C200 VP.n0 VSUBS 0.04619f
C201 VP.t9 VSUBS 1.95933f
C202 VP.n1 VSUBS 0.062897f
C203 VP.n2 VSUBS 0.035035f
C204 VP.t3 VSUBS 1.95933f
C205 VP.n3 VSUBS 0.715347f
C206 VP.n4 VSUBS 0.035035f
C207 VP.n5 VSUBS 0.029049f
C208 VP.n6 VSUBS 0.035035f
C209 VP.t2 VSUBS 1.95933f
C210 VP.n7 VSUBS 0.065296f
C211 VP.n8 VSUBS 0.035035f
C212 VP.n9 VSUBS 0.065296f
C213 VP.n10 VSUBS 0.035035f
C214 VP.t4 VSUBS 1.95933f
C215 VP.n11 VSUBS 0.035387f
C216 VP.n12 VSUBS 0.035035f
C217 VP.t0 VSUBS 1.95933f
C218 VP.n13 VSUBS 0.835722f
C219 VP.n14 VSUBS 0.04619f
C220 VP.t1 VSUBS 1.95933f
C221 VP.n15 VSUBS 0.062897f
C222 VP.n16 VSUBS 0.035035f
C223 VP.t5 VSUBS 1.95933f
C224 VP.n17 VSUBS 0.715347f
C225 VP.n18 VSUBS 0.035035f
C226 VP.n19 VSUBS 0.029049f
C227 VP.n20 VSUBS 0.035035f
C228 VP.t7 VSUBS 1.95933f
C229 VP.n21 VSUBS 0.065296f
C230 VP.n22 VSUBS 0.035035f
C231 VP.n23 VSUBS 0.065296f
C232 VP.t6 VSUBS 2.27034f
C233 VP.n24 VSUBS 0.786508f
C234 VP.t8 VSUBS 1.95933f
C235 VP.n25 VSUBS 0.810128f
C236 VP.n26 VSUBS 0.038217f
C237 VP.n27 VSUBS 0.344083f
C238 VP.n28 VSUBS 0.035035f
C239 VP.n29 VSUBS 0.035035f
C240 VP.n30 VSUBS 0.067896f
C241 VP.n31 VSUBS 0.029049f
C242 VP.n32 VSUBS 0.070639f
C243 VP.n33 VSUBS 0.035035f
C244 VP.n34 VSUBS 0.035035f
C245 VP.n35 VSUBS 0.035035f
C246 VP.n36 VSUBS 0.748405f
C247 VP.n37 VSUBS 0.065296f
C248 VP.n38 VSUBS 0.070639f
C249 VP.n39 VSUBS 0.035035f
C250 VP.n40 VSUBS 0.035035f
C251 VP.n41 VSUBS 0.035035f
C252 VP.n42 VSUBS 0.067896f
C253 VP.n43 VSUBS 0.065296f
C254 VP.n44 VSUBS 0.038217f
C255 VP.n45 VSUBS 0.035035f
C256 VP.n46 VSUBS 0.035035f
C257 VP.n47 VSUBS 0.060138f
C258 VP.n48 VSUBS 0.0693f
C259 VP.n49 VSUBS 0.035387f
C260 VP.n50 VSUBS 0.035035f
C261 VP.n51 VSUBS 0.035035f
C262 VP.n52 VSUBS 0.035035f
C263 VP.n53 VSUBS 0.065296f
C264 VP.n54 VSUBS 0.043375f
C265 VP.n55 VSUBS 0.835722f
C266 VP.n56 VSUBS 1.98875f
C267 VP.n57 VSUBS 2.01364f
C268 VP.n58 VSUBS 0.04619f
C269 VP.n59 VSUBS 0.043375f
C270 VP.n60 VSUBS 0.065296f
C271 VP.n61 VSUBS 0.062897f
C272 VP.n62 VSUBS 0.035035f
C273 VP.n63 VSUBS 0.035035f
C274 VP.n64 VSUBS 0.035035f
C275 VP.n65 VSUBS 0.0693f
C276 VP.n66 VSUBS 0.060138f
C277 VP.n67 VSUBS 0.715347f
C278 VP.n68 VSUBS 0.038217f
C279 VP.n69 VSUBS 0.035035f
C280 VP.n70 VSUBS 0.035035f
C281 VP.n71 VSUBS 0.035035f
C282 VP.n72 VSUBS 0.067896f
C283 VP.n73 VSUBS 0.029049f
C284 VP.n74 VSUBS 0.070639f
C285 VP.n75 VSUBS 0.035035f
C286 VP.n76 VSUBS 0.035035f
C287 VP.n77 VSUBS 0.035035f
C288 VP.n78 VSUBS 0.748405f
C289 VP.n79 VSUBS 0.065296f
C290 VP.n80 VSUBS 0.070639f
C291 VP.n81 VSUBS 0.035035f
C292 VP.n82 VSUBS 0.035035f
C293 VP.n83 VSUBS 0.035035f
C294 VP.n84 VSUBS 0.067896f
C295 VP.n85 VSUBS 0.065296f
C296 VP.n86 VSUBS 0.038217f
C297 VP.n87 VSUBS 0.035035f
C298 VP.n88 VSUBS 0.035035f
C299 VP.n89 VSUBS 0.060138f
C300 VP.n90 VSUBS 0.0693f
C301 VP.n91 VSUBS 0.035387f
C302 VP.n92 VSUBS 0.035035f
C303 VP.n93 VSUBS 0.035035f
C304 VP.n94 VSUBS 0.035035f
C305 VP.n95 VSUBS 0.065296f
C306 VP.n96 VSUBS 0.043375f
C307 VP.n97 VSUBS 0.835722f
C308 VP.n98 VSUBS 0.06066f
C309 B.n0 VSUBS 0.009626f
C310 B.n1 VSUBS 0.009626f
C311 B.n2 VSUBS 0.014236f
C312 B.n3 VSUBS 0.010909f
C313 B.n4 VSUBS 0.010909f
C314 B.n5 VSUBS 0.010909f
C315 B.n6 VSUBS 0.010909f
C316 B.n7 VSUBS 0.010909f
C317 B.n8 VSUBS 0.010909f
C318 B.n9 VSUBS 0.010909f
C319 B.n10 VSUBS 0.010909f
C320 B.n11 VSUBS 0.010909f
C321 B.n12 VSUBS 0.010909f
C322 B.n13 VSUBS 0.010909f
C323 B.n14 VSUBS 0.010909f
C324 B.n15 VSUBS 0.010909f
C325 B.n16 VSUBS 0.010909f
C326 B.n17 VSUBS 0.010909f
C327 B.n18 VSUBS 0.010909f
C328 B.n19 VSUBS 0.010909f
C329 B.n20 VSUBS 0.010909f
C330 B.n21 VSUBS 0.010909f
C331 B.n22 VSUBS 0.010909f
C332 B.n23 VSUBS 0.010909f
C333 B.n24 VSUBS 0.010909f
C334 B.n25 VSUBS 0.010909f
C335 B.n26 VSUBS 0.010909f
C336 B.n27 VSUBS 0.010909f
C337 B.n28 VSUBS 0.010909f
C338 B.n29 VSUBS 0.010909f
C339 B.n30 VSUBS 0.010909f
C340 B.n31 VSUBS 0.010909f
C341 B.n32 VSUBS 0.010909f
C342 B.n33 VSUBS 0.025538f
C343 B.n34 VSUBS 0.010909f
C344 B.n35 VSUBS 0.010909f
C345 B.n36 VSUBS 0.010909f
C346 B.n37 VSUBS 0.010909f
C347 B.n38 VSUBS 0.010909f
C348 B.n39 VSUBS 0.010909f
C349 B.n40 VSUBS 0.010909f
C350 B.n41 VSUBS 0.010909f
C351 B.n42 VSUBS 0.010909f
C352 B.n43 VSUBS 0.010909f
C353 B.n44 VSUBS 0.010909f
C354 B.n45 VSUBS 0.010909f
C355 B.n46 VSUBS 0.010909f
C356 B.n47 VSUBS 0.010909f
C357 B.t1 VSUBS 0.361758f
C358 B.t2 VSUBS 0.395506f
C359 B.t0 VSUBS 1.52557f
C360 B.n48 VSUBS 0.219001f
C361 B.n49 VSUBS 0.112084f
C362 B.n50 VSUBS 0.010909f
C363 B.n51 VSUBS 0.010909f
C364 B.n52 VSUBS 0.010909f
C365 B.n53 VSUBS 0.010909f
C366 B.t10 VSUBS 0.361756f
C367 B.t11 VSUBS 0.395503f
C368 B.t9 VSUBS 1.52557f
C369 B.n54 VSUBS 0.219005f
C370 B.n55 VSUBS 0.112087f
C371 B.n56 VSUBS 0.025276f
C372 B.n57 VSUBS 0.010909f
C373 B.n58 VSUBS 0.010909f
C374 B.n59 VSUBS 0.010909f
C375 B.n60 VSUBS 0.010909f
C376 B.n61 VSUBS 0.010909f
C377 B.n62 VSUBS 0.010909f
C378 B.n63 VSUBS 0.010909f
C379 B.n64 VSUBS 0.010909f
C380 B.n65 VSUBS 0.010909f
C381 B.n66 VSUBS 0.010909f
C382 B.n67 VSUBS 0.010909f
C383 B.n68 VSUBS 0.010909f
C384 B.n69 VSUBS 0.010909f
C385 B.n70 VSUBS 0.010909f
C386 B.n71 VSUBS 0.024196f
C387 B.n72 VSUBS 0.010909f
C388 B.n73 VSUBS 0.010909f
C389 B.n74 VSUBS 0.010909f
C390 B.n75 VSUBS 0.010909f
C391 B.n76 VSUBS 0.010909f
C392 B.n77 VSUBS 0.010909f
C393 B.n78 VSUBS 0.010909f
C394 B.n79 VSUBS 0.010909f
C395 B.n80 VSUBS 0.010909f
C396 B.n81 VSUBS 0.010909f
C397 B.n82 VSUBS 0.010909f
C398 B.n83 VSUBS 0.010909f
C399 B.n84 VSUBS 0.010909f
C400 B.n85 VSUBS 0.010909f
C401 B.n86 VSUBS 0.010909f
C402 B.n87 VSUBS 0.010909f
C403 B.n88 VSUBS 0.010909f
C404 B.n89 VSUBS 0.010909f
C405 B.n90 VSUBS 0.010909f
C406 B.n91 VSUBS 0.010909f
C407 B.n92 VSUBS 0.010909f
C408 B.n93 VSUBS 0.010909f
C409 B.n94 VSUBS 0.010909f
C410 B.n95 VSUBS 0.010909f
C411 B.n96 VSUBS 0.010909f
C412 B.n97 VSUBS 0.010909f
C413 B.n98 VSUBS 0.010909f
C414 B.n99 VSUBS 0.010909f
C415 B.n100 VSUBS 0.010909f
C416 B.n101 VSUBS 0.010909f
C417 B.n102 VSUBS 0.010909f
C418 B.n103 VSUBS 0.010909f
C419 B.n104 VSUBS 0.010909f
C420 B.n105 VSUBS 0.010909f
C421 B.n106 VSUBS 0.010909f
C422 B.n107 VSUBS 0.010909f
C423 B.n108 VSUBS 0.010909f
C424 B.n109 VSUBS 0.010909f
C425 B.n110 VSUBS 0.010909f
C426 B.n111 VSUBS 0.010909f
C427 B.n112 VSUBS 0.010909f
C428 B.n113 VSUBS 0.010909f
C429 B.n114 VSUBS 0.010909f
C430 B.n115 VSUBS 0.010909f
C431 B.n116 VSUBS 0.010909f
C432 B.n117 VSUBS 0.010909f
C433 B.n118 VSUBS 0.010909f
C434 B.n119 VSUBS 0.010909f
C435 B.n120 VSUBS 0.010909f
C436 B.n121 VSUBS 0.010909f
C437 B.n122 VSUBS 0.010909f
C438 B.n123 VSUBS 0.010909f
C439 B.n124 VSUBS 0.010909f
C440 B.n125 VSUBS 0.010909f
C441 B.n126 VSUBS 0.010909f
C442 B.n127 VSUBS 0.010909f
C443 B.n128 VSUBS 0.010909f
C444 B.n129 VSUBS 0.010909f
C445 B.n130 VSUBS 0.010909f
C446 B.n131 VSUBS 0.010909f
C447 B.n132 VSUBS 0.010909f
C448 B.n133 VSUBS 0.010909f
C449 B.n134 VSUBS 0.024196f
C450 B.n135 VSUBS 0.010909f
C451 B.n136 VSUBS 0.010909f
C452 B.n137 VSUBS 0.010909f
C453 B.n138 VSUBS 0.010909f
C454 B.n139 VSUBS 0.010909f
C455 B.n140 VSUBS 0.010909f
C456 B.n141 VSUBS 0.010909f
C457 B.n142 VSUBS 0.010909f
C458 B.n143 VSUBS 0.010909f
C459 B.n144 VSUBS 0.010909f
C460 B.n145 VSUBS 0.010909f
C461 B.n146 VSUBS 0.010909f
C462 B.n147 VSUBS 0.010909f
C463 B.n148 VSUBS 0.00754f
C464 B.n149 VSUBS 0.010909f
C465 B.n150 VSUBS 0.010909f
C466 B.n151 VSUBS 0.010909f
C467 B.n152 VSUBS 0.010909f
C468 B.n153 VSUBS 0.010909f
C469 B.t5 VSUBS 0.361758f
C470 B.t4 VSUBS 0.395506f
C471 B.t3 VSUBS 1.52557f
C472 B.n154 VSUBS 0.219001f
C473 B.n155 VSUBS 0.112084f
C474 B.n156 VSUBS 0.010909f
C475 B.n157 VSUBS 0.010909f
C476 B.n158 VSUBS 0.010909f
C477 B.n159 VSUBS 0.010909f
C478 B.n160 VSUBS 0.010909f
C479 B.n161 VSUBS 0.010909f
C480 B.n162 VSUBS 0.010909f
C481 B.n163 VSUBS 0.010909f
C482 B.n164 VSUBS 0.010909f
C483 B.n165 VSUBS 0.010909f
C484 B.n166 VSUBS 0.010909f
C485 B.n167 VSUBS 0.010909f
C486 B.n168 VSUBS 0.010909f
C487 B.n169 VSUBS 0.025538f
C488 B.n170 VSUBS 0.010909f
C489 B.n171 VSUBS 0.010909f
C490 B.n172 VSUBS 0.010909f
C491 B.n173 VSUBS 0.010909f
C492 B.n174 VSUBS 0.010909f
C493 B.n175 VSUBS 0.010909f
C494 B.n176 VSUBS 0.010909f
C495 B.n177 VSUBS 0.010909f
C496 B.n178 VSUBS 0.010909f
C497 B.n179 VSUBS 0.010909f
C498 B.n180 VSUBS 0.010909f
C499 B.n181 VSUBS 0.010909f
C500 B.n182 VSUBS 0.010909f
C501 B.n183 VSUBS 0.010909f
C502 B.n184 VSUBS 0.010909f
C503 B.n185 VSUBS 0.010909f
C504 B.n186 VSUBS 0.010909f
C505 B.n187 VSUBS 0.010909f
C506 B.n188 VSUBS 0.010909f
C507 B.n189 VSUBS 0.010909f
C508 B.n190 VSUBS 0.010909f
C509 B.n191 VSUBS 0.010909f
C510 B.n192 VSUBS 0.010909f
C511 B.n193 VSUBS 0.010909f
C512 B.n194 VSUBS 0.010909f
C513 B.n195 VSUBS 0.010909f
C514 B.n196 VSUBS 0.010909f
C515 B.n197 VSUBS 0.010909f
C516 B.n198 VSUBS 0.010909f
C517 B.n199 VSUBS 0.010909f
C518 B.n200 VSUBS 0.010909f
C519 B.n201 VSUBS 0.010909f
C520 B.n202 VSUBS 0.010909f
C521 B.n203 VSUBS 0.010909f
C522 B.n204 VSUBS 0.010909f
C523 B.n205 VSUBS 0.010909f
C524 B.n206 VSUBS 0.010909f
C525 B.n207 VSUBS 0.010909f
C526 B.n208 VSUBS 0.010909f
C527 B.n209 VSUBS 0.010909f
C528 B.n210 VSUBS 0.010909f
C529 B.n211 VSUBS 0.010909f
C530 B.n212 VSUBS 0.010909f
C531 B.n213 VSUBS 0.010909f
C532 B.n214 VSUBS 0.010909f
C533 B.n215 VSUBS 0.010909f
C534 B.n216 VSUBS 0.010909f
C535 B.n217 VSUBS 0.010909f
C536 B.n218 VSUBS 0.010909f
C537 B.n219 VSUBS 0.010909f
C538 B.n220 VSUBS 0.010909f
C539 B.n221 VSUBS 0.010909f
C540 B.n222 VSUBS 0.010909f
C541 B.n223 VSUBS 0.010909f
C542 B.n224 VSUBS 0.010909f
C543 B.n225 VSUBS 0.010909f
C544 B.n226 VSUBS 0.010909f
C545 B.n227 VSUBS 0.010909f
C546 B.n228 VSUBS 0.010909f
C547 B.n229 VSUBS 0.010909f
C548 B.n230 VSUBS 0.010909f
C549 B.n231 VSUBS 0.010909f
C550 B.n232 VSUBS 0.010909f
C551 B.n233 VSUBS 0.010909f
C552 B.n234 VSUBS 0.010909f
C553 B.n235 VSUBS 0.010909f
C554 B.n236 VSUBS 0.010909f
C555 B.n237 VSUBS 0.010909f
C556 B.n238 VSUBS 0.010909f
C557 B.n239 VSUBS 0.010909f
C558 B.n240 VSUBS 0.010909f
C559 B.n241 VSUBS 0.010909f
C560 B.n242 VSUBS 0.010909f
C561 B.n243 VSUBS 0.010909f
C562 B.n244 VSUBS 0.010909f
C563 B.n245 VSUBS 0.010909f
C564 B.n246 VSUBS 0.010909f
C565 B.n247 VSUBS 0.010909f
C566 B.n248 VSUBS 0.010909f
C567 B.n249 VSUBS 0.010909f
C568 B.n250 VSUBS 0.010909f
C569 B.n251 VSUBS 0.010909f
C570 B.n252 VSUBS 0.010909f
C571 B.n253 VSUBS 0.010909f
C572 B.n254 VSUBS 0.010909f
C573 B.n255 VSUBS 0.010909f
C574 B.n256 VSUBS 0.010909f
C575 B.n257 VSUBS 0.010909f
C576 B.n258 VSUBS 0.010909f
C577 B.n259 VSUBS 0.010909f
C578 B.n260 VSUBS 0.010909f
C579 B.n261 VSUBS 0.010909f
C580 B.n262 VSUBS 0.010909f
C581 B.n263 VSUBS 0.010909f
C582 B.n264 VSUBS 0.010909f
C583 B.n265 VSUBS 0.010909f
C584 B.n266 VSUBS 0.010909f
C585 B.n267 VSUBS 0.010909f
C586 B.n268 VSUBS 0.010909f
C587 B.n269 VSUBS 0.010909f
C588 B.n270 VSUBS 0.010909f
C589 B.n271 VSUBS 0.010909f
C590 B.n272 VSUBS 0.010909f
C591 B.n273 VSUBS 0.010909f
C592 B.n274 VSUBS 0.010909f
C593 B.n275 VSUBS 0.010909f
C594 B.n276 VSUBS 0.010909f
C595 B.n277 VSUBS 0.010909f
C596 B.n278 VSUBS 0.010909f
C597 B.n279 VSUBS 0.010909f
C598 B.n280 VSUBS 0.010909f
C599 B.n281 VSUBS 0.010909f
C600 B.n282 VSUBS 0.010909f
C601 B.n283 VSUBS 0.010909f
C602 B.n284 VSUBS 0.010909f
C603 B.n285 VSUBS 0.010909f
C604 B.n286 VSUBS 0.010909f
C605 B.n287 VSUBS 0.010909f
C606 B.n288 VSUBS 0.010909f
C607 B.n289 VSUBS 0.010909f
C608 B.n290 VSUBS 0.024196f
C609 B.n291 VSUBS 0.024196f
C610 B.n292 VSUBS 0.025538f
C611 B.n293 VSUBS 0.010909f
C612 B.n294 VSUBS 0.010909f
C613 B.n295 VSUBS 0.010909f
C614 B.n296 VSUBS 0.010909f
C615 B.n297 VSUBS 0.010909f
C616 B.n298 VSUBS 0.010909f
C617 B.n299 VSUBS 0.010909f
C618 B.n300 VSUBS 0.010909f
C619 B.n301 VSUBS 0.010909f
C620 B.n302 VSUBS 0.010909f
C621 B.n303 VSUBS 0.010909f
C622 B.n304 VSUBS 0.010909f
C623 B.n305 VSUBS 0.010909f
C624 B.n306 VSUBS 0.010909f
C625 B.n307 VSUBS 0.010909f
C626 B.n308 VSUBS 0.010909f
C627 B.n309 VSUBS 0.010909f
C628 B.n310 VSUBS 0.010909f
C629 B.n311 VSUBS 0.010909f
C630 B.n312 VSUBS 0.010909f
C631 B.n313 VSUBS 0.010909f
C632 B.n314 VSUBS 0.010909f
C633 B.n315 VSUBS 0.010909f
C634 B.n316 VSUBS 0.010909f
C635 B.n317 VSUBS 0.010909f
C636 B.n318 VSUBS 0.010909f
C637 B.n319 VSUBS 0.010909f
C638 B.n320 VSUBS 0.010909f
C639 B.n321 VSUBS 0.010909f
C640 B.n322 VSUBS 0.010909f
C641 B.n323 VSUBS 0.010909f
C642 B.n324 VSUBS 0.010909f
C643 B.n325 VSUBS 0.010909f
C644 B.n326 VSUBS 0.010909f
C645 B.n327 VSUBS 0.010909f
C646 B.n328 VSUBS 0.010909f
C647 B.n329 VSUBS 0.010909f
C648 B.n330 VSUBS 0.010909f
C649 B.n331 VSUBS 0.010909f
C650 B.n332 VSUBS 0.010909f
C651 B.n333 VSUBS 0.010909f
C652 B.n334 VSUBS 0.00754f
C653 B.n335 VSUBS 0.025276f
C654 B.n336 VSUBS 0.008824f
C655 B.n337 VSUBS 0.010909f
C656 B.n338 VSUBS 0.010909f
C657 B.n339 VSUBS 0.010909f
C658 B.n340 VSUBS 0.010909f
C659 B.n341 VSUBS 0.010909f
C660 B.n342 VSUBS 0.010909f
C661 B.n343 VSUBS 0.010909f
C662 B.n344 VSUBS 0.010909f
C663 B.n345 VSUBS 0.010909f
C664 B.n346 VSUBS 0.010909f
C665 B.n347 VSUBS 0.010909f
C666 B.t8 VSUBS 0.361756f
C667 B.t7 VSUBS 0.395503f
C668 B.t6 VSUBS 1.52557f
C669 B.n348 VSUBS 0.219005f
C670 B.n349 VSUBS 0.112087f
C671 B.n350 VSUBS 0.025276f
C672 B.n351 VSUBS 0.008824f
C673 B.n352 VSUBS 0.010909f
C674 B.n353 VSUBS 0.010909f
C675 B.n354 VSUBS 0.010909f
C676 B.n355 VSUBS 0.010909f
C677 B.n356 VSUBS 0.010909f
C678 B.n357 VSUBS 0.010909f
C679 B.n358 VSUBS 0.010909f
C680 B.n359 VSUBS 0.010909f
C681 B.n360 VSUBS 0.010909f
C682 B.n361 VSUBS 0.010909f
C683 B.n362 VSUBS 0.010909f
C684 B.n363 VSUBS 0.010909f
C685 B.n364 VSUBS 0.010909f
C686 B.n365 VSUBS 0.010909f
C687 B.n366 VSUBS 0.010909f
C688 B.n367 VSUBS 0.010909f
C689 B.n368 VSUBS 0.010909f
C690 B.n369 VSUBS 0.010909f
C691 B.n370 VSUBS 0.010909f
C692 B.n371 VSUBS 0.010909f
C693 B.n372 VSUBS 0.010909f
C694 B.n373 VSUBS 0.010909f
C695 B.n374 VSUBS 0.010909f
C696 B.n375 VSUBS 0.010909f
C697 B.n376 VSUBS 0.010909f
C698 B.n377 VSUBS 0.010909f
C699 B.n378 VSUBS 0.010909f
C700 B.n379 VSUBS 0.010909f
C701 B.n380 VSUBS 0.010909f
C702 B.n381 VSUBS 0.010909f
C703 B.n382 VSUBS 0.010909f
C704 B.n383 VSUBS 0.010909f
C705 B.n384 VSUBS 0.010909f
C706 B.n385 VSUBS 0.010909f
C707 B.n386 VSUBS 0.010909f
C708 B.n387 VSUBS 0.010909f
C709 B.n388 VSUBS 0.010909f
C710 B.n389 VSUBS 0.010909f
C711 B.n390 VSUBS 0.010909f
C712 B.n391 VSUBS 0.010909f
C713 B.n392 VSUBS 0.010909f
C714 B.n393 VSUBS 0.010909f
C715 B.n394 VSUBS 0.010909f
C716 B.n395 VSUBS 0.025538f
C717 B.n396 VSUBS 0.024196f
C718 B.n397 VSUBS 0.025538f
C719 B.n398 VSUBS 0.010909f
C720 B.n399 VSUBS 0.010909f
C721 B.n400 VSUBS 0.010909f
C722 B.n401 VSUBS 0.010909f
C723 B.n402 VSUBS 0.010909f
C724 B.n403 VSUBS 0.010909f
C725 B.n404 VSUBS 0.010909f
C726 B.n405 VSUBS 0.010909f
C727 B.n406 VSUBS 0.010909f
C728 B.n407 VSUBS 0.010909f
C729 B.n408 VSUBS 0.010909f
C730 B.n409 VSUBS 0.010909f
C731 B.n410 VSUBS 0.010909f
C732 B.n411 VSUBS 0.010909f
C733 B.n412 VSUBS 0.010909f
C734 B.n413 VSUBS 0.010909f
C735 B.n414 VSUBS 0.010909f
C736 B.n415 VSUBS 0.010909f
C737 B.n416 VSUBS 0.010909f
C738 B.n417 VSUBS 0.010909f
C739 B.n418 VSUBS 0.010909f
C740 B.n419 VSUBS 0.010909f
C741 B.n420 VSUBS 0.010909f
C742 B.n421 VSUBS 0.010909f
C743 B.n422 VSUBS 0.010909f
C744 B.n423 VSUBS 0.010909f
C745 B.n424 VSUBS 0.010909f
C746 B.n425 VSUBS 0.010909f
C747 B.n426 VSUBS 0.010909f
C748 B.n427 VSUBS 0.010909f
C749 B.n428 VSUBS 0.010909f
C750 B.n429 VSUBS 0.010909f
C751 B.n430 VSUBS 0.010909f
C752 B.n431 VSUBS 0.010909f
C753 B.n432 VSUBS 0.010909f
C754 B.n433 VSUBS 0.010909f
C755 B.n434 VSUBS 0.010909f
C756 B.n435 VSUBS 0.010909f
C757 B.n436 VSUBS 0.010909f
C758 B.n437 VSUBS 0.010909f
C759 B.n438 VSUBS 0.010909f
C760 B.n439 VSUBS 0.010909f
C761 B.n440 VSUBS 0.010909f
C762 B.n441 VSUBS 0.010909f
C763 B.n442 VSUBS 0.010909f
C764 B.n443 VSUBS 0.010909f
C765 B.n444 VSUBS 0.010909f
C766 B.n445 VSUBS 0.010909f
C767 B.n446 VSUBS 0.010909f
C768 B.n447 VSUBS 0.010909f
C769 B.n448 VSUBS 0.010909f
C770 B.n449 VSUBS 0.010909f
C771 B.n450 VSUBS 0.010909f
C772 B.n451 VSUBS 0.010909f
C773 B.n452 VSUBS 0.010909f
C774 B.n453 VSUBS 0.010909f
C775 B.n454 VSUBS 0.010909f
C776 B.n455 VSUBS 0.010909f
C777 B.n456 VSUBS 0.010909f
C778 B.n457 VSUBS 0.010909f
C779 B.n458 VSUBS 0.010909f
C780 B.n459 VSUBS 0.010909f
C781 B.n460 VSUBS 0.010909f
C782 B.n461 VSUBS 0.010909f
C783 B.n462 VSUBS 0.010909f
C784 B.n463 VSUBS 0.010909f
C785 B.n464 VSUBS 0.010909f
C786 B.n465 VSUBS 0.010909f
C787 B.n466 VSUBS 0.010909f
C788 B.n467 VSUBS 0.010909f
C789 B.n468 VSUBS 0.010909f
C790 B.n469 VSUBS 0.010909f
C791 B.n470 VSUBS 0.010909f
C792 B.n471 VSUBS 0.010909f
C793 B.n472 VSUBS 0.010909f
C794 B.n473 VSUBS 0.010909f
C795 B.n474 VSUBS 0.010909f
C796 B.n475 VSUBS 0.010909f
C797 B.n476 VSUBS 0.010909f
C798 B.n477 VSUBS 0.010909f
C799 B.n478 VSUBS 0.010909f
C800 B.n479 VSUBS 0.010909f
C801 B.n480 VSUBS 0.010909f
C802 B.n481 VSUBS 0.010909f
C803 B.n482 VSUBS 0.010909f
C804 B.n483 VSUBS 0.010909f
C805 B.n484 VSUBS 0.010909f
C806 B.n485 VSUBS 0.010909f
C807 B.n486 VSUBS 0.010909f
C808 B.n487 VSUBS 0.010909f
C809 B.n488 VSUBS 0.010909f
C810 B.n489 VSUBS 0.010909f
C811 B.n490 VSUBS 0.010909f
C812 B.n491 VSUBS 0.010909f
C813 B.n492 VSUBS 0.010909f
C814 B.n493 VSUBS 0.010909f
C815 B.n494 VSUBS 0.010909f
C816 B.n495 VSUBS 0.010909f
C817 B.n496 VSUBS 0.010909f
C818 B.n497 VSUBS 0.010909f
C819 B.n498 VSUBS 0.010909f
C820 B.n499 VSUBS 0.010909f
C821 B.n500 VSUBS 0.010909f
C822 B.n501 VSUBS 0.010909f
C823 B.n502 VSUBS 0.010909f
C824 B.n503 VSUBS 0.010909f
C825 B.n504 VSUBS 0.010909f
C826 B.n505 VSUBS 0.010909f
C827 B.n506 VSUBS 0.010909f
C828 B.n507 VSUBS 0.010909f
C829 B.n508 VSUBS 0.010909f
C830 B.n509 VSUBS 0.010909f
C831 B.n510 VSUBS 0.010909f
C832 B.n511 VSUBS 0.010909f
C833 B.n512 VSUBS 0.010909f
C834 B.n513 VSUBS 0.010909f
C835 B.n514 VSUBS 0.010909f
C836 B.n515 VSUBS 0.010909f
C837 B.n516 VSUBS 0.010909f
C838 B.n517 VSUBS 0.010909f
C839 B.n518 VSUBS 0.010909f
C840 B.n519 VSUBS 0.010909f
C841 B.n520 VSUBS 0.010909f
C842 B.n521 VSUBS 0.010909f
C843 B.n522 VSUBS 0.010909f
C844 B.n523 VSUBS 0.010909f
C845 B.n524 VSUBS 0.010909f
C846 B.n525 VSUBS 0.010909f
C847 B.n526 VSUBS 0.010909f
C848 B.n527 VSUBS 0.010909f
C849 B.n528 VSUBS 0.010909f
C850 B.n529 VSUBS 0.010909f
C851 B.n530 VSUBS 0.010909f
C852 B.n531 VSUBS 0.010909f
C853 B.n532 VSUBS 0.010909f
C854 B.n533 VSUBS 0.010909f
C855 B.n534 VSUBS 0.010909f
C856 B.n535 VSUBS 0.010909f
C857 B.n536 VSUBS 0.010909f
C858 B.n537 VSUBS 0.010909f
C859 B.n538 VSUBS 0.010909f
C860 B.n539 VSUBS 0.010909f
C861 B.n540 VSUBS 0.010909f
C862 B.n541 VSUBS 0.010909f
C863 B.n542 VSUBS 0.010909f
C864 B.n543 VSUBS 0.010909f
C865 B.n544 VSUBS 0.010909f
C866 B.n545 VSUBS 0.010909f
C867 B.n546 VSUBS 0.010909f
C868 B.n547 VSUBS 0.010909f
C869 B.n548 VSUBS 0.010909f
C870 B.n549 VSUBS 0.010909f
C871 B.n550 VSUBS 0.010909f
C872 B.n551 VSUBS 0.010909f
C873 B.n552 VSUBS 0.010909f
C874 B.n553 VSUBS 0.010909f
C875 B.n554 VSUBS 0.010909f
C876 B.n555 VSUBS 0.010909f
C877 B.n556 VSUBS 0.010909f
C878 B.n557 VSUBS 0.010909f
C879 B.n558 VSUBS 0.010909f
C880 B.n559 VSUBS 0.010909f
C881 B.n560 VSUBS 0.010909f
C882 B.n561 VSUBS 0.010909f
C883 B.n562 VSUBS 0.010909f
C884 B.n563 VSUBS 0.010909f
C885 B.n564 VSUBS 0.010909f
C886 B.n565 VSUBS 0.010909f
C887 B.n566 VSUBS 0.010909f
C888 B.n567 VSUBS 0.010909f
C889 B.n568 VSUBS 0.010909f
C890 B.n569 VSUBS 0.010909f
C891 B.n570 VSUBS 0.010909f
C892 B.n571 VSUBS 0.010909f
C893 B.n572 VSUBS 0.010909f
C894 B.n573 VSUBS 0.010909f
C895 B.n574 VSUBS 0.010909f
C896 B.n575 VSUBS 0.010909f
C897 B.n576 VSUBS 0.010909f
C898 B.n577 VSUBS 0.010909f
C899 B.n578 VSUBS 0.010909f
C900 B.n579 VSUBS 0.010909f
C901 B.n580 VSUBS 0.010909f
C902 B.n581 VSUBS 0.010909f
C903 B.n582 VSUBS 0.010909f
C904 B.n583 VSUBS 0.010909f
C905 B.n584 VSUBS 0.024196f
C906 B.n585 VSUBS 0.025538f
C907 B.n586 VSUBS 0.025538f
C908 B.n587 VSUBS 0.010909f
C909 B.n588 VSUBS 0.010909f
C910 B.n589 VSUBS 0.010909f
C911 B.n590 VSUBS 0.010909f
C912 B.n591 VSUBS 0.010909f
C913 B.n592 VSUBS 0.010909f
C914 B.n593 VSUBS 0.010909f
C915 B.n594 VSUBS 0.010909f
C916 B.n595 VSUBS 0.010909f
C917 B.n596 VSUBS 0.010909f
C918 B.n597 VSUBS 0.010909f
C919 B.n598 VSUBS 0.010909f
C920 B.n599 VSUBS 0.010909f
C921 B.n600 VSUBS 0.010909f
C922 B.n601 VSUBS 0.010909f
C923 B.n602 VSUBS 0.010909f
C924 B.n603 VSUBS 0.010909f
C925 B.n604 VSUBS 0.010909f
C926 B.n605 VSUBS 0.010909f
C927 B.n606 VSUBS 0.010909f
C928 B.n607 VSUBS 0.010909f
C929 B.n608 VSUBS 0.010909f
C930 B.n609 VSUBS 0.010909f
C931 B.n610 VSUBS 0.010909f
C932 B.n611 VSUBS 0.010909f
C933 B.n612 VSUBS 0.010909f
C934 B.n613 VSUBS 0.010909f
C935 B.n614 VSUBS 0.010909f
C936 B.n615 VSUBS 0.010909f
C937 B.n616 VSUBS 0.010909f
C938 B.n617 VSUBS 0.010909f
C939 B.n618 VSUBS 0.010909f
C940 B.n619 VSUBS 0.010909f
C941 B.n620 VSUBS 0.010909f
C942 B.n621 VSUBS 0.010909f
C943 B.n622 VSUBS 0.010909f
C944 B.n623 VSUBS 0.010909f
C945 B.n624 VSUBS 0.010909f
C946 B.n625 VSUBS 0.010909f
C947 B.n626 VSUBS 0.010909f
C948 B.n627 VSUBS 0.00754f
C949 B.n628 VSUBS 0.010909f
C950 B.n629 VSUBS 0.010909f
C951 B.n630 VSUBS 0.008824f
C952 B.n631 VSUBS 0.010909f
C953 B.n632 VSUBS 0.010909f
C954 B.n633 VSUBS 0.010909f
C955 B.n634 VSUBS 0.010909f
C956 B.n635 VSUBS 0.010909f
C957 B.n636 VSUBS 0.010909f
C958 B.n637 VSUBS 0.010909f
C959 B.n638 VSUBS 0.010909f
C960 B.n639 VSUBS 0.010909f
C961 B.n640 VSUBS 0.010909f
C962 B.n641 VSUBS 0.010909f
C963 B.n642 VSUBS 0.008824f
C964 B.n643 VSUBS 0.025276f
C965 B.n644 VSUBS 0.00754f
C966 B.n645 VSUBS 0.010909f
C967 B.n646 VSUBS 0.010909f
C968 B.n647 VSUBS 0.010909f
C969 B.n648 VSUBS 0.010909f
C970 B.n649 VSUBS 0.010909f
C971 B.n650 VSUBS 0.010909f
C972 B.n651 VSUBS 0.010909f
C973 B.n652 VSUBS 0.010909f
C974 B.n653 VSUBS 0.010909f
C975 B.n654 VSUBS 0.010909f
C976 B.n655 VSUBS 0.010909f
C977 B.n656 VSUBS 0.010909f
C978 B.n657 VSUBS 0.010909f
C979 B.n658 VSUBS 0.010909f
C980 B.n659 VSUBS 0.010909f
C981 B.n660 VSUBS 0.010909f
C982 B.n661 VSUBS 0.010909f
C983 B.n662 VSUBS 0.010909f
C984 B.n663 VSUBS 0.010909f
C985 B.n664 VSUBS 0.010909f
C986 B.n665 VSUBS 0.010909f
C987 B.n666 VSUBS 0.010909f
C988 B.n667 VSUBS 0.010909f
C989 B.n668 VSUBS 0.010909f
C990 B.n669 VSUBS 0.010909f
C991 B.n670 VSUBS 0.010909f
C992 B.n671 VSUBS 0.010909f
C993 B.n672 VSUBS 0.010909f
C994 B.n673 VSUBS 0.010909f
C995 B.n674 VSUBS 0.010909f
C996 B.n675 VSUBS 0.010909f
C997 B.n676 VSUBS 0.010909f
C998 B.n677 VSUBS 0.010909f
C999 B.n678 VSUBS 0.010909f
C1000 B.n679 VSUBS 0.010909f
C1001 B.n680 VSUBS 0.010909f
C1002 B.n681 VSUBS 0.010909f
C1003 B.n682 VSUBS 0.010909f
C1004 B.n683 VSUBS 0.010909f
C1005 B.n684 VSUBS 0.010909f
C1006 B.n685 VSUBS 0.010909f
C1007 B.n686 VSUBS 0.025538f
C1008 B.n687 VSUBS 0.024196f
C1009 B.n688 VSUBS 0.024196f
C1010 B.n689 VSUBS 0.010909f
C1011 B.n690 VSUBS 0.010909f
C1012 B.n691 VSUBS 0.010909f
C1013 B.n692 VSUBS 0.010909f
C1014 B.n693 VSUBS 0.010909f
C1015 B.n694 VSUBS 0.010909f
C1016 B.n695 VSUBS 0.010909f
C1017 B.n696 VSUBS 0.010909f
C1018 B.n697 VSUBS 0.010909f
C1019 B.n698 VSUBS 0.010909f
C1020 B.n699 VSUBS 0.010909f
C1021 B.n700 VSUBS 0.010909f
C1022 B.n701 VSUBS 0.010909f
C1023 B.n702 VSUBS 0.010909f
C1024 B.n703 VSUBS 0.010909f
C1025 B.n704 VSUBS 0.010909f
C1026 B.n705 VSUBS 0.010909f
C1027 B.n706 VSUBS 0.010909f
C1028 B.n707 VSUBS 0.010909f
C1029 B.n708 VSUBS 0.010909f
C1030 B.n709 VSUBS 0.010909f
C1031 B.n710 VSUBS 0.010909f
C1032 B.n711 VSUBS 0.010909f
C1033 B.n712 VSUBS 0.010909f
C1034 B.n713 VSUBS 0.010909f
C1035 B.n714 VSUBS 0.010909f
C1036 B.n715 VSUBS 0.010909f
C1037 B.n716 VSUBS 0.010909f
C1038 B.n717 VSUBS 0.010909f
C1039 B.n718 VSUBS 0.010909f
C1040 B.n719 VSUBS 0.010909f
C1041 B.n720 VSUBS 0.010909f
C1042 B.n721 VSUBS 0.010909f
C1043 B.n722 VSUBS 0.010909f
C1044 B.n723 VSUBS 0.010909f
C1045 B.n724 VSUBS 0.010909f
C1046 B.n725 VSUBS 0.010909f
C1047 B.n726 VSUBS 0.010909f
C1048 B.n727 VSUBS 0.010909f
C1049 B.n728 VSUBS 0.010909f
C1050 B.n729 VSUBS 0.010909f
C1051 B.n730 VSUBS 0.010909f
C1052 B.n731 VSUBS 0.010909f
C1053 B.n732 VSUBS 0.010909f
C1054 B.n733 VSUBS 0.010909f
C1055 B.n734 VSUBS 0.010909f
C1056 B.n735 VSUBS 0.010909f
C1057 B.n736 VSUBS 0.010909f
C1058 B.n737 VSUBS 0.010909f
C1059 B.n738 VSUBS 0.010909f
C1060 B.n739 VSUBS 0.010909f
C1061 B.n740 VSUBS 0.010909f
C1062 B.n741 VSUBS 0.010909f
C1063 B.n742 VSUBS 0.010909f
C1064 B.n743 VSUBS 0.010909f
C1065 B.n744 VSUBS 0.010909f
C1066 B.n745 VSUBS 0.010909f
C1067 B.n746 VSUBS 0.010909f
C1068 B.n747 VSUBS 0.010909f
C1069 B.n748 VSUBS 0.010909f
C1070 B.n749 VSUBS 0.010909f
C1071 B.n750 VSUBS 0.010909f
C1072 B.n751 VSUBS 0.010909f
C1073 B.n752 VSUBS 0.010909f
C1074 B.n753 VSUBS 0.010909f
C1075 B.n754 VSUBS 0.010909f
C1076 B.n755 VSUBS 0.010909f
C1077 B.n756 VSUBS 0.010909f
C1078 B.n757 VSUBS 0.010909f
C1079 B.n758 VSUBS 0.010909f
C1080 B.n759 VSUBS 0.010909f
C1081 B.n760 VSUBS 0.010909f
C1082 B.n761 VSUBS 0.010909f
C1083 B.n762 VSUBS 0.010909f
C1084 B.n763 VSUBS 0.010909f
C1085 B.n764 VSUBS 0.010909f
C1086 B.n765 VSUBS 0.010909f
C1087 B.n766 VSUBS 0.010909f
C1088 B.n767 VSUBS 0.010909f
C1089 B.n768 VSUBS 0.010909f
C1090 B.n769 VSUBS 0.010909f
C1091 B.n770 VSUBS 0.010909f
C1092 B.n771 VSUBS 0.010909f
C1093 B.n772 VSUBS 0.010909f
C1094 B.n773 VSUBS 0.010909f
C1095 B.n774 VSUBS 0.010909f
C1096 B.n775 VSUBS 0.010909f
C1097 B.n776 VSUBS 0.010909f
C1098 B.n777 VSUBS 0.010909f
C1099 B.n778 VSUBS 0.010909f
C1100 B.n779 VSUBS 0.014236f
C1101 B.n780 VSUBS 0.015165f
C1102 B.n781 VSUBS 0.030158f
.ends

