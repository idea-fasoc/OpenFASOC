* NGSPICE file created from diff_pair_sample_1592.ext - technology: sky130A

.subckt diff_pair_sample_1592 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=0 ps=0 w=8.52 l=2.42
X1 VDD1.t5 VP.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=1.4058 ps=8.85 w=8.52 l=2.42
X2 VDD1.t4 VP.t1 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=1.4058 ps=8.85 w=8.52 l=2.42
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=0 ps=0 w=8.52 l=2.42
X4 VTAIL.t5 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=1.4058 ps=8.85 w=8.52 l=2.42
X5 VDD2.t5 VN.t0 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=1.4058 ps=8.85 w=8.52 l=2.42
X6 VDD1.t2 VP.t3 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=3.3228 ps=17.82 w=8.52 l=2.42
X7 VDD2.t4 VN.t1 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=3.3228 ps=17.82 w=8.52 l=2.42
X8 VDD2.t3 VN.t2 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=1.4058 ps=8.85 w=8.52 l=2.42
X9 VDD2.t2 VN.t3 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=3.3228 ps=17.82 w=8.52 l=2.42
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=0 ps=0 w=8.52 l=2.42
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3228 pd=17.82 as=0 ps=0 w=8.52 l=2.42
X12 VTAIL.t7 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=1.4058 ps=8.85 w=8.52 l=2.42
X13 VTAIL.t2 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=1.4058 ps=8.85 w=8.52 l=2.42
X14 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=1.4058 ps=8.85 w=8.52 l=2.42
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4058 pd=8.85 as=3.3228 ps=17.82 w=8.52 l=2.42
R0 B.n695 B.n694 585
R1 B.n257 B.n112 585
R2 B.n256 B.n255 585
R3 B.n254 B.n253 585
R4 B.n252 B.n251 585
R5 B.n250 B.n249 585
R6 B.n248 B.n247 585
R7 B.n246 B.n245 585
R8 B.n244 B.n243 585
R9 B.n242 B.n241 585
R10 B.n240 B.n239 585
R11 B.n238 B.n237 585
R12 B.n236 B.n235 585
R13 B.n234 B.n233 585
R14 B.n232 B.n231 585
R15 B.n230 B.n229 585
R16 B.n228 B.n227 585
R17 B.n226 B.n225 585
R18 B.n224 B.n223 585
R19 B.n222 B.n221 585
R20 B.n220 B.n219 585
R21 B.n218 B.n217 585
R22 B.n216 B.n215 585
R23 B.n214 B.n213 585
R24 B.n212 B.n211 585
R25 B.n210 B.n209 585
R26 B.n208 B.n207 585
R27 B.n206 B.n205 585
R28 B.n204 B.n203 585
R29 B.n202 B.n201 585
R30 B.n200 B.n199 585
R31 B.n197 B.n196 585
R32 B.n195 B.n194 585
R33 B.n193 B.n192 585
R34 B.n191 B.n190 585
R35 B.n189 B.n188 585
R36 B.n187 B.n186 585
R37 B.n185 B.n184 585
R38 B.n183 B.n182 585
R39 B.n181 B.n180 585
R40 B.n179 B.n178 585
R41 B.n176 B.n175 585
R42 B.n174 B.n173 585
R43 B.n172 B.n171 585
R44 B.n170 B.n169 585
R45 B.n168 B.n167 585
R46 B.n166 B.n165 585
R47 B.n164 B.n163 585
R48 B.n162 B.n161 585
R49 B.n160 B.n159 585
R50 B.n158 B.n157 585
R51 B.n156 B.n155 585
R52 B.n154 B.n153 585
R53 B.n152 B.n151 585
R54 B.n150 B.n149 585
R55 B.n148 B.n147 585
R56 B.n146 B.n145 585
R57 B.n144 B.n143 585
R58 B.n142 B.n141 585
R59 B.n140 B.n139 585
R60 B.n138 B.n137 585
R61 B.n136 B.n135 585
R62 B.n134 B.n133 585
R63 B.n132 B.n131 585
R64 B.n130 B.n129 585
R65 B.n128 B.n127 585
R66 B.n126 B.n125 585
R67 B.n124 B.n123 585
R68 B.n122 B.n121 585
R69 B.n120 B.n119 585
R70 B.n118 B.n117 585
R71 B.n75 B.n74 585
R72 B.n693 B.n76 585
R73 B.n698 B.n76 585
R74 B.n692 B.n691 585
R75 B.n691 B.n72 585
R76 B.n690 B.n71 585
R77 B.n704 B.n71 585
R78 B.n689 B.n70 585
R79 B.n705 B.n70 585
R80 B.n688 B.n69 585
R81 B.n706 B.n69 585
R82 B.n687 B.n686 585
R83 B.n686 B.n65 585
R84 B.n685 B.n64 585
R85 B.n712 B.n64 585
R86 B.n684 B.n63 585
R87 B.n713 B.n63 585
R88 B.n683 B.n62 585
R89 B.n714 B.n62 585
R90 B.n682 B.n681 585
R91 B.n681 B.n58 585
R92 B.n680 B.n57 585
R93 B.n720 B.n57 585
R94 B.n679 B.n56 585
R95 B.n721 B.n56 585
R96 B.n678 B.n55 585
R97 B.n722 B.n55 585
R98 B.n677 B.n676 585
R99 B.n676 B.n51 585
R100 B.n675 B.n50 585
R101 B.n728 B.n50 585
R102 B.n674 B.n49 585
R103 B.n729 B.n49 585
R104 B.n673 B.n48 585
R105 B.n730 B.n48 585
R106 B.n672 B.n671 585
R107 B.n671 B.n44 585
R108 B.n670 B.n43 585
R109 B.n736 B.n43 585
R110 B.n669 B.n42 585
R111 B.n737 B.n42 585
R112 B.n668 B.n41 585
R113 B.n738 B.n41 585
R114 B.n667 B.n666 585
R115 B.n666 B.n37 585
R116 B.n665 B.n36 585
R117 B.n744 B.n36 585
R118 B.n664 B.n35 585
R119 B.n745 B.n35 585
R120 B.n663 B.n34 585
R121 B.n746 B.n34 585
R122 B.n662 B.n661 585
R123 B.n661 B.n30 585
R124 B.n660 B.n29 585
R125 B.n752 B.n29 585
R126 B.n659 B.n28 585
R127 B.n753 B.n28 585
R128 B.n658 B.n27 585
R129 B.n754 B.n27 585
R130 B.n657 B.n656 585
R131 B.n656 B.n23 585
R132 B.n655 B.n22 585
R133 B.n760 B.n22 585
R134 B.n654 B.n21 585
R135 B.n761 B.n21 585
R136 B.n653 B.n20 585
R137 B.n762 B.n20 585
R138 B.n652 B.n651 585
R139 B.n651 B.n16 585
R140 B.n650 B.n15 585
R141 B.n768 B.n15 585
R142 B.n649 B.n14 585
R143 B.n769 B.n14 585
R144 B.n648 B.n13 585
R145 B.n770 B.n13 585
R146 B.n647 B.n646 585
R147 B.n646 B.n12 585
R148 B.n645 B.n644 585
R149 B.n645 B.n8 585
R150 B.n643 B.n7 585
R151 B.n777 B.n7 585
R152 B.n642 B.n6 585
R153 B.n778 B.n6 585
R154 B.n641 B.n5 585
R155 B.n779 B.n5 585
R156 B.n640 B.n639 585
R157 B.n639 B.n4 585
R158 B.n638 B.n258 585
R159 B.n638 B.n637 585
R160 B.n628 B.n259 585
R161 B.n260 B.n259 585
R162 B.n630 B.n629 585
R163 B.n631 B.n630 585
R164 B.n627 B.n265 585
R165 B.n265 B.n264 585
R166 B.n626 B.n625 585
R167 B.n625 B.n624 585
R168 B.n267 B.n266 585
R169 B.n268 B.n267 585
R170 B.n617 B.n616 585
R171 B.n618 B.n617 585
R172 B.n615 B.n273 585
R173 B.n273 B.n272 585
R174 B.n614 B.n613 585
R175 B.n613 B.n612 585
R176 B.n275 B.n274 585
R177 B.n276 B.n275 585
R178 B.n605 B.n604 585
R179 B.n606 B.n605 585
R180 B.n603 B.n281 585
R181 B.n281 B.n280 585
R182 B.n602 B.n601 585
R183 B.n601 B.n600 585
R184 B.n283 B.n282 585
R185 B.n284 B.n283 585
R186 B.n593 B.n592 585
R187 B.n594 B.n593 585
R188 B.n591 B.n289 585
R189 B.n289 B.n288 585
R190 B.n590 B.n589 585
R191 B.n589 B.n588 585
R192 B.n291 B.n290 585
R193 B.n292 B.n291 585
R194 B.n581 B.n580 585
R195 B.n582 B.n581 585
R196 B.n579 B.n297 585
R197 B.n297 B.n296 585
R198 B.n578 B.n577 585
R199 B.n577 B.n576 585
R200 B.n299 B.n298 585
R201 B.n300 B.n299 585
R202 B.n569 B.n568 585
R203 B.n570 B.n569 585
R204 B.n567 B.n305 585
R205 B.n305 B.n304 585
R206 B.n566 B.n565 585
R207 B.n565 B.n564 585
R208 B.n307 B.n306 585
R209 B.n308 B.n307 585
R210 B.n557 B.n556 585
R211 B.n558 B.n557 585
R212 B.n555 B.n313 585
R213 B.n313 B.n312 585
R214 B.n554 B.n553 585
R215 B.n553 B.n552 585
R216 B.n315 B.n314 585
R217 B.n316 B.n315 585
R218 B.n545 B.n544 585
R219 B.n546 B.n545 585
R220 B.n543 B.n320 585
R221 B.n324 B.n320 585
R222 B.n542 B.n541 585
R223 B.n541 B.n540 585
R224 B.n322 B.n321 585
R225 B.n323 B.n322 585
R226 B.n533 B.n532 585
R227 B.n534 B.n533 585
R228 B.n531 B.n329 585
R229 B.n329 B.n328 585
R230 B.n530 B.n529 585
R231 B.n529 B.n528 585
R232 B.n331 B.n330 585
R233 B.n332 B.n331 585
R234 B.n521 B.n520 585
R235 B.n522 B.n521 585
R236 B.n335 B.n334 585
R237 B.n380 B.n379 585
R238 B.n381 B.n377 585
R239 B.n377 B.n336 585
R240 B.n383 B.n382 585
R241 B.n385 B.n376 585
R242 B.n388 B.n387 585
R243 B.n389 B.n375 585
R244 B.n391 B.n390 585
R245 B.n393 B.n374 585
R246 B.n396 B.n395 585
R247 B.n397 B.n373 585
R248 B.n399 B.n398 585
R249 B.n401 B.n372 585
R250 B.n404 B.n403 585
R251 B.n405 B.n371 585
R252 B.n407 B.n406 585
R253 B.n409 B.n370 585
R254 B.n412 B.n411 585
R255 B.n413 B.n369 585
R256 B.n415 B.n414 585
R257 B.n417 B.n368 585
R258 B.n420 B.n419 585
R259 B.n421 B.n367 585
R260 B.n423 B.n422 585
R261 B.n425 B.n366 585
R262 B.n428 B.n427 585
R263 B.n429 B.n365 585
R264 B.n431 B.n430 585
R265 B.n433 B.n364 585
R266 B.n436 B.n435 585
R267 B.n437 B.n361 585
R268 B.n440 B.n439 585
R269 B.n442 B.n360 585
R270 B.n445 B.n444 585
R271 B.n446 B.n359 585
R272 B.n448 B.n447 585
R273 B.n450 B.n358 585
R274 B.n453 B.n452 585
R275 B.n454 B.n357 585
R276 B.n456 B.n455 585
R277 B.n458 B.n356 585
R278 B.n461 B.n460 585
R279 B.n462 B.n352 585
R280 B.n464 B.n463 585
R281 B.n466 B.n351 585
R282 B.n469 B.n468 585
R283 B.n470 B.n350 585
R284 B.n472 B.n471 585
R285 B.n474 B.n349 585
R286 B.n477 B.n476 585
R287 B.n478 B.n348 585
R288 B.n480 B.n479 585
R289 B.n482 B.n347 585
R290 B.n485 B.n484 585
R291 B.n486 B.n346 585
R292 B.n488 B.n487 585
R293 B.n490 B.n345 585
R294 B.n493 B.n492 585
R295 B.n494 B.n344 585
R296 B.n496 B.n495 585
R297 B.n498 B.n343 585
R298 B.n501 B.n500 585
R299 B.n502 B.n342 585
R300 B.n504 B.n503 585
R301 B.n506 B.n341 585
R302 B.n509 B.n508 585
R303 B.n510 B.n340 585
R304 B.n512 B.n511 585
R305 B.n514 B.n339 585
R306 B.n515 B.n338 585
R307 B.n518 B.n517 585
R308 B.n519 B.n337 585
R309 B.n337 B.n336 585
R310 B.n524 B.n523 585
R311 B.n523 B.n522 585
R312 B.n525 B.n333 585
R313 B.n333 B.n332 585
R314 B.n527 B.n526 585
R315 B.n528 B.n527 585
R316 B.n327 B.n326 585
R317 B.n328 B.n327 585
R318 B.n536 B.n535 585
R319 B.n535 B.n534 585
R320 B.n537 B.n325 585
R321 B.n325 B.n323 585
R322 B.n539 B.n538 585
R323 B.n540 B.n539 585
R324 B.n319 B.n318 585
R325 B.n324 B.n319 585
R326 B.n548 B.n547 585
R327 B.n547 B.n546 585
R328 B.n549 B.n317 585
R329 B.n317 B.n316 585
R330 B.n551 B.n550 585
R331 B.n552 B.n551 585
R332 B.n311 B.n310 585
R333 B.n312 B.n311 585
R334 B.n560 B.n559 585
R335 B.n559 B.n558 585
R336 B.n561 B.n309 585
R337 B.n309 B.n308 585
R338 B.n563 B.n562 585
R339 B.n564 B.n563 585
R340 B.n303 B.n302 585
R341 B.n304 B.n303 585
R342 B.n572 B.n571 585
R343 B.n571 B.n570 585
R344 B.n573 B.n301 585
R345 B.n301 B.n300 585
R346 B.n575 B.n574 585
R347 B.n576 B.n575 585
R348 B.n295 B.n294 585
R349 B.n296 B.n295 585
R350 B.n584 B.n583 585
R351 B.n583 B.n582 585
R352 B.n585 B.n293 585
R353 B.n293 B.n292 585
R354 B.n587 B.n586 585
R355 B.n588 B.n587 585
R356 B.n287 B.n286 585
R357 B.n288 B.n287 585
R358 B.n596 B.n595 585
R359 B.n595 B.n594 585
R360 B.n597 B.n285 585
R361 B.n285 B.n284 585
R362 B.n599 B.n598 585
R363 B.n600 B.n599 585
R364 B.n279 B.n278 585
R365 B.n280 B.n279 585
R366 B.n608 B.n607 585
R367 B.n607 B.n606 585
R368 B.n609 B.n277 585
R369 B.n277 B.n276 585
R370 B.n611 B.n610 585
R371 B.n612 B.n611 585
R372 B.n271 B.n270 585
R373 B.n272 B.n271 585
R374 B.n620 B.n619 585
R375 B.n619 B.n618 585
R376 B.n621 B.n269 585
R377 B.n269 B.n268 585
R378 B.n623 B.n622 585
R379 B.n624 B.n623 585
R380 B.n263 B.n262 585
R381 B.n264 B.n263 585
R382 B.n633 B.n632 585
R383 B.n632 B.n631 585
R384 B.n634 B.n261 585
R385 B.n261 B.n260 585
R386 B.n636 B.n635 585
R387 B.n637 B.n636 585
R388 B.n3 B.n0 585
R389 B.n4 B.n3 585
R390 B.n776 B.n1 585
R391 B.n777 B.n776 585
R392 B.n775 B.n774 585
R393 B.n775 B.n8 585
R394 B.n773 B.n9 585
R395 B.n12 B.n9 585
R396 B.n772 B.n771 585
R397 B.n771 B.n770 585
R398 B.n11 B.n10 585
R399 B.n769 B.n11 585
R400 B.n767 B.n766 585
R401 B.n768 B.n767 585
R402 B.n765 B.n17 585
R403 B.n17 B.n16 585
R404 B.n764 B.n763 585
R405 B.n763 B.n762 585
R406 B.n19 B.n18 585
R407 B.n761 B.n19 585
R408 B.n759 B.n758 585
R409 B.n760 B.n759 585
R410 B.n757 B.n24 585
R411 B.n24 B.n23 585
R412 B.n756 B.n755 585
R413 B.n755 B.n754 585
R414 B.n26 B.n25 585
R415 B.n753 B.n26 585
R416 B.n751 B.n750 585
R417 B.n752 B.n751 585
R418 B.n749 B.n31 585
R419 B.n31 B.n30 585
R420 B.n748 B.n747 585
R421 B.n747 B.n746 585
R422 B.n33 B.n32 585
R423 B.n745 B.n33 585
R424 B.n743 B.n742 585
R425 B.n744 B.n743 585
R426 B.n741 B.n38 585
R427 B.n38 B.n37 585
R428 B.n740 B.n739 585
R429 B.n739 B.n738 585
R430 B.n40 B.n39 585
R431 B.n737 B.n40 585
R432 B.n735 B.n734 585
R433 B.n736 B.n735 585
R434 B.n733 B.n45 585
R435 B.n45 B.n44 585
R436 B.n732 B.n731 585
R437 B.n731 B.n730 585
R438 B.n47 B.n46 585
R439 B.n729 B.n47 585
R440 B.n727 B.n726 585
R441 B.n728 B.n727 585
R442 B.n725 B.n52 585
R443 B.n52 B.n51 585
R444 B.n724 B.n723 585
R445 B.n723 B.n722 585
R446 B.n54 B.n53 585
R447 B.n721 B.n54 585
R448 B.n719 B.n718 585
R449 B.n720 B.n719 585
R450 B.n717 B.n59 585
R451 B.n59 B.n58 585
R452 B.n716 B.n715 585
R453 B.n715 B.n714 585
R454 B.n61 B.n60 585
R455 B.n713 B.n61 585
R456 B.n711 B.n710 585
R457 B.n712 B.n711 585
R458 B.n709 B.n66 585
R459 B.n66 B.n65 585
R460 B.n708 B.n707 585
R461 B.n707 B.n706 585
R462 B.n68 B.n67 585
R463 B.n705 B.n68 585
R464 B.n703 B.n702 585
R465 B.n704 B.n703 585
R466 B.n701 B.n73 585
R467 B.n73 B.n72 585
R468 B.n700 B.n699 585
R469 B.n699 B.n698 585
R470 B.n780 B.n779 585
R471 B.n778 B.n2 585
R472 B.n699 B.n75 521.33
R473 B.n695 B.n76 521.33
R474 B.n521 B.n337 521.33
R475 B.n523 B.n335 521.33
R476 B.n115 B.t14 292.606
R477 B.n113 B.t10 292.606
R478 B.n353 B.t6 292.606
R479 B.n362 B.t17 292.606
R480 B.n113 B.t12 275.231
R481 B.n353 B.t9 275.231
R482 B.n115 B.t15 275.231
R483 B.n362 B.t19 275.231
R484 B.n697 B.n696 256.663
R485 B.n697 B.n111 256.663
R486 B.n697 B.n110 256.663
R487 B.n697 B.n109 256.663
R488 B.n697 B.n108 256.663
R489 B.n697 B.n107 256.663
R490 B.n697 B.n106 256.663
R491 B.n697 B.n105 256.663
R492 B.n697 B.n104 256.663
R493 B.n697 B.n103 256.663
R494 B.n697 B.n102 256.663
R495 B.n697 B.n101 256.663
R496 B.n697 B.n100 256.663
R497 B.n697 B.n99 256.663
R498 B.n697 B.n98 256.663
R499 B.n697 B.n97 256.663
R500 B.n697 B.n96 256.663
R501 B.n697 B.n95 256.663
R502 B.n697 B.n94 256.663
R503 B.n697 B.n93 256.663
R504 B.n697 B.n92 256.663
R505 B.n697 B.n91 256.663
R506 B.n697 B.n90 256.663
R507 B.n697 B.n89 256.663
R508 B.n697 B.n88 256.663
R509 B.n697 B.n87 256.663
R510 B.n697 B.n86 256.663
R511 B.n697 B.n85 256.663
R512 B.n697 B.n84 256.663
R513 B.n697 B.n83 256.663
R514 B.n697 B.n82 256.663
R515 B.n697 B.n81 256.663
R516 B.n697 B.n80 256.663
R517 B.n697 B.n79 256.663
R518 B.n697 B.n78 256.663
R519 B.n697 B.n77 256.663
R520 B.n378 B.n336 256.663
R521 B.n384 B.n336 256.663
R522 B.n386 B.n336 256.663
R523 B.n392 B.n336 256.663
R524 B.n394 B.n336 256.663
R525 B.n400 B.n336 256.663
R526 B.n402 B.n336 256.663
R527 B.n408 B.n336 256.663
R528 B.n410 B.n336 256.663
R529 B.n416 B.n336 256.663
R530 B.n418 B.n336 256.663
R531 B.n424 B.n336 256.663
R532 B.n426 B.n336 256.663
R533 B.n432 B.n336 256.663
R534 B.n434 B.n336 256.663
R535 B.n441 B.n336 256.663
R536 B.n443 B.n336 256.663
R537 B.n449 B.n336 256.663
R538 B.n451 B.n336 256.663
R539 B.n457 B.n336 256.663
R540 B.n459 B.n336 256.663
R541 B.n465 B.n336 256.663
R542 B.n467 B.n336 256.663
R543 B.n473 B.n336 256.663
R544 B.n475 B.n336 256.663
R545 B.n481 B.n336 256.663
R546 B.n483 B.n336 256.663
R547 B.n489 B.n336 256.663
R548 B.n491 B.n336 256.663
R549 B.n497 B.n336 256.663
R550 B.n499 B.n336 256.663
R551 B.n505 B.n336 256.663
R552 B.n507 B.n336 256.663
R553 B.n513 B.n336 256.663
R554 B.n516 B.n336 256.663
R555 B.n782 B.n781 256.663
R556 B.n114 B.t13 221.898
R557 B.n354 B.t8 221.898
R558 B.n116 B.t16 221.898
R559 B.n363 B.t18 221.898
R560 B.n119 B.n118 163.367
R561 B.n123 B.n122 163.367
R562 B.n127 B.n126 163.367
R563 B.n131 B.n130 163.367
R564 B.n135 B.n134 163.367
R565 B.n139 B.n138 163.367
R566 B.n143 B.n142 163.367
R567 B.n147 B.n146 163.367
R568 B.n151 B.n150 163.367
R569 B.n155 B.n154 163.367
R570 B.n159 B.n158 163.367
R571 B.n163 B.n162 163.367
R572 B.n167 B.n166 163.367
R573 B.n171 B.n170 163.367
R574 B.n175 B.n174 163.367
R575 B.n180 B.n179 163.367
R576 B.n184 B.n183 163.367
R577 B.n188 B.n187 163.367
R578 B.n192 B.n191 163.367
R579 B.n196 B.n195 163.367
R580 B.n201 B.n200 163.367
R581 B.n205 B.n204 163.367
R582 B.n209 B.n208 163.367
R583 B.n213 B.n212 163.367
R584 B.n217 B.n216 163.367
R585 B.n221 B.n220 163.367
R586 B.n225 B.n224 163.367
R587 B.n229 B.n228 163.367
R588 B.n233 B.n232 163.367
R589 B.n237 B.n236 163.367
R590 B.n241 B.n240 163.367
R591 B.n245 B.n244 163.367
R592 B.n249 B.n248 163.367
R593 B.n253 B.n252 163.367
R594 B.n255 B.n112 163.367
R595 B.n521 B.n331 163.367
R596 B.n529 B.n331 163.367
R597 B.n529 B.n329 163.367
R598 B.n533 B.n329 163.367
R599 B.n533 B.n322 163.367
R600 B.n541 B.n322 163.367
R601 B.n541 B.n320 163.367
R602 B.n545 B.n320 163.367
R603 B.n545 B.n315 163.367
R604 B.n553 B.n315 163.367
R605 B.n553 B.n313 163.367
R606 B.n557 B.n313 163.367
R607 B.n557 B.n307 163.367
R608 B.n565 B.n307 163.367
R609 B.n565 B.n305 163.367
R610 B.n569 B.n305 163.367
R611 B.n569 B.n299 163.367
R612 B.n577 B.n299 163.367
R613 B.n577 B.n297 163.367
R614 B.n581 B.n297 163.367
R615 B.n581 B.n291 163.367
R616 B.n589 B.n291 163.367
R617 B.n589 B.n289 163.367
R618 B.n593 B.n289 163.367
R619 B.n593 B.n283 163.367
R620 B.n601 B.n283 163.367
R621 B.n601 B.n281 163.367
R622 B.n605 B.n281 163.367
R623 B.n605 B.n275 163.367
R624 B.n613 B.n275 163.367
R625 B.n613 B.n273 163.367
R626 B.n617 B.n273 163.367
R627 B.n617 B.n267 163.367
R628 B.n625 B.n267 163.367
R629 B.n625 B.n265 163.367
R630 B.n630 B.n265 163.367
R631 B.n630 B.n259 163.367
R632 B.n638 B.n259 163.367
R633 B.n639 B.n638 163.367
R634 B.n639 B.n5 163.367
R635 B.n6 B.n5 163.367
R636 B.n7 B.n6 163.367
R637 B.n645 B.n7 163.367
R638 B.n646 B.n645 163.367
R639 B.n646 B.n13 163.367
R640 B.n14 B.n13 163.367
R641 B.n15 B.n14 163.367
R642 B.n651 B.n15 163.367
R643 B.n651 B.n20 163.367
R644 B.n21 B.n20 163.367
R645 B.n22 B.n21 163.367
R646 B.n656 B.n22 163.367
R647 B.n656 B.n27 163.367
R648 B.n28 B.n27 163.367
R649 B.n29 B.n28 163.367
R650 B.n661 B.n29 163.367
R651 B.n661 B.n34 163.367
R652 B.n35 B.n34 163.367
R653 B.n36 B.n35 163.367
R654 B.n666 B.n36 163.367
R655 B.n666 B.n41 163.367
R656 B.n42 B.n41 163.367
R657 B.n43 B.n42 163.367
R658 B.n671 B.n43 163.367
R659 B.n671 B.n48 163.367
R660 B.n49 B.n48 163.367
R661 B.n50 B.n49 163.367
R662 B.n676 B.n50 163.367
R663 B.n676 B.n55 163.367
R664 B.n56 B.n55 163.367
R665 B.n57 B.n56 163.367
R666 B.n681 B.n57 163.367
R667 B.n681 B.n62 163.367
R668 B.n63 B.n62 163.367
R669 B.n64 B.n63 163.367
R670 B.n686 B.n64 163.367
R671 B.n686 B.n69 163.367
R672 B.n70 B.n69 163.367
R673 B.n71 B.n70 163.367
R674 B.n691 B.n71 163.367
R675 B.n691 B.n76 163.367
R676 B.n379 B.n377 163.367
R677 B.n383 B.n377 163.367
R678 B.n387 B.n385 163.367
R679 B.n391 B.n375 163.367
R680 B.n395 B.n393 163.367
R681 B.n399 B.n373 163.367
R682 B.n403 B.n401 163.367
R683 B.n407 B.n371 163.367
R684 B.n411 B.n409 163.367
R685 B.n415 B.n369 163.367
R686 B.n419 B.n417 163.367
R687 B.n423 B.n367 163.367
R688 B.n427 B.n425 163.367
R689 B.n431 B.n365 163.367
R690 B.n435 B.n433 163.367
R691 B.n440 B.n361 163.367
R692 B.n444 B.n442 163.367
R693 B.n448 B.n359 163.367
R694 B.n452 B.n450 163.367
R695 B.n456 B.n357 163.367
R696 B.n460 B.n458 163.367
R697 B.n464 B.n352 163.367
R698 B.n468 B.n466 163.367
R699 B.n472 B.n350 163.367
R700 B.n476 B.n474 163.367
R701 B.n480 B.n348 163.367
R702 B.n484 B.n482 163.367
R703 B.n488 B.n346 163.367
R704 B.n492 B.n490 163.367
R705 B.n496 B.n344 163.367
R706 B.n500 B.n498 163.367
R707 B.n504 B.n342 163.367
R708 B.n508 B.n506 163.367
R709 B.n512 B.n340 163.367
R710 B.n515 B.n514 163.367
R711 B.n517 B.n337 163.367
R712 B.n523 B.n333 163.367
R713 B.n527 B.n333 163.367
R714 B.n527 B.n327 163.367
R715 B.n535 B.n327 163.367
R716 B.n535 B.n325 163.367
R717 B.n539 B.n325 163.367
R718 B.n539 B.n319 163.367
R719 B.n547 B.n319 163.367
R720 B.n547 B.n317 163.367
R721 B.n551 B.n317 163.367
R722 B.n551 B.n311 163.367
R723 B.n559 B.n311 163.367
R724 B.n559 B.n309 163.367
R725 B.n563 B.n309 163.367
R726 B.n563 B.n303 163.367
R727 B.n571 B.n303 163.367
R728 B.n571 B.n301 163.367
R729 B.n575 B.n301 163.367
R730 B.n575 B.n295 163.367
R731 B.n583 B.n295 163.367
R732 B.n583 B.n293 163.367
R733 B.n587 B.n293 163.367
R734 B.n587 B.n287 163.367
R735 B.n595 B.n287 163.367
R736 B.n595 B.n285 163.367
R737 B.n599 B.n285 163.367
R738 B.n599 B.n279 163.367
R739 B.n607 B.n279 163.367
R740 B.n607 B.n277 163.367
R741 B.n611 B.n277 163.367
R742 B.n611 B.n271 163.367
R743 B.n619 B.n271 163.367
R744 B.n619 B.n269 163.367
R745 B.n623 B.n269 163.367
R746 B.n623 B.n263 163.367
R747 B.n632 B.n263 163.367
R748 B.n632 B.n261 163.367
R749 B.n636 B.n261 163.367
R750 B.n636 B.n3 163.367
R751 B.n780 B.n3 163.367
R752 B.n776 B.n2 163.367
R753 B.n776 B.n775 163.367
R754 B.n775 B.n9 163.367
R755 B.n771 B.n9 163.367
R756 B.n771 B.n11 163.367
R757 B.n767 B.n11 163.367
R758 B.n767 B.n17 163.367
R759 B.n763 B.n17 163.367
R760 B.n763 B.n19 163.367
R761 B.n759 B.n19 163.367
R762 B.n759 B.n24 163.367
R763 B.n755 B.n24 163.367
R764 B.n755 B.n26 163.367
R765 B.n751 B.n26 163.367
R766 B.n751 B.n31 163.367
R767 B.n747 B.n31 163.367
R768 B.n747 B.n33 163.367
R769 B.n743 B.n33 163.367
R770 B.n743 B.n38 163.367
R771 B.n739 B.n38 163.367
R772 B.n739 B.n40 163.367
R773 B.n735 B.n40 163.367
R774 B.n735 B.n45 163.367
R775 B.n731 B.n45 163.367
R776 B.n731 B.n47 163.367
R777 B.n727 B.n47 163.367
R778 B.n727 B.n52 163.367
R779 B.n723 B.n52 163.367
R780 B.n723 B.n54 163.367
R781 B.n719 B.n54 163.367
R782 B.n719 B.n59 163.367
R783 B.n715 B.n59 163.367
R784 B.n715 B.n61 163.367
R785 B.n711 B.n61 163.367
R786 B.n711 B.n66 163.367
R787 B.n707 B.n66 163.367
R788 B.n707 B.n68 163.367
R789 B.n703 B.n68 163.367
R790 B.n703 B.n73 163.367
R791 B.n699 B.n73 163.367
R792 B.n522 B.n336 96.4847
R793 B.n698 B.n697 96.4847
R794 B.n77 B.n75 71.676
R795 B.n119 B.n78 71.676
R796 B.n123 B.n79 71.676
R797 B.n127 B.n80 71.676
R798 B.n131 B.n81 71.676
R799 B.n135 B.n82 71.676
R800 B.n139 B.n83 71.676
R801 B.n143 B.n84 71.676
R802 B.n147 B.n85 71.676
R803 B.n151 B.n86 71.676
R804 B.n155 B.n87 71.676
R805 B.n159 B.n88 71.676
R806 B.n163 B.n89 71.676
R807 B.n167 B.n90 71.676
R808 B.n171 B.n91 71.676
R809 B.n175 B.n92 71.676
R810 B.n180 B.n93 71.676
R811 B.n184 B.n94 71.676
R812 B.n188 B.n95 71.676
R813 B.n192 B.n96 71.676
R814 B.n196 B.n97 71.676
R815 B.n201 B.n98 71.676
R816 B.n205 B.n99 71.676
R817 B.n209 B.n100 71.676
R818 B.n213 B.n101 71.676
R819 B.n217 B.n102 71.676
R820 B.n221 B.n103 71.676
R821 B.n225 B.n104 71.676
R822 B.n229 B.n105 71.676
R823 B.n233 B.n106 71.676
R824 B.n237 B.n107 71.676
R825 B.n241 B.n108 71.676
R826 B.n245 B.n109 71.676
R827 B.n249 B.n110 71.676
R828 B.n253 B.n111 71.676
R829 B.n696 B.n112 71.676
R830 B.n696 B.n695 71.676
R831 B.n255 B.n111 71.676
R832 B.n252 B.n110 71.676
R833 B.n248 B.n109 71.676
R834 B.n244 B.n108 71.676
R835 B.n240 B.n107 71.676
R836 B.n236 B.n106 71.676
R837 B.n232 B.n105 71.676
R838 B.n228 B.n104 71.676
R839 B.n224 B.n103 71.676
R840 B.n220 B.n102 71.676
R841 B.n216 B.n101 71.676
R842 B.n212 B.n100 71.676
R843 B.n208 B.n99 71.676
R844 B.n204 B.n98 71.676
R845 B.n200 B.n97 71.676
R846 B.n195 B.n96 71.676
R847 B.n191 B.n95 71.676
R848 B.n187 B.n94 71.676
R849 B.n183 B.n93 71.676
R850 B.n179 B.n92 71.676
R851 B.n174 B.n91 71.676
R852 B.n170 B.n90 71.676
R853 B.n166 B.n89 71.676
R854 B.n162 B.n88 71.676
R855 B.n158 B.n87 71.676
R856 B.n154 B.n86 71.676
R857 B.n150 B.n85 71.676
R858 B.n146 B.n84 71.676
R859 B.n142 B.n83 71.676
R860 B.n138 B.n82 71.676
R861 B.n134 B.n81 71.676
R862 B.n130 B.n80 71.676
R863 B.n126 B.n79 71.676
R864 B.n122 B.n78 71.676
R865 B.n118 B.n77 71.676
R866 B.n378 B.n335 71.676
R867 B.n384 B.n383 71.676
R868 B.n387 B.n386 71.676
R869 B.n392 B.n391 71.676
R870 B.n395 B.n394 71.676
R871 B.n400 B.n399 71.676
R872 B.n403 B.n402 71.676
R873 B.n408 B.n407 71.676
R874 B.n411 B.n410 71.676
R875 B.n416 B.n415 71.676
R876 B.n419 B.n418 71.676
R877 B.n424 B.n423 71.676
R878 B.n427 B.n426 71.676
R879 B.n432 B.n431 71.676
R880 B.n435 B.n434 71.676
R881 B.n441 B.n440 71.676
R882 B.n444 B.n443 71.676
R883 B.n449 B.n448 71.676
R884 B.n452 B.n451 71.676
R885 B.n457 B.n456 71.676
R886 B.n460 B.n459 71.676
R887 B.n465 B.n464 71.676
R888 B.n468 B.n467 71.676
R889 B.n473 B.n472 71.676
R890 B.n476 B.n475 71.676
R891 B.n481 B.n480 71.676
R892 B.n484 B.n483 71.676
R893 B.n489 B.n488 71.676
R894 B.n492 B.n491 71.676
R895 B.n497 B.n496 71.676
R896 B.n500 B.n499 71.676
R897 B.n505 B.n504 71.676
R898 B.n508 B.n507 71.676
R899 B.n513 B.n512 71.676
R900 B.n516 B.n515 71.676
R901 B.n379 B.n378 71.676
R902 B.n385 B.n384 71.676
R903 B.n386 B.n375 71.676
R904 B.n393 B.n392 71.676
R905 B.n394 B.n373 71.676
R906 B.n401 B.n400 71.676
R907 B.n402 B.n371 71.676
R908 B.n409 B.n408 71.676
R909 B.n410 B.n369 71.676
R910 B.n417 B.n416 71.676
R911 B.n418 B.n367 71.676
R912 B.n425 B.n424 71.676
R913 B.n426 B.n365 71.676
R914 B.n433 B.n432 71.676
R915 B.n434 B.n361 71.676
R916 B.n442 B.n441 71.676
R917 B.n443 B.n359 71.676
R918 B.n450 B.n449 71.676
R919 B.n451 B.n357 71.676
R920 B.n458 B.n457 71.676
R921 B.n459 B.n352 71.676
R922 B.n466 B.n465 71.676
R923 B.n467 B.n350 71.676
R924 B.n474 B.n473 71.676
R925 B.n475 B.n348 71.676
R926 B.n482 B.n481 71.676
R927 B.n483 B.n346 71.676
R928 B.n490 B.n489 71.676
R929 B.n491 B.n344 71.676
R930 B.n498 B.n497 71.676
R931 B.n499 B.n342 71.676
R932 B.n506 B.n505 71.676
R933 B.n507 B.n340 71.676
R934 B.n514 B.n513 71.676
R935 B.n517 B.n516 71.676
R936 B.n781 B.n780 71.676
R937 B.n781 B.n2 71.676
R938 B.n177 B.n116 59.5399
R939 B.n198 B.n114 59.5399
R940 B.n355 B.n354 59.5399
R941 B.n438 B.n363 59.5399
R942 B.n522 B.n332 54.223
R943 B.n528 B.n332 54.223
R944 B.n528 B.n328 54.223
R945 B.n534 B.n328 54.223
R946 B.n534 B.n323 54.223
R947 B.n540 B.n323 54.223
R948 B.n540 B.n324 54.223
R949 B.n546 B.n316 54.223
R950 B.n552 B.n316 54.223
R951 B.n552 B.n312 54.223
R952 B.n558 B.n312 54.223
R953 B.n558 B.n308 54.223
R954 B.n564 B.n308 54.223
R955 B.n564 B.n304 54.223
R956 B.n570 B.n304 54.223
R957 B.n570 B.n300 54.223
R958 B.n576 B.n300 54.223
R959 B.n582 B.n296 54.223
R960 B.n582 B.n292 54.223
R961 B.n588 B.n292 54.223
R962 B.n588 B.n288 54.223
R963 B.n594 B.n288 54.223
R964 B.n594 B.n284 54.223
R965 B.n600 B.n284 54.223
R966 B.n606 B.n280 54.223
R967 B.n606 B.n276 54.223
R968 B.n612 B.n276 54.223
R969 B.n612 B.n272 54.223
R970 B.n618 B.n272 54.223
R971 B.n618 B.n268 54.223
R972 B.n624 B.n268 54.223
R973 B.n631 B.n264 54.223
R974 B.n631 B.n260 54.223
R975 B.n637 B.n260 54.223
R976 B.n637 B.n4 54.223
R977 B.n779 B.n4 54.223
R978 B.n779 B.n778 54.223
R979 B.n778 B.n777 54.223
R980 B.n777 B.n8 54.223
R981 B.n12 B.n8 54.223
R982 B.n770 B.n12 54.223
R983 B.n770 B.n769 54.223
R984 B.n768 B.n16 54.223
R985 B.n762 B.n16 54.223
R986 B.n762 B.n761 54.223
R987 B.n761 B.n760 54.223
R988 B.n760 B.n23 54.223
R989 B.n754 B.n23 54.223
R990 B.n754 B.n753 54.223
R991 B.n752 B.n30 54.223
R992 B.n746 B.n30 54.223
R993 B.n746 B.n745 54.223
R994 B.n745 B.n744 54.223
R995 B.n744 B.n37 54.223
R996 B.n738 B.n37 54.223
R997 B.n738 B.n737 54.223
R998 B.n736 B.n44 54.223
R999 B.n730 B.n44 54.223
R1000 B.n730 B.n729 54.223
R1001 B.n729 B.n728 54.223
R1002 B.n728 B.n51 54.223
R1003 B.n722 B.n51 54.223
R1004 B.n722 B.n721 54.223
R1005 B.n721 B.n720 54.223
R1006 B.n720 B.n58 54.223
R1007 B.n714 B.n58 54.223
R1008 B.n713 B.n712 54.223
R1009 B.n712 B.n65 54.223
R1010 B.n706 B.n65 54.223
R1011 B.n706 B.n705 54.223
R1012 B.n705 B.n704 54.223
R1013 B.n704 B.n72 54.223
R1014 B.n698 B.n72 54.223
R1015 B.n116 B.n115 53.3338
R1016 B.n114 B.n113 53.3338
R1017 B.n354 B.n353 53.3338
R1018 B.n363 B.n362 53.3338
R1019 B.n624 B.t1 46.2491
R1020 B.t2 B.n768 46.2491
R1021 B.n600 B.t4 41.4648
R1022 B.t0 B.n752 41.4648
R1023 B.n576 B.t5 36.6805
R1024 B.t3 B.n736 36.6805
R1025 B.n524 B.n334 33.8737
R1026 B.n520 B.n519 33.8737
R1027 B.n694 B.n693 33.8737
R1028 B.n700 B.n74 33.8737
R1029 B.n546 B.t7 33.4909
R1030 B.n714 B.t11 33.4909
R1031 B.n324 B.t7 20.7326
R1032 B.t11 B.n713 20.7326
R1033 B B.n782 18.0485
R1034 B.t5 B.n296 17.5431
R1035 B.n737 B.t3 17.5431
R1036 B.t4 B.n280 12.7587
R1037 B.n753 B.t0 12.7587
R1038 B.n525 B.n524 10.6151
R1039 B.n526 B.n525 10.6151
R1040 B.n526 B.n326 10.6151
R1041 B.n536 B.n326 10.6151
R1042 B.n537 B.n536 10.6151
R1043 B.n538 B.n537 10.6151
R1044 B.n538 B.n318 10.6151
R1045 B.n548 B.n318 10.6151
R1046 B.n549 B.n548 10.6151
R1047 B.n550 B.n549 10.6151
R1048 B.n550 B.n310 10.6151
R1049 B.n560 B.n310 10.6151
R1050 B.n561 B.n560 10.6151
R1051 B.n562 B.n561 10.6151
R1052 B.n562 B.n302 10.6151
R1053 B.n572 B.n302 10.6151
R1054 B.n573 B.n572 10.6151
R1055 B.n574 B.n573 10.6151
R1056 B.n574 B.n294 10.6151
R1057 B.n584 B.n294 10.6151
R1058 B.n585 B.n584 10.6151
R1059 B.n586 B.n585 10.6151
R1060 B.n586 B.n286 10.6151
R1061 B.n596 B.n286 10.6151
R1062 B.n597 B.n596 10.6151
R1063 B.n598 B.n597 10.6151
R1064 B.n598 B.n278 10.6151
R1065 B.n608 B.n278 10.6151
R1066 B.n609 B.n608 10.6151
R1067 B.n610 B.n609 10.6151
R1068 B.n610 B.n270 10.6151
R1069 B.n620 B.n270 10.6151
R1070 B.n621 B.n620 10.6151
R1071 B.n622 B.n621 10.6151
R1072 B.n622 B.n262 10.6151
R1073 B.n633 B.n262 10.6151
R1074 B.n634 B.n633 10.6151
R1075 B.n635 B.n634 10.6151
R1076 B.n635 B.n0 10.6151
R1077 B.n380 B.n334 10.6151
R1078 B.n381 B.n380 10.6151
R1079 B.n382 B.n381 10.6151
R1080 B.n382 B.n376 10.6151
R1081 B.n388 B.n376 10.6151
R1082 B.n389 B.n388 10.6151
R1083 B.n390 B.n389 10.6151
R1084 B.n390 B.n374 10.6151
R1085 B.n396 B.n374 10.6151
R1086 B.n397 B.n396 10.6151
R1087 B.n398 B.n397 10.6151
R1088 B.n398 B.n372 10.6151
R1089 B.n404 B.n372 10.6151
R1090 B.n405 B.n404 10.6151
R1091 B.n406 B.n405 10.6151
R1092 B.n406 B.n370 10.6151
R1093 B.n412 B.n370 10.6151
R1094 B.n413 B.n412 10.6151
R1095 B.n414 B.n413 10.6151
R1096 B.n414 B.n368 10.6151
R1097 B.n420 B.n368 10.6151
R1098 B.n421 B.n420 10.6151
R1099 B.n422 B.n421 10.6151
R1100 B.n422 B.n366 10.6151
R1101 B.n428 B.n366 10.6151
R1102 B.n429 B.n428 10.6151
R1103 B.n430 B.n429 10.6151
R1104 B.n430 B.n364 10.6151
R1105 B.n436 B.n364 10.6151
R1106 B.n437 B.n436 10.6151
R1107 B.n439 B.n360 10.6151
R1108 B.n445 B.n360 10.6151
R1109 B.n446 B.n445 10.6151
R1110 B.n447 B.n446 10.6151
R1111 B.n447 B.n358 10.6151
R1112 B.n453 B.n358 10.6151
R1113 B.n454 B.n453 10.6151
R1114 B.n455 B.n454 10.6151
R1115 B.n455 B.n356 10.6151
R1116 B.n462 B.n461 10.6151
R1117 B.n463 B.n462 10.6151
R1118 B.n463 B.n351 10.6151
R1119 B.n469 B.n351 10.6151
R1120 B.n470 B.n469 10.6151
R1121 B.n471 B.n470 10.6151
R1122 B.n471 B.n349 10.6151
R1123 B.n477 B.n349 10.6151
R1124 B.n478 B.n477 10.6151
R1125 B.n479 B.n478 10.6151
R1126 B.n479 B.n347 10.6151
R1127 B.n485 B.n347 10.6151
R1128 B.n486 B.n485 10.6151
R1129 B.n487 B.n486 10.6151
R1130 B.n487 B.n345 10.6151
R1131 B.n493 B.n345 10.6151
R1132 B.n494 B.n493 10.6151
R1133 B.n495 B.n494 10.6151
R1134 B.n495 B.n343 10.6151
R1135 B.n501 B.n343 10.6151
R1136 B.n502 B.n501 10.6151
R1137 B.n503 B.n502 10.6151
R1138 B.n503 B.n341 10.6151
R1139 B.n509 B.n341 10.6151
R1140 B.n510 B.n509 10.6151
R1141 B.n511 B.n510 10.6151
R1142 B.n511 B.n339 10.6151
R1143 B.n339 B.n338 10.6151
R1144 B.n518 B.n338 10.6151
R1145 B.n519 B.n518 10.6151
R1146 B.n520 B.n330 10.6151
R1147 B.n530 B.n330 10.6151
R1148 B.n531 B.n530 10.6151
R1149 B.n532 B.n531 10.6151
R1150 B.n532 B.n321 10.6151
R1151 B.n542 B.n321 10.6151
R1152 B.n543 B.n542 10.6151
R1153 B.n544 B.n543 10.6151
R1154 B.n544 B.n314 10.6151
R1155 B.n554 B.n314 10.6151
R1156 B.n555 B.n554 10.6151
R1157 B.n556 B.n555 10.6151
R1158 B.n556 B.n306 10.6151
R1159 B.n566 B.n306 10.6151
R1160 B.n567 B.n566 10.6151
R1161 B.n568 B.n567 10.6151
R1162 B.n568 B.n298 10.6151
R1163 B.n578 B.n298 10.6151
R1164 B.n579 B.n578 10.6151
R1165 B.n580 B.n579 10.6151
R1166 B.n580 B.n290 10.6151
R1167 B.n590 B.n290 10.6151
R1168 B.n591 B.n590 10.6151
R1169 B.n592 B.n591 10.6151
R1170 B.n592 B.n282 10.6151
R1171 B.n602 B.n282 10.6151
R1172 B.n603 B.n602 10.6151
R1173 B.n604 B.n603 10.6151
R1174 B.n604 B.n274 10.6151
R1175 B.n614 B.n274 10.6151
R1176 B.n615 B.n614 10.6151
R1177 B.n616 B.n615 10.6151
R1178 B.n616 B.n266 10.6151
R1179 B.n626 B.n266 10.6151
R1180 B.n627 B.n626 10.6151
R1181 B.n629 B.n627 10.6151
R1182 B.n629 B.n628 10.6151
R1183 B.n628 B.n258 10.6151
R1184 B.n640 B.n258 10.6151
R1185 B.n641 B.n640 10.6151
R1186 B.n642 B.n641 10.6151
R1187 B.n643 B.n642 10.6151
R1188 B.n644 B.n643 10.6151
R1189 B.n647 B.n644 10.6151
R1190 B.n648 B.n647 10.6151
R1191 B.n649 B.n648 10.6151
R1192 B.n650 B.n649 10.6151
R1193 B.n652 B.n650 10.6151
R1194 B.n653 B.n652 10.6151
R1195 B.n654 B.n653 10.6151
R1196 B.n655 B.n654 10.6151
R1197 B.n657 B.n655 10.6151
R1198 B.n658 B.n657 10.6151
R1199 B.n659 B.n658 10.6151
R1200 B.n660 B.n659 10.6151
R1201 B.n662 B.n660 10.6151
R1202 B.n663 B.n662 10.6151
R1203 B.n664 B.n663 10.6151
R1204 B.n665 B.n664 10.6151
R1205 B.n667 B.n665 10.6151
R1206 B.n668 B.n667 10.6151
R1207 B.n669 B.n668 10.6151
R1208 B.n670 B.n669 10.6151
R1209 B.n672 B.n670 10.6151
R1210 B.n673 B.n672 10.6151
R1211 B.n674 B.n673 10.6151
R1212 B.n675 B.n674 10.6151
R1213 B.n677 B.n675 10.6151
R1214 B.n678 B.n677 10.6151
R1215 B.n679 B.n678 10.6151
R1216 B.n680 B.n679 10.6151
R1217 B.n682 B.n680 10.6151
R1218 B.n683 B.n682 10.6151
R1219 B.n684 B.n683 10.6151
R1220 B.n685 B.n684 10.6151
R1221 B.n687 B.n685 10.6151
R1222 B.n688 B.n687 10.6151
R1223 B.n689 B.n688 10.6151
R1224 B.n690 B.n689 10.6151
R1225 B.n692 B.n690 10.6151
R1226 B.n693 B.n692 10.6151
R1227 B.n774 B.n1 10.6151
R1228 B.n774 B.n773 10.6151
R1229 B.n773 B.n772 10.6151
R1230 B.n772 B.n10 10.6151
R1231 B.n766 B.n10 10.6151
R1232 B.n766 B.n765 10.6151
R1233 B.n765 B.n764 10.6151
R1234 B.n764 B.n18 10.6151
R1235 B.n758 B.n18 10.6151
R1236 B.n758 B.n757 10.6151
R1237 B.n757 B.n756 10.6151
R1238 B.n756 B.n25 10.6151
R1239 B.n750 B.n25 10.6151
R1240 B.n750 B.n749 10.6151
R1241 B.n749 B.n748 10.6151
R1242 B.n748 B.n32 10.6151
R1243 B.n742 B.n32 10.6151
R1244 B.n742 B.n741 10.6151
R1245 B.n741 B.n740 10.6151
R1246 B.n740 B.n39 10.6151
R1247 B.n734 B.n39 10.6151
R1248 B.n734 B.n733 10.6151
R1249 B.n733 B.n732 10.6151
R1250 B.n732 B.n46 10.6151
R1251 B.n726 B.n46 10.6151
R1252 B.n726 B.n725 10.6151
R1253 B.n725 B.n724 10.6151
R1254 B.n724 B.n53 10.6151
R1255 B.n718 B.n53 10.6151
R1256 B.n718 B.n717 10.6151
R1257 B.n717 B.n716 10.6151
R1258 B.n716 B.n60 10.6151
R1259 B.n710 B.n60 10.6151
R1260 B.n710 B.n709 10.6151
R1261 B.n709 B.n708 10.6151
R1262 B.n708 B.n67 10.6151
R1263 B.n702 B.n67 10.6151
R1264 B.n702 B.n701 10.6151
R1265 B.n701 B.n700 10.6151
R1266 B.n117 B.n74 10.6151
R1267 B.n120 B.n117 10.6151
R1268 B.n121 B.n120 10.6151
R1269 B.n124 B.n121 10.6151
R1270 B.n125 B.n124 10.6151
R1271 B.n128 B.n125 10.6151
R1272 B.n129 B.n128 10.6151
R1273 B.n132 B.n129 10.6151
R1274 B.n133 B.n132 10.6151
R1275 B.n136 B.n133 10.6151
R1276 B.n137 B.n136 10.6151
R1277 B.n140 B.n137 10.6151
R1278 B.n141 B.n140 10.6151
R1279 B.n144 B.n141 10.6151
R1280 B.n145 B.n144 10.6151
R1281 B.n148 B.n145 10.6151
R1282 B.n149 B.n148 10.6151
R1283 B.n152 B.n149 10.6151
R1284 B.n153 B.n152 10.6151
R1285 B.n156 B.n153 10.6151
R1286 B.n157 B.n156 10.6151
R1287 B.n160 B.n157 10.6151
R1288 B.n161 B.n160 10.6151
R1289 B.n164 B.n161 10.6151
R1290 B.n165 B.n164 10.6151
R1291 B.n168 B.n165 10.6151
R1292 B.n169 B.n168 10.6151
R1293 B.n172 B.n169 10.6151
R1294 B.n173 B.n172 10.6151
R1295 B.n176 B.n173 10.6151
R1296 B.n181 B.n178 10.6151
R1297 B.n182 B.n181 10.6151
R1298 B.n185 B.n182 10.6151
R1299 B.n186 B.n185 10.6151
R1300 B.n189 B.n186 10.6151
R1301 B.n190 B.n189 10.6151
R1302 B.n193 B.n190 10.6151
R1303 B.n194 B.n193 10.6151
R1304 B.n197 B.n194 10.6151
R1305 B.n202 B.n199 10.6151
R1306 B.n203 B.n202 10.6151
R1307 B.n206 B.n203 10.6151
R1308 B.n207 B.n206 10.6151
R1309 B.n210 B.n207 10.6151
R1310 B.n211 B.n210 10.6151
R1311 B.n214 B.n211 10.6151
R1312 B.n215 B.n214 10.6151
R1313 B.n218 B.n215 10.6151
R1314 B.n219 B.n218 10.6151
R1315 B.n222 B.n219 10.6151
R1316 B.n223 B.n222 10.6151
R1317 B.n226 B.n223 10.6151
R1318 B.n227 B.n226 10.6151
R1319 B.n230 B.n227 10.6151
R1320 B.n231 B.n230 10.6151
R1321 B.n234 B.n231 10.6151
R1322 B.n235 B.n234 10.6151
R1323 B.n238 B.n235 10.6151
R1324 B.n239 B.n238 10.6151
R1325 B.n242 B.n239 10.6151
R1326 B.n243 B.n242 10.6151
R1327 B.n246 B.n243 10.6151
R1328 B.n247 B.n246 10.6151
R1329 B.n250 B.n247 10.6151
R1330 B.n251 B.n250 10.6151
R1331 B.n254 B.n251 10.6151
R1332 B.n256 B.n254 10.6151
R1333 B.n257 B.n256 10.6151
R1334 B.n694 B.n257 10.6151
R1335 B.n438 B.n437 9.36635
R1336 B.n461 B.n355 9.36635
R1337 B.n177 B.n176 9.36635
R1338 B.n199 B.n198 9.36635
R1339 B.n782 B.n0 8.11757
R1340 B.n782 B.n1 8.11757
R1341 B.t1 B.n264 7.9744
R1342 B.n769 B.t2 7.9744
R1343 B.n439 B.n438 1.24928
R1344 B.n356 B.n355 1.24928
R1345 B.n178 B.n177 1.24928
R1346 B.n198 B.n197 1.24928
R1347 VP.n11 VP.n8 161.3
R1348 VP.n13 VP.n12 161.3
R1349 VP.n14 VP.n7 161.3
R1350 VP.n16 VP.n15 161.3
R1351 VP.n17 VP.n6 161.3
R1352 VP.n37 VP.n0 161.3
R1353 VP.n36 VP.n35 161.3
R1354 VP.n34 VP.n1 161.3
R1355 VP.n33 VP.n32 161.3
R1356 VP.n31 VP.n2 161.3
R1357 VP.n30 VP.n29 161.3
R1358 VP.n28 VP.n3 161.3
R1359 VP.n27 VP.n26 161.3
R1360 VP.n25 VP.n4 161.3
R1361 VP.n24 VP.n23 161.3
R1362 VP.n22 VP.n5 161.3
R1363 VP.n9 VP.t0 119.316
R1364 VP.n21 VP.n20 98.6123
R1365 VP.n39 VP.n38 98.6123
R1366 VP.n19 VP.n18 98.6123
R1367 VP.n30 VP.t4 84.8484
R1368 VP.n20 VP.t1 84.8484
R1369 VP.n38 VP.t3 84.8484
R1370 VP.n10 VP.t2 84.8484
R1371 VP.n18 VP.t5 84.8484
R1372 VP.n26 VP.n25 52.6866
R1373 VP.n32 VP.n1 52.6866
R1374 VP.n12 VP.n7 52.6866
R1375 VP.n10 VP.n9 48.1102
R1376 VP.n21 VP.n19 45.3443
R1377 VP.n25 VP.n24 28.4674
R1378 VP.n36 VP.n1 28.4674
R1379 VP.n16 VP.n7 28.4674
R1380 VP.n24 VP.n5 24.5923
R1381 VP.n26 VP.n3 24.5923
R1382 VP.n30 VP.n3 24.5923
R1383 VP.n31 VP.n30 24.5923
R1384 VP.n32 VP.n31 24.5923
R1385 VP.n37 VP.n36 24.5923
R1386 VP.n17 VP.n16 24.5923
R1387 VP.n11 VP.n10 24.5923
R1388 VP.n12 VP.n11 24.5923
R1389 VP.n20 VP.n5 12.2964
R1390 VP.n38 VP.n37 12.2964
R1391 VP.n18 VP.n17 12.2964
R1392 VP.n9 VP.n8 6.67081
R1393 VP.n19 VP.n6 0.278335
R1394 VP.n22 VP.n21 0.278335
R1395 VP.n39 VP.n0 0.278335
R1396 VP.n13 VP.n8 0.189894
R1397 VP.n14 VP.n13 0.189894
R1398 VP.n15 VP.n14 0.189894
R1399 VP.n15 VP.n6 0.189894
R1400 VP.n23 VP.n22 0.189894
R1401 VP.n23 VP.n4 0.189894
R1402 VP.n27 VP.n4 0.189894
R1403 VP.n28 VP.n27 0.189894
R1404 VP.n29 VP.n28 0.189894
R1405 VP.n29 VP.n2 0.189894
R1406 VP.n33 VP.n2 0.189894
R1407 VP.n34 VP.n33 0.189894
R1408 VP.n35 VP.n34 0.189894
R1409 VP.n35 VP.n0 0.189894
R1410 VP VP.n39 0.153485
R1411 VTAIL.n186 VTAIL.n146 289.615
R1412 VTAIL.n42 VTAIL.n2 289.615
R1413 VTAIL.n140 VTAIL.n100 289.615
R1414 VTAIL.n92 VTAIL.n52 289.615
R1415 VTAIL.n161 VTAIL.n160 185
R1416 VTAIL.n158 VTAIL.n157 185
R1417 VTAIL.n167 VTAIL.n166 185
R1418 VTAIL.n169 VTAIL.n168 185
R1419 VTAIL.n154 VTAIL.n153 185
R1420 VTAIL.n175 VTAIL.n174 185
R1421 VTAIL.n178 VTAIL.n177 185
R1422 VTAIL.n176 VTAIL.n150 185
R1423 VTAIL.n183 VTAIL.n149 185
R1424 VTAIL.n185 VTAIL.n184 185
R1425 VTAIL.n187 VTAIL.n186 185
R1426 VTAIL.n17 VTAIL.n16 185
R1427 VTAIL.n14 VTAIL.n13 185
R1428 VTAIL.n23 VTAIL.n22 185
R1429 VTAIL.n25 VTAIL.n24 185
R1430 VTAIL.n10 VTAIL.n9 185
R1431 VTAIL.n31 VTAIL.n30 185
R1432 VTAIL.n34 VTAIL.n33 185
R1433 VTAIL.n32 VTAIL.n6 185
R1434 VTAIL.n39 VTAIL.n5 185
R1435 VTAIL.n41 VTAIL.n40 185
R1436 VTAIL.n43 VTAIL.n42 185
R1437 VTAIL.n141 VTAIL.n140 185
R1438 VTAIL.n139 VTAIL.n138 185
R1439 VTAIL.n137 VTAIL.n103 185
R1440 VTAIL.n107 VTAIL.n104 185
R1441 VTAIL.n132 VTAIL.n131 185
R1442 VTAIL.n130 VTAIL.n129 185
R1443 VTAIL.n109 VTAIL.n108 185
R1444 VTAIL.n124 VTAIL.n123 185
R1445 VTAIL.n122 VTAIL.n121 185
R1446 VTAIL.n113 VTAIL.n112 185
R1447 VTAIL.n116 VTAIL.n115 185
R1448 VTAIL.n93 VTAIL.n92 185
R1449 VTAIL.n91 VTAIL.n90 185
R1450 VTAIL.n89 VTAIL.n55 185
R1451 VTAIL.n59 VTAIL.n56 185
R1452 VTAIL.n84 VTAIL.n83 185
R1453 VTAIL.n82 VTAIL.n81 185
R1454 VTAIL.n61 VTAIL.n60 185
R1455 VTAIL.n76 VTAIL.n75 185
R1456 VTAIL.n74 VTAIL.n73 185
R1457 VTAIL.n65 VTAIL.n64 185
R1458 VTAIL.n68 VTAIL.n67 185
R1459 VTAIL.t1 VTAIL.n159 149.524
R1460 VTAIL.t10 VTAIL.n15 149.524
R1461 VTAIL.t6 VTAIL.n114 149.524
R1462 VTAIL.t3 VTAIL.n66 149.524
R1463 VTAIL.n160 VTAIL.n157 104.615
R1464 VTAIL.n167 VTAIL.n157 104.615
R1465 VTAIL.n168 VTAIL.n167 104.615
R1466 VTAIL.n168 VTAIL.n153 104.615
R1467 VTAIL.n175 VTAIL.n153 104.615
R1468 VTAIL.n177 VTAIL.n175 104.615
R1469 VTAIL.n177 VTAIL.n176 104.615
R1470 VTAIL.n176 VTAIL.n149 104.615
R1471 VTAIL.n185 VTAIL.n149 104.615
R1472 VTAIL.n186 VTAIL.n185 104.615
R1473 VTAIL.n16 VTAIL.n13 104.615
R1474 VTAIL.n23 VTAIL.n13 104.615
R1475 VTAIL.n24 VTAIL.n23 104.615
R1476 VTAIL.n24 VTAIL.n9 104.615
R1477 VTAIL.n31 VTAIL.n9 104.615
R1478 VTAIL.n33 VTAIL.n31 104.615
R1479 VTAIL.n33 VTAIL.n32 104.615
R1480 VTAIL.n32 VTAIL.n5 104.615
R1481 VTAIL.n41 VTAIL.n5 104.615
R1482 VTAIL.n42 VTAIL.n41 104.615
R1483 VTAIL.n140 VTAIL.n139 104.615
R1484 VTAIL.n139 VTAIL.n103 104.615
R1485 VTAIL.n107 VTAIL.n103 104.615
R1486 VTAIL.n131 VTAIL.n107 104.615
R1487 VTAIL.n131 VTAIL.n130 104.615
R1488 VTAIL.n130 VTAIL.n108 104.615
R1489 VTAIL.n123 VTAIL.n108 104.615
R1490 VTAIL.n123 VTAIL.n122 104.615
R1491 VTAIL.n122 VTAIL.n112 104.615
R1492 VTAIL.n115 VTAIL.n112 104.615
R1493 VTAIL.n92 VTAIL.n91 104.615
R1494 VTAIL.n91 VTAIL.n55 104.615
R1495 VTAIL.n59 VTAIL.n55 104.615
R1496 VTAIL.n83 VTAIL.n59 104.615
R1497 VTAIL.n83 VTAIL.n82 104.615
R1498 VTAIL.n82 VTAIL.n60 104.615
R1499 VTAIL.n75 VTAIL.n60 104.615
R1500 VTAIL.n75 VTAIL.n74 104.615
R1501 VTAIL.n74 VTAIL.n64 104.615
R1502 VTAIL.n67 VTAIL.n64 104.615
R1503 VTAIL.n160 VTAIL.t1 52.3082
R1504 VTAIL.n16 VTAIL.t10 52.3082
R1505 VTAIL.n115 VTAIL.t6 52.3082
R1506 VTAIL.n67 VTAIL.t3 52.3082
R1507 VTAIL.n99 VTAIL.n98 46.7624
R1508 VTAIL.n51 VTAIL.n50 46.7624
R1509 VTAIL.n1 VTAIL.n0 46.7622
R1510 VTAIL.n49 VTAIL.n48 46.7622
R1511 VTAIL.n191 VTAIL.n190 32.1853
R1512 VTAIL.n47 VTAIL.n46 32.1853
R1513 VTAIL.n145 VTAIL.n144 32.1853
R1514 VTAIL.n97 VTAIL.n96 32.1853
R1515 VTAIL.n51 VTAIL.n49 24.4531
R1516 VTAIL.n191 VTAIL.n145 22.0824
R1517 VTAIL.n184 VTAIL.n183 13.1884
R1518 VTAIL.n40 VTAIL.n39 13.1884
R1519 VTAIL.n138 VTAIL.n137 13.1884
R1520 VTAIL.n90 VTAIL.n89 13.1884
R1521 VTAIL.n182 VTAIL.n150 12.8005
R1522 VTAIL.n187 VTAIL.n148 12.8005
R1523 VTAIL.n38 VTAIL.n6 12.8005
R1524 VTAIL.n43 VTAIL.n4 12.8005
R1525 VTAIL.n141 VTAIL.n102 12.8005
R1526 VTAIL.n136 VTAIL.n104 12.8005
R1527 VTAIL.n93 VTAIL.n54 12.8005
R1528 VTAIL.n88 VTAIL.n56 12.8005
R1529 VTAIL.n179 VTAIL.n178 12.0247
R1530 VTAIL.n188 VTAIL.n146 12.0247
R1531 VTAIL.n35 VTAIL.n34 12.0247
R1532 VTAIL.n44 VTAIL.n2 12.0247
R1533 VTAIL.n142 VTAIL.n100 12.0247
R1534 VTAIL.n133 VTAIL.n132 12.0247
R1535 VTAIL.n94 VTAIL.n52 12.0247
R1536 VTAIL.n85 VTAIL.n84 12.0247
R1537 VTAIL.n174 VTAIL.n152 11.249
R1538 VTAIL.n30 VTAIL.n8 11.249
R1539 VTAIL.n129 VTAIL.n106 11.249
R1540 VTAIL.n81 VTAIL.n58 11.249
R1541 VTAIL.n173 VTAIL.n154 10.4732
R1542 VTAIL.n29 VTAIL.n10 10.4732
R1543 VTAIL.n128 VTAIL.n109 10.4732
R1544 VTAIL.n80 VTAIL.n61 10.4732
R1545 VTAIL.n161 VTAIL.n159 10.2747
R1546 VTAIL.n17 VTAIL.n15 10.2747
R1547 VTAIL.n116 VTAIL.n114 10.2747
R1548 VTAIL.n68 VTAIL.n66 10.2747
R1549 VTAIL.n170 VTAIL.n169 9.69747
R1550 VTAIL.n26 VTAIL.n25 9.69747
R1551 VTAIL.n125 VTAIL.n124 9.69747
R1552 VTAIL.n77 VTAIL.n76 9.69747
R1553 VTAIL.n190 VTAIL.n189 9.45567
R1554 VTAIL.n46 VTAIL.n45 9.45567
R1555 VTAIL.n144 VTAIL.n143 9.45567
R1556 VTAIL.n96 VTAIL.n95 9.45567
R1557 VTAIL.n189 VTAIL.n188 9.3005
R1558 VTAIL.n148 VTAIL.n147 9.3005
R1559 VTAIL.n163 VTAIL.n162 9.3005
R1560 VTAIL.n165 VTAIL.n164 9.3005
R1561 VTAIL.n156 VTAIL.n155 9.3005
R1562 VTAIL.n171 VTAIL.n170 9.3005
R1563 VTAIL.n173 VTAIL.n172 9.3005
R1564 VTAIL.n152 VTAIL.n151 9.3005
R1565 VTAIL.n180 VTAIL.n179 9.3005
R1566 VTAIL.n182 VTAIL.n181 9.3005
R1567 VTAIL.n45 VTAIL.n44 9.3005
R1568 VTAIL.n4 VTAIL.n3 9.3005
R1569 VTAIL.n19 VTAIL.n18 9.3005
R1570 VTAIL.n21 VTAIL.n20 9.3005
R1571 VTAIL.n12 VTAIL.n11 9.3005
R1572 VTAIL.n27 VTAIL.n26 9.3005
R1573 VTAIL.n29 VTAIL.n28 9.3005
R1574 VTAIL.n8 VTAIL.n7 9.3005
R1575 VTAIL.n36 VTAIL.n35 9.3005
R1576 VTAIL.n38 VTAIL.n37 9.3005
R1577 VTAIL.n118 VTAIL.n117 9.3005
R1578 VTAIL.n120 VTAIL.n119 9.3005
R1579 VTAIL.n111 VTAIL.n110 9.3005
R1580 VTAIL.n126 VTAIL.n125 9.3005
R1581 VTAIL.n128 VTAIL.n127 9.3005
R1582 VTAIL.n106 VTAIL.n105 9.3005
R1583 VTAIL.n134 VTAIL.n133 9.3005
R1584 VTAIL.n136 VTAIL.n135 9.3005
R1585 VTAIL.n143 VTAIL.n142 9.3005
R1586 VTAIL.n102 VTAIL.n101 9.3005
R1587 VTAIL.n70 VTAIL.n69 9.3005
R1588 VTAIL.n72 VTAIL.n71 9.3005
R1589 VTAIL.n63 VTAIL.n62 9.3005
R1590 VTAIL.n78 VTAIL.n77 9.3005
R1591 VTAIL.n80 VTAIL.n79 9.3005
R1592 VTAIL.n58 VTAIL.n57 9.3005
R1593 VTAIL.n86 VTAIL.n85 9.3005
R1594 VTAIL.n88 VTAIL.n87 9.3005
R1595 VTAIL.n95 VTAIL.n94 9.3005
R1596 VTAIL.n54 VTAIL.n53 9.3005
R1597 VTAIL.n166 VTAIL.n156 8.92171
R1598 VTAIL.n22 VTAIL.n12 8.92171
R1599 VTAIL.n121 VTAIL.n111 8.92171
R1600 VTAIL.n73 VTAIL.n63 8.92171
R1601 VTAIL.n165 VTAIL.n158 8.14595
R1602 VTAIL.n21 VTAIL.n14 8.14595
R1603 VTAIL.n120 VTAIL.n113 8.14595
R1604 VTAIL.n72 VTAIL.n65 8.14595
R1605 VTAIL.n162 VTAIL.n161 7.3702
R1606 VTAIL.n18 VTAIL.n17 7.3702
R1607 VTAIL.n117 VTAIL.n116 7.3702
R1608 VTAIL.n69 VTAIL.n68 7.3702
R1609 VTAIL.n162 VTAIL.n158 5.81868
R1610 VTAIL.n18 VTAIL.n14 5.81868
R1611 VTAIL.n117 VTAIL.n113 5.81868
R1612 VTAIL.n69 VTAIL.n65 5.81868
R1613 VTAIL.n166 VTAIL.n165 5.04292
R1614 VTAIL.n22 VTAIL.n21 5.04292
R1615 VTAIL.n121 VTAIL.n120 5.04292
R1616 VTAIL.n73 VTAIL.n72 5.04292
R1617 VTAIL.n169 VTAIL.n156 4.26717
R1618 VTAIL.n25 VTAIL.n12 4.26717
R1619 VTAIL.n124 VTAIL.n111 4.26717
R1620 VTAIL.n76 VTAIL.n63 4.26717
R1621 VTAIL.n170 VTAIL.n154 3.49141
R1622 VTAIL.n26 VTAIL.n10 3.49141
R1623 VTAIL.n125 VTAIL.n109 3.49141
R1624 VTAIL.n77 VTAIL.n61 3.49141
R1625 VTAIL.n163 VTAIL.n159 2.84303
R1626 VTAIL.n19 VTAIL.n15 2.84303
R1627 VTAIL.n118 VTAIL.n114 2.84303
R1628 VTAIL.n70 VTAIL.n66 2.84303
R1629 VTAIL.n174 VTAIL.n173 2.71565
R1630 VTAIL.n30 VTAIL.n29 2.71565
R1631 VTAIL.n129 VTAIL.n128 2.71565
R1632 VTAIL.n81 VTAIL.n80 2.71565
R1633 VTAIL.n97 VTAIL.n51 2.37119
R1634 VTAIL.n145 VTAIL.n99 2.37119
R1635 VTAIL.n49 VTAIL.n47 2.37119
R1636 VTAIL.n0 VTAIL.t11 2.32444
R1637 VTAIL.n0 VTAIL.t0 2.32444
R1638 VTAIL.n48 VTAIL.t8 2.32444
R1639 VTAIL.n48 VTAIL.t7 2.32444
R1640 VTAIL.n98 VTAIL.t9 2.32444
R1641 VTAIL.n98 VTAIL.t5 2.32444
R1642 VTAIL.n50 VTAIL.t4 2.32444
R1643 VTAIL.n50 VTAIL.t2 2.32444
R1644 VTAIL.n178 VTAIL.n152 1.93989
R1645 VTAIL.n190 VTAIL.n146 1.93989
R1646 VTAIL.n34 VTAIL.n8 1.93989
R1647 VTAIL.n46 VTAIL.n2 1.93989
R1648 VTAIL.n144 VTAIL.n100 1.93989
R1649 VTAIL.n132 VTAIL.n106 1.93989
R1650 VTAIL.n96 VTAIL.n52 1.93989
R1651 VTAIL.n84 VTAIL.n58 1.93989
R1652 VTAIL VTAIL.n191 1.72033
R1653 VTAIL.n99 VTAIL.n97 1.65567
R1654 VTAIL.n47 VTAIL.n1 1.65567
R1655 VTAIL.n179 VTAIL.n150 1.16414
R1656 VTAIL.n188 VTAIL.n187 1.16414
R1657 VTAIL.n35 VTAIL.n6 1.16414
R1658 VTAIL.n44 VTAIL.n43 1.16414
R1659 VTAIL.n142 VTAIL.n141 1.16414
R1660 VTAIL.n133 VTAIL.n104 1.16414
R1661 VTAIL.n94 VTAIL.n93 1.16414
R1662 VTAIL.n85 VTAIL.n56 1.16414
R1663 VTAIL VTAIL.n1 0.651362
R1664 VTAIL.n183 VTAIL.n182 0.388379
R1665 VTAIL.n184 VTAIL.n148 0.388379
R1666 VTAIL.n39 VTAIL.n38 0.388379
R1667 VTAIL.n40 VTAIL.n4 0.388379
R1668 VTAIL.n138 VTAIL.n102 0.388379
R1669 VTAIL.n137 VTAIL.n136 0.388379
R1670 VTAIL.n90 VTAIL.n54 0.388379
R1671 VTAIL.n89 VTAIL.n88 0.388379
R1672 VTAIL.n164 VTAIL.n163 0.155672
R1673 VTAIL.n164 VTAIL.n155 0.155672
R1674 VTAIL.n171 VTAIL.n155 0.155672
R1675 VTAIL.n172 VTAIL.n171 0.155672
R1676 VTAIL.n172 VTAIL.n151 0.155672
R1677 VTAIL.n180 VTAIL.n151 0.155672
R1678 VTAIL.n181 VTAIL.n180 0.155672
R1679 VTAIL.n181 VTAIL.n147 0.155672
R1680 VTAIL.n189 VTAIL.n147 0.155672
R1681 VTAIL.n20 VTAIL.n19 0.155672
R1682 VTAIL.n20 VTAIL.n11 0.155672
R1683 VTAIL.n27 VTAIL.n11 0.155672
R1684 VTAIL.n28 VTAIL.n27 0.155672
R1685 VTAIL.n28 VTAIL.n7 0.155672
R1686 VTAIL.n36 VTAIL.n7 0.155672
R1687 VTAIL.n37 VTAIL.n36 0.155672
R1688 VTAIL.n37 VTAIL.n3 0.155672
R1689 VTAIL.n45 VTAIL.n3 0.155672
R1690 VTAIL.n143 VTAIL.n101 0.155672
R1691 VTAIL.n135 VTAIL.n101 0.155672
R1692 VTAIL.n135 VTAIL.n134 0.155672
R1693 VTAIL.n134 VTAIL.n105 0.155672
R1694 VTAIL.n127 VTAIL.n105 0.155672
R1695 VTAIL.n127 VTAIL.n126 0.155672
R1696 VTAIL.n126 VTAIL.n110 0.155672
R1697 VTAIL.n119 VTAIL.n110 0.155672
R1698 VTAIL.n119 VTAIL.n118 0.155672
R1699 VTAIL.n95 VTAIL.n53 0.155672
R1700 VTAIL.n87 VTAIL.n53 0.155672
R1701 VTAIL.n87 VTAIL.n86 0.155672
R1702 VTAIL.n86 VTAIL.n57 0.155672
R1703 VTAIL.n79 VTAIL.n57 0.155672
R1704 VTAIL.n79 VTAIL.n78 0.155672
R1705 VTAIL.n78 VTAIL.n62 0.155672
R1706 VTAIL.n71 VTAIL.n62 0.155672
R1707 VTAIL.n71 VTAIL.n70 0.155672
R1708 VDD1.n40 VDD1.n0 289.615
R1709 VDD1.n85 VDD1.n45 289.615
R1710 VDD1.n41 VDD1.n40 185
R1711 VDD1.n39 VDD1.n38 185
R1712 VDD1.n37 VDD1.n3 185
R1713 VDD1.n7 VDD1.n4 185
R1714 VDD1.n32 VDD1.n31 185
R1715 VDD1.n30 VDD1.n29 185
R1716 VDD1.n9 VDD1.n8 185
R1717 VDD1.n24 VDD1.n23 185
R1718 VDD1.n22 VDD1.n21 185
R1719 VDD1.n13 VDD1.n12 185
R1720 VDD1.n16 VDD1.n15 185
R1721 VDD1.n60 VDD1.n59 185
R1722 VDD1.n57 VDD1.n56 185
R1723 VDD1.n66 VDD1.n65 185
R1724 VDD1.n68 VDD1.n67 185
R1725 VDD1.n53 VDD1.n52 185
R1726 VDD1.n74 VDD1.n73 185
R1727 VDD1.n77 VDD1.n76 185
R1728 VDD1.n75 VDD1.n49 185
R1729 VDD1.n82 VDD1.n48 185
R1730 VDD1.n84 VDD1.n83 185
R1731 VDD1.n86 VDD1.n85 185
R1732 VDD1.t5 VDD1.n14 149.524
R1733 VDD1.t4 VDD1.n58 149.524
R1734 VDD1.n40 VDD1.n39 104.615
R1735 VDD1.n39 VDD1.n3 104.615
R1736 VDD1.n7 VDD1.n3 104.615
R1737 VDD1.n31 VDD1.n7 104.615
R1738 VDD1.n31 VDD1.n30 104.615
R1739 VDD1.n30 VDD1.n8 104.615
R1740 VDD1.n23 VDD1.n8 104.615
R1741 VDD1.n23 VDD1.n22 104.615
R1742 VDD1.n22 VDD1.n12 104.615
R1743 VDD1.n15 VDD1.n12 104.615
R1744 VDD1.n59 VDD1.n56 104.615
R1745 VDD1.n66 VDD1.n56 104.615
R1746 VDD1.n67 VDD1.n66 104.615
R1747 VDD1.n67 VDD1.n52 104.615
R1748 VDD1.n74 VDD1.n52 104.615
R1749 VDD1.n76 VDD1.n74 104.615
R1750 VDD1.n76 VDD1.n75 104.615
R1751 VDD1.n75 VDD1.n48 104.615
R1752 VDD1.n84 VDD1.n48 104.615
R1753 VDD1.n85 VDD1.n84 104.615
R1754 VDD1.n91 VDD1.n90 63.9783
R1755 VDD1.n93 VDD1.n92 63.441
R1756 VDD1.n15 VDD1.t5 52.3082
R1757 VDD1.n59 VDD1.t4 52.3082
R1758 VDD1 VDD1.n44 50.7003
R1759 VDD1.n91 VDD1.n89 50.5868
R1760 VDD1.n93 VDD1.n91 40.5332
R1761 VDD1.n38 VDD1.n37 13.1884
R1762 VDD1.n83 VDD1.n82 13.1884
R1763 VDD1.n41 VDD1.n2 12.8005
R1764 VDD1.n36 VDD1.n4 12.8005
R1765 VDD1.n81 VDD1.n49 12.8005
R1766 VDD1.n86 VDD1.n47 12.8005
R1767 VDD1.n42 VDD1.n0 12.0247
R1768 VDD1.n33 VDD1.n32 12.0247
R1769 VDD1.n78 VDD1.n77 12.0247
R1770 VDD1.n87 VDD1.n45 12.0247
R1771 VDD1.n29 VDD1.n6 11.249
R1772 VDD1.n73 VDD1.n51 11.249
R1773 VDD1.n28 VDD1.n9 10.4732
R1774 VDD1.n72 VDD1.n53 10.4732
R1775 VDD1.n16 VDD1.n14 10.2747
R1776 VDD1.n60 VDD1.n58 10.2747
R1777 VDD1.n25 VDD1.n24 9.69747
R1778 VDD1.n69 VDD1.n68 9.69747
R1779 VDD1.n44 VDD1.n43 9.45567
R1780 VDD1.n89 VDD1.n88 9.45567
R1781 VDD1.n18 VDD1.n17 9.3005
R1782 VDD1.n20 VDD1.n19 9.3005
R1783 VDD1.n11 VDD1.n10 9.3005
R1784 VDD1.n26 VDD1.n25 9.3005
R1785 VDD1.n28 VDD1.n27 9.3005
R1786 VDD1.n6 VDD1.n5 9.3005
R1787 VDD1.n34 VDD1.n33 9.3005
R1788 VDD1.n36 VDD1.n35 9.3005
R1789 VDD1.n43 VDD1.n42 9.3005
R1790 VDD1.n2 VDD1.n1 9.3005
R1791 VDD1.n88 VDD1.n87 9.3005
R1792 VDD1.n47 VDD1.n46 9.3005
R1793 VDD1.n62 VDD1.n61 9.3005
R1794 VDD1.n64 VDD1.n63 9.3005
R1795 VDD1.n55 VDD1.n54 9.3005
R1796 VDD1.n70 VDD1.n69 9.3005
R1797 VDD1.n72 VDD1.n71 9.3005
R1798 VDD1.n51 VDD1.n50 9.3005
R1799 VDD1.n79 VDD1.n78 9.3005
R1800 VDD1.n81 VDD1.n80 9.3005
R1801 VDD1.n21 VDD1.n11 8.92171
R1802 VDD1.n65 VDD1.n55 8.92171
R1803 VDD1.n20 VDD1.n13 8.14595
R1804 VDD1.n64 VDD1.n57 8.14595
R1805 VDD1.n17 VDD1.n16 7.3702
R1806 VDD1.n61 VDD1.n60 7.3702
R1807 VDD1.n17 VDD1.n13 5.81868
R1808 VDD1.n61 VDD1.n57 5.81868
R1809 VDD1.n21 VDD1.n20 5.04292
R1810 VDD1.n65 VDD1.n64 5.04292
R1811 VDD1.n24 VDD1.n11 4.26717
R1812 VDD1.n68 VDD1.n55 4.26717
R1813 VDD1.n25 VDD1.n9 3.49141
R1814 VDD1.n69 VDD1.n53 3.49141
R1815 VDD1.n62 VDD1.n58 2.84303
R1816 VDD1.n18 VDD1.n14 2.84303
R1817 VDD1.n29 VDD1.n28 2.71565
R1818 VDD1.n73 VDD1.n72 2.71565
R1819 VDD1.n92 VDD1.t3 2.32444
R1820 VDD1.n92 VDD1.t0 2.32444
R1821 VDD1.n90 VDD1.t1 2.32444
R1822 VDD1.n90 VDD1.t2 2.32444
R1823 VDD1.n44 VDD1.n0 1.93989
R1824 VDD1.n32 VDD1.n6 1.93989
R1825 VDD1.n77 VDD1.n51 1.93989
R1826 VDD1.n89 VDD1.n45 1.93989
R1827 VDD1.n42 VDD1.n41 1.16414
R1828 VDD1.n33 VDD1.n4 1.16414
R1829 VDD1.n78 VDD1.n49 1.16414
R1830 VDD1.n87 VDD1.n86 1.16414
R1831 VDD1 VDD1.n93 0.534983
R1832 VDD1.n38 VDD1.n2 0.388379
R1833 VDD1.n37 VDD1.n36 0.388379
R1834 VDD1.n82 VDD1.n81 0.388379
R1835 VDD1.n83 VDD1.n47 0.388379
R1836 VDD1.n43 VDD1.n1 0.155672
R1837 VDD1.n35 VDD1.n1 0.155672
R1838 VDD1.n35 VDD1.n34 0.155672
R1839 VDD1.n34 VDD1.n5 0.155672
R1840 VDD1.n27 VDD1.n5 0.155672
R1841 VDD1.n27 VDD1.n26 0.155672
R1842 VDD1.n26 VDD1.n10 0.155672
R1843 VDD1.n19 VDD1.n10 0.155672
R1844 VDD1.n19 VDD1.n18 0.155672
R1845 VDD1.n63 VDD1.n62 0.155672
R1846 VDD1.n63 VDD1.n54 0.155672
R1847 VDD1.n70 VDD1.n54 0.155672
R1848 VDD1.n71 VDD1.n70 0.155672
R1849 VDD1.n71 VDD1.n50 0.155672
R1850 VDD1.n79 VDD1.n50 0.155672
R1851 VDD1.n80 VDD1.n79 0.155672
R1852 VDD1.n80 VDD1.n46 0.155672
R1853 VDD1.n88 VDD1.n46 0.155672
R1854 VN.n25 VN.n14 161.3
R1855 VN.n24 VN.n23 161.3
R1856 VN.n22 VN.n15 161.3
R1857 VN.n21 VN.n20 161.3
R1858 VN.n19 VN.n16 161.3
R1859 VN.n11 VN.n0 161.3
R1860 VN.n10 VN.n9 161.3
R1861 VN.n8 VN.n1 161.3
R1862 VN.n7 VN.n6 161.3
R1863 VN.n5 VN.n2 161.3
R1864 VN.n3 VN.t2 119.316
R1865 VN.n17 VN.t3 119.316
R1866 VN.n13 VN.n12 98.6123
R1867 VN.n27 VN.n26 98.6123
R1868 VN.n4 VN.t5 84.8484
R1869 VN.n12 VN.t1 84.8484
R1870 VN.n18 VN.t4 84.8484
R1871 VN.n26 VN.t0 84.8484
R1872 VN.n6 VN.n1 52.6866
R1873 VN.n20 VN.n15 52.6866
R1874 VN.n4 VN.n3 48.1102
R1875 VN.n18 VN.n17 48.1102
R1876 VN VN.n27 45.6232
R1877 VN.n10 VN.n1 28.4674
R1878 VN.n24 VN.n15 28.4674
R1879 VN.n5 VN.n4 24.5923
R1880 VN.n6 VN.n5 24.5923
R1881 VN.n11 VN.n10 24.5923
R1882 VN.n20 VN.n19 24.5923
R1883 VN.n19 VN.n18 24.5923
R1884 VN.n25 VN.n24 24.5923
R1885 VN.n12 VN.n11 12.2964
R1886 VN.n26 VN.n25 12.2964
R1887 VN.n17 VN.n16 6.67081
R1888 VN.n3 VN.n2 6.67081
R1889 VN.n27 VN.n14 0.278335
R1890 VN.n13 VN.n0 0.278335
R1891 VN.n23 VN.n14 0.189894
R1892 VN.n23 VN.n22 0.189894
R1893 VN.n22 VN.n21 0.189894
R1894 VN.n21 VN.n16 0.189894
R1895 VN.n7 VN.n2 0.189894
R1896 VN.n8 VN.n7 0.189894
R1897 VN.n9 VN.n8 0.189894
R1898 VN.n9 VN.n0 0.189894
R1899 VN VN.n13 0.153485
R1900 VDD2.n87 VDD2.n47 289.615
R1901 VDD2.n40 VDD2.n0 289.615
R1902 VDD2.n88 VDD2.n87 185
R1903 VDD2.n86 VDD2.n85 185
R1904 VDD2.n84 VDD2.n50 185
R1905 VDD2.n54 VDD2.n51 185
R1906 VDD2.n79 VDD2.n78 185
R1907 VDD2.n77 VDD2.n76 185
R1908 VDD2.n56 VDD2.n55 185
R1909 VDD2.n71 VDD2.n70 185
R1910 VDD2.n69 VDD2.n68 185
R1911 VDD2.n60 VDD2.n59 185
R1912 VDD2.n63 VDD2.n62 185
R1913 VDD2.n15 VDD2.n14 185
R1914 VDD2.n12 VDD2.n11 185
R1915 VDD2.n21 VDD2.n20 185
R1916 VDD2.n23 VDD2.n22 185
R1917 VDD2.n8 VDD2.n7 185
R1918 VDD2.n29 VDD2.n28 185
R1919 VDD2.n32 VDD2.n31 185
R1920 VDD2.n30 VDD2.n4 185
R1921 VDD2.n37 VDD2.n3 185
R1922 VDD2.n39 VDD2.n38 185
R1923 VDD2.n41 VDD2.n40 185
R1924 VDD2.t5 VDD2.n61 149.524
R1925 VDD2.t3 VDD2.n13 149.524
R1926 VDD2.n87 VDD2.n86 104.615
R1927 VDD2.n86 VDD2.n50 104.615
R1928 VDD2.n54 VDD2.n50 104.615
R1929 VDD2.n78 VDD2.n54 104.615
R1930 VDD2.n78 VDD2.n77 104.615
R1931 VDD2.n77 VDD2.n55 104.615
R1932 VDD2.n70 VDD2.n55 104.615
R1933 VDD2.n70 VDD2.n69 104.615
R1934 VDD2.n69 VDD2.n59 104.615
R1935 VDD2.n62 VDD2.n59 104.615
R1936 VDD2.n14 VDD2.n11 104.615
R1937 VDD2.n21 VDD2.n11 104.615
R1938 VDD2.n22 VDD2.n21 104.615
R1939 VDD2.n22 VDD2.n7 104.615
R1940 VDD2.n29 VDD2.n7 104.615
R1941 VDD2.n31 VDD2.n29 104.615
R1942 VDD2.n31 VDD2.n30 104.615
R1943 VDD2.n30 VDD2.n3 104.615
R1944 VDD2.n39 VDD2.n3 104.615
R1945 VDD2.n40 VDD2.n39 104.615
R1946 VDD2.n46 VDD2.n45 63.9783
R1947 VDD2 VDD2.n93 63.9755
R1948 VDD2.n62 VDD2.t5 52.3082
R1949 VDD2.n14 VDD2.t3 52.3082
R1950 VDD2.n46 VDD2.n44 50.5868
R1951 VDD2.n92 VDD2.n91 48.8641
R1952 VDD2.n92 VDD2.n46 38.7649
R1953 VDD2.n85 VDD2.n84 13.1884
R1954 VDD2.n38 VDD2.n37 13.1884
R1955 VDD2.n88 VDD2.n49 12.8005
R1956 VDD2.n83 VDD2.n51 12.8005
R1957 VDD2.n36 VDD2.n4 12.8005
R1958 VDD2.n41 VDD2.n2 12.8005
R1959 VDD2.n89 VDD2.n47 12.0247
R1960 VDD2.n80 VDD2.n79 12.0247
R1961 VDD2.n33 VDD2.n32 12.0247
R1962 VDD2.n42 VDD2.n0 12.0247
R1963 VDD2.n76 VDD2.n53 11.249
R1964 VDD2.n28 VDD2.n6 11.249
R1965 VDD2.n75 VDD2.n56 10.4732
R1966 VDD2.n27 VDD2.n8 10.4732
R1967 VDD2.n63 VDD2.n61 10.2747
R1968 VDD2.n15 VDD2.n13 10.2747
R1969 VDD2.n72 VDD2.n71 9.69747
R1970 VDD2.n24 VDD2.n23 9.69747
R1971 VDD2.n91 VDD2.n90 9.45567
R1972 VDD2.n44 VDD2.n43 9.45567
R1973 VDD2.n65 VDD2.n64 9.3005
R1974 VDD2.n67 VDD2.n66 9.3005
R1975 VDD2.n58 VDD2.n57 9.3005
R1976 VDD2.n73 VDD2.n72 9.3005
R1977 VDD2.n75 VDD2.n74 9.3005
R1978 VDD2.n53 VDD2.n52 9.3005
R1979 VDD2.n81 VDD2.n80 9.3005
R1980 VDD2.n83 VDD2.n82 9.3005
R1981 VDD2.n90 VDD2.n89 9.3005
R1982 VDD2.n49 VDD2.n48 9.3005
R1983 VDD2.n43 VDD2.n42 9.3005
R1984 VDD2.n2 VDD2.n1 9.3005
R1985 VDD2.n17 VDD2.n16 9.3005
R1986 VDD2.n19 VDD2.n18 9.3005
R1987 VDD2.n10 VDD2.n9 9.3005
R1988 VDD2.n25 VDD2.n24 9.3005
R1989 VDD2.n27 VDD2.n26 9.3005
R1990 VDD2.n6 VDD2.n5 9.3005
R1991 VDD2.n34 VDD2.n33 9.3005
R1992 VDD2.n36 VDD2.n35 9.3005
R1993 VDD2.n68 VDD2.n58 8.92171
R1994 VDD2.n20 VDD2.n10 8.92171
R1995 VDD2.n67 VDD2.n60 8.14595
R1996 VDD2.n19 VDD2.n12 8.14595
R1997 VDD2.n64 VDD2.n63 7.3702
R1998 VDD2.n16 VDD2.n15 7.3702
R1999 VDD2.n64 VDD2.n60 5.81868
R2000 VDD2.n16 VDD2.n12 5.81868
R2001 VDD2.n68 VDD2.n67 5.04292
R2002 VDD2.n20 VDD2.n19 5.04292
R2003 VDD2.n71 VDD2.n58 4.26717
R2004 VDD2.n23 VDD2.n10 4.26717
R2005 VDD2.n72 VDD2.n56 3.49141
R2006 VDD2.n24 VDD2.n8 3.49141
R2007 VDD2.n17 VDD2.n13 2.84303
R2008 VDD2.n65 VDD2.n61 2.84303
R2009 VDD2.n76 VDD2.n75 2.71565
R2010 VDD2.n28 VDD2.n27 2.71565
R2011 VDD2.n93 VDD2.t1 2.32444
R2012 VDD2.n93 VDD2.t2 2.32444
R2013 VDD2.n45 VDD2.t0 2.32444
R2014 VDD2.n45 VDD2.t4 2.32444
R2015 VDD2.n91 VDD2.n47 1.93989
R2016 VDD2.n79 VDD2.n53 1.93989
R2017 VDD2.n32 VDD2.n6 1.93989
R2018 VDD2.n44 VDD2.n0 1.93989
R2019 VDD2 VDD2.n92 1.83671
R2020 VDD2.n89 VDD2.n88 1.16414
R2021 VDD2.n80 VDD2.n51 1.16414
R2022 VDD2.n33 VDD2.n4 1.16414
R2023 VDD2.n42 VDD2.n41 1.16414
R2024 VDD2.n85 VDD2.n49 0.388379
R2025 VDD2.n84 VDD2.n83 0.388379
R2026 VDD2.n37 VDD2.n36 0.388379
R2027 VDD2.n38 VDD2.n2 0.388379
R2028 VDD2.n90 VDD2.n48 0.155672
R2029 VDD2.n82 VDD2.n48 0.155672
R2030 VDD2.n82 VDD2.n81 0.155672
R2031 VDD2.n81 VDD2.n52 0.155672
R2032 VDD2.n74 VDD2.n52 0.155672
R2033 VDD2.n74 VDD2.n73 0.155672
R2034 VDD2.n73 VDD2.n57 0.155672
R2035 VDD2.n66 VDD2.n57 0.155672
R2036 VDD2.n66 VDD2.n65 0.155672
R2037 VDD2.n18 VDD2.n17 0.155672
R2038 VDD2.n18 VDD2.n9 0.155672
R2039 VDD2.n25 VDD2.n9 0.155672
R2040 VDD2.n26 VDD2.n25 0.155672
R2041 VDD2.n26 VDD2.n5 0.155672
R2042 VDD2.n34 VDD2.n5 0.155672
R2043 VDD2.n35 VDD2.n34 0.155672
R2044 VDD2.n35 VDD2.n1 0.155672
R2045 VDD2.n43 VDD2.n1 0.155672
C0 VDD2 VN 4.81603f
C1 VDD1 VDD2 1.33646f
C2 VDD1 VN 0.150826f
C3 VTAIL VP 5.09829f
C4 VTAIL VDD2 6.4598f
C5 VTAIL VN 5.08405f
C6 VP VDD2 0.443107f
C7 VDD1 VTAIL 6.40951f
C8 VP VN 6.10274f
C9 VDD1 VP 5.10572f
C10 VDD2 B 5.231028f
C11 VDD1 B 5.349606f
C12 VTAIL B 6.312391f
C13 VN B 12.07618f
C14 VP B 10.729935f
C15 VDD2.n0 B 0.027518f
C16 VDD2.n1 B 0.021656f
C17 VDD2.n2 B 0.011637f
C18 VDD2.n3 B 0.027506f
C19 VDD2.n4 B 0.012322f
C20 VDD2.n5 B 0.021656f
C21 VDD2.n6 B 0.011637f
C22 VDD2.n7 B 0.027506f
C23 VDD2.n8 B 0.012322f
C24 VDD2.n9 B 0.021656f
C25 VDD2.n10 B 0.011637f
C26 VDD2.n11 B 0.027506f
C27 VDD2.n12 B 0.012322f
C28 VDD2.n13 B 0.127216f
C29 VDD2.t3 B 0.046056f
C30 VDD2.n14 B 0.02063f
C31 VDD2.n15 B 0.019445f
C32 VDD2.n16 B 0.011637f
C33 VDD2.n17 B 0.757304f
C34 VDD2.n18 B 0.021656f
C35 VDD2.n19 B 0.011637f
C36 VDD2.n20 B 0.012322f
C37 VDD2.n21 B 0.027506f
C38 VDD2.n22 B 0.027506f
C39 VDD2.n23 B 0.012322f
C40 VDD2.n24 B 0.011637f
C41 VDD2.n25 B 0.021656f
C42 VDD2.n26 B 0.021656f
C43 VDD2.n27 B 0.011637f
C44 VDD2.n28 B 0.012322f
C45 VDD2.n29 B 0.027506f
C46 VDD2.n30 B 0.027506f
C47 VDD2.n31 B 0.027506f
C48 VDD2.n32 B 0.012322f
C49 VDD2.n33 B 0.011637f
C50 VDD2.n34 B 0.021656f
C51 VDD2.n35 B 0.021656f
C52 VDD2.n36 B 0.011637f
C53 VDD2.n37 B 0.011979f
C54 VDD2.n38 B 0.011979f
C55 VDD2.n39 B 0.027506f
C56 VDD2.n40 B 0.054378f
C57 VDD2.n41 B 0.012322f
C58 VDD2.n42 B 0.011637f
C59 VDD2.n43 B 0.050058f
C60 VDD2.n44 B 0.050373f
C61 VDD2.t0 B 0.145808f
C62 VDD2.t4 B 0.145808f
C63 VDD2.n45 B 1.27167f
C64 VDD2.n46 B 2.06453f
C65 VDD2.n47 B 0.027518f
C66 VDD2.n48 B 0.021656f
C67 VDD2.n49 B 0.011637f
C68 VDD2.n50 B 0.027506f
C69 VDD2.n51 B 0.012322f
C70 VDD2.n52 B 0.021656f
C71 VDD2.n53 B 0.011637f
C72 VDD2.n54 B 0.027506f
C73 VDD2.n55 B 0.027506f
C74 VDD2.n56 B 0.012322f
C75 VDD2.n57 B 0.021656f
C76 VDD2.n58 B 0.011637f
C77 VDD2.n59 B 0.027506f
C78 VDD2.n60 B 0.012322f
C79 VDD2.n61 B 0.127216f
C80 VDD2.t5 B 0.046056f
C81 VDD2.n62 B 0.02063f
C82 VDD2.n63 B 0.019445f
C83 VDD2.n64 B 0.011637f
C84 VDD2.n65 B 0.757304f
C85 VDD2.n66 B 0.021656f
C86 VDD2.n67 B 0.011637f
C87 VDD2.n68 B 0.012322f
C88 VDD2.n69 B 0.027506f
C89 VDD2.n70 B 0.027506f
C90 VDD2.n71 B 0.012322f
C91 VDD2.n72 B 0.011637f
C92 VDD2.n73 B 0.021656f
C93 VDD2.n74 B 0.021656f
C94 VDD2.n75 B 0.011637f
C95 VDD2.n76 B 0.012322f
C96 VDD2.n77 B 0.027506f
C97 VDD2.n78 B 0.027506f
C98 VDD2.n79 B 0.012322f
C99 VDD2.n80 B 0.011637f
C100 VDD2.n81 B 0.021656f
C101 VDD2.n82 B 0.021656f
C102 VDD2.n83 B 0.011637f
C103 VDD2.n84 B 0.011979f
C104 VDD2.n85 B 0.011979f
C105 VDD2.n86 B 0.027506f
C106 VDD2.n87 B 0.054378f
C107 VDD2.n88 B 0.012322f
C108 VDD2.n89 B 0.011637f
C109 VDD2.n90 B 0.050058f
C110 VDD2.n91 B 0.044849f
C111 VDD2.n92 B 1.94135f
C112 VDD2.t1 B 0.145808f
C113 VDD2.t2 B 0.145808f
C114 VDD2.n93 B 1.27164f
C115 VN.n0 B 0.033601f
C116 VN.t1 B 1.41512f
C117 VN.n1 B 0.026159f
C118 VN.n2 B 0.241708f
C119 VN.t5 B 1.41512f
C120 VN.t2 B 1.60733f
C121 VN.n3 B 0.563155f
C122 VN.n4 B 0.598027f
C123 VN.n5 B 0.047264f
C124 VN.n6 B 0.045274f
C125 VN.n7 B 0.025488f
C126 VN.n8 B 0.025488f
C127 VN.n9 B 0.025488f
C128 VN.n10 B 0.049933f
C129 VN.n11 B 0.035598f
C130 VN.n12 B 0.59619f
C131 VN.n13 B 0.038606f
C132 VN.n14 B 0.033601f
C133 VN.t0 B 1.41512f
C134 VN.n15 B 0.026159f
C135 VN.n16 B 0.241708f
C136 VN.t4 B 1.41512f
C137 VN.t3 B 1.60733f
C138 VN.n17 B 0.563155f
C139 VN.n18 B 0.598027f
C140 VN.n19 B 0.047264f
C141 VN.n20 B 0.045274f
C142 VN.n21 B 0.025488f
C143 VN.n22 B 0.025488f
C144 VN.n23 B 0.025488f
C145 VN.n24 B 0.049933f
C146 VN.n25 B 0.035598f
C147 VN.n26 B 0.59619f
C148 VN.n27 B 1.23493f
C149 VDD1.n0 B 0.027808f
C150 VDD1.n1 B 0.021885f
C151 VDD1.n2 B 0.01176f
C152 VDD1.n3 B 0.027796f
C153 VDD1.n4 B 0.012452f
C154 VDD1.n5 B 0.021885f
C155 VDD1.n6 B 0.01176f
C156 VDD1.n7 B 0.027796f
C157 VDD1.n8 B 0.027796f
C158 VDD1.n9 B 0.012452f
C159 VDD1.n10 B 0.021885f
C160 VDD1.n11 B 0.01176f
C161 VDD1.n12 B 0.027796f
C162 VDD1.n13 B 0.012452f
C163 VDD1.n14 B 0.128558f
C164 VDD1.t5 B 0.046541f
C165 VDD1.n15 B 0.020847f
C166 VDD1.n16 B 0.01965f
C167 VDD1.n17 B 0.01176f
C168 VDD1.n18 B 0.76529f
C169 VDD1.n19 B 0.021885f
C170 VDD1.n20 B 0.01176f
C171 VDD1.n21 B 0.012452f
C172 VDD1.n22 B 0.027796f
C173 VDD1.n23 B 0.027796f
C174 VDD1.n24 B 0.012452f
C175 VDD1.n25 B 0.01176f
C176 VDD1.n26 B 0.021885f
C177 VDD1.n27 B 0.021885f
C178 VDD1.n28 B 0.01176f
C179 VDD1.n29 B 0.012452f
C180 VDD1.n30 B 0.027796f
C181 VDD1.n31 B 0.027796f
C182 VDD1.n32 B 0.012452f
C183 VDD1.n33 B 0.01176f
C184 VDD1.n34 B 0.021885f
C185 VDD1.n35 B 0.021885f
C186 VDD1.n36 B 0.01176f
C187 VDD1.n37 B 0.012106f
C188 VDD1.n38 B 0.012106f
C189 VDD1.n39 B 0.027796f
C190 VDD1.n40 B 0.054952f
C191 VDD1.n41 B 0.012452f
C192 VDD1.n42 B 0.01176f
C193 VDD1.n43 B 0.050586f
C194 VDD1.n44 B 0.051538f
C195 VDD1.n45 B 0.027808f
C196 VDD1.n46 B 0.021885f
C197 VDD1.n47 B 0.01176f
C198 VDD1.n48 B 0.027796f
C199 VDD1.n49 B 0.012452f
C200 VDD1.n50 B 0.021885f
C201 VDD1.n51 B 0.01176f
C202 VDD1.n52 B 0.027796f
C203 VDD1.n53 B 0.012452f
C204 VDD1.n54 B 0.021885f
C205 VDD1.n55 B 0.01176f
C206 VDD1.n56 B 0.027796f
C207 VDD1.n57 B 0.012452f
C208 VDD1.n58 B 0.128558f
C209 VDD1.t4 B 0.046541f
C210 VDD1.n59 B 0.020847f
C211 VDD1.n60 B 0.01965f
C212 VDD1.n61 B 0.01176f
C213 VDD1.n62 B 0.76529f
C214 VDD1.n63 B 0.021885f
C215 VDD1.n64 B 0.01176f
C216 VDD1.n65 B 0.012452f
C217 VDD1.n66 B 0.027796f
C218 VDD1.n67 B 0.027796f
C219 VDD1.n68 B 0.012452f
C220 VDD1.n69 B 0.01176f
C221 VDD1.n70 B 0.021885f
C222 VDD1.n71 B 0.021885f
C223 VDD1.n72 B 0.01176f
C224 VDD1.n73 B 0.012452f
C225 VDD1.n74 B 0.027796f
C226 VDD1.n75 B 0.027796f
C227 VDD1.n76 B 0.027796f
C228 VDD1.n77 B 0.012452f
C229 VDD1.n78 B 0.01176f
C230 VDD1.n79 B 0.021885f
C231 VDD1.n80 B 0.021885f
C232 VDD1.n81 B 0.01176f
C233 VDD1.n82 B 0.012106f
C234 VDD1.n83 B 0.012106f
C235 VDD1.n84 B 0.027796f
C236 VDD1.n85 B 0.054952f
C237 VDD1.n86 B 0.012452f
C238 VDD1.n87 B 0.01176f
C239 VDD1.n88 B 0.050586f
C240 VDD1.n89 B 0.050904f
C241 VDD1.t1 B 0.147345f
C242 VDD1.t2 B 0.147345f
C243 VDD1.n90 B 1.28508f
C244 VDD1.n91 B 2.18836f
C245 VDD1.t3 B 0.147345f
C246 VDD1.t0 B 0.147345f
C247 VDD1.n92 B 1.2818f
C248 VDD1.n93 B 2.15856f
C249 VTAIL.t11 B 0.167851f
C250 VTAIL.t0 B 0.167851f
C251 VTAIL.n0 B 1.3904f
C252 VTAIL.n1 B 0.421521f
C253 VTAIL.n2 B 0.031678f
C254 VTAIL.n3 B 0.02493f
C255 VTAIL.n4 B 0.013396f
C256 VTAIL.n5 B 0.031665f
C257 VTAIL.n6 B 0.014185f
C258 VTAIL.n7 B 0.02493f
C259 VTAIL.n8 B 0.013396f
C260 VTAIL.n9 B 0.031665f
C261 VTAIL.n10 B 0.014185f
C262 VTAIL.n11 B 0.02493f
C263 VTAIL.n12 B 0.013396f
C264 VTAIL.n13 B 0.031665f
C265 VTAIL.n14 B 0.014185f
C266 VTAIL.n15 B 0.146449f
C267 VTAIL.t10 B 0.053018f
C268 VTAIL.n16 B 0.023748f
C269 VTAIL.n17 B 0.022384f
C270 VTAIL.n18 B 0.013396f
C271 VTAIL.n19 B 0.871792f
C272 VTAIL.n20 B 0.02493f
C273 VTAIL.n21 B 0.013396f
C274 VTAIL.n22 B 0.014185f
C275 VTAIL.n23 B 0.031665f
C276 VTAIL.n24 B 0.031665f
C277 VTAIL.n25 B 0.014185f
C278 VTAIL.n26 B 0.013396f
C279 VTAIL.n27 B 0.02493f
C280 VTAIL.n28 B 0.02493f
C281 VTAIL.n29 B 0.013396f
C282 VTAIL.n30 B 0.014185f
C283 VTAIL.n31 B 0.031665f
C284 VTAIL.n32 B 0.031665f
C285 VTAIL.n33 B 0.031665f
C286 VTAIL.n34 B 0.014185f
C287 VTAIL.n35 B 0.013396f
C288 VTAIL.n36 B 0.02493f
C289 VTAIL.n37 B 0.02493f
C290 VTAIL.n38 B 0.013396f
C291 VTAIL.n39 B 0.01379f
C292 VTAIL.n40 B 0.01379f
C293 VTAIL.n41 B 0.031665f
C294 VTAIL.n42 B 0.062599f
C295 VTAIL.n43 B 0.014185f
C296 VTAIL.n44 B 0.013396f
C297 VTAIL.n45 B 0.057625f
C298 VTAIL.n46 B 0.034415f
C299 VTAIL.n47 B 0.344695f
C300 VTAIL.t8 B 0.167851f
C301 VTAIL.t7 B 0.167851f
C302 VTAIL.n48 B 1.3904f
C303 VTAIL.n49 B 1.73627f
C304 VTAIL.t4 B 0.167851f
C305 VTAIL.t2 B 0.167851f
C306 VTAIL.n50 B 1.39041f
C307 VTAIL.n51 B 1.73626f
C308 VTAIL.n52 B 0.031678f
C309 VTAIL.n53 B 0.02493f
C310 VTAIL.n54 B 0.013396f
C311 VTAIL.n55 B 0.031665f
C312 VTAIL.n56 B 0.014185f
C313 VTAIL.n57 B 0.02493f
C314 VTAIL.n58 B 0.013396f
C315 VTAIL.n59 B 0.031665f
C316 VTAIL.n60 B 0.031665f
C317 VTAIL.n61 B 0.014185f
C318 VTAIL.n62 B 0.02493f
C319 VTAIL.n63 B 0.013396f
C320 VTAIL.n64 B 0.031665f
C321 VTAIL.n65 B 0.014185f
C322 VTAIL.n66 B 0.146449f
C323 VTAIL.t3 B 0.053018f
C324 VTAIL.n67 B 0.023748f
C325 VTAIL.n68 B 0.022384f
C326 VTAIL.n69 B 0.013396f
C327 VTAIL.n70 B 0.871792f
C328 VTAIL.n71 B 0.02493f
C329 VTAIL.n72 B 0.013396f
C330 VTAIL.n73 B 0.014185f
C331 VTAIL.n74 B 0.031665f
C332 VTAIL.n75 B 0.031665f
C333 VTAIL.n76 B 0.014185f
C334 VTAIL.n77 B 0.013396f
C335 VTAIL.n78 B 0.02493f
C336 VTAIL.n79 B 0.02493f
C337 VTAIL.n80 B 0.013396f
C338 VTAIL.n81 B 0.014185f
C339 VTAIL.n82 B 0.031665f
C340 VTAIL.n83 B 0.031665f
C341 VTAIL.n84 B 0.014185f
C342 VTAIL.n85 B 0.013396f
C343 VTAIL.n86 B 0.02493f
C344 VTAIL.n87 B 0.02493f
C345 VTAIL.n88 B 0.013396f
C346 VTAIL.n89 B 0.01379f
C347 VTAIL.n90 B 0.01379f
C348 VTAIL.n91 B 0.031665f
C349 VTAIL.n92 B 0.062599f
C350 VTAIL.n93 B 0.014185f
C351 VTAIL.n94 B 0.013396f
C352 VTAIL.n95 B 0.057625f
C353 VTAIL.n96 B 0.034415f
C354 VTAIL.n97 B 0.344695f
C355 VTAIL.t9 B 0.167851f
C356 VTAIL.t5 B 0.167851f
C357 VTAIL.n98 B 1.39041f
C358 VTAIL.n99 B 0.559669f
C359 VTAIL.n100 B 0.031678f
C360 VTAIL.n101 B 0.02493f
C361 VTAIL.n102 B 0.013396f
C362 VTAIL.n103 B 0.031665f
C363 VTAIL.n104 B 0.014185f
C364 VTAIL.n105 B 0.02493f
C365 VTAIL.n106 B 0.013396f
C366 VTAIL.n107 B 0.031665f
C367 VTAIL.n108 B 0.031665f
C368 VTAIL.n109 B 0.014185f
C369 VTAIL.n110 B 0.02493f
C370 VTAIL.n111 B 0.013396f
C371 VTAIL.n112 B 0.031665f
C372 VTAIL.n113 B 0.014185f
C373 VTAIL.n114 B 0.146449f
C374 VTAIL.t6 B 0.053018f
C375 VTAIL.n115 B 0.023748f
C376 VTAIL.n116 B 0.022384f
C377 VTAIL.n117 B 0.013396f
C378 VTAIL.n118 B 0.871792f
C379 VTAIL.n119 B 0.02493f
C380 VTAIL.n120 B 0.013396f
C381 VTAIL.n121 B 0.014185f
C382 VTAIL.n122 B 0.031665f
C383 VTAIL.n123 B 0.031665f
C384 VTAIL.n124 B 0.014185f
C385 VTAIL.n125 B 0.013396f
C386 VTAIL.n126 B 0.02493f
C387 VTAIL.n127 B 0.02493f
C388 VTAIL.n128 B 0.013396f
C389 VTAIL.n129 B 0.014185f
C390 VTAIL.n130 B 0.031665f
C391 VTAIL.n131 B 0.031665f
C392 VTAIL.n132 B 0.014185f
C393 VTAIL.n133 B 0.013396f
C394 VTAIL.n134 B 0.02493f
C395 VTAIL.n135 B 0.02493f
C396 VTAIL.n136 B 0.013396f
C397 VTAIL.n137 B 0.01379f
C398 VTAIL.n138 B 0.01379f
C399 VTAIL.n139 B 0.031665f
C400 VTAIL.n140 B 0.062599f
C401 VTAIL.n141 B 0.014185f
C402 VTAIL.n142 B 0.013396f
C403 VTAIL.n143 B 0.057625f
C404 VTAIL.n144 B 0.034415f
C405 VTAIL.n145 B 1.33084f
C406 VTAIL.n146 B 0.031678f
C407 VTAIL.n147 B 0.02493f
C408 VTAIL.n148 B 0.013396f
C409 VTAIL.n149 B 0.031665f
C410 VTAIL.n150 B 0.014185f
C411 VTAIL.n151 B 0.02493f
C412 VTAIL.n152 B 0.013396f
C413 VTAIL.n153 B 0.031665f
C414 VTAIL.n154 B 0.014185f
C415 VTAIL.n155 B 0.02493f
C416 VTAIL.n156 B 0.013396f
C417 VTAIL.n157 B 0.031665f
C418 VTAIL.n158 B 0.014185f
C419 VTAIL.n159 B 0.146449f
C420 VTAIL.t1 B 0.053018f
C421 VTAIL.n160 B 0.023748f
C422 VTAIL.n161 B 0.022384f
C423 VTAIL.n162 B 0.013396f
C424 VTAIL.n163 B 0.871792f
C425 VTAIL.n164 B 0.02493f
C426 VTAIL.n165 B 0.013396f
C427 VTAIL.n166 B 0.014185f
C428 VTAIL.n167 B 0.031665f
C429 VTAIL.n168 B 0.031665f
C430 VTAIL.n169 B 0.014185f
C431 VTAIL.n170 B 0.013396f
C432 VTAIL.n171 B 0.02493f
C433 VTAIL.n172 B 0.02493f
C434 VTAIL.n173 B 0.013396f
C435 VTAIL.n174 B 0.014185f
C436 VTAIL.n175 B 0.031665f
C437 VTAIL.n176 B 0.031665f
C438 VTAIL.n177 B 0.031665f
C439 VTAIL.n178 B 0.014185f
C440 VTAIL.n179 B 0.013396f
C441 VTAIL.n180 B 0.02493f
C442 VTAIL.n181 B 0.02493f
C443 VTAIL.n182 B 0.013396f
C444 VTAIL.n183 B 0.01379f
C445 VTAIL.n184 B 0.01379f
C446 VTAIL.n185 B 0.031665f
C447 VTAIL.n186 B 0.062599f
C448 VTAIL.n187 B 0.014185f
C449 VTAIL.n188 B 0.013396f
C450 VTAIL.n189 B 0.057625f
C451 VTAIL.n190 B 0.034415f
C452 VTAIL.n191 B 1.27856f
C453 VP.n0 B 0.034308f
C454 VP.t3 B 1.44489f
C455 VP.n1 B 0.026709f
C456 VP.n2 B 0.026024f
C457 VP.t4 B 1.44489f
C458 VP.n3 B 0.048259f
C459 VP.n4 B 0.026024f
C460 VP.n5 B 0.036347f
C461 VP.n6 B 0.034308f
C462 VP.t5 B 1.44489f
C463 VP.n7 B 0.026709f
C464 VP.n8 B 0.246792f
C465 VP.t2 B 1.44489f
C466 VP.t0 B 1.64114f
C467 VP.n9 B 0.575002f
C468 VP.n10 B 0.610607f
C469 VP.n11 B 0.048259f
C470 VP.n12 B 0.046226f
C471 VP.n13 B 0.026024f
C472 VP.n14 B 0.026024f
C473 VP.n15 B 0.026024f
C474 VP.n16 B 0.050983f
C475 VP.n17 B 0.036347f
C476 VP.n18 B 0.608731f
C477 VP.n19 B 1.2467f
C478 VP.t1 B 1.44489f
C479 VP.n20 B 0.608731f
C480 VP.n21 B 1.26739f
C481 VP.n22 B 0.034308f
C482 VP.n23 B 0.026024f
C483 VP.n24 B 0.050983f
C484 VP.n25 B 0.026709f
C485 VP.n26 B 0.046226f
C486 VP.n27 B 0.026024f
C487 VP.n28 B 0.026024f
C488 VP.n29 B 0.026024f
C489 VP.n30 B 0.549499f
C490 VP.n31 B 0.048259f
C491 VP.n32 B 0.046226f
C492 VP.n33 B 0.026024f
C493 VP.n34 B 0.026024f
C494 VP.n35 B 0.026024f
C495 VP.n36 B 0.050983f
C496 VP.n37 B 0.036347f
C497 VP.n38 B 0.608731f
C498 VP.n39 B 0.039418f
.ends

