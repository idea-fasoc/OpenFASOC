* NGSPICE file created from diff_pair_sample_1519.ext - technology: sky130A

.subckt diff_pair_sample_1519 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=0 ps=0 w=4.64 l=3.96
X1 B.t8 B.t6 B.t7 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=0 ps=0 w=4.64 l=3.96
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=1.8096 ps=10.06 w=4.64 l=3.96
X3 B.t5 B.t3 B.t4 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=0 ps=0 w=4.64 l=3.96
X4 VDD1.t1 VP.t0 VTAIL.t1 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=1.8096 ps=10.06 w=4.64 l=3.96
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=1.8096 ps=10.06 w=4.64 l=3.96
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=1.8096 ps=10.06 w=4.64 l=3.96
X7 B.t2 B.t0 B.t1 w_n2686_n1896# sky130_fd_pr__pfet_01v8 ad=1.8096 pd=10.06 as=0 ps=0 w=4.64 l=3.96
R0 B.n249 B.n82 585
R1 B.n248 B.n247 585
R2 B.n246 B.n83 585
R3 B.n245 B.n244 585
R4 B.n243 B.n84 585
R5 B.n242 B.n241 585
R6 B.n240 B.n85 585
R7 B.n239 B.n238 585
R8 B.n237 B.n86 585
R9 B.n236 B.n235 585
R10 B.n234 B.n87 585
R11 B.n233 B.n232 585
R12 B.n231 B.n88 585
R13 B.n230 B.n229 585
R14 B.n228 B.n89 585
R15 B.n227 B.n226 585
R16 B.n225 B.n90 585
R17 B.n224 B.n223 585
R18 B.n222 B.n91 585
R19 B.n221 B.n220 585
R20 B.n218 B.n92 585
R21 B.n217 B.n216 585
R22 B.n215 B.n95 585
R23 B.n214 B.n213 585
R24 B.n212 B.n96 585
R25 B.n211 B.n210 585
R26 B.n209 B.n97 585
R27 B.n208 B.n207 585
R28 B.n206 B.n98 585
R29 B.n204 B.n203 585
R30 B.n202 B.n101 585
R31 B.n201 B.n200 585
R32 B.n199 B.n102 585
R33 B.n198 B.n197 585
R34 B.n196 B.n103 585
R35 B.n195 B.n194 585
R36 B.n193 B.n104 585
R37 B.n192 B.n191 585
R38 B.n190 B.n105 585
R39 B.n189 B.n188 585
R40 B.n187 B.n106 585
R41 B.n186 B.n185 585
R42 B.n184 B.n107 585
R43 B.n183 B.n182 585
R44 B.n181 B.n108 585
R45 B.n180 B.n179 585
R46 B.n178 B.n109 585
R47 B.n177 B.n176 585
R48 B.n175 B.n110 585
R49 B.n251 B.n250 585
R50 B.n252 B.n81 585
R51 B.n254 B.n253 585
R52 B.n255 B.n80 585
R53 B.n257 B.n256 585
R54 B.n258 B.n79 585
R55 B.n260 B.n259 585
R56 B.n261 B.n78 585
R57 B.n263 B.n262 585
R58 B.n264 B.n77 585
R59 B.n266 B.n265 585
R60 B.n267 B.n76 585
R61 B.n269 B.n268 585
R62 B.n270 B.n75 585
R63 B.n272 B.n271 585
R64 B.n273 B.n74 585
R65 B.n275 B.n274 585
R66 B.n276 B.n73 585
R67 B.n278 B.n277 585
R68 B.n279 B.n72 585
R69 B.n281 B.n280 585
R70 B.n282 B.n71 585
R71 B.n284 B.n283 585
R72 B.n285 B.n70 585
R73 B.n287 B.n286 585
R74 B.n288 B.n69 585
R75 B.n290 B.n289 585
R76 B.n291 B.n68 585
R77 B.n293 B.n292 585
R78 B.n294 B.n67 585
R79 B.n296 B.n295 585
R80 B.n297 B.n66 585
R81 B.n299 B.n298 585
R82 B.n300 B.n65 585
R83 B.n302 B.n301 585
R84 B.n303 B.n64 585
R85 B.n305 B.n304 585
R86 B.n306 B.n63 585
R87 B.n308 B.n307 585
R88 B.n309 B.n62 585
R89 B.n311 B.n310 585
R90 B.n312 B.n61 585
R91 B.n314 B.n313 585
R92 B.n315 B.n60 585
R93 B.n317 B.n316 585
R94 B.n318 B.n59 585
R95 B.n320 B.n319 585
R96 B.n321 B.n58 585
R97 B.n323 B.n322 585
R98 B.n324 B.n57 585
R99 B.n326 B.n325 585
R100 B.n327 B.n56 585
R101 B.n329 B.n328 585
R102 B.n330 B.n55 585
R103 B.n332 B.n331 585
R104 B.n333 B.n54 585
R105 B.n335 B.n334 585
R106 B.n336 B.n53 585
R107 B.n338 B.n337 585
R108 B.n339 B.n52 585
R109 B.n341 B.n340 585
R110 B.n342 B.n51 585
R111 B.n344 B.n343 585
R112 B.n345 B.n50 585
R113 B.n347 B.n346 585
R114 B.n348 B.n49 585
R115 B.n350 B.n349 585
R116 B.n351 B.n48 585
R117 B.n426 B.n425 585
R118 B.n424 B.n19 585
R119 B.n423 B.n422 585
R120 B.n421 B.n20 585
R121 B.n420 B.n419 585
R122 B.n418 B.n21 585
R123 B.n417 B.n416 585
R124 B.n415 B.n22 585
R125 B.n414 B.n413 585
R126 B.n412 B.n23 585
R127 B.n411 B.n410 585
R128 B.n409 B.n24 585
R129 B.n408 B.n407 585
R130 B.n406 B.n25 585
R131 B.n405 B.n404 585
R132 B.n403 B.n26 585
R133 B.n402 B.n401 585
R134 B.n400 B.n27 585
R135 B.n399 B.n398 585
R136 B.n397 B.n28 585
R137 B.n396 B.n395 585
R138 B.n394 B.n29 585
R139 B.n393 B.n392 585
R140 B.n391 B.n33 585
R141 B.n390 B.n389 585
R142 B.n388 B.n34 585
R143 B.n387 B.n386 585
R144 B.n385 B.n35 585
R145 B.n384 B.n383 585
R146 B.n381 B.n36 585
R147 B.n380 B.n379 585
R148 B.n378 B.n39 585
R149 B.n377 B.n376 585
R150 B.n375 B.n40 585
R151 B.n374 B.n373 585
R152 B.n372 B.n41 585
R153 B.n371 B.n370 585
R154 B.n369 B.n42 585
R155 B.n368 B.n367 585
R156 B.n366 B.n43 585
R157 B.n365 B.n364 585
R158 B.n363 B.n44 585
R159 B.n362 B.n361 585
R160 B.n360 B.n45 585
R161 B.n359 B.n358 585
R162 B.n357 B.n46 585
R163 B.n356 B.n355 585
R164 B.n354 B.n47 585
R165 B.n353 B.n352 585
R166 B.n427 B.n18 585
R167 B.n429 B.n428 585
R168 B.n430 B.n17 585
R169 B.n432 B.n431 585
R170 B.n433 B.n16 585
R171 B.n435 B.n434 585
R172 B.n436 B.n15 585
R173 B.n438 B.n437 585
R174 B.n439 B.n14 585
R175 B.n441 B.n440 585
R176 B.n442 B.n13 585
R177 B.n444 B.n443 585
R178 B.n445 B.n12 585
R179 B.n447 B.n446 585
R180 B.n448 B.n11 585
R181 B.n450 B.n449 585
R182 B.n451 B.n10 585
R183 B.n453 B.n452 585
R184 B.n454 B.n9 585
R185 B.n456 B.n455 585
R186 B.n457 B.n8 585
R187 B.n459 B.n458 585
R188 B.n460 B.n7 585
R189 B.n462 B.n461 585
R190 B.n463 B.n6 585
R191 B.n465 B.n464 585
R192 B.n466 B.n5 585
R193 B.n468 B.n467 585
R194 B.n469 B.n4 585
R195 B.n471 B.n470 585
R196 B.n472 B.n3 585
R197 B.n474 B.n473 585
R198 B.n475 B.n0 585
R199 B.n2 B.n1 585
R200 B.n127 B.n126 585
R201 B.n129 B.n128 585
R202 B.n130 B.n125 585
R203 B.n132 B.n131 585
R204 B.n133 B.n124 585
R205 B.n135 B.n134 585
R206 B.n136 B.n123 585
R207 B.n138 B.n137 585
R208 B.n139 B.n122 585
R209 B.n141 B.n140 585
R210 B.n142 B.n121 585
R211 B.n144 B.n143 585
R212 B.n145 B.n120 585
R213 B.n147 B.n146 585
R214 B.n148 B.n119 585
R215 B.n150 B.n149 585
R216 B.n151 B.n118 585
R217 B.n153 B.n152 585
R218 B.n154 B.n117 585
R219 B.n156 B.n155 585
R220 B.n157 B.n116 585
R221 B.n159 B.n158 585
R222 B.n160 B.n115 585
R223 B.n162 B.n161 585
R224 B.n163 B.n114 585
R225 B.n165 B.n164 585
R226 B.n166 B.n113 585
R227 B.n168 B.n167 585
R228 B.n169 B.n112 585
R229 B.n171 B.n170 585
R230 B.n172 B.n111 585
R231 B.n174 B.n173 585
R232 B.n173 B.n110 516.524
R233 B.n251 B.n82 516.524
R234 B.n353 B.n48 516.524
R235 B.n427 B.n426 516.524
R236 B.n93 B.t4 328.32
R237 B.n37 B.t8 328.32
R238 B.n99 B.t1 328.32
R239 B.n30 B.t11 328.32
R240 B.n477 B.n476 256.663
R241 B.n94 B.t5 245.12
R242 B.n38 B.t7 245.12
R243 B.n100 B.t2 245.12
R244 B.n31 B.t10 245.12
R245 B.n99 B.t0 237.702
R246 B.n93 B.t3 237.702
R247 B.n37 B.t6 237.702
R248 B.n30 B.t9 237.702
R249 B.n476 B.n475 235.042
R250 B.n476 B.n2 235.042
R251 B.n177 B.n110 163.367
R252 B.n178 B.n177 163.367
R253 B.n179 B.n178 163.367
R254 B.n179 B.n108 163.367
R255 B.n183 B.n108 163.367
R256 B.n184 B.n183 163.367
R257 B.n185 B.n184 163.367
R258 B.n185 B.n106 163.367
R259 B.n189 B.n106 163.367
R260 B.n190 B.n189 163.367
R261 B.n191 B.n190 163.367
R262 B.n191 B.n104 163.367
R263 B.n195 B.n104 163.367
R264 B.n196 B.n195 163.367
R265 B.n197 B.n196 163.367
R266 B.n197 B.n102 163.367
R267 B.n201 B.n102 163.367
R268 B.n202 B.n201 163.367
R269 B.n203 B.n202 163.367
R270 B.n203 B.n98 163.367
R271 B.n208 B.n98 163.367
R272 B.n209 B.n208 163.367
R273 B.n210 B.n209 163.367
R274 B.n210 B.n96 163.367
R275 B.n214 B.n96 163.367
R276 B.n215 B.n214 163.367
R277 B.n216 B.n215 163.367
R278 B.n216 B.n92 163.367
R279 B.n221 B.n92 163.367
R280 B.n222 B.n221 163.367
R281 B.n223 B.n222 163.367
R282 B.n223 B.n90 163.367
R283 B.n227 B.n90 163.367
R284 B.n228 B.n227 163.367
R285 B.n229 B.n228 163.367
R286 B.n229 B.n88 163.367
R287 B.n233 B.n88 163.367
R288 B.n234 B.n233 163.367
R289 B.n235 B.n234 163.367
R290 B.n235 B.n86 163.367
R291 B.n239 B.n86 163.367
R292 B.n240 B.n239 163.367
R293 B.n241 B.n240 163.367
R294 B.n241 B.n84 163.367
R295 B.n245 B.n84 163.367
R296 B.n246 B.n245 163.367
R297 B.n247 B.n246 163.367
R298 B.n247 B.n82 163.367
R299 B.n349 B.n48 163.367
R300 B.n349 B.n348 163.367
R301 B.n348 B.n347 163.367
R302 B.n347 B.n50 163.367
R303 B.n343 B.n50 163.367
R304 B.n343 B.n342 163.367
R305 B.n342 B.n341 163.367
R306 B.n341 B.n52 163.367
R307 B.n337 B.n52 163.367
R308 B.n337 B.n336 163.367
R309 B.n336 B.n335 163.367
R310 B.n335 B.n54 163.367
R311 B.n331 B.n54 163.367
R312 B.n331 B.n330 163.367
R313 B.n330 B.n329 163.367
R314 B.n329 B.n56 163.367
R315 B.n325 B.n56 163.367
R316 B.n325 B.n324 163.367
R317 B.n324 B.n323 163.367
R318 B.n323 B.n58 163.367
R319 B.n319 B.n58 163.367
R320 B.n319 B.n318 163.367
R321 B.n318 B.n317 163.367
R322 B.n317 B.n60 163.367
R323 B.n313 B.n60 163.367
R324 B.n313 B.n312 163.367
R325 B.n312 B.n311 163.367
R326 B.n311 B.n62 163.367
R327 B.n307 B.n62 163.367
R328 B.n307 B.n306 163.367
R329 B.n306 B.n305 163.367
R330 B.n305 B.n64 163.367
R331 B.n301 B.n64 163.367
R332 B.n301 B.n300 163.367
R333 B.n300 B.n299 163.367
R334 B.n299 B.n66 163.367
R335 B.n295 B.n66 163.367
R336 B.n295 B.n294 163.367
R337 B.n294 B.n293 163.367
R338 B.n293 B.n68 163.367
R339 B.n289 B.n68 163.367
R340 B.n289 B.n288 163.367
R341 B.n288 B.n287 163.367
R342 B.n287 B.n70 163.367
R343 B.n283 B.n70 163.367
R344 B.n283 B.n282 163.367
R345 B.n282 B.n281 163.367
R346 B.n281 B.n72 163.367
R347 B.n277 B.n72 163.367
R348 B.n277 B.n276 163.367
R349 B.n276 B.n275 163.367
R350 B.n275 B.n74 163.367
R351 B.n271 B.n74 163.367
R352 B.n271 B.n270 163.367
R353 B.n270 B.n269 163.367
R354 B.n269 B.n76 163.367
R355 B.n265 B.n76 163.367
R356 B.n265 B.n264 163.367
R357 B.n264 B.n263 163.367
R358 B.n263 B.n78 163.367
R359 B.n259 B.n78 163.367
R360 B.n259 B.n258 163.367
R361 B.n258 B.n257 163.367
R362 B.n257 B.n80 163.367
R363 B.n253 B.n80 163.367
R364 B.n253 B.n252 163.367
R365 B.n252 B.n251 163.367
R366 B.n426 B.n19 163.367
R367 B.n422 B.n19 163.367
R368 B.n422 B.n421 163.367
R369 B.n421 B.n420 163.367
R370 B.n420 B.n21 163.367
R371 B.n416 B.n21 163.367
R372 B.n416 B.n415 163.367
R373 B.n415 B.n414 163.367
R374 B.n414 B.n23 163.367
R375 B.n410 B.n23 163.367
R376 B.n410 B.n409 163.367
R377 B.n409 B.n408 163.367
R378 B.n408 B.n25 163.367
R379 B.n404 B.n25 163.367
R380 B.n404 B.n403 163.367
R381 B.n403 B.n402 163.367
R382 B.n402 B.n27 163.367
R383 B.n398 B.n27 163.367
R384 B.n398 B.n397 163.367
R385 B.n397 B.n396 163.367
R386 B.n396 B.n29 163.367
R387 B.n392 B.n29 163.367
R388 B.n392 B.n391 163.367
R389 B.n391 B.n390 163.367
R390 B.n390 B.n34 163.367
R391 B.n386 B.n34 163.367
R392 B.n386 B.n385 163.367
R393 B.n385 B.n384 163.367
R394 B.n384 B.n36 163.367
R395 B.n379 B.n36 163.367
R396 B.n379 B.n378 163.367
R397 B.n378 B.n377 163.367
R398 B.n377 B.n40 163.367
R399 B.n373 B.n40 163.367
R400 B.n373 B.n372 163.367
R401 B.n372 B.n371 163.367
R402 B.n371 B.n42 163.367
R403 B.n367 B.n42 163.367
R404 B.n367 B.n366 163.367
R405 B.n366 B.n365 163.367
R406 B.n365 B.n44 163.367
R407 B.n361 B.n44 163.367
R408 B.n361 B.n360 163.367
R409 B.n360 B.n359 163.367
R410 B.n359 B.n46 163.367
R411 B.n355 B.n46 163.367
R412 B.n355 B.n354 163.367
R413 B.n354 B.n353 163.367
R414 B.n428 B.n427 163.367
R415 B.n428 B.n17 163.367
R416 B.n432 B.n17 163.367
R417 B.n433 B.n432 163.367
R418 B.n434 B.n433 163.367
R419 B.n434 B.n15 163.367
R420 B.n438 B.n15 163.367
R421 B.n439 B.n438 163.367
R422 B.n440 B.n439 163.367
R423 B.n440 B.n13 163.367
R424 B.n444 B.n13 163.367
R425 B.n445 B.n444 163.367
R426 B.n446 B.n445 163.367
R427 B.n446 B.n11 163.367
R428 B.n450 B.n11 163.367
R429 B.n451 B.n450 163.367
R430 B.n452 B.n451 163.367
R431 B.n452 B.n9 163.367
R432 B.n456 B.n9 163.367
R433 B.n457 B.n456 163.367
R434 B.n458 B.n457 163.367
R435 B.n458 B.n7 163.367
R436 B.n462 B.n7 163.367
R437 B.n463 B.n462 163.367
R438 B.n464 B.n463 163.367
R439 B.n464 B.n5 163.367
R440 B.n468 B.n5 163.367
R441 B.n469 B.n468 163.367
R442 B.n470 B.n469 163.367
R443 B.n470 B.n3 163.367
R444 B.n474 B.n3 163.367
R445 B.n475 B.n474 163.367
R446 B.n126 B.n2 163.367
R447 B.n129 B.n126 163.367
R448 B.n130 B.n129 163.367
R449 B.n131 B.n130 163.367
R450 B.n131 B.n124 163.367
R451 B.n135 B.n124 163.367
R452 B.n136 B.n135 163.367
R453 B.n137 B.n136 163.367
R454 B.n137 B.n122 163.367
R455 B.n141 B.n122 163.367
R456 B.n142 B.n141 163.367
R457 B.n143 B.n142 163.367
R458 B.n143 B.n120 163.367
R459 B.n147 B.n120 163.367
R460 B.n148 B.n147 163.367
R461 B.n149 B.n148 163.367
R462 B.n149 B.n118 163.367
R463 B.n153 B.n118 163.367
R464 B.n154 B.n153 163.367
R465 B.n155 B.n154 163.367
R466 B.n155 B.n116 163.367
R467 B.n159 B.n116 163.367
R468 B.n160 B.n159 163.367
R469 B.n161 B.n160 163.367
R470 B.n161 B.n114 163.367
R471 B.n165 B.n114 163.367
R472 B.n166 B.n165 163.367
R473 B.n167 B.n166 163.367
R474 B.n167 B.n112 163.367
R475 B.n171 B.n112 163.367
R476 B.n172 B.n171 163.367
R477 B.n173 B.n172 163.367
R478 B.n100 B.n99 83.2005
R479 B.n94 B.n93 83.2005
R480 B.n38 B.n37 83.2005
R481 B.n31 B.n30 83.2005
R482 B.n205 B.n100 59.5399
R483 B.n219 B.n94 59.5399
R484 B.n382 B.n38 59.5399
R485 B.n32 B.n31 59.5399
R486 B.n425 B.n18 33.5615
R487 B.n352 B.n351 33.5615
R488 B.n250 B.n249 33.5615
R489 B.n175 B.n174 33.5615
R490 B B.n477 18.0485
R491 B.n429 B.n18 10.6151
R492 B.n430 B.n429 10.6151
R493 B.n431 B.n430 10.6151
R494 B.n431 B.n16 10.6151
R495 B.n435 B.n16 10.6151
R496 B.n436 B.n435 10.6151
R497 B.n437 B.n436 10.6151
R498 B.n437 B.n14 10.6151
R499 B.n441 B.n14 10.6151
R500 B.n442 B.n441 10.6151
R501 B.n443 B.n442 10.6151
R502 B.n443 B.n12 10.6151
R503 B.n447 B.n12 10.6151
R504 B.n448 B.n447 10.6151
R505 B.n449 B.n448 10.6151
R506 B.n449 B.n10 10.6151
R507 B.n453 B.n10 10.6151
R508 B.n454 B.n453 10.6151
R509 B.n455 B.n454 10.6151
R510 B.n455 B.n8 10.6151
R511 B.n459 B.n8 10.6151
R512 B.n460 B.n459 10.6151
R513 B.n461 B.n460 10.6151
R514 B.n461 B.n6 10.6151
R515 B.n465 B.n6 10.6151
R516 B.n466 B.n465 10.6151
R517 B.n467 B.n466 10.6151
R518 B.n467 B.n4 10.6151
R519 B.n471 B.n4 10.6151
R520 B.n472 B.n471 10.6151
R521 B.n473 B.n472 10.6151
R522 B.n473 B.n0 10.6151
R523 B.n425 B.n424 10.6151
R524 B.n424 B.n423 10.6151
R525 B.n423 B.n20 10.6151
R526 B.n419 B.n20 10.6151
R527 B.n419 B.n418 10.6151
R528 B.n418 B.n417 10.6151
R529 B.n417 B.n22 10.6151
R530 B.n413 B.n22 10.6151
R531 B.n413 B.n412 10.6151
R532 B.n412 B.n411 10.6151
R533 B.n411 B.n24 10.6151
R534 B.n407 B.n24 10.6151
R535 B.n407 B.n406 10.6151
R536 B.n406 B.n405 10.6151
R537 B.n405 B.n26 10.6151
R538 B.n401 B.n26 10.6151
R539 B.n401 B.n400 10.6151
R540 B.n400 B.n399 10.6151
R541 B.n399 B.n28 10.6151
R542 B.n395 B.n394 10.6151
R543 B.n394 B.n393 10.6151
R544 B.n393 B.n33 10.6151
R545 B.n389 B.n33 10.6151
R546 B.n389 B.n388 10.6151
R547 B.n388 B.n387 10.6151
R548 B.n387 B.n35 10.6151
R549 B.n383 B.n35 10.6151
R550 B.n381 B.n380 10.6151
R551 B.n380 B.n39 10.6151
R552 B.n376 B.n39 10.6151
R553 B.n376 B.n375 10.6151
R554 B.n375 B.n374 10.6151
R555 B.n374 B.n41 10.6151
R556 B.n370 B.n41 10.6151
R557 B.n370 B.n369 10.6151
R558 B.n369 B.n368 10.6151
R559 B.n368 B.n43 10.6151
R560 B.n364 B.n43 10.6151
R561 B.n364 B.n363 10.6151
R562 B.n363 B.n362 10.6151
R563 B.n362 B.n45 10.6151
R564 B.n358 B.n45 10.6151
R565 B.n358 B.n357 10.6151
R566 B.n357 B.n356 10.6151
R567 B.n356 B.n47 10.6151
R568 B.n352 B.n47 10.6151
R569 B.n351 B.n350 10.6151
R570 B.n350 B.n49 10.6151
R571 B.n346 B.n49 10.6151
R572 B.n346 B.n345 10.6151
R573 B.n345 B.n344 10.6151
R574 B.n344 B.n51 10.6151
R575 B.n340 B.n51 10.6151
R576 B.n340 B.n339 10.6151
R577 B.n339 B.n338 10.6151
R578 B.n338 B.n53 10.6151
R579 B.n334 B.n53 10.6151
R580 B.n334 B.n333 10.6151
R581 B.n333 B.n332 10.6151
R582 B.n332 B.n55 10.6151
R583 B.n328 B.n55 10.6151
R584 B.n328 B.n327 10.6151
R585 B.n327 B.n326 10.6151
R586 B.n326 B.n57 10.6151
R587 B.n322 B.n57 10.6151
R588 B.n322 B.n321 10.6151
R589 B.n321 B.n320 10.6151
R590 B.n320 B.n59 10.6151
R591 B.n316 B.n59 10.6151
R592 B.n316 B.n315 10.6151
R593 B.n315 B.n314 10.6151
R594 B.n314 B.n61 10.6151
R595 B.n310 B.n61 10.6151
R596 B.n310 B.n309 10.6151
R597 B.n309 B.n308 10.6151
R598 B.n308 B.n63 10.6151
R599 B.n304 B.n63 10.6151
R600 B.n304 B.n303 10.6151
R601 B.n303 B.n302 10.6151
R602 B.n302 B.n65 10.6151
R603 B.n298 B.n65 10.6151
R604 B.n298 B.n297 10.6151
R605 B.n297 B.n296 10.6151
R606 B.n296 B.n67 10.6151
R607 B.n292 B.n67 10.6151
R608 B.n292 B.n291 10.6151
R609 B.n291 B.n290 10.6151
R610 B.n290 B.n69 10.6151
R611 B.n286 B.n69 10.6151
R612 B.n286 B.n285 10.6151
R613 B.n285 B.n284 10.6151
R614 B.n284 B.n71 10.6151
R615 B.n280 B.n71 10.6151
R616 B.n280 B.n279 10.6151
R617 B.n279 B.n278 10.6151
R618 B.n278 B.n73 10.6151
R619 B.n274 B.n73 10.6151
R620 B.n274 B.n273 10.6151
R621 B.n273 B.n272 10.6151
R622 B.n272 B.n75 10.6151
R623 B.n268 B.n75 10.6151
R624 B.n268 B.n267 10.6151
R625 B.n267 B.n266 10.6151
R626 B.n266 B.n77 10.6151
R627 B.n262 B.n77 10.6151
R628 B.n262 B.n261 10.6151
R629 B.n261 B.n260 10.6151
R630 B.n260 B.n79 10.6151
R631 B.n256 B.n79 10.6151
R632 B.n256 B.n255 10.6151
R633 B.n255 B.n254 10.6151
R634 B.n254 B.n81 10.6151
R635 B.n250 B.n81 10.6151
R636 B.n127 B.n1 10.6151
R637 B.n128 B.n127 10.6151
R638 B.n128 B.n125 10.6151
R639 B.n132 B.n125 10.6151
R640 B.n133 B.n132 10.6151
R641 B.n134 B.n133 10.6151
R642 B.n134 B.n123 10.6151
R643 B.n138 B.n123 10.6151
R644 B.n139 B.n138 10.6151
R645 B.n140 B.n139 10.6151
R646 B.n140 B.n121 10.6151
R647 B.n144 B.n121 10.6151
R648 B.n145 B.n144 10.6151
R649 B.n146 B.n145 10.6151
R650 B.n146 B.n119 10.6151
R651 B.n150 B.n119 10.6151
R652 B.n151 B.n150 10.6151
R653 B.n152 B.n151 10.6151
R654 B.n152 B.n117 10.6151
R655 B.n156 B.n117 10.6151
R656 B.n157 B.n156 10.6151
R657 B.n158 B.n157 10.6151
R658 B.n158 B.n115 10.6151
R659 B.n162 B.n115 10.6151
R660 B.n163 B.n162 10.6151
R661 B.n164 B.n163 10.6151
R662 B.n164 B.n113 10.6151
R663 B.n168 B.n113 10.6151
R664 B.n169 B.n168 10.6151
R665 B.n170 B.n169 10.6151
R666 B.n170 B.n111 10.6151
R667 B.n174 B.n111 10.6151
R668 B.n176 B.n175 10.6151
R669 B.n176 B.n109 10.6151
R670 B.n180 B.n109 10.6151
R671 B.n181 B.n180 10.6151
R672 B.n182 B.n181 10.6151
R673 B.n182 B.n107 10.6151
R674 B.n186 B.n107 10.6151
R675 B.n187 B.n186 10.6151
R676 B.n188 B.n187 10.6151
R677 B.n188 B.n105 10.6151
R678 B.n192 B.n105 10.6151
R679 B.n193 B.n192 10.6151
R680 B.n194 B.n193 10.6151
R681 B.n194 B.n103 10.6151
R682 B.n198 B.n103 10.6151
R683 B.n199 B.n198 10.6151
R684 B.n200 B.n199 10.6151
R685 B.n200 B.n101 10.6151
R686 B.n204 B.n101 10.6151
R687 B.n207 B.n206 10.6151
R688 B.n207 B.n97 10.6151
R689 B.n211 B.n97 10.6151
R690 B.n212 B.n211 10.6151
R691 B.n213 B.n212 10.6151
R692 B.n213 B.n95 10.6151
R693 B.n217 B.n95 10.6151
R694 B.n218 B.n217 10.6151
R695 B.n220 B.n91 10.6151
R696 B.n224 B.n91 10.6151
R697 B.n225 B.n224 10.6151
R698 B.n226 B.n225 10.6151
R699 B.n226 B.n89 10.6151
R700 B.n230 B.n89 10.6151
R701 B.n231 B.n230 10.6151
R702 B.n232 B.n231 10.6151
R703 B.n232 B.n87 10.6151
R704 B.n236 B.n87 10.6151
R705 B.n237 B.n236 10.6151
R706 B.n238 B.n237 10.6151
R707 B.n238 B.n85 10.6151
R708 B.n242 B.n85 10.6151
R709 B.n243 B.n242 10.6151
R710 B.n244 B.n243 10.6151
R711 B.n244 B.n83 10.6151
R712 B.n248 B.n83 10.6151
R713 B.n249 B.n248 10.6151
R714 B.n477 B.n0 8.11757
R715 B.n477 B.n1 8.11757
R716 B.n395 B.n32 6.5566
R717 B.n383 B.n382 6.5566
R718 B.n206 B.n205 6.5566
R719 B.n219 B.n218 6.5566
R720 B.n32 B.n28 4.05904
R721 B.n382 B.n381 4.05904
R722 B.n205 B.n204 4.05904
R723 B.n220 B.n219 4.05904
R724 VN VN.t0 105.831
R725 VN VN.t1 63.9512
R726 VTAIL.n90 VTAIL.n72 756.745
R727 VTAIL.n18 VTAIL.n0 756.745
R728 VTAIL.n66 VTAIL.n48 756.745
R729 VTAIL.n42 VTAIL.n24 756.745
R730 VTAIL.n81 VTAIL.n80 585
R731 VTAIL.n83 VTAIL.n82 585
R732 VTAIL.n76 VTAIL.n75 585
R733 VTAIL.n89 VTAIL.n88 585
R734 VTAIL.n91 VTAIL.n90 585
R735 VTAIL.n9 VTAIL.n8 585
R736 VTAIL.n11 VTAIL.n10 585
R737 VTAIL.n4 VTAIL.n3 585
R738 VTAIL.n17 VTAIL.n16 585
R739 VTAIL.n19 VTAIL.n18 585
R740 VTAIL.n67 VTAIL.n66 585
R741 VTAIL.n65 VTAIL.n64 585
R742 VTAIL.n52 VTAIL.n51 585
R743 VTAIL.n59 VTAIL.n58 585
R744 VTAIL.n57 VTAIL.n56 585
R745 VTAIL.n43 VTAIL.n42 585
R746 VTAIL.n41 VTAIL.n40 585
R747 VTAIL.n28 VTAIL.n27 585
R748 VTAIL.n35 VTAIL.n34 585
R749 VTAIL.n33 VTAIL.n32 585
R750 VTAIL.n79 VTAIL.t2 328.587
R751 VTAIL.n7 VTAIL.t1 328.587
R752 VTAIL.n55 VTAIL.t0 328.587
R753 VTAIL.n31 VTAIL.t3 328.587
R754 VTAIL.n82 VTAIL.n81 171.744
R755 VTAIL.n82 VTAIL.n75 171.744
R756 VTAIL.n89 VTAIL.n75 171.744
R757 VTAIL.n90 VTAIL.n89 171.744
R758 VTAIL.n10 VTAIL.n9 171.744
R759 VTAIL.n10 VTAIL.n3 171.744
R760 VTAIL.n17 VTAIL.n3 171.744
R761 VTAIL.n18 VTAIL.n17 171.744
R762 VTAIL.n66 VTAIL.n65 171.744
R763 VTAIL.n65 VTAIL.n51 171.744
R764 VTAIL.n58 VTAIL.n51 171.744
R765 VTAIL.n58 VTAIL.n57 171.744
R766 VTAIL.n42 VTAIL.n41 171.744
R767 VTAIL.n41 VTAIL.n27 171.744
R768 VTAIL.n34 VTAIL.n27 171.744
R769 VTAIL.n34 VTAIL.n33 171.744
R770 VTAIL.n81 VTAIL.t2 85.8723
R771 VTAIL.n9 VTAIL.t1 85.8723
R772 VTAIL.n57 VTAIL.t0 85.8723
R773 VTAIL.n33 VTAIL.t3 85.8723
R774 VTAIL.n95 VTAIL.n94 33.7369
R775 VTAIL.n23 VTAIL.n22 33.7369
R776 VTAIL.n71 VTAIL.n70 33.7369
R777 VTAIL.n47 VTAIL.n46 33.7369
R778 VTAIL.n47 VTAIL.n23 23.7634
R779 VTAIL.n95 VTAIL.n71 20.0652
R780 VTAIL.n80 VTAIL.n79 16.3651
R781 VTAIL.n8 VTAIL.n7 16.3651
R782 VTAIL.n56 VTAIL.n55 16.3651
R783 VTAIL.n32 VTAIL.n31 16.3651
R784 VTAIL.n83 VTAIL.n78 12.8005
R785 VTAIL.n11 VTAIL.n6 12.8005
R786 VTAIL.n59 VTAIL.n54 12.8005
R787 VTAIL.n35 VTAIL.n30 12.8005
R788 VTAIL.n84 VTAIL.n76 12.0247
R789 VTAIL.n12 VTAIL.n4 12.0247
R790 VTAIL.n60 VTAIL.n52 12.0247
R791 VTAIL.n36 VTAIL.n28 12.0247
R792 VTAIL.n88 VTAIL.n87 11.249
R793 VTAIL.n16 VTAIL.n15 11.249
R794 VTAIL.n64 VTAIL.n63 11.249
R795 VTAIL.n40 VTAIL.n39 11.249
R796 VTAIL.n91 VTAIL.n74 10.4732
R797 VTAIL.n19 VTAIL.n2 10.4732
R798 VTAIL.n67 VTAIL.n50 10.4732
R799 VTAIL.n43 VTAIL.n26 10.4732
R800 VTAIL.n92 VTAIL.n72 9.69747
R801 VTAIL.n20 VTAIL.n0 9.69747
R802 VTAIL.n68 VTAIL.n48 9.69747
R803 VTAIL.n44 VTAIL.n24 9.69747
R804 VTAIL.n94 VTAIL.n93 9.45567
R805 VTAIL.n22 VTAIL.n21 9.45567
R806 VTAIL.n70 VTAIL.n69 9.45567
R807 VTAIL.n46 VTAIL.n45 9.45567
R808 VTAIL.n93 VTAIL.n92 9.3005
R809 VTAIL.n74 VTAIL.n73 9.3005
R810 VTAIL.n87 VTAIL.n86 9.3005
R811 VTAIL.n85 VTAIL.n84 9.3005
R812 VTAIL.n78 VTAIL.n77 9.3005
R813 VTAIL.n21 VTAIL.n20 9.3005
R814 VTAIL.n2 VTAIL.n1 9.3005
R815 VTAIL.n15 VTAIL.n14 9.3005
R816 VTAIL.n13 VTAIL.n12 9.3005
R817 VTAIL.n6 VTAIL.n5 9.3005
R818 VTAIL.n69 VTAIL.n68 9.3005
R819 VTAIL.n50 VTAIL.n49 9.3005
R820 VTAIL.n63 VTAIL.n62 9.3005
R821 VTAIL.n61 VTAIL.n60 9.3005
R822 VTAIL.n54 VTAIL.n53 9.3005
R823 VTAIL.n45 VTAIL.n44 9.3005
R824 VTAIL.n26 VTAIL.n25 9.3005
R825 VTAIL.n39 VTAIL.n38 9.3005
R826 VTAIL.n37 VTAIL.n36 9.3005
R827 VTAIL.n30 VTAIL.n29 9.3005
R828 VTAIL.n94 VTAIL.n72 4.26717
R829 VTAIL.n22 VTAIL.n0 4.26717
R830 VTAIL.n70 VTAIL.n48 4.26717
R831 VTAIL.n46 VTAIL.n24 4.26717
R832 VTAIL.n79 VTAIL.n77 3.73474
R833 VTAIL.n7 VTAIL.n5 3.73474
R834 VTAIL.n55 VTAIL.n53 3.73474
R835 VTAIL.n31 VTAIL.n29 3.73474
R836 VTAIL.n92 VTAIL.n91 3.49141
R837 VTAIL.n20 VTAIL.n19 3.49141
R838 VTAIL.n68 VTAIL.n67 3.49141
R839 VTAIL.n44 VTAIL.n43 3.49141
R840 VTAIL.n88 VTAIL.n74 2.71565
R841 VTAIL.n16 VTAIL.n2 2.71565
R842 VTAIL.n64 VTAIL.n50 2.71565
R843 VTAIL.n40 VTAIL.n26 2.71565
R844 VTAIL.n71 VTAIL.n47 2.31947
R845 VTAIL.n87 VTAIL.n76 1.93989
R846 VTAIL.n15 VTAIL.n4 1.93989
R847 VTAIL.n63 VTAIL.n52 1.93989
R848 VTAIL.n39 VTAIL.n28 1.93989
R849 VTAIL VTAIL.n23 1.45309
R850 VTAIL.n84 VTAIL.n83 1.16414
R851 VTAIL.n12 VTAIL.n11 1.16414
R852 VTAIL.n60 VTAIL.n59 1.16414
R853 VTAIL.n36 VTAIL.n35 1.16414
R854 VTAIL VTAIL.n95 0.866879
R855 VTAIL.n80 VTAIL.n78 0.388379
R856 VTAIL.n8 VTAIL.n6 0.388379
R857 VTAIL.n56 VTAIL.n54 0.388379
R858 VTAIL.n32 VTAIL.n30 0.388379
R859 VTAIL.n85 VTAIL.n77 0.155672
R860 VTAIL.n86 VTAIL.n85 0.155672
R861 VTAIL.n86 VTAIL.n73 0.155672
R862 VTAIL.n93 VTAIL.n73 0.155672
R863 VTAIL.n13 VTAIL.n5 0.155672
R864 VTAIL.n14 VTAIL.n13 0.155672
R865 VTAIL.n14 VTAIL.n1 0.155672
R866 VTAIL.n21 VTAIL.n1 0.155672
R867 VTAIL.n69 VTAIL.n49 0.155672
R868 VTAIL.n62 VTAIL.n49 0.155672
R869 VTAIL.n62 VTAIL.n61 0.155672
R870 VTAIL.n61 VTAIL.n53 0.155672
R871 VTAIL.n45 VTAIL.n25 0.155672
R872 VTAIL.n38 VTAIL.n25 0.155672
R873 VTAIL.n38 VTAIL.n37 0.155672
R874 VTAIL.n37 VTAIL.n29 0.155672
R875 VDD2.n41 VDD2.n23 756.745
R876 VDD2.n18 VDD2.n0 756.745
R877 VDD2.n42 VDD2.n41 585
R878 VDD2.n40 VDD2.n39 585
R879 VDD2.n27 VDD2.n26 585
R880 VDD2.n34 VDD2.n33 585
R881 VDD2.n32 VDD2.n31 585
R882 VDD2.n9 VDD2.n8 585
R883 VDD2.n11 VDD2.n10 585
R884 VDD2.n4 VDD2.n3 585
R885 VDD2.n17 VDD2.n16 585
R886 VDD2.n19 VDD2.n18 585
R887 VDD2.n30 VDD2.t1 328.587
R888 VDD2.n7 VDD2.t0 328.587
R889 VDD2.n41 VDD2.n40 171.744
R890 VDD2.n40 VDD2.n26 171.744
R891 VDD2.n33 VDD2.n26 171.744
R892 VDD2.n33 VDD2.n32 171.744
R893 VDD2.n10 VDD2.n9 171.744
R894 VDD2.n10 VDD2.n3 171.744
R895 VDD2.n17 VDD2.n3 171.744
R896 VDD2.n18 VDD2.n17 171.744
R897 VDD2.n32 VDD2.t1 85.8723
R898 VDD2.n9 VDD2.t0 85.8723
R899 VDD2.n46 VDD2.n22 85.4716
R900 VDD2.n46 VDD2.n45 50.4157
R901 VDD2.n31 VDD2.n30 16.3651
R902 VDD2.n8 VDD2.n7 16.3651
R903 VDD2.n34 VDD2.n29 12.8005
R904 VDD2.n11 VDD2.n6 12.8005
R905 VDD2.n35 VDD2.n27 12.0247
R906 VDD2.n12 VDD2.n4 12.0247
R907 VDD2.n39 VDD2.n38 11.249
R908 VDD2.n16 VDD2.n15 11.249
R909 VDD2.n42 VDD2.n25 10.4732
R910 VDD2.n19 VDD2.n2 10.4732
R911 VDD2.n43 VDD2.n23 9.69747
R912 VDD2.n20 VDD2.n0 9.69747
R913 VDD2.n45 VDD2.n44 9.45567
R914 VDD2.n22 VDD2.n21 9.45567
R915 VDD2.n44 VDD2.n43 9.3005
R916 VDD2.n25 VDD2.n24 9.3005
R917 VDD2.n38 VDD2.n37 9.3005
R918 VDD2.n36 VDD2.n35 9.3005
R919 VDD2.n29 VDD2.n28 9.3005
R920 VDD2.n21 VDD2.n20 9.3005
R921 VDD2.n2 VDD2.n1 9.3005
R922 VDD2.n15 VDD2.n14 9.3005
R923 VDD2.n13 VDD2.n12 9.3005
R924 VDD2.n6 VDD2.n5 9.3005
R925 VDD2.n45 VDD2.n23 4.26717
R926 VDD2.n22 VDD2.n0 4.26717
R927 VDD2.n30 VDD2.n28 3.73474
R928 VDD2.n7 VDD2.n5 3.73474
R929 VDD2.n43 VDD2.n42 3.49141
R930 VDD2.n20 VDD2.n19 3.49141
R931 VDD2.n39 VDD2.n25 2.71565
R932 VDD2.n16 VDD2.n2 2.71565
R933 VDD2.n38 VDD2.n27 1.93989
R934 VDD2.n15 VDD2.n4 1.93989
R935 VDD2.n35 VDD2.n34 1.16414
R936 VDD2.n12 VDD2.n11 1.16414
R937 VDD2 VDD2.n46 0.983259
R938 VDD2.n31 VDD2.n29 0.388379
R939 VDD2.n8 VDD2.n6 0.388379
R940 VDD2.n44 VDD2.n24 0.155672
R941 VDD2.n37 VDD2.n24 0.155672
R942 VDD2.n37 VDD2.n36 0.155672
R943 VDD2.n36 VDD2.n28 0.155672
R944 VDD2.n13 VDD2.n5 0.155672
R945 VDD2.n14 VDD2.n13 0.155672
R946 VDD2.n14 VDD2.n1 0.155672
R947 VDD2.n21 VDD2.n1 0.155672
R948 VP.n0 VP.t1 106.017
R949 VP.n0 VP.t0 63.3305
R950 VP VP.n0 0.62124
R951 VDD1.n18 VDD1.n0 756.745
R952 VDD1.n41 VDD1.n23 756.745
R953 VDD1.n19 VDD1.n18 585
R954 VDD1.n17 VDD1.n16 585
R955 VDD1.n4 VDD1.n3 585
R956 VDD1.n11 VDD1.n10 585
R957 VDD1.n9 VDD1.n8 585
R958 VDD1.n32 VDD1.n31 585
R959 VDD1.n34 VDD1.n33 585
R960 VDD1.n27 VDD1.n26 585
R961 VDD1.n40 VDD1.n39 585
R962 VDD1.n42 VDD1.n41 585
R963 VDD1.n7 VDD1.t0 328.587
R964 VDD1.n30 VDD1.t1 328.587
R965 VDD1.n18 VDD1.n17 171.744
R966 VDD1.n17 VDD1.n3 171.744
R967 VDD1.n10 VDD1.n3 171.744
R968 VDD1.n10 VDD1.n9 171.744
R969 VDD1.n33 VDD1.n32 171.744
R970 VDD1.n33 VDD1.n26 171.744
R971 VDD1.n40 VDD1.n26 171.744
R972 VDD1.n41 VDD1.n40 171.744
R973 VDD1 VDD1.n45 86.921
R974 VDD1.n9 VDD1.t0 85.8723
R975 VDD1.n32 VDD1.t1 85.8723
R976 VDD1 VDD1.n22 51.3984
R977 VDD1.n8 VDD1.n7 16.3651
R978 VDD1.n31 VDD1.n30 16.3651
R979 VDD1.n11 VDD1.n6 12.8005
R980 VDD1.n34 VDD1.n29 12.8005
R981 VDD1.n12 VDD1.n4 12.0247
R982 VDD1.n35 VDD1.n27 12.0247
R983 VDD1.n16 VDD1.n15 11.249
R984 VDD1.n39 VDD1.n38 11.249
R985 VDD1.n19 VDD1.n2 10.4732
R986 VDD1.n42 VDD1.n25 10.4732
R987 VDD1.n20 VDD1.n0 9.69747
R988 VDD1.n43 VDD1.n23 9.69747
R989 VDD1.n22 VDD1.n21 9.45567
R990 VDD1.n45 VDD1.n44 9.45567
R991 VDD1.n21 VDD1.n20 9.3005
R992 VDD1.n2 VDD1.n1 9.3005
R993 VDD1.n15 VDD1.n14 9.3005
R994 VDD1.n13 VDD1.n12 9.3005
R995 VDD1.n6 VDD1.n5 9.3005
R996 VDD1.n44 VDD1.n43 9.3005
R997 VDD1.n25 VDD1.n24 9.3005
R998 VDD1.n38 VDD1.n37 9.3005
R999 VDD1.n36 VDD1.n35 9.3005
R1000 VDD1.n29 VDD1.n28 9.3005
R1001 VDD1.n22 VDD1.n0 4.26717
R1002 VDD1.n45 VDD1.n23 4.26717
R1003 VDD1.n7 VDD1.n5 3.73474
R1004 VDD1.n30 VDD1.n28 3.73474
R1005 VDD1.n20 VDD1.n19 3.49141
R1006 VDD1.n43 VDD1.n42 3.49141
R1007 VDD1.n16 VDD1.n2 2.71565
R1008 VDD1.n39 VDD1.n25 2.71565
R1009 VDD1.n15 VDD1.n4 1.93989
R1010 VDD1.n38 VDD1.n27 1.93989
R1011 VDD1.n12 VDD1.n11 1.16414
R1012 VDD1.n35 VDD1.n34 1.16414
R1013 VDD1.n8 VDD1.n6 0.388379
R1014 VDD1.n31 VDD1.n29 0.388379
R1015 VDD1.n21 VDD1.n1 0.155672
R1016 VDD1.n14 VDD1.n1 0.155672
R1017 VDD1.n14 VDD1.n13 0.155672
R1018 VDD1.n13 VDD1.n5 0.155672
R1019 VDD1.n36 VDD1.n28 0.155672
R1020 VDD1.n37 VDD1.n36 0.155672
R1021 VDD1.n37 VDD1.n24 0.155672
R1022 VDD1.n44 VDD1.n24 0.155672
C0 B VTAIL 2.33636f
C1 VTAIL VN 1.53997f
C2 VDD1 VDD2 0.827739f
C3 w_n2686_n1896# VTAIL 1.78415f
C4 B VDD1 1.28758f
C5 B VDD2 1.33007f
C6 VDD1 VN 0.152998f
C7 VDD2 VN 1.29584f
C8 B VN 1.19459f
C9 VDD1 w_n2686_n1896# 1.43035f
C10 w_n2686_n1896# VDD2 1.47265f
C11 B w_n2686_n1896# 8.2368f
C12 w_n2686_n1896# VN 3.69289f
C13 VTAIL VP 1.55438f
C14 VDD1 VP 1.53572f
C15 VDD2 VP 0.394172f
C16 B VP 1.76728f
C17 VP VN 4.72691f
C18 w_n2686_n1896# VP 4.03787f
C19 VDD1 VTAIL 3.53079f
C20 VTAIL VDD2 3.59266f
C21 VDD2 VSUBS 0.749359f
C22 VDD1 VSUBS 2.668975f
C23 VTAIL VSUBS 0.540864f
C24 VN VSUBS 6.00562f
C25 VP VSUBS 1.668217f
C26 B VSUBS 4.061018f
C27 w_n2686_n1896# VSUBS 63.916103f
C28 VDD1.n0 VSUBS 0.01686f
C29 VDD1.n1 VSUBS 0.015403f
C30 VDD1.n2 VSUBS 0.008277f
C31 VDD1.n3 VSUBS 0.019563f
C32 VDD1.n4 VSUBS 0.008764f
C33 VDD1.n5 VSUBS 0.256933f
C34 VDD1.n6 VSUBS 0.008277f
C35 VDD1.t0 VSUBS 0.042675f
C36 VDD1.n7 VSUBS 0.062519f
C37 VDD1.n8 VSUBS 0.012394f
C38 VDD1.n9 VSUBS 0.014673f
C39 VDD1.n10 VSUBS 0.019563f
C40 VDD1.n11 VSUBS 0.008764f
C41 VDD1.n12 VSUBS 0.008277f
C42 VDD1.n13 VSUBS 0.015403f
C43 VDD1.n14 VSUBS 0.015403f
C44 VDD1.n15 VSUBS 0.008277f
C45 VDD1.n16 VSUBS 0.008764f
C46 VDD1.n17 VSUBS 0.019563f
C47 VDD1.n18 VSUBS 0.047141f
C48 VDD1.n19 VSUBS 0.008764f
C49 VDD1.n20 VSUBS 0.008277f
C50 VDD1.n21 VSUBS 0.037286f
C51 VDD1.n22 VSUBS 0.035889f
C52 VDD1.n23 VSUBS 0.01686f
C53 VDD1.n24 VSUBS 0.015403f
C54 VDD1.n25 VSUBS 0.008277f
C55 VDD1.n26 VSUBS 0.019563f
C56 VDD1.n27 VSUBS 0.008764f
C57 VDD1.n28 VSUBS 0.256933f
C58 VDD1.n29 VSUBS 0.008277f
C59 VDD1.t1 VSUBS 0.042675f
C60 VDD1.n30 VSUBS 0.062519f
C61 VDD1.n31 VSUBS 0.012394f
C62 VDD1.n32 VSUBS 0.014673f
C63 VDD1.n33 VSUBS 0.019563f
C64 VDD1.n34 VSUBS 0.008764f
C65 VDD1.n35 VSUBS 0.008277f
C66 VDD1.n36 VSUBS 0.015403f
C67 VDD1.n37 VSUBS 0.015403f
C68 VDD1.n38 VSUBS 0.008277f
C69 VDD1.n39 VSUBS 0.008764f
C70 VDD1.n40 VSUBS 0.019563f
C71 VDD1.n41 VSUBS 0.047141f
C72 VDD1.n42 VSUBS 0.008764f
C73 VDD1.n43 VSUBS 0.008277f
C74 VDD1.n44 VSUBS 0.037286f
C75 VDD1.n45 VSUBS 0.379859f
C76 VP.t1 VSUBS 3.02485f
C77 VP.t0 VSUBS 2.1414f
C78 VP.n0 VSUBS 3.38101f
C79 VDD2.n0 VSUBS 0.017628f
C80 VDD2.n1 VSUBS 0.016105f
C81 VDD2.n2 VSUBS 0.008654f
C82 VDD2.n3 VSUBS 0.020455f
C83 VDD2.n4 VSUBS 0.009163f
C84 VDD2.n5 VSUBS 0.268641f
C85 VDD2.n6 VSUBS 0.008654f
C86 VDD2.t0 VSUBS 0.04462f
C87 VDD2.n7 VSUBS 0.065368f
C88 VDD2.n8 VSUBS 0.012958f
C89 VDD2.n9 VSUBS 0.015341f
C90 VDD2.n10 VSUBS 0.020455f
C91 VDD2.n11 VSUBS 0.009163f
C92 VDD2.n12 VSUBS 0.008654f
C93 VDD2.n13 VSUBS 0.016105f
C94 VDD2.n14 VSUBS 0.016105f
C95 VDD2.n15 VSUBS 0.008654f
C96 VDD2.n16 VSUBS 0.009163f
C97 VDD2.n17 VSUBS 0.020455f
C98 VDD2.n18 VSUBS 0.049289f
C99 VDD2.n19 VSUBS 0.009163f
C100 VDD2.n20 VSUBS 0.008654f
C101 VDD2.n21 VSUBS 0.038985f
C102 VDD2.n22 VSUBS 0.363426f
C103 VDD2.n23 VSUBS 0.017628f
C104 VDD2.n24 VSUBS 0.016105f
C105 VDD2.n25 VSUBS 0.008654f
C106 VDD2.n26 VSUBS 0.020455f
C107 VDD2.n27 VSUBS 0.009163f
C108 VDD2.n28 VSUBS 0.268641f
C109 VDD2.n29 VSUBS 0.008654f
C110 VDD2.t1 VSUBS 0.04462f
C111 VDD2.n30 VSUBS 0.065368f
C112 VDD2.n31 VSUBS 0.012958f
C113 VDD2.n32 VSUBS 0.015341f
C114 VDD2.n33 VSUBS 0.020455f
C115 VDD2.n34 VSUBS 0.009163f
C116 VDD2.n35 VSUBS 0.008654f
C117 VDD2.n36 VSUBS 0.016105f
C118 VDD2.n37 VSUBS 0.016105f
C119 VDD2.n38 VSUBS 0.008654f
C120 VDD2.n39 VSUBS 0.009163f
C121 VDD2.n40 VSUBS 0.020455f
C122 VDD2.n41 VSUBS 0.049289f
C123 VDD2.n42 VSUBS 0.009163f
C124 VDD2.n43 VSUBS 0.008654f
C125 VDD2.n44 VSUBS 0.038985f
C126 VDD2.n45 VSUBS 0.035937f
C127 VDD2.n46 VSUBS 1.64837f
C128 VTAIL.n0 VSUBS 0.026277f
C129 VTAIL.n1 VSUBS 0.024006f
C130 VTAIL.n2 VSUBS 0.012899f
C131 VTAIL.n3 VSUBS 0.03049f
C132 VTAIL.n4 VSUBS 0.013658f
C133 VTAIL.n5 VSUBS 0.400434f
C134 VTAIL.n6 VSUBS 0.012899f
C135 VTAIL.t1 VSUBS 0.06651f
C136 VTAIL.n7 VSUBS 0.097438f
C137 VTAIL.n8 VSUBS 0.019316f
C138 VTAIL.n9 VSUBS 0.022867f
C139 VTAIL.n10 VSUBS 0.03049f
C140 VTAIL.n11 VSUBS 0.013658f
C141 VTAIL.n12 VSUBS 0.012899f
C142 VTAIL.n13 VSUBS 0.024006f
C143 VTAIL.n14 VSUBS 0.024006f
C144 VTAIL.n15 VSUBS 0.012899f
C145 VTAIL.n16 VSUBS 0.013658f
C146 VTAIL.n17 VSUBS 0.03049f
C147 VTAIL.n18 VSUBS 0.073471f
C148 VTAIL.n19 VSUBS 0.013658f
C149 VTAIL.n20 VSUBS 0.012899f
C150 VTAIL.n21 VSUBS 0.058111f
C151 VTAIL.n22 VSUBS 0.037012f
C152 VTAIL.n23 VSUBS 1.34197f
C153 VTAIL.n24 VSUBS 0.026277f
C154 VTAIL.n25 VSUBS 0.024006f
C155 VTAIL.n26 VSUBS 0.012899f
C156 VTAIL.n27 VSUBS 0.03049f
C157 VTAIL.n28 VSUBS 0.013658f
C158 VTAIL.n29 VSUBS 0.400434f
C159 VTAIL.n30 VSUBS 0.012899f
C160 VTAIL.t3 VSUBS 0.06651f
C161 VTAIL.n31 VSUBS 0.097438f
C162 VTAIL.n32 VSUBS 0.019316f
C163 VTAIL.n33 VSUBS 0.022867f
C164 VTAIL.n34 VSUBS 0.03049f
C165 VTAIL.n35 VSUBS 0.013658f
C166 VTAIL.n36 VSUBS 0.012899f
C167 VTAIL.n37 VSUBS 0.024006f
C168 VTAIL.n38 VSUBS 0.024006f
C169 VTAIL.n39 VSUBS 0.012899f
C170 VTAIL.n40 VSUBS 0.013658f
C171 VTAIL.n41 VSUBS 0.03049f
C172 VTAIL.n42 VSUBS 0.073471f
C173 VTAIL.n43 VSUBS 0.013658f
C174 VTAIL.n44 VSUBS 0.012899f
C175 VTAIL.n45 VSUBS 0.058111f
C176 VTAIL.n46 VSUBS 0.037012f
C177 VTAIL.n47 VSUBS 1.40898f
C178 VTAIL.n48 VSUBS 0.026277f
C179 VTAIL.n49 VSUBS 0.024006f
C180 VTAIL.n50 VSUBS 0.012899f
C181 VTAIL.n51 VSUBS 0.03049f
C182 VTAIL.n52 VSUBS 0.013658f
C183 VTAIL.n53 VSUBS 0.400434f
C184 VTAIL.n54 VSUBS 0.012899f
C185 VTAIL.t0 VSUBS 0.06651f
C186 VTAIL.n55 VSUBS 0.097438f
C187 VTAIL.n56 VSUBS 0.019316f
C188 VTAIL.n57 VSUBS 0.022867f
C189 VTAIL.n58 VSUBS 0.03049f
C190 VTAIL.n59 VSUBS 0.013658f
C191 VTAIL.n60 VSUBS 0.012899f
C192 VTAIL.n61 VSUBS 0.024006f
C193 VTAIL.n62 VSUBS 0.024006f
C194 VTAIL.n63 VSUBS 0.012899f
C195 VTAIL.n64 VSUBS 0.013658f
C196 VTAIL.n65 VSUBS 0.03049f
C197 VTAIL.n66 VSUBS 0.073471f
C198 VTAIL.n67 VSUBS 0.013658f
C199 VTAIL.n68 VSUBS 0.012899f
C200 VTAIL.n69 VSUBS 0.058111f
C201 VTAIL.n70 VSUBS 0.037012f
C202 VTAIL.n71 VSUBS 1.12292f
C203 VTAIL.n72 VSUBS 0.026277f
C204 VTAIL.n73 VSUBS 0.024006f
C205 VTAIL.n74 VSUBS 0.012899f
C206 VTAIL.n75 VSUBS 0.03049f
C207 VTAIL.n76 VSUBS 0.013658f
C208 VTAIL.n77 VSUBS 0.400434f
C209 VTAIL.n78 VSUBS 0.012899f
C210 VTAIL.t2 VSUBS 0.06651f
C211 VTAIL.n79 VSUBS 0.097438f
C212 VTAIL.n80 VSUBS 0.019316f
C213 VTAIL.n81 VSUBS 0.022867f
C214 VTAIL.n82 VSUBS 0.03049f
C215 VTAIL.n83 VSUBS 0.013658f
C216 VTAIL.n84 VSUBS 0.012899f
C217 VTAIL.n85 VSUBS 0.024006f
C218 VTAIL.n86 VSUBS 0.024006f
C219 VTAIL.n87 VSUBS 0.012899f
C220 VTAIL.n88 VSUBS 0.013658f
C221 VTAIL.n89 VSUBS 0.03049f
C222 VTAIL.n90 VSUBS 0.073471f
C223 VTAIL.n91 VSUBS 0.013658f
C224 VTAIL.n92 VSUBS 0.012899f
C225 VTAIL.n93 VSUBS 0.058111f
C226 VTAIL.n94 VSUBS 0.037012f
C227 VTAIL.n95 VSUBS 1.01056f
C228 VN.t1 VSUBS 2.06264f
C229 VN.t0 VSUBS 2.90283f
C230 B.n0 VSUBS 0.007264f
C231 B.n1 VSUBS 0.007264f
C232 B.n2 VSUBS 0.010743f
C233 B.n3 VSUBS 0.008232f
C234 B.n4 VSUBS 0.008232f
C235 B.n5 VSUBS 0.008232f
C236 B.n6 VSUBS 0.008232f
C237 B.n7 VSUBS 0.008232f
C238 B.n8 VSUBS 0.008232f
C239 B.n9 VSUBS 0.008232f
C240 B.n10 VSUBS 0.008232f
C241 B.n11 VSUBS 0.008232f
C242 B.n12 VSUBS 0.008232f
C243 B.n13 VSUBS 0.008232f
C244 B.n14 VSUBS 0.008232f
C245 B.n15 VSUBS 0.008232f
C246 B.n16 VSUBS 0.008232f
C247 B.n17 VSUBS 0.008232f
C248 B.n18 VSUBS 0.019485f
C249 B.n19 VSUBS 0.008232f
C250 B.n20 VSUBS 0.008232f
C251 B.n21 VSUBS 0.008232f
C252 B.n22 VSUBS 0.008232f
C253 B.n23 VSUBS 0.008232f
C254 B.n24 VSUBS 0.008232f
C255 B.n25 VSUBS 0.008232f
C256 B.n26 VSUBS 0.008232f
C257 B.n27 VSUBS 0.008232f
C258 B.n28 VSUBS 0.00569f
C259 B.n29 VSUBS 0.008232f
C260 B.t10 VSUBS 0.079096f
C261 B.t11 VSUBS 0.116395f
C262 B.t9 VSUBS 1.04904f
C263 B.n30 VSUBS 0.194195f
C264 B.n31 VSUBS 0.158927f
C265 B.n32 VSUBS 0.019073f
C266 B.n33 VSUBS 0.008232f
C267 B.n34 VSUBS 0.008232f
C268 B.n35 VSUBS 0.008232f
C269 B.n36 VSUBS 0.008232f
C270 B.t7 VSUBS 0.079098f
C271 B.t8 VSUBS 0.116396f
C272 B.t6 VSUBS 1.04904f
C273 B.n37 VSUBS 0.194194f
C274 B.n38 VSUBS 0.158925f
C275 B.n39 VSUBS 0.008232f
C276 B.n40 VSUBS 0.008232f
C277 B.n41 VSUBS 0.008232f
C278 B.n42 VSUBS 0.008232f
C279 B.n43 VSUBS 0.008232f
C280 B.n44 VSUBS 0.008232f
C281 B.n45 VSUBS 0.008232f
C282 B.n46 VSUBS 0.008232f
C283 B.n47 VSUBS 0.008232f
C284 B.n48 VSUBS 0.019485f
C285 B.n49 VSUBS 0.008232f
C286 B.n50 VSUBS 0.008232f
C287 B.n51 VSUBS 0.008232f
C288 B.n52 VSUBS 0.008232f
C289 B.n53 VSUBS 0.008232f
C290 B.n54 VSUBS 0.008232f
C291 B.n55 VSUBS 0.008232f
C292 B.n56 VSUBS 0.008232f
C293 B.n57 VSUBS 0.008232f
C294 B.n58 VSUBS 0.008232f
C295 B.n59 VSUBS 0.008232f
C296 B.n60 VSUBS 0.008232f
C297 B.n61 VSUBS 0.008232f
C298 B.n62 VSUBS 0.008232f
C299 B.n63 VSUBS 0.008232f
C300 B.n64 VSUBS 0.008232f
C301 B.n65 VSUBS 0.008232f
C302 B.n66 VSUBS 0.008232f
C303 B.n67 VSUBS 0.008232f
C304 B.n68 VSUBS 0.008232f
C305 B.n69 VSUBS 0.008232f
C306 B.n70 VSUBS 0.008232f
C307 B.n71 VSUBS 0.008232f
C308 B.n72 VSUBS 0.008232f
C309 B.n73 VSUBS 0.008232f
C310 B.n74 VSUBS 0.008232f
C311 B.n75 VSUBS 0.008232f
C312 B.n76 VSUBS 0.008232f
C313 B.n77 VSUBS 0.008232f
C314 B.n78 VSUBS 0.008232f
C315 B.n79 VSUBS 0.008232f
C316 B.n80 VSUBS 0.008232f
C317 B.n81 VSUBS 0.008232f
C318 B.n82 VSUBS 0.019739f
C319 B.n83 VSUBS 0.008232f
C320 B.n84 VSUBS 0.008232f
C321 B.n85 VSUBS 0.008232f
C322 B.n86 VSUBS 0.008232f
C323 B.n87 VSUBS 0.008232f
C324 B.n88 VSUBS 0.008232f
C325 B.n89 VSUBS 0.008232f
C326 B.n90 VSUBS 0.008232f
C327 B.n91 VSUBS 0.008232f
C328 B.n92 VSUBS 0.008232f
C329 B.t5 VSUBS 0.079098f
C330 B.t4 VSUBS 0.116396f
C331 B.t3 VSUBS 1.04904f
C332 B.n93 VSUBS 0.194194f
C333 B.n94 VSUBS 0.158925f
C334 B.n95 VSUBS 0.008232f
C335 B.n96 VSUBS 0.008232f
C336 B.n97 VSUBS 0.008232f
C337 B.n98 VSUBS 0.008232f
C338 B.t2 VSUBS 0.079096f
C339 B.t1 VSUBS 0.116395f
C340 B.t0 VSUBS 1.04904f
C341 B.n99 VSUBS 0.194195f
C342 B.n100 VSUBS 0.158927f
C343 B.n101 VSUBS 0.008232f
C344 B.n102 VSUBS 0.008232f
C345 B.n103 VSUBS 0.008232f
C346 B.n104 VSUBS 0.008232f
C347 B.n105 VSUBS 0.008232f
C348 B.n106 VSUBS 0.008232f
C349 B.n107 VSUBS 0.008232f
C350 B.n108 VSUBS 0.008232f
C351 B.n109 VSUBS 0.008232f
C352 B.n110 VSUBS 0.019739f
C353 B.n111 VSUBS 0.008232f
C354 B.n112 VSUBS 0.008232f
C355 B.n113 VSUBS 0.008232f
C356 B.n114 VSUBS 0.008232f
C357 B.n115 VSUBS 0.008232f
C358 B.n116 VSUBS 0.008232f
C359 B.n117 VSUBS 0.008232f
C360 B.n118 VSUBS 0.008232f
C361 B.n119 VSUBS 0.008232f
C362 B.n120 VSUBS 0.008232f
C363 B.n121 VSUBS 0.008232f
C364 B.n122 VSUBS 0.008232f
C365 B.n123 VSUBS 0.008232f
C366 B.n124 VSUBS 0.008232f
C367 B.n125 VSUBS 0.008232f
C368 B.n126 VSUBS 0.008232f
C369 B.n127 VSUBS 0.008232f
C370 B.n128 VSUBS 0.008232f
C371 B.n129 VSUBS 0.008232f
C372 B.n130 VSUBS 0.008232f
C373 B.n131 VSUBS 0.008232f
C374 B.n132 VSUBS 0.008232f
C375 B.n133 VSUBS 0.008232f
C376 B.n134 VSUBS 0.008232f
C377 B.n135 VSUBS 0.008232f
C378 B.n136 VSUBS 0.008232f
C379 B.n137 VSUBS 0.008232f
C380 B.n138 VSUBS 0.008232f
C381 B.n139 VSUBS 0.008232f
C382 B.n140 VSUBS 0.008232f
C383 B.n141 VSUBS 0.008232f
C384 B.n142 VSUBS 0.008232f
C385 B.n143 VSUBS 0.008232f
C386 B.n144 VSUBS 0.008232f
C387 B.n145 VSUBS 0.008232f
C388 B.n146 VSUBS 0.008232f
C389 B.n147 VSUBS 0.008232f
C390 B.n148 VSUBS 0.008232f
C391 B.n149 VSUBS 0.008232f
C392 B.n150 VSUBS 0.008232f
C393 B.n151 VSUBS 0.008232f
C394 B.n152 VSUBS 0.008232f
C395 B.n153 VSUBS 0.008232f
C396 B.n154 VSUBS 0.008232f
C397 B.n155 VSUBS 0.008232f
C398 B.n156 VSUBS 0.008232f
C399 B.n157 VSUBS 0.008232f
C400 B.n158 VSUBS 0.008232f
C401 B.n159 VSUBS 0.008232f
C402 B.n160 VSUBS 0.008232f
C403 B.n161 VSUBS 0.008232f
C404 B.n162 VSUBS 0.008232f
C405 B.n163 VSUBS 0.008232f
C406 B.n164 VSUBS 0.008232f
C407 B.n165 VSUBS 0.008232f
C408 B.n166 VSUBS 0.008232f
C409 B.n167 VSUBS 0.008232f
C410 B.n168 VSUBS 0.008232f
C411 B.n169 VSUBS 0.008232f
C412 B.n170 VSUBS 0.008232f
C413 B.n171 VSUBS 0.008232f
C414 B.n172 VSUBS 0.008232f
C415 B.n173 VSUBS 0.019485f
C416 B.n174 VSUBS 0.019485f
C417 B.n175 VSUBS 0.019739f
C418 B.n176 VSUBS 0.008232f
C419 B.n177 VSUBS 0.008232f
C420 B.n178 VSUBS 0.008232f
C421 B.n179 VSUBS 0.008232f
C422 B.n180 VSUBS 0.008232f
C423 B.n181 VSUBS 0.008232f
C424 B.n182 VSUBS 0.008232f
C425 B.n183 VSUBS 0.008232f
C426 B.n184 VSUBS 0.008232f
C427 B.n185 VSUBS 0.008232f
C428 B.n186 VSUBS 0.008232f
C429 B.n187 VSUBS 0.008232f
C430 B.n188 VSUBS 0.008232f
C431 B.n189 VSUBS 0.008232f
C432 B.n190 VSUBS 0.008232f
C433 B.n191 VSUBS 0.008232f
C434 B.n192 VSUBS 0.008232f
C435 B.n193 VSUBS 0.008232f
C436 B.n194 VSUBS 0.008232f
C437 B.n195 VSUBS 0.008232f
C438 B.n196 VSUBS 0.008232f
C439 B.n197 VSUBS 0.008232f
C440 B.n198 VSUBS 0.008232f
C441 B.n199 VSUBS 0.008232f
C442 B.n200 VSUBS 0.008232f
C443 B.n201 VSUBS 0.008232f
C444 B.n202 VSUBS 0.008232f
C445 B.n203 VSUBS 0.008232f
C446 B.n204 VSUBS 0.00569f
C447 B.n205 VSUBS 0.019073f
C448 B.n206 VSUBS 0.006659f
C449 B.n207 VSUBS 0.008232f
C450 B.n208 VSUBS 0.008232f
C451 B.n209 VSUBS 0.008232f
C452 B.n210 VSUBS 0.008232f
C453 B.n211 VSUBS 0.008232f
C454 B.n212 VSUBS 0.008232f
C455 B.n213 VSUBS 0.008232f
C456 B.n214 VSUBS 0.008232f
C457 B.n215 VSUBS 0.008232f
C458 B.n216 VSUBS 0.008232f
C459 B.n217 VSUBS 0.008232f
C460 B.n218 VSUBS 0.006659f
C461 B.n219 VSUBS 0.019073f
C462 B.n220 VSUBS 0.00569f
C463 B.n221 VSUBS 0.008232f
C464 B.n222 VSUBS 0.008232f
C465 B.n223 VSUBS 0.008232f
C466 B.n224 VSUBS 0.008232f
C467 B.n225 VSUBS 0.008232f
C468 B.n226 VSUBS 0.008232f
C469 B.n227 VSUBS 0.008232f
C470 B.n228 VSUBS 0.008232f
C471 B.n229 VSUBS 0.008232f
C472 B.n230 VSUBS 0.008232f
C473 B.n231 VSUBS 0.008232f
C474 B.n232 VSUBS 0.008232f
C475 B.n233 VSUBS 0.008232f
C476 B.n234 VSUBS 0.008232f
C477 B.n235 VSUBS 0.008232f
C478 B.n236 VSUBS 0.008232f
C479 B.n237 VSUBS 0.008232f
C480 B.n238 VSUBS 0.008232f
C481 B.n239 VSUBS 0.008232f
C482 B.n240 VSUBS 0.008232f
C483 B.n241 VSUBS 0.008232f
C484 B.n242 VSUBS 0.008232f
C485 B.n243 VSUBS 0.008232f
C486 B.n244 VSUBS 0.008232f
C487 B.n245 VSUBS 0.008232f
C488 B.n246 VSUBS 0.008232f
C489 B.n247 VSUBS 0.008232f
C490 B.n248 VSUBS 0.008232f
C491 B.n249 VSUBS 0.018793f
C492 B.n250 VSUBS 0.020432f
C493 B.n251 VSUBS 0.019485f
C494 B.n252 VSUBS 0.008232f
C495 B.n253 VSUBS 0.008232f
C496 B.n254 VSUBS 0.008232f
C497 B.n255 VSUBS 0.008232f
C498 B.n256 VSUBS 0.008232f
C499 B.n257 VSUBS 0.008232f
C500 B.n258 VSUBS 0.008232f
C501 B.n259 VSUBS 0.008232f
C502 B.n260 VSUBS 0.008232f
C503 B.n261 VSUBS 0.008232f
C504 B.n262 VSUBS 0.008232f
C505 B.n263 VSUBS 0.008232f
C506 B.n264 VSUBS 0.008232f
C507 B.n265 VSUBS 0.008232f
C508 B.n266 VSUBS 0.008232f
C509 B.n267 VSUBS 0.008232f
C510 B.n268 VSUBS 0.008232f
C511 B.n269 VSUBS 0.008232f
C512 B.n270 VSUBS 0.008232f
C513 B.n271 VSUBS 0.008232f
C514 B.n272 VSUBS 0.008232f
C515 B.n273 VSUBS 0.008232f
C516 B.n274 VSUBS 0.008232f
C517 B.n275 VSUBS 0.008232f
C518 B.n276 VSUBS 0.008232f
C519 B.n277 VSUBS 0.008232f
C520 B.n278 VSUBS 0.008232f
C521 B.n279 VSUBS 0.008232f
C522 B.n280 VSUBS 0.008232f
C523 B.n281 VSUBS 0.008232f
C524 B.n282 VSUBS 0.008232f
C525 B.n283 VSUBS 0.008232f
C526 B.n284 VSUBS 0.008232f
C527 B.n285 VSUBS 0.008232f
C528 B.n286 VSUBS 0.008232f
C529 B.n287 VSUBS 0.008232f
C530 B.n288 VSUBS 0.008232f
C531 B.n289 VSUBS 0.008232f
C532 B.n290 VSUBS 0.008232f
C533 B.n291 VSUBS 0.008232f
C534 B.n292 VSUBS 0.008232f
C535 B.n293 VSUBS 0.008232f
C536 B.n294 VSUBS 0.008232f
C537 B.n295 VSUBS 0.008232f
C538 B.n296 VSUBS 0.008232f
C539 B.n297 VSUBS 0.008232f
C540 B.n298 VSUBS 0.008232f
C541 B.n299 VSUBS 0.008232f
C542 B.n300 VSUBS 0.008232f
C543 B.n301 VSUBS 0.008232f
C544 B.n302 VSUBS 0.008232f
C545 B.n303 VSUBS 0.008232f
C546 B.n304 VSUBS 0.008232f
C547 B.n305 VSUBS 0.008232f
C548 B.n306 VSUBS 0.008232f
C549 B.n307 VSUBS 0.008232f
C550 B.n308 VSUBS 0.008232f
C551 B.n309 VSUBS 0.008232f
C552 B.n310 VSUBS 0.008232f
C553 B.n311 VSUBS 0.008232f
C554 B.n312 VSUBS 0.008232f
C555 B.n313 VSUBS 0.008232f
C556 B.n314 VSUBS 0.008232f
C557 B.n315 VSUBS 0.008232f
C558 B.n316 VSUBS 0.008232f
C559 B.n317 VSUBS 0.008232f
C560 B.n318 VSUBS 0.008232f
C561 B.n319 VSUBS 0.008232f
C562 B.n320 VSUBS 0.008232f
C563 B.n321 VSUBS 0.008232f
C564 B.n322 VSUBS 0.008232f
C565 B.n323 VSUBS 0.008232f
C566 B.n324 VSUBS 0.008232f
C567 B.n325 VSUBS 0.008232f
C568 B.n326 VSUBS 0.008232f
C569 B.n327 VSUBS 0.008232f
C570 B.n328 VSUBS 0.008232f
C571 B.n329 VSUBS 0.008232f
C572 B.n330 VSUBS 0.008232f
C573 B.n331 VSUBS 0.008232f
C574 B.n332 VSUBS 0.008232f
C575 B.n333 VSUBS 0.008232f
C576 B.n334 VSUBS 0.008232f
C577 B.n335 VSUBS 0.008232f
C578 B.n336 VSUBS 0.008232f
C579 B.n337 VSUBS 0.008232f
C580 B.n338 VSUBS 0.008232f
C581 B.n339 VSUBS 0.008232f
C582 B.n340 VSUBS 0.008232f
C583 B.n341 VSUBS 0.008232f
C584 B.n342 VSUBS 0.008232f
C585 B.n343 VSUBS 0.008232f
C586 B.n344 VSUBS 0.008232f
C587 B.n345 VSUBS 0.008232f
C588 B.n346 VSUBS 0.008232f
C589 B.n347 VSUBS 0.008232f
C590 B.n348 VSUBS 0.008232f
C591 B.n349 VSUBS 0.008232f
C592 B.n350 VSUBS 0.008232f
C593 B.n351 VSUBS 0.019485f
C594 B.n352 VSUBS 0.019739f
C595 B.n353 VSUBS 0.019739f
C596 B.n354 VSUBS 0.008232f
C597 B.n355 VSUBS 0.008232f
C598 B.n356 VSUBS 0.008232f
C599 B.n357 VSUBS 0.008232f
C600 B.n358 VSUBS 0.008232f
C601 B.n359 VSUBS 0.008232f
C602 B.n360 VSUBS 0.008232f
C603 B.n361 VSUBS 0.008232f
C604 B.n362 VSUBS 0.008232f
C605 B.n363 VSUBS 0.008232f
C606 B.n364 VSUBS 0.008232f
C607 B.n365 VSUBS 0.008232f
C608 B.n366 VSUBS 0.008232f
C609 B.n367 VSUBS 0.008232f
C610 B.n368 VSUBS 0.008232f
C611 B.n369 VSUBS 0.008232f
C612 B.n370 VSUBS 0.008232f
C613 B.n371 VSUBS 0.008232f
C614 B.n372 VSUBS 0.008232f
C615 B.n373 VSUBS 0.008232f
C616 B.n374 VSUBS 0.008232f
C617 B.n375 VSUBS 0.008232f
C618 B.n376 VSUBS 0.008232f
C619 B.n377 VSUBS 0.008232f
C620 B.n378 VSUBS 0.008232f
C621 B.n379 VSUBS 0.008232f
C622 B.n380 VSUBS 0.008232f
C623 B.n381 VSUBS 0.00569f
C624 B.n382 VSUBS 0.019073f
C625 B.n383 VSUBS 0.006659f
C626 B.n384 VSUBS 0.008232f
C627 B.n385 VSUBS 0.008232f
C628 B.n386 VSUBS 0.008232f
C629 B.n387 VSUBS 0.008232f
C630 B.n388 VSUBS 0.008232f
C631 B.n389 VSUBS 0.008232f
C632 B.n390 VSUBS 0.008232f
C633 B.n391 VSUBS 0.008232f
C634 B.n392 VSUBS 0.008232f
C635 B.n393 VSUBS 0.008232f
C636 B.n394 VSUBS 0.008232f
C637 B.n395 VSUBS 0.006659f
C638 B.n396 VSUBS 0.008232f
C639 B.n397 VSUBS 0.008232f
C640 B.n398 VSUBS 0.008232f
C641 B.n399 VSUBS 0.008232f
C642 B.n400 VSUBS 0.008232f
C643 B.n401 VSUBS 0.008232f
C644 B.n402 VSUBS 0.008232f
C645 B.n403 VSUBS 0.008232f
C646 B.n404 VSUBS 0.008232f
C647 B.n405 VSUBS 0.008232f
C648 B.n406 VSUBS 0.008232f
C649 B.n407 VSUBS 0.008232f
C650 B.n408 VSUBS 0.008232f
C651 B.n409 VSUBS 0.008232f
C652 B.n410 VSUBS 0.008232f
C653 B.n411 VSUBS 0.008232f
C654 B.n412 VSUBS 0.008232f
C655 B.n413 VSUBS 0.008232f
C656 B.n414 VSUBS 0.008232f
C657 B.n415 VSUBS 0.008232f
C658 B.n416 VSUBS 0.008232f
C659 B.n417 VSUBS 0.008232f
C660 B.n418 VSUBS 0.008232f
C661 B.n419 VSUBS 0.008232f
C662 B.n420 VSUBS 0.008232f
C663 B.n421 VSUBS 0.008232f
C664 B.n422 VSUBS 0.008232f
C665 B.n423 VSUBS 0.008232f
C666 B.n424 VSUBS 0.008232f
C667 B.n425 VSUBS 0.019739f
C668 B.n426 VSUBS 0.019739f
C669 B.n427 VSUBS 0.019485f
C670 B.n428 VSUBS 0.008232f
C671 B.n429 VSUBS 0.008232f
C672 B.n430 VSUBS 0.008232f
C673 B.n431 VSUBS 0.008232f
C674 B.n432 VSUBS 0.008232f
C675 B.n433 VSUBS 0.008232f
C676 B.n434 VSUBS 0.008232f
C677 B.n435 VSUBS 0.008232f
C678 B.n436 VSUBS 0.008232f
C679 B.n437 VSUBS 0.008232f
C680 B.n438 VSUBS 0.008232f
C681 B.n439 VSUBS 0.008232f
C682 B.n440 VSUBS 0.008232f
C683 B.n441 VSUBS 0.008232f
C684 B.n442 VSUBS 0.008232f
C685 B.n443 VSUBS 0.008232f
C686 B.n444 VSUBS 0.008232f
C687 B.n445 VSUBS 0.008232f
C688 B.n446 VSUBS 0.008232f
C689 B.n447 VSUBS 0.008232f
C690 B.n448 VSUBS 0.008232f
C691 B.n449 VSUBS 0.008232f
C692 B.n450 VSUBS 0.008232f
C693 B.n451 VSUBS 0.008232f
C694 B.n452 VSUBS 0.008232f
C695 B.n453 VSUBS 0.008232f
C696 B.n454 VSUBS 0.008232f
C697 B.n455 VSUBS 0.008232f
C698 B.n456 VSUBS 0.008232f
C699 B.n457 VSUBS 0.008232f
C700 B.n458 VSUBS 0.008232f
C701 B.n459 VSUBS 0.008232f
C702 B.n460 VSUBS 0.008232f
C703 B.n461 VSUBS 0.008232f
C704 B.n462 VSUBS 0.008232f
C705 B.n463 VSUBS 0.008232f
C706 B.n464 VSUBS 0.008232f
C707 B.n465 VSUBS 0.008232f
C708 B.n466 VSUBS 0.008232f
C709 B.n467 VSUBS 0.008232f
C710 B.n468 VSUBS 0.008232f
C711 B.n469 VSUBS 0.008232f
C712 B.n470 VSUBS 0.008232f
C713 B.n471 VSUBS 0.008232f
C714 B.n472 VSUBS 0.008232f
C715 B.n473 VSUBS 0.008232f
C716 B.n474 VSUBS 0.008232f
C717 B.n475 VSUBS 0.010743f
C718 B.n476 VSUBS 0.011444f
C719 B.n477 VSUBS 0.022757f
.ends

