* NGSPICE file created from diff_pair_sample_0488.ext - technology: sky130A

.subckt diff_pair_sample_0488 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=3.89
X1 VTAIL.t5 VP.t0 VDD1.t7 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=3.89
X2 VDD1.t6 VP.t1 VTAIL.t3 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=3.89
X3 B.t11 B.t9 B.t10 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=3.89
X4 B.t8 B.t6 B.t7 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=3.89
X5 VTAIL.t14 VN.t1 VDD2.t2 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X6 VTAIL.t7 VP.t2 VDD1.t5 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=3.89
X7 VTAIL.t6 VP.t3 VDD1.t4 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X8 VDD1.t3 VP.t4 VTAIL.t0 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X9 VDD1.t2 VP.t5 VTAIL.t1 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X10 VDD2.t1 VN.t2 VTAIL.t13 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X11 VTAIL.t12 VN.t3 VDD2.t0 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=3.89
X12 VDD2.t5 VN.t4 VTAIL.t11 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=3.89
X13 B.t5 B.t3 B.t4 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=3.89
X14 B.t2 B.t0 B.t1 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=3.89
X15 VDD1.t1 VP.t6 VTAIL.t2 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=3.89
X16 VTAIL.t4 VP.t7 VDD1.t0 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X17 VTAIL.t10 VN.t5 VDD2.t4 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X18 VDD2.t7 VN.t6 VTAIL.t9 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=2.90565 ps=17.94 w=17.61 l=3.89
X19 VDD2.t6 VN.t7 VTAIL.t8 w_n5190_n4490# sky130_fd_pr__pfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=3.89
R0 VN.n76 VN.n75 161.3
R1 VN.n74 VN.n40 161.3
R2 VN.n73 VN.n72 161.3
R3 VN.n71 VN.n41 161.3
R4 VN.n70 VN.n69 161.3
R5 VN.n68 VN.n42 161.3
R6 VN.n67 VN.n66 161.3
R7 VN.n65 VN.n43 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n61 VN.n44 161.3
R10 VN.n60 VN.n59 161.3
R11 VN.n58 VN.n45 161.3
R12 VN.n57 VN.n56 161.3
R13 VN.n55 VN.n46 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n47 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n1 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n2 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n3 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n4 161.3
R25 VN.n25 VN.n24 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n48 VN.t4 142.212
R35 VN.n9 VN.t0 142.212
R36 VN.n10 VN.t6 109.102
R37 VN.n23 VN.t1 109.102
R38 VN.n0 VN.t7 109.102
R39 VN.n49 VN.t5 109.102
R40 VN.n62 VN.t2 109.102
R41 VN.n39 VN.t3 109.102
R42 VN.n38 VN.n0 86.1527
R43 VN.n77 VN.n39 86.1527
R44 VN VN.n77 61.4374
R45 VN.n49 VN.n48 57.4697
R46 VN.n10 VN.n9 57.4697
R47 VN.n17 VN.n16 56.5193
R48 VN.n56 VN.n55 56.5193
R49 VN.n30 VN.n29 43.4072
R50 VN.n69 VN.n68 43.4072
R51 VN.n30 VN.n2 37.5796
R52 VN.n69 VN.n41 37.5796
R53 VN.n11 VN.n8 24.4675
R54 VN.n15 VN.n8 24.4675
R55 VN.n16 VN.n15 24.4675
R56 VN.n17 VN.n6 24.4675
R57 VN.n21 VN.n6 24.4675
R58 VN.n22 VN.n21 24.4675
R59 VN.n24 VN.n4 24.4675
R60 VN.n28 VN.n4 24.4675
R61 VN.n29 VN.n28 24.4675
R62 VN.n34 VN.n2 24.4675
R63 VN.n35 VN.n34 24.4675
R64 VN.n36 VN.n35 24.4675
R65 VN.n55 VN.n54 24.4675
R66 VN.n54 VN.n47 24.4675
R67 VN.n50 VN.n47 24.4675
R68 VN.n68 VN.n67 24.4675
R69 VN.n67 VN.n43 24.4675
R70 VN.n63 VN.n43 24.4675
R71 VN.n61 VN.n60 24.4675
R72 VN.n60 VN.n45 24.4675
R73 VN.n56 VN.n45 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n73 24.4675
R76 VN.n73 VN.n41 24.4675
R77 VN.n11 VN.n10 17.6167
R78 VN.n23 VN.n22 17.6167
R79 VN.n50 VN.n49 17.6167
R80 VN.n62 VN.n61 17.6167
R81 VN.n24 VN.n23 6.85126
R82 VN.n63 VN.n62 6.85126
R83 VN.n36 VN.n0 3.91522
R84 VN.n75 VN.n39 3.91522
R85 VN.n51 VN.n48 2.44109
R86 VN.n12 VN.n9 2.44109
R87 VN.n77 VN.n76 0.354971
R88 VN.n38 VN.n37 0.354971
R89 VN VN.n38 0.26696
R90 VN.n76 VN.n40 0.189894
R91 VN.n72 VN.n40 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n70 0.189894
R94 VN.n70 VN.n42 0.189894
R95 VN.n66 VN.n42 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n64 0.189894
R98 VN.n64 VN.n44 0.189894
R99 VN.n59 VN.n44 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n57 0.189894
R102 VN.n57 VN.n46 0.189894
R103 VN.n53 VN.n46 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n51 0.189894
R106 VN.n13 VN.n12 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n14 VN.n7 0.189894
R109 VN.n18 VN.n7 0.189894
R110 VN.n19 VN.n18 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n20 VN.n5 0.189894
R113 VN.n25 VN.n5 0.189894
R114 VN.n26 VN.n25 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n27 VN.n3 0.189894
R117 VN.n31 VN.n3 0.189894
R118 VN.n32 VN.n31 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n33 VN.n1 0.189894
R121 VN.n37 VN.n1 0.189894
R122 VDD2.n2 VDD2.n1 72.5311
R123 VDD2.n2 VDD2.n0 72.5311
R124 VDD2 VDD2.n5 72.5283
R125 VDD2.n4 VDD2.n3 70.7677
R126 VDD2.n4 VDD2.n2 55.267
R127 VDD2 VDD2.n4 1.87766
R128 VDD2.n5 VDD2.t4 1.84633
R129 VDD2.n5 VDD2.t5 1.84633
R130 VDD2.n3 VDD2.t0 1.84633
R131 VDD2.n3 VDD2.t1 1.84633
R132 VDD2.n1 VDD2.t2 1.84633
R133 VDD2.n1 VDD2.t6 1.84633
R134 VDD2.n0 VDD2.t3 1.84633
R135 VDD2.n0 VDD2.t7 1.84633
R136 VTAIL.n786 VTAIL.n694 756.745
R137 VTAIL.n94 VTAIL.n2 756.745
R138 VTAIL.n192 VTAIL.n100 756.745
R139 VTAIL.n292 VTAIL.n200 756.745
R140 VTAIL.n688 VTAIL.n596 756.745
R141 VTAIL.n588 VTAIL.n496 756.745
R142 VTAIL.n490 VTAIL.n398 756.745
R143 VTAIL.n390 VTAIL.n298 756.745
R144 VTAIL.n727 VTAIL.n726 585
R145 VTAIL.n729 VTAIL.n728 585
R146 VTAIL.n722 VTAIL.n721 585
R147 VTAIL.n735 VTAIL.n734 585
R148 VTAIL.n737 VTAIL.n736 585
R149 VTAIL.n718 VTAIL.n717 585
R150 VTAIL.n743 VTAIL.n742 585
R151 VTAIL.n745 VTAIL.n744 585
R152 VTAIL.n714 VTAIL.n713 585
R153 VTAIL.n751 VTAIL.n750 585
R154 VTAIL.n753 VTAIL.n752 585
R155 VTAIL.n710 VTAIL.n709 585
R156 VTAIL.n759 VTAIL.n758 585
R157 VTAIL.n761 VTAIL.n760 585
R158 VTAIL.n706 VTAIL.n705 585
R159 VTAIL.n768 VTAIL.n767 585
R160 VTAIL.n769 VTAIL.n704 585
R161 VTAIL.n771 VTAIL.n770 585
R162 VTAIL.n702 VTAIL.n701 585
R163 VTAIL.n777 VTAIL.n776 585
R164 VTAIL.n779 VTAIL.n778 585
R165 VTAIL.n698 VTAIL.n697 585
R166 VTAIL.n785 VTAIL.n784 585
R167 VTAIL.n787 VTAIL.n786 585
R168 VTAIL.n35 VTAIL.n34 585
R169 VTAIL.n37 VTAIL.n36 585
R170 VTAIL.n30 VTAIL.n29 585
R171 VTAIL.n43 VTAIL.n42 585
R172 VTAIL.n45 VTAIL.n44 585
R173 VTAIL.n26 VTAIL.n25 585
R174 VTAIL.n51 VTAIL.n50 585
R175 VTAIL.n53 VTAIL.n52 585
R176 VTAIL.n22 VTAIL.n21 585
R177 VTAIL.n59 VTAIL.n58 585
R178 VTAIL.n61 VTAIL.n60 585
R179 VTAIL.n18 VTAIL.n17 585
R180 VTAIL.n67 VTAIL.n66 585
R181 VTAIL.n69 VTAIL.n68 585
R182 VTAIL.n14 VTAIL.n13 585
R183 VTAIL.n76 VTAIL.n75 585
R184 VTAIL.n77 VTAIL.n12 585
R185 VTAIL.n79 VTAIL.n78 585
R186 VTAIL.n10 VTAIL.n9 585
R187 VTAIL.n85 VTAIL.n84 585
R188 VTAIL.n87 VTAIL.n86 585
R189 VTAIL.n6 VTAIL.n5 585
R190 VTAIL.n93 VTAIL.n92 585
R191 VTAIL.n95 VTAIL.n94 585
R192 VTAIL.n133 VTAIL.n132 585
R193 VTAIL.n135 VTAIL.n134 585
R194 VTAIL.n128 VTAIL.n127 585
R195 VTAIL.n141 VTAIL.n140 585
R196 VTAIL.n143 VTAIL.n142 585
R197 VTAIL.n124 VTAIL.n123 585
R198 VTAIL.n149 VTAIL.n148 585
R199 VTAIL.n151 VTAIL.n150 585
R200 VTAIL.n120 VTAIL.n119 585
R201 VTAIL.n157 VTAIL.n156 585
R202 VTAIL.n159 VTAIL.n158 585
R203 VTAIL.n116 VTAIL.n115 585
R204 VTAIL.n165 VTAIL.n164 585
R205 VTAIL.n167 VTAIL.n166 585
R206 VTAIL.n112 VTAIL.n111 585
R207 VTAIL.n174 VTAIL.n173 585
R208 VTAIL.n175 VTAIL.n110 585
R209 VTAIL.n177 VTAIL.n176 585
R210 VTAIL.n108 VTAIL.n107 585
R211 VTAIL.n183 VTAIL.n182 585
R212 VTAIL.n185 VTAIL.n184 585
R213 VTAIL.n104 VTAIL.n103 585
R214 VTAIL.n191 VTAIL.n190 585
R215 VTAIL.n193 VTAIL.n192 585
R216 VTAIL.n233 VTAIL.n232 585
R217 VTAIL.n235 VTAIL.n234 585
R218 VTAIL.n228 VTAIL.n227 585
R219 VTAIL.n241 VTAIL.n240 585
R220 VTAIL.n243 VTAIL.n242 585
R221 VTAIL.n224 VTAIL.n223 585
R222 VTAIL.n249 VTAIL.n248 585
R223 VTAIL.n251 VTAIL.n250 585
R224 VTAIL.n220 VTAIL.n219 585
R225 VTAIL.n257 VTAIL.n256 585
R226 VTAIL.n259 VTAIL.n258 585
R227 VTAIL.n216 VTAIL.n215 585
R228 VTAIL.n265 VTAIL.n264 585
R229 VTAIL.n267 VTAIL.n266 585
R230 VTAIL.n212 VTAIL.n211 585
R231 VTAIL.n274 VTAIL.n273 585
R232 VTAIL.n275 VTAIL.n210 585
R233 VTAIL.n277 VTAIL.n276 585
R234 VTAIL.n208 VTAIL.n207 585
R235 VTAIL.n283 VTAIL.n282 585
R236 VTAIL.n285 VTAIL.n284 585
R237 VTAIL.n204 VTAIL.n203 585
R238 VTAIL.n291 VTAIL.n290 585
R239 VTAIL.n293 VTAIL.n292 585
R240 VTAIL.n689 VTAIL.n688 585
R241 VTAIL.n687 VTAIL.n686 585
R242 VTAIL.n600 VTAIL.n599 585
R243 VTAIL.n681 VTAIL.n680 585
R244 VTAIL.n679 VTAIL.n678 585
R245 VTAIL.n604 VTAIL.n603 585
R246 VTAIL.n608 VTAIL.n606 585
R247 VTAIL.n673 VTAIL.n672 585
R248 VTAIL.n671 VTAIL.n670 585
R249 VTAIL.n610 VTAIL.n609 585
R250 VTAIL.n665 VTAIL.n664 585
R251 VTAIL.n663 VTAIL.n662 585
R252 VTAIL.n614 VTAIL.n613 585
R253 VTAIL.n657 VTAIL.n656 585
R254 VTAIL.n655 VTAIL.n654 585
R255 VTAIL.n618 VTAIL.n617 585
R256 VTAIL.n649 VTAIL.n648 585
R257 VTAIL.n647 VTAIL.n646 585
R258 VTAIL.n622 VTAIL.n621 585
R259 VTAIL.n641 VTAIL.n640 585
R260 VTAIL.n639 VTAIL.n638 585
R261 VTAIL.n626 VTAIL.n625 585
R262 VTAIL.n633 VTAIL.n632 585
R263 VTAIL.n631 VTAIL.n630 585
R264 VTAIL.n589 VTAIL.n588 585
R265 VTAIL.n587 VTAIL.n586 585
R266 VTAIL.n500 VTAIL.n499 585
R267 VTAIL.n581 VTAIL.n580 585
R268 VTAIL.n579 VTAIL.n578 585
R269 VTAIL.n504 VTAIL.n503 585
R270 VTAIL.n508 VTAIL.n506 585
R271 VTAIL.n573 VTAIL.n572 585
R272 VTAIL.n571 VTAIL.n570 585
R273 VTAIL.n510 VTAIL.n509 585
R274 VTAIL.n565 VTAIL.n564 585
R275 VTAIL.n563 VTAIL.n562 585
R276 VTAIL.n514 VTAIL.n513 585
R277 VTAIL.n557 VTAIL.n556 585
R278 VTAIL.n555 VTAIL.n554 585
R279 VTAIL.n518 VTAIL.n517 585
R280 VTAIL.n549 VTAIL.n548 585
R281 VTAIL.n547 VTAIL.n546 585
R282 VTAIL.n522 VTAIL.n521 585
R283 VTAIL.n541 VTAIL.n540 585
R284 VTAIL.n539 VTAIL.n538 585
R285 VTAIL.n526 VTAIL.n525 585
R286 VTAIL.n533 VTAIL.n532 585
R287 VTAIL.n531 VTAIL.n530 585
R288 VTAIL.n491 VTAIL.n490 585
R289 VTAIL.n489 VTAIL.n488 585
R290 VTAIL.n402 VTAIL.n401 585
R291 VTAIL.n483 VTAIL.n482 585
R292 VTAIL.n481 VTAIL.n480 585
R293 VTAIL.n406 VTAIL.n405 585
R294 VTAIL.n410 VTAIL.n408 585
R295 VTAIL.n475 VTAIL.n474 585
R296 VTAIL.n473 VTAIL.n472 585
R297 VTAIL.n412 VTAIL.n411 585
R298 VTAIL.n467 VTAIL.n466 585
R299 VTAIL.n465 VTAIL.n464 585
R300 VTAIL.n416 VTAIL.n415 585
R301 VTAIL.n459 VTAIL.n458 585
R302 VTAIL.n457 VTAIL.n456 585
R303 VTAIL.n420 VTAIL.n419 585
R304 VTAIL.n451 VTAIL.n450 585
R305 VTAIL.n449 VTAIL.n448 585
R306 VTAIL.n424 VTAIL.n423 585
R307 VTAIL.n443 VTAIL.n442 585
R308 VTAIL.n441 VTAIL.n440 585
R309 VTAIL.n428 VTAIL.n427 585
R310 VTAIL.n435 VTAIL.n434 585
R311 VTAIL.n433 VTAIL.n432 585
R312 VTAIL.n391 VTAIL.n390 585
R313 VTAIL.n389 VTAIL.n388 585
R314 VTAIL.n302 VTAIL.n301 585
R315 VTAIL.n383 VTAIL.n382 585
R316 VTAIL.n381 VTAIL.n380 585
R317 VTAIL.n306 VTAIL.n305 585
R318 VTAIL.n310 VTAIL.n308 585
R319 VTAIL.n375 VTAIL.n374 585
R320 VTAIL.n373 VTAIL.n372 585
R321 VTAIL.n312 VTAIL.n311 585
R322 VTAIL.n367 VTAIL.n366 585
R323 VTAIL.n365 VTAIL.n364 585
R324 VTAIL.n316 VTAIL.n315 585
R325 VTAIL.n359 VTAIL.n358 585
R326 VTAIL.n357 VTAIL.n356 585
R327 VTAIL.n320 VTAIL.n319 585
R328 VTAIL.n351 VTAIL.n350 585
R329 VTAIL.n349 VTAIL.n348 585
R330 VTAIL.n324 VTAIL.n323 585
R331 VTAIL.n343 VTAIL.n342 585
R332 VTAIL.n341 VTAIL.n340 585
R333 VTAIL.n328 VTAIL.n327 585
R334 VTAIL.n335 VTAIL.n334 585
R335 VTAIL.n333 VTAIL.n332 585
R336 VTAIL.n725 VTAIL.t8 327.466
R337 VTAIL.n33 VTAIL.t15 327.466
R338 VTAIL.n131 VTAIL.t3 327.466
R339 VTAIL.n231 VTAIL.t7 327.466
R340 VTAIL.n629 VTAIL.t2 327.466
R341 VTAIL.n529 VTAIL.t5 327.466
R342 VTAIL.n431 VTAIL.t11 327.466
R343 VTAIL.n331 VTAIL.t12 327.466
R344 VTAIL.n728 VTAIL.n727 171.744
R345 VTAIL.n728 VTAIL.n721 171.744
R346 VTAIL.n735 VTAIL.n721 171.744
R347 VTAIL.n736 VTAIL.n735 171.744
R348 VTAIL.n736 VTAIL.n717 171.744
R349 VTAIL.n743 VTAIL.n717 171.744
R350 VTAIL.n744 VTAIL.n743 171.744
R351 VTAIL.n744 VTAIL.n713 171.744
R352 VTAIL.n751 VTAIL.n713 171.744
R353 VTAIL.n752 VTAIL.n751 171.744
R354 VTAIL.n752 VTAIL.n709 171.744
R355 VTAIL.n759 VTAIL.n709 171.744
R356 VTAIL.n760 VTAIL.n759 171.744
R357 VTAIL.n760 VTAIL.n705 171.744
R358 VTAIL.n768 VTAIL.n705 171.744
R359 VTAIL.n769 VTAIL.n768 171.744
R360 VTAIL.n770 VTAIL.n769 171.744
R361 VTAIL.n770 VTAIL.n701 171.744
R362 VTAIL.n777 VTAIL.n701 171.744
R363 VTAIL.n778 VTAIL.n777 171.744
R364 VTAIL.n778 VTAIL.n697 171.744
R365 VTAIL.n785 VTAIL.n697 171.744
R366 VTAIL.n786 VTAIL.n785 171.744
R367 VTAIL.n36 VTAIL.n35 171.744
R368 VTAIL.n36 VTAIL.n29 171.744
R369 VTAIL.n43 VTAIL.n29 171.744
R370 VTAIL.n44 VTAIL.n43 171.744
R371 VTAIL.n44 VTAIL.n25 171.744
R372 VTAIL.n51 VTAIL.n25 171.744
R373 VTAIL.n52 VTAIL.n51 171.744
R374 VTAIL.n52 VTAIL.n21 171.744
R375 VTAIL.n59 VTAIL.n21 171.744
R376 VTAIL.n60 VTAIL.n59 171.744
R377 VTAIL.n60 VTAIL.n17 171.744
R378 VTAIL.n67 VTAIL.n17 171.744
R379 VTAIL.n68 VTAIL.n67 171.744
R380 VTAIL.n68 VTAIL.n13 171.744
R381 VTAIL.n76 VTAIL.n13 171.744
R382 VTAIL.n77 VTAIL.n76 171.744
R383 VTAIL.n78 VTAIL.n77 171.744
R384 VTAIL.n78 VTAIL.n9 171.744
R385 VTAIL.n85 VTAIL.n9 171.744
R386 VTAIL.n86 VTAIL.n85 171.744
R387 VTAIL.n86 VTAIL.n5 171.744
R388 VTAIL.n93 VTAIL.n5 171.744
R389 VTAIL.n94 VTAIL.n93 171.744
R390 VTAIL.n134 VTAIL.n133 171.744
R391 VTAIL.n134 VTAIL.n127 171.744
R392 VTAIL.n141 VTAIL.n127 171.744
R393 VTAIL.n142 VTAIL.n141 171.744
R394 VTAIL.n142 VTAIL.n123 171.744
R395 VTAIL.n149 VTAIL.n123 171.744
R396 VTAIL.n150 VTAIL.n149 171.744
R397 VTAIL.n150 VTAIL.n119 171.744
R398 VTAIL.n157 VTAIL.n119 171.744
R399 VTAIL.n158 VTAIL.n157 171.744
R400 VTAIL.n158 VTAIL.n115 171.744
R401 VTAIL.n165 VTAIL.n115 171.744
R402 VTAIL.n166 VTAIL.n165 171.744
R403 VTAIL.n166 VTAIL.n111 171.744
R404 VTAIL.n174 VTAIL.n111 171.744
R405 VTAIL.n175 VTAIL.n174 171.744
R406 VTAIL.n176 VTAIL.n175 171.744
R407 VTAIL.n176 VTAIL.n107 171.744
R408 VTAIL.n183 VTAIL.n107 171.744
R409 VTAIL.n184 VTAIL.n183 171.744
R410 VTAIL.n184 VTAIL.n103 171.744
R411 VTAIL.n191 VTAIL.n103 171.744
R412 VTAIL.n192 VTAIL.n191 171.744
R413 VTAIL.n234 VTAIL.n233 171.744
R414 VTAIL.n234 VTAIL.n227 171.744
R415 VTAIL.n241 VTAIL.n227 171.744
R416 VTAIL.n242 VTAIL.n241 171.744
R417 VTAIL.n242 VTAIL.n223 171.744
R418 VTAIL.n249 VTAIL.n223 171.744
R419 VTAIL.n250 VTAIL.n249 171.744
R420 VTAIL.n250 VTAIL.n219 171.744
R421 VTAIL.n257 VTAIL.n219 171.744
R422 VTAIL.n258 VTAIL.n257 171.744
R423 VTAIL.n258 VTAIL.n215 171.744
R424 VTAIL.n265 VTAIL.n215 171.744
R425 VTAIL.n266 VTAIL.n265 171.744
R426 VTAIL.n266 VTAIL.n211 171.744
R427 VTAIL.n274 VTAIL.n211 171.744
R428 VTAIL.n275 VTAIL.n274 171.744
R429 VTAIL.n276 VTAIL.n275 171.744
R430 VTAIL.n276 VTAIL.n207 171.744
R431 VTAIL.n283 VTAIL.n207 171.744
R432 VTAIL.n284 VTAIL.n283 171.744
R433 VTAIL.n284 VTAIL.n203 171.744
R434 VTAIL.n291 VTAIL.n203 171.744
R435 VTAIL.n292 VTAIL.n291 171.744
R436 VTAIL.n688 VTAIL.n687 171.744
R437 VTAIL.n687 VTAIL.n599 171.744
R438 VTAIL.n680 VTAIL.n599 171.744
R439 VTAIL.n680 VTAIL.n679 171.744
R440 VTAIL.n679 VTAIL.n603 171.744
R441 VTAIL.n608 VTAIL.n603 171.744
R442 VTAIL.n672 VTAIL.n608 171.744
R443 VTAIL.n672 VTAIL.n671 171.744
R444 VTAIL.n671 VTAIL.n609 171.744
R445 VTAIL.n664 VTAIL.n609 171.744
R446 VTAIL.n664 VTAIL.n663 171.744
R447 VTAIL.n663 VTAIL.n613 171.744
R448 VTAIL.n656 VTAIL.n613 171.744
R449 VTAIL.n656 VTAIL.n655 171.744
R450 VTAIL.n655 VTAIL.n617 171.744
R451 VTAIL.n648 VTAIL.n617 171.744
R452 VTAIL.n648 VTAIL.n647 171.744
R453 VTAIL.n647 VTAIL.n621 171.744
R454 VTAIL.n640 VTAIL.n621 171.744
R455 VTAIL.n640 VTAIL.n639 171.744
R456 VTAIL.n639 VTAIL.n625 171.744
R457 VTAIL.n632 VTAIL.n625 171.744
R458 VTAIL.n632 VTAIL.n631 171.744
R459 VTAIL.n588 VTAIL.n587 171.744
R460 VTAIL.n587 VTAIL.n499 171.744
R461 VTAIL.n580 VTAIL.n499 171.744
R462 VTAIL.n580 VTAIL.n579 171.744
R463 VTAIL.n579 VTAIL.n503 171.744
R464 VTAIL.n508 VTAIL.n503 171.744
R465 VTAIL.n572 VTAIL.n508 171.744
R466 VTAIL.n572 VTAIL.n571 171.744
R467 VTAIL.n571 VTAIL.n509 171.744
R468 VTAIL.n564 VTAIL.n509 171.744
R469 VTAIL.n564 VTAIL.n563 171.744
R470 VTAIL.n563 VTAIL.n513 171.744
R471 VTAIL.n556 VTAIL.n513 171.744
R472 VTAIL.n556 VTAIL.n555 171.744
R473 VTAIL.n555 VTAIL.n517 171.744
R474 VTAIL.n548 VTAIL.n517 171.744
R475 VTAIL.n548 VTAIL.n547 171.744
R476 VTAIL.n547 VTAIL.n521 171.744
R477 VTAIL.n540 VTAIL.n521 171.744
R478 VTAIL.n540 VTAIL.n539 171.744
R479 VTAIL.n539 VTAIL.n525 171.744
R480 VTAIL.n532 VTAIL.n525 171.744
R481 VTAIL.n532 VTAIL.n531 171.744
R482 VTAIL.n490 VTAIL.n489 171.744
R483 VTAIL.n489 VTAIL.n401 171.744
R484 VTAIL.n482 VTAIL.n401 171.744
R485 VTAIL.n482 VTAIL.n481 171.744
R486 VTAIL.n481 VTAIL.n405 171.744
R487 VTAIL.n410 VTAIL.n405 171.744
R488 VTAIL.n474 VTAIL.n410 171.744
R489 VTAIL.n474 VTAIL.n473 171.744
R490 VTAIL.n473 VTAIL.n411 171.744
R491 VTAIL.n466 VTAIL.n411 171.744
R492 VTAIL.n466 VTAIL.n465 171.744
R493 VTAIL.n465 VTAIL.n415 171.744
R494 VTAIL.n458 VTAIL.n415 171.744
R495 VTAIL.n458 VTAIL.n457 171.744
R496 VTAIL.n457 VTAIL.n419 171.744
R497 VTAIL.n450 VTAIL.n419 171.744
R498 VTAIL.n450 VTAIL.n449 171.744
R499 VTAIL.n449 VTAIL.n423 171.744
R500 VTAIL.n442 VTAIL.n423 171.744
R501 VTAIL.n442 VTAIL.n441 171.744
R502 VTAIL.n441 VTAIL.n427 171.744
R503 VTAIL.n434 VTAIL.n427 171.744
R504 VTAIL.n434 VTAIL.n433 171.744
R505 VTAIL.n390 VTAIL.n389 171.744
R506 VTAIL.n389 VTAIL.n301 171.744
R507 VTAIL.n382 VTAIL.n301 171.744
R508 VTAIL.n382 VTAIL.n381 171.744
R509 VTAIL.n381 VTAIL.n305 171.744
R510 VTAIL.n310 VTAIL.n305 171.744
R511 VTAIL.n374 VTAIL.n310 171.744
R512 VTAIL.n374 VTAIL.n373 171.744
R513 VTAIL.n373 VTAIL.n311 171.744
R514 VTAIL.n366 VTAIL.n311 171.744
R515 VTAIL.n366 VTAIL.n365 171.744
R516 VTAIL.n365 VTAIL.n315 171.744
R517 VTAIL.n358 VTAIL.n315 171.744
R518 VTAIL.n358 VTAIL.n357 171.744
R519 VTAIL.n357 VTAIL.n319 171.744
R520 VTAIL.n350 VTAIL.n319 171.744
R521 VTAIL.n350 VTAIL.n349 171.744
R522 VTAIL.n349 VTAIL.n323 171.744
R523 VTAIL.n342 VTAIL.n323 171.744
R524 VTAIL.n342 VTAIL.n341 171.744
R525 VTAIL.n341 VTAIL.n327 171.744
R526 VTAIL.n334 VTAIL.n327 171.744
R527 VTAIL.n334 VTAIL.n333 171.744
R528 VTAIL.n727 VTAIL.t8 85.8723
R529 VTAIL.n35 VTAIL.t15 85.8723
R530 VTAIL.n133 VTAIL.t3 85.8723
R531 VTAIL.n233 VTAIL.t7 85.8723
R532 VTAIL.n631 VTAIL.t2 85.8723
R533 VTAIL.n531 VTAIL.t5 85.8723
R534 VTAIL.n433 VTAIL.t11 85.8723
R535 VTAIL.n333 VTAIL.t12 85.8723
R536 VTAIL.n595 VTAIL.n594 54.0889
R537 VTAIL.n397 VTAIL.n396 54.0889
R538 VTAIL.n1 VTAIL.n0 54.0887
R539 VTAIL.n199 VTAIL.n198 54.0887
R540 VTAIL.n791 VTAIL.n790 33.9308
R541 VTAIL.n99 VTAIL.n98 33.9308
R542 VTAIL.n197 VTAIL.n196 33.9308
R543 VTAIL.n297 VTAIL.n296 33.9308
R544 VTAIL.n693 VTAIL.n692 33.9308
R545 VTAIL.n593 VTAIL.n592 33.9308
R546 VTAIL.n495 VTAIL.n494 33.9308
R547 VTAIL.n395 VTAIL.n394 33.9308
R548 VTAIL.n791 VTAIL.n693 31.1858
R549 VTAIL.n395 VTAIL.n297 31.1858
R550 VTAIL.n726 VTAIL.n725 16.3895
R551 VTAIL.n34 VTAIL.n33 16.3895
R552 VTAIL.n132 VTAIL.n131 16.3895
R553 VTAIL.n232 VTAIL.n231 16.3895
R554 VTAIL.n630 VTAIL.n629 16.3895
R555 VTAIL.n530 VTAIL.n529 16.3895
R556 VTAIL.n432 VTAIL.n431 16.3895
R557 VTAIL.n332 VTAIL.n331 16.3895
R558 VTAIL.n771 VTAIL.n702 13.1884
R559 VTAIL.n79 VTAIL.n10 13.1884
R560 VTAIL.n177 VTAIL.n108 13.1884
R561 VTAIL.n277 VTAIL.n208 13.1884
R562 VTAIL.n606 VTAIL.n604 13.1884
R563 VTAIL.n506 VTAIL.n504 13.1884
R564 VTAIL.n408 VTAIL.n406 13.1884
R565 VTAIL.n308 VTAIL.n306 13.1884
R566 VTAIL.n729 VTAIL.n724 12.8005
R567 VTAIL.n772 VTAIL.n704 12.8005
R568 VTAIL.n776 VTAIL.n775 12.8005
R569 VTAIL.n37 VTAIL.n32 12.8005
R570 VTAIL.n80 VTAIL.n12 12.8005
R571 VTAIL.n84 VTAIL.n83 12.8005
R572 VTAIL.n135 VTAIL.n130 12.8005
R573 VTAIL.n178 VTAIL.n110 12.8005
R574 VTAIL.n182 VTAIL.n181 12.8005
R575 VTAIL.n235 VTAIL.n230 12.8005
R576 VTAIL.n278 VTAIL.n210 12.8005
R577 VTAIL.n282 VTAIL.n281 12.8005
R578 VTAIL.n678 VTAIL.n677 12.8005
R579 VTAIL.n674 VTAIL.n673 12.8005
R580 VTAIL.n633 VTAIL.n628 12.8005
R581 VTAIL.n578 VTAIL.n577 12.8005
R582 VTAIL.n574 VTAIL.n573 12.8005
R583 VTAIL.n533 VTAIL.n528 12.8005
R584 VTAIL.n480 VTAIL.n479 12.8005
R585 VTAIL.n476 VTAIL.n475 12.8005
R586 VTAIL.n435 VTAIL.n430 12.8005
R587 VTAIL.n380 VTAIL.n379 12.8005
R588 VTAIL.n376 VTAIL.n375 12.8005
R589 VTAIL.n335 VTAIL.n330 12.8005
R590 VTAIL.n730 VTAIL.n722 12.0247
R591 VTAIL.n767 VTAIL.n766 12.0247
R592 VTAIL.n779 VTAIL.n700 12.0247
R593 VTAIL.n38 VTAIL.n30 12.0247
R594 VTAIL.n75 VTAIL.n74 12.0247
R595 VTAIL.n87 VTAIL.n8 12.0247
R596 VTAIL.n136 VTAIL.n128 12.0247
R597 VTAIL.n173 VTAIL.n172 12.0247
R598 VTAIL.n185 VTAIL.n106 12.0247
R599 VTAIL.n236 VTAIL.n228 12.0247
R600 VTAIL.n273 VTAIL.n272 12.0247
R601 VTAIL.n285 VTAIL.n206 12.0247
R602 VTAIL.n681 VTAIL.n602 12.0247
R603 VTAIL.n670 VTAIL.n607 12.0247
R604 VTAIL.n634 VTAIL.n626 12.0247
R605 VTAIL.n581 VTAIL.n502 12.0247
R606 VTAIL.n570 VTAIL.n507 12.0247
R607 VTAIL.n534 VTAIL.n526 12.0247
R608 VTAIL.n483 VTAIL.n404 12.0247
R609 VTAIL.n472 VTAIL.n409 12.0247
R610 VTAIL.n436 VTAIL.n428 12.0247
R611 VTAIL.n383 VTAIL.n304 12.0247
R612 VTAIL.n372 VTAIL.n309 12.0247
R613 VTAIL.n336 VTAIL.n328 12.0247
R614 VTAIL.n734 VTAIL.n733 11.249
R615 VTAIL.n765 VTAIL.n706 11.249
R616 VTAIL.n780 VTAIL.n698 11.249
R617 VTAIL.n42 VTAIL.n41 11.249
R618 VTAIL.n73 VTAIL.n14 11.249
R619 VTAIL.n88 VTAIL.n6 11.249
R620 VTAIL.n140 VTAIL.n139 11.249
R621 VTAIL.n171 VTAIL.n112 11.249
R622 VTAIL.n186 VTAIL.n104 11.249
R623 VTAIL.n240 VTAIL.n239 11.249
R624 VTAIL.n271 VTAIL.n212 11.249
R625 VTAIL.n286 VTAIL.n204 11.249
R626 VTAIL.n682 VTAIL.n600 11.249
R627 VTAIL.n669 VTAIL.n610 11.249
R628 VTAIL.n638 VTAIL.n637 11.249
R629 VTAIL.n582 VTAIL.n500 11.249
R630 VTAIL.n569 VTAIL.n510 11.249
R631 VTAIL.n538 VTAIL.n537 11.249
R632 VTAIL.n484 VTAIL.n402 11.249
R633 VTAIL.n471 VTAIL.n412 11.249
R634 VTAIL.n440 VTAIL.n439 11.249
R635 VTAIL.n384 VTAIL.n302 11.249
R636 VTAIL.n371 VTAIL.n312 11.249
R637 VTAIL.n340 VTAIL.n339 11.249
R638 VTAIL.n737 VTAIL.n720 10.4732
R639 VTAIL.n762 VTAIL.n761 10.4732
R640 VTAIL.n784 VTAIL.n783 10.4732
R641 VTAIL.n45 VTAIL.n28 10.4732
R642 VTAIL.n70 VTAIL.n69 10.4732
R643 VTAIL.n92 VTAIL.n91 10.4732
R644 VTAIL.n143 VTAIL.n126 10.4732
R645 VTAIL.n168 VTAIL.n167 10.4732
R646 VTAIL.n190 VTAIL.n189 10.4732
R647 VTAIL.n243 VTAIL.n226 10.4732
R648 VTAIL.n268 VTAIL.n267 10.4732
R649 VTAIL.n290 VTAIL.n289 10.4732
R650 VTAIL.n686 VTAIL.n685 10.4732
R651 VTAIL.n666 VTAIL.n665 10.4732
R652 VTAIL.n641 VTAIL.n624 10.4732
R653 VTAIL.n586 VTAIL.n585 10.4732
R654 VTAIL.n566 VTAIL.n565 10.4732
R655 VTAIL.n541 VTAIL.n524 10.4732
R656 VTAIL.n488 VTAIL.n487 10.4732
R657 VTAIL.n468 VTAIL.n467 10.4732
R658 VTAIL.n443 VTAIL.n426 10.4732
R659 VTAIL.n388 VTAIL.n387 10.4732
R660 VTAIL.n368 VTAIL.n367 10.4732
R661 VTAIL.n343 VTAIL.n326 10.4732
R662 VTAIL.n738 VTAIL.n718 9.69747
R663 VTAIL.n758 VTAIL.n708 9.69747
R664 VTAIL.n787 VTAIL.n696 9.69747
R665 VTAIL.n46 VTAIL.n26 9.69747
R666 VTAIL.n66 VTAIL.n16 9.69747
R667 VTAIL.n95 VTAIL.n4 9.69747
R668 VTAIL.n144 VTAIL.n124 9.69747
R669 VTAIL.n164 VTAIL.n114 9.69747
R670 VTAIL.n193 VTAIL.n102 9.69747
R671 VTAIL.n244 VTAIL.n224 9.69747
R672 VTAIL.n264 VTAIL.n214 9.69747
R673 VTAIL.n293 VTAIL.n202 9.69747
R674 VTAIL.n689 VTAIL.n598 9.69747
R675 VTAIL.n662 VTAIL.n612 9.69747
R676 VTAIL.n642 VTAIL.n622 9.69747
R677 VTAIL.n589 VTAIL.n498 9.69747
R678 VTAIL.n562 VTAIL.n512 9.69747
R679 VTAIL.n542 VTAIL.n522 9.69747
R680 VTAIL.n491 VTAIL.n400 9.69747
R681 VTAIL.n464 VTAIL.n414 9.69747
R682 VTAIL.n444 VTAIL.n424 9.69747
R683 VTAIL.n391 VTAIL.n300 9.69747
R684 VTAIL.n364 VTAIL.n314 9.69747
R685 VTAIL.n344 VTAIL.n324 9.69747
R686 VTAIL.n790 VTAIL.n789 9.45567
R687 VTAIL.n98 VTAIL.n97 9.45567
R688 VTAIL.n196 VTAIL.n195 9.45567
R689 VTAIL.n296 VTAIL.n295 9.45567
R690 VTAIL.n692 VTAIL.n691 9.45567
R691 VTAIL.n592 VTAIL.n591 9.45567
R692 VTAIL.n494 VTAIL.n493 9.45567
R693 VTAIL.n394 VTAIL.n393 9.45567
R694 VTAIL.n789 VTAIL.n788 9.3005
R695 VTAIL.n696 VTAIL.n695 9.3005
R696 VTAIL.n783 VTAIL.n782 9.3005
R697 VTAIL.n781 VTAIL.n780 9.3005
R698 VTAIL.n700 VTAIL.n699 9.3005
R699 VTAIL.n775 VTAIL.n774 9.3005
R700 VTAIL.n747 VTAIL.n746 9.3005
R701 VTAIL.n716 VTAIL.n715 9.3005
R702 VTAIL.n741 VTAIL.n740 9.3005
R703 VTAIL.n739 VTAIL.n738 9.3005
R704 VTAIL.n720 VTAIL.n719 9.3005
R705 VTAIL.n733 VTAIL.n732 9.3005
R706 VTAIL.n731 VTAIL.n730 9.3005
R707 VTAIL.n724 VTAIL.n723 9.3005
R708 VTAIL.n749 VTAIL.n748 9.3005
R709 VTAIL.n712 VTAIL.n711 9.3005
R710 VTAIL.n755 VTAIL.n754 9.3005
R711 VTAIL.n757 VTAIL.n756 9.3005
R712 VTAIL.n708 VTAIL.n707 9.3005
R713 VTAIL.n763 VTAIL.n762 9.3005
R714 VTAIL.n765 VTAIL.n764 9.3005
R715 VTAIL.n766 VTAIL.n703 9.3005
R716 VTAIL.n773 VTAIL.n772 9.3005
R717 VTAIL.n97 VTAIL.n96 9.3005
R718 VTAIL.n4 VTAIL.n3 9.3005
R719 VTAIL.n91 VTAIL.n90 9.3005
R720 VTAIL.n89 VTAIL.n88 9.3005
R721 VTAIL.n8 VTAIL.n7 9.3005
R722 VTAIL.n83 VTAIL.n82 9.3005
R723 VTAIL.n55 VTAIL.n54 9.3005
R724 VTAIL.n24 VTAIL.n23 9.3005
R725 VTAIL.n49 VTAIL.n48 9.3005
R726 VTAIL.n47 VTAIL.n46 9.3005
R727 VTAIL.n28 VTAIL.n27 9.3005
R728 VTAIL.n41 VTAIL.n40 9.3005
R729 VTAIL.n39 VTAIL.n38 9.3005
R730 VTAIL.n32 VTAIL.n31 9.3005
R731 VTAIL.n57 VTAIL.n56 9.3005
R732 VTAIL.n20 VTAIL.n19 9.3005
R733 VTAIL.n63 VTAIL.n62 9.3005
R734 VTAIL.n65 VTAIL.n64 9.3005
R735 VTAIL.n16 VTAIL.n15 9.3005
R736 VTAIL.n71 VTAIL.n70 9.3005
R737 VTAIL.n73 VTAIL.n72 9.3005
R738 VTAIL.n74 VTAIL.n11 9.3005
R739 VTAIL.n81 VTAIL.n80 9.3005
R740 VTAIL.n195 VTAIL.n194 9.3005
R741 VTAIL.n102 VTAIL.n101 9.3005
R742 VTAIL.n189 VTAIL.n188 9.3005
R743 VTAIL.n187 VTAIL.n186 9.3005
R744 VTAIL.n106 VTAIL.n105 9.3005
R745 VTAIL.n181 VTAIL.n180 9.3005
R746 VTAIL.n153 VTAIL.n152 9.3005
R747 VTAIL.n122 VTAIL.n121 9.3005
R748 VTAIL.n147 VTAIL.n146 9.3005
R749 VTAIL.n145 VTAIL.n144 9.3005
R750 VTAIL.n126 VTAIL.n125 9.3005
R751 VTAIL.n139 VTAIL.n138 9.3005
R752 VTAIL.n137 VTAIL.n136 9.3005
R753 VTAIL.n130 VTAIL.n129 9.3005
R754 VTAIL.n155 VTAIL.n154 9.3005
R755 VTAIL.n118 VTAIL.n117 9.3005
R756 VTAIL.n161 VTAIL.n160 9.3005
R757 VTAIL.n163 VTAIL.n162 9.3005
R758 VTAIL.n114 VTAIL.n113 9.3005
R759 VTAIL.n169 VTAIL.n168 9.3005
R760 VTAIL.n171 VTAIL.n170 9.3005
R761 VTAIL.n172 VTAIL.n109 9.3005
R762 VTAIL.n179 VTAIL.n178 9.3005
R763 VTAIL.n295 VTAIL.n294 9.3005
R764 VTAIL.n202 VTAIL.n201 9.3005
R765 VTAIL.n289 VTAIL.n288 9.3005
R766 VTAIL.n287 VTAIL.n286 9.3005
R767 VTAIL.n206 VTAIL.n205 9.3005
R768 VTAIL.n281 VTAIL.n280 9.3005
R769 VTAIL.n253 VTAIL.n252 9.3005
R770 VTAIL.n222 VTAIL.n221 9.3005
R771 VTAIL.n247 VTAIL.n246 9.3005
R772 VTAIL.n245 VTAIL.n244 9.3005
R773 VTAIL.n226 VTAIL.n225 9.3005
R774 VTAIL.n239 VTAIL.n238 9.3005
R775 VTAIL.n237 VTAIL.n236 9.3005
R776 VTAIL.n230 VTAIL.n229 9.3005
R777 VTAIL.n255 VTAIL.n254 9.3005
R778 VTAIL.n218 VTAIL.n217 9.3005
R779 VTAIL.n261 VTAIL.n260 9.3005
R780 VTAIL.n263 VTAIL.n262 9.3005
R781 VTAIL.n214 VTAIL.n213 9.3005
R782 VTAIL.n269 VTAIL.n268 9.3005
R783 VTAIL.n271 VTAIL.n270 9.3005
R784 VTAIL.n272 VTAIL.n209 9.3005
R785 VTAIL.n279 VTAIL.n278 9.3005
R786 VTAIL.n616 VTAIL.n615 9.3005
R787 VTAIL.n659 VTAIL.n658 9.3005
R788 VTAIL.n661 VTAIL.n660 9.3005
R789 VTAIL.n612 VTAIL.n611 9.3005
R790 VTAIL.n667 VTAIL.n666 9.3005
R791 VTAIL.n669 VTAIL.n668 9.3005
R792 VTAIL.n607 VTAIL.n605 9.3005
R793 VTAIL.n675 VTAIL.n674 9.3005
R794 VTAIL.n691 VTAIL.n690 9.3005
R795 VTAIL.n598 VTAIL.n597 9.3005
R796 VTAIL.n685 VTAIL.n684 9.3005
R797 VTAIL.n683 VTAIL.n682 9.3005
R798 VTAIL.n602 VTAIL.n601 9.3005
R799 VTAIL.n677 VTAIL.n676 9.3005
R800 VTAIL.n653 VTAIL.n652 9.3005
R801 VTAIL.n651 VTAIL.n650 9.3005
R802 VTAIL.n620 VTAIL.n619 9.3005
R803 VTAIL.n645 VTAIL.n644 9.3005
R804 VTAIL.n643 VTAIL.n642 9.3005
R805 VTAIL.n624 VTAIL.n623 9.3005
R806 VTAIL.n637 VTAIL.n636 9.3005
R807 VTAIL.n635 VTAIL.n634 9.3005
R808 VTAIL.n628 VTAIL.n627 9.3005
R809 VTAIL.n516 VTAIL.n515 9.3005
R810 VTAIL.n559 VTAIL.n558 9.3005
R811 VTAIL.n561 VTAIL.n560 9.3005
R812 VTAIL.n512 VTAIL.n511 9.3005
R813 VTAIL.n567 VTAIL.n566 9.3005
R814 VTAIL.n569 VTAIL.n568 9.3005
R815 VTAIL.n507 VTAIL.n505 9.3005
R816 VTAIL.n575 VTAIL.n574 9.3005
R817 VTAIL.n591 VTAIL.n590 9.3005
R818 VTAIL.n498 VTAIL.n497 9.3005
R819 VTAIL.n585 VTAIL.n584 9.3005
R820 VTAIL.n583 VTAIL.n582 9.3005
R821 VTAIL.n502 VTAIL.n501 9.3005
R822 VTAIL.n577 VTAIL.n576 9.3005
R823 VTAIL.n553 VTAIL.n552 9.3005
R824 VTAIL.n551 VTAIL.n550 9.3005
R825 VTAIL.n520 VTAIL.n519 9.3005
R826 VTAIL.n545 VTAIL.n544 9.3005
R827 VTAIL.n543 VTAIL.n542 9.3005
R828 VTAIL.n524 VTAIL.n523 9.3005
R829 VTAIL.n537 VTAIL.n536 9.3005
R830 VTAIL.n535 VTAIL.n534 9.3005
R831 VTAIL.n528 VTAIL.n527 9.3005
R832 VTAIL.n418 VTAIL.n417 9.3005
R833 VTAIL.n461 VTAIL.n460 9.3005
R834 VTAIL.n463 VTAIL.n462 9.3005
R835 VTAIL.n414 VTAIL.n413 9.3005
R836 VTAIL.n469 VTAIL.n468 9.3005
R837 VTAIL.n471 VTAIL.n470 9.3005
R838 VTAIL.n409 VTAIL.n407 9.3005
R839 VTAIL.n477 VTAIL.n476 9.3005
R840 VTAIL.n493 VTAIL.n492 9.3005
R841 VTAIL.n400 VTAIL.n399 9.3005
R842 VTAIL.n487 VTAIL.n486 9.3005
R843 VTAIL.n485 VTAIL.n484 9.3005
R844 VTAIL.n404 VTAIL.n403 9.3005
R845 VTAIL.n479 VTAIL.n478 9.3005
R846 VTAIL.n455 VTAIL.n454 9.3005
R847 VTAIL.n453 VTAIL.n452 9.3005
R848 VTAIL.n422 VTAIL.n421 9.3005
R849 VTAIL.n447 VTAIL.n446 9.3005
R850 VTAIL.n445 VTAIL.n444 9.3005
R851 VTAIL.n426 VTAIL.n425 9.3005
R852 VTAIL.n439 VTAIL.n438 9.3005
R853 VTAIL.n437 VTAIL.n436 9.3005
R854 VTAIL.n430 VTAIL.n429 9.3005
R855 VTAIL.n318 VTAIL.n317 9.3005
R856 VTAIL.n361 VTAIL.n360 9.3005
R857 VTAIL.n363 VTAIL.n362 9.3005
R858 VTAIL.n314 VTAIL.n313 9.3005
R859 VTAIL.n369 VTAIL.n368 9.3005
R860 VTAIL.n371 VTAIL.n370 9.3005
R861 VTAIL.n309 VTAIL.n307 9.3005
R862 VTAIL.n377 VTAIL.n376 9.3005
R863 VTAIL.n393 VTAIL.n392 9.3005
R864 VTAIL.n300 VTAIL.n299 9.3005
R865 VTAIL.n387 VTAIL.n386 9.3005
R866 VTAIL.n385 VTAIL.n384 9.3005
R867 VTAIL.n304 VTAIL.n303 9.3005
R868 VTAIL.n379 VTAIL.n378 9.3005
R869 VTAIL.n355 VTAIL.n354 9.3005
R870 VTAIL.n353 VTAIL.n352 9.3005
R871 VTAIL.n322 VTAIL.n321 9.3005
R872 VTAIL.n347 VTAIL.n346 9.3005
R873 VTAIL.n345 VTAIL.n344 9.3005
R874 VTAIL.n326 VTAIL.n325 9.3005
R875 VTAIL.n339 VTAIL.n338 9.3005
R876 VTAIL.n337 VTAIL.n336 9.3005
R877 VTAIL.n330 VTAIL.n329 9.3005
R878 VTAIL.n742 VTAIL.n741 8.92171
R879 VTAIL.n757 VTAIL.n710 8.92171
R880 VTAIL.n788 VTAIL.n694 8.92171
R881 VTAIL.n50 VTAIL.n49 8.92171
R882 VTAIL.n65 VTAIL.n18 8.92171
R883 VTAIL.n96 VTAIL.n2 8.92171
R884 VTAIL.n148 VTAIL.n147 8.92171
R885 VTAIL.n163 VTAIL.n116 8.92171
R886 VTAIL.n194 VTAIL.n100 8.92171
R887 VTAIL.n248 VTAIL.n247 8.92171
R888 VTAIL.n263 VTAIL.n216 8.92171
R889 VTAIL.n294 VTAIL.n200 8.92171
R890 VTAIL.n690 VTAIL.n596 8.92171
R891 VTAIL.n661 VTAIL.n614 8.92171
R892 VTAIL.n646 VTAIL.n645 8.92171
R893 VTAIL.n590 VTAIL.n496 8.92171
R894 VTAIL.n561 VTAIL.n514 8.92171
R895 VTAIL.n546 VTAIL.n545 8.92171
R896 VTAIL.n492 VTAIL.n398 8.92171
R897 VTAIL.n463 VTAIL.n416 8.92171
R898 VTAIL.n448 VTAIL.n447 8.92171
R899 VTAIL.n392 VTAIL.n298 8.92171
R900 VTAIL.n363 VTAIL.n316 8.92171
R901 VTAIL.n348 VTAIL.n347 8.92171
R902 VTAIL.n745 VTAIL.n716 8.14595
R903 VTAIL.n754 VTAIL.n753 8.14595
R904 VTAIL.n53 VTAIL.n24 8.14595
R905 VTAIL.n62 VTAIL.n61 8.14595
R906 VTAIL.n151 VTAIL.n122 8.14595
R907 VTAIL.n160 VTAIL.n159 8.14595
R908 VTAIL.n251 VTAIL.n222 8.14595
R909 VTAIL.n260 VTAIL.n259 8.14595
R910 VTAIL.n658 VTAIL.n657 8.14595
R911 VTAIL.n649 VTAIL.n620 8.14595
R912 VTAIL.n558 VTAIL.n557 8.14595
R913 VTAIL.n549 VTAIL.n520 8.14595
R914 VTAIL.n460 VTAIL.n459 8.14595
R915 VTAIL.n451 VTAIL.n422 8.14595
R916 VTAIL.n360 VTAIL.n359 8.14595
R917 VTAIL.n351 VTAIL.n322 8.14595
R918 VTAIL.n746 VTAIL.n714 7.3702
R919 VTAIL.n750 VTAIL.n712 7.3702
R920 VTAIL.n54 VTAIL.n22 7.3702
R921 VTAIL.n58 VTAIL.n20 7.3702
R922 VTAIL.n152 VTAIL.n120 7.3702
R923 VTAIL.n156 VTAIL.n118 7.3702
R924 VTAIL.n252 VTAIL.n220 7.3702
R925 VTAIL.n256 VTAIL.n218 7.3702
R926 VTAIL.n654 VTAIL.n616 7.3702
R927 VTAIL.n650 VTAIL.n618 7.3702
R928 VTAIL.n554 VTAIL.n516 7.3702
R929 VTAIL.n550 VTAIL.n518 7.3702
R930 VTAIL.n456 VTAIL.n418 7.3702
R931 VTAIL.n452 VTAIL.n420 7.3702
R932 VTAIL.n356 VTAIL.n318 7.3702
R933 VTAIL.n352 VTAIL.n320 7.3702
R934 VTAIL.n749 VTAIL.n714 6.59444
R935 VTAIL.n750 VTAIL.n749 6.59444
R936 VTAIL.n57 VTAIL.n22 6.59444
R937 VTAIL.n58 VTAIL.n57 6.59444
R938 VTAIL.n155 VTAIL.n120 6.59444
R939 VTAIL.n156 VTAIL.n155 6.59444
R940 VTAIL.n255 VTAIL.n220 6.59444
R941 VTAIL.n256 VTAIL.n255 6.59444
R942 VTAIL.n654 VTAIL.n653 6.59444
R943 VTAIL.n653 VTAIL.n618 6.59444
R944 VTAIL.n554 VTAIL.n553 6.59444
R945 VTAIL.n553 VTAIL.n518 6.59444
R946 VTAIL.n456 VTAIL.n455 6.59444
R947 VTAIL.n455 VTAIL.n420 6.59444
R948 VTAIL.n356 VTAIL.n355 6.59444
R949 VTAIL.n355 VTAIL.n320 6.59444
R950 VTAIL.n746 VTAIL.n745 5.81868
R951 VTAIL.n753 VTAIL.n712 5.81868
R952 VTAIL.n54 VTAIL.n53 5.81868
R953 VTAIL.n61 VTAIL.n20 5.81868
R954 VTAIL.n152 VTAIL.n151 5.81868
R955 VTAIL.n159 VTAIL.n118 5.81868
R956 VTAIL.n252 VTAIL.n251 5.81868
R957 VTAIL.n259 VTAIL.n218 5.81868
R958 VTAIL.n657 VTAIL.n616 5.81868
R959 VTAIL.n650 VTAIL.n649 5.81868
R960 VTAIL.n557 VTAIL.n516 5.81868
R961 VTAIL.n550 VTAIL.n549 5.81868
R962 VTAIL.n459 VTAIL.n418 5.81868
R963 VTAIL.n452 VTAIL.n451 5.81868
R964 VTAIL.n359 VTAIL.n318 5.81868
R965 VTAIL.n352 VTAIL.n351 5.81868
R966 VTAIL.n742 VTAIL.n716 5.04292
R967 VTAIL.n754 VTAIL.n710 5.04292
R968 VTAIL.n790 VTAIL.n694 5.04292
R969 VTAIL.n50 VTAIL.n24 5.04292
R970 VTAIL.n62 VTAIL.n18 5.04292
R971 VTAIL.n98 VTAIL.n2 5.04292
R972 VTAIL.n148 VTAIL.n122 5.04292
R973 VTAIL.n160 VTAIL.n116 5.04292
R974 VTAIL.n196 VTAIL.n100 5.04292
R975 VTAIL.n248 VTAIL.n222 5.04292
R976 VTAIL.n260 VTAIL.n216 5.04292
R977 VTAIL.n296 VTAIL.n200 5.04292
R978 VTAIL.n692 VTAIL.n596 5.04292
R979 VTAIL.n658 VTAIL.n614 5.04292
R980 VTAIL.n646 VTAIL.n620 5.04292
R981 VTAIL.n592 VTAIL.n496 5.04292
R982 VTAIL.n558 VTAIL.n514 5.04292
R983 VTAIL.n546 VTAIL.n520 5.04292
R984 VTAIL.n494 VTAIL.n398 5.04292
R985 VTAIL.n460 VTAIL.n416 5.04292
R986 VTAIL.n448 VTAIL.n422 5.04292
R987 VTAIL.n394 VTAIL.n298 5.04292
R988 VTAIL.n360 VTAIL.n316 5.04292
R989 VTAIL.n348 VTAIL.n322 5.04292
R990 VTAIL.n741 VTAIL.n718 4.26717
R991 VTAIL.n758 VTAIL.n757 4.26717
R992 VTAIL.n788 VTAIL.n787 4.26717
R993 VTAIL.n49 VTAIL.n26 4.26717
R994 VTAIL.n66 VTAIL.n65 4.26717
R995 VTAIL.n96 VTAIL.n95 4.26717
R996 VTAIL.n147 VTAIL.n124 4.26717
R997 VTAIL.n164 VTAIL.n163 4.26717
R998 VTAIL.n194 VTAIL.n193 4.26717
R999 VTAIL.n247 VTAIL.n224 4.26717
R1000 VTAIL.n264 VTAIL.n263 4.26717
R1001 VTAIL.n294 VTAIL.n293 4.26717
R1002 VTAIL.n690 VTAIL.n689 4.26717
R1003 VTAIL.n662 VTAIL.n661 4.26717
R1004 VTAIL.n645 VTAIL.n622 4.26717
R1005 VTAIL.n590 VTAIL.n589 4.26717
R1006 VTAIL.n562 VTAIL.n561 4.26717
R1007 VTAIL.n545 VTAIL.n522 4.26717
R1008 VTAIL.n492 VTAIL.n491 4.26717
R1009 VTAIL.n464 VTAIL.n463 4.26717
R1010 VTAIL.n447 VTAIL.n424 4.26717
R1011 VTAIL.n392 VTAIL.n391 4.26717
R1012 VTAIL.n364 VTAIL.n363 4.26717
R1013 VTAIL.n347 VTAIL.n324 4.26717
R1014 VTAIL.n725 VTAIL.n723 3.70982
R1015 VTAIL.n33 VTAIL.n31 3.70982
R1016 VTAIL.n131 VTAIL.n129 3.70982
R1017 VTAIL.n231 VTAIL.n229 3.70982
R1018 VTAIL.n629 VTAIL.n627 3.70982
R1019 VTAIL.n529 VTAIL.n527 3.70982
R1020 VTAIL.n431 VTAIL.n429 3.70982
R1021 VTAIL.n331 VTAIL.n329 3.70982
R1022 VTAIL.n397 VTAIL.n395 3.63843
R1023 VTAIL.n495 VTAIL.n397 3.63843
R1024 VTAIL.n595 VTAIL.n593 3.63843
R1025 VTAIL.n693 VTAIL.n595 3.63843
R1026 VTAIL.n297 VTAIL.n199 3.63843
R1027 VTAIL.n199 VTAIL.n197 3.63843
R1028 VTAIL.n99 VTAIL.n1 3.63843
R1029 VTAIL VTAIL.n791 3.58024
R1030 VTAIL.n738 VTAIL.n737 3.49141
R1031 VTAIL.n761 VTAIL.n708 3.49141
R1032 VTAIL.n784 VTAIL.n696 3.49141
R1033 VTAIL.n46 VTAIL.n45 3.49141
R1034 VTAIL.n69 VTAIL.n16 3.49141
R1035 VTAIL.n92 VTAIL.n4 3.49141
R1036 VTAIL.n144 VTAIL.n143 3.49141
R1037 VTAIL.n167 VTAIL.n114 3.49141
R1038 VTAIL.n190 VTAIL.n102 3.49141
R1039 VTAIL.n244 VTAIL.n243 3.49141
R1040 VTAIL.n267 VTAIL.n214 3.49141
R1041 VTAIL.n290 VTAIL.n202 3.49141
R1042 VTAIL.n686 VTAIL.n598 3.49141
R1043 VTAIL.n665 VTAIL.n612 3.49141
R1044 VTAIL.n642 VTAIL.n641 3.49141
R1045 VTAIL.n586 VTAIL.n498 3.49141
R1046 VTAIL.n565 VTAIL.n512 3.49141
R1047 VTAIL.n542 VTAIL.n541 3.49141
R1048 VTAIL.n488 VTAIL.n400 3.49141
R1049 VTAIL.n467 VTAIL.n414 3.49141
R1050 VTAIL.n444 VTAIL.n443 3.49141
R1051 VTAIL.n388 VTAIL.n300 3.49141
R1052 VTAIL.n367 VTAIL.n314 3.49141
R1053 VTAIL.n344 VTAIL.n343 3.49141
R1054 VTAIL.n734 VTAIL.n720 2.71565
R1055 VTAIL.n762 VTAIL.n706 2.71565
R1056 VTAIL.n783 VTAIL.n698 2.71565
R1057 VTAIL.n42 VTAIL.n28 2.71565
R1058 VTAIL.n70 VTAIL.n14 2.71565
R1059 VTAIL.n91 VTAIL.n6 2.71565
R1060 VTAIL.n140 VTAIL.n126 2.71565
R1061 VTAIL.n168 VTAIL.n112 2.71565
R1062 VTAIL.n189 VTAIL.n104 2.71565
R1063 VTAIL.n240 VTAIL.n226 2.71565
R1064 VTAIL.n268 VTAIL.n212 2.71565
R1065 VTAIL.n289 VTAIL.n204 2.71565
R1066 VTAIL.n685 VTAIL.n600 2.71565
R1067 VTAIL.n666 VTAIL.n610 2.71565
R1068 VTAIL.n638 VTAIL.n624 2.71565
R1069 VTAIL.n585 VTAIL.n500 2.71565
R1070 VTAIL.n566 VTAIL.n510 2.71565
R1071 VTAIL.n538 VTAIL.n524 2.71565
R1072 VTAIL.n487 VTAIL.n402 2.71565
R1073 VTAIL.n468 VTAIL.n412 2.71565
R1074 VTAIL.n440 VTAIL.n426 2.71565
R1075 VTAIL.n387 VTAIL.n302 2.71565
R1076 VTAIL.n368 VTAIL.n312 2.71565
R1077 VTAIL.n340 VTAIL.n326 2.71565
R1078 VTAIL.n733 VTAIL.n722 1.93989
R1079 VTAIL.n767 VTAIL.n765 1.93989
R1080 VTAIL.n780 VTAIL.n779 1.93989
R1081 VTAIL.n41 VTAIL.n30 1.93989
R1082 VTAIL.n75 VTAIL.n73 1.93989
R1083 VTAIL.n88 VTAIL.n87 1.93989
R1084 VTAIL.n139 VTAIL.n128 1.93989
R1085 VTAIL.n173 VTAIL.n171 1.93989
R1086 VTAIL.n186 VTAIL.n185 1.93989
R1087 VTAIL.n239 VTAIL.n228 1.93989
R1088 VTAIL.n273 VTAIL.n271 1.93989
R1089 VTAIL.n286 VTAIL.n285 1.93989
R1090 VTAIL.n682 VTAIL.n681 1.93989
R1091 VTAIL.n670 VTAIL.n669 1.93989
R1092 VTAIL.n637 VTAIL.n626 1.93989
R1093 VTAIL.n582 VTAIL.n581 1.93989
R1094 VTAIL.n570 VTAIL.n569 1.93989
R1095 VTAIL.n537 VTAIL.n526 1.93989
R1096 VTAIL.n484 VTAIL.n483 1.93989
R1097 VTAIL.n472 VTAIL.n471 1.93989
R1098 VTAIL.n439 VTAIL.n428 1.93989
R1099 VTAIL.n384 VTAIL.n383 1.93989
R1100 VTAIL.n372 VTAIL.n371 1.93989
R1101 VTAIL.n339 VTAIL.n328 1.93989
R1102 VTAIL.n0 VTAIL.t9 1.84633
R1103 VTAIL.n0 VTAIL.t14 1.84633
R1104 VTAIL.n198 VTAIL.t0 1.84633
R1105 VTAIL.n198 VTAIL.t6 1.84633
R1106 VTAIL.n594 VTAIL.t1 1.84633
R1107 VTAIL.n594 VTAIL.t4 1.84633
R1108 VTAIL.n396 VTAIL.t13 1.84633
R1109 VTAIL.n396 VTAIL.t10 1.84633
R1110 VTAIL.n730 VTAIL.n729 1.16414
R1111 VTAIL.n766 VTAIL.n704 1.16414
R1112 VTAIL.n776 VTAIL.n700 1.16414
R1113 VTAIL.n38 VTAIL.n37 1.16414
R1114 VTAIL.n74 VTAIL.n12 1.16414
R1115 VTAIL.n84 VTAIL.n8 1.16414
R1116 VTAIL.n136 VTAIL.n135 1.16414
R1117 VTAIL.n172 VTAIL.n110 1.16414
R1118 VTAIL.n182 VTAIL.n106 1.16414
R1119 VTAIL.n236 VTAIL.n235 1.16414
R1120 VTAIL.n272 VTAIL.n210 1.16414
R1121 VTAIL.n282 VTAIL.n206 1.16414
R1122 VTAIL.n678 VTAIL.n602 1.16414
R1123 VTAIL.n673 VTAIL.n607 1.16414
R1124 VTAIL.n634 VTAIL.n633 1.16414
R1125 VTAIL.n578 VTAIL.n502 1.16414
R1126 VTAIL.n573 VTAIL.n507 1.16414
R1127 VTAIL.n534 VTAIL.n533 1.16414
R1128 VTAIL.n480 VTAIL.n404 1.16414
R1129 VTAIL.n475 VTAIL.n409 1.16414
R1130 VTAIL.n436 VTAIL.n435 1.16414
R1131 VTAIL.n380 VTAIL.n304 1.16414
R1132 VTAIL.n375 VTAIL.n309 1.16414
R1133 VTAIL.n336 VTAIL.n335 1.16414
R1134 VTAIL.n593 VTAIL.n495 0.470328
R1135 VTAIL.n197 VTAIL.n99 0.470328
R1136 VTAIL.n726 VTAIL.n724 0.388379
R1137 VTAIL.n772 VTAIL.n771 0.388379
R1138 VTAIL.n775 VTAIL.n702 0.388379
R1139 VTAIL.n34 VTAIL.n32 0.388379
R1140 VTAIL.n80 VTAIL.n79 0.388379
R1141 VTAIL.n83 VTAIL.n10 0.388379
R1142 VTAIL.n132 VTAIL.n130 0.388379
R1143 VTAIL.n178 VTAIL.n177 0.388379
R1144 VTAIL.n181 VTAIL.n108 0.388379
R1145 VTAIL.n232 VTAIL.n230 0.388379
R1146 VTAIL.n278 VTAIL.n277 0.388379
R1147 VTAIL.n281 VTAIL.n208 0.388379
R1148 VTAIL.n677 VTAIL.n604 0.388379
R1149 VTAIL.n674 VTAIL.n606 0.388379
R1150 VTAIL.n630 VTAIL.n628 0.388379
R1151 VTAIL.n577 VTAIL.n504 0.388379
R1152 VTAIL.n574 VTAIL.n506 0.388379
R1153 VTAIL.n530 VTAIL.n528 0.388379
R1154 VTAIL.n479 VTAIL.n406 0.388379
R1155 VTAIL.n476 VTAIL.n408 0.388379
R1156 VTAIL.n432 VTAIL.n430 0.388379
R1157 VTAIL.n379 VTAIL.n306 0.388379
R1158 VTAIL.n376 VTAIL.n308 0.388379
R1159 VTAIL.n332 VTAIL.n330 0.388379
R1160 VTAIL.n731 VTAIL.n723 0.155672
R1161 VTAIL.n732 VTAIL.n731 0.155672
R1162 VTAIL.n732 VTAIL.n719 0.155672
R1163 VTAIL.n739 VTAIL.n719 0.155672
R1164 VTAIL.n740 VTAIL.n739 0.155672
R1165 VTAIL.n740 VTAIL.n715 0.155672
R1166 VTAIL.n747 VTAIL.n715 0.155672
R1167 VTAIL.n748 VTAIL.n747 0.155672
R1168 VTAIL.n748 VTAIL.n711 0.155672
R1169 VTAIL.n755 VTAIL.n711 0.155672
R1170 VTAIL.n756 VTAIL.n755 0.155672
R1171 VTAIL.n756 VTAIL.n707 0.155672
R1172 VTAIL.n763 VTAIL.n707 0.155672
R1173 VTAIL.n764 VTAIL.n763 0.155672
R1174 VTAIL.n764 VTAIL.n703 0.155672
R1175 VTAIL.n773 VTAIL.n703 0.155672
R1176 VTAIL.n774 VTAIL.n773 0.155672
R1177 VTAIL.n774 VTAIL.n699 0.155672
R1178 VTAIL.n781 VTAIL.n699 0.155672
R1179 VTAIL.n782 VTAIL.n781 0.155672
R1180 VTAIL.n782 VTAIL.n695 0.155672
R1181 VTAIL.n789 VTAIL.n695 0.155672
R1182 VTAIL.n39 VTAIL.n31 0.155672
R1183 VTAIL.n40 VTAIL.n39 0.155672
R1184 VTAIL.n40 VTAIL.n27 0.155672
R1185 VTAIL.n47 VTAIL.n27 0.155672
R1186 VTAIL.n48 VTAIL.n47 0.155672
R1187 VTAIL.n48 VTAIL.n23 0.155672
R1188 VTAIL.n55 VTAIL.n23 0.155672
R1189 VTAIL.n56 VTAIL.n55 0.155672
R1190 VTAIL.n56 VTAIL.n19 0.155672
R1191 VTAIL.n63 VTAIL.n19 0.155672
R1192 VTAIL.n64 VTAIL.n63 0.155672
R1193 VTAIL.n64 VTAIL.n15 0.155672
R1194 VTAIL.n71 VTAIL.n15 0.155672
R1195 VTAIL.n72 VTAIL.n71 0.155672
R1196 VTAIL.n72 VTAIL.n11 0.155672
R1197 VTAIL.n81 VTAIL.n11 0.155672
R1198 VTAIL.n82 VTAIL.n81 0.155672
R1199 VTAIL.n82 VTAIL.n7 0.155672
R1200 VTAIL.n89 VTAIL.n7 0.155672
R1201 VTAIL.n90 VTAIL.n89 0.155672
R1202 VTAIL.n90 VTAIL.n3 0.155672
R1203 VTAIL.n97 VTAIL.n3 0.155672
R1204 VTAIL.n137 VTAIL.n129 0.155672
R1205 VTAIL.n138 VTAIL.n137 0.155672
R1206 VTAIL.n138 VTAIL.n125 0.155672
R1207 VTAIL.n145 VTAIL.n125 0.155672
R1208 VTAIL.n146 VTAIL.n145 0.155672
R1209 VTAIL.n146 VTAIL.n121 0.155672
R1210 VTAIL.n153 VTAIL.n121 0.155672
R1211 VTAIL.n154 VTAIL.n153 0.155672
R1212 VTAIL.n154 VTAIL.n117 0.155672
R1213 VTAIL.n161 VTAIL.n117 0.155672
R1214 VTAIL.n162 VTAIL.n161 0.155672
R1215 VTAIL.n162 VTAIL.n113 0.155672
R1216 VTAIL.n169 VTAIL.n113 0.155672
R1217 VTAIL.n170 VTAIL.n169 0.155672
R1218 VTAIL.n170 VTAIL.n109 0.155672
R1219 VTAIL.n179 VTAIL.n109 0.155672
R1220 VTAIL.n180 VTAIL.n179 0.155672
R1221 VTAIL.n180 VTAIL.n105 0.155672
R1222 VTAIL.n187 VTAIL.n105 0.155672
R1223 VTAIL.n188 VTAIL.n187 0.155672
R1224 VTAIL.n188 VTAIL.n101 0.155672
R1225 VTAIL.n195 VTAIL.n101 0.155672
R1226 VTAIL.n237 VTAIL.n229 0.155672
R1227 VTAIL.n238 VTAIL.n237 0.155672
R1228 VTAIL.n238 VTAIL.n225 0.155672
R1229 VTAIL.n245 VTAIL.n225 0.155672
R1230 VTAIL.n246 VTAIL.n245 0.155672
R1231 VTAIL.n246 VTAIL.n221 0.155672
R1232 VTAIL.n253 VTAIL.n221 0.155672
R1233 VTAIL.n254 VTAIL.n253 0.155672
R1234 VTAIL.n254 VTAIL.n217 0.155672
R1235 VTAIL.n261 VTAIL.n217 0.155672
R1236 VTAIL.n262 VTAIL.n261 0.155672
R1237 VTAIL.n262 VTAIL.n213 0.155672
R1238 VTAIL.n269 VTAIL.n213 0.155672
R1239 VTAIL.n270 VTAIL.n269 0.155672
R1240 VTAIL.n270 VTAIL.n209 0.155672
R1241 VTAIL.n279 VTAIL.n209 0.155672
R1242 VTAIL.n280 VTAIL.n279 0.155672
R1243 VTAIL.n280 VTAIL.n205 0.155672
R1244 VTAIL.n287 VTAIL.n205 0.155672
R1245 VTAIL.n288 VTAIL.n287 0.155672
R1246 VTAIL.n288 VTAIL.n201 0.155672
R1247 VTAIL.n295 VTAIL.n201 0.155672
R1248 VTAIL.n691 VTAIL.n597 0.155672
R1249 VTAIL.n684 VTAIL.n597 0.155672
R1250 VTAIL.n684 VTAIL.n683 0.155672
R1251 VTAIL.n683 VTAIL.n601 0.155672
R1252 VTAIL.n676 VTAIL.n601 0.155672
R1253 VTAIL.n676 VTAIL.n675 0.155672
R1254 VTAIL.n675 VTAIL.n605 0.155672
R1255 VTAIL.n668 VTAIL.n605 0.155672
R1256 VTAIL.n668 VTAIL.n667 0.155672
R1257 VTAIL.n667 VTAIL.n611 0.155672
R1258 VTAIL.n660 VTAIL.n611 0.155672
R1259 VTAIL.n660 VTAIL.n659 0.155672
R1260 VTAIL.n659 VTAIL.n615 0.155672
R1261 VTAIL.n652 VTAIL.n615 0.155672
R1262 VTAIL.n652 VTAIL.n651 0.155672
R1263 VTAIL.n651 VTAIL.n619 0.155672
R1264 VTAIL.n644 VTAIL.n619 0.155672
R1265 VTAIL.n644 VTAIL.n643 0.155672
R1266 VTAIL.n643 VTAIL.n623 0.155672
R1267 VTAIL.n636 VTAIL.n623 0.155672
R1268 VTAIL.n636 VTAIL.n635 0.155672
R1269 VTAIL.n635 VTAIL.n627 0.155672
R1270 VTAIL.n591 VTAIL.n497 0.155672
R1271 VTAIL.n584 VTAIL.n497 0.155672
R1272 VTAIL.n584 VTAIL.n583 0.155672
R1273 VTAIL.n583 VTAIL.n501 0.155672
R1274 VTAIL.n576 VTAIL.n501 0.155672
R1275 VTAIL.n576 VTAIL.n575 0.155672
R1276 VTAIL.n575 VTAIL.n505 0.155672
R1277 VTAIL.n568 VTAIL.n505 0.155672
R1278 VTAIL.n568 VTAIL.n567 0.155672
R1279 VTAIL.n567 VTAIL.n511 0.155672
R1280 VTAIL.n560 VTAIL.n511 0.155672
R1281 VTAIL.n560 VTAIL.n559 0.155672
R1282 VTAIL.n559 VTAIL.n515 0.155672
R1283 VTAIL.n552 VTAIL.n515 0.155672
R1284 VTAIL.n552 VTAIL.n551 0.155672
R1285 VTAIL.n551 VTAIL.n519 0.155672
R1286 VTAIL.n544 VTAIL.n519 0.155672
R1287 VTAIL.n544 VTAIL.n543 0.155672
R1288 VTAIL.n543 VTAIL.n523 0.155672
R1289 VTAIL.n536 VTAIL.n523 0.155672
R1290 VTAIL.n536 VTAIL.n535 0.155672
R1291 VTAIL.n535 VTAIL.n527 0.155672
R1292 VTAIL.n493 VTAIL.n399 0.155672
R1293 VTAIL.n486 VTAIL.n399 0.155672
R1294 VTAIL.n486 VTAIL.n485 0.155672
R1295 VTAIL.n485 VTAIL.n403 0.155672
R1296 VTAIL.n478 VTAIL.n403 0.155672
R1297 VTAIL.n478 VTAIL.n477 0.155672
R1298 VTAIL.n477 VTAIL.n407 0.155672
R1299 VTAIL.n470 VTAIL.n407 0.155672
R1300 VTAIL.n470 VTAIL.n469 0.155672
R1301 VTAIL.n469 VTAIL.n413 0.155672
R1302 VTAIL.n462 VTAIL.n413 0.155672
R1303 VTAIL.n462 VTAIL.n461 0.155672
R1304 VTAIL.n461 VTAIL.n417 0.155672
R1305 VTAIL.n454 VTAIL.n417 0.155672
R1306 VTAIL.n454 VTAIL.n453 0.155672
R1307 VTAIL.n453 VTAIL.n421 0.155672
R1308 VTAIL.n446 VTAIL.n421 0.155672
R1309 VTAIL.n446 VTAIL.n445 0.155672
R1310 VTAIL.n445 VTAIL.n425 0.155672
R1311 VTAIL.n438 VTAIL.n425 0.155672
R1312 VTAIL.n438 VTAIL.n437 0.155672
R1313 VTAIL.n437 VTAIL.n429 0.155672
R1314 VTAIL.n393 VTAIL.n299 0.155672
R1315 VTAIL.n386 VTAIL.n299 0.155672
R1316 VTAIL.n386 VTAIL.n385 0.155672
R1317 VTAIL.n385 VTAIL.n303 0.155672
R1318 VTAIL.n378 VTAIL.n303 0.155672
R1319 VTAIL.n378 VTAIL.n377 0.155672
R1320 VTAIL.n377 VTAIL.n307 0.155672
R1321 VTAIL.n370 VTAIL.n307 0.155672
R1322 VTAIL.n370 VTAIL.n369 0.155672
R1323 VTAIL.n369 VTAIL.n313 0.155672
R1324 VTAIL.n362 VTAIL.n313 0.155672
R1325 VTAIL.n362 VTAIL.n361 0.155672
R1326 VTAIL.n361 VTAIL.n317 0.155672
R1327 VTAIL.n354 VTAIL.n317 0.155672
R1328 VTAIL.n354 VTAIL.n353 0.155672
R1329 VTAIL.n353 VTAIL.n321 0.155672
R1330 VTAIL.n346 VTAIL.n321 0.155672
R1331 VTAIL.n346 VTAIL.n345 0.155672
R1332 VTAIL.n345 VTAIL.n325 0.155672
R1333 VTAIL.n338 VTAIL.n325 0.155672
R1334 VTAIL.n338 VTAIL.n337 0.155672
R1335 VTAIL.n337 VTAIL.n329 0.155672
R1336 VTAIL VTAIL.n1 0.0586897
R1337 VP.n26 VP.n25 161.3
R1338 VP.n27 VP.n22 161.3
R1339 VP.n29 VP.n28 161.3
R1340 VP.n30 VP.n21 161.3
R1341 VP.n32 VP.n31 161.3
R1342 VP.n33 VP.n20 161.3
R1343 VP.n35 VP.n34 161.3
R1344 VP.n36 VP.n19 161.3
R1345 VP.n39 VP.n38 161.3
R1346 VP.n40 VP.n18 161.3
R1347 VP.n42 VP.n41 161.3
R1348 VP.n43 VP.n17 161.3
R1349 VP.n45 VP.n44 161.3
R1350 VP.n46 VP.n16 161.3
R1351 VP.n48 VP.n47 161.3
R1352 VP.n49 VP.n15 161.3
R1353 VP.n51 VP.n50 161.3
R1354 VP.n95 VP.n94 161.3
R1355 VP.n93 VP.n1 161.3
R1356 VP.n92 VP.n91 161.3
R1357 VP.n90 VP.n2 161.3
R1358 VP.n89 VP.n88 161.3
R1359 VP.n87 VP.n3 161.3
R1360 VP.n86 VP.n85 161.3
R1361 VP.n84 VP.n4 161.3
R1362 VP.n83 VP.n82 161.3
R1363 VP.n80 VP.n5 161.3
R1364 VP.n79 VP.n78 161.3
R1365 VP.n77 VP.n6 161.3
R1366 VP.n76 VP.n75 161.3
R1367 VP.n74 VP.n7 161.3
R1368 VP.n73 VP.n72 161.3
R1369 VP.n71 VP.n8 161.3
R1370 VP.n70 VP.n69 161.3
R1371 VP.n67 VP.n9 161.3
R1372 VP.n66 VP.n65 161.3
R1373 VP.n64 VP.n10 161.3
R1374 VP.n63 VP.n62 161.3
R1375 VP.n61 VP.n11 161.3
R1376 VP.n60 VP.n59 161.3
R1377 VP.n58 VP.n12 161.3
R1378 VP.n57 VP.n56 161.3
R1379 VP.n55 VP.n13 161.3
R1380 VP.n23 VP.t0 142.212
R1381 VP.n54 VP.t2 109.102
R1382 VP.n68 VP.t4 109.102
R1383 VP.n81 VP.t3 109.102
R1384 VP.n0 VP.t1 109.102
R1385 VP.n14 VP.t6 109.102
R1386 VP.n37 VP.t7 109.102
R1387 VP.n24 VP.t5 109.102
R1388 VP.n54 VP.n53 86.1527
R1389 VP.n96 VP.n0 86.1527
R1390 VP.n52 VP.n14 86.1527
R1391 VP.n53 VP.n52 61.2721
R1392 VP.n24 VP.n23 57.4697
R1393 VP.n75 VP.n74 56.5193
R1394 VP.n31 VP.n30 56.5193
R1395 VP.n62 VP.n61 43.4072
R1396 VP.n88 VP.n87 43.4072
R1397 VP.n44 VP.n43 43.4072
R1398 VP.n61 VP.n60 37.5796
R1399 VP.n88 VP.n2 37.5796
R1400 VP.n44 VP.n16 37.5796
R1401 VP.n56 VP.n55 24.4675
R1402 VP.n56 VP.n12 24.4675
R1403 VP.n60 VP.n12 24.4675
R1404 VP.n62 VP.n10 24.4675
R1405 VP.n66 VP.n10 24.4675
R1406 VP.n67 VP.n66 24.4675
R1407 VP.n69 VP.n8 24.4675
R1408 VP.n73 VP.n8 24.4675
R1409 VP.n74 VP.n73 24.4675
R1410 VP.n75 VP.n6 24.4675
R1411 VP.n79 VP.n6 24.4675
R1412 VP.n80 VP.n79 24.4675
R1413 VP.n82 VP.n4 24.4675
R1414 VP.n86 VP.n4 24.4675
R1415 VP.n87 VP.n86 24.4675
R1416 VP.n92 VP.n2 24.4675
R1417 VP.n93 VP.n92 24.4675
R1418 VP.n94 VP.n93 24.4675
R1419 VP.n48 VP.n16 24.4675
R1420 VP.n49 VP.n48 24.4675
R1421 VP.n50 VP.n49 24.4675
R1422 VP.n31 VP.n20 24.4675
R1423 VP.n35 VP.n20 24.4675
R1424 VP.n36 VP.n35 24.4675
R1425 VP.n38 VP.n18 24.4675
R1426 VP.n42 VP.n18 24.4675
R1427 VP.n43 VP.n42 24.4675
R1428 VP.n25 VP.n22 24.4675
R1429 VP.n29 VP.n22 24.4675
R1430 VP.n30 VP.n29 24.4675
R1431 VP.n69 VP.n68 17.6167
R1432 VP.n81 VP.n80 17.6167
R1433 VP.n37 VP.n36 17.6167
R1434 VP.n25 VP.n24 17.6167
R1435 VP.n68 VP.n67 6.85126
R1436 VP.n82 VP.n81 6.85126
R1437 VP.n38 VP.n37 6.85126
R1438 VP.n55 VP.n54 3.91522
R1439 VP.n94 VP.n0 3.91522
R1440 VP.n50 VP.n14 3.91522
R1441 VP.n26 VP.n23 2.44108
R1442 VP.n52 VP.n51 0.354971
R1443 VP.n53 VP.n13 0.354971
R1444 VP.n96 VP.n95 0.354971
R1445 VP VP.n96 0.26696
R1446 VP.n27 VP.n26 0.189894
R1447 VP.n28 VP.n27 0.189894
R1448 VP.n28 VP.n21 0.189894
R1449 VP.n32 VP.n21 0.189894
R1450 VP.n33 VP.n32 0.189894
R1451 VP.n34 VP.n33 0.189894
R1452 VP.n34 VP.n19 0.189894
R1453 VP.n39 VP.n19 0.189894
R1454 VP.n40 VP.n39 0.189894
R1455 VP.n41 VP.n40 0.189894
R1456 VP.n41 VP.n17 0.189894
R1457 VP.n45 VP.n17 0.189894
R1458 VP.n46 VP.n45 0.189894
R1459 VP.n47 VP.n46 0.189894
R1460 VP.n47 VP.n15 0.189894
R1461 VP.n51 VP.n15 0.189894
R1462 VP.n57 VP.n13 0.189894
R1463 VP.n58 VP.n57 0.189894
R1464 VP.n59 VP.n58 0.189894
R1465 VP.n59 VP.n11 0.189894
R1466 VP.n63 VP.n11 0.189894
R1467 VP.n64 VP.n63 0.189894
R1468 VP.n65 VP.n64 0.189894
R1469 VP.n65 VP.n9 0.189894
R1470 VP.n70 VP.n9 0.189894
R1471 VP.n71 VP.n70 0.189894
R1472 VP.n72 VP.n71 0.189894
R1473 VP.n72 VP.n7 0.189894
R1474 VP.n76 VP.n7 0.189894
R1475 VP.n77 VP.n76 0.189894
R1476 VP.n78 VP.n77 0.189894
R1477 VP.n78 VP.n5 0.189894
R1478 VP.n83 VP.n5 0.189894
R1479 VP.n84 VP.n83 0.189894
R1480 VP.n85 VP.n84 0.189894
R1481 VP.n85 VP.n3 0.189894
R1482 VP.n89 VP.n3 0.189894
R1483 VP.n90 VP.n89 0.189894
R1484 VP.n91 VP.n90 0.189894
R1485 VP.n91 VP.n1 0.189894
R1486 VP.n95 VP.n1 0.189894
R1487 VDD1 VDD1.n0 72.6448
R1488 VDD1.n3 VDD1.n2 72.5311
R1489 VDD1.n3 VDD1.n1 72.5311
R1490 VDD1.n5 VDD1.n4 70.7675
R1491 VDD1.n5 VDD1.n3 55.85
R1492 VDD1.n4 VDD1.t0 1.84633
R1493 VDD1.n4 VDD1.t1 1.84633
R1494 VDD1.n0 VDD1.t7 1.84633
R1495 VDD1.n0 VDD1.t2 1.84633
R1496 VDD1.n2 VDD1.t4 1.84633
R1497 VDD1.n2 VDD1.t6 1.84633
R1498 VDD1.n1 VDD1.t5 1.84633
R1499 VDD1.n1 VDD1.t3 1.84633
R1500 VDD1 VDD1.n5 1.76128
R1501 B.n783 B.n104 585
R1502 B.n785 B.n784 585
R1503 B.n786 B.n103 585
R1504 B.n788 B.n787 585
R1505 B.n789 B.n102 585
R1506 B.n791 B.n790 585
R1507 B.n792 B.n101 585
R1508 B.n794 B.n793 585
R1509 B.n795 B.n100 585
R1510 B.n797 B.n796 585
R1511 B.n798 B.n99 585
R1512 B.n800 B.n799 585
R1513 B.n801 B.n98 585
R1514 B.n803 B.n802 585
R1515 B.n804 B.n97 585
R1516 B.n806 B.n805 585
R1517 B.n807 B.n96 585
R1518 B.n809 B.n808 585
R1519 B.n810 B.n95 585
R1520 B.n812 B.n811 585
R1521 B.n813 B.n94 585
R1522 B.n815 B.n814 585
R1523 B.n816 B.n93 585
R1524 B.n818 B.n817 585
R1525 B.n819 B.n92 585
R1526 B.n821 B.n820 585
R1527 B.n822 B.n91 585
R1528 B.n824 B.n823 585
R1529 B.n825 B.n90 585
R1530 B.n827 B.n826 585
R1531 B.n828 B.n89 585
R1532 B.n830 B.n829 585
R1533 B.n831 B.n88 585
R1534 B.n833 B.n832 585
R1535 B.n834 B.n87 585
R1536 B.n836 B.n835 585
R1537 B.n837 B.n86 585
R1538 B.n839 B.n838 585
R1539 B.n840 B.n85 585
R1540 B.n842 B.n841 585
R1541 B.n843 B.n84 585
R1542 B.n845 B.n844 585
R1543 B.n846 B.n83 585
R1544 B.n848 B.n847 585
R1545 B.n849 B.n82 585
R1546 B.n851 B.n850 585
R1547 B.n852 B.n81 585
R1548 B.n854 B.n853 585
R1549 B.n855 B.n80 585
R1550 B.n857 B.n856 585
R1551 B.n858 B.n79 585
R1552 B.n860 B.n859 585
R1553 B.n861 B.n78 585
R1554 B.n863 B.n862 585
R1555 B.n864 B.n77 585
R1556 B.n866 B.n865 585
R1557 B.n867 B.n76 585
R1558 B.n869 B.n868 585
R1559 B.n871 B.n73 585
R1560 B.n873 B.n872 585
R1561 B.n874 B.n72 585
R1562 B.n876 B.n875 585
R1563 B.n877 B.n71 585
R1564 B.n879 B.n878 585
R1565 B.n880 B.n70 585
R1566 B.n882 B.n881 585
R1567 B.n883 B.n69 585
R1568 B.n885 B.n884 585
R1569 B.n887 B.n886 585
R1570 B.n888 B.n65 585
R1571 B.n890 B.n889 585
R1572 B.n891 B.n64 585
R1573 B.n893 B.n892 585
R1574 B.n894 B.n63 585
R1575 B.n896 B.n895 585
R1576 B.n897 B.n62 585
R1577 B.n899 B.n898 585
R1578 B.n900 B.n61 585
R1579 B.n902 B.n901 585
R1580 B.n903 B.n60 585
R1581 B.n905 B.n904 585
R1582 B.n906 B.n59 585
R1583 B.n908 B.n907 585
R1584 B.n909 B.n58 585
R1585 B.n911 B.n910 585
R1586 B.n912 B.n57 585
R1587 B.n914 B.n913 585
R1588 B.n915 B.n56 585
R1589 B.n917 B.n916 585
R1590 B.n918 B.n55 585
R1591 B.n920 B.n919 585
R1592 B.n921 B.n54 585
R1593 B.n923 B.n922 585
R1594 B.n924 B.n53 585
R1595 B.n926 B.n925 585
R1596 B.n927 B.n52 585
R1597 B.n929 B.n928 585
R1598 B.n930 B.n51 585
R1599 B.n932 B.n931 585
R1600 B.n933 B.n50 585
R1601 B.n935 B.n934 585
R1602 B.n936 B.n49 585
R1603 B.n938 B.n937 585
R1604 B.n939 B.n48 585
R1605 B.n941 B.n940 585
R1606 B.n942 B.n47 585
R1607 B.n944 B.n943 585
R1608 B.n945 B.n46 585
R1609 B.n947 B.n946 585
R1610 B.n948 B.n45 585
R1611 B.n950 B.n949 585
R1612 B.n951 B.n44 585
R1613 B.n953 B.n952 585
R1614 B.n954 B.n43 585
R1615 B.n956 B.n955 585
R1616 B.n957 B.n42 585
R1617 B.n959 B.n958 585
R1618 B.n960 B.n41 585
R1619 B.n962 B.n961 585
R1620 B.n963 B.n40 585
R1621 B.n965 B.n964 585
R1622 B.n966 B.n39 585
R1623 B.n968 B.n967 585
R1624 B.n969 B.n38 585
R1625 B.n971 B.n970 585
R1626 B.n972 B.n37 585
R1627 B.n782 B.n781 585
R1628 B.n780 B.n105 585
R1629 B.n779 B.n778 585
R1630 B.n777 B.n106 585
R1631 B.n776 B.n775 585
R1632 B.n774 B.n107 585
R1633 B.n773 B.n772 585
R1634 B.n771 B.n108 585
R1635 B.n770 B.n769 585
R1636 B.n768 B.n109 585
R1637 B.n767 B.n766 585
R1638 B.n765 B.n110 585
R1639 B.n764 B.n763 585
R1640 B.n762 B.n111 585
R1641 B.n761 B.n760 585
R1642 B.n759 B.n112 585
R1643 B.n758 B.n757 585
R1644 B.n756 B.n113 585
R1645 B.n755 B.n754 585
R1646 B.n753 B.n114 585
R1647 B.n752 B.n751 585
R1648 B.n750 B.n115 585
R1649 B.n749 B.n748 585
R1650 B.n747 B.n116 585
R1651 B.n746 B.n745 585
R1652 B.n744 B.n117 585
R1653 B.n743 B.n742 585
R1654 B.n741 B.n118 585
R1655 B.n740 B.n739 585
R1656 B.n738 B.n119 585
R1657 B.n737 B.n736 585
R1658 B.n735 B.n120 585
R1659 B.n734 B.n733 585
R1660 B.n732 B.n121 585
R1661 B.n731 B.n730 585
R1662 B.n729 B.n122 585
R1663 B.n728 B.n727 585
R1664 B.n726 B.n123 585
R1665 B.n725 B.n724 585
R1666 B.n723 B.n124 585
R1667 B.n722 B.n721 585
R1668 B.n720 B.n125 585
R1669 B.n719 B.n718 585
R1670 B.n717 B.n126 585
R1671 B.n716 B.n715 585
R1672 B.n714 B.n127 585
R1673 B.n713 B.n712 585
R1674 B.n711 B.n128 585
R1675 B.n710 B.n709 585
R1676 B.n708 B.n129 585
R1677 B.n707 B.n706 585
R1678 B.n705 B.n130 585
R1679 B.n704 B.n703 585
R1680 B.n702 B.n131 585
R1681 B.n701 B.n700 585
R1682 B.n699 B.n132 585
R1683 B.n698 B.n697 585
R1684 B.n696 B.n133 585
R1685 B.n695 B.n694 585
R1686 B.n693 B.n134 585
R1687 B.n692 B.n691 585
R1688 B.n690 B.n135 585
R1689 B.n689 B.n688 585
R1690 B.n687 B.n136 585
R1691 B.n686 B.n685 585
R1692 B.n684 B.n137 585
R1693 B.n683 B.n682 585
R1694 B.n681 B.n138 585
R1695 B.n680 B.n679 585
R1696 B.n678 B.n139 585
R1697 B.n677 B.n676 585
R1698 B.n675 B.n140 585
R1699 B.n674 B.n673 585
R1700 B.n672 B.n141 585
R1701 B.n671 B.n670 585
R1702 B.n669 B.n142 585
R1703 B.n668 B.n667 585
R1704 B.n666 B.n143 585
R1705 B.n665 B.n664 585
R1706 B.n663 B.n144 585
R1707 B.n662 B.n661 585
R1708 B.n660 B.n145 585
R1709 B.n659 B.n658 585
R1710 B.n657 B.n146 585
R1711 B.n656 B.n655 585
R1712 B.n654 B.n147 585
R1713 B.n653 B.n652 585
R1714 B.n651 B.n148 585
R1715 B.n650 B.n649 585
R1716 B.n648 B.n149 585
R1717 B.n647 B.n646 585
R1718 B.n645 B.n150 585
R1719 B.n644 B.n643 585
R1720 B.n642 B.n151 585
R1721 B.n641 B.n640 585
R1722 B.n639 B.n152 585
R1723 B.n638 B.n637 585
R1724 B.n636 B.n153 585
R1725 B.n635 B.n634 585
R1726 B.n633 B.n154 585
R1727 B.n632 B.n631 585
R1728 B.n630 B.n155 585
R1729 B.n629 B.n628 585
R1730 B.n627 B.n156 585
R1731 B.n626 B.n625 585
R1732 B.n624 B.n157 585
R1733 B.n623 B.n622 585
R1734 B.n621 B.n158 585
R1735 B.n620 B.n619 585
R1736 B.n618 B.n159 585
R1737 B.n617 B.n616 585
R1738 B.n615 B.n160 585
R1739 B.n614 B.n613 585
R1740 B.n612 B.n161 585
R1741 B.n611 B.n610 585
R1742 B.n609 B.n162 585
R1743 B.n608 B.n607 585
R1744 B.n606 B.n163 585
R1745 B.n605 B.n604 585
R1746 B.n603 B.n164 585
R1747 B.n602 B.n601 585
R1748 B.n600 B.n165 585
R1749 B.n599 B.n598 585
R1750 B.n597 B.n166 585
R1751 B.n596 B.n595 585
R1752 B.n594 B.n167 585
R1753 B.n593 B.n592 585
R1754 B.n591 B.n168 585
R1755 B.n590 B.n589 585
R1756 B.n588 B.n169 585
R1757 B.n587 B.n586 585
R1758 B.n585 B.n170 585
R1759 B.n584 B.n583 585
R1760 B.n582 B.n171 585
R1761 B.n581 B.n580 585
R1762 B.n579 B.n172 585
R1763 B.n578 B.n577 585
R1764 B.n576 B.n173 585
R1765 B.n575 B.n574 585
R1766 B.n573 B.n174 585
R1767 B.n572 B.n571 585
R1768 B.n381 B.n242 585
R1769 B.n383 B.n382 585
R1770 B.n384 B.n241 585
R1771 B.n386 B.n385 585
R1772 B.n387 B.n240 585
R1773 B.n389 B.n388 585
R1774 B.n390 B.n239 585
R1775 B.n392 B.n391 585
R1776 B.n393 B.n238 585
R1777 B.n395 B.n394 585
R1778 B.n396 B.n237 585
R1779 B.n398 B.n397 585
R1780 B.n399 B.n236 585
R1781 B.n401 B.n400 585
R1782 B.n402 B.n235 585
R1783 B.n404 B.n403 585
R1784 B.n405 B.n234 585
R1785 B.n407 B.n406 585
R1786 B.n408 B.n233 585
R1787 B.n410 B.n409 585
R1788 B.n411 B.n232 585
R1789 B.n413 B.n412 585
R1790 B.n414 B.n231 585
R1791 B.n416 B.n415 585
R1792 B.n417 B.n230 585
R1793 B.n419 B.n418 585
R1794 B.n420 B.n229 585
R1795 B.n422 B.n421 585
R1796 B.n423 B.n228 585
R1797 B.n425 B.n424 585
R1798 B.n426 B.n227 585
R1799 B.n428 B.n427 585
R1800 B.n429 B.n226 585
R1801 B.n431 B.n430 585
R1802 B.n432 B.n225 585
R1803 B.n434 B.n433 585
R1804 B.n435 B.n224 585
R1805 B.n437 B.n436 585
R1806 B.n438 B.n223 585
R1807 B.n440 B.n439 585
R1808 B.n441 B.n222 585
R1809 B.n443 B.n442 585
R1810 B.n444 B.n221 585
R1811 B.n446 B.n445 585
R1812 B.n447 B.n220 585
R1813 B.n449 B.n448 585
R1814 B.n450 B.n219 585
R1815 B.n452 B.n451 585
R1816 B.n453 B.n218 585
R1817 B.n455 B.n454 585
R1818 B.n456 B.n217 585
R1819 B.n458 B.n457 585
R1820 B.n459 B.n216 585
R1821 B.n461 B.n460 585
R1822 B.n462 B.n215 585
R1823 B.n464 B.n463 585
R1824 B.n465 B.n214 585
R1825 B.n467 B.n466 585
R1826 B.n469 B.n211 585
R1827 B.n471 B.n470 585
R1828 B.n472 B.n210 585
R1829 B.n474 B.n473 585
R1830 B.n475 B.n209 585
R1831 B.n477 B.n476 585
R1832 B.n478 B.n208 585
R1833 B.n480 B.n479 585
R1834 B.n481 B.n207 585
R1835 B.n483 B.n482 585
R1836 B.n485 B.n484 585
R1837 B.n486 B.n203 585
R1838 B.n488 B.n487 585
R1839 B.n489 B.n202 585
R1840 B.n491 B.n490 585
R1841 B.n492 B.n201 585
R1842 B.n494 B.n493 585
R1843 B.n495 B.n200 585
R1844 B.n497 B.n496 585
R1845 B.n498 B.n199 585
R1846 B.n500 B.n499 585
R1847 B.n501 B.n198 585
R1848 B.n503 B.n502 585
R1849 B.n504 B.n197 585
R1850 B.n506 B.n505 585
R1851 B.n507 B.n196 585
R1852 B.n509 B.n508 585
R1853 B.n510 B.n195 585
R1854 B.n512 B.n511 585
R1855 B.n513 B.n194 585
R1856 B.n515 B.n514 585
R1857 B.n516 B.n193 585
R1858 B.n518 B.n517 585
R1859 B.n519 B.n192 585
R1860 B.n521 B.n520 585
R1861 B.n522 B.n191 585
R1862 B.n524 B.n523 585
R1863 B.n525 B.n190 585
R1864 B.n527 B.n526 585
R1865 B.n528 B.n189 585
R1866 B.n530 B.n529 585
R1867 B.n531 B.n188 585
R1868 B.n533 B.n532 585
R1869 B.n534 B.n187 585
R1870 B.n536 B.n535 585
R1871 B.n537 B.n186 585
R1872 B.n539 B.n538 585
R1873 B.n540 B.n185 585
R1874 B.n542 B.n541 585
R1875 B.n543 B.n184 585
R1876 B.n545 B.n544 585
R1877 B.n546 B.n183 585
R1878 B.n548 B.n547 585
R1879 B.n549 B.n182 585
R1880 B.n551 B.n550 585
R1881 B.n552 B.n181 585
R1882 B.n554 B.n553 585
R1883 B.n555 B.n180 585
R1884 B.n557 B.n556 585
R1885 B.n558 B.n179 585
R1886 B.n560 B.n559 585
R1887 B.n561 B.n178 585
R1888 B.n563 B.n562 585
R1889 B.n564 B.n177 585
R1890 B.n566 B.n565 585
R1891 B.n567 B.n176 585
R1892 B.n569 B.n568 585
R1893 B.n570 B.n175 585
R1894 B.n380 B.n379 585
R1895 B.n378 B.n243 585
R1896 B.n377 B.n376 585
R1897 B.n375 B.n244 585
R1898 B.n374 B.n373 585
R1899 B.n372 B.n245 585
R1900 B.n371 B.n370 585
R1901 B.n369 B.n246 585
R1902 B.n368 B.n367 585
R1903 B.n366 B.n247 585
R1904 B.n365 B.n364 585
R1905 B.n363 B.n248 585
R1906 B.n362 B.n361 585
R1907 B.n360 B.n249 585
R1908 B.n359 B.n358 585
R1909 B.n357 B.n250 585
R1910 B.n356 B.n355 585
R1911 B.n354 B.n251 585
R1912 B.n353 B.n352 585
R1913 B.n351 B.n252 585
R1914 B.n350 B.n349 585
R1915 B.n348 B.n253 585
R1916 B.n347 B.n346 585
R1917 B.n345 B.n254 585
R1918 B.n344 B.n343 585
R1919 B.n342 B.n255 585
R1920 B.n341 B.n340 585
R1921 B.n339 B.n256 585
R1922 B.n338 B.n337 585
R1923 B.n336 B.n257 585
R1924 B.n335 B.n334 585
R1925 B.n333 B.n258 585
R1926 B.n332 B.n331 585
R1927 B.n330 B.n259 585
R1928 B.n329 B.n328 585
R1929 B.n327 B.n260 585
R1930 B.n326 B.n325 585
R1931 B.n324 B.n261 585
R1932 B.n323 B.n322 585
R1933 B.n321 B.n262 585
R1934 B.n320 B.n319 585
R1935 B.n318 B.n263 585
R1936 B.n317 B.n316 585
R1937 B.n315 B.n264 585
R1938 B.n314 B.n313 585
R1939 B.n312 B.n265 585
R1940 B.n311 B.n310 585
R1941 B.n309 B.n266 585
R1942 B.n308 B.n307 585
R1943 B.n306 B.n267 585
R1944 B.n305 B.n304 585
R1945 B.n303 B.n268 585
R1946 B.n302 B.n301 585
R1947 B.n300 B.n269 585
R1948 B.n299 B.n298 585
R1949 B.n297 B.n270 585
R1950 B.n296 B.n295 585
R1951 B.n294 B.n271 585
R1952 B.n293 B.n292 585
R1953 B.n291 B.n272 585
R1954 B.n290 B.n289 585
R1955 B.n288 B.n273 585
R1956 B.n287 B.n286 585
R1957 B.n285 B.n274 585
R1958 B.n284 B.n283 585
R1959 B.n282 B.n275 585
R1960 B.n281 B.n280 585
R1961 B.n279 B.n276 585
R1962 B.n278 B.n277 585
R1963 B.n2 B.n0 585
R1964 B.n1077 B.n1 585
R1965 B.n1076 B.n1075 585
R1966 B.n1074 B.n3 585
R1967 B.n1073 B.n1072 585
R1968 B.n1071 B.n4 585
R1969 B.n1070 B.n1069 585
R1970 B.n1068 B.n5 585
R1971 B.n1067 B.n1066 585
R1972 B.n1065 B.n6 585
R1973 B.n1064 B.n1063 585
R1974 B.n1062 B.n7 585
R1975 B.n1061 B.n1060 585
R1976 B.n1059 B.n8 585
R1977 B.n1058 B.n1057 585
R1978 B.n1056 B.n9 585
R1979 B.n1055 B.n1054 585
R1980 B.n1053 B.n10 585
R1981 B.n1052 B.n1051 585
R1982 B.n1050 B.n11 585
R1983 B.n1049 B.n1048 585
R1984 B.n1047 B.n12 585
R1985 B.n1046 B.n1045 585
R1986 B.n1044 B.n13 585
R1987 B.n1043 B.n1042 585
R1988 B.n1041 B.n14 585
R1989 B.n1040 B.n1039 585
R1990 B.n1038 B.n15 585
R1991 B.n1037 B.n1036 585
R1992 B.n1035 B.n16 585
R1993 B.n1034 B.n1033 585
R1994 B.n1032 B.n17 585
R1995 B.n1031 B.n1030 585
R1996 B.n1029 B.n18 585
R1997 B.n1028 B.n1027 585
R1998 B.n1026 B.n19 585
R1999 B.n1025 B.n1024 585
R2000 B.n1023 B.n20 585
R2001 B.n1022 B.n1021 585
R2002 B.n1020 B.n21 585
R2003 B.n1019 B.n1018 585
R2004 B.n1017 B.n22 585
R2005 B.n1016 B.n1015 585
R2006 B.n1014 B.n23 585
R2007 B.n1013 B.n1012 585
R2008 B.n1011 B.n24 585
R2009 B.n1010 B.n1009 585
R2010 B.n1008 B.n25 585
R2011 B.n1007 B.n1006 585
R2012 B.n1005 B.n26 585
R2013 B.n1004 B.n1003 585
R2014 B.n1002 B.n27 585
R2015 B.n1001 B.n1000 585
R2016 B.n999 B.n28 585
R2017 B.n998 B.n997 585
R2018 B.n996 B.n29 585
R2019 B.n995 B.n994 585
R2020 B.n993 B.n30 585
R2021 B.n992 B.n991 585
R2022 B.n990 B.n31 585
R2023 B.n989 B.n988 585
R2024 B.n987 B.n32 585
R2025 B.n986 B.n985 585
R2026 B.n984 B.n33 585
R2027 B.n983 B.n982 585
R2028 B.n981 B.n34 585
R2029 B.n980 B.n979 585
R2030 B.n978 B.n35 585
R2031 B.n977 B.n976 585
R2032 B.n975 B.n36 585
R2033 B.n974 B.n973 585
R2034 B.n1079 B.n1078 585
R2035 B.n204 B.t2 558.653
R2036 B.n74 B.t7 558.653
R2037 B.n212 B.t11 558.653
R2038 B.n66 B.t4 558.653
R2039 B.n381 B.n380 511.721
R2040 B.n974 B.n37 511.721
R2041 B.n572 B.n175 511.721
R2042 B.n783 B.n782 511.721
R2043 B.n205 B.t1 476.81
R2044 B.n75 B.t8 476.81
R2045 B.n213 B.t10 476.81
R2046 B.n67 B.t5 476.81
R2047 B.n204 B.t0 318.512
R2048 B.n212 B.t9 318.512
R2049 B.n66 B.t3 318.512
R2050 B.n74 B.t6 318.512
R2051 B.n380 B.n243 163.367
R2052 B.n376 B.n243 163.367
R2053 B.n376 B.n375 163.367
R2054 B.n375 B.n374 163.367
R2055 B.n374 B.n245 163.367
R2056 B.n370 B.n245 163.367
R2057 B.n370 B.n369 163.367
R2058 B.n369 B.n368 163.367
R2059 B.n368 B.n247 163.367
R2060 B.n364 B.n247 163.367
R2061 B.n364 B.n363 163.367
R2062 B.n363 B.n362 163.367
R2063 B.n362 B.n249 163.367
R2064 B.n358 B.n249 163.367
R2065 B.n358 B.n357 163.367
R2066 B.n357 B.n356 163.367
R2067 B.n356 B.n251 163.367
R2068 B.n352 B.n251 163.367
R2069 B.n352 B.n351 163.367
R2070 B.n351 B.n350 163.367
R2071 B.n350 B.n253 163.367
R2072 B.n346 B.n253 163.367
R2073 B.n346 B.n345 163.367
R2074 B.n345 B.n344 163.367
R2075 B.n344 B.n255 163.367
R2076 B.n340 B.n255 163.367
R2077 B.n340 B.n339 163.367
R2078 B.n339 B.n338 163.367
R2079 B.n338 B.n257 163.367
R2080 B.n334 B.n257 163.367
R2081 B.n334 B.n333 163.367
R2082 B.n333 B.n332 163.367
R2083 B.n332 B.n259 163.367
R2084 B.n328 B.n259 163.367
R2085 B.n328 B.n327 163.367
R2086 B.n327 B.n326 163.367
R2087 B.n326 B.n261 163.367
R2088 B.n322 B.n261 163.367
R2089 B.n322 B.n321 163.367
R2090 B.n321 B.n320 163.367
R2091 B.n320 B.n263 163.367
R2092 B.n316 B.n263 163.367
R2093 B.n316 B.n315 163.367
R2094 B.n315 B.n314 163.367
R2095 B.n314 B.n265 163.367
R2096 B.n310 B.n265 163.367
R2097 B.n310 B.n309 163.367
R2098 B.n309 B.n308 163.367
R2099 B.n308 B.n267 163.367
R2100 B.n304 B.n267 163.367
R2101 B.n304 B.n303 163.367
R2102 B.n303 B.n302 163.367
R2103 B.n302 B.n269 163.367
R2104 B.n298 B.n269 163.367
R2105 B.n298 B.n297 163.367
R2106 B.n297 B.n296 163.367
R2107 B.n296 B.n271 163.367
R2108 B.n292 B.n271 163.367
R2109 B.n292 B.n291 163.367
R2110 B.n291 B.n290 163.367
R2111 B.n290 B.n273 163.367
R2112 B.n286 B.n273 163.367
R2113 B.n286 B.n285 163.367
R2114 B.n285 B.n284 163.367
R2115 B.n284 B.n275 163.367
R2116 B.n280 B.n275 163.367
R2117 B.n280 B.n279 163.367
R2118 B.n279 B.n278 163.367
R2119 B.n278 B.n2 163.367
R2120 B.n1078 B.n2 163.367
R2121 B.n1078 B.n1077 163.367
R2122 B.n1077 B.n1076 163.367
R2123 B.n1076 B.n3 163.367
R2124 B.n1072 B.n3 163.367
R2125 B.n1072 B.n1071 163.367
R2126 B.n1071 B.n1070 163.367
R2127 B.n1070 B.n5 163.367
R2128 B.n1066 B.n5 163.367
R2129 B.n1066 B.n1065 163.367
R2130 B.n1065 B.n1064 163.367
R2131 B.n1064 B.n7 163.367
R2132 B.n1060 B.n7 163.367
R2133 B.n1060 B.n1059 163.367
R2134 B.n1059 B.n1058 163.367
R2135 B.n1058 B.n9 163.367
R2136 B.n1054 B.n9 163.367
R2137 B.n1054 B.n1053 163.367
R2138 B.n1053 B.n1052 163.367
R2139 B.n1052 B.n11 163.367
R2140 B.n1048 B.n11 163.367
R2141 B.n1048 B.n1047 163.367
R2142 B.n1047 B.n1046 163.367
R2143 B.n1046 B.n13 163.367
R2144 B.n1042 B.n13 163.367
R2145 B.n1042 B.n1041 163.367
R2146 B.n1041 B.n1040 163.367
R2147 B.n1040 B.n15 163.367
R2148 B.n1036 B.n15 163.367
R2149 B.n1036 B.n1035 163.367
R2150 B.n1035 B.n1034 163.367
R2151 B.n1034 B.n17 163.367
R2152 B.n1030 B.n17 163.367
R2153 B.n1030 B.n1029 163.367
R2154 B.n1029 B.n1028 163.367
R2155 B.n1028 B.n19 163.367
R2156 B.n1024 B.n19 163.367
R2157 B.n1024 B.n1023 163.367
R2158 B.n1023 B.n1022 163.367
R2159 B.n1022 B.n21 163.367
R2160 B.n1018 B.n21 163.367
R2161 B.n1018 B.n1017 163.367
R2162 B.n1017 B.n1016 163.367
R2163 B.n1016 B.n23 163.367
R2164 B.n1012 B.n23 163.367
R2165 B.n1012 B.n1011 163.367
R2166 B.n1011 B.n1010 163.367
R2167 B.n1010 B.n25 163.367
R2168 B.n1006 B.n25 163.367
R2169 B.n1006 B.n1005 163.367
R2170 B.n1005 B.n1004 163.367
R2171 B.n1004 B.n27 163.367
R2172 B.n1000 B.n27 163.367
R2173 B.n1000 B.n999 163.367
R2174 B.n999 B.n998 163.367
R2175 B.n998 B.n29 163.367
R2176 B.n994 B.n29 163.367
R2177 B.n994 B.n993 163.367
R2178 B.n993 B.n992 163.367
R2179 B.n992 B.n31 163.367
R2180 B.n988 B.n31 163.367
R2181 B.n988 B.n987 163.367
R2182 B.n987 B.n986 163.367
R2183 B.n986 B.n33 163.367
R2184 B.n982 B.n33 163.367
R2185 B.n982 B.n981 163.367
R2186 B.n981 B.n980 163.367
R2187 B.n980 B.n35 163.367
R2188 B.n976 B.n35 163.367
R2189 B.n976 B.n975 163.367
R2190 B.n975 B.n974 163.367
R2191 B.n382 B.n381 163.367
R2192 B.n382 B.n241 163.367
R2193 B.n386 B.n241 163.367
R2194 B.n387 B.n386 163.367
R2195 B.n388 B.n387 163.367
R2196 B.n388 B.n239 163.367
R2197 B.n392 B.n239 163.367
R2198 B.n393 B.n392 163.367
R2199 B.n394 B.n393 163.367
R2200 B.n394 B.n237 163.367
R2201 B.n398 B.n237 163.367
R2202 B.n399 B.n398 163.367
R2203 B.n400 B.n399 163.367
R2204 B.n400 B.n235 163.367
R2205 B.n404 B.n235 163.367
R2206 B.n405 B.n404 163.367
R2207 B.n406 B.n405 163.367
R2208 B.n406 B.n233 163.367
R2209 B.n410 B.n233 163.367
R2210 B.n411 B.n410 163.367
R2211 B.n412 B.n411 163.367
R2212 B.n412 B.n231 163.367
R2213 B.n416 B.n231 163.367
R2214 B.n417 B.n416 163.367
R2215 B.n418 B.n417 163.367
R2216 B.n418 B.n229 163.367
R2217 B.n422 B.n229 163.367
R2218 B.n423 B.n422 163.367
R2219 B.n424 B.n423 163.367
R2220 B.n424 B.n227 163.367
R2221 B.n428 B.n227 163.367
R2222 B.n429 B.n428 163.367
R2223 B.n430 B.n429 163.367
R2224 B.n430 B.n225 163.367
R2225 B.n434 B.n225 163.367
R2226 B.n435 B.n434 163.367
R2227 B.n436 B.n435 163.367
R2228 B.n436 B.n223 163.367
R2229 B.n440 B.n223 163.367
R2230 B.n441 B.n440 163.367
R2231 B.n442 B.n441 163.367
R2232 B.n442 B.n221 163.367
R2233 B.n446 B.n221 163.367
R2234 B.n447 B.n446 163.367
R2235 B.n448 B.n447 163.367
R2236 B.n448 B.n219 163.367
R2237 B.n452 B.n219 163.367
R2238 B.n453 B.n452 163.367
R2239 B.n454 B.n453 163.367
R2240 B.n454 B.n217 163.367
R2241 B.n458 B.n217 163.367
R2242 B.n459 B.n458 163.367
R2243 B.n460 B.n459 163.367
R2244 B.n460 B.n215 163.367
R2245 B.n464 B.n215 163.367
R2246 B.n465 B.n464 163.367
R2247 B.n466 B.n465 163.367
R2248 B.n466 B.n211 163.367
R2249 B.n471 B.n211 163.367
R2250 B.n472 B.n471 163.367
R2251 B.n473 B.n472 163.367
R2252 B.n473 B.n209 163.367
R2253 B.n477 B.n209 163.367
R2254 B.n478 B.n477 163.367
R2255 B.n479 B.n478 163.367
R2256 B.n479 B.n207 163.367
R2257 B.n483 B.n207 163.367
R2258 B.n484 B.n483 163.367
R2259 B.n484 B.n203 163.367
R2260 B.n488 B.n203 163.367
R2261 B.n489 B.n488 163.367
R2262 B.n490 B.n489 163.367
R2263 B.n490 B.n201 163.367
R2264 B.n494 B.n201 163.367
R2265 B.n495 B.n494 163.367
R2266 B.n496 B.n495 163.367
R2267 B.n496 B.n199 163.367
R2268 B.n500 B.n199 163.367
R2269 B.n501 B.n500 163.367
R2270 B.n502 B.n501 163.367
R2271 B.n502 B.n197 163.367
R2272 B.n506 B.n197 163.367
R2273 B.n507 B.n506 163.367
R2274 B.n508 B.n507 163.367
R2275 B.n508 B.n195 163.367
R2276 B.n512 B.n195 163.367
R2277 B.n513 B.n512 163.367
R2278 B.n514 B.n513 163.367
R2279 B.n514 B.n193 163.367
R2280 B.n518 B.n193 163.367
R2281 B.n519 B.n518 163.367
R2282 B.n520 B.n519 163.367
R2283 B.n520 B.n191 163.367
R2284 B.n524 B.n191 163.367
R2285 B.n525 B.n524 163.367
R2286 B.n526 B.n525 163.367
R2287 B.n526 B.n189 163.367
R2288 B.n530 B.n189 163.367
R2289 B.n531 B.n530 163.367
R2290 B.n532 B.n531 163.367
R2291 B.n532 B.n187 163.367
R2292 B.n536 B.n187 163.367
R2293 B.n537 B.n536 163.367
R2294 B.n538 B.n537 163.367
R2295 B.n538 B.n185 163.367
R2296 B.n542 B.n185 163.367
R2297 B.n543 B.n542 163.367
R2298 B.n544 B.n543 163.367
R2299 B.n544 B.n183 163.367
R2300 B.n548 B.n183 163.367
R2301 B.n549 B.n548 163.367
R2302 B.n550 B.n549 163.367
R2303 B.n550 B.n181 163.367
R2304 B.n554 B.n181 163.367
R2305 B.n555 B.n554 163.367
R2306 B.n556 B.n555 163.367
R2307 B.n556 B.n179 163.367
R2308 B.n560 B.n179 163.367
R2309 B.n561 B.n560 163.367
R2310 B.n562 B.n561 163.367
R2311 B.n562 B.n177 163.367
R2312 B.n566 B.n177 163.367
R2313 B.n567 B.n566 163.367
R2314 B.n568 B.n567 163.367
R2315 B.n568 B.n175 163.367
R2316 B.n573 B.n572 163.367
R2317 B.n574 B.n573 163.367
R2318 B.n574 B.n173 163.367
R2319 B.n578 B.n173 163.367
R2320 B.n579 B.n578 163.367
R2321 B.n580 B.n579 163.367
R2322 B.n580 B.n171 163.367
R2323 B.n584 B.n171 163.367
R2324 B.n585 B.n584 163.367
R2325 B.n586 B.n585 163.367
R2326 B.n586 B.n169 163.367
R2327 B.n590 B.n169 163.367
R2328 B.n591 B.n590 163.367
R2329 B.n592 B.n591 163.367
R2330 B.n592 B.n167 163.367
R2331 B.n596 B.n167 163.367
R2332 B.n597 B.n596 163.367
R2333 B.n598 B.n597 163.367
R2334 B.n598 B.n165 163.367
R2335 B.n602 B.n165 163.367
R2336 B.n603 B.n602 163.367
R2337 B.n604 B.n603 163.367
R2338 B.n604 B.n163 163.367
R2339 B.n608 B.n163 163.367
R2340 B.n609 B.n608 163.367
R2341 B.n610 B.n609 163.367
R2342 B.n610 B.n161 163.367
R2343 B.n614 B.n161 163.367
R2344 B.n615 B.n614 163.367
R2345 B.n616 B.n615 163.367
R2346 B.n616 B.n159 163.367
R2347 B.n620 B.n159 163.367
R2348 B.n621 B.n620 163.367
R2349 B.n622 B.n621 163.367
R2350 B.n622 B.n157 163.367
R2351 B.n626 B.n157 163.367
R2352 B.n627 B.n626 163.367
R2353 B.n628 B.n627 163.367
R2354 B.n628 B.n155 163.367
R2355 B.n632 B.n155 163.367
R2356 B.n633 B.n632 163.367
R2357 B.n634 B.n633 163.367
R2358 B.n634 B.n153 163.367
R2359 B.n638 B.n153 163.367
R2360 B.n639 B.n638 163.367
R2361 B.n640 B.n639 163.367
R2362 B.n640 B.n151 163.367
R2363 B.n644 B.n151 163.367
R2364 B.n645 B.n644 163.367
R2365 B.n646 B.n645 163.367
R2366 B.n646 B.n149 163.367
R2367 B.n650 B.n149 163.367
R2368 B.n651 B.n650 163.367
R2369 B.n652 B.n651 163.367
R2370 B.n652 B.n147 163.367
R2371 B.n656 B.n147 163.367
R2372 B.n657 B.n656 163.367
R2373 B.n658 B.n657 163.367
R2374 B.n658 B.n145 163.367
R2375 B.n662 B.n145 163.367
R2376 B.n663 B.n662 163.367
R2377 B.n664 B.n663 163.367
R2378 B.n664 B.n143 163.367
R2379 B.n668 B.n143 163.367
R2380 B.n669 B.n668 163.367
R2381 B.n670 B.n669 163.367
R2382 B.n670 B.n141 163.367
R2383 B.n674 B.n141 163.367
R2384 B.n675 B.n674 163.367
R2385 B.n676 B.n675 163.367
R2386 B.n676 B.n139 163.367
R2387 B.n680 B.n139 163.367
R2388 B.n681 B.n680 163.367
R2389 B.n682 B.n681 163.367
R2390 B.n682 B.n137 163.367
R2391 B.n686 B.n137 163.367
R2392 B.n687 B.n686 163.367
R2393 B.n688 B.n687 163.367
R2394 B.n688 B.n135 163.367
R2395 B.n692 B.n135 163.367
R2396 B.n693 B.n692 163.367
R2397 B.n694 B.n693 163.367
R2398 B.n694 B.n133 163.367
R2399 B.n698 B.n133 163.367
R2400 B.n699 B.n698 163.367
R2401 B.n700 B.n699 163.367
R2402 B.n700 B.n131 163.367
R2403 B.n704 B.n131 163.367
R2404 B.n705 B.n704 163.367
R2405 B.n706 B.n705 163.367
R2406 B.n706 B.n129 163.367
R2407 B.n710 B.n129 163.367
R2408 B.n711 B.n710 163.367
R2409 B.n712 B.n711 163.367
R2410 B.n712 B.n127 163.367
R2411 B.n716 B.n127 163.367
R2412 B.n717 B.n716 163.367
R2413 B.n718 B.n717 163.367
R2414 B.n718 B.n125 163.367
R2415 B.n722 B.n125 163.367
R2416 B.n723 B.n722 163.367
R2417 B.n724 B.n723 163.367
R2418 B.n724 B.n123 163.367
R2419 B.n728 B.n123 163.367
R2420 B.n729 B.n728 163.367
R2421 B.n730 B.n729 163.367
R2422 B.n730 B.n121 163.367
R2423 B.n734 B.n121 163.367
R2424 B.n735 B.n734 163.367
R2425 B.n736 B.n735 163.367
R2426 B.n736 B.n119 163.367
R2427 B.n740 B.n119 163.367
R2428 B.n741 B.n740 163.367
R2429 B.n742 B.n741 163.367
R2430 B.n742 B.n117 163.367
R2431 B.n746 B.n117 163.367
R2432 B.n747 B.n746 163.367
R2433 B.n748 B.n747 163.367
R2434 B.n748 B.n115 163.367
R2435 B.n752 B.n115 163.367
R2436 B.n753 B.n752 163.367
R2437 B.n754 B.n753 163.367
R2438 B.n754 B.n113 163.367
R2439 B.n758 B.n113 163.367
R2440 B.n759 B.n758 163.367
R2441 B.n760 B.n759 163.367
R2442 B.n760 B.n111 163.367
R2443 B.n764 B.n111 163.367
R2444 B.n765 B.n764 163.367
R2445 B.n766 B.n765 163.367
R2446 B.n766 B.n109 163.367
R2447 B.n770 B.n109 163.367
R2448 B.n771 B.n770 163.367
R2449 B.n772 B.n771 163.367
R2450 B.n772 B.n107 163.367
R2451 B.n776 B.n107 163.367
R2452 B.n777 B.n776 163.367
R2453 B.n778 B.n777 163.367
R2454 B.n778 B.n105 163.367
R2455 B.n782 B.n105 163.367
R2456 B.n970 B.n37 163.367
R2457 B.n970 B.n969 163.367
R2458 B.n969 B.n968 163.367
R2459 B.n968 B.n39 163.367
R2460 B.n964 B.n39 163.367
R2461 B.n964 B.n963 163.367
R2462 B.n963 B.n962 163.367
R2463 B.n962 B.n41 163.367
R2464 B.n958 B.n41 163.367
R2465 B.n958 B.n957 163.367
R2466 B.n957 B.n956 163.367
R2467 B.n956 B.n43 163.367
R2468 B.n952 B.n43 163.367
R2469 B.n952 B.n951 163.367
R2470 B.n951 B.n950 163.367
R2471 B.n950 B.n45 163.367
R2472 B.n946 B.n45 163.367
R2473 B.n946 B.n945 163.367
R2474 B.n945 B.n944 163.367
R2475 B.n944 B.n47 163.367
R2476 B.n940 B.n47 163.367
R2477 B.n940 B.n939 163.367
R2478 B.n939 B.n938 163.367
R2479 B.n938 B.n49 163.367
R2480 B.n934 B.n49 163.367
R2481 B.n934 B.n933 163.367
R2482 B.n933 B.n932 163.367
R2483 B.n932 B.n51 163.367
R2484 B.n928 B.n51 163.367
R2485 B.n928 B.n927 163.367
R2486 B.n927 B.n926 163.367
R2487 B.n926 B.n53 163.367
R2488 B.n922 B.n53 163.367
R2489 B.n922 B.n921 163.367
R2490 B.n921 B.n920 163.367
R2491 B.n920 B.n55 163.367
R2492 B.n916 B.n55 163.367
R2493 B.n916 B.n915 163.367
R2494 B.n915 B.n914 163.367
R2495 B.n914 B.n57 163.367
R2496 B.n910 B.n57 163.367
R2497 B.n910 B.n909 163.367
R2498 B.n909 B.n908 163.367
R2499 B.n908 B.n59 163.367
R2500 B.n904 B.n59 163.367
R2501 B.n904 B.n903 163.367
R2502 B.n903 B.n902 163.367
R2503 B.n902 B.n61 163.367
R2504 B.n898 B.n61 163.367
R2505 B.n898 B.n897 163.367
R2506 B.n897 B.n896 163.367
R2507 B.n896 B.n63 163.367
R2508 B.n892 B.n63 163.367
R2509 B.n892 B.n891 163.367
R2510 B.n891 B.n890 163.367
R2511 B.n890 B.n65 163.367
R2512 B.n886 B.n65 163.367
R2513 B.n886 B.n885 163.367
R2514 B.n885 B.n69 163.367
R2515 B.n881 B.n69 163.367
R2516 B.n881 B.n880 163.367
R2517 B.n880 B.n879 163.367
R2518 B.n879 B.n71 163.367
R2519 B.n875 B.n71 163.367
R2520 B.n875 B.n874 163.367
R2521 B.n874 B.n873 163.367
R2522 B.n873 B.n73 163.367
R2523 B.n868 B.n73 163.367
R2524 B.n868 B.n867 163.367
R2525 B.n867 B.n866 163.367
R2526 B.n866 B.n77 163.367
R2527 B.n862 B.n77 163.367
R2528 B.n862 B.n861 163.367
R2529 B.n861 B.n860 163.367
R2530 B.n860 B.n79 163.367
R2531 B.n856 B.n79 163.367
R2532 B.n856 B.n855 163.367
R2533 B.n855 B.n854 163.367
R2534 B.n854 B.n81 163.367
R2535 B.n850 B.n81 163.367
R2536 B.n850 B.n849 163.367
R2537 B.n849 B.n848 163.367
R2538 B.n848 B.n83 163.367
R2539 B.n844 B.n83 163.367
R2540 B.n844 B.n843 163.367
R2541 B.n843 B.n842 163.367
R2542 B.n842 B.n85 163.367
R2543 B.n838 B.n85 163.367
R2544 B.n838 B.n837 163.367
R2545 B.n837 B.n836 163.367
R2546 B.n836 B.n87 163.367
R2547 B.n832 B.n87 163.367
R2548 B.n832 B.n831 163.367
R2549 B.n831 B.n830 163.367
R2550 B.n830 B.n89 163.367
R2551 B.n826 B.n89 163.367
R2552 B.n826 B.n825 163.367
R2553 B.n825 B.n824 163.367
R2554 B.n824 B.n91 163.367
R2555 B.n820 B.n91 163.367
R2556 B.n820 B.n819 163.367
R2557 B.n819 B.n818 163.367
R2558 B.n818 B.n93 163.367
R2559 B.n814 B.n93 163.367
R2560 B.n814 B.n813 163.367
R2561 B.n813 B.n812 163.367
R2562 B.n812 B.n95 163.367
R2563 B.n808 B.n95 163.367
R2564 B.n808 B.n807 163.367
R2565 B.n807 B.n806 163.367
R2566 B.n806 B.n97 163.367
R2567 B.n802 B.n97 163.367
R2568 B.n802 B.n801 163.367
R2569 B.n801 B.n800 163.367
R2570 B.n800 B.n99 163.367
R2571 B.n796 B.n99 163.367
R2572 B.n796 B.n795 163.367
R2573 B.n795 B.n794 163.367
R2574 B.n794 B.n101 163.367
R2575 B.n790 B.n101 163.367
R2576 B.n790 B.n789 163.367
R2577 B.n789 B.n788 163.367
R2578 B.n788 B.n103 163.367
R2579 B.n784 B.n103 163.367
R2580 B.n784 B.n783 163.367
R2581 B.n205 B.n204 81.8429
R2582 B.n213 B.n212 81.8429
R2583 B.n67 B.n66 81.8429
R2584 B.n75 B.n74 81.8429
R2585 B.n206 B.n205 59.5399
R2586 B.n468 B.n213 59.5399
R2587 B.n68 B.n67 59.5399
R2588 B.n870 B.n75 59.5399
R2589 B.n973 B.n972 33.2493
R2590 B.n781 B.n104 33.2493
R2591 B.n571 B.n570 33.2493
R2592 B.n379 B.n242 33.2493
R2593 B B.n1079 18.0485
R2594 B.n972 B.n971 10.6151
R2595 B.n971 B.n38 10.6151
R2596 B.n967 B.n38 10.6151
R2597 B.n967 B.n966 10.6151
R2598 B.n966 B.n965 10.6151
R2599 B.n965 B.n40 10.6151
R2600 B.n961 B.n40 10.6151
R2601 B.n961 B.n960 10.6151
R2602 B.n960 B.n959 10.6151
R2603 B.n959 B.n42 10.6151
R2604 B.n955 B.n42 10.6151
R2605 B.n955 B.n954 10.6151
R2606 B.n954 B.n953 10.6151
R2607 B.n953 B.n44 10.6151
R2608 B.n949 B.n44 10.6151
R2609 B.n949 B.n948 10.6151
R2610 B.n948 B.n947 10.6151
R2611 B.n947 B.n46 10.6151
R2612 B.n943 B.n46 10.6151
R2613 B.n943 B.n942 10.6151
R2614 B.n942 B.n941 10.6151
R2615 B.n941 B.n48 10.6151
R2616 B.n937 B.n48 10.6151
R2617 B.n937 B.n936 10.6151
R2618 B.n936 B.n935 10.6151
R2619 B.n935 B.n50 10.6151
R2620 B.n931 B.n50 10.6151
R2621 B.n931 B.n930 10.6151
R2622 B.n930 B.n929 10.6151
R2623 B.n929 B.n52 10.6151
R2624 B.n925 B.n52 10.6151
R2625 B.n925 B.n924 10.6151
R2626 B.n924 B.n923 10.6151
R2627 B.n923 B.n54 10.6151
R2628 B.n919 B.n54 10.6151
R2629 B.n919 B.n918 10.6151
R2630 B.n918 B.n917 10.6151
R2631 B.n917 B.n56 10.6151
R2632 B.n913 B.n56 10.6151
R2633 B.n913 B.n912 10.6151
R2634 B.n912 B.n911 10.6151
R2635 B.n911 B.n58 10.6151
R2636 B.n907 B.n58 10.6151
R2637 B.n907 B.n906 10.6151
R2638 B.n906 B.n905 10.6151
R2639 B.n905 B.n60 10.6151
R2640 B.n901 B.n60 10.6151
R2641 B.n901 B.n900 10.6151
R2642 B.n900 B.n899 10.6151
R2643 B.n899 B.n62 10.6151
R2644 B.n895 B.n62 10.6151
R2645 B.n895 B.n894 10.6151
R2646 B.n894 B.n893 10.6151
R2647 B.n893 B.n64 10.6151
R2648 B.n889 B.n64 10.6151
R2649 B.n889 B.n888 10.6151
R2650 B.n888 B.n887 10.6151
R2651 B.n884 B.n883 10.6151
R2652 B.n883 B.n882 10.6151
R2653 B.n882 B.n70 10.6151
R2654 B.n878 B.n70 10.6151
R2655 B.n878 B.n877 10.6151
R2656 B.n877 B.n876 10.6151
R2657 B.n876 B.n72 10.6151
R2658 B.n872 B.n72 10.6151
R2659 B.n872 B.n871 10.6151
R2660 B.n869 B.n76 10.6151
R2661 B.n865 B.n76 10.6151
R2662 B.n865 B.n864 10.6151
R2663 B.n864 B.n863 10.6151
R2664 B.n863 B.n78 10.6151
R2665 B.n859 B.n78 10.6151
R2666 B.n859 B.n858 10.6151
R2667 B.n858 B.n857 10.6151
R2668 B.n857 B.n80 10.6151
R2669 B.n853 B.n80 10.6151
R2670 B.n853 B.n852 10.6151
R2671 B.n852 B.n851 10.6151
R2672 B.n851 B.n82 10.6151
R2673 B.n847 B.n82 10.6151
R2674 B.n847 B.n846 10.6151
R2675 B.n846 B.n845 10.6151
R2676 B.n845 B.n84 10.6151
R2677 B.n841 B.n84 10.6151
R2678 B.n841 B.n840 10.6151
R2679 B.n840 B.n839 10.6151
R2680 B.n839 B.n86 10.6151
R2681 B.n835 B.n86 10.6151
R2682 B.n835 B.n834 10.6151
R2683 B.n834 B.n833 10.6151
R2684 B.n833 B.n88 10.6151
R2685 B.n829 B.n88 10.6151
R2686 B.n829 B.n828 10.6151
R2687 B.n828 B.n827 10.6151
R2688 B.n827 B.n90 10.6151
R2689 B.n823 B.n90 10.6151
R2690 B.n823 B.n822 10.6151
R2691 B.n822 B.n821 10.6151
R2692 B.n821 B.n92 10.6151
R2693 B.n817 B.n92 10.6151
R2694 B.n817 B.n816 10.6151
R2695 B.n816 B.n815 10.6151
R2696 B.n815 B.n94 10.6151
R2697 B.n811 B.n94 10.6151
R2698 B.n811 B.n810 10.6151
R2699 B.n810 B.n809 10.6151
R2700 B.n809 B.n96 10.6151
R2701 B.n805 B.n96 10.6151
R2702 B.n805 B.n804 10.6151
R2703 B.n804 B.n803 10.6151
R2704 B.n803 B.n98 10.6151
R2705 B.n799 B.n98 10.6151
R2706 B.n799 B.n798 10.6151
R2707 B.n798 B.n797 10.6151
R2708 B.n797 B.n100 10.6151
R2709 B.n793 B.n100 10.6151
R2710 B.n793 B.n792 10.6151
R2711 B.n792 B.n791 10.6151
R2712 B.n791 B.n102 10.6151
R2713 B.n787 B.n102 10.6151
R2714 B.n787 B.n786 10.6151
R2715 B.n786 B.n785 10.6151
R2716 B.n785 B.n104 10.6151
R2717 B.n571 B.n174 10.6151
R2718 B.n575 B.n174 10.6151
R2719 B.n576 B.n575 10.6151
R2720 B.n577 B.n576 10.6151
R2721 B.n577 B.n172 10.6151
R2722 B.n581 B.n172 10.6151
R2723 B.n582 B.n581 10.6151
R2724 B.n583 B.n582 10.6151
R2725 B.n583 B.n170 10.6151
R2726 B.n587 B.n170 10.6151
R2727 B.n588 B.n587 10.6151
R2728 B.n589 B.n588 10.6151
R2729 B.n589 B.n168 10.6151
R2730 B.n593 B.n168 10.6151
R2731 B.n594 B.n593 10.6151
R2732 B.n595 B.n594 10.6151
R2733 B.n595 B.n166 10.6151
R2734 B.n599 B.n166 10.6151
R2735 B.n600 B.n599 10.6151
R2736 B.n601 B.n600 10.6151
R2737 B.n601 B.n164 10.6151
R2738 B.n605 B.n164 10.6151
R2739 B.n606 B.n605 10.6151
R2740 B.n607 B.n606 10.6151
R2741 B.n607 B.n162 10.6151
R2742 B.n611 B.n162 10.6151
R2743 B.n612 B.n611 10.6151
R2744 B.n613 B.n612 10.6151
R2745 B.n613 B.n160 10.6151
R2746 B.n617 B.n160 10.6151
R2747 B.n618 B.n617 10.6151
R2748 B.n619 B.n618 10.6151
R2749 B.n619 B.n158 10.6151
R2750 B.n623 B.n158 10.6151
R2751 B.n624 B.n623 10.6151
R2752 B.n625 B.n624 10.6151
R2753 B.n625 B.n156 10.6151
R2754 B.n629 B.n156 10.6151
R2755 B.n630 B.n629 10.6151
R2756 B.n631 B.n630 10.6151
R2757 B.n631 B.n154 10.6151
R2758 B.n635 B.n154 10.6151
R2759 B.n636 B.n635 10.6151
R2760 B.n637 B.n636 10.6151
R2761 B.n637 B.n152 10.6151
R2762 B.n641 B.n152 10.6151
R2763 B.n642 B.n641 10.6151
R2764 B.n643 B.n642 10.6151
R2765 B.n643 B.n150 10.6151
R2766 B.n647 B.n150 10.6151
R2767 B.n648 B.n647 10.6151
R2768 B.n649 B.n648 10.6151
R2769 B.n649 B.n148 10.6151
R2770 B.n653 B.n148 10.6151
R2771 B.n654 B.n653 10.6151
R2772 B.n655 B.n654 10.6151
R2773 B.n655 B.n146 10.6151
R2774 B.n659 B.n146 10.6151
R2775 B.n660 B.n659 10.6151
R2776 B.n661 B.n660 10.6151
R2777 B.n661 B.n144 10.6151
R2778 B.n665 B.n144 10.6151
R2779 B.n666 B.n665 10.6151
R2780 B.n667 B.n666 10.6151
R2781 B.n667 B.n142 10.6151
R2782 B.n671 B.n142 10.6151
R2783 B.n672 B.n671 10.6151
R2784 B.n673 B.n672 10.6151
R2785 B.n673 B.n140 10.6151
R2786 B.n677 B.n140 10.6151
R2787 B.n678 B.n677 10.6151
R2788 B.n679 B.n678 10.6151
R2789 B.n679 B.n138 10.6151
R2790 B.n683 B.n138 10.6151
R2791 B.n684 B.n683 10.6151
R2792 B.n685 B.n684 10.6151
R2793 B.n685 B.n136 10.6151
R2794 B.n689 B.n136 10.6151
R2795 B.n690 B.n689 10.6151
R2796 B.n691 B.n690 10.6151
R2797 B.n691 B.n134 10.6151
R2798 B.n695 B.n134 10.6151
R2799 B.n696 B.n695 10.6151
R2800 B.n697 B.n696 10.6151
R2801 B.n697 B.n132 10.6151
R2802 B.n701 B.n132 10.6151
R2803 B.n702 B.n701 10.6151
R2804 B.n703 B.n702 10.6151
R2805 B.n703 B.n130 10.6151
R2806 B.n707 B.n130 10.6151
R2807 B.n708 B.n707 10.6151
R2808 B.n709 B.n708 10.6151
R2809 B.n709 B.n128 10.6151
R2810 B.n713 B.n128 10.6151
R2811 B.n714 B.n713 10.6151
R2812 B.n715 B.n714 10.6151
R2813 B.n715 B.n126 10.6151
R2814 B.n719 B.n126 10.6151
R2815 B.n720 B.n719 10.6151
R2816 B.n721 B.n720 10.6151
R2817 B.n721 B.n124 10.6151
R2818 B.n725 B.n124 10.6151
R2819 B.n726 B.n725 10.6151
R2820 B.n727 B.n726 10.6151
R2821 B.n727 B.n122 10.6151
R2822 B.n731 B.n122 10.6151
R2823 B.n732 B.n731 10.6151
R2824 B.n733 B.n732 10.6151
R2825 B.n733 B.n120 10.6151
R2826 B.n737 B.n120 10.6151
R2827 B.n738 B.n737 10.6151
R2828 B.n739 B.n738 10.6151
R2829 B.n739 B.n118 10.6151
R2830 B.n743 B.n118 10.6151
R2831 B.n744 B.n743 10.6151
R2832 B.n745 B.n744 10.6151
R2833 B.n745 B.n116 10.6151
R2834 B.n749 B.n116 10.6151
R2835 B.n750 B.n749 10.6151
R2836 B.n751 B.n750 10.6151
R2837 B.n751 B.n114 10.6151
R2838 B.n755 B.n114 10.6151
R2839 B.n756 B.n755 10.6151
R2840 B.n757 B.n756 10.6151
R2841 B.n757 B.n112 10.6151
R2842 B.n761 B.n112 10.6151
R2843 B.n762 B.n761 10.6151
R2844 B.n763 B.n762 10.6151
R2845 B.n763 B.n110 10.6151
R2846 B.n767 B.n110 10.6151
R2847 B.n768 B.n767 10.6151
R2848 B.n769 B.n768 10.6151
R2849 B.n769 B.n108 10.6151
R2850 B.n773 B.n108 10.6151
R2851 B.n774 B.n773 10.6151
R2852 B.n775 B.n774 10.6151
R2853 B.n775 B.n106 10.6151
R2854 B.n779 B.n106 10.6151
R2855 B.n780 B.n779 10.6151
R2856 B.n781 B.n780 10.6151
R2857 B.n383 B.n242 10.6151
R2858 B.n384 B.n383 10.6151
R2859 B.n385 B.n384 10.6151
R2860 B.n385 B.n240 10.6151
R2861 B.n389 B.n240 10.6151
R2862 B.n390 B.n389 10.6151
R2863 B.n391 B.n390 10.6151
R2864 B.n391 B.n238 10.6151
R2865 B.n395 B.n238 10.6151
R2866 B.n396 B.n395 10.6151
R2867 B.n397 B.n396 10.6151
R2868 B.n397 B.n236 10.6151
R2869 B.n401 B.n236 10.6151
R2870 B.n402 B.n401 10.6151
R2871 B.n403 B.n402 10.6151
R2872 B.n403 B.n234 10.6151
R2873 B.n407 B.n234 10.6151
R2874 B.n408 B.n407 10.6151
R2875 B.n409 B.n408 10.6151
R2876 B.n409 B.n232 10.6151
R2877 B.n413 B.n232 10.6151
R2878 B.n414 B.n413 10.6151
R2879 B.n415 B.n414 10.6151
R2880 B.n415 B.n230 10.6151
R2881 B.n419 B.n230 10.6151
R2882 B.n420 B.n419 10.6151
R2883 B.n421 B.n420 10.6151
R2884 B.n421 B.n228 10.6151
R2885 B.n425 B.n228 10.6151
R2886 B.n426 B.n425 10.6151
R2887 B.n427 B.n426 10.6151
R2888 B.n427 B.n226 10.6151
R2889 B.n431 B.n226 10.6151
R2890 B.n432 B.n431 10.6151
R2891 B.n433 B.n432 10.6151
R2892 B.n433 B.n224 10.6151
R2893 B.n437 B.n224 10.6151
R2894 B.n438 B.n437 10.6151
R2895 B.n439 B.n438 10.6151
R2896 B.n439 B.n222 10.6151
R2897 B.n443 B.n222 10.6151
R2898 B.n444 B.n443 10.6151
R2899 B.n445 B.n444 10.6151
R2900 B.n445 B.n220 10.6151
R2901 B.n449 B.n220 10.6151
R2902 B.n450 B.n449 10.6151
R2903 B.n451 B.n450 10.6151
R2904 B.n451 B.n218 10.6151
R2905 B.n455 B.n218 10.6151
R2906 B.n456 B.n455 10.6151
R2907 B.n457 B.n456 10.6151
R2908 B.n457 B.n216 10.6151
R2909 B.n461 B.n216 10.6151
R2910 B.n462 B.n461 10.6151
R2911 B.n463 B.n462 10.6151
R2912 B.n463 B.n214 10.6151
R2913 B.n467 B.n214 10.6151
R2914 B.n470 B.n469 10.6151
R2915 B.n470 B.n210 10.6151
R2916 B.n474 B.n210 10.6151
R2917 B.n475 B.n474 10.6151
R2918 B.n476 B.n475 10.6151
R2919 B.n476 B.n208 10.6151
R2920 B.n480 B.n208 10.6151
R2921 B.n481 B.n480 10.6151
R2922 B.n482 B.n481 10.6151
R2923 B.n486 B.n485 10.6151
R2924 B.n487 B.n486 10.6151
R2925 B.n487 B.n202 10.6151
R2926 B.n491 B.n202 10.6151
R2927 B.n492 B.n491 10.6151
R2928 B.n493 B.n492 10.6151
R2929 B.n493 B.n200 10.6151
R2930 B.n497 B.n200 10.6151
R2931 B.n498 B.n497 10.6151
R2932 B.n499 B.n498 10.6151
R2933 B.n499 B.n198 10.6151
R2934 B.n503 B.n198 10.6151
R2935 B.n504 B.n503 10.6151
R2936 B.n505 B.n504 10.6151
R2937 B.n505 B.n196 10.6151
R2938 B.n509 B.n196 10.6151
R2939 B.n510 B.n509 10.6151
R2940 B.n511 B.n510 10.6151
R2941 B.n511 B.n194 10.6151
R2942 B.n515 B.n194 10.6151
R2943 B.n516 B.n515 10.6151
R2944 B.n517 B.n516 10.6151
R2945 B.n517 B.n192 10.6151
R2946 B.n521 B.n192 10.6151
R2947 B.n522 B.n521 10.6151
R2948 B.n523 B.n522 10.6151
R2949 B.n523 B.n190 10.6151
R2950 B.n527 B.n190 10.6151
R2951 B.n528 B.n527 10.6151
R2952 B.n529 B.n528 10.6151
R2953 B.n529 B.n188 10.6151
R2954 B.n533 B.n188 10.6151
R2955 B.n534 B.n533 10.6151
R2956 B.n535 B.n534 10.6151
R2957 B.n535 B.n186 10.6151
R2958 B.n539 B.n186 10.6151
R2959 B.n540 B.n539 10.6151
R2960 B.n541 B.n540 10.6151
R2961 B.n541 B.n184 10.6151
R2962 B.n545 B.n184 10.6151
R2963 B.n546 B.n545 10.6151
R2964 B.n547 B.n546 10.6151
R2965 B.n547 B.n182 10.6151
R2966 B.n551 B.n182 10.6151
R2967 B.n552 B.n551 10.6151
R2968 B.n553 B.n552 10.6151
R2969 B.n553 B.n180 10.6151
R2970 B.n557 B.n180 10.6151
R2971 B.n558 B.n557 10.6151
R2972 B.n559 B.n558 10.6151
R2973 B.n559 B.n178 10.6151
R2974 B.n563 B.n178 10.6151
R2975 B.n564 B.n563 10.6151
R2976 B.n565 B.n564 10.6151
R2977 B.n565 B.n176 10.6151
R2978 B.n569 B.n176 10.6151
R2979 B.n570 B.n569 10.6151
R2980 B.n379 B.n378 10.6151
R2981 B.n378 B.n377 10.6151
R2982 B.n377 B.n244 10.6151
R2983 B.n373 B.n244 10.6151
R2984 B.n373 B.n372 10.6151
R2985 B.n372 B.n371 10.6151
R2986 B.n371 B.n246 10.6151
R2987 B.n367 B.n246 10.6151
R2988 B.n367 B.n366 10.6151
R2989 B.n366 B.n365 10.6151
R2990 B.n365 B.n248 10.6151
R2991 B.n361 B.n248 10.6151
R2992 B.n361 B.n360 10.6151
R2993 B.n360 B.n359 10.6151
R2994 B.n359 B.n250 10.6151
R2995 B.n355 B.n250 10.6151
R2996 B.n355 B.n354 10.6151
R2997 B.n354 B.n353 10.6151
R2998 B.n353 B.n252 10.6151
R2999 B.n349 B.n252 10.6151
R3000 B.n349 B.n348 10.6151
R3001 B.n348 B.n347 10.6151
R3002 B.n347 B.n254 10.6151
R3003 B.n343 B.n254 10.6151
R3004 B.n343 B.n342 10.6151
R3005 B.n342 B.n341 10.6151
R3006 B.n341 B.n256 10.6151
R3007 B.n337 B.n256 10.6151
R3008 B.n337 B.n336 10.6151
R3009 B.n336 B.n335 10.6151
R3010 B.n335 B.n258 10.6151
R3011 B.n331 B.n258 10.6151
R3012 B.n331 B.n330 10.6151
R3013 B.n330 B.n329 10.6151
R3014 B.n329 B.n260 10.6151
R3015 B.n325 B.n260 10.6151
R3016 B.n325 B.n324 10.6151
R3017 B.n324 B.n323 10.6151
R3018 B.n323 B.n262 10.6151
R3019 B.n319 B.n262 10.6151
R3020 B.n319 B.n318 10.6151
R3021 B.n318 B.n317 10.6151
R3022 B.n317 B.n264 10.6151
R3023 B.n313 B.n264 10.6151
R3024 B.n313 B.n312 10.6151
R3025 B.n312 B.n311 10.6151
R3026 B.n311 B.n266 10.6151
R3027 B.n307 B.n266 10.6151
R3028 B.n307 B.n306 10.6151
R3029 B.n306 B.n305 10.6151
R3030 B.n305 B.n268 10.6151
R3031 B.n301 B.n268 10.6151
R3032 B.n301 B.n300 10.6151
R3033 B.n300 B.n299 10.6151
R3034 B.n299 B.n270 10.6151
R3035 B.n295 B.n270 10.6151
R3036 B.n295 B.n294 10.6151
R3037 B.n294 B.n293 10.6151
R3038 B.n293 B.n272 10.6151
R3039 B.n289 B.n272 10.6151
R3040 B.n289 B.n288 10.6151
R3041 B.n288 B.n287 10.6151
R3042 B.n287 B.n274 10.6151
R3043 B.n283 B.n274 10.6151
R3044 B.n283 B.n282 10.6151
R3045 B.n282 B.n281 10.6151
R3046 B.n281 B.n276 10.6151
R3047 B.n277 B.n276 10.6151
R3048 B.n277 B.n0 10.6151
R3049 B.n1075 B.n1 10.6151
R3050 B.n1075 B.n1074 10.6151
R3051 B.n1074 B.n1073 10.6151
R3052 B.n1073 B.n4 10.6151
R3053 B.n1069 B.n4 10.6151
R3054 B.n1069 B.n1068 10.6151
R3055 B.n1068 B.n1067 10.6151
R3056 B.n1067 B.n6 10.6151
R3057 B.n1063 B.n6 10.6151
R3058 B.n1063 B.n1062 10.6151
R3059 B.n1062 B.n1061 10.6151
R3060 B.n1061 B.n8 10.6151
R3061 B.n1057 B.n8 10.6151
R3062 B.n1057 B.n1056 10.6151
R3063 B.n1056 B.n1055 10.6151
R3064 B.n1055 B.n10 10.6151
R3065 B.n1051 B.n10 10.6151
R3066 B.n1051 B.n1050 10.6151
R3067 B.n1050 B.n1049 10.6151
R3068 B.n1049 B.n12 10.6151
R3069 B.n1045 B.n12 10.6151
R3070 B.n1045 B.n1044 10.6151
R3071 B.n1044 B.n1043 10.6151
R3072 B.n1043 B.n14 10.6151
R3073 B.n1039 B.n14 10.6151
R3074 B.n1039 B.n1038 10.6151
R3075 B.n1038 B.n1037 10.6151
R3076 B.n1037 B.n16 10.6151
R3077 B.n1033 B.n16 10.6151
R3078 B.n1033 B.n1032 10.6151
R3079 B.n1032 B.n1031 10.6151
R3080 B.n1031 B.n18 10.6151
R3081 B.n1027 B.n18 10.6151
R3082 B.n1027 B.n1026 10.6151
R3083 B.n1026 B.n1025 10.6151
R3084 B.n1025 B.n20 10.6151
R3085 B.n1021 B.n20 10.6151
R3086 B.n1021 B.n1020 10.6151
R3087 B.n1020 B.n1019 10.6151
R3088 B.n1019 B.n22 10.6151
R3089 B.n1015 B.n22 10.6151
R3090 B.n1015 B.n1014 10.6151
R3091 B.n1014 B.n1013 10.6151
R3092 B.n1013 B.n24 10.6151
R3093 B.n1009 B.n24 10.6151
R3094 B.n1009 B.n1008 10.6151
R3095 B.n1008 B.n1007 10.6151
R3096 B.n1007 B.n26 10.6151
R3097 B.n1003 B.n26 10.6151
R3098 B.n1003 B.n1002 10.6151
R3099 B.n1002 B.n1001 10.6151
R3100 B.n1001 B.n28 10.6151
R3101 B.n997 B.n28 10.6151
R3102 B.n997 B.n996 10.6151
R3103 B.n996 B.n995 10.6151
R3104 B.n995 B.n30 10.6151
R3105 B.n991 B.n30 10.6151
R3106 B.n991 B.n990 10.6151
R3107 B.n990 B.n989 10.6151
R3108 B.n989 B.n32 10.6151
R3109 B.n985 B.n32 10.6151
R3110 B.n985 B.n984 10.6151
R3111 B.n984 B.n983 10.6151
R3112 B.n983 B.n34 10.6151
R3113 B.n979 B.n34 10.6151
R3114 B.n979 B.n978 10.6151
R3115 B.n978 B.n977 10.6151
R3116 B.n977 B.n36 10.6151
R3117 B.n973 B.n36 10.6151
R3118 B.n887 B.n68 9.36635
R3119 B.n870 B.n869 9.36635
R3120 B.n468 B.n467 9.36635
R3121 B.n485 B.n206 9.36635
R3122 B.n1079 B.n0 2.81026
R3123 B.n1079 B.n1 2.81026
R3124 B.n884 B.n68 1.24928
R3125 B.n871 B.n870 1.24928
R3126 B.n469 B.n468 1.24928
R3127 B.n482 B.n206 1.24928
C0 VN VTAIL 13.962501f
C1 VDD1 VN 0.153716f
C2 VN B 1.59134f
C3 w_n5190_n4490# VN 11.024199f
C4 VDD2 VN 13.414901f
C5 VDD1 VTAIL 10.1995f
C6 VN VP 10.278099f
C7 VTAIL B 7.455979f
C8 w_n5190_n4490# VTAIL 5.53794f
C9 VDD2 VTAIL 10.2626f
C10 VTAIL VP 13.9766f
C11 VDD1 B 2.19473f
C12 w_n5190_n4490# VDD1 2.51318f
C13 w_n5190_n4490# B 13.6627f
C14 VDD1 VDD2 2.44482f
C15 VDD1 VP 13.9157f
C16 VDD2 B 2.33134f
C17 B VP 2.73406f
C18 w_n5190_n4490# VDD2 2.682f
C19 w_n5190_n4490# VP 11.7018f
C20 VDD2 VP 0.656596f
C21 VDD2 VSUBS 2.61997f
C22 VDD1 VSUBS 3.48732f
C23 VTAIL VSUBS 1.823556f
C24 VN VSUBS 8.64397f
C25 VP VSUBS 5.107593f
C26 B VSUBS 6.915059f
C27 w_n5190_n4490# VSUBS 0.285056p
C28 B.n0 VSUBS 0.004666f
C29 B.n1 VSUBS 0.004666f
C30 B.n2 VSUBS 0.007379f
C31 B.n3 VSUBS 0.007379f
C32 B.n4 VSUBS 0.007379f
C33 B.n5 VSUBS 0.007379f
C34 B.n6 VSUBS 0.007379f
C35 B.n7 VSUBS 0.007379f
C36 B.n8 VSUBS 0.007379f
C37 B.n9 VSUBS 0.007379f
C38 B.n10 VSUBS 0.007379f
C39 B.n11 VSUBS 0.007379f
C40 B.n12 VSUBS 0.007379f
C41 B.n13 VSUBS 0.007379f
C42 B.n14 VSUBS 0.007379f
C43 B.n15 VSUBS 0.007379f
C44 B.n16 VSUBS 0.007379f
C45 B.n17 VSUBS 0.007379f
C46 B.n18 VSUBS 0.007379f
C47 B.n19 VSUBS 0.007379f
C48 B.n20 VSUBS 0.007379f
C49 B.n21 VSUBS 0.007379f
C50 B.n22 VSUBS 0.007379f
C51 B.n23 VSUBS 0.007379f
C52 B.n24 VSUBS 0.007379f
C53 B.n25 VSUBS 0.007379f
C54 B.n26 VSUBS 0.007379f
C55 B.n27 VSUBS 0.007379f
C56 B.n28 VSUBS 0.007379f
C57 B.n29 VSUBS 0.007379f
C58 B.n30 VSUBS 0.007379f
C59 B.n31 VSUBS 0.007379f
C60 B.n32 VSUBS 0.007379f
C61 B.n33 VSUBS 0.007379f
C62 B.n34 VSUBS 0.007379f
C63 B.n35 VSUBS 0.007379f
C64 B.n36 VSUBS 0.007379f
C65 B.n37 VSUBS 0.018066f
C66 B.n38 VSUBS 0.007379f
C67 B.n39 VSUBS 0.007379f
C68 B.n40 VSUBS 0.007379f
C69 B.n41 VSUBS 0.007379f
C70 B.n42 VSUBS 0.007379f
C71 B.n43 VSUBS 0.007379f
C72 B.n44 VSUBS 0.007379f
C73 B.n45 VSUBS 0.007379f
C74 B.n46 VSUBS 0.007379f
C75 B.n47 VSUBS 0.007379f
C76 B.n48 VSUBS 0.007379f
C77 B.n49 VSUBS 0.007379f
C78 B.n50 VSUBS 0.007379f
C79 B.n51 VSUBS 0.007379f
C80 B.n52 VSUBS 0.007379f
C81 B.n53 VSUBS 0.007379f
C82 B.n54 VSUBS 0.007379f
C83 B.n55 VSUBS 0.007379f
C84 B.n56 VSUBS 0.007379f
C85 B.n57 VSUBS 0.007379f
C86 B.n58 VSUBS 0.007379f
C87 B.n59 VSUBS 0.007379f
C88 B.n60 VSUBS 0.007379f
C89 B.n61 VSUBS 0.007379f
C90 B.n62 VSUBS 0.007379f
C91 B.n63 VSUBS 0.007379f
C92 B.n64 VSUBS 0.007379f
C93 B.n65 VSUBS 0.007379f
C94 B.t5 VSUBS 0.360297f
C95 B.t4 VSUBS 0.409597f
C96 B.t3 VSUBS 3.29996f
C97 B.n66 VSUBS 0.655893f
C98 B.n67 VSUBS 0.347044f
C99 B.n68 VSUBS 0.017096f
C100 B.n69 VSUBS 0.007379f
C101 B.n70 VSUBS 0.007379f
C102 B.n71 VSUBS 0.007379f
C103 B.n72 VSUBS 0.007379f
C104 B.n73 VSUBS 0.007379f
C105 B.t8 VSUBS 0.360301f
C106 B.t7 VSUBS 0.4096f
C107 B.t6 VSUBS 3.29996f
C108 B.n74 VSUBS 0.65589f
C109 B.n75 VSUBS 0.34704f
C110 B.n76 VSUBS 0.007379f
C111 B.n77 VSUBS 0.007379f
C112 B.n78 VSUBS 0.007379f
C113 B.n79 VSUBS 0.007379f
C114 B.n80 VSUBS 0.007379f
C115 B.n81 VSUBS 0.007379f
C116 B.n82 VSUBS 0.007379f
C117 B.n83 VSUBS 0.007379f
C118 B.n84 VSUBS 0.007379f
C119 B.n85 VSUBS 0.007379f
C120 B.n86 VSUBS 0.007379f
C121 B.n87 VSUBS 0.007379f
C122 B.n88 VSUBS 0.007379f
C123 B.n89 VSUBS 0.007379f
C124 B.n90 VSUBS 0.007379f
C125 B.n91 VSUBS 0.007379f
C126 B.n92 VSUBS 0.007379f
C127 B.n93 VSUBS 0.007379f
C128 B.n94 VSUBS 0.007379f
C129 B.n95 VSUBS 0.007379f
C130 B.n96 VSUBS 0.007379f
C131 B.n97 VSUBS 0.007379f
C132 B.n98 VSUBS 0.007379f
C133 B.n99 VSUBS 0.007379f
C134 B.n100 VSUBS 0.007379f
C135 B.n101 VSUBS 0.007379f
C136 B.n102 VSUBS 0.007379f
C137 B.n103 VSUBS 0.007379f
C138 B.n104 VSUBS 0.017209f
C139 B.n105 VSUBS 0.007379f
C140 B.n106 VSUBS 0.007379f
C141 B.n107 VSUBS 0.007379f
C142 B.n108 VSUBS 0.007379f
C143 B.n109 VSUBS 0.007379f
C144 B.n110 VSUBS 0.007379f
C145 B.n111 VSUBS 0.007379f
C146 B.n112 VSUBS 0.007379f
C147 B.n113 VSUBS 0.007379f
C148 B.n114 VSUBS 0.007379f
C149 B.n115 VSUBS 0.007379f
C150 B.n116 VSUBS 0.007379f
C151 B.n117 VSUBS 0.007379f
C152 B.n118 VSUBS 0.007379f
C153 B.n119 VSUBS 0.007379f
C154 B.n120 VSUBS 0.007379f
C155 B.n121 VSUBS 0.007379f
C156 B.n122 VSUBS 0.007379f
C157 B.n123 VSUBS 0.007379f
C158 B.n124 VSUBS 0.007379f
C159 B.n125 VSUBS 0.007379f
C160 B.n126 VSUBS 0.007379f
C161 B.n127 VSUBS 0.007379f
C162 B.n128 VSUBS 0.007379f
C163 B.n129 VSUBS 0.007379f
C164 B.n130 VSUBS 0.007379f
C165 B.n131 VSUBS 0.007379f
C166 B.n132 VSUBS 0.007379f
C167 B.n133 VSUBS 0.007379f
C168 B.n134 VSUBS 0.007379f
C169 B.n135 VSUBS 0.007379f
C170 B.n136 VSUBS 0.007379f
C171 B.n137 VSUBS 0.007379f
C172 B.n138 VSUBS 0.007379f
C173 B.n139 VSUBS 0.007379f
C174 B.n140 VSUBS 0.007379f
C175 B.n141 VSUBS 0.007379f
C176 B.n142 VSUBS 0.007379f
C177 B.n143 VSUBS 0.007379f
C178 B.n144 VSUBS 0.007379f
C179 B.n145 VSUBS 0.007379f
C180 B.n146 VSUBS 0.007379f
C181 B.n147 VSUBS 0.007379f
C182 B.n148 VSUBS 0.007379f
C183 B.n149 VSUBS 0.007379f
C184 B.n150 VSUBS 0.007379f
C185 B.n151 VSUBS 0.007379f
C186 B.n152 VSUBS 0.007379f
C187 B.n153 VSUBS 0.007379f
C188 B.n154 VSUBS 0.007379f
C189 B.n155 VSUBS 0.007379f
C190 B.n156 VSUBS 0.007379f
C191 B.n157 VSUBS 0.007379f
C192 B.n158 VSUBS 0.007379f
C193 B.n159 VSUBS 0.007379f
C194 B.n160 VSUBS 0.007379f
C195 B.n161 VSUBS 0.007379f
C196 B.n162 VSUBS 0.007379f
C197 B.n163 VSUBS 0.007379f
C198 B.n164 VSUBS 0.007379f
C199 B.n165 VSUBS 0.007379f
C200 B.n166 VSUBS 0.007379f
C201 B.n167 VSUBS 0.007379f
C202 B.n168 VSUBS 0.007379f
C203 B.n169 VSUBS 0.007379f
C204 B.n170 VSUBS 0.007379f
C205 B.n171 VSUBS 0.007379f
C206 B.n172 VSUBS 0.007379f
C207 B.n173 VSUBS 0.007379f
C208 B.n174 VSUBS 0.007379f
C209 B.n175 VSUBS 0.018066f
C210 B.n176 VSUBS 0.007379f
C211 B.n177 VSUBS 0.007379f
C212 B.n178 VSUBS 0.007379f
C213 B.n179 VSUBS 0.007379f
C214 B.n180 VSUBS 0.007379f
C215 B.n181 VSUBS 0.007379f
C216 B.n182 VSUBS 0.007379f
C217 B.n183 VSUBS 0.007379f
C218 B.n184 VSUBS 0.007379f
C219 B.n185 VSUBS 0.007379f
C220 B.n186 VSUBS 0.007379f
C221 B.n187 VSUBS 0.007379f
C222 B.n188 VSUBS 0.007379f
C223 B.n189 VSUBS 0.007379f
C224 B.n190 VSUBS 0.007379f
C225 B.n191 VSUBS 0.007379f
C226 B.n192 VSUBS 0.007379f
C227 B.n193 VSUBS 0.007379f
C228 B.n194 VSUBS 0.007379f
C229 B.n195 VSUBS 0.007379f
C230 B.n196 VSUBS 0.007379f
C231 B.n197 VSUBS 0.007379f
C232 B.n198 VSUBS 0.007379f
C233 B.n199 VSUBS 0.007379f
C234 B.n200 VSUBS 0.007379f
C235 B.n201 VSUBS 0.007379f
C236 B.n202 VSUBS 0.007379f
C237 B.n203 VSUBS 0.007379f
C238 B.t1 VSUBS 0.360301f
C239 B.t2 VSUBS 0.4096f
C240 B.t0 VSUBS 3.29996f
C241 B.n204 VSUBS 0.65589f
C242 B.n205 VSUBS 0.34704f
C243 B.n206 VSUBS 0.017096f
C244 B.n207 VSUBS 0.007379f
C245 B.n208 VSUBS 0.007379f
C246 B.n209 VSUBS 0.007379f
C247 B.n210 VSUBS 0.007379f
C248 B.n211 VSUBS 0.007379f
C249 B.t10 VSUBS 0.360297f
C250 B.t11 VSUBS 0.409597f
C251 B.t9 VSUBS 3.29996f
C252 B.n212 VSUBS 0.655893f
C253 B.n213 VSUBS 0.347044f
C254 B.n214 VSUBS 0.007379f
C255 B.n215 VSUBS 0.007379f
C256 B.n216 VSUBS 0.007379f
C257 B.n217 VSUBS 0.007379f
C258 B.n218 VSUBS 0.007379f
C259 B.n219 VSUBS 0.007379f
C260 B.n220 VSUBS 0.007379f
C261 B.n221 VSUBS 0.007379f
C262 B.n222 VSUBS 0.007379f
C263 B.n223 VSUBS 0.007379f
C264 B.n224 VSUBS 0.007379f
C265 B.n225 VSUBS 0.007379f
C266 B.n226 VSUBS 0.007379f
C267 B.n227 VSUBS 0.007379f
C268 B.n228 VSUBS 0.007379f
C269 B.n229 VSUBS 0.007379f
C270 B.n230 VSUBS 0.007379f
C271 B.n231 VSUBS 0.007379f
C272 B.n232 VSUBS 0.007379f
C273 B.n233 VSUBS 0.007379f
C274 B.n234 VSUBS 0.007379f
C275 B.n235 VSUBS 0.007379f
C276 B.n236 VSUBS 0.007379f
C277 B.n237 VSUBS 0.007379f
C278 B.n238 VSUBS 0.007379f
C279 B.n239 VSUBS 0.007379f
C280 B.n240 VSUBS 0.007379f
C281 B.n241 VSUBS 0.007379f
C282 B.n242 VSUBS 0.018066f
C283 B.n243 VSUBS 0.007379f
C284 B.n244 VSUBS 0.007379f
C285 B.n245 VSUBS 0.007379f
C286 B.n246 VSUBS 0.007379f
C287 B.n247 VSUBS 0.007379f
C288 B.n248 VSUBS 0.007379f
C289 B.n249 VSUBS 0.007379f
C290 B.n250 VSUBS 0.007379f
C291 B.n251 VSUBS 0.007379f
C292 B.n252 VSUBS 0.007379f
C293 B.n253 VSUBS 0.007379f
C294 B.n254 VSUBS 0.007379f
C295 B.n255 VSUBS 0.007379f
C296 B.n256 VSUBS 0.007379f
C297 B.n257 VSUBS 0.007379f
C298 B.n258 VSUBS 0.007379f
C299 B.n259 VSUBS 0.007379f
C300 B.n260 VSUBS 0.007379f
C301 B.n261 VSUBS 0.007379f
C302 B.n262 VSUBS 0.007379f
C303 B.n263 VSUBS 0.007379f
C304 B.n264 VSUBS 0.007379f
C305 B.n265 VSUBS 0.007379f
C306 B.n266 VSUBS 0.007379f
C307 B.n267 VSUBS 0.007379f
C308 B.n268 VSUBS 0.007379f
C309 B.n269 VSUBS 0.007379f
C310 B.n270 VSUBS 0.007379f
C311 B.n271 VSUBS 0.007379f
C312 B.n272 VSUBS 0.007379f
C313 B.n273 VSUBS 0.007379f
C314 B.n274 VSUBS 0.007379f
C315 B.n275 VSUBS 0.007379f
C316 B.n276 VSUBS 0.007379f
C317 B.n277 VSUBS 0.007379f
C318 B.n278 VSUBS 0.007379f
C319 B.n279 VSUBS 0.007379f
C320 B.n280 VSUBS 0.007379f
C321 B.n281 VSUBS 0.007379f
C322 B.n282 VSUBS 0.007379f
C323 B.n283 VSUBS 0.007379f
C324 B.n284 VSUBS 0.007379f
C325 B.n285 VSUBS 0.007379f
C326 B.n286 VSUBS 0.007379f
C327 B.n287 VSUBS 0.007379f
C328 B.n288 VSUBS 0.007379f
C329 B.n289 VSUBS 0.007379f
C330 B.n290 VSUBS 0.007379f
C331 B.n291 VSUBS 0.007379f
C332 B.n292 VSUBS 0.007379f
C333 B.n293 VSUBS 0.007379f
C334 B.n294 VSUBS 0.007379f
C335 B.n295 VSUBS 0.007379f
C336 B.n296 VSUBS 0.007379f
C337 B.n297 VSUBS 0.007379f
C338 B.n298 VSUBS 0.007379f
C339 B.n299 VSUBS 0.007379f
C340 B.n300 VSUBS 0.007379f
C341 B.n301 VSUBS 0.007379f
C342 B.n302 VSUBS 0.007379f
C343 B.n303 VSUBS 0.007379f
C344 B.n304 VSUBS 0.007379f
C345 B.n305 VSUBS 0.007379f
C346 B.n306 VSUBS 0.007379f
C347 B.n307 VSUBS 0.007379f
C348 B.n308 VSUBS 0.007379f
C349 B.n309 VSUBS 0.007379f
C350 B.n310 VSUBS 0.007379f
C351 B.n311 VSUBS 0.007379f
C352 B.n312 VSUBS 0.007379f
C353 B.n313 VSUBS 0.007379f
C354 B.n314 VSUBS 0.007379f
C355 B.n315 VSUBS 0.007379f
C356 B.n316 VSUBS 0.007379f
C357 B.n317 VSUBS 0.007379f
C358 B.n318 VSUBS 0.007379f
C359 B.n319 VSUBS 0.007379f
C360 B.n320 VSUBS 0.007379f
C361 B.n321 VSUBS 0.007379f
C362 B.n322 VSUBS 0.007379f
C363 B.n323 VSUBS 0.007379f
C364 B.n324 VSUBS 0.007379f
C365 B.n325 VSUBS 0.007379f
C366 B.n326 VSUBS 0.007379f
C367 B.n327 VSUBS 0.007379f
C368 B.n328 VSUBS 0.007379f
C369 B.n329 VSUBS 0.007379f
C370 B.n330 VSUBS 0.007379f
C371 B.n331 VSUBS 0.007379f
C372 B.n332 VSUBS 0.007379f
C373 B.n333 VSUBS 0.007379f
C374 B.n334 VSUBS 0.007379f
C375 B.n335 VSUBS 0.007379f
C376 B.n336 VSUBS 0.007379f
C377 B.n337 VSUBS 0.007379f
C378 B.n338 VSUBS 0.007379f
C379 B.n339 VSUBS 0.007379f
C380 B.n340 VSUBS 0.007379f
C381 B.n341 VSUBS 0.007379f
C382 B.n342 VSUBS 0.007379f
C383 B.n343 VSUBS 0.007379f
C384 B.n344 VSUBS 0.007379f
C385 B.n345 VSUBS 0.007379f
C386 B.n346 VSUBS 0.007379f
C387 B.n347 VSUBS 0.007379f
C388 B.n348 VSUBS 0.007379f
C389 B.n349 VSUBS 0.007379f
C390 B.n350 VSUBS 0.007379f
C391 B.n351 VSUBS 0.007379f
C392 B.n352 VSUBS 0.007379f
C393 B.n353 VSUBS 0.007379f
C394 B.n354 VSUBS 0.007379f
C395 B.n355 VSUBS 0.007379f
C396 B.n356 VSUBS 0.007379f
C397 B.n357 VSUBS 0.007379f
C398 B.n358 VSUBS 0.007379f
C399 B.n359 VSUBS 0.007379f
C400 B.n360 VSUBS 0.007379f
C401 B.n361 VSUBS 0.007379f
C402 B.n362 VSUBS 0.007379f
C403 B.n363 VSUBS 0.007379f
C404 B.n364 VSUBS 0.007379f
C405 B.n365 VSUBS 0.007379f
C406 B.n366 VSUBS 0.007379f
C407 B.n367 VSUBS 0.007379f
C408 B.n368 VSUBS 0.007379f
C409 B.n369 VSUBS 0.007379f
C410 B.n370 VSUBS 0.007379f
C411 B.n371 VSUBS 0.007379f
C412 B.n372 VSUBS 0.007379f
C413 B.n373 VSUBS 0.007379f
C414 B.n374 VSUBS 0.007379f
C415 B.n375 VSUBS 0.007379f
C416 B.n376 VSUBS 0.007379f
C417 B.n377 VSUBS 0.007379f
C418 B.n378 VSUBS 0.007379f
C419 B.n379 VSUBS 0.016875f
C420 B.n380 VSUBS 0.016875f
C421 B.n381 VSUBS 0.018066f
C422 B.n382 VSUBS 0.007379f
C423 B.n383 VSUBS 0.007379f
C424 B.n384 VSUBS 0.007379f
C425 B.n385 VSUBS 0.007379f
C426 B.n386 VSUBS 0.007379f
C427 B.n387 VSUBS 0.007379f
C428 B.n388 VSUBS 0.007379f
C429 B.n389 VSUBS 0.007379f
C430 B.n390 VSUBS 0.007379f
C431 B.n391 VSUBS 0.007379f
C432 B.n392 VSUBS 0.007379f
C433 B.n393 VSUBS 0.007379f
C434 B.n394 VSUBS 0.007379f
C435 B.n395 VSUBS 0.007379f
C436 B.n396 VSUBS 0.007379f
C437 B.n397 VSUBS 0.007379f
C438 B.n398 VSUBS 0.007379f
C439 B.n399 VSUBS 0.007379f
C440 B.n400 VSUBS 0.007379f
C441 B.n401 VSUBS 0.007379f
C442 B.n402 VSUBS 0.007379f
C443 B.n403 VSUBS 0.007379f
C444 B.n404 VSUBS 0.007379f
C445 B.n405 VSUBS 0.007379f
C446 B.n406 VSUBS 0.007379f
C447 B.n407 VSUBS 0.007379f
C448 B.n408 VSUBS 0.007379f
C449 B.n409 VSUBS 0.007379f
C450 B.n410 VSUBS 0.007379f
C451 B.n411 VSUBS 0.007379f
C452 B.n412 VSUBS 0.007379f
C453 B.n413 VSUBS 0.007379f
C454 B.n414 VSUBS 0.007379f
C455 B.n415 VSUBS 0.007379f
C456 B.n416 VSUBS 0.007379f
C457 B.n417 VSUBS 0.007379f
C458 B.n418 VSUBS 0.007379f
C459 B.n419 VSUBS 0.007379f
C460 B.n420 VSUBS 0.007379f
C461 B.n421 VSUBS 0.007379f
C462 B.n422 VSUBS 0.007379f
C463 B.n423 VSUBS 0.007379f
C464 B.n424 VSUBS 0.007379f
C465 B.n425 VSUBS 0.007379f
C466 B.n426 VSUBS 0.007379f
C467 B.n427 VSUBS 0.007379f
C468 B.n428 VSUBS 0.007379f
C469 B.n429 VSUBS 0.007379f
C470 B.n430 VSUBS 0.007379f
C471 B.n431 VSUBS 0.007379f
C472 B.n432 VSUBS 0.007379f
C473 B.n433 VSUBS 0.007379f
C474 B.n434 VSUBS 0.007379f
C475 B.n435 VSUBS 0.007379f
C476 B.n436 VSUBS 0.007379f
C477 B.n437 VSUBS 0.007379f
C478 B.n438 VSUBS 0.007379f
C479 B.n439 VSUBS 0.007379f
C480 B.n440 VSUBS 0.007379f
C481 B.n441 VSUBS 0.007379f
C482 B.n442 VSUBS 0.007379f
C483 B.n443 VSUBS 0.007379f
C484 B.n444 VSUBS 0.007379f
C485 B.n445 VSUBS 0.007379f
C486 B.n446 VSUBS 0.007379f
C487 B.n447 VSUBS 0.007379f
C488 B.n448 VSUBS 0.007379f
C489 B.n449 VSUBS 0.007379f
C490 B.n450 VSUBS 0.007379f
C491 B.n451 VSUBS 0.007379f
C492 B.n452 VSUBS 0.007379f
C493 B.n453 VSUBS 0.007379f
C494 B.n454 VSUBS 0.007379f
C495 B.n455 VSUBS 0.007379f
C496 B.n456 VSUBS 0.007379f
C497 B.n457 VSUBS 0.007379f
C498 B.n458 VSUBS 0.007379f
C499 B.n459 VSUBS 0.007379f
C500 B.n460 VSUBS 0.007379f
C501 B.n461 VSUBS 0.007379f
C502 B.n462 VSUBS 0.007379f
C503 B.n463 VSUBS 0.007379f
C504 B.n464 VSUBS 0.007379f
C505 B.n465 VSUBS 0.007379f
C506 B.n466 VSUBS 0.007379f
C507 B.n467 VSUBS 0.006945f
C508 B.n468 VSUBS 0.017096f
C509 B.n469 VSUBS 0.004123f
C510 B.n470 VSUBS 0.007379f
C511 B.n471 VSUBS 0.007379f
C512 B.n472 VSUBS 0.007379f
C513 B.n473 VSUBS 0.007379f
C514 B.n474 VSUBS 0.007379f
C515 B.n475 VSUBS 0.007379f
C516 B.n476 VSUBS 0.007379f
C517 B.n477 VSUBS 0.007379f
C518 B.n478 VSUBS 0.007379f
C519 B.n479 VSUBS 0.007379f
C520 B.n480 VSUBS 0.007379f
C521 B.n481 VSUBS 0.007379f
C522 B.n482 VSUBS 0.004123f
C523 B.n483 VSUBS 0.007379f
C524 B.n484 VSUBS 0.007379f
C525 B.n485 VSUBS 0.006945f
C526 B.n486 VSUBS 0.007379f
C527 B.n487 VSUBS 0.007379f
C528 B.n488 VSUBS 0.007379f
C529 B.n489 VSUBS 0.007379f
C530 B.n490 VSUBS 0.007379f
C531 B.n491 VSUBS 0.007379f
C532 B.n492 VSUBS 0.007379f
C533 B.n493 VSUBS 0.007379f
C534 B.n494 VSUBS 0.007379f
C535 B.n495 VSUBS 0.007379f
C536 B.n496 VSUBS 0.007379f
C537 B.n497 VSUBS 0.007379f
C538 B.n498 VSUBS 0.007379f
C539 B.n499 VSUBS 0.007379f
C540 B.n500 VSUBS 0.007379f
C541 B.n501 VSUBS 0.007379f
C542 B.n502 VSUBS 0.007379f
C543 B.n503 VSUBS 0.007379f
C544 B.n504 VSUBS 0.007379f
C545 B.n505 VSUBS 0.007379f
C546 B.n506 VSUBS 0.007379f
C547 B.n507 VSUBS 0.007379f
C548 B.n508 VSUBS 0.007379f
C549 B.n509 VSUBS 0.007379f
C550 B.n510 VSUBS 0.007379f
C551 B.n511 VSUBS 0.007379f
C552 B.n512 VSUBS 0.007379f
C553 B.n513 VSUBS 0.007379f
C554 B.n514 VSUBS 0.007379f
C555 B.n515 VSUBS 0.007379f
C556 B.n516 VSUBS 0.007379f
C557 B.n517 VSUBS 0.007379f
C558 B.n518 VSUBS 0.007379f
C559 B.n519 VSUBS 0.007379f
C560 B.n520 VSUBS 0.007379f
C561 B.n521 VSUBS 0.007379f
C562 B.n522 VSUBS 0.007379f
C563 B.n523 VSUBS 0.007379f
C564 B.n524 VSUBS 0.007379f
C565 B.n525 VSUBS 0.007379f
C566 B.n526 VSUBS 0.007379f
C567 B.n527 VSUBS 0.007379f
C568 B.n528 VSUBS 0.007379f
C569 B.n529 VSUBS 0.007379f
C570 B.n530 VSUBS 0.007379f
C571 B.n531 VSUBS 0.007379f
C572 B.n532 VSUBS 0.007379f
C573 B.n533 VSUBS 0.007379f
C574 B.n534 VSUBS 0.007379f
C575 B.n535 VSUBS 0.007379f
C576 B.n536 VSUBS 0.007379f
C577 B.n537 VSUBS 0.007379f
C578 B.n538 VSUBS 0.007379f
C579 B.n539 VSUBS 0.007379f
C580 B.n540 VSUBS 0.007379f
C581 B.n541 VSUBS 0.007379f
C582 B.n542 VSUBS 0.007379f
C583 B.n543 VSUBS 0.007379f
C584 B.n544 VSUBS 0.007379f
C585 B.n545 VSUBS 0.007379f
C586 B.n546 VSUBS 0.007379f
C587 B.n547 VSUBS 0.007379f
C588 B.n548 VSUBS 0.007379f
C589 B.n549 VSUBS 0.007379f
C590 B.n550 VSUBS 0.007379f
C591 B.n551 VSUBS 0.007379f
C592 B.n552 VSUBS 0.007379f
C593 B.n553 VSUBS 0.007379f
C594 B.n554 VSUBS 0.007379f
C595 B.n555 VSUBS 0.007379f
C596 B.n556 VSUBS 0.007379f
C597 B.n557 VSUBS 0.007379f
C598 B.n558 VSUBS 0.007379f
C599 B.n559 VSUBS 0.007379f
C600 B.n560 VSUBS 0.007379f
C601 B.n561 VSUBS 0.007379f
C602 B.n562 VSUBS 0.007379f
C603 B.n563 VSUBS 0.007379f
C604 B.n564 VSUBS 0.007379f
C605 B.n565 VSUBS 0.007379f
C606 B.n566 VSUBS 0.007379f
C607 B.n567 VSUBS 0.007379f
C608 B.n568 VSUBS 0.007379f
C609 B.n569 VSUBS 0.007379f
C610 B.n570 VSUBS 0.018066f
C611 B.n571 VSUBS 0.016875f
C612 B.n572 VSUBS 0.016875f
C613 B.n573 VSUBS 0.007379f
C614 B.n574 VSUBS 0.007379f
C615 B.n575 VSUBS 0.007379f
C616 B.n576 VSUBS 0.007379f
C617 B.n577 VSUBS 0.007379f
C618 B.n578 VSUBS 0.007379f
C619 B.n579 VSUBS 0.007379f
C620 B.n580 VSUBS 0.007379f
C621 B.n581 VSUBS 0.007379f
C622 B.n582 VSUBS 0.007379f
C623 B.n583 VSUBS 0.007379f
C624 B.n584 VSUBS 0.007379f
C625 B.n585 VSUBS 0.007379f
C626 B.n586 VSUBS 0.007379f
C627 B.n587 VSUBS 0.007379f
C628 B.n588 VSUBS 0.007379f
C629 B.n589 VSUBS 0.007379f
C630 B.n590 VSUBS 0.007379f
C631 B.n591 VSUBS 0.007379f
C632 B.n592 VSUBS 0.007379f
C633 B.n593 VSUBS 0.007379f
C634 B.n594 VSUBS 0.007379f
C635 B.n595 VSUBS 0.007379f
C636 B.n596 VSUBS 0.007379f
C637 B.n597 VSUBS 0.007379f
C638 B.n598 VSUBS 0.007379f
C639 B.n599 VSUBS 0.007379f
C640 B.n600 VSUBS 0.007379f
C641 B.n601 VSUBS 0.007379f
C642 B.n602 VSUBS 0.007379f
C643 B.n603 VSUBS 0.007379f
C644 B.n604 VSUBS 0.007379f
C645 B.n605 VSUBS 0.007379f
C646 B.n606 VSUBS 0.007379f
C647 B.n607 VSUBS 0.007379f
C648 B.n608 VSUBS 0.007379f
C649 B.n609 VSUBS 0.007379f
C650 B.n610 VSUBS 0.007379f
C651 B.n611 VSUBS 0.007379f
C652 B.n612 VSUBS 0.007379f
C653 B.n613 VSUBS 0.007379f
C654 B.n614 VSUBS 0.007379f
C655 B.n615 VSUBS 0.007379f
C656 B.n616 VSUBS 0.007379f
C657 B.n617 VSUBS 0.007379f
C658 B.n618 VSUBS 0.007379f
C659 B.n619 VSUBS 0.007379f
C660 B.n620 VSUBS 0.007379f
C661 B.n621 VSUBS 0.007379f
C662 B.n622 VSUBS 0.007379f
C663 B.n623 VSUBS 0.007379f
C664 B.n624 VSUBS 0.007379f
C665 B.n625 VSUBS 0.007379f
C666 B.n626 VSUBS 0.007379f
C667 B.n627 VSUBS 0.007379f
C668 B.n628 VSUBS 0.007379f
C669 B.n629 VSUBS 0.007379f
C670 B.n630 VSUBS 0.007379f
C671 B.n631 VSUBS 0.007379f
C672 B.n632 VSUBS 0.007379f
C673 B.n633 VSUBS 0.007379f
C674 B.n634 VSUBS 0.007379f
C675 B.n635 VSUBS 0.007379f
C676 B.n636 VSUBS 0.007379f
C677 B.n637 VSUBS 0.007379f
C678 B.n638 VSUBS 0.007379f
C679 B.n639 VSUBS 0.007379f
C680 B.n640 VSUBS 0.007379f
C681 B.n641 VSUBS 0.007379f
C682 B.n642 VSUBS 0.007379f
C683 B.n643 VSUBS 0.007379f
C684 B.n644 VSUBS 0.007379f
C685 B.n645 VSUBS 0.007379f
C686 B.n646 VSUBS 0.007379f
C687 B.n647 VSUBS 0.007379f
C688 B.n648 VSUBS 0.007379f
C689 B.n649 VSUBS 0.007379f
C690 B.n650 VSUBS 0.007379f
C691 B.n651 VSUBS 0.007379f
C692 B.n652 VSUBS 0.007379f
C693 B.n653 VSUBS 0.007379f
C694 B.n654 VSUBS 0.007379f
C695 B.n655 VSUBS 0.007379f
C696 B.n656 VSUBS 0.007379f
C697 B.n657 VSUBS 0.007379f
C698 B.n658 VSUBS 0.007379f
C699 B.n659 VSUBS 0.007379f
C700 B.n660 VSUBS 0.007379f
C701 B.n661 VSUBS 0.007379f
C702 B.n662 VSUBS 0.007379f
C703 B.n663 VSUBS 0.007379f
C704 B.n664 VSUBS 0.007379f
C705 B.n665 VSUBS 0.007379f
C706 B.n666 VSUBS 0.007379f
C707 B.n667 VSUBS 0.007379f
C708 B.n668 VSUBS 0.007379f
C709 B.n669 VSUBS 0.007379f
C710 B.n670 VSUBS 0.007379f
C711 B.n671 VSUBS 0.007379f
C712 B.n672 VSUBS 0.007379f
C713 B.n673 VSUBS 0.007379f
C714 B.n674 VSUBS 0.007379f
C715 B.n675 VSUBS 0.007379f
C716 B.n676 VSUBS 0.007379f
C717 B.n677 VSUBS 0.007379f
C718 B.n678 VSUBS 0.007379f
C719 B.n679 VSUBS 0.007379f
C720 B.n680 VSUBS 0.007379f
C721 B.n681 VSUBS 0.007379f
C722 B.n682 VSUBS 0.007379f
C723 B.n683 VSUBS 0.007379f
C724 B.n684 VSUBS 0.007379f
C725 B.n685 VSUBS 0.007379f
C726 B.n686 VSUBS 0.007379f
C727 B.n687 VSUBS 0.007379f
C728 B.n688 VSUBS 0.007379f
C729 B.n689 VSUBS 0.007379f
C730 B.n690 VSUBS 0.007379f
C731 B.n691 VSUBS 0.007379f
C732 B.n692 VSUBS 0.007379f
C733 B.n693 VSUBS 0.007379f
C734 B.n694 VSUBS 0.007379f
C735 B.n695 VSUBS 0.007379f
C736 B.n696 VSUBS 0.007379f
C737 B.n697 VSUBS 0.007379f
C738 B.n698 VSUBS 0.007379f
C739 B.n699 VSUBS 0.007379f
C740 B.n700 VSUBS 0.007379f
C741 B.n701 VSUBS 0.007379f
C742 B.n702 VSUBS 0.007379f
C743 B.n703 VSUBS 0.007379f
C744 B.n704 VSUBS 0.007379f
C745 B.n705 VSUBS 0.007379f
C746 B.n706 VSUBS 0.007379f
C747 B.n707 VSUBS 0.007379f
C748 B.n708 VSUBS 0.007379f
C749 B.n709 VSUBS 0.007379f
C750 B.n710 VSUBS 0.007379f
C751 B.n711 VSUBS 0.007379f
C752 B.n712 VSUBS 0.007379f
C753 B.n713 VSUBS 0.007379f
C754 B.n714 VSUBS 0.007379f
C755 B.n715 VSUBS 0.007379f
C756 B.n716 VSUBS 0.007379f
C757 B.n717 VSUBS 0.007379f
C758 B.n718 VSUBS 0.007379f
C759 B.n719 VSUBS 0.007379f
C760 B.n720 VSUBS 0.007379f
C761 B.n721 VSUBS 0.007379f
C762 B.n722 VSUBS 0.007379f
C763 B.n723 VSUBS 0.007379f
C764 B.n724 VSUBS 0.007379f
C765 B.n725 VSUBS 0.007379f
C766 B.n726 VSUBS 0.007379f
C767 B.n727 VSUBS 0.007379f
C768 B.n728 VSUBS 0.007379f
C769 B.n729 VSUBS 0.007379f
C770 B.n730 VSUBS 0.007379f
C771 B.n731 VSUBS 0.007379f
C772 B.n732 VSUBS 0.007379f
C773 B.n733 VSUBS 0.007379f
C774 B.n734 VSUBS 0.007379f
C775 B.n735 VSUBS 0.007379f
C776 B.n736 VSUBS 0.007379f
C777 B.n737 VSUBS 0.007379f
C778 B.n738 VSUBS 0.007379f
C779 B.n739 VSUBS 0.007379f
C780 B.n740 VSUBS 0.007379f
C781 B.n741 VSUBS 0.007379f
C782 B.n742 VSUBS 0.007379f
C783 B.n743 VSUBS 0.007379f
C784 B.n744 VSUBS 0.007379f
C785 B.n745 VSUBS 0.007379f
C786 B.n746 VSUBS 0.007379f
C787 B.n747 VSUBS 0.007379f
C788 B.n748 VSUBS 0.007379f
C789 B.n749 VSUBS 0.007379f
C790 B.n750 VSUBS 0.007379f
C791 B.n751 VSUBS 0.007379f
C792 B.n752 VSUBS 0.007379f
C793 B.n753 VSUBS 0.007379f
C794 B.n754 VSUBS 0.007379f
C795 B.n755 VSUBS 0.007379f
C796 B.n756 VSUBS 0.007379f
C797 B.n757 VSUBS 0.007379f
C798 B.n758 VSUBS 0.007379f
C799 B.n759 VSUBS 0.007379f
C800 B.n760 VSUBS 0.007379f
C801 B.n761 VSUBS 0.007379f
C802 B.n762 VSUBS 0.007379f
C803 B.n763 VSUBS 0.007379f
C804 B.n764 VSUBS 0.007379f
C805 B.n765 VSUBS 0.007379f
C806 B.n766 VSUBS 0.007379f
C807 B.n767 VSUBS 0.007379f
C808 B.n768 VSUBS 0.007379f
C809 B.n769 VSUBS 0.007379f
C810 B.n770 VSUBS 0.007379f
C811 B.n771 VSUBS 0.007379f
C812 B.n772 VSUBS 0.007379f
C813 B.n773 VSUBS 0.007379f
C814 B.n774 VSUBS 0.007379f
C815 B.n775 VSUBS 0.007379f
C816 B.n776 VSUBS 0.007379f
C817 B.n777 VSUBS 0.007379f
C818 B.n778 VSUBS 0.007379f
C819 B.n779 VSUBS 0.007379f
C820 B.n780 VSUBS 0.007379f
C821 B.n781 VSUBS 0.017731f
C822 B.n782 VSUBS 0.016875f
C823 B.n783 VSUBS 0.018066f
C824 B.n784 VSUBS 0.007379f
C825 B.n785 VSUBS 0.007379f
C826 B.n786 VSUBS 0.007379f
C827 B.n787 VSUBS 0.007379f
C828 B.n788 VSUBS 0.007379f
C829 B.n789 VSUBS 0.007379f
C830 B.n790 VSUBS 0.007379f
C831 B.n791 VSUBS 0.007379f
C832 B.n792 VSUBS 0.007379f
C833 B.n793 VSUBS 0.007379f
C834 B.n794 VSUBS 0.007379f
C835 B.n795 VSUBS 0.007379f
C836 B.n796 VSUBS 0.007379f
C837 B.n797 VSUBS 0.007379f
C838 B.n798 VSUBS 0.007379f
C839 B.n799 VSUBS 0.007379f
C840 B.n800 VSUBS 0.007379f
C841 B.n801 VSUBS 0.007379f
C842 B.n802 VSUBS 0.007379f
C843 B.n803 VSUBS 0.007379f
C844 B.n804 VSUBS 0.007379f
C845 B.n805 VSUBS 0.007379f
C846 B.n806 VSUBS 0.007379f
C847 B.n807 VSUBS 0.007379f
C848 B.n808 VSUBS 0.007379f
C849 B.n809 VSUBS 0.007379f
C850 B.n810 VSUBS 0.007379f
C851 B.n811 VSUBS 0.007379f
C852 B.n812 VSUBS 0.007379f
C853 B.n813 VSUBS 0.007379f
C854 B.n814 VSUBS 0.007379f
C855 B.n815 VSUBS 0.007379f
C856 B.n816 VSUBS 0.007379f
C857 B.n817 VSUBS 0.007379f
C858 B.n818 VSUBS 0.007379f
C859 B.n819 VSUBS 0.007379f
C860 B.n820 VSUBS 0.007379f
C861 B.n821 VSUBS 0.007379f
C862 B.n822 VSUBS 0.007379f
C863 B.n823 VSUBS 0.007379f
C864 B.n824 VSUBS 0.007379f
C865 B.n825 VSUBS 0.007379f
C866 B.n826 VSUBS 0.007379f
C867 B.n827 VSUBS 0.007379f
C868 B.n828 VSUBS 0.007379f
C869 B.n829 VSUBS 0.007379f
C870 B.n830 VSUBS 0.007379f
C871 B.n831 VSUBS 0.007379f
C872 B.n832 VSUBS 0.007379f
C873 B.n833 VSUBS 0.007379f
C874 B.n834 VSUBS 0.007379f
C875 B.n835 VSUBS 0.007379f
C876 B.n836 VSUBS 0.007379f
C877 B.n837 VSUBS 0.007379f
C878 B.n838 VSUBS 0.007379f
C879 B.n839 VSUBS 0.007379f
C880 B.n840 VSUBS 0.007379f
C881 B.n841 VSUBS 0.007379f
C882 B.n842 VSUBS 0.007379f
C883 B.n843 VSUBS 0.007379f
C884 B.n844 VSUBS 0.007379f
C885 B.n845 VSUBS 0.007379f
C886 B.n846 VSUBS 0.007379f
C887 B.n847 VSUBS 0.007379f
C888 B.n848 VSUBS 0.007379f
C889 B.n849 VSUBS 0.007379f
C890 B.n850 VSUBS 0.007379f
C891 B.n851 VSUBS 0.007379f
C892 B.n852 VSUBS 0.007379f
C893 B.n853 VSUBS 0.007379f
C894 B.n854 VSUBS 0.007379f
C895 B.n855 VSUBS 0.007379f
C896 B.n856 VSUBS 0.007379f
C897 B.n857 VSUBS 0.007379f
C898 B.n858 VSUBS 0.007379f
C899 B.n859 VSUBS 0.007379f
C900 B.n860 VSUBS 0.007379f
C901 B.n861 VSUBS 0.007379f
C902 B.n862 VSUBS 0.007379f
C903 B.n863 VSUBS 0.007379f
C904 B.n864 VSUBS 0.007379f
C905 B.n865 VSUBS 0.007379f
C906 B.n866 VSUBS 0.007379f
C907 B.n867 VSUBS 0.007379f
C908 B.n868 VSUBS 0.007379f
C909 B.n869 VSUBS 0.006945f
C910 B.n870 VSUBS 0.017096f
C911 B.n871 VSUBS 0.004123f
C912 B.n872 VSUBS 0.007379f
C913 B.n873 VSUBS 0.007379f
C914 B.n874 VSUBS 0.007379f
C915 B.n875 VSUBS 0.007379f
C916 B.n876 VSUBS 0.007379f
C917 B.n877 VSUBS 0.007379f
C918 B.n878 VSUBS 0.007379f
C919 B.n879 VSUBS 0.007379f
C920 B.n880 VSUBS 0.007379f
C921 B.n881 VSUBS 0.007379f
C922 B.n882 VSUBS 0.007379f
C923 B.n883 VSUBS 0.007379f
C924 B.n884 VSUBS 0.004123f
C925 B.n885 VSUBS 0.007379f
C926 B.n886 VSUBS 0.007379f
C927 B.n887 VSUBS 0.006945f
C928 B.n888 VSUBS 0.007379f
C929 B.n889 VSUBS 0.007379f
C930 B.n890 VSUBS 0.007379f
C931 B.n891 VSUBS 0.007379f
C932 B.n892 VSUBS 0.007379f
C933 B.n893 VSUBS 0.007379f
C934 B.n894 VSUBS 0.007379f
C935 B.n895 VSUBS 0.007379f
C936 B.n896 VSUBS 0.007379f
C937 B.n897 VSUBS 0.007379f
C938 B.n898 VSUBS 0.007379f
C939 B.n899 VSUBS 0.007379f
C940 B.n900 VSUBS 0.007379f
C941 B.n901 VSUBS 0.007379f
C942 B.n902 VSUBS 0.007379f
C943 B.n903 VSUBS 0.007379f
C944 B.n904 VSUBS 0.007379f
C945 B.n905 VSUBS 0.007379f
C946 B.n906 VSUBS 0.007379f
C947 B.n907 VSUBS 0.007379f
C948 B.n908 VSUBS 0.007379f
C949 B.n909 VSUBS 0.007379f
C950 B.n910 VSUBS 0.007379f
C951 B.n911 VSUBS 0.007379f
C952 B.n912 VSUBS 0.007379f
C953 B.n913 VSUBS 0.007379f
C954 B.n914 VSUBS 0.007379f
C955 B.n915 VSUBS 0.007379f
C956 B.n916 VSUBS 0.007379f
C957 B.n917 VSUBS 0.007379f
C958 B.n918 VSUBS 0.007379f
C959 B.n919 VSUBS 0.007379f
C960 B.n920 VSUBS 0.007379f
C961 B.n921 VSUBS 0.007379f
C962 B.n922 VSUBS 0.007379f
C963 B.n923 VSUBS 0.007379f
C964 B.n924 VSUBS 0.007379f
C965 B.n925 VSUBS 0.007379f
C966 B.n926 VSUBS 0.007379f
C967 B.n927 VSUBS 0.007379f
C968 B.n928 VSUBS 0.007379f
C969 B.n929 VSUBS 0.007379f
C970 B.n930 VSUBS 0.007379f
C971 B.n931 VSUBS 0.007379f
C972 B.n932 VSUBS 0.007379f
C973 B.n933 VSUBS 0.007379f
C974 B.n934 VSUBS 0.007379f
C975 B.n935 VSUBS 0.007379f
C976 B.n936 VSUBS 0.007379f
C977 B.n937 VSUBS 0.007379f
C978 B.n938 VSUBS 0.007379f
C979 B.n939 VSUBS 0.007379f
C980 B.n940 VSUBS 0.007379f
C981 B.n941 VSUBS 0.007379f
C982 B.n942 VSUBS 0.007379f
C983 B.n943 VSUBS 0.007379f
C984 B.n944 VSUBS 0.007379f
C985 B.n945 VSUBS 0.007379f
C986 B.n946 VSUBS 0.007379f
C987 B.n947 VSUBS 0.007379f
C988 B.n948 VSUBS 0.007379f
C989 B.n949 VSUBS 0.007379f
C990 B.n950 VSUBS 0.007379f
C991 B.n951 VSUBS 0.007379f
C992 B.n952 VSUBS 0.007379f
C993 B.n953 VSUBS 0.007379f
C994 B.n954 VSUBS 0.007379f
C995 B.n955 VSUBS 0.007379f
C996 B.n956 VSUBS 0.007379f
C997 B.n957 VSUBS 0.007379f
C998 B.n958 VSUBS 0.007379f
C999 B.n959 VSUBS 0.007379f
C1000 B.n960 VSUBS 0.007379f
C1001 B.n961 VSUBS 0.007379f
C1002 B.n962 VSUBS 0.007379f
C1003 B.n963 VSUBS 0.007379f
C1004 B.n964 VSUBS 0.007379f
C1005 B.n965 VSUBS 0.007379f
C1006 B.n966 VSUBS 0.007379f
C1007 B.n967 VSUBS 0.007379f
C1008 B.n968 VSUBS 0.007379f
C1009 B.n969 VSUBS 0.007379f
C1010 B.n970 VSUBS 0.007379f
C1011 B.n971 VSUBS 0.007379f
C1012 B.n972 VSUBS 0.018066f
C1013 B.n973 VSUBS 0.016875f
C1014 B.n974 VSUBS 0.016875f
C1015 B.n975 VSUBS 0.007379f
C1016 B.n976 VSUBS 0.007379f
C1017 B.n977 VSUBS 0.007379f
C1018 B.n978 VSUBS 0.007379f
C1019 B.n979 VSUBS 0.007379f
C1020 B.n980 VSUBS 0.007379f
C1021 B.n981 VSUBS 0.007379f
C1022 B.n982 VSUBS 0.007379f
C1023 B.n983 VSUBS 0.007379f
C1024 B.n984 VSUBS 0.007379f
C1025 B.n985 VSUBS 0.007379f
C1026 B.n986 VSUBS 0.007379f
C1027 B.n987 VSUBS 0.007379f
C1028 B.n988 VSUBS 0.007379f
C1029 B.n989 VSUBS 0.007379f
C1030 B.n990 VSUBS 0.007379f
C1031 B.n991 VSUBS 0.007379f
C1032 B.n992 VSUBS 0.007379f
C1033 B.n993 VSUBS 0.007379f
C1034 B.n994 VSUBS 0.007379f
C1035 B.n995 VSUBS 0.007379f
C1036 B.n996 VSUBS 0.007379f
C1037 B.n997 VSUBS 0.007379f
C1038 B.n998 VSUBS 0.007379f
C1039 B.n999 VSUBS 0.007379f
C1040 B.n1000 VSUBS 0.007379f
C1041 B.n1001 VSUBS 0.007379f
C1042 B.n1002 VSUBS 0.007379f
C1043 B.n1003 VSUBS 0.007379f
C1044 B.n1004 VSUBS 0.007379f
C1045 B.n1005 VSUBS 0.007379f
C1046 B.n1006 VSUBS 0.007379f
C1047 B.n1007 VSUBS 0.007379f
C1048 B.n1008 VSUBS 0.007379f
C1049 B.n1009 VSUBS 0.007379f
C1050 B.n1010 VSUBS 0.007379f
C1051 B.n1011 VSUBS 0.007379f
C1052 B.n1012 VSUBS 0.007379f
C1053 B.n1013 VSUBS 0.007379f
C1054 B.n1014 VSUBS 0.007379f
C1055 B.n1015 VSUBS 0.007379f
C1056 B.n1016 VSUBS 0.007379f
C1057 B.n1017 VSUBS 0.007379f
C1058 B.n1018 VSUBS 0.007379f
C1059 B.n1019 VSUBS 0.007379f
C1060 B.n1020 VSUBS 0.007379f
C1061 B.n1021 VSUBS 0.007379f
C1062 B.n1022 VSUBS 0.007379f
C1063 B.n1023 VSUBS 0.007379f
C1064 B.n1024 VSUBS 0.007379f
C1065 B.n1025 VSUBS 0.007379f
C1066 B.n1026 VSUBS 0.007379f
C1067 B.n1027 VSUBS 0.007379f
C1068 B.n1028 VSUBS 0.007379f
C1069 B.n1029 VSUBS 0.007379f
C1070 B.n1030 VSUBS 0.007379f
C1071 B.n1031 VSUBS 0.007379f
C1072 B.n1032 VSUBS 0.007379f
C1073 B.n1033 VSUBS 0.007379f
C1074 B.n1034 VSUBS 0.007379f
C1075 B.n1035 VSUBS 0.007379f
C1076 B.n1036 VSUBS 0.007379f
C1077 B.n1037 VSUBS 0.007379f
C1078 B.n1038 VSUBS 0.007379f
C1079 B.n1039 VSUBS 0.007379f
C1080 B.n1040 VSUBS 0.007379f
C1081 B.n1041 VSUBS 0.007379f
C1082 B.n1042 VSUBS 0.007379f
C1083 B.n1043 VSUBS 0.007379f
C1084 B.n1044 VSUBS 0.007379f
C1085 B.n1045 VSUBS 0.007379f
C1086 B.n1046 VSUBS 0.007379f
C1087 B.n1047 VSUBS 0.007379f
C1088 B.n1048 VSUBS 0.007379f
C1089 B.n1049 VSUBS 0.007379f
C1090 B.n1050 VSUBS 0.007379f
C1091 B.n1051 VSUBS 0.007379f
C1092 B.n1052 VSUBS 0.007379f
C1093 B.n1053 VSUBS 0.007379f
C1094 B.n1054 VSUBS 0.007379f
C1095 B.n1055 VSUBS 0.007379f
C1096 B.n1056 VSUBS 0.007379f
C1097 B.n1057 VSUBS 0.007379f
C1098 B.n1058 VSUBS 0.007379f
C1099 B.n1059 VSUBS 0.007379f
C1100 B.n1060 VSUBS 0.007379f
C1101 B.n1061 VSUBS 0.007379f
C1102 B.n1062 VSUBS 0.007379f
C1103 B.n1063 VSUBS 0.007379f
C1104 B.n1064 VSUBS 0.007379f
C1105 B.n1065 VSUBS 0.007379f
C1106 B.n1066 VSUBS 0.007379f
C1107 B.n1067 VSUBS 0.007379f
C1108 B.n1068 VSUBS 0.007379f
C1109 B.n1069 VSUBS 0.007379f
C1110 B.n1070 VSUBS 0.007379f
C1111 B.n1071 VSUBS 0.007379f
C1112 B.n1072 VSUBS 0.007379f
C1113 B.n1073 VSUBS 0.007379f
C1114 B.n1074 VSUBS 0.007379f
C1115 B.n1075 VSUBS 0.007379f
C1116 B.n1076 VSUBS 0.007379f
C1117 B.n1077 VSUBS 0.007379f
C1118 B.n1078 VSUBS 0.007379f
C1119 B.n1079 VSUBS 0.016708f
C1120 VDD1.t7 VSUBS 0.438955f
C1121 VDD1.t2 VSUBS 0.438955f
C1122 VDD1.n0 VSUBS 3.67619f
C1123 VDD1.t5 VSUBS 0.438955f
C1124 VDD1.t3 VSUBS 0.438955f
C1125 VDD1.n1 VSUBS 3.6741f
C1126 VDD1.t4 VSUBS 0.438955f
C1127 VDD1.t6 VSUBS 0.438955f
C1128 VDD1.n2 VSUBS 3.6741f
C1129 VDD1.n3 VSUBS 6.28363f
C1130 VDD1.t0 VSUBS 0.438955f
C1131 VDD1.t1 VSUBS 0.438955f
C1132 VDD1.n4 VSUBS 3.64556f
C1133 VDD1.n5 VSUBS 5.21098f
C1134 VP.t1 VSUBS 4.22541f
C1135 VP.n0 VSUBS 1.54365f
C1136 VP.n1 VSUBS 0.022435f
C1137 VP.n2 VSUBS 0.045124f
C1138 VP.n3 VSUBS 0.022435f
C1139 VP.n4 VSUBS 0.041813f
C1140 VP.n5 VSUBS 0.022435f
C1141 VP.t3 VSUBS 4.22541f
C1142 VP.n6 VSUBS 0.041813f
C1143 VP.n7 VSUBS 0.022435f
C1144 VP.n8 VSUBS 0.041813f
C1145 VP.n9 VSUBS 0.022435f
C1146 VP.t4 VSUBS 4.22541f
C1147 VP.n10 VSUBS 0.041813f
C1148 VP.n11 VSUBS 0.022435f
C1149 VP.n12 VSUBS 0.041813f
C1150 VP.n13 VSUBS 0.036209f
C1151 VP.t2 VSUBS 4.22541f
C1152 VP.t6 VSUBS 4.22541f
C1153 VP.n14 VSUBS 1.54365f
C1154 VP.n15 VSUBS 0.022435f
C1155 VP.n16 VSUBS 0.045124f
C1156 VP.n17 VSUBS 0.022435f
C1157 VP.n18 VSUBS 0.041813f
C1158 VP.n19 VSUBS 0.022435f
C1159 VP.t7 VSUBS 4.22541f
C1160 VP.n20 VSUBS 0.041813f
C1161 VP.n21 VSUBS 0.022435f
C1162 VP.n22 VSUBS 0.041813f
C1163 VP.t0 VSUBS 4.60672f
C1164 VP.n23 VSUBS 1.46871f
C1165 VP.t5 VSUBS 4.22541f
C1166 VP.n24 VSUBS 1.54225f
C1167 VP.n25 VSUBS 0.036032f
C1168 VP.n26 VSUBS 0.290393f
C1169 VP.n27 VSUBS 0.022435f
C1170 VP.n28 VSUBS 0.022435f
C1171 VP.n29 VSUBS 0.041813f
C1172 VP.n30 VSUBS 0.03275f
C1173 VP.n31 VSUBS 0.03275f
C1174 VP.n32 VSUBS 0.022435f
C1175 VP.n33 VSUBS 0.022435f
C1176 VP.n34 VSUBS 0.022435f
C1177 VP.n35 VSUBS 0.041813f
C1178 VP.n36 VSUBS 0.036032f
C1179 VP.n37 VSUBS 1.45629f
C1180 VP.n38 VSUBS 0.026949f
C1181 VP.n39 VSUBS 0.022435f
C1182 VP.n40 VSUBS 0.022435f
C1183 VP.n41 VSUBS 0.022435f
C1184 VP.n42 VSUBS 0.041813f
C1185 VP.n43 VSUBS 0.043792f
C1186 VP.n44 VSUBS 0.018397f
C1187 VP.n45 VSUBS 0.022435f
C1188 VP.n46 VSUBS 0.022435f
C1189 VP.n47 VSUBS 0.022435f
C1190 VP.n48 VSUBS 0.041813f
C1191 VP.n49 VSUBS 0.041813f
C1192 VP.n50 VSUBS 0.024472f
C1193 VP.n51 VSUBS 0.036209f
C1194 VP.n52 VSUBS 1.70564f
C1195 VP.n53 VSUBS 1.71881f
C1196 VP.n54 VSUBS 1.54365f
C1197 VP.n55 VSUBS 0.024472f
C1198 VP.n56 VSUBS 0.041813f
C1199 VP.n57 VSUBS 0.022435f
C1200 VP.n58 VSUBS 0.022435f
C1201 VP.n59 VSUBS 0.022435f
C1202 VP.n60 VSUBS 0.045124f
C1203 VP.n61 VSUBS 0.018397f
C1204 VP.n62 VSUBS 0.043792f
C1205 VP.n63 VSUBS 0.022435f
C1206 VP.n64 VSUBS 0.022435f
C1207 VP.n65 VSUBS 0.022435f
C1208 VP.n66 VSUBS 0.041813f
C1209 VP.n67 VSUBS 0.026949f
C1210 VP.n68 VSUBS 1.45629f
C1211 VP.n69 VSUBS 0.036032f
C1212 VP.n70 VSUBS 0.022435f
C1213 VP.n71 VSUBS 0.022435f
C1214 VP.n72 VSUBS 0.022435f
C1215 VP.n73 VSUBS 0.041813f
C1216 VP.n74 VSUBS 0.03275f
C1217 VP.n75 VSUBS 0.03275f
C1218 VP.n76 VSUBS 0.022435f
C1219 VP.n77 VSUBS 0.022435f
C1220 VP.n78 VSUBS 0.022435f
C1221 VP.n79 VSUBS 0.041813f
C1222 VP.n80 VSUBS 0.036032f
C1223 VP.n81 VSUBS 1.45629f
C1224 VP.n82 VSUBS 0.026949f
C1225 VP.n83 VSUBS 0.022435f
C1226 VP.n84 VSUBS 0.022435f
C1227 VP.n85 VSUBS 0.022435f
C1228 VP.n86 VSUBS 0.041813f
C1229 VP.n87 VSUBS 0.043792f
C1230 VP.n88 VSUBS 0.018397f
C1231 VP.n89 VSUBS 0.022435f
C1232 VP.n90 VSUBS 0.022435f
C1233 VP.n91 VSUBS 0.022435f
C1234 VP.n92 VSUBS 0.041813f
C1235 VP.n93 VSUBS 0.041813f
C1236 VP.n94 VSUBS 0.024472f
C1237 VP.n95 VSUBS 0.036209f
C1238 VP.n96 VSUBS 0.069325f
C1239 VTAIL.t9 VSUBS 0.341156f
C1240 VTAIL.t14 VSUBS 0.341156f
C1241 VTAIL.n0 VSUBS 2.68824f
C1242 VTAIL.n1 VSUBS 0.878942f
C1243 VTAIL.n2 VSUBS 0.027354f
C1244 VTAIL.n3 VSUBS 0.024515f
C1245 VTAIL.n4 VSUBS 0.013174f
C1246 VTAIL.n5 VSUBS 0.031137f
C1247 VTAIL.n6 VSUBS 0.013948f
C1248 VTAIL.n7 VSUBS 0.024515f
C1249 VTAIL.n8 VSUBS 0.013174f
C1250 VTAIL.n9 VSUBS 0.031137f
C1251 VTAIL.n10 VSUBS 0.013561f
C1252 VTAIL.n11 VSUBS 0.024515f
C1253 VTAIL.n12 VSUBS 0.013948f
C1254 VTAIL.n13 VSUBS 0.031137f
C1255 VTAIL.n14 VSUBS 0.013948f
C1256 VTAIL.n15 VSUBS 0.024515f
C1257 VTAIL.n16 VSUBS 0.013174f
C1258 VTAIL.n17 VSUBS 0.031137f
C1259 VTAIL.n18 VSUBS 0.013948f
C1260 VTAIL.n19 VSUBS 0.024515f
C1261 VTAIL.n20 VSUBS 0.013174f
C1262 VTAIL.n21 VSUBS 0.031137f
C1263 VTAIL.n22 VSUBS 0.013948f
C1264 VTAIL.n23 VSUBS 0.024515f
C1265 VTAIL.n24 VSUBS 0.013174f
C1266 VTAIL.n25 VSUBS 0.031137f
C1267 VTAIL.n26 VSUBS 0.013948f
C1268 VTAIL.n27 VSUBS 0.024515f
C1269 VTAIL.n28 VSUBS 0.013174f
C1270 VTAIL.n29 VSUBS 0.031137f
C1271 VTAIL.n30 VSUBS 0.013948f
C1272 VTAIL.n31 VSUBS 1.85584f
C1273 VTAIL.n32 VSUBS 0.013174f
C1274 VTAIL.t15 VSUBS 0.066818f
C1275 VTAIL.n33 VSUBS 0.191685f
C1276 VTAIL.n34 VSUBS 0.019808f
C1277 VTAIL.n35 VSUBS 0.023353f
C1278 VTAIL.n36 VSUBS 0.031137f
C1279 VTAIL.n37 VSUBS 0.013948f
C1280 VTAIL.n38 VSUBS 0.013174f
C1281 VTAIL.n39 VSUBS 0.024515f
C1282 VTAIL.n40 VSUBS 0.024515f
C1283 VTAIL.n41 VSUBS 0.013174f
C1284 VTAIL.n42 VSUBS 0.013948f
C1285 VTAIL.n43 VSUBS 0.031137f
C1286 VTAIL.n44 VSUBS 0.031137f
C1287 VTAIL.n45 VSUBS 0.013948f
C1288 VTAIL.n46 VSUBS 0.013174f
C1289 VTAIL.n47 VSUBS 0.024515f
C1290 VTAIL.n48 VSUBS 0.024515f
C1291 VTAIL.n49 VSUBS 0.013174f
C1292 VTAIL.n50 VSUBS 0.013948f
C1293 VTAIL.n51 VSUBS 0.031137f
C1294 VTAIL.n52 VSUBS 0.031137f
C1295 VTAIL.n53 VSUBS 0.013948f
C1296 VTAIL.n54 VSUBS 0.013174f
C1297 VTAIL.n55 VSUBS 0.024515f
C1298 VTAIL.n56 VSUBS 0.024515f
C1299 VTAIL.n57 VSUBS 0.013174f
C1300 VTAIL.n58 VSUBS 0.013948f
C1301 VTAIL.n59 VSUBS 0.031137f
C1302 VTAIL.n60 VSUBS 0.031137f
C1303 VTAIL.n61 VSUBS 0.013948f
C1304 VTAIL.n62 VSUBS 0.013174f
C1305 VTAIL.n63 VSUBS 0.024515f
C1306 VTAIL.n64 VSUBS 0.024515f
C1307 VTAIL.n65 VSUBS 0.013174f
C1308 VTAIL.n66 VSUBS 0.013948f
C1309 VTAIL.n67 VSUBS 0.031137f
C1310 VTAIL.n68 VSUBS 0.031137f
C1311 VTAIL.n69 VSUBS 0.013948f
C1312 VTAIL.n70 VSUBS 0.013174f
C1313 VTAIL.n71 VSUBS 0.024515f
C1314 VTAIL.n72 VSUBS 0.024515f
C1315 VTAIL.n73 VSUBS 0.013174f
C1316 VTAIL.n74 VSUBS 0.013174f
C1317 VTAIL.n75 VSUBS 0.013948f
C1318 VTAIL.n76 VSUBS 0.031137f
C1319 VTAIL.n77 VSUBS 0.031137f
C1320 VTAIL.n78 VSUBS 0.031137f
C1321 VTAIL.n79 VSUBS 0.013561f
C1322 VTAIL.n80 VSUBS 0.013174f
C1323 VTAIL.n81 VSUBS 0.024515f
C1324 VTAIL.n82 VSUBS 0.024515f
C1325 VTAIL.n83 VSUBS 0.013174f
C1326 VTAIL.n84 VSUBS 0.013948f
C1327 VTAIL.n85 VSUBS 0.031137f
C1328 VTAIL.n86 VSUBS 0.031137f
C1329 VTAIL.n87 VSUBS 0.013948f
C1330 VTAIL.n88 VSUBS 0.013174f
C1331 VTAIL.n89 VSUBS 0.024515f
C1332 VTAIL.n90 VSUBS 0.024515f
C1333 VTAIL.n91 VSUBS 0.013174f
C1334 VTAIL.n92 VSUBS 0.013948f
C1335 VTAIL.n93 VSUBS 0.031137f
C1336 VTAIL.n94 VSUBS 0.076801f
C1337 VTAIL.n95 VSUBS 0.013948f
C1338 VTAIL.n96 VSUBS 0.013174f
C1339 VTAIL.n97 VSUBS 0.05968f
C1340 VTAIL.n98 VSUBS 0.038776f
C1341 VTAIL.n99 VSUBS 0.34713f
C1342 VTAIL.n100 VSUBS 0.027354f
C1343 VTAIL.n101 VSUBS 0.024515f
C1344 VTAIL.n102 VSUBS 0.013174f
C1345 VTAIL.n103 VSUBS 0.031137f
C1346 VTAIL.n104 VSUBS 0.013948f
C1347 VTAIL.n105 VSUBS 0.024515f
C1348 VTAIL.n106 VSUBS 0.013174f
C1349 VTAIL.n107 VSUBS 0.031137f
C1350 VTAIL.n108 VSUBS 0.013561f
C1351 VTAIL.n109 VSUBS 0.024515f
C1352 VTAIL.n110 VSUBS 0.013948f
C1353 VTAIL.n111 VSUBS 0.031137f
C1354 VTAIL.n112 VSUBS 0.013948f
C1355 VTAIL.n113 VSUBS 0.024515f
C1356 VTAIL.n114 VSUBS 0.013174f
C1357 VTAIL.n115 VSUBS 0.031137f
C1358 VTAIL.n116 VSUBS 0.013948f
C1359 VTAIL.n117 VSUBS 0.024515f
C1360 VTAIL.n118 VSUBS 0.013174f
C1361 VTAIL.n119 VSUBS 0.031137f
C1362 VTAIL.n120 VSUBS 0.013948f
C1363 VTAIL.n121 VSUBS 0.024515f
C1364 VTAIL.n122 VSUBS 0.013174f
C1365 VTAIL.n123 VSUBS 0.031137f
C1366 VTAIL.n124 VSUBS 0.013948f
C1367 VTAIL.n125 VSUBS 0.024515f
C1368 VTAIL.n126 VSUBS 0.013174f
C1369 VTAIL.n127 VSUBS 0.031137f
C1370 VTAIL.n128 VSUBS 0.013948f
C1371 VTAIL.n129 VSUBS 1.85584f
C1372 VTAIL.n130 VSUBS 0.013174f
C1373 VTAIL.t3 VSUBS 0.066818f
C1374 VTAIL.n131 VSUBS 0.191685f
C1375 VTAIL.n132 VSUBS 0.019808f
C1376 VTAIL.n133 VSUBS 0.023353f
C1377 VTAIL.n134 VSUBS 0.031137f
C1378 VTAIL.n135 VSUBS 0.013948f
C1379 VTAIL.n136 VSUBS 0.013174f
C1380 VTAIL.n137 VSUBS 0.024515f
C1381 VTAIL.n138 VSUBS 0.024515f
C1382 VTAIL.n139 VSUBS 0.013174f
C1383 VTAIL.n140 VSUBS 0.013948f
C1384 VTAIL.n141 VSUBS 0.031137f
C1385 VTAIL.n142 VSUBS 0.031137f
C1386 VTAIL.n143 VSUBS 0.013948f
C1387 VTAIL.n144 VSUBS 0.013174f
C1388 VTAIL.n145 VSUBS 0.024515f
C1389 VTAIL.n146 VSUBS 0.024515f
C1390 VTAIL.n147 VSUBS 0.013174f
C1391 VTAIL.n148 VSUBS 0.013948f
C1392 VTAIL.n149 VSUBS 0.031137f
C1393 VTAIL.n150 VSUBS 0.031137f
C1394 VTAIL.n151 VSUBS 0.013948f
C1395 VTAIL.n152 VSUBS 0.013174f
C1396 VTAIL.n153 VSUBS 0.024515f
C1397 VTAIL.n154 VSUBS 0.024515f
C1398 VTAIL.n155 VSUBS 0.013174f
C1399 VTAIL.n156 VSUBS 0.013948f
C1400 VTAIL.n157 VSUBS 0.031137f
C1401 VTAIL.n158 VSUBS 0.031137f
C1402 VTAIL.n159 VSUBS 0.013948f
C1403 VTAIL.n160 VSUBS 0.013174f
C1404 VTAIL.n161 VSUBS 0.024515f
C1405 VTAIL.n162 VSUBS 0.024515f
C1406 VTAIL.n163 VSUBS 0.013174f
C1407 VTAIL.n164 VSUBS 0.013948f
C1408 VTAIL.n165 VSUBS 0.031137f
C1409 VTAIL.n166 VSUBS 0.031137f
C1410 VTAIL.n167 VSUBS 0.013948f
C1411 VTAIL.n168 VSUBS 0.013174f
C1412 VTAIL.n169 VSUBS 0.024515f
C1413 VTAIL.n170 VSUBS 0.024515f
C1414 VTAIL.n171 VSUBS 0.013174f
C1415 VTAIL.n172 VSUBS 0.013174f
C1416 VTAIL.n173 VSUBS 0.013948f
C1417 VTAIL.n174 VSUBS 0.031137f
C1418 VTAIL.n175 VSUBS 0.031137f
C1419 VTAIL.n176 VSUBS 0.031137f
C1420 VTAIL.n177 VSUBS 0.013561f
C1421 VTAIL.n178 VSUBS 0.013174f
C1422 VTAIL.n179 VSUBS 0.024515f
C1423 VTAIL.n180 VSUBS 0.024515f
C1424 VTAIL.n181 VSUBS 0.013174f
C1425 VTAIL.n182 VSUBS 0.013948f
C1426 VTAIL.n183 VSUBS 0.031137f
C1427 VTAIL.n184 VSUBS 0.031137f
C1428 VTAIL.n185 VSUBS 0.013948f
C1429 VTAIL.n186 VSUBS 0.013174f
C1430 VTAIL.n187 VSUBS 0.024515f
C1431 VTAIL.n188 VSUBS 0.024515f
C1432 VTAIL.n189 VSUBS 0.013174f
C1433 VTAIL.n190 VSUBS 0.013948f
C1434 VTAIL.n191 VSUBS 0.031137f
C1435 VTAIL.n192 VSUBS 0.076801f
C1436 VTAIL.n193 VSUBS 0.013948f
C1437 VTAIL.n194 VSUBS 0.013174f
C1438 VTAIL.n195 VSUBS 0.05968f
C1439 VTAIL.n196 VSUBS 0.038776f
C1440 VTAIL.n197 VSUBS 0.34713f
C1441 VTAIL.t0 VSUBS 0.341156f
C1442 VTAIL.t6 VSUBS 0.341156f
C1443 VTAIL.n198 VSUBS 2.68824f
C1444 VTAIL.n199 VSUBS 1.16172f
C1445 VTAIL.n200 VSUBS 0.027354f
C1446 VTAIL.n201 VSUBS 0.024515f
C1447 VTAIL.n202 VSUBS 0.013174f
C1448 VTAIL.n203 VSUBS 0.031137f
C1449 VTAIL.n204 VSUBS 0.013948f
C1450 VTAIL.n205 VSUBS 0.024515f
C1451 VTAIL.n206 VSUBS 0.013174f
C1452 VTAIL.n207 VSUBS 0.031137f
C1453 VTAIL.n208 VSUBS 0.013561f
C1454 VTAIL.n209 VSUBS 0.024515f
C1455 VTAIL.n210 VSUBS 0.013948f
C1456 VTAIL.n211 VSUBS 0.031137f
C1457 VTAIL.n212 VSUBS 0.013948f
C1458 VTAIL.n213 VSUBS 0.024515f
C1459 VTAIL.n214 VSUBS 0.013174f
C1460 VTAIL.n215 VSUBS 0.031137f
C1461 VTAIL.n216 VSUBS 0.013948f
C1462 VTAIL.n217 VSUBS 0.024515f
C1463 VTAIL.n218 VSUBS 0.013174f
C1464 VTAIL.n219 VSUBS 0.031137f
C1465 VTAIL.n220 VSUBS 0.013948f
C1466 VTAIL.n221 VSUBS 0.024515f
C1467 VTAIL.n222 VSUBS 0.013174f
C1468 VTAIL.n223 VSUBS 0.031137f
C1469 VTAIL.n224 VSUBS 0.013948f
C1470 VTAIL.n225 VSUBS 0.024515f
C1471 VTAIL.n226 VSUBS 0.013174f
C1472 VTAIL.n227 VSUBS 0.031137f
C1473 VTAIL.n228 VSUBS 0.013948f
C1474 VTAIL.n229 VSUBS 1.85584f
C1475 VTAIL.n230 VSUBS 0.013174f
C1476 VTAIL.t7 VSUBS 0.066818f
C1477 VTAIL.n231 VSUBS 0.191685f
C1478 VTAIL.n232 VSUBS 0.019808f
C1479 VTAIL.n233 VSUBS 0.023353f
C1480 VTAIL.n234 VSUBS 0.031137f
C1481 VTAIL.n235 VSUBS 0.013948f
C1482 VTAIL.n236 VSUBS 0.013174f
C1483 VTAIL.n237 VSUBS 0.024515f
C1484 VTAIL.n238 VSUBS 0.024515f
C1485 VTAIL.n239 VSUBS 0.013174f
C1486 VTAIL.n240 VSUBS 0.013948f
C1487 VTAIL.n241 VSUBS 0.031137f
C1488 VTAIL.n242 VSUBS 0.031137f
C1489 VTAIL.n243 VSUBS 0.013948f
C1490 VTAIL.n244 VSUBS 0.013174f
C1491 VTAIL.n245 VSUBS 0.024515f
C1492 VTAIL.n246 VSUBS 0.024515f
C1493 VTAIL.n247 VSUBS 0.013174f
C1494 VTAIL.n248 VSUBS 0.013948f
C1495 VTAIL.n249 VSUBS 0.031137f
C1496 VTAIL.n250 VSUBS 0.031137f
C1497 VTAIL.n251 VSUBS 0.013948f
C1498 VTAIL.n252 VSUBS 0.013174f
C1499 VTAIL.n253 VSUBS 0.024515f
C1500 VTAIL.n254 VSUBS 0.024515f
C1501 VTAIL.n255 VSUBS 0.013174f
C1502 VTAIL.n256 VSUBS 0.013948f
C1503 VTAIL.n257 VSUBS 0.031137f
C1504 VTAIL.n258 VSUBS 0.031137f
C1505 VTAIL.n259 VSUBS 0.013948f
C1506 VTAIL.n260 VSUBS 0.013174f
C1507 VTAIL.n261 VSUBS 0.024515f
C1508 VTAIL.n262 VSUBS 0.024515f
C1509 VTAIL.n263 VSUBS 0.013174f
C1510 VTAIL.n264 VSUBS 0.013948f
C1511 VTAIL.n265 VSUBS 0.031137f
C1512 VTAIL.n266 VSUBS 0.031137f
C1513 VTAIL.n267 VSUBS 0.013948f
C1514 VTAIL.n268 VSUBS 0.013174f
C1515 VTAIL.n269 VSUBS 0.024515f
C1516 VTAIL.n270 VSUBS 0.024515f
C1517 VTAIL.n271 VSUBS 0.013174f
C1518 VTAIL.n272 VSUBS 0.013174f
C1519 VTAIL.n273 VSUBS 0.013948f
C1520 VTAIL.n274 VSUBS 0.031137f
C1521 VTAIL.n275 VSUBS 0.031137f
C1522 VTAIL.n276 VSUBS 0.031137f
C1523 VTAIL.n277 VSUBS 0.013561f
C1524 VTAIL.n278 VSUBS 0.013174f
C1525 VTAIL.n279 VSUBS 0.024515f
C1526 VTAIL.n280 VSUBS 0.024515f
C1527 VTAIL.n281 VSUBS 0.013174f
C1528 VTAIL.n282 VSUBS 0.013948f
C1529 VTAIL.n283 VSUBS 0.031137f
C1530 VTAIL.n284 VSUBS 0.031137f
C1531 VTAIL.n285 VSUBS 0.013948f
C1532 VTAIL.n286 VSUBS 0.013174f
C1533 VTAIL.n287 VSUBS 0.024515f
C1534 VTAIL.n288 VSUBS 0.024515f
C1535 VTAIL.n289 VSUBS 0.013174f
C1536 VTAIL.n290 VSUBS 0.013948f
C1537 VTAIL.n291 VSUBS 0.031137f
C1538 VTAIL.n292 VSUBS 0.076801f
C1539 VTAIL.n293 VSUBS 0.013948f
C1540 VTAIL.n294 VSUBS 0.013174f
C1541 VTAIL.n295 VSUBS 0.05968f
C1542 VTAIL.n296 VSUBS 0.038776f
C1543 VTAIL.n297 VSUBS 2.12962f
C1544 VTAIL.n298 VSUBS 0.027354f
C1545 VTAIL.n299 VSUBS 0.024515f
C1546 VTAIL.n300 VSUBS 0.013174f
C1547 VTAIL.n301 VSUBS 0.031137f
C1548 VTAIL.n302 VSUBS 0.013948f
C1549 VTAIL.n303 VSUBS 0.024515f
C1550 VTAIL.n304 VSUBS 0.013174f
C1551 VTAIL.n305 VSUBS 0.031137f
C1552 VTAIL.n306 VSUBS 0.013561f
C1553 VTAIL.n307 VSUBS 0.024515f
C1554 VTAIL.n308 VSUBS 0.013561f
C1555 VTAIL.n309 VSUBS 0.013174f
C1556 VTAIL.n310 VSUBS 0.031137f
C1557 VTAIL.n311 VSUBS 0.031137f
C1558 VTAIL.n312 VSUBS 0.013948f
C1559 VTAIL.n313 VSUBS 0.024515f
C1560 VTAIL.n314 VSUBS 0.013174f
C1561 VTAIL.n315 VSUBS 0.031137f
C1562 VTAIL.n316 VSUBS 0.013948f
C1563 VTAIL.n317 VSUBS 0.024515f
C1564 VTAIL.n318 VSUBS 0.013174f
C1565 VTAIL.n319 VSUBS 0.031137f
C1566 VTAIL.n320 VSUBS 0.013948f
C1567 VTAIL.n321 VSUBS 0.024515f
C1568 VTAIL.n322 VSUBS 0.013174f
C1569 VTAIL.n323 VSUBS 0.031137f
C1570 VTAIL.n324 VSUBS 0.013948f
C1571 VTAIL.n325 VSUBS 0.024515f
C1572 VTAIL.n326 VSUBS 0.013174f
C1573 VTAIL.n327 VSUBS 0.031137f
C1574 VTAIL.n328 VSUBS 0.013948f
C1575 VTAIL.n329 VSUBS 1.85584f
C1576 VTAIL.n330 VSUBS 0.013174f
C1577 VTAIL.t12 VSUBS 0.066818f
C1578 VTAIL.n331 VSUBS 0.191685f
C1579 VTAIL.n332 VSUBS 0.019808f
C1580 VTAIL.n333 VSUBS 0.023353f
C1581 VTAIL.n334 VSUBS 0.031137f
C1582 VTAIL.n335 VSUBS 0.013948f
C1583 VTAIL.n336 VSUBS 0.013174f
C1584 VTAIL.n337 VSUBS 0.024515f
C1585 VTAIL.n338 VSUBS 0.024515f
C1586 VTAIL.n339 VSUBS 0.013174f
C1587 VTAIL.n340 VSUBS 0.013948f
C1588 VTAIL.n341 VSUBS 0.031137f
C1589 VTAIL.n342 VSUBS 0.031137f
C1590 VTAIL.n343 VSUBS 0.013948f
C1591 VTAIL.n344 VSUBS 0.013174f
C1592 VTAIL.n345 VSUBS 0.024515f
C1593 VTAIL.n346 VSUBS 0.024515f
C1594 VTAIL.n347 VSUBS 0.013174f
C1595 VTAIL.n348 VSUBS 0.013948f
C1596 VTAIL.n349 VSUBS 0.031137f
C1597 VTAIL.n350 VSUBS 0.031137f
C1598 VTAIL.n351 VSUBS 0.013948f
C1599 VTAIL.n352 VSUBS 0.013174f
C1600 VTAIL.n353 VSUBS 0.024515f
C1601 VTAIL.n354 VSUBS 0.024515f
C1602 VTAIL.n355 VSUBS 0.013174f
C1603 VTAIL.n356 VSUBS 0.013948f
C1604 VTAIL.n357 VSUBS 0.031137f
C1605 VTAIL.n358 VSUBS 0.031137f
C1606 VTAIL.n359 VSUBS 0.013948f
C1607 VTAIL.n360 VSUBS 0.013174f
C1608 VTAIL.n361 VSUBS 0.024515f
C1609 VTAIL.n362 VSUBS 0.024515f
C1610 VTAIL.n363 VSUBS 0.013174f
C1611 VTAIL.n364 VSUBS 0.013948f
C1612 VTAIL.n365 VSUBS 0.031137f
C1613 VTAIL.n366 VSUBS 0.031137f
C1614 VTAIL.n367 VSUBS 0.013948f
C1615 VTAIL.n368 VSUBS 0.013174f
C1616 VTAIL.n369 VSUBS 0.024515f
C1617 VTAIL.n370 VSUBS 0.024515f
C1618 VTAIL.n371 VSUBS 0.013174f
C1619 VTAIL.n372 VSUBS 0.013948f
C1620 VTAIL.n373 VSUBS 0.031137f
C1621 VTAIL.n374 VSUBS 0.031137f
C1622 VTAIL.n375 VSUBS 0.013948f
C1623 VTAIL.n376 VSUBS 0.013174f
C1624 VTAIL.n377 VSUBS 0.024515f
C1625 VTAIL.n378 VSUBS 0.024515f
C1626 VTAIL.n379 VSUBS 0.013174f
C1627 VTAIL.n380 VSUBS 0.013948f
C1628 VTAIL.n381 VSUBS 0.031137f
C1629 VTAIL.n382 VSUBS 0.031137f
C1630 VTAIL.n383 VSUBS 0.013948f
C1631 VTAIL.n384 VSUBS 0.013174f
C1632 VTAIL.n385 VSUBS 0.024515f
C1633 VTAIL.n386 VSUBS 0.024515f
C1634 VTAIL.n387 VSUBS 0.013174f
C1635 VTAIL.n388 VSUBS 0.013948f
C1636 VTAIL.n389 VSUBS 0.031137f
C1637 VTAIL.n390 VSUBS 0.076801f
C1638 VTAIL.n391 VSUBS 0.013948f
C1639 VTAIL.n392 VSUBS 0.013174f
C1640 VTAIL.n393 VSUBS 0.05968f
C1641 VTAIL.n394 VSUBS 0.038776f
C1642 VTAIL.n395 VSUBS 2.12962f
C1643 VTAIL.t13 VSUBS 0.341156f
C1644 VTAIL.t10 VSUBS 0.341156f
C1645 VTAIL.n396 VSUBS 2.68825f
C1646 VTAIL.n397 VSUBS 1.16171f
C1647 VTAIL.n398 VSUBS 0.027354f
C1648 VTAIL.n399 VSUBS 0.024515f
C1649 VTAIL.n400 VSUBS 0.013174f
C1650 VTAIL.n401 VSUBS 0.031137f
C1651 VTAIL.n402 VSUBS 0.013948f
C1652 VTAIL.n403 VSUBS 0.024515f
C1653 VTAIL.n404 VSUBS 0.013174f
C1654 VTAIL.n405 VSUBS 0.031137f
C1655 VTAIL.n406 VSUBS 0.013561f
C1656 VTAIL.n407 VSUBS 0.024515f
C1657 VTAIL.n408 VSUBS 0.013561f
C1658 VTAIL.n409 VSUBS 0.013174f
C1659 VTAIL.n410 VSUBS 0.031137f
C1660 VTAIL.n411 VSUBS 0.031137f
C1661 VTAIL.n412 VSUBS 0.013948f
C1662 VTAIL.n413 VSUBS 0.024515f
C1663 VTAIL.n414 VSUBS 0.013174f
C1664 VTAIL.n415 VSUBS 0.031137f
C1665 VTAIL.n416 VSUBS 0.013948f
C1666 VTAIL.n417 VSUBS 0.024515f
C1667 VTAIL.n418 VSUBS 0.013174f
C1668 VTAIL.n419 VSUBS 0.031137f
C1669 VTAIL.n420 VSUBS 0.013948f
C1670 VTAIL.n421 VSUBS 0.024515f
C1671 VTAIL.n422 VSUBS 0.013174f
C1672 VTAIL.n423 VSUBS 0.031137f
C1673 VTAIL.n424 VSUBS 0.013948f
C1674 VTAIL.n425 VSUBS 0.024515f
C1675 VTAIL.n426 VSUBS 0.013174f
C1676 VTAIL.n427 VSUBS 0.031137f
C1677 VTAIL.n428 VSUBS 0.013948f
C1678 VTAIL.n429 VSUBS 1.85584f
C1679 VTAIL.n430 VSUBS 0.013174f
C1680 VTAIL.t11 VSUBS 0.066818f
C1681 VTAIL.n431 VSUBS 0.191685f
C1682 VTAIL.n432 VSUBS 0.019808f
C1683 VTAIL.n433 VSUBS 0.023353f
C1684 VTAIL.n434 VSUBS 0.031137f
C1685 VTAIL.n435 VSUBS 0.013948f
C1686 VTAIL.n436 VSUBS 0.013174f
C1687 VTAIL.n437 VSUBS 0.024515f
C1688 VTAIL.n438 VSUBS 0.024515f
C1689 VTAIL.n439 VSUBS 0.013174f
C1690 VTAIL.n440 VSUBS 0.013948f
C1691 VTAIL.n441 VSUBS 0.031137f
C1692 VTAIL.n442 VSUBS 0.031137f
C1693 VTAIL.n443 VSUBS 0.013948f
C1694 VTAIL.n444 VSUBS 0.013174f
C1695 VTAIL.n445 VSUBS 0.024515f
C1696 VTAIL.n446 VSUBS 0.024515f
C1697 VTAIL.n447 VSUBS 0.013174f
C1698 VTAIL.n448 VSUBS 0.013948f
C1699 VTAIL.n449 VSUBS 0.031137f
C1700 VTAIL.n450 VSUBS 0.031137f
C1701 VTAIL.n451 VSUBS 0.013948f
C1702 VTAIL.n452 VSUBS 0.013174f
C1703 VTAIL.n453 VSUBS 0.024515f
C1704 VTAIL.n454 VSUBS 0.024515f
C1705 VTAIL.n455 VSUBS 0.013174f
C1706 VTAIL.n456 VSUBS 0.013948f
C1707 VTAIL.n457 VSUBS 0.031137f
C1708 VTAIL.n458 VSUBS 0.031137f
C1709 VTAIL.n459 VSUBS 0.013948f
C1710 VTAIL.n460 VSUBS 0.013174f
C1711 VTAIL.n461 VSUBS 0.024515f
C1712 VTAIL.n462 VSUBS 0.024515f
C1713 VTAIL.n463 VSUBS 0.013174f
C1714 VTAIL.n464 VSUBS 0.013948f
C1715 VTAIL.n465 VSUBS 0.031137f
C1716 VTAIL.n466 VSUBS 0.031137f
C1717 VTAIL.n467 VSUBS 0.013948f
C1718 VTAIL.n468 VSUBS 0.013174f
C1719 VTAIL.n469 VSUBS 0.024515f
C1720 VTAIL.n470 VSUBS 0.024515f
C1721 VTAIL.n471 VSUBS 0.013174f
C1722 VTAIL.n472 VSUBS 0.013948f
C1723 VTAIL.n473 VSUBS 0.031137f
C1724 VTAIL.n474 VSUBS 0.031137f
C1725 VTAIL.n475 VSUBS 0.013948f
C1726 VTAIL.n476 VSUBS 0.013174f
C1727 VTAIL.n477 VSUBS 0.024515f
C1728 VTAIL.n478 VSUBS 0.024515f
C1729 VTAIL.n479 VSUBS 0.013174f
C1730 VTAIL.n480 VSUBS 0.013948f
C1731 VTAIL.n481 VSUBS 0.031137f
C1732 VTAIL.n482 VSUBS 0.031137f
C1733 VTAIL.n483 VSUBS 0.013948f
C1734 VTAIL.n484 VSUBS 0.013174f
C1735 VTAIL.n485 VSUBS 0.024515f
C1736 VTAIL.n486 VSUBS 0.024515f
C1737 VTAIL.n487 VSUBS 0.013174f
C1738 VTAIL.n488 VSUBS 0.013948f
C1739 VTAIL.n489 VSUBS 0.031137f
C1740 VTAIL.n490 VSUBS 0.076801f
C1741 VTAIL.n491 VSUBS 0.013948f
C1742 VTAIL.n492 VSUBS 0.013174f
C1743 VTAIL.n493 VSUBS 0.05968f
C1744 VTAIL.n494 VSUBS 0.038776f
C1745 VTAIL.n495 VSUBS 0.34713f
C1746 VTAIL.n496 VSUBS 0.027354f
C1747 VTAIL.n497 VSUBS 0.024515f
C1748 VTAIL.n498 VSUBS 0.013174f
C1749 VTAIL.n499 VSUBS 0.031137f
C1750 VTAIL.n500 VSUBS 0.013948f
C1751 VTAIL.n501 VSUBS 0.024515f
C1752 VTAIL.n502 VSUBS 0.013174f
C1753 VTAIL.n503 VSUBS 0.031137f
C1754 VTAIL.n504 VSUBS 0.013561f
C1755 VTAIL.n505 VSUBS 0.024515f
C1756 VTAIL.n506 VSUBS 0.013561f
C1757 VTAIL.n507 VSUBS 0.013174f
C1758 VTAIL.n508 VSUBS 0.031137f
C1759 VTAIL.n509 VSUBS 0.031137f
C1760 VTAIL.n510 VSUBS 0.013948f
C1761 VTAIL.n511 VSUBS 0.024515f
C1762 VTAIL.n512 VSUBS 0.013174f
C1763 VTAIL.n513 VSUBS 0.031137f
C1764 VTAIL.n514 VSUBS 0.013948f
C1765 VTAIL.n515 VSUBS 0.024515f
C1766 VTAIL.n516 VSUBS 0.013174f
C1767 VTAIL.n517 VSUBS 0.031137f
C1768 VTAIL.n518 VSUBS 0.013948f
C1769 VTAIL.n519 VSUBS 0.024515f
C1770 VTAIL.n520 VSUBS 0.013174f
C1771 VTAIL.n521 VSUBS 0.031137f
C1772 VTAIL.n522 VSUBS 0.013948f
C1773 VTAIL.n523 VSUBS 0.024515f
C1774 VTAIL.n524 VSUBS 0.013174f
C1775 VTAIL.n525 VSUBS 0.031137f
C1776 VTAIL.n526 VSUBS 0.013948f
C1777 VTAIL.n527 VSUBS 1.85584f
C1778 VTAIL.n528 VSUBS 0.013174f
C1779 VTAIL.t5 VSUBS 0.066818f
C1780 VTAIL.n529 VSUBS 0.191685f
C1781 VTAIL.n530 VSUBS 0.019808f
C1782 VTAIL.n531 VSUBS 0.023353f
C1783 VTAIL.n532 VSUBS 0.031137f
C1784 VTAIL.n533 VSUBS 0.013948f
C1785 VTAIL.n534 VSUBS 0.013174f
C1786 VTAIL.n535 VSUBS 0.024515f
C1787 VTAIL.n536 VSUBS 0.024515f
C1788 VTAIL.n537 VSUBS 0.013174f
C1789 VTAIL.n538 VSUBS 0.013948f
C1790 VTAIL.n539 VSUBS 0.031137f
C1791 VTAIL.n540 VSUBS 0.031137f
C1792 VTAIL.n541 VSUBS 0.013948f
C1793 VTAIL.n542 VSUBS 0.013174f
C1794 VTAIL.n543 VSUBS 0.024515f
C1795 VTAIL.n544 VSUBS 0.024515f
C1796 VTAIL.n545 VSUBS 0.013174f
C1797 VTAIL.n546 VSUBS 0.013948f
C1798 VTAIL.n547 VSUBS 0.031137f
C1799 VTAIL.n548 VSUBS 0.031137f
C1800 VTAIL.n549 VSUBS 0.013948f
C1801 VTAIL.n550 VSUBS 0.013174f
C1802 VTAIL.n551 VSUBS 0.024515f
C1803 VTAIL.n552 VSUBS 0.024515f
C1804 VTAIL.n553 VSUBS 0.013174f
C1805 VTAIL.n554 VSUBS 0.013948f
C1806 VTAIL.n555 VSUBS 0.031137f
C1807 VTAIL.n556 VSUBS 0.031137f
C1808 VTAIL.n557 VSUBS 0.013948f
C1809 VTAIL.n558 VSUBS 0.013174f
C1810 VTAIL.n559 VSUBS 0.024515f
C1811 VTAIL.n560 VSUBS 0.024515f
C1812 VTAIL.n561 VSUBS 0.013174f
C1813 VTAIL.n562 VSUBS 0.013948f
C1814 VTAIL.n563 VSUBS 0.031137f
C1815 VTAIL.n564 VSUBS 0.031137f
C1816 VTAIL.n565 VSUBS 0.013948f
C1817 VTAIL.n566 VSUBS 0.013174f
C1818 VTAIL.n567 VSUBS 0.024515f
C1819 VTAIL.n568 VSUBS 0.024515f
C1820 VTAIL.n569 VSUBS 0.013174f
C1821 VTAIL.n570 VSUBS 0.013948f
C1822 VTAIL.n571 VSUBS 0.031137f
C1823 VTAIL.n572 VSUBS 0.031137f
C1824 VTAIL.n573 VSUBS 0.013948f
C1825 VTAIL.n574 VSUBS 0.013174f
C1826 VTAIL.n575 VSUBS 0.024515f
C1827 VTAIL.n576 VSUBS 0.024515f
C1828 VTAIL.n577 VSUBS 0.013174f
C1829 VTAIL.n578 VSUBS 0.013948f
C1830 VTAIL.n579 VSUBS 0.031137f
C1831 VTAIL.n580 VSUBS 0.031137f
C1832 VTAIL.n581 VSUBS 0.013948f
C1833 VTAIL.n582 VSUBS 0.013174f
C1834 VTAIL.n583 VSUBS 0.024515f
C1835 VTAIL.n584 VSUBS 0.024515f
C1836 VTAIL.n585 VSUBS 0.013174f
C1837 VTAIL.n586 VSUBS 0.013948f
C1838 VTAIL.n587 VSUBS 0.031137f
C1839 VTAIL.n588 VSUBS 0.076801f
C1840 VTAIL.n589 VSUBS 0.013948f
C1841 VTAIL.n590 VSUBS 0.013174f
C1842 VTAIL.n591 VSUBS 0.05968f
C1843 VTAIL.n592 VSUBS 0.038776f
C1844 VTAIL.n593 VSUBS 0.34713f
C1845 VTAIL.t1 VSUBS 0.341156f
C1846 VTAIL.t4 VSUBS 0.341156f
C1847 VTAIL.n594 VSUBS 2.68825f
C1848 VTAIL.n595 VSUBS 1.16171f
C1849 VTAIL.n596 VSUBS 0.027354f
C1850 VTAIL.n597 VSUBS 0.024515f
C1851 VTAIL.n598 VSUBS 0.013174f
C1852 VTAIL.n599 VSUBS 0.031137f
C1853 VTAIL.n600 VSUBS 0.013948f
C1854 VTAIL.n601 VSUBS 0.024515f
C1855 VTAIL.n602 VSUBS 0.013174f
C1856 VTAIL.n603 VSUBS 0.031137f
C1857 VTAIL.n604 VSUBS 0.013561f
C1858 VTAIL.n605 VSUBS 0.024515f
C1859 VTAIL.n606 VSUBS 0.013561f
C1860 VTAIL.n607 VSUBS 0.013174f
C1861 VTAIL.n608 VSUBS 0.031137f
C1862 VTAIL.n609 VSUBS 0.031137f
C1863 VTAIL.n610 VSUBS 0.013948f
C1864 VTAIL.n611 VSUBS 0.024515f
C1865 VTAIL.n612 VSUBS 0.013174f
C1866 VTAIL.n613 VSUBS 0.031137f
C1867 VTAIL.n614 VSUBS 0.013948f
C1868 VTAIL.n615 VSUBS 0.024515f
C1869 VTAIL.n616 VSUBS 0.013174f
C1870 VTAIL.n617 VSUBS 0.031137f
C1871 VTAIL.n618 VSUBS 0.013948f
C1872 VTAIL.n619 VSUBS 0.024515f
C1873 VTAIL.n620 VSUBS 0.013174f
C1874 VTAIL.n621 VSUBS 0.031137f
C1875 VTAIL.n622 VSUBS 0.013948f
C1876 VTAIL.n623 VSUBS 0.024515f
C1877 VTAIL.n624 VSUBS 0.013174f
C1878 VTAIL.n625 VSUBS 0.031137f
C1879 VTAIL.n626 VSUBS 0.013948f
C1880 VTAIL.n627 VSUBS 1.85584f
C1881 VTAIL.n628 VSUBS 0.013174f
C1882 VTAIL.t2 VSUBS 0.066818f
C1883 VTAIL.n629 VSUBS 0.191685f
C1884 VTAIL.n630 VSUBS 0.019808f
C1885 VTAIL.n631 VSUBS 0.023353f
C1886 VTAIL.n632 VSUBS 0.031137f
C1887 VTAIL.n633 VSUBS 0.013948f
C1888 VTAIL.n634 VSUBS 0.013174f
C1889 VTAIL.n635 VSUBS 0.024515f
C1890 VTAIL.n636 VSUBS 0.024515f
C1891 VTAIL.n637 VSUBS 0.013174f
C1892 VTAIL.n638 VSUBS 0.013948f
C1893 VTAIL.n639 VSUBS 0.031137f
C1894 VTAIL.n640 VSUBS 0.031137f
C1895 VTAIL.n641 VSUBS 0.013948f
C1896 VTAIL.n642 VSUBS 0.013174f
C1897 VTAIL.n643 VSUBS 0.024515f
C1898 VTAIL.n644 VSUBS 0.024515f
C1899 VTAIL.n645 VSUBS 0.013174f
C1900 VTAIL.n646 VSUBS 0.013948f
C1901 VTAIL.n647 VSUBS 0.031137f
C1902 VTAIL.n648 VSUBS 0.031137f
C1903 VTAIL.n649 VSUBS 0.013948f
C1904 VTAIL.n650 VSUBS 0.013174f
C1905 VTAIL.n651 VSUBS 0.024515f
C1906 VTAIL.n652 VSUBS 0.024515f
C1907 VTAIL.n653 VSUBS 0.013174f
C1908 VTAIL.n654 VSUBS 0.013948f
C1909 VTAIL.n655 VSUBS 0.031137f
C1910 VTAIL.n656 VSUBS 0.031137f
C1911 VTAIL.n657 VSUBS 0.013948f
C1912 VTAIL.n658 VSUBS 0.013174f
C1913 VTAIL.n659 VSUBS 0.024515f
C1914 VTAIL.n660 VSUBS 0.024515f
C1915 VTAIL.n661 VSUBS 0.013174f
C1916 VTAIL.n662 VSUBS 0.013948f
C1917 VTAIL.n663 VSUBS 0.031137f
C1918 VTAIL.n664 VSUBS 0.031137f
C1919 VTAIL.n665 VSUBS 0.013948f
C1920 VTAIL.n666 VSUBS 0.013174f
C1921 VTAIL.n667 VSUBS 0.024515f
C1922 VTAIL.n668 VSUBS 0.024515f
C1923 VTAIL.n669 VSUBS 0.013174f
C1924 VTAIL.n670 VSUBS 0.013948f
C1925 VTAIL.n671 VSUBS 0.031137f
C1926 VTAIL.n672 VSUBS 0.031137f
C1927 VTAIL.n673 VSUBS 0.013948f
C1928 VTAIL.n674 VSUBS 0.013174f
C1929 VTAIL.n675 VSUBS 0.024515f
C1930 VTAIL.n676 VSUBS 0.024515f
C1931 VTAIL.n677 VSUBS 0.013174f
C1932 VTAIL.n678 VSUBS 0.013948f
C1933 VTAIL.n679 VSUBS 0.031137f
C1934 VTAIL.n680 VSUBS 0.031137f
C1935 VTAIL.n681 VSUBS 0.013948f
C1936 VTAIL.n682 VSUBS 0.013174f
C1937 VTAIL.n683 VSUBS 0.024515f
C1938 VTAIL.n684 VSUBS 0.024515f
C1939 VTAIL.n685 VSUBS 0.013174f
C1940 VTAIL.n686 VSUBS 0.013948f
C1941 VTAIL.n687 VSUBS 0.031137f
C1942 VTAIL.n688 VSUBS 0.076801f
C1943 VTAIL.n689 VSUBS 0.013948f
C1944 VTAIL.n690 VSUBS 0.013174f
C1945 VTAIL.n691 VSUBS 0.05968f
C1946 VTAIL.n692 VSUBS 0.038776f
C1947 VTAIL.n693 VSUBS 2.12962f
C1948 VTAIL.n694 VSUBS 0.027354f
C1949 VTAIL.n695 VSUBS 0.024515f
C1950 VTAIL.n696 VSUBS 0.013174f
C1951 VTAIL.n697 VSUBS 0.031137f
C1952 VTAIL.n698 VSUBS 0.013948f
C1953 VTAIL.n699 VSUBS 0.024515f
C1954 VTAIL.n700 VSUBS 0.013174f
C1955 VTAIL.n701 VSUBS 0.031137f
C1956 VTAIL.n702 VSUBS 0.013561f
C1957 VTAIL.n703 VSUBS 0.024515f
C1958 VTAIL.n704 VSUBS 0.013948f
C1959 VTAIL.n705 VSUBS 0.031137f
C1960 VTAIL.n706 VSUBS 0.013948f
C1961 VTAIL.n707 VSUBS 0.024515f
C1962 VTAIL.n708 VSUBS 0.013174f
C1963 VTAIL.n709 VSUBS 0.031137f
C1964 VTAIL.n710 VSUBS 0.013948f
C1965 VTAIL.n711 VSUBS 0.024515f
C1966 VTAIL.n712 VSUBS 0.013174f
C1967 VTAIL.n713 VSUBS 0.031137f
C1968 VTAIL.n714 VSUBS 0.013948f
C1969 VTAIL.n715 VSUBS 0.024515f
C1970 VTAIL.n716 VSUBS 0.013174f
C1971 VTAIL.n717 VSUBS 0.031137f
C1972 VTAIL.n718 VSUBS 0.013948f
C1973 VTAIL.n719 VSUBS 0.024515f
C1974 VTAIL.n720 VSUBS 0.013174f
C1975 VTAIL.n721 VSUBS 0.031137f
C1976 VTAIL.n722 VSUBS 0.013948f
C1977 VTAIL.n723 VSUBS 1.85584f
C1978 VTAIL.n724 VSUBS 0.013174f
C1979 VTAIL.t8 VSUBS 0.066818f
C1980 VTAIL.n725 VSUBS 0.191685f
C1981 VTAIL.n726 VSUBS 0.019808f
C1982 VTAIL.n727 VSUBS 0.023353f
C1983 VTAIL.n728 VSUBS 0.031137f
C1984 VTAIL.n729 VSUBS 0.013948f
C1985 VTAIL.n730 VSUBS 0.013174f
C1986 VTAIL.n731 VSUBS 0.024515f
C1987 VTAIL.n732 VSUBS 0.024515f
C1988 VTAIL.n733 VSUBS 0.013174f
C1989 VTAIL.n734 VSUBS 0.013948f
C1990 VTAIL.n735 VSUBS 0.031137f
C1991 VTAIL.n736 VSUBS 0.031137f
C1992 VTAIL.n737 VSUBS 0.013948f
C1993 VTAIL.n738 VSUBS 0.013174f
C1994 VTAIL.n739 VSUBS 0.024515f
C1995 VTAIL.n740 VSUBS 0.024515f
C1996 VTAIL.n741 VSUBS 0.013174f
C1997 VTAIL.n742 VSUBS 0.013948f
C1998 VTAIL.n743 VSUBS 0.031137f
C1999 VTAIL.n744 VSUBS 0.031137f
C2000 VTAIL.n745 VSUBS 0.013948f
C2001 VTAIL.n746 VSUBS 0.013174f
C2002 VTAIL.n747 VSUBS 0.024515f
C2003 VTAIL.n748 VSUBS 0.024515f
C2004 VTAIL.n749 VSUBS 0.013174f
C2005 VTAIL.n750 VSUBS 0.013948f
C2006 VTAIL.n751 VSUBS 0.031137f
C2007 VTAIL.n752 VSUBS 0.031137f
C2008 VTAIL.n753 VSUBS 0.013948f
C2009 VTAIL.n754 VSUBS 0.013174f
C2010 VTAIL.n755 VSUBS 0.024515f
C2011 VTAIL.n756 VSUBS 0.024515f
C2012 VTAIL.n757 VSUBS 0.013174f
C2013 VTAIL.n758 VSUBS 0.013948f
C2014 VTAIL.n759 VSUBS 0.031137f
C2015 VTAIL.n760 VSUBS 0.031137f
C2016 VTAIL.n761 VSUBS 0.013948f
C2017 VTAIL.n762 VSUBS 0.013174f
C2018 VTAIL.n763 VSUBS 0.024515f
C2019 VTAIL.n764 VSUBS 0.024515f
C2020 VTAIL.n765 VSUBS 0.013174f
C2021 VTAIL.n766 VSUBS 0.013174f
C2022 VTAIL.n767 VSUBS 0.013948f
C2023 VTAIL.n768 VSUBS 0.031137f
C2024 VTAIL.n769 VSUBS 0.031137f
C2025 VTAIL.n770 VSUBS 0.031137f
C2026 VTAIL.n771 VSUBS 0.013561f
C2027 VTAIL.n772 VSUBS 0.013174f
C2028 VTAIL.n773 VSUBS 0.024515f
C2029 VTAIL.n774 VSUBS 0.024515f
C2030 VTAIL.n775 VSUBS 0.013174f
C2031 VTAIL.n776 VSUBS 0.013948f
C2032 VTAIL.n777 VSUBS 0.031137f
C2033 VTAIL.n778 VSUBS 0.031137f
C2034 VTAIL.n779 VSUBS 0.013948f
C2035 VTAIL.n780 VSUBS 0.013174f
C2036 VTAIL.n781 VSUBS 0.024515f
C2037 VTAIL.n782 VSUBS 0.024515f
C2038 VTAIL.n783 VSUBS 0.013174f
C2039 VTAIL.n784 VSUBS 0.013948f
C2040 VTAIL.n785 VSUBS 0.031137f
C2041 VTAIL.n786 VSUBS 0.076801f
C2042 VTAIL.n787 VSUBS 0.013948f
C2043 VTAIL.n788 VSUBS 0.013174f
C2044 VTAIL.n789 VSUBS 0.05968f
C2045 VTAIL.n790 VSUBS 0.038776f
C2046 VTAIL.n791 VSUBS 2.12502f
C2047 VDD2.t3 VSUBS 0.439188f
C2048 VDD2.t7 VSUBS 0.439188f
C2049 VDD2.n0 VSUBS 3.67605f
C2050 VDD2.t2 VSUBS 0.439188f
C2051 VDD2.t6 VSUBS 0.439188f
C2052 VDD2.n1 VSUBS 3.67605f
C2053 VDD2.n2 VSUBS 6.2223f
C2054 VDD2.t0 VSUBS 0.439188f
C2055 VDD2.t1 VSUBS 0.439188f
C2056 VDD2.n3 VSUBS 3.64751f
C2057 VDD2.n4 VSUBS 5.17366f
C2058 VDD2.t4 VSUBS 0.439188f
C2059 VDD2.t5 VSUBS 0.439188f
C2060 VDD2.n5 VSUBS 3.67599f
C2061 VN.t7 VSUBS 3.90978f
C2062 VN.n0 VSUBS 1.42834f
C2063 VN.n1 VSUBS 0.020759f
C2064 VN.n2 VSUBS 0.041753f
C2065 VN.n3 VSUBS 0.020759f
C2066 VN.n4 VSUBS 0.038689f
C2067 VN.n5 VSUBS 0.020759f
C2068 VN.t1 VSUBS 3.90978f
C2069 VN.n6 VSUBS 0.038689f
C2070 VN.n7 VSUBS 0.020759f
C2071 VN.n8 VSUBS 0.038689f
C2072 VN.t0 VSUBS 4.26261f
C2073 VN.n9 VSUBS 1.35899f
C2074 VN.t6 VSUBS 3.90978f
C2075 VN.n10 VSUBS 1.42705f
C2076 VN.n11 VSUBS 0.033341f
C2077 VN.n12 VSUBS 0.2687f
C2078 VN.n13 VSUBS 0.020759f
C2079 VN.n14 VSUBS 0.020759f
C2080 VN.n15 VSUBS 0.038689f
C2081 VN.n16 VSUBS 0.030304f
C2082 VN.n17 VSUBS 0.030304f
C2083 VN.n18 VSUBS 0.020759f
C2084 VN.n19 VSUBS 0.020759f
C2085 VN.n20 VSUBS 0.020759f
C2086 VN.n21 VSUBS 0.038689f
C2087 VN.n22 VSUBS 0.033341f
C2088 VN.n23 VSUBS 1.3475f
C2089 VN.n24 VSUBS 0.024936f
C2090 VN.n25 VSUBS 0.020759f
C2091 VN.n26 VSUBS 0.020759f
C2092 VN.n27 VSUBS 0.020759f
C2093 VN.n28 VSUBS 0.038689f
C2094 VN.n29 VSUBS 0.040521f
C2095 VN.n30 VSUBS 0.017023f
C2096 VN.n31 VSUBS 0.020759f
C2097 VN.n32 VSUBS 0.020759f
C2098 VN.n33 VSUBS 0.020759f
C2099 VN.n34 VSUBS 0.038689f
C2100 VN.n35 VSUBS 0.038689f
C2101 VN.n36 VSUBS 0.022644f
C2102 VN.n37 VSUBS 0.033504f
C2103 VN.n38 VSUBS 0.064146f
C2104 VN.t3 VSUBS 3.90978f
C2105 VN.n39 VSUBS 1.42834f
C2106 VN.n40 VSUBS 0.020759f
C2107 VN.n41 VSUBS 0.041753f
C2108 VN.n42 VSUBS 0.020759f
C2109 VN.n43 VSUBS 0.038689f
C2110 VN.n44 VSUBS 0.020759f
C2111 VN.t2 VSUBS 3.90978f
C2112 VN.n45 VSUBS 0.038689f
C2113 VN.n46 VSUBS 0.020759f
C2114 VN.n47 VSUBS 0.038689f
C2115 VN.t4 VSUBS 4.26261f
C2116 VN.n48 VSUBS 1.35899f
C2117 VN.t5 VSUBS 3.90978f
C2118 VN.n49 VSUBS 1.42705f
C2119 VN.n50 VSUBS 0.033341f
C2120 VN.n51 VSUBS 0.2687f
C2121 VN.n52 VSUBS 0.020759f
C2122 VN.n53 VSUBS 0.020759f
C2123 VN.n54 VSUBS 0.038689f
C2124 VN.n55 VSUBS 0.030304f
C2125 VN.n56 VSUBS 0.030304f
C2126 VN.n57 VSUBS 0.020759f
C2127 VN.n58 VSUBS 0.020759f
C2128 VN.n59 VSUBS 0.020759f
C2129 VN.n60 VSUBS 0.038689f
C2130 VN.n61 VSUBS 0.033341f
C2131 VN.n62 VSUBS 1.3475f
C2132 VN.n63 VSUBS 0.024936f
C2133 VN.n64 VSUBS 0.020759f
C2134 VN.n65 VSUBS 0.020759f
C2135 VN.n66 VSUBS 0.020759f
C2136 VN.n67 VSUBS 0.038689f
C2137 VN.n68 VSUBS 0.040521f
C2138 VN.n69 VSUBS 0.017023f
C2139 VN.n70 VSUBS 0.020759f
C2140 VN.n71 VSUBS 0.020759f
C2141 VN.n72 VSUBS 0.020759f
C2142 VN.n73 VSUBS 0.038689f
C2143 VN.n74 VSUBS 0.038689f
C2144 VN.n75 VSUBS 0.022644f
C2145 VN.n76 VSUBS 0.033504f
C2146 VN.n77 VSUBS 1.58618f
.ends

