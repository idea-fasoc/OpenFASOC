* NGSPICE file created from diff_pair_sample_1403.ext - technology: sky130A

.subckt diff_pair_sample_1403 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X1 VTAIL.t11 VN.t1 VDD2.t6 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X2 B.t11 B.t9 B.t10 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=0 ps=0 w=19.6 l=0.23
X3 VDD2.t5 VN.t2 VTAIL.t10 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=7.644 ps=39.98 w=19.6 l=0.23
X4 VDD1.t7 VP.t0 VTAIL.t2 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X5 VTAIL.t1 VP.t1 VDD1.t6 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X6 VTAIL.t15 VN.t3 VDD2.t4 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X7 VDD1.t5 VP.t2 VTAIL.t4 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=7.644 ps=39.98 w=19.6 l=0.23
X8 B.t8 B.t6 B.t7 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=0 ps=0 w=19.6 l=0.23
X9 VTAIL.t5 VP.t3 VDD1.t4 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=3.234 ps=19.93 w=19.6 l=0.23
X10 VTAIL.t6 VP.t4 VDD1.t3 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X11 VDD2.t3 VN.t4 VTAIL.t13 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=7.644 ps=39.98 w=19.6 l=0.23
X12 B.t5 B.t3 B.t4 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=0 ps=0 w=19.6 l=0.23
X13 VDD1.t2 VP.t5 VTAIL.t7 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X14 VTAIL.t0 VP.t6 VDD1.t1 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=3.234 ps=19.93 w=19.6 l=0.23
X15 VTAIL.t8 VN.t5 VDD2.t2 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=3.234 ps=19.93 w=19.6 l=0.23
X16 VTAIL.t14 VN.t6 VDD2.t1 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=3.234 ps=19.93 w=19.6 l=0.23
X17 B.t2 B.t0 B.t1 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=7.644 pd=39.98 as=0 ps=0 w=19.6 l=0.23
X18 VDD2.t0 VN.t7 VTAIL.t9 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=3.234 ps=19.93 w=19.6 l=0.23
X19 VDD1.t0 VP.t7 VTAIL.t3 w_n1530_n4888# sky130_fd_pr__pfet_01v8 ad=3.234 pd=19.93 as=7.644 ps=39.98 w=19.6 l=0.23
R0 VN.n5 VN.t2 2241.71
R1 VN.n1 VN.t6 2241.71
R2 VN.n12 VN.t5 2241.71
R3 VN.n8 VN.t4 2241.71
R4 VN.n4 VN.t1 2192.05
R5 VN.n2 VN.t7 2192.05
R6 VN.n11 VN.t0 2192.05
R7 VN.n9 VN.t3 2192.05
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN VN.n13 46.0403
R15 VN.n3 VN.n2 40.8975
R16 VN.n4 VN.n3 40.8975
R17 VN.n11 VN.n10 40.8975
R18 VN.n10 VN.n9 40.8975
R19 VN.n2 VN.n1 32.1338
R20 VN.n5 VN.n4 32.1338
R21 VN.n12 VN.n11 32.1338
R22 VN.n9 VN.n8 32.1338
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VTAIL.n882 VTAIL.n778 756.745
R27 VTAIL.n106 VTAIL.n2 756.745
R28 VTAIL.n216 VTAIL.n112 756.745
R29 VTAIL.n328 VTAIL.n224 756.745
R30 VTAIL.n772 VTAIL.n668 756.745
R31 VTAIL.n660 VTAIL.n556 756.745
R32 VTAIL.n550 VTAIL.n446 756.745
R33 VTAIL.n438 VTAIL.n334 756.745
R34 VTAIL.n815 VTAIL.n814 585
R35 VTAIL.n817 VTAIL.n816 585
R36 VTAIL.n810 VTAIL.n809 585
R37 VTAIL.n823 VTAIL.n822 585
R38 VTAIL.n825 VTAIL.n824 585
R39 VTAIL.n806 VTAIL.n805 585
R40 VTAIL.n831 VTAIL.n830 585
R41 VTAIL.n833 VTAIL.n832 585
R42 VTAIL.n802 VTAIL.n801 585
R43 VTAIL.n839 VTAIL.n838 585
R44 VTAIL.n841 VTAIL.n840 585
R45 VTAIL.n798 VTAIL.n797 585
R46 VTAIL.n847 VTAIL.n846 585
R47 VTAIL.n849 VTAIL.n848 585
R48 VTAIL.n794 VTAIL.n793 585
R49 VTAIL.n856 VTAIL.n855 585
R50 VTAIL.n857 VTAIL.n792 585
R51 VTAIL.n859 VTAIL.n858 585
R52 VTAIL.n790 VTAIL.n789 585
R53 VTAIL.n865 VTAIL.n864 585
R54 VTAIL.n867 VTAIL.n866 585
R55 VTAIL.n786 VTAIL.n785 585
R56 VTAIL.n873 VTAIL.n872 585
R57 VTAIL.n875 VTAIL.n874 585
R58 VTAIL.n782 VTAIL.n781 585
R59 VTAIL.n881 VTAIL.n880 585
R60 VTAIL.n883 VTAIL.n882 585
R61 VTAIL.n39 VTAIL.n38 585
R62 VTAIL.n41 VTAIL.n40 585
R63 VTAIL.n34 VTAIL.n33 585
R64 VTAIL.n47 VTAIL.n46 585
R65 VTAIL.n49 VTAIL.n48 585
R66 VTAIL.n30 VTAIL.n29 585
R67 VTAIL.n55 VTAIL.n54 585
R68 VTAIL.n57 VTAIL.n56 585
R69 VTAIL.n26 VTAIL.n25 585
R70 VTAIL.n63 VTAIL.n62 585
R71 VTAIL.n65 VTAIL.n64 585
R72 VTAIL.n22 VTAIL.n21 585
R73 VTAIL.n71 VTAIL.n70 585
R74 VTAIL.n73 VTAIL.n72 585
R75 VTAIL.n18 VTAIL.n17 585
R76 VTAIL.n80 VTAIL.n79 585
R77 VTAIL.n81 VTAIL.n16 585
R78 VTAIL.n83 VTAIL.n82 585
R79 VTAIL.n14 VTAIL.n13 585
R80 VTAIL.n89 VTAIL.n88 585
R81 VTAIL.n91 VTAIL.n90 585
R82 VTAIL.n10 VTAIL.n9 585
R83 VTAIL.n97 VTAIL.n96 585
R84 VTAIL.n99 VTAIL.n98 585
R85 VTAIL.n6 VTAIL.n5 585
R86 VTAIL.n105 VTAIL.n104 585
R87 VTAIL.n107 VTAIL.n106 585
R88 VTAIL.n149 VTAIL.n148 585
R89 VTAIL.n151 VTAIL.n150 585
R90 VTAIL.n144 VTAIL.n143 585
R91 VTAIL.n157 VTAIL.n156 585
R92 VTAIL.n159 VTAIL.n158 585
R93 VTAIL.n140 VTAIL.n139 585
R94 VTAIL.n165 VTAIL.n164 585
R95 VTAIL.n167 VTAIL.n166 585
R96 VTAIL.n136 VTAIL.n135 585
R97 VTAIL.n173 VTAIL.n172 585
R98 VTAIL.n175 VTAIL.n174 585
R99 VTAIL.n132 VTAIL.n131 585
R100 VTAIL.n181 VTAIL.n180 585
R101 VTAIL.n183 VTAIL.n182 585
R102 VTAIL.n128 VTAIL.n127 585
R103 VTAIL.n190 VTAIL.n189 585
R104 VTAIL.n191 VTAIL.n126 585
R105 VTAIL.n193 VTAIL.n192 585
R106 VTAIL.n124 VTAIL.n123 585
R107 VTAIL.n199 VTAIL.n198 585
R108 VTAIL.n201 VTAIL.n200 585
R109 VTAIL.n120 VTAIL.n119 585
R110 VTAIL.n207 VTAIL.n206 585
R111 VTAIL.n209 VTAIL.n208 585
R112 VTAIL.n116 VTAIL.n115 585
R113 VTAIL.n215 VTAIL.n214 585
R114 VTAIL.n217 VTAIL.n216 585
R115 VTAIL.n261 VTAIL.n260 585
R116 VTAIL.n263 VTAIL.n262 585
R117 VTAIL.n256 VTAIL.n255 585
R118 VTAIL.n269 VTAIL.n268 585
R119 VTAIL.n271 VTAIL.n270 585
R120 VTAIL.n252 VTAIL.n251 585
R121 VTAIL.n277 VTAIL.n276 585
R122 VTAIL.n279 VTAIL.n278 585
R123 VTAIL.n248 VTAIL.n247 585
R124 VTAIL.n285 VTAIL.n284 585
R125 VTAIL.n287 VTAIL.n286 585
R126 VTAIL.n244 VTAIL.n243 585
R127 VTAIL.n293 VTAIL.n292 585
R128 VTAIL.n295 VTAIL.n294 585
R129 VTAIL.n240 VTAIL.n239 585
R130 VTAIL.n302 VTAIL.n301 585
R131 VTAIL.n303 VTAIL.n238 585
R132 VTAIL.n305 VTAIL.n304 585
R133 VTAIL.n236 VTAIL.n235 585
R134 VTAIL.n311 VTAIL.n310 585
R135 VTAIL.n313 VTAIL.n312 585
R136 VTAIL.n232 VTAIL.n231 585
R137 VTAIL.n319 VTAIL.n318 585
R138 VTAIL.n321 VTAIL.n320 585
R139 VTAIL.n228 VTAIL.n227 585
R140 VTAIL.n327 VTAIL.n326 585
R141 VTAIL.n329 VTAIL.n328 585
R142 VTAIL.n773 VTAIL.n772 585
R143 VTAIL.n771 VTAIL.n770 585
R144 VTAIL.n672 VTAIL.n671 585
R145 VTAIL.n765 VTAIL.n764 585
R146 VTAIL.n763 VTAIL.n762 585
R147 VTAIL.n676 VTAIL.n675 585
R148 VTAIL.n757 VTAIL.n756 585
R149 VTAIL.n755 VTAIL.n754 585
R150 VTAIL.n680 VTAIL.n679 585
R151 VTAIL.n684 VTAIL.n682 585
R152 VTAIL.n749 VTAIL.n748 585
R153 VTAIL.n747 VTAIL.n746 585
R154 VTAIL.n686 VTAIL.n685 585
R155 VTAIL.n741 VTAIL.n740 585
R156 VTAIL.n739 VTAIL.n738 585
R157 VTAIL.n690 VTAIL.n689 585
R158 VTAIL.n733 VTAIL.n732 585
R159 VTAIL.n731 VTAIL.n730 585
R160 VTAIL.n694 VTAIL.n693 585
R161 VTAIL.n725 VTAIL.n724 585
R162 VTAIL.n723 VTAIL.n722 585
R163 VTAIL.n698 VTAIL.n697 585
R164 VTAIL.n717 VTAIL.n716 585
R165 VTAIL.n715 VTAIL.n714 585
R166 VTAIL.n702 VTAIL.n701 585
R167 VTAIL.n709 VTAIL.n708 585
R168 VTAIL.n707 VTAIL.n706 585
R169 VTAIL.n661 VTAIL.n660 585
R170 VTAIL.n659 VTAIL.n658 585
R171 VTAIL.n560 VTAIL.n559 585
R172 VTAIL.n653 VTAIL.n652 585
R173 VTAIL.n651 VTAIL.n650 585
R174 VTAIL.n564 VTAIL.n563 585
R175 VTAIL.n645 VTAIL.n644 585
R176 VTAIL.n643 VTAIL.n642 585
R177 VTAIL.n568 VTAIL.n567 585
R178 VTAIL.n572 VTAIL.n570 585
R179 VTAIL.n637 VTAIL.n636 585
R180 VTAIL.n635 VTAIL.n634 585
R181 VTAIL.n574 VTAIL.n573 585
R182 VTAIL.n629 VTAIL.n628 585
R183 VTAIL.n627 VTAIL.n626 585
R184 VTAIL.n578 VTAIL.n577 585
R185 VTAIL.n621 VTAIL.n620 585
R186 VTAIL.n619 VTAIL.n618 585
R187 VTAIL.n582 VTAIL.n581 585
R188 VTAIL.n613 VTAIL.n612 585
R189 VTAIL.n611 VTAIL.n610 585
R190 VTAIL.n586 VTAIL.n585 585
R191 VTAIL.n605 VTAIL.n604 585
R192 VTAIL.n603 VTAIL.n602 585
R193 VTAIL.n590 VTAIL.n589 585
R194 VTAIL.n597 VTAIL.n596 585
R195 VTAIL.n595 VTAIL.n594 585
R196 VTAIL.n551 VTAIL.n550 585
R197 VTAIL.n549 VTAIL.n548 585
R198 VTAIL.n450 VTAIL.n449 585
R199 VTAIL.n543 VTAIL.n542 585
R200 VTAIL.n541 VTAIL.n540 585
R201 VTAIL.n454 VTAIL.n453 585
R202 VTAIL.n535 VTAIL.n534 585
R203 VTAIL.n533 VTAIL.n532 585
R204 VTAIL.n458 VTAIL.n457 585
R205 VTAIL.n462 VTAIL.n460 585
R206 VTAIL.n527 VTAIL.n526 585
R207 VTAIL.n525 VTAIL.n524 585
R208 VTAIL.n464 VTAIL.n463 585
R209 VTAIL.n519 VTAIL.n518 585
R210 VTAIL.n517 VTAIL.n516 585
R211 VTAIL.n468 VTAIL.n467 585
R212 VTAIL.n511 VTAIL.n510 585
R213 VTAIL.n509 VTAIL.n508 585
R214 VTAIL.n472 VTAIL.n471 585
R215 VTAIL.n503 VTAIL.n502 585
R216 VTAIL.n501 VTAIL.n500 585
R217 VTAIL.n476 VTAIL.n475 585
R218 VTAIL.n495 VTAIL.n494 585
R219 VTAIL.n493 VTAIL.n492 585
R220 VTAIL.n480 VTAIL.n479 585
R221 VTAIL.n487 VTAIL.n486 585
R222 VTAIL.n485 VTAIL.n484 585
R223 VTAIL.n439 VTAIL.n438 585
R224 VTAIL.n437 VTAIL.n436 585
R225 VTAIL.n338 VTAIL.n337 585
R226 VTAIL.n431 VTAIL.n430 585
R227 VTAIL.n429 VTAIL.n428 585
R228 VTAIL.n342 VTAIL.n341 585
R229 VTAIL.n423 VTAIL.n422 585
R230 VTAIL.n421 VTAIL.n420 585
R231 VTAIL.n346 VTAIL.n345 585
R232 VTAIL.n350 VTAIL.n348 585
R233 VTAIL.n415 VTAIL.n414 585
R234 VTAIL.n413 VTAIL.n412 585
R235 VTAIL.n352 VTAIL.n351 585
R236 VTAIL.n407 VTAIL.n406 585
R237 VTAIL.n405 VTAIL.n404 585
R238 VTAIL.n356 VTAIL.n355 585
R239 VTAIL.n399 VTAIL.n398 585
R240 VTAIL.n397 VTAIL.n396 585
R241 VTAIL.n360 VTAIL.n359 585
R242 VTAIL.n391 VTAIL.n390 585
R243 VTAIL.n389 VTAIL.n388 585
R244 VTAIL.n364 VTAIL.n363 585
R245 VTAIL.n383 VTAIL.n382 585
R246 VTAIL.n381 VTAIL.n380 585
R247 VTAIL.n368 VTAIL.n367 585
R248 VTAIL.n375 VTAIL.n374 585
R249 VTAIL.n373 VTAIL.n372 585
R250 VTAIL.n813 VTAIL.t10 327.466
R251 VTAIL.n37 VTAIL.t14 327.466
R252 VTAIL.n147 VTAIL.t4 327.466
R253 VTAIL.n259 VTAIL.t0 327.466
R254 VTAIL.n705 VTAIL.t3 327.466
R255 VTAIL.n593 VTAIL.t5 327.466
R256 VTAIL.n483 VTAIL.t13 327.466
R257 VTAIL.n371 VTAIL.t8 327.466
R258 VTAIL.n816 VTAIL.n815 171.744
R259 VTAIL.n816 VTAIL.n809 171.744
R260 VTAIL.n823 VTAIL.n809 171.744
R261 VTAIL.n824 VTAIL.n823 171.744
R262 VTAIL.n824 VTAIL.n805 171.744
R263 VTAIL.n831 VTAIL.n805 171.744
R264 VTAIL.n832 VTAIL.n831 171.744
R265 VTAIL.n832 VTAIL.n801 171.744
R266 VTAIL.n839 VTAIL.n801 171.744
R267 VTAIL.n840 VTAIL.n839 171.744
R268 VTAIL.n840 VTAIL.n797 171.744
R269 VTAIL.n847 VTAIL.n797 171.744
R270 VTAIL.n848 VTAIL.n847 171.744
R271 VTAIL.n848 VTAIL.n793 171.744
R272 VTAIL.n856 VTAIL.n793 171.744
R273 VTAIL.n857 VTAIL.n856 171.744
R274 VTAIL.n858 VTAIL.n857 171.744
R275 VTAIL.n858 VTAIL.n789 171.744
R276 VTAIL.n865 VTAIL.n789 171.744
R277 VTAIL.n866 VTAIL.n865 171.744
R278 VTAIL.n866 VTAIL.n785 171.744
R279 VTAIL.n873 VTAIL.n785 171.744
R280 VTAIL.n874 VTAIL.n873 171.744
R281 VTAIL.n874 VTAIL.n781 171.744
R282 VTAIL.n881 VTAIL.n781 171.744
R283 VTAIL.n882 VTAIL.n881 171.744
R284 VTAIL.n40 VTAIL.n39 171.744
R285 VTAIL.n40 VTAIL.n33 171.744
R286 VTAIL.n47 VTAIL.n33 171.744
R287 VTAIL.n48 VTAIL.n47 171.744
R288 VTAIL.n48 VTAIL.n29 171.744
R289 VTAIL.n55 VTAIL.n29 171.744
R290 VTAIL.n56 VTAIL.n55 171.744
R291 VTAIL.n56 VTAIL.n25 171.744
R292 VTAIL.n63 VTAIL.n25 171.744
R293 VTAIL.n64 VTAIL.n63 171.744
R294 VTAIL.n64 VTAIL.n21 171.744
R295 VTAIL.n71 VTAIL.n21 171.744
R296 VTAIL.n72 VTAIL.n71 171.744
R297 VTAIL.n72 VTAIL.n17 171.744
R298 VTAIL.n80 VTAIL.n17 171.744
R299 VTAIL.n81 VTAIL.n80 171.744
R300 VTAIL.n82 VTAIL.n81 171.744
R301 VTAIL.n82 VTAIL.n13 171.744
R302 VTAIL.n89 VTAIL.n13 171.744
R303 VTAIL.n90 VTAIL.n89 171.744
R304 VTAIL.n90 VTAIL.n9 171.744
R305 VTAIL.n97 VTAIL.n9 171.744
R306 VTAIL.n98 VTAIL.n97 171.744
R307 VTAIL.n98 VTAIL.n5 171.744
R308 VTAIL.n105 VTAIL.n5 171.744
R309 VTAIL.n106 VTAIL.n105 171.744
R310 VTAIL.n150 VTAIL.n149 171.744
R311 VTAIL.n150 VTAIL.n143 171.744
R312 VTAIL.n157 VTAIL.n143 171.744
R313 VTAIL.n158 VTAIL.n157 171.744
R314 VTAIL.n158 VTAIL.n139 171.744
R315 VTAIL.n165 VTAIL.n139 171.744
R316 VTAIL.n166 VTAIL.n165 171.744
R317 VTAIL.n166 VTAIL.n135 171.744
R318 VTAIL.n173 VTAIL.n135 171.744
R319 VTAIL.n174 VTAIL.n173 171.744
R320 VTAIL.n174 VTAIL.n131 171.744
R321 VTAIL.n181 VTAIL.n131 171.744
R322 VTAIL.n182 VTAIL.n181 171.744
R323 VTAIL.n182 VTAIL.n127 171.744
R324 VTAIL.n190 VTAIL.n127 171.744
R325 VTAIL.n191 VTAIL.n190 171.744
R326 VTAIL.n192 VTAIL.n191 171.744
R327 VTAIL.n192 VTAIL.n123 171.744
R328 VTAIL.n199 VTAIL.n123 171.744
R329 VTAIL.n200 VTAIL.n199 171.744
R330 VTAIL.n200 VTAIL.n119 171.744
R331 VTAIL.n207 VTAIL.n119 171.744
R332 VTAIL.n208 VTAIL.n207 171.744
R333 VTAIL.n208 VTAIL.n115 171.744
R334 VTAIL.n215 VTAIL.n115 171.744
R335 VTAIL.n216 VTAIL.n215 171.744
R336 VTAIL.n262 VTAIL.n261 171.744
R337 VTAIL.n262 VTAIL.n255 171.744
R338 VTAIL.n269 VTAIL.n255 171.744
R339 VTAIL.n270 VTAIL.n269 171.744
R340 VTAIL.n270 VTAIL.n251 171.744
R341 VTAIL.n277 VTAIL.n251 171.744
R342 VTAIL.n278 VTAIL.n277 171.744
R343 VTAIL.n278 VTAIL.n247 171.744
R344 VTAIL.n285 VTAIL.n247 171.744
R345 VTAIL.n286 VTAIL.n285 171.744
R346 VTAIL.n286 VTAIL.n243 171.744
R347 VTAIL.n293 VTAIL.n243 171.744
R348 VTAIL.n294 VTAIL.n293 171.744
R349 VTAIL.n294 VTAIL.n239 171.744
R350 VTAIL.n302 VTAIL.n239 171.744
R351 VTAIL.n303 VTAIL.n302 171.744
R352 VTAIL.n304 VTAIL.n303 171.744
R353 VTAIL.n304 VTAIL.n235 171.744
R354 VTAIL.n311 VTAIL.n235 171.744
R355 VTAIL.n312 VTAIL.n311 171.744
R356 VTAIL.n312 VTAIL.n231 171.744
R357 VTAIL.n319 VTAIL.n231 171.744
R358 VTAIL.n320 VTAIL.n319 171.744
R359 VTAIL.n320 VTAIL.n227 171.744
R360 VTAIL.n327 VTAIL.n227 171.744
R361 VTAIL.n328 VTAIL.n327 171.744
R362 VTAIL.n772 VTAIL.n771 171.744
R363 VTAIL.n771 VTAIL.n671 171.744
R364 VTAIL.n764 VTAIL.n671 171.744
R365 VTAIL.n764 VTAIL.n763 171.744
R366 VTAIL.n763 VTAIL.n675 171.744
R367 VTAIL.n756 VTAIL.n675 171.744
R368 VTAIL.n756 VTAIL.n755 171.744
R369 VTAIL.n755 VTAIL.n679 171.744
R370 VTAIL.n684 VTAIL.n679 171.744
R371 VTAIL.n748 VTAIL.n684 171.744
R372 VTAIL.n748 VTAIL.n747 171.744
R373 VTAIL.n747 VTAIL.n685 171.744
R374 VTAIL.n740 VTAIL.n685 171.744
R375 VTAIL.n740 VTAIL.n739 171.744
R376 VTAIL.n739 VTAIL.n689 171.744
R377 VTAIL.n732 VTAIL.n689 171.744
R378 VTAIL.n732 VTAIL.n731 171.744
R379 VTAIL.n731 VTAIL.n693 171.744
R380 VTAIL.n724 VTAIL.n693 171.744
R381 VTAIL.n724 VTAIL.n723 171.744
R382 VTAIL.n723 VTAIL.n697 171.744
R383 VTAIL.n716 VTAIL.n697 171.744
R384 VTAIL.n716 VTAIL.n715 171.744
R385 VTAIL.n715 VTAIL.n701 171.744
R386 VTAIL.n708 VTAIL.n701 171.744
R387 VTAIL.n708 VTAIL.n707 171.744
R388 VTAIL.n660 VTAIL.n659 171.744
R389 VTAIL.n659 VTAIL.n559 171.744
R390 VTAIL.n652 VTAIL.n559 171.744
R391 VTAIL.n652 VTAIL.n651 171.744
R392 VTAIL.n651 VTAIL.n563 171.744
R393 VTAIL.n644 VTAIL.n563 171.744
R394 VTAIL.n644 VTAIL.n643 171.744
R395 VTAIL.n643 VTAIL.n567 171.744
R396 VTAIL.n572 VTAIL.n567 171.744
R397 VTAIL.n636 VTAIL.n572 171.744
R398 VTAIL.n636 VTAIL.n635 171.744
R399 VTAIL.n635 VTAIL.n573 171.744
R400 VTAIL.n628 VTAIL.n573 171.744
R401 VTAIL.n628 VTAIL.n627 171.744
R402 VTAIL.n627 VTAIL.n577 171.744
R403 VTAIL.n620 VTAIL.n577 171.744
R404 VTAIL.n620 VTAIL.n619 171.744
R405 VTAIL.n619 VTAIL.n581 171.744
R406 VTAIL.n612 VTAIL.n581 171.744
R407 VTAIL.n612 VTAIL.n611 171.744
R408 VTAIL.n611 VTAIL.n585 171.744
R409 VTAIL.n604 VTAIL.n585 171.744
R410 VTAIL.n604 VTAIL.n603 171.744
R411 VTAIL.n603 VTAIL.n589 171.744
R412 VTAIL.n596 VTAIL.n589 171.744
R413 VTAIL.n596 VTAIL.n595 171.744
R414 VTAIL.n550 VTAIL.n549 171.744
R415 VTAIL.n549 VTAIL.n449 171.744
R416 VTAIL.n542 VTAIL.n449 171.744
R417 VTAIL.n542 VTAIL.n541 171.744
R418 VTAIL.n541 VTAIL.n453 171.744
R419 VTAIL.n534 VTAIL.n453 171.744
R420 VTAIL.n534 VTAIL.n533 171.744
R421 VTAIL.n533 VTAIL.n457 171.744
R422 VTAIL.n462 VTAIL.n457 171.744
R423 VTAIL.n526 VTAIL.n462 171.744
R424 VTAIL.n526 VTAIL.n525 171.744
R425 VTAIL.n525 VTAIL.n463 171.744
R426 VTAIL.n518 VTAIL.n463 171.744
R427 VTAIL.n518 VTAIL.n517 171.744
R428 VTAIL.n517 VTAIL.n467 171.744
R429 VTAIL.n510 VTAIL.n467 171.744
R430 VTAIL.n510 VTAIL.n509 171.744
R431 VTAIL.n509 VTAIL.n471 171.744
R432 VTAIL.n502 VTAIL.n471 171.744
R433 VTAIL.n502 VTAIL.n501 171.744
R434 VTAIL.n501 VTAIL.n475 171.744
R435 VTAIL.n494 VTAIL.n475 171.744
R436 VTAIL.n494 VTAIL.n493 171.744
R437 VTAIL.n493 VTAIL.n479 171.744
R438 VTAIL.n486 VTAIL.n479 171.744
R439 VTAIL.n486 VTAIL.n485 171.744
R440 VTAIL.n438 VTAIL.n437 171.744
R441 VTAIL.n437 VTAIL.n337 171.744
R442 VTAIL.n430 VTAIL.n337 171.744
R443 VTAIL.n430 VTAIL.n429 171.744
R444 VTAIL.n429 VTAIL.n341 171.744
R445 VTAIL.n422 VTAIL.n341 171.744
R446 VTAIL.n422 VTAIL.n421 171.744
R447 VTAIL.n421 VTAIL.n345 171.744
R448 VTAIL.n350 VTAIL.n345 171.744
R449 VTAIL.n414 VTAIL.n350 171.744
R450 VTAIL.n414 VTAIL.n413 171.744
R451 VTAIL.n413 VTAIL.n351 171.744
R452 VTAIL.n406 VTAIL.n351 171.744
R453 VTAIL.n406 VTAIL.n405 171.744
R454 VTAIL.n405 VTAIL.n355 171.744
R455 VTAIL.n398 VTAIL.n355 171.744
R456 VTAIL.n398 VTAIL.n397 171.744
R457 VTAIL.n397 VTAIL.n359 171.744
R458 VTAIL.n390 VTAIL.n359 171.744
R459 VTAIL.n390 VTAIL.n389 171.744
R460 VTAIL.n389 VTAIL.n363 171.744
R461 VTAIL.n382 VTAIL.n363 171.744
R462 VTAIL.n382 VTAIL.n381 171.744
R463 VTAIL.n381 VTAIL.n367 171.744
R464 VTAIL.n374 VTAIL.n367 171.744
R465 VTAIL.n374 VTAIL.n373 171.744
R466 VTAIL.n815 VTAIL.t10 85.8723
R467 VTAIL.n39 VTAIL.t14 85.8723
R468 VTAIL.n149 VTAIL.t4 85.8723
R469 VTAIL.n261 VTAIL.t0 85.8723
R470 VTAIL.n707 VTAIL.t3 85.8723
R471 VTAIL.n595 VTAIL.t5 85.8723
R472 VTAIL.n485 VTAIL.t13 85.8723
R473 VTAIL.n373 VTAIL.t8 85.8723
R474 VTAIL.n667 VTAIL.n666 49.8795
R475 VTAIL.n445 VTAIL.n444 49.8795
R476 VTAIL.n1 VTAIL.n0 49.8793
R477 VTAIL.n223 VTAIL.n222 49.8793
R478 VTAIL.n887 VTAIL.n886 30.6338
R479 VTAIL.n111 VTAIL.n110 30.6338
R480 VTAIL.n221 VTAIL.n220 30.6338
R481 VTAIL.n333 VTAIL.n332 30.6338
R482 VTAIL.n777 VTAIL.n776 30.6338
R483 VTAIL.n665 VTAIL.n664 30.6338
R484 VTAIL.n555 VTAIL.n554 30.6338
R485 VTAIL.n443 VTAIL.n442 30.6338
R486 VTAIL.n887 VTAIL.n777 29.7462
R487 VTAIL.n443 VTAIL.n333 29.7462
R488 VTAIL.n814 VTAIL.n813 16.3895
R489 VTAIL.n38 VTAIL.n37 16.3895
R490 VTAIL.n148 VTAIL.n147 16.3895
R491 VTAIL.n260 VTAIL.n259 16.3895
R492 VTAIL.n706 VTAIL.n705 16.3895
R493 VTAIL.n594 VTAIL.n593 16.3895
R494 VTAIL.n484 VTAIL.n483 16.3895
R495 VTAIL.n372 VTAIL.n371 16.3895
R496 VTAIL.n859 VTAIL.n790 13.1884
R497 VTAIL.n83 VTAIL.n14 13.1884
R498 VTAIL.n193 VTAIL.n124 13.1884
R499 VTAIL.n305 VTAIL.n236 13.1884
R500 VTAIL.n682 VTAIL.n680 13.1884
R501 VTAIL.n570 VTAIL.n568 13.1884
R502 VTAIL.n460 VTAIL.n458 13.1884
R503 VTAIL.n348 VTAIL.n346 13.1884
R504 VTAIL.n817 VTAIL.n812 12.8005
R505 VTAIL.n860 VTAIL.n792 12.8005
R506 VTAIL.n864 VTAIL.n863 12.8005
R507 VTAIL.n41 VTAIL.n36 12.8005
R508 VTAIL.n84 VTAIL.n16 12.8005
R509 VTAIL.n88 VTAIL.n87 12.8005
R510 VTAIL.n151 VTAIL.n146 12.8005
R511 VTAIL.n194 VTAIL.n126 12.8005
R512 VTAIL.n198 VTAIL.n197 12.8005
R513 VTAIL.n263 VTAIL.n258 12.8005
R514 VTAIL.n306 VTAIL.n238 12.8005
R515 VTAIL.n310 VTAIL.n309 12.8005
R516 VTAIL.n754 VTAIL.n753 12.8005
R517 VTAIL.n750 VTAIL.n749 12.8005
R518 VTAIL.n709 VTAIL.n704 12.8005
R519 VTAIL.n642 VTAIL.n641 12.8005
R520 VTAIL.n638 VTAIL.n637 12.8005
R521 VTAIL.n597 VTAIL.n592 12.8005
R522 VTAIL.n532 VTAIL.n531 12.8005
R523 VTAIL.n528 VTAIL.n527 12.8005
R524 VTAIL.n487 VTAIL.n482 12.8005
R525 VTAIL.n420 VTAIL.n419 12.8005
R526 VTAIL.n416 VTAIL.n415 12.8005
R527 VTAIL.n375 VTAIL.n370 12.8005
R528 VTAIL.n818 VTAIL.n810 12.0247
R529 VTAIL.n855 VTAIL.n854 12.0247
R530 VTAIL.n867 VTAIL.n788 12.0247
R531 VTAIL.n42 VTAIL.n34 12.0247
R532 VTAIL.n79 VTAIL.n78 12.0247
R533 VTAIL.n91 VTAIL.n12 12.0247
R534 VTAIL.n152 VTAIL.n144 12.0247
R535 VTAIL.n189 VTAIL.n188 12.0247
R536 VTAIL.n201 VTAIL.n122 12.0247
R537 VTAIL.n264 VTAIL.n256 12.0247
R538 VTAIL.n301 VTAIL.n300 12.0247
R539 VTAIL.n313 VTAIL.n234 12.0247
R540 VTAIL.n757 VTAIL.n678 12.0247
R541 VTAIL.n746 VTAIL.n683 12.0247
R542 VTAIL.n710 VTAIL.n702 12.0247
R543 VTAIL.n645 VTAIL.n566 12.0247
R544 VTAIL.n634 VTAIL.n571 12.0247
R545 VTAIL.n598 VTAIL.n590 12.0247
R546 VTAIL.n535 VTAIL.n456 12.0247
R547 VTAIL.n524 VTAIL.n461 12.0247
R548 VTAIL.n488 VTAIL.n480 12.0247
R549 VTAIL.n423 VTAIL.n344 12.0247
R550 VTAIL.n412 VTAIL.n349 12.0247
R551 VTAIL.n376 VTAIL.n368 12.0247
R552 VTAIL.n822 VTAIL.n821 11.249
R553 VTAIL.n853 VTAIL.n794 11.249
R554 VTAIL.n868 VTAIL.n786 11.249
R555 VTAIL.n46 VTAIL.n45 11.249
R556 VTAIL.n77 VTAIL.n18 11.249
R557 VTAIL.n92 VTAIL.n10 11.249
R558 VTAIL.n156 VTAIL.n155 11.249
R559 VTAIL.n187 VTAIL.n128 11.249
R560 VTAIL.n202 VTAIL.n120 11.249
R561 VTAIL.n268 VTAIL.n267 11.249
R562 VTAIL.n299 VTAIL.n240 11.249
R563 VTAIL.n314 VTAIL.n232 11.249
R564 VTAIL.n758 VTAIL.n676 11.249
R565 VTAIL.n745 VTAIL.n686 11.249
R566 VTAIL.n714 VTAIL.n713 11.249
R567 VTAIL.n646 VTAIL.n564 11.249
R568 VTAIL.n633 VTAIL.n574 11.249
R569 VTAIL.n602 VTAIL.n601 11.249
R570 VTAIL.n536 VTAIL.n454 11.249
R571 VTAIL.n523 VTAIL.n464 11.249
R572 VTAIL.n492 VTAIL.n491 11.249
R573 VTAIL.n424 VTAIL.n342 11.249
R574 VTAIL.n411 VTAIL.n352 11.249
R575 VTAIL.n380 VTAIL.n379 11.249
R576 VTAIL.n825 VTAIL.n808 10.4732
R577 VTAIL.n850 VTAIL.n849 10.4732
R578 VTAIL.n872 VTAIL.n871 10.4732
R579 VTAIL.n49 VTAIL.n32 10.4732
R580 VTAIL.n74 VTAIL.n73 10.4732
R581 VTAIL.n96 VTAIL.n95 10.4732
R582 VTAIL.n159 VTAIL.n142 10.4732
R583 VTAIL.n184 VTAIL.n183 10.4732
R584 VTAIL.n206 VTAIL.n205 10.4732
R585 VTAIL.n271 VTAIL.n254 10.4732
R586 VTAIL.n296 VTAIL.n295 10.4732
R587 VTAIL.n318 VTAIL.n317 10.4732
R588 VTAIL.n762 VTAIL.n761 10.4732
R589 VTAIL.n742 VTAIL.n741 10.4732
R590 VTAIL.n717 VTAIL.n700 10.4732
R591 VTAIL.n650 VTAIL.n649 10.4732
R592 VTAIL.n630 VTAIL.n629 10.4732
R593 VTAIL.n605 VTAIL.n588 10.4732
R594 VTAIL.n540 VTAIL.n539 10.4732
R595 VTAIL.n520 VTAIL.n519 10.4732
R596 VTAIL.n495 VTAIL.n478 10.4732
R597 VTAIL.n428 VTAIL.n427 10.4732
R598 VTAIL.n408 VTAIL.n407 10.4732
R599 VTAIL.n383 VTAIL.n366 10.4732
R600 VTAIL.n826 VTAIL.n806 9.69747
R601 VTAIL.n846 VTAIL.n796 9.69747
R602 VTAIL.n875 VTAIL.n784 9.69747
R603 VTAIL.n50 VTAIL.n30 9.69747
R604 VTAIL.n70 VTAIL.n20 9.69747
R605 VTAIL.n99 VTAIL.n8 9.69747
R606 VTAIL.n160 VTAIL.n140 9.69747
R607 VTAIL.n180 VTAIL.n130 9.69747
R608 VTAIL.n209 VTAIL.n118 9.69747
R609 VTAIL.n272 VTAIL.n252 9.69747
R610 VTAIL.n292 VTAIL.n242 9.69747
R611 VTAIL.n321 VTAIL.n230 9.69747
R612 VTAIL.n765 VTAIL.n674 9.69747
R613 VTAIL.n738 VTAIL.n688 9.69747
R614 VTAIL.n718 VTAIL.n698 9.69747
R615 VTAIL.n653 VTAIL.n562 9.69747
R616 VTAIL.n626 VTAIL.n576 9.69747
R617 VTAIL.n606 VTAIL.n586 9.69747
R618 VTAIL.n543 VTAIL.n452 9.69747
R619 VTAIL.n516 VTAIL.n466 9.69747
R620 VTAIL.n496 VTAIL.n476 9.69747
R621 VTAIL.n431 VTAIL.n340 9.69747
R622 VTAIL.n404 VTAIL.n354 9.69747
R623 VTAIL.n384 VTAIL.n364 9.69747
R624 VTAIL.n886 VTAIL.n885 9.45567
R625 VTAIL.n110 VTAIL.n109 9.45567
R626 VTAIL.n220 VTAIL.n219 9.45567
R627 VTAIL.n332 VTAIL.n331 9.45567
R628 VTAIL.n776 VTAIL.n775 9.45567
R629 VTAIL.n664 VTAIL.n663 9.45567
R630 VTAIL.n554 VTAIL.n553 9.45567
R631 VTAIL.n442 VTAIL.n441 9.45567
R632 VTAIL.n885 VTAIL.n884 9.3005
R633 VTAIL.n879 VTAIL.n878 9.3005
R634 VTAIL.n877 VTAIL.n876 9.3005
R635 VTAIL.n784 VTAIL.n783 9.3005
R636 VTAIL.n871 VTAIL.n870 9.3005
R637 VTAIL.n869 VTAIL.n868 9.3005
R638 VTAIL.n788 VTAIL.n787 9.3005
R639 VTAIL.n863 VTAIL.n862 9.3005
R640 VTAIL.n835 VTAIL.n834 9.3005
R641 VTAIL.n804 VTAIL.n803 9.3005
R642 VTAIL.n829 VTAIL.n828 9.3005
R643 VTAIL.n827 VTAIL.n826 9.3005
R644 VTAIL.n808 VTAIL.n807 9.3005
R645 VTAIL.n821 VTAIL.n820 9.3005
R646 VTAIL.n819 VTAIL.n818 9.3005
R647 VTAIL.n812 VTAIL.n811 9.3005
R648 VTAIL.n837 VTAIL.n836 9.3005
R649 VTAIL.n800 VTAIL.n799 9.3005
R650 VTAIL.n843 VTAIL.n842 9.3005
R651 VTAIL.n845 VTAIL.n844 9.3005
R652 VTAIL.n796 VTAIL.n795 9.3005
R653 VTAIL.n851 VTAIL.n850 9.3005
R654 VTAIL.n853 VTAIL.n852 9.3005
R655 VTAIL.n854 VTAIL.n791 9.3005
R656 VTAIL.n861 VTAIL.n860 9.3005
R657 VTAIL.n780 VTAIL.n779 9.3005
R658 VTAIL.n109 VTAIL.n108 9.3005
R659 VTAIL.n103 VTAIL.n102 9.3005
R660 VTAIL.n101 VTAIL.n100 9.3005
R661 VTAIL.n8 VTAIL.n7 9.3005
R662 VTAIL.n95 VTAIL.n94 9.3005
R663 VTAIL.n93 VTAIL.n92 9.3005
R664 VTAIL.n12 VTAIL.n11 9.3005
R665 VTAIL.n87 VTAIL.n86 9.3005
R666 VTAIL.n59 VTAIL.n58 9.3005
R667 VTAIL.n28 VTAIL.n27 9.3005
R668 VTAIL.n53 VTAIL.n52 9.3005
R669 VTAIL.n51 VTAIL.n50 9.3005
R670 VTAIL.n32 VTAIL.n31 9.3005
R671 VTAIL.n45 VTAIL.n44 9.3005
R672 VTAIL.n43 VTAIL.n42 9.3005
R673 VTAIL.n36 VTAIL.n35 9.3005
R674 VTAIL.n61 VTAIL.n60 9.3005
R675 VTAIL.n24 VTAIL.n23 9.3005
R676 VTAIL.n67 VTAIL.n66 9.3005
R677 VTAIL.n69 VTAIL.n68 9.3005
R678 VTAIL.n20 VTAIL.n19 9.3005
R679 VTAIL.n75 VTAIL.n74 9.3005
R680 VTAIL.n77 VTAIL.n76 9.3005
R681 VTAIL.n78 VTAIL.n15 9.3005
R682 VTAIL.n85 VTAIL.n84 9.3005
R683 VTAIL.n4 VTAIL.n3 9.3005
R684 VTAIL.n219 VTAIL.n218 9.3005
R685 VTAIL.n213 VTAIL.n212 9.3005
R686 VTAIL.n211 VTAIL.n210 9.3005
R687 VTAIL.n118 VTAIL.n117 9.3005
R688 VTAIL.n205 VTAIL.n204 9.3005
R689 VTAIL.n203 VTAIL.n202 9.3005
R690 VTAIL.n122 VTAIL.n121 9.3005
R691 VTAIL.n197 VTAIL.n196 9.3005
R692 VTAIL.n169 VTAIL.n168 9.3005
R693 VTAIL.n138 VTAIL.n137 9.3005
R694 VTAIL.n163 VTAIL.n162 9.3005
R695 VTAIL.n161 VTAIL.n160 9.3005
R696 VTAIL.n142 VTAIL.n141 9.3005
R697 VTAIL.n155 VTAIL.n154 9.3005
R698 VTAIL.n153 VTAIL.n152 9.3005
R699 VTAIL.n146 VTAIL.n145 9.3005
R700 VTAIL.n171 VTAIL.n170 9.3005
R701 VTAIL.n134 VTAIL.n133 9.3005
R702 VTAIL.n177 VTAIL.n176 9.3005
R703 VTAIL.n179 VTAIL.n178 9.3005
R704 VTAIL.n130 VTAIL.n129 9.3005
R705 VTAIL.n185 VTAIL.n184 9.3005
R706 VTAIL.n187 VTAIL.n186 9.3005
R707 VTAIL.n188 VTAIL.n125 9.3005
R708 VTAIL.n195 VTAIL.n194 9.3005
R709 VTAIL.n114 VTAIL.n113 9.3005
R710 VTAIL.n331 VTAIL.n330 9.3005
R711 VTAIL.n325 VTAIL.n324 9.3005
R712 VTAIL.n323 VTAIL.n322 9.3005
R713 VTAIL.n230 VTAIL.n229 9.3005
R714 VTAIL.n317 VTAIL.n316 9.3005
R715 VTAIL.n315 VTAIL.n314 9.3005
R716 VTAIL.n234 VTAIL.n233 9.3005
R717 VTAIL.n309 VTAIL.n308 9.3005
R718 VTAIL.n281 VTAIL.n280 9.3005
R719 VTAIL.n250 VTAIL.n249 9.3005
R720 VTAIL.n275 VTAIL.n274 9.3005
R721 VTAIL.n273 VTAIL.n272 9.3005
R722 VTAIL.n254 VTAIL.n253 9.3005
R723 VTAIL.n267 VTAIL.n266 9.3005
R724 VTAIL.n265 VTAIL.n264 9.3005
R725 VTAIL.n258 VTAIL.n257 9.3005
R726 VTAIL.n283 VTAIL.n282 9.3005
R727 VTAIL.n246 VTAIL.n245 9.3005
R728 VTAIL.n289 VTAIL.n288 9.3005
R729 VTAIL.n291 VTAIL.n290 9.3005
R730 VTAIL.n242 VTAIL.n241 9.3005
R731 VTAIL.n297 VTAIL.n296 9.3005
R732 VTAIL.n299 VTAIL.n298 9.3005
R733 VTAIL.n300 VTAIL.n237 9.3005
R734 VTAIL.n307 VTAIL.n306 9.3005
R735 VTAIL.n226 VTAIL.n225 9.3005
R736 VTAIL.n692 VTAIL.n691 9.3005
R737 VTAIL.n735 VTAIL.n734 9.3005
R738 VTAIL.n737 VTAIL.n736 9.3005
R739 VTAIL.n688 VTAIL.n687 9.3005
R740 VTAIL.n743 VTAIL.n742 9.3005
R741 VTAIL.n745 VTAIL.n744 9.3005
R742 VTAIL.n683 VTAIL.n681 9.3005
R743 VTAIL.n751 VTAIL.n750 9.3005
R744 VTAIL.n775 VTAIL.n774 9.3005
R745 VTAIL.n670 VTAIL.n669 9.3005
R746 VTAIL.n769 VTAIL.n768 9.3005
R747 VTAIL.n767 VTAIL.n766 9.3005
R748 VTAIL.n674 VTAIL.n673 9.3005
R749 VTAIL.n761 VTAIL.n760 9.3005
R750 VTAIL.n759 VTAIL.n758 9.3005
R751 VTAIL.n678 VTAIL.n677 9.3005
R752 VTAIL.n753 VTAIL.n752 9.3005
R753 VTAIL.n729 VTAIL.n728 9.3005
R754 VTAIL.n727 VTAIL.n726 9.3005
R755 VTAIL.n696 VTAIL.n695 9.3005
R756 VTAIL.n721 VTAIL.n720 9.3005
R757 VTAIL.n719 VTAIL.n718 9.3005
R758 VTAIL.n700 VTAIL.n699 9.3005
R759 VTAIL.n713 VTAIL.n712 9.3005
R760 VTAIL.n711 VTAIL.n710 9.3005
R761 VTAIL.n704 VTAIL.n703 9.3005
R762 VTAIL.n580 VTAIL.n579 9.3005
R763 VTAIL.n623 VTAIL.n622 9.3005
R764 VTAIL.n625 VTAIL.n624 9.3005
R765 VTAIL.n576 VTAIL.n575 9.3005
R766 VTAIL.n631 VTAIL.n630 9.3005
R767 VTAIL.n633 VTAIL.n632 9.3005
R768 VTAIL.n571 VTAIL.n569 9.3005
R769 VTAIL.n639 VTAIL.n638 9.3005
R770 VTAIL.n663 VTAIL.n662 9.3005
R771 VTAIL.n558 VTAIL.n557 9.3005
R772 VTAIL.n657 VTAIL.n656 9.3005
R773 VTAIL.n655 VTAIL.n654 9.3005
R774 VTAIL.n562 VTAIL.n561 9.3005
R775 VTAIL.n649 VTAIL.n648 9.3005
R776 VTAIL.n647 VTAIL.n646 9.3005
R777 VTAIL.n566 VTAIL.n565 9.3005
R778 VTAIL.n641 VTAIL.n640 9.3005
R779 VTAIL.n617 VTAIL.n616 9.3005
R780 VTAIL.n615 VTAIL.n614 9.3005
R781 VTAIL.n584 VTAIL.n583 9.3005
R782 VTAIL.n609 VTAIL.n608 9.3005
R783 VTAIL.n607 VTAIL.n606 9.3005
R784 VTAIL.n588 VTAIL.n587 9.3005
R785 VTAIL.n601 VTAIL.n600 9.3005
R786 VTAIL.n599 VTAIL.n598 9.3005
R787 VTAIL.n592 VTAIL.n591 9.3005
R788 VTAIL.n470 VTAIL.n469 9.3005
R789 VTAIL.n513 VTAIL.n512 9.3005
R790 VTAIL.n515 VTAIL.n514 9.3005
R791 VTAIL.n466 VTAIL.n465 9.3005
R792 VTAIL.n521 VTAIL.n520 9.3005
R793 VTAIL.n523 VTAIL.n522 9.3005
R794 VTAIL.n461 VTAIL.n459 9.3005
R795 VTAIL.n529 VTAIL.n528 9.3005
R796 VTAIL.n553 VTAIL.n552 9.3005
R797 VTAIL.n448 VTAIL.n447 9.3005
R798 VTAIL.n547 VTAIL.n546 9.3005
R799 VTAIL.n545 VTAIL.n544 9.3005
R800 VTAIL.n452 VTAIL.n451 9.3005
R801 VTAIL.n539 VTAIL.n538 9.3005
R802 VTAIL.n537 VTAIL.n536 9.3005
R803 VTAIL.n456 VTAIL.n455 9.3005
R804 VTAIL.n531 VTAIL.n530 9.3005
R805 VTAIL.n507 VTAIL.n506 9.3005
R806 VTAIL.n505 VTAIL.n504 9.3005
R807 VTAIL.n474 VTAIL.n473 9.3005
R808 VTAIL.n499 VTAIL.n498 9.3005
R809 VTAIL.n497 VTAIL.n496 9.3005
R810 VTAIL.n478 VTAIL.n477 9.3005
R811 VTAIL.n491 VTAIL.n490 9.3005
R812 VTAIL.n489 VTAIL.n488 9.3005
R813 VTAIL.n482 VTAIL.n481 9.3005
R814 VTAIL.n358 VTAIL.n357 9.3005
R815 VTAIL.n401 VTAIL.n400 9.3005
R816 VTAIL.n403 VTAIL.n402 9.3005
R817 VTAIL.n354 VTAIL.n353 9.3005
R818 VTAIL.n409 VTAIL.n408 9.3005
R819 VTAIL.n411 VTAIL.n410 9.3005
R820 VTAIL.n349 VTAIL.n347 9.3005
R821 VTAIL.n417 VTAIL.n416 9.3005
R822 VTAIL.n441 VTAIL.n440 9.3005
R823 VTAIL.n336 VTAIL.n335 9.3005
R824 VTAIL.n435 VTAIL.n434 9.3005
R825 VTAIL.n433 VTAIL.n432 9.3005
R826 VTAIL.n340 VTAIL.n339 9.3005
R827 VTAIL.n427 VTAIL.n426 9.3005
R828 VTAIL.n425 VTAIL.n424 9.3005
R829 VTAIL.n344 VTAIL.n343 9.3005
R830 VTAIL.n419 VTAIL.n418 9.3005
R831 VTAIL.n395 VTAIL.n394 9.3005
R832 VTAIL.n393 VTAIL.n392 9.3005
R833 VTAIL.n362 VTAIL.n361 9.3005
R834 VTAIL.n387 VTAIL.n386 9.3005
R835 VTAIL.n385 VTAIL.n384 9.3005
R836 VTAIL.n366 VTAIL.n365 9.3005
R837 VTAIL.n379 VTAIL.n378 9.3005
R838 VTAIL.n377 VTAIL.n376 9.3005
R839 VTAIL.n370 VTAIL.n369 9.3005
R840 VTAIL.n830 VTAIL.n829 8.92171
R841 VTAIL.n845 VTAIL.n798 8.92171
R842 VTAIL.n876 VTAIL.n782 8.92171
R843 VTAIL.n54 VTAIL.n53 8.92171
R844 VTAIL.n69 VTAIL.n22 8.92171
R845 VTAIL.n100 VTAIL.n6 8.92171
R846 VTAIL.n164 VTAIL.n163 8.92171
R847 VTAIL.n179 VTAIL.n132 8.92171
R848 VTAIL.n210 VTAIL.n116 8.92171
R849 VTAIL.n276 VTAIL.n275 8.92171
R850 VTAIL.n291 VTAIL.n244 8.92171
R851 VTAIL.n322 VTAIL.n228 8.92171
R852 VTAIL.n766 VTAIL.n672 8.92171
R853 VTAIL.n737 VTAIL.n690 8.92171
R854 VTAIL.n722 VTAIL.n721 8.92171
R855 VTAIL.n654 VTAIL.n560 8.92171
R856 VTAIL.n625 VTAIL.n578 8.92171
R857 VTAIL.n610 VTAIL.n609 8.92171
R858 VTAIL.n544 VTAIL.n450 8.92171
R859 VTAIL.n515 VTAIL.n468 8.92171
R860 VTAIL.n500 VTAIL.n499 8.92171
R861 VTAIL.n432 VTAIL.n338 8.92171
R862 VTAIL.n403 VTAIL.n356 8.92171
R863 VTAIL.n388 VTAIL.n387 8.92171
R864 VTAIL.n833 VTAIL.n804 8.14595
R865 VTAIL.n842 VTAIL.n841 8.14595
R866 VTAIL.n880 VTAIL.n879 8.14595
R867 VTAIL.n57 VTAIL.n28 8.14595
R868 VTAIL.n66 VTAIL.n65 8.14595
R869 VTAIL.n104 VTAIL.n103 8.14595
R870 VTAIL.n167 VTAIL.n138 8.14595
R871 VTAIL.n176 VTAIL.n175 8.14595
R872 VTAIL.n214 VTAIL.n213 8.14595
R873 VTAIL.n279 VTAIL.n250 8.14595
R874 VTAIL.n288 VTAIL.n287 8.14595
R875 VTAIL.n326 VTAIL.n325 8.14595
R876 VTAIL.n770 VTAIL.n769 8.14595
R877 VTAIL.n734 VTAIL.n733 8.14595
R878 VTAIL.n725 VTAIL.n696 8.14595
R879 VTAIL.n658 VTAIL.n657 8.14595
R880 VTAIL.n622 VTAIL.n621 8.14595
R881 VTAIL.n613 VTAIL.n584 8.14595
R882 VTAIL.n548 VTAIL.n547 8.14595
R883 VTAIL.n512 VTAIL.n511 8.14595
R884 VTAIL.n503 VTAIL.n474 8.14595
R885 VTAIL.n436 VTAIL.n435 8.14595
R886 VTAIL.n400 VTAIL.n399 8.14595
R887 VTAIL.n391 VTAIL.n362 8.14595
R888 VTAIL.n834 VTAIL.n802 7.3702
R889 VTAIL.n838 VTAIL.n800 7.3702
R890 VTAIL.n883 VTAIL.n780 7.3702
R891 VTAIL.n886 VTAIL.n778 7.3702
R892 VTAIL.n58 VTAIL.n26 7.3702
R893 VTAIL.n62 VTAIL.n24 7.3702
R894 VTAIL.n107 VTAIL.n4 7.3702
R895 VTAIL.n110 VTAIL.n2 7.3702
R896 VTAIL.n168 VTAIL.n136 7.3702
R897 VTAIL.n172 VTAIL.n134 7.3702
R898 VTAIL.n217 VTAIL.n114 7.3702
R899 VTAIL.n220 VTAIL.n112 7.3702
R900 VTAIL.n280 VTAIL.n248 7.3702
R901 VTAIL.n284 VTAIL.n246 7.3702
R902 VTAIL.n329 VTAIL.n226 7.3702
R903 VTAIL.n332 VTAIL.n224 7.3702
R904 VTAIL.n776 VTAIL.n668 7.3702
R905 VTAIL.n773 VTAIL.n670 7.3702
R906 VTAIL.n730 VTAIL.n692 7.3702
R907 VTAIL.n726 VTAIL.n694 7.3702
R908 VTAIL.n664 VTAIL.n556 7.3702
R909 VTAIL.n661 VTAIL.n558 7.3702
R910 VTAIL.n618 VTAIL.n580 7.3702
R911 VTAIL.n614 VTAIL.n582 7.3702
R912 VTAIL.n554 VTAIL.n446 7.3702
R913 VTAIL.n551 VTAIL.n448 7.3702
R914 VTAIL.n508 VTAIL.n470 7.3702
R915 VTAIL.n504 VTAIL.n472 7.3702
R916 VTAIL.n442 VTAIL.n334 7.3702
R917 VTAIL.n439 VTAIL.n336 7.3702
R918 VTAIL.n396 VTAIL.n358 7.3702
R919 VTAIL.n392 VTAIL.n360 7.3702
R920 VTAIL.n837 VTAIL.n802 6.59444
R921 VTAIL.n838 VTAIL.n837 6.59444
R922 VTAIL.n884 VTAIL.n883 6.59444
R923 VTAIL.n884 VTAIL.n778 6.59444
R924 VTAIL.n61 VTAIL.n26 6.59444
R925 VTAIL.n62 VTAIL.n61 6.59444
R926 VTAIL.n108 VTAIL.n107 6.59444
R927 VTAIL.n108 VTAIL.n2 6.59444
R928 VTAIL.n171 VTAIL.n136 6.59444
R929 VTAIL.n172 VTAIL.n171 6.59444
R930 VTAIL.n218 VTAIL.n217 6.59444
R931 VTAIL.n218 VTAIL.n112 6.59444
R932 VTAIL.n283 VTAIL.n248 6.59444
R933 VTAIL.n284 VTAIL.n283 6.59444
R934 VTAIL.n330 VTAIL.n329 6.59444
R935 VTAIL.n330 VTAIL.n224 6.59444
R936 VTAIL.n774 VTAIL.n668 6.59444
R937 VTAIL.n774 VTAIL.n773 6.59444
R938 VTAIL.n730 VTAIL.n729 6.59444
R939 VTAIL.n729 VTAIL.n694 6.59444
R940 VTAIL.n662 VTAIL.n556 6.59444
R941 VTAIL.n662 VTAIL.n661 6.59444
R942 VTAIL.n618 VTAIL.n617 6.59444
R943 VTAIL.n617 VTAIL.n582 6.59444
R944 VTAIL.n552 VTAIL.n446 6.59444
R945 VTAIL.n552 VTAIL.n551 6.59444
R946 VTAIL.n508 VTAIL.n507 6.59444
R947 VTAIL.n507 VTAIL.n472 6.59444
R948 VTAIL.n440 VTAIL.n334 6.59444
R949 VTAIL.n440 VTAIL.n439 6.59444
R950 VTAIL.n396 VTAIL.n395 6.59444
R951 VTAIL.n395 VTAIL.n360 6.59444
R952 VTAIL.n834 VTAIL.n833 5.81868
R953 VTAIL.n841 VTAIL.n800 5.81868
R954 VTAIL.n880 VTAIL.n780 5.81868
R955 VTAIL.n58 VTAIL.n57 5.81868
R956 VTAIL.n65 VTAIL.n24 5.81868
R957 VTAIL.n104 VTAIL.n4 5.81868
R958 VTAIL.n168 VTAIL.n167 5.81868
R959 VTAIL.n175 VTAIL.n134 5.81868
R960 VTAIL.n214 VTAIL.n114 5.81868
R961 VTAIL.n280 VTAIL.n279 5.81868
R962 VTAIL.n287 VTAIL.n246 5.81868
R963 VTAIL.n326 VTAIL.n226 5.81868
R964 VTAIL.n770 VTAIL.n670 5.81868
R965 VTAIL.n733 VTAIL.n692 5.81868
R966 VTAIL.n726 VTAIL.n725 5.81868
R967 VTAIL.n658 VTAIL.n558 5.81868
R968 VTAIL.n621 VTAIL.n580 5.81868
R969 VTAIL.n614 VTAIL.n613 5.81868
R970 VTAIL.n548 VTAIL.n448 5.81868
R971 VTAIL.n511 VTAIL.n470 5.81868
R972 VTAIL.n504 VTAIL.n503 5.81868
R973 VTAIL.n436 VTAIL.n336 5.81868
R974 VTAIL.n399 VTAIL.n358 5.81868
R975 VTAIL.n392 VTAIL.n391 5.81868
R976 VTAIL.n830 VTAIL.n804 5.04292
R977 VTAIL.n842 VTAIL.n798 5.04292
R978 VTAIL.n879 VTAIL.n782 5.04292
R979 VTAIL.n54 VTAIL.n28 5.04292
R980 VTAIL.n66 VTAIL.n22 5.04292
R981 VTAIL.n103 VTAIL.n6 5.04292
R982 VTAIL.n164 VTAIL.n138 5.04292
R983 VTAIL.n176 VTAIL.n132 5.04292
R984 VTAIL.n213 VTAIL.n116 5.04292
R985 VTAIL.n276 VTAIL.n250 5.04292
R986 VTAIL.n288 VTAIL.n244 5.04292
R987 VTAIL.n325 VTAIL.n228 5.04292
R988 VTAIL.n769 VTAIL.n672 5.04292
R989 VTAIL.n734 VTAIL.n690 5.04292
R990 VTAIL.n722 VTAIL.n696 5.04292
R991 VTAIL.n657 VTAIL.n560 5.04292
R992 VTAIL.n622 VTAIL.n578 5.04292
R993 VTAIL.n610 VTAIL.n584 5.04292
R994 VTAIL.n547 VTAIL.n450 5.04292
R995 VTAIL.n512 VTAIL.n468 5.04292
R996 VTAIL.n500 VTAIL.n474 5.04292
R997 VTAIL.n435 VTAIL.n338 5.04292
R998 VTAIL.n400 VTAIL.n356 5.04292
R999 VTAIL.n388 VTAIL.n362 5.04292
R1000 VTAIL.n829 VTAIL.n806 4.26717
R1001 VTAIL.n846 VTAIL.n845 4.26717
R1002 VTAIL.n876 VTAIL.n875 4.26717
R1003 VTAIL.n53 VTAIL.n30 4.26717
R1004 VTAIL.n70 VTAIL.n69 4.26717
R1005 VTAIL.n100 VTAIL.n99 4.26717
R1006 VTAIL.n163 VTAIL.n140 4.26717
R1007 VTAIL.n180 VTAIL.n179 4.26717
R1008 VTAIL.n210 VTAIL.n209 4.26717
R1009 VTAIL.n275 VTAIL.n252 4.26717
R1010 VTAIL.n292 VTAIL.n291 4.26717
R1011 VTAIL.n322 VTAIL.n321 4.26717
R1012 VTAIL.n766 VTAIL.n765 4.26717
R1013 VTAIL.n738 VTAIL.n737 4.26717
R1014 VTAIL.n721 VTAIL.n698 4.26717
R1015 VTAIL.n654 VTAIL.n653 4.26717
R1016 VTAIL.n626 VTAIL.n625 4.26717
R1017 VTAIL.n609 VTAIL.n586 4.26717
R1018 VTAIL.n544 VTAIL.n543 4.26717
R1019 VTAIL.n516 VTAIL.n515 4.26717
R1020 VTAIL.n499 VTAIL.n476 4.26717
R1021 VTAIL.n432 VTAIL.n431 4.26717
R1022 VTAIL.n404 VTAIL.n403 4.26717
R1023 VTAIL.n387 VTAIL.n364 4.26717
R1024 VTAIL.n813 VTAIL.n811 3.70982
R1025 VTAIL.n37 VTAIL.n35 3.70982
R1026 VTAIL.n147 VTAIL.n145 3.70982
R1027 VTAIL.n259 VTAIL.n257 3.70982
R1028 VTAIL.n705 VTAIL.n703 3.70982
R1029 VTAIL.n593 VTAIL.n591 3.70982
R1030 VTAIL.n483 VTAIL.n481 3.70982
R1031 VTAIL.n371 VTAIL.n369 3.70982
R1032 VTAIL.n826 VTAIL.n825 3.49141
R1033 VTAIL.n849 VTAIL.n796 3.49141
R1034 VTAIL.n872 VTAIL.n784 3.49141
R1035 VTAIL.n50 VTAIL.n49 3.49141
R1036 VTAIL.n73 VTAIL.n20 3.49141
R1037 VTAIL.n96 VTAIL.n8 3.49141
R1038 VTAIL.n160 VTAIL.n159 3.49141
R1039 VTAIL.n183 VTAIL.n130 3.49141
R1040 VTAIL.n206 VTAIL.n118 3.49141
R1041 VTAIL.n272 VTAIL.n271 3.49141
R1042 VTAIL.n295 VTAIL.n242 3.49141
R1043 VTAIL.n318 VTAIL.n230 3.49141
R1044 VTAIL.n762 VTAIL.n674 3.49141
R1045 VTAIL.n741 VTAIL.n688 3.49141
R1046 VTAIL.n718 VTAIL.n717 3.49141
R1047 VTAIL.n650 VTAIL.n562 3.49141
R1048 VTAIL.n629 VTAIL.n576 3.49141
R1049 VTAIL.n606 VTAIL.n605 3.49141
R1050 VTAIL.n540 VTAIL.n452 3.49141
R1051 VTAIL.n519 VTAIL.n466 3.49141
R1052 VTAIL.n496 VTAIL.n495 3.49141
R1053 VTAIL.n428 VTAIL.n340 3.49141
R1054 VTAIL.n407 VTAIL.n354 3.49141
R1055 VTAIL.n384 VTAIL.n383 3.49141
R1056 VTAIL.n822 VTAIL.n808 2.71565
R1057 VTAIL.n850 VTAIL.n794 2.71565
R1058 VTAIL.n871 VTAIL.n786 2.71565
R1059 VTAIL.n46 VTAIL.n32 2.71565
R1060 VTAIL.n74 VTAIL.n18 2.71565
R1061 VTAIL.n95 VTAIL.n10 2.71565
R1062 VTAIL.n156 VTAIL.n142 2.71565
R1063 VTAIL.n184 VTAIL.n128 2.71565
R1064 VTAIL.n205 VTAIL.n120 2.71565
R1065 VTAIL.n268 VTAIL.n254 2.71565
R1066 VTAIL.n296 VTAIL.n240 2.71565
R1067 VTAIL.n317 VTAIL.n232 2.71565
R1068 VTAIL.n761 VTAIL.n676 2.71565
R1069 VTAIL.n742 VTAIL.n686 2.71565
R1070 VTAIL.n714 VTAIL.n700 2.71565
R1071 VTAIL.n649 VTAIL.n564 2.71565
R1072 VTAIL.n630 VTAIL.n574 2.71565
R1073 VTAIL.n602 VTAIL.n588 2.71565
R1074 VTAIL.n539 VTAIL.n454 2.71565
R1075 VTAIL.n520 VTAIL.n464 2.71565
R1076 VTAIL.n492 VTAIL.n478 2.71565
R1077 VTAIL.n427 VTAIL.n342 2.71565
R1078 VTAIL.n408 VTAIL.n352 2.71565
R1079 VTAIL.n380 VTAIL.n366 2.71565
R1080 VTAIL.n821 VTAIL.n810 1.93989
R1081 VTAIL.n855 VTAIL.n853 1.93989
R1082 VTAIL.n868 VTAIL.n867 1.93989
R1083 VTAIL.n45 VTAIL.n34 1.93989
R1084 VTAIL.n79 VTAIL.n77 1.93989
R1085 VTAIL.n92 VTAIL.n91 1.93989
R1086 VTAIL.n155 VTAIL.n144 1.93989
R1087 VTAIL.n189 VTAIL.n187 1.93989
R1088 VTAIL.n202 VTAIL.n201 1.93989
R1089 VTAIL.n267 VTAIL.n256 1.93989
R1090 VTAIL.n301 VTAIL.n299 1.93989
R1091 VTAIL.n314 VTAIL.n313 1.93989
R1092 VTAIL.n758 VTAIL.n757 1.93989
R1093 VTAIL.n746 VTAIL.n745 1.93989
R1094 VTAIL.n713 VTAIL.n702 1.93989
R1095 VTAIL.n646 VTAIL.n645 1.93989
R1096 VTAIL.n634 VTAIL.n633 1.93989
R1097 VTAIL.n601 VTAIL.n590 1.93989
R1098 VTAIL.n536 VTAIL.n535 1.93989
R1099 VTAIL.n524 VTAIL.n523 1.93989
R1100 VTAIL.n491 VTAIL.n480 1.93989
R1101 VTAIL.n424 VTAIL.n423 1.93989
R1102 VTAIL.n412 VTAIL.n411 1.93989
R1103 VTAIL.n379 VTAIL.n368 1.93989
R1104 VTAIL.n0 VTAIL.t9 1.65892
R1105 VTAIL.n0 VTAIL.t11 1.65892
R1106 VTAIL.n222 VTAIL.t7 1.65892
R1107 VTAIL.n222 VTAIL.t6 1.65892
R1108 VTAIL.n666 VTAIL.t2 1.65892
R1109 VTAIL.n666 VTAIL.t1 1.65892
R1110 VTAIL.n444 VTAIL.t12 1.65892
R1111 VTAIL.n444 VTAIL.t15 1.65892
R1112 VTAIL.n818 VTAIL.n817 1.16414
R1113 VTAIL.n854 VTAIL.n792 1.16414
R1114 VTAIL.n864 VTAIL.n788 1.16414
R1115 VTAIL.n42 VTAIL.n41 1.16414
R1116 VTAIL.n78 VTAIL.n16 1.16414
R1117 VTAIL.n88 VTAIL.n12 1.16414
R1118 VTAIL.n152 VTAIL.n151 1.16414
R1119 VTAIL.n188 VTAIL.n126 1.16414
R1120 VTAIL.n198 VTAIL.n122 1.16414
R1121 VTAIL.n264 VTAIL.n263 1.16414
R1122 VTAIL.n300 VTAIL.n238 1.16414
R1123 VTAIL.n310 VTAIL.n234 1.16414
R1124 VTAIL.n754 VTAIL.n678 1.16414
R1125 VTAIL.n749 VTAIL.n683 1.16414
R1126 VTAIL.n710 VTAIL.n709 1.16414
R1127 VTAIL.n642 VTAIL.n566 1.16414
R1128 VTAIL.n637 VTAIL.n571 1.16414
R1129 VTAIL.n598 VTAIL.n597 1.16414
R1130 VTAIL.n532 VTAIL.n456 1.16414
R1131 VTAIL.n527 VTAIL.n461 1.16414
R1132 VTAIL.n488 VTAIL.n487 1.16414
R1133 VTAIL.n420 VTAIL.n344 1.16414
R1134 VTAIL.n415 VTAIL.n349 1.16414
R1135 VTAIL.n376 VTAIL.n375 1.16414
R1136 VTAIL.n445 VTAIL.n443 0.483259
R1137 VTAIL.n555 VTAIL.n445 0.483259
R1138 VTAIL.n667 VTAIL.n665 0.483259
R1139 VTAIL.n777 VTAIL.n667 0.483259
R1140 VTAIL.n333 VTAIL.n223 0.483259
R1141 VTAIL.n223 VTAIL.n221 0.483259
R1142 VTAIL.n111 VTAIL.n1 0.483259
R1143 VTAIL.n665 VTAIL.n555 0.470328
R1144 VTAIL.n221 VTAIL.n111 0.470328
R1145 VTAIL VTAIL.n887 0.425069
R1146 VTAIL.n814 VTAIL.n812 0.388379
R1147 VTAIL.n860 VTAIL.n859 0.388379
R1148 VTAIL.n863 VTAIL.n790 0.388379
R1149 VTAIL.n38 VTAIL.n36 0.388379
R1150 VTAIL.n84 VTAIL.n83 0.388379
R1151 VTAIL.n87 VTAIL.n14 0.388379
R1152 VTAIL.n148 VTAIL.n146 0.388379
R1153 VTAIL.n194 VTAIL.n193 0.388379
R1154 VTAIL.n197 VTAIL.n124 0.388379
R1155 VTAIL.n260 VTAIL.n258 0.388379
R1156 VTAIL.n306 VTAIL.n305 0.388379
R1157 VTAIL.n309 VTAIL.n236 0.388379
R1158 VTAIL.n753 VTAIL.n680 0.388379
R1159 VTAIL.n750 VTAIL.n682 0.388379
R1160 VTAIL.n706 VTAIL.n704 0.388379
R1161 VTAIL.n641 VTAIL.n568 0.388379
R1162 VTAIL.n638 VTAIL.n570 0.388379
R1163 VTAIL.n594 VTAIL.n592 0.388379
R1164 VTAIL.n531 VTAIL.n458 0.388379
R1165 VTAIL.n528 VTAIL.n460 0.388379
R1166 VTAIL.n484 VTAIL.n482 0.388379
R1167 VTAIL.n419 VTAIL.n346 0.388379
R1168 VTAIL.n416 VTAIL.n348 0.388379
R1169 VTAIL.n372 VTAIL.n370 0.388379
R1170 VTAIL.n819 VTAIL.n811 0.155672
R1171 VTAIL.n820 VTAIL.n819 0.155672
R1172 VTAIL.n820 VTAIL.n807 0.155672
R1173 VTAIL.n827 VTAIL.n807 0.155672
R1174 VTAIL.n828 VTAIL.n827 0.155672
R1175 VTAIL.n828 VTAIL.n803 0.155672
R1176 VTAIL.n835 VTAIL.n803 0.155672
R1177 VTAIL.n836 VTAIL.n835 0.155672
R1178 VTAIL.n836 VTAIL.n799 0.155672
R1179 VTAIL.n843 VTAIL.n799 0.155672
R1180 VTAIL.n844 VTAIL.n843 0.155672
R1181 VTAIL.n844 VTAIL.n795 0.155672
R1182 VTAIL.n851 VTAIL.n795 0.155672
R1183 VTAIL.n852 VTAIL.n851 0.155672
R1184 VTAIL.n852 VTAIL.n791 0.155672
R1185 VTAIL.n861 VTAIL.n791 0.155672
R1186 VTAIL.n862 VTAIL.n861 0.155672
R1187 VTAIL.n862 VTAIL.n787 0.155672
R1188 VTAIL.n869 VTAIL.n787 0.155672
R1189 VTAIL.n870 VTAIL.n869 0.155672
R1190 VTAIL.n870 VTAIL.n783 0.155672
R1191 VTAIL.n877 VTAIL.n783 0.155672
R1192 VTAIL.n878 VTAIL.n877 0.155672
R1193 VTAIL.n878 VTAIL.n779 0.155672
R1194 VTAIL.n885 VTAIL.n779 0.155672
R1195 VTAIL.n43 VTAIL.n35 0.155672
R1196 VTAIL.n44 VTAIL.n43 0.155672
R1197 VTAIL.n44 VTAIL.n31 0.155672
R1198 VTAIL.n51 VTAIL.n31 0.155672
R1199 VTAIL.n52 VTAIL.n51 0.155672
R1200 VTAIL.n52 VTAIL.n27 0.155672
R1201 VTAIL.n59 VTAIL.n27 0.155672
R1202 VTAIL.n60 VTAIL.n59 0.155672
R1203 VTAIL.n60 VTAIL.n23 0.155672
R1204 VTAIL.n67 VTAIL.n23 0.155672
R1205 VTAIL.n68 VTAIL.n67 0.155672
R1206 VTAIL.n68 VTAIL.n19 0.155672
R1207 VTAIL.n75 VTAIL.n19 0.155672
R1208 VTAIL.n76 VTAIL.n75 0.155672
R1209 VTAIL.n76 VTAIL.n15 0.155672
R1210 VTAIL.n85 VTAIL.n15 0.155672
R1211 VTAIL.n86 VTAIL.n85 0.155672
R1212 VTAIL.n86 VTAIL.n11 0.155672
R1213 VTAIL.n93 VTAIL.n11 0.155672
R1214 VTAIL.n94 VTAIL.n93 0.155672
R1215 VTAIL.n94 VTAIL.n7 0.155672
R1216 VTAIL.n101 VTAIL.n7 0.155672
R1217 VTAIL.n102 VTAIL.n101 0.155672
R1218 VTAIL.n102 VTAIL.n3 0.155672
R1219 VTAIL.n109 VTAIL.n3 0.155672
R1220 VTAIL.n153 VTAIL.n145 0.155672
R1221 VTAIL.n154 VTAIL.n153 0.155672
R1222 VTAIL.n154 VTAIL.n141 0.155672
R1223 VTAIL.n161 VTAIL.n141 0.155672
R1224 VTAIL.n162 VTAIL.n161 0.155672
R1225 VTAIL.n162 VTAIL.n137 0.155672
R1226 VTAIL.n169 VTAIL.n137 0.155672
R1227 VTAIL.n170 VTAIL.n169 0.155672
R1228 VTAIL.n170 VTAIL.n133 0.155672
R1229 VTAIL.n177 VTAIL.n133 0.155672
R1230 VTAIL.n178 VTAIL.n177 0.155672
R1231 VTAIL.n178 VTAIL.n129 0.155672
R1232 VTAIL.n185 VTAIL.n129 0.155672
R1233 VTAIL.n186 VTAIL.n185 0.155672
R1234 VTAIL.n186 VTAIL.n125 0.155672
R1235 VTAIL.n195 VTAIL.n125 0.155672
R1236 VTAIL.n196 VTAIL.n195 0.155672
R1237 VTAIL.n196 VTAIL.n121 0.155672
R1238 VTAIL.n203 VTAIL.n121 0.155672
R1239 VTAIL.n204 VTAIL.n203 0.155672
R1240 VTAIL.n204 VTAIL.n117 0.155672
R1241 VTAIL.n211 VTAIL.n117 0.155672
R1242 VTAIL.n212 VTAIL.n211 0.155672
R1243 VTAIL.n212 VTAIL.n113 0.155672
R1244 VTAIL.n219 VTAIL.n113 0.155672
R1245 VTAIL.n265 VTAIL.n257 0.155672
R1246 VTAIL.n266 VTAIL.n265 0.155672
R1247 VTAIL.n266 VTAIL.n253 0.155672
R1248 VTAIL.n273 VTAIL.n253 0.155672
R1249 VTAIL.n274 VTAIL.n273 0.155672
R1250 VTAIL.n274 VTAIL.n249 0.155672
R1251 VTAIL.n281 VTAIL.n249 0.155672
R1252 VTAIL.n282 VTAIL.n281 0.155672
R1253 VTAIL.n282 VTAIL.n245 0.155672
R1254 VTAIL.n289 VTAIL.n245 0.155672
R1255 VTAIL.n290 VTAIL.n289 0.155672
R1256 VTAIL.n290 VTAIL.n241 0.155672
R1257 VTAIL.n297 VTAIL.n241 0.155672
R1258 VTAIL.n298 VTAIL.n297 0.155672
R1259 VTAIL.n298 VTAIL.n237 0.155672
R1260 VTAIL.n307 VTAIL.n237 0.155672
R1261 VTAIL.n308 VTAIL.n307 0.155672
R1262 VTAIL.n308 VTAIL.n233 0.155672
R1263 VTAIL.n315 VTAIL.n233 0.155672
R1264 VTAIL.n316 VTAIL.n315 0.155672
R1265 VTAIL.n316 VTAIL.n229 0.155672
R1266 VTAIL.n323 VTAIL.n229 0.155672
R1267 VTAIL.n324 VTAIL.n323 0.155672
R1268 VTAIL.n324 VTAIL.n225 0.155672
R1269 VTAIL.n331 VTAIL.n225 0.155672
R1270 VTAIL.n775 VTAIL.n669 0.155672
R1271 VTAIL.n768 VTAIL.n669 0.155672
R1272 VTAIL.n768 VTAIL.n767 0.155672
R1273 VTAIL.n767 VTAIL.n673 0.155672
R1274 VTAIL.n760 VTAIL.n673 0.155672
R1275 VTAIL.n760 VTAIL.n759 0.155672
R1276 VTAIL.n759 VTAIL.n677 0.155672
R1277 VTAIL.n752 VTAIL.n677 0.155672
R1278 VTAIL.n752 VTAIL.n751 0.155672
R1279 VTAIL.n751 VTAIL.n681 0.155672
R1280 VTAIL.n744 VTAIL.n681 0.155672
R1281 VTAIL.n744 VTAIL.n743 0.155672
R1282 VTAIL.n743 VTAIL.n687 0.155672
R1283 VTAIL.n736 VTAIL.n687 0.155672
R1284 VTAIL.n736 VTAIL.n735 0.155672
R1285 VTAIL.n735 VTAIL.n691 0.155672
R1286 VTAIL.n728 VTAIL.n691 0.155672
R1287 VTAIL.n728 VTAIL.n727 0.155672
R1288 VTAIL.n727 VTAIL.n695 0.155672
R1289 VTAIL.n720 VTAIL.n695 0.155672
R1290 VTAIL.n720 VTAIL.n719 0.155672
R1291 VTAIL.n719 VTAIL.n699 0.155672
R1292 VTAIL.n712 VTAIL.n699 0.155672
R1293 VTAIL.n712 VTAIL.n711 0.155672
R1294 VTAIL.n711 VTAIL.n703 0.155672
R1295 VTAIL.n663 VTAIL.n557 0.155672
R1296 VTAIL.n656 VTAIL.n557 0.155672
R1297 VTAIL.n656 VTAIL.n655 0.155672
R1298 VTAIL.n655 VTAIL.n561 0.155672
R1299 VTAIL.n648 VTAIL.n561 0.155672
R1300 VTAIL.n648 VTAIL.n647 0.155672
R1301 VTAIL.n647 VTAIL.n565 0.155672
R1302 VTAIL.n640 VTAIL.n565 0.155672
R1303 VTAIL.n640 VTAIL.n639 0.155672
R1304 VTAIL.n639 VTAIL.n569 0.155672
R1305 VTAIL.n632 VTAIL.n569 0.155672
R1306 VTAIL.n632 VTAIL.n631 0.155672
R1307 VTAIL.n631 VTAIL.n575 0.155672
R1308 VTAIL.n624 VTAIL.n575 0.155672
R1309 VTAIL.n624 VTAIL.n623 0.155672
R1310 VTAIL.n623 VTAIL.n579 0.155672
R1311 VTAIL.n616 VTAIL.n579 0.155672
R1312 VTAIL.n616 VTAIL.n615 0.155672
R1313 VTAIL.n615 VTAIL.n583 0.155672
R1314 VTAIL.n608 VTAIL.n583 0.155672
R1315 VTAIL.n608 VTAIL.n607 0.155672
R1316 VTAIL.n607 VTAIL.n587 0.155672
R1317 VTAIL.n600 VTAIL.n587 0.155672
R1318 VTAIL.n600 VTAIL.n599 0.155672
R1319 VTAIL.n599 VTAIL.n591 0.155672
R1320 VTAIL.n553 VTAIL.n447 0.155672
R1321 VTAIL.n546 VTAIL.n447 0.155672
R1322 VTAIL.n546 VTAIL.n545 0.155672
R1323 VTAIL.n545 VTAIL.n451 0.155672
R1324 VTAIL.n538 VTAIL.n451 0.155672
R1325 VTAIL.n538 VTAIL.n537 0.155672
R1326 VTAIL.n537 VTAIL.n455 0.155672
R1327 VTAIL.n530 VTAIL.n455 0.155672
R1328 VTAIL.n530 VTAIL.n529 0.155672
R1329 VTAIL.n529 VTAIL.n459 0.155672
R1330 VTAIL.n522 VTAIL.n459 0.155672
R1331 VTAIL.n522 VTAIL.n521 0.155672
R1332 VTAIL.n521 VTAIL.n465 0.155672
R1333 VTAIL.n514 VTAIL.n465 0.155672
R1334 VTAIL.n514 VTAIL.n513 0.155672
R1335 VTAIL.n513 VTAIL.n469 0.155672
R1336 VTAIL.n506 VTAIL.n469 0.155672
R1337 VTAIL.n506 VTAIL.n505 0.155672
R1338 VTAIL.n505 VTAIL.n473 0.155672
R1339 VTAIL.n498 VTAIL.n473 0.155672
R1340 VTAIL.n498 VTAIL.n497 0.155672
R1341 VTAIL.n497 VTAIL.n477 0.155672
R1342 VTAIL.n490 VTAIL.n477 0.155672
R1343 VTAIL.n490 VTAIL.n489 0.155672
R1344 VTAIL.n489 VTAIL.n481 0.155672
R1345 VTAIL.n441 VTAIL.n335 0.155672
R1346 VTAIL.n434 VTAIL.n335 0.155672
R1347 VTAIL.n434 VTAIL.n433 0.155672
R1348 VTAIL.n433 VTAIL.n339 0.155672
R1349 VTAIL.n426 VTAIL.n339 0.155672
R1350 VTAIL.n426 VTAIL.n425 0.155672
R1351 VTAIL.n425 VTAIL.n343 0.155672
R1352 VTAIL.n418 VTAIL.n343 0.155672
R1353 VTAIL.n418 VTAIL.n417 0.155672
R1354 VTAIL.n417 VTAIL.n347 0.155672
R1355 VTAIL.n410 VTAIL.n347 0.155672
R1356 VTAIL.n410 VTAIL.n409 0.155672
R1357 VTAIL.n409 VTAIL.n353 0.155672
R1358 VTAIL.n402 VTAIL.n353 0.155672
R1359 VTAIL.n402 VTAIL.n401 0.155672
R1360 VTAIL.n401 VTAIL.n357 0.155672
R1361 VTAIL.n394 VTAIL.n357 0.155672
R1362 VTAIL.n394 VTAIL.n393 0.155672
R1363 VTAIL.n393 VTAIL.n361 0.155672
R1364 VTAIL.n386 VTAIL.n361 0.155672
R1365 VTAIL.n386 VTAIL.n385 0.155672
R1366 VTAIL.n385 VTAIL.n365 0.155672
R1367 VTAIL.n378 VTAIL.n365 0.155672
R1368 VTAIL.n378 VTAIL.n377 0.155672
R1369 VTAIL.n377 VTAIL.n369 0.155672
R1370 VTAIL VTAIL.n1 0.0586897
R1371 VDD2.n2 VDD2.n1 66.7441
R1372 VDD2.n2 VDD2.n0 66.7441
R1373 VDD2 VDD2.n5 66.7413
R1374 VDD2.n4 VDD2.n3 66.5583
R1375 VDD2.n4 VDD2.n2 42.7843
R1376 VDD2.n5 VDD2.t4 1.65892
R1377 VDD2.n5 VDD2.t3 1.65892
R1378 VDD2.n3 VDD2.t2 1.65892
R1379 VDD2.n3 VDD2.t7 1.65892
R1380 VDD2.n1 VDD2.t6 1.65892
R1381 VDD2.n1 VDD2.t5 1.65892
R1382 VDD2.n0 VDD2.t1 1.65892
R1383 VDD2.n0 VDD2.t0 1.65892
R1384 VDD2 VDD2.n4 0.300069
R1385 B.n140 B.t6 2282.23
R1386 B.n132 B.t9 2282.23
R1387 B.n50 B.t0 2282.23
R1388 B.n42 B.t3 2282.23
R1389 B.n409 B.n100 585
R1390 B.n408 B.n407 585
R1391 B.n406 B.n101 585
R1392 B.n405 B.n404 585
R1393 B.n403 B.n102 585
R1394 B.n402 B.n401 585
R1395 B.n400 B.n103 585
R1396 B.n399 B.n398 585
R1397 B.n397 B.n104 585
R1398 B.n396 B.n395 585
R1399 B.n394 B.n105 585
R1400 B.n393 B.n392 585
R1401 B.n391 B.n106 585
R1402 B.n390 B.n389 585
R1403 B.n388 B.n107 585
R1404 B.n387 B.n386 585
R1405 B.n385 B.n108 585
R1406 B.n384 B.n383 585
R1407 B.n382 B.n109 585
R1408 B.n381 B.n380 585
R1409 B.n379 B.n110 585
R1410 B.n378 B.n377 585
R1411 B.n376 B.n111 585
R1412 B.n375 B.n374 585
R1413 B.n373 B.n112 585
R1414 B.n372 B.n371 585
R1415 B.n370 B.n113 585
R1416 B.n369 B.n368 585
R1417 B.n367 B.n114 585
R1418 B.n366 B.n365 585
R1419 B.n364 B.n115 585
R1420 B.n363 B.n362 585
R1421 B.n361 B.n116 585
R1422 B.n360 B.n359 585
R1423 B.n358 B.n117 585
R1424 B.n357 B.n356 585
R1425 B.n355 B.n118 585
R1426 B.n354 B.n353 585
R1427 B.n352 B.n119 585
R1428 B.n351 B.n350 585
R1429 B.n349 B.n120 585
R1430 B.n348 B.n347 585
R1431 B.n346 B.n121 585
R1432 B.n345 B.n344 585
R1433 B.n343 B.n122 585
R1434 B.n342 B.n341 585
R1435 B.n340 B.n123 585
R1436 B.n339 B.n338 585
R1437 B.n337 B.n124 585
R1438 B.n336 B.n335 585
R1439 B.n334 B.n125 585
R1440 B.n333 B.n332 585
R1441 B.n331 B.n126 585
R1442 B.n330 B.n329 585
R1443 B.n328 B.n127 585
R1444 B.n327 B.n326 585
R1445 B.n325 B.n128 585
R1446 B.n324 B.n323 585
R1447 B.n322 B.n129 585
R1448 B.n321 B.n320 585
R1449 B.n319 B.n130 585
R1450 B.n318 B.n317 585
R1451 B.n316 B.n131 585
R1452 B.n315 B.n314 585
R1453 B.n313 B.n312 585
R1454 B.n311 B.n135 585
R1455 B.n310 B.n309 585
R1456 B.n308 B.n136 585
R1457 B.n307 B.n306 585
R1458 B.n305 B.n137 585
R1459 B.n304 B.n303 585
R1460 B.n302 B.n138 585
R1461 B.n301 B.n300 585
R1462 B.n298 B.n139 585
R1463 B.n297 B.n296 585
R1464 B.n295 B.n142 585
R1465 B.n294 B.n293 585
R1466 B.n292 B.n143 585
R1467 B.n291 B.n290 585
R1468 B.n289 B.n144 585
R1469 B.n288 B.n287 585
R1470 B.n286 B.n145 585
R1471 B.n285 B.n284 585
R1472 B.n283 B.n146 585
R1473 B.n282 B.n281 585
R1474 B.n280 B.n147 585
R1475 B.n279 B.n278 585
R1476 B.n277 B.n148 585
R1477 B.n276 B.n275 585
R1478 B.n274 B.n149 585
R1479 B.n273 B.n272 585
R1480 B.n271 B.n150 585
R1481 B.n270 B.n269 585
R1482 B.n268 B.n151 585
R1483 B.n267 B.n266 585
R1484 B.n265 B.n152 585
R1485 B.n264 B.n263 585
R1486 B.n262 B.n153 585
R1487 B.n261 B.n260 585
R1488 B.n259 B.n154 585
R1489 B.n258 B.n257 585
R1490 B.n256 B.n155 585
R1491 B.n255 B.n254 585
R1492 B.n253 B.n156 585
R1493 B.n252 B.n251 585
R1494 B.n250 B.n157 585
R1495 B.n249 B.n248 585
R1496 B.n247 B.n158 585
R1497 B.n246 B.n245 585
R1498 B.n244 B.n159 585
R1499 B.n243 B.n242 585
R1500 B.n241 B.n160 585
R1501 B.n240 B.n239 585
R1502 B.n238 B.n161 585
R1503 B.n237 B.n236 585
R1504 B.n235 B.n162 585
R1505 B.n234 B.n233 585
R1506 B.n232 B.n163 585
R1507 B.n231 B.n230 585
R1508 B.n229 B.n164 585
R1509 B.n228 B.n227 585
R1510 B.n226 B.n165 585
R1511 B.n225 B.n224 585
R1512 B.n223 B.n166 585
R1513 B.n222 B.n221 585
R1514 B.n220 B.n167 585
R1515 B.n219 B.n218 585
R1516 B.n217 B.n168 585
R1517 B.n216 B.n215 585
R1518 B.n214 B.n169 585
R1519 B.n213 B.n212 585
R1520 B.n211 B.n170 585
R1521 B.n210 B.n209 585
R1522 B.n208 B.n171 585
R1523 B.n207 B.n206 585
R1524 B.n205 B.n172 585
R1525 B.n204 B.n203 585
R1526 B.n411 B.n410 585
R1527 B.n412 B.n99 585
R1528 B.n414 B.n413 585
R1529 B.n415 B.n98 585
R1530 B.n417 B.n416 585
R1531 B.n418 B.n97 585
R1532 B.n420 B.n419 585
R1533 B.n421 B.n96 585
R1534 B.n423 B.n422 585
R1535 B.n424 B.n95 585
R1536 B.n426 B.n425 585
R1537 B.n427 B.n94 585
R1538 B.n429 B.n428 585
R1539 B.n430 B.n93 585
R1540 B.n432 B.n431 585
R1541 B.n433 B.n92 585
R1542 B.n435 B.n434 585
R1543 B.n436 B.n91 585
R1544 B.n438 B.n437 585
R1545 B.n439 B.n90 585
R1546 B.n441 B.n440 585
R1547 B.n442 B.n89 585
R1548 B.n444 B.n443 585
R1549 B.n445 B.n88 585
R1550 B.n447 B.n446 585
R1551 B.n448 B.n87 585
R1552 B.n450 B.n449 585
R1553 B.n451 B.n86 585
R1554 B.n453 B.n452 585
R1555 B.n454 B.n85 585
R1556 B.n456 B.n455 585
R1557 B.n457 B.n84 585
R1558 B.n459 B.n458 585
R1559 B.n460 B.n83 585
R1560 B.n667 B.n10 585
R1561 B.n666 B.n665 585
R1562 B.n664 B.n11 585
R1563 B.n663 B.n662 585
R1564 B.n661 B.n12 585
R1565 B.n660 B.n659 585
R1566 B.n658 B.n13 585
R1567 B.n657 B.n656 585
R1568 B.n655 B.n14 585
R1569 B.n654 B.n653 585
R1570 B.n652 B.n15 585
R1571 B.n651 B.n650 585
R1572 B.n649 B.n16 585
R1573 B.n648 B.n647 585
R1574 B.n646 B.n17 585
R1575 B.n645 B.n644 585
R1576 B.n643 B.n18 585
R1577 B.n642 B.n641 585
R1578 B.n640 B.n19 585
R1579 B.n639 B.n638 585
R1580 B.n637 B.n20 585
R1581 B.n636 B.n635 585
R1582 B.n634 B.n21 585
R1583 B.n633 B.n632 585
R1584 B.n631 B.n22 585
R1585 B.n630 B.n629 585
R1586 B.n628 B.n23 585
R1587 B.n627 B.n626 585
R1588 B.n625 B.n24 585
R1589 B.n624 B.n623 585
R1590 B.n622 B.n25 585
R1591 B.n621 B.n620 585
R1592 B.n619 B.n26 585
R1593 B.n618 B.n617 585
R1594 B.n616 B.n27 585
R1595 B.n615 B.n614 585
R1596 B.n613 B.n28 585
R1597 B.n612 B.n611 585
R1598 B.n610 B.n29 585
R1599 B.n609 B.n608 585
R1600 B.n607 B.n30 585
R1601 B.n606 B.n605 585
R1602 B.n604 B.n31 585
R1603 B.n603 B.n602 585
R1604 B.n601 B.n32 585
R1605 B.n600 B.n599 585
R1606 B.n598 B.n33 585
R1607 B.n597 B.n596 585
R1608 B.n595 B.n34 585
R1609 B.n594 B.n593 585
R1610 B.n592 B.n35 585
R1611 B.n591 B.n590 585
R1612 B.n589 B.n36 585
R1613 B.n588 B.n587 585
R1614 B.n586 B.n37 585
R1615 B.n585 B.n584 585
R1616 B.n583 B.n38 585
R1617 B.n582 B.n581 585
R1618 B.n580 B.n39 585
R1619 B.n579 B.n578 585
R1620 B.n577 B.n40 585
R1621 B.n576 B.n575 585
R1622 B.n574 B.n41 585
R1623 B.n573 B.n572 585
R1624 B.n571 B.n570 585
R1625 B.n569 B.n45 585
R1626 B.n568 B.n567 585
R1627 B.n566 B.n46 585
R1628 B.n565 B.n564 585
R1629 B.n563 B.n47 585
R1630 B.n562 B.n561 585
R1631 B.n560 B.n48 585
R1632 B.n559 B.n558 585
R1633 B.n556 B.n49 585
R1634 B.n555 B.n554 585
R1635 B.n553 B.n52 585
R1636 B.n552 B.n551 585
R1637 B.n550 B.n53 585
R1638 B.n549 B.n548 585
R1639 B.n547 B.n54 585
R1640 B.n546 B.n545 585
R1641 B.n544 B.n55 585
R1642 B.n543 B.n542 585
R1643 B.n541 B.n56 585
R1644 B.n540 B.n539 585
R1645 B.n538 B.n57 585
R1646 B.n537 B.n536 585
R1647 B.n535 B.n58 585
R1648 B.n534 B.n533 585
R1649 B.n532 B.n59 585
R1650 B.n531 B.n530 585
R1651 B.n529 B.n60 585
R1652 B.n528 B.n527 585
R1653 B.n526 B.n61 585
R1654 B.n525 B.n524 585
R1655 B.n523 B.n62 585
R1656 B.n522 B.n521 585
R1657 B.n520 B.n63 585
R1658 B.n519 B.n518 585
R1659 B.n517 B.n64 585
R1660 B.n516 B.n515 585
R1661 B.n514 B.n65 585
R1662 B.n513 B.n512 585
R1663 B.n511 B.n66 585
R1664 B.n510 B.n509 585
R1665 B.n508 B.n67 585
R1666 B.n507 B.n506 585
R1667 B.n505 B.n68 585
R1668 B.n504 B.n503 585
R1669 B.n502 B.n69 585
R1670 B.n501 B.n500 585
R1671 B.n499 B.n70 585
R1672 B.n498 B.n497 585
R1673 B.n496 B.n71 585
R1674 B.n495 B.n494 585
R1675 B.n493 B.n72 585
R1676 B.n492 B.n491 585
R1677 B.n490 B.n73 585
R1678 B.n489 B.n488 585
R1679 B.n487 B.n74 585
R1680 B.n486 B.n485 585
R1681 B.n484 B.n75 585
R1682 B.n483 B.n482 585
R1683 B.n481 B.n76 585
R1684 B.n480 B.n479 585
R1685 B.n478 B.n77 585
R1686 B.n477 B.n476 585
R1687 B.n475 B.n78 585
R1688 B.n474 B.n473 585
R1689 B.n472 B.n79 585
R1690 B.n471 B.n470 585
R1691 B.n469 B.n80 585
R1692 B.n468 B.n467 585
R1693 B.n466 B.n81 585
R1694 B.n465 B.n464 585
R1695 B.n463 B.n82 585
R1696 B.n462 B.n461 585
R1697 B.n669 B.n668 585
R1698 B.n670 B.n9 585
R1699 B.n672 B.n671 585
R1700 B.n673 B.n8 585
R1701 B.n675 B.n674 585
R1702 B.n676 B.n7 585
R1703 B.n678 B.n677 585
R1704 B.n679 B.n6 585
R1705 B.n681 B.n680 585
R1706 B.n682 B.n5 585
R1707 B.n684 B.n683 585
R1708 B.n685 B.n4 585
R1709 B.n687 B.n686 585
R1710 B.n688 B.n3 585
R1711 B.n690 B.n689 585
R1712 B.n691 B.n0 585
R1713 B.n2 B.n1 585
R1714 B.n181 B.n180 585
R1715 B.n183 B.n182 585
R1716 B.n184 B.n179 585
R1717 B.n186 B.n185 585
R1718 B.n187 B.n178 585
R1719 B.n189 B.n188 585
R1720 B.n190 B.n177 585
R1721 B.n192 B.n191 585
R1722 B.n193 B.n176 585
R1723 B.n195 B.n194 585
R1724 B.n196 B.n175 585
R1725 B.n198 B.n197 585
R1726 B.n199 B.n174 585
R1727 B.n201 B.n200 585
R1728 B.n202 B.n173 585
R1729 B.n132 B.t10 523.447
R1730 B.n50 B.t2 523.447
R1731 B.n140 B.t7 523.447
R1732 B.n42 B.t5 523.447
R1733 B.n204 B.n173 516.524
R1734 B.n410 B.n409 516.524
R1735 B.n462 B.n83 516.524
R1736 B.n668 B.n667 516.524
R1737 B.n133 B.t11 512.586
R1738 B.n51 B.t1 512.586
R1739 B.n141 B.t8 512.586
R1740 B.n43 B.t4 512.586
R1741 B.n693 B.n692 256.663
R1742 B.n692 B.n691 235.042
R1743 B.n692 B.n2 235.042
R1744 B.n205 B.n204 163.367
R1745 B.n206 B.n205 163.367
R1746 B.n206 B.n171 163.367
R1747 B.n210 B.n171 163.367
R1748 B.n211 B.n210 163.367
R1749 B.n212 B.n211 163.367
R1750 B.n212 B.n169 163.367
R1751 B.n216 B.n169 163.367
R1752 B.n217 B.n216 163.367
R1753 B.n218 B.n217 163.367
R1754 B.n218 B.n167 163.367
R1755 B.n222 B.n167 163.367
R1756 B.n223 B.n222 163.367
R1757 B.n224 B.n223 163.367
R1758 B.n224 B.n165 163.367
R1759 B.n228 B.n165 163.367
R1760 B.n229 B.n228 163.367
R1761 B.n230 B.n229 163.367
R1762 B.n230 B.n163 163.367
R1763 B.n234 B.n163 163.367
R1764 B.n235 B.n234 163.367
R1765 B.n236 B.n235 163.367
R1766 B.n236 B.n161 163.367
R1767 B.n240 B.n161 163.367
R1768 B.n241 B.n240 163.367
R1769 B.n242 B.n241 163.367
R1770 B.n242 B.n159 163.367
R1771 B.n246 B.n159 163.367
R1772 B.n247 B.n246 163.367
R1773 B.n248 B.n247 163.367
R1774 B.n248 B.n157 163.367
R1775 B.n252 B.n157 163.367
R1776 B.n253 B.n252 163.367
R1777 B.n254 B.n253 163.367
R1778 B.n254 B.n155 163.367
R1779 B.n258 B.n155 163.367
R1780 B.n259 B.n258 163.367
R1781 B.n260 B.n259 163.367
R1782 B.n260 B.n153 163.367
R1783 B.n264 B.n153 163.367
R1784 B.n265 B.n264 163.367
R1785 B.n266 B.n265 163.367
R1786 B.n266 B.n151 163.367
R1787 B.n270 B.n151 163.367
R1788 B.n271 B.n270 163.367
R1789 B.n272 B.n271 163.367
R1790 B.n272 B.n149 163.367
R1791 B.n276 B.n149 163.367
R1792 B.n277 B.n276 163.367
R1793 B.n278 B.n277 163.367
R1794 B.n278 B.n147 163.367
R1795 B.n282 B.n147 163.367
R1796 B.n283 B.n282 163.367
R1797 B.n284 B.n283 163.367
R1798 B.n284 B.n145 163.367
R1799 B.n288 B.n145 163.367
R1800 B.n289 B.n288 163.367
R1801 B.n290 B.n289 163.367
R1802 B.n290 B.n143 163.367
R1803 B.n294 B.n143 163.367
R1804 B.n295 B.n294 163.367
R1805 B.n296 B.n295 163.367
R1806 B.n296 B.n139 163.367
R1807 B.n301 B.n139 163.367
R1808 B.n302 B.n301 163.367
R1809 B.n303 B.n302 163.367
R1810 B.n303 B.n137 163.367
R1811 B.n307 B.n137 163.367
R1812 B.n308 B.n307 163.367
R1813 B.n309 B.n308 163.367
R1814 B.n309 B.n135 163.367
R1815 B.n313 B.n135 163.367
R1816 B.n314 B.n313 163.367
R1817 B.n314 B.n131 163.367
R1818 B.n318 B.n131 163.367
R1819 B.n319 B.n318 163.367
R1820 B.n320 B.n319 163.367
R1821 B.n320 B.n129 163.367
R1822 B.n324 B.n129 163.367
R1823 B.n325 B.n324 163.367
R1824 B.n326 B.n325 163.367
R1825 B.n326 B.n127 163.367
R1826 B.n330 B.n127 163.367
R1827 B.n331 B.n330 163.367
R1828 B.n332 B.n331 163.367
R1829 B.n332 B.n125 163.367
R1830 B.n336 B.n125 163.367
R1831 B.n337 B.n336 163.367
R1832 B.n338 B.n337 163.367
R1833 B.n338 B.n123 163.367
R1834 B.n342 B.n123 163.367
R1835 B.n343 B.n342 163.367
R1836 B.n344 B.n343 163.367
R1837 B.n344 B.n121 163.367
R1838 B.n348 B.n121 163.367
R1839 B.n349 B.n348 163.367
R1840 B.n350 B.n349 163.367
R1841 B.n350 B.n119 163.367
R1842 B.n354 B.n119 163.367
R1843 B.n355 B.n354 163.367
R1844 B.n356 B.n355 163.367
R1845 B.n356 B.n117 163.367
R1846 B.n360 B.n117 163.367
R1847 B.n361 B.n360 163.367
R1848 B.n362 B.n361 163.367
R1849 B.n362 B.n115 163.367
R1850 B.n366 B.n115 163.367
R1851 B.n367 B.n366 163.367
R1852 B.n368 B.n367 163.367
R1853 B.n368 B.n113 163.367
R1854 B.n372 B.n113 163.367
R1855 B.n373 B.n372 163.367
R1856 B.n374 B.n373 163.367
R1857 B.n374 B.n111 163.367
R1858 B.n378 B.n111 163.367
R1859 B.n379 B.n378 163.367
R1860 B.n380 B.n379 163.367
R1861 B.n380 B.n109 163.367
R1862 B.n384 B.n109 163.367
R1863 B.n385 B.n384 163.367
R1864 B.n386 B.n385 163.367
R1865 B.n386 B.n107 163.367
R1866 B.n390 B.n107 163.367
R1867 B.n391 B.n390 163.367
R1868 B.n392 B.n391 163.367
R1869 B.n392 B.n105 163.367
R1870 B.n396 B.n105 163.367
R1871 B.n397 B.n396 163.367
R1872 B.n398 B.n397 163.367
R1873 B.n398 B.n103 163.367
R1874 B.n402 B.n103 163.367
R1875 B.n403 B.n402 163.367
R1876 B.n404 B.n403 163.367
R1877 B.n404 B.n101 163.367
R1878 B.n408 B.n101 163.367
R1879 B.n409 B.n408 163.367
R1880 B.n458 B.n83 163.367
R1881 B.n458 B.n457 163.367
R1882 B.n457 B.n456 163.367
R1883 B.n456 B.n85 163.367
R1884 B.n452 B.n85 163.367
R1885 B.n452 B.n451 163.367
R1886 B.n451 B.n450 163.367
R1887 B.n450 B.n87 163.367
R1888 B.n446 B.n87 163.367
R1889 B.n446 B.n445 163.367
R1890 B.n445 B.n444 163.367
R1891 B.n444 B.n89 163.367
R1892 B.n440 B.n89 163.367
R1893 B.n440 B.n439 163.367
R1894 B.n439 B.n438 163.367
R1895 B.n438 B.n91 163.367
R1896 B.n434 B.n91 163.367
R1897 B.n434 B.n433 163.367
R1898 B.n433 B.n432 163.367
R1899 B.n432 B.n93 163.367
R1900 B.n428 B.n93 163.367
R1901 B.n428 B.n427 163.367
R1902 B.n427 B.n426 163.367
R1903 B.n426 B.n95 163.367
R1904 B.n422 B.n95 163.367
R1905 B.n422 B.n421 163.367
R1906 B.n421 B.n420 163.367
R1907 B.n420 B.n97 163.367
R1908 B.n416 B.n97 163.367
R1909 B.n416 B.n415 163.367
R1910 B.n415 B.n414 163.367
R1911 B.n414 B.n99 163.367
R1912 B.n410 B.n99 163.367
R1913 B.n667 B.n666 163.367
R1914 B.n666 B.n11 163.367
R1915 B.n662 B.n11 163.367
R1916 B.n662 B.n661 163.367
R1917 B.n661 B.n660 163.367
R1918 B.n660 B.n13 163.367
R1919 B.n656 B.n13 163.367
R1920 B.n656 B.n655 163.367
R1921 B.n655 B.n654 163.367
R1922 B.n654 B.n15 163.367
R1923 B.n650 B.n15 163.367
R1924 B.n650 B.n649 163.367
R1925 B.n649 B.n648 163.367
R1926 B.n648 B.n17 163.367
R1927 B.n644 B.n17 163.367
R1928 B.n644 B.n643 163.367
R1929 B.n643 B.n642 163.367
R1930 B.n642 B.n19 163.367
R1931 B.n638 B.n19 163.367
R1932 B.n638 B.n637 163.367
R1933 B.n637 B.n636 163.367
R1934 B.n636 B.n21 163.367
R1935 B.n632 B.n21 163.367
R1936 B.n632 B.n631 163.367
R1937 B.n631 B.n630 163.367
R1938 B.n630 B.n23 163.367
R1939 B.n626 B.n23 163.367
R1940 B.n626 B.n625 163.367
R1941 B.n625 B.n624 163.367
R1942 B.n624 B.n25 163.367
R1943 B.n620 B.n25 163.367
R1944 B.n620 B.n619 163.367
R1945 B.n619 B.n618 163.367
R1946 B.n618 B.n27 163.367
R1947 B.n614 B.n27 163.367
R1948 B.n614 B.n613 163.367
R1949 B.n613 B.n612 163.367
R1950 B.n612 B.n29 163.367
R1951 B.n608 B.n29 163.367
R1952 B.n608 B.n607 163.367
R1953 B.n607 B.n606 163.367
R1954 B.n606 B.n31 163.367
R1955 B.n602 B.n31 163.367
R1956 B.n602 B.n601 163.367
R1957 B.n601 B.n600 163.367
R1958 B.n600 B.n33 163.367
R1959 B.n596 B.n33 163.367
R1960 B.n596 B.n595 163.367
R1961 B.n595 B.n594 163.367
R1962 B.n594 B.n35 163.367
R1963 B.n590 B.n35 163.367
R1964 B.n590 B.n589 163.367
R1965 B.n589 B.n588 163.367
R1966 B.n588 B.n37 163.367
R1967 B.n584 B.n37 163.367
R1968 B.n584 B.n583 163.367
R1969 B.n583 B.n582 163.367
R1970 B.n582 B.n39 163.367
R1971 B.n578 B.n39 163.367
R1972 B.n578 B.n577 163.367
R1973 B.n577 B.n576 163.367
R1974 B.n576 B.n41 163.367
R1975 B.n572 B.n41 163.367
R1976 B.n572 B.n571 163.367
R1977 B.n571 B.n45 163.367
R1978 B.n567 B.n45 163.367
R1979 B.n567 B.n566 163.367
R1980 B.n566 B.n565 163.367
R1981 B.n565 B.n47 163.367
R1982 B.n561 B.n47 163.367
R1983 B.n561 B.n560 163.367
R1984 B.n560 B.n559 163.367
R1985 B.n559 B.n49 163.367
R1986 B.n554 B.n49 163.367
R1987 B.n554 B.n553 163.367
R1988 B.n553 B.n552 163.367
R1989 B.n552 B.n53 163.367
R1990 B.n548 B.n53 163.367
R1991 B.n548 B.n547 163.367
R1992 B.n547 B.n546 163.367
R1993 B.n546 B.n55 163.367
R1994 B.n542 B.n55 163.367
R1995 B.n542 B.n541 163.367
R1996 B.n541 B.n540 163.367
R1997 B.n540 B.n57 163.367
R1998 B.n536 B.n57 163.367
R1999 B.n536 B.n535 163.367
R2000 B.n535 B.n534 163.367
R2001 B.n534 B.n59 163.367
R2002 B.n530 B.n59 163.367
R2003 B.n530 B.n529 163.367
R2004 B.n529 B.n528 163.367
R2005 B.n528 B.n61 163.367
R2006 B.n524 B.n61 163.367
R2007 B.n524 B.n523 163.367
R2008 B.n523 B.n522 163.367
R2009 B.n522 B.n63 163.367
R2010 B.n518 B.n63 163.367
R2011 B.n518 B.n517 163.367
R2012 B.n517 B.n516 163.367
R2013 B.n516 B.n65 163.367
R2014 B.n512 B.n65 163.367
R2015 B.n512 B.n511 163.367
R2016 B.n511 B.n510 163.367
R2017 B.n510 B.n67 163.367
R2018 B.n506 B.n67 163.367
R2019 B.n506 B.n505 163.367
R2020 B.n505 B.n504 163.367
R2021 B.n504 B.n69 163.367
R2022 B.n500 B.n69 163.367
R2023 B.n500 B.n499 163.367
R2024 B.n499 B.n498 163.367
R2025 B.n498 B.n71 163.367
R2026 B.n494 B.n71 163.367
R2027 B.n494 B.n493 163.367
R2028 B.n493 B.n492 163.367
R2029 B.n492 B.n73 163.367
R2030 B.n488 B.n73 163.367
R2031 B.n488 B.n487 163.367
R2032 B.n487 B.n486 163.367
R2033 B.n486 B.n75 163.367
R2034 B.n482 B.n75 163.367
R2035 B.n482 B.n481 163.367
R2036 B.n481 B.n480 163.367
R2037 B.n480 B.n77 163.367
R2038 B.n476 B.n77 163.367
R2039 B.n476 B.n475 163.367
R2040 B.n475 B.n474 163.367
R2041 B.n474 B.n79 163.367
R2042 B.n470 B.n79 163.367
R2043 B.n470 B.n469 163.367
R2044 B.n469 B.n468 163.367
R2045 B.n468 B.n81 163.367
R2046 B.n464 B.n81 163.367
R2047 B.n464 B.n463 163.367
R2048 B.n463 B.n462 163.367
R2049 B.n668 B.n9 163.367
R2050 B.n672 B.n9 163.367
R2051 B.n673 B.n672 163.367
R2052 B.n674 B.n673 163.367
R2053 B.n674 B.n7 163.367
R2054 B.n678 B.n7 163.367
R2055 B.n679 B.n678 163.367
R2056 B.n680 B.n679 163.367
R2057 B.n680 B.n5 163.367
R2058 B.n684 B.n5 163.367
R2059 B.n685 B.n684 163.367
R2060 B.n686 B.n685 163.367
R2061 B.n686 B.n3 163.367
R2062 B.n690 B.n3 163.367
R2063 B.n691 B.n690 163.367
R2064 B.n181 B.n2 163.367
R2065 B.n182 B.n181 163.367
R2066 B.n182 B.n179 163.367
R2067 B.n186 B.n179 163.367
R2068 B.n187 B.n186 163.367
R2069 B.n188 B.n187 163.367
R2070 B.n188 B.n177 163.367
R2071 B.n192 B.n177 163.367
R2072 B.n193 B.n192 163.367
R2073 B.n194 B.n193 163.367
R2074 B.n194 B.n175 163.367
R2075 B.n198 B.n175 163.367
R2076 B.n199 B.n198 163.367
R2077 B.n200 B.n199 163.367
R2078 B.n200 B.n173 163.367
R2079 B.n299 B.n141 59.5399
R2080 B.n134 B.n133 59.5399
R2081 B.n557 B.n51 59.5399
R2082 B.n44 B.n43 59.5399
R2083 B.n669 B.n10 33.5615
R2084 B.n461 B.n460 33.5615
R2085 B.n411 B.n100 33.5615
R2086 B.n203 B.n202 33.5615
R2087 B B.n693 18.0485
R2088 B.n141 B.n140 10.8611
R2089 B.n133 B.n132 10.8611
R2090 B.n51 B.n50 10.8611
R2091 B.n43 B.n42 10.8611
R2092 B.n670 B.n669 10.6151
R2093 B.n671 B.n670 10.6151
R2094 B.n671 B.n8 10.6151
R2095 B.n675 B.n8 10.6151
R2096 B.n676 B.n675 10.6151
R2097 B.n677 B.n676 10.6151
R2098 B.n677 B.n6 10.6151
R2099 B.n681 B.n6 10.6151
R2100 B.n682 B.n681 10.6151
R2101 B.n683 B.n682 10.6151
R2102 B.n683 B.n4 10.6151
R2103 B.n687 B.n4 10.6151
R2104 B.n688 B.n687 10.6151
R2105 B.n689 B.n688 10.6151
R2106 B.n689 B.n0 10.6151
R2107 B.n665 B.n10 10.6151
R2108 B.n665 B.n664 10.6151
R2109 B.n664 B.n663 10.6151
R2110 B.n663 B.n12 10.6151
R2111 B.n659 B.n12 10.6151
R2112 B.n659 B.n658 10.6151
R2113 B.n658 B.n657 10.6151
R2114 B.n657 B.n14 10.6151
R2115 B.n653 B.n14 10.6151
R2116 B.n653 B.n652 10.6151
R2117 B.n652 B.n651 10.6151
R2118 B.n651 B.n16 10.6151
R2119 B.n647 B.n16 10.6151
R2120 B.n647 B.n646 10.6151
R2121 B.n646 B.n645 10.6151
R2122 B.n645 B.n18 10.6151
R2123 B.n641 B.n18 10.6151
R2124 B.n641 B.n640 10.6151
R2125 B.n640 B.n639 10.6151
R2126 B.n639 B.n20 10.6151
R2127 B.n635 B.n20 10.6151
R2128 B.n635 B.n634 10.6151
R2129 B.n634 B.n633 10.6151
R2130 B.n633 B.n22 10.6151
R2131 B.n629 B.n22 10.6151
R2132 B.n629 B.n628 10.6151
R2133 B.n628 B.n627 10.6151
R2134 B.n627 B.n24 10.6151
R2135 B.n623 B.n24 10.6151
R2136 B.n623 B.n622 10.6151
R2137 B.n622 B.n621 10.6151
R2138 B.n621 B.n26 10.6151
R2139 B.n617 B.n26 10.6151
R2140 B.n617 B.n616 10.6151
R2141 B.n616 B.n615 10.6151
R2142 B.n615 B.n28 10.6151
R2143 B.n611 B.n28 10.6151
R2144 B.n611 B.n610 10.6151
R2145 B.n610 B.n609 10.6151
R2146 B.n609 B.n30 10.6151
R2147 B.n605 B.n30 10.6151
R2148 B.n605 B.n604 10.6151
R2149 B.n604 B.n603 10.6151
R2150 B.n603 B.n32 10.6151
R2151 B.n599 B.n32 10.6151
R2152 B.n599 B.n598 10.6151
R2153 B.n598 B.n597 10.6151
R2154 B.n597 B.n34 10.6151
R2155 B.n593 B.n34 10.6151
R2156 B.n593 B.n592 10.6151
R2157 B.n592 B.n591 10.6151
R2158 B.n591 B.n36 10.6151
R2159 B.n587 B.n36 10.6151
R2160 B.n587 B.n586 10.6151
R2161 B.n586 B.n585 10.6151
R2162 B.n585 B.n38 10.6151
R2163 B.n581 B.n38 10.6151
R2164 B.n581 B.n580 10.6151
R2165 B.n580 B.n579 10.6151
R2166 B.n579 B.n40 10.6151
R2167 B.n575 B.n40 10.6151
R2168 B.n575 B.n574 10.6151
R2169 B.n574 B.n573 10.6151
R2170 B.n570 B.n569 10.6151
R2171 B.n569 B.n568 10.6151
R2172 B.n568 B.n46 10.6151
R2173 B.n564 B.n46 10.6151
R2174 B.n564 B.n563 10.6151
R2175 B.n563 B.n562 10.6151
R2176 B.n562 B.n48 10.6151
R2177 B.n558 B.n48 10.6151
R2178 B.n556 B.n555 10.6151
R2179 B.n555 B.n52 10.6151
R2180 B.n551 B.n52 10.6151
R2181 B.n551 B.n550 10.6151
R2182 B.n550 B.n549 10.6151
R2183 B.n549 B.n54 10.6151
R2184 B.n545 B.n54 10.6151
R2185 B.n545 B.n544 10.6151
R2186 B.n544 B.n543 10.6151
R2187 B.n543 B.n56 10.6151
R2188 B.n539 B.n56 10.6151
R2189 B.n539 B.n538 10.6151
R2190 B.n538 B.n537 10.6151
R2191 B.n537 B.n58 10.6151
R2192 B.n533 B.n58 10.6151
R2193 B.n533 B.n532 10.6151
R2194 B.n532 B.n531 10.6151
R2195 B.n531 B.n60 10.6151
R2196 B.n527 B.n60 10.6151
R2197 B.n527 B.n526 10.6151
R2198 B.n526 B.n525 10.6151
R2199 B.n525 B.n62 10.6151
R2200 B.n521 B.n62 10.6151
R2201 B.n521 B.n520 10.6151
R2202 B.n520 B.n519 10.6151
R2203 B.n519 B.n64 10.6151
R2204 B.n515 B.n64 10.6151
R2205 B.n515 B.n514 10.6151
R2206 B.n514 B.n513 10.6151
R2207 B.n513 B.n66 10.6151
R2208 B.n509 B.n66 10.6151
R2209 B.n509 B.n508 10.6151
R2210 B.n508 B.n507 10.6151
R2211 B.n507 B.n68 10.6151
R2212 B.n503 B.n68 10.6151
R2213 B.n503 B.n502 10.6151
R2214 B.n502 B.n501 10.6151
R2215 B.n501 B.n70 10.6151
R2216 B.n497 B.n70 10.6151
R2217 B.n497 B.n496 10.6151
R2218 B.n496 B.n495 10.6151
R2219 B.n495 B.n72 10.6151
R2220 B.n491 B.n72 10.6151
R2221 B.n491 B.n490 10.6151
R2222 B.n490 B.n489 10.6151
R2223 B.n489 B.n74 10.6151
R2224 B.n485 B.n74 10.6151
R2225 B.n485 B.n484 10.6151
R2226 B.n484 B.n483 10.6151
R2227 B.n483 B.n76 10.6151
R2228 B.n479 B.n76 10.6151
R2229 B.n479 B.n478 10.6151
R2230 B.n478 B.n477 10.6151
R2231 B.n477 B.n78 10.6151
R2232 B.n473 B.n78 10.6151
R2233 B.n473 B.n472 10.6151
R2234 B.n472 B.n471 10.6151
R2235 B.n471 B.n80 10.6151
R2236 B.n467 B.n80 10.6151
R2237 B.n467 B.n466 10.6151
R2238 B.n466 B.n465 10.6151
R2239 B.n465 B.n82 10.6151
R2240 B.n461 B.n82 10.6151
R2241 B.n460 B.n459 10.6151
R2242 B.n459 B.n84 10.6151
R2243 B.n455 B.n84 10.6151
R2244 B.n455 B.n454 10.6151
R2245 B.n454 B.n453 10.6151
R2246 B.n453 B.n86 10.6151
R2247 B.n449 B.n86 10.6151
R2248 B.n449 B.n448 10.6151
R2249 B.n448 B.n447 10.6151
R2250 B.n447 B.n88 10.6151
R2251 B.n443 B.n88 10.6151
R2252 B.n443 B.n442 10.6151
R2253 B.n442 B.n441 10.6151
R2254 B.n441 B.n90 10.6151
R2255 B.n437 B.n90 10.6151
R2256 B.n437 B.n436 10.6151
R2257 B.n436 B.n435 10.6151
R2258 B.n435 B.n92 10.6151
R2259 B.n431 B.n92 10.6151
R2260 B.n431 B.n430 10.6151
R2261 B.n430 B.n429 10.6151
R2262 B.n429 B.n94 10.6151
R2263 B.n425 B.n94 10.6151
R2264 B.n425 B.n424 10.6151
R2265 B.n424 B.n423 10.6151
R2266 B.n423 B.n96 10.6151
R2267 B.n419 B.n96 10.6151
R2268 B.n419 B.n418 10.6151
R2269 B.n418 B.n417 10.6151
R2270 B.n417 B.n98 10.6151
R2271 B.n413 B.n98 10.6151
R2272 B.n413 B.n412 10.6151
R2273 B.n412 B.n411 10.6151
R2274 B.n180 B.n1 10.6151
R2275 B.n183 B.n180 10.6151
R2276 B.n184 B.n183 10.6151
R2277 B.n185 B.n184 10.6151
R2278 B.n185 B.n178 10.6151
R2279 B.n189 B.n178 10.6151
R2280 B.n190 B.n189 10.6151
R2281 B.n191 B.n190 10.6151
R2282 B.n191 B.n176 10.6151
R2283 B.n195 B.n176 10.6151
R2284 B.n196 B.n195 10.6151
R2285 B.n197 B.n196 10.6151
R2286 B.n197 B.n174 10.6151
R2287 B.n201 B.n174 10.6151
R2288 B.n202 B.n201 10.6151
R2289 B.n203 B.n172 10.6151
R2290 B.n207 B.n172 10.6151
R2291 B.n208 B.n207 10.6151
R2292 B.n209 B.n208 10.6151
R2293 B.n209 B.n170 10.6151
R2294 B.n213 B.n170 10.6151
R2295 B.n214 B.n213 10.6151
R2296 B.n215 B.n214 10.6151
R2297 B.n215 B.n168 10.6151
R2298 B.n219 B.n168 10.6151
R2299 B.n220 B.n219 10.6151
R2300 B.n221 B.n220 10.6151
R2301 B.n221 B.n166 10.6151
R2302 B.n225 B.n166 10.6151
R2303 B.n226 B.n225 10.6151
R2304 B.n227 B.n226 10.6151
R2305 B.n227 B.n164 10.6151
R2306 B.n231 B.n164 10.6151
R2307 B.n232 B.n231 10.6151
R2308 B.n233 B.n232 10.6151
R2309 B.n233 B.n162 10.6151
R2310 B.n237 B.n162 10.6151
R2311 B.n238 B.n237 10.6151
R2312 B.n239 B.n238 10.6151
R2313 B.n239 B.n160 10.6151
R2314 B.n243 B.n160 10.6151
R2315 B.n244 B.n243 10.6151
R2316 B.n245 B.n244 10.6151
R2317 B.n245 B.n158 10.6151
R2318 B.n249 B.n158 10.6151
R2319 B.n250 B.n249 10.6151
R2320 B.n251 B.n250 10.6151
R2321 B.n251 B.n156 10.6151
R2322 B.n255 B.n156 10.6151
R2323 B.n256 B.n255 10.6151
R2324 B.n257 B.n256 10.6151
R2325 B.n257 B.n154 10.6151
R2326 B.n261 B.n154 10.6151
R2327 B.n262 B.n261 10.6151
R2328 B.n263 B.n262 10.6151
R2329 B.n263 B.n152 10.6151
R2330 B.n267 B.n152 10.6151
R2331 B.n268 B.n267 10.6151
R2332 B.n269 B.n268 10.6151
R2333 B.n269 B.n150 10.6151
R2334 B.n273 B.n150 10.6151
R2335 B.n274 B.n273 10.6151
R2336 B.n275 B.n274 10.6151
R2337 B.n275 B.n148 10.6151
R2338 B.n279 B.n148 10.6151
R2339 B.n280 B.n279 10.6151
R2340 B.n281 B.n280 10.6151
R2341 B.n281 B.n146 10.6151
R2342 B.n285 B.n146 10.6151
R2343 B.n286 B.n285 10.6151
R2344 B.n287 B.n286 10.6151
R2345 B.n287 B.n144 10.6151
R2346 B.n291 B.n144 10.6151
R2347 B.n292 B.n291 10.6151
R2348 B.n293 B.n292 10.6151
R2349 B.n293 B.n142 10.6151
R2350 B.n297 B.n142 10.6151
R2351 B.n298 B.n297 10.6151
R2352 B.n300 B.n138 10.6151
R2353 B.n304 B.n138 10.6151
R2354 B.n305 B.n304 10.6151
R2355 B.n306 B.n305 10.6151
R2356 B.n306 B.n136 10.6151
R2357 B.n310 B.n136 10.6151
R2358 B.n311 B.n310 10.6151
R2359 B.n312 B.n311 10.6151
R2360 B.n316 B.n315 10.6151
R2361 B.n317 B.n316 10.6151
R2362 B.n317 B.n130 10.6151
R2363 B.n321 B.n130 10.6151
R2364 B.n322 B.n321 10.6151
R2365 B.n323 B.n322 10.6151
R2366 B.n323 B.n128 10.6151
R2367 B.n327 B.n128 10.6151
R2368 B.n328 B.n327 10.6151
R2369 B.n329 B.n328 10.6151
R2370 B.n329 B.n126 10.6151
R2371 B.n333 B.n126 10.6151
R2372 B.n334 B.n333 10.6151
R2373 B.n335 B.n334 10.6151
R2374 B.n335 B.n124 10.6151
R2375 B.n339 B.n124 10.6151
R2376 B.n340 B.n339 10.6151
R2377 B.n341 B.n340 10.6151
R2378 B.n341 B.n122 10.6151
R2379 B.n345 B.n122 10.6151
R2380 B.n346 B.n345 10.6151
R2381 B.n347 B.n346 10.6151
R2382 B.n347 B.n120 10.6151
R2383 B.n351 B.n120 10.6151
R2384 B.n352 B.n351 10.6151
R2385 B.n353 B.n352 10.6151
R2386 B.n353 B.n118 10.6151
R2387 B.n357 B.n118 10.6151
R2388 B.n358 B.n357 10.6151
R2389 B.n359 B.n358 10.6151
R2390 B.n359 B.n116 10.6151
R2391 B.n363 B.n116 10.6151
R2392 B.n364 B.n363 10.6151
R2393 B.n365 B.n364 10.6151
R2394 B.n365 B.n114 10.6151
R2395 B.n369 B.n114 10.6151
R2396 B.n370 B.n369 10.6151
R2397 B.n371 B.n370 10.6151
R2398 B.n371 B.n112 10.6151
R2399 B.n375 B.n112 10.6151
R2400 B.n376 B.n375 10.6151
R2401 B.n377 B.n376 10.6151
R2402 B.n377 B.n110 10.6151
R2403 B.n381 B.n110 10.6151
R2404 B.n382 B.n381 10.6151
R2405 B.n383 B.n382 10.6151
R2406 B.n383 B.n108 10.6151
R2407 B.n387 B.n108 10.6151
R2408 B.n388 B.n387 10.6151
R2409 B.n389 B.n388 10.6151
R2410 B.n389 B.n106 10.6151
R2411 B.n393 B.n106 10.6151
R2412 B.n394 B.n393 10.6151
R2413 B.n395 B.n394 10.6151
R2414 B.n395 B.n104 10.6151
R2415 B.n399 B.n104 10.6151
R2416 B.n400 B.n399 10.6151
R2417 B.n401 B.n400 10.6151
R2418 B.n401 B.n102 10.6151
R2419 B.n405 B.n102 10.6151
R2420 B.n406 B.n405 10.6151
R2421 B.n407 B.n406 10.6151
R2422 B.n407 B.n100 10.6151
R2423 B.n693 B.n0 8.11757
R2424 B.n693 B.n1 8.11757
R2425 B.n570 B.n44 6.5566
R2426 B.n558 B.n557 6.5566
R2427 B.n300 B.n299 6.5566
R2428 B.n312 B.n134 6.5566
R2429 B.n573 B.n44 4.05904
R2430 B.n557 B.n556 4.05904
R2431 B.n299 B.n298 4.05904
R2432 B.n315 B.n134 4.05904
R2433 VP.n13 VP.t2 2241.71
R2434 VP.n9 VP.t6 2241.71
R2435 VP.n2 VP.t3 2241.71
R2436 VP.n6 VP.t7 2241.71
R2437 VP.n12 VP.t4 2192.05
R2438 VP.n10 VP.t5 2192.05
R2439 VP.n3 VP.t0 2192.05
R2440 VP.n5 VP.t1 2192.05
R2441 VP.n2 VP.n1 161.489
R2442 VP.n14 VP.n13 161.3
R2443 VP.n4 VP.n1 161.3
R2444 VP.n7 VP.n6 161.3
R2445 VP.n11 VP.n0 161.3
R2446 VP.n9 VP.n8 161.3
R2447 VP.n8 VP.n7 45.6596
R2448 VP.n11 VP.n10 40.8975
R2449 VP.n12 VP.n11 40.8975
R2450 VP.n4 VP.n3 40.8975
R2451 VP.n5 VP.n4 40.8975
R2452 VP.n10 VP.n9 32.1338
R2453 VP.n13 VP.n12 32.1338
R2454 VP.n3 VP.n2 32.1338
R2455 VP.n6 VP.n5 32.1338
R2456 VP.n7 VP.n1 0.189894
R2457 VP.n8 VP.n0 0.189894
R2458 VP.n14 VP.n0 0.189894
R2459 VP VP.n14 0.0516364
R2460 VDD1 VDD1.n0 66.8578
R2461 VDD1.n3 VDD1.n2 66.7441
R2462 VDD1.n3 VDD1.n1 66.7441
R2463 VDD1.n5 VDD1.n4 66.5581
R2464 VDD1.n5 VDD1.n3 43.3673
R2465 VDD1.n4 VDD1.t6 1.65892
R2466 VDD1.n4 VDD1.t0 1.65892
R2467 VDD1.n0 VDD1.t4 1.65892
R2468 VDD1.n0 VDD1.t7 1.65892
R2469 VDD1.n2 VDD1.t3 1.65892
R2470 VDD1.n2 VDD1.t5 1.65892
R2471 VDD1.n1 VDD1.t1 1.65892
R2472 VDD1.n1 VDD1.t2 1.65892
R2473 VDD1 VDD1.n5 0.18369
C0 VTAIL VN 3.62302f
C1 w_n1530_n4888# VP 2.78944f
C2 VDD1 w_n1530_n4888# 1.30386f
C3 VP VN 6.17279f
C4 VDD1 VN 0.14675f
C5 w_n1530_n4888# VDD2 1.31957f
C6 VTAIL VP 3.63712f
C7 w_n1530_n4888# B 8.66623f
C8 VTAIL VDD1 28.9961f
C9 VDD2 VN 4.41966f
C10 B VN 0.75614f
C11 VTAIL VDD2 29.0346f
C12 VTAIL B 5.28948f
C13 VDD1 VP 4.5395f
C14 VDD2 VP 0.266784f
C15 VDD1 VDD2 0.597203f
C16 B VP 1.06476f
C17 VDD1 B 1.13113f
C18 B VDD2 1.15366f
C19 w_n1530_n4888# VN 2.5978f
C20 VTAIL w_n1530_n4888# 6.28954f
C21 VDD2 VSUBS 1.659694f
C22 VDD1 VSUBS 1.869053f
C23 VTAIL VSUBS 0.869895f
C24 VN VSUBS 5.34001f
C25 VP VSUBS 1.460068f
C26 B VSUBS 2.990289f
C27 w_n1530_n4888# VSUBS 91.340996f
C28 VDD1.t4 VSUBS 0.57022f
C29 VDD1.t7 VSUBS 0.57022f
C30 VDD1.n0 VSUBS 4.77567f
C31 VDD1.t1 VSUBS 0.57022f
C32 VDD1.t2 VSUBS 0.57022f
C33 VDD1.n1 VSUBS 4.77417f
C34 VDD1.t3 VSUBS 0.57022f
C35 VDD1.t5 VSUBS 0.57022f
C36 VDD1.n2 VSUBS 4.77417f
C37 VDD1.n3 VSUBS 4.45353f
C38 VDD1.t6 VSUBS 0.57022f
C39 VDD1.t0 VSUBS 0.57022f
C40 VDD1.n4 VSUBS 4.77181f
C41 VDD1.n5 VSUBS 4.48024f
C42 VP.n0 VSUBS 0.070586f
C43 VP.t4 VSUBS 0.896609f
C44 VP.t5 VSUBS 0.896609f
C45 VP.t6 VSUBS 0.904187f
C46 VP.n1 VSUBS 0.158912f
C47 VP.t1 VSUBS 0.896609f
C48 VP.t0 VSUBS 0.896609f
C49 VP.t3 VSUBS 0.904187f
C50 VP.n2 VSUBS 0.36063f
C51 VP.n3 VSUBS 0.339031f
C52 VP.n4 VSUBS 0.026027f
C53 VP.n5 VSUBS 0.339031f
C54 VP.t7 VSUBS 0.904187f
C55 VP.n6 VSUBS 0.360526f
C56 VP.n7 VSUBS 3.33655f
C57 VP.n8 VSUBS 3.39196f
C58 VP.n9 VSUBS 0.360526f
C59 VP.n10 VSUBS 0.339031f
C60 VP.n11 VSUBS 0.026027f
C61 VP.n12 VSUBS 0.339031f
C62 VP.t2 VSUBS 0.904187f
C63 VP.n13 VSUBS 0.360526f
C64 VP.n14 VSUBS 0.054702f
C65 B.n0 VSUBS 0.007369f
C66 B.n1 VSUBS 0.007369f
C67 B.n2 VSUBS 0.010898f
C68 B.n3 VSUBS 0.008351f
C69 B.n4 VSUBS 0.008351f
C70 B.n5 VSUBS 0.008351f
C71 B.n6 VSUBS 0.008351f
C72 B.n7 VSUBS 0.008351f
C73 B.n8 VSUBS 0.008351f
C74 B.n9 VSUBS 0.008351f
C75 B.n10 VSUBS 0.020024f
C76 B.n11 VSUBS 0.008351f
C77 B.n12 VSUBS 0.008351f
C78 B.n13 VSUBS 0.008351f
C79 B.n14 VSUBS 0.008351f
C80 B.n15 VSUBS 0.008351f
C81 B.n16 VSUBS 0.008351f
C82 B.n17 VSUBS 0.008351f
C83 B.n18 VSUBS 0.008351f
C84 B.n19 VSUBS 0.008351f
C85 B.n20 VSUBS 0.008351f
C86 B.n21 VSUBS 0.008351f
C87 B.n22 VSUBS 0.008351f
C88 B.n23 VSUBS 0.008351f
C89 B.n24 VSUBS 0.008351f
C90 B.n25 VSUBS 0.008351f
C91 B.n26 VSUBS 0.008351f
C92 B.n27 VSUBS 0.008351f
C93 B.n28 VSUBS 0.008351f
C94 B.n29 VSUBS 0.008351f
C95 B.n30 VSUBS 0.008351f
C96 B.n31 VSUBS 0.008351f
C97 B.n32 VSUBS 0.008351f
C98 B.n33 VSUBS 0.008351f
C99 B.n34 VSUBS 0.008351f
C100 B.n35 VSUBS 0.008351f
C101 B.n36 VSUBS 0.008351f
C102 B.n37 VSUBS 0.008351f
C103 B.n38 VSUBS 0.008351f
C104 B.n39 VSUBS 0.008351f
C105 B.n40 VSUBS 0.008351f
C106 B.n41 VSUBS 0.008351f
C107 B.t4 VSUBS 0.465406f
C108 B.t5 VSUBS 0.473518f
C109 B.t3 VSUBS 0.206623f
C110 B.n42 VSUBS 0.458387f
C111 B.n43 VSUBS 0.402907f
C112 B.n44 VSUBS 0.019349f
C113 B.n45 VSUBS 0.008351f
C114 B.n46 VSUBS 0.008351f
C115 B.n47 VSUBS 0.008351f
C116 B.n48 VSUBS 0.008351f
C117 B.n49 VSUBS 0.008351f
C118 B.t1 VSUBS 0.46541f
C119 B.t2 VSUBS 0.473523f
C120 B.t0 VSUBS 0.206623f
C121 B.n50 VSUBS 0.458383f
C122 B.n51 VSUBS 0.402902f
C123 B.n52 VSUBS 0.008351f
C124 B.n53 VSUBS 0.008351f
C125 B.n54 VSUBS 0.008351f
C126 B.n55 VSUBS 0.008351f
C127 B.n56 VSUBS 0.008351f
C128 B.n57 VSUBS 0.008351f
C129 B.n58 VSUBS 0.008351f
C130 B.n59 VSUBS 0.008351f
C131 B.n60 VSUBS 0.008351f
C132 B.n61 VSUBS 0.008351f
C133 B.n62 VSUBS 0.008351f
C134 B.n63 VSUBS 0.008351f
C135 B.n64 VSUBS 0.008351f
C136 B.n65 VSUBS 0.008351f
C137 B.n66 VSUBS 0.008351f
C138 B.n67 VSUBS 0.008351f
C139 B.n68 VSUBS 0.008351f
C140 B.n69 VSUBS 0.008351f
C141 B.n70 VSUBS 0.008351f
C142 B.n71 VSUBS 0.008351f
C143 B.n72 VSUBS 0.008351f
C144 B.n73 VSUBS 0.008351f
C145 B.n74 VSUBS 0.008351f
C146 B.n75 VSUBS 0.008351f
C147 B.n76 VSUBS 0.008351f
C148 B.n77 VSUBS 0.008351f
C149 B.n78 VSUBS 0.008351f
C150 B.n79 VSUBS 0.008351f
C151 B.n80 VSUBS 0.008351f
C152 B.n81 VSUBS 0.008351f
C153 B.n82 VSUBS 0.008351f
C154 B.n83 VSUBS 0.019767f
C155 B.n84 VSUBS 0.008351f
C156 B.n85 VSUBS 0.008351f
C157 B.n86 VSUBS 0.008351f
C158 B.n87 VSUBS 0.008351f
C159 B.n88 VSUBS 0.008351f
C160 B.n89 VSUBS 0.008351f
C161 B.n90 VSUBS 0.008351f
C162 B.n91 VSUBS 0.008351f
C163 B.n92 VSUBS 0.008351f
C164 B.n93 VSUBS 0.008351f
C165 B.n94 VSUBS 0.008351f
C166 B.n95 VSUBS 0.008351f
C167 B.n96 VSUBS 0.008351f
C168 B.n97 VSUBS 0.008351f
C169 B.n98 VSUBS 0.008351f
C170 B.n99 VSUBS 0.008351f
C171 B.n100 VSUBS 0.019064f
C172 B.n101 VSUBS 0.008351f
C173 B.n102 VSUBS 0.008351f
C174 B.n103 VSUBS 0.008351f
C175 B.n104 VSUBS 0.008351f
C176 B.n105 VSUBS 0.008351f
C177 B.n106 VSUBS 0.008351f
C178 B.n107 VSUBS 0.008351f
C179 B.n108 VSUBS 0.008351f
C180 B.n109 VSUBS 0.008351f
C181 B.n110 VSUBS 0.008351f
C182 B.n111 VSUBS 0.008351f
C183 B.n112 VSUBS 0.008351f
C184 B.n113 VSUBS 0.008351f
C185 B.n114 VSUBS 0.008351f
C186 B.n115 VSUBS 0.008351f
C187 B.n116 VSUBS 0.008351f
C188 B.n117 VSUBS 0.008351f
C189 B.n118 VSUBS 0.008351f
C190 B.n119 VSUBS 0.008351f
C191 B.n120 VSUBS 0.008351f
C192 B.n121 VSUBS 0.008351f
C193 B.n122 VSUBS 0.008351f
C194 B.n123 VSUBS 0.008351f
C195 B.n124 VSUBS 0.008351f
C196 B.n125 VSUBS 0.008351f
C197 B.n126 VSUBS 0.008351f
C198 B.n127 VSUBS 0.008351f
C199 B.n128 VSUBS 0.008351f
C200 B.n129 VSUBS 0.008351f
C201 B.n130 VSUBS 0.008351f
C202 B.n131 VSUBS 0.008351f
C203 B.t11 VSUBS 0.46541f
C204 B.t10 VSUBS 0.473523f
C205 B.t9 VSUBS 0.206623f
C206 B.n132 VSUBS 0.458383f
C207 B.n133 VSUBS 0.402902f
C208 B.n134 VSUBS 0.019349f
C209 B.n135 VSUBS 0.008351f
C210 B.n136 VSUBS 0.008351f
C211 B.n137 VSUBS 0.008351f
C212 B.n138 VSUBS 0.008351f
C213 B.n139 VSUBS 0.008351f
C214 B.t8 VSUBS 0.465406f
C215 B.t7 VSUBS 0.473518f
C216 B.t6 VSUBS 0.206623f
C217 B.n140 VSUBS 0.458387f
C218 B.n141 VSUBS 0.402907f
C219 B.n142 VSUBS 0.008351f
C220 B.n143 VSUBS 0.008351f
C221 B.n144 VSUBS 0.008351f
C222 B.n145 VSUBS 0.008351f
C223 B.n146 VSUBS 0.008351f
C224 B.n147 VSUBS 0.008351f
C225 B.n148 VSUBS 0.008351f
C226 B.n149 VSUBS 0.008351f
C227 B.n150 VSUBS 0.008351f
C228 B.n151 VSUBS 0.008351f
C229 B.n152 VSUBS 0.008351f
C230 B.n153 VSUBS 0.008351f
C231 B.n154 VSUBS 0.008351f
C232 B.n155 VSUBS 0.008351f
C233 B.n156 VSUBS 0.008351f
C234 B.n157 VSUBS 0.008351f
C235 B.n158 VSUBS 0.008351f
C236 B.n159 VSUBS 0.008351f
C237 B.n160 VSUBS 0.008351f
C238 B.n161 VSUBS 0.008351f
C239 B.n162 VSUBS 0.008351f
C240 B.n163 VSUBS 0.008351f
C241 B.n164 VSUBS 0.008351f
C242 B.n165 VSUBS 0.008351f
C243 B.n166 VSUBS 0.008351f
C244 B.n167 VSUBS 0.008351f
C245 B.n168 VSUBS 0.008351f
C246 B.n169 VSUBS 0.008351f
C247 B.n170 VSUBS 0.008351f
C248 B.n171 VSUBS 0.008351f
C249 B.n172 VSUBS 0.008351f
C250 B.n173 VSUBS 0.019767f
C251 B.n174 VSUBS 0.008351f
C252 B.n175 VSUBS 0.008351f
C253 B.n176 VSUBS 0.008351f
C254 B.n177 VSUBS 0.008351f
C255 B.n178 VSUBS 0.008351f
C256 B.n179 VSUBS 0.008351f
C257 B.n180 VSUBS 0.008351f
C258 B.n181 VSUBS 0.008351f
C259 B.n182 VSUBS 0.008351f
C260 B.n183 VSUBS 0.008351f
C261 B.n184 VSUBS 0.008351f
C262 B.n185 VSUBS 0.008351f
C263 B.n186 VSUBS 0.008351f
C264 B.n187 VSUBS 0.008351f
C265 B.n188 VSUBS 0.008351f
C266 B.n189 VSUBS 0.008351f
C267 B.n190 VSUBS 0.008351f
C268 B.n191 VSUBS 0.008351f
C269 B.n192 VSUBS 0.008351f
C270 B.n193 VSUBS 0.008351f
C271 B.n194 VSUBS 0.008351f
C272 B.n195 VSUBS 0.008351f
C273 B.n196 VSUBS 0.008351f
C274 B.n197 VSUBS 0.008351f
C275 B.n198 VSUBS 0.008351f
C276 B.n199 VSUBS 0.008351f
C277 B.n200 VSUBS 0.008351f
C278 B.n201 VSUBS 0.008351f
C279 B.n202 VSUBS 0.019767f
C280 B.n203 VSUBS 0.020024f
C281 B.n204 VSUBS 0.020024f
C282 B.n205 VSUBS 0.008351f
C283 B.n206 VSUBS 0.008351f
C284 B.n207 VSUBS 0.008351f
C285 B.n208 VSUBS 0.008351f
C286 B.n209 VSUBS 0.008351f
C287 B.n210 VSUBS 0.008351f
C288 B.n211 VSUBS 0.008351f
C289 B.n212 VSUBS 0.008351f
C290 B.n213 VSUBS 0.008351f
C291 B.n214 VSUBS 0.008351f
C292 B.n215 VSUBS 0.008351f
C293 B.n216 VSUBS 0.008351f
C294 B.n217 VSUBS 0.008351f
C295 B.n218 VSUBS 0.008351f
C296 B.n219 VSUBS 0.008351f
C297 B.n220 VSUBS 0.008351f
C298 B.n221 VSUBS 0.008351f
C299 B.n222 VSUBS 0.008351f
C300 B.n223 VSUBS 0.008351f
C301 B.n224 VSUBS 0.008351f
C302 B.n225 VSUBS 0.008351f
C303 B.n226 VSUBS 0.008351f
C304 B.n227 VSUBS 0.008351f
C305 B.n228 VSUBS 0.008351f
C306 B.n229 VSUBS 0.008351f
C307 B.n230 VSUBS 0.008351f
C308 B.n231 VSUBS 0.008351f
C309 B.n232 VSUBS 0.008351f
C310 B.n233 VSUBS 0.008351f
C311 B.n234 VSUBS 0.008351f
C312 B.n235 VSUBS 0.008351f
C313 B.n236 VSUBS 0.008351f
C314 B.n237 VSUBS 0.008351f
C315 B.n238 VSUBS 0.008351f
C316 B.n239 VSUBS 0.008351f
C317 B.n240 VSUBS 0.008351f
C318 B.n241 VSUBS 0.008351f
C319 B.n242 VSUBS 0.008351f
C320 B.n243 VSUBS 0.008351f
C321 B.n244 VSUBS 0.008351f
C322 B.n245 VSUBS 0.008351f
C323 B.n246 VSUBS 0.008351f
C324 B.n247 VSUBS 0.008351f
C325 B.n248 VSUBS 0.008351f
C326 B.n249 VSUBS 0.008351f
C327 B.n250 VSUBS 0.008351f
C328 B.n251 VSUBS 0.008351f
C329 B.n252 VSUBS 0.008351f
C330 B.n253 VSUBS 0.008351f
C331 B.n254 VSUBS 0.008351f
C332 B.n255 VSUBS 0.008351f
C333 B.n256 VSUBS 0.008351f
C334 B.n257 VSUBS 0.008351f
C335 B.n258 VSUBS 0.008351f
C336 B.n259 VSUBS 0.008351f
C337 B.n260 VSUBS 0.008351f
C338 B.n261 VSUBS 0.008351f
C339 B.n262 VSUBS 0.008351f
C340 B.n263 VSUBS 0.008351f
C341 B.n264 VSUBS 0.008351f
C342 B.n265 VSUBS 0.008351f
C343 B.n266 VSUBS 0.008351f
C344 B.n267 VSUBS 0.008351f
C345 B.n268 VSUBS 0.008351f
C346 B.n269 VSUBS 0.008351f
C347 B.n270 VSUBS 0.008351f
C348 B.n271 VSUBS 0.008351f
C349 B.n272 VSUBS 0.008351f
C350 B.n273 VSUBS 0.008351f
C351 B.n274 VSUBS 0.008351f
C352 B.n275 VSUBS 0.008351f
C353 B.n276 VSUBS 0.008351f
C354 B.n277 VSUBS 0.008351f
C355 B.n278 VSUBS 0.008351f
C356 B.n279 VSUBS 0.008351f
C357 B.n280 VSUBS 0.008351f
C358 B.n281 VSUBS 0.008351f
C359 B.n282 VSUBS 0.008351f
C360 B.n283 VSUBS 0.008351f
C361 B.n284 VSUBS 0.008351f
C362 B.n285 VSUBS 0.008351f
C363 B.n286 VSUBS 0.008351f
C364 B.n287 VSUBS 0.008351f
C365 B.n288 VSUBS 0.008351f
C366 B.n289 VSUBS 0.008351f
C367 B.n290 VSUBS 0.008351f
C368 B.n291 VSUBS 0.008351f
C369 B.n292 VSUBS 0.008351f
C370 B.n293 VSUBS 0.008351f
C371 B.n294 VSUBS 0.008351f
C372 B.n295 VSUBS 0.008351f
C373 B.n296 VSUBS 0.008351f
C374 B.n297 VSUBS 0.008351f
C375 B.n298 VSUBS 0.005772f
C376 B.n299 VSUBS 0.019349f
C377 B.n300 VSUBS 0.006755f
C378 B.n301 VSUBS 0.008351f
C379 B.n302 VSUBS 0.008351f
C380 B.n303 VSUBS 0.008351f
C381 B.n304 VSUBS 0.008351f
C382 B.n305 VSUBS 0.008351f
C383 B.n306 VSUBS 0.008351f
C384 B.n307 VSUBS 0.008351f
C385 B.n308 VSUBS 0.008351f
C386 B.n309 VSUBS 0.008351f
C387 B.n310 VSUBS 0.008351f
C388 B.n311 VSUBS 0.008351f
C389 B.n312 VSUBS 0.006755f
C390 B.n313 VSUBS 0.008351f
C391 B.n314 VSUBS 0.008351f
C392 B.n315 VSUBS 0.005772f
C393 B.n316 VSUBS 0.008351f
C394 B.n317 VSUBS 0.008351f
C395 B.n318 VSUBS 0.008351f
C396 B.n319 VSUBS 0.008351f
C397 B.n320 VSUBS 0.008351f
C398 B.n321 VSUBS 0.008351f
C399 B.n322 VSUBS 0.008351f
C400 B.n323 VSUBS 0.008351f
C401 B.n324 VSUBS 0.008351f
C402 B.n325 VSUBS 0.008351f
C403 B.n326 VSUBS 0.008351f
C404 B.n327 VSUBS 0.008351f
C405 B.n328 VSUBS 0.008351f
C406 B.n329 VSUBS 0.008351f
C407 B.n330 VSUBS 0.008351f
C408 B.n331 VSUBS 0.008351f
C409 B.n332 VSUBS 0.008351f
C410 B.n333 VSUBS 0.008351f
C411 B.n334 VSUBS 0.008351f
C412 B.n335 VSUBS 0.008351f
C413 B.n336 VSUBS 0.008351f
C414 B.n337 VSUBS 0.008351f
C415 B.n338 VSUBS 0.008351f
C416 B.n339 VSUBS 0.008351f
C417 B.n340 VSUBS 0.008351f
C418 B.n341 VSUBS 0.008351f
C419 B.n342 VSUBS 0.008351f
C420 B.n343 VSUBS 0.008351f
C421 B.n344 VSUBS 0.008351f
C422 B.n345 VSUBS 0.008351f
C423 B.n346 VSUBS 0.008351f
C424 B.n347 VSUBS 0.008351f
C425 B.n348 VSUBS 0.008351f
C426 B.n349 VSUBS 0.008351f
C427 B.n350 VSUBS 0.008351f
C428 B.n351 VSUBS 0.008351f
C429 B.n352 VSUBS 0.008351f
C430 B.n353 VSUBS 0.008351f
C431 B.n354 VSUBS 0.008351f
C432 B.n355 VSUBS 0.008351f
C433 B.n356 VSUBS 0.008351f
C434 B.n357 VSUBS 0.008351f
C435 B.n358 VSUBS 0.008351f
C436 B.n359 VSUBS 0.008351f
C437 B.n360 VSUBS 0.008351f
C438 B.n361 VSUBS 0.008351f
C439 B.n362 VSUBS 0.008351f
C440 B.n363 VSUBS 0.008351f
C441 B.n364 VSUBS 0.008351f
C442 B.n365 VSUBS 0.008351f
C443 B.n366 VSUBS 0.008351f
C444 B.n367 VSUBS 0.008351f
C445 B.n368 VSUBS 0.008351f
C446 B.n369 VSUBS 0.008351f
C447 B.n370 VSUBS 0.008351f
C448 B.n371 VSUBS 0.008351f
C449 B.n372 VSUBS 0.008351f
C450 B.n373 VSUBS 0.008351f
C451 B.n374 VSUBS 0.008351f
C452 B.n375 VSUBS 0.008351f
C453 B.n376 VSUBS 0.008351f
C454 B.n377 VSUBS 0.008351f
C455 B.n378 VSUBS 0.008351f
C456 B.n379 VSUBS 0.008351f
C457 B.n380 VSUBS 0.008351f
C458 B.n381 VSUBS 0.008351f
C459 B.n382 VSUBS 0.008351f
C460 B.n383 VSUBS 0.008351f
C461 B.n384 VSUBS 0.008351f
C462 B.n385 VSUBS 0.008351f
C463 B.n386 VSUBS 0.008351f
C464 B.n387 VSUBS 0.008351f
C465 B.n388 VSUBS 0.008351f
C466 B.n389 VSUBS 0.008351f
C467 B.n390 VSUBS 0.008351f
C468 B.n391 VSUBS 0.008351f
C469 B.n392 VSUBS 0.008351f
C470 B.n393 VSUBS 0.008351f
C471 B.n394 VSUBS 0.008351f
C472 B.n395 VSUBS 0.008351f
C473 B.n396 VSUBS 0.008351f
C474 B.n397 VSUBS 0.008351f
C475 B.n398 VSUBS 0.008351f
C476 B.n399 VSUBS 0.008351f
C477 B.n400 VSUBS 0.008351f
C478 B.n401 VSUBS 0.008351f
C479 B.n402 VSUBS 0.008351f
C480 B.n403 VSUBS 0.008351f
C481 B.n404 VSUBS 0.008351f
C482 B.n405 VSUBS 0.008351f
C483 B.n406 VSUBS 0.008351f
C484 B.n407 VSUBS 0.008351f
C485 B.n408 VSUBS 0.008351f
C486 B.n409 VSUBS 0.020024f
C487 B.n410 VSUBS 0.019767f
C488 B.n411 VSUBS 0.020727f
C489 B.n412 VSUBS 0.008351f
C490 B.n413 VSUBS 0.008351f
C491 B.n414 VSUBS 0.008351f
C492 B.n415 VSUBS 0.008351f
C493 B.n416 VSUBS 0.008351f
C494 B.n417 VSUBS 0.008351f
C495 B.n418 VSUBS 0.008351f
C496 B.n419 VSUBS 0.008351f
C497 B.n420 VSUBS 0.008351f
C498 B.n421 VSUBS 0.008351f
C499 B.n422 VSUBS 0.008351f
C500 B.n423 VSUBS 0.008351f
C501 B.n424 VSUBS 0.008351f
C502 B.n425 VSUBS 0.008351f
C503 B.n426 VSUBS 0.008351f
C504 B.n427 VSUBS 0.008351f
C505 B.n428 VSUBS 0.008351f
C506 B.n429 VSUBS 0.008351f
C507 B.n430 VSUBS 0.008351f
C508 B.n431 VSUBS 0.008351f
C509 B.n432 VSUBS 0.008351f
C510 B.n433 VSUBS 0.008351f
C511 B.n434 VSUBS 0.008351f
C512 B.n435 VSUBS 0.008351f
C513 B.n436 VSUBS 0.008351f
C514 B.n437 VSUBS 0.008351f
C515 B.n438 VSUBS 0.008351f
C516 B.n439 VSUBS 0.008351f
C517 B.n440 VSUBS 0.008351f
C518 B.n441 VSUBS 0.008351f
C519 B.n442 VSUBS 0.008351f
C520 B.n443 VSUBS 0.008351f
C521 B.n444 VSUBS 0.008351f
C522 B.n445 VSUBS 0.008351f
C523 B.n446 VSUBS 0.008351f
C524 B.n447 VSUBS 0.008351f
C525 B.n448 VSUBS 0.008351f
C526 B.n449 VSUBS 0.008351f
C527 B.n450 VSUBS 0.008351f
C528 B.n451 VSUBS 0.008351f
C529 B.n452 VSUBS 0.008351f
C530 B.n453 VSUBS 0.008351f
C531 B.n454 VSUBS 0.008351f
C532 B.n455 VSUBS 0.008351f
C533 B.n456 VSUBS 0.008351f
C534 B.n457 VSUBS 0.008351f
C535 B.n458 VSUBS 0.008351f
C536 B.n459 VSUBS 0.008351f
C537 B.n460 VSUBS 0.019767f
C538 B.n461 VSUBS 0.020024f
C539 B.n462 VSUBS 0.020024f
C540 B.n463 VSUBS 0.008351f
C541 B.n464 VSUBS 0.008351f
C542 B.n465 VSUBS 0.008351f
C543 B.n466 VSUBS 0.008351f
C544 B.n467 VSUBS 0.008351f
C545 B.n468 VSUBS 0.008351f
C546 B.n469 VSUBS 0.008351f
C547 B.n470 VSUBS 0.008351f
C548 B.n471 VSUBS 0.008351f
C549 B.n472 VSUBS 0.008351f
C550 B.n473 VSUBS 0.008351f
C551 B.n474 VSUBS 0.008351f
C552 B.n475 VSUBS 0.008351f
C553 B.n476 VSUBS 0.008351f
C554 B.n477 VSUBS 0.008351f
C555 B.n478 VSUBS 0.008351f
C556 B.n479 VSUBS 0.008351f
C557 B.n480 VSUBS 0.008351f
C558 B.n481 VSUBS 0.008351f
C559 B.n482 VSUBS 0.008351f
C560 B.n483 VSUBS 0.008351f
C561 B.n484 VSUBS 0.008351f
C562 B.n485 VSUBS 0.008351f
C563 B.n486 VSUBS 0.008351f
C564 B.n487 VSUBS 0.008351f
C565 B.n488 VSUBS 0.008351f
C566 B.n489 VSUBS 0.008351f
C567 B.n490 VSUBS 0.008351f
C568 B.n491 VSUBS 0.008351f
C569 B.n492 VSUBS 0.008351f
C570 B.n493 VSUBS 0.008351f
C571 B.n494 VSUBS 0.008351f
C572 B.n495 VSUBS 0.008351f
C573 B.n496 VSUBS 0.008351f
C574 B.n497 VSUBS 0.008351f
C575 B.n498 VSUBS 0.008351f
C576 B.n499 VSUBS 0.008351f
C577 B.n500 VSUBS 0.008351f
C578 B.n501 VSUBS 0.008351f
C579 B.n502 VSUBS 0.008351f
C580 B.n503 VSUBS 0.008351f
C581 B.n504 VSUBS 0.008351f
C582 B.n505 VSUBS 0.008351f
C583 B.n506 VSUBS 0.008351f
C584 B.n507 VSUBS 0.008351f
C585 B.n508 VSUBS 0.008351f
C586 B.n509 VSUBS 0.008351f
C587 B.n510 VSUBS 0.008351f
C588 B.n511 VSUBS 0.008351f
C589 B.n512 VSUBS 0.008351f
C590 B.n513 VSUBS 0.008351f
C591 B.n514 VSUBS 0.008351f
C592 B.n515 VSUBS 0.008351f
C593 B.n516 VSUBS 0.008351f
C594 B.n517 VSUBS 0.008351f
C595 B.n518 VSUBS 0.008351f
C596 B.n519 VSUBS 0.008351f
C597 B.n520 VSUBS 0.008351f
C598 B.n521 VSUBS 0.008351f
C599 B.n522 VSUBS 0.008351f
C600 B.n523 VSUBS 0.008351f
C601 B.n524 VSUBS 0.008351f
C602 B.n525 VSUBS 0.008351f
C603 B.n526 VSUBS 0.008351f
C604 B.n527 VSUBS 0.008351f
C605 B.n528 VSUBS 0.008351f
C606 B.n529 VSUBS 0.008351f
C607 B.n530 VSUBS 0.008351f
C608 B.n531 VSUBS 0.008351f
C609 B.n532 VSUBS 0.008351f
C610 B.n533 VSUBS 0.008351f
C611 B.n534 VSUBS 0.008351f
C612 B.n535 VSUBS 0.008351f
C613 B.n536 VSUBS 0.008351f
C614 B.n537 VSUBS 0.008351f
C615 B.n538 VSUBS 0.008351f
C616 B.n539 VSUBS 0.008351f
C617 B.n540 VSUBS 0.008351f
C618 B.n541 VSUBS 0.008351f
C619 B.n542 VSUBS 0.008351f
C620 B.n543 VSUBS 0.008351f
C621 B.n544 VSUBS 0.008351f
C622 B.n545 VSUBS 0.008351f
C623 B.n546 VSUBS 0.008351f
C624 B.n547 VSUBS 0.008351f
C625 B.n548 VSUBS 0.008351f
C626 B.n549 VSUBS 0.008351f
C627 B.n550 VSUBS 0.008351f
C628 B.n551 VSUBS 0.008351f
C629 B.n552 VSUBS 0.008351f
C630 B.n553 VSUBS 0.008351f
C631 B.n554 VSUBS 0.008351f
C632 B.n555 VSUBS 0.008351f
C633 B.n556 VSUBS 0.005772f
C634 B.n557 VSUBS 0.019349f
C635 B.n558 VSUBS 0.006755f
C636 B.n559 VSUBS 0.008351f
C637 B.n560 VSUBS 0.008351f
C638 B.n561 VSUBS 0.008351f
C639 B.n562 VSUBS 0.008351f
C640 B.n563 VSUBS 0.008351f
C641 B.n564 VSUBS 0.008351f
C642 B.n565 VSUBS 0.008351f
C643 B.n566 VSUBS 0.008351f
C644 B.n567 VSUBS 0.008351f
C645 B.n568 VSUBS 0.008351f
C646 B.n569 VSUBS 0.008351f
C647 B.n570 VSUBS 0.006755f
C648 B.n571 VSUBS 0.008351f
C649 B.n572 VSUBS 0.008351f
C650 B.n573 VSUBS 0.005772f
C651 B.n574 VSUBS 0.008351f
C652 B.n575 VSUBS 0.008351f
C653 B.n576 VSUBS 0.008351f
C654 B.n577 VSUBS 0.008351f
C655 B.n578 VSUBS 0.008351f
C656 B.n579 VSUBS 0.008351f
C657 B.n580 VSUBS 0.008351f
C658 B.n581 VSUBS 0.008351f
C659 B.n582 VSUBS 0.008351f
C660 B.n583 VSUBS 0.008351f
C661 B.n584 VSUBS 0.008351f
C662 B.n585 VSUBS 0.008351f
C663 B.n586 VSUBS 0.008351f
C664 B.n587 VSUBS 0.008351f
C665 B.n588 VSUBS 0.008351f
C666 B.n589 VSUBS 0.008351f
C667 B.n590 VSUBS 0.008351f
C668 B.n591 VSUBS 0.008351f
C669 B.n592 VSUBS 0.008351f
C670 B.n593 VSUBS 0.008351f
C671 B.n594 VSUBS 0.008351f
C672 B.n595 VSUBS 0.008351f
C673 B.n596 VSUBS 0.008351f
C674 B.n597 VSUBS 0.008351f
C675 B.n598 VSUBS 0.008351f
C676 B.n599 VSUBS 0.008351f
C677 B.n600 VSUBS 0.008351f
C678 B.n601 VSUBS 0.008351f
C679 B.n602 VSUBS 0.008351f
C680 B.n603 VSUBS 0.008351f
C681 B.n604 VSUBS 0.008351f
C682 B.n605 VSUBS 0.008351f
C683 B.n606 VSUBS 0.008351f
C684 B.n607 VSUBS 0.008351f
C685 B.n608 VSUBS 0.008351f
C686 B.n609 VSUBS 0.008351f
C687 B.n610 VSUBS 0.008351f
C688 B.n611 VSUBS 0.008351f
C689 B.n612 VSUBS 0.008351f
C690 B.n613 VSUBS 0.008351f
C691 B.n614 VSUBS 0.008351f
C692 B.n615 VSUBS 0.008351f
C693 B.n616 VSUBS 0.008351f
C694 B.n617 VSUBS 0.008351f
C695 B.n618 VSUBS 0.008351f
C696 B.n619 VSUBS 0.008351f
C697 B.n620 VSUBS 0.008351f
C698 B.n621 VSUBS 0.008351f
C699 B.n622 VSUBS 0.008351f
C700 B.n623 VSUBS 0.008351f
C701 B.n624 VSUBS 0.008351f
C702 B.n625 VSUBS 0.008351f
C703 B.n626 VSUBS 0.008351f
C704 B.n627 VSUBS 0.008351f
C705 B.n628 VSUBS 0.008351f
C706 B.n629 VSUBS 0.008351f
C707 B.n630 VSUBS 0.008351f
C708 B.n631 VSUBS 0.008351f
C709 B.n632 VSUBS 0.008351f
C710 B.n633 VSUBS 0.008351f
C711 B.n634 VSUBS 0.008351f
C712 B.n635 VSUBS 0.008351f
C713 B.n636 VSUBS 0.008351f
C714 B.n637 VSUBS 0.008351f
C715 B.n638 VSUBS 0.008351f
C716 B.n639 VSUBS 0.008351f
C717 B.n640 VSUBS 0.008351f
C718 B.n641 VSUBS 0.008351f
C719 B.n642 VSUBS 0.008351f
C720 B.n643 VSUBS 0.008351f
C721 B.n644 VSUBS 0.008351f
C722 B.n645 VSUBS 0.008351f
C723 B.n646 VSUBS 0.008351f
C724 B.n647 VSUBS 0.008351f
C725 B.n648 VSUBS 0.008351f
C726 B.n649 VSUBS 0.008351f
C727 B.n650 VSUBS 0.008351f
C728 B.n651 VSUBS 0.008351f
C729 B.n652 VSUBS 0.008351f
C730 B.n653 VSUBS 0.008351f
C731 B.n654 VSUBS 0.008351f
C732 B.n655 VSUBS 0.008351f
C733 B.n656 VSUBS 0.008351f
C734 B.n657 VSUBS 0.008351f
C735 B.n658 VSUBS 0.008351f
C736 B.n659 VSUBS 0.008351f
C737 B.n660 VSUBS 0.008351f
C738 B.n661 VSUBS 0.008351f
C739 B.n662 VSUBS 0.008351f
C740 B.n663 VSUBS 0.008351f
C741 B.n664 VSUBS 0.008351f
C742 B.n665 VSUBS 0.008351f
C743 B.n666 VSUBS 0.008351f
C744 B.n667 VSUBS 0.020024f
C745 B.n668 VSUBS 0.019767f
C746 B.n669 VSUBS 0.019767f
C747 B.n670 VSUBS 0.008351f
C748 B.n671 VSUBS 0.008351f
C749 B.n672 VSUBS 0.008351f
C750 B.n673 VSUBS 0.008351f
C751 B.n674 VSUBS 0.008351f
C752 B.n675 VSUBS 0.008351f
C753 B.n676 VSUBS 0.008351f
C754 B.n677 VSUBS 0.008351f
C755 B.n678 VSUBS 0.008351f
C756 B.n679 VSUBS 0.008351f
C757 B.n680 VSUBS 0.008351f
C758 B.n681 VSUBS 0.008351f
C759 B.n682 VSUBS 0.008351f
C760 B.n683 VSUBS 0.008351f
C761 B.n684 VSUBS 0.008351f
C762 B.n685 VSUBS 0.008351f
C763 B.n686 VSUBS 0.008351f
C764 B.n687 VSUBS 0.008351f
C765 B.n688 VSUBS 0.008351f
C766 B.n689 VSUBS 0.008351f
C767 B.n690 VSUBS 0.008351f
C768 B.n691 VSUBS 0.010898f
C769 B.n692 VSUBS 0.011609f
C770 B.n693 VSUBS 0.023086f
C771 VDD2.t1 VSUBS 0.570835f
C772 VDD2.t0 VSUBS 0.570835f
C773 VDD2.n0 VSUBS 4.77932f
C774 VDD2.t6 VSUBS 0.570835f
C775 VDD2.t5 VSUBS 0.570835f
C776 VDD2.n1 VSUBS 4.77932f
C777 VDD2.n2 VSUBS 4.37986f
C778 VDD2.t2 VSUBS 0.570835f
C779 VDD2.t7 VSUBS 0.570835f
C780 VDD2.n3 VSUBS 4.77698f
C781 VDD2.n4 VSUBS 4.44122f
C782 VDD2.t4 VSUBS 0.570835f
C783 VDD2.t3 VSUBS 0.570835f
C784 VDD2.n5 VSUBS 4.77927f
C785 VTAIL.t9 VSUBS 0.465775f
C786 VTAIL.t11 VSUBS 0.465775f
C787 VTAIL.n0 VSUBS 3.6955f
C788 VTAIL.n1 VSUBS 0.824482f
C789 VTAIL.n2 VSUBS 0.032917f
C790 VTAIL.n3 VSUBS 0.030072f
C791 VTAIL.n4 VSUBS 0.016159f
C792 VTAIL.n5 VSUBS 0.038195f
C793 VTAIL.n6 VSUBS 0.01711f
C794 VTAIL.n7 VSUBS 0.030072f
C795 VTAIL.n8 VSUBS 0.016159f
C796 VTAIL.n9 VSUBS 0.038195f
C797 VTAIL.n10 VSUBS 0.01711f
C798 VTAIL.n11 VSUBS 0.030072f
C799 VTAIL.n12 VSUBS 0.016159f
C800 VTAIL.n13 VSUBS 0.038195f
C801 VTAIL.n14 VSUBS 0.016635f
C802 VTAIL.n15 VSUBS 0.030072f
C803 VTAIL.n16 VSUBS 0.01711f
C804 VTAIL.n17 VSUBS 0.038195f
C805 VTAIL.n18 VSUBS 0.01711f
C806 VTAIL.n19 VSUBS 0.030072f
C807 VTAIL.n20 VSUBS 0.016159f
C808 VTAIL.n21 VSUBS 0.038195f
C809 VTAIL.n22 VSUBS 0.01711f
C810 VTAIL.n23 VSUBS 0.030072f
C811 VTAIL.n24 VSUBS 0.016159f
C812 VTAIL.n25 VSUBS 0.038195f
C813 VTAIL.n26 VSUBS 0.01711f
C814 VTAIL.n27 VSUBS 0.030072f
C815 VTAIL.n28 VSUBS 0.016159f
C816 VTAIL.n29 VSUBS 0.038195f
C817 VTAIL.n30 VSUBS 0.01711f
C818 VTAIL.n31 VSUBS 0.030072f
C819 VTAIL.n32 VSUBS 0.016159f
C820 VTAIL.n33 VSUBS 0.038195f
C821 VTAIL.n34 VSUBS 0.01711f
C822 VTAIL.n35 VSUBS 2.54817f
C823 VTAIL.n36 VSUBS 0.016159f
C824 VTAIL.t14 VSUBS 0.082112f
C825 VTAIL.n37 VSUBS 0.252786f
C826 VTAIL.n38 VSUBS 0.024298f
C827 VTAIL.n39 VSUBS 0.028646f
C828 VTAIL.n40 VSUBS 0.038195f
C829 VTAIL.n41 VSUBS 0.01711f
C830 VTAIL.n42 VSUBS 0.016159f
C831 VTAIL.n43 VSUBS 0.030072f
C832 VTAIL.n44 VSUBS 0.030072f
C833 VTAIL.n45 VSUBS 0.016159f
C834 VTAIL.n46 VSUBS 0.01711f
C835 VTAIL.n47 VSUBS 0.038195f
C836 VTAIL.n48 VSUBS 0.038195f
C837 VTAIL.n49 VSUBS 0.01711f
C838 VTAIL.n50 VSUBS 0.016159f
C839 VTAIL.n51 VSUBS 0.030072f
C840 VTAIL.n52 VSUBS 0.030072f
C841 VTAIL.n53 VSUBS 0.016159f
C842 VTAIL.n54 VSUBS 0.01711f
C843 VTAIL.n55 VSUBS 0.038195f
C844 VTAIL.n56 VSUBS 0.038195f
C845 VTAIL.n57 VSUBS 0.01711f
C846 VTAIL.n58 VSUBS 0.016159f
C847 VTAIL.n59 VSUBS 0.030072f
C848 VTAIL.n60 VSUBS 0.030072f
C849 VTAIL.n61 VSUBS 0.016159f
C850 VTAIL.n62 VSUBS 0.01711f
C851 VTAIL.n63 VSUBS 0.038195f
C852 VTAIL.n64 VSUBS 0.038195f
C853 VTAIL.n65 VSUBS 0.01711f
C854 VTAIL.n66 VSUBS 0.016159f
C855 VTAIL.n67 VSUBS 0.030072f
C856 VTAIL.n68 VSUBS 0.030072f
C857 VTAIL.n69 VSUBS 0.016159f
C858 VTAIL.n70 VSUBS 0.01711f
C859 VTAIL.n71 VSUBS 0.038195f
C860 VTAIL.n72 VSUBS 0.038195f
C861 VTAIL.n73 VSUBS 0.01711f
C862 VTAIL.n74 VSUBS 0.016159f
C863 VTAIL.n75 VSUBS 0.030072f
C864 VTAIL.n76 VSUBS 0.030072f
C865 VTAIL.n77 VSUBS 0.016159f
C866 VTAIL.n78 VSUBS 0.016159f
C867 VTAIL.n79 VSUBS 0.01711f
C868 VTAIL.n80 VSUBS 0.038195f
C869 VTAIL.n81 VSUBS 0.038195f
C870 VTAIL.n82 VSUBS 0.038195f
C871 VTAIL.n83 VSUBS 0.016635f
C872 VTAIL.n84 VSUBS 0.016159f
C873 VTAIL.n85 VSUBS 0.030072f
C874 VTAIL.n86 VSUBS 0.030072f
C875 VTAIL.n87 VSUBS 0.016159f
C876 VTAIL.n88 VSUBS 0.01711f
C877 VTAIL.n89 VSUBS 0.038195f
C878 VTAIL.n90 VSUBS 0.038195f
C879 VTAIL.n91 VSUBS 0.01711f
C880 VTAIL.n92 VSUBS 0.016159f
C881 VTAIL.n93 VSUBS 0.030072f
C882 VTAIL.n94 VSUBS 0.030072f
C883 VTAIL.n95 VSUBS 0.016159f
C884 VTAIL.n96 VSUBS 0.01711f
C885 VTAIL.n97 VSUBS 0.038195f
C886 VTAIL.n98 VSUBS 0.038195f
C887 VTAIL.n99 VSUBS 0.01711f
C888 VTAIL.n100 VSUBS 0.016159f
C889 VTAIL.n101 VSUBS 0.030072f
C890 VTAIL.n102 VSUBS 0.030072f
C891 VTAIL.n103 VSUBS 0.016159f
C892 VTAIL.n104 VSUBS 0.01711f
C893 VTAIL.n105 VSUBS 0.038195f
C894 VTAIL.n106 VSUBS 0.092038f
C895 VTAIL.n107 VSUBS 0.01711f
C896 VTAIL.n108 VSUBS 0.016159f
C897 VTAIL.n109 VSUBS 0.066224f
C898 VTAIL.n110 VSUBS 0.046163f
C899 VTAIL.n111 VSUBS 0.116136f
C900 VTAIL.n112 VSUBS 0.032917f
C901 VTAIL.n113 VSUBS 0.030072f
C902 VTAIL.n114 VSUBS 0.016159f
C903 VTAIL.n115 VSUBS 0.038195f
C904 VTAIL.n116 VSUBS 0.01711f
C905 VTAIL.n117 VSUBS 0.030072f
C906 VTAIL.n118 VSUBS 0.016159f
C907 VTAIL.n119 VSUBS 0.038195f
C908 VTAIL.n120 VSUBS 0.01711f
C909 VTAIL.n121 VSUBS 0.030072f
C910 VTAIL.n122 VSUBS 0.016159f
C911 VTAIL.n123 VSUBS 0.038195f
C912 VTAIL.n124 VSUBS 0.016635f
C913 VTAIL.n125 VSUBS 0.030072f
C914 VTAIL.n126 VSUBS 0.01711f
C915 VTAIL.n127 VSUBS 0.038195f
C916 VTAIL.n128 VSUBS 0.01711f
C917 VTAIL.n129 VSUBS 0.030072f
C918 VTAIL.n130 VSUBS 0.016159f
C919 VTAIL.n131 VSUBS 0.038195f
C920 VTAIL.n132 VSUBS 0.01711f
C921 VTAIL.n133 VSUBS 0.030072f
C922 VTAIL.n134 VSUBS 0.016159f
C923 VTAIL.n135 VSUBS 0.038195f
C924 VTAIL.n136 VSUBS 0.01711f
C925 VTAIL.n137 VSUBS 0.030072f
C926 VTAIL.n138 VSUBS 0.016159f
C927 VTAIL.n139 VSUBS 0.038195f
C928 VTAIL.n140 VSUBS 0.01711f
C929 VTAIL.n141 VSUBS 0.030072f
C930 VTAIL.n142 VSUBS 0.016159f
C931 VTAIL.n143 VSUBS 0.038195f
C932 VTAIL.n144 VSUBS 0.01711f
C933 VTAIL.n145 VSUBS 2.54817f
C934 VTAIL.n146 VSUBS 0.016159f
C935 VTAIL.t4 VSUBS 0.082112f
C936 VTAIL.n147 VSUBS 0.252786f
C937 VTAIL.n148 VSUBS 0.024298f
C938 VTAIL.n149 VSUBS 0.028646f
C939 VTAIL.n150 VSUBS 0.038195f
C940 VTAIL.n151 VSUBS 0.01711f
C941 VTAIL.n152 VSUBS 0.016159f
C942 VTAIL.n153 VSUBS 0.030072f
C943 VTAIL.n154 VSUBS 0.030072f
C944 VTAIL.n155 VSUBS 0.016159f
C945 VTAIL.n156 VSUBS 0.01711f
C946 VTAIL.n157 VSUBS 0.038195f
C947 VTAIL.n158 VSUBS 0.038195f
C948 VTAIL.n159 VSUBS 0.01711f
C949 VTAIL.n160 VSUBS 0.016159f
C950 VTAIL.n161 VSUBS 0.030072f
C951 VTAIL.n162 VSUBS 0.030072f
C952 VTAIL.n163 VSUBS 0.016159f
C953 VTAIL.n164 VSUBS 0.01711f
C954 VTAIL.n165 VSUBS 0.038195f
C955 VTAIL.n166 VSUBS 0.038195f
C956 VTAIL.n167 VSUBS 0.01711f
C957 VTAIL.n168 VSUBS 0.016159f
C958 VTAIL.n169 VSUBS 0.030072f
C959 VTAIL.n170 VSUBS 0.030072f
C960 VTAIL.n171 VSUBS 0.016159f
C961 VTAIL.n172 VSUBS 0.01711f
C962 VTAIL.n173 VSUBS 0.038195f
C963 VTAIL.n174 VSUBS 0.038195f
C964 VTAIL.n175 VSUBS 0.01711f
C965 VTAIL.n176 VSUBS 0.016159f
C966 VTAIL.n177 VSUBS 0.030072f
C967 VTAIL.n178 VSUBS 0.030072f
C968 VTAIL.n179 VSUBS 0.016159f
C969 VTAIL.n180 VSUBS 0.01711f
C970 VTAIL.n181 VSUBS 0.038195f
C971 VTAIL.n182 VSUBS 0.038195f
C972 VTAIL.n183 VSUBS 0.01711f
C973 VTAIL.n184 VSUBS 0.016159f
C974 VTAIL.n185 VSUBS 0.030072f
C975 VTAIL.n186 VSUBS 0.030072f
C976 VTAIL.n187 VSUBS 0.016159f
C977 VTAIL.n188 VSUBS 0.016159f
C978 VTAIL.n189 VSUBS 0.01711f
C979 VTAIL.n190 VSUBS 0.038195f
C980 VTAIL.n191 VSUBS 0.038195f
C981 VTAIL.n192 VSUBS 0.038195f
C982 VTAIL.n193 VSUBS 0.016635f
C983 VTAIL.n194 VSUBS 0.016159f
C984 VTAIL.n195 VSUBS 0.030072f
C985 VTAIL.n196 VSUBS 0.030072f
C986 VTAIL.n197 VSUBS 0.016159f
C987 VTAIL.n198 VSUBS 0.01711f
C988 VTAIL.n199 VSUBS 0.038195f
C989 VTAIL.n200 VSUBS 0.038195f
C990 VTAIL.n201 VSUBS 0.01711f
C991 VTAIL.n202 VSUBS 0.016159f
C992 VTAIL.n203 VSUBS 0.030072f
C993 VTAIL.n204 VSUBS 0.030072f
C994 VTAIL.n205 VSUBS 0.016159f
C995 VTAIL.n206 VSUBS 0.01711f
C996 VTAIL.n207 VSUBS 0.038195f
C997 VTAIL.n208 VSUBS 0.038195f
C998 VTAIL.n209 VSUBS 0.01711f
C999 VTAIL.n210 VSUBS 0.016159f
C1000 VTAIL.n211 VSUBS 0.030072f
C1001 VTAIL.n212 VSUBS 0.030072f
C1002 VTAIL.n213 VSUBS 0.016159f
C1003 VTAIL.n214 VSUBS 0.01711f
C1004 VTAIL.n215 VSUBS 0.038195f
C1005 VTAIL.n216 VSUBS 0.092038f
C1006 VTAIL.n217 VSUBS 0.01711f
C1007 VTAIL.n218 VSUBS 0.016159f
C1008 VTAIL.n219 VSUBS 0.066224f
C1009 VTAIL.n220 VSUBS 0.046163f
C1010 VTAIL.n221 VSUBS 0.116136f
C1011 VTAIL.t7 VSUBS 0.465775f
C1012 VTAIL.t6 VSUBS 0.465775f
C1013 VTAIL.n222 VSUBS 3.6955f
C1014 VTAIL.n223 VSUBS 0.865623f
C1015 VTAIL.n224 VSUBS 0.032917f
C1016 VTAIL.n225 VSUBS 0.030072f
C1017 VTAIL.n226 VSUBS 0.016159f
C1018 VTAIL.n227 VSUBS 0.038195f
C1019 VTAIL.n228 VSUBS 0.01711f
C1020 VTAIL.n229 VSUBS 0.030072f
C1021 VTAIL.n230 VSUBS 0.016159f
C1022 VTAIL.n231 VSUBS 0.038195f
C1023 VTAIL.n232 VSUBS 0.01711f
C1024 VTAIL.n233 VSUBS 0.030072f
C1025 VTAIL.n234 VSUBS 0.016159f
C1026 VTAIL.n235 VSUBS 0.038195f
C1027 VTAIL.n236 VSUBS 0.016635f
C1028 VTAIL.n237 VSUBS 0.030072f
C1029 VTAIL.n238 VSUBS 0.01711f
C1030 VTAIL.n239 VSUBS 0.038195f
C1031 VTAIL.n240 VSUBS 0.01711f
C1032 VTAIL.n241 VSUBS 0.030072f
C1033 VTAIL.n242 VSUBS 0.016159f
C1034 VTAIL.n243 VSUBS 0.038195f
C1035 VTAIL.n244 VSUBS 0.01711f
C1036 VTAIL.n245 VSUBS 0.030072f
C1037 VTAIL.n246 VSUBS 0.016159f
C1038 VTAIL.n247 VSUBS 0.038195f
C1039 VTAIL.n248 VSUBS 0.01711f
C1040 VTAIL.n249 VSUBS 0.030072f
C1041 VTAIL.n250 VSUBS 0.016159f
C1042 VTAIL.n251 VSUBS 0.038195f
C1043 VTAIL.n252 VSUBS 0.01711f
C1044 VTAIL.n253 VSUBS 0.030072f
C1045 VTAIL.n254 VSUBS 0.016159f
C1046 VTAIL.n255 VSUBS 0.038195f
C1047 VTAIL.n256 VSUBS 0.01711f
C1048 VTAIL.n257 VSUBS 2.54817f
C1049 VTAIL.n258 VSUBS 0.016159f
C1050 VTAIL.t0 VSUBS 0.082112f
C1051 VTAIL.n259 VSUBS 0.252786f
C1052 VTAIL.n260 VSUBS 0.024298f
C1053 VTAIL.n261 VSUBS 0.028646f
C1054 VTAIL.n262 VSUBS 0.038195f
C1055 VTAIL.n263 VSUBS 0.01711f
C1056 VTAIL.n264 VSUBS 0.016159f
C1057 VTAIL.n265 VSUBS 0.030072f
C1058 VTAIL.n266 VSUBS 0.030072f
C1059 VTAIL.n267 VSUBS 0.016159f
C1060 VTAIL.n268 VSUBS 0.01711f
C1061 VTAIL.n269 VSUBS 0.038195f
C1062 VTAIL.n270 VSUBS 0.038195f
C1063 VTAIL.n271 VSUBS 0.01711f
C1064 VTAIL.n272 VSUBS 0.016159f
C1065 VTAIL.n273 VSUBS 0.030072f
C1066 VTAIL.n274 VSUBS 0.030072f
C1067 VTAIL.n275 VSUBS 0.016159f
C1068 VTAIL.n276 VSUBS 0.01711f
C1069 VTAIL.n277 VSUBS 0.038195f
C1070 VTAIL.n278 VSUBS 0.038195f
C1071 VTAIL.n279 VSUBS 0.01711f
C1072 VTAIL.n280 VSUBS 0.016159f
C1073 VTAIL.n281 VSUBS 0.030072f
C1074 VTAIL.n282 VSUBS 0.030072f
C1075 VTAIL.n283 VSUBS 0.016159f
C1076 VTAIL.n284 VSUBS 0.01711f
C1077 VTAIL.n285 VSUBS 0.038195f
C1078 VTAIL.n286 VSUBS 0.038195f
C1079 VTAIL.n287 VSUBS 0.01711f
C1080 VTAIL.n288 VSUBS 0.016159f
C1081 VTAIL.n289 VSUBS 0.030072f
C1082 VTAIL.n290 VSUBS 0.030072f
C1083 VTAIL.n291 VSUBS 0.016159f
C1084 VTAIL.n292 VSUBS 0.01711f
C1085 VTAIL.n293 VSUBS 0.038195f
C1086 VTAIL.n294 VSUBS 0.038195f
C1087 VTAIL.n295 VSUBS 0.01711f
C1088 VTAIL.n296 VSUBS 0.016159f
C1089 VTAIL.n297 VSUBS 0.030072f
C1090 VTAIL.n298 VSUBS 0.030072f
C1091 VTAIL.n299 VSUBS 0.016159f
C1092 VTAIL.n300 VSUBS 0.016159f
C1093 VTAIL.n301 VSUBS 0.01711f
C1094 VTAIL.n302 VSUBS 0.038195f
C1095 VTAIL.n303 VSUBS 0.038195f
C1096 VTAIL.n304 VSUBS 0.038195f
C1097 VTAIL.n305 VSUBS 0.016635f
C1098 VTAIL.n306 VSUBS 0.016159f
C1099 VTAIL.n307 VSUBS 0.030072f
C1100 VTAIL.n308 VSUBS 0.030072f
C1101 VTAIL.n309 VSUBS 0.016159f
C1102 VTAIL.n310 VSUBS 0.01711f
C1103 VTAIL.n311 VSUBS 0.038195f
C1104 VTAIL.n312 VSUBS 0.038195f
C1105 VTAIL.n313 VSUBS 0.01711f
C1106 VTAIL.n314 VSUBS 0.016159f
C1107 VTAIL.n315 VSUBS 0.030072f
C1108 VTAIL.n316 VSUBS 0.030072f
C1109 VTAIL.n317 VSUBS 0.016159f
C1110 VTAIL.n318 VSUBS 0.01711f
C1111 VTAIL.n319 VSUBS 0.038195f
C1112 VTAIL.n320 VSUBS 0.038195f
C1113 VTAIL.n321 VSUBS 0.01711f
C1114 VTAIL.n322 VSUBS 0.016159f
C1115 VTAIL.n323 VSUBS 0.030072f
C1116 VTAIL.n324 VSUBS 0.030072f
C1117 VTAIL.n325 VSUBS 0.016159f
C1118 VTAIL.n326 VSUBS 0.01711f
C1119 VTAIL.n327 VSUBS 0.038195f
C1120 VTAIL.n328 VSUBS 0.092038f
C1121 VTAIL.n329 VSUBS 0.01711f
C1122 VTAIL.n330 VSUBS 0.016159f
C1123 VTAIL.n331 VSUBS 0.066224f
C1124 VTAIL.n332 VSUBS 0.046163f
C1125 VTAIL.n333 VSUBS 2.16315f
C1126 VTAIL.n334 VSUBS 0.032917f
C1127 VTAIL.n335 VSUBS 0.030072f
C1128 VTAIL.n336 VSUBS 0.016159f
C1129 VTAIL.n337 VSUBS 0.038195f
C1130 VTAIL.n338 VSUBS 0.01711f
C1131 VTAIL.n339 VSUBS 0.030072f
C1132 VTAIL.n340 VSUBS 0.016159f
C1133 VTAIL.n341 VSUBS 0.038195f
C1134 VTAIL.n342 VSUBS 0.01711f
C1135 VTAIL.n343 VSUBS 0.030072f
C1136 VTAIL.n344 VSUBS 0.016159f
C1137 VTAIL.n345 VSUBS 0.038195f
C1138 VTAIL.n346 VSUBS 0.016635f
C1139 VTAIL.n347 VSUBS 0.030072f
C1140 VTAIL.n348 VSUBS 0.016635f
C1141 VTAIL.n349 VSUBS 0.016159f
C1142 VTAIL.n350 VSUBS 0.038195f
C1143 VTAIL.n351 VSUBS 0.038195f
C1144 VTAIL.n352 VSUBS 0.01711f
C1145 VTAIL.n353 VSUBS 0.030072f
C1146 VTAIL.n354 VSUBS 0.016159f
C1147 VTAIL.n355 VSUBS 0.038195f
C1148 VTAIL.n356 VSUBS 0.01711f
C1149 VTAIL.n357 VSUBS 0.030072f
C1150 VTAIL.n358 VSUBS 0.016159f
C1151 VTAIL.n359 VSUBS 0.038195f
C1152 VTAIL.n360 VSUBS 0.01711f
C1153 VTAIL.n361 VSUBS 0.030072f
C1154 VTAIL.n362 VSUBS 0.016159f
C1155 VTAIL.n363 VSUBS 0.038195f
C1156 VTAIL.n364 VSUBS 0.01711f
C1157 VTAIL.n365 VSUBS 0.030072f
C1158 VTAIL.n366 VSUBS 0.016159f
C1159 VTAIL.n367 VSUBS 0.038195f
C1160 VTAIL.n368 VSUBS 0.01711f
C1161 VTAIL.n369 VSUBS 2.54816f
C1162 VTAIL.n370 VSUBS 0.016159f
C1163 VTAIL.t8 VSUBS 0.082112f
C1164 VTAIL.n371 VSUBS 0.252786f
C1165 VTAIL.n372 VSUBS 0.024298f
C1166 VTAIL.n373 VSUBS 0.028646f
C1167 VTAIL.n374 VSUBS 0.038195f
C1168 VTAIL.n375 VSUBS 0.01711f
C1169 VTAIL.n376 VSUBS 0.016159f
C1170 VTAIL.n377 VSUBS 0.030072f
C1171 VTAIL.n378 VSUBS 0.030072f
C1172 VTAIL.n379 VSUBS 0.016159f
C1173 VTAIL.n380 VSUBS 0.01711f
C1174 VTAIL.n381 VSUBS 0.038195f
C1175 VTAIL.n382 VSUBS 0.038195f
C1176 VTAIL.n383 VSUBS 0.01711f
C1177 VTAIL.n384 VSUBS 0.016159f
C1178 VTAIL.n385 VSUBS 0.030072f
C1179 VTAIL.n386 VSUBS 0.030072f
C1180 VTAIL.n387 VSUBS 0.016159f
C1181 VTAIL.n388 VSUBS 0.01711f
C1182 VTAIL.n389 VSUBS 0.038195f
C1183 VTAIL.n390 VSUBS 0.038195f
C1184 VTAIL.n391 VSUBS 0.01711f
C1185 VTAIL.n392 VSUBS 0.016159f
C1186 VTAIL.n393 VSUBS 0.030072f
C1187 VTAIL.n394 VSUBS 0.030072f
C1188 VTAIL.n395 VSUBS 0.016159f
C1189 VTAIL.n396 VSUBS 0.01711f
C1190 VTAIL.n397 VSUBS 0.038195f
C1191 VTAIL.n398 VSUBS 0.038195f
C1192 VTAIL.n399 VSUBS 0.01711f
C1193 VTAIL.n400 VSUBS 0.016159f
C1194 VTAIL.n401 VSUBS 0.030072f
C1195 VTAIL.n402 VSUBS 0.030072f
C1196 VTAIL.n403 VSUBS 0.016159f
C1197 VTAIL.n404 VSUBS 0.01711f
C1198 VTAIL.n405 VSUBS 0.038195f
C1199 VTAIL.n406 VSUBS 0.038195f
C1200 VTAIL.n407 VSUBS 0.01711f
C1201 VTAIL.n408 VSUBS 0.016159f
C1202 VTAIL.n409 VSUBS 0.030072f
C1203 VTAIL.n410 VSUBS 0.030072f
C1204 VTAIL.n411 VSUBS 0.016159f
C1205 VTAIL.n412 VSUBS 0.01711f
C1206 VTAIL.n413 VSUBS 0.038195f
C1207 VTAIL.n414 VSUBS 0.038195f
C1208 VTAIL.n415 VSUBS 0.01711f
C1209 VTAIL.n416 VSUBS 0.016159f
C1210 VTAIL.n417 VSUBS 0.030072f
C1211 VTAIL.n418 VSUBS 0.030072f
C1212 VTAIL.n419 VSUBS 0.016159f
C1213 VTAIL.n420 VSUBS 0.01711f
C1214 VTAIL.n421 VSUBS 0.038195f
C1215 VTAIL.n422 VSUBS 0.038195f
C1216 VTAIL.n423 VSUBS 0.01711f
C1217 VTAIL.n424 VSUBS 0.016159f
C1218 VTAIL.n425 VSUBS 0.030072f
C1219 VTAIL.n426 VSUBS 0.030072f
C1220 VTAIL.n427 VSUBS 0.016159f
C1221 VTAIL.n428 VSUBS 0.01711f
C1222 VTAIL.n429 VSUBS 0.038195f
C1223 VTAIL.n430 VSUBS 0.038195f
C1224 VTAIL.n431 VSUBS 0.01711f
C1225 VTAIL.n432 VSUBS 0.016159f
C1226 VTAIL.n433 VSUBS 0.030072f
C1227 VTAIL.n434 VSUBS 0.030072f
C1228 VTAIL.n435 VSUBS 0.016159f
C1229 VTAIL.n436 VSUBS 0.01711f
C1230 VTAIL.n437 VSUBS 0.038195f
C1231 VTAIL.n438 VSUBS 0.092038f
C1232 VTAIL.n439 VSUBS 0.01711f
C1233 VTAIL.n440 VSUBS 0.016159f
C1234 VTAIL.n441 VSUBS 0.066224f
C1235 VTAIL.n442 VSUBS 0.046163f
C1236 VTAIL.n443 VSUBS 2.16315f
C1237 VTAIL.t12 VSUBS 0.465775f
C1238 VTAIL.t15 VSUBS 0.465775f
C1239 VTAIL.n444 VSUBS 3.69552f
C1240 VTAIL.n445 VSUBS 0.865601f
C1241 VTAIL.n446 VSUBS 0.032917f
C1242 VTAIL.n447 VSUBS 0.030072f
C1243 VTAIL.n448 VSUBS 0.016159f
C1244 VTAIL.n449 VSUBS 0.038195f
C1245 VTAIL.n450 VSUBS 0.01711f
C1246 VTAIL.n451 VSUBS 0.030072f
C1247 VTAIL.n452 VSUBS 0.016159f
C1248 VTAIL.n453 VSUBS 0.038195f
C1249 VTAIL.n454 VSUBS 0.01711f
C1250 VTAIL.n455 VSUBS 0.030072f
C1251 VTAIL.n456 VSUBS 0.016159f
C1252 VTAIL.n457 VSUBS 0.038195f
C1253 VTAIL.n458 VSUBS 0.016635f
C1254 VTAIL.n459 VSUBS 0.030072f
C1255 VTAIL.n460 VSUBS 0.016635f
C1256 VTAIL.n461 VSUBS 0.016159f
C1257 VTAIL.n462 VSUBS 0.038195f
C1258 VTAIL.n463 VSUBS 0.038195f
C1259 VTAIL.n464 VSUBS 0.01711f
C1260 VTAIL.n465 VSUBS 0.030072f
C1261 VTAIL.n466 VSUBS 0.016159f
C1262 VTAIL.n467 VSUBS 0.038195f
C1263 VTAIL.n468 VSUBS 0.01711f
C1264 VTAIL.n469 VSUBS 0.030072f
C1265 VTAIL.n470 VSUBS 0.016159f
C1266 VTAIL.n471 VSUBS 0.038195f
C1267 VTAIL.n472 VSUBS 0.01711f
C1268 VTAIL.n473 VSUBS 0.030072f
C1269 VTAIL.n474 VSUBS 0.016159f
C1270 VTAIL.n475 VSUBS 0.038195f
C1271 VTAIL.n476 VSUBS 0.01711f
C1272 VTAIL.n477 VSUBS 0.030072f
C1273 VTAIL.n478 VSUBS 0.016159f
C1274 VTAIL.n479 VSUBS 0.038195f
C1275 VTAIL.n480 VSUBS 0.01711f
C1276 VTAIL.n481 VSUBS 2.54816f
C1277 VTAIL.n482 VSUBS 0.016159f
C1278 VTAIL.t13 VSUBS 0.082112f
C1279 VTAIL.n483 VSUBS 0.252786f
C1280 VTAIL.n484 VSUBS 0.024298f
C1281 VTAIL.n485 VSUBS 0.028646f
C1282 VTAIL.n486 VSUBS 0.038195f
C1283 VTAIL.n487 VSUBS 0.01711f
C1284 VTAIL.n488 VSUBS 0.016159f
C1285 VTAIL.n489 VSUBS 0.030072f
C1286 VTAIL.n490 VSUBS 0.030072f
C1287 VTAIL.n491 VSUBS 0.016159f
C1288 VTAIL.n492 VSUBS 0.01711f
C1289 VTAIL.n493 VSUBS 0.038195f
C1290 VTAIL.n494 VSUBS 0.038195f
C1291 VTAIL.n495 VSUBS 0.01711f
C1292 VTAIL.n496 VSUBS 0.016159f
C1293 VTAIL.n497 VSUBS 0.030072f
C1294 VTAIL.n498 VSUBS 0.030072f
C1295 VTAIL.n499 VSUBS 0.016159f
C1296 VTAIL.n500 VSUBS 0.01711f
C1297 VTAIL.n501 VSUBS 0.038195f
C1298 VTAIL.n502 VSUBS 0.038195f
C1299 VTAIL.n503 VSUBS 0.01711f
C1300 VTAIL.n504 VSUBS 0.016159f
C1301 VTAIL.n505 VSUBS 0.030072f
C1302 VTAIL.n506 VSUBS 0.030072f
C1303 VTAIL.n507 VSUBS 0.016159f
C1304 VTAIL.n508 VSUBS 0.01711f
C1305 VTAIL.n509 VSUBS 0.038195f
C1306 VTAIL.n510 VSUBS 0.038195f
C1307 VTAIL.n511 VSUBS 0.01711f
C1308 VTAIL.n512 VSUBS 0.016159f
C1309 VTAIL.n513 VSUBS 0.030072f
C1310 VTAIL.n514 VSUBS 0.030072f
C1311 VTAIL.n515 VSUBS 0.016159f
C1312 VTAIL.n516 VSUBS 0.01711f
C1313 VTAIL.n517 VSUBS 0.038195f
C1314 VTAIL.n518 VSUBS 0.038195f
C1315 VTAIL.n519 VSUBS 0.01711f
C1316 VTAIL.n520 VSUBS 0.016159f
C1317 VTAIL.n521 VSUBS 0.030072f
C1318 VTAIL.n522 VSUBS 0.030072f
C1319 VTAIL.n523 VSUBS 0.016159f
C1320 VTAIL.n524 VSUBS 0.01711f
C1321 VTAIL.n525 VSUBS 0.038195f
C1322 VTAIL.n526 VSUBS 0.038195f
C1323 VTAIL.n527 VSUBS 0.01711f
C1324 VTAIL.n528 VSUBS 0.016159f
C1325 VTAIL.n529 VSUBS 0.030072f
C1326 VTAIL.n530 VSUBS 0.030072f
C1327 VTAIL.n531 VSUBS 0.016159f
C1328 VTAIL.n532 VSUBS 0.01711f
C1329 VTAIL.n533 VSUBS 0.038195f
C1330 VTAIL.n534 VSUBS 0.038195f
C1331 VTAIL.n535 VSUBS 0.01711f
C1332 VTAIL.n536 VSUBS 0.016159f
C1333 VTAIL.n537 VSUBS 0.030072f
C1334 VTAIL.n538 VSUBS 0.030072f
C1335 VTAIL.n539 VSUBS 0.016159f
C1336 VTAIL.n540 VSUBS 0.01711f
C1337 VTAIL.n541 VSUBS 0.038195f
C1338 VTAIL.n542 VSUBS 0.038195f
C1339 VTAIL.n543 VSUBS 0.01711f
C1340 VTAIL.n544 VSUBS 0.016159f
C1341 VTAIL.n545 VSUBS 0.030072f
C1342 VTAIL.n546 VSUBS 0.030072f
C1343 VTAIL.n547 VSUBS 0.016159f
C1344 VTAIL.n548 VSUBS 0.01711f
C1345 VTAIL.n549 VSUBS 0.038195f
C1346 VTAIL.n550 VSUBS 0.092038f
C1347 VTAIL.n551 VSUBS 0.01711f
C1348 VTAIL.n552 VSUBS 0.016159f
C1349 VTAIL.n553 VSUBS 0.066224f
C1350 VTAIL.n554 VSUBS 0.046163f
C1351 VTAIL.n555 VSUBS 0.116136f
C1352 VTAIL.n556 VSUBS 0.032917f
C1353 VTAIL.n557 VSUBS 0.030072f
C1354 VTAIL.n558 VSUBS 0.016159f
C1355 VTAIL.n559 VSUBS 0.038195f
C1356 VTAIL.n560 VSUBS 0.01711f
C1357 VTAIL.n561 VSUBS 0.030072f
C1358 VTAIL.n562 VSUBS 0.016159f
C1359 VTAIL.n563 VSUBS 0.038195f
C1360 VTAIL.n564 VSUBS 0.01711f
C1361 VTAIL.n565 VSUBS 0.030072f
C1362 VTAIL.n566 VSUBS 0.016159f
C1363 VTAIL.n567 VSUBS 0.038195f
C1364 VTAIL.n568 VSUBS 0.016635f
C1365 VTAIL.n569 VSUBS 0.030072f
C1366 VTAIL.n570 VSUBS 0.016635f
C1367 VTAIL.n571 VSUBS 0.016159f
C1368 VTAIL.n572 VSUBS 0.038195f
C1369 VTAIL.n573 VSUBS 0.038195f
C1370 VTAIL.n574 VSUBS 0.01711f
C1371 VTAIL.n575 VSUBS 0.030072f
C1372 VTAIL.n576 VSUBS 0.016159f
C1373 VTAIL.n577 VSUBS 0.038195f
C1374 VTAIL.n578 VSUBS 0.01711f
C1375 VTAIL.n579 VSUBS 0.030072f
C1376 VTAIL.n580 VSUBS 0.016159f
C1377 VTAIL.n581 VSUBS 0.038195f
C1378 VTAIL.n582 VSUBS 0.01711f
C1379 VTAIL.n583 VSUBS 0.030072f
C1380 VTAIL.n584 VSUBS 0.016159f
C1381 VTAIL.n585 VSUBS 0.038195f
C1382 VTAIL.n586 VSUBS 0.01711f
C1383 VTAIL.n587 VSUBS 0.030072f
C1384 VTAIL.n588 VSUBS 0.016159f
C1385 VTAIL.n589 VSUBS 0.038195f
C1386 VTAIL.n590 VSUBS 0.01711f
C1387 VTAIL.n591 VSUBS 2.54816f
C1388 VTAIL.n592 VSUBS 0.016159f
C1389 VTAIL.t5 VSUBS 0.082112f
C1390 VTAIL.n593 VSUBS 0.252786f
C1391 VTAIL.n594 VSUBS 0.024298f
C1392 VTAIL.n595 VSUBS 0.028646f
C1393 VTAIL.n596 VSUBS 0.038195f
C1394 VTAIL.n597 VSUBS 0.01711f
C1395 VTAIL.n598 VSUBS 0.016159f
C1396 VTAIL.n599 VSUBS 0.030072f
C1397 VTAIL.n600 VSUBS 0.030072f
C1398 VTAIL.n601 VSUBS 0.016159f
C1399 VTAIL.n602 VSUBS 0.01711f
C1400 VTAIL.n603 VSUBS 0.038195f
C1401 VTAIL.n604 VSUBS 0.038195f
C1402 VTAIL.n605 VSUBS 0.01711f
C1403 VTAIL.n606 VSUBS 0.016159f
C1404 VTAIL.n607 VSUBS 0.030072f
C1405 VTAIL.n608 VSUBS 0.030072f
C1406 VTAIL.n609 VSUBS 0.016159f
C1407 VTAIL.n610 VSUBS 0.01711f
C1408 VTAIL.n611 VSUBS 0.038195f
C1409 VTAIL.n612 VSUBS 0.038195f
C1410 VTAIL.n613 VSUBS 0.01711f
C1411 VTAIL.n614 VSUBS 0.016159f
C1412 VTAIL.n615 VSUBS 0.030072f
C1413 VTAIL.n616 VSUBS 0.030072f
C1414 VTAIL.n617 VSUBS 0.016159f
C1415 VTAIL.n618 VSUBS 0.01711f
C1416 VTAIL.n619 VSUBS 0.038195f
C1417 VTAIL.n620 VSUBS 0.038195f
C1418 VTAIL.n621 VSUBS 0.01711f
C1419 VTAIL.n622 VSUBS 0.016159f
C1420 VTAIL.n623 VSUBS 0.030072f
C1421 VTAIL.n624 VSUBS 0.030072f
C1422 VTAIL.n625 VSUBS 0.016159f
C1423 VTAIL.n626 VSUBS 0.01711f
C1424 VTAIL.n627 VSUBS 0.038195f
C1425 VTAIL.n628 VSUBS 0.038195f
C1426 VTAIL.n629 VSUBS 0.01711f
C1427 VTAIL.n630 VSUBS 0.016159f
C1428 VTAIL.n631 VSUBS 0.030072f
C1429 VTAIL.n632 VSUBS 0.030072f
C1430 VTAIL.n633 VSUBS 0.016159f
C1431 VTAIL.n634 VSUBS 0.01711f
C1432 VTAIL.n635 VSUBS 0.038195f
C1433 VTAIL.n636 VSUBS 0.038195f
C1434 VTAIL.n637 VSUBS 0.01711f
C1435 VTAIL.n638 VSUBS 0.016159f
C1436 VTAIL.n639 VSUBS 0.030072f
C1437 VTAIL.n640 VSUBS 0.030072f
C1438 VTAIL.n641 VSUBS 0.016159f
C1439 VTAIL.n642 VSUBS 0.01711f
C1440 VTAIL.n643 VSUBS 0.038195f
C1441 VTAIL.n644 VSUBS 0.038195f
C1442 VTAIL.n645 VSUBS 0.01711f
C1443 VTAIL.n646 VSUBS 0.016159f
C1444 VTAIL.n647 VSUBS 0.030072f
C1445 VTAIL.n648 VSUBS 0.030072f
C1446 VTAIL.n649 VSUBS 0.016159f
C1447 VTAIL.n650 VSUBS 0.01711f
C1448 VTAIL.n651 VSUBS 0.038195f
C1449 VTAIL.n652 VSUBS 0.038195f
C1450 VTAIL.n653 VSUBS 0.01711f
C1451 VTAIL.n654 VSUBS 0.016159f
C1452 VTAIL.n655 VSUBS 0.030072f
C1453 VTAIL.n656 VSUBS 0.030072f
C1454 VTAIL.n657 VSUBS 0.016159f
C1455 VTAIL.n658 VSUBS 0.01711f
C1456 VTAIL.n659 VSUBS 0.038195f
C1457 VTAIL.n660 VSUBS 0.092038f
C1458 VTAIL.n661 VSUBS 0.01711f
C1459 VTAIL.n662 VSUBS 0.016159f
C1460 VTAIL.n663 VSUBS 0.066224f
C1461 VTAIL.n664 VSUBS 0.046163f
C1462 VTAIL.n665 VSUBS 0.116136f
C1463 VTAIL.t2 VSUBS 0.465775f
C1464 VTAIL.t1 VSUBS 0.465775f
C1465 VTAIL.n666 VSUBS 3.69552f
C1466 VTAIL.n667 VSUBS 0.865601f
C1467 VTAIL.n668 VSUBS 0.032917f
C1468 VTAIL.n669 VSUBS 0.030072f
C1469 VTAIL.n670 VSUBS 0.016159f
C1470 VTAIL.n671 VSUBS 0.038195f
C1471 VTAIL.n672 VSUBS 0.01711f
C1472 VTAIL.n673 VSUBS 0.030072f
C1473 VTAIL.n674 VSUBS 0.016159f
C1474 VTAIL.n675 VSUBS 0.038195f
C1475 VTAIL.n676 VSUBS 0.01711f
C1476 VTAIL.n677 VSUBS 0.030072f
C1477 VTAIL.n678 VSUBS 0.016159f
C1478 VTAIL.n679 VSUBS 0.038195f
C1479 VTAIL.n680 VSUBS 0.016635f
C1480 VTAIL.n681 VSUBS 0.030072f
C1481 VTAIL.n682 VSUBS 0.016635f
C1482 VTAIL.n683 VSUBS 0.016159f
C1483 VTAIL.n684 VSUBS 0.038195f
C1484 VTAIL.n685 VSUBS 0.038195f
C1485 VTAIL.n686 VSUBS 0.01711f
C1486 VTAIL.n687 VSUBS 0.030072f
C1487 VTAIL.n688 VSUBS 0.016159f
C1488 VTAIL.n689 VSUBS 0.038195f
C1489 VTAIL.n690 VSUBS 0.01711f
C1490 VTAIL.n691 VSUBS 0.030072f
C1491 VTAIL.n692 VSUBS 0.016159f
C1492 VTAIL.n693 VSUBS 0.038195f
C1493 VTAIL.n694 VSUBS 0.01711f
C1494 VTAIL.n695 VSUBS 0.030072f
C1495 VTAIL.n696 VSUBS 0.016159f
C1496 VTAIL.n697 VSUBS 0.038195f
C1497 VTAIL.n698 VSUBS 0.01711f
C1498 VTAIL.n699 VSUBS 0.030072f
C1499 VTAIL.n700 VSUBS 0.016159f
C1500 VTAIL.n701 VSUBS 0.038195f
C1501 VTAIL.n702 VSUBS 0.01711f
C1502 VTAIL.n703 VSUBS 2.54816f
C1503 VTAIL.n704 VSUBS 0.016159f
C1504 VTAIL.t3 VSUBS 0.082112f
C1505 VTAIL.n705 VSUBS 0.252786f
C1506 VTAIL.n706 VSUBS 0.024298f
C1507 VTAIL.n707 VSUBS 0.028646f
C1508 VTAIL.n708 VSUBS 0.038195f
C1509 VTAIL.n709 VSUBS 0.01711f
C1510 VTAIL.n710 VSUBS 0.016159f
C1511 VTAIL.n711 VSUBS 0.030072f
C1512 VTAIL.n712 VSUBS 0.030072f
C1513 VTAIL.n713 VSUBS 0.016159f
C1514 VTAIL.n714 VSUBS 0.01711f
C1515 VTAIL.n715 VSUBS 0.038195f
C1516 VTAIL.n716 VSUBS 0.038195f
C1517 VTAIL.n717 VSUBS 0.01711f
C1518 VTAIL.n718 VSUBS 0.016159f
C1519 VTAIL.n719 VSUBS 0.030072f
C1520 VTAIL.n720 VSUBS 0.030072f
C1521 VTAIL.n721 VSUBS 0.016159f
C1522 VTAIL.n722 VSUBS 0.01711f
C1523 VTAIL.n723 VSUBS 0.038195f
C1524 VTAIL.n724 VSUBS 0.038195f
C1525 VTAIL.n725 VSUBS 0.01711f
C1526 VTAIL.n726 VSUBS 0.016159f
C1527 VTAIL.n727 VSUBS 0.030072f
C1528 VTAIL.n728 VSUBS 0.030072f
C1529 VTAIL.n729 VSUBS 0.016159f
C1530 VTAIL.n730 VSUBS 0.01711f
C1531 VTAIL.n731 VSUBS 0.038195f
C1532 VTAIL.n732 VSUBS 0.038195f
C1533 VTAIL.n733 VSUBS 0.01711f
C1534 VTAIL.n734 VSUBS 0.016159f
C1535 VTAIL.n735 VSUBS 0.030072f
C1536 VTAIL.n736 VSUBS 0.030072f
C1537 VTAIL.n737 VSUBS 0.016159f
C1538 VTAIL.n738 VSUBS 0.01711f
C1539 VTAIL.n739 VSUBS 0.038195f
C1540 VTAIL.n740 VSUBS 0.038195f
C1541 VTAIL.n741 VSUBS 0.01711f
C1542 VTAIL.n742 VSUBS 0.016159f
C1543 VTAIL.n743 VSUBS 0.030072f
C1544 VTAIL.n744 VSUBS 0.030072f
C1545 VTAIL.n745 VSUBS 0.016159f
C1546 VTAIL.n746 VSUBS 0.01711f
C1547 VTAIL.n747 VSUBS 0.038195f
C1548 VTAIL.n748 VSUBS 0.038195f
C1549 VTAIL.n749 VSUBS 0.01711f
C1550 VTAIL.n750 VSUBS 0.016159f
C1551 VTAIL.n751 VSUBS 0.030072f
C1552 VTAIL.n752 VSUBS 0.030072f
C1553 VTAIL.n753 VSUBS 0.016159f
C1554 VTAIL.n754 VSUBS 0.01711f
C1555 VTAIL.n755 VSUBS 0.038195f
C1556 VTAIL.n756 VSUBS 0.038195f
C1557 VTAIL.n757 VSUBS 0.01711f
C1558 VTAIL.n758 VSUBS 0.016159f
C1559 VTAIL.n759 VSUBS 0.030072f
C1560 VTAIL.n760 VSUBS 0.030072f
C1561 VTAIL.n761 VSUBS 0.016159f
C1562 VTAIL.n762 VSUBS 0.01711f
C1563 VTAIL.n763 VSUBS 0.038195f
C1564 VTAIL.n764 VSUBS 0.038195f
C1565 VTAIL.n765 VSUBS 0.01711f
C1566 VTAIL.n766 VSUBS 0.016159f
C1567 VTAIL.n767 VSUBS 0.030072f
C1568 VTAIL.n768 VSUBS 0.030072f
C1569 VTAIL.n769 VSUBS 0.016159f
C1570 VTAIL.n770 VSUBS 0.01711f
C1571 VTAIL.n771 VSUBS 0.038195f
C1572 VTAIL.n772 VSUBS 0.092038f
C1573 VTAIL.n773 VSUBS 0.01711f
C1574 VTAIL.n774 VSUBS 0.016159f
C1575 VTAIL.n775 VSUBS 0.066224f
C1576 VTAIL.n776 VSUBS 0.046163f
C1577 VTAIL.n777 VSUBS 2.16315f
C1578 VTAIL.n778 VSUBS 0.032917f
C1579 VTAIL.n779 VSUBS 0.030072f
C1580 VTAIL.n780 VSUBS 0.016159f
C1581 VTAIL.n781 VSUBS 0.038195f
C1582 VTAIL.n782 VSUBS 0.01711f
C1583 VTAIL.n783 VSUBS 0.030072f
C1584 VTAIL.n784 VSUBS 0.016159f
C1585 VTAIL.n785 VSUBS 0.038195f
C1586 VTAIL.n786 VSUBS 0.01711f
C1587 VTAIL.n787 VSUBS 0.030072f
C1588 VTAIL.n788 VSUBS 0.016159f
C1589 VTAIL.n789 VSUBS 0.038195f
C1590 VTAIL.n790 VSUBS 0.016635f
C1591 VTAIL.n791 VSUBS 0.030072f
C1592 VTAIL.n792 VSUBS 0.01711f
C1593 VTAIL.n793 VSUBS 0.038195f
C1594 VTAIL.n794 VSUBS 0.01711f
C1595 VTAIL.n795 VSUBS 0.030072f
C1596 VTAIL.n796 VSUBS 0.016159f
C1597 VTAIL.n797 VSUBS 0.038195f
C1598 VTAIL.n798 VSUBS 0.01711f
C1599 VTAIL.n799 VSUBS 0.030072f
C1600 VTAIL.n800 VSUBS 0.016159f
C1601 VTAIL.n801 VSUBS 0.038195f
C1602 VTAIL.n802 VSUBS 0.01711f
C1603 VTAIL.n803 VSUBS 0.030072f
C1604 VTAIL.n804 VSUBS 0.016159f
C1605 VTAIL.n805 VSUBS 0.038195f
C1606 VTAIL.n806 VSUBS 0.01711f
C1607 VTAIL.n807 VSUBS 0.030072f
C1608 VTAIL.n808 VSUBS 0.016159f
C1609 VTAIL.n809 VSUBS 0.038195f
C1610 VTAIL.n810 VSUBS 0.01711f
C1611 VTAIL.n811 VSUBS 2.54817f
C1612 VTAIL.n812 VSUBS 0.016159f
C1613 VTAIL.t10 VSUBS 0.082112f
C1614 VTAIL.n813 VSUBS 0.252786f
C1615 VTAIL.n814 VSUBS 0.024298f
C1616 VTAIL.n815 VSUBS 0.028646f
C1617 VTAIL.n816 VSUBS 0.038195f
C1618 VTAIL.n817 VSUBS 0.01711f
C1619 VTAIL.n818 VSUBS 0.016159f
C1620 VTAIL.n819 VSUBS 0.030072f
C1621 VTAIL.n820 VSUBS 0.030072f
C1622 VTAIL.n821 VSUBS 0.016159f
C1623 VTAIL.n822 VSUBS 0.01711f
C1624 VTAIL.n823 VSUBS 0.038195f
C1625 VTAIL.n824 VSUBS 0.038195f
C1626 VTAIL.n825 VSUBS 0.01711f
C1627 VTAIL.n826 VSUBS 0.016159f
C1628 VTAIL.n827 VSUBS 0.030072f
C1629 VTAIL.n828 VSUBS 0.030072f
C1630 VTAIL.n829 VSUBS 0.016159f
C1631 VTAIL.n830 VSUBS 0.01711f
C1632 VTAIL.n831 VSUBS 0.038195f
C1633 VTAIL.n832 VSUBS 0.038195f
C1634 VTAIL.n833 VSUBS 0.01711f
C1635 VTAIL.n834 VSUBS 0.016159f
C1636 VTAIL.n835 VSUBS 0.030072f
C1637 VTAIL.n836 VSUBS 0.030072f
C1638 VTAIL.n837 VSUBS 0.016159f
C1639 VTAIL.n838 VSUBS 0.01711f
C1640 VTAIL.n839 VSUBS 0.038195f
C1641 VTAIL.n840 VSUBS 0.038195f
C1642 VTAIL.n841 VSUBS 0.01711f
C1643 VTAIL.n842 VSUBS 0.016159f
C1644 VTAIL.n843 VSUBS 0.030072f
C1645 VTAIL.n844 VSUBS 0.030072f
C1646 VTAIL.n845 VSUBS 0.016159f
C1647 VTAIL.n846 VSUBS 0.01711f
C1648 VTAIL.n847 VSUBS 0.038195f
C1649 VTAIL.n848 VSUBS 0.038195f
C1650 VTAIL.n849 VSUBS 0.01711f
C1651 VTAIL.n850 VSUBS 0.016159f
C1652 VTAIL.n851 VSUBS 0.030072f
C1653 VTAIL.n852 VSUBS 0.030072f
C1654 VTAIL.n853 VSUBS 0.016159f
C1655 VTAIL.n854 VSUBS 0.016159f
C1656 VTAIL.n855 VSUBS 0.01711f
C1657 VTAIL.n856 VSUBS 0.038195f
C1658 VTAIL.n857 VSUBS 0.038195f
C1659 VTAIL.n858 VSUBS 0.038195f
C1660 VTAIL.n859 VSUBS 0.016635f
C1661 VTAIL.n860 VSUBS 0.016159f
C1662 VTAIL.n861 VSUBS 0.030072f
C1663 VTAIL.n862 VSUBS 0.030072f
C1664 VTAIL.n863 VSUBS 0.016159f
C1665 VTAIL.n864 VSUBS 0.01711f
C1666 VTAIL.n865 VSUBS 0.038195f
C1667 VTAIL.n866 VSUBS 0.038195f
C1668 VTAIL.n867 VSUBS 0.01711f
C1669 VTAIL.n868 VSUBS 0.016159f
C1670 VTAIL.n869 VSUBS 0.030072f
C1671 VTAIL.n870 VSUBS 0.030072f
C1672 VTAIL.n871 VSUBS 0.016159f
C1673 VTAIL.n872 VSUBS 0.01711f
C1674 VTAIL.n873 VSUBS 0.038195f
C1675 VTAIL.n874 VSUBS 0.038195f
C1676 VTAIL.n875 VSUBS 0.01711f
C1677 VTAIL.n876 VSUBS 0.016159f
C1678 VTAIL.n877 VSUBS 0.030072f
C1679 VTAIL.n878 VSUBS 0.030072f
C1680 VTAIL.n879 VSUBS 0.016159f
C1681 VTAIL.n880 VSUBS 0.01711f
C1682 VTAIL.n881 VSUBS 0.038195f
C1683 VTAIL.n882 VSUBS 0.092038f
C1684 VTAIL.n883 VSUBS 0.01711f
C1685 VTAIL.n884 VSUBS 0.016159f
C1686 VTAIL.n885 VSUBS 0.066224f
C1687 VTAIL.n886 VSUBS 0.046163f
C1688 VTAIL.n887 VSUBS 2.15751f
C1689 VN.n0 VSUBS 0.155224f
C1690 VN.t1 VSUBS 0.875797f
C1691 VN.t7 VSUBS 0.875797f
C1692 VN.t6 VSUBS 0.883199f
C1693 VN.n1 VSUBS 0.352259f
C1694 VN.n2 VSUBS 0.331161f
C1695 VN.n3 VSUBS 0.025423f
C1696 VN.n4 VSUBS 0.331161f
C1697 VN.t2 VSUBS 0.883199f
C1698 VN.n5 VSUBS 0.352158f
C1699 VN.n6 VSUBS 0.053432f
C1700 VN.n7 VSUBS 0.155224f
C1701 VN.t5 VSUBS 0.883199f
C1702 VN.t0 VSUBS 0.875797f
C1703 VN.t3 VSUBS 0.875797f
C1704 VN.t4 VSUBS 0.883199f
C1705 VN.n8 VSUBS 0.352259f
C1706 VN.n9 VSUBS 0.331161f
C1707 VN.n10 VSUBS 0.025423f
C1708 VN.n11 VSUBS 0.331161f
C1709 VN.n12 VSUBS 0.352158f
C1710 VN.n13 VSUBS 3.30414f
.ends

