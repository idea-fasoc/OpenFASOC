* NGSPICE file created from diff_pair_sample_1674.ext - technology: sky130A

.subckt diff_pair_sample_1674 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0 ps=0 w=5.18 l=1.09
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=0.8547 pd=5.51 as=2.0202 ps=11.14 w=5.18 l=1.09
X2 VTAIL.t6 VP.t1 VDD1.t2 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0.8547 ps=5.51 w=5.18 l=1.09
X3 VDD1.t1 VP.t2 VTAIL.t5 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=0.8547 pd=5.51 as=2.0202 ps=11.14 w=5.18 l=1.09
X4 B.t8 B.t6 B.t7 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0 ps=0 w=5.18 l=1.09
X5 VDD2.t3 VN.t0 VTAIL.t1 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=0.8547 pd=5.51 as=2.0202 ps=11.14 w=5.18 l=1.09
X6 VDD2.t2 VN.t1 VTAIL.t2 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=0.8547 pd=5.51 as=2.0202 ps=11.14 w=5.18 l=1.09
X7 VTAIL.t3 VN.t2 VDD2.t1 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0.8547 ps=5.51 w=5.18 l=1.09
X8 B.t5 B.t3 B.t4 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0 ps=0 w=5.18 l=1.09
X9 VTAIL.t0 VN.t3 VDD2.t0 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0.8547 ps=5.51 w=5.18 l=1.09
X10 VTAIL.t4 VP.t3 VDD1.t0 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0.8547 ps=5.51 w=5.18 l=1.09
X11 B.t2 B.t0 B.t1 w_n1822_n2004# sky130_fd_pr__pfet_01v8 ad=2.0202 pd=11.14 as=0 ps=0 w=5.18 l=1.09
R0 B.n213 B.n212 585
R1 B.n211 B.n64 585
R2 B.n210 B.n209 585
R3 B.n208 B.n65 585
R4 B.n207 B.n206 585
R5 B.n205 B.n66 585
R6 B.n204 B.n203 585
R7 B.n202 B.n67 585
R8 B.n201 B.n200 585
R9 B.n199 B.n68 585
R10 B.n198 B.n197 585
R11 B.n196 B.n69 585
R12 B.n195 B.n194 585
R13 B.n193 B.n70 585
R14 B.n192 B.n191 585
R15 B.n190 B.n71 585
R16 B.n189 B.n188 585
R17 B.n187 B.n72 585
R18 B.n186 B.n185 585
R19 B.n184 B.n73 585
R20 B.n183 B.n182 585
R21 B.n181 B.n74 585
R22 B.n180 B.n179 585
R23 B.n175 B.n75 585
R24 B.n174 B.n173 585
R25 B.n172 B.n76 585
R26 B.n171 B.n170 585
R27 B.n169 B.n77 585
R28 B.n168 B.n167 585
R29 B.n166 B.n78 585
R30 B.n165 B.n164 585
R31 B.n162 B.n79 585
R32 B.n161 B.n160 585
R33 B.n159 B.n82 585
R34 B.n158 B.n157 585
R35 B.n156 B.n83 585
R36 B.n155 B.n154 585
R37 B.n153 B.n84 585
R38 B.n152 B.n151 585
R39 B.n150 B.n85 585
R40 B.n149 B.n148 585
R41 B.n147 B.n86 585
R42 B.n146 B.n145 585
R43 B.n144 B.n87 585
R44 B.n143 B.n142 585
R45 B.n141 B.n88 585
R46 B.n140 B.n139 585
R47 B.n138 B.n89 585
R48 B.n137 B.n136 585
R49 B.n135 B.n90 585
R50 B.n134 B.n133 585
R51 B.n132 B.n91 585
R52 B.n131 B.n130 585
R53 B.n214 B.n63 585
R54 B.n216 B.n215 585
R55 B.n217 B.n62 585
R56 B.n219 B.n218 585
R57 B.n220 B.n61 585
R58 B.n222 B.n221 585
R59 B.n223 B.n60 585
R60 B.n225 B.n224 585
R61 B.n226 B.n59 585
R62 B.n228 B.n227 585
R63 B.n229 B.n58 585
R64 B.n231 B.n230 585
R65 B.n232 B.n57 585
R66 B.n234 B.n233 585
R67 B.n235 B.n56 585
R68 B.n237 B.n236 585
R69 B.n238 B.n55 585
R70 B.n240 B.n239 585
R71 B.n241 B.n54 585
R72 B.n243 B.n242 585
R73 B.n244 B.n53 585
R74 B.n246 B.n245 585
R75 B.n247 B.n52 585
R76 B.n249 B.n248 585
R77 B.n250 B.n51 585
R78 B.n252 B.n251 585
R79 B.n253 B.n50 585
R80 B.n255 B.n254 585
R81 B.n256 B.n49 585
R82 B.n258 B.n257 585
R83 B.n259 B.n48 585
R84 B.n261 B.n260 585
R85 B.n262 B.n47 585
R86 B.n264 B.n263 585
R87 B.n265 B.n46 585
R88 B.n267 B.n266 585
R89 B.n268 B.n45 585
R90 B.n270 B.n269 585
R91 B.n271 B.n44 585
R92 B.n273 B.n272 585
R93 B.n274 B.n43 585
R94 B.n276 B.n275 585
R95 B.n357 B.n12 585
R96 B.n356 B.n355 585
R97 B.n354 B.n13 585
R98 B.n353 B.n352 585
R99 B.n351 B.n14 585
R100 B.n350 B.n349 585
R101 B.n348 B.n15 585
R102 B.n347 B.n346 585
R103 B.n345 B.n16 585
R104 B.n344 B.n343 585
R105 B.n342 B.n17 585
R106 B.n341 B.n340 585
R107 B.n339 B.n18 585
R108 B.n338 B.n337 585
R109 B.n336 B.n19 585
R110 B.n335 B.n334 585
R111 B.n333 B.n20 585
R112 B.n332 B.n331 585
R113 B.n330 B.n21 585
R114 B.n329 B.n328 585
R115 B.n327 B.n22 585
R116 B.n326 B.n325 585
R117 B.n323 B.n23 585
R118 B.n322 B.n321 585
R119 B.n320 B.n26 585
R120 B.n319 B.n318 585
R121 B.n317 B.n27 585
R122 B.n316 B.n315 585
R123 B.n314 B.n28 585
R124 B.n313 B.n312 585
R125 B.n311 B.n29 585
R126 B.n309 B.n308 585
R127 B.n307 B.n32 585
R128 B.n306 B.n305 585
R129 B.n304 B.n33 585
R130 B.n303 B.n302 585
R131 B.n301 B.n34 585
R132 B.n300 B.n299 585
R133 B.n298 B.n35 585
R134 B.n297 B.n296 585
R135 B.n295 B.n36 585
R136 B.n294 B.n293 585
R137 B.n292 B.n37 585
R138 B.n291 B.n290 585
R139 B.n289 B.n38 585
R140 B.n288 B.n287 585
R141 B.n286 B.n39 585
R142 B.n285 B.n284 585
R143 B.n283 B.n40 585
R144 B.n282 B.n281 585
R145 B.n280 B.n41 585
R146 B.n279 B.n278 585
R147 B.n277 B.n42 585
R148 B.n359 B.n358 585
R149 B.n360 B.n11 585
R150 B.n362 B.n361 585
R151 B.n363 B.n10 585
R152 B.n365 B.n364 585
R153 B.n366 B.n9 585
R154 B.n368 B.n367 585
R155 B.n369 B.n8 585
R156 B.n371 B.n370 585
R157 B.n372 B.n7 585
R158 B.n374 B.n373 585
R159 B.n375 B.n6 585
R160 B.n377 B.n376 585
R161 B.n378 B.n5 585
R162 B.n380 B.n379 585
R163 B.n381 B.n4 585
R164 B.n383 B.n382 585
R165 B.n384 B.n3 585
R166 B.n386 B.n385 585
R167 B.n387 B.n0 585
R168 B.n2 B.n1 585
R169 B.n102 B.n101 585
R170 B.n104 B.n103 585
R171 B.n105 B.n100 585
R172 B.n107 B.n106 585
R173 B.n108 B.n99 585
R174 B.n110 B.n109 585
R175 B.n111 B.n98 585
R176 B.n113 B.n112 585
R177 B.n114 B.n97 585
R178 B.n116 B.n115 585
R179 B.n117 B.n96 585
R180 B.n119 B.n118 585
R181 B.n120 B.n95 585
R182 B.n122 B.n121 585
R183 B.n123 B.n94 585
R184 B.n125 B.n124 585
R185 B.n126 B.n93 585
R186 B.n128 B.n127 585
R187 B.n129 B.n92 585
R188 B.n130 B.n129 497.305
R189 B.n212 B.n63 497.305
R190 B.n277 B.n276 497.305
R191 B.n358 B.n357 497.305
R192 B.n80 B.t0 318.031
R193 B.n176 B.t6 318.031
R194 B.n30 B.t9 318.031
R195 B.n24 B.t3 318.031
R196 B.n176 B.t7 281.248
R197 B.n30 B.t11 281.248
R198 B.n80 B.t1 281.248
R199 B.n24 B.t5 281.248
R200 B.n389 B.n388 256.663
R201 B.n177 B.t8 253.708
R202 B.n31 B.t10 253.708
R203 B.n81 B.t2 253.708
R204 B.n25 B.t4 253.708
R205 B.n388 B.n387 235.042
R206 B.n388 B.n2 235.042
R207 B.n130 B.n91 163.367
R208 B.n134 B.n91 163.367
R209 B.n135 B.n134 163.367
R210 B.n136 B.n135 163.367
R211 B.n136 B.n89 163.367
R212 B.n140 B.n89 163.367
R213 B.n141 B.n140 163.367
R214 B.n142 B.n141 163.367
R215 B.n142 B.n87 163.367
R216 B.n146 B.n87 163.367
R217 B.n147 B.n146 163.367
R218 B.n148 B.n147 163.367
R219 B.n148 B.n85 163.367
R220 B.n152 B.n85 163.367
R221 B.n153 B.n152 163.367
R222 B.n154 B.n153 163.367
R223 B.n154 B.n83 163.367
R224 B.n158 B.n83 163.367
R225 B.n159 B.n158 163.367
R226 B.n160 B.n159 163.367
R227 B.n160 B.n79 163.367
R228 B.n165 B.n79 163.367
R229 B.n166 B.n165 163.367
R230 B.n167 B.n166 163.367
R231 B.n167 B.n77 163.367
R232 B.n171 B.n77 163.367
R233 B.n172 B.n171 163.367
R234 B.n173 B.n172 163.367
R235 B.n173 B.n75 163.367
R236 B.n180 B.n75 163.367
R237 B.n181 B.n180 163.367
R238 B.n182 B.n181 163.367
R239 B.n182 B.n73 163.367
R240 B.n186 B.n73 163.367
R241 B.n187 B.n186 163.367
R242 B.n188 B.n187 163.367
R243 B.n188 B.n71 163.367
R244 B.n192 B.n71 163.367
R245 B.n193 B.n192 163.367
R246 B.n194 B.n193 163.367
R247 B.n194 B.n69 163.367
R248 B.n198 B.n69 163.367
R249 B.n199 B.n198 163.367
R250 B.n200 B.n199 163.367
R251 B.n200 B.n67 163.367
R252 B.n204 B.n67 163.367
R253 B.n205 B.n204 163.367
R254 B.n206 B.n205 163.367
R255 B.n206 B.n65 163.367
R256 B.n210 B.n65 163.367
R257 B.n211 B.n210 163.367
R258 B.n212 B.n211 163.367
R259 B.n276 B.n43 163.367
R260 B.n272 B.n43 163.367
R261 B.n272 B.n271 163.367
R262 B.n271 B.n270 163.367
R263 B.n270 B.n45 163.367
R264 B.n266 B.n45 163.367
R265 B.n266 B.n265 163.367
R266 B.n265 B.n264 163.367
R267 B.n264 B.n47 163.367
R268 B.n260 B.n47 163.367
R269 B.n260 B.n259 163.367
R270 B.n259 B.n258 163.367
R271 B.n258 B.n49 163.367
R272 B.n254 B.n49 163.367
R273 B.n254 B.n253 163.367
R274 B.n253 B.n252 163.367
R275 B.n252 B.n51 163.367
R276 B.n248 B.n51 163.367
R277 B.n248 B.n247 163.367
R278 B.n247 B.n246 163.367
R279 B.n246 B.n53 163.367
R280 B.n242 B.n53 163.367
R281 B.n242 B.n241 163.367
R282 B.n241 B.n240 163.367
R283 B.n240 B.n55 163.367
R284 B.n236 B.n55 163.367
R285 B.n236 B.n235 163.367
R286 B.n235 B.n234 163.367
R287 B.n234 B.n57 163.367
R288 B.n230 B.n57 163.367
R289 B.n230 B.n229 163.367
R290 B.n229 B.n228 163.367
R291 B.n228 B.n59 163.367
R292 B.n224 B.n59 163.367
R293 B.n224 B.n223 163.367
R294 B.n223 B.n222 163.367
R295 B.n222 B.n61 163.367
R296 B.n218 B.n61 163.367
R297 B.n218 B.n217 163.367
R298 B.n217 B.n216 163.367
R299 B.n216 B.n63 163.367
R300 B.n357 B.n356 163.367
R301 B.n356 B.n13 163.367
R302 B.n352 B.n13 163.367
R303 B.n352 B.n351 163.367
R304 B.n351 B.n350 163.367
R305 B.n350 B.n15 163.367
R306 B.n346 B.n15 163.367
R307 B.n346 B.n345 163.367
R308 B.n345 B.n344 163.367
R309 B.n344 B.n17 163.367
R310 B.n340 B.n17 163.367
R311 B.n340 B.n339 163.367
R312 B.n339 B.n338 163.367
R313 B.n338 B.n19 163.367
R314 B.n334 B.n19 163.367
R315 B.n334 B.n333 163.367
R316 B.n333 B.n332 163.367
R317 B.n332 B.n21 163.367
R318 B.n328 B.n21 163.367
R319 B.n328 B.n327 163.367
R320 B.n327 B.n326 163.367
R321 B.n326 B.n23 163.367
R322 B.n321 B.n23 163.367
R323 B.n321 B.n320 163.367
R324 B.n320 B.n319 163.367
R325 B.n319 B.n27 163.367
R326 B.n315 B.n27 163.367
R327 B.n315 B.n314 163.367
R328 B.n314 B.n313 163.367
R329 B.n313 B.n29 163.367
R330 B.n308 B.n29 163.367
R331 B.n308 B.n307 163.367
R332 B.n307 B.n306 163.367
R333 B.n306 B.n33 163.367
R334 B.n302 B.n33 163.367
R335 B.n302 B.n301 163.367
R336 B.n301 B.n300 163.367
R337 B.n300 B.n35 163.367
R338 B.n296 B.n35 163.367
R339 B.n296 B.n295 163.367
R340 B.n295 B.n294 163.367
R341 B.n294 B.n37 163.367
R342 B.n290 B.n37 163.367
R343 B.n290 B.n289 163.367
R344 B.n289 B.n288 163.367
R345 B.n288 B.n39 163.367
R346 B.n284 B.n39 163.367
R347 B.n284 B.n283 163.367
R348 B.n283 B.n282 163.367
R349 B.n282 B.n41 163.367
R350 B.n278 B.n41 163.367
R351 B.n278 B.n277 163.367
R352 B.n358 B.n11 163.367
R353 B.n362 B.n11 163.367
R354 B.n363 B.n362 163.367
R355 B.n364 B.n363 163.367
R356 B.n364 B.n9 163.367
R357 B.n368 B.n9 163.367
R358 B.n369 B.n368 163.367
R359 B.n370 B.n369 163.367
R360 B.n370 B.n7 163.367
R361 B.n374 B.n7 163.367
R362 B.n375 B.n374 163.367
R363 B.n376 B.n375 163.367
R364 B.n376 B.n5 163.367
R365 B.n380 B.n5 163.367
R366 B.n381 B.n380 163.367
R367 B.n382 B.n381 163.367
R368 B.n382 B.n3 163.367
R369 B.n386 B.n3 163.367
R370 B.n387 B.n386 163.367
R371 B.n101 B.n2 163.367
R372 B.n104 B.n101 163.367
R373 B.n105 B.n104 163.367
R374 B.n106 B.n105 163.367
R375 B.n106 B.n99 163.367
R376 B.n110 B.n99 163.367
R377 B.n111 B.n110 163.367
R378 B.n112 B.n111 163.367
R379 B.n112 B.n97 163.367
R380 B.n116 B.n97 163.367
R381 B.n117 B.n116 163.367
R382 B.n118 B.n117 163.367
R383 B.n118 B.n95 163.367
R384 B.n122 B.n95 163.367
R385 B.n123 B.n122 163.367
R386 B.n124 B.n123 163.367
R387 B.n124 B.n93 163.367
R388 B.n128 B.n93 163.367
R389 B.n129 B.n128 163.367
R390 B.n163 B.n81 59.5399
R391 B.n178 B.n177 59.5399
R392 B.n310 B.n31 59.5399
R393 B.n324 B.n25 59.5399
R394 B.n359 B.n12 32.3127
R395 B.n275 B.n42 32.3127
R396 B.n214 B.n213 32.3127
R397 B.n131 B.n92 32.3127
R398 B.n81 B.n80 27.5399
R399 B.n177 B.n176 27.5399
R400 B.n31 B.n30 27.5399
R401 B.n25 B.n24 27.5399
R402 B B.n389 18.0485
R403 B.n360 B.n359 10.6151
R404 B.n361 B.n360 10.6151
R405 B.n361 B.n10 10.6151
R406 B.n365 B.n10 10.6151
R407 B.n366 B.n365 10.6151
R408 B.n367 B.n366 10.6151
R409 B.n367 B.n8 10.6151
R410 B.n371 B.n8 10.6151
R411 B.n372 B.n371 10.6151
R412 B.n373 B.n372 10.6151
R413 B.n373 B.n6 10.6151
R414 B.n377 B.n6 10.6151
R415 B.n378 B.n377 10.6151
R416 B.n379 B.n378 10.6151
R417 B.n379 B.n4 10.6151
R418 B.n383 B.n4 10.6151
R419 B.n384 B.n383 10.6151
R420 B.n385 B.n384 10.6151
R421 B.n385 B.n0 10.6151
R422 B.n355 B.n12 10.6151
R423 B.n355 B.n354 10.6151
R424 B.n354 B.n353 10.6151
R425 B.n353 B.n14 10.6151
R426 B.n349 B.n14 10.6151
R427 B.n349 B.n348 10.6151
R428 B.n348 B.n347 10.6151
R429 B.n347 B.n16 10.6151
R430 B.n343 B.n16 10.6151
R431 B.n343 B.n342 10.6151
R432 B.n342 B.n341 10.6151
R433 B.n341 B.n18 10.6151
R434 B.n337 B.n18 10.6151
R435 B.n337 B.n336 10.6151
R436 B.n336 B.n335 10.6151
R437 B.n335 B.n20 10.6151
R438 B.n331 B.n20 10.6151
R439 B.n331 B.n330 10.6151
R440 B.n330 B.n329 10.6151
R441 B.n329 B.n22 10.6151
R442 B.n325 B.n22 10.6151
R443 B.n323 B.n322 10.6151
R444 B.n322 B.n26 10.6151
R445 B.n318 B.n26 10.6151
R446 B.n318 B.n317 10.6151
R447 B.n317 B.n316 10.6151
R448 B.n316 B.n28 10.6151
R449 B.n312 B.n28 10.6151
R450 B.n312 B.n311 10.6151
R451 B.n309 B.n32 10.6151
R452 B.n305 B.n32 10.6151
R453 B.n305 B.n304 10.6151
R454 B.n304 B.n303 10.6151
R455 B.n303 B.n34 10.6151
R456 B.n299 B.n34 10.6151
R457 B.n299 B.n298 10.6151
R458 B.n298 B.n297 10.6151
R459 B.n297 B.n36 10.6151
R460 B.n293 B.n36 10.6151
R461 B.n293 B.n292 10.6151
R462 B.n292 B.n291 10.6151
R463 B.n291 B.n38 10.6151
R464 B.n287 B.n38 10.6151
R465 B.n287 B.n286 10.6151
R466 B.n286 B.n285 10.6151
R467 B.n285 B.n40 10.6151
R468 B.n281 B.n40 10.6151
R469 B.n281 B.n280 10.6151
R470 B.n280 B.n279 10.6151
R471 B.n279 B.n42 10.6151
R472 B.n275 B.n274 10.6151
R473 B.n274 B.n273 10.6151
R474 B.n273 B.n44 10.6151
R475 B.n269 B.n44 10.6151
R476 B.n269 B.n268 10.6151
R477 B.n268 B.n267 10.6151
R478 B.n267 B.n46 10.6151
R479 B.n263 B.n46 10.6151
R480 B.n263 B.n262 10.6151
R481 B.n262 B.n261 10.6151
R482 B.n261 B.n48 10.6151
R483 B.n257 B.n48 10.6151
R484 B.n257 B.n256 10.6151
R485 B.n256 B.n255 10.6151
R486 B.n255 B.n50 10.6151
R487 B.n251 B.n50 10.6151
R488 B.n251 B.n250 10.6151
R489 B.n250 B.n249 10.6151
R490 B.n249 B.n52 10.6151
R491 B.n245 B.n52 10.6151
R492 B.n245 B.n244 10.6151
R493 B.n244 B.n243 10.6151
R494 B.n243 B.n54 10.6151
R495 B.n239 B.n54 10.6151
R496 B.n239 B.n238 10.6151
R497 B.n238 B.n237 10.6151
R498 B.n237 B.n56 10.6151
R499 B.n233 B.n56 10.6151
R500 B.n233 B.n232 10.6151
R501 B.n232 B.n231 10.6151
R502 B.n231 B.n58 10.6151
R503 B.n227 B.n58 10.6151
R504 B.n227 B.n226 10.6151
R505 B.n226 B.n225 10.6151
R506 B.n225 B.n60 10.6151
R507 B.n221 B.n60 10.6151
R508 B.n221 B.n220 10.6151
R509 B.n220 B.n219 10.6151
R510 B.n219 B.n62 10.6151
R511 B.n215 B.n62 10.6151
R512 B.n215 B.n214 10.6151
R513 B.n102 B.n1 10.6151
R514 B.n103 B.n102 10.6151
R515 B.n103 B.n100 10.6151
R516 B.n107 B.n100 10.6151
R517 B.n108 B.n107 10.6151
R518 B.n109 B.n108 10.6151
R519 B.n109 B.n98 10.6151
R520 B.n113 B.n98 10.6151
R521 B.n114 B.n113 10.6151
R522 B.n115 B.n114 10.6151
R523 B.n115 B.n96 10.6151
R524 B.n119 B.n96 10.6151
R525 B.n120 B.n119 10.6151
R526 B.n121 B.n120 10.6151
R527 B.n121 B.n94 10.6151
R528 B.n125 B.n94 10.6151
R529 B.n126 B.n125 10.6151
R530 B.n127 B.n126 10.6151
R531 B.n127 B.n92 10.6151
R532 B.n132 B.n131 10.6151
R533 B.n133 B.n132 10.6151
R534 B.n133 B.n90 10.6151
R535 B.n137 B.n90 10.6151
R536 B.n138 B.n137 10.6151
R537 B.n139 B.n138 10.6151
R538 B.n139 B.n88 10.6151
R539 B.n143 B.n88 10.6151
R540 B.n144 B.n143 10.6151
R541 B.n145 B.n144 10.6151
R542 B.n145 B.n86 10.6151
R543 B.n149 B.n86 10.6151
R544 B.n150 B.n149 10.6151
R545 B.n151 B.n150 10.6151
R546 B.n151 B.n84 10.6151
R547 B.n155 B.n84 10.6151
R548 B.n156 B.n155 10.6151
R549 B.n157 B.n156 10.6151
R550 B.n157 B.n82 10.6151
R551 B.n161 B.n82 10.6151
R552 B.n162 B.n161 10.6151
R553 B.n164 B.n78 10.6151
R554 B.n168 B.n78 10.6151
R555 B.n169 B.n168 10.6151
R556 B.n170 B.n169 10.6151
R557 B.n170 B.n76 10.6151
R558 B.n174 B.n76 10.6151
R559 B.n175 B.n174 10.6151
R560 B.n179 B.n175 10.6151
R561 B.n183 B.n74 10.6151
R562 B.n184 B.n183 10.6151
R563 B.n185 B.n184 10.6151
R564 B.n185 B.n72 10.6151
R565 B.n189 B.n72 10.6151
R566 B.n190 B.n189 10.6151
R567 B.n191 B.n190 10.6151
R568 B.n191 B.n70 10.6151
R569 B.n195 B.n70 10.6151
R570 B.n196 B.n195 10.6151
R571 B.n197 B.n196 10.6151
R572 B.n197 B.n68 10.6151
R573 B.n201 B.n68 10.6151
R574 B.n202 B.n201 10.6151
R575 B.n203 B.n202 10.6151
R576 B.n203 B.n66 10.6151
R577 B.n207 B.n66 10.6151
R578 B.n208 B.n207 10.6151
R579 B.n209 B.n208 10.6151
R580 B.n209 B.n64 10.6151
R581 B.n213 B.n64 10.6151
R582 B.n389 B.n0 8.11757
R583 B.n389 B.n1 8.11757
R584 B.n324 B.n323 6.5566
R585 B.n311 B.n310 6.5566
R586 B.n164 B.n163 6.5566
R587 B.n179 B.n178 6.5566
R588 B.n325 B.n324 4.05904
R589 B.n310 B.n309 4.05904
R590 B.n163 B.n162 4.05904
R591 B.n178 B.n74 4.05904
R592 VP.n0 VP.t3 169.178
R593 VP.n0 VP.t2 169.089
R594 VP.n2 VP.t1 150.571
R595 VP.n3 VP.t0 150.571
R596 VP.n4 VP.n3 80.6037
R597 VP.n2 VP.n1 80.6037
R598 VP.n1 VP.n0 67.8365
R599 VP.n3 VP.n2 48.2005
R600 VP.n4 VP.n1 0.380177
R601 VP VP.n4 0.146778
R602 VTAIL.n218 VTAIL.n196 756.745
R603 VTAIL.n22 VTAIL.n0 756.745
R604 VTAIL.n50 VTAIL.n28 756.745
R605 VTAIL.n78 VTAIL.n56 756.745
R606 VTAIL.n190 VTAIL.n168 756.745
R607 VTAIL.n162 VTAIL.n140 756.745
R608 VTAIL.n134 VTAIL.n112 756.745
R609 VTAIL.n106 VTAIL.n84 756.745
R610 VTAIL.n204 VTAIL.n203 585
R611 VTAIL.n209 VTAIL.n208 585
R612 VTAIL.n211 VTAIL.n210 585
R613 VTAIL.n200 VTAIL.n199 585
R614 VTAIL.n217 VTAIL.n216 585
R615 VTAIL.n219 VTAIL.n218 585
R616 VTAIL.n8 VTAIL.n7 585
R617 VTAIL.n13 VTAIL.n12 585
R618 VTAIL.n15 VTAIL.n14 585
R619 VTAIL.n4 VTAIL.n3 585
R620 VTAIL.n21 VTAIL.n20 585
R621 VTAIL.n23 VTAIL.n22 585
R622 VTAIL.n36 VTAIL.n35 585
R623 VTAIL.n41 VTAIL.n40 585
R624 VTAIL.n43 VTAIL.n42 585
R625 VTAIL.n32 VTAIL.n31 585
R626 VTAIL.n49 VTAIL.n48 585
R627 VTAIL.n51 VTAIL.n50 585
R628 VTAIL.n64 VTAIL.n63 585
R629 VTAIL.n69 VTAIL.n68 585
R630 VTAIL.n71 VTAIL.n70 585
R631 VTAIL.n60 VTAIL.n59 585
R632 VTAIL.n77 VTAIL.n76 585
R633 VTAIL.n79 VTAIL.n78 585
R634 VTAIL.n191 VTAIL.n190 585
R635 VTAIL.n189 VTAIL.n188 585
R636 VTAIL.n172 VTAIL.n171 585
R637 VTAIL.n183 VTAIL.n182 585
R638 VTAIL.n181 VTAIL.n180 585
R639 VTAIL.n176 VTAIL.n175 585
R640 VTAIL.n163 VTAIL.n162 585
R641 VTAIL.n161 VTAIL.n160 585
R642 VTAIL.n144 VTAIL.n143 585
R643 VTAIL.n155 VTAIL.n154 585
R644 VTAIL.n153 VTAIL.n152 585
R645 VTAIL.n148 VTAIL.n147 585
R646 VTAIL.n135 VTAIL.n134 585
R647 VTAIL.n133 VTAIL.n132 585
R648 VTAIL.n116 VTAIL.n115 585
R649 VTAIL.n127 VTAIL.n126 585
R650 VTAIL.n125 VTAIL.n124 585
R651 VTAIL.n120 VTAIL.n119 585
R652 VTAIL.n107 VTAIL.n106 585
R653 VTAIL.n105 VTAIL.n104 585
R654 VTAIL.n88 VTAIL.n87 585
R655 VTAIL.n99 VTAIL.n98 585
R656 VTAIL.n97 VTAIL.n96 585
R657 VTAIL.n92 VTAIL.n91 585
R658 VTAIL.n205 VTAIL.t1 327.856
R659 VTAIL.n9 VTAIL.t3 327.856
R660 VTAIL.n37 VTAIL.t7 327.856
R661 VTAIL.n65 VTAIL.t6 327.856
R662 VTAIL.n177 VTAIL.t5 327.856
R663 VTAIL.n149 VTAIL.t4 327.856
R664 VTAIL.n121 VTAIL.t2 327.856
R665 VTAIL.n93 VTAIL.t0 327.856
R666 VTAIL.n209 VTAIL.n203 171.744
R667 VTAIL.n210 VTAIL.n209 171.744
R668 VTAIL.n210 VTAIL.n199 171.744
R669 VTAIL.n217 VTAIL.n199 171.744
R670 VTAIL.n218 VTAIL.n217 171.744
R671 VTAIL.n13 VTAIL.n7 171.744
R672 VTAIL.n14 VTAIL.n13 171.744
R673 VTAIL.n14 VTAIL.n3 171.744
R674 VTAIL.n21 VTAIL.n3 171.744
R675 VTAIL.n22 VTAIL.n21 171.744
R676 VTAIL.n41 VTAIL.n35 171.744
R677 VTAIL.n42 VTAIL.n41 171.744
R678 VTAIL.n42 VTAIL.n31 171.744
R679 VTAIL.n49 VTAIL.n31 171.744
R680 VTAIL.n50 VTAIL.n49 171.744
R681 VTAIL.n69 VTAIL.n63 171.744
R682 VTAIL.n70 VTAIL.n69 171.744
R683 VTAIL.n70 VTAIL.n59 171.744
R684 VTAIL.n77 VTAIL.n59 171.744
R685 VTAIL.n78 VTAIL.n77 171.744
R686 VTAIL.n190 VTAIL.n189 171.744
R687 VTAIL.n189 VTAIL.n171 171.744
R688 VTAIL.n182 VTAIL.n171 171.744
R689 VTAIL.n182 VTAIL.n181 171.744
R690 VTAIL.n181 VTAIL.n175 171.744
R691 VTAIL.n162 VTAIL.n161 171.744
R692 VTAIL.n161 VTAIL.n143 171.744
R693 VTAIL.n154 VTAIL.n143 171.744
R694 VTAIL.n154 VTAIL.n153 171.744
R695 VTAIL.n153 VTAIL.n147 171.744
R696 VTAIL.n134 VTAIL.n133 171.744
R697 VTAIL.n133 VTAIL.n115 171.744
R698 VTAIL.n126 VTAIL.n115 171.744
R699 VTAIL.n126 VTAIL.n125 171.744
R700 VTAIL.n125 VTAIL.n119 171.744
R701 VTAIL.n106 VTAIL.n105 171.744
R702 VTAIL.n105 VTAIL.n87 171.744
R703 VTAIL.n98 VTAIL.n87 171.744
R704 VTAIL.n98 VTAIL.n97 171.744
R705 VTAIL.n97 VTAIL.n91 171.744
R706 VTAIL.t1 VTAIL.n203 85.8723
R707 VTAIL.t3 VTAIL.n7 85.8723
R708 VTAIL.t7 VTAIL.n35 85.8723
R709 VTAIL.t6 VTAIL.n63 85.8723
R710 VTAIL.t5 VTAIL.n175 85.8723
R711 VTAIL.t4 VTAIL.n147 85.8723
R712 VTAIL.t2 VTAIL.n119 85.8723
R713 VTAIL.t0 VTAIL.n91 85.8723
R714 VTAIL.n223 VTAIL.n222 30.246
R715 VTAIL.n27 VTAIL.n26 30.246
R716 VTAIL.n55 VTAIL.n54 30.246
R717 VTAIL.n83 VTAIL.n82 30.246
R718 VTAIL.n195 VTAIL.n194 30.246
R719 VTAIL.n167 VTAIL.n166 30.246
R720 VTAIL.n139 VTAIL.n138 30.246
R721 VTAIL.n111 VTAIL.n110 30.246
R722 VTAIL.n223 VTAIL.n195 18.0565
R723 VTAIL.n111 VTAIL.n83 18.0565
R724 VTAIL.n205 VTAIL.n204 16.381
R725 VTAIL.n9 VTAIL.n8 16.381
R726 VTAIL.n37 VTAIL.n36 16.381
R727 VTAIL.n65 VTAIL.n64 16.381
R728 VTAIL.n177 VTAIL.n176 16.381
R729 VTAIL.n149 VTAIL.n148 16.381
R730 VTAIL.n121 VTAIL.n120 16.381
R731 VTAIL.n93 VTAIL.n92 16.381
R732 VTAIL.n208 VTAIL.n207 12.8005
R733 VTAIL.n12 VTAIL.n11 12.8005
R734 VTAIL.n40 VTAIL.n39 12.8005
R735 VTAIL.n68 VTAIL.n67 12.8005
R736 VTAIL.n180 VTAIL.n179 12.8005
R737 VTAIL.n152 VTAIL.n151 12.8005
R738 VTAIL.n124 VTAIL.n123 12.8005
R739 VTAIL.n96 VTAIL.n95 12.8005
R740 VTAIL.n211 VTAIL.n202 12.0247
R741 VTAIL.n15 VTAIL.n6 12.0247
R742 VTAIL.n43 VTAIL.n34 12.0247
R743 VTAIL.n71 VTAIL.n62 12.0247
R744 VTAIL.n183 VTAIL.n174 12.0247
R745 VTAIL.n155 VTAIL.n146 12.0247
R746 VTAIL.n127 VTAIL.n118 12.0247
R747 VTAIL.n99 VTAIL.n90 12.0247
R748 VTAIL.n212 VTAIL.n200 11.249
R749 VTAIL.n16 VTAIL.n4 11.249
R750 VTAIL.n44 VTAIL.n32 11.249
R751 VTAIL.n72 VTAIL.n60 11.249
R752 VTAIL.n184 VTAIL.n172 11.249
R753 VTAIL.n156 VTAIL.n144 11.249
R754 VTAIL.n128 VTAIL.n116 11.249
R755 VTAIL.n100 VTAIL.n88 11.249
R756 VTAIL.n216 VTAIL.n215 10.4732
R757 VTAIL.n20 VTAIL.n19 10.4732
R758 VTAIL.n48 VTAIL.n47 10.4732
R759 VTAIL.n76 VTAIL.n75 10.4732
R760 VTAIL.n188 VTAIL.n187 10.4732
R761 VTAIL.n160 VTAIL.n159 10.4732
R762 VTAIL.n132 VTAIL.n131 10.4732
R763 VTAIL.n104 VTAIL.n103 10.4732
R764 VTAIL.n219 VTAIL.n198 9.69747
R765 VTAIL.n23 VTAIL.n2 9.69747
R766 VTAIL.n51 VTAIL.n30 9.69747
R767 VTAIL.n79 VTAIL.n58 9.69747
R768 VTAIL.n191 VTAIL.n170 9.69747
R769 VTAIL.n163 VTAIL.n142 9.69747
R770 VTAIL.n135 VTAIL.n114 9.69747
R771 VTAIL.n107 VTAIL.n86 9.69747
R772 VTAIL.n222 VTAIL.n221 9.45567
R773 VTAIL.n26 VTAIL.n25 9.45567
R774 VTAIL.n54 VTAIL.n53 9.45567
R775 VTAIL.n82 VTAIL.n81 9.45567
R776 VTAIL.n194 VTAIL.n193 9.45567
R777 VTAIL.n166 VTAIL.n165 9.45567
R778 VTAIL.n138 VTAIL.n137 9.45567
R779 VTAIL.n110 VTAIL.n109 9.45567
R780 VTAIL.n221 VTAIL.n220 9.3005
R781 VTAIL.n198 VTAIL.n197 9.3005
R782 VTAIL.n215 VTAIL.n214 9.3005
R783 VTAIL.n213 VTAIL.n212 9.3005
R784 VTAIL.n202 VTAIL.n201 9.3005
R785 VTAIL.n207 VTAIL.n206 9.3005
R786 VTAIL.n25 VTAIL.n24 9.3005
R787 VTAIL.n2 VTAIL.n1 9.3005
R788 VTAIL.n19 VTAIL.n18 9.3005
R789 VTAIL.n17 VTAIL.n16 9.3005
R790 VTAIL.n6 VTAIL.n5 9.3005
R791 VTAIL.n11 VTAIL.n10 9.3005
R792 VTAIL.n53 VTAIL.n52 9.3005
R793 VTAIL.n30 VTAIL.n29 9.3005
R794 VTAIL.n47 VTAIL.n46 9.3005
R795 VTAIL.n45 VTAIL.n44 9.3005
R796 VTAIL.n34 VTAIL.n33 9.3005
R797 VTAIL.n39 VTAIL.n38 9.3005
R798 VTAIL.n81 VTAIL.n80 9.3005
R799 VTAIL.n58 VTAIL.n57 9.3005
R800 VTAIL.n75 VTAIL.n74 9.3005
R801 VTAIL.n73 VTAIL.n72 9.3005
R802 VTAIL.n62 VTAIL.n61 9.3005
R803 VTAIL.n67 VTAIL.n66 9.3005
R804 VTAIL.n193 VTAIL.n192 9.3005
R805 VTAIL.n170 VTAIL.n169 9.3005
R806 VTAIL.n187 VTAIL.n186 9.3005
R807 VTAIL.n185 VTAIL.n184 9.3005
R808 VTAIL.n174 VTAIL.n173 9.3005
R809 VTAIL.n179 VTAIL.n178 9.3005
R810 VTAIL.n165 VTAIL.n164 9.3005
R811 VTAIL.n142 VTAIL.n141 9.3005
R812 VTAIL.n159 VTAIL.n158 9.3005
R813 VTAIL.n157 VTAIL.n156 9.3005
R814 VTAIL.n146 VTAIL.n145 9.3005
R815 VTAIL.n151 VTAIL.n150 9.3005
R816 VTAIL.n137 VTAIL.n136 9.3005
R817 VTAIL.n114 VTAIL.n113 9.3005
R818 VTAIL.n131 VTAIL.n130 9.3005
R819 VTAIL.n129 VTAIL.n128 9.3005
R820 VTAIL.n118 VTAIL.n117 9.3005
R821 VTAIL.n123 VTAIL.n122 9.3005
R822 VTAIL.n109 VTAIL.n108 9.3005
R823 VTAIL.n86 VTAIL.n85 9.3005
R824 VTAIL.n103 VTAIL.n102 9.3005
R825 VTAIL.n101 VTAIL.n100 9.3005
R826 VTAIL.n90 VTAIL.n89 9.3005
R827 VTAIL.n95 VTAIL.n94 9.3005
R828 VTAIL.n220 VTAIL.n196 8.92171
R829 VTAIL.n24 VTAIL.n0 8.92171
R830 VTAIL.n52 VTAIL.n28 8.92171
R831 VTAIL.n80 VTAIL.n56 8.92171
R832 VTAIL.n192 VTAIL.n168 8.92171
R833 VTAIL.n164 VTAIL.n140 8.92171
R834 VTAIL.n136 VTAIL.n112 8.92171
R835 VTAIL.n108 VTAIL.n84 8.92171
R836 VTAIL.n222 VTAIL.n196 5.04292
R837 VTAIL.n26 VTAIL.n0 5.04292
R838 VTAIL.n54 VTAIL.n28 5.04292
R839 VTAIL.n82 VTAIL.n56 5.04292
R840 VTAIL.n194 VTAIL.n168 5.04292
R841 VTAIL.n166 VTAIL.n140 5.04292
R842 VTAIL.n138 VTAIL.n112 5.04292
R843 VTAIL.n110 VTAIL.n84 5.04292
R844 VTAIL.n220 VTAIL.n219 4.26717
R845 VTAIL.n24 VTAIL.n23 4.26717
R846 VTAIL.n52 VTAIL.n51 4.26717
R847 VTAIL.n80 VTAIL.n79 4.26717
R848 VTAIL.n192 VTAIL.n191 4.26717
R849 VTAIL.n164 VTAIL.n163 4.26717
R850 VTAIL.n136 VTAIL.n135 4.26717
R851 VTAIL.n108 VTAIL.n107 4.26717
R852 VTAIL.n178 VTAIL.n177 3.71853
R853 VTAIL.n150 VTAIL.n149 3.71853
R854 VTAIL.n122 VTAIL.n121 3.71853
R855 VTAIL.n94 VTAIL.n93 3.71853
R856 VTAIL.n206 VTAIL.n205 3.71853
R857 VTAIL.n10 VTAIL.n9 3.71853
R858 VTAIL.n38 VTAIL.n37 3.71853
R859 VTAIL.n66 VTAIL.n65 3.71853
R860 VTAIL.n216 VTAIL.n198 3.49141
R861 VTAIL.n20 VTAIL.n2 3.49141
R862 VTAIL.n48 VTAIL.n30 3.49141
R863 VTAIL.n76 VTAIL.n58 3.49141
R864 VTAIL.n188 VTAIL.n170 3.49141
R865 VTAIL.n160 VTAIL.n142 3.49141
R866 VTAIL.n132 VTAIL.n114 3.49141
R867 VTAIL.n104 VTAIL.n86 3.49141
R868 VTAIL.n215 VTAIL.n200 2.71565
R869 VTAIL.n19 VTAIL.n4 2.71565
R870 VTAIL.n47 VTAIL.n32 2.71565
R871 VTAIL.n75 VTAIL.n60 2.71565
R872 VTAIL.n187 VTAIL.n172 2.71565
R873 VTAIL.n159 VTAIL.n144 2.71565
R874 VTAIL.n131 VTAIL.n116 2.71565
R875 VTAIL.n103 VTAIL.n88 2.71565
R876 VTAIL.n212 VTAIL.n211 1.93989
R877 VTAIL.n16 VTAIL.n15 1.93989
R878 VTAIL.n44 VTAIL.n43 1.93989
R879 VTAIL.n72 VTAIL.n71 1.93989
R880 VTAIL.n184 VTAIL.n183 1.93989
R881 VTAIL.n156 VTAIL.n155 1.93989
R882 VTAIL.n128 VTAIL.n127 1.93989
R883 VTAIL.n100 VTAIL.n99 1.93989
R884 VTAIL.n139 VTAIL.n111 1.22464
R885 VTAIL.n195 VTAIL.n167 1.22464
R886 VTAIL.n83 VTAIL.n55 1.22464
R887 VTAIL.n208 VTAIL.n202 1.16414
R888 VTAIL.n12 VTAIL.n6 1.16414
R889 VTAIL.n40 VTAIL.n34 1.16414
R890 VTAIL.n68 VTAIL.n62 1.16414
R891 VTAIL.n180 VTAIL.n174 1.16414
R892 VTAIL.n152 VTAIL.n146 1.16414
R893 VTAIL.n124 VTAIL.n118 1.16414
R894 VTAIL.n96 VTAIL.n90 1.16414
R895 VTAIL VTAIL.n27 0.670759
R896 VTAIL VTAIL.n223 0.554379
R897 VTAIL.n167 VTAIL.n139 0.470328
R898 VTAIL.n55 VTAIL.n27 0.470328
R899 VTAIL.n207 VTAIL.n204 0.388379
R900 VTAIL.n11 VTAIL.n8 0.388379
R901 VTAIL.n39 VTAIL.n36 0.388379
R902 VTAIL.n67 VTAIL.n64 0.388379
R903 VTAIL.n179 VTAIL.n176 0.388379
R904 VTAIL.n151 VTAIL.n148 0.388379
R905 VTAIL.n123 VTAIL.n120 0.388379
R906 VTAIL.n95 VTAIL.n92 0.388379
R907 VTAIL.n206 VTAIL.n201 0.155672
R908 VTAIL.n213 VTAIL.n201 0.155672
R909 VTAIL.n214 VTAIL.n213 0.155672
R910 VTAIL.n214 VTAIL.n197 0.155672
R911 VTAIL.n221 VTAIL.n197 0.155672
R912 VTAIL.n10 VTAIL.n5 0.155672
R913 VTAIL.n17 VTAIL.n5 0.155672
R914 VTAIL.n18 VTAIL.n17 0.155672
R915 VTAIL.n18 VTAIL.n1 0.155672
R916 VTAIL.n25 VTAIL.n1 0.155672
R917 VTAIL.n38 VTAIL.n33 0.155672
R918 VTAIL.n45 VTAIL.n33 0.155672
R919 VTAIL.n46 VTAIL.n45 0.155672
R920 VTAIL.n46 VTAIL.n29 0.155672
R921 VTAIL.n53 VTAIL.n29 0.155672
R922 VTAIL.n66 VTAIL.n61 0.155672
R923 VTAIL.n73 VTAIL.n61 0.155672
R924 VTAIL.n74 VTAIL.n73 0.155672
R925 VTAIL.n74 VTAIL.n57 0.155672
R926 VTAIL.n81 VTAIL.n57 0.155672
R927 VTAIL.n193 VTAIL.n169 0.155672
R928 VTAIL.n186 VTAIL.n169 0.155672
R929 VTAIL.n186 VTAIL.n185 0.155672
R930 VTAIL.n185 VTAIL.n173 0.155672
R931 VTAIL.n178 VTAIL.n173 0.155672
R932 VTAIL.n165 VTAIL.n141 0.155672
R933 VTAIL.n158 VTAIL.n141 0.155672
R934 VTAIL.n158 VTAIL.n157 0.155672
R935 VTAIL.n157 VTAIL.n145 0.155672
R936 VTAIL.n150 VTAIL.n145 0.155672
R937 VTAIL.n137 VTAIL.n113 0.155672
R938 VTAIL.n130 VTAIL.n113 0.155672
R939 VTAIL.n130 VTAIL.n129 0.155672
R940 VTAIL.n129 VTAIL.n117 0.155672
R941 VTAIL.n122 VTAIL.n117 0.155672
R942 VTAIL.n109 VTAIL.n85 0.155672
R943 VTAIL.n102 VTAIL.n85 0.155672
R944 VTAIL.n102 VTAIL.n101 0.155672
R945 VTAIL.n101 VTAIL.n89 0.155672
R946 VTAIL.n94 VTAIL.n89 0.155672
R947 VDD1 VDD1.n1 127.769
R948 VDD1 VDD1.n0 95.4496
R949 VDD1.n0 VDD1.t0 6.2756
R950 VDD1.n0 VDD1.t1 6.2756
R951 VDD1.n1 VDD1.t2 6.2756
R952 VDD1.n1 VDD1.t3 6.2756
R953 VN.n0 VN.t2 169.178
R954 VN.n1 VN.t1 169.178
R955 VN.n1 VN.t3 169.089
R956 VN.n0 VN.t0 169.089
R957 VN VN.n1 68.1221
R958 VN VN.n0 31.2622
R959 VDD2.n2 VDD2.n0 127.245
R960 VDD2.n2 VDD2.n1 95.3914
R961 VDD2.n1 VDD2.t0 6.2756
R962 VDD2.n1 VDD2.t2 6.2756
R963 VDD2.n0 VDD2.t1 6.2756
R964 VDD2.n0 VDD2.t3 6.2756
R965 VDD2 VDD2.n2 0.0586897
C0 w_n1822_n2004# VDD2 0.990848f
C1 VP VDD1 1.94734f
C2 B VTAIL 2.14375f
C3 VN VTAIL 1.8232f
C4 VDD1 VDD2 0.660055f
C5 VN B 0.746938f
C6 w_n1822_n2004# VTAIL 2.37975f
C7 VP VDD2 0.302645f
C8 B w_n1822_n2004# 5.47912f
C9 VDD1 VTAIL 3.50906f
C10 VN w_n1822_n2004# 2.66609f
C11 B VDD1 0.811536f
C12 VP VTAIL 1.83731f
C13 VN VDD1 0.14808f
C14 VTAIL VDD2 3.55315f
C15 B VP 1.12223f
C16 w_n1822_n2004# VDD1 0.968429f
C17 VN VP 3.83489f
C18 B VDD2 0.839188f
C19 VN VDD2 1.79715f
C20 VP w_n1822_n2004# 2.89642f
C21 VDD2 VSUBS 0.515331f
C22 VDD1 VSUBS 2.774327f
C23 VTAIL VSUBS 0.493836f
C24 VN VSUBS 3.89667f
C25 VP VSUBS 1.165674f
C26 B VSUBS 2.28392f
C27 w_n1822_n2004# VSUBS 45.7176f
C28 VDD2.t1 VSUBS 0.074607f
C29 VDD2.t3 VSUBS 0.074607f
C30 VDD2.n0 VSUBS 0.698727f
C31 VDD2.t0 VSUBS 0.074607f
C32 VDD2.t2 VSUBS 0.074607f
C33 VDD2.n1 VSUBS 0.472247f
C34 VDD2.n2 VSUBS 2.05478f
C35 VN.t2 VSUBS 0.659033f
C36 VN.t0 VSUBS 0.65885f
C37 VN.n0 VSUBS 0.532962f
C38 VN.t1 VSUBS 0.659033f
C39 VN.t3 VSUBS 0.65885f
C40 VN.n1 VSUBS 1.27997f
C41 VDD1.t0 VSUBS 0.071203f
C42 VDD1.t1 VSUBS 0.071203f
C43 VDD1.n0 VSUBS 0.450915f
C44 VDD1.t2 VSUBS 0.071203f
C45 VDD1.t3 VSUBS 0.071203f
C46 VDD1.n1 VSUBS 0.678538f
C47 VTAIL.n0 VSUBS 0.020861f
C48 VTAIL.n1 VSUBS 0.020151f
C49 VTAIL.n2 VSUBS 0.010828f
C50 VTAIL.n3 VSUBS 0.025594f
C51 VTAIL.n4 VSUBS 0.011465f
C52 VTAIL.n5 VSUBS 0.020151f
C53 VTAIL.n6 VSUBS 0.010828f
C54 VTAIL.n7 VSUBS 0.019195f
C55 VTAIL.n8 VSUBS 0.016257f
C56 VTAIL.t3 VSUBS 0.054998f
C57 VTAIL.n9 VSUBS 0.084287f
C58 VTAIL.n10 VSUBS 0.387056f
C59 VTAIL.n11 VSUBS 0.010828f
C60 VTAIL.n12 VSUBS 0.011465f
C61 VTAIL.n13 VSUBS 0.025594f
C62 VTAIL.n14 VSUBS 0.025594f
C63 VTAIL.n15 VSUBS 0.011465f
C64 VTAIL.n16 VSUBS 0.010828f
C65 VTAIL.n17 VSUBS 0.020151f
C66 VTAIL.n18 VSUBS 0.020151f
C67 VTAIL.n19 VSUBS 0.010828f
C68 VTAIL.n20 VSUBS 0.011465f
C69 VTAIL.n21 VSUBS 0.025594f
C70 VTAIL.n22 VSUBS 0.057599f
C71 VTAIL.n23 VSUBS 0.011465f
C72 VTAIL.n24 VSUBS 0.010828f
C73 VTAIL.n25 VSUBS 0.043824f
C74 VTAIL.n26 VSUBS 0.028685f
C75 VTAIL.n27 VSUBS 0.089684f
C76 VTAIL.n28 VSUBS 0.020861f
C77 VTAIL.n29 VSUBS 0.020151f
C78 VTAIL.n30 VSUBS 0.010828f
C79 VTAIL.n31 VSUBS 0.025594f
C80 VTAIL.n32 VSUBS 0.011465f
C81 VTAIL.n33 VSUBS 0.020151f
C82 VTAIL.n34 VSUBS 0.010828f
C83 VTAIL.n35 VSUBS 0.019195f
C84 VTAIL.n36 VSUBS 0.016257f
C85 VTAIL.t7 VSUBS 0.054998f
C86 VTAIL.n37 VSUBS 0.084287f
C87 VTAIL.n38 VSUBS 0.387056f
C88 VTAIL.n39 VSUBS 0.010828f
C89 VTAIL.n40 VSUBS 0.011465f
C90 VTAIL.n41 VSUBS 0.025594f
C91 VTAIL.n42 VSUBS 0.025594f
C92 VTAIL.n43 VSUBS 0.011465f
C93 VTAIL.n44 VSUBS 0.010828f
C94 VTAIL.n45 VSUBS 0.020151f
C95 VTAIL.n46 VSUBS 0.020151f
C96 VTAIL.n47 VSUBS 0.010828f
C97 VTAIL.n48 VSUBS 0.011465f
C98 VTAIL.n49 VSUBS 0.025594f
C99 VTAIL.n50 VSUBS 0.057599f
C100 VTAIL.n51 VSUBS 0.011465f
C101 VTAIL.n52 VSUBS 0.010828f
C102 VTAIL.n53 VSUBS 0.043824f
C103 VTAIL.n54 VSUBS 0.028685f
C104 VTAIL.n55 VSUBS 0.125647f
C105 VTAIL.n56 VSUBS 0.020861f
C106 VTAIL.n57 VSUBS 0.020151f
C107 VTAIL.n58 VSUBS 0.010828f
C108 VTAIL.n59 VSUBS 0.025594f
C109 VTAIL.n60 VSUBS 0.011465f
C110 VTAIL.n61 VSUBS 0.020151f
C111 VTAIL.n62 VSUBS 0.010828f
C112 VTAIL.n63 VSUBS 0.019195f
C113 VTAIL.n64 VSUBS 0.016257f
C114 VTAIL.t6 VSUBS 0.054998f
C115 VTAIL.n65 VSUBS 0.084287f
C116 VTAIL.n66 VSUBS 0.387056f
C117 VTAIL.n67 VSUBS 0.010828f
C118 VTAIL.n68 VSUBS 0.011465f
C119 VTAIL.n69 VSUBS 0.025594f
C120 VTAIL.n70 VSUBS 0.025594f
C121 VTAIL.n71 VSUBS 0.011465f
C122 VTAIL.n72 VSUBS 0.010828f
C123 VTAIL.n73 VSUBS 0.020151f
C124 VTAIL.n74 VSUBS 0.020151f
C125 VTAIL.n75 VSUBS 0.010828f
C126 VTAIL.n76 VSUBS 0.011465f
C127 VTAIL.n77 VSUBS 0.025594f
C128 VTAIL.n78 VSUBS 0.057599f
C129 VTAIL.n79 VSUBS 0.011465f
C130 VTAIL.n80 VSUBS 0.010828f
C131 VTAIL.n81 VSUBS 0.043824f
C132 VTAIL.n82 VSUBS 0.028685f
C133 VTAIL.n83 VSUBS 0.73829f
C134 VTAIL.n84 VSUBS 0.020861f
C135 VTAIL.n85 VSUBS 0.020151f
C136 VTAIL.n86 VSUBS 0.010828f
C137 VTAIL.n87 VSUBS 0.025594f
C138 VTAIL.n88 VSUBS 0.011465f
C139 VTAIL.n89 VSUBS 0.020151f
C140 VTAIL.n90 VSUBS 0.010828f
C141 VTAIL.n91 VSUBS 0.019195f
C142 VTAIL.n92 VSUBS 0.016257f
C143 VTAIL.t0 VSUBS 0.054998f
C144 VTAIL.n93 VSUBS 0.084287f
C145 VTAIL.n94 VSUBS 0.387056f
C146 VTAIL.n95 VSUBS 0.010828f
C147 VTAIL.n96 VSUBS 0.011465f
C148 VTAIL.n97 VSUBS 0.025594f
C149 VTAIL.n98 VSUBS 0.025594f
C150 VTAIL.n99 VSUBS 0.011465f
C151 VTAIL.n100 VSUBS 0.010828f
C152 VTAIL.n101 VSUBS 0.020151f
C153 VTAIL.n102 VSUBS 0.020151f
C154 VTAIL.n103 VSUBS 0.010828f
C155 VTAIL.n104 VSUBS 0.011465f
C156 VTAIL.n105 VSUBS 0.025594f
C157 VTAIL.n106 VSUBS 0.057599f
C158 VTAIL.n107 VSUBS 0.011465f
C159 VTAIL.n108 VSUBS 0.010828f
C160 VTAIL.n109 VSUBS 0.043824f
C161 VTAIL.n110 VSUBS 0.028685f
C162 VTAIL.n111 VSUBS 0.73829f
C163 VTAIL.n112 VSUBS 0.020861f
C164 VTAIL.n113 VSUBS 0.020151f
C165 VTAIL.n114 VSUBS 0.010828f
C166 VTAIL.n115 VSUBS 0.025594f
C167 VTAIL.n116 VSUBS 0.011465f
C168 VTAIL.n117 VSUBS 0.020151f
C169 VTAIL.n118 VSUBS 0.010828f
C170 VTAIL.n119 VSUBS 0.019195f
C171 VTAIL.n120 VSUBS 0.016257f
C172 VTAIL.t2 VSUBS 0.054998f
C173 VTAIL.n121 VSUBS 0.084287f
C174 VTAIL.n122 VSUBS 0.387056f
C175 VTAIL.n123 VSUBS 0.010828f
C176 VTAIL.n124 VSUBS 0.011465f
C177 VTAIL.n125 VSUBS 0.025594f
C178 VTAIL.n126 VSUBS 0.025594f
C179 VTAIL.n127 VSUBS 0.011465f
C180 VTAIL.n128 VSUBS 0.010828f
C181 VTAIL.n129 VSUBS 0.020151f
C182 VTAIL.n130 VSUBS 0.020151f
C183 VTAIL.n131 VSUBS 0.010828f
C184 VTAIL.n132 VSUBS 0.011465f
C185 VTAIL.n133 VSUBS 0.025594f
C186 VTAIL.n134 VSUBS 0.057599f
C187 VTAIL.n135 VSUBS 0.011465f
C188 VTAIL.n136 VSUBS 0.010828f
C189 VTAIL.n137 VSUBS 0.043824f
C190 VTAIL.n138 VSUBS 0.028685f
C191 VTAIL.n139 VSUBS 0.125647f
C192 VTAIL.n140 VSUBS 0.020861f
C193 VTAIL.n141 VSUBS 0.020151f
C194 VTAIL.n142 VSUBS 0.010828f
C195 VTAIL.n143 VSUBS 0.025594f
C196 VTAIL.n144 VSUBS 0.011465f
C197 VTAIL.n145 VSUBS 0.020151f
C198 VTAIL.n146 VSUBS 0.010828f
C199 VTAIL.n147 VSUBS 0.019195f
C200 VTAIL.n148 VSUBS 0.016257f
C201 VTAIL.t4 VSUBS 0.054998f
C202 VTAIL.n149 VSUBS 0.084287f
C203 VTAIL.n150 VSUBS 0.387056f
C204 VTAIL.n151 VSUBS 0.010828f
C205 VTAIL.n152 VSUBS 0.011465f
C206 VTAIL.n153 VSUBS 0.025594f
C207 VTAIL.n154 VSUBS 0.025594f
C208 VTAIL.n155 VSUBS 0.011465f
C209 VTAIL.n156 VSUBS 0.010828f
C210 VTAIL.n157 VSUBS 0.020151f
C211 VTAIL.n158 VSUBS 0.020151f
C212 VTAIL.n159 VSUBS 0.010828f
C213 VTAIL.n160 VSUBS 0.011465f
C214 VTAIL.n161 VSUBS 0.025594f
C215 VTAIL.n162 VSUBS 0.057599f
C216 VTAIL.n163 VSUBS 0.011465f
C217 VTAIL.n164 VSUBS 0.010828f
C218 VTAIL.n165 VSUBS 0.043824f
C219 VTAIL.n166 VSUBS 0.028685f
C220 VTAIL.n167 VSUBS 0.125647f
C221 VTAIL.n168 VSUBS 0.020861f
C222 VTAIL.n169 VSUBS 0.020151f
C223 VTAIL.n170 VSUBS 0.010828f
C224 VTAIL.n171 VSUBS 0.025594f
C225 VTAIL.n172 VSUBS 0.011465f
C226 VTAIL.n173 VSUBS 0.020151f
C227 VTAIL.n174 VSUBS 0.010828f
C228 VTAIL.n175 VSUBS 0.019195f
C229 VTAIL.n176 VSUBS 0.016257f
C230 VTAIL.t5 VSUBS 0.054998f
C231 VTAIL.n177 VSUBS 0.084287f
C232 VTAIL.n178 VSUBS 0.387056f
C233 VTAIL.n179 VSUBS 0.010828f
C234 VTAIL.n180 VSUBS 0.011465f
C235 VTAIL.n181 VSUBS 0.025594f
C236 VTAIL.n182 VSUBS 0.025594f
C237 VTAIL.n183 VSUBS 0.011465f
C238 VTAIL.n184 VSUBS 0.010828f
C239 VTAIL.n185 VSUBS 0.020151f
C240 VTAIL.n186 VSUBS 0.020151f
C241 VTAIL.n187 VSUBS 0.010828f
C242 VTAIL.n188 VSUBS 0.011465f
C243 VTAIL.n189 VSUBS 0.025594f
C244 VTAIL.n190 VSUBS 0.057599f
C245 VTAIL.n191 VSUBS 0.011465f
C246 VTAIL.n192 VSUBS 0.010828f
C247 VTAIL.n193 VSUBS 0.043824f
C248 VTAIL.n194 VSUBS 0.028685f
C249 VTAIL.n195 VSUBS 0.73829f
C250 VTAIL.n196 VSUBS 0.020861f
C251 VTAIL.n197 VSUBS 0.020151f
C252 VTAIL.n198 VSUBS 0.010828f
C253 VTAIL.n199 VSUBS 0.025594f
C254 VTAIL.n200 VSUBS 0.011465f
C255 VTAIL.n201 VSUBS 0.020151f
C256 VTAIL.n202 VSUBS 0.010828f
C257 VTAIL.n203 VSUBS 0.019195f
C258 VTAIL.n204 VSUBS 0.016257f
C259 VTAIL.t1 VSUBS 0.054998f
C260 VTAIL.n205 VSUBS 0.084287f
C261 VTAIL.n206 VSUBS 0.387056f
C262 VTAIL.n207 VSUBS 0.010828f
C263 VTAIL.n208 VSUBS 0.011465f
C264 VTAIL.n209 VSUBS 0.025594f
C265 VTAIL.n210 VSUBS 0.025594f
C266 VTAIL.n211 VSUBS 0.011465f
C267 VTAIL.n212 VSUBS 0.010828f
C268 VTAIL.n213 VSUBS 0.020151f
C269 VTAIL.n214 VSUBS 0.020151f
C270 VTAIL.n215 VSUBS 0.010828f
C271 VTAIL.n216 VSUBS 0.011465f
C272 VTAIL.n217 VSUBS 0.025594f
C273 VTAIL.n218 VSUBS 0.057599f
C274 VTAIL.n219 VSUBS 0.011465f
C275 VTAIL.n220 VSUBS 0.010828f
C276 VTAIL.n221 VSUBS 0.043824f
C277 VTAIL.n222 VSUBS 0.028685f
C278 VTAIL.n223 VSUBS 0.69477f
C279 VP.t2 VSUBS 0.684754f
C280 VP.t3 VSUBS 0.684944f
C281 VP.n0 VSUBS 1.31523f
C282 VP.n1 VSUBS 2.00107f
C283 VP.t1 VSUBS 0.650744f
C284 VP.n2 VSUBS 0.310518f
C285 VP.t0 VSUBS 0.650744f
C286 VP.n3 VSUBS 0.310518f
C287 VP.n4 VSUBS 0.050231f
C288 B.n0 VSUBS 0.008214f
C289 B.n1 VSUBS 0.008214f
C290 B.n2 VSUBS 0.012148f
C291 B.n3 VSUBS 0.009309f
C292 B.n4 VSUBS 0.009309f
C293 B.n5 VSUBS 0.009309f
C294 B.n6 VSUBS 0.009309f
C295 B.n7 VSUBS 0.009309f
C296 B.n8 VSUBS 0.009309f
C297 B.n9 VSUBS 0.009309f
C298 B.n10 VSUBS 0.009309f
C299 B.n11 VSUBS 0.009309f
C300 B.n12 VSUBS 0.022429f
C301 B.n13 VSUBS 0.009309f
C302 B.n14 VSUBS 0.009309f
C303 B.n15 VSUBS 0.009309f
C304 B.n16 VSUBS 0.009309f
C305 B.n17 VSUBS 0.009309f
C306 B.n18 VSUBS 0.009309f
C307 B.n19 VSUBS 0.009309f
C308 B.n20 VSUBS 0.009309f
C309 B.n21 VSUBS 0.009309f
C310 B.n22 VSUBS 0.009309f
C311 B.n23 VSUBS 0.009309f
C312 B.t4 VSUBS 0.100255f
C313 B.t5 VSUBS 0.116487f
C314 B.t3 VSUBS 0.339869f
C315 B.n24 VSUBS 0.20963f
C316 B.n25 VSUBS 0.179047f
C317 B.n26 VSUBS 0.009309f
C318 B.n27 VSUBS 0.009309f
C319 B.n28 VSUBS 0.009309f
C320 B.n29 VSUBS 0.009309f
C321 B.t10 VSUBS 0.100257f
C322 B.t11 VSUBS 0.116489f
C323 B.t9 VSUBS 0.339869f
C324 B.n30 VSUBS 0.209628f
C325 B.n31 VSUBS 0.179045f
C326 B.n32 VSUBS 0.009309f
C327 B.n33 VSUBS 0.009309f
C328 B.n34 VSUBS 0.009309f
C329 B.n35 VSUBS 0.009309f
C330 B.n36 VSUBS 0.009309f
C331 B.n37 VSUBS 0.009309f
C332 B.n38 VSUBS 0.009309f
C333 B.n39 VSUBS 0.009309f
C334 B.n40 VSUBS 0.009309f
C335 B.n41 VSUBS 0.009309f
C336 B.n42 VSUBS 0.022429f
C337 B.n43 VSUBS 0.009309f
C338 B.n44 VSUBS 0.009309f
C339 B.n45 VSUBS 0.009309f
C340 B.n46 VSUBS 0.009309f
C341 B.n47 VSUBS 0.009309f
C342 B.n48 VSUBS 0.009309f
C343 B.n49 VSUBS 0.009309f
C344 B.n50 VSUBS 0.009309f
C345 B.n51 VSUBS 0.009309f
C346 B.n52 VSUBS 0.009309f
C347 B.n53 VSUBS 0.009309f
C348 B.n54 VSUBS 0.009309f
C349 B.n55 VSUBS 0.009309f
C350 B.n56 VSUBS 0.009309f
C351 B.n57 VSUBS 0.009309f
C352 B.n58 VSUBS 0.009309f
C353 B.n59 VSUBS 0.009309f
C354 B.n60 VSUBS 0.009309f
C355 B.n61 VSUBS 0.009309f
C356 B.n62 VSUBS 0.009309f
C357 B.n63 VSUBS 0.02083f
C358 B.n64 VSUBS 0.009309f
C359 B.n65 VSUBS 0.009309f
C360 B.n66 VSUBS 0.009309f
C361 B.n67 VSUBS 0.009309f
C362 B.n68 VSUBS 0.009309f
C363 B.n69 VSUBS 0.009309f
C364 B.n70 VSUBS 0.009309f
C365 B.n71 VSUBS 0.009309f
C366 B.n72 VSUBS 0.009309f
C367 B.n73 VSUBS 0.009309f
C368 B.n74 VSUBS 0.006434f
C369 B.n75 VSUBS 0.009309f
C370 B.n76 VSUBS 0.009309f
C371 B.n77 VSUBS 0.009309f
C372 B.n78 VSUBS 0.009309f
C373 B.n79 VSUBS 0.009309f
C374 B.t2 VSUBS 0.100255f
C375 B.t1 VSUBS 0.116487f
C376 B.t0 VSUBS 0.339869f
C377 B.n80 VSUBS 0.20963f
C378 B.n81 VSUBS 0.179047f
C379 B.n82 VSUBS 0.009309f
C380 B.n83 VSUBS 0.009309f
C381 B.n84 VSUBS 0.009309f
C382 B.n85 VSUBS 0.009309f
C383 B.n86 VSUBS 0.009309f
C384 B.n87 VSUBS 0.009309f
C385 B.n88 VSUBS 0.009309f
C386 B.n89 VSUBS 0.009309f
C387 B.n90 VSUBS 0.009309f
C388 B.n91 VSUBS 0.009309f
C389 B.n92 VSUBS 0.02083f
C390 B.n93 VSUBS 0.009309f
C391 B.n94 VSUBS 0.009309f
C392 B.n95 VSUBS 0.009309f
C393 B.n96 VSUBS 0.009309f
C394 B.n97 VSUBS 0.009309f
C395 B.n98 VSUBS 0.009309f
C396 B.n99 VSUBS 0.009309f
C397 B.n100 VSUBS 0.009309f
C398 B.n101 VSUBS 0.009309f
C399 B.n102 VSUBS 0.009309f
C400 B.n103 VSUBS 0.009309f
C401 B.n104 VSUBS 0.009309f
C402 B.n105 VSUBS 0.009309f
C403 B.n106 VSUBS 0.009309f
C404 B.n107 VSUBS 0.009309f
C405 B.n108 VSUBS 0.009309f
C406 B.n109 VSUBS 0.009309f
C407 B.n110 VSUBS 0.009309f
C408 B.n111 VSUBS 0.009309f
C409 B.n112 VSUBS 0.009309f
C410 B.n113 VSUBS 0.009309f
C411 B.n114 VSUBS 0.009309f
C412 B.n115 VSUBS 0.009309f
C413 B.n116 VSUBS 0.009309f
C414 B.n117 VSUBS 0.009309f
C415 B.n118 VSUBS 0.009309f
C416 B.n119 VSUBS 0.009309f
C417 B.n120 VSUBS 0.009309f
C418 B.n121 VSUBS 0.009309f
C419 B.n122 VSUBS 0.009309f
C420 B.n123 VSUBS 0.009309f
C421 B.n124 VSUBS 0.009309f
C422 B.n125 VSUBS 0.009309f
C423 B.n126 VSUBS 0.009309f
C424 B.n127 VSUBS 0.009309f
C425 B.n128 VSUBS 0.009309f
C426 B.n129 VSUBS 0.02083f
C427 B.n130 VSUBS 0.022429f
C428 B.n131 VSUBS 0.022429f
C429 B.n132 VSUBS 0.009309f
C430 B.n133 VSUBS 0.009309f
C431 B.n134 VSUBS 0.009309f
C432 B.n135 VSUBS 0.009309f
C433 B.n136 VSUBS 0.009309f
C434 B.n137 VSUBS 0.009309f
C435 B.n138 VSUBS 0.009309f
C436 B.n139 VSUBS 0.009309f
C437 B.n140 VSUBS 0.009309f
C438 B.n141 VSUBS 0.009309f
C439 B.n142 VSUBS 0.009309f
C440 B.n143 VSUBS 0.009309f
C441 B.n144 VSUBS 0.009309f
C442 B.n145 VSUBS 0.009309f
C443 B.n146 VSUBS 0.009309f
C444 B.n147 VSUBS 0.009309f
C445 B.n148 VSUBS 0.009309f
C446 B.n149 VSUBS 0.009309f
C447 B.n150 VSUBS 0.009309f
C448 B.n151 VSUBS 0.009309f
C449 B.n152 VSUBS 0.009309f
C450 B.n153 VSUBS 0.009309f
C451 B.n154 VSUBS 0.009309f
C452 B.n155 VSUBS 0.009309f
C453 B.n156 VSUBS 0.009309f
C454 B.n157 VSUBS 0.009309f
C455 B.n158 VSUBS 0.009309f
C456 B.n159 VSUBS 0.009309f
C457 B.n160 VSUBS 0.009309f
C458 B.n161 VSUBS 0.009309f
C459 B.n162 VSUBS 0.006434f
C460 B.n163 VSUBS 0.021568f
C461 B.n164 VSUBS 0.007529f
C462 B.n165 VSUBS 0.009309f
C463 B.n166 VSUBS 0.009309f
C464 B.n167 VSUBS 0.009309f
C465 B.n168 VSUBS 0.009309f
C466 B.n169 VSUBS 0.009309f
C467 B.n170 VSUBS 0.009309f
C468 B.n171 VSUBS 0.009309f
C469 B.n172 VSUBS 0.009309f
C470 B.n173 VSUBS 0.009309f
C471 B.n174 VSUBS 0.009309f
C472 B.n175 VSUBS 0.009309f
C473 B.t8 VSUBS 0.100257f
C474 B.t7 VSUBS 0.116489f
C475 B.t6 VSUBS 0.339869f
C476 B.n176 VSUBS 0.209628f
C477 B.n177 VSUBS 0.179045f
C478 B.n178 VSUBS 0.021568f
C479 B.n179 VSUBS 0.007529f
C480 B.n180 VSUBS 0.009309f
C481 B.n181 VSUBS 0.009309f
C482 B.n182 VSUBS 0.009309f
C483 B.n183 VSUBS 0.009309f
C484 B.n184 VSUBS 0.009309f
C485 B.n185 VSUBS 0.009309f
C486 B.n186 VSUBS 0.009309f
C487 B.n187 VSUBS 0.009309f
C488 B.n188 VSUBS 0.009309f
C489 B.n189 VSUBS 0.009309f
C490 B.n190 VSUBS 0.009309f
C491 B.n191 VSUBS 0.009309f
C492 B.n192 VSUBS 0.009309f
C493 B.n193 VSUBS 0.009309f
C494 B.n194 VSUBS 0.009309f
C495 B.n195 VSUBS 0.009309f
C496 B.n196 VSUBS 0.009309f
C497 B.n197 VSUBS 0.009309f
C498 B.n198 VSUBS 0.009309f
C499 B.n199 VSUBS 0.009309f
C500 B.n200 VSUBS 0.009309f
C501 B.n201 VSUBS 0.009309f
C502 B.n202 VSUBS 0.009309f
C503 B.n203 VSUBS 0.009309f
C504 B.n204 VSUBS 0.009309f
C505 B.n205 VSUBS 0.009309f
C506 B.n206 VSUBS 0.009309f
C507 B.n207 VSUBS 0.009309f
C508 B.n208 VSUBS 0.009309f
C509 B.n209 VSUBS 0.009309f
C510 B.n210 VSUBS 0.009309f
C511 B.n211 VSUBS 0.009309f
C512 B.n212 VSUBS 0.022429f
C513 B.n213 VSUBS 0.021318f
C514 B.n214 VSUBS 0.021941f
C515 B.n215 VSUBS 0.009309f
C516 B.n216 VSUBS 0.009309f
C517 B.n217 VSUBS 0.009309f
C518 B.n218 VSUBS 0.009309f
C519 B.n219 VSUBS 0.009309f
C520 B.n220 VSUBS 0.009309f
C521 B.n221 VSUBS 0.009309f
C522 B.n222 VSUBS 0.009309f
C523 B.n223 VSUBS 0.009309f
C524 B.n224 VSUBS 0.009309f
C525 B.n225 VSUBS 0.009309f
C526 B.n226 VSUBS 0.009309f
C527 B.n227 VSUBS 0.009309f
C528 B.n228 VSUBS 0.009309f
C529 B.n229 VSUBS 0.009309f
C530 B.n230 VSUBS 0.009309f
C531 B.n231 VSUBS 0.009309f
C532 B.n232 VSUBS 0.009309f
C533 B.n233 VSUBS 0.009309f
C534 B.n234 VSUBS 0.009309f
C535 B.n235 VSUBS 0.009309f
C536 B.n236 VSUBS 0.009309f
C537 B.n237 VSUBS 0.009309f
C538 B.n238 VSUBS 0.009309f
C539 B.n239 VSUBS 0.009309f
C540 B.n240 VSUBS 0.009309f
C541 B.n241 VSUBS 0.009309f
C542 B.n242 VSUBS 0.009309f
C543 B.n243 VSUBS 0.009309f
C544 B.n244 VSUBS 0.009309f
C545 B.n245 VSUBS 0.009309f
C546 B.n246 VSUBS 0.009309f
C547 B.n247 VSUBS 0.009309f
C548 B.n248 VSUBS 0.009309f
C549 B.n249 VSUBS 0.009309f
C550 B.n250 VSUBS 0.009309f
C551 B.n251 VSUBS 0.009309f
C552 B.n252 VSUBS 0.009309f
C553 B.n253 VSUBS 0.009309f
C554 B.n254 VSUBS 0.009309f
C555 B.n255 VSUBS 0.009309f
C556 B.n256 VSUBS 0.009309f
C557 B.n257 VSUBS 0.009309f
C558 B.n258 VSUBS 0.009309f
C559 B.n259 VSUBS 0.009309f
C560 B.n260 VSUBS 0.009309f
C561 B.n261 VSUBS 0.009309f
C562 B.n262 VSUBS 0.009309f
C563 B.n263 VSUBS 0.009309f
C564 B.n264 VSUBS 0.009309f
C565 B.n265 VSUBS 0.009309f
C566 B.n266 VSUBS 0.009309f
C567 B.n267 VSUBS 0.009309f
C568 B.n268 VSUBS 0.009309f
C569 B.n269 VSUBS 0.009309f
C570 B.n270 VSUBS 0.009309f
C571 B.n271 VSUBS 0.009309f
C572 B.n272 VSUBS 0.009309f
C573 B.n273 VSUBS 0.009309f
C574 B.n274 VSUBS 0.009309f
C575 B.n275 VSUBS 0.02083f
C576 B.n276 VSUBS 0.02083f
C577 B.n277 VSUBS 0.022429f
C578 B.n278 VSUBS 0.009309f
C579 B.n279 VSUBS 0.009309f
C580 B.n280 VSUBS 0.009309f
C581 B.n281 VSUBS 0.009309f
C582 B.n282 VSUBS 0.009309f
C583 B.n283 VSUBS 0.009309f
C584 B.n284 VSUBS 0.009309f
C585 B.n285 VSUBS 0.009309f
C586 B.n286 VSUBS 0.009309f
C587 B.n287 VSUBS 0.009309f
C588 B.n288 VSUBS 0.009309f
C589 B.n289 VSUBS 0.009309f
C590 B.n290 VSUBS 0.009309f
C591 B.n291 VSUBS 0.009309f
C592 B.n292 VSUBS 0.009309f
C593 B.n293 VSUBS 0.009309f
C594 B.n294 VSUBS 0.009309f
C595 B.n295 VSUBS 0.009309f
C596 B.n296 VSUBS 0.009309f
C597 B.n297 VSUBS 0.009309f
C598 B.n298 VSUBS 0.009309f
C599 B.n299 VSUBS 0.009309f
C600 B.n300 VSUBS 0.009309f
C601 B.n301 VSUBS 0.009309f
C602 B.n302 VSUBS 0.009309f
C603 B.n303 VSUBS 0.009309f
C604 B.n304 VSUBS 0.009309f
C605 B.n305 VSUBS 0.009309f
C606 B.n306 VSUBS 0.009309f
C607 B.n307 VSUBS 0.009309f
C608 B.n308 VSUBS 0.009309f
C609 B.n309 VSUBS 0.006434f
C610 B.n310 VSUBS 0.021568f
C611 B.n311 VSUBS 0.007529f
C612 B.n312 VSUBS 0.009309f
C613 B.n313 VSUBS 0.009309f
C614 B.n314 VSUBS 0.009309f
C615 B.n315 VSUBS 0.009309f
C616 B.n316 VSUBS 0.009309f
C617 B.n317 VSUBS 0.009309f
C618 B.n318 VSUBS 0.009309f
C619 B.n319 VSUBS 0.009309f
C620 B.n320 VSUBS 0.009309f
C621 B.n321 VSUBS 0.009309f
C622 B.n322 VSUBS 0.009309f
C623 B.n323 VSUBS 0.007529f
C624 B.n324 VSUBS 0.021568f
C625 B.n325 VSUBS 0.006434f
C626 B.n326 VSUBS 0.009309f
C627 B.n327 VSUBS 0.009309f
C628 B.n328 VSUBS 0.009309f
C629 B.n329 VSUBS 0.009309f
C630 B.n330 VSUBS 0.009309f
C631 B.n331 VSUBS 0.009309f
C632 B.n332 VSUBS 0.009309f
C633 B.n333 VSUBS 0.009309f
C634 B.n334 VSUBS 0.009309f
C635 B.n335 VSUBS 0.009309f
C636 B.n336 VSUBS 0.009309f
C637 B.n337 VSUBS 0.009309f
C638 B.n338 VSUBS 0.009309f
C639 B.n339 VSUBS 0.009309f
C640 B.n340 VSUBS 0.009309f
C641 B.n341 VSUBS 0.009309f
C642 B.n342 VSUBS 0.009309f
C643 B.n343 VSUBS 0.009309f
C644 B.n344 VSUBS 0.009309f
C645 B.n345 VSUBS 0.009309f
C646 B.n346 VSUBS 0.009309f
C647 B.n347 VSUBS 0.009309f
C648 B.n348 VSUBS 0.009309f
C649 B.n349 VSUBS 0.009309f
C650 B.n350 VSUBS 0.009309f
C651 B.n351 VSUBS 0.009309f
C652 B.n352 VSUBS 0.009309f
C653 B.n353 VSUBS 0.009309f
C654 B.n354 VSUBS 0.009309f
C655 B.n355 VSUBS 0.009309f
C656 B.n356 VSUBS 0.009309f
C657 B.n357 VSUBS 0.022429f
C658 B.n358 VSUBS 0.02083f
C659 B.n359 VSUBS 0.02083f
C660 B.n360 VSUBS 0.009309f
C661 B.n361 VSUBS 0.009309f
C662 B.n362 VSUBS 0.009309f
C663 B.n363 VSUBS 0.009309f
C664 B.n364 VSUBS 0.009309f
C665 B.n365 VSUBS 0.009309f
C666 B.n366 VSUBS 0.009309f
C667 B.n367 VSUBS 0.009309f
C668 B.n368 VSUBS 0.009309f
C669 B.n369 VSUBS 0.009309f
C670 B.n370 VSUBS 0.009309f
C671 B.n371 VSUBS 0.009309f
C672 B.n372 VSUBS 0.009309f
C673 B.n373 VSUBS 0.009309f
C674 B.n374 VSUBS 0.009309f
C675 B.n375 VSUBS 0.009309f
C676 B.n376 VSUBS 0.009309f
C677 B.n377 VSUBS 0.009309f
C678 B.n378 VSUBS 0.009309f
C679 B.n379 VSUBS 0.009309f
C680 B.n380 VSUBS 0.009309f
C681 B.n381 VSUBS 0.009309f
C682 B.n382 VSUBS 0.009309f
C683 B.n383 VSUBS 0.009309f
C684 B.n384 VSUBS 0.009309f
C685 B.n385 VSUBS 0.009309f
C686 B.n386 VSUBS 0.009309f
C687 B.n387 VSUBS 0.012148f
C688 B.n388 VSUBS 0.01294f
C689 B.n389 VSUBS 0.025733f
.ends

