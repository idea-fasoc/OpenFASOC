* NGSPICE file created from diff_pair_sample_1143.ext - technology: sky130A

.subckt diff_pair_sample_1143 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t1 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X1 VTAIL.t17 VP.t1 VDD1.t3 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X2 VTAIL.t16 VP.t2 VDD1.t6 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X3 B.t11 B.t9 B.t10 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0 ps=0 w=4.85 l=3.42
X4 VTAIL.t1 VN.t0 VDD2.t9 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X5 VDD2.t8 VN.t1 VTAIL.t2 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X6 VDD2.t7 VN.t2 VTAIL.t5 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0.80025 ps=5.18 w=4.85 l=3.42
X7 B.t8 B.t6 B.t7 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0 ps=0 w=4.85 l=3.42
X8 VDD2.t6 VN.t3 VTAIL.t0 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X9 VDD1.t4 VP.t3 VTAIL.t15 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X10 VTAIL.t8 VN.t4 VDD2.t5 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X11 VTAIL.t14 VP.t4 VDD1.t5 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X12 VDD2.t4 VN.t5 VTAIL.t7 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=1.8915 ps=10.48 w=4.85 l=3.42
X13 VTAIL.t19 VN.t6 VDD2.t3 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X14 VDD1.t7 VP.t5 VTAIL.t13 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0.80025 ps=5.18 w=4.85 l=3.42
X15 VDD1.t0 VP.t6 VTAIL.t12 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
X16 VDD1.t2 VP.t7 VTAIL.t11 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0.80025 ps=5.18 w=4.85 l=3.42
X17 B.t5 B.t3 B.t4 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0 ps=0 w=4.85 l=3.42
X18 B.t2 B.t0 B.t1 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0 ps=0 w=4.85 l=3.42
X19 VDD2.t2 VN.t7 VTAIL.t4 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=1.8915 pd=10.48 as=0.80025 ps=5.18 w=4.85 l=3.42
X20 VDD2.t1 VN.t8 VTAIL.t6 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=1.8915 ps=10.48 w=4.85 l=3.42
X21 VDD1.t9 VP.t8 VTAIL.t10 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=1.8915 ps=10.48 w=4.85 l=3.42
X22 VDD1.t8 VP.t9 VTAIL.t9 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=1.8915 ps=10.48 w=4.85 l=3.42
X23 VTAIL.t3 VN.t9 VDD2.t0 w_n5470_n1938# sky130_fd_pr__pfet_01v8 ad=0.80025 pd=5.18 as=0.80025 ps=5.18 w=4.85 l=3.42
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n53 VP.n21 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n20 161.3
R17 VP.n58 VP.n57 161.3
R18 VP.n59 VP.n19 161.3
R19 VP.n61 VP.n60 161.3
R20 VP.n62 VP.n18 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n112 VP.n111 161.3
R23 VP.n110 VP.n1 161.3
R24 VP.n109 VP.n108 161.3
R25 VP.n107 VP.n2 161.3
R26 VP.n106 VP.n105 161.3
R27 VP.n104 VP.n3 161.3
R28 VP.n103 VP.n102 161.3
R29 VP.n101 VP.n4 161.3
R30 VP.n100 VP.n99 161.3
R31 VP.n98 VP.n5 161.3
R32 VP.n97 VP.n96 161.3
R33 VP.n95 VP.n6 161.3
R34 VP.n94 VP.n93 161.3
R35 VP.n92 VP.n7 161.3
R36 VP.n91 VP.n90 161.3
R37 VP.n89 VP.n88 161.3
R38 VP.n87 VP.n9 161.3
R39 VP.n86 VP.n85 161.3
R40 VP.n84 VP.n10 161.3
R41 VP.n83 VP.n82 161.3
R42 VP.n81 VP.n11 161.3
R43 VP.n80 VP.n79 161.3
R44 VP.n78 VP.n12 161.3
R45 VP.n77 VP.n76 161.3
R46 VP.n75 VP.n13 161.3
R47 VP.n74 VP.n73 161.3
R48 VP.n72 VP.n14 161.3
R49 VP.n71 VP.n70 161.3
R50 VP.n69 VP.n15 161.3
R51 VP.n68 VP.n67 161.3
R52 VP.n66 VP.n16 77.8339
R53 VP.n113 VP.n0 77.8339
R54 VP.n65 VP.n17 77.8339
R55 VP.n30 VP.t5 67.9561
R56 VP.n74 VP.n14 52.6342
R57 VP.n82 VP.n10 52.6342
R58 VP.n97 VP.n6 52.6342
R59 VP.n105 VP.n2 52.6342
R60 VP.n57 VP.n19 52.6342
R61 VP.n49 VP.n23 52.6342
R62 VP.n34 VP.n27 52.6342
R63 VP.n66 VP.n65 52.2607
R64 VP.n30 VP.n29 50.1549
R65 VP.n4 VP.t2 34.1774
R66 VP.n12 VP.t4 34.1774
R67 VP.n16 VP.t7 34.1774
R68 VP.n8 VP.t3 34.1774
R69 VP.n0 VP.t8 34.1774
R70 VP.n29 VP.t1 34.1774
R71 VP.n21 VP.t0 34.1774
R72 VP.n17 VP.t9 34.1774
R73 VP.n25 VP.t6 34.1774
R74 VP.n70 VP.n14 28.3526
R75 VP.n86 VP.n10 28.3526
R76 VP.n93 VP.n6 28.3526
R77 VP.n109 VP.n2 28.3526
R78 VP.n61 VP.n19 28.3526
R79 VP.n45 VP.n23 28.3526
R80 VP.n38 VP.n27 28.3526
R81 VP.n69 VP.n68 24.4675
R82 VP.n70 VP.n69 24.4675
R83 VP.n75 VP.n74 24.4675
R84 VP.n76 VP.n75 24.4675
R85 VP.n76 VP.n12 24.4675
R86 VP.n80 VP.n12 24.4675
R87 VP.n81 VP.n80 24.4675
R88 VP.n82 VP.n81 24.4675
R89 VP.n87 VP.n86 24.4675
R90 VP.n88 VP.n87 24.4675
R91 VP.n92 VP.n91 24.4675
R92 VP.n93 VP.n92 24.4675
R93 VP.n98 VP.n97 24.4675
R94 VP.n99 VP.n98 24.4675
R95 VP.n99 VP.n4 24.4675
R96 VP.n103 VP.n4 24.4675
R97 VP.n104 VP.n103 24.4675
R98 VP.n105 VP.n104 24.4675
R99 VP.n110 VP.n109 24.4675
R100 VP.n111 VP.n110 24.4675
R101 VP.n62 VP.n61 24.4675
R102 VP.n63 VP.n62 24.4675
R103 VP.n50 VP.n49 24.4675
R104 VP.n51 VP.n50 24.4675
R105 VP.n51 VP.n21 24.4675
R106 VP.n55 VP.n21 24.4675
R107 VP.n56 VP.n55 24.4675
R108 VP.n57 VP.n56 24.4675
R109 VP.n39 VP.n38 24.4675
R110 VP.n40 VP.n39 24.4675
R111 VP.n44 VP.n43 24.4675
R112 VP.n45 VP.n44 24.4675
R113 VP.n32 VP.n29 24.4675
R114 VP.n33 VP.n32 24.4675
R115 VP.n34 VP.n33 24.4675
R116 VP.n68 VP.n16 12.234
R117 VP.n88 VP.n8 12.234
R118 VP.n91 VP.n8 12.234
R119 VP.n111 VP.n0 12.234
R120 VP.n63 VP.n17 12.234
R121 VP.n40 VP.n25 12.234
R122 VP.n43 VP.n25 12.234
R123 VP.n31 VP.n30 3.07681
R124 VP.n65 VP.n64 0.354971
R125 VP.n67 VP.n66 0.354971
R126 VP.n113 VP.n112 0.354971
R127 VP VP.n113 0.26696
R128 VP.n31 VP.n28 0.189894
R129 VP.n35 VP.n28 0.189894
R130 VP.n36 VP.n35 0.189894
R131 VP.n37 VP.n36 0.189894
R132 VP.n37 VP.n26 0.189894
R133 VP.n41 VP.n26 0.189894
R134 VP.n42 VP.n41 0.189894
R135 VP.n42 VP.n24 0.189894
R136 VP.n46 VP.n24 0.189894
R137 VP.n47 VP.n46 0.189894
R138 VP.n48 VP.n47 0.189894
R139 VP.n48 VP.n22 0.189894
R140 VP.n52 VP.n22 0.189894
R141 VP.n53 VP.n52 0.189894
R142 VP.n54 VP.n53 0.189894
R143 VP.n54 VP.n20 0.189894
R144 VP.n58 VP.n20 0.189894
R145 VP.n59 VP.n58 0.189894
R146 VP.n60 VP.n59 0.189894
R147 VP.n60 VP.n18 0.189894
R148 VP.n64 VP.n18 0.189894
R149 VP.n67 VP.n15 0.189894
R150 VP.n71 VP.n15 0.189894
R151 VP.n72 VP.n71 0.189894
R152 VP.n73 VP.n72 0.189894
R153 VP.n73 VP.n13 0.189894
R154 VP.n77 VP.n13 0.189894
R155 VP.n78 VP.n77 0.189894
R156 VP.n79 VP.n78 0.189894
R157 VP.n79 VP.n11 0.189894
R158 VP.n83 VP.n11 0.189894
R159 VP.n84 VP.n83 0.189894
R160 VP.n85 VP.n84 0.189894
R161 VP.n85 VP.n9 0.189894
R162 VP.n89 VP.n9 0.189894
R163 VP.n90 VP.n89 0.189894
R164 VP.n90 VP.n7 0.189894
R165 VP.n94 VP.n7 0.189894
R166 VP.n95 VP.n94 0.189894
R167 VP.n96 VP.n95 0.189894
R168 VP.n96 VP.n5 0.189894
R169 VP.n100 VP.n5 0.189894
R170 VP.n101 VP.n100 0.189894
R171 VP.n102 VP.n101 0.189894
R172 VP.n102 VP.n3 0.189894
R173 VP.n106 VP.n3 0.189894
R174 VP.n107 VP.n106 0.189894
R175 VP.n108 VP.n107 0.189894
R176 VP.n108 VP.n1 0.189894
R177 VP.n112 VP.n1 0.189894
R178 VDD1.n1 VDD1.t7 109.017
R179 VDD1.n3 VDD1.t2 109.017
R180 VDD1.n5 VDD1.n4 101.453
R181 VDD1.n1 VDD1.n0 99.0832
R182 VDD1.n7 VDD1.n6 99.0831
R183 VDD1.n3 VDD1.n2 99.083
R184 VDD1.n7 VDD1.n5 45.4513
R185 VDD1.n6 VDD1.t1 6.70256
R186 VDD1.n6 VDD1.t8 6.70256
R187 VDD1.n0 VDD1.t3 6.70256
R188 VDD1.n0 VDD1.t0 6.70256
R189 VDD1.n4 VDD1.t6 6.70256
R190 VDD1.n4 VDD1.t9 6.70256
R191 VDD1.n2 VDD1.t5 6.70256
R192 VDD1.n2 VDD1.t4 6.70256
R193 VDD1 VDD1.n7 2.36688
R194 VDD1 VDD1.n1 0.866879
R195 VDD1.n5 VDD1.n3 0.753344
R196 VTAIL.n11 VTAIL.t7 89.1064
R197 VTAIL.n16 VTAIL.t9 89.1063
R198 VTAIL.n17 VTAIL.t6 89.1063
R199 VTAIL.n2 VTAIL.t10 89.1063
R200 VTAIL.n15 VTAIL.n14 82.4044
R201 VTAIL.n13 VTAIL.n12 82.4044
R202 VTAIL.n10 VTAIL.n9 82.4044
R203 VTAIL.n8 VTAIL.n7 82.4044
R204 VTAIL.n19 VTAIL.n18 82.4042
R205 VTAIL.n1 VTAIL.n0 82.4042
R206 VTAIL.n4 VTAIL.n3 82.4042
R207 VTAIL.n6 VTAIL.n5 82.4042
R208 VTAIL.n8 VTAIL.n6 23.0134
R209 VTAIL.n17 VTAIL.n16 19.7807
R210 VTAIL.n18 VTAIL.t0 6.70256
R211 VTAIL.n18 VTAIL.t8 6.70256
R212 VTAIL.n0 VTAIL.t4 6.70256
R213 VTAIL.n0 VTAIL.t3 6.70256
R214 VTAIL.n3 VTAIL.t15 6.70256
R215 VTAIL.n3 VTAIL.t16 6.70256
R216 VTAIL.n5 VTAIL.t11 6.70256
R217 VTAIL.n5 VTAIL.t14 6.70256
R218 VTAIL.n14 VTAIL.t12 6.70256
R219 VTAIL.n14 VTAIL.t18 6.70256
R220 VTAIL.n12 VTAIL.t13 6.70256
R221 VTAIL.n12 VTAIL.t17 6.70256
R222 VTAIL.n9 VTAIL.t2 6.70256
R223 VTAIL.n9 VTAIL.t1 6.70256
R224 VTAIL.n7 VTAIL.t5 6.70256
R225 VTAIL.n7 VTAIL.t19 6.70256
R226 VTAIL.n10 VTAIL.n8 3.23326
R227 VTAIL.n11 VTAIL.n10 3.23326
R228 VTAIL.n15 VTAIL.n13 3.23326
R229 VTAIL.n16 VTAIL.n15 3.23326
R230 VTAIL.n6 VTAIL.n4 3.23326
R231 VTAIL.n4 VTAIL.n2 3.23326
R232 VTAIL.n19 VTAIL.n17 3.23326
R233 VTAIL VTAIL.n1 2.48326
R234 VTAIL.n13 VTAIL.n11 2.08671
R235 VTAIL.n2 VTAIL.n1 2.08671
R236 VTAIL VTAIL.n19 0.7505
R237 B.n397 B.n144 585
R238 B.n396 B.n395 585
R239 B.n394 B.n145 585
R240 B.n393 B.n392 585
R241 B.n391 B.n146 585
R242 B.n390 B.n389 585
R243 B.n388 B.n147 585
R244 B.n387 B.n386 585
R245 B.n385 B.n148 585
R246 B.n384 B.n383 585
R247 B.n382 B.n149 585
R248 B.n381 B.n380 585
R249 B.n379 B.n150 585
R250 B.n378 B.n377 585
R251 B.n376 B.n151 585
R252 B.n375 B.n374 585
R253 B.n373 B.n152 585
R254 B.n372 B.n371 585
R255 B.n370 B.n153 585
R256 B.n369 B.n368 585
R257 B.n367 B.n154 585
R258 B.n366 B.n365 585
R259 B.n361 B.n155 585
R260 B.n360 B.n359 585
R261 B.n358 B.n156 585
R262 B.n357 B.n356 585
R263 B.n355 B.n157 585
R264 B.n354 B.n353 585
R265 B.n352 B.n158 585
R266 B.n351 B.n350 585
R267 B.n348 B.n159 585
R268 B.n347 B.n346 585
R269 B.n345 B.n162 585
R270 B.n344 B.n343 585
R271 B.n342 B.n163 585
R272 B.n341 B.n340 585
R273 B.n339 B.n164 585
R274 B.n338 B.n337 585
R275 B.n336 B.n165 585
R276 B.n335 B.n334 585
R277 B.n333 B.n166 585
R278 B.n332 B.n331 585
R279 B.n330 B.n167 585
R280 B.n329 B.n328 585
R281 B.n327 B.n168 585
R282 B.n326 B.n325 585
R283 B.n324 B.n169 585
R284 B.n323 B.n322 585
R285 B.n321 B.n170 585
R286 B.n320 B.n319 585
R287 B.n318 B.n171 585
R288 B.n399 B.n398 585
R289 B.n400 B.n143 585
R290 B.n402 B.n401 585
R291 B.n403 B.n142 585
R292 B.n405 B.n404 585
R293 B.n406 B.n141 585
R294 B.n408 B.n407 585
R295 B.n409 B.n140 585
R296 B.n411 B.n410 585
R297 B.n412 B.n139 585
R298 B.n414 B.n413 585
R299 B.n415 B.n138 585
R300 B.n417 B.n416 585
R301 B.n418 B.n137 585
R302 B.n420 B.n419 585
R303 B.n421 B.n136 585
R304 B.n423 B.n422 585
R305 B.n424 B.n135 585
R306 B.n426 B.n425 585
R307 B.n427 B.n134 585
R308 B.n429 B.n428 585
R309 B.n430 B.n133 585
R310 B.n432 B.n431 585
R311 B.n433 B.n132 585
R312 B.n435 B.n434 585
R313 B.n436 B.n131 585
R314 B.n438 B.n437 585
R315 B.n439 B.n130 585
R316 B.n441 B.n440 585
R317 B.n442 B.n129 585
R318 B.n444 B.n443 585
R319 B.n445 B.n128 585
R320 B.n447 B.n446 585
R321 B.n448 B.n127 585
R322 B.n450 B.n449 585
R323 B.n451 B.n126 585
R324 B.n453 B.n452 585
R325 B.n454 B.n125 585
R326 B.n456 B.n455 585
R327 B.n457 B.n124 585
R328 B.n459 B.n458 585
R329 B.n460 B.n123 585
R330 B.n462 B.n461 585
R331 B.n463 B.n122 585
R332 B.n465 B.n464 585
R333 B.n466 B.n121 585
R334 B.n468 B.n467 585
R335 B.n469 B.n120 585
R336 B.n471 B.n470 585
R337 B.n472 B.n119 585
R338 B.n474 B.n473 585
R339 B.n475 B.n118 585
R340 B.n477 B.n476 585
R341 B.n478 B.n117 585
R342 B.n480 B.n479 585
R343 B.n481 B.n116 585
R344 B.n483 B.n482 585
R345 B.n484 B.n115 585
R346 B.n486 B.n485 585
R347 B.n487 B.n114 585
R348 B.n489 B.n488 585
R349 B.n490 B.n113 585
R350 B.n492 B.n491 585
R351 B.n493 B.n112 585
R352 B.n495 B.n494 585
R353 B.n496 B.n111 585
R354 B.n498 B.n497 585
R355 B.n499 B.n110 585
R356 B.n501 B.n500 585
R357 B.n502 B.n109 585
R358 B.n504 B.n503 585
R359 B.n505 B.n108 585
R360 B.n507 B.n506 585
R361 B.n508 B.n107 585
R362 B.n510 B.n509 585
R363 B.n511 B.n106 585
R364 B.n513 B.n512 585
R365 B.n514 B.n105 585
R366 B.n516 B.n515 585
R367 B.n517 B.n104 585
R368 B.n519 B.n518 585
R369 B.n520 B.n103 585
R370 B.n522 B.n521 585
R371 B.n523 B.n102 585
R372 B.n525 B.n524 585
R373 B.n526 B.n101 585
R374 B.n528 B.n527 585
R375 B.n529 B.n100 585
R376 B.n531 B.n530 585
R377 B.n532 B.n99 585
R378 B.n534 B.n533 585
R379 B.n535 B.n98 585
R380 B.n537 B.n536 585
R381 B.n538 B.n97 585
R382 B.n540 B.n539 585
R383 B.n541 B.n96 585
R384 B.n543 B.n542 585
R385 B.n544 B.n95 585
R386 B.n546 B.n545 585
R387 B.n547 B.n94 585
R388 B.n549 B.n548 585
R389 B.n550 B.n93 585
R390 B.n552 B.n551 585
R391 B.n553 B.n92 585
R392 B.n555 B.n554 585
R393 B.n556 B.n91 585
R394 B.n558 B.n557 585
R395 B.n559 B.n90 585
R396 B.n561 B.n560 585
R397 B.n562 B.n89 585
R398 B.n564 B.n563 585
R399 B.n565 B.n88 585
R400 B.n567 B.n566 585
R401 B.n568 B.n87 585
R402 B.n570 B.n569 585
R403 B.n571 B.n86 585
R404 B.n573 B.n572 585
R405 B.n574 B.n85 585
R406 B.n576 B.n575 585
R407 B.n577 B.n84 585
R408 B.n579 B.n578 585
R409 B.n580 B.n83 585
R410 B.n582 B.n581 585
R411 B.n583 B.n82 585
R412 B.n585 B.n584 585
R413 B.n586 B.n81 585
R414 B.n588 B.n587 585
R415 B.n589 B.n80 585
R416 B.n591 B.n590 585
R417 B.n592 B.n79 585
R418 B.n594 B.n593 585
R419 B.n595 B.n78 585
R420 B.n597 B.n596 585
R421 B.n598 B.n77 585
R422 B.n600 B.n599 585
R423 B.n601 B.n76 585
R424 B.n603 B.n602 585
R425 B.n604 B.n75 585
R426 B.n606 B.n605 585
R427 B.n607 B.n74 585
R428 B.n609 B.n608 585
R429 B.n610 B.n73 585
R430 B.n612 B.n611 585
R431 B.n613 B.n72 585
R432 B.n615 B.n614 585
R433 B.n616 B.n71 585
R434 B.n618 B.n617 585
R435 B.n619 B.n70 585
R436 B.n621 B.n620 585
R437 B.n622 B.n69 585
R438 B.n700 B.n39 585
R439 B.n699 B.n698 585
R440 B.n697 B.n40 585
R441 B.n696 B.n695 585
R442 B.n694 B.n41 585
R443 B.n693 B.n692 585
R444 B.n691 B.n42 585
R445 B.n690 B.n689 585
R446 B.n688 B.n43 585
R447 B.n687 B.n686 585
R448 B.n685 B.n44 585
R449 B.n684 B.n683 585
R450 B.n682 B.n45 585
R451 B.n681 B.n680 585
R452 B.n679 B.n46 585
R453 B.n678 B.n677 585
R454 B.n676 B.n47 585
R455 B.n675 B.n674 585
R456 B.n673 B.n48 585
R457 B.n672 B.n671 585
R458 B.n670 B.n49 585
R459 B.n668 B.n667 585
R460 B.n666 B.n52 585
R461 B.n665 B.n664 585
R462 B.n663 B.n53 585
R463 B.n662 B.n661 585
R464 B.n660 B.n54 585
R465 B.n659 B.n658 585
R466 B.n657 B.n55 585
R467 B.n656 B.n655 585
R468 B.n654 B.n653 585
R469 B.n652 B.n59 585
R470 B.n651 B.n650 585
R471 B.n649 B.n60 585
R472 B.n648 B.n647 585
R473 B.n646 B.n61 585
R474 B.n645 B.n644 585
R475 B.n643 B.n62 585
R476 B.n642 B.n641 585
R477 B.n640 B.n63 585
R478 B.n639 B.n638 585
R479 B.n637 B.n64 585
R480 B.n636 B.n635 585
R481 B.n634 B.n65 585
R482 B.n633 B.n632 585
R483 B.n631 B.n66 585
R484 B.n630 B.n629 585
R485 B.n628 B.n67 585
R486 B.n627 B.n626 585
R487 B.n625 B.n68 585
R488 B.n624 B.n623 585
R489 B.n702 B.n701 585
R490 B.n703 B.n38 585
R491 B.n705 B.n704 585
R492 B.n706 B.n37 585
R493 B.n708 B.n707 585
R494 B.n709 B.n36 585
R495 B.n711 B.n710 585
R496 B.n712 B.n35 585
R497 B.n714 B.n713 585
R498 B.n715 B.n34 585
R499 B.n717 B.n716 585
R500 B.n718 B.n33 585
R501 B.n720 B.n719 585
R502 B.n721 B.n32 585
R503 B.n723 B.n722 585
R504 B.n724 B.n31 585
R505 B.n726 B.n725 585
R506 B.n727 B.n30 585
R507 B.n729 B.n728 585
R508 B.n730 B.n29 585
R509 B.n732 B.n731 585
R510 B.n733 B.n28 585
R511 B.n735 B.n734 585
R512 B.n736 B.n27 585
R513 B.n738 B.n737 585
R514 B.n739 B.n26 585
R515 B.n741 B.n740 585
R516 B.n742 B.n25 585
R517 B.n744 B.n743 585
R518 B.n745 B.n24 585
R519 B.n747 B.n746 585
R520 B.n748 B.n23 585
R521 B.n750 B.n749 585
R522 B.n751 B.n22 585
R523 B.n753 B.n752 585
R524 B.n754 B.n21 585
R525 B.n756 B.n755 585
R526 B.n757 B.n20 585
R527 B.n759 B.n758 585
R528 B.n760 B.n19 585
R529 B.n762 B.n761 585
R530 B.n763 B.n18 585
R531 B.n765 B.n764 585
R532 B.n766 B.n17 585
R533 B.n768 B.n767 585
R534 B.n769 B.n16 585
R535 B.n771 B.n770 585
R536 B.n772 B.n15 585
R537 B.n774 B.n773 585
R538 B.n775 B.n14 585
R539 B.n777 B.n776 585
R540 B.n778 B.n13 585
R541 B.n780 B.n779 585
R542 B.n781 B.n12 585
R543 B.n783 B.n782 585
R544 B.n784 B.n11 585
R545 B.n786 B.n785 585
R546 B.n787 B.n10 585
R547 B.n789 B.n788 585
R548 B.n790 B.n9 585
R549 B.n792 B.n791 585
R550 B.n793 B.n8 585
R551 B.n795 B.n794 585
R552 B.n796 B.n7 585
R553 B.n798 B.n797 585
R554 B.n799 B.n6 585
R555 B.n801 B.n800 585
R556 B.n802 B.n5 585
R557 B.n804 B.n803 585
R558 B.n805 B.n4 585
R559 B.n807 B.n806 585
R560 B.n808 B.n3 585
R561 B.n810 B.n809 585
R562 B.n811 B.n0 585
R563 B.n2 B.n1 585
R564 B.n209 B.n208 585
R565 B.n210 B.n207 585
R566 B.n212 B.n211 585
R567 B.n213 B.n206 585
R568 B.n215 B.n214 585
R569 B.n216 B.n205 585
R570 B.n218 B.n217 585
R571 B.n219 B.n204 585
R572 B.n221 B.n220 585
R573 B.n222 B.n203 585
R574 B.n224 B.n223 585
R575 B.n225 B.n202 585
R576 B.n227 B.n226 585
R577 B.n228 B.n201 585
R578 B.n230 B.n229 585
R579 B.n231 B.n200 585
R580 B.n233 B.n232 585
R581 B.n234 B.n199 585
R582 B.n236 B.n235 585
R583 B.n237 B.n198 585
R584 B.n239 B.n238 585
R585 B.n240 B.n197 585
R586 B.n242 B.n241 585
R587 B.n243 B.n196 585
R588 B.n245 B.n244 585
R589 B.n246 B.n195 585
R590 B.n248 B.n247 585
R591 B.n249 B.n194 585
R592 B.n251 B.n250 585
R593 B.n252 B.n193 585
R594 B.n254 B.n253 585
R595 B.n255 B.n192 585
R596 B.n257 B.n256 585
R597 B.n258 B.n191 585
R598 B.n260 B.n259 585
R599 B.n261 B.n190 585
R600 B.n263 B.n262 585
R601 B.n264 B.n189 585
R602 B.n266 B.n265 585
R603 B.n267 B.n188 585
R604 B.n269 B.n268 585
R605 B.n270 B.n187 585
R606 B.n272 B.n271 585
R607 B.n273 B.n186 585
R608 B.n275 B.n274 585
R609 B.n276 B.n185 585
R610 B.n278 B.n277 585
R611 B.n279 B.n184 585
R612 B.n281 B.n280 585
R613 B.n282 B.n183 585
R614 B.n284 B.n283 585
R615 B.n285 B.n182 585
R616 B.n287 B.n286 585
R617 B.n288 B.n181 585
R618 B.n290 B.n289 585
R619 B.n291 B.n180 585
R620 B.n293 B.n292 585
R621 B.n294 B.n179 585
R622 B.n296 B.n295 585
R623 B.n297 B.n178 585
R624 B.n299 B.n298 585
R625 B.n300 B.n177 585
R626 B.n302 B.n301 585
R627 B.n303 B.n176 585
R628 B.n305 B.n304 585
R629 B.n306 B.n175 585
R630 B.n308 B.n307 585
R631 B.n309 B.n174 585
R632 B.n311 B.n310 585
R633 B.n312 B.n173 585
R634 B.n314 B.n313 585
R635 B.n315 B.n172 585
R636 B.n317 B.n316 585
R637 B.n316 B.n171 444.452
R638 B.n398 B.n397 444.452
R639 B.n624 B.n69 444.452
R640 B.n702 B.n39 444.452
R641 B.n813 B.n812 256.663
R642 B.n160 B.t3 243.197
R643 B.n362 B.t0 243.197
R644 B.n56 B.t9 243.197
R645 B.n50 B.t6 243.197
R646 B.n812 B.n811 235.042
R647 B.n812 B.n2 235.042
R648 B.n362 B.t1 189.194
R649 B.n56 B.t11 189.194
R650 B.n160 B.t4 189.189
R651 B.n50 B.t8 189.189
R652 B.n320 B.n171 163.367
R653 B.n321 B.n320 163.367
R654 B.n322 B.n321 163.367
R655 B.n322 B.n169 163.367
R656 B.n326 B.n169 163.367
R657 B.n327 B.n326 163.367
R658 B.n328 B.n327 163.367
R659 B.n328 B.n167 163.367
R660 B.n332 B.n167 163.367
R661 B.n333 B.n332 163.367
R662 B.n334 B.n333 163.367
R663 B.n334 B.n165 163.367
R664 B.n338 B.n165 163.367
R665 B.n339 B.n338 163.367
R666 B.n340 B.n339 163.367
R667 B.n340 B.n163 163.367
R668 B.n344 B.n163 163.367
R669 B.n345 B.n344 163.367
R670 B.n346 B.n345 163.367
R671 B.n346 B.n159 163.367
R672 B.n351 B.n159 163.367
R673 B.n352 B.n351 163.367
R674 B.n353 B.n352 163.367
R675 B.n353 B.n157 163.367
R676 B.n357 B.n157 163.367
R677 B.n358 B.n357 163.367
R678 B.n359 B.n358 163.367
R679 B.n359 B.n155 163.367
R680 B.n366 B.n155 163.367
R681 B.n367 B.n366 163.367
R682 B.n368 B.n367 163.367
R683 B.n368 B.n153 163.367
R684 B.n372 B.n153 163.367
R685 B.n373 B.n372 163.367
R686 B.n374 B.n373 163.367
R687 B.n374 B.n151 163.367
R688 B.n378 B.n151 163.367
R689 B.n379 B.n378 163.367
R690 B.n380 B.n379 163.367
R691 B.n380 B.n149 163.367
R692 B.n384 B.n149 163.367
R693 B.n385 B.n384 163.367
R694 B.n386 B.n385 163.367
R695 B.n386 B.n147 163.367
R696 B.n390 B.n147 163.367
R697 B.n391 B.n390 163.367
R698 B.n392 B.n391 163.367
R699 B.n392 B.n145 163.367
R700 B.n396 B.n145 163.367
R701 B.n397 B.n396 163.367
R702 B.n620 B.n69 163.367
R703 B.n620 B.n619 163.367
R704 B.n619 B.n618 163.367
R705 B.n618 B.n71 163.367
R706 B.n614 B.n71 163.367
R707 B.n614 B.n613 163.367
R708 B.n613 B.n612 163.367
R709 B.n612 B.n73 163.367
R710 B.n608 B.n73 163.367
R711 B.n608 B.n607 163.367
R712 B.n607 B.n606 163.367
R713 B.n606 B.n75 163.367
R714 B.n602 B.n75 163.367
R715 B.n602 B.n601 163.367
R716 B.n601 B.n600 163.367
R717 B.n600 B.n77 163.367
R718 B.n596 B.n77 163.367
R719 B.n596 B.n595 163.367
R720 B.n595 B.n594 163.367
R721 B.n594 B.n79 163.367
R722 B.n590 B.n79 163.367
R723 B.n590 B.n589 163.367
R724 B.n589 B.n588 163.367
R725 B.n588 B.n81 163.367
R726 B.n584 B.n81 163.367
R727 B.n584 B.n583 163.367
R728 B.n583 B.n582 163.367
R729 B.n582 B.n83 163.367
R730 B.n578 B.n83 163.367
R731 B.n578 B.n577 163.367
R732 B.n577 B.n576 163.367
R733 B.n576 B.n85 163.367
R734 B.n572 B.n85 163.367
R735 B.n572 B.n571 163.367
R736 B.n571 B.n570 163.367
R737 B.n570 B.n87 163.367
R738 B.n566 B.n87 163.367
R739 B.n566 B.n565 163.367
R740 B.n565 B.n564 163.367
R741 B.n564 B.n89 163.367
R742 B.n560 B.n89 163.367
R743 B.n560 B.n559 163.367
R744 B.n559 B.n558 163.367
R745 B.n558 B.n91 163.367
R746 B.n554 B.n91 163.367
R747 B.n554 B.n553 163.367
R748 B.n553 B.n552 163.367
R749 B.n552 B.n93 163.367
R750 B.n548 B.n93 163.367
R751 B.n548 B.n547 163.367
R752 B.n547 B.n546 163.367
R753 B.n546 B.n95 163.367
R754 B.n542 B.n95 163.367
R755 B.n542 B.n541 163.367
R756 B.n541 B.n540 163.367
R757 B.n540 B.n97 163.367
R758 B.n536 B.n97 163.367
R759 B.n536 B.n535 163.367
R760 B.n535 B.n534 163.367
R761 B.n534 B.n99 163.367
R762 B.n530 B.n99 163.367
R763 B.n530 B.n529 163.367
R764 B.n529 B.n528 163.367
R765 B.n528 B.n101 163.367
R766 B.n524 B.n101 163.367
R767 B.n524 B.n523 163.367
R768 B.n523 B.n522 163.367
R769 B.n522 B.n103 163.367
R770 B.n518 B.n103 163.367
R771 B.n518 B.n517 163.367
R772 B.n517 B.n516 163.367
R773 B.n516 B.n105 163.367
R774 B.n512 B.n105 163.367
R775 B.n512 B.n511 163.367
R776 B.n511 B.n510 163.367
R777 B.n510 B.n107 163.367
R778 B.n506 B.n107 163.367
R779 B.n506 B.n505 163.367
R780 B.n505 B.n504 163.367
R781 B.n504 B.n109 163.367
R782 B.n500 B.n109 163.367
R783 B.n500 B.n499 163.367
R784 B.n499 B.n498 163.367
R785 B.n498 B.n111 163.367
R786 B.n494 B.n111 163.367
R787 B.n494 B.n493 163.367
R788 B.n493 B.n492 163.367
R789 B.n492 B.n113 163.367
R790 B.n488 B.n113 163.367
R791 B.n488 B.n487 163.367
R792 B.n487 B.n486 163.367
R793 B.n486 B.n115 163.367
R794 B.n482 B.n115 163.367
R795 B.n482 B.n481 163.367
R796 B.n481 B.n480 163.367
R797 B.n480 B.n117 163.367
R798 B.n476 B.n117 163.367
R799 B.n476 B.n475 163.367
R800 B.n475 B.n474 163.367
R801 B.n474 B.n119 163.367
R802 B.n470 B.n119 163.367
R803 B.n470 B.n469 163.367
R804 B.n469 B.n468 163.367
R805 B.n468 B.n121 163.367
R806 B.n464 B.n121 163.367
R807 B.n464 B.n463 163.367
R808 B.n463 B.n462 163.367
R809 B.n462 B.n123 163.367
R810 B.n458 B.n123 163.367
R811 B.n458 B.n457 163.367
R812 B.n457 B.n456 163.367
R813 B.n456 B.n125 163.367
R814 B.n452 B.n125 163.367
R815 B.n452 B.n451 163.367
R816 B.n451 B.n450 163.367
R817 B.n450 B.n127 163.367
R818 B.n446 B.n127 163.367
R819 B.n446 B.n445 163.367
R820 B.n445 B.n444 163.367
R821 B.n444 B.n129 163.367
R822 B.n440 B.n129 163.367
R823 B.n440 B.n439 163.367
R824 B.n439 B.n438 163.367
R825 B.n438 B.n131 163.367
R826 B.n434 B.n131 163.367
R827 B.n434 B.n433 163.367
R828 B.n433 B.n432 163.367
R829 B.n432 B.n133 163.367
R830 B.n428 B.n133 163.367
R831 B.n428 B.n427 163.367
R832 B.n427 B.n426 163.367
R833 B.n426 B.n135 163.367
R834 B.n422 B.n135 163.367
R835 B.n422 B.n421 163.367
R836 B.n421 B.n420 163.367
R837 B.n420 B.n137 163.367
R838 B.n416 B.n137 163.367
R839 B.n416 B.n415 163.367
R840 B.n415 B.n414 163.367
R841 B.n414 B.n139 163.367
R842 B.n410 B.n139 163.367
R843 B.n410 B.n409 163.367
R844 B.n409 B.n408 163.367
R845 B.n408 B.n141 163.367
R846 B.n404 B.n141 163.367
R847 B.n404 B.n403 163.367
R848 B.n403 B.n402 163.367
R849 B.n402 B.n143 163.367
R850 B.n398 B.n143 163.367
R851 B.n698 B.n39 163.367
R852 B.n698 B.n697 163.367
R853 B.n697 B.n696 163.367
R854 B.n696 B.n41 163.367
R855 B.n692 B.n41 163.367
R856 B.n692 B.n691 163.367
R857 B.n691 B.n690 163.367
R858 B.n690 B.n43 163.367
R859 B.n686 B.n43 163.367
R860 B.n686 B.n685 163.367
R861 B.n685 B.n684 163.367
R862 B.n684 B.n45 163.367
R863 B.n680 B.n45 163.367
R864 B.n680 B.n679 163.367
R865 B.n679 B.n678 163.367
R866 B.n678 B.n47 163.367
R867 B.n674 B.n47 163.367
R868 B.n674 B.n673 163.367
R869 B.n673 B.n672 163.367
R870 B.n672 B.n49 163.367
R871 B.n667 B.n49 163.367
R872 B.n667 B.n666 163.367
R873 B.n666 B.n665 163.367
R874 B.n665 B.n53 163.367
R875 B.n661 B.n53 163.367
R876 B.n661 B.n660 163.367
R877 B.n660 B.n659 163.367
R878 B.n659 B.n55 163.367
R879 B.n655 B.n55 163.367
R880 B.n655 B.n654 163.367
R881 B.n654 B.n59 163.367
R882 B.n650 B.n59 163.367
R883 B.n650 B.n649 163.367
R884 B.n649 B.n648 163.367
R885 B.n648 B.n61 163.367
R886 B.n644 B.n61 163.367
R887 B.n644 B.n643 163.367
R888 B.n643 B.n642 163.367
R889 B.n642 B.n63 163.367
R890 B.n638 B.n63 163.367
R891 B.n638 B.n637 163.367
R892 B.n637 B.n636 163.367
R893 B.n636 B.n65 163.367
R894 B.n632 B.n65 163.367
R895 B.n632 B.n631 163.367
R896 B.n631 B.n630 163.367
R897 B.n630 B.n67 163.367
R898 B.n626 B.n67 163.367
R899 B.n626 B.n625 163.367
R900 B.n625 B.n624 163.367
R901 B.n703 B.n702 163.367
R902 B.n704 B.n703 163.367
R903 B.n704 B.n37 163.367
R904 B.n708 B.n37 163.367
R905 B.n709 B.n708 163.367
R906 B.n710 B.n709 163.367
R907 B.n710 B.n35 163.367
R908 B.n714 B.n35 163.367
R909 B.n715 B.n714 163.367
R910 B.n716 B.n715 163.367
R911 B.n716 B.n33 163.367
R912 B.n720 B.n33 163.367
R913 B.n721 B.n720 163.367
R914 B.n722 B.n721 163.367
R915 B.n722 B.n31 163.367
R916 B.n726 B.n31 163.367
R917 B.n727 B.n726 163.367
R918 B.n728 B.n727 163.367
R919 B.n728 B.n29 163.367
R920 B.n732 B.n29 163.367
R921 B.n733 B.n732 163.367
R922 B.n734 B.n733 163.367
R923 B.n734 B.n27 163.367
R924 B.n738 B.n27 163.367
R925 B.n739 B.n738 163.367
R926 B.n740 B.n739 163.367
R927 B.n740 B.n25 163.367
R928 B.n744 B.n25 163.367
R929 B.n745 B.n744 163.367
R930 B.n746 B.n745 163.367
R931 B.n746 B.n23 163.367
R932 B.n750 B.n23 163.367
R933 B.n751 B.n750 163.367
R934 B.n752 B.n751 163.367
R935 B.n752 B.n21 163.367
R936 B.n756 B.n21 163.367
R937 B.n757 B.n756 163.367
R938 B.n758 B.n757 163.367
R939 B.n758 B.n19 163.367
R940 B.n762 B.n19 163.367
R941 B.n763 B.n762 163.367
R942 B.n764 B.n763 163.367
R943 B.n764 B.n17 163.367
R944 B.n768 B.n17 163.367
R945 B.n769 B.n768 163.367
R946 B.n770 B.n769 163.367
R947 B.n770 B.n15 163.367
R948 B.n774 B.n15 163.367
R949 B.n775 B.n774 163.367
R950 B.n776 B.n775 163.367
R951 B.n776 B.n13 163.367
R952 B.n780 B.n13 163.367
R953 B.n781 B.n780 163.367
R954 B.n782 B.n781 163.367
R955 B.n782 B.n11 163.367
R956 B.n786 B.n11 163.367
R957 B.n787 B.n786 163.367
R958 B.n788 B.n787 163.367
R959 B.n788 B.n9 163.367
R960 B.n792 B.n9 163.367
R961 B.n793 B.n792 163.367
R962 B.n794 B.n793 163.367
R963 B.n794 B.n7 163.367
R964 B.n798 B.n7 163.367
R965 B.n799 B.n798 163.367
R966 B.n800 B.n799 163.367
R967 B.n800 B.n5 163.367
R968 B.n804 B.n5 163.367
R969 B.n805 B.n804 163.367
R970 B.n806 B.n805 163.367
R971 B.n806 B.n3 163.367
R972 B.n810 B.n3 163.367
R973 B.n811 B.n810 163.367
R974 B.n208 B.n2 163.367
R975 B.n208 B.n207 163.367
R976 B.n212 B.n207 163.367
R977 B.n213 B.n212 163.367
R978 B.n214 B.n213 163.367
R979 B.n214 B.n205 163.367
R980 B.n218 B.n205 163.367
R981 B.n219 B.n218 163.367
R982 B.n220 B.n219 163.367
R983 B.n220 B.n203 163.367
R984 B.n224 B.n203 163.367
R985 B.n225 B.n224 163.367
R986 B.n226 B.n225 163.367
R987 B.n226 B.n201 163.367
R988 B.n230 B.n201 163.367
R989 B.n231 B.n230 163.367
R990 B.n232 B.n231 163.367
R991 B.n232 B.n199 163.367
R992 B.n236 B.n199 163.367
R993 B.n237 B.n236 163.367
R994 B.n238 B.n237 163.367
R995 B.n238 B.n197 163.367
R996 B.n242 B.n197 163.367
R997 B.n243 B.n242 163.367
R998 B.n244 B.n243 163.367
R999 B.n244 B.n195 163.367
R1000 B.n248 B.n195 163.367
R1001 B.n249 B.n248 163.367
R1002 B.n250 B.n249 163.367
R1003 B.n250 B.n193 163.367
R1004 B.n254 B.n193 163.367
R1005 B.n255 B.n254 163.367
R1006 B.n256 B.n255 163.367
R1007 B.n256 B.n191 163.367
R1008 B.n260 B.n191 163.367
R1009 B.n261 B.n260 163.367
R1010 B.n262 B.n261 163.367
R1011 B.n262 B.n189 163.367
R1012 B.n266 B.n189 163.367
R1013 B.n267 B.n266 163.367
R1014 B.n268 B.n267 163.367
R1015 B.n268 B.n187 163.367
R1016 B.n272 B.n187 163.367
R1017 B.n273 B.n272 163.367
R1018 B.n274 B.n273 163.367
R1019 B.n274 B.n185 163.367
R1020 B.n278 B.n185 163.367
R1021 B.n279 B.n278 163.367
R1022 B.n280 B.n279 163.367
R1023 B.n280 B.n183 163.367
R1024 B.n284 B.n183 163.367
R1025 B.n285 B.n284 163.367
R1026 B.n286 B.n285 163.367
R1027 B.n286 B.n181 163.367
R1028 B.n290 B.n181 163.367
R1029 B.n291 B.n290 163.367
R1030 B.n292 B.n291 163.367
R1031 B.n292 B.n179 163.367
R1032 B.n296 B.n179 163.367
R1033 B.n297 B.n296 163.367
R1034 B.n298 B.n297 163.367
R1035 B.n298 B.n177 163.367
R1036 B.n302 B.n177 163.367
R1037 B.n303 B.n302 163.367
R1038 B.n304 B.n303 163.367
R1039 B.n304 B.n175 163.367
R1040 B.n308 B.n175 163.367
R1041 B.n309 B.n308 163.367
R1042 B.n310 B.n309 163.367
R1043 B.n310 B.n173 163.367
R1044 B.n314 B.n173 163.367
R1045 B.n315 B.n314 163.367
R1046 B.n316 B.n315 163.367
R1047 B.n363 B.t2 116.466
R1048 B.n57 B.t10 116.466
R1049 B.n161 B.t5 116.462
R1050 B.n51 B.t7 116.462
R1051 B.n161 B.n160 72.7278
R1052 B.n363 B.n362 72.7278
R1053 B.n57 B.n56 72.7278
R1054 B.n51 B.n50 72.7278
R1055 B.n349 B.n161 59.5399
R1056 B.n364 B.n363 59.5399
R1057 B.n58 B.n57 59.5399
R1058 B.n669 B.n51 59.5399
R1059 B.n701 B.n700 28.8785
R1060 B.n623 B.n622 28.8785
R1061 B.n318 B.n317 28.8785
R1062 B.n399 B.n144 28.8785
R1063 B B.n813 18.0485
R1064 B.n701 B.n38 10.6151
R1065 B.n705 B.n38 10.6151
R1066 B.n706 B.n705 10.6151
R1067 B.n707 B.n706 10.6151
R1068 B.n707 B.n36 10.6151
R1069 B.n711 B.n36 10.6151
R1070 B.n712 B.n711 10.6151
R1071 B.n713 B.n712 10.6151
R1072 B.n713 B.n34 10.6151
R1073 B.n717 B.n34 10.6151
R1074 B.n718 B.n717 10.6151
R1075 B.n719 B.n718 10.6151
R1076 B.n719 B.n32 10.6151
R1077 B.n723 B.n32 10.6151
R1078 B.n724 B.n723 10.6151
R1079 B.n725 B.n724 10.6151
R1080 B.n725 B.n30 10.6151
R1081 B.n729 B.n30 10.6151
R1082 B.n730 B.n729 10.6151
R1083 B.n731 B.n730 10.6151
R1084 B.n731 B.n28 10.6151
R1085 B.n735 B.n28 10.6151
R1086 B.n736 B.n735 10.6151
R1087 B.n737 B.n736 10.6151
R1088 B.n737 B.n26 10.6151
R1089 B.n741 B.n26 10.6151
R1090 B.n742 B.n741 10.6151
R1091 B.n743 B.n742 10.6151
R1092 B.n743 B.n24 10.6151
R1093 B.n747 B.n24 10.6151
R1094 B.n748 B.n747 10.6151
R1095 B.n749 B.n748 10.6151
R1096 B.n749 B.n22 10.6151
R1097 B.n753 B.n22 10.6151
R1098 B.n754 B.n753 10.6151
R1099 B.n755 B.n754 10.6151
R1100 B.n755 B.n20 10.6151
R1101 B.n759 B.n20 10.6151
R1102 B.n760 B.n759 10.6151
R1103 B.n761 B.n760 10.6151
R1104 B.n761 B.n18 10.6151
R1105 B.n765 B.n18 10.6151
R1106 B.n766 B.n765 10.6151
R1107 B.n767 B.n766 10.6151
R1108 B.n767 B.n16 10.6151
R1109 B.n771 B.n16 10.6151
R1110 B.n772 B.n771 10.6151
R1111 B.n773 B.n772 10.6151
R1112 B.n773 B.n14 10.6151
R1113 B.n777 B.n14 10.6151
R1114 B.n778 B.n777 10.6151
R1115 B.n779 B.n778 10.6151
R1116 B.n779 B.n12 10.6151
R1117 B.n783 B.n12 10.6151
R1118 B.n784 B.n783 10.6151
R1119 B.n785 B.n784 10.6151
R1120 B.n785 B.n10 10.6151
R1121 B.n789 B.n10 10.6151
R1122 B.n790 B.n789 10.6151
R1123 B.n791 B.n790 10.6151
R1124 B.n791 B.n8 10.6151
R1125 B.n795 B.n8 10.6151
R1126 B.n796 B.n795 10.6151
R1127 B.n797 B.n796 10.6151
R1128 B.n797 B.n6 10.6151
R1129 B.n801 B.n6 10.6151
R1130 B.n802 B.n801 10.6151
R1131 B.n803 B.n802 10.6151
R1132 B.n803 B.n4 10.6151
R1133 B.n807 B.n4 10.6151
R1134 B.n808 B.n807 10.6151
R1135 B.n809 B.n808 10.6151
R1136 B.n809 B.n0 10.6151
R1137 B.n700 B.n699 10.6151
R1138 B.n699 B.n40 10.6151
R1139 B.n695 B.n40 10.6151
R1140 B.n695 B.n694 10.6151
R1141 B.n694 B.n693 10.6151
R1142 B.n693 B.n42 10.6151
R1143 B.n689 B.n42 10.6151
R1144 B.n689 B.n688 10.6151
R1145 B.n688 B.n687 10.6151
R1146 B.n687 B.n44 10.6151
R1147 B.n683 B.n44 10.6151
R1148 B.n683 B.n682 10.6151
R1149 B.n682 B.n681 10.6151
R1150 B.n681 B.n46 10.6151
R1151 B.n677 B.n46 10.6151
R1152 B.n677 B.n676 10.6151
R1153 B.n676 B.n675 10.6151
R1154 B.n675 B.n48 10.6151
R1155 B.n671 B.n48 10.6151
R1156 B.n671 B.n670 10.6151
R1157 B.n668 B.n52 10.6151
R1158 B.n664 B.n52 10.6151
R1159 B.n664 B.n663 10.6151
R1160 B.n663 B.n662 10.6151
R1161 B.n662 B.n54 10.6151
R1162 B.n658 B.n54 10.6151
R1163 B.n658 B.n657 10.6151
R1164 B.n657 B.n656 10.6151
R1165 B.n653 B.n652 10.6151
R1166 B.n652 B.n651 10.6151
R1167 B.n651 B.n60 10.6151
R1168 B.n647 B.n60 10.6151
R1169 B.n647 B.n646 10.6151
R1170 B.n646 B.n645 10.6151
R1171 B.n645 B.n62 10.6151
R1172 B.n641 B.n62 10.6151
R1173 B.n641 B.n640 10.6151
R1174 B.n640 B.n639 10.6151
R1175 B.n639 B.n64 10.6151
R1176 B.n635 B.n64 10.6151
R1177 B.n635 B.n634 10.6151
R1178 B.n634 B.n633 10.6151
R1179 B.n633 B.n66 10.6151
R1180 B.n629 B.n66 10.6151
R1181 B.n629 B.n628 10.6151
R1182 B.n628 B.n627 10.6151
R1183 B.n627 B.n68 10.6151
R1184 B.n623 B.n68 10.6151
R1185 B.n622 B.n621 10.6151
R1186 B.n621 B.n70 10.6151
R1187 B.n617 B.n70 10.6151
R1188 B.n617 B.n616 10.6151
R1189 B.n616 B.n615 10.6151
R1190 B.n615 B.n72 10.6151
R1191 B.n611 B.n72 10.6151
R1192 B.n611 B.n610 10.6151
R1193 B.n610 B.n609 10.6151
R1194 B.n609 B.n74 10.6151
R1195 B.n605 B.n74 10.6151
R1196 B.n605 B.n604 10.6151
R1197 B.n604 B.n603 10.6151
R1198 B.n603 B.n76 10.6151
R1199 B.n599 B.n76 10.6151
R1200 B.n599 B.n598 10.6151
R1201 B.n598 B.n597 10.6151
R1202 B.n597 B.n78 10.6151
R1203 B.n593 B.n78 10.6151
R1204 B.n593 B.n592 10.6151
R1205 B.n592 B.n591 10.6151
R1206 B.n591 B.n80 10.6151
R1207 B.n587 B.n80 10.6151
R1208 B.n587 B.n586 10.6151
R1209 B.n586 B.n585 10.6151
R1210 B.n585 B.n82 10.6151
R1211 B.n581 B.n82 10.6151
R1212 B.n581 B.n580 10.6151
R1213 B.n580 B.n579 10.6151
R1214 B.n579 B.n84 10.6151
R1215 B.n575 B.n84 10.6151
R1216 B.n575 B.n574 10.6151
R1217 B.n574 B.n573 10.6151
R1218 B.n573 B.n86 10.6151
R1219 B.n569 B.n86 10.6151
R1220 B.n569 B.n568 10.6151
R1221 B.n568 B.n567 10.6151
R1222 B.n567 B.n88 10.6151
R1223 B.n563 B.n88 10.6151
R1224 B.n563 B.n562 10.6151
R1225 B.n562 B.n561 10.6151
R1226 B.n561 B.n90 10.6151
R1227 B.n557 B.n90 10.6151
R1228 B.n557 B.n556 10.6151
R1229 B.n556 B.n555 10.6151
R1230 B.n555 B.n92 10.6151
R1231 B.n551 B.n92 10.6151
R1232 B.n551 B.n550 10.6151
R1233 B.n550 B.n549 10.6151
R1234 B.n549 B.n94 10.6151
R1235 B.n545 B.n94 10.6151
R1236 B.n545 B.n544 10.6151
R1237 B.n544 B.n543 10.6151
R1238 B.n543 B.n96 10.6151
R1239 B.n539 B.n96 10.6151
R1240 B.n539 B.n538 10.6151
R1241 B.n538 B.n537 10.6151
R1242 B.n537 B.n98 10.6151
R1243 B.n533 B.n98 10.6151
R1244 B.n533 B.n532 10.6151
R1245 B.n532 B.n531 10.6151
R1246 B.n531 B.n100 10.6151
R1247 B.n527 B.n100 10.6151
R1248 B.n527 B.n526 10.6151
R1249 B.n526 B.n525 10.6151
R1250 B.n525 B.n102 10.6151
R1251 B.n521 B.n102 10.6151
R1252 B.n521 B.n520 10.6151
R1253 B.n520 B.n519 10.6151
R1254 B.n519 B.n104 10.6151
R1255 B.n515 B.n104 10.6151
R1256 B.n515 B.n514 10.6151
R1257 B.n514 B.n513 10.6151
R1258 B.n513 B.n106 10.6151
R1259 B.n509 B.n106 10.6151
R1260 B.n509 B.n508 10.6151
R1261 B.n508 B.n507 10.6151
R1262 B.n507 B.n108 10.6151
R1263 B.n503 B.n108 10.6151
R1264 B.n503 B.n502 10.6151
R1265 B.n502 B.n501 10.6151
R1266 B.n501 B.n110 10.6151
R1267 B.n497 B.n110 10.6151
R1268 B.n497 B.n496 10.6151
R1269 B.n496 B.n495 10.6151
R1270 B.n495 B.n112 10.6151
R1271 B.n491 B.n112 10.6151
R1272 B.n491 B.n490 10.6151
R1273 B.n490 B.n489 10.6151
R1274 B.n489 B.n114 10.6151
R1275 B.n485 B.n114 10.6151
R1276 B.n485 B.n484 10.6151
R1277 B.n484 B.n483 10.6151
R1278 B.n483 B.n116 10.6151
R1279 B.n479 B.n116 10.6151
R1280 B.n479 B.n478 10.6151
R1281 B.n478 B.n477 10.6151
R1282 B.n477 B.n118 10.6151
R1283 B.n473 B.n118 10.6151
R1284 B.n473 B.n472 10.6151
R1285 B.n472 B.n471 10.6151
R1286 B.n471 B.n120 10.6151
R1287 B.n467 B.n120 10.6151
R1288 B.n467 B.n466 10.6151
R1289 B.n466 B.n465 10.6151
R1290 B.n465 B.n122 10.6151
R1291 B.n461 B.n122 10.6151
R1292 B.n461 B.n460 10.6151
R1293 B.n460 B.n459 10.6151
R1294 B.n459 B.n124 10.6151
R1295 B.n455 B.n124 10.6151
R1296 B.n455 B.n454 10.6151
R1297 B.n454 B.n453 10.6151
R1298 B.n453 B.n126 10.6151
R1299 B.n449 B.n126 10.6151
R1300 B.n449 B.n448 10.6151
R1301 B.n448 B.n447 10.6151
R1302 B.n447 B.n128 10.6151
R1303 B.n443 B.n128 10.6151
R1304 B.n443 B.n442 10.6151
R1305 B.n442 B.n441 10.6151
R1306 B.n441 B.n130 10.6151
R1307 B.n437 B.n130 10.6151
R1308 B.n437 B.n436 10.6151
R1309 B.n436 B.n435 10.6151
R1310 B.n435 B.n132 10.6151
R1311 B.n431 B.n132 10.6151
R1312 B.n431 B.n430 10.6151
R1313 B.n430 B.n429 10.6151
R1314 B.n429 B.n134 10.6151
R1315 B.n425 B.n134 10.6151
R1316 B.n425 B.n424 10.6151
R1317 B.n424 B.n423 10.6151
R1318 B.n423 B.n136 10.6151
R1319 B.n419 B.n136 10.6151
R1320 B.n419 B.n418 10.6151
R1321 B.n418 B.n417 10.6151
R1322 B.n417 B.n138 10.6151
R1323 B.n413 B.n138 10.6151
R1324 B.n413 B.n412 10.6151
R1325 B.n412 B.n411 10.6151
R1326 B.n411 B.n140 10.6151
R1327 B.n407 B.n140 10.6151
R1328 B.n407 B.n406 10.6151
R1329 B.n406 B.n405 10.6151
R1330 B.n405 B.n142 10.6151
R1331 B.n401 B.n142 10.6151
R1332 B.n401 B.n400 10.6151
R1333 B.n400 B.n399 10.6151
R1334 B.n209 B.n1 10.6151
R1335 B.n210 B.n209 10.6151
R1336 B.n211 B.n210 10.6151
R1337 B.n211 B.n206 10.6151
R1338 B.n215 B.n206 10.6151
R1339 B.n216 B.n215 10.6151
R1340 B.n217 B.n216 10.6151
R1341 B.n217 B.n204 10.6151
R1342 B.n221 B.n204 10.6151
R1343 B.n222 B.n221 10.6151
R1344 B.n223 B.n222 10.6151
R1345 B.n223 B.n202 10.6151
R1346 B.n227 B.n202 10.6151
R1347 B.n228 B.n227 10.6151
R1348 B.n229 B.n228 10.6151
R1349 B.n229 B.n200 10.6151
R1350 B.n233 B.n200 10.6151
R1351 B.n234 B.n233 10.6151
R1352 B.n235 B.n234 10.6151
R1353 B.n235 B.n198 10.6151
R1354 B.n239 B.n198 10.6151
R1355 B.n240 B.n239 10.6151
R1356 B.n241 B.n240 10.6151
R1357 B.n241 B.n196 10.6151
R1358 B.n245 B.n196 10.6151
R1359 B.n246 B.n245 10.6151
R1360 B.n247 B.n246 10.6151
R1361 B.n247 B.n194 10.6151
R1362 B.n251 B.n194 10.6151
R1363 B.n252 B.n251 10.6151
R1364 B.n253 B.n252 10.6151
R1365 B.n253 B.n192 10.6151
R1366 B.n257 B.n192 10.6151
R1367 B.n258 B.n257 10.6151
R1368 B.n259 B.n258 10.6151
R1369 B.n259 B.n190 10.6151
R1370 B.n263 B.n190 10.6151
R1371 B.n264 B.n263 10.6151
R1372 B.n265 B.n264 10.6151
R1373 B.n265 B.n188 10.6151
R1374 B.n269 B.n188 10.6151
R1375 B.n270 B.n269 10.6151
R1376 B.n271 B.n270 10.6151
R1377 B.n271 B.n186 10.6151
R1378 B.n275 B.n186 10.6151
R1379 B.n276 B.n275 10.6151
R1380 B.n277 B.n276 10.6151
R1381 B.n277 B.n184 10.6151
R1382 B.n281 B.n184 10.6151
R1383 B.n282 B.n281 10.6151
R1384 B.n283 B.n282 10.6151
R1385 B.n283 B.n182 10.6151
R1386 B.n287 B.n182 10.6151
R1387 B.n288 B.n287 10.6151
R1388 B.n289 B.n288 10.6151
R1389 B.n289 B.n180 10.6151
R1390 B.n293 B.n180 10.6151
R1391 B.n294 B.n293 10.6151
R1392 B.n295 B.n294 10.6151
R1393 B.n295 B.n178 10.6151
R1394 B.n299 B.n178 10.6151
R1395 B.n300 B.n299 10.6151
R1396 B.n301 B.n300 10.6151
R1397 B.n301 B.n176 10.6151
R1398 B.n305 B.n176 10.6151
R1399 B.n306 B.n305 10.6151
R1400 B.n307 B.n306 10.6151
R1401 B.n307 B.n174 10.6151
R1402 B.n311 B.n174 10.6151
R1403 B.n312 B.n311 10.6151
R1404 B.n313 B.n312 10.6151
R1405 B.n313 B.n172 10.6151
R1406 B.n317 B.n172 10.6151
R1407 B.n319 B.n318 10.6151
R1408 B.n319 B.n170 10.6151
R1409 B.n323 B.n170 10.6151
R1410 B.n324 B.n323 10.6151
R1411 B.n325 B.n324 10.6151
R1412 B.n325 B.n168 10.6151
R1413 B.n329 B.n168 10.6151
R1414 B.n330 B.n329 10.6151
R1415 B.n331 B.n330 10.6151
R1416 B.n331 B.n166 10.6151
R1417 B.n335 B.n166 10.6151
R1418 B.n336 B.n335 10.6151
R1419 B.n337 B.n336 10.6151
R1420 B.n337 B.n164 10.6151
R1421 B.n341 B.n164 10.6151
R1422 B.n342 B.n341 10.6151
R1423 B.n343 B.n342 10.6151
R1424 B.n343 B.n162 10.6151
R1425 B.n347 B.n162 10.6151
R1426 B.n348 B.n347 10.6151
R1427 B.n350 B.n158 10.6151
R1428 B.n354 B.n158 10.6151
R1429 B.n355 B.n354 10.6151
R1430 B.n356 B.n355 10.6151
R1431 B.n356 B.n156 10.6151
R1432 B.n360 B.n156 10.6151
R1433 B.n361 B.n360 10.6151
R1434 B.n365 B.n361 10.6151
R1435 B.n369 B.n154 10.6151
R1436 B.n370 B.n369 10.6151
R1437 B.n371 B.n370 10.6151
R1438 B.n371 B.n152 10.6151
R1439 B.n375 B.n152 10.6151
R1440 B.n376 B.n375 10.6151
R1441 B.n377 B.n376 10.6151
R1442 B.n377 B.n150 10.6151
R1443 B.n381 B.n150 10.6151
R1444 B.n382 B.n381 10.6151
R1445 B.n383 B.n382 10.6151
R1446 B.n383 B.n148 10.6151
R1447 B.n387 B.n148 10.6151
R1448 B.n388 B.n387 10.6151
R1449 B.n389 B.n388 10.6151
R1450 B.n389 B.n146 10.6151
R1451 B.n393 B.n146 10.6151
R1452 B.n394 B.n393 10.6151
R1453 B.n395 B.n394 10.6151
R1454 B.n395 B.n144 10.6151
R1455 B.n813 B.n0 8.11757
R1456 B.n813 B.n1 8.11757
R1457 B.n669 B.n668 6.5566
R1458 B.n656 B.n58 6.5566
R1459 B.n350 B.n349 6.5566
R1460 B.n365 B.n364 6.5566
R1461 B.n670 B.n669 4.05904
R1462 B.n653 B.n58 4.05904
R1463 B.n349 B.n348 4.05904
R1464 B.n364 B.n154 4.05904
R1465 VN.n96 VN.n95 161.3
R1466 VN.n94 VN.n50 161.3
R1467 VN.n93 VN.n92 161.3
R1468 VN.n91 VN.n51 161.3
R1469 VN.n90 VN.n89 161.3
R1470 VN.n88 VN.n52 161.3
R1471 VN.n87 VN.n86 161.3
R1472 VN.n85 VN.n53 161.3
R1473 VN.n84 VN.n83 161.3
R1474 VN.n82 VN.n54 161.3
R1475 VN.n81 VN.n80 161.3
R1476 VN.n79 VN.n55 161.3
R1477 VN.n78 VN.n77 161.3
R1478 VN.n76 VN.n56 161.3
R1479 VN.n75 VN.n74 161.3
R1480 VN.n73 VN.n72 161.3
R1481 VN.n71 VN.n58 161.3
R1482 VN.n70 VN.n69 161.3
R1483 VN.n68 VN.n59 161.3
R1484 VN.n67 VN.n66 161.3
R1485 VN.n65 VN.n60 161.3
R1486 VN.n64 VN.n63 161.3
R1487 VN.n47 VN.n46 161.3
R1488 VN.n45 VN.n1 161.3
R1489 VN.n44 VN.n43 161.3
R1490 VN.n42 VN.n2 161.3
R1491 VN.n41 VN.n40 161.3
R1492 VN.n39 VN.n3 161.3
R1493 VN.n38 VN.n37 161.3
R1494 VN.n36 VN.n4 161.3
R1495 VN.n35 VN.n34 161.3
R1496 VN.n33 VN.n5 161.3
R1497 VN.n32 VN.n31 161.3
R1498 VN.n30 VN.n6 161.3
R1499 VN.n29 VN.n28 161.3
R1500 VN.n27 VN.n7 161.3
R1501 VN.n26 VN.n25 161.3
R1502 VN.n24 VN.n23 161.3
R1503 VN.n22 VN.n9 161.3
R1504 VN.n21 VN.n20 161.3
R1505 VN.n19 VN.n10 161.3
R1506 VN.n18 VN.n17 161.3
R1507 VN.n16 VN.n11 161.3
R1508 VN.n15 VN.n14 161.3
R1509 VN.n48 VN.n0 77.8339
R1510 VN.n97 VN.n49 77.8339
R1511 VN.n62 VN.t5 67.9562
R1512 VN.n13 VN.t7 67.9562
R1513 VN.n17 VN.n10 52.6342
R1514 VN.n32 VN.n6 52.6342
R1515 VN.n40 VN.n2 52.6342
R1516 VN.n66 VN.n59 52.6342
R1517 VN.n81 VN.n55 52.6342
R1518 VN.n89 VN.n51 52.6342
R1519 VN VN.n97 52.4261
R1520 VN.n13 VN.n12 50.1549
R1521 VN.n62 VN.n61 50.1549
R1522 VN.n4 VN.t4 34.1774
R1523 VN.n12 VN.t9 34.1774
R1524 VN.n8 VN.t3 34.1774
R1525 VN.n0 VN.t8 34.1774
R1526 VN.n53 VN.t6 34.1774
R1527 VN.n61 VN.t0 34.1774
R1528 VN.n57 VN.t1 34.1774
R1529 VN.n49 VN.t2 34.1774
R1530 VN.n21 VN.n10 28.3526
R1531 VN.n28 VN.n6 28.3526
R1532 VN.n44 VN.n2 28.3526
R1533 VN.n70 VN.n59 28.3526
R1534 VN.n77 VN.n55 28.3526
R1535 VN.n93 VN.n51 28.3526
R1536 VN.n15 VN.n12 24.4675
R1537 VN.n16 VN.n15 24.4675
R1538 VN.n17 VN.n16 24.4675
R1539 VN.n22 VN.n21 24.4675
R1540 VN.n23 VN.n22 24.4675
R1541 VN.n27 VN.n26 24.4675
R1542 VN.n28 VN.n27 24.4675
R1543 VN.n33 VN.n32 24.4675
R1544 VN.n34 VN.n33 24.4675
R1545 VN.n34 VN.n4 24.4675
R1546 VN.n38 VN.n4 24.4675
R1547 VN.n39 VN.n38 24.4675
R1548 VN.n40 VN.n39 24.4675
R1549 VN.n45 VN.n44 24.4675
R1550 VN.n46 VN.n45 24.4675
R1551 VN.n66 VN.n65 24.4675
R1552 VN.n65 VN.n64 24.4675
R1553 VN.n64 VN.n61 24.4675
R1554 VN.n77 VN.n76 24.4675
R1555 VN.n76 VN.n75 24.4675
R1556 VN.n72 VN.n71 24.4675
R1557 VN.n71 VN.n70 24.4675
R1558 VN.n89 VN.n88 24.4675
R1559 VN.n88 VN.n87 24.4675
R1560 VN.n87 VN.n53 24.4675
R1561 VN.n83 VN.n53 24.4675
R1562 VN.n83 VN.n82 24.4675
R1563 VN.n82 VN.n81 24.4675
R1564 VN.n95 VN.n94 24.4675
R1565 VN.n94 VN.n93 24.4675
R1566 VN.n23 VN.n8 12.234
R1567 VN.n26 VN.n8 12.234
R1568 VN.n46 VN.n0 12.234
R1569 VN.n75 VN.n57 12.234
R1570 VN.n72 VN.n57 12.234
R1571 VN.n95 VN.n49 12.234
R1572 VN.n63 VN.n62 3.07682
R1573 VN.n14 VN.n13 3.07682
R1574 VN.n97 VN.n96 0.354971
R1575 VN.n48 VN.n47 0.354971
R1576 VN VN.n48 0.26696
R1577 VN.n96 VN.n50 0.189894
R1578 VN.n92 VN.n50 0.189894
R1579 VN.n92 VN.n91 0.189894
R1580 VN.n91 VN.n90 0.189894
R1581 VN.n90 VN.n52 0.189894
R1582 VN.n86 VN.n52 0.189894
R1583 VN.n86 VN.n85 0.189894
R1584 VN.n85 VN.n84 0.189894
R1585 VN.n84 VN.n54 0.189894
R1586 VN.n80 VN.n54 0.189894
R1587 VN.n80 VN.n79 0.189894
R1588 VN.n79 VN.n78 0.189894
R1589 VN.n78 VN.n56 0.189894
R1590 VN.n74 VN.n56 0.189894
R1591 VN.n74 VN.n73 0.189894
R1592 VN.n73 VN.n58 0.189894
R1593 VN.n69 VN.n58 0.189894
R1594 VN.n69 VN.n68 0.189894
R1595 VN.n68 VN.n67 0.189894
R1596 VN.n67 VN.n60 0.189894
R1597 VN.n63 VN.n60 0.189894
R1598 VN.n14 VN.n11 0.189894
R1599 VN.n18 VN.n11 0.189894
R1600 VN.n19 VN.n18 0.189894
R1601 VN.n20 VN.n19 0.189894
R1602 VN.n20 VN.n9 0.189894
R1603 VN.n24 VN.n9 0.189894
R1604 VN.n25 VN.n24 0.189894
R1605 VN.n25 VN.n7 0.189894
R1606 VN.n29 VN.n7 0.189894
R1607 VN.n30 VN.n29 0.189894
R1608 VN.n31 VN.n30 0.189894
R1609 VN.n31 VN.n5 0.189894
R1610 VN.n35 VN.n5 0.189894
R1611 VN.n36 VN.n35 0.189894
R1612 VN.n37 VN.n36 0.189894
R1613 VN.n37 VN.n3 0.189894
R1614 VN.n41 VN.n3 0.189894
R1615 VN.n42 VN.n41 0.189894
R1616 VN.n43 VN.n42 0.189894
R1617 VN.n43 VN.n1 0.189894
R1618 VN.n47 VN.n1 0.189894
R1619 VDD2.n1 VDD2.t2 109.017
R1620 VDD2.n4 VDD2.t7 105.785
R1621 VDD2.n3 VDD2.n2 101.453
R1622 VDD2 VDD2.n7 101.45
R1623 VDD2.n6 VDD2.n5 99.0832
R1624 VDD2.n1 VDD2.n0 99.083
R1625 VDD2.n4 VDD2.n3 43.2519
R1626 VDD2.n7 VDD2.t9 6.70256
R1627 VDD2.n7 VDD2.t4 6.70256
R1628 VDD2.n5 VDD2.t3 6.70256
R1629 VDD2.n5 VDD2.t8 6.70256
R1630 VDD2.n2 VDD2.t5 6.70256
R1631 VDD2.n2 VDD2.t1 6.70256
R1632 VDD2.n0 VDD2.t0 6.70256
R1633 VDD2.n0 VDD2.t6 6.70256
R1634 VDD2.n6 VDD2.n4 3.23326
R1635 VDD2 VDD2.n6 0.866879
R1636 VDD2.n3 VDD2.n1 0.753344
C0 VTAIL VDD2 7.91104f
C1 VN VP 8.2841f
C2 B w_n5470_n1938# 9.939429f
C3 VDD2 w_n5470_n1938# 2.79514f
C4 VN B 1.46569f
C5 VN VDD2 4.850049f
C6 VTAIL w_n5470_n1938# 2.34605f
C7 VDD1 VP 5.37941f
C8 VTAIL VN 6.4591f
C9 VDD1 B 2.22533f
C10 VDD1 VDD2 2.70803f
C11 VN w_n5470_n1938# 11.838f
C12 VTAIL VDD1 7.85263f
C13 VDD1 w_n5470_n1938# 2.60928f
C14 VP B 2.67194f
C15 VDD1 VN 0.159077f
C16 VP VDD2 0.692262f
C17 VDD2 B 2.37532f
C18 VTAIL VP 6.473259f
C19 VP w_n5470_n1938# 12.5526f
C20 VTAIL B 2.3389f
C21 VDD2 VSUBS 2.417474f
C22 VDD1 VSUBS 2.146155f
C23 VTAIL VSUBS 0.742813f
C24 VN VSUBS 8.80811f
C25 VP VSUBS 4.659995f
C26 B VSUBS 5.424492f
C27 w_n5470_n1938# VSUBS 0.132921p
C28 VDD2.t2 VSUBS 1.21576f
C29 VDD2.t0 VSUBS 0.140518f
C30 VDD2.t6 VSUBS 0.140518f
C31 VDD2.n0 VSUBS 0.872811f
C32 VDD2.n1 VSUBS 2.02402f
C33 VDD2.t5 VSUBS 0.140518f
C34 VDD2.t1 VSUBS 0.140518f
C35 VDD2.n2 VSUBS 0.90164f
C36 VDD2.n3 VSUBS 4.50763f
C37 VDD2.t7 VSUBS 1.18537f
C38 VDD2.n4 VSUBS 4.46551f
C39 VDD2.t3 VSUBS 0.140518f
C40 VDD2.t8 VSUBS 0.140518f
C41 VDD2.n5 VSUBS 0.872815f
C42 VDD2.n6 VSUBS 1.0418f
C43 VDD2.t9 VSUBS 0.140518f
C44 VDD2.t4 VSUBS 0.140518f
C45 VDD2.n7 VSUBS 0.901589f
C46 VN.t8 VSUBS 1.50511f
C47 VN.n0 VSUBS 0.706669f
C48 VN.n1 VSUBS 0.034768f
C49 VN.n2 VSUBS 0.035775f
C50 VN.n3 VSUBS 0.034768f
C51 VN.t4 VSUBS 1.50511f
C52 VN.n4 VSUBS 0.603527f
C53 VN.n5 VSUBS 0.034768f
C54 VN.n6 VSUBS 0.035775f
C55 VN.n7 VSUBS 0.034768f
C56 VN.t3 VSUBS 1.50511f
C57 VN.n8 VSUBS 0.57072f
C58 VN.n9 VSUBS 0.034768f
C59 VN.n10 VSUBS 0.035775f
C60 VN.n11 VSUBS 0.034768f
C61 VN.t9 VSUBS 1.50511f
C62 VN.n12 VSUBS 0.708341f
C63 VN.t7 VSUBS 1.9178f
C64 VN.n13 VSUBS 0.669579f
C65 VN.n14 VSUBS 0.424646f
C66 VN.n15 VSUBS 0.064799f
C67 VN.n16 VSUBS 0.064799f
C68 VN.n17 VSUBS 0.06206f
C69 VN.n18 VSUBS 0.034768f
C70 VN.n19 VSUBS 0.034768f
C71 VN.n20 VSUBS 0.034768f
C72 VN.n21 VSUBS 0.068482f
C73 VN.n22 VSUBS 0.064799f
C74 VN.n23 VSUBS 0.048803f
C75 VN.n24 VSUBS 0.034768f
C76 VN.n25 VSUBS 0.034768f
C77 VN.n26 VSUBS 0.048803f
C78 VN.n27 VSUBS 0.064799f
C79 VN.n28 VSUBS 0.068482f
C80 VN.n29 VSUBS 0.034768f
C81 VN.n30 VSUBS 0.034768f
C82 VN.n31 VSUBS 0.034768f
C83 VN.n32 VSUBS 0.06206f
C84 VN.n33 VSUBS 0.064799f
C85 VN.n34 VSUBS 0.064799f
C86 VN.n35 VSUBS 0.034768f
C87 VN.n36 VSUBS 0.034768f
C88 VN.n37 VSUBS 0.034768f
C89 VN.n38 VSUBS 0.064799f
C90 VN.n39 VSUBS 0.064799f
C91 VN.n40 VSUBS 0.06206f
C92 VN.n41 VSUBS 0.034768f
C93 VN.n42 VSUBS 0.034768f
C94 VN.n43 VSUBS 0.034768f
C95 VN.n44 VSUBS 0.068482f
C96 VN.n45 VSUBS 0.064799f
C97 VN.n46 VSUBS 0.048803f
C98 VN.n47 VSUBS 0.056115f
C99 VN.n48 VSUBS 0.089246f
C100 VN.t2 VSUBS 1.50511f
C101 VN.n49 VSUBS 0.706669f
C102 VN.n50 VSUBS 0.034768f
C103 VN.n51 VSUBS 0.035775f
C104 VN.n52 VSUBS 0.034768f
C105 VN.t6 VSUBS 1.50511f
C106 VN.n53 VSUBS 0.603527f
C107 VN.n54 VSUBS 0.034768f
C108 VN.n55 VSUBS 0.035775f
C109 VN.n56 VSUBS 0.034768f
C110 VN.t1 VSUBS 1.50511f
C111 VN.n57 VSUBS 0.57072f
C112 VN.n58 VSUBS 0.034768f
C113 VN.n59 VSUBS 0.035775f
C114 VN.n60 VSUBS 0.034768f
C115 VN.t0 VSUBS 1.50511f
C116 VN.n61 VSUBS 0.708341f
C117 VN.t5 VSUBS 1.9178f
C118 VN.n62 VSUBS 0.669579f
C119 VN.n63 VSUBS 0.424646f
C120 VN.n64 VSUBS 0.064799f
C121 VN.n65 VSUBS 0.064799f
C122 VN.n66 VSUBS 0.06206f
C123 VN.n67 VSUBS 0.034768f
C124 VN.n68 VSUBS 0.034768f
C125 VN.n69 VSUBS 0.034768f
C126 VN.n70 VSUBS 0.068482f
C127 VN.n71 VSUBS 0.064799f
C128 VN.n72 VSUBS 0.048803f
C129 VN.n73 VSUBS 0.034768f
C130 VN.n74 VSUBS 0.034768f
C131 VN.n75 VSUBS 0.048803f
C132 VN.n76 VSUBS 0.064799f
C133 VN.n77 VSUBS 0.068482f
C134 VN.n78 VSUBS 0.034768f
C135 VN.n79 VSUBS 0.034768f
C136 VN.n80 VSUBS 0.034768f
C137 VN.n81 VSUBS 0.06206f
C138 VN.n82 VSUBS 0.064799f
C139 VN.n83 VSUBS 0.064799f
C140 VN.n84 VSUBS 0.034768f
C141 VN.n85 VSUBS 0.034768f
C142 VN.n86 VSUBS 0.034768f
C143 VN.n87 VSUBS 0.064799f
C144 VN.n88 VSUBS 0.064799f
C145 VN.n89 VSUBS 0.06206f
C146 VN.n90 VSUBS 0.034768f
C147 VN.n91 VSUBS 0.034768f
C148 VN.n92 VSUBS 0.034768f
C149 VN.n93 VSUBS 0.068482f
C150 VN.n94 VSUBS 0.064799f
C151 VN.n95 VSUBS 0.048803f
C152 VN.n96 VSUBS 0.056115f
C153 VN.n97 VSUBS 2.12587f
C154 B.n0 VSUBS 0.011028f
C155 B.n1 VSUBS 0.011028f
C156 B.n2 VSUBS 0.01631f
C157 B.n3 VSUBS 0.012498f
C158 B.n4 VSUBS 0.012498f
C159 B.n5 VSUBS 0.012498f
C160 B.n6 VSUBS 0.012498f
C161 B.n7 VSUBS 0.012498f
C162 B.n8 VSUBS 0.012498f
C163 B.n9 VSUBS 0.012498f
C164 B.n10 VSUBS 0.012498f
C165 B.n11 VSUBS 0.012498f
C166 B.n12 VSUBS 0.012498f
C167 B.n13 VSUBS 0.012498f
C168 B.n14 VSUBS 0.012498f
C169 B.n15 VSUBS 0.012498f
C170 B.n16 VSUBS 0.012498f
C171 B.n17 VSUBS 0.012498f
C172 B.n18 VSUBS 0.012498f
C173 B.n19 VSUBS 0.012498f
C174 B.n20 VSUBS 0.012498f
C175 B.n21 VSUBS 0.012498f
C176 B.n22 VSUBS 0.012498f
C177 B.n23 VSUBS 0.012498f
C178 B.n24 VSUBS 0.012498f
C179 B.n25 VSUBS 0.012498f
C180 B.n26 VSUBS 0.012498f
C181 B.n27 VSUBS 0.012498f
C182 B.n28 VSUBS 0.012498f
C183 B.n29 VSUBS 0.012498f
C184 B.n30 VSUBS 0.012498f
C185 B.n31 VSUBS 0.012498f
C186 B.n32 VSUBS 0.012498f
C187 B.n33 VSUBS 0.012498f
C188 B.n34 VSUBS 0.012498f
C189 B.n35 VSUBS 0.012498f
C190 B.n36 VSUBS 0.012498f
C191 B.n37 VSUBS 0.012498f
C192 B.n38 VSUBS 0.012498f
C193 B.n39 VSUBS 0.027691f
C194 B.n40 VSUBS 0.012498f
C195 B.n41 VSUBS 0.012498f
C196 B.n42 VSUBS 0.012498f
C197 B.n43 VSUBS 0.012498f
C198 B.n44 VSUBS 0.012498f
C199 B.n45 VSUBS 0.012498f
C200 B.n46 VSUBS 0.012498f
C201 B.n47 VSUBS 0.012498f
C202 B.n48 VSUBS 0.012498f
C203 B.n49 VSUBS 0.012498f
C204 B.t7 VSUBS 0.240133f
C205 B.t8 VSUBS 0.283561f
C206 B.t6 VSUBS 1.42897f
C207 B.n50 VSUBS 0.192977f
C208 B.n51 VSUBS 0.130797f
C209 B.n52 VSUBS 0.012498f
C210 B.n53 VSUBS 0.012498f
C211 B.n54 VSUBS 0.012498f
C212 B.n55 VSUBS 0.012498f
C213 B.t10 VSUBS 0.240133f
C214 B.t11 VSUBS 0.28356f
C215 B.t9 VSUBS 1.42897f
C216 B.n56 VSUBS 0.192978f
C217 B.n57 VSUBS 0.130797f
C218 B.n58 VSUBS 0.028957f
C219 B.n59 VSUBS 0.012498f
C220 B.n60 VSUBS 0.012498f
C221 B.n61 VSUBS 0.012498f
C222 B.n62 VSUBS 0.012498f
C223 B.n63 VSUBS 0.012498f
C224 B.n64 VSUBS 0.012498f
C225 B.n65 VSUBS 0.012498f
C226 B.n66 VSUBS 0.012498f
C227 B.n67 VSUBS 0.012498f
C228 B.n68 VSUBS 0.012498f
C229 B.n69 VSUBS 0.026346f
C230 B.n70 VSUBS 0.012498f
C231 B.n71 VSUBS 0.012498f
C232 B.n72 VSUBS 0.012498f
C233 B.n73 VSUBS 0.012498f
C234 B.n74 VSUBS 0.012498f
C235 B.n75 VSUBS 0.012498f
C236 B.n76 VSUBS 0.012498f
C237 B.n77 VSUBS 0.012498f
C238 B.n78 VSUBS 0.012498f
C239 B.n79 VSUBS 0.012498f
C240 B.n80 VSUBS 0.012498f
C241 B.n81 VSUBS 0.012498f
C242 B.n82 VSUBS 0.012498f
C243 B.n83 VSUBS 0.012498f
C244 B.n84 VSUBS 0.012498f
C245 B.n85 VSUBS 0.012498f
C246 B.n86 VSUBS 0.012498f
C247 B.n87 VSUBS 0.012498f
C248 B.n88 VSUBS 0.012498f
C249 B.n89 VSUBS 0.012498f
C250 B.n90 VSUBS 0.012498f
C251 B.n91 VSUBS 0.012498f
C252 B.n92 VSUBS 0.012498f
C253 B.n93 VSUBS 0.012498f
C254 B.n94 VSUBS 0.012498f
C255 B.n95 VSUBS 0.012498f
C256 B.n96 VSUBS 0.012498f
C257 B.n97 VSUBS 0.012498f
C258 B.n98 VSUBS 0.012498f
C259 B.n99 VSUBS 0.012498f
C260 B.n100 VSUBS 0.012498f
C261 B.n101 VSUBS 0.012498f
C262 B.n102 VSUBS 0.012498f
C263 B.n103 VSUBS 0.012498f
C264 B.n104 VSUBS 0.012498f
C265 B.n105 VSUBS 0.012498f
C266 B.n106 VSUBS 0.012498f
C267 B.n107 VSUBS 0.012498f
C268 B.n108 VSUBS 0.012498f
C269 B.n109 VSUBS 0.012498f
C270 B.n110 VSUBS 0.012498f
C271 B.n111 VSUBS 0.012498f
C272 B.n112 VSUBS 0.012498f
C273 B.n113 VSUBS 0.012498f
C274 B.n114 VSUBS 0.012498f
C275 B.n115 VSUBS 0.012498f
C276 B.n116 VSUBS 0.012498f
C277 B.n117 VSUBS 0.012498f
C278 B.n118 VSUBS 0.012498f
C279 B.n119 VSUBS 0.012498f
C280 B.n120 VSUBS 0.012498f
C281 B.n121 VSUBS 0.012498f
C282 B.n122 VSUBS 0.012498f
C283 B.n123 VSUBS 0.012498f
C284 B.n124 VSUBS 0.012498f
C285 B.n125 VSUBS 0.012498f
C286 B.n126 VSUBS 0.012498f
C287 B.n127 VSUBS 0.012498f
C288 B.n128 VSUBS 0.012498f
C289 B.n129 VSUBS 0.012498f
C290 B.n130 VSUBS 0.012498f
C291 B.n131 VSUBS 0.012498f
C292 B.n132 VSUBS 0.012498f
C293 B.n133 VSUBS 0.012498f
C294 B.n134 VSUBS 0.012498f
C295 B.n135 VSUBS 0.012498f
C296 B.n136 VSUBS 0.012498f
C297 B.n137 VSUBS 0.012498f
C298 B.n138 VSUBS 0.012498f
C299 B.n139 VSUBS 0.012498f
C300 B.n140 VSUBS 0.012498f
C301 B.n141 VSUBS 0.012498f
C302 B.n142 VSUBS 0.012498f
C303 B.n143 VSUBS 0.012498f
C304 B.n144 VSUBS 0.026021f
C305 B.n145 VSUBS 0.012498f
C306 B.n146 VSUBS 0.012498f
C307 B.n147 VSUBS 0.012498f
C308 B.n148 VSUBS 0.012498f
C309 B.n149 VSUBS 0.012498f
C310 B.n150 VSUBS 0.012498f
C311 B.n151 VSUBS 0.012498f
C312 B.n152 VSUBS 0.012498f
C313 B.n153 VSUBS 0.012498f
C314 B.n154 VSUBS 0.008639f
C315 B.n155 VSUBS 0.012498f
C316 B.n156 VSUBS 0.012498f
C317 B.n157 VSUBS 0.012498f
C318 B.n158 VSUBS 0.012498f
C319 B.n159 VSUBS 0.012498f
C320 B.t5 VSUBS 0.240133f
C321 B.t4 VSUBS 0.283561f
C322 B.t3 VSUBS 1.42897f
C323 B.n160 VSUBS 0.192977f
C324 B.n161 VSUBS 0.130797f
C325 B.n162 VSUBS 0.012498f
C326 B.n163 VSUBS 0.012498f
C327 B.n164 VSUBS 0.012498f
C328 B.n165 VSUBS 0.012498f
C329 B.n166 VSUBS 0.012498f
C330 B.n167 VSUBS 0.012498f
C331 B.n168 VSUBS 0.012498f
C332 B.n169 VSUBS 0.012498f
C333 B.n170 VSUBS 0.012498f
C334 B.n171 VSUBS 0.027691f
C335 B.n172 VSUBS 0.012498f
C336 B.n173 VSUBS 0.012498f
C337 B.n174 VSUBS 0.012498f
C338 B.n175 VSUBS 0.012498f
C339 B.n176 VSUBS 0.012498f
C340 B.n177 VSUBS 0.012498f
C341 B.n178 VSUBS 0.012498f
C342 B.n179 VSUBS 0.012498f
C343 B.n180 VSUBS 0.012498f
C344 B.n181 VSUBS 0.012498f
C345 B.n182 VSUBS 0.012498f
C346 B.n183 VSUBS 0.012498f
C347 B.n184 VSUBS 0.012498f
C348 B.n185 VSUBS 0.012498f
C349 B.n186 VSUBS 0.012498f
C350 B.n187 VSUBS 0.012498f
C351 B.n188 VSUBS 0.012498f
C352 B.n189 VSUBS 0.012498f
C353 B.n190 VSUBS 0.012498f
C354 B.n191 VSUBS 0.012498f
C355 B.n192 VSUBS 0.012498f
C356 B.n193 VSUBS 0.012498f
C357 B.n194 VSUBS 0.012498f
C358 B.n195 VSUBS 0.012498f
C359 B.n196 VSUBS 0.012498f
C360 B.n197 VSUBS 0.012498f
C361 B.n198 VSUBS 0.012498f
C362 B.n199 VSUBS 0.012498f
C363 B.n200 VSUBS 0.012498f
C364 B.n201 VSUBS 0.012498f
C365 B.n202 VSUBS 0.012498f
C366 B.n203 VSUBS 0.012498f
C367 B.n204 VSUBS 0.012498f
C368 B.n205 VSUBS 0.012498f
C369 B.n206 VSUBS 0.012498f
C370 B.n207 VSUBS 0.012498f
C371 B.n208 VSUBS 0.012498f
C372 B.n209 VSUBS 0.012498f
C373 B.n210 VSUBS 0.012498f
C374 B.n211 VSUBS 0.012498f
C375 B.n212 VSUBS 0.012498f
C376 B.n213 VSUBS 0.012498f
C377 B.n214 VSUBS 0.012498f
C378 B.n215 VSUBS 0.012498f
C379 B.n216 VSUBS 0.012498f
C380 B.n217 VSUBS 0.012498f
C381 B.n218 VSUBS 0.012498f
C382 B.n219 VSUBS 0.012498f
C383 B.n220 VSUBS 0.012498f
C384 B.n221 VSUBS 0.012498f
C385 B.n222 VSUBS 0.012498f
C386 B.n223 VSUBS 0.012498f
C387 B.n224 VSUBS 0.012498f
C388 B.n225 VSUBS 0.012498f
C389 B.n226 VSUBS 0.012498f
C390 B.n227 VSUBS 0.012498f
C391 B.n228 VSUBS 0.012498f
C392 B.n229 VSUBS 0.012498f
C393 B.n230 VSUBS 0.012498f
C394 B.n231 VSUBS 0.012498f
C395 B.n232 VSUBS 0.012498f
C396 B.n233 VSUBS 0.012498f
C397 B.n234 VSUBS 0.012498f
C398 B.n235 VSUBS 0.012498f
C399 B.n236 VSUBS 0.012498f
C400 B.n237 VSUBS 0.012498f
C401 B.n238 VSUBS 0.012498f
C402 B.n239 VSUBS 0.012498f
C403 B.n240 VSUBS 0.012498f
C404 B.n241 VSUBS 0.012498f
C405 B.n242 VSUBS 0.012498f
C406 B.n243 VSUBS 0.012498f
C407 B.n244 VSUBS 0.012498f
C408 B.n245 VSUBS 0.012498f
C409 B.n246 VSUBS 0.012498f
C410 B.n247 VSUBS 0.012498f
C411 B.n248 VSUBS 0.012498f
C412 B.n249 VSUBS 0.012498f
C413 B.n250 VSUBS 0.012498f
C414 B.n251 VSUBS 0.012498f
C415 B.n252 VSUBS 0.012498f
C416 B.n253 VSUBS 0.012498f
C417 B.n254 VSUBS 0.012498f
C418 B.n255 VSUBS 0.012498f
C419 B.n256 VSUBS 0.012498f
C420 B.n257 VSUBS 0.012498f
C421 B.n258 VSUBS 0.012498f
C422 B.n259 VSUBS 0.012498f
C423 B.n260 VSUBS 0.012498f
C424 B.n261 VSUBS 0.012498f
C425 B.n262 VSUBS 0.012498f
C426 B.n263 VSUBS 0.012498f
C427 B.n264 VSUBS 0.012498f
C428 B.n265 VSUBS 0.012498f
C429 B.n266 VSUBS 0.012498f
C430 B.n267 VSUBS 0.012498f
C431 B.n268 VSUBS 0.012498f
C432 B.n269 VSUBS 0.012498f
C433 B.n270 VSUBS 0.012498f
C434 B.n271 VSUBS 0.012498f
C435 B.n272 VSUBS 0.012498f
C436 B.n273 VSUBS 0.012498f
C437 B.n274 VSUBS 0.012498f
C438 B.n275 VSUBS 0.012498f
C439 B.n276 VSUBS 0.012498f
C440 B.n277 VSUBS 0.012498f
C441 B.n278 VSUBS 0.012498f
C442 B.n279 VSUBS 0.012498f
C443 B.n280 VSUBS 0.012498f
C444 B.n281 VSUBS 0.012498f
C445 B.n282 VSUBS 0.012498f
C446 B.n283 VSUBS 0.012498f
C447 B.n284 VSUBS 0.012498f
C448 B.n285 VSUBS 0.012498f
C449 B.n286 VSUBS 0.012498f
C450 B.n287 VSUBS 0.012498f
C451 B.n288 VSUBS 0.012498f
C452 B.n289 VSUBS 0.012498f
C453 B.n290 VSUBS 0.012498f
C454 B.n291 VSUBS 0.012498f
C455 B.n292 VSUBS 0.012498f
C456 B.n293 VSUBS 0.012498f
C457 B.n294 VSUBS 0.012498f
C458 B.n295 VSUBS 0.012498f
C459 B.n296 VSUBS 0.012498f
C460 B.n297 VSUBS 0.012498f
C461 B.n298 VSUBS 0.012498f
C462 B.n299 VSUBS 0.012498f
C463 B.n300 VSUBS 0.012498f
C464 B.n301 VSUBS 0.012498f
C465 B.n302 VSUBS 0.012498f
C466 B.n303 VSUBS 0.012498f
C467 B.n304 VSUBS 0.012498f
C468 B.n305 VSUBS 0.012498f
C469 B.n306 VSUBS 0.012498f
C470 B.n307 VSUBS 0.012498f
C471 B.n308 VSUBS 0.012498f
C472 B.n309 VSUBS 0.012498f
C473 B.n310 VSUBS 0.012498f
C474 B.n311 VSUBS 0.012498f
C475 B.n312 VSUBS 0.012498f
C476 B.n313 VSUBS 0.012498f
C477 B.n314 VSUBS 0.012498f
C478 B.n315 VSUBS 0.012498f
C479 B.n316 VSUBS 0.026346f
C480 B.n317 VSUBS 0.026346f
C481 B.n318 VSUBS 0.027691f
C482 B.n319 VSUBS 0.012498f
C483 B.n320 VSUBS 0.012498f
C484 B.n321 VSUBS 0.012498f
C485 B.n322 VSUBS 0.012498f
C486 B.n323 VSUBS 0.012498f
C487 B.n324 VSUBS 0.012498f
C488 B.n325 VSUBS 0.012498f
C489 B.n326 VSUBS 0.012498f
C490 B.n327 VSUBS 0.012498f
C491 B.n328 VSUBS 0.012498f
C492 B.n329 VSUBS 0.012498f
C493 B.n330 VSUBS 0.012498f
C494 B.n331 VSUBS 0.012498f
C495 B.n332 VSUBS 0.012498f
C496 B.n333 VSUBS 0.012498f
C497 B.n334 VSUBS 0.012498f
C498 B.n335 VSUBS 0.012498f
C499 B.n336 VSUBS 0.012498f
C500 B.n337 VSUBS 0.012498f
C501 B.n338 VSUBS 0.012498f
C502 B.n339 VSUBS 0.012498f
C503 B.n340 VSUBS 0.012498f
C504 B.n341 VSUBS 0.012498f
C505 B.n342 VSUBS 0.012498f
C506 B.n343 VSUBS 0.012498f
C507 B.n344 VSUBS 0.012498f
C508 B.n345 VSUBS 0.012498f
C509 B.n346 VSUBS 0.012498f
C510 B.n347 VSUBS 0.012498f
C511 B.n348 VSUBS 0.008639f
C512 B.n349 VSUBS 0.028957f
C513 B.n350 VSUBS 0.010109f
C514 B.n351 VSUBS 0.012498f
C515 B.n352 VSUBS 0.012498f
C516 B.n353 VSUBS 0.012498f
C517 B.n354 VSUBS 0.012498f
C518 B.n355 VSUBS 0.012498f
C519 B.n356 VSUBS 0.012498f
C520 B.n357 VSUBS 0.012498f
C521 B.n358 VSUBS 0.012498f
C522 B.n359 VSUBS 0.012498f
C523 B.n360 VSUBS 0.012498f
C524 B.n361 VSUBS 0.012498f
C525 B.t2 VSUBS 0.240133f
C526 B.t1 VSUBS 0.28356f
C527 B.t0 VSUBS 1.42897f
C528 B.n362 VSUBS 0.192978f
C529 B.n363 VSUBS 0.130797f
C530 B.n364 VSUBS 0.028957f
C531 B.n365 VSUBS 0.010109f
C532 B.n366 VSUBS 0.012498f
C533 B.n367 VSUBS 0.012498f
C534 B.n368 VSUBS 0.012498f
C535 B.n369 VSUBS 0.012498f
C536 B.n370 VSUBS 0.012498f
C537 B.n371 VSUBS 0.012498f
C538 B.n372 VSUBS 0.012498f
C539 B.n373 VSUBS 0.012498f
C540 B.n374 VSUBS 0.012498f
C541 B.n375 VSUBS 0.012498f
C542 B.n376 VSUBS 0.012498f
C543 B.n377 VSUBS 0.012498f
C544 B.n378 VSUBS 0.012498f
C545 B.n379 VSUBS 0.012498f
C546 B.n380 VSUBS 0.012498f
C547 B.n381 VSUBS 0.012498f
C548 B.n382 VSUBS 0.012498f
C549 B.n383 VSUBS 0.012498f
C550 B.n384 VSUBS 0.012498f
C551 B.n385 VSUBS 0.012498f
C552 B.n386 VSUBS 0.012498f
C553 B.n387 VSUBS 0.012498f
C554 B.n388 VSUBS 0.012498f
C555 B.n389 VSUBS 0.012498f
C556 B.n390 VSUBS 0.012498f
C557 B.n391 VSUBS 0.012498f
C558 B.n392 VSUBS 0.012498f
C559 B.n393 VSUBS 0.012498f
C560 B.n394 VSUBS 0.012498f
C561 B.n395 VSUBS 0.012498f
C562 B.n396 VSUBS 0.012498f
C563 B.n397 VSUBS 0.027691f
C564 B.n398 VSUBS 0.026346f
C565 B.n399 VSUBS 0.028017f
C566 B.n400 VSUBS 0.012498f
C567 B.n401 VSUBS 0.012498f
C568 B.n402 VSUBS 0.012498f
C569 B.n403 VSUBS 0.012498f
C570 B.n404 VSUBS 0.012498f
C571 B.n405 VSUBS 0.012498f
C572 B.n406 VSUBS 0.012498f
C573 B.n407 VSUBS 0.012498f
C574 B.n408 VSUBS 0.012498f
C575 B.n409 VSUBS 0.012498f
C576 B.n410 VSUBS 0.012498f
C577 B.n411 VSUBS 0.012498f
C578 B.n412 VSUBS 0.012498f
C579 B.n413 VSUBS 0.012498f
C580 B.n414 VSUBS 0.012498f
C581 B.n415 VSUBS 0.012498f
C582 B.n416 VSUBS 0.012498f
C583 B.n417 VSUBS 0.012498f
C584 B.n418 VSUBS 0.012498f
C585 B.n419 VSUBS 0.012498f
C586 B.n420 VSUBS 0.012498f
C587 B.n421 VSUBS 0.012498f
C588 B.n422 VSUBS 0.012498f
C589 B.n423 VSUBS 0.012498f
C590 B.n424 VSUBS 0.012498f
C591 B.n425 VSUBS 0.012498f
C592 B.n426 VSUBS 0.012498f
C593 B.n427 VSUBS 0.012498f
C594 B.n428 VSUBS 0.012498f
C595 B.n429 VSUBS 0.012498f
C596 B.n430 VSUBS 0.012498f
C597 B.n431 VSUBS 0.012498f
C598 B.n432 VSUBS 0.012498f
C599 B.n433 VSUBS 0.012498f
C600 B.n434 VSUBS 0.012498f
C601 B.n435 VSUBS 0.012498f
C602 B.n436 VSUBS 0.012498f
C603 B.n437 VSUBS 0.012498f
C604 B.n438 VSUBS 0.012498f
C605 B.n439 VSUBS 0.012498f
C606 B.n440 VSUBS 0.012498f
C607 B.n441 VSUBS 0.012498f
C608 B.n442 VSUBS 0.012498f
C609 B.n443 VSUBS 0.012498f
C610 B.n444 VSUBS 0.012498f
C611 B.n445 VSUBS 0.012498f
C612 B.n446 VSUBS 0.012498f
C613 B.n447 VSUBS 0.012498f
C614 B.n448 VSUBS 0.012498f
C615 B.n449 VSUBS 0.012498f
C616 B.n450 VSUBS 0.012498f
C617 B.n451 VSUBS 0.012498f
C618 B.n452 VSUBS 0.012498f
C619 B.n453 VSUBS 0.012498f
C620 B.n454 VSUBS 0.012498f
C621 B.n455 VSUBS 0.012498f
C622 B.n456 VSUBS 0.012498f
C623 B.n457 VSUBS 0.012498f
C624 B.n458 VSUBS 0.012498f
C625 B.n459 VSUBS 0.012498f
C626 B.n460 VSUBS 0.012498f
C627 B.n461 VSUBS 0.012498f
C628 B.n462 VSUBS 0.012498f
C629 B.n463 VSUBS 0.012498f
C630 B.n464 VSUBS 0.012498f
C631 B.n465 VSUBS 0.012498f
C632 B.n466 VSUBS 0.012498f
C633 B.n467 VSUBS 0.012498f
C634 B.n468 VSUBS 0.012498f
C635 B.n469 VSUBS 0.012498f
C636 B.n470 VSUBS 0.012498f
C637 B.n471 VSUBS 0.012498f
C638 B.n472 VSUBS 0.012498f
C639 B.n473 VSUBS 0.012498f
C640 B.n474 VSUBS 0.012498f
C641 B.n475 VSUBS 0.012498f
C642 B.n476 VSUBS 0.012498f
C643 B.n477 VSUBS 0.012498f
C644 B.n478 VSUBS 0.012498f
C645 B.n479 VSUBS 0.012498f
C646 B.n480 VSUBS 0.012498f
C647 B.n481 VSUBS 0.012498f
C648 B.n482 VSUBS 0.012498f
C649 B.n483 VSUBS 0.012498f
C650 B.n484 VSUBS 0.012498f
C651 B.n485 VSUBS 0.012498f
C652 B.n486 VSUBS 0.012498f
C653 B.n487 VSUBS 0.012498f
C654 B.n488 VSUBS 0.012498f
C655 B.n489 VSUBS 0.012498f
C656 B.n490 VSUBS 0.012498f
C657 B.n491 VSUBS 0.012498f
C658 B.n492 VSUBS 0.012498f
C659 B.n493 VSUBS 0.012498f
C660 B.n494 VSUBS 0.012498f
C661 B.n495 VSUBS 0.012498f
C662 B.n496 VSUBS 0.012498f
C663 B.n497 VSUBS 0.012498f
C664 B.n498 VSUBS 0.012498f
C665 B.n499 VSUBS 0.012498f
C666 B.n500 VSUBS 0.012498f
C667 B.n501 VSUBS 0.012498f
C668 B.n502 VSUBS 0.012498f
C669 B.n503 VSUBS 0.012498f
C670 B.n504 VSUBS 0.012498f
C671 B.n505 VSUBS 0.012498f
C672 B.n506 VSUBS 0.012498f
C673 B.n507 VSUBS 0.012498f
C674 B.n508 VSUBS 0.012498f
C675 B.n509 VSUBS 0.012498f
C676 B.n510 VSUBS 0.012498f
C677 B.n511 VSUBS 0.012498f
C678 B.n512 VSUBS 0.012498f
C679 B.n513 VSUBS 0.012498f
C680 B.n514 VSUBS 0.012498f
C681 B.n515 VSUBS 0.012498f
C682 B.n516 VSUBS 0.012498f
C683 B.n517 VSUBS 0.012498f
C684 B.n518 VSUBS 0.012498f
C685 B.n519 VSUBS 0.012498f
C686 B.n520 VSUBS 0.012498f
C687 B.n521 VSUBS 0.012498f
C688 B.n522 VSUBS 0.012498f
C689 B.n523 VSUBS 0.012498f
C690 B.n524 VSUBS 0.012498f
C691 B.n525 VSUBS 0.012498f
C692 B.n526 VSUBS 0.012498f
C693 B.n527 VSUBS 0.012498f
C694 B.n528 VSUBS 0.012498f
C695 B.n529 VSUBS 0.012498f
C696 B.n530 VSUBS 0.012498f
C697 B.n531 VSUBS 0.012498f
C698 B.n532 VSUBS 0.012498f
C699 B.n533 VSUBS 0.012498f
C700 B.n534 VSUBS 0.012498f
C701 B.n535 VSUBS 0.012498f
C702 B.n536 VSUBS 0.012498f
C703 B.n537 VSUBS 0.012498f
C704 B.n538 VSUBS 0.012498f
C705 B.n539 VSUBS 0.012498f
C706 B.n540 VSUBS 0.012498f
C707 B.n541 VSUBS 0.012498f
C708 B.n542 VSUBS 0.012498f
C709 B.n543 VSUBS 0.012498f
C710 B.n544 VSUBS 0.012498f
C711 B.n545 VSUBS 0.012498f
C712 B.n546 VSUBS 0.012498f
C713 B.n547 VSUBS 0.012498f
C714 B.n548 VSUBS 0.012498f
C715 B.n549 VSUBS 0.012498f
C716 B.n550 VSUBS 0.012498f
C717 B.n551 VSUBS 0.012498f
C718 B.n552 VSUBS 0.012498f
C719 B.n553 VSUBS 0.012498f
C720 B.n554 VSUBS 0.012498f
C721 B.n555 VSUBS 0.012498f
C722 B.n556 VSUBS 0.012498f
C723 B.n557 VSUBS 0.012498f
C724 B.n558 VSUBS 0.012498f
C725 B.n559 VSUBS 0.012498f
C726 B.n560 VSUBS 0.012498f
C727 B.n561 VSUBS 0.012498f
C728 B.n562 VSUBS 0.012498f
C729 B.n563 VSUBS 0.012498f
C730 B.n564 VSUBS 0.012498f
C731 B.n565 VSUBS 0.012498f
C732 B.n566 VSUBS 0.012498f
C733 B.n567 VSUBS 0.012498f
C734 B.n568 VSUBS 0.012498f
C735 B.n569 VSUBS 0.012498f
C736 B.n570 VSUBS 0.012498f
C737 B.n571 VSUBS 0.012498f
C738 B.n572 VSUBS 0.012498f
C739 B.n573 VSUBS 0.012498f
C740 B.n574 VSUBS 0.012498f
C741 B.n575 VSUBS 0.012498f
C742 B.n576 VSUBS 0.012498f
C743 B.n577 VSUBS 0.012498f
C744 B.n578 VSUBS 0.012498f
C745 B.n579 VSUBS 0.012498f
C746 B.n580 VSUBS 0.012498f
C747 B.n581 VSUBS 0.012498f
C748 B.n582 VSUBS 0.012498f
C749 B.n583 VSUBS 0.012498f
C750 B.n584 VSUBS 0.012498f
C751 B.n585 VSUBS 0.012498f
C752 B.n586 VSUBS 0.012498f
C753 B.n587 VSUBS 0.012498f
C754 B.n588 VSUBS 0.012498f
C755 B.n589 VSUBS 0.012498f
C756 B.n590 VSUBS 0.012498f
C757 B.n591 VSUBS 0.012498f
C758 B.n592 VSUBS 0.012498f
C759 B.n593 VSUBS 0.012498f
C760 B.n594 VSUBS 0.012498f
C761 B.n595 VSUBS 0.012498f
C762 B.n596 VSUBS 0.012498f
C763 B.n597 VSUBS 0.012498f
C764 B.n598 VSUBS 0.012498f
C765 B.n599 VSUBS 0.012498f
C766 B.n600 VSUBS 0.012498f
C767 B.n601 VSUBS 0.012498f
C768 B.n602 VSUBS 0.012498f
C769 B.n603 VSUBS 0.012498f
C770 B.n604 VSUBS 0.012498f
C771 B.n605 VSUBS 0.012498f
C772 B.n606 VSUBS 0.012498f
C773 B.n607 VSUBS 0.012498f
C774 B.n608 VSUBS 0.012498f
C775 B.n609 VSUBS 0.012498f
C776 B.n610 VSUBS 0.012498f
C777 B.n611 VSUBS 0.012498f
C778 B.n612 VSUBS 0.012498f
C779 B.n613 VSUBS 0.012498f
C780 B.n614 VSUBS 0.012498f
C781 B.n615 VSUBS 0.012498f
C782 B.n616 VSUBS 0.012498f
C783 B.n617 VSUBS 0.012498f
C784 B.n618 VSUBS 0.012498f
C785 B.n619 VSUBS 0.012498f
C786 B.n620 VSUBS 0.012498f
C787 B.n621 VSUBS 0.012498f
C788 B.n622 VSUBS 0.026346f
C789 B.n623 VSUBS 0.027691f
C790 B.n624 VSUBS 0.027691f
C791 B.n625 VSUBS 0.012498f
C792 B.n626 VSUBS 0.012498f
C793 B.n627 VSUBS 0.012498f
C794 B.n628 VSUBS 0.012498f
C795 B.n629 VSUBS 0.012498f
C796 B.n630 VSUBS 0.012498f
C797 B.n631 VSUBS 0.012498f
C798 B.n632 VSUBS 0.012498f
C799 B.n633 VSUBS 0.012498f
C800 B.n634 VSUBS 0.012498f
C801 B.n635 VSUBS 0.012498f
C802 B.n636 VSUBS 0.012498f
C803 B.n637 VSUBS 0.012498f
C804 B.n638 VSUBS 0.012498f
C805 B.n639 VSUBS 0.012498f
C806 B.n640 VSUBS 0.012498f
C807 B.n641 VSUBS 0.012498f
C808 B.n642 VSUBS 0.012498f
C809 B.n643 VSUBS 0.012498f
C810 B.n644 VSUBS 0.012498f
C811 B.n645 VSUBS 0.012498f
C812 B.n646 VSUBS 0.012498f
C813 B.n647 VSUBS 0.012498f
C814 B.n648 VSUBS 0.012498f
C815 B.n649 VSUBS 0.012498f
C816 B.n650 VSUBS 0.012498f
C817 B.n651 VSUBS 0.012498f
C818 B.n652 VSUBS 0.012498f
C819 B.n653 VSUBS 0.008639f
C820 B.n654 VSUBS 0.012498f
C821 B.n655 VSUBS 0.012498f
C822 B.n656 VSUBS 0.010109f
C823 B.n657 VSUBS 0.012498f
C824 B.n658 VSUBS 0.012498f
C825 B.n659 VSUBS 0.012498f
C826 B.n660 VSUBS 0.012498f
C827 B.n661 VSUBS 0.012498f
C828 B.n662 VSUBS 0.012498f
C829 B.n663 VSUBS 0.012498f
C830 B.n664 VSUBS 0.012498f
C831 B.n665 VSUBS 0.012498f
C832 B.n666 VSUBS 0.012498f
C833 B.n667 VSUBS 0.012498f
C834 B.n668 VSUBS 0.010109f
C835 B.n669 VSUBS 0.028957f
C836 B.n670 VSUBS 0.008639f
C837 B.n671 VSUBS 0.012498f
C838 B.n672 VSUBS 0.012498f
C839 B.n673 VSUBS 0.012498f
C840 B.n674 VSUBS 0.012498f
C841 B.n675 VSUBS 0.012498f
C842 B.n676 VSUBS 0.012498f
C843 B.n677 VSUBS 0.012498f
C844 B.n678 VSUBS 0.012498f
C845 B.n679 VSUBS 0.012498f
C846 B.n680 VSUBS 0.012498f
C847 B.n681 VSUBS 0.012498f
C848 B.n682 VSUBS 0.012498f
C849 B.n683 VSUBS 0.012498f
C850 B.n684 VSUBS 0.012498f
C851 B.n685 VSUBS 0.012498f
C852 B.n686 VSUBS 0.012498f
C853 B.n687 VSUBS 0.012498f
C854 B.n688 VSUBS 0.012498f
C855 B.n689 VSUBS 0.012498f
C856 B.n690 VSUBS 0.012498f
C857 B.n691 VSUBS 0.012498f
C858 B.n692 VSUBS 0.012498f
C859 B.n693 VSUBS 0.012498f
C860 B.n694 VSUBS 0.012498f
C861 B.n695 VSUBS 0.012498f
C862 B.n696 VSUBS 0.012498f
C863 B.n697 VSUBS 0.012498f
C864 B.n698 VSUBS 0.012498f
C865 B.n699 VSUBS 0.012498f
C866 B.n700 VSUBS 0.027691f
C867 B.n701 VSUBS 0.026346f
C868 B.n702 VSUBS 0.026346f
C869 B.n703 VSUBS 0.012498f
C870 B.n704 VSUBS 0.012498f
C871 B.n705 VSUBS 0.012498f
C872 B.n706 VSUBS 0.012498f
C873 B.n707 VSUBS 0.012498f
C874 B.n708 VSUBS 0.012498f
C875 B.n709 VSUBS 0.012498f
C876 B.n710 VSUBS 0.012498f
C877 B.n711 VSUBS 0.012498f
C878 B.n712 VSUBS 0.012498f
C879 B.n713 VSUBS 0.012498f
C880 B.n714 VSUBS 0.012498f
C881 B.n715 VSUBS 0.012498f
C882 B.n716 VSUBS 0.012498f
C883 B.n717 VSUBS 0.012498f
C884 B.n718 VSUBS 0.012498f
C885 B.n719 VSUBS 0.012498f
C886 B.n720 VSUBS 0.012498f
C887 B.n721 VSUBS 0.012498f
C888 B.n722 VSUBS 0.012498f
C889 B.n723 VSUBS 0.012498f
C890 B.n724 VSUBS 0.012498f
C891 B.n725 VSUBS 0.012498f
C892 B.n726 VSUBS 0.012498f
C893 B.n727 VSUBS 0.012498f
C894 B.n728 VSUBS 0.012498f
C895 B.n729 VSUBS 0.012498f
C896 B.n730 VSUBS 0.012498f
C897 B.n731 VSUBS 0.012498f
C898 B.n732 VSUBS 0.012498f
C899 B.n733 VSUBS 0.012498f
C900 B.n734 VSUBS 0.012498f
C901 B.n735 VSUBS 0.012498f
C902 B.n736 VSUBS 0.012498f
C903 B.n737 VSUBS 0.012498f
C904 B.n738 VSUBS 0.012498f
C905 B.n739 VSUBS 0.012498f
C906 B.n740 VSUBS 0.012498f
C907 B.n741 VSUBS 0.012498f
C908 B.n742 VSUBS 0.012498f
C909 B.n743 VSUBS 0.012498f
C910 B.n744 VSUBS 0.012498f
C911 B.n745 VSUBS 0.012498f
C912 B.n746 VSUBS 0.012498f
C913 B.n747 VSUBS 0.012498f
C914 B.n748 VSUBS 0.012498f
C915 B.n749 VSUBS 0.012498f
C916 B.n750 VSUBS 0.012498f
C917 B.n751 VSUBS 0.012498f
C918 B.n752 VSUBS 0.012498f
C919 B.n753 VSUBS 0.012498f
C920 B.n754 VSUBS 0.012498f
C921 B.n755 VSUBS 0.012498f
C922 B.n756 VSUBS 0.012498f
C923 B.n757 VSUBS 0.012498f
C924 B.n758 VSUBS 0.012498f
C925 B.n759 VSUBS 0.012498f
C926 B.n760 VSUBS 0.012498f
C927 B.n761 VSUBS 0.012498f
C928 B.n762 VSUBS 0.012498f
C929 B.n763 VSUBS 0.012498f
C930 B.n764 VSUBS 0.012498f
C931 B.n765 VSUBS 0.012498f
C932 B.n766 VSUBS 0.012498f
C933 B.n767 VSUBS 0.012498f
C934 B.n768 VSUBS 0.012498f
C935 B.n769 VSUBS 0.012498f
C936 B.n770 VSUBS 0.012498f
C937 B.n771 VSUBS 0.012498f
C938 B.n772 VSUBS 0.012498f
C939 B.n773 VSUBS 0.012498f
C940 B.n774 VSUBS 0.012498f
C941 B.n775 VSUBS 0.012498f
C942 B.n776 VSUBS 0.012498f
C943 B.n777 VSUBS 0.012498f
C944 B.n778 VSUBS 0.012498f
C945 B.n779 VSUBS 0.012498f
C946 B.n780 VSUBS 0.012498f
C947 B.n781 VSUBS 0.012498f
C948 B.n782 VSUBS 0.012498f
C949 B.n783 VSUBS 0.012498f
C950 B.n784 VSUBS 0.012498f
C951 B.n785 VSUBS 0.012498f
C952 B.n786 VSUBS 0.012498f
C953 B.n787 VSUBS 0.012498f
C954 B.n788 VSUBS 0.012498f
C955 B.n789 VSUBS 0.012498f
C956 B.n790 VSUBS 0.012498f
C957 B.n791 VSUBS 0.012498f
C958 B.n792 VSUBS 0.012498f
C959 B.n793 VSUBS 0.012498f
C960 B.n794 VSUBS 0.012498f
C961 B.n795 VSUBS 0.012498f
C962 B.n796 VSUBS 0.012498f
C963 B.n797 VSUBS 0.012498f
C964 B.n798 VSUBS 0.012498f
C965 B.n799 VSUBS 0.012498f
C966 B.n800 VSUBS 0.012498f
C967 B.n801 VSUBS 0.012498f
C968 B.n802 VSUBS 0.012498f
C969 B.n803 VSUBS 0.012498f
C970 B.n804 VSUBS 0.012498f
C971 B.n805 VSUBS 0.012498f
C972 B.n806 VSUBS 0.012498f
C973 B.n807 VSUBS 0.012498f
C974 B.n808 VSUBS 0.012498f
C975 B.n809 VSUBS 0.012498f
C976 B.n810 VSUBS 0.012498f
C977 B.n811 VSUBS 0.01631f
C978 B.n812 VSUBS 0.017374f
C979 B.n813 VSUBS 0.03455f
C980 VTAIL.t4 VSUBS 0.139254f
C981 VTAIL.t3 VSUBS 0.139254f
C982 VTAIL.n0 VSUBS 0.754527f
C983 VTAIL.n1 VSUBS 1.14848f
C984 VTAIL.t10 VSUBS 1.05947f
C985 VTAIL.n2 VSUBS 1.31113f
C986 VTAIL.t15 VSUBS 0.139254f
C987 VTAIL.t16 VSUBS 0.139254f
C988 VTAIL.n3 VSUBS 0.754527f
C989 VTAIL.n4 VSUBS 1.37052f
C990 VTAIL.t11 VSUBS 0.139254f
C991 VTAIL.t14 VSUBS 0.139254f
C992 VTAIL.n5 VSUBS 0.754527f
C993 VTAIL.n6 VSUBS 2.73205f
C994 VTAIL.t5 VSUBS 0.139254f
C995 VTAIL.t19 VSUBS 0.139254f
C996 VTAIL.n7 VSUBS 0.754532f
C997 VTAIL.n8 VSUBS 2.73205f
C998 VTAIL.t2 VSUBS 0.139254f
C999 VTAIL.t1 VSUBS 0.139254f
C1000 VTAIL.n9 VSUBS 0.754532f
C1001 VTAIL.n10 VSUBS 1.37052f
C1002 VTAIL.t7 VSUBS 1.05947f
C1003 VTAIL.n11 VSUBS 1.31112f
C1004 VTAIL.t13 VSUBS 0.139254f
C1005 VTAIL.t17 VSUBS 0.139254f
C1006 VTAIL.n12 VSUBS 0.754532f
C1007 VTAIL.n13 VSUBS 1.23628f
C1008 VTAIL.t12 VSUBS 0.139254f
C1009 VTAIL.t18 VSUBS 0.139254f
C1010 VTAIL.n14 VSUBS 0.754532f
C1011 VTAIL.n15 VSUBS 1.37052f
C1012 VTAIL.t9 VSUBS 1.05947f
C1013 VTAIL.n16 VSUBS 2.42842f
C1014 VTAIL.t6 VSUBS 1.05947f
C1015 VTAIL.n17 VSUBS 2.42842f
C1016 VTAIL.t0 VSUBS 0.139254f
C1017 VTAIL.t8 VSUBS 0.139254f
C1018 VTAIL.n18 VSUBS 0.754527f
C1019 VTAIL.n19 VSUBS 1.07985f
C1020 VDD1.t7 VSUBS 1.2137f
C1021 VDD1.t3 VSUBS 0.140279f
C1022 VDD1.t0 VSUBS 0.140279f
C1023 VDD1.n0 VSUBS 0.871332f
C1024 VDD1.n1 VSUBS 2.03283f
C1025 VDD1.t2 VSUBS 1.21369f
C1026 VDD1.t5 VSUBS 0.140279f
C1027 VDD1.t4 VSUBS 0.140279f
C1028 VDD1.n2 VSUBS 0.871328f
C1029 VDD1.n3 VSUBS 2.02058f
C1030 VDD1.t6 VSUBS 0.140279f
C1031 VDD1.t9 VSUBS 0.140279f
C1032 VDD1.n4 VSUBS 0.900108f
C1033 VDD1.n5 VSUBS 4.70623f
C1034 VDD1.t1 VSUBS 0.140279f
C1035 VDD1.t8 VSUBS 0.140279f
C1036 VDD1.n6 VSUBS 0.871327f
C1037 VDD1.n7 VSUBS 4.59538f
C1038 VP.t8 VSUBS 1.69887f
C1039 VP.n0 VSUBS 0.797643f
C1040 VP.n1 VSUBS 0.039244f
C1041 VP.n2 VSUBS 0.04038f
C1042 VP.n3 VSUBS 0.039244f
C1043 VP.t2 VSUBS 1.69887f
C1044 VP.n4 VSUBS 0.681223f
C1045 VP.n5 VSUBS 0.039244f
C1046 VP.n6 VSUBS 0.04038f
C1047 VP.n7 VSUBS 0.039244f
C1048 VP.t3 VSUBS 1.69887f
C1049 VP.n8 VSUBS 0.644192f
C1050 VP.n9 VSUBS 0.039244f
C1051 VP.n10 VSUBS 0.04038f
C1052 VP.n11 VSUBS 0.039244f
C1053 VP.t4 VSUBS 1.69887f
C1054 VP.n12 VSUBS 0.681223f
C1055 VP.n13 VSUBS 0.039244f
C1056 VP.n14 VSUBS 0.04038f
C1057 VP.n15 VSUBS 0.039244f
C1058 VP.t7 VSUBS 1.69887f
C1059 VP.n16 VSUBS 0.797643f
C1060 VP.t9 VSUBS 1.69887f
C1061 VP.n17 VSUBS 0.797643f
C1062 VP.n18 VSUBS 0.039244f
C1063 VP.n19 VSUBS 0.04038f
C1064 VP.n20 VSUBS 0.039244f
C1065 VP.t0 VSUBS 1.69887f
C1066 VP.n21 VSUBS 0.681223f
C1067 VP.n22 VSUBS 0.039244f
C1068 VP.n23 VSUBS 0.04038f
C1069 VP.n24 VSUBS 0.039244f
C1070 VP.t6 VSUBS 1.69887f
C1071 VP.n25 VSUBS 0.644192f
C1072 VP.n26 VSUBS 0.039244f
C1073 VP.n27 VSUBS 0.04038f
C1074 VP.n28 VSUBS 0.039244f
C1075 VP.t1 VSUBS 1.69887f
C1076 VP.n29 VSUBS 0.79953f
C1077 VP.t5 VSUBS 2.16469f
C1078 VP.n30 VSUBS 0.755778f
C1079 VP.n31 VSUBS 0.479314f
C1080 VP.n32 VSUBS 0.073141f
C1081 VP.n33 VSUBS 0.073141f
C1082 VP.n34 VSUBS 0.070049f
C1083 VP.n35 VSUBS 0.039244f
C1084 VP.n36 VSUBS 0.039244f
C1085 VP.n37 VSUBS 0.039244f
C1086 VP.n38 VSUBS 0.077298f
C1087 VP.n39 VSUBS 0.073141f
C1088 VP.n40 VSUBS 0.055086f
C1089 VP.n41 VSUBS 0.039244f
C1090 VP.n42 VSUBS 0.039244f
C1091 VP.n43 VSUBS 0.055086f
C1092 VP.n44 VSUBS 0.073141f
C1093 VP.n45 VSUBS 0.077298f
C1094 VP.n46 VSUBS 0.039244f
C1095 VP.n47 VSUBS 0.039244f
C1096 VP.n48 VSUBS 0.039244f
C1097 VP.n49 VSUBS 0.070049f
C1098 VP.n50 VSUBS 0.073141f
C1099 VP.n51 VSUBS 0.073141f
C1100 VP.n52 VSUBS 0.039244f
C1101 VP.n53 VSUBS 0.039244f
C1102 VP.n54 VSUBS 0.039244f
C1103 VP.n55 VSUBS 0.073141f
C1104 VP.n56 VSUBS 0.073141f
C1105 VP.n57 VSUBS 0.070049f
C1106 VP.n58 VSUBS 0.039244f
C1107 VP.n59 VSUBS 0.039244f
C1108 VP.n60 VSUBS 0.039244f
C1109 VP.n61 VSUBS 0.077298f
C1110 VP.n62 VSUBS 0.073141f
C1111 VP.n63 VSUBS 0.055086f
C1112 VP.n64 VSUBS 0.063339f
C1113 VP.n65 VSUBS 2.38373f
C1114 VP.n66 VSUBS 2.41072f
C1115 VP.n67 VSUBS 0.063339f
C1116 VP.n68 VSUBS 0.055086f
C1117 VP.n69 VSUBS 0.073141f
C1118 VP.n70 VSUBS 0.077298f
C1119 VP.n71 VSUBS 0.039244f
C1120 VP.n72 VSUBS 0.039244f
C1121 VP.n73 VSUBS 0.039244f
C1122 VP.n74 VSUBS 0.070049f
C1123 VP.n75 VSUBS 0.073141f
C1124 VP.n76 VSUBS 0.073141f
C1125 VP.n77 VSUBS 0.039244f
C1126 VP.n78 VSUBS 0.039244f
C1127 VP.n79 VSUBS 0.039244f
C1128 VP.n80 VSUBS 0.073141f
C1129 VP.n81 VSUBS 0.073141f
C1130 VP.n82 VSUBS 0.070049f
C1131 VP.n83 VSUBS 0.039244f
C1132 VP.n84 VSUBS 0.039244f
C1133 VP.n85 VSUBS 0.039244f
C1134 VP.n86 VSUBS 0.077298f
C1135 VP.n87 VSUBS 0.073141f
C1136 VP.n88 VSUBS 0.055086f
C1137 VP.n89 VSUBS 0.039244f
C1138 VP.n90 VSUBS 0.039244f
C1139 VP.n91 VSUBS 0.055086f
C1140 VP.n92 VSUBS 0.073141f
C1141 VP.n93 VSUBS 0.077298f
C1142 VP.n94 VSUBS 0.039244f
C1143 VP.n95 VSUBS 0.039244f
C1144 VP.n96 VSUBS 0.039244f
C1145 VP.n97 VSUBS 0.070049f
C1146 VP.n98 VSUBS 0.073141f
C1147 VP.n99 VSUBS 0.073141f
C1148 VP.n100 VSUBS 0.039244f
C1149 VP.n101 VSUBS 0.039244f
C1150 VP.n102 VSUBS 0.039244f
C1151 VP.n103 VSUBS 0.073141f
C1152 VP.n104 VSUBS 0.073141f
C1153 VP.n105 VSUBS 0.070049f
C1154 VP.n106 VSUBS 0.039244f
C1155 VP.n107 VSUBS 0.039244f
C1156 VP.n108 VSUBS 0.039244f
C1157 VP.n109 VSUBS 0.077298f
C1158 VP.n110 VSUBS 0.073141f
C1159 VP.n111 VSUBS 0.055086f
C1160 VP.n112 VSUBS 0.063339f
C1161 VP.n113 VSUBS 0.100735f
.ends

