* NGSPICE file created from diff_pair_sample_0298.ext - technology: sky130A

.subckt diff_pair_sample_0298 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=3.2175 ps=17.28 w=8.25 l=0.97
X1 VDD1.t0 VP.t1 VTAIL.t2 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=3.2175 ps=17.28 w=8.25 l=0.97
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=3.2175 ps=17.28 w=8.25 l=0.97
X3 B.t11 B.t9 B.t10 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=0 ps=0 w=8.25 l=0.97
X4 B.t8 B.t6 B.t7 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=0 ps=0 w=8.25 l=0.97
X5 B.t5 B.t3 B.t4 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=0 ps=0 w=8.25 l=0.97
X6 B.t2 B.t0 B.t1 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=0 ps=0 w=8.25 l=0.97
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1490_n2622# sky130_fd_pr__pfet_01v8 ad=3.2175 pd=17.28 as=3.2175 ps=17.28 w=8.25 l=0.97
R0 VP.n0 VP.t1 444.529
R1 VP.n0 VP.t0 407.022
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 70.2914
R4 VTAIL.n3 VTAIL.t3 70.2913
R5 VTAIL.n0 VTAIL.t1 70.2913
R6 VTAIL.n2 VTAIL.t2 70.2913
R7 VTAIL.n1 VTAIL.n0 21.7376
R8 VTAIL.n3 VTAIL.n2 20.6169
R9 VTAIL.n2 VTAIL.n1 1.03067
R10 VTAIL VTAIL.n0 0.80869
R11 VTAIL VTAIL.n3 0.222483
R12 VDD1 VDD1.t1 120.805
R13 VDD1 VDD1.t0 87.3085
R14 VN VN.t1 444.909
R15 VN VN.t0 407.072
R16 VDD2.n0 VDD2.t1 120.001
R17 VDD2.n0 VDD2.t0 86.9701
R18 VDD2 VDD2.n0 0.338862
R19 B.n240 B.n65 585
R20 B.n239 B.n238 585
R21 B.n237 B.n66 585
R22 B.n236 B.n235 585
R23 B.n234 B.n67 585
R24 B.n233 B.n232 585
R25 B.n231 B.n68 585
R26 B.n230 B.n229 585
R27 B.n228 B.n69 585
R28 B.n227 B.n226 585
R29 B.n225 B.n70 585
R30 B.n224 B.n223 585
R31 B.n222 B.n71 585
R32 B.n221 B.n220 585
R33 B.n219 B.n72 585
R34 B.n218 B.n217 585
R35 B.n216 B.n73 585
R36 B.n215 B.n214 585
R37 B.n213 B.n74 585
R38 B.n212 B.n211 585
R39 B.n210 B.n75 585
R40 B.n209 B.n208 585
R41 B.n207 B.n76 585
R42 B.n206 B.n205 585
R43 B.n204 B.n77 585
R44 B.n203 B.n202 585
R45 B.n201 B.n78 585
R46 B.n200 B.n199 585
R47 B.n198 B.n79 585
R48 B.n197 B.n196 585
R49 B.n195 B.n80 585
R50 B.n194 B.n193 585
R51 B.n189 B.n81 585
R52 B.n188 B.n187 585
R53 B.n186 B.n82 585
R54 B.n185 B.n184 585
R55 B.n183 B.n83 585
R56 B.n182 B.n181 585
R57 B.n180 B.n84 585
R58 B.n179 B.n178 585
R59 B.n176 B.n85 585
R60 B.n175 B.n174 585
R61 B.n173 B.n88 585
R62 B.n172 B.n171 585
R63 B.n170 B.n89 585
R64 B.n169 B.n168 585
R65 B.n167 B.n90 585
R66 B.n166 B.n165 585
R67 B.n164 B.n91 585
R68 B.n163 B.n162 585
R69 B.n161 B.n92 585
R70 B.n160 B.n159 585
R71 B.n158 B.n93 585
R72 B.n157 B.n156 585
R73 B.n155 B.n94 585
R74 B.n154 B.n153 585
R75 B.n152 B.n95 585
R76 B.n151 B.n150 585
R77 B.n149 B.n96 585
R78 B.n148 B.n147 585
R79 B.n146 B.n97 585
R80 B.n145 B.n144 585
R81 B.n143 B.n98 585
R82 B.n142 B.n141 585
R83 B.n140 B.n99 585
R84 B.n139 B.n138 585
R85 B.n137 B.n100 585
R86 B.n136 B.n135 585
R87 B.n134 B.n101 585
R88 B.n133 B.n132 585
R89 B.n131 B.n102 585
R90 B.n242 B.n241 585
R91 B.n243 B.n64 585
R92 B.n245 B.n244 585
R93 B.n246 B.n63 585
R94 B.n248 B.n247 585
R95 B.n249 B.n62 585
R96 B.n251 B.n250 585
R97 B.n252 B.n61 585
R98 B.n254 B.n253 585
R99 B.n255 B.n60 585
R100 B.n257 B.n256 585
R101 B.n258 B.n59 585
R102 B.n260 B.n259 585
R103 B.n261 B.n58 585
R104 B.n263 B.n262 585
R105 B.n264 B.n57 585
R106 B.n266 B.n265 585
R107 B.n267 B.n56 585
R108 B.n269 B.n268 585
R109 B.n270 B.n55 585
R110 B.n272 B.n271 585
R111 B.n273 B.n54 585
R112 B.n275 B.n274 585
R113 B.n276 B.n53 585
R114 B.n278 B.n277 585
R115 B.n279 B.n52 585
R116 B.n281 B.n280 585
R117 B.n282 B.n51 585
R118 B.n284 B.n283 585
R119 B.n285 B.n50 585
R120 B.n287 B.n286 585
R121 B.n288 B.n49 585
R122 B.n397 B.n396 585
R123 B.n395 B.n10 585
R124 B.n394 B.n393 585
R125 B.n392 B.n11 585
R126 B.n391 B.n390 585
R127 B.n389 B.n12 585
R128 B.n388 B.n387 585
R129 B.n386 B.n13 585
R130 B.n385 B.n384 585
R131 B.n383 B.n14 585
R132 B.n382 B.n381 585
R133 B.n380 B.n15 585
R134 B.n379 B.n378 585
R135 B.n377 B.n16 585
R136 B.n376 B.n375 585
R137 B.n374 B.n17 585
R138 B.n373 B.n372 585
R139 B.n371 B.n18 585
R140 B.n370 B.n369 585
R141 B.n368 B.n19 585
R142 B.n367 B.n366 585
R143 B.n365 B.n20 585
R144 B.n364 B.n363 585
R145 B.n362 B.n21 585
R146 B.n361 B.n360 585
R147 B.n359 B.n22 585
R148 B.n358 B.n357 585
R149 B.n356 B.n23 585
R150 B.n355 B.n354 585
R151 B.n353 B.n24 585
R152 B.n352 B.n351 585
R153 B.n349 B.n25 585
R154 B.n348 B.n347 585
R155 B.n346 B.n28 585
R156 B.n345 B.n344 585
R157 B.n343 B.n29 585
R158 B.n342 B.n341 585
R159 B.n340 B.n30 585
R160 B.n339 B.n338 585
R161 B.n337 B.n31 585
R162 B.n335 B.n334 585
R163 B.n333 B.n34 585
R164 B.n332 B.n331 585
R165 B.n330 B.n35 585
R166 B.n329 B.n328 585
R167 B.n327 B.n36 585
R168 B.n326 B.n325 585
R169 B.n324 B.n37 585
R170 B.n323 B.n322 585
R171 B.n321 B.n38 585
R172 B.n320 B.n319 585
R173 B.n318 B.n39 585
R174 B.n317 B.n316 585
R175 B.n315 B.n40 585
R176 B.n314 B.n313 585
R177 B.n312 B.n41 585
R178 B.n311 B.n310 585
R179 B.n309 B.n42 585
R180 B.n308 B.n307 585
R181 B.n306 B.n43 585
R182 B.n305 B.n304 585
R183 B.n303 B.n44 585
R184 B.n302 B.n301 585
R185 B.n300 B.n45 585
R186 B.n299 B.n298 585
R187 B.n297 B.n46 585
R188 B.n296 B.n295 585
R189 B.n294 B.n47 585
R190 B.n293 B.n292 585
R191 B.n291 B.n48 585
R192 B.n290 B.n289 585
R193 B.n398 B.n9 585
R194 B.n400 B.n399 585
R195 B.n401 B.n8 585
R196 B.n403 B.n402 585
R197 B.n404 B.n7 585
R198 B.n406 B.n405 585
R199 B.n407 B.n6 585
R200 B.n409 B.n408 585
R201 B.n410 B.n5 585
R202 B.n412 B.n411 585
R203 B.n413 B.n4 585
R204 B.n415 B.n414 585
R205 B.n416 B.n3 585
R206 B.n418 B.n417 585
R207 B.n419 B.n0 585
R208 B.n2 B.n1 585
R209 B.n110 B.n109 585
R210 B.n112 B.n111 585
R211 B.n113 B.n108 585
R212 B.n115 B.n114 585
R213 B.n116 B.n107 585
R214 B.n118 B.n117 585
R215 B.n119 B.n106 585
R216 B.n121 B.n120 585
R217 B.n122 B.n105 585
R218 B.n124 B.n123 585
R219 B.n125 B.n104 585
R220 B.n127 B.n126 585
R221 B.n128 B.n103 585
R222 B.n130 B.n129 585
R223 B.n131 B.n130 530.939
R224 B.n242 B.n65 530.939
R225 B.n290 B.n49 530.939
R226 B.n396 B.n9 530.939
R227 B.n86 B.t3 407.693
R228 B.n190 B.t0 407.693
R229 B.n32 B.t6 407.693
R230 B.n26 B.t9 407.693
R231 B.n421 B.n420 256.663
R232 B.n420 B.n419 235.042
R233 B.n420 B.n2 235.042
R234 B.n132 B.n131 163.367
R235 B.n132 B.n101 163.367
R236 B.n136 B.n101 163.367
R237 B.n137 B.n136 163.367
R238 B.n138 B.n137 163.367
R239 B.n138 B.n99 163.367
R240 B.n142 B.n99 163.367
R241 B.n143 B.n142 163.367
R242 B.n144 B.n143 163.367
R243 B.n144 B.n97 163.367
R244 B.n148 B.n97 163.367
R245 B.n149 B.n148 163.367
R246 B.n150 B.n149 163.367
R247 B.n150 B.n95 163.367
R248 B.n154 B.n95 163.367
R249 B.n155 B.n154 163.367
R250 B.n156 B.n155 163.367
R251 B.n156 B.n93 163.367
R252 B.n160 B.n93 163.367
R253 B.n161 B.n160 163.367
R254 B.n162 B.n161 163.367
R255 B.n162 B.n91 163.367
R256 B.n166 B.n91 163.367
R257 B.n167 B.n166 163.367
R258 B.n168 B.n167 163.367
R259 B.n168 B.n89 163.367
R260 B.n172 B.n89 163.367
R261 B.n173 B.n172 163.367
R262 B.n174 B.n173 163.367
R263 B.n174 B.n85 163.367
R264 B.n179 B.n85 163.367
R265 B.n180 B.n179 163.367
R266 B.n181 B.n180 163.367
R267 B.n181 B.n83 163.367
R268 B.n185 B.n83 163.367
R269 B.n186 B.n185 163.367
R270 B.n187 B.n186 163.367
R271 B.n187 B.n81 163.367
R272 B.n194 B.n81 163.367
R273 B.n195 B.n194 163.367
R274 B.n196 B.n195 163.367
R275 B.n196 B.n79 163.367
R276 B.n200 B.n79 163.367
R277 B.n201 B.n200 163.367
R278 B.n202 B.n201 163.367
R279 B.n202 B.n77 163.367
R280 B.n206 B.n77 163.367
R281 B.n207 B.n206 163.367
R282 B.n208 B.n207 163.367
R283 B.n208 B.n75 163.367
R284 B.n212 B.n75 163.367
R285 B.n213 B.n212 163.367
R286 B.n214 B.n213 163.367
R287 B.n214 B.n73 163.367
R288 B.n218 B.n73 163.367
R289 B.n219 B.n218 163.367
R290 B.n220 B.n219 163.367
R291 B.n220 B.n71 163.367
R292 B.n224 B.n71 163.367
R293 B.n225 B.n224 163.367
R294 B.n226 B.n225 163.367
R295 B.n226 B.n69 163.367
R296 B.n230 B.n69 163.367
R297 B.n231 B.n230 163.367
R298 B.n232 B.n231 163.367
R299 B.n232 B.n67 163.367
R300 B.n236 B.n67 163.367
R301 B.n237 B.n236 163.367
R302 B.n238 B.n237 163.367
R303 B.n238 B.n65 163.367
R304 B.n286 B.n49 163.367
R305 B.n286 B.n285 163.367
R306 B.n285 B.n284 163.367
R307 B.n284 B.n51 163.367
R308 B.n280 B.n51 163.367
R309 B.n280 B.n279 163.367
R310 B.n279 B.n278 163.367
R311 B.n278 B.n53 163.367
R312 B.n274 B.n53 163.367
R313 B.n274 B.n273 163.367
R314 B.n273 B.n272 163.367
R315 B.n272 B.n55 163.367
R316 B.n268 B.n55 163.367
R317 B.n268 B.n267 163.367
R318 B.n267 B.n266 163.367
R319 B.n266 B.n57 163.367
R320 B.n262 B.n57 163.367
R321 B.n262 B.n261 163.367
R322 B.n261 B.n260 163.367
R323 B.n260 B.n59 163.367
R324 B.n256 B.n59 163.367
R325 B.n256 B.n255 163.367
R326 B.n255 B.n254 163.367
R327 B.n254 B.n61 163.367
R328 B.n250 B.n61 163.367
R329 B.n250 B.n249 163.367
R330 B.n249 B.n248 163.367
R331 B.n248 B.n63 163.367
R332 B.n244 B.n63 163.367
R333 B.n244 B.n243 163.367
R334 B.n243 B.n242 163.367
R335 B.n396 B.n395 163.367
R336 B.n395 B.n394 163.367
R337 B.n394 B.n11 163.367
R338 B.n390 B.n11 163.367
R339 B.n390 B.n389 163.367
R340 B.n389 B.n388 163.367
R341 B.n388 B.n13 163.367
R342 B.n384 B.n13 163.367
R343 B.n384 B.n383 163.367
R344 B.n383 B.n382 163.367
R345 B.n382 B.n15 163.367
R346 B.n378 B.n15 163.367
R347 B.n378 B.n377 163.367
R348 B.n377 B.n376 163.367
R349 B.n376 B.n17 163.367
R350 B.n372 B.n17 163.367
R351 B.n372 B.n371 163.367
R352 B.n371 B.n370 163.367
R353 B.n370 B.n19 163.367
R354 B.n366 B.n19 163.367
R355 B.n366 B.n365 163.367
R356 B.n365 B.n364 163.367
R357 B.n364 B.n21 163.367
R358 B.n360 B.n21 163.367
R359 B.n360 B.n359 163.367
R360 B.n359 B.n358 163.367
R361 B.n358 B.n23 163.367
R362 B.n354 B.n23 163.367
R363 B.n354 B.n353 163.367
R364 B.n353 B.n352 163.367
R365 B.n352 B.n25 163.367
R366 B.n347 B.n25 163.367
R367 B.n347 B.n346 163.367
R368 B.n346 B.n345 163.367
R369 B.n345 B.n29 163.367
R370 B.n341 B.n29 163.367
R371 B.n341 B.n340 163.367
R372 B.n340 B.n339 163.367
R373 B.n339 B.n31 163.367
R374 B.n334 B.n31 163.367
R375 B.n334 B.n333 163.367
R376 B.n333 B.n332 163.367
R377 B.n332 B.n35 163.367
R378 B.n328 B.n35 163.367
R379 B.n328 B.n327 163.367
R380 B.n327 B.n326 163.367
R381 B.n326 B.n37 163.367
R382 B.n322 B.n37 163.367
R383 B.n322 B.n321 163.367
R384 B.n321 B.n320 163.367
R385 B.n320 B.n39 163.367
R386 B.n316 B.n39 163.367
R387 B.n316 B.n315 163.367
R388 B.n315 B.n314 163.367
R389 B.n314 B.n41 163.367
R390 B.n310 B.n41 163.367
R391 B.n310 B.n309 163.367
R392 B.n309 B.n308 163.367
R393 B.n308 B.n43 163.367
R394 B.n304 B.n43 163.367
R395 B.n304 B.n303 163.367
R396 B.n303 B.n302 163.367
R397 B.n302 B.n45 163.367
R398 B.n298 B.n45 163.367
R399 B.n298 B.n297 163.367
R400 B.n297 B.n296 163.367
R401 B.n296 B.n47 163.367
R402 B.n292 B.n47 163.367
R403 B.n292 B.n291 163.367
R404 B.n291 B.n290 163.367
R405 B.n400 B.n9 163.367
R406 B.n401 B.n400 163.367
R407 B.n402 B.n401 163.367
R408 B.n402 B.n7 163.367
R409 B.n406 B.n7 163.367
R410 B.n407 B.n406 163.367
R411 B.n408 B.n407 163.367
R412 B.n408 B.n5 163.367
R413 B.n412 B.n5 163.367
R414 B.n413 B.n412 163.367
R415 B.n414 B.n413 163.367
R416 B.n414 B.n3 163.367
R417 B.n418 B.n3 163.367
R418 B.n419 B.n418 163.367
R419 B.n109 B.n2 163.367
R420 B.n112 B.n109 163.367
R421 B.n113 B.n112 163.367
R422 B.n114 B.n113 163.367
R423 B.n114 B.n107 163.367
R424 B.n118 B.n107 163.367
R425 B.n119 B.n118 163.367
R426 B.n120 B.n119 163.367
R427 B.n120 B.n105 163.367
R428 B.n124 B.n105 163.367
R429 B.n125 B.n124 163.367
R430 B.n126 B.n125 163.367
R431 B.n126 B.n103 163.367
R432 B.n130 B.n103 163.367
R433 B.n190 B.t1 135.459
R434 B.n32 B.t8 135.459
R435 B.n86 B.t4 135.451
R436 B.n26 B.t11 135.451
R437 B.n191 B.t2 110.248
R438 B.n33 B.t7 110.248
R439 B.n87 B.t5 110.239
R440 B.n27 B.t10 110.239
R441 B.n177 B.n87 59.5399
R442 B.n192 B.n191 59.5399
R443 B.n336 B.n33 59.5399
R444 B.n350 B.n27 59.5399
R445 B.n398 B.n397 34.4981
R446 B.n289 B.n288 34.4981
R447 B.n241 B.n240 34.4981
R448 B.n129 B.n102 34.4981
R449 B.n87 B.n86 25.2126
R450 B.n191 B.n190 25.2126
R451 B.n33 B.n32 25.2126
R452 B.n27 B.n26 25.2126
R453 B B.n421 18.0485
R454 B.n399 B.n398 10.6151
R455 B.n399 B.n8 10.6151
R456 B.n403 B.n8 10.6151
R457 B.n404 B.n403 10.6151
R458 B.n405 B.n404 10.6151
R459 B.n405 B.n6 10.6151
R460 B.n409 B.n6 10.6151
R461 B.n410 B.n409 10.6151
R462 B.n411 B.n410 10.6151
R463 B.n411 B.n4 10.6151
R464 B.n415 B.n4 10.6151
R465 B.n416 B.n415 10.6151
R466 B.n417 B.n416 10.6151
R467 B.n417 B.n0 10.6151
R468 B.n397 B.n10 10.6151
R469 B.n393 B.n10 10.6151
R470 B.n393 B.n392 10.6151
R471 B.n392 B.n391 10.6151
R472 B.n391 B.n12 10.6151
R473 B.n387 B.n12 10.6151
R474 B.n387 B.n386 10.6151
R475 B.n386 B.n385 10.6151
R476 B.n385 B.n14 10.6151
R477 B.n381 B.n14 10.6151
R478 B.n381 B.n380 10.6151
R479 B.n380 B.n379 10.6151
R480 B.n379 B.n16 10.6151
R481 B.n375 B.n16 10.6151
R482 B.n375 B.n374 10.6151
R483 B.n374 B.n373 10.6151
R484 B.n373 B.n18 10.6151
R485 B.n369 B.n18 10.6151
R486 B.n369 B.n368 10.6151
R487 B.n368 B.n367 10.6151
R488 B.n367 B.n20 10.6151
R489 B.n363 B.n20 10.6151
R490 B.n363 B.n362 10.6151
R491 B.n362 B.n361 10.6151
R492 B.n361 B.n22 10.6151
R493 B.n357 B.n22 10.6151
R494 B.n357 B.n356 10.6151
R495 B.n356 B.n355 10.6151
R496 B.n355 B.n24 10.6151
R497 B.n351 B.n24 10.6151
R498 B.n349 B.n348 10.6151
R499 B.n348 B.n28 10.6151
R500 B.n344 B.n28 10.6151
R501 B.n344 B.n343 10.6151
R502 B.n343 B.n342 10.6151
R503 B.n342 B.n30 10.6151
R504 B.n338 B.n30 10.6151
R505 B.n338 B.n337 10.6151
R506 B.n335 B.n34 10.6151
R507 B.n331 B.n34 10.6151
R508 B.n331 B.n330 10.6151
R509 B.n330 B.n329 10.6151
R510 B.n329 B.n36 10.6151
R511 B.n325 B.n36 10.6151
R512 B.n325 B.n324 10.6151
R513 B.n324 B.n323 10.6151
R514 B.n323 B.n38 10.6151
R515 B.n319 B.n38 10.6151
R516 B.n319 B.n318 10.6151
R517 B.n318 B.n317 10.6151
R518 B.n317 B.n40 10.6151
R519 B.n313 B.n40 10.6151
R520 B.n313 B.n312 10.6151
R521 B.n312 B.n311 10.6151
R522 B.n311 B.n42 10.6151
R523 B.n307 B.n42 10.6151
R524 B.n307 B.n306 10.6151
R525 B.n306 B.n305 10.6151
R526 B.n305 B.n44 10.6151
R527 B.n301 B.n44 10.6151
R528 B.n301 B.n300 10.6151
R529 B.n300 B.n299 10.6151
R530 B.n299 B.n46 10.6151
R531 B.n295 B.n46 10.6151
R532 B.n295 B.n294 10.6151
R533 B.n294 B.n293 10.6151
R534 B.n293 B.n48 10.6151
R535 B.n289 B.n48 10.6151
R536 B.n288 B.n287 10.6151
R537 B.n287 B.n50 10.6151
R538 B.n283 B.n50 10.6151
R539 B.n283 B.n282 10.6151
R540 B.n282 B.n281 10.6151
R541 B.n281 B.n52 10.6151
R542 B.n277 B.n52 10.6151
R543 B.n277 B.n276 10.6151
R544 B.n276 B.n275 10.6151
R545 B.n275 B.n54 10.6151
R546 B.n271 B.n54 10.6151
R547 B.n271 B.n270 10.6151
R548 B.n270 B.n269 10.6151
R549 B.n269 B.n56 10.6151
R550 B.n265 B.n56 10.6151
R551 B.n265 B.n264 10.6151
R552 B.n264 B.n263 10.6151
R553 B.n263 B.n58 10.6151
R554 B.n259 B.n58 10.6151
R555 B.n259 B.n258 10.6151
R556 B.n258 B.n257 10.6151
R557 B.n257 B.n60 10.6151
R558 B.n253 B.n60 10.6151
R559 B.n253 B.n252 10.6151
R560 B.n252 B.n251 10.6151
R561 B.n251 B.n62 10.6151
R562 B.n247 B.n62 10.6151
R563 B.n247 B.n246 10.6151
R564 B.n246 B.n245 10.6151
R565 B.n245 B.n64 10.6151
R566 B.n241 B.n64 10.6151
R567 B.n110 B.n1 10.6151
R568 B.n111 B.n110 10.6151
R569 B.n111 B.n108 10.6151
R570 B.n115 B.n108 10.6151
R571 B.n116 B.n115 10.6151
R572 B.n117 B.n116 10.6151
R573 B.n117 B.n106 10.6151
R574 B.n121 B.n106 10.6151
R575 B.n122 B.n121 10.6151
R576 B.n123 B.n122 10.6151
R577 B.n123 B.n104 10.6151
R578 B.n127 B.n104 10.6151
R579 B.n128 B.n127 10.6151
R580 B.n129 B.n128 10.6151
R581 B.n133 B.n102 10.6151
R582 B.n134 B.n133 10.6151
R583 B.n135 B.n134 10.6151
R584 B.n135 B.n100 10.6151
R585 B.n139 B.n100 10.6151
R586 B.n140 B.n139 10.6151
R587 B.n141 B.n140 10.6151
R588 B.n141 B.n98 10.6151
R589 B.n145 B.n98 10.6151
R590 B.n146 B.n145 10.6151
R591 B.n147 B.n146 10.6151
R592 B.n147 B.n96 10.6151
R593 B.n151 B.n96 10.6151
R594 B.n152 B.n151 10.6151
R595 B.n153 B.n152 10.6151
R596 B.n153 B.n94 10.6151
R597 B.n157 B.n94 10.6151
R598 B.n158 B.n157 10.6151
R599 B.n159 B.n158 10.6151
R600 B.n159 B.n92 10.6151
R601 B.n163 B.n92 10.6151
R602 B.n164 B.n163 10.6151
R603 B.n165 B.n164 10.6151
R604 B.n165 B.n90 10.6151
R605 B.n169 B.n90 10.6151
R606 B.n170 B.n169 10.6151
R607 B.n171 B.n170 10.6151
R608 B.n171 B.n88 10.6151
R609 B.n175 B.n88 10.6151
R610 B.n176 B.n175 10.6151
R611 B.n178 B.n84 10.6151
R612 B.n182 B.n84 10.6151
R613 B.n183 B.n182 10.6151
R614 B.n184 B.n183 10.6151
R615 B.n184 B.n82 10.6151
R616 B.n188 B.n82 10.6151
R617 B.n189 B.n188 10.6151
R618 B.n193 B.n189 10.6151
R619 B.n197 B.n80 10.6151
R620 B.n198 B.n197 10.6151
R621 B.n199 B.n198 10.6151
R622 B.n199 B.n78 10.6151
R623 B.n203 B.n78 10.6151
R624 B.n204 B.n203 10.6151
R625 B.n205 B.n204 10.6151
R626 B.n205 B.n76 10.6151
R627 B.n209 B.n76 10.6151
R628 B.n210 B.n209 10.6151
R629 B.n211 B.n210 10.6151
R630 B.n211 B.n74 10.6151
R631 B.n215 B.n74 10.6151
R632 B.n216 B.n215 10.6151
R633 B.n217 B.n216 10.6151
R634 B.n217 B.n72 10.6151
R635 B.n221 B.n72 10.6151
R636 B.n222 B.n221 10.6151
R637 B.n223 B.n222 10.6151
R638 B.n223 B.n70 10.6151
R639 B.n227 B.n70 10.6151
R640 B.n228 B.n227 10.6151
R641 B.n229 B.n228 10.6151
R642 B.n229 B.n68 10.6151
R643 B.n233 B.n68 10.6151
R644 B.n234 B.n233 10.6151
R645 B.n235 B.n234 10.6151
R646 B.n235 B.n66 10.6151
R647 B.n239 B.n66 10.6151
R648 B.n240 B.n239 10.6151
R649 B.n421 B.n0 8.11757
R650 B.n421 B.n1 8.11757
R651 B.n350 B.n349 7.18099
R652 B.n337 B.n336 7.18099
R653 B.n178 B.n177 7.18099
R654 B.n193 B.n192 7.18099
R655 B.n351 B.n350 3.43465
R656 B.n336 B.n335 3.43465
R657 B.n177 B.n176 3.43465
R658 B.n192 B.n80 3.43465
C0 VDD2 VP 0.265709f
C1 VDD1 VP 1.71035f
C2 VTAIL VN 1.29312f
C3 VP B 1.02957f
C4 VTAIL w_n1490_n2622# 2.27288f
C5 VDD2 VDD1 0.488111f
C6 VP VN 3.98924f
C7 VDD2 B 1.20151f
C8 VDD1 B 1.18508f
C9 VP w_n1490_n2622# 2.02713f
C10 VDD2 VN 1.59614f
C11 VDD1 VN 0.148712f
C12 VDD2 w_n1490_n2622# 1.33509f
C13 VTAIL VP 1.30752f
C14 B VN 0.729851f
C15 VDD1 w_n1490_n2622# 1.32772f
C16 B w_n1490_n2622# 6.00082f
C17 VDD2 VTAIL 4.11412f
C18 VDD1 VTAIL 4.0757f
C19 VN w_n1490_n2622# 1.84084f
C20 VTAIL B 2.16525f
C21 VDD2 VSUBS 0.625732f
C22 VDD1 VSUBS 2.739871f
C23 VTAIL VSUBS 0.656115f
C24 VN VSUBS 3.92855f
C25 VP VSUBS 1.044368f
C26 B VSUBS 2.377986f
C27 w_n1490_n2622# VSUBS 48.436897f
C28 B.n0 VSUBS 0.006934f
C29 B.n1 VSUBS 0.006934f
C30 B.n2 VSUBS 0.010256f
C31 B.n3 VSUBS 0.007859f
C32 B.n4 VSUBS 0.007859f
C33 B.n5 VSUBS 0.007859f
C34 B.n6 VSUBS 0.007859f
C35 B.n7 VSUBS 0.007859f
C36 B.n8 VSUBS 0.007859f
C37 B.n9 VSUBS 0.018416f
C38 B.n10 VSUBS 0.007859f
C39 B.n11 VSUBS 0.007859f
C40 B.n12 VSUBS 0.007859f
C41 B.n13 VSUBS 0.007859f
C42 B.n14 VSUBS 0.007859f
C43 B.n15 VSUBS 0.007859f
C44 B.n16 VSUBS 0.007859f
C45 B.n17 VSUBS 0.007859f
C46 B.n18 VSUBS 0.007859f
C47 B.n19 VSUBS 0.007859f
C48 B.n20 VSUBS 0.007859f
C49 B.n21 VSUBS 0.007859f
C50 B.n22 VSUBS 0.007859f
C51 B.n23 VSUBS 0.007859f
C52 B.n24 VSUBS 0.007859f
C53 B.n25 VSUBS 0.007859f
C54 B.t10 VSUBS 0.287266f
C55 B.t11 VSUBS 0.298691f
C56 B.t9 VSUBS 0.389785f
C57 B.n26 VSUBS 0.129557f
C58 B.n27 VSUBS 0.072588f
C59 B.n28 VSUBS 0.007859f
C60 B.n29 VSUBS 0.007859f
C61 B.n30 VSUBS 0.007859f
C62 B.n31 VSUBS 0.007859f
C63 B.t7 VSUBS 0.287263f
C64 B.t8 VSUBS 0.298688f
C65 B.t6 VSUBS 0.389785f
C66 B.n32 VSUBS 0.129559f
C67 B.n33 VSUBS 0.072591f
C68 B.n34 VSUBS 0.007859f
C69 B.n35 VSUBS 0.007859f
C70 B.n36 VSUBS 0.007859f
C71 B.n37 VSUBS 0.007859f
C72 B.n38 VSUBS 0.007859f
C73 B.n39 VSUBS 0.007859f
C74 B.n40 VSUBS 0.007859f
C75 B.n41 VSUBS 0.007859f
C76 B.n42 VSUBS 0.007859f
C77 B.n43 VSUBS 0.007859f
C78 B.n44 VSUBS 0.007859f
C79 B.n45 VSUBS 0.007859f
C80 B.n46 VSUBS 0.007859f
C81 B.n47 VSUBS 0.007859f
C82 B.n48 VSUBS 0.007859f
C83 B.n49 VSUBS 0.018416f
C84 B.n50 VSUBS 0.007859f
C85 B.n51 VSUBS 0.007859f
C86 B.n52 VSUBS 0.007859f
C87 B.n53 VSUBS 0.007859f
C88 B.n54 VSUBS 0.007859f
C89 B.n55 VSUBS 0.007859f
C90 B.n56 VSUBS 0.007859f
C91 B.n57 VSUBS 0.007859f
C92 B.n58 VSUBS 0.007859f
C93 B.n59 VSUBS 0.007859f
C94 B.n60 VSUBS 0.007859f
C95 B.n61 VSUBS 0.007859f
C96 B.n62 VSUBS 0.007859f
C97 B.n63 VSUBS 0.007859f
C98 B.n64 VSUBS 0.007859f
C99 B.n65 VSUBS 0.019723f
C100 B.n66 VSUBS 0.007859f
C101 B.n67 VSUBS 0.007859f
C102 B.n68 VSUBS 0.007859f
C103 B.n69 VSUBS 0.007859f
C104 B.n70 VSUBS 0.007859f
C105 B.n71 VSUBS 0.007859f
C106 B.n72 VSUBS 0.007859f
C107 B.n73 VSUBS 0.007859f
C108 B.n74 VSUBS 0.007859f
C109 B.n75 VSUBS 0.007859f
C110 B.n76 VSUBS 0.007859f
C111 B.n77 VSUBS 0.007859f
C112 B.n78 VSUBS 0.007859f
C113 B.n79 VSUBS 0.007859f
C114 B.n80 VSUBS 0.005201f
C115 B.n81 VSUBS 0.007859f
C116 B.n82 VSUBS 0.007859f
C117 B.n83 VSUBS 0.007859f
C118 B.n84 VSUBS 0.007859f
C119 B.n85 VSUBS 0.007859f
C120 B.t5 VSUBS 0.287266f
C121 B.t4 VSUBS 0.298691f
C122 B.t3 VSUBS 0.389785f
C123 B.n86 VSUBS 0.129557f
C124 B.n87 VSUBS 0.072588f
C125 B.n88 VSUBS 0.007859f
C126 B.n89 VSUBS 0.007859f
C127 B.n90 VSUBS 0.007859f
C128 B.n91 VSUBS 0.007859f
C129 B.n92 VSUBS 0.007859f
C130 B.n93 VSUBS 0.007859f
C131 B.n94 VSUBS 0.007859f
C132 B.n95 VSUBS 0.007859f
C133 B.n96 VSUBS 0.007859f
C134 B.n97 VSUBS 0.007859f
C135 B.n98 VSUBS 0.007859f
C136 B.n99 VSUBS 0.007859f
C137 B.n100 VSUBS 0.007859f
C138 B.n101 VSUBS 0.007859f
C139 B.n102 VSUBS 0.019723f
C140 B.n103 VSUBS 0.007859f
C141 B.n104 VSUBS 0.007859f
C142 B.n105 VSUBS 0.007859f
C143 B.n106 VSUBS 0.007859f
C144 B.n107 VSUBS 0.007859f
C145 B.n108 VSUBS 0.007859f
C146 B.n109 VSUBS 0.007859f
C147 B.n110 VSUBS 0.007859f
C148 B.n111 VSUBS 0.007859f
C149 B.n112 VSUBS 0.007859f
C150 B.n113 VSUBS 0.007859f
C151 B.n114 VSUBS 0.007859f
C152 B.n115 VSUBS 0.007859f
C153 B.n116 VSUBS 0.007859f
C154 B.n117 VSUBS 0.007859f
C155 B.n118 VSUBS 0.007859f
C156 B.n119 VSUBS 0.007859f
C157 B.n120 VSUBS 0.007859f
C158 B.n121 VSUBS 0.007859f
C159 B.n122 VSUBS 0.007859f
C160 B.n123 VSUBS 0.007859f
C161 B.n124 VSUBS 0.007859f
C162 B.n125 VSUBS 0.007859f
C163 B.n126 VSUBS 0.007859f
C164 B.n127 VSUBS 0.007859f
C165 B.n128 VSUBS 0.007859f
C166 B.n129 VSUBS 0.018416f
C167 B.n130 VSUBS 0.018416f
C168 B.n131 VSUBS 0.019723f
C169 B.n132 VSUBS 0.007859f
C170 B.n133 VSUBS 0.007859f
C171 B.n134 VSUBS 0.007859f
C172 B.n135 VSUBS 0.007859f
C173 B.n136 VSUBS 0.007859f
C174 B.n137 VSUBS 0.007859f
C175 B.n138 VSUBS 0.007859f
C176 B.n139 VSUBS 0.007859f
C177 B.n140 VSUBS 0.007859f
C178 B.n141 VSUBS 0.007859f
C179 B.n142 VSUBS 0.007859f
C180 B.n143 VSUBS 0.007859f
C181 B.n144 VSUBS 0.007859f
C182 B.n145 VSUBS 0.007859f
C183 B.n146 VSUBS 0.007859f
C184 B.n147 VSUBS 0.007859f
C185 B.n148 VSUBS 0.007859f
C186 B.n149 VSUBS 0.007859f
C187 B.n150 VSUBS 0.007859f
C188 B.n151 VSUBS 0.007859f
C189 B.n152 VSUBS 0.007859f
C190 B.n153 VSUBS 0.007859f
C191 B.n154 VSUBS 0.007859f
C192 B.n155 VSUBS 0.007859f
C193 B.n156 VSUBS 0.007859f
C194 B.n157 VSUBS 0.007859f
C195 B.n158 VSUBS 0.007859f
C196 B.n159 VSUBS 0.007859f
C197 B.n160 VSUBS 0.007859f
C198 B.n161 VSUBS 0.007859f
C199 B.n162 VSUBS 0.007859f
C200 B.n163 VSUBS 0.007859f
C201 B.n164 VSUBS 0.007859f
C202 B.n165 VSUBS 0.007859f
C203 B.n166 VSUBS 0.007859f
C204 B.n167 VSUBS 0.007859f
C205 B.n168 VSUBS 0.007859f
C206 B.n169 VSUBS 0.007859f
C207 B.n170 VSUBS 0.007859f
C208 B.n171 VSUBS 0.007859f
C209 B.n172 VSUBS 0.007859f
C210 B.n173 VSUBS 0.007859f
C211 B.n174 VSUBS 0.007859f
C212 B.n175 VSUBS 0.007859f
C213 B.n176 VSUBS 0.005201f
C214 B.n177 VSUBS 0.018208f
C215 B.n178 VSUBS 0.006588f
C216 B.n179 VSUBS 0.007859f
C217 B.n180 VSUBS 0.007859f
C218 B.n181 VSUBS 0.007859f
C219 B.n182 VSUBS 0.007859f
C220 B.n183 VSUBS 0.007859f
C221 B.n184 VSUBS 0.007859f
C222 B.n185 VSUBS 0.007859f
C223 B.n186 VSUBS 0.007859f
C224 B.n187 VSUBS 0.007859f
C225 B.n188 VSUBS 0.007859f
C226 B.n189 VSUBS 0.007859f
C227 B.t2 VSUBS 0.287263f
C228 B.t1 VSUBS 0.298688f
C229 B.t0 VSUBS 0.389785f
C230 B.n190 VSUBS 0.129559f
C231 B.n191 VSUBS 0.072591f
C232 B.n192 VSUBS 0.018208f
C233 B.n193 VSUBS 0.006588f
C234 B.n194 VSUBS 0.007859f
C235 B.n195 VSUBS 0.007859f
C236 B.n196 VSUBS 0.007859f
C237 B.n197 VSUBS 0.007859f
C238 B.n198 VSUBS 0.007859f
C239 B.n199 VSUBS 0.007859f
C240 B.n200 VSUBS 0.007859f
C241 B.n201 VSUBS 0.007859f
C242 B.n202 VSUBS 0.007859f
C243 B.n203 VSUBS 0.007859f
C244 B.n204 VSUBS 0.007859f
C245 B.n205 VSUBS 0.007859f
C246 B.n206 VSUBS 0.007859f
C247 B.n207 VSUBS 0.007859f
C248 B.n208 VSUBS 0.007859f
C249 B.n209 VSUBS 0.007859f
C250 B.n210 VSUBS 0.007859f
C251 B.n211 VSUBS 0.007859f
C252 B.n212 VSUBS 0.007859f
C253 B.n213 VSUBS 0.007859f
C254 B.n214 VSUBS 0.007859f
C255 B.n215 VSUBS 0.007859f
C256 B.n216 VSUBS 0.007859f
C257 B.n217 VSUBS 0.007859f
C258 B.n218 VSUBS 0.007859f
C259 B.n219 VSUBS 0.007859f
C260 B.n220 VSUBS 0.007859f
C261 B.n221 VSUBS 0.007859f
C262 B.n222 VSUBS 0.007859f
C263 B.n223 VSUBS 0.007859f
C264 B.n224 VSUBS 0.007859f
C265 B.n225 VSUBS 0.007859f
C266 B.n226 VSUBS 0.007859f
C267 B.n227 VSUBS 0.007859f
C268 B.n228 VSUBS 0.007859f
C269 B.n229 VSUBS 0.007859f
C270 B.n230 VSUBS 0.007859f
C271 B.n231 VSUBS 0.007859f
C272 B.n232 VSUBS 0.007859f
C273 B.n233 VSUBS 0.007859f
C274 B.n234 VSUBS 0.007859f
C275 B.n235 VSUBS 0.007859f
C276 B.n236 VSUBS 0.007859f
C277 B.n237 VSUBS 0.007859f
C278 B.n238 VSUBS 0.007859f
C279 B.n239 VSUBS 0.007859f
C280 B.n240 VSUBS 0.018844f
C281 B.n241 VSUBS 0.019295f
C282 B.n242 VSUBS 0.018416f
C283 B.n243 VSUBS 0.007859f
C284 B.n244 VSUBS 0.007859f
C285 B.n245 VSUBS 0.007859f
C286 B.n246 VSUBS 0.007859f
C287 B.n247 VSUBS 0.007859f
C288 B.n248 VSUBS 0.007859f
C289 B.n249 VSUBS 0.007859f
C290 B.n250 VSUBS 0.007859f
C291 B.n251 VSUBS 0.007859f
C292 B.n252 VSUBS 0.007859f
C293 B.n253 VSUBS 0.007859f
C294 B.n254 VSUBS 0.007859f
C295 B.n255 VSUBS 0.007859f
C296 B.n256 VSUBS 0.007859f
C297 B.n257 VSUBS 0.007859f
C298 B.n258 VSUBS 0.007859f
C299 B.n259 VSUBS 0.007859f
C300 B.n260 VSUBS 0.007859f
C301 B.n261 VSUBS 0.007859f
C302 B.n262 VSUBS 0.007859f
C303 B.n263 VSUBS 0.007859f
C304 B.n264 VSUBS 0.007859f
C305 B.n265 VSUBS 0.007859f
C306 B.n266 VSUBS 0.007859f
C307 B.n267 VSUBS 0.007859f
C308 B.n268 VSUBS 0.007859f
C309 B.n269 VSUBS 0.007859f
C310 B.n270 VSUBS 0.007859f
C311 B.n271 VSUBS 0.007859f
C312 B.n272 VSUBS 0.007859f
C313 B.n273 VSUBS 0.007859f
C314 B.n274 VSUBS 0.007859f
C315 B.n275 VSUBS 0.007859f
C316 B.n276 VSUBS 0.007859f
C317 B.n277 VSUBS 0.007859f
C318 B.n278 VSUBS 0.007859f
C319 B.n279 VSUBS 0.007859f
C320 B.n280 VSUBS 0.007859f
C321 B.n281 VSUBS 0.007859f
C322 B.n282 VSUBS 0.007859f
C323 B.n283 VSUBS 0.007859f
C324 B.n284 VSUBS 0.007859f
C325 B.n285 VSUBS 0.007859f
C326 B.n286 VSUBS 0.007859f
C327 B.n287 VSUBS 0.007859f
C328 B.n288 VSUBS 0.018416f
C329 B.n289 VSUBS 0.019723f
C330 B.n290 VSUBS 0.019723f
C331 B.n291 VSUBS 0.007859f
C332 B.n292 VSUBS 0.007859f
C333 B.n293 VSUBS 0.007859f
C334 B.n294 VSUBS 0.007859f
C335 B.n295 VSUBS 0.007859f
C336 B.n296 VSUBS 0.007859f
C337 B.n297 VSUBS 0.007859f
C338 B.n298 VSUBS 0.007859f
C339 B.n299 VSUBS 0.007859f
C340 B.n300 VSUBS 0.007859f
C341 B.n301 VSUBS 0.007859f
C342 B.n302 VSUBS 0.007859f
C343 B.n303 VSUBS 0.007859f
C344 B.n304 VSUBS 0.007859f
C345 B.n305 VSUBS 0.007859f
C346 B.n306 VSUBS 0.007859f
C347 B.n307 VSUBS 0.007859f
C348 B.n308 VSUBS 0.007859f
C349 B.n309 VSUBS 0.007859f
C350 B.n310 VSUBS 0.007859f
C351 B.n311 VSUBS 0.007859f
C352 B.n312 VSUBS 0.007859f
C353 B.n313 VSUBS 0.007859f
C354 B.n314 VSUBS 0.007859f
C355 B.n315 VSUBS 0.007859f
C356 B.n316 VSUBS 0.007859f
C357 B.n317 VSUBS 0.007859f
C358 B.n318 VSUBS 0.007859f
C359 B.n319 VSUBS 0.007859f
C360 B.n320 VSUBS 0.007859f
C361 B.n321 VSUBS 0.007859f
C362 B.n322 VSUBS 0.007859f
C363 B.n323 VSUBS 0.007859f
C364 B.n324 VSUBS 0.007859f
C365 B.n325 VSUBS 0.007859f
C366 B.n326 VSUBS 0.007859f
C367 B.n327 VSUBS 0.007859f
C368 B.n328 VSUBS 0.007859f
C369 B.n329 VSUBS 0.007859f
C370 B.n330 VSUBS 0.007859f
C371 B.n331 VSUBS 0.007859f
C372 B.n332 VSUBS 0.007859f
C373 B.n333 VSUBS 0.007859f
C374 B.n334 VSUBS 0.007859f
C375 B.n335 VSUBS 0.005201f
C376 B.n336 VSUBS 0.018208f
C377 B.n337 VSUBS 0.006588f
C378 B.n338 VSUBS 0.007859f
C379 B.n339 VSUBS 0.007859f
C380 B.n340 VSUBS 0.007859f
C381 B.n341 VSUBS 0.007859f
C382 B.n342 VSUBS 0.007859f
C383 B.n343 VSUBS 0.007859f
C384 B.n344 VSUBS 0.007859f
C385 B.n345 VSUBS 0.007859f
C386 B.n346 VSUBS 0.007859f
C387 B.n347 VSUBS 0.007859f
C388 B.n348 VSUBS 0.007859f
C389 B.n349 VSUBS 0.006588f
C390 B.n350 VSUBS 0.018208f
C391 B.n351 VSUBS 0.005201f
C392 B.n352 VSUBS 0.007859f
C393 B.n353 VSUBS 0.007859f
C394 B.n354 VSUBS 0.007859f
C395 B.n355 VSUBS 0.007859f
C396 B.n356 VSUBS 0.007859f
C397 B.n357 VSUBS 0.007859f
C398 B.n358 VSUBS 0.007859f
C399 B.n359 VSUBS 0.007859f
C400 B.n360 VSUBS 0.007859f
C401 B.n361 VSUBS 0.007859f
C402 B.n362 VSUBS 0.007859f
C403 B.n363 VSUBS 0.007859f
C404 B.n364 VSUBS 0.007859f
C405 B.n365 VSUBS 0.007859f
C406 B.n366 VSUBS 0.007859f
C407 B.n367 VSUBS 0.007859f
C408 B.n368 VSUBS 0.007859f
C409 B.n369 VSUBS 0.007859f
C410 B.n370 VSUBS 0.007859f
C411 B.n371 VSUBS 0.007859f
C412 B.n372 VSUBS 0.007859f
C413 B.n373 VSUBS 0.007859f
C414 B.n374 VSUBS 0.007859f
C415 B.n375 VSUBS 0.007859f
C416 B.n376 VSUBS 0.007859f
C417 B.n377 VSUBS 0.007859f
C418 B.n378 VSUBS 0.007859f
C419 B.n379 VSUBS 0.007859f
C420 B.n380 VSUBS 0.007859f
C421 B.n381 VSUBS 0.007859f
C422 B.n382 VSUBS 0.007859f
C423 B.n383 VSUBS 0.007859f
C424 B.n384 VSUBS 0.007859f
C425 B.n385 VSUBS 0.007859f
C426 B.n386 VSUBS 0.007859f
C427 B.n387 VSUBS 0.007859f
C428 B.n388 VSUBS 0.007859f
C429 B.n389 VSUBS 0.007859f
C430 B.n390 VSUBS 0.007859f
C431 B.n391 VSUBS 0.007859f
C432 B.n392 VSUBS 0.007859f
C433 B.n393 VSUBS 0.007859f
C434 B.n394 VSUBS 0.007859f
C435 B.n395 VSUBS 0.007859f
C436 B.n396 VSUBS 0.019723f
C437 B.n397 VSUBS 0.019723f
C438 B.n398 VSUBS 0.018416f
C439 B.n399 VSUBS 0.007859f
C440 B.n400 VSUBS 0.007859f
C441 B.n401 VSUBS 0.007859f
C442 B.n402 VSUBS 0.007859f
C443 B.n403 VSUBS 0.007859f
C444 B.n404 VSUBS 0.007859f
C445 B.n405 VSUBS 0.007859f
C446 B.n406 VSUBS 0.007859f
C447 B.n407 VSUBS 0.007859f
C448 B.n408 VSUBS 0.007859f
C449 B.n409 VSUBS 0.007859f
C450 B.n410 VSUBS 0.007859f
C451 B.n411 VSUBS 0.007859f
C452 B.n412 VSUBS 0.007859f
C453 B.n413 VSUBS 0.007859f
C454 B.n414 VSUBS 0.007859f
C455 B.n415 VSUBS 0.007859f
C456 B.n416 VSUBS 0.007859f
C457 B.n417 VSUBS 0.007859f
C458 B.n418 VSUBS 0.007859f
C459 B.n419 VSUBS 0.010256f
C460 B.n420 VSUBS 0.010925f
C461 B.n421 VSUBS 0.021725f
C462 VDD2.t1 VSUBS 1.18815f
C463 VDD2.t0 VSUBS 0.929529f
C464 VDD2.n0 VSUBS 1.93892f
C465 VN.t0 VSUBS 0.78867f
C466 VN.t1 VSUBS 0.890485f
C467 VDD1.t0 VSUBS 0.918468f
C468 VDD1.t1 VSUBS 1.18756f
C469 VTAIL.t1 VSUBS 1.45748f
C470 VTAIL.n0 VSUBS 1.74493f
C471 VTAIL.t0 VSUBS 1.45749f
C472 VTAIL.n1 VSUBS 1.7629f
C473 VTAIL.t2 VSUBS 1.45748f
C474 VTAIL.n2 VSUBS 1.67212f
C475 VTAIL.t3 VSUBS 1.45748f
C476 VTAIL.n3 VSUBS 1.60665f
C477 VP.t1 VSUBS 1.34577f
C478 VP.t0 VSUBS 1.19533f
C479 VP.n0 VSUBS 3.43594f
.ends

