* NGSPICE file created from tg_sample_0009.ext - technology: sky130A

.subckt tg_sample_0009 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t27 VOUT.t26 VOUT.t27 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.3036 pd=2.17 as=0 ps=0 w=1.84 l=0.26
X1 VOUT.t25 VOUT.t24 VOUT.t25 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.3036 pd=2.17 as=0 ps=0 w=1.84 l=0.26
X2 VOUT.t23 VOUT.t21 VOUT.t22 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X3 VSS.t16 VSS.t14 VSS.t15 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X4 VOUT.t20 VOUT.t19 VOUT.t20 VCC.t2 sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=0 ps=0 w=13.44 l=0.21
X5 VOUT.t18 VOUT.t17 VOUT.t18 VCC.t1 sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=0 ps=0 w=13.44 l=0.21
X6 VCC.t16 VCC.t14 VCC.t15 VCC.t8 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
X7 VSS.t13 VSS.t10 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X8 VOUT.t16 VOUT.t15 VOUT.t16 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.3036 pd=2.17 as=0 ps=0 w=1.84 l=0.26
X9 VSS.t9 VSS.t7 VSS.t8 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X10 VOUT.t14 VOUT.t13 VOUT.t14 VCC.t2 sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=0 ps=0 w=13.44 l=0.21
X11 VOUT.t12 VOUT.t10 VOUT.t11 VCC.t0 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
X12 VCC.t13 VCC.t11 VCC.t12 VCC.t4 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
X13 VOUT.t9 VOUT.t7 VOUT.t8 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X14 VOUT.t6 VOUT.t5 VOUT.t6 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.3036 pd=2.17 as=0 ps=0 w=1.84 l=0.26
X15 VSS.t6 VSS.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=0.26
X16 VOUT.t4 VOUT.t3 VOUT.t4 VCC.t1 sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=0 ps=0 w=13.44 l=0.21
X17 VCC.t10 VCC.t7 VCC.t9 VCC.t8 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
X18 VOUT.t2 VOUT.t0 VOUT.t1 VCC.t0 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
X19 VCC.t6 VCC.t3 VCC.t5 VCC.t4 sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=0.21
R0 VOUT.n177 VOUT.t10 1733.95
R1 VOUT.n179 VOUT.t19 1733.95
R2 VOUT.n168 VOUT.t0 1733.95
R3 VOUT.n170 VOUT.t13 1733.95
R4 VOUT.n178 VOUT.t3 1691.59
R5 VOUT.n169 VOUT.t17 1691.59
R6 VOUT.n120 VOUT.n118 756.745
R7 VOUT.n333 VOUT.n265 756.745
R8 VOUT.n251 VOUT.n183 756.745
R9 VOUT.n90 VOUT.n22 756.745
R10 VOUT.n167 VOUT.n166 585
R11 VOUT.n98 VOUT.n97 585
R12 VOUT.n161 VOUT.n160 585
R13 VOUT.n159 VOUT.n158 585
R14 VOUT.n102 VOUT.n101 585
R15 VOUT.n153 VOUT.n152 585
R16 VOUT.n151 VOUT.n150 585
R17 VOUT.n106 VOUT.n105 585
R18 VOUT.n145 VOUT.n144 585
R19 VOUT.n143 VOUT.n108 585
R20 VOUT.n142 VOUT.n141 585
R21 VOUT.n111 VOUT.n109 585
R22 VOUT.n136 VOUT.n135 585
R23 VOUT.n134 VOUT.n133 585
R24 VOUT.n115 VOUT.n114 585
R25 VOUT.n128 VOUT.n127 585
R26 VOUT.n126 VOUT.n125 585
R27 VOUT.n119 VOUT.n118 585
R28 VOUT.n290 VOUT.n289 585
R29 VOUT.n292 VOUT.n291 585
R30 VOUT.n285 VOUT.n284 585
R31 VOUT.n298 VOUT.n297 585
R32 VOUT.n300 VOUT.n299 585
R33 VOUT.n281 VOUT.n280 585
R34 VOUT.n307 VOUT.n306 585
R35 VOUT.n308 VOUT.n279 585
R36 VOUT.n310 VOUT.n309 585
R37 VOUT.n277 VOUT.n276 585
R38 VOUT.n316 VOUT.n315 585
R39 VOUT.n318 VOUT.n317 585
R40 VOUT.n273 VOUT.n272 585
R41 VOUT.n324 VOUT.n323 585
R42 VOUT.n326 VOUT.n325 585
R43 VOUT.n269 VOUT.n268 585
R44 VOUT.n332 VOUT.n331 585
R45 VOUT.n334 VOUT.n333 585
R46 VOUT.n208 VOUT.n207 585
R47 VOUT.n210 VOUT.n209 585
R48 VOUT.n203 VOUT.n202 585
R49 VOUT.n216 VOUT.n215 585
R50 VOUT.n218 VOUT.n217 585
R51 VOUT.n199 VOUT.n198 585
R52 VOUT.n225 VOUT.n224 585
R53 VOUT.n226 VOUT.n197 585
R54 VOUT.n228 VOUT.n227 585
R55 VOUT.n195 VOUT.n194 585
R56 VOUT.n234 VOUT.n233 585
R57 VOUT.n236 VOUT.n235 585
R58 VOUT.n191 VOUT.n190 585
R59 VOUT.n242 VOUT.n241 585
R60 VOUT.n244 VOUT.n243 585
R61 VOUT.n187 VOUT.n186 585
R62 VOUT.n250 VOUT.n249 585
R63 VOUT.n252 VOUT.n251 585
R64 VOUT.n47 VOUT.n46 585
R65 VOUT.n49 VOUT.n48 585
R66 VOUT.n42 VOUT.n41 585
R67 VOUT.n55 VOUT.n54 585
R68 VOUT.n57 VOUT.n56 585
R69 VOUT.n38 VOUT.n37 585
R70 VOUT.n64 VOUT.n63 585
R71 VOUT.n65 VOUT.n36 585
R72 VOUT.n67 VOUT.n66 585
R73 VOUT.n34 VOUT.n33 585
R74 VOUT.n73 VOUT.n72 585
R75 VOUT.n75 VOUT.n74 585
R76 VOUT.n30 VOUT.n29 585
R77 VOUT.n81 VOUT.n80 585
R78 VOUT.n83 VOUT.n82 585
R79 VOUT.n26 VOUT.n25 585
R80 VOUT.n89 VOUT.n88 585
R81 VOUT.n91 VOUT.n90 585
R82 VOUT.n174 VOUT.t24 340.714
R83 VOUT.n172 VOUT.t21 340.714
R84 VOUT.n2 VOUT.t26 340.714
R85 VOUT.n0 VOUT.t7 340.714
R86 VOUT.t14 VOUT.n96 329.036
R87 VOUT.n288 VOUT.t12 329.036
R88 VOUT.n206 VOUT.t2 329.036
R89 VOUT.n45 VOUT.t20 329.036
R90 VOUT.n173 VOUT.t5 291.055
R91 VOUT.n1 VOUT.t15 291.055
R92 VOUT.n351 VOUT.n349 289.615
R93 VOUT.n343 VOUT.n340 289.615
R94 VOUT.n15 VOUT.n13 289.615
R95 VOUT.n7 VOUT.n5 289.615
R96 VOUT.n352 VOUT.n351 185
R97 VOUT.n345 VOUT.n340 185
R98 VOUT.n16 VOUT.n15 185
R99 VOUT.n8 VOUT.n7 185
R100 VOUT.n167 VOUT.n97 171.744
R101 VOUT.n160 VOUT.n97 171.744
R102 VOUT.n160 VOUT.n159 171.744
R103 VOUT.n159 VOUT.n101 171.744
R104 VOUT.n152 VOUT.n101 171.744
R105 VOUT.n152 VOUT.n151 171.744
R106 VOUT.n151 VOUT.n105 171.744
R107 VOUT.n144 VOUT.n105 171.744
R108 VOUT.n144 VOUT.n143 171.744
R109 VOUT.n143 VOUT.n142 171.744
R110 VOUT.n142 VOUT.n109 171.744
R111 VOUT.n135 VOUT.n109 171.744
R112 VOUT.n135 VOUT.n134 171.744
R113 VOUT.n134 VOUT.n114 171.744
R114 VOUT.n127 VOUT.n114 171.744
R115 VOUT.n127 VOUT.n126 171.744
R116 VOUT.n126 VOUT.n118 171.744
R117 VOUT.n291 VOUT.n290 171.744
R118 VOUT.n291 VOUT.n284 171.744
R119 VOUT.n298 VOUT.n284 171.744
R120 VOUT.n299 VOUT.n298 171.744
R121 VOUT.n299 VOUT.n280 171.744
R122 VOUT.n307 VOUT.n280 171.744
R123 VOUT.n308 VOUT.n307 171.744
R124 VOUT.n309 VOUT.n308 171.744
R125 VOUT.n309 VOUT.n276 171.744
R126 VOUT.n316 VOUT.n276 171.744
R127 VOUT.n317 VOUT.n316 171.744
R128 VOUT.n317 VOUT.n272 171.744
R129 VOUT.n324 VOUT.n272 171.744
R130 VOUT.n325 VOUT.n324 171.744
R131 VOUT.n325 VOUT.n268 171.744
R132 VOUT.n332 VOUT.n268 171.744
R133 VOUT.n333 VOUT.n332 171.744
R134 VOUT.n209 VOUT.n208 171.744
R135 VOUT.n209 VOUT.n202 171.744
R136 VOUT.n216 VOUT.n202 171.744
R137 VOUT.n217 VOUT.n216 171.744
R138 VOUT.n217 VOUT.n198 171.744
R139 VOUT.n225 VOUT.n198 171.744
R140 VOUT.n226 VOUT.n225 171.744
R141 VOUT.n227 VOUT.n226 171.744
R142 VOUT.n227 VOUT.n194 171.744
R143 VOUT.n234 VOUT.n194 171.744
R144 VOUT.n235 VOUT.n234 171.744
R145 VOUT.n235 VOUT.n190 171.744
R146 VOUT.n242 VOUT.n190 171.744
R147 VOUT.n243 VOUT.n242 171.744
R148 VOUT.n243 VOUT.n186 171.744
R149 VOUT.n250 VOUT.n186 171.744
R150 VOUT.n251 VOUT.n250 171.744
R151 VOUT.n48 VOUT.n47 171.744
R152 VOUT.n48 VOUT.n41 171.744
R153 VOUT.n55 VOUT.n41 171.744
R154 VOUT.n56 VOUT.n55 171.744
R155 VOUT.n56 VOUT.n37 171.744
R156 VOUT.n64 VOUT.n37 171.744
R157 VOUT.n65 VOUT.n64 171.744
R158 VOUT.n66 VOUT.n65 171.744
R159 VOUT.n66 VOUT.n33 171.744
R160 VOUT.n73 VOUT.n33 171.744
R161 VOUT.n74 VOUT.n73 171.744
R162 VOUT.n74 VOUT.n29 171.744
R163 VOUT.n81 VOUT.n29 171.744
R164 VOUT.n82 VOUT.n81 171.744
R165 VOUT.n82 VOUT.n25 171.744
R166 VOUT.n89 VOUT.n25 171.744
R167 VOUT.n90 VOUT.n89 171.744
R168 VOUT.t23 VOUT.n350 164.876
R169 VOUT.t25 VOUT.n346 164.876
R170 VOUT.n14 VOUT.t27 164.876
R171 VOUT.t9 VOUT.n6 164.876
R172 VOUT.n175 VOUT.n172 161.489
R173 VOUT.n180 VOUT.n177 161.489
R174 VOUT.n171 VOUT.n168 161.489
R175 VOUT.n3 VOUT.n0 161.489
R176 VOUT.n175 VOUT.n174 161.3
R177 VOUT.n180 VOUT.n179 161.3
R178 VOUT.n171 VOUT.n170 161.3
R179 VOUT.n3 VOUT.n2 161.3
R180 VOUT.n347 VOUT.n20 102.587
R181 VOUT.n361 VOUT.n360 102.587
R182 VOUT.n356 VOUT.n348 86.4166
R183 VOUT.n363 VOUT.n362 85.9079
R184 VOUT.t14 VOUT.n167 85.8723
R185 VOUT.n290 VOUT.t12 85.8723
R186 VOUT.n208 VOUT.t2 85.8723
R187 VOUT.n47 VOUT.t20 85.8723
R188 VOUT.n260 VOUT.n259 69.9534
R189 VOUT.n263 VOUT.n262 69.9534
R190 VOUT.n338 VOUT.n264 53.7401
R191 VOUT.n258 VOUT.n257 53.2746
R192 VOUT.n342 VOUT.n20 52.4758
R193 VOUT.n360 VOUT.n19 52.4758
R194 VOUT.n351 VOUT.t23 52.3082
R195 VOUT.t25 VOUT.n340 52.3082
R196 VOUT.n15 VOUT.t27 52.3082
R197 VOUT.n7 VOUT.t9 52.3082
R198 VOUT.n260 VOUT.n95 47.0024
R199 VOUT.n262 VOUT.n94 47.0024
R200 VOUT.n174 VOUT.n173 36.5157
R201 VOUT.n173 VOUT.n172 36.5157
R202 VOUT.n179 VOUT.n178 36.5157
R203 VOUT.n178 VOUT.n177 36.5157
R204 VOUT.n170 VOUT.n169 36.5157
R205 VOUT.n169 VOUT.n168 36.5157
R206 VOUT.n2 VOUT.n1 36.5157
R207 VOUT.n1 VOUT.n0 36.5157
R208 VOUT.n356 VOUT.n355 35.2884
R209 VOUT.n12 VOUT.n11 35.2884
R210 VOUT.n338 VOUT.n337 29.8581
R211 VOUT.n256 VOUT.n255 29.8581
R212 VOUT.n262 VOUT.n261 17.2979
R213 VOUT.n352 VOUT.n350 14.7318
R214 VOUT.n346 VOUT.n345 14.7318
R215 VOUT.n16 VOUT.n14 14.7318
R216 VOUT.n8 VOUT.n6 14.7318
R217 VOUT.n145 VOUT.n108 13.1884
R218 VOUT.n310 VOUT.n277 13.1884
R219 VOUT.n228 VOUT.n195 13.1884
R220 VOUT.n67 VOUT.n34 13.1884
R221 VOUT.n146 VOUT.n106 12.8005
R222 VOUT.n141 VOUT.n110 12.8005
R223 VOUT.n311 VOUT.n279 12.8005
R224 VOUT.n315 VOUT.n314 12.8005
R225 VOUT.n353 VOUT.n349 12.8005
R226 VOUT.n344 VOUT.n343 12.8005
R227 VOUT.n17 VOUT.n13 12.8005
R228 VOUT.n9 VOUT.n5 12.8005
R229 VOUT.n229 VOUT.n197 12.8005
R230 VOUT.n233 VOUT.n232 12.8005
R231 VOUT.n68 VOUT.n36 12.8005
R232 VOUT.n72 VOUT.n71 12.8005
R233 VOUT.n359 VOUT.n20 12.3626
R234 VOUT.n150 VOUT.n149 12.0247
R235 VOUT.n140 VOUT.n111 12.0247
R236 VOUT.n306 VOUT.n305 12.0247
R237 VOUT.n318 VOUT.n275 12.0247
R238 VOUT.n224 VOUT.n223 12.0247
R239 VOUT.n236 VOUT.n193 12.0247
R240 VOUT.n63 VOUT.n62 12.0247
R241 VOUT.n75 VOUT.n32 12.0247
R242 VOUT.n153 VOUT.n104 11.249
R243 VOUT.n137 VOUT.n136 11.249
R244 VOUT.n304 VOUT.n281 11.249
R245 VOUT.n319 VOUT.n273 11.249
R246 VOUT.n222 VOUT.n199 11.249
R247 VOUT.n237 VOUT.n191 11.249
R248 VOUT.n61 VOUT.n38 11.249
R249 VOUT.n76 VOUT.n30 11.249
R250 VOUT.n348 VOUT.t25 10.7614
R251 VOUT.n348 VOUT.t6 10.7614
R252 VOUT.t6 VOUT.n347 10.7614
R253 VOUT.n347 VOUT.t22 10.7614
R254 VOUT.t16 VOUT.n361 10.7614
R255 VOUT.n361 VOUT.t8 10.7614
R256 VOUT.n362 VOUT.t27 10.7614
R257 VOUT.n362 VOUT.t16 10.7614
R258 VOUT.n166 VOUT.n96 10.7239
R259 VOUT.n289 VOUT.n288 10.7239
R260 VOUT.n207 VOUT.n206 10.7239
R261 VOUT.n46 VOUT.n45 10.7239
R262 VOUT.n154 VOUT.n102 10.4732
R263 VOUT.n133 VOUT.n113 10.4732
R264 VOUT.n301 VOUT.n300 10.4732
R265 VOUT.n323 VOUT.n322 10.4732
R266 VOUT.n219 VOUT.n218 10.4732
R267 VOUT.n241 VOUT.n240 10.4732
R268 VOUT.n58 VOUT.n57 10.4732
R269 VOUT.n80 VOUT.n79 10.4732
R270 VOUT.n182 VGP 10.2901
R271 VOUT.n158 VOUT.n157 9.69747
R272 VOUT.n132 VOUT.n115 9.69747
R273 VOUT.n297 VOUT.n283 9.69747
R274 VOUT.n326 VOUT.n271 9.69747
R275 VOUT.n215 VOUT.n201 9.69747
R276 VOUT.n244 VOUT.n189 9.69747
R277 VOUT.n54 VOUT.n40 9.69747
R278 VOUT.n83 VOUT.n28 9.69747
R279 VOUT.n122 VOUT.n95 9.45567
R280 VOUT.n337 VOUT.n336 9.45567
R281 VOUT.n355 VOUT.n354 9.45567
R282 VOUT.n342 VOUT.n341 9.45567
R283 VOUT.n19 VOUT.n18 9.45567
R284 VOUT.n11 VOUT.n10 9.45567
R285 VOUT.n255 VOUT.n254 9.45567
R286 VOUT.n94 VOUT.n93 9.45567
R287 VOUT.n122 VOUT.n121 9.3005
R288 VOUT.n117 VOUT.n116 9.3005
R289 VOUT.n130 VOUT.n129 9.3005
R290 VOUT.n132 VOUT.n131 9.3005
R291 VOUT.n113 VOUT.n112 9.3005
R292 VOUT.n138 VOUT.n137 9.3005
R293 VOUT.n140 VOUT.n139 9.3005
R294 VOUT.n110 VOUT.n107 9.3005
R295 VOUT.n165 VOUT.n164 9.3005
R296 VOUT.n163 VOUT.n162 9.3005
R297 VOUT.n100 VOUT.n99 9.3005
R298 VOUT.n157 VOUT.n156 9.3005
R299 VOUT.n155 VOUT.n154 9.3005
R300 VOUT.n104 VOUT.n103 9.3005
R301 VOUT.n149 VOUT.n148 9.3005
R302 VOUT.n147 VOUT.n146 9.3005
R303 VOUT.n124 VOUT.n123 9.3005
R304 VOUT.n336 VOUT.n335 9.3005
R305 VOUT.n330 VOUT.n329 9.3005
R306 VOUT.n328 VOUT.n327 9.3005
R307 VOUT.n271 VOUT.n270 9.3005
R308 VOUT.n322 VOUT.n321 9.3005
R309 VOUT.n320 VOUT.n319 9.3005
R310 VOUT.n275 VOUT.n274 9.3005
R311 VOUT.n314 VOUT.n313 9.3005
R312 VOUT.n287 VOUT.n286 9.3005
R313 VOUT.n294 VOUT.n293 9.3005
R314 VOUT.n296 VOUT.n295 9.3005
R315 VOUT.n283 VOUT.n282 9.3005
R316 VOUT.n302 VOUT.n301 9.3005
R317 VOUT.n304 VOUT.n303 9.3005
R318 VOUT.n305 VOUT.n278 9.3005
R319 VOUT.n312 VOUT.n311 9.3005
R320 VOUT.n267 VOUT.n266 9.3005
R321 VOUT.n354 VOUT.n353 9.3005
R322 VOUT.n344 VOUT.n341 9.3005
R323 VOUT.n18 VOUT.n17 9.3005
R324 VOUT.n10 VOUT.n9 9.3005
R325 VOUT.n254 VOUT.n253 9.3005
R326 VOUT.n248 VOUT.n247 9.3005
R327 VOUT.n246 VOUT.n245 9.3005
R328 VOUT.n189 VOUT.n188 9.3005
R329 VOUT.n240 VOUT.n239 9.3005
R330 VOUT.n238 VOUT.n237 9.3005
R331 VOUT.n193 VOUT.n192 9.3005
R332 VOUT.n232 VOUT.n231 9.3005
R333 VOUT.n205 VOUT.n204 9.3005
R334 VOUT.n212 VOUT.n211 9.3005
R335 VOUT.n214 VOUT.n213 9.3005
R336 VOUT.n201 VOUT.n200 9.3005
R337 VOUT.n220 VOUT.n219 9.3005
R338 VOUT.n222 VOUT.n221 9.3005
R339 VOUT.n223 VOUT.n196 9.3005
R340 VOUT.n230 VOUT.n229 9.3005
R341 VOUT.n185 VOUT.n184 9.3005
R342 VOUT.n93 VOUT.n92 9.3005
R343 VOUT.n87 VOUT.n86 9.3005
R344 VOUT.n85 VOUT.n84 9.3005
R345 VOUT.n28 VOUT.n27 9.3005
R346 VOUT.n79 VOUT.n78 9.3005
R347 VOUT.n77 VOUT.n76 9.3005
R348 VOUT.n32 VOUT.n31 9.3005
R349 VOUT.n71 VOUT.n70 9.3005
R350 VOUT.n44 VOUT.n43 9.3005
R351 VOUT.n51 VOUT.n50 9.3005
R352 VOUT.n53 VOUT.n52 9.3005
R353 VOUT.n40 VOUT.n39 9.3005
R354 VOUT.n59 VOUT.n58 9.3005
R355 VOUT.n61 VOUT.n60 9.3005
R356 VOUT.n62 VOUT.n35 9.3005
R357 VOUT.n69 VOUT.n68 9.3005
R358 VOUT.n24 VOUT.n23 9.3005
R359 VOUT.n181 VOUT.n176 9.18554
R360 VOUT.n161 VOUT.n100 8.92171
R361 VOUT.n129 VOUT.n128 8.92171
R362 VOUT.n296 VOUT.n285 8.92171
R363 VOUT.n327 VOUT.n269 8.92171
R364 VOUT.n214 VOUT.n203 8.92171
R365 VOUT.n245 VOUT.n187 8.92171
R366 VOUT.n53 VOUT.n42 8.92171
R367 VOUT.n84 VOUT.n26 8.92171
R368 VOUT.n162 VOUT.n98 8.14595
R369 VOUT.n125 VOUT.n117 8.14595
R370 VOUT.n293 VOUT.n292 8.14595
R371 VOUT.n331 VOUT.n330 8.14595
R372 VOUT.n211 VOUT.n210 8.14595
R373 VOUT.n249 VOUT.n248 8.14595
R374 VOUT.n50 VOUT.n49 8.14595
R375 VOUT.n88 VOUT.n87 8.14595
R376 VOUT.n166 VOUT.n165 7.3702
R377 VOUT.n124 VOUT.n119 7.3702
R378 VOUT.n120 VOUT.n95 7.3702
R379 VOUT.n289 VOUT.n287 7.3702
R380 VOUT.n334 VOUT.n267 7.3702
R381 VOUT.n337 VOUT.n265 7.3702
R382 VOUT.n207 VOUT.n205 7.3702
R383 VOUT.n252 VOUT.n185 7.3702
R384 VOUT.n255 VOUT.n183 7.3702
R385 VOUT.n46 VOUT.n44 7.3702
R386 VOUT.n91 VOUT.n24 7.3702
R387 VOUT.n94 VOUT.n22 7.3702
R388 VOUT.n121 VOUT.n119 6.59444
R389 VOUT.n121 VOUT.n120 6.59444
R390 VOUT.n335 VOUT.n334 6.59444
R391 VOUT.n335 VOUT.n265 6.59444
R392 VOUT.n253 VOUT.n252 6.59444
R393 VOUT.n253 VOUT.n183 6.59444
R394 VOUT.n92 VOUT.n91 6.59444
R395 VOUT.n92 VOUT.n22 6.59444
R396 VOUT.n339 VOUT.n21 6.46171
R397 VOUT.n4 VGN 5.90067
R398 VOUT.n165 VOUT.n98 5.81868
R399 VOUT.n125 VOUT.n124 5.81868
R400 VOUT.n292 VOUT.n287 5.81868
R401 VOUT.n331 VOUT.n267 5.81868
R402 VOUT.n210 VOUT.n205 5.81868
R403 VOUT.n249 VOUT.n185 5.81868
R404 VOUT.n49 VOUT.n44 5.81868
R405 VOUT.n88 VOUT.n24 5.81868
R406 VOUT.n354 VOUT.n350 5.62509
R407 VOUT.n346 VOUT.n341 5.62509
R408 VOUT.n18 VOUT.n14 5.62509
R409 VOUT.n10 VOUT.n6 5.62509
R410 VOUT.n257 VOUT.n182 5.09533
R411 VOUT.n256 VOUT.n21 5.06947
R412 VOUT.n358 VOUT.n12 5.06539
R413 VOUT.n162 VOUT.n161 5.04292
R414 VOUT.n128 VOUT.n117 5.04292
R415 VOUT.n293 VOUT.n285 5.04292
R416 VOUT.n330 VOUT.n269 5.04292
R417 VOUT.n211 VOUT.n203 5.04292
R418 VOUT.n248 VOUT.n187 5.04292
R419 VOUT.n50 VOUT.n42 5.04292
R420 VOUT.n87 VOUT.n26 5.04292
R421 VOUT.n176 VOUT.n175 4.9683
R422 VOUT.n181 VOUT.n180 4.93989
R423 VOUT.n339 VOUT.n338 4.88412
R424 VOUT.n357 VOUT.n356 4.88412
R425 VIN VOUT.n4 4.83671
R426 VOUT.n359 VOUT.n358 4.5005
R427 VOUT.n261 VOUT.n21 4.5005
R428 VOUT.n158 VOUT.n100 4.26717
R429 VOUT.n129 VOUT.n115 4.26717
R430 VOUT.n297 VOUT.n296 4.26717
R431 VOUT.n327 VOUT.n326 4.26717
R432 VOUT.n215 VOUT.n214 4.26717
R433 VOUT.n245 VOUT.n244 4.26717
R434 VOUT.n54 VOUT.n53 4.26717
R435 VOUT.n84 VOUT.n83 4.26717
R436 VOUT.n157 VOUT.n102 3.49141
R437 VOUT.n133 VOUT.n132 3.49141
R438 VOUT.n300 VOUT.n283 3.49141
R439 VOUT.n323 VOUT.n271 3.49141
R440 VOUT.n218 VOUT.n201 3.49141
R441 VOUT.n241 VOUT.n189 3.49141
R442 VOUT.n57 VOUT.n40 3.49141
R443 VOUT.n80 VOUT.n28 3.49141
R444 VOUT.n154 VOUT.n153 2.71565
R445 VOUT.n136 VOUT.n113 2.71565
R446 VOUT.n301 VOUT.n281 2.71565
R447 VOUT.n322 VOUT.n273 2.71565
R448 VOUT.n219 VOUT.n199 2.71565
R449 VOUT.n240 VOUT.n191 2.71565
R450 VOUT.n58 VOUT.n38 2.71565
R451 VOUT.n79 VOUT.n30 2.71565
R452 VOUT.n259 VOUT.t18 2.41903
R453 VOUT.n259 VOUT.t1 2.41903
R454 VOUT.n264 VOUT.t20 2.41903
R455 VOUT.n264 VOUT.t4 2.41903
R456 VOUT.n258 VOUT.t14 2.41903
R457 VOUT.t18 VOUT.n258 2.41903
R458 VOUT.t4 VOUT.n263 2.41903
R459 VOUT.n263 VOUT.t11 2.41903
R460 VOUT.n164 VOUT.n96 2.41282
R461 VOUT.n288 VOUT.n286 2.41282
R462 VOUT.n206 VOUT.n204 2.41282
R463 VOUT.n45 VOUT.n43 2.41282
R464 VOUT.n150 VOUT.n104 1.93989
R465 VOUT.n137 VOUT.n111 1.93989
R466 VOUT.n306 VOUT.n304 1.93989
R467 VOUT.n319 VOUT.n318 1.93989
R468 VOUT.n224 VOUT.n222 1.93989
R469 VOUT.n237 VOUT.n236 1.93989
R470 VOUT.n63 VOUT.n61 1.93989
R471 VOUT.n76 VOUT.n75 1.93989
R472 VOUT.n357 VOUT.n339 1.68608
R473 VOUT.n149 VOUT.n106 1.16414
R474 VOUT.n141 VOUT.n140 1.16414
R475 VOUT.n305 VOUT.n279 1.16414
R476 VOUT.n315 VOUT.n275 1.16414
R477 VOUT.n355 VOUT.n349 1.16414
R478 VOUT.n343 VOUT.n342 1.16414
R479 VOUT.n19 VOUT.n13 1.16414
R480 VOUT.n11 VOUT.n5 1.16414
R481 VOUT.n223 VOUT.n197 1.16414
R482 VOUT.n233 VOUT.n193 1.16414
R483 VOUT.n62 VOUT.n36 1.16414
R484 VOUT.n72 VOUT.n32 1.16414
R485 VOUT.n358 VOUT.n357 1.11094
R486 VOUT.n360 VOUT.n359 0.595328
R487 VOUT.n363 VOUT.n12 0.509121
R488 VOUT.n257 VOUT.n256 0.466017
R489 VOUT.n146 VOUT.n145 0.388379
R490 VOUT.n110 VOUT.n108 0.388379
R491 VOUT.n311 VOUT.n310 0.388379
R492 VOUT.n314 VOUT.n277 0.388379
R493 VOUT.n353 VOUT.n352 0.388379
R494 VOUT.n345 VOUT.n344 0.388379
R495 VOUT.n17 VOUT.n16 0.388379
R496 VOUT.n9 VOUT.n8 0.388379
R497 VOUT.n229 VOUT.n228 0.388379
R498 VOUT.n232 VOUT.n195 0.388379
R499 VOUT.n68 VOUT.n67 0.388379
R500 VOUT.n71 VOUT.n34 0.388379
R501 VOUT VOUT.n260 0.353948
R502 VOUT.n176 VOUT.n4 0.282952
R503 VOUT.n261 VOUT 0.263431
R504 VIN VOUT.n363 0.259121
R505 VOUT.n182 VOUT.n181 0.258175
R506 VOUT.n164 VOUT.n163 0.155672
R507 VOUT.n163 VOUT.n99 0.155672
R508 VOUT.n156 VOUT.n99 0.155672
R509 VOUT.n156 VOUT.n155 0.155672
R510 VOUT.n155 VOUT.n103 0.155672
R511 VOUT.n148 VOUT.n103 0.155672
R512 VOUT.n148 VOUT.n147 0.155672
R513 VOUT.n147 VOUT.n107 0.155672
R514 VOUT.n139 VOUT.n107 0.155672
R515 VOUT.n139 VOUT.n138 0.155672
R516 VOUT.n138 VOUT.n112 0.155672
R517 VOUT.n131 VOUT.n112 0.155672
R518 VOUT.n131 VOUT.n130 0.155672
R519 VOUT.n130 VOUT.n116 0.155672
R520 VOUT.n123 VOUT.n116 0.155672
R521 VOUT.n123 VOUT.n122 0.155672
R522 VOUT.n294 VOUT.n286 0.155672
R523 VOUT.n295 VOUT.n294 0.155672
R524 VOUT.n295 VOUT.n282 0.155672
R525 VOUT.n302 VOUT.n282 0.155672
R526 VOUT.n303 VOUT.n302 0.155672
R527 VOUT.n303 VOUT.n278 0.155672
R528 VOUT.n312 VOUT.n278 0.155672
R529 VOUT.n313 VOUT.n312 0.155672
R530 VOUT.n313 VOUT.n274 0.155672
R531 VOUT.n320 VOUT.n274 0.155672
R532 VOUT.n321 VOUT.n320 0.155672
R533 VOUT.n321 VOUT.n270 0.155672
R534 VOUT.n328 VOUT.n270 0.155672
R535 VOUT.n329 VOUT.n328 0.155672
R536 VOUT.n329 VOUT.n266 0.155672
R537 VOUT.n336 VOUT.n266 0.155672
R538 VOUT.n212 VOUT.n204 0.155672
R539 VOUT.n213 VOUT.n212 0.155672
R540 VOUT.n213 VOUT.n200 0.155672
R541 VOUT.n220 VOUT.n200 0.155672
R542 VOUT.n221 VOUT.n220 0.155672
R543 VOUT.n221 VOUT.n196 0.155672
R544 VOUT.n230 VOUT.n196 0.155672
R545 VOUT.n231 VOUT.n230 0.155672
R546 VOUT.n231 VOUT.n192 0.155672
R547 VOUT.n238 VOUT.n192 0.155672
R548 VOUT.n239 VOUT.n238 0.155672
R549 VOUT.n239 VOUT.n188 0.155672
R550 VOUT.n246 VOUT.n188 0.155672
R551 VOUT.n247 VOUT.n246 0.155672
R552 VOUT.n247 VOUT.n184 0.155672
R553 VOUT.n254 VOUT.n184 0.155672
R554 VOUT.n51 VOUT.n43 0.155672
R555 VOUT.n52 VOUT.n51 0.155672
R556 VOUT.n52 VOUT.n39 0.155672
R557 VOUT.n59 VOUT.n39 0.155672
R558 VOUT.n60 VOUT.n59 0.155672
R559 VOUT.n60 VOUT.n35 0.155672
R560 VOUT.n69 VOUT.n35 0.155672
R561 VOUT.n70 VOUT.n69 0.155672
R562 VOUT.n70 VOUT.n31 0.155672
R563 VOUT.n77 VOUT.n31 0.155672
R564 VOUT.n78 VOUT.n77 0.155672
R565 VOUT.n78 VOUT.n27 0.155672
R566 VOUT.n85 VOUT.n27 0.155672
R567 VOUT.n86 VOUT.n85 0.155672
R568 VOUT.n86 VOUT.n23 0.155672
R569 VOUT.n93 VOUT.n23 0.155672
R570 VGN VOUT.n3 0.127394
R571 VGP VOUT.n171 0.0989849
R572 VSS.n121 VSS.n50 586.196
R573 VSS.n72 VSS.n48 586.196
R574 VSS.n213 VSS.n25 586.196
R575 VSS.n216 VSS.n10 586.196
R576 VSS.n51 VSS.n50 585
R577 VSS.n50 VSS.n49 585
R578 VSS.n126 VSS.n125 585
R579 VSS.n127 VSS.n126 585
R580 VSS.n42 VSS.n41 585
R581 VSS.n43 VSS.n42 585
R582 VSS.n139 VSS.n138 585
R583 VSS.n138 VSS.n137 585
R584 VSS.n39 VSS.n38 585
R585 VSS.n136 VSS.n38 585
R586 VSS.n144 VSS.n143 585
R587 VSS.n145 VSS.n144 585
R588 VSS.n36 VSS.n35 585
R589 VSS.n146 VSS.n36 585
R590 VSS.n149 VSS.n148 585
R591 VSS.n148 VSS.n147 585
R592 VSS.n33 VSS.n32 585
R593 VSS.n32 VSS.n30 585
R594 VSS.n155 VSS.n154 585
R595 VSS.n156 VSS.n155 585
R596 VSS.n29 VSS.n28 585
R597 VSS.n157 VSS.n29 585
R598 VSS.n160 VSS.n159 585
R599 VSS.n159 VSS.n158 585
R600 VSS.n161 VSS.n25 585
R601 VSS.n25 VSS.n13 585
R602 VSS.n219 VSS.n10 585
R603 VSS.n13 VSS.n10 585
R604 VSS.n220 VSS.n9 585
R605 VSS.n158 VSS.n9 585
R606 VSS.n221 VSS.n8 585
R607 VSS.n157 VSS.n8 585
R608 VSS.n31 VSS.n6 585
R609 VSS.n156 VSS.n31 585
R610 VSS.n225 VSS.n5 585
R611 VSS.n30 VSS.n5 585
R612 VSS.n226 VSS.n4 585
R613 VSS.n147 VSS.n4 585
R614 VSS.n227 VSS.n3 585
R615 VSS.n146 VSS.n3 585
R616 VSS.n37 VSS.n2 585
R617 VSS.n145 VSS.n37 585
R618 VSS.n135 VSS.n134 585
R619 VSS.n136 VSS.n135 585
R620 VSS.n45 VSS.n44 585
R621 VSS.n137 VSS.n44 585
R622 VSS.n130 VSS.n129 585
R623 VSS.n129 VSS.n43 585
R624 VSS.n128 VSS.n47 585
R625 VSS.n128 VSS.n127 585
R626 VSS.n70 VSS.n48 585
R627 VSS.n49 VSS.n48 585
R628 VSS.n217 VSS.n216 585
R629 VSS.n12 VSS.n11 585
R630 VSS.n168 VSS.n167 585
R631 VSS.n171 VSS.n170 585
R632 VSS.n173 VSS.n172 585
R633 VSS.n175 VSS.n174 585
R634 VSS.n177 VSS.n176 585
R635 VSS.n179 VSS.n178 585
R636 VSS.n181 VSS.n180 585
R637 VSS.n183 VSS.n182 585
R638 VSS.n185 VSS.n184 585
R639 VSS.n187 VSS.n186 585
R640 VSS.n189 VSS.n188 585
R641 VSS.n191 VSS.n190 585
R642 VSS.n193 VSS.n192 585
R643 VSS.n196 VSS.n195 585
R644 VSS.n198 VSS.n197 585
R645 VSS.n200 VSS.n199 585
R646 VSS.n202 VSS.n201 585
R647 VSS.n204 VSS.n203 585
R648 VSS.n206 VSS.n205 585
R649 VSS.n208 VSS.n207 585
R650 VSS.n210 VSS.n209 585
R651 VSS.n211 VSS.n26 585
R652 VSS.n213 VSS.n212 585
R653 VSS.n214 VSS.n213 585
R654 VSS.n122 VSS.n121 585
R655 VSS.n53 VSS.n52 585
R656 VSS.n118 VSS.n117 585
R657 VSS.n119 VSS.n118 585
R658 VSS.n116 VSS.n65 585
R659 VSS.n115 VSS.n114 585
R660 VSS.n113 VSS.n112 585
R661 VSS.n111 VSS.n110 585
R662 VSS.n109 VSS.n108 585
R663 VSS.n107 VSS.n106 585
R664 VSS.n105 VSS.n104 585
R665 VSS.n102 VSS.n101 585
R666 VSS.n100 VSS.n99 585
R667 VSS.n98 VSS.n97 585
R668 VSS.n96 VSS.n95 585
R669 VSS.n94 VSS.n93 585
R670 VSS.n92 VSS.n91 585
R671 VSS.n90 VSS.n89 585
R672 VSS.n88 VSS.n87 585
R673 VSS.n86 VSS.n85 585
R674 VSS.n84 VSS.n83 585
R675 VSS.n82 VSS.n81 585
R676 VSS.n80 VSS.n79 585
R677 VSS.n77 VSS.n76 585
R678 VSS.n75 VSS.n74 585
R679 VSS.n73 VSS.n72 585
R680 VSS.n163 VSS.t7 393
R681 VSS.n165 VSS.t3 393
R682 VSS.n68 VSS.t14 393
R683 VSS.n66 VSS.t10 393
R684 VSS.n119 VSS.n49 342.13
R685 VSS.n214 VSS.n13 342.13
R686 VSS.n215 VSS.n214 256.663
R687 VSS.n214 VSS.n14 256.663
R688 VSS.n214 VSS.n15 256.663
R689 VSS.n214 VSS.n16 256.663
R690 VSS.n214 VSS.n17 256.663
R691 VSS.n214 VSS.n18 256.663
R692 VSS.n214 VSS.n19 256.663
R693 VSS.n214 VSS.n20 256.663
R694 VSS.n214 VSS.n21 256.663
R695 VSS.n214 VSS.n22 256.663
R696 VSS.n214 VSS.n23 256.663
R697 VSS.n214 VSS.n24 256.663
R698 VSS.n120 VSS.n119 256.663
R699 VSS.n119 VSS.n54 256.663
R700 VSS.n119 VSS.n55 256.663
R701 VSS.n119 VSS.n56 256.663
R702 VSS.n119 VSS.n57 256.663
R703 VSS.n119 VSS.n58 256.663
R704 VSS.n119 VSS.n59 256.663
R705 VSS.n119 VSS.n60 256.663
R706 VSS.n119 VSS.n61 256.663
R707 VSS.n119 VSS.n62 256.663
R708 VSS.n119 VSS.n63 256.663
R709 VSS.n119 VSS.n64 256.663
R710 VSS.n126 VSS.n50 240.244
R711 VSS.n126 VSS.n42 240.244
R712 VSS.n138 VSS.n42 240.244
R713 VSS.n138 VSS.n38 240.244
R714 VSS.n144 VSS.n38 240.244
R715 VSS.n144 VSS.n36 240.244
R716 VSS.n148 VSS.n36 240.244
R717 VSS.n148 VSS.n32 240.244
R718 VSS.n155 VSS.n32 240.244
R719 VSS.n155 VSS.n29 240.244
R720 VSS.n159 VSS.n29 240.244
R721 VSS.n159 VSS.n25 240.244
R722 VSS.n128 VSS.n48 240.244
R723 VSS.n129 VSS.n128 240.244
R724 VSS.n129 VSS.n44 240.244
R725 VSS.n135 VSS.n44 240.244
R726 VSS.n135 VSS.n37 240.244
R727 VSS.n37 VSS.n3 240.244
R728 VSS.n4 VSS.n3 240.244
R729 VSS.n5 VSS.n4 240.244
R730 VSS.n31 VSS.n5 240.244
R731 VSS.n31 VSS.n8 240.244
R732 VSS.n9 VSS.n8 240.244
R733 VSS.n10 VSS.n9 240.244
R734 VSS.n127 VSS.n49 207.352
R735 VSS.n137 VSS.n43 207.352
R736 VSS.n137 VSS.n136 207.352
R737 VSS.n147 VSS.n30 207.352
R738 VSS.n156 VSS.n30 207.352
R739 VSS.n157 VSS.n156 207.352
R740 VSS.n158 VSS.n13 207.352
R741 VSS.t11 VSS.n43 182.47
R742 VSS.t1 VSS.n146 174.175
R743 VSS.n158 VSS.t4 165.881
R744 VSS.n118 VSS.n53 163.367
R745 VSS.n118 VSS.n65 163.367
R746 VSS.n114 VSS.n113 163.367
R747 VSS.n110 VSS.n109 163.367
R748 VSS.n106 VSS.n105 163.367
R749 VSS.n101 VSS.n100 163.367
R750 VSS.n97 VSS.n96 163.367
R751 VSS.n93 VSS.n92 163.367
R752 VSS.n89 VSS.n88 163.367
R753 VSS.n85 VSS.n84 163.367
R754 VSS.n81 VSS.n80 163.367
R755 VSS.n76 VSS.n75 163.367
R756 VSS.n213 VSS.n26 163.367
R757 VSS.n209 VSS.n208 163.367
R758 VSS.n205 VSS.n204 163.367
R759 VSS.n201 VSS.n200 163.367
R760 VSS.n197 VSS.n196 163.367
R761 VSS.n192 VSS.n191 163.367
R762 VSS.n188 VSS.n187 163.367
R763 VSS.n184 VSS.n183 163.367
R764 VSS.n180 VSS.n179 163.367
R765 VSS.n176 VSS.n175 163.367
R766 VSS.n172 VSS.n171 163.367
R767 VSS.n167 VSS.n12 163.367
R768 VSS.t0 VSS.n145 136.852
R769 VSS.n163 VSS.t8 131.357
R770 VSS.n165 VSS.t5 131.357
R771 VSS.n68 VSS.t16 131.357
R772 VSS.n66 VSS.t13 131.357
R773 VSS.n164 VSS.t9 119.915
R774 VSS.n166 VSS.t6 119.915
R775 VSS.n69 VSS.t15 119.915
R776 VSS.n67 VSS.t12 119.915
R777 VSS.n145 VSS.t2 107.823
R778 VSS.n136 VSS.t2 99.5292
R779 VSS.n121 VSS.n120 71.676
R780 VSS.n65 VSS.n54 71.676
R781 VSS.n113 VSS.n55 71.676
R782 VSS.n109 VSS.n56 71.676
R783 VSS.n105 VSS.n57 71.676
R784 VSS.n100 VSS.n58 71.676
R785 VSS.n96 VSS.n59 71.676
R786 VSS.n92 VSS.n60 71.676
R787 VSS.n88 VSS.n61 71.676
R788 VSS.n84 VSS.n62 71.676
R789 VSS.n80 VSS.n63 71.676
R790 VSS.n75 VSS.n64 71.676
R791 VSS.n209 VSS.n24 71.676
R792 VSS.n205 VSS.n23 71.676
R793 VSS.n201 VSS.n22 71.676
R794 VSS.n197 VSS.n21 71.676
R795 VSS.n192 VSS.n20 71.676
R796 VSS.n188 VSS.n19 71.676
R797 VSS.n184 VSS.n18 71.676
R798 VSS.n180 VSS.n17 71.676
R799 VSS.n176 VSS.n16 71.676
R800 VSS.n172 VSS.n15 71.676
R801 VSS.n167 VSS.n14 71.676
R802 VSS.n216 VSS.n215 71.676
R803 VSS.n215 VSS.n12 71.676
R804 VSS.n171 VSS.n14 71.676
R805 VSS.n175 VSS.n15 71.676
R806 VSS.n179 VSS.n16 71.676
R807 VSS.n183 VSS.n17 71.676
R808 VSS.n187 VSS.n18 71.676
R809 VSS.n191 VSS.n19 71.676
R810 VSS.n196 VSS.n20 71.676
R811 VSS.n200 VSS.n21 71.676
R812 VSS.n204 VSS.n22 71.676
R813 VSS.n208 VSS.n23 71.676
R814 VSS.n26 VSS.n24 71.676
R815 VSS.n120 VSS.n53 71.676
R816 VSS.n114 VSS.n54 71.676
R817 VSS.n110 VSS.n55 71.676
R818 VSS.n106 VSS.n56 71.676
R819 VSS.n101 VSS.n57 71.676
R820 VSS.n97 VSS.n58 71.676
R821 VSS.n93 VSS.n59 71.676
R822 VSS.n89 VSS.n60 71.676
R823 VSS.n85 VSS.n61 71.676
R824 VSS.n81 VSS.n62 71.676
R825 VSS.n76 VSS.n63 71.676
R826 VSS.n72 VSS.n64 71.676
R827 VSS.n146 VSS.t0 70.5
R828 VSS.n194 VSS.n164 47.5157
R829 VSS.n169 VSS.n166 47.5157
R830 VSS.t4 VSS.n157 41.4708
R831 VSS.n78 VSS.n69 34.3278
R832 VSS.n103 VSS.n67 34.3278
R833 VSS.n147 VSS.t1 33.1768
R834 VSS.n212 VSS.n162 28.2837
R835 VSS.n218 VSS.n217 28.2837
R836 VSS.n123 VSS.n122 28.2837
R837 VSS.n73 VSS.n71 28.2837
R838 VSS.n127 VSS.t11 24.8827
R839 VSS.n125 VSS.n51 19.3944
R840 VSS.n125 VSS.n41 19.3944
R841 VSS.n139 VSS.n41 19.3944
R842 VSS.n139 VSS.n39 19.3944
R843 VSS.n143 VSS.n39 19.3944
R844 VSS.n143 VSS.n35 19.3944
R845 VSS.n149 VSS.n35 19.3944
R846 VSS.n149 VSS.n33 19.3944
R847 VSS.n154 VSS.n33 19.3944
R848 VSS.n154 VSS.n28 19.3944
R849 VSS.n160 VSS.n28 19.3944
R850 VSS.n161 VSS.n160 19.3944
R851 VSS.n70 VSS.n47 19.3944
R852 VSS.n130 VSS.n47 19.3944
R853 VSS.n130 VSS.n45 19.3944
R854 VSS.n134 VSS.n45 19.3944
R855 VSS.n134 VSS.n2 19.3944
R856 VSS.n227 VSS.n2 19.3944
R857 VSS.n227 VSS.n226 19.3944
R858 VSS.n226 VSS.n225 19.3944
R859 VSS.n225 VSS.n6 19.3944
R860 VSS.n221 VSS.n6 19.3944
R861 VSS.n221 VSS.n220 19.3944
R862 VSS.n220 VSS.n219 19.3944
R863 VSS.n164 VSS.n163 11.4429
R864 VSS.n166 VSS.n165 11.4429
R865 VSS.n69 VSS.n68 11.4429
R866 VSS.n67 VSS.n66 11.4429
R867 VSS.n212 VSS.n211 10.6151
R868 VSS.n211 VSS.n210 10.6151
R869 VSS.n210 VSS.n207 10.6151
R870 VSS.n207 VSS.n206 10.6151
R871 VSS.n206 VSS.n203 10.6151
R872 VSS.n203 VSS.n202 10.6151
R873 VSS.n202 VSS.n199 10.6151
R874 VSS.n199 VSS.n198 10.6151
R875 VSS.n198 VSS.n195 10.6151
R876 VSS.n193 VSS.n190 10.6151
R877 VSS.n190 VSS.n189 10.6151
R878 VSS.n189 VSS.n186 10.6151
R879 VSS.n186 VSS.n185 10.6151
R880 VSS.n185 VSS.n182 10.6151
R881 VSS.n182 VSS.n181 10.6151
R882 VSS.n181 VSS.n178 10.6151
R883 VSS.n178 VSS.n177 10.6151
R884 VSS.n177 VSS.n174 10.6151
R885 VSS.n174 VSS.n173 10.6151
R886 VSS.n173 VSS.n170 10.6151
R887 VSS.n168 VSS.n11 10.6151
R888 VSS.n217 VSS.n11 10.6151
R889 VSS.n122 VSS.n52 10.6151
R890 VSS.n117 VSS.n52 10.6151
R891 VSS.n117 VSS.n116 10.6151
R892 VSS.n116 VSS.n115 10.6151
R893 VSS.n115 VSS.n112 10.6151
R894 VSS.n112 VSS.n111 10.6151
R895 VSS.n111 VSS.n108 10.6151
R896 VSS.n108 VSS.n107 10.6151
R897 VSS.n107 VSS.n104 10.6151
R898 VSS.n102 VSS.n99 10.6151
R899 VSS.n99 VSS.n98 10.6151
R900 VSS.n98 VSS.n95 10.6151
R901 VSS.n95 VSS.n94 10.6151
R902 VSS.n94 VSS.n91 10.6151
R903 VSS.n91 VSS.n90 10.6151
R904 VSS.n90 VSS.n87 10.6151
R905 VSS.n87 VSS.n86 10.6151
R906 VSS.n86 VSS.n83 10.6151
R907 VSS.n83 VSS.n82 10.6151
R908 VSS.n82 VSS.n79 10.6151
R909 VSS.n77 VSS.n74 10.6151
R910 VSS.n74 VSS.n73 10.6151
R911 VSS.n226 VSS.n0 9.3005
R912 VSS.n225 VSS.n224 9.3005
R913 VSS.n223 VSS.n6 9.3005
R914 VSS.n222 VSS.n221 9.3005
R915 VSS.n220 VSS.n7 9.3005
R916 VSS.n219 VSS.n218 9.3005
R917 VSS.n123 VSS.n51 9.3005
R918 VSS.n125 VSS.n124 9.3005
R919 VSS.n41 VSS.n40 9.3005
R920 VSS.n140 VSS.n139 9.3005
R921 VSS.n141 VSS.n39 9.3005
R922 VSS.n143 VSS.n142 9.3005
R923 VSS.n35 VSS.n34 9.3005
R924 VSS.n150 VSS.n149 9.3005
R925 VSS.n151 VSS.n33 9.3005
R926 VSS.n154 VSS.n153 9.3005
R927 VSS.n152 VSS.n28 9.3005
R928 VSS.n160 VSS.n27 9.3005
R929 VSS.n162 VSS.n161 9.3005
R930 VSS.n47 VSS.n46 9.3005
R931 VSS.n131 VSS.n130 9.3005
R932 VSS.n132 VSS.n45 9.3005
R933 VSS.n134 VSS.n133 9.3005
R934 VSS.n2 VSS.n1 9.3005
R935 VSS.n71 VSS.n70 9.3005
R936 VSS.n228 VSS.n227 9.3005
R937 VSS.n170 VSS.n169 6.7127
R938 VSS.n79 VSS.n78 6.7127
R939 VSS.n195 VSS.n194 6.0883
R940 VSS.n104 VSS.n103 6.0883
R941 VSS.n194 VSS.n193 4.52733
R942 VSS.n103 VSS.n102 4.52733
R943 VSS.n169 VSS.n168 3.90294
R944 VSS.n78 VSS.n77 3.90294
R945 VSS.n224 VSS.n0 0.152939
R946 VSS.n224 VSS.n223 0.152939
R947 VSS.n223 VSS.n222 0.152939
R948 VSS.n222 VSS.n7 0.152939
R949 VSS.n218 VSS.n7 0.152939
R950 VSS.n124 VSS.n123 0.152939
R951 VSS.n124 VSS.n40 0.152939
R952 VSS.n140 VSS.n40 0.152939
R953 VSS.n141 VSS.n140 0.152939
R954 VSS.n142 VSS.n141 0.152939
R955 VSS.n142 VSS.n34 0.152939
R956 VSS.n150 VSS.n34 0.152939
R957 VSS.n151 VSS.n150 0.152939
R958 VSS.n153 VSS.n151 0.152939
R959 VSS.n153 VSS.n152 0.152939
R960 VSS.n152 VSS.n27 0.152939
R961 VSS.n162 VSS.n27 0.152939
R962 VSS.n71 VSS.n46 0.152939
R963 VSS.n131 VSS.n46 0.152939
R964 VSS.n132 VSS.n131 0.152939
R965 VSS.n133 VSS.n132 0.152939
R966 VSS.n133 VSS.n1 0.152939
R967 VSS.n228 VSS.n1 0.13922
R968 VSS VSS.n0 0.0767195
R969 VSS VSS.n228 0.063
R970 VCC.n355 VCC.t14 1775.88
R971 VCC.n331 VCC.t7 1775.88
R972 VCC.n88 VCC.t11 1775.88
R973 VCC.n85 VCC.t3 1775.88
R974 VCC.n355 VCC.t15 412.048
R975 VCC.n331 VCC.t9 412.048
R976 VCC.n88 VCC.t13 412.048
R977 VCC.n85 VCC.t6 412.048
R978 VCC.n356 VCC.t16 401.575
R979 VCC.n332 VCC.t10 401.575
R980 VCC.n89 VCC.t12 401.575
R981 VCC.n86 VCC.t5 401.575
R982 VCC.n547 VCC.n9 386.341
R983 VCC.n545 VCC.n13 386.341
R984 VCC.n82 VCC.n31 386.341
R985 VCC.n271 VCC.n32 386.341
R986 VCC.n545 VCC.n544 185
R987 VCC.n546 VCC.n545 185
R988 VCC.n14 VCC.n12 185
R989 VCC.n12 VCC.n10 185
R990 VCC.n306 VCC.n305 185
R991 VCC.n305 VCC.n304 185
R992 VCC.n17 VCC.n16 185
R993 VCC.n302 VCC.n17 185
R994 VCC.n300 VCC.n299 185
R995 VCC.n301 VCC.n300 185
R996 VCC.n19 VCC.n18 185
R997 VCC.n23 VCC.n18 185
R998 VCC.n295 VCC.n294 185
R999 VCC.n294 VCC.n293 185
R1000 VCC.n22 VCC.n21 185
R1001 VCC.n290 VCC.n22 185
R1002 VCC.n288 VCC.n287 185
R1003 VCC.n289 VCC.n288 185
R1004 VCC.n28 VCC.n27 185
R1005 VCC.n27 VCC.n26 185
R1006 VCC.n283 VCC.n282 185
R1007 VCC.n282 VCC.n281 185
R1008 VCC.n31 VCC.n30 185
R1009 VCC.n83 VCC.n31 185
R1010 VCC.n34 VCC.n32 185
R1011 VCC.n83 VCC.n32 185
R1012 VCC.n280 VCC.n279 185
R1013 VCC.n281 VCC.n280 185
R1014 VCC.n35 VCC.n33 185
R1015 VCC.n33 VCC.n26 185
R1016 VCC.n275 VCC.n24 185
R1017 VCC.n289 VCC.n24 185
R1018 VCC.n291 VCC.n25 185
R1019 VCC.n291 VCC.n290 185
R1020 VCC.n292 VCC.n2 185
R1021 VCC.n293 VCC.n292 185
R1022 VCC.n555 VCC.n3 185
R1023 VCC.n23 VCC.n3 185
R1024 VCC.n554 VCC.n4 185
R1025 VCC.n301 VCC.n4 185
R1026 VCC.n553 VCC.n5 185
R1027 VCC.n302 VCC.n5 185
R1028 VCC.n303 VCC.n6 185
R1029 VCC.n304 VCC.n303 185
R1030 VCC.n549 VCC.n8 185
R1031 VCC.n10 VCC.n8 185
R1032 VCC.n548 VCC.n547 185
R1033 VCC.n547 VCC.n546 185
R1034 VCC.n542 VCC.n13 185
R1035 VCC.n541 VCC.n540 185
R1036 VCC.n538 VCC.n309 185
R1037 VCC.n536 VCC.n535 185
R1038 VCC.n534 VCC.n310 185
R1039 VCC.n533 VCC.n532 185
R1040 VCC.n530 VCC.n311 185
R1041 VCC.n528 VCC.n527 185
R1042 VCC.n526 VCC.n312 185
R1043 VCC.n525 VCC.n524 185
R1044 VCC.n522 VCC.n313 185
R1045 VCC.n520 VCC.n519 185
R1046 VCC.n518 VCC.n314 185
R1047 VCC.n517 VCC.n516 185
R1048 VCC.n514 VCC.n315 185
R1049 VCC.n512 VCC.n511 185
R1050 VCC.n510 VCC.n316 185
R1051 VCC.n509 VCC.n508 185
R1052 VCC.n506 VCC.n317 185
R1053 VCC.n504 VCC.n503 185
R1054 VCC.n502 VCC.n318 185
R1055 VCC.n501 VCC.n500 185
R1056 VCC.n498 VCC.n319 185
R1057 VCC.n496 VCC.n495 185
R1058 VCC.n494 VCC.n320 185
R1059 VCC.n493 VCC.n492 185
R1060 VCC.n490 VCC.n321 185
R1061 VCC.n488 VCC.n487 185
R1062 VCC.n486 VCC.n322 185
R1063 VCC.n485 VCC.n484 185
R1064 VCC.n482 VCC.n323 185
R1065 VCC.n480 VCC.n479 185
R1066 VCC.n478 VCC.n324 185
R1067 VCC.n477 VCC.n476 185
R1068 VCC.n474 VCC.n325 185
R1069 VCC.n472 VCC.n471 185
R1070 VCC.n470 VCC.n326 185
R1071 VCC.n469 VCC.n468 185
R1072 VCC.n466 VCC.n327 185
R1073 VCC.n464 VCC.n463 185
R1074 VCC.n462 VCC.n328 185
R1075 VCC.n461 VCC.n460 185
R1076 VCC.n458 VCC.n329 185
R1077 VCC.n456 VCC.n455 185
R1078 VCC.n453 VCC.n330 185
R1079 VCC.n452 VCC.n451 185
R1080 VCC.n449 VCC.n333 185
R1081 VCC.n447 VCC.n446 185
R1082 VCC.n445 VCC.n334 185
R1083 VCC.n444 VCC.n443 185
R1084 VCC.n441 VCC.n335 185
R1085 VCC.n439 VCC.n438 185
R1086 VCC.n437 VCC.n336 185
R1087 VCC.n436 VCC.n435 185
R1088 VCC.n433 VCC.n337 185
R1089 VCC.n431 VCC.n430 185
R1090 VCC.n429 VCC.n338 185
R1091 VCC.n428 VCC.n427 185
R1092 VCC.n425 VCC.n339 185
R1093 VCC.n423 VCC.n422 185
R1094 VCC.n421 VCC.n340 185
R1095 VCC.n420 VCC.n419 185
R1096 VCC.n417 VCC.n341 185
R1097 VCC.n415 VCC.n414 185
R1098 VCC.n413 VCC.n342 185
R1099 VCC.n412 VCC.n411 185
R1100 VCC.n409 VCC.n343 185
R1101 VCC.n407 VCC.n406 185
R1102 VCC.n405 VCC.n344 185
R1103 VCC.n404 VCC.n403 185
R1104 VCC.n401 VCC.n345 185
R1105 VCC.n399 VCC.n398 185
R1106 VCC.n397 VCC.n346 185
R1107 VCC.n396 VCC.n395 185
R1108 VCC.n393 VCC.n347 185
R1109 VCC.n391 VCC.n390 185
R1110 VCC.n389 VCC.n348 185
R1111 VCC.n388 VCC.n387 185
R1112 VCC.n385 VCC.n349 185
R1113 VCC.n383 VCC.n382 185
R1114 VCC.n381 VCC.n350 185
R1115 VCC.n380 VCC.n379 185
R1116 VCC.n377 VCC.n351 185
R1117 VCC.n375 VCC.n374 185
R1118 VCC.n373 VCC.n352 185
R1119 VCC.n372 VCC.n371 185
R1120 VCC.n369 VCC.n353 185
R1121 VCC.n367 VCC.n366 185
R1122 VCC.n365 VCC.n354 185
R1123 VCC.n364 VCC.n363 185
R1124 VCC.n361 VCC.n360 185
R1125 VCC.n359 VCC.n9 185
R1126 VCC.n272 VCC.n271 185
R1127 VCC.n37 VCC.n36 185
R1128 VCC.n268 VCC.n267 185
R1129 VCC.n269 VCC.n268 185
R1130 VCC.n266 VCC.n84 185
R1131 VCC.n265 VCC.n264 185
R1132 VCC.n263 VCC.n262 185
R1133 VCC.n261 VCC.n260 185
R1134 VCC.n259 VCC.n258 185
R1135 VCC.n257 VCC.n256 185
R1136 VCC.n255 VCC.n254 185
R1137 VCC.n253 VCC.n252 185
R1138 VCC.n251 VCC.n250 185
R1139 VCC.n249 VCC.n248 185
R1140 VCC.n247 VCC.n246 185
R1141 VCC.n245 VCC.n244 185
R1142 VCC.n243 VCC.n242 185
R1143 VCC.n241 VCC.n240 185
R1144 VCC.n239 VCC.n238 185
R1145 VCC.n237 VCC.n236 185
R1146 VCC.n235 VCC.n234 185
R1147 VCC.n233 VCC.n232 185
R1148 VCC.n231 VCC.n230 185
R1149 VCC.n229 VCC.n228 185
R1150 VCC.n227 VCC.n226 185
R1151 VCC.n225 VCC.n224 185
R1152 VCC.n223 VCC.n222 185
R1153 VCC.n221 VCC.n220 185
R1154 VCC.n219 VCC.n218 185
R1155 VCC.n217 VCC.n216 185
R1156 VCC.n215 VCC.n214 185
R1157 VCC.n213 VCC.n212 185
R1158 VCC.n211 VCC.n210 185
R1159 VCC.n209 VCC.n208 185
R1160 VCC.n207 VCC.n206 185
R1161 VCC.n205 VCC.n204 185
R1162 VCC.n203 VCC.n202 185
R1163 VCC.n201 VCC.n200 185
R1164 VCC.n199 VCC.n198 185
R1165 VCC.n197 VCC.n196 185
R1166 VCC.n195 VCC.n194 185
R1167 VCC.n193 VCC.n192 185
R1168 VCC.n191 VCC.n190 185
R1169 VCC.n189 VCC.n188 185
R1170 VCC.n187 VCC.n186 185
R1171 VCC.n185 VCC.n184 185
R1172 VCC.n183 VCC.n182 185
R1173 VCC.n181 VCC.n180 185
R1174 VCC.n179 VCC.n178 185
R1175 VCC.n176 VCC.n175 185
R1176 VCC.n174 VCC.n173 185
R1177 VCC.n172 VCC.n171 185
R1178 VCC.n170 VCC.n169 185
R1179 VCC.n168 VCC.n167 185
R1180 VCC.n166 VCC.n165 185
R1181 VCC.n164 VCC.n163 185
R1182 VCC.n162 VCC.n161 185
R1183 VCC.n160 VCC.n159 185
R1184 VCC.n158 VCC.n157 185
R1185 VCC.n156 VCC.n155 185
R1186 VCC.n154 VCC.n153 185
R1187 VCC.n152 VCC.n151 185
R1188 VCC.n150 VCC.n149 185
R1189 VCC.n148 VCC.n147 185
R1190 VCC.n146 VCC.n145 185
R1191 VCC.n144 VCC.n143 185
R1192 VCC.n142 VCC.n141 185
R1193 VCC.n140 VCC.n139 185
R1194 VCC.n138 VCC.n137 185
R1195 VCC.n136 VCC.n135 185
R1196 VCC.n134 VCC.n133 185
R1197 VCC.n132 VCC.n131 185
R1198 VCC.n130 VCC.n129 185
R1199 VCC.n128 VCC.n127 185
R1200 VCC.n126 VCC.n125 185
R1201 VCC.n124 VCC.n123 185
R1202 VCC.n122 VCC.n121 185
R1203 VCC.n120 VCC.n119 185
R1204 VCC.n118 VCC.n117 185
R1205 VCC.n116 VCC.n115 185
R1206 VCC.n114 VCC.n113 185
R1207 VCC.n112 VCC.n111 185
R1208 VCC.n110 VCC.n109 185
R1209 VCC.n108 VCC.n107 185
R1210 VCC.n106 VCC.n105 185
R1211 VCC.n104 VCC.n103 185
R1212 VCC.n102 VCC.n101 185
R1213 VCC.n100 VCC.n99 185
R1214 VCC.n98 VCC.n97 185
R1215 VCC.n96 VCC.n95 185
R1216 VCC.n94 VCC.n93 185
R1217 VCC.n92 VCC.n91 185
R1218 VCC.n90 VCC.n82 185
R1219 VCC.n269 VCC.n82 185
R1220 VCC.n282 VCC.n31 146.341
R1221 VCC.n282 VCC.n27 146.341
R1222 VCC.n288 VCC.n27 146.341
R1223 VCC.n288 VCC.n22 146.341
R1224 VCC.n294 VCC.n22 146.341
R1225 VCC.n294 VCC.n18 146.341
R1226 VCC.n300 VCC.n18 146.341
R1227 VCC.n300 VCC.n17 146.341
R1228 VCC.n305 VCC.n17 146.341
R1229 VCC.n305 VCC.n12 146.341
R1230 VCC.n545 VCC.n12 146.341
R1231 VCC.n280 VCC.n32 146.341
R1232 VCC.n280 VCC.n33 146.341
R1233 VCC.n33 VCC.n24 146.341
R1234 VCC.n291 VCC.n24 146.341
R1235 VCC.n292 VCC.n291 146.341
R1236 VCC.n292 VCC.n3 146.341
R1237 VCC.n4 VCC.n3 146.341
R1238 VCC.n5 VCC.n4 146.341
R1239 VCC.n303 VCC.n5 146.341
R1240 VCC.n303 VCC.n8 146.341
R1241 VCC.n547 VCC.n8 146.341
R1242 VCC.n363 VCC.n361 99.5127
R1243 VCC.n367 VCC.n354 99.5127
R1244 VCC.n371 VCC.n369 99.5127
R1245 VCC.n375 VCC.n352 99.5127
R1246 VCC.n379 VCC.n377 99.5127
R1247 VCC.n383 VCC.n350 99.5127
R1248 VCC.n387 VCC.n385 99.5127
R1249 VCC.n391 VCC.n348 99.5127
R1250 VCC.n395 VCC.n393 99.5127
R1251 VCC.n399 VCC.n346 99.5127
R1252 VCC.n403 VCC.n401 99.5127
R1253 VCC.n407 VCC.n344 99.5127
R1254 VCC.n411 VCC.n409 99.5127
R1255 VCC.n415 VCC.n342 99.5127
R1256 VCC.n419 VCC.n417 99.5127
R1257 VCC.n423 VCC.n340 99.5127
R1258 VCC.n427 VCC.n425 99.5127
R1259 VCC.n431 VCC.n338 99.5127
R1260 VCC.n435 VCC.n433 99.5127
R1261 VCC.n439 VCC.n336 99.5127
R1262 VCC.n443 VCC.n441 99.5127
R1263 VCC.n447 VCC.n334 99.5127
R1264 VCC.n451 VCC.n449 99.5127
R1265 VCC.n456 VCC.n330 99.5127
R1266 VCC.n460 VCC.n458 99.5127
R1267 VCC.n464 VCC.n328 99.5127
R1268 VCC.n468 VCC.n466 99.5127
R1269 VCC.n472 VCC.n326 99.5127
R1270 VCC.n476 VCC.n474 99.5127
R1271 VCC.n480 VCC.n324 99.5127
R1272 VCC.n484 VCC.n482 99.5127
R1273 VCC.n488 VCC.n322 99.5127
R1274 VCC.n492 VCC.n490 99.5127
R1275 VCC.n496 VCC.n320 99.5127
R1276 VCC.n500 VCC.n498 99.5127
R1277 VCC.n504 VCC.n318 99.5127
R1278 VCC.n508 VCC.n506 99.5127
R1279 VCC.n512 VCC.n316 99.5127
R1280 VCC.n516 VCC.n514 99.5127
R1281 VCC.n520 VCC.n314 99.5127
R1282 VCC.n524 VCC.n522 99.5127
R1283 VCC.n528 VCC.n312 99.5127
R1284 VCC.n532 VCC.n530 99.5127
R1285 VCC.n536 VCC.n310 99.5127
R1286 VCC.n540 VCC.n538 99.5127
R1287 VCC.n268 VCC.n37 99.5127
R1288 VCC.n268 VCC.n84 99.5127
R1289 VCC.n264 VCC.n263 99.5127
R1290 VCC.n260 VCC.n259 99.5127
R1291 VCC.n256 VCC.n255 99.5127
R1292 VCC.n252 VCC.n251 99.5127
R1293 VCC.n248 VCC.n247 99.5127
R1294 VCC.n244 VCC.n243 99.5127
R1295 VCC.n240 VCC.n239 99.5127
R1296 VCC.n236 VCC.n235 99.5127
R1297 VCC.n232 VCC.n231 99.5127
R1298 VCC.n228 VCC.n227 99.5127
R1299 VCC.n224 VCC.n223 99.5127
R1300 VCC.n220 VCC.n219 99.5127
R1301 VCC.n216 VCC.n215 99.5127
R1302 VCC.n212 VCC.n211 99.5127
R1303 VCC.n208 VCC.n207 99.5127
R1304 VCC.n204 VCC.n203 99.5127
R1305 VCC.n200 VCC.n199 99.5127
R1306 VCC.n196 VCC.n195 99.5127
R1307 VCC.n192 VCC.n191 99.5127
R1308 VCC.n188 VCC.n187 99.5127
R1309 VCC.n184 VCC.n183 99.5127
R1310 VCC.n180 VCC.n179 99.5127
R1311 VCC.n175 VCC.n174 99.5127
R1312 VCC.n171 VCC.n170 99.5127
R1313 VCC.n167 VCC.n166 99.5127
R1314 VCC.n163 VCC.n162 99.5127
R1315 VCC.n159 VCC.n158 99.5127
R1316 VCC.n155 VCC.n154 99.5127
R1317 VCC.n151 VCC.n150 99.5127
R1318 VCC.n147 VCC.n146 99.5127
R1319 VCC.n143 VCC.n142 99.5127
R1320 VCC.n139 VCC.n138 99.5127
R1321 VCC.n135 VCC.n134 99.5127
R1322 VCC.n131 VCC.n130 99.5127
R1323 VCC.n127 VCC.n126 99.5127
R1324 VCC.n123 VCC.n122 99.5127
R1325 VCC.n119 VCC.n118 99.5127
R1326 VCC.n115 VCC.n114 99.5127
R1327 VCC.n111 VCC.n110 99.5127
R1328 VCC.n107 VCC.n106 99.5127
R1329 VCC.n103 VCC.n102 99.5127
R1330 VCC.n99 VCC.n98 99.5127
R1331 VCC.n95 VCC.n94 99.5127
R1332 VCC.n91 VCC.n82 99.5127
R1333 VCC.n539 VCC.n11 72.8958
R1334 VCC.n537 VCC.n11 72.8958
R1335 VCC.n531 VCC.n11 72.8958
R1336 VCC.n529 VCC.n11 72.8958
R1337 VCC.n523 VCC.n11 72.8958
R1338 VCC.n521 VCC.n11 72.8958
R1339 VCC.n515 VCC.n11 72.8958
R1340 VCC.n513 VCC.n11 72.8958
R1341 VCC.n507 VCC.n11 72.8958
R1342 VCC.n505 VCC.n11 72.8958
R1343 VCC.n499 VCC.n11 72.8958
R1344 VCC.n497 VCC.n11 72.8958
R1345 VCC.n491 VCC.n11 72.8958
R1346 VCC.n489 VCC.n11 72.8958
R1347 VCC.n483 VCC.n11 72.8958
R1348 VCC.n481 VCC.n11 72.8958
R1349 VCC.n475 VCC.n11 72.8958
R1350 VCC.n473 VCC.n11 72.8958
R1351 VCC.n467 VCC.n11 72.8958
R1352 VCC.n465 VCC.n11 72.8958
R1353 VCC.n459 VCC.n11 72.8958
R1354 VCC.n457 VCC.n11 72.8958
R1355 VCC.n450 VCC.n11 72.8958
R1356 VCC.n448 VCC.n11 72.8958
R1357 VCC.n442 VCC.n11 72.8958
R1358 VCC.n440 VCC.n11 72.8958
R1359 VCC.n434 VCC.n11 72.8958
R1360 VCC.n432 VCC.n11 72.8958
R1361 VCC.n426 VCC.n11 72.8958
R1362 VCC.n424 VCC.n11 72.8958
R1363 VCC.n418 VCC.n11 72.8958
R1364 VCC.n416 VCC.n11 72.8958
R1365 VCC.n410 VCC.n11 72.8958
R1366 VCC.n408 VCC.n11 72.8958
R1367 VCC.n402 VCC.n11 72.8958
R1368 VCC.n400 VCC.n11 72.8958
R1369 VCC.n394 VCC.n11 72.8958
R1370 VCC.n392 VCC.n11 72.8958
R1371 VCC.n386 VCC.n11 72.8958
R1372 VCC.n384 VCC.n11 72.8958
R1373 VCC.n378 VCC.n11 72.8958
R1374 VCC.n376 VCC.n11 72.8958
R1375 VCC.n370 VCC.n11 72.8958
R1376 VCC.n368 VCC.n11 72.8958
R1377 VCC.n362 VCC.n11 72.8958
R1378 VCC.n358 VCC.n11 72.8958
R1379 VCC.n270 VCC.n269 72.8958
R1380 VCC.n269 VCC.n38 72.8958
R1381 VCC.n269 VCC.n39 72.8958
R1382 VCC.n269 VCC.n40 72.8958
R1383 VCC.n269 VCC.n41 72.8958
R1384 VCC.n269 VCC.n42 72.8958
R1385 VCC.n269 VCC.n43 72.8958
R1386 VCC.n269 VCC.n44 72.8958
R1387 VCC.n269 VCC.n45 72.8958
R1388 VCC.n269 VCC.n46 72.8958
R1389 VCC.n269 VCC.n47 72.8958
R1390 VCC.n269 VCC.n48 72.8958
R1391 VCC.n269 VCC.n49 72.8958
R1392 VCC.n269 VCC.n50 72.8958
R1393 VCC.n269 VCC.n51 72.8958
R1394 VCC.n269 VCC.n52 72.8958
R1395 VCC.n269 VCC.n53 72.8958
R1396 VCC.n269 VCC.n54 72.8958
R1397 VCC.n269 VCC.n55 72.8958
R1398 VCC.n269 VCC.n56 72.8958
R1399 VCC.n269 VCC.n57 72.8958
R1400 VCC.n269 VCC.n58 72.8958
R1401 VCC.n269 VCC.n59 72.8958
R1402 VCC.n269 VCC.n60 72.8958
R1403 VCC.n269 VCC.n61 72.8958
R1404 VCC.n269 VCC.n62 72.8958
R1405 VCC.n269 VCC.n63 72.8958
R1406 VCC.n269 VCC.n64 72.8958
R1407 VCC.n269 VCC.n65 72.8958
R1408 VCC.n269 VCC.n66 72.8958
R1409 VCC.n269 VCC.n67 72.8958
R1410 VCC.n269 VCC.n68 72.8958
R1411 VCC.n269 VCC.n69 72.8958
R1412 VCC.n269 VCC.n70 72.8958
R1413 VCC.n269 VCC.n71 72.8958
R1414 VCC.n269 VCC.n72 72.8958
R1415 VCC.n269 VCC.n73 72.8958
R1416 VCC.n269 VCC.n74 72.8958
R1417 VCC.n269 VCC.n75 72.8958
R1418 VCC.n269 VCC.n76 72.8958
R1419 VCC.n269 VCC.n77 72.8958
R1420 VCC.n269 VCC.n78 72.8958
R1421 VCC.n269 VCC.n79 72.8958
R1422 VCC.n269 VCC.n80 72.8958
R1423 VCC.n269 VCC.n81 72.8958
R1424 VCC.n357 VCC.n356 44.4126
R1425 VCC.n454 VCC.n332 44.4126
R1426 VCC.n361 VCC.n358 39.2114
R1427 VCC.n362 VCC.n354 39.2114
R1428 VCC.n369 VCC.n368 39.2114
R1429 VCC.n370 VCC.n352 39.2114
R1430 VCC.n377 VCC.n376 39.2114
R1431 VCC.n378 VCC.n350 39.2114
R1432 VCC.n385 VCC.n384 39.2114
R1433 VCC.n386 VCC.n348 39.2114
R1434 VCC.n393 VCC.n392 39.2114
R1435 VCC.n394 VCC.n346 39.2114
R1436 VCC.n401 VCC.n400 39.2114
R1437 VCC.n402 VCC.n344 39.2114
R1438 VCC.n409 VCC.n408 39.2114
R1439 VCC.n410 VCC.n342 39.2114
R1440 VCC.n417 VCC.n416 39.2114
R1441 VCC.n418 VCC.n340 39.2114
R1442 VCC.n425 VCC.n424 39.2114
R1443 VCC.n426 VCC.n338 39.2114
R1444 VCC.n433 VCC.n432 39.2114
R1445 VCC.n434 VCC.n336 39.2114
R1446 VCC.n441 VCC.n440 39.2114
R1447 VCC.n442 VCC.n334 39.2114
R1448 VCC.n449 VCC.n448 39.2114
R1449 VCC.n450 VCC.n330 39.2114
R1450 VCC.n458 VCC.n457 39.2114
R1451 VCC.n459 VCC.n328 39.2114
R1452 VCC.n466 VCC.n465 39.2114
R1453 VCC.n467 VCC.n326 39.2114
R1454 VCC.n474 VCC.n473 39.2114
R1455 VCC.n475 VCC.n324 39.2114
R1456 VCC.n482 VCC.n481 39.2114
R1457 VCC.n483 VCC.n322 39.2114
R1458 VCC.n490 VCC.n489 39.2114
R1459 VCC.n491 VCC.n320 39.2114
R1460 VCC.n498 VCC.n497 39.2114
R1461 VCC.n499 VCC.n318 39.2114
R1462 VCC.n506 VCC.n505 39.2114
R1463 VCC.n507 VCC.n316 39.2114
R1464 VCC.n514 VCC.n513 39.2114
R1465 VCC.n515 VCC.n314 39.2114
R1466 VCC.n522 VCC.n521 39.2114
R1467 VCC.n523 VCC.n312 39.2114
R1468 VCC.n530 VCC.n529 39.2114
R1469 VCC.n531 VCC.n310 39.2114
R1470 VCC.n538 VCC.n537 39.2114
R1471 VCC.n539 VCC.n13 39.2114
R1472 VCC.n271 VCC.n270 39.2114
R1473 VCC.n84 VCC.n38 39.2114
R1474 VCC.n263 VCC.n39 39.2114
R1475 VCC.n259 VCC.n40 39.2114
R1476 VCC.n255 VCC.n41 39.2114
R1477 VCC.n251 VCC.n42 39.2114
R1478 VCC.n247 VCC.n43 39.2114
R1479 VCC.n243 VCC.n44 39.2114
R1480 VCC.n239 VCC.n45 39.2114
R1481 VCC.n235 VCC.n46 39.2114
R1482 VCC.n231 VCC.n47 39.2114
R1483 VCC.n227 VCC.n48 39.2114
R1484 VCC.n223 VCC.n49 39.2114
R1485 VCC.n219 VCC.n50 39.2114
R1486 VCC.n215 VCC.n51 39.2114
R1487 VCC.n211 VCC.n52 39.2114
R1488 VCC.n207 VCC.n53 39.2114
R1489 VCC.n203 VCC.n54 39.2114
R1490 VCC.n199 VCC.n55 39.2114
R1491 VCC.n195 VCC.n56 39.2114
R1492 VCC.n191 VCC.n57 39.2114
R1493 VCC.n187 VCC.n58 39.2114
R1494 VCC.n183 VCC.n59 39.2114
R1495 VCC.n179 VCC.n60 39.2114
R1496 VCC.n174 VCC.n61 39.2114
R1497 VCC.n170 VCC.n62 39.2114
R1498 VCC.n166 VCC.n63 39.2114
R1499 VCC.n162 VCC.n64 39.2114
R1500 VCC.n158 VCC.n65 39.2114
R1501 VCC.n154 VCC.n66 39.2114
R1502 VCC.n150 VCC.n67 39.2114
R1503 VCC.n146 VCC.n68 39.2114
R1504 VCC.n142 VCC.n69 39.2114
R1505 VCC.n138 VCC.n70 39.2114
R1506 VCC.n134 VCC.n71 39.2114
R1507 VCC.n130 VCC.n72 39.2114
R1508 VCC.n126 VCC.n73 39.2114
R1509 VCC.n122 VCC.n74 39.2114
R1510 VCC.n118 VCC.n75 39.2114
R1511 VCC.n114 VCC.n76 39.2114
R1512 VCC.n110 VCC.n77 39.2114
R1513 VCC.n106 VCC.n78 39.2114
R1514 VCC.n102 VCC.n79 39.2114
R1515 VCC.n98 VCC.n80 39.2114
R1516 VCC.n94 VCC.n81 39.2114
R1517 VCC.n540 VCC.n539 39.2114
R1518 VCC.n537 VCC.n536 39.2114
R1519 VCC.n532 VCC.n531 39.2114
R1520 VCC.n529 VCC.n528 39.2114
R1521 VCC.n524 VCC.n523 39.2114
R1522 VCC.n521 VCC.n520 39.2114
R1523 VCC.n516 VCC.n515 39.2114
R1524 VCC.n513 VCC.n512 39.2114
R1525 VCC.n508 VCC.n507 39.2114
R1526 VCC.n505 VCC.n504 39.2114
R1527 VCC.n500 VCC.n499 39.2114
R1528 VCC.n497 VCC.n496 39.2114
R1529 VCC.n492 VCC.n491 39.2114
R1530 VCC.n489 VCC.n488 39.2114
R1531 VCC.n484 VCC.n483 39.2114
R1532 VCC.n481 VCC.n480 39.2114
R1533 VCC.n476 VCC.n475 39.2114
R1534 VCC.n473 VCC.n472 39.2114
R1535 VCC.n468 VCC.n467 39.2114
R1536 VCC.n465 VCC.n464 39.2114
R1537 VCC.n460 VCC.n459 39.2114
R1538 VCC.n457 VCC.n456 39.2114
R1539 VCC.n451 VCC.n450 39.2114
R1540 VCC.n448 VCC.n447 39.2114
R1541 VCC.n443 VCC.n442 39.2114
R1542 VCC.n440 VCC.n439 39.2114
R1543 VCC.n435 VCC.n434 39.2114
R1544 VCC.n432 VCC.n431 39.2114
R1545 VCC.n427 VCC.n426 39.2114
R1546 VCC.n424 VCC.n423 39.2114
R1547 VCC.n419 VCC.n418 39.2114
R1548 VCC.n416 VCC.n415 39.2114
R1549 VCC.n411 VCC.n410 39.2114
R1550 VCC.n408 VCC.n407 39.2114
R1551 VCC.n403 VCC.n402 39.2114
R1552 VCC.n400 VCC.n399 39.2114
R1553 VCC.n395 VCC.n394 39.2114
R1554 VCC.n392 VCC.n391 39.2114
R1555 VCC.n387 VCC.n386 39.2114
R1556 VCC.n384 VCC.n383 39.2114
R1557 VCC.n379 VCC.n378 39.2114
R1558 VCC.n376 VCC.n375 39.2114
R1559 VCC.n371 VCC.n370 39.2114
R1560 VCC.n368 VCC.n367 39.2114
R1561 VCC.n363 VCC.n362 39.2114
R1562 VCC.n358 VCC.n9 39.2114
R1563 VCC.n270 VCC.n37 39.2114
R1564 VCC.n264 VCC.n38 39.2114
R1565 VCC.n260 VCC.n39 39.2114
R1566 VCC.n256 VCC.n40 39.2114
R1567 VCC.n252 VCC.n41 39.2114
R1568 VCC.n248 VCC.n42 39.2114
R1569 VCC.n244 VCC.n43 39.2114
R1570 VCC.n240 VCC.n44 39.2114
R1571 VCC.n236 VCC.n45 39.2114
R1572 VCC.n232 VCC.n46 39.2114
R1573 VCC.n228 VCC.n47 39.2114
R1574 VCC.n224 VCC.n48 39.2114
R1575 VCC.n220 VCC.n49 39.2114
R1576 VCC.n216 VCC.n50 39.2114
R1577 VCC.n212 VCC.n51 39.2114
R1578 VCC.n208 VCC.n52 39.2114
R1579 VCC.n204 VCC.n53 39.2114
R1580 VCC.n200 VCC.n54 39.2114
R1581 VCC.n196 VCC.n55 39.2114
R1582 VCC.n192 VCC.n56 39.2114
R1583 VCC.n188 VCC.n57 39.2114
R1584 VCC.n184 VCC.n58 39.2114
R1585 VCC.n180 VCC.n59 39.2114
R1586 VCC.n175 VCC.n60 39.2114
R1587 VCC.n171 VCC.n61 39.2114
R1588 VCC.n167 VCC.n62 39.2114
R1589 VCC.n163 VCC.n63 39.2114
R1590 VCC.n159 VCC.n64 39.2114
R1591 VCC.n155 VCC.n65 39.2114
R1592 VCC.n151 VCC.n66 39.2114
R1593 VCC.n147 VCC.n67 39.2114
R1594 VCC.n143 VCC.n68 39.2114
R1595 VCC.n139 VCC.n69 39.2114
R1596 VCC.n135 VCC.n70 39.2114
R1597 VCC.n131 VCC.n71 39.2114
R1598 VCC.n127 VCC.n72 39.2114
R1599 VCC.n123 VCC.n73 39.2114
R1600 VCC.n119 VCC.n74 39.2114
R1601 VCC.n115 VCC.n75 39.2114
R1602 VCC.n111 VCC.n76 39.2114
R1603 VCC.n107 VCC.n77 39.2114
R1604 VCC.n103 VCC.n78 39.2114
R1605 VCC.n99 VCC.n79 39.2114
R1606 VCC.n95 VCC.n80 39.2114
R1607 VCC.n91 VCC.n81 39.2114
R1608 VCC.n359 VCC.n7 30.7874
R1609 VCC.n543 VCC.n542 30.7874
R1610 VCC.n273 VCC.n272 30.7874
R1611 VCC.n90 VCC.n29 30.7874
R1612 VCC.n177 VCC.n89 29.2853
R1613 VCC.n87 VCC.n86 29.2853
R1614 VCC.n269 VCC.n83 24.0854
R1615 VCC.n546 VCC.n11 24.0854
R1616 VCC.n283 VCC.n30 19.3944
R1617 VCC.n283 VCC.n28 19.3944
R1618 VCC.n287 VCC.n28 19.3944
R1619 VCC.n287 VCC.n21 19.3944
R1620 VCC.n295 VCC.n21 19.3944
R1621 VCC.n295 VCC.n19 19.3944
R1622 VCC.n299 VCC.n19 19.3944
R1623 VCC.n299 VCC.n16 19.3944
R1624 VCC.n306 VCC.n16 19.3944
R1625 VCC.n306 VCC.n14 19.3944
R1626 VCC.n544 VCC.n14 19.3944
R1627 VCC.n279 VCC.n34 19.3944
R1628 VCC.n279 VCC.n35 19.3944
R1629 VCC.n275 VCC.n35 19.3944
R1630 VCC.n275 VCC.n25 19.3944
R1631 VCC.n25 VCC.n2 19.3944
R1632 VCC.n555 VCC.n2 19.3944
R1633 VCC.n555 VCC.n554 19.3944
R1634 VCC.n554 VCC.n553 19.3944
R1635 VCC.n553 VCC.n6 19.3944
R1636 VCC.n549 VCC.n6 19.3944
R1637 VCC.n549 VCC.n548 19.3944
R1638 VCC.n281 VCC.n26 14.2519
R1639 VCC.n289 VCC.n26 14.2519
R1640 VCC.n290 VCC.n289 14.2519
R1641 VCC.n302 VCC.n301 14.2519
R1642 VCC.n304 VCC.n302 14.2519
R1643 VCC.n546 VCC.n10 14.2519
R1644 VCC.n293 VCC.t2 13.8244
R1645 VCC.t1 VCC.n23 12.6843
R1646 VCC.n301 VCC.t0 11.5442
R1647 VCC.n83 VCC.t4 10.9741
R1648 VCC.n360 VCC.n359 10.6151
R1649 VCC.n365 VCC.n364 10.6151
R1650 VCC.n366 VCC.n365 10.6151
R1651 VCC.n366 VCC.n353 10.6151
R1652 VCC.n372 VCC.n353 10.6151
R1653 VCC.n373 VCC.n372 10.6151
R1654 VCC.n374 VCC.n373 10.6151
R1655 VCC.n374 VCC.n351 10.6151
R1656 VCC.n380 VCC.n351 10.6151
R1657 VCC.n381 VCC.n380 10.6151
R1658 VCC.n382 VCC.n381 10.6151
R1659 VCC.n382 VCC.n349 10.6151
R1660 VCC.n388 VCC.n349 10.6151
R1661 VCC.n389 VCC.n388 10.6151
R1662 VCC.n390 VCC.n389 10.6151
R1663 VCC.n390 VCC.n347 10.6151
R1664 VCC.n396 VCC.n347 10.6151
R1665 VCC.n397 VCC.n396 10.6151
R1666 VCC.n398 VCC.n397 10.6151
R1667 VCC.n398 VCC.n345 10.6151
R1668 VCC.n404 VCC.n345 10.6151
R1669 VCC.n405 VCC.n404 10.6151
R1670 VCC.n406 VCC.n405 10.6151
R1671 VCC.n406 VCC.n343 10.6151
R1672 VCC.n412 VCC.n343 10.6151
R1673 VCC.n413 VCC.n412 10.6151
R1674 VCC.n414 VCC.n413 10.6151
R1675 VCC.n414 VCC.n341 10.6151
R1676 VCC.n420 VCC.n341 10.6151
R1677 VCC.n421 VCC.n420 10.6151
R1678 VCC.n422 VCC.n421 10.6151
R1679 VCC.n422 VCC.n339 10.6151
R1680 VCC.n428 VCC.n339 10.6151
R1681 VCC.n429 VCC.n428 10.6151
R1682 VCC.n430 VCC.n429 10.6151
R1683 VCC.n430 VCC.n337 10.6151
R1684 VCC.n436 VCC.n337 10.6151
R1685 VCC.n437 VCC.n436 10.6151
R1686 VCC.n438 VCC.n437 10.6151
R1687 VCC.n438 VCC.n335 10.6151
R1688 VCC.n444 VCC.n335 10.6151
R1689 VCC.n445 VCC.n444 10.6151
R1690 VCC.n446 VCC.n445 10.6151
R1691 VCC.n446 VCC.n333 10.6151
R1692 VCC.n452 VCC.n333 10.6151
R1693 VCC.n453 VCC.n452 10.6151
R1694 VCC.n455 VCC.n329 10.6151
R1695 VCC.n461 VCC.n329 10.6151
R1696 VCC.n462 VCC.n461 10.6151
R1697 VCC.n463 VCC.n462 10.6151
R1698 VCC.n463 VCC.n327 10.6151
R1699 VCC.n469 VCC.n327 10.6151
R1700 VCC.n470 VCC.n469 10.6151
R1701 VCC.n471 VCC.n470 10.6151
R1702 VCC.n471 VCC.n325 10.6151
R1703 VCC.n477 VCC.n325 10.6151
R1704 VCC.n478 VCC.n477 10.6151
R1705 VCC.n479 VCC.n478 10.6151
R1706 VCC.n479 VCC.n323 10.6151
R1707 VCC.n485 VCC.n323 10.6151
R1708 VCC.n486 VCC.n485 10.6151
R1709 VCC.n487 VCC.n486 10.6151
R1710 VCC.n487 VCC.n321 10.6151
R1711 VCC.n493 VCC.n321 10.6151
R1712 VCC.n494 VCC.n493 10.6151
R1713 VCC.n495 VCC.n494 10.6151
R1714 VCC.n495 VCC.n319 10.6151
R1715 VCC.n501 VCC.n319 10.6151
R1716 VCC.n502 VCC.n501 10.6151
R1717 VCC.n503 VCC.n502 10.6151
R1718 VCC.n503 VCC.n317 10.6151
R1719 VCC.n509 VCC.n317 10.6151
R1720 VCC.n510 VCC.n509 10.6151
R1721 VCC.n511 VCC.n510 10.6151
R1722 VCC.n511 VCC.n315 10.6151
R1723 VCC.n517 VCC.n315 10.6151
R1724 VCC.n518 VCC.n517 10.6151
R1725 VCC.n519 VCC.n518 10.6151
R1726 VCC.n519 VCC.n313 10.6151
R1727 VCC.n525 VCC.n313 10.6151
R1728 VCC.n526 VCC.n525 10.6151
R1729 VCC.n527 VCC.n526 10.6151
R1730 VCC.n527 VCC.n311 10.6151
R1731 VCC.n533 VCC.n311 10.6151
R1732 VCC.n534 VCC.n533 10.6151
R1733 VCC.n535 VCC.n534 10.6151
R1734 VCC.n535 VCC.n309 10.6151
R1735 VCC.n541 VCC.n309 10.6151
R1736 VCC.n542 VCC.n541 10.6151
R1737 VCC.n272 VCC.n36 10.6151
R1738 VCC.n267 VCC.n266 10.6151
R1739 VCC.n266 VCC.n265 10.6151
R1740 VCC.n265 VCC.n262 10.6151
R1741 VCC.n262 VCC.n261 10.6151
R1742 VCC.n261 VCC.n258 10.6151
R1743 VCC.n258 VCC.n257 10.6151
R1744 VCC.n257 VCC.n254 10.6151
R1745 VCC.n254 VCC.n253 10.6151
R1746 VCC.n253 VCC.n250 10.6151
R1747 VCC.n250 VCC.n249 10.6151
R1748 VCC.n249 VCC.n246 10.6151
R1749 VCC.n246 VCC.n245 10.6151
R1750 VCC.n245 VCC.n242 10.6151
R1751 VCC.n242 VCC.n241 10.6151
R1752 VCC.n241 VCC.n238 10.6151
R1753 VCC.n238 VCC.n237 10.6151
R1754 VCC.n237 VCC.n234 10.6151
R1755 VCC.n234 VCC.n233 10.6151
R1756 VCC.n233 VCC.n230 10.6151
R1757 VCC.n230 VCC.n229 10.6151
R1758 VCC.n229 VCC.n226 10.6151
R1759 VCC.n226 VCC.n225 10.6151
R1760 VCC.n225 VCC.n222 10.6151
R1761 VCC.n222 VCC.n221 10.6151
R1762 VCC.n221 VCC.n218 10.6151
R1763 VCC.n218 VCC.n217 10.6151
R1764 VCC.n217 VCC.n214 10.6151
R1765 VCC.n214 VCC.n213 10.6151
R1766 VCC.n213 VCC.n210 10.6151
R1767 VCC.n210 VCC.n209 10.6151
R1768 VCC.n209 VCC.n206 10.6151
R1769 VCC.n206 VCC.n205 10.6151
R1770 VCC.n205 VCC.n202 10.6151
R1771 VCC.n202 VCC.n201 10.6151
R1772 VCC.n201 VCC.n198 10.6151
R1773 VCC.n198 VCC.n197 10.6151
R1774 VCC.n197 VCC.n194 10.6151
R1775 VCC.n194 VCC.n193 10.6151
R1776 VCC.n193 VCC.n190 10.6151
R1777 VCC.n190 VCC.n189 10.6151
R1778 VCC.n189 VCC.n186 10.6151
R1779 VCC.n186 VCC.n185 10.6151
R1780 VCC.n185 VCC.n182 10.6151
R1781 VCC.n182 VCC.n181 10.6151
R1782 VCC.n181 VCC.n178 10.6151
R1783 VCC.n176 VCC.n173 10.6151
R1784 VCC.n173 VCC.n172 10.6151
R1785 VCC.n172 VCC.n169 10.6151
R1786 VCC.n169 VCC.n168 10.6151
R1787 VCC.n168 VCC.n165 10.6151
R1788 VCC.n165 VCC.n164 10.6151
R1789 VCC.n164 VCC.n161 10.6151
R1790 VCC.n161 VCC.n160 10.6151
R1791 VCC.n160 VCC.n157 10.6151
R1792 VCC.n157 VCC.n156 10.6151
R1793 VCC.n156 VCC.n153 10.6151
R1794 VCC.n153 VCC.n152 10.6151
R1795 VCC.n152 VCC.n149 10.6151
R1796 VCC.n149 VCC.n148 10.6151
R1797 VCC.n148 VCC.n145 10.6151
R1798 VCC.n145 VCC.n144 10.6151
R1799 VCC.n144 VCC.n141 10.6151
R1800 VCC.n141 VCC.n140 10.6151
R1801 VCC.n140 VCC.n137 10.6151
R1802 VCC.n137 VCC.n136 10.6151
R1803 VCC.n136 VCC.n133 10.6151
R1804 VCC.n133 VCC.n132 10.6151
R1805 VCC.n132 VCC.n129 10.6151
R1806 VCC.n129 VCC.n128 10.6151
R1807 VCC.n128 VCC.n125 10.6151
R1808 VCC.n125 VCC.n124 10.6151
R1809 VCC.n124 VCC.n121 10.6151
R1810 VCC.n121 VCC.n120 10.6151
R1811 VCC.n120 VCC.n117 10.6151
R1812 VCC.n117 VCC.n116 10.6151
R1813 VCC.n116 VCC.n113 10.6151
R1814 VCC.n113 VCC.n112 10.6151
R1815 VCC.n112 VCC.n109 10.6151
R1816 VCC.n109 VCC.n108 10.6151
R1817 VCC.n108 VCC.n105 10.6151
R1818 VCC.n105 VCC.n104 10.6151
R1819 VCC.n104 VCC.n101 10.6151
R1820 VCC.n101 VCC.n100 10.6151
R1821 VCC.n100 VCC.n97 10.6151
R1822 VCC.n97 VCC.n96 10.6151
R1823 VCC.n96 VCC.n93 10.6151
R1824 VCC.n93 VCC.n92 10.6151
R1825 VCC.n92 VCC.n90 10.6151
R1826 VCC.n356 VCC.n355 10.4732
R1827 VCC.n332 VCC.n331 10.4732
R1828 VCC.n89 VCC.n88 10.4732
R1829 VCC.n86 VCC.n85 10.4732
R1830 VCC.n454 VCC.n453 9.83465
R1831 VCC.n178 VCC.n177 9.83465
R1832 VCC.n554 VCC.n0 9.3005
R1833 VCC.n553 VCC.n552 9.3005
R1834 VCC.n551 VCC.n6 9.3005
R1835 VCC.n550 VCC.n549 9.3005
R1836 VCC.n548 VCC.n7 9.3005
R1837 VCC.n284 VCC.n283 9.3005
R1838 VCC.n285 VCC.n28 9.3005
R1839 VCC.n287 VCC.n286 9.3005
R1840 VCC.n21 VCC.n20 9.3005
R1841 VCC.n296 VCC.n295 9.3005
R1842 VCC.n297 VCC.n19 9.3005
R1843 VCC.n299 VCC.n298 9.3005
R1844 VCC.n16 VCC.n15 9.3005
R1845 VCC.n307 VCC.n306 9.3005
R1846 VCC.n308 VCC.n14 9.3005
R1847 VCC.n544 VCC.n543 9.3005
R1848 VCC.n30 VCC.n29 9.3005
R1849 VCC.n273 VCC.n34 9.3005
R1850 VCC.n279 VCC.n278 9.3005
R1851 VCC.n277 VCC.n35 9.3005
R1852 VCC.n276 VCC.n275 9.3005
R1853 VCC.n274 VCC.n25 9.3005
R1854 VCC.n2 VCC.n1 9.3005
R1855 VCC VCC.n555 9.3005
R1856 VCC.n360 VCC.n357 7.96148
R1857 VCC.n87 VCC.n36 7.96148
R1858 VCC.t8 VCC.n10 7.83878
R1859 VCC.n304 VCC.t8 6.41364
R1860 VCC.n281 VCC.t4 3.27833
R1861 VCC.n23 VCC.t0 2.70827
R1862 VCC.n364 VCC.n357 2.65416
R1863 VCC.n267 VCC.n87 2.65416
R1864 VCC.n293 VCC.t1 1.56816
R1865 VCC.n455 VCC.n454 0.780988
R1866 VCC.n177 VCC.n176 0.780988
R1867 VCC.n290 VCC.t2 0.428043
R1868 VCC VCC.n0 0.152939
R1869 VCC.n552 VCC.n0 0.152939
R1870 VCC.n552 VCC.n551 0.152939
R1871 VCC.n551 VCC.n550 0.152939
R1872 VCC.n550 VCC.n7 0.152939
R1873 VCC.n284 VCC.n29 0.152939
R1874 VCC.n285 VCC.n284 0.152939
R1875 VCC.n286 VCC.n285 0.152939
R1876 VCC.n286 VCC.n20 0.152939
R1877 VCC.n296 VCC.n20 0.152939
R1878 VCC.n297 VCC.n296 0.152939
R1879 VCC.n298 VCC.n297 0.152939
R1880 VCC.n298 VCC.n15 0.152939
R1881 VCC.n307 VCC.n15 0.152939
R1882 VCC.n308 VCC.n307 0.152939
R1883 VCC.n543 VCC.n308 0.152939
R1884 VCC.n278 VCC.n273 0.152939
R1885 VCC.n278 VCC.n277 0.152939
R1886 VCC.n277 VCC.n276 0.152939
R1887 VCC.n276 VCC.n274 0.152939
R1888 VCC.n274 VCC.n1 0.152939
R1889 VCC VCC.n1 0.1255
C0 VCC VOUT 8.94991f
C1 VOUT VSS 6.484709f
C2 VGP VSS 0.085018f
C3 VGN VSS 0.027265f
C4 VIN VSS 0.020864f
C5 VCC VSS 35.574257f
C6 VCC.n0 VSS 0.004192f
C7 VCC.n1 VSS 0.004652f
C8 VCC.n2 VSS 0.003374f
C9 VCC.n3 VSS 0.004192f
C10 VCC.n4 VSS 0.004192f
C11 VCC.n5 VSS 0.004192f
C12 VCC.n6 VSS 0.003374f
C13 VCC.n7 VSS 0.014004f
C14 VCC.n8 VSS 0.004192f
C15 VCC.n9 VSS 0.008058f
C16 VCC.n10 VSS 0.264072f
C17 VCC.n11 VSS 0.638884f
C18 VCC.n12 VSS 0.004192f
C19 VCC.n13 VSS 0.008058f
C20 VCC.n14 VSS 0.003374f
C21 VCC.n15 VSS 0.004192f
C22 VCC.n16 VSS 0.003374f
C23 VCC.n17 VSS 0.004192f
C24 VCC.t0 VSS 0.170369f
C25 VCC.n18 VSS 0.004192f
C26 VCC.n19 VSS 0.003374f
C27 VCC.n20 VSS 0.004192f
C28 VCC.n21 VSS 0.003374f
C29 VCC.n22 VSS 0.004192f
C30 VCC.t2 VSS 0.170369f
C31 VCC.n23 VSS 0.183999f
C32 VCC.t1 VSS 0.170369f
C33 VCC.n24 VSS 0.004192f
C34 VCC.n25 VSS 0.003374f
C35 VCC.n26 VSS 0.340738f
C36 VCC.n27 VSS 0.004192f
C37 VCC.n28 VSS 0.003374f
C38 VCC.n29 VSS 0.014004f
C39 VCC.n30 VSS 0.0028f
C40 VCC.n31 VSS 0.008247f
C41 VCC.t4 VSS 0.170369f
C42 VCC.n32 VSS 0.008247f
C43 VCC.n33 VSS 0.004192f
C44 VCC.n34 VSS 0.0028f
C45 VCC.n35 VSS 0.003374f
C46 VCC.n36 VSS 0.002494f
C47 VCC.n37 VSS 0.00285f
C48 VCC.n82 VSS 0.008058f
C49 VCC.n83 VSS 0.419108f
C50 VCC.n84 VSS 0.00285f
C51 VCC.t5 VSS 0.099161f
C52 VCC.t6 VSS 0.101764f
C53 VCC.t3 VSS 0.044426f
C54 VCC.n85 VSS 0.117132f
C55 VCC.n86 VSS 0.103839f
C56 VCC.n87 VSS 0.003972f
C57 VCC.t12 VSS 0.099161f
C58 VCC.t13 VSS 0.101764f
C59 VCC.t11 VSS 0.044426f
C60 VCC.n88 VSS 0.117132f
C61 VCC.n89 VSS 0.103839f
C62 VCC.n90 VSS 0.005738f
C63 VCC.n91 VSS 0.00285f
C64 VCC.n92 VSS 0.00285f
C65 VCC.n93 VSS 0.00285f
C66 VCC.n94 VSS 0.00285f
C67 VCC.n95 VSS 0.00285f
C68 VCC.n96 VSS 0.00285f
C69 VCC.n97 VSS 0.00285f
C70 VCC.n98 VSS 0.00285f
C71 VCC.n99 VSS 0.00285f
C72 VCC.n100 VSS 0.00285f
C73 VCC.n101 VSS 0.00285f
C74 VCC.n102 VSS 0.00285f
C75 VCC.n103 VSS 0.00285f
C76 VCC.n104 VSS 0.00285f
C77 VCC.n105 VSS 0.00285f
C78 VCC.n106 VSS 0.00285f
C79 VCC.n107 VSS 0.00285f
C80 VCC.n108 VSS 0.00285f
C81 VCC.n109 VSS 0.00285f
C82 VCC.n110 VSS 0.00285f
C83 VCC.n111 VSS 0.00285f
C84 VCC.n112 VSS 0.00285f
C85 VCC.n113 VSS 0.00285f
C86 VCC.n114 VSS 0.00285f
C87 VCC.n115 VSS 0.00285f
C88 VCC.n116 VSS 0.00285f
C89 VCC.n117 VSS 0.00285f
C90 VCC.n118 VSS 0.00285f
C91 VCC.n119 VSS 0.00285f
C92 VCC.n120 VSS 0.00285f
C93 VCC.n121 VSS 0.00285f
C94 VCC.n122 VSS 0.00285f
C95 VCC.n123 VSS 0.00285f
C96 VCC.n124 VSS 0.00285f
C97 VCC.n125 VSS 0.00285f
C98 VCC.n126 VSS 0.00285f
C99 VCC.n127 VSS 0.00285f
C100 VCC.n128 VSS 0.00285f
C101 VCC.n129 VSS 0.00285f
C102 VCC.n130 VSS 0.00285f
C103 VCC.n131 VSS 0.00285f
C104 VCC.n132 VSS 0.00285f
C105 VCC.n133 VSS 0.00285f
C106 VCC.n134 VSS 0.00285f
C107 VCC.n135 VSS 0.00285f
C108 VCC.n136 VSS 0.00285f
C109 VCC.n137 VSS 0.00285f
C110 VCC.n138 VSS 0.00285f
C111 VCC.n139 VSS 0.00285f
C112 VCC.n140 VSS 0.00285f
C113 VCC.n141 VSS 0.00285f
C114 VCC.n142 VSS 0.00285f
C115 VCC.n143 VSS 0.00285f
C116 VCC.n144 VSS 0.00285f
C117 VCC.n145 VSS 0.00285f
C118 VCC.n146 VSS 0.00285f
C119 VCC.n147 VSS 0.00285f
C120 VCC.n148 VSS 0.00285f
C121 VCC.n149 VSS 0.00285f
C122 VCC.n150 VSS 0.00285f
C123 VCC.n151 VSS 0.00285f
C124 VCC.n152 VSS 0.00285f
C125 VCC.n153 VSS 0.00285f
C126 VCC.n154 VSS 0.00285f
C127 VCC.n155 VSS 0.00285f
C128 VCC.n156 VSS 0.00285f
C129 VCC.n157 VSS 0.00285f
C130 VCC.n158 VSS 0.00285f
C131 VCC.n159 VSS 0.00285f
C132 VCC.n160 VSS 0.00285f
C133 VCC.n161 VSS 0.00285f
C134 VCC.n162 VSS 0.00285f
C135 VCC.n163 VSS 0.00285f
C136 VCC.n164 VSS 0.00285f
C137 VCC.n165 VSS 0.00285f
C138 VCC.n166 VSS 0.00285f
C139 VCC.n167 VSS 0.00285f
C140 VCC.n168 VSS 0.00285f
C141 VCC.n169 VSS 0.00285f
C142 VCC.n170 VSS 0.00285f
C143 VCC.n171 VSS 0.00285f
C144 VCC.n172 VSS 0.00285f
C145 VCC.n173 VSS 0.00285f
C146 VCC.n174 VSS 0.00285f
C147 VCC.n175 VSS 0.00285f
C148 VCC.n176 VSS 0.00153f
C149 VCC.n177 VSS 0.003972f
C150 VCC.n178 VSS 0.002745f
C151 VCC.n179 VSS 0.00285f
C152 VCC.n180 VSS 0.00285f
C153 VCC.n181 VSS 0.00285f
C154 VCC.n182 VSS 0.00285f
C155 VCC.n183 VSS 0.00285f
C156 VCC.n184 VSS 0.00285f
C157 VCC.n185 VSS 0.00285f
C158 VCC.n186 VSS 0.00285f
C159 VCC.n187 VSS 0.00285f
C160 VCC.n188 VSS 0.00285f
C161 VCC.n189 VSS 0.00285f
C162 VCC.n190 VSS 0.00285f
C163 VCC.n191 VSS 0.00285f
C164 VCC.n192 VSS 0.00285f
C165 VCC.n193 VSS 0.00285f
C166 VCC.n194 VSS 0.00285f
C167 VCC.n195 VSS 0.00285f
C168 VCC.n196 VSS 0.00285f
C169 VCC.n197 VSS 0.00285f
C170 VCC.n198 VSS 0.00285f
C171 VCC.n199 VSS 0.00285f
C172 VCC.n200 VSS 0.00285f
C173 VCC.n201 VSS 0.00285f
C174 VCC.n202 VSS 0.00285f
C175 VCC.n203 VSS 0.00285f
C176 VCC.n204 VSS 0.00285f
C177 VCC.n205 VSS 0.00285f
C178 VCC.n206 VSS 0.00285f
C179 VCC.n207 VSS 0.00285f
C180 VCC.n208 VSS 0.00285f
C181 VCC.n209 VSS 0.00285f
C182 VCC.n210 VSS 0.00285f
C183 VCC.n211 VSS 0.00285f
C184 VCC.n212 VSS 0.00285f
C185 VCC.n213 VSS 0.00285f
C186 VCC.n214 VSS 0.00285f
C187 VCC.n215 VSS 0.00285f
C188 VCC.n216 VSS 0.00285f
C189 VCC.n217 VSS 0.00285f
C190 VCC.n218 VSS 0.00285f
C191 VCC.n219 VSS 0.00285f
C192 VCC.n220 VSS 0.00285f
C193 VCC.n221 VSS 0.00285f
C194 VCC.n222 VSS 0.00285f
C195 VCC.n223 VSS 0.00285f
C196 VCC.n224 VSS 0.00285f
C197 VCC.n225 VSS 0.00285f
C198 VCC.n226 VSS 0.00285f
C199 VCC.n227 VSS 0.00285f
C200 VCC.n228 VSS 0.00285f
C201 VCC.n229 VSS 0.00285f
C202 VCC.n230 VSS 0.00285f
C203 VCC.n231 VSS 0.00285f
C204 VCC.n232 VSS 0.00285f
C205 VCC.n233 VSS 0.00285f
C206 VCC.n234 VSS 0.00285f
C207 VCC.n235 VSS 0.00285f
C208 VCC.n236 VSS 0.00285f
C209 VCC.n237 VSS 0.00285f
C210 VCC.n238 VSS 0.00285f
C211 VCC.n239 VSS 0.00285f
C212 VCC.n240 VSS 0.00285f
C213 VCC.n241 VSS 0.00285f
C214 VCC.n242 VSS 0.00285f
C215 VCC.n243 VSS 0.00285f
C216 VCC.n244 VSS 0.00285f
C217 VCC.n245 VSS 0.00285f
C218 VCC.n246 VSS 0.00285f
C219 VCC.n247 VSS 0.00285f
C220 VCC.n248 VSS 0.00285f
C221 VCC.n249 VSS 0.00285f
C222 VCC.n250 VSS 0.00285f
C223 VCC.n251 VSS 0.00285f
C224 VCC.n252 VSS 0.00285f
C225 VCC.n253 VSS 0.00285f
C226 VCC.n254 VSS 0.00285f
C227 VCC.n255 VSS 0.00285f
C228 VCC.n256 VSS 0.00285f
C229 VCC.n257 VSS 0.00285f
C230 VCC.n258 VSS 0.00285f
C231 VCC.n259 VSS 0.00285f
C232 VCC.n260 VSS 0.00285f
C233 VCC.n261 VSS 0.00285f
C234 VCC.n262 VSS 0.00285f
C235 VCC.n263 VSS 0.00285f
C236 VCC.n264 VSS 0.00285f
C237 VCC.n265 VSS 0.00285f
C238 VCC.n266 VSS 0.00285f
C239 VCC.n267 VSS 0.001781f
C240 VCC.n268 VSS 0.00285f
C241 VCC.n269 VSS 0.638884f
C242 VCC.n271 VSS 0.008058f
C243 VCC.n272 VSS 0.005738f
C244 VCC.n273 VSS 0.014004f
C245 VCC.n274 VSS 0.004192f
C246 VCC.n275 VSS 0.003374f
C247 VCC.n276 VSS 0.004192f
C248 VCC.n277 VSS 0.004192f
C249 VCC.n278 VSS 0.004192f
C250 VCC.n279 VSS 0.003374f
C251 VCC.n280 VSS 0.004192f
C252 VCC.n281 VSS 0.209554f
C253 VCC.n282 VSS 0.004192f
C254 VCC.n283 VSS 0.003374f
C255 VCC.n284 VSS 0.004192f
C256 VCC.n285 VSS 0.004192f
C257 VCC.n286 VSS 0.004192f
C258 VCC.n287 VSS 0.003374f
C259 VCC.n288 VSS 0.004192f
C260 VCC.n289 VSS 0.340738f
C261 VCC.n290 VSS 0.17548f
C262 VCC.n291 VSS 0.004192f
C263 VCC.n292 VSS 0.004192f
C264 VCC.n293 VSS 0.183999f
C265 VCC.n294 VSS 0.004192f
C266 VCC.n295 VSS 0.003374f
C267 VCC.n296 VSS 0.004192f
C268 VCC.n297 VSS 0.004192f
C269 VCC.n298 VSS 0.004192f
C270 VCC.n299 VSS 0.003374f
C271 VCC.n300 VSS 0.004192f
C272 VCC.n301 VSS 0.308368f
C273 VCC.n302 VSS 0.340738f
C274 VCC.t8 VSS 0.170369f
C275 VCC.n303 VSS 0.004192f
C276 VCC.n304 VSS 0.247035f
C277 VCC.n305 VSS 0.004192f
C278 VCC.n306 VSS 0.003374f
C279 VCC.n307 VSS 0.004192f
C280 VCC.n308 VSS 0.004192f
C281 VCC.n309 VSS 0.00285f
C282 VCC.n310 VSS 0.00285f
C283 VCC.n311 VSS 0.00285f
C284 VCC.n312 VSS 0.00285f
C285 VCC.n313 VSS 0.00285f
C286 VCC.n314 VSS 0.00285f
C287 VCC.n315 VSS 0.00285f
C288 VCC.n316 VSS 0.00285f
C289 VCC.n317 VSS 0.00285f
C290 VCC.n318 VSS 0.00285f
C291 VCC.n319 VSS 0.00285f
C292 VCC.n320 VSS 0.00285f
C293 VCC.n321 VSS 0.00285f
C294 VCC.n322 VSS 0.00285f
C295 VCC.n323 VSS 0.00285f
C296 VCC.n324 VSS 0.00285f
C297 VCC.n325 VSS 0.00285f
C298 VCC.n326 VSS 0.00285f
C299 VCC.n327 VSS 0.00285f
C300 VCC.n328 VSS 0.00285f
C301 VCC.n329 VSS 0.00285f
C302 VCC.n330 VSS 0.00285f
C303 VCC.t10 VSS 0.099161f
C304 VCC.t9 VSS 0.101764f
C305 VCC.t7 VSS 0.044426f
C306 VCC.n331 VSS 0.117132f
C307 VCC.n332 VSS 0.105154f
C308 VCC.n333 VSS 0.00285f
C309 VCC.n334 VSS 0.00285f
C310 VCC.n335 VSS 0.00285f
C311 VCC.n336 VSS 0.00285f
C312 VCC.n337 VSS 0.00285f
C313 VCC.n338 VSS 0.00285f
C314 VCC.n339 VSS 0.00285f
C315 VCC.n340 VSS 0.00285f
C316 VCC.n341 VSS 0.00285f
C317 VCC.n342 VSS 0.00285f
C318 VCC.n343 VSS 0.00285f
C319 VCC.n344 VSS 0.00285f
C320 VCC.n345 VSS 0.00285f
C321 VCC.n346 VSS 0.00285f
C322 VCC.n347 VSS 0.00285f
C323 VCC.n348 VSS 0.00285f
C324 VCC.n349 VSS 0.00285f
C325 VCC.n350 VSS 0.00285f
C326 VCC.n351 VSS 0.00285f
C327 VCC.n352 VSS 0.00285f
C328 VCC.n353 VSS 0.00285f
C329 VCC.n354 VSS 0.00285f
C330 VCC.t16 VSS 0.099161f
C331 VCC.t15 VSS 0.101764f
C332 VCC.t14 VSS 0.044426f
C333 VCC.n355 VSS 0.117132f
C334 VCC.n356 VSS 0.105154f
C335 VCC.n357 VSS 0.005288f
C336 VCC.n359 VSS 0.005738f
C337 VCC.n360 VSS 0.002494f
C338 VCC.n361 VSS 0.00285f
C339 VCC.n363 VSS 0.00285f
C340 VCC.n364 VSS 0.001781f
C341 VCC.n365 VSS 0.00285f
C342 VCC.n366 VSS 0.00285f
C343 VCC.n367 VSS 0.00285f
C344 VCC.n369 VSS 0.00285f
C345 VCC.n371 VSS 0.00285f
C346 VCC.n372 VSS 0.00285f
C347 VCC.n373 VSS 0.00285f
C348 VCC.n374 VSS 0.00285f
C349 VCC.n375 VSS 0.00285f
C350 VCC.n377 VSS 0.00285f
C351 VCC.n379 VSS 0.00285f
C352 VCC.n380 VSS 0.00285f
C353 VCC.n381 VSS 0.00285f
C354 VCC.n382 VSS 0.00285f
C355 VCC.n383 VSS 0.00285f
C356 VCC.n385 VSS 0.00285f
C357 VCC.n387 VSS 0.00285f
C358 VCC.n388 VSS 0.00285f
C359 VCC.n389 VSS 0.00285f
C360 VCC.n390 VSS 0.00285f
C361 VCC.n391 VSS 0.00285f
C362 VCC.n393 VSS 0.00285f
C363 VCC.n395 VSS 0.00285f
C364 VCC.n396 VSS 0.00285f
C365 VCC.n397 VSS 0.00285f
C366 VCC.n398 VSS 0.00285f
C367 VCC.n399 VSS 0.00285f
C368 VCC.n401 VSS 0.00285f
C369 VCC.n403 VSS 0.00285f
C370 VCC.n404 VSS 0.00285f
C371 VCC.n405 VSS 0.00285f
C372 VCC.n406 VSS 0.00285f
C373 VCC.n407 VSS 0.00285f
C374 VCC.n409 VSS 0.00285f
C375 VCC.n411 VSS 0.00285f
C376 VCC.n412 VSS 0.00285f
C377 VCC.n413 VSS 0.00285f
C378 VCC.n414 VSS 0.00285f
C379 VCC.n415 VSS 0.00285f
C380 VCC.n417 VSS 0.00285f
C381 VCC.n419 VSS 0.00285f
C382 VCC.n420 VSS 0.00285f
C383 VCC.n421 VSS 0.00285f
C384 VCC.n422 VSS 0.00285f
C385 VCC.n423 VSS 0.00285f
C386 VCC.n425 VSS 0.00285f
C387 VCC.n427 VSS 0.00285f
C388 VCC.n428 VSS 0.00285f
C389 VCC.n429 VSS 0.00285f
C390 VCC.n430 VSS 0.00285f
C391 VCC.n431 VSS 0.00285f
C392 VCC.n433 VSS 0.00285f
C393 VCC.n435 VSS 0.00285f
C394 VCC.n436 VSS 0.00285f
C395 VCC.n437 VSS 0.00285f
C396 VCC.n438 VSS 0.00285f
C397 VCC.n439 VSS 0.00285f
C398 VCC.n441 VSS 0.00285f
C399 VCC.n443 VSS 0.00285f
C400 VCC.n444 VSS 0.00285f
C401 VCC.n445 VSS 0.00285f
C402 VCC.n446 VSS 0.00285f
C403 VCC.n447 VSS 0.00285f
C404 VCC.n449 VSS 0.00285f
C405 VCC.n451 VSS 0.00285f
C406 VCC.n452 VSS 0.00285f
C407 VCC.n453 VSS 0.002745f
C408 VCC.n454 VSS 0.005288f
C409 VCC.n455 VSS 0.00153f
C410 VCC.n456 VSS 0.00285f
C411 VCC.n458 VSS 0.00285f
C412 VCC.n460 VSS 0.00285f
C413 VCC.n461 VSS 0.00285f
C414 VCC.n462 VSS 0.00285f
C415 VCC.n463 VSS 0.00285f
C416 VCC.n464 VSS 0.00285f
C417 VCC.n466 VSS 0.00285f
C418 VCC.n468 VSS 0.00285f
C419 VCC.n469 VSS 0.00285f
C420 VCC.n470 VSS 0.00285f
C421 VCC.n471 VSS 0.00285f
C422 VCC.n472 VSS 0.00285f
C423 VCC.n474 VSS 0.00285f
C424 VCC.n476 VSS 0.00285f
C425 VCC.n477 VSS 0.00285f
C426 VCC.n478 VSS 0.00285f
C427 VCC.n479 VSS 0.00285f
C428 VCC.n480 VSS 0.00285f
C429 VCC.n482 VSS 0.00285f
C430 VCC.n484 VSS 0.00285f
C431 VCC.n485 VSS 0.00285f
C432 VCC.n486 VSS 0.00285f
C433 VCC.n487 VSS 0.00285f
C434 VCC.n488 VSS 0.00285f
C435 VCC.n490 VSS 0.00285f
C436 VCC.n492 VSS 0.00285f
C437 VCC.n493 VSS 0.00285f
C438 VCC.n494 VSS 0.00285f
C439 VCC.n495 VSS 0.00285f
C440 VCC.n496 VSS 0.00285f
C441 VCC.n498 VSS 0.00285f
C442 VCC.n500 VSS 0.00285f
C443 VCC.n501 VSS 0.00285f
C444 VCC.n502 VSS 0.00285f
C445 VCC.n503 VSS 0.00285f
C446 VCC.n504 VSS 0.00285f
C447 VCC.n506 VSS 0.00285f
C448 VCC.n508 VSS 0.00285f
C449 VCC.n509 VSS 0.00285f
C450 VCC.n510 VSS 0.00285f
C451 VCC.n511 VSS 0.00285f
C452 VCC.n512 VSS 0.00285f
C453 VCC.n514 VSS 0.00285f
C454 VCC.n516 VSS 0.00285f
C455 VCC.n517 VSS 0.00285f
C456 VCC.n518 VSS 0.00285f
C457 VCC.n519 VSS 0.00285f
C458 VCC.n520 VSS 0.00285f
C459 VCC.n522 VSS 0.00285f
C460 VCC.n524 VSS 0.00285f
C461 VCC.n525 VSS 0.00285f
C462 VCC.n526 VSS 0.00285f
C463 VCC.n527 VSS 0.00285f
C464 VCC.n528 VSS 0.00285f
C465 VCC.n530 VSS 0.00285f
C466 VCC.n532 VSS 0.00285f
C467 VCC.n533 VSS 0.00285f
C468 VCC.n534 VSS 0.00285f
C469 VCC.n535 VSS 0.00285f
C470 VCC.n536 VSS 0.00285f
C471 VCC.n538 VSS 0.00285f
C472 VCC.n540 VSS 0.00285f
C473 VCC.n541 VSS 0.00285f
C474 VCC.n542 VSS 0.005738f
C475 VCC.n543 VSS 0.014004f
C476 VCC.n544 VSS 0.0028f
C477 VCC.n545 VSS 0.008247f
C478 VCC.n546 VSS 0.458293f
C479 VCC.n547 VSS 0.008247f
C480 VCC.n548 VSS 0.0028f
C481 VCC.n549 VSS 0.003374f
C482 VCC.n550 VSS 0.004192f
C483 VCC.n551 VSS 0.004192f
C484 VCC.n552 VSS 0.004192f
C485 VCC.n553 VSS 0.003374f
C486 VCC.n554 VSS 0.003374f
C487 VCC.n555 VSS 0.003374f
C488 VOUT.t7 VSS 0.020098f
C489 VOUT.n0 VSS 0.017266f
C490 VOUT.t26 VSS 0.020098f
C491 VOUT.t15 VSS 0.017996f
C492 VOUT.n1 VSS 0.013634f
C493 VOUT.n2 VSS 0.017247f
C494 VOUT.n3 VSS 0.027601f
C495 VOUT.n4 VSS 0.062912f
C496 VOUT.n5 VSS 0.006713f
C497 VOUT.n6 VSS 0.015735f
C498 VOUT.t9 VSS 0.011196f
C499 VOUT.n7 VSS 0.011604f
C500 VOUT.n8 VSS 0.003288f
C501 VOUT.n9 VSS 0.002669f
C502 VOUT.n10 VSS 0.030873f
C503 VOUT.n11 VSS 0.007359f
C504 VOUT.n12 VSS 0.031452f
C505 VOUT.t27 VSS 0.018417f
C506 VOUT.t8 VSS 0.007221f
C507 VOUT.n13 VSS 0.006713f
C508 VOUT.n14 VSS 0.015735f
C509 VOUT.n15 VSS 0.011604f
C510 VOUT.n16 VSS 0.003288f
C511 VOUT.n17 VSS 0.002669f
C512 VOUT.n18 VSS 0.030873f
C513 VOUT.n19 VSS 0.010958f
C514 VOUT.n20 VSS 0.135637f
C515 VOUT.n21 VSS 0.121527f
C516 VOUT.t20 VSS 0.066363f
C517 VOUT.n22 VSS 0.005352f
C518 VOUT.n23 VSS 0.004966f
C519 VOUT.n24 VSS 0.002669f
C520 VOUT.n25 VSS 0.006308f
C521 VOUT.n26 VSS 0.002826f
C522 VOUT.n27 VSS 0.004966f
C523 VOUT.n28 VSS 0.002669f
C524 VOUT.n29 VSS 0.006308f
C525 VOUT.n30 VSS 0.002826f
C526 VOUT.n31 VSS 0.004966f
C527 VOUT.n32 VSS 0.002669f
C528 VOUT.n33 VSS 0.006308f
C529 VOUT.n34 VSS 0.002747f
C530 VOUT.n35 VSS 0.004966f
C531 VOUT.n36 VSS 0.002826f
C532 VOUT.n37 VSS 0.006308f
C533 VOUT.n38 VSS 0.002826f
C534 VOUT.n39 VSS 0.004966f
C535 VOUT.n40 VSS 0.002669f
C536 VOUT.n41 VSS 0.006308f
C537 VOUT.n42 VSS 0.002826f
C538 VOUT.n43 VSS 0.275351f
C539 VOUT.n44 VSS 0.002669f
C540 VOUT.n45 VSS 0.042346f
C541 VOUT.n46 VSS 0.004745f
C542 VOUT.n47 VSS 0.004731f
C543 VOUT.n48 VSS 0.006308f
C544 VOUT.n49 VSS 0.002826f
C545 VOUT.n50 VSS 0.002669f
C546 VOUT.n51 VSS 0.004966f
C547 VOUT.n52 VSS 0.004966f
C548 VOUT.n53 VSS 0.002669f
C549 VOUT.n54 VSS 0.002826f
C550 VOUT.n55 VSS 0.006308f
C551 VOUT.n56 VSS 0.006308f
C552 VOUT.n57 VSS 0.002826f
C553 VOUT.n58 VSS 0.002669f
C554 VOUT.n59 VSS 0.004966f
C555 VOUT.n60 VSS 0.004966f
C556 VOUT.n61 VSS 0.002669f
C557 VOUT.n62 VSS 0.002669f
C558 VOUT.n63 VSS 0.002826f
C559 VOUT.n64 VSS 0.006308f
C560 VOUT.n65 VSS 0.006308f
C561 VOUT.n66 VSS 0.006308f
C562 VOUT.n67 VSS 0.002747f
C563 VOUT.n68 VSS 0.002669f
C564 VOUT.n69 VSS 0.004966f
C565 VOUT.n70 VSS 0.004966f
C566 VOUT.n71 VSS 0.002669f
C567 VOUT.n72 VSS 0.002826f
C568 VOUT.n73 VSS 0.006308f
C569 VOUT.n74 VSS 0.006308f
C570 VOUT.n75 VSS 0.002826f
C571 VOUT.n76 VSS 0.002669f
C572 VOUT.n77 VSS 0.004966f
C573 VOUT.n78 VSS 0.004966f
C574 VOUT.n79 VSS 0.002669f
C575 VOUT.n80 VSS 0.002826f
C576 VOUT.n81 VSS 0.006308f
C577 VOUT.n82 VSS 0.006308f
C578 VOUT.n83 VSS 0.002826f
C579 VOUT.n84 VSS 0.002669f
C580 VOUT.n85 VSS 0.004966f
C581 VOUT.n86 VSS 0.004966f
C582 VOUT.n87 VSS 0.002669f
C583 VOUT.n88 VSS 0.002826f
C584 VOUT.n89 VSS 0.006308f
C585 VOUT.n90 VSS 0.014913f
C586 VOUT.n91 VSS 0.002826f
C587 VOUT.n92 VSS 0.002669f
C588 VOUT.n93 VSS 0.010665f
C589 VOUT.n94 VSS 0.011058f
C590 VOUT.n95 VSS 0.011058f
C591 VOUT.n96 VSS 0.042346f
C592 VOUT.n97 VSS 0.006308f
C593 VOUT.n98 VSS 0.002826f
C594 VOUT.n99 VSS 0.004966f
C595 VOUT.n100 VSS 0.002669f
C596 VOUT.n101 VSS 0.006308f
C597 VOUT.n102 VSS 0.002826f
C598 VOUT.n103 VSS 0.004966f
C599 VOUT.n104 VSS 0.002669f
C600 VOUT.n105 VSS 0.006308f
C601 VOUT.n106 VSS 0.002826f
C602 VOUT.n107 VSS 0.004966f
C603 VOUT.n108 VSS 0.002747f
C604 VOUT.n109 VSS 0.006308f
C605 VOUT.n110 VSS 0.002669f
C606 VOUT.n111 VSS 0.002826f
C607 VOUT.n112 VSS 0.004966f
C608 VOUT.n113 VSS 0.002669f
C609 VOUT.n114 VSS 0.006308f
C610 VOUT.n115 VSS 0.002826f
C611 VOUT.n116 VSS 0.004966f
C612 VOUT.n117 VSS 0.002669f
C613 VOUT.n118 VSS 0.014913f
C614 VOUT.n119 VSS 0.002826f
C615 VOUT.n120 VSS 0.005352f
C616 VOUT.n121 VSS 0.002669f
C617 VOUT.n122 VSS 0.010665f
C618 VOUT.n123 VSS 0.004966f
C619 VOUT.n124 VSS 0.002669f
C620 VOUT.n125 VSS 0.002826f
C621 VOUT.n126 VSS 0.006308f
C622 VOUT.n127 VSS 0.006308f
C623 VOUT.n128 VSS 0.002826f
C624 VOUT.n129 VSS 0.002669f
C625 VOUT.n130 VSS 0.004966f
C626 VOUT.n131 VSS 0.004966f
C627 VOUT.n132 VSS 0.002669f
C628 VOUT.n133 VSS 0.002826f
C629 VOUT.n134 VSS 0.006308f
C630 VOUT.n135 VSS 0.006308f
C631 VOUT.n136 VSS 0.002826f
C632 VOUT.n137 VSS 0.002669f
C633 VOUT.n138 VSS 0.004966f
C634 VOUT.n139 VSS 0.004966f
C635 VOUT.n140 VSS 0.002669f
C636 VOUT.n141 VSS 0.002826f
C637 VOUT.n142 VSS 0.006308f
C638 VOUT.n143 VSS 0.006308f
C639 VOUT.n144 VSS 0.006308f
C640 VOUT.n145 VSS 0.002747f
C641 VOUT.n146 VSS 0.002669f
C642 VOUT.n147 VSS 0.004966f
C643 VOUT.n148 VSS 0.004966f
C644 VOUT.n149 VSS 0.002669f
C645 VOUT.n150 VSS 0.002826f
C646 VOUT.n151 VSS 0.006308f
C647 VOUT.n152 VSS 0.006308f
C648 VOUT.n153 VSS 0.002826f
C649 VOUT.n154 VSS 0.002669f
C650 VOUT.n155 VSS 0.004966f
C651 VOUT.n156 VSS 0.004966f
C652 VOUT.n157 VSS 0.002669f
C653 VOUT.n158 VSS 0.002826f
C654 VOUT.n159 VSS 0.006308f
C655 VOUT.n160 VSS 0.006308f
C656 VOUT.n161 VSS 0.002826f
C657 VOUT.n162 VSS 0.002669f
C658 VOUT.n163 VSS 0.004966f
C659 VOUT.n164 VSS 0.275351f
C660 VOUT.n165 VSS 0.002669f
C661 VOUT.n166 VSS 0.004745f
C662 VOUT.n167 VSS 0.004731f
C663 VOUT.t14 VSS 0.066363f
C664 VOUT.t0 VSS 0.102442f
C665 VOUT.n168 VSS 0.044297f
C666 VOUT.t13 VSS 0.102442f
C667 VOUT.t17 VSS 0.101447f
C668 VOUT.n169 VSS 0.040737f
C669 VOUT.n170 VSS 0.044279f
C670 VOUT.n171 VSS 0.025837f
C671 VOUT.t21 VSS 0.020098f
C672 VOUT.n172 VSS 0.017266f
C673 VOUT.t24 VSS 0.020098f
C674 VOUT.t5 VSS 0.017996f
C675 VOUT.n173 VSS 0.013634f
C676 VOUT.n174 VSS 0.017247f
C677 VOUT.n175 VSS 0.049079f
C678 VOUT.n176 VSS 0.165647f
C679 VOUT.t10 VSS 0.102442f
C680 VOUT.n177 VSS 0.044297f
C681 VOUT.t19 VSS 0.102442f
C682 VOUT.t3 VSS 0.101447f
C683 VOUT.n178 VSS 0.040737f
C684 VOUT.n179 VSS 0.044279f
C685 VOUT.n180 VSS 0.046861f
C686 VOUT.n181 VSS 0.167564f
C687 VOUT.n182 VSS 0.189639f
C688 VOUT.n183 VSS 0.005352f
C689 VOUT.n184 VSS 0.004966f
C690 VOUT.n185 VSS 0.002669f
C691 VOUT.n186 VSS 0.006308f
C692 VOUT.n187 VSS 0.002826f
C693 VOUT.n188 VSS 0.004966f
C694 VOUT.n189 VSS 0.002669f
C695 VOUT.n190 VSS 0.006308f
C696 VOUT.n191 VSS 0.002826f
C697 VOUT.n192 VSS 0.004966f
C698 VOUT.n193 VSS 0.002669f
C699 VOUT.n194 VSS 0.006308f
C700 VOUT.n195 VSS 0.002747f
C701 VOUT.n196 VSS 0.004966f
C702 VOUT.n197 VSS 0.002826f
C703 VOUT.n198 VSS 0.006308f
C704 VOUT.n199 VSS 0.002826f
C705 VOUT.n200 VSS 0.004966f
C706 VOUT.n201 VSS 0.002669f
C707 VOUT.n202 VSS 0.006308f
C708 VOUT.n203 VSS 0.002826f
C709 VOUT.n204 VSS 0.275351f
C710 VOUT.n205 VSS 0.002669f
C711 VOUT.t2 VSS 0.013616f
C712 VOUT.n206 VSS 0.042346f
C713 VOUT.n207 VSS 0.004745f
C714 VOUT.n208 VSS 0.004731f
C715 VOUT.n209 VSS 0.006308f
C716 VOUT.n210 VSS 0.002826f
C717 VOUT.n211 VSS 0.002669f
C718 VOUT.n212 VSS 0.004966f
C719 VOUT.n213 VSS 0.004966f
C720 VOUT.n214 VSS 0.002669f
C721 VOUT.n215 VSS 0.002826f
C722 VOUT.n216 VSS 0.006308f
C723 VOUT.n217 VSS 0.006308f
C724 VOUT.n218 VSS 0.002826f
C725 VOUT.n219 VSS 0.002669f
C726 VOUT.n220 VSS 0.004966f
C727 VOUT.n221 VSS 0.004966f
C728 VOUT.n222 VSS 0.002669f
C729 VOUT.n223 VSS 0.002669f
C730 VOUT.n224 VSS 0.002826f
C731 VOUT.n225 VSS 0.006308f
C732 VOUT.n226 VSS 0.006308f
C733 VOUT.n227 VSS 0.006308f
C734 VOUT.n228 VSS 0.002747f
C735 VOUT.n229 VSS 0.002669f
C736 VOUT.n230 VSS 0.004966f
C737 VOUT.n231 VSS 0.004966f
C738 VOUT.n232 VSS 0.002669f
C739 VOUT.n233 VSS 0.002826f
C740 VOUT.n234 VSS 0.006308f
C741 VOUT.n235 VSS 0.006308f
C742 VOUT.n236 VSS 0.002826f
C743 VOUT.n237 VSS 0.002669f
C744 VOUT.n238 VSS 0.004966f
C745 VOUT.n239 VSS 0.004966f
C746 VOUT.n240 VSS 0.002669f
C747 VOUT.n241 VSS 0.002826f
C748 VOUT.n242 VSS 0.006308f
C749 VOUT.n243 VSS 0.006308f
C750 VOUT.n244 VSS 0.002826f
C751 VOUT.n245 VSS 0.002669f
C752 VOUT.n246 VSS 0.004966f
C753 VOUT.n247 VSS 0.004966f
C754 VOUT.n248 VSS 0.002669f
C755 VOUT.n249 VSS 0.002826f
C756 VOUT.n250 VSS 0.006308f
C757 VOUT.n251 VSS 0.014913f
C758 VOUT.n252 VSS 0.002826f
C759 VOUT.n253 VSS 0.002669f
C760 VOUT.n254 VSS 0.010665f
C761 VOUT.n255 VSS 0.007458f
C762 VOUT.n256 VSS 0.029699f
C763 VOUT.n257 VSS 0.152048f
C764 VOUT.n258 VSS 0.387121f
C765 VOUT.t18 VSS 0.105493f
C766 VOUT.t1 VSS 0.052746f
C767 VOUT.n259 VSS 0.417273f
C768 VOUT.n260 VSS 0.126743f
C769 VOUT.n261 VSS 0.149983f
C770 VOUT.n262 VSS 0.272567f
C771 VOUT.t11 VSS 0.052746f
C772 VOUT.n263 VSS 0.417273f
C773 VOUT.t4 VSS 0.105493f
C774 VOUT.n264 VSS 0.388313f
C775 VOUT.n265 VSS 0.005352f
C776 VOUT.n266 VSS 0.004966f
C777 VOUT.n267 VSS 0.002669f
C778 VOUT.n268 VSS 0.006308f
C779 VOUT.n269 VSS 0.002826f
C780 VOUT.n270 VSS 0.004966f
C781 VOUT.n271 VSS 0.002669f
C782 VOUT.n272 VSS 0.006308f
C783 VOUT.n273 VSS 0.002826f
C784 VOUT.n274 VSS 0.004966f
C785 VOUT.n275 VSS 0.002669f
C786 VOUT.n276 VSS 0.006308f
C787 VOUT.n277 VSS 0.002747f
C788 VOUT.n278 VSS 0.004966f
C789 VOUT.n279 VSS 0.002826f
C790 VOUT.n280 VSS 0.006308f
C791 VOUT.n281 VSS 0.002826f
C792 VOUT.n282 VSS 0.004966f
C793 VOUT.n283 VSS 0.002669f
C794 VOUT.n284 VSS 0.006308f
C795 VOUT.n285 VSS 0.002826f
C796 VOUT.n286 VSS 0.275351f
C797 VOUT.n287 VSS 0.002669f
C798 VOUT.t12 VSS 0.013616f
C799 VOUT.n288 VSS 0.042346f
C800 VOUT.n289 VSS 0.004745f
C801 VOUT.n290 VSS 0.004731f
C802 VOUT.n291 VSS 0.006308f
C803 VOUT.n292 VSS 0.002826f
C804 VOUT.n293 VSS 0.002669f
C805 VOUT.n294 VSS 0.004966f
C806 VOUT.n295 VSS 0.004966f
C807 VOUT.n296 VSS 0.002669f
C808 VOUT.n297 VSS 0.002826f
C809 VOUT.n298 VSS 0.006308f
C810 VOUT.n299 VSS 0.006308f
C811 VOUT.n300 VSS 0.002826f
C812 VOUT.n301 VSS 0.002669f
C813 VOUT.n302 VSS 0.004966f
C814 VOUT.n303 VSS 0.004966f
C815 VOUT.n304 VSS 0.002669f
C816 VOUT.n305 VSS 0.002669f
C817 VOUT.n306 VSS 0.002826f
C818 VOUT.n307 VSS 0.006308f
C819 VOUT.n308 VSS 0.006308f
C820 VOUT.n309 VSS 0.006308f
C821 VOUT.n310 VSS 0.002747f
C822 VOUT.n311 VSS 0.002669f
C823 VOUT.n312 VSS 0.004966f
C824 VOUT.n313 VSS 0.004966f
C825 VOUT.n314 VSS 0.002669f
C826 VOUT.n315 VSS 0.002826f
C827 VOUT.n316 VSS 0.006308f
C828 VOUT.n317 VSS 0.006308f
C829 VOUT.n318 VSS 0.002826f
C830 VOUT.n319 VSS 0.002669f
C831 VOUT.n320 VSS 0.004966f
C832 VOUT.n321 VSS 0.004966f
C833 VOUT.n322 VSS 0.002669f
C834 VOUT.n323 VSS 0.002826f
C835 VOUT.n324 VSS 0.006308f
C836 VOUT.n325 VSS 0.006308f
C837 VOUT.n326 VSS 0.002826f
C838 VOUT.n327 VSS 0.002669f
C839 VOUT.n328 VSS 0.004966f
C840 VOUT.n329 VSS 0.004966f
C841 VOUT.n330 VSS 0.002669f
C842 VOUT.n331 VSS 0.002826f
C843 VOUT.n332 VSS 0.006308f
C844 VOUT.n333 VSS 0.014913f
C845 VOUT.n334 VSS 0.002826f
C846 VOUT.n335 VSS 0.002669f
C847 VOUT.n336 VSS 0.010665f
C848 VOUT.n337 VSS 0.007458f
C849 VOUT.n338 VSS 0.165669f
C850 VOUT.n339 VSS 0.136172f
C851 VOUT.n340 VSS 0.011604f
C852 VOUT.n341 VSS 0.030873f
C853 VOUT.n342 VSS 0.010958f
C854 VOUT.n343 VSS 0.006713f
C855 VOUT.n344 VSS 0.002669f
C856 VOUT.n345 VSS 0.003288f
C857 VOUT.n346 VSS 0.015735f
C858 VOUT.t25 VSS 0.018417f
C859 VOUT.t22 VSS 0.007221f
C860 VOUT.n347 VSS 0.04631f
C861 VOUT.t6 VSS 0.014443f
C862 VOUT.n348 VSS 0.040003f
C863 VOUT.n349 VSS 0.006713f
C864 VOUT.n350 VSS 0.015735f
C865 VOUT.t23 VSS 0.011196f
C866 VOUT.n351 VSS 0.011604f
C867 VOUT.n352 VSS 0.003288f
C868 VOUT.n353 VSS 0.002669f
C869 VOUT.n354 VSS 0.030873f
C870 VOUT.n355 VSS 0.007359f
C871 VOUT.n356 VSS 0.083941f
C872 VOUT.n357 VSS 0.064266f
C873 VOUT.n358 VSS 0.049509f
C874 VOUT.n359 VSS 0.074663f
C875 VOUT.n360 VSS 0.07097f
C876 VOUT.n361 VSS 0.04631f
C877 VOUT.t16 VSS 0.014443f
C878 VOUT.n362 VSS 0.03969f
C879 VOUT.n363 VSS 0.047186f
.ends

