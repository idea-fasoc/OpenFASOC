* NGSPICE file created from diff_pair_sample_1238.ext - technology: sky130A

.subckt diff_pair_sample_1238 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=3.74
X1 VTAIL.t19 VP.t0 VDD1.t1 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X2 VDD1.t2 VP.t1 VTAIL.t18 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=3.74
X3 VDD2.t9 VN.t0 VTAIL.t2 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=3.74
X4 VDD2.t8 VN.t1 VTAIL.t7 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X5 VTAIL.t17 VP.t2 VDD1.t3 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X6 VDD1.t0 VP.t3 VTAIL.t16 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=3.74
X7 VTAIL.t15 VP.t4 VDD1.t4 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X8 VDD2.t7 VN.t2 VTAIL.t4 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=3.74
X9 VTAIL.t1 VN.t3 VDD2.t6 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X10 VDD2.t5 VN.t4 VTAIL.t0 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=3.74
X11 VTAIL.t3 VN.t5 VDD2.t4 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X12 VTAIL.t9 VN.t6 VDD2.t3 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X13 VDD1.t5 VP.t5 VTAIL.t14 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X14 B.t8 B.t6 B.t7 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=3.74
X15 VDD2.t2 VN.t7 VTAIL.t5 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X16 VDD2.t1 VN.t8 VTAIL.t8 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=3.74
X17 VDD1.t8 VP.t6 VTAIL.t13 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X18 VDD1.t7 VP.t7 VTAIL.t12 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=3.74
X19 VTAIL.t6 VN.t9 VDD2.t0 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X20 B.t5 B.t3 B.t4 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=3.74
X21 B.t2 B.t0 B.t1 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=3.74
X22 VTAIL.t11 VP.t8 VDD1.t9 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=3.74
X23 VDD1.t6 VP.t9 VTAIL.t10 w_n5854_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=3.74
R0 B.n845 B.n108 585
R1 B.n847 B.n846 585
R2 B.n848 B.n107 585
R3 B.n850 B.n849 585
R4 B.n851 B.n106 585
R5 B.n853 B.n852 585
R6 B.n854 B.n105 585
R7 B.n856 B.n855 585
R8 B.n857 B.n104 585
R9 B.n859 B.n858 585
R10 B.n860 B.n103 585
R11 B.n862 B.n861 585
R12 B.n863 B.n102 585
R13 B.n865 B.n864 585
R14 B.n866 B.n101 585
R15 B.n868 B.n867 585
R16 B.n869 B.n100 585
R17 B.n871 B.n870 585
R18 B.n872 B.n99 585
R19 B.n874 B.n873 585
R20 B.n875 B.n98 585
R21 B.n877 B.n876 585
R22 B.n878 B.n97 585
R23 B.n880 B.n879 585
R24 B.n881 B.n96 585
R25 B.n883 B.n882 585
R26 B.n884 B.n95 585
R27 B.n886 B.n885 585
R28 B.n887 B.n94 585
R29 B.n889 B.n888 585
R30 B.n890 B.n93 585
R31 B.n892 B.n891 585
R32 B.n893 B.n92 585
R33 B.n895 B.n894 585
R34 B.n896 B.n91 585
R35 B.n898 B.n897 585
R36 B.n899 B.n90 585
R37 B.n901 B.n900 585
R38 B.n902 B.n89 585
R39 B.n904 B.n903 585
R40 B.n905 B.n88 585
R41 B.n907 B.n906 585
R42 B.n908 B.n87 585
R43 B.n910 B.n909 585
R44 B.n911 B.n86 585
R45 B.n913 B.n912 585
R46 B.n914 B.n85 585
R47 B.n916 B.n915 585
R48 B.n917 B.n84 585
R49 B.n919 B.n918 585
R50 B.n920 B.n83 585
R51 B.n922 B.n921 585
R52 B.n923 B.n82 585
R53 B.n925 B.n924 585
R54 B.n926 B.n81 585
R55 B.n928 B.n927 585
R56 B.n929 B.n80 585
R57 B.n931 B.n930 585
R58 B.n933 B.n77 585
R59 B.n935 B.n934 585
R60 B.n936 B.n76 585
R61 B.n938 B.n937 585
R62 B.n939 B.n75 585
R63 B.n941 B.n940 585
R64 B.n942 B.n74 585
R65 B.n944 B.n943 585
R66 B.n945 B.n71 585
R67 B.n948 B.n947 585
R68 B.n949 B.n70 585
R69 B.n951 B.n950 585
R70 B.n952 B.n69 585
R71 B.n954 B.n953 585
R72 B.n955 B.n68 585
R73 B.n957 B.n956 585
R74 B.n958 B.n67 585
R75 B.n960 B.n959 585
R76 B.n961 B.n66 585
R77 B.n963 B.n962 585
R78 B.n964 B.n65 585
R79 B.n966 B.n965 585
R80 B.n967 B.n64 585
R81 B.n969 B.n968 585
R82 B.n970 B.n63 585
R83 B.n972 B.n971 585
R84 B.n973 B.n62 585
R85 B.n975 B.n974 585
R86 B.n976 B.n61 585
R87 B.n978 B.n977 585
R88 B.n979 B.n60 585
R89 B.n981 B.n980 585
R90 B.n982 B.n59 585
R91 B.n984 B.n983 585
R92 B.n985 B.n58 585
R93 B.n987 B.n986 585
R94 B.n988 B.n57 585
R95 B.n990 B.n989 585
R96 B.n991 B.n56 585
R97 B.n993 B.n992 585
R98 B.n994 B.n55 585
R99 B.n996 B.n995 585
R100 B.n997 B.n54 585
R101 B.n999 B.n998 585
R102 B.n1000 B.n53 585
R103 B.n1002 B.n1001 585
R104 B.n1003 B.n52 585
R105 B.n1005 B.n1004 585
R106 B.n1006 B.n51 585
R107 B.n1008 B.n1007 585
R108 B.n1009 B.n50 585
R109 B.n1011 B.n1010 585
R110 B.n1012 B.n49 585
R111 B.n1014 B.n1013 585
R112 B.n1015 B.n48 585
R113 B.n1017 B.n1016 585
R114 B.n1018 B.n47 585
R115 B.n1020 B.n1019 585
R116 B.n1021 B.n46 585
R117 B.n1023 B.n1022 585
R118 B.n1024 B.n45 585
R119 B.n1026 B.n1025 585
R120 B.n1027 B.n44 585
R121 B.n1029 B.n1028 585
R122 B.n1030 B.n43 585
R123 B.n1032 B.n1031 585
R124 B.n1033 B.n42 585
R125 B.n844 B.n843 585
R126 B.n842 B.n109 585
R127 B.n841 B.n840 585
R128 B.n839 B.n110 585
R129 B.n838 B.n837 585
R130 B.n836 B.n111 585
R131 B.n835 B.n834 585
R132 B.n833 B.n112 585
R133 B.n832 B.n831 585
R134 B.n830 B.n113 585
R135 B.n829 B.n828 585
R136 B.n827 B.n114 585
R137 B.n826 B.n825 585
R138 B.n824 B.n115 585
R139 B.n823 B.n822 585
R140 B.n821 B.n116 585
R141 B.n820 B.n819 585
R142 B.n818 B.n117 585
R143 B.n817 B.n816 585
R144 B.n815 B.n118 585
R145 B.n814 B.n813 585
R146 B.n812 B.n119 585
R147 B.n811 B.n810 585
R148 B.n809 B.n120 585
R149 B.n808 B.n807 585
R150 B.n806 B.n121 585
R151 B.n805 B.n804 585
R152 B.n803 B.n122 585
R153 B.n802 B.n801 585
R154 B.n800 B.n123 585
R155 B.n799 B.n798 585
R156 B.n797 B.n124 585
R157 B.n796 B.n795 585
R158 B.n794 B.n125 585
R159 B.n793 B.n792 585
R160 B.n791 B.n126 585
R161 B.n790 B.n789 585
R162 B.n788 B.n127 585
R163 B.n787 B.n786 585
R164 B.n785 B.n128 585
R165 B.n784 B.n783 585
R166 B.n782 B.n129 585
R167 B.n781 B.n780 585
R168 B.n779 B.n130 585
R169 B.n778 B.n777 585
R170 B.n776 B.n131 585
R171 B.n775 B.n774 585
R172 B.n773 B.n132 585
R173 B.n772 B.n771 585
R174 B.n770 B.n133 585
R175 B.n769 B.n768 585
R176 B.n767 B.n134 585
R177 B.n766 B.n765 585
R178 B.n764 B.n135 585
R179 B.n763 B.n762 585
R180 B.n761 B.n136 585
R181 B.n760 B.n759 585
R182 B.n758 B.n137 585
R183 B.n757 B.n756 585
R184 B.n755 B.n138 585
R185 B.n754 B.n753 585
R186 B.n752 B.n139 585
R187 B.n751 B.n750 585
R188 B.n749 B.n140 585
R189 B.n748 B.n747 585
R190 B.n746 B.n141 585
R191 B.n745 B.n744 585
R192 B.n743 B.n142 585
R193 B.n742 B.n741 585
R194 B.n740 B.n143 585
R195 B.n739 B.n738 585
R196 B.n737 B.n144 585
R197 B.n736 B.n735 585
R198 B.n734 B.n145 585
R199 B.n733 B.n732 585
R200 B.n731 B.n146 585
R201 B.n730 B.n729 585
R202 B.n728 B.n147 585
R203 B.n727 B.n726 585
R204 B.n725 B.n148 585
R205 B.n724 B.n723 585
R206 B.n722 B.n149 585
R207 B.n721 B.n720 585
R208 B.n719 B.n150 585
R209 B.n718 B.n717 585
R210 B.n716 B.n151 585
R211 B.n715 B.n714 585
R212 B.n713 B.n152 585
R213 B.n712 B.n711 585
R214 B.n710 B.n153 585
R215 B.n709 B.n708 585
R216 B.n707 B.n154 585
R217 B.n706 B.n705 585
R218 B.n704 B.n155 585
R219 B.n703 B.n702 585
R220 B.n701 B.n156 585
R221 B.n700 B.n699 585
R222 B.n698 B.n157 585
R223 B.n697 B.n696 585
R224 B.n695 B.n158 585
R225 B.n694 B.n693 585
R226 B.n692 B.n159 585
R227 B.n691 B.n690 585
R228 B.n689 B.n160 585
R229 B.n688 B.n687 585
R230 B.n686 B.n161 585
R231 B.n685 B.n684 585
R232 B.n683 B.n162 585
R233 B.n682 B.n681 585
R234 B.n680 B.n163 585
R235 B.n679 B.n678 585
R236 B.n677 B.n164 585
R237 B.n676 B.n675 585
R238 B.n674 B.n165 585
R239 B.n673 B.n672 585
R240 B.n671 B.n166 585
R241 B.n670 B.n669 585
R242 B.n668 B.n167 585
R243 B.n667 B.n666 585
R244 B.n665 B.n168 585
R245 B.n664 B.n663 585
R246 B.n662 B.n169 585
R247 B.n661 B.n660 585
R248 B.n659 B.n170 585
R249 B.n658 B.n657 585
R250 B.n656 B.n171 585
R251 B.n655 B.n654 585
R252 B.n653 B.n172 585
R253 B.n652 B.n651 585
R254 B.n650 B.n173 585
R255 B.n649 B.n648 585
R256 B.n647 B.n174 585
R257 B.n646 B.n645 585
R258 B.n644 B.n175 585
R259 B.n643 B.n642 585
R260 B.n641 B.n176 585
R261 B.n640 B.n639 585
R262 B.n638 B.n177 585
R263 B.n637 B.n636 585
R264 B.n635 B.n178 585
R265 B.n634 B.n633 585
R266 B.n632 B.n179 585
R267 B.n631 B.n630 585
R268 B.n629 B.n180 585
R269 B.n628 B.n627 585
R270 B.n626 B.n181 585
R271 B.n625 B.n624 585
R272 B.n623 B.n182 585
R273 B.n622 B.n621 585
R274 B.n620 B.n183 585
R275 B.n619 B.n618 585
R276 B.n617 B.n184 585
R277 B.n616 B.n615 585
R278 B.n614 B.n185 585
R279 B.n613 B.n612 585
R280 B.n611 B.n186 585
R281 B.n610 B.n609 585
R282 B.n608 B.n187 585
R283 B.n607 B.n606 585
R284 B.n605 B.n188 585
R285 B.n604 B.n603 585
R286 B.n415 B.n414 585
R287 B.n416 B.n255 585
R288 B.n418 B.n417 585
R289 B.n419 B.n254 585
R290 B.n421 B.n420 585
R291 B.n422 B.n253 585
R292 B.n424 B.n423 585
R293 B.n425 B.n252 585
R294 B.n427 B.n426 585
R295 B.n428 B.n251 585
R296 B.n430 B.n429 585
R297 B.n431 B.n250 585
R298 B.n433 B.n432 585
R299 B.n434 B.n249 585
R300 B.n436 B.n435 585
R301 B.n437 B.n248 585
R302 B.n439 B.n438 585
R303 B.n440 B.n247 585
R304 B.n442 B.n441 585
R305 B.n443 B.n246 585
R306 B.n445 B.n444 585
R307 B.n446 B.n245 585
R308 B.n448 B.n447 585
R309 B.n449 B.n244 585
R310 B.n451 B.n450 585
R311 B.n452 B.n243 585
R312 B.n454 B.n453 585
R313 B.n455 B.n242 585
R314 B.n457 B.n456 585
R315 B.n458 B.n241 585
R316 B.n460 B.n459 585
R317 B.n461 B.n240 585
R318 B.n463 B.n462 585
R319 B.n464 B.n239 585
R320 B.n466 B.n465 585
R321 B.n467 B.n238 585
R322 B.n469 B.n468 585
R323 B.n470 B.n237 585
R324 B.n472 B.n471 585
R325 B.n473 B.n236 585
R326 B.n475 B.n474 585
R327 B.n476 B.n235 585
R328 B.n478 B.n477 585
R329 B.n479 B.n234 585
R330 B.n481 B.n480 585
R331 B.n482 B.n233 585
R332 B.n484 B.n483 585
R333 B.n485 B.n232 585
R334 B.n487 B.n486 585
R335 B.n488 B.n231 585
R336 B.n490 B.n489 585
R337 B.n491 B.n230 585
R338 B.n493 B.n492 585
R339 B.n494 B.n229 585
R340 B.n496 B.n495 585
R341 B.n497 B.n228 585
R342 B.n499 B.n498 585
R343 B.n500 B.n225 585
R344 B.n503 B.n502 585
R345 B.n504 B.n224 585
R346 B.n506 B.n505 585
R347 B.n507 B.n223 585
R348 B.n509 B.n508 585
R349 B.n510 B.n222 585
R350 B.n512 B.n511 585
R351 B.n513 B.n221 585
R352 B.n515 B.n514 585
R353 B.n517 B.n516 585
R354 B.n518 B.n217 585
R355 B.n520 B.n519 585
R356 B.n521 B.n216 585
R357 B.n523 B.n522 585
R358 B.n524 B.n215 585
R359 B.n526 B.n525 585
R360 B.n527 B.n214 585
R361 B.n529 B.n528 585
R362 B.n530 B.n213 585
R363 B.n532 B.n531 585
R364 B.n533 B.n212 585
R365 B.n535 B.n534 585
R366 B.n536 B.n211 585
R367 B.n538 B.n537 585
R368 B.n539 B.n210 585
R369 B.n541 B.n540 585
R370 B.n542 B.n209 585
R371 B.n544 B.n543 585
R372 B.n545 B.n208 585
R373 B.n547 B.n546 585
R374 B.n548 B.n207 585
R375 B.n550 B.n549 585
R376 B.n551 B.n206 585
R377 B.n553 B.n552 585
R378 B.n554 B.n205 585
R379 B.n556 B.n555 585
R380 B.n557 B.n204 585
R381 B.n559 B.n558 585
R382 B.n560 B.n203 585
R383 B.n562 B.n561 585
R384 B.n563 B.n202 585
R385 B.n565 B.n564 585
R386 B.n566 B.n201 585
R387 B.n568 B.n567 585
R388 B.n569 B.n200 585
R389 B.n571 B.n570 585
R390 B.n572 B.n199 585
R391 B.n574 B.n573 585
R392 B.n575 B.n198 585
R393 B.n577 B.n576 585
R394 B.n578 B.n197 585
R395 B.n580 B.n579 585
R396 B.n581 B.n196 585
R397 B.n583 B.n582 585
R398 B.n584 B.n195 585
R399 B.n586 B.n585 585
R400 B.n587 B.n194 585
R401 B.n589 B.n588 585
R402 B.n590 B.n193 585
R403 B.n592 B.n591 585
R404 B.n593 B.n192 585
R405 B.n595 B.n594 585
R406 B.n596 B.n191 585
R407 B.n598 B.n597 585
R408 B.n599 B.n190 585
R409 B.n601 B.n600 585
R410 B.n602 B.n189 585
R411 B.n413 B.n256 585
R412 B.n412 B.n411 585
R413 B.n410 B.n257 585
R414 B.n409 B.n408 585
R415 B.n407 B.n258 585
R416 B.n406 B.n405 585
R417 B.n404 B.n259 585
R418 B.n403 B.n402 585
R419 B.n401 B.n260 585
R420 B.n400 B.n399 585
R421 B.n398 B.n261 585
R422 B.n397 B.n396 585
R423 B.n395 B.n262 585
R424 B.n394 B.n393 585
R425 B.n392 B.n263 585
R426 B.n391 B.n390 585
R427 B.n389 B.n264 585
R428 B.n388 B.n387 585
R429 B.n386 B.n265 585
R430 B.n385 B.n384 585
R431 B.n383 B.n266 585
R432 B.n382 B.n381 585
R433 B.n380 B.n267 585
R434 B.n379 B.n378 585
R435 B.n377 B.n268 585
R436 B.n376 B.n375 585
R437 B.n374 B.n269 585
R438 B.n373 B.n372 585
R439 B.n371 B.n270 585
R440 B.n370 B.n369 585
R441 B.n368 B.n271 585
R442 B.n367 B.n366 585
R443 B.n365 B.n272 585
R444 B.n364 B.n363 585
R445 B.n362 B.n273 585
R446 B.n361 B.n360 585
R447 B.n359 B.n274 585
R448 B.n358 B.n357 585
R449 B.n356 B.n275 585
R450 B.n355 B.n354 585
R451 B.n353 B.n276 585
R452 B.n352 B.n351 585
R453 B.n350 B.n277 585
R454 B.n349 B.n348 585
R455 B.n347 B.n278 585
R456 B.n346 B.n345 585
R457 B.n344 B.n279 585
R458 B.n343 B.n342 585
R459 B.n341 B.n280 585
R460 B.n340 B.n339 585
R461 B.n338 B.n281 585
R462 B.n337 B.n336 585
R463 B.n335 B.n282 585
R464 B.n334 B.n333 585
R465 B.n332 B.n283 585
R466 B.n331 B.n330 585
R467 B.n329 B.n284 585
R468 B.n328 B.n327 585
R469 B.n326 B.n285 585
R470 B.n325 B.n324 585
R471 B.n323 B.n286 585
R472 B.n322 B.n321 585
R473 B.n320 B.n287 585
R474 B.n319 B.n318 585
R475 B.n317 B.n288 585
R476 B.n316 B.n315 585
R477 B.n314 B.n289 585
R478 B.n313 B.n312 585
R479 B.n311 B.n290 585
R480 B.n310 B.n309 585
R481 B.n308 B.n291 585
R482 B.n307 B.n306 585
R483 B.n305 B.n292 585
R484 B.n304 B.n303 585
R485 B.n302 B.n293 585
R486 B.n301 B.n300 585
R487 B.n299 B.n294 585
R488 B.n298 B.n297 585
R489 B.n296 B.n295 585
R490 B.n2 B.n0 585
R491 B.n1153 B.n1 585
R492 B.n1152 B.n1151 585
R493 B.n1150 B.n3 585
R494 B.n1149 B.n1148 585
R495 B.n1147 B.n4 585
R496 B.n1146 B.n1145 585
R497 B.n1144 B.n5 585
R498 B.n1143 B.n1142 585
R499 B.n1141 B.n6 585
R500 B.n1140 B.n1139 585
R501 B.n1138 B.n7 585
R502 B.n1137 B.n1136 585
R503 B.n1135 B.n8 585
R504 B.n1134 B.n1133 585
R505 B.n1132 B.n9 585
R506 B.n1131 B.n1130 585
R507 B.n1129 B.n10 585
R508 B.n1128 B.n1127 585
R509 B.n1126 B.n11 585
R510 B.n1125 B.n1124 585
R511 B.n1123 B.n12 585
R512 B.n1122 B.n1121 585
R513 B.n1120 B.n13 585
R514 B.n1119 B.n1118 585
R515 B.n1117 B.n14 585
R516 B.n1116 B.n1115 585
R517 B.n1114 B.n15 585
R518 B.n1113 B.n1112 585
R519 B.n1111 B.n16 585
R520 B.n1110 B.n1109 585
R521 B.n1108 B.n17 585
R522 B.n1107 B.n1106 585
R523 B.n1105 B.n18 585
R524 B.n1104 B.n1103 585
R525 B.n1102 B.n19 585
R526 B.n1101 B.n1100 585
R527 B.n1099 B.n20 585
R528 B.n1098 B.n1097 585
R529 B.n1096 B.n21 585
R530 B.n1095 B.n1094 585
R531 B.n1093 B.n22 585
R532 B.n1092 B.n1091 585
R533 B.n1090 B.n23 585
R534 B.n1089 B.n1088 585
R535 B.n1087 B.n24 585
R536 B.n1086 B.n1085 585
R537 B.n1084 B.n25 585
R538 B.n1083 B.n1082 585
R539 B.n1081 B.n26 585
R540 B.n1080 B.n1079 585
R541 B.n1078 B.n27 585
R542 B.n1077 B.n1076 585
R543 B.n1075 B.n28 585
R544 B.n1074 B.n1073 585
R545 B.n1072 B.n29 585
R546 B.n1071 B.n1070 585
R547 B.n1069 B.n30 585
R548 B.n1068 B.n1067 585
R549 B.n1066 B.n31 585
R550 B.n1065 B.n1064 585
R551 B.n1063 B.n32 585
R552 B.n1062 B.n1061 585
R553 B.n1060 B.n33 585
R554 B.n1059 B.n1058 585
R555 B.n1057 B.n34 585
R556 B.n1056 B.n1055 585
R557 B.n1054 B.n35 585
R558 B.n1053 B.n1052 585
R559 B.n1051 B.n36 585
R560 B.n1050 B.n1049 585
R561 B.n1048 B.n37 585
R562 B.n1047 B.n1046 585
R563 B.n1045 B.n38 585
R564 B.n1044 B.n1043 585
R565 B.n1042 B.n39 585
R566 B.n1041 B.n1040 585
R567 B.n1039 B.n40 585
R568 B.n1038 B.n1037 585
R569 B.n1036 B.n41 585
R570 B.n1035 B.n1034 585
R571 B.n1155 B.n1154 585
R572 B.n218 B.t5 552.835
R573 B.n78 B.t10 552.835
R574 B.n226 B.t2 552.835
R575 B.n72 B.t7 552.835
R576 B.n414 B.n413 482.89
R577 B.n1034 B.n1033 482.89
R578 B.n604 B.n189 482.89
R579 B.n845 B.n844 482.89
R580 B.n219 B.t4 473.901
R581 B.n79 B.t11 473.901
R582 B.n227 B.t1 473.901
R583 B.n73 B.t8 473.901
R584 B.n218 B.t3 321.807
R585 B.n226 B.t0 321.807
R586 B.n72 B.t6 321.807
R587 B.n78 B.t9 321.807
R588 B.n413 B.n412 163.367
R589 B.n412 B.n257 163.367
R590 B.n408 B.n257 163.367
R591 B.n408 B.n407 163.367
R592 B.n407 B.n406 163.367
R593 B.n406 B.n259 163.367
R594 B.n402 B.n259 163.367
R595 B.n402 B.n401 163.367
R596 B.n401 B.n400 163.367
R597 B.n400 B.n261 163.367
R598 B.n396 B.n261 163.367
R599 B.n396 B.n395 163.367
R600 B.n395 B.n394 163.367
R601 B.n394 B.n263 163.367
R602 B.n390 B.n263 163.367
R603 B.n390 B.n389 163.367
R604 B.n389 B.n388 163.367
R605 B.n388 B.n265 163.367
R606 B.n384 B.n265 163.367
R607 B.n384 B.n383 163.367
R608 B.n383 B.n382 163.367
R609 B.n382 B.n267 163.367
R610 B.n378 B.n267 163.367
R611 B.n378 B.n377 163.367
R612 B.n377 B.n376 163.367
R613 B.n376 B.n269 163.367
R614 B.n372 B.n269 163.367
R615 B.n372 B.n371 163.367
R616 B.n371 B.n370 163.367
R617 B.n370 B.n271 163.367
R618 B.n366 B.n271 163.367
R619 B.n366 B.n365 163.367
R620 B.n365 B.n364 163.367
R621 B.n364 B.n273 163.367
R622 B.n360 B.n273 163.367
R623 B.n360 B.n359 163.367
R624 B.n359 B.n358 163.367
R625 B.n358 B.n275 163.367
R626 B.n354 B.n275 163.367
R627 B.n354 B.n353 163.367
R628 B.n353 B.n352 163.367
R629 B.n352 B.n277 163.367
R630 B.n348 B.n277 163.367
R631 B.n348 B.n347 163.367
R632 B.n347 B.n346 163.367
R633 B.n346 B.n279 163.367
R634 B.n342 B.n279 163.367
R635 B.n342 B.n341 163.367
R636 B.n341 B.n340 163.367
R637 B.n340 B.n281 163.367
R638 B.n336 B.n281 163.367
R639 B.n336 B.n335 163.367
R640 B.n335 B.n334 163.367
R641 B.n334 B.n283 163.367
R642 B.n330 B.n283 163.367
R643 B.n330 B.n329 163.367
R644 B.n329 B.n328 163.367
R645 B.n328 B.n285 163.367
R646 B.n324 B.n285 163.367
R647 B.n324 B.n323 163.367
R648 B.n323 B.n322 163.367
R649 B.n322 B.n287 163.367
R650 B.n318 B.n287 163.367
R651 B.n318 B.n317 163.367
R652 B.n317 B.n316 163.367
R653 B.n316 B.n289 163.367
R654 B.n312 B.n289 163.367
R655 B.n312 B.n311 163.367
R656 B.n311 B.n310 163.367
R657 B.n310 B.n291 163.367
R658 B.n306 B.n291 163.367
R659 B.n306 B.n305 163.367
R660 B.n305 B.n304 163.367
R661 B.n304 B.n293 163.367
R662 B.n300 B.n293 163.367
R663 B.n300 B.n299 163.367
R664 B.n299 B.n298 163.367
R665 B.n298 B.n295 163.367
R666 B.n295 B.n2 163.367
R667 B.n1154 B.n2 163.367
R668 B.n1154 B.n1153 163.367
R669 B.n1153 B.n1152 163.367
R670 B.n1152 B.n3 163.367
R671 B.n1148 B.n3 163.367
R672 B.n1148 B.n1147 163.367
R673 B.n1147 B.n1146 163.367
R674 B.n1146 B.n5 163.367
R675 B.n1142 B.n5 163.367
R676 B.n1142 B.n1141 163.367
R677 B.n1141 B.n1140 163.367
R678 B.n1140 B.n7 163.367
R679 B.n1136 B.n7 163.367
R680 B.n1136 B.n1135 163.367
R681 B.n1135 B.n1134 163.367
R682 B.n1134 B.n9 163.367
R683 B.n1130 B.n9 163.367
R684 B.n1130 B.n1129 163.367
R685 B.n1129 B.n1128 163.367
R686 B.n1128 B.n11 163.367
R687 B.n1124 B.n11 163.367
R688 B.n1124 B.n1123 163.367
R689 B.n1123 B.n1122 163.367
R690 B.n1122 B.n13 163.367
R691 B.n1118 B.n13 163.367
R692 B.n1118 B.n1117 163.367
R693 B.n1117 B.n1116 163.367
R694 B.n1116 B.n15 163.367
R695 B.n1112 B.n15 163.367
R696 B.n1112 B.n1111 163.367
R697 B.n1111 B.n1110 163.367
R698 B.n1110 B.n17 163.367
R699 B.n1106 B.n17 163.367
R700 B.n1106 B.n1105 163.367
R701 B.n1105 B.n1104 163.367
R702 B.n1104 B.n19 163.367
R703 B.n1100 B.n19 163.367
R704 B.n1100 B.n1099 163.367
R705 B.n1099 B.n1098 163.367
R706 B.n1098 B.n21 163.367
R707 B.n1094 B.n21 163.367
R708 B.n1094 B.n1093 163.367
R709 B.n1093 B.n1092 163.367
R710 B.n1092 B.n23 163.367
R711 B.n1088 B.n23 163.367
R712 B.n1088 B.n1087 163.367
R713 B.n1087 B.n1086 163.367
R714 B.n1086 B.n25 163.367
R715 B.n1082 B.n25 163.367
R716 B.n1082 B.n1081 163.367
R717 B.n1081 B.n1080 163.367
R718 B.n1080 B.n27 163.367
R719 B.n1076 B.n27 163.367
R720 B.n1076 B.n1075 163.367
R721 B.n1075 B.n1074 163.367
R722 B.n1074 B.n29 163.367
R723 B.n1070 B.n29 163.367
R724 B.n1070 B.n1069 163.367
R725 B.n1069 B.n1068 163.367
R726 B.n1068 B.n31 163.367
R727 B.n1064 B.n31 163.367
R728 B.n1064 B.n1063 163.367
R729 B.n1063 B.n1062 163.367
R730 B.n1062 B.n33 163.367
R731 B.n1058 B.n33 163.367
R732 B.n1058 B.n1057 163.367
R733 B.n1057 B.n1056 163.367
R734 B.n1056 B.n35 163.367
R735 B.n1052 B.n35 163.367
R736 B.n1052 B.n1051 163.367
R737 B.n1051 B.n1050 163.367
R738 B.n1050 B.n37 163.367
R739 B.n1046 B.n37 163.367
R740 B.n1046 B.n1045 163.367
R741 B.n1045 B.n1044 163.367
R742 B.n1044 B.n39 163.367
R743 B.n1040 B.n39 163.367
R744 B.n1040 B.n1039 163.367
R745 B.n1039 B.n1038 163.367
R746 B.n1038 B.n41 163.367
R747 B.n1034 B.n41 163.367
R748 B.n414 B.n255 163.367
R749 B.n418 B.n255 163.367
R750 B.n419 B.n418 163.367
R751 B.n420 B.n419 163.367
R752 B.n420 B.n253 163.367
R753 B.n424 B.n253 163.367
R754 B.n425 B.n424 163.367
R755 B.n426 B.n425 163.367
R756 B.n426 B.n251 163.367
R757 B.n430 B.n251 163.367
R758 B.n431 B.n430 163.367
R759 B.n432 B.n431 163.367
R760 B.n432 B.n249 163.367
R761 B.n436 B.n249 163.367
R762 B.n437 B.n436 163.367
R763 B.n438 B.n437 163.367
R764 B.n438 B.n247 163.367
R765 B.n442 B.n247 163.367
R766 B.n443 B.n442 163.367
R767 B.n444 B.n443 163.367
R768 B.n444 B.n245 163.367
R769 B.n448 B.n245 163.367
R770 B.n449 B.n448 163.367
R771 B.n450 B.n449 163.367
R772 B.n450 B.n243 163.367
R773 B.n454 B.n243 163.367
R774 B.n455 B.n454 163.367
R775 B.n456 B.n455 163.367
R776 B.n456 B.n241 163.367
R777 B.n460 B.n241 163.367
R778 B.n461 B.n460 163.367
R779 B.n462 B.n461 163.367
R780 B.n462 B.n239 163.367
R781 B.n466 B.n239 163.367
R782 B.n467 B.n466 163.367
R783 B.n468 B.n467 163.367
R784 B.n468 B.n237 163.367
R785 B.n472 B.n237 163.367
R786 B.n473 B.n472 163.367
R787 B.n474 B.n473 163.367
R788 B.n474 B.n235 163.367
R789 B.n478 B.n235 163.367
R790 B.n479 B.n478 163.367
R791 B.n480 B.n479 163.367
R792 B.n480 B.n233 163.367
R793 B.n484 B.n233 163.367
R794 B.n485 B.n484 163.367
R795 B.n486 B.n485 163.367
R796 B.n486 B.n231 163.367
R797 B.n490 B.n231 163.367
R798 B.n491 B.n490 163.367
R799 B.n492 B.n491 163.367
R800 B.n492 B.n229 163.367
R801 B.n496 B.n229 163.367
R802 B.n497 B.n496 163.367
R803 B.n498 B.n497 163.367
R804 B.n498 B.n225 163.367
R805 B.n503 B.n225 163.367
R806 B.n504 B.n503 163.367
R807 B.n505 B.n504 163.367
R808 B.n505 B.n223 163.367
R809 B.n509 B.n223 163.367
R810 B.n510 B.n509 163.367
R811 B.n511 B.n510 163.367
R812 B.n511 B.n221 163.367
R813 B.n515 B.n221 163.367
R814 B.n516 B.n515 163.367
R815 B.n516 B.n217 163.367
R816 B.n520 B.n217 163.367
R817 B.n521 B.n520 163.367
R818 B.n522 B.n521 163.367
R819 B.n522 B.n215 163.367
R820 B.n526 B.n215 163.367
R821 B.n527 B.n526 163.367
R822 B.n528 B.n527 163.367
R823 B.n528 B.n213 163.367
R824 B.n532 B.n213 163.367
R825 B.n533 B.n532 163.367
R826 B.n534 B.n533 163.367
R827 B.n534 B.n211 163.367
R828 B.n538 B.n211 163.367
R829 B.n539 B.n538 163.367
R830 B.n540 B.n539 163.367
R831 B.n540 B.n209 163.367
R832 B.n544 B.n209 163.367
R833 B.n545 B.n544 163.367
R834 B.n546 B.n545 163.367
R835 B.n546 B.n207 163.367
R836 B.n550 B.n207 163.367
R837 B.n551 B.n550 163.367
R838 B.n552 B.n551 163.367
R839 B.n552 B.n205 163.367
R840 B.n556 B.n205 163.367
R841 B.n557 B.n556 163.367
R842 B.n558 B.n557 163.367
R843 B.n558 B.n203 163.367
R844 B.n562 B.n203 163.367
R845 B.n563 B.n562 163.367
R846 B.n564 B.n563 163.367
R847 B.n564 B.n201 163.367
R848 B.n568 B.n201 163.367
R849 B.n569 B.n568 163.367
R850 B.n570 B.n569 163.367
R851 B.n570 B.n199 163.367
R852 B.n574 B.n199 163.367
R853 B.n575 B.n574 163.367
R854 B.n576 B.n575 163.367
R855 B.n576 B.n197 163.367
R856 B.n580 B.n197 163.367
R857 B.n581 B.n580 163.367
R858 B.n582 B.n581 163.367
R859 B.n582 B.n195 163.367
R860 B.n586 B.n195 163.367
R861 B.n587 B.n586 163.367
R862 B.n588 B.n587 163.367
R863 B.n588 B.n193 163.367
R864 B.n592 B.n193 163.367
R865 B.n593 B.n592 163.367
R866 B.n594 B.n593 163.367
R867 B.n594 B.n191 163.367
R868 B.n598 B.n191 163.367
R869 B.n599 B.n598 163.367
R870 B.n600 B.n599 163.367
R871 B.n600 B.n189 163.367
R872 B.n605 B.n604 163.367
R873 B.n606 B.n605 163.367
R874 B.n606 B.n187 163.367
R875 B.n610 B.n187 163.367
R876 B.n611 B.n610 163.367
R877 B.n612 B.n611 163.367
R878 B.n612 B.n185 163.367
R879 B.n616 B.n185 163.367
R880 B.n617 B.n616 163.367
R881 B.n618 B.n617 163.367
R882 B.n618 B.n183 163.367
R883 B.n622 B.n183 163.367
R884 B.n623 B.n622 163.367
R885 B.n624 B.n623 163.367
R886 B.n624 B.n181 163.367
R887 B.n628 B.n181 163.367
R888 B.n629 B.n628 163.367
R889 B.n630 B.n629 163.367
R890 B.n630 B.n179 163.367
R891 B.n634 B.n179 163.367
R892 B.n635 B.n634 163.367
R893 B.n636 B.n635 163.367
R894 B.n636 B.n177 163.367
R895 B.n640 B.n177 163.367
R896 B.n641 B.n640 163.367
R897 B.n642 B.n641 163.367
R898 B.n642 B.n175 163.367
R899 B.n646 B.n175 163.367
R900 B.n647 B.n646 163.367
R901 B.n648 B.n647 163.367
R902 B.n648 B.n173 163.367
R903 B.n652 B.n173 163.367
R904 B.n653 B.n652 163.367
R905 B.n654 B.n653 163.367
R906 B.n654 B.n171 163.367
R907 B.n658 B.n171 163.367
R908 B.n659 B.n658 163.367
R909 B.n660 B.n659 163.367
R910 B.n660 B.n169 163.367
R911 B.n664 B.n169 163.367
R912 B.n665 B.n664 163.367
R913 B.n666 B.n665 163.367
R914 B.n666 B.n167 163.367
R915 B.n670 B.n167 163.367
R916 B.n671 B.n670 163.367
R917 B.n672 B.n671 163.367
R918 B.n672 B.n165 163.367
R919 B.n676 B.n165 163.367
R920 B.n677 B.n676 163.367
R921 B.n678 B.n677 163.367
R922 B.n678 B.n163 163.367
R923 B.n682 B.n163 163.367
R924 B.n683 B.n682 163.367
R925 B.n684 B.n683 163.367
R926 B.n684 B.n161 163.367
R927 B.n688 B.n161 163.367
R928 B.n689 B.n688 163.367
R929 B.n690 B.n689 163.367
R930 B.n690 B.n159 163.367
R931 B.n694 B.n159 163.367
R932 B.n695 B.n694 163.367
R933 B.n696 B.n695 163.367
R934 B.n696 B.n157 163.367
R935 B.n700 B.n157 163.367
R936 B.n701 B.n700 163.367
R937 B.n702 B.n701 163.367
R938 B.n702 B.n155 163.367
R939 B.n706 B.n155 163.367
R940 B.n707 B.n706 163.367
R941 B.n708 B.n707 163.367
R942 B.n708 B.n153 163.367
R943 B.n712 B.n153 163.367
R944 B.n713 B.n712 163.367
R945 B.n714 B.n713 163.367
R946 B.n714 B.n151 163.367
R947 B.n718 B.n151 163.367
R948 B.n719 B.n718 163.367
R949 B.n720 B.n719 163.367
R950 B.n720 B.n149 163.367
R951 B.n724 B.n149 163.367
R952 B.n725 B.n724 163.367
R953 B.n726 B.n725 163.367
R954 B.n726 B.n147 163.367
R955 B.n730 B.n147 163.367
R956 B.n731 B.n730 163.367
R957 B.n732 B.n731 163.367
R958 B.n732 B.n145 163.367
R959 B.n736 B.n145 163.367
R960 B.n737 B.n736 163.367
R961 B.n738 B.n737 163.367
R962 B.n738 B.n143 163.367
R963 B.n742 B.n143 163.367
R964 B.n743 B.n742 163.367
R965 B.n744 B.n743 163.367
R966 B.n744 B.n141 163.367
R967 B.n748 B.n141 163.367
R968 B.n749 B.n748 163.367
R969 B.n750 B.n749 163.367
R970 B.n750 B.n139 163.367
R971 B.n754 B.n139 163.367
R972 B.n755 B.n754 163.367
R973 B.n756 B.n755 163.367
R974 B.n756 B.n137 163.367
R975 B.n760 B.n137 163.367
R976 B.n761 B.n760 163.367
R977 B.n762 B.n761 163.367
R978 B.n762 B.n135 163.367
R979 B.n766 B.n135 163.367
R980 B.n767 B.n766 163.367
R981 B.n768 B.n767 163.367
R982 B.n768 B.n133 163.367
R983 B.n772 B.n133 163.367
R984 B.n773 B.n772 163.367
R985 B.n774 B.n773 163.367
R986 B.n774 B.n131 163.367
R987 B.n778 B.n131 163.367
R988 B.n779 B.n778 163.367
R989 B.n780 B.n779 163.367
R990 B.n780 B.n129 163.367
R991 B.n784 B.n129 163.367
R992 B.n785 B.n784 163.367
R993 B.n786 B.n785 163.367
R994 B.n786 B.n127 163.367
R995 B.n790 B.n127 163.367
R996 B.n791 B.n790 163.367
R997 B.n792 B.n791 163.367
R998 B.n792 B.n125 163.367
R999 B.n796 B.n125 163.367
R1000 B.n797 B.n796 163.367
R1001 B.n798 B.n797 163.367
R1002 B.n798 B.n123 163.367
R1003 B.n802 B.n123 163.367
R1004 B.n803 B.n802 163.367
R1005 B.n804 B.n803 163.367
R1006 B.n804 B.n121 163.367
R1007 B.n808 B.n121 163.367
R1008 B.n809 B.n808 163.367
R1009 B.n810 B.n809 163.367
R1010 B.n810 B.n119 163.367
R1011 B.n814 B.n119 163.367
R1012 B.n815 B.n814 163.367
R1013 B.n816 B.n815 163.367
R1014 B.n816 B.n117 163.367
R1015 B.n820 B.n117 163.367
R1016 B.n821 B.n820 163.367
R1017 B.n822 B.n821 163.367
R1018 B.n822 B.n115 163.367
R1019 B.n826 B.n115 163.367
R1020 B.n827 B.n826 163.367
R1021 B.n828 B.n827 163.367
R1022 B.n828 B.n113 163.367
R1023 B.n832 B.n113 163.367
R1024 B.n833 B.n832 163.367
R1025 B.n834 B.n833 163.367
R1026 B.n834 B.n111 163.367
R1027 B.n838 B.n111 163.367
R1028 B.n839 B.n838 163.367
R1029 B.n840 B.n839 163.367
R1030 B.n840 B.n109 163.367
R1031 B.n844 B.n109 163.367
R1032 B.n1033 B.n1032 163.367
R1033 B.n1032 B.n43 163.367
R1034 B.n1028 B.n43 163.367
R1035 B.n1028 B.n1027 163.367
R1036 B.n1027 B.n1026 163.367
R1037 B.n1026 B.n45 163.367
R1038 B.n1022 B.n45 163.367
R1039 B.n1022 B.n1021 163.367
R1040 B.n1021 B.n1020 163.367
R1041 B.n1020 B.n47 163.367
R1042 B.n1016 B.n47 163.367
R1043 B.n1016 B.n1015 163.367
R1044 B.n1015 B.n1014 163.367
R1045 B.n1014 B.n49 163.367
R1046 B.n1010 B.n49 163.367
R1047 B.n1010 B.n1009 163.367
R1048 B.n1009 B.n1008 163.367
R1049 B.n1008 B.n51 163.367
R1050 B.n1004 B.n51 163.367
R1051 B.n1004 B.n1003 163.367
R1052 B.n1003 B.n1002 163.367
R1053 B.n1002 B.n53 163.367
R1054 B.n998 B.n53 163.367
R1055 B.n998 B.n997 163.367
R1056 B.n997 B.n996 163.367
R1057 B.n996 B.n55 163.367
R1058 B.n992 B.n55 163.367
R1059 B.n992 B.n991 163.367
R1060 B.n991 B.n990 163.367
R1061 B.n990 B.n57 163.367
R1062 B.n986 B.n57 163.367
R1063 B.n986 B.n985 163.367
R1064 B.n985 B.n984 163.367
R1065 B.n984 B.n59 163.367
R1066 B.n980 B.n59 163.367
R1067 B.n980 B.n979 163.367
R1068 B.n979 B.n978 163.367
R1069 B.n978 B.n61 163.367
R1070 B.n974 B.n61 163.367
R1071 B.n974 B.n973 163.367
R1072 B.n973 B.n972 163.367
R1073 B.n972 B.n63 163.367
R1074 B.n968 B.n63 163.367
R1075 B.n968 B.n967 163.367
R1076 B.n967 B.n966 163.367
R1077 B.n966 B.n65 163.367
R1078 B.n962 B.n65 163.367
R1079 B.n962 B.n961 163.367
R1080 B.n961 B.n960 163.367
R1081 B.n960 B.n67 163.367
R1082 B.n956 B.n67 163.367
R1083 B.n956 B.n955 163.367
R1084 B.n955 B.n954 163.367
R1085 B.n954 B.n69 163.367
R1086 B.n950 B.n69 163.367
R1087 B.n950 B.n949 163.367
R1088 B.n949 B.n948 163.367
R1089 B.n948 B.n71 163.367
R1090 B.n943 B.n71 163.367
R1091 B.n943 B.n942 163.367
R1092 B.n942 B.n941 163.367
R1093 B.n941 B.n75 163.367
R1094 B.n937 B.n75 163.367
R1095 B.n937 B.n936 163.367
R1096 B.n936 B.n935 163.367
R1097 B.n935 B.n77 163.367
R1098 B.n930 B.n77 163.367
R1099 B.n930 B.n929 163.367
R1100 B.n929 B.n928 163.367
R1101 B.n928 B.n81 163.367
R1102 B.n924 B.n81 163.367
R1103 B.n924 B.n923 163.367
R1104 B.n923 B.n922 163.367
R1105 B.n922 B.n83 163.367
R1106 B.n918 B.n83 163.367
R1107 B.n918 B.n917 163.367
R1108 B.n917 B.n916 163.367
R1109 B.n916 B.n85 163.367
R1110 B.n912 B.n85 163.367
R1111 B.n912 B.n911 163.367
R1112 B.n911 B.n910 163.367
R1113 B.n910 B.n87 163.367
R1114 B.n906 B.n87 163.367
R1115 B.n906 B.n905 163.367
R1116 B.n905 B.n904 163.367
R1117 B.n904 B.n89 163.367
R1118 B.n900 B.n89 163.367
R1119 B.n900 B.n899 163.367
R1120 B.n899 B.n898 163.367
R1121 B.n898 B.n91 163.367
R1122 B.n894 B.n91 163.367
R1123 B.n894 B.n893 163.367
R1124 B.n893 B.n892 163.367
R1125 B.n892 B.n93 163.367
R1126 B.n888 B.n93 163.367
R1127 B.n888 B.n887 163.367
R1128 B.n887 B.n886 163.367
R1129 B.n886 B.n95 163.367
R1130 B.n882 B.n95 163.367
R1131 B.n882 B.n881 163.367
R1132 B.n881 B.n880 163.367
R1133 B.n880 B.n97 163.367
R1134 B.n876 B.n97 163.367
R1135 B.n876 B.n875 163.367
R1136 B.n875 B.n874 163.367
R1137 B.n874 B.n99 163.367
R1138 B.n870 B.n99 163.367
R1139 B.n870 B.n869 163.367
R1140 B.n869 B.n868 163.367
R1141 B.n868 B.n101 163.367
R1142 B.n864 B.n101 163.367
R1143 B.n864 B.n863 163.367
R1144 B.n863 B.n862 163.367
R1145 B.n862 B.n103 163.367
R1146 B.n858 B.n103 163.367
R1147 B.n858 B.n857 163.367
R1148 B.n857 B.n856 163.367
R1149 B.n856 B.n105 163.367
R1150 B.n852 B.n105 163.367
R1151 B.n852 B.n851 163.367
R1152 B.n851 B.n850 163.367
R1153 B.n850 B.n107 163.367
R1154 B.n846 B.n107 163.367
R1155 B.n846 B.n845 163.367
R1156 B.n219 B.n218 78.9338
R1157 B.n227 B.n226 78.9338
R1158 B.n73 B.n72 78.9338
R1159 B.n79 B.n78 78.9338
R1160 B.n220 B.n219 59.5399
R1161 B.n501 B.n227 59.5399
R1162 B.n946 B.n73 59.5399
R1163 B.n932 B.n79 59.5399
R1164 B.n1035 B.n42 31.3761
R1165 B.n843 B.n108 31.3761
R1166 B.n603 B.n602 31.3761
R1167 B.n415 B.n256 31.3761
R1168 B B.n1155 18.0485
R1169 B.n1031 B.n42 10.6151
R1170 B.n1031 B.n1030 10.6151
R1171 B.n1030 B.n1029 10.6151
R1172 B.n1029 B.n44 10.6151
R1173 B.n1025 B.n44 10.6151
R1174 B.n1025 B.n1024 10.6151
R1175 B.n1024 B.n1023 10.6151
R1176 B.n1023 B.n46 10.6151
R1177 B.n1019 B.n46 10.6151
R1178 B.n1019 B.n1018 10.6151
R1179 B.n1018 B.n1017 10.6151
R1180 B.n1017 B.n48 10.6151
R1181 B.n1013 B.n48 10.6151
R1182 B.n1013 B.n1012 10.6151
R1183 B.n1012 B.n1011 10.6151
R1184 B.n1011 B.n50 10.6151
R1185 B.n1007 B.n50 10.6151
R1186 B.n1007 B.n1006 10.6151
R1187 B.n1006 B.n1005 10.6151
R1188 B.n1005 B.n52 10.6151
R1189 B.n1001 B.n52 10.6151
R1190 B.n1001 B.n1000 10.6151
R1191 B.n1000 B.n999 10.6151
R1192 B.n999 B.n54 10.6151
R1193 B.n995 B.n54 10.6151
R1194 B.n995 B.n994 10.6151
R1195 B.n994 B.n993 10.6151
R1196 B.n993 B.n56 10.6151
R1197 B.n989 B.n56 10.6151
R1198 B.n989 B.n988 10.6151
R1199 B.n988 B.n987 10.6151
R1200 B.n987 B.n58 10.6151
R1201 B.n983 B.n58 10.6151
R1202 B.n983 B.n982 10.6151
R1203 B.n982 B.n981 10.6151
R1204 B.n981 B.n60 10.6151
R1205 B.n977 B.n60 10.6151
R1206 B.n977 B.n976 10.6151
R1207 B.n976 B.n975 10.6151
R1208 B.n975 B.n62 10.6151
R1209 B.n971 B.n62 10.6151
R1210 B.n971 B.n970 10.6151
R1211 B.n970 B.n969 10.6151
R1212 B.n969 B.n64 10.6151
R1213 B.n965 B.n64 10.6151
R1214 B.n965 B.n964 10.6151
R1215 B.n964 B.n963 10.6151
R1216 B.n963 B.n66 10.6151
R1217 B.n959 B.n66 10.6151
R1218 B.n959 B.n958 10.6151
R1219 B.n958 B.n957 10.6151
R1220 B.n957 B.n68 10.6151
R1221 B.n953 B.n68 10.6151
R1222 B.n953 B.n952 10.6151
R1223 B.n952 B.n951 10.6151
R1224 B.n951 B.n70 10.6151
R1225 B.n947 B.n70 10.6151
R1226 B.n945 B.n944 10.6151
R1227 B.n944 B.n74 10.6151
R1228 B.n940 B.n74 10.6151
R1229 B.n940 B.n939 10.6151
R1230 B.n939 B.n938 10.6151
R1231 B.n938 B.n76 10.6151
R1232 B.n934 B.n76 10.6151
R1233 B.n934 B.n933 10.6151
R1234 B.n931 B.n80 10.6151
R1235 B.n927 B.n80 10.6151
R1236 B.n927 B.n926 10.6151
R1237 B.n926 B.n925 10.6151
R1238 B.n925 B.n82 10.6151
R1239 B.n921 B.n82 10.6151
R1240 B.n921 B.n920 10.6151
R1241 B.n920 B.n919 10.6151
R1242 B.n919 B.n84 10.6151
R1243 B.n915 B.n84 10.6151
R1244 B.n915 B.n914 10.6151
R1245 B.n914 B.n913 10.6151
R1246 B.n913 B.n86 10.6151
R1247 B.n909 B.n86 10.6151
R1248 B.n909 B.n908 10.6151
R1249 B.n908 B.n907 10.6151
R1250 B.n907 B.n88 10.6151
R1251 B.n903 B.n88 10.6151
R1252 B.n903 B.n902 10.6151
R1253 B.n902 B.n901 10.6151
R1254 B.n901 B.n90 10.6151
R1255 B.n897 B.n90 10.6151
R1256 B.n897 B.n896 10.6151
R1257 B.n896 B.n895 10.6151
R1258 B.n895 B.n92 10.6151
R1259 B.n891 B.n92 10.6151
R1260 B.n891 B.n890 10.6151
R1261 B.n890 B.n889 10.6151
R1262 B.n889 B.n94 10.6151
R1263 B.n885 B.n94 10.6151
R1264 B.n885 B.n884 10.6151
R1265 B.n884 B.n883 10.6151
R1266 B.n883 B.n96 10.6151
R1267 B.n879 B.n96 10.6151
R1268 B.n879 B.n878 10.6151
R1269 B.n878 B.n877 10.6151
R1270 B.n877 B.n98 10.6151
R1271 B.n873 B.n98 10.6151
R1272 B.n873 B.n872 10.6151
R1273 B.n872 B.n871 10.6151
R1274 B.n871 B.n100 10.6151
R1275 B.n867 B.n100 10.6151
R1276 B.n867 B.n866 10.6151
R1277 B.n866 B.n865 10.6151
R1278 B.n865 B.n102 10.6151
R1279 B.n861 B.n102 10.6151
R1280 B.n861 B.n860 10.6151
R1281 B.n860 B.n859 10.6151
R1282 B.n859 B.n104 10.6151
R1283 B.n855 B.n104 10.6151
R1284 B.n855 B.n854 10.6151
R1285 B.n854 B.n853 10.6151
R1286 B.n853 B.n106 10.6151
R1287 B.n849 B.n106 10.6151
R1288 B.n849 B.n848 10.6151
R1289 B.n848 B.n847 10.6151
R1290 B.n847 B.n108 10.6151
R1291 B.n603 B.n188 10.6151
R1292 B.n607 B.n188 10.6151
R1293 B.n608 B.n607 10.6151
R1294 B.n609 B.n608 10.6151
R1295 B.n609 B.n186 10.6151
R1296 B.n613 B.n186 10.6151
R1297 B.n614 B.n613 10.6151
R1298 B.n615 B.n614 10.6151
R1299 B.n615 B.n184 10.6151
R1300 B.n619 B.n184 10.6151
R1301 B.n620 B.n619 10.6151
R1302 B.n621 B.n620 10.6151
R1303 B.n621 B.n182 10.6151
R1304 B.n625 B.n182 10.6151
R1305 B.n626 B.n625 10.6151
R1306 B.n627 B.n626 10.6151
R1307 B.n627 B.n180 10.6151
R1308 B.n631 B.n180 10.6151
R1309 B.n632 B.n631 10.6151
R1310 B.n633 B.n632 10.6151
R1311 B.n633 B.n178 10.6151
R1312 B.n637 B.n178 10.6151
R1313 B.n638 B.n637 10.6151
R1314 B.n639 B.n638 10.6151
R1315 B.n639 B.n176 10.6151
R1316 B.n643 B.n176 10.6151
R1317 B.n644 B.n643 10.6151
R1318 B.n645 B.n644 10.6151
R1319 B.n645 B.n174 10.6151
R1320 B.n649 B.n174 10.6151
R1321 B.n650 B.n649 10.6151
R1322 B.n651 B.n650 10.6151
R1323 B.n651 B.n172 10.6151
R1324 B.n655 B.n172 10.6151
R1325 B.n656 B.n655 10.6151
R1326 B.n657 B.n656 10.6151
R1327 B.n657 B.n170 10.6151
R1328 B.n661 B.n170 10.6151
R1329 B.n662 B.n661 10.6151
R1330 B.n663 B.n662 10.6151
R1331 B.n663 B.n168 10.6151
R1332 B.n667 B.n168 10.6151
R1333 B.n668 B.n667 10.6151
R1334 B.n669 B.n668 10.6151
R1335 B.n669 B.n166 10.6151
R1336 B.n673 B.n166 10.6151
R1337 B.n674 B.n673 10.6151
R1338 B.n675 B.n674 10.6151
R1339 B.n675 B.n164 10.6151
R1340 B.n679 B.n164 10.6151
R1341 B.n680 B.n679 10.6151
R1342 B.n681 B.n680 10.6151
R1343 B.n681 B.n162 10.6151
R1344 B.n685 B.n162 10.6151
R1345 B.n686 B.n685 10.6151
R1346 B.n687 B.n686 10.6151
R1347 B.n687 B.n160 10.6151
R1348 B.n691 B.n160 10.6151
R1349 B.n692 B.n691 10.6151
R1350 B.n693 B.n692 10.6151
R1351 B.n693 B.n158 10.6151
R1352 B.n697 B.n158 10.6151
R1353 B.n698 B.n697 10.6151
R1354 B.n699 B.n698 10.6151
R1355 B.n699 B.n156 10.6151
R1356 B.n703 B.n156 10.6151
R1357 B.n704 B.n703 10.6151
R1358 B.n705 B.n704 10.6151
R1359 B.n705 B.n154 10.6151
R1360 B.n709 B.n154 10.6151
R1361 B.n710 B.n709 10.6151
R1362 B.n711 B.n710 10.6151
R1363 B.n711 B.n152 10.6151
R1364 B.n715 B.n152 10.6151
R1365 B.n716 B.n715 10.6151
R1366 B.n717 B.n716 10.6151
R1367 B.n717 B.n150 10.6151
R1368 B.n721 B.n150 10.6151
R1369 B.n722 B.n721 10.6151
R1370 B.n723 B.n722 10.6151
R1371 B.n723 B.n148 10.6151
R1372 B.n727 B.n148 10.6151
R1373 B.n728 B.n727 10.6151
R1374 B.n729 B.n728 10.6151
R1375 B.n729 B.n146 10.6151
R1376 B.n733 B.n146 10.6151
R1377 B.n734 B.n733 10.6151
R1378 B.n735 B.n734 10.6151
R1379 B.n735 B.n144 10.6151
R1380 B.n739 B.n144 10.6151
R1381 B.n740 B.n739 10.6151
R1382 B.n741 B.n740 10.6151
R1383 B.n741 B.n142 10.6151
R1384 B.n745 B.n142 10.6151
R1385 B.n746 B.n745 10.6151
R1386 B.n747 B.n746 10.6151
R1387 B.n747 B.n140 10.6151
R1388 B.n751 B.n140 10.6151
R1389 B.n752 B.n751 10.6151
R1390 B.n753 B.n752 10.6151
R1391 B.n753 B.n138 10.6151
R1392 B.n757 B.n138 10.6151
R1393 B.n758 B.n757 10.6151
R1394 B.n759 B.n758 10.6151
R1395 B.n759 B.n136 10.6151
R1396 B.n763 B.n136 10.6151
R1397 B.n764 B.n763 10.6151
R1398 B.n765 B.n764 10.6151
R1399 B.n765 B.n134 10.6151
R1400 B.n769 B.n134 10.6151
R1401 B.n770 B.n769 10.6151
R1402 B.n771 B.n770 10.6151
R1403 B.n771 B.n132 10.6151
R1404 B.n775 B.n132 10.6151
R1405 B.n776 B.n775 10.6151
R1406 B.n777 B.n776 10.6151
R1407 B.n777 B.n130 10.6151
R1408 B.n781 B.n130 10.6151
R1409 B.n782 B.n781 10.6151
R1410 B.n783 B.n782 10.6151
R1411 B.n783 B.n128 10.6151
R1412 B.n787 B.n128 10.6151
R1413 B.n788 B.n787 10.6151
R1414 B.n789 B.n788 10.6151
R1415 B.n789 B.n126 10.6151
R1416 B.n793 B.n126 10.6151
R1417 B.n794 B.n793 10.6151
R1418 B.n795 B.n794 10.6151
R1419 B.n795 B.n124 10.6151
R1420 B.n799 B.n124 10.6151
R1421 B.n800 B.n799 10.6151
R1422 B.n801 B.n800 10.6151
R1423 B.n801 B.n122 10.6151
R1424 B.n805 B.n122 10.6151
R1425 B.n806 B.n805 10.6151
R1426 B.n807 B.n806 10.6151
R1427 B.n807 B.n120 10.6151
R1428 B.n811 B.n120 10.6151
R1429 B.n812 B.n811 10.6151
R1430 B.n813 B.n812 10.6151
R1431 B.n813 B.n118 10.6151
R1432 B.n817 B.n118 10.6151
R1433 B.n818 B.n817 10.6151
R1434 B.n819 B.n818 10.6151
R1435 B.n819 B.n116 10.6151
R1436 B.n823 B.n116 10.6151
R1437 B.n824 B.n823 10.6151
R1438 B.n825 B.n824 10.6151
R1439 B.n825 B.n114 10.6151
R1440 B.n829 B.n114 10.6151
R1441 B.n830 B.n829 10.6151
R1442 B.n831 B.n830 10.6151
R1443 B.n831 B.n112 10.6151
R1444 B.n835 B.n112 10.6151
R1445 B.n836 B.n835 10.6151
R1446 B.n837 B.n836 10.6151
R1447 B.n837 B.n110 10.6151
R1448 B.n841 B.n110 10.6151
R1449 B.n842 B.n841 10.6151
R1450 B.n843 B.n842 10.6151
R1451 B.n416 B.n415 10.6151
R1452 B.n417 B.n416 10.6151
R1453 B.n417 B.n254 10.6151
R1454 B.n421 B.n254 10.6151
R1455 B.n422 B.n421 10.6151
R1456 B.n423 B.n422 10.6151
R1457 B.n423 B.n252 10.6151
R1458 B.n427 B.n252 10.6151
R1459 B.n428 B.n427 10.6151
R1460 B.n429 B.n428 10.6151
R1461 B.n429 B.n250 10.6151
R1462 B.n433 B.n250 10.6151
R1463 B.n434 B.n433 10.6151
R1464 B.n435 B.n434 10.6151
R1465 B.n435 B.n248 10.6151
R1466 B.n439 B.n248 10.6151
R1467 B.n440 B.n439 10.6151
R1468 B.n441 B.n440 10.6151
R1469 B.n441 B.n246 10.6151
R1470 B.n445 B.n246 10.6151
R1471 B.n446 B.n445 10.6151
R1472 B.n447 B.n446 10.6151
R1473 B.n447 B.n244 10.6151
R1474 B.n451 B.n244 10.6151
R1475 B.n452 B.n451 10.6151
R1476 B.n453 B.n452 10.6151
R1477 B.n453 B.n242 10.6151
R1478 B.n457 B.n242 10.6151
R1479 B.n458 B.n457 10.6151
R1480 B.n459 B.n458 10.6151
R1481 B.n459 B.n240 10.6151
R1482 B.n463 B.n240 10.6151
R1483 B.n464 B.n463 10.6151
R1484 B.n465 B.n464 10.6151
R1485 B.n465 B.n238 10.6151
R1486 B.n469 B.n238 10.6151
R1487 B.n470 B.n469 10.6151
R1488 B.n471 B.n470 10.6151
R1489 B.n471 B.n236 10.6151
R1490 B.n475 B.n236 10.6151
R1491 B.n476 B.n475 10.6151
R1492 B.n477 B.n476 10.6151
R1493 B.n477 B.n234 10.6151
R1494 B.n481 B.n234 10.6151
R1495 B.n482 B.n481 10.6151
R1496 B.n483 B.n482 10.6151
R1497 B.n483 B.n232 10.6151
R1498 B.n487 B.n232 10.6151
R1499 B.n488 B.n487 10.6151
R1500 B.n489 B.n488 10.6151
R1501 B.n489 B.n230 10.6151
R1502 B.n493 B.n230 10.6151
R1503 B.n494 B.n493 10.6151
R1504 B.n495 B.n494 10.6151
R1505 B.n495 B.n228 10.6151
R1506 B.n499 B.n228 10.6151
R1507 B.n500 B.n499 10.6151
R1508 B.n502 B.n224 10.6151
R1509 B.n506 B.n224 10.6151
R1510 B.n507 B.n506 10.6151
R1511 B.n508 B.n507 10.6151
R1512 B.n508 B.n222 10.6151
R1513 B.n512 B.n222 10.6151
R1514 B.n513 B.n512 10.6151
R1515 B.n514 B.n513 10.6151
R1516 B.n518 B.n517 10.6151
R1517 B.n519 B.n518 10.6151
R1518 B.n519 B.n216 10.6151
R1519 B.n523 B.n216 10.6151
R1520 B.n524 B.n523 10.6151
R1521 B.n525 B.n524 10.6151
R1522 B.n525 B.n214 10.6151
R1523 B.n529 B.n214 10.6151
R1524 B.n530 B.n529 10.6151
R1525 B.n531 B.n530 10.6151
R1526 B.n531 B.n212 10.6151
R1527 B.n535 B.n212 10.6151
R1528 B.n536 B.n535 10.6151
R1529 B.n537 B.n536 10.6151
R1530 B.n537 B.n210 10.6151
R1531 B.n541 B.n210 10.6151
R1532 B.n542 B.n541 10.6151
R1533 B.n543 B.n542 10.6151
R1534 B.n543 B.n208 10.6151
R1535 B.n547 B.n208 10.6151
R1536 B.n548 B.n547 10.6151
R1537 B.n549 B.n548 10.6151
R1538 B.n549 B.n206 10.6151
R1539 B.n553 B.n206 10.6151
R1540 B.n554 B.n553 10.6151
R1541 B.n555 B.n554 10.6151
R1542 B.n555 B.n204 10.6151
R1543 B.n559 B.n204 10.6151
R1544 B.n560 B.n559 10.6151
R1545 B.n561 B.n560 10.6151
R1546 B.n561 B.n202 10.6151
R1547 B.n565 B.n202 10.6151
R1548 B.n566 B.n565 10.6151
R1549 B.n567 B.n566 10.6151
R1550 B.n567 B.n200 10.6151
R1551 B.n571 B.n200 10.6151
R1552 B.n572 B.n571 10.6151
R1553 B.n573 B.n572 10.6151
R1554 B.n573 B.n198 10.6151
R1555 B.n577 B.n198 10.6151
R1556 B.n578 B.n577 10.6151
R1557 B.n579 B.n578 10.6151
R1558 B.n579 B.n196 10.6151
R1559 B.n583 B.n196 10.6151
R1560 B.n584 B.n583 10.6151
R1561 B.n585 B.n584 10.6151
R1562 B.n585 B.n194 10.6151
R1563 B.n589 B.n194 10.6151
R1564 B.n590 B.n589 10.6151
R1565 B.n591 B.n590 10.6151
R1566 B.n591 B.n192 10.6151
R1567 B.n595 B.n192 10.6151
R1568 B.n596 B.n595 10.6151
R1569 B.n597 B.n596 10.6151
R1570 B.n597 B.n190 10.6151
R1571 B.n601 B.n190 10.6151
R1572 B.n602 B.n601 10.6151
R1573 B.n411 B.n256 10.6151
R1574 B.n411 B.n410 10.6151
R1575 B.n410 B.n409 10.6151
R1576 B.n409 B.n258 10.6151
R1577 B.n405 B.n258 10.6151
R1578 B.n405 B.n404 10.6151
R1579 B.n404 B.n403 10.6151
R1580 B.n403 B.n260 10.6151
R1581 B.n399 B.n260 10.6151
R1582 B.n399 B.n398 10.6151
R1583 B.n398 B.n397 10.6151
R1584 B.n397 B.n262 10.6151
R1585 B.n393 B.n262 10.6151
R1586 B.n393 B.n392 10.6151
R1587 B.n392 B.n391 10.6151
R1588 B.n391 B.n264 10.6151
R1589 B.n387 B.n264 10.6151
R1590 B.n387 B.n386 10.6151
R1591 B.n386 B.n385 10.6151
R1592 B.n385 B.n266 10.6151
R1593 B.n381 B.n266 10.6151
R1594 B.n381 B.n380 10.6151
R1595 B.n380 B.n379 10.6151
R1596 B.n379 B.n268 10.6151
R1597 B.n375 B.n268 10.6151
R1598 B.n375 B.n374 10.6151
R1599 B.n374 B.n373 10.6151
R1600 B.n373 B.n270 10.6151
R1601 B.n369 B.n270 10.6151
R1602 B.n369 B.n368 10.6151
R1603 B.n368 B.n367 10.6151
R1604 B.n367 B.n272 10.6151
R1605 B.n363 B.n272 10.6151
R1606 B.n363 B.n362 10.6151
R1607 B.n362 B.n361 10.6151
R1608 B.n361 B.n274 10.6151
R1609 B.n357 B.n274 10.6151
R1610 B.n357 B.n356 10.6151
R1611 B.n356 B.n355 10.6151
R1612 B.n355 B.n276 10.6151
R1613 B.n351 B.n276 10.6151
R1614 B.n351 B.n350 10.6151
R1615 B.n350 B.n349 10.6151
R1616 B.n349 B.n278 10.6151
R1617 B.n345 B.n278 10.6151
R1618 B.n345 B.n344 10.6151
R1619 B.n344 B.n343 10.6151
R1620 B.n343 B.n280 10.6151
R1621 B.n339 B.n280 10.6151
R1622 B.n339 B.n338 10.6151
R1623 B.n338 B.n337 10.6151
R1624 B.n337 B.n282 10.6151
R1625 B.n333 B.n282 10.6151
R1626 B.n333 B.n332 10.6151
R1627 B.n332 B.n331 10.6151
R1628 B.n331 B.n284 10.6151
R1629 B.n327 B.n284 10.6151
R1630 B.n327 B.n326 10.6151
R1631 B.n326 B.n325 10.6151
R1632 B.n325 B.n286 10.6151
R1633 B.n321 B.n286 10.6151
R1634 B.n321 B.n320 10.6151
R1635 B.n320 B.n319 10.6151
R1636 B.n319 B.n288 10.6151
R1637 B.n315 B.n288 10.6151
R1638 B.n315 B.n314 10.6151
R1639 B.n314 B.n313 10.6151
R1640 B.n313 B.n290 10.6151
R1641 B.n309 B.n290 10.6151
R1642 B.n309 B.n308 10.6151
R1643 B.n308 B.n307 10.6151
R1644 B.n307 B.n292 10.6151
R1645 B.n303 B.n292 10.6151
R1646 B.n303 B.n302 10.6151
R1647 B.n302 B.n301 10.6151
R1648 B.n301 B.n294 10.6151
R1649 B.n297 B.n294 10.6151
R1650 B.n297 B.n296 10.6151
R1651 B.n296 B.n0 10.6151
R1652 B.n1151 B.n1 10.6151
R1653 B.n1151 B.n1150 10.6151
R1654 B.n1150 B.n1149 10.6151
R1655 B.n1149 B.n4 10.6151
R1656 B.n1145 B.n4 10.6151
R1657 B.n1145 B.n1144 10.6151
R1658 B.n1144 B.n1143 10.6151
R1659 B.n1143 B.n6 10.6151
R1660 B.n1139 B.n6 10.6151
R1661 B.n1139 B.n1138 10.6151
R1662 B.n1138 B.n1137 10.6151
R1663 B.n1137 B.n8 10.6151
R1664 B.n1133 B.n8 10.6151
R1665 B.n1133 B.n1132 10.6151
R1666 B.n1132 B.n1131 10.6151
R1667 B.n1131 B.n10 10.6151
R1668 B.n1127 B.n10 10.6151
R1669 B.n1127 B.n1126 10.6151
R1670 B.n1126 B.n1125 10.6151
R1671 B.n1125 B.n12 10.6151
R1672 B.n1121 B.n12 10.6151
R1673 B.n1121 B.n1120 10.6151
R1674 B.n1120 B.n1119 10.6151
R1675 B.n1119 B.n14 10.6151
R1676 B.n1115 B.n14 10.6151
R1677 B.n1115 B.n1114 10.6151
R1678 B.n1114 B.n1113 10.6151
R1679 B.n1113 B.n16 10.6151
R1680 B.n1109 B.n16 10.6151
R1681 B.n1109 B.n1108 10.6151
R1682 B.n1108 B.n1107 10.6151
R1683 B.n1107 B.n18 10.6151
R1684 B.n1103 B.n18 10.6151
R1685 B.n1103 B.n1102 10.6151
R1686 B.n1102 B.n1101 10.6151
R1687 B.n1101 B.n20 10.6151
R1688 B.n1097 B.n20 10.6151
R1689 B.n1097 B.n1096 10.6151
R1690 B.n1096 B.n1095 10.6151
R1691 B.n1095 B.n22 10.6151
R1692 B.n1091 B.n22 10.6151
R1693 B.n1091 B.n1090 10.6151
R1694 B.n1090 B.n1089 10.6151
R1695 B.n1089 B.n24 10.6151
R1696 B.n1085 B.n24 10.6151
R1697 B.n1085 B.n1084 10.6151
R1698 B.n1084 B.n1083 10.6151
R1699 B.n1083 B.n26 10.6151
R1700 B.n1079 B.n26 10.6151
R1701 B.n1079 B.n1078 10.6151
R1702 B.n1078 B.n1077 10.6151
R1703 B.n1077 B.n28 10.6151
R1704 B.n1073 B.n28 10.6151
R1705 B.n1073 B.n1072 10.6151
R1706 B.n1072 B.n1071 10.6151
R1707 B.n1071 B.n30 10.6151
R1708 B.n1067 B.n30 10.6151
R1709 B.n1067 B.n1066 10.6151
R1710 B.n1066 B.n1065 10.6151
R1711 B.n1065 B.n32 10.6151
R1712 B.n1061 B.n32 10.6151
R1713 B.n1061 B.n1060 10.6151
R1714 B.n1060 B.n1059 10.6151
R1715 B.n1059 B.n34 10.6151
R1716 B.n1055 B.n34 10.6151
R1717 B.n1055 B.n1054 10.6151
R1718 B.n1054 B.n1053 10.6151
R1719 B.n1053 B.n36 10.6151
R1720 B.n1049 B.n36 10.6151
R1721 B.n1049 B.n1048 10.6151
R1722 B.n1048 B.n1047 10.6151
R1723 B.n1047 B.n38 10.6151
R1724 B.n1043 B.n38 10.6151
R1725 B.n1043 B.n1042 10.6151
R1726 B.n1042 B.n1041 10.6151
R1727 B.n1041 B.n40 10.6151
R1728 B.n1037 B.n40 10.6151
R1729 B.n1037 B.n1036 10.6151
R1730 B.n1036 B.n1035 10.6151
R1731 B.n946 B.n945 6.5566
R1732 B.n933 B.n932 6.5566
R1733 B.n502 B.n501 6.5566
R1734 B.n514 B.n220 6.5566
R1735 B.n947 B.n946 4.05904
R1736 B.n932 B.n931 4.05904
R1737 B.n501 B.n500 4.05904
R1738 B.n517 B.n220 4.05904
R1739 B.n1155 B.n0 2.81026
R1740 B.n1155 B.n1 2.81026
R1741 VP.n33 VP.n32 161.3
R1742 VP.n34 VP.n29 161.3
R1743 VP.n36 VP.n35 161.3
R1744 VP.n37 VP.n28 161.3
R1745 VP.n39 VP.n38 161.3
R1746 VP.n40 VP.n27 161.3
R1747 VP.n42 VP.n41 161.3
R1748 VP.n43 VP.n26 161.3
R1749 VP.n45 VP.n44 161.3
R1750 VP.n46 VP.n25 161.3
R1751 VP.n48 VP.n47 161.3
R1752 VP.n49 VP.n24 161.3
R1753 VP.n51 VP.n50 161.3
R1754 VP.n52 VP.n23 161.3
R1755 VP.n54 VP.n53 161.3
R1756 VP.n55 VP.n22 161.3
R1757 VP.n58 VP.n57 161.3
R1758 VP.n59 VP.n21 161.3
R1759 VP.n61 VP.n60 161.3
R1760 VP.n62 VP.n20 161.3
R1761 VP.n64 VP.n63 161.3
R1762 VP.n65 VP.n19 161.3
R1763 VP.n67 VP.n66 161.3
R1764 VP.n68 VP.n18 161.3
R1765 VP.n70 VP.n69 161.3
R1766 VP.n125 VP.n124 161.3
R1767 VP.n123 VP.n1 161.3
R1768 VP.n122 VP.n121 161.3
R1769 VP.n120 VP.n2 161.3
R1770 VP.n119 VP.n118 161.3
R1771 VP.n117 VP.n3 161.3
R1772 VP.n116 VP.n115 161.3
R1773 VP.n114 VP.n4 161.3
R1774 VP.n113 VP.n112 161.3
R1775 VP.n110 VP.n5 161.3
R1776 VP.n109 VP.n108 161.3
R1777 VP.n107 VP.n6 161.3
R1778 VP.n106 VP.n105 161.3
R1779 VP.n104 VP.n7 161.3
R1780 VP.n103 VP.n102 161.3
R1781 VP.n101 VP.n8 161.3
R1782 VP.n100 VP.n99 161.3
R1783 VP.n98 VP.n9 161.3
R1784 VP.n97 VP.n96 161.3
R1785 VP.n95 VP.n10 161.3
R1786 VP.n94 VP.n93 161.3
R1787 VP.n92 VP.n11 161.3
R1788 VP.n91 VP.n90 161.3
R1789 VP.n89 VP.n12 161.3
R1790 VP.n88 VP.n87 161.3
R1791 VP.n85 VP.n13 161.3
R1792 VP.n84 VP.n83 161.3
R1793 VP.n82 VP.n14 161.3
R1794 VP.n81 VP.n80 161.3
R1795 VP.n79 VP.n15 161.3
R1796 VP.n78 VP.n77 161.3
R1797 VP.n76 VP.n16 161.3
R1798 VP.n75 VP.n74 161.3
R1799 VP.n30 VP.t7 145.398
R1800 VP.n99 VP.t5 112.51
R1801 VP.n73 VP.t9 112.51
R1802 VP.n86 VP.t2 112.51
R1803 VP.n111 VP.t0 112.51
R1804 VP.n0 VP.t3 112.51
R1805 VP.n44 VP.t6 112.51
R1806 VP.n17 VP.t1 112.51
R1807 VP.n56 VP.t4 112.51
R1808 VP.n31 VP.t8 112.51
R1809 VP.n73 VP.n72 83.3598
R1810 VP.n126 VP.n0 83.3598
R1811 VP.n71 VP.n17 83.3598
R1812 VP.n31 VP.n30 71.5921
R1813 VP.n72 VP.n71 63.5488
R1814 VP.n80 VP.n79 50.7491
R1815 VP.n118 VP.n2 50.7491
R1816 VP.n63 VP.n19 50.7491
R1817 VP.n93 VP.n92 43.9677
R1818 VP.n105 VP.n6 43.9677
R1819 VP.n50 VP.n23 43.9677
R1820 VP.n38 VP.n37 43.9677
R1821 VP.n93 VP.n10 37.1863
R1822 VP.n105 VP.n104 37.1863
R1823 VP.n50 VP.n49 37.1863
R1824 VP.n38 VP.n27 37.1863
R1825 VP.n80 VP.n14 30.405
R1826 VP.n118 VP.n117 30.405
R1827 VP.n63 VP.n62 30.405
R1828 VP.n74 VP.n16 24.5923
R1829 VP.n78 VP.n16 24.5923
R1830 VP.n79 VP.n78 24.5923
R1831 VP.n84 VP.n14 24.5923
R1832 VP.n85 VP.n84 24.5923
R1833 VP.n87 VP.n12 24.5923
R1834 VP.n91 VP.n12 24.5923
R1835 VP.n92 VP.n91 24.5923
R1836 VP.n97 VP.n10 24.5923
R1837 VP.n98 VP.n97 24.5923
R1838 VP.n99 VP.n98 24.5923
R1839 VP.n99 VP.n8 24.5923
R1840 VP.n103 VP.n8 24.5923
R1841 VP.n104 VP.n103 24.5923
R1842 VP.n109 VP.n6 24.5923
R1843 VP.n110 VP.n109 24.5923
R1844 VP.n112 VP.n110 24.5923
R1845 VP.n116 VP.n4 24.5923
R1846 VP.n117 VP.n116 24.5923
R1847 VP.n122 VP.n2 24.5923
R1848 VP.n123 VP.n122 24.5923
R1849 VP.n124 VP.n123 24.5923
R1850 VP.n67 VP.n19 24.5923
R1851 VP.n68 VP.n67 24.5923
R1852 VP.n69 VP.n68 24.5923
R1853 VP.n54 VP.n23 24.5923
R1854 VP.n55 VP.n54 24.5923
R1855 VP.n57 VP.n55 24.5923
R1856 VP.n61 VP.n21 24.5923
R1857 VP.n62 VP.n61 24.5923
R1858 VP.n42 VP.n27 24.5923
R1859 VP.n43 VP.n42 24.5923
R1860 VP.n44 VP.n43 24.5923
R1861 VP.n44 VP.n25 24.5923
R1862 VP.n48 VP.n25 24.5923
R1863 VP.n49 VP.n48 24.5923
R1864 VP.n32 VP.n29 24.5923
R1865 VP.n36 VP.n29 24.5923
R1866 VP.n37 VP.n36 24.5923
R1867 VP.n86 VP.n85 21.1495
R1868 VP.n111 VP.n4 21.1495
R1869 VP.n56 VP.n21 21.1495
R1870 VP.n74 VP.n73 6.88621
R1871 VP.n124 VP.n0 6.88621
R1872 VP.n69 VP.n17 6.88621
R1873 VP.n87 VP.n86 3.44336
R1874 VP.n112 VP.n111 3.44336
R1875 VP.n57 VP.n56 3.44336
R1876 VP.n32 VP.n31 3.44336
R1877 VP.n33 VP.n30 3.23942
R1878 VP.n71 VP.n70 0.354861
R1879 VP.n75 VP.n72 0.354861
R1880 VP.n126 VP.n125 0.354861
R1881 VP VP.n126 0.267071
R1882 VP.n34 VP.n33 0.189894
R1883 VP.n35 VP.n34 0.189894
R1884 VP.n35 VP.n28 0.189894
R1885 VP.n39 VP.n28 0.189894
R1886 VP.n40 VP.n39 0.189894
R1887 VP.n41 VP.n40 0.189894
R1888 VP.n41 VP.n26 0.189894
R1889 VP.n45 VP.n26 0.189894
R1890 VP.n46 VP.n45 0.189894
R1891 VP.n47 VP.n46 0.189894
R1892 VP.n47 VP.n24 0.189894
R1893 VP.n51 VP.n24 0.189894
R1894 VP.n52 VP.n51 0.189894
R1895 VP.n53 VP.n52 0.189894
R1896 VP.n53 VP.n22 0.189894
R1897 VP.n58 VP.n22 0.189894
R1898 VP.n59 VP.n58 0.189894
R1899 VP.n60 VP.n59 0.189894
R1900 VP.n60 VP.n20 0.189894
R1901 VP.n64 VP.n20 0.189894
R1902 VP.n65 VP.n64 0.189894
R1903 VP.n66 VP.n65 0.189894
R1904 VP.n66 VP.n18 0.189894
R1905 VP.n70 VP.n18 0.189894
R1906 VP.n76 VP.n75 0.189894
R1907 VP.n77 VP.n76 0.189894
R1908 VP.n77 VP.n15 0.189894
R1909 VP.n81 VP.n15 0.189894
R1910 VP.n82 VP.n81 0.189894
R1911 VP.n83 VP.n82 0.189894
R1912 VP.n83 VP.n13 0.189894
R1913 VP.n88 VP.n13 0.189894
R1914 VP.n89 VP.n88 0.189894
R1915 VP.n90 VP.n89 0.189894
R1916 VP.n90 VP.n11 0.189894
R1917 VP.n94 VP.n11 0.189894
R1918 VP.n95 VP.n94 0.189894
R1919 VP.n96 VP.n95 0.189894
R1920 VP.n96 VP.n9 0.189894
R1921 VP.n100 VP.n9 0.189894
R1922 VP.n101 VP.n100 0.189894
R1923 VP.n102 VP.n101 0.189894
R1924 VP.n102 VP.n7 0.189894
R1925 VP.n106 VP.n7 0.189894
R1926 VP.n107 VP.n106 0.189894
R1927 VP.n108 VP.n107 0.189894
R1928 VP.n108 VP.n5 0.189894
R1929 VP.n113 VP.n5 0.189894
R1930 VP.n114 VP.n113 0.189894
R1931 VP.n115 VP.n114 0.189894
R1932 VP.n115 VP.n3 0.189894
R1933 VP.n119 VP.n3 0.189894
R1934 VP.n120 VP.n119 0.189894
R1935 VP.n121 VP.n120 0.189894
R1936 VP.n121 VP.n1 0.189894
R1937 VP.n125 VP.n1 0.189894
R1938 VDD1.n92 VDD1.n0 756.745
R1939 VDD1.n191 VDD1.n99 756.745
R1940 VDD1.n93 VDD1.n92 585
R1941 VDD1.n91 VDD1.n90 585
R1942 VDD1.n4 VDD1.n3 585
R1943 VDD1.n85 VDD1.n84 585
R1944 VDD1.n83 VDD1.n82 585
R1945 VDD1.n8 VDD1.n7 585
R1946 VDD1.n12 VDD1.n10 585
R1947 VDD1.n77 VDD1.n76 585
R1948 VDD1.n75 VDD1.n74 585
R1949 VDD1.n14 VDD1.n13 585
R1950 VDD1.n69 VDD1.n68 585
R1951 VDD1.n67 VDD1.n66 585
R1952 VDD1.n18 VDD1.n17 585
R1953 VDD1.n61 VDD1.n60 585
R1954 VDD1.n59 VDD1.n58 585
R1955 VDD1.n22 VDD1.n21 585
R1956 VDD1.n53 VDD1.n52 585
R1957 VDD1.n51 VDD1.n50 585
R1958 VDD1.n26 VDD1.n25 585
R1959 VDD1.n45 VDD1.n44 585
R1960 VDD1.n43 VDD1.n42 585
R1961 VDD1.n30 VDD1.n29 585
R1962 VDD1.n37 VDD1.n36 585
R1963 VDD1.n35 VDD1.n34 585
R1964 VDD1.n132 VDD1.n131 585
R1965 VDD1.n134 VDD1.n133 585
R1966 VDD1.n127 VDD1.n126 585
R1967 VDD1.n140 VDD1.n139 585
R1968 VDD1.n142 VDD1.n141 585
R1969 VDD1.n123 VDD1.n122 585
R1970 VDD1.n148 VDD1.n147 585
R1971 VDD1.n150 VDD1.n149 585
R1972 VDD1.n119 VDD1.n118 585
R1973 VDD1.n156 VDD1.n155 585
R1974 VDD1.n158 VDD1.n157 585
R1975 VDD1.n115 VDD1.n114 585
R1976 VDD1.n164 VDD1.n163 585
R1977 VDD1.n166 VDD1.n165 585
R1978 VDD1.n111 VDD1.n110 585
R1979 VDD1.n173 VDD1.n172 585
R1980 VDD1.n174 VDD1.n109 585
R1981 VDD1.n176 VDD1.n175 585
R1982 VDD1.n107 VDD1.n106 585
R1983 VDD1.n182 VDD1.n181 585
R1984 VDD1.n184 VDD1.n183 585
R1985 VDD1.n103 VDD1.n102 585
R1986 VDD1.n190 VDD1.n189 585
R1987 VDD1.n192 VDD1.n191 585
R1988 VDD1.n33 VDD1.t7 327.466
R1989 VDD1.n130 VDD1.t6 327.466
R1990 VDD1.n92 VDD1.n91 171.744
R1991 VDD1.n91 VDD1.n3 171.744
R1992 VDD1.n84 VDD1.n3 171.744
R1993 VDD1.n84 VDD1.n83 171.744
R1994 VDD1.n83 VDD1.n7 171.744
R1995 VDD1.n12 VDD1.n7 171.744
R1996 VDD1.n76 VDD1.n12 171.744
R1997 VDD1.n76 VDD1.n75 171.744
R1998 VDD1.n75 VDD1.n13 171.744
R1999 VDD1.n68 VDD1.n13 171.744
R2000 VDD1.n68 VDD1.n67 171.744
R2001 VDD1.n67 VDD1.n17 171.744
R2002 VDD1.n60 VDD1.n17 171.744
R2003 VDD1.n60 VDD1.n59 171.744
R2004 VDD1.n59 VDD1.n21 171.744
R2005 VDD1.n52 VDD1.n21 171.744
R2006 VDD1.n52 VDD1.n51 171.744
R2007 VDD1.n51 VDD1.n25 171.744
R2008 VDD1.n44 VDD1.n25 171.744
R2009 VDD1.n44 VDD1.n43 171.744
R2010 VDD1.n43 VDD1.n29 171.744
R2011 VDD1.n36 VDD1.n29 171.744
R2012 VDD1.n36 VDD1.n35 171.744
R2013 VDD1.n133 VDD1.n132 171.744
R2014 VDD1.n133 VDD1.n126 171.744
R2015 VDD1.n140 VDD1.n126 171.744
R2016 VDD1.n141 VDD1.n140 171.744
R2017 VDD1.n141 VDD1.n122 171.744
R2018 VDD1.n148 VDD1.n122 171.744
R2019 VDD1.n149 VDD1.n148 171.744
R2020 VDD1.n149 VDD1.n118 171.744
R2021 VDD1.n156 VDD1.n118 171.744
R2022 VDD1.n157 VDD1.n156 171.744
R2023 VDD1.n157 VDD1.n114 171.744
R2024 VDD1.n164 VDD1.n114 171.744
R2025 VDD1.n165 VDD1.n164 171.744
R2026 VDD1.n165 VDD1.n110 171.744
R2027 VDD1.n173 VDD1.n110 171.744
R2028 VDD1.n174 VDD1.n173 171.744
R2029 VDD1.n175 VDD1.n174 171.744
R2030 VDD1.n175 VDD1.n106 171.744
R2031 VDD1.n182 VDD1.n106 171.744
R2032 VDD1.n183 VDD1.n182 171.744
R2033 VDD1.n183 VDD1.n102 171.744
R2034 VDD1.n190 VDD1.n102 171.744
R2035 VDD1.n191 VDD1.n190 171.744
R2036 VDD1.n35 VDD1.t7 85.8723
R2037 VDD1.n132 VDD1.t6 85.8723
R2038 VDD1.n199 VDD1.n198 70.4345
R2039 VDD1.n98 VDD1.n97 67.8586
R2040 VDD1.n201 VDD1.n200 67.8584
R2041 VDD1.n197 VDD1.n196 67.8584
R2042 VDD1.n201 VDD1.n199 57.7703
R2043 VDD1.n98 VDD1.n96 51.2091
R2044 VDD1.n197 VDD1.n195 51.2091
R2045 VDD1.n34 VDD1.n33 16.3895
R2046 VDD1.n131 VDD1.n130 16.3895
R2047 VDD1.n10 VDD1.n8 13.1884
R2048 VDD1.n176 VDD1.n107 13.1884
R2049 VDD1.n82 VDD1.n81 12.8005
R2050 VDD1.n78 VDD1.n77 12.8005
R2051 VDD1.n37 VDD1.n32 12.8005
R2052 VDD1.n134 VDD1.n129 12.8005
R2053 VDD1.n177 VDD1.n109 12.8005
R2054 VDD1.n181 VDD1.n180 12.8005
R2055 VDD1.n85 VDD1.n6 12.0247
R2056 VDD1.n74 VDD1.n11 12.0247
R2057 VDD1.n38 VDD1.n30 12.0247
R2058 VDD1.n135 VDD1.n127 12.0247
R2059 VDD1.n172 VDD1.n171 12.0247
R2060 VDD1.n184 VDD1.n105 12.0247
R2061 VDD1.n86 VDD1.n4 11.249
R2062 VDD1.n73 VDD1.n14 11.249
R2063 VDD1.n42 VDD1.n41 11.249
R2064 VDD1.n139 VDD1.n138 11.249
R2065 VDD1.n170 VDD1.n111 11.249
R2066 VDD1.n185 VDD1.n103 11.249
R2067 VDD1.n90 VDD1.n89 10.4732
R2068 VDD1.n70 VDD1.n69 10.4732
R2069 VDD1.n45 VDD1.n28 10.4732
R2070 VDD1.n142 VDD1.n125 10.4732
R2071 VDD1.n167 VDD1.n166 10.4732
R2072 VDD1.n189 VDD1.n188 10.4732
R2073 VDD1.n93 VDD1.n2 9.69747
R2074 VDD1.n66 VDD1.n16 9.69747
R2075 VDD1.n46 VDD1.n26 9.69747
R2076 VDD1.n143 VDD1.n123 9.69747
R2077 VDD1.n163 VDD1.n113 9.69747
R2078 VDD1.n192 VDD1.n101 9.69747
R2079 VDD1.n96 VDD1.n95 9.45567
R2080 VDD1.n195 VDD1.n194 9.45567
R2081 VDD1.n20 VDD1.n19 9.3005
R2082 VDD1.n63 VDD1.n62 9.3005
R2083 VDD1.n65 VDD1.n64 9.3005
R2084 VDD1.n16 VDD1.n15 9.3005
R2085 VDD1.n71 VDD1.n70 9.3005
R2086 VDD1.n73 VDD1.n72 9.3005
R2087 VDD1.n11 VDD1.n9 9.3005
R2088 VDD1.n79 VDD1.n78 9.3005
R2089 VDD1.n95 VDD1.n94 9.3005
R2090 VDD1.n2 VDD1.n1 9.3005
R2091 VDD1.n89 VDD1.n88 9.3005
R2092 VDD1.n87 VDD1.n86 9.3005
R2093 VDD1.n6 VDD1.n5 9.3005
R2094 VDD1.n81 VDD1.n80 9.3005
R2095 VDD1.n57 VDD1.n56 9.3005
R2096 VDD1.n55 VDD1.n54 9.3005
R2097 VDD1.n24 VDD1.n23 9.3005
R2098 VDD1.n49 VDD1.n48 9.3005
R2099 VDD1.n47 VDD1.n46 9.3005
R2100 VDD1.n28 VDD1.n27 9.3005
R2101 VDD1.n41 VDD1.n40 9.3005
R2102 VDD1.n39 VDD1.n38 9.3005
R2103 VDD1.n32 VDD1.n31 9.3005
R2104 VDD1.n194 VDD1.n193 9.3005
R2105 VDD1.n101 VDD1.n100 9.3005
R2106 VDD1.n188 VDD1.n187 9.3005
R2107 VDD1.n186 VDD1.n185 9.3005
R2108 VDD1.n105 VDD1.n104 9.3005
R2109 VDD1.n180 VDD1.n179 9.3005
R2110 VDD1.n152 VDD1.n151 9.3005
R2111 VDD1.n121 VDD1.n120 9.3005
R2112 VDD1.n146 VDD1.n145 9.3005
R2113 VDD1.n144 VDD1.n143 9.3005
R2114 VDD1.n125 VDD1.n124 9.3005
R2115 VDD1.n138 VDD1.n137 9.3005
R2116 VDD1.n136 VDD1.n135 9.3005
R2117 VDD1.n129 VDD1.n128 9.3005
R2118 VDD1.n154 VDD1.n153 9.3005
R2119 VDD1.n117 VDD1.n116 9.3005
R2120 VDD1.n160 VDD1.n159 9.3005
R2121 VDD1.n162 VDD1.n161 9.3005
R2122 VDD1.n113 VDD1.n112 9.3005
R2123 VDD1.n168 VDD1.n167 9.3005
R2124 VDD1.n170 VDD1.n169 9.3005
R2125 VDD1.n171 VDD1.n108 9.3005
R2126 VDD1.n178 VDD1.n177 9.3005
R2127 VDD1.n94 VDD1.n0 8.92171
R2128 VDD1.n65 VDD1.n18 8.92171
R2129 VDD1.n50 VDD1.n49 8.92171
R2130 VDD1.n147 VDD1.n146 8.92171
R2131 VDD1.n162 VDD1.n115 8.92171
R2132 VDD1.n193 VDD1.n99 8.92171
R2133 VDD1.n62 VDD1.n61 8.14595
R2134 VDD1.n53 VDD1.n24 8.14595
R2135 VDD1.n150 VDD1.n121 8.14595
R2136 VDD1.n159 VDD1.n158 8.14595
R2137 VDD1.n58 VDD1.n20 7.3702
R2138 VDD1.n54 VDD1.n22 7.3702
R2139 VDD1.n151 VDD1.n119 7.3702
R2140 VDD1.n155 VDD1.n117 7.3702
R2141 VDD1.n58 VDD1.n57 6.59444
R2142 VDD1.n57 VDD1.n22 6.59444
R2143 VDD1.n154 VDD1.n119 6.59444
R2144 VDD1.n155 VDD1.n154 6.59444
R2145 VDD1.n61 VDD1.n20 5.81868
R2146 VDD1.n54 VDD1.n53 5.81868
R2147 VDD1.n151 VDD1.n150 5.81868
R2148 VDD1.n158 VDD1.n117 5.81868
R2149 VDD1.n96 VDD1.n0 5.04292
R2150 VDD1.n62 VDD1.n18 5.04292
R2151 VDD1.n50 VDD1.n24 5.04292
R2152 VDD1.n147 VDD1.n121 5.04292
R2153 VDD1.n159 VDD1.n115 5.04292
R2154 VDD1.n195 VDD1.n99 5.04292
R2155 VDD1.n94 VDD1.n93 4.26717
R2156 VDD1.n66 VDD1.n65 4.26717
R2157 VDD1.n49 VDD1.n26 4.26717
R2158 VDD1.n146 VDD1.n123 4.26717
R2159 VDD1.n163 VDD1.n162 4.26717
R2160 VDD1.n193 VDD1.n192 4.26717
R2161 VDD1.n33 VDD1.n31 3.70982
R2162 VDD1.n130 VDD1.n128 3.70982
R2163 VDD1.n90 VDD1.n2 3.49141
R2164 VDD1.n69 VDD1.n16 3.49141
R2165 VDD1.n46 VDD1.n45 3.49141
R2166 VDD1.n143 VDD1.n142 3.49141
R2167 VDD1.n166 VDD1.n113 3.49141
R2168 VDD1.n189 VDD1.n101 3.49141
R2169 VDD1.n89 VDD1.n4 2.71565
R2170 VDD1.n70 VDD1.n14 2.71565
R2171 VDD1.n42 VDD1.n28 2.71565
R2172 VDD1.n139 VDD1.n125 2.71565
R2173 VDD1.n167 VDD1.n111 2.71565
R2174 VDD1.n188 VDD1.n103 2.71565
R2175 VDD1 VDD1.n201 2.57378
R2176 VDD1.n86 VDD1.n85 1.93989
R2177 VDD1.n74 VDD1.n73 1.93989
R2178 VDD1.n41 VDD1.n30 1.93989
R2179 VDD1.n138 VDD1.n127 1.93989
R2180 VDD1.n172 VDD1.n170 1.93989
R2181 VDD1.n185 VDD1.n184 1.93989
R2182 VDD1.n200 VDD1.t4 1.86218
R2183 VDD1.n200 VDD1.t2 1.86218
R2184 VDD1.n97 VDD1.t9 1.86218
R2185 VDD1.n97 VDD1.t8 1.86218
R2186 VDD1.n198 VDD1.t1 1.86218
R2187 VDD1.n198 VDD1.t0 1.86218
R2188 VDD1.n196 VDD1.t3 1.86218
R2189 VDD1.n196 VDD1.t5 1.86218
R2190 VDD1.n82 VDD1.n6 1.16414
R2191 VDD1.n77 VDD1.n11 1.16414
R2192 VDD1.n38 VDD1.n37 1.16414
R2193 VDD1.n135 VDD1.n134 1.16414
R2194 VDD1.n171 VDD1.n109 1.16414
R2195 VDD1.n181 VDD1.n105 1.16414
R2196 VDD1 VDD1.n98 0.935845
R2197 VDD1.n199 VDD1.n197 0.822309
R2198 VDD1.n81 VDD1.n8 0.388379
R2199 VDD1.n78 VDD1.n10 0.388379
R2200 VDD1.n34 VDD1.n32 0.388379
R2201 VDD1.n131 VDD1.n129 0.388379
R2202 VDD1.n177 VDD1.n176 0.388379
R2203 VDD1.n180 VDD1.n107 0.388379
R2204 VDD1.n95 VDD1.n1 0.155672
R2205 VDD1.n88 VDD1.n1 0.155672
R2206 VDD1.n88 VDD1.n87 0.155672
R2207 VDD1.n87 VDD1.n5 0.155672
R2208 VDD1.n80 VDD1.n5 0.155672
R2209 VDD1.n80 VDD1.n79 0.155672
R2210 VDD1.n79 VDD1.n9 0.155672
R2211 VDD1.n72 VDD1.n9 0.155672
R2212 VDD1.n72 VDD1.n71 0.155672
R2213 VDD1.n71 VDD1.n15 0.155672
R2214 VDD1.n64 VDD1.n15 0.155672
R2215 VDD1.n64 VDD1.n63 0.155672
R2216 VDD1.n63 VDD1.n19 0.155672
R2217 VDD1.n56 VDD1.n19 0.155672
R2218 VDD1.n56 VDD1.n55 0.155672
R2219 VDD1.n55 VDD1.n23 0.155672
R2220 VDD1.n48 VDD1.n23 0.155672
R2221 VDD1.n48 VDD1.n47 0.155672
R2222 VDD1.n47 VDD1.n27 0.155672
R2223 VDD1.n40 VDD1.n27 0.155672
R2224 VDD1.n40 VDD1.n39 0.155672
R2225 VDD1.n39 VDD1.n31 0.155672
R2226 VDD1.n136 VDD1.n128 0.155672
R2227 VDD1.n137 VDD1.n136 0.155672
R2228 VDD1.n137 VDD1.n124 0.155672
R2229 VDD1.n144 VDD1.n124 0.155672
R2230 VDD1.n145 VDD1.n144 0.155672
R2231 VDD1.n145 VDD1.n120 0.155672
R2232 VDD1.n152 VDD1.n120 0.155672
R2233 VDD1.n153 VDD1.n152 0.155672
R2234 VDD1.n153 VDD1.n116 0.155672
R2235 VDD1.n160 VDD1.n116 0.155672
R2236 VDD1.n161 VDD1.n160 0.155672
R2237 VDD1.n161 VDD1.n112 0.155672
R2238 VDD1.n168 VDD1.n112 0.155672
R2239 VDD1.n169 VDD1.n168 0.155672
R2240 VDD1.n169 VDD1.n108 0.155672
R2241 VDD1.n178 VDD1.n108 0.155672
R2242 VDD1.n179 VDD1.n178 0.155672
R2243 VDD1.n179 VDD1.n104 0.155672
R2244 VDD1.n186 VDD1.n104 0.155672
R2245 VDD1.n187 VDD1.n186 0.155672
R2246 VDD1.n187 VDD1.n100 0.155672
R2247 VDD1.n194 VDD1.n100 0.155672
R2248 VTAIL.n400 VTAIL.n308 756.745
R2249 VTAIL.n94 VTAIL.n2 756.745
R2250 VTAIL.n302 VTAIL.n210 756.745
R2251 VTAIL.n200 VTAIL.n108 756.745
R2252 VTAIL.n341 VTAIL.n340 585
R2253 VTAIL.n343 VTAIL.n342 585
R2254 VTAIL.n336 VTAIL.n335 585
R2255 VTAIL.n349 VTAIL.n348 585
R2256 VTAIL.n351 VTAIL.n350 585
R2257 VTAIL.n332 VTAIL.n331 585
R2258 VTAIL.n357 VTAIL.n356 585
R2259 VTAIL.n359 VTAIL.n358 585
R2260 VTAIL.n328 VTAIL.n327 585
R2261 VTAIL.n365 VTAIL.n364 585
R2262 VTAIL.n367 VTAIL.n366 585
R2263 VTAIL.n324 VTAIL.n323 585
R2264 VTAIL.n373 VTAIL.n372 585
R2265 VTAIL.n375 VTAIL.n374 585
R2266 VTAIL.n320 VTAIL.n319 585
R2267 VTAIL.n382 VTAIL.n381 585
R2268 VTAIL.n383 VTAIL.n318 585
R2269 VTAIL.n385 VTAIL.n384 585
R2270 VTAIL.n316 VTAIL.n315 585
R2271 VTAIL.n391 VTAIL.n390 585
R2272 VTAIL.n393 VTAIL.n392 585
R2273 VTAIL.n312 VTAIL.n311 585
R2274 VTAIL.n399 VTAIL.n398 585
R2275 VTAIL.n401 VTAIL.n400 585
R2276 VTAIL.n35 VTAIL.n34 585
R2277 VTAIL.n37 VTAIL.n36 585
R2278 VTAIL.n30 VTAIL.n29 585
R2279 VTAIL.n43 VTAIL.n42 585
R2280 VTAIL.n45 VTAIL.n44 585
R2281 VTAIL.n26 VTAIL.n25 585
R2282 VTAIL.n51 VTAIL.n50 585
R2283 VTAIL.n53 VTAIL.n52 585
R2284 VTAIL.n22 VTAIL.n21 585
R2285 VTAIL.n59 VTAIL.n58 585
R2286 VTAIL.n61 VTAIL.n60 585
R2287 VTAIL.n18 VTAIL.n17 585
R2288 VTAIL.n67 VTAIL.n66 585
R2289 VTAIL.n69 VTAIL.n68 585
R2290 VTAIL.n14 VTAIL.n13 585
R2291 VTAIL.n76 VTAIL.n75 585
R2292 VTAIL.n77 VTAIL.n12 585
R2293 VTAIL.n79 VTAIL.n78 585
R2294 VTAIL.n10 VTAIL.n9 585
R2295 VTAIL.n85 VTAIL.n84 585
R2296 VTAIL.n87 VTAIL.n86 585
R2297 VTAIL.n6 VTAIL.n5 585
R2298 VTAIL.n93 VTAIL.n92 585
R2299 VTAIL.n95 VTAIL.n94 585
R2300 VTAIL.n303 VTAIL.n302 585
R2301 VTAIL.n301 VTAIL.n300 585
R2302 VTAIL.n214 VTAIL.n213 585
R2303 VTAIL.n295 VTAIL.n294 585
R2304 VTAIL.n293 VTAIL.n292 585
R2305 VTAIL.n218 VTAIL.n217 585
R2306 VTAIL.n222 VTAIL.n220 585
R2307 VTAIL.n287 VTAIL.n286 585
R2308 VTAIL.n285 VTAIL.n284 585
R2309 VTAIL.n224 VTAIL.n223 585
R2310 VTAIL.n279 VTAIL.n278 585
R2311 VTAIL.n277 VTAIL.n276 585
R2312 VTAIL.n228 VTAIL.n227 585
R2313 VTAIL.n271 VTAIL.n270 585
R2314 VTAIL.n269 VTAIL.n268 585
R2315 VTAIL.n232 VTAIL.n231 585
R2316 VTAIL.n263 VTAIL.n262 585
R2317 VTAIL.n261 VTAIL.n260 585
R2318 VTAIL.n236 VTAIL.n235 585
R2319 VTAIL.n255 VTAIL.n254 585
R2320 VTAIL.n253 VTAIL.n252 585
R2321 VTAIL.n240 VTAIL.n239 585
R2322 VTAIL.n247 VTAIL.n246 585
R2323 VTAIL.n245 VTAIL.n244 585
R2324 VTAIL.n201 VTAIL.n200 585
R2325 VTAIL.n199 VTAIL.n198 585
R2326 VTAIL.n112 VTAIL.n111 585
R2327 VTAIL.n193 VTAIL.n192 585
R2328 VTAIL.n191 VTAIL.n190 585
R2329 VTAIL.n116 VTAIL.n115 585
R2330 VTAIL.n120 VTAIL.n118 585
R2331 VTAIL.n185 VTAIL.n184 585
R2332 VTAIL.n183 VTAIL.n182 585
R2333 VTAIL.n122 VTAIL.n121 585
R2334 VTAIL.n177 VTAIL.n176 585
R2335 VTAIL.n175 VTAIL.n174 585
R2336 VTAIL.n126 VTAIL.n125 585
R2337 VTAIL.n169 VTAIL.n168 585
R2338 VTAIL.n167 VTAIL.n166 585
R2339 VTAIL.n130 VTAIL.n129 585
R2340 VTAIL.n161 VTAIL.n160 585
R2341 VTAIL.n159 VTAIL.n158 585
R2342 VTAIL.n134 VTAIL.n133 585
R2343 VTAIL.n153 VTAIL.n152 585
R2344 VTAIL.n151 VTAIL.n150 585
R2345 VTAIL.n138 VTAIL.n137 585
R2346 VTAIL.n145 VTAIL.n144 585
R2347 VTAIL.n143 VTAIL.n142 585
R2348 VTAIL.n339 VTAIL.t0 327.466
R2349 VTAIL.n33 VTAIL.t16 327.466
R2350 VTAIL.n243 VTAIL.t18 327.466
R2351 VTAIL.n141 VTAIL.t4 327.466
R2352 VTAIL.n342 VTAIL.n341 171.744
R2353 VTAIL.n342 VTAIL.n335 171.744
R2354 VTAIL.n349 VTAIL.n335 171.744
R2355 VTAIL.n350 VTAIL.n349 171.744
R2356 VTAIL.n350 VTAIL.n331 171.744
R2357 VTAIL.n357 VTAIL.n331 171.744
R2358 VTAIL.n358 VTAIL.n357 171.744
R2359 VTAIL.n358 VTAIL.n327 171.744
R2360 VTAIL.n365 VTAIL.n327 171.744
R2361 VTAIL.n366 VTAIL.n365 171.744
R2362 VTAIL.n366 VTAIL.n323 171.744
R2363 VTAIL.n373 VTAIL.n323 171.744
R2364 VTAIL.n374 VTAIL.n373 171.744
R2365 VTAIL.n374 VTAIL.n319 171.744
R2366 VTAIL.n382 VTAIL.n319 171.744
R2367 VTAIL.n383 VTAIL.n382 171.744
R2368 VTAIL.n384 VTAIL.n383 171.744
R2369 VTAIL.n384 VTAIL.n315 171.744
R2370 VTAIL.n391 VTAIL.n315 171.744
R2371 VTAIL.n392 VTAIL.n391 171.744
R2372 VTAIL.n392 VTAIL.n311 171.744
R2373 VTAIL.n399 VTAIL.n311 171.744
R2374 VTAIL.n400 VTAIL.n399 171.744
R2375 VTAIL.n36 VTAIL.n35 171.744
R2376 VTAIL.n36 VTAIL.n29 171.744
R2377 VTAIL.n43 VTAIL.n29 171.744
R2378 VTAIL.n44 VTAIL.n43 171.744
R2379 VTAIL.n44 VTAIL.n25 171.744
R2380 VTAIL.n51 VTAIL.n25 171.744
R2381 VTAIL.n52 VTAIL.n51 171.744
R2382 VTAIL.n52 VTAIL.n21 171.744
R2383 VTAIL.n59 VTAIL.n21 171.744
R2384 VTAIL.n60 VTAIL.n59 171.744
R2385 VTAIL.n60 VTAIL.n17 171.744
R2386 VTAIL.n67 VTAIL.n17 171.744
R2387 VTAIL.n68 VTAIL.n67 171.744
R2388 VTAIL.n68 VTAIL.n13 171.744
R2389 VTAIL.n76 VTAIL.n13 171.744
R2390 VTAIL.n77 VTAIL.n76 171.744
R2391 VTAIL.n78 VTAIL.n77 171.744
R2392 VTAIL.n78 VTAIL.n9 171.744
R2393 VTAIL.n85 VTAIL.n9 171.744
R2394 VTAIL.n86 VTAIL.n85 171.744
R2395 VTAIL.n86 VTAIL.n5 171.744
R2396 VTAIL.n93 VTAIL.n5 171.744
R2397 VTAIL.n94 VTAIL.n93 171.744
R2398 VTAIL.n302 VTAIL.n301 171.744
R2399 VTAIL.n301 VTAIL.n213 171.744
R2400 VTAIL.n294 VTAIL.n213 171.744
R2401 VTAIL.n294 VTAIL.n293 171.744
R2402 VTAIL.n293 VTAIL.n217 171.744
R2403 VTAIL.n222 VTAIL.n217 171.744
R2404 VTAIL.n286 VTAIL.n222 171.744
R2405 VTAIL.n286 VTAIL.n285 171.744
R2406 VTAIL.n285 VTAIL.n223 171.744
R2407 VTAIL.n278 VTAIL.n223 171.744
R2408 VTAIL.n278 VTAIL.n277 171.744
R2409 VTAIL.n277 VTAIL.n227 171.744
R2410 VTAIL.n270 VTAIL.n227 171.744
R2411 VTAIL.n270 VTAIL.n269 171.744
R2412 VTAIL.n269 VTAIL.n231 171.744
R2413 VTAIL.n262 VTAIL.n231 171.744
R2414 VTAIL.n262 VTAIL.n261 171.744
R2415 VTAIL.n261 VTAIL.n235 171.744
R2416 VTAIL.n254 VTAIL.n235 171.744
R2417 VTAIL.n254 VTAIL.n253 171.744
R2418 VTAIL.n253 VTAIL.n239 171.744
R2419 VTAIL.n246 VTAIL.n239 171.744
R2420 VTAIL.n246 VTAIL.n245 171.744
R2421 VTAIL.n200 VTAIL.n199 171.744
R2422 VTAIL.n199 VTAIL.n111 171.744
R2423 VTAIL.n192 VTAIL.n111 171.744
R2424 VTAIL.n192 VTAIL.n191 171.744
R2425 VTAIL.n191 VTAIL.n115 171.744
R2426 VTAIL.n120 VTAIL.n115 171.744
R2427 VTAIL.n184 VTAIL.n120 171.744
R2428 VTAIL.n184 VTAIL.n183 171.744
R2429 VTAIL.n183 VTAIL.n121 171.744
R2430 VTAIL.n176 VTAIL.n121 171.744
R2431 VTAIL.n176 VTAIL.n175 171.744
R2432 VTAIL.n175 VTAIL.n125 171.744
R2433 VTAIL.n168 VTAIL.n125 171.744
R2434 VTAIL.n168 VTAIL.n167 171.744
R2435 VTAIL.n167 VTAIL.n129 171.744
R2436 VTAIL.n160 VTAIL.n129 171.744
R2437 VTAIL.n160 VTAIL.n159 171.744
R2438 VTAIL.n159 VTAIL.n133 171.744
R2439 VTAIL.n152 VTAIL.n133 171.744
R2440 VTAIL.n152 VTAIL.n151 171.744
R2441 VTAIL.n151 VTAIL.n137 171.744
R2442 VTAIL.n144 VTAIL.n137 171.744
R2443 VTAIL.n144 VTAIL.n143 171.744
R2444 VTAIL.n341 VTAIL.t0 85.8723
R2445 VTAIL.n35 VTAIL.t16 85.8723
R2446 VTAIL.n245 VTAIL.t18 85.8723
R2447 VTAIL.n143 VTAIL.t4 85.8723
R2448 VTAIL.n209 VTAIL.n208 51.1798
R2449 VTAIL.n207 VTAIL.n206 51.1798
R2450 VTAIL.n107 VTAIL.n106 51.1798
R2451 VTAIL.n105 VTAIL.n104 51.1798
R2452 VTAIL.n407 VTAIL.n406 51.1796
R2453 VTAIL.n1 VTAIL.n0 51.1796
R2454 VTAIL.n101 VTAIL.n100 51.1796
R2455 VTAIL.n103 VTAIL.n102 51.1796
R2456 VTAIL.n105 VTAIL.n103 34.4358
R2457 VTAIL.n405 VTAIL.n404 31.0217
R2458 VTAIL.n99 VTAIL.n98 31.0217
R2459 VTAIL.n307 VTAIL.n306 31.0217
R2460 VTAIL.n205 VTAIL.n204 31.0217
R2461 VTAIL.n405 VTAIL.n307 30.9272
R2462 VTAIL.n340 VTAIL.n339 16.3895
R2463 VTAIL.n34 VTAIL.n33 16.3895
R2464 VTAIL.n244 VTAIL.n243 16.3895
R2465 VTAIL.n142 VTAIL.n141 16.3895
R2466 VTAIL.n385 VTAIL.n316 13.1884
R2467 VTAIL.n79 VTAIL.n10 13.1884
R2468 VTAIL.n220 VTAIL.n218 13.1884
R2469 VTAIL.n118 VTAIL.n116 13.1884
R2470 VTAIL.n343 VTAIL.n338 12.8005
R2471 VTAIL.n386 VTAIL.n318 12.8005
R2472 VTAIL.n390 VTAIL.n389 12.8005
R2473 VTAIL.n37 VTAIL.n32 12.8005
R2474 VTAIL.n80 VTAIL.n12 12.8005
R2475 VTAIL.n84 VTAIL.n83 12.8005
R2476 VTAIL.n292 VTAIL.n291 12.8005
R2477 VTAIL.n288 VTAIL.n287 12.8005
R2478 VTAIL.n247 VTAIL.n242 12.8005
R2479 VTAIL.n190 VTAIL.n189 12.8005
R2480 VTAIL.n186 VTAIL.n185 12.8005
R2481 VTAIL.n145 VTAIL.n140 12.8005
R2482 VTAIL.n344 VTAIL.n336 12.0247
R2483 VTAIL.n381 VTAIL.n380 12.0247
R2484 VTAIL.n393 VTAIL.n314 12.0247
R2485 VTAIL.n38 VTAIL.n30 12.0247
R2486 VTAIL.n75 VTAIL.n74 12.0247
R2487 VTAIL.n87 VTAIL.n8 12.0247
R2488 VTAIL.n295 VTAIL.n216 12.0247
R2489 VTAIL.n284 VTAIL.n221 12.0247
R2490 VTAIL.n248 VTAIL.n240 12.0247
R2491 VTAIL.n193 VTAIL.n114 12.0247
R2492 VTAIL.n182 VTAIL.n119 12.0247
R2493 VTAIL.n146 VTAIL.n138 12.0247
R2494 VTAIL.n348 VTAIL.n347 11.249
R2495 VTAIL.n379 VTAIL.n320 11.249
R2496 VTAIL.n394 VTAIL.n312 11.249
R2497 VTAIL.n42 VTAIL.n41 11.249
R2498 VTAIL.n73 VTAIL.n14 11.249
R2499 VTAIL.n88 VTAIL.n6 11.249
R2500 VTAIL.n296 VTAIL.n214 11.249
R2501 VTAIL.n283 VTAIL.n224 11.249
R2502 VTAIL.n252 VTAIL.n251 11.249
R2503 VTAIL.n194 VTAIL.n112 11.249
R2504 VTAIL.n181 VTAIL.n122 11.249
R2505 VTAIL.n150 VTAIL.n149 11.249
R2506 VTAIL.n351 VTAIL.n334 10.4732
R2507 VTAIL.n376 VTAIL.n375 10.4732
R2508 VTAIL.n398 VTAIL.n397 10.4732
R2509 VTAIL.n45 VTAIL.n28 10.4732
R2510 VTAIL.n70 VTAIL.n69 10.4732
R2511 VTAIL.n92 VTAIL.n91 10.4732
R2512 VTAIL.n300 VTAIL.n299 10.4732
R2513 VTAIL.n280 VTAIL.n279 10.4732
R2514 VTAIL.n255 VTAIL.n238 10.4732
R2515 VTAIL.n198 VTAIL.n197 10.4732
R2516 VTAIL.n178 VTAIL.n177 10.4732
R2517 VTAIL.n153 VTAIL.n136 10.4732
R2518 VTAIL.n352 VTAIL.n332 9.69747
R2519 VTAIL.n372 VTAIL.n322 9.69747
R2520 VTAIL.n401 VTAIL.n310 9.69747
R2521 VTAIL.n46 VTAIL.n26 9.69747
R2522 VTAIL.n66 VTAIL.n16 9.69747
R2523 VTAIL.n95 VTAIL.n4 9.69747
R2524 VTAIL.n303 VTAIL.n212 9.69747
R2525 VTAIL.n276 VTAIL.n226 9.69747
R2526 VTAIL.n256 VTAIL.n236 9.69747
R2527 VTAIL.n201 VTAIL.n110 9.69747
R2528 VTAIL.n174 VTAIL.n124 9.69747
R2529 VTAIL.n154 VTAIL.n134 9.69747
R2530 VTAIL.n404 VTAIL.n403 9.45567
R2531 VTAIL.n98 VTAIL.n97 9.45567
R2532 VTAIL.n306 VTAIL.n305 9.45567
R2533 VTAIL.n204 VTAIL.n203 9.45567
R2534 VTAIL.n403 VTAIL.n402 9.3005
R2535 VTAIL.n310 VTAIL.n309 9.3005
R2536 VTAIL.n397 VTAIL.n396 9.3005
R2537 VTAIL.n395 VTAIL.n394 9.3005
R2538 VTAIL.n314 VTAIL.n313 9.3005
R2539 VTAIL.n389 VTAIL.n388 9.3005
R2540 VTAIL.n361 VTAIL.n360 9.3005
R2541 VTAIL.n330 VTAIL.n329 9.3005
R2542 VTAIL.n355 VTAIL.n354 9.3005
R2543 VTAIL.n353 VTAIL.n352 9.3005
R2544 VTAIL.n334 VTAIL.n333 9.3005
R2545 VTAIL.n347 VTAIL.n346 9.3005
R2546 VTAIL.n345 VTAIL.n344 9.3005
R2547 VTAIL.n338 VTAIL.n337 9.3005
R2548 VTAIL.n363 VTAIL.n362 9.3005
R2549 VTAIL.n326 VTAIL.n325 9.3005
R2550 VTAIL.n369 VTAIL.n368 9.3005
R2551 VTAIL.n371 VTAIL.n370 9.3005
R2552 VTAIL.n322 VTAIL.n321 9.3005
R2553 VTAIL.n377 VTAIL.n376 9.3005
R2554 VTAIL.n379 VTAIL.n378 9.3005
R2555 VTAIL.n380 VTAIL.n317 9.3005
R2556 VTAIL.n387 VTAIL.n386 9.3005
R2557 VTAIL.n97 VTAIL.n96 9.3005
R2558 VTAIL.n4 VTAIL.n3 9.3005
R2559 VTAIL.n91 VTAIL.n90 9.3005
R2560 VTAIL.n89 VTAIL.n88 9.3005
R2561 VTAIL.n8 VTAIL.n7 9.3005
R2562 VTAIL.n83 VTAIL.n82 9.3005
R2563 VTAIL.n55 VTAIL.n54 9.3005
R2564 VTAIL.n24 VTAIL.n23 9.3005
R2565 VTAIL.n49 VTAIL.n48 9.3005
R2566 VTAIL.n47 VTAIL.n46 9.3005
R2567 VTAIL.n28 VTAIL.n27 9.3005
R2568 VTAIL.n41 VTAIL.n40 9.3005
R2569 VTAIL.n39 VTAIL.n38 9.3005
R2570 VTAIL.n32 VTAIL.n31 9.3005
R2571 VTAIL.n57 VTAIL.n56 9.3005
R2572 VTAIL.n20 VTAIL.n19 9.3005
R2573 VTAIL.n63 VTAIL.n62 9.3005
R2574 VTAIL.n65 VTAIL.n64 9.3005
R2575 VTAIL.n16 VTAIL.n15 9.3005
R2576 VTAIL.n71 VTAIL.n70 9.3005
R2577 VTAIL.n73 VTAIL.n72 9.3005
R2578 VTAIL.n74 VTAIL.n11 9.3005
R2579 VTAIL.n81 VTAIL.n80 9.3005
R2580 VTAIL.n230 VTAIL.n229 9.3005
R2581 VTAIL.n273 VTAIL.n272 9.3005
R2582 VTAIL.n275 VTAIL.n274 9.3005
R2583 VTAIL.n226 VTAIL.n225 9.3005
R2584 VTAIL.n281 VTAIL.n280 9.3005
R2585 VTAIL.n283 VTAIL.n282 9.3005
R2586 VTAIL.n221 VTAIL.n219 9.3005
R2587 VTAIL.n289 VTAIL.n288 9.3005
R2588 VTAIL.n305 VTAIL.n304 9.3005
R2589 VTAIL.n212 VTAIL.n211 9.3005
R2590 VTAIL.n299 VTAIL.n298 9.3005
R2591 VTAIL.n297 VTAIL.n296 9.3005
R2592 VTAIL.n216 VTAIL.n215 9.3005
R2593 VTAIL.n291 VTAIL.n290 9.3005
R2594 VTAIL.n267 VTAIL.n266 9.3005
R2595 VTAIL.n265 VTAIL.n264 9.3005
R2596 VTAIL.n234 VTAIL.n233 9.3005
R2597 VTAIL.n259 VTAIL.n258 9.3005
R2598 VTAIL.n257 VTAIL.n256 9.3005
R2599 VTAIL.n238 VTAIL.n237 9.3005
R2600 VTAIL.n251 VTAIL.n250 9.3005
R2601 VTAIL.n249 VTAIL.n248 9.3005
R2602 VTAIL.n242 VTAIL.n241 9.3005
R2603 VTAIL.n128 VTAIL.n127 9.3005
R2604 VTAIL.n171 VTAIL.n170 9.3005
R2605 VTAIL.n173 VTAIL.n172 9.3005
R2606 VTAIL.n124 VTAIL.n123 9.3005
R2607 VTAIL.n179 VTAIL.n178 9.3005
R2608 VTAIL.n181 VTAIL.n180 9.3005
R2609 VTAIL.n119 VTAIL.n117 9.3005
R2610 VTAIL.n187 VTAIL.n186 9.3005
R2611 VTAIL.n203 VTAIL.n202 9.3005
R2612 VTAIL.n110 VTAIL.n109 9.3005
R2613 VTAIL.n197 VTAIL.n196 9.3005
R2614 VTAIL.n195 VTAIL.n194 9.3005
R2615 VTAIL.n114 VTAIL.n113 9.3005
R2616 VTAIL.n189 VTAIL.n188 9.3005
R2617 VTAIL.n165 VTAIL.n164 9.3005
R2618 VTAIL.n163 VTAIL.n162 9.3005
R2619 VTAIL.n132 VTAIL.n131 9.3005
R2620 VTAIL.n157 VTAIL.n156 9.3005
R2621 VTAIL.n155 VTAIL.n154 9.3005
R2622 VTAIL.n136 VTAIL.n135 9.3005
R2623 VTAIL.n149 VTAIL.n148 9.3005
R2624 VTAIL.n147 VTAIL.n146 9.3005
R2625 VTAIL.n140 VTAIL.n139 9.3005
R2626 VTAIL.n356 VTAIL.n355 8.92171
R2627 VTAIL.n371 VTAIL.n324 8.92171
R2628 VTAIL.n402 VTAIL.n308 8.92171
R2629 VTAIL.n50 VTAIL.n49 8.92171
R2630 VTAIL.n65 VTAIL.n18 8.92171
R2631 VTAIL.n96 VTAIL.n2 8.92171
R2632 VTAIL.n304 VTAIL.n210 8.92171
R2633 VTAIL.n275 VTAIL.n228 8.92171
R2634 VTAIL.n260 VTAIL.n259 8.92171
R2635 VTAIL.n202 VTAIL.n108 8.92171
R2636 VTAIL.n173 VTAIL.n126 8.92171
R2637 VTAIL.n158 VTAIL.n157 8.92171
R2638 VTAIL.n359 VTAIL.n330 8.14595
R2639 VTAIL.n368 VTAIL.n367 8.14595
R2640 VTAIL.n53 VTAIL.n24 8.14595
R2641 VTAIL.n62 VTAIL.n61 8.14595
R2642 VTAIL.n272 VTAIL.n271 8.14595
R2643 VTAIL.n263 VTAIL.n234 8.14595
R2644 VTAIL.n170 VTAIL.n169 8.14595
R2645 VTAIL.n161 VTAIL.n132 8.14595
R2646 VTAIL.n360 VTAIL.n328 7.3702
R2647 VTAIL.n364 VTAIL.n326 7.3702
R2648 VTAIL.n54 VTAIL.n22 7.3702
R2649 VTAIL.n58 VTAIL.n20 7.3702
R2650 VTAIL.n268 VTAIL.n230 7.3702
R2651 VTAIL.n264 VTAIL.n232 7.3702
R2652 VTAIL.n166 VTAIL.n128 7.3702
R2653 VTAIL.n162 VTAIL.n130 7.3702
R2654 VTAIL.n363 VTAIL.n328 6.59444
R2655 VTAIL.n364 VTAIL.n363 6.59444
R2656 VTAIL.n57 VTAIL.n22 6.59444
R2657 VTAIL.n58 VTAIL.n57 6.59444
R2658 VTAIL.n268 VTAIL.n267 6.59444
R2659 VTAIL.n267 VTAIL.n232 6.59444
R2660 VTAIL.n166 VTAIL.n165 6.59444
R2661 VTAIL.n165 VTAIL.n130 6.59444
R2662 VTAIL.n360 VTAIL.n359 5.81868
R2663 VTAIL.n367 VTAIL.n326 5.81868
R2664 VTAIL.n54 VTAIL.n53 5.81868
R2665 VTAIL.n61 VTAIL.n20 5.81868
R2666 VTAIL.n271 VTAIL.n230 5.81868
R2667 VTAIL.n264 VTAIL.n263 5.81868
R2668 VTAIL.n169 VTAIL.n128 5.81868
R2669 VTAIL.n162 VTAIL.n161 5.81868
R2670 VTAIL.n356 VTAIL.n330 5.04292
R2671 VTAIL.n368 VTAIL.n324 5.04292
R2672 VTAIL.n404 VTAIL.n308 5.04292
R2673 VTAIL.n50 VTAIL.n24 5.04292
R2674 VTAIL.n62 VTAIL.n18 5.04292
R2675 VTAIL.n98 VTAIL.n2 5.04292
R2676 VTAIL.n306 VTAIL.n210 5.04292
R2677 VTAIL.n272 VTAIL.n228 5.04292
R2678 VTAIL.n260 VTAIL.n234 5.04292
R2679 VTAIL.n204 VTAIL.n108 5.04292
R2680 VTAIL.n170 VTAIL.n126 5.04292
R2681 VTAIL.n158 VTAIL.n132 5.04292
R2682 VTAIL.n355 VTAIL.n332 4.26717
R2683 VTAIL.n372 VTAIL.n371 4.26717
R2684 VTAIL.n402 VTAIL.n401 4.26717
R2685 VTAIL.n49 VTAIL.n26 4.26717
R2686 VTAIL.n66 VTAIL.n65 4.26717
R2687 VTAIL.n96 VTAIL.n95 4.26717
R2688 VTAIL.n304 VTAIL.n303 4.26717
R2689 VTAIL.n276 VTAIL.n275 4.26717
R2690 VTAIL.n259 VTAIL.n236 4.26717
R2691 VTAIL.n202 VTAIL.n201 4.26717
R2692 VTAIL.n174 VTAIL.n173 4.26717
R2693 VTAIL.n157 VTAIL.n134 4.26717
R2694 VTAIL.n339 VTAIL.n337 3.70982
R2695 VTAIL.n33 VTAIL.n31 3.70982
R2696 VTAIL.n243 VTAIL.n241 3.70982
R2697 VTAIL.n141 VTAIL.n139 3.70982
R2698 VTAIL.n107 VTAIL.n105 3.50912
R2699 VTAIL.n205 VTAIL.n107 3.50912
R2700 VTAIL.n209 VTAIL.n207 3.50912
R2701 VTAIL.n307 VTAIL.n209 3.50912
R2702 VTAIL.n103 VTAIL.n101 3.50912
R2703 VTAIL.n101 VTAIL.n99 3.50912
R2704 VTAIL.n407 VTAIL.n405 3.50912
R2705 VTAIL.n352 VTAIL.n351 3.49141
R2706 VTAIL.n375 VTAIL.n322 3.49141
R2707 VTAIL.n398 VTAIL.n310 3.49141
R2708 VTAIL.n46 VTAIL.n45 3.49141
R2709 VTAIL.n69 VTAIL.n16 3.49141
R2710 VTAIL.n92 VTAIL.n4 3.49141
R2711 VTAIL.n300 VTAIL.n212 3.49141
R2712 VTAIL.n279 VTAIL.n226 3.49141
R2713 VTAIL.n256 VTAIL.n255 3.49141
R2714 VTAIL.n198 VTAIL.n110 3.49141
R2715 VTAIL.n177 VTAIL.n124 3.49141
R2716 VTAIL.n154 VTAIL.n153 3.49141
R2717 VTAIL.n348 VTAIL.n334 2.71565
R2718 VTAIL.n376 VTAIL.n320 2.71565
R2719 VTAIL.n397 VTAIL.n312 2.71565
R2720 VTAIL.n42 VTAIL.n28 2.71565
R2721 VTAIL.n70 VTAIL.n14 2.71565
R2722 VTAIL.n91 VTAIL.n6 2.71565
R2723 VTAIL.n299 VTAIL.n214 2.71565
R2724 VTAIL.n280 VTAIL.n224 2.71565
R2725 VTAIL.n252 VTAIL.n238 2.71565
R2726 VTAIL.n197 VTAIL.n112 2.71565
R2727 VTAIL.n178 VTAIL.n122 2.71565
R2728 VTAIL.n150 VTAIL.n136 2.71565
R2729 VTAIL VTAIL.n1 2.69016
R2730 VTAIL.n207 VTAIL.n205 2.22464
R2731 VTAIL.n99 VTAIL.n1 2.22464
R2732 VTAIL.n347 VTAIL.n336 1.93989
R2733 VTAIL.n381 VTAIL.n379 1.93989
R2734 VTAIL.n394 VTAIL.n393 1.93989
R2735 VTAIL.n41 VTAIL.n30 1.93989
R2736 VTAIL.n75 VTAIL.n73 1.93989
R2737 VTAIL.n88 VTAIL.n87 1.93989
R2738 VTAIL.n296 VTAIL.n295 1.93989
R2739 VTAIL.n284 VTAIL.n283 1.93989
R2740 VTAIL.n251 VTAIL.n240 1.93989
R2741 VTAIL.n194 VTAIL.n193 1.93989
R2742 VTAIL.n182 VTAIL.n181 1.93989
R2743 VTAIL.n149 VTAIL.n138 1.93989
R2744 VTAIL.n406 VTAIL.t7 1.86218
R2745 VTAIL.n406 VTAIL.t6 1.86218
R2746 VTAIL.n0 VTAIL.t8 1.86218
R2747 VTAIL.n0 VTAIL.t3 1.86218
R2748 VTAIL.n100 VTAIL.t14 1.86218
R2749 VTAIL.n100 VTAIL.t19 1.86218
R2750 VTAIL.n102 VTAIL.t10 1.86218
R2751 VTAIL.n102 VTAIL.t17 1.86218
R2752 VTAIL.n208 VTAIL.t13 1.86218
R2753 VTAIL.n208 VTAIL.t15 1.86218
R2754 VTAIL.n206 VTAIL.t12 1.86218
R2755 VTAIL.n206 VTAIL.t11 1.86218
R2756 VTAIL.n106 VTAIL.t5 1.86218
R2757 VTAIL.n106 VTAIL.t9 1.86218
R2758 VTAIL.n104 VTAIL.t2 1.86218
R2759 VTAIL.n104 VTAIL.t1 1.86218
R2760 VTAIL.n344 VTAIL.n343 1.16414
R2761 VTAIL.n380 VTAIL.n318 1.16414
R2762 VTAIL.n390 VTAIL.n314 1.16414
R2763 VTAIL.n38 VTAIL.n37 1.16414
R2764 VTAIL.n74 VTAIL.n12 1.16414
R2765 VTAIL.n84 VTAIL.n8 1.16414
R2766 VTAIL.n292 VTAIL.n216 1.16414
R2767 VTAIL.n287 VTAIL.n221 1.16414
R2768 VTAIL.n248 VTAIL.n247 1.16414
R2769 VTAIL.n190 VTAIL.n114 1.16414
R2770 VTAIL.n185 VTAIL.n119 1.16414
R2771 VTAIL.n146 VTAIL.n145 1.16414
R2772 VTAIL VTAIL.n407 0.819465
R2773 VTAIL.n340 VTAIL.n338 0.388379
R2774 VTAIL.n386 VTAIL.n385 0.388379
R2775 VTAIL.n389 VTAIL.n316 0.388379
R2776 VTAIL.n34 VTAIL.n32 0.388379
R2777 VTAIL.n80 VTAIL.n79 0.388379
R2778 VTAIL.n83 VTAIL.n10 0.388379
R2779 VTAIL.n291 VTAIL.n218 0.388379
R2780 VTAIL.n288 VTAIL.n220 0.388379
R2781 VTAIL.n244 VTAIL.n242 0.388379
R2782 VTAIL.n189 VTAIL.n116 0.388379
R2783 VTAIL.n186 VTAIL.n118 0.388379
R2784 VTAIL.n142 VTAIL.n140 0.388379
R2785 VTAIL.n345 VTAIL.n337 0.155672
R2786 VTAIL.n346 VTAIL.n345 0.155672
R2787 VTAIL.n346 VTAIL.n333 0.155672
R2788 VTAIL.n353 VTAIL.n333 0.155672
R2789 VTAIL.n354 VTAIL.n353 0.155672
R2790 VTAIL.n354 VTAIL.n329 0.155672
R2791 VTAIL.n361 VTAIL.n329 0.155672
R2792 VTAIL.n362 VTAIL.n361 0.155672
R2793 VTAIL.n362 VTAIL.n325 0.155672
R2794 VTAIL.n369 VTAIL.n325 0.155672
R2795 VTAIL.n370 VTAIL.n369 0.155672
R2796 VTAIL.n370 VTAIL.n321 0.155672
R2797 VTAIL.n377 VTAIL.n321 0.155672
R2798 VTAIL.n378 VTAIL.n377 0.155672
R2799 VTAIL.n378 VTAIL.n317 0.155672
R2800 VTAIL.n387 VTAIL.n317 0.155672
R2801 VTAIL.n388 VTAIL.n387 0.155672
R2802 VTAIL.n388 VTAIL.n313 0.155672
R2803 VTAIL.n395 VTAIL.n313 0.155672
R2804 VTAIL.n396 VTAIL.n395 0.155672
R2805 VTAIL.n396 VTAIL.n309 0.155672
R2806 VTAIL.n403 VTAIL.n309 0.155672
R2807 VTAIL.n39 VTAIL.n31 0.155672
R2808 VTAIL.n40 VTAIL.n39 0.155672
R2809 VTAIL.n40 VTAIL.n27 0.155672
R2810 VTAIL.n47 VTAIL.n27 0.155672
R2811 VTAIL.n48 VTAIL.n47 0.155672
R2812 VTAIL.n48 VTAIL.n23 0.155672
R2813 VTAIL.n55 VTAIL.n23 0.155672
R2814 VTAIL.n56 VTAIL.n55 0.155672
R2815 VTAIL.n56 VTAIL.n19 0.155672
R2816 VTAIL.n63 VTAIL.n19 0.155672
R2817 VTAIL.n64 VTAIL.n63 0.155672
R2818 VTAIL.n64 VTAIL.n15 0.155672
R2819 VTAIL.n71 VTAIL.n15 0.155672
R2820 VTAIL.n72 VTAIL.n71 0.155672
R2821 VTAIL.n72 VTAIL.n11 0.155672
R2822 VTAIL.n81 VTAIL.n11 0.155672
R2823 VTAIL.n82 VTAIL.n81 0.155672
R2824 VTAIL.n82 VTAIL.n7 0.155672
R2825 VTAIL.n89 VTAIL.n7 0.155672
R2826 VTAIL.n90 VTAIL.n89 0.155672
R2827 VTAIL.n90 VTAIL.n3 0.155672
R2828 VTAIL.n97 VTAIL.n3 0.155672
R2829 VTAIL.n305 VTAIL.n211 0.155672
R2830 VTAIL.n298 VTAIL.n211 0.155672
R2831 VTAIL.n298 VTAIL.n297 0.155672
R2832 VTAIL.n297 VTAIL.n215 0.155672
R2833 VTAIL.n290 VTAIL.n215 0.155672
R2834 VTAIL.n290 VTAIL.n289 0.155672
R2835 VTAIL.n289 VTAIL.n219 0.155672
R2836 VTAIL.n282 VTAIL.n219 0.155672
R2837 VTAIL.n282 VTAIL.n281 0.155672
R2838 VTAIL.n281 VTAIL.n225 0.155672
R2839 VTAIL.n274 VTAIL.n225 0.155672
R2840 VTAIL.n274 VTAIL.n273 0.155672
R2841 VTAIL.n273 VTAIL.n229 0.155672
R2842 VTAIL.n266 VTAIL.n229 0.155672
R2843 VTAIL.n266 VTAIL.n265 0.155672
R2844 VTAIL.n265 VTAIL.n233 0.155672
R2845 VTAIL.n258 VTAIL.n233 0.155672
R2846 VTAIL.n258 VTAIL.n257 0.155672
R2847 VTAIL.n257 VTAIL.n237 0.155672
R2848 VTAIL.n250 VTAIL.n237 0.155672
R2849 VTAIL.n250 VTAIL.n249 0.155672
R2850 VTAIL.n249 VTAIL.n241 0.155672
R2851 VTAIL.n203 VTAIL.n109 0.155672
R2852 VTAIL.n196 VTAIL.n109 0.155672
R2853 VTAIL.n196 VTAIL.n195 0.155672
R2854 VTAIL.n195 VTAIL.n113 0.155672
R2855 VTAIL.n188 VTAIL.n113 0.155672
R2856 VTAIL.n188 VTAIL.n187 0.155672
R2857 VTAIL.n187 VTAIL.n117 0.155672
R2858 VTAIL.n180 VTAIL.n117 0.155672
R2859 VTAIL.n180 VTAIL.n179 0.155672
R2860 VTAIL.n179 VTAIL.n123 0.155672
R2861 VTAIL.n172 VTAIL.n123 0.155672
R2862 VTAIL.n172 VTAIL.n171 0.155672
R2863 VTAIL.n171 VTAIL.n127 0.155672
R2864 VTAIL.n164 VTAIL.n127 0.155672
R2865 VTAIL.n164 VTAIL.n163 0.155672
R2866 VTAIL.n163 VTAIL.n131 0.155672
R2867 VTAIL.n156 VTAIL.n131 0.155672
R2868 VTAIL.n156 VTAIL.n155 0.155672
R2869 VTAIL.n155 VTAIL.n135 0.155672
R2870 VTAIL.n148 VTAIL.n135 0.155672
R2871 VTAIL.n148 VTAIL.n147 0.155672
R2872 VTAIL.n147 VTAIL.n139 0.155672
R2873 VN.n108 VN.n107 161.3
R2874 VN.n106 VN.n56 161.3
R2875 VN.n105 VN.n104 161.3
R2876 VN.n103 VN.n57 161.3
R2877 VN.n102 VN.n101 161.3
R2878 VN.n100 VN.n58 161.3
R2879 VN.n99 VN.n98 161.3
R2880 VN.n97 VN.n59 161.3
R2881 VN.n96 VN.n95 161.3
R2882 VN.n94 VN.n60 161.3
R2883 VN.n93 VN.n92 161.3
R2884 VN.n91 VN.n62 161.3
R2885 VN.n90 VN.n89 161.3
R2886 VN.n88 VN.n63 161.3
R2887 VN.n87 VN.n86 161.3
R2888 VN.n85 VN.n64 161.3
R2889 VN.n84 VN.n83 161.3
R2890 VN.n82 VN.n65 161.3
R2891 VN.n81 VN.n80 161.3
R2892 VN.n79 VN.n66 161.3
R2893 VN.n78 VN.n77 161.3
R2894 VN.n76 VN.n67 161.3
R2895 VN.n75 VN.n74 161.3
R2896 VN.n73 VN.n68 161.3
R2897 VN.n72 VN.n71 161.3
R2898 VN.n53 VN.n52 161.3
R2899 VN.n51 VN.n1 161.3
R2900 VN.n50 VN.n49 161.3
R2901 VN.n48 VN.n2 161.3
R2902 VN.n47 VN.n46 161.3
R2903 VN.n45 VN.n3 161.3
R2904 VN.n44 VN.n43 161.3
R2905 VN.n42 VN.n4 161.3
R2906 VN.n41 VN.n40 161.3
R2907 VN.n38 VN.n5 161.3
R2908 VN.n37 VN.n36 161.3
R2909 VN.n35 VN.n6 161.3
R2910 VN.n34 VN.n33 161.3
R2911 VN.n32 VN.n7 161.3
R2912 VN.n31 VN.n30 161.3
R2913 VN.n29 VN.n8 161.3
R2914 VN.n28 VN.n27 161.3
R2915 VN.n26 VN.n9 161.3
R2916 VN.n25 VN.n24 161.3
R2917 VN.n23 VN.n10 161.3
R2918 VN.n22 VN.n21 161.3
R2919 VN.n20 VN.n11 161.3
R2920 VN.n19 VN.n18 161.3
R2921 VN.n17 VN.n12 161.3
R2922 VN.n16 VN.n15 161.3
R2923 VN.n69 VN.t2 145.398
R2924 VN.n13 VN.t8 145.398
R2925 VN.n27 VN.t1 112.51
R2926 VN.n14 VN.t5 112.51
R2927 VN.n39 VN.t9 112.51
R2928 VN.n0 VN.t4 112.51
R2929 VN.n83 VN.t7 112.51
R2930 VN.n70 VN.t6 112.51
R2931 VN.n61 VN.t3 112.51
R2932 VN.n55 VN.t0 112.51
R2933 VN.n54 VN.n0 83.3598
R2934 VN.n109 VN.n55 83.3598
R2935 VN.n14 VN.n13 71.5921
R2936 VN.n70 VN.n69 71.5921
R2937 VN VN.n109 63.714
R2938 VN.n46 VN.n2 50.7491
R2939 VN.n101 VN.n57 50.7491
R2940 VN.n21 VN.n20 43.9677
R2941 VN.n33 VN.n6 43.9677
R2942 VN.n77 VN.n76 43.9677
R2943 VN.n89 VN.n62 43.9677
R2944 VN.n21 VN.n10 37.1863
R2945 VN.n33 VN.n32 37.1863
R2946 VN.n77 VN.n66 37.1863
R2947 VN.n89 VN.n88 37.1863
R2948 VN.n46 VN.n45 30.405
R2949 VN.n101 VN.n100 30.405
R2950 VN.n15 VN.n12 24.5923
R2951 VN.n19 VN.n12 24.5923
R2952 VN.n20 VN.n19 24.5923
R2953 VN.n25 VN.n10 24.5923
R2954 VN.n26 VN.n25 24.5923
R2955 VN.n27 VN.n26 24.5923
R2956 VN.n27 VN.n8 24.5923
R2957 VN.n31 VN.n8 24.5923
R2958 VN.n32 VN.n31 24.5923
R2959 VN.n37 VN.n6 24.5923
R2960 VN.n38 VN.n37 24.5923
R2961 VN.n40 VN.n38 24.5923
R2962 VN.n44 VN.n4 24.5923
R2963 VN.n45 VN.n44 24.5923
R2964 VN.n50 VN.n2 24.5923
R2965 VN.n51 VN.n50 24.5923
R2966 VN.n52 VN.n51 24.5923
R2967 VN.n76 VN.n75 24.5923
R2968 VN.n75 VN.n68 24.5923
R2969 VN.n71 VN.n68 24.5923
R2970 VN.n88 VN.n87 24.5923
R2971 VN.n87 VN.n64 24.5923
R2972 VN.n83 VN.n64 24.5923
R2973 VN.n83 VN.n82 24.5923
R2974 VN.n82 VN.n81 24.5923
R2975 VN.n81 VN.n66 24.5923
R2976 VN.n100 VN.n99 24.5923
R2977 VN.n99 VN.n59 24.5923
R2978 VN.n95 VN.n94 24.5923
R2979 VN.n94 VN.n93 24.5923
R2980 VN.n93 VN.n62 24.5923
R2981 VN.n107 VN.n106 24.5923
R2982 VN.n106 VN.n105 24.5923
R2983 VN.n105 VN.n57 24.5923
R2984 VN.n39 VN.n4 21.1495
R2985 VN.n61 VN.n59 21.1495
R2986 VN.n52 VN.n0 6.88621
R2987 VN.n107 VN.n55 6.88621
R2988 VN.n15 VN.n14 3.44336
R2989 VN.n40 VN.n39 3.44336
R2990 VN.n71 VN.n70 3.44336
R2991 VN.n95 VN.n61 3.44336
R2992 VN.n72 VN.n69 3.23944
R2993 VN.n16 VN.n13 3.23944
R2994 VN.n109 VN.n108 0.354861
R2995 VN.n54 VN.n53 0.354861
R2996 VN VN.n54 0.267071
R2997 VN.n108 VN.n56 0.189894
R2998 VN.n104 VN.n56 0.189894
R2999 VN.n104 VN.n103 0.189894
R3000 VN.n103 VN.n102 0.189894
R3001 VN.n102 VN.n58 0.189894
R3002 VN.n98 VN.n58 0.189894
R3003 VN.n98 VN.n97 0.189894
R3004 VN.n97 VN.n96 0.189894
R3005 VN.n96 VN.n60 0.189894
R3006 VN.n92 VN.n60 0.189894
R3007 VN.n92 VN.n91 0.189894
R3008 VN.n91 VN.n90 0.189894
R3009 VN.n90 VN.n63 0.189894
R3010 VN.n86 VN.n63 0.189894
R3011 VN.n86 VN.n85 0.189894
R3012 VN.n85 VN.n84 0.189894
R3013 VN.n84 VN.n65 0.189894
R3014 VN.n80 VN.n65 0.189894
R3015 VN.n80 VN.n79 0.189894
R3016 VN.n79 VN.n78 0.189894
R3017 VN.n78 VN.n67 0.189894
R3018 VN.n74 VN.n67 0.189894
R3019 VN.n74 VN.n73 0.189894
R3020 VN.n73 VN.n72 0.189894
R3021 VN.n17 VN.n16 0.189894
R3022 VN.n18 VN.n17 0.189894
R3023 VN.n18 VN.n11 0.189894
R3024 VN.n22 VN.n11 0.189894
R3025 VN.n23 VN.n22 0.189894
R3026 VN.n24 VN.n23 0.189894
R3027 VN.n24 VN.n9 0.189894
R3028 VN.n28 VN.n9 0.189894
R3029 VN.n29 VN.n28 0.189894
R3030 VN.n30 VN.n29 0.189894
R3031 VN.n30 VN.n7 0.189894
R3032 VN.n34 VN.n7 0.189894
R3033 VN.n35 VN.n34 0.189894
R3034 VN.n36 VN.n35 0.189894
R3035 VN.n36 VN.n5 0.189894
R3036 VN.n41 VN.n5 0.189894
R3037 VN.n42 VN.n41 0.189894
R3038 VN.n43 VN.n42 0.189894
R3039 VN.n43 VN.n3 0.189894
R3040 VN.n47 VN.n3 0.189894
R3041 VN.n48 VN.n47 0.189894
R3042 VN.n49 VN.n48 0.189894
R3043 VN.n49 VN.n1 0.189894
R3044 VN.n53 VN.n1 0.189894
R3045 VDD2.n193 VDD2.n101 756.745
R3046 VDD2.n92 VDD2.n0 756.745
R3047 VDD2.n194 VDD2.n193 585
R3048 VDD2.n192 VDD2.n191 585
R3049 VDD2.n105 VDD2.n104 585
R3050 VDD2.n186 VDD2.n185 585
R3051 VDD2.n184 VDD2.n183 585
R3052 VDD2.n109 VDD2.n108 585
R3053 VDD2.n113 VDD2.n111 585
R3054 VDD2.n178 VDD2.n177 585
R3055 VDD2.n176 VDD2.n175 585
R3056 VDD2.n115 VDD2.n114 585
R3057 VDD2.n170 VDD2.n169 585
R3058 VDD2.n168 VDD2.n167 585
R3059 VDD2.n119 VDD2.n118 585
R3060 VDD2.n162 VDD2.n161 585
R3061 VDD2.n160 VDD2.n159 585
R3062 VDD2.n123 VDD2.n122 585
R3063 VDD2.n154 VDD2.n153 585
R3064 VDD2.n152 VDD2.n151 585
R3065 VDD2.n127 VDD2.n126 585
R3066 VDD2.n146 VDD2.n145 585
R3067 VDD2.n144 VDD2.n143 585
R3068 VDD2.n131 VDD2.n130 585
R3069 VDD2.n138 VDD2.n137 585
R3070 VDD2.n136 VDD2.n135 585
R3071 VDD2.n33 VDD2.n32 585
R3072 VDD2.n35 VDD2.n34 585
R3073 VDD2.n28 VDD2.n27 585
R3074 VDD2.n41 VDD2.n40 585
R3075 VDD2.n43 VDD2.n42 585
R3076 VDD2.n24 VDD2.n23 585
R3077 VDD2.n49 VDD2.n48 585
R3078 VDD2.n51 VDD2.n50 585
R3079 VDD2.n20 VDD2.n19 585
R3080 VDD2.n57 VDD2.n56 585
R3081 VDD2.n59 VDD2.n58 585
R3082 VDD2.n16 VDD2.n15 585
R3083 VDD2.n65 VDD2.n64 585
R3084 VDD2.n67 VDD2.n66 585
R3085 VDD2.n12 VDD2.n11 585
R3086 VDD2.n74 VDD2.n73 585
R3087 VDD2.n75 VDD2.n10 585
R3088 VDD2.n77 VDD2.n76 585
R3089 VDD2.n8 VDD2.n7 585
R3090 VDD2.n83 VDD2.n82 585
R3091 VDD2.n85 VDD2.n84 585
R3092 VDD2.n4 VDD2.n3 585
R3093 VDD2.n91 VDD2.n90 585
R3094 VDD2.n93 VDD2.n92 585
R3095 VDD2.n134 VDD2.t9 327.466
R3096 VDD2.n31 VDD2.t1 327.466
R3097 VDD2.n193 VDD2.n192 171.744
R3098 VDD2.n192 VDD2.n104 171.744
R3099 VDD2.n185 VDD2.n104 171.744
R3100 VDD2.n185 VDD2.n184 171.744
R3101 VDD2.n184 VDD2.n108 171.744
R3102 VDD2.n113 VDD2.n108 171.744
R3103 VDD2.n177 VDD2.n113 171.744
R3104 VDD2.n177 VDD2.n176 171.744
R3105 VDD2.n176 VDD2.n114 171.744
R3106 VDD2.n169 VDD2.n114 171.744
R3107 VDD2.n169 VDD2.n168 171.744
R3108 VDD2.n168 VDD2.n118 171.744
R3109 VDD2.n161 VDD2.n118 171.744
R3110 VDD2.n161 VDD2.n160 171.744
R3111 VDD2.n160 VDD2.n122 171.744
R3112 VDD2.n153 VDD2.n122 171.744
R3113 VDD2.n153 VDD2.n152 171.744
R3114 VDD2.n152 VDD2.n126 171.744
R3115 VDD2.n145 VDD2.n126 171.744
R3116 VDD2.n145 VDD2.n144 171.744
R3117 VDD2.n144 VDD2.n130 171.744
R3118 VDD2.n137 VDD2.n130 171.744
R3119 VDD2.n137 VDD2.n136 171.744
R3120 VDD2.n34 VDD2.n33 171.744
R3121 VDD2.n34 VDD2.n27 171.744
R3122 VDD2.n41 VDD2.n27 171.744
R3123 VDD2.n42 VDD2.n41 171.744
R3124 VDD2.n42 VDD2.n23 171.744
R3125 VDD2.n49 VDD2.n23 171.744
R3126 VDD2.n50 VDD2.n49 171.744
R3127 VDD2.n50 VDD2.n19 171.744
R3128 VDD2.n57 VDD2.n19 171.744
R3129 VDD2.n58 VDD2.n57 171.744
R3130 VDD2.n58 VDD2.n15 171.744
R3131 VDD2.n65 VDD2.n15 171.744
R3132 VDD2.n66 VDD2.n65 171.744
R3133 VDD2.n66 VDD2.n11 171.744
R3134 VDD2.n74 VDD2.n11 171.744
R3135 VDD2.n75 VDD2.n74 171.744
R3136 VDD2.n76 VDD2.n75 171.744
R3137 VDD2.n76 VDD2.n7 171.744
R3138 VDD2.n83 VDD2.n7 171.744
R3139 VDD2.n84 VDD2.n83 171.744
R3140 VDD2.n84 VDD2.n3 171.744
R3141 VDD2.n91 VDD2.n3 171.744
R3142 VDD2.n92 VDD2.n91 171.744
R3143 VDD2.n136 VDD2.t9 85.8723
R3144 VDD2.n33 VDD2.t1 85.8723
R3145 VDD2.n100 VDD2.n99 70.4345
R3146 VDD2 VDD2.n201 70.4317
R3147 VDD2.n200 VDD2.n199 67.8586
R3148 VDD2.n98 VDD2.n97 67.8584
R3149 VDD2.n198 VDD2.n100 55.433
R3150 VDD2.n98 VDD2.n96 51.2091
R3151 VDD2.n198 VDD2.n197 47.7005
R3152 VDD2.n135 VDD2.n134 16.3895
R3153 VDD2.n32 VDD2.n31 16.3895
R3154 VDD2.n111 VDD2.n109 13.1884
R3155 VDD2.n77 VDD2.n8 13.1884
R3156 VDD2.n183 VDD2.n182 12.8005
R3157 VDD2.n179 VDD2.n178 12.8005
R3158 VDD2.n138 VDD2.n133 12.8005
R3159 VDD2.n35 VDD2.n30 12.8005
R3160 VDD2.n78 VDD2.n10 12.8005
R3161 VDD2.n82 VDD2.n81 12.8005
R3162 VDD2.n186 VDD2.n107 12.0247
R3163 VDD2.n175 VDD2.n112 12.0247
R3164 VDD2.n139 VDD2.n131 12.0247
R3165 VDD2.n36 VDD2.n28 12.0247
R3166 VDD2.n73 VDD2.n72 12.0247
R3167 VDD2.n85 VDD2.n6 12.0247
R3168 VDD2.n187 VDD2.n105 11.249
R3169 VDD2.n174 VDD2.n115 11.249
R3170 VDD2.n143 VDD2.n142 11.249
R3171 VDD2.n40 VDD2.n39 11.249
R3172 VDD2.n71 VDD2.n12 11.249
R3173 VDD2.n86 VDD2.n4 11.249
R3174 VDD2.n191 VDD2.n190 10.4732
R3175 VDD2.n171 VDD2.n170 10.4732
R3176 VDD2.n146 VDD2.n129 10.4732
R3177 VDD2.n43 VDD2.n26 10.4732
R3178 VDD2.n68 VDD2.n67 10.4732
R3179 VDD2.n90 VDD2.n89 10.4732
R3180 VDD2.n194 VDD2.n103 9.69747
R3181 VDD2.n167 VDD2.n117 9.69747
R3182 VDD2.n147 VDD2.n127 9.69747
R3183 VDD2.n44 VDD2.n24 9.69747
R3184 VDD2.n64 VDD2.n14 9.69747
R3185 VDD2.n93 VDD2.n2 9.69747
R3186 VDD2.n197 VDD2.n196 9.45567
R3187 VDD2.n96 VDD2.n95 9.45567
R3188 VDD2.n121 VDD2.n120 9.3005
R3189 VDD2.n164 VDD2.n163 9.3005
R3190 VDD2.n166 VDD2.n165 9.3005
R3191 VDD2.n117 VDD2.n116 9.3005
R3192 VDD2.n172 VDD2.n171 9.3005
R3193 VDD2.n174 VDD2.n173 9.3005
R3194 VDD2.n112 VDD2.n110 9.3005
R3195 VDD2.n180 VDD2.n179 9.3005
R3196 VDD2.n196 VDD2.n195 9.3005
R3197 VDD2.n103 VDD2.n102 9.3005
R3198 VDD2.n190 VDD2.n189 9.3005
R3199 VDD2.n188 VDD2.n187 9.3005
R3200 VDD2.n107 VDD2.n106 9.3005
R3201 VDD2.n182 VDD2.n181 9.3005
R3202 VDD2.n158 VDD2.n157 9.3005
R3203 VDD2.n156 VDD2.n155 9.3005
R3204 VDD2.n125 VDD2.n124 9.3005
R3205 VDD2.n150 VDD2.n149 9.3005
R3206 VDD2.n148 VDD2.n147 9.3005
R3207 VDD2.n129 VDD2.n128 9.3005
R3208 VDD2.n142 VDD2.n141 9.3005
R3209 VDD2.n140 VDD2.n139 9.3005
R3210 VDD2.n133 VDD2.n132 9.3005
R3211 VDD2.n95 VDD2.n94 9.3005
R3212 VDD2.n2 VDD2.n1 9.3005
R3213 VDD2.n89 VDD2.n88 9.3005
R3214 VDD2.n87 VDD2.n86 9.3005
R3215 VDD2.n6 VDD2.n5 9.3005
R3216 VDD2.n81 VDD2.n80 9.3005
R3217 VDD2.n53 VDD2.n52 9.3005
R3218 VDD2.n22 VDD2.n21 9.3005
R3219 VDD2.n47 VDD2.n46 9.3005
R3220 VDD2.n45 VDD2.n44 9.3005
R3221 VDD2.n26 VDD2.n25 9.3005
R3222 VDD2.n39 VDD2.n38 9.3005
R3223 VDD2.n37 VDD2.n36 9.3005
R3224 VDD2.n30 VDD2.n29 9.3005
R3225 VDD2.n55 VDD2.n54 9.3005
R3226 VDD2.n18 VDD2.n17 9.3005
R3227 VDD2.n61 VDD2.n60 9.3005
R3228 VDD2.n63 VDD2.n62 9.3005
R3229 VDD2.n14 VDD2.n13 9.3005
R3230 VDD2.n69 VDD2.n68 9.3005
R3231 VDD2.n71 VDD2.n70 9.3005
R3232 VDD2.n72 VDD2.n9 9.3005
R3233 VDD2.n79 VDD2.n78 9.3005
R3234 VDD2.n195 VDD2.n101 8.92171
R3235 VDD2.n166 VDD2.n119 8.92171
R3236 VDD2.n151 VDD2.n150 8.92171
R3237 VDD2.n48 VDD2.n47 8.92171
R3238 VDD2.n63 VDD2.n16 8.92171
R3239 VDD2.n94 VDD2.n0 8.92171
R3240 VDD2.n163 VDD2.n162 8.14595
R3241 VDD2.n154 VDD2.n125 8.14595
R3242 VDD2.n51 VDD2.n22 8.14595
R3243 VDD2.n60 VDD2.n59 8.14595
R3244 VDD2.n159 VDD2.n121 7.3702
R3245 VDD2.n155 VDD2.n123 7.3702
R3246 VDD2.n52 VDD2.n20 7.3702
R3247 VDD2.n56 VDD2.n18 7.3702
R3248 VDD2.n159 VDD2.n158 6.59444
R3249 VDD2.n158 VDD2.n123 6.59444
R3250 VDD2.n55 VDD2.n20 6.59444
R3251 VDD2.n56 VDD2.n55 6.59444
R3252 VDD2.n162 VDD2.n121 5.81868
R3253 VDD2.n155 VDD2.n154 5.81868
R3254 VDD2.n52 VDD2.n51 5.81868
R3255 VDD2.n59 VDD2.n18 5.81868
R3256 VDD2.n197 VDD2.n101 5.04292
R3257 VDD2.n163 VDD2.n119 5.04292
R3258 VDD2.n151 VDD2.n125 5.04292
R3259 VDD2.n48 VDD2.n22 5.04292
R3260 VDD2.n60 VDD2.n16 5.04292
R3261 VDD2.n96 VDD2.n0 5.04292
R3262 VDD2.n195 VDD2.n194 4.26717
R3263 VDD2.n167 VDD2.n166 4.26717
R3264 VDD2.n150 VDD2.n127 4.26717
R3265 VDD2.n47 VDD2.n24 4.26717
R3266 VDD2.n64 VDD2.n63 4.26717
R3267 VDD2.n94 VDD2.n93 4.26717
R3268 VDD2.n134 VDD2.n132 3.70982
R3269 VDD2.n31 VDD2.n29 3.70982
R3270 VDD2.n200 VDD2.n198 3.50912
R3271 VDD2.n191 VDD2.n103 3.49141
R3272 VDD2.n170 VDD2.n117 3.49141
R3273 VDD2.n147 VDD2.n146 3.49141
R3274 VDD2.n44 VDD2.n43 3.49141
R3275 VDD2.n67 VDD2.n14 3.49141
R3276 VDD2.n90 VDD2.n2 3.49141
R3277 VDD2.n190 VDD2.n105 2.71565
R3278 VDD2.n171 VDD2.n115 2.71565
R3279 VDD2.n143 VDD2.n129 2.71565
R3280 VDD2.n40 VDD2.n26 2.71565
R3281 VDD2.n68 VDD2.n12 2.71565
R3282 VDD2.n89 VDD2.n4 2.71565
R3283 VDD2.n187 VDD2.n186 1.93989
R3284 VDD2.n175 VDD2.n174 1.93989
R3285 VDD2.n142 VDD2.n131 1.93989
R3286 VDD2.n39 VDD2.n28 1.93989
R3287 VDD2.n73 VDD2.n71 1.93989
R3288 VDD2.n86 VDD2.n85 1.93989
R3289 VDD2.n201 VDD2.t3 1.86218
R3290 VDD2.n201 VDD2.t7 1.86218
R3291 VDD2.n199 VDD2.t6 1.86218
R3292 VDD2.n199 VDD2.t2 1.86218
R3293 VDD2.n99 VDD2.t0 1.86218
R3294 VDD2.n99 VDD2.t5 1.86218
R3295 VDD2.n97 VDD2.t4 1.86218
R3296 VDD2.n97 VDD2.t8 1.86218
R3297 VDD2.n183 VDD2.n107 1.16414
R3298 VDD2.n178 VDD2.n112 1.16414
R3299 VDD2.n139 VDD2.n138 1.16414
R3300 VDD2.n36 VDD2.n35 1.16414
R3301 VDD2.n72 VDD2.n10 1.16414
R3302 VDD2.n82 VDD2.n6 1.16414
R3303 VDD2 VDD2.n200 0.935845
R3304 VDD2.n100 VDD2.n98 0.822309
R3305 VDD2.n182 VDD2.n109 0.388379
R3306 VDD2.n179 VDD2.n111 0.388379
R3307 VDD2.n135 VDD2.n133 0.388379
R3308 VDD2.n32 VDD2.n30 0.388379
R3309 VDD2.n78 VDD2.n77 0.388379
R3310 VDD2.n81 VDD2.n8 0.388379
R3311 VDD2.n196 VDD2.n102 0.155672
R3312 VDD2.n189 VDD2.n102 0.155672
R3313 VDD2.n189 VDD2.n188 0.155672
R3314 VDD2.n188 VDD2.n106 0.155672
R3315 VDD2.n181 VDD2.n106 0.155672
R3316 VDD2.n181 VDD2.n180 0.155672
R3317 VDD2.n180 VDD2.n110 0.155672
R3318 VDD2.n173 VDD2.n110 0.155672
R3319 VDD2.n173 VDD2.n172 0.155672
R3320 VDD2.n172 VDD2.n116 0.155672
R3321 VDD2.n165 VDD2.n116 0.155672
R3322 VDD2.n165 VDD2.n164 0.155672
R3323 VDD2.n164 VDD2.n120 0.155672
R3324 VDD2.n157 VDD2.n120 0.155672
R3325 VDD2.n157 VDD2.n156 0.155672
R3326 VDD2.n156 VDD2.n124 0.155672
R3327 VDD2.n149 VDD2.n124 0.155672
R3328 VDD2.n149 VDD2.n148 0.155672
R3329 VDD2.n148 VDD2.n128 0.155672
R3330 VDD2.n141 VDD2.n128 0.155672
R3331 VDD2.n141 VDD2.n140 0.155672
R3332 VDD2.n140 VDD2.n132 0.155672
R3333 VDD2.n37 VDD2.n29 0.155672
R3334 VDD2.n38 VDD2.n37 0.155672
R3335 VDD2.n38 VDD2.n25 0.155672
R3336 VDD2.n45 VDD2.n25 0.155672
R3337 VDD2.n46 VDD2.n45 0.155672
R3338 VDD2.n46 VDD2.n21 0.155672
R3339 VDD2.n53 VDD2.n21 0.155672
R3340 VDD2.n54 VDD2.n53 0.155672
R3341 VDD2.n54 VDD2.n17 0.155672
R3342 VDD2.n61 VDD2.n17 0.155672
R3343 VDD2.n62 VDD2.n61 0.155672
R3344 VDD2.n62 VDD2.n13 0.155672
R3345 VDD2.n69 VDD2.n13 0.155672
R3346 VDD2.n70 VDD2.n69 0.155672
R3347 VDD2.n70 VDD2.n9 0.155672
R3348 VDD2.n79 VDD2.n9 0.155672
R3349 VDD2.n80 VDD2.n79 0.155672
R3350 VDD2.n80 VDD2.n5 0.155672
R3351 VDD2.n87 VDD2.n5 0.155672
R3352 VDD2.n88 VDD2.n87 0.155672
R3353 VDD2.n88 VDD2.n1 0.155672
R3354 VDD2.n95 VDD2.n1 0.155672
C0 VDD1 B 3.36372f
C1 VDD2 B 3.52603f
C2 VDD1 VP 16.835302f
C3 w_n5854_n4460# B 13.9941f
C4 VDD2 VP 0.728979f
C5 B VN 1.64221f
C6 w_n5854_n4460# VP 13.718901f
C7 VP VN 11.0807f
C8 B VTAIL 5.46229f
C9 VDD1 VDD2 2.91634f
C10 VP VTAIL 17.1508f
C11 w_n5854_n4460# VDD1 3.58823f
C12 VDD1 VN 0.156125f
C13 w_n5854_n4460# VDD2 3.79104f
C14 VDD2 VN 16.2665f
C15 VDD1 VTAIL 13.0963f
C16 w_n5854_n4460# VN 12.9532f
C17 VDD2 VTAIL 13.155f
C18 w_n5854_n4460# VTAIL 4.10318f
C19 VN VTAIL 17.136f
C20 B VP 2.93604f
C21 VDD2 VSUBS 2.68896f
C22 VDD1 VSUBS 2.567404f
C23 VTAIL VSUBS 1.757516f
C24 VN VSUBS 9.756379f
C25 VP VSUBS 5.886122f
C26 B VSUBS 7.239938f
C27 w_n5854_n4460# VSUBS 0.319418p
C28 VDD2.n0 VSUBS 0.03083f
C29 VDD2.n1 VSUBS 0.0293f
C30 VDD2.n2 VSUBS 0.015744f
C31 VDD2.n3 VSUBS 0.037214f
C32 VDD2.n4 VSUBS 0.016671f
C33 VDD2.n5 VSUBS 0.0293f
C34 VDD2.n6 VSUBS 0.015744f
C35 VDD2.n7 VSUBS 0.037214f
C36 VDD2.n8 VSUBS 0.016208f
C37 VDD2.n9 VSUBS 0.0293f
C38 VDD2.n10 VSUBS 0.016671f
C39 VDD2.n11 VSUBS 0.037214f
C40 VDD2.n12 VSUBS 0.016671f
C41 VDD2.n13 VSUBS 0.0293f
C42 VDD2.n14 VSUBS 0.015744f
C43 VDD2.n15 VSUBS 0.037214f
C44 VDD2.n16 VSUBS 0.016671f
C45 VDD2.n17 VSUBS 0.0293f
C46 VDD2.n18 VSUBS 0.015744f
C47 VDD2.n19 VSUBS 0.037214f
C48 VDD2.n20 VSUBS 0.016671f
C49 VDD2.n21 VSUBS 0.0293f
C50 VDD2.n22 VSUBS 0.015744f
C51 VDD2.n23 VSUBS 0.037214f
C52 VDD2.n24 VSUBS 0.016671f
C53 VDD2.n25 VSUBS 0.0293f
C54 VDD2.n26 VSUBS 0.015744f
C55 VDD2.n27 VSUBS 0.037214f
C56 VDD2.n28 VSUBS 0.016671f
C57 VDD2.n29 VSUBS 2.19808f
C58 VDD2.n30 VSUBS 0.015744f
C59 VDD2.t1 VSUBS 0.079848f
C60 VDD2.n31 VSUBS 0.227799f
C61 VDD2.n32 VSUBS 0.023674f
C62 VDD2.n33 VSUBS 0.027911f
C63 VDD2.n34 VSUBS 0.037214f
C64 VDD2.n35 VSUBS 0.016671f
C65 VDD2.n36 VSUBS 0.015744f
C66 VDD2.n37 VSUBS 0.0293f
C67 VDD2.n38 VSUBS 0.0293f
C68 VDD2.n39 VSUBS 0.015744f
C69 VDD2.n40 VSUBS 0.016671f
C70 VDD2.n41 VSUBS 0.037214f
C71 VDD2.n42 VSUBS 0.037214f
C72 VDD2.n43 VSUBS 0.016671f
C73 VDD2.n44 VSUBS 0.015744f
C74 VDD2.n45 VSUBS 0.0293f
C75 VDD2.n46 VSUBS 0.0293f
C76 VDD2.n47 VSUBS 0.015744f
C77 VDD2.n48 VSUBS 0.016671f
C78 VDD2.n49 VSUBS 0.037214f
C79 VDD2.n50 VSUBS 0.037214f
C80 VDD2.n51 VSUBS 0.016671f
C81 VDD2.n52 VSUBS 0.015744f
C82 VDD2.n53 VSUBS 0.0293f
C83 VDD2.n54 VSUBS 0.0293f
C84 VDD2.n55 VSUBS 0.015744f
C85 VDD2.n56 VSUBS 0.016671f
C86 VDD2.n57 VSUBS 0.037214f
C87 VDD2.n58 VSUBS 0.037214f
C88 VDD2.n59 VSUBS 0.016671f
C89 VDD2.n60 VSUBS 0.015744f
C90 VDD2.n61 VSUBS 0.0293f
C91 VDD2.n62 VSUBS 0.0293f
C92 VDD2.n63 VSUBS 0.015744f
C93 VDD2.n64 VSUBS 0.016671f
C94 VDD2.n65 VSUBS 0.037214f
C95 VDD2.n66 VSUBS 0.037214f
C96 VDD2.n67 VSUBS 0.016671f
C97 VDD2.n68 VSUBS 0.015744f
C98 VDD2.n69 VSUBS 0.0293f
C99 VDD2.n70 VSUBS 0.0293f
C100 VDD2.n71 VSUBS 0.015744f
C101 VDD2.n72 VSUBS 0.015744f
C102 VDD2.n73 VSUBS 0.016671f
C103 VDD2.n74 VSUBS 0.037214f
C104 VDD2.n75 VSUBS 0.037214f
C105 VDD2.n76 VSUBS 0.037214f
C106 VDD2.n77 VSUBS 0.016208f
C107 VDD2.n78 VSUBS 0.015744f
C108 VDD2.n79 VSUBS 0.0293f
C109 VDD2.n80 VSUBS 0.0293f
C110 VDD2.n81 VSUBS 0.015744f
C111 VDD2.n82 VSUBS 0.016671f
C112 VDD2.n83 VSUBS 0.037214f
C113 VDD2.n84 VSUBS 0.037214f
C114 VDD2.n85 VSUBS 0.016671f
C115 VDD2.n86 VSUBS 0.015744f
C116 VDD2.n87 VSUBS 0.0293f
C117 VDD2.n88 VSUBS 0.0293f
C118 VDD2.n89 VSUBS 0.015744f
C119 VDD2.n90 VSUBS 0.016671f
C120 VDD2.n91 VSUBS 0.037214f
C121 VDD2.n92 VSUBS 0.085444f
C122 VDD2.n93 VSUBS 0.016671f
C123 VDD2.n94 VSUBS 0.015744f
C124 VDD2.n95 VSUBS 0.065324f
C125 VDD2.n96 VSUBS 0.089406f
C126 VDD2.t4 VSUBS 0.404264f
C127 VDD2.t8 VSUBS 0.404264f
C128 VDD2.n97 VSUBS 3.33869f
C129 VDD2.n98 VSUBS 1.35199f
C130 VDD2.t0 VSUBS 0.404264f
C131 VDD2.t5 VSUBS 0.404264f
C132 VDD2.n99 VSUBS 3.38145f
C133 VDD2.n100 VSUBS 4.83418f
C134 VDD2.n101 VSUBS 0.03083f
C135 VDD2.n102 VSUBS 0.0293f
C136 VDD2.n103 VSUBS 0.015744f
C137 VDD2.n104 VSUBS 0.037214f
C138 VDD2.n105 VSUBS 0.016671f
C139 VDD2.n106 VSUBS 0.0293f
C140 VDD2.n107 VSUBS 0.015744f
C141 VDD2.n108 VSUBS 0.037214f
C142 VDD2.n109 VSUBS 0.016208f
C143 VDD2.n110 VSUBS 0.0293f
C144 VDD2.n111 VSUBS 0.016208f
C145 VDD2.n112 VSUBS 0.015744f
C146 VDD2.n113 VSUBS 0.037214f
C147 VDD2.n114 VSUBS 0.037214f
C148 VDD2.n115 VSUBS 0.016671f
C149 VDD2.n116 VSUBS 0.0293f
C150 VDD2.n117 VSUBS 0.015744f
C151 VDD2.n118 VSUBS 0.037214f
C152 VDD2.n119 VSUBS 0.016671f
C153 VDD2.n120 VSUBS 0.0293f
C154 VDD2.n121 VSUBS 0.015744f
C155 VDD2.n122 VSUBS 0.037214f
C156 VDD2.n123 VSUBS 0.016671f
C157 VDD2.n124 VSUBS 0.0293f
C158 VDD2.n125 VSUBS 0.015744f
C159 VDD2.n126 VSUBS 0.037214f
C160 VDD2.n127 VSUBS 0.016671f
C161 VDD2.n128 VSUBS 0.0293f
C162 VDD2.n129 VSUBS 0.015744f
C163 VDD2.n130 VSUBS 0.037214f
C164 VDD2.n131 VSUBS 0.016671f
C165 VDD2.n132 VSUBS 2.19808f
C166 VDD2.n133 VSUBS 0.015744f
C167 VDD2.t9 VSUBS 0.079848f
C168 VDD2.n134 VSUBS 0.227799f
C169 VDD2.n135 VSUBS 0.023674f
C170 VDD2.n136 VSUBS 0.027911f
C171 VDD2.n137 VSUBS 0.037214f
C172 VDD2.n138 VSUBS 0.016671f
C173 VDD2.n139 VSUBS 0.015744f
C174 VDD2.n140 VSUBS 0.0293f
C175 VDD2.n141 VSUBS 0.0293f
C176 VDD2.n142 VSUBS 0.015744f
C177 VDD2.n143 VSUBS 0.016671f
C178 VDD2.n144 VSUBS 0.037214f
C179 VDD2.n145 VSUBS 0.037214f
C180 VDD2.n146 VSUBS 0.016671f
C181 VDD2.n147 VSUBS 0.015744f
C182 VDD2.n148 VSUBS 0.0293f
C183 VDD2.n149 VSUBS 0.0293f
C184 VDD2.n150 VSUBS 0.015744f
C185 VDD2.n151 VSUBS 0.016671f
C186 VDD2.n152 VSUBS 0.037214f
C187 VDD2.n153 VSUBS 0.037214f
C188 VDD2.n154 VSUBS 0.016671f
C189 VDD2.n155 VSUBS 0.015744f
C190 VDD2.n156 VSUBS 0.0293f
C191 VDD2.n157 VSUBS 0.0293f
C192 VDD2.n158 VSUBS 0.015744f
C193 VDD2.n159 VSUBS 0.016671f
C194 VDD2.n160 VSUBS 0.037214f
C195 VDD2.n161 VSUBS 0.037214f
C196 VDD2.n162 VSUBS 0.016671f
C197 VDD2.n163 VSUBS 0.015744f
C198 VDD2.n164 VSUBS 0.0293f
C199 VDD2.n165 VSUBS 0.0293f
C200 VDD2.n166 VSUBS 0.015744f
C201 VDD2.n167 VSUBS 0.016671f
C202 VDD2.n168 VSUBS 0.037214f
C203 VDD2.n169 VSUBS 0.037214f
C204 VDD2.n170 VSUBS 0.016671f
C205 VDD2.n171 VSUBS 0.015744f
C206 VDD2.n172 VSUBS 0.0293f
C207 VDD2.n173 VSUBS 0.0293f
C208 VDD2.n174 VSUBS 0.015744f
C209 VDD2.n175 VSUBS 0.016671f
C210 VDD2.n176 VSUBS 0.037214f
C211 VDD2.n177 VSUBS 0.037214f
C212 VDD2.n178 VSUBS 0.016671f
C213 VDD2.n179 VSUBS 0.015744f
C214 VDD2.n180 VSUBS 0.0293f
C215 VDD2.n181 VSUBS 0.0293f
C216 VDD2.n182 VSUBS 0.015744f
C217 VDD2.n183 VSUBS 0.016671f
C218 VDD2.n184 VSUBS 0.037214f
C219 VDD2.n185 VSUBS 0.037214f
C220 VDD2.n186 VSUBS 0.016671f
C221 VDD2.n187 VSUBS 0.015744f
C222 VDD2.n188 VSUBS 0.0293f
C223 VDD2.n189 VSUBS 0.0293f
C224 VDD2.n190 VSUBS 0.015744f
C225 VDD2.n191 VSUBS 0.016671f
C226 VDD2.n192 VSUBS 0.037214f
C227 VDD2.n193 VSUBS 0.085444f
C228 VDD2.n194 VSUBS 0.016671f
C229 VDD2.n195 VSUBS 0.015744f
C230 VDD2.n196 VSUBS 0.065324f
C231 VDD2.n197 VSUBS 0.062938f
C232 VDD2.n198 VSUBS 4.39295f
C233 VDD2.t6 VSUBS 0.404264f
C234 VDD2.t2 VSUBS 0.404264f
C235 VDD2.n199 VSUBS 3.3387f
C236 VDD2.n200 VSUBS 1.00204f
C237 VDD2.t3 VSUBS 0.404264f
C238 VDD2.t7 VSUBS 0.404264f
C239 VDD2.n201 VSUBS 3.38138f
C240 VN.t4 VSUBS 3.71642f
C241 VN.n0 VSUBS 1.36236f
C242 VN.n1 VSUBS 0.020703f
C243 VN.n2 VSUBS 0.037611f
C244 VN.n3 VSUBS 0.020703f
C245 VN.n4 VSUBS 0.035739f
C246 VN.n5 VSUBS 0.020703f
C247 VN.n6 VSUBS 0.040063f
C248 VN.n7 VSUBS 0.020703f
C249 VN.n8 VSUBS 0.038392f
C250 VN.n9 VSUBS 0.020703f
C251 VN.t1 VSUBS 3.71642f
C252 VN.n10 VSUBS 0.041474f
C253 VN.n11 VSUBS 0.020703f
C254 VN.n12 VSUBS 0.038392f
C255 VN.t8 VSUBS 4.04229f
C256 VN.n13 VSUBS 1.28536f
C257 VN.t5 VSUBS 3.71642f
C258 VN.n14 VSUBS 1.34859f
C259 VN.n15 VSUBS 0.022093f
C260 VN.n16 VSUBS 0.262814f
C261 VN.n17 VSUBS 0.020703f
C262 VN.n18 VSUBS 0.020703f
C263 VN.n19 VSUBS 0.038392f
C264 VN.n20 VSUBS 0.040063f
C265 VN.n21 VSUBS 0.017047f
C266 VN.n22 VSUBS 0.020703f
C267 VN.n23 VSUBS 0.020703f
C268 VN.n24 VSUBS 0.020703f
C269 VN.n25 VSUBS 0.038392f
C270 VN.n26 VSUBS 0.038392f
C271 VN.n27 VSUBS 1.30131f
C272 VN.n28 VSUBS 0.020703f
C273 VN.n29 VSUBS 0.020703f
C274 VN.n30 VSUBS 0.020703f
C275 VN.n31 VSUBS 0.038392f
C276 VN.n32 VSUBS 0.041474f
C277 VN.n33 VSUBS 0.017047f
C278 VN.n34 VSUBS 0.020703f
C279 VN.n35 VSUBS 0.020703f
C280 VN.n36 VSUBS 0.020703f
C281 VN.n37 VSUBS 0.038392f
C282 VN.n38 VSUBS 0.038392f
C283 VN.t9 VSUBS 3.71642f
C284 VN.n39 VSUBS 1.28187f
C285 VN.n40 VSUBS 0.022093f
C286 VN.n41 VSUBS 0.020703f
C287 VN.n42 VSUBS 0.020703f
C288 VN.n43 VSUBS 0.020703f
C289 VN.n44 VSUBS 0.038392f
C290 VN.n45 VSUBS 0.041146f
C291 VN.n46 VSUBS 0.019826f
C292 VN.n47 VSUBS 0.020703f
C293 VN.n48 VSUBS 0.020703f
C294 VN.n49 VSUBS 0.020703f
C295 VN.n50 VSUBS 0.038392f
C296 VN.n51 VSUBS 0.038392f
C297 VN.n52 VSUBS 0.024746f
C298 VN.n53 VSUBS 0.033409f
C299 VN.n54 VSUBS 0.060249f
C300 VN.t0 VSUBS 3.71642f
C301 VN.n55 VSUBS 1.36236f
C302 VN.n56 VSUBS 0.020703f
C303 VN.n57 VSUBS 0.037611f
C304 VN.n58 VSUBS 0.020703f
C305 VN.n59 VSUBS 0.035739f
C306 VN.n60 VSUBS 0.020703f
C307 VN.t3 VSUBS 3.71642f
C308 VN.n61 VSUBS 1.28187f
C309 VN.n62 VSUBS 0.040063f
C310 VN.n63 VSUBS 0.020703f
C311 VN.n64 VSUBS 0.038392f
C312 VN.n65 VSUBS 0.020703f
C313 VN.t7 VSUBS 3.71642f
C314 VN.n66 VSUBS 0.041474f
C315 VN.n67 VSUBS 0.020703f
C316 VN.n68 VSUBS 0.038392f
C317 VN.t2 VSUBS 4.04229f
C318 VN.n69 VSUBS 1.28536f
C319 VN.t6 VSUBS 3.71642f
C320 VN.n70 VSUBS 1.34859f
C321 VN.n71 VSUBS 0.022093f
C322 VN.n72 VSUBS 0.262814f
C323 VN.n73 VSUBS 0.020703f
C324 VN.n74 VSUBS 0.020703f
C325 VN.n75 VSUBS 0.038392f
C326 VN.n76 VSUBS 0.040063f
C327 VN.n77 VSUBS 0.017047f
C328 VN.n78 VSUBS 0.020703f
C329 VN.n79 VSUBS 0.020703f
C330 VN.n80 VSUBS 0.020703f
C331 VN.n81 VSUBS 0.038392f
C332 VN.n82 VSUBS 0.038392f
C333 VN.n83 VSUBS 1.30131f
C334 VN.n84 VSUBS 0.020703f
C335 VN.n85 VSUBS 0.020703f
C336 VN.n86 VSUBS 0.020703f
C337 VN.n87 VSUBS 0.038392f
C338 VN.n88 VSUBS 0.041474f
C339 VN.n89 VSUBS 0.017047f
C340 VN.n90 VSUBS 0.020703f
C341 VN.n91 VSUBS 0.020703f
C342 VN.n92 VSUBS 0.020703f
C343 VN.n93 VSUBS 0.038392f
C344 VN.n94 VSUBS 0.038392f
C345 VN.n95 VSUBS 0.022093f
C346 VN.n96 VSUBS 0.020703f
C347 VN.n97 VSUBS 0.020703f
C348 VN.n98 VSUBS 0.020703f
C349 VN.n99 VSUBS 0.038392f
C350 VN.n100 VSUBS 0.041146f
C351 VN.n101 VSUBS 0.019826f
C352 VN.n102 VSUBS 0.020703f
C353 VN.n103 VSUBS 0.020703f
C354 VN.n104 VSUBS 0.020703f
C355 VN.n105 VSUBS 0.038392f
C356 VN.n106 VSUBS 0.038392f
C357 VN.n107 VSUBS 0.024746f
C358 VN.n108 VSUBS 0.033409f
C359 VN.n109 VSUBS 1.65482f
C360 VTAIL.t8 VSUBS 0.389513f
C361 VTAIL.t3 VSUBS 0.389513f
C362 VTAIL.n0 VSUBS 3.03572f
C363 VTAIL.n1 VSUBS 1.15101f
C364 VTAIL.n2 VSUBS 0.029705f
C365 VTAIL.n3 VSUBS 0.028231f
C366 VTAIL.n4 VSUBS 0.01517f
C367 VTAIL.n5 VSUBS 0.035857f
C368 VTAIL.n6 VSUBS 0.016062f
C369 VTAIL.n7 VSUBS 0.028231f
C370 VTAIL.n8 VSUBS 0.01517f
C371 VTAIL.n9 VSUBS 0.035857f
C372 VTAIL.n10 VSUBS 0.015616f
C373 VTAIL.n11 VSUBS 0.028231f
C374 VTAIL.n12 VSUBS 0.016062f
C375 VTAIL.n13 VSUBS 0.035857f
C376 VTAIL.n14 VSUBS 0.016062f
C377 VTAIL.n15 VSUBS 0.028231f
C378 VTAIL.n16 VSUBS 0.01517f
C379 VTAIL.n17 VSUBS 0.035857f
C380 VTAIL.n18 VSUBS 0.016062f
C381 VTAIL.n19 VSUBS 0.028231f
C382 VTAIL.n20 VSUBS 0.01517f
C383 VTAIL.n21 VSUBS 0.035857f
C384 VTAIL.n22 VSUBS 0.016062f
C385 VTAIL.n23 VSUBS 0.028231f
C386 VTAIL.n24 VSUBS 0.01517f
C387 VTAIL.n25 VSUBS 0.035857f
C388 VTAIL.n26 VSUBS 0.016062f
C389 VTAIL.n27 VSUBS 0.028231f
C390 VTAIL.n28 VSUBS 0.01517f
C391 VTAIL.n29 VSUBS 0.035857f
C392 VTAIL.n30 VSUBS 0.016062f
C393 VTAIL.n31 VSUBS 2.11787f
C394 VTAIL.n32 VSUBS 0.01517f
C395 VTAIL.t16 VSUBS 0.076934f
C396 VTAIL.n33 VSUBS 0.219487f
C397 VTAIL.n34 VSUBS 0.02281f
C398 VTAIL.n35 VSUBS 0.026892f
C399 VTAIL.n36 VSUBS 0.035857f
C400 VTAIL.n37 VSUBS 0.016062f
C401 VTAIL.n38 VSUBS 0.01517f
C402 VTAIL.n39 VSUBS 0.028231f
C403 VTAIL.n40 VSUBS 0.028231f
C404 VTAIL.n41 VSUBS 0.01517f
C405 VTAIL.n42 VSUBS 0.016062f
C406 VTAIL.n43 VSUBS 0.035857f
C407 VTAIL.n44 VSUBS 0.035857f
C408 VTAIL.n45 VSUBS 0.016062f
C409 VTAIL.n46 VSUBS 0.01517f
C410 VTAIL.n47 VSUBS 0.028231f
C411 VTAIL.n48 VSUBS 0.028231f
C412 VTAIL.n49 VSUBS 0.01517f
C413 VTAIL.n50 VSUBS 0.016062f
C414 VTAIL.n51 VSUBS 0.035857f
C415 VTAIL.n52 VSUBS 0.035857f
C416 VTAIL.n53 VSUBS 0.016062f
C417 VTAIL.n54 VSUBS 0.01517f
C418 VTAIL.n55 VSUBS 0.028231f
C419 VTAIL.n56 VSUBS 0.028231f
C420 VTAIL.n57 VSUBS 0.01517f
C421 VTAIL.n58 VSUBS 0.016062f
C422 VTAIL.n59 VSUBS 0.035857f
C423 VTAIL.n60 VSUBS 0.035857f
C424 VTAIL.n61 VSUBS 0.016062f
C425 VTAIL.n62 VSUBS 0.01517f
C426 VTAIL.n63 VSUBS 0.028231f
C427 VTAIL.n64 VSUBS 0.028231f
C428 VTAIL.n65 VSUBS 0.01517f
C429 VTAIL.n66 VSUBS 0.016062f
C430 VTAIL.n67 VSUBS 0.035857f
C431 VTAIL.n68 VSUBS 0.035857f
C432 VTAIL.n69 VSUBS 0.016062f
C433 VTAIL.n70 VSUBS 0.01517f
C434 VTAIL.n71 VSUBS 0.028231f
C435 VTAIL.n72 VSUBS 0.028231f
C436 VTAIL.n73 VSUBS 0.01517f
C437 VTAIL.n74 VSUBS 0.01517f
C438 VTAIL.n75 VSUBS 0.016062f
C439 VTAIL.n76 VSUBS 0.035857f
C440 VTAIL.n77 VSUBS 0.035857f
C441 VTAIL.n78 VSUBS 0.035857f
C442 VTAIL.n79 VSUBS 0.015616f
C443 VTAIL.n80 VSUBS 0.01517f
C444 VTAIL.n81 VSUBS 0.028231f
C445 VTAIL.n82 VSUBS 0.028231f
C446 VTAIL.n83 VSUBS 0.01517f
C447 VTAIL.n84 VSUBS 0.016062f
C448 VTAIL.n85 VSUBS 0.035857f
C449 VTAIL.n86 VSUBS 0.035857f
C450 VTAIL.n87 VSUBS 0.016062f
C451 VTAIL.n88 VSUBS 0.01517f
C452 VTAIL.n89 VSUBS 0.028231f
C453 VTAIL.n90 VSUBS 0.028231f
C454 VTAIL.n91 VSUBS 0.01517f
C455 VTAIL.n92 VSUBS 0.016062f
C456 VTAIL.n93 VSUBS 0.035857f
C457 VTAIL.n94 VSUBS 0.082326f
C458 VTAIL.n95 VSUBS 0.016062f
C459 VTAIL.n96 VSUBS 0.01517f
C460 VTAIL.n97 VSUBS 0.06294f
C461 VTAIL.n98 VSUBS 0.04113f
C462 VTAIL.n99 VSUBS 0.544294f
C463 VTAIL.t14 VSUBS 0.389513f
C464 VTAIL.t19 VSUBS 0.389513f
C465 VTAIL.n100 VSUBS 3.03572f
C466 VTAIL.n101 VSUBS 1.34236f
C467 VTAIL.t10 VSUBS 0.389513f
C468 VTAIL.t17 VSUBS 0.389513f
C469 VTAIL.n102 VSUBS 3.03572f
C470 VTAIL.n103 VSUBS 3.41421f
C471 VTAIL.t2 VSUBS 0.389513f
C472 VTAIL.t1 VSUBS 0.389513f
C473 VTAIL.n104 VSUBS 3.03574f
C474 VTAIL.n105 VSUBS 3.41419f
C475 VTAIL.t5 VSUBS 0.389513f
C476 VTAIL.t9 VSUBS 0.389513f
C477 VTAIL.n106 VSUBS 3.03574f
C478 VTAIL.n107 VSUBS 1.34234f
C479 VTAIL.n108 VSUBS 0.029705f
C480 VTAIL.n109 VSUBS 0.028231f
C481 VTAIL.n110 VSUBS 0.01517f
C482 VTAIL.n111 VSUBS 0.035857f
C483 VTAIL.n112 VSUBS 0.016062f
C484 VTAIL.n113 VSUBS 0.028231f
C485 VTAIL.n114 VSUBS 0.01517f
C486 VTAIL.n115 VSUBS 0.035857f
C487 VTAIL.n116 VSUBS 0.015616f
C488 VTAIL.n117 VSUBS 0.028231f
C489 VTAIL.n118 VSUBS 0.015616f
C490 VTAIL.n119 VSUBS 0.01517f
C491 VTAIL.n120 VSUBS 0.035857f
C492 VTAIL.n121 VSUBS 0.035857f
C493 VTAIL.n122 VSUBS 0.016062f
C494 VTAIL.n123 VSUBS 0.028231f
C495 VTAIL.n124 VSUBS 0.01517f
C496 VTAIL.n125 VSUBS 0.035857f
C497 VTAIL.n126 VSUBS 0.016062f
C498 VTAIL.n127 VSUBS 0.028231f
C499 VTAIL.n128 VSUBS 0.01517f
C500 VTAIL.n129 VSUBS 0.035857f
C501 VTAIL.n130 VSUBS 0.016062f
C502 VTAIL.n131 VSUBS 0.028231f
C503 VTAIL.n132 VSUBS 0.01517f
C504 VTAIL.n133 VSUBS 0.035857f
C505 VTAIL.n134 VSUBS 0.016062f
C506 VTAIL.n135 VSUBS 0.028231f
C507 VTAIL.n136 VSUBS 0.01517f
C508 VTAIL.n137 VSUBS 0.035857f
C509 VTAIL.n138 VSUBS 0.016062f
C510 VTAIL.n139 VSUBS 2.11787f
C511 VTAIL.n140 VSUBS 0.01517f
C512 VTAIL.t4 VSUBS 0.076934f
C513 VTAIL.n141 VSUBS 0.219487f
C514 VTAIL.n142 VSUBS 0.02281f
C515 VTAIL.n143 VSUBS 0.026892f
C516 VTAIL.n144 VSUBS 0.035857f
C517 VTAIL.n145 VSUBS 0.016062f
C518 VTAIL.n146 VSUBS 0.01517f
C519 VTAIL.n147 VSUBS 0.028231f
C520 VTAIL.n148 VSUBS 0.028231f
C521 VTAIL.n149 VSUBS 0.01517f
C522 VTAIL.n150 VSUBS 0.016062f
C523 VTAIL.n151 VSUBS 0.035857f
C524 VTAIL.n152 VSUBS 0.035857f
C525 VTAIL.n153 VSUBS 0.016062f
C526 VTAIL.n154 VSUBS 0.01517f
C527 VTAIL.n155 VSUBS 0.028231f
C528 VTAIL.n156 VSUBS 0.028231f
C529 VTAIL.n157 VSUBS 0.01517f
C530 VTAIL.n158 VSUBS 0.016062f
C531 VTAIL.n159 VSUBS 0.035857f
C532 VTAIL.n160 VSUBS 0.035857f
C533 VTAIL.n161 VSUBS 0.016062f
C534 VTAIL.n162 VSUBS 0.01517f
C535 VTAIL.n163 VSUBS 0.028231f
C536 VTAIL.n164 VSUBS 0.028231f
C537 VTAIL.n165 VSUBS 0.01517f
C538 VTAIL.n166 VSUBS 0.016062f
C539 VTAIL.n167 VSUBS 0.035857f
C540 VTAIL.n168 VSUBS 0.035857f
C541 VTAIL.n169 VSUBS 0.016062f
C542 VTAIL.n170 VSUBS 0.01517f
C543 VTAIL.n171 VSUBS 0.028231f
C544 VTAIL.n172 VSUBS 0.028231f
C545 VTAIL.n173 VSUBS 0.01517f
C546 VTAIL.n174 VSUBS 0.016062f
C547 VTAIL.n175 VSUBS 0.035857f
C548 VTAIL.n176 VSUBS 0.035857f
C549 VTAIL.n177 VSUBS 0.016062f
C550 VTAIL.n178 VSUBS 0.01517f
C551 VTAIL.n179 VSUBS 0.028231f
C552 VTAIL.n180 VSUBS 0.028231f
C553 VTAIL.n181 VSUBS 0.01517f
C554 VTAIL.n182 VSUBS 0.016062f
C555 VTAIL.n183 VSUBS 0.035857f
C556 VTAIL.n184 VSUBS 0.035857f
C557 VTAIL.n185 VSUBS 0.016062f
C558 VTAIL.n186 VSUBS 0.01517f
C559 VTAIL.n187 VSUBS 0.028231f
C560 VTAIL.n188 VSUBS 0.028231f
C561 VTAIL.n189 VSUBS 0.01517f
C562 VTAIL.n190 VSUBS 0.016062f
C563 VTAIL.n191 VSUBS 0.035857f
C564 VTAIL.n192 VSUBS 0.035857f
C565 VTAIL.n193 VSUBS 0.016062f
C566 VTAIL.n194 VSUBS 0.01517f
C567 VTAIL.n195 VSUBS 0.028231f
C568 VTAIL.n196 VSUBS 0.028231f
C569 VTAIL.n197 VSUBS 0.01517f
C570 VTAIL.n198 VSUBS 0.016062f
C571 VTAIL.n199 VSUBS 0.035857f
C572 VTAIL.n200 VSUBS 0.082326f
C573 VTAIL.n201 VSUBS 0.016062f
C574 VTAIL.n202 VSUBS 0.01517f
C575 VTAIL.n203 VSUBS 0.06294f
C576 VTAIL.n204 VSUBS 0.04113f
C577 VTAIL.n205 VSUBS 0.544294f
C578 VTAIL.t12 VSUBS 0.389513f
C579 VTAIL.t11 VSUBS 0.389513f
C580 VTAIL.n206 VSUBS 3.03574f
C581 VTAIL.n207 VSUBS 1.22549f
C582 VTAIL.t13 VSUBS 0.389513f
C583 VTAIL.t15 VSUBS 0.389513f
C584 VTAIL.n208 VSUBS 3.03574f
C585 VTAIL.n209 VSUBS 1.34234f
C586 VTAIL.n210 VSUBS 0.029705f
C587 VTAIL.n211 VSUBS 0.028231f
C588 VTAIL.n212 VSUBS 0.01517f
C589 VTAIL.n213 VSUBS 0.035857f
C590 VTAIL.n214 VSUBS 0.016062f
C591 VTAIL.n215 VSUBS 0.028231f
C592 VTAIL.n216 VSUBS 0.01517f
C593 VTAIL.n217 VSUBS 0.035857f
C594 VTAIL.n218 VSUBS 0.015616f
C595 VTAIL.n219 VSUBS 0.028231f
C596 VTAIL.n220 VSUBS 0.015616f
C597 VTAIL.n221 VSUBS 0.01517f
C598 VTAIL.n222 VSUBS 0.035857f
C599 VTAIL.n223 VSUBS 0.035857f
C600 VTAIL.n224 VSUBS 0.016062f
C601 VTAIL.n225 VSUBS 0.028231f
C602 VTAIL.n226 VSUBS 0.01517f
C603 VTAIL.n227 VSUBS 0.035857f
C604 VTAIL.n228 VSUBS 0.016062f
C605 VTAIL.n229 VSUBS 0.028231f
C606 VTAIL.n230 VSUBS 0.01517f
C607 VTAIL.n231 VSUBS 0.035857f
C608 VTAIL.n232 VSUBS 0.016062f
C609 VTAIL.n233 VSUBS 0.028231f
C610 VTAIL.n234 VSUBS 0.01517f
C611 VTAIL.n235 VSUBS 0.035857f
C612 VTAIL.n236 VSUBS 0.016062f
C613 VTAIL.n237 VSUBS 0.028231f
C614 VTAIL.n238 VSUBS 0.01517f
C615 VTAIL.n239 VSUBS 0.035857f
C616 VTAIL.n240 VSUBS 0.016062f
C617 VTAIL.n241 VSUBS 2.11787f
C618 VTAIL.n242 VSUBS 0.01517f
C619 VTAIL.t18 VSUBS 0.076934f
C620 VTAIL.n243 VSUBS 0.219487f
C621 VTAIL.n244 VSUBS 0.02281f
C622 VTAIL.n245 VSUBS 0.026892f
C623 VTAIL.n246 VSUBS 0.035857f
C624 VTAIL.n247 VSUBS 0.016062f
C625 VTAIL.n248 VSUBS 0.01517f
C626 VTAIL.n249 VSUBS 0.028231f
C627 VTAIL.n250 VSUBS 0.028231f
C628 VTAIL.n251 VSUBS 0.01517f
C629 VTAIL.n252 VSUBS 0.016062f
C630 VTAIL.n253 VSUBS 0.035857f
C631 VTAIL.n254 VSUBS 0.035857f
C632 VTAIL.n255 VSUBS 0.016062f
C633 VTAIL.n256 VSUBS 0.01517f
C634 VTAIL.n257 VSUBS 0.028231f
C635 VTAIL.n258 VSUBS 0.028231f
C636 VTAIL.n259 VSUBS 0.01517f
C637 VTAIL.n260 VSUBS 0.016062f
C638 VTAIL.n261 VSUBS 0.035857f
C639 VTAIL.n262 VSUBS 0.035857f
C640 VTAIL.n263 VSUBS 0.016062f
C641 VTAIL.n264 VSUBS 0.01517f
C642 VTAIL.n265 VSUBS 0.028231f
C643 VTAIL.n266 VSUBS 0.028231f
C644 VTAIL.n267 VSUBS 0.01517f
C645 VTAIL.n268 VSUBS 0.016062f
C646 VTAIL.n269 VSUBS 0.035857f
C647 VTAIL.n270 VSUBS 0.035857f
C648 VTAIL.n271 VSUBS 0.016062f
C649 VTAIL.n272 VSUBS 0.01517f
C650 VTAIL.n273 VSUBS 0.028231f
C651 VTAIL.n274 VSUBS 0.028231f
C652 VTAIL.n275 VSUBS 0.01517f
C653 VTAIL.n276 VSUBS 0.016062f
C654 VTAIL.n277 VSUBS 0.035857f
C655 VTAIL.n278 VSUBS 0.035857f
C656 VTAIL.n279 VSUBS 0.016062f
C657 VTAIL.n280 VSUBS 0.01517f
C658 VTAIL.n281 VSUBS 0.028231f
C659 VTAIL.n282 VSUBS 0.028231f
C660 VTAIL.n283 VSUBS 0.01517f
C661 VTAIL.n284 VSUBS 0.016062f
C662 VTAIL.n285 VSUBS 0.035857f
C663 VTAIL.n286 VSUBS 0.035857f
C664 VTAIL.n287 VSUBS 0.016062f
C665 VTAIL.n288 VSUBS 0.01517f
C666 VTAIL.n289 VSUBS 0.028231f
C667 VTAIL.n290 VSUBS 0.028231f
C668 VTAIL.n291 VSUBS 0.01517f
C669 VTAIL.n292 VSUBS 0.016062f
C670 VTAIL.n293 VSUBS 0.035857f
C671 VTAIL.n294 VSUBS 0.035857f
C672 VTAIL.n295 VSUBS 0.016062f
C673 VTAIL.n296 VSUBS 0.01517f
C674 VTAIL.n297 VSUBS 0.028231f
C675 VTAIL.n298 VSUBS 0.028231f
C676 VTAIL.n299 VSUBS 0.01517f
C677 VTAIL.n300 VSUBS 0.016062f
C678 VTAIL.n301 VSUBS 0.035857f
C679 VTAIL.n302 VSUBS 0.082326f
C680 VTAIL.n303 VSUBS 0.016062f
C681 VTAIL.n304 VSUBS 0.01517f
C682 VTAIL.n305 VSUBS 0.06294f
C683 VTAIL.n306 VSUBS 0.04113f
C684 VTAIL.n307 VSUBS 2.41382f
C685 VTAIL.n308 VSUBS 0.029705f
C686 VTAIL.n309 VSUBS 0.028231f
C687 VTAIL.n310 VSUBS 0.01517f
C688 VTAIL.n311 VSUBS 0.035857f
C689 VTAIL.n312 VSUBS 0.016062f
C690 VTAIL.n313 VSUBS 0.028231f
C691 VTAIL.n314 VSUBS 0.01517f
C692 VTAIL.n315 VSUBS 0.035857f
C693 VTAIL.n316 VSUBS 0.015616f
C694 VTAIL.n317 VSUBS 0.028231f
C695 VTAIL.n318 VSUBS 0.016062f
C696 VTAIL.n319 VSUBS 0.035857f
C697 VTAIL.n320 VSUBS 0.016062f
C698 VTAIL.n321 VSUBS 0.028231f
C699 VTAIL.n322 VSUBS 0.01517f
C700 VTAIL.n323 VSUBS 0.035857f
C701 VTAIL.n324 VSUBS 0.016062f
C702 VTAIL.n325 VSUBS 0.028231f
C703 VTAIL.n326 VSUBS 0.01517f
C704 VTAIL.n327 VSUBS 0.035857f
C705 VTAIL.n328 VSUBS 0.016062f
C706 VTAIL.n329 VSUBS 0.028231f
C707 VTAIL.n330 VSUBS 0.01517f
C708 VTAIL.n331 VSUBS 0.035857f
C709 VTAIL.n332 VSUBS 0.016062f
C710 VTAIL.n333 VSUBS 0.028231f
C711 VTAIL.n334 VSUBS 0.01517f
C712 VTAIL.n335 VSUBS 0.035857f
C713 VTAIL.n336 VSUBS 0.016062f
C714 VTAIL.n337 VSUBS 2.11787f
C715 VTAIL.n338 VSUBS 0.01517f
C716 VTAIL.t0 VSUBS 0.076934f
C717 VTAIL.n339 VSUBS 0.219487f
C718 VTAIL.n340 VSUBS 0.02281f
C719 VTAIL.n341 VSUBS 0.026892f
C720 VTAIL.n342 VSUBS 0.035857f
C721 VTAIL.n343 VSUBS 0.016062f
C722 VTAIL.n344 VSUBS 0.01517f
C723 VTAIL.n345 VSUBS 0.028231f
C724 VTAIL.n346 VSUBS 0.028231f
C725 VTAIL.n347 VSUBS 0.01517f
C726 VTAIL.n348 VSUBS 0.016062f
C727 VTAIL.n349 VSUBS 0.035857f
C728 VTAIL.n350 VSUBS 0.035857f
C729 VTAIL.n351 VSUBS 0.016062f
C730 VTAIL.n352 VSUBS 0.01517f
C731 VTAIL.n353 VSUBS 0.028231f
C732 VTAIL.n354 VSUBS 0.028231f
C733 VTAIL.n355 VSUBS 0.01517f
C734 VTAIL.n356 VSUBS 0.016062f
C735 VTAIL.n357 VSUBS 0.035857f
C736 VTAIL.n358 VSUBS 0.035857f
C737 VTAIL.n359 VSUBS 0.016062f
C738 VTAIL.n360 VSUBS 0.01517f
C739 VTAIL.n361 VSUBS 0.028231f
C740 VTAIL.n362 VSUBS 0.028231f
C741 VTAIL.n363 VSUBS 0.01517f
C742 VTAIL.n364 VSUBS 0.016062f
C743 VTAIL.n365 VSUBS 0.035857f
C744 VTAIL.n366 VSUBS 0.035857f
C745 VTAIL.n367 VSUBS 0.016062f
C746 VTAIL.n368 VSUBS 0.01517f
C747 VTAIL.n369 VSUBS 0.028231f
C748 VTAIL.n370 VSUBS 0.028231f
C749 VTAIL.n371 VSUBS 0.01517f
C750 VTAIL.n372 VSUBS 0.016062f
C751 VTAIL.n373 VSUBS 0.035857f
C752 VTAIL.n374 VSUBS 0.035857f
C753 VTAIL.n375 VSUBS 0.016062f
C754 VTAIL.n376 VSUBS 0.01517f
C755 VTAIL.n377 VSUBS 0.028231f
C756 VTAIL.n378 VSUBS 0.028231f
C757 VTAIL.n379 VSUBS 0.01517f
C758 VTAIL.n380 VSUBS 0.01517f
C759 VTAIL.n381 VSUBS 0.016062f
C760 VTAIL.n382 VSUBS 0.035857f
C761 VTAIL.n383 VSUBS 0.035857f
C762 VTAIL.n384 VSUBS 0.035857f
C763 VTAIL.n385 VSUBS 0.015616f
C764 VTAIL.n386 VSUBS 0.01517f
C765 VTAIL.n387 VSUBS 0.028231f
C766 VTAIL.n388 VSUBS 0.028231f
C767 VTAIL.n389 VSUBS 0.01517f
C768 VTAIL.n390 VSUBS 0.016062f
C769 VTAIL.n391 VSUBS 0.035857f
C770 VTAIL.n392 VSUBS 0.035857f
C771 VTAIL.n393 VSUBS 0.016062f
C772 VTAIL.n394 VSUBS 0.01517f
C773 VTAIL.n395 VSUBS 0.028231f
C774 VTAIL.n396 VSUBS 0.028231f
C775 VTAIL.n397 VSUBS 0.01517f
C776 VTAIL.n398 VSUBS 0.016062f
C777 VTAIL.n399 VSUBS 0.035857f
C778 VTAIL.n400 VSUBS 0.082326f
C779 VTAIL.n401 VSUBS 0.016062f
C780 VTAIL.n402 VSUBS 0.01517f
C781 VTAIL.n403 VSUBS 0.06294f
C782 VTAIL.n404 VSUBS 0.04113f
C783 VTAIL.n405 VSUBS 2.41382f
C784 VTAIL.t7 VSUBS 0.389513f
C785 VTAIL.t6 VSUBS 0.389513f
C786 VTAIL.n406 VSUBS 3.03572f
C787 VTAIL.n407 VSUBS 1.09769f
C788 VDD1.n0 VSUBS 0.030823f
C789 VDD1.n1 VSUBS 0.029294f
C790 VDD1.n2 VSUBS 0.015741f
C791 VDD1.n3 VSUBS 0.037207f
C792 VDD1.n4 VSUBS 0.016667f
C793 VDD1.n5 VSUBS 0.029294f
C794 VDD1.n6 VSUBS 0.015741f
C795 VDD1.n7 VSUBS 0.037207f
C796 VDD1.n8 VSUBS 0.016204f
C797 VDD1.n9 VSUBS 0.029294f
C798 VDD1.n10 VSUBS 0.016204f
C799 VDD1.n11 VSUBS 0.015741f
C800 VDD1.n12 VSUBS 0.037207f
C801 VDD1.n13 VSUBS 0.037207f
C802 VDD1.n14 VSUBS 0.016667f
C803 VDD1.n15 VSUBS 0.029294f
C804 VDD1.n16 VSUBS 0.015741f
C805 VDD1.n17 VSUBS 0.037207f
C806 VDD1.n18 VSUBS 0.016667f
C807 VDD1.n19 VSUBS 0.029294f
C808 VDD1.n20 VSUBS 0.015741f
C809 VDD1.n21 VSUBS 0.037207f
C810 VDD1.n22 VSUBS 0.016667f
C811 VDD1.n23 VSUBS 0.029294f
C812 VDD1.n24 VSUBS 0.015741f
C813 VDD1.n25 VSUBS 0.037207f
C814 VDD1.n26 VSUBS 0.016667f
C815 VDD1.n27 VSUBS 0.029294f
C816 VDD1.n28 VSUBS 0.015741f
C817 VDD1.n29 VSUBS 0.037207f
C818 VDD1.n30 VSUBS 0.016667f
C819 VDD1.n31 VSUBS 2.19762f
C820 VDD1.n32 VSUBS 0.015741f
C821 VDD1.t7 VSUBS 0.079831f
C822 VDD1.n33 VSUBS 0.227752f
C823 VDD1.n34 VSUBS 0.023669f
C824 VDD1.n35 VSUBS 0.027905f
C825 VDD1.n36 VSUBS 0.037207f
C826 VDD1.n37 VSUBS 0.016667f
C827 VDD1.n38 VSUBS 0.015741f
C828 VDD1.n39 VSUBS 0.029294f
C829 VDD1.n40 VSUBS 0.029294f
C830 VDD1.n41 VSUBS 0.015741f
C831 VDD1.n42 VSUBS 0.016667f
C832 VDD1.n43 VSUBS 0.037207f
C833 VDD1.n44 VSUBS 0.037207f
C834 VDD1.n45 VSUBS 0.016667f
C835 VDD1.n46 VSUBS 0.015741f
C836 VDD1.n47 VSUBS 0.029294f
C837 VDD1.n48 VSUBS 0.029294f
C838 VDD1.n49 VSUBS 0.015741f
C839 VDD1.n50 VSUBS 0.016667f
C840 VDD1.n51 VSUBS 0.037207f
C841 VDD1.n52 VSUBS 0.037207f
C842 VDD1.n53 VSUBS 0.016667f
C843 VDD1.n54 VSUBS 0.015741f
C844 VDD1.n55 VSUBS 0.029294f
C845 VDD1.n56 VSUBS 0.029294f
C846 VDD1.n57 VSUBS 0.015741f
C847 VDD1.n58 VSUBS 0.016667f
C848 VDD1.n59 VSUBS 0.037207f
C849 VDD1.n60 VSUBS 0.037207f
C850 VDD1.n61 VSUBS 0.016667f
C851 VDD1.n62 VSUBS 0.015741f
C852 VDD1.n63 VSUBS 0.029294f
C853 VDD1.n64 VSUBS 0.029294f
C854 VDD1.n65 VSUBS 0.015741f
C855 VDD1.n66 VSUBS 0.016667f
C856 VDD1.n67 VSUBS 0.037207f
C857 VDD1.n68 VSUBS 0.037207f
C858 VDD1.n69 VSUBS 0.016667f
C859 VDD1.n70 VSUBS 0.015741f
C860 VDD1.n71 VSUBS 0.029294f
C861 VDD1.n72 VSUBS 0.029294f
C862 VDD1.n73 VSUBS 0.015741f
C863 VDD1.n74 VSUBS 0.016667f
C864 VDD1.n75 VSUBS 0.037207f
C865 VDD1.n76 VSUBS 0.037207f
C866 VDD1.n77 VSUBS 0.016667f
C867 VDD1.n78 VSUBS 0.015741f
C868 VDD1.n79 VSUBS 0.029294f
C869 VDD1.n80 VSUBS 0.029294f
C870 VDD1.n81 VSUBS 0.015741f
C871 VDD1.n82 VSUBS 0.016667f
C872 VDD1.n83 VSUBS 0.037207f
C873 VDD1.n84 VSUBS 0.037207f
C874 VDD1.n85 VSUBS 0.016667f
C875 VDD1.n86 VSUBS 0.015741f
C876 VDD1.n87 VSUBS 0.029294f
C877 VDD1.n88 VSUBS 0.029294f
C878 VDD1.n89 VSUBS 0.015741f
C879 VDD1.n90 VSUBS 0.016667f
C880 VDD1.n91 VSUBS 0.037207f
C881 VDD1.n92 VSUBS 0.085426f
C882 VDD1.n93 VSUBS 0.016667f
C883 VDD1.n94 VSUBS 0.015741f
C884 VDD1.n95 VSUBS 0.06531f
C885 VDD1.n96 VSUBS 0.089388f
C886 VDD1.t9 VSUBS 0.404181f
C887 VDD1.t8 VSUBS 0.404181f
C888 VDD1.n97 VSUBS 3.33801f
C889 VDD1.n98 VSUBS 1.36159f
C890 VDD1.n99 VSUBS 0.030823f
C891 VDD1.n100 VSUBS 0.029294f
C892 VDD1.n101 VSUBS 0.015741f
C893 VDD1.n102 VSUBS 0.037207f
C894 VDD1.n103 VSUBS 0.016667f
C895 VDD1.n104 VSUBS 0.029294f
C896 VDD1.n105 VSUBS 0.015741f
C897 VDD1.n106 VSUBS 0.037207f
C898 VDD1.n107 VSUBS 0.016204f
C899 VDD1.n108 VSUBS 0.029294f
C900 VDD1.n109 VSUBS 0.016667f
C901 VDD1.n110 VSUBS 0.037207f
C902 VDD1.n111 VSUBS 0.016667f
C903 VDD1.n112 VSUBS 0.029294f
C904 VDD1.n113 VSUBS 0.015741f
C905 VDD1.n114 VSUBS 0.037207f
C906 VDD1.n115 VSUBS 0.016667f
C907 VDD1.n116 VSUBS 0.029294f
C908 VDD1.n117 VSUBS 0.015741f
C909 VDD1.n118 VSUBS 0.037207f
C910 VDD1.n119 VSUBS 0.016667f
C911 VDD1.n120 VSUBS 0.029294f
C912 VDD1.n121 VSUBS 0.015741f
C913 VDD1.n122 VSUBS 0.037207f
C914 VDD1.n123 VSUBS 0.016667f
C915 VDD1.n124 VSUBS 0.029294f
C916 VDD1.n125 VSUBS 0.015741f
C917 VDD1.n126 VSUBS 0.037207f
C918 VDD1.n127 VSUBS 0.016667f
C919 VDD1.n128 VSUBS 2.19762f
C920 VDD1.n129 VSUBS 0.015741f
C921 VDD1.t6 VSUBS 0.079831f
C922 VDD1.n130 VSUBS 0.227752f
C923 VDD1.n131 VSUBS 0.023669f
C924 VDD1.n132 VSUBS 0.027905f
C925 VDD1.n133 VSUBS 0.037207f
C926 VDD1.n134 VSUBS 0.016667f
C927 VDD1.n135 VSUBS 0.015741f
C928 VDD1.n136 VSUBS 0.029294f
C929 VDD1.n137 VSUBS 0.029294f
C930 VDD1.n138 VSUBS 0.015741f
C931 VDD1.n139 VSUBS 0.016667f
C932 VDD1.n140 VSUBS 0.037207f
C933 VDD1.n141 VSUBS 0.037207f
C934 VDD1.n142 VSUBS 0.016667f
C935 VDD1.n143 VSUBS 0.015741f
C936 VDD1.n144 VSUBS 0.029294f
C937 VDD1.n145 VSUBS 0.029294f
C938 VDD1.n146 VSUBS 0.015741f
C939 VDD1.n147 VSUBS 0.016667f
C940 VDD1.n148 VSUBS 0.037207f
C941 VDD1.n149 VSUBS 0.037207f
C942 VDD1.n150 VSUBS 0.016667f
C943 VDD1.n151 VSUBS 0.015741f
C944 VDD1.n152 VSUBS 0.029294f
C945 VDD1.n153 VSUBS 0.029294f
C946 VDD1.n154 VSUBS 0.015741f
C947 VDD1.n155 VSUBS 0.016667f
C948 VDD1.n156 VSUBS 0.037207f
C949 VDD1.n157 VSUBS 0.037207f
C950 VDD1.n158 VSUBS 0.016667f
C951 VDD1.n159 VSUBS 0.015741f
C952 VDD1.n160 VSUBS 0.029294f
C953 VDD1.n161 VSUBS 0.029294f
C954 VDD1.n162 VSUBS 0.015741f
C955 VDD1.n163 VSUBS 0.016667f
C956 VDD1.n164 VSUBS 0.037207f
C957 VDD1.n165 VSUBS 0.037207f
C958 VDD1.n166 VSUBS 0.016667f
C959 VDD1.n167 VSUBS 0.015741f
C960 VDD1.n168 VSUBS 0.029294f
C961 VDD1.n169 VSUBS 0.029294f
C962 VDD1.n170 VSUBS 0.015741f
C963 VDD1.n171 VSUBS 0.015741f
C964 VDD1.n172 VSUBS 0.016667f
C965 VDD1.n173 VSUBS 0.037207f
C966 VDD1.n174 VSUBS 0.037207f
C967 VDD1.n175 VSUBS 0.037207f
C968 VDD1.n176 VSUBS 0.016204f
C969 VDD1.n177 VSUBS 0.015741f
C970 VDD1.n178 VSUBS 0.029294f
C971 VDD1.n179 VSUBS 0.029294f
C972 VDD1.n180 VSUBS 0.015741f
C973 VDD1.n181 VSUBS 0.016667f
C974 VDD1.n182 VSUBS 0.037207f
C975 VDD1.n183 VSUBS 0.037207f
C976 VDD1.n184 VSUBS 0.016667f
C977 VDD1.n185 VSUBS 0.015741f
C978 VDD1.n186 VSUBS 0.029294f
C979 VDD1.n187 VSUBS 0.029294f
C980 VDD1.n188 VSUBS 0.015741f
C981 VDD1.n189 VSUBS 0.016667f
C982 VDD1.n190 VSUBS 0.037207f
C983 VDD1.n191 VSUBS 0.085426f
C984 VDD1.n192 VSUBS 0.016667f
C985 VDD1.n193 VSUBS 0.015741f
C986 VDD1.n194 VSUBS 0.06531f
C987 VDD1.n195 VSUBS 0.089388f
C988 VDD1.t3 VSUBS 0.404181f
C989 VDD1.t5 VSUBS 0.404181f
C990 VDD1.n196 VSUBS 3.338f
C991 VDD1.n197 VSUBS 1.35172f
C992 VDD1.t1 VSUBS 0.404181f
C993 VDD1.t0 VSUBS 0.404181f
C994 VDD1.n198 VSUBS 3.38075f
C995 VDD1.n199 VSUBS 5.02113f
C996 VDD1.t4 VSUBS 0.404181f
C997 VDD1.t2 VSUBS 0.404181f
C998 VDD1.n200 VSUBS 3.338f
C999 VDD1.n201 VSUBS 5.09434f
C1000 VP.t3 VSUBS 3.9899f
C1001 VP.n0 VSUBS 1.46262f
C1002 VP.n1 VSUBS 0.022227f
C1003 VP.n2 VSUBS 0.040378f
C1004 VP.n3 VSUBS 0.022227f
C1005 VP.n4 VSUBS 0.038369f
C1006 VP.n5 VSUBS 0.022227f
C1007 VP.n6 VSUBS 0.043011f
C1008 VP.n7 VSUBS 0.022227f
C1009 VP.n8 VSUBS 0.041217f
C1010 VP.n9 VSUBS 0.022227f
C1011 VP.t5 VSUBS 3.9899f
C1012 VP.n10 VSUBS 0.044525f
C1013 VP.n11 VSUBS 0.022227f
C1014 VP.n12 VSUBS 0.041217f
C1015 VP.n13 VSUBS 0.022227f
C1016 VP.t2 VSUBS 3.9899f
C1017 VP.n14 VSUBS 0.044174f
C1018 VP.n15 VSUBS 0.022227f
C1019 VP.n16 VSUBS 0.041217f
C1020 VP.t1 VSUBS 3.9899f
C1021 VP.n17 VSUBS 1.46262f
C1022 VP.n18 VSUBS 0.022227f
C1023 VP.n19 VSUBS 0.040378f
C1024 VP.n20 VSUBS 0.022227f
C1025 VP.n21 VSUBS 0.038369f
C1026 VP.n22 VSUBS 0.022227f
C1027 VP.n23 VSUBS 0.043011f
C1028 VP.n24 VSUBS 0.022227f
C1029 VP.n25 VSUBS 0.041217f
C1030 VP.n26 VSUBS 0.022227f
C1031 VP.t6 VSUBS 3.9899f
C1032 VP.n27 VSUBS 0.044525f
C1033 VP.n28 VSUBS 0.022227f
C1034 VP.n29 VSUBS 0.041217f
C1035 VP.t7 VSUBS 4.33974f
C1036 VP.n30 VSUBS 1.37995f
C1037 VP.t8 VSUBS 3.9899f
C1038 VP.n31 VSUBS 1.44783f
C1039 VP.n32 VSUBS 0.023718f
C1040 VP.n33 VSUBS 0.282154f
C1041 VP.n34 VSUBS 0.022227f
C1042 VP.n35 VSUBS 0.022227f
C1043 VP.n36 VSUBS 0.041217f
C1044 VP.n37 VSUBS 0.043011f
C1045 VP.n38 VSUBS 0.018301f
C1046 VP.n39 VSUBS 0.022227f
C1047 VP.n40 VSUBS 0.022227f
C1048 VP.n41 VSUBS 0.022227f
C1049 VP.n42 VSUBS 0.041217f
C1050 VP.n43 VSUBS 0.041217f
C1051 VP.n44 VSUBS 1.39707f
C1052 VP.n45 VSUBS 0.022227f
C1053 VP.n46 VSUBS 0.022227f
C1054 VP.n47 VSUBS 0.022227f
C1055 VP.n48 VSUBS 0.041217f
C1056 VP.n49 VSUBS 0.044525f
C1057 VP.n50 VSUBS 0.018301f
C1058 VP.n51 VSUBS 0.022227f
C1059 VP.n52 VSUBS 0.022227f
C1060 VP.n53 VSUBS 0.022227f
C1061 VP.n54 VSUBS 0.041217f
C1062 VP.n55 VSUBS 0.041217f
C1063 VP.t4 VSUBS 3.9899f
C1064 VP.n56 VSUBS 1.3762f
C1065 VP.n57 VSUBS 0.023718f
C1066 VP.n58 VSUBS 0.022227f
C1067 VP.n59 VSUBS 0.022227f
C1068 VP.n60 VSUBS 0.022227f
C1069 VP.n61 VSUBS 0.041217f
C1070 VP.n62 VSUBS 0.044174f
C1071 VP.n63 VSUBS 0.021285f
C1072 VP.n64 VSUBS 0.022227f
C1073 VP.n65 VSUBS 0.022227f
C1074 VP.n66 VSUBS 0.022227f
C1075 VP.n67 VSUBS 0.041217f
C1076 VP.n68 VSUBS 0.041217f
C1077 VP.n69 VSUBS 0.026567f
C1078 VP.n70 VSUBS 0.035868f
C1079 VP.n71 VSUBS 1.76817f
C1080 VP.n72 VSUBS 1.78078f
C1081 VP.t9 VSUBS 3.9899f
C1082 VP.n73 VSUBS 1.46262f
C1083 VP.n74 VSUBS 0.026567f
C1084 VP.n75 VSUBS 0.035868f
C1085 VP.n76 VSUBS 0.022227f
C1086 VP.n77 VSUBS 0.022227f
C1087 VP.n78 VSUBS 0.041217f
C1088 VP.n79 VSUBS 0.040378f
C1089 VP.n80 VSUBS 0.021285f
C1090 VP.n81 VSUBS 0.022227f
C1091 VP.n82 VSUBS 0.022227f
C1092 VP.n83 VSUBS 0.022227f
C1093 VP.n84 VSUBS 0.041217f
C1094 VP.n85 VSUBS 0.038369f
C1095 VP.n86 VSUBS 1.3762f
C1096 VP.n87 VSUBS 0.023718f
C1097 VP.n88 VSUBS 0.022227f
C1098 VP.n89 VSUBS 0.022227f
C1099 VP.n90 VSUBS 0.022227f
C1100 VP.n91 VSUBS 0.041217f
C1101 VP.n92 VSUBS 0.043011f
C1102 VP.n93 VSUBS 0.018301f
C1103 VP.n94 VSUBS 0.022227f
C1104 VP.n95 VSUBS 0.022227f
C1105 VP.n96 VSUBS 0.022227f
C1106 VP.n97 VSUBS 0.041217f
C1107 VP.n98 VSUBS 0.041217f
C1108 VP.n99 VSUBS 1.39707f
C1109 VP.n100 VSUBS 0.022227f
C1110 VP.n101 VSUBS 0.022227f
C1111 VP.n102 VSUBS 0.022227f
C1112 VP.n103 VSUBS 0.041217f
C1113 VP.n104 VSUBS 0.044525f
C1114 VP.n105 VSUBS 0.018301f
C1115 VP.n106 VSUBS 0.022227f
C1116 VP.n107 VSUBS 0.022227f
C1117 VP.n108 VSUBS 0.022227f
C1118 VP.n109 VSUBS 0.041217f
C1119 VP.n110 VSUBS 0.041217f
C1120 VP.t0 VSUBS 3.9899f
C1121 VP.n111 VSUBS 1.3762f
C1122 VP.n112 VSUBS 0.023718f
C1123 VP.n113 VSUBS 0.022227f
C1124 VP.n114 VSUBS 0.022227f
C1125 VP.n115 VSUBS 0.022227f
C1126 VP.n116 VSUBS 0.041217f
C1127 VP.n117 VSUBS 0.044174f
C1128 VP.n118 VSUBS 0.021285f
C1129 VP.n119 VSUBS 0.022227f
C1130 VP.n120 VSUBS 0.022227f
C1131 VP.n121 VSUBS 0.022227f
C1132 VP.n122 VSUBS 0.041217f
C1133 VP.n123 VSUBS 0.041217f
C1134 VP.n124 VSUBS 0.026567f
C1135 VP.n125 VSUBS 0.035868f
C1136 VP.n126 VSUBS 0.064683f
C1137 B.n0 VSUBS 0.004845f
C1138 B.n1 VSUBS 0.004845f
C1139 B.n2 VSUBS 0.007662f
C1140 B.n3 VSUBS 0.007662f
C1141 B.n4 VSUBS 0.007662f
C1142 B.n5 VSUBS 0.007662f
C1143 B.n6 VSUBS 0.007662f
C1144 B.n7 VSUBS 0.007662f
C1145 B.n8 VSUBS 0.007662f
C1146 B.n9 VSUBS 0.007662f
C1147 B.n10 VSUBS 0.007662f
C1148 B.n11 VSUBS 0.007662f
C1149 B.n12 VSUBS 0.007662f
C1150 B.n13 VSUBS 0.007662f
C1151 B.n14 VSUBS 0.007662f
C1152 B.n15 VSUBS 0.007662f
C1153 B.n16 VSUBS 0.007662f
C1154 B.n17 VSUBS 0.007662f
C1155 B.n18 VSUBS 0.007662f
C1156 B.n19 VSUBS 0.007662f
C1157 B.n20 VSUBS 0.007662f
C1158 B.n21 VSUBS 0.007662f
C1159 B.n22 VSUBS 0.007662f
C1160 B.n23 VSUBS 0.007662f
C1161 B.n24 VSUBS 0.007662f
C1162 B.n25 VSUBS 0.007662f
C1163 B.n26 VSUBS 0.007662f
C1164 B.n27 VSUBS 0.007662f
C1165 B.n28 VSUBS 0.007662f
C1166 B.n29 VSUBS 0.007662f
C1167 B.n30 VSUBS 0.007662f
C1168 B.n31 VSUBS 0.007662f
C1169 B.n32 VSUBS 0.007662f
C1170 B.n33 VSUBS 0.007662f
C1171 B.n34 VSUBS 0.007662f
C1172 B.n35 VSUBS 0.007662f
C1173 B.n36 VSUBS 0.007662f
C1174 B.n37 VSUBS 0.007662f
C1175 B.n38 VSUBS 0.007662f
C1176 B.n39 VSUBS 0.007662f
C1177 B.n40 VSUBS 0.007662f
C1178 B.n41 VSUBS 0.007662f
C1179 B.n42 VSUBS 0.01789f
C1180 B.n43 VSUBS 0.007662f
C1181 B.n44 VSUBS 0.007662f
C1182 B.n45 VSUBS 0.007662f
C1183 B.n46 VSUBS 0.007662f
C1184 B.n47 VSUBS 0.007662f
C1185 B.n48 VSUBS 0.007662f
C1186 B.n49 VSUBS 0.007662f
C1187 B.n50 VSUBS 0.007662f
C1188 B.n51 VSUBS 0.007662f
C1189 B.n52 VSUBS 0.007662f
C1190 B.n53 VSUBS 0.007662f
C1191 B.n54 VSUBS 0.007662f
C1192 B.n55 VSUBS 0.007662f
C1193 B.n56 VSUBS 0.007662f
C1194 B.n57 VSUBS 0.007662f
C1195 B.n58 VSUBS 0.007662f
C1196 B.n59 VSUBS 0.007662f
C1197 B.n60 VSUBS 0.007662f
C1198 B.n61 VSUBS 0.007662f
C1199 B.n62 VSUBS 0.007662f
C1200 B.n63 VSUBS 0.007662f
C1201 B.n64 VSUBS 0.007662f
C1202 B.n65 VSUBS 0.007662f
C1203 B.n66 VSUBS 0.007662f
C1204 B.n67 VSUBS 0.007662f
C1205 B.n68 VSUBS 0.007662f
C1206 B.n69 VSUBS 0.007662f
C1207 B.n70 VSUBS 0.007662f
C1208 B.n71 VSUBS 0.007662f
C1209 B.t8 VSUBS 0.369941f
C1210 B.t7 VSUBS 0.41949f
C1211 B.t6 VSUBS 3.25976f
C1212 B.n72 VSUBS 0.669891f
C1213 B.n73 VSUBS 0.357955f
C1214 B.n74 VSUBS 0.007662f
C1215 B.n75 VSUBS 0.007662f
C1216 B.n76 VSUBS 0.007662f
C1217 B.n77 VSUBS 0.007662f
C1218 B.t11 VSUBS 0.369945f
C1219 B.t10 VSUBS 0.419493f
C1220 B.t9 VSUBS 3.25976f
C1221 B.n78 VSUBS 0.669888f
C1222 B.n79 VSUBS 0.357951f
C1223 B.n80 VSUBS 0.007662f
C1224 B.n81 VSUBS 0.007662f
C1225 B.n82 VSUBS 0.007662f
C1226 B.n83 VSUBS 0.007662f
C1227 B.n84 VSUBS 0.007662f
C1228 B.n85 VSUBS 0.007662f
C1229 B.n86 VSUBS 0.007662f
C1230 B.n87 VSUBS 0.007662f
C1231 B.n88 VSUBS 0.007662f
C1232 B.n89 VSUBS 0.007662f
C1233 B.n90 VSUBS 0.007662f
C1234 B.n91 VSUBS 0.007662f
C1235 B.n92 VSUBS 0.007662f
C1236 B.n93 VSUBS 0.007662f
C1237 B.n94 VSUBS 0.007662f
C1238 B.n95 VSUBS 0.007662f
C1239 B.n96 VSUBS 0.007662f
C1240 B.n97 VSUBS 0.007662f
C1241 B.n98 VSUBS 0.007662f
C1242 B.n99 VSUBS 0.007662f
C1243 B.n100 VSUBS 0.007662f
C1244 B.n101 VSUBS 0.007662f
C1245 B.n102 VSUBS 0.007662f
C1246 B.n103 VSUBS 0.007662f
C1247 B.n104 VSUBS 0.007662f
C1248 B.n105 VSUBS 0.007662f
C1249 B.n106 VSUBS 0.007662f
C1250 B.n107 VSUBS 0.007662f
C1251 B.n108 VSUBS 0.016948f
C1252 B.n109 VSUBS 0.007662f
C1253 B.n110 VSUBS 0.007662f
C1254 B.n111 VSUBS 0.007662f
C1255 B.n112 VSUBS 0.007662f
C1256 B.n113 VSUBS 0.007662f
C1257 B.n114 VSUBS 0.007662f
C1258 B.n115 VSUBS 0.007662f
C1259 B.n116 VSUBS 0.007662f
C1260 B.n117 VSUBS 0.007662f
C1261 B.n118 VSUBS 0.007662f
C1262 B.n119 VSUBS 0.007662f
C1263 B.n120 VSUBS 0.007662f
C1264 B.n121 VSUBS 0.007662f
C1265 B.n122 VSUBS 0.007662f
C1266 B.n123 VSUBS 0.007662f
C1267 B.n124 VSUBS 0.007662f
C1268 B.n125 VSUBS 0.007662f
C1269 B.n126 VSUBS 0.007662f
C1270 B.n127 VSUBS 0.007662f
C1271 B.n128 VSUBS 0.007662f
C1272 B.n129 VSUBS 0.007662f
C1273 B.n130 VSUBS 0.007662f
C1274 B.n131 VSUBS 0.007662f
C1275 B.n132 VSUBS 0.007662f
C1276 B.n133 VSUBS 0.007662f
C1277 B.n134 VSUBS 0.007662f
C1278 B.n135 VSUBS 0.007662f
C1279 B.n136 VSUBS 0.007662f
C1280 B.n137 VSUBS 0.007662f
C1281 B.n138 VSUBS 0.007662f
C1282 B.n139 VSUBS 0.007662f
C1283 B.n140 VSUBS 0.007662f
C1284 B.n141 VSUBS 0.007662f
C1285 B.n142 VSUBS 0.007662f
C1286 B.n143 VSUBS 0.007662f
C1287 B.n144 VSUBS 0.007662f
C1288 B.n145 VSUBS 0.007662f
C1289 B.n146 VSUBS 0.007662f
C1290 B.n147 VSUBS 0.007662f
C1291 B.n148 VSUBS 0.007662f
C1292 B.n149 VSUBS 0.007662f
C1293 B.n150 VSUBS 0.007662f
C1294 B.n151 VSUBS 0.007662f
C1295 B.n152 VSUBS 0.007662f
C1296 B.n153 VSUBS 0.007662f
C1297 B.n154 VSUBS 0.007662f
C1298 B.n155 VSUBS 0.007662f
C1299 B.n156 VSUBS 0.007662f
C1300 B.n157 VSUBS 0.007662f
C1301 B.n158 VSUBS 0.007662f
C1302 B.n159 VSUBS 0.007662f
C1303 B.n160 VSUBS 0.007662f
C1304 B.n161 VSUBS 0.007662f
C1305 B.n162 VSUBS 0.007662f
C1306 B.n163 VSUBS 0.007662f
C1307 B.n164 VSUBS 0.007662f
C1308 B.n165 VSUBS 0.007662f
C1309 B.n166 VSUBS 0.007662f
C1310 B.n167 VSUBS 0.007662f
C1311 B.n168 VSUBS 0.007662f
C1312 B.n169 VSUBS 0.007662f
C1313 B.n170 VSUBS 0.007662f
C1314 B.n171 VSUBS 0.007662f
C1315 B.n172 VSUBS 0.007662f
C1316 B.n173 VSUBS 0.007662f
C1317 B.n174 VSUBS 0.007662f
C1318 B.n175 VSUBS 0.007662f
C1319 B.n176 VSUBS 0.007662f
C1320 B.n177 VSUBS 0.007662f
C1321 B.n178 VSUBS 0.007662f
C1322 B.n179 VSUBS 0.007662f
C1323 B.n180 VSUBS 0.007662f
C1324 B.n181 VSUBS 0.007662f
C1325 B.n182 VSUBS 0.007662f
C1326 B.n183 VSUBS 0.007662f
C1327 B.n184 VSUBS 0.007662f
C1328 B.n185 VSUBS 0.007662f
C1329 B.n186 VSUBS 0.007662f
C1330 B.n187 VSUBS 0.007662f
C1331 B.n188 VSUBS 0.007662f
C1332 B.n189 VSUBS 0.01789f
C1333 B.n190 VSUBS 0.007662f
C1334 B.n191 VSUBS 0.007662f
C1335 B.n192 VSUBS 0.007662f
C1336 B.n193 VSUBS 0.007662f
C1337 B.n194 VSUBS 0.007662f
C1338 B.n195 VSUBS 0.007662f
C1339 B.n196 VSUBS 0.007662f
C1340 B.n197 VSUBS 0.007662f
C1341 B.n198 VSUBS 0.007662f
C1342 B.n199 VSUBS 0.007662f
C1343 B.n200 VSUBS 0.007662f
C1344 B.n201 VSUBS 0.007662f
C1345 B.n202 VSUBS 0.007662f
C1346 B.n203 VSUBS 0.007662f
C1347 B.n204 VSUBS 0.007662f
C1348 B.n205 VSUBS 0.007662f
C1349 B.n206 VSUBS 0.007662f
C1350 B.n207 VSUBS 0.007662f
C1351 B.n208 VSUBS 0.007662f
C1352 B.n209 VSUBS 0.007662f
C1353 B.n210 VSUBS 0.007662f
C1354 B.n211 VSUBS 0.007662f
C1355 B.n212 VSUBS 0.007662f
C1356 B.n213 VSUBS 0.007662f
C1357 B.n214 VSUBS 0.007662f
C1358 B.n215 VSUBS 0.007662f
C1359 B.n216 VSUBS 0.007662f
C1360 B.n217 VSUBS 0.007662f
C1361 B.t4 VSUBS 0.369945f
C1362 B.t5 VSUBS 0.419493f
C1363 B.t3 VSUBS 3.25976f
C1364 B.n218 VSUBS 0.669888f
C1365 B.n219 VSUBS 0.357951f
C1366 B.n220 VSUBS 0.017753f
C1367 B.n221 VSUBS 0.007662f
C1368 B.n222 VSUBS 0.007662f
C1369 B.n223 VSUBS 0.007662f
C1370 B.n224 VSUBS 0.007662f
C1371 B.n225 VSUBS 0.007662f
C1372 B.t1 VSUBS 0.369941f
C1373 B.t2 VSUBS 0.41949f
C1374 B.t0 VSUBS 3.25976f
C1375 B.n226 VSUBS 0.669891f
C1376 B.n227 VSUBS 0.357955f
C1377 B.n228 VSUBS 0.007662f
C1378 B.n229 VSUBS 0.007662f
C1379 B.n230 VSUBS 0.007662f
C1380 B.n231 VSUBS 0.007662f
C1381 B.n232 VSUBS 0.007662f
C1382 B.n233 VSUBS 0.007662f
C1383 B.n234 VSUBS 0.007662f
C1384 B.n235 VSUBS 0.007662f
C1385 B.n236 VSUBS 0.007662f
C1386 B.n237 VSUBS 0.007662f
C1387 B.n238 VSUBS 0.007662f
C1388 B.n239 VSUBS 0.007662f
C1389 B.n240 VSUBS 0.007662f
C1390 B.n241 VSUBS 0.007662f
C1391 B.n242 VSUBS 0.007662f
C1392 B.n243 VSUBS 0.007662f
C1393 B.n244 VSUBS 0.007662f
C1394 B.n245 VSUBS 0.007662f
C1395 B.n246 VSUBS 0.007662f
C1396 B.n247 VSUBS 0.007662f
C1397 B.n248 VSUBS 0.007662f
C1398 B.n249 VSUBS 0.007662f
C1399 B.n250 VSUBS 0.007662f
C1400 B.n251 VSUBS 0.007662f
C1401 B.n252 VSUBS 0.007662f
C1402 B.n253 VSUBS 0.007662f
C1403 B.n254 VSUBS 0.007662f
C1404 B.n255 VSUBS 0.007662f
C1405 B.n256 VSUBS 0.01704f
C1406 B.n257 VSUBS 0.007662f
C1407 B.n258 VSUBS 0.007662f
C1408 B.n259 VSUBS 0.007662f
C1409 B.n260 VSUBS 0.007662f
C1410 B.n261 VSUBS 0.007662f
C1411 B.n262 VSUBS 0.007662f
C1412 B.n263 VSUBS 0.007662f
C1413 B.n264 VSUBS 0.007662f
C1414 B.n265 VSUBS 0.007662f
C1415 B.n266 VSUBS 0.007662f
C1416 B.n267 VSUBS 0.007662f
C1417 B.n268 VSUBS 0.007662f
C1418 B.n269 VSUBS 0.007662f
C1419 B.n270 VSUBS 0.007662f
C1420 B.n271 VSUBS 0.007662f
C1421 B.n272 VSUBS 0.007662f
C1422 B.n273 VSUBS 0.007662f
C1423 B.n274 VSUBS 0.007662f
C1424 B.n275 VSUBS 0.007662f
C1425 B.n276 VSUBS 0.007662f
C1426 B.n277 VSUBS 0.007662f
C1427 B.n278 VSUBS 0.007662f
C1428 B.n279 VSUBS 0.007662f
C1429 B.n280 VSUBS 0.007662f
C1430 B.n281 VSUBS 0.007662f
C1431 B.n282 VSUBS 0.007662f
C1432 B.n283 VSUBS 0.007662f
C1433 B.n284 VSUBS 0.007662f
C1434 B.n285 VSUBS 0.007662f
C1435 B.n286 VSUBS 0.007662f
C1436 B.n287 VSUBS 0.007662f
C1437 B.n288 VSUBS 0.007662f
C1438 B.n289 VSUBS 0.007662f
C1439 B.n290 VSUBS 0.007662f
C1440 B.n291 VSUBS 0.007662f
C1441 B.n292 VSUBS 0.007662f
C1442 B.n293 VSUBS 0.007662f
C1443 B.n294 VSUBS 0.007662f
C1444 B.n295 VSUBS 0.007662f
C1445 B.n296 VSUBS 0.007662f
C1446 B.n297 VSUBS 0.007662f
C1447 B.n298 VSUBS 0.007662f
C1448 B.n299 VSUBS 0.007662f
C1449 B.n300 VSUBS 0.007662f
C1450 B.n301 VSUBS 0.007662f
C1451 B.n302 VSUBS 0.007662f
C1452 B.n303 VSUBS 0.007662f
C1453 B.n304 VSUBS 0.007662f
C1454 B.n305 VSUBS 0.007662f
C1455 B.n306 VSUBS 0.007662f
C1456 B.n307 VSUBS 0.007662f
C1457 B.n308 VSUBS 0.007662f
C1458 B.n309 VSUBS 0.007662f
C1459 B.n310 VSUBS 0.007662f
C1460 B.n311 VSUBS 0.007662f
C1461 B.n312 VSUBS 0.007662f
C1462 B.n313 VSUBS 0.007662f
C1463 B.n314 VSUBS 0.007662f
C1464 B.n315 VSUBS 0.007662f
C1465 B.n316 VSUBS 0.007662f
C1466 B.n317 VSUBS 0.007662f
C1467 B.n318 VSUBS 0.007662f
C1468 B.n319 VSUBS 0.007662f
C1469 B.n320 VSUBS 0.007662f
C1470 B.n321 VSUBS 0.007662f
C1471 B.n322 VSUBS 0.007662f
C1472 B.n323 VSUBS 0.007662f
C1473 B.n324 VSUBS 0.007662f
C1474 B.n325 VSUBS 0.007662f
C1475 B.n326 VSUBS 0.007662f
C1476 B.n327 VSUBS 0.007662f
C1477 B.n328 VSUBS 0.007662f
C1478 B.n329 VSUBS 0.007662f
C1479 B.n330 VSUBS 0.007662f
C1480 B.n331 VSUBS 0.007662f
C1481 B.n332 VSUBS 0.007662f
C1482 B.n333 VSUBS 0.007662f
C1483 B.n334 VSUBS 0.007662f
C1484 B.n335 VSUBS 0.007662f
C1485 B.n336 VSUBS 0.007662f
C1486 B.n337 VSUBS 0.007662f
C1487 B.n338 VSUBS 0.007662f
C1488 B.n339 VSUBS 0.007662f
C1489 B.n340 VSUBS 0.007662f
C1490 B.n341 VSUBS 0.007662f
C1491 B.n342 VSUBS 0.007662f
C1492 B.n343 VSUBS 0.007662f
C1493 B.n344 VSUBS 0.007662f
C1494 B.n345 VSUBS 0.007662f
C1495 B.n346 VSUBS 0.007662f
C1496 B.n347 VSUBS 0.007662f
C1497 B.n348 VSUBS 0.007662f
C1498 B.n349 VSUBS 0.007662f
C1499 B.n350 VSUBS 0.007662f
C1500 B.n351 VSUBS 0.007662f
C1501 B.n352 VSUBS 0.007662f
C1502 B.n353 VSUBS 0.007662f
C1503 B.n354 VSUBS 0.007662f
C1504 B.n355 VSUBS 0.007662f
C1505 B.n356 VSUBS 0.007662f
C1506 B.n357 VSUBS 0.007662f
C1507 B.n358 VSUBS 0.007662f
C1508 B.n359 VSUBS 0.007662f
C1509 B.n360 VSUBS 0.007662f
C1510 B.n361 VSUBS 0.007662f
C1511 B.n362 VSUBS 0.007662f
C1512 B.n363 VSUBS 0.007662f
C1513 B.n364 VSUBS 0.007662f
C1514 B.n365 VSUBS 0.007662f
C1515 B.n366 VSUBS 0.007662f
C1516 B.n367 VSUBS 0.007662f
C1517 B.n368 VSUBS 0.007662f
C1518 B.n369 VSUBS 0.007662f
C1519 B.n370 VSUBS 0.007662f
C1520 B.n371 VSUBS 0.007662f
C1521 B.n372 VSUBS 0.007662f
C1522 B.n373 VSUBS 0.007662f
C1523 B.n374 VSUBS 0.007662f
C1524 B.n375 VSUBS 0.007662f
C1525 B.n376 VSUBS 0.007662f
C1526 B.n377 VSUBS 0.007662f
C1527 B.n378 VSUBS 0.007662f
C1528 B.n379 VSUBS 0.007662f
C1529 B.n380 VSUBS 0.007662f
C1530 B.n381 VSUBS 0.007662f
C1531 B.n382 VSUBS 0.007662f
C1532 B.n383 VSUBS 0.007662f
C1533 B.n384 VSUBS 0.007662f
C1534 B.n385 VSUBS 0.007662f
C1535 B.n386 VSUBS 0.007662f
C1536 B.n387 VSUBS 0.007662f
C1537 B.n388 VSUBS 0.007662f
C1538 B.n389 VSUBS 0.007662f
C1539 B.n390 VSUBS 0.007662f
C1540 B.n391 VSUBS 0.007662f
C1541 B.n392 VSUBS 0.007662f
C1542 B.n393 VSUBS 0.007662f
C1543 B.n394 VSUBS 0.007662f
C1544 B.n395 VSUBS 0.007662f
C1545 B.n396 VSUBS 0.007662f
C1546 B.n397 VSUBS 0.007662f
C1547 B.n398 VSUBS 0.007662f
C1548 B.n399 VSUBS 0.007662f
C1549 B.n400 VSUBS 0.007662f
C1550 B.n401 VSUBS 0.007662f
C1551 B.n402 VSUBS 0.007662f
C1552 B.n403 VSUBS 0.007662f
C1553 B.n404 VSUBS 0.007662f
C1554 B.n405 VSUBS 0.007662f
C1555 B.n406 VSUBS 0.007662f
C1556 B.n407 VSUBS 0.007662f
C1557 B.n408 VSUBS 0.007662f
C1558 B.n409 VSUBS 0.007662f
C1559 B.n410 VSUBS 0.007662f
C1560 B.n411 VSUBS 0.007662f
C1561 B.n412 VSUBS 0.007662f
C1562 B.n413 VSUBS 0.01704f
C1563 B.n414 VSUBS 0.01789f
C1564 B.n415 VSUBS 0.01789f
C1565 B.n416 VSUBS 0.007662f
C1566 B.n417 VSUBS 0.007662f
C1567 B.n418 VSUBS 0.007662f
C1568 B.n419 VSUBS 0.007662f
C1569 B.n420 VSUBS 0.007662f
C1570 B.n421 VSUBS 0.007662f
C1571 B.n422 VSUBS 0.007662f
C1572 B.n423 VSUBS 0.007662f
C1573 B.n424 VSUBS 0.007662f
C1574 B.n425 VSUBS 0.007662f
C1575 B.n426 VSUBS 0.007662f
C1576 B.n427 VSUBS 0.007662f
C1577 B.n428 VSUBS 0.007662f
C1578 B.n429 VSUBS 0.007662f
C1579 B.n430 VSUBS 0.007662f
C1580 B.n431 VSUBS 0.007662f
C1581 B.n432 VSUBS 0.007662f
C1582 B.n433 VSUBS 0.007662f
C1583 B.n434 VSUBS 0.007662f
C1584 B.n435 VSUBS 0.007662f
C1585 B.n436 VSUBS 0.007662f
C1586 B.n437 VSUBS 0.007662f
C1587 B.n438 VSUBS 0.007662f
C1588 B.n439 VSUBS 0.007662f
C1589 B.n440 VSUBS 0.007662f
C1590 B.n441 VSUBS 0.007662f
C1591 B.n442 VSUBS 0.007662f
C1592 B.n443 VSUBS 0.007662f
C1593 B.n444 VSUBS 0.007662f
C1594 B.n445 VSUBS 0.007662f
C1595 B.n446 VSUBS 0.007662f
C1596 B.n447 VSUBS 0.007662f
C1597 B.n448 VSUBS 0.007662f
C1598 B.n449 VSUBS 0.007662f
C1599 B.n450 VSUBS 0.007662f
C1600 B.n451 VSUBS 0.007662f
C1601 B.n452 VSUBS 0.007662f
C1602 B.n453 VSUBS 0.007662f
C1603 B.n454 VSUBS 0.007662f
C1604 B.n455 VSUBS 0.007662f
C1605 B.n456 VSUBS 0.007662f
C1606 B.n457 VSUBS 0.007662f
C1607 B.n458 VSUBS 0.007662f
C1608 B.n459 VSUBS 0.007662f
C1609 B.n460 VSUBS 0.007662f
C1610 B.n461 VSUBS 0.007662f
C1611 B.n462 VSUBS 0.007662f
C1612 B.n463 VSUBS 0.007662f
C1613 B.n464 VSUBS 0.007662f
C1614 B.n465 VSUBS 0.007662f
C1615 B.n466 VSUBS 0.007662f
C1616 B.n467 VSUBS 0.007662f
C1617 B.n468 VSUBS 0.007662f
C1618 B.n469 VSUBS 0.007662f
C1619 B.n470 VSUBS 0.007662f
C1620 B.n471 VSUBS 0.007662f
C1621 B.n472 VSUBS 0.007662f
C1622 B.n473 VSUBS 0.007662f
C1623 B.n474 VSUBS 0.007662f
C1624 B.n475 VSUBS 0.007662f
C1625 B.n476 VSUBS 0.007662f
C1626 B.n477 VSUBS 0.007662f
C1627 B.n478 VSUBS 0.007662f
C1628 B.n479 VSUBS 0.007662f
C1629 B.n480 VSUBS 0.007662f
C1630 B.n481 VSUBS 0.007662f
C1631 B.n482 VSUBS 0.007662f
C1632 B.n483 VSUBS 0.007662f
C1633 B.n484 VSUBS 0.007662f
C1634 B.n485 VSUBS 0.007662f
C1635 B.n486 VSUBS 0.007662f
C1636 B.n487 VSUBS 0.007662f
C1637 B.n488 VSUBS 0.007662f
C1638 B.n489 VSUBS 0.007662f
C1639 B.n490 VSUBS 0.007662f
C1640 B.n491 VSUBS 0.007662f
C1641 B.n492 VSUBS 0.007662f
C1642 B.n493 VSUBS 0.007662f
C1643 B.n494 VSUBS 0.007662f
C1644 B.n495 VSUBS 0.007662f
C1645 B.n496 VSUBS 0.007662f
C1646 B.n497 VSUBS 0.007662f
C1647 B.n498 VSUBS 0.007662f
C1648 B.n499 VSUBS 0.007662f
C1649 B.n500 VSUBS 0.005296f
C1650 B.n501 VSUBS 0.017753f
C1651 B.n502 VSUBS 0.006197f
C1652 B.n503 VSUBS 0.007662f
C1653 B.n504 VSUBS 0.007662f
C1654 B.n505 VSUBS 0.007662f
C1655 B.n506 VSUBS 0.007662f
C1656 B.n507 VSUBS 0.007662f
C1657 B.n508 VSUBS 0.007662f
C1658 B.n509 VSUBS 0.007662f
C1659 B.n510 VSUBS 0.007662f
C1660 B.n511 VSUBS 0.007662f
C1661 B.n512 VSUBS 0.007662f
C1662 B.n513 VSUBS 0.007662f
C1663 B.n514 VSUBS 0.006197f
C1664 B.n515 VSUBS 0.007662f
C1665 B.n516 VSUBS 0.007662f
C1666 B.n517 VSUBS 0.005296f
C1667 B.n518 VSUBS 0.007662f
C1668 B.n519 VSUBS 0.007662f
C1669 B.n520 VSUBS 0.007662f
C1670 B.n521 VSUBS 0.007662f
C1671 B.n522 VSUBS 0.007662f
C1672 B.n523 VSUBS 0.007662f
C1673 B.n524 VSUBS 0.007662f
C1674 B.n525 VSUBS 0.007662f
C1675 B.n526 VSUBS 0.007662f
C1676 B.n527 VSUBS 0.007662f
C1677 B.n528 VSUBS 0.007662f
C1678 B.n529 VSUBS 0.007662f
C1679 B.n530 VSUBS 0.007662f
C1680 B.n531 VSUBS 0.007662f
C1681 B.n532 VSUBS 0.007662f
C1682 B.n533 VSUBS 0.007662f
C1683 B.n534 VSUBS 0.007662f
C1684 B.n535 VSUBS 0.007662f
C1685 B.n536 VSUBS 0.007662f
C1686 B.n537 VSUBS 0.007662f
C1687 B.n538 VSUBS 0.007662f
C1688 B.n539 VSUBS 0.007662f
C1689 B.n540 VSUBS 0.007662f
C1690 B.n541 VSUBS 0.007662f
C1691 B.n542 VSUBS 0.007662f
C1692 B.n543 VSUBS 0.007662f
C1693 B.n544 VSUBS 0.007662f
C1694 B.n545 VSUBS 0.007662f
C1695 B.n546 VSUBS 0.007662f
C1696 B.n547 VSUBS 0.007662f
C1697 B.n548 VSUBS 0.007662f
C1698 B.n549 VSUBS 0.007662f
C1699 B.n550 VSUBS 0.007662f
C1700 B.n551 VSUBS 0.007662f
C1701 B.n552 VSUBS 0.007662f
C1702 B.n553 VSUBS 0.007662f
C1703 B.n554 VSUBS 0.007662f
C1704 B.n555 VSUBS 0.007662f
C1705 B.n556 VSUBS 0.007662f
C1706 B.n557 VSUBS 0.007662f
C1707 B.n558 VSUBS 0.007662f
C1708 B.n559 VSUBS 0.007662f
C1709 B.n560 VSUBS 0.007662f
C1710 B.n561 VSUBS 0.007662f
C1711 B.n562 VSUBS 0.007662f
C1712 B.n563 VSUBS 0.007662f
C1713 B.n564 VSUBS 0.007662f
C1714 B.n565 VSUBS 0.007662f
C1715 B.n566 VSUBS 0.007662f
C1716 B.n567 VSUBS 0.007662f
C1717 B.n568 VSUBS 0.007662f
C1718 B.n569 VSUBS 0.007662f
C1719 B.n570 VSUBS 0.007662f
C1720 B.n571 VSUBS 0.007662f
C1721 B.n572 VSUBS 0.007662f
C1722 B.n573 VSUBS 0.007662f
C1723 B.n574 VSUBS 0.007662f
C1724 B.n575 VSUBS 0.007662f
C1725 B.n576 VSUBS 0.007662f
C1726 B.n577 VSUBS 0.007662f
C1727 B.n578 VSUBS 0.007662f
C1728 B.n579 VSUBS 0.007662f
C1729 B.n580 VSUBS 0.007662f
C1730 B.n581 VSUBS 0.007662f
C1731 B.n582 VSUBS 0.007662f
C1732 B.n583 VSUBS 0.007662f
C1733 B.n584 VSUBS 0.007662f
C1734 B.n585 VSUBS 0.007662f
C1735 B.n586 VSUBS 0.007662f
C1736 B.n587 VSUBS 0.007662f
C1737 B.n588 VSUBS 0.007662f
C1738 B.n589 VSUBS 0.007662f
C1739 B.n590 VSUBS 0.007662f
C1740 B.n591 VSUBS 0.007662f
C1741 B.n592 VSUBS 0.007662f
C1742 B.n593 VSUBS 0.007662f
C1743 B.n594 VSUBS 0.007662f
C1744 B.n595 VSUBS 0.007662f
C1745 B.n596 VSUBS 0.007662f
C1746 B.n597 VSUBS 0.007662f
C1747 B.n598 VSUBS 0.007662f
C1748 B.n599 VSUBS 0.007662f
C1749 B.n600 VSUBS 0.007662f
C1750 B.n601 VSUBS 0.007662f
C1751 B.n602 VSUBS 0.01789f
C1752 B.n603 VSUBS 0.01704f
C1753 B.n604 VSUBS 0.01704f
C1754 B.n605 VSUBS 0.007662f
C1755 B.n606 VSUBS 0.007662f
C1756 B.n607 VSUBS 0.007662f
C1757 B.n608 VSUBS 0.007662f
C1758 B.n609 VSUBS 0.007662f
C1759 B.n610 VSUBS 0.007662f
C1760 B.n611 VSUBS 0.007662f
C1761 B.n612 VSUBS 0.007662f
C1762 B.n613 VSUBS 0.007662f
C1763 B.n614 VSUBS 0.007662f
C1764 B.n615 VSUBS 0.007662f
C1765 B.n616 VSUBS 0.007662f
C1766 B.n617 VSUBS 0.007662f
C1767 B.n618 VSUBS 0.007662f
C1768 B.n619 VSUBS 0.007662f
C1769 B.n620 VSUBS 0.007662f
C1770 B.n621 VSUBS 0.007662f
C1771 B.n622 VSUBS 0.007662f
C1772 B.n623 VSUBS 0.007662f
C1773 B.n624 VSUBS 0.007662f
C1774 B.n625 VSUBS 0.007662f
C1775 B.n626 VSUBS 0.007662f
C1776 B.n627 VSUBS 0.007662f
C1777 B.n628 VSUBS 0.007662f
C1778 B.n629 VSUBS 0.007662f
C1779 B.n630 VSUBS 0.007662f
C1780 B.n631 VSUBS 0.007662f
C1781 B.n632 VSUBS 0.007662f
C1782 B.n633 VSUBS 0.007662f
C1783 B.n634 VSUBS 0.007662f
C1784 B.n635 VSUBS 0.007662f
C1785 B.n636 VSUBS 0.007662f
C1786 B.n637 VSUBS 0.007662f
C1787 B.n638 VSUBS 0.007662f
C1788 B.n639 VSUBS 0.007662f
C1789 B.n640 VSUBS 0.007662f
C1790 B.n641 VSUBS 0.007662f
C1791 B.n642 VSUBS 0.007662f
C1792 B.n643 VSUBS 0.007662f
C1793 B.n644 VSUBS 0.007662f
C1794 B.n645 VSUBS 0.007662f
C1795 B.n646 VSUBS 0.007662f
C1796 B.n647 VSUBS 0.007662f
C1797 B.n648 VSUBS 0.007662f
C1798 B.n649 VSUBS 0.007662f
C1799 B.n650 VSUBS 0.007662f
C1800 B.n651 VSUBS 0.007662f
C1801 B.n652 VSUBS 0.007662f
C1802 B.n653 VSUBS 0.007662f
C1803 B.n654 VSUBS 0.007662f
C1804 B.n655 VSUBS 0.007662f
C1805 B.n656 VSUBS 0.007662f
C1806 B.n657 VSUBS 0.007662f
C1807 B.n658 VSUBS 0.007662f
C1808 B.n659 VSUBS 0.007662f
C1809 B.n660 VSUBS 0.007662f
C1810 B.n661 VSUBS 0.007662f
C1811 B.n662 VSUBS 0.007662f
C1812 B.n663 VSUBS 0.007662f
C1813 B.n664 VSUBS 0.007662f
C1814 B.n665 VSUBS 0.007662f
C1815 B.n666 VSUBS 0.007662f
C1816 B.n667 VSUBS 0.007662f
C1817 B.n668 VSUBS 0.007662f
C1818 B.n669 VSUBS 0.007662f
C1819 B.n670 VSUBS 0.007662f
C1820 B.n671 VSUBS 0.007662f
C1821 B.n672 VSUBS 0.007662f
C1822 B.n673 VSUBS 0.007662f
C1823 B.n674 VSUBS 0.007662f
C1824 B.n675 VSUBS 0.007662f
C1825 B.n676 VSUBS 0.007662f
C1826 B.n677 VSUBS 0.007662f
C1827 B.n678 VSUBS 0.007662f
C1828 B.n679 VSUBS 0.007662f
C1829 B.n680 VSUBS 0.007662f
C1830 B.n681 VSUBS 0.007662f
C1831 B.n682 VSUBS 0.007662f
C1832 B.n683 VSUBS 0.007662f
C1833 B.n684 VSUBS 0.007662f
C1834 B.n685 VSUBS 0.007662f
C1835 B.n686 VSUBS 0.007662f
C1836 B.n687 VSUBS 0.007662f
C1837 B.n688 VSUBS 0.007662f
C1838 B.n689 VSUBS 0.007662f
C1839 B.n690 VSUBS 0.007662f
C1840 B.n691 VSUBS 0.007662f
C1841 B.n692 VSUBS 0.007662f
C1842 B.n693 VSUBS 0.007662f
C1843 B.n694 VSUBS 0.007662f
C1844 B.n695 VSUBS 0.007662f
C1845 B.n696 VSUBS 0.007662f
C1846 B.n697 VSUBS 0.007662f
C1847 B.n698 VSUBS 0.007662f
C1848 B.n699 VSUBS 0.007662f
C1849 B.n700 VSUBS 0.007662f
C1850 B.n701 VSUBS 0.007662f
C1851 B.n702 VSUBS 0.007662f
C1852 B.n703 VSUBS 0.007662f
C1853 B.n704 VSUBS 0.007662f
C1854 B.n705 VSUBS 0.007662f
C1855 B.n706 VSUBS 0.007662f
C1856 B.n707 VSUBS 0.007662f
C1857 B.n708 VSUBS 0.007662f
C1858 B.n709 VSUBS 0.007662f
C1859 B.n710 VSUBS 0.007662f
C1860 B.n711 VSUBS 0.007662f
C1861 B.n712 VSUBS 0.007662f
C1862 B.n713 VSUBS 0.007662f
C1863 B.n714 VSUBS 0.007662f
C1864 B.n715 VSUBS 0.007662f
C1865 B.n716 VSUBS 0.007662f
C1866 B.n717 VSUBS 0.007662f
C1867 B.n718 VSUBS 0.007662f
C1868 B.n719 VSUBS 0.007662f
C1869 B.n720 VSUBS 0.007662f
C1870 B.n721 VSUBS 0.007662f
C1871 B.n722 VSUBS 0.007662f
C1872 B.n723 VSUBS 0.007662f
C1873 B.n724 VSUBS 0.007662f
C1874 B.n725 VSUBS 0.007662f
C1875 B.n726 VSUBS 0.007662f
C1876 B.n727 VSUBS 0.007662f
C1877 B.n728 VSUBS 0.007662f
C1878 B.n729 VSUBS 0.007662f
C1879 B.n730 VSUBS 0.007662f
C1880 B.n731 VSUBS 0.007662f
C1881 B.n732 VSUBS 0.007662f
C1882 B.n733 VSUBS 0.007662f
C1883 B.n734 VSUBS 0.007662f
C1884 B.n735 VSUBS 0.007662f
C1885 B.n736 VSUBS 0.007662f
C1886 B.n737 VSUBS 0.007662f
C1887 B.n738 VSUBS 0.007662f
C1888 B.n739 VSUBS 0.007662f
C1889 B.n740 VSUBS 0.007662f
C1890 B.n741 VSUBS 0.007662f
C1891 B.n742 VSUBS 0.007662f
C1892 B.n743 VSUBS 0.007662f
C1893 B.n744 VSUBS 0.007662f
C1894 B.n745 VSUBS 0.007662f
C1895 B.n746 VSUBS 0.007662f
C1896 B.n747 VSUBS 0.007662f
C1897 B.n748 VSUBS 0.007662f
C1898 B.n749 VSUBS 0.007662f
C1899 B.n750 VSUBS 0.007662f
C1900 B.n751 VSUBS 0.007662f
C1901 B.n752 VSUBS 0.007662f
C1902 B.n753 VSUBS 0.007662f
C1903 B.n754 VSUBS 0.007662f
C1904 B.n755 VSUBS 0.007662f
C1905 B.n756 VSUBS 0.007662f
C1906 B.n757 VSUBS 0.007662f
C1907 B.n758 VSUBS 0.007662f
C1908 B.n759 VSUBS 0.007662f
C1909 B.n760 VSUBS 0.007662f
C1910 B.n761 VSUBS 0.007662f
C1911 B.n762 VSUBS 0.007662f
C1912 B.n763 VSUBS 0.007662f
C1913 B.n764 VSUBS 0.007662f
C1914 B.n765 VSUBS 0.007662f
C1915 B.n766 VSUBS 0.007662f
C1916 B.n767 VSUBS 0.007662f
C1917 B.n768 VSUBS 0.007662f
C1918 B.n769 VSUBS 0.007662f
C1919 B.n770 VSUBS 0.007662f
C1920 B.n771 VSUBS 0.007662f
C1921 B.n772 VSUBS 0.007662f
C1922 B.n773 VSUBS 0.007662f
C1923 B.n774 VSUBS 0.007662f
C1924 B.n775 VSUBS 0.007662f
C1925 B.n776 VSUBS 0.007662f
C1926 B.n777 VSUBS 0.007662f
C1927 B.n778 VSUBS 0.007662f
C1928 B.n779 VSUBS 0.007662f
C1929 B.n780 VSUBS 0.007662f
C1930 B.n781 VSUBS 0.007662f
C1931 B.n782 VSUBS 0.007662f
C1932 B.n783 VSUBS 0.007662f
C1933 B.n784 VSUBS 0.007662f
C1934 B.n785 VSUBS 0.007662f
C1935 B.n786 VSUBS 0.007662f
C1936 B.n787 VSUBS 0.007662f
C1937 B.n788 VSUBS 0.007662f
C1938 B.n789 VSUBS 0.007662f
C1939 B.n790 VSUBS 0.007662f
C1940 B.n791 VSUBS 0.007662f
C1941 B.n792 VSUBS 0.007662f
C1942 B.n793 VSUBS 0.007662f
C1943 B.n794 VSUBS 0.007662f
C1944 B.n795 VSUBS 0.007662f
C1945 B.n796 VSUBS 0.007662f
C1946 B.n797 VSUBS 0.007662f
C1947 B.n798 VSUBS 0.007662f
C1948 B.n799 VSUBS 0.007662f
C1949 B.n800 VSUBS 0.007662f
C1950 B.n801 VSUBS 0.007662f
C1951 B.n802 VSUBS 0.007662f
C1952 B.n803 VSUBS 0.007662f
C1953 B.n804 VSUBS 0.007662f
C1954 B.n805 VSUBS 0.007662f
C1955 B.n806 VSUBS 0.007662f
C1956 B.n807 VSUBS 0.007662f
C1957 B.n808 VSUBS 0.007662f
C1958 B.n809 VSUBS 0.007662f
C1959 B.n810 VSUBS 0.007662f
C1960 B.n811 VSUBS 0.007662f
C1961 B.n812 VSUBS 0.007662f
C1962 B.n813 VSUBS 0.007662f
C1963 B.n814 VSUBS 0.007662f
C1964 B.n815 VSUBS 0.007662f
C1965 B.n816 VSUBS 0.007662f
C1966 B.n817 VSUBS 0.007662f
C1967 B.n818 VSUBS 0.007662f
C1968 B.n819 VSUBS 0.007662f
C1969 B.n820 VSUBS 0.007662f
C1970 B.n821 VSUBS 0.007662f
C1971 B.n822 VSUBS 0.007662f
C1972 B.n823 VSUBS 0.007662f
C1973 B.n824 VSUBS 0.007662f
C1974 B.n825 VSUBS 0.007662f
C1975 B.n826 VSUBS 0.007662f
C1976 B.n827 VSUBS 0.007662f
C1977 B.n828 VSUBS 0.007662f
C1978 B.n829 VSUBS 0.007662f
C1979 B.n830 VSUBS 0.007662f
C1980 B.n831 VSUBS 0.007662f
C1981 B.n832 VSUBS 0.007662f
C1982 B.n833 VSUBS 0.007662f
C1983 B.n834 VSUBS 0.007662f
C1984 B.n835 VSUBS 0.007662f
C1985 B.n836 VSUBS 0.007662f
C1986 B.n837 VSUBS 0.007662f
C1987 B.n838 VSUBS 0.007662f
C1988 B.n839 VSUBS 0.007662f
C1989 B.n840 VSUBS 0.007662f
C1990 B.n841 VSUBS 0.007662f
C1991 B.n842 VSUBS 0.007662f
C1992 B.n843 VSUBS 0.017982f
C1993 B.n844 VSUBS 0.01704f
C1994 B.n845 VSUBS 0.01789f
C1995 B.n846 VSUBS 0.007662f
C1996 B.n847 VSUBS 0.007662f
C1997 B.n848 VSUBS 0.007662f
C1998 B.n849 VSUBS 0.007662f
C1999 B.n850 VSUBS 0.007662f
C2000 B.n851 VSUBS 0.007662f
C2001 B.n852 VSUBS 0.007662f
C2002 B.n853 VSUBS 0.007662f
C2003 B.n854 VSUBS 0.007662f
C2004 B.n855 VSUBS 0.007662f
C2005 B.n856 VSUBS 0.007662f
C2006 B.n857 VSUBS 0.007662f
C2007 B.n858 VSUBS 0.007662f
C2008 B.n859 VSUBS 0.007662f
C2009 B.n860 VSUBS 0.007662f
C2010 B.n861 VSUBS 0.007662f
C2011 B.n862 VSUBS 0.007662f
C2012 B.n863 VSUBS 0.007662f
C2013 B.n864 VSUBS 0.007662f
C2014 B.n865 VSUBS 0.007662f
C2015 B.n866 VSUBS 0.007662f
C2016 B.n867 VSUBS 0.007662f
C2017 B.n868 VSUBS 0.007662f
C2018 B.n869 VSUBS 0.007662f
C2019 B.n870 VSUBS 0.007662f
C2020 B.n871 VSUBS 0.007662f
C2021 B.n872 VSUBS 0.007662f
C2022 B.n873 VSUBS 0.007662f
C2023 B.n874 VSUBS 0.007662f
C2024 B.n875 VSUBS 0.007662f
C2025 B.n876 VSUBS 0.007662f
C2026 B.n877 VSUBS 0.007662f
C2027 B.n878 VSUBS 0.007662f
C2028 B.n879 VSUBS 0.007662f
C2029 B.n880 VSUBS 0.007662f
C2030 B.n881 VSUBS 0.007662f
C2031 B.n882 VSUBS 0.007662f
C2032 B.n883 VSUBS 0.007662f
C2033 B.n884 VSUBS 0.007662f
C2034 B.n885 VSUBS 0.007662f
C2035 B.n886 VSUBS 0.007662f
C2036 B.n887 VSUBS 0.007662f
C2037 B.n888 VSUBS 0.007662f
C2038 B.n889 VSUBS 0.007662f
C2039 B.n890 VSUBS 0.007662f
C2040 B.n891 VSUBS 0.007662f
C2041 B.n892 VSUBS 0.007662f
C2042 B.n893 VSUBS 0.007662f
C2043 B.n894 VSUBS 0.007662f
C2044 B.n895 VSUBS 0.007662f
C2045 B.n896 VSUBS 0.007662f
C2046 B.n897 VSUBS 0.007662f
C2047 B.n898 VSUBS 0.007662f
C2048 B.n899 VSUBS 0.007662f
C2049 B.n900 VSUBS 0.007662f
C2050 B.n901 VSUBS 0.007662f
C2051 B.n902 VSUBS 0.007662f
C2052 B.n903 VSUBS 0.007662f
C2053 B.n904 VSUBS 0.007662f
C2054 B.n905 VSUBS 0.007662f
C2055 B.n906 VSUBS 0.007662f
C2056 B.n907 VSUBS 0.007662f
C2057 B.n908 VSUBS 0.007662f
C2058 B.n909 VSUBS 0.007662f
C2059 B.n910 VSUBS 0.007662f
C2060 B.n911 VSUBS 0.007662f
C2061 B.n912 VSUBS 0.007662f
C2062 B.n913 VSUBS 0.007662f
C2063 B.n914 VSUBS 0.007662f
C2064 B.n915 VSUBS 0.007662f
C2065 B.n916 VSUBS 0.007662f
C2066 B.n917 VSUBS 0.007662f
C2067 B.n918 VSUBS 0.007662f
C2068 B.n919 VSUBS 0.007662f
C2069 B.n920 VSUBS 0.007662f
C2070 B.n921 VSUBS 0.007662f
C2071 B.n922 VSUBS 0.007662f
C2072 B.n923 VSUBS 0.007662f
C2073 B.n924 VSUBS 0.007662f
C2074 B.n925 VSUBS 0.007662f
C2075 B.n926 VSUBS 0.007662f
C2076 B.n927 VSUBS 0.007662f
C2077 B.n928 VSUBS 0.007662f
C2078 B.n929 VSUBS 0.007662f
C2079 B.n930 VSUBS 0.007662f
C2080 B.n931 VSUBS 0.005296f
C2081 B.n932 VSUBS 0.017753f
C2082 B.n933 VSUBS 0.006197f
C2083 B.n934 VSUBS 0.007662f
C2084 B.n935 VSUBS 0.007662f
C2085 B.n936 VSUBS 0.007662f
C2086 B.n937 VSUBS 0.007662f
C2087 B.n938 VSUBS 0.007662f
C2088 B.n939 VSUBS 0.007662f
C2089 B.n940 VSUBS 0.007662f
C2090 B.n941 VSUBS 0.007662f
C2091 B.n942 VSUBS 0.007662f
C2092 B.n943 VSUBS 0.007662f
C2093 B.n944 VSUBS 0.007662f
C2094 B.n945 VSUBS 0.006197f
C2095 B.n946 VSUBS 0.017753f
C2096 B.n947 VSUBS 0.005296f
C2097 B.n948 VSUBS 0.007662f
C2098 B.n949 VSUBS 0.007662f
C2099 B.n950 VSUBS 0.007662f
C2100 B.n951 VSUBS 0.007662f
C2101 B.n952 VSUBS 0.007662f
C2102 B.n953 VSUBS 0.007662f
C2103 B.n954 VSUBS 0.007662f
C2104 B.n955 VSUBS 0.007662f
C2105 B.n956 VSUBS 0.007662f
C2106 B.n957 VSUBS 0.007662f
C2107 B.n958 VSUBS 0.007662f
C2108 B.n959 VSUBS 0.007662f
C2109 B.n960 VSUBS 0.007662f
C2110 B.n961 VSUBS 0.007662f
C2111 B.n962 VSUBS 0.007662f
C2112 B.n963 VSUBS 0.007662f
C2113 B.n964 VSUBS 0.007662f
C2114 B.n965 VSUBS 0.007662f
C2115 B.n966 VSUBS 0.007662f
C2116 B.n967 VSUBS 0.007662f
C2117 B.n968 VSUBS 0.007662f
C2118 B.n969 VSUBS 0.007662f
C2119 B.n970 VSUBS 0.007662f
C2120 B.n971 VSUBS 0.007662f
C2121 B.n972 VSUBS 0.007662f
C2122 B.n973 VSUBS 0.007662f
C2123 B.n974 VSUBS 0.007662f
C2124 B.n975 VSUBS 0.007662f
C2125 B.n976 VSUBS 0.007662f
C2126 B.n977 VSUBS 0.007662f
C2127 B.n978 VSUBS 0.007662f
C2128 B.n979 VSUBS 0.007662f
C2129 B.n980 VSUBS 0.007662f
C2130 B.n981 VSUBS 0.007662f
C2131 B.n982 VSUBS 0.007662f
C2132 B.n983 VSUBS 0.007662f
C2133 B.n984 VSUBS 0.007662f
C2134 B.n985 VSUBS 0.007662f
C2135 B.n986 VSUBS 0.007662f
C2136 B.n987 VSUBS 0.007662f
C2137 B.n988 VSUBS 0.007662f
C2138 B.n989 VSUBS 0.007662f
C2139 B.n990 VSUBS 0.007662f
C2140 B.n991 VSUBS 0.007662f
C2141 B.n992 VSUBS 0.007662f
C2142 B.n993 VSUBS 0.007662f
C2143 B.n994 VSUBS 0.007662f
C2144 B.n995 VSUBS 0.007662f
C2145 B.n996 VSUBS 0.007662f
C2146 B.n997 VSUBS 0.007662f
C2147 B.n998 VSUBS 0.007662f
C2148 B.n999 VSUBS 0.007662f
C2149 B.n1000 VSUBS 0.007662f
C2150 B.n1001 VSUBS 0.007662f
C2151 B.n1002 VSUBS 0.007662f
C2152 B.n1003 VSUBS 0.007662f
C2153 B.n1004 VSUBS 0.007662f
C2154 B.n1005 VSUBS 0.007662f
C2155 B.n1006 VSUBS 0.007662f
C2156 B.n1007 VSUBS 0.007662f
C2157 B.n1008 VSUBS 0.007662f
C2158 B.n1009 VSUBS 0.007662f
C2159 B.n1010 VSUBS 0.007662f
C2160 B.n1011 VSUBS 0.007662f
C2161 B.n1012 VSUBS 0.007662f
C2162 B.n1013 VSUBS 0.007662f
C2163 B.n1014 VSUBS 0.007662f
C2164 B.n1015 VSUBS 0.007662f
C2165 B.n1016 VSUBS 0.007662f
C2166 B.n1017 VSUBS 0.007662f
C2167 B.n1018 VSUBS 0.007662f
C2168 B.n1019 VSUBS 0.007662f
C2169 B.n1020 VSUBS 0.007662f
C2170 B.n1021 VSUBS 0.007662f
C2171 B.n1022 VSUBS 0.007662f
C2172 B.n1023 VSUBS 0.007662f
C2173 B.n1024 VSUBS 0.007662f
C2174 B.n1025 VSUBS 0.007662f
C2175 B.n1026 VSUBS 0.007662f
C2176 B.n1027 VSUBS 0.007662f
C2177 B.n1028 VSUBS 0.007662f
C2178 B.n1029 VSUBS 0.007662f
C2179 B.n1030 VSUBS 0.007662f
C2180 B.n1031 VSUBS 0.007662f
C2181 B.n1032 VSUBS 0.007662f
C2182 B.n1033 VSUBS 0.01789f
C2183 B.n1034 VSUBS 0.01704f
C2184 B.n1035 VSUBS 0.01704f
C2185 B.n1036 VSUBS 0.007662f
C2186 B.n1037 VSUBS 0.007662f
C2187 B.n1038 VSUBS 0.007662f
C2188 B.n1039 VSUBS 0.007662f
C2189 B.n1040 VSUBS 0.007662f
C2190 B.n1041 VSUBS 0.007662f
C2191 B.n1042 VSUBS 0.007662f
C2192 B.n1043 VSUBS 0.007662f
C2193 B.n1044 VSUBS 0.007662f
C2194 B.n1045 VSUBS 0.007662f
C2195 B.n1046 VSUBS 0.007662f
C2196 B.n1047 VSUBS 0.007662f
C2197 B.n1048 VSUBS 0.007662f
C2198 B.n1049 VSUBS 0.007662f
C2199 B.n1050 VSUBS 0.007662f
C2200 B.n1051 VSUBS 0.007662f
C2201 B.n1052 VSUBS 0.007662f
C2202 B.n1053 VSUBS 0.007662f
C2203 B.n1054 VSUBS 0.007662f
C2204 B.n1055 VSUBS 0.007662f
C2205 B.n1056 VSUBS 0.007662f
C2206 B.n1057 VSUBS 0.007662f
C2207 B.n1058 VSUBS 0.007662f
C2208 B.n1059 VSUBS 0.007662f
C2209 B.n1060 VSUBS 0.007662f
C2210 B.n1061 VSUBS 0.007662f
C2211 B.n1062 VSUBS 0.007662f
C2212 B.n1063 VSUBS 0.007662f
C2213 B.n1064 VSUBS 0.007662f
C2214 B.n1065 VSUBS 0.007662f
C2215 B.n1066 VSUBS 0.007662f
C2216 B.n1067 VSUBS 0.007662f
C2217 B.n1068 VSUBS 0.007662f
C2218 B.n1069 VSUBS 0.007662f
C2219 B.n1070 VSUBS 0.007662f
C2220 B.n1071 VSUBS 0.007662f
C2221 B.n1072 VSUBS 0.007662f
C2222 B.n1073 VSUBS 0.007662f
C2223 B.n1074 VSUBS 0.007662f
C2224 B.n1075 VSUBS 0.007662f
C2225 B.n1076 VSUBS 0.007662f
C2226 B.n1077 VSUBS 0.007662f
C2227 B.n1078 VSUBS 0.007662f
C2228 B.n1079 VSUBS 0.007662f
C2229 B.n1080 VSUBS 0.007662f
C2230 B.n1081 VSUBS 0.007662f
C2231 B.n1082 VSUBS 0.007662f
C2232 B.n1083 VSUBS 0.007662f
C2233 B.n1084 VSUBS 0.007662f
C2234 B.n1085 VSUBS 0.007662f
C2235 B.n1086 VSUBS 0.007662f
C2236 B.n1087 VSUBS 0.007662f
C2237 B.n1088 VSUBS 0.007662f
C2238 B.n1089 VSUBS 0.007662f
C2239 B.n1090 VSUBS 0.007662f
C2240 B.n1091 VSUBS 0.007662f
C2241 B.n1092 VSUBS 0.007662f
C2242 B.n1093 VSUBS 0.007662f
C2243 B.n1094 VSUBS 0.007662f
C2244 B.n1095 VSUBS 0.007662f
C2245 B.n1096 VSUBS 0.007662f
C2246 B.n1097 VSUBS 0.007662f
C2247 B.n1098 VSUBS 0.007662f
C2248 B.n1099 VSUBS 0.007662f
C2249 B.n1100 VSUBS 0.007662f
C2250 B.n1101 VSUBS 0.007662f
C2251 B.n1102 VSUBS 0.007662f
C2252 B.n1103 VSUBS 0.007662f
C2253 B.n1104 VSUBS 0.007662f
C2254 B.n1105 VSUBS 0.007662f
C2255 B.n1106 VSUBS 0.007662f
C2256 B.n1107 VSUBS 0.007662f
C2257 B.n1108 VSUBS 0.007662f
C2258 B.n1109 VSUBS 0.007662f
C2259 B.n1110 VSUBS 0.007662f
C2260 B.n1111 VSUBS 0.007662f
C2261 B.n1112 VSUBS 0.007662f
C2262 B.n1113 VSUBS 0.007662f
C2263 B.n1114 VSUBS 0.007662f
C2264 B.n1115 VSUBS 0.007662f
C2265 B.n1116 VSUBS 0.007662f
C2266 B.n1117 VSUBS 0.007662f
C2267 B.n1118 VSUBS 0.007662f
C2268 B.n1119 VSUBS 0.007662f
C2269 B.n1120 VSUBS 0.007662f
C2270 B.n1121 VSUBS 0.007662f
C2271 B.n1122 VSUBS 0.007662f
C2272 B.n1123 VSUBS 0.007662f
C2273 B.n1124 VSUBS 0.007662f
C2274 B.n1125 VSUBS 0.007662f
C2275 B.n1126 VSUBS 0.007662f
C2276 B.n1127 VSUBS 0.007662f
C2277 B.n1128 VSUBS 0.007662f
C2278 B.n1129 VSUBS 0.007662f
C2279 B.n1130 VSUBS 0.007662f
C2280 B.n1131 VSUBS 0.007662f
C2281 B.n1132 VSUBS 0.007662f
C2282 B.n1133 VSUBS 0.007662f
C2283 B.n1134 VSUBS 0.007662f
C2284 B.n1135 VSUBS 0.007662f
C2285 B.n1136 VSUBS 0.007662f
C2286 B.n1137 VSUBS 0.007662f
C2287 B.n1138 VSUBS 0.007662f
C2288 B.n1139 VSUBS 0.007662f
C2289 B.n1140 VSUBS 0.007662f
C2290 B.n1141 VSUBS 0.007662f
C2291 B.n1142 VSUBS 0.007662f
C2292 B.n1143 VSUBS 0.007662f
C2293 B.n1144 VSUBS 0.007662f
C2294 B.n1145 VSUBS 0.007662f
C2295 B.n1146 VSUBS 0.007662f
C2296 B.n1147 VSUBS 0.007662f
C2297 B.n1148 VSUBS 0.007662f
C2298 B.n1149 VSUBS 0.007662f
C2299 B.n1150 VSUBS 0.007662f
C2300 B.n1151 VSUBS 0.007662f
C2301 B.n1152 VSUBS 0.007662f
C2302 B.n1153 VSUBS 0.007662f
C2303 B.n1154 VSUBS 0.007662f
C2304 B.n1155 VSUBS 0.01735f
.ends

