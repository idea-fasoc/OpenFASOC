* NGSPICE file created from diff_pair_sample_1560.ext - technology: sky130A

.subckt diff_pair_sample_1560 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X1 VTAIL.t11 VP.t1 VDD1.t8 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X2 VTAIL.t4 VN.t0 VDD2.t9 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X3 VDD1.t7 VP.t2 VTAIL.t15 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=1.2
X4 VDD2.t8 VN.t1 VTAIL.t7 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=1.2
X5 VDD2.t7 VN.t2 VTAIL.t0 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X6 VTAIL.t5 VN.t3 VDD2.t6 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X7 B.t11 B.t9 B.t10 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=1.2
X8 VDD2.t5 VN.t4 VTAIL.t1 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=1.2
X9 VDD1.t6 VP.t3 VTAIL.t16 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=1.2
X10 VDD1.t5 VP.t4 VTAIL.t12 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=1.2
X11 VDD2.t4 VN.t5 VTAIL.t6 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=1.2
X12 VTAIL.t2 VN.t6 VDD2.t3 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X13 VDD1.t4 VP.t5 VTAIL.t17 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=1.2
X14 VDD2.t2 VN.t7 VTAIL.t8 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X15 B.t8 B.t6 B.t7 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=1.2
X16 VTAIL.t13 VP.t6 VDD1.t3 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X17 VTAIL.t14 VP.t7 VDD1.t2 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X18 VDD1.t1 VP.t8 VTAIL.t18 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X19 VTAIL.t19 VP.t9 VDD1.t0 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X20 VDD2.t1 VN.t8 VTAIL.t3 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=1.2
X21 B.t5 B.t3 B.t4 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=1.2
X22 VTAIL.t9 VN.t9 VDD2.t0 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=1.2
X23 B.t2 B.t0 B.t1 w_n2806_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=1.2
R0 VP.n15 VP.n14 161.3
R1 VP.n16 VP.n11 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n20 VP.n19 161.3
R4 VP.n21 VP.n9 161.3
R5 VP.n23 VP.n22 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n26 VP.n7 161.3
R8 VP.n46 VP.n0 161.3
R9 VP.n45 VP.n44 161.3
R10 VP.n43 VP.n42 161.3
R11 VP.n41 VP.n2 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n38 VP.n37 161.3
R14 VP.n36 VP.n4 161.3
R15 VP.n35 VP.n34 161.3
R16 VP.n33 VP.n32 161.3
R17 VP.n31 VP.n6 161.3
R18 VP.n13 VP.t5 102.323
R19 VP.n30 VP.t4 83.3463
R20 VP.n47 VP.t2 83.3463
R21 VP.n27 VP.t3 83.3463
R22 VP.n28 VP.n27 80.6037
R23 VP.n48 VP.n47 80.6037
R24 VP.n30 VP.n29 80.6037
R25 VP.n5 VP.t6 50.4097
R26 VP.n3 VP.t8 50.4097
R27 VP.n1 VP.t7 50.4097
R28 VP.n8 VP.t1 50.4097
R29 VP.n10 VP.t0 50.4097
R30 VP.n12 VP.t9 50.4097
R31 VP.n13 VP.n12 43.9705
R32 VP.n36 VP.n35 41.9503
R33 VP.n42 VP.n41 41.9503
R34 VP.n22 VP.n21 41.9503
R35 VP.n16 VP.n15 41.9503
R36 VP.n37 VP.n36 39.0365
R37 VP.n41 VP.n40 39.0365
R38 VP.n21 VP.n20 39.0365
R39 VP.n17 VP.n16 39.0365
R40 VP.n29 VP.n28 38.437
R41 VP.n32 VP.n31 36.1227
R42 VP.n46 VP.n45 36.1227
R43 VP.n26 VP.n25 36.1227
R44 VP.n31 VP.n30 30.6732
R45 VP.n47 VP.n46 30.6732
R46 VP.n27 VP.n26 30.6732
R47 VP.n14 VP.n13 29.5703
R48 VP.n35 VP.n5 13.702
R49 VP.n42 VP.n1 13.702
R50 VP.n22 VP.n8 13.702
R51 VP.n15 VP.n12 13.702
R52 VP.n37 VP.n3 12.234
R53 VP.n40 VP.n3 12.234
R54 VP.n17 VP.n10 12.234
R55 VP.n20 VP.n10 12.234
R56 VP.n32 VP.n5 10.766
R57 VP.n45 VP.n1 10.766
R58 VP.n25 VP.n8 10.766
R59 VP.n28 VP.n7 0.285035
R60 VP.n29 VP.n6 0.285035
R61 VP.n48 VP.n0 0.285035
R62 VP.n14 VP.n11 0.189894
R63 VP.n18 VP.n11 0.189894
R64 VP.n19 VP.n18 0.189894
R65 VP.n19 VP.n9 0.189894
R66 VP.n23 VP.n9 0.189894
R67 VP.n24 VP.n23 0.189894
R68 VP.n24 VP.n7 0.189894
R69 VP.n33 VP.n6 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n4 0.189894
R72 VP.n38 VP.n4 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n43 VP.n2 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n44 VP.n0 0.189894
R78 VP VP.n48 0.146778
R79 VTAIL.n56 VTAIL.n50 756.745
R80 VTAIL.n8 VTAIL.n2 756.745
R81 VTAIL.n44 VTAIL.n38 756.745
R82 VTAIL.n28 VTAIL.n22 756.745
R83 VTAIL.n55 VTAIL.n54 585
R84 VTAIL.n57 VTAIL.n56 585
R85 VTAIL.n7 VTAIL.n6 585
R86 VTAIL.n9 VTAIL.n8 585
R87 VTAIL.n45 VTAIL.n44 585
R88 VTAIL.n43 VTAIL.n42 585
R89 VTAIL.n29 VTAIL.n28 585
R90 VTAIL.n27 VTAIL.n26 585
R91 VTAIL.n53 VTAIL.t3 355.474
R92 VTAIL.n5 VTAIL.t15 355.474
R93 VTAIL.n41 VTAIL.t16 355.474
R94 VTAIL.n25 VTAIL.t1 355.474
R95 VTAIL.n56 VTAIL.n55 171.744
R96 VTAIL.n8 VTAIL.n7 171.744
R97 VTAIL.n44 VTAIL.n43 171.744
R98 VTAIL.n28 VTAIL.n27 171.744
R99 VTAIL.n37 VTAIL.n36 137.174
R100 VTAIL.n35 VTAIL.n34 137.174
R101 VTAIL.n21 VTAIL.n20 137.174
R102 VTAIL.n19 VTAIL.n18 137.174
R103 VTAIL.n63 VTAIL.n62 137.174
R104 VTAIL.n1 VTAIL.n0 137.174
R105 VTAIL.n15 VTAIL.n14 137.174
R106 VTAIL.n17 VTAIL.n16 137.174
R107 VTAIL.n55 VTAIL.t3 85.8723
R108 VTAIL.n7 VTAIL.t15 85.8723
R109 VTAIL.n43 VTAIL.t16 85.8723
R110 VTAIL.n27 VTAIL.t1 85.8723
R111 VTAIL.n61 VTAIL.n60 34.3187
R112 VTAIL.n13 VTAIL.n12 34.3187
R113 VTAIL.n49 VTAIL.n48 34.3187
R114 VTAIL.n33 VTAIL.n32 34.3187
R115 VTAIL.n19 VTAIL.n17 17.1686
R116 VTAIL.n61 VTAIL.n49 15.8496
R117 VTAIL.n54 VTAIL.n53 15.8418
R118 VTAIL.n6 VTAIL.n5 15.8418
R119 VTAIL.n42 VTAIL.n41 15.8418
R120 VTAIL.n26 VTAIL.n25 15.8418
R121 VTAIL.n62 VTAIL.t0 12.9507
R122 VTAIL.n62 VTAIL.t4 12.9507
R123 VTAIL.n0 VTAIL.t6 12.9507
R124 VTAIL.n0 VTAIL.t5 12.9507
R125 VTAIL.n14 VTAIL.t18 12.9507
R126 VTAIL.n14 VTAIL.t14 12.9507
R127 VTAIL.n16 VTAIL.t12 12.9507
R128 VTAIL.n16 VTAIL.t13 12.9507
R129 VTAIL.n36 VTAIL.t10 12.9507
R130 VTAIL.n36 VTAIL.t11 12.9507
R131 VTAIL.n34 VTAIL.t17 12.9507
R132 VTAIL.n34 VTAIL.t19 12.9507
R133 VTAIL.n20 VTAIL.t8 12.9507
R134 VTAIL.n20 VTAIL.t2 12.9507
R135 VTAIL.n18 VTAIL.t7 12.9507
R136 VTAIL.n18 VTAIL.t9 12.9507
R137 VTAIL.n57 VTAIL.n52 12.8005
R138 VTAIL.n9 VTAIL.n4 12.8005
R139 VTAIL.n45 VTAIL.n40 12.8005
R140 VTAIL.n29 VTAIL.n24 12.8005
R141 VTAIL.n58 VTAIL.n50 12.0247
R142 VTAIL.n10 VTAIL.n2 12.0247
R143 VTAIL.n46 VTAIL.n38 12.0247
R144 VTAIL.n30 VTAIL.n22 12.0247
R145 VTAIL.n60 VTAIL.n59 9.45567
R146 VTAIL.n12 VTAIL.n11 9.45567
R147 VTAIL.n48 VTAIL.n47 9.45567
R148 VTAIL.n32 VTAIL.n31 9.45567
R149 VTAIL.n59 VTAIL.n58 9.3005
R150 VTAIL.n52 VTAIL.n51 9.3005
R151 VTAIL.n11 VTAIL.n10 9.3005
R152 VTAIL.n4 VTAIL.n3 9.3005
R153 VTAIL.n47 VTAIL.n46 9.3005
R154 VTAIL.n40 VTAIL.n39 9.3005
R155 VTAIL.n31 VTAIL.n30 9.3005
R156 VTAIL.n24 VTAIL.n23 9.3005
R157 VTAIL.n41 VTAIL.n39 4.29255
R158 VTAIL.n25 VTAIL.n23 4.29255
R159 VTAIL.n53 VTAIL.n51 4.29255
R160 VTAIL.n5 VTAIL.n3 4.29255
R161 VTAIL.n60 VTAIL.n50 1.93989
R162 VTAIL.n12 VTAIL.n2 1.93989
R163 VTAIL.n48 VTAIL.n38 1.93989
R164 VTAIL.n32 VTAIL.n22 1.93989
R165 VTAIL.n21 VTAIL.n19 1.31947
R166 VTAIL.n33 VTAIL.n21 1.31947
R167 VTAIL.n37 VTAIL.n35 1.31947
R168 VTAIL.n49 VTAIL.n37 1.31947
R169 VTAIL.n17 VTAIL.n15 1.31947
R170 VTAIL.n15 VTAIL.n13 1.31947
R171 VTAIL.n63 VTAIL.n61 1.31947
R172 VTAIL.n58 VTAIL.n57 1.16414
R173 VTAIL.n10 VTAIL.n9 1.16414
R174 VTAIL.n46 VTAIL.n45 1.16414
R175 VTAIL.n30 VTAIL.n29 1.16414
R176 VTAIL.n35 VTAIL.n33 1.12981
R177 VTAIL.n13 VTAIL.n1 1.12981
R178 VTAIL VTAIL.n1 1.04791
R179 VTAIL.n54 VTAIL.n52 0.388379
R180 VTAIL.n6 VTAIL.n4 0.388379
R181 VTAIL.n42 VTAIL.n40 0.388379
R182 VTAIL.n26 VTAIL.n24 0.388379
R183 VTAIL VTAIL.n63 0.272052
R184 VTAIL.n59 VTAIL.n51 0.155672
R185 VTAIL.n11 VTAIL.n3 0.155672
R186 VTAIL.n47 VTAIL.n39 0.155672
R187 VTAIL.n31 VTAIL.n23 0.155672
R188 VDD1.n6 VDD1.n0 756.745
R189 VDD1.n19 VDD1.n13 756.745
R190 VDD1.n7 VDD1.n6 585
R191 VDD1.n5 VDD1.n4 585
R192 VDD1.n18 VDD1.n17 585
R193 VDD1.n20 VDD1.n19 585
R194 VDD1.n3 VDD1.t4 355.474
R195 VDD1.n16 VDD1.t5 355.474
R196 VDD1.n6 VDD1.n5 171.744
R197 VDD1.n19 VDD1.n18 171.744
R198 VDD1.n27 VDD1.n26 154.787
R199 VDD1.n12 VDD1.n11 153.853
R200 VDD1.n29 VDD1.n28 153.853
R201 VDD1.n25 VDD1.n24 153.853
R202 VDD1.n5 VDD1.t4 85.8723
R203 VDD1.n18 VDD1.t5 85.8723
R204 VDD1.n12 VDD1.n10 52.3164
R205 VDD1.n25 VDD1.n23 52.3164
R206 VDD1.n29 VDD1.n27 33.3867
R207 VDD1.n4 VDD1.n3 15.8418
R208 VDD1.n17 VDD1.n16 15.8418
R209 VDD1.n28 VDD1.t8 12.9507
R210 VDD1.n28 VDD1.t6 12.9507
R211 VDD1.n11 VDD1.t0 12.9507
R212 VDD1.n11 VDD1.t9 12.9507
R213 VDD1.n26 VDD1.t2 12.9507
R214 VDD1.n26 VDD1.t7 12.9507
R215 VDD1.n24 VDD1.t3 12.9507
R216 VDD1.n24 VDD1.t1 12.9507
R217 VDD1.n7 VDD1.n2 12.8005
R218 VDD1.n20 VDD1.n15 12.8005
R219 VDD1.n8 VDD1.n0 12.0247
R220 VDD1.n21 VDD1.n13 12.0247
R221 VDD1.n10 VDD1.n9 9.45567
R222 VDD1.n23 VDD1.n22 9.45567
R223 VDD1.n9 VDD1.n8 9.3005
R224 VDD1.n2 VDD1.n1 9.3005
R225 VDD1.n22 VDD1.n21 9.3005
R226 VDD1.n15 VDD1.n14 9.3005
R227 VDD1.n3 VDD1.n1 4.29255
R228 VDD1.n16 VDD1.n14 4.29255
R229 VDD1.n10 VDD1.n0 1.93989
R230 VDD1.n23 VDD1.n13 1.93989
R231 VDD1.n8 VDD1.n7 1.16414
R232 VDD1.n21 VDD1.n20 1.16414
R233 VDD1 VDD1.n29 0.931535
R234 VDD1 VDD1.n12 0.388431
R235 VDD1.n4 VDD1.n2 0.388379
R236 VDD1.n17 VDD1.n15 0.388379
R237 VDD1.n27 VDD1.n25 0.274895
R238 VDD1.n9 VDD1.n1 0.155672
R239 VDD1.n22 VDD1.n14 0.155672
R240 VN.n41 VN.n22 161.3
R241 VN.n40 VN.n39 161.3
R242 VN.n38 VN.n37 161.3
R243 VN.n36 VN.n24 161.3
R244 VN.n35 VN.n34 161.3
R245 VN.n33 VN.n32 161.3
R246 VN.n31 VN.n26 161.3
R247 VN.n30 VN.n29 161.3
R248 VN.n19 VN.n0 161.3
R249 VN.n18 VN.n17 161.3
R250 VN.n16 VN.n15 161.3
R251 VN.n14 VN.n2 161.3
R252 VN.n13 VN.n12 161.3
R253 VN.n11 VN.n10 161.3
R254 VN.n9 VN.n4 161.3
R255 VN.n8 VN.n7 161.3
R256 VN.n6 VN.t5 102.323
R257 VN.n28 VN.t4 102.323
R258 VN.n20 VN.t8 83.3463
R259 VN.n42 VN.t1 83.3463
R260 VN.n43 VN.n42 80.6037
R261 VN.n21 VN.n20 80.6037
R262 VN.n5 VN.t3 50.4097
R263 VN.n3 VN.t2 50.4097
R264 VN.n1 VN.t0 50.4097
R265 VN.n27 VN.t6 50.4097
R266 VN.n25 VN.t7 50.4097
R267 VN.n23 VN.t9 50.4097
R268 VN.n6 VN.n5 43.9705
R269 VN.n28 VN.n27 43.9705
R270 VN.n9 VN.n8 41.9503
R271 VN.n15 VN.n14 41.9503
R272 VN.n31 VN.n30 41.9503
R273 VN.n37 VN.n36 41.9503
R274 VN.n10 VN.n9 39.0365
R275 VN.n14 VN.n13 39.0365
R276 VN.n32 VN.n31 39.0365
R277 VN.n36 VN.n35 39.0365
R278 VN VN.n43 38.7225
R279 VN.n19 VN.n18 36.1227
R280 VN.n41 VN.n40 36.1227
R281 VN.n20 VN.n19 30.6732
R282 VN.n42 VN.n41 30.6732
R283 VN.n29 VN.n28 29.5703
R284 VN.n7 VN.n6 29.5703
R285 VN.n8 VN.n5 13.702
R286 VN.n15 VN.n1 13.702
R287 VN.n30 VN.n27 13.702
R288 VN.n37 VN.n23 13.702
R289 VN.n10 VN.n3 12.234
R290 VN.n13 VN.n3 12.234
R291 VN.n35 VN.n25 12.234
R292 VN.n32 VN.n25 12.234
R293 VN.n18 VN.n1 10.766
R294 VN.n40 VN.n23 10.766
R295 VN.n43 VN.n22 0.285035
R296 VN.n21 VN.n0 0.285035
R297 VN.n39 VN.n22 0.189894
R298 VN.n39 VN.n38 0.189894
R299 VN.n38 VN.n24 0.189894
R300 VN.n34 VN.n24 0.189894
R301 VN.n34 VN.n33 0.189894
R302 VN.n33 VN.n26 0.189894
R303 VN.n29 VN.n26 0.189894
R304 VN.n7 VN.n4 0.189894
R305 VN.n11 VN.n4 0.189894
R306 VN.n12 VN.n11 0.189894
R307 VN.n12 VN.n2 0.189894
R308 VN.n16 VN.n2 0.189894
R309 VN.n17 VN.n16 0.189894
R310 VN.n17 VN.n0 0.189894
R311 VN VN.n21 0.146778
R312 VDD2.n21 VDD2.n15 756.745
R313 VDD2.n6 VDD2.n0 756.745
R314 VDD2.n22 VDD2.n21 585
R315 VDD2.n20 VDD2.n19 585
R316 VDD2.n5 VDD2.n4 585
R317 VDD2.n7 VDD2.n6 585
R318 VDD2.n18 VDD2.t8 355.474
R319 VDD2.n3 VDD2.t4 355.474
R320 VDD2.n21 VDD2.n20 171.744
R321 VDD2.n6 VDD2.n5 171.744
R322 VDD2.n14 VDD2.n13 154.787
R323 VDD2 VDD2.n29 154.785
R324 VDD2.n28 VDD2.n27 153.853
R325 VDD2.n12 VDD2.n11 153.853
R326 VDD2.n20 VDD2.t8 85.8723
R327 VDD2.n5 VDD2.t4 85.8723
R328 VDD2.n12 VDD2.n10 52.3164
R329 VDD2.n26 VDD2.n25 50.9975
R330 VDD2.n26 VDD2.n14 32.1442
R331 VDD2.n19 VDD2.n18 15.8418
R332 VDD2.n4 VDD2.n3 15.8418
R333 VDD2.n29 VDD2.t3 12.9507
R334 VDD2.n29 VDD2.t5 12.9507
R335 VDD2.n27 VDD2.t0 12.9507
R336 VDD2.n27 VDD2.t2 12.9507
R337 VDD2.n13 VDD2.t9 12.9507
R338 VDD2.n13 VDD2.t1 12.9507
R339 VDD2.n11 VDD2.t6 12.9507
R340 VDD2.n11 VDD2.t7 12.9507
R341 VDD2.n22 VDD2.n17 12.8005
R342 VDD2.n7 VDD2.n2 12.8005
R343 VDD2.n23 VDD2.n15 12.0247
R344 VDD2.n8 VDD2.n0 12.0247
R345 VDD2.n25 VDD2.n24 9.45567
R346 VDD2.n10 VDD2.n9 9.45567
R347 VDD2.n24 VDD2.n23 9.3005
R348 VDD2.n17 VDD2.n16 9.3005
R349 VDD2.n9 VDD2.n8 9.3005
R350 VDD2.n2 VDD2.n1 9.3005
R351 VDD2.n18 VDD2.n16 4.29255
R352 VDD2.n3 VDD2.n1 4.29255
R353 VDD2.n25 VDD2.n15 1.93989
R354 VDD2.n10 VDD2.n0 1.93989
R355 VDD2.n28 VDD2.n26 1.31947
R356 VDD2.n23 VDD2.n22 1.16414
R357 VDD2.n8 VDD2.n7 1.16414
R358 VDD2 VDD2.n28 0.388431
R359 VDD2.n19 VDD2.n17 0.388379
R360 VDD2.n4 VDD2.n2 0.388379
R361 VDD2.n14 VDD2.n12 0.274895
R362 VDD2.n24 VDD2.n16 0.155672
R363 VDD2.n9 VDD2.n1 0.155672
R364 B.n334 B.n333 585
R365 B.n335 B.n42 585
R366 B.n337 B.n336 585
R367 B.n338 B.n41 585
R368 B.n340 B.n339 585
R369 B.n341 B.n40 585
R370 B.n343 B.n342 585
R371 B.n344 B.n39 585
R372 B.n346 B.n345 585
R373 B.n347 B.n38 585
R374 B.n349 B.n348 585
R375 B.n350 B.n37 585
R376 B.n352 B.n351 585
R377 B.n353 B.n34 585
R378 B.n356 B.n355 585
R379 B.n357 B.n33 585
R380 B.n359 B.n358 585
R381 B.n360 B.n32 585
R382 B.n362 B.n361 585
R383 B.n363 B.n31 585
R384 B.n365 B.n364 585
R385 B.n366 B.n27 585
R386 B.n368 B.n367 585
R387 B.n369 B.n26 585
R388 B.n371 B.n370 585
R389 B.n372 B.n25 585
R390 B.n374 B.n373 585
R391 B.n375 B.n24 585
R392 B.n377 B.n376 585
R393 B.n378 B.n23 585
R394 B.n380 B.n379 585
R395 B.n381 B.n22 585
R396 B.n383 B.n382 585
R397 B.n384 B.n21 585
R398 B.n386 B.n385 585
R399 B.n387 B.n20 585
R400 B.n389 B.n388 585
R401 B.n332 B.n43 585
R402 B.n331 B.n330 585
R403 B.n329 B.n44 585
R404 B.n328 B.n327 585
R405 B.n326 B.n45 585
R406 B.n325 B.n324 585
R407 B.n323 B.n46 585
R408 B.n322 B.n321 585
R409 B.n320 B.n47 585
R410 B.n319 B.n318 585
R411 B.n317 B.n48 585
R412 B.n316 B.n315 585
R413 B.n314 B.n49 585
R414 B.n313 B.n312 585
R415 B.n311 B.n50 585
R416 B.n310 B.n309 585
R417 B.n308 B.n51 585
R418 B.n307 B.n306 585
R419 B.n305 B.n52 585
R420 B.n304 B.n303 585
R421 B.n302 B.n53 585
R422 B.n301 B.n300 585
R423 B.n299 B.n54 585
R424 B.n298 B.n297 585
R425 B.n296 B.n55 585
R426 B.n295 B.n294 585
R427 B.n293 B.n56 585
R428 B.n292 B.n291 585
R429 B.n290 B.n57 585
R430 B.n289 B.n288 585
R431 B.n287 B.n58 585
R432 B.n286 B.n285 585
R433 B.n284 B.n59 585
R434 B.n283 B.n282 585
R435 B.n281 B.n60 585
R436 B.n280 B.n279 585
R437 B.n278 B.n61 585
R438 B.n277 B.n276 585
R439 B.n275 B.n62 585
R440 B.n274 B.n273 585
R441 B.n272 B.n63 585
R442 B.n271 B.n270 585
R443 B.n269 B.n64 585
R444 B.n268 B.n267 585
R445 B.n266 B.n65 585
R446 B.n265 B.n264 585
R447 B.n263 B.n66 585
R448 B.n262 B.n261 585
R449 B.n260 B.n67 585
R450 B.n259 B.n258 585
R451 B.n257 B.n68 585
R452 B.n256 B.n255 585
R453 B.n254 B.n69 585
R454 B.n253 B.n252 585
R455 B.n251 B.n70 585
R456 B.n250 B.n249 585
R457 B.n248 B.n71 585
R458 B.n247 B.n246 585
R459 B.n245 B.n72 585
R460 B.n244 B.n243 585
R461 B.n242 B.n73 585
R462 B.n241 B.n240 585
R463 B.n239 B.n74 585
R464 B.n238 B.n237 585
R465 B.n236 B.n75 585
R466 B.n235 B.n234 585
R467 B.n233 B.n76 585
R468 B.n232 B.n231 585
R469 B.n230 B.n77 585
R470 B.n229 B.n228 585
R471 B.n227 B.n78 585
R472 B.n168 B.n167 585
R473 B.n169 B.n98 585
R474 B.n171 B.n170 585
R475 B.n172 B.n97 585
R476 B.n174 B.n173 585
R477 B.n175 B.n96 585
R478 B.n177 B.n176 585
R479 B.n178 B.n95 585
R480 B.n180 B.n179 585
R481 B.n181 B.n94 585
R482 B.n183 B.n182 585
R483 B.n184 B.n93 585
R484 B.n186 B.n185 585
R485 B.n187 B.n90 585
R486 B.n190 B.n189 585
R487 B.n191 B.n89 585
R488 B.n193 B.n192 585
R489 B.n194 B.n88 585
R490 B.n196 B.n195 585
R491 B.n197 B.n87 585
R492 B.n199 B.n198 585
R493 B.n200 B.n86 585
R494 B.n205 B.n204 585
R495 B.n206 B.n85 585
R496 B.n208 B.n207 585
R497 B.n209 B.n84 585
R498 B.n211 B.n210 585
R499 B.n212 B.n83 585
R500 B.n214 B.n213 585
R501 B.n215 B.n82 585
R502 B.n217 B.n216 585
R503 B.n218 B.n81 585
R504 B.n220 B.n219 585
R505 B.n221 B.n80 585
R506 B.n223 B.n222 585
R507 B.n224 B.n79 585
R508 B.n226 B.n225 585
R509 B.n166 B.n99 585
R510 B.n165 B.n164 585
R511 B.n163 B.n100 585
R512 B.n162 B.n161 585
R513 B.n160 B.n101 585
R514 B.n159 B.n158 585
R515 B.n157 B.n102 585
R516 B.n156 B.n155 585
R517 B.n154 B.n103 585
R518 B.n153 B.n152 585
R519 B.n151 B.n104 585
R520 B.n150 B.n149 585
R521 B.n148 B.n105 585
R522 B.n147 B.n146 585
R523 B.n145 B.n106 585
R524 B.n144 B.n143 585
R525 B.n142 B.n107 585
R526 B.n141 B.n140 585
R527 B.n139 B.n108 585
R528 B.n138 B.n137 585
R529 B.n136 B.n109 585
R530 B.n135 B.n134 585
R531 B.n133 B.n110 585
R532 B.n132 B.n131 585
R533 B.n130 B.n111 585
R534 B.n129 B.n128 585
R535 B.n127 B.n112 585
R536 B.n126 B.n125 585
R537 B.n124 B.n113 585
R538 B.n123 B.n122 585
R539 B.n121 B.n114 585
R540 B.n120 B.n119 585
R541 B.n118 B.n115 585
R542 B.n117 B.n116 585
R543 B.n2 B.n0 585
R544 B.n441 B.n1 585
R545 B.n440 B.n439 585
R546 B.n438 B.n3 585
R547 B.n437 B.n436 585
R548 B.n435 B.n4 585
R549 B.n434 B.n433 585
R550 B.n432 B.n5 585
R551 B.n431 B.n430 585
R552 B.n429 B.n6 585
R553 B.n428 B.n427 585
R554 B.n426 B.n7 585
R555 B.n425 B.n424 585
R556 B.n423 B.n8 585
R557 B.n422 B.n421 585
R558 B.n420 B.n9 585
R559 B.n419 B.n418 585
R560 B.n417 B.n10 585
R561 B.n416 B.n415 585
R562 B.n414 B.n11 585
R563 B.n413 B.n412 585
R564 B.n411 B.n12 585
R565 B.n410 B.n409 585
R566 B.n408 B.n13 585
R567 B.n407 B.n406 585
R568 B.n405 B.n14 585
R569 B.n404 B.n403 585
R570 B.n402 B.n15 585
R571 B.n401 B.n400 585
R572 B.n399 B.n16 585
R573 B.n398 B.n397 585
R574 B.n396 B.n17 585
R575 B.n395 B.n394 585
R576 B.n393 B.n18 585
R577 B.n392 B.n391 585
R578 B.n390 B.n19 585
R579 B.n443 B.n442 585
R580 B.n167 B.n166 516.524
R581 B.n388 B.n19 516.524
R582 B.n225 B.n78 516.524
R583 B.n333 B.n332 516.524
R584 B.n201 B.t0 254.525
R585 B.n91 B.t6 254.525
R586 B.n28 B.t3 254.525
R587 B.n35 B.t9 254.525
R588 B.n201 B.t2 254.119
R589 B.n35 B.t10 254.119
R590 B.n91 B.t8 254.118
R591 B.n28 B.t4 254.118
R592 B.n202 B.t1 224.446
R593 B.n36 B.t11 224.446
R594 B.n92 B.t7 224.446
R595 B.n29 B.t5 224.446
R596 B.n166 B.n165 163.367
R597 B.n165 B.n100 163.367
R598 B.n161 B.n100 163.367
R599 B.n161 B.n160 163.367
R600 B.n160 B.n159 163.367
R601 B.n159 B.n102 163.367
R602 B.n155 B.n102 163.367
R603 B.n155 B.n154 163.367
R604 B.n154 B.n153 163.367
R605 B.n153 B.n104 163.367
R606 B.n149 B.n104 163.367
R607 B.n149 B.n148 163.367
R608 B.n148 B.n147 163.367
R609 B.n147 B.n106 163.367
R610 B.n143 B.n106 163.367
R611 B.n143 B.n142 163.367
R612 B.n142 B.n141 163.367
R613 B.n141 B.n108 163.367
R614 B.n137 B.n108 163.367
R615 B.n137 B.n136 163.367
R616 B.n136 B.n135 163.367
R617 B.n135 B.n110 163.367
R618 B.n131 B.n110 163.367
R619 B.n131 B.n130 163.367
R620 B.n130 B.n129 163.367
R621 B.n129 B.n112 163.367
R622 B.n125 B.n112 163.367
R623 B.n125 B.n124 163.367
R624 B.n124 B.n123 163.367
R625 B.n123 B.n114 163.367
R626 B.n119 B.n114 163.367
R627 B.n119 B.n118 163.367
R628 B.n118 B.n117 163.367
R629 B.n117 B.n2 163.367
R630 B.n442 B.n2 163.367
R631 B.n442 B.n441 163.367
R632 B.n441 B.n440 163.367
R633 B.n440 B.n3 163.367
R634 B.n436 B.n3 163.367
R635 B.n436 B.n435 163.367
R636 B.n435 B.n434 163.367
R637 B.n434 B.n5 163.367
R638 B.n430 B.n5 163.367
R639 B.n430 B.n429 163.367
R640 B.n429 B.n428 163.367
R641 B.n428 B.n7 163.367
R642 B.n424 B.n7 163.367
R643 B.n424 B.n423 163.367
R644 B.n423 B.n422 163.367
R645 B.n422 B.n9 163.367
R646 B.n418 B.n9 163.367
R647 B.n418 B.n417 163.367
R648 B.n417 B.n416 163.367
R649 B.n416 B.n11 163.367
R650 B.n412 B.n11 163.367
R651 B.n412 B.n411 163.367
R652 B.n411 B.n410 163.367
R653 B.n410 B.n13 163.367
R654 B.n406 B.n13 163.367
R655 B.n406 B.n405 163.367
R656 B.n405 B.n404 163.367
R657 B.n404 B.n15 163.367
R658 B.n400 B.n15 163.367
R659 B.n400 B.n399 163.367
R660 B.n399 B.n398 163.367
R661 B.n398 B.n17 163.367
R662 B.n394 B.n17 163.367
R663 B.n394 B.n393 163.367
R664 B.n393 B.n392 163.367
R665 B.n392 B.n19 163.367
R666 B.n167 B.n98 163.367
R667 B.n171 B.n98 163.367
R668 B.n172 B.n171 163.367
R669 B.n173 B.n172 163.367
R670 B.n173 B.n96 163.367
R671 B.n177 B.n96 163.367
R672 B.n178 B.n177 163.367
R673 B.n179 B.n178 163.367
R674 B.n179 B.n94 163.367
R675 B.n183 B.n94 163.367
R676 B.n184 B.n183 163.367
R677 B.n185 B.n184 163.367
R678 B.n185 B.n90 163.367
R679 B.n190 B.n90 163.367
R680 B.n191 B.n190 163.367
R681 B.n192 B.n191 163.367
R682 B.n192 B.n88 163.367
R683 B.n196 B.n88 163.367
R684 B.n197 B.n196 163.367
R685 B.n198 B.n197 163.367
R686 B.n198 B.n86 163.367
R687 B.n205 B.n86 163.367
R688 B.n206 B.n205 163.367
R689 B.n207 B.n206 163.367
R690 B.n207 B.n84 163.367
R691 B.n211 B.n84 163.367
R692 B.n212 B.n211 163.367
R693 B.n213 B.n212 163.367
R694 B.n213 B.n82 163.367
R695 B.n217 B.n82 163.367
R696 B.n218 B.n217 163.367
R697 B.n219 B.n218 163.367
R698 B.n219 B.n80 163.367
R699 B.n223 B.n80 163.367
R700 B.n224 B.n223 163.367
R701 B.n225 B.n224 163.367
R702 B.n229 B.n78 163.367
R703 B.n230 B.n229 163.367
R704 B.n231 B.n230 163.367
R705 B.n231 B.n76 163.367
R706 B.n235 B.n76 163.367
R707 B.n236 B.n235 163.367
R708 B.n237 B.n236 163.367
R709 B.n237 B.n74 163.367
R710 B.n241 B.n74 163.367
R711 B.n242 B.n241 163.367
R712 B.n243 B.n242 163.367
R713 B.n243 B.n72 163.367
R714 B.n247 B.n72 163.367
R715 B.n248 B.n247 163.367
R716 B.n249 B.n248 163.367
R717 B.n249 B.n70 163.367
R718 B.n253 B.n70 163.367
R719 B.n254 B.n253 163.367
R720 B.n255 B.n254 163.367
R721 B.n255 B.n68 163.367
R722 B.n259 B.n68 163.367
R723 B.n260 B.n259 163.367
R724 B.n261 B.n260 163.367
R725 B.n261 B.n66 163.367
R726 B.n265 B.n66 163.367
R727 B.n266 B.n265 163.367
R728 B.n267 B.n266 163.367
R729 B.n267 B.n64 163.367
R730 B.n271 B.n64 163.367
R731 B.n272 B.n271 163.367
R732 B.n273 B.n272 163.367
R733 B.n273 B.n62 163.367
R734 B.n277 B.n62 163.367
R735 B.n278 B.n277 163.367
R736 B.n279 B.n278 163.367
R737 B.n279 B.n60 163.367
R738 B.n283 B.n60 163.367
R739 B.n284 B.n283 163.367
R740 B.n285 B.n284 163.367
R741 B.n285 B.n58 163.367
R742 B.n289 B.n58 163.367
R743 B.n290 B.n289 163.367
R744 B.n291 B.n290 163.367
R745 B.n291 B.n56 163.367
R746 B.n295 B.n56 163.367
R747 B.n296 B.n295 163.367
R748 B.n297 B.n296 163.367
R749 B.n297 B.n54 163.367
R750 B.n301 B.n54 163.367
R751 B.n302 B.n301 163.367
R752 B.n303 B.n302 163.367
R753 B.n303 B.n52 163.367
R754 B.n307 B.n52 163.367
R755 B.n308 B.n307 163.367
R756 B.n309 B.n308 163.367
R757 B.n309 B.n50 163.367
R758 B.n313 B.n50 163.367
R759 B.n314 B.n313 163.367
R760 B.n315 B.n314 163.367
R761 B.n315 B.n48 163.367
R762 B.n319 B.n48 163.367
R763 B.n320 B.n319 163.367
R764 B.n321 B.n320 163.367
R765 B.n321 B.n46 163.367
R766 B.n325 B.n46 163.367
R767 B.n326 B.n325 163.367
R768 B.n327 B.n326 163.367
R769 B.n327 B.n44 163.367
R770 B.n331 B.n44 163.367
R771 B.n332 B.n331 163.367
R772 B.n388 B.n387 163.367
R773 B.n387 B.n386 163.367
R774 B.n386 B.n21 163.367
R775 B.n382 B.n21 163.367
R776 B.n382 B.n381 163.367
R777 B.n381 B.n380 163.367
R778 B.n380 B.n23 163.367
R779 B.n376 B.n23 163.367
R780 B.n376 B.n375 163.367
R781 B.n375 B.n374 163.367
R782 B.n374 B.n25 163.367
R783 B.n370 B.n25 163.367
R784 B.n370 B.n369 163.367
R785 B.n369 B.n368 163.367
R786 B.n368 B.n27 163.367
R787 B.n364 B.n27 163.367
R788 B.n364 B.n363 163.367
R789 B.n363 B.n362 163.367
R790 B.n362 B.n32 163.367
R791 B.n358 B.n32 163.367
R792 B.n358 B.n357 163.367
R793 B.n357 B.n356 163.367
R794 B.n356 B.n34 163.367
R795 B.n351 B.n34 163.367
R796 B.n351 B.n350 163.367
R797 B.n350 B.n349 163.367
R798 B.n349 B.n38 163.367
R799 B.n345 B.n38 163.367
R800 B.n345 B.n344 163.367
R801 B.n344 B.n343 163.367
R802 B.n343 B.n40 163.367
R803 B.n339 B.n40 163.367
R804 B.n339 B.n338 163.367
R805 B.n338 B.n337 163.367
R806 B.n337 B.n42 163.367
R807 B.n333 B.n42 163.367
R808 B.n203 B.n202 59.5399
R809 B.n188 B.n92 59.5399
R810 B.n30 B.n29 59.5399
R811 B.n354 B.n36 59.5399
R812 B.n390 B.n389 33.5615
R813 B.n334 B.n43 33.5615
R814 B.n227 B.n226 33.5615
R815 B.n168 B.n99 33.5615
R816 B.n202 B.n201 29.6732
R817 B.n92 B.n91 29.6732
R818 B.n29 B.n28 29.6732
R819 B.n36 B.n35 29.6732
R820 B B.n443 18.0485
R821 B.n389 B.n20 10.6151
R822 B.n385 B.n20 10.6151
R823 B.n385 B.n384 10.6151
R824 B.n384 B.n383 10.6151
R825 B.n383 B.n22 10.6151
R826 B.n379 B.n22 10.6151
R827 B.n379 B.n378 10.6151
R828 B.n378 B.n377 10.6151
R829 B.n377 B.n24 10.6151
R830 B.n373 B.n24 10.6151
R831 B.n373 B.n372 10.6151
R832 B.n372 B.n371 10.6151
R833 B.n371 B.n26 10.6151
R834 B.n367 B.n366 10.6151
R835 B.n366 B.n365 10.6151
R836 B.n365 B.n31 10.6151
R837 B.n361 B.n31 10.6151
R838 B.n361 B.n360 10.6151
R839 B.n360 B.n359 10.6151
R840 B.n359 B.n33 10.6151
R841 B.n355 B.n33 10.6151
R842 B.n353 B.n352 10.6151
R843 B.n352 B.n37 10.6151
R844 B.n348 B.n37 10.6151
R845 B.n348 B.n347 10.6151
R846 B.n347 B.n346 10.6151
R847 B.n346 B.n39 10.6151
R848 B.n342 B.n39 10.6151
R849 B.n342 B.n341 10.6151
R850 B.n341 B.n340 10.6151
R851 B.n340 B.n41 10.6151
R852 B.n336 B.n41 10.6151
R853 B.n336 B.n335 10.6151
R854 B.n335 B.n334 10.6151
R855 B.n228 B.n227 10.6151
R856 B.n228 B.n77 10.6151
R857 B.n232 B.n77 10.6151
R858 B.n233 B.n232 10.6151
R859 B.n234 B.n233 10.6151
R860 B.n234 B.n75 10.6151
R861 B.n238 B.n75 10.6151
R862 B.n239 B.n238 10.6151
R863 B.n240 B.n239 10.6151
R864 B.n240 B.n73 10.6151
R865 B.n244 B.n73 10.6151
R866 B.n245 B.n244 10.6151
R867 B.n246 B.n245 10.6151
R868 B.n246 B.n71 10.6151
R869 B.n250 B.n71 10.6151
R870 B.n251 B.n250 10.6151
R871 B.n252 B.n251 10.6151
R872 B.n252 B.n69 10.6151
R873 B.n256 B.n69 10.6151
R874 B.n257 B.n256 10.6151
R875 B.n258 B.n257 10.6151
R876 B.n258 B.n67 10.6151
R877 B.n262 B.n67 10.6151
R878 B.n263 B.n262 10.6151
R879 B.n264 B.n263 10.6151
R880 B.n264 B.n65 10.6151
R881 B.n268 B.n65 10.6151
R882 B.n269 B.n268 10.6151
R883 B.n270 B.n269 10.6151
R884 B.n270 B.n63 10.6151
R885 B.n274 B.n63 10.6151
R886 B.n275 B.n274 10.6151
R887 B.n276 B.n275 10.6151
R888 B.n276 B.n61 10.6151
R889 B.n280 B.n61 10.6151
R890 B.n281 B.n280 10.6151
R891 B.n282 B.n281 10.6151
R892 B.n282 B.n59 10.6151
R893 B.n286 B.n59 10.6151
R894 B.n287 B.n286 10.6151
R895 B.n288 B.n287 10.6151
R896 B.n288 B.n57 10.6151
R897 B.n292 B.n57 10.6151
R898 B.n293 B.n292 10.6151
R899 B.n294 B.n293 10.6151
R900 B.n294 B.n55 10.6151
R901 B.n298 B.n55 10.6151
R902 B.n299 B.n298 10.6151
R903 B.n300 B.n299 10.6151
R904 B.n300 B.n53 10.6151
R905 B.n304 B.n53 10.6151
R906 B.n305 B.n304 10.6151
R907 B.n306 B.n305 10.6151
R908 B.n306 B.n51 10.6151
R909 B.n310 B.n51 10.6151
R910 B.n311 B.n310 10.6151
R911 B.n312 B.n311 10.6151
R912 B.n312 B.n49 10.6151
R913 B.n316 B.n49 10.6151
R914 B.n317 B.n316 10.6151
R915 B.n318 B.n317 10.6151
R916 B.n318 B.n47 10.6151
R917 B.n322 B.n47 10.6151
R918 B.n323 B.n322 10.6151
R919 B.n324 B.n323 10.6151
R920 B.n324 B.n45 10.6151
R921 B.n328 B.n45 10.6151
R922 B.n329 B.n328 10.6151
R923 B.n330 B.n329 10.6151
R924 B.n330 B.n43 10.6151
R925 B.n169 B.n168 10.6151
R926 B.n170 B.n169 10.6151
R927 B.n170 B.n97 10.6151
R928 B.n174 B.n97 10.6151
R929 B.n175 B.n174 10.6151
R930 B.n176 B.n175 10.6151
R931 B.n176 B.n95 10.6151
R932 B.n180 B.n95 10.6151
R933 B.n181 B.n180 10.6151
R934 B.n182 B.n181 10.6151
R935 B.n182 B.n93 10.6151
R936 B.n186 B.n93 10.6151
R937 B.n187 B.n186 10.6151
R938 B.n189 B.n89 10.6151
R939 B.n193 B.n89 10.6151
R940 B.n194 B.n193 10.6151
R941 B.n195 B.n194 10.6151
R942 B.n195 B.n87 10.6151
R943 B.n199 B.n87 10.6151
R944 B.n200 B.n199 10.6151
R945 B.n204 B.n200 10.6151
R946 B.n208 B.n85 10.6151
R947 B.n209 B.n208 10.6151
R948 B.n210 B.n209 10.6151
R949 B.n210 B.n83 10.6151
R950 B.n214 B.n83 10.6151
R951 B.n215 B.n214 10.6151
R952 B.n216 B.n215 10.6151
R953 B.n216 B.n81 10.6151
R954 B.n220 B.n81 10.6151
R955 B.n221 B.n220 10.6151
R956 B.n222 B.n221 10.6151
R957 B.n222 B.n79 10.6151
R958 B.n226 B.n79 10.6151
R959 B.n164 B.n99 10.6151
R960 B.n164 B.n163 10.6151
R961 B.n163 B.n162 10.6151
R962 B.n162 B.n101 10.6151
R963 B.n158 B.n101 10.6151
R964 B.n158 B.n157 10.6151
R965 B.n157 B.n156 10.6151
R966 B.n156 B.n103 10.6151
R967 B.n152 B.n103 10.6151
R968 B.n152 B.n151 10.6151
R969 B.n151 B.n150 10.6151
R970 B.n150 B.n105 10.6151
R971 B.n146 B.n105 10.6151
R972 B.n146 B.n145 10.6151
R973 B.n145 B.n144 10.6151
R974 B.n144 B.n107 10.6151
R975 B.n140 B.n107 10.6151
R976 B.n140 B.n139 10.6151
R977 B.n139 B.n138 10.6151
R978 B.n138 B.n109 10.6151
R979 B.n134 B.n109 10.6151
R980 B.n134 B.n133 10.6151
R981 B.n133 B.n132 10.6151
R982 B.n132 B.n111 10.6151
R983 B.n128 B.n111 10.6151
R984 B.n128 B.n127 10.6151
R985 B.n127 B.n126 10.6151
R986 B.n126 B.n113 10.6151
R987 B.n122 B.n113 10.6151
R988 B.n122 B.n121 10.6151
R989 B.n121 B.n120 10.6151
R990 B.n120 B.n115 10.6151
R991 B.n116 B.n115 10.6151
R992 B.n116 B.n0 10.6151
R993 B.n439 B.n1 10.6151
R994 B.n439 B.n438 10.6151
R995 B.n438 B.n437 10.6151
R996 B.n437 B.n4 10.6151
R997 B.n433 B.n4 10.6151
R998 B.n433 B.n432 10.6151
R999 B.n432 B.n431 10.6151
R1000 B.n431 B.n6 10.6151
R1001 B.n427 B.n6 10.6151
R1002 B.n427 B.n426 10.6151
R1003 B.n426 B.n425 10.6151
R1004 B.n425 B.n8 10.6151
R1005 B.n421 B.n8 10.6151
R1006 B.n421 B.n420 10.6151
R1007 B.n420 B.n419 10.6151
R1008 B.n419 B.n10 10.6151
R1009 B.n415 B.n10 10.6151
R1010 B.n415 B.n414 10.6151
R1011 B.n414 B.n413 10.6151
R1012 B.n413 B.n12 10.6151
R1013 B.n409 B.n12 10.6151
R1014 B.n409 B.n408 10.6151
R1015 B.n408 B.n407 10.6151
R1016 B.n407 B.n14 10.6151
R1017 B.n403 B.n14 10.6151
R1018 B.n403 B.n402 10.6151
R1019 B.n402 B.n401 10.6151
R1020 B.n401 B.n16 10.6151
R1021 B.n397 B.n16 10.6151
R1022 B.n397 B.n396 10.6151
R1023 B.n396 B.n395 10.6151
R1024 B.n395 B.n18 10.6151
R1025 B.n391 B.n18 10.6151
R1026 B.n391 B.n390 10.6151
R1027 B.n367 B.n30 6.5566
R1028 B.n355 B.n354 6.5566
R1029 B.n189 B.n188 6.5566
R1030 B.n204 B.n203 6.5566
R1031 B.n30 B.n26 4.05904
R1032 B.n354 B.n353 4.05904
R1033 B.n188 B.n187 4.05904
R1034 B.n203 B.n85 4.05904
R1035 B.n443 B.n0 2.81026
R1036 B.n443 B.n1 2.81026
C0 VN w_n2806_n1470# 5.39857f
C1 w_n2806_n1470# VDD2 1.62506f
C2 VTAIL VDD1 4.88963f
C3 w_n2806_n1470# B 5.54102f
C4 VTAIL w_n2806_n1470# 1.58308f
C5 w_n2806_n1470# VDD1 1.55491f
C6 VN VP 4.58516f
C7 VDD2 VP 0.41012f
C8 B VP 1.41603f
C9 VN VDD2 2.16627f
C10 VTAIL VP 2.77482f
C11 VN B 0.817267f
C12 VDD2 B 1.26628f
C13 VTAIL VN 2.76063f
C14 VTAIL VDD2 4.93284f
C15 VTAIL B 1.15941f
C16 VDD1 VP 2.41839f
C17 w_n2806_n1470# VP 5.75638f
C18 VN VDD1 0.155554f
C19 VDD1 VDD2 1.27554f
C20 VDD1 B 1.20266f
C21 VDD2 VSUBS 1.05828f
C22 VDD1 VSUBS 1.054251f
C23 VTAIL VSUBS 0.406577f
C24 VN VSUBS 5.227611f
C25 VP VSUBS 1.959738f
C26 B VSUBS 2.678399f
C27 w_n2806_n1470# VSUBS 52.4273f
C28 B.n0 VSUBS 0.005081f
C29 B.n1 VSUBS 0.005081f
C30 B.n2 VSUBS 0.008035f
C31 B.n3 VSUBS 0.008035f
C32 B.n4 VSUBS 0.008035f
C33 B.n5 VSUBS 0.008035f
C34 B.n6 VSUBS 0.008035f
C35 B.n7 VSUBS 0.008035f
C36 B.n8 VSUBS 0.008035f
C37 B.n9 VSUBS 0.008035f
C38 B.n10 VSUBS 0.008035f
C39 B.n11 VSUBS 0.008035f
C40 B.n12 VSUBS 0.008035f
C41 B.n13 VSUBS 0.008035f
C42 B.n14 VSUBS 0.008035f
C43 B.n15 VSUBS 0.008035f
C44 B.n16 VSUBS 0.008035f
C45 B.n17 VSUBS 0.008035f
C46 B.n18 VSUBS 0.008035f
C47 B.n19 VSUBS 0.018613f
C48 B.n20 VSUBS 0.008035f
C49 B.n21 VSUBS 0.008035f
C50 B.n22 VSUBS 0.008035f
C51 B.n23 VSUBS 0.008035f
C52 B.n24 VSUBS 0.008035f
C53 B.n25 VSUBS 0.008035f
C54 B.n26 VSUBS 0.005554f
C55 B.n27 VSUBS 0.008035f
C56 B.t5 VSUBS 0.044664f
C57 B.t4 VSUBS 0.053384f
C58 B.t3 VSUBS 0.165148f
C59 B.n28 VSUBS 0.095248f
C60 B.n29 VSUBS 0.086134f
C61 B.n30 VSUBS 0.018617f
C62 B.n31 VSUBS 0.008035f
C63 B.n32 VSUBS 0.008035f
C64 B.n33 VSUBS 0.008035f
C65 B.n34 VSUBS 0.008035f
C66 B.t11 VSUBS 0.044665f
C67 B.t10 VSUBS 0.053384f
C68 B.t9 VSUBS 0.165148f
C69 B.n35 VSUBS 0.095248f
C70 B.n36 VSUBS 0.086133f
C71 B.n37 VSUBS 0.008035f
C72 B.n38 VSUBS 0.008035f
C73 B.n39 VSUBS 0.008035f
C74 B.n40 VSUBS 0.008035f
C75 B.n41 VSUBS 0.008035f
C76 B.n42 VSUBS 0.008035f
C77 B.n43 VSUBS 0.019537f
C78 B.n44 VSUBS 0.008035f
C79 B.n45 VSUBS 0.008035f
C80 B.n46 VSUBS 0.008035f
C81 B.n47 VSUBS 0.008035f
C82 B.n48 VSUBS 0.008035f
C83 B.n49 VSUBS 0.008035f
C84 B.n50 VSUBS 0.008035f
C85 B.n51 VSUBS 0.008035f
C86 B.n52 VSUBS 0.008035f
C87 B.n53 VSUBS 0.008035f
C88 B.n54 VSUBS 0.008035f
C89 B.n55 VSUBS 0.008035f
C90 B.n56 VSUBS 0.008035f
C91 B.n57 VSUBS 0.008035f
C92 B.n58 VSUBS 0.008035f
C93 B.n59 VSUBS 0.008035f
C94 B.n60 VSUBS 0.008035f
C95 B.n61 VSUBS 0.008035f
C96 B.n62 VSUBS 0.008035f
C97 B.n63 VSUBS 0.008035f
C98 B.n64 VSUBS 0.008035f
C99 B.n65 VSUBS 0.008035f
C100 B.n66 VSUBS 0.008035f
C101 B.n67 VSUBS 0.008035f
C102 B.n68 VSUBS 0.008035f
C103 B.n69 VSUBS 0.008035f
C104 B.n70 VSUBS 0.008035f
C105 B.n71 VSUBS 0.008035f
C106 B.n72 VSUBS 0.008035f
C107 B.n73 VSUBS 0.008035f
C108 B.n74 VSUBS 0.008035f
C109 B.n75 VSUBS 0.008035f
C110 B.n76 VSUBS 0.008035f
C111 B.n77 VSUBS 0.008035f
C112 B.n78 VSUBS 0.018613f
C113 B.n79 VSUBS 0.008035f
C114 B.n80 VSUBS 0.008035f
C115 B.n81 VSUBS 0.008035f
C116 B.n82 VSUBS 0.008035f
C117 B.n83 VSUBS 0.008035f
C118 B.n84 VSUBS 0.008035f
C119 B.n85 VSUBS 0.005554f
C120 B.n86 VSUBS 0.008035f
C121 B.n87 VSUBS 0.008035f
C122 B.n88 VSUBS 0.008035f
C123 B.n89 VSUBS 0.008035f
C124 B.n90 VSUBS 0.008035f
C125 B.t7 VSUBS 0.044664f
C126 B.t8 VSUBS 0.053384f
C127 B.t6 VSUBS 0.165148f
C128 B.n91 VSUBS 0.095248f
C129 B.n92 VSUBS 0.086134f
C130 B.n93 VSUBS 0.008035f
C131 B.n94 VSUBS 0.008035f
C132 B.n95 VSUBS 0.008035f
C133 B.n96 VSUBS 0.008035f
C134 B.n97 VSUBS 0.008035f
C135 B.n98 VSUBS 0.008035f
C136 B.n99 VSUBS 0.018613f
C137 B.n100 VSUBS 0.008035f
C138 B.n101 VSUBS 0.008035f
C139 B.n102 VSUBS 0.008035f
C140 B.n103 VSUBS 0.008035f
C141 B.n104 VSUBS 0.008035f
C142 B.n105 VSUBS 0.008035f
C143 B.n106 VSUBS 0.008035f
C144 B.n107 VSUBS 0.008035f
C145 B.n108 VSUBS 0.008035f
C146 B.n109 VSUBS 0.008035f
C147 B.n110 VSUBS 0.008035f
C148 B.n111 VSUBS 0.008035f
C149 B.n112 VSUBS 0.008035f
C150 B.n113 VSUBS 0.008035f
C151 B.n114 VSUBS 0.008035f
C152 B.n115 VSUBS 0.008035f
C153 B.n116 VSUBS 0.008035f
C154 B.n117 VSUBS 0.008035f
C155 B.n118 VSUBS 0.008035f
C156 B.n119 VSUBS 0.008035f
C157 B.n120 VSUBS 0.008035f
C158 B.n121 VSUBS 0.008035f
C159 B.n122 VSUBS 0.008035f
C160 B.n123 VSUBS 0.008035f
C161 B.n124 VSUBS 0.008035f
C162 B.n125 VSUBS 0.008035f
C163 B.n126 VSUBS 0.008035f
C164 B.n127 VSUBS 0.008035f
C165 B.n128 VSUBS 0.008035f
C166 B.n129 VSUBS 0.008035f
C167 B.n130 VSUBS 0.008035f
C168 B.n131 VSUBS 0.008035f
C169 B.n132 VSUBS 0.008035f
C170 B.n133 VSUBS 0.008035f
C171 B.n134 VSUBS 0.008035f
C172 B.n135 VSUBS 0.008035f
C173 B.n136 VSUBS 0.008035f
C174 B.n137 VSUBS 0.008035f
C175 B.n138 VSUBS 0.008035f
C176 B.n139 VSUBS 0.008035f
C177 B.n140 VSUBS 0.008035f
C178 B.n141 VSUBS 0.008035f
C179 B.n142 VSUBS 0.008035f
C180 B.n143 VSUBS 0.008035f
C181 B.n144 VSUBS 0.008035f
C182 B.n145 VSUBS 0.008035f
C183 B.n146 VSUBS 0.008035f
C184 B.n147 VSUBS 0.008035f
C185 B.n148 VSUBS 0.008035f
C186 B.n149 VSUBS 0.008035f
C187 B.n150 VSUBS 0.008035f
C188 B.n151 VSUBS 0.008035f
C189 B.n152 VSUBS 0.008035f
C190 B.n153 VSUBS 0.008035f
C191 B.n154 VSUBS 0.008035f
C192 B.n155 VSUBS 0.008035f
C193 B.n156 VSUBS 0.008035f
C194 B.n157 VSUBS 0.008035f
C195 B.n158 VSUBS 0.008035f
C196 B.n159 VSUBS 0.008035f
C197 B.n160 VSUBS 0.008035f
C198 B.n161 VSUBS 0.008035f
C199 B.n162 VSUBS 0.008035f
C200 B.n163 VSUBS 0.008035f
C201 B.n164 VSUBS 0.008035f
C202 B.n165 VSUBS 0.008035f
C203 B.n166 VSUBS 0.018613f
C204 B.n167 VSUBS 0.019672f
C205 B.n168 VSUBS 0.019672f
C206 B.n169 VSUBS 0.008035f
C207 B.n170 VSUBS 0.008035f
C208 B.n171 VSUBS 0.008035f
C209 B.n172 VSUBS 0.008035f
C210 B.n173 VSUBS 0.008035f
C211 B.n174 VSUBS 0.008035f
C212 B.n175 VSUBS 0.008035f
C213 B.n176 VSUBS 0.008035f
C214 B.n177 VSUBS 0.008035f
C215 B.n178 VSUBS 0.008035f
C216 B.n179 VSUBS 0.008035f
C217 B.n180 VSUBS 0.008035f
C218 B.n181 VSUBS 0.008035f
C219 B.n182 VSUBS 0.008035f
C220 B.n183 VSUBS 0.008035f
C221 B.n184 VSUBS 0.008035f
C222 B.n185 VSUBS 0.008035f
C223 B.n186 VSUBS 0.008035f
C224 B.n187 VSUBS 0.005554f
C225 B.n188 VSUBS 0.018617f
C226 B.n189 VSUBS 0.006499f
C227 B.n190 VSUBS 0.008035f
C228 B.n191 VSUBS 0.008035f
C229 B.n192 VSUBS 0.008035f
C230 B.n193 VSUBS 0.008035f
C231 B.n194 VSUBS 0.008035f
C232 B.n195 VSUBS 0.008035f
C233 B.n196 VSUBS 0.008035f
C234 B.n197 VSUBS 0.008035f
C235 B.n198 VSUBS 0.008035f
C236 B.n199 VSUBS 0.008035f
C237 B.n200 VSUBS 0.008035f
C238 B.t1 VSUBS 0.044665f
C239 B.t2 VSUBS 0.053384f
C240 B.t0 VSUBS 0.165148f
C241 B.n201 VSUBS 0.095248f
C242 B.n202 VSUBS 0.086133f
C243 B.n203 VSUBS 0.018617f
C244 B.n204 VSUBS 0.006499f
C245 B.n205 VSUBS 0.008035f
C246 B.n206 VSUBS 0.008035f
C247 B.n207 VSUBS 0.008035f
C248 B.n208 VSUBS 0.008035f
C249 B.n209 VSUBS 0.008035f
C250 B.n210 VSUBS 0.008035f
C251 B.n211 VSUBS 0.008035f
C252 B.n212 VSUBS 0.008035f
C253 B.n213 VSUBS 0.008035f
C254 B.n214 VSUBS 0.008035f
C255 B.n215 VSUBS 0.008035f
C256 B.n216 VSUBS 0.008035f
C257 B.n217 VSUBS 0.008035f
C258 B.n218 VSUBS 0.008035f
C259 B.n219 VSUBS 0.008035f
C260 B.n220 VSUBS 0.008035f
C261 B.n221 VSUBS 0.008035f
C262 B.n222 VSUBS 0.008035f
C263 B.n223 VSUBS 0.008035f
C264 B.n224 VSUBS 0.008035f
C265 B.n225 VSUBS 0.019672f
C266 B.n226 VSUBS 0.019672f
C267 B.n227 VSUBS 0.018613f
C268 B.n228 VSUBS 0.008035f
C269 B.n229 VSUBS 0.008035f
C270 B.n230 VSUBS 0.008035f
C271 B.n231 VSUBS 0.008035f
C272 B.n232 VSUBS 0.008035f
C273 B.n233 VSUBS 0.008035f
C274 B.n234 VSUBS 0.008035f
C275 B.n235 VSUBS 0.008035f
C276 B.n236 VSUBS 0.008035f
C277 B.n237 VSUBS 0.008035f
C278 B.n238 VSUBS 0.008035f
C279 B.n239 VSUBS 0.008035f
C280 B.n240 VSUBS 0.008035f
C281 B.n241 VSUBS 0.008035f
C282 B.n242 VSUBS 0.008035f
C283 B.n243 VSUBS 0.008035f
C284 B.n244 VSUBS 0.008035f
C285 B.n245 VSUBS 0.008035f
C286 B.n246 VSUBS 0.008035f
C287 B.n247 VSUBS 0.008035f
C288 B.n248 VSUBS 0.008035f
C289 B.n249 VSUBS 0.008035f
C290 B.n250 VSUBS 0.008035f
C291 B.n251 VSUBS 0.008035f
C292 B.n252 VSUBS 0.008035f
C293 B.n253 VSUBS 0.008035f
C294 B.n254 VSUBS 0.008035f
C295 B.n255 VSUBS 0.008035f
C296 B.n256 VSUBS 0.008035f
C297 B.n257 VSUBS 0.008035f
C298 B.n258 VSUBS 0.008035f
C299 B.n259 VSUBS 0.008035f
C300 B.n260 VSUBS 0.008035f
C301 B.n261 VSUBS 0.008035f
C302 B.n262 VSUBS 0.008035f
C303 B.n263 VSUBS 0.008035f
C304 B.n264 VSUBS 0.008035f
C305 B.n265 VSUBS 0.008035f
C306 B.n266 VSUBS 0.008035f
C307 B.n267 VSUBS 0.008035f
C308 B.n268 VSUBS 0.008035f
C309 B.n269 VSUBS 0.008035f
C310 B.n270 VSUBS 0.008035f
C311 B.n271 VSUBS 0.008035f
C312 B.n272 VSUBS 0.008035f
C313 B.n273 VSUBS 0.008035f
C314 B.n274 VSUBS 0.008035f
C315 B.n275 VSUBS 0.008035f
C316 B.n276 VSUBS 0.008035f
C317 B.n277 VSUBS 0.008035f
C318 B.n278 VSUBS 0.008035f
C319 B.n279 VSUBS 0.008035f
C320 B.n280 VSUBS 0.008035f
C321 B.n281 VSUBS 0.008035f
C322 B.n282 VSUBS 0.008035f
C323 B.n283 VSUBS 0.008035f
C324 B.n284 VSUBS 0.008035f
C325 B.n285 VSUBS 0.008035f
C326 B.n286 VSUBS 0.008035f
C327 B.n287 VSUBS 0.008035f
C328 B.n288 VSUBS 0.008035f
C329 B.n289 VSUBS 0.008035f
C330 B.n290 VSUBS 0.008035f
C331 B.n291 VSUBS 0.008035f
C332 B.n292 VSUBS 0.008035f
C333 B.n293 VSUBS 0.008035f
C334 B.n294 VSUBS 0.008035f
C335 B.n295 VSUBS 0.008035f
C336 B.n296 VSUBS 0.008035f
C337 B.n297 VSUBS 0.008035f
C338 B.n298 VSUBS 0.008035f
C339 B.n299 VSUBS 0.008035f
C340 B.n300 VSUBS 0.008035f
C341 B.n301 VSUBS 0.008035f
C342 B.n302 VSUBS 0.008035f
C343 B.n303 VSUBS 0.008035f
C344 B.n304 VSUBS 0.008035f
C345 B.n305 VSUBS 0.008035f
C346 B.n306 VSUBS 0.008035f
C347 B.n307 VSUBS 0.008035f
C348 B.n308 VSUBS 0.008035f
C349 B.n309 VSUBS 0.008035f
C350 B.n310 VSUBS 0.008035f
C351 B.n311 VSUBS 0.008035f
C352 B.n312 VSUBS 0.008035f
C353 B.n313 VSUBS 0.008035f
C354 B.n314 VSUBS 0.008035f
C355 B.n315 VSUBS 0.008035f
C356 B.n316 VSUBS 0.008035f
C357 B.n317 VSUBS 0.008035f
C358 B.n318 VSUBS 0.008035f
C359 B.n319 VSUBS 0.008035f
C360 B.n320 VSUBS 0.008035f
C361 B.n321 VSUBS 0.008035f
C362 B.n322 VSUBS 0.008035f
C363 B.n323 VSUBS 0.008035f
C364 B.n324 VSUBS 0.008035f
C365 B.n325 VSUBS 0.008035f
C366 B.n326 VSUBS 0.008035f
C367 B.n327 VSUBS 0.008035f
C368 B.n328 VSUBS 0.008035f
C369 B.n329 VSUBS 0.008035f
C370 B.n330 VSUBS 0.008035f
C371 B.n331 VSUBS 0.008035f
C372 B.n332 VSUBS 0.018613f
C373 B.n333 VSUBS 0.019672f
C374 B.n334 VSUBS 0.018748f
C375 B.n335 VSUBS 0.008035f
C376 B.n336 VSUBS 0.008035f
C377 B.n337 VSUBS 0.008035f
C378 B.n338 VSUBS 0.008035f
C379 B.n339 VSUBS 0.008035f
C380 B.n340 VSUBS 0.008035f
C381 B.n341 VSUBS 0.008035f
C382 B.n342 VSUBS 0.008035f
C383 B.n343 VSUBS 0.008035f
C384 B.n344 VSUBS 0.008035f
C385 B.n345 VSUBS 0.008035f
C386 B.n346 VSUBS 0.008035f
C387 B.n347 VSUBS 0.008035f
C388 B.n348 VSUBS 0.008035f
C389 B.n349 VSUBS 0.008035f
C390 B.n350 VSUBS 0.008035f
C391 B.n351 VSUBS 0.008035f
C392 B.n352 VSUBS 0.008035f
C393 B.n353 VSUBS 0.005554f
C394 B.n354 VSUBS 0.018617f
C395 B.n355 VSUBS 0.006499f
C396 B.n356 VSUBS 0.008035f
C397 B.n357 VSUBS 0.008035f
C398 B.n358 VSUBS 0.008035f
C399 B.n359 VSUBS 0.008035f
C400 B.n360 VSUBS 0.008035f
C401 B.n361 VSUBS 0.008035f
C402 B.n362 VSUBS 0.008035f
C403 B.n363 VSUBS 0.008035f
C404 B.n364 VSUBS 0.008035f
C405 B.n365 VSUBS 0.008035f
C406 B.n366 VSUBS 0.008035f
C407 B.n367 VSUBS 0.006499f
C408 B.n368 VSUBS 0.008035f
C409 B.n369 VSUBS 0.008035f
C410 B.n370 VSUBS 0.008035f
C411 B.n371 VSUBS 0.008035f
C412 B.n372 VSUBS 0.008035f
C413 B.n373 VSUBS 0.008035f
C414 B.n374 VSUBS 0.008035f
C415 B.n375 VSUBS 0.008035f
C416 B.n376 VSUBS 0.008035f
C417 B.n377 VSUBS 0.008035f
C418 B.n378 VSUBS 0.008035f
C419 B.n379 VSUBS 0.008035f
C420 B.n380 VSUBS 0.008035f
C421 B.n381 VSUBS 0.008035f
C422 B.n382 VSUBS 0.008035f
C423 B.n383 VSUBS 0.008035f
C424 B.n384 VSUBS 0.008035f
C425 B.n385 VSUBS 0.008035f
C426 B.n386 VSUBS 0.008035f
C427 B.n387 VSUBS 0.008035f
C428 B.n388 VSUBS 0.019672f
C429 B.n389 VSUBS 0.019672f
C430 B.n390 VSUBS 0.018613f
C431 B.n391 VSUBS 0.008035f
C432 B.n392 VSUBS 0.008035f
C433 B.n393 VSUBS 0.008035f
C434 B.n394 VSUBS 0.008035f
C435 B.n395 VSUBS 0.008035f
C436 B.n396 VSUBS 0.008035f
C437 B.n397 VSUBS 0.008035f
C438 B.n398 VSUBS 0.008035f
C439 B.n399 VSUBS 0.008035f
C440 B.n400 VSUBS 0.008035f
C441 B.n401 VSUBS 0.008035f
C442 B.n402 VSUBS 0.008035f
C443 B.n403 VSUBS 0.008035f
C444 B.n404 VSUBS 0.008035f
C445 B.n405 VSUBS 0.008035f
C446 B.n406 VSUBS 0.008035f
C447 B.n407 VSUBS 0.008035f
C448 B.n408 VSUBS 0.008035f
C449 B.n409 VSUBS 0.008035f
C450 B.n410 VSUBS 0.008035f
C451 B.n411 VSUBS 0.008035f
C452 B.n412 VSUBS 0.008035f
C453 B.n413 VSUBS 0.008035f
C454 B.n414 VSUBS 0.008035f
C455 B.n415 VSUBS 0.008035f
C456 B.n416 VSUBS 0.008035f
C457 B.n417 VSUBS 0.008035f
C458 B.n418 VSUBS 0.008035f
C459 B.n419 VSUBS 0.008035f
C460 B.n420 VSUBS 0.008035f
C461 B.n421 VSUBS 0.008035f
C462 B.n422 VSUBS 0.008035f
C463 B.n423 VSUBS 0.008035f
C464 B.n424 VSUBS 0.008035f
C465 B.n425 VSUBS 0.008035f
C466 B.n426 VSUBS 0.008035f
C467 B.n427 VSUBS 0.008035f
C468 B.n428 VSUBS 0.008035f
C469 B.n429 VSUBS 0.008035f
C470 B.n430 VSUBS 0.008035f
C471 B.n431 VSUBS 0.008035f
C472 B.n432 VSUBS 0.008035f
C473 B.n433 VSUBS 0.008035f
C474 B.n434 VSUBS 0.008035f
C475 B.n435 VSUBS 0.008035f
C476 B.n436 VSUBS 0.008035f
C477 B.n437 VSUBS 0.008035f
C478 B.n438 VSUBS 0.008035f
C479 B.n439 VSUBS 0.008035f
C480 B.n440 VSUBS 0.008035f
C481 B.n441 VSUBS 0.008035f
C482 B.n442 VSUBS 0.008035f
C483 B.n443 VSUBS 0.018194f
C484 VDD2.n0 VSUBS 0.024929f
C485 VDD2.n1 VSUBS 0.167329f
C486 VDD2.n2 VSUBS 0.01268f
C487 VDD2.t4 VSUBS 0.066978f
C488 VDD2.n3 VSUBS 0.078655f
C489 VDD2.n4 VSUBS 0.017671f
C490 VDD2.n5 VSUBS 0.022478f
C491 VDD2.n6 VSUBS 0.069152f
C492 VDD2.n7 VSUBS 0.013426f
C493 VDD2.n8 VSUBS 0.01268f
C494 VDD2.n9 VSUBS 0.058088f
C495 VDD2.n10 VSUBS 0.054723f
C496 VDD2.t6 VSUBS 0.046803f
C497 VDD2.t7 VSUBS 0.046803f
C498 VDD2.n11 VSUBS 0.228848f
C499 VDD2.n12 VSUBS 0.543704f
C500 VDD2.t9 VSUBS 0.046803f
C501 VDD2.t1 VSUBS 0.046803f
C502 VDD2.n13 VSUBS 0.231611f
C503 VDD2.n14 VSUBS 1.60399f
C504 VDD2.n15 VSUBS 0.024929f
C505 VDD2.n16 VSUBS 0.167329f
C506 VDD2.n17 VSUBS 0.01268f
C507 VDD2.t8 VSUBS 0.066978f
C508 VDD2.n18 VSUBS 0.078655f
C509 VDD2.n19 VSUBS 0.017671f
C510 VDD2.n20 VSUBS 0.022478f
C511 VDD2.n21 VSUBS 0.069152f
C512 VDD2.n22 VSUBS 0.013426f
C513 VDD2.n23 VSUBS 0.01268f
C514 VDD2.n24 VSUBS 0.058088f
C515 VDD2.n25 VSUBS 0.050998f
C516 VDD2.n26 VSUBS 1.50215f
C517 VDD2.t0 VSUBS 0.046803f
C518 VDD2.t2 VSUBS 0.046803f
C519 VDD2.n27 VSUBS 0.228849f
C520 VDD2.n28 VSUBS 0.406314f
C521 VDD2.t3 VSUBS 0.046803f
C522 VDD2.t5 VSUBS 0.046803f
C523 VDD2.n29 VSUBS 0.231598f
C524 VN.n0 VSUBS 0.080575f
C525 VN.t0 VSUBS 0.442017f
C526 VN.n1 VSUBS 0.225465f
C527 VN.n2 VSUBS 0.060384f
C528 VN.t2 VSUBS 0.442017f
C529 VN.n3 VSUBS 0.225465f
C530 VN.n4 VSUBS 0.060384f
C531 VN.t3 VSUBS 0.442017f
C532 VN.n5 VSUBS 0.30352f
C533 VN.t5 VSUBS 0.61796f
C534 VN.n6 VSUBS 0.324516f
C535 VN.n7 VSUBS 0.311064f
C536 VN.n8 VSUBS 0.094578f
C537 VN.n9 VSUBS 0.048992f
C538 VN.n10 VSUBS 0.093055f
C539 VN.n11 VSUBS 0.060384f
C540 VN.n12 VSUBS 0.060384f
C541 VN.n13 VSUBS 0.093055f
C542 VN.n14 VSUBS 0.048992f
C543 VN.n15 VSUBS 0.094578f
C544 VN.n16 VSUBS 0.060384f
C545 VN.n17 VSUBS 0.060384f
C546 VN.n18 VSUBS 0.090749f
C547 VN.n19 VSUBS 0.03774f
C548 VN.t8 VSUBS 0.553029f
C549 VN.n20 VSUBS 0.336242f
C550 VN.n21 VSUBS 0.056552f
C551 VN.n22 VSUBS 0.080575f
C552 VN.t9 VSUBS 0.442017f
C553 VN.n23 VSUBS 0.225465f
C554 VN.n24 VSUBS 0.060384f
C555 VN.t7 VSUBS 0.442017f
C556 VN.n25 VSUBS 0.225465f
C557 VN.n26 VSUBS 0.060384f
C558 VN.t6 VSUBS 0.442017f
C559 VN.n27 VSUBS 0.30352f
C560 VN.t4 VSUBS 0.61796f
C561 VN.n28 VSUBS 0.324516f
C562 VN.n29 VSUBS 0.311064f
C563 VN.n30 VSUBS 0.094578f
C564 VN.n31 VSUBS 0.048992f
C565 VN.n32 VSUBS 0.093055f
C566 VN.n33 VSUBS 0.060384f
C567 VN.n34 VSUBS 0.060384f
C568 VN.n35 VSUBS 0.093055f
C569 VN.n36 VSUBS 0.048992f
C570 VN.n37 VSUBS 0.094578f
C571 VN.n38 VSUBS 0.060384f
C572 VN.n39 VSUBS 0.060384f
C573 VN.n40 VSUBS 0.090749f
C574 VN.n41 VSUBS 0.03774f
C575 VN.t1 VSUBS 0.553029f
C576 VN.n42 VSUBS 0.336242f
C577 VN.n43 VSUBS 2.19582f
C578 VDD1.n0 VSUBS 0.02532f
C579 VDD1.n1 VSUBS 0.169957f
C580 VDD1.n2 VSUBS 0.012879f
C581 VDD1.t4 VSUBS 0.06803f
C582 VDD1.n3 VSUBS 0.07989f
C583 VDD1.n4 VSUBS 0.017949f
C584 VDD1.n5 VSUBS 0.022831f
C585 VDD1.n6 VSUBS 0.070238f
C586 VDD1.n7 VSUBS 0.013636f
C587 VDD1.n8 VSUBS 0.012879f
C588 VDD1.n9 VSUBS 0.059f
C589 VDD1.n10 VSUBS 0.055582f
C590 VDD1.t0 VSUBS 0.047538f
C591 VDD1.t9 VSUBS 0.047538f
C592 VDD1.n11 VSUBS 0.232442f
C593 VDD1.n12 VSUBS 0.558983f
C594 VDD1.n13 VSUBS 0.02532f
C595 VDD1.n14 VSUBS 0.169957f
C596 VDD1.n15 VSUBS 0.012879f
C597 VDD1.t5 VSUBS 0.06803f
C598 VDD1.n16 VSUBS 0.07989f
C599 VDD1.n17 VSUBS 0.017949f
C600 VDD1.n18 VSUBS 0.022831f
C601 VDD1.n19 VSUBS 0.070238f
C602 VDD1.n20 VSUBS 0.013636f
C603 VDD1.n21 VSUBS 0.012879f
C604 VDD1.n22 VSUBS 0.059f
C605 VDD1.n23 VSUBS 0.055582f
C606 VDD1.t3 VSUBS 0.047538f
C607 VDD1.t1 VSUBS 0.047538f
C608 VDD1.n24 VSUBS 0.232441f
C609 VDD1.n25 VSUBS 0.552241f
C610 VDD1.t2 VSUBS 0.047538f
C611 VDD1.t7 VSUBS 0.047538f
C612 VDD1.n26 VSUBS 0.235247f
C613 VDD1.n27 VSUBS 1.70873f
C614 VDD1.t8 VSUBS 0.047538f
C615 VDD1.t6 VSUBS 0.047538f
C616 VDD1.n28 VSUBS 0.232441f
C617 VDD1.n29 VSUBS 1.84893f
C618 VTAIL.t6 VSUBS 0.063065f
C619 VTAIL.t5 VSUBS 0.063065f
C620 VTAIL.n0 VSUBS 0.263789f
C621 VTAIL.n1 VSUBS 0.596973f
C622 VTAIL.n2 VSUBS 0.03359f
C623 VTAIL.n3 VSUBS 0.225466f
C624 VTAIL.n4 VSUBS 0.017085f
C625 VTAIL.t15 VSUBS 0.090249f
C626 VTAIL.n5 VSUBS 0.105983f
C627 VTAIL.n6 VSUBS 0.023811f
C628 VTAIL.n7 VSUBS 0.030287f
C629 VTAIL.n8 VSUBS 0.093179f
C630 VTAIL.n9 VSUBS 0.01809f
C631 VTAIL.n10 VSUBS 0.017085f
C632 VTAIL.n11 VSUBS 0.07827f
C633 VTAIL.n12 VSUBS 0.046798f
C634 VTAIL.n13 VSUBS 0.280682f
C635 VTAIL.t18 VSUBS 0.063065f
C636 VTAIL.t14 VSUBS 0.063065f
C637 VTAIL.n14 VSUBS 0.263789f
C638 VTAIL.n15 VSUBS 0.644223f
C639 VTAIL.t12 VSUBS 0.063065f
C640 VTAIL.t13 VSUBS 0.063065f
C641 VTAIL.n16 VSUBS 0.263789f
C642 VTAIL.n17 VSUBS 1.43293f
C643 VTAIL.t7 VSUBS 0.063065f
C644 VTAIL.t9 VSUBS 0.063065f
C645 VTAIL.n18 VSUBS 0.263791f
C646 VTAIL.n19 VSUBS 1.43293f
C647 VTAIL.t8 VSUBS 0.063065f
C648 VTAIL.t2 VSUBS 0.063065f
C649 VTAIL.n20 VSUBS 0.263791f
C650 VTAIL.n21 VSUBS 0.644222f
C651 VTAIL.n22 VSUBS 0.03359f
C652 VTAIL.n23 VSUBS 0.225466f
C653 VTAIL.n24 VSUBS 0.017085f
C654 VTAIL.t1 VSUBS 0.090249f
C655 VTAIL.n25 VSUBS 0.105983f
C656 VTAIL.n26 VSUBS 0.023811f
C657 VTAIL.n27 VSUBS 0.030287f
C658 VTAIL.n28 VSUBS 0.093179f
C659 VTAIL.n29 VSUBS 0.01809f
C660 VTAIL.n30 VSUBS 0.017085f
C661 VTAIL.n31 VSUBS 0.07827f
C662 VTAIL.n32 VSUBS 0.046798f
C663 VTAIL.n33 VSUBS 0.280682f
C664 VTAIL.t17 VSUBS 0.063065f
C665 VTAIL.t19 VSUBS 0.063065f
C666 VTAIL.n34 VSUBS 0.263791f
C667 VTAIL.n35 VSUBS 0.624792f
C668 VTAIL.t10 VSUBS 0.063065f
C669 VTAIL.t11 VSUBS 0.063065f
C670 VTAIL.n36 VSUBS 0.263791f
C671 VTAIL.n37 VSUBS 0.644222f
C672 VTAIL.n38 VSUBS 0.03359f
C673 VTAIL.n39 VSUBS 0.225466f
C674 VTAIL.n40 VSUBS 0.017085f
C675 VTAIL.t16 VSUBS 0.090249f
C676 VTAIL.n41 VSUBS 0.105983f
C677 VTAIL.n42 VSUBS 0.023811f
C678 VTAIL.n43 VSUBS 0.030287f
C679 VTAIL.n44 VSUBS 0.093179f
C680 VTAIL.n45 VSUBS 0.01809f
C681 VTAIL.n46 VSUBS 0.017085f
C682 VTAIL.n47 VSUBS 0.07827f
C683 VTAIL.n48 VSUBS 0.046798f
C684 VTAIL.n49 VSUBS 0.95369f
C685 VTAIL.n50 VSUBS 0.03359f
C686 VTAIL.n51 VSUBS 0.225466f
C687 VTAIL.n52 VSUBS 0.017085f
C688 VTAIL.t3 VSUBS 0.090249f
C689 VTAIL.n53 VSUBS 0.105983f
C690 VTAIL.n54 VSUBS 0.023811f
C691 VTAIL.n55 VSUBS 0.030287f
C692 VTAIL.n56 VSUBS 0.093179f
C693 VTAIL.n57 VSUBS 0.01809f
C694 VTAIL.n58 VSUBS 0.017085f
C695 VTAIL.n59 VSUBS 0.07827f
C696 VTAIL.n60 VSUBS 0.046798f
C697 VTAIL.n61 VSUBS 0.95369f
C698 VTAIL.t0 VSUBS 0.063065f
C699 VTAIL.t4 VSUBS 0.063065f
C700 VTAIL.n62 VSUBS 0.263789f
C701 VTAIL.n63 VSUBS 0.536915f
C702 VP.n0 VSUBS 0.084275f
C703 VP.t7 VSUBS 0.462314f
C704 VP.n1 VSUBS 0.235818f
C705 VP.n2 VSUBS 0.063157f
C706 VP.t8 VSUBS 0.462314f
C707 VP.n3 VSUBS 0.235818f
C708 VP.n4 VSUBS 0.063157f
C709 VP.t6 VSUBS 0.462314f
C710 VP.n5 VSUBS 0.235818f
C711 VP.n6 VSUBS 0.084275f
C712 VP.n7 VSUBS 0.084275f
C713 VP.t3 VSUBS 0.578424f
C714 VP.t1 VSUBS 0.462314f
C715 VP.n8 VSUBS 0.235818f
C716 VP.n9 VSUBS 0.063157f
C717 VP.t0 VSUBS 0.462314f
C718 VP.n10 VSUBS 0.235818f
C719 VP.n11 VSUBS 0.063157f
C720 VP.t9 VSUBS 0.462314f
C721 VP.n12 VSUBS 0.317457f
C722 VP.t5 VSUBS 0.646336f
C723 VP.n13 VSUBS 0.339418f
C724 VP.n14 VSUBS 0.325348f
C725 VP.n15 VSUBS 0.098921f
C726 VP.n16 VSUBS 0.051242f
C727 VP.n17 VSUBS 0.097328f
C728 VP.n18 VSUBS 0.063157f
C729 VP.n19 VSUBS 0.063157f
C730 VP.n20 VSUBS 0.097328f
C731 VP.n21 VSUBS 0.051242f
C732 VP.n22 VSUBS 0.098921f
C733 VP.n23 VSUBS 0.063157f
C734 VP.n24 VSUBS 0.063157f
C735 VP.n25 VSUBS 0.094916f
C736 VP.n26 VSUBS 0.039473f
C737 VP.n27 VSUBS 0.351682f
C738 VP.n28 VSUBS 2.26064f
C739 VP.n29 VSUBS 2.3197f
C740 VP.t4 VSUBS 0.578424f
C741 VP.n30 VSUBS 0.351682f
C742 VP.n31 VSUBS 0.039473f
C743 VP.n32 VSUBS 0.094916f
C744 VP.n33 VSUBS 0.063157f
C745 VP.n34 VSUBS 0.063157f
C746 VP.n35 VSUBS 0.098921f
C747 VP.n36 VSUBS 0.051242f
C748 VP.n37 VSUBS 0.097328f
C749 VP.n38 VSUBS 0.063157f
C750 VP.n39 VSUBS 0.063157f
C751 VP.n40 VSUBS 0.097328f
C752 VP.n41 VSUBS 0.051242f
C753 VP.n42 VSUBS 0.098921f
C754 VP.n43 VSUBS 0.063157f
C755 VP.n44 VSUBS 0.063157f
C756 VP.n45 VSUBS 0.094916f
C757 VP.n46 VSUBS 0.039473f
C758 VP.t2 VSUBS 0.578424f
C759 VP.n47 VSUBS 0.351682f
C760 VP.n48 VSUBS 0.059149f
.ends

