* NGSPICE file created from diff_pair_sample_1703.ext - technology: sky130A

.subckt diff_pair_sample_1703 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X1 VDD1.t9 VP.t0 VTAIL.t8 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X2 VTAIL.t9 VP.t1 VDD1.t8 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X3 VDD2.t2 VN.t1 VTAIL.t18 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=2.91
X4 B.t11 B.t9 B.t10 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=2.91
X5 VTAIL.t17 VN.t2 VDD2.t1 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X6 B.t8 B.t6 B.t7 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=2.91
X7 VDD1.t7 VP.t2 VTAIL.t7 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=2.91
X8 VDD2.t0 VN.t3 VTAIL.t16 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=2.91
X9 VTAIL.t15 VN.t4 VDD2.t5 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X10 B.t5 B.t3 B.t4 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=2.91
X11 VDD1.t6 VP.t3 VTAIL.t5 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X12 VTAIL.t14 VN.t5 VDD2.t4 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X13 VDD2.t9 VN.t6 VTAIL.t13 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=2.91
X14 VDD1.t5 VP.t4 VTAIL.t0 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=2.91
X15 VDD2.t8 VN.t7 VTAIL.t12 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=2.91
X16 VDD2.t7 VN.t8 VTAIL.t11 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X17 VTAIL.t6 VP.t5 VDD1.t4 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X18 VTAIL.t1 VP.t6 VDD1.t3 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X19 VTAIL.t4 VP.t7 VDD1.t2 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X20 VDD2.t6 VN.t9 VTAIL.t10 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=2.96505 ps=18.3 w=17.97 l=2.91
X21 VDD1.t1 VP.t8 VTAIL.t3 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=2.96505 ps=18.3 w=17.97 l=2.91
X22 B.t2 B.t0 B.t1 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=7.0083 pd=36.72 as=0 ps=0 w=17.97 l=2.91
X23 VDD1.t0 VP.t9 VTAIL.t2 w_n4858_n4562# sky130_fd_pr__pfet_01v8 ad=2.96505 pd=18.3 as=7.0083 ps=36.72 w=17.97 l=2.91
R0 VN.n54 VN.t3 180.657
R1 VN.n11 VN.t6 180.657
R2 VN.n84 VN.n83 161.3
R3 VN.n82 VN.n44 161.3
R4 VN.n81 VN.n80 161.3
R5 VN.n79 VN.n45 161.3
R6 VN.n78 VN.n77 161.3
R7 VN.n76 VN.n46 161.3
R8 VN.n74 VN.n73 161.3
R9 VN.n72 VN.n47 161.3
R10 VN.n71 VN.n70 161.3
R11 VN.n69 VN.n48 161.3
R12 VN.n68 VN.n67 161.3
R13 VN.n66 VN.n49 161.3
R14 VN.n65 VN.n64 161.3
R15 VN.n63 VN.n50 161.3
R16 VN.n62 VN.n61 161.3
R17 VN.n60 VN.n51 161.3
R18 VN.n59 VN.n58 161.3
R19 VN.n57 VN.n52 161.3
R20 VN.n56 VN.n55 161.3
R21 VN.n41 VN.n40 161.3
R22 VN.n39 VN.n1 161.3
R23 VN.n38 VN.n37 161.3
R24 VN.n36 VN.n2 161.3
R25 VN.n35 VN.n34 161.3
R26 VN.n33 VN.n3 161.3
R27 VN.n31 VN.n30 161.3
R28 VN.n29 VN.n4 161.3
R29 VN.n28 VN.n27 161.3
R30 VN.n26 VN.n5 161.3
R31 VN.n25 VN.n24 161.3
R32 VN.n23 VN.n6 161.3
R33 VN.n22 VN.n21 161.3
R34 VN.n20 VN.n7 161.3
R35 VN.n19 VN.n18 161.3
R36 VN.n17 VN.n8 161.3
R37 VN.n16 VN.n15 161.3
R38 VN.n14 VN.n9 161.3
R39 VN.n13 VN.n12 161.3
R40 VN.n21 VN.t8 148.825
R41 VN.n10 VN.t4 148.825
R42 VN.n32 VN.t5 148.825
R43 VN.n0 VN.t7 148.825
R44 VN.n64 VN.t9 148.825
R45 VN.n53 VN.t0 148.825
R46 VN.n75 VN.t2 148.825
R47 VN.n43 VN.t1 148.825
R48 VN.n42 VN.n0 66.5791
R49 VN.n85 VN.n43 66.5791
R50 VN.n11 VN.n10 62.0865
R51 VN.n54 VN.n53 62.0865
R52 VN VN.n85 59.642
R53 VN.n38 VN.n2 54.0911
R54 VN.n81 VN.n45 54.0911
R55 VN.n15 VN.n8 52.1486
R56 VN.n27 VN.n26 52.1486
R57 VN.n58 VN.n51 52.1486
R58 VN.n70 VN.n69 52.1486
R59 VN.n19 VN.n8 28.8382
R60 VN.n26 VN.n25 28.8382
R61 VN.n62 VN.n51 28.8382
R62 VN.n69 VN.n68 28.8382
R63 VN.n39 VN.n38 26.8957
R64 VN.n82 VN.n81 26.8957
R65 VN.n14 VN.n13 24.4675
R66 VN.n15 VN.n14 24.4675
R67 VN.n20 VN.n19 24.4675
R68 VN.n21 VN.n20 24.4675
R69 VN.n21 VN.n6 24.4675
R70 VN.n25 VN.n6 24.4675
R71 VN.n27 VN.n4 24.4675
R72 VN.n31 VN.n4 24.4675
R73 VN.n34 VN.n33 24.4675
R74 VN.n34 VN.n2 24.4675
R75 VN.n40 VN.n39 24.4675
R76 VN.n58 VN.n57 24.4675
R77 VN.n57 VN.n56 24.4675
R78 VN.n68 VN.n49 24.4675
R79 VN.n64 VN.n49 24.4675
R80 VN.n64 VN.n63 24.4675
R81 VN.n63 VN.n62 24.4675
R82 VN.n77 VN.n45 24.4675
R83 VN.n77 VN.n76 24.4675
R84 VN.n74 VN.n47 24.4675
R85 VN.n70 VN.n47 24.4675
R86 VN.n83 VN.n82 24.4675
R87 VN.n40 VN.n0 23.4888
R88 VN.n83 VN.n43 23.4888
R89 VN.n33 VN.n32 12.7233
R90 VN.n76 VN.n75 12.7233
R91 VN.n13 VN.n10 11.7447
R92 VN.n32 VN.n31 11.7447
R93 VN.n56 VN.n53 11.7447
R94 VN.n75 VN.n74 11.7447
R95 VN.n55 VN.n54 5.2926
R96 VN.n12 VN.n11 5.2926
R97 VN.n85 VN.n84 0.354971
R98 VN.n42 VN.n41 0.354971
R99 VN VN.n42 0.26696
R100 VN.n84 VN.n44 0.189894
R101 VN.n80 VN.n44 0.189894
R102 VN.n80 VN.n79 0.189894
R103 VN.n79 VN.n78 0.189894
R104 VN.n78 VN.n46 0.189894
R105 VN.n73 VN.n46 0.189894
R106 VN.n73 VN.n72 0.189894
R107 VN.n72 VN.n71 0.189894
R108 VN.n71 VN.n48 0.189894
R109 VN.n67 VN.n48 0.189894
R110 VN.n67 VN.n66 0.189894
R111 VN.n66 VN.n65 0.189894
R112 VN.n65 VN.n50 0.189894
R113 VN.n61 VN.n50 0.189894
R114 VN.n61 VN.n60 0.189894
R115 VN.n60 VN.n59 0.189894
R116 VN.n59 VN.n52 0.189894
R117 VN.n55 VN.n52 0.189894
R118 VN.n12 VN.n9 0.189894
R119 VN.n16 VN.n9 0.189894
R120 VN.n17 VN.n16 0.189894
R121 VN.n18 VN.n17 0.189894
R122 VN.n18 VN.n7 0.189894
R123 VN.n22 VN.n7 0.189894
R124 VN.n23 VN.n22 0.189894
R125 VN.n24 VN.n23 0.189894
R126 VN.n24 VN.n5 0.189894
R127 VN.n28 VN.n5 0.189894
R128 VN.n29 VN.n28 0.189894
R129 VN.n30 VN.n29 0.189894
R130 VN.n30 VN.n3 0.189894
R131 VN.n35 VN.n3 0.189894
R132 VN.n36 VN.n35 0.189894
R133 VN.n37 VN.n36 0.189894
R134 VN.n37 VN.n1 0.189894
R135 VN.n41 VN.n1 0.189894
R136 VDD2.n1 VDD2.t9 75.1978
R137 VDD2.n3 VDD2.n2 72.6354
R138 VDD2 VDD2.n7 72.6326
R139 VDD2.n4 VDD2.t2 72.405
R140 VDD2.n6 VDD2.n5 70.5961
R141 VDD2.n1 VDD2.n0 70.5959
R142 VDD2.n4 VDD2.n3 52.4739
R143 VDD2.n6 VDD2.n4 2.7936
R144 VDD2.n7 VDD2.t3 1.80935
R145 VDD2.n7 VDD2.t0 1.80935
R146 VDD2.n5 VDD2.t1 1.80935
R147 VDD2.n5 VDD2.t6 1.80935
R148 VDD2.n2 VDD2.t4 1.80935
R149 VDD2.n2 VDD2.t8 1.80935
R150 VDD2.n0 VDD2.t5 1.80935
R151 VDD2.n0 VDD2.t7 1.80935
R152 VDD2 VDD2.n6 0.756965
R153 VDD2.n3 VDD2.n1 0.64343
R154 VTAIL.n11 VTAIL.t16 55.7262
R155 VTAIL.n17 VTAIL.t12 55.726
R156 VTAIL.n2 VTAIL.t2 55.726
R157 VTAIL.n16 VTAIL.t0 55.726
R158 VTAIL.n15 VTAIL.n14 53.9174
R159 VTAIL.n13 VTAIL.n12 53.9174
R160 VTAIL.n10 VTAIL.n9 53.9174
R161 VTAIL.n8 VTAIL.n7 53.9174
R162 VTAIL.n19 VTAIL.n18 53.9171
R163 VTAIL.n1 VTAIL.n0 53.9171
R164 VTAIL.n4 VTAIL.n3 53.9171
R165 VTAIL.n6 VTAIL.n5 53.9171
R166 VTAIL.n8 VTAIL.n6 33.4445
R167 VTAIL.n17 VTAIL.n16 30.6514
R168 VTAIL.n10 VTAIL.n8 2.7936
R169 VTAIL.n11 VTAIL.n10 2.7936
R170 VTAIL.n15 VTAIL.n13 2.7936
R171 VTAIL.n16 VTAIL.n15 2.7936
R172 VTAIL.n6 VTAIL.n4 2.7936
R173 VTAIL.n4 VTAIL.n2 2.7936
R174 VTAIL.n19 VTAIL.n17 2.7936
R175 VTAIL VTAIL.n1 2.15352
R176 VTAIL.n13 VTAIL.n11 1.86688
R177 VTAIL.n2 VTAIL.n1 1.86688
R178 VTAIL.n18 VTAIL.t11 1.80935
R179 VTAIL.n18 VTAIL.t14 1.80935
R180 VTAIL.n0 VTAIL.t13 1.80935
R181 VTAIL.n0 VTAIL.t15 1.80935
R182 VTAIL.n3 VTAIL.t8 1.80935
R183 VTAIL.n3 VTAIL.t1 1.80935
R184 VTAIL.n5 VTAIL.t3 1.80935
R185 VTAIL.n5 VTAIL.t6 1.80935
R186 VTAIL.n14 VTAIL.t5 1.80935
R187 VTAIL.n14 VTAIL.t9 1.80935
R188 VTAIL.n12 VTAIL.t7 1.80935
R189 VTAIL.n12 VTAIL.t4 1.80935
R190 VTAIL.n9 VTAIL.t10 1.80935
R191 VTAIL.n9 VTAIL.t19 1.80935
R192 VTAIL.n7 VTAIL.t18 1.80935
R193 VTAIL.n7 VTAIL.t17 1.80935
R194 VTAIL VTAIL.n19 0.640586
R195 VP.n25 VP.t2 180.657
R196 VP.n27 VP.n26 161.3
R197 VP.n28 VP.n23 161.3
R198 VP.n30 VP.n29 161.3
R199 VP.n31 VP.n22 161.3
R200 VP.n33 VP.n32 161.3
R201 VP.n34 VP.n21 161.3
R202 VP.n36 VP.n35 161.3
R203 VP.n37 VP.n20 161.3
R204 VP.n39 VP.n38 161.3
R205 VP.n40 VP.n19 161.3
R206 VP.n42 VP.n41 161.3
R207 VP.n43 VP.n18 161.3
R208 VP.n45 VP.n44 161.3
R209 VP.n47 VP.n17 161.3
R210 VP.n49 VP.n48 161.3
R211 VP.n50 VP.n16 161.3
R212 VP.n52 VP.n51 161.3
R213 VP.n53 VP.n15 161.3
R214 VP.n55 VP.n54 161.3
R215 VP.n97 VP.n96 161.3
R216 VP.n95 VP.n1 161.3
R217 VP.n94 VP.n93 161.3
R218 VP.n92 VP.n2 161.3
R219 VP.n91 VP.n90 161.3
R220 VP.n89 VP.n3 161.3
R221 VP.n87 VP.n86 161.3
R222 VP.n85 VP.n4 161.3
R223 VP.n84 VP.n83 161.3
R224 VP.n82 VP.n5 161.3
R225 VP.n81 VP.n80 161.3
R226 VP.n79 VP.n6 161.3
R227 VP.n78 VP.n77 161.3
R228 VP.n76 VP.n7 161.3
R229 VP.n75 VP.n74 161.3
R230 VP.n73 VP.n8 161.3
R231 VP.n72 VP.n71 161.3
R232 VP.n70 VP.n9 161.3
R233 VP.n69 VP.n68 161.3
R234 VP.n67 VP.n66 161.3
R235 VP.n65 VP.n11 161.3
R236 VP.n64 VP.n63 161.3
R237 VP.n62 VP.n12 161.3
R238 VP.n61 VP.n60 161.3
R239 VP.n59 VP.n13 161.3
R240 VP.n77 VP.t0 148.825
R241 VP.n58 VP.t8 148.825
R242 VP.n10 VP.t5 148.825
R243 VP.n88 VP.t6 148.825
R244 VP.n0 VP.t9 148.825
R245 VP.n35 VP.t3 148.825
R246 VP.n14 VP.t4 148.825
R247 VP.n46 VP.t1 148.825
R248 VP.n24 VP.t7 148.825
R249 VP.n58 VP.n57 66.5791
R250 VP.n98 VP.n0 66.5791
R251 VP.n56 VP.n14 66.5791
R252 VP.n25 VP.n24 62.0865
R253 VP.n57 VP.n56 59.4766
R254 VP.n64 VP.n12 54.0911
R255 VP.n94 VP.n2 54.0911
R256 VP.n52 VP.n16 54.0911
R257 VP.n71 VP.n8 52.1486
R258 VP.n83 VP.n82 52.1486
R259 VP.n41 VP.n40 52.1486
R260 VP.n29 VP.n22 52.1486
R261 VP.n75 VP.n8 28.8382
R262 VP.n82 VP.n81 28.8382
R263 VP.n40 VP.n39 28.8382
R264 VP.n33 VP.n22 28.8382
R265 VP.n60 VP.n12 26.8957
R266 VP.n95 VP.n94 26.8957
R267 VP.n53 VP.n52 26.8957
R268 VP.n60 VP.n59 24.4675
R269 VP.n65 VP.n64 24.4675
R270 VP.n66 VP.n65 24.4675
R271 VP.n70 VP.n69 24.4675
R272 VP.n71 VP.n70 24.4675
R273 VP.n76 VP.n75 24.4675
R274 VP.n77 VP.n76 24.4675
R275 VP.n77 VP.n6 24.4675
R276 VP.n81 VP.n6 24.4675
R277 VP.n83 VP.n4 24.4675
R278 VP.n87 VP.n4 24.4675
R279 VP.n90 VP.n89 24.4675
R280 VP.n90 VP.n2 24.4675
R281 VP.n96 VP.n95 24.4675
R282 VP.n54 VP.n53 24.4675
R283 VP.n41 VP.n18 24.4675
R284 VP.n45 VP.n18 24.4675
R285 VP.n48 VP.n47 24.4675
R286 VP.n48 VP.n16 24.4675
R287 VP.n34 VP.n33 24.4675
R288 VP.n35 VP.n34 24.4675
R289 VP.n35 VP.n20 24.4675
R290 VP.n39 VP.n20 24.4675
R291 VP.n28 VP.n27 24.4675
R292 VP.n29 VP.n28 24.4675
R293 VP.n59 VP.n58 23.4888
R294 VP.n96 VP.n0 23.4888
R295 VP.n54 VP.n14 23.4888
R296 VP.n66 VP.n10 12.7233
R297 VP.n89 VP.n88 12.7233
R298 VP.n47 VP.n46 12.7233
R299 VP.n69 VP.n10 11.7447
R300 VP.n88 VP.n87 11.7447
R301 VP.n46 VP.n45 11.7447
R302 VP.n27 VP.n24 11.7447
R303 VP.n26 VP.n25 5.29256
R304 VP.n56 VP.n55 0.354971
R305 VP.n57 VP.n13 0.354971
R306 VP.n98 VP.n97 0.354971
R307 VP VP.n98 0.26696
R308 VP.n26 VP.n23 0.189894
R309 VP.n30 VP.n23 0.189894
R310 VP.n31 VP.n30 0.189894
R311 VP.n32 VP.n31 0.189894
R312 VP.n32 VP.n21 0.189894
R313 VP.n36 VP.n21 0.189894
R314 VP.n37 VP.n36 0.189894
R315 VP.n38 VP.n37 0.189894
R316 VP.n38 VP.n19 0.189894
R317 VP.n42 VP.n19 0.189894
R318 VP.n43 VP.n42 0.189894
R319 VP.n44 VP.n43 0.189894
R320 VP.n44 VP.n17 0.189894
R321 VP.n49 VP.n17 0.189894
R322 VP.n50 VP.n49 0.189894
R323 VP.n51 VP.n50 0.189894
R324 VP.n51 VP.n15 0.189894
R325 VP.n55 VP.n15 0.189894
R326 VP.n61 VP.n13 0.189894
R327 VP.n62 VP.n61 0.189894
R328 VP.n63 VP.n62 0.189894
R329 VP.n63 VP.n11 0.189894
R330 VP.n67 VP.n11 0.189894
R331 VP.n68 VP.n67 0.189894
R332 VP.n68 VP.n9 0.189894
R333 VP.n72 VP.n9 0.189894
R334 VP.n73 VP.n72 0.189894
R335 VP.n74 VP.n73 0.189894
R336 VP.n74 VP.n7 0.189894
R337 VP.n78 VP.n7 0.189894
R338 VP.n79 VP.n78 0.189894
R339 VP.n80 VP.n79 0.189894
R340 VP.n80 VP.n5 0.189894
R341 VP.n84 VP.n5 0.189894
R342 VP.n85 VP.n84 0.189894
R343 VP.n86 VP.n85 0.189894
R344 VP.n86 VP.n3 0.189894
R345 VP.n91 VP.n3 0.189894
R346 VP.n92 VP.n91 0.189894
R347 VP.n93 VP.n92 0.189894
R348 VP.n93 VP.n1 0.189894
R349 VP.n97 VP.n1 0.189894
R350 VDD1.n1 VDD1.t7 75.1981
R351 VDD1.n3 VDD1.t1 75.1978
R352 VDD1.n5 VDD1.n4 72.6354
R353 VDD1.n1 VDD1.n0 70.5961
R354 VDD1.n7 VDD1.n6 70.596
R355 VDD1.n3 VDD1.n2 70.5959
R356 VDD1.n7 VDD1.n5 54.4535
R357 VDD1 VDD1.n7 2.03714
R358 VDD1.n6 VDD1.t8 1.80935
R359 VDD1.n6 VDD1.t5 1.80935
R360 VDD1.n0 VDD1.t2 1.80935
R361 VDD1.n0 VDD1.t6 1.80935
R362 VDD1.n4 VDD1.t3 1.80935
R363 VDD1.n4 VDD1.t0 1.80935
R364 VDD1.n2 VDD1.t4 1.80935
R365 VDD1.n2 VDD1.t9 1.80935
R366 VDD1 VDD1.n1 0.756965
R367 VDD1.n5 VDD1.n3 0.64343
R368 B.n558 B.n169 585
R369 B.n557 B.n556 585
R370 B.n555 B.n170 585
R371 B.n554 B.n553 585
R372 B.n552 B.n171 585
R373 B.n551 B.n550 585
R374 B.n549 B.n172 585
R375 B.n548 B.n547 585
R376 B.n546 B.n173 585
R377 B.n545 B.n544 585
R378 B.n543 B.n174 585
R379 B.n542 B.n541 585
R380 B.n540 B.n175 585
R381 B.n539 B.n538 585
R382 B.n537 B.n176 585
R383 B.n536 B.n535 585
R384 B.n534 B.n177 585
R385 B.n533 B.n532 585
R386 B.n531 B.n178 585
R387 B.n530 B.n529 585
R388 B.n528 B.n179 585
R389 B.n527 B.n526 585
R390 B.n525 B.n180 585
R391 B.n524 B.n523 585
R392 B.n522 B.n181 585
R393 B.n521 B.n520 585
R394 B.n519 B.n182 585
R395 B.n518 B.n517 585
R396 B.n516 B.n183 585
R397 B.n515 B.n514 585
R398 B.n513 B.n184 585
R399 B.n512 B.n511 585
R400 B.n510 B.n185 585
R401 B.n509 B.n508 585
R402 B.n507 B.n186 585
R403 B.n506 B.n505 585
R404 B.n504 B.n187 585
R405 B.n503 B.n502 585
R406 B.n501 B.n188 585
R407 B.n500 B.n499 585
R408 B.n498 B.n189 585
R409 B.n497 B.n496 585
R410 B.n495 B.n190 585
R411 B.n494 B.n493 585
R412 B.n492 B.n191 585
R413 B.n491 B.n490 585
R414 B.n489 B.n192 585
R415 B.n488 B.n487 585
R416 B.n486 B.n193 585
R417 B.n485 B.n484 585
R418 B.n483 B.n194 585
R419 B.n482 B.n481 585
R420 B.n480 B.n195 585
R421 B.n479 B.n478 585
R422 B.n477 B.n196 585
R423 B.n476 B.n475 585
R424 B.n474 B.n197 585
R425 B.n473 B.n472 585
R426 B.n471 B.n198 585
R427 B.n470 B.n469 585
R428 B.n465 B.n199 585
R429 B.n464 B.n463 585
R430 B.n462 B.n200 585
R431 B.n461 B.n460 585
R432 B.n459 B.n201 585
R433 B.n458 B.n457 585
R434 B.n456 B.n202 585
R435 B.n455 B.n454 585
R436 B.n453 B.n203 585
R437 B.n451 B.n450 585
R438 B.n449 B.n206 585
R439 B.n448 B.n447 585
R440 B.n446 B.n207 585
R441 B.n445 B.n444 585
R442 B.n443 B.n208 585
R443 B.n442 B.n441 585
R444 B.n440 B.n209 585
R445 B.n439 B.n438 585
R446 B.n437 B.n210 585
R447 B.n436 B.n435 585
R448 B.n434 B.n211 585
R449 B.n433 B.n432 585
R450 B.n431 B.n212 585
R451 B.n430 B.n429 585
R452 B.n428 B.n213 585
R453 B.n427 B.n426 585
R454 B.n425 B.n214 585
R455 B.n424 B.n423 585
R456 B.n422 B.n215 585
R457 B.n421 B.n420 585
R458 B.n419 B.n216 585
R459 B.n418 B.n417 585
R460 B.n416 B.n217 585
R461 B.n415 B.n414 585
R462 B.n413 B.n218 585
R463 B.n412 B.n411 585
R464 B.n410 B.n219 585
R465 B.n409 B.n408 585
R466 B.n407 B.n220 585
R467 B.n406 B.n405 585
R468 B.n404 B.n221 585
R469 B.n403 B.n402 585
R470 B.n401 B.n222 585
R471 B.n400 B.n399 585
R472 B.n398 B.n223 585
R473 B.n397 B.n396 585
R474 B.n395 B.n224 585
R475 B.n394 B.n393 585
R476 B.n392 B.n225 585
R477 B.n391 B.n390 585
R478 B.n389 B.n226 585
R479 B.n388 B.n387 585
R480 B.n386 B.n227 585
R481 B.n385 B.n384 585
R482 B.n383 B.n228 585
R483 B.n382 B.n381 585
R484 B.n380 B.n229 585
R485 B.n379 B.n378 585
R486 B.n377 B.n230 585
R487 B.n376 B.n375 585
R488 B.n374 B.n231 585
R489 B.n373 B.n372 585
R490 B.n371 B.n232 585
R491 B.n370 B.n369 585
R492 B.n368 B.n233 585
R493 B.n367 B.n366 585
R494 B.n365 B.n234 585
R495 B.n364 B.n363 585
R496 B.n560 B.n559 585
R497 B.n561 B.n168 585
R498 B.n563 B.n562 585
R499 B.n564 B.n167 585
R500 B.n566 B.n565 585
R501 B.n567 B.n166 585
R502 B.n569 B.n568 585
R503 B.n570 B.n165 585
R504 B.n572 B.n571 585
R505 B.n573 B.n164 585
R506 B.n575 B.n574 585
R507 B.n576 B.n163 585
R508 B.n578 B.n577 585
R509 B.n579 B.n162 585
R510 B.n581 B.n580 585
R511 B.n582 B.n161 585
R512 B.n584 B.n583 585
R513 B.n585 B.n160 585
R514 B.n587 B.n586 585
R515 B.n588 B.n159 585
R516 B.n590 B.n589 585
R517 B.n591 B.n158 585
R518 B.n593 B.n592 585
R519 B.n594 B.n157 585
R520 B.n596 B.n595 585
R521 B.n597 B.n156 585
R522 B.n599 B.n598 585
R523 B.n600 B.n155 585
R524 B.n602 B.n601 585
R525 B.n603 B.n154 585
R526 B.n605 B.n604 585
R527 B.n606 B.n153 585
R528 B.n608 B.n607 585
R529 B.n609 B.n152 585
R530 B.n611 B.n610 585
R531 B.n612 B.n151 585
R532 B.n614 B.n613 585
R533 B.n615 B.n150 585
R534 B.n617 B.n616 585
R535 B.n618 B.n149 585
R536 B.n620 B.n619 585
R537 B.n621 B.n148 585
R538 B.n623 B.n622 585
R539 B.n624 B.n147 585
R540 B.n626 B.n625 585
R541 B.n627 B.n146 585
R542 B.n629 B.n628 585
R543 B.n630 B.n145 585
R544 B.n632 B.n631 585
R545 B.n633 B.n144 585
R546 B.n635 B.n634 585
R547 B.n636 B.n143 585
R548 B.n638 B.n637 585
R549 B.n639 B.n142 585
R550 B.n641 B.n640 585
R551 B.n642 B.n141 585
R552 B.n644 B.n643 585
R553 B.n645 B.n140 585
R554 B.n647 B.n646 585
R555 B.n648 B.n139 585
R556 B.n650 B.n649 585
R557 B.n651 B.n138 585
R558 B.n653 B.n652 585
R559 B.n654 B.n137 585
R560 B.n656 B.n655 585
R561 B.n657 B.n136 585
R562 B.n659 B.n658 585
R563 B.n660 B.n135 585
R564 B.n662 B.n661 585
R565 B.n663 B.n134 585
R566 B.n665 B.n664 585
R567 B.n666 B.n133 585
R568 B.n668 B.n667 585
R569 B.n669 B.n132 585
R570 B.n671 B.n670 585
R571 B.n672 B.n131 585
R572 B.n674 B.n673 585
R573 B.n675 B.n130 585
R574 B.n677 B.n676 585
R575 B.n678 B.n129 585
R576 B.n680 B.n679 585
R577 B.n681 B.n128 585
R578 B.n683 B.n682 585
R579 B.n684 B.n127 585
R580 B.n686 B.n685 585
R581 B.n687 B.n126 585
R582 B.n689 B.n688 585
R583 B.n690 B.n125 585
R584 B.n692 B.n691 585
R585 B.n693 B.n124 585
R586 B.n695 B.n694 585
R587 B.n696 B.n123 585
R588 B.n698 B.n697 585
R589 B.n699 B.n122 585
R590 B.n701 B.n700 585
R591 B.n702 B.n121 585
R592 B.n704 B.n703 585
R593 B.n705 B.n120 585
R594 B.n707 B.n706 585
R595 B.n708 B.n119 585
R596 B.n710 B.n709 585
R597 B.n711 B.n118 585
R598 B.n713 B.n712 585
R599 B.n714 B.n117 585
R600 B.n716 B.n715 585
R601 B.n717 B.n116 585
R602 B.n719 B.n718 585
R603 B.n720 B.n115 585
R604 B.n722 B.n721 585
R605 B.n723 B.n114 585
R606 B.n725 B.n724 585
R607 B.n726 B.n113 585
R608 B.n728 B.n727 585
R609 B.n729 B.n112 585
R610 B.n731 B.n730 585
R611 B.n732 B.n111 585
R612 B.n734 B.n733 585
R613 B.n735 B.n110 585
R614 B.n737 B.n736 585
R615 B.n738 B.n109 585
R616 B.n740 B.n739 585
R617 B.n741 B.n108 585
R618 B.n743 B.n742 585
R619 B.n744 B.n107 585
R620 B.n746 B.n745 585
R621 B.n747 B.n106 585
R622 B.n749 B.n748 585
R623 B.n750 B.n105 585
R624 B.n752 B.n751 585
R625 B.n753 B.n104 585
R626 B.n755 B.n754 585
R627 B.n756 B.n103 585
R628 B.n950 B.n949 585
R629 B.n948 B.n35 585
R630 B.n947 B.n946 585
R631 B.n945 B.n36 585
R632 B.n944 B.n943 585
R633 B.n942 B.n37 585
R634 B.n941 B.n940 585
R635 B.n939 B.n38 585
R636 B.n938 B.n937 585
R637 B.n936 B.n39 585
R638 B.n935 B.n934 585
R639 B.n933 B.n40 585
R640 B.n932 B.n931 585
R641 B.n930 B.n41 585
R642 B.n929 B.n928 585
R643 B.n927 B.n42 585
R644 B.n926 B.n925 585
R645 B.n924 B.n43 585
R646 B.n923 B.n922 585
R647 B.n921 B.n44 585
R648 B.n920 B.n919 585
R649 B.n918 B.n45 585
R650 B.n917 B.n916 585
R651 B.n915 B.n46 585
R652 B.n914 B.n913 585
R653 B.n912 B.n47 585
R654 B.n911 B.n910 585
R655 B.n909 B.n48 585
R656 B.n908 B.n907 585
R657 B.n906 B.n49 585
R658 B.n905 B.n904 585
R659 B.n903 B.n50 585
R660 B.n902 B.n901 585
R661 B.n900 B.n51 585
R662 B.n899 B.n898 585
R663 B.n897 B.n52 585
R664 B.n896 B.n895 585
R665 B.n894 B.n53 585
R666 B.n893 B.n892 585
R667 B.n891 B.n54 585
R668 B.n890 B.n889 585
R669 B.n888 B.n55 585
R670 B.n887 B.n886 585
R671 B.n885 B.n56 585
R672 B.n884 B.n883 585
R673 B.n882 B.n57 585
R674 B.n881 B.n880 585
R675 B.n879 B.n58 585
R676 B.n878 B.n877 585
R677 B.n876 B.n59 585
R678 B.n875 B.n874 585
R679 B.n873 B.n60 585
R680 B.n872 B.n871 585
R681 B.n870 B.n61 585
R682 B.n869 B.n868 585
R683 B.n867 B.n62 585
R684 B.n866 B.n865 585
R685 B.n864 B.n63 585
R686 B.n863 B.n862 585
R687 B.n861 B.n860 585
R688 B.n859 B.n67 585
R689 B.n858 B.n857 585
R690 B.n856 B.n68 585
R691 B.n855 B.n854 585
R692 B.n853 B.n69 585
R693 B.n852 B.n851 585
R694 B.n850 B.n70 585
R695 B.n849 B.n848 585
R696 B.n847 B.n71 585
R697 B.n845 B.n844 585
R698 B.n843 B.n74 585
R699 B.n842 B.n841 585
R700 B.n840 B.n75 585
R701 B.n839 B.n838 585
R702 B.n837 B.n76 585
R703 B.n836 B.n835 585
R704 B.n834 B.n77 585
R705 B.n833 B.n832 585
R706 B.n831 B.n78 585
R707 B.n830 B.n829 585
R708 B.n828 B.n79 585
R709 B.n827 B.n826 585
R710 B.n825 B.n80 585
R711 B.n824 B.n823 585
R712 B.n822 B.n81 585
R713 B.n821 B.n820 585
R714 B.n819 B.n82 585
R715 B.n818 B.n817 585
R716 B.n816 B.n83 585
R717 B.n815 B.n814 585
R718 B.n813 B.n84 585
R719 B.n812 B.n811 585
R720 B.n810 B.n85 585
R721 B.n809 B.n808 585
R722 B.n807 B.n86 585
R723 B.n806 B.n805 585
R724 B.n804 B.n87 585
R725 B.n803 B.n802 585
R726 B.n801 B.n88 585
R727 B.n800 B.n799 585
R728 B.n798 B.n89 585
R729 B.n797 B.n796 585
R730 B.n795 B.n90 585
R731 B.n794 B.n793 585
R732 B.n792 B.n91 585
R733 B.n791 B.n790 585
R734 B.n789 B.n92 585
R735 B.n788 B.n787 585
R736 B.n786 B.n93 585
R737 B.n785 B.n784 585
R738 B.n783 B.n94 585
R739 B.n782 B.n781 585
R740 B.n780 B.n95 585
R741 B.n779 B.n778 585
R742 B.n777 B.n96 585
R743 B.n776 B.n775 585
R744 B.n774 B.n97 585
R745 B.n773 B.n772 585
R746 B.n771 B.n98 585
R747 B.n770 B.n769 585
R748 B.n768 B.n99 585
R749 B.n767 B.n766 585
R750 B.n765 B.n100 585
R751 B.n764 B.n763 585
R752 B.n762 B.n101 585
R753 B.n761 B.n760 585
R754 B.n759 B.n102 585
R755 B.n758 B.n757 585
R756 B.n951 B.n34 585
R757 B.n953 B.n952 585
R758 B.n954 B.n33 585
R759 B.n956 B.n955 585
R760 B.n957 B.n32 585
R761 B.n959 B.n958 585
R762 B.n960 B.n31 585
R763 B.n962 B.n961 585
R764 B.n963 B.n30 585
R765 B.n965 B.n964 585
R766 B.n966 B.n29 585
R767 B.n968 B.n967 585
R768 B.n969 B.n28 585
R769 B.n971 B.n970 585
R770 B.n972 B.n27 585
R771 B.n974 B.n973 585
R772 B.n975 B.n26 585
R773 B.n977 B.n976 585
R774 B.n978 B.n25 585
R775 B.n980 B.n979 585
R776 B.n981 B.n24 585
R777 B.n983 B.n982 585
R778 B.n984 B.n23 585
R779 B.n986 B.n985 585
R780 B.n987 B.n22 585
R781 B.n989 B.n988 585
R782 B.n990 B.n21 585
R783 B.n992 B.n991 585
R784 B.n993 B.n20 585
R785 B.n995 B.n994 585
R786 B.n996 B.n19 585
R787 B.n998 B.n997 585
R788 B.n999 B.n18 585
R789 B.n1001 B.n1000 585
R790 B.n1002 B.n17 585
R791 B.n1004 B.n1003 585
R792 B.n1005 B.n16 585
R793 B.n1007 B.n1006 585
R794 B.n1008 B.n15 585
R795 B.n1010 B.n1009 585
R796 B.n1011 B.n14 585
R797 B.n1013 B.n1012 585
R798 B.n1014 B.n13 585
R799 B.n1016 B.n1015 585
R800 B.n1017 B.n12 585
R801 B.n1019 B.n1018 585
R802 B.n1020 B.n11 585
R803 B.n1022 B.n1021 585
R804 B.n1023 B.n10 585
R805 B.n1025 B.n1024 585
R806 B.n1026 B.n9 585
R807 B.n1028 B.n1027 585
R808 B.n1029 B.n8 585
R809 B.n1031 B.n1030 585
R810 B.n1032 B.n7 585
R811 B.n1034 B.n1033 585
R812 B.n1035 B.n6 585
R813 B.n1037 B.n1036 585
R814 B.n1038 B.n5 585
R815 B.n1040 B.n1039 585
R816 B.n1041 B.n4 585
R817 B.n1043 B.n1042 585
R818 B.n1044 B.n3 585
R819 B.n1046 B.n1045 585
R820 B.n1047 B.n0 585
R821 B.n2 B.n1 585
R822 B.n268 B.n267 585
R823 B.n269 B.n266 585
R824 B.n271 B.n270 585
R825 B.n272 B.n265 585
R826 B.n274 B.n273 585
R827 B.n275 B.n264 585
R828 B.n277 B.n276 585
R829 B.n278 B.n263 585
R830 B.n280 B.n279 585
R831 B.n281 B.n262 585
R832 B.n283 B.n282 585
R833 B.n284 B.n261 585
R834 B.n286 B.n285 585
R835 B.n287 B.n260 585
R836 B.n289 B.n288 585
R837 B.n290 B.n259 585
R838 B.n292 B.n291 585
R839 B.n293 B.n258 585
R840 B.n295 B.n294 585
R841 B.n296 B.n257 585
R842 B.n298 B.n297 585
R843 B.n299 B.n256 585
R844 B.n301 B.n300 585
R845 B.n302 B.n255 585
R846 B.n304 B.n303 585
R847 B.n305 B.n254 585
R848 B.n307 B.n306 585
R849 B.n308 B.n253 585
R850 B.n310 B.n309 585
R851 B.n311 B.n252 585
R852 B.n313 B.n312 585
R853 B.n314 B.n251 585
R854 B.n316 B.n315 585
R855 B.n317 B.n250 585
R856 B.n319 B.n318 585
R857 B.n320 B.n249 585
R858 B.n322 B.n321 585
R859 B.n323 B.n248 585
R860 B.n325 B.n324 585
R861 B.n326 B.n247 585
R862 B.n328 B.n327 585
R863 B.n329 B.n246 585
R864 B.n331 B.n330 585
R865 B.n332 B.n245 585
R866 B.n334 B.n333 585
R867 B.n335 B.n244 585
R868 B.n337 B.n336 585
R869 B.n338 B.n243 585
R870 B.n340 B.n339 585
R871 B.n341 B.n242 585
R872 B.n343 B.n342 585
R873 B.n344 B.n241 585
R874 B.n346 B.n345 585
R875 B.n347 B.n240 585
R876 B.n349 B.n348 585
R877 B.n350 B.n239 585
R878 B.n352 B.n351 585
R879 B.n353 B.n238 585
R880 B.n355 B.n354 585
R881 B.n356 B.n237 585
R882 B.n358 B.n357 585
R883 B.n359 B.n236 585
R884 B.n361 B.n360 585
R885 B.n362 B.n235 585
R886 B.n364 B.n235 458.866
R887 B.n560 B.n169 458.866
R888 B.n758 B.n103 458.866
R889 B.n951 B.n950 458.866
R890 B.n204 B.t3 357.296
R891 B.n466 B.t6 357.296
R892 B.n72 B.t0 357.296
R893 B.n64 B.t9 357.296
R894 B.n1049 B.n1048 256.663
R895 B.n1048 B.n1047 235.042
R896 B.n1048 B.n2 235.042
R897 B.n466 B.t7 174.667
R898 B.n72 B.t2 174.667
R899 B.n204 B.t4 174.644
R900 B.n64 B.t11 174.644
R901 B.n365 B.n364 163.367
R902 B.n366 B.n365 163.367
R903 B.n366 B.n233 163.367
R904 B.n370 B.n233 163.367
R905 B.n371 B.n370 163.367
R906 B.n372 B.n371 163.367
R907 B.n372 B.n231 163.367
R908 B.n376 B.n231 163.367
R909 B.n377 B.n376 163.367
R910 B.n378 B.n377 163.367
R911 B.n378 B.n229 163.367
R912 B.n382 B.n229 163.367
R913 B.n383 B.n382 163.367
R914 B.n384 B.n383 163.367
R915 B.n384 B.n227 163.367
R916 B.n388 B.n227 163.367
R917 B.n389 B.n388 163.367
R918 B.n390 B.n389 163.367
R919 B.n390 B.n225 163.367
R920 B.n394 B.n225 163.367
R921 B.n395 B.n394 163.367
R922 B.n396 B.n395 163.367
R923 B.n396 B.n223 163.367
R924 B.n400 B.n223 163.367
R925 B.n401 B.n400 163.367
R926 B.n402 B.n401 163.367
R927 B.n402 B.n221 163.367
R928 B.n406 B.n221 163.367
R929 B.n407 B.n406 163.367
R930 B.n408 B.n407 163.367
R931 B.n408 B.n219 163.367
R932 B.n412 B.n219 163.367
R933 B.n413 B.n412 163.367
R934 B.n414 B.n413 163.367
R935 B.n414 B.n217 163.367
R936 B.n418 B.n217 163.367
R937 B.n419 B.n418 163.367
R938 B.n420 B.n419 163.367
R939 B.n420 B.n215 163.367
R940 B.n424 B.n215 163.367
R941 B.n425 B.n424 163.367
R942 B.n426 B.n425 163.367
R943 B.n426 B.n213 163.367
R944 B.n430 B.n213 163.367
R945 B.n431 B.n430 163.367
R946 B.n432 B.n431 163.367
R947 B.n432 B.n211 163.367
R948 B.n436 B.n211 163.367
R949 B.n437 B.n436 163.367
R950 B.n438 B.n437 163.367
R951 B.n438 B.n209 163.367
R952 B.n442 B.n209 163.367
R953 B.n443 B.n442 163.367
R954 B.n444 B.n443 163.367
R955 B.n444 B.n207 163.367
R956 B.n448 B.n207 163.367
R957 B.n449 B.n448 163.367
R958 B.n450 B.n449 163.367
R959 B.n450 B.n203 163.367
R960 B.n455 B.n203 163.367
R961 B.n456 B.n455 163.367
R962 B.n457 B.n456 163.367
R963 B.n457 B.n201 163.367
R964 B.n461 B.n201 163.367
R965 B.n462 B.n461 163.367
R966 B.n463 B.n462 163.367
R967 B.n463 B.n199 163.367
R968 B.n470 B.n199 163.367
R969 B.n471 B.n470 163.367
R970 B.n472 B.n471 163.367
R971 B.n472 B.n197 163.367
R972 B.n476 B.n197 163.367
R973 B.n477 B.n476 163.367
R974 B.n478 B.n477 163.367
R975 B.n478 B.n195 163.367
R976 B.n482 B.n195 163.367
R977 B.n483 B.n482 163.367
R978 B.n484 B.n483 163.367
R979 B.n484 B.n193 163.367
R980 B.n488 B.n193 163.367
R981 B.n489 B.n488 163.367
R982 B.n490 B.n489 163.367
R983 B.n490 B.n191 163.367
R984 B.n494 B.n191 163.367
R985 B.n495 B.n494 163.367
R986 B.n496 B.n495 163.367
R987 B.n496 B.n189 163.367
R988 B.n500 B.n189 163.367
R989 B.n501 B.n500 163.367
R990 B.n502 B.n501 163.367
R991 B.n502 B.n187 163.367
R992 B.n506 B.n187 163.367
R993 B.n507 B.n506 163.367
R994 B.n508 B.n507 163.367
R995 B.n508 B.n185 163.367
R996 B.n512 B.n185 163.367
R997 B.n513 B.n512 163.367
R998 B.n514 B.n513 163.367
R999 B.n514 B.n183 163.367
R1000 B.n518 B.n183 163.367
R1001 B.n519 B.n518 163.367
R1002 B.n520 B.n519 163.367
R1003 B.n520 B.n181 163.367
R1004 B.n524 B.n181 163.367
R1005 B.n525 B.n524 163.367
R1006 B.n526 B.n525 163.367
R1007 B.n526 B.n179 163.367
R1008 B.n530 B.n179 163.367
R1009 B.n531 B.n530 163.367
R1010 B.n532 B.n531 163.367
R1011 B.n532 B.n177 163.367
R1012 B.n536 B.n177 163.367
R1013 B.n537 B.n536 163.367
R1014 B.n538 B.n537 163.367
R1015 B.n538 B.n175 163.367
R1016 B.n542 B.n175 163.367
R1017 B.n543 B.n542 163.367
R1018 B.n544 B.n543 163.367
R1019 B.n544 B.n173 163.367
R1020 B.n548 B.n173 163.367
R1021 B.n549 B.n548 163.367
R1022 B.n550 B.n549 163.367
R1023 B.n550 B.n171 163.367
R1024 B.n554 B.n171 163.367
R1025 B.n555 B.n554 163.367
R1026 B.n556 B.n555 163.367
R1027 B.n556 B.n169 163.367
R1028 B.n754 B.n103 163.367
R1029 B.n754 B.n753 163.367
R1030 B.n753 B.n752 163.367
R1031 B.n752 B.n105 163.367
R1032 B.n748 B.n105 163.367
R1033 B.n748 B.n747 163.367
R1034 B.n747 B.n746 163.367
R1035 B.n746 B.n107 163.367
R1036 B.n742 B.n107 163.367
R1037 B.n742 B.n741 163.367
R1038 B.n741 B.n740 163.367
R1039 B.n740 B.n109 163.367
R1040 B.n736 B.n109 163.367
R1041 B.n736 B.n735 163.367
R1042 B.n735 B.n734 163.367
R1043 B.n734 B.n111 163.367
R1044 B.n730 B.n111 163.367
R1045 B.n730 B.n729 163.367
R1046 B.n729 B.n728 163.367
R1047 B.n728 B.n113 163.367
R1048 B.n724 B.n113 163.367
R1049 B.n724 B.n723 163.367
R1050 B.n723 B.n722 163.367
R1051 B.n722 B.n115 163.367
R1052 B.n718 B.n115 163.367
R1053 B.n718 B.n717 163.367
R1054 B.n717 B.n716 163.367
R1055 B.n716 B.n117 163.367
R1056 B.n712 B.n117 163.367
R1057 B.n712 B.n711 163.367
R1058 B.n711 B.n710 163.367
R1059 B.n710 B.n119 163.367
R1060 B.n706 B.n119 163.367
R1061 B.n706 B.n705 163.367
R1062 B.n705 B.n704 163.367
R1063 B.n704 B.n121 163.367
R1064 B.n700 B.n121 163.367
R1065 B.n700 B.n699 163.367
R1066 B.n699 B.n698 163.367
R1067 B.n698 B.n123 163.367
R1068 B.n694 B.n123 163.367
R1069 B.n694 B.n693 163.367
R1070 B.n693 B.n692 163.367
R1071 B.n692 B.n125 163.367
R1072 B.n688 B.n125 163.367
R1073 B.n688 B.n687 163.367
R1074 B.n687 B.n686 163.367
R1075 B.n686 B.n127 163.367
R1076 B.n682 B.n127 163.367
R1077 B.n682 B.n681 163.367
R1078 B.n681 B.n680 163.367
R1079 B.n680 B.n129 163.367
R1080 B.n676 B.n129 163.367
R1081 B.n676 B.n675 163.367
R1082 B.n675 B.n674 163.367
R1083 B.n674 B.n131 163.367
R1084 B.n670 B.n131 163.367
R1085 B.n670 B.n669 163.367
R1086 B.n669 B.n668 163.367
R1087 B.n668 B.n133 163.367
R1088 B.n664 B.n133 163.367
R1089 B.n664 B.n663 163.367
R1090 B.n663 B.n662 163.367
R1091 B.n662 B.n135 163.367
R1092 B.n658 B.n135 163.367
R1093 B.n658 B.n657 163.367
R1094 B.n657 B.n656 163.367
R1095 B.n656 B.n137 163.367
R1096 B.n652 B.n137 163.367
R1097 B.n652 B.n651 163.367
R1098 B.n651 B.n650 163.367
R1099 B.n650 B.n139 163.367
R1100 B.n646 B.n139 163.367
R1101 B.n646 B.n645 163.367
R1102 B.n645 B.n644 163.367
R1103 B.n644 B.n141 163.367
R1104 B.n640 B.n141 163.367
R1105 B.n640 B.n639 163.367
R1106 B.n639 B.n638 163.367
R1107 B.n638 B.n143 163.367
R1108 B.n634 B.n143 163.367
R1109 B.n634 B.n633 163.367
R1110 B.n633 B.n632 163.367
R1111 B.n632 B.n145 163.367
R1112 B.n628 B.n145 163.367
R1113 B.n628 B.n627 163.367
R1114 B.n627 B.n626 163.367
R1115 B.n626 B.n147 163.367
R1116 B.n622 B.n147 163.367
R1117 B.n622 B.n621 163.367
R1118 B.n621 B.n620 163.367
R1119 B.n620 B.n149 163.367
R1120 B.n616 B.n149 163.367
R1121 B.n616 B.n615 163.367
R1122 B.n615 B.n614 163.367
R1123 B.n614 B.n151 163.367
R1124 B.n610 B.n151 163.367
R1125 B.n610 B.n609 163.367
R1126 B.n609 B.n608 163.367
R1127 B.n608 B.n153 163.367
R1128 B.n604 B.n153 163.367
R1129 B.n604 B.n603 163.367
R1130 B.n603 B.n602 163.367
R1131 B.n602 B.n155 163.367
R1132 B.n598 B.n155 163.367
R1133 B.n598 B.n597 163.367
R1134 B.n597 B.n596 163.367
R1135 B.n596 B.n157 163.367
R1136 B.n592 B.n157 163.367
R1137 B.n592 B.n591 163.367
R1138 B.n591 B.n590 163.367
R1139 B.n590 B.n159 163.367
R1140 B.n586 B.n159 163.367
R1141 B.n586 B.n585 163.367
R1142 B.n585 B.n584 163.367
R1143 B.n584 B.n161 163.367
R1144 B.n580 B.n161 163.367
R1145 B.n580 B.n579 163.367
R1146 B.n579 B.n578 163.367
R1147 B.n578 B.n163 163.367
R1148 B.n574 B.n163 163.367
R1149 B.n574 B.n573 163.367
R1150 B.n573 B.n572 163.367
R1151 B.n572 B.n165 163.367
R1152 B.n568 B.n165 163.367
R1153 B.n568 B.n567 163.367
R1154 B.n567 B.n566 163.367
R1155 B.n566 B.n167 163.367
R1156 B.n562 B.n167 163.367
R1157 B.n562 B.n561 163.367
R1158 B.n561 B.n560 163.367
R1159 B.n950 B.n35 163.367
R1160 B.n946 B.n35 163.367
R1161 B.n946 B.n945 163.367
R1162 B.n945 B.n944 163.367
R1163 B.n944 B.n37 163.367
R1164 B.n940 B.n37 163.367
R1165 B.n940 B.n939 163.367
R1166 B.n939 B.n938 163.367
R1167 B.n938 B.n39 163.367
R1168 B.n934 B.n39 163.367
R1169 B.n934 B.n933 163.367
R1170 B.n933 B.n932 163.367
R1171 B.n932 B.n41 163.367
R1172 B.n928 B.n41 163.367
R1173 B.n928 B.n927 163.367
R1174 B.n927 B.n926 163.367
R1175 B.n926 B.n43 163.367
R1176 B.n922 B.n43 163.367
R1177 B.n922 B.n921 163.367
R1178 B.n921 B.n920 163.367
R1179 B.n920 B.n45 163.367
R1180 B.n916 B.n45 163.367
R1181 B.n916 B.n915 163.367
R1182 B.n915 B.n914 163.367
R1183 B.n914 B.n47 163.367
R1184 B.n910 B.n47 163.367
R1185 B.n910 B.n909 163.367
R1186 B.n909 B.n908 163.367
R1187 B.n908 B.n49 163.367
R1188 B.n904 B.n49 163.367
R1189 B.n904 B.n903 163.367
R1190 B.n903 B.n902 163.367
R1191 B.n902 B.n51 163.367
R1192 B.n898 B.n51 163.367
R1193 B.n898 B.n897 163.367
R1194 B.n897 B.n896 163.367
R1195 B.n896 B.n53 163.367
R1196 B.n892 B.n53 163.367
R1197 B.n892 B.n891 163.367
R1198 B.n891 B.n890 163.367
R1199 B.n890 B.n55 163.367
R1200 B.n886 B.n55 163.367
R1201 B.n886 B.n885 163.367
R1202 B.n885 B.n884 163.367
R1203 B.n884 B.n57 163.367
R1204 B.n880 B.n57 163.367
R1205 B.n880 B.n879 163.367
R1206 B.n879 B.n878 163.367
R1207 B.n878 B.n59 163.367
R1208 B.n874 B.n59 163.367
R1209 B.n874 B.n873 163.367
R1210 B.n873 B.n872 163.367
R1211 B.n872 B.n61 163.367
R1212 B.n868 B.n61 163.367
R1213 B.n868 B.n867 163.367
R1214 B.n867 B.n866 163.367
R1215 B.n866 B.n63 163.367
R1216 B.n862 B.n63 163.367
R1217 B.n862 B.n861 163.367
R1218 B.n861 B.n67 163.367
R1219 B.n857 B.n67 163.367
R1220 B.n857 B.n856 163.367
R1221 B.n856 B.n855 163.367
R1222 B.n855 B.n69 163.367
R1223 B.n851 B.n69 163.367
R1224 B.n851 B.n850 163.367
R1225 B.n850 B.n849 163.367
R1226 B.n849 B.n71 163.367
R1227 B.n844 B.n71 163.367
R1228 B.n844 B.n843 163.367
R1229 B.n843 B.n842 163.367
R1230 B.n842 B.n75 163.367
R1231 B.n838 B.n75 163.367
R1232 B.n838 B.n837 163.367
R1233 B.n837 B.n836 163.367
R1234 B.n836 B.n77 163.367
R1235 B.n832 B.n77 163.367
R1236 B.n832 B.n831 163.367
R1237 B.n831 B.n830 163.367
R1238 B.n830 B.n79 163.367
R1239 B.n826 B.n79 163.367
R1240 B.n826 B.n825 163.367
R1241 B.n825 B.n824 163.367
R1242 B.n824 B.n81 163.367
R1243 B.n820 B.n81 163.367
R1244 B.n820 B.n819 163.367
R1245 B.n819 B.n818 163.367
R1246 B.n818 B.n83 163.367
R1247 B.n814 B.n83 163.367
R1248 B.n814 B.n813 163.367
R1249 B.n813 B.n812 163.367
R1250 B.n812 B.n85 163.367
R1251 B.n808 B.n85 163.367
R1252 B.n808 B.n807 163.367
R1253 B.n807 B.n806 163.367
R1254 B.n806 B.n87 163.367
R1255 B.n802 B.n87 163.367
R1256 B.n802 B.n801 163.367
R1257 B.n801 B.n800 163.367
R1258 B.n800 B.n89 163.367
R1259 B.n796 B.n89 163.367
R1260 B.n796 B.n795 163.367
R1261 B.n795 B.n794 163.367
R1262 B.n794 B.n91 163.367
R1263 B.n790 B.n91 163.367
R1264 B.n790 B.n789 163.367
R1265 B.n789 B.n788 163.367
R1266 B.n788 B.n93 163.367
R1267 B.n784 B.n93 163.367
R1268 B.n784 B.n783 163.367
R1269 B.n783 B.n782 163.367
R1270 B.n782 B.n95 163.367
R1271 B.n778 B.n95 163.367
R1272 B.n778 B.n777 163.367
R1273 B.n777 B.n776 163.367
R1274 B.n776 B.n97 163.367
R1275 B.n772 B.n97 163.367
R1276 B.n772 B.n771 163.367
R1277 B.n771 B.n770 163.367
R1278 B.n770 B.n99 163.367
R1279 B.n766 B.n99 163.367
R1280 B.n766 B.n765 163.367
R1281 B.n765 B.n764 163.367
R1282 B.n764 B.n101 163.367
R1283 B.n760 B.n101 163.367
R1284 B.n760 B.n759 163.367
R1285 B.n759 B.n758 163.367
R1286 B.n952 B.n951 163.367
R1287 B.n952 B.n33 163.367
R1288 B.n956 B.n33 163.367
R1289 B.n957 B.n956 163.367
R1290 B.n958 B.n957 163.367
R1291 B.n958 B.n31 163.367
R1292 B.n962 B.n31 163.367
R1293 B.n963 B.n962 163.367
R1294 B.n964 B.n963 163.367
R1295 B.n964 B.n29 163.367
R1296 B.n968 B.n29 163.367
R1297 B.n969 B.n968 163.367
R1298 B.n970 B.n969 163.367
R1299 B.n970 B.n27 163.367
R1300 B.n974 B.n27 163.367
R1301 B.n975 B.n974 163.367
R1302 B.n976 B.n975 163.367
R1303 B.n976 B.n25 163.367
R1304 B.n980 B.n25 163.367
R1305 B.n981 B.n980 163.367
R1306 B.n982 B.n981 163.367
R1307 B.n982 B.n23 163.367
R1308 B.n986 B.n23 163.367
R1309 B.n987 B.n986 163.367
R1310 B.n988 B.n987 163.367
R1311 B.n988 B.n21 163.367
R1312 B.n992 B.n21 163.367
R1313 B.n993 B.n992 163.367
R1314 B.n994 B.n993 163.367
R1315 B.n994 B.n19 163.367
R1316 B.n998 B.n19 163.367
R1317 B.n999 B.n998 163.367
R1318 B.n1000 B.n999 163.367
R1319 B.n1000 B.n17 163.367
R1320 B.n1004 B.n17 163.367
R1321 B.n1005 B.n1004 163.367
R1322 B.n1006 B.n1005 163.367
R1323 B.n1006 B.n15 163.367
R1324 B.n1010 B.n15 163.367
R1325 B.n1011 B.n1010 163.367
R1326 B.n1012 B.n1011 163.367
R1327 B.n1012 B.n13 163.367
R1328 B.n1016 B.n13 163.367
R1329 B.n1017 B.n1016 163.367
R1330 B.n1018 B.n1017 163.367
R1331 B.n1018 B.n11 163.367
R1332 B.n1022 B.n11 163.367
R1333 B.n1023 B.n1022 163.367
R1334 B.n1024 B.n1023 163.367
R1335 B.n1024 B.n9 163.367
R1336 B.n1028 B.n9 163.367
R1337 B.n1029 B.n1028 163.367
R1338 B.n1030 B.n1029 163.367
R1339 B.n1030 B.n7 163.367
R1340 B.n1034 B.n7 163.367
R1341 B.n1035 B.n1034 163.367
R1342 B.n1036 B.n1035 163.367
R1343 B.n1036 B.n5 163.367
R1344 B.n1040 B.n5 163.367
R1345 B.n1041 B.n1040 163.367
R1346 B.n1042 B.n1041 163.367
R1347 B.n1042 B.n3 163.367
R1348 B.n1046 B.n3 163.367
R1349 B.n1047 B.n1046 163.367
R1350 B.n268 B.n2 163.367
R1351 B.n269 B.n268 163.367
R1352 B.n270 B.n269 163.367
R1353 B.n270 B.n265 163.367
R1354 B.n274 B.n265 163.367
R1355 B.n275 B.n274 163.367
R1356 B.n276 B.n275 163.367
R1357 B.n276 B.n263 163.367
R1358 B.n280 B.n263 163.367
R1359 B.n281 B.n280 163.367
R1360 B.n282 B.n281 163.367
R1361 B.n282 B.n261 163.367
R1362 B.n286 B.n261 163.367
R1363 B.n287 B.n286 163.367
R1364 B.n288 B.n287 163.367
R1365 B.n288 B.n259 163.367
R1366 B.n292 B.n259 163.367
R1367 B.n293 B.n292 163.367
R1368 B.n294 B.n293 163.367
R1369 B.n294 B.n257 163.367
R1370 B.n298 B.n257 163.367
R1371 B.n299 B.n298 163.367
R1372 B.n300 B.n299 163.367
R1373 B.n300 B.n255 163.367
R1374 B.n304 B.n255 163.367
R1375 B.n305 B.n304 163.367
R1376 B.n306 B.n305 163.367
R1377 B.n306 B.n253 163.367
R1378 B.n310 B.n253 163.367
R1379 B.n311 B.n310 163.367
R1380 B.n312 B.n311 163.367
R1381 B.n312 B.n251 163.367
R1382 B.n316 B.n251 163.367
R1383 B.n317 B.n316 163.367
R1384 B.n318 B.n317 163.367
R1385 B.n318 B.n249 163.367
R1386 B.n322 B.n249 163.367
R1387 B.n323 B.n322 163.367
R1388 B.n324 B.n323 163.367
R1389 B.n324 B.n247 163.367
R1390 B.n328 B.n247 163.367
R1391 B.n329 B.n328 163.367
R1392 B.n330 B.n329 163.367
R1393 B.n330 B.n245 163.367
R1394 B.n334 B.n245 163.367
R1395 B.n335 B.n334 163.367
R1396 B.n336 B.n335 163.367
R1397 B.n336 B.n243 163.367
R1398 B.n340 B.n243 163.367
R1399 B.n341 B.n340 163.367
R1400 B.n342 B.n341 163.367
R1401 B.n342 B.n241 163.367
R1402 B.n346 B.n241 163.367
R1403 B.n347 B.n346 163.367
R1404 B.n348 B.n347 163.367
R1405 B.n348 B.n239 163.367
R1406 B.n352 B.n239 163.367
R1407 B.n353 B.n352 163.367
R1408 B.n354 B.n353 163.367
R1409 B.n354 B.n237 163.367
R1410 B.n358 B.n237 163.367
R1411 B.n359 B.n358 163.367
R1412 B.n360 B.n359 163.367
R1413 B.n360 B.n235 163.367
R1414 B.n467 B.t8 111.832
R1415 B.n73 B.t1 111.832
R1416 B.n205 B.t5 111.808
R1417 B.n65 B.t10 111.808
R1418 B.n205 B.n204 62.8369
R1419 B.n467 B.n466 62.8369
R1420 B.n73 B.n72 62.8369
R1421 B.n65 B.n64 62.8369
R1422 B.n452 B.n205 59.5399
R1423 B.n468 B.n467 59.5399
R1424 B.n846 B.n73 59.5399
R1425 B.n66 B.n65 59.5399
R1426 B.n949 B.n34 29.8151
R1427 B.n757 B.n756 29.8151
R1428 B.n363 B.n362 29.8151
R1429 B.n559 B.n558 29.8151
R1430 B B.n1049 18.0485
R1431 B.n953 B.n34 10.6151
R1432 B.n954 B.n953 10.6151
R1433 B.n955 B.n954 10.6151
R1434 B.n955 B.n32 10.6151
R1435 B.n959 B.n32 10.6151
R1436 B.n960 B.n959 10.6151
R1437 B.n961 B.n960 10.6151
R1438 B.n961 B.n30 10.6151
R1439 B.n965 B.n30 10.6151
R1440 B.n966 B.n965 10.6151
R1441 B.n967 B.n966 10.6151
R1442 B.n967 B.n28 10.6151
R1443 B.n971 B.n28 10.6151
R1444 B.n972 B.n971 10.6151
R1445 B.n973 B.n972 10.6151
R1446 B.n973 B.n26 10.6151
R1447 B.n977 B.n26 10.6151
R1448 B.n978 B.n977 10.6151
R1449 B.n979 B.n978 10.6151
R1450 B.n979 B.n24 10.6151
R1451 B.n983 B.n24 10.6151
R1452 B.n984 B.n983 10.6151
R1453 B.n985 B.n984 10.6151
R1454 B.n985 B.n22 10.6151
R1455 B.n989 B.n22 10.6151
R1456 B.n990 B.n989 10.6151
R1457 B.n991 B.n990 10.6151
R1458 B.n991 B.n20 10.6151
R1459 B.n995 B.n20 10.6151
R1460 B.n996 B.n995 10.6151
R1461 B.n997 B.n996 10.6151
R1462 B.n997 B.n18 10.6151
R1463 B.n1001 B.n18 10.6151
R1464 B.n1002 B.n1001 10.6151
R1465 B.n1003 B.n1002 10.6151
R1466 B.n1003 B.n16 10.6151
R1467 B.n1007 B.n16 10.6151
R1468 B.n1008 B.n1007 10.6151
R1469 B.n1009 B.n1008 10.6151
R1470 B.n1009 B.n14 10.6151
R1471 B.n1013 B.n14 10.6151
R1472 B.n1014 B.n1013 10.6151
R1473 B.n1015 B.n1014 10.6151
R1474 B.n1015 B.n12 10.6151
R1475 B.n1019 B.n12 10.6151
R1476 B.n1020 B.n1019 10.6151
R1477 B.n1021 B.n1020 10.6151
R1478 B.n1021 B.n10 10.6151
R1479 B.n1025 B.n10 10.6151
R1480 B.n1026 B.n1025 10.6151
R1481 B.n1027 B.n1026 10.6151
R1482 B.n1027 B.n8 10.6151
R1483 B.n1031 B.n8 10.6151
R1484 B.n1032 B.n1031 10.6151
R1485 B.n1033 B.n1032 10.6151
R1486 B.n1033 B.n6 10.6151
R1487 B.n1037 B.n6 10.6151
R1488 B.n1038 B.n1037 10.6151
R1489 B.n1039 B.n1038 10.6151
R1490 B.n1039 B.n4 10.6151
R1491 B.n1043 B.n4 10.6151
R1492 B.n1044 B.n1043 10.6151
R1493 B.n1045 B.n1044 10.6151
R1494 B.n1045 B.n0 10.6151
R1495 B.n949 B.n948 10.6151
R1496 B.n948 B.n947 10.6151
R1497 B.n947 B.n36 10.6151
R1498 B.n943 B.n36 10.6151
R1499 B.n943 B.n942 10.6151
R1500 B.n942 B.n941 10.6151
R1501 B.n941 B.n38 10.6151
R1502 B.n937 B.n38 10.6151
R1503 B.n937 B.n936 10.6151
R1504 B.n936 B.n935 10.6151
R1505 B.n935 B.n40 10.6151
R1506 B.n931 B.n40 10.6151
R1507 B.n931 B.n930 10.6151
R1508 B.n930 B.n929 10.6151
R1509 B.n929 B.n42 10.6151
R1510 B.n925 B.n42 10.6151
R1511 B.n925 B.n924 10.6151
R1512 B.n924 B.n923 10.6151
R1513 B.n923 B.n44 10.6151
R1514 B.n919 B.n44 10.6151
R1515 B.n919 B.n918 10.6151
R1516 B.n918 B.n917 10.6151
R1517 B.n917 B.n46 10.6151
R1518 B.n913 B.n46 10.6151
R1519 B.n913 B.n912 10.6151
R1520 B.n912 B.n911 10.6151
R1521 B.n911 B.n48 10.6151
R1522 B.n907 B.n48 10.6151
R1523 B.n907 B.n906 10.6151
R1524 B.n906 B.n905 10.6151
R1525 B.n905 B.n50 10.6151
R1526 B.n901 B.n50 10.6151
R1527 B.n901 B.n900 10.6151
R1528 B.n900 B.n899 10.6151
R1529 B.n899 B.n52 10.6151
R1530 B.n895 B.n52 10.6151
R1531 B.n895 B.n894 10.6151
R1532 B.n894 B.n893 10.6151
R1533 B.n893 B.n54 10.6151
R1534 B.n889 B.n54 10.6151
R1535 B.n889 B.n888 10.6151
R1536 B.n888 B.n887 10.6151
R1537 B.n887 B.n56 10.6151
R1538 B.n883 B.n56 10.6151
R1539 B.n883 B.n882 10.6151
R1540 B.n882 B.n881 10.6151
R1541 B.n881 B.n58 10.6151
R1542 B.n877 B.n58 10.6151
R1543 B.n877 B.n876 10.6151
R1544 B.n876 B.n875 10.6151
R1545 B.n875 B.n60 10.6151
R1546 B.n871 B.n60 10.6151
R1547 B.n871 B.n870 10.6151
R1548 B.n870 B.n869 10.6151
R1549 B.n869 B.n62 10.6151
R1550 B.n865 B.n62 10.6151
R1551 B.n865 B.n864 10.6151
R1552 B.n864 B.n863 10.6151
R1553 B.n860 B.n859 10.6151
R1554 B.n859 B.n858 10.6151
R1555 B.n858 B.n68 10.6151
R1556 B.n854 B.n68 10.6151
R1557 B.n854 B.n853 10.6151
R1558 B.n853 B.n852 10.6151
R1559 B.n852 B.n70 10.6151
R1560 B.n848 B.n70 10.6151
R1561 B.n848 B.n847 10.6151
R1562 B.n845 B.n74 10.6151
R1563 B.n841 B.n74 10.6151
R1564 B.n841 B.n840 10.6151
R1565 B.n840 B.n839 10.6151
R1566 B.n839 B.n76 10.6151
R1567 B.n835 B.n76 10.6151
R1568 B.n835 B.n834 10.6151
R1569 B.n834 B.n833 10.6151
R1570 B.n833 B.n78 10.6151
R1571 B.n829 B.n78 10.6151
R1572 B.n829 B.n828 10.6151
R1573 B.n828 B.n827 10.6151
R1574 B.n827 B.n80 10.6151
R1575 B.n823 B.n80 10.6151
R1576 B.n823 B.n822 10.6151
R1577 B.n822 B.n821 10.6151
R1578 B.n821 B.n82 10.6151
R1579 B.n817 B.n82 10.6151
R1580 B.n817 B.n816 10.6151
R1581 B.n816 B.n815 10.6151
R1582 B.n815 B.n84 10.6151
R1583 B.n811 B.n84 10.6151
R1584 B.n811 B.n810 10.6151
R1585 B.n810 B.n809 10.6151
R1586 B.n809 B.n86 10.6151
R1587 B.n805 B.n86 10.6151
R1588 B.n805 B.n804 10.6151
R1589 B.n804 B.n803 10.6151
R1590 B.n803 B.n88 10.6151
R1591 B.n799 B.n88 10.6151
R1592 B.n799 B.n798 10.6151
R1593 B.n798 B.n797 10.6151
R1594 B.n797 B.n90 10.6151
R1595 B.n793 B.n90 10.6151
R1596 B.n793 B.n792 10.6151
R1597 B.n792 B.n791 10.6151
R1598 B.n791 B.n92 10.6151
R1599 B.n787 B.n92 10.6151
R1600 B.n787 B.n786 10.6151
R1601 B.n786 B.n785 10.6151
R1602 B.n785 B.n94 10.6151
R1603 B.n781 B.n94 10.6151
R1604 B.n781 B.n780 10.6151
R1605 B.n780 B.n779 10.6151
R1606 B.n779 B.n96 10.6151
R1607 B.n775 B.n96 10.6151
R1608 B.n775 B.n774 10.6151
R1609 B.n774 B.n773 10.6151
R1610 B.n773 B.n98 10.6151
R1611 B.n769 B.n98 10.6151
R1612 B.n769 B.n768 10.6151
R1613 B.n768 B.n767 10.6151
R1614 B.n767 B.n100 10.6151
R1615 B.n763 B.n100 10.6151
R1616 B.n763 B.n762 10.6151
R1617 B.n762 B.n761 10.6151
R1618 B.n761 B.n102 10.6151
R1619 B.n757 B.n102 10.6151
R1620 B.n756 B.n755 10.6151
R1621 B.n755 B.n104 10.6151
R1622 B.n751 B.n104 10.6151
R1623 B.n751 B.n750 10.6151
R1624 B.n750 B.n749 10.6151
R1625 B.n749 B.n106 10.6151
R1626 B.n745 B.n106 10.6151
R1627 B.n745 B.n744 10.6151
R1628 B.n744 B.n743 10.6151
R1629 B.n743 B.n108 10.6151
R1630 B.n739 B.n108 10.6151
R1631 B.n739 B.n738 10.6151
R1632 B.n738 B.n737 10.6151
R1633 B.n737 B.n110 10.6151
R1634 B.n733 B.n110 10.6151
R1635 B.n733 B.n732 10.6151
R1636 B.n732 B.n731 10.6151
R1637 B.n731 B.n112 10.6151
R1638 B.n727 B.n112 10.6151
R1639 B.n727 B.n726 10.6151
R1640 B.n726 B.n725 10.6151
R1641 B.n725 B.n114 10.6151
R1642 B.n721 B.n114 10.6151
R1643 B.n721 B.n720 10.6151
R1644 B.n720 B.n719 10.6151
R1645 B.n719 B.n116 10.6151
R1646 B.n715 B.n116 10.6151
R1647 B.n715 B.n714 10.6151
R1648 B.n714 B.n713 10.6151
R1649 B.n713 B.n118 10.6151
R1650 B.n709 B.n118 10.6151
R1651 B.n709 B.n708 10.6151
R1652 B.n708 B.n707 10.6151
R1653 B.n707 B.n120 10.6151
R1654 B.n703 B.n120 10.6151
R1655 B.n703 B.n702 10.6151
R1656 B.n702 B.n701 10.6151
R1657 B.n701 B.n122 10.6151
R1658 B.n697 B.n122 10.6151
R1659 B.n697 B.n696 10.6151
R1660 B.n696 B.n695 10.6151
R1661 B.n695 B.n124 10.6151
R1662 B.n691 B.n124 10.6151
R1663 B.n691 B.n690 10.6151
R1664 B.n690 B.n689 10.6151
R1665 B.n689 B.n126 10.6151
R1666 B.n685 B.n126 10.6151
R1667 B.n685 B.n684 10.6151
R1668 B.n684 B.n683 10.6151
R1669 B.n683 B.n128 10.6151
R1670 B.n679 B.n128 10.6151
R1671 B.n679 B.n678 10.6151
R1672 B.n678 B.n677 10.6151
R1673 B.n677 B.n130 10.6151
R1674 B.n673 B.n130 10.6151
R1675 B.n673 B.n672 10.6151
R1676 B.n672 B.n671 10.6151
R1677 B.n671 B.n132 10.6151
R1678 B.n667 B.n132 10.6151
R1679 B.n667 B.n666 10.6151
R1680 B.n666 B.n665 10.6151
R1681 B.n665 B.n134 10.6151
R1682 B.n661 B.n134 10.6151
R1683 B.n661 B.n660 10.6151
R1684 B.n660 B.n659 10.6151
R1685 B.n659 B.n136 10.6151
R1686 B.n655 B.n136 10.6151
R1687 B.n655 B.n654 10.6151
R1688 B.n654 B.n653 10.6151
R1689 B.n653 B.n138 10.6151
R1690 B.n649 B.n138 10.6151
R1691 B.n649 B.n648 10.6151
R1692 B.n648 B.n647 10.6151
R1693 B.n647 B.n140 10.6151
R1694 B.n643 B.n140 10.6151
R1695 B.n643 B.n642 10.6151
R1696 B.n642 B.n641 10.6151
R1697 B.n641 B.n142 10.6151
R1698 B.n637 B.n142 10.6151
R1699 B.n637 B.n636 10.6151
R1700 B.n636 B.n635 10.6151
R1701 B.n635 B.n144 10.6151
R1702 B.n631 B.n144 10.6151
R1703 B.n631 B.n630 10.6151
R1704 B.n630 B.n629 10.6151
R1705 B.n629 B.n146 10.6151
R1706 B.n625 B.n146 10.6151
R1707 B.n625 B.n624 10.6151
R1708 B.n624 B.n623 10.6151
R1709 B.n623 B.n148 10.6151
R1710 B.n619 B.n148 10.6151
R1711 B.n619 B.n618 10.6151
R1712 B.n618 B.n617 10.6151
R1713 B.n617 B.n150 10.6151
R1714 B.n613 B.n150 10.6151
R1715 B.n613 B.n612 10.6151
R1716 B.n612 B.n611 10.6151
R1717 B.n611 B.n152 10.6151
R1718 B.n607 B.n152 10.6151
R1719 B.n607 B.n606 10.6151
R1720 B.n606 B.n605 10.6151
R1721 B.n605 B.n154 10.6151
R1722 B.n601 B.n154 10.6151
R1723 B.n601 B.n600 10.6151
R1724 B.n600 B.n599 10.6151
R1725 B.n599 B.n156 10.6151
R1726 B.n595 B.n156 10.6151
R1727 B.n595 B.n594 10.6151
R1728 B.n594 B.n593 10.6151
R1729 B.n593 B.n158 10.6151
R1730 B.n589 B.n158 10.6151
R1731 B.n589 B.n588 10.6151
R1732 B.n588 B.n587 10.6151
R1733 B.n587 B.n160 10.6151
R1734 B.n583 B.n160 10.6151
R1735 B.n583 B.n582 10.6151
R1736 B.n582 B.n581 10.6151
R1737 B.n581 B.n162 10.6151
R1738 B.n577 B.n162 10.6151
R1739 B.n577 B.n576 10.6151
R1740 B.n576 B.n575 10.6151
R1741 B.n575 B.n164 10.6151
R1742 B.n571 B.n164 10.6151
R1743 B.n571 B.n570 10.6151
R1744 B.n570 B.n569 10.6151
R1745 B.n569 B.n166 10.6151
R1746 B.n565 B.n166 10.6151
R1747 B.n565 B.n564 10.6151
R1748 B.n564 B.n563 10.6151
R1749 B.n563 B.n168 10.6151
R1750 B.n559 B.n168 10.6151
R1751 B.n267 B.n1 10.6151
R1752 B.n267 B.n266 10.6151
R1753 B.n271 B.n266 10.6151
R1754 B.n272 B.n271 10.6151
R1755 B.n273 B.n272 10.6151
R1756 B.n273 B.n264 10.6151
R1757 B.n277 B.n264 10.6151
R1758 B.n278 B.n277 10.6151
R1759 B.n279 B.n278 10.6151
R1760 B.n279 B.n262 10.6151
R1761 B.n283 B.n262 10.6151
R1762 B.n284 B.n283 10.6151
R1763 B.n285 B.n284 10.6151
R1764 B.n285 B.n260 10.6151
R1765 B.n289 B.n260 10.6151
R1766 B.n290 B.n289 10.6151
R1767 B.n291 B.n290 10.6151
R1768 B.n291 B.n258 10.6151
R1769 B.n295 B.n258 10.6151
R1770 B.n296 B.n295 10.6151
R1771 B.n297 B.n296 10.6151
R1772 B.n297 B.n256 10.6151
R1773 B.n301 B.n256 10.6151
R1774 B.n302 B.n301 10.6151
R1775 B.n303 B.n302 10.6151
R1776 B.n303 B.n254 10.6151
R1777 B.n307 B.n254 10.6151
R1778 B.n308 B.n307 10.6151
R1779 B.n309 B.n308 10.6151
R1780 B.n309 B.n252 10.6151
R1781 B.n313 B.n252 10.6151
R1782 B.n314 B.n313 10.6151
R1783 B.n315 B.n314 10.6151
R1784 B.n315 B.n250 10.6151
R1785 B.n319 B.n250 10.6151
R1786 B.n320 B.n319 10.6151
R1787 B.n321 B.n320 10.6151
R1788 B.n321 B.n248 10.6151
R1789 B.n325 B.n248 10.6151
R1790 B.n326 B.n325 10.6151
R1791 B.n327 B.n326 10.6151
R1792 B.n327 B.n246 10.6151
R1793 B.n331 B.n246 10.6151
R1794 B.n332 B.n331 10.6151
R1795 B.n333 B.n332 10.6151
R1796 B.n333 B.n244 10.6151
R1797 B.n337 B.n244 10.6151
R1798 B.n338 B.n337 10.6151
R1799 B.n339 B.n338 10.6151
R1800 B.n339 B.n242 10.6151
R1801 B.n343 B.n242 10.6151
R1802 B.n344 B.n343 10.6151
R1803 B.n345 B.n344 10.6151
R1804 B.n345 B.n240 10.6151
R1805 B.n349 B.n240 10.6151
R1806 B.n350 B.n349 10.6151
R1807 B.n351 B.n350 10.6151
R1808 B.n351 B.n238 10.6151
R1809 B.n355 B.n238 10.6151
R1810 B.n356 B.n355 10.6151
R1811 B.n357 B.n356 10.6151
R1812 B.n357 B.n236 10.6151
R1813 B.n361 B.n236 10.6151
R1814 B.n362 B.n361 10.6151
R1815 B.n363 B.n234 10.6151
R1816 B.n367 B.n234 10.6151
R1817 B.n368 B.n367 10.6151
R1818 B.n369 B.n368 10.6151
R1819 B.n369 B.n232 10.6151
R1820 B.n373 B.n232 10.6151
R1821 B.n374 B.n373 10.6151
R1822 B.n375 B.n374 10.6151
R1823 B.n375 B.n230 10.6151
R1824 B.n379 B.n230 10.6151
R1825 B.n380 B.n379 10.6151
R1826 B.n381 B.n380 10.6151
R1827 B.n381 B.n228 10.6151
R1828 B.n385 B.n228 10.6151
R1829 B.n386 B.n385 10.6151
R1830 B.n387 B.n386 10.6151
R1831 B.n387 B.n226 10.6151
R1832 B.n391 B.n226 10.6151
R1833 B.n392 B.n391 10.6151
R1834 B.n393 B.n392 10.6151
R1835 B.n393 B.n224 10.6151
R1836 B.n397 B.n224 10.6151
R1837 B.n398 B.n397 10.6151
R1838 B.n399 B.n398 10.6151
R1839 B.n399 B.n222 10.6151
R1840 B.n403 B.n222 10.6151
R1841 B.n404 B.n403 10.6151
R1842 B.n405 B.n404 10.6151
R1843 B.n405 B.n220 10.6151
R1844 B.n409 B.n220 10.6151
R1845 B.n410 B.n409 10.6151
R1846 B.n411 B.n410 10.6151
R1847 B.n411 B.n218 10.6151
R1848 B.n415 B.n218 10.6151
R1849 B.n416 B.n415 10.6151
R1850 B.n417 B.n416 10.6151
R1851 B.n417 B.n216 10.6151
R1852 B.n421 B.n216 10.6151
R1853 B.n422 B.n421 10.6151
R1854 B.n423 B.n422 10.6151
R1855 B.n423 B.n214 10.6151
R1856 B.n427 B.n214 10.6151
R1857 B.n428 B.n427 10.6151
R1858 B.n429 B.n428 10.6151
R1859 B.n429 B.n212 10.6151
R1860 B.n433 B.n212 10.6151
R1861 B.n434 B.n433 10.6151
R1862 B.n435 B.n434 10.6151
R1863 B.n435 B.n210 10.6151
R1864 B.n439 B.n210 10.6151
R1865 B.n440 B.n439 10.6151
R1866 B.n441 B.n440 10.6151
R1867 B.n441 B.n208 10.6151
R1868 B.n445 B.n208 10.6151
R1869 B.n446 B.n445 10.6151
R1870 B.n447 B.n446 10.6151
R1871 B.n447 B.n206 10.6151
R1872 B.n451 B.n206 10.6151
R1873 B.n454 B.n453 10.6151
R1874 B.n454 B.n202 10.6151
R1875 B.n458 B.n202 10.6151
R1876 B.n459 B.n458 10.6151
R1877 B.n460 B.n459 10.6151
R1878 B.n460 B.n200 10.6151
R1879 B.n464 B.n200 10.6151
R1880 B.n465 B.n464 10.6151
R1881 B.n469 B.n465 10.6151
R1882 B.n473 B.n198 10.6151
R1883 B.n474 B.n473 10.6151
R1884 B.n475 B.n474 10.6151
R1885 B.n475 B.n196 10.6151
R1886 B.n479 B.n196 10.6151
R1887 B.n480 B.n479 10.6151
R1888 B.n481 B.n480 10.6151
R1889 B.n481 B.n194 10.6151
R1890 B.n485 B.n194 10.6151
R1891 B.n486 B.n485 10.6151
R1892 B.n487 B.n486 10.6151
R1893 B.n487 B.n192 10.6151
R1894 B.n491 B.n192 10.6151
R1895 B.n492 B.n491 10.6151
R1896 B.n493 B.n492 10.6151
R1897 B.n493 B.n190 10.6151
R1898 B.n497 B.n190 10.6151
R1899 B.n498 B.n497 10.6151
R1900 B.n499 B.n498 10.6151
R1901 B.n499 B.n188 10.6151
R1902 B.n503 B.n188 10.6151
R1903 B.n504 B.n503 10.6151
R1904 B.n505 B.n504 10.6151
R1905 B.n505 B.n186 10.6151
R1906 B.n509 B.n186 10.6151
R1907 B.n510 B.n509 10.6151
R1908 B.n511 B.n510 10.6151
R1909 B.n511 B.n184 10.6151
R1910 B.n515 B.n184 10.6151
R1911 B.n516 B.n515 10.6151
R1912 B.n517 B.n516 10.6151
R1913 B.n517 B.n182 10.6151
R1914 B.n521 B.n182 10.6151
R1915 B.n522 B.n521 10.6151
R1916 B.n523 B.n522 10.6151
R1917 B.n523 B.n180 10.6151
R1918 B.n527 B.n180 10.6151
R1919 B.n528 B.n527 10.6151
R1920 B.n529 B.n528 10.6151
R1921 B.n529 B.n178 10.6151
R1922 B.n533 B.n178 10.6151
R1923 B.n534 B.n533 10.6151
R1924 B.n535 B.n534 10.6151
R1925 B.n535 B.n176 10.6151
R1926 B.n539 B.n176 10.6151
R1927 B.n540 B.n539 10.6151
R1928 B.n541 B.n540 10.6151
R1929 B.n541 B.n174 10.6151
R1930 B.n545 B.n174 10.6151
R1931 B.n546 B.n545 10.6151
R1932 B.n547 B.n546 10.6151
R1933 B.n547 B.n172 10.6151
R1934 B.n551 B.n172 10.6151
R1935 B.n552 B.n551 10.6151
R1936 B.n553 B.n552 10.6151
R1937 B.n553 B.n170 10.6151
R1938 B.n557 B.n170 10.6151
R1939 B.n558 B.n557 10.6151
R1940 B.n863 B.n66 9.36635
R1941 B.n846 B.n845 9.36635
R1942 B.n452 B.n451 9.36635
R1943 B.n468 B.n198 9.36635
R1944 B.n1049 B.n0 8.11757
R1945 B.n1049 B.n1 8.11757
R1946 B.n860 B.n66 1.24928
R1947 B.n847 B.n846 1.24928
R1948 B.n453 B.n452 1.24928
R1949 B.n469 B.n468 1.24928
C0 w_n4858_n4562# VN 10.597401f
C1 w_n4858_n4562# VDD1 3.31957f
C2 B VN 1.43228f
C3 B VDD1 3.07664f
C4 VTAIL VN 16.567099f
C5 VDD1 VTAIL 13.092401f
C6 VP VN 9.96237f
C7 VDD1 VP 16.5241f
C8 VDD2 VN 16.0594f
C9 VDD1 VDD2 2.37705f
C10 w_n4858_n4562# B 12.7421f
C11 w_n4858_n4562# VTAIL 4.07836f
C12 B VTAIL 5.22064f
C13 w_n4858_n4562# VP 11.230901f
C14 B VP 2.49916f
C15 VP VTAIL 16.5814f
C16 w_n4858_n4562# VDD2 3.47923f
C17 B VDD2 3.20663f
C18 VDD2 VTAIL 13.144501f
C19 VP VDD2 0.623584f
C20 VDD1 VN 0.154092f
C21 VDD2 VSUBS 2.40334f
C22 VDD1 VSUBS 2.243401f
C23 VTAIL VSUBS 1.589632f
C24 VN VSUBS 8.42284f
C25 VP VSUBS 4.862926f
C26 B VSUBS 6.255851f
C27 w_n4858_n4562# VSUBS 0.271018p
C28 B.n0 VSUBS 0.007014f
C29 B.n1 VSUBS 0.007014f
C30 B.n2 VSUBS 0.010374f
C31 B.n3 VSUBS 0.007949f
C32 B.n4 VSUBS 0.007949f
C33 B.n5 VSUBS 0.007949f
C34 B.n6 VSUBS 0.007949f
C35 B.n7 VSUBS 0.007949f
C36 B.n8 VSUBS 0.007949f
C37 B.n9 VSUBS 0.007949f
C38 B.n10 VSUBS 0.007949f
C39 B.n11 VSUBS 0.007949f
C40 B.n12 VSUBS 0.007949f
C41 B.n13 VSUBS 0.007949f
C42 B.n14 VSUBS 0.007949f
C43 B.n15 VSUBS 0.007949f
C44 B.n16 VSUBS 0.007949f
C45 B.n17 VSUBS 0.007949f
C46 B.n18 VSUBS 0.007949f
C47 B.n19 VSUBS 0.007949f
C48 B.n20 VSUBS 0.007949f
C49 B.n21 VSUBS 0.007949f
C50 B.n22 VSUBS 0.007949f
C51 B.n23 VSUBS 0.007949f
C52 B.n24 VSUBS 0.007949f
C53 B.n25 VSUBS 0.007949f
C54 B.n26 VSUBS 0.007949f
C55 B.n27 VSUBS 0.007949f
C56 B.n28 VSUBS 0.007949f
C57 B.n29 VSUBS 0.007949f
C58 B.n30 VSUBS 0.007949f
C59 B.n31 VSUBS 0.007949f
C60 B.n32 VSUBS 0.007949f
C61 B.n33 VSUBS 0.007949f
C62 B.n34 VSUBS 0.017197f
C63 B.n35 VSUBS 0.007949f
C64 B.n36 VSUBS 0.007949f
C65 B.n37 VSUBS 0.007949f
C66 B.n38 VSUBS 0.007949f
C67 B.n39 VSUBS 0.007949f
C68 B.n40 VSUBS 0.007949f
C69 B.n41 VSUBS 0.007949f
C70 B.n42 VSUBS 0.007949f
C71 B.n43 VSUBS 0.007949f
C72 B.n44 VSUBS 0.007949f
C73 B.n45 VSUBS 0.007949f
C74 B.n46 VSUBS 0.007949f
C75 B.n47 VSUBS 0.007949f
C76 B.n48 VSUBS 0.007949f
C77 B.n49 VSUBS 0.007949f
C78 B.n50 VSUBS 0.007949f
C79 B.n51 VSUBS 0.007949f
C80 B.n52 VSUBS 0.007949f
C81 B.n53 VSUBS 0.007949f
C82 B.n54 VSUBS 0.007949f
C83 B.n55 VSUBS 0.007949f
C84 B.n56 VSUBS 0.007949f
C85 B.n57 VSUBS 0.007949f
C86 B.n58 VSUBS 0.007949f
C87 B.n59 VSUBS 0.007949f
C88 B.n60 VSUBS 0.007949f
C89 B.n61 VSUBS 0.007949f
C90 B.n62 VSUBS 0.007949f
C91 B.n63 VSUBS 0.007949f
C92 B.t10 VSUBS 0.688886f
C93 B.t11 VSUBS 0.714787f
C94 B.t9 VSUBS 2.65641f
C95 B.n64 VSUBS 0.408404f
C96 B.n65 VSUBS 0.083326f
C97 B.n66 VSUBS 0.018418f
C98 B.n67 VSUBS 0.007949f
C99 B.n68 VSUBS 0.007949f
C100 B.n69 VSUBS 0.007949f
C101 B.n70 VSUBS 0.007949f
C102 B.n71 VSUBS 0.007949f
C103 B.t1 VSUBS 0.688862f
C104 B.t2 VSUBS 0.714768f
C105 B.t0 VSUBS 2.65641f
C106 B.n72 VSUBS 0.408423f
C107 B.n73 VSUBS 0.08335f
C108 B.n74 VSUBS 0.007949f
C109 B.n75 VSUBS 0.007949f
C110 B.n76 VSUBS 0.007949f
C111 B.n77 VSUBS 0.007949f
C112 B.n78 VSUBS 0.007949f
C113 B.n79 VSUBS 0.007949f
C114 B.n80 VSUBS 0.007949f
C115 B.n81 VSUBS 0.007949f
C116 B.n82 VSUBS 0.007949f
C117 B.n83 VSUBS 0.007949f
C118 B.n84 VSUBS 0.007949f
C119 B.n85 VSUBS 0.007949f
C120 B.n86 VSUBS 0.007949f
C121 B.n87 VSUBS 0.007949f
C122 B.n88 VSUBS 0.007949f
C123 B.n89 VSUBS 0.007949f
C124 B.n90 VSUBS 0.007949f
C125 B.n91 VSUBS 0.007949f
C126 B.n92 VSUBS 0.007949f
C127 B.n93 VSUBS 0.007949f
C128 B.n94 VSUBS 0.007949f
C129 B.n95 VSUBS 0.007949f
C130 B.n96 VSUBS 0.007949f
C131 B.n97 VSUBS 0.007949f
C132 B.n98 VSUBS 0.007949f
C133 B.n99 VSUBS 0.007949f
C134 B.n100 VSUBS 0.007949f
C135 B.n101 VSUBS 0.007949f
C136 B.n102 VSUBS 0.007949f
C137 B.n103 VSUBS 0.017197f
C138 B.n104 VSUBS 0.007949f
C139 B.n105 VSUBS 0.007949f
C140 B.n106 VSUBS 0.007949f
C141 B.n107 VSUBS 0.007949f
C142 B.n108 VSUBS 0.007949f
C143 B.n109 VSUBS 0.007949f
C144 B.n110 VSUBS 0.007949f
C145 B.n111 VSUBS 0.007949f
C146 B.n112 VSUBS 0.007949f
C147 B.n113 VSUBS 0.007949f
C148 B.n114 VSUBS 0.007949f
C149 B.n115 VSUBS 0.007949f
C150 B.n116 VSUBS 0.007949f
C151 B.n117 VSUBS 0.007949f
C152 B.n118 VSUBS 0.007949f
C153 B.n119 VSUBS 0.007949f
C154 B.n120 VSUBS 0.007949f
C155 B.n121 VSUBS 0.007949f
C156 B.n122 VSUBS 0.007949f
C157 B.n123 VSUBS 0.007949f
C158 B.n124 VSUBS 0.007949f
C159 B.n125 VSUBS 0.007949f
C160 B.n126 VSUBS 0.007949f
C161 B.n127 VSUBS 0.007949f
C162 B.n128 VSUBS 0.007949f
C163 B.n129 VSUBS 0.007949f
C164 B.n130 VSUBS 0.007949f
C165 B.n131 VSUBS 0.007949f
C166 B.n132 VSUBS 0.007949f
C167 B.n133 VSUBS 0.007949f
C168 B.n134 VSUBS 0.007949f
C169 B.n135 VSUBS 0.007949f
C170 B.n136 VSUBS 0.007949f
C171 B.n137 VSUBS 0.007949f
C172 B.n138 VSUBS 0.007949f
C173 B.n139 VSUBS 0.007949f
C174 B.n140 VSUBS 0.007949f
C175 B.n141 VSUBS 0.007949f
C176 B.n142 VSUBS 0.007949f
C177 B.n143 VSUBS 0.007949f
C178 B.n144 VSUBS 0.007949f
C179 B.n145 VSUBS 0.007949f
C180 B.n146 VSUBS 0.007949f
C181 B.n147 VSUBS 0.007949f
C182 B.n148 VSUBS 0.007949f
C183 B.n149 VSUBS 0.007949f
C184 B.n150 VSUBS 0.007949f
C185 B.n151 VSUBS 0.007949f
C186 B.n152 VSUBS 0.007949f
C187 B.n153 VSUBS 0.007949f
C188 B.n154 VSUBS 0.007949f
C189 B.n155 VSUBS 0.007949f
C190 B.n156 VSUBS 0.007949f
C191 B.n157 VSUBS 0.007949f
C192 B.n158 VSUBS 0.007949f
C193 B.n159 VSUBS 0.007949f
C194 B.n160 VSUBS 0.007949f
C195 B.n161 VSUBS 0.007949f
C196 B.n162 VSUBS 0.007949f
C197 B.n163 VSUBS 0.007949f
C198 B.n164 VSUBS 0.007949f
C199 B.n165 VSUBS 0.007949f
C200 B.n166 VSUBS 0.007949f
C201 B.n167 VSUBS 0.007949f
C202 B.n168 VSUBS 0.007949f
C203 B.n169 VSUBS 0.017874f
C204 B.n170 VSUBS 0.007949f
C205 B.n171 VSUBS 0.007949f
C206 B.n172 VSUBS 0.007949f
C207 B.n173 VSUBS 0.007949f
C208 B.n174 VSUBS 0.007949f
C209 B.n175 VSUBS 0.007949f
C210 B.n176 VSUBS 0.007949f
C211 B.n177 VSUBS 0.007949f
C212 B.n178 VSUBS 0.007949f
C213 B.n179 VSUBS 0.007949f
C214 B.n180 VSUBS 0.007949f
C215 B.n181 VSUBS 0.007949f
C216 B.n182 VSUBS 0.007949f
C217 B.n183 VSUBS 0.007949f
C218 B.n184 VSUBS 0.007949f
C219 B.n185 VSUBS 0.007949f
C220 B.n186 VSUBS 0.007949f
C221 B.n187 VSUBS 0.007949f
C222 B.n188 VSUBS 0.007949f
C223 B.n189 VSUBS 0.007949f
C224 B.n190 VSUBS 0.007949f
C225 B.n191 VSUBS 0.007949f
C226 B.n192 VSUBS 0.007949f
C227 B.n193 VSUBS 0.007949f
C228 B.n194 VSUBS 0.007949f
C229 B.n195 VSUBS 0.007949f
C230 B.n196 VSUBS 0.007949f
C231 B.n197 VSUBS 0.007949f
C232 B.n198 VSUBS 0.007482f
C233 B.n199 VSUBS 0.007949f
C234 B.n200 VSUBS 0.007949f
C235 B.n201 VSUBS 0.007949f
C236 B.n202 VSUBS 0.007949f
C237 B.n203 VSUBS 0.007949f
C238 B.t5 VSUBS 0.688886f
C239 B.t4 VSUBS 0.714787f
C240 B.t3 VSUBS 2.65641f
C241 B.n204 VSUBS 0.408404f
C242 B.n205 VSUBS 0.083326f
C243 B.n206 VSUBS 0.007949f
C244 B.n207 VSUBS 0.007949f
C245 B.n208 VSUBS 0.007949f
C246 B.n209 VSUBS 0.007949f
C247 B.n210 VSUBS 0.007949f
C248 B.n211 VSUBS 0.007949f
C249 B.n212 VSUBS 0.007949f
C250 B.n213 VSUBS 0.007949f
C251 B.n214 VSUBS 0.007949f
C252 B.n215 VSUBS 0.007949f
C253 B.n216 VSUBS 0.007949f
C254 B.n217 VSUBS 0.007949f
C255 B.n218 VSUBS 0.007949f
C256 B.n219 VSUBS 0.007949f
C257 B.n220 VSUBS 0.007949f
C258 B.n221 VSUBS 0.007949f
C259 B.n222 VSUBS 0.007949f
C260 B.n223 VSUBS 0.007949f
C261 B.n224 VSUBS 0.007949f
C262 B.n225 VSUBS 0.007949f
C263 B.n226 VSUBS 0.007949f
C264 B.n227 VSUBS 0.007949f
C265 B.n228 VSUBS 0.007949f
C266 B.n229 VSUBS 0.007949f
C267 B.n230 VSUBS 0.007949f
C268 B.n231 VSUBS 0.007949f
C269 B.n232 VSUBS 0.007949f
C270 B.n233 VSUBS 0.007949f
C271 B.n234 VSUBS 0.007949f
C272 B.n235 VSUBS 0.017197f
C273 B.n236 VSUBS 0.007949f
C274 B.n237 VSUBS 0.007949f
C275 B.n238 VSUBS 0.007949f
C276 B.n239 VSUBS 0.007949f
C277 B.n240 VSUBS 0.007949f
C278 B.n241 VSUBS 0.007949f
C279 B.n242 VSUBS 0.007949f
C280 B.n243 VSUBS 0.007949f
C281 B.n244 VSUBS 0.007949f
C282 B.n245 VSUBS 0.007949f
C283 B.n246 VSUBS 0.007949f
C284 B.n247 VSUBS 0.007949f
C285 B.n248 VSUBS 0.007949f
C286 B.n249 VSUBS 0.007949f
C287 B.n250 VSUBS 0.007949f
C288 B.n251 VSUBS 0.007949f
C289 B.n252 VSUBS 0.007949f
C290 B.n253 VSUBS 0.007949f
C291 B.n254 VSUBS 0.007949f
C292 B.n255 VSUBS 0.007949f
C293 B.n256 VSUBS 0.007949f
C294 B.n257 VSUBS 0.007949f
C295 B.n258 VSUBS 0.007949f
C296 B.n259 VSUBS 0.007949f
C297 B.n260 VSUBS 0.007949f
C298 B.n261 VSUBS 0.007949f
C299 B.n262 VSUBS 0.007949f
C300 B.n263 VSUBS 0.007949f
C301 B.n264 VSUBS 0.007949f
C302 B.n265 VSUBS 0.007949f
C303 B.n266 VSUBS 0.007949f
C304 B.n267 VSUBS 0.007949f
C305 B.n268 VSUBS 0.007949f
C306 B.n269 VSUBS 0.007949f
C307 B.n270 VSUBS 0.007949f
C308 B.n271 VSUBS 0.007949f
C309 B.n272 VSUBS 0.007949f
C310 B.n273 VSUBS 0.007949f
C311 B.n274 VSUBS 0.007949f
C312 B.n275 VSUBS 0.007949f
C313 B.n276 VSUBS 0.007949f
C314 B.n277 VSUBS 0.007949f
C315 B.n278 VSUBS 0.007949f
C316 B.n279 VSUBS 0.007949f
C317 B.n280 VSUBS 0.007949f
C318 B.n281 VSUBS 0.007949f
C319 B.n282 VSUBS 0.007949f
C320 B.n283 VSUBS 0.007949f
C321 B.n284 VSUBS 0.007949f
C322 B.n285 VSUBS 0.007949f
C323 B.n286 VSUBS 0.007949f
C324 B.n287 VSUBS 0.007949f
C325 B.n288 VSUBS 0.007949f
C326 B.n289 VSUBS 0.007949f
C327 B.n290 VSUBS 0.007949f
C328 B.n291 VSUBS 0.007949f
C329 B.n292 VSUBS 0.007949f
C330 B.n293 VSUBS 0.007949f
C331 B.n294 VSUBS 0.007949f
C332 B.n295 VSUBS 0.007949f
C333 B.n296 VSUBS 0.007949f
C334 B.n297 VSUBS 0.007949f
C335 B.n298 VSUBS 0.007949f
C336 B.n299 VSUBS 0.007949f
C337 B.n300 VSUBS 0.007949f
C338 B.n301 VSUBS 0.007949f
C339 B.n302 VSUBS 0.007949f
C340 B.n303 VSUBS 0.007949f
C341 B.n304 VSUBS 0.007949f
C342 B.n305 VSUBS 0.007949f
C343 B.n306 VSUBS 0.007949f
C344 B.n307 VSUBS 0.007949f
C345 B.n308 VSUBS 0.007949f
C346 B.n309 VSUBS 0.007949f
C347 B.n310 VSUBS 0.007949f
C348 B.n311 VSUBS 0.007949f
C349 B.n312 VSUBS 0.007949f
C350 B.n313 VSUBS 0.007949f
C351 B.n314 VSUBS 0.007949f
C352 B.n315 VSUBS 0.007949f
C353 B.n316 VSUBS 0.007949f
C354 B.n317 VSUBS 0.007949f
C355 B.n318 VSUBS 0.007949f
C356 B.n319 VSUBS 0.007949f
C357 B.n320 VSUBS 0.007949f
C358 B.n321 VSUBS 0.007949f
C359 B.n322 VSUBS 0.007949f
C360 B.n323 VSUBS 0.007949f
C361 B.n324 VSUBS 0.007949f
C362 B.n325 VSUBS 0.007949f
C363 B.n326 VSUBS 0.007949f
C364 B.n327 VSUBS 0.007949f
C365 B.n328 VSUBS 0.007949f
C366 B.n329 VSUBS 0.007949f
C367 B.n330 VSUBS 0.007949f
C368 B.n331 VSUBS 0.007949f
C369 B.n332 VSUBS 0.007949f
C370 B.n333 VSUBS 0.007949f
C371 B.n334 VSUBS 0.007949f
C372 B.n335 VSUBS 0.007949f
C373 B.n336 VSUBS 0.007949f
C374 B.n337 VSUBS 0.007949f
C375 B.n338 VSUBS 0.007949f
C376 B.n339 VSUBS 0.007949f
C377 B.n340 VSUBS 0.007949f
C378 B.n341 VSUBS 0.007949f
C379 B.n342 VSUBS 0.007949f
C380 B.n343 VSUBS 0.007949f
C381 B.n344 VSUBS 0.007949f
C382 B.n345 VSUBS 0.007949f
C383 B.n346 VSUBS 0.007949f
C384 B.n347 VSUBS 0.007949f
C385 B.n348 VSUBS 0.007949f
C386 B.n349 VSUBS 0.007949f
C387 B.n350 VSUBS 0.007949f
C388 B.n351 VSUBS 0.007949f
C389 B.n352 VSUBS 0.007949f
C390 B.n353 VSUBS 0.007949f
C391 B.n354 VSUBS 0.007949f
C392 B.n355 VSUBS 0.007949f
C393 B.n356 VSUBS 0.007949f
C394 B.n357 VSUBS 0.007949f
C395 B.n358 VSUBS 0.007949f
C396 B.n359 VSUBS 0.007949f
C397 B.n360 VSUBS 0.007949f
C398 B.n361 VSUBS 0.007949f
C399 B.n362 VSUBS 0.017197f
C400 B.n363 VSUBS 0.017874f
C401 B.n364 VSUBS 0.017874f
C402 B.n365 VSUBS 0.007949f
C403 B.n366 VSUBS 0.007949f
C404 B.n367 VSUBS 0.007949f
C405 B.n368 VSUBS 0.007949f
C406 B.n369 VSUBS 0.007949f
C407 B.n370 VSUBS 0.007949f
C408 B.n371 VSUBS 0.007949f
C409 B.n372 VSUBS 0.007949f
C410 B.n373 VSUBS 0.007949f
C411 B.n374 VSUBS 0.007949f
C412 B.n375 VSUBS 0.007949f
C413 B.n376 VSUBS 0.007949f
C414 B.n377 VSUBS 0.007949f
C415 B.n378 VSUBS 0.007949f
C416 B.n379 VSUBS 0.007949f
C417 B.n380 VSUBS 0.007949f
C418 B.n381 VSUBS 0.007949f
C419 B.n382 VSUBS 0.007949f
C420 B.n383 VSUBS 0.007949f
C421 B.n384 VSUBS 0.007949f
C422 B.n385 VSUBS 0.007949f
C423 B.n386 VSUBS 0.007949f
C424 B.n387 VSUBS 0.007949f
C425 B.n388 VSUBS 0.007949f
C426 B.n389 VSUBS 0.007949f
C427 B.n390 VSUBS 0.007949f
C428 B.n391 VSUBS 0.007949f
C429 B.n392 VSUBS 0.007949f
C430 B.n393 VSUBS 0.007949f
C431 B.n394 VSUBS 0.007949f
C432 B.n395 VSUBS 0.007949f
C433 B.n396 VSUBS 0.007949f
C434 B.n397 VSUBS 0.007949f
C435 B.n398 VSUBS 0.007949f
C436 B.n399 VSUBS 0.007949f
C437 B.n400 VSUBS 0.007949f
C438 B.n401 VSUBS 0.007949f
C439 B.n402 VSUBS 0.007949f
C440 B.n403 VSUBS 0.007949f
C441 B.n404 VSUBS 0.007949f
C442 B.n405 VSUBS 0.007949f
C443 B.n406 VSUBS 0.007949f
C444 B.n407 VSUBS 0.007949f
C445 B.n408 VSUBS 0.007949f
C446 B.n409 VSUBS 0.007949f
C447 B.n410 VSUBS 0.007949f
C448 B.n411 VSUBS 0.007949f
C449 B.n412 VSUBS 0.007949f
C450 B.n413 VSUBS 0.007949f
C451 B.n414 VSUBS 0.007949f
C452 B.n415 VSUBS 0.007949f
C453 B.n416 VSUBS 0.007949f
C454 B.n417 VSUBS 0.007949f
C455 B.n418 VSUBS 0.007949f
C456 B.n419 VSUBS 0.007949f
C457 B.n420 VSUBS 0.007949f
C458 B.n421 VSUBS 0.007949f
C459 B.n422 VSUBS 0.007949f
C460 B.n423 VSUBS 0.007949f
C461 B.n424 VSUBS 0.007949f
C462 B.n425 VSUBS 0.007949f
C463 B.n426 VSUBS 0.007949f
C464 B.n427 VSUBS 0.007949f
C465 B.n428 VSUBS 0.007949f
C466 B.n429 VSUBS 0.007949f
C467 B.n430 VSUBS 0.007949f
C468 B.n431 VSUBS 0.007949f
C469 B.n432 VSUBS 0.007949f
C470 B.n433 VSUBS 0.007949f
C471 B.n434 VSUBS 0.007949f
C472 B.n435 VSUBS 0.007949f
C473 B.n436 VSUBS 0.007949f
C474 B.n437 VSUBS 0.007949f
C475 B.n438 VSUBS 0.007949f
C476 B.n439 VSUBS 0.007949f
C477 B.n440 VSUBS 0.007949f
C478 B.n441 VSUBS 0.007949f
C479 B.n442 VSUBS 0.007949f
C480 B.n443 VSUBS 0.007949f
C481 B.n444 VSUBS 0.007949f
C482 B.n445 VSUBS 0.007949f
C483 B.n446 VSUBS 0.007949f
C484 B.n447 VSUBS 0.007949f
C485 B.n448 VSUBS 0.007949f
C486 B.n449 VSUBS 0.007949f
C487 B.n450 VSUBS 0.007949f
C488 B.n451 VSUBS 0.007482f
C489 B.n452 VSUBS 0.018418f
C490 B.n453 VSUBS 0.004442f
C491 B.n454 VSUBS 0.007949f
C492 B.n455 VSUBS 0.007949f
C493 B.n456 VSUBS 0.007949f
C494 B.n457 VSUBS 0.007949f
C495 B.n458 VSUBS 0.007949f
C496 B.n459 VSUBS 0.007949f
C497 B.n460 VSUBS 0.007949f
C498 B.n461 VSUBS 0.007949f
C499 B.n462 VSUBS 0.007949f
C500 B.n463 VSUBS 0.007949f
C501 B.n464 VSUBS 0.007949f
C502 B.n465 VSUBS 0.007949f
C503 B.t8 VSUBS 0.688862f
C504 B.t7 VSUBS 0.714768f
C505 B.t6 VSUBS 2.65641f
C506 B.n466 VSUBS 0.408423f
C507 B.n467 VSUBS 0.08335f
C508 B.n468 VSUBS 0.018418f
C509 B.n469 VSUBS 0.004442f
C510 B.n470 VSUBS 0.007949f
C511 B.n471 VSUBS 0.007949f
C512 B.n472 VSUBS 0.007949f
C513 B.n473 VSUBS 0.007949f
C514 B.n474 VSUBS 0.007949f
C515 B.n475 VSUBS 0.007949f
C516 B.n476 VSUBS 0.007949f
C517 B.n477 VSUBS 0.007949f
C518 B.n478 VSUBS 0.007949f
C519 B.n479 VSUBS 0.007949f
C520 B.n480 VSUBS 0.007949f
C521 B.n481 VSUBS 0.007949f
C522 B.n482 VSUBS 0.007949f
C523 B.n483 VSUBS 0.007949f
C524 B.n484 VSUBS 0.007949f
C525 B.n485 VSUBS 0.007949f
C526 B.n486 VSUBS 0.007949f
C527 B.n487 VSUBS 0.007949f
C528 B.n488 VSUBS 0.007949f
C529 B.n489 VSUBS 0.007949f
C530 B.n490 VSUBS 0.007949f
C531 B.n491 VSUBS 0.007949f
C532 B.n492 VSUBS 0.007949f
C533 B.n493 VSUBS 0.007949f
C534 B.n494 VSUBS 0.007949f
C535 B.n495 VSUBS 0.007949f
C536 B.n496 VSUBS 0.007949f
C537 B.n497 VSUBS 0.007949f
C538 B.n498 VSUBS 0.007949f
C539 B.n499 VSUBS 0.007949f
C540 B.n500 VSUBS 0.007949f
C541 B.n501 VSUBS 0.007949f
C542 B.n502 VSUBS 0.007949f
C543 B.n503 VSUBS 0.007949f
C544 B.n504 VSUBS 0.007949f
C545 B.n505 VSUBS 0.007949f
C546 B.n506 VSUBS 0.007949f
C547 B.n507 VSUBS 0.007949f
C548 B.n508 VSUBS 0.007949f
C549 B.n509 VSUBS 0.007949f
C550 B.n510 VSUBS 0.007949f
C551 B.n511 VSUBS 0.007949f
C552 B.n512 VSUBS 0.007949f
C553 B.n513 VSUBS 0.007949f
C554 B.n514 VSUBS 0.007949f
C555 B.n515 VSUBS 0.007949f
C556 B.n516 VSUBS 0.007949f
C557 B.n517 VSUBS 0.007949f
C558 B.n518 VSUBS 0.007949f
C559 B.n519 VSUBS 0.007949f
C560 B.n520 VSUBS 0.007949f
C561 B.n521 VSUBS 0.007949f
C562 B.n522 VSUBS 0.007949f
C563 B.n523 VSUBS 0.007949f
C564 B.n524 VSUBS 0.007949f
C565 B.n525 VSUBS 0.007949f
C566 B.n526 VSUBS 0.007949f
C567 B.n527 VSUBS 0.007949f
C568 B.n528 VSUBS 0.007949f
C569 B.n529 VSUBS 0.007949f
C570 B.n530 VSUBS 0.007949f
C571 B.n531 VSUBS 0.007949f
C572 B.n532 VSUBS 0.007949f
C573 B.n533 VSUBS 0.007949f
C574 B.n534 VSUBS 0.007949f
C575 B.n535 VSUBS 0.007949f
C576 B.n536 VSUBS 0.007949f
C577 B.n537 VSUBS 0.007949f
C578 B.n538 VSUBS 0.007949f
C579 B.n539 VSUBS 0.007949f
C580 B.n540 VSUBS 0.007949f
C581 B.n541 VSUBS 0.007949f
C582 B.n542 VSUBS 0.007949f
C583 B.n543 VSUBS 0.007949f
C584 B.n544 VSUBS 0.007949f
C585 B.n545 VSUBS 0.007949f
C586 B.n546 VSUBS 0.007949f
C587 B.n547 VSUBS 0.007949f
C588 B.n548 VSUBS 0.007949f
C589 B.n549 VSUBS 0.007949f
C590 B.n550 VSUBS 0.007949f
C591 B.n551 VSUBS 0.007949f
C592 B.n552 VSUBS 0.007949f
C593 B.n553 VSUBS 0.007949f
C594 B.n554 VSUBS 0.007949f
C595 B.n555 VSUBS 0.007949f
C596 B.n556 VSUBS 0.007949f
C597 B.n557 VSUBS 0.007949f
C598 B.n558 VSUBS 0.016845f
C599 B.n559 VSUBS 0.018226f
C600 B.n560 VSUBS 0.017197f
C601 B.n561 VSUBS 0.007949f
C602 B.n562 VSUBS 0.007949f
C603 B.n563 VSUBS 0.007949f
C604 B.n564 VSUBS 0.007949f
C605 B.n565 VSUBS 0.007949f
C606 B.n566 VSUBS 0.007949f
C607 B.n567 VSUBS 0.007949f
C608 B.n568 VSUBS 0.007949f
C609 B.n569 VSUBS 0.007949f
C610 B.n570 VSUBS 0.007949f
C611 B.n571 VSUBS 0.007949f
C612 B.n572 VSUBS 0.007949f
C613 B.n573 VSUBS 0.007949f
C614 B.n574 VSUBS 0.007949f
C615 B.n575 VSUBS 0.007949f
C616 B.n576 VSUBS 0.007949f
C617 B.n577 VSUBS 0.007949f
C618 B.n578 VSUBS 0.007949f
C619 B.n579 VSUBS 0.007949f
C620 B.n580 VSUBS 0.007949f
C621 B.n581 VSUBS 0.007949f
C622 B.n582 VSUBS 0.007949f
C623 B.n583 VSUBS 0.007949f
C624 B.n584 VSUBS 0.007949f
C625 B.n585 VSUBS 0.007949f
C626 B.n586 VSUBS 0.007949f
C627 B.n587 VSUBS 0.007949f
C628 B.n588 VSUBS 0.007949f
C629 B.n589 VSUBS 0.007949f
C630 B.n590 VSUBS 0.007949f
C631 B.n591 VSUBS 0.007949f
C632 B.n592 VSUBS 0.007949f
C633 B.n593 VSUBS 0.007949f
C634 B.n594 VSUBS 0.007949f
C635 B.n595 VSUBS 0.007949f
C636 B.n596 VSUBS 0.007949f
C637 B.n597 VSUBS 0.007949f
C638 B.n598 VSUBS 0.007949f
C639 B.n599 VSUBS 0.007949f
C640 B.n600 VSUBS 0.007949f
C641 B.n601 VSUBS 0.007949f
C642 B.n602 VSUBS 0.007949f
C643 B.n603 VSUBS 0.007949f
C644 B.n604 VSUBS 0.007949f
C645 B.n605 VSUBS 0.007949f
C646 B.n606 VSUBS 0.007949f
C647 B.n607 VSUBS 0.007949f
C648 B.n608 VSUBS 0.007949f
C649 B.n609 VSUBS 0.007949f
C650 B.n610 VSUBS 0.007949f
C651 B.n611 VSUBS 0.007949f
C652 B.n612 VSUBS 0.007949f
C653 B.n613 VSUBS 0.007949f
C654 B.n614 VSUBS 0.007949f
C655 B.n615 VSUBS 0.007949f
C656 B.n616 VSUBS 0.007949f
C657 B.n617 VSUBS 0.007949f
C658 B.n618 VSUBS 0.007949f
C659 B.n619 VSUBS 0.007949f
C660 B.n620 VSUBS 0.007949f
C661 B.n621 VSUBS 0.007949f
C662 B.n622 VSUBS 0.007949f
C663 B.n623 VSUBS 0.007949f
C664 B.n624 VSUBS 0.007949f
C665 B.n625 VSUBS 0.007949f
C666 B.n626 VSUBS 0.007949f
C667 B.n627 VSUBS 0.007949f
C668 B.n628 VSUBS 0.007949f
C669 B.n629 VSUBS 0.007949f
C670 B.n630 VSUBS 0.007949f
C671 B.n631 VSUBS 0.007949f
C672 B.n632 VSUBS 0.007949f
C673 B.n633 VSUBS 0.007949f
C674 B.n634 VSUBS 0.007949f
C675 B.n635 VSUBS 0.007949f
C676 B.n636 VSUBS 0.007949f
C677 B.n637 VSUBS 0.007949f
C678 B.n638 VSUBS 0.007949f
C679 B.n639 VSUBS 0.007949f
C680 B.n640 VSUBS 0.007949f
C681 B.n641 VSUBS 0.007949f
C682 B.n642 VSUBS 0.007949f
C683 B.n643 VSUBS 0.007949f
C684 B.n644 VSUBS 0.007949f
C685 B.n645 VSUBS 0.007949f
C686 B.n646 VSUBS 0.007949f
C687 B.n647 VSUBS 0.007949f
C688 B.n648 VSUBS 0.007949f
C689 B.n649 VSUBS 0.007949f
C690 B.n650 VSUBS 0.007949f
C691 B.n651 VSUBS 0.007949f
C692 B.n652 VSUBS 0.007949f
C693 B.n653 VSUBS 0.007949f
C694 B.n654 VSUBS 0.007949f
C695 B.n655 VSUBS 0.007949f
C696 B.n656 VSUBS 0.007949f
C697 B.n657 VSUBS 0.007949f
C698 B.n658 VSUBS 0.007949f
C699 B.n659 VSUBS 0.007949f
C700 B.n660 VSUBS 0.007949f
C701 B.n661 VSUBS 0.007949f
C702 B.n662 VSUBS 0.007949f
C703 B.n663 VSUBS 0.007949f
C704 B.n664 VSUBS 0.007949f
C705 B.n665 VSUBS 0.007949f
C706 B.n666 VSUBS 0.007949f
C707 B.n667 VSUBS 0.007949f
C708 B.n668 VSUBS 0.007949f
C709 B.n669 VSUBS 0.007949f
C710 B.n670 VSUBS 0.007949f
C711 B.n671 VSUBS 0.007949f
C712 B.n672 VSUBS 0.007949f
C713 B.n673 VSUBS 0.007949f
C714 B.n674 VSUBS 0.007949f
C715 B.n675 VSUBS 0.007949f
C716 B.n676 VSUBS 0.007949f
C717 B.n677 VSUBS 0.007949f
C718 B.n678 VSUBS 0.007949f
C719 B.n679 VSUBS 0.007949f
C720 B.n680 VSUBS 0.007949f
C721 B.n681 VSUBS 0.007949f
C722 B.n682 VSUBS 0.007949f
C723 B.n683 VSUBS 0.007949f
C724 B.n684 VSUBS 0.007949f
C725 B.n685 VSUBS 0.007949f
C726 B.n686 VSUBS 0.007949f
C727 B.n687 VSUBS 0.007949f
C728 B.n688 VSUBS 0.007949f
C729 B.n689 VSUBS 0.007949f
C730 B.n690 VSUBS 0.007949f
C731 B.n691 VSUBS 0.007949f
C732 B.n692 VSUBS 0.007949f
C733 B.n693 VSUBS 0.007949f
C734 B.n694 VSUBS 0.007949f
C735 B.n695 VSUBS 0.007949f
C736 B.n696 VSUBS 0.007949f
C737 B.n697 VSUBS 0.007949f
C738 B.n698 VSUBS 0.007949f
C739 B.n699 VSUBS 0.007949f
C740 B.n700 VSUBS 0.007949f
C741 B.n701 VSUBS 0.007949f
C742 B.n702 VSUBS 0.007949f
C743 B.n703 VSUBS 0.007949f
C744 B.n704 VSUBS 0.007949f
C745 B.n705 VSUBS 0.007949f
C746 B.n706 VSUBS 0.007949f
C747 B.n707 VSUBS 0.007949f
C748 B.n708 VSUBS 0.007949f
C749 B.n709 VSUBS 0.007949f
C750 B.n710 VSUBS 0.007949f
C751 B.n711 VSUBS 0.007949f
C752 B.n712 VSUBS 0.007949f
C753 B.n713 VSUBS 0.007949f
C754 B.n714 VSUBS 0.007949f
C755 B.n715 VSUBS 0.007949f
C756 B.n716 VSUBS 0.007949f
C757 B.n717 VSUBS 0.007949f
C758 B.n718 VSUBS 0.007949f
C759 B.n719 VSUBS 0.007949f
C760 B.n720 VSUBS 0.007949f
C761 B.n721 VSUBS 0.007949f
C762 B.n722 VSUBS 0.007949f
C763 B.n723 VSUBS 0.007949f
C764 B.n724 VSUBS 0.007949f
C765 B.n725 VSUBS 0.007949f
C766 B.n726 VSUBS 0.007949f
C767 B.n727 VSUBS 0.007949f
C768 B.n728 VSUBS 0.007949f
C769 B.n729 VSUBS 0.007949f
C770 B.n730 VSUBS 0.007949f
C771 B.n731 VSUBS 0.007949f
C772 B.n732 VSUBS 0.007949f
C773 B.n733 VSUBS 0.007949f
C774 B.n734 VSUBS 0.007949f
C775 B.n735 VSUBS 0.007949f
C776 B.n736 VSUBS 0.007949f
C777 B.n737 VSUBS 0.007949f
C778 B.n738 VSUBS 0.007949f
C779 B.n739 VSUBS 0.007949f
C780 B.n740 VSUBS 0.007949f
C781 B.n741 VSUBS 0.007949f
C782 B.n742 VSUBS 0.007949f
C783 B.n743 VSUBS 0.007949f
C784 B.n744 VSUBS 0.007949f
C785 B.n745 VSUBS 0.007949f
C786 B.n746 VSUBS 0.007949f
C787 B.n747 VSUBS 0.007949f
C788 B.n748 VSUBS 0.007949f
C789 B.n749 VSUBS 0.007949f
C790 B.n750 VSUBS 0.007949f
C791 B.n751 VSUBS 0.007949f
C792 B.n752 VSUBS 0.007949f
C793 B.n753 VSUBS 0.007949f
C794 B.n754 VSUBS 0.007949f
C795 B.n755 VSUBS 0.007949f
C796 B.n756 VSUBS 0.017197f
C797 B.n757 VSUBS 0.017874f
C798 B.n758 VSUBS 0.017874f
C799 B.n759 VSUBS 0.007949f
C800 B.n760 VSUBS 0.007949f
C801 B.n761 VSUBS 0.007949f
C802 B.n762 VSUBS 0.007949f
C803 B.n763 VSUBS 0.007949f
C804 B.n764 VSUBS 0.007949f
C805 B.n765 VSUBS 0.007949f
C806 B.n766 VSUBS 0.007949f
C807 B.n767 VSUBS 0.007949f
C808 B.n768 VSUBS 0.007949f
C809 B.n769 VSUBS 0.007949f
C810 B.n770 VSUBS 0.007949f
C811 B.n771 VSUBS 0.007949f
C812 B.n772 VSUBS 0.007949f
C813 B.n773 VSUBS 0.007949f
C814 B.n774 VSUBS 0.007949f
C815 B.n775 VSUBS 0.007949f
C816 B.n776 VSUBS 0.007949f
C817 B.n777 VSUBS 0.007949f
C818 B.n778 VSUBS 0.007949f
C819 B.n779 VSUBS 0.007949f
C820 B.n780 VSUBS 0.007949f
C821 B.n781 VSUBS 0.007949f
C822 B.n782 VSUBS 0.007949f
C823 B.n783 VSUBS 0.007949f
C824 B.n784 VSUBS 0.007949f
C825 B.n785 VSUBS 0.007949f
C826 B.n786 VSUBS 0.007949f
C827 B.n787 VSUBS 0.007949f
C828 B.n788 VSUBS 0.007949f
C829 B.n789 VSUBS 0.007949f
C830 B.n790 VSUBS 0.007949f
C831 B.n791 VSUBS 0.007949f
C832 B.n792 VSUBS 0.007949f
C833 B.n793 VSUBS 0.007949f
C834 B.n794 VSUBS 0.007949f
C835 B.n795 VSUBS 0.007949f
C836 B.n796 VSUBS 0.007949f
C837 B.n797 VSUBS 0.007949f
C838 B.n798 VSUBS 0.007949f
C839 B.n799 VSUBS 0.007949f
C840 B.n800 VSUBS 0.007949f
C841 B.n801 VSUBS 0.007949f
C842 B.n802 VSUBS 0.007949f
C843 B.n803 VSUBS 0.007949f
C844 B.n804 VSUBS 0.007949f
C845 B.n805 VSUBS 0.007949f
C846 B.n806 VSUBS 0.007949f
C847 B.n807 VSUBS 0.007949f
C848 B.n808 VSUBS 0.007949f
C849 B.n809 VSUBS 0.007949f
C850 B.n810 VSUBS 0.007949f
C851 B.n811 VSUBS 0.007949f
C852 B.n812 VSUBS 0.007949f
C853 B.n813 VSUBS 0.007949f
C854 B.n814 VSUBS 0.007949f
C855 B.n815 VSUBS 0.007949f
C856 B.n816 VSUBS 0.007949f
C857 B.n817 VSUBS 0.007949f
C858 B.n818 VSUBS 0.007949f
C859 B.n819 VSUBS 0.007949f
C860 B.n820 VSUBS 0.007949f
C861 B.n821 VSUBS 0.007949f
C862 B.n822 VSUBS 0.007949f
C863 B.n823 VSUBS 0.007949f
C864 B.n824 VSUBS 0.007949f
C865 B.n825 VSUBS 0.007949f
C866 B.n826 VSUBS 0.007949f
C867 B.n827 VSUBS 0.007949f
C868 B.n828 VSUBS 0.007949f
C869 B.n829 VSUBS 0.007949f
C870 B.n830 VSUBS 0.007949f
C871 B.n831 VSUBS 0.007949f
C872 B.n832 VSUBS 0.007949f
C873 B.n833 VSUBS 0.007949f
C874 B.n834 VSUBS 0.007949f
C875 B.n835 VSUBS 0.007949f
C876 B.n836 VSUBS 0.007949f
C877 B.n837 VSUBS 0.007949f
C878 B.n838 VSUBS 0.007949f
C879 B.n839 VSUBS 0.007949f
C880 B.n840 VSUBS 0.007949f
C881 B.n841 VSUBS 0.007949f
C882 B.n842 VSUBS 0.007949f
C883 B.n843 VSUBS 0.007949f
C884 B.n844 VSUBS 0.007949f
C885 B.n845 VSUBS 0.007482f
C886 B.n846 VSUBS 0.018418f
C887 B.n847 VSUBS 0.004442f
C888 B.n848 VSUBS 0.007949f
C889 B.n849 VSUBS 0.007949f
C890 B.n850 VSUBS 0.007949f
C891 B.n851 VSUBS 0.007949f
C892 B.n852 VSUBS 0.007949f
C893 B.n853 VSUBS 0.007949f
C894 B.n854 VSUBS 0.007949f
C895 B.n855 VSUBS 0.007949f
C896 B.n856 VSUBS 0.007949f
C897 B.n857 VSUBS 0.007949f
C898 B.n858 VSUBS 0.007949f
C899 B.n859 VSUBS 0.007949f
C900 B.n860 VSUBS 0.004442f
C901 B.n861 VSUBS 0.007949f
C902 B.n862 VSUBS 0.007949f
C903 B.n863 VSUBS 0.007482f
C904 B.n864 VSUBS 0.007949f
C905 B.n865 VSUBS 0.007949f
C906 B.n866 VSUBS 0.007949f
C907 B.n867 VSUBS 0.007949f
C908 B.n868 VSUBS 0.007949f
C909 B.n869 VSUBS 0.007949f
C910 B.n870 VSUBS 0.007949f
C911 B.n871 VSUBS 0.007949f
C912 B.n872 VSUBS 0.007949f
C913 B.n873 VSUBS 0.007949f
C914 B.n874 VSUBS 0.007949f
C915 B.n875 VSUBS 0.007949f
C916 B.n876 VSUBS 0.007949f
C917 B.n877 VSUBS 0.007949f
C918 B.n878 VSUBS 0.007949f
C919 B.n879 VSUBS 0.007949f
C920 B.n880 VSUBS 0.007949f
C921 B.n881 VSUBS 0.007949f
C922 B.n882 VSUBS 0.007949f
C923 B.n883 VSUBS 0.007949f
C924 B.n884 VSUBS 0.007949f
C925 B.n885 VSUBS 0.007949f
C926 B.n886 VSUBS 0.007949f
C927 B.n887 VSUBS 0.007949f
C928 B.n888 VSUBS 0.007949f
C929 B.n889 VSUBS 0.007949f
C930 B.n890 VSUBS 0.007949f
C931 B.n891 VSUBS 0.007949f
C932 B.n892 VSUBS 0.007949f
C933 B.n893 VSUBS 0.007949f
C934 B.n894 VSUBS 0.007949f
C935 B.n895 VSUBS 0.007949f
C936 B.n896 VSUBS 0.007949f
C937 B.n897 VSUBS 0.007949f
C938 B.n898 VSUBS 0.007949f
C939 B.n899 VSUBS 0.007949f
C940 B.n900 VSUBS 0.007949f
C941 B.n901 VSUBS 0.007949f
C942 B.n902 VSUBS 0.007949f
C943 B.n903 VSUBS 0.007949f
C944 B.n904 VSUBS 0.007949f
C945 B.n905 VSUBS 0.007949f
C946 B.n906 VSUBS 0.007949f
C947 B.n907 VSUBS 0.007949f
C948 B.n908 VSUBS 0.007949f
C949 B.n909 VSUBS 0.007949f
C950 B.n910 VSUBS 0.007949f
C951 B.n911 VSUBS 0.007949f
C952 B.n912 VSUBS 0.007949f
C953 B.n913 VSUBS 0.007949f
C954 B.n914 VSUBS 0.007949f
C955 B.n915 VSUBS 0.007949f
C956 B.n916 VSUBS 0.007949f
C957 B.n917 VSUBS 0.007949f
C958 B.n918 VSUBS 0.007949f
C959 B.n919 VSUBS 0.007949f
C960 B.n920 VSUBS 0.007949f
C961 B.n921 VSUBS 0.007949f
C962 B.n922 VSUBS 0.007949f
C963 B.n923 VSUBS 0.007949f
C964 B.n924 VSUBS 0.007949f
C965 B.n925 VSUBS 0.007949f
C966 B.n926 VSUBS 0.007949f
C967 B.n927 VSUBS 0.007949f
C968 B.n928 VSUBS 0.007949f
C969 B.n929 VSUBS 0.007949f
C970 B.n930 VSUBS 0.007949f
C971 B.n931 VSUBS 0.007949f
C972 B.n932 VSUBS 0.007949f
C973 B.n933 VSUBS 0.007949f
C974 B.n934 VSUBS 0.007949f
C975 B.n935 VSUBS 0.007949f
C976 B.n936 VSUBS 0.007949f
C977 B.n937 VSUBS 0.007949f
C978 B.n938 VSUBS 0.007949f
C979 B.n939 VSUBS 0.007949f
C980 B.n940 VSUBS 0.007949f
C981 B.n941 VSUBS 0.007949f
C982 B.n942 VSUBS 0.007949f
C983 B.n943 VSUBS 0.007949f
C984 B.n944 VSUBS 0.007949f
C985 B.n945 VSUBS 0.007949f
C986 B.n946 VSUBS 0.007949f
C987 B.n947 VSUBS 0.007949f
C988 B.n948 VSUBS 0.007949f
C989 B.n949 VSUBS 0.017874f
C990 B.n950 VSUBS 0.017874f
C991 B.n951 VSUBS 0.017197f
C992 B.n952 VSUBS 0.007949f
C993 B.n953 VSUBS 0.007949f
C994 B.n954 VSUBS 0.007949f
C995 B.n955 VSUBS 0.007949f
C996 B.n956 VSUBS 0.007949f
C997 B.n957 VSUBS 0.007949f
C998 B.n958 VSUBS 0.007949f
C999 B.n959 VSUBS 0.007949f
C1000 B.n960 VSUBS 0.007949f
C1001 B.n961 VSUBS 0.007949f
C1002 B.n962 VSUBS 0.007949f
C1003 B.n963 VSUBS 0.007949f
C1004 B.n964 VSUBS 0.007949f
C1005 B.n965 VSUBS 0.007949f
C1006 B.n966 VSUBS 0.007949f
C1007 B.n967 VSUBS 0.007949f
C1008 B.n968 VSUBS 0.007949f
C1009 B.n969 VSUBS 0.007949f
C1010 B.n970 VSUBS 0.007949f
C1011 B.n971 VSUBS 0.007949f
C1012 B.n972 VSUBS 0.007949f
C1013 B.n973 VSUBS 0.007949f
C1014 B.n974 VSUBS 0.007949f
C1015 B.n975 VSUBS 0.007949f
C1016 B.n976 VSUBS 0.007949f
C1017 B.n977 VSUBS 0.007949f
C1018 B.n978 VSUBS 0.007949f
C1019 B.n979 VSUBS 0.007949f
C1020 B.n980 VSUBS 0.007949f
C1021 B.n981 VSUBS 0.007949f
C1022 B.n982 VSUBS 0.007949f
C1023 B.n983 VSUBS 0.007949f
C1024 B.n984 VSUBS 0.007949f
C1025 B.n985 VSUBS 0.007949f
C1026 B.n986 VSUBS 0.007949f
C1027 B.n987 VSUBS 0.007949f
C1028 B.n988 VSUBS 0.007949f
C1029 B.n989 VSUBS 0.007949f
C1030 B.n990 VSUBS 0.007949f
C1031 B.n991 VSUBS 0.007949f
C1032 B.n992 VSUBS 0.007949f
C1033 B.n993 VSUBS 0.007949f
C1034 B.n994 VSUBS 0.007949f
C1035 B.n995 VSUBS 0.007949f
C1036 B.n996 VSUBS 0.007949f
C1037 B.n997 VSUBS 0.007949f
C1038 B.n998 VSUBS 0.007949f
C1039 B.n999 VSUBS 0.007949f
C1040 B.n1000 VSUBS 0.007949f
C1041 B.n1001 VSUBS 0.007949f
C1042 B.n1002 VSUBS 0.007949f
C1043 B.n1003 VSUBS 0.007949f
C1044 B.n1004 VSUBS 0.007949f
C1045 B.n1005 VSUBS 0.007949f
C1046 B.n1006 VSUBS 0.007949f
C1047 B.n1007 VSUBS 0.007949f
C1048 B.n1008 VSUBS 0.007949f
C1049 B.n1009 VSUBS 0.007949f
C1050 B.n1010 VSUBS 0.007949f
C1051 B.n1011 VSUBS 0.007949f
C1052 B.n1012 VSUBS 0.007949f
C1053 B.n1013 VSUBS 0.007949f
C1054 B.n1014 VSUBS 0.007949f
C1055 B.n1015 VSUBS 0.007949f
C1056 B.n1016 VSUBS 0.007949f
C1057 B.n1017 VSUBS 0.007949f
C1058 B.n1018 VSUBS 0.007949f
C1059 B.n1019 VSUBS 0.007949f
C1060 B.n1020 VSUBS 0.007949f
C1061 B.n1021 VSUBS 0.007949f
C1062 B.n1022 VSUBS 0.007949f
C1063 B.n1023 VSUBS 0.007949f
C1064 B.n1024 VSUBS 0.007949f
C1065 B.n1025 VSUBS 0.007949f
C1066 B.n1026 VSUBS 0.007949f
C1067 B.n1027 VSUBS 0.007949f
C1068 B.n1028 VSUBS 0.007949f
C1069 B.n1029 VSUBS 0.007949f
C1070 B.n1030 VSUBS 0.007949f
C1071 B.n1031 VSUBS 0.007949f
C1072 B.n1032 VSUBS 0.007949f
C1073 B.n1033 VSUBS 0.007949f
C1074 B.n1034 VSUBS 0.007949f
C1075 B.n1035 VSUBS 0.007949f
C1076 B.n1036 VSUBS 0.007949f
C1077 B.n1037 VSUBS 0.007949f
C1078 B.n1038 VSUBS 0.007949f
C1079 B.n1039 VSUBS 0.007949f
C1080 B.n1040 VSUBS 0.007949f
C1081 B.n1041 VSUBS 0.007949f
C1082 B.n1042 VSUBS 0.007949f
C1083 B.n1043 VSUBS 0.007949f
C1084 B.n1044 VSUBS 0.007949f
C1085 B.n1045 VSUBS 0.007949f
C1086 B.n1046 VSUBS 0.007949f
C1087 B.n1047 VSUBS 0.010374f
C1088 B.n1048 VSUBS 0.01105f
C1089 B.n1049 VSUBS 0.021975f
C1090 VDD1.t7 VSUBS 4.41373f
C1091 VDD1.t2 VSUBS 0.40544f
C1092 VDD1.t6 VSUBS 0.40544f
C1093 VDD1.n0 VSUBS 3.37543f
C1094 VDD1.n1 VSUBS 1.77255f
C1095 VDD1.t1 VSUBS 4.41373f
C1096 VDD1.t4 VSUBS 0.40544f
C1097 VDD1.t9 VSUBS 0.40544f
C1098 VDD1.n2 VSUBS 3.37543f
C1099 VDD1.n3 VSUBS 1.76314f
C1100 VDD1.t3 VSUBS 0.40544f
C1101 VDD1.t0 VSUBS 0.40544f
C1102 VDD1.n4 VSUBS 3.40383f
C1103 VDD1.n5 VSUBS 4.40073f
C1104 VDD1.t8 VSUBS 0.40544f
C1105 VDD1.t5 VSUBS 0.40544f
C1106 VDD1.n6 VSUBS 3.37542f
C1107 VDD1.n7 VSUBS 4.60553f
C1108 VP.t9 VSUBS 3.65044f
C1109 VP.n0 VSUBS 1.36704f
C1110 VP.n1 VSUBS 0.02538f
C1111 VP.n2 VSUBS 0.044486f
C1112 VP.n3 VSUBS 0.02538f
C1113 VP.t6 VSUBS 3.65044f
C1114 VP.n4 VSUBS 0.047302f
C1115 VP.n5 VSUBS 0.02538f
C1116 VP.n6 VSUBS 0.047302f
C1117 VP.n7 VSUBS 0.02538f
C1118 VP.t0 VSUBS 3.65044f
C1119 VP.n8 VSUBS 0.025635f
C1120 VP.n9 VSUBS 0.02538f
C1121 VP.t5 VSUBS 3.65044f
C1122 VP.n10 VSUBS 1.26316f
C1123 VP.n11 VSUBS 0.02538f
C1124 VP.n12 VSUBS 0.027718f
C1125 VP.n13 VSUBS 0.040963f
C1126 VP.t8 VSUBS 3.65044f
C1127 VP.t4 VSUBS 3.65044f
C1128 VP.n14 VSUBS 1.36704f
C1129 VP.n15 VSUBS 0.02538f
C1130 VP.n16 VSUBS 0.044486f
C1131 VP.n17 VSUBS 0.02538f
C1132 VP.t1 VSUBS 3.65044f
C1133 VP.n18 VSUBS 0.047302f
C1134 VP.n19 VSUBS 0.02538f
C1135 VP.n20 VSUBS 0.047302f
C1136 VP.n21 VSUBS 0.02538f
C1137 VP.t3 VSUBS 3.65044f
C1138 VP.n22 VSUBS 0.025635f
C1139 VP.n23 VSUBS 0.02538f
C1140 VP.t7 VSUBS 3.65044f
C1141 VP.n24 VSUBS 1.34217f
C1142 VP.t2 VSUBS 3.90312f
C1143 VP.n25 VSUBS 1.30888f
C1144 VP.n26 VSUBS 0.270118f
C1145 VP.n27 VSUBS 0.035159f
C1146 VP.n28 VSUBS 0.047302f
C1147 VP.n29 VSUBS 0.045565f
C1148 VP.n30 VSUBS 0.02538f
C1149 VP.n31 VSUBS 0.02538f
C1150 VP.n32 VSUBS 0.02538f
C1151 VP.n33 VSUBS 0.050203f
C1152 VP.n34 VSUBS 0.047302f
C1153 VP.n35 VSUBS 1.28711f
C1154 VP.n36 VSUBS 0.02538f
C1155 VP.n37 VSUBS 0.02538f
C1156 VP.n38 VSUBS 0.02538f
C1157 VP.n39 VSUBS 0.050203f
C1158 VP.n40 VSUBS 0.025635f
C1159 VP.n41 VSUBS 0.045565f
C1160 VP.n42 VSUBS 0.02538f
C1161 VP.n43 VSUBS 0.02538f
C1162 VP.n44 VSUBS 0.02538f
C1163 VP.n45 VSUBS 0.035159f
C1164 VP.n46 VSUBS 1.26316f
C1165 VP.n47 VSUBS 0.036093f
C1166 VP.n48 VSUBS 0.047302f
C1167 VP.n49 VSUBS 0.02538f
C1168 VP.n50 VSUBS 0.02538f
C1169 VP.n51 VSUBS 0.02538f
C1170 VP.n52 VSUBS 0.027718f
C1171 VP.n53 VSUBS 0.049199f
C1172 VP.n54 VSUBS 0.046368f
C1173 VP.n55 VSUBS 0.040963f
C1174 VP.n56 VSUBS 1.82306f
C1175 VP.n57 VSUBS 1.8384f
C1176 VP.n58 VSUBS 1.36704f
C1177 VP.n59 VSUBS 0.046368f
C1178 VP.n60 VSUBS 0.049199f
C1179 VP.n61 VSUBS 0.02538f
C1180 VP.n62 VSUBS 0.02538f
C1181 VP.n63 VSUBS 0.02538f
C1182 VP.n64 VSUBS 0.044486f
C1183 VP.n65 VSUBS 0.047302f
C1184 VP.n66 VSUBS 0.036093f
C1185 VP.n67 VSUBS 0.02538f
C1186 VP.n68 VSUBS 0.02538f
C1187 VP.n69 VSUBS 0.035159f
C1188 VP.n70 VSUBS 0.047302f
C1189 VP.n71 VSUBS 0.045565f
C1190 VP.n72 VSUBS 0.02538f
C1191 VP.n73 VSUBS 0.02538f
C1192 VP.n74 VSUBS 0.02538f
C1193 VP.n75 VSUBS 0.050203f
C1194 VP.n76 VSUBS 0.047302f
C1195 VP.n77 VSUBS 1.28711f
C1196 VP.n78 VSUBS 0.02538f
C1197 VP.n79 VSUBS 0.02538f
C1198 VP.n80 VSUBS 0.02538f
C1199 VP.n81 VSUBS 0.050203f
C1200 VP.n82 VSUBS 0.025635f
C1201 VP.n83 VSUBS 0.045565f
C1202 VP.n84 VSUBS 0.02538f
C1203 VP.n85 VSUBS 0.02538f
C1204 VP.n86 VSUBS 0.02538f
C1205 VP.n87 VSUBS 0.035159f
C1206 VP.n88 VSUBS 1.26316f
C1207 VP.n89 VSUBS 0.036093f
C1208 VP.n90 VSUBS 0.047302f
C1209 VP.n91 VSUBS 0.02538f
C1210 VP.n92 VSUBS 0.02538f
C1211 VP.n93 VSUBS 0.02538f
C1212 VP.n94 VSUBS 0.027718f
C1213 VP.n95 VSUBS 0.049199f
C1214 VP.n96 VSUBS 0.046368f
C1215 VP.n97 VSUBS 0.040963f
C1216 VP.n98 VSUBS 0.047874f
C1217 VTAIL.t13 VSUBS 0.391193f
C1218 VTAIL.t15 VSUBS 0.391193f
C1219 VTAIL.n0 VSUBS 3.09277f
C1220 VTAIL.n1 VSUBS 1.01892f
C1221 VTAIL.t2 VSUBS 4.03734f
C1222 VTAIL.n2 VSUBS 1.19807f
C1223 VTAIL.t8 VSUBS 0.391193f
C1224 VTAIL.t1 VSUBS 0.391193f
C1225 VTAIL.n3 VSUBS 3.09277f
C1226 VTAIL.n4 VSUBS 1.158f
C1227 VTAIL.t3 VSUBS 0.391193f
C1228 VTAIL.t6 VSUBS 0.391193f
C1229 VTAIL.n5 VSUBS 3.09277f
C1230 VTAIL.n6 VSUBS 3.15524f
C1231 VTAIL.t18 VSUBS 0.391193f
C1232 VTAIL.t17 VSUBS 0.391193f
C1233 VTAIL.n7 VSUBS 3.09278f
C1234 VTAIL.n8 VSUBS 3.15524f
C1235 VTAIL.t10 VSUBS 0.391193f
C1236 VTAIL.t19 VSUBS 0.391193f
C1237 VTAIL.n9 VSUBS 3.09278f
C1238 VTAIL.n10 VSUBS 1.158f
C1239 VTAIL.t16 VSUBS 4.03734f
C1240 VTAIL.n11 VSUBS 1.19806f
C1241 VTAIL.t7 VSUBS 0.391193f
C1242 VTAIL.t4 VSUBS 0.391193f
C1243 VTAIL.n12 VSUBS 3.09278f
C1244 VTAIL.n13 VSUBS 1.07574f
C1245 VTAIL.t5 VSUBS 0.391193f
C1246 VTAIL.t9 VSUBS 0.391193f
C1247 VTAIL.n14 VSUBS 3.09278f
C1248 VTAIL.n15 VSUBS 1.158f
C1249 VTAIL.t0 VSUBS 4.03734f
C1250 VTAIL.n16 VSUBS 3.02964f
C1251 VTAIL.t12 VSUBS 4.03734f
C1252 VTAIL.n17 VSUBS 3.02964f
C1253 VTAIL.t11 VSUBS 0.391193f
C1254 VTAIL.t14 VSUBS 0.391193f
C1255 VTAIL.n18 VSUBS 3.09277f
C1256 VTAIL.n19 VSUBS 0.96689f
C1257 VDD2.t9 VSUBS 4.41435f
C1258 VDD2.t5 VSUBS 0.405498f
C1259 VDD2.t7 VSUBS 0.405498f
C1260 VDD2.n0 VSUBS 3.37591f
C1261 VDD2.n1 VSUBS 1.76339f
C1262 VDD2.t4 VSUBS 0.405498f
C1263 VDD2.t8 VSUBS 0.405498f
C1264 VDD2.n2 VSUBS 3.40432f
C1265 VDD2.n3 VSUBS 4.24461f
C1266 VDD2.t2 VSUBS 4.37998f
C1267 VDD2.n4 VSUBS 4.57189f
C1268 VDD2.t1 VSUBS 0.405498f
C1269 VDD2.t6 VSUBS 0.405498f
C1270 VDD2.n5 VSUBS 3.37592f
C1271 VDD2.n6 VSUBS 0.881721f
C1272 VDD2.t3 VSUBS 0.405498f
C1273 VDD2.t0 VSUBS 0.405498f
C1274 VDD2.n7 VSUBS 3.40425f
C1275 VN.t7 VSUBS 3.42335f
C1276 VN.n0 VSUBS 1.282f
C1277 VN.n1 VSUBS 0.023801f
C1278 VN.n2 VSUBS 0.041719f
C1279 VN.n3 VSUBS 0.023801f
C1280 VN.t5 VSUBS 3.42335f
C1281 VN.n4 VSUBS 0.04436f
C1282 VN.n5 VSUBS 0.023801f
C1283 VN.n6 VSUBS 0.04436f
C1284 VN.n7 VSUBS 0.023801f
C1285 VN.t8 VSUBS 3.42335f
C1286 VN.n8 VSUBS 0.024041f
C1287 VN.n9 VSUBS 0.023801f
C1288 VN.t4 VSUBS 3.42335f
C1289 VN.n10 VSUBS 1.25868f
C1290 VN.t6 VSUBS 3.66031f
C1291 VN.n11 VSUBS 1.22746f
C1292 VN.n12 VSUBS 0.253314f
C1293 VN.n13 VSUBS 0.032971f
C1294 VN.n14 VSUBS 0.04436f
C1295 VN.n15 VSUBS 0.04273f
C1296 VN.n16 VSUBS 0.023801f
C1297 VN.n17 VSUBS 0.023801f
C1298 VN.n18 VSUBS 0.023801f
C1299 VN.n19 VSUBS 0.04708f
C1300 VN.n20 VSUBS 0.04436f
C1301 VN.n21 VSUBS 1.20704f
C1302 VN.n22 VSUBS 0.023801f
C1303 VN.n23 VSUBS 0.023801f
C1304 VN.n24 VSUBS 0.023801f
C1305 VN.n25 VSUBS 0.04708f
C1306 VN.n26 VSUBS 0.024041f
C1307 VN.n27 VSUBS 0.04273f
C1308 VN.n28 VSUBS 0.023801f
C1309 VN.n29 VSUBS 0.023801f
C1310 VN.n30 VSUBS 0.023801f
C1311 VN.n31 VSUBS 0.032971f
C1312 VN.n32 VSUBS 1.18458f
C1313 VN.n33 VSUBS 0.033847f
C1314 VN.n34 VSUBS 0.04436f
C1315 VN.n35 VSUBS 0.023801f
C1316 VN.n36 VSUBS 0.023801f
C1317 VN.n37 VSUBS 0.023801f
C1318 VN.n38 VSUBS 0.025994f
C1319 VN.n39 VSUBS 0.046138f
C1320 VN.n40 VSUBS 0.043484f
C1321 VN.n41 VSUBS 0.038415f
C1322 VN.n42 VSUBS 0.044896f
C1323 VN.t1 VSUBS 3.42335f
C1324 VN.n43 VSUBS 1.282f
C1325 VN.n44 VSUBS 0.023801f
C1326 VN.n45 VSUBS 0.041719f
C1327 VN.n46 VSUBS 0.023801f
C1328 VN.t2 VSUBS 3.42335f
C1329 VN.n47 VSUBS 0.04436f
C1330 VN.n48 VSUBS 0.023801f
C1331 VN.n49 VSUBS 0.04436f
C1332 VN.n50 VSUBS 0.023801f
C1333 VN.t9 VSUBS 3.42335f
C1334 VN.n51 VSUBS 0.024041f
C1335 VN.n52 VSUBS 0.023801f
C1336 VN.t0 VSUBS 3.42335f
C1337 VN.n53 VSUBS 1.25868f
C1338 VN.t3 VSUBS 3.66031f
C1339 VN.n54 VSUBS 1.22746f
C1340 VN.n55 VSUBS 0.253314f
C1341 VN.n56 VSUBS 0.032971f
C1342 VN.n57 VSUBS 0.04436f
C1343 VN.n58 VSUBS 0.04273f
C1344 VN.n59 VSUBS 0.023801f
C1345 VN.n60 VSUBS 0.023801f
C1346 VN.n61 VSUBS 0.023801f
C1347 VN.n62 VSUBS 0.04708f
C1348 VN.n63 VSUBS 0.04436f
C1349 VN.n64 VSUBS 1.20704f
C1350 VN.n65 VSUBS 0.023801f
C1351 VN.n66 VSUBS 0.023801f
C1352 VN.n67 VSUBS 0.023801f
C1353 VN.n68 VSUBS 0.04708f
C1354 VN.n69 VSUBS 0.024041f
C1355 VN.n70 VSUBS 0.04273f
C1356 VN.n71 VSUBS 0.023801f
C1357 VN.n72 VSUBS 0.023801f
C1358 VN.n73 VSUBS 0.023801f
C1359 VN.n74 VSUBS 0.032971f
C1360 VN.n75 VSUBS 1.18458f
C1361 VN.n76 VSUBS 0.033847f
C1362 VN.n77 VSUBS 0.04436f
C1363 VN.n78 VSUBS 0.023801f
C1364 VN.n79 VSUBS 0.023801f
C1365 VN.n80 VSUBS 0.023801f
C1366 VN.n81 VSUBS 0.025994f
C1367 VN.n82 VSUBS 0.046138f
C1368 VN.n83 VSUBS 0.043484f
C1369 VN.n84 VSUBS 0.038415f
C1370 VN.n85 VSUBS 1.71885f
.ends

