* NGSPICE file created from tg_sample_0004.ext - technology: sky130A

.subckt tg_sample_0004 VIN VGN VGP VSS VCC VOUT
X0 VIN.t7 VGP.t0 VOUT.t4 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.54
X1 VIN.t2 VGN.t0 VOUT.t2 VSS.t3 sky130_fd_pr__nfet_01v8 ad=2.3727 pd=14.71 as=2.3727 ps=14.71 w=14.38 l=2.98
X2 VOUT.t1 VGN.t1 VIN.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=2.3727 pd=14.71 as=5.6082 ps=29.54 w=14.38 l=2.98
X3 VIN.t6 VGP.t1 VOUT.t5 VCC.t2 sky130_fd_pr__pfet_01v8 ad=2.7495 pd=14.88 as=1.16325 ps=7.38 w=7.05 l=2.54
X4 VOUT.t0 VGN.t2 VIN.t0 VSS.t1 sky130_fd_pr__nfet_01v8 ad=2.3727 pd=14.71 as=2.3727 ps=14.71 w=14.38 l=2.98
X5 VIN.t3 VGN.t3 VOUT.t3 VSS.t0 sky130_fd_pr__nfet_01v8 ad=5.6082 pd=29.54 as=2.3727 ps=14.71 w=14.38 l=2.98
X6 VCC.t11 VCC.t8 VCC.t10 VCC.t9 sky130_fd_pr__pfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.54
X7 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.54
X8 VOUT.t6 VGP.t2 VIN.t5 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.16325 pd=7.38 as=2.7495 ps=14.88 w=7.05 l=2.54
X9 VOUT.t7 VGP.t3 VIN.t4 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.54
X10 VSS.t11 VSS.t8 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=2.98
X11 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=5.6082 pd=29.54 as=0 ps=0 w=14.38 l=2.98
R0 VGP.n26 VGP.n0 161.3
R1 VGP.n25 VGP.n24 161.3
R2 VGP.n23 VGP.n1 161.3
R3 VGP.n22 VGP.n21 161.3
R4 VGP.n20 VGP.n2 161.3
R5 VGP.n19 VGP.n18 161.3
R6 VGP.n17 VGP.n16 161.3
R7 VGP.n15 VGP.n4 161.3
R8 VGP.n14 VGP.n13 161.3
R9 VGP.n12 VGP.n5 161.3
R10 VGP.n11 VGP.n10 161.3
R11 VGP.n9 VGP.n6 161.3
R12 VGP.n28 VGP.n27 108.066
R13 VGP.n7 VGP.t2 98.0515
R14 VGP.n8 VGP.t0 66.8922
R15 VGP.n3 VGP.t3 66.8922
R16 VGP.n27 VGP.t1 66.8922
R17 VGP.n8 VGP.n7 63.437
R18 VGP.n14 VGP.n5 56.5193
R19 VGP.n21 VGP.n1 52.1486
R20 VGP.n21 VGP.n20 28.8382
R21 VGP.n10 VGP.n5 24.4675
R22 VGP.n10 VGP.n9 24.4675
R23 VGP.n20 VGP.n19 24.4675
R24 VGP.n16 VGP.n15 24.4675
R25 VGP.n15 VGP.n14 24.4675
R26 VGP.n26 VGP.n25 24.4675
R27 VGP.n25 VGP.n1 24.4675
R28 VGP.n19 VGP.n3 15.4147
R29 VGP.n9 VGP.n8 9.05329
R30 VGP.n16 VGP.n3 9.05329
R31 VGP.n7 VGP.n6 7.31035
R32 VGP.n27 VGP.n26 2.69187
R33 VGP.n28 VGP.n0 0.278367
R34 VGP.n24 VGP.n0 0.189894
R35 VGP.n24 VGP.n23 0.189894
R36 VGP.n23 VGP.n22 0.189894
R37 VGP.n22 VGP.n2 0.189894
R38 VGP.n18 VGP.n2 0.189894
R39 VGP.n18 VGP.n17 0.189894
R40 VGP.n17 VGP.n4 0.189894
R41 VGP.n13 VGP.n4 0.189894
R42 VGP.n13 VGP.n12 0.189894
R43 VGP.n12 VGP.n11 0.189894
R44 VGP.n11 VGP.n6 0.189894
R45 VGP VGP.n28 0.174287
R46 VOUT.n2 VOUT.n0 88.6584
R47 VOUT.n2 VOUT.n1 86.1831
R48 VOUT.n5 VOUT.n3 65.7587
R49 VOUT.n5 VOUT.n4 62.9053
R50 VOUT VOUT.n5 12.5652
R51 VOUT.n1 VOUT.t4 4.61114
R52 VOUT.n1 VOUT.t6 4.61114
R53 VOUT.n0 VOUT.t5 4.61114
R54 VOUT.n0 VOUT.t7 4.61114
R55 VOUT.n4 VOUT.t2 1.37741
R56 VOUT.n4 VOUT.t1 1.37741
R57 VOUT.n3 VOUT.t3 1.37741
R58 VOUT.n3 VOUT.t0 1.37741
R59 VOUT VOUT.n2 1.35826
R60 VIN.n1 VIN.t5 76.5903
R61 VIN.n2 VIN.t6 74.1159
R62 VIN.n1 VIN.n0 69.5055
R63 VIN.n4 VIN.t1 50.4568
R64 VIN.n5 VIN.t3 47.6033
R65 VIN.n4 VIN.n3 46.2265
R66 VIN VIN.n2 11.7462
R67 VIN.n0 VIN.t4 4.61114
R68 VIN.n0 VIN.t7 4.61114
R69 VIN.n5 VIN.n4 2.85395
R70 VIN.n2 VIN.n1 2.47464
R71 VIN.n3 VIN.t0 1.37741
R72 VIN.n3 VIN.t2 1.37741
R73 VIN VIN.n5 0.00481034
R74 VCC.n390 VCC.n28 395.123
R75 VCC.n339 VCC.n338 395.123
R76 VCC.n205 VCC.n135 395.123
R77 VCC.n207 VCC.n133 395.123
R78 VCC.n44 VCC.t8 274.846
R79 VCC.n148 VCC.t4 274.846
R80 VCC.n338 VCC.n337 185
R81 VCC.n338 VCC.n30 185
R82 VCC.n336 VCC.n48 185
R83 VCC.n328 VCC.n48 185
R84 VCC.n53 VCC.n49 185
R85 VCC.n329 VCC.n53 185
R86 VCC.n332 VCC.n331 185
R87 VCC.n331 VCC.n330 185
R88 VCC.n52 VCC.n51 185
R89 VCC.n327 VCC.n52 185
R90 VCC.n324 VCC.n323 185
R91 VCC.n325 VCC.n324 185
R92 VCC.n56 VCC.n55 185
R93 VCC.n55 VCC.n54 185
R94 VCC.n319 VCC.n318 185
R95 VCC.n318 VCC.n317 185
R96 VCC.n59 VCC.n58 185
R97 VCC.n316 VCC.n59 185
R98 VCC.n313 VCC.n312 185
R99 VCC.n314 VCC.n313 185
R100 VCC.n62 VCC.n61 185
R101 VCC.n61 VCC.n60 185
R102 VCC.n308 VCC.n307 185
R103 VCC.n307 VCC.n306 185
R104 VCC.n65 VCC.n64 185
R105 VCC.n305 VCC.n65 185
R106 VCC.n302 VCC.n301 185
R107 VCC.n303 VCC.n302 185
R108 VCC.n68 VCC.n67 185
R109 VCC.n67 VCC.n66 185
R110 VCC.n297 VCC.n296 185
R111 VCC.n296 VCC.n295 185
R112 VCC.n71 VCC.n70 185
R113 VCC.n294 VCC.n71 185
R114 VCC.n291 VCC.n290 185
R115 VCC.n292 VCC.n291 185
R116 VCC.n74 VCC.n73 185
R117 VCC.n73 VCC.n72 185
R118 VCC.n286 VCC.n285 185
R119 VCC.n285 VCC.n284 185
R120 VCC.n77 VCC.n76 185
R121 VCC.n283 VCC.n77 185
R122 VCC.n88 VCC.n86 185
R123 VCC.n86 VCC.n78 185
R124 VCC.n272 VCC.n271 185
R125 VCC.n273 VCC.n272 185
R126 VCC.n87 VCC.n85 185
R127 VCC.n274 VCC.n85 185
R128 VCC.n266 VCC.n265 185
R129 VCC.n265 VCC.n84 185
R130 VCC.n264 VCC.n90 185
R131 VCC.n264 VCC.n263 185
R132 VCC.n101 VCC.n91 185
R133 VCC.n92 VCC.n91 185
R134 VCC.n254 VCC.n253 185
R135 VCC.n255 VCC.n254 185
R136 VCC.n100 VCC.n99 185
R137 VCC.n99 VCC.n98 185
R138 VCC.n248 VCC.n247 185
R139 VCC.n247 VCC.n246 185
R140 VCC.n104 VCC.n103 185
R141 VCC.n105 VCC.n104 185
R142 VCC.n237 VCC.n236 185
R143 VCC.n238 VCC.n237 185
R144 VCC.n113 VCC.n112 185
R145 VCC.n112 VCC.n111 185
R146 VCC.n232 VCC.n231 185
R147 VCC.n231 VCC.n230 185
R148 VCC.n116 VCC.n115 185
R149 VCC.n117 VCC.n116 185
R150 VCC.n221 VCC.n220 185
R151 VCC.n222 VCC.n221 185
R152 VCC.n125 VCC.n124 185
R153 VCC.n124 VCC.n123 185
R154 VCC.n216 VCC.n215 185
R155 VCC.n215 VCC.n214 185
R156 VCC.n128 VCC.n127 185
R157 VCC.n129 VCC.n128 185
R158 VCC.n205 VCC.n204 185
R159 VCC.n206 VCC.n205 185
R160 VCC.n208 VCC.n207 185
R161 VCC.n207 VCC.n206 185
R162 VCC.n131 VCC.n130 185
R163 VCC.n130 VCC.n129 185
R164 VCC.n213 VCC.n212 185
R165 VCC.n214 VCC.n213 185
R166 VCC.n122 VCC.n121 185
R167 VCC.n123 VCC.n122 185
R168 VCC.n224 VCC.n223 185
R169 VCC.n223 VCC.n222 185
R170 VCC.n119 VCC.n118 185
R171 VCC.n118 VCC.n117 185
R172 VCC.n229 VCC.n228 185
R173 VCC.n230 VCC.n229 185
R174 VCC.n110 VCC.n109 185
R175 VCC.n111 VCC.n110 185
R176 VCC.n240 VCC.n239 185
R177 VCC.n239 VCC.n238 185
R178 VCC.n107 VCC.n106 185
R179 VCC.n106 VCC.n105 185
R180 VCC.n245 VCC.n244 185
R181 VCC.n246 VCC.n245 185
R182 VCC.n97 VCC.n96 185
R183 VCC.n98 VCC.n97 185
R184 VCC.n257 VCC.n256 185
R185 VCC.n256 VCC.n255 185
R186 VCC.n94 VCC.n93 185
R187 VCC.n93 VCC.n92 185
R188 VCC.n262 VCC.n261 185
R189 VCC.n263 VCC.n262 185
R190 VCC.n83 VCC.n82 185
R191 VCC.n84 VCC.n83 185
R192 VCC.n276 VCC.n275 185
R193 VCC.n275 VCC.n274 185
R194 VCC.n80 VCC.n79 185
R195 VCC.n273 VCC.n79 185
R196 VCC.n281 VCC.n280 185
R197 VCC.n281 VCC.n78 185
R198 VCC.n282 VCC.n2 185
R199 VCC.n283 VCC.n282 185
R200 VCC.n420 VCC.n3 185
R201 VCC.n284 VCC.n3 185
R202 VCC.n419 VCC.n4 185
R203 VCC.n72 VCC.n4 185
R204 VCC.n418 VCC.n5 185
R205 VCC.n292 VCC.n5 185
R206 VCC.n293 VCC.n6 185
R207 VCC.n294 VCC.n293 185
R208 VCC.n414 VCC.n8 185
R209 VCC.n295 VCC.n8 185
R210 VCC.n413 VCC.n9 185
R211 VCC.n66 VCC.n9 185
R212 VCC.n412 VCC.n10 185
R213 VCC.n303 VCC.n10 185
R214 VCC.n304 VCC.n11 185
R215 VCC.n305 VCC.n304 185
R216 VCC.n408 VCC.n13 185
R217 VCC.n306 VCC.n13 185
R218 VCC.n407 VCC.n14 185
R219 VCC.n60 VCC.n14 185
R220 VCC.n406 VCC.n15 185
R221 VCC.n314 VCC.n15 185
R222 VCC.n315 VCC.n16 185
R223 VCC.n316 VCC.n315 185
R224 VCC.n402 VCC.n18 185
R225 VCC.n317 VCC.n18 185
R226 VCC.n401 VCC.n19 185
R227 VCC.n54 VCC.n19 185
R228 VCC.n400 VCC.n20 185
R229 VCC.n325 VCC.n20 185
R230 VCC.n326 VCC.n21 185
R231 VCC.n327 VCC.n326 185
R232 VCC.n396 VCC.n23 185
R233 VCC.n330 VCC.n23 185
R234 VCC.n395 VCC.n24 185
R235 VCC.n329 VCC.n24 185
R236 VCC.n394 VCC.n25 185
R237 VCC.n328 VCC.n25 185
R238 VCC.n28 VCC.n26 185
R239 VCC.n30 VCC.n28 185
R240 VCC.n340 VCC.n339 185
R241 VCC.n342 VCC.n341 185
R242 VCC.n344 VCC.n343 185
R243 VCC.n346 VCC.n345 185
R244 VCC.n348 VCC.n347 185
R245 VCC.n350 VCC.n349 185
R246 VCC.n352 VCC.n351 185
R247 VCC.n354 VCC.n353 185
R248 VCC.n356 VCC.n355 185
R249 VCC.n358 VCC.n357 185
R250 VCC.n360 VCC.n359 185
R251 VCC.n362 VCC.n361 185
R252 VCC.n364 VCC.n363 185
R253 VCC.n366 VCC.n365 185
R254 VCC.n368 VCC.n367 185
R255 VCC.n370 VCC.n369 185
R256 VCC.n372 VCC.n371 185
R257 VCC.n374 VCC.n373 185
R258 VCC.n376 VCC.n375 185
R259 VCC.n378 VCC.n377 185
R260 VCC.n380 VCC.n379 185
R261 VCC.n382 VCC.n381 185
R262 VCC.n384 VCC.n383 185
R263 VCC.n385 VCC.n43 185
R264 VCC.n387 VCC.n386 185
R265 VCC.n29 VCC.n27 185
R266 VCC.n391 VCC.n390 185
R267 VCC.n390 VCC.n389 185
R268 VCC.n133 VCC.n132 185
R269 VCC.n152 VCC.n151 185
R270 VCC.n154 VCC.n147 185
R271 VCC.n147 VCC.n134 185
R272 VCC.n156 VCC.n155 185
R273 VCC.n158 VCC.n146 185
R274 VCC.n161 VCC.n160 185
R275 VCC.n162 VCC.n145 185
R276 VCC.n164 VCC.n163 185
R277 VCC.n166 VCC.n144 185
R278 VCC.n169 VCC.n168 185
R279 VCC.n170 VCC.n143 185
R280 VCC.n172 VCC.n171 185
R281 VCC.n174 VCC.n142 185
R282 VCC.n177 VCC.n176 185
R283 VCC.n178 VCC.n141 185
R284 VCC.n180 VCC.n179 185
R285 VCC.n182 VCC.n140 185
R286 VCC.n185 VCC.n184 185
R287 VCC.n186 VCC.n139 185
R288 VCC.n188 VCC.n187 185
R289 VCC.n190 VCC.n138 185
R290 VCC.n193 VCC.n192 185
R291 VCC.n194 VCC.n137 185
R292 VCC.n196 VCC.n195 185
R293 VCC.n198 VCC.n136 185
R294 VCC.n201 VCC.n200 185
R295 VCC.n202 VCC.n135 185
R296 VCC.n44 VCC.t10 170.094
R297 VCC.n148 VCC.t7 170.094
R298 VCC.n205 VCC.n128 146.341
R299 VCC.n215 VCC.n128 146.341
R300 VCC.n215 VCC.n124 146.341
R301 VCC.n221 VCC.n124 146.341
R302 VCC.n221 VCC.n116 146.341
R303 VCC.n231 VCC.n116 146.341
R304 VCC.n231 VCC.n112 146.341
R305 VCC.n237 VCC.n112 146.341
R306 VCC.n237 VCC.n104 146.341
R307 VCC.n247 VCC.n104 146.341
R308 VCC.n247 VCC.n99 146.341
R309 VCC.n254 VCC.n99 146.341
R310 VCC.n254 VCC.n91 146.341
R311 VCC.n264 VCC.n91 146.341
R312 VCC.n265 VCC.n264 146.341
R313 VCC.n265 VCC.n85 146.341
R314 VCC.n272 VCC.n85 146.341
R315 VCC.n272 VCC.n86 146.341
R316 VCC.n86 VCC.n77 146.341
R317 VCC.n285 VCC.n77 146.341
R318 VCC.n285 VCC.n73 146.341
R319 VCC.n291 VCC.n73 146.341
R320 VCC.n291 VCC.n71 146.341
R321 VCC.n296 VCC.n71 146.341
R322 VCC.n296 VCC.n67 146.341
R323 VCC.n302 VCC.n67 146.341
R324 VCC.n302 VCC.n65 146.341
R325 VCC.n307 VCC.n65 146.341
R326 VCC.n307 VCC.n61 146.341
R327 VCC.n313 VCC.n61 146.341
R328 VCC.n313 VCC.n59 146.341
R329 VCC.n318 VCC.n59 146.341
R330 VCC.n318 VCC.n55 146.341
R331 VCC.n324 VCC.n55 146.341
R332 VCC.n324 VCC.n52 146.341
R333 VCC.n331 VCC.n52 146.341
R334 VCC.n331 VCC.n53 146.341
R335 VCC.n53 VCC.n48 146.341
R336 VCC.n338 VCC.n48 146.341
R337 VCC.n207 VCC.n130 146.341
R338 VCC.n213 VCC.n130 146.341
R339 VCC.n213 VCC.n122 146.341
R340 VCC.n223 VCC.n122 146.341
R341 VCC.n223 VCC.n118 146.341
R342 VCC.n229 VCC.n118 146.341
R343 VCC.n229 VCC.n110 146.341
R344 VCC.n239 VCC.n110 146.341
R345 VCC.n239 VCC.n106 146.341
R346 VCC.n245 VCC.n106 146.341
R347 VCC.n245 VCC.n97 146.341
R348 VCC.n256 VCC.n97 146.341
R349 VCC.n256 VCC.n93 146.341
R350 VCC.n262 VCC.n93 146.341
R351 VCC.n262 VCC.n83 146.341
R352 VCC.n275 VCC.n83 146.341
R353 VCC.n275 VCC.n79 146.341
R354 VCC.n281 VCC.n79 146.341
R355 VCC.n282 VCC.n281 146.341
R356 VCC.n282 VCC.n3 146.341
R357 VCC.n4 VCC.n3 146.341
R358 VCC.n5 VCC.n4 146.341
R359 VCC.n293 VCC.n5 146.341
R360 VCC.n293 VCC.n8 146.341
R361 VCC.n9 VCC.n8 146.341
R362 VCC.n10 VCC.n9 146.341
R363 VCC.n304 VCC.n10 146.341
R364 VCC.n304 VCC.n13 146.341
R365 VCC.n14 VCC.n13 146.341
R366 VCC.n15 VCC.n14 146.341
R367 VCC.n315 VCC.n15 146.341
R368 VCC.n315 VCC.n18 146.341
R369 VCC.n19 VCC.n18 146.341
R370 VCC.n20 VCC.n19 146.341
R371 VCC.n326 VCC.n20 146.341
R372 VCC.n326 VCC.n23 146.341
R373 VCC.n24 VCC.n23 146.341
R374 VCC.n25 VCC.n24 146.341
R375 VCC.n28 VCC.n25 146.341
R376 VCC.n45 VCC.t11 114.433
R377 VCC.n149 VCC.t6 114.433
R378 VCC.n390 VCC.n29 99.5127
R379 VCC.n387 VCC.n43 99.5127
R380 VCC.n383 VCC.n382 99.5127
R381 VCC.n379 VCC.n378 99.5127
R382 VCC.n375 VCC.n374 99.5127
R383 VCC.n371 VCC.n370 99.5127
R384 VCC.n367 VCC.n366 99.5127
R385 VCC.n363 VCC.n362 99.5127
R386 VCC.n359 VCC.n358 99.5127
R387 VCC.n355 VCC.n354 99.5127
R388 VCC.n351 VCC.n350 99.5127
R389 VCC.n347 VCC.n346 99.5127
R390 VCC.n343 VCC.n342 99.5127
R391 VCC.n151 VCC.n147 99.5127
R392 VCC.n156 VCC.n147 99.5127
R393 VCC.n160 VCC.n158 99.5127
R394 VCC.n164 VCC.n145 99.5127
R395 VCC.n168 VCC.n166 99.5127
R396 VCC.n172 VCC.n143 99.5127
R397 VCC.n176 VCC.n174 99.5127
R398 VCC.n180 VCC.n141 99.5127
R399 VCC.n184 VCC.n182 99.5127
R400 VCC.n188 VCC.n139 99.5127
R401 VCC.n192 VCC.n190 99.5127
R402 VCC.n196 VCC.n137 99.5127
R403 VCC.n200 VCC.n198 99.5127
R404 VCC.n206 VCC.n134 77.4647
R405 VCC.n389 VCC.n30 77.4647
R406 VCC.n389 VCC.n31 72.8958
R407 VCC.n389 VCC.n32 72.8958
R408 VCC.n389 VCC.n33 72.8958
R409 VCC.n389 VCC.n34 72.8958
R410 VCC.n389 VCC.n35 72.8958
R411 VCC.n389 VCC.n36 72.8958
R412 VCC.n389 VCC.n37 72.8958
R413 VCC.n389 VCC.n38 72.8958
R414 VCC.n389 VCC.n39 72.8958
R415 VCC.n389 VCC.n40 72.8958
R416 VCC.n389 VCC.n41 72.8958
R417 VCC.n389 VCC.n42 72.8958
R418 VCC.n389 VCC.n388 72.8958
R419 VCC.n150 VCC.n134 72.8958
R420 VCC.n157 VCC.n134 72.8958
R421 VCC.n159 VCC.n134 72.8958
R422 VCC.n165 VCC.n134 72.8958
R423 VCC.n167 VCC.n134 72.8958
R424 VCC.n173 VCC.n134 72.8958
R425 VCC.n175 VCC.n134 72.8958
R426 VCC.n181 VCC.n134 72.8958
R427 VCC.n183 VCC.n134 72.8958
R428 VCC.n189 VCC.n134 72.8958
R429 VCC.n191 VCC.n134 72.8958
R430 VCC.n197 VCC.n134 72.8958
R431 VCC.n199 VCC.n134 72.8958
R432 VCC.n45 VCC.n44 55.6611
R433 VCC.n149 VCC.n148 55.6611
R434 VCC.n206 VCC.n129 42.5632
R435 VCC.n214 VCC.n129 42.5632
R436 VCC.n222 VCC.n123 42.5632
R437 VCC.n222 VCC.n117 42.5632
R438 VCC.n230 VCC.n117 42.5632
R439 VCC.n230 VCC.n111 42.5632
R440 VCC.n238 VCC.n111 42.5632
R441 VCC.n238 VCC.n105 42.5632
R442 VCC.n246 VCC.n105 42.5632
R443 VCC.n255 VCC.n98 42.5632
R444 VCC.n255 VCC.n92 42.5632
R445 VCC.n263 VCC.n92 42.5632
R446 VCC.n263 VCC.n84 42.5632
R447 VCC.n274 VCC.n84 42.5632
R448 VCC.n273 VCC.n78 42.5632
R449 VCC.n283 VCC.n78 42.5632
R450 VCC.n284 VCC.n283 42.5632
R451 VCC.n284 VCC.n72 42.5632
R452 VCC.n292 VCC.n72 42.5632
R453 VCC.n295 VCC.n294 42.5632
R454 VCC.n295 VCC.n66 42.5632
R455 VCC.n303 VCC.n66 42.5632
R456 VCC.n305 VCC.n303 42.5632
R457 VCC.n306 VCC.n305 42.5632
R458 VCC.n314 VCC.n60 42.5632
R459 VCC.n316 VCC.n314 42.5632
R460 VCC.n317 VCC.n316 42.5632
R461 VCC.n317 VCC.n54 42.5632
R462 VCC.n325 VCC.n54 42.5632
R463 VCC.n327 VCC.n325 42.5632
R464 VCC.n330 VCC.n327 42.5632
R465 VCC.n329 VCC.n328 42.5632
R466 VCC.n328 VCC.n30 42.5632
R467 VCC.n214 VCC.t5 41.2863
R468 VCC.t9 VCC.n329 41.2863
R469 VCC.n388 VCC.n387 39.2114
R470 VCC.n383 VCC.n42 39.2114
R471 VCC.n379 VCC.n41 39.2114
R472 VCC.n375 VCC.n40 39.2114
R473 VCC.n371 VCC.n39 39.2114
R474 VCC.n367 VCC.n38 39.2114
R475 VCC.n363 VCC.n37 39.2114
R476 VCC.n359 VCC.n36 39.2114
R477 VCC.n355 VCC.n35 39.2114
R478 VCC.n351 VCC.n34 39.2114
R479 VCC.n347 VCC.n33 39.2114
R480 VCC.n343 VCC.n32 39.2114
R481 VCC.n339 VCC.n31 39.2114
R482 VCC.n150 VCC.n133 39.2114
R483 VCC.n157 VCC.n156 39.2114
R484 VCC.n160 VCC.n159 39.2114
R485 VCC.n165 VCC.n164 39.2114
R486 VCC.n168 VCC.n167 39.2114
R487 VCC.n173 VCC.n172 39.2114
R488 VCC.n176 VCC.n175 39.2114
R489 VCC.n181 VCC.n180 39.2114
R490 VCC.n184 VCC.n183 39.2114
R491 VCC.n189 VCC.n188 39.2114
R492 VCC.n192 VCC.n191 39.2114
R493 VCC.n197 VCC.n196 39.2114
R494 VCC.n200 VCC.n199 39.2114
R495 VCC.n342 VCC.n31 39.2114
R496 VCC.n346 VCC.n32 39.2114
R497 VCC.n350 VCC.n33 39.2114
R498 VCC.n354 VCC.n34 39.2114
R499 VCC.n358 VCC.n35 39.2114
R500 VCC.n362 VCC.n36 39.2114
R501 VCC.n366 VCC.n37 39.2114
R502 VCC.n370 VCC.n38 39.2114
R503 VCC.n374 VCC.n39 39.2114
R504 VCC.n378 VCC.n40 39.2114
R505 VCC.n382 VCC.n41 39.2114
R506 VCC.n43 VCC.n42 39.2114
R507 VCC.n388 VCC.n29 39.2114
R508 VCC.n151 VCC.n150 39.2114
R509 VCC.n158 VCC.n157 39.2114
R510 VCC.n159 VCC.n145 39.2114
R511 VCC.n166 VCC.n165 39.2114
R512 VCC.n167 VCC.n143 39.2114
R513 VCC.n174 VCC.n173 39.2114
R514 VCC.n175 VCC.n141 39.2114
R515 VCC.n182 VCC.n181 39.2114
R516 VCC.n183 VCC.n139 39.2114
R517 VCC.n190 VCC.n189 39.2114
R518 VCC.n191 VCC.n137 39.2114
R519 VCC.n198 VCC.n197 39.2114
R520 VCC.n199 VCC.n135 39.2114
R521 VCC.n246 VCC.t2 37.8813
R522 VCC.t1 VCC.n60 37.8813
R523 VCC.n392 VCC.n391 29.7145
R524 VCC.n340 VCC.n47 29.7145
R525 VCC.n209 VCC.n132 29.7145
R526 VCC.n203 VCC.n202 29.7145
R527 VCC.n46 VCC.n45 29.2853
R528 VCC.n153 VCC.n149 29.2853
R529 VCC.n274 VCC.t0 26.815
R530 VCC.n294 VCC.t3 26.815
R531 VCC.n204 VCC.n127 19.3944
R532 VCC.n216 VCC.n127 19.3944
R533 VCC.n216 VCC.n125 19.3944
R534 VCC.n220 VCC.n125 19.3944
R535 VCC.n220 VCC.n115 19.3944
R536 VCC.n232 VCC.n115 19.3944
R537 VCC.n232 VCC.n113 19.3944
R538 VCC.n236 VCC.n113 19.3944
R539 VCC.n236 VCC.n103 19.3944
R540 VCC.n248 VCC.n103 19.3944
R541 VCC.n248 VCC.n100 19.3944
R542 VCC.n253 VCC.n100 19.3944
R543 VCC.n253 VCC.n101 19.3944
R544 VCC.n101 VCC.n90 19.3944
R545 VCC.n266 VCC.n90 19.3944
R546 VCC.n266 VCC.n87 19.3944
R547 VCC.n271 VCC.n87 19.3944
R548 VCC.n271 VCC.n88 19.3944
R549 VCC.n88 VCC.n76 19.3944
R550 VCC.n286 VCC.n76 19.3944
R551 VCC.n286 VCC.n74 19.3944
R552 VCC.n290 VCC.n74 19.3944
R553 VCC.n290 VCC.n70 19.3944
R554 VCC.n297 VCC.n70 19.3944
R555 VCC.n297 VCC.n68 19.3944
R556 VCC.n301 VCC.n68 19.3944
R557 VCC.n301 VCC.n64 19.3944
R558 VCC.n308 VCC.n64 19.3944
R559 VCC.n308 VCC.n62 19.3944
R560 VCC.n312 VCC.n62 19.3944
R561 VCC.n312 VCC.n58 19.3944
R562 VCC.n319 VCC.n58 19.3944
R563 VCC.n319 VCC.n56 19.3944
R564 VCC.n323 VCC.n56 19.3944
R565 VCC.n323 VCC.n51 19.3944
R566 VCC.n332 VCC.n51 19.3944
R567 VCC.n332 VCC.n49 19.3944
R568 VCC.n336 VCC.n49 19.3944
R569 VCC.n337 VCC.n336 19.3944
R570 VCC.n208 VCC.n131 19.3944
R571 VCC.n212 VCC.n131 19.3944
R572 VCC.n212 VCC.n121 19.3944
R573 VCC.n224 VCC.n121 19.3944
R574 VCC.n224 VCC.n119 19.3944
R575 VCC.n228 VCC.n119 19.3944
R576 VCC.n228 VCC.n109 19.3944
R577 VCC.n240 VCC.n109 19.3944
R578 VCC.n240 VCC.n107 19.3944
R579 VCC.n244 VCC.n107 19.3944
R580 VCC.n244 VCC.n96 19.3944
R581 VCC.n257 VCC.n96 19.3944
R582 VCC.n257 VCC.n94 19.3944
R583 VCC.n261 VCC.n94 19.3944
R584 VCC.n261 VCC.n82 19.3944
R585 VCC.n276 VCC.n82 19.3944
R586 VCC.n276 VCC.n80 19.3944
R587 VCC.n280 VCC.n80 19.3944
R588 VCC.n280 VCC.n2 19.3944
R589 VCC.n420 VCC.n2 19.3944
R590 VCC.n420 VCC.n419 19.3944
R591 VCC.n419 VCC.n418 19.3944
R592 VCC.n418 VCC.n6 19.3944
R593 VCC.n414 VCC.n6 19.3944
R594 VCC.n414 VCC.n413 19.3944
R595 VCC.n413 VCC.n412 19.3944
R596 VCC.n412 VCC.n11 19.3944
R597 VCC.n408 VCC.n11 19.3944
R598 VCC.n408 VCC.n407 19.3944
R599 VCC.n407 VCC.n406 19.3944
R600 VCC.n406 VCC.n16 19.3944
R601 VCC.n402 VCC.n16 19.3944
R602 VCC.n402 VCC.n401 19.3944
R603 VCC.n401 VCC.n400 19.3944
R604 VCC.n400 VCC.n21 19.3944
R605 VCC.n396 VCC.n21 19.3944
R606 VCC.n396 VCC.n395 19.3944
R607 VCC.n395 VCC.n394 19.3944
R608 VCC.n394 VCC.n26 19.3944
R609 VCC.t0 VCC.n273 15.7487
R610 VCC.t3 VCC.n292 15.7487
R611 VCC.n391 VCC.n27 10.6151
R612 VCC.n386 VCC.n385 10.6151
R613 VCC.n385 VCC.n384 10.6151
R614 VCC.n384 VCC.n381 10.6151
R615 VCC.n381 VCC.n380 10.6151
R616 VCC.n380 VCC.n377 10.6151
R617 VCC.n377 VCC.n376 10.6151
R618 VCC.n376 VCC.n373 10.6151
R619 VCC.n373 VCC.n372 10.6151
R620 VCC.n372 VCC.n369 10.6151
R621 VCC.n369 VCC.n368 10.6151
R622 VCC.n368 VCC.n365 10.6151
R623 VCC.n365 VCC.n364 10.6151
R624 VCC.n364 VCC.n361 10.6151
R625 VCC.n361 VCC.n360 10.6151
R626 VCC.n360 VCC.n357 10.6151
R627 VCC.n357 VCC.n356 10.6151
R628 VCC.n356 VCC.n353 10.6151
R629 VCC.n353 VCC.n352 10.6151
R630 VCC.n352 VCC.n349 10.6151
R631 VCC.n349 VCC.n348 10.6151
R632 VCC.n348 VCC.n345 10.6151
R633 VCC.n345 VCC.n344 10.6151
R634 VCC.n344 VCC.n341 10.6151
R635 VCC.n341 VCC.n340 10.6151
R636 VCC.n152 VCC.n132 10.6151
R637 VCC.n155 VCC.n154 10.6151
R638 VCC.n155 VCC.n146 10.6151
R639 VCC.n161 VCC.n146 10.6151
R640 VCC.n162 VCC.n161 10.6151
R641 VCC.n163 VCC.n162 10.6151
R642 VCC.n163 VCC.n144 10.6151
R643 VCC.n169 VCC.n144 10.6151
R644 VCC.n170 VCC.n169 10.6151
R645 VCC.n171 VCC.n170 10.6151
R646 VCC.n171 VCC.n142 10.6151
R647 VCC.n177 VCC.n142 10.6151
R648 VCC.n178 VCC.n177 10.6151
R649 VCC.n179 VCC.n178 10.6151
R650 VCC.n179 VCC.n140 10.6151
R651 VCC.n185 VCC.n140 10.6151
R652 VCC.n186 VCC.n185 10.6151
R653 VCC.n187 VCC.n186 10.6151
R654 VCC.n187 VCC.n138 10.6151
R655 VCC.n193 VCC.n138 10.6151
R656 VCC.n194 VCC.n193 10.6151
R657 VCC.n195 VCC.n194 10.6151
R658 VCC.n195 VCC.n136 10.6151
R659 VCC.n201 VCC.n136 10.6151
R660 VCC.n202 VCC.n201 10.6151
R661 VCC.n419 VCC.n0 9.3005
R662 VCC.n418 VCC.n417 9.3005
R663 VCC.n416 VCC.n6 9.3005
R664 VCC.n415 VCC.n414 9.3005
R665 VCC.n413 VCC.n7 9.3005
R666 VCC.n412 VCC.n411 9.3005
R667 VCC.n410 VCC.n11 9.3005
R668 VCC.n409 VCC.n408 9.3005
R669 VCC.n407 VCC.n12 9.3005
R670 VCC.n406 VCC.n405 9.3005
R671 VCC.n404 VCC.n16 9.3005
R672 VCC.n403 VCC.n402 9.3005
R673 VCC.n401 VCC.n17 9.3005
R674 VCC.n400 VCC.n399 9.3005
R675 VCC.n398 VCC.n21 9.3005
R676 VCC.n397 VCC.n396 9.3005
R677 VCC.n395 VCC.n22 9.3005
R678 VCC.n394 VCC.n393 9.3005
R679 VCC.n392 VCC.n26 9.3005
R680 VCC.n127 VCC.n126 9.3005
R681 VCC.n217 VCC.n216 9.3005
R682 VCC.n218 VCC.n125 9.3005
R683 VCC.n220 VCC.n219 9.3005
R684 VCC.n115 VCC.n114 9.3005
R685 VCC.n233 VCC.n232 9.3005
R686 VCC.n234 VCC.n113 9.3005
R687 VCC.n236 VCC.n235 9.3005
R688 VCC.n103 VCC.n102 9.3005
R689 VCC.n249 VCC.n248 9.3005
R690 VCC.n250 VCC.n100 9.3005
R691 VCC.n253 VCC.n252 9.3005
R692 VCC.n251 VCC.n101 9.3005
R693 VCC.n90 VCC.n89 9.3005
R694 VCC.n267 VCC.n266 9.3005
R695 VCC.n268 VCC.n87 9.3005
R696 VCC.n271 VCC.n270 9.3005
R697 VCC.n269 VCC.n88 9.3005
R698 VCC.n76 VCC.n75 9.3005
R699 VCC.n287 VCC.n286 9.3005
R700 VCC.n288 VCC.n74 9.3005
R701 VCC.n290 VCC.n289 9.3005
R702 VCC.n70 VCC.n69 9.3005
R703 VCC.n298 VCC.n297 9.3005
R704 VCC.n299 VCC.n68 9.3005
R705 VCC.n301 VCC.n300 9.3005
R706 VCC.n64 VCC.n63 9.3005
R707 VCC.n309 VCC.n308 9.3005
R708 VCC.n310 VCC.n62 9.3005
R709 VCC.n312 VCC.n311 9.3005
R710 VCC.n58 VCC.n57 9.3005
R711 VCC.n320 VCC.n319 9.3005
R712 VCC.n321 VCC.n56 9.3005
R713 VCC.n323 VCC.n322 9.3005
R714 VCC.n51 VCC.n50 9.3005
R715 VCC.n333 VCC.n332 9.3005
R716 VCC.n334 VCC.n49 9.3005
R717 VCC.n336 VCC.n335 9.3005
R718 VCC.n337 VCC.n47 9.3005
R719 VCC.n204 VCC.n203 9.3005
R720 VCC.n209 VCC.n208 9.3005
R721 VCC.n210 VCC.n131 9.3005
R722 VCC.n212 VCC.n211 9.3005
R723 VCC.n121 VCC.n120 9.3005
R724 VCC.n225 VCC.n224 9.3005
R725 VCC.n226 VCC.n119 9.3005
R726 VCC.n228 VCC.n227 9.3005
R727 VCC.n109 VCC.n108 9.3005
R728 VCC.n241 VCC.n240 9.3005
R729 VCC.n242 VCC.n107 9.3005
R730 VCC.n244 VCC.n243 9.3005
R731 VCC.n96 VCC.n95 9.3005
R732 VCC.n258 VCC.n257 9.3005
R733 VCC.n259 VCC.n94 9.3005
R734 VCC.n261 VCC.n260 9.3005
R735 VCC.n82 VCC.n81 9.3005
R736 VCC.n277 VCC.n276 9.3005
R737 VCC.n278 VCC.n80 9.3005
R738 VCC.n280 VCC.n279 9.3005
R739 VCC.n2 VCC.n1 9.3005
R740 VCC VCC.n420 9.3005
R741 VCC.n46 VCC.n27 6.5566
R742 VCC.n153 VCC.n152 6.5566
R743 VCC.t2 VCC.n98 4.6824
R744 VCC.n306 VCC.t1 4.6824
R745 VCC.n386 VCC.n46 4.05904
R746 VCC.n154 VCC.n153 4.05904
R747 VCC.t5 VCC.n123 1.27738
R748 VCC.n330 VCC.t9 1.27738
R749 VCC VCC.n0 0.152939
R750 VCC.n417 VCC.n0 0.152939
R751 VCC.n417 VCC.n416 0.152939
R752 VCC.n416 VCC.n415 0.152939
R753 VCC.n415 VCC.n7 0.152939
R754 VCC.n411 VCC.n7 0.152939
R755 VCC.n411 VCC.n410 0.152939
R756 VCC.n410 VCC.n409 0.152939
R757 VCC.n409 VCC.n12 0.152939
R758 VCC.n405 VCC.n12 0.152939
R759 VCC.n405 VCC.n404 0.152939
R760 VCC.n404 VCC.n403 0.152939
R761 VCC.n403 VCC.n17 0.152939
R762 VCC.n399 VCC.n17 0.152939
R763 VCC.n399 VCC.n398 0.152939
R764 VCC.n398 VCC.n397 0.152939
R765 VCC.n397 VCC.n22 0.152939
R766 VCC.n393 VCC.n22 0.152939
R767 VCC.n393 VCC.n392 0.152939
R768 VCC.n203 VCC.n126 0.152939
R769 VCC.n217 VCC.n126 0.152939
R770 VCC.n218 VCC.n217 0.152939
R771 VCC.n219 VCC.n218 0.152939
R772 VCC.n219 VCC.n114 0.152939
R773 VCC.n233 VCC.n114 0.152939
R774 VCC.n234 VCC.n233 0.152939
R775 VCC.n235 VCC.n234 0.152939
R776 VCC.n235 VCC.n102 0.152939
R777 VCC.n249 VCC.n102 0.152939
R778 VCC.n250 VCC.n249 0.152939
R779 VCC.n252 VCC.n250 0.152939
R780 VCC.n252 VCC.n251 0.152939
R781 VCC.n251 VCC.n89 0.152939
R782 VCC.n267 VCC.n89 0.152939
R783 VCC.n268 VCC.n267 0.152939
R784 VCC.n270 VCC.n268 0.152939
R785 VCC.n270 VCC.n269 0.152939
R786 VCC.n269 VCC.n75 0.152939
R787 VCC.n287 VCC.n75 0.152939
R788 VCC.n288 VCC.n287 0.152939
R789 VCC.n289 VCC.n288 0.152939
R790 VCC.n289 VCC.n69 0.152939
R791 VCC.n298 VCC.n69 0.152939
R792 VCC.n299 VCC.n298 0.152939
R793 VCC.n300 VCC.n299 0.152939
R794 VCC.n300 VCC.n63 0.152939
R795 VCC.n309 VCC.n63 0.152939
R796 VCC.n310 VCC.n309 0.152939
R797 VCC.n311 VCC.n310 0.152939
R798 VCC.n311 VCC.n57 0.152939
R799 VCC.n320 VCC.n57 0.152939
R800 VCC.n321 VCC.n320 0.152939
R801 VCC.n322 VCC.n321 0.152939
R802 VCC.n322 VCC.n50 0.152939
R803 VCC.n333 VCC.n50 0.152939
R804 VCC.n334 VCC.n333 0.152939
R805 VCC.n335 VCC.n334 0.152939
R806 VCC.n335 VCC.n47 0.152939
R807 VCC.n210 VCC.n209 0.152939
R808 VCC.n211 VCC.n210 0.152939
R809 VCC.n211 VCC.n120 0.152939
R810 VCC.n225 VCC.n120 0.152939
R811 VCC.n226 VCC.n225 0.152939
R812 VCC.n227 VCC.n226 0.152939
R813 VCC.n227 VCC.n108 0.152939
R814 VCC.n241 VCC.n108 0.152939
R815 VCC.n242 VCC.n241 0.152939
R816 VCC.n243 VCC.n242 0.152939
R817 VCC.n243 VCC.n95 0.152939
R818 VCC.n258 VCC.n95 0.152939
R819 VCC.n259 VCC.n258 0.152939
R820 VCC.n260 VCC.n259 0.152939
R821 VCC.n260 VCC.n81 0.152939
R822 VCC.n277 VCC.n81 0.152939
R823 VCC.n278 VCC.n277 0.152939
R824 VCC.n279 VCC.n278 0.152939
R825 VCC.n279 VCC.n1 0.152939
R826 VCC VCC.n1 0.1255
R827 VGN.n29 VGN.n28 161.3
R828 VGN.n27 VGN.n1 161.3
R829 VGN.n26 VGN.n25 161.3
R830 VGN.n24 VGN.n2 161.3
R831 VGN.n23 VGN.n22 161.3
R832 VGN.n21 VGN.n3 161.3
R833 VGN.n19 VGN.n18 161.3
R834 VGN.n17 VGN.n4 161.3
R835 VGN.n16 VGN.n15 161.3
R836 VGN.n14 VGN.n5 161.3
R837 VGN.n13 VGN.n12 161.3
R838 VGN.n11 VGN.n6 161.3
R839 VGN.n10 VGN.n9 161.3
R840 VGN.n7 VGN.t1 147.981
R841 VGN.n8 VGN.t0 116.296
R842 VGN.n20 VGN.t2 116.296
R843 VGN.n0 VGN.t3 116.296
R844 VGN.n30 VGN.n0 67.2516
R845 VGN.n8 VGN.n7 66.0814
R846 VGN.n26 VGN.n2 56.4773
R847 VGN.n14 VGN.n13 40.4106
R848 VGN.n15 VGN.n14 40.4106
R849 VGN.n13 VGN.n6 24.3439
R850 VGN.n9 VGN.n6 24.3439
R851 VGN.n22 VGN.n2 24.3439
R852 VGN.n22 VGN.n21 24.3439
R853 VGN.n19 VGN.n4 24.3439
R854 VGN.n15 VGN.n4 24.3439
R855 VGN.n28 VGN.n27 24.3439
R856 VGN.n27 VGN.n26 24.3439
R857 VGN.n28 VGN.n0 22.6399
R858 VGN.n21 VGN.n20 16.7975
R859 VGN.n9 VGN.n8 7.54696
R860 VGN.n20 VGN.n19 7.54696
R861 VGN.n10 VGN.n7 5.37324
R862 VGN.n30 VGN.n29 0.355081
R863 VGN VGN.n30 0.336926
R864 VGN.n29 VGN.n1 0.189894
R865 VGN.n25 VGN.n1 0.189894
R866 VGN.n25 VGN.n24 0.189894
R867 VGN.n24 VGN.n23 0.189894
R868 VGN.n23 VGN.n3 0.189894
R869 VGN.n18 VGN.n3 0.189894
R870 VGN.n18 VGN.n17 0.189894
R871 VGN.n17 VGN.n16 0.189894
R872 VGN.n16 VGN.n5 0.189894
R873 VGN.n12 VGN.n5 0.189894
R874 VGN.n12 VGN.n11 0.189894
R875 VGN.n11 VGN.n10 0.189894
R876 VSS.n291 VSS.n162 651.062
R877 VSS.n289 VSS.n164 651.062
R878 VSS.n534 VSS.n57 651.062
R879 VSS.n537 VSS.n30 651.062
R880 VSS.n292 VSS.n291 585
R881 VSS.n291 VSS.n290 585
R882 VSS.n160 VSS.n159 585
R883 VSS.n159 VSS.n157 585
R884 VSS.n297 VSS.n296 585
R885 VSS.n298 VSS.n297 585
R886 VSS.n151 VSS.n150 585
R887 VSS.n158 VSS.n151 585
R888 VSS.n308 VSS.n307 585
R889 VSS.n307 VSS.n306 585
R890 VSS.n148 VSS.n147 585
R891 VSS.n147 VSS.n146 585
R892 VSS.n313 VSS.n312 585
R893 VSS.n314 VSS.n313 585
R894 VSS.n139 VSS.n138 585
R895 VSS.n140 VSS.n139 585
R896 VSS.n324 VSS.n323 585
R897 VSS.n323 VSS.n322 585
R898 VSS.n136 VSS.n135 585
R899 VSS.n135 VSS.n134 585
R900 VSS.n329 VSS.n328 585
R901 VSS.n330 VSS.n329 585
R902 VSS.n127 VSS.n126 585
R903 VSS.n128 VSS.n127 585
R904 VSS.n340 VSS.n339 585
R905 VSS.n339 VSS.n338 585
R906 VSS.n124 VSS.n123 585
R907 VSS.n123 VSS.n122 585
R908 VSS.n345 VSS.n344 585
R909 VSS.n346 VSS.n345 585
R910 VSS.n115 VSS.n114 585
R911 VSS.n116 VSS.n115 585
R912 VSS.n356 VSS.n355 585
R913 VSS.n355 VSS.n354 585
R914 VSS.n112 VSS.n111 585
R915 VSS.n111 VSS.n109 585
R916 VSS.n361 VSS.n360 585
R917 VSS.n362 VSS.n361 585
R918 VSS.n101 VSS.n100 585
R919 VSS.n110 VSS.n101 585
R920 VSS.n373 VSS.n372 585
R921 VSS.n372 VSS.n371 585
R922 VSS.n98 VSS.n97 585
R923 VSS.n97 VSS.n95 585
R924 VSS.n378 VSS.n377 585
R925 VSS.n379 VSS.n378 585
R926 VSS.n94 VSS.n93 585
R927 VSS.n380 VSS.n94 585
R928 VSS.n384 VSS.n383 585
R929 VSS.n383 VSS.n382 585
R930 VSS.n91 VSS.n90 585
R931 VSS.n381 VSS.n90 585
R932 VSS.n389 VSS.n388 585
R933 VSS.n390 VSS.n389 585
R934 VSS.n88 VSS.n87 585
R935 VSS.n391 VSS.n88 585
R936 VSS.n394 VSS.n393 585
R937 VSS.n393 VSS.n392 585
R938 VSS.n85 VSS.n84 585
R939 VSS.n84 VSS.n82 585
R940 VSS.n399 VSS.n398 585
R941 VSS.n400 VSS.n399 585
R942 VSS.n81 VSS.n80 585
R943 VSS.n401 VSS.n81 585
R944 VSS.n404 VSS.n403 585
R945 VSS.n403 VSS.n402 585
R946 VSS.n78 VSS.n77 585
R947 VSS.n77 VSS.n75 585
R948 VSS.n409 VSS.n408 585
R949 VSS.n410 VSS.n409 585
R950 VSS.n74 VSS.n73 585
R951 VSS.n411 VSS.n74 585
R952 VSS.n414 VSS.n413 585
R953 VSS.n413 VSS.n412 585
R954 VSS.n71 VSS.n70 585
R955 VSS.n70 VSS.n68 585
R956 VSS.n419 VSS.n418 585
R957 VSS.n420 VSS.n419 585
R958 VSS.n67 VSS.n66 585
R959 VSS.n421 VSS.n67 585
R960 VSS.n425 VSS.n424 585
R961 VSS.n424 VSS.n423 585
R962 VSS.n64 VSS.n63 585
R963 VSS.n422 VSS.n63 585
R964 VSS.n431 VSS.n430 585
R965 VSS.n432 VSS.n431 585
R966 VSS.n61 VSS.n60 585
R967 VSS.n433 VSS.n61 585
R968 VSS.n436 VSS.n435 585
R969 VSS.n435 VSS.n434 585
R970 VSS.n437 VSS.n57 585
R971 VSS.n57 VSS.n33 585
R972 VSS.n540 VSS.n30 585
R973 VSS.n33 VSS.n30 585
R974 VSS.n541 VSS.n29 585
R975 VSS.n434 VSS.n29 585
R976 VSS.n542 VSS.n28 585
R977 VSS.n433 VSS.n28 585
R978 VSS.n62 VSS.n26 585
R979 VSS.n432 VSS.n62 585
R980 VSS.n546 VSS.n25 585
R981 VSS.n422 VSS.n25 585
R982 VSS.n547 VSS.n24 585
R983 VSS.n423 VSS.n24 585
R984 VSS.n548 VSS.n23 585
R985 VSS.n421 VSS.n23 585
R986 VSS.n69 VSS.n21 585
R987 VSS.n420 VSS.n69 585
R988 VSS.n552 VSS.n20 585
R989 VSS.n68 VSS.n20 585
R990 VSS.n553 VSS.n19 585
R991 VSS.n412 VSS.n19 585
R992 VSS.n554 VSS.n18 585
R993 VSS.n411 VSS.n18 585
R994 VSS.n76 VSS.n16 585
R995 VSS.n410 VSS.n76 585
R996 VSS.n558 VSS.n15 585
R997 VSS.n75 VSS.n15 585
R998 VSS.n559 VSS.n14 585
R999 VSS.n402 VSS.n14 585
R1000 VSS.n560 VSS.n13 585
R1001 VSS.n401 VSS.n13 585
R1002 VSS.n83 VSS.n11 585
R1003 VSS.n400 VSS.n83 585
R1004 VSS.n564 VSS.n10 585
R1005 VSS.n82 VSS.n10 585
R1006 VSS.n565 VSS.n9 585
R1007 VSS.n392 VSS.n9 585
R1008 VSS.n566 VSS.n8 585
R1009 VSS.n391 VSS.n8 585
R1010 VSS.n89 VSS.n6 585
R1011 VSS.n390 VSS.n89 585
R1012 VSS.n570 VSS.n5 585
R1013 VSS.n381 VSS.n5 585
R1014 VSS.n571 VSS.n4 585
R1015 VSS.n382 VSS.n4 585
R1016 VSS.n572 VSS.n3 585
R1017 VSS.n380 VSS.n3 585
R1018 VSS.n96 VSS.n2 585
R1019 VSS.n379 VSS.n96 585
R1020 VSS.n105 VSS.n103 585
R1021 VSS.n103 VSS.n95 585
R1022 VSS.n370 VSS.n369 585
R1023 VSS.n371 VSS.n370 585
R1024 VSS.n104 VSS.n102 585
R1025 VSS.n110 VSS.n102 585
R1026 VSS.n364 VSS.n363 585
R1027 VSS.n363 VSS.n362 585
R1028 VSS.n108 VSS.n107 585
R1029 VSS.n109 VSS.n108 585
R1030 VSS.n353 VSS.n352 585
R1031 VSS.n354 VSS.n353 585
R1032 VSS.n118 VSS.n117 585
R1033 VSS.n117 VSS.n116 585
R1034 VSS.n348 VSS.n347 585
R1035 VSS.n347 VSS.n346 585
R1036 VSS.n121 VSS.n120 585
R1037 VSS.n122 VSS.n121 585
R1038 VSS.n337 VSS.n336 585
R1039 VSS.n338 VSS.n337 585
R1040 VSS.n130 VSS.n129 585
R1041 VSS.n129 VSS.n128 585
R1042 VSS.n332 VSS.n331 585
R1043 VSS.n331 VSS.n330 585
R1044 VSS.n133 VSS.n132 585
R1045 VSS.n134 VSS.n133 585
R1046 VSS.n321 VSS.n320 585
R1047 VSS.n322 VSS.n321 585
R1048 VSS.n142 VSS.n141 585
R1049 VSS.n141 VSS.n140 585
R1050 VSS.n316 VSS.n315 585
R1051 VSS.n315 VSS.n314 585
R1052 VSS.n145 VSS.n144 585
R1053 VSS.n146 VSS.n145 585
R1054 VSS.n305 VSS.n304 585
R1055 VSS.n306 VSS.n305 585
R1056 VSS.n153 VSS.n152 585
R1057 VSS.n158 VSS.n152 585
R1058 VSS.n300 VSS.n299 585
R1059 VSS.n299 VSS.n298 585
R1060 VSS.n156 VSS.n155 585
R1061 VSS.n157 VSS.n156 585
R1062 VSS.n289 VSS.n288 585
R1063 VSS.n290 VSS.n289 585
R1064 VSS.n538 VSS.n537 585
R1065 VSS.n32 VSS.n31 585
R1066 VSS.n443 VSS.n442 585
R1067 VSS.n445 VSS.n444 585
R1068 VSS.n447 VSS.n446 585
R1069 VSS.n449 VSS.n448 585
R1070 VSS.n451 VSS.n450 585
R1071 VSS.n453 VSS.n452 585
R1072 VSS.n455 VSS.n454 585
R1073 VSS.n457 VSS.n456 585
R1074 VSS.n459 VSS.n458 585
R1075 VSS.n461 VSS.n460 585
R1076 VSS.n463 VSS.n462 585
R1077 VSS.n465 VSS.n464 585
R1078 VSS.n467 VSS.n466 585
R1079 VSS.n469 VSS.n468 585
R1080 VSS.n471 VSS.n470 585
R1081 VSS.n473 VSS.n472 585
R1082 VSS.n475 VSS.n474 585
R1083 VSS.n477 VSS.n476 585
R1084 VSS.n479 VSS.n478 585
R1085 VSS.n481 VSS.n480 585
R1086 VSS.n483 VSS.n482 585
R1087 VSS.n485 VSS.n484 585
R1088 VSS.n487 VSS.n486 585
R1089 VSS.n489 VSS.n488 585
R1090 VSS.n491 VSS.n490 585
R1091 VSS.n493 VSS.n492 585
R1092 VSS.n495 VSS.n494 585
R1093 VSS.n497 VSS.n496 585
R1094 VSS.n499 VSS.n498 585
R1095 VSS.n501 VSS.n500 585
R1096 VSS.n503 VSS.n502 585
R1097 VSS.n505 VSS.n504 585
R1098 VSS.n507 VSS.n506 585
R1099 VSS.n509 VSS.n508 585
R1100 VSS.n511 VSS.n510 585
R1101 VSS.n513 VSS.n512 585
R1102 VSS.n515 VSS.n514 585
R1103 VSS.n517 VSS.n516 585
R1104 VSS.n519 VSS.n518 585
R1105 VSS.n521 VSS.n520 585
R1106 VSS.n523 VSS.n522 585
R1107 VSS.n525 VSS.n524 585
R1108 VSS.n527 VSS.n526 585
R1109 VSS.n529 VSS.n528 585
R1110 VSS.n531 VSS.n530 585
R1111 VSS.n532 VSS.n58 585
R1112 VSS.n534 VSS.n533 585
R1113 VSS.n535 VSS.n534 585
R1114 VSS.n162 VSS.n161 585
R1115 VSS.n193 VSS.n191 585
R1116 VSS.n194 VSS.n190 585
R1117 VSS.n194 VSS.n163 585
R1118 VSS.n197 VSS.n196 585
R1119 VSS.n198 VSS.n189 585
R1120 VSS.n200 VSS.n199 585
R1121 VSS.n202 VSS.n188 585
R1122 VSS.n205 VSS.n204 585
R1123 VSS.n206 VSS.n187 585
R1124 VSS.n208 VSS.n207 585
R1125 VSS.n210 VSS.n186 585
R1126 VSS.n213 VSS.n212 585
R1127 VSS.n214 VSS.n185 585
R1128 VSS.n216 VSS.n215 585
R1129 VSS.n218 VSS.n184 585
R1130 VSS.n221 VSS.n220 585
R1131 VSS.n222 VSS.n183 585
R1132 VSS.n224 VSS.n223 585
R1133 VSS.n226 VSS.n182 585
R1134 VSS.n229 VSS.n228 585
R1135 VSS.n230 VSS.n181 585
R1136 VSS.n232 VSS.n231 585
R1137 VSS.n234 VSS.n180 585
R1138 VSS.n237 VSS.n236 585
R1139 VSS.n238 VSS.n179 585
R1140 VSS.n240 VSS.n239 585
R1141 VSS.n242 VSS.n178 585
R1142 VSS.n245 VSS.n244 585
R1143 VSS.n246 VSS.n177 585
R1144 VSS.n248 VSS.n247 585
R1145 VSS.n250 VSS.n176 585
R1146 VSS.n253 VSS.n252 585
R1147 VSS.n254 VSS.n175 585
R1148 VSS.n256 VSS.n255 585
R1149 VSS.n258 VSS.n174 585
R1150 VSS.n261 VSS.n260 585
R1151 VSS.n262 VSS.n173 585
R1152 VSS.n264 VSS.n263 585
R1153 VSS.n266 VSS.n172 585
R1154 VSS.n269 VSS.n268 585
R1155 VSS.n270 VSS.n171 585
R1156 VSS.n272 VSS.n271 585
R1157 VSS.n274 VSS.n170 585
R1158 VSS.n277 VSS.n276 585
R1159 VSS.n278 VSS.n169 585
R1160 VSS.n280 VSS.n279 585
R1161 VSS.n282 VSS.n168 585
R1162 VSS.n285 VSS.n284 585
R1163 VSS.n286 VSS.n164 585
R1164 VSS.n439 VSS.t8 324.851
R1165 VSS.n165 VSS.t4 324.851
R1166 VSS.n536 VSS.n535 256.663
R1167 VSS.n535 VSS.n34 256.663
R1168 VSS.n535 VSS.n35 256.663
R1169 VSS.n535 VSS.n36 256.663
R1170 VSS.n535 VSS.n37 256.663
R1171 VSS.n535 VSS.n38 256.663
R1172 VSS.n535 VSS.n39 256.663
R1173 VSS.n535 VSS.n40 256.663
R1174 VSS.n535 VSS.n41 256.663
R1175 VSS.n535 VSS.n42 256.663
R1176 VSS.n535 VSS.n43 256.663
R1177 VSS.n535 VSS.n44 256.663
R1178 VSS.n535 VSS.n45 256.663
R1179 VSS.n535 VSS.n46 256.663
R1180 VSS.n535 VSS.n47 256.663
R1181 VSS.n535 VSS.n48 256.663
R1182 VSS.n535 VSS.n49 256.663
R1183 VSS.n535 VSS.n50 256.663
R1184 VSS.n535 VSS.n51 256.663
R1185 VSS.n535 VSS.n52 256.663
R1186 VSS.n535 VSS.n53 256.663
R1187 VSS.n535 VSS.n54 256.663
R1188 VSS.n535 VSS.n55 256.663
R1189 VSS.n535 VSS.n56 256.663
R1190 VSS.n192 VSS.n163 256.663
R1191 VSS.n195 VSS.n163 256.663
R1192 VSS.n201 VSS.n163 256.663
R1193 VSS.n203 VSS.n163 256.663
R1194 VSS.n209 VSS.n163 256.663
R1195 VSS.n211 VSS.n163 256.663
R1196 VSS.n217 VSS.n163 256.663
R1197 VSS.n219 VSS.n163 256.663
R1198 VSS.n225 VSS.n163 256.663
R1199 VSS.n227 VSS.n163 256.663
R1200 VSS.n233 VSS.n163 256.663
R1201 VSS.n235 VSS.n163 256.663
R1202 VSS.n241 VSS.n163 256.663
R1203 VSS.n243 VSS.n163 256.663
R1204 VSS.n249 VSS.n163 256.663
R1205 VSS.n251 VSS.n163 256.663
R1206 VSS.n257 VSS.n163 256.663
R1207 VSS.n259 VSS.n163 256.663
R1208 VSS.n265 VSS.n163 256.663
R1209 VSS.n267 VSS.n163 256.663
R1210 VSS.n273 VSS.n163 256.663
R1211 VSS.n275 VSS.n163 256.663
R1212 VSS.n281 VSS.n163 256.663
R1213 VSS.n283 VSS.n163 256.663
R1214 VSS.n291 VSS.n159 240.244
R1215 VSS.n297 VSS.n159 240.244
R1216 VSS.n297 VSS.n151 240.244
R1217 VSS.n307 VSS.n151 240.244
R1218 VSS.n307 VSS.n147 240.244
R1219 VSS.n313 VSS.n147 240.244
R1220 VSS.n313 VSS.n139 240.244
R1221 VSS.n323 VSS.n139 240.244
R1222 VSS.n323 VSS.n135 240.244
R1223 VSS.n329 VSS.n135 240.244
R1224 VSS.n329 VSS.n127 240.244
R1225 VSS.n339 VSS.n127 240.244
R1226 VSS.n339 VSS.n123 240.244
R1227 VSS.n345 VSS.n123 240.244
R1228 VSS.n345 VSS.n115 240.244
R1229 VSS.n355 VSS.n115 240.244
R1230 VSS.n355 VSS.n111 240.244
R1231 VSS.n361 VSS.n111 240.244
R1232 VSS.n361 VSS.n101 240.244
R1233 VSS.n372 VSS.n101 240.244
R1234 VSS.n372 VSS.n97 240.244
R1235 VSS.n378 VSS.n97 240.244
R1236 VSS.n378 VSS.n94 240.244
R1237 VSS.n383 VSS.n94 240.244
R1238 VSS.n383 VSS.n90 240.244
R1239 VSS.n389 VSS.n90 240.244
R1240 VSS.n389 VSS.n88 240.244
R1241 VSS.n393 VSS.n88 240.244
R1242 VSS.n393 VSS.n84 240.244
R1243 VSS.n399 VSS.n84 240.244
R1244 VSS.n399 VSS.n81 240.244
R1245 VSS.n403 VSS.n81 240.244
R1246 VSS.n403 VSS.n77 240.244
R1247 VSS.n409 VSS.n77 240.244
R1248 VSS.n409 VSS.n74 240.244
R1249 VSS.n413 VSS.n74 240.244
R1250 VSS.n413 VSS.n70 240.244
R1251 VSS.n419 VSS.n70 240.244
R1252 VSS.n419 VSS.n67 240.244
R1253 VSS.n424 VSS.n67 240.244
R1254 VSS.n424 VSS.n63 240.244
R1255 VSS.n431 VSS.n63 240.244
R1256 VSS.n431 VSS.n61 240.244
R1257 VSS.n435 VSS.n61 240.244
R1258 VSS.n435 VSS.n57 240.244
R1259 VSS.n289 VSS.n156 240.244
R1260 VSS.n299 VSS.n156 240.244
R1261 VSS.n299 VSS.n152 240.244
R1262 VSS.n305 VSS.n152 240.244
R1263 VSS.n305 VSS.n145 240.244
R1264 VSS.n315 VSS.n145 240.244
R1265 VSS.n315 VSS.n141 240.244
R1266 VSS.n321 VSS.n141 240.244
R1267 VSS.n321 VSS.n133 240.244
R1268 VSS.n331 VSS.n133 240.244
R1269 VSS.n331 VSS.n129 240.244
R1270 VSS.n337 VSS.n129 240.244
R1271 VSS.n337 VSS.n121 240.244
R1272 VSS.n347 VSS.n121 240.244
R1273 VSS.n347 VSS.n117 240.244
R1274 VSS.n353 VSS.n117 240.244
R1275 VSS.n353 VSS.n108 240.244
R1276 VSS.n363 VSS.n108 240.244
R1277 VSS.n363 VSS.n102 240.244
R1278 VSS.n370 VSS.n102 240.244
R1279 VSS.n370 VSS.n103 240.244
R1280 VSS.n103 VSS.n96 240.244
R1281 VSS.n96 VSS.n3 240.244
R1282 VSS.n4 VSS.n3 240.244
R1283 VSS.n5 VSS.n4 240.244
R1284 VSS.n89 VSS.n5 240.244
R1285 VSS.n89 VSS.n8 240.244
R1286 VSS.n9 VSS.n8 240.244
R1287 VSS.n10 VSS.n9 240.244
R1288 VSS.n83 VSS.n10 240.244
R1289 VSS.n83 VSS.n13 240.244
R1290 VSS.n14 VSS.n13 240.244
R1291 VSS.n15 VSS.n14 240.244
R1292 VSS.n76 VSS.n15 240.244
R1293 VSS.n76 VSS.n18 240.244
R1294 VSS.n19 VSS.n18 240.244
R1295 VSS.n20 VSS.n19 240.244
R1296 VSS.n69 VSS.n20 240.244
R1297 VSS.n69 VSS.n23 240.244
R1298 VSS.n24 VSS.n23 240.244
R1299 VSS.n25 VSS.n24 240.244
R1300 VSS.n62 VSS.n25 240.244
R1301 VSS.n62 VSS.n28 240.244
R1302 VSS.n29 VSS.n28 240.244
R1303 VSS.n30 VSS.n29 240.244
R1304 VSS.n290 VSS.n163 199.474
R1305 VSS.n535 VSS.n33 199.474
R1306 VSS.n194 VSS.n193 163.367
R1307 VSS.n196 VSS.n194 163.367
R1308 VSS.n200 VSS.n189 163.367
R1309 VSS.n204 VSS.n202 163.367
R1310 VSS.n208 VSS.n187 163.367
R1311 VSS.n212 VSS.n210 163.367
R1312 VSS.n216 VSS.n185 163.367
R1313 VSS.n220 VSS.n218 163.367
R1314 VSS.n224 VSS.n183 163.367
R1315 VSS.n228 VSS.n226 163.367
R1316 VSS.n232 VSS.n181 163.367
R1317 VSS.n236 VSS.n234 163.367
R1318 VSS.n240 VSS.n179 163.367
R1319 VSS.n244 VSS.n242 163.367
R1320 VSS.n248 VSS.n177 163.367
R1321 VSS.n252 VSS.n250 163.367
R1322 VSS.n256 VSS.n175 163.367
R1323 VSS.n260 VSS.n258 163.367
R1324 VSS.n264 VSS.n173 163.367
R1325 VSS.n268 VSS.n266 163.367
R1326 VSS.n272 VSS.n171 163.367
R1327 VSS.n276 VSS.n274 163.367
R1328 VSS.n280 VSS.n169 163.367
R1329 VSS.n284 VSS.n282 163.367
R1330 VSS.n534 VSS.n58 163.367
R1331 VSS.n530 VSS.n529 163.367
R1332 VSS.n526 VSS.n525 163.367
R1333 VSS.n522 VSS.n521 163.367
R1334 VSS.n518 VSS.n517 163.367
R1335 VSS.n514 VSS.n513 163.367
R1336 VSS.n510 VSS.n509 163.367
R1337 VSS.n506 VSS.n505 163.367
R1338 VSS.n502 VSS.n501 163.367
R1339 VSS.n498 VSS.n497 163.367
R1340 VSS.n494 VSS.n493 163.367
R1341 VSS.n490 VSS.n489 163.367
R1342 VSS.n486 VSS.n485 163.367
R1343 VSS.n482 VSS.n481 163.367
R1344 VSS.n478 VSS.n477 163.367
R1345 VSS.n474 VSS.n473 163.367
R1346 VSS.n470 VSS.n469 163.367
R1347 VSS.n466 VSS.n465 163.367
R1348 VSS.n462 VSS.n461 163.367
R1349 VSS.n458 VSS.n457 163.367
R1350 VSS.n454 VSS.n453 163.367
R1351 VSS.n450 VSS.n449 163.367
R1352 VSS.n446 VSS.n445 163.367
R1353 VSS.n442 VSS.n32 163.367
R1354 VSS.n439 VSS.t10 133.635
R1355 VSS.n165 VSS.t7 133.635
R1356 VSS.n290 VSS.n157 115.974
R1357 VSS.n298 VSS.n157 115.974
R1358 VSS.n298 VSS.n158 115.974
R1359 VSS.n306 VSS.n146 115.974
R1360 VSS.n314 VSS.n146 115.974
R1361 VSS.n314 VSS.n140 115.974
R1362 VSS.n322 VSS.n140 115.974
R1363 VSS.n322 VSS.n134 115.974
R1364 VSS.n330 VSS.n134 115.974
R1365 VSS.n330 VSS.n128 115.974
R1366 VSS.n338 VSS.n128 115.974
R1367 VSS.n346 VSS.n122 115.974
R1368 VSS.n346 VSS.n116 115.974
R1369 VSS.n354 VSS.n116 115.974
R1370 VSS.n354 VSS.n109 115.974
R1371 VSS.n362 VSS.n109 115.974
R1372 VSS.n362 VSS.n110 115.974
R1373 VSS.n371 VSS.n95 115.974
R1374 VSS.n379 VSS.n95 115.974
R1375 VSS.n380 VSS.n379 115.974
R1376 VSS.n382 VSS.n380 115.974
R1377 VSS.n382 VSS.n381 115.974
R1378 VSS.n391 VSS.n390 115.974
R1379 VSS.n392 VSS.n391 115.974
R1380 VSS.n392 VSS.n82 115.974
R1381 VSS.n400 VSS.n82 115.974
R1382 VSS.n401 VSS.n400 115.974
R1383 VSS.n402 VSS.n401 115.974
R1384 VSS.n410 VSS.n75 115.974
R1385 VSS.n411 VSS.n410 115.974
R1386 VSS.n412 VSS.n411 115.974
R1387 VSS.n412 VSS.n68 115.974
R1388 VSS.n420 VSS.n68 115.974
R1389 VSS.n421 VSS.n420 115.974
R1390 VSS.n423 VSS.n421 115.974
R1391 VSS.n423 VSS.n422 115.974
R1392 VSS.n433 VSS.n432 115.974
R1393 VSS.n434 VSS.n433 115.974
R1394 VSS.n434 VSS.n33 115.974
R1395 VSS.n371 VSS.t1 93.9383
R1396 VSS.n381 VSS.t3 93.9383
R1397 VSS.n158 VSS.t5 89.2994
R1398 VSS.n432 VSS.t9 89.2994
R1399 VSS.n192 VSS.n162 71.676
R1400 VSS.n196 VSS.n195 71.676
R1401 VSS.n201 VSS.n200 71.676
R1402 VSS.n204 VSS.n203 71.676
R1403 VSS.n209 VSS.n208 71.676
R1404 VSS.n212 VSS.n211 71.676
R1405 VSS.n217 VSS.n216 71.676
R1406 VSS.n220 VSS.n219 71.676
R1407 VSS.n225 VSS.n224 71.676
R1408 VSS.n228 VSS.n227 71.676
R1409 VSS.n233 VSS.n232 71.676
R1410 VSS.n236 VSS.n235 71.676
R1411 VSS.n241 VSS.n240 71.676
R1412 VSS.n244 VSS.n243 71.676
R1413 VSS.n249 VSS.n248 71.676
R1414 VSS.n252 VSS.n251 71.676
R1415 VSS.n257 VSS.n256 71.676
R1416 VSS.n260 VSS.n259 71.676
R1417 VSS.n265 VSS.n264 71.676
R1418 VSS.n268 VSS.n267 71.676
R1419 VSS.n273 VSS.n272 71.676
R1420 VSS.n276 VSS.n275 71.676
R1421 VSS.n281 VSS.n280 71.676
R1422 VSS.n284 VSS.n283 71.676
R1423 VSS.n530 VSS.n56 71.676
R1424 VSS.n526 VSS.n55 71.676
R1425 VSS.n522 VSS.n54 71.676
R1426 VSS.n518 VSS.n53 71.676
R1427 VSS.n514 VSS.n52 71.676
R1428 VSS.n510 VSS.n51 71.676
R1429 VSS.n506 VSS.n50 71.676
R1430 VSS.n502 VSS.n49 71.676
R1431 VSS.n498 VSS.n48 71.676
R1432 VSS.n494 VSS.n47 71.676
R1433 VSS.n490 VSS.n46 71.676
R1434 VSS.n486 VSS.n45 71.676
R1435 VSS.n482 VSS.n44 71.676
R1436 VSS.n478 VSS.n43 71.676
R1437 VSS.n474 VSS.n42 71.676
R1438 VSS.n470 VSS.n41 71.676
R1439 VSS.n466 VSS.n40 71.676
R1440 VSS.n462 VSS.n39 71.676
R1441 VSS.n458 VSS.n38 71.676
R1442 VSS.n454 VSS.n37 71.676
R1443 VSS.n450 VSS.n36 71.676
R1444 VSS.n446 VSS.n35 71.676
R1445 VSS.n442 VSS.n34 71.676
R1446 VSS.n537 VSS.n536 71.676
R1447 VSS.n536 VSS.n32 71.676
R1448 VSS.n445 VSS.n34 71.676
R1449 VSS.n449 VSS.n35 71.676
R1450 VSS.n453 VSS.n36 71.676
R1451 VSS.n457 VSS.n37 71.676
R1452 VSS.n461 VSS.n38 71.676
R1453 VSS.n465 VSS.n39 71.676
R1454 VSS.n469 VSS.n40 71.676
R1455 VSS.n473 VSS.n41 71.676
R1456 VSS.n477 VSS.n42 71.676
R1457 VSS.n481 VSS.n43 71.676
R1458 VSS.n485 VSS.n44 71.676
R1459 VSS.n489 VSS.n45 71.676
R1460 VSS.n493 VSS.n46 71.676
R1461 VSS.n497 VSS.n47 71.676
R1462 VSS.n501 VSS.n48 71.676
R1463 VSS.n505 VSS.n49 71.676
R1464 VSS.n509 VSS.n50 71.676
R1465 VSS.n513 VSS.n51 71.676
R1466 VSS.n517 VSS.n52 71.676
R1467 VSS.n521 VSS.n53 71.676
R1468 VSS.n525 VSS.n54 71.676
R1469 VSS.n529 VSS.n55 71.676
R1470 VSS.n58 VSS.n56 71.676
R1471 VSS.n193 VSS.n192 71.676
R1472 VSS.n195 VSS.n189 71.676
R1473 VSS.n202 VSS.n201 71.676
R1474 VSS.n203 VSS.n187 71.676
R1475 VSS.n210 VSS.n209 71.676
R1476 VSS.n211 VSS.n185 71.676
R1477 VSS.n218 VSS.n217 71.676
R1478 VSS.n219 VSS.n183 71.676
R1479 VSS.n226 VSS.n225 71.676
R1480 VSS.n227 VSS.n181 71.676
R1481 VSS.n234 VSS.n233 71.676
R1482 VSS.n235 VSS.n179 71.676
R1483 VSS.n242 VSS.n241 71.676
R1484 VSS.n243 VSS.n177 71.676
R1485 VSS.n250 VSS.n249 71.676
R1486 VSS.n251 VSS.n175 71.676
R1487 VSS.n258 VSS.n257 71.676
R1488 VSS.n259 VSS.n173 71.676
R1489 VSS.n266 VSS.n265 71.676
R1490 VSS.n267 VSS.n171 71.676
R1491 VSS.n274 VSS.n273 71.676
R1492 VSS.n275 VSS.n169 71.676
R1493 VSS.n282 VSS.n281 71.676
R1494 VSS.n283 VSS.n164 71.676
R1495 VSS.n440 VSS.t11 69.441
R1496 VSS.n166 VSS.t6 69.441
R1497 VSS.n338 VSS.t0 66.1049
R1498 VSS.t2 VSS.n75 66.1049
R1499 VSS.n440 VSS.n439 64.1944
R1500 VSS.n166 VSS.n165 64.1944
R1501 VSS.t0 VSS.n122 49.8687
R1502 VSS.n402 VSS.t2 49.8687
R1503 VSS.n441 VSS.n440 34.3278
R1504 VSS.n167 VSS.n166 34.3278
R1505 VSS.n533 VSS.n438 31.4164
R1506 VSS.n539 VSS.n538 31.4164
R1507 VSS.n293 VSS.n161 31.4164
R1508 VSS.n287 VSS.n286 31.4164
R1509 VSS.n306 VSS.t5 26.6742
R1510 VSS.n422 VSS.t9 26.6742
R1511 VSS.n110 VSS.t1 22.0353
R1512 VSS.n390 VSS.t3 22.0353
R1513 VSS.n292 VSS.n160 19.3944
R1514 VSS.n296 VSS.n160 19.3944
R1515 VSS.n296 VSS.n150 19.3944
R1516 VSS.n308 VSS.n150 19.3944
R1517 VSS.n308 VSS.n148 19.3944
R1518 VSS.n312 VSS.n148 19.3944
R1519 VSS.n312 VSS.n138 19.3944
R1520 VSS.n324 VSS.n138 19.3944
R1521 VSS.n324 VSS.n136 19.3944
R1522 VSS.n328 VSS.n136 19.3944
R1523 VSS.n328 VSS.n126 19.3944
R1524 VSS.n340 VSS.n126 19.3944
R1525 VSS.n340 VSS.n124 19.3944
R1526 VSS.n344 VSS.n124 19.3944
R1527 VSS.n344 VSS.n114 19.3944
R1528 VSS.n356 VSS.n114 19.3944
R1529 VSS.n356 VSS.n112 19.3944
R1530 VSS.n360 VSS.n112 19.3944
R1531 VSS.n360 VSS.n100 19.3944
R1532 VSS.n373 VSS.n100 19.3944
R1533 VSS.n373 VSS.n98 19.3944
R1534 VSS.n377 VSS.n98 19.3944
R1535 VSS.n377 VSS.n93 19.3944
R1536 VSS.n384 VSS.n93 19.3944
R1537 VSS.n384 VSS.n91 19.3944
R1538 VSS.n388 VSS.n91 19.3944
R1539 VSS.n388 VSS.n87 19.3944
R1540 VSS.n394 VSS.n87 19.3944
R1541 VSS.n394 VSS.n85 19.3944
R1542 VSS.n398 VSS.n85 19.3944
R1543 VSS.n398 VSS.n80 19.3944
R1544 VSS.n404 VSS.n80 19.3944
R1545 VSS.n404 VSS.n78 19.3944
R1546 VSS.n408 VSS.n78 19.3944
R1547 VSS.n408 VSS.n73 19.3944
R1548 VSS.n414 VSS.n73 19.3944
R1549 VSS.n414 VSS.n71 19.3944
R1550 VSS.n418 VSS.n71 19.3944
R1551 VSS.n418 VSS.n66 19.3944
R1552 VSS.n425 VSS.n66 19.3944
R1553 VSS.n425 VSS.n64 19.3944
R1554 VSS.n430 VSS.n64 19.3944
R1555 VSS.n430 VSS.n60 19.3944
R1556 VSS.n436 VSS.n60 19.3944
R1557 VSS.n437 VSS.n436 19.3944
R1558 VSS.n288 VSS.n155 19.3944
R1559 VSS.n300 VSS.n155 19.3944
R1560 VSS.n300 VSS.n153 19.3944
R1561 VSS.n304 VSS.n153 19.3944
R1562 VSS.n304 VSS.n144 19.3944
R1563 VSS.n316 VSS.n144 19.3944
R1564 VSS.n316 VSS.n142 19.3944
R1565 VSS.n320 VSS.n142 19.3944
R1566 VSS.n320 VSS.n132 19.3944
R1567 VSS.n332 VSS.n132 19.3944
R1568 VSS.n332 VSS.n130 19.3944
R1569 VSS.n336 VSS.n130 19.3944
R1570 VSS.n336 VSS.n120 19.3944
R1571 VSS.n348 VSS.n120 19.3944
R1572 VSS.n348 VSS.n118 19.3944
R1573 VSS.n352 VSS.n118 19.3944
R1574 VSS.n352 VSS.n107 19.3944
R1575 VSS.n364 VSS.n107 19.3944
R1576 VSS.n364 VSS.n104 19.3944
R1577 VSS.n369 VSS.n104 19.3944
R1578 VSS.n369 VSS.n105 19.3944
R1579 VSS.n105 VSS.n2 19.3944
R1580 VSS.n572 VSS.n2 19.3944
R1581 VSS.n572 VSS.n571 19.3944
R1582 VSS.n571 VSS.n570 19.3944
R1583 VSS.n570 VSS.n6 19.3944
R1584 VSS.n566 VSS.n6 19.3944
R1585 VSS.n566 VSS.n565 19.3944
R1586 VSS.n565 VSS.n564 19.3944
R1587 VSS.n564 VSS.n11 19.3944
R1588 VSS.n560 VSS.n11 19.3944
R1589 VSS.n560 VSS.n559 19.3944
R1590 VSS.n559 VSS.n558 19.3944
R1591 VSS.n558 VSS.n16 19.3944
R1592 VSS.n554 VSS.n16 19.3944
R1593 VSS.n554 VSS.n553 19.3944
R1594 VSS.n553 VSS.n552 19.3944
R1595 VSS.n552 VSS.n21 19.3944
R1596 VSS.n548 VSS.n21 19.3944
R1597 VSS.n548 VSS.n547 19.3944
R1598 VSS.n547 VSS.n546 19.3944
R1599 VSS.n546 VSS.n26 19.3944
R1600 VSS.n542 VSS.n26 19.3944
R1601 VSS.n542 VSS.n541 19.3944
R1602 VSS.n541 VSS.n540 19.3944
R1603 VSS.n533 VSS.n532 10.6151
R1604 VSS.n532 VSS.n531 10.6151
R1605 VSS.n531 VSS.n528 10.6151
R1606 VSS.n528 VSS.n527 10.6151
R1607 VSS.n527 VSS.n524 10.6151
R1608 VSS.n524 VSS.n523 10.6151
R1609 VSS.n523 VSS.n520 10.6151
R1610 VSS.n520 VSS.n519 10.6151
R1611 VSS.n519 VSS.n516 10.6151
R1612 VSS.n516 VSS.n515 10.6151
R1613 VSS.n515 VSS.n512 10.6151
R1614 VSS.n512 VSS.n511 10.6151
R1615 VSS.n511 VSS.n508 10.6151
R1616 VSS.n508 VSS.n507 10.6151
R1617 VSS.n507 VSS.n504 10.6151
R1618 VSS.n504 VSS.n503 10.6151
R1619 VSS.n503 VSS.n500 10.6151
R1620 VSS.n500 VSS.n499 10.6151
R1621 VSS.n499 VSS.n496 10.6151
R1622 VSS.n496 VSS.n495 10.6151
R1623 VSS.n495 VSS.n492 10.6151
R1624 VSS.n492 VSS.n491 10.6151
R1625 VSS.n491 VSS.n488 10.6151
R1626 VSS.n488 VSS.n487 10.6151
R1627 VSS.n487 VSS.n484 10.6151
R1628 VSS.n484 VSS.n483 10.6151
R1629 VSS.n483 VSS.n480 10.6151
R1630 VSS.n480 VSS.n479 10.6151
R1631 VSS.n479 VSS.n476 10.6151
R1632 VSS.n476 VSS.n475 10.6151
R1633 VSS.n475 VSS.n472 10.6151
R1634 VSS.n472 VSS.n471 10.6151
R1635 VSS.n471 VSS.n468 10.6151
R1636 VSS.n468 VSS.n467 10.6151
R1637 VSS.n467 VSS.n464 10.6151
R1638 VSS.n464 VSS.n463 10.6151
R1639 VSS.n463 VSS.n460 10.6151
R1640 VSS.n460 VSS.n459 10.6151
R1641 VSS.n459 VSS.n456 10.6151
R1642 VSS.n456 VSS.n455 10.6151
R1643 VSS.n455 VSS.n452 10.6151
R1644 VSS.n452 VSS.n451 10.6151
R1645 VSS.n451 VSS.n448 10.6151
R1646 VSS.n448 VSS.n447 10.6151
R1647 VSS.n447 VSS.n444 10.6151
R1648 VSS.n444 VSS.n443 10.6151
R1649 VSS.n538 VSS.n31 10.6151
R1650 VSS.n191 VSS.n161 10.6151
R1651 VSS.n191 VSS.n190 10.6151
R1652 VSS.n197 VSS.n190 10.6151
R1653 VSS.n198 VSS.n197 10.6151
R1654 VSS.n199 VSS.n198 10.6151
R1655 VSS.n199 VSS.n188 10.6151
R1656 VSS.n205 VSS.n188 10.6151
R1657 VSS.n206 VSS.n205 10.6151
R1658 VSS.n207 VSS.n206 10.6151
R1659 VSS.n207 VSS.n186 10.6151
R1660 VSS.n213 VSS.n186 10.6151
R1661 VSS.n214 VSS.n213 10.6151
R1662 VSS.n215 VSS.n214 10.6151
R1663 VSS.n215 VSS.n184 10.6151
R1664 VSS.n221 VSS.n184 10.6151
R1665 VSS.n222 VSS.n221 10.6151
R1666 VSS.n223 VSS.n222 10.6151
R1667 VSS.n223 VSS.n182 10.6151
R1668 VSS.n229 VSS.n182 10.6151
R1669 VSS.n230 VSS.n229 10.6151
R1670 VSS.n231 VSS.n230 10.6151
R1671 VSS.n231 VSS.n180 10.6151
R1672 VSS.n237 VSS.n180 10.6151
R1673 VSS.n238 VSS.n237 10.6151
R1674 VSS.n239 VSS.n238 10.6151
R1675 VSS.n239 VSS.n178 10.6151
R1676 VSS.n245 VSS.n178 10.6151
R1677 VSS.n246 VSS.n245 10.6151
R1678 VSS.n247 VSS.n246 10.6151
R1679 VSS.n247 VSS.n176 10.6151
R1680 VSS.n253 VSS.n176 10.6151
R1681 VSS.n254 VSS.n253 10.6151
R1682 VSS.n255 VSS.n254 10.6151
R1683 VSS.n255 VSS.n174 10.6151
R1684 VSS.n261 VSS.n174 10.6151
R1685 VSS.n262 VSS.n261 10.6151
R1686 VSS.n263 VSS.n262 10.6151
R1687 VSS.n263 VSS.n172 10.6151
R1688 VSS.n269 VSS.n172 10.6151
R1689 VSS.n270 VSS.n269 10.6151
R1690 VSS.n271 VSS.n270 10.6151
R1691 VSS.n271 VSS.n170 10.6151
R1692 VSS.n277 VSS.n170 10.6151
R1693 VSS.n278 VSS.n277 10.6151
R1694 VSS.n279 VSS.n278 10.6151
R1695 VSS.n279 VSS.n168 10.6151
R1696 VSS.n286 VSS.n285 10.6151
R1697 VSS.n571 VSS.n0 9.3005
R1698 VSS.n570 VSS.n569 9.3005
R1699 VSS.n568 VSS.n6 9.3005
R1700 VSS.n567 VSS.n566 9.3005
R1701 VSS.n565 VSS.n7 9.3005
R1702 VSS.n564 VSS.n563 9.3005
R1703 VSS.n562 VSS.n11 9.3005
R1704 VSS.n561 VSS.n560 9.3005
R1705 VSS.n559 VSS.n12 9.3005
R1706 VSS.n558 VSS.n557 9.3005
R1707 VSS.n556 VSS.n16 9.3005
R1708 VSS.n555 VSS.n554 9.3005
R1709 VSS.n553 VSS.n17 9.3005
R1710 VSS.n552 VSS.n551 9.3005
R1711 VSS.n550 VSS.n21 9.3005
R1712 VSS.n549 VSS.n548 9.3005
R1713 VSS.n547 VSS.n22 9.3005
R1714 VSS.n546 VSS.n545 9.3005
R1715 VSS.n544 VSS.n26 9.3005
R1716 VSS.n543 VSS.n542 9.3005
R1717 VSS.n541 VSS.n27 9.3005
R1718 VSS.n540 VSS.n539 9.3005
R1719 VSS.n293 VSS.n292 9.3005
R1720 VSS.n294 VSS.n160 9.3005
R1721 VSS.n296 VSS.n295 9.3005
R1722 VSS.n150 VSS.n149 9.3005
R1723 VSS.n309 VSS.n308 9.3005
R1724 VSS.n310 VSS.n148 9.3005
R1725 VSS.n312 VSS.n311 9.3005
R1726 VSS.n138 VSS.n137 9.3005
R1727 VSS.n325 VSS.n324 9.3005
R1728 VSS.n326 VSS.n136 9.3005
R1729 VSS.n328 VSS.n327 9.3005
R1730 VSS.n126 VSS.n125 9.3005
R1731 VSS.n341 VSS.n340 9.3005
R1732 VSS.n342 VSS.n124 9.3005
R1733 VSS.n344 VSS.n343 9.3005
R1734 VSS.n114 VSS.n113 9.3005
R1735 VSS.n357 VSS.n356 9.3005
R1736 VSS.n358 VSS.n112 9.3005
R1737 VSS.n360 VSS.n359 9.3005
R1738 VSS.n100 VSS.n99 9.3005
R1739 VSS.n374 VSS.n373 9.3005
R1740 VSS.n375 VSS.n98 9.3005
R1741 VSS.n377 VSS.n376 9.3005
R1742 VSS.n93 VSS.n92 9.3005
R1743 VSS.n385 VSS.n384 9.3005
R1744 VSS.n386 VSS.n91 9.3005
R1745 VSS.n388 VSS.n387 9.3005
R1746 VSS.n87 VSS.n86 9.3005
R1747 VSS.n395 VSS.n394 9.3005
R1748 VSS.n396 VSS.n85 9.3005
R1749 VSS.n398 VSS.n397 9.3005
R1750 VSS.n80 VSS.n79 9.3005
R1751 VSS.n405 VSS.n404 9.3005
R1752 VSS.n406 VSS.n78 9.3005
R1753 VSS.n408 VSS.n407 9.3005
R1754 VSS.n73 VSS.n72 9.3005
R1755 VSS.n415 VSS.n414 9.3005
R1756 VSS.n416 VSS.n71 9.3005
R1757 VSS.n418 VSS.n417 9.3005
R1758 VSS.n66 VSS.n65 9.3005
R1759 VSS.n426 VSS.n425 9.3005
R1760 VSS.n427 VSS.n64 9.3005
R1761 VSS.n430 VSS.n429 9.3005
R1762 VSS.n428 VSS.n60 9.3005
R1763 VSS.n436 VSS.n59 9.3005
R1764 VSS.n438 VSS.n437 9.3005
R1765 VSS.n155 VSS.n154 9.3005
R1766 VSS.n301 VSS.n300 9.3005
R1767 VSS.n302 VSS.n153 9.3005
R1768 VSS.n304 VSS.n303 9.3005
R1769 VSS.n144 VSS.n143 9.3005
R1770 VSS.n317 VSS.n316 9.3005
R1771 VSS.n318 VSS.n142 9.3005
R1772 VSS.n320 VSS.n319 9.3005
R1773 VSS.n132 VSS.n131 9.3005
R1774 VSS.n333 VSS.n332 9.3005
R1775 VSS.n334 VSS.n130 9.3005
R1776 VSS.n336 VSS.n335 9.3005
R1777 VSS.n120 VSS.n119 9.3005
R1778 VSS.n349 VSS.n348 9.3005
R1779 VSS.n350 VSS.n118 9.3005
R1780 VSS.n352 VSS.n351 9.3005
R1781 VSS.n107 VSS.n106 9.3005
R1782 VSS.n365 VSS.n364 9.3005
R1783 VSS.n366 VSS.n104 9.3005
R1784 VSS.n369 VSS.n368 9.3005
R1785 VSS.n367 VSS.n105 9.3005
R1786 VSS.n2 VSS.n1 9.3005
R1787 VSS.n288 VSS.n287 9.3005
R1788 VSS VSS.n572 9.3005
R1789 VSS.n441 VSS.n31 8.89806
R1790 VSS.n285 VSS.n167 8.89806
R1791 VSS.n443 VSS.n441 1.71757
R1792 VSS.n168 VSS.n167 1.71757
R1793 VSS VSS.n0 0.152939
R1794 VSS.n569 VSS.n0 0.152939
R1795 VSS.n569 VSS.n568 0.152939
R1796 VSS.n568 VSS.n567 0.152939
R1797 VSS.n567 VSS.n7 0.152939
R1798 VSS.n563 VSS.n7 0.152939
R1799 VSS.n563 VSS.n562 0.152939
R1800 VSS.n562 VSS.n561 0.152939
R1801 VSS.n561 VSS.n12 0.152939
R1802 VSS.n557 VSS.n12 0.152939
R1803 VSS.n557 VSS.n556 0.152939
R1804 VSS.n556 VSS.n555 0.152939
R1805 VSS.n555 VSS.n17 0.152939
R1806 VSS.n551 VSS.n17 0.152939
R1807 VSS.n551 VSS.n550 0.152939
R1808 VSS.n550 VSS.n549 0.152939
R1809 VSS.n549 VSS.n22 0.152939
R1810 VSS.n545 VSS.n22 0.152939
R1811 VSS.n545 VSS.n544 0.152939
R1812 VSS.n544 VSS.n543 0.152939
R1813 VSS.n543 VSS.n27 0.152939
R1814 VSS.n539 VSS.n27 0.152939
R1815 VSS.n294 VSS.n293 0.152939
R1816 VSS.n295 VSS.n294 0.152939
R1817 VSS.n295 VSS.n149 0.152939
R1818 VSS.n309 VSS.n149 0.152939
R1819 VSS.n310 VSS.n309 0.152939
R1820 VSS.n311 VSS.n310 0.152939
R1821 VSS.n311 VSS.n137 0.152939
R1822 VSS.n325 VSS.n137 0.152939
R1823 VSS.n326 VSS.n325 0.152939
R1824 VSS.n327 VSS.n326 0.152939
R1825 VSS.n327 VSS.n125 0.152939
R1826 VSS.n341 VSS.n125 0.152939
R1827 VSS.n342 VSS.n341 0.152939
R1828 VSS.n343 VSS.n342 0.152939
R1829 VSS.n343 VSS.n113 0.152939
R1830 VSS.n357 VSS.n113 0.152939
R1831 VSS.n358 VSS.n357 0.152939
R1832 VSS.n359 VSS.n358 0.152939
R1833 VSS.n359 VSS.n99 0.152939
R1834 VSS.n374 VSS.n99 0.152939
R1835 VSS.n375 VSS.n374 0.152939
R1836 VSS.n376 VSS.n375 0.152939
R1837 VSS.n376 VSS.n92 0.152939
R1838 VSS.n385 VSS.n92 0.152939
R1839 VSS.n386 VSS.n385 0.152939
R1840 VSS.n387 VSS.n386 0.152939
R1841 VSS.n387 VSS.n86 0.152939
R1842 VSS.n395 VSS.n86 0.152939
R1843 VSS.n396 VSS.n395 0.152939
R1844 VSS.n397 VSS.n396 0.152939
R1845 VSS.n397 VSS.n79 0.152939
R1846 VSS.n405 VSS.n79 0.152939
R1847 VSS.n406 VSS.n405 0.152939
R1848 VSS.n407 VSS.n406 0.152939
R1849 VSS.n407 VSS.n72 0.152939
R1850 VSS.n415 VSS.n72 0.152939
R1851 VSS.n416 VSS.n415 0.152939
R1852 VSS.n417 VSS.n416 0.152939
R1853 VSS.n417 VSS.n65 0.152939
R1854 VSS.n426 VSS.n65 0.152939
R1855 VSS.n427 VSS.n426 0.152939
R1856 VSS.n429 VSS.n427 0.152939
R1857 VSS.n429 VSS.n428 0.152939
R1858 VSS.n428 VSS.n59 0.152939
R1859 VSS.n438 VSS.n59 0.152939
R1860 VSS.n287 VSS.n154 0.152939
R1861 VSS.n301 VSS.n154 0.152939
R1862 VSS.n302 VSS.n301 0.152939
R1863 VSS.n303 VSS.n302 0.152939
R1864 VSS.n303 VSS.n143 0.152939
R1865 VSS.n317 VSS.n143 0.152939
R1866 VSS.n318 VSS.n317 0.152939
R1867 VSS.n319 VSS.n318 0.152939
R1868 VSS.n319 VSS.n131 0.152939
R1869 VSS.n333 VSS.n131 0.152939
R1870 VSS.n334 VSS.n333 0.152939
R1871 VSS.n335 VSS.n334 0.152939
R1872 VSS.n335 VSS.n119 0.152939
R1873 VSS.n349 VSS.n119 0.152939
R1874 VSS.n350 VSS.n349 0.152939
R1875 VSS.n351 VSS.n350 0.152939
R1876 VSS.n351 VSS.n106 0.152939
R1877 VSS.n365 VSS.n106 0.152939
R1878 VSS.n366 VSS.n365 0.152939
R1879 VSS.n368 VSS.n366 0.152939
R1880 VSS.n368 VSS.n367 0.152939
R1881 VSS.n367 VSS.n1 0.152939
R1882 VSS VSS.n1 0.1255
C0 VGN VOUT 4.83106f
C1 VGN VCC 0.047271f
C2 VOUT VCC 1.57787f
C3 VGN VGP 0.038f
C4 VOUT VGP 2.36121f
C5 VGP VCC 4.19161f
C6 VGN VIN 5.37865f
C7 VOUT VIN 5.14834f
C8 VIN VCC 1.67493f
C9 VGP VIN 2.87283f
C10 VGN VSS 6.26762f
C11 VOUT VSS 2.003088f
C12 VIN VSS 3.461631f
C13 VGP VSS 1.408172f
C14 VCC VSS 32.998955f
C15 VGN.t3 VSS 1.70715f
C16 VGN.n0 VSS 0.656395f
C17 VGN.n1 VSS 0.014553f
C18 VGN.n2 VSS 0.023787f
C19 VGN.n3 VSS 0.014553f
C20 VGN.t2 VSS 1.70715f
C21 VGN.n4 VSS 0.027259f
C22 VGN.n5 VSS 0.014553f
C23 VGN.n6 VSS 0.027259f
C24 VGN.t1 VSS 1.85606f
C25 VGN.n7 VSS 0.622867f
C26 VGN.t0 VSS 1.70715f
C27 VGN.n8 VSS 0.640004f
C28 VGN.n9 VSS 0.017972f
C29 VGN.n10 VSS 0.15635f
C30 VGN.n11 VSS 0.014553f
C31 VGN.n12 VSS 0.014553f
C32 VGN.n13 VSS 0.029078f
C33 VGN.n14 VSS 0.011776f
C34 VGN.n15 VSS 0.029078f
C35 VGN.n16 VSS 0.014553f
C36 VGN.n17 VSS 0.014553f
C37 VGN.n18 VSS 0.014553f
C38 VGN.n19 VSS 0.017972f
C39 VGN.n20 VSS 0.596014f
C40 VGN.n21 VSS 0.023086f
C41 VGN.n22 VSS 0.027259f
C42 VGN.n23 VSS 0.014553f
C43 VGN.n24 VSS 0.014553f
C44 VGN.n25 VSS 0.014553f
C45 VGN.n26 VSS 0.018886f
C46 VGN.n27 VSS 0.027259f
C47 VGN.n28 VSS 0.026316f
C48 VGN.n29 VSS 0.023491f
C49 VGN.n30 VSS 0.033694f
C50 VCC.n0 VSS 0.002302f
C51 VCC.n1 VSS 0.002555f
C52 VCC.n2 VSS 0.001853f
C53 VCC.n3 VSS 0.002302f
C54 VCC.n4 VSS 0.002302f
C55 VCC.n5 VSS 0.002302f
C56 VCC.n6 VSS 0.001853f
C57 VCC.n7 VSS 0.002302f
C58 VCC.n8 VSS 0.002302f
C59 VCC.n9 VSS 0.002302f
C60 VCC.n10 VSS 0.002302f
C61 VCC.n11 VSS 0.001853f
C62 VCC.n12 VSS 0.002302f
C63 VCC.n13 VSS 0.002302f
C64 VCC.n14 VSS 0.002302f
C65 VCC.n15 VSS 0.002302f
C66 VCC.n16 VSS 0.001853f
C67 VCC.n17 VSS 0.002302f
C68 VCC.n18 VSS 0.002302f
C69 VCC.n19 VSS 0.002302f
C70 VCC.n20 VSS 0.002302f
C71 VCC.n21 VSS 0.001853f
C72 VCC.n22 VSS 0.002302f
C73 VCC.n23 VSS 0.002302f
C74 VCC.n24 VSS 0.002302f
C75 VCC.n25 VSS 0.002302f
C76 VCC.n26 VSS 0.001538f
C77 VCC.n27 VSS 0.001266f
C78 VCC.n28 VSS 0.004567f
C79 VCC.n29 VSS 0.001566f
C80 VCC.n30 VSS 0.08836f
C81 VCC.n43 VSS 0.001566f
C82 VCC.t11 VSS 0.047552f
C83 VCC.t10 VSS 0.052019f
C84 VCC.t8 VSS 0.187712f
C85 VCC.n44 VSS 0.029121f
C86 VCC.n45 VSS 0.014439f
C87 VCC.n46 VSS 0.002182f
C88 VCC.n47 VSS 0.007903f
C89 VCC.n48 VSS 0.002302f
C90 VCC.n49 VSS 0.001853f
C91 VCC.n50 VSS 0.002302f
C92 VCC.n51 VSS 0.001853f
C93 VCC.n52 VSS 0.002302f
C94 VCC.n53 VSS 0.002302f
C95 VCC.n54 VSS 0.062667f
C96 VCC.n55 VSS 0.002302f
C97 VCC.n56 VSS 0.001853f
C98 VCC.n57 VSS 0.002302f
C99 VCC.n58 VSS 0.001853f
C100 VCC.n59 VSS 0.002302f
C101 VCC.n60 VSS 0.05922f
C102 VCC.n61 VSS 0.002302f
C103 VCC.n62 VSS 0.001853f
C104 VCC.n63 VSS 0.002302f
C105 VCC.n64 VSS 0.001853f
C106 VCC.n65 VSS 0.002302f
C107 VCC.n66 VSS 0.062667f
C108 VCC.n67 VSS 0.002302f
C109 VCC.n68 VSS 0.001853f
C110 VCC.n69 VSS 0.002302f
C111 VCC.n70 VSS 0.001853f
C112 VCC.n71 VSS 0.002302f
C113 VCC.n72 VSS 0.062667f
C114 VCC.n73 VSS 0.002302f
C115 VCC.n74 VSS 0.001853f
C116 VCC.n75 VSS 0.002302f
C117 VCC.n76 VSS 0.001853f
C118 VCC.n77 VSS 0.002302f
C119 VCC.n78 VSS 0.062667f
C120 VCC.n79 VSS 0.002302f
C121 VCC.n80 VSS 0.001853f
C122 VCC.n81 VSS 0.002302f
C123 VCC.n82 VSS 0.001853f
C124 VCC.n83 VSS 0.002302f
C125 VCC.n84 VSS 0.062667f
C126 VCC.n85 VSS 0.002302f
C127 VCC.n86 VSS 0.002302f
C128 VCC.n87 VSS 0.001853f
C129 VCC.n88 VSS 0.001853f
C130 VCC.n89 VSS 0.002302f
C131 VCC.n90 VSS 0.001853f
C132 VCC.n91 VSS 0.002302f
C133 VCC.n92 VSS 0.062667f
C134 VCC.n93 VSS 0.002302f
C135 VCC.n94 VSS 0.001853f
C136 VCC.n95 VSS 0.002302f
C137 VCC.n96 VSS 0.001853f
C138 VCC.n97 VSS 0.002302f
C139 VCC.n98 VSS 0.03478f
C140 VCC.n99 VSS 0.002302f
C141 VCC.n100 VSS 0.001853f
C142 VCC.n101 VSS 0.001853f
C143 VCC.n102 VSS 0.002302f
C144 VCC.n103 VSS 0.001853f
C145 VCC.n104 VSS 0.002302f
C146 VCC.n105 VSS 0.062667f
C147 VCC.t2 VSS 0.031333f
C148 VCC.n106 VSS 0.002302f
C149 VCC.n107 VSS 0.001853f
C150 VCC.n108 VSS 0.002302f
C151 VCC.n109 VSS 0.001853f
C152 VCC.n110 VSS 0.002302f
C153 VCC.n111 VSS 0.062667f
C154 VCC.n112 VSS 0.002302f
C155 VCC.n113 VSS 0.001853f
C156 VCC.n114 VSS 0.002302f
C157 VCC.n115 VSS 0.001853f
C158 VCC.n116 VSS 0.002302f
C159 VCC.n117 VSS 0.062667f
C160 VCC.n118 VSS 0.002302f
C161 VCC.n119 VSS 0.001853f
C162 VCC.n120 VSS 0.002302f
C163 VCC.n121 VSS 0.001853f
C164 VCC.n122 VSS 0.002302f
C165 VCC.n123 VSS 0.032273f
C166 VCC.n124 VSS 0.002302f
C167 VCC.n125 VSS 0.001853f
C168 VCC.n126 VSS 0.002302f
C169 VCC.n127 VSS 0.001853f
C170 VCC.n128 VSS 0.002302f
C171 VCC.n129 VSS 0.062667f
C172 VCC.t5 VSS 0.031333f
C173 VCC.n130 VSS 0.002302f
C174 VCC.n131 VSS 0.001853f
C175 VCC.n132 VSS 0.003079f
C176 VCC.n133 VSS 0.004527f
C177 VCC.n134 VSS 0.121574f
C178 VCC.n135 VSS 0.004527f
C179 VCC.n136 VSS 0.001566f
C180 VCC.n137 VSS 0.001566f
C181 VCC.n138 VSS 0.001566f
C182 VCC.n139 VSS 0.001566f
C183 VCC.n140 VSS 0.001566f
C184 VCC.n141 VSS 0.001566f
C185 VCC.n142 VSS 0.001566f
C186 VCC.n143 VSS 0.001566f
C187 VCC.n144 VSS 0.001566f
C188 VCC.n145 VSS 0.001566f
C189 VCC.n146 VSS 0.001566f
C190 VCC.n147 VSS 0.001566f
C191 VCC.t6 VSS 0.047552f
C192 VCC.t7 VSS 0.052019f
C193 VCC.t4 VSS 0.187712f
C194 VCC.n148 VSS 0.029121f
C195 VCC.n149 VSS 0.014439f
C196 VCC.n151 VSS 0.001566f
C197 VCC.n152 VSS 0.001266f
C198 VCC.n153 VSS 0.002182f
C199 VCC.n154 VSS 0.001082f
C200 VCC.n155 VSS 0.001566f
C201 VCC.n156 VSS 0.001566f
C202 VCC.n158 VSS 0.001566f
C203 VCC.n160 VSS 0.001566f
C204 VCC.n161 VSS 0.001566f
C205 VCC.n162 VSS 0.001566f
C206 VCC.n163 VSS 0.001566f
C207 VCC.n164 VSS 0.001566f
C208 VCC.n166 VSS 0.001566f
C209 VCC.n168 VSS 0.001566f
C210 VCC.n169 VSS 0.001566f
C211 VCC.n170 VSS 0.001566f
C212 VCC.n171 VSS 0.001566f
C213 VCC.n172 VSS 0.001566f
C214 VCC.n174 VSS 0.001566f
C215 VCC.n176 VSS 0.001566f
C216 VCC.n177 VSS 0.001566f
C217 VCC.n178 VSS 0.001566f
C218 VCC.n179 VSS 0.001566f
C219 VCC.n180 VSS 0.001566f
C220 VCC.n182 VSS 0.001566f
C221 VCC.n184 VSS 0.001566f
C222 VCC.n185 VSS 0.001566f
C223 VCC.n186 VSS 0.001566f
C224 VCC.n187 VSS 0.001566f
C225 VCC.n188 VSS 0.001566f
C226 VCC.n190 VSS 0.001566f
C227 VCC.n192 VSS 0.001566f
C228 VCC.n193 VSS 0.001566f
C229 VCC.n194 VSS 0.001566f
C230 VCC.n195 VSS 0.001566f
C231 VCC.n196 VSS 0.001566f
C232 VCC.n198 VSS 0.001566f
C233 VCC.n200 VSS 0.001566f
C234 VCC.n201 VSS 0.001566f
C235 VCC.n202 VSS 0.003079f
C236 VCC.n203 VSS 0.007903f
C237 VCC.n204 VSS 0.001538f
C238 VCC.n205 VSS 0.004567f
C239 VCC.n206 VSS 0.08836f
C240 VCC.n207 VSS 0.004567f
C241 VCC.n208 VSS 0.001538f
C242 VCC.n209 VSS 0.007903f
C243 VCC.n210 VSS 0.002302f
C244 VCC.n211 VSS 0.002302f
C245 VCC.n212 VSS 0.001853f
C246 VCC.n213 VSS 0.002302f
C247 VCC.n214 VSS 0.061727f
C248 VCC.n215 VSS 0.002302f
C249 VCC.n216 VSS 0.001853f
C250 VCC.n217 VSS 0.002302f
C251 VCC.n218 VSS 0.002302f
C252 VCC.n219 VSS 0.002302f
C253 VCC.n220 VSS 0.001853f
C254 VCC.n221 VSS 0.002302f
C255 VCC.n222 VSS 0.062667f
C256 VCC.n223 VSS 0.002302f
C257 VCC.n224 VSS 0.001853f
C258 VCC.n225 VSS 0.002302f
C259 VCC.n226 VSS 0.002302f
C260 VCC.n227 VSS 0.002302f
C261 VCC.n228 VSS 0.001853f
C262 VCC.n229 VSS 0.002302f
C263 VCC.n230 VSS 0.062667f
C264 VCC.n231 VSS 0.002302f
C265 VCC.n232 VSS 0.001853f
C266 VCC.n233 VSS 0.002302f
C267 VCC.n234 VSS 0.002302f
C268 VCC.n235 VSS 0.002302f
C269 VCC.n236 VSS 0.001853f
C270 VCC.n237 VSS 0.002302f
C271 VCC.n238 VSS 0.062667f
C272 VCC.n239 VSS 0.002302f
C273 VCC.n240 VSS 0.001853f
C274 VCC.n241 VSS 0.002302f
C275 VCC.n242 VSS 0.002302f
C276 VCC.n243 VSS 0.002302f
C277 VCC.n244 VSS 0.001853f
C278 VCC.n245 VSS 0.002302f
C279 VCC.n246 VSS 0.05922f
C280 VCC.n247 VSS 0.002302f
C281 VCC.n248 VSS 0.001853f
C282 VCC.n249 VSS 0.002302f
C283 VCC.n250 VSS 0.002302f
C284 VCC.n251 VSS 0.002302f
C285 VCC.n252 VSS 0.002302f
C286 VCC.n253 VSS 0.001853f
C287 VCC.n254 VSS 0.002302f
C288 VCC.n255 VSS 0.062667f
C289 VCC.n256 VSS 0.002302f
C290 VCC.n257 VSS 0.001853f
C291 VCC.n258 VSS 0.002302f
C292 VCC.n259 VSS 0.002302f
C293 VCC.n260 VSS 0.002302f
C294 VCC.n261 VSS 0.001853f
C295 VCC.n262 VSS 0.002302f
C296 VCC.n263 VSS 0.062667f
C297 VCC.n264 VSS 0.002302f
C298 VCC.n265 VSS 0.002302f
C299 VCC.n266 VSS 0.001853f
C300 VCC.n267 VSS 0.002302f
C301 VCC.n268 VSS 0.002302f
C302 VCC.n269 VSS 0.002302f
C303 VCC.n270 VSS 0.002302f
C304 VCC.n271 VSS 0.001853f
C305 VCC.n272 VSS 0.002302f
C306 VCC.n273 VSS 0.042927f
C307 VCC.t0 VSS 0.031333f
C308 VCC.n274 VSS 0.051074f
C309 VCC.n275 VSS 0.002302f
C310 VCC.n276 VSS 0.001853f
C311 VCC.n277 VSS 0.002302f
C312 VCC.n278 VSS 0.002302f
C313 VCC.n279 VSS 0.002302f
C314 VCC.n280 VSS 0.001853f
C315 VCC.n281 VSS 0.002302f
C316 VCC.n282 VSS 0.002302f
C317 VCC.n283 VSS 0.062667f
C318 VCC.n284 VSS 0.062667f
C319 VCC.n285 VSS 0.002302f
C320 VCC.n286 VSS 0.001853f
C321 VCC.n287 VSS 0.002302f
C322 VCC.n288 VSS 0.002302f
C323 VCC.n289 VSS 0.002302f
C324 VCC.n290 VSS 0.001853f
C325 VCC.n291 VSS 0.002302f
C326 VCC.n292 VSS 0.042927f
C327 VCC.t3 VSS 0.031333f
C328 VCC.n293 VSS 0.002302f
C329 VCC.n294 VSS 0.051074f
C330 VCC.n295 VSS 0.062667f
C331 VCC.n296 VSS 0.002302f
C332 VCC.n297 VSS 0.001853f
C333 VCC.n298 VSS 0.002302f
C334 VCC.n299 VSS 0.002302f
C335 VCC.n300 VSS 0.002302f
C336 VCC.n301 VSS 0.001853f
C337 VCC.n302 VSS 0.002302f
C338 VCC.n303 VSS 0.062667f
C339 VCC.n304 VSS 0.002302f
C340 VCC.n305 VSS 0.062667f
C341 VCC.t1 VSS 0.031333f
C342 VCC.n306 VSS 0.03478f
C343 VCC.n307 VSS 0.002302f
C344 VCC.n308 VSS 0.001853f
C345 VCC.n309 VSS 0.002302f
C346 VCC.n310 VSS 0.002302f
C347 VCC.n311 VSS 0.002302f
C348 VCC.n312 VSS 0.001853f
C349 VCC.n313 VSS 0.002302f
C350 VCC.n314 VSS 0.062667f
C351 VCC.n315 VSS 0.002302f
C352 VCC.n316 VSS 0.062667f
C353 VCC.n317 VSS 0.062667f
C354 VCC.n318 VSS 0.002302f
C355 VCC.n319 VSS 0.001853f
C356 VCC.n320 VSS 0.002302f
C357 VCC.n321 VSS 0.002302f
C358 VCC.n322 VSS 0.002302f
C359 VCC.n323 VSS 0.001853f
C360 VCC.n324 VSS 0.002302f
C361 VCC.n325 VSS 0.062667f
C362 VCC.n326 VSS 0.002302f
C363 VCC.n327 VSS 0.062667f
C364 VCC.n328 VSS 0.062667f
C365 VCC.n329 VSS 0.061727f
C366 VCC.t9 VSS 0.031333f
C367 VCC.n330 VSS 0.032273f
C368 VCC.n331 VSS 0.002302f
C369 VCC.n332 VSS 0.001853f
C370 VCC.n333 VSS 0.002302f
C371 VCC.n334 VSS 0.002302f
C372 VCC.n335 VSS 0.002302f
C373 VCC.n336 VSS 0.001853f
C374 VCC.n337 VSS 0.001538f
C375 VCC.n338 VSS 0.004567f
C376 VCC.n339 VSS 0.004527f
C377 VCC.n340 VSS 0.003079f
C378 VCC.n341 VSS 0.001566f
C379 VCC.n342 VSS 0.001566f
C380 VCC.n343 VSS 0.001566f
C381 VCC.n344 VSS 0.001566f
C382 VCC.n345 VSS 0.001566f
C383 VCC.n346 VSS 0.001566f
C384 VCC.n347 VSS 0.001566f
C385 VCC.n348 VSS 0.001566f
C386 VCC.n349 VSS 0.001566f
C387 VCC.n350 VSS 0.001566f
C388 VCC.n351 VSS 0.001566f
C389 VCC.n352 VSS 0.001566f
C390 VCC.n353 VSS 0.001566f
C391 VCC.n354 VSS 0.001566f
C392 VCC.n355 VSS 0.001566f
C393 VCC.n356 VSS 0.001566f
C394 VCC.n357 VSS 0.001566f
C395 VCC.n358 VSS 0.001566f
C396 VCC.n359 VSS 0.001566f
C397 VCC.n360 VSS 0.001566f
C398 VCC.n361 VSS 0.001566f
C399 VCC.n362 VSS 0.001566f
C400 VCC.n363 VSS 0.001566f
C401 VCC.n364 VSS 0.001566f
C402 VCC.n365 VSS 0.001566f
C403 VCC.n366 VSS 0.001566f
C404 VCC.n367 VSS 0.001566f
C405 VCC.n368 VSS 0.001566f
C406 VCC.n369 VSS 0.001566f
C407 VCC.n370 VSS 0.001566f
C408 VCC.n371 VSS 0.001566f
C409 VCC.n372 VSS 0.001566f
C410 VCC.n373 VSS 0.001566f
C411 VCC.n374 VSS 0.001566f
C412 VCC.n375 VSS 0.001566f
C413 VCC.n376 VSS 0.001566f
C414 VCC.n377 VSS 0.001566f
C415 VCC.n378 VSS 0.001566f
C416 VCC.n379 VSS 0.001566f
C417 VCC.n380 VSS 0.001566f
C418 VCC.n381 VSS 0.001566f
C419 VCC.n382 VSS 0.001566f
C420 VCC.n383 VSS 0.001566f
C421 VCC.n384 VSS 0.001566f
C422 VCC.n385 VSS 0.001566f
C423 VCC.n386 VSS 0.001082f
C424 VCC.n387 VSS 0.001566f
C425 VCC.n389 VSS 0.121574f
C426 VCC.n390 VSS 0.004527f
C427 VCC.n391 VSS 0.003079f
C428 VCC.n392 VSS 0.007903f
C429 VCC.n393 VSS 0.002302f
C430 VCC.n394 VSS 0.001853f
C431 VCC.n395 VSS 0.001853f
C432 VCC.n396 VSS 0.001853f
C433 VCC.n397 VSS 0.002302f
C434 VCC.n398 VSS 0.002302f
C435 VCC.n399 VSS 0.002302f
C436 VCC.n400 VSS 0.001853f
C437 VCC.n401 VSS 0.001853f
C438 VCC.n402 VSS 0.001853f
C439 VCC.n403 VSS 0.002302f
C440 VCC.n404 VSS 0.002302f
C441 VCC.n405 VSS 0.002302f
C442 VCC.n406 VSS 0.001853f
C443 VCC.n407 VSS 0.001853f
C444 VCC.n408 VSS 0.001853f
C445 VCC.n409 VSS 0.002302f
C446 VCC.n410 VSS 0.002302f
C447 VCC.n411 VSS 0.002302f
C448 VCC.n412 VSS 0.001853f
C449 VCC.n413 VSS 0.001853f
C450 VCC.n414 VSS 0.001853f
C451 VCC.n415 VSS 0.002302f
C452 VCC.n416 VSS 0.002302f
C453 VCC.n417 VSS 0.002302f
C454 VCC.n418 VSS 0.001853f
C455 VCC.n419 VSS 0.001853f
C456 VCC.n420 VSS 0.001853f
C457 VIN.t5 VSS 0.904311f
C458 VIN.t4 VSS 0.10523f
C459 VIN.t7 VSS 0.10523f
C460 VIN.n0 VSS 0.650228f
C461 VIN.n1 VSS 1.23915f
C462 VIN.t6 VSS 0.885461f
C463 VIN.n2 VSS 0.810787f
C464 VIN.t1 VSS 2.42843f
C465 VIN.t0 VSS 0.21464f
C466 VIN.t2 VSS 0.21464f
C467 VIN.n3 VSS 1.88411f
C468 VIN.n4 VSS 0.930891f
C469 VIN.t3 VSS 2.40428f
C470 VIN.n5 VSS 0.419753f
C471 VOUT.t5 VSS 0.139935f
C472 VOUT.t7 VSS 0.139935f
C473 VOUT.n0 VSS 0.989892f
C474 VOUT.t4 VSS 0.139935f
C475 VOUT.t6 VSS 0.139935f
C476 VOUT.n1 VSS 0.966459f
C477 VOUT.n2 VSS 1.55524f
C478 VOUT.t3 VSS 0.285429f
C479 VOUT.t0 VSS 0.285429f
C480 VOUT.n3 VSS 2.60625f
C481 VOUT.t2 VSS 0.285429f
C482 VOUT.t1 VSS 0.285429f
C483 VOUT.n4 VSS 2.57696f
C484 VOUT.n5 VSS 1.49794f
C485 VGP.n0 VSS 0.039188f
C486 VGP.t1 VSS 1.42113f
C487 VGP.n1 VSS 0.053363f
C488 VGP.n2 VSS 0.029724f
C489 VGP.t3 VSS 1.42113f
C490 VGP.n3 VSS 0.524568f
C491 VGP.n4 VSS 0.029724f
C492 VGP.n5 VSS 0.043392f
C493 VGP.n6 VSS 0.284563f
C494 VGP.t0 VSS 1.42113f
C495 VGP.t2 VSS 1.64436f
C496 VGP.n7 VSS 0.595425f
C497 VGP.n8 VSS 0.606086f
C498 VGP.n9 VSS 0.038166f
C499 VGP.n10 VSS 0.055398f
C500 VGP.n11 VSS 0.029724f
C501 VGP.n12 VSS 0.029724f
C502 VGP.n13 VSS 0.029724f
C503 VGP.n14 VSS 0.043392f
C504 VGP.n15 VSS 0.055398f
C505 VGP.n16 VSS 0.038166f
C506 VGP.n17 VSS 0.029724f
C507 VGP.n18 VSS 0.029724f
C508 VGP.n19 VSS 0.045277f
C509 VGP.n20 VSS 0.058796f
C510 VGP.n21 VSS 0.030023f
C511 VGP.n22 VSS 0.029724f
C512 VGP.n23 VSS 0.029724f
C513 VGP.n24 VSS 0.029724f
C514 VGP.n25 VSS 0.055398f
C515 VGP.n26 VSS 0.031055f
C516 VGP.n27 VSS 0.610498f
C517 VGP.n28 VSS 0.055371f
.ends

