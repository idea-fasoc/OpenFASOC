* NGSPICE file created from diff_pair_sample_0926.ext - technology: sky130A

.subckt diff_pair_sample_0926 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=3.71
X1 VDD2.t9 VN.t0 VTAIL.t17 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=3.71
X2 VDD2.t8 VN.t1 VTAIL.t6 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=3.71
X3 B.t11 B.t9 B.t10 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=3.71
X4 VDD2.t7 VN.t2 VTAIL.t1 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X5 VDD1.t8 VP.t1 VTAIL.t12 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=3.71
X6 VTAIL.t9 VP.t2 VDD1.t7 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X7 VDD1.t6 VP.t3 VTAIL.t8 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X8 B.t8 B.t6 B.t7 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=3.71
X9 VTAIL.t19 VN.t3 VDD2.t6 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X10 VDD2.t5 VN.t4 VTAIL.t0 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=3.71
X11 VDD2.t4 VN.t5 VTAIL.t5 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=3.71
X12 VTAIL.t18 VN.t6 VDD2.t3 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X13 VTAIL.t2 VN.t7 VDD2.t2 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X14 VTAIL.t13 VP.t4 VDD1.t5 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X15 VTAIL.t15 VP.t5 VDD1.t4 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X16 VDD1.t3 VP.t6 VTAIL.t16 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=3.71
X17 VDD2.t1 VN.t8 VTAIL.t3 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X18 B.t5 B.t3 B.t4 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=3.71
X19 VDD1.t2 VP.t7 VTAIL.t7 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=3.71
X20 VTAIL.t4 VN.t9 VDD2.t0 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X21 VDD1.t1 VP.t8 VTAIL.t11 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
X22 B.t2 B.t0 B.t1 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=3.71
X23 VTAIL.t10 VP.t9 VDD1.t0 w_n5818_n1158# sky130_fd_pr__pfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=3.71
R0 VP.n33 VP.n32 161.3
R1 VP.n34 VP.n29 161.3
R2 VP.n36 VP.n35 161.3
R3 VP.n37 VP.n28 161.3
R4 VP.n39 VP.n38 161.3
R5 VP.n40 VP.n27 161.3
R6 VP.n42 VP.n41 161.3
R7 VP.n43 VP.n26 161.3
R8 VP.n45 VP.n44 161.3
R9 VP.n46 VP.n25 161.3
R10 VP.n48 VP.n47 161.3
R11 VP.n49 VP.n24 161.3
R12 VP.n51 VP.n50 161.3
R13 VP.n52 VP.n23 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n22 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n21 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n20 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n19 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n68 VP.n18 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n125 VP.n124 161.3
R26 VP.n123 VP.n1 161.3
R27 VP.n122 VP.n121 161.3
R28 VP.n120 VP.n2 161.3
R29 VP.n119 VP.n118 161.3
R30 VP.n117 VP.n3 161.3
R31 VP.n116 VP.n115 161.3
R32 VP.n114 VP.n4 161.3
R33 VP.n113 VP.n112 161.3
R34 VP.n110 VP.n5 161.3
R35 VP.n109 VP.n108 161.3
R36 VP.n107 VP.n6 161.3
R37 VP.n106 VP.n105 161.3
R38 VP.n104 VP.n7 161.3
R39 VP.n103 VP.n102 161.3
R40 VP.n101 VP.n8 161.3
R41 VP.n100 VP.n99 161.3
R42 VP.n98 VP.n9 161.3
R43 VP.n97 VP.n96 161.3
R44 VP.n95 VP.n10 161.3
R45 VP.n94 VP.n93 161.3
R46 VP.n92 VP.n11 161.3
R47 VP.n91 VP.n90 161.3
R48 VP.n89 VP.n12 161.3
R49 VP.n88 VP.n87 161.3
R50 VP.n85 VP.n13 161.3
R51 VP.n84 VP.n83 161.3
R52 VP.n82 VP.n14 161.3
R53 VP.n81 VP.n80 161.3
R54 VP.n79 VP.n15 161.3
R55 VP.n78 VP.n77 161.3
R56 VP.n76 VP.n16 161.3
R57 VP.n75 VP.n74 161.3
R58 VP.n73 VP.n72 86.1527
R59 VP.n126 VP.n0 86.1527
R60 VP.n71 VP.n17 86.1527
R61 VP.n31 VP.n30 72.9615
R62 VP.n72 VP.n71 50.8251
R63 VP.n80 VP.n79 46.321
R64 VP.n118 VP.n2 46.321
R65 VP.n63 VP.n19 46.321
R66 VP.n93 VP.n92 42.4359
R67 VP.n105 VP.n6 42.4359
R68 VP.n50 VP.n23 42.4359
R69 VP.n38 VP.n37 42.4359
R70 VP.n93 VP.n10 38.5509
R71 VP.n105 VP.n104 38.5509
R72 VP.n50 VP.n49 38.5509
R73 VP.n38 VP.n27 38.5509
R74 VP.n30 VP.t6 38.2987
R75 VP.n80 VP.n14 34.6658
R76 VP.n118 VP.n117 34.6658
R77 VP.n63 VP.n62 34.6658
R78 VP.n74 VP.n16 24.4675
R79 VP.n78 VP.n16 24.4675
R80 VP.n79 VP.n78 24.4675
R81 VP.n84 VP.n14 24.4675
R82 VP.n85 VP.n84 24.4675
R83 VP.n87 VP.n12 24.4675
R84 VP.n91 VP.n12 24.4675
R85 VP.n92 VP.n91 24.4675
R86 VP.n97 VP.n10 24.4675
R87 VP.n98 VP.n97 24.4675
R88 VP.n99 VP.n98 24.4675
R89 VP.n99 VP.n8 24.4675
R90 VP.n103 VP.n8 24.4675
R91 VP.n104 VP.n103 24.4675
R92 VP.n109 VP.n6 24.4675
R93 VP.n110 VP.n109 24.4675
R94 VP.n112 VP.n110 24.4675
R95 VP.n116 VP.n4 24.4675
R96 VP.n117 VP.n116 24.4675
R97 VP.n122 VP.n2 24.4675
R98 VP.n123 VP.n122 24.4675
R99 VP.n124 VP.n123 24.4675
R100 VP.n67 VP.n19 24.4675
R101 VP.n68 VP.n67 24.4675
R102 VP.n69 VP.n68 24.4675
R103 VP.n54 VP.n23 24.4675
R104 VP.n55 VP.n54 24.4675
R105 VP.n57 VP.n55 24.4675
R106 VP.n61 VP.n21 24.4675
R107 VP.n62 VP.n61 24.4675
R108 VP.n42 VP.n27 24.4675
R109 VP.n43 VP.n42 24.4675
R110 VP.n44 VP.n43 24.4675
R111 VP.n44 VP.n25 24.4675
R112 VP.n48 VP.n25 24.4675
R113 VP.n49 VP.n48 24.4675
R114 VP.n32 VP.n29 24.4675
R115 VP.n36 VP.n29 24.4675
R116 VP.n37 VP.n36 24.4675
R117 VP.n86 VP.n85 22.5101
R118 VP.n111 VP.n4 22.5101
R119 VP.n56 VP.n21 22.5101
R120 VP.n99 VP.t8 6.17166
R121 VP.n73 VP.t1 6.17166
R122 VP.n86 VP.t5 6.17166
R123 VP.n111 VP.t9 6.17166
R124 VP.n0 VP.t7 6.17166
R125 VP.n44 VP.t3 6.17166
R126 VP.n17 VP.t0 6.17166
R127 VP.n56 VP.t2 6.17166
R128 VP.n31 VP.t4 6.17166
R129 VP.n74 VP.n73 3.91522
R130 VP.n124 VP.n0 3.91522
R131 VP.n69 VP.n17 3.91522
R132 VP.n33 VP.n30 3.3454
R133 VP.n87 VP.n86 1.95786
R134 VP.n112 VP.n111 1.95786
R135 VP.n57 VP.n56 1.95786
R136 VP.n32 VP.n31 1.95786
R137 VP.n71 VP.n70 0.354971
R138 VP.n75 VP.n72 0.354971
R139 VP.n126 VP.n125 0.354971
R140 VP VP.n126 0.26696
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n28 0.189894
R144 VP.n39 VP.n28 0.189894
R145 VP.n40 VP.n39 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n41 VP.n26 0.189894
R148 VP.n45 VP.n26 0.189894
R149 VP.n46 VP.n45 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n47 VP.n24 0.189894
R152 VP.n51 VP.n24 0.189894
R153 VP.n52 VP.n51 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n53 VP.n22 0.189894
R156 VP.n58 VP.n22 0.189894
R157 VP.n59 VP.n58 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n60 VP.n20 0.189894
R160 VP.n64 VP.n20 0.189894
R161 VP.n65 VP.n64 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n66 VP.n18 0.189894
R164 VP.n70 VP.n18 0.189894
R165 VP.n76 VP.n75 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n77 VP.n15 0.189894
R168 VP.n81 VP.n15 0.189894
R169 VP.n82 VP.n81 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n83 VP.n13 0.189894
R172 VP.n88 VP.n13 0.189894
R173 VP.n89 VP.n88 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n90 VP.n11 0.189894
R176 VP.n94 VP.n11 0.189894
R177 VP.n95 VP.n94 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n96 VP.n9 0.189894
R180 VP.n100 VP.n9 0.189894
R181 VP.n101 VP.n100 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n102 VP.n7 0.189894
R184 VP.n106 VP.n7 0.189894
R185 VP.n107 VP.n106 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n108 VP.n5 0.189894
R188 VP.n113 VP.n5 0.189894
R189 VP.n114 VP.n113 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n115 VP.n3 0.189894
R192 VP.n119 VP.n3 0.189894
R193 VP.n120 VP.n119 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n121 VP.n1 0.189894
R196 VP.n125 VP.n1 0.189894
R197 VTAIL.n16 VTAIL.t14 656.701
R198 VTAIL.n11 VTAIL.t5 656.701
R199 VTAIL.n17 VTAIL.t6 656.699
R200 VTAIL.n2 VTAIL.t7 656.699
R201 VTAIL.n15 VTAIL.n14 622.485
R202 VTAIL.n13 VTAIL.n12 622.485
R203 VTAIL.n10 VTAIL.n9 622.485
R204 VTAIL.n8 VTAIL.n7 622.485
R205 VTAIL.n19 VTAIL.n18 622.484
R206 VTAIL.n1 VTAIL.n0 622.484
R207 VTAIL.n4 VTAIL.n3 622.484
R208 VTAIL.n6 VTAIL.n5 622.484
R209 VTAIL.n18 VTAIL.t1 34.2163
R210 VTAIL.n18 VTAIL.t2 34.2163
R211 VTAIL.n0 VTAIL.t0 34.2163
R212 VTAIL.n0 VTAIL.t4 34.2163
R213 VTAIL.n3 VTAIL.t11 34.2163
R214 VTAIL.n3 VTAIL.t10 34.2163
R215 VTAIL.n5 VTAIL.t12 34.2163
R216 VTAIL.n5 VTAIL.t15 34.2163
R217 VTAIL.n14 VTAIL.t8 34.2163
R218 VTAIL.n14 VTAIL.t9 34.2163
R219 VTAIL.n12 VTAIL.t16 34.2163
R220 VTAIL.n12 VTAIL.t13 34.2163
R221 VTAIL.n9 VTAIL.t3 34.2163
R222 VTAIL.n9 VTAIL.t18 34.2163
R223 VTAIL.n7 VTAIL.t17 34.2163
R224 VTAIL.n7 VTAIL.t19 34.2163
R225 VTAIL.n8 VTAIL.n6 20.1514
R226 VTAIL.n17 VTAIL.n16 16.6686
R227 VTAIL.n10 VTAIL.n8 3.48326
R228 VTAIL.n11 VTAIL.n10 3.48326
R229 VTAIL.n15 VTAIL.n13 3.48326
R230 VTAIL.n16 VTAIL.n15 3.48326
R231 VTAIL.n6 VTAIL.n4 3.48326
R232 VTAIL.n4 VTAIL.n2 3.48326
R233 VTAIL.n19 VTAIL.n17 3.48326
R234 VTAIL VTAIL.n1 2.67076
R235 VTAIL.n13 VTAIL.n11 2.21171
R236 VTAIL.n2 VTAIL.n1 2.21171
R237 VTAIL VTAIL.n19 0.813
R238 VDD1.n1 VDD1.t3 676.861
R239 VDD1.n3 VDD1.t8 676.861
R240 VDD1.n5 VDD1.n4 641.718
R241 VDD1.n7 VDD1.n6 639.163
R242 VDD1.n1 VDD1.n0 639.163
R243 VDD1.n3 VDD1.n2 639.163
R244 VDD1.n7 VDD1.n5 43.4018
R245 VDD1.n6 VDD1.t7 34.2163
R246 VDD1.n6 VDD1.t9 34.2163
R247 VDD1.n0 VDD1.t5 34.2163
R248 VDD1.n0 VDD1.t6 34.2163
R249 VDD1.n4 VDD1.t0 34.2163
R250 VDD1.n4 VDD1.t2 34.2163
R251 VDD1.n2 VDD1.t4 34.2163
R252 VDD1.n2 VDD1.t1 34.2163
R253 VDD1 VDD1.n7 2.55438
R254 VDD1 VDD1.n1 0.929379
R255 VDD1.n5 VDD1.n3 0.815844
R256 VN.n108 VN.n107 161.3
R257 VN.n106 VN.n56 161.3
R258 VN.n105 VN.n104 161.3
R259 VN.n103 VN.n57 161.3
R260 VN.n102 VN.n101 161.3
R261 VN.n100 VN.n58 161.3
R262 VN.n99 VN.n98 161.3
R263 VN.n97 VN.n59 161.3
R264 VN.n96 VN.n95 161.3
R265 VN.n94 VN.n60 161.3
R266 VN.n93 VN.n92 161.3
R267 VN.n91 VN.n62 161.3
R268 VN.n90 VN.n89 161.3
R269 VN.n88 VN.n63 161.3
R270 VN.n87 VN.n86 161.3
R271 VN.n85 VN.n64 161.3
R272 VN.n84 VN.n83 161.3
R273 VN.n82 VN.n65 161.3
R274 VN.n81 VN.n80 161.3
R275 VN.n79 VN.n66 161.3
R276 VN.n78 VN.n77 161.3
R277 VN.n76 VN.n67 161.3
R278 VN.n75 VN.n74 161.3
R279 VN.n73 VN.n68 161.3
R280 VN.n72 VN.n71 161.3
R281 VN.n53 VN.n52 161.3
R282 VN.n51 VN.n1 161.3
R283 VN.n50 VN.n49 161.3
R284 VN.n48 VN.n2 161.3
R285 VN.n47 VN.n46 161.3
R286 VN.n45 VN.n3 161.3
R287 VN.n44 VN.n43 161.3
R288 VN.n42 VN.n4 161.3
R289 VN.n41 VN.n40 161.3
R290 VN.n38 VN.n5 161.3
R291 VN.n37 VN.n36 161.3
R292 VN.n35 VN.n6 161.3
R293 VN.n34 VN.n33 161.3
R294 VN.n32 VN.n7 161.3
R295 VN.n31 VN.n30 161.3
R296 VN.n29 VN.n8 161.3
R297 VN.n28 VN.n27 161.3
R298 VN.n26 VN.n9 161.3
R299 VN.n25 VN.n24 161.3
R300 VN.n23 VN.n10 161.3
R301 VN.n22 VN.n21 161.3
R302 VN.n20 VN.n11 161.3
R303 VN.n19 VN.n18 161.3
R304 VN.n17 VN.n12 161.3
R305 VN.n16 VN.n15 161.3
R306 VN.n54 VN.n0 86.1527
R307 VN.n109 VN.n55 86.1527
R308 VN.n14 VN.n13 72.9614
R309 VN.n70 VN.n69 72.9614
R310 VN VN.n109 50.9904
R311 VN.n46 VN.n2 46.321
R312 VN.n101 VN.n57 46.321
R313 VN.n21 VN.n20 42.4359
R314 VN.n33 VN.n6 42.4359
R315 VN.n77 VN.n76 42.4359
R316 VN.n89 VN.n62 42.4359
R317 VN.n21 VN.n10 38.5509
R318 VN.n33 VN.n32 38.5509
R319 VN.n77 VN.n66 38.5509
R320 VN.n89 VN.n88 38.5509
R321 VN.n69 VN.t5 38.2989
R322 VN.n13 VN.t4 38.2989
R323 VN.n46 VN.n45 34.6658
R324 VN.n101 VN.n100 34.6658
R325 VN.n15 VN.n12 24.4675
R326 VN.n19 VN.n12 24.4675
R327 VN.n20 VN.n19 24.4675
R328 VN.n25 VN.n10 24.4675
R329 VN.n26 VN.n25 24.4675
R330 VN.n27 VN.n26 24.4675
R331 VN.n27 VN.n8 24.4675
R332 VN.n31 VN.n8 24.4675
R333 VN.n32 VN.n31 24.4675
R334 VN.n37 VN.n6 24.4675
R335 VN.n38 VN.n37 24.4675
R336 VN.n40 VN.n38 24.4675
R337 VN.n44 VN.n4 24.4675
R338 VN.n45 VN.n44 24.4675
R339 VN.n50 VN.n2 24.4675
R340 VN.n51 VN.n50 24.4675
R341 VN.n52 VN.n51 24.4675
R342 VN.n76 VN.n75 24.4675
R343 VN.n75 VN.n68 24.4675
R344 VN.n71 VN.n68 24.4675
R345 VN.n88 VN.n87 24.4675
R346 VN.n87 VN.n64 24.4675
R347 VN.n83 VN.n64 24.4675
R348 VN.n83 VN.n82 24.4675
R349 VN.n82 VN.n81 24.4675
R350 VN.n81 VN.n66 24.4675
R351 VN.n100 VN.n99 24.4675
R352 VN.n99 VN.n59 24.4675
R353 VN.n95 VN.n94 24.4675
R354 VN.n94 VN.n93 24.4675
R355 VN.n93 VN.n62 24.4675
R356 VN.n107 VN.n106 24.4675
R357 VN.n106 VN.n105 24.4675
R358 VN.n105 VN.n57 24.4675
R359 VN.n39 VN.n4 22.5101
R360 VN.n61 VN.n59 22.5101
R361 VN.n27 VN.t2 6.17166
R362 VN.n14 VN.t9 6.17166
R363 VN.n39 VN.t7 6.17166
R364 VN.n0 VN.t1 6.17166
R365 VN.n83 VN.t8 6.17166
R366 VN.n70 VN.t6 6.17166
R367 VN.n61 VN.t3 6.17166
R368 VN.n55 VN.t0 6.17166
R369 VN.n52 VN.n0 3.91522
R370 VN.n107 VN.n55 3.91522
R371 VN.n72 VN.n69 3.34541
R372 VN.n16 VN.n13 3.34541
R373 VN.n15 VN.n14 1.95786
R374 VN.n40 VN.n39 1.95786
R375 VN.n71 VN.n70 1.95786
R376 VN.n95 VN.n61 1.95786
R377 VN.n109 VN.n108 0.354971
R378 VN.n54 VN.n53 0.354971
R379 VN VN.n54 0.26696
R380 VN.n108 VN.n56 0.189894
R381 VN.n104 VN.n56 0.189894
R382 VN.n104 VN.n103 0.189894
R383 VN.n103 VN.n102 0.189894
R384 VN.n102 VN.n58 0.189894
R385 VN.n98 VN.n58 0.189894
R386 VN.n98 VN.n97 0.189894
R387 VN.n97 VN.n96 0.189894
R388 VN.n96 VN.n60 0.189894
R389 VN.n92 VN.n60 0.189894
R390 VN.n92 VN.n91 0.189894
R391 VN.n91 VN.n90 0.189894
R392 VN.n90 VN.n63 0.189894
R393 VN.n86 VN.n63 0.189894
R394 VN.n86 VN.n85 0.189894
R395 VN.n85 VN.n84 0.189894
R396 VN.n84 VN.n65 0.189894
R397 VN.n80 VN.n65 0.189894
R398 VN.n80 VN.n79 0.189894
R399 VN.n79 VN.n78 0.189894
R400 VN.n78 VN.n67 0.189894
R401 VN.n74 VN.n67 0.189894
R402 VN.n74 VN.n73 0.189894
R403 VN.n73 VN.n72 0.189894
R404 VN.n17 VN.n16 0.189894
R405 VN.n18 VN.n17 0.189894
R406 VN.n18 VN.n11 0.189894
R407 VN.n22 VN.n11 0.189894
R408 VN.n23 VN.n22 0.189894
R409 VN.n24 VN.n23 0.189894
R410 VN.n24 VN.n9 0.189894
R411 VN.n28 VN.n9 0.189894
R412 VN.n29 VN.n28 0.189894
R413 VN.n30 VN.n29 0.189894
R414 VN.n30 VN.n7 0.189894
R415 VN.n34 VN.n7 0.189894
R416 VN.n35 VN.n34 0.189894
R417 VN.n36 VN.n35 0.189894
R418 VN.n36 VN.n5 0.189894
R419 VN.n41 VN.n5 0.189894
R420 VN.n42 VN.n41 0.189894
R421 VN.n43 VN.n42 0.189894
R422 VN.n43 VN.n3 0.189894
R423 VN.n47 VN.n3 0.189894
R424 VN.n48 VN.n47 0.189894
R425 VN.n49 VN.n48 0.189894
R426 VN.n49 VN.n1 0.189894
R427 VN.n53 VN.n1 0.189894
R428 VDD2.n1 VDD2.t5 676.861
R429 VDD2.n4 VDD2.t9 673.379
R430 VDD2.n3 VDD2.n2 641.718
R431 VDD2 VDD2.n7 641.717
R432 VDD2.n6 VDD2.n5 639.163
R433 VDD2.n1 VDD2.n0 639.163
R434 VDD2.n4 VDD2.n3 41.0774
R435 VDD2.n7 VDD2.t3 34.2163
R436 VDD2.n7 VDD2.t4 34.2163
R437 VDD2.n5 VDD2.t6 34.2163
R438 VDD2.n5 VDD2.t1 34.2163
R439 VDD2.n2 VDD2.t2 34.2163
R440 VDD2.n2 VDD2.t8 34.2163
R441 VDD2.n0 VDD2.t0 34.2163
R442 VDD2.n0 VDD2.t7 34.2163
R443 VDD2.n6 VDD2.n4 3.48326
R444 VDD2 VDD2.n6 0.929379
R445 VDD2.n3 VDD2.n1 0.815844
R446 B.n150 B.t7 725.689
R447 B.n340 B.t10 725.689
R448 B.n54 B.t2 725.689
R449 B.n46 B.t5 725.689
R450 B.n151 B.t8 647.337
R451 B.n341 B.t11 647.337
R452 B.n55 B.t1 647.337
R453 B.n47 B.t4 647.337
R454 B.n357 B.n140 585
R455 B.n356 B.n355 585
R456 B.n354 B.n141 585
R457 B.n353 B.n352 585
R458 B.n351 B.n142 585
R459 B.n350 B.n349 585
R460 B.n348 B.n143 585
R461 B.n347 B.n346 585
R462 B.n345 B.n144 585
R463 B.n344 B.n343 585
R464 B.n339 B.n145 585
R465 B.n338 B.n337 585
R466 B.n336 B.n146 585
R467 B.n335 B.n334 585
R468 B.n333 B.n147 585
R469 B.n332 B.n331 585
R470 B.n330 B.n148 585
R471 B.n329 B.n328 585
R472 B.n327 B.n149 585
R473 B.n325 B.n324 585
R474 B.n323 B.n152 585
R475 B.n322 B.n321 585
R476 B.n320 B.n153 585
R477 B.n319 B.n318 585
R478 B.n317 B.n154 585
R479 B.n316 B.n315 585
R480 B.n314 B.n155 585
R481 B.n313 B.n312 585
R482 B.n359 B.n358 585
R483 B.n360 B.n139 585
R484 B.n362 B.n361 585
R485 B.n363 B.n138 585
R486 B.n365 B.n364 585
R487 B.n366 B.n137 585
R488 B.n368 B.n367 585
R489 B.n369 B.n136 585
R490 B.n371 B.n370 585
R491 B.n372 B.n135 585
R492 B.n374 B.n373 585
R493 B.n375 B.n134 585
R494 B.n377 B.n376 585
R495 B.n378 B.n133 585
R496 B.n380 B.n379 585
R497 B.n381 B.n132 585
R498 B.n383 B.n382 585
R499 B.n384 B.n131 585
R500 B.n386 B.n385 585
R501 B.n387 B.n130 585
R502 B.n389 B.n388 585
R503 B.n390 B.n129 585
R504 B.n392 B.n391 585
R505 B.n393 B.n128 585
R506 B.n395 B.n394 585
R507 B.n396 B.n127 585
R508 B.n398 B.n397 585
R509 B.n399 B.n126 585
R510 B.n401 B.n400 585
R511 B.n402 B.n125 585
R512 B.n404 B.n403 585
R513 B.n405 B.n124 585
R514 B.n407 B.n406 585
R515 B.n408 B.n123 585
R516 B.n410 B.n409 585
R517 B.n411 B.n122 585
R518 B.n413 B.n412 585
R519 B.n414 B.n121 585
R520 B.n416 B.n415 585
R521 B.n417 B.n120 585
R522 B.n419 B.n418 585
R523 B.n420 B.n119 585
R524 B.n422 B.n421 585
R525 B.n423 B.n118 585
R526 B.n425 B.n424 585
R527 B.n426 B.n117 585
R528 B.n428 B.n427 585
R529 B.n429 B.n116 585
R530 B.n431 B.n430 585
R531 B.n432 B.n115 585
R532 B.n434 B.n433 585
R533 B.n435 B.n114 585
R534 B.n437 B.n436 585
R535 B.n438 B.n113 585
R536 B.n440 B.n439 585
R537 B.n441 B.n112 585
R538 B.n443 B.n442 585
R539 B.n444 B.n111 585
R540 B.n446 B.n445 585
R541 B.n447 B.n110 585
R542 B.n449 B.n448 585
R543 B.n450 B.n109 585
R544 B.n452 B.n451 585
R545 B.n453 B.n108 585
R546 B.n455 B.n454 585
R547 B.n456 B.n107 585
R548 B.n458 B.n457 585
R549 B.n459 B.n106 585
R550 B.n461 B.n460 585
R551 B.n462 B.n105 585
R552 B.n464 B.n463 585
R553 B.n465 B.n104 585
R554 B.n467 B.n466 585
R555 B.n468 B.n103 585
R556 B.n470 B.n469 585
R557 B.n471 B.n102 585
R558 B.n473 B.n472 585
R559 B.n474 B.n101 585
R560 B.n476 B.n475 585
R561 B.n477 B.n100 585
R562 B.n479 B.n478 585
R563 B.n480 B.n99 585
R564 B.n482 B.n481 585
R565 B.n483 B.n98 585
R566 B.n485 B.n484 585
R567 B.n486 B.n97 585
R568 B.n488 B.n487 585
R569 B.n489 B.n96 585
R570 B.n491 B.n490 585
R571 B.n492 B.n95 585
R572 B.n494 B.n493 585
R573 B.n495 B.n94 585
R574 B.n497 B.n496 585
R575 B.n498 B.n93 585
R576 B.n500 B.n499 585
R577 B.n501 B.n92 585
R578 B.n503 B.n502 585
R579 B.n504 B.n91 585
R580 B.n506 B.n505 585
R581 B.n507 B.n90 585
R582 B.n509 B.n508 585
R583 B.n510 B.n89 585
R584 B.n512 B.n511 585
R585 B.n513 B.n88 585
R586 B.n515 B.n514 585
R587 B.n516 B.n87 585
R588 B.n518 B.n517 585
R589 B.n519 B.n86 585
R590 B.n521 B.n520 585
R591 B.n522 B.n85 585
R592 B.n524 B.n523 585
R593 B.n525 B.n84 585
R594 B.n527 B.n526 585
R595 B.n528 B.n83 585
R596 B.n530 B.n529 585
R597 B.n531 B.n82 585
R598 B.n533 B.n532 585
R599 B.n534 B.n81 585
R600 B.n536 B.n535 585
R601 B.n537 B.n80 585
R602 B.n539 B.n538 585
R603 B.n540 B.n79 585
R604 B.n542 B.n541 585
R605 B.n543 B.n78 585
R606 B.n545 B.n544 585
R607 B.n546 B.n77 585
R608 B.n548 B.n547 585
R609 B.n549 B.n76 585
R610 B.n551 B.n550 585
R611 B.n552 B.n75 585
R612 B.n554 B.n553 585
R613 B.n555 B.n74 585
R614 B.n557 B.n556 585
R615 B.n558 B.n73 585
R616 B.n560 B.n559 585
R617 B.n561 B.n72 585
R618 B.n563 B.n562 585
R619 B.n564 B.n71 585
R620 B.n566 B.n565 585
R621 B.n567 B.n70 585
R622 B.n569 B.n568 585
R623 B.n570 B.n69 585
R624 B.n572 B.n571 585
R625 B.n573 B.n68 585
R626 B.n575 B.n574 585
R627 B.n576 B.n67 585
R628 B.n578 B.n577 585
R629 B.n579 B.n66 585
R630 B.n581 B.n580 585
R631 B.n582 B.n65 585
R632 B.n584 B.n583 585
R633 B.n585 B.n64 585
R634 B.n587 B.n586 585
R635 B.n588 B.n63 585
R636 B.n590 B.n589 585
R637 B.n591 B.n62 585
R638 B.n593 B.n592 585
R639 B.n594 B.n61 585
R640 B.n596 B.n595 585
R641 B.n597 B.n60 585
R642 B.n641 B.n640 585
R643 B.n639 B.n42 585
R644 B.n638 B.n637 585
R645 B.n636 B.n43 585
R646 B.n635 B.n634 585
R647 B.n633 B.n44 585
R648 B.n632 B.n631 585
R649 B.n630 B.n45 585
R650 B.n629 B.n628 585
R651 B.n627 B.n626 585
R652 B.n625 B.n49 585
R653 B.n624 B.n623 585
R654 B.n622 B.n50 585
R655 B.n621 B.n620 585
R656 B.n619 B.n51 585
R657 B.n618 B.n617 585
R658 B.n616 B.n52 585
R659 B.n615 B.n614 585
R660 B.n613 B.n53 585
R661 B.n611 B.n610 585
R662 B.n609 B.n56 585
R663 B.n608 B.n607 585
R664 B.n606 B.n57 585
R665 B.n605 B.n604 585
R666 B.n603 B.n58 585
R667 B.n602 B.n601 585
R668 B.n600 B.n59 585
R669 B.n599 B.n598 585
R670 B.n642 B.n41 585
R671 B.n644 B.n643 585
R672 B.n645 B.n40 585
R673 B.n647 B.n646 585
R674 B.n648 B.n39 585
R675 B.n650 B.n649 585
R676 B.n651 B.n38 585
R677 B.n653 B.n652 585
R678 B.n654 B.n37 585
R679 B.n656 B.n655 585
R680 B.n657 B.n36 585
R681 B.n659 B.n658 585
R682 B.n660 B.n35 585
R683 B.n662 B.n661 585
R684 B.n663 B.n34 585
R685 B.n665 B.n664 585
R686 B.n666 B.n33 585
R687 B.n668 B.n667 585
R688 B.n669 B.n32 585
R689 B.n671 B.n670 585
R690 B.n672 B.n31 585
R691 B.n674 B.n673 585
R692 B.n675 B.n30 585
R693 B.n677 B.n676 585
R694 B.n678 B.n29 585
R695 B.n680 B.n679 585
R696 B.n681 B.n28 585
R697 B.n683 B.n682 585
R698 B.n684 B.n27 585
R699 B.n686 B.n685 585
R700 B.n687 B.n26 585
R701 B.n689 B.n688 585
R702 B.n690 B.n25 585
R703 B.n692 B.n691 585
R704 B.n693 B.n24 585
R705 B.n695 B.n694 585
R706 B.n696 B.n23 585
R707 B.n698 B.n697 585
R708 B.n699 B.n22 585
R709 B.n701 B.n700 585
R710 B.n702 B.n21 585
R711 B.n704 B.n703 585
R712 B.n705 B.n20 585
R713 B.n707 B.n706 585
R714 B.n708 B.n19 585
R715 B.n710 B.n709 585
R716 B.n711 B.n18 585
R717 B.n713 B.n712 585
R718 B.n714 B.n17 585
R719 B.n716 B.n715 585
R720 B.n717 B.n16 585
R721 B.n719 B.n718 585
R722 B.n720 B.n15 585
R723 B.n722 B.n721 585
R724 B.n723 B.n14 585
R725 B.n725 B.n724 585
R726 B.n726 B.n13 585
R727 B.n728 B.n727 585
R728 B.n729 B.n12 585
R729 B.n731 B.n730 585
R730 B.n732 B.n11 585
R731 B.n734 B.n733 585
R732 B.n735 B.n10 585
R733 B.n737 B.n736 585
R734 B.n738 B.n9 585
R735 B.n740 B.n739 585
R736 B.n741 B.n8 585
R737 B.n743 B.n742 585
R738 B.n744 B.n7 585
R739 B.n746 B.n745 585
R740 B.n747 B.n6 585
R741 B.n749 B.n748 585
R742 B.n750 B.n5 585
R743 B.n752 B.n751 585
R744 B.n753 B.n4 585
R745 B.n755 B.n754 585
R746 B.n756 B.n3 585
R747 B.n758 B.n757 585
R748 B.n759 B.n0 585
R749 B.n2 B.n1 585
R750 B.n196 B.n195 585
R751 B.n197 B.n194 585
R752 B.n199 B.n198 585
R753 B.n200 B.n193 585
R754 B.n202 B.n201 585
R755 B.n203 B.n192 585
R756 B.n205 B.n204 585
R757 B.n206 B.n191 585
R758 B.n208 B.n207 585
R759 B.n209 B.n190 585
R760 B.n211 B.n210 585
R761 B.n212 B.n189 585
R762 B.n214 B.n213 585
R763 B.n215 B.n188 585
R764 B.n217 B.n216 585
R765 B.n218 B.n187 585
R766 B.n220 B.n219 585
R767 B.n221 B.n186 585
R768 B.n223 B.n222 585
R769 B.n224 B.n185 585
R770 B.n226 B.n225 585
R771 B.n227 B.n184 585
R772 B.n229 B.n228 585
R773 B.n230 B.n183 585
R774 B.n232 B.n231 585
R775 B.n233 B.n182 585
R776 B.n235 B.n234 585
R777 B.n236 B.n181 585
R778 B.n238 B.n237 585
R779 B.n239 B.n180 585
R780 B.n241 B.n240 585
R781 B.n242 B.n179 585
R782 B.n244 B.n243 585
R783 B.n245 B.n178 585
R784 B.n247 B.n246 585
R785 B.n248 B.n177 585
R786 B.n250 B.n249 585
R787 B.n251 B.n176 585
R788 B.n253 B.n252 585
R789 B.n254 B.n175 585
R790 B.n256 B.n255 585
R791 B.n257 B.n174 585
R792 B.n259 B.n258 585
R793 B.n260 B.n173 585
R794 B.n262 B.n261 585
R795 B.n263 B.n172 585
R796 B.n265 B.n264 585
R797 B.n266 B.n171 585
R798 B.n268 B.n267 585
R799 B.n269 B.n170 585
R800 B.n271 B.n270 585
R801 B.n272 B.n169 585
R802 B.n274 B.n273 585
R803 B.n275 B.n168 585
R804 B.n277 B.n276 585
R805 B.n278 B.n167 585
R806 B.n280 B.n279 585
R807 B.n281 B.n166 585
R808 B.n283 B.n282 585
R809 B.n284 B.n165 585
R810 B.n286 B.n285 585
R811 B.n287 B.n164 585
R812 B.n289 B.n288 585
R813 B.n290 B.n163 585
R814 B.n292 B.n291 585
R815 B.n293 B.n162 585
R816 B.n295 B.n294 585
R817 B.n296 B.n161 585
R818 B.n298 B.n297 585
R819 B.n299 B.n160 585
R820 B.n301 B.n300 585
R821 B.n302 B.n159 585
R822 B.n304 B.n303 585
R823 B.n305 B.n158 585
R824 B.n307 B.n306 585
R825 B.n308 B.n157 585
R826 B.n310 B.n309 585
R827 B.n311 B.n156 585
R828 B.n312 B.n311 468.476
R829 B.n358 B.n357 468.476
R830 B.n598 B.n597 468.476
R831 B.n640 B.n41 468.476
R832 B.n761 B.n760 256.663
R833 B.n760 B.n759 235.042
R834 B.n760 B.n2 235.042
R835 B.n150 B.t6 209.957
R836 B.n340 B.t9 209.957
R837 B.n54 B.t0 209.957
R838 B.n46 B.t3 209.957
R839 B.n312 B.n155 163.367
R840 B.n316 B.n155 163.367
R841 B.n317 B.n316 163.367
R842 B.n318 B.n317 163.367
R843 B.n318 B.n153 163.367
R844 B.n322 B.n153 163.367
R845 B.n323 B.n322 163.367
R846 B.n324 B.n323 163.367
R847 B.n324 B.n149 163.367
R848 B.n329 B.n149 163.367
R849 B.n330 B.n329 163.367
R850 B.n331 B.n330 163.367
R851 B.n331 B.n147 163.367
R852 B.n335 B.n147 163.367
R853 B.n336 B.n335 163.367
R854 B.n337 B.n336 163.367
R855 B.n337 B.n145 163.367
R856 B.n344 B.n145 163.367
R857 B.n345 B.n344 163.367
R858 B.n346 B.n345 163.367
R859 B.n346 B.n143 163.367
R860 B.n350 B.n143 163.367
R861 B.n351 B.n350 163.367
R862 B.n352 B.n351 163.367
R863 B.n352 B.n141 163.367
R864 B.n356 B.n141 163.367
R865 B.n357 B.n356 163.367
R866 B.n597 B.n596 163.367
R867 B.n596 B.n61 163.367
R868 B.n592 B.n61 163.367
R869 B.n592 B.n591 163.367
R870 B.n591 B.n590 163.367
R871 B.n590 B.n63 163.367
R872 B.n586 B.n63 163.367
R873 B.n586 B.n585 163.367
R874 B.n585 B.n584 163.367
R875 B.n584 B.n65 163.367
R876 B.n580 B.n65 163.367
R877 B.n580 B.n579 163.367
R878 B.n579 B.n578 163.367
R879 B.n578 B.n67 163.367
R880 B.n574 B.n67 163.367
R881 B.n574 B.n573 163.367
R882 B.n573 B.n572 163.367
R883 B.n572 B.n69 163.367
R884 B.n568 B.n69 163.367
R885 B.n568 B.n567 163.367
R886 B.n567 B.n566 163.367
R887 B.n566 B.n71 163.367
R888 B.n562 B.n71 163.367
R889 B.n562 B.n561 163.367
R890 B.n561 B.n560 163.367
R891 B.n560 B.n73 163.367
R892 B.n556 B.n73 163.367
R893 B.n556 B.n555 163.367
R894 B.n555 B.n554 163.367
R895 B.n554 B.n75 163.367
R896 B.n550 B.n75 163.367
R897 B.n550 B.n549 163.367
R898 B.n549 B.n548 163.367
R899 B.n548 B.n77 163.367
R900 B.n544 B.n77 163.367
R901 B.n544 B.n543 163.367
R902 B.n543 B.n542 163.367
R903 B.n542 B.n79 163.367
R904 B.n538 B.n79 163.367
R905 B.n538 B.n537 163.367
R906 B.n537 B.n536 163.367
R907 B.n536 B.n81 163.367
R908 B.n532 B.n81 163.367
R909 B.n532 B.n531 163.367
R910 B.n531 B.n530 163.367
R911 B.n530 B.n83 163.367
R912 B.n526 B.n83 163.367
R913 B.n526 B.n525 163.367
R914 B.n525 B.n524 163.367
R915 B.n524 B.n85 163.367
R916 B.n520 B.n85 163.367
R917 B.n520 B.n519 163.367
R918 B.n519 B.n518 163.367
R919 B.n518 B.n87 163.367
R920 B.n514 B.n87 163.367
R921 B.n514 B.n513 163.367
R922 B.n513 B.n512 163.367
R923 B.n512 B.n89 163.367
R924 B.n508 B.n89 163.367
R925 B.n508 B.n507 163.367
R926 B.n507 B.n506 163.367
R927 B.n506 B.n91 163.367
R928 B.n502 B.n91 163.367
R929 B.n502 B.n501 163.367
R930 B.n501 B.n500 163.367
R931 B.n500 B.n93 163.367
R932 B.n496 B.n93 163.367
R933 B.n496 B.n495 163.367
R934 B.n495 B.n494 163.367
R935 B.n494 B.n95 163.367
R936 B.n490 B.n95 163.367
R937 B.n490 B.n489 163.367
R938 B.n489 B.n488 163.367
R939 B.n488 B.n97 163.367
R940 B.n484 B.n97 163.367
R941 B.n484 B.n483 163.367
R942 B.n483 B.n482 163.367
R943 B.n482 B.n99 163.367
R944 B.n478 B.n99 163.367
R945 B.n478 B.n477 163.367
R946 B.n477 B.n476 163.367
R947 B.n476 B.n101 163.367
R948 B.n472 B.n101 163.367
R949 B.n472 B.n471 163.367
R950 B.n471 B.n470 163.367
R951 B.n470 B.n103 163.367
R952 B.n466 B.n103 163.367
R953 B.n466 B.n465 163.367
R954 B.n465 B.n464 163.367
R955 B.n464 B.n105 163.367
R956 B.n460 B.n105 163.367
R957 B.n460 B.n459 163.367
R958 B.n459 B.n458 163.367
R959 B.n458 B.n107 163.367
R960 B.n454 B.n107 163.367
R961 B.n454 B.n453 163.367
R962 B.n453 B.n452 163.367
R963 B.n452 B.n109 163.367
R964 B.n448 B.n109 163.367
R965 B.n448 B.n447 163.367
R966 B.n447 B.n446 163.367
R967 B.n446 B.n111 163.367
R968 B.n442 B.n111 163.367
R969 B.n442 B.n441 163.367
R970 B.n441 B.n440 163.367
R971 B.n440 B.n113 163.367
R972 B.n436 B.n113 163.367
R973 B.n436 B.n435 163.367
R974 B.n435 B.n434 163.367
R975 B.n434 B.n115 163.367
R976 B.n430 B.n115 163.367
R977 B.n430 B.n429 163.367
R978 B.n429 B.n428 163.367
R979 B.n428 B.n117 163.367
R980 B.n424 B.n117 163.367
R981 B.n424 B.n423 163.367
R982 B.n423 B.n422 163.367
R983 B.n422 B.n119 163.367
R984 B.n418 B.n119 163.367
R985 B.n418 B.n417 163.367
R986 B.n417 B.n416 163.367
R987 B.n416 B.n121 163.367
R988 B.n412 B.n121 163.367
R989 B.n412 B.n411 163.367
R990 B.n411 B.n410 163.367
R991 B.n410 B.n123 163.367
R992 B.n406 B.n123 163.367
R993 B.n406 B.n405 163.367
R994 B.n405 B.n404 163.367
R995 B.n404 B.n125 163.367
R996 B.n400 B.n125 163.367
R997 B.n400 B.n399 163.367
R998 B.n399 B.n398 163.367
R999 B.n398 B.n127 163.367
R1000 B.n394 B.n127 163.367
R1001 B.n394 B.n393 163.367
R1002 B.n393 B.n392 163.367
R1003 B.n392 B.n129 163.367
R1004 B.n388 B.n129 163.367
R1005 B.n388 B.n387 163.367
R1006 B.n387 B.n386 163.367
R1007 B.n386 B.n131 163.367
R1008 B.n382 B.n131 163.367
R1009 B.n382 B.n381 163.367
R1010 B.n381 B.n380 163.367
R1011 B.n380 B.n133 163.367
R1012 B.n376 B.n133 163.367
R1013 B.n376 B.n375 163.367
R1014 B.n375 B.n374 163.367
R1015 B.n374 B.n135 163.367
R1016 B.n370 B.n135 163.367
R1017 B.n370 B.n369 163.367
R1018 B.n369 B.n368 163.367
R1019 B.n368 B.n137 163.367
R1020 B.n364 B.n137 163.367
R1021 B.n364 B.n363 163.367
R1022 B.n363 B.n362 163.367
R1023 B.n362 B.n139 163.367
R1024 B.n358 B.n139 163.367
R1025 B.n640 B.n639 163.367
R1026 B.n639 B.n638 163.367
R1027 B.n638 B.n43 163.367
R1028 B.n634 B.n43 163.367
R1029 B.n634 B.n633 163.367
R1030 B.n633 B.n632 163.367
R1031 B.n632 B.n45 163.367
R1032 B.n628 B.n45 163.367
R1033 B.n628 B.n627 163.367
R1034 B.n627 B.n49 163.367
R1035 B.n623 B.n49 163.367
R1036 B.n623 B.n622 163.367
R1037 B.n622 B.n621 163.367
R1038 B.n621 B.n51 163.367
R1039 B.n617 B.n51 163.367
R1040 B.n617 B.n616 163.367
R1041 B.n616 B.n615 163.367
R1042 B.n615 B.n53 163.367
R1043 B.n610 B.n53 163.367
R1044 B.n610 B.n609 163.367
R1045 B.n609 B.n608 163.367
R1046 B.n608 B.n57 163.367
R1047 B.n604 B.n57 163.367
R1048 B.n604 B.n603 163.367
R1049 B.n603 B.n602 163.367
R1050 B.n602 B.n59 163.367
R1051 B.n598 B.n59 163.367
R1052 B.n644 B.n41 163.367
R1053 B.n645 B.n644 163.367
R1054 B.n646 B.n645 163.367
R1055 B.n646 B.n39 163.367
R1056 B.n650 B.n39 163.367
R1057 B.n651 B.n650 163.367
R1058 B.n652 B.n651 163.367
R1059 B.n652 B.n37 163.367
R1060 B.n656 B.n37 163.367
R1061 B.n657 B.n656 163.367
R1062 B.n658 B.n657 163.367
R1063 B.n658 B.n35 163.367
R1064 B.n662 B.n35 163.367
R1065 B.n663 B.n662 163.367
R1066 B.n664 B.n663 163.367
R1067 B.n664 B.n33 163.367
R1068 B.n668 B.n33 163.367
R1069 B.n669 B.n668 163.367
R1070 B.n670 B.n669 163.367
R1071 B.n670 B.n31 163.367
R1072 B.n674 B.n31 163.367
R1073 B.n675 B.n674 163.367
R1074 B.n676 B.n675 163.367
R1075 B.n676 B.n29 163.367
R1076 B.n680 B.n29 163.367
R1077 B.n681 B.n680 163.367
R1078 B.n682 B.n681 163.367
R1079 B.n682 B.n27 163.367
R1080 B.n686 B.n27 163.367
R1081 B.n687 B.n686 163.367
R1082 B.n688 B.n687 163.367
R1083 B.n688 B.n25 163.367
R1084 B.n692 B.n25 163.367
R1085 B.n693 B.n692 163.367
R1086 B.n694 B.n693 163.367
R1087 B.n694 B.n23 163.367
R1088 B.n698 B.n23 163.367
R1089 B.n699 B.n698 163.367
R1090 B.n700 B.n699 163.367
R1091 B.n700 B.n21 163.367
R1092 B.n704 B.n21 163.367
R1093 B.n705 B.n704 163.367
R1094 B.n706 B.n705 163.367
R1095 B.n706 B.n19 163.367
R1096 B.n710 B.n19 163.367
R1097 B.n711 B.n710 163.367
R1098 B.n712 B.n711 163.367
R1099 B.n712 B.n17 163.367
R1100 B.n716 B.n17 163.367
R1101 B.n717 B.n716 163.367
R1102 B.n718 B.n717 163.367
R1103 B.n718 B.n15 163.367
R1104 B.n722 B.n15 163.367
R1105 B.n723 B.n722 163.367
R1106 B.n724 B.n723 163.367
R1107 B.n724 B.n13 163.367
R1108 B.n728 B.n13 163.367
R1109 B.n729 B.n728 163.367
R1110 B.n730 B.n729 163.367
R1111 B.n730 B.n11 163.367
R1112 B.n734 B.n11 163.367
R1113 B.n735 B.n734 163.367
R1114 B.n736 B.n735 163.367
R1115 B.n736 B.n9 163.367
R1116 B.n740 B.n9 163.367
R1117 B.n741 B.n740 163.367
R1118 B.n742 B.n741 163.367
R1119 B.n742 B.n7 163.367
R1120 B.n746 B.n7 163.367
R1121 B.n747 B.n746 163.367
R1122 B.n748 B.n747 163.367
R1123 B.n748 B.n5 163.367
R1124 B.n752 B.n5 163.367
R1125 B.n753 B.n752 163.367
R1126 B.n754 B.n753 163.367
R1127 B.n754 B.n3 163.367
R1128 B.n758 B.n3 163.367
R1129 B.n759 B.n758 163.367
R1130 B.n196 B.n2 163.367
R1131 B.n197 B.n196 163.367
R1132 B.n198 B.n197 163.367
R1133 B.n198 B.n193 163.367
R1134 B.n202 B.n193 163.367
R1135 B.n203 B.n202 163.367
R1136 B.n204 B.n203 163.367
R1137 B.n204 B.n191 163.367
R1138 B.n208 B.n191 163.367
R1139 B.n209 B.n208 163.367
R1140 B.n210 B.n209 163.367
R1141 B.n210 B.n189 163.367
R1142 B.n214 B.n189 163.367
R1143 B.n215 B.n214 163.367
R1144 B.n216 B.n215 163.367
R1145 B.n216 B.n187 163.367
R1146 B.n220 B.n187 163.367
R1147 B.n221 B.n220 163.367
R1148 B.n222 B.n221 163.367
R1149 B.n222 B.n185 163.367
R1150 B.n226 B.n185 163.367
R1151 B.n227 B.n226 163.367
R1152 B.n228 B.n227 163.367
R1153 B.n228 B.n183 163.367
R1154 B.n232 B.n183 163.367
R1155 B.n233 B.n232 163.367
R1156 B.n234 B.n233 163.367
R1157 B.n234 B.n181 163.367
R1158 B.n238 B.n181 163.367
R1159 B.n239 B.n238 163.367
R1160 B.n240 B.n239 163.367
R1161 B.n240 B.n179 163.367
R1162 B.n244 B.n179 163.367
R1163 B.n245 B.n244 163.367
R1164 B.n246 B.n245 163.367
R1165 B.n246 B.n177 163.367
R1166 B.n250 B.n177 163.367
R1167 B.n251 B.n250 163.367
R1168 B.n252 B.n251 163.367
R1169 B.n252 B.n175 163.367
R1170 B.n256 B.n175 163.367
R1171 B.n257 B.n256 163.367
R1172 B.n258 B.n257 163.367
R1173 B.n258 B.n173 163.367
R1174 B.n262 B.n173 163.367
R1175 B.n263 B.n262 163.367
R1176 B.n264 B.n263 163.367
R1177 B.n264 B.n171 163.367
R1178 B.n268 B.n171 163.367
R1179 B.n269 B.n268 163.367
R1180 B.n270 B.n269 163.367
R1181 B.n270 B.n169 163.367
R1182 B.n274 B.n169 163.367
R1183 B.n275 B.n274 163.367
R1184 B.n276 B.n275 163.367
R1185 B.n276 B.n167 163.367
R1186 B.n280 B.n167 163.367
R1187 B.n281 B.n280 163.367
R1188 B.n282 B.n281 163.367
R1189 B.n282 B.n165 163.367
R1190 B.n286 B.n165 163.367
R1191 B.n287 B.n286 163.367
R1192 B.n288 B.n287 163.367
R1193 B.n288 B.n163 163.367
R1194 B.n292 B.n163 163.367
R1195 B.n293 B.n292 163.367
R1196 B.n294 B.n293 163.367
R1197 B.n294 B.n161 163.367
R1198 B.n298 B.n161 163.367
R1199 B.n299 B.n298 163.367
R1200 B.n300 B.n299 163.367
R1201 B.n300 B.n159 163.367
R1202 B.n304 B.n159 163.367
R1203 B.n305 B.n304 163.367
R1204 B.n306 B.n305 163.367
R1205 B.n306 B.n157 163.367
R1206 B.n310 B.n157 163.367
R1207 B.n311 B.n310 163.367
R1208 B.n151 B.n150 78.352
R1209 B.n341 B.n340 78.352
R1210 B.n55 B.n54 78.352
R1211 B.n47 B.n46 78.352
R1212 B.n326 B.n151 59.5399
R1213 B.n342 B.n341 59.5399
R1214 B.n612 B.n55 59.5399
R1215 B.n48 B.n47 59.5399
R1216 B.n642 B.n641 30.4395
R1217 B.n599 B.n60 30.4395
R1218 B.n359 B.n140 30.4395
R1219 B.n313 B.n156 30.4395
R1220 B B.n761 18.0485
R1221 B.n643 B.n642 10.6151
R1222 B.n643 B.n40 10.6151
R1223 B.n647 B.n40 10.6151
R1224 B.n648 B.n647 10.6151
R1225 B.n649 B.n648 10.6151
R1226 B.n649 B.n38 10.6151
R1227 B.n653 B.n38 10.6151
R1228 B.n654 B.n653 10.6151
R1229 B.n655 B.n654 10.6151
R1230 B.n655 B.n36 10.6151
R1231 B.n659 B.n36 10.6151
R1232 B.n660 B.n659 10.6151
R1233 B.n661 B.n660 10.6151
R1234 B.n661 B.n34 10.6151
R1235 B.n665 B.n34 10.6151
R1236 B.n666 B.n665 10.6151
R1237 B.n667 B.n666 10.6151
R1238 B.n667 B.n32 10.6151
R1239 B.n671 B.n32 10.6151
R1240 B.n672 B.n671 10.6151
R1241 B.n673 B.n672 10.6151
R1242 B.n673 B.n30 10.6151
R1243 B.n677 B.n30 10.6151
R1244 B.n678 B.n677 10.6151
R1245 B.n679 B.n678 10.6151
R1246 B.n679 B.n28 10.6151
R1247 B.n683 B.n28 10.6151
R1248 B.n684 B.n683 10.6151
R1249 B.n685 B.n684 10.6151
R1250 B.n685 B.n26 10.6151
R1251 B.n689 B.n26 10.6151
R1252 B.n690 B.n689 10.6151
R1253 B.n691 B.n690 10.6151
R1254 B.n691 B.n24 10.6151
R1255 B.n695 B.n24 10.6151
R1256 B.n696 B.n695 10.6151
R1257 B.n697 B.n696 10.6151
R1258 B.n697 B.n22 10.6151
R1259 B.n701 B.n22 10.6151
R1260 B.n702 B.n701 10.6151
R1261 B.n703 B.n702 10.6151
R1262 B.n703 B.n20 10.6151
R1263 B.n707 B.n20 10.6151
R1264 B.n708 B.n707 10.6151
R1265 B.n709 B.n708 10.6151
R1266 B.n709 B.n18 10.6151
R1267 B.n713 B.n18 10.6151
R1268 B.n714 B.n713 10.6151
R1269 B.n715 B.n714 10.6151
R1270 B.n715 B.n16 10.6151
R1271 B.n719 B.n16 10.6151
R1272 B.n720 B.n719 10.6151
R1273 B.n721 B.n720 10.6151
R1274 B.n721 B.n14 10.6151
R1275 B.n725 B.n14 10.6151
R1276 B.n726 B.n725 10.6151
R1277 B.n727 B.n726 10.6151
R1278 B.n727 B.n12 10.6151
R1279 B.n731 B.n12 10.6151
R1280 B.n732 B.n731 10.6151
R1281 B.n733 B.n732 10.6151
R1282 B.n733 B.n10 10.6151
R1283 B.n737 B.n10 10.6151
R1284 B.n738 B.n737 10.6151
R1285 B.n739 B.n738 10.6151
R1286 B.n739 B.n8 10.6151
R1287 B.n743 B.n8 10.6151
R1288 B.n744 B.n743 10.6151
R1289 B.n745 B.n744 10.6151
R1290 B.n745 B.n6 10.6151
R1291 B.n749 B.n6 10.6151
R1292 B.n750 B.n749 10.6151
R1293 B.n751 B.n750 10.6151
R1294 B.n751 B.n4 10.6151
R1295 B.n755 B.n4 10.6151
R1296 B.n756 B.n755 10.6151
R1297 B.n757 B.n756 10.6151
R1298 B.n757 B.n0 10.6151
R1299 B.n641 B.n42 10.6151
R1300 B.n637 B.n42 10.6151
R1301 B.n637 B.n636 10.6151
R1302 B.n636 B.n635 10.6151
R1303 B.n635 B.n44 10.6151
R1304 B.n631 B.n44 10.6151
R1305 B.n631 B.n630 10.6151
R1306 B.n630 B.n629 10.6151
R1307 B.n626 B.n625 10.6151
R1308 B.n625 B.n624 10.6151
R1309 B.n624 B.n50 10.6151
R1310 B.n620 B.n50 10.6151
R1311 B.n620 B.n619 10.6151
R1312 B.n619 B.n618 10.6151
R1313 B.n618 B.n52 10.6151
R1314 B.n614 B.n52 10.6151
R1315 B.n614 B.n613 10.6151
R1316 B.n611 B.n56 10.6151
R1317 B.n607 B.n56 10.6151
R1318 B.n607 B.n606 10.6151
R1319 B.n606 B.n605 10.6151
R1320 B.n605 B.n58 10.6151
R1321 B.n601 B.n58 10.6151
R1322 B.n601 B.n600 10.6151
R1323 B.n600 B.n599 10.6151
R1324 B.n595 B.n60 10.6151
R1325 B.n595 B.n594 10.6151
R1326 B.n594 B.n593 10.6151
R1327 B.n593 B.n62 10.6151
R1328 B.n589 B.n62 10.6151
R1329 B.n589 B.n588 10.6151
R1330 B.n588 B.n587 10.6151
R1331 B.n587 B.n64 10.6151
R1332 B.n583 B.n64 10.6151
R1333 B.n583 B.n582 10.6151
R1334 B.n582 B.n581 10.6151
R1335 B.n581 B.n66 10.6151
R1336 B.n577 B.n66 10.6151
R1337 B.n577 B.n576 10.6151
R1338 B.n576 B.n575 10.6151
R1339 B.n575 B.n68 10.6151
R1340 B.n571 B.n68 10.6151
R1341 B.n571 B.n570 10.6151
R1342 B.n570 B.n569 10.6151
R1343 B.n569 B.n70 10.6151
R1344 B.n565 B.n70 10.6151
R1345 B.n565 B.n564 10.6151
R1346 B.n564 B.n563 10.6151
R1347 B.n563 B.n72 10.6151
R1348 B.n559 B.n72 10.6151
R1349 B.n559 B.n558 10.6151
R1350 B.n558 B.n557 10.6151
R1351 B.n557 B.n74 10.6151
R1352 B.n553 B.n74 10.6151
R1353 B.n553 B.n552 10.6151
R1354 B.n552 B.n551 10.6151
R1355 B.n551 B.n76 10.6151
R1356 B.n547 B.n76 10.6151
R1357 B.n547 B.n546 10.6151
R1358 B.n546 B.n545 10.6151
R1359 B.n545 B.n78 10.6151
R1360 B.n541 B.n78 10.6151
R1361 B.n541 B.n540 10.6151
R1362 B.n540 B.n539 10.6151
R1363 B.n539 B.n80 10.6151
R1364 B.n535 B.n80 10.6151
R1365 B.n535 B.n534 10.6151
R1366 B.n534 B.n533 10.6151
R1367 B.n533 B.n82 10.6151
R1368 B.n529 B.n82 10.6151
R1369 B.n529 B.n528 10.6151
R1370 B.n528 B.n527 10.6151
R1371 B.n527 B.n84 10.6151
R1372 B.n523 B.n84 10.6151
R1373 B.n523 B.n522 10.6151
R1374 B.n522 B.n521 10.6151
R1375 B.n521 B.n86 10.6151
R1376 B.n517 B.n86 10.6151
R1377 B.n517 B.n516 10.6151
R1378 B.n516 B.n515 10.6151
R1379 B.n515 B.n88 10.6151
R1380 B.n511 B.n88 10.6151
R1381 B.n511 B.n510 10.6151
R1382 B.n510 B.n509 10.6151
R1383 B.n509 B.n90 10.6151
R1384 B.n505 B.n90 10.6151
R1385 B.n505 B.n504 10.6151
R1386 B.n504 B.n503 10.6151
R1387 B.n503 B.n92 10.6151
R1388 B.n499 B.n92 10.6151
R1389 B.n499 B.n498 10.6151
R1390 B.n498 B.n497 10.6151
R1391 B.n497 B.n94 10.6151
R1392 B.n493 B.n94 10.6151
R1393 B.n493 B.n492 10.6151
R1394 B.n492 B.n491 10.6151
R1395 B.n491 B.n96 10.6151
R1396 B.n487 B.n96 10.6151
R1397 B.n487 B.n486 10.6151
R1398 B.n486 B.n485 10.6151
R1399 B.n485 B.n98 10.6151
R1400 B.n481 B.n98 10.6151
R1401 B.n481 B.n480 10.6151
R1402 B.n480 B.n479 10.6151
R1403 B.n479 B.n100 10.6151
R1404 B.n475 B.n100 10.6151
R1405 B.n475 B.n474 10.6151
R1406 B.n474 B.n473 10.6151
R1407 B.n473 B.n102 10.6151
R1408 B.n469 B.n102 10.6151
R1409 B.n469 B.n468 10.6151
R1410 B.n468 B.n467 10.6151
R1411 B.n467 B.n104 10.6151
R1412 B.n463 B.n104 10.6151
R1413 B.n463 B.n462 10.6151
R1414 B.n462 B.n461 10.6151
R1415 B.n461 B.n106 10.6151
R1416 B.n457 B.n106 10.6151
R1417 B.n457 B.n456 10.6151
R1418 B.n456 B.n455 10.6151
R1419 B.n455 B.n108 10.6151
R1420 B.n451 B.n108 10.6151
R1421 B.n451 B.n450 10.6151
R1422 B.n450 B.n449 10.6151
R1423 B.n449 B.n110 10.6151
R1424 B.n445 B.n110 10.6151
R1425 B.n445 B.n444 10.6151
R1426 B.n444 B.n443 10.6151
R1427 B.n443 B.n112 10.6151
R1428 B.n439 B.n112 10.6151
R1429 B.n439 B.n438 10.6151
R1430 B.n438 B.n437 10.6151
R1431 B.n437 B.n114 10.6151
R1432 B.n433 B.n114 10.6151
R1433 B.n433 B.n432 10.6151
R1434 B.n432 B.n431 10.6151
R1435 B.n431 B.n116 10.6151
R1436 B.n427 B.n116 10.6151
R1437 B.n427 B.n426 10.6151
R1438 B.n426 B.n425 10.6151
R1439 B.n425 B.n118 10.6151
R1440 B.n421 B.n118 10.6151
R1441 B.n421 B.n420 10.6151
R1442 B.n420 B.n419 10.6151
R1443 B.n419 B.n120 10.6151
R1444 B.n415 B.n120 10.6151
R1445 B.n415 B.n414 10.6151
R1446 B.n414 B.n413 10.6151
R1447 B.n413 B.n122 10.6151
R1448 B.n409 B.n122 10.6151
R1449 B.n409 B.n408 10.6151
R1450 B.n408 B.n407 10.6151
R1451 B.n407 B.n124 10.6151
R1452 B.n403 B.n124 10.6151
R1453 B.n403 B.n402 10.6151
R1454 B.n402 B.n401 10.6151
R1455 B.n401 B.n126 10.6151
R1456 B.n397 B.n126 10.6151
R1457 B.n397 B.n396 10.6151
R1458 B.n396 B.n395 10.6151
R1459 B.n395 B.n128 10.6151
R1460 B.n391 B.n128 10.6151
R1461 B.n391 B.n390 10.6151
R1462 B.n390 B.n389 10.6151
R1463 B.n389 B.n130 10.6151
R1464 B.n385 B.n130 10.6151
R1465 B.n385 B.n384 10.6151
R1466 B.n384 B.n383 10.6151
R1467 B.n383 B.n132 10.6151
R1468 B.n379 B.n132 10.6151
R1469 B.n379 B.n378 10.6151
R1470 B.n378 B.n377 10.6151
R1471 B.n377 B.n134 10.6151
R1472 B.n373 B.n134 10.6151
R1473 B.n373 B.n372 10.6151
R1474 B.n372 B.n371 10.6151
R1475 B.n371 B.n136 10.6151
R1476 B.n367 B.n136 10.6151
R1477 B.n367 B.n366 10.6151
R1478 B.n366 B.n365 10.6151
R1479 B.n365 B.n138 10.6151
R1480 B.n361 B.n138 10.6151
R1481 B.n361 B.n360 10.6151
R1482 B.n360 B.n359 10.6151
R1483 B.n195 B.n1 10.6151
R1484 B.n195 B.n194 10.6151
R1485 B.n199 B.n194 10.6151
R1486 B.n200 B.n199 10.6151
R1487 B.n201 B.n200 10.6151
R1488 B.n201 B.n192 10.6151
R1489 B.n205 B.n192 10.6151
R1490 B.n206 B.n205 10.6151
R1491 B.n207 B.n206 10.6151
R1492 B.n207 B.n190 10.6151
R1493 B.n211 B.n190 10.6151
R1494 B.n212 B.n211 10.6151
R1495 B.n213 B.n212 10.6151
R1496 B.n213 B.n188 10.6151
R1497 B.n217 B.n188 10.6151
R1498 B.n218 B.n217 10.6151
R1499 B.n219 B.n218 10.6151
R1500 B.n219 B.n186 10.6151
R1501 B.n223 B.n186 10.6151
R1502 B.n224 B.n223 10.6151
R1503 B.n225 B.n224 10.6151
R1504 B.n225 B.n184 10.6151
R1505 B.n229 B.n184 10.6151
R1506 B.n230 B.n229 10.6151
R1507 B.n231 B.n230 10.6151
R1508 B.n231 B.n182 10.6151
R1509 B.n235 B.n182 10.6151
R1510 B.n236 B.n235 10.6151
R1511 B.n237 B.n236 10.6151
R1512 B.n237 B.n180 10.6151
R1513 B.n241 B.n180 10.6151
R1514 B.n242 B.n241 10.6151
R1515 B.n243 B.n242 10.6151
R1516 B.n243 B.n178 10.6151
R1517 B.n247 B.n178 10.6151
R1518 B.n248 B.n247 10.6151
R1519 B.n249 B.n248 10.6151
R1520 B.n249 B.n176 10.6151
R1521 B.n253 B.n176 10.6151
R1522 B.n254 B.n253 10.6151
R1523 B.n255 B.n254 10.6151
R1524 B.n255 B.n174 10.6151
R1525 B.n259 B.n174 10.6151
R1526 B.n260 B.n259 10.6151
R1527 B.n261 B.n260 10.6151
R1528 B.n261 B.n172 10.6151
R1529 B.n265 B.n172 10.6151
R1530 B.n266 B.n265 10.6151
R1531 B.n267 B.n266 10.6151
R1532 B.n267 B.n170 10.6151
R1533 B.n271 B.n170 10.6151
R1534 B.n272 B.n271 10.6151
R1535 B.n273 B.n272 10.6151
R1536 B.n273 B.n168 10.6151
R1537 B.n277 B.n168 10.6151
R1538 B.n278 B.n277 10.6151
R1539 B.n279 B.n278 10.6151
R1540 B.n279 B.n166 10.6151
R1541 B.n283 B.n166 10.6151
R1542 B.n284 B.n283 10.6151
R1543 B.n285 B.n284 10.6151
R1544 B.n285 B.n164 10.6151
R1545 B.n289 B.n164 10.6151
R1546 B.n290 B.n289 10.6151
R1547 B.n291 B.n290 10.6151
R1548 B.n291 B.n162 10.6151
R1549 B.n295 B.n162 10.6151
R1550 B.n296 B.n295 10.6151
R1551 B.n297 B.n296 10.6151
R1552 B.n297 B.n160 10.6151
R1553 B.n301 B.n160 10.6151
R1554 B.n302 B.n301 10.6151
R1555 B.n303 B.n302 10.6151
R1556 B.n303 B.n158 10.6151
R1557 B.n307 B.n158 10.6151
R1558 B.n308 B.n307 10.6151
R1559 B.n309 B.n308 10.6151
R1560 B.n309 B.n156 10.6151
R1561 B.n314 B.n313 10.6151
R1562 B.n315 B.n314 10.6151
R1563 B.n315 B.n154 10.6151
R1564 B.n319 B.n154 10.6151
R1565 B.n320 B.n319 10.6151
R1566 B.n321 B.n320 10.6151
R1567 B.n321 B.n152 10.6151
R1568 B.n325 B.n152 10.6151
R1569 B.n328 B.n327 10.6151
R1570 B.n328 B.n148 10.6151
R1571 B.n332 B.n148 10.6151
R1572 B.n333 B.n332 10.6151
R1573 B.n334 B.n333 10.6151
R1574 B.n334 B.n146 10.6151
R1575 B.n338 B.n146 10.6151
R1576 B.n339 B.n338 10.6151
R1577 B.n343 B.n339 10.6151
R1578 B.n347 B.n144 10.6151
R1579 B.n348 B.n347 10.6151
R1580 B.n349 B.n348 10.6151
R1581 B.n349 B.n142 10.6151
R1582 B.n353 B.n142 10.6151
R1583 B.n354 B.n353 10.6151
R1584 B.n355 B.n354 10.6151
R1585 B.n355 B.n140 10.6151
R1586 B.n629 B.n48 9.36635
R1587 B.n612 B.n611 9.36635
R1588 B.n326 B.n325 9.36635
R1589 B.n342 B.n144 9.36635
R1590 B.n761 B.n0 8.11757
R1591 B.n761 B.n1 8.11757
R1592 B.n626 B.n48 1.24928
R1593 B.n613 B.n612 1.24928
R1594 B.n327 B.n326 1.24928
R1595 B.n343 B.n342 1.24928
C0 w_n5818_n1158# VTAIL 1.79422f
C1 VDD2 VP 0.734958f
C2 B VDD2 2.18151f
C3 VDD1 VDD2 2.89477f
C4 VDD2 VN 1.42249f
C5 B VP 2.69187f
C6 VDD2 w_n5818_n1158# 2.64028f
C7 VDD1 VP 1.98777f
C8 VP VN 7.9998f
C9 VDD1 B 2.01952f
C10 VDD2 VTAIL 6.67888f
C11 B VN 1.40753f
C12 VDD1 VN 0.163639f
C13 VP w_n5818_n1158# 13.4349f
C14 B w_n5818_n1158# 9.471709f
C15 VDD1 w_n5818_n1158# 2.44014f
C16 VP VTAIL 3.68727f
C17 w_n5818_n1158# VN 12.682f
C18 B VTAIL 1.29644f
C19 VDD1 VTAIL 6.61783f
C20 VTAIL VN 3.67313f
C21 VDD2 VSUBS 2.381571f
C22 VDD1 VSUBS 2.201568f
C23 VTAIL VSUBS 0.71901f
C24 VN VSUBS 10.33607f
C25 VP VSUBS 4.887106f
C26 B VSUBS 5.437582f
C27 w_n5818_n1158# VSUBS 86.9209f
C28 B.n0 VSUBS 0.014824f
C29 B.n1 VSUBS 0.014824f
C30 B.n2 VSUBS 0.021924f
C31 B.n3 VSUBS 0.016801f
C32 B.n4 VSUBS 0.016801f
C33 B.n5 VSUBS 0.016801f
C34 B.n6 VSUBS 0.016801f
C35 B.n7 VSUBS 0.016801f
C36 B.n8 VSUBS 0.016801f
C37 B.n9 VSUBS 0.016801f
C38 B.n10 VSUBS 0.016801f
C39 B.n11 VSUBS 0.016801f
C40 B.n12 VSUBS 0.016801f
C41 B.n13 VSUBS 0.016801f
C42 B.n14 VSUBS 0.016801f
C43 B.n15 VSUBS 0.016801f
C44 B.n16 VSUBS 0.016801f
C45 B.n17 VSUBS 0.016801f
C46 B.n18 VSUBS 0.016801f
C47 B.n19 VSUBS 0.016801f
C48 B.n20 VSUBS 0.016801f
C49 B.n21 VSUBS 0.016801f
C50 B.n22 VSUBS 0.016801f
C51 B.n23 VSUBS 0.016801f
C52 B.n24 VSUBS 0.016801f
C53 B.n25 VSUBS 0.016801f
C54 B.n26 VSUBS 0.016801f
C55 B.n27 VSUBS 0.016801f
C56 B.n28 VSUBS 0.016801f
C57 B.n29 VSUBS 0.016801f
C58 B.n30 VSUBS 0.016801f
C59 B.n31 VSUBS 0.016801f
C60 B.n32 VSUBS 0.016801f
C61 B.n33 VSUBS 0.016801f
C62 B.n34 VSUBS 0.016801f
C63 B.n35 VSUBS 0.016801f
C64 B.n36 VSUBS 0.016801f
C65 B.n37 VSUBS 0.016801f
C66 B.n38 VSUBS 0.016801f
C67 B.n39 VSUBS 0.016801f
C68 B.n40 VSUBS 0.016801f
C69 B.n41 VSUBS 0.036541f
C70 B.n42 VSUBS 0.016801f
C71 B.n43 VSUBS 0.016801f
C72 B.n44 VSUBS 0.016801f
C73 B.n45 VSUBS 0.016801f
C74 B.t4 VSUBS 0.044239f
C75 B.t5 VSUBS 0.054482f
C76 B.t3 VSUBS 0.425138f
C77 B.n46 VSUBS 0.177729f
C78 B.n47 VSUBS 0.118834f
C79 B.n48 VSUBS 0.038925f
C80 B.n49 VSUBS 0.016801f
C81 B.n50 VSUBS 0.016801f
C82 B.n51 VSUBS 0.016801f
C83 B.n52 VSUBS 0.016801f
C84 B.n53 VSUBS 0.016801f
C85 B.t1 VSUBS 0.044239f
C86 B.t2 VSUBS 0.054482f
C87 B.t0 VSUBS 0.425138f
C88 B.n54 VSUBS 0.177729f
C89 B.n55 VSUBS 0.118834f
C90 B.n56 VSUBS 0.016801f
C91 B.n57 VSUBS 0.016801f
C92 B.n58 VSUBS 0.016801f
C93 B.n59 VSUBS 0.016801f
C94 B.n60 VSUBS 0.036541f
C95 B.n61 VSUBS 0.016801f
C96 B.n62 VSUBS 0.016801f
C97 B.n63 VSUBS 0.016801f
C98 B.n64 VSUBS 0.016801f
C99 B.n65 VSUBS 0.016801f
C100 B.n66 VSUBS 0.016801f
C101 B.n67 VSUBS 0.016801f
C102 B.n68 VSUBS 0.016801f
C103 B.n69 VSUBS 0.016801f
C104 B.n70 VSUBS 0.016801f
C105 B.n71 VSUBS 0.016801f
C106 B.n72 VSUBS 0.016801f
C107 B.n73 VSUBS 0.016801f
C108 B.n74 VSUBS 0.016801f
C109 B.n75 VSUBS 0.016801f
C110 B.n76 VSUBS 0.016801f
C111 B.n77 VSUBS 0.016801f
C112 B.n78 VSUBS 0.016801f
C113 B.n79 VSUBS 0.016801f
C114 B.n80 VSUBS 0.016801f
C115 B.n81 VSUBS 0.016801f
C116 B.n82 VSUBS 0.016801f
C117 B.n83 VSUBS 0.016801f
C118 B.n84 VSUBS 0.016801f
C119 B.n85 VSUBS 0.016801f
C120 B.n86 VSUBS 0.016801f
C121 B.n87 VSUBS 0.016801f
C122 B.n88 VSUBS 0.016801f
C123 B.n89 VSUBS 0.016801f
C124 B.n90 VSUBS 0.016801f
C125 B.n91 VSUBS 0.016801f
C126 B.n92 VSUBS 0.016801f
C127 B.n93 VSUBS 0.016801f
C128 B.n94 VSUBS 0.016801f
C129 B.n95 VSUBS 0.016801f
C130 B.n96 VSUBS 0.016801f
C131 B.n97 VSUBS 0.016801f
C132 B.n98 VSUBS 0.016801f
C133 B.n99 VSUBS 0.016801f
C134 B.n100 VSUBS 0.016801f
C135 B.n101 VSUBS 0.016801f
C136 B.n102 VSUBS 0.016801f
C137 B.n103 VSUBS 0.016801f
C138 B.n104 VSUBS 0.016801f
C139 B.n105 VSUBS 0.016801f
C140 B.n106 VSUBS 0.016801f
C141 B.n107 VSUBS 0.016801f
C142 B.n108 VSUBS 0.016801f
C143 B.n109 VSUBS 0.016801f
C144 B.n110 VSUBS 0.016801f
C145 B.n111 VSUBS 0.016801f
C146 B.n112 VSUBS 0.016801f
C147 B.n113 VSUBS 0.016801f
C148 B.n114 VSUBS 0.016801f
C149 B.n115 VSUBS 0.016801f
C150 B.n116 VSUBS 0.016801f
C151 B.n117 VSUBS 0.016801f
C152 B.n118 VSUBS 0.016801f
C153 B.n119 VSUBS 0.016801f
C154 B.n120 VSUBS 0.016801f
C155 B.n121 VSUBS 0.016801f
C156 B.n122 VSUBS 0.016801f
C157 B.n123 VSUBS 0.016801f
C158 B.n124 VSUBS 0.016801f
C159 B.n125 VSUBS 0.016801f
C160 B.n126 VSUBS 0.016801f
C161 B.n127 VSUBS 0.016801f
C162 B.n128 VSUBS 0.016801f
C163 B.n129 VSUBS 0.016801f
C164 B.n130 VSUBS 0.016801f
C165 B.n131 VSUBS 0.016801f
C166 B.n132 VSUBS 0.016801f
C167 B.n133 VSUBS 0.016801f
C168 B.n134 VSUBS 0.016801f
C169 B.n135 VSUBS 0.016801f
C170 B.n136 VSUBS 0.016801f
C171 B.n137 VSUBS 0.016801f
C172 B.n138 VSUBS 0.016801f
C173 B.n139 VSUBS 0.016801f
C174 B.n140 VSUBS 0.036437f
C175 B.n141 VSUBS 0.016801f
C176 B.n142 VSUBS 0.016801f
C177 B.n143 VSUBS 0.016801f
C178 B.n144 VSUBS 0.015812f
C179 B.n145 VSUBS 0.016801f
C180 B.n146 VSUBS 0.016801f
C181 B.n147 VSUBS 0.016801f
C182 B.n148 VSUBS 0.016801f
C183 B.n149 VSUBS 0.016801f
C184 B.t8 VSUBS 0.044239f
C185 B.t7 VSUBS 0.054482f
C186 B.t6 VSUBS 0.425138f
C187 B.n150 VSUBS 0.177729f
C188 B.n151 VSUBS 0.118834f
C189 B.n152 VSUBS 0.016801f
C190 B.n153 VSUBS 0.016801f
C191 B.n154 VSUBS 0.016801f
C192 B.n155 VSUBS 0.016801f
C193 B.n156 VSUBS 0.036541f
C194 B.n157 VSUBS 0.016801f
C195 B.n158 VSUBS 0.016801f
C196 B.n159 VSUBS 0.016801f
C197 B.n160 VSUBS 0.016801f
C198 B.n161 VSUBS 0.016801f
C199 B.n162 VSUBS 0.016801f
C200 B.n163 VSUBS 0.016801f
C201 B.n164 VSUBS 0.016801f
C202 B.n165 VSUBS 0.016801f
C203 B.n166 VSUBS 0.016801f
C204 B.n167 VSUBS 0.016801f
C205 B.n168 VSUBS 0.016801f
C206 B.n169 VSUBS 0.016801f
C207 B.n170 VSUBS 0.016801f
C208 B.n171 VSUBS 0.016801f
C209 B.n172 VSUBS 0.016801f
C210 B.n173 VSUBS 0.016801f
C211 B.n174 VSUBS 0.016801f
C212 B.n175 VSUBS 0.016801f
C213 B.n176 VSUBS 0.016801f
C214 B.n177 VSUBS 0.016801f
C215 B.n178 VSUBS 0.016801f
C216 B.n179 VSUBS 0.016801f
C217 B.n180 VSUBS 0.016801f
C218 B.n181 VSUBS 0.016801f
C219 B.n182 VSUBS 0.016801f
C220 B.n183 VSUBS 0.016801f
C221 B.n184 VSUBS 0.016801f
C222 B.n185 VSUBS 0.016801f
C223 B.n186 VSUBS 0.016801f
C224 B.n187 VSUBS 0.016801f
C225 B.n188 VSUBS 0.016801f
C226 B.n189 VSUBS 0.016801f
C227 B.n190 VSUBS 0.016801f
C228 B.n191 VSUBS 0.016801f
C229 B.n192 VSUBS 0.016801f
C230 B.n193 VSUBS 0.016801f
C231 B.n194 VSUBS 0.016801f
C232 B.n195 VSUBS 0.016801f
C233 B.n196 VSUBS 0.016801f
C234 B.n197 VSUBS 0.016801f
C235 B.n198 VSUBS 0.016801f
C236 B.n199 VSUBS 0.016801f
C237 B.n200 VSUBS 0.016801f
C238 B.n201 VSUBS 0.016801f
C239 B.n202 VSUBS 0.016801f
C240 B.n203 VSUBS 0.016801f
C241 B.n204 VSUBS 0.016801f
C242 B.n205 VSUBS 0.016801f
C243 B.n206 VSUBS 0.016801f
C244 B.n207 VSUBS 0.016801f
C245 B.n208 VSUBS 0.016801f
C246 B.n209 VSUBS 0.016801f
C247 B.n210 VSUBS 0.016801f
C248 B.n211 VSUBS 0.016801f
C249 B.n212 VSUBS 0.016801f
C250 B.n213 VSUBS 0.016801f
C251 B.n214 VSUBS 0.016801f
C252 B.n215 VSUBS 0.016801f
C253 B.n216 VSUBS 0.016801f
C254 B.n217 VSUBS 0.016801f
C255 B.n218 VSUBS 0.016801f
C256 B.n219 VSUBS 0.016801f
C257 B.n220 VSUBS 0.016801f
C258 B.n221 VSUBS 0.016801f
C259 B.n222 VSUBS 0.016801f
C260 B.n223 VSUBS 0.016801f
C261 B.n224 VSUBS 0.016801f
C262 B.n225 VSUBS 0.016801f
C263 B.n226 VSUBS 0.016801f
C264 B.n227 VSUBS 0.016801f
C265 B.n228 VSUBS 0.016801f
C266 B.n229 VSUBS 0.016801f
C267 B.n230 VSUBS 0.016801f
C268 B.n231 VSUBS 0.016801f
C269 B.n232 VSUBS 0.016801f
C270 B.n233 VSUBS 0.016801f
C271 B.n234 VSUBS 0.016801f
C272 B.n235 VSUBS 0.016801f
C273 B.n236 VSUBS 0.016801f
C274 B.n237 VSUBS 0.016801f
C275 B.n238 VSUBS 0.016801f
C276 B.n239 VSUBS 0.016801f
C277 B.n240 VSUBS 0.016801f
C278 B.n241 VSUBS 0.016801f
C279 B.n242 VSUBS 0.016801f
C280 B.n243 VSUBS 0.016801f
C281 B.n244 VSUBS 0.016801f
C282 B.n245 VSUBS 0.016801f
C283 B.n246 VSUBS 0.016801f
C284 B.n247 VSUBS 0.016801f
C285 B.n248 VSUBS 0.016801f
C286 B.n249 VSUBS 0.016801f
C287 B.n250 VSUBS 0.016801f
C288 B.n251 VSUBS 0.016801f
C289 B.n252 VSUBS 0.016801f
C290 B.n253 VSUBS 0.016801f
C291 B.n254 VSUBS 0.016801f
C292 B.n255 VSUBS 0.016801f
C293 B.n256 VSUBS 0.016801f
C294 B.n257 VSUBS 0.016801f
C295 B.n258 VSUBS 0.016801f
C296 B.n259 VSUBS 0.016801f
C297 B.n260 VSUBS 0.016801f
C298 B.n261 VSUBS 0.016801f
C299 B.n262 VSUBS 0.016801f
C300 B.n263 VSUBS 0.016801f
C301 B.n264 VSUBS 0.016801f
C302 B.n265 VSUBS 0.016801f
C303 B.n266 VSUBS 0.016801f
C304 B.n267 VSUBS 0.016801f
C305 B.n268 VSUBS 0.016801f
C306 B.n269 VSUBS 0.016801f
C307 B.n270 VSUBS 0.016801f
C308 B.n271 VSUBS 0.016801f
C309 B.n272 VSUBS 0.016801f
C310 B.n273 VSUBS 0.016801f
C311 B.n274 VSUBS 0.016801f
C312 B.n275 VSUBS 0.016801f
C313 B.n276 VSUBS 0.016801f
C314 B.n277 VSUBS 0.016801f
C315 B.n278 VSUBS 0.016801f
C316 B.n279 VSUBS 0.016801f
C317 B.n280 VSUBS 0.016801f
C318 B.n281 VSUBS 0.016801f
C319 B.n282 VSUBS 0.016801f
C320 B.n283 VSUBS 0.016801f
C321 B.n284 VSUBS 0.016801f
C322 B.n285 VSUBS 0.016801f
C323 B.n286 VSUBS 0.016801f
C324 B.n287 VSUBS 0.016801f
C325 B.n288 VSUBS 0.016801f
C326 B.n289 VSUBS 0.016801f
C327 B.n290 VSUBS 0.016801f
C328 B.n291 VSUBS 0.016801f
C329 B.n292 VSUBS 0.016801f
C330 B.n293 VSUBS 0.016801f
C331 B.n294 VSUBS 0.016801f
C332 B.n295 VSUBS 0.016801f
C333 B.n296 VSUBS 0.016801f
C334 B.n297 VSUBS 0.016801f
C335 B.n298 VSUBS 0.016801f
C336 B.n299 VSUBS 0.016801f
C337 B.n300 VSUBS 0.016801f
C338 B.n301 VSUBS 0.016801f
C339 B.n302 VSUBS 0.016801f
C340 B.n303 VSUBS 0.016801f
C341 B.n304 VSUBS 0.016801f
C342 B.n305 VSUBS 0.016801f
C343 B.n306 VSUBS 0.016801f
C344 B.n307 VSUBS 0.016801f
C345 B.n308 VSUBS 0.016801f
C346 B.n309 VSUBS 0.016801f
C347 B.n310 VSUBS 0.016801f
C348 B.n311 VSUBS 0.036541f
C349 B.n312 VSUBS 0.038567f
C350 B.n313 VSUBS 0.038567f
C351 B.n314 VSUBS 0.016801f
C352 B.n315 VSUBS 0.016801f
C353 B.n316 VSUBS 0.016801f
C354 B.n317 VSUBS 0.016801f
C355 B.n318 VSUBS 0.016801f
C356 B.n319 VSUBS 0.016801f
C357 B.n320 VSUBS 0.016801f
C358 B.n321 VSUBS 0.016801f
C359 B.n322 VSUBS 0.016801f
C360 B.n323 VSUBS 0.016801f
C361 B.n324 VSUBS 0.016801f
C362 B.n325 VSUBS 0.015812f
C363 B.n326 VSUBS 0.038925f
C364 B.n327 VSUBS 0.009389f
C365 B.n328 VSUBS 0.016801f
C366 B.n329 VSUBS 0.016801f
C367 B.n330 VSUBS 0.016801f
C368 B.n331 VSUBS 0.016801f
C369 B.n332 VSUBS 0.016801f
C370 B.n333 VSUBS 0.016801f
C371 B.n334 VSUBS 0.016801f
C372 B.n335 VSUBS 0.016801f
C373 B.n336 VSUBS 0.016801f
C374 B.n337 VSUBS 0.016801f
C375 B.n338 VSUBS 0.016801f
C376 B.n339 VSUBS 0.016801f
C377 B.t11 VSUBS 0.044239f
C378 B.t10 VSUBS 0.054482f
C379 B.t9 VSUBS 0.425138f
C380 B.n340 VSUBS 0.177729f
C381 B.n341 VSUBS 0.118834f
C382 B.n342 VSUBS 0.038925f
C383 B.n343 VSUBS 0.009389f
C384 B.n344 VSUBS 0.016801f
C385 B.n345 VSUBS 0.016801f
C386 B.n346 VSUBS 0.016801f
C387 B.n347 VSUBS 0.016801f
C388 B.n348 VSUBS 0.016801f
C389 B.n349 VSUBS 0.016801f
C390 B.n350 VSUBS 0.016801f
C391 B.n351 VSUBS 0.016801f
C392 B.n352 VSUBS 0.016801f
C393 B.n353 VSUBS 0.016801f
C394 B.n354 VSUBS 0.016801f
C395 B.n355 VSUBS 0.016801f
C396 B.n356 VSUBS 0.016801f
C397 B.n357 VSUBS 0.038567f
C398 B.n358 VSUBS 0.036541f
C399 B.n359 VSUBS 0.038671f
C400 B.n360 VSUBS 0.016801f
C401 B.n361 VSUBS 0.016801f
C402 B.n362 VSUBS 0.016801f
C403 B.n363 VSUBS 0.016801f
C404 B.n364 VSUBS 0.016801f
C405 B.n365 VSUBS 0.016801f
C406 B.n366 VSUBS 0.016801f
C407 B.n367 VSUBS 0.016801f
C408 B.n368 VSUBS 0.016801f
C409 B.n369 VSUBS 0.016801f
C410 B.n370 VSUBS 0.016801f
C411 B.n371 VSUBS 0.016801f
C412 B.n372 VSUBS 0.016801f
C413 B.n373 VSUBS 0.016801f
C414 B.n374 VSUBS 0.016801f
C415 B.n375 VSUBS 0.016801f
C416 B.n376 VSUBS 0.016801f
C417 B.n377 VSUBS 0.016801f
C418 B.n378 VSUBS 0.016801f
C419 B.n379 VSUBS 0.016801f
C420 B.n380 VSUBS 0.016801f
C421 B.n381 VSUBS 0.016801f
C422 B.n382 VSUBS 0.016801f
C423 B.n383 VSUBS 0.016801f
C424 B.n384 VSUBS 0.016801f
C425 B.n385 VSUBS 0.016801f
C426 B.n386 VSUBS 0.016801f
C427 B.n387 VSUBS 0.016801f
C428 B.n388 VSUBS 0.016801f
C429 B.n389 VSUBS 0.016801f
C430 B.n390 VSUBS 0.016801f
C431 B.n391 VSUBS 0.016801f
C432 B.n392 VSUBS 0.016801f
C433 B.n393 VSUBS 0.016801f
C434 B.n394 VSUBS 0.016801f
C435 B.n395 VSUBS 0.016801f
C436 B.n396 VSUBS 0.016801f
C437 B.n397 VSUBS 0.016801f
C438 B.n398 VSUBS 0.016801f
C439 B.n399 VSUBS 0.016801f
C440 B.n400 VSUBS 0.016801f
C441 B.n401 VSUBS 0.016801f
C442 B.n402 VSUBS 0.016801f
C443 B.n403 VSUBS 0.016801f
C444 B.n404 VSUBS 0.016801f
C445 B.n405 VSUBS 0.016801f
C446 B.n406 VSUBS 0.016801f
C447 B.n407 VSUBS 0.016801f
C448 B.n408 VSUBS 0.016801f
C449 B.n409 VSUBS 0.016801f
C450 B.n410 VSUBS 0.016801f
C451 B.n411 VSUBS 0.016801f
C452 B.n412 VSUBS 0.016801f
C453 B.n413 VSUBS 0.016801f
C454 B.n414 VSUBS 0.016801f
C455 B.n415 VSUBS 0.016801f
C456 B.n416 VSUBS 0.016801f
C457 B.n417 VSUBS 0.016801f
C458 B.n418 VSUBS 0.016801f
C459 B.n419 VSUBS 0.016801f
C460 B.n420 VSUBS 0.016801f
C461 B.n421 VSUBS 0.016801f
C462 B.n422 VSUBS 0.016801f
C463 B.n423 VSUBS 0.016801f
C464 B.n424 VSUBS 0.016801f
C465 B.n425 VSUBS 0.016801f
C466 B.n426 VSUBS 0.016801f
C467 B.n427 VSUBS 0.016801f
C468 B.n428 VSUBS 0.016801f
C469 B.n429 VSUBS 0.016801f
C470 B.n430 VSUBS 0.016801f
C471 B.n431 VSUBS 0.016801f
C472 B.n432 VSUBS 0.016801f
C473 B.n433 VSUBS 0.016801f
C474 B.n434 VSUBS 0.016801f
C475 B.n435 VSUBS 0.016801f
C476 B.n436 VSUBS 0.016801f
C477 B.n437 VSUBS 0.016801f
C478 B.n438 VSUBS 0.016801f
C479 B.n439 VSUBS 0.016801f
C480 B.n440 VSUBS 0.016801f
C481 B.n441 VSUBS 0.016801f
C482 B.n442 VSUBS 0.016801f
C483 B.n443 VSUBS 0.016801f
C484 B.n444 VSUBS 0.016801f
C485 B.n445 VSUBS 0.016801f
C486 B.n446 VSUBS 0.016801f
C487 B.n447 VSUBS 0.016801f
C488 B.n448 VSUBS 0.016801f
C489 B.n449 VSUBS 0.016801f
C490 B.n450 VSUBS 0.016801f
C491 B.n451 VSUBS 0.016801f
C492 B.n452 VSUBS 0.016801f
C493 B.n453 VSUBS 0.016801f
C494 B.n454 VSUBS 0.016801f
C495 B.n455 VSUBS 0.016801f
C496 B.n456 VSUBS 0.016801f
C497 B.n457 VSUBS 0.016801f
C498 B.n458 VSUBS 0.016801f
C499 B.n459 VSUBS 0.016801f
C500 B.n460 VSUBS 0.016801f
C501 B.n461 VSUBS 0.016801f
C502 B.n462 VSUBS 0.016801f
C503 B.n463 VSUBS 0.016801f
C504 B.n464 VSUBS 0.016801f
C505 B.n465 VSUBS 0.016801f
C506 B.n466 VSUBS 0.016801f
C507 B.n467 VSUBS 0.016801f
C508 B.n468 VSUBS 0.016801f
C509 B.n469 VSUBS 0.016801f
C510 B.n470 VSUBS 0.016801f
C511 B.n471 VSUBS 0.016801f
C512 B.n472 VSUBS 0.016801f
C513 B.n473 VSUBS 0.016801f
C514 B.n474 VSUBS 0.016801f
C515 B.n475 VSUBS 0.016801f
C516 B.n476 VSUBS 0.016801f
C517 B.n477 VSUBS 0.016801f
C518 B.n478 VSUBS 0.016801f
C519 B.n479 VSUBS 0.016801f
C520 B.n480 VSUBS 0.016801f
C521 B.n481 VSUBS 0.016801f
C522 B.n482 VSUBS 0.016801f
C523 B.n483 VSUBS 0.016801f
C524 B.n484 VSUBS 0.016801f
C525 B.n485 VSUBS 0.016801f
C526 B.n486 VSUBS 0.016801f
C527 B.n487 VSUBS 0.016801f
C528 B.n488 VSUBS 0.016801f
C529 B.n489 VSUBS 0.016801f
C530 B.n490 VSUBS 0.016801f
C531 B.n491 VSUBS 0.016801f
C532 B.n492 VSUBS 0.016801f
C533 B.n493 VSUBS 0.016801f
C534 B.n494 VSUBS 0.016801f
C535 B.n495 VSUBS 0.016801f
C536 B.n496 VSUBS 0.016801f
C537 B.n497 VSUBS 0.016801f
C538 B.n498 VSUBS 0.016801f
C539 B.n499 VSUBS 0.016801f
C540 B.n500 VSUBS 0.016801f
C541 B.n501 VSUBS 0.016801f
C542 B.n502 VSUBS 0.016801f
C543 B.n503 VSUBS 0.016801f
C544 B.n504 VSUBS 0.016801f
C545 B.n505 VSUBS 0.016801f
C546 B.n506 VSUBS 0.016801f
C547 B.n507 VSUBS 0.016801f
C548 B.n508 VSUBS 0.016801f
C549 B.n509 VSUBS 0.016801f
C550 B.n510 VSUBS 0.016801f
C551 B.n511 VSUBS 0.016801f
C552 B.n512 VSUBS 0.016801f
C553 B.n513 VSUBS 0.016801f
C554 B.n514 VSUBS 0.016801f
C555 B.n515 VSUBS 0.016801f
C556 B.n516 VSUBS 0.016801f
C557 B.n517 VSUBS 0.016801f
C558 B.n518 VSUBS 0.016801f
C559 B.n519 VSUBS 0.016801f
C560 B.n520 VSUBS 0.016801f
C561 B.n521 VSUBS 0.016801f
C562 B.n522 VSUBS 0.016801f
C563 B.n523 VSUBS 0.016801f
C564 B.n524 VSUBS 0.016801f
C565 B.n525 VSUBS 0.016801f
C566 B.n526 VSUBS 0.016801f
C567 B.n527 VSUBS 0.016801f
C568 B.n528 VSUBS 0.016801f
C569 B.n529 VSUBS 0.016801f
C570 B.n530 VSUBS 0.016801f
C571 B.n531 VSUBS 0.016801f
C572 B.n532 VSUBS 0.016801f
C573 B.n533 VSUBS 0.016801f
C574 B.n534 VSUBS 0.016801f
C575 B.n535 VSUBS 0.016801f
C576 B.n536 VSUBS 0.016801f
C577 B.n537 VSUBS 0.016801f
C578 B.n538 VSUBS 0.016801f
C579 B.n539 VSUBS 0.016801f
C580 B.n540 VSUBS 0.016801f
C581 B.n541 VSUBS 0.016801f
C582 B.n542 VSUBS 0.016801f
C583 B.n543 VSUBS 0.016801f
C584 B.n544 VSUBS 0.016801f
C585 B.n545 VSUBS 0.016801f
C586 B.n546 VSUBS 0.016801f
C587 B.n547 VSUBS 0.016801f
C588 B.n548 VSUBS 0.016801f
C589 B.n549 VSUBS 0.016801f
C590 B.n550 VSUBS 0.016801f
C591 B.n551 VSUBS 0.016801f
C592 B.n552 VSUBS 0.016801f
C593 B.n553 VSUBS 0.016801f
C594 B.n554 VSUBS 0.016801f
C595 B.n555 VSUBS 0.016801f
C596 B.n556 VSUBS 0.016801f
C597 B.n557 VSUBS 0.016801f
C598 B.n558 VSUBS 0.016801f
C599 B.n559 VSUBS 0.016801f
C600 B.n560 VSUBS 0.016801f
C601 B.n561 VSUBS 0.016801f
C602 B.n562 VSUBS 0.016801f
C603 B.n563 VSUBS 0.016801f
C604 B.n564 VSUBS 0.016801f
C605 B.n565 VSUBS 0.016801f
C606 B.n566 VSUBS 0.016801f
C607 B.n567 VSUBS 0.016801f
C608 B.n568 VSUBS 0.016801f
C609 B.n569 VSUBS 0.016801f
C610 B.n570 VSUBS 0.016801f
C611 B.n571 VSUBS 0.016801f
C612 B.n572 VSUBS 0.016801f
C613 B.n573 VSUBS 0.016801f
C614 B.n574 VSUBS 0.016801f
C615 B.n575 VSUBS 0.016801f
C616 B.n576 VSUBS 0.016801f
C617 B.n577 VSUBS 0.016801f
C618 B.n578 VSUBS 0.016801f
C619 B.n579 VSUBS 0.016801f
C620 B.n580 VSUBS 0.016801f
C621 B.n581 VSUBS 0.016801f
C622 B.n582 VSUBS 0.016801f
C623 B.n583 VSUBS 0.016801f
C624 B.n584 VSUBS 0.016801f
C625 B.n585 VSUBS 0.016801f
C626 B.n586 VSUBS 0.016801f
C627 B.n587 VSUBS 0.016801f
C628 B.n588 VSUBS 0.016801f
C629 B.n589 VSUBS 0.016801f
C630 B.n590 VSUBS 0.016801f
C631 B.n591 VSUBS 0.016801f
C632 B.n592 VSUBS 0.016801f
C633 B.n593 VSUBS 0.016801f
C634 B.n594 VSUBS 0.016801f
C635 B.n595 VSUBS 0.016801f
C636 B.n596 VSUBS 0.016801f
C637 B.n597 VSUBS 0.036541f
C638 B.n598 VSUBS 0.038567f
C639 B.n599 VSUBS 0.038567f
C640 B.n600 VSUBS 0.016801f
C641 B.n601 VSUBS 0.016801f
C642 B.n602 VSUBS 0.016801f
C643 B.n603 VSUBS 0.016801f
C644 B.n604 VSUBS 0.016801f
C645 B.n605 VSUBS 0.016801f
C646 B.n606 VSUBS 0.016801f
C647 B.n607 VSUBS 0.016801f
C648 B.n608 VSUBS 0.016801f
C649 B.n609 VSUBS 0.016801f
C650 B.n610 VSUBS 0.016801f
C651 B.n611 VSUBS 0.015812f
C652 B.n612 VSUBS 0.038925f
C653 B.n613 VSUBS 0.009389f
C654 B.n614 VSUBS 0.016801f
C655 B.n615 VSUBS 0.016801f
C656 B.n616 VSUBS 0.016801f
C657 B.n617 VSUBS 0.016801f
C658 B.n618 VSUBS 0.016801f
C659 B.n619 VSUBS 0.016801f
C660 B.n620 VSUBS 0.016801f
C661 B.n621 VSUBS 0.016801f
C662 B.n622 VSUBS 0.016801f
C663 B.n623 VSUBS 0.016801f
C664 B.n624 VSUBS 0.016801f
C665 B.n625 VSUBS 0.016801f
C666 B.n626 VSUBS 0.009389f
C667 B.n627 VSUBS 0.016801f
C668 B.n628 VSUBS 0.016801f
C669 B.n629 VSUBS 0.015812f
C670 B.n630 VSUBS 0.016801f
C671 B.n631 VSUBS 0.016801f
C672 B.n632 VSUBS 0.016801f
C673 B.n633 VSUBS 0.016801f
C674 B.n634 VSUBS 0.016801f
C675 B.n635 VSUBS 0.016801f
C676 B.n636 VSUBS 0.016801f
C677 B.n637 VSUBS 0.016801f
C678 B.n638 VSUBS 0.016801f
C679 B.n639 VSUBS 0.016801f
C680 B.n640 VSUBS 0.038567f
C681 B.n641 VSUBS 0.038567f
C682 B.n642 VSUBS 0.036541f
C683 B.n643 VSUBS 0.016801f
C684 B.n644 VSUBS 0.016801f
C685 B.n645 VSUBS 0.016801f
C686 B.n646 VSUBS 0.016801f
C687 B.n647 VSUBS 0.016801f
C688 B.n648 VSUBS 0.016801f
C689 B.n649 VSUBS 0.016801f
C690 B.n650 VSUBS 0.016801f
C691 B.n651 VSUBS 0.016801f
C692 B.n652 VSUBS 0.016801f
C693 B.n653 VSUBS 0.016801f
C694 B.n654 VSUBS 0.016801f
C695 B.n655 VSUBS 0.016801f
C696 B.n656 VSUBS 0.016801f
C697 B.n657 VSUBS 0.016801f
C698 B.n658 VSUBS 0.016801f
C699 B.n659 VSUBS 0.016801f
C700 B.n660 VSUBS 0.016801f
C701 B.n661 VSUBS 0.016801f
C702 B.n662 VSUBS 0.016801f
C703 B.n663 VSUBS 0.016801f
C704 B.n664 VSUBS 0.016801f
C705 B.n665 VSUBS 0.016801f
C706 B.n666 VSUBS 0.016801f
C707 B.n667 VSUBS 0.016801f
C708 B.n668 VSUBS 0.016801f
C709 B.n669 VSUBS 0.016801f
C710 B.n670 VSUBS 0.016801f
C711 B.n671 VSUBS 0.016801f
C712 B.n672 VSUBS 0.016801f
C713 B.n673 VSUBS 0.016801f
C714 B.n674 VSUBS 0.016801f
C715 B.n675 VSUBS 0.016801f
C716 B.n676 VSUBS 0.016801f
C717 B.n677 VSUBS 0.016801f
C718 B.n678 VSUBS 0.016801f
C719 B.n679 VSUBS 0.016801f
C720 B.n680 VSUBS 0.016801f
C721 B.n681 VSUBS 0.016801f
C722 B.n682 VSUBS 0.016801f
C723 B.n683 VSUBS 0.016801f
C724 B.n684 VSUBS 0.016801f
C725 B.n685 VSUBS 0.016801f
C726 B.n686 VSUBS 0.016801f
C727 B.n687 VSUBS 0.016801f
C728 B.n688 VSUBS 0.016801f
C729 B.n689 VSUBS 0.016801f
C730 B.n690 VSUBS 0.016801f
C731 B.n691 VSUBS 0.016801f
C732 B.n692 VSUBS 0.016801f
C733 B.n693 VSUBS 0.016801f
C734 B.n694 VSUBS 0.016801f
C735 B.n695 VSUBS 0.016801f
C736 B.n696 VSUBS 0.016801f
C737 B.n697 VSUBS 0.016801f
C738 B.n698 VSUBS 0.016801f
C739 B.n699 VSUBS 0.016801f
C740 B.n700 VSUBS 0.016801f
C741 B.n701 VSUBS 0.016801f
C742 B.n702 VSUBS 0.016801f
C743 B.n703 VSUBS 0.016801f
C744 B.n704 VSUBS 0.016801f
C745 B.n705 VSUBS 0.016801f
C746 B.n706 VSUBS 0.016801f
C747 B.n707 VSUBS 0.016801f
C748 B.n708 VSUBS 0.016801f
C749 B.n709 VSUBS 0.016801f
C750 B.n710 VSUBS 0.016801f
C751 B.n711 VSUBS 0.016801f
C752 B.n712 VSUBS 0.016801f
C753 B.n713 VSUBS 0.016801f
C754 B.n714 VSUBS 0.016801f
C755 B.n715 VSUBS 0.016801f
C756 B.n716 VSUBS 0.016801f
C757 B.n717 VSUBS 0.016801f
C758 B.n718 VSUBS 0.016801f
C759 B.n719 VSUBS 0.016801f
C760 B.n720 VSUBS 0.016801f
C761 B.n721 VSUBS 0.016801f
C762 B.n722 VSUBS 0.016801f
C763 B.n723 VSUBS 0.016801f
C764 B.n724 VSUBS 0.016801f
C765 B.n725 VSUBS 0.016801f
C766 B.n726 VSUBS 0.016801f
C767 B.n727 VSUBS 0.016801f
C768 B.n728 VSUBS 0.016801f
C769 B.n729 VSUBS 0.016801f
C770 B.n730 VSUBS 0.016801f
C771 B.n731 VSUBS 0.016801f
C772 B.n732 VSUBS 0.016801f
C773 B.n733 VSUBS 0.016801f
C774 B.n734 VSUBS 0.016801f
C775 B.n735 VSUBS 0.016801f
C776 B.n736 VSUBS 0.016801f
C777 B.n737 VSUBS 0.016801f
C778 B.n738 VSUBS 0.016801f
C779 B.n739 VSUBS 0.016801f
C780 B.n740 VSUBS 0.016801f
C781 B.n741 VSUBS 0.016801f
C782 B.n742 VSUBS 0.016801f
C783 B.n743 VSUBS 0.016801f
C784 B.n744 VSUBS 0.016801f
C785 B.n745 VSUBS 0.016801f
C786 B.n746 VSUBS 0.016801f
C787 B.n747 VSUBS 0.016801f
C788 B.n748 VSUBS 0.016801f
C789 B.n749 VSUBS 0.016801f
C790 B.n750 VSUBS 0.016801f
C791 B.n751 VSUBS 0.016801f
C792 B.n752 VSUBS 0.016801f
C793 B.n753 VSUBS 0.016801f
C794 B.n754 VSUBS 0.016801f
C795 B.n755 VSUBS 0.016801f
C796 B.n756 VSUBS 0.016801f
C797 B.n757 VSUBS 0.016801f
C798 B.n758 VSUBS 0.016801f
C799 B.n759 VSUBS 0.021924f
C800 B.n760 VSUBS 0.023355f
C801 B.n761 VSUBS 0.046443f
C802 VDD2.t5 VSUBS 0.169173f
C803 VDD2.t0 VSUBS 0.031682f
C804 VDD2.t7 VSUBS 0.031682f
C805 VDD2.n0 VSUBS 0.085678f
C806 VDD2.n1 VSUBS 1.7255f
C807 VDD2.t2 VSUBS 0.031682f
C808 VDD2.t8 VSUBS 0.031682f
C809 VDD2.n2 VSUBS 0.090307f
C810 VDD2.n3 VSUBS 4.76378f
C811 VDD2.t9 VSUBS 0.164949f
C812 VDD2.n4 VSUBS 4.41808f
C813 VDD2.t6 VSUBS 0.031682f
C814 VDD2.t1 VSUBS 0.031682f
C815 VDD2.n5 VSUBS 0.085678f
C816 VDD2.n6 VSUBS 0.923073f
C817 VDD2.t3 VSUBS 0.031682f
C818 VDD2.t4 VSUBS 0.031682f
C819 VDD2.n7 VSUBS 0.090299f
C820 VN.t1 VSUBS 0.366143f
C821 VN.n0 VSUBS 0.453197f
C822 VN.n1 VSUBS 0.057106f
C823 VN.n2 VSUBS 0.108907f
C824 VN.n3 VSUBS 0.057106f
C825 VN.n4 VSUBS 0.102229f
C826 VN.n5 VSUBS 0.057106f
C827 VN.n6 VSUBS 0.112213f
C828 VN.n7 VSUBS 0.057106f
C829 VN.n8 VSUBS 0.106432f
C830 VN.n9 VSUBS 0.057106f
C831 VN.t2 VSUBS 0.366143f
C832 VN.n10 VSUBS 0.114491f
C833 VN.n11 VSUBS 0.057106f
C834 VN.n12 VSUBS 0.106432f
C835 VN.t4 VSUBS 0.933614f
C836 VN.n13 VSUBS 0.569694f
C837 VN.t9 VSUBS 0.366143f
C838 VN.n14 VSUBS 0.42325f
C839 VN.n15 VSUBS 0.05809f
C840 VN.n16 VSUBS 0.725776f
C841 VN.n17 VSUBS 0.057106f
C842 VN.n18 VSUBS 0.057106f
C843 VN.n19 VSUBS 0.106432f
C844 VN.n20 VSUBS 0.112213f
C845 VN.n21 VSUBS 0.046459f
C846 VN.n22 VSUBS 0.057106f
C847 VN.n23 VSUBS 0.057106f
C848 VN.n24 VSUBS 0.057106f
C849 VN.n25 VSUBS 0.106432f
C850 VN.n26 VSUBS 0.106432f
C851 VN.n27 VSUBS 0.294452f
C852 VN.n28 VSUBS 0.057106f
C853 VN.n29 VSUBS 0.057106f
C854 VN.n30 VSUBS 0.057106f
C855 VN.n31 VSUBS 0.106432f
C856 VN.n32 VSUBS 0.114491f
C857 VN.n33 VSUBS 0.046459f
C858 VN.n34 VSUBS 0.057106f
C859 VN.n35 VSUBS 0.057106f
C860 VN.n36 VSUBS 0.057106f
C861 VN.n37 VSUBS 0.106432f
C862 VN.n38 VSUBS 0.106432f
C863 VN.t7 VSUBS 0.366143f
C864 VN.n39 VSUBS 0.240566f
C865 VN.n40 VSUBS 0.05809f
C866 VN.n41 VSUBS 0.057106f
C867 VN.n42 VSUBS 0.057106f
C868 VN.n43 VSUBS 0.057106f
C869 VN.n44 VSUBS 0.106432f
C870 VN.n45 VSUBS 0.115394f
C871 VN.n46 VSUBS 0.048861f
C872 VN.n47 VSUBS 0.057106f
C873 VN.n48 VSUBS 0.057106f
C874 VN.n49 VSUBS 0.057106f
C875 VN.n50 VSUBS 0.106432f
C876 VN.n51 VSUBS 0.106432f
C877 VN.n52 VSUBS 0.062293f
C878 VN.n53 VSUBS 0.092169f
C879 VN.n54 VSUBS 0.17085f
C880 VN.t0 VSUBS 0.366143f
C881 VN.n55 VSUBS 0.453197f
C882 VN.n56 VSUBS 0.057106f
C883 VN.n57 VSUBS 0.108907f
C884 VN.n58 VSUBS 0.057106f
C885 VN.n59 VSUBS 0.102229f
C886 VN.n60 VSUBS 0.057106f
C887 VN.t3 VSUBS 0.366143f
C888 VN.n61 VSUBS 0.240566f
C889 VN.n62 VSUBS 0.112213f
C890 VN.n63 VSUBS 0.057106f
C891 VN.n64 VSUBS 0.106432f
C892 VN.n65 VSUBS 0.057106f
C893 VN.t8 VSUBS 0.366143f
C894 VN.n66 VSUBS 0.114491f
C895 VN.n67 VSUBS 0.057106f
C896 VN.n68 VSUBS 0.106432f
C897 VN.t5 VSUBS 0.933614f
C898 VN.n69 VSUBS 0.569694f
C899 VN.t6 VSUBS 0.366143f
C900 VN.n70 VSUBS 0.42325f
C901 VN.n71 VSUBS 0.05809f
C902 VN.n72 VSUBS 0.725776f
C903 VN.n73 VSUBS 0.057106f
C904 VN.n74 VSUBS 0.057106f
C905 VN.n75 VSUBS 0.106432f
C906 VN.n76 VSUBS 0.112213f
C907 VN.n77 VSUBS 0.046459f
C908 VN.n78 VSUBS 0.057106f
C909 VN.n79 VSUBS 0.057106f
C910 VN.n80 VSUBS 0.057106f
C911 VN.n81 VSUBS 0.106432f
C912 VN.n82 VSUBS 0.106432f
C913 VN.n83 VSUBS 0.294452f
C914 VN.n84 VSUBS 0.057106f
C915 VN.n85 VSUBS 0.057106f
C916 VN.n86 VSUBS 0.057106f
C917 VN.n87 VSUBS 0.106432f
C918 VN.n88 VSUBS 0.114491f
C919 VN.n89 VSUBS 0.046459f
C920 VN.n90 VSUBS 0.057106f
C921 VN.n91 VSUBS 0.057106f
C922 VN.n92 VSUBS 0.057106f
C923 VN.n93 VSUBS 0.106432f
C924 VN.n94 VSUBS 0.106432f
C925 VN.n95 VSUBS 0.05809f
C926 VN.n96 VSUBS 0.057106f
C927 VN.n97 VSUBS 0.057106f
C928 VN.n98 VSUBS 0.057106f
C929 VN.n99 VSUBS 0.106432f
C930 VN.n100 VSUBS 0.115394f
C931 VN.n101 VSUBS 0.048861f
C932 VN.n102 VSUBS 0.057106f
C933 VN.n103 VSUBS 0.057106f
C934 VN.n104 VSUBS 0.057106f
C935 VN.n105 VSUBS 0.106432f
C936 VN.n106 VSUBS 0.106432f
C937 VN.n107 VSUBS 0.062293f
C938 VN.n108 VSUBS 0.092169f
C939 VN.n109 VSUBS 3.38122f
C940 VDD1.t3 VSUBS 0.16155f
C941 VDD1.t5 VSUBS 0.030254f
C942 VDD1.t6 VSUBS 0.030254f
C943 VDD1.n0 VSUBS 0.081818f
C944 VDD1.n1 VSUBS 1.66135f
C945 VDD1.t8 VSUBS 0.16155f
C946 VDD1.t4 VSUBS 0.030254f
C947 VDD1.t1 VSUBS 0.030254f
C948 VDD1.n2 VSUBS 0.081818f
C949 VDD1.n3 VSUBS 1.64775f
C950 VDD1.t0 VSUBS 0.030254f
C951 VDD1.t2 VSUBS 0.030254f
C952 VDD1.n4 VSUBS 0.086238f
C953 VDD1.n5 VSUBS 4.78114f
C954 VDD1.t7 VSUBS 0.030254f
C955 VDD1.t9 VSUBS 0.030254f
C956 VDD1.n6 VSUBS 0.081818f
C957 VDD1.n7 VSUBS 4.46068f
C958 VTAIL.t0 VSUBS 0.033751f
C959 VTAIL.t4 VSUBS 0.033751f
C960 VTAIL.n0 VSUBS 0.08228f
C961 VTAIL.n1 VSUBS 0.999321f
C962 VTAIL.t7 VSUBS 0.167004f
C963 VTAIL.n2 VSUBS 1.12435f
C964 VTAIL.t11 VSUBS 0.033751f
C965 VTAIL.t10 VSUBS 0.033751f
C966 VTAIL.n3 VSUBS 0.08228f
C967 VTAIL.n4 VSUBS 1.30123f
C968 VTAIL.t12 VSUBS 0.033751f
C969 VTAIL.t15 VSUBS 0.033751f
C970 VTAIL.n5 VSUBS 0.08228f
C971 VTAIL.n6 VSUBS 2.53512f
C972 VTAIL.t17 VSUBS 0.033751f
C973 VTAIL.t19 VSUBS 0.033751f
C974 VTAIL.n7 VSUBS 0.08228f
C975 VTAIL.n8 VSUBS 2.53512f
C976 VTAIL.t3 VSUBS 0.033751f
C977 VTAIL.t18 VSUBS 0.033751f
C978 VTAIL.n9 VSUBS 0.08228f
C979 VTAIL.n10 VSUBS 1.30123f
C980 VTAIL.t5 VSUBS 0.167005f
C981 VTAIL.n11 VSUBS 1.12435f
C982 VTAIL.t16 VSUBS 0.033751f
C983 VTAIL.t13 VSUBS 0.033751f
C984 VTAIL.n12 VSUBS 0.08228f
C985 VTAIL.n13 VSUBS 1.11703f
C986 VTAIL.t8 VSUBS 0.033751f
C987 VTAIL.t9 VSUBS 0.033751f
C988 VTAIL.n14 VSUBS 0.08228f
C989 VTAIL.n15 VSUBS 1.30123f
C990 VTAIL.t14 VSUBS 0.167005f
C991 VTAIL.n16 VSUBS 2.03791f
C992 VTAIL.t6 VSUBS 0.167004f
C993 VTAIL.n17 VSUBS 2.03791f
C994 VTAIL.t1 VSUBS 0.033751f
C995 VTAIL.t2 VSUBS 0.033751f
C996 VTAIL.n18 VSUBS 0.08228f
C997 VTAIL.n19 VSUBS 0.9144f
C998 VP.t7 VSUBS 0.41854f
C999 VP.n0 VSUBS 0.518052f
C1000 VP.n1 VSUBS 0.065279f
C1001 VP.n2 VSUBS 0.124492f
C1002 VP.n3 VSUBS 0.065279f
C1003 VP.n4 VSUBS 0.116858f
C1004 VP.n5 VSUBS 0.065279f
C1005 VP.n6 VSUBS 0.128271f
C1006 VP.n7 VSUBS 0.065279f
C1007 VP.n8 VSUBS 0.121663f
C1008 VP.n9 VSUBS 0.065279f
C1009 VP.t8 VSUBS 0.41854f
C1010 VP.n10 VSUBS 0.130875f
C1011 VP.n11 VSUBS 0.065279f
C1012 VP.n12 VSUBS 0.121663f
C1013 VP.n13 VSUBS 0.065279f
C1014 VP.t5 VSUBS 0.41854f
C1015 VP.n14 VSUBS 0.131908f
C1016 VP.n15 VSUBS 0.065279f
C1017 VP.n16 VSUBS 0.121663f
C1018 VP.t0 VSUBS 0.41854f
C1019 VP.n17 VSUBS 0.518052f
C1020 VP.n18 VSUBS 0.065279f
C1021 VP.n19 VSUBS 0.124492f
C1022 VP.n20 VSUBS 0.065279f
C1023 VP.n21 VSUBS 0.116858f
C1024 VP.n22 VSUBS 0.065279f
C1025 VP.n23 VSUBS 0.128271f
C1026 VP.n24 VSUBS 0.065279f
C1027 VP.n25 VSUBS 0.121663f
C1028 VP.n26 VSUBS 0.065279f
C1029 VP.t3 VSUBS 0.41854f
C1030 VP.n27 VSUBS 0.130875f
C1031 VP.n28 VSUBS 0.065279f
C1032 VP.n29 VSUBS 0.121663f
C1033 VP.t6 VSUBS 1.06722f
C1034 VP.n30 VSUBS 0.651221f
C1035 VP.t4 VSUBS 0.41854f
C1036 VP.n31 VSUBS 0.483819f
C1037 VP.n32 VSUBS 0.066403f
C1038 VP.n33 VSUBS 0.82964f
C1039 VP.n34 VSUBS 0.065279f
C1040 VP.n35 VSUBS 0.065279f
C1041 VP.n36 VSUBS 0.121663f
C1042 VP.n37 VSUBS 0.128271f
C1043 VP.n38 VSUBS 0.053108f
C1044 VP.n39 VSUBS 0.065279f
C1045 VP.n40 VSUBS 0.065279f
C1046 VP.n41 VSUBS 0.065279f
C1047 VP.n42 VSUBS 0.121663f
C1048 VP.n43 VSUBS 0.121663f
C1049 VP.n44 VSUBS 0.336589f
C1050 VP.n45 VSUBS 0.065279f
C1051 VP.n46 VSUBS 0.065279f
C1052 VP.n47 VSUBS 0.065279f
C1053 VP.n48 VSUBS 0.121663f
C1054 VP.n49 VSUBS 0.130875f
C1055 VP.n50 VSUBS 0.053108f
C1056 VP.n51 VSUBS 0.065279f
C1057 VP.n52 VSUBS 0.065279f
C1058 VP.n53 VSUBS 0.065279f
C1059 VP.n54 VSUBS 0.121663f
C1060 VP.n55 VSUBS 0.121663f
C1061 VP.t2 VSUBS 0.41854f
C1062 VP.n56 VSUBS 0.274992f
C1063 VP.n57 VSUBS 0.066403f
C1064 VP.n58 VSUBS 0.065279f
C1065 VP.n59 VSUBS 0.065279f
C1066 VP.n60 VSUBS 0.065279f
C1067 VP.n61 VSUBS 0.121663f
C1068 VP.n62 VSUBS 0.131908f
C1069 VP.n63 VSUBS 0.055854f
C1070 VP.n64 VSUBS 0.065279f
C1071 VP.n65 VSUBS 0.065279f
C1072 VP.n66 VSUBS 0.065279f
C1073 VP.n67 VSUBS 0.121663f
C1074 VP.n68 VSUBS 0.121663f
C1075 VP.n69 VSUBS 0.071208f
C1076 VP.n70 VSUBS 0.105359f
C1077 VP.n71 VSUBS 3.83853f
C1078 VP.n72 VSUBS 3.8847f
C1079 VP.t1 VSUBS 0.41854f
C1080 VP.n73 VSUBS 0.518052f
C1081 VP.n74 VSUBS 0.071208f
C1082 VP.n75 VSUBS 0.105359f
C1083 VP.n76 VSUBS 0.065279f
C1084 VP.n77 VSUBS 0.065279f
C1085 VP.n78 VSUBS 0.121663f
C1086 VP.n79 VSUBS 0.124492f
C1087 VP.n80 VSUBS 0.055854f
C1088 VP.n81 VSUBS 0.065279f
C1089 VP.n82 VSUBS 0.065279f
C1090 VP.n83 VSUBS 0.065279f
C1091 VP.n84 VSUBS 0.121663f
C1092 VP.n85 VSUBS 0.116858f
C1093 VP.n86 VSUBS 0.274992f
C1094 VP.n87 VSUBS 0.066403f
C1095 VP.n88 VSUBS 0.065279f
C1096 VP.n89 VSUBS 0.065279f
C1097 VP.n90 VSUBS 0.065279f
C1098 VP.n91 VSUBS 0.121663f
C1099 VP.n92 VSUBS 0.128271f
C1100 VP.n93 VSUBS 0.053108f
C1101 VP.n94 VSUBS 0.065279f
C1102 VP.n95 VSUBS 0.065279f
C1103 VP.n96 VSUBS 0.065279f
C1104 VP.n97 VSUBS 0.121663f
C1105 VP.n98 VSUBS 0.121663f
C1106 VP.n99 VSUBS 0.336589f
C1107 VP.n100 VSUBS 0.065279f
C1108 VP.n101 VSUBS 0.065279f
C1109 VP.n102 VSUBS 0.065279f
C1110 VP.n103 VSUBS 0.121663f
C1111 VP.n104 VSUBS 0.130875f
C1112 VP.n105 VSUBS 0.053108f
C1113 VP.n106 VSUBS 0.065279f
C1114 VP.n107 VSUBS 0.065279f
C1115 VP.n108 VSUBS 0.065279f
C1116 VP.n109 VSUBS 0.121663f
C1117 VP.n110 VSUBS 0.121663f
C1118 VP.t9 VSUBS 0.41854f
C1119 VP.n111 VSUBS 0.274992f
C1120 VP.n112 VSUBS 0.066403f
C1121 VP.n113 VSUBS 0.065279f
C1122 VP.n114 VSUBS 0.065279f
C1123 VP.n115 VSUBS 0.065279f
C1124 VP.n116 VSUBS 0.121663f
C1125 VP.n117 VSUBS 0.131908f
C1126 VP.n118 VSUBS 0.055854f
C1127 VP.n119 VSUBS 0.065279f
C1128 VP.n120 VSUBS 0.065279f
C1129 VP.n121 VSUBS 0.065279f
C1130 VP.n122 VSUBS 0.121663f
C1131 VP.n123 VSUBS 0.121663f
C1132 VP.n124 VSUBS 0.071208f
C1133 VP.n125 VSUBS 0.105359f
C1134 VP.n126 VSUBS 0.195299f
.ends

