* NGSPICE file created from diff_pair_sample_1603.ext - technology: sky130A

.subckt diff_pair_sample_1603 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=2.6481 ps=14.36 w=6.79 l=3.17
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=2.6481 ps=14.36 w=6.79 l=3.17
X2 B.t11 B.t9 B.t10 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=0 ps=0 w=6.79 l=3.17
X3 B.t8 B.t6 B.t7 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=0 ps=0 w=6.79 l=3.17
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=2.6481 ps=14.36 w=6.79 l=3.17
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=2.6481 ps=14.36 w=6.79 l=3.17
X6 B.t5 B.t3 B.t4 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=0 ps=0 w=6.79 l=3.17
X7 B.t2 B.t0 B.t1 w_n2370_n2326# sky130_fd_pr__pfet_01v8 ad=2.6481 pd=14.36 as=0 ps=0 w=6.79 l=3.17
R0 VN VN.t1 132.537
R1 VN VN.t0 90.9352
R2 VTAIL.n138 VTAIL.n108 756.745
R3 VTAIL.n30 VTAIL.n0 756.745
R4 VTAIL.n102 VTAIL.n72 756.745
R5 VTAIL.n66 VTAIL.n36 756.745
R6 VTAIL.n121 VTAIL.n120 585
R7 VTAIL.n123 VTAIL.n122 585
R8 VTAIL.n116 VTAIL.n115 585
R9 VTAIL.n129 VTAIL.n128 585
R10 VTAIL.n131 VTAIL.n130 585
R11 VTAIL.n112 VTAIL.n111 585
R12 VTAIL.n137 VTAIL.n136 585
R13 VTAIL.n139 VTAIL.n138 585
R14 VTAIL.n13 VTAIL.n12 585
R15 VTAIL.n15 VTAIL.n14 585
R16 VTAIL.n8 VTAIL.n7 585
R17 VTAIL.n21 VTAIL.n20 585
R18 VTAIL.n23 VTAIL.n22 585
R19 VTAIL.n4 VTAIL.n3 585
R20 VTAIL.n29 VTAIL.n28 585
R21 VTAIL.n31 VTAIL.n30 585
R22 VTAIL.n103 VTAIL.n102 585
R23 VTAIL.n101 VTAIL.n100 585
R24 VTAIL.n76 VTAIL.n75 585
R25 VTAIL.n95 VTAIL.n94 585
R26 VTAIL.n93 VTAIL.n92 585
R27 VTAIL.n80 VTAIL.n79 585
R28 VTAIL.n87 VTAIL.n86 585
R29 VTAIL.n85 VTAIL.n84 585
R30 VTAIL.n67 VTAIL.n66 585
R31 VTAIL.n65 VTAIL.n64 585
R32 VTAIL.n40 VTAIL.n39 585
R33 VTAIL.n59 VTAIL.n58 585
R34 VTAIL.n57 VTAIL.n56 585
R35 VTAIL.n44 VTAIL.n43 585
R36 VTAIL.n51 VTAIL.n50 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n119 VTAIL.t3 327.514
R39 VTAIL.n11 VTAIL.t1 327.514
R40 VTAIL.n83 VTAIL.t0 327.514
R41 VTAIL.n47 VTAIL.t2 327.514
R42 VTAIL.n122 VTAIL.n121 171.744
R43 VTAIL.n122 VTAIL.n115 171.744
R44 VTAIL.n129 VTAIL.n115 171.744
R45 VTAIL.n130 VTAIL.n129 171.744
R46 VTAIL.n130 VTAIL.n111 171.744
R47 VTAIL.n137 VTAIL.n111 171.744
R48 VTAIL.n138 VTAIL.n137 171.744
R49 VTAIL.n14 VTAIL.n13 171.744
R50 VTAIL.n14 VTAIL.n7 171.744
R51 VTAIL.n21 VTAIL.n7 171.744
R52 VTAIL.n22 VTAIL.n21 171.744
R53 VTAIL.n22 VTAIL.n3 171.744
R54 VTAIL.n29 VTAIL.n3 171.744
R55 VTAIL.n30 VTAIL.n29 171.744
R56 VTAIL.n102 VTAIL.n101 171.744
R57 VTAIL.n101 VTAIL.n75 171.744
R58 VTAIL.n94 VTAIL.n75 171.744
R59 VTAIL.n94 VTAIL.n93 171.744
R60 VTAIL.n93 VTAIL.n79 171.744
R61 VTAIL.n86 VTAIL.n79 171.744
R62 VTAIL.n86 VTAIL.n85 171.744
R63 VTAIL.n66 VTAIL.n65 171.744
R64 VTAIL.n65 VTAIL.n39 171.744
R65 VTAIL.n58 VTAIL.n39 171.744
R66 VTAIL.n58 VTAIL.n57 171.744
R67 VTAIL.n57 VTAIL.n43 171.744
R68 VTAIL.n50 VTAIL.n43 171.744
R69 VTAIL.n50 VTAIL.n49 171.744
R70 VTAIL.n121 VTAIL.t3 85.8723
R71 VTAIL.n13 VTAIL.t1 85.8723
R72 VTAIL.n85 VTAIL.t0 85.8723
R73 VTAIL.n49 VTAIL.t2 85.8723
R74 VTAIL.n143 VTAIL.n142 33.5429
R75 VTAIL.n35 VTAIL.n34 33.5429
R76 VTAIL.n107 VTAIL.n106 33.5429
R77 VTAIL.n71 VTAIL.n70 33.5429
R78 VTAIL.n71 VTAIL.n35 24.2548
R79 VTAIL.n143 VTAIL.n107 21.2376
R80 VTAIL.n120 VTAIL.n119 16.3884
R81 VTAIL.n12 VTAIL.n11 16.3884
R82 VTAIL.n84 VTAIL.n83 16.3884
R83 VTAIL.n48 VTAIL.n47 16.3884
R84 VTAIL.n123 VTAIL.n118 12.8005
R85 VTAIL.n15 VTAIL.n10 12.8005
R86 VTAIL.n87 VTAIL.n82 12.8005
R87 VTAIL.n51 VTAIL.n46 12.8005
R88 VTAIL.n124 VTAIL.n116 12.0247
R89 VTAIL.n16 VTAIL.n8 12.0247
R90 VTAIL.n88 VTAIL.n80 12.0247
R91 VTAIL.n52 VTAIL.n44 12.0247
R92 VTAIL.n128 VTAIL.n127 11.249
R93 VTAIL.n20 VTAIL.n19 11.249
R94 VTAIL.n92 VTAIL.n91 11.249
R95 VTAIL.n56 VTAIL.n55 11.249
R96 VTAIL.n131 VTAIL.n114 10.4732
R97 VTAIL.n23 VTAIL.n6 10.4732
R98 VTAIL.n95 VTAIL.n78 10.4732
R99 VTAIL.n59 VTAIL.n42 10.4732
R100 VTAIL.n132 VTAIL.n112 9.69747
R101 VTAIL.n24 VTAIL.n4 9.69747
R102 VTAIL.n96 VTAIL.n76 9.69747
R103 VTAIL.n60 VTAIL.n40 9.69747
R104 VTAIL.n142 VTAIL.n141 9.45567
R105 VTAIL.n34 VTAIL.n33 9.45567
R106 VTAIL.n106 VTAIL.n105 9.45567
R107 VTAIL.n70 VTAIL.n69 9.45567
R108 VTAIL.n110 VTAIL.n109 9.3005
R109 VTAIL.n135 VTAIL.n134 9.3005
R110 VTAIL.n133 VTAIL.n132 9.3005
R111 VTAIL.n114 VTAIL.n113 9.3005
R112 VTAIL.n127 VTAIL.n126 9.3005
R113 VTAIL.n125 VTAIL.n124 9.3005
R114 VTAIL.n118 VTAIL.n117 9.3005
R115 VTAIL.n141 VTAIL.n140 9.3005
R116 VTAIL.n2 VTAIL.n1 9.3005
R117 VTAIL.n27 VTAIL.n26 9.3005
R118 VTAIL.n25 VTAIL.n24 9.3005
R119 VTAIL.n6 VTAIL.n5 9.3005
R120 VTAIL.n19 VTAIL.n18 9.3005
R121 VTAIL.n17 VTAIL.n16 9.3005
R122 VTAIL.n10 VTAIL.n9 9.3005
R123 VTAIL.n33 VTAIL.n32 9.3005
R124 VTAIL.n105 VTAIL.n104 9.3005
R125 VTAIL.n74 VTAIL.n73 9.3005
R126 VTAIL.n99 VTAIL.n98 9.3005
R127 VTAIL.n97 VTAIL.n96 9.3005
R128 VTAIL.n78 VTAIL.n77 9.3005
R129 VTAIL.n91 VTAIL.n90 9.3005
R130 VTAIL.n89 VTAIL.n88 9.3005
R131 VTAIL.n82 VTAIL.n81 9.3005
R132 VTAIL.n69 VTAIL.n68 9.3005
R133 VTAIL.n38 VTAIL.n37 9.3005
R134 VTAIL.n63 VTAIL.n62 9.3005
R135 VTAIL.n61 VTAIL.n60 9.3005
R136 VTAIL.n42 VTAIL.n41 9.3005
R137 VTAIL.n55 VTAIL.n54 9.3005
R138 VTAIL.n53 VTAIL.n52 9.3005
R139 VTAIL.n46 VTAIL.n45 9.3005
R140 VTAIL.n136 VTAIL.n135 8.92171
R141 VTAIL.n28 VTAIL.n27 8.92171
R142 VTAIL.n100 VTAIL.n99 8.92171
R143 VTAIL.n64 VTAIL.n63 8.92171
R144 VTAIL.n139 VTAIL.n110 8.14595
R145 VTAIL.n31 VTAIL.n2 8.14595
R146 VTAIL.n103 VTAIL.n74 8.14595
R147 VTAIL.n67 VTAIL.n38 8.14595
R148 VTAIL.n140 VTAIL.n108 7.3702
R149 VTAIL.n32 VTAIL.n0 7.3702
R150 VTAIL.n104 VTAIL.n72 7.3702
R151 VTAIL.n68 VTAIL.n36 7.3702
R152 VTAIL.n142 VTAIL.n108 6.59444
R153 VTAIL.n34 VTAIL.n0 6.59444
R154 VTAIL.n106 VTAIL.n72 6.59444
R155 VTAIL.n70 VTAIL.n36 6.59444
R156 VTAIL.n140 VTAIL.n139 5.81868
R157 VTAIL.n32 VTAIL.n31 5.81868
R158 VTAIL.n104 VTAIL.n103 5.81868
R159 VTAIL.n68 VTAIL.n67 5.81868
R160 VTAIL.n136 VTAIL.n110 5.04292
R161 VTAIL.n28 VTAIL.n2 5.04292
R162 VTAIL.n100 VTAIL.n74 5.04292
R163 VTAIL.n64 VTAIL.n38 5.04292
R164 VTAIL.n135 VTAIL.n112 4.26717
R165 VTAIL.n27 VTAIL.n4 4.26717
R166 VTAIL.n99 VTAIL.n76 4.26717
R167 VTAIL.n63 VTAIL.n40 4.26717
R168 VTAIL.n119 VTAIL.n117 3.71088
R169 VTAIL.n11 VTAIL.n9 3.71088
R170 VTAIL.n83 VTAIL.n81 3.71088
R171 VTAIL.n47 VTAIL.n45 3.71088
R172 VTAIL.n132 VTAIL.n131 3.49141
R173 VTAIL.n24 VTAIL.n23 3.49141
R174 VTAIL.n96 VTAIL.n95 3.49141
R175 VTAIL.n60 VTAIL.n59 3.49141
R176 VTAIL.n128 VTAIL.n114 2.71565
R177 VTAIL.n20 VTAIL.n6 2.71565
R178 VTAIL.n92 VTAIL.n78 2.71565
R179 VTAIL.n56 VTAIL.n42 2.71565
R180 VTAIL.n107 VTAIL.n71 1.97895
R181 VTAIL.n127 VTAIL.n116 1.93989
R182 VTAIL.n19 VTAIL.n8 1.93989
R183 VTAIL.n91 VTAIL.n80 1.93989
R184 VTAIL.n55 VTAIL.n44 1.93989
R185 VTAIL VTAIL.n35 1.28283
R186 VTAIL.n124 VTAIL.n123 1.16414
R187 VTAIL.n16 VTAIL.n15 1.16414
R188 VTAIL.n88 VTAIL.n87 1.16414
R189 VTAIL.n52 VTAIL.n51 1.16414
R190 VTAIL VTAIL.n143 0.696621
R191 VTAIL.n120 VTAIL.n118 0.388379
R192 VTAIL.n12 VTAIL.n10 0.388379
R193 VTAIL.n84 VTAIL.n82 0.388379
R194 VTAIL.n48 VTAIL.n46 0.388379
R195 VTAIL.n125 VTAIL.n117 0.155672
R196 VTAIL.n126 VTAIL.n125 0.155672
R197 VTAIL.n126 VTAIL.n113 0.155672
R198 VTAIL.n133 VTAIL.n113 0.155672
R199 VTAIL.n134 VTAIL.n133 0.155672
R200 VTAIL.n134 VTAIL.n109 0.155672
R201 VTAIL.n141 VTAIL.n109 0.155672
R202 VTAIL.n17 VTAIL.n9 0.155672
R203 VTAIL.n18 VTAIL.n17 0.155672
R204 VTAIL.n18 VTAIL.n5 0.155672
R205 VTAIL.n25 VTAIL.n5 0.155672
R206 VTAIL.n26 VTAIL.n25 0.155672
R207 VTAIL.n26 VTAIL.n1 0.155672
R208 VTAIL.n33 VTAIL.n1 0.155672
R209 VTAIL.n105 VTAIL.n73 0.155672
R210 VTAIL.n98 VTAIL.n73 0.155672
R211 VTAIL.n98 VTAIL.n97 0.155672
R212 VTAIL.n97 VTAIL.n77 0.155672
R213 VTAIL.n90 VTAIL.n77 0.155672
R214 VTAIL.n90 VTAIL.n89 0.155672
R215 VTAIL.n89 VTAIL.n81 0.155672
R216 VTAIL.n69 VTAIL.n37 0.155672
R217 VTAIL.n62 VTAIL.n37 0.155672
R218 VTAIL.n62 VTAIL.n61 0.155672
R219 VTAIL.n61 VTAIL.n41 0.155672
R220 VTAIL.n54 VTAIL.n41 0.155672
R221 VTAIL.n54 VTAIL.n53 0.155672
R222 VTAIL.n53 VTAIL.n45 0.155672
R223 VDD2.n65 VDD2.n35 756.745
R224 VDD2.n30 VDD2.n0 756.745
R225 VDD2.n66 VDD2.n65 585
R226 VDD2.n64 VDD2.n63 585
R227 VDD2.n39 VDD2.n38 585
R228 VDD2.n58 VDD2.n57 585
R229 VDD2.n56 VDD2.n55 585
R230 VDD2.n43 VDD2.n42 585
R231 VDD2.n50 VDD2.n49 585
R232 VDD2.n48 VDD2.n47 585
R233 VDD2.n13 VDD2.n12 585
R234 VDD2.n15 VDD2.n14 585
R235 VDD2.n8 VDD2.n7 585
R236 VDD2.n21 VDD2.n20 585
R237 VDD2.n23 VDD2.n22 585
R238 VDD2.n4 VDD2.n3 585
R239 VDD2.n29 VDD2.n28 585
R240 VDD2.n31 VDD2.n30 585
R241 VDD2.n46 VDD2.t0 327.514
R242 VDD2.n11 VDD2.t1 327.514
R243 VDD2.n65 VDD2.n64 171.744
R244 VDD2.n64 VDD2.n38 171.744
R245 VDD2.n57 VDD2.n38 171.744
R246 VDD2.n57 VDD2.n56 171.744
R247 VDD2.n56 VDD2.n42 171.744
R248 VDD2.n49 VDD2.n42 171.744
R249 VDD2.n49 VDD2.n48 171.744
R250 VDD2.n14 VDD2.n13 171.744
R251 VDD2.n14 VDD2.n7 171.744
R252 VDD2.n21 VDD2.n7 171.744
R253 VDD2.n22 VDD2.n21 171.744
R254 VDD2.n22 VDD2.n3 171.744
R255 VDD2.n29 VDD2.n3 171.744
R256 VDD2.n30 VDD2.n29 171.744
R257 VDD2.n48 VDD2.t0 85.8723
R258 VDD2.n13 VDD2.t1 85.8723
R259 VDD2.n70 VDD2.n34 85.7691
R260 VDD2.n70 VDD2.n69 50.2217
R261 VDD2.n12 VDD2.n11 16.3884
R262 VDD2.n47 VDD2.n46 16.3884
R263 VDD2.n50 VDD2.n45 12.8005
R264 VDD2.n15 VDD2.n10 12.8005
R265 VDD2.n51 VDD2.n43 12.0247
R266 VDD2.n16 VDD2.n8 12.0247
R267 VDD2.n55 VDD2.n54 11.249
R268 VDD2.n20 VDD2.n19 11.249
R269 VDD2.n58 VDD2.n41 10.4732
R270 VDD2.n23 VDD2.n6 10.4732
R271 VDD2.n59 VDD2.n39 9.69747
R272 VDD2.n24 VDD2.n4 9.69747
R273 VDD2.n69 VDD2.n68 9.45567
R274 VDD2.n34 VDD2.n33 9.45567
R275 VDD2.n68 VDD2.n67 9.3005
R276 VDD2.n37 VDD2.n36 9.3005
R277 VDD2.n62 VDD2.n61 9.3005
R278 VDD2.n60 VDD2.n59 9.3005
R279 VDD2.n41 VDD2.n40 9.3005
R280 VDD2.n54 VDD2.n53 9.3005
R281 VDD2.n52 VDD2.n51 9.3005
R282 VDD2.n45 VDD2.n44 9.3005
R283 VDD2.n2 VDD2.n1 9.3005
R284 VDD2.n27 VDD2.n26 9.3005
R285 VDD2.n25 VDD2.n24 9.3005
R286 VDD2.n6 VDD2.n5 9.3005
R287 VDD2.n19 VDD2.n18 9.3005
R288 VDD2.n17 VDD2.n16 9.3005
R289 VDD2.n10 VDD2.n9 9.3005
R290 VDD2.n33 VDD2.n32 9.3005
R291 VDD2.n63 VDD2.n62 8.92171
R292 VDD2.n28 VDD2.n27 8.92171
R293 VDD2.n66 VDD2.n37 8.14595
R294 VDD2.n31 VDD2.n2 8.14595
R295 VDD2.n67 VDD2.n35 7.3702
R296 VDD2.n32 VDD2.n0 7.3702
R297 VDD2.n69 VDD2.n35 6.59444
R298 VDD2.n34 VDD2.n0 6.59444
R299 VDD2.n67 VDD2.n66 5.81868
R300 VDD2.n32 VDD2.n31 5.81868
R301 VDD2.n63 VDD2.n37 5.04292
R302 VDD2.n28 VDD2.n2 5.04292
R303 VDD2.n62 VDD2.n39 4.26717
R304 VDD2.n27 VDD2.n4 4.26717
R305 VDD2.n46 VDD2.n44 3.71088
R306 VDD2.n11 VDD2.n9 3.71088
R307 VDD2.n59 VDD2.n58 3.49141
R308 VDD2.n24 VDD2.n23 3.49141
R309 VDD2.n55 VDD2.n41 2.71565
R310 VDD2.n20 VDD2.n6 2.71565
R311 VDD2.n54 VDD2.n43 1.93989
R312 VDD2.n19 VDD2.n8 1.93989
R313 VDD2.n51 VDD2.n50 1.16414
R314 VDD2.n16 VDD2.n15 1.16414
R315 VDD2 VDD2.n70 0.813
R316 VDD2.n47 VDD2.n45 0.388379
R317 VDD2.n12 VDD2.n10 0.388379
R318 VDD2.n68 VDD2.n36 0.155672
R319 VDD2.n61 VDD2.n36 0.155672
R320 VDD2.n61 VDD2.n60 0.155672
R321 VDD2.n60 VDD2.n40 0.155672
R322 VDD2.n53 VDD2.n40 0.155672
R323 VDD2.n53 VDD2.n52 0.155672
R324 VDD2.n52 VDD2.n44 0.155672
R325 VDD2.n17 VDD2.n9 0.155672
R326 VDD2.n18 VDD2.n17 0.155672
R327 VDD2.n18 VDD2.n5 0.155672
R328 VDD2.n25 VDD2.n5 0.155672
R329 VDD2.n26 VDD2.n25 0.155672
R330 VDD2.n26 VDD2.n1 0.155672
R331 VDD2.n33 VDD2.n1 0.155672
R332 VP.n0 VP.t1 132.631
R333 VP.n0 VP.t0 90.4094
R334 VP VP.n0 0.52637
R335 VDD1.n30 VDD1.n0 756.745
R336 VDD1.n65 VDD1.n35 756.745
R337 VDD1.n31 VDD1.n30 585
R338 VDD1.n29 VDD1.n28 585
R339 VDD1.n4 VDD1.n3 585
R340 VDD1.n23 VDD1.n22 585
R341 VDD1.n21 VDD1.n20 585
R342 VDD1.n8 VDD1.n7 585
R343 VDD1.n15 VDD1.n14 585
R344 VDD1.n13 VDD1.n12 585
R345 VDD1.n48 VDD1.n47 585
R346 VDD1.n50 VDD1.n49 585
R347 VDD1.n43 VDD1.n42 585
R348 VDD1.n56 VDD1.n55 585
R349 VDD1.n58 VDD1.n57 585
R350 VDD1.n39 VDD1.n38 585
R351 VDD1.n64 VDD1.n63 585
R352 VDD1.n66 VDD1.n65 585
R353 VDD1.n11 VDD1.t0 327.514
R354 VDD1.n46 VDD1.t1 327.514
R355 VDD1.n30 VDD1.n29 171.744
R356 VDD1.n29 VDD1.n3 171.744
R357 VDD1.n22 VDD1.n3 171.744
R358 VDD1.n22 VDD1.n21 171.744
R359 VDD1.n21 VDD1.n7 171.744
R360 VDD1.n14 VDD1.n7 171.744
R361 VDD1.n14 VDD1.n13 171.744
R362 VDD1.n49 VDD1.n48 171.744
R363 VDD1.n49 VDD1.n42 171.744
R364 VDD1.n56 VDD1.n42 171.744
R365 VDD1.n57 VDD1.n56 171.744
R366 VDD1.n57 VDD1.n38 171.744
R367 VDD1.n64 VDD1.n38 171.744
R368 VDD1.n65 VDD1.n64 171.744
R369 VDD1 VDD1.n69 87.0482
R370 VDD1.n13 VDD1.t0 85.8723
R371 VDD1.n48 VDD1.t1 85.8723
R372 VDD1 VDD1.n34 51.0342
R373 VDD1.n47 VDD1.n46 16.3884
R374 VDD1.n12 VDD1.n11 16.3884
R375 VDD1.n15 VDD1.n10 12.8005
R376 VDD1.n50 VDD1.n45 12.8005
R377 VDD1.n16 VDD1.n8 12.0247
R378 VDD1.n51 VDD1.n43 12.0247
R379 VDD1.n20 VDD1.n19 11.249
R380 VDD1.n55 VDD1.n54 11.249
R381 VDD1.n23 VDD1.n6 10.4732
R382 VDD1.n58 VDD1.n41 10.4732
R383 VDD1.n24 VDD1.n4 9.69747
R384 VDD1.n59 VDD1.n39 9.69747
R385 VDD1.n34 VDD1.n33 9.45567
R386 VDD1.n69 VDD1.n68 9.45567
R387 VDD1.n33 VDD1.n32 9.3005
R388 VDD1.n2 VDD1.n1 9.3005
R389 VDD1.n27 VDD1.n26 9.3005
R390 VDD1.n25 VDD1.n24 9.3005
R391 VDD1.n6 VDD1.n5 9.3005
R392 VDD1.n19 VDD1.n18 9.3005
R393 VDD1.n17 VDD1.n16 9.3005
R394 VDD1.n10 VDD1.n9 9.3005
R395 VDD1.n37 VDD1.n36 9.3005
R396 VDD1.n62 VDD1.n61 9.3005
R397 VDD1.n60 VDD1.n59 9.3005
R398 VDD1.n41 VDD1.n40 9.3005
R399 VDD1.n54 VDD1.n53 9.3005
R400 VDD1.n52 VDD1.n51 9.3005
R401 VDD1.n45 VDD1.n44 9.3005
R402 VDD1.n68 VDD1.n67 9.3005
R403 VDD1.n28 VDD1.n27 8.92171
R404 VDD1.n63 VDD1.n62 8.92171
R405 VDD1.n31 VDD1.n2 8.14595
R406 VDD1.n66 VDD1.n37 8.14595
R407 VDD1.n32 VDD1.n0 7.3702
R408 VDD1.n67 VDD1.n35 7.3702
R409 VDD1.n34 VDD1.n0 6.59444
R410 VDD1.n69 VDD1.n35 6.59444
R411 VDD1.n32 VDD1.n31 5.81868
R412 VDD1.n67 VDD1.n66 5.81868
R413 VDD1.n28 VDD1.n2 5.04292
R414 VDD1.n63 VDD1.n37 5.04292
R415 VDD1.n27 VDD1.n4 4.26717
R416 VDD1.n62 VDD1.n39 4.26717
R417 VDD1.n11 VDD1.n9 3.71088
R418 VDD1.n46 VDD1.n44 3.71088
R419 VDD1.n24 VDD1.n23 3.49141
R420 VDD1.n59 VDD1.n58 3.49141
R421 VDD1.n20 VDD1.n6 2.71565
R422 VDD1.n55 VDD1.n41 2.71565
R423 VDD1.n19 VDD1.n8 1.93989
R424 VDD1.n54 VDD1.n43 1.93989
R425 VDD1.n16 VDD1.n15 1.16414
R426 VDD1.n51 VDD1.n50 1.16414
R427 VDD1.n12 VDD1.n10 0.388379
R428 VDD1.n47 VDD1.n45 0.388379
R429 VDD1.n33 VDD1.n1 0.155672
R430 VDD1.n26 VDD1.n1 0.155672
R431 VDD1.n26 VDD1.n25 0.155672
R432 VDD1.n25 VDD1.n5 0.155672
R433 VDD1.n18 VDD1.n5 0.155672
R434 VDD1.n18 VDD1.n17 0.155672
R435 VDD1.n17 VDD1.n9 0.155672
R436 VDD1.n52 VDD1.n44 0.155672
R437 VDD1.n53 VDD1.n52 0.155672
R438 VDD1.n53 VDD1.n40 0.155672
R439 VDD1.n60 VDD1.n40 0.155672
R440 VDD1.n61 VDD1.n60 0.155672
R441 VDD1.n61 VDD1.n36 0.155672
R442 VDD1.n68 VDD1.n36 0.155672
R443 B.n264 B.n263 585
R444 B.n262 B.n81 585
R445 B.n261 B.n260 585
R446 B.n259 B.n82 585
R447 B.n258 B.n257 585
R448 B.n256 B.n83 585
R449 B.n255 B.n254 585
R450 B.n253 B.n84 585
R451 B.n252 B.n251 585
R452 B.n250 B.n85 585
R453 B.n249 B.n248 585
R454 B.n247 B.n86 585
R455 B.n246 B.n245 585
R456 B.n244 B.n87 585
R457 B.n243 B.n242 585
R458 B.n241 B.n88 585
R459 B.n240 B.n239 585
R460 B.n238 B.n89 585
R461 B.n237 B.n236 585
R462 B.n235 B.n90 585
R463 B.n234 B.n233 585
R464 B.n232 B.n91 585
R465 B.n231 B.n230 585
R466 B.n229 B.n92 585
R467 B.n228 B.n227 585
R468 B.n226 B.n93 585
R469 B.n224 B.n223 585
R470 B.n222 B.n96 585
R471 B.n221 B.n220 585
R472 B.n219 B.n97 585
R473 B.n218 B.n217 585
R474 B.n216 B.n98 585
R475 B.n215 B.n214 585
R476 B.n213 B.n99 585
R477 B.n212 B.n211 585
R478 B.n210 B.n100 585
R479 B.n209 B.n208 585
R480 B.n204 B.n101 585
R481 B.n203 B.n202 585
R482 B.n201 B.n102 585
R483 B.n200 B.n199 585
R484 B.n198 B.n103 585
R485 B.n197 B.n196 585
R486 B.n195 B.n104 585
R487 B.n194 B.n193 585
R488 B.n192 B.n105 585
R489 B.n191 B.n190 585
R490 B.n189 B.n106 585
R491 B.n188 B.n187 585
R492 B.n186 B.n107 585
R493 B.n185 B.n184 585
R494 B.n183 B.n108 585
R495 B.n182 B.n181 585
R496 B.n180 B.n109 585
R497 B.n179 B.n178 585
R498 B.n177 B.n110 585
R499 B.n176 B.n175 585
R500 B.n174 B.n111 585
R501 B.n173 B.n172 585
R502 B.n171 B.n112 585
R503 B.n170 B.n169 585
R504 B.n168 B.n113 585
R505 B.n265 B.n80 585
R506 B.n267 B.n266 585
R507 B.n268 B.n79 585
R508 B.n270 B.n269 585
R509 B.n271 B.n78 585
R510 B.n273 B.n272 585
R511 B.n274 B.n77 585
R512 B.n276 B.n275 585
R513 B.n277 B.n76 585
R514 B.n279 B.n278 585
R515 B.n280 B.n75 585
R516 B.n282 B.n281 585
R517 B.n283 B.n74 585
R518 B.n285 B.n284 585
R519 B.n286 B.n73 585
R520 B.n288 B.n287 585
R521 B.n289 B.n72 585
R522 B.n291 B.n290 585
R523 B.n292 B.n71 585
R524 B.n294 B.n293 585
R525 B.n295 B.n70 585
R526 B.n297 B.n296 585
R527 B.n298 B.n69 585
R528 B.n300 B.n299 585
R529 B.n301 B.n68 585
R530 B.n303 B.n302 585
R531 B.n304 B.n67 585
R532 B.n306 B.n305 585
R533 B.n307 B.n66 585
R534 B.n309 B.n308 585
R535 B.n310 B.n65 585
R536 B.n312 B.n311 585
R537 B.n313 B.n64 585
R538 B.n315 B.n314 585
R539 B.n316 B.n63 585
R540 B.n318 B.n317 585
R541 B.n319 B.n62 585
R542 B.n321 B.n320 585
R543 B.n322 B.n61 585
R544 B.n324 B.n323 585
R545 B.n325 B.n60 585
R546 B.n327 B.n326 585
R547 B.n328 B.n59 585
R548 B.n330 B.n329 585
R549 B.n331 B.n58 585
R550 B.n333 B.n332 585
R551 B.n334 B.n57 585
R552 B.n336 B.n335 585
R553 B.n337 B.n56 585
R554 B.n339 B.n338 585
R555 B.n340 B.n55 585
R556 B.n342 B.n341 585
R557 B.n343 B.n54 585
R558 B.n345 B.n344 585
R559 B.n346 B.n53 585
R560 B.n348 B.n347 585
R561 B.n349 B.n52 585
R562 B.n351 B.n350 585
R563 B.n445 B.n16 585
R564 B.n444 B.n443 585
R565 B.n442 B.n17 585
R566 B.n441 B.n440 585
R567 B.n439 B.n18 585
R568 B.n438 B.n437 585
R569 B.n436 B.n19 585
R570 B.n435 B.n434 585
R571 B.n433 B.n20 585
R572 B.n432 B.n431 585
R573 B.n430 B.n21 585
R574 B.n429 B.n428 585
R575 B.n427 B.n22 585
R576 B.n426 B.n425 585
R577 B.n424 B.n23 585
R578 B.n423 B.n422 585
R579 B.n421 B.n24 585
R580 B.n420 B.n419 585
R581 B.n418 B.n25 585
R582 B.n417 B.n416 585
R583 B.n415 B.n26 585
R584 B.n414 B.n413 585
R585 B.n412 B.n27 585
R586 B.n411 B.n410 585
R587 B.n409 B.n28 585
R588 B.n408 B.n407 585
R589 B.n405 B.n29 585
R590 B.n404 B.n403 585
R591 B.n402 B.n32 585
R592 B.n401 B.n400 585
R593 B.n399 B.n33 585
R594 B.n398 B.n397 585
R595 B.n396 B.n34 585
R596 B.n395 B.n394 585
R597 B.n393 B.n35 585
R598 B.n392 B.n391 585
R599 B.n390 B.n389 585
R600 B.n388 B.n39 585
R601 B.n387 B.n386 585
R602 B.n385 B.n40 585
R603 B.n384 B.n383 585
R604 B.n382 B.n41 585
R605 B.n381 B.n380 585
R606 B.n379 B.n42 585
R607 B.n378 B.n377 585
R608 B.n376 B.n43 585
R609 B.n375 B.n374 585
R610 B.n373 B.n44 585
R611 B.n372 B.n371 585
R612 B.n370 B.n45 585
R613 B.n369 B.n368 585
R614 B.n367 B.n46 585
R615 B.n366 B.n365 585
R616 B.n364 B.n47 585
R617 B.n363 B.n362 585
R618 B.n361 B.n48 585
R619 B.n360 B.n359 585
R620 B.n358 B.n49 585
R621 B.n357 B.n356 585
R622 B.n355 B.n50 585
R623 B.n354 B.n353 585
R624 B.n352 B.n51 585
R625 B.n447 B.n446 585
R626 B.n448 B.n15 585
R627 B.n450 B.n449 585
R628 B.n451 B.n14 585
R629 B.n453 B.n452 585
R630 B.n454 B.n13 585
R631 B.n456 B.n455 585
R632 B.n457 B.n12 585
R633 B.n459 B.n458 585
R634 B.n460 B.n11 585
R635 B.n462 B.n461 585
R636 B.n463 B.n10 585
R637 B.n465 B.n464 585
R638 B.n466 B.n9 585
R639 B.n468 B.n467 585
R640 B.n469 B.n8 585
R641 B.n471 B.n470 585
R642 B.n472 B.n7 585
R643 B.n474 B.n473 585
R644 B.n475 B.n6 585
R645 B.n477 B.n476 585
R646 B.n478 B.n5 585
R647 B.n480 B.n479 585
R648 B.n481 B.n4 585
R649 B.n483 B.n482 585
R650 B.n484 B.n3 585
R651 B.n486 B.n485 585
R652 B.n487 B.n0 585
R653 B.n2 B.n1 585
R654 B.n128 B.n127 585
R655 B.n129 B.n126 585
R656 B.n131 B.n130 585
R657 B.n132 B.n125 585
R658 B.n134 B.n133 585
R659 B.n135 B.n124 585
R660 B.n137 B.n136 585
R661 B.n138 B.n123 585
R662 B.n140 B.n139 585
R663 B.n141 B.n122 585
R664 B.n143 B.n142 585
R665 B.n144 B.n121 585
R666 B.n146 B.n145 585
R667 B.n147 B.n120 585
R668 B.n149 B.n148 585
R669 B.n150 B.n119 585
R670 B.n152 B.n151 585
R671 B.n153 B.n118 585
R672 B.n155 B.n154 585
R673 B.n156 B.n117 585
R674 B.n158 B.n157 585
R675 B.n159 B.n116 585
R676 B.n161 B.n160 585
R677 B.n162 B.n115 585
R678 B.n164 B.n163 585
R679 B.n165 B.n114 585
R680 B.n167 B.n166 585
R681 B.n166 B.n113 545.355
R682 B.n265 B.n264 545.355
R683 B.n350 B.n51 545.355
R684 B.n446 B.n445 545.355
R685 B.n94 B.t10 350.199
R686 B.n36 B.t8 350.199
R687 B.n205 B.t4 350.199
R688 B.n30 B.t2 350.199
R689 B.n95 B.t11 282.32
R690 B.n37 B.t7 282.32
R691 B.n206 B.t5 282.32
R692 B.n31 B.t1 282.32
R693 B.n205 B.t3 260.392
R694 B.n94 B.t9 260.392
R695 B.n36 B.t6 260.392
R696 B.n30 B.t0 260.392
R697 B.n489 B.n488 256.663
R698 B.n488 B.n487 235.042
R699 B.n488 B.n2 235.042
R700 B.n170 B.n113 163.367
R701 B.n171 B.n170 163.367
R702 B.n172 B.n171 163.367
R703 B.n172 B.n111 163.367
R704 B.n176 B.n111 163.367
R705 B.n177 B.n176 163.367
R706 B.n178 B.n177 163.367
R707 B.n178 B.n109 163.367
R708 B.n182 B.n109 163.367
R709 B.n183 B.n182 163.367
R710 B.n184 B.n183 163.367
R711 B.n184 B.n107 163.367
R712 B.n188 B.n107 163.367
R713 B.n189 B.n188 163.367
R714 B.n190 B.n189 163.367
R715 B.n190 B.n105 163.367
R716 B.n194 B.n105 163.367
R717 B.n195 B.n194 163.367
R718 B.n196 B.n195 163.367
R719 B.n196 B.n103 163.367
R720 B.n200 B.n103 163.367
R721 B.n201 B.n200 163.367
R722 B.n202 B.n201 163.367
R723 B.n202 B.n101 163.367
R724 B.n209 B.n101 163.367
R725 B.n210 B.n209 163.367
R726 B.n211 B.n210 163.367
R727 B.n211 B.n99 163.367
R728 B.n215 B.n99 163.367
R729 B.n216 B.n215 163.367
R730 B.n217 B.n216 163.367
R731 B.n217 B.n97 163.367
R732 B.n221 B.n97 163.367
R733 B.n222 B.n221 163.367
R734 B.n223 B.n222 163.367
R735 B.n223 B.n93 163.367
R736 B.n228 B.n93 163.367
R737 B.n229 B.n228 163.367
R738 B.n230 B.n229 163.367
R739 B.n230 B.n91 163.367
R740 B.n234 B.n91 163.367
R741 B.n235 B.n234 163.367
R742 B.n236 B.n235 163.367
R743 B.n236 B.n89 163.367
R744 B.n240 B.n89 163.367
R745 B.n241 B.n240 163.367
R746 B.n242 B.n241 163.367
R747 B.n242 B.n87 163.367
R748 B.n246 B.n87 163.367
R749 B.n247 B.n246 163.367
R750 B.n248 B.n247 163.367
R751 B.n248 B.n85 163.367
R752 B.n252 B.n85 163.367
R753 B.n253 B.n252 163.367
R754 B.n254 B.n253 163.367
R755 B.n254 B.n83 163.367
R756 B.n258 B.n83 163.367
R757 B.n259 B.n258 163.367
R758 B.n260 B.n259 163.367
R759 B.n260 B.n81 163.367
R760 B.n264 B.n81 163.367
R761 B.n350 B.n349 163.367
R762 B.n349 B.n348 163.367
R763 B.n348 B.n53 163.367
R764 B.n344 B.n53 163.367
R765 B.n344 B.n343 163.367
R766 B.n343 B.n342 163.367
R767 B.n342 B.n55 163.367
R768 B.n338 B.n55 163.367
R769 B.n338 B.n337 163.367
R770 B.n337 B.n336 163.367
R771 B.n336 B.n57 163.367
R772 B.n332 B.n57 163.367
R773 B.n332 B.n331 163.367
R774 B.n331 B.n330 163.367
R775 B.n330 B.n59 163.367
R776 B.n326 B.n59 163.367
R777 B.n326 B.n325 163.367
R778 B.n325 B.n324 163.367
R779 B.n324 B.n61 163.367
R780 B.n320 B.n61 163.367
R781 B.n320 B.n319 163.367
R782 B.n319 B.n318 163.367
R783 B.n318 B.n63 163.367
R784 B.n314 B.n63 163.367
R785 B.n314 B.n313 163.367
R786 B.n313 B.n312 163.367
R787 B.n312 B.n65 163.367
R788 B.n308 B.n65 163.367
R789 B.n308 B.n307 163.367
R790 B.n307 B.n306 163.367
R791 B.n306 B.n67 163.367
R792 B.n302 B.n67 163.367
R793 B.n302 B.n301 163.367
R794 B.n301 B.n300 163.367
R795 B.n300 B.n69 163.367
R796 B.n296 B.n69 163.367
R797 B.n296 B.n295 163.367
R798 B.n295 B.n294 163.367
R799 B.n294 B.n71 163.367
R800 B.n290 B.n71 163.367
R801 B.n290 B.n289 163.367
R802 B.n289 B.n288 163.367
R803 B.n288 B.n73 163.367
R804 B.n284 B.n73 163.367
R805 B.n284 B.n283 163.367
R806 B.n283 B.n282 163.367
R807 B.n282 B.n75 163.367
R808 B.n278 B.n75 163.367
R809 B.n278 B.n277 163.367
R810 B.n277 B.n276 163.367
R811 B.n276 B.n77 163.367
R812 B.n272 B.n77 163.367
R813 B.n272 B.n271 163.367
R814 B.n271 B.n270 163.367
R815 B.n270 B.n79 163.367
R816 B.n266 B.n79 163.367
R817 B.n266 B.n265 163.367
R818 B.n445 B.n444 163.367
R819 B.n444 B.n17 163.367
R820 B.n440 B.n17 163.367
R821 B.n440 B.n439 163.367
R822 B.n439 B.n438 163.367
R823 B.n438 B.n19 163.367
R824 B.n434 B.n19 163.367
R825 B.n434 B.n433 163.367
R826 B.n433 B.n432 163.367
R827 B.n432 B.n21 163.367
R828 B.n428 B.n21 163.367
R829 B.n428 B.n427 163.367
R830 B.n427 B.n426 163.367
R831 B.n426 B.n23 163.367
R832 B.n422 B.n23 163.367
R833 B.n422 B.n421 163.367
R834 B.n421 B.n420 163.367
R835 B.n420 B.n25 163.367
R836 B.n416 B.n25 163.367
R837 B.n416 B.n415 163.367
R838 B.n415 B.n414 163.367
R839 B.n414 B.n27 163.367
R840 B.n410 B.n27 163.367
R841 B.n410 B.n409 163.367
R842 B.n409 B.n408 163.367
R843 B.n408 B.n29 163.367
R844 B.n403 B.n29 163.367
R845 B.n403 B.n402 163.367
R846 B.n402 B.n401 163.367
R847 B.n401 B.n33 163.367
R848 B.n397 B.n33 163.367
R849 B.n397 B.n396 163.367
R850 B.n396 B.n395 163.367
R851 B.n395 B.n35 163.367
R852 B.n391 B.n35 163.367
R853 B.n391 B.n390 163.367
R854 B.n390 B.n39 163.367
R855 B.n386 B.n39 163.367
R856 B.n386 B.n385 163.367
R857 B.n385 B.n384 163.367
R858 B.n384 B.n41 163.367
R859 B.n380 B.n41 163.367
R860 B.n380 B.n379 163.367
R861 B.n379 B.n378 163.367
R862 B.n378 B.n43 163.367
R863 B.n374 B.n43 163.367
R864 B.n374 B.n373 163.367
R865 B.n373 B.n372 163.367
R866 B.n372 B.n45 163.367
R867 B.n368 B.n45 163.367
R868 B.n368 B.n367 163.367
R869 B.n367 B.n366 163.367
R870 B.n366 B.n47 163.367
R871 B.n362 B.n47 163.367
R872 B.n362 B.n361 163.367
R873 B.n361 B.n360 163.367
R874 B.n360 B.n49 163.367
R875 B.n356 B.n49 163.367
R876 B.n356 B.n355 163.367
R877 B.n355 B.n354 163.367
R878 B.n354 B.n51 163.367
R879 B.n446 B.n15 163.367
R880 B.n450 B.n15 163.367
R881 B.n451 B.n450 163.367
R882 B.n452 B.n451 163.367
R883 B.n452 B.n13 163.367
R884 B.n456 B.n13 163.367
R885 B.n457 B.n456 163.367
R886 B.n458 B.n457 163.367
R887 B.n458 B.n11 163.367
R888 B.n462 B.n11 163.367
R889 B.n463 B.n462 163.367
R890 B.n464 B.n463 163.367
R891 B.n464 B.n9 163.367
R892 B.n468 B.n9 163.367
R893 B.n469 B.n468 163.367
R894 B.n470 B.n469 163.367
R895 B.n470 B.n7 163.367
R896 B.n474 B.n7 163.367
R897 B.n475 B.n474 163.367
R898 B.n476 B.n475 163.367
R899 B.n476 B.n5 163.367
R900 B.n480 B.n5 163.367
R901 B.n481 B.n480 163.367
R902 B.n482 B.n481 163.367
R903 B.n482 B.n3 163.367
R904 B.n486 B.n3 163.367
R905 B.n487 B.n486 163.367
R906 B.n128 B.n2 163.367
R907 B.n129 B.n128 163.367
R908 B.n130 B.n129 163.367
R909 B.n130 B.n125 163.367
R910 B.n134 B.n125 163.367
R911 B.n135 B.n134 163.367
R912 B.n136 B.n135 163.367
R913 B.n136 B.n123 163.367
R914 B.n140 B.n123 163.367
R915 B.n141 B.n140 163.367
R916 B.n142 B.n141 163.367
R917 B.n142 B.n121 163.367
R918 B.n146 B.n121 163.367
R919 B.n147 B.n146 163.367
R920 B.n148 B.n147 163.367
R921 B.n148 B.n119 163.367
R922 B.n152 B.n119 163.367
R923 B.n153 B.n152 163.367
R924 B.n154 B.n153 163.367
R925 B.n154 B.n117 163.367
R926 B.n158 B.n117 163.367
R927 B.n159 B.n158 163.367
R928 B.n160 B.n159 163.367
R929 B.n160 B.n115 163.367
R930 B.n164 B.n115 163.367
R931 B.n165 B.n164 163.367
R932 B.n166 B.n165 163.367
R933 B.n206 B.n205 67.8793
R934 B.n95 B.n94 67.8793
R935 B.n37 B.n36 67.8793
R936 B.n31 B.n30 67.8793
R937 B.n207 B.n206 59.5399
R938 B.n225 B.n95 59.5399
R939 B.n38 B.n37 59.5399
R940 B.n406 B.n31 59.5399
R941 B.n263 B.n80 35.4346
R942 B.n447 B.n16 35.4346
R943 B.n352 B.n351 35.4346
R944 B.n168 B.n167 35.4346
R945 B B.n489 18.0485
R946 B.n448 B.n447 10.6151
R947 B.n449 B.n448 10.6151
R948 B.n449 B.n14 10.6151
R949 B.n453 B.n14 10.6151
R950 B.n454 B.n453 10.6151
R951 B.n455 B.n454 10.6151
R952 B.n455 B.n12 10.6151
R953 B.n459 B.n12 10.6151
R954 B.n460 B.n459 10.6151
R955 B.n461 B.n460 10.6151
R956 B.n461 B.n10 10.6151
R957 B.n465 B.n10 10.6151
R958 B.n466 B.n465 10.6151
R959 B.n467 B.n466 10.6151
R960 B.n467 B.n8 10.6151
R961 B.n471 B.n8 10.6151
R962 B.n472 B.n471 10.6151
R963 B.n473 B.n472 10.6151
R964 B.n473 B.n6 10.6151
R965 B.n477 B.n6 10.6151
R966 B.n478 B.n477 10.6151
R967 B.n479 B.n478 10.6151
R968 B.n479 B.n4 10.6151
R969 B.n483 B.n4 10.6151
R970 B.n484 B.n483 10.6151
R971 B.n485 B.n484 10.6151
R972 B.n485 B.n0 10.6151
R973 B.n443 B.n16 10.6151
R974 B.n443 B.n442 10.6151
R975 B.n442 B.n441 10.6151
R976 B.n441 B.n18 10.6151
R977 B.n437 B.n18 10.6151
R978 B.n437 B.n436 10.6151
R979 B.n436 B.n435 10.6151
R980 B.n435 B.n20 10.6151
R981 B.n431 B.n20 10.6151
R982 B.n431 B.n430 10.6151
R983 B.n430 B.n429 10.6151
R984 B.n429 B.n22 10.6151
R985 B.n425 B.n22 10.6151
R986 B.n425 B.n424 10.6151
R987 B.n424 B.n423 10.6151
R988 B.n423 B.n24 10.6151
R989 B.n419 B.n24 10.6151
R990 B.n419 B.n418 10.6151
R991 B.n418 B.n417 10.6151
R992 B.n417 B.n26 10.6151
R993 B.n413 B.n26 10.6151
R994 B.n413 B.n412 10.6151
R995 B.n412 B.n411 10.6151
R996 B.n411 B.n28 10.6151
R997 B.n407 B.n28 10.6151
R998 B.n405 B.n404 10.6151
R999 B.n404 B.n32 10.6151
R1000 B.n400 B.n32 10.6151
R1001 B.n400 B.n399 10.6151
R1002 B.n399 B.n398 10.6151
R1003 B.n398 B.n34 10.6151
R1004 B.n394 B.n34 10.6151
R1005 B.n394 B.n393 10.6151
R1006 B.n393 B.n392 10.6151
R1007 B.n389 B.n388 10.6151
R1008 B.n388 B.n387 10.6151
R1009 B.n387 B.n40 10.6151
R1010 B.n383 B.n40 10.6151
R1011 B.n383 B.n382 10.6151
R1012 B.n382 B.n381 10.6151
R1013 B.n381 B.n42 10.6151
R1014 B.n377 B.n42 10.6151
R1015 B.n377 B.n376 10.6151
R1016 B.n376 B.n375 10.6151
R1017 B.n375 B.n44 10.6151
R1018 B.n371 B.n44 10.6151
R1019 B.n371 B.n370 10.6151
R1020 B.n370 B.n369 10.6151
R1021 B.n369 B.n46 10.6151
R1022 B.n365 B.n46 10.6151
R1023 B.n365 B.n364 10.6151
R1024 B.n364 B.n363 10.6151
R1025 B.n363 B.n48 10.6151
R1026 B.n359 B.n48 10.6151
R1027 B.n359 B.n358 10.6151
R1028 B.n358 B.n357 10.6151
R1029 B.n357 B.n50 10.6151
R1030 B.n353 B.n50 10.6151
R1031 B.n353 B.n352 10.6151
R1032 B.n351 B.n52 10.6151
R1033 B.n347 B.n52 10.6151
R1034 B.n347 B.n346 10.6151
R1035 B.n346 B.n345 10.6151
R1036 B.n345 B.n54 10.6151
R1037 B.n341 B.n54 10.6151
R1038 B.n341 B.n340 10.6151
R1039 B.n340 B.n339 10.6151
R1040 B.n339 B.n56 10.6151
R1041 B.n335 B.n56 10.6151
R1042 B.n335 B.n334 10.6151
R1043 B.n334 B.n333 10.6151
R1044 B.n333 B.n58 10.6151
R1045 B.n329 B.n58 10.6151
R1046 B.n329 B.n328 10.6151
R1047 B.n328 B.n327 10.6151
R1048 B.n327 B.n60 10.6151
R1049 B.n323 B.n60 10.6151
R1050 B.n323 B.n322 10.6151
R1051 B.n322 B.n321 10.6151
R1052 B.n321 B.n62 10.6151
R1053 B.n317 B.n62 10.6151
R1054 B.n317 B.n316 10.6151
R1055 B.n316 B.n315 10.6151
R1056 B.n315 B.n64 10.6151
R1057 B.n311 B.n64 10.6151
R1058 B.n311 B.n310 10.6151
R1059 B.n310 B.n309 10.6151
R1060 B.n309 B.n66 10.6151
R1061 B.n305 B.n66 10.6151
R1062 B.n305 B.n304 10.6151
R1063 B.n304 B.n303 10.6151
R1064 B.n303 B.n68 10.6151
R1065 B.n299 B.n68 10.6151
R1066 B.n299 B.n298 10.6151
R1067 B.n298 B.n297 10.6151
R1068 B.n297 B.n70 10.6151
R1069 B.n293 B.n70 10.6151
R1070 B.n293 B.n292 10.6151
R1071 B.n292 B.n291 10.6151
R1072 B.n291 B.n72 10.6151
R1073 B.n287 B.n72 10.6151
R1074 B.n287 B.n286 10.6151
R1075 B.n286 B.n285 10.6151
R1076 B.n285 B.n74 10.6151
R1077 B.n281 B.n74 10.6151
R1078 B.n281 B.n280 10.6151
R1079 B.n280 B.n279 10.6151
R1080 B.n279 B.n76 10.6151
R1081 B.n275 B.n76 10.6151
R1082 B.n275 B.n274 10.6151
R1083 B.n274 B.n273 10.6151
R1084 B.n273 B.n78 10.6151
R1085 B.n269 B.n78 10.6151
R1086 B.n269 B.n268 10.6151
R1087 B.n268 B.n267 10.6151
R1088 B.n267 B.n80 10.6151
R1089 B.n127 B.n1 10.6151
R1090 B.n127 B.n126 10.6151
R1091 B.n131 B.n126 10.6151
R1092 B.n132 B.n131 10.6151
R1093 B.n133 B.n132 10.6151
R1094 B.n133 B.n124 10.6151
R1095 B.n137 B.n124 10.6151
R1096 B.n138 B.n137 10.6151
R1097 B.n139 B.n138 10.6151
R1098 B.n139 B.n122 10.6151
R1099 B.n143 B.n122 10.6151
R1100 B.n144 B.n143 10.6151
R1101 B.n145 B.n144 10.6151
R1102 B.n145 B.n120 10.6151
R1103 B.n149 B.n120 10.6151
R1104 B.n150 B.n149 10.6151
R1105 B.n151 B.n150 10.6151
R1106 B.n151 B.n118 10.6151
R1107 B.n155 B.n118 10.6151
R1108 B.n156 B.n155 10.6151
R1109 B.n157 B.n156 10.6151
R1110 B.n157 B.n116 10.6151
R1111 B.n161 B.n116 10.6151
R1112 B.n162 B.n161 10.6151
R1113 B.n163 B.n162 10.6151
R1114 B.n163 B.n114 10.6151
R1115 B.n167 B.n114 10.6151
R1116 B.n169 B.n168 10.6151
R1117 B.n169 B.n112 10.6151
R1118 B.n173 B.n112 10.6151
R1119 B.n174 B.n173 10.6151
R1120 B.n175 B.n174 10.6151
R1121 B.n175 B.n110 10.6151
R1122 B.n179 B.n110 10.6151
R1123 B.n180 B.n179 10.6151
R1124 B.n181 B.n180 10.6151
R1125 B.n181 B.n108 10.6151
R1126 B.n185 B.n108 10.6151
R1127 B.n186 B.n185 10.6151
R1128 B.n187 B.n186 10.6151
R1129 B.n187 B.n106 10.6151
R1130 B.n191 B.n106 10.6151
R1131 B.n192 B.n191 10.6151
R1132 B.n193 B.n192 10.6151
R1133 B.n193 B.n104 10.6151
R1134 B.n197 B.n104 10.6151
R1135 B.n198 B.n197 10.6151
R1136 B.n199 B.n198 10.6151
R1137 B.n199 B.n102 10.6151
R1138 B.n203 B.n102 10.6151
R1139 B.n204 B.n203 10.6151
R1140 B.n208 B.n204 10.6151
R1141 B.n212 B.n100 10.6151
R1142 B.n213 B.n212 10.6151
R1143 B.n214 B.n213 10.6151
R1144 B.n214 B.n98 10.6151
R1145 B.n218 B.n98 10.6151
R1146 B.n219 B.n218 10.6151
R1147 B.n220 B.n219 10.6151
R1148 B.n220 B.n96 10.6151
R1149 B.n224 B.n96 10.6151
R1150 B.n227 B.n226 10.6151
R1151 B.n227 B.n92 10.6151
R1152 B.n231 B.n92 10.6151
R1153 B.n232 B.n231 10.6151
R1154 B.n233 B.n232 10.6151
R1155 B.n233 B.n90 10.6151
R1156 B.n237 B.n90 10.6151
R1157 B.n238 B.n237 10.6151
R1158 B.n239 B.n238 10.6151
R1159 B.n239 B.n88 10.6151
R1160 B.n243 B.n88 10.6151
R1161 B.n244 B.n243 10.6151
R1162 B.n245 B.n244 10.6151
R1163 B.n245 B.n86 10.6151
R1164 B.n249 B.n86 10.6151
R1165 B.n250 B.n249 10.6151
R1166 B.n251 B.n250 10.6151
R1167 B.n251 B.n84 10.6151
R1168 B.n255 B.n84 10.6151
R1169 B.n256 B.n255 10.6151
R1170 B.n257 B.n256 10.6151
R1171 B.n257 B.n82 10.6151
R1172 B.n261 B.n82 10.6151
R1173 B.n262 B.n261 10.6151
R1174 B.n263 B.n262 10.6151
R1175 B.n407 B.n406 9.36635
R1176 B.n389 B.n38 9.36635
R1177 B.n208 B.n207 9.36635
R1178 B.n226 B.n225 9.36635
R1179 B.n489 B.n0 8.11757
R1180 B.n489 B.n1 8.11757
R1181 B.n406 B.n405 1.24928
R1182 B.n392 B.n38 1.24928
R1183 B.n207 B.n100 1.24928
R1184 B.n225 B.n224 1.24928
C0 VDD2 VDD1 0.743463f
C1 VN VP 4.76235f
C2 VP VTAIL 1.78228f
C3 VP VDD1 1.93328f
C4 VN B 1.08288f
C5 VN w_n2370_n2326# 3.24214f
C6 B VTAIL 2.66164f
C7 VP VDD2 0.356653f
C8 VTAIL w_n2370_n2326# 2.04012f
C9 B VDD1 1.36541f
C10 w_n2370_n2326# VDD1 1.48685f
C11 B VDD2 1.40057f
C12 VDD2 w_n2370_n2326# 1.51977f
C13 B VP 1.58351f
C14 VP w_n2370_n2326# 3.54526f
C15 VN VTAIL 1.76809f
C16 VN VDD1 0.148384f
C17 VTAIL VDD1 3.8352f
C18 B w_n2370_n2326# 7.96929f
C19 VN VDD2 1.72652f
C20 VDD2 VTAIL 3.89115f
C21 VDD2 VSUBS 0.730579f
C22 VDD1 VSUBS 2.512518f
C23 VTAIL VSUBS 0.614118f
C24 VN VSUBS 5.65446f
C25 VP VSUBS 1.54105f
C26 B VSUBS 3.887442f
C27 w_n2370_n2326# VSUBS 68.6257f
C28 B.n0 VSUBS 0.006464f
C29 B.n1 VSUBS 0.006464f
C30 B.n2 VSUBS 0.00956f
C31 B.n3 VSUBS 0.007326f
C32 B.n4 VSUBS 0.007326f
C33 B.n5 VSUBS 0.007326f
C34 B.n6 VSUBS 0.007326f
C35 B.n7 VSUBS 0.007326f
C36 B.n8 VSUBS 0.007326f
C37 B.n9 VSUBS 0.007326f
C38 B.n10 VSUBS 0.007326f
C39 B.n11 VSUBS 0.007326f
C40 B.n12 VSUBS 0.007326f
C41 B.n13 VSUBS 0.007326f
C42 B.n14 VSUBS 0.007326f
C43 B.n15 VSUBS 0.007326f
C44 B.n16 VSUBS 0.018556f
C45 B.n17 VSUBS 0.007326f
C46 B.n18 VSUBS 0.007326f
C47 B.n19 VSUBS 0.007326f
C48 B.n20 VSUBS 0.007326f
C49 B.n21 VSUBS 0.007326f
C50 B.n22 VSUBS 0.007326f
C51 B.n23 VSUBS 0.007326f
C52 B.n24 VSUBS 0.007326f
C53 B.n25 VSUBS 0.007326f
C54 B.n26 VSUBS 0.007326f
C55 B.n27 VSUBS 0.007326f
C56 B.n28 VSUBS 0.007326f
C57 B.n29 VSUBS 0.007326f
C58 B.t1 VSUBS 0.108709f
C59 B.t2 VSUBS 0.141772f
C60 B.t0 VSUBS 1.06952f
C61 B.n30 VSUBS 0.235201f
C62 B.n31 VSUBS 0.181025f
C63 B.n32 VSUBS 0.007326f
C64 B.n33 VSUBS 0.007326f
C65 B.n34 VSUBS 0.007326f
C66 B.n35 VSUBS 0.007326f
C67 B.t7 VSUBS 0.108711f
C68 B.t8 VSUBS 0.141774f
C69 B.t6 VSUBS 1.06952f
C70 B.n36 VSUBS 0.2352f
C71 B.n37 VSUBS 0.181023f
C72 B.n38 VSUBS 0.016973f
C73 B.n39 VSUBS 0.007326f
C74 B.n40 VSUBS 0.007326f
C75 B.n41 VSUBS 0.007326f
C76 B.n42 VSUBS 0.007326f
C77 B.n43 VSUBS 0.007326f
C78 B.n44 VSUBS 0.007326f
C79 B.n45 VSUBS 0.007326f
C80 B.n46 VSUBS 0.007326f
C81 B.n47 VSUBS 0.007326f
C82 B.n48 VSUBS 0.007326f
C83 B.n49 VSUBS 0.007326f
C84 B.n50 VSUBS 0.007326f
C85 B.n51 VSUBS 0.018556f
C86 B.n52 VSUBS 0.007326f
C87 B.n53 VSUBS 0.007326f
C88 B.n54 VSUBS 0.007326f
C89 B.n55 VSUBS 0.007326f
C90 B.n56 VSUBS 0.007326f
C91 B.n57 VSUBS 0.007326f
C92 B.n58 VSUBS 0.007326f
C93 B.n59 VSUBS 0.007326f
C94 B.n60 VSUBS 0.007326f
C95 B.n61 VSUBS 0.007326f
C96 B.n62 VSUBS 0.007326f
C97 B.n63 VSUBS 0.007326f
C98 B.n64 VSUBS 0.007326f
C99 B.n65 VSUBS 0.007326f
C100 B.n66 VSUBS 0.007326f
C101 B.n67 VSUBS 0.007326f
C102 B.n68 VSUBS 0.007326f
C103 B.n69 VSUBS 0.007326f
C104 B.n70 VSUBS 0.007326f
C105 B.n71 VSUBS 0.007326f
C106 B.n72 VSUBS 0.007326f
C107 B.n73 VSUBS 0.007326f
C108 B.n74 VSUBS 0.007326f
C109 B.n75 VSUBS 0.007326f
C110 B.n76 VSUBS 0.007326f
C111 B.n77 VSUBS 0.007326f
C112 B.n78 VSUBS 0.007326f
C113 B.n79 VSUBS 0.007326f
C114 B.n80 VSUBS 0.018439f
C115 B.n81 VSUBS 0.007326f
C116 B.n82 VSUBS 0.007326f
C117 B.n83 VSUBS 0.007326f
C118 B.n84 VSUBS 0.007326f
C119 B.n85 VSUBS 0.007326f
C120 B.n86 VSUBS 0.007326f
C121 B.n87 VSUBS 0.007326f
C122 B.n88 VSUBS 0.007326f
C123 B.n89 VSUBS 0.007326f
C124 B.n90 VSUBS 0.007326f
C125 B.n91 VSUBS 0.007326f
C126 B.n92 VSUBS 0.007326f
C127 B.n93 VSUBS 0.007326f
C128 B.t11 VSUBS 0.108711f
C129 B.t10 VSUBS 0.141774f
C130 B.t9 VSUBS 1.06952f
C131 B.n94 VSUBS 0.2352f
C132 B.n95 VSUBS 0.181023f
C133 B.n96 VSUBS 0.007326f
C134 B.n97 VSUBS 0.007326f
C135 B.n98 VSUBS 0.007326f
C136 B.n99 VSUBS 0.007326f
C137 B.n100 VSUBS 0.004094f
C138 B.n101 VSUBS 0.007326f
C139 B.n102 VSUBS 0.007326f
C140 B.n103 VSUBS 0.007326f
C141 B.n104 VSUBS 0.007326f
C142 B.n105 VSUBS 0.007326f
C143 B.n106 VSUBS 0.007326f
C144 B.n107 VSUBS 0.007326f
C145 B.n108 VSUBS 0.007326f
C146 B.n109 VSUBS 0.007326f
C147 B.n110 VSUBS 0.007326f
C148 B.n111 VSUBS 0.007326f
C149 B.n112 VSUBS 0.007326f
C150 B.n113 VSUBS 0.018556f
C151 B.n114 VSUBS 0.007326f
C152 B.n115 VSUBS 0.007326f
C153 B.n116 VSUBS 0.007326f
C154 B.n117 VSUBS 0.007326f
C155 B.n118 VSUBS 0.007326f
C156 B.n119 VSUBS 0.007326f
C157 B.n120 VSUBS 0.007326f
C158 B.n121 VSUBS 0.007326f
C159 B.n122 VSUBS 0.007326f
C160 B.n123 VSUBS 0.007326f
C161 B.n124 VSUBS 0.007326f
C162 B.n125 VSUBS 0.007326f
C163 B.n126 VSUBS 0.007326f
C164 B.n127 VSUBS 0.007326f
C165 B.n128 VSUBS 0.007326f
C166 B.n129 VSUBS 0.007326f
C167 B.n130 VSUBS 0.007326f
C168 B.n131 VSUBS 0.007326f
C169 B.n132 VSUBS 0.007326f
C170 B.n133 VSUBS 0.007326f
C171 B.n134 VSUBS 0.007326f
C172 B.n135 VSUBS 0.007326f
C173 B.n136 VSUBS 0.007326f
C174 B.n137 VSUBS 0.007326f
C175 B.n138 VSUBS 0.007326f
C176 B.n139 VSUBS 0.007326f
C177 B.n140 VSUBS 0.007326f
C178 B.n141 VSUBS 0.007326f
C179 B.n142 VSUBS 0.007326f
C180 B.n143 VSUBS 0.007326f
C181 B.n144 VSUBS 0.007326f
C182 B.n145 VSUBS 0.007326f
C183 B.n146 VSUBS 0.007326f
C184 B.n147 VSUBS 0.007326f
C185 B.n148 VSUBS 0.007326f
C186 B.n149 VSUBS 0.007326f
C187 B.n150 VSUBS 0.007326f
C188 B.n151 VSUBS 0.007326f
C189 B.n152 VSUBS 0.007326f
C190 B.n153 VSUBS 0.007326f
C191 B.n154 VSUBS 0.007326f
C192 B.n155 VSUBS 0.007326f
C193 B.n156 VSUBS 0.007326f
C194 B.n157 VSUBS 0.007326f
C195 B.n158 VSUBS 0.007326f
C196 B.n159 VSUBS 0.007326f
C197 B.n160 VSUBS 0.007326f
C198 B.n161 VSUBS 0.007326f
C199 B.n162 VSUBS 0.007326f
C200 B.n163 VSUBS 0.007326f
C201 B.n164 VSUBS 0.007326f
C202 B.n165 VSUBS 0.007326f
C203 B.n166 VSUBS 0.017642f
C204 B.n167 VSUBS 0.017642f
C205 B.n168 VSUBS 0.018556f
C206 B.n169 VSUBS 0.007326f
C207 B.n170 VSUBS 0.007326f
C208 B.n171 VSUBS 0.007326f
C209 B.n172 VSUBS 0.007326f
C210 B.n173 VSUBS 0.007326f
C211 B.n174 VSUBS 0.007326f
C212 B.n175 VSUBS 0.007326f
C213 B.n176 VSUBS 0.007326f
C214 B.n177 VSUBS 0.007326f
C215 B.n178 VSUBS 0.007326f
C216 B.n179 VSUBS 0.007326f
C217 B.n180 VSUBS 0.007326f
C218 B.n181 VSUBS 0.007326f
C219 B.n182 VSUBS 0.007326f
C220 B.n183 VSUBS 0.007326f
C221 B.n184 VSUBS 0.007326f
C222 B.n185 VSUBS 0.007326f
C223 B.n186 VSUBS 0.007326f
C224 B.n187 VSUBS 0.007326f
C225 B.n188 VSUBS 0.007326f
C226 B.n189 VSUBS 0.007326f
C227 B.n190 VSUBS 0.007326f
C228 B.n191 VSUBS 0.007326f
C229 B.n192 VSUBS 0.007326f
C230 B.n193 VSUBS 0.007326f
C231 B.n194 VSUBS 0.007326f
C232 B.n195 VSUBS 0.007326f
C233 B.n196 VSUBS 0.007326f
C234 B.n197 VSUBS 0.007326f
C235 B.n198 VSUBS 0.007326f
C236 B.n199 VSUBS 0.007326f
C237 B.n200 VSUBS 0.007326f
C238 B.n201 VSUBS 0.007326f
C239 B.n202 VSUBS 0.007326f
C240 B.n203 VSUBS 0.007326f
C241 B.n204 VSUBS 0.007326f
C242 B.t5 VSUBS 0.108709f
C243 B.t4 VSUBS 0.141772f
C244 B.t3 VSUBS 1.06952f
C245 B.n205 VSUBS 0.235201f
C246 B.n206 VSUBS 0.181025f
C247 B.n207 VSUBS 0.016973f
C248 B.n208 VSUBS 0.006895f
C249 B.n209 VSUBS 0.007326f
C250 B.n210 VSUBS 0.007326f
C251 B.n211 VSUBS 0.007326f
C252 B.n212 VSUBS 0.007326f
C253 B.n213 VSUBS 0.007326f
C254 B.n214 VSUBS 0.007326f
C255 B.n215 VSUBS 0.007326f
C256 B.n216 VSUBS 0.007326f
C257 B.n217 VSUBS 0.007326f
C258 B.n218 VSUBS 0.007326f
C259 B.n219 VSUBS 0.007326f
C260 B.n220 VSUBS 0.007326f
C261 B.n221 VSUBS 0.007326f
C262 B.n222 VSUBS 0.007326f
C263 B.n223 VSUBS 0.007326f
C264 B.n224 VSUBS 0.004094f
C265 B.n225 VSUBS 0.016973f
C266 B.n226 VSUBS 0.006895f
C267 B.n227 VSUBS 0.007326f
C268 B.n228 VSUBS 0.007326f
C269 B.n229 VSUBS 0.007326f
C270 B.n230 VSUBS 0.007326f
C271 B.n231 VSUBS 0.007326f
C272 B.n232 VSUBS 0.007326f
C273 B.n233 VSUBS 0.007326f
C274 B.n234 VSUBS 0.007326f
C275 B.n235 VSUBS 0.007326f
C276 B.n236 VSUBS 0.007326f
C277 B.n237 VSUBS 0.007326f
C278 B.n238 VSUBS 0.007326f
C279 B.n239 VSUBS 0.007326f
C280 B.n240 VSUBS 0.007326f
C281 B.n241 VSUBS 0.007326f
C282 B.n242 VSUBS 0.007326f
C283 B.n243 VSUBS 0.007326f
C284 B.n244 VSUBS 0.007326f
C285 B.n245 VSUBS 0.007326f
C286 B.n246 VSUBS 0.007326f
C287 B.n247 VSUBS 0.007326f
C288 B.n248 VSUBS 0.007326f
C289 B.n249 VSUBS 0.007326f
C290 B.n250 VSUBS 0.007326f
C291 B.n251 VSUBS 0.007326f
C292 B.n252 VSUBS 0.007326f
C293 B.n253 VSUBS 0.007326f
C294 B.n254 VSUBS 0.007326f
C295 B.n255 VSUBS 0.007326f
C296 B.n256 VSUBS 0.007326f
C297 B.n257 VSUBS 0.007326f
C298 B.n258 VSUBS 0.007326f
C299 B.n259 VSUBS 0.007326f
C300 B.n260 VSUBS 0.007326f
C301 B.n261 VSUBS 0.007326f
C302 B.n262 VSUBS 0.007326f
C303 B.n263 VSUBS 0.017758f
C304 B.n264 VSUBS 0.018556f
C305 B.n265 VSUBS 0.017642f
C306 B.n266 VSUBS 0.007326f
C307 B.n267 VSUBS 0.007326f
C308 B.n268 VSUBS 0.007326f
C309 B.n269 VSUBS 0.007326f
C310 B.n270 VSUBS 0.007326f
C311 B.n271 VSUBS 0.007326f
C312 B.n272 VSUBS 0.007326f
C313 B.n273 VSUBS 0.007326f
C314 B.n274 VSUBS 0.007326f
C315 B.n275 VSUBS 0.007326f
C316 B.n276 VSUBS 0.007326f
C317 B.n277 VSUBS 0.007326f
C318 B.n278 VSUBS 0.007326f
C319 B.n279 VSUBS 0.007326f
C320 B.n280 VSUBS 0.007326f
C321 B.n281 VSUBS 0.007326f
C322 B.n282 VSUBS 0.007326f
C323 B.n283 VSUBS 0.007326f
C324 B.n284 VSUBS 0.007326f
C325 B.n285 VSUBS 0.007326f
C326 B.n286 VSUBS 0.007326f
C327 B.n287 VSUBS 0.007326f
C328 B.n288 VSUBS 0.007326f
C329 B.n289 VSUBS 0.007326f
C330 B.n290 VSUBS 0.007326f
C331 B.n291 VSUBS 0.007326f
C332 B.n292 VSUBS 0.007326f
C333 B.n293 VSUBS 0.007326f
C334 B.n294 VSUBS 0.007326f
C335 B.n295 VSUBS 0.007326f
C336 B.n296 VSUBS 0.007326f
C337 B.n297 VSUBS 0.007326f
C338 B.n298 VSUBS 0.007326f
C339 B.n299 VSUBS 0.007326f
C340 B.n300 VSUBS 0.007326f
C341 B.n301 VSUBS 0.007326f
C342 B.n302 VSUBS 0.007326f
C343 B.n303 VSUBS 0.007326f
C344 B.n304 VSUBS 0.007326f
C345 B.n305 VSUBS 0.007326f
C346 B.n306 VSUBS 0.007326f
C347 B.n307 VSUBS 0.007326f
C348 B.n308 VSUBS 0.007326f
C349 B.n309 VSUBS 0.007326f
C350 B.n310 VSUBS 0.007326f
C351 B.n311 VSUBS 0.007326f
C352 B.n312 VSUBS 0.007326f
C353 B.n313 VSUBS 0.007326f
C354 B.n314 VSUBS 0.007326f
C355 B.n315 VSUBS 0.007326f
C356 B.n316 VSUBS 0.007326f
C357 B.n317 VSUBS 0.007326f
C358 B.n318 VSUBS 0.007326f
C359 B.n319 VSUBS 0.007326f
C360 B.n320 VSUBS 0.007326f
C361 B.n321 VSUBS 0.007326f
C362 B.n322 VSUBS 0.007326f
C363 B.n323 VSUBS 0.007326f
C364 B.n324 VSUBS 0.007326f
C365 B.n325 VSUBS 0.007326f
C366 B.n326 VSUBS 0.007326f
C367 B.n327 VSUBS 0.007326f
C368 B.n328 VSUBS 0.007326f
C369 B.n329 VSUBS 0.007326f
C370 B.n330 VSUBS 0.007326f
C371 B.n331 VSUBS 0.007326f
C372 B.n332 VSUBS 0.007326f
C373 B.n333 VSUBS 0.007326f
C374 B.n334 VSUBS 0.007326f
C375 B.n335 VSUBS 0.007326f
C376 B.n336 VSUBS 0.007326f
C377 B.n337 VSUBS 0.007326f
C378 B.n338 VSUBS 0.007326f
C379 B.n339 VSUBS 0.007326f
C380 B.n340 VSUBS 0.007326f
C381 B.n341 VSUBS 0.007326f
C382 B.n342 VSUBS 0.007326f
C383 B.n343 VSUBS 0.007326f
C384 B.n344 VSUBS 0.007326f
C385 B.n345 VSUBS 0.007326f
C386 B.n346 VSUBS 0.007326f
C387 B.n347 VSUBS 0.007326f
C388 B.n348 VSUBS 0.007326f
C389 B.n349 VSUBS 0.007326f
C390 B.n350 VSUBS 0.017642f
C391 B.n351 VSUBS 0.017642f
C392 B.n352 VSUBS 0.018556f
C393 B.n353 VSUBS 0.007326f
C394 B.n354 VSUBS 0.007326f
C395 B.n355 VSUBS 0.007326f
C396 B.n356 VSUBS 0.007326f
C397 B.n357 VSUBS 0.007326f
C398 B.n358 VSUBS 0.007326f
C399 B.n359 VSUBS 0.007326f
C400 B.n360 VSUBS 0.007326f
C401 B.n361 VSUBS 0.007326f
C402 B.n362 VSUBS 0.007326f
C403 B.n363 VSUBS 0.007326f
C404 B.n364 VSUBS 0.007326f
C405 B.n365 VSUBS 0.007326f
C406 B.n366 VSUBS 0.007326f
C407 B.n367 VSUBS 0.007326f
C408 B.n368 VSUBS 0.007326f
C409 B.n369 VSUBS 0.007326f
C410 B.n370 VSUBS 0.007326f
C411 B.n371 VSUBS 0.007326f
C412 B.n372 VSUBS 0.007326f
C413 B.n373 VSUBS 0.007326f
C414 B.n374 VSUBS 0.007326f
C415 B.n375 VSUBS 0.007326f
C416 B.n376 VSUBS 0.007326f
C417 B.n377 VSUBS 0.007326f
C418 B.n378 VSUBS 0.007326f
C419 B.n379 VSUBS 0.007326f
C420 B.n380 VSUBS 0.007326f
C421 B.n381 VSUBS 0.007326f
C422 B.n382 VSUBS 0.007326f
C423 B.n383 VSUBS 0.007326f
C424 B.n384 VSUBS 0.007326f
C425 B.n385 VSUBS 0.007326f
C426 B.n386 VSUBS 0.007326f
C427 B.n387 VSUBS 0.007326f
C428 B.n388 VSUBS 0.007326f
C429 B.n389 VSUBS 0.006895f
C430 B.n390 VSUBS 0.007326f
C431 B.n391 VSUBS 0.007326f
C432 B.n392 VSUBS 0.004094f
C433 B.n393 VSUBS 0.007326f
C434 B.n394 VSUBS 0.007326f
C435 B.n395 VSUBS 0.007326f
C436 B.n396 VSUBS 0.007326f
C437 B.n397 VSUBS 0.007326f
C438 B.n398 VSUBS 0.007326f
C439 B.n399 VSUBS 0.007326f
C440 B.n400 VSUBS 0.007326f
C441 B.n401 VSUBS 0.007326f
C442 B.n402 VSUBS 0.007326f
C443 B.n403 VSUBS 0.007326f
C444 B.n404 VSUBS 0.007326f
C445 B.n405 VSUBS 0.004094f
C446 B.n406 VSUBS 0.016973f
C447 B.n407 VSUBS 0.006895f
C448 B.n408 VSUBS 0.007326f
C449 B.n409 VSUBS 0.007326f
C450 B.n410 VSUBS 0.007326f
C451 B.n411 VSUBS 0.007326f
C452 B.n412 VSUBS 0.007326f
C453 B.n413 VSUBS 0.007326f
C454 B.n414 VSUBS 0.007326f
C455 B.n415 VSUBS 0.007326f
C456 B.n416 VSUBS 0.007326f
C457 B.n417 VSUBS 0.007326f
C458 B.n418 VSUBS 0.007326f
C459 B.n419 VSUBS 0.007326f
C460 B.n420 VSUBS 0.007326f
C461 B.n421 VSUBS 0.007326f
C462 B.n422 VSUBS 0.007326f
C463 B.n423 VSUBS 0.007326f
C464 B.n424 VSUBS 0.007326f
C465 B.n425 VSUBS 0.007326f
C466 B.n426 VSUBS 0.007326f
C467 B.n427 VSUBS 0.007326f
C468 B.n428 VSUBS 0.007326f
C469 B.n429 VSUBS 0.007326f
C470 B.n430 VSUBS 0.007326f
C471 B.n431 VSUBS 0.007326f
C472 B.n432 VSUBS 0.007326f
C473 B.n433 VSUBS 0.007326f
C474 B.n434 VSUBS 0.007326f
C475 B.n435 VSUBS 0.007326f
C476 B.n436 VSUBS 0.007326f
C477 B.n437 VSUBS 0.007326f
C478 B.n438 VSUBS 0.007326f
C479 B.n439 VSUBS 0.007326f
C480 B.n440 VSUBS 0.007326f
C481 B.n441 VSUBS 0.007326f
C482 B.n442 VSUBS 0.007326f
C483 B.n443 VSUBS 0.007326f
C484 B.n444 VSUBS 0.007326f
C485 B.n445 VSUBS 0.018556f
C486 B.n446 VSUBS 0.017642f
C487 B.n447 VSUBS 0.017642f
C488 B.n448 VSUBS 0.007326f
C489 B.n449 VSUBS 0.007326f
C490 B.n450 VSUBS 0.007326f
C491 B.n451 VSUBS 0.007326f
C492 B.n452 VSUBS 0.007326f
C493 B.n453 VSUBS 0.007326f
C494 B.n454 VSUBS 0.007326f
C495 B.n455 VSUBS 0.007326f
C496 B.n456 VSUBS 0.007326f
C497 B.n457 VSUBS 0.007326f
C498 B.n458 VSUBS 0.007326f
C499 B.n459 VSUBS 0.007326f
C500 B.n460 VSUBS 0.007326f
C501 B.n461 VSUBS 0.007326f
C502 B.n462 VSUBS 0.007326f
C503 B.n463 VSUBS 0.007326f
C504 B.n464 VSUBS 0.007326f
C505 B.n465 VSUBS 0.007326f
C506 B.n466 VSUBS 0.007326f
C507 B.n467 VSUBS 0.007326f
C508 B.n468 VSUBS 0.007326f
C509 B.n469 VSUBS 0.007326f
C510 B.n470 VSUBS 0.007326f
C511 B.n471 VSUBS 0.007326f
C512 B.n472 VSUBS 0.007326f
C513 B.n473 VSUBS 0.007326f
C514 B.n474 VSUBS 0.007326f
C515 B.n475 VSUBS 0.007326f
C516 B.n476 VSUBS 0.007326f
C517 B.n477 VSUBS 0.007326f
C518 B.n478 VSUBS 0.007326f
C519 B.n479 VSUBS 0.007326f
C520 B.n480 VSUBS 0.007326f
C521 B.n481 VSUBS 0.007326f
C522 B.n482 VSUBS 0.007326f
C523 B.n483 VSUBS 0.007326f
C524 B.n484 VSUBS 0.007326f
C525 B.n485 VSUBS 0.007326f
C526 B.n486 VSUBS 0.007326f
C527 B.n487 VSUBS 0.00956f
C528 B.n488 VSUBS 0.010184f
C529 B.n489 VSUBS 0.020251f
C530 VDD1.n0 VSUBS 0.016008f
C531 VDD1.n1 VSUBS 0.014027f
C532 VDD1.n2 VSUBS 0.007538f
C533 VDD1.n3 VSUBS 0.017816f
C534 VDD1.n4 VSUBS 0.007981f
C535 VDD1.n5 VSUBS 0.014027f
C536 VDD1.n6 VSUBS 0.007538f
C537 VDD1.n7 VSUBS 0.017816f
C538 VDD1.n8 VSUBS 0.007981f
C539 VDD1.n9 VSUBS 0.372291f
C540 VDD1.n10 VSUBS 0.007538f
C541 VDD1.t0 VSUBS 0.038144f
C542 VDD1.n11 VSUBS 0.065192f
C543 VDD1.n12 VSUBS 0.011332f
C544 VDD1.n13 VSUBS 0.013362f
C545 VDD1.n14 VSUBS 0.017816f
C546 VDD1.n15 VSUBS 0.007981f
C547 VDD1.n16 VSUBS 0.007538f
C548 VDD1.n17 VSUBS 0.014027f
C549 VDD1.n18 VSUBS 0.014027f
C550 VDD1.n19 VSUBS 0.007538f
C551 VDD1.n20 VSUBS 0.007981f
C552 VDD1.n21 VSUBS 0.017816f
C553 VDD1.n22 VSUBS 0.017816f
C554 VDD1.n23 VSUBS 0.007981f
C555 VDD1.n24 VSUBS 0.007538f
C556 VDD1.n25 VSUBS 0.014027f
C557 VDD1.n26 VSUBS 0.014027f
C558 VDD1.n27 VSUBS 0.007538f
C559 VDD1.n28 VSUBS 0.007981f
C560 VDD1.n29 VSUBS 0.017816f
C561 VDD1.n30 VSUBS 0.04516f
C562 VDD1.n31 VSUBS 0.007981f
C563 VDD1.n32 VSUBS 0.007538f
C564 VDD1.n33 VSUBS 0.033765f
C565 VDD1.n34 VSUBS 0.033543f
C566 VDD1.n35 VSUBS 0.016008f
C567 VDD1.n36 VSUBS 0.014027f
C568 VDD1.n37 VSUBS 0.007538f
C569 VDD1.n38 VSUBS 0.017816f
C570 VDD1.n39 VSUBS 0.007981f
C571 VDD1.n40 VSUBS 0.014027f
C572 VDD1.n41 VSUBS 0.007538f
C573 VDD1.n42 VSUBS 0.017816f
C574 VDD1.n43 VSUBS 0.007981f
C575 VDD1.n44 VSUBS 0.372291f
C576 VDD1.n45 VSUBS 0.007538f
C577 VDD1.t1 VSUBS 0.038144f
C578 VDD1.n46 VSUBS 0.065192f
C579 VDD1.n47 VSUBS 0.011332f
C580 VDD1.n48 VSUBS 0.013362f
C581 VDD1.n49 VSUBS 0.017816f
C582 VDD1.n50 VSUBS 0.007981f
C583 VDD1.n51 VSUBS 0.007538f
C584 VDD1.n52 VSUBS 0.014027f
C585 VDD1.n53 VSUBS 0.014027f
C586 VDD1.n54 VSUBS 0.007538f
C587 VDD1.n55 VSUBS 0.007981f
C588 VDD1.n56 VSUBS 0.017816f
C589 VDD1.n57 VSUBS 0.017816f
C590 VDD1.n58 VSUBS 0.007981f
C591 VDD1.n59 VSUBS 0.007538f
C592 VDD1.n60 VSUBS 0.014027f
C593 VDD1.n61 VSUBS 0.014027f
C594 VDD1.n62 VSUBS 0.007538f
C595 VDD1.n63 VSUBS 0.007981f
C596 VDD1.n64 VSUBS 0.017816f
C597 VDD1.n65 VSUBS 0.04516f
C598 VDD1.n66 VSUBS 0.007981f
C599 VDD1.n67 VSUBS 0.007538f
C600 VDD1.n68 VSUBS 0.033765f
C601 VDD1.n69 VSUBS 0.357289f
C602 VP.t1 VSUBS 2.77459f
C603 VP.t0 VSUBS 2.13838f
C604 VP.n0 VSUBS 3.28411f
C605 VDD2.n0 VSUBS 0.016657f
C606 VDD2.n1 VSUBS 0.014595f
C607 VDD2.n2 VSUBS 0.007843f
C608 VDD2.n3 VSUBS 0.018538f
C609 VDD2.n4 VSUBS 0.008304f
C610 VDD2.n5 VSUBS 0.014595f
C611 VDD2.n6 VSUBS 0.007843f
C612 VDD2.n7 VSUBS 0.018538f
C613 VDD2.n8 VSUBS 0.008304f
C614 VDD2.n9 VSUBS 0.387369f
C615 VDD2.n10 VSUBS 0.007843f
C616 VDD2.t1 VSUBS 0.039689f
C617 VDD2.n11 VSUBS 0.067832f
C618 VDD2.n12 VSUBS 0.011791f
C619 VDD2.n13 VSUBS 0.013903f
C620 VDD2.n14 VSUBS 0.018538f
C621 VDD2.n15 VSUBS 0.008304f
C622 VDD2.n16 VSUBS 0.007843f
C623 VDD2.n17 VSUBS 0.014595f
C624 VDD2.n18 VSUBS 0.014595f
C625 VDD2.n19 VSUBS 0.007843f
C626 VDD2.n20 VSUBS 0.008304f
C627 VDD2.n21 VSUBS 0.018538f
C628 VDD2.n22 VSUBS 0.018538f
C629 VDD2.n23 VSUBS 0.008304f
C630 VDD2.n24 VSUBS 0.007843f
C631 VDD2.n25 VSUBS 0.014595f
C632 VDD2.n26 VSUBS 0.014595f
C633 VDD2.n27 VSUBS 0.007843f
C634 VDD2.n28 VSUBS 0.008304f
C635 VDD2.n29 VSUBS 0.018538f
C636 VDD2.n30 VSUBS 0.046988f
C637 VDD2.n31 VSUBS 0.008304f
C638 VDD2.n32 VSUBS 0.007843f
C639 VDD2.n33 VSUBS 0.035132f
C640 VDD2.n34 VSUBS 0.343544f
C641 VDD2.n35 VSUBS 0.016657f
C642 VDD2.n36 VSUBS 0.014595f
C643 VDD2.n37 VSUBS 0.007843f
C644 VDD2.n38 VSUBS 0.018538f
C645 VDD2.n39 VSUBS 0.008304f
C646 VDD2.n40 VSUBS 0.014595f
C647 VDD2.n41 VSUBS 0.007843f
C648 VDD2.n42 VSUBS 0.018538f
C649 VDD2.n43 VSUBS 0.008304f
C650 VDD2.n44 VSUBS 0.387369f
C651 VDD2.n45 VSUBS 0.007843f
C652 VDD2.t0 VSUBS 0.039689f
C653 VDD2.n46 VSUBS 0.067832f
C654 VDD2.n47 VSUBS 0.011791f
C655 VDD2.n48 VSUBS 0.013903f
C656 VDD2.n49 VSUBS 0.018538f
C657 VDD2.n50 VSUBS 0.008304f
C658 VDD2.n51 VSUBS 0.007843f
C659 VDD2.n52 VSUBS 0.014595f
C660 VDD2.n53 VSUBS 0.014595f
C661 VDD2.n54 VSUBS 0.007843f
C662 VDD2.n55 VSUBS 0.008304f
C663 VDD2.n56 VSUBS 0.018538f
C664 VDD2.n57 VSUBS 0.018538f
C665 VDD2.n58 VSUBS 0.008304f
C666 VDD2.n59 VSUBS 0.007843f
C667 VDD2.n60 VSUBS 0.014595f
C668 VDD2.n61 VSUBS 0.014595f
C669 VDD2.n62 VSUBS 0.007843f
C670 VDD2.n63 VSUBS 0.008304f
C671 VDD2.n64 VSUBS 0.018538f
C672 VDD2.n65 VSUBS 0.046988f
C673 VDD2.n66 VSUBS 0.008304f
C674 VDD2.n67 VSUBS 0.007843f
C675 VDD2.n68 VSUBS 0.035132f
C676 VDD2.n69 VSUBS 0.033833f
C677 VDD2.n70 VSUBS 1.53498f
C678 VTAIL.n0 VSUBS 0.029414f
C679 VTAIL.n1 VSUBS 0.025774f
C680 VTAIL.n2 VSUBS 0.01385f
C681 VTAIL.n3 VSUBS 0.032736f
C682 VTAIL.n4 VSUBS 0.014664f
C683 VTAIL.n5 VSUBS 0.025774f
C684 VTAIL.n6 VSUBS 0.01385f
C685 VTAIL.n7 VSUBS 0.032736f
C686 VTAIL.n8 VSUBS 0.014664f
C687 VTAIL.n9 VSUBS 0.684048f
C688 VTAIL.n10 VSUBS 0.01385f
C689 VTAIL.t1 VSUBS 0.070085f
C690 VTAIL.n11 VSUBS 0.119784f
C691 VTAIL.n12 VSUBS 0.020821f
C692 VTAIL.n13 VSUBS 0.024552f
C693 VTAIL.n14 VSUBS 0.032736f
C694 VTAIL.n15 VSUBS 0.014664f
C695 VTAIL.n16 VSUBS 0.01385f
C696 VTAIL.n17 VSUBS 0.025774f
C697 VTAIL.n18 VSUBS 0.025774f
C698 VTAIL.n19 VSUBS 0.01385f
C699 VTAIL.n20 VSUBS 0.014664f
C700 VTAIL.n21 VSUBS 0.032736f
C701 VTAIL.n22 VSUBS 0.032736f
C702 VTAIL.n23 VSUBS 0.014664f
C703 VTAIL.n24 VSUBS 0.01385f
C704 VTAIL.n25 VSUBS 0.025774f
C705 VTAIL.n26 VSUBS 0.025774f
C706 VTAIL.n27 VSUBS 0.01385f
C707 VTAIL.n28 VSUBS 0.014664f
C708 VTAIL.n29 VSUBS 0.032736f
C709 VTAIL.n30 VSUBS 0.082976f
C710 VTAIL.n31 VSUBS 0.014664f
C711 VTAIL.n32 VSUBS 0.01385f
C712 VTAIL.n33 VSUBS 0.062039f
C713 VTAIL.n34 VSUBS 0.041968f
C714 VTAIL.n35 VSUBS 1.46729f
C715 VTAIL.n36 VSUBS 0.029414f
C716 VTAIL.n37 VSUBS 0.025774f
C717 VTAIL.n38 VSUBS 0.01385f
C718 VTAIL.n39 VSUBS 0.032736f
C719 VTAIL.n40 VSUBS 0.014664f
C720 VTAIL.n41 VSUBS 0.025774f
C721 VTAIL.n42 VSUBS 0.01385f
C722 VTAIL.n43 VSUBS 0.032736f
C723 VTAIL.n44 VSUBS 0.014664f
C724 VTAIL.n45 VSUBS 0.684047f
C725 VTAIL.n46 VSUBS 0.01385f
C726 VTAIL.t2 VSUBS 0.070085f
C727 VTAIL.n47 VSUBS 0.119784f
C728 VTAIL.n48 VSUBS 0.020821f
C729 VTAIL.n49 VSUBS 0.024552f
C730 VTAIL.n50 VSUBS 0.032736f
C731 VTAIL.n51 VSUBS 0.014664f
C732 VTAIL.n52 VSUBS 0.01385f
C733 VTAIL.n53 VSUBS 0.025774f
C734 VTAIL.n54 VSUBS 0.025774f
C735 VTAIL.n55 VSUBS 0.01385f
C736 VTAIL.n56 VSUBS 0.014664f
C737 VTAIL.n57 VSUBS 0.032736f
C738 VTAIL.n58 VSUBS 0.032736f
C739 VTAIL.n59 VSUBS 0.014664f
C740 VTAIL.n60 VSUBS 0.01385f
C741 VTAIL.n61 VSUBS 0.025774f
C742 VTAIL.n62 VSUBS 0.025774f
C743 VTAIL.n63 VSUBS 0.01385f
C744 VTAIL.n64 VSUBS 0.014664f
C745 VTAIL.n65 VSUBS 0.032736f
C746 VTAIL.n66 VSUBS 0.082976f
C747 VTAIL.n67 VSUBS 0.014664f
C748 VTAIL.n68 VSUBS 0.01385f
C749 VTAIL.n69 VSUBS 0.062039f
C750 VTAIL.n70 VSUBS 0.041968f
C751 VTAIL.n71 VSUBS 1.5251f
C752 VTAIL.n72 VSUBS 0.029414f
C753 VTAIL.n73 VSUBS 0.025774f
C754 VTAIL.n74 VSUBS 0.01385f
C755 VTAIL.n75 VSUBS 0.032736f
C756 VTAIL.n76 VSUBS 0.014664f
C757 VTAIL.n77 VSUBS 0.025774f
C758 VTAIL.n78 VSUBS 0.01385f
C759 VTAIL.n79 VSUBS 0.032736f
C760 VTAIL.n80 VSUBS 0.014664f
C761 VTAIL.n81 VSUBS 0.684047f
C762 VTAIL.n82 VSUBS 0.01385f
C763 VTAIL.t0 VSUBS 0.070085f
C764 VTAIL.n83 VSUBS 0.119784f
C765 VTAIL.n84 VSUBS 0.020821f
C766 VTAIL.n85 VSUBS 0.024552f
C767 VTAIL.n86 VSUBS 0.032736f
C768 VTAIL.n87 VSUBS 0.014664f
C769 VTAIL.n88 VSUBS 0.01385f
C770 VTAIL.n89 VSUBS 0.025774f
C771 VTAIL.n90 VSUBS 0.025774f
C772 VTAIL.n91 VSUBS 0.01385f
C773 VTAIL.n92 VSUBS 0.014664f
C774 VTAIL.n93 VSUBS 0.032736f
C775 VTAIL.n94 VSUBS 0.032736f
C776 VTAIL.n95 VSUBS 0.014664f
C777 VTAIL.n96 VSUBS 0.01385f
C778 VTAIL.n97 VSUBS 0.025774f
C779 VTAIL.n98 VSUBS 0.025774f
C780 VTAIL.n99 VSUBS 0.01385f
C781 VTAIL.n100 VSUBS 0.014664f
C782 VTAIL.n101 VSUBS 0.032736f
C783 VTAIL.n102 VSUBS 0.082976f
C784 VTAIL.n103 VSUBS 0.014664f
C785 VTAIL.n104 VSUBS 0.01385f
C786 VTAIL.n105 VSUBS 0.062039f
C787 VTAIL.n106 VSUBS 0.041968f
C788 VTAIL.n107 VSUBS 1.27452f
C789 VTAIL.n108 VSUBS 0.029414f
C790 VTAIL.n109 VSUBS 0.025774f
C791 VTAIL.n110 VSUBS 0.01385f
C792 VTAIL.n111 VSUBS 0.032736f
C793 VTAIL.n112 VSUBS 0.014664f
C794 VTAIL.n113 VSUBS 0.025774f
C795 VTAIL.n114 VSUBS 0.01385f
C796 VTAIL.n115 VSUBS 0.032736f
C797 VTAIL.n116 VSUBS 0.014664f
C798 VTAIL.n117 VSUBS 0.684048f
C799 VTAIL.n118 VSUBS 0.01385f
C800 VTAIL.t3 VSUBS 0.070085f
C801 VTAIL.n119 VSUBS 0.119784f
C802 VTAIL.n120 VSUBS 0.020821f
C803 VTAIL.n121 VSUBS 0.024552f
C804 VTAIL.n122 VSUBS 0.032736f
C805 VTAIL.n123 VSUBS 0.014664f
C806 VTAIL.n124 VSUBS 0.01385f
C807 VTAIL.n125 VSUBS 0.025774f
C808 VTAIL.n126 VSUBS 0.025774f
C809 VTAIL.n127 VSUBS 0.01385f
C810 VTAIL.n128 VSUBS 0.014664f
C811 VTAIL.n129 VSUBS 0.032736f
C812 VTAIL.n130 VSUBS 0.032736f
C813 VTAIL.n131 VSUBS 0.014664f
C814 VTAIL.n132 VSUBS 0.01385f
C815 VTAIL.n133 VSUBS 0.025774f
C816 VTAIL.n134 VSUBS 0.025774f
C817 VTAIL.n135 VSUBS 0.01385f
C818 VTAIL.n136 VSUBS 0.014664f
C819 VTAIL.n137 VSUBS 0.032736f
C820 VTAIL.n138 VSUBS 0.082976f
C821 VTAIL.n139 VSUBS 0.014664f
C822 VTAIL.n140 VSUBS 0.01385f
C823 VTAIL.n141 VSUBS 0.062039f
C824 VTAIL.n142 VSUBS 0.041968f
C825 VTAIL.n143 VSUBS 1.16802f
C826 VN.t0 VSUBS 2.05427f
C827 VN.t1 VSUBS 2.66102f
.ends

