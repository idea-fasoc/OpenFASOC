* NGSPICE file created from diff_pair_sample_1797.ext - technology: sky130A

.subckt diff_pair_sample_1797 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=1.7394 ps=9.7 w=4.46 l=0.43
X1 B.t11 B.t9 B.t10 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=0 ps=0 w=4.46 l=0.43
X2 B.t8 B.t6 B.t7 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=0 ps=0 w=4.46 l=0.43
X3 B.t5 B.t3 B.t4 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=0 ps=0 w=4.46 l=0.43
X4 B.t2 B.t0 B.t1 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=0 ps=0 w=4.46 l=0.43
X5 VDD2.t1 VN.t0 VTAIL.t1 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=1.7394 ps=9.7 w=4.46 l=0.43
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=1.7394 ps=9.7 w=4.46 l=0.43
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n1274_n1864# sky130_fd_pr__pfet_01v8 ad=1.7394 pd=9.7 as=1.7394 ps=9.7 w=4.46 l=0.43
R0 VP.n0 VP.t0 535.828
R1 VP.n0 VP.t1 502.623
R2 VP VP.n0 0.0516364
R3 VTAIL.n90 VTAIL.n72 756.745
R4 VTAIL.n18 VTAIL.n0 756.745
R5 VTAIL.n66 VTAIL.n48 756.745
R6 VTAIL.n42 VTAIL.n24 756.745
R7 VTAIL.n81 VTAIL.n80 585
R8 VTAIL.n83 VTAIL.n82 585
R9 VTAIL.n76 VTAIL.n75 585
R10 VTAIL.n89 VTAIL.n88 585
R11 VTAIL.n91 VTAIL.n90 585
R12 VTAIL.n9 VTAIL.n8 585
R13 VTAIL.n11 VTAIL.n10 585
R14 VTAIL.n4 VTAIL.n3 585
R15 VTAIL.n17 VTAIL.n16 585
R16 VTAIL.n19 VTAIL.n18 585
R17 VTAIL.n67 VTAIL.n66 585
R18 VTAIL.n65 VTAIL.n64 585
R19 VTAIL.n52 VTAIL.n51 585
R20 VTAIL.n59 VTAIL.n58 585
R21 VTAIL.n57 VTAIL.n56 585
R22 VTAIL.n43 VTAIL.n42 585
R23 VTAIL.n41 VTAIL.n40 585
R24 VTAIL.n28 VTAIL.n27 585
R25 VTAIL.n35 VTAIL.n34 585
R26 VTAIL.n33 VTAIL.n32 585
R27 VTAIL.n79 VTAIL.t1 328.587
R28 VTAIL.n7 VTAIL.t3 328.587
R29 VTAIL.n55 VTAIL.t2 328.587
R30 VTAIL.n31 VTAIL.t0 328.587
R31 VTAIL.n82 VTAIL.n81 171.744
R32 VTAIL.n82 VTAIL.n75 171.744
R33 VTAIL.n89 VTAIL.n75 171.744
R34 VTAIL.n90 VTAIL.n89 171.744
R35 VTAIL.n10 VTAIL.n9 171.744
R36 VTAIL.n10 VTAIL.n3 171.744
R37 VTAIL.n17 VTAIL.n3 171.744
R38 VTAIL.n18 VTAIL.n17 171.744
R39 VTAIL.n66 VTAIL.n65 171.744
R40 VTAIL.n65 VTAIL.n51 171.744
R41 VTAIL.n58 VTAIL.n51 171.744
R42 VTAIL.n58 VTAIL.n57 171.744
R43 VTAIL.n42 VTAIL.n41 171.744
R44 VTAIL.n41 VTAIL.n27 171.744
R45 VTAIL.n34 VTAIL.n27 171.744
R46 VTAIL.n34 VTAIL.n33 171.744
R47 VTAIL.n81 VTAIL.t1 85.8723
R48 VTAIL.n9 VTAIL.t3 85.8723
R49 VTAIL.n57 VTAIL.t2 85.8723
R50 VTAIL.n33 VTAIL.t0 85.8723
R51 VTAIL.n95 VTAIL.n94 30.246
R52 VTAIL.n23 VTAIL.n22 30.246
R53 VTAIL.n71 VTAIL.n70 30.246
R54 VTAIL.n47 VTAIL.n46 30.246
R55 VTAIL.n47 VTAIL.n23 17.5393
R56 VTAIL.n95 VTAIL.n71 16.8841
R57 VTAIL.n80 VTAIL.n79 16.3651
R58 VTAIL.n8 VTAIL.n7 16.3651
R59 VTAIL.n56 VTAIL.n55 16.3651
R60 VTAIL.n32 VTAIL.n31 16.3651
R61 VTAIL.n83 VTAIL.n78 12.8005
R62 VTAIL.n11 VTAIL.n6 12.8005
R63 VTAIL.n59 VTAIL.n54 12.8005
R64 VTAIL.n35 VTAIL.n30 12.8005
R65 VTAIL.n84 VTAIL.n76 12.0247
R66 VTAIL.n12 VTAIL.n4 12.0247
R67 VTAIL.n60 VTAIL.n52 12.0247
R68 VTAIL.n36 VTAIL.n28 12.0247
R69 VTAIL.n88 VTAIL.n87 11.249
R70 VTAIL.n16 VTAIL.n15 11.249
R71 VTAIL.n64 VTAIL.n63 11.249
R72 VTAIL.n40 VTAIL.n39 11.249
R73 VTAIL.n91 VTAIL.n74 10.4732
R74 VTAIL.n19 VTAIL.n2 10.4732
R75 VTAIL.n67 VTAIL.n50 10.4732
R76 VTAIL.n43 VTAIL.n26 10.4732
R77 VTAIL.n92 VTAIL.n72 9.69747
R78 VTAIL.n20 VTAIL.n0 9.69747
R79 VTAIL.n68 VTAIL.n48 9.69747
R80 VTAIL.n44 VTAIL.n24 9.69747
R81 VTAIL.n94 VTAIL.n93 9.45567
R82 VTAIL.n22 VTAIL.n21 9.45567
R83 VTAIL.n70 VTAIL.n69 9.45567
R84 VTAIL.n46 VTAIL.n45 9.45567
R85 VTAIL.n93 VTAIL.n92 9.3005
R86 VTAIL.n74 VTAIL.n73 9.3005
R87 VTAIL.n87 VTAIL.n86 9.3005
R88 VTAIL.n85 VTAIL.n84 9.3005
R89 VTAIL.n78 VTAIL.n77 9.3005
R90 VTAIL.n21 VTAIL.n20 9.3005
R91 VTAIL.n2 VTAIL.n1 9.3005
R92 VTAIL.n15 VTAIL.n14 9.3005
R93 VTAIL.n13 VTAIL.n12 9.3005
R94 VTAIL.n6 VTAIL.n5 9.3005
R95 VTAIL.n69 VTAIL.n68 9.3005
R96 VTAIL.n50 VTAIL.n49 9.3005
R97 VTAIL.n63 VTAIL.n62 9.3005
R98 VTAIL.n61 VTAIL.n60 9.3005
R99 VTAIL.n54 VTAIL.n53 9.3005
R100 VTAIL.n45 VTAIL.n44 9.3005
R101 VTAIL.n26 VTAIL.n25 9.3005
R102 VTAIL.n39 VTAIL.n38 9.3005
R103 VTAIL.n37 VTAIL.n36 9.3005
R104 VTAIL.n30 VTAIL.n29 9.3005
R105 VTAIL.n94 VTAIL.n72 4.26717
R106 VTAIL.n22 VTAIL.n0 4.26717
R107 VTAIL.n70 VTAIL.n48 4.26717
R108 VTAIL.n46 VTAIL.n24 4.26717
R109 VTAIL.n79 VTAIL.n77 3.73474
R110 VTAIL.n7 VTAIL.n5 3.73474
R111 VTAIL.n55 VTAIL.n53 3.73474
R112 VTAIL.n31 VTAIL.n29 3.73474
R113 VTAIL.n92 VTAIL.n91 3.49141
R114 VTAIL.n20 VTAIL.n19 3.49141
R115 VTAIL.n68 VTAIL.n67 3.49141
R116 VTAIL.n44 VTAIL.n43 3.49141
R117 VTAIL.n88 VTAIL.n74 2.71565
R118 VTAIL.n16 VTAIL.n2 2.71565
R119 VTAIL.n64 VTAIL.n50 2.71565
R120 VTAIL.n40 VTAIL.n26 2.71565
R121 VTAIL.n87 VTAIL.n76 1.93989
R122 VTAIL.n15 VTAIL.n4 1.93989
R123 VTAIL.n63 VTAIL.n52 1.93989
R124 VTAIL.n39 VTAIL.n28 1.93989
R125 VTAIL.n84 VTAIL.n83 1.16414
R126 VTAIL.n12 VTAIL.n11 1.16414
R127 VTAIL.n60 VTAIL.n59 1.16414
R128 VTAIL.n36 VTAIL.n35 1.16414
R129 VTAIL.n71 VTAIL.n47 0.797914
R130 VTAIL VTAIL.n23 0.69231
R131 VTAIL.n80 VTAIL.n78 0.388379
R132 VTAIL.n8 VTAIL.n6 0.388379
R133 VTAIL.n56 VTAIL.n54 0.388379
R134 VTAIL.n32 VTAIL.n30 0.388379
R135 VTAIL.n85 VTAIL.n77 0.155672
R136 VTAIL.n86 VTAIL.n85 0.155672
R137 VTAIL.n86 VTAIL.n73 0.155672
R138 VTAIL.n93 VTAIL.n73 0.155672
R139 VTAIL.n13 VTAIL.n5 0.155672
R140 VTAIL.n14 VTAIL.n13 0.155672
R141 VTAIL.n14 VTAIL.n1 0.155672
R142 VTAIL.n21 VTAIL.n1 0.155672
R143 VTAIL.n69 VTAIL.n49 0.155672
R144 VTAIL.n62 VTAIL.n49 0.155672
R145 VTAIL.n62 VTAIL.n61 0.155672
R146 VTAIL.n61 VTAIL.n53 0.155672
R147 VTAIL.n45 VTAIL.n25 0.155672
R148 VTAIL.n38 VTAIL.n25 0.155672
R149 VTAIL.n38 VTAIL.n37 0.155672
R150 VTAIL.n37 VTAIL.n29 0.155672
R151 VTAIL VTAIL.n95 0.106103
R152 VDD1.n18 VDD1.n0 756.745
R153 VDD1.n41 VDD1.n23 756.745
R154 VDD1.n19 VDD1.n18 585
R155 VDD1.n17 VDD1.n16 585
R156 VDD1.n4 VDD1.n3 585
R157 VDD1.n11 VDD1.n10 585
R158 VDD1.n9 VDD1.n8 585
R159 VDD1.n32 VDD1.n31 585
R160 VDD1.n34 VDD1.n33 585
R161 VDD1.n27 VDD1.n26 585
R162 VDD1.n40 VDD1.n39 585
R163 VDD1.n42 VDD1.n41 585
R164 VDD1.n7 VDD1.t1 328.587
R165 VDD1.n30 VDD1.t0 328.587
R166 VDD1.n18 VDD1.n17 171.744
R167 VDD1.n17 VDD1.n3 171.744
R168 VDD1.n10 VDD1.n3 171.744
R169 VDD1.n10 VDD1.n9 171.744
R170 VDD1.n33 VDD1.n32 171.744
R171 VDD1.n33 VDD1.n26 171.744
R172 VDD1.n40 VDD1.n26 171.744
R173 VDD1.n41 VDD1.n40 171.744
R174 VDD1.n9 VDD1.t1 85.8723
R175 VDD1.n32 VDD1.t0 85.8723
R176 VDD1 VDD1.n45 76.4452
R177 VDD1 VDD1.n22 47.1467
R178 VDD1.n8 VDD1.n7 16.3651
R179 VDD1.n31 VDD1.n30 16.3651
R180 VDD1.n11 VDD1.n6 12.8005
R181 VDD1.n34 VDD1.n29 12.8005
R182 VDD1.n12 VDD1.n4 12.0247
R183 VDD1.n35 VDD1.n27 12.0247
R184 VDD1.n16 VDD1.n15 11.249
R185 VDD1.n39 VDD1.n38 11.249
R186 VDD1.n19 VDD1.n2 10.4732
R187 VDD1.n42 VDD1.n25 10.4732
R188 VDD1.n20 VDD1.n0 9.69747
R189 VDD1.n43 VDD1.n23 9.69747
R190 VDD1.n22 VDD1.n21 9.45567
R191 VDD1.n45 VDD1.n44 9.45567
R192 VDD1.n21 VDD1.n20 9.3005
R193 VDD1.n2 VDD1.n1 9.3005
R194 VDD1.n15 VDD1.n14 9.3005
R195 VDD1.n13 VDD1.n12 9.3005
R196 VDD1.n6 VDD1.n5 9.3005
R197 VDD1.n44 VDD1.n43 9.3005
R198 VDD1.n25 VDD1.n24 9.3005
R199 VDD1.n38 VDD1.n37 9.3005
R200 VDD1.n36 VDD1.n35 9.3005
R201 VDD1.n29 VDD1.n28 9.3005
R202 VDD1.n22 VDD1.n0 4.26717
R203 VDD1.n45 VDD1.n23 4.26717
R204 VDD1.n7 VDD1.n5 3.73474
R205 VDD1.n30 VDD1.n28 3.73474
R206 VDD1.n20 VDD1.n19 3.49141
R207 VDD1.n43 VDD1.n42 3.49141
R208 VDD1.n16 VDD1.n2 2.71565
R209 VDD1.n39 VDD1.n25 2.71565
R210 VDD1.n15 VDD1.n4 1.93989
R211 VDD1.n38 VDD1.n27 1.93989
R212 VDD1.n12 VDD1.n11 1.16414
R213 VDD1.n35 VDD1.n34 1.16414
R214 VDD1.n8 VDD1.n6 0.388379
R215 VDD1.n31 VDD1.n29 0.388379
R216 VDD1.n21 VDD1.n1 0.155672
R217 VDD1.n14 VDD1.n1 0.155672
R218 VDD1.n14 VDD1.n13 0.155672
R219 VDD1.n13 VDD1.n5 0.155672
R220 VDD1.n36 VDD1.n28 0.155672
R221 VDD1.n37 VDD1.n36 0.155672
R222 VDD1.n37 VDD1.n24 0.155672
R223 VDD1.n44 VDD1.n24 0.155672
R224 B.n175 B.n50 585
R225 B.n174 B.n173 585
R226 B.n172 B.n51 585
R227 B.n171 B.n170 585
R228 B.n169 B.n52 585
R229 B.n168 B.n167 585
R230 B.n166 B.n53 585
R231 B.n165 B.n164 585
R232 B.n163 B.n54 585
R233 B.n162 B.n161 585
R234 B.n160 B.n55 585
R235 B.n159 B.n158 585
R236 B.n157 B.n56 585
R237 B.n156 B.n155 585
R238 B.n154 B.n57 585
R239 B.n153 B.n152 585
R240 B.n151 B.n58 585
R241 B.n150 B.n149 585
R242 B.n148 B.n59 585
R243 B.n147 B.n146 585
R244 B.n145 B.n144 585
R245 B.n143 B.n63 585
R246 B.n142 B.n141 585
R247 B.n140 B.n64 585
R248 B.n139 B.n138 585
R249 B.n137 B.n65 585
R250 B.n136 B.n135 585
R251 B.n134 B.n66 585
R252 B.n133 B.n132 585
R253 B.n130 B.n67 585
R254 B.n129 B.n128 585
R255 B.n127 B.n70 585
R256 B.n126 B.n125 585
R257 B.n124 B.n71 585
R258 B.n123 B.n122 585
R259 B.n121 B.n72 585
R260 B.n120 B.n119 585
R261 B.n118 B.n73 585
R262 B.n117 B.n116 585
R263 B.n115 B.n74 585
R264 B.n114 B.n113 585
R265 B.n112 B.n75 585
R266 B.n111 B.n110 585
R267 B.n109 B.n76 585
R268 B.n108 B.n107 585
R269 B.n106 B.n77 585
R270 B.n105 B.n104 585
R271 B.n103 B.n78 585
R272 B.n102 B.n101 585
R273 B.n177 B.n176 585
R274 B.n178 B.n49 585
R275 B.n180 B.n179 585
R276 B.n181 B.n48 585
R277 B.n183 B.n182 585
R278 B.n184 B.n47 585
R279 B.n186 B.n185 585
R280 B.n187 B.n46 585
R281 B.n189 B.n188 585
R282 B.n190 B.n45 585
R283 B.n192 B.n191 585
R284 B.n193 B.n44 585
R285 B.n195 B.n194 585
R286 B.n196 B.n43 585
R287 B.n198 B.n197 585
R288 B.n199 B.n42 585
R289 B.n201 B.n200 585
R290 B.n202 B.n41 585
R291 B.n204 B.n203 585
R292 B.n205 B.n40 585
R293 B.n207 B.n206 585
R294 B.n208 B.n39 585
R295 B.n210 B.n209 585
R296 B.n211 B.n38 585
R297 B.n213 B.n212 585
R298 B.n214 B.n37 585
R299 B.n289 B.n8 585
R300 B.n288 B.n287 585
R301 B.n286 B.n9 585
R302 B.n285 B.n284 585
R303 B.n283 B.n10 585
R304 B.n282 B.n281 585
R305 B.n280 B.n11 585
R306 B.n279 B.n278 585
R307 B.n277 B.n12 585
R308 B.n276 B.n275 585
R309 B.n274 B.n13 585
R310 B.n273 B.n272 585
R311 B.n271 B.n14 585
R312 B.n270 B.n269 585
R313 B.n268 B.n15 585
R314 B.n267 B.n266 585
R315 B.n265 B.n16 585
R316 B.n264 B.n263 585
R317 B.n262 B.n17 585
R318 B.n261 B.n260 585
R319 B.n259 B.n258 585
R320 B.n257 B.n21 585
R321 B.n256 B.n255 585
R322 B.n254 B.n22 585
R323 B.n253 B.n252 585
R324 B.n251 B.n23 585
R325 B.n250 B.n249 585
R326 B.n248 B.n24 585
R327 B.n247 B.n246 585
R328 B.n244 B.n25 585
R329 B.n243 B.n242 585
R330 B.n241 B.n28 585
R331 B.n240 B.n239 585
R332 B.n238 B.n29 585
R333 B.n237 B.n236 585
R334 B.n235 B.n30 585
R335 B.n234 B.n233 585
R336 B.n232 B.n31 585
R337 B.n231 B.n230 585
R338 B.n229 B.n32 585
R339 B.n228 B.n227 585
R340 B.n226 B.n33 585
R341 B.n225 B.n224 585
R342 B.n223 B.n34 585
R343 B.n222 B.n221 585
R344 B.n220 B.n35 585
R345 B.n219 B.n218 585
R346 B.n217 B.n36 585
R347 B.n216 B.n215 585
R348 B.n291 B.n290 585
R349 B.n292 B.n7 585
R350 B.n294 B.n293 585
R351 B.n295 B.n6 585
R352 B.n297 B.n296 585
R353 B.n298 B.n5 585
R354 B.n300 B.n299 585
R355 B.n301 B.n4 585
R356 B.n303 B.n302 585
R357 B.n304 B.n3 585
R358 B.n306 B.n305 585
R359 B.n307 B.n0 585
R360 B.n2 B.n1 585
R361 B.n85 B.n84 585
R362 B.n87 B.n86 585
R363 B.n88 B.n83 585
R364 B.n90 B.n89 585
R365 B.n91 B.n82 585
R366 B.n93 B.n92 585
R367 B.n94 B.n81 585
R368 B.n96 B.n95 585
R369 B.n97 B.n80 585
R370 B.n99 B.n98 585
R371 B.n100 B.n79 585
R372 B.n102 B.n79 478.086
R373 B.n176 B.n175 478.086
R374 B.n216 B.n37 478.086
R375 B.n290 B.n289 478.086
R376 B.n68 B.t6 458.337
R377 B.n60 B.t0 458.337
R378 B.n26 B.t9 458.337
R379 B.n18 B.t3 458.337
R380 B.n309 B.n308 256.663
R381 B.n60 B.t1 256.368
R382 B.n26 B.t11 256.368
R383 B.n68 B.t7 256.368
R384 B.n18 B.t5 256.368
R385 B.n61 B.t2 241.63
R386 B.n27 B.t10 241.63
R387 B.n69 B.t8 241.63
R388 B.n19 B.t4 241.63
R389 B.n308 B.n307 235.042
R390 B.n308 B.n2 235.042
R391 B.n103 B.n102 163.367
R392 B.n104 B.n103 163.367
R393 B.n104 B.n77 163.367
R394 B.n108 B.n77 163.367
R395 B.n109 B.n108 163.367
R396 B.n110 B.n109 163.367
R397 B.n110 B.n75 163.367
R398 B.n114 B.n75 163.367
R399 B.n115 B.n114 163.367
R400 B.n116 B.n115 163.367
R401 B.n116 B.n73 163.367
R402 B.n120 B.n73 163.367
R403 B.n121 B.n120 163.367
R404 B.n122 B.n121 163.367
R405 B.n122 B.n71 163.367
R406 B.n126 B.n71 163.367
R407 B.n127 B.n126 163.367
R408 B.n128 B.n127 163.367
R409 B.n128 B.n67 163.367
R410 B.n133 B.n67 163.367
R411 B.n134 B.n133 163.367
R412 B.n135 B.n134 163.367
R413 B.n135 B.n65 163.367
R414 B.n139 B.n65 163.367
R415 B.n140 B.n139 163.367
R416 B.n141 B.n140 163.367
R417 B.n141 B.n63 163.367
R418 B.n145 B.n63 163.367
R419 B.n146 B.n145 163.367
R420 B.n146 B.n59 163.367
R421 B.n150 B.n59 163.367
R422 B.n151 B.n150 163.367
R423 B.n152 B.n151 163.367
R424 B.n152 B.n57 163.367
R425 B.n156 B.n57 163.367
R426 B.n157 B.n156 163.367
R427 B.n158 B.n157 163.367
R428 B.n158 B.n55 163.367
R429 B.n162 B.n55 163.367
R430 B.n163 B.n162 163.367
R431 B.n164 B.n163 163.367
R432 B.n164 B.n53 163.367
R433 B.n168 B.n53 163.367
R434 B.n169 B.n168 163.367
R435 B.n170 B.n169 163.367
R436 B.n170 B.n51 163.367
R437 B.n174 B.n51 163.367
R438 B.n175 B.n174 163.367
R439 B.n212 B.n37 163.367
R440 B.n212 B.n211 163.367
R441 B.n211 B.n210 163.367
R442 B.n210 B.n39 163.367
R443 B.n206 B.n39 163.367
R444 B.n206 B.n205 163.367
R445 B.n205 B.n204 163.367
R446 B.n204 B.n41 163.367
R447 B.n200 B.n41 163.367
R448 B.n200 B.n199 163.367
R449 B.n199 B.n198 163.367
R450 B.n198 B.n43 163.367
R451 B.n194 B.n43 163.367
R452 B.n194 B.n193 163.367
R453 B.n193 B.n192 163.367
R454 B.n192 B.n45 163.367
R455 B.n188 B.n45 163.367
R456 B.n188 B.n187 163.367
R457 B.n187 B.n186 163.367
R458 B.n186 B.n47 163.367
R459 B.n182 B.n47 163.367
R460 B.n182 B.n181 163.367
R461 B.n181 B.n180 163.367
R462 B.n180 B.n49 163.367
R463 B.n176 B.n49 163.367
R464 B.n289 B.n288 163.367
R465 B.n288 B.n9 163.367
R466 B.n284 B.n9 163.367
R467 B.n284 B.n283 163.367
R468 B.n283 B.n282 163.367
R469 B.n282 B.n11 163.367
R470 B.n278 B.n11 163.367
R471 B.n278 B.n277 163.367
R472 B.n277 B.n276 163.367
R473 B.n276 B.n13 163.367
R474 B.n272 B.n13 163.367
R475 B.n272 B.n271 163.367
R476 B.n271 B.n270 163.367
R477 B.n270 B.n15 163.367
R478 B.n266 B.n15 163.367
R479 B.n266 B.n265 163.367
R480 B.n265 B.n264 163.367
R481 B.n264 B.n17 163.367
R482 B.n260 B.n17 163.367
R483 B.n260 B.n259 163.367
R484 B.n259 B.n21 163.367
R485 B.n255 B.n21 163.367
R486 B.n255 B.n254 163.367
R487 B.n254 B.n253 163.367
R488 B.n253 B.n23 163.367
R489 B.n249 B.n23 163.367
R490 B.n249 B.n248 163.367
R491 B.n248 B.n247 163.367
R492 B.n247 B.n25 163.367
R493 B.n242 B.n25 163.367
R494 B.n242 B.n241 163.367
R495 B.n241 B.n240 163.367
R496 B.n240 B.n29 163.367
R497 B.n236 B.n29 163.367
R498 B.n236 B.n235 163.367
R499 B.n235 B.n234 163.367
R500 B.n234 B.n31 163.367
R501 B.n230 B.n31 163.367
R502 B.n230 B.n229 163.367
R503 B.n229 B.n228 163.367
R504 B.n228 B.n33 163.367
R505 B.n224 B.n33 163.367
R506 B.n224 B.n223 163.367
R507 B.n223 B.n222 163.367
R508 B.n222 B.n35 163.367
R509 B.n218 B.n35 163.367
R510 B.n218 B.n217 163.367
R511 B.n217 B.n216 163.367
R512 B.n290 B.n7 163.367
R513 B.n294 B.n7 163.367
R514 B.n295 B.n294 163.367
R515 B.n296 B.n295 163.367
R516 B.n296 B.n5 163.367
R517 B.n300 B.n5 163.367
R518 B.n301 B.n300 163.367
R519 B.n302 B.n301 163.367
R520 B.n302 B.n3 163.367
R521 B.n306 B.n3 163.367
R522 B.n307 B.n306 163.367
R523 B.n85 B.n2 163.367
R524 B.n86 B.n85 163.367
R525 B.n86 B.n83 163.367
R526 B.n90 B.n83 163.367
R527 B.n91 B.n90 163.367
R528 B.n92 B.n91 163.367
R529 B.n92 B.n81 163.367
R530 B.n96 B.n81 163.367
R531 B.n97 B.n96 163.367
R532 B.n98 B.n97 163.367
R533 B.n98 B.n79 163.367
R534 B.n131 B.n69 59.5399
R535 B.n62 B.n61 59.5399
R536 B.n245 B.n27 59.5399
R537 B.n20 B.n19 59.5399
R538 B.n291 B.n8 31.0639
R539 B.n215 B.n214 31.0639
R540 B.n177 B.n50 31.0639
R541 B.n101 B.n100 31.0639
R542 B B.n309 18.0485
R543 B.n69 B.n68 14.7399
R544 B.n61 B.n60 14.7399
R545 B.n27 B.n26 14.7399
R546 B.n19 B.n18 14.7399
R547 B.n292 B.n291 10.6151
R548 B.n293 B.n292 10.6151
R549 B.n293 B.n6 10.6151
R550 B.n297 B.n6 10.6151
R551 B.n298 B.n297 10.6151
R552 B.n299 B.n298 10.6151
R553 B.n299 B.n4 10.6151
R554 B.n303 B.n4 10.6151
R555 B.n304 B.n303 10.6151
R556 B.n305 B.n304 10.6151
R557 B.n305 B.n0 10.6151
R558 B.n287 B.n8 10.6151
R559 B.n287 B.n286 10.6151
R560 B.n286 B.n285 10.6151
R561 B.n285 B.n10 10.6151
R562 B.n281 B.n10 10.6151
R563 B.n281 B.n280 10.6151
R564 B.n280 B.n279 10.6151
R565 B.n279 B.n12 10.6151
R566 B.n275 B.n12 10.6151
R567 B.n275 B.n274 10.6151
R568 B.n274 B.n273 10.6151
R569 B.n273 B.n14 10.6151
R570 B.n269 B.n14 10.6151
R571 B.n269 B.n268 10.6151
R572 B.n268 B.n267 10.6151
R573 B.n267 B.n16 10.6151
R574 B.n263 B.n16 10.6151
R575 B.n263 B.n262 10.6151
R576 B.n262 B.n261 10.6151
R577 B.n258 B.n257 10.6151
R578 B.n257 B.n256 10.6151
R579 B.n256 B.n22 10.6151
R580 B.n252 B.n22 10.6151
R581 B.n252 B.n251 10.6151
R582 B.n251 B.n250 10.6151
R583 B.n250 B.n24 10.6151
R584 B.n246 B.n24 10.6151
R585 B.n244 B.n243 10.6151
R586 B.n243 B.n28 10.6151
R587 B.n239 B.n28 10.6151
R588 B.n239 B.n238 10.6151
R589 B.n238 B.n237 10.6151
R590 B.n237 B.n30 10.6151
R591 B.n233 B.n30 10.6151
R592 B.n233 B.n232 10.6151
R593 B.n232 B.n231 10.6151
R594 B.n231 B.n32 10.6151
R595 B.n227 B.n32 10.6151
R596 B.n227 B.n226 10.6151
R597 B.n226 B.n225 10.6151
R598 B.n225 B.n34 10.6151
R599 B.n221 B.n34 10.6151
R600 B.n221 B.n220 10.6151
R601 B.n220 B.n219 10.6151
R602 B.n219 B.n36 10.6151
R603 B.n215 B.n36 10.6151
R604 B.n214 B.n213 10.6151
R605 B.n213 B.n38 10.6151
R606 B.n209 B.n38 10.6151
R607 B.n209 B.n208 10.6151
R608 B.n208 B.n207 10.6151
R609 B.n207 B.n40 10.6151
R610 B.n203 B.n40 10.6151
R611 B.n203 B.n202 10.6151
R612 B.n202 B.n201 10.6151
R613 B.n201 B.n42 10.6151
R614 B.n197 B.n42 10.6151
R615 B.n197 B.n196 10.6151
R616 B.n196 B.n195 10.6151
R617 B.n195 B.n44 10.6151
R618 B.n191 B.n44 10.6151
R619 B.n191 B.n190 10.6151
R620 B.n190 B.n189 10.6151
R621 B.n189 B.n46 10.6151
R622 B.n185 B.n46 10.6151
R623 B.n185 B.n184 10.6151
R624 B.n184 B.n183 10.6151
R625 B.n183 B.n48 10.6151
R626 B.n179 B.n48 10.6151
R627 B.n179 B.n178 10.6151
R628 B.n178 B.n177 10.6151
R629 B.n84 B.n1 10.6151
R630 B.n87 B.n84 10.6151
R631 B.n88 B.n87 10.6151
R632 B.n89 B.n88 10.6151
R633 B.n89 B.n82 10.6151
R634 B.n93 B.n82 10.6151
R635 B.n94 B.n93 10.6151
R636 B.n95 B.n94 10.6151
R637 B.n95 B.n80 10.6151
R638 B.n99 B.n80 10.6151
R639 B.n100 B.n99 10.6151
R640 B.n101 B.n78 10.6151
R641 B.n105 B.n78 10.6151
R642 B.n106 B.n105 10.6151
R643 B.n107 B.n106 10.6151
R644 B.n107 B.n76 10.6151
R645 B.n111 B.n76 10.6151
R646 B.n112 B.n111 10.6151
R647 B.n113 B.n112 10.6151
R648 B.n113 B.n74 10.6151
R649 B.n117 B.n74 10.6151
R650 B.n118 B.n117 10.6151
R651 B.n119 B.n118 10.6151
R652 B.n119 B.n72 10.6151
R653 B.n123 B.n72 10.6151
R654 B.n124 B.n123 10.6151
R655 B.n125 B.n124 10.6151
R656 B.n125 B.n70 10.6151
R657 B.n129 B.n70 10.6151
R658 B.n130 B.n129 10.6151
R659 B.n132 B.n66 10.6151
R660 B.n136 B.n66 10.6151
R661 B.n137 B.n136 10.6151
R662 B.n138 B.n137 10.6151
R663 B.n138 B.n64 10.6151
R664 B.n142 B.n64 10.6151
R665 B.n143 B.n142 10.6151
R666 B.n144 B.n143 10.6151
R667 B.n148 B.n147 10.6151
R668 B.n149 B.n148 10.6151
R669 B.n149 B.n58 10.6151
R670 B.n153 B.n58 10.6151
R671 B.n154 B.n153 10.6151
R672 B.n155 B.n154 10.6151
R673 B.n155 B.n56 10.6151
R674 B.n159 B.n56 10.6151
R675 B.n160 B.n159 10.6151
R676 B.n161 B.n160 10.6151
R677 B.n161 B.n54 10.6151
R678 B.n165 B.n54 10.6151
R679 B.n166 B.n165 10.6151
R680 B.n167 B.n166 10.6151
R681 B.n167 B.n52 10.6151
R682 B.n171 B.n52 10.6151
R683 B.n172 B.n171 10.6151
R684 B.n173 B.n172 10.6151
R685 B.n173 B.n50 10.6151
R686 B.n309 B.n0 8.11757
R687 B.n309 B.n1 8.11757
R688 B.n258 B.n20 7.18099
R689 B.n246 B.n245 7.18099
R690 B.n132 B.n131 7.18099
R691 B.n144 B.n62 7.18099
R692 B.n261 B.n20 3.43465
R693 B.n245 B.n244 3.43465
R694 B.n131 B.n130 3.43465
R695 B.n147 B.n62 3.43465
R696 VN VN.t1 536.208
R697 VN VN.t0 502.675
R698 VDD2.n41 VDD2.n23 756.745
R699 VDD2.n18 VDD2.n0 756.745
R700 VDD2.n42 VDD2.n41 585
R701 VDD2.n40 VDD2.n39 585
R702 VDD2.n27 VDD2.n26 585
R703 VDD2.n34 VDD2.n33 585
R704 VDD2.n32 VDD2.n31 585
R705 VDD2.n9 VDD2.n8 585
R706 VDD2.n11 VDD2.n10 585
R707 VDD2.n4 VDD2.n3 585
R708 VDD2.n17 VDD2.n16 585
R709 VDD2.n19 VDD2.n18 585
R710 VDD2.n30 VDD2.t0 328.587
R711 VDD2.n7 VDD2.t1 328.587
R712 VDD2.n41 VDD2.n40 171.744
R713 VDD2.n40 VDD2.n26 171.744
R714 VDD2.n33 VDD2.n26 171.744
R715 VDD2.n33 VDD2.n32 171.744
R716 VDD2.n10 VDD2.n9 171.744
R717 VDD2.n10 VDD2.n3 171.744
R718 VDD2.n17 VDD2.n3 171.744
R719 VDD2.n18 VDD2.n17 171.744
R720 VDD2.n32 VDD2.t0 85.8723
R721 VDD2.n9 VDD2.t1 85.8723
R722 VDD2.n46 VDD2.n22 75.7566
R723 VDD2.n46 VDD2.n45 46.9247
R724 VDD2.n31 VDD2.n30 16.3651
R725 VDD2.n8 VDD2.n7 16.3651
R726 VDD2.n34 VDD2.n29 12.8005
R727 VDD2.n11 VDD2.n6 12.8005
R728 VDD2.n35 VDD2.n27 12.0247
R729 VDD2.n12 VDD2.n4 12.0247
R730 VDD2.n39 VDD2.n38 11.249
R731 VDD2.n16 VDD2.n15 11.249
R732 VDD2.n42 VDD2.n25 10.4732
R733 VDD2.n19 VDD2.n2 10.4732
R734 VDD2.n43 VDD2.n23 9.69747
R735 VDD2.n20 VDD2.n0 9.69747
R736 VDD2.n45 VDD2.n44 9.45567
R737 VDD2.n22 VDD2.n21 9.45567
R738 VDD2.n44 VDD2.n43 9.3005
R739 VDD2.n25 VDD2.n24 9.3005
R740 VDD2.n38 VDD2.n37 9.3005
R741 VDD2.n36 VDD2.n35 9.3005
R742 VDD2.n29 VDD2.n28 9.3005
R743 VDD2.n21 VDD2.n20 9.3005
R744 VDD2.n2 VDD2.n1 9.3005
R745 VDD2.n15 VDD2.n14 9.3005
R746 VDD2.n13 VDD2.n12 9.3005
R747 VDD2.n6 VDD2.n5 9.3005
R748 VDD2.n45 VDD2.n23 4.26717
R749 VDD2.n22 VDD2.n0 4.26717
R750 VDD2.n30 VDD2.n28 3.73474
R751 VDD2.n7 VDD2.n5 3.73474
R752 VDD2.n43 VDD2.n42 3.49141
R753 VDD2.n20 VDD2.n19 3.49141
R754 VDD2.n39 VDD2.n25 2.71565
R755 VDD2.n16 VDD2.n2 2.71565
R756 VDD2.n38 VDD2.n27 1.93989
R757 VDD2.n15 VDD2.n4 1.93989
R758 VDD2.n35 VDD2.n34 1.16414
R759 VDD2.n12 VDD2.n11 1.16414
R760 VDD2.n31 VDD2.n29 0.388379
R761 VDD2.n8 VDD2.n6 0.388379
R762 VDD2 VDD2.n46 0.222483
R763 VDD2.n44 VDD2.n24 0.155672
R764 VDD2.n37 VDD2.n24 0.155672
R765 VDD2.n37 VDD2.n36 0.155672
R766 VDD2.n36 VDD2.n28 0.155672
R767 VDD2.n13 VDD2.n5 0.155672
R768 VDD2.n14 VDD2.n13 0.155672
R769 VDD2.n14 VDD2.n1 0.155672
R770 VDD2.n21 VDD2.n1 0.155672
C0 VDD1 B 0.828145f
C1 VN VTAIL 0.599191f
C2 VP VTAIL 0.61352f
C3 VDD1 w_n1274_n1864# 0.977945f
C4 B VTAIL 1.24713f
C5 VN VDD2 0.760797f
C6 VDD2 VP 0.247153f
C7 w_n1274_n1864# VTAIL 1.66686f
C8 B VDD2 0.840902f
C9 VN VP 3.04659f
C10 VN B 0.591996f
C11 VDD2 w_n1274_n1864# 0.979576f
C12 B VP 0.842284f
C13 VN w_n1274_n1864# 1.43312f
C14 w_n1274_n1864# VP 1.59044f
C15 B w_n1274_n1864# 4.34997f
C16 VDD1 VTAIL 3.07329f
C17 VDD1 VDD2 0.43512f
C18 VDD1 VN 0.152799f
C19 VDD2 VTAIL 3.10906f
C20 VDD1 VP 0.85296f
C21 VDD2 VSUBS 0.45954f
C22 VDD1 VSUBS 1.88674f
C23 VTAIL VSUBS 0.141825f
C24 VN VSUBS 3.57581f
C25 VP VSUBS 0.679984f
C26 B VSUBS 1.592416f
C27 w_n1274_n1864# VSUBS 29.8269f
C28 VDD2.n0 VSUBS 0.018034f
C29 VDD2.n1 VSUBS 0.01771f
C30 VDD2.n2 VSUBS 0.009517f
C31 VDD2.n3 VSUBS 0.022494f
C32 VDD2.n4 VSUBS 0.010076f
C33 VDD2.n5 VSUBS 0.281939f
C34 VDD2.n6 VSUBS 0.009517f
C35 VDD2.t1 VSUBS 0.048566f
C36 VDD2.n7 VSUBS 0.070449f
C37 VDD2.n8 VSUBS 0.01425f
C38 VDD2.n9 VSUBS 0.01687f
C39 VDD2.n10 VSUBS 0.022494f
C40 VDD2.n11 VSUBS 0.010076f
C41 VDD2.n12 VSUBS 0.009517f
C42 VDD2.n13 VSUBS 0.01771f
C43 VDD2.n14 VSUBS 0.01771f
C44 VDD2.n15 VSUBS 0.009517f
C45 VDD2.n16 VSUBS 0.010076f
C46 VDD2.n17 VSUBS 0.022494f
C47 VDD2.n18 VSUBS 0.0496f
C48 VDD2.n19 VSUBS 0.010076f
C49 VDD2.n20 VSUBS 0.009517f
C50 VDD2.n21 VSUBS 0.038517f
C51 VDD2.n22 VSUBS 0.265655f
C52 VDD2.n23 VSUBS 0.018034f
C53 VDD2.n24 VSUBS 0.01771f
C54 VDD2.n25 VSUBS 0.009517f
C55 VDD2.n26 VSUBS 0.022494f
C56 VDD2.n27 VSUBS 0.010076f
C57 VDD2.n28 VSUBS 0.281939f
C58 VDD2.n29 VSUBS 0.009517f
C59 VDD2.t0 VSUBS 0.048566f
C60 VDD2.n30 VSUBS 0.070449f
C61 VDD2.n31 VSUBS 0.01425f
C62 VDD2.n32 VSUBS 0.01687f
C63 VDD2.n33 VSUBS 0.022494f
C64 VDD2.n34 VSUBS 0.010076f
C65 VDD2.n35 VSUBS 0.009517f
C66 VDD2.n36 VSUBS 0.01771f
C67 VDD2.n37 VSUBS 0.01771f
C68 VDD2.n38 VSUBS 0.009517f
C69 VDD2.n39 VSUBS 0.010076f
C70 VDD2.n40 VSUBS 0.022494f
C71 VDD2.n41 VSUBS 0.0496f
C72 VDD2.n42 VSUBS 0.010076f
C73 VDD2.n43 VSUBS 0.009517f
C74 VDD2.n44 VSUBS 0.038517f
C75 VDD2.n45 VSUBS 0.036901f
C76 VDD2.n46 VSUBS 1.27214f
C77 VN.t0 VSUBS 0.268f
C78 VN.t1 VSUBS 0.343647f
C79 B.n0 VSUBS 0.006404f
C80 B.n1 VSUBS 0.006404f
C81 B.n2 VSUBS 0.009471f
C82 B.n3 VSUBS 0.007257f
C83 B.n4 VSUBS 0.007257f
C84 B.n5 VSUBS 0.007257f
C85 B.n6 VSUBS 0.007257f
C86 B.n7 VSUBS 0.007257f
C87 B.n8 VSUBS 0.017084f
C88 B.n9 VSUBS 0.007257f
C89 B.n10 VSUBS 0.007257f
C90 B.n11 VSUBS 0.007257f
C91 B.n12 VSUBS 0.007257f
C92 B.n13 VSUBS 0.007257f
C93 B.n14 VSUBS 0.007257f
C94 B.n15 VSUBS 0.007257f
C95 B.n16 VSUBS 0.007257f
C96 B.n17 VSUBS 0.007257f
C97 B.t4 VSUBS 0.066399f
C98 B.t5 VSUBS 0.07279f
C99 B.t3 VSUBS 0.084962f
C100 B.n18 VSUBS 0.131864f
C101 B.n19 VSUBS 0.121527f
C102 B.n20 VSUBS 0.016815f
C103 B.n21 VSUBS 0.007257f
C104 B.n22 VSUBS 0.007257f
C105 B.n23 VSUBS 0.007257f
C106 B.n24 VSUBS 0.007257f
C107 B.n25 VSUBS 0.007257f
C108 B.t10 VSUBS 0.0664f
C109 B.t11 VSUBS 0.072792f
C110 B.t9 VSUBS 0.084962f
C111 B.n26 VSUBS 0.131863f
C112 B.n27 VSUBS 0.121526f
C113 B.n28 VSUBS 0.007257f
C114 B.n29 VSUBS 0.007257f
C115 B.n30 VSUBS 0.007257f
C116 B.n31 VSUBS 0.007257f
C117 B.n32 VSUBS 0.007257f
C118 B.n33 VSUBS 0.007257f
C119 B.n34 VSUBS 0.007257f
C120 B.n35 VSUBS 0.007257f
C121 B.n36 VSUBS 0.007257f
C122 B.n37 VSUBS 0.015787f
C123 B.n38 VSUBS 0.007257f
C124 B.n39 VSUBS 0.007257f
C125 B.n40 VSUBS 0.007257f
C126 B.n41 VSUBS 0.007257f
C127 B.n42 VSUBS 0.007257f
C128 B.n43 VSUBS 0.007257f
C129 B.n44 VSUBS 0.007257f
C130 B.n45 VSUBS 0.007257f
C131 B.n46 VSUBS 0.007257f
C132 B.n47 VSUBS 0.007257f
C133 B.n48 VSUBS 0.007257f
C134 B.n49 VSUBS 0.007257f
C135 B.n50 VSUBS 0.016183f
C136 B.n51 VSUBS 0.007257f
C137 B.n52 VSUBS 0.007257f
C138 B.n53 VSUBS 0.007257f
C139 B.n54 VSUBS 0.007257f
C140 B.n55 VSUBS 0.007257f
C141 B.n56 VSUBS 0.007257f
C142 B.n57 VSUBS 0.007257f
C143 B.n58 VSUBS 0.007257f
C144 B.n59 VSUBS 0.007257f
C145 B.t2 VSUBS 0.0664f
C146 B.t1 VSUBS 0.072792f
C147 B.t0 VSUBS 0.084962f
C148 B.n60 VSUBS 0.131863f
C149 B.n61 VSUBS 0.121526f
C150 B.n62 VSUBS 0.016815f
C151 B.n63 VSUBS 0.007257f
C152 B.n64 VSUBS 0.007257f
C153 B.n65 VSUBS 0.007257f
C154 B.n66 VSUBS 0.007257f
C155 B.n67 VSUBS 0.007257f
C156 B.t8 VSUBS 0.066399f
C157 B.t7 VSUBS 0.07279f
C158 B.t6 VSUBS 0.084962f
C159 B.n68 VSUBS 0.131864f
C160 B.n69 VSUBS 0.121527f
C161 B.n70 VSUBS 0.007257f
C162 B.n71 VSUBS 0.007257f
C163 B.n72 VSUBS 0.007257f
C164 B.n73 VSUBS 0.007257f
C165 B.n74 VSUBS 0.007257f
C166 B.n75 VSUBS 0.007257f
C167 B.n76 VSUBS 0.007257f
C168 B.n77 VSUBS 0.007257f
C169 B.n78 VSUBS 0.007257f
C170 B.n79 VSUBS 0.015787f
C171 B.n80 VSUBS 0.007257f
C172 B.n81 VSUBS 0.007257f
C173 B.n82 VSUBS 0.007257f
C174 B.n83 VSUBS 0.007257f
C175 B.n84 VSUBS 0.007257f
C176 B.n85 VSUBS 0.007257f
C177 B.n86 VSUBS 0.007257f
C178 B.n87 VSUBS 0.007257f
C179 B.n88 VSUBS 0.007257f
C180 B.n89 VSUBS 0.007257f
C181 B.n90 VSUBS 0.007257f
C182 B.n91 VSUBS 0.007257f
C183 B.n92 VSUBS 0.007257f
C184 B.n93 VSUBS 0.007257f
C185 B.n94 VSUBS 0.007257f
C186 B.n95 VSUBS 0.007257f
C187 B.n96 VSUBS 0.007257f
C188 B.n97 VSUBS 0.007257f
C189 B.n98 VSUBS 0.007257f
C190 B.n99 VSUBS 0.007257f
C191 B.n100 VSUBS 0.015787f
C192 B.n101 VSUBS 0.017084f
C193 B.n102 VSUBS 0.017084f
C194 B.n103 VSUBS 0.007257f
C195 B.n104 VSUBS 0.007257f
C196 B.n105 VSUBS 0.007257f
C197 B.n106 VSUBS 0.007257f
C198 B.n107 VSUBS 0.007257f
C199 B.n108 VSUBS 0.007257f
C200 B.n109 VSUBS 0.007257f
C201 B.n110 VSUBS 0.007257f
C202 B.n111 VSUBS 0.007257f
C203 B.n112 VSUBS 0.007257f
C204 B.n113 VSUBS 0.007257f
C205 B.n114 VSUBS 0.007257f
C206 B.n115 VSUBS 0.007257f
C207 B.n116 VSUBS 0.007257f
C208 B.n117 VSUBS 0.007257f
C209 B.n118 VSUBS 0.007257f
C210 B.n119 VSUBS 0.007257f
C211 B.n120 VSUBS 0.007257f
C212 B.n121 VSUBS 0.007257f
C213 B.n122 VSUBS 0.007257f
C214 B.n123 VSUBS 0.007257f
C215 B.n124 VSUBS 0.007257f
C216 B.n125 VSUBS 0.007257f
C217 B.n126 VSUBS 0.007257f
C218 B.n127 VSUBS 0.007257f
C219 B.n128 VSUBS 0.007257f
C220 B.n129 VSUBS 0.007257f
C221 B.n130 VSUBS 0.004803f
C222 B.n131 VSUBS 0.016815f
C223 B.n132 VSUBS 0.006083f
C224 B.n133 VSUBS 0.007257f
C225 B.n134 VSUBS 0.007257f
C226 B.n135 VSUBS 0.007257f
C227 B.n136 VSUBS 0.007257f
C228 B.n137 VSUBS 0.007257f
C229 B.n138 VSUBS 0.007257f
C230 B.n139 VSUBS 0.007257f
C231 B.n140 VSUBS 0.007257f
C232 B.n141 VSUBS 0.007257f
C233 B.n142 VSUBS 0.007257f
C234 B.n143 VSUBS 0.007257f
C235 B.n144 VSUBS 0.006083f
C236 B.n145 VSUBS 0.007257f
C237 B.n146 VSUBS 0.007257f
C238 B.n147 VSUBS 0.004803f
C239 B.n148 VSUBS 0.007257f
C240 B.n149 VSUBS 0.007257f
C241 B.n150 VSUBS 0.007257f
C242 B.n151 VSUBS 0.007257f
C243 B.n152 VSUBS 0.007257f
C244 B.n153 VSUBS 0.007257f
C245 B.n154 VSUBS 0.007257f
C246 B.n155 VSUBS 0.007257f
C247 B.n156 VSUBS 0.007257f
C248 B.n157 VSUBS 0.007257f
C249 B.n158 VSUBS 0.007257f
C250 B.n159 VSUBS 0.007257f
C251 B.n160 VSUBS 0.007257f
C252 B.n161 VSUBS 0.007257f
C253 B.n162 VSUBS 0.007257f
C254 B.n163 VSUBS 0.007257f
C255 B.n164 VSUBS 0.007257f
C256 B.n165 VSUBS 0.007257f
C257 B.n166 VSUBS 0.007257f
C258 B.n167 VSUBS 0.007257f
C259 B.n168 VSUBS 0.007257f
C260 B.n169 VSUBS 0.007257f
C261 B.n170 VSUBS 0.007257f
C262 B.n171 VSUBS 0.007257f
C263 B.n172 VSUBS 0.007257f
C264 B.n173 VSUBS 0.007257f
C265 B.n174 VSUBS 0.007257f
C266 B.n175 VSUBS 0.017084f
C267 B.n176 VSUBS 0.015787f
C268 B.n177 VSUBS 0.016689f
C269 B.n178 VSUBS 0.007257f
C270 B.n179 VSUBS 0.007257f
C271 B.n180 VSUBS 0.007257f
C272 B.n181 VSUBS 0.007257f
C273 B.n182 VSUBS 0.007257f
C274 B.n183 VSUBS 0.007257f
C275 B.n184 VSUBS 0.007257f
C276 B.n185 VSUBS 0.007257f
C277 B.n186 VSUBS 0.007257f
C278 B.n187 VSUBS 0.007257f
C279 B.n188 VSUBS 0.007257f
C280 B.n189 VSUBS 0.007257f
C281 B.n190 VSUBS 0.007257f
C282 B.n191 VSUBS 0.007257f
C283 B.n192 VSUBS 0.007257f
C284 B.n193 VSUBS 0.007257f
C285 B.n194 VSUBS 0.007257f
C286 B.n195 VSUBS 0.007257f
C287 B.n196 VSUBS 0.007257f
C288 B.n197 VSUBS 0.007257f
C289 B.n198 VSUBS 0.007257f
C290 B.n199 VSUBS 0.007257f
C291 B.n200 VSUBS 0.007257f
C292 B.n201 VSUBS 0.007257f
C293 B.n202 VSUBS 0.007257f
C294 B.n203 VSUBS 0.007257f
C295 B.n204 VSUBS 0.007257f
C296 B.n205 VSUBS 0.007257f
C297 B.n206 VSUBS 0.007257f
C298 B.n207 VSUBS 0.007257f
C299 B.n208 VSUBS 0.007257f
C300 B.n209 VSUBS 0.007257f
C301 B.n210 VSUBS 0.007257f
C302 B.n211 VSUBS 0.007257f
C303 B.n212 VSUBS 0.007257f
C304 B.n213 VSUBS 0.007257f
C305 B.n214 VSUBS 0.015787f
C306 B.n215 VSUBS 0.017084f
C307 B.n216 VSUBS 0.017084f
C308 B.n217 VSUBS 0.007257f
C309 B.n218 VSUBS 0.007257f
C310 B.n219 VSUBS 0.007257f
C311 B.n220 VSUBS 0.007257f
C312 B.n221 VSUBS 0.007257f
C313 B.n222 VSUBS 0.007257f
C314 B.n223 VSUBS 0.007257f
C315 B.n224 VSUBS 0.007257f
C316 B.n225 VSUBS 0.007257f
C317 B.n226 VSUBS 0.007257f
C318 B.n227 VSUBS 0.007257f
C319 B.n228 VSUBS 0.007257f
C320 B.n229 VSUBS 0.007257f
C321 B.n230 VSUBS 0.007257f
C322 B.n231 VSUBS 0.007257f
C323 B.n232 VSUBS 0.007257f
C324 B.n233 VSUBS 0.007257f
C325 B.n234 VSUBS 0.007257f
C326 B.n235 VSUBS 0.007257f
C327 B.n236 VSUBS 0.007257f
C328 B.n237 VSUBS 0.007257f
C329 B.n238 VSUBS 0.007257f
C330 B.n239 VSUBS 0.007257f
C331 B.n240 VSUBS 0.007257f
C332 B.n241 VSUBS 0.007257f
C333 B.n242 VSUBS 0.007257f
C334 B.n243 VSUBS 0.007257f
C335 B.n244 VSUBS 0.004803f
C336 B.n245 VSUBS 0.016815f
C337 B.n246 VSUBS 0.006083f
C338 B.n247 VSUBS 0.007257f
C339 B.n248 VSUBS 0.007257f
C340 B.n249 VSUBS 0.007257f
C341 B.n250 VSUBS 0.007257f
C342 B.n251 VSUBS 0.007257f
C343 B.n252 VSUBS 0.007257f
C344 B.n253 VSUBS 0.007257f
C345 B.n254 VSUBS 0.007257f
C346 B.n255 VSUBS 0.007257f
C347 B.n256 VSUBS 0.007257f
C348 B.n257 VSUBS 0.007257f
C349 B.n258 VSUBS 0.006083f
C350 B.n259 VSUBS 0.007257f
C351 B.n260 VSUBS 0.007257f
C352 B.n261 VSUBS 0.004803f
C353 B.n262 VSUBS 0.007257f
C354 B.n263 VSUBS 0.007257f
C355 B.n264 VSUBS 0.007257f
C356 B.n265 VSUBS 0.007257f
C357 B.n266 VSUBS 0.007257f
C358 B.n267 VSUBS 0.007257f
C359 B.n268 VSUBS 0.007257f
C360 B.n269 VSUBS 0.007257f
C361 B.n270 VSUBS 0.007257f
C362 B.n271 VSUBS 0.007257f
C363 B.n272 VSUBS 0.007257f
C364 B.n273 VSUBS 0.007257f
C365 B.n274 VSUBS 0.007257f
C366 B.n275 VSUBS 0.007257f
C367 B.n276 VSUBS 0.007257f
C368 B.n277 VSUBS 0.007257f
C369 B.n278 VSUBS 0.007257f
C370 B.n279 VSUBS 0.007257f
C371 B.n280 VSUBS 0.007257f
C372 B.n281 VSUBS 0.007257f
C373 B.n282 VSUBS 0.007257f
C374 B.n283 VSUBS 0.007257f
C375 B.n284 VSUBS 0.007257f
C376 B.n285 VSUBS 0.007257f
C377 B.n286 VSUBS 0.007257f
C378 B.n287 VSUBS 0.007257f
C379 B.n288 VSUBS 0.007257f
C380 B.n289 VSUBS 0.017084f
C381 B.n290 VSUBS 0.015787f
C382 B.n291 VSUBS 0.015787f
C383 B.n292 VSUBS 0.007257f
C384 B.n293 VSUBS 0.007257f
C385 B.n294 VSUBS 0.007257f
C386 B.n295 VSUBS 0.007257f
C387 B.n296 VSUBS 0.007257f
C388 B.n297 VSUBS 0.007257f
C389 B.n298 VSUBS 0.007257f
C390 B.n299 VSUBS 0.007257f
C391 B.n300 VSUBS 0.007257f
C392 B.n301 VSUBS 0.007257f
C393 B.n302 VSUBS 0.007257f
C394 B.n303 VSUBS 0.007257f
C395 B.n304 VSUBS 0.007257f
C396 B.n305 VSUBS 0.007257f
C397 B.n306 VSUBS 0.007257f
C398 B.n307 VSUBS 0.009471f
C399 B.n308 VSUBS 0.010088f
C400 B.n309 VSUBS 0.020062f
C401 VDD1.n0 VSUBS 0.017662f
C402 VDD1.n1 VSUBS 0.017344f
C403 VDD1.n2 VSUBS 0.00932f
C404 VDD1.n3 VSUBS 0.022029f
C405 VDD1.n4 VSUBS 0.009868f
C406 VDD1.n5 VSUBS 0.276113f
C407 VDD1.n6 VSUBS 0.00932f
C408 VDD1.t1 VSUBS 0.047562f
C409 VDD1.n7 VSUBS 0.068993f
C410 VDD1.n8 VSUBS 0.013956f
C411 VDD1.n9 VSUBS 0.016522f
C412 VDD1.n10 VSUBS 0.022029f
C413 VDD1.n11 VSUBS 0.009868f
C414 VDD1.n12 VSUBS 0.00932f
C415 VDD1.n13 VSUBS 0.017344f
C416 VDD1.n14 VSUBS 0.017344f
C417 VDD1.n15 VSUBS 0.00932f
C418 VDD1.n16 VSUBS 0.009868f
C419 VDD1.n17 VSUBS 0.022029f
C420 VDD1.n18 VSUBS 0.048575f
C421 VDD1.n19 VSUBS 0.009868f
C422 VDD1.n20 VSUBS 0.00932f
C423 VDD1.n21 VSUBS 0.037721f
C424 VDD1.n22 VSUBS 0.036347f
C425 VDD1.n23 VSUBS 0.017662f
C426 VDD1.n24 VSUBS 0.017344f
C427 VDD1.n25 VSUBS 0.00932f
C428 VDD1.n26 VSUBS 0.022029f
C429 VDD1.n27 VSUBS 0.009868f
C430 VDD1.n28 VSUBS 0.276113f
C431 VDD1.n29 VSUBS 0.00932f
C432 VDD1.t0 VSUBS 0.047562f
C433 VDD1.n30 VSUBS 0.068993f
C434 VDD1.n31 VSUBS 0.013956f
C435 VDD1.n32 VSUBS 0.016522f
C436 VDD1.n33 VSUBS 0.022029f
C437 VDD1.n34 VSUBS 0.009868f
C438 VDD1.n35 VSUBS 0.00932f
C439 VDD1.n36 VSUBS 0.017344f
C440 VDD1.n37 VSUBS 0.017344f
C441 VDD1.n38 VSUBS 0.00932f
C442 VDD1.n39 VSUBS 0.009868f
C443 VDD1.n40 VSUBS 0.022029f
C444 VDD1.n41 VSUBS 0.048575f
C445 VDD1.n42 VSUBS 0.009868f
C446 VDD1.n43 VSUBS 0.00932f
C447 VDD1.n44 VSUBS 0.037721f
C448 VDD1.n45 VSUBS 0.279174f
C449 VTAIL.n0 VSUBS 0.020742f
C450 VTAIL.n1 VSUBS 0.020369f
C451 VTAIL.n2 VSUBS 0.010945f
C452 VTAIL.n3 VSUBS 0.025871f
C453 VTAIL.n4 VSUBS 0.011589f
C454 VTAIL.n5 VSUBS 0.324262f
C455 VTAIL.n6 VSUBS 0.010945f
C456 VTAIL.t3 VSUBS 0.055857f
C457 VTAIL.n7 VSUBS 0.081024f
C458 VTAIL.n8 VSUBS 0.016389f
C459 VTAIL.n9 VSUBS 0.019403f
C460 VTAIL.n10 VSUBS 0.025871f
C461 VTAIL.n11 VSUBS 0.011589f
C462 VTAIL.n12 VSUBS 0.010945f
C463 VTAIL.n13 VSUBS 0.020369f
C464 VTAIL.n14 VSUBS 0.020369f
C465 VTAIL.n15 VSUBS 0.010945f
C466 VTAIL.n16 VSUBS 0.011589f
C467 VTAIL.n17 VSUBS 0.025871f
C468 VTAIL.n18 VSUBS 0.057046f
C469 VTAIL.n19 VSUBS 0.011589f
C470 VTAIL.n20 VSUBS 0.010945f
C471 VTAIL.n21 VSUBS 0.044299f
C472 VTAIL.n22 VSUBS 0.028352f
C473 VTAIL.n23 VSUBS 0.677396f
C474 VTAIL.n24 VSUBS 0.020742f
C475 VTAIL.n25 VSUBS 0.020369f
C476 VTAIL.n26 VSUBS 0.010945f
C477 VTAIL.n27 VSUBS 0.025871f
C478 VTAIL.n28 VSUBS 0.011589f
C479 VTAIL.n29 VSUBS 0.324262f
C480 VTAIL.n30 VSUBS 0.010945f
C481 VTAIL.t0 VSUBS 0.055857f
C482 VTAIL.n31 VSUBS 0.081024f
C483 VTAIL.n32 VSUBS 0.016389f
C484 VTAIL.n33 VSUBS 0.019403f
C485 VTAIL.n34 VSUBS 0.025871f
C486 VTAIL.n35 VSUBS 0.011589f
C487 VTAIL.n36 VSUBS 0.010945f
C488 VTAIL.n37 VSUBS 0.020369f
C489 VTAIL.n38 VSUBS 0.020369f
C490 VTAIL.n39 VSUBS 0.010945f
C491 VTAIL.n40 VSUBS 0.011589f
C492 VTAIL.n41 VSUBS 0.025871f
C493 VTAIL.n42 VSUBS 0.057046f
C494 VTAIL.n43 VSUBS 0.011589f
C495 VTAIL.n44 VSUBS 0.010945f
C496 VTAIL.n45 VSUBS 0.044299f
C497 VTAIL.n46 VSUBS 0.028352f
C498 VTAIL.n47 VSUBS 0.684327f
C499 VTAIL.n48 VSUBS 0.020742f
C500 VTAIL.n49 VSUBS 0.020369f
C501 VTAIL.n50 VSUBS 0.010945f
C502 VTAIL.n51 VSUBS 0.025871f
C503 VTAIL.n52 VSUBS 0.011589f
C504 VTAIL.n53 VSUBS 0.324262f
C505 VTAIL.n54 VSUBS 0.010945f
C506 VTAIL.t2 VSUBS 0.055857f
C507 VTAIL.n55 VSUBS 0.081024f
C508 VTAIL.n56 VSUBS 0.016389f
C509 VTAIL.n57 VSUBS 0.019403f
C510 VTAIL.n58 VSUBS 0.025871f
C511 VTAIL.n59 VSUBS 0.011589f
C512 VTAIL.n60 VSUBS 0.010945f
C513 VTAIL.n61 VSUBS 0.020369f
C514 VTAIL.n62 VSUBS 0.020369f
C515 VTAIL.n63 VSUBS 0.010945f
C516 VTAIL.n64 VSUBS 0.011589f
C517 VTAIL.n65 VSUBS 0.025871f
C518 VTAIL.n66 VSUBS 0.057046f
C519 VTAIL.n67 VSUBS 0.011589f
C520 VTAIL.n68 VSUBS 0.010945f
C521 VTAIL.n69 VSUBS 0.044299f
C522 VTAIL.n70 VSUBS 0.028352f
C523 VTAIL.n71 VSUBS 0.641326f
C524 VTAIL.n72 VSUBS 0.020742f
C525 VTAIL.n73 VSUBS 0.020369f
C526 VTAIL.n74 VSUBS 0.010945f
C527 VTAIL.n75 VSUBS 0.025871f
C528 VTAIL.n76 VSUBS 0.011589f
C529 VTAIL.n77 VSUBS 0.324262f
C530 VTAIL.n78 VSUBS 0.010945f
C531 VTAIL.t1 VSUBS 0.055857f
C532 VTAIL.n79 VSUBS 0.081024f
C533 VTAIL.n80 VSUBS 0.016389f
C534 VTAIL.n81 VSUBS 0.019403f
C535 VTAIL.n82 VSUBS 0.025871f
C536 VTAIL.n83 VSUBS 0.011589f
C537 VTAIL.n84 VSUBS 0.010945f
C538 VTAIL.n85 VSUBS 0.020369f
C539 VTAIL.n86 VSUBS 0.020369f
C540 VTAIL.n87 VSUBS 0.010945f
C541 VTAIL.n88 VSUBS 0.011589f
C542 VTAIL.n89 VSUBS 0.025871f
C543 VTAIL.n90 VSUBS 0.057046f
C544 VTAIL.n91 VSUBS 0.011589f
C545 VTAIL.n92 VSUBS 0.010945f
C546 VTAIL.n93 VSUBS 0.044299f
C547 VTAIL.n94 VSUBS 0.028352f
C548 VTAIL.n95 VSUBS 0.595921f
C549 VP.t0 VSUBS 0.347854f
C550 VP.t1 VSUBS 0.273264f
C551 VP.n0 VSUBS 2.37124f
.ends

