* NGSPICE file created from diff_pair_sample_0680.ext - technology: sky130A

.subckt diff_pair_sample_0680 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=2.43045 ps=15.06 w=14.73 l=3.66
X1 VDD1.t2 VP.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X2 VTAIL.t13 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X3 VDD2.t7 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=5.7447 ps=30.24 w=14.73 l=3.66
X4 VDD1.t4 VP.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X5 VDD1.t1 VP.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=5.7447 ps=30.24 w=14.73 l=3.66
X6 VTAIL.t10 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X7 VDD1.t7 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=5.7447 ps=30.24 w=14.73 l=3.66
X8 VDD2.t6 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X9 VTAIL.t7 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=2.43045 ps=15.06 w=14.73 l=3.66
X10 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X11 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
X12 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=0 ps=0 w=14.73 l=3.66
X13 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=2.43045 ps=15.06 w=14.73 l=3.66
X14 VDD2.t1 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=5.7447 ps=30.24 w=14.73 l=3.66
X15 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=0 ps=0 w=14.73 l=3.66
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=0 ps=0 w=14.73 l=3.66
X17 VTAIL.t8 VP.t7 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=2.43045 ps=15.06 w=14.73 l=3.66
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7447 pd=30.24 as=0 ps=0 w=14.73 l=3.66
X19 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.43045 pd=15.06 as=2.43045 ps=15.06 w=14.73 l=3.66
R0 VP.n22 VP.n19 161.3
R1 VP.n24 VP.n23 161.3
R2 VP.n25 VP.n18 161.3
R3 VP.n27 VP.n26 161.3
R4 VP.n28 VP.n17 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n31 VP.n16 161.3
R7 VP.n34 VP.n33 161.3
R8 VP.n35 VP.n15 161.3
R9 VP.n37 VP.n36 161.3
R10 VP.n38 VP.n14 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n41 VP.n13 161.3
R13 VP.n43 VP.n42 161.3
R14 VP.n44 VP.n12 161.3
R15 VP.n84 VP.n0 161.3
R16 VP.n83 VP.n82 161.3
R17 VP.n81 VP.n1 161.3
R18 VP.n80 VP.n79 161.3
R19 VP.n78 VP.n2 161.3
R20 VP.n77 VP.n76 161.3
R21 VP.n75 VP.n3 161.3
R22 VP.n74 VP.n73 161.3
R23 VP.n71 VP.n4 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n68 VP.n5 161.3
R26 VP.n67 VP.n66 161.3
R27 VP.n65 VP.n6 161.3
R28 VP.n64 VP.n63 161.3
R29 VP.n62 VP.n7 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n58 VP.n8 161.3
R32 VP.n57 VP.n56 161.3
R33 VP.n55 VP.n9 161.3
R34 VP.n54 VP.n53 161.3
R35 VP.n52 VP.n10 161.3
R36 VP.n51 VP.n50 161.3
R37 VP.n49 VP.n11 161.3
R38 VP.n21 VP.t0 129.172
R39 VP.n47 VP.t7 96.9931
R40 VP.n59 VP.t1 96.9931
R41 VP.n72 VP.t2 96.9931
R42 VP.n85 VP.t6 96.9931
R43 VP.n45 VP.t4 96.9931
R44 VP.n32 VP.t5 96.9931
R45 VP.n20 VP.t3 96.9931
R46 VP.n48 VP.n47 58.4488
R47 VP.n86 VP.n85 58.4488
R48 VP.n46 VP.n45 58.4488
R49 VP.n48 VP.n46 58.1404
R50 VP.n21 VP.n20 50.7163
R51 VP.n53 VP.n9 41.4647
R52 VP.n79 VP.n78 41.4647
R53 VP.n39 VP.n38 41.4647
R54 VP.n66 VP.n65 40.4934
R55 VP.n66 VP.n5 40.4934
R56 VP.n26 VP.n17 40.4934
R57 VP.n26 VP.n25 40.4934
R58 VP.n53 VP.n52 39.5221
R59 VP.n79 VP.n1 39.5221
R60 VP.n39 VP.n13 39.5221
R61 VP.n51 VP.n11 24.4675
R62 VP.n52 VP.n51 24.4675
R63 VP.n57 VP.n9 24.4675
R64 VP.n58 VP.n57 24.4675
R65 VP.n60 VP.n58 24.4675
R66 VP.n64 VP.n7 24.4675
R67 VP.n65 VP.n64 24.4675
R68 VP.n70 VP.n5 24.4675
R69 VP.n71 VP.n70 24.4675
R70 VP.n73 VP.n3 24.4675
R71 VP.n77 VP.n3 24.4675
R72 VP.n78 VP.n77 24.4675
R73 VP.n83 VP.n1 24.4675
R74 VP.n84 VP.n83 24.4675
R75 VP.n43 VP.n13 24.4675
R76 VP.n44 VP.n43 24.4675
R77 VP.n30 VP.n17 24.4675
R78 VP.n31 VP.n30 24.4675
R79 VP.n33 VP.n15 24.4675
R80 VP.n37 VP.n15 24.4675
R81 VP.n38 VP.n37 24.4675
R82 VP.n24 VP.n19 24.4675
R83 VP.n25 VP.n24 24.4675
R84 VP.n59 VP.n7 24.2228
R85 VP.n72 VP.n71 24.2228
R86 VP.n32 VP.n31 24.2228
R87 VP.n20 VP.n19 24.2228
R88 VP.n47 VP.n11 23.7335
R89 VP.n85 VP.n84 23.7335
R90 VP.n45 VP.n44 23.7335
R91 VP.n22 VP.n21 2.55161
R92 VP.n46 VP.n12 0.417535
R93 VP.n49 VP.n48 0.417535
R94 VP.n86 VP.n0 0.417535
R95 VP VP.n86 0.394291
R96 VP.n60 VP.n59 0.24517
R97 VP.n73 VP.n72 0.24517
R98 VP.n33 VP.n32 0.24517
R99 VP.n23 VP.n22 0.189894
R100 VP.n23 VP.n18 0.189894
R101 VP.n27 VP.n18 0.189894
R102 VP.n28 VP.n27 0.189894
R103 VP.n29 VP.n28 0.189894
R104 VP.n29 VP.n16 0.189894
R105 VP.n34 VP.n16 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n14 0.189894
R109 VP.n40 VP.n14 0.189894
R110 VP.n41 VP.n40 0.189894
R111 VP.n42 VP.n41 0.189894
R112 VP.n42 VP.n12 0.189894
R113 VP.n50 VP.n49 0.189894
R114 VP.n50 VP.n10 0.189894
R115 VP.n54 VP.n10 0.189894
R116 VP.n55 VP.n54 0.189894
R117 VP.n56 VP.n55 0.189894
R118 VP.n56 VP.n8 0.189894
R119 VP.n61 VP.n8 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n63 VP.n62 0.189894
R122 VP.n63 VP.n6 0.189894
R123 VP.n67 VP.n6 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n69 VP.n68 0.189894
R126 VP.n69 VP.n4 0.189894
R127 VP.n74 VP.n4 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n76 VP.n75 0.189894
R130 VP.n76 VP.n2 0.189894
R131 VP.n80 VP.n2 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n82 VP.n81 0.189894
R134 VP.n82 VP.n0 0.189894
R135 VDD1 VDD1.n0 64.4446
R136 VDD1.n3 VDD1.n2 64.3309
R137 VDD1.n3 VDD1.n1 64.3309
R138 VDD1.n5 VDD1.n4 62.6664
R139 VDD1.n5 VDD1.n3 52.475
R140 VDD1 VDD1.n5 1.66214
R141 VDD1.n4 VDD1.t0 1.3447
R142 VDD1.n4 VDD1.t1 1.3447
R143 VDD1.n0 VDD1.t3 1.3447
R144 VDD1.n0 VDD1.t4 1.3447
R145 VDD1.n2 VDD1.t5 1.3447
R146 VDD1.n2 VDD1.t7 1.3447
R147 VDD1.n1 VDD1.t6 1.3447
R148 VDD1.n1 VDD1.t2 1.3447
R149 VTAIL.n658 VTAIL.n582 289.615
R150 VTAIL.n78 VTAIL.n2 289.615
R151 VTAIL.n160 VTAIL.n84 289.615
R152 VTAIL.n244 VTAIL.n168 289.615
R153 VTAIL.n576 VTAIL.n500 289.615
R154 VTAIL.n492 VTAIL.n416 289.615
R155 VTAIL.n410 VTAIL.n334 289.615
R156 VTAIL.n326 VTAIL.n250 289.615
R157 VTAIL.n609 VTAIL.n608 185
R158 VTAIL.n606 VTAIL.n605 185
R159 VTAIL.n615 VTAIL.n614 185
R160 VTAIL.n617 VTAIL.n616 185
R161 VTAIL.n602 VTAIL.n601 185
R162 VTAIL.n623 VTAIL.n622 185
R163 VTAIL.n625 VTAIL.n624 185
R164 VTAIL.n598 VTAIL.n597 185
R165 VTAIL.n631 VTAIL.n630 185
R166 VTAIL.n633 VTAIL.n632 185
R167 VTAIL.n594 VTAIL.n593 185
R168 VTAIL.n639 VTAIL.n638 185
R169 VTAIL.n641 VTAIL.n640 185
R170 VTAIL.n590 VTAIL.n589 185
R171 VTAIL.n647 VTAIL.n646 185
R172 VTAIL.n650 VTAIL.n649 185
R173 VTAIL.n648 VTAIL.n586 185
R174 VTAIL.n655 VTAIL.n585 185
R175 VTAIL.n657 VTAIL.n656 185
R176 VTAIL.n659 VTAIL.n658 185
R177 VTAIL.n29 VTAIL.n28 185
R178 VTAIL.n26 VTAIL.n25 185
R179 VTAIL.n35 VTAIL.n34 185
R180 VTAIL.n37 VTAIL.n36 185
R181 VTAIL.n22 VTAIL.n21 185
R182 VTAIL.n43 VTAIL.n42 185
R183 VTAIL.n45 VTAIL.n44 185
R184 VTAIL.n18 VTAIL.n17 185
R185 VTAIL.n51 VTAIL.n50 185
R186 VTAIL.n53 VTAIL.n52 185
R187 VTAIL.n14 VTAIL.n13 185
R188 VTAIL.n59 VTAIL.n58 185
R189 VTAIL.n61 VTAIL.n60 185
R190 VTAIL.n10 VTAIL.n9 185
R191 VTAIL.n67 VTAIL.n66 185
R192 VTAIL.n70 VTAIL.n69 185
R193 VTAIL.n68 VTAIL.n6 185
R194 VTAIL.n75 VTAIL.n5 185
R195 VTAIL.n77 VTAIL.n76 185
R196 VTAIL.n79 VTAIL.n78 185
R197 VTAIL.n111 VTAIL.n110 185
R198 VTAIL.n108 VTAIL.n107 185
R199 VTAIL.n117 VTAIL.n116 185
R200 VTAIL.n119 VTAIL.n118 185
R201 VTAIL.n104 VTAIL.n103 185
R202 VTAIL.n125 VTAIL.n124 185
R203 VTAIL.n127 VTAIL.n126 185
R204 VTAIL.n100 VTAIL.n99 185
R205 VTAIL.n133 VTAIL.n132 185
R206 VTAIL.n135 VTAIL.n134 185
R207 VTAIL.n96 VTAIL.n95 185
R208 VTAIL.n141 VTAIL.n140 185
R209 VTAIL.n143 VTAIL.n142 185
R210 VTAIL.n92 VTAIL.n91 185
R211 VTAIL.n149 VTAIL.n148 185
R212 VTAIL.n152 VTAIL.n151 185
R213 VTAIL.n150 VTAIL.n88 185
R214 VTAIL.n157 VTAIL.n87 185
R215 VTAIL.n159 VTAIL.n158 185
R216 VTAIL.n161 VTAIL.n160 185
R217 VTAIL.n195 VTAIL.n194 185
R218 VTAIL.n192 VTAIL.n191 185
R219 VTAIL.n201 VTAIL.n200 185
R220 VTAIL.n203 VTAIL.n202 185
R221 VTAIL.n188 VTAIL.n187 185
R222 VTAIL.n209 VTAIL.n208 185
R223 VTAIL.n211 VTAIL.n210 185
R224 VTAIL.n184 VTAIL.n183 185
R225 VTAIL.n217 VTAIL.n216 185
R226 VTAIL.n219 VTAIL.n218 185
R227 VTAIL.n180 VTAIL.n179 185
R228 VTAIL.n225 VTAIL.n224 185
R229 VTAIL.n227 VTAIL.n226 185
R230 VTAIL.n176 VTAIL.n175 185
R231 VTAIL.n233 VTAIL.n232 185
R232 VTAIL.n236 VTAIL.n235 185
R233 VTAIL.n234 VTAIL.n172 185
R234 VTAIL.n241 VTAIL.n171 185
R235 VTAIL.n243 VTAIL.n242 185
R236 VTAIL.n245 VTAIL.n244 185
R237 VTAIL.n577 VTAIL.n576 185
R238 VTAIL.n575 VTAIL.n574 185
R239 VTAIL.n573 VTAIL.n503 185
R240 VTAIL.n507 VTAIL.n504 185
R241 VTAIL.n568 VTAIL.n567 185
R242 VTAIL.n566 VTAIL.n565 185
R243 VTAIL.n509 VTAIL.n508 185
R244 VTAIL.n560 VTAIL.n559 185
R245 VTAIL.n558 VTAIL.n557 185
R246 VTAIL.n513 VTAIL.n512 185
R247 VTAIL.n552 VTAIL.n551 185
R248 VTAIL.n550 VTAIL.n549 185
R249 VTAIL.n517 VTAIL.n516 185
R250 VTAIL.n544 VTAIL.n543 185
R251 VTAIL.n542 VTAIL.n541 185
R252 VTAIL.n521 VTAIL.n520 185
R253 VTAIL.n536 VTAIL.n535 185
R254 VTAIL.n534 VTAIL.n533 185
R255 VTAIL.n525 VTAIL.n524 185
R256 VTAIL.n528 VTAIL.n527 185
R257 VTAIL.n493 VTAIL.n492 185
R258 VTAIL.n491 VTAIL.n490 185
R259 VTAIL.n489 VTAIL.n419 185
R260 VTAIL.n423 VTAIL.n420 185
R261 VTAIL.n484 VTAIL.n483 185
R262 VTAIL.n482 VTAIL.n481 185
R263 VTAIL.n425 VTAIL.n424 185
R264 VTAIL.n476 VTAIL.n475 185
R265 VTAIL.n474 VTAIL.n473 185
R266 VTAIL.n429 VTAIL.n428 185
R267 VTAIL.n468 VTAIL.n467 185
R268 VTAIL.n466 VTAIL.n465 185
R269 VTAIL.n433 VTAIL.n432 185
R270 VTAIL.n460 VTAIL.n459 185
R271 VTAIL.n458 VTAIL.n457 185
R272 VTAIL.n437 VTAIL.n436 185
R273 VTAIL.n452 VTAIL.n451 185
R274 VTAIL.n450 VTAIL.n449 185
R275 VTAIL.n441 VTAIL.n440 185
R276 VTAIL.n444 VTAIL.n443 185
R277 VTAIL.n411 VTAIL.n410 185
R278 VTAIL.n409 VTAIL.n408 185
R279 VTAIL.n407 VTAIL.n337 185
R280 VTAIL.n341 VTAIL.n338 185
R281 VTAIL.n402 VTAIL.n401 185
R282 VTAIL.n400 VTAIL.n399 185
R283 VTAIL.n343 VTAIL.n342 185
R284 VTAIL.n394 VTAIL.n393 185
R285 VTAIL.n392 VTAIL.n391 185
R286 VTAIL.n347 VTAIL.n346 185
R287 VTAIL.n386 VTAIL.n385 185
R288 VTAIL.n384 VTAIL.n383 185
R289 VTAIL.n351 VTAIL.n350 185
R290 VTAIL.n378 VTAIL.n377 185
R291 VTAIL.n376 VTAIL.n375 185
R292 VTAIL.n355 VTAIL.n354 185
R293 VTAIL.n370 VTAIL.n369 185
R294 VTAIL.n368 VTAIL.n367 185
R295 VTAIL.n359 VTAIL.n358 185
R296 VTAIL.n362 VTAIL.n361 185
R297 VTAIL.n327 VTAIL.n326 185
R298 VTAIL.n325 VTAIL.n324 185
R299 VTAIL.n323 VTAIL.n253 185
R300 VTAIL.n257 VTAIL.n254 185
R301 VTAIL.n318 VTAIL.n317 185
R302 VTAIL.n316 VTAIL.n315 185
R303 VTAIL.n259 VTAIL.n258 185
R304 VTAIL.n310 VTAIL.n309 185
R305 VTAIL.n308 VTAIL.n307 185
R306 VTAIL.n263 VTAIL.n262 185
R307 VTAIL.n302 VTAIL.n301 185
R308 VTAIL.n300 VTAIL.n299 185
R309 VTAIL.n267 VTAIL.n266 185
R310 VTAIL.n294 VTAIL.n293 185
R311 VTAIL.n292 VTAIL.n291 185
R312 VTAIL.n271 VTAIL.n270 185
R313 VTAIL.n286 VTAIL.n285 185
R314 VTAIL.n284 VTAIL.n283 185
R315 VTAIL.n275 VTAIL.n274 185
R316 VTAIL.n278 VTAIL.n277 185
R317 VTAIL.t11 VTAIL.n526 147.659
R318 VTAIL.t15 VTAIL.n442 147.659
R319 VTAIL.t5 VTAIL.n360 147.659
R320 VTAIL.t7 VTAIL.n276 147.659
R321 VTAIL.t2 VTAIL.n607 147.659
R322 VTAIL.t1 VTAIL.n27 147.659
R323 VTAIL.t9 VTAIL.n109 147.659
R324 VTAIL.t8 VTAIL.n193 147.659
R325 VTAIL.n608 VTAIL.n605 104.615
R326 VTAIL.n615 VTAIL.n605 104.615
R327 VTAIL.n616 VTAIL.n615 104.615
R328 VTAIL.n616 VTAIL.n601 104.615
R329 VTAIL.n623 VTAIL.n601 104.615
R330 VTAIL.n624 VTAIL.n623 104.615
R331 VTAIL.n624 VTAIL.n597 104.615
R332 VTAIL.n631 VTAIL.n597 104.615
R333 VTAIL.n632 VTAIL.n631 104.615
R334 VTAIL.n632 VTAIL.n593 104.615
R335 VTAIL.n639 VTAIL.n593 104.615
R336 VTAIL.n640 VTAIL.n639 104.615
R337 VTAIL.n640 VTAIL.n589 104.615
R338 VTAIL.n647 VTAIL.n589 104.615
R339 VTAIL.n649 VTAIL.n647 104.615
R340 VTAIL.n649 VTAIL.n648 104.615
R341 VTAIL.n648 VTAIL.n585 104.615
R342 VTAIL.n657 VTAIL.n585 104.615
R343 VTAIL.n658 VTAIL.n657 104.615
R344 VTAIL.n28 VTAIL.n25 104.615
R345 VTAIL.n35 VTAIL.n25 104.615
R346 VTAIL.n36 VTAIL.n35 104.615
R347 VTAIL.n36 VTAIL.n21 104.615
R348 VTAIL.n43 VTAIL.n21 104.615
R349 VTAIL.n44 VTAIL.n43 104.615
R350 VTAIL.n44 VTAIL.n17 104.615
R351 VTAIL.n51 VTAIL.n17 104.615
R352 VTAIL.n52 VTAIL.n51 104.615
R353 VTAIL.n52 VTAIL.n13 104.615
R354 VTAIL.n59 VTAIL.n13 104.615
R355 VTAIL.n60 VTAIL.n59 104.615
R356 VTAIL.n60 VTAIL.n9 104.615
R357 VTAIL.n67 VTAIL.n9 104.615
R358 VTAIL.n69 VTAIL.n67 104.615
R359 VTAIL.n69 VTAIL.n68 104.615
R360 VTAIL.n68 VTAIL.n5 104.615
R361 VTAIL.n77 VTAIL.n5 104.615
R362 VTAIL.n78 VTAIL.n77 104.615
R363 VTAIL.n110 VTAIL.n107 104.615
R364 VTAIL.n117 VTAIL.n107 104.615
R365 VTAIL.n118 VTAIL.n117 104.615
R366 VTAIL.n118 VTAIL.n103 104.615
R367 VTAIL.n125 VTAIL.n103 104.615
R368 VTAIL.n126 VTAIL.n125 104.615
R369 VTAIL.n126 VTAIL.n99 104.615
R370 VTAIL.n133 VTAIL.n99 104.615
R371 VTAIL.n134 VTAIL.n133 104.615
R372 VTAIL.n134 VTAIL.n95 104.615
R373 VTAIL.n141 VTAIL.n95 104.615
R374 VTAIL.n142 VTAIL.n141 104.615
R375 VTAIL.n142 VTAIL.n91 104.615
R376 VTAIL.n149 VTAIL.n91 104.615
R377 VTAIL.n151 VTAIL.n149 104.615
R378 VTAIL.n151 VTAIL.n150 104.615
R379 VTAIL.n150 VTAIL.n87 104.615
R380 VTAIL.n159 VTAIL.n87 104.615
R381 VTAIL.n160 VTAIL.n159 104.615
R382 VTAIL.n194 VTAIL.n191 104.615
R383 VTAIL.n201 VTAIL.n191 104.615
R384 VTAIL.n202 VTAIL.n201 104.615
R385 VTAIL.n202 VTAIL.n187 104.615
R386 VTAIL.n209 VTAIL.n187 104.615
R387 VTAIL.n210 VTAIL.n209 104.615
R388 VTAIL.n210 VTAIL.n183 104.615
R389 VTAIL.n217 VTAIL.n183 104.615
R390 VTAIL.n218 VTAIL.n217 104.615
R391 VTAIL.n218 VTAIL.n179 104.615
R392 VTAIL.n225 VTAIL.n179 104.615
R393 VTAIL.n226 VTAIL.n225 104.615
R394 VTAIL.n226 VTAIL.n175 104.615
R395 VTAIL.n233 VTAIL.n175 104.615
R396 VTAIL.n235 VTAIL.n233 104.615
R397 VTAIL.n235 VTAIL.n234 104.615
R398 VTAIL.n234 VTAIL.n171 104.615
R399 VTAIL.n243 VTAIL.n171 104.615
R400 VTAIL.n244 VTAIL.n243 104.615
R401 VTAIL.n576 VTAIL.n575 104.615
R402 VTAIL.n575 VTAIL.n503 104.615
R403 VTAIL.n507 VTAIL.n503 104.615
R404 VTAIL.n567 VTAIL.n507 104.615
R405 VTAIL.n567 VTAIL.n566 104.615
R406 VTAIL.n566 VTAIL.n508 104.615
R407 VTAIL.n559 VTAIL.n508 104.615
R408 VTAIL.n559 VTAIL.n558 104.615
R409 VTAIL.n558 VTAIL.n512 104.615
R410 VTAIL.n551 VTAIL.n512 104.615
R411 VTAIL.n551 VTAIL.n550 104.615
R412 VTAIL.n550 VTAIL.n516 104.615
R413 VTAIL.n543 VTAIL.n516 104.615
R414 VTAIL.n543 VTAIL.n542 104.615
R415 VTAIL.n542 VTAIL.n520 104.615
R416 VTAIL.n535 VTAIL.n520 104.615
R417 VTAIL.n535 VTAIL.n534 104.615
R418 VTAIL.n534 VTAIL.n524 104.615
R419 VTAIL.n527 VTAIL.n524 104.615
R420 VTAIL.n492 VTAIL.n491 104.615
R421 VTAIL.n491 VTAIL.n419 104.615
R422 VTAIL.n423 VTAIL.n419 104.615
R423 VTAIL.n483 VTAIL.n423 104.615
R424 VTAIL.n483 VTAIL.n482 104.615
R425 VTAIL.n482 VTAIL.n424 104.615
R426 VTAIL.n475 VTAIL.n424 104.615
R427 VTAIL.n475 VTAIL.n474 104.615
R428 VTAIL.n474 VTAIL.n428 104.615
R429 VTAIL.n467 VTAIL.n428 104.615
R430 VTAIL.n467 VTAIL.n466 104.615
R431 VTAIL.n466 VTAIL.n432 104.615
R432 VTAIL.n459 VTAIL.n432 104.615
R433 VTAIL.n459 VTAIL.n458 104.615
R434 VTAIL.n458 VTAIL.n436 104.615
R435 VTAIL.n451 VTAIL.n436 104.615
R436 VTAIL.n451 VTAIL.n450 104.615
R437 VTAIL.n450 VTAIL.n440 104.615
R438 VTAIL.n443 VTAIL.n440 104.615
R439 VTAIL.n410 VTAIL.n409 104.615
R440 VTAIL.n409 VTAIL.n337 104.615
R441 VTAIL.n341 VTAIL.n337 104.615
R442 VTAIL.n401 VTAIL.n341 104.615
R443 VTAIL.n401 VTAIL.n400 104.615
R444 VTAIL.n400 VTAIL.n342 104.615
R445 VTAIL.n393 VTAIL.n342 104.615
R446 VTAIL.n393 VTAIL.n392 104.615
R447 VTAIL.n392 VTAIL.n346 104.615
R448 VTAIL.n385 VTAIL.n346 104.615
R449 VTAIL.n385 VTAIL.n384 104.615
R450 VTAIL.n384 VTAIL.n350 104.615
R451 VTAIL.n377 VTAIL.n350 104.615
R452 VTAIL.n377 VTAIL.n376 104.615
R453 VTAIL.n376 VTAIL.n354 104.615
R454 VTAIL.n369 VTAIL.n354 104.615
R455 VTAIL.n369 VTAIL.n368 104.615
R456 VTAIL.n368 VTAIL.n358 104.615
R457 VTAIL.n361 VTAIL.n358 104.615
R458 VTAIL.n326 VTAIL.n325 104.615
R459 VTAIL.n325 VTAIL.n253 104.615
R460 VTAIL.n257 VTAIL.n253 104.615
R461 VTAIL.n317 VTAIL.n257 104.615
R462 VTAIL.n317 VTAIL.n316 104.615
R463 VTAIL.n316 VTAIL.n258 104.615
R464 VTAIL.n309 VTAIL.n258 104.615
R465 VTAIL.n309 VTAIL.n308 104.615
R466 VTAIL.n308 VTAIL.n262 104.615
R467 VTAIL.n301 VTAIL.n262 104.615
R468 VTAIL.n301 VTAIL.n300 104.615
R469 VTAIL.n300 VTAIL.n266 104.615
R470 VTAIL.n293 VTAIL.n266 104.615
R471 VTAIL.n293 VTAIL.n292 104.615
R472 VTAIL.n292 VTAIL.n270 104.615
R473 VTAIL.n285 VTAIL.n270 104.615
R474 VTAIL.n285 VTAIL.n284 104.615
R475 VTAIL.n284 VTAIL.n274 104.615
R476 VTAIL.n277 VTAIL.n274 104.615
R477 VTAIL.n608 VTAIL.t2 52.3082
R478 VTAIL.n28 VTAIL.t1 52.3082
R479 VTAIL.n110 VTAIL.t9 52.3082
R480 VTAIL.n194 VTAIL.t8 52.3082
R481 VTAIL.n527 VTAIL.t11 52.3082
R482 VTAIL.n443 VTAIL.t15 52.3082
R483 VTAIL.n361 VTAIL.t5 52.3082
R484 VTAIL.n277 VTAIL.t7 52.3082
R485 VTAIL.n499 VTAIL.n498 45.9878
R486 VTAIL.n333 VTAIL.n332 45.9878
R487 VTAIL.n1 VTAIL.n0 45.9876
R488 VTAIL.n167 VTAIL.n166 45.9876
R489 VTAIL.n663 VTAIL.n662 33.9308
R490 VTAIL.n83 VTAIL.n82 33.9308
R491 VTAIL.n165 VTAIL.n164 33.9308
R492 VTAIL.n249 VTAIL.n248 33.9308
R493 VTAIL.n581 VTAIL.n580 33.9308
R494 VTAIL.n497 VTAIL.n496 33.9308
R495 VTAIL.n415 VTAIL.n414 33.9308
R496 VTAIL.n331 VTAIL.n330 33.9308
R497 VTAIL.n663 VTAIL.n581 28.5048
R498 VTAIL.n331 VTAIL.n249 28.5048
R499 VTAIL.n609 VTAIL.n607 15.6677
R500 VTAIL.n29 VTAIL.n27 15.6677
R501 VTAIL.n111 VTAIL.n109 15.6677
R502 VTAIL.n195 VTAIL.n193 15.6677
R503 VTAIL.n528 VTAIL.n526 15.6677
R504 VTAIL.n444 VTAIL.n442 15.6677
R505 VTAIL.n362 VTAIL.n360 15.6677
R506 VTAIL.n278 VTAIL.n276 15.6677
R507 VTAIL.n656 VTAIL.n655 13.1884
R508 VTAIL.n76 VTAIL.n75 13.1884
R509 VTAIL.n158 VTAIL.n157 13.1884
R510 VTAIL.n242 VTAIL.n241 13.1884
R511 VTAIL.n574 VTAIL.n573 13.1884
R512 VTAIL.n490 VTAIL.n489 13.1884
R513 VTAIL.n408 VTAIL.n407 13.1884
R514 VTAIL.n324 VTAIL.n323 13.1884
R515 VTAIL.n610 VTAIL.n606 12.8005
R516 VTAIL.n654 VTAIL.n586 12.8005
R517 VTAIL.n659 VTAIL.n584 12.8005
R518 VTAIL.n30 VTAIL.n26 12.8005
R519 VTAIL.n74 VTAIL.n6 12.8005
R520 VTAIL.n79 VTAIL.n4 12.8005
R521 VTAIL.n112 VTAIL.n108 12.8005
R522 VTAIL.n156 VTAIL.n88 12.8005
R523 VTAIL.n161 VTAIL.n86 12.8005
R524 VTAIL.n196 VTAIL.n192 12.8005
R525 VTAIL.n240 VTAIL.n172 12.8005
R526 VTAIL.n245 VTAIL.n170 12.8005
R527 VTAIL.n577 VTAIL.n502 12.8005
R528 VTAIL.n572 VTAIL.n504 12.8005
R529 VTAIL.n529 VTAIL.n525 12.8005
R530 VTAIL.n493 VTAIL.n418 12.8005
R531 VTAIL.n488 VTAIL.n420 12.8005
R532 VTAIL.n445 VTAIL.n441 12.8005
R533 VTAIL.n411 VTAIL.n336 12.8005
R534 VTAIL.n406 VTAIL.n338 12.8005
R535 VTAIL.n363 VTAIL.n359 12.8005
R536 VTAIL.n327 VTAIL.n252 12.8005
R537 VTAIL.n322 VTAIL.n254 12.8005
R538 VTAIL.n279 VTAIL.n275 12.8005
R539 VTAIL.n614 VTAIL.n613 12.0247
R540 VTAIL.n651 VTAIL.n650 12.0247
R541 VTAIL.n660 VTAIL.n582 12.0247
R542 VTAIL.n34 VTAIL.n33 12.0247
R543 VTAIL.n71 VTAIL.n70 12.0247
R544 VTAIL.n80 VTAIL.n2 12.0247
R545 VTAIL.n116 VTAIL.n115 12.0247
R546 VTAIL.n153 VTAIL.n152 12.0247
R547 VTAIL.n162 VTAIL.n84 12.0247
R548 VTAIL.n200 VTAIL.n199 12.0247
R549 VTAIL.n237 VTAIL.n236 12.0247
R550 VTAIL.n246 VTAIL.n168 12.0247
R551 VTAIL.n578 VTAIL.n500 12.0247
R552 VTAIL.n569 VTAIL.n568 12.0247
R553 VTAIL.n533 VTAIL.n532 12.0247
R554 VTAIL.n494 VTAIL.n416 12.0247
R555 VTAIL.n485 VTAIL.n484 12.0247
R556 VTAIL.n449 VTAIL.n448 12.0247
R557 VTAIL.n412 VTAIL.n334 12.0247
R558 VTAIL.n403 VTAIL.n402 12.0247
R559 VTAIL.n367 VTAIL.n366 12.0247
R560 VTAIL.n328 VTAIL.n250 12.0247
R561 VTAIL.n319 VTAIL.n318 12.0247
R562 VTAIL.n283 VTAIL.n282 12.0247
R563 VTAIL.n617 VTAIL.n604 11.249
R564 VTAIL.n646 VTAIL.n588 11.249
R565 VTAIL.n37 VTAIL.n24 11.249
R566 VTAIL.n66 VTAIL.n8 11.249
R567 VTAIL.n119 VTAIL.n106 11.249
R568 VTAIL.n148 VTAIL.n90 11.249
R569 VTAIL.n203 VTAIL.n190 11.249
R570 VTAIL.n232 VTAIL.n174 11.249
R571 VTAIL.n565 VTAIL.n506 11.249
R572 VTAIL.n536 VTAIL.n523 11.249
R573 VTAIL.n481 VTAIL.n422 11.249
R574 VTAIL.n452 VTAIL.n439 11.249
R575 VTAIL.n399 VTAIL.n340 11.249
R576 VTAIL.n370 VTAIL.n357 11.249
R577 VTAIL.n315 VTAIL.n256 11.249
R578 VTAIL.n286 VTAIL.n273 11.249
R579 VTAIL.n618 VTAIL.n602 10.4732
R580 VTAIL.n645 VTAIL.n590 10.4732
R581 VTAIL.n38 VTAIL.n22 10.4732
R582 VTAIL.n65 VTAIL.n10 10.4732
R583 VTAIL.n120 VTAIL.n104 10.4732
R584 VTAIL.n147 VTAIL.n92 10.4732
R585 VTAIL.n204 VTAIL.n188 10.4732
R586 VTAIL.n231 VTAIL.n176 10.4732
R587 VTAIL.n564 VTAIL.n509 10.4732
R588 VTAIL.n537 VTAIL.n521 10.4732
R589 VTAIL.n480 VTAIL.n425 10.4732
R590 VTAIL.n453 VTAIL.n437 10.4732
R591 VTAIL.n398 VTAIL.n343 10.4732
R592 VTAIL.n371 VTAIL.n355 10.4732
R593 VTAIL.n314 VTAIL.n259 10.4732
R594 VTAIL.n287 VTAIL.n271 10.4732
R595 VTAIL.n622 VTAIL.n621 9.69747
R596 VTAIL.n642 VTAIL.n641 9.69747
R597 VTAIL.n42 VTAIL.n41 9.69747
R598 VTAIL.n62 VTAIL.n61 9.69747
R599 VTAIL.n124 VTAIL.n123 9.69747
R600 VTAIL.n144 VTAIL.n143 9.69747
R601 VTAIL.n208 VTAIL.n207 9.69747
R602 VTAIL.n228 VTAIL.n227 9.69747
R603 VTAIL.n561 VTAIL.n560 9.69747
R604 VTAIL.n541 VTAIL.n540 9.69747
R605 VTAIL.n477 VTAIL.n476 9.69747
R606 VTAIL.n457 VTAIL.n456 9.69747
R607 VTAIL.n395 VTAIL.n394 9.69747
R608 VTAIL.n375 VTAIL.n374 9.69747
R609 VTAIL.n311 VTAIL.n310 9.69747
R610 VTAIL.n291 VTAIL.n290 9.69747
R611 VTAIL.n662 VTAIL.n661 9.45567
R612 VTAIL.n82 VTAIL.n81 9.45567
R613 VTAIL.n164 VTAIL.n163 9.45567
R614 VTAIL.n248 VTAIL.n247 9.45567
R615 VTAIL.n580 VTAIL.n579 9.45567
R616 VTAIL.n496 VTAIL.n495 9.45567
R617 VTAIL.n414 VTAIL.n413 9.45567
R618 VTAIL.n330 VTAIL.n329 9.45567
R619 VTAIL.n661 VTAIL.n660 9.3005
R620 VTAIL.n584 VTAIL.n583 9.3005
R621 VTAIL.n629 VTAIL.n628 9.3005
R622 VTAIL.n627 VTAIL.n626 9.3005
R623 VTAIL.n600 VTAIL.n599 9.3005
R624 VTAIL.n621 VTAIL.n620 9.3005
R625 VTAIL.n619 VTAIL.n618 9.3005
R626 VTAIL.n604 VTAIL.n603 9.3005
R627 VTAIL.n613 VTAIL.n612 9.3005
R628 VTAIL.n611 VTAIL.n610 9.3005
R629 VTAIL.n596 VTAIL.n595 9.3005
R630 VTAIL.n635 VTAIL.n634 9.3005
R631 VTAIL.n637 VTAIL.n636 9.3005
R632 VTAIL.n592 VTAIL.n591 9.3005
R633 VTAIL.n643 VTAIL.n642 9.3005
R634 VTAIL.n645 VTAIL.n644 9.3005
R635 VTAIL.n588 VTAIL.n587 9.3005
R636 VTAIL.n652 VTAIL.n651 9.3005
R637 VTAIL.n654 VTAIL.n653 9.3005
R638 VTAIL.n81 VTAIL.n80 9.3005
R639 VTAIL.n4 VTAIL.n3 9.3005
R640 VTAIL.n49 VTAIL.n48 9.3005
R641 VTAIL.n47 VTAIL.n46 9.3005
R642 VTAIL.n20 VTAIL.n19 9.3005
R643 VTAIL.n41 VTAIL.n40 9.3005
R644 VTAIL.n39 VTAIL.n38 9.3005
R645 VTAIL.n24 VTAIL.n23 9.3005
R646 VTAIL.n33 VTAIL.n32 9.3005
R647 VTAIL.n31 VTAIL.n30 9.3005
R648 VTAIL.n16 VTAIL.n15 9.3005
R649 VTAIL.n55 VTAIL.n54 9.3005
R650 VTAIL.n57 VTAIL.n56 9.3005
R651 VTAIL.n12 VTAIL.n11 9.3005
R652 VTAIL.n63 VTAIL.n62 9.3005
R653 VTAIL.n65 VTAIL.n64 9.3005
R654 VTAIL.n8 VTAIL.n7 9.3005
R655 VTAIL.n72 VTAIL.n71 9.3005
R656 VTAIL.n74 VTAIL.n73 9.3005
R657 VTAIL.n163 VTAIL.n162 9.3005
R658 VTAIL.n86 VTAIL.n85 9.3005
R659 VTAIL.n131 VTAIL.n130 9.3005
R660 VTAIL.n129 VTAIL.n128 9.3005
R661 VTAIL.n102 VTAIL.n101 9.3005
R662 VTAIL.n123 VTAIL.n122 9.3005
R663 VTAIL.n121 VTAIL.n120 9.3005
R664 VTAIL.n106 VTAIL.n105 9.3005
R665 VTAIL.n115 VTAIL.n114 9.3005
R666 VTAIL.n113 VTAIL.n112 9.3005
R667 VTAIL.n98 VTAIL.n97 9.3005
R668 VTAIL.n137 VTAIL.n136 9.3005
R669 VTAIL.n139 VTAIL.n138 9.3005
R670 VTAIL.n94 VTAIL.n93 9.3005
R671 VTAIL.n145 VTAIL.n144 9.3005
R672 VTAIL.n147 VTAIL.n146 9.3005
R673 VTAIL.n90 VTAIL.n89 9.3005
R674 VTAIL.n154 VTAIL.n153 9.3005
R675 VTAIL.n156 VTAIL.n155 9.3005
R676 VTAIL.n247 VTAIL.n246 9.3005
R677 VTAIL.n170 VTAIL.n169 9.3005
R678 VTAIL.n215 VTAIL.n214 9.3005
R679 VTAIL.n213 VTAIL.n212 9.3005
R680 VTAIL.n186 VTAIL.n185 9.3005
R681 VTAIL.n207 VTAIL.n206 9.3005
R682 VTAIL.n205 VTAIL.n204 9.3005
R683 VTAIL.n190 VTAIL.n189 9.3005
R684 VTAIL.n199 VTAIL.n198 9.3005
R685 VTAIL.n197 VTAIL.n196 9.3005
R686 VTAIL.n182 VTAIL.n181 9.3005
R687 VTAIL.n221 VTAIL.n220 9.3005
R688 VTAIL.n223 VTAIL.n222 9.3005
R689 VTAIL.n178 VTAIL.n177 9.3005
R690 VTAIL.n229 VTAIL.n228 9.3005
R691 VTAIL.n231 VTAIL.n230 9.3005
R692 VTAIL.n174 VTAIL.n173 9.3005
R693 VTAIL.n238 VTAIL.n237 9.3005
R694 VTAIL.n240 VTAIL.n239 9.3005
R695 VTAIL.n554 VTAIL.n553 9.3005
R696 VTAIL.n556 VTAIL.n555 9.3005
R697 VTAIL.n511 VTAIL.n510 9.3005
R698 VTAIL.n562 VTAIL.n561 9.3005
R699 VTAIL.n564 VTAIL.n563 9.3005
R700 VTAIL.n506 VTAIL.n505 9.3005
R701 VTAIL.n570 VTAIL.n569 9.3005
R702 VTAIL.n572 VTAIL.n571 9.3005
R703 VTAIL.n579 VTAIL.n578 9.3005
R704 VTAIL.n502 VTAIL.n501 9.3005
R705 VTAIL.n515 VTAIL.n514 9.3005
R706 VTAIL.n548 VTAIL.n547 9.3005
R707 VTAIL.n546 VTAIL.n545 9.3005
R708 VTAIL.n519 VTAIL.n518 9.3005
R709 VTAIL.n540 VTAIL.n539 9.3005
R710 VTAIL.n538 VTAIL.n537 9.3005
R711 VTAIL.n523 VTAIL.n522 9.3005
R712 VTAIL.n532 VTAIL.n531 9.3005
R713 VTAIL.n530 VTAIL.n529 9.3005
R714 VTAIL.n470 VTAIL.n469 9.3005
R715 VTAIL.n472 VTAIL.n471 9.3005
R716 VTAIL.n427 VTAIL.n426 9.3005
R717 VTAIL.n478 VTAIL.n477 9.3005
R718 VTAIL.n480 VTAIL.n479 9.3005
R719 VTAIL.n422 VTAIL.n421 9.3005
R720 VTAIL.n486 VTAIL.n485 9.3005
R721 VTAIL.n488 VTAIL.n487 9.3005
R722 VTAIL.n495 VTAIL.n494 9.3005
R723 VTAIL.n418 VTAIL.n417 9.3005
R724 VTAIL.n431 VTAIL.n430 9.3005
R725 VTAIL.n464 VTAIL.n463 9.3005
R726 VTAIL.n462 VTAIL.n461 9.3005
R727 VTAIL.n435 VTAIL.n434 9.3005
R728 VTAIL.n456 VTAIL.n455 9.3005
R729 VTAIL.n454 VTAIL.n453 9.3005
R730 VTAIL.n439 VTAIL.n438 9.3005
R731 VTAIL.n448 VTAIL.n447 9.3005
R732 VTAIL.n446 VTAIL.n445 9.3005
R733 VTAIL.n388 VTAIL.n387 9.3005
R734 VTAIL.n390 VTAIL.n389 9.3005
R735 VTAIL.n345 VTAIL.n344 9.3005
R736 VTAIL.n396 VTAIL.n395 9.3005
R737 VTAIL.n398 VTAIL.n397 9.3005
R738 VTAIL.n340 VTAIL.n339 9.3005
R739 VTAIL.n404 VTAIL.n403 9.3005
R740 VTAIL.n406 VTAIL.n405 9.3005
R741 VTAIL.n413 VTAIL.n412 9.3005
R742 VTAIL.n336 VTAIL.n335 9.3005
R743 VTAIL.n349 VTAIL.n348 9.3005
R744 VTAIL.n382 VTAIL.n381 9.3005
R745 VTAIL.n380 VTAIL.n379 9.3005
R746 VTAIL.n353 VTAIL.n352 9.3005
R747 VTAIL.n374 VTAIL.n373 9.3005
R748 VTAIL.n372 VTAIL.n371 9.3005
R749 VTAIL.n357 VTAIL.n356 9.3005
R750 VTAIL.n366 VTAIL.n365 9.3005
R751 VTAIL.n364 VTAIL.n363 9.3005
R752 VTAIL.n304 VTAIL.n303 9.3005
R753 VTAIL.n306 VTAIL.n305 9.3005
R754 VTAIL.n261 VTAIL.n260 9.3005
R755 VTAIL.n312 VTAIL.n311 9.3005
R756 VTAIL.n314 VTAIL.n313 9.3005
R757 VTAIL.n256 VTAIL.n255 9.3005
R758 VTAIL.n320 VTAIL.n319 9.3005
R759 VTAIL.n322 VTAIL.n321 9.3005
R760 VTAIL.n329 VTAIL.n328 9.3005
R761 VTAIL.n252 VTAIL.n251 9.3005
R762 VTAIL.n265 VTAIL.n264 9.3005
R763 VTAIL.n298 VTAIL.n297 9.3005
R764 VTAIL.n296 VTAIL.n295 9.3005
R765 VTAIL.n269 VTAIL.n268 9.3005
R766 VTAIL.n290 VTAIL.n289 9.3005
R767 VTAIL.n288 VTAIL.n287 9.3005
R768 VTAIL.n273 VTAIL.n272 9.3005
R769 VTAIL.n282 VTAIL.n281 9.3005
R770 VTAIL.n280 VTAIL.n279 9.3005
R771 VTAIL.n625 VTAIL.n600 8.92171
R772 VTAIL.n638 VTAIL.n592 8.92171
R773 VTAIL.n45 VTAIL.n20 8.92171
R774 VTAIL.n58 VTAIL.n12 8.92171
R775 VTAIL.n127 VTAIL.n102 8.92171
R776 VTAIL.n140 VTAIL.n94 8.92171
R777 VTAIL.n211 VTAIL.n186 8.92171
R778 VTAIL.n224 VTAIL.n178 8.92171
R779 VTAIL.n557 VTAIL.n511 8.92171
R780 VTAIL.n544 VTAIL.n519 8.92171
R781 VTAIL.n473 VTAIL.n427 8.92171
R782 VTAIL.n460 VTAIL.n435 8.92171
R783 VTAIL.n391 VTAIL.n345 8.92171
R784 VTAIL.n378 VTAIL.n353 8.92171
R785 VTAIL.n307 VTAIL.n261 8.92171
R786 VTAIL.n294 VTAIL.n269 8.92171
R787 VTAIL.n626 VTAIL.n598 8.14595
R788 VTAIL.n637 VTAIL.n594 8.14595
R789 VTAIL.n46 VTAIL.n18 8.14595
R790 VTAIL.n57 VTAIL.n14 8.14595
R791 VTAIL.n128 VTAIL.n100 8.14595
R792 VTAIL.n139 VTAIL.n96 8.14595
R793 VTAIL.n212 VTAIL.n184 8.14595
R794 VTAIL.n223 VTAIL.n180 8.14595
R795 VTAIL.n556 VTAIL.n513 8.14595
R796 VTAIL.n545 VTAIL.n517 8.14595
R797 VTAIL.n472 VTAIL.n429 8.14595
R798 VTAIL.n461 VTAIL.n433 8.14595
R799 VTAIL.n390 VTAIL.n347 8.14595
R800 VTAIL.n379 VTAIL.n351 8.14595
R801 VTAIL.n306 VTAIL.n263 8.14595
R802 VTAIL.n295 VTAIL.n267 8.14595
R803 VTAIL.n630 VTAIL.n629 7.3702
R804 VTAIL.n634 VTAIL.n633 7.3702
R805 VTAIL.n50 VTAIL.n49 7.3702
R806 VTAIL.n54 VTAIL.n53 7.3702
R807 VTAIL.n132 VTAIL.n131 7.3702
R808 VTAIL.n136 VTAIL.n135 7.3702
R809 VTAIL.n216 VTAIL.n215 7.3702
R810 VTAIL.n220 VTAIL.n219 7.3702
R811 VTAIL.n553 VTAIL.n552 7.3702
R812 VTAIL.n549 VTAIL.n548 7.3702
R813 VTAIL.n469 VTAIL.n468 7.3702
R814 VTAIL.n465 VTAIL.n464 7.3702
R815 VTAIL.n387 VTAIL.n386 7.3702
R816 VTAIL.n383 VTAIL.n382 7.3702
R817 VTAIL.n303 VTAIL.n302 7.3702
R818 VTAIL.n299 VTAIL.n298 7.3702
R819 VTAIL.n630 VTAIL.n596 6.59444
R820 VTAIL.n633 VTAIL.n596 6.59444
R821 VTAIL.n50 VTAIL.n16 6.59444
R822 VTAIL.n53 VTAIL.n16 6.59444
R823 VTAIL.n132 VTAIL.n98 6.59444
R824 VTAIL.n135 VTAIL.n98 6.59444
R825 VTAIL.n216 VTAIL.n182 6.59444
R826 VTAIL.n219 VTAIL.n182 6.59444
R827 VTAIL.n552 VTAIL.n515 6.59444
R828 VTAIL.n549 VTAIL.n515 6.59444
R829 VTAIL.n468 VTAIL.n431 6.59444
R830 VTAIL.n465 VTAIL.n431 6.59444
R831 VTAIL.n386 VTAIL.n349 6.59444
R832 VTAIL.n383 VTAIL.n349 6.59444
R833 VTAIL.n302 VTAIL.n265 6.59444
R834 VTAIL.n299 VTAIL.n265 6.59444
R835 VTAIL.n629 VTAIL.n598 5.81868
R836 VTAIL.n634 VTAIL.n594 5.81868
R837 VTAIL.n49 VTAIL.n18 5.81868
R838 VTAIL.n54 VTAIL.n14 5.81868
R839 VTAIL.n131 VTAIL.n100 5.81868
R840 VTAIL.n136 VTAIL.n96 5.81868
R841 VTAIL.n215 VTAIL.n184 5.81868
R842 VTAIL.n220 VTAIL.n180 5.81868
R843 VTAIL.n553 VTAIL.n513 5.81868
R844 VTAIL.n548 VTAIL.n517 5.81868
R845 VTAIL.n469 VTAIL.n429 5.81868
R846 VTAIL.n464 VTAIL.n433 5.81868
R847 VTAIL.n387 VTAIL.n347 5.81868
R848 VTAIL.n382 VTAIL.n351 5.81868
R849 VTAIL.n303 VTAIL.n263 5.81868
R850 VTAIL.n298 VTAIL.n267 5.81868
R851 VTAIL.n626 VTAIL.n625 5.04292
R852 VTAIL.n638 VTAIL.n637 5.04292
R853 VTAIL.n46 VTAIL.n45 5.04292
R854 VTAIL.n58 VTAIL.n57 5.04292
R855 VTAIL.n128 VTAIL.n127 5.04292
R856 VTAIL.n140 VTAIL.n139 5.04292
R857 VTAIL.n212 VTAIL.n211 5.04292
R858 VTAIL.n224 VTAIL.n223 5.04292
R859 VTAIL.n557 VTAIL.n556 5.04292
R860 VTAIL.n545 VTAIL.n544 5.04292
R861 VTAIL.n473 VTAIL.n472 5.04292
R862 VTAIL.n461 VTAIL.n460 5.04292
R863 VTAIL.n391 VTAIL.n390 5.04292
R864 VTAIL.n379 VTAIL.n378 5.04292
R865 VTAIL.n307 VTAIL.n306 5.04292
R866 VTAIL.n295 VTAIL.n294 5.04292
R867 VTAIL.n530 VTAIL.n526 4.38563
R868 VTAIL.n446 VTAIL.n442 4.38563
R869 VTAIL.n364 VTAIL.n360 4.38563
R870 VTAIL.n280 VTAIL.n276 4.38563
R871 VTAIL.n611 VTAIL.n607 4.38563
R872 VTAIL.n31 VTAIL.n27 4.38563
R873 VTAIL.n113 VTAIL.n109 4.38563
R874 VTAIL.n197 VTAIL.n193 4.38563
R875 VTAIL.n622 VTAIL.n600 4.26717
R876 VTAIL.n641 VTAIL.n592 4.26717
R877 VTAIL.n42 VTAIL.n20 4.26717
R878 VTAIL.n61 VTAIL.n12 4.26717
R879 VTAIL.n124 VTAIL.n102 4.26717
R880 VTAIL.n143 VTAIL.n94 4.26717
R881 VTAIL.n208 VTAIL.n186 4.26717
R882 VTAIL.n227 VTAIL.n178 4.26717
R883 VTAIL.n560 VTAIL.n511 4.26717
R884 VTAIL.n541 VTAIL.n519 4.26717
R885 VTAIL.n476 VTAIL.n427 4.26717
R886 VTAIL.n457 VTAIL.n435 4.26717
R887 VTAIL.n394 VTAIL.n345 4.26717
R888 VTAIL.n375 VTAIL.n353 4.26717
R889 VTAIL.n310 VTAIL.n261 4.26717
R890 VTAIL.n291 VTAIL.n269 4.26717
R891 VTAIL.n621 VTAIL.n602 3.49141
R892 VTAIL.n642 VTAIL.n590 3.49141
R893 VTAIL.n41 VTAIL.n22 3.49141
R894 VTAIL.n62 VTAIL.n10 3.49141
R895 VTAIL.n123 VTAIL.n104 3.49141
R896 VTAIL.n144 VTAIL.n92 3.49141
R897 VTAIL.n207 VTAIL.n188 3.49141
R898 VTAIL.n228 VTAIL.n176 3.49141
R899 VTAIL.n561 VTAIL.n509 3.49141
R900 VTAIL.n540 VTAIL.n521 3.49141
R901 VTAIL.n477 VTAIL.n425 3.49141
R902 VTAIL.n456 VTAIL.n437 3.49141
R903 VTAIL.n395 VTAIL.n343 3.49141
R904 VTAIL.n374 VTAIL.n355 3.49141
R905 VTAIL.n311 VTAIL.n259 3.49141
R906 VTAIL.n290 VTAIL.n271 3.49141
R907 VTAIL.n333 VTAIL.n331 3.44016
R908 VTAIL.n415 VTAIL.n333 3.44016
R909 VTAIL.n499 VTAIL.n497 3.44016
R910 VTAIL.n581 VTAIL.n499 3.44016
R911 VTAIL.n249 VTAIL.n167 3.44016
R912 VTAIL.n167 VTAIL.n165 3.44016
R913 VTAIL.n83 VTAIL.n1 3.44016
R914 VTAIL VTAIL.n663 3.38197
R915 VTAIL.n618 VTAIL.n617 2.71565
R916 VTAIL.n646 VTAIL.n645 2.71565
R917 VTAIL.n38 VTAIL.n37 2.71565
R918 VTAIL.n66 VTAIL.n65 2.71565
R919 VTAIL.n120 VTAIL.n119 2.71565
R920 VTAIL.n148 VTAIL.n147 2.71565
R921 VTAIL.n204 VTAIL.n203 2.71565
R922 VTAIL.n232 VTAIL.n231 2.71565
R923 VTAIL.n565 VTAIL.n564 2.71565
R924 VTAIL.n537 VTAIL.n536 2.71565
R925 VTAIL.n481 VTAIL.n480 2.71565
R926 VTAIL.n453 VTAIL.n452 2.71565
R927 VTAIL.n399 VTAIL.n398 2.71565
R928 VTAIL.n371 VTAIL.n370 2.71565
R929 VTAIL.n315 VTAIL.n314 2.71565
R930 VTAIL.n287 VTAIL.n286 2.71565
R931 VTAIL.n614 VTAIL.n604 1.93989
R932 VTAIL.n650 VTAIL.n588 1.93989
R933 VTAIL.n662 VTAIL.n582 1.93989
R934 VTAIL.n34 VTAIL.n24 1.93989
R935 VTAIL.n70 VTAIL.n8 1.93989
R936 VTAIL.n82 VTAIL.n2 1.93989
R937 VTAIL.n116 VTAIL.n106 1.93989
R938 VTAIL.n152 VTAIL.n90 1.93989
R939 VTAIL.n164 VTAIL.n84 1.93989
R940 VTAIL.n200 VTAIL.n190 1.93989
R941 VTAIL.n236 VTAIL.n174 1.93989
R942 VTAIL.n248 VTAIL.n168 1.93989
R943 VTAIL.n580 VTAIL.n500 1.93989
R944 VTAIL.n568 VTAIL.n506 1.93989
R945 VTAIL.n533 VTAIL.n523 1.93989
R946 VTAIL.n496 VTAIL.n416 1.93989
R947 VTAIL.n484 VTAIL.n422 1.93989
R948 VTAIL.n449 VTAIL.n439 1.93989
R949 VTAIL.n414 VTAIL.n334 1.93989
R950 VTAIL.n402 VTAIL.n340 1.93989
R951 VTAIL.n367 VTAIL.n357 1.93989
R952 VTAIL.n330 VTAIL.n250 1.93989
R953 VTAIL.n318 VTAIL.n256 1.93989
R954 VTAIL.n283 VTAIL.n273 1.93989
R955 VTAIL.n0 VTAIL.t3 1.3447
R956 VTAIL.n0 VTAIL.t4 1.3447
R957 VTAIL.n166 VTAIL.t14 1.3447
R958 VTAIL.n166 VTAIL.t13 1.3447
R959 VTAIL.n498 VTAIL.t12 1.3447
R960 VTAIL.n498 VTAIL.t10 1.3447
R961 VTAIL.n332 VTAIL.t6 1.3447
R962 VTAIL.n332 VTAIL.t0 1.3447
R963 VTAIL.n613 VTAIL.n606 1.16414
R964 VTAIL.n651 VTAIL.n586 1.16414
R965 VTAIL.n660 VTAIL.n659 1.16414
R966 VTAIL.n33 VTAIL.n26 1.16414
R967 VTAIL.n71 VTAIL.n6 1.16414
R968 VTAIL.n80 VTAIL.n79 1.16414
R969 VTAIL.n115 VTAIL.n108 1.16414
R970 VTAIL.n153 VTAIL.n88 1.16414
R971 VTAIL.n162 VTAIL.n161 1.16414
R972 VTAIL.n199 VTAIL.n192 1.16414
R973 VTAIL.n237 VTAIL.n172 1.16414
R974 VTAIL.n246 VTAIL.n245 1.16414
R975 VTAIL.n578 VTAIL.n577 1.16414
R976 VTAIL.n569 VTAIL.n504 1.16414
R977 VTAIL.n532 VTAIL.n525 1.16414
R978 VTAIL.n494 VTAIL.n493 1.16414
R979 VTAIL.n485 VTAIL.n420 1.16414
R980 VTAIL.n448 VTAIL.n441 1.16414
R981 VTAIL.n412 VTAIL.n411 1.16414
R982 VTAIL.n403 VTAIL.n338 1.16414
R983 VTAIL.n366 VTAIL.n359 1.16414
R984 VTAIL.n328 VTAIL.n327 1.16414
R985 VTAIL.n319 VTAIL.n254 1.16414
R986 VTAIL.n282 VTAIL.n275 1.16414
R987 VTAIL.n497 VTAIL.n415 0.470328
R988 VTAIL.n165 VTAIL.n83 0.470328
R989 VTAIL.n610 VTAIL.n609 0.388379
R990 VTAIL.n655 VTAIL.n654 0.388379
R991 VTAIL.n656 VTAIL.n584 0.388379
R992 VTAIL.n30 VTAIL.n29 0.388379
R993 VTAIL.n75 VTAIL.n74 0.388379
R994 VTAIL.n76 VTAIL.n4 0.388379
R995 VTAIL.n112 VTAIL.n111 0.388379
R996 VTAIL.n157 VTAIL.n156 0.388379
R997 VTAIL.n158 VTAIL.n86 0.388379
R998 VTAIL.n196 VTAIL.n195 0.388379
R999 VTAIL.n241 VTAIL.n240 0.388379
R1000 VTAIL.n242 VTAIL.n170 0.388379
R1001 VTAIL.n574 VTAIL.n502 0.388379
R1002 VTAIL.n573 VTAIL.n572 0.388379
R1003 VTAIL.n529 VTAIL.n528 0.388379
R1004 VTAIL.n490 VTAIL.n418 0.388379
R1005 VTAIL.n489 VTAIL.n488 0.388379
R1006 VTAIL.n445 VTAIL.n444 0.388379
R1007 VTAIL.n408 VTAIL.n336 0.388379
R1008 VTAIL.n407 VTAIL.n406 0.388379
R1009 VTAIL.n363 VTAIL.n362 0.388379
R1010 VTAIL.n324 VTAIL.n252 0.388379
R1011 VTAIL.n323 VTAIL.n322 0.388379
R1012 VTAIL.n279 VTAIL.n278 0.388379
R1013 VTAIL.n612 VTAIL.n611 0.155672
R1014 VTAIL.n612 VTAIL.n603 0.155672
R1015 VTAIL.n619 VTAIL.n603 0.155672
R1016 VTAIL.n620 VTAIL.n619 0.155672
R1017 VTAIL.n620 VTAIL.n599 0.155672
R1018 VTAIL.n627 VTAIL.n599 0.155672
R1019 VTAIL.n628 VTAIL.n627 0.155672
R1020 VTAIL.n628 VTAIL.n595 0.155672
R1021 VTAIL.n635 VTAIL.n595 0.155672
R1022 VTAIL.n636 VTAIL.n635 0.155672
R1023 VTAIL.n636 VTAIL.n591 0.155672
R1024 VTAIL.n643 VTAIL.n591 0.155672
R1025 VTAIL.n644 VTAIL.n643 0.155672
R1026 VTAIL.n644 VTAIL.n587 0.155672
R1027 VTAIL.n652 VTAIL.n587 0.155672
R1028 VTAIL.n653 VTAIL.n652 0.155672
R1029 VTAIL.n653 VTAIL.n583 0.155672
R1030 VTAIL.n661 VTAIL.n583 0.155672
R1031 VTAIL.n32 VTAIL.n31 0.155672
R1032 VTAIL.n32 VTAIL.n23 0.155672
R1033 VTAIL.n39 VTAIL.n23 0.155672
R1034 VTAIL.n40 VTAIL.n39 0.155672
R1035 VTAIL.n40 VTAIL.n19 0.155672
R1036 VTAIL.n47 VTAIL.n19 0.155672
R1037 VTAIL.n48 VTAIL.n47 0.155672
R1038 VTAIL.n48 VTAIL.n15 0.155672
R1039 VTAIL.n55 VTAIL.n15 0.155672
R1040 VTAIL.n56 VTAIL.n55 0.155672
R1041 VTAIL.n56 VTAIL.n11 0.155672
R1042 VTAIL.n63 VTAIL.n11 0.155672
R1043 VTAIL.n64 VTAIL.n63 0.155672
R1044 VTAIL.n64 VTAIL.n7 0.155672
R1045 VTAIL.n72 VTAIL.n7 0.155672
R1046 VTAIL.n73 VTAIL.n72 0.155672
R1047 VTAIL.n73 VTAIL.n3 0.155672
R1048 VTAIL.n81 VTAIL.n3 0.155672
R1049 VTAIL.n114 VTAIL.n113 0.155672
R1050 VTAIL.n114 VTAIL.n105 0.155672
R1051 VTAIL.n121 VTAIL.n105 0.155672
R1052 VTAIL.n122 VTAIL.n121 0.155672
R1053 VTAIL.n122 VTAIL.n101 0.155672
R1054 VTAIL.n129 VTAIL.n101 0.155672
R1055 VTAIL.n130 VTAIL.n129 0.155672
R1056 VTAIL.n130 VTAIL.n97 0.155672
R1057 VTAIL.n137 VTAIL.n97 0.155672
R1058 VTAIL.n138 VTAIL.n137 0.155672
R1059 VTAIL.n138 VTAIL.n93 0.155672
R1060 VTAIL.n145 VTAIL.n93 0.155672
R1061 VTAIL.n146 VTAIL.n145 0.155672
R1062 VTAIL.n146 VTAIL.n89 0.155672
R1063 VTAIL.n154 VTAIL.n89 0.155672
R1064 VTAIL.n155 VTAIL.n154 0.155672
R1065 VTAIL.n155 VTAIL.n85 0.155672
R1066 VTAIL.n163 VTAIL.n85 0.155672
R1067 VTAIL.n198 VTAIL.n197 0.155672
R1068 VTAIL.n198 VTAIL.n189 0.155672
R1069 VTAIL.n205 VTAIL.n189 0.155672
R1070 VTAIL.n206 VTAIL.n205 0.155672
R1071 VTAIL.n206 VTAIL.n185 0.155672
R1072 VTAIL.n213 VTAIL.n185 0.155672
R1073 VTAIL.n214 VTAIL.n213 0.155672
R1074 VTAIL.n214 VTAIL.n181 0.155672
R1075 VTAIL.n221 VTAIL.n181 0.155672
R1076 VTAIL.n222 VTAIL.n221 0.155672
R1077 VTAIL.n222 VTAIL.n177 0.155672
R1078 VTAIL.n229 VTAIL.n177 0.155672
R1079 VTAIL.n230 VTAIL.n229 0.155672
R1080 VTAIL.n230 VTAIL.n173 0.155672
R1081 VTAIL.n238 VTAIL.n173 0.155672
R1082 VTAIL.n239 VTAIL.n238 0.155672
R1083 VTAIL.n239 VTAIL.n169 0.155672
R1084 VTAIL.n247 VTAIL.n169 0.155672
R1085 VTAIL.n579 VTAIL.n501 0.155672
R1086 VTAIL.n571 VTAIL.n501 0.155672
R1087 VTAIL.n571 VTAIL.n570 0.155672
R1088 VTAIL.n570 VTAIL.n505 0.155672
R1089 VTAIL.n563 VTAIL.n505 0.155672
R1090 VTAIL.n563 VTAIL.n562 0.155672
R1091 VTAIL.n562 VTAIL.n510 0.155672
R1092 VTAIL.n555 VTAIL.n510 0.155672
R1093 VTAIL.n555 VTAIL.n554 0.155672
R1094 VTAIL.n554 VTAIL.n514 0.155672
R1095 VTAIL.n547 VTAIL.n514 0.155672
R1096 VTAIL.n547 VTAIL.n546 0.155672
R1097 VTAIL.n546 VTAIL.n518 0.155672
R1098 VTAIL.n539 VTAIL.n518 0.155672
R1099 VTAIL.n539 VTAIL.n538 0.155672
R1100 VTAIL.n538 VTAIL.n522 0.155672
R1101 VTAIL.n531 VTAIL.n522 0.155672
R1102 VTAIL.n531 VTAIL.n530 0.155672
R1103 VTAIL.n495 VTAIL.n417 0.155672
R1104 VTAIL.n487 VTAIL.n417 0.155672
R1105 VTAIL.n487 VTAIL.n486 0.155672
R1106 VTAIL.n486 VTAIL.n421 0.155672
R1107 VTAIL.n479 VTAIL.n421 0.155672
R1108 VTAIL.n479 VTAIL.n478 0.155672
R1109 VTAIL.n478 VTAIL.n426 0.155672
R1110 VTAIL.n471 VTAIL.n426 0.155672
R1111 VTAIL.n471 VTAIL.n470 0.155672
R1112 VTAIL.n470 VTAIL.n430 0.155672
R1113 VTAIL.n463 VTAIL.n430 0.155672
R1114 VTAIL.n463 VTAIL.n462 0.155672
R1115 VTAIL.n462 VTAIL.n434 0.155672
R1116 VTAIL.n455 VTAIL.n434 0.155672
R1117 VTAIL.n455 VTAIL.n454 0.155672
R1118 VTAIL.n454 VTAIL.n438 0.155672
R1119 VTAIL.n447 VTAIL.n438 0.155672
R1120 VTAIL.n447 VTAIL.n446 0.155672
R1121 VTAIL.n413 VTAIL.n335 0.155672
R1122 VTAIL.n405 VTAIL.n335 0.155672
R1123 VTAIL.n405 VTAIL.n404 0.155672
R1124 VTAIL.n404 VTAIL.n339 0.155672
R1125 VTAIL.n397 VTAIL.n339 0.155672
R1126 VTAIL.n397 VTAIL.n396 0.155672
R1127 VTAIL.n396 VTAIL.n344 0.155672
R1128 VTAIL.n389 VTAIL.n344 0.155672
R1129 VTAIL.n389 VTAIL.n388 0.155672
R1130 VTAIL.n388 VTAIL.n348 0.155672
R1131 VTAIL.n381 VTAIL.n348 0.155672
R1132 VTAIL.n381 VTAIL.n380 0.155672
R1133 VTAIL.n380 VTAIL.n352 0.155672
R1134 VTAIL.n373 VTAIL.n352 0.155672
R1135 VTAIL.n373 VTAIL.n372 0.155672
R1136 VTAIL.n372 VTAIL.n356 0.155672
R1137 VTAIL.n365 VTAIL.n356 0.155672
R1138 VTAIL.n365 VTAIL.n364 0.155672
R1139 VTAIL.n329 VTAIL.n251 0.155672
R1140 VTAIL.n321 VTAIL.n251 0.155672
R1141 VTAIL.n321 VTAIL.n320 0.155672
R1142 VTAIL.n320 VTAIL.n255 0.155672
R1143 VTAIL.n313 VTAIL.n255 0.155672
R1144 VTAIL.n313 VTAIL.n312 0.155672
R1145 VTAIL.n312 VTAIL.n260 0.155672
R1146 VTAIL.n305 VTAIL.n260 0.155672
R1147 VTAIL.n305 VTAIL.n304 0.155672
R1148 VTAIL.n304 VTAIL.n264 0.155672
R1149 VTAIL.n297 VTAIL.n264 0.155672
R1150 VTAIL.n297 VTAIL.n296 0.155672
R1151 VTAIL.n296 VTAIL.n268 0.155672
R1152 VTAIL.n289 VTAIL.n268 0.155672
R1153 VTAIL.n289 VTAIL.n288 0.155672
R1154 VTAIL.n288 VTAIL.n272 0.155672
R1155 VTAIL.n281 VTAIL.n272 0.155672
R1156 VTAIL.n281 VTAIL.n280 0.155672
R1157 VTAIL VTAIL.n1 0.0586897
R1158 B.n1092 B.n1091 585
R1159 B.n1093 B.n1092 585
R1160 B.n395 B.n177 585
R1161 B.n394 B.n393 585
R1162 B.n392 B.n391 585
R1163 B.n390 B.n389 585
R1164 B.n388 B.n387 585
R1165 B.n386 B.n385 585
R1166 B.n384 B.n383 585
R1167 B.n382 B.n381 585
R1168 B.n380 B.n379 585
R1169 B.n378 B.n377 585
R1170 B.n376 B.n375 585
R1171 B.n374 B.n373 585
R1172 B.n372 B.n371 585
R1173 B.n370 B.n369 585
R1174 B.n368 B.n367 585
R1175 B.n366 B.n365 585
R1176 B.n364 B.n363 585
R1177 B.n362 B.n361 585
R1178 B.n360 B.n359 585
R1179 B.n358 B.n357 585
R1180 B.n356 B.n355 585
R1181 B.n354 B.n353 585
R1182 B.n352 B.n351 585
R1183 B.n350 B.n349 585
R1184 B.n348 B.n347 585
R1185 B.n346 B.n345 585
R1186 B.n344 B.n343 585
R1187 B.n342 B.n341 585
R1188 B.n340 B.n339 585
R1189 B.n338 B.n337 585
R1190 B.n336 B.n335 585
R1191 B.n334 B.n333 585
R1192 B.n332 B.n331 585
R1193 B.n330 B.n329 585
R1194 B.n328 B.n327 585
R1195 B.n326 B.n325 585
R1196 B.n324 B.n323 585
R1197 B.n322 B.n321 585
R1198 B.n320 B.n319 585
R1199 B.n318 B.n317 585
R1200 B.n316 B.n315 585
R1201 B.n314 B.n313 585
R1202 B.n312 B.n311 585
R1203 B.n310 B.n309 585
R1204 B.n308 B.n307 585
R1205 B.n306 B.n305 585
R1206 B.n304 B.n303 585
R1207 B.n302 B.n301 585
R1208 B.n300 B.n299 585
R1209 B.n297 B.n296 585
R1210 B.n295 B.n294 585
R1211 B.n293 B.n292 585
R1212 B.n291 B.n290 585
R1213 B.n289 B.n288 585
R1214 B.n287 B.n286 585
R1215 B.n285 B.n284 585
R1216 B.n283 B.n282 585
R1217 B.n281 B.n280 585
R1218 B.n279 B.n278 585
R1219 B.n277 B.n276 585
R1220 B.n275 B.n274 585
R1221 B.n273 B.n272 585
R1222 B.n271 B.n270 585
R1223 B.n269 B.n268 585
R1224 B.n267 B.n266 585
R1225 B.n265 B.n264 585
R1226 B.n263 B.n262 585
R1227 B.n261 B.n260 585
R1228 B.n259 B.n258 585
R1229 B.n257 B.n256 585
R1230 B.n255 B.n254 585
R1231 B.n253 B.n252 585
R1232 B.n251 B.n250 585
R1233 B.n249 B.n248 585
R1234 B.n247 B.n246 585
R1235 B.n245 B.n244 585
R1236 B.n243 B.n242 585
R1237 B.n241 B.n240 585
R1238 B.n239 B.n238 585
R1239 B.n237 B.n236 585
R1240 B.n235 B.n234 585
R1241 B.n233 B.n232 585
R1242 B.n231 B.n230 585
R1243 B.n229 B.n228 585
R1244 B.n227 B.n226 585
R1245 B.n225 B.n224 585
R1246 B.n223 B.n222 585
R1247 B.n221 B.n220 585
R1248 B.n219 B.n218 585
R1249 B.n217 B.n216 585
R1250 B.n215 B.n214 585
R1251 B.n213 B.n212 585
R1252 B.n211 B.n210 585
R1253 B.n209 B.n208 585
R1254 B.n207 B.n206 585
R1255 B.n205 B.n204 585
R1256 B.n203 B.n202 585
R1257 B.n201 B.n200 585
R1258 B.n199 B.n198 585
R1259 B.n197 B.n196 585
R1260 B.n195 B.n194 585
R1261 B.n193 B.n192 585
R1262 B.n191 B.n190 585
R1263 B.n189 B.n188 585
R1264 B.n187 B.n186 585
R1265 B.n185 B.n184 585
R1266 B.n123 B.n122 585
R1267 B.n1096 B.n1095 585
R1268 B.n1090 B.n178 585
R1269 B.n178 B.n120 585
R1270 B.n1089 B.n119 585
R1271 B.n1100 B.n119 585
R1272 B.n1088 B.n118 585
R1273 B.n1101 B.n118 585
R1274 B.n1087 B.n117 585
R1275 B.n1102 B.n117 585
R1276 B.n1086 B.n1085 585
R1277 B.n1085 B.n113 585
R1278 B.n1084 B.n112 585
R1279 B.n1108 B.n112 585
R1280 B.n1083 B.n111 585
R1281 B.n1109 B.n111 585
R1282 B.n1082 B.n110 585
R1283 B.n1110 B.n110 585
R1284 B.n1081 B.n1080 585
R1285 B.n1080 B.n106 585
R1286 B.n1079 B.n105 585
R1287 B.n1116 B.n105 585
R1288 B.n1078 B.n104 585
R1289 B.n1117 B.n104 585
R1290 B.n1077 B.n103 585
R1291 B.n1118 B.n103 585
R1292 B.n1076 B.n1075 585
R1293 B.n1075 B.n99 585
R1294 B.n1074 B.n98 585
R1295 B.n1124 B.n98 585
R1296 B.n1073 B.n97 585
R1297 B.n1125 B.n97 585
R1298 B.n1072 B.n96 585
R1299 B.n1126 B.n96 585
R1300 B.n1071 B.n1070 585
R1301 B.n1070 B.n92 585
R1302 B.n1069 B.n91 585
R1303 B.n1132 B.n91 585
R1304 B.n1068 B.n90 585
R1305 B.n1133 B.n90 585
R1306 B.n1067 B.n89 585
R1307 B.n1134 B.n89 585
R1308 B.n1066 B.n1065 585
R1309 B.n1065 B.n85 585
R1310 B.n1064 B.n84 585
R1311 B.n1140 B.n84 585
R1312 B.n1063 B.n83 585
R1313 B.n1141 B.n83 585
R1314 B.n1062 B.n82 585
R1315 B.n1142 B.n82 585
R1316 B.n1061 B.n1060 585
R1317 B.n1060 B.n81 585
R1318 B.n1059 B.n77 585
R1319 B.n1148 B.n77 585
R1320 B.n1058 B.n76 585
R1321 B.n1149 B.n76 585
R1322 B.n1057 B.n75 585
R1323 B.n1150 B.n75 585
R1324 B.n1056 B.n1055 585
R1325 B.n1055 B.n71 585
R1326 B.n1054 B.n70 585
R1327 B.n1156 B.n70 585
R1328 B.n1053 B.n69 585
R1329 B.n1157 B.n69 585
R1330 B.n1052 B.n68 585
R1331 B.n1158 B.n68 585
R1332 B.n1051 B.n1050 585
R1333 B.n1050 B.n64 585
R1334 B.n1049 B.n63 585
R1335 B.n1164 B.n63 585
R1336 B.n1048 B.n62 585
R1337 B.n1165 B.n62 585
R1338 B.n1047 B.n61 585
R1339 B.n1166 B.n61 585
R1340 B.n1046 B.n1045 585
R1341 B.n1045 B.n60 585
R1342 B.n1044 B.n56 585
R1343 B.n1172 B.n56 585
R1344 B.n1043 B.n55 585
R1345 B.n1173 B.n55 585
R1346 B.n1042 B.n54 585
R1347 B.n1174 B.n54 585
R1348 B.n1041 B.n1040 585
R1349 B.n1040 B.n50 585
R1350 B.n1039 B.n49 585
R1351 B.n1180 B.n49 585
R1352 B.n1038 B.n48 585
R1353 B.n1181 B.n48 585
R1354 B.n1037 B.n47 585
R1355 B.n1182 B.n47 585
R1356 B.n1036 B.n1035 585
R1357 B.n1035 B.n43 585
R1358 B.n1034 B.n42 585
R1359 B.n1188 B.n42 585
R1360 B.n1033 B.n41 585
R1361 B.n1189 B.n41 585
R1362 B.n1032 B.n40 585
R1363 B.n1190 B.n40 585
R1364 B.n1031 B.n1030 585
R1365 B.n1030 B.n36 585
R1366 B.n1029 B.n35 585
R1367 B.n1196 B.n35 585
R1368 B.n1028 B.n34 585
R1369 B.n1197 B.n34 585
R1370 B.n1027 B.n33 585
R1371 B.n1198 B.n33 585
R1372 B.n1026 B.n1025 585
R1373 B.n1025 B.n29 585
R1374 B.n1024 B.n28 585
R1375 B.n1204 B.n28 585
R1376 B.n1023 B.n27 585
R1377 B.n1205 B.n27 585
R1378 B.n1022 B.n26 585
R1379 B.n1206 B.n26 585
R1380 B.n1021 B.n1020 585
R1381 B.n1020 B.n22 585
R1382 B.n1019 B.n21 585
R1383 B.n1212 B.n21 585
R1384 B.n1018 B.n20 585
R1385 B.n1213 B.n20 585
R1386 B.n1017 B.n19 585
R1387 B.n1214 B.n19 585
R1388 B.n1016 B.n1015 585
R1389 B.n1015 B.n15 585
R1390 B.n1014 B.n14 585
R1391 B.n1220 B.n14 585
R1392 B.n1013 B.n13 585
R1393 B.n1221 B.n13 585
R1394 B.n1012 B.n12 585
R1395 B.n1222 B.n12 585
R1396 B.n1011 B.n1010 585
R1397 B.n1010 B.n8 585
R1398 B.n1009 B.n7 585
R1399 B.n1228 B.n7 585
R1400 B.n1008 B.n6 585
R1401 B.n1229 B.n6 585
R1402 B.n1007 B.n5 585
R1403 B.n1230 B.n5 585
R1404 B.n1006 B.n1005 585
R1405 B.n1005 B.n4 585
R1406 B.n1004 B.n396 585
R1407 B.n1004 B.n1003 585
R1408 B.n994 B.n397 585
R1409 B.n398 B.n397 585
R1410 B.n996 B.n995 585
R1411 B.n997 B.n996 585
R1412 B.n993 B.n403 585
R1413 B.n403 B.n402 585
R1414 B.n992 B.n991 585
R1415 B.n991 B.n990 585
R1416 B.n405 B.n404 585
R1417 B.n406 B.n405 585
R1418 B.n983 B.n982 585
R1419 B.n984 B.n983 585
R1420 B.n981 B.n411 585
R1421 B.n411 B.n410 585
R1422 B.n980 B.n979 585
R1423 B.n979 B.n978 585
R1424 B.n413 B.n412 585
R1425 B.n414 B.n413 585
R1426 B.n971 B.n970 585
R1427 B.n972 B.n971 585
R1428 B.n969 B.n419 585
R1429 B.n419 B.n418 585
R1430 B.n968 B.n967 585
R1431 B.n967 B.n966 585
R1432 B.n421 B.n420 585
R1433 B.n422 B.n421 585
R1434 B.n959 B.n958 585
R1435 B.n960 B.n959 585
R1436 B.n957 B.n427 585
R1437 B.n427 B.n426 585
R1438 B.n956 B.n955 585
R1439 B.n955 B.n954 585
R1440 B.n429 B.n428 585
R1441 B.n430 B.n429 585
R1442 B.n947 B.n946 585
R1443 B.n948 B.n947 585
R1444 B.n945 B.n435 585
R1445 B.n435 B.n434 585
R1446 B.n944 B.n943 585
R1447 B.n943 B.n942 585
R1448 B.n437 B.n436 585
R1449 B.n438 B.n437 585
R1450 B.n935 B.n934 585
R1451 B.n936 B.n935 585
R1452 B.n933 B.n443 585
R1453 B.n443 B.n442 585
R1454 B.n932 B.n931 585
R1455 B.n931 B.n930 585
R1456 B.n445 B.n444 585
R1457 B.n446 B.n445 585
R1458 B.n923 B.n922 585
R1459 B.n924 B.n923 585
R1460 B.n921 B.n451 585
R1461 B.n451 B.n450 585
R1462 B.n920 B.n919 585
R1463 B.n919 B.n918 585
R1464 B.n453 B.n452 585
R1465 B.n911 B.n453 585
R1466 B.n910 B.n909 585
R1467 B.n912 B.n910 585
R1468 B.n908 B.n458 585
R1469 B.n458 B.n457 585
R1470 B.n907 B.n906 585
R1471 B.n906 B.n905 585
R1472 B.n460 B.n459 585
R1473 B.n461 B.n460 585
R1474 B.n898 B.n897 585
R1475 B.n899 B.n898 585
R1476 B.n896 B.n466 585
R1477 B.n466 B.n465 585
R1478 B.n895 B.n894 585
R1479 B.n894 B.n893 585
R1480 B.n468 B.n467 585
R1481 B.n469 B.n468 585
R1482 B.n886 B.n885 585
R1483 B.n887 B.n886 585
R1484 B.n884 B.n474 585
R1485 B.n474 B.n473 585
R1486 B.n883 B.n882 585
R1487 B.n882 B.n881 585
R1488 B.n476 B.n475 585
R1489 B.n874 B.n476 585
R1490 B.n873 B.n872 585
R1491 B.n875 B.n873 585
R1492 B.n871 B.n481 585
R1493 B.n481 B.n480 585
R1494 B.n870 B.n869 585
R1495 B.n869 B.n868 585
R1496 B.n483 B.n482 585
R1497 B.n484 B.n483 585
R1498 B.n861 B.n860 585
R1499 B.n862 B.n861 585
R1500 B.n859 B.n489 585
R1501 B.n489 B.n488 585
R1502 B.n858 B.n857 585
R1503 B.n857 B.n856 585
R1504 B.n491 B.n490 585
R1505 B.n492 B.n491 585
R1506 B.n849 B.n848 585
R1507 B.n850 B.n849 585
R1508 B.n847 B.n497 585
R1509 B.n497 B.n496 585
R1510 B.n846 B.n845 585
R1511 B.n845 B.n844 585
R1512 B.n499 B.n498 585
R1513 B.n500 B.n499 585
R1514 B.n837 B.n836 585
R1515 B.n838 B.n837 585
R1516 B.n835 B.n505 585
R1517 B.n505 B.n504 585
R1518 B.n834 B.n833 585
R1519 B.n833 B.n832 585
R1520 B.n507 B.n506 585
R1521 B.n508 B.n507 585
R1522 B.n825 B.n824 585
R1523 B.n826 B.n825 585
R1524 B.n823 B.n513 585
R1525 B.n513 B.n512 585
R1526 B.n822 B.n821 585
R1527 B.n821 B.n820 585
R1528 B.n515 B.n514 585
R1529 B.n516 B.n515 585
R1530 B.n813 B.n812 585
R1531 B.n814 B.n813 585
R1532 B.n811 B.n521 585
R1533 B.n521 B.n520 585
R1534 B.n810 B.n809 585
R1535 B.n809 B.n808 585
R1536 B.n523 B.n522 585
R1537 B.n524 B.n523 585
R1538 B.n804 B.n803 585
R1539 B.n527 B.n526 585
R1540 B.n800 B.n799 585
R1541 B.n801 B.n800 585
R1542 B.n798 B.n581 585
R1543 B.n797 B.n796 585
R1544 B.n795 B.n794 585
R1545 B.n793 B.n792 585
R1546 B.n791 B.n790 585
R1547 B.n789 B.n788 585
R1548 B.n787 B.n786 585
R1549 B.n785 B.n784 585
R1550 B.n783 B.n782 585
R1551 B.n781 B.n780 585
R1552 B.n779 B.n778 585
R1553 B.n777 B.n776 585
R1554 B.n775 B.n774 585
R1555 B.n773 B.n772 585
R1556 B.n771 B.n770 585
R1557 B.n769 B.n768 585
R1558 B.n767 B.n766 585
R1559 B.n765 B.n764 585
R1560 B.n763 B.n762 585
R1561 B.n761 B.n760 585
R1562 B.n759 B.n758 585
R1563 B.n757 B.n756 585
R1564 B.n755 B.n754 585
R1565 B.n753 B.n752 585
R1566 B.n751 B.n750 585
R1567 B.n749 B.n748 585
R1568 B.n747 B.n746 585
R1569 B.n745 B.n744 585
R1570 B.n743 B.n742 585
R1571 B.n741 B.n740 585
R1572 B.n739 B.n738 585
R1573 B.n737 B.n736 585
R1574 B.n735 B.n734 585
R1575 B.n733 B.n732 585
R1576 B.n731 B.n730 585
R1577 B.n729 B.n728 585
R1578 B.n727 B.n726 585
R1579 B.n725 B.n724 585
R1580 B.n723 B.n722 585
R1581 B.n721 B.n720 585
R1582 B.n719 B.n718 585
R1583 B.n717 B.n716 585
R1584 B.n715 B.n714 585
R1585 B.n713 B.n712 585
R1586 B.n711 B.n710 585
R1587 B.n709 B.n708 585
R1588 B.n707 B.n706 585
R1589 B.n704 B.n703 585
R1590 B.n702 B.n701 585
R1591 B.n700 B.n699 585
R1592 B.n698 B.n697 585
R1593 B.n696 B.n695 585
R1594 B.n694 B.n693 585
R1595 B.n692 B.n691 585
R1596 B.n690 B.n689 585
R1597 B.n688 B.n687 585
R1598 B.n686 B.n685 585
R1599 B.n684 B.n683 585
R1600 B.n682 B.n681 585
R1601 B.n680 B.n679 585
R1602 B.n678 B.n677 585
R1603 B.n676 B.n675 585
R1604 B.n674 B.n673 585
R1605 B.n672 B.n671 585
R1606 B.n670 B.n669 585
R1607 B.n668 B.n667 585
R1608 B.n666 B.n665 585
R1609 B.n664 B.n663 585
R1610 B.n662 B.n661 585
R1611 B.n660 B.n659 585
R1612 B.n658 B.n657 585
R1613 B.n656 B.n655 585
R1614 B.n654 B.n653 585
R1615 B.n652 B.n651 585
R1616 B.n650 B.n649 585
R1617 B.n648 B.n647 585
R1618 B.n646 B.n645 585
R1619 B.n644 B.n643 585
R1620 B.n642 B.n641 585
R1621 B.n640 B.n639 585
R1622 B.n638 B.n637 585
R1623 B.n636 B.n635 585
R1624 B.n634 B.n633 585
R1625 B.n632 B.n631 585
R1626 B.n630 B.n629 585
R1627 B.n628 B.n627 585
R1628 B.n626 B.n625 585
R1629 B.n624 B.n623 585
R1630 B.n622 B.n621 585
R1631 B.n620 B.n619 585
R1632 B.n618 B.n617 585
R1633 B.n616 B.n615 585
R1634 B.n614 B.n613 585
R1635 B.n612 B.n611 585
R1636 B.n610 B.n609 585
R1637 B.n608 B.n607 585
R1638 B.n606 B.n605 585
R1639 B.n604 B.n603 585
R1640 B.n602 B.n601 585
R1641 B.n600 B.n599 585
R1642 B.n598 B.n597 585
R1643 B.n596 B.n595 585
R1644 B.n594 B.n593 585
R1645 B.n592 B.n591 585
R1646 B.n590 B.n589 585
R1647 B.n588 B.n587 585
R1648 B.n805 B.n525 585
R1649 B.n525 B.n524 585
R1650 B.n807 B.n806 585
R1651 B.n808 B.n807 585
R1652 B.n519 B.n518 585
R1653 B.n520 B.n519 585
R1654 B.n816 B.n815 585
R1655 B.n815 B.n814 585
R1656 B.n817 B.n517 585
R1657 B.n517 B.n516 585
R1658 B.n819 B.n818 585
R1659 B.n820 B.n819 585
R1660 B.n511 B.n510 585
R1661 B.n512 B.n511 585
R1662 B.n828 B.n827 585
R1663 B.n827 B.n826 585
R1664 B.n829 B.n509 585
R1665 B.n509 B.n508 585
R1666 B.n831 B.n830 585
R1667 B.n832 B.n831 585
R1668 B.n503 B.n502 585
R1669 B.n504 B.n503 585
R1670 B.n840 B.n839 585
R1671 B.n839 B.n838 585
R1672 B.n841 B.n501 585
R1673 B.n501 B.n500 585
R1674 B.n843 B.n842 585
R1675 B.n844 B.n843 585
R1676 B.n495 B.n494 585
R1677 B.n496 B.n495 585
R1678 B.n852 B.n851 585
R1679 B.n851 B.n850 585
R1680 B.n853 B.n493 585
R1681 B.n493 B.n492 585
R1682 B.n855 B.n854 585
R1683 B.n856 B.n855 585
R1684 B.n487 B.n486 585
R1685 B.n488 B.n487 585
R1686 B.n864 B.n863 585
R1687 B.n863 B.n862 585
R1688 B.n865 B.n485 585
R1689 B.n485 B.n484 585
R1690 B.n867 B.n866 585
R1691 B.n868 B.n867 585
R1692 B.n479 B.n478 585
R1693 B.n480 B.n479 585
R1694 B.n877 B.n876 585
R1695 B.n876 B.n875 585
R1696 B.n878 B.n477 585
R1697 B.n874 B.n477 585
R1698 B.n880 B.n879 585
R1699 B.n881 B.n880 585
R1700 B.n472 B.n471 585
R1701 B.n473 B.n472 585
R1702 B.n889 B.n888 585
R1703 B.n888 B.n887 585
R1704 B.n890 B.n470 585
R1705 B.n470 B.n469 585
R1706 B.n892 B.n891 585
R1707 B.n893 B.n892 585
R1708 B.n464 B.n463 585
R1709 B.n465 B.n464 585
R1710 B.n901 B.n900 585
R1711 B.n900 B.n899 585
R1712 B.n902 B.n462 585
R1713 B.n462 B.n461 585
R1714 B.n904 B.n903 585
R1715 B.n905 B.n904 585
R1716 B.n456 B.n455 585
R1717 B.n457 B.n456 585
R1718 B.n914 B.n913 585
R1719 B.n913 B.n912 585
R1720 B.n915 B.n454 585
R1721 B.n911 B.n454 585
R1722 B.n917 B.n916 585
R1723 B.n918 B.n917 585
R1724 B.n449 B.n448 585
R1725 B.n450 B.n449 585
R1726 B.n926 B.n925 585
R1727 B.n925 B.n924 585
R1728 B.n927 B.n447 585
R1729 B.n447 B.n446 585
R1730 B.n929 B.n928 585
R1731 B.n930 B.n929 585
R1732 B.n441 B.n440 585
R1733 B.n442 B.n441 585
R1734 B.n938 B.n937 585
R1735 B.n937 B.n936 585
R1736 B.n939 B.n439 585
R1737 B.n439 B.n438 585
R1738 B.n941 B.n940 585
R1739 B.n942 B.n941 585
R1740 B.n433 B.n432 585
R1741 B.n434 B.n433 585
R1742 B.n950 B.n949 585
R1743 B.n949 B.n948 585
R1744 B.n951 B.n431 585
R1745 B.n431 B.n430 585
R1746 B.n953 B.n952 585
R1747 B.n954 B.n953 585
R1748 B.n425 B.n424 585
R1749 B.n426 B.n425 585
R1750 B.n962 B.n961 585
R1751 B.n961 B.n960 585
R1752 B.n963 B.n423 585
R1753 B.n423 B.n422 585
R1754 B.n965 B.n964 585
R1755 B.n966 B.n965 585
R1756 B.n417 B.n416 585
R1757 B.n418 B.n417 585
R1758 B.n974 B.n973 585
R1759 B.n973 B.n972 585
R1760 B.n975 B.n415 585
R1761 B.n415 B.n414 585
R1762 B.n977 B.n976 585
R1763 B.n978 B.n977 585
R1764 B.n409 B.n408 585
R1765 B.n410 B.n409 585
R1766 B.n986 B.n985 585
R1767 B.n985 B.n984 585
R1768 B.n987 B.n407 585
R1769 B.n407 B.n406 585
R1770 B.n989 B.n988 585
R1771 B.n990 B.n989 585
R1772 B.n401 B.n400 585
R1773 B.n402 B.n401 585
R1774 B.n999 B.n998 585
R1775 B.n998 B.n997 585
R1776 B.n1000 B.n399 585
R1777 B.n399 B.n398 585
R1778 B.n1002 B.n1001 585
R1779 B.n1003 B.n1002 585
R1780 B.n2 B.n0 585
R1781 B.n4 B.n2 585
R1782 B.n3 B.n1 585
R1783 B.n1229 B.n3 585
R1784 B.n1227 B.n1226 585
R1785 B.n1228 B.n1227 585
R1786 B.n1225 B.n9 585
R1787 B.n9 B.n8 585
R1788 B.n1224 B.n1223 585
R1789 B.n1223 B.n1222 585
R1790 B.n11 B.n10 585
R1791 B.n1221 B.n11 585
R1792 B.n1219 B.n1218 585
R1793 B.n1220 B.n1219 585
R1794 B.n1217 B.n16 585
R1795 B.n16 B.n15 585
R1796 B.n1216 B.n1215 585
R1797 B.n1215 B.n1214 585
R1798 B.n18 B.n17 585
R1799 B.n1213 B.n18 585
R1800 B.n1211 B.n1210 585
R1801 B.n1212 B.n1211 585
R1802 B.n1209 B.n23 585
R1803 B.n23 B.n22 585
R1804 B.n1208 B.n1207 585
R1805 B.n1207 B.n1206 585
R1806 B.n25 B.n24 585
R1807 B.n1205 B.n25 585
R1808 B.n1203 B.n1202 585
R1809 B.n1204 B.n1203 585
R1810 B.n1201 B.n30 585
R1811 B.n30 B.n29 585
R1812 B.n1200 B.n1199 585
R1813 B.n1199 B.n1198 585
R1814 B.n32 B.n31 585
R1815 B.n1197 B.n32 585
R1816 B.n1195 B.n1194 585
R1817 B.n1196 B.n1195 585
R1818 B.n1193 B.n37 585
R1819 B.n37 B.n36 585
R1820 B.n1192 B.n1191 585
R1821 B.n1191 B.n1190 585
R1822 B.n39 B.n38 585
R1823 B.n1189 B.n39 585
R1824 B.n1187 B.n1186 585
R1825 B.n1188 B.n1187 585
R1826 B.n1185 B.n44 585
R1827 B.n44 B.n43 585
R1828 B.n1184 B.n1183 585
R1829 B.n1183 B.n1182 585
R1830 B.n46 B.n45 585
R1831 B.n1181 B.n46 585
R1832 B.n1179 B.n1178 585
R1833 B.n1180 B.n1179 585
R1834 B.n1177 B.n51 585
R1835 B.n51 B.n50 585
R1836 B.n1176 B.n1175 585
R1837 B.n1175 B.n1174 585
R1838 B.n53 B.n52 585
R1839 B.n1173 B.n53 585
R1840 B.n1171 B.n1170 585
R1841 B.n1172 B.n1171 585
R1842 B.n1169 B.n57 585
R1843 B.n60 B.n57 585
R1844 B.n1168 B.n1167 585
R1845 B.n1167 B.n1166 585
R1846 B.n59 B.n58 585
R1847 B.n1165 B.n59 585
R1848 B.n1163 B.n1162 585
R1849 B.n1164 B.n1163 585
R1850 B.n1161 B.n65 585
R1851 B.n65 B.n64 585
R1852 B.n1160 B.n1159 585
R1853 B.n1159 B.n1158 585
R1854 B.n67 B.n66 585
R1855 B.n1157 B.n67 585
R1856 B.n1155 B.n1154 585
R1857 B.n1156 B.n1155 585
R1858 B.n1153 B.n72 585
R1859 B.n72 B.n71 585
R1860 B.n1152 B.n1151 585
R1861 B.n1151 B.n1150 585
R1862 B.n74 B.n73 585
R1863 B.n1149 B.n74 585
R1864 B.n1147 B.n1146 585
R1865 B.n1148 B.n1147 585
R1866 B.n1145 B.n78 585
R1867 B.n81 B.n78 585
R1868 B.n1144 B.n1143 585
R1869 B.n1143 B.n1142 585
R1870 B.n80 B.n79 585
R1871 B.n1141 B.n80 585
R1872 B.n1139 B.n1138 585
R1873 B.n1140 B.n1139 585
R1874 B.n1137 B.n86 585
R1875 B.n86 B.n85 585
R1876 B.n1136 B.n1135 585
R1877 B.n1135 B.n1134 585
R1878 B.n88 B.n87 585
R1879 B.n1133 B.n88 585
R1880 B.n1131 B.n1130 585
R1881 B.n1132 B.n1131 585
R1882 B.n1129 B.n93 585
R1883 B.n93 B.n92 585
R1884 B.n1128 B.n1127 585
R1885 B.n1127 B.n1126 585
R1886 B.n95 B.n94 585
R1887 B.n1125 B.n95 585
R1888 B.n1123 B.n1122 585
R1889 B.n1124 B.n1123 585
R1890 B.n1121 B.n100 585
R1891 B.n100 B.n99 585
R1892 B.n1120 B.n1119 585
R1893 B.n1119 B.n1118 585
R1894 B.n102 B.n101 585
R1895 B.n1117 B.n102 585
R1896 B.n1115 B.n1114 585
R1897 B.n1116 B.n1115 585
R1898 B.n1113 B.n107 585
R1899 B.n107 B.n106 585
R1900 B.n1112 B.n1111 585
R1901 B.n1111 B.n1110 585
R1902 B.n109 B.n108 585
R1903 B.n1109 B.n109 585
R1904 B.n1107 B.n1106 585
R1905 B.n1108 B.n1107 585
R1906 B.n1105 B.n114 585
R1907 B.n114 B.n113 585
R1908 B.n1104 B.n1103 585
R1909 B.n1103 B.n1102 585
R1910 B.n116 B.n115 585
R1911 B.n1101 B.n116 585
R1912 B.n1099 B.n1098 585
R1913 B.n1100 B.n1099 585
R1914 B.n1097 B.n121 585
R1915 B.n121 B.n120 585
R1916 B.n1232 B.n1231 585
R1917 B.n1231 B.n1230 585
R1918 B.n803 B.n525 454.062
R1919 B.n1095 B.n121 454.062
R1920 B.n587 B.n523 454.062
R1921 B.n1092 B.n178 454.062
R1922 B.n584 B.t21 406.433
R1923 B.n179 B.t10 406.433
R1924 B.n582 B.t15 406.433
R1925 B.n181 B.t17 406.433
R1926 B.n585 B.t20 329.051
R1927 B.n180 B.t11 329.051
R1928 B.n583 B.t14 329.051
R1929 B.n182 B.t18 329.051
R1930 B.n584 B.t19 306.224
R1931 B.n582 B.t12 306.224
R1932 B.n181 B.t16 306.224
R1933 B.n179 B.t8 306.224
R1934 B.n1093 B.n176 256.663
R1935 B.n1093 B.n175 256.663
R1936 B.n1093 B.n174 256.663
R1937 B.n1093 B.n173 256.663
R1938 B.n1093 B.n172 256.663
R1939 B.n1093 B.n171 256.663
R1940 B.n1093 B.n170 256.663
R1941 B.n1093 B.n169 256.663
R1942 B.n1093 B.n168 256.663
R1943 B.n1093 B.n167 256.663
R1944 B.n1093 B.n166 256.663
R1945 B.n1093 B.n165 256.663
R1946 B.n1093 B.n164 256.663
R1947 B.n1093 B.n163 256.663
R1948 B.n1093 B.n162 256.663
R1949 B.n1093 B.n161 256.663
R1950 B.n1093 B.n160 256.663
R1951 B.n1093 B.n159 256.663
R1952 B.n1093 B.n158 256.663
R1953 B.n1093 B.n157 256.663
R1954 B.n1093 B.n156 256.663
R1955 B.n1093 B.n155 256.663
R1956 B.n1093 B.n154 256.663
R1957 B.n1093 B.n153 256.663
R1958 B.n1093 B.n152 256.663
R1959 B.n1093 B.n151 256.663
R1960 B.n1093 B.n150 256.663
R1961 B.n1093 B.n149 256.663
R1962 B.n1093 B.n148 256.663
R1963 B.n1093 B.n147 256.663
R1964 B.n1093 B.n146 256.663
R1965 B.n1093 B.n145 256.663
R1966 B.n1093 B.n144 256.663
R1967 B.n1093 B.n143 256.663
R1968 B.n1093 B.n142 256.663
R1969 B.n1093 B.n141 256.663
R1970 B.n1093 B.n140 256.663
R1971 B.n1093 B.n139 256.663
R1972 B.n1093 B.n138 256.663
R1973 B.n1093 B.n137 256.663
R1974 B.n1093 B.n136 256.663
R1975 B.n1093 B.n135 256.663
R1976 B.n1093 B.n134 256.663
R1977 B.n1093 B.n133 256.663
R1978 B.n1093 B.n132 256.663
R1979 B.n1093 B.n131 256.663
R1980 B.n1093 B.n130 256.663
R1981 B.n1093 B.n129 256.663
R1982 B.n1093 B.n128 256.663
R1983 B.n1093 B.n127 256.663
R1984 B.n1093 B.n126 256.663
R1985 B.n1093 B.n125 256.663
R1986 B.n1093 B.n124 256.663
R1987 B.n1094 B.n1093 256.663
R1988 B.n802 B.n801 256.663
R1989 B.n801 B.n528 256.663
R1990 B.n801 B.n529 256.663
R1991 B.n801 B.n530 256.663
R1992 B.n801 B.n531 256.663
R1993 B.n801 B.n532 256.663
R1994 B.n801 B.n533 256.663
R1995 B.n801 B.n534 256.663
R1996 B.n801 B.n535 256.663
R1997 B.n801 B.n536 256.663
R1998 B.n801 B.n537 256.663
R1999 B.n801 B.n538 256.663
R2000 B.n801 B.n539 256.663
R2001 B.n801 B.n540 256.663
R2002 B.n801 B.n541 256.663
R2003 B.n801 B.n542 256.663
R2004 B.n801 B.n543 256.663
R2005 B.n801 B.n544 256.663
R2006 B.n801 B.n545 256.663
R2007 B.n801 B.n546 256.663
R2008 B.n801 B.n547 256.663
R2009 B.n801 B.n548 256.663
R2010 B.n801 B.n549 256.663
R2011 B.n801 B.n550 256.663
R2012 B.n801 B.n551 256.663
R2013 B.n801 B.n552 256.663
R2014 B.n801 B.n553 256.663
R2015 B.n801 B.n554 256.663
R2016 B.n801 B.n555 256.663
R2017 B.n801 B.n556 256.663
R2018 B.n801 B.n557 256.663
R2019 B.n801 B.n558 256.663
R2020 B.n801 B.n559 256.663
R2021 B.n801 B.n560 256.663
R2022 B.n801 B.n561 256.663
R2023 B.n801 B.n562 256.663
R2024 B.n801 B.n563 256.663
R2025 B.n801 B.n564 256.663
R2026 B.n801 B.n565 256.663
R2027 B.n801 B.n566 256.663
R2028 B.n801 B.n567 256.663
R2029 B.n801 B.n568 256.663
R2030 B.n801 B.n569 256.663
R2031 B.n801 B.n570 256.663
R2032 B.n801 B.n571 256.663
R2033 B.n801 B.n572 256.663
R2034 B.n801 B.n573 256.663
R2035 B.n801 B.n574 256.663
R2036 B.n801 B.n575 256.663
R2037 B.n801 B.n576 256.663
R2038 B.n801 B.n577 256.663
R2039 B.n801 B.n578 256.663
R2040 B.n801 B.n579 256.663
R2041 B.n801 B.n580 256.663
R2042 B.n807 B.n525 163.367
R2043 B.n807 B.n519 163.367
R2044 B.n815 B.n519 163.367
R2045 B.n815 B.n517 163.367
R2046 B.n819 B.n517 163.367
R2047 B.n819 B.n511 163.367
R2048 B.n827 B.n511 163.367
R2049 B.n827 B.n509 163.367
R2050 B.n831 B.n509 163.367
R2051 B.n831 B.n503 163.367
R2052 B.n839 B.n503 163.367
R2053 B.n839 B.n501 163.367
R2054 B.n843 B.n501 163.367
R2055 B.n843 B.n495 163.367
R2056 B.n851 B.n495 163.367
R2057 B.n851 B.n493 163.367
R2058 B.n855 B.n493 163.367
R2059 B.n855 B.n487 163.367
R2060 B.n863 B.n487 163.367
R2061 B.n863 B.n485 163.367
R2062 B.n867 B.n485 163.367
R2063 B.n867 B.n479 163.367
R2064 B.n876 B.n479 163.367
R2065 B.n876 B.n477 163.367
R2066 B.n880 B.n477 163.367
R2067 B.n880 B.n472 163.367
R2068 B.n888 B.n472 163.367
R2069 B.n888 B.n470 163.367
R2070 B.n892 B.n470 163.367
R2071 B.n892 B.n464 163.367
R2072 B.n900 B.n464 163.367
R2073 B.n900 B.n462 163.367
R2074 B.n904 B.n462 163.367
R2075 B.n904 B.n456 163.367
R2076 B.n913 B.n456 163.367
R2077 B.n913 B.n454 163.367
R2078 B.n917 B.n454 163.367
R2079 B.n917 B.n449 163.367
R2080 B.n925 B.n449 163.367
R2081 B.n925 B.n447 163.367
R2082 B.n929 B.n447 163.367
R2083 B.n929 B.n441 163.367
R2084 B.n937 B.n441 163.367
R2085 B.n937 B.n439 163.367
R2086 B.n941 B.n439 163.367
R2087 B.n941 B.n433 163.367
R2088 B.n949 B.n433 163.367
R2089 B.n949 B.n431 163.367
R2090 B.n953 B.n431 163.367
R2091 B.n953 B.n425 163.367
R2092 B.n961 B.n425 163.367
R2093 B.n961 B.n423 163.367
R2094 B.n965 B.n423 163.367
R2095 B.n965 B.n417 163.367
R2096 B.n973 B.n417 163.367
R2097 B.n973 B.n415 163.367
R2098 B.n977 B.n415 163.367
R2099 B.n977 B.n409 163.367
R2100 B.n985 B.n409 163.367
R2101 B.n985 B.n407 163.367
R2102 B.n989 B.n407 163.367
R2103 B.n989 B.n401 163.367
R2104 B.n998 B.n401 163.367
R2105 B.n998 B.n399 163.367
R2106 B.n1002 B.n399 163.367
R2107 B.n1002 B.n2 163.367
R2108 B.n1231 B.n2 163.367
R2109 B.n1231 B.n3 163.367
R2110 B.n1227 B.n3 163.367
R2111 B.n1227 B.n9 163.367
R2112 B.n1223 B.n9 163.367
R2113 B.n1223 B.n11 163.367
R2114 B.n1219 B.n11 163.367
R2115 B.n1219 B.n16 163.367
R2116 B.n1215 B.n16 163.367
R2117 B.n1215 B.n18 163.367
R2118 B.n1211 B.n18 163.367
R2119 B.n1211 B.n23 163.367
R2120 B.n1207 B.n23 163.367
R2121 B.n1207 B.n25 163.367
R2122 B.n1203 B.n25 163.367
R2123 B.n1203 B.n30 163.367
R2124 B.n1199 B.n30 163.367
R2125 B.n1199 B.n32 163.367
R2126 B.n1195 B.n32 163.367
R2127 B.n1195 B.n37 163.367
R2128 B.n1191 B.n37 163.367
R2129 B.n1191 B.n39 163.367
R2130 B.n1187 B.n39 163.367
R2131 B.n1187 B.n44 163.367
R2132 B.n1183 B.n44 163.367
R2133 B.n1183 B.n46 163.367
R2134 B.n1179 B.n46 163.367
R2135 B.n1179 B.n51 163.367
R2136 B.n1175 B.n51 163.367
R2137 B.n1175 B.n53 163.367
R2138 B.n1171 B.n53 163.367
R2139 B.n1171 B.n57 163.367
R2140 B.n1167 B.n57 163.367
R2141 B.n1167 B.n59 163.367
R2142 B.n1163 B.n59 163.367
R2143 B.n1163 B.n65 163.367
R2144 B.n1159 B.n65 163.367
R2145 B.n1159 B.n67 163.367
R2146 B.n1155 B.n67 163.367
R2147 B.n1155 B.n72 163.367
R2148 B.n1151 B.n72 163.367
R2149 B.n1151 B.n74 163.367
R2150 B.n1147 B.n74 163.367
R2151 B.n1147 B.n78 163.367
R2152 B.n1143 B.n78 163.367
R2153 B.n1143 B.n80 163.367
R2154 B.n1139 B.n80 163.367
R2155 B.n1139 B.n86 163.367
R2156 B.n1135 B.n86 163.367
R2157 B.n1135 B.n88 163.367
R2158 B.n1131 B.n88 163.367
R2159 B.n1131 B.n93 163.367
R2160 B.n1127 B.n93 163.367
R2161 B.n1127 B.n95 163.367
R2162 B.n1123 B.n95 163.367
R2163 B.n1123 B.n100 163.367
R2164 B.n1119 B.n100 163.367
R2165 B.n1119 B.n102 163.367
R2166 B.n1115 B.n102 163.367
R2167 B.n1115 B.n107 163.367
R2168 B.n1111 B.n107 163.367
R2169 B.n1111 B.n109 163.367
R2170 B.n1107 B.n109 163.367
R2171 B.n1107 B.n114 163.367
R2172 B.n1103 B.n114 163.367
R2173 B.n1103 B.n116 163.367
R2174 B.n1099 B.n116 163.367
R2175 B.n1099 B.n121 163.367
R2176 B.n800 B.n527 163.367
R2177 B.n800 B.n581 163.367
R2178 B.n796 B.n795 163.367
R2179 B.n792 B.n791 163.367
R2180 B.n788 B.n787 163.367
R2181 B.n784 B.n783 163.367
R2182 B.n780 B.n779 163.367
R2183 B.n776 B.n775 163.367
R2184 B.n772 B.n771 163.367
R2185 B.n768 B.n767 163.367
R2186 B.n764 B.n763 163.367
R2187 B.n760 B.n759 163.367
R2188 B.n756 B.n755 163.367
R2189 B.n752 B.n751 163.367
R2190 B.n748 B.n747 163.367
R2191 B.n744 B.n743 163.367
R2192 B.n740 B.n739 163.367
R2193 B.n736 B.n735 163.367
R2194 B.n732 B.n731 163.367
R2195 B.n728 B.n727 163.367
R2196 B.n724 B.n723 163.367
R2197 B.n720 B.n719 163.367
R2198 B.n716 B.n715 163.367
R2199 B.n712 B.n711 163.367
R2200 B.n708 B.n707 163.367
R2201 B.n703 B.n702 163.367
R2202 B.n699 B.n698 163.367
R2203 B.n695 B.n694 163.367
R2204 B.n691 B.n690 163.367
R2205 B.n687 B.n686 163.367
R2206 B.n683 B.n682 163.367
R2207 B.n679 B.n678 163.367
R2208 B.n675 B.n674 163.367
R2209 B.n671 B.n670 163.367
R2210 B.n667 B.n666 163.367
R2211 B.n663 B.n662 163.367
R2212 B.n659 B.n658 163.367
R2213 B.n655 B.n654 163.367
R2214 B.n651 B.n650 163.367
R2215 B.n647 B.n646 163.367
R2216 B.n643 B.n642 163.367
R2217 B.n639 B.n638 163.367
R2218 B.n635 B.n634 163.367
R2219 B.n631 B.n630 163.367
R2220 B.n627 B.n626 163.367
R2221 B.n623 B.n622 163.367
R2222 B.n619 B.n618 163.367
R2223 B.n615 B.n614 163.367
R2224 B.n611 B.n610 163.367
R2225 B.n607 B.n606 163.367
R2226 B.n603 B.n602 163.367
R2227 B.n599 B.n598 163.367
R2228 B.n595 B.n594 163.367
R2229 B.n591 B.n590 163.367
R2230 B.n809 B.n523 163.367
R2231 B.n809 B.n521 163.367
R2232 B.n813 B.n521 163.367
R2233 B.n813 B.n515 163.367
R2234 B.n821 B.n515 163.367
R2235 B.n821 B.n513 163.367
R2236 B.n825 B.n513 163.367
R2237 B.n825 B.n507 163.367
R2238 B.n833 B.n507 163.367
R2239 B.n833 B.n505 163.367
R2240 B.n837 B.n505 163.367
R2241 B.n837 B.n499 163.367
R2242 B.n845 B.n499 163.367
R2243 B.n845 B.n497 163.367
R2244 B.n849 B.n497 163.367
R2245 B.n849 B.n491 163.367
R2246 B.n857 B.n491 163.367
R2247 B.n857 B.n489 163.367
R2248 B.n861 B.n489 163.367
R2249 B.n861 B.n483 163.367
R2250 B.n869 B.n483 163.367
R2251 B.n869 B.n481 163.367
R2252 B.n873 B.n481 163.367
R2253 B.n873 B.n476 163.367
R2254 B.n882 B.n476 163.367
R2255 B.n882 B.n474 163.367
R2256 B.n886 B.n474 163.367
R2257 B.n886 B.n468 163.367
R2258 B.n894 B.n468 163.367
R2259 B.n894 B.n466 163.367
R2260 B.n898 B.n466 163.367
R2261 B.n898 B.n460 163.367
R2262 B.n906 B.n460 163.367
R2263 B.n906 B.n458 163.367
R2264 B.n910 B.n458 163.367
R2265 B.n910 B.n453 163.367
R2266 B.n919 B.n453 163.367
R2267 B.n919 B.n451 163.367
R2268 B.n923 B.n451 163.367
R2269 B.n923 B.n445 163.367
R2270 B.n931 B.n445 163.367
R2271 B.n931 B.n443 163.367
R2272 B.n935 B.n443 163.367
R2273 B.n935 B.n437 163.367
R2274 B.n943 B.n437 163.367
R2275 B.n943 B.n435 163.367
R2276 B.n947 B.n435 163.367
R2277 B.n947 B.n429 163.367
R2278 B.n955 B.n429 163.367
R2279 B.n955 B.n427 163.367
R2280 B.n959 B.n427 163.367
R2281 B.n959 B.n421 163.367
R2282 B.n967 B.n421 163.367
R2283 B.n967 B.n419 163.367
R2284 B.n971 B.n419 163.367
R2285 B.n971 B.n413 163.367
R2286 B.n979 B.n413 163.367
R2287 B.n979 B.n411 163.367
R2288 B.n983 B.n411 163.367
R2289 B.n983 B.n405 163.367
R2290 B.n991 B.n405 163.367
R2291 B.n991 B.n403 163.367
R2292 B.n996 B.n403 163.367
R2293 B.n996 B.n397 163.367
R2294 B.n1004 B.n397 163.367
R2295 B.n1005 B.n1004 163.367
R2296 B.n1005 B.n5 163.367
R2297 B.n6 B.n5 163.367
R2298 B.n7 B.n6 163.367
R2299 B.n1010 B.n7 163.367
R2300 B.n1010 B.n12 163.367
R2301 B.n13 B.n12 163.367
R2302 B.n14 B.n13 163.367
R2303 B.n1015 B.n14 163.367
R2304 B.n1015 B.n19 163.367
R2305 B.n20 B.n19 163.367
R2306 B.n21 B.n20 163.367
R2307 B.n1020 B.n21 163.367
R2308 B.n1020 B.n26 163.367
R2309 B.n27 B.n26 163.367
R2310 B.n28 B.n27 163.367
R2311 B.n1025 B.n28 163.367
R2312 B.n1025 B.n33 163.367
R2313 B.n34 B.n33 163.367
R2314 B.n35 B.n34 163.367
R2315 B.n1030 B.n35 163.367
R2316 B.n1030 B.n40 163.367
R2317 B.n41 B.n40 163.367
R2318 B.n42 B.n41 163.367
R2319 B.n1035 B.n42 163.367
R2320 B.n1035 B.n47 163.367
R2321 B.n48 B.n47 163.367
R2322 B.n49 B.n48 163.367
R2323 B.n1040 B.n49 163.367
R2324 B.n1040 B.n54 163.367
R2325 B.n55 B.n54 163.367
R2326 B.n56 B.n55 163.367
R2327 B.n1045 B.n56 163.367
R2328 B.n1045 B.n61 163.367
R2329 B.n62 B.n61 163.367
R2330 B.n63 B.n62 163.367
R2331 B.n1050 B.n63 163.367
R2332 B.n1050 B.n68 163.367
R2333 B.n69 B.n68 163.367
R2334 B.n70 B.n69 163.367
R2335 B.n1055 B.n70 163.367
R2336 B.n1055 B.n75 163.367
R2337 B.n76 B.n75 163.367
R2338 B.n77 B.n76 163.367
R2339 B.n1060 B.n77 163.367
R2340 B.n1060 B.n82 163.367
R2341 B.n83 B.n82 163.367
R2342 B.n84 B.n83 163.367
R2343 B.n1065 B.n84 163.367
R2344 B.n1065 B.n89 163.367
R2345 B.n90 B.n89 163.367
R2346 B.n91 B.n90 163.367
R2347 B.n1070 B.n91 163.367
R2348 B.n1070 B.n96 163.367
R2349 B.n97 B.n96 163.367
R2350 B.n98 B.n97 163.367
R2351 B.n1075 B.n98 163.367
R2352 B.n1075 B.n103 163.367
R2353 B.n104 B.n103 163.367
R2354 B.n105 B.n104 163.367
R2355 B.n1080 B.n105 163.367
R2356 B.n1080 B.n110 163.367
R2357 B.n111 B.n110 163.367
R2358 B.n112 B.n111 163.367
R2359 B.n1085 B.n112 163.367
R2360 B.n1085 B.n117 163.367
R2361 B.n118 B.n117 163.367
R2362 B.n119 B.n118 163.367
R2363 B.n178 B.n119 163.367
R2364 B.n184 B.n123 163.367
R2365 B.n188 B.n187 163.367
R2366 B.n192 B.n191 163.367
R2367 B.n196 B.n195 163.367
R2368 B.n200 B.n199 163.367
R2369 B.n204 B.n203 163.367
R2370 B.n208 B.n207 163.367
R2371 B.n212 B.n211 163.367
R2372 B.n216 B.n215 163.367
R2373 B.n220 B.n219 163.367
R2374 B.n224 B.n223 163.367
R2375 B.n228 B.n227 163.367
R2376 B.n232 B.n231 163.367
R2377 B.n236 B.n235 163.367
R2378 B.n240 B.n239 163.367
R2379 B.n244 B.n243 163.367
R2380 B.n248 B.n247 163.367
R2381 B.n252 B.n251 163.367
R2382 B.n256 B.n255 163.367
R2383 B.n260 B.n259 163.367
R2384 B.n264 B.n263 163.367
R2385 B.n268 B.n267 163.367
R2386 B.n272 B.n271 163.367
R2387 B.n276 B.n275 163.367
R2388 B.n280 B.n279 163.367
R2389 B.n284 B.n283 163.367
R2390 B.n288 B.n287 163.367
R2391 B.n292 B.n291 163.367
R2392 B.n296 B.n295 163.367
R2393 B.n301 B.n300 163.367
R2394 B.n305 B.n304 163.367
R2395 B.n309 B.n308 163.367
R2396 B.n313 B.n312 163.367
R2397 B.n317 B.n316 163.367
R2398 B.n321 B.n320 163.367
R2399 B.n325 B.n324 163.367
R2400 B.n329 B.n328 163.367
R2401 B.n333 B.n332 163.367
R2402 B.n337 B.n336 163.367
R2403 B.n341 B.n340 163.367
R2404 B.n345 B.n344 163.367
R2405 B.n349 B.n348 163.367
R2406 B.n353 B.n352 163.367
R2407 B.n357 B.n356 163.367
R2408 B.n361 B.n360 163.367
R2409 B.n365 B.n364 163.367
R2410 B.n369 B.n368 163.367
R2411 B.n373 B.n372 163.367
R2412 B.n377 B.n376 163.367
R2413 B.n381 B.n380 163.367
R2414 B.n385 B.n384 163.367
R2415 B.n389 B.n388 163.367
R2416 B.n393 B.n392 163.367
R2417 B.n1092 B.n177 163.367
R2418 B.n585 B.n584 77.3823
R2419 B.n583 B.n582 77.3823
R2420 B.n182 B.n181 77.3823
R2421 B.n180 B.n179 77.3823
R2422 B.n803 B.n802 71.676
R2423 B.n581 B.n528 71.676
R2424 B.n795 B.n529 71.676
R2425 B.n791 B.n530 71.676
R2426 B.n787 B.n531 71.676
R2427 B.n783 B.n532 71.676
R2428 B.n779 B.n533 71.676
R2429 B.n775 B.n534 71.676
R2430 B.n771 B.n535 71.676
R2431 B.n767 B.n536 71.676
R2432 B.n763 B.n537 71.676
R2433 B.n759 B.n538 71.676
R2434 B.n755 B.n539 71.676
R2435 B.n751 B.n540 71.676
R2436 B.n747 B.n541 71.676
R2437 B.n743 B.n542 71.676
R2438 B.n739 B.n543 71.676
R2439 B.n735 B.n544 71.676
R2440 B.n731 B.n545 71.676
R2441 B.n727 B.n546 71.676
R2442 B.n723 B.n547 71.676
R2443 B.n719 B.n548 71.676
R2444 B.n715 B.n549 71.676
R2445 B.n711 B.n550 71.676
R2446 B.n707 B.n551 71.676
R2447 B.n702 B.n552 71.676
R2448 B.n698 B.n553 71.676
R2449 B.n694 B.n554 71.676
R2450 B.n690 B.n555 71.676
R2451 B.n686 B.n556 71.676
R2452 B.n682 B.n557 71.676
R2453 B.n678 B.n558 71.676
R2454 B.n674 B.n559 71.676
R2455 B.n670 B.n560 71.676
R2456 B.n666 B.n561 71.676
R2457 B.n662 B.n562 71.676
R2458 B.n658 B.n563 71.676
R2459 B.n654 B.n564 71.676
R2460 B.n650 B.n565 71.676
R2461 B.n646 B.n566 71.676
R2462 B.n642 B.n567 71.676
R2463 B.n638 B.n568 71.676
R2464 B.n634 B.n569 71.676
R2465 B.n630 B.n570 71.676
R2466 B.n626 B.n571 71.676
R2467 B.n622 B.n572 71.676
R2468 B.n618 B.n573 71.676
R2469 B.n614 B.n574 71.676
R2470 B.n610 B.n575 71.676
R2471 B.n606 B.n576 71.676
R2472 B.n602 B.n577 71.676
R2473 B.n598 B.n578 71.676
R2474 B.n594 B.n579 71.676
R2475 B.n590 B.n580 71.676
R2476 B.n1095 B.n1094 71.676
R2477 B.n184 B.n124 71.676
R2478 B.n188 B.n125 71.676
R2479 B.n192 B.n126 71.676
R2480 B.n196 B.n127 71.676
R2481 B.n200 B.n128 71.676
R2482 B.n204 B.n129 71.676
R2483 B.n208 B.n130 71.676
R2484 B.n212 B.n131 71.676
R2485 B.n216 B.n132 71.676
R2486 B.n220 B.n133 71.676
R2487 B.n224 B.n134 71.676
R2488 B.n228 B.n135 71.676
R2489 B.n232 B.n136 71.676
R2490 B.n236 B.n137 71.676
R2491 B.n240 B.n138 71.676
R2492 B.n244 B.n139 71.676
R2493 B.n248 B.n140 71.676
R2494 B.n252 B.n141 71.676
R2495 B.n256 B.n142 71.676
R2496 B.n260 B.n143 71.676
R2497 B.n264 B.n144 71.676
R2498 B.n268 B.n145 71.676
R2499 B.n272 B.n146 71.676
R2500 B.n276 B.n147 71.676
R2501 B.n280 B.n148 71.676
R2502 B.n284 B.n149 71.676
R2503 B.n288 B.n150 71.676
R2504 B.n292 B.n151 71.676
R2505 B.n296 B.n152 71.676
R2506 B.n301 B.n153 71.676
R2507 B.n305 B.n154 71.676
R2508 B.n309 B.n155 71.676
R2509 B.n313 B.n156 71.676
R2510 B.n317 B.n157 71.676
R2511 B.n321 B.n158 71.676
R2512 B.n325 B.n159 71.676
R2513 B.n329 B.n160 71.676
R2514 B.n333 B.n161 71.676
R2515 B.n337 B.n162 71.676
R2516 B.n341 B.n163 71.676
R2517 B.n345 B.n164 71.676
R2518 B.n349 B.n165 71.676
R2519 B.n353 B.n166 71.676
R2520 B.n357 B.n167 71.676
R2521 B.n361 B.n168 71.676
R2522 B.n365 B.n169 71.676
R2523 B.n369 B.n170 71.676
R2524 B.n373 B.n171 71.676
R2525 B.n377 B.n172 71.676
R2526 B.n381 B.n173 71.676
R2527 B.n385 B.n174 71.676
R2528 B.n389 B.n175 71.676
R2529 B.n393 B.n176 71.676
R2530 B.n177 B.n176 71.676
R2531 B.n392 B.n175 71.676
R2532 B.n388 B.n174 71.676
R2533 B.n384 B.n173 71.676
R2534 B.n380 B.n172 71.676
R2535 B.n376 B.n171 71.676
R2536 B.n372 B.n170 71.676
R2537 B.n368 B.n169 71.676
R2538 B.n364 B.n168 71.676
R2539 B.n360 B.n167 71.676
R2540 B.n356 B.n166 71.676
R2541 B.n352 B.n165 71.676
R2542 B.n348 B.n164 71.676
R2543 B.n344 B.n163 71.676
R2544 B.n340 B.n162 71.676
R2545 B.n336 B.n161 71.676
R2546 B.n332 B.n160 71.676
R2547 B.n328 B.n159 71.676
R2548 B.n324 B.n158 71.676
R2549 B.n320 B.n157 71.676
R2550 B.n316 B.n156 71.676
R2551 B.n312 B.n155 71.676
R2552 B.n308 B.n154 71.676
R2553 B.n304 B.n153 71.676
R2554 B.n300 B.n152 71.676
R2555 B.n295 B.n151 71.676
R2556 B.n291 B.n150 71.676
R2557 B.n287 B.n149 71.676
R2558 B.n283 B.n148 71.676
R2559 B.n279 B.n147 71.676
R2560 B.n275 B.n146 71.676
R2561 B.n271 B.n145 71.676
R2562 B.n267 B.n144 71.676
R2563 B.n263 B.n143 71.676
R2564 B.n259 B.n142 71.676
R2565 B.n255 B.n141 71.676
R2566 B.n251 B.n140 71.676
R2567 B.n247 B.n139 71.676
R2568 B.n243 B.n138 71.676
R2569 B.n239 B.n137 71.676
R2570 B.n235 B.n136 71.676
R2571 B.n231 B.n135 71.676
R2572 B.n227 B.n134 71.676
R2573 B.n223 B.n133 71.676
R2574 B.n219 B.n132 71.676
R2575 B.n215 B.n131 71.676
R2576 B.n211 B.n130 71.676
R2577 B.n207 B.n129 71.676
R2578 B.n203 B.n128 71.676
R2579 B.n199 B.n127 71.676
R2580 B.n195 B.n126 71.676
R2581 B.n191 B.n125 71.676
R2582 B.n187 B.n124 71.676
R2583 B.n1094 B.n123 71.676
R2584 B.n802 B.n527 71.676
R2585 B.n796 B.n528 71.676
R2586 B.n792 B.n529 71.676
R2587 B.n788 B.n530 71.676
R2588 B.n784 B.n531 71.676
R2589 B.n780 B.n532 71.676
R2590 B.n776 B.n533 71.676
R2591 B.n772 B.n534 71.676
R2592 B.n768 B.n535 71.676
R2593 B.n764 B.n536 71.676
R2594 B.n760 B.n537 71.676
R2595 B.n756 B.n538 71.676
R2596 B.n752 B.n539 71.676
R2597 B.n748 B.n540 71.676
R2598 B.n744 B.n541 71.676
R2599 B.n740 B.n542 71.676
R2600 B.n736 B.n543 71.676
R2601 B.n732 B.n544 71.676
R2602 B.n728 B.n545 71.676
R2603 B.n724 B.n546 71.676
R2604 B.n720 B.n547 71.676
R2605 B.n716 B.n548 71.676
R2606 B.n712 B.n549 71.676
R2607 B.n708 B.n550 71.676
R2608 B.n703 B.n551 71.676
R2609 B.n699 B.n552 71.676
R2610 B.n695 B.n553 71.676
R2611 B.n691 B.n554 71.676
R2612 B.n687 B.n555 71.676
R2613 B.n683 B.n556 71.676
R2614 B.n679 B.n557 71.676
R2615 B.n675 B.n558 71.676
R2616 B.n671 B.n559 71.676
R2617 B.n667 B.n560 71.676
R2618 B.n663 B.n561 71.676
R2619 B.n659 B.n562 71.676
R2620 B.n655 B.n563 71.676
R2621 B.n651 B.n564 71.676
R2622 B.n647 B.n565 71.676
R2623 B.n643 B.n566 71.676
R2624 B.n639 B.n567 71.676
R2625 B.n635 B.n568 71.676
R2626 B.n631 B.n569 71.676
R2627 B.n627 B.n570 71.676
R2628 B.n623 B.n571 71.676
R2629 B.n619 B.n572 71.676
R2630 B.n615 B.n573 71.676
R2631 B.n611 B.n574 71.676
R2632 B.n607 B.n575 71.676
R2633 B.n603 B.n576 71.676
R2634 B.n599 B.n577 71.676
R2635 B.n595 B.n578 71.676
R2636 B.n591 B.n579 71.676
R2637 B.n587 B.n580 71.676
R2638 B.n801 B.n524 59.9355
R2639 B.n1093 B.n120 59.9355
R2640 B.n586 B.n585 59.5399
R2641 B.n705 B.n583 59.5399
R2642 B.n183 B.n182 59.5399
R2643 B.n298 B.n180 59.5399
R2644 B.n808 B.n524 37.3912
R2645 B.n808 B.n520 37.3912
R2646 B.n814 B.n520 37.3912
R2647 B.n814 B.n516 37.3912
R2648 B.n820 B.n516 37.3912
R2649 B.n820 B.n512 37.3912
R2650 B.n826 B.n512 37.3912
R2651 B.n826 B.n508 37.3912
R2652 B.n832 B.n508 37.3912
R2653 B.n838 B.n504 37.3912
R2654 B.n838 B.n500 37.3912
R2655 B.n844 B.n500 37.3912
R2656 B.n844 B.n496 37.3912
R2657 B.n850 B.n496 37.3912
R2658 B.n850 B.n492 37.3912
R2659 B.n856 B.n492 37.3912
R2660 B.n856 B.n488 37.3912
R2661 B.n862 B.n488 37.3912
R2662 B.n862 B.n484 37.3912
R2663 B.n868 B.n484 37.3912
R2664 B.n868 B.n480 37.3912
R2665 B.n875 B.n480 37.3912
R2666 B.n875 B.n874 37.3912
R2667 B.n881 B.n473 37.3912
R2668 B.n887 B.n473 37.3912
R2669 B.n887 B.n469 37.3912
R2670 B.n893 B.n469 37.3912
R2671 B.n893 B.n465 37.3912
R2672 B.n899 B.n465 37.3912
R2673 B.n899 B.n461 37.3912
R2674 B.n905 B.n461 37.3912
R2675 B.n905 B.n457 37.3912
R2676 B.n912 B.n457 37.3912
R2677 B.n912 B.n911 37.3912
R2678 B.n918 B.n450 37.3912
R2679 B.n924 B.n450 37.3912
R2680 B.n924 B.n446 37.3912
R2681 B.n930 B.n446 37.3912
R2682 B.n930 B.n442 37.3912
R2683 B.n936 B.n442 37.3912
R2684 B.n936 B.n438 37.3912
R2685 B.n942 B.n438 37.3912
R2686 B.n942 B.n434 37.3912
R2687 B.n948 B.n434 37.3912
R2688 B.n954 B.n430 37.3912
R2689 B.n954 B.n426 37.3912
R2690 B.n960 B.n426 37.3912
R2691 B.n960 B.n422 37.3912
R2692 B.n966 B.n422 37.3912
R2693 B.n966 B.n418 37.3912
R2694 B.n972 B.n418 37.3912
R2695 B.n972 B.n414 37.3912
R2696 B.n978 B.n414 37.3912
R2697 B.n978 B.n410 37.3912
R2698 B.n984 B.n410 37.3912
R2699 B.n990 B.n406 37.3912
R2700 B.n990 B.n402 37.3912
R2701 B.n997 B.n402 37.3912
R2702 B.n997 B.n398 37.3912
R2703 B.n1003 B.n398 37.3912
R2704 B.n1003 B.n4 37.3912
R2705 B.n1230 B.n4 37.3912
R2706 B.n1230 B.n1229 37.3912
R2707 B.n1229 B.n1228 37.3912
R2708 B.n1228 B.n8 37.3912
R2709 B.n1222 B.n8 37.3912
R2710 B.n1222 B.n1221 37.3912
R2711 B.n1221 B.n1220 37.3912
R2712 B.n1220 B.n15 37.3912
R2713 B.n1214 B.n1213 37.3912
R2714 B.n1213 B.n1212 37.3912
R2715 B.n1212 B.n22 37.3912
R2716 B.n1206 B.n22 37.3912
R2717 B.n1206 B.n1205 37.3912
R2718 B.n1205 B.n1204 37.3912
R2719 B.n1204 B.n29 37.3912
R2720 B.n1198 B.n29 37.3912
R2721 B.n1198 B.n1197 37.3912
R2722 B.n1197 B.n1196 37.3912
R2723 B.n1196 B.n36 37.3912
R2724 B.n1190 B.n1189 37.3912
R2725 B.n1189 B.n1188 37.3912
R2726 B.n1188 B.n43 37.3912
R2727 B.n1182 B.n43 37.3912
R2728 B.n1182 B.n1181 37.3912
R2729 B.n1181 B.n1180 37.3912
R2730 B.n1180 B.n50 37.3912
R2731 B.n1174 B.n50 37.3912
R2732 B.n1174 B.n1173 37.3912
R2733 B.n1173 B.n1172 37.3912
R2734 B.n1166 B.n60 37.3912
R2735 B.n1166 B.n1165 37.3912
R2736 B.n1165 B.n1164 37.3912
R2737 B.n1164 B.n64 37.3912
R2738 B.n1158 B.n64 37.3912
R2739 B.n1158 B.n1157 37.3912
R2740 B.n1157 B.n1156 37.3912
R2741 B.n1156 B.n71 37.3912
R2742 B.n1150 B.n71 37.3912
R2743 B.n1150 B.n1149 37.3912
R2744 B.n1149 B.n1148 37.3912
R2745 B.n1142 B.n81 37.3912
R2746 B.n1142 B.n1141 37.3912
R2747 B.n1141 B.n1140 37.3912
R2748 B.n1140 B.n85 37.3912
R2749 B.n1134 B.n85 37.3912
R2750 B.n1134 B.n1133 37.3912
R2751 B.n1133 B.n1132 37.3912
R2752 B.n1132 B.n92 37.3912
R2753 B.n1126 B.n92 37.3912
R2754 B.n1126 B.n1125 37.3912
R2755 B.n1125 B.n1124 37.3912
R2756 B.n1124 B.n99 37.3912
R2757 B.n1118 B.n99 37.3912
R2758 B.n1118 B.n1117 37.3912
R2759 B.n1116 B.n106 37.3912
R2760 B.n1110 B.n106 37.3912
R2761 B.n1110 B.n1109 37.3912
R2762 B.n1109 B.n1108 37.3912
R2763 B.n1108 B.n113 37.3912
R2764 B.n1102 B.n113 37.3912
R2765 B.n1102 B.n1101 37.3912
R2766 B.n1101 B.n1100 37.3912
R2767 B.n1100 B.n120 37.3912
R2768 B.n918 B.t6 35.1917
R2769 B.n1172 B.t4 35.1917
R2770 B.n948 B.t0 29.6931
R2771 B.n1190 B.t3 29.6931
R2772 B.n1097 B.n1096 29.5029
R2773 B.n588 B.n522 29.5029
R2774 B.n805 B.n804 29.5029
R2775 B.n1091 B.n1090 29.5029
R2776 B.n881 B.t7 25.2942
R2777 B.n1148 B.t2 25.2942
R2778 B.t13 B.n504 23.0947
R2779 B.n1117 B.t9 23.0947
R2780 B.n984 B.t5 19.7956
R2781 B.n1214 B.t1 19.7956
R2782 B B.n1232 18.0485
R2783 B.t5 B.n406 17.5961
R2784 B.t1 B.n15 17.5961
R2785 B.n832 B.t13 14.2969
R2786 B.t9 B.n1116 14.2969
R2787 B.n874 B.t7 12.0975
R2788 B.n81 B.t2 12.0975
R2789 B.n1096 B.n122 10.6151
R2790 B.n185 B.n122 10.6151
R2791 B.n186 B.n185 10.6151
R2792 B.n189 B.n186 10.6151
R2793 B.n190 B.n189 10.6151
R2794 B.n193 B.n190 10.6151
R2795 B.n194 B.n193 10.6151
R2796 B.n197 B.n194 10.6151
R2797 B.n198 B.n197 10.6151
R2798 B.n201 B.n198 10.6151
R2799 B.n202 B.n201 10.6151
R2800 B.n205 B.n202 10.6151
R2801 B.n206 B.n205 10.6151
R2802 B.n209 B.n206 10.6151
R2803 B.n210 B.n209 10.6151
R2804 B.n213 B.n210 10.6151
R2805 B.n214 B.n213 10.6151
R2806 B.n217 B.n214 10.6151
R2807 B.n218 B.n217 10.6151
R2808 B.n221 B.n218 10.6151
R2809 B.n222 B.n221 10.6151
R2810 B.n225 B.n222 10.6151
R2811 B.n226 B.n225 10.6151
R2812 B.n229 B.n226 10.6151
R2813 B.n230 B.n229 10.6151
R2814 B.n233 B.n230 10.6151
R2815 B.n234 B.n233 10.6151
R2816 B.n237 B.n234 10.6151
R2817 B.n238 B.n237 10.6151
R2818 B.n241 B.n238 10.6151
R2819 B.n242 B.n241 10.6151
R2820 B.n245 B.n242 10.6151
R2821 B.n246 B.n245 10.6151
R2822 B.n249 B.n246 10.6151
R2823 B.n250 B.n249 10.6151
R2824 B.n253 B.n250 10.6151
R2825 B.n254 B.n253 10.6151
R2826 B.n257 B.n254 10.6151
R2827 B.n258 B.n257 10.6151
R2828 B.n261 B.n258 10.6151
R2829 B.n262 B.n261 10.6151
R2830 B.n265 B.n262 10.6151
R2831 B.n266 B.n265 10.6151
R2832 B.n269 B.n266 10.6151
R2833 B.n270 B.n269 10.6151
R2834 B.n273 B.n270 10.6151
R2835 B.n274 B.n273 10.6151
R2836 B.n277 B.n274 10.6151
R2837 B.n278 B.n277 10.6151
R2838 B.n282 B.n281 10.6151
R2839 B.n285 B.n282 10.6151
R2840 B.n286 B.n285 10.6151
R2841 B.n289 B.n286 10.6151
R2842 B.n290 B.n289 10.6151
R2843 B.n293 B.n290 10.6151
R2844 B.n294 B.n293 10.6151
R2845 B.n297 B.n294 10.6151
R2846 B.n302 B.n299 10.6151
R2847 B.n303 B.n302 10.6151
R2848 B.n306 B.n303 10.6151
R2849 B.n307 B.n306 10.6151
R2850 B.n310 B.n307 10.6151
R2851 B.n311 B.n310 10.6151
R2852 B.n314 B.n311 10.6151
R2853 B.n315 B.n314 10.6151
R2854 B.n318 B.n315 10.6151
R2855 B.n319 B.n318 10.6151
R2856 B.n322 B.n319 10.6151
R2857 B.n323 B.n322 10.6151
R2858 B.n326 B.n323 10.6151
R2859 B.n327 B.n326 10.6151
R2860 B.n330 B.n327 10.6151
R2861 B.n331 B.n330 10.6151
R2862 B.n334 B.n331 10.6151
R2863 B.n335 B.n334 10.6151
R2864 B.n338 B.n335 10.6151
R2865 B.n339 B.n338 10.6151
R2866 B.n342 B.n339 10.6151
R2867 B.n343 B.n342 10.6151
R2868 B.n346 B.n343 10.6151
R2869 B.n347 B.n346 10.6151
R2870 B.n350 B.n347 10.6151
R2871 B.n351 B.n350 10.6151
R2872 B.n354 B.n351 10.6151
R2873 B.n355 B.n354 10.6151
R2874 B.n358 B.n355 10.6151
R2875 B.n359 B.n358 10.6151
R2876 B.n362 B.n359 10.6151
R2877 B.n363 B.n362 10.6151
R2878 B.n366 B.n363 10.6151
R2879 B.n367 B.n366 10.6151
R2880 B.n370 B.n367 10.6151
R2881 B.n371 B.n370 10.6151
R2882 B.n374 B.n371 10.6151
R2883 B.n375 B.n374 10.6151
R2884 B.n378 B.n375 10.6151
R2885 B.n379 B.n378 10.6151
R2886 B.n382 B.n379 10.6151
R2887 B.n383 B.n382 10.6151
R2888 B.n386 B.n383 10.6151
R2889 B.n387 B.n386 10.6151
R2890 B.n390 B.n387 10.6151
R2891 B.n391 B.n390 10.6151
R2892 B.n394 B.n391 10.6151
R2893 B.n395 B.n394 10.6151
R2894 B.n1091 B.n395 10.6151
R2895 B.n810 B.n522 10.6151
R2896 B.n811 B.n810 10.6151
R2897 B.n812 B.n811 10.6151
R2898 B.n812 B.n514 10.6151
R2899 B.n822 B.n514 10.6151
R2900 B.n823 B.n822 10.6151
R2901 B.n824 B.n823 10.6151
R2902 B.n824 B.n506 10.6151
R2903 B.n834 B.n506 10.6151
R2904 B.n835 B.n834 10.6151
R2905 B.n836 B.n835 10.6151
R2906 B.n836 B.n498 10.6151
R2907 B.n846 B.n498 10.6151
R2908 B.n847 B.n846 10.6151
R2909 B.n848 B.n847 10.6151
R2910 B.n848 B.n490 10.6151
R2911 B.n858 B.n490 10.6151
R2912 B.n859 B.n858 10.6151
R2913 B.n860 B.n859 10.6151
R2914 B.n860 B.n482 10.6151
R2915 B.n870 B.n482 10.6151
R2916 B.n871 B.n870 10.6151
R2917 B.n872 B.n871 10.6151
R2918 B.n872 B.n475 10.6151
R2919 B.n883 B.n475 10.6151
R2920 B.n884 B.n883 10.6151
R2921 B.n885 B.n884 10.6151
R2922 B.n885 B.n467 10.6151
R2923 B.n895 B.n467 10.6151
R2924 B.n896 B.n895 10.6151
R2925 B.n897 B.n896 10.6151
R2926 B.n897 B.n459 10.6151
R2927 B.n907 B.n459 10.6151
R2928 B.n908 B.n907 10.6151
R2929 B.n909 B.n908 10.6151
R2930 B.n909 B.n452 10.6151
R2931 B.n920 B.n452 10.6151
R2932 B.n921 B.n920 10.6151
R2933 B.n922 B.n921 10.6151
R2934 B.n922 B.n444 10.6151
R2935 B.n932 B.n444 10.6151
R2936 B.n933 B.n932 10.6151
R2937 B.n934 B.n933 10.6151
R2938 B.n934 B.n436 10.6151
R2939 B.n944 B.n436 10.6151
R2940 B.n945 B.n944 10.6151
R2941 B.n946 B.n945 10.6151
R2942 B.n946 B.n428 10.6151
R2943 B.n956 B.n428 10.6151
R2944 B.n957 B.n956 10.6151
R2945 B.n958 B.n957 10.6151
R2946 B.n958 B.n420 10.6151
R2947 B.n968 B.n420 10.6151
R2948 B.n969 B.n968 10.6151
R2949 B.n970 B.n969 10.6151
R2950 B.n970 B.n412 10.6151
R2951 B.n980 B.n412 10.6151
R2952 B.n981 B.n980 10.6151
R2953 B.n982 B.n981 10.6151
R2954 B.n982 B.n404 10.6151
R2955 B.n992 B.n404 10.6151
R2956 B.n993 B.n992 10.6151
R2957 B.n995 B.n993 10.6151
R2958 B.n995 B.n994 10.6151
R2959 B.n994 B.n396 10.6151
R2960 B.n1006 B.n396 10.6151
R2961 B.n1007 B.n1006 10.6151
R2962 B.n1008 B.n1007 10.6151
R2963 B.n1009 B.n1008 10.6151
R2964 B.n1011 B.n1009 10.6151
R2965 B.n1012 B.n1011 10.6151
R2966 B.n1013 B.n1012 10.6151
R2967 B.n1014 B.n1013 10.6151
R2968 B.n1016 B.n1014 10.6151
R2969 B.n1017 B.n1016 10.6151
R2970 B.n1018 B.n1017 10.6151
R2971 B.n1019 B.n1018 10.6151
R2972 B.n1021 B.n1019 10.6151
R2973 B.n1022 B.n1021 10.6151
R2974 B.n1023 B.n1022 10.6151
R2975 B.n1024 B.n1023 10.6151
R2976 B.n1026 B.n1024 10.6151
R2977 B.n1027 B.n1026 10.6151
R2978 B.n1028 B.n1027 10.6151
R2979 B.n1029 B.n1028 10.6151
R2980 B.n1031 B.n1029 10.6151
R2981 B.n1032 B.n1031 10.6151
R2982 B.n1033 B.n1032 10.6151
R2983 B.n1034 B.n1033 10.6151
R2984 B.n1036 B.n1034 10.6151
R2985 B.n1037 B.n1036 10.6151
R2986 B.n1038 B.n1037 10.6151
R2987 B.n1039 B.n1038 10.6151
R2988 B.n1041 B.n1039 10.6151
R2989 B.n1042 B.n1041 10.6151
R2990 B.n1043 B.n1042 10.6151
R2991 B.n1044 B.n1043 10.6151
R2992 B.n1046 B.n1044 10.6151
R2993 B.n1047 B.n1046 10.6151
R2994 B.n1048 B.n1047 10.6151
R2995 B.n1049 B.n1048 10.6151
R2996 B.n1051 B.n1049 10.6151
R2997 B.n1052 B.n1051 10.6151
R2998 B.n1053 B.n1052 10.6151
R2999 B.n1054 B.n1053 10.6151
R3000 B.n1056 B.n1054 10.6151
R3001 B.n1057 B.n1056 10.6151
R3002 B.n1058 B.n1057 10.6151
R3003 B.n1059 B.n1058 10.6151
R3004 B.n1061 B.n1059 10.6151
R3005 B.n1062 B.n1061 10.6151
R3006 B.n1063 B.n1062 10.6151
R3007 B.n1064 B.n1063 10.6151
R3008 B.n1066 B.n1064 10.6151
R3009 B.n1067 B.n1066 10.6151
R3010 B.n1068 B.n1067 10.6151
R3011 B.n1069 B.n1068 10.6151
R3012 B.n1071 B.n1069 10.6151
R3013 B.n1072 B.n1071 10.6151
R3014 B.n1073 B.n1072 10.6151
R3015 B.n1074 B.n1073 10.6151
R3016 B.n1076 B.n1074 10.6151
R3017 B.n1077 B.n1076 10.6151
R3018 B.n1078 B.n1077 10.6151
R3019 B.n1079 B.n1078 10.6151
R3020 B.n1081 B.n1079 10.6151
R3021 B.n1082 B.n1081 10.6151
R3022 B.n1083 B.n1082 10.6151
R3023 B.n1084 B.n1083 10.6151
R3024 B.n1086 B.n1084 10.6151
R3025 B.n1087 B.n1086 10.6151
R3026 B.n1088 B.n1087 10.6151
R3027 B.n1089 B.n1088 10.6151
R3028 B.n1090 B.n1089 10.6151
R3029 B.n804 B.n526 10.6151
R3030 B.n799 B.n526 10.6151
R3031 B.n799 B.n798 10.6151
R3032 B.n798 B.n797 10.6151
R3033 B.n797 B.n794 10.6151
R3034 B.n794 B.n793 10.6151
R3035 B.n793 B.n790 10.6151
R3036 B.n790 B.n789 10.6151
R3037 B.n789 B.n786 10.6151
R3038 B.n786 B.n785 10.6151
R3039 B.n785 B.n782 10.6151
R3040 B.n782 B.n781 10.6151
R3041 B.n781 B.n778 10.6151
R3042 B.n778 B.n777 10.6151
R3043 B.n777 B.n774 10.6151
R3044 B.n774 B.n773 10.6151
R3045 B.n773 B.n770 10.6151
R3046 B.n770 B.n769 10.6151
R3047 B.n769 B.n766 10.6151
R3048 B.n766 B.n765 10.6151
R3049 B.n765 B.n762 10.6151
R3050 B.n762 B.n761 10.6151
R3051 B.n761 B.n758 10.6151
R3052 B.n758 B.n757 10.6151
R3053 B.n757 B.n754 10.6151
R3054 B.n754 B.n753 10.6151
R3055 B.n753 B.n750 10.6151
R3056 B.n750 B.n749 10.6151
R3057 B.n749 B.n746 10.6151
R3058 B.n746 B.n745 10.6151
R3059 B.n745 B.n742 10.6151
R3060 B.n742 B.n741 10.6151
R3061 B.n741 B.n738 10.6151
R3062 B.n738 B.n737 10.6151
R3063 B.n737 B.n734 10.6151
R3064 B.n734 B.n733 10.6151
R3065 B.n733 B.n730 10.6151
R3066 B.n730 B.n729 10.6151
R3067 B.n729 B.n726 10.6151
R3068 B.n726 B.n725 10.6151
R3069 B.n725 B.n722 10.6151
R3070 B.n722 B.n721 10.6151
R3071 B.n721 B.n718 10.6151
R3072 B.n718 B.n717 10.6151
R3073 B.n717 B.n714 10.6151
R3074 B.n714 B.n713 10.6151
R3075 B.n713 B.n710 10.6151
R3076 B.n710 B.n709 10.6151
R3077 B.n709 B.n706 10.6151
R3078 B.n704 B.n701 10.6151
R3079 B.n701 B.n700 10.6151
R3080 B.n700 B.n697 10.6151
R3081 B.n697 B.n696 10.6151
R3082 B.n696 B.n693 10.6151
R3083 B.n693 B.n692 10.6151
R3084 B.n692 B.n689 10.6151
R3085 B.n689 B.n688 10.6151
R3086 B.n685 B.n684 10.6151
R3087 B.n684 B.n681 10.6151
R3088 B.n681 B.n680 10.6151
R3089 B.n680 B.n677 10.6151
R3090 B.n677 B.n676 10.6151
R3091 B.n676 B.n673 10.6151
R3092 B.n673 B.n672 10.6151
R3093 B.n672 B.n669 10.6151
R3094 B.n669 B.n668 10.6151
R3095 B.n668 B.n665 10.6151
R3096 B.n665 B.n664 10.6151
R3097 B.n664 B.n661 10.6151
R3098 B.n661 B.n660 10.6151
R3099 B.n660 B.n657 10.6151
R3100 B.n657 B.n656 10.6151
R3101 B.n656 B.n653 10.6151
R3102 B.n653 B.n652 10.6151
R3103 B.n652 B.n649 10.6151
R3104 B.n649 B.n648 10.6151
R3105 B.n648 B.n645 10.6151
R3106 B.n645 B.n644 10.6151
R3107 B.n644 B.n641 10.6151
R3108 B.n641 B.n640 10.6151
R3109 B.n640 B.n637 10.6151
R3110 B.n637 B.n636 10.6151
R3111 B.n636 B.n633 10.6151
R3112 B.n633 B.n632 10.6151
R3113 B.n632 B.n629 10.6151
R3114 B.n629 B.n628 10.6151
R3115 B.n628 B.n625 10.6151
R3116 B.n625 B.n624 10.6151
R3117 B.n624 B.n621 10.6151
R3118 B.n621 B.n620 10.6151
R3119 B.n620 B.n617 10.6151
R3120 B.n617 B.n616 10.6151
R3121 B.n616 B.n613 10.6151
R3122 B.n613 B.n612 10.6151
R3123 B.n612 B.n609 10.6151
R3124 B.n609 B.n608 10.6151
R3125 B.n608 B.n605 10.6151
R3126 B.n605 B.n604 10.6151
R3127 B.n604 B.n601 10.6151
R3128 B.n601 B.n600 10.6151
R3129 B.n600 B.n597 10.6151
R3130 B.n597 B.n596 10.6151
R3131 B.n596 B.n593 10.6151
R3132 B.n593 B.n592 10.6151
R3133 B.n592 B.n589 10.6151
R3134 B.n589 B.n588 10.6151
R3135 B.n806 B.n805 10.6151
R3136 B.n806 B.n518 10.6151
R3137 B.n816 B.n518 10.6151
R3138 B.n817 B.n816 10.6151
R3139 B.n818 B.n817 10.6151
R3140 B.n818 B.n510 10.6151
R3141 B.n828 B.n510 10.6151
R3142 B.n829 B.n828 10.6151
R3143 B.n830 B.n829 10.6151
R3144 B.n830 B.n502 10.6151
R3145 B.n840 B.n502 10.6151
R3146 B.n841 B.n840 10.6151
R3147 B.n842 B.n841 10.6151
R3148 B.n842 B.n494 10.6151
R3149 B.n852 B.n494 10.6151
R3150 B.n853 B.n852 10.6151
R3151 B.n854 B.n853 10.6151
R3152 B.n854 B.n486 10.6151
R3153 B.n864 B.n486 10.6151
R3154 B.n865 B.n864 10.6151
R3155 B.n866 B.n865 10.6151
R3156 B.n866 B.n478 10.6151
R3157 B.n877 B.n478 10.6151
R3158 B.n878 B.n877 10.6151
R3159 B.n879 B.n878 10.6151
R3160 B.n879 B.n471 10.6151
R3161 B.n889 B.n471 10.6151
R3162 B.n890 B.n889 10.6151
R3163 B.n891 B.n890 10.6151
R3164 B.n891 B.n463 10.6151
R3165 B.n901 B.n463 10.6151
R3166 B.n902 B.n901 10.6151
R3167 B.n903 B.n902 10.6151
R3168 B.n903 B.n455 10.6151
R3169 B.n914 B.n455 10.6151
R3170 B.n915 B.n914 10.6151
R3171 B.n916 B.n915 10.6151
R3172 B.n916 B.n448 10.6151
R3173 B.n926 B.n448 10.6151
R3174 B.n927 B.n926 10.6151
R3175 B.n928 B.n927 10.6151
R3176 B.n928 B.n440 10.6151
R3177 B.n938 B.n440 10.6151
R3178 B.n939 B.n938 10.6151
R3179 B.n940 B.n939 10.6151
R3180 B.n940 B.n432 10.6151
R3181 B.n950 B.n432 10.6151
R3182 B.n951 B.n950 10.6151
R3183 B.n952 B.n951 10.6151
R3184 B.n952 B.n424 10.6151
R3185 B.n962 B.n424 10.6151
R3186 B.n963 B.n962 10.6151
R3187 B.n964 B.n963 10.6151
R3188 B.n964 B.n416 10.6151
R3189 B.n974 B.n416 10.6151
R3190 B.n975 B.n974 10.6151
R3191 B.n976 B.n975 10.6151
R3192 B.n976 B.n408 10.6151
R3193 B.n986 B.n408 10.6151
R3194 B.n987 B.n986 10.6151
R3195 B.n988 B.n987 10.6151
R3196 B.n988 B.n400 10.6151
R3197 B.n999 B.n400 10.6151
R3198 B.n1000 B.n999 10.6151
R3199 B.n1001 B.n1000 10.6151
R3200 B.n1001 B.n0 10.6151
R3201 B.n1226 B.n1 10.6151
R3202 B.n1226 B.n1225 10.6151
R3203 B.n1225 B.n1224 10.6151
R3204 B.n1224 B.n10 10.6151
R3205 B.n1218 B.n10 10.6151
R3206 B.n1218 B.n1217 10.6151
R3207 B.n1217 B.n1216 10.6151
R3208 B.n1216 B.n17 10.6151
R3209 B.n1210 B.n17 10.6151
R3210 B.n1210 B.n1209 10.6151
R3211 B.n1209 B.n1208 10.6151
R3212 B.n1208 B.n24 10.6151
R3213 B.n1202 B.n24 10.6151
R3214 B.n1202 B.n1201 10.6151
R3215 B.n1201 B.n1200 10.6151
R3216 B.n1200 B.n31 10.6151
R3217 B.n1194 B.n31 10.6151
R3218 B.n1194 B.n1193 10.6151
R3219 B.n1193 B.n1192 10.6151
R3220 B.n1192 B.n38 10.6151
R3221 B.n1186 B.n38 10.6151
R3222 B.n1186 B.n1185 10.6151
R3223 B.n1185 B.n1184 10.6151
R3224 B.n1184 B.n45 10.6151
R3225 B.n1178 B.n45 10.6151
R3226 B.n1178 B.n1177 10.6151
R3227 B.n1177 B.n1176 10.6151
R3228 B.n1176 B.n52 10.6151
R3229 B.n1170 B.n52 10.6151
R3230 B.n1170 B.n1169 10.6151
R3231 B.n1169 B.n1168 10.6151
R3232 B.n1168 B.n58 10.6151
R3233 B.n1162 B.n58 10.6151
R3234 B.n1162 B.n1161 10.6151
R3235 B.n1161 B.n1160 10.6151
R3236 B.n1160 B.n66 10.6151
R3237 B.n1154 B.n66 10.6151
R3238 B.n1154 B.n1153 10.6151
R3239 B.n1153 B.n1152 10.6151
R3240 B.n1152 B.n73 10.6151
R3241 B.n1146 B.n73 10.6151
R3242 B.n1146 B.n1145 10.6151
R3243 B.n1145 B.n1144 10.6151
R3244 B.n1144 B.n79 10.6151
R3245 B.n1138 B.n79 10.6151
R3246 B.n1138 B.n1137 10.6151
R3247 B.n1137 B.n1136 10.6151
R3248 B.n1136 B.n87 10.6151
R3249 B.n1130 B.n87 10.6151
R3250 B.n1130 B.n1129 10.6151
R3251 B.n1129 B.n1128 10.6151
R3252 B.n1128 B.n94 10.6151
R3253 B.n1122 B.n94 10.6151
R3254 B.n1122 B.n1121 10.6151
R3255 B.n1121 B.n1120 10.6151
R3256 B.n1120 B.n101 10.6151
R3257 B.n1114 B.n101 10.6151
R3258 B.n1114 B.n1113 10.6151
R3259 B.n1113 B.n1112 10.6151
R3260 B.n1112 B.n108 10.6151
R3261 B.n1106 B.n108 10.6151
R3262 B.n1106 B.n1105 10.6151
R3263 B.n1105 B.n1104 10.6151
R3264 B.n1104 B.n115 10.6151
R3265 B.n1098 B.n115 10.6151
R3266 B.n1098 B.n1097 10.6151
R3267 B.t0 B.n430 7.69858
R3268 B.t3 B.n36 7.69858
R3269 B.n281 B.n183 6.5566
R3270 B.n298 B.n297 6.5566
R3271 B.n705 B.n704 6.5566
R3272 B.n688 B.n586 6.5566
R3273 B.n278 B.n183 4.05904
R3274 B.n299 B.n298 4.05904
R3275 B.n706 B.n705 4.05904
R3276 B.n685 B.n586 4.05904
R3277 B.n1232 B.n0 2.81026
R3278 B.n1232 B.n1 2.81026
R3279 B.n911 B.t6 2.19995
R3280 B.n60 B.t4 2.19995
R3281 VN.n67 VN.n35 161.3
R3282 VN.n66 VN.n65 161.3
R3283 VN.n64 VN.n36 161.3
R3284 VN.n63 VN.n62 161.3
R3285 VN.n61 VN.n37 161.3
R3286 VN.n60 VN.n59 161.3
R3287 VN.n58 VN.n38 161.3
R3288 VN.n57 VN.n56 161.3
R3289 VN.n54 VN.n39 161.3
R3290 VN.n53 VN.n52 161.3
R3291 VN.n51 VN.n40 161.3
R3292 VN.n50 VN.n49 161.3
R3293 VN.n48 VN.n41 161.3
R3294 VN.n47 VN.n46 161.3
R3295 VN.n45 VN.n42 161.3
R3296 VN.n32 VN.n0 161.3
R3297 VN.n31 VN.n30 161.3
R3298 VN.n29 VN.n1 161.3
R3299 VN.n28 VN.n27 161.3
R3300 VN.n26 VN.n2 161.3
R3301 VN.n25 VN.n24 161.3
R3302 VN.n23 VN.n3 161.3
R3303 VN.n22 VN.n21 161.3
R3304 VN.n19 VN.n4 161.3
R3305 VN.n18 VN.n17 161.3
R3306 VN.n16 VN.n5 161.3
R3307 VN.n15 VN.n14 161.3
R3308 VN.n13 VN.n6 161.3
R3309 VN.n12 VN.n11 161.3
R3310 VN.n10 VN.n7 161.3
R3311 VN.n9 VN.t5 129.172
R3312 VN.n44 VN.t6 129.172
R3313 VN.n8 VN.t4 96.9931
R3314 VN.n20 VN.t3 96.9931
R3315 VN.n33 VN.t0 96.9931
R3316 VN.n43 VN.t7 96.9931
R3317 VN.n55 VN.t1 96.9931
R3318 VN.n68 VN.t2 96.9931
R3319 VN.n34 VN.n33 58.4488
R3320 VN.n69 VN.n68 58.4488
R3321 VN VN.n69 58.1784
R3322 VN.n9 VN.n8 50.7162
R3323 VN.n44 VN.n43 50.7162
R3324 VN.n27 VN.n26 41.4647
R3325 VN.n62 VN.n61 41.4647
R3326 VN.n14 VN.n13 40.4934
R3327 VN.n14 VN.n5 40.4934
R3328 VN.n49 VN.n48 40.4934
R3329 VN.n49 VN.n40 40.4934
R3330 VN.n27 VN.n1 39.5221
R3331 VN.n62 VN.n36 39.5221
R3332 VN.n12 VN.n7 24.4675
R3333 VN.n13 VN.n12 24.4675
R3334 VN.n18 VN.n5 24.4675
R3335 VN.n19 VN.n18 24.4675
R3336 VN.n21 VN.n3 24.4675
R3337 VN.n25 VN.n3 24.4675
R3338 VN.n26 VN.n25 24.4675
R3339 VN.n31 VN.n1 24.4675
R3340 VN.n32 VN.n31 24.4675
R3341 VN.n48 VN.n47 24.4675
R3342 VN.n47 VN.n42 24.4675
R3343 VN.n61 VN.n60 24.4675
R3344 VN.n60 VN.n38 24.4675
R3345 VN.n56 VN.n38 24.4675
R3346 VN.n54 VN.n53 24.4675
R3347 VN.n53 VN.n40 24.4675
R3348 VN.n67 VN.n66 24.4675
R3349 VN.n66 VN.n36 24.4675
R3350 VN.n8 VN.n7 24.2228
R3351 VN.n20 VN.n19 24.2228
R3352 VN.n43 VN.n42 24.2228
R3353 VN.n55 VN.n54 24.2228
R3354 VN.n33 VN.n32 23.7335
R3355 VN.n68 VN.n67 23.7335
R3356 VN.n45 VN.n44 2.55164
R3357 VN.n10 VN.n9 2.55164
R3358 VN.n69 VN.n35 0.417535
R3359 VN.n34 VN.n0 0.417535
R3360 VN VN.n34 0.394291
R3361 VN.n21 VN.n20 0.24517
R3362 VN.n56 VN.n55 0.24517
R3363 VN.n65 VN.n35 0.189894
R3364 VN.n65 VN.n64 0.189894
R3365 VN.n64 VN.n63 0.189894
R3366 VN.n63 VN.n37 0.189894
R3367 VN.n59 VN.n37 0.189894
R3368 VN.n59 VN.n58 0.189894
R3369 VN.n58 VN.n57 0.189894
R3370 VN.n57 VN.n39 0.189894
R3371 VN.n52 VN.n39 0.189894
R3372 VN.n52 VN.n51 0.189894
R3373 VN.n51 VN.n50 0.189894
R3374 VN.n50 VN.n41 0.189894
R3375 VN.n46 VN.n41 0.189894
R3376 VN.n46 VN.n45 0.189894
R3377 VN.n11 VN.n10 0.189894
R3378 VN.n11 VN.n6 0.189894
R3379 VN.n15 VN.n6 0.189894
R3380 VN.n16 VN.n15 0.189894
R3381 VN.n17 VN.n16 0.189894
R3382 VN.n17 VN.n4 0.189894
R3383 VN.n22 VN.n4 0.189894
R3384 VN.n23 VN.n22 0.189894
R3385 VN.n24 VN.n23 0.189894
R3386 VN.n24 VN.n2 0.189894
R3387 VN.n28 VN.n2 0.189894
R3388 VN.n29 VN.n28 0.189894
R3389 VN.n30 VN.n29 0.189894
R3390 VN.n30 VN.n0 0.189894
R3391 VDD2.n2 VDD2.n1 64.3309
R3392 VDD2.n2 VDD2.n0 64.3309
R3393 VDD2 VDD2.n5 64.328
R3394 VDD2.n4 VDD2.n3 62.6665
R3395 VDD2.n4 VDD2.n2 51.892
R3396 VDD2 VDD2.n4 1.77852
R3397 VDD2.n5 VDD2.t0 1.3447
R3398 VDD2.n5 VDD2.t1 1.3447
R3399 VDD2.n3 VDD2.t5 1.3447
R3400 VDD2.n3 VDD2.t6 1.3447
R3401 VDD2.n1 VDD2.t4 1.3447
R3402 VDD2.n1 VDD2.t7 1.3447
R3403 VDD2.n0 VDD2.t2 1.3447
R3404 VDD2.n0 VDD2.t3 1.3447
C0 VP VDD1 11.6832f
C1 VN VTAIL 11.822701f
C2 VN VDD1 0.153221f
C3 VP VN 9.47022f
C4 VTAIL VDD2 9.352281f
C5 VDD1 VDD2 2.32426f
C6 VP VDD2 0.632043f
C7 VN VDD2 11.2063f
C8 VTAIL VDD1 9.29076f
C9 VP VTAIL 11.8368f
C10 VDD2 B 6.653831f
C11 VDD1 B 7.204293f
C12 VTAIL B 12.844375f
C13 VN B 19.83506f
C14 VP B 18.469343f
C15 VDD2.t2 B 0.311992f
C16 VDD2.t3 B 0.311992f
C17 VDD2.n0 B 2.83705f
C18 VDD2.t4 B 0.311992f
C19 VDD2.t7 B 0.311992f
C20 VDD2.n1 B 2.83705f
C21 VDD2.n2 B 4.34999f
C22 VDD2.t5 B 0.311992f
C23 VDD2.t6 B 0.311992f
C24 VDD2.n3 B 2.81975f
C25 VDD2.n4 B 3.77491f
C26 VDD2.t0 B 0.311992f
C27 VDD2.t1 B 0.311992f
C28 VDD2.n5 B 2.83701f
C29 VN.n0 B 0.032325f
C30 VN.t0 B 2.53766f
C31 VN.n1 B 0.034316f
C32 VN.n2 B 0.017185f
C33 VN.n3 B 0.032029f
C34 VN.n4 B 0.017185f
C35 VN.t3 B 2.53766f
C36 VN.n5 B 0.034155f
C37 VN.n6 B 0.017185f
C38 VN.n7 B 0.03187f
C39 VN.t5 B 2.79045f
C40 VN.t4 B 2.53766f
C41 VN.n8 B 0.951125f
C42 VN.n9 B 0.907144f
C43 VN.n10 B 0.219399f
C44 VN.n11 B 0.017185f
C45 VN.n12 B 0.032029f
C46 VN.n13 B 0.034155f
C47 VN.n14 B 0.013892f
C48 VN.n15 B 0.017185f
C49 VN.n16 B 0.017185f
C50 VN.n17 B 0.017185f
C51 VN.n18 B 0.032029f
C52 VN.n19 B 0.03187f
C53 VN.n20 B 0.881284f
C54 VN.n21 B 0.016373f
C55 VN.n22 B 0.017185f
C56 VN.n23 B 0.017185f
C57 VN.n24 B 0.017185f
C58 VN.n25 B 0.032029f
C59 VN.n26 B 0.033972f
C60 VN.n27 B 0.013915f
C61 VN.n28 B 0.017185f
C62 VN.n29 B 0.017185f
C63 VN.n30 B 0.017185f
C64 VN.n31 B 0.032029f
C65 VN.n32 B 0.031553f
C66 VN.n33 B 0.956328f
C67 VN.n34 B 0.049048f
C68 VN.n35 B 0.032325f
C69 VN.t2 B 2.53766f
C70 VN.n36 B 0.034316f
C71 VN.n37 B 0.017185f
C72 VN.n38 B 0.032029f
C73 VN.n39 B 0.017185f
C74 VN.t1 B 2.53766f
C75 VN.n40 B 0.034155f
C76 VN.n41 B 0.017185f
C77 VN.n42 B 0.03187f
C78 VN.t6 B 2.79045f
C79 VN.t7 B 2.53766f
C80 VN.n43 B 0.951125f
C81 VN.n44 B 0.907144f
C82 VN.n45 B 0.219399f
C83 VN.n46 B 0.017185f
C84 VN.n47 B 0.032029f
C85 VN.n48 B 0.034155f
C86 VN.n49 B 0.013892f
C87 VN.n50 B 0.017185f
C88 VN.n51 B 0.017185f
C89 VN.n52 B 0.017185f
C90 VN.n53 B 0.032029f
C91 VN.n54 B 0.03187f
C92 VN.n55 B 0.881284f
C93 VN.n56 B 0.016373f
C94 VN.n57 B 0.017185f
C95 VN.n58 B 0.017185f
C96 VN.n59 B 0.017185f
C97 VN.n60 B 0.032029f
C98 VN.n61 B 0.033972f
C99 VN.n62 B 0.013915f
C100 VN.n63 B 0.017185f
C101 VN.n64 B 0.017185f
C102 VN.n65 B 0.017185f
C103 VN.n66 B 0.032029f
C104 VN.n67 B 0.031553f
C105 VN.n68 B 0.956328f
C106 VN.n69 B 1.22597f
C107 VTAIL.t3 B 0.2305f
C108 VTAIL.t4 B 0.2305f
C109 VTAIL.n0 B 2.02642f
C110 VTAIL.n1 B 0.413486f
C111 VTAIL.n2 B 0.026364f
C112 VTAIL.n3 B 0.019802f
C113 VTAIL.n4 B 0.010641f
C114 VTAIL.n5 B 0.025151f
C115 VTAIL.n6 B 0.011267f
C116 VTAIL.n7 B 0.019802f
C117 VTAIL.n8 B 0.010641f
C118 VTAIL.n9 B 0.025151f
C119 VTAIL.n10 B 0.011267f
C120 VTAIL.n11 B 0.019802f
C121 VTAIL.n12 B 0.010641f
C122 VTAIL.n13 B 0.025151f
C123 VTAIL.n14 B 0.011267f
C124 VTAIL.n15 B 0.019802f
C125 VTAIL.n16 B 0.010641f
C126 VTAIL.n17 B 0.025151f
C127 VTAIL.n18 B 0.011267f
C128 VTAIL.n19 B 0.019802f
C129 VTAIL.n20 B 0.010641f
C130 VTAIL.n21 B 0.025151f
C131 VTAIL.n22 B 0.011267f
C132 VTAIL.n23 B 0.019802f
C133 VTAIL.n24 B 0.010641f
C134 VTAIL.n25 B 0.025151f
C135 VTAIL.n26 B 0.011267f
C136 VTAIL.n27 B 0.127814f
C137 VTAIL.t1 B 0.041453f
C138 VTAIL.n28 B 0.018863f
C139 VTAIL.n29 B 0.014858f
C140 VTAIL.n30 B 0.010641f
C141 VTAIL.n31 B 1.26386f
C142 VTAIL.n32 B 0.019802f
C143 VTAIL.n33 B 0.010641f
C144 VTAIL.n34 B 0.011267f
C145 VTAIL.n35 B 0.025151f
C146 VTAIL.n36 B 0.025151f
C147 VTAIL.n37 B 0.011267f
C148 VTAIL.n38 B 0.010641f
C149 VTAIL.n39 B 0.019802f
C150 VTAIL.n40 B 0.019802f
C151 VTAIL.n41 B 0.010641f
C152 VTAIL.n42 B 0.011267f
C153 VTAIL.n43 B 0.025151f
C154 VTAIL.n44 B 0.025151f
C155 VTAIL.n45 B 0.011267f
C156 VTAIL.n46 B 0.010641f
C157 VTAIL.n47 B 0.019802f
C158 VTAIL.n48 B 0.019802f
C159 VTAIL.n49 B 0.010641f
C160 VTAIL.n50 B 0.011267f
C161 VTAIL.n51 B 0.025151f
C162 VTAIL.n52 B 0.025151f
C163 VTAIL.n53 B 0.011267f
C164 VTAIL.n54 B 0.010641f
C165 VTAIL.n55 B 0.019802f
C166 VTAIL.n56 B 0.019802f
C167 VTAIL.n57 B 0.010641f
C168 VTAIL.n58 B 0.011267f
C169 VTAIL.n59 B 0.025151f
C170 VTAIL.n60 B 0.025151f
C171 VTAIL.n61 B 0.011267f
C172 VTAIL.n62 B 0.010641f
C173 VTAIL.n63 B 0.019802f
C174 VTAIL.n64 B 0.019802f
C175 VTAIL.n65 B 0.010641f
C176 VTAIL.n66 B 0.011267f
C177 VTAIL.n67 B 0.025151f
C178 VTAIL.n68 B 0.025151f
C179 VTAIL.n69 B 0.025151f
C180 VTAIL.n70 B 0.011267f
C181 VTAIL.n71 B 0.010641f
C182 VTAIL.n72 B 0.019802f
C183 VTAIL.n73 B 0.019802f
C184 VTAIL.n74 B 0.010641f
C185 VTAIL.n75 B 0.010954f
C186 VTAIL.n76 B 0.010954f
C187 VTAIL.n77 B 0.025151f
C188 VTAIL.n78 B 0.051849f
C189 VTAIL.n79 B 0.011267f
C190 VTAIL.n80 B 0.010641f
C191 VTAIL.n81 B 0.048207f
C192 VTAIL.n82 B 0.028818f
C193 VTAIL.n83 B 0.267742f
C194 VTAIL.n84 B 0.026364f
C195 VTAIL.n85 B 0.019802f
C196 VTAIL.n86 B 0.010641f
C197 VTAIL.n87 B 0.025151f
C198 VTAIL.n88 B 0.011267f
C199 VTAIL.n89 B 0.019802f
C200 VTAIL.n90 B 0.010641f
C201 VTAIL.n91 B 0.025151f
C202 VTAIL.n92 B 0.011267f
C203 VTAIL.n93 B 0.019802f
C204 VTAIL.n94 B 0.010641f
C205 VTAIL.n95 B 0.025151f
C206 VTAIL.n96 B 0.011267f
C207 VTAIL.n97 B 0.019802f
C208 VTAIL.n98 B 0.010641f
C209 VTAIL.n99 B 0.025151f
C210 VTAIL.n100 B 0.011267f
C211 VTAIL.n101 B 0.019802f
C212 VTAIL.n102 B 0.010641f
C213 VTAIL.n103 B 0.025151f
C214 VTAIL.n104 B 0.011267f
C215 VTAIL.n105 B 0.019802f
C216 VTAIL.n106 B 0.010641f
C217 VTAIL.n107 B 0.025151f
C218 VTAIL.n108 B 0.011267f
C219 VTAIL.n109 B 0.127814f
C220 VTAIL.t9 B 0.041453f
C221 VTAIL.n110 B 0.018863f
C222 VTAIL.n111 B 0.014858f
C223 VTAIL.n112 B 0.010641f
C224 VTAIL.n113 B 1.26386f
C225 VTAIL.n114 B 0.019802f
C226 VTAIL.n115 B 0.010641f
C227 VTAIL.n116 B 0.011267f
C228 VTAIL.n117 B 0.025151f
C229 VTAIL.n118 B 0.025151f
C230 VTAIL.n119 B 0.011267f
C231 VTAIL.n120 B 0.010641f
C232 VTAIL.n121 B 0.019802f
C233 VTAIL.n122 B 0.019802f
C234 VTAIL.n123 B 0.010641f
C235 VTAIL.n124 B 0.011267f
C236 VTAIL.n125 B 0.025151f
C237 VTAIL.n126 B 0.025151f
C238 VTAIL.n127 B 0.011267f
C239 VTAIL.n128 B 0.010641f
C240 VTAIL.n129 B 0.019802f
C241 VTAIL.n130 B 0.019802f
C242 VTAIL.n131 B 0.010641f
C243 VTAIL.n132 B 0.011267f
C244 VTAIL.n133 B 0.025151f
C245 VTAIL.n134 B 0.025151f
C246 VTAIL.n135 B 0.011267f
C247 VTAIL.n136 B 0.010641f
C248 VTAIL.n137 B 0.019802f
C249 VTAIL.n138 B 0.019802f
C250 VTAIL.n139 B 0.010641f
C251 VTAIL.n140 B 0.011267f
C252 VTAIL.n141 B 0.025151f
C253 VTAIL.n142 B 0.025151f
C254 VTAIL.n143 B 0.011267f
C255 VTAIL.n144 B 0.010641f
C256 VTAIL.n145 B 0.019802f
C257 VTAIL.n146 B 0.019802f
C258 VTAIL.n147 B 0.010641f
C259 VTAIL.n148 B 0.011267f
C260 VTAIL.n149 B 0.025151f
C261 VTAIL.n150 B 0.025151f
C262 VTAIL.n151 B 0.025151f
C263 VTAIL.n152 B 0.011267f
C264 VTAIL.n153 B 0.010641f
C265 VTAIL.n154 B 0.019802f
C266 VTAIL.n155 B 0.019802f
C267 VTAIL.n156 B 0.010641f
C268 VTAIL.n157 B 0.010954f
C269 VTAIL.n158 B 0.010954f
C270 VTAIL.n159 B 0.025151f
C271 VTAIL.n160 B 0.051849f
C272 VTAIL.n161 B 0.011267f
C273 VTAIL.n162 B 0.010641f
C274 VTAIL.n163 B 0.048207f
C275 VTAIL.n164 B 0.028818f
C276 VTAIL.n165 B 0.267742f
C277 VTAIL.t14 B 0.2305f
C278 VTAIL.t13 B 0.2305f
C279 VTAIL.n166 B 2.02642f
C280 VTAIL.n167 B 0.629248f
C281 VTAIL.n168 B 0.026364f
C282 VTAIL.n169 B 0.019802f
C283 VTAIL.n170 B 0.010641f
C284 VTAIL.n171 B 0.025151f
C285 VTAIL.n172 B 0.011267f
C286 VTAIL.n173 B 0.019802f
C287 VTAIL.n174 B 0.010641f
C288 VTAIL.n175 B 0.025151f
C289 VTAIL.n176 B 0.011267f
C290 VTAIL.n177 B 0.019802f
C291 VTAIL.n178 B 0.010641f
C292 VTAIL.n179 B 0.025151f
C293 VTAIL.n180 B 0.011267f
C294 VTAIL.n181 B 0.019802f
C295 VTAIL.n182 B 0.010641f
C296 VTAIL.n183 B 0.025151f
C297 VTAIL.n184 B 0.011267f
C298 VTAIL.n185 B 0.019802f
C299 VTAIL.n186 B 0.010641f
C300 VTAIL.n187 B 0.025151f
C301 VTAIL.n188 B 0.011267f
C302 VTAIL.n189 B 0.019802f
C303 VTAIL.n190 B 0.010641f
C304 VTAIL.n191 B 0.025151f
C305 VTAIL.n192 B 0.011267f
C306 VTAIL.n193 B 0.127814f
C307 VTAIL.t8 B 0.041453f
C308 VTAIL.n194 B 0.018863f
C309 VTAIL.n195 B 0.014858f
C310 VTAIL.n196 B 0.010641f
C311 VTAIL.n197 B 1.26386f
C312 VTAIL.n198 B 0.019802f
C313 VTAIL.n199 B 0.010641f
C314 VTAIL.n200 B 0.011267f
C315 VTAIL.n201 B 0.025151f
C316 VTAIL.n202 B 0.025151f
C317 VTAIL.n203 B 0.011267f
C318 VTAIL.n204 B 0.010641f
C319 VTAIL.n205 B 0.019802f
C320 VTAIL.n206 B 0.019802f
C321 VTAIL.n207 B 0.010641f
C322 VTAIL.n208 B 0.011267f
C323 VTAIL.n209 B 0.025151f
C324 VTAIL.n210 B 0.025151f
C325 VTAIL.n211 B 0.011267f
C326 VTAIL.n212 B 0.010641f
C327 VTAIL.n213 B 0.019802f
C328 VTAIL.n214 B 0.019802f
C329 VTAIL.n215 B 0.010641f
C330 VTAIL.n216 B 0.011267f
C331 VTAIL.n217 B 0.025151f
C332 VTAIL.n218 B 0.025151f
C333 VTAIL.n219 B 0.011267f
C334 VTAIL.n220 B 0.010641f
C335 VTAIL.n221 B 0.019802f
C336 VTAIL.n222 B 0.019802f
C337 VTAIL.n223 B 0.010641f
C338 VTAIL.n224 B 0.011267f
C339 VTAIL.n225 B 0.025151f
C340 VTAIL.n226 B 0.025151f
C341 VTAIL.n227 B 0.011267f
C342 VTAIL.n228 B 0.010641f
C343 VTAIL.n229 B 0.019802f
C344 VTAIL.n230 B 0.019802f
C345 VTAIL.n231 B 0.010641f
C346 VTAIL.n232 B 0.011267f
C347 VTAIL.n233 B 0.025151f
C348 VTAIL.n234 B 0.025151f
C349 VTAIL.n235 B 0.025151f
C350 VTAIL.n236 B 0.011267f
C351 VTAIL.n237 B 0.010641f
C352 VTAIL.n238 B 0.019802f
C353 VTAIL.n239 B 0.019802f
C354 VTAIL.n240 B 0.010641f
C355 VTAIL.n241 B 0.010954f
C356 VTAIL.n242 B 0.010954f
C357 VTAIL.n243 B 0.025151f
C358 VTAIL.n244 B 0.051849f
C359 VTAIL.n245 B 0.011267f
C360 VTAIL.n246 B 0.010641f
C361 VTAIL.n247 B 0.048207f
C362 VTAIL.n248 B 0.028818f
C363 VTAIL.n249 B 1.53647f
C364 VTAIL.n250 B 0.026364f
C365 VTAIL.n251 B 0.019802f
C366 VTAIL.n252 B 0.010641f
C367 VTAIL.n253 B 0.025151f
C368 VTAIL.n254 B 0.011267f
C369 VTAIL.n255 B 0.019802f
C370 VTAIL.n256 B 0.010641f
C371 VTAIL.n257 B 0.025151f
C372 VTAIL.n258 B 0.025151f
C373 VTAIL.n259 B 0.011267f
C374 VTAIL.n260 B 0.019802f
C375 VTAIL.n261 B 0.010641f
C376 VTAIL.n262 B 0.025151f
C377 VTAIL.n263 B 0.011267f
C378 VTAIL.n264 B 0.019802f
C379 VTAIL.n265 B 0.010641f
C380 VTAIL.n266 B 0.025151f
C381 VTAIL.n267 B 0.011267f
C382 VTAIL.n268 B 0.019802f
C383 VTAIL.n269 B 0.010641f
C384 VTAIL.n270 B 0.025151f
C385 VTAIL.n271 B 0.011267f
C386 VTAIL.n272 B 0.019802f
C387 VTAIL.n273 B 0.010641f
C388 VTAIL.n274 B 0.025151f
C389 VTAIL.n275 B 0.011267f
C390 VTAIL.n276 B 0.127814f
C391 VTAIL.t7 B 0.041453f
C392 VTAIL.n277 B 0.018863f
C393 VTAIL.n278 B 0.014858f
C394 VTAIL.n279 B 0.010641f
C395 VTAIL.n280 B 1.26386f
C396 VTAIL.n281 B 0.019802f
C397 VTAIL.n282 B 0.010641f
C398 VTAIL.n283 B 0.011267f
C399 VTAIL.n284 B 0.025151f
C400 VTAIL.n285 B 0.025151f
C401 VTAIL.n286 B 0.011267f
C402 VTAIL.n287 B 0.010641f
C403 VTAIL.n288 B 0.019802f
C404 VTAIL.n289 B 0.019802f
C405 VTAIL.n290 B 0.010641f
C406 VTAIL.n291 B 0.011267f
C407 VTAIL.n292 B 0.025151f
C408 VTAIL.n293 B 0.025151f
C409 VTAIL.n294 B 0.011267f
C410 VTAIL.n295 B 0.010641f
C411 VTAIL.n296 B 0.019802f
C412 VTAIL.n297 B 0.019802f
C413 VTAIL.n298 B 0.010641f
C414 VTAIL.n299 B 0.011267f
C415 VTAIL.n300 B 0.025151f
C416 VTAIL.n301 B 0.025151f
C417 VTAIL.n302 B 0.011267f
C418 VTAIL.n303 B 0.010641f
C419 VTAIL.n304 B 0.019802f
C420 VTAIL.n305 B 0.019802f
C421 VTAIL.n306 B 0.010641f
C422 VTAIL.n307 B 0.011267f
C423 VTAIL.n308 B 0.025151f
C424 VTAIL.n309 B 0.025151f
C425 VTAIL.n310 B 0.011267f
C426 VTAIL.n311 B 0.010641f
C427 VTAIL.n312 B 0.019802f
C428 VTAIL.n313 B 0.019802f
C429 VTAIL.n314 B 0.010641f
C430 VTAIL.n315 B 0.011267f
C431 VTAIL.n316 B 0.025151f
C432 VTAIL.n317 B 0.025151f
C433 VTAIL.n318 B 0.011267f
C434 VTAIL.n319 B 0.010641f
C435 VTAIL.n320 B 0.019802f
C436 VTAIL.n321 B 0.019802f
C437 VTAIL.n322 B 0.010641f
C438 VTAIL.n323 B 0.010954f
C439 VTAIL.n324 B 0.010954f
C440 VTAIL.n325 B 0.025151f
C441 VTAIL.n326 B 0.051849f
C442 VTAIL.n327 B 0.011267f
C443 VTAIL.n328 B 0.010641f
C444 VTAIL.n329 B 0.048207f
C445 VTAIL.n330 B 0.028818f
C446 VTAIL.n331 B 1.53647f
C447 VTAIL.t6 B 0.2305f
C448 VTAIL.t0 B 0.2305f
C449 VTAIL.n332 B 2.02643f
C450 VTAIL.n333 B 0.629238f
C451 VTAIL.n334 B 0.026364f
C452 VTAIL.n335 B 0.019802f
C453 VTAIL.n336 B 0.010641f
C454 VTAIL.n337 B 0.025151f
C455 VTAIL.n338 B 0.011267f
C456 VTAIL.n339 B 0.019802f
C457 VTAIL.n340 B 0.010641f
C458 VTAIL.n341 B 0.025151f
C459 VTAIL.n342 B 0.025151f
C460 VTAIL.n343 B 0.011267f
C461 VTAIL.n344 B 0.019802f
C462 VTAIL.n345 B 0.010641f
C463 VTAIL.n346 B 0.025151f
C464 VTAIL.n347 B 0.011267f
C465 VTAIL.n348 B 0.019802f
C466 VTAIL.n349 B 0.010641f
C467 VTAIL.n350 B 0.025151f
C468 VTAIL.n351 B 0.011267f
C469 VTAIL.n352 B 0.019802f
C470 VTAIL.n353 B 0.010641f
C471 VTAIL.n354 B 0.025151f
C472 VTAIL.n355 B 0.011267f
C473 VTAIL.n356 B 0.019802f
C474 VTAIL.n357 B 0.010641f
C475 VTAIL.n358 B 0.025151f
C476 VTAIL.n359 B 0.011267f
C477 VTAIL.n360 B 0.127814f
C478 VTAIL.t5 B 0.041453f
C479 VTAIL.n361 B 0.018863f
C480 VTAIL.n362 B 0.014858f
C481 VTAIL.n363 B 0.010641f
C482 VTAIL.n364 B 1.26386f
C483 VTAIL.n365 B 0.019802f
C484 VTAIL.n366 B 0.010641f
C485 VTAIL.n367 B 0.011267f
C486 VTAIL.n368 B 0.025151f
C487 VTAIL.n369 B 0.025151f
C488 VTAIL.n370 B 0.011267f
C489 VTAIL.n371 B 0.010641f
C490 VTAIL.n372 B 0.019802f
C491 VTAIL.n373 B 0.019802f
C492 VTAIL.n374 B 0.010641f
C493 VTAIL.n375 B 0.011267f
C494 VTAIL.n376 B 0.025151f
C495 VTAIL.n377 B 0.025151f
C496 VTAIL.n378 B 0.011267f
C497 VTAIL.n379 B 0.010641f
C498 VTAIL.n380 B 0.019802f
C499 VTAIL.n381 B 0.019802f
C500 VTAIL.n382 B 0.010641f
C501 VTAIL.n383 B 0.011267f
C502 VTAIL.n384 B 0.025151f
C503 VTAIL.n385 B 0.025151f
C504 VTAIL.n386 B 0.011267f
C505 VTAIL.n387 B 0.010641f
C506 VTAIL.n388 B 0.019802f
C507 VTAIL.n389 B 0.019802f
C508 VTAIL.n390 B 0.010641f
C509 VTAIL.n391 B 0.011267f
C510 VTAIL.n392 B 0.025151f
C511 VTAIL.n393 B 0.025151f
C512 VTAIL.n394 B 0.011267f
C513 VTAIL.n395 B 0.010641f
C514 VTAIL.n396 B 0.019802f
C515 VTAIL.n397 B 0.019802f
C516 VTAIL.n398 B 0.010641f
C517 VTAIL.n399 B 0.011267f
C518 VTAIL.n400 B 0.025151f
C519 VTAIL.n401 B 0.025151f
C520 VTAIL.n402 B 0.011267f
C521 VTAIL.n403 B 0.010641f
C522 VTAIL.n404 B 0.019802f
C523 VTAIL.n405 B 0.019802f
C524 VTAIL.n406 B 0.010641f
C525 VTAIL.n407 B 0.010954f
C526 VTAIL.n408 B 0.010954f
C527 VTAIL.n409 B 0.025151f
C528 VTAIL.n410 B 0.051849f
C529 VTAIL.n411 B 0.011267f
C530 VTAIL.n412 B 0.010641f
C531 VTAIL.n413 B 0.048207f
C532 VTAIL.n414 B 0.028818f
C533 VTAIL.n415 B 0.267742f
C534 VTAIL.n416 B 0.026364f
C535 VTAIL.n417 B 0.019802f
C536 VTAIL.n418 B 0.010641f
C537 VTAIL.n419 B 0.025151f
C538 VTAIL.n420 B 0.011267f
C539 VTAIL.n421 B 0.019802f
C540 VTAIL.n422 B 0.010641f
C541 VTAIL.n423 B 0.025151f
C542 VTAIL.n424 B 0.025151f
C543 VTAIL.n425 B 0.011267f
C544 VTAIL.n426 B 0.019802f
C545 VTAIL.n427 B 0.010641f
C546 VTAIL.n428 B 0.025151f
C547 VTAIL.n429 B 0.011267f
C548 VTAIL.n430 B 0.019802f
C549 VTAIL.n431 B 0.010641f
C550 VTAIL.n432 B 0.025151f
C551 VTAIL.n433 B 0.011267f
C552 VTAIL.n434 B 0.019802f
C553 VTAIL.n435 B 0.010641f
C554 VTAIL.n436 B 0.025151f
C555 VTAIL.n437 B 0.011267f
C556 VTAIL.n438 B 0.019802f
C557 VTAIL.n439 B 0.010641f
C558 VTAIL.n440 B 0.025151f
C559 VTAIL.n441 B 0.011267f
C560 VTAIL.n442 B 0.127814f
C561 VTAIL.t15 B 0.041453f
C562 VTAIL.n443 B 0.018863f
C563 VTAIL.n444 B 0.014858f
C564 VTAIL.n445 B 0.010641f
C565 VTAIL.n446 B 1.26386f
C566 VTAIL.n447 B 0.019802f
C567 VTAIL.n448 B 0.010641f
C568 VTAIL.n449 B 0.011267f
C569 VTAIL.n450 B 0.025151f
C570 VTAIL.n451 B 0.025151f
C571 VTAIL.n452 B 0.011267f
C572 VTAIL.n453 B 0.010641f
C573 VTAIL.n454 B 0.019802f
C574 VTAIL.n455 B 0.019802f
C575 VTAIL.n456 B 0.010641f
C576 VTAIL.n457 B 0.011267f
C577 VTAIL.n458 B 0.025151f
C578 VTAIL.n459 B 0.025151f
C579 VTAIL.n460 B 0.011267f
C580 VTAIL.n461 B 0.010641f
C581 VTAIL.n462 B 0.019802f
C582 VTAIL.n463 B 0.019802f
C583 VTAIL.n464 B 0.010641f
C584 VTAIL.n465 B 0.011267f
C585 VTAIL.n466 B 0.025151f
C586 VTAIL.n467 B 0.025151f
C587 VTAIL.n468 B 0.011267f
C588 VTAIL.n469 B 0.010641f
C589 VTAIL.n470 B 0.019802f
C590 VTAIL.n471 B 0.019802f
C591 VTAIL.n472 B 0.010641f
C592 VTAIL.n473 B 0.011267f
C593 VTAIL.n474 B 0.025151f
C594 VTAIL.n475 B 0.025151f
C595 VTAIL.n476 B 0.011267f
C596 VTAIL.n477 B 0.010641f
C597 VTAIL.n478 B 0.019802f
C598 VTAIL.n479 B 0.019802f
C599 VTAIL.n480 B 0.010641f
C600 VTAIL.n481 B 0.011267f
C601 VTAIL.n482 B 0.025151f
C602 VTAIL.n483 B 0.025151f
C603 VTAIL.n484 B 0.011267f
C604 VTAIL.n485 B 0.010641f
C605 VTAIL.n486 B 0.019802f
C606 VTAIL.n487 B 0.019802f
C607 VTAIL.n488 B 0.010641f
C608 VTAIL.n489 B 0.010954f
C609 VTAIL.n490 B 0.010954f
C610 VTAIL.n491 B 0.025151f
C611 VTAIL.n492 B 0.051849f
C612 VTAIL.n493 B 0.011267f
C613 VTAIL.n494 B 0.010641f
C614 VTAIL.n495 B 0.048207f
C615 VTAIL.n496 B 0.028818f
C616 VTAIL.n497 B 0.267742f
C617 VTAIL.t12 B 0.2305f
C618 VTAIL.t10 B 0.2305f
C619 VTAIL.n498 B 2.02643f
C620 VTAIL.n499 B 0.629238f
C621 VTAIL.n500 B 0.026364f
C622 VTAIL.n501 B 0.019802f
C623 VTAIL.n502 B 0.010641f
C624 VTAIL.n503 B 0.025151f
C625 VTAIL.n504 B 0.011267f
C626 VTAIL.n505 B 0.019802f
C627 VTAIL.n506 B 0.010641f
C628 VTAIL.n507 B 0.025151f
C629 VTAIL.n508 B 0.025151f
C630 VTAIL.n509 B 0.011267f
C631 VTAIL.n510 B 0.019802f
C632 VTAIL.n511 B 0.010641f
C633 VTAIL.n512 B 0.025151f
C634 VTAIL.n513 B 0.011267f
C635 VTAIL.n514 B 0.019802f
C636 VTAIL.n515 B 0.010641f
C637 VTAIL.n516 B 0.025151f
C638 VTAIL.n517 B 0.011267f
C639 VTAIL.n518 B 0.019802f
C640 VTAIL.n519 B 0.010641f
C641 VTAIL.n520 B 0.025151f
C642 VTAIL.n521 B 0.011267f
C643 VTAIL.n522 B 0.019802f
C644 VTAIL.n523 B 0.010641f
C645 VTAIL.n524 B 0.025151f
C646 VTAIL.n525 B 0.011267f
C647 VTAIL.n526 B 0.127814f
C648 VTAIL.t11 B 0.041453f
C649 VTAIL.n527 B 0.018863f
C650 VTAIL.n528 B 0.014858f
C651 VTAIL.n529 B 0.010641f
C652 VTAIL.n530 B 1.26386f
C653 VTAIL.n531 B 0.019802f
C654 VTAIL.n532 B 0.010641f
C655 VTAIL.n533 B 0.011267f
C656 VTAIL.n534 B 0.025151f
C657 VTAIL.n535 B 0.025151f
C658 VTAIL.n536 B 0.011267f
C659 VTAIL.n537 B 0.010641f
C660 VTAIL.n538 B 0.019802f
C661 VTAIL.n539 B 0.019802f
C662 VTAIL.n540 B 0.010641f
C663 VTAIL.n541 B 0.011267f
C664 VTAIL.n542 B 0.025151f
C665 VTAIL.n543 B 0.025151f
C666 VTAIL.n544 B 0.011267f
C667 VTAIL.n545 B 0.010641f
C668 VTAIL.n546 B 0.019802f
C669 VTAIL.n547 B 0.019802f
C670 VTAIL.n548 B 0.010641f
C671 VTAIL.n549 B 0.011267f
C672 VTAIL.n550 B 0.025151f
C673 VTAIL.n551 B 0.025151f
C674 VTAIL.n552 B 0.011267f
C675 VTAIL.n553 B 0.010641f
C676 VTAIL.n554 B 0.019802f
C677 VTAIL.n555 B 0.019802f
C678 VTAIL.n556 B 0.010641f
C679 VTAIL.n557 B 0.011267f
C680 VTAIL.n558 B 0.025151f
C681 VTAIL.n559 B 0.025151f
C682 VTAIL.n560 B 0.011267f
C683 VTAIL.n561 B 0.010641f
C684 VTAIL.n562 B 0.019802f
C685 VTAIL.n563 B 0.019802f
C686 VTAIL.n564 B 0.010641f
C687 VTAIL.n565 B 0.011267f
C688 VTAIL.n566 B 0.025151f
C689 VTAIL.n567 B 0.025151f
C690 VTAIL.n568 B 0.011267f
C691 VTAIL.n569 B 0.010641f
C692 VTAIL.n570 B 0.019802f
C693 VTAIL.n571 B 0.019802f
C694 VTAIL.n572 B 0.010641f
C695 VTAIL.n573 B 0.010954f
C696 VTAIL.n574 B 0.010954f
C697 VTAIL.n575 B 0.025151f
C698 VTAIL.n576 B 0.051849f
C699 VTAIL.n577 B 0.011267f
C700 VTAIL.n578 B 0.010641f
C701 VTAIL.n579 B 0.048207f
C702 VTAIL.n580 B 0.028818f
C703 VTAIL.n581 B 1.53647f
C704 VTAIL.n582 B 0.026364f
C705 VTAIL.n583 B 0.019802f
C706 VTAIL.n584 B 0.010641f
C707 VTAIL.n585 B 0.025151f
C708 VTAIL.n586 B 0.011267f
C709 VTAIL.n587 B 0.019802f
C710 VTAIL.n588 B 0.010641f
C711 VTAIL.n589 B 0.025151f
C712 VTAIL.n590 B 0.011267f
C713 VTAIL.n591 B 0.019802f
C714 VTAIL.n592 B 0.010641f
C715 VTAIL.n593 B 0.025151f
C716 VTAIL.n594 B 0.011267f
C717 VTAIL.n595 B 0.019802f
C718 VTAIL.n596 B 0.010641f
C719 VTAIL.n597 B 0.025151f
C720 VTAIL.n598 B 0.011267f
C721 VTAIL.n599 B 0.019802f
C722 VTAIL.n600 B 0.010641f
C723 VTAIL.n601 B 0.025151f
C724 VTAIL.n602 B 0.011267f
C725 VTAIL.n603 B 0.019802f
C726 VTAIL.n604 B 0.010641f
C727 VTAIL.n605 B 0.025151f
C728 VTAIL.n606 B 0.011267f
C729 VTAIL.n607 B 0.127814f
C730 VTAIL.t2 B 0.041453f
C731 VTAIL.n608 B 0.018863f
C732 VTAIL.n609 B 0.014858f
C733 VTAIL.n610 B 0.010641f
C734 VTAIL.n611 B 1.26386f
C735 VTAIL.n612 B 0.019802f
C736 VTAIL.n613 B 0.010641f
C737 VTAIL.n614 B 0.011267f
C738 VTAIL.n615 B 0.025151f
C739 VTAIL.n616 B 0.025151f
C740 VTAIL.n617 B 0.011267f
C741 VTAIL.n618 B 0.010641f
C742 VTAIL.n619 B 0.019802f
C743 VTAIL.n620 B 0.019802f
C744 VTAIL.n621 B 0.010641f
C745 VTAIL.n622 B 0.011267f
C746 VTAIL.n623 B 0.025151f
C747 VTAIL.n624 B 0.025151f
C748 VTAIL.n625 B 0.011267f
C749 VTAIL.n626 B 0.010641f
C750 VTAIL.n627 B 0.019802f
C751 VTAIL.n628 B 0.019802f
C752 VTAIL.n629 B 0.010641f
C753 VTAIL.n630 B 0.011267f
C754 VTAIL.n631 B 0.025151f
C755 VTAIL.n632 B 0.025151f
C756 VTAIL.n633 B 0.011267f
C757 VTAIL.n634 B 0.010641f
C758 VTAIL.n635 B 0.019802f
C759 VTAIL.n636 B 0.019802f
C760 VTAIL.n637 B 0.010641f
C761 VTAIL.n638 B 0.011267f
C762 VTAIL.n639 B 0.025151f
C763 VTAIL.n640 B 0.025151f
C764 VTAIL.n641 B 0.011267f
C765 VTAIL.n642 B 0.010641f
C766 VTAIL.n643 B 0.019802f
C767 VTAIL.n644 B 0.019802f
C768 VTAIL.n645 B 0.010641f
C769 VTAIL.n646 B 0.011267f
C770 VTAIL.n647 B 0.025151f
C771 VTAIL.n648 B 0.025151f
C772 VTAIL.n649 B 0.025151f
C773 VTAIL.n650 B 0.011267f
C774 VTAIL.n651 B 0.010641f
C775 VTAIL.n652 B 0.019802f
C776 VTAIL.n653 B 0.019802f
C777 VTAIL.n654 B 0.010641f
C778 VTAIL.n655 B 0.010954f
C779 VTAIL.n656 B 0.010954f
C780 VTAIL.n657 B 0.025151f
C781 VTAIL.n658 B 0.051849f
C782 VTAIL.n659 B 0.011267f
C783 VTAIL.n660 B 0.010641f
C784 VTAIL.n661 B 0.048207f
C785 VTAIL.n662 B 0.028818f
C786 VTAIL.n663 B 1.53276f
C787 VDD1.t3 B 0.316076f
C788 VDD1.t4 B 0.316076f
C789 VDD1.n0 B 2.87562f
C790 VDD1.t6 B 0.316076f
C791 VDD1.t2 B 0.316076f
C792 VDD1.n1 B 2.87418f
C793 VDD1.t5 B 0.316076f
C794 VDD1.t7 B 0.316076f
C795 VDD1.n2 B 2.87418f
C796 VDD1.n3 B 4.46278f
C797 VDD1.t0 B 0.316076f
C798 VDD1.t1 B 0.316076f
C799 VDD1.n4 B 2.85665f
C800 VDD1.n5 B 3.85858f
C801 VP.n0 B 0.032847f
C802 VP.t6 B 2.57862f
C803 VP.n1 B 0.03487f
C804 VP.n2 B 0.017462f
C805 VP.n3 B 0.032545f
C806 VP.n4 B 0.017462f
C807 VP.t2 B 2.57862f
C808 VP.n5 B 0.034706f
C809 VP.n6 B 0.017462f
C810 VP.n7 B 0.032384f
C811 VP.n8 B 0.017462f
C812 VP.n9 B 0.03452f
C813 VP.n10 B 0.017462f
C814 VP.n11 B 0.032063f
C815 VP.n12 B 0.032847f
C816 VP.t4 B 2.57862f
C817 VP.n13 B 0.03487f
C818 VP.n14 B 0.017462f
C819 VP.n15 B 0.032545f
C820 VP.n16 B 0.017462f
C821 VP.t5 B 2.57862f
C822 VP.n17 B 0.034706f
C823 VP.n18 B 0.017462f
C824 VP.n19 B 0.032384f
C825 VP.t0 B 2.83548f
C826 VP.t3 B 2.57862f
C827 VP.n20 B 0.966476f
C828 VP.n21 B 0.921788f
C829 VP.n22 B 0.222941f
C830 VP.n23 B 0.017462f
C831 VP.n24 B 0.032545f
C832 VP.n25 B 0.034706f
C833 VP.n26 B 0.014117f
C834 VP.n27 B 0.017462f
C835 VP.n28 B 0.017462f
C836 VP.n29 B 0.017462f
C837 VP.n30 B 0.032545f
C838 VP.n31 B 0.032384f
C839 VP.n32 B 0.895508f
C840 VP.n33 B 0.016638f
C841 VP.n34 B 0.017462f
C842 VP.n35 B 0.017462f
C843 VP.n36 B 0.017462f
C844 VP.n37 B 0.032545f
C845 VP.n38 B 0.03452f
C846 VP.n39 B 0.014139f
C847 VP.n40 B 0.017462f
C848 VP.n41 B 0.017462f
C849 VP.n42 B 0.017462f
C850 VP.n43 B 0.032545f
C851 VP.n44 B 0.032063f
C852 VP.n45 B 0.971763f
C853 VP.n46 B 1.24167f
C854 VP.t7 B 2.57862f
C855 VP.n47 B 0.971763f
C856 VP.n48 B 1.25247f
C857 VP.n49 B 0.032847f
C858 VP.n50 B 0.017462f
C859 VP.n51 B 0.032545f
C860 VP.n52 B 0.03487f
C861 VP.n53 B 0.014139f
C862 VP.n54 B 0.017462f
C863 VP.n55 B 0.017462f
C864 VP.n56 B 0.017462f
C865 VP.n57 B 0.032545f
C866 VP.n58 B 0.032545f
C867 VP.t1 B 2.57862f
C868 VP.n59 B 0.895508f
C869 VP.n60 B 0.016638f
C870 VP.n61 B 0.017462f
C871 VP.n62 B 0.017462f
C872 VP.n63 B 0.017462f
C873 VP.n64 B 0.032545f
C874 VP.n65 B 0.034706f
C875 VP.n66 B 0.014117f
C876 VP.n67 B 0.017462f
C877 VP.n68 B 0.017462f
C878 VP.n69 B 0.017462f
C879 VP.n70 B 0.032545f
C880 VP.n71 B 0.032384f
C881 VP.n72 B 0.895508f
C882 VP.n73 B 0.016638f
C883 VP.n74 B 0.017462f
C884 VP.n75 B 0.017462f
C885 VP.n76 B 0.017462f
C886 VP.n77 B 0.032545f
C887 VP.n78 B 0.03452f
C888 VP.n79 B 0.014139f
C889 VP.n80 B 0.017462f
C890 VP.n81 B 0.017462f
C891 VP.n82 B 0.017462f
C892 VP.n83 B 0.032545f
C893 VP.n84 B 0.032063f
C894 VP.n85 B 0.971763f
C895 VP.n86 B 0.049839f
.ends

